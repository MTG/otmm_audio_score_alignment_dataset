BZh91AY&SY�ɉ<�y_�pp���� ����a|_  �
� �  
U  P  @
��*@     P �@�$ �$�J�!
��UQ	 R����Jk%*��AUIP�(P�(T�J�J�     h (@   �w 2�&��F�����(=�m���택�������� pu�ޙǵ��T���x�]�
` �5�Znf��qeЭ8�u��+�p �êu��@��=QC�/cF���C@��z  �@� � ў�Tť�{t�[�*������Gs���s�ҽ��s��z Q�$�sǆ����	;�i�{�r�����[�y��3�ݵ�v�� 
�\�:czoy��;
�z�W�       f�M=�E��1����᜜�� )n�9=�93�W�Η�q�G8A�|�����s� 9�r�3�<�� 2}����s����e����=�ӏ
���s��fN��x��zQT ��  @   㺀<���g6�[��<�� G:O]G=�{���tU�׮�FO���8>��<c.�&#�� �}�&[��ɂY�]����@=��&,���evr���    >�  �� i�2}�.0�0n��gT�� ���X�J�/�9�{��>�����si��@"��R��L�����=�C�1��`��D� G�ۘ=�9���`�U       �z�M��U2�0Fz	� %0����)�2hё�1F���=UR�b`	� &L�تT�ISF�=FM  i�@�"���E6�R�@�  ��  ���T�2�e=OT�d�=4��O�'����k������l=���׾���EU�5p(���QQU?�EU�h�*���"����U]_��L""���?�@�*��L���O�U�ՈC���d���fF�5�Nlȫkn���cQ��Ti�n/�BWC�gM�؞&�5d���M���>R��<䫾[x�
���Q]7ǡ7��I�F;��č�t�	1�[^���6���nTR��ۻ����7�%��k���R�z�v|�ǐwW�>��[>pS=�����&���G,y��炥Ct�r�N"���q≯�p��mՍl���B��r�Ic&*��#_���`�A$Dg���7:��՜C��r��8-�|�7Rz��ӣV��,��t�}6U��%��٧������1��߹M�������x�k#/��L؁2#��;�x5���GB]kWJ'�TD�F4�b����E�D$����^q���wOw"�6�,�,C&4}�讜�)ԅ����}����>Z�E�p�i����������e���E) h6�&,�e���A��42���4�t���x��O5���ܖh5�5C��L_H��p�}ÞC�{XL���p��).){�2o3��Y˳�ۻ��^��\�vu^	}��{;���xZ�Z��9�9�ˊ�"��]��I���6��$�Y
5��$'�I<c��14�bvw=���H��#繯��j�lJ����j�	��+��$4cJ��D��8�{�&�愹nU��3�驏Fy2,�x��l�W��ӻZ��c!r�,!��8��ƐR��K��>Z[���.9�ڇA��قx�0X�MBNV�5;7:���'VAo�Ou$%��v�>}��s�k�j�3u=;����T�>�	q�>N6�c�a&ք�,5�}|�̹��lٹЛ��s�:�u�����'/gߺ9G����x��vz�!,&&]���ۺQ�zj��Y.�.cYE@Gc�+��/>"�H����hٸ�8�-w}�n"��{5ѩh�T�`�)�h}_RXl���ӓf�X����>�x�^',���S#����۹ڬ`��a
}ǈ_#LG�˾DQ���y1�g�Hh������9�)���sPT�"s���8�Ny�IA@�1�7���r<�eŎo�y�G�<M�c	Md.y}�����$o1I�̜Ӣ%G�i���%MK���%�Dh�!�\�u	YQCpN-@����]
{y�.mY�v�0r����XQc����)9Q�o0\�)8v8ϼ.�߹��U�߳o��SӜX�Q��u�W�^���I�&U�P� �
��}�#����?�Ͼ����`�1&	�S��������å �aA��Zj��#1�$@��N�s��ӯg���D*����A:W.'r��U��i'Glx�k�`9�N��qF8	�(@C����0OcY1��/;D�������8/���N���Լ��"eY^�k�3�ud�%��wM>�d����¬N���Hjy�<m\���M��,�d7r��f��9�%�c&"2��s�5�E�+��,F��붹��u���rU�}5�y	ף��hӮ������7ӛ7|uF5�ש�u$������~�������LM���|���X�1y��j1;VJj5�BZ-ۼ�^��z�|v��#�;ވ]�VDA"A
F��=�N[�㦩t����qn'(�qU}W�E��o7��y��,���z�շO5��E����DF�u)�eD]����&TV;�q��� 4ch�j��D$tTU<�:0�oxpOuj�/��|s$�7�1]��TX�,����!%�'�uW�4氂��y�,i�	P<������X�Q6�Ȧ	�%�X�ÝMb�%�<&p��"@�2�	$�uv����ÙŎ�&u8�L�eɛ ����c�Fc���O��J��(�U�ξ;����F��� �1�j���C�8��mŐ�
"��g>X��sv�|.:��%�RtYP08�s���)�0K�F$�X�V;���a޷��(Gx.!�=��^2Bs����;�^}uk���̀��B���h��>I�8�X�$�]:<�c!A4�Pਐ,�*d�z*#��4�PC֮���lv���歯�j<�ۭ��%����=��*wN��ّlN���|��ݼǥN�8�NQ������3ܞ�j�s��^F��U7-��.�E��~p�,�!8�����C�gP�^;��C�E^R�ђ^N��S�ιN��ESr^�]X��癜8����	�� ��8)w�U�N,j�X���,���$^��6������ ��sH�we�9�H��0��Gp�,)^#��d8G��%iJ�����'����$	�ț^$^���U�͛���6sϧ#+E�PA FSLHX��Lp2a�VuY��Ν��n���=�3|��'8^W���[(��kz6��8\�o*@�q<�ڟ�w�27�.(��>�Nw��n���<�'^���q��C�;��c5j��"����
�3����o��cn!�Տ��}�Z��I���D[��^ڽ�����,P�"HPR	{J\M�P*d��d	q���I�\�9�恵�w��"jy��}q�_h ���f�9�SA��OX���`B'���@fT�f6�	�!,H`�ҟ2�Z/eg19Ճ��ɘ�'pd�I^"Q�2"ޣ��ɼb^�D��m�%�{ۍ��+yy������u�o\�]��ޕI���"o���:j����!9��!�	�o���̻y<&��q���丶�	���{�����S���47i���1���)����'Rո�E
n+QP�B��������s���L|�|یW7:KLS����K���;4����Ny��%�%�����|��v��7X����J4��i���w�G�X��x�1�q3��ΠJDPl��tHG̺s���o����A��PcM,|�i0�&d"h��{h����Ӝۼ<v��ϛ��~��h��K1-���ދSӢ�������P����\����J�7@��tF�hr����Z'
�<�K�C��!�'E��ix��3�o�+�q��
dC�l���'yx�>�k�O5AAk�74�T�RrZ>ʳI�8��m[��CLh`�ŋ�y�4��������I��8#�<���t����L�v���"���t�c�u��6Q.����d��5���0CR�
�F�E4��#æ6�G�a�[�w�Z�.K�Hflճ0�Ih|�a������ٚT�!�(pvx��DY.;3��Pu&(�V�����1}��q9Ō���78��(2�p#'�}�����+tFE������h�ǔG���Į=(��Y/ER�M�V"��7�8��o���X�v���\����X2�nBdk>lK�	ۻ�ƱE�G!�c19,�I�	N=�#ࡺ�u6��=� x�!�pNY��'vڶt�,����[+������j|W�[��M�+/����/ܔ�l����8�O�����U�7"����h���;�o=���]:��?p���o*�����Yc�5h$�p��1�a�բ}Y	
L`��a,j�^Q*��d��&Q8�4�xjG+78�;L�)�x��{�d��)1��J��iρ�sx�(n�ϻ��l��1�O���{�<��KMV�1���*B*������jsO��(�jA�h�e:`�K���Z!'1���g<�(K<H���&&S��Ba�&sZ�fD\"q�	4����h�6�H,���`K�@aBQ�d�	�C�����l�+
)�`�
�}}�F滘���[�dϦ�|��� 4e��b�N�iW�&0������H�1;���ھ�G2b�F�O��E�3U|s��n�C�3n]%��
�3&q`>�a�P�k��ʘ	�"��r���\U !��"ĝ\�}w��/N��Z���'3�T�N�"n�r���,b�	�&�p�d�aa��F�ki�R:���w�y�h�P�Y�l�q�'㚇�>���\�CPO��;���78��V]hh[��ē�t���|����W��L.�ߑ�o1˝�O&Su��$J4�����*B��]���_Q�ND�6�/Ӽ7'uނ|^��[����{:滯^�v�ן"��3��m德b�bF�f|�N9��w���W�z�"#��^;2�N�s��%*�	�L�����9���S�U���s\���5��7��Ӽ�s�:;��4>�	�`�1LD�D<���Ê�.g���ֵ�WDj������9�;���������<H;��!$т`�K��k̈�d\ȶ�p�	9T�>S��9;��F	�(�g�b�nu��&��X�1��x�#]�yv�2H�W:Vƻ/���aqg��Q�if4;_<}ׄ�¼!��yĐ!�8���d�g���4+#	�f��E	ܩ�5QQ�lbH,�:��,=C���bi�,!y�ST��C���/3�
SC��İ����(42$0��I���顣���9�'�⒧��,k�������h�ߵ��������YA!�b"�k��J�9�S��#�!«]Q��D�SDsdM2�mB�N�P���#y��$W4�����u1t�	ƚ�iN=F�	G�B>��	��s�g3����2����:�	��#��8���i(�.)w=�w�㽓׻�}�F	%�����Է��Q:'��Y˩��4�����Ƕ����.%V=������r<�˯[�l8�S�$�Las���y�}o2!�~Y׽��vBU���*��ѵ��t�]��gG����%��{�?g"����j=P�]�Xs��=ǘ�e:�hwP浚	�u���¶qc#(#! R�j�V	��x�XsR�,�؞�M�;.O|��f���Ic>QW�z��۾�M"f$�@V4��1����,����a�ַ�O�^q=�*�][���˻:��ϻ���F|U������ϸ��o��׻��t�Ӛ���58�>�4�9�<����;����d�퓜';�7��}i�/{��<����@<�\��X�T�N��M�ﶎ��ʤ��}��D��Q�̉������I1�9�0Hɋ����bK���s�����1�ӉB���Ӈ�w(ʆB��SV�!	��ōM��_��#y�9��0DF�gQ�C "�	 �y3q�O��^��g��Q��V��(D08����&.��(�N|�vh��%��{ε����o��'~�:y��ξ#xkB�9V��r]�k�����sm����No����|s��B��;�q������C�&)\@�P�L�$5��K�Ά�c,�6�P�/�Lփ�%	BR����w���)��g=��W;�w�¡��,S�|��<��(�ث\�>���ʕ�y���y��V�����F���k��$'~�s^n��������]Hŉ$�}�r^��`���qjX�?c�,]�y_wp��gxro<��|�C����qH'$n25��'�]�]۝dXt��Pi!��_x}�<Sx��[uM֖�xNo���mb(����˗�7�!7���l�p�>F4�aV0Y��L��s("H
>�z�upz��W��W�q2xN]DJ�".^j�|�q}y�w��ya�@�P���a!t�ӈ��3��$c�i���y��|�[��H7'u{��5hąǻ��so�ǋ�"^�O�Ḙ���N�m�h�,[�*c�_U�f4�#��sNHC&D��Zy�|�wrs�{�.�cO���YkM�����RE��o��w�'��������>�| 3�@�  k �m#l �`�8f� � �Jr�.�   �s�H  ��   -���    6  �n�ؗ2��&8J�/ �햪+ U� �sF'��T��ўV��+��8}�Umr9�Y�P�6�'ju�-��:��hc��\��3�5*�*�����X�,�n@�l�kv����e��^�tAm,�VI^Z�*��6�:�$��3�ݑ��� �ݱ�����5�[6UUR�����5�k;p�R/C����r:��q�^St�x.�F���u<��z�MdC�mp�;�Hri�����-�m��;(���m��-�)�ݻU�\�k�����mv��u\���fz;:d&�v7%7T���b=��챤
�T���A��f�k��%�`:�t�v��Oe0�v[UƏ-+�5,m�&��f�.V�h���3����jՎs;h��n��t��uv��Ɓ�ا���p���d�ٕ9�msT�T�mI�p 6)0�����WLAt�YGvJ�U�^�jzR;#9�lṝ4�3�{ioI�nҳ��r�/.�:+k���k�!=�۰#QvU�%)��K�[Um=�(7m��(݃�Q�t�[p� A�-�&��̃�!��gQ�Z�HqP����gl�F.i��� ��������6��Mw+͹5�R��r�ɻo-c� gY�4[t�mo�t�X�9�z�kq�G#����v�7jhqs�ҽ�u���zZT˺� ����W�R�*������V
�*q�0#�o- �X��<�+6�kj�y@j����U+�uScp�rC����ŷ���
���<ۮ�}��ĊP�F���t�Z�m�D�f���դ�\�l��	a:xkp6�ѐ��N��m�m�D9T��g<O��3�p8��mm+�z����W*���[���im�Z�aX
S�uJ�r��WD����v�P�j�]�T�6,u��r���nv�rv��g�=����B1�xƚ}W���� �����'����.ָ�)�ծ�d�Kuu@uV(��l����q�6�R�T�pᶶ�����H�ā��&�cH�$^�W�I�< ���A�nA���6�8m�,�-��� BꪪU�u����}�}��nI_>��Z�����Tq�4�WPcւ&U�eWʪ�@UQ@p�-�mnM��t��ݷU�!)ې�Jڪ���̊��y�Kn�0m�6�s[v ��;��[Zk5�A[US(�ꝹP(�����Gg�(��`��`sv�u]�j�7�Q��k/odwk�n��s�������\fAS���럁��e��k7j�mbTr�t�;��
���w%n[u��\�e�m>�~(/�����d�;u����˦��҄�=��d)�`�ۮ���T��6��#nBQ7��� pJNL�m��!i2BFf�i��JD�����!&ݵ���qv�A�}�W��*�Tq�:M�@evj��s��!� D��\���<��H�'Z�_���'>�.L>@����_D��0X��=�b�`���]�n�4���͔��R�UU��ҨiB@q�M�u��K�^{��̎	��yx7=�r����\�UQEW*��n�}
�Mb]��M�`h��`�v�6���H�-�Hf���m�m� �K'Ygv��m��`��v�����>��9���Q�T l�@�*ܭ�PUR�����-����m�6��e��� I�֞�Զ�e��E��Vô�@-��
[vۮ���i�q��Ή�"�;���m�'-M�=�5l�z��6:�l]&N�v���\[��j�����6�'kغ��n��]f0�����*�r��	��<\90�3�yb���t]�v���:�==n�knB�ϻ<�n�l�f�V��q֘�IݜJ�[Ai��i�t:cN��fu��gC�$<�{M�h3�G�N�l�;b��˶�W��u�m�^-ѓ7=n�::U��K�6�<�3gȅ[R\MB�((-����.ы��m����wi+9���g`��j��7W!Idո��9�g�y�;[uVm`؛Xv;0tmr��N�xڰ0�۔����Uq��Ղ%�B��N�r�Լ���6���ռ��1�̪�@mX����eyj�v�j�}�R�q��.�f�=�]���(�<¦�<om�j�Y��	�㙝��퍁]�]� j��ݡ6Ն�פ�
�[*pK����We�UZ\�}�ζ�떺�Z�(�%�����։l��mD#<�t]J�G�5��cxv�i6�]sͣ�U�n�i�����r� �Իo��vz�z�v�n��^C8lb��qUUG� Slq۷
��6�݀U� ;!�6�資M�9i�����5*�[[��d��˴���K�l�!0����I�WH$�bu�����z�7�]un��X��[ַ)���r�
��UV�Z@7e��ު8�����r�`(�
��Br��u9j4mٶ�:v�[@��8��gV�\g.��]�j�[Q���J���L����Q��g^ܑ��	֖�Y��	[mcZ��p��PG���!��"ͺ���%Z��y�e^���j�yzPݚ�
��N��kqĠ6��B�v4nԯ	X�kn�i4���pj��W"Q�nb��@N��i-�n��U����lqƞ���3pGWS(��9Z�@:Bmrf��T�r�svdܯe�;r �!uR�v��8(*�E��y��ĩ����um�"�ؒ�Ȭ���YP��������tXH8��m6�VݯV�b��΋:���	��I���]��W*��t���c���ᶵ[2��]5�mlOJn�.C�iRp���J��x�V�`�,jWg��غ�̆M�۠=6��-r����U�sb�^�H�]����Ȑ$-i4�6Zl]Z�V�N݆�� �U���.z��m;�G���V�uV�1!2�W���e..���(n�{f��K�%�Ԝ�i����W��t+��;UJ�[1����lq�n���&4��Y����E�[veo6�U�hHm=W \�%n�VYe�%�"$6��	=U�6Ͳe���۰-�-���`*�h�;[�� ��Q�8��nݸ'UR� p� �v�HI\�^Q�n�9����v����k̀�l��||	��m��$�9�J�{Z��L�%�4�UUTgPX�]c������<��I��,��*��]c禚����C�����ݮ`�j����h¹�x�%�ܑ�m�ލp$9��Q�,�2k���㦪�-m	����l3N�V���
��
����}¿UQ�m[  rN9��jAK�ɲՆ�ʭuUR�媪�eN*��VHֵ۳V��R���  �I�nYv��j���^۶Z�V�h��[���`pn�	��ZU�ey�
�Z�̞m�������q!��.�F��[Ms֥��؊�r� �Si�UP�煪��-�ml�\���'sm#�$�p�]�)-�6㚫�R8j���nÙ+j@l�28p�  P��h�����P۱UA�ekj�Z���<�a�Ą�����WuJܹ��E�N�^^\k%�$�\Ը���S��|�y��`� �U�
��]���j�J�c=�uѩ�Bw/]�W!Wm�N	ieUCa���� m����0my���8H6Zc������q���6�&��V�A�)�Q�[��	jr�UuYFܤ�c�r�k��.��;��.j1%���)(R@l�iT�=�4pP��j�e��p �UUҒ�M�����W��W��Od���k�졬1�hl�=�8��P���\�XU�����6Ϧg=���[\�&�<�	H��η���be�zj{.H�N|u�>;�&��"D�u���g;^�iyI�Q1 -�ک"K��YV�m�ݦ��� Gm,��k�+khGƙ�g���͞ʽp�ۡz �이�v��[�PRI&s�bV�eݔ���f�1��N��~��gc�Oۘ�b��]�+6��V�L�"� ��k3�ְմ��-����
�6*�[��ɍ�-r�#n���nuҶ�Zvu����&V���t�˲��c�Uj���J�vx`:�c"��9����^UU�mڣ�ڍK����Z�]�����l ��C�H*�R���A���va Hp�M��m�N�[v�9��t�f�i m�6^��j���=J��4P [v�l�sm�Hm�LH���%皪��6�b3����k�6�5��M�FC���l ��+���_-@TVP�4u�Z�hM+hֲ�+��5i$��UU*�l;T��.e��1M�,��Be[˵�����,����Ҭڪ��b8B���l��]�6*�������m�[Uu���U~���,�UPj��	�����PI�n۰ �22�����*���ԙ��zƌL���˓m�V�2�ь����UO0l=jݶݔ:��9v��UV�Z�$��F�Nlِ;��k�B��<��,"jW�O+t�P��f�v�K���^A�V��J	ס��`�m�u�!�R���h���Wi$Ma��5	�\D�����95@�n5�`��.ve]��B���n����W���h[�Ŷ@ $��\�ۃl'��Ǐ�
U垇mG	(@[/2ù��*e��+N˖uS� ���`!��Gl�Al�mS` ���n�UUI���}�㴫�ّQ��OuWPJ�کsl�ؖ�k�KF��M"�}U�R�������㢝�e����y����*����iUs������{����@p���> �d�|T�   ��lH� hC���B��Ȃ��c� ��|aQS�m$GH���S\O���>mA�x��A�A���� �Fx �8��LC2EHs!> }BP��H Ї6��� ��`�OAQ�N�,H�ȑ�� ��'�#�BA�⏃�,��?	�>?AU~�$2A!�Mq��z�U`>�'� jj�]>*�EH�"��~"�h���}@ӄ����&��$�J��W�#�OW�*�X8}P8���,��P�C��W����G�E_��J a�<	C���H߈:�'��1G�iF=�������]'�҉�W�8 �Q�H�~p O�}~
�TE�4���d#,d-#�)q�"'�_���B�)E� VRDq�>��)���XBM�E�(Ĵ�
��PM2��HH�D�JSS(Ġ�%R�D��_]",H�/��Y ��G��⫩�Z
�H9�`�)DH�Rd*�)KJ��.� ��2(�Ax�ϿbP��%(P�fb`�M
����	�$�@����"�*"H��fG���"�
�K �nE� (������)*�"��� ��� x���])hGi�"?��EU�;�_��>��G�[�?�D̰�'���HI�(�MF��ޝ��A��S(	B�Cc�4�H��@����{�W�?����}�<�\��l��N[K��Ŵp���n�ս��:�ܙ��m���G=s�F�+v�s.ݫ'��6��%����q�����|��-��ԡ���^vLfu�@ܚz����;gSe�n]�e�&+j5;0�;OJH�g���c,�nn6!�`�5�Fyy�S9��ƴq�n�|k�t�9;5i�5Phʬ��LR���jLX67'c��Y�ܝ�� �/C�(��:uF-U�n���Zi9�M���8l؍-��ͪ��z�;i�'	�,6�m\�+NG�f%3���cpWy�z�Z����T�/F�4X8�9��m�y1L�]�� ҇ 6�T�mX�jݴY�K6�g�SN�m�)5�1�r�A�e�<������Y��62�s��쬱�kՕ��bS�+Ƨ�DX�#�qt�ՓI��!bY�ն�H'-�:�JN,����#.�l9�l�&�xq��"z6�E���l��Gh8�\�� ���x)ӶzU�\��M��^A�מI��V.K���9���Yƞ�h�2<�lc�CQ��ݞ1�:[+/1�9�H���6��1ۧ�.c�����v���oX������֭�۠Cfq�vm�kxyŷI��8�:v�5����=�c��d乺�^�3��]��>#��xl�ŒgP�d1=reVU�a��nm�1�I05�V#r&v���3��OX�̐F��lF��i˃;6Da6�u8�s���6���vM��ri�$������
v�i�Hףr��>,�9N�cn<<��y�[2nM�zv��n9ܝ�{n�gj�"Гγ�u��u�^{�ŉ{:��Ơ�H�u<Í�/��;8$����ׂ͸��:����S,������a��9s(hCGf��(6�0���k3����o��)�2[��rP8ڝ�*���̰��n��o�8�b�b�V��c�2��a��G����P��s63㭼�wف�w�Oaګm�]�v����,"OY2�!F��6�NZ�� ����30��� �����_�Q8���8�����&�OE$}>�@ڼS��1�>i|�u�v�!cvVzSK/^�h���L:J��UN'7G0Yj��C��q��\�p�/=���뭫v%�v��nٶwA����S�mݰ��>:$9y��qI\��l��-����u:
ឝb�U�׹�g;�vݺ�8��í��"�0`ܥi�ݝ�n)�G-��D8�pu�si�e]�:�y]�;���c��m��S=�s�uƥI'Il������s0�9�p�)x�ڃY"JLL7=�>^�6rxE�`��&'��-E]�{�%�zT�������A:8`tܶ��)�n�� �w<��X�ό~��oX��v���7cm���X�ό~���s�>\�z�:��j��ʶ�`w>0��� {�� ��vV��sbM4+Wv�Ҷ`��, ������������̠?*��O���8mY��vq�cKX:�����ݮ���vw8. ò䘄;�M����e�� {�� ��vV�s� ߯�`�O�+i5mڣ+��K���o�#�ɂ�fE�:~������~� =����v���V�n��M��s� ߯ܰ��x����ur�l�uc�E	�`��,�����t���K�d0�;��e�P���V�X�w<~�e`�|`���?W�D����.��M�wd �m�{u��,��s��]�.n��mWRNqBʐ�%RƲQ+b��ė}��5%����_�`���\�z�:n�T�M��u�}���7�>0��x����_��$E�)n�Ƅ'bcJـ}��nU}���Q2LFEbe����\�ŕdi`Hp��_e`w>0��w4�n�t�ڵwl�{����+ ���o�|`�]��bj۱Ҧ��~�e`w>0w�i�%�}�Ԓ;���L�p�Pj�ql팓�F��Z����/�����]>9�"�n���j���$�`w>0�ό ����{���u
�_Z�������0�ݕ��UW䃺G�}�X�ό��Ϋ���趭�m� {�� ���'ꪤ�#���� ޲�W:�h�Гv6��=��+ ���o_�`}� F,��1*�o�R]6xZ��*lcn������ {�� ���MI.����H�j�e�r1���R!�vm������ӍZD��NrJ�լ:�X	��b�`�ܰ��x�s�V�����E�[���jݳ =��}�>0������|�f"���*j��7�|`u�,'��p�� Ww���B�cwv�l�p�(�;nx����fe���� =�]����M]+m`}���>��X�ό޾�W��F�ʁqtU��NS�Uͺץ���M�g�Ft�]�Z��.�=��='��z�h��m�Z�-�n]�N;
C��a��Q��a��lM������:�i1p]��@�W3�v�]���̑b�^�-g�۸I�urn^�[���r��	���sh�i�q�ڑ;��Iͱݤ�7@$g���u�9#�*�p��v�R�BnK��[�T��aS�{���}�n�;>��ð���g$��_Ã��;�V�7!&�&��CL��M˫WmZcn�m֤�K�`�>0�}� ���}e�ն�	7UUW<����L��nx�� �+�:��g͐JQ@E��U�/w��ԗ~���>��,��j���T��U�3VpD$��o��y�9�}�� ����7�\��Wn��E��v���À}�^=�� ��8�
#Ա~�֭ޭ�K��ۋc3oV�<;uU�]�,�]yp�����$�ڮaWd��p�^��q�vA�p���l�n�&ـw��d���x6�߄̈!9Dƌ�@��*WuTDBE��� �v���xq��C�˹wuo��TRV��=��w��}�>0��,�u4��!60Mݵwl��_��N�ގ�}� ���z�:��m�;������}���>�ݕ�{���>��������GK�,t�t�9[kRKӎ��'M�"az��8ޝ�l�6r��#���U�Z�%Z���_����=���7�|`�rW�Lt��m�l�>�ό�ό~������g���nմ15wl�=����/��"!TW�/�����W��?'j�m��Wl�7�|`u�,���=�|`wyYg[m]���m�{��y�w��o���=�}1�U$��W	�V��;LӤ����T��]-���+q\�nV��s'n����X{��ό�ό�uv��lt&ݵj��;���T���/ �0���#r����v4�0/Ix{��s� �s� ߯����閏����;���>���*����`�C�l�*$7�=�`��Z�E4]64ـ}��� �(x�΁����f^��9wS$���]bp$�s�;]EŻx7k�5ش!y���泖��9��%m����}� �s� ���,z�ԟ;�m�&�ـo�ܰ������X�ό ��VZ��[��V+m`u�,�ܰw>0��� {�߮������E%m��ܰ�|`��,����uGV+_������f^�Vd�̼8�fqp
�P�������>T�A�I%�T�r�깛#��@u��J1�K�1���d��s��\��F���=�lKě��;e�g�������Z׋���u�6:�v�ٍ�yN3r��۵s�]���;k�{.^u1O��;�o�f�^��["Cѐcb^���{d�.Cl�dȥ��//�ɘ;��7/��r��P�K�޽\��	�`�1��6�SQ(R�E)ZB--T��ޙ��,'����j���WQ�SesF8����J���v�.�t�x;\q<LZ�Z���n��6�c���� ��"�;��}����ό﯒���tƏɍX�w>0�>0�>0���޾�/��:)�鱦����;���=��{�u�]���ue�wl�3�xp��Ɍ�{8��+�/�}%`����c�+y_|����we}�s��wvW��0�Xm��&r�����L=�o�ݬ]��ݵ�̝�V�y]�.KRN^�r��fq}�e��ff�Q�������U9��յ�n[�{��f`�@1	�6��=��|����t���~���Ckꝅ-v�eY����:���>��}����f��_C�ʝ�V:����ʌ�����#338��reRʫV\I6\��]Fffq}�e����_fT8�f.·�m��ѼHq��ld���7h���v��N�vg�=�m�\�-��<֖�w����UWwwe|}����+|�]}v�`պ�ڪ�K=��q	A���<m�}�e���ג:Ȩnݶ1�����w�ݟ����r<h5&o�5jJ��=�i�D4������A�:@�;��Ɵ�s�k)h��>I�J "J֓�|�	�tRg���t�	������6#�Ė$�`�$���cf8�8%��h!�I��_S�p���.�/4l��`������aʏp�napO'�q������79�mw�
�<}�qf�"�>��|}��|�<O���8{�R�L�>9��:u$�¤���wp�����Z��X�70;��f�>!%L3	)>$��L$n�C^���������$�XLG�U��
�Y���ŭ�k�y�8y�d��di1&�=�0m`o�s��p�fU�3�x�D"��_������_ �Q�}D�T|E����QC30SpTS�� �����W��}��
d� �O{��R�������)vﺊ3��ؤ+"rٹ�Y�F~��ߴ�,JS�w���);����JȀBN���B�
=�AMV�ͫ*n���9������{�)JRw�{��������({���JS�{w�����{+�vݺ���F��{n�n�\{`���{=��Z��sy��e���3�~��JRw���%)O����({�{�'�JR�s��k�R��;ذ�����qf�z����|��>��\R���}�x>JR�3��\R���}�x>JK0����~��U�%J�,��,�#?w���JS�{��R'{����D/Nc�D �A	�uE2e]�.iU�3��8>JP��=�u�)JN����JS�{�u�(I���� L`ӣt0���	�TT��0O Z�~�%)Os���ֳu���Z޷��R���{���$B[�7��F���(��2�g�؀�/��۴�=0�nw�ι�7�Y9�X�#��kv�{\����h1}�V*�z����>��\R���}�x>JR�=�y�iJN�����)|��j����Y��Vk{��({�{��)����R���}�x>JR�s�{�
�$g~�����G,�n�Ř%���8�)I����|���=��┥{�{��R��ޙ�s\�����[��z���
�����JS����R�=���JW�{�qJR��}�����[q��ۦqf	f?��70R�~%����p~JR�~��)JRw���%)OO�Xpa������A��& eZ��9H�g��:�6EnY���r�iLf{8`��>��l\�tH�n��֒�b
�ώ���*
E�ݮ2��Wh�a�/9�\[l\;7C]��N,蝒鱳�:���c��Z8�L�!u�3ko`��5�WKn�����o�-йA��l��m��7��-�࡙����l.vMЙ�]��uѥ]`�;�b�A]/Zn�~�fa�����$��8B*D�y"����ɈhuA���YIbuŹx�ݲ�M�*���l�Z6oY���)J߾����R���w��)JN�����)�{�u�+0K߾�"��e���Yvm��qf	b|�wۀҔ��{���������
m�GD�"�B�N�ʹ�RU��Y�K�$BZ�w�:D �N[��%?�!����߸>JR�{��)JV����ʢ��B�.�Ř%�y��u�)J�����)����j��t�A���I��SuJ�Q5{��({���J�?{���)JR~����%)O����)?.�~��'<om�E��[ ��D5=vi�u��)�\cW5�7a�+�۟��~����kz0��s��)����);����JS�w���B�����`�a��?����Z:EevJ�0K0����� � ��4�:�+�Q�37��R�=�����)J{��� 9)I�;�����nf�z޷��|��;��~��({�����Os�)I����%)O��&��JA*��$���3��w�%)Os��\R������%)��m�"D ��P�L�Ys%+��s{��JS�u���({�{��������({�{�����������{�����V����xy��[r�{��ֹm�����y������l��m���)JR~��߸>JR�{�{�R��6�	t�A�|�r!B[��UUasVIJɫꏈ�6��H"
�����)�}�u�)JN�����f%�#��Gs��K!Yv���({�{���������|Ԩ�,�JFS�a��#1	��ւӎb6�@Ӂ`�J�bx8�'����)Jw���(����n)�����%��8��<���┥'}�{��R���]�qJD�|Q�!B��|�V���Z����oz┥'}�{��R�>}��qJR�����|��>��{�)JR~@{�~�{��g�˻!B;8;���F�<���k���0u�p�햲��n�}�G��y���R���~�)JP��{����ߺ���������%)O���
R��Aa*욫��B�
6������䧾뿳�R���������Ϻ�s��R�����Wvfn��F��k��8>JR�~����);�{��+J|���8�)I�{��%)O��')�+����*躺�B�Bx��|��>�})I�{��%(>
��v�$�S5�!	�X,t_ �G� �s�k�R������?ZK%�N]3�0K0���縔����a�R��;�u�)J���"D-�����Q7ET��Ƹz{=��=�Z;)�ݐu��=i��d՝�g�S��g3 -R4��嶕�'k��,�~��|��>���8�)I�{���R����┥Ͼ���k��Fh��a����)J{���JRw���%)O��{�R��������a���~�R7%#%��k��,�,;�{�������)O�L��~ފ:D �M���!B]��s5eٸ��o[�����)�����)JN����)J{�]�qJ� 䟻��������Z3��a[�5�[ַ�R��������B����┥'������)�����)JN�EH�X
@j������h�oz����k���N�V�g%�uh�{m����Kg[���uU��3s��!��7p�ι�d4w۫������cZ�N�c���=p�Ny��e�!�9�n��D�Xul�����}�@���*����x��W�4q;�zOf8�P��e�`�Yx :��͑;i���.���'�kl�.��sd���uA����0��f�UH���<`%||v�0q��[�s�����7l-���@W���gͺ�V��w����\���֎z�_���)J~��g�);�{���������);�{���)�ze�wz7���kuf����R������R��{�)JRw��}��JS�� *!.�9�%՗wv*&��:D �/����JR�����>H��}�(!<m�GH���JT���^��o|R���I���o�>JR�{��8�)I�{��|��/����JFw��G'��e��uŘ%�w�ÊR������JR����"��:D �^m̈\(*�eQT�
�� �ۭ�x�nو��Ʉ�p[��lO`VE]qT��[%��	f	a��߿i�JR��}���)I�}���)��i��Y�Xs�Gib(���m�<��/����Sݿ~(i�P!�'y��q\h�8�A	�l*Q��'|��%)O���8�)I߽�x>Bҟ>�Z3�7�o,5�����JR�����%)O���R������%)K��|R��?d��jf�XXR�.�t�Af>R������%)K��|R��O1�t�A�qH��+����	����)JRw�{������{�)JRw�{���)��{�┥'ϵ�s�n���ڷ�i�^�`kc�6��^ݵ����]�*�؍{d!�Ж���is�|��?6}�o�R������C�)��w��)JN�����)��V��Q�e++n[��Y�X~����Ř)O���)JRw���%)K��|Q,�#>���&��#�d�cr�8�)��w��)JN����� x�3
�eP�L�BTp�p�@�p�/{߻┥'~��}�Ř%�~��ȗ�L�r�c��`�`$������)}���R�����a�R�>{��8�)I�b�[ٽo����淾�����{�)JP'}���>JR��׽�)JRw�{�������~�w�;-���n͛=c��=�d8fspZv�ú$��	حV6��3,�5��{�ލ��{┥'}���>JR���{�R������@<��/������������)QY��wQ�Y�Y�=M�Z(��!-ǻ�"D#5��JR��}����J{��w]޳y�-kyZֵ��qJR��}�x>JR�����J(0�I�����|��;�~���ß����T�v�,jIt�,J/���┥'~���%)O~��)Bk��A�\@���J~4�PM�z|�>~��%)K�n�T�j���\�����B����y)@~T�;��~�)JR~���p|��/���┥'�~�TA�]�ѻ[|���Ӌlv{nF�v���g��J����]l�.��),I�6Gj$�cv�8��=���qJR�����|��/����B_fV9Q�!Bm�4��QtM�{��{8�)I���$
R��{�)JR|�������{�Q�ÿ�!}?%iecn�k��Y�Y����|R�����{�!P)O~��8�)I����%)O�}ٖ���vo+z�[޷�)K�Y2O}���JS����R��}�{��R��1	Nk��B����ڙV��UU�^����JS߽�n)JQ�$O������R�����┥'߾����)Jw��{����h��3X�t��S�1,�L�Q`ks#��u1F�ԯ"(�B ԯ<����+o�s��Cl)��푯$&}���<s�\(��k12_��ь����&x������6!�"��>6l�w��CR���\q���Q{���Q�ςl,!9>�>-�Q������>b��8a��c�s�7����&�YVŕ����c���i")ل�3[ѥKBm܄oG��Nc`T�m�O�>C�9`QCy|��9��&BF���Ey�Ya�j5��X)���7A,À�ӊ���4PG�p�,���D!�b��
��0�M@a������~^����?*1mR�؄
�'"�r��s���u�R b�i[$;$I5�F\�<C�ŷ4�bS)����l��:���':�n��s�!A�4:K=r���c�����j6�<O����`>��:���xq��\ێ̘̪>j�wO9y��O;Sv.�i9�@I�e�ayポ�DG�"�&��Y8Kϵ�c����Ɣi!����us��8#r�wٲ5��\��g�� ���ʸ�ifut;]���C�x&�v�d�la��Qeĝ����7lr�r���7/�����$�1�g��HG��݁Q�Dn9A5(�A[TLr�l�Ɯ���99����vț��qƅ��gt�i�-�:�l�e���l���	5��ۂ��93O�۱�ޅرlnݑ���]���c�7n��6uJ�,nԫS4<e�E5q�.���u����
�l�B�7n�m��۳'O���Q<�uWW.�is������].�٭&�C��N��g,�#��- rK���M�����X^�zJ�ZZfv!`�(�-��!�X�8�z{7;b��2�a��I�����S`���d0�e�6|/��乗:�rm$���gmt��U[$m��n�7Gh��4������ay8W3C\b�%��ږn�{Ue�����2<c�74����tn�{'��,��P�vH�:�'ٖ������q�j�7d���e����]�Al�"�k���+Шp�՗������6Ի�3���eۗBq%!�*勠�v7�� ���r�]��bq9����91���X����[cce÷����ym�T8�.5�������#��u�B���L�����v��c�(����H15k�Z$.4�t���[v�Ƕg�1<�U����VR'��qvq����mg6�.қ� K��s���ڃ�^W:�������޺�V�=-=k�f����tm�+��
a7bĉ��%j��*�c/�ve[�h��Ʈ�l�''NG (=�J�rK��U�6띱;+pn�Avnњbsp%���M ~���@=E=�|4Q4������}�DOD1AT@~ �Q����o_�<r�+rn�C�NF݅�g�������7���[ќx�N��gU��x��$`�b�,v���	��5�[�q��`]U��;v��gj���,6�r�����'e�D�ol��v�\�P��e0Xy�l@9��B`��..�صn�r����
��3���2����c�8�TR�<����{����u��Q��[Q$+D�:�A����W���Rw�������Ø9|q����;Vy�;gb�Ɓ怹�\��C�wu}Ɵ���h-kZַqJR�������)�����)JO�}׽�<��=���┥'���VsusWrR�j���B��X�?�L�����`�)Jw���qJP!w|Q�"!	)�]�7Jo8�)I��u�p|��=���8�?�I��~���R�����8�)C�c�IT:خ�T�|�J��!Fz��)JRy�{���������i=�X�GH�	�
�]TZ�n���┥'�����)B;�{�R������>JR���}��)I���wy��m�vv�m�8�4k����[x$Ә��D����W*������Zt����~%)O�׽�)H]���o*�����R�w���EJv�\ͩWW7uW<������vo�&@p�B � ��qE-s���]���@��9��㝝�	V�����h�,{��?P}/��'��h�"\e����.�յ����&�u�x�|gCbb�ݞ��U�˶�n��˷���XUS�8h�`�M�=:`R����-]Ю����wl�팘�u�<]�/KA[����v��ny_����^Z��Ʈ��[X�L��޸�?c}Ԓ�DB_�Og��Ҫ���ʙ��p��nx�@<���<����ΉB���ɻ��E���M�����:�<>Y򈪈P���!)o��:��<���UwArww7wކ����	f����y�@�Ss��
���{�r*R��ڕm�ݵ�w��UUU{�|`�tK��qi\aeU��%e:�)XS�a�=���n�Z��uӭi��VH18�H�q��S� ����*tc�N�a�w�E�N�n��X� <o���H��v����Gwj��'I7J�����,t��}W�����l�n���ot�� �3�D@g���6�������خj�b�xP��{�Ӡ<w��]���W�		,
~qT��W�^o���]����֭���jT���@�e��j��%���>�O�`��h!2��ջue� �iU��E��Q+�th��Eb�mD�Kh���d�0��U���X�n���&�K����GP�p瀖�W@+WwW7wށ�s�!B�R�y�@x�N �ފ��Y2�K�\�rw-�k �&C@�s�ꪪ'I7@�^9��.]�J����������
!,�8`���}/����'I��;�D�w6�������� ��@ԔA	G��� ���=��tJ	��	A�ß�|���N�\�V!5+MJ��>���AD%�6�cu.O!�i�r��V�)���yۗWk�b�J��M\&v�H��j�t��zxSF<u��3ɊƍYkq�F���pg����p8�}�ηKe�uӱ=�t���:�k��L�u��9m����V;%�iJ�2��c�����h�y�x�Ӌ�����-x.�=�=vSD�a�̹��+��(��������7�n!�B�J�BA�7ulqtL�ΰ��jm�I
*��r������ҩ���m]\��*�������|g@�e�+�P�&�����Jlӿ֭�{�C@�t��'�M�>��g����aj��?:bwI+y���镀Ot������� ���$�P�e��*�m��0?Q=�n���� ���+�{�0�(]Dn��C��n�{�}/���(Q0�����;Ӏ?c}�������d�y1�n�n//cA���D�y���w���[�������v>�D��&���'�d4�r,{�ڪ�=��	�q�*��ջI��hz�X�#�"%B�ym��fV9�����Q�TD��&���\����.��x����{Վx	1��Ss�3�N�v7n�U������t�wL���_E������n�}AҬ,��	����w�N��>��	�&�.�x��������'qZ�n6�u(,)����M:�����ں�u�1es[s����gdA�Wt�f��:�X�?6��>��\�����P�^��ʶ�I[X�o���>��\��>��<J!E���E��vݷ�˺^�{�v��J$<�P��eD��B�<�EZ����>�I���V
:i �vդ��~������s�6��"��Η�Ot���T�V�+��hu�\ J�x��@�sp��:�B�����������-��ւ�v�O<�wI]ͱs��ʓI�X�X����T�U�ww{�>��\�|d%
:���J +�c��v
��{�|����@<��t�X�?6��S�Hy;4l�j�T�� �{�:ެk��Q=�n���v��c��L�_8t��X�?c}�Nc�**x�>�l�}�y��~�,�����)��J��'�M�>^�x�c��z�� ؅k���
�M]M��vA��`y�i���+9
��V�%��r<�\쳗��`�`�֣U�e�Kw�/?�&�l��Z޾�?W�;����
:b�t;jӷx��kJ�߃�_E�w{z��u�I$BQ!�����%؄U[�I7��{�,��7J���t�d�k@��K��0�ci�k����7@�{��'M��_E�w���Q�vݶЩ�ot��^ ~���N�^U���r�}��|�Y��#��~1��7�aKQk��qұ�*��c��R�f��'��VG��.q)����^�ݡ���Z���@����d�U��s��
��k��Ξ�����#�vQ.����K:�k�:rm�i�������s��=���kQ�c���:x`��s�F��B�q�c�8��c-�ĭ�(F�^&޹�qxD|�e@�k
lEO\�����g9��l�:T�m�U%-Ma���fcԩ����(gn,�[=�v�Z�+��k��S�ny��d�d9g��H��{��|�o��t���ۼ��M� ��j�V���K��K�E�l@�%o+@����
 �{!G��{\sw�wRJdǳsFͪ���uw3Ug �{��Nd�߫�=�!�w�� ޮ�����vۻot
�_��tx�L����Q��N��ށ�ZUL�ڲPZ.�J�����Dg�������?�R^���~	��X��U��܀��7�[0�Iu��y:�v�Y��qX�3�Y�1�[����m��}=�n�}�W��_����'�.������e�v�U߾��x{��b�b��D��<S��m>�z8sb`�1t��Z@������@����|�}��ެsȈ���JL��jn��ITU_z��� ���鰒I
Q&e=���{���jA��WUu7H��� ����z�� y���(Q}� =�v��؁�$��޼s��""c|���|��s�<��B̈́��UE2B,�T�LC�o��l�[��/���|s9���`�lO`�ww��$K��Gkڮn�f�x��ހ}�w���)$�t�}�\WQ����;m�ot��� ~v���X�?c}��%)DB�l�"v�H�����n;ݞ���;��G611U~����7��2q�
4qЛ8�{Q��`i�(p�0�?P��U���. �M}��.�%2	C7�؈$���N�)06F��kϵ�o�Me�}���)�����ּ�xf�:52Y+�cI���m�hs1�ur��9��l�;u�LX�bJ$�����<�����^f��!����!gϾ|��N�b��B@�$K8�R��l/Lˑ�̊bJ0�$4���bD�98v��L�Ú�&h��B�Qo�SW�ɇ�K���y���ޯ�mE ��4��P�A��|�~T꣯��AXQ"�+�DWj����m4�4���?��U��@�t��t�.!�um���-���u�X�I�˺^=�E�zA�*����L�ݵ�Ot��%O�� ~�nzެs�>�c�V��F�x;^b��9���"I;�ڬgRv�&�m=��ۘNe-;��{ޯ��b�1�U|������<�g�%�%
Cq���C�(�&�]U��+��� �����l���z�7\��P�3�,�lLC�I^f-w8`�&��J
"!%&�n� �{�:��n�R\sw3Ug%
C�7ހ�M�*��{��VА$I`�N��Yv:v�m[{�O[s�
"�;g@��g ~���5`}������JJ�����I����s�g)�Jf�b{r�Eu$�u�cj�ᙆY��خ��f��x��i�>yl���R�Q�3Վx^9e%�R�����Ӝ0	�t��X�L���������PĪ[�-	�ՖـOt��g��!B����΁��g y�Ni�I6ąV]��+���_E�N��>��OI7@>����J�v�wM�\���΁��
!-ǽ\sw{���j�JT,�r�tT�Ws7b.�=E+ �n�Xֹ�����U���sp�qf�9���9��J��H�a��%�+�{fďs���u�+C����u���_}�p?�]�0��"v�*�6�-%kv^ŸS�e�ln��m3���������4���u6��C�i��i��0�D㍈�e����	��\�3�۟����]�v��\�I�=IF��.a�2�a��p��1T�[���q�9�ݏ�u��e-��`�e��z����t˅��	��yw2T�ҙ��p�s� ���z�,N��t�l-$��[�Ҷ� ���?~��"�$��=:eeW�7�Q�En�v��m�m�@�Ss���:~D(!%&k�.��w@����R��AN����X�L����+ ��7@����}�����L*ĭ�M��@�t��
���Ot��w���'��h�)j4~�n����#�+��]]�WQJ��l�i]���[���@t��o�I��۬wI�z�,y�1DDt�p�����U��V�ZߞUߺ�����Pq�0Qq���x�C�p:���+���|������;�� ��K)�n���Mݵ�OI��'���~�wI���X��`�컈�wn�$�a��_����t����Q�{�����t�
��i]� ��7@��� ���'��Z�？��Z�Ԯ$�9qA�k�Í<�!�<u�y��1:h�BbЪ�>_�k�e���6�ݷ���XN���TN�tHժ%�� ����=Ϝ��[8��@�V9�D��K(.�0��i�׋@�t��'�&鿿W�p ri��9{�����E�}�T�U)]$�iZ�u�Ot��w���'�ȴ
�U_N�X��6�hS5jeM�5}���< J">yM�@~���3��z{@"fe]u!���pb����[y�gY�]������ܓ��Cm��sиԄ�6�E�����7��=����3;��@�sp��1��Yd�v��|Iw�i��`����7@�wK�>�r-�K�����ww3Wk�{��zӘ뀢(>��w�i�/|����IU&R�%��,���1� ��=�����I)�$���ttj�Ej���64��Ӝ�@�
>̶p��ށ��:��d�;��n�/yx�g���ɬ��kq�q���W:�b�bPT�*�s00,�a�*Q�RM�8t�-�1�ށ��:ԡGd7^�N�٥��۲JD�u2U]�ͷ�ꄢT(Q'��� ��4�f[9��H?j7T͒Z��S*n���@����wI��;��zI7@>��T�&�&��J��~���!�{��zI7��L(�f�pٳ��*�n�L�]���������63ww��������@C@>6���Y1�<��њ�',�ڝ���F��C�[ps'S�_q��tk���r�o�Ҿ��xݭ�ճJs�/[�[���q�
*��W�#8�&㝚�3��<���mڧ;���RZ�;mȚ�Q҃�v��E�޼��n�=^�d�����6ܝgj�Z��:v^���%n���$�r{Q��+z˷R��=�hK�Pl�ۣk���գp�<�Jm��N��,��l��c'w�& ��k�##�W1�G,c���KBR]�p�l�i���j��L�
���-��&�aj�V�[�һf�w��/t��L����� �*.�*���ݍ����/?P�d4����t��F�T�V�*��ӷxt��s��$��oE��N�U�4�oxt�[8�o���u��J"" ���y�@�is2��EH�.�jj��nM�>^���2���t�QC���nмr�G/����:�w�ŷ]r��
���ۦ�bO�eKlu5F��K�Iv|�p��΁�e�aB�]�����ѳ�Fҹ����W3W\1�s��BQp)���Fg-��<}�O�� }�)ұ\M�$�I<�Z����t��S>�ݮ ����bn�*\��T�j�욫8�"'7w{�=9�\1�s�ؘ�|Ӏ6,ڝ
�sw(�������u�6I����c�8�o� ����b}��؎��C�tz��s�\ؙR���6�v�ď��eV{{��a;�ǳڴ;w�wG"�=�p�=$��|�%��tl:ae$�4��-���I&�/Ix�d4���B�U�WD�t�jj�����>�7\*!l
L�_���o/߷�}�����|��.拙��R���_z0��7k�n��N��e��6��@>����]�UU�M+w�I&C@��{�0	$��|���ԗ�����AF��JGk%���ǭ��^z᮸��	ãq�r�.aq�����뗇L�t�o0�=�p�$�n�����������Pr�UWWd�Y�m����	)=9�\ww�t{-�ؙ�4*��+S5wwwwށ����$�!���UA�s�$�tH�d�*�b�.˛��DB���΁�c��]�{�<����L�B@d����IOE�9�s��_~_{�Ѭ�6�ѭ���9yW�}�U�Cwwy������:�l�"�47�5���;{W��؎'��x<ۋ��!K�]��
�M	U�e]�t���X�M����ݷ)DB��>.�y���R����Қ��@>x��!���=��. �o�Ԣ&C�nĩ6nꪪ�QuW|wovz{$��o� �tx�r�wJ��ݻ���Šw��p�}���"!�nz�l����b�m�۬I&�ӣ�'{��<�߾��*��d��蘐�&(d�[-$�q���7���e:�1|Ϫ���
H�����=��3x3�07Ȉx�B]�"0��F���.�3��,��\&y���=(s "�Y�a��m�d3:͇�_�2� 9�|ͬB�}рs9$�Z�@A"�5���X8��X5��f��9{����!��֚��k.0Q0��$�g�R$�c�1�ʤ
"�2H�|��ᙃF�ŐB�M��L2��Ǿ�~�K)m�۲�ʰ����
��j��< h�.yR�8]�;�Xg��<qge!ή�*gn 뮲�;+ћml��'7 ttkq<���ͳ�u +�vU`���q.:���:	6�Z�h�$��5Ⱥv�^*�����5���)K�nm����L�sr�Ѫ��׭�rG��m��cM���Ye��[lrA]��b@9��X^NgOCL`��kIb�;s�nE��QmFx��v���:�#˲���y�����W"��k�d�7!�I�2�0(R�G.��{s��c���`�E�dzo9�Ƙ�����K��̭�m���v�ǹ�f7l��y,�l�g��Y�l�<n��N�<�]`�tkH;% e6�m�m]�d2�z6���C�m1�շ�Q=���iEuWa=I�tk2����1���f�b^;#����ٯ�F�\۬��:s�.+��ڵ��:3D�k݄s�-���6��a��Mf�n ����(��{o<vG��h]Abݶ�M�r$��}�GQt!fk4t;��3�u�dL��ln��I��&��u�D�\�\�c�nR
Ԣ��ʵ]:���67J�t�n��s�MیKWJ����9�1NCi��n�+��|���k���ӡ���C���������L�t8����������=N�׋�6p�ے�
N���t��ƈ��gdn6K,�qƞ�g�&Rp�K�㳷9�g.5�C��
�tRA�m��c�=�/��Mm�nMH��pd���g���kr�����"�9^��ºo]�%�հnCQ�s;q�WYyN3���a�4=��] N�W\�1�(&��n��xK;[=���[��@ax��O^wk��.B;5�y� 0J6�M��r[YҵJ��h��r�������6 ����V74��ir
�N*��Ur��(%��1fm����^�<i�����Sz����vt�K�"8�W�����:4Qf� >.���^���Ś�6��VՕ�Z������Ȍ������� u���U��x�����T~���@`�8a�0�i��+Z�I]r�8��ȳT�i��t8ѵ�[bLY�B���w@�l��n�vs\q΀�s�v-�N�ʗ/g�s��U��A�)���J���˱��ڕ�d��ck+q=��������C#���4-���-�nn�͘u%���u&��l�Ց��cs���yj*T���tk��rm�J0v�Hz<e��'!C�Y,%uK��-Ŋ�b��H�N�ə�����&)T��6���W[�[[��J�۶Mn��^��=5���������퍺I7m��hN� �[s�3���"#~J�wy���rQ;E\/ց�i��}#�h�XwI����j���n��Q�̑4���������wt��zG�}#�h�]$��2��;��]������ �tx�L���t��>�B%m�N��T�]���f;�����ox�f7ށ�/���P'bi�$�D�DnY*�K=�׎u\����)�=����-I�ظ�f��W5W\���>�|\3�QHz[��n΢�T�e��Mڙ��p�f[9�*�Q�I
l˶��{����$���Ʈ�]+M�Wl�;�M����>�2��x��]���i��{�wG�}:d4��0�I��,JSe+�t�o �t�h�p�;�&�ӣ�;�H��>d��ѱ��7n�ŶD�_7M'0<��{;k�ױ�#X�3�3;<����&�}� g���;��ހ|�ޥ��>i��L̦�YUu7*f�����>�a$��{^� ���=����s57r+�nں�v�� �tx��!���TQ���c1p�`So���{�ʽޓt��J���t��}��t�[8~�}�l���p�墩T�!�]��J�a�w�� ��M�>S���vC@��U*Ie��w��?[��z��w]�Fy����_'���n���18<���i��&�'l�>�۠|�%���!�{��}^�t����5An�+����럓'ُ�t�zp����<�abQ���7c�x�ݐ�=�p�����7@�zK�'�WQ���������9��p����}/p>�I*�)N�:4��a�s9�-�UI���ZhZKH0`��h*��1���kDe�?	�=x
��_�����_��$�T�6�i	ݶ`���t�}ݐ�;��}�Q)n���I�I-�w=y�m��9M��;Dm�\��v��ћ�[�gZv��J�1+M�j�M�;v���:^�ݐ�;��owM��%)�;�W*��w38��
$�{�ð�g����l���ٓ��CV���.��ht��7���_��S���vC@�n�R�s6�ue�U��lOُ~�:��~�q�(P�>.��e5*�]+�ujj��ϛ������>[�5%�����Jf<;�|~��U��%�]���&h#	��u�U�OW!=�z⊆�H#]�p���p�[���c���%&��n���^0K�̝\���9�t�
�%0']�\lus�Kt쐖n�����:ی��5�{rsf��E��י�lɛZ���A+�[R����T��hyr��=�t�x�������ۡi��������']k�%��[��Z��Y.AO��˳�v"R�����\@W��t��H��3қ��G��;�;lƬ��X�M�*�I�]�jK�����1�p��}؄DDG�l��pcvW��~�WI�op�'t��7�t� ~n�}��;�"!%0�"L�I�����i
�۬�I��=#��ߒ���`1�p��ʩEMMUT�s�(J����}�;�V�wM�	Q(�Q:N��MPշ�o��-�W���e`�t� ��<����]b-!��g'n�:��Fx��y�����i�#svgeu�uwcM�7���t��>�t� ��<�UT���@��]_蓫�m����r�����y��)���@t��=m� ��m�@���sa!%f��b�]ڙ]\��������[s�=�X�JQ(
:M$��w�����"�=�X�|�%������S�.�W{��{�V U~���4�H��9��Y���iݥ��mvSu熞��JK{4��v5��Խ��9�2�v$����ݴ��۬��M��G�oyȪ�@�t��=�J��t�v��.ɫ��@>�L�<�����p����Jb����Nͩ�Wv\��[�*�����<����/�}H��F�P⎓	�$]:-P�C�2�)�:0t#!��D(�.��=�@�o�7�IҷI۱�&���+���t��>��n�}��T�����n�IJV��H*�U�X��M�*���#�7�r-�镩.����(�vQ��BQ$�%J�u�.��K�M'�mˮl:��s+p��2�r�]�7n�[���/ ߹ȴ{�VUW�>��n�GM&�T;lm��s�z����}�c�@�|�r!(�f*��UJ�Zi^�-�镀}�t���/ ߹ȴ(�V]Kݴ����">����}>n�~�nzG!y!Ja�P$�H��!J�,RNiP1	�s���t��Vʶ��Э����^ DB��X�{���}�}��| ���=Z8��g���q�h�o9�hݭ�s�����o:+m�+����\\���3������{�V��_���H��:�]J�t&�v�o3��t��7��t�7|��n{��J���۩)N�ک$��m����t�H��9��t��>��wN�ۻV�@���������=����؄��S�~��(ڸ����]�uw|��nz�A	'�z��{ހ|�� �^"P�ؘG  ��F ��V��X���)���~�w�V
����Oc7:�Wi���=d;]��f�Ìnܛ8�Ly�gnɹ��ҍe-�M]h��nzۯ5;ZC��n۸�N�;/F皞v�i����q��&ܖ�Ӗ���<��ܚ�s����/ev����K�Z��4uݬ>o�7=�nš���/odyòl]y\�*��Wk�ۮ�g�A�r5�=.�ϴn��݂;x�'RM�슕R���0���������w:{ev���n �@�l��%n5�A�:6�hy�lZ����:����6�㪴�߳�=?����n��^W�g��@�E.˩c������u�w�ӽ�2zwv�ۗ�=3����T���v���$�g��@�镀w��t�K��S�˻n˫Wn��r-��V��M�?|����z��RlI�;V�<x��X{�7@�I/ ��"�'�E�Wwt�X��]-;�۷gY'�F���/=����0������eR����U��1]
�m�Wm���M�>RK�7��ZwL���:�SwMP]��/8�����ˈ�F�����G�舿U��}��U��{Õ}����
d�(�F��ՁD�]�w\�m��@���p!����}>n����.:k�V�%{��{�V�{��/7\����{=����U75W2M�U�ｏ�bDG�7k�}��=�|\R�i� *&�\T\�ER�u71I�˲��
��z5���
ҫ�Z\�!E[C+PO��V�Y*��7%U���=9�\�׎z���bd��z�^��5j�M]U*����Ϣ�;�2���7@�zK���R�):hmիO3��t��;�t�?���cF2FYHFf!Q1/�l*C7�����5��P��g�G�%58@D�I>	�0�����'�@�&��Q4E��ޤyF�?)�m0��|��K�����#O���Q�6P��f��1�kx`��1�/(bS�9`p���?"o���2��������JF�	I!
 V$8ɴe����0�E���hw!�b�`& �y�q�L�a�D�Uљ��I^!�p<g|��X5��<�3��&C��a�`nH���%L�ӏ�Ǟo���"�_u�ԙ�2fL>"ؗϻW��(}W �H�4���*����O���C�}����+��G�D"!%���k�{��bmL���DȪ�j���"_��z��� ��㞀{�<k�߮QV[mZ��ˤ�g�E�� ��t��K
`,�ɭ��Ou��=#v�ŋc��um�pC�{\��k�:���M�W�m�}�{�<��M��G�z�aq��S�c�w��{�<��H��������g�E�z�˲�X����Bn�x}|�K�6yȴ���}(�q�&�v$�v����^��w<����+�ާUS���J+}G�. ��~��|���a��v��Y�wui[�g��@=���M�>]?MIC;>?O�ʂ�D���H�,l9�{�ݝ��n5ɨ�v.��ok��T�~���������V�/�:O�{��ˤ�~�E�uH j�ZJ����+�|��>���ߝ�= �c�lBJd�\V���j���j��=;�\�;�hwG�{���ȩKt���%uvU�p5(���ݞ�6����}�jS�����j���dܢh�3]�'���{��ށ���w<�΀�	DZ�D	!x�C#�d!�����ۀf􋥔�C7�� X��ug�V�++�����Ubuk�Փ�/�Vi ��'u����+s��,�#/$a���EGg�'h���ۓ�f��m��y��|d3Yh�����z�\s؝�OUk�,I��c].;rf훗7�K�N'�].�N1{ut��W�,mPOn��,�h�r:]��ql���Ʋ�y�+�y�����4��� ��Z��8M��2�pV���̒e!#R`���ݪn8J�U&T�R����fM��c��9�M���\����uɺ�.G�at��m�߀߽�t��������oo�?j�EmҺ�j���U���$�d솀wtxw�n��zԻ�m�wV�V�����vC@;�>�D�x��ӻ���yHڵWrM��Z��a���|���l���=R����ZJ���ڻo ��M�>]%�'d4����r �W�Y�����iݗ��ϝ��t�s��9ֻU۷����hò������2���m�����<���f;ԡ%���z��I��.j�I��.��q��IC���`30�0,\,a1�k�(��>?_ �x��>�n���T�Ze�t�t�{��{�<��)y=��<�i�<¥�җaJf�����~(S�~���\�c�:��|�N]m�����ot�����C@;�<�{�����3��ҵ{
Og��lJ8���.�(8�kV�W��RYj�WGb����+$��Is�~�ˉwG�}�t���^ w��D��m
�bum^a�� ���ˤ�g�C@��uj+��um;o �{��U�=�u�b� ��Y�]��4����U���n���v���>�n�_��f;�j�J^cߺ���3Z�*�L�j���_��6Q/wo�<ǽ�6�<��TUՔ]]�� J`�v�/L�z�t����Ln ��]vv�.SAutSe'Cuj�Uuv4���G�{��$� ߤ�h�iEuq��v�I���=�t� �G�o�d4�����2Uh��jmL�j���������3��|��>�<Ss*���cnڤ�o ߤ�h�<�}��y_@��Jb�J�K�0�!&H��GtJ���|Qؤ};_}| �x$��j��j�˪��p�m� �ُ� �����5DBI?�/� lm�b���TJ��Ym�jsOp^��y����닸s"��py�^�����6ߟ���z����>3�۾�	�9�7C�i��ot�� ߽� �%���}�_�F�&uQ(ER���>�L�4�����ݺ��� ���R���&��ƕ��@:H���n�t���vC@�(��h�wlI���7���G�o�� �#�2�$�)�
w��ȯu���o{��-��m0�mã�9ӹ�sX|0�_3�4-���vq*������dK�g=���m��L�M��4��Q2�h㳹��/��^���5�I��
���W�	��^M��d��n�qh��	4����m�i�ZAs�<�'�Rj�6�����[t���pa�8�2Uj�ݔ��X�z��ݳ1*{%�{0M�a9]�V#���f�D�!�!S�����`V���YU��Γ�7ng������m�����[u���;-�Jղ�Һh�N�m�@'�x�ݐ��<}zu&�.�b�۶�
��7�솀t���t� ���bL�{GKf������k�: �v�}�}鰦G���>�>i���52J��Ssuw��
!%?{��������t��{�x�Ueթ�tս��<~�d4�� ߽ϽS�{7IR���T��BU�r�us��z^;���r�%kHt�/c�BYଅ�����t�tRM:Wm�zL�4I��M�	$x��"R��RN�]�+{��N��� }x/��y}��Uw�{�U���x�Eu�7v�������>����IL����@7wo�|��ҏ�hv t�ot�� ߻�ˤ��U/�}7@��&�.�[M�T�m��vC@�t��o��tޑ��٭R&`ҁMȪIUE�6��Q9󫃤���<���H/2��P^p�p�"?1�b.��>�^��M�zG�o�솁+�T�ˊ�v�$��7�t� ��x���h^��x�F*Ln��T�ҹ��@=��w�g��P�Z����(h��CA|P�p+b��x}'���Â�S�N�I�W7w��ID��}Ӡd��p��}����%}┢:�H�ut�V���^�{^��f��}��::�-D�м������GZ M۝h�n+m���gu��q'�e���j�Hn�$�Vۼ~�7@=�����^'�������%�ww}����a(�3���@�������uB���T�������Wur�����Ɓ��/ ߧM�zG����	]:Ct�؝����~�<����|�py��Bf���D3>�^�\Ix�G����j�F���t� ��x��d4/Ix������PŠ;n��pb���e���q��klM]���.u�cH���X�c�n�pE5otޑ��ݐ�<�%���/T�MM��I&�U]� �1�v~'7k�}��z�7|��-�JWT�*n�����7\�6��bd�ݾ����>�d�u-��I4U�� �����w�3�=�S����7�ɭ���WN�M��@=��s�h^�uʾ}�{�xw���@S�O���2U� ��-���I�2R�$$�	36�sBѤ�2N�,�2������((�!���y�ʹ'��M0�9d�b��i�����Q�g�>�)�]A`U�F	�$��L~:�5���&�6DZ� �X��R��	>i���4R�X"����hK�DeV���D�DEU��7T�g���~�}a����ݙad<qSs��C���0�<��ֵ(' �9sbU0��-�>A2�5͚�Nl�Y� �&)�u��뵡�4�
��} �F��������iV���"����� ��x�C0�[2|#���" ���G�7N�0W����Z��ie|��XK��L8k4@h$�4�H�w���<,1���98�F��>��<����f�~fh�4�U�z��8�&	�fe�(h�4�Z,-jm�e�&�����;���L��cFg0(}�;'m-��ڵ����ƚ�I�$�%�I2�]��ݬ���\�gb��;ϳ��嚣Ypv:t��6<�����B1ج�7.�0��$��������dͧqP��㷍k��6��G&�́qd4cV��Q�.�uh�:Zs��&�Ls-q���wkQv���u��wI�Ww�������DN&1%�n=��+5��<kq�wv�z7�<!��l�^5#�Q8�]Wc�z3��Ƣ�K��59=)]@{��l�xq�i�Z��v�m�e��ny�\�96Z���N�3 �/Oqǎ�oFv�6�[2s�S��v�6�n�D�|�0���M���ɡv{Zݯ@p��n[���&ͭ���"r�D�h'����"k��C�v{S����3����/(�l��9�)���ψ�s+�m����3vgU��W۵nˡ�5�-�f��9J���e�%�Ҧ,���y4���������u{ub�;g3�x�S�h���hr]�[�!�����Eʊ��.�묝�,.�{r�vɰ�Yy����U�ܧ&I��.�X��eY������n˂�N�7t�RT���\��d2�1�涓��6�v�*�)�}n�X��v�`Wk�Q��⫷gb�ʴ�/
ض�8�̭�Քۃ;3�R�uҹ�M/[v��'=��5:a!�`�.��c�r��[��$v�m-�$�e�������A{��혶&5�4��<vNz��Ͳ���V:��'KͺMZ :���u��P�g�z	�Q����j=/=c�Z��lW�]r�nt�k�<�"��n2�A�v��q��:n�=ڬ��pT*�97�[P�즘;�nù�����+'�;Z{C �m��׫r
u �p�u��.�YNѰ3�1Sm��-ɑ j3���j8��W����)�A��x�󭉰v��T^����l+]��`��;��9��U�l)���.Sl�Krz�
��m���:�힉B���7g^������H6���ƍ���V��JD��a��s�0�ø��S����pQ��� mVP�Y�e1FWbO��U�� ⡿��s+<��"�^'GQ�%��R�YJ�Nň�;<U�Fy�v�^3]�9F�RN�Ա�M�v��FmAv�&0r�Z�#�ȏ)��ƹS�K�Y1�&�su���U%<��=�Fψ���$;csA`�۬���A�g����=�D���mdwhx��{n0�D��tcF;d�͎�Ok=	j����`���MF�Y����8��{<�X�Ԙ5V��L��{��{ǹ[����v��*���2A���6�����ݫ�r������V�Cvܹzx@�+rԜ�m�;��-��^����� ==��7Iݍfb�<�%�zI��H�{��@��;�R�]�IۺI�w�}�&��#�=��Z���C�F*T��:.��V�@=���"�<�%�t�t�Z:�ڻ�RI3v���{2۞��
2��t=��@>�w�5Fc6f��L�E�	���˜�7=�gu�CN�g��u�طg�'b�L�9ۭw��+������i���r��x�$ހ}��Wd1�ݞ��;SKjԗuD��޷�U����y�$D�TSz�t���9��@O����ZM��@>� ��ȴ/t��I7@�JM%۷t�j��x��E�y{��zI���x���'V��UuE�9���c��
=��������[s�=��*��J�nPR��N;n�gNL������v�q�<ѼK��n�TJן����-e��)*n�M[��I7@>� ��񚾐�ǵ�5�:�2j�n�U�j��ޑ����X�$�?��GTM��&�n���wL���M�K~K�T%
ӵ﷽ �� ~�KE'BW4T��w�CRIO��� ����=������'�]M:�%�X���Xޒn�w�<��"�>��x[*���╓SJ��VP�t����A#��[��n�%"�&:*�ej	�0�5=v�n���hm�����{��@�_E�}�&����Q�v�[m�HV��e�=�
!L��{<ٻ��{�@���45i�۫nƳ1hK����M������n�g�8�����6�V�X�$� �tx��CCꏮ'��ߠ���Ͽs�w���t�4:���;���w�<��!�}/��>�&��!*�*�Iݖ�wB�E�/7�l*�ݒ-��n^��7a�n��J�n;y��ۢ���!�}/��>�&�� �tx���ԫJ��6�p�>��`t�t���w9�URS �gjjv�EuTT���\�7�ހw�<��"�>�p�'�\���i�����ot���{��@����{�w��TܒV��Z����35w�=��}�p���@>�;�	\!Dx�;��n���g����m�w��q��i͵�S��e�w9���
 <�(<�ա�s��ӹ���P��"�]��N�nW�s�p�&yc�wh�⢧�`*m��MC���Ѭ�(�ۃ�l\:���ǫ�wۀ��9�)���u���v8 8������q�]��nj�(r]�³�c����ތ��e���2E7���D�u9"��șm��t�|�9ʂ�L=����vٺ��n��g��\�ƉC�k���y�w7Mɫ���[�[��k�4����n�}� �s�h�Чd�V��-[f�I7@�{����΁�����2=:�����eڥot.�׀w�d4��Ӥ���\�m��4�;h�w�w�ȴ��Ӥ��Oz�)]Jc�Ʈ޼Z����n���K�;�Ⱥ��"'[Ҕ����&�3a1tLՖ�m5�>�bɣ;�wC���إ�u�t��	nEuTT��5g@���z��u�3�m��!짳�30�ڻ������任�������(F�V�O@G��K��Ym�@̬s�>x�zy���]ڔ�۴�J���r-�_E��Dϵ���zq�p��M�]\�ܗWv5��@���`zI���/ ��"�:�D�(��
��m��I���/ ��"�>�8`wDQU�(Nհ��
˭�q�)�m�v)9�v�P�vS5�]�q�	ȉU�*�T��Iyė_��5#���@���}'M�>�ˮ;m��I[�����"�>�8`I&���`����XҫMSV޼Z���*����yxz*��� � ���BIz$���]^� ����@1̺�R�)��b�����t�%��2����R��v�V�m��^��
���'_E�}'M�9Px��R�U�G1�$��l�(�E��m�:B��6�
\�n�%�պni+T�Kn���C@�}�E�/ 'ޢ�6��ݺ���4�u�Y�$N�^������;�_Z��t�Э��	;��zK�;�r-u�X��
��]�w6�����S����;ݞ�����	CP�^S�w�}'���t��-�m�xw9�:�,����9�u�1��TQT���\�X6���v�R��[�<�Þ<�FNf7Nܝ7��H�v震J���X��V޼Z�����7[�o/vz �gjjv�K*��K�]��}'M�"���wzd4	��`�R��4�I!���/IxwL��:�,�$�ޔ�V�M��L�����/�N���� ��}�}%��������ڶ��W�h����7ހ�M� �c�:Q�	s+������n�v���M5���6te��aF�i��wM@�a|����"�R��=g�u�v���hv��U6�c˱È�󒐺��Moop�	��CZ��ܽn:��z�ӣ��]a饭�etj{�+����*ڀ)p�L���Vt��C�T�Z��s�9WN�8���n��졞ϠA�0���B7Kmv�h����mcd�g�0��!!��|��n�w������mp7�]w����ZH9�,�Ӊ��9{$s�֣G��;��ހ��� �e�?��}!��� ����-�n�ݺ�ot	�`�9��� ��>�aDD��0u5�t�R����x���+��IL�[���ݞ �򑩤Ֆ�&�\��o��WE�}�&��"�=�r- 蒊�X���Z��m`zI��Ȱ{��@�}�yD�����v]]Г���3�R���w=�-֫�9��40��7Y��/U����殛� m6�@���s�h���>��tzRhQYn��mڧwn�}�{�p��
�0�U$A�`�P��D�.��{�=�}�|�sRP�Cw���7j�m:k-�\�X�$�z�X��s�<�˥C�B˹&��x�^n��r�g�y�=�c��,)7e[�N�;{�O\� ��"�'_E�w���w�D���lv�B)R�.9)�ݞ�a��t�4���1]��s�i�2�V�q���m��U�n�k ��"�'_E�w���O\� ��
�S't��׋@�}�I7@���s�hD�Wr�N���'��k ��M�"������ ���sX�� �!�bC$)A3AR�	���PT��ӣ-	�F1�Q_>ܮHDD�d$�JA-2�r+��I-�Q<��v�#���%�AB��`h�U�
�f�6I�G۞nL<ІIA40���Da�������� ��"�-ٴV�p$K�,b�=�Ş�0�L"�8cV����.��i'�#�Y�d	JDR��0C
4�Q��DI��3*(+,Í�·�dṦћw�K0�Dpq�#**�H
���Ȋ.O#TF��,���()!�!`,ZV��<Nb1�ٛ�f�4RD�-C$E7.%��:�3��Z$dBF&5�;p��gxZ5�h�I����
z*�P��>�:UؿA~
�.�O�� §�Ȟ�DO�}	UI,�؅1ԡ'3���=�M� ϼj����v$��ot�%��9�:�,�I7@��;ID�n��wv� ��ȴ	��`zI�^��zt+v�mc�1�1�]j
�T�N�������e�A��\oLN�F:��|}��� �Xi�}}5���x��ހ����.�6�vz-�2l�	.䚻��6�{�B�6sv�7{��V9�b�v�������zK�=��Z���I����J�*v*��M���_�s{�:�{<�m���P��A��04�@H0�����?o_�g*߽�4�YhU7*��:��<�rn�=r,��!�}���괝*K�ӻ"��mv�{<s���S���NN5nn��uX{��uUІ�j텺wwWt�m`t�t	�`�u�X���7���-w7wހ�M�5BS&7�Ӡk���>��{�$�L����gff��M�\�������t��xj��)�f���nV��	=GۻM�+n��u�Xޒn������=PR���4�������E�/ ��d4	��r��H`�K��0�D�w��߭v�&�yc`[������x.���&z�a ��1�����L�ڹpy��H�i�h�Ӭv�:;�!�M�[pfi�%j�u��][Z����b��gF.6�G���i��d\S��V�s��v/�3y����m<���Y4�/�4�J��Z�p�i�H��.y��g�݇XU^�U�r'pF��Ԇ�[]�h:غ;d{��kq�]E�o;����f���"TM�cB��UZB�͞��8��y���;3�ܼ-�(���[��y#�gT���n���f>3�<�s�>��z���I\(b�Ui��k �t�h���>�&��"�$�KIGCi�j���N�� ����O\� �t�: ܒ�i�v]U)��SUs��J"'�w~���<ُ��+���i�(���i���Ȱ�u�X�I�C�~Eݖ5L_�]��vr��잹4�c�֎�`�ݢ�n���u���d�6�nګWm`�2���o��!}!�[���Cْ�]���귻5�^U�u�s�����:�r�&�wK�;�d4T;PWJ�7J��X�t�%��d4	��x��\�W�諙���CT(Q����77y�@yX�<���>��R��P�EՍ��X��u�X�t	�`S���V#��t��l��9���)s�l؍�A�⣐N�8���XΣz��I�j�E�SJ����	�&�zK�'��h)�V���X�:&�x�o�ԒP�M�ݞ����c�jJ!L��5S[Qq2U�M���nV���|gMp�C�@P'	
$�8�Sݪ���7w7��j�Ih���UW7*��灩O�w�tݽ8wI��"�}PJ�[n��H�{�M�$��I��?�n-��USD�D����*�R����rn5�sշ ��Х�i�9T���m�;O8ً�V٠t��۠E$��!�I0g�j�
�-Z������@rۮj�
����tݽ8ٍ���"dr`�Lֈ�EJʻ.���i�v��t��E$��ߗQ5L�Ʃ�i�Q��Ӏy���-��}��1�`��'h�#��w�M�D(��6;V+N��`wI�RK�:G�hG��PUݖ��T�D�)2�֪h��� 
^8���Z6�nֻqv�*t���ˢ�_�X��ot���t���$�I�t�S�KcUv�wWwn���Z�� �:n����@�[��lw��@��87��6"IL�����og�z�F��[�Ym�*ն`'M�$�'�cw�z
��4��֪��V���fj����lBOw�g�7v���>��!(Jd9�M�Q(Sw3w9N��ڌtiR<vݜq���v����c���.c�i�KnݎɰnFIG�䵉7[��v�ޖ����q�(����<�j�'ZӶ���%ۋX��Y��{lFB�-���J�i�%TE�lh�vRJ)p��b��ϱ��h��}�pO8s���g��$�];�up<l�FSjxո�+���u�7��݅�m��zd�Ѷ�2Wm���R���{���n셑1���u�nM�ca�� ��`e��	ة��XsԖ�i*V$�ራ�[m6�O���۶p7������ݞ��-j�+T\��+����g6&L�{ށ��� ڠ>RRRՎ��Ҵ�f'��K�`s�	#��BQq�άJ؁&��K�`s�	#�'���˩aI��MU���	��-H�N���Ir,�����V�S�^V5�jWt㷗v�c�K�qD!h ���Ӯtj�?/}�����f���1hGw��)%���Z�j��]�ۢ�[f;�n�j\Q�\��� ~�nzn�ͅ
!L����%U��T�]U��l��p��-H�N���r��J6RB�C����=E�I0	ޓt?�W�[[�\�D�m���T�첻|��۶p��z��p���@��)y�<n�K�9wF�F�y���n֧����zV��D�n��x$uա{%����n��7M� o/��A�e�ߛ������l@�m�˹0;���@�0	=&�t�\.�ۤ�����\���~�<����r�(`(��A�bT	h�I�
	AH�
�	R`��AG��۝�t	/����]:N�ۺm؞f-H�I�7@��/TB���u����m�MV�I%]�M]��7ށ�������@��g ϛ&�5�������UM܊B��p�{FM��\b6�u�X]N�/m��lOa���U�[��ot]��z>�@�G�t��r�jĮ�'iح������p}���d�:�&���m���T�캞�'�{v��Ǐ�'1� �y�Z��%-X����I�V�q��@��u�=��s�؄�P
"�Ҫ`qS��{�\��?���F�� V�������>�@�Gd��uEL���wE&���]��ڻ:��n�E5>{g�q���a�n���۱V&ƨI��;��-�0���UUW�"�����'�n��j����3����n�˺^�G�h�-Ej�hE��Vـ{�&�����}����⮥Zv��SwJ��˺^����p�=�I�/*��v�Z��v+w�}��-�8����2sp�l>�s�;"fH�2�a�3�F,�����>��t����:��A�Z�(�D�3Hf4�ܜ
9+�RD�D<3W��������I�<s����LD2��TU��77��W��;07���*ۭa��"�E��`���)����ך����h�j����0�J0�&�rbF`�Q(�cKD�
�b�4L�ٖ�-�ӃȈlL2й�,DEC��V��C�!�6ț-k��;���>�٫,]'J_eHѲr�ȣ /p5$l�����.�%�`�HwP��&��',i�H�'27�͆Va�DS��z����&MCe��u P�0��9+��T���>u/��a2��Jr*�33��K�q���L3"�N6�����T�w���!����-�����A�`՝/��E�������X�������bȝ���Z��*�t���ӹ�k�e���Փ,HѮ9�{g��%d;V��]N%�t[��ج�����'�۱6˻d�֝�QĀ�]
��ug��gj4��n���nA�k� =�]��<m�݊�!{��q�\$��c<�׳[���t���lVS.�ȯ�y6�rv8��V#�\��:���vK��v�U�X:j�d]�����<�������ƴ����Qq�[hqM�F��#4
̩ͧ�u����W��l{n3˓���m�nǎ+�78��Z3��}<lO�U����9FWp�y��y�\Y9����nw��dּ̖Fv�SB��iѮn0��lp��,e@X��bu���2[�D{��3�����6���fG�;=�/Ff����ӏU���`�%�㋴�>��&[�^�F�u����QObw ]���ru.�F���s7�����Ժ4�^9M�\v�Ǳ�0Ӷ9j��\�a��NAԫA�ۭ�&n�&8�m���f�0�-r��3�u����c�XӜQ�;�v/&%x-�����f�9Zg2�&kS�&����T�W���m�ɋ����l��i9Lu���k��*�T�^�0v�'�)}m���ke�QGtv�4ʺє��Z��!;�ŵ[p6�Q�ݮKa4���C�ZXYv��Ʊ��;3���q=4���o�����9_�8�1����p�2HS�!��;n]s>�؍��H�K6�1B3�kM��gd�֗6ɰ�:AɷX��;slohi�G'�W��<̕�����ĸv���z�O�������f��^ח��	 �裊^u�7n��u�4����t�<�����W���;@\�ݞ8�\����,��ݞmL�<,"c��O�r��\55\��0ZWh�뛇�llZ������Υ�i���m����KdH�:�;s��������h9]ۣ)�#;d�μپ��>3���6�ޘ�<H�e�͙ٗ.H햶�;������������~�#
�(�C����*���'�1@�+>�Qf_s���'lJ�얥Rn�b���#�n	"h��%�U]����*��L�\��v3���z�6�bo&՜n�6c� �6��̽��[�gx����ķ�j'q\v�k&�]�|��N���\/��q��V-ob�ݭ���Ý�Ȅ.�ȝ�a�׌l�W�6�iΞ8�����<��/�,�$����!��vu�J��)F��rCں%����g���{n����*
�2��	R�����T�g�mu��q��3�f�v��mɺ���_�zp}���d�:�y�9��4��cc@���f�M�9wK�>�s�>n���2}���ۨ6Z[��@�O��>�}����7@��2�[(m�m��I��>�}����n�˺^ OW��n�n��;��b�>�� ��&����z>�@�а�B]���;�UVQbzt:���gl%�������J�8���b7&��I[f�ޟ�۠r}��-�0	_�]J�Ռ7t��������@�&�sRB�4�	Q������@{��ﱾ�aDL�LN��T�S*n�蚺�ͷ��>n��=�I�.�x�R%(�V�%M����l(�n�N�{��9���IO�x�zNj�ڪWe�&虵svp}�n�˺^����p�;��%4�r��.t�Q�;��X�,�3:켷V�[��V��	x��Q�Z}e�v�J�~6ߙ�u�;�x�|ݳT$�!�o{�=��R�QweU�JQ3w\�w�{�
Q2{v�����'1�5D�kMj�n�Lͫ�����nޜ�c}�	$��� �H����g{�\��޹��*\�S.E5wHU5vp}�n�˺^����p�%|wT�R�d��5Wށ���l$�(ǽ�O�{v���1��z|KJ�.��uq2���g�㣎�\�f�nL��.����<�5V�����6ӫV�۱[�}E�}#�ﻦ�wG�N�T�p�;�֩��׋@�G�t�������IK��cT$�'M6`��� ����E�}#��ԹZ����fd�����CR����� �m����wە��`�8%"r�Q��Dd!��O:5DɎ�weU�T�$��>�}����t��ԗ���!,mV8�(�m�[��B+�j�<�ۢ�m�Z���+#-��8Z�H��R[��J��i];�Š}#��$� ���w>�@�t��t�%nm���w�""Jd{|���>n���� ��;��ڵot���>�}��
"g۷� ����b���wstLԅ�eݷ�os��p�7���wG�{�)\b����k^-�0�o� ��|����"����~@ݷ�q-]]T#En��S�hӷ�8�ʝ!�$R[�s\�/�ct�ݷ9u�>:��;7��z��V�u�h\�;A�7=��Sm��I�μ���6�l�q����f�v��۔t;	ۮ�Ĩjtܫ�˴r��-ƕ9x�+h�nx=�K�c���A��h��:�s�9�'/������O׳v��a�7U�==��o;� ؞�]h�{����<�e�MmK�Lr� �pv���p �J�����r]=p�\�]��c@�q\!$�'M6x	��n�wtx�9��ފ�+W1[I"�[ot���%2{v�g�{v����{��L��(7fj����T��� ����@�����n�wtx�Ht�wt�Һ�9=��3�@31�aB��n�vz���ڭ�q3WT�SWg ��7@;�<��@�G}ĕWE$�ۮj��O퍌�qݵ�&����ѣA���Å�|��)c�2�����G�zG�hH�t���}�Z9�jh���ɪ�����r""�(S���0��t���>�Eu+�n��*캞�'�|ݳ�c�}�BS#oo ����EC�V�V�����n�wtxO9����W*�r���fʪ��3�{�Ӡ}#�����t�H���MC�2�u�m�9��}jk��]���v�z-�l��l���hmv�m�J�M���0�|`�c�@31�6�n�Jں���s4��g@����=��ހfc��-�����p�%nm���n�w��|�;.�\7�8�NS�H�J.!GN������1|zY2仺i��+{���8`����]�}�zQh���+N�.��8`���=�I����S���U0�ë�aW6�����6��z�)���8����,�E?�H��l.��]����}#�ޝ7@;�<}�u�v�N�!�;l�;Ӧ�wG�O�� ����J8Wuq;V�cV�@;�<}�>0��҂�D�ګ�T���TDD)�o�>n�ʽ�����|�e�d��!��$$��iD|�Dvo���z�`�Z��Wdӵ���
G�t� ���	<��\���BG�1�#���K"j6����Nw^:�ɚq����z����J��l���0��VـwN���'��>0	���j$��b�[V6�@;�<O<8s/����DL�h��дYI�+���0�|`�$� ���H��W���C�4�p�3}�f;�lDB��|g >2[��ժ�.�f�vp�o�g5���l��/�<�!(x�L�
�e�Iv]��,M�d�^+#mH�n2 ���\s]u�nѥm�`�3�u��v�(e�[C�ʷ��cA`fՒ�la_K�6��w	�gOfch�*ʹ�tA�H��ux�Ӏ�\�n8e�wcj�	��y��=�b����~��Cv-G!�A{N�4��/
�:c�.NCY�k��c��)��x[a-n]�Zx�.�ִ��.{��b�O�`3��[�	)�,ky�=n��'�����7&��\[ry�]�Ŵҙ�Qd�*��*�&l.�:�������=�>0��t��]w�i6�T���	�|`��OI����H;ґ�\+ح���;�� ��7@=:<{ό��wi.����Wm�I�tӣ�'����;��L���K�m����T��n�� ���	�>0}ό�:n���"IV��M=�]���Bq��=r�*[Ӳ��j�6�s���'��R���<WF�B���������?�v`�����]J뮌޵��̷�/*���:���t��"	X���������Q!��Ԗ��E����7g ow{�=-��:s� �s� �@�+.;��P�.���2[u�1�À{2��j�{����A�ɥm�M�;�w�t���c|g@ǻ��-���d�j-L�� �t�Lz��pnF1�;]�ۆ�uf��x᭎t4Ҭ"��:V�6+��H�}��zKn�;!����*]�����m���&��� �s� ���I�F�V��T��c���#�_;��r�}�%Rh��7�٧R��j�3[�u1��c��yP�aʔ��	�l�9���A�C�q��4&͎��#����]�PO[��K��cI��tC[�� �/ 1����fFkck�`aԺ<xmNEG��E�g��*m�1Q��Đf\dM�	
D�j����o���4�W�Ù���c�ā��1��h(>y�1~T�*�1���ou�˛��x�mb_}]{Ϛt�EE[��>�xSA��~2p~�4$�\�����7�����߾�aoE�R3���y�aw��U|�>�6IAY�E[9p�@�x'�	�M56�&� �'�����4W�va�Bt`��*��F��h�������Y~γ��ǘe�ˍ� �m�>:b�j9�AQ1��Hz}��8���0^��E��6�D�_������C�'��>+衳���g�(�CB"���R$JAЁ舁�|A� A�#���7@��&�����t�n����/�e��=���?!B������=�)���YI;VƝ��@��I��#�:s� <}�:��������>v�똞u�T+Y��;��m���V����;[�մ����e�m&��I����<�6�c�p�2f���Z��ot�G�zs� ���y��݄�Ob
ݺT]ܓv��������À{}�� �n��r,�n�,m4���4�� �ޓt����XBZ�~3Q�����ѣ��03�82�7'�Ht�%�๮"�?
�^y��\��TN��Q�I�tQvـ{����$x[�pf^a(��&��Mܹs¯N��w �R��c=��
�rӶ<:�b;+�H�[X(A���m�_����c�����RIvC=�{�=�����q4�������-���)��p�۠$x}JWR����cN��t��$x�8`�2�l-\����ɻ8�(����=ݾ��ٗ� ��a3E2�PZcm�t���� �s� ����
��
"�۩�j)U]\�]���n�EZ��XȜ�.`����]�r����m�ݗ�f��k9ì�:�5�9Ӵ=�]n��gn��^d��ܻh�L�ٓe.���:ܖ'���yz���m�E���/)������|�'>:�Goi[e½��H[q��K�v"��X{[���ܻ��W>a�g`�H7�鍸yu�n�k�q�x�d�t�N^�d�;��d�^i���lvF��?�w0�2�N>+P%*QN���k�؇[m��A��H{�/I%�X�8)���2��V�t��|�?�όݗ� �3��������d[֓*��i'��t���� �#�;�\�
d�i�j�;�����8�7{��<�镀{���'t�J�JaM��-��I�t��=�|`ޓt�Xtm;���v��;�X�ό{�n�zH��B���[�G\v�kj���1�@��ţ�3�jY�x3ێ�)(�AX���"�F�+%�8�����ozM���t������k5���7��y����6�X��� .���՝�wʼ��xr����nU�IPJ㶅`�E��� ���L��s� ߻��prw��*�m��L��s� ߻���G��WM������V�ގ����<w�=�|\b""��@'��ZWyy���,�:�U�w�۱�����x��泚Nn��"&j�.ݖ���?����ӣ�=�X�όwJ#h�aN��Wv�@:tx�镀{���7���~��,�]�v;���LN���{Õ}����$~0���(N��^�'���y�W~��Wϝ�:�ԫj��ok@���:n�t����V w/]��cC��bvp���@Ԣ^����=���^�����?WI�Dd@՞�(cv+=��n[h۰��.-����\�e����y����vE��� ���}�+ �y�oޓt�w�t;i�]���L�����zM�� }<�v�I۵i'��t�~�M����e`]\��W�Гv�� ߽�t+����}�V �	T�(D��H̍UD����*����~oەw�$��$��+UWSUWހc�|a{�tyl��ٽ�+	iV�ܫ���8���̚��6v(�����p��gx8�&Y�V	2��V���cL��ށ��X����;�f�b#�Kݮ�ٔ���W4X;b�w��{�� ߻��N� ���sT%�A���w3e�d�S7dݜ�=��;�
g<���c�g �kL��usTj��������׷�3��+ �y�o��7@���膛b���U�o ��2�w���n�t��%��,c�?X�?��),�Ԯ!�R2�&ӤZU��l �ԗm�^�M�p�ͭ�v��<xK(6ć	Li��`�t��ɇ�A����v-Ir#�R�]��˶�ݵSؕ�o`�&�fÁ�t.N�w
l��(���Pp�7g�����Q)���l��r� @ض��I7
RY�h�Ɉ��ۊ�cf9�Nۀ�I-��=lЍ2��j%�*ݞS5��W� 0M ����|���xc�&���l-�Z�,e3��v=r��*\����c�ȁ}ߍ�����{���ӣ�7�X�W&�|4Sv�� ߧM���t��=�|`�U�.�$�um�m����t��=�|`����]��_�4����7�X�ό~�7@:tx�%]J�~�]�v�V�k@���<}�<w�;�>.���8�Y�έ��m{d�ڡ0�"�y��7C���b\�}p�]��chB���:�������t�G�o�2�w��%A]�����*�*j��x�Q0�
!U~!���LCPI��!�1 !N���w_>p�]��0��M�:��[�l�n��U�o ��X�ό~�7@;�x�-RPjГNդ�V��0�t� ���L���ɫB�C�j�[l�7��t�G�o�2����������Tl�X�$ӥyqJ��0]�۱�V2�@Ruq�ê5�qy�\�8'msNi�wH���V�s� ߧM�>�ꉡ�c@ݦ�x��+ ���o�M����WR�c���^���_{���^|�{�G��)��#�}��U���W߾��*��乤ƇjժlV�~�n�wH��镀}���>��Wwj�i���M�wH��镀}���7�&�/�a�����i�E,HEn�8�
������:7[���qq���Ŵy��ݺq۶�:����Z��ze`w>0��M�� ztV��FI��I<��8`��t�G�}�L�(=]\�b�v����B��~�n�wH��镅�όwB�1]�t:m؝�����2����	~uT�X��P:u�04ՃZ��e�b�%qQ
!
}����y��7u"��-�m��{�X�ό~�7@;���~�]������n�*�pG.H��ֻ��؃�����:5�.2�i�n[�l���۝Sud���|nޜ�c}�cw�;�2��q|�cBj��6+f�����<{�V�s� ��Q]����i���m�wH���V�s� �zM�>�9e�Jݶ�J�[x���.����=#��I��#�N��&]��(�����.����D/����W~���Ͼ��Z�W���ֈ"������������T�W|�EG��A�PT�������jR�G?�kO��܈"�����_�\�����������������~���{��������������g�R��DDD~������EU���"�����C�������_��iBP�""?��߯�ߧ�?���W�du~���5��ũ}Ji��w���9�T�!Q%HQ%FTIBI`�THaD�`�Q%H!D�P���D�Q$�RYQ!	Q eD��BE�&I!D�Q$�R�TIaD�HVTHQ�TI�Q�AaD�eD�IVIA�Q�T%D��T�I%�R	Q"TI%D�I	!D�Q&TH�Q&@ !D�IYQ%IFTIFHHBTIVTIFTIDI�RPeD� %D��PI !D�	Q!	Q% �!D�TJH�%D�JfB`"B	 !  $$		P��PH	QBBBBQ		U�$!Y	BD��`!! ��D������B 		����`%d$	 $������BF��d @�HHU��BQBQV��$ Aa`$@��	@��H�$B$%	BU���%IY	BA�!	���$�� ��@$%AU��Ud d%U 	E$ @��@`%VBU	@��$!QBQ� ` D$$@�!BXP����� BB!	��D�����&BdY	B@��%���$Dd!ae!	d!F@���� � ��	 %�)��"�	dBX	IB@!@ !Q�$A�%��YU�!IBd�)P$$	HBA�$@�d$W��@�V@�B$ � � a	`IBD�%d	R@�B 	R�!	� 	BI%dd!dR�PX%�I�bQ%!%�`���R %D�%D�TL��5���������}�������������������{��_���"<����o�?�EU��=���/�}��U�EU������ ����G��3338G?��A�F���O���
\0Uo����?����DU����_�����}7��*����*����l����������_�Ϧ�~�>�."����A�}ߞ����AW�?�o�����AW/�����������_��PVI��Sg��|��` �����aw�@��� =:��*�A� g���m����8N�݀+�F�XLAZ݇��<�{]�dd �Ϩ � (EH)��%)��;c�J�t�Z R�N��:�;�   V�B�
m�Ԁ֍Cl�ho    ꢉv�;��A���o6 �o�}���>GsA� �l�pg��=;��9�Wڷ�o�꯽�W����6�rs�T��P�}�R��}�Uͪ�.n�t����aJ\:9��`y��`w��}�� �m�6�v 9*"[�G��+U���^���J_;� Rl(�ݹJP>�{(������J<��
R�)��7w)J9�a��w:R�=� �
[۔���JMf�� t�����t�=���:P)tΚQNvJP���s�
{��=�p=
Q۹� 3e� ��E��k�
*�i��n�F+�N����/��C݁������ϟC|�=�O^��������E>�}��>��Z�  ���m�>(�-�>����N�C�`�q�>��]�;���C݁�}���  �m�lP �} ���[g|�n��|��{�j
;�f���G�`l����9��|À ��s�̀�:��mx���9w�O'�:�}�՚Ozw ͏���2�  �;`(��� �P���_ ��������{{o�����1!ϰw۾��{�ҍ.�� �{�  >������t�[Z�1o�}�71�0q{������7�g��;�:>��o>�x      ���6�)P  "{J������h i�R�=6�P  ���U�E  ���U$�R�i�42DHCR������=�������������ԟ}�|?g���@
���w� �*�O� U���� EX��
���>dI�t?���fof�SDkt��{U�C�K�W;\��؞|]��B��+w�R�q�s�D�/�)�m��7��R��f�Sw�e�I��c9�L�S�[�)ͤ��fd��5��s%�X]�s4�h٣��tj�Cg��{S��a*N$	,H�F�2뛹��g��{O3\�}�n$�3�]M$x�<q,Y�,7����>�ӻ�e�]���[]���s��!	�8ˇ�Ip߻�Jc=׆��B��)n�$%(z���ѧ�a����� ��j7̄%+��X\5_՛�U����[�=��=�j�ޝ�1}l�o�vs��3�y�u�!<�Ew��xϕ����k;Y{{�|ZcyA��8{��5�1#s7�����o��潆��y��{O�J�<�R|�)%��3$��֘R0�Ɔ5��)�P�$l��0�
�#P���-tVm�B���	��!�B`a� X%(&;aq�1�IH5�`V��o���!��
BC�a��Ґ�a�D� �"�Cc��F)��Y�8�m��@�����$I�b\&���7ᰱ��@l�revAb$��0����p�����K��4xЏ�A
c����1߱+���$�ߚ��.Zj%���Gz�Fi|=w������1���z[n�}8��[y�]s��GsM�g��Ѹ�^l��=e2���I�\����⨥��f��E<��f�pO;�}k�fl��f��8aL��o=�,�9�9S�T+�VU�Zj�_,���[Y|�9=�ϝ,�Y��J3�	.��&��/P��>���ݫ�,1����|�_�*c.R�Jd)�)�
"B��[�1�;���*������>V�By�<y��s^C@�|&���P�~���<9琥&<��->��笡3����'�����IL�)�.0�+
˽V9}'�7�Hf�\u3d3Z	LȎ�c<Yo��-_����>������֔����nr�[~s�K������^�3?<�sV�}�z�v*�k�S�Tkq��V�t��q�K%��T����<����sz�|�Ѽ�5Nv�[� R�]�EY��TU��y�`��!R�� 2$bF���S�(d@�xD����W	F�0�߼=�L�L0�N�^>|O�6�OO��\޹O=��=ֱ)J�YT*������]�>�E[�|�¯{\ߵ��n��ܧ�Wi�%j�:w7��+�]c�9ھ��x닽6w�����mT:���hSs�Z���5t��||P�d��&�Y�gץ�N�)]���Tͤ.9�}4j�R���Z�at9�ѹ��7�<��^l#HW� K����5Öp۳wȐ�N3�5�.q42,��\e0�I�%3Ё4d᠏���]S^jy�{����]�j���#31��V����)v���h��B�����dK�8�ͻ�RK�2X繗�Nz�1��!�}s�{��"��s3Æf1޽���m��o���^w���/9k:���m�r�s9T+}��ͽ[f�[�����_u��v���(N����¿��e.v���\okn�A�����y���w�j�W�Τ=C߷�n�;&�����On|��[��~��/p���kRZ{).�o/��K�-��cD��kS���M��y ��UcZ�_s�y�f{�����F޳�i��=tl�X���u��y�7��CЅ&��Nx4��ޒY��]�S�P��D�jӁs2�{��y�5(M�� �¤h`he�������Aƒ�(a��21�P$�`�#2%�v{��y��p���3�>��Нv�����0��h�r������W����]������x�@�qrt���
�����k�3$����ڪ��،k���f]'�֫������OrV����,_|��F��R�K7�s�$�K�.$!�%��6�C˪���W~��R���\�R���/�����ݜ>+~��]�G(�eu���]r�|#�Iּa�	���Y���z%�bB�!R�ʡ`�\�j���;߱q�����)��!B�h��VZa
&���,JP�T�SU��Q1 ��aR���$��	$D�X� �cp"�$L�L�����{�ۭ���F>oЅa�W;<�מ����_4l��y�cM�o�0ӛ�F�eIy�y8�<��e|C�G4n�e����M�|��/ֲ�����y޿����N�/��ev�(�ܭ�U��/� H��5�n$����K��i�f_��}���U�����W;[V�]X�٭�\��6a��&sfs�����U�Wo>/��3�����	r��
��Y�˧�f#af=w�g�t!MV������ff
�	s1֔��Nh���)
p3w��d���p��q#\=�I�M^xiӯL��l�����l�·뭓�����2\	8�f���fKT��%�|�Q�B������c���պk6�	�K�B�]%��F<_I��#�'�M��I����f�9y0��0�9�{�톎s>5�,p4jq� �0a�+��n�&�Q�=C�?%,�����,_g�V]�]��;����sY�
V�#�f��W{g�I|��0�g;���N���Q:��������-��%j�
u�NR���k~}9ܵ2����)T|_�g8r�xxq�%�Ny�!��sHs����q%LbT"H��ĸ����H�w�#7�'���#���xx���.:[��n���L�%5u&�sm�۳�Y�$�<�k�����+��m<&�tI�Y����4n�Z6z=
ᭌ�)�![#bhXV^2�<���׼�<��/����9��yܲn�v>;hZ&ow�8�ggs��v�+)���T-U�+>���n��=�����y�a�<cS�G�S�l��o����aJV��7l��S`D���0�$��K
\�B,LR64"C�b�X�ŁBWL,bJ�Bč��U� !Yq%����!,��I(���YL;8yI��$BŻ8b;|�C���16��i7 ����x1B��7�߆��x抻8�o		�SVZ�R$H�BHaS �b%BkP�C!��6z�.��������_nd<��_v���m��3�.��ꍳw�U�2�
�]�|G+�����j�3�]೉�9�C�y��W^�y����6�3�<˹�_����ʺ*��8��"��U
�ޯ���0�/�����禖\�㵴w�ƻ�.�Nb���TWë�(�S���%(�G5鰗5���XR7�\��hd
d������e�D�� B��XR�`L�XVVP�&L7r��7Ŝ3FC��&�i�[ߢ�@��w�.�{��
�y'�KXV�ЗRp7�5.��GICR�JS��7}[i��bg�q�{v�p&f��o{�3��<�OM�m�1.���o%�0,�&���w�\�=�����P��nV�w���V�Bv�/T�2��������u�r_IB$#Isɞy� F$=ѽ��(U��ʟؾYήl�t���ma�p�c�[�s�L�y����s5̇����FY��z=�K9`��{l4d���p��L4��!��1tm���)�QN��(ɋ�n��n���U�T�ݮЖm�Nc��B��>�ow9ھ���I�B�/vs�]J��y�nmo�о���'8v��wj4u�B��)]�R� ��u�]|���h���*+�Ӽ��q���ߎWh�yE��ݾ�ނUBYx�9���]��ܾ���39]��}���v�Svw���ʛ�WI|R�)�t���%|*����3�Ը�i�R�mu5Y�];ڻ��ݮVя3�>����vkl�6�dB�.h���}����g�&������[!Q�"�"Leۭ]B��G<��<�3\�a1"D��(J��+
a)��$�qwG�m�L�.H�!�#c ����ޮ��og��=3g��.u����r�ġ��H��;���:,}�u�9\�����r�8�\�C��h��3�����;�����)r���B�Y\���}���ZKv��/���{\��W�no۔R���֯�vڬ�>�tv_���P����L�5㰗<�9�I7�/�Gˬ=�J]�ҺIR`E�XP10�vԅ����#b�v�.��9���|'O5�33�}����R�k��򯮘)ǊJa����r79|���zJdH'�	�%�3.����B��y�Y�M� K���`C�.i�C�F\�B��B���&�ܑ�W�ň�<��0�7�R���yA����yE*QV�\sn��9�y�Ba˭2�.0�X��� �[�=��Xo�������%� Ms��xf��.{�5Y�IL��*��_E}ʣ�ݺ���z��9k��/+��/]�P��3��:)���#��S39�q�<��<fl���\&p�ޘЊR��\	p!IsɣZ_2����6{CW^����8hن�֙sA(�dh@��(K�j4˜���|#q%�������.�)��\x�>�q�|Y|6��QH��(EЊaJ2�.d��\K���N&%�\BP�`F��Mh6�֝�dq���4 ��)F0��ˆ���
F�*8	�&<�L]&�p4�Ny�D+�2Hh�f]��a{B�=�[�f��7���)�����&����	G�3N�Ժ�ۤ��6g���,�$�j��7&!r�~��盔�7���%�?��I�%|+4%���^)%�R������~?>K)!�,Yi��e7Z���3�.�&��F�|?{�}�{�[In�`�k����2�&$..YE�r�}������߳:�U������\�Ta��l��՛�<�V^���s��h���ګ���Ϟ��sV�eo��7���N.��Xm/���g��q�s{�C7��as^�5�����d�l�d1.]�4@�Zy_e>I���ӯ���[Y\�3���efUf&
�X������F��f%^���0���[7��sҼi��Bu�S��U����fe��	BZ�q!aI4k��6a͙�D܍-aR	#Y	�����M�7��C'7�s�L)�%�.�nu�&*�m<������ U��r������\�w�̣W��|Vt.e�W��)�<��M�X�i�r�Iԅe�vK���u���rˆ��˽rf��xH��w��\8a��|�0�aCF���z��.�j>�4l�$��2��6�h@��3\�����:�i�s�4n�$���!tq�nf�t���A��q=OasZv���	w�Q��Ć���U�ąH��!4�!pbBT0�n��#hٳN������>��d���N�>>T��YK.�G�>��8ng9���Or�[9��7��2��=�xI(B�#�d��4�Дaq!P�7G,#L6D5 J�b@��
�A0t�*��4�v����
h7�pލ��,'Y��?UUUUUUUTUUUTTUAUUZ�MHEqS֍O ��6h˶M���s��[���=Ǝz�ٹ�%2��UҚs��v�����Ű�Ψ��zF��y���'p�$3��	�a��9�I�to��v�M�j��fU"���v��N�wf�m�!Ƨ+t ���<=*�XܽyE���Y��Z5P���#L�V,�� Ua"s���dўm�
�	��p��+MUW2յ��t�vtc�,T%Ad�6�FS��uV\�5�Q-�\J��(�����Pk��W�t�kV��M�y�m����W��7`�mp�į��*�s�R
��Mn8A���&0�z}�Α�Wh��-[\�l�ۣ�� �ܛ/��j���).�
�j�`�h��\����V��8\P5lI3�����jڷj�hʪ����)��,PԘ}b�
��RXS�c�U.u��l4�`�ݶ���f�{1T��� ��ں�(���}<�ۈ�:iI�꭪��S�67U9C��X�᜵��`*�%�<l$U�6��Gj�-�n x�\���@AKUU�*�QP���;��"U��*�kfkV�.'e�y���fh�1UG���5A��-����=�ټ���Vh��an���(-��pJ��$i���U�K�������a)MV$�PWm�R[��fEu$!,j��W�Keawe2�Pr;��[��x2)Ӻ�.����m�֋���J��vj�k�ۖɎ��5�ƃ�z������T�?
;ʼ��m���,���g�n)����=�)as�t�6n�:��J�I��X�4+a]34*���39i5	i#�B3 ���E�Z�#�-��ˀ�o�tftey�j{�'`�`�/�cH�mz5��e�V�W���B�c�cr�Vk�M]�X�אYq�*&Y�*;*�j2�lh�݋�O�����&��U�Qȩ	�L#�Qt��Ys�,ʪ�.��D�,LKd����CiL�Z�Ƃ�� �vn\�#X�IJ�Z�B5j���������_�]c	s�n��(�O#�Iۘxnr#�{u�3�m�Lg�f({J�e�+�^m��.S�=�眍�c>��]S����n6QL�nW�Sn��2��6�����m�IrCjuY�+]��s�4Ic�g�}S�!�мr`6�q	����NM�b�n!�;J�/5."ƚ�ɬs��86k��h-&nK�
�\k�4�6��[��4i-t�����l.ƅU-h��[�OJ�t��Ī�@,���cX��;i�ؠ�j�0+�qNg<��v��HU�
�����5uTy���+U�l�j��U[Ua��_\�����M�	�66�^�c)��bRڼ	��4XݯX��]�W5�GE�* �Rr�"U����`�d����f
��Ӏ�`'�]�����8���J��Q�mҠ9F����Zp��.W��U|�x�k���*���
Z��
��5�P宂�����
V�M�� <|��z���y�Ʈ��.�
�/����r��
�j����gA\je]b�y�釳��p���w2��R�TR+�Iu�Wdn�hT�0�TN�ͧ\[kUUWU[�Ğv�ޝ��-�jh��@sj�����*�]nա�hW�V���'U�Rl*�mUǊ	��#T�!qU��@����ml%��@6����Tb��me�Qp�č�s4(i����JJ���8A�L�R�`���V�B �@ы)��rͺ�p�1�٧v�%f���T���:��{a�ֳ۳��C�����D،C![����(�Y�YM<d���Bv��0g�IN�@��Q!�X:[Z��R��´7bh�����S�O TUl*�ѩS�f��TOmTSZ
�-,�lZf�x���b���1�޹N,���n��ƳM�����e%]Pa�͹n`�����UU@pG�*uZ�Uj�5Z���T�m�`�^ˬi���ݥ`
� �C�પ�Ѣ��\�������gO- �x�Y���Ӗڨ8�U���{lƮ� U�I�,J���yٚ�B�j���Du������g��W*�P��*UX����`�88^��������v�u����*�W�B[.��+MB��`b�b��APtԻ���U�g���L�]�:^.f�v�5�p+*�WUJ�W]%vD�J�$�=��� \]_U|`�u����^_U�<�Q̨�*�U��Q�b �b������f�R�UUUpM��\ǫ�E�rX�W�lp��S�&E�[�� +�P�UUlpUc

���>q��v���i3����*��(Hw-����U��uN궪-����U%�T�@�1=���w/]�����c�=���<J`���� D���j�UU($��`Aڭ�����In�SUԤ�*�R�
����L�U���5��j��,����P pl�5�Tj^э��p���yq���UU�@*�URUҭU*ԥ̝-R���Z���&����9�Ag����i�TD�Qvv� Uf)t.RE�ˆ�4P��W�V	,�,W�E��S�Kj�Ul�iyjU���V���i{j����n�Ut���UU����@UUV�UUUU��V�uWU��@O(UU:*�`�U����@�yU�+�X��P��U-J�V�b�OT;:Nj��0L�������`B����Vڨ
�P��;(i�[U�UU[+d#d���^���j�����u�8j��2�WUmUK�j����PppS�C*�PUUUUV� [U
�b�;TPUHE��Ԫ��ۭ�֨�U�Q�
���*�j�'d-�=K��������YV�*�UU��nI'=n�򍱴X����q����#&�mWmZ5P���;U&B�]UU]UT������u��
����@UK@R�PյU����-l]c��k.9R(.��20
����f���V�++���UcPQ�ܮi��j�W�v庪�V����'T��UUU@UU*�UR
������UU�[l�x����عV`��UZ��@A�R�Z���A��VʠR�2�V��UT�R�UUT����PUU]UUUR���C� ����j��Z��衺�5R�U�(�Y*�S�mJ�c�����>��r�c5T�vn�=��  �jU�:��䋓�K 9���U[���J�J�UUl��E�h�9��U���Ucs�Vm�2	�J7<N�k]���/���U���]���U�L�.��t���.��R�>�9�a�[�0{	j�.%���;k�h��*���k�eUX
�%+j@���
^Z����6T2�_*��T*�i��J�Skj���*�-�����UUݐ 6'P�fV)j��j���
���tTkL�:����ݸ^��J�V��˔�U��J�P��UV6HA{m[]Y��?����
��pNñMմ@K[�Z�;�Cd�9���u���V�$UUVQ�.�M�`:yZ�T������#B5����%�p]��ʶ�4��Q��.S�8�-�Z�u\�>��u=r��e� W�*��ݮ���q1b�c��F�Dn��q�x���k=T�����X˺m�UA�ʤF�1l�h��K�F������:����r��ڪ���t�&�P%ZU�g�3/�z����-����c`�:!�U��rKti�d[���o{ǀ)�F�@���:���)Un�ּ���痗`��[�]�`UX�ܺ\��O�L�'+�8���ڸ
��e.Z�5mO;L�U��L��8���q�*�@�X���oz�5�TL�´��`�U�UQ����Uuc8��^�� �M���Ysm���lV9�r ��9֤���(�+[UJr���j�]�UUu+F˱ ��l�"�������*��U��R�+��D�j9�p�$�mt�6�F"킓a��f�
B�X���M������R��P�.v���S����`EUC%��.y֓���[S��j�\�]�z�/56�]UJ�UV�HZ�j��˄�63E-T����������9q��ʄЪ���X ��3�h�L"�T2 *�jj�AUR�K٬N�vm�J�R�ˍK�f\�3����RYV��f�uiɫ�]��{O�; vu+�jn���� �ANd�+T�d�`��e���3�k�b���V���
-��
������"#���m���,&�q�dP�UM�Ii\�ꐔ���v�%��u�Hnּ�j�=3�d���[3��'!�$���d5�k'/I����j�Ji��UUUUUUhEwk�R���ې��*\�	OKc@�$����X*�y�G����H�cz4l�q�K�]��v�ŵ�ʴ�xɴ���ݑ�@]�;Q��ͣ�b�u�T�AnnX݆��s����6b:��n���n�FƄY��Sz���V���5�n��8��15�N����ոՌ*�R�K��nF�*��bٹ���lhMh� (��[UUB-�� ��	sUٮp#��!*�]��TU�h�[m��}��yZ������iV�m<�ګ�y'd)j����U������������+��R(�5�n+X�P�Z���[TUUUT���UT�:
�J��y �����Av�,UU�UX��*�UmUWU�٪�� UX�^@�h*�h��j 
�]�`)�u]J�TmlZ�j
%V
v孞�����_V͵yw#0�rˠ(b���穫kj�ڭ���[�d��+�S�M�UUUUUUK��UUU�m@���.u��d�‧�Ѫ:�%��6s�Arj6�_x'�m�$?�T��	PS�F��BA6��A��0P�D�#M�TJ?��d$  ���0D�
z`�� ؈��A6 � ��*4\)�P�RQp���BAСpT���H@�P���'���b:P6���� ń6� | U>P�_�8�Y b��+� �?*`��"|+����)�x�l6��y�(�8l_� ���{�'�+UH'��� 0Q &��]��華�"��Q> �iT�������~Tw�*<<J�E �T��������hWh��� z���� EH�HVĂ! �<_Q[����*+�<���U�C�h�	$�$! F1��D�X@����"�B	+ B$�@�F�!$�`�Q�P�@���(���� �e��b�R-��H��"@"�$	dIJZ��,H!$�!*��Uأ�b�#��!�{��@����R��	m�`�� m@�=t��P1D��+�⮑B�����*��~(.-h����> C�`
���?� ~��*E�8�aD
�`�C�����}�;L�nin��*o�vt� �^ڥ�Ý ��
�m]��KXh�b��c�7E�H����2vi���(��,��@���d� hI�N2�v숛;W���m�A�tXaP�싋�`�ͤv��hgj��2�j�*�n����`�@��{���-�e8��.à�M��vɊz��5c�1�r۔y�GvyM��<t��M�k+��
���F���s5�/6lZ��)��N�F�q��2��.]�\���J2n��:D�OEe{[x�(m�E��.���dn�z �����G�<��dt#�9��5%���.�4\ʤ�T�[@t��Sխ�n�m"[�v��6��C	4+F2�u�F�j����Х�H��5��6	Y��͠$%�ūdQW�Wv|���#�H-�8�p��^J��#�
�K�4h��ܬ-��Jk�1R����:c@{4i`&��]�uSj�#-+t�m�lr��7b��`	�Hf���fc��Z��2�6�]�%��X��'���O-h�Փ�9���l��\�a^�&t��r�e
����#a�m�ȵ=�+Yz*5��YQ�0�#+�3/l�ǰ���1�]283��1b�L���c�]!]�*�m�Y���"Y��Tͤ���V����c�i�y޷Vֺ��"W��q��Gm.ݱ�-�0�6.��6\�f`�Q�:�*=�v &N�9ˀQ$�îX8�y|W��I����K��@�n֎5i�AB.�4�ЖWlcJ�\93��x8��gent�� �`aT����q�nm�+��
�FS^Y��������HDR�ٌ���W(�;u�JN�f�Jc 27�YE9��Vn{qɦ�&�$��6��m(�Uk���f0�th��=u���fmM�`�=	f��0�ZՖ�ҕ��z큹B��t��N�����du+pv�-Vu658B��cv�k��.��L��\�n��x�nu��\�l-��\�2�{��>U 5�A:8��(�� �'�?�|�§�&��t�N��wO�����t"����*u�-���k��Sůhx���-h�jt�c<�NI�	 Q'���s�p#�>��q�9��lg�T��`��vN�8��$�Mu�ƷJ�ɸ�,��N�G�����:!�zk3���&�<�dl;�'&z�q��O s^Қ�(%@���Q�5�4H��!�i��ʍU�0]qT3:=�'N������_Ox�K��)����f��������C`ܫ�es�]�_�J�]���M�f͙X��`n�u���������=B60wM���8�K�}�G�~�T���L��P�Z�i&�ZlV� ��w�un��9$��8�K�'n����ݶ�ZM��:�e��e`[%�\��WbbW+��ݫh�w�rI��ql��I{�[��T�J���I�Y\��Z%��.Bnړ5&0��Y]�T�
CM3/ ���=��π_���	/c��v^7fV����CmYwi�ݻ�;/c��ܔPB
	�JI	$�"%L�ڕ_R"���9�2�.�x$jR�
�I�-�v��:���	�2��][�^���X���պvS�Cn�	6e`]����XWv^ l�I��64۬��^�k ����$ٕ�z��b�此�41*�v�&nY�s���c'=����d�^ͺ w�L�`��ht��)��lV�o��f�ݗ�I�+ �엀w�HЍ��]+v�Zv��:�%�l��:�%��Ƴޓ�Z{�~�Ƕ���w�{��vnI���s���H�ŭU�A��޾�\�ܓ��f��OJ�)�V?��M���/ �5�uvK�$ٕ�s����Mج�m����k �엀I�+ �엀�[��*k���a1�pךOu���'=�"C���6�^:�dauԱp�`���f���/ �fV��/ �5�n��][�e�wlw�I�+=�}_$j�z�������x�bLt��e��l�:�%�/c�=�}�Z�޼���!Դ7t�n��]��6^��ܓ���f�y�~"�E"1`�J*0J'ʎ}�oy�'��g��Z���n��ۼ��^;�Wd�e�w�rk���Wc���$�,6��k�e֢��K�= ��Wj���3w@m����bVЭ�;�Wd�e�w視�V�׀v�C�{����m�Wd�e�w�uvK�'u� �j)�(MЬB�˻w�l�����xy/H�`�޼f�)7B��������U}Ko}��=#�uvK�;/c�v����5i��n�	��uvK�;/c��l��S��|#�;����3��pvr��u�5�B0��I�6[��u��:�D����jn�q���ҍ���k)1V	.�hF��)e�v��2�!Xe��c;�ۥ)qt�L���L�]�sä�9$q,��^�6Qm*1s���5��68�3N�8�Om�筶�����ֆy�<�����iv�8귱��%�����3ݴs��㮘Y{fLy�������Y�I1<_vV�4cPv!�zl^��K��I�\�- ^0v@�֐�+�Z��#��L�r}�������� �/ ���IԴ4�`7J�.�����~���H����=#�j엀wn�����mۦ�m��6^7\0]����� �ԀvR����7eۼ/I�0�޼��;�:���9�����U��V�Wd���;�:���&�꯾�{��Y��GMD8n�,1\�6V$˵u-��Xa�pj^�Z{PĎ�'�٠���v�o�y���/ ��������V�׀OF�M�R`:e�.�n����f�︉��$(�a%sE�5t�GD�E-d�,a
h�p�ud���\�;OT"*g_)�xe�w�nܔ?�����M0V� �{��/ 콎���x�IB���n�lv�X����[{�^���xWd�m�Xv$�i��St����ٮ5�uvK�&�ŀuvK��(CiҷV�j�N\�2ks3�ƪ��˷En\���sk�lq���=
��wV����i�k �엀M�� �엀vk�`���J-� Mح�6�,��^ٮ5�uvK�9�mH��Ż,vճ �엀v{��w7�"� �!8�{[�+�9��vG���`һt�ح�ݻ�;5ư��x�p�:�%�/T�lT��컶��:�%�u� �엀vk�`���E���fZk���2c�y.�M�^��#04,��URar�\�f�+*e-3����^^�uvK�;5ư��x�IB���n�66�Wd���_$o��X��� ��v$���n��]��;5ư��x�p�:�%�Z#Be�E]��Ӷ���/ ��W�}��@��	�M��}����'>������n�n�	��z������o��X{r,�4]+Te��ݥ�sB�&&��v���5�6�f-M��b�t�)���R�3z��y�n����;ۑ`u� �`�U��ݖƕ�;�xf���܋ ��Wd�f�N����ӻ.���X�p�:�%�����rSE]�V��ӻ��	��uvK�;/c���^ l�RM$�M�'M�ـuvK�;/c���^7\0�~_}�R�����j�IA�`�\9d	vMTMU�c��	n��P�Z�m�'M�2,��ӀwcpӸ�		t�O%�r[����ڂvd�K��zT�l���wZ�=`�+8ޡ�K�,f9��n7#��;QOmvr2�TAm�y�ϒ�!�=����,Դ�Dpl٢�cz�j�Hz�;ln��01���$F^�jXMoE�%�(q��ȣ��++j|��sӤ=�_0���@�-����\9�4҅�v�k�v[�E��6z�������"��Wk�|~�����/ ��Wd� �hD��vR�t�v��:�%�u� �엀vk�`���"���݊��u� �엀vk�`]��m@�W)���;jـuvK�;5Ƴ�%۹�I)���K��M�y���ٛ��{���<78n�Jn�9Ēճ*�$�:E9v�v�M�u78�n�%S��:�Y���%��ԣ�9�'S����V���1,��vʝ���:�v�~���9�m�����(�3-����W��s���E�mi�� 9�r�Ξ��`@@ K~���ݶ�{����`yw@�zr+�b���Ijٕx�K��w�$�Tp�I%7s���9�
p* ¬2ݙ� <��8�]Q��$���s�%�L�ĒK���^ڳ[�����t M܇8�Z�ʼI%ٹ�K�UU�0W���H:b����2���R�e�g�q��m�<r��S��BQ	a�P̍��dݤ����I-Q��$�f�k�I-W"�����o@nk�Υ�3{�ӏ.�W�wio�y�q$��y^$���s�}U{��u�n�G*ܵ37@�s���[o�>����>n�f��8ss2�|L4��9L�B���B�S^�~�8<6�)���}b�׎��n���NR�?4<3��l�#wIzg�lK	'��%���(�ᤀ�9�m�qcb},�.@�=-]�w������������nG���_B���3['��y�g���x�$.��绛	3��G|"<��'���t�������M��$�4:�0�'$^�֦��̫�.N������	-)8h�5�	�V��BG\I�%�2���-�TĘ��H�Ê<�!�S{��foDɬ	u9�h�곜�,�J�?���.$��!�7Z�-�]�����h#i]l��	4]h3͉���h۩gG��A6S�%%��8� ��b��@|"��x	��� @�H�$HH�a#,&��C�)Kpp@M��O�B �+�U_V�gNq$�lʼI%�L�ӢfSv�eN� ��� 9�r�ؒճ*�%������Ny�q$����,�s	�Ŧn� ����`�� <���q$����I)�1Z��V��t�8R�[a��n9�@Ӈu�,�\�V���f�7O3Q��Kk3�����:��ٹ�K�8_���v�����$���C�Ѷ,2�3t {�z�w���^$��܇8�Z�ʼ�]�JD�G��Jښ(�;��}�� �޹{��L�Ē[7#\�I)?�ϛv6�+wx�Ju�\�Ij�*�$����8���z��@`���$`��E��<� �Vk���ݶ�>+_���Zms�%�L�Ē[��Ӟ;Ԓ���x�Ko��Ko�㤛�Vs��`H	'g�w%�Ɓ9.5��+�ntt{%g���L0��f6-��-L���܍s�%��W�$�^��$��2�A�=��h�1��6U������	%;�q$�lʼI%��w�$��:.�9%���8� ����`��I%��w�$�cq,I$��(`�`��g+{���u7@�}���/��{�/}�sk�p*%b�n̼I%��w�$����g��I/l��Ij�홻m�a��g̢A����o֓Lyo(fb���Y� �ە���r�<[�X�[�F.��Ӫ�H� @���׮d;h*�]����'0�N"�f{cf�"N��z2��t�5���۱��;�2'#d�x�)�i;�}�]��; ��pQY?@��'Ʈ� 8x��V��l��Z���:���X]�����L�@Mu��n�x��Hkh熻���̗�Mh�[r��2��}f�Kɖp����0�-��|ᯃ4�� �Rכ�`ĺ]5�&LЋc4cB���b4PWw�8ߒĒS���KT�W�$�=��Ē\�[Fr�&]\� �޹{�T�W�$�=��Ē��KIshߊ�]9"�]���`��St {��;��[�bI)��s�%݂ş2��Bn�cV��$����8�[-�bI)��s��9�� s���+k�j�l��i%��$��UU_W�s�z�Q{�W�$��q;� �ou�i�m�n�:�:��=���&,9�DM��m�t��N��j�.�j˱!+bĒS���KV̫��=���~��~��� �}����K�M�ֵ9�m����߈��%T��ϯ[&k\�Iv[�ĒS���=_U~��>�����m�vf� ����Ē��$�w!�$���W�$��/���ˌcE�}�xq�� �r�Ijٕx�Kc��I%5 �M�9�ɺ 9�r�����n��c�q$��Ex�K��UV����u�%`�x�ǫD�cbn�nK�<cZj���j{L����f.+"�]���9�R�$�Ǳ�8�]W"�I%;�q$��[����*�5ٛ��>�����I)��s�%�fU�I)��*��6U����t s�z������H�+ n-h�Ichdd"P"A$XA#��r	 �<"�9�����m����g9m��u��V�-�h웠?�o��^� �Ϻ���>������� >�s}�����U����:���������vw���������[o�QΚ��S55l��ݯ3�.��sG<dleQ���\�z�a���?��W��J��֡��������s�%ێZĒSw!���QOe^$��|)\���G)�`m�mת��/I�9Ē�{*�$�f�k��Uݥ�����k����� s�}{�ճ+ ���8�K�9�m �h�M�˶��wfVٮ5�snE����`$`�h)��g�s���',�]:n�c�;�Xf��͹7fV�ٕ�~���t�ג�6�4��QZ�.��hM�lP;��v:�c���f�s�X�ٚ$������S�o��|`ve`ݙXf���ٔ�һtt�]��Mٕ�����X�?5�snE�E6�$�v튝:�ݺ�;�2��q�=Iv_��I�(DAZ��;lM�f���$�n̬?/�}UW�{?^){�m�6
Һm;m`~�۞������������ʞ�~8}��&}TQ�����)j��.E�xJka�X[��.:7vi�sk���,�b��"�a���	eč�� �Ŏ����ƺ��a&���e��m����*M�\���Jh���k���\v���m!��Ns���<�ƍ��i��b10l���Ip��G9�ܪ�\4���4LYfֽ�Ԍ�� 献��q�:�i^����C���e^!6�+nv��]���P��O�t��bx�2���<<�1p$	��%�!u�s�7>^�����$��g_Y|_jPB�����?��g��G��qT�����J�K�|�,�m� ���RG}��:��x{�K���r�;��X��$��m��0}]��5�:��x���"��?^��}ϷP�pի���_~�������_�~���?���U.�g����=�t�e�M&�"ջ�=<�`��<p�?5�qI/ �dD��c�`pLv:٦�k���i�Eq��]����v"5�Q~��7[�

��3.�ݷ����95ư)%�u� ��Ri]��Z�*������w�$��KМH�I`z�FLF	B�,�!$4�-F�57�/fNw7�����7veg��P�<[hM�U��i�k ��X�p�Ԕ��X�?5��K"��e��]����L�I=��wuư=T�~�� �QC<��)�V��l�7ve`�d�5�:��^�{$�R����$��Iٻ\-	M/;mPL�Q�͉;ZlHs
:����YHv����v�n��-����^���d�V=�^R��n���ڵm��ql����6\��6Oe`��{�H��e;)�i�6��ջ�6\��'������)�P�D�`QA0C��@!���;�:����"�r�n��ln�;v����|�Or���;�8�K���/G<�*��*M+�j��m��`������z���,��+ ;��\7m	l�u.nŀ��ņLJJ�D{;M)���Ɗ���:x;{��۩��*|���{׀M��ٕ������(�y��t4+wi[�mȳ�_$l���;�w�qI/=_$�J*�M6�]�m`Oe`�������Uޯ߿^�ߟ� ��N Wl�-�m�ݺ���}K�s����^68`J�����՘b��� ���@n���'ݟw7A�4,n�ʻ�>_��o �wN���߽��.�=��X%�w�l�1��][��疶¯^����0l�;�,�ӳ��[���r��I�"�ƯF������wc��{���� �=��z@EA�c6vN��{Ǘ��~�'�}s��S޼mȳ�UW�U�y*Wt;I��-� �y�ղ^�ﾤ�/�X�?6�[R�ӤӷN�m���
~Ts�w��ܓ�s��'���������~}���������k��Y�.���}�{�ܓ�~��?O$�~���nI���rA=�N}Ё L�|8l9jP��B:JB7��,�N��###a�0dX1 LB%B5�T"����B$@�#�H1�����B�5V�$�[	��N��� XFJK���Mj\IAp8KzӋ~y7��twǋ>i���AC��6�Ww�BZ�b�I#������Bq��.���@!`1�% FRT�"��J,+
9�V4{,�#=-'W�`�z�B$c�ZF0$�����\�G.1��V#�"�!A!A�B1�HQ��^q`_uD��a	'��$4��Hē�r�r`拚��������j*^H�1$H�I<@�����x�r훘َ��`lפ�f�_T�F�!� I���g����O!�6B'$b�a!� E�`aѵ��F$"I$a	H�$��#"H0��)`s���$$RFH�Dw�㎆_�i)y����ִ{�A���,#'wc��wi!̳BO�{��V 8�x99�Uφ�-k�l����9خ��[u�xq�I�4c:��qD[�ܷ�x�&{QF�x�S<:�pf6�եEV��&�1,+f"Yu�#aT��K�6�C�����FN`���@��`Ws�IV�.�qBV �Լ����R5�,�6�^7��'���.�tP�-7Kpc۵�Z���3���Q��v3�K�λJ�탯hh���2��Gh�Ŏɍ�Z�nl���1�+5��6�b��1��`�4L���CK熰<O��.���:9���=�;Nh�� nF۪�3���.�0$a�IAݥ'��e��ӛ���L���Ũ�%Y[k�e�f#eU4���x8�
r�nNN.�f��ܘC�2.y�%klͤ��m�&��9�2V��Ԙ(<�4�����I��Ƿ3n)�nɋ-��64lE�$ddް����d�pwl[3˶�ø�����$����4]5,��#)�t�o���2ԭډ-�%u�lX�ۓ[g���k1O "&��t�q
�Dpb�"��լ�p�綠kk�s:�Gl3��D��[����9Q��S�:�X2.�:�`$�˛�K�cm�,�ͪr� nk��3u��͏Z�\�c���m6��Ξ̑�MRT��^X���e�΄��\p�3�E��\+�M�Ur�6��Z:��L�1	������E��]p�J�K[��[�03�����2aƖ ��ql�3�j�ݺ��d`Ž��R��7	645��nc�t^�v_2��� ���9�3l��� �bh:ظW.�].J���Xn���U��LF3wI��<Lb�H��C.��e'(�x ����7	`9�p����k6 'kR���M���	7\٪g	�pE1XFj�CfkP�n(�ruͮ{���H�VYbLW89SK�K*���-l�l��nڸ�GR7�����5f��`��VmP�t.���Ll)>f��겗���Ͳts"ln3m�9#t�����*��:^�G-l��q�|��]�@5UD�xtT�¿ ����S� �Q�O~#��?�C#���ͭkH�KI�1�"R��lr�Dv��)�6c-z��B{{[&����U�®V��SGWI�*"�G�����71z�휯�S^�����M�x���.�	ez�A��e��sp��E-�v�qΪ�2ʄ(�.jF �5q����y]���;^a�M���10�jcD���]�9E6ޘ�:B�a1n-�I�ְ�.��I��__��sg)'����!�b�46�m�l��K�'��(v�#�3Q��c�'K�VYK}��SkN����� 콎��%��靖=.y`k�ؐ��'M:m�����;�W�}I��^�s� ݎ���H�=��C��HTէwm��j��x�ذ�}_��������O���9$�l�e������������~0�q���%���������Z��s���n���W��k�j��x�p��9�*�i�%f�i`�PZAa.��HZ"�.�R 36�Zh\j.#��:OL{i�v
���8�?5��Gշ�z����(�%�߾�f��"dK��o��r%�bX�wM��0��D��h�]f�v��bX�'���6��SB�+$Q)	Ya�M�X�@�`B-� �HaCJ$���&��}�ND�,K�{�ͧ"X�%��~�uv��� �DȖ%��{l��,��`Ot�zk�^�������r%�bX�}���9�ı=���ӑ,K����nӑ,Kľ|���jG[�ry��ҝ)��)���ݧ"X�%��~�uv��bX�'��{v��bX��dO��?M�#)ҝ)����y�qW8f�.o�>	bX�'��}��r%�bX"��w�iȖ%�bw�ٴ�Kı>�]��O�Jt�Jt��{}�&j��&U�We��rny7)�I��H�:	��솆{K�p������K���W����+����MzX��]��r%�bX����m9ı,O��{v� �DȖ%��u�����t�Jt�O������83��ҹ�t�Kı=����r*�bX�}���9ı,O~���m9ı,O~�{v���X�%�{߯Ku�]XkPљ�kSiȖ%�b{��۴�Kı=��iȖ5�B��"X�k���r%�bX����m9ı,K���Kfai�Mf�35��K�ȫ"}�}���r%�bX�w��M�"X�%�߾�fӑ,K!�����<:@�n���ma�1֫�� �'����pIC�}��iؖ%�b{�{ͧ"X�%��u�u�ND�,�N���'�rJ���b�G]�j�i2�1�QApSg�&�U��1���I#�m�s5�˚̙��ND�,K�}�ͧ"X�%����6��bX�'����l@9ı,O{���9ı,K����÷WV����f�ӑ,K�����NE �,K����6��bX�'���6��bX�'~�ݻNA �,K��zy�.*����:|:S�:S�����6��bX�'��{�ND�@,K�k�ݧ"X�%����6��bX�����w�����9w�>)ҟ��D�]��6��bX�'�뿮ӑ,K�����ND�,� (�<6�� �(H����k6��bX������&y���F���å:S��k��ND�,K�AT�����<�bX�'����ͧ"X�%��}��ӑ��N������{X�m3�r�m�q��{`�+���SyG��P��ͣ�P�$zI��o&�C[��l��:|:S�:S��Ͼݧ"X�%��u�u�ND�,K����� �Kı;��۴�Kı�����ٮ�e2�o�>)ҝ)ǝ���m9�"dK��fӑ,K���~�v��bX�'�k��NA'Jt�Jt����=��fr���:r%�bX���w6��bX�'~�{v��` X�'�k��ND�,K���Ο��N���{m?_snsz��k��r%�` X��_v�9ı,O>�{v��bX�'����m9İ�=Ͼ�m9ı,K�����ˬ�.��u����Kı<�]��r%�bX~F~�k6�D�,K��fӑ,K�����iȖ%�bq����g�l�V��,
aЎ��%��,�J8餸�u�k5��M
���]ͨ�n�A�fՌB�c�P�jVjQ�A�݊<��v��حG�����ve��7��uo:X+T*�[3��
��.�	��ݹ��#C����\;����g�Z�n�6��9�A�c�c���H�f�L�- ���#��I��oR�6Ī������R�0���]/I$�;�D|e�I��ĻT�Y����!mu�*%�ش�q��a0\��3O���J�ڄ�:���t�Kı;�w�WiȖ%�b{�}��r%�bX��_v�P�Kı<�]��å:S�:~�������Q�.�uv��bX�'���ͧ"X�%�ߵ�nӑ,K���w�iȖ%�b{߷�|��IN��N�����lpg���ֵv��bX�'~�{v��bX�'�k��ND��,O;�����Kı=Ͼ�m9ı,K�{ze�335�h�ֵ���K����w�iȖ%�b{߷�]�"X�%��}�siȖ%��'~�ݻND�,K�=�S�\�[�Z�Z��]�"X�%���uv��bX��Q"����ٴ�%�bX��~�ND�,Kϵ�ݧ"X�%�|�ӗ�Wh-���]O��+M�#2��0=�V)��X`���Z�F1���>���kFZ�֥��j�<�bX�'���ͧ"X�%����nӑ,K���w�`��bX�'��}��r%�bX��e����֮kFeֵ�u��r%�bX�}���9�"�+��%���ݧ"X�%���uv��bX�'���ͧ"H���zk�~}�����s�p.�O���bX��߿fӑ,K��o��ND�@�,O���m9ı,N���m9:S�:S���z{�ݮ�J�Uj�:|�bX�؞w��WiȖ%�b}��siȖ%�bw���ӑ,K��=���O�Jt�Jt������æ�.Weֵv��bX�'���6��bX�'~�xm9ı,O���m9ı,O;�����Kı/�{���5���-�Q�v�YV��(ۍYM�g[�^���$��عMUY�cl�fs3Ti���O���bX�����Kı>�����Kı<�����,K��;�����N��N�߾�f��m�`sVyӑ,K��;��ӐAKı<���ӑ,K��;��ӑ,K�����  �%�b_���t˙�ܺԺ.f�iȖ%�by߷�]�"X�%��w�ͧ"X�i�dQ�$T�t��]��2&D����"X�%��w��ӑ,K��>���3j��[�O�Jt��Ӻ�?n����Kı;�{�iȖ%�b}��siȖ%�
؞w��WiȖ%�N������QnYu\ڻΟ��N,N����r%�bX"'���6��bX�'��}��r%�bX�g{��r%:S�:}�����eZZ�]3&��
"���Z����]2�%1��m6vjZ4a)`�e��Y5u�Ѵ�Kı>�����Kı<���ӑ,K��;��� �Kı;�{�iȖ%�by�;~�k
�Wy��ҝ)ҝ?����r �bX�w]��r%�bX�����Kı>�����O�D�/Mz~���O�T����O�,K���~�v��bX�'~��6��`�bX�g{��r%�bX����W}>)ҝ)���{�k4̣��V���bX؝����r%�bX�g{��r%�bX����WiȖ%��4 &�4���U2'o�ӑ,Kޛ��ߥ2G�fkQF{���^���>�����Kı=���ӑ,K����nӑ,K���w�ӑ,K�?�N�������f:�&JX�"<��x���a��m�Xm��5V�;���ok��ܺ����k6�D�,K����]�"X�%��u�ݧ"X�%�߾����bX�'���6��bX�'��/ݚ�۴]���t�t�Jt�O޾�|NDBı,N��xm9ı,O���m9ı,O{�����OʤȘ�N������c�]�J�Ο��ı?w��m9ı,O���m9�[���o��ND�,K��{�ND�Jt�K���XOb7\��uY�O�%���u�ݧ"X�%��u�u�ND�,K��{�ND�,K�}�gå:S�:}���ˍ�*+|ND�,K����6��bX� ���6��bX�'~��6��bX�'��{v��bX�&#� G���50�-�P
�۲<�q���WZ�Ws����\O�Gv�
���.h^�����ϕNJ�2�������Yf��)��ׯQj�dmPa��×��E�ܼ�,��f�y\�n{'0���z|��^���P����e��g�n�Ɠuj��FihY��JҔ��Me]B`�,�uM*�\ZZ���)B�n��ч0ib�S&�zf\��&^���+�p��\��]Y�B�m�`���.�v̨�]�!Ah��z^:�b�t���t�<�=4Gl�;"��|�5�X����ND�,K��xm9ı,O�����Kı<��fӑ)ҝ)���{�k4̭Ѡ��t�t�,K��xm9[ı>�۴�Kı<��fӑ,K��;��ӇJt�Jt����j�(�t�ı,O����9ı,O;��Y��Kı>�����Kı;�{��O�Jt�Jt�����[�����]��r%�`'��}��r%�bX�g{��r%�bX�����K��T"w_�~ͧ"X�%��v��!���Ȼ�>^��צ�?������Kı ^����r%�bX�g{��r%�bX�w��WiȖ%�b_9�Ƈ�un,Ѻc$G
:Gi�l^�S�"+=r�Fڻ.����Z�h�GK�6�WY��r%�bX�����Kı=�۴�Kı<����9ı,O���6��bX�%�߉HwRk2�Y����Ѵ�Kı=�۴�<���DJBA��n�M[ ��P���h �J�YH8j�ؘE�A]�D�]�����bX��o��ӑ,K��?}�6��bX�'~�xm9Jt�Jt��Ox��2��Ο�%�by߷�]�"X�%��}��ӑ,(�@2&D�����Kı>��߮ӑ,K������hˣZ��k2�Z�ND�,K���ͧ"X�%�߾��"X�%��u�ݧ"X� *��~�uv��bX�'��}�#6�F�Wy��ҝ)ҝ=���M�"X�%� ��{v��bX�'����m9ı,O���m9ı,�������^��:\���3�.���0���6��ь�B�s]Z����;�Wϵ4L�ɨeT�å:S�:~����O�Kı=��iȖ%�b}��sh �bX�'~�}�ND�,K�=�;��h]Z�ͳ|���N��N�}���r%�bX�g{��r%�bX����m9ı,O����9�ȅ�M���}� Sp9�{���T�,N��߳iȖ%�bw�ٴ�K��|K7u���$�f�ć�u%��!c @ Ѕ)"F,#$��	�d�o1�"�e�\'��a���-�-�-C|!��<�n��i�fL�f�Kɠ��$E�$v�k��kA_��#����@�"g=�)����0�A����wo<����O�a!7n�ۄJH$�$B0 ܶL+�a	�h��ܑ"��!���}�m,K�))!"H�^%�ۜ�tKuL�c�=��d!"DѺH��{��.$�}|X�	64�;�K�G�<�� �m���h�	bR&[�X҃B$<�l4�B Ĝb����ӆ"���D�_D�P���x��x�� h��� � �=CGڈt��k�]�"X�%��o��ND�,K�~��_X0�9˛Wy��ҝ)��%�߾�fӑ,K����nӑ,K���o��ND�,K��{�ND�)ҝ/߿�a7��suջf���ҝ,K�뽻ND�,K�����9ı,O���m9ı,N����9�)ҝ=��g�M�B��,fC�b���P2�ZB2�م��k[�rb��I$�`���Ι�U·Ο��N���߷�]�"X�%��w�ͧ"X�%�ߵ�݇� ��"X�'k����Mzk�����|�#�:�]�9ı,O���m9ı,N����9ı,O����9ı,O;�����Uı<���]SFd4ja�&���ND�,K�k��ND�,K�뽻ND���"dOw�v��bX�'s��ٴ�Kı/��l�YsP�2ɚ�kWiȖ%��X�w]��r%�bX����WiȖ%�b}��siȖ%�S�H@BDYb�y�'~�;v��bX�%����nkE5�]]h��]�"X�%��~�uv��bX�"	�w�ͧ"X�%�ߵ�nӑ,K����nӑ,K���}���?AB0�7�kا��4�WW�Aq�خm�g�v�P�ϝ'w_R��&��dCduv�D�,K�����r%�bX��_v�9ı,O����9ı,O{�����Kı/�[>��5u3\�k5n��ND�,K�k�ݧ"X�%��u�ݧ"X�%��~�uv��bX�'���6���bX���)�u�sW.]\���r%�bX�w]��r%�bX����WiȖ6%��w�ͧ"X�%��u�nӑ,K���vnw&���U�t�t�J����t��?��9ı,N�~ͧ"X�%��u�ݧ"X�%��u�ݧ"X�%��ϻ��80msu]|���N��N�����r%�bX~�}��]��,K���_�]�"X�%���o�v��bX�����}C�}8��L�X�\����x�V����CIk���5��n���ȹ�H�0��s.� �ږ[��$u56/Wk45Ք���7.��Fu	�U0�)��,#W�%ڔ\j$b�����ݺ�5q��F6�ga1�:�=iF6�ۢ�ǰtǇ���e��me�^x:����ʁ����
�S:���k�4Xa�Hp��f#~I��;�1�6�h��L�WZl��v5̡� ��;[����ݦ.J;h�ȸ�;�>�
Ja�	���r%�bX��k���ND�,K��{v��bX�'�����r%�bX��۴�Kı/��l�YsP�2ə��]�"X�%��뽻N@ı>���.ӑ,K��u�ݧ"X�%��u�ݧ !bX�%����r�CU��o�>)ҝ)����{��9ı,N�]��r%�6%��u�ݧ"X�%��뽻ND�,K�	��6Ը(��s��>)ҝ)����"X�%��u�ݧ"X�%��뽻ND�,�>���.ӑ,Kľ}i��T��6����å:S�:}����r%�bX)�뽻ND�,K�~�r�9ı,N�{��r%�bXϹ/-�b�{BR���c��`�)�9Ƥ��[.À\�Q�z�4�:���H˗Y�֦ӑ,K��u�ݧ"X�%���o��9ı,N�]�ڇ"X�%��u�ݧ"X�%���nw&]e�kD.kSZ��r%�bX�}�����(��$�Z!?�мE^ X�%����}v��bX�'�뿮ӑ,K��u�ݧ"X�%��ϻ�)�G��k��O�Jt�Jt���Ο,K����nӑ,A�,O���m9ı,O>��ͧ"X�%��~�e�S4�j[�O�Jt�$'IN�}��M�$���6$�H��߳I�$���u�ݧ"X�%�|�{d�e�e�2ٚ�f�ӑ,K��;��ӑ,K��w9��Kı>�۴�Kı;��۴�Kı>����ѫ�彮����Ps�m�d^"����t�cVS_﹞�%žbE�>ww����Psh��0'����bX���ӛND�,K�뽻ND�,K�}�@�Kı>�����e:S�:_�~���m�F���>X�%��u�ݧ"X�%�߾��"X�%��w�ͧ"X�%��~��Ӑ�)ҝ)��~��o�\����V�ӑ,K���w�ӑ,K��;��ӑ,�p"�p��bxx��,O�k���r%�bX�{��]�"X�%����tɆk.f]f]h�r%�bX������Kı>�_v]�"X�%��뽻ND�,�=����O�Jt�Jt������6˪�"X�%������9ı,P�u�ݧ"X�%��~�fӑ,K��w�w�>)ҝ)���~��J��9X��Fu��� ]k]��f�L�A�9���!�����`ִT�t�t�Jt��۴�Kı=����r%�bX�ϻ��~ �DȖ%�ߵ���9�צ�?>��ڑ�L�hk(��>^���,O=��6��6%�bw>�siȖ%�b{��v��bX�'��{v��N��N���}�l�Aƴ�*y���ı,O���6��bX�'�뽗iȖ"�%��u�ݧ"X�%���fӇJt�Jt����˦Ѩ8�2��:r%�`�b{��v��bX�'��{v��bX�'��}�ND�,]�D�P��w7��ӑ,KĽ�w�n�[�hܗΟ��N�����o�Ȗ%�`���fӑ,K��>�siȖ%�b{��v��bX�'�M{����k7�0\�^Gq�-V��V�]�N�u.x�n����=�����.�Z�K�]�"X�%���fӑ,K��>�siȖ%�b{��v�	�L�bX�~���iȖ%�b}�IHo?s	�.M���r%�bX�g��m9ȁ2&D�>�_�K��Kı>��߮ӑ,K����iȟ�H���:S������k�)-��;Ο�%�b}��~�iȖ%�b{�w�iȖ%�by�wٴ�Kı>ϻ��r%:S�:~�����3G=b��R���ŉb��u�ݧ"X�%���fӑ,K��>�siȖ%��*�O����|���N��N�Ͽ���	���r%�bX�{��m9ı,?+뿿f�Ȗ%�b}��~�iȖ%�b{�w�iȖ%�bq}D �l@, %5��C��G���M.���'�LX,.6��ٚҜT�q�n��VQ� .&�Ֆ�jْ�Rm*�c�&�ݶ�[.חq��h�±�� ����CLk�ټ�K�i��,� �6d���Nڅ�`���@홖}��B��#����iλ�X��d�2q:�N2�녻�ݞ�N�=� ���HgGQ�C�ݣV���e�"��U�R=G �%e7ޏw~�N�>��<8�Yw�Fn��HM��<<[a�$�r񵷝-���ă�:}�k`�\�ja֦ӑ,K��?w�m9ı,O}�{.ӑ,K����nӑ,K���|��å:S�:_������5�-R��m9ı,O}�{.ӐVı,N����9ı,O=��6��bX�'s��6���bX��v}ٚ��E�Y�5sR�9ı,N����9ı,O=��6��bX�'s��6��bX�'�뽗iȖ%�b_=�v^��3R��Xj�WiȖ%��'���6��bX�'s��6��bX�'�뽗iȖ%�� b�?w�]�"X�%����P<�0��h�֬�å:S���{�ND�,K���˴�Kı;��۴�Kı;����Kķ�9x>�K�h����jc�&	R|a��g��rA�C��:VY�t�`����
[E���å:S�:{���|���bX�'~�{v��bX�'~�}��(�_"dK�����6��bX�'g߿wɣ0Ԅ]��w�|�5�Mx���nӐ�PJ*�Ȗ%�߾�fӑ,K��}��ӑ,K�����9ı<��][�a3Z�ND�,K�k��ND�,K��{�ND�����?w]�.ӑ,K���~�v��bX�%��L�՚�4[fkY��ND�,T,N���m9ı,N���.ӑ,K����nӑ,K�k��ND�,K����՚�vF����å:S�:{���|��Kİ� ǿ�s��yı,O����iȖ%�b}��siȖ%�b_=)�I�-�2cU�u�\���p�wm�rU�����5�F1�������͘��5f�j]�"X�%��{�ͧ"X�%��u�ݧ"X�%��w�ͧ"X�%������9ı,K�����]Y0Թu�ɬ��r%�bX��]��r"%�b}�w���Kı>�_v]�"X�%��{�ͧ bX�'��JC�ֵΎ����:|:S�:S����w�>X�%������9�`�HDiB$
�FF@�@� �D�0��ƤE�q@�"r&���ӑ,K���_~�gå:S�:{�����3-��f���bX�X��_v]�"X�%��o�iȖ%�bw�w�iȖ%�by�����ҝ)ҝ?O{~K6�b��ZԻND�,K�u�nӑ,K�G�k��ND�,K�u�ݧ"X�%��u�e�r%�bX���v�R]k(]^���Z:�䓩�L��n��k�]4�Ur��N��4��i.�G{���D�,O��{v��bX�'�뽻ND�,K���˴�Kı=�~�m9�)ҝ/��}�c-��-2�t�t�,K�{�ͧ!�V(9"X���K��Kı>ϻ�6��bX�'�~��Ο��N��~϶��v��[sSiȖ%�bw�}�v��bX�'���ͧ"X�"�dL������Kı=����ND�,K�>�ݙM[���f���K��K�U�=Ͼ�m9ı,N���6��bX�'�w}�ND�,q�1`0�i����ݗiȖ%�b^�m;{�3%��f��n��ND�,K�}�ͧ"X�%��H(>��?M��,K�����]�"X�%��}�siȖ%�b}�ߦ^�h��Ƙ�&֕���������b���.͍�,0@vkiQ��p)�c�Z�Ο"X�%��u�ݧ"X�%��u�e�r%�bX�g{��"�%�bX�����å:S�:{���͍�T0.k���Kı;��N@�,K��{�ND�,K�}�ͧ"X�%��{�ͧ"~Qr�D�:~���	�5���un�kZ�iȖ%�bw��~�ND�,K�}�ͧ"X�%��{�ͧ"X�%��u�e�r%�bX�w��Զms����:|:S�:S���y��O�X�%��{�ͧ"X�%��u�e�r%�b���u�ݧ"X�%�|�zS6k�m���:|:S�:S��}���9ı,N���.ӑ,K����nӑ,K����nӑ,K��u�k�S�Mq�ۤ�2R&�����c[u(f�l�C{v<H��$`E�$!	�3�D�!	�˔a$3
�P�Ʉ��@1�&P�փ�bI�D�xR�,�BI��<y�g_<��}�-��-�%Uc�jBl�BB.����@!$�`A�HF#"�H1b������I3)k�Z��,��1H�ZrՒ,�ٰ�B����r�$����p-k�V�VV`Bws)�m����`Zm��"�D�-��c������<.�0�,�ݻ횝۵��<�(KnB\�ҁ���
в˵؞�����3:��.�{�k��n-ۣ��sI�'cs��m�h S]G�HM�̀�D7R=v.���=�U�yw;����m�4"K	aHqUn�f�GpP�bVǒs���.Ӟ T���|x�eW������xq�:��vv�k&�N4� �°n��yv�h5�+��`��$Z�˳�q٘��Es��9d�Y���pf�1km�� 2�$�j�j�	Mr ����t#m��SQ��,�����h�%��i��O���4;��Ŕf�t��ͥ��lq����6����=�L�`�r�q��f�h�.�e��/<�V��zS��J��mT�٣cSB�����GZc�R`季-��&G�N�Y�!<����fL;<�js+��Rp�n��j��s�� ��m�4��I�8
8W�1m��h6m8�d6��Z�Wfn;�)5�F� j[-T�R�Tۖ����ViӍ��pT��rn��ev�V�ˀ��ۑۜ�q��'���q�e&�[���r[񋅉���.-���P�iU�Y�j�\is(e)Tj�f̀oY�gM��W9��\��bH�j��¬fj	0��
����ź4�k����X\�@m�hv\*Y3v�+�J�dշ:8���Wmȯdݓ$[k�VѤ��n�� s�XV+��a�I�pŝF�!ud����gF��[��C�4.;=M���Ǯ����m��[�Ŕc�H��a��tܵ;cgIσG-�@s
آ���*nΌk{=���sd�1ۨC�h�Ѧ��R�<�X�h�XD-��*GWd��#�����콁.�(�y���F�Sv��t�r�X�n
(���ʜ܎d�x5�8�v潉��Q��xή�kE��ժv� MF�Gl��U�;rp�lW7:y3�(!�z��]r�K�묱�1vfEw�45,/@͹�֋����E��|h�>
�� " ><�� ���4S�6����k6���Ť[*���̈3vٰ�F�B���ŭ :\�� ��жe�X�h�0���6:���a5� v�3�Nśe����X�8� &iHx0��SW]>bs���6B�5�b�C0
+�nnv�=�z�����RNՎ�"�b;y�f� ���y�jf�YK���i��(����gpsbF�R�(�Y�c2��N'wj��0�����c��)�Y�lq�u�뚵�C���Q3�t�������&�mMM�"X�%����e�r%�bX�w]��r%�bX��]��~X��L�bX����ӑ,K�����f�j��Rk5f��]�"X�%��u�ݧ"X�%�ߵ�ݧ"X�%��{�ͧ"X�%�ߵޗiȟ�H&DȖ%�}i�}u�ٸ�.�O���5�O��߻iȖ%�b}��iȖ%�bw�w��r%�bX�w]��r%�bX�{���߀�j�-�å:Rt�O���ͧ"X�%�ߵޗiȖ%�b}�w�iȖ%�bw�w�iȖ%�bw�~��-�e��o�>)ҝ)�ߵޗiȖ%�b{�w�iȖ%�bw�w�iȖ%�b}��۴�Kı>��(_��rWn�0��M��%x2;����=e�X5]�m��e�t���R���F�Y5�.ӑ,K��}��ӑ,K����nӑ,K����n��O"dK���~�]�"X�%������̥�՚�LfkWiȖ%�bw�}۴�0�T��7ı3��nӑ,K����K��Kı;�w�iȖ%�c/���,��3�m��y��ҝ)Ҝw��nӑ,K���K��K �,N�{��r%�bX����m9ı)��>������QGf���ҝ)����K��Kı;��siȖ%�b{߷ٴ�Kű;�w�iȖ%��O�{}�2�ʤ�hܗΟ��O�W������
�}3� ���X���m��]�ܤ\Л�.�H����m��L.�ٷm�#8\�c%�d ��������Ir,{{�������׀zy%E��c��i�V�K�g���H���/{׀M��?|��DL�6�E��m��=�<,)%�M�	�XA"��8��9�s�N�ŀmM�*�wM�LN�ذ?W����׀~����$���s��;�?|�t�4:l��n�	��`��~��۞��˖��hn�+m�4�`�oL��vEl�J\OBBv�PS�b�q-j�ۥWB����I�v�%Ȱ	��XRK�z_��ժ_���T�46;��	��Y�#������,K�`U�F[`����hjذ���M�������s���J:-շWi���~���^��X�~��&߿K�:��FFw�1����:I@���`F�:$70�,k���:D��+"�X�,$(��-��CQ-�B!���
B���C#�Q��]�~-׿�f䟽���%˰���m`\� �{�E$�-�������M|
�V	�q�a
����A�4��.e&)g�����į]du��+��6� �Ix[%�\� ڒ,��X�ۢ�WclXRK�U$yOz�z��M���9#��WM[��e��w�E�^%Ȱ�ԗ��԰/{׀�R����ۺt����%ȰMq�)%�z������T��N펛�X&�������f�}�}w$���`�M߲�����h2�B���B�&u�1�WG!Yeu.m3�D���h2��jc�c	��]J;#xY��˭�Y��$(���j\��MV�1*\Fhkk�zɶ��s����j璞]�A���j�)yy@e퐸����d
�:s;u�&��s/lR����fl-,b2��3�eL���q��H�RaŶX�jR� �L8�e>ww��{zo��,Er��;d���i���;l��ųEjAi�b�LƔ]r�p�ʀ�;��}�۫o��	.Eﾮ ��X�%��.�V�i�6��K�"�^ɮ5�K��f�"��߻-)?d�͚�jf]7x�����95ư�|�$�ۑ`��wawWuiv��JwrZ�=���6�XRK�6�&U�e�m�M+�M��$��G�.��z�	�rέ��p��[��4��L���8*�9�x�قW��Nq(�EҏN�܀�cuZ��XeȰ���ou�^���޿y`}�R�.�;)�V��xRK�R�������Uٷ�Z�9.E��<�U_~���������ƛ�x���X�"����(),�c����hwm,�������`����"�^��%�5lv6���]��� M������޾���$�45����^��c��u��0;����^4/��=l�Y��J���7:��U����vk�`\��\@O{� ݢT�#���ڮ�������;�=�{����"�^~��5ǝ]Z�&�՗e���_��l��P��EU(�$H�!�F��)
Q�$�
����$!BD 2���H�R�h�#K�U_eVW�R<��x��%�rG)���Ll���Iz{� ���x�r��'u���o����4���F�;f�K�`���I�K�Is� �2��z�j,I�1�����,�\�]�n9s.�G-�vӏYc{b:,X�F2���Mڶ� ��`��`c�꯾����uA{�[��[�ݴ;���{68`�"�&�g��_]�⼽�6�e��Wli��~���0Kذ��X�\0��C��ӵWH�m�Ի�<��~K ���UT��$��@ �	dW��T}�J�'/ ݢ&O���V�I��0��X�����~:�~��Mp��yo��EZ;2�8�c�+l[*��gi
��f& ���*y��m��y�uv�X�\0d� ��}\A=��=��CUt�i��� 7dx&�`��X�\3�W߾����]"��&�
�v����f����V�x�[j�:��M1�v��Է�<�6?���?}U��.�g��޻V؁���m]� �����������I����ܓ߽�f�'�(���� B"1��S�E� �D	�ȩ"����/�6hO^�v�)�)�$�՛�T:`n�@��Ek���f�9̉{-G�� �,xxT��7Tq�X�:������l�n�p'�.�]č����c�Ok�$�*��@u���`+nZ�Q���ϱh��`��NLmqS�ݮ�O�!F�a�.�`��4��l&�Bj3iLR#,A�Ќ���i���[]Kp�B����)��F�A���RXeqn̹�$��.
���둍M����r�w�7��%�1v��qe&��>F���b�"�Ca,��E:��}<�Mp�6l���q۞XQN�ڤU�,V��95�?Wԑ�Oe`ny`k�~��#v����h��t2�f�Oe`�ذ	/b�'u� �6�զ�����`��`^ŀN��{�ܬz?P�]5i��h��X�Ȱ	ݙXݙX��X�� �)1`�i] ��%�Q�yC��u
.u��ݣ:���s�ăޞOx6��`�]I6��{+ ��+ ��� $�����J41;v���0	6ed9@����&�N�ɝ��w$�w��8g꯾H��O+V�-[*ݻj��<�M� ��2��c��v�+Li��lx$p�$�U)��7|�J�u��ȺE��x$p�=UU_U{�<p	.y`���x��:�?[��\͡���J�s�Y��,�����n�t��.���hF+t6��!�XX�]'t1�g ���n�ŀI��{����������=f���b�kl�7ob�$��8`k�$pk�n�wV�-��N܋ �x�y~8�l�T�%!hl�Pk`ЅYH�ÙM�Ѡ]9�Q2,"2�-LW0�5q@3i2R�)h�B�BK�Gsar�˳3���e0 ݒ��5`�3�r�	r�.h���� ��.3T	%m��!"ҖR�������(kY���fa��u��1"HXSZ	m d�W#@���a�R��4�X@��[*(lع�)n��Y��a)�!����L�oT�J�$	�0�HBA�$i��a��.��g��<T�2ҡ1Y�)_o�YB̺�t0�4�(�OAJ�H�a$�!"�b#O�@�ှ��@�x�"���(�{�kٹ'�g�]�'�}�d��n�Һ.��0=U�.��� ����{�\0�J�S����0��n�ŀl��8`%#Ҝ��K�5M*'W���3r�h���yOfg�8�okb� �1���%��Wl�\����0���R;b�)���6�M�?W�W����ޏ��{��*iEi�J��m��8`5� ݽ� 6lx{F�jP�t��T1�f�\0'��]�'�{�� } �0b� B��[����������������X��X�c�9.E�lٕ�z~<�����Ҳ��Gh�K�u(����b�35,��5[H�]p�XA�v��{Ȣ�\ ��x%Ȱ�2��ذ��v�J��i�t�ـr\� ٳ+ ݽ� �\3�U}�G}
g��T;i5M��X�=��n�ŀ6<��XE���)!��hm����R��, ����r,R�3� x����wn��'li����r,���nI���rO�iAO`
"B#������,��E4�Ad$ �YP0����cPVAG>o.Xh˔%%�˨@5���ҁ-ym+ce#1ijFS����s�V7g�d��B%�g��HU����8:���Nm��vGF��˘����#�94�I@Բ�H�:x��-�qk� �ƹ�Фg������e�us�Q���W���q�.�f�L�^P�5�2f�bY�t)����j7 T�vUb ��o���;�yKE��&��iC6��ѳ4�P�l1164]m#�ERfI��d��<�m���`�p�5n��}_q=<�Ѕ5�4�i����6k��v^ odx%ȰF�:�t����e�m���x�c��%�_��	��`c�/�6�Wt�V�� ٱ��"�6k��v^ w����E۶�ժj��9.E�I���x�������N+tF\2����WR6�Қ�\�d�Y�&���lG���5 ���Jڳa6:j�e����jݗ�l�WN��P��{���}���YK*�d2�ܓ��f�p�Z�)"F�P�L�,@ ��O~澛�yۑ`$��V�i�ҫ���m��8`�"�6I��jݗ�otV��m�Aҍʞ�ӯ���� ���`�e��� �CJj&��[j�.��L������'���\<�����~��u�#�Xd�,e�5Ф�B�[���/l�7��F91S��+4f2Seح���� ղ^�{�&V68�S��wB)�k 7dx%�Xd�X��, �wg�զ�v間Y�nIϳ߮����7,�E���ذd� �%4:�7N�[k ݓ+ ��ŀ�<R���:�g��銓b�`���7��`�������|���nɕ�{����3`v��(F�K�f�({s�ܽ�d;C���tc�hfD��E"�M\������r^ŀM�+ �ݗ�w�$�ϭ;bn��m�%�X�e`�ذ	#�z�&��mZUv�ul���{���7��`#��{ J�#�N����;.�n���X{&Vɟ}w'�ޘa	�dXF4XIIe��1I0�`S)	��d%��l!)XHY-%*C�*99��_�_0m՗at��k �c��{����7��`�ﾪ���4{��4.��[h�OgP������k���b�Np�"ι�D����6߻���w�2�]�xd����T�[��m�m`�̬V��l���,߾H�6R���ؕ�Wt��ݗ�qwS6�� �ٕ��H���]$텷x�x%�X�fV��/ ��	YV��b.�����`ݙX��Xd�*�����!�bYĊli����~֊�P/ ]Q۞,XsAg�ݗ	��W	���׆�t�����ΈR�dT׵��+���Tvb��]���Y��+�q�r[]����6��=��;8A�qx��籣S�ǃ8*���,b��b`L�ۇ��J�c�v5Z^���#1V[���ɣ
$�1�J���f��S��}f�xcr�N3g],Ф6�ن��t�&�m4� ST����!�d�qo.�g�+�k�bh9��X����]���e<���9�������^;0kkc�MX+O�Eح�7\0-�x�p�9�2�l�V�tպmZ.�4ـj���'c�ɳ+ �� �wg�զ���Av��_}�/l�w���'u� �nE�rh�M�����{&V;�{r,v�, �ҭ��7��!6 �%[s���̼��X'us��k��i��阅�*��ƦB�����ɕ�N܋ �d��4R+i�j�u���jnI��}�~�Z	�J-�7fV7\0�D����ڶ�m�� ���Xz����=��s�h˖���m�[����X�p�&���'c� mJ��P$���n�	��w�� ���s�N����ͱ̤4�����l��ֶ���h�A�tn,��̋�\��s�M�h�T6�v�,v8`�e`u� 9]��i7n������� �+ �����$rkU���7t퍳 �+ ��3~���@�R�:B����`!���i�(�U��w�ܓ�{����5l�۫��i��u����$�S޼��XvL�*Ԥ�C�iҤ��ݳ �%Ȱ�2��p�'@ڀ]YX�C@�]ҠI҃�FR�5�sV�6���QbmE�u�8׭+]�-�l�9.E�Nɕ�n�;�;F��n��V�j�wm`veg�����$~0O8`�"�}��$��ί��%B�n�	���9.E�rk��&V�&QV6�tݴ:T�f vH�Mp�7d��TϪ��蠒FB��$��b�>��|�M���B��
��RM��\0�X�\0vG�M+\�튮�[�����8�c�;<.��DVc�"��ٟ�kg�i�v�s�(]T�G"��>��O ��p��X���,���I��֝ l.۬{��G�r^ŀlٕ�EZ��ht���J���c�9/b�7�e`��wtIQ>�;��m[w�r\� ��+ ��.���F]Ɨ֭�ղ���'ve`��N�ŀr\� T��F�+���k1���i O9���p��3�MJK�ᴗZ��K�0"� B"�J��lHI$g����� �)	b�i]�!!8� B&a.��!L6�XR�����qf��%�.���[;wq�ș�|	P�Rd�oy����.���>���嬮Q��˾|�1[�>����|�$瑒�cʡX��>~�5�f���!�� H՗�|8�xm�R�A��d�XF�3 @�
+�x�)�$!�d`I	'���y�J�yIsWn��nf�֩O 1��l ^Z1�Ғ*Ip�e`@�d �cP���,���##75X!�"b���$�w�E�C�%\o����Cq�7p�M�]�0�P�)�s�%��a�i�#ă	6�>@>>O0׃M�7u��_����M�f�jg0���>��N02,
�+Ayͩ��S��I!0!x���CG����b�bA�)*� B$a��$� ��hSa�,&�7&��B1|�E��n�.���"�϶C��a� 0��9�p����HOНӯn��˿�����mQS�i �B1y�C��*B.�D��(�c6Ktt�)[�=ɺ�P��t*n��D��Y̋�<���X]�aō 1M�R�Z�k�¯<�^)�x���ǋӦB���y9�՜`���]�7K;���T:�&����88�R��q��̓*:Y[[�6��s`���7�yK��j��V��vݝNyà�m�]�qI���fU�hl�W;�i�q��b����6y]x�:���9���gx����X���� \f�bKhH�n��h.WH�hҤPf���j��q�ж�\���*��(v���j7k=t��a��n�p�0�m�힁y6|��Am+]��3Ult�O��g��U��.U�9��$�ϋ�m>'l\p�6wm�K�z��	DŢ��ӎ���!ˮ���5�S�Whp���D�Ak��sfڇ��|�+T�m
YTCPc�L�M
��OV;�ŝ1��v�s���]P.�ϴ
��ݓ*�En��x�v9��q)��9V��te��H(�V���pl����6��j���O4�q��`�E�r"m�7c$'�q�M�=�]�l�+lN�!'u�UJ�Ԝ�K8�^7@�j,Ŗn{@�v,V��NTd��VX�m���� �izmx��<�DN��:{iym]��ˬ婪лRr;��3ѻK;��"�N�=�'b��g" �>���9t�c�K�R�5й0��l93���n�+��H�Z�A:�jĀt�+YpQ2�S�����;���B�g�u�X8.]i�X�A�FeN��
R��sa�J�A.{745�[/>�z���ӎ�bNt��l�l�-�F�l��g`y)���f��F�G�t�aJI���W�4nں�q�5=���˹��=nL�8�pP�E��5��&q�G;	�r�nˈ��lS��wXk9|/m��G���PkiH�f��/W�:�<�Ʌծ����7/Q�.���(�m�A���V��ќ*�:�Anw�t�����
)Oh���� ~4�	��p#"�B�At)��� x��z>�^F{ h�R\�-i��Ȍh�r@s�#r�i��k^�ܑ��]���`<� 3�$h���`�ւ��ʓAtE���:�e�j��,ΖB��m2R�q���F��ROe-���3��Wt��mV��9yE1P�W6Hul�7�k�p\��@u�h]Z�!c��8f�x�^�j#�E��p>ݶ�"1��bⶑ��%5�Z���w�$�%����1X�1�v�=!D&�\ٻ���r�nY��UŰuQ�Ze�5f�`��J�fum��yp	�ذK�~����=��X���>�ڻm7eҡ�`u� �$�X�`7T���Uաݳ ��2��`���rF�0�N�ۺv�ـl�+ �� n��.G�`��A]4�M�Cav�`�p�=U��|���vI��{ｶ����j3���4u�8|����M�[ dۭ���P�kqh�t��2���v� I�<��,�L�WI�lT{��i'ljۼ��Y���W�v�������ܙ��su� �r,��F+���lm[.�I2��p�$�%ȰjB:�-�ڦ�j�n�-��`G��X�e`�`i�v�n˥Cl�$�%Ȱ	$��7u� ���wr���ڧ�n�&��jx/-T�xw.����\�6��"y���?�T��M1\��o|��շ�I��n뇫ﾮ �����5^av�`���`$��7u� 7�<�8`��K�N�)�T�E�u�n��nI=�ﵹ߼�B! �i�W�}_||(��`�L�*5Hˡջ�B�cM�W�WԔ�y���� �ٕ�n�ŀs��D���۠Bm���X�2��ذ�c�5-��rٱV٦Z�H�V	��
ٴl��5�X�\qXg�P�Ƿg8��+6�>�ٳ+ ݽ� 7��r, ��#��I�LIZ�[�v�,���W�$g��_��M�X���ئ���6��[k 7v<v�X{�K����K�X��$���*uj���	��s߾ٹ'��]�Ê��B�O=��܆��ڱ�6ـsd��&�ŀ�;0��X��+����O��yR���W [ԌD�Pղ�!�C[�1��.ڳ1%q�π{�����c�'c�ɳ+ �F�)�'e'�Wl�l��ǟ�#������'u�=�w��*=��C�TI��{ny`��N�ŀݏ �ѣ��wc�ն���9��Eݗ��ǁ꯾^�<�ka�M�;bajՉ� ��/ 7�;{ɮ�V��m�r�ú�[�f(�k�w��!ڝ7;eF�$8��Д�6�!�[�3���X�,2����R[�˲��L�]�vRt���Z�8Sc%�	�&��D��b��e�m�W�ɷGn�ڑ;
�lnS�g0��h��@����j@�T�d�F�5�v%���S��00;u],i{�'q[	ko<�.%���f�[ulӠr���c�-���s͸8�N��,݃�������b۶��9.��N٩��G!�-�Dn�40��m��|�m�� ��v�, �uO�M]��ӫT���'u�5#�3+ �� �v<�)���6Վ����+ �� ���	�p�;�ԗv�N��N˶� �� ���	�p�9$��5Q�JwI�N�J�����	�p�96e`ob�?U}_}_lq
��i���2�Z՝
ر�k������7gl-Im9p�h�:F�+
��kf�{���rl��'ob����ǀs�jC���sq��um���RI���bA`AXD�H�$!��_�_]J��V%ݗ��<v�, �H���cN��b�X]�x���	�ذn̬v)�t��v�t�7x���	�p�96e`��`;�|��;t�Wm��"�96e`ob�ݏ 6�Ge�;tZcV*���lV1�ƈ��&��KRJ��1X�fa
�3,�6��j����L�n�`wc�'c��.��n�c��.۬n�`�c�'c�ɳ+ �l�����7l��ǀN��� l��B�" �a	
��)@/���nI������Q2ݰL�T�$��95� �ٕ�ou� 7��wIT�];��V���+ [��p����,�{B_n�GIdX��7ZS�/9���nV윁���6\�u9՗�щU��`�ذ����,��+ �Ԙ%C���n�v��ݗ�I�;&V�ތ9տ!����ۼ�{�ɕ�ou� ����9��p�v5bwcl���ɕ�ou� ������W�UU}����{�.��n�`ۻwv+n��`]�x%�X&̬�/Oa~)Ym&ݤ�Fm���Y�Q`��S:��-ԝ�\��C7��V�i41�M��pl��9/b�96ez��� �s� �*�vZ���1&��{ɳ+ ��ŀݏ 憻B���ݰV���fV��� 7��{ޒ^|ۻ[�wjҷX��,Wv^�{�ɕ�wjL���M�7Jݻ�;/b�9/b�7�e`��M#�H�EKF�.+ܴ�����c5�j������.1��cOM=j� �Ǳ���!��X��<�Ht竳�//Og��yk��� q����{ 23r���T.�=83��Gi�q��)���-�V�R���g�N�M]�����4���K�y���7F..Q��$�疛�^�N5h���nC�����4�Ӹ�;:�e3����ϝ��av�ċa�f�j��K�(��<p��<`�	K��#�V�"���6:����_���2��p���}\A��������XՉݍ��X�X�`RK�9.E��#�]{�lWM�t���X��`RK��%�G� ����"�v�v�մ�+v��T��Mp�7d��7��sM;Q��(Wn�Mp�6l��7��j�/ �
�DWXy3aŭHj�-�\l�1�` 0��K�B�k��0rb���Ae��p�-��͙X�\0Se���`�ٟ���.fe��rO|�_M�E�!"�H#f*�I�엀oob�;6eg�����`촄؋t�l�"���9/b�96e`���`}v�M�t��x���|��w�~0�p�5we�]�\)����e��Mp�7ob�5we�^��ëoߡ�!97�.Eє��Ʈ���v�5��6�,��v��nݱHvi.y�1���I�N��n��$��j���9.E�rk��GwI��m�j��5we��"�95� ݽ� �M;��ЄZI��9#��0t��M�R6���>����!�<%4���t`D"@�E0� F�I���Y�i݁9RQ�B���dp���0!BȗD$�0�r�vkSZ�,X��t�ڤ6���I!J&%�!���$$Yhn�!m$!�y
O#��835n��s��`�! ��O8I0&ap ��!	 @�V�����[*%ZA��*�"@! D��&��&A��V�+��P,0n�C�8am#
JXXTA6n�XM�Bii!�]�ڭń1���4�
�  ���!x�70�a\i���	 ���r�m��  ���� h��Q��~�xDW�T~QA 6����.US~y��w$���ٹ'<�P�J�)uvƛ0H�ou� ջ/ ����S*�*�U�Wj�0�`�e���`�� ����:��p�Z7��q�l�RcA��n�#v�W�BQL)vꍺ���4ـjݗ�r^ŀrGW�}�c�	����V�Eۼ��,�W�$w�~0	.y`�ǀqv}p�즪�V6�m`�� ݽ� 7v<��X�u;i��V۴7l�7����O=��nIϳ߮���`�,�# V+'N��l�?_���>�{�?7[�l���< ��x��<�g��{����!�5n�bA6�����mZJ��'#cI����Ȉ�[���2�3\Ū���X68`��ݏ 憡�N��0lp�W�|��� l�x�g����7jz�-4[e6���f�� wv<=_}I{c�vy��;+fR����'j�6`wc�'u� ��w\0�[�*�V�.��'u� ��n�`w~��">0J&L���ٓP�5�c�s���pˊ{�E]��jK��,2l"Ҋ(�\2�ٲ�D��Pn-"�#0�FxCT\��<qƭm��;5�G����F�b�n���yyL��/(w�7;��zh��`6-��
��σ�^Wm�%z�b�SuE�1���|�\�2��F��,���]��=R��y�*n*nW�ѱy�����u���v�1��g�w�%��r!(<f��vy�����k���n]V�O��M��:��2��X�;j���4�~0�p�5n��9.E�IWm�t�m��`���K�`��D�;��Ս�m�j��5we��"�95� ��ޕ�|��7e��M�����9�w�~0�`�e���4B��]��k ��\0[��Kذ	4�yI�i&충���V�뀱P<m�H]�kl
�紨��Q�V�)]����v鉵wvـou� �ݗ�r^�ﾪ��?ʞ�_?��C�z&��7$���ٿ@H�Q%��gܸ{0�`wbK�*�V���x%�X68`�p�:�e�[>�:c�mX�-��諭����M��ջ/ 佋 ���m	��6�-�0�`]�x%�X;<��o���[R���Y��u%&��ܲ�d����3�L�(.�ֱ�mTMA�Y�n��`]�x&�`�p�7��oJԇ)�WcuvZC�x&�g�����#��� ���v^{��#�%!�Š`ӫ��ـvy��7��zFHD�	B2��0�@�a�$"�`�P����;��`�l��۫n݃m��l��W�R�3��O^ɮ68`�ٔ�;bT�[��w�un��9#�͎��xA%+������Ф�sv:����u&F t�B5m�6���i��P��"��6w�|���x68`�e�]�x��)�c�6[�e��Mp�UW�|���-�� ��~�|��wZ{�ў�Z��\.f��Wv^�r,�\0�[�]���M�C�x�K���;������}7$�"��1�(`!)3eW@��u�ٹ'<���*��n���ۼ��X&�`�e����MI-���0aJ۷]����C�:!x�4Z����E;���5�E��J��i:WV�0Mp�5n��5we��"�7���)��m[�ݻVـjݗ�ݏ �ɮv��|��CJ��� ��x%Ȱ��UUIw���"�׀�(E;47e���r\� �c��v^���o߿�|���^X�̳*+|�����������9.E�J����xkl���9m���FkYWP�V:!������hja�5IJ����k̼4�xARq�X�v{v��r��ս=�|���i��m
a���r�&�<v����خ���3f�+aԂ�S�����SY��#�����їBŰ�i������ua���m���Ŕ&Ҥ΍r�huc��ن��Y������g�ݶ���lH�6΁p�W0�޲w|�;��ì��A�}�F���v�m�6�]�,nvd�-��uͲ1m	�A�W4Cg����/{��{���"�W�}_}���� }8s�C-�4U���m��x���@=��,�~��&�ŀoJԇW�ƾ�wI�x�Ȱv�X�ذ���t6�4O��m�J�k �nE�E�/ ;ݏ �{����5m�v�[���0	ۑ`{��ob�9���m��	��#����[jhVmWjx��D�Ԁh��z��2��(��A��Mb�%CJ��X��x�ذv8`�"��J)�4�l����	��d���T��f�8`�Ȱ.���U�������`�[t���wc�N܋ ����"���7`�;m5t�m�;f;�v^v^���wfx�""��N۵e�Mۤ�v^v^��6�,�U_w\B�n8�c>:����������#q&f�E�#\:�8 �h�I6ԉR�4"4�[�^��ŀM����[��M�ݍڤ��w�s��W{��qM��E�/ ����5m�ݻNڻl�'��]�9|�����H#@ E"d�M\���ܓ�=��rO>�ˤ66��˷H���ݗ�E�/ �u��_W�|�����*C��]�J�
��vK�=_W��<���,��� 6���cn�-��V�ڴ\F��F#e�u���݆��s]���0�OV�+uzt�n�vۼ��� �{��ŀE�/ �)�զ��;V����	��`��X]��v�,�W�}_$DE+¦�N覚����;�<��%���X�ذo�*r��Һ�v�[X����z���,Kذ?}�Ur���"LQ{�ڎ�_w[�ܓߤ�-�m0�e'm�X;���`��XSe��J�j�'V��
c�����C�g�m��r�I�H��T����٬�:�x[����ؓ���0	/b�9�ذ������~��l��`���]lb��N�X�XV�)��lp�$�� ;6RE5n���Wav� �l��0��%�\��5I��9�!V�t��I�M�n�lp�&�ŀun��"엀M��:�i;e+-���	��`]�x]��v8`���N�Kp��|d>4�g2�y>0���:�/�(U�HI����I�D�� E�����@`�$",
�Ba		@v�L�Ea$a	��e���,�).�5��oc�(KiIH����4kM��!��v�X�9q�sZM�&��@�AL�c!�0�!Ĝ���XBl��o{�D�`�"	�D�6B��2H�BB0�@�	��_@�0���I!"�%-�34�����|�y�߻������D�|�,X��FY!XP��b�)0 JjF"��"@�Q! �$$2)XB$���!�۰�-m���H6���ͳz�6JR�]fa,�(�a#Bm7"�a		��oa���3]]��nQ�9 �0+D�	�����T�6V
B �Ga)HB2F��!��	F1�I)d����1����Y4J�+
ĉ,#M�h�
� W��O����� �m���;���(n$�F�ݧgh�̝bE���^��5��9���Лv�Y1���yE�퍝 &���:�JKZ0-�:�t,!37WKBP�rm����;J���ã��}P+����9:��릦r��n1�<V��8�z�8������x�j�-=��`�a�t�ْ�)^LJZz^���;M<Z�yz��J��G%;=t@\X6�[)��[`���^�N}nL��q#ҝ�=g�z�S�,������n[m�
����ѭ�Jv��z�����ɍ�B�:�R����nڙ���F����;Tn۵Ȼ"k۬�����.��8�Έ��<h�=��5��L:.�Τ������+&������ں�W\�ux��1jꀋ�8&A����H���<5�PFc E�-�u#e`K���IG�1f=ttp�cX��t��p��;y�~��`$��`V�ep��-Z�L�.�I�IYٞ[)nh�=T�7q3::-�6�;p�ۊ�]-�ո<g�Ѳ�t�l�gX�R�E�e�`�4U]�J�o"S�Dʹ̘�7�%�P�X玺��'3��`���
g-�C�L��<��!D�6��KBe�Y{5�x�[k�i�3R����8wnc.�ɞ�^y ��V�ӳS�ma�6|��M1�YI���[E�)B����v��b��a@z7��b����=�A�E���PqToGgrvM�J����q�gF��Iv\m�͂%a��lM5;M�YS )��geb��f���mK7��2���C��狃�8�Z����k6:i�+EP݌�g�����:���s��¼�!���y7h(��V���y���/6���R�Շ3`�o/�CjóXuIy�FX�0����W�70���R�[;E%�n�(N�7!�.<a{u�D���L�ոM�b�m:x�Ƴӵ�a�3��6�/U���kl&���AK�����ϓ�Vָ�4+�b�L12���u՘d�dɫ��I�> <���l<j"��@�M���1�<Uq�@ׂ�z�y�����z�;9M��-�l�v�_WVZ{Q��T5�֋h�Ǻ�$�n�D�k�P�!tk��3��ʠ�ֈqj�F/+���T��L+vL�r׋^�MB�Onb�����X�,����Bз@�n�e���c��v�.9*7dj�����.�g�����8��e4\�S�8����[�j�ٱ�bL��.��1�zK:tX���hU��JP���k�5"��LXZ�Л摆��.��[�0��{���M��h��C�E�����x]��v8`ob�9���7C�u`���vK�9��M�� �����UU~�������ۺt[E'v��g���&�ŀuwe�vK�7���[��uhv��f6�,�v^d�|�=�0�W�������N�X�XV�.�x68`ob�9-j��Z-����+��t�UKq�X�I����ƍ�$�\e�g�فbf4b]6�����sum���M�� �ݗ�snB�)�!ն]k5�f���}7�D����!�]�4z��Z��5�nI�����'�Ϲ��$��_��g��$���ٽ[~�~0��x]��lp�5jZA}ao��؝���nO^��������eA4��;���7x]��mȰ	��un��6�{l9LK��m���+P����K���V��t��J���h(U����7�#s6���r,n�`[���UUq��׀n���|��n����vـM���W�}UT��O^����ឯ�7}^ʺ��vZv��6`���n��*<(� H*2�����}�}��?7�� Wd��j�1��uwn��e���N܋ �ݗ�qM�4S��	�Lv��9�� �T����'��{ nҭ��4��nf��ὄKv�T�P�)pJ\e����v�C�`ϰ�Y��$4�7���?OP;��{͎TKH/�-�S��n������`ۑ`�%��Dҍ��Cn�t�o 콋 �܋U%�׀'��5	������[m�X���c���׀ݚܛT��<_���}�ܓ�o�m�V�4ݦ�m�d���<�����Ix�4�M��e��.��-�R�Z98�-�qI�˨��W]N�l�v&:��� n�x[��)%�vK�
� /�c��`�o �v^~��ꪤ��{׀yo�x����H;�����շxT�� ��^����6O<�O^$GN�n��e�ۼ.�x[%�n��"�/ �Դ���'�ӻ�n������rz�T�� ��^ϫ��dM,K�ؔfc�R��R# ��Tn6�)$c�&XM[��ԋ�BK;cBMl�]�-a��-�j@��%B����;f!ɫ@rrݜa�n0=�Ұ�*��L�ķE��Zn�^+��۾�I��+�Vp	�-ź���d���Tհ�:; ��K�Q�̽�Ε ���t�r���43%bPr�5.Ѯ�`�*���'j,�H��HMePe7�'t�I�w^�7`����>�#5��M��;[�s`��G*מ�s��Qam�pQ�p��t\`^�� �܋ ��^ wv<�jI
�#�n�ۼ�3���}������׀����e�����#v��e�Wv�v��0-�� ;���0쩖	+O�v&:��� wv<-�x$p��}U�/^�׀=��uo�ۻv]��Eݗ�rG.� ���	�I�ݵt]�쫻C���-!˓c�۲�,�9���l/�}�oki� vX4c��b�i�h��w�;<�`we�[�����	 ���vշlAv� ��/����~�F��x]�x�x�KH/��u`���ۼ��/ ��/���R]����׀oMN�F�+��4;w�Eݗ�s�� ��/ ����9��4��Q0�wi��9��{���׳�| �<����	4���:��{I٣*ك��ә�\�M�8�ͳ\����l-Ƿ��4�Qk`we^ wv<.�}\A��� �A��H�c.�c�n�^ wv<.��8`��� V�|�o�ۻw35��>�=��I���f�6�IU)�p1"�"Ć(|a@>���O��;#�Ihbv��6�n�X��	�r� ���<��y`��W�պM�m[H��'u�0wc�'ob�8���sh�.�����nm���+лM#�̳.Еn��	5�y1Av�ьj�ZL��M�f^���}��	�p�8���N�`��)N�X]1���	�ឤ��=x���x���i�v�wb�S�;i� �/ ��U��c�&������.�cwbi���_U|�{�U���}��nO<��@��*F"X ӧ��N������(���Um۫��ǀM���^d��o�����7��R4�����563-��r�a,����$�:0b�[w:��m�˶�	�p�8���E�*�wc�M�.���t6�6�;{��8���	����H��:���tݷm!�k �����/ ����� թin�wV�ڴ�n� ����'u� �ob��W�T�{=W�l"wIy�]���4&� ����vU�]�xk>�P}�}u5KU���mK��,Q�hʈK�[��qrQ':��&�5MD@P�ږ�#����H�'n:�=fvN���v�獜cԮ-��d+��a��0P����OVf9�b�)�����J-���Z�����@X2�n����F�h�Yn�d^�܅ǁ�n
"�S�Y£�n��";���킲y�g��F�:�8l/-��vM�ӧC��I�����Y=�u�e�e��y��x �MZ���O��[sӧ�1tٗ��Էk^�W
� ��{�`we^�ݗ�N��֨e!ZN��+v'm`we^��/ �����Z�/�;�[)]۫�:�%���w�"�&�`wv���Ֆ�t����� �nE�M�(�:�%��H-�T;E��0��,n�F��/ ���ԧp`�H~ѷN��c�s�u�<�snv�{�3-�]r�T#5A�K�\ݼ{z09����i-��T��\��4M�9|���E
�m:AZ$�����rO��~��}����mjwJթM+-+v���k���ŀI{)`]��t6��E�S�'m6`��XSe^�ݗ�I�{Z����v��M��E6U�]�x��s��`6�iq;�I�4�غ��%TjI���G������hy�ٗ&��̠pR3T�fn���{/ �\0v�,)�� +�`/�-��ۺ��x��s��`M�xv^ N�tˤ�C�[m� �o߮�_}���`�i�p�xis1��ע3��;"ը]Y ����� �b�# �����V-H���55���&��kB�i��D��!��1~����4��uO�H�,`0Bl���p�3e�frk�h��n!"V�C�珞�o[�g�O-�$(KL�˓2�5��fM�,h縩��&��Y @�)�2��G.��>]k���ӽ����73�0d#"�!�d�cJK	tI��S��zз���c�'�᯶�2�d@�BB! �BU$	��Z�6K����5���[��-H�H�BB$����0��>!��3�	w�����v�a7��z�����uc��h��R�F�.��Ȟ[����8k1-e4�L`H� %��f���Y�kM��^S1����'�$�dP B0@ �!�4�BH�ٽo�-H�!�4>���@��`@�"���+�������x���A�����;5�:T�S�&z⩈%c F@da$�� �D��>UC�W��Q 8��9s�rN}����}� �9p�9TS�o}��[{<�v8`~����n��E���utĬe�&��.�x�p�;�ذ�e^ٮ�WP�N�"�U;����M��.
T+[��{<�u�]�#��!���^5:-"ݡ7x�p�;�ذ�e_��� ��z��JwIk�YO��m�{{��8�%���=�$n���RH�WN­:M��zG�0.�x��`��X���Г��w@�� �엀I{��Ł}J�������}"`:��4b��GowI�+�}��м(͖��g`^ŀw��`k�`]��}��}>�����%j�!��G�HD���F�5�d�,���٥54Z�rE��y�ą�m��s� �\� �������\A��?^��s�3�.pg*�E:���YF{���#�g� ����9�ذZ-Q+�t�J�-$�рqwe��� �ob�&�`���"&�J�ʷhM�;0v�,m쥀qwe��m;�����?���`�`#�`]�x�p�*�����ң�(��B#�f��s�rS��yd�kqQ�z���f�V�z^�����a�9�ѭcv�nH�]�smoi+l�,�m�s7$DM�lP��fLl�2�Ď��E�ݲ��b�̰��:�p�m�� ���2up�C��@3�9Ecf�\lz']O#�&����_[���it�Hl
ۊq��1��[I�������GZ9��P��\�̲��$��;�I0��{�i
b�����sL��d�q�1N�<�u���-p���
Y�f�զS�?{��p.�Mp�9�ذ�8_ʝ�&�ӫNۼ�d�Kذ��Xe�w����x�c�۷j�[���ͽ� �ٌ�8�K�	5JHc�&[�[�m`[%��1�V�x�ذ	6�����ݷw`ۼ�f3 ��/ �{�r, �!(��9����u�ѐ ��,�6��!�C,vPvj���['S�1����M�T�x�ذ�Ȱ͘�v}��?0q�%u� ����y�M;�ЈR+���� ^�S2�=��`Se���wIs�,'e���Ȱ��XT�x��X�E1T�]�i�v���;�:���'ob�7�"�;4p�N�T�&�.�n����	�ذ�Ȱ/����[~���No�>�1vK��V���\�bʛu�Y��F�s��[�`�<aj.Ͱ_�*vƆn�����ŀl��8�%�����m"۶���ŀl��8�%���`���\)�g.��[}��og��71��"�`�BA���Gj"�����}۹'�g���{}��+j���c��;m`]��	�ذ��,f��6�;�DӥeՉ�w�N�ŀz����<��~k ���?��'�)�ɚ P�
D��ŹŲ���{vD��۲𽉢l0��S���o�;-��uwe�5ư.�x��X{���I��ݻ����x�q���^v^��ŀvh�t�ZI�t��� �엀Eݗ�w��`5ư{�/��Amӱ�ۼ.���<�>��I����]�Ӆ!�# �B) � �!� ��@�{���䓝�t�jkZ��v���]����XWd�.��շ�?~9����FSKܴ	'[�!ȦbnGs��#4�պƎ4�P#2� ���ӧm��w�'��XWd�.�W�}��޼("���ݫ.ڱZv��:�%�we�]����Y��������i�QwVߏy����x�q���^��t�WH��wi��:�%�/c���^v^��Qg�6�j��;�x��� �엀Eݗ�uvK�'ݪ>�|W�F)�ZH��\2\��ٙ-�bK��YJ�A��CiAν�-��V6	53�.b�Ġ��f.+gk�R;�z�N�am�����>��ϐ3/���ü5�wX#�ႆ���g��	e���y[��MGT6aLf�H�a�
�2�$�c��4��$���#��8Iʽ�V�b<ݸ���"Jn�v����R�Rݳa4�HX�H��'j�D[,m�;�b�!�K���P=U<Q�<��V�fj�Z�Srr�^^^pa���n-ѓ`�F᱓q�E���\�	�Q��Ҧq��������n��:�%���� n�-:�Jۤ�ۼ-�xWd���;�:�%����ڦ���[w�uvK�;/c�?|���� ���v��$ݻ�6+w�v^�xd�m�XWv^բ*O�'em14�w�qvK�&�ŀuwe������S�n>�����4���5⣷oJ�l���z�D�j�بA�b�d��	\QwV�m�XWv^�{�]��hm&$�����;n��:����W+�W��H���lI$�!A�H0�_UUVq��.� �{��QeW`��ۼ�f3 �엀M�� ����6h�];)�`�v]ݶ`Se�ob�5vK�;6c0[�h��t���0�w�M�� ��/ 콎����	�&[�j�Wi�wk�㵪�y.8��(�ѫ�ܿk}/��]6����bA�-�����;�� �}��;/c��l�m�X���ݻ�6&� 콎����	��`�%�ۤV�,N�]�v+I�xT�x�M�@H`�U&{}�y�'>Ͼ�nI���4��n�6�n�	5� ��/ ��Se��m&$��O��u�j엀v\�����	$��?�;�����Km�12�Ij�.�t�z��X��Z�O6[YMv;	q�r��(�m
�v�w��;�:���$�+ ��/ �������v]�n�����${��V�׀r\��[�h��t���L��&ɕ�j엀r\�����Ceccn��[u�j���9.Gx�xUr�UW�)
V.6̡�`Е�H$�0��
��-i�Bp�*~�M?I?~y�y����ss�5�lM��r;�8���$�+ �ݗ��~�_�h�5elC@3�J���1lf����Ŏ�z�L�k��4f�j��V��ۼ�l�I2�]�~����[�į�˿�v��ۼl�Y꯾H�g� �y��6^Άҡ�Uu>��v���5we�����6^ɳ+ ��R�6���j�����������׀rl��5vK�9�8N��I�-�v��:���������גI�{��{�y�rO�
����E_��
����*��TU�@
��� U� �*��P��! *��`�AF
� �AR
�D`�D@��
�*P**T �@@��
�@���X*��X* �E��R
�X�`�D��B
�Q`�EV
�P �EX*V*�@ *F
�U��H*
�  �EH�R
�Q��`�AX*��B�R*�X*H*E* B
�D
�
�D"�V
�QH* �D
�U �AR�b�E
�  �@X*F
�E��E
�A"�EF
�`*`�E �AA �@Tb*T
�Q  �EPR
�QP
�Q*��b�@@
�
�
��F
�@*�DX
�*`�EU��@ �D���H*��X
� �@X��P��`�AH
�V
�@��A`�A`*
�
�R�����D`�D`**X��F
���@
�A * ��H��P�� *
���@H��A��`*
�  *F*���DX
� �@�b* ��`*V�*V"� 
�DH*`*@b*`�E��A@��AH
�*���A * �H���
�"+?�TU�pQW��*�� Uj���TU� 
��� U����@E_� �*�@
���
����PVI��KOdA1��` �����aO� z���9��!jśs�Ю�>Ozހ�:t� u��띭;kkZ�d�D���Zʃ�B@�k� گ�
���� hU�h(+JV�
��!#EZ( 4(H�@֔�   5�QF����kJ�\     �N�B�TR��q:�o �t�>���=�^�{zQ��Vk�(寽gG�a�d��`;�F�����'\ Pמ���`;�򯣻���C��c�1�������mx� 2�{��� {��5
��� KB�
9�ZP�x���>W��=�}�������Q�J��8=�|�������:o��G�Oi�p==��C�a�� ����}<�=w�[6� ���á�X:n�}h|��/gs������=x�z�C�o�Tp��4H
_`j�E7���Ϸ��e��>��zt��`iN�޵B��/v�)�u��<Jt�<����Jzt짦��gG��ޱ�@�kJ
 ��= 'OM(9�=3nOJ{�N��{��S�y�4AJ{�4��r��z�@���A�:tS�w=4�� �<4 @ K@ 7 \����bh�M-��|y��� =]�����CC�{�v�;J��o��}>À�@c�`t����e�dx��;�.�����`;�謲x���>����� � �uY���#% j�1�j�^>���@�Ӑ�<����/fm�A�`�|�@ӝ����ؓ�;g�d1�Z ��<�6���xYn�|��á�`���7�Z)���{{ �`�{�  ?BT�ԩJ� hت�Sڨ0F3*R���R�� �M���ڥR� �4�j�5)J0  �jT$F��x�����X���������}�}�Ͼϵ�  *���� �� U?� ��� 
��  U` *��_�����&�n�O�%WN����珜aR5!M�e8<<<Y�$H�a7	�z��_���%3[9�9�|捳�Ͳ�����XF%"V1��%X��$f�|_&��/�6�asP��[n2\��1��Z�	���8a0�֘x��a�/+(fC[?�x������&��Y�B��6�)����y�ĻRƐ���6^o��g�͞��.����o~�ږ��3n��K+���kkB�d���y���K�&�6rn���:��cK���D]���6�#��\�M���!RP�%�.�d���2O�;q�[�TA;~����ia��i��s3�m�y�I���B@�2�Z����a���M߾y1��9����h�b�>[���o�L3�ˎ}�=�+�k|���rg7�k��#�i����P�T��9)F����(�L}'�o5�g��7��Ǜ�5�a-�Msg���N�5|<SSÏ��2o��4�%]���ϋ�O��>r�����
dZ&f�I廄�'���¡)��~��lʹ��k!c
²�'���HM4�q!4�/��ω�W���y��!s6B�dO>ߌ႟�>��z}��a�ŋ#��������e��G������3��a�����������zI.y
��l���$bh�W0���%�\���՞>�u�5|0�Þ��o�|.�H�n�����S=�x��=�5�j��ωq |f�zJF���h��HP������/���(��6���!�����M}�<_Z���g�|��]������w���PHL�+f��}>כ2�o=��]���d��fy������Ʊ��/��߿y�Ɲ[��
w9����_���5{x^N�&/�}��~B���ၝX`,k&��z��~:�}���!����=��͏2��5���H\e�5����<��}>��]���{e�ÌI����Ѻ_�f�S5Xl�}�>]y˹w�������K��?>�
��?I?p�?�O��#�~�߰��J��r�w99����/����"c��ڛ��~�ӛ�g����'��0ó�c��;'���	�}"Gc���UP�F��a4!w�<י��78�k~������^(xo>����g���5��M:�ueIBn�<����2�N�2��_�ߟލ&�����O��꿐�l�gq?�︳&0�kϳ����n�M�gQ�~��~�sz���d�	C?���=������4zN}��'!�YV�N������uc����I�q�;�8i�8�ݯ��u4.�]�B��z� ��wG�}��~�RR\IL��P��,�I~�]��c��ٺz�����!k�C@�4n]�!I���y�5��� Si*�E.RQ��Mc�jB��`IJ�`B�D
.��;��I�.�\�?�'?��S��%���t����}�/�Ƈ��]X%�~�z~_�a���pNf���9�����=�V{��߻��<�ɰ�C��]�˓��$���5o��y��]�S���I����S5��&���o\���#�5�<��M.`B��>��@��l��:7tFr���\	L"M^D�ݘ���xK��B��H0a�f����^���I�?��?���C�Ϻ���;��jR�������l�f�I|�כ!��Hq��rp[	z3��gɿ}��tS<��Q����ą�Ă �L6!F��$�7�7��������1����o�K��o	�I5��Nx��kws��Ë�Ĕ���Y�.��F0�m˴�y5��羙�B�Y�=�����J��ae�|ׇ7��=��K�a<<�<������K�.l P��K��Q0�XI.�W4m%rd�!Yc%�Iq#,�H�&�u�#�,7x����3������X>��g����/����p��RY!B˞Sr���<<%��d5�0c��=�I���'��|��n���3_۟�~��~>>�9��o:������i�����%߸����{ۜ�e�j��~x}1=�៍y���l��%³[�M�ѯ���<޼���Ӛ�^C�9��	3�SY���>n<|�|�.f�Bja�}�{�!Ys�~��<�i
h!`T�!T�#vB��.VQ�e�®J��8�����*,Y Jlk`J��B���)/�k5}ݞ�!�,H0j�JaHBK�jȼvC�o^�7��F��ˢv(�Р�ڿ������rÁ�g�-��%ndd�S,�\ ��	C����7i.�\�J�e��fs!�)�g/�))����TÎ<=��W!sN��r��ׂj2$��"B���49ߌ��1}ȿ}�2>����H	sY�$,)��M,�4=8pcLѷ�����z���	p�.��4.�%XY��t$ФI�]M$,HB�)!( J�hL3|7|8o�j�ny4f���g�#rn~�w��/����>{'Oϻ�~���fB�)|��瓼O�Hib�'m��@��.I.kl���t��0p�$� BP��5�qJD"���L4V,"H�pӳn�P�Z&͚6s��ǁ ��vS������ �1֡���Ô���8D���[M���x{��� �Lu����9�<�S�n]$����/9��X�
{�nP�B��1�!\t0���e��uB���4v���gݓ��2���\L��K6aa��7�~��<�=jBK�	�����f���U<�,%�;Y��}��au|�y)8�	��� ��zW�of�M��w�\=��p&f{�,�xhc]y���ߚ�'�籘�nxg����(����È��~�;ޟ�o���\�ni�Д湜fN�'�߅1�5�5�~��[}̌7�ҏ�6���4"HA���.^.��D��.R_8"e��urs�؎��*�ӟ!5�n'��|�K������>0�t�Ս���u�g��wgف;qkX�3�G�����߻�Nǘ��t?3����}�y�yɬM���ɞj<�7Ze�l,Iw<M!/��q�	�u�Ϲ��5������,u��9�݉y��ns�n5��a���?=��7帛�����}�R�nˇ9C��0M���3�<�/<�BZzf�rl�%3���O{��5������P*!ܮ�gbgRmZ��;bR`�>2�5c&uv�O����1���o2�P�%�+|���>���4q��˿_��~W��g�8/�l��?_�~]�k3��9�_M&�qI�>/��}�����#���٢\������13fG��	�2Χj���O����ܿ^�}��}�`}�ߍ>��N����9�����џ�e�O�>������։W/л���fxf��џ{�4������M*/N�<�Q2;9޿t�k���S��]޵�w.j��|�qM�1f�o�>q�;{�[h����9>s�~�~xL��ٸ'�dy��v}�|�ךMw���D/����	����xl���C
_�p�f�9�߾�{��,��ԙ2vw~�{}�\���1����e뿏������g�5�>�������o��і瞲����B�P�!w��g����Y澬"���
�����\�OSR��[�>��曃0a4xˁ�h߬.1!&��w�s���ٿ'����L��%��w�;��>~�%���~�20����2%�KH��؎��D�j���������[,�Ǖ�	�!,��?|�-ީ�Y�w0�7��8k�&�N�f�p嶖��Yu��N���'��p�g���V/���}����A�>�;��ǆa�Í-��w���eOu��>�Y�{	��&[�̼�q�>ᖽ��)�5i�/�����N3��7�5��s^��Z��GY�3��+��g�,5��(F3��W؅��_�k���z��uN��7�;[��<珆�/�)F��g����	�9~{�.%�2R�۶S��%ç��v�ˌ�˄Ǆu�$a�)�%b��K�k����5=8y�l�B� ��/��8�BC]�5���i}Ü�f�]2����JeRj�Ys�y&k�Hq(bFeU�d�4˄)���H���� Jʓ��湻������<#s\�$�<��d_<޾�F�e�.�q8Xx���8�ϵ���D��[�(P�:K�5X(r��+M9��/�f���i/�߻��~?u�15�&�w�s��d���^�����~��f���<��[�G[�ؙ9���r�s��m6̈́�a-���g�>t%��#����!5c����-p�0���x�3�f^rp�x����쬷M!�F�鷏<%4��a������ևz08c��a��[�E%��)w�!RB0�`P20p9
a��b��L3F�i�8��nk!���f��NB2槗����N�u�����ҝ�'�܇�k������]y�5�_��A��΋�r�����3=(C���s>ÎȒ��}�<ך�NT8}gGy��w���d��ɬs�u�����|�՗8ώc I�r,�a�-�		I��r����a���*p с�"E#��>�7L���D.CXB��ީ��*B0x�no�]{�y��-�1c�f9{��7��+�L0�Ϳ![��
n�Ͼ�>�ݖ_>������5��ţF,�4TƄ���Y���6v����Kĳ39ͥ\��a|&̆˗4��Ɓ�����I	/'*�P!�����Ry�6�dH /�H�b	HT������8%%^�~O%��B�D�%�4����|,�_8|��L$�7��
�<ԕ#t�\ CD
g��}��G��0�g�<�����jo�����aᇡ�=M�y���'8l�
pq!�*K(JB�|��&����1�!q)���ky�K�X�
FA�9�s�%5�ԇ#!�w�ir�,a(�&fl�!|xĦ.�<8M;٢S�%�]o\޷�����Noesb�͇�>��߷��w�|2n��޽��t�&^O�}����1�z�w����:���?s����l/�?~Y�0L�۽k�w���kɋ�,i�^p���x{�$�7�����r��#�F:H`0�܆���f�����zϔ��L�u'���W8�?��g��T��8�f�a�wxk~�ޛ9�:!��$$�$d{��f�����~��6y�}��x^g�sSd��P�4�HlHI�\1 �Q"!��L@�$�"����%�aS�BD G��T��,bFbXD"��LR�!�4fk~n��='!w�sϴi�pѳ�=��<9yĔ�ߚ����®�Wa	������O/7<yf᱗{�M��ٗsy����#��9.S���[#�<X��q�a�����\�g�Sv�t���l1�\,*\6���\�.GP����Șԅ`B��k0�y���hѳ׌=��Sc�L=6kg�/�����O69�R����ֽ�F��Ͼ�&��R8k:�c7s���a�b�����0�O<�h1��χ��0��N�$D��<��&�
jSa��7�h�]���$K��z6�/b3Y��e�9�xg�n��9	&�^BJ{�������UUUUUUUV�ꪪ�������
����������U���
��Z�����)�э�U�-*u�byZ�U�p[^�ظ n�ݪ�g�a���ҕ�����Y�l�J���U��_ ����������Z(��$�e���r�E��VU� �^`��T�E*�[���I���%1��ې��s,UUU!e�(eAa5����/�9�v�6yd�Fԛ=7H�V�M�*ܬ�M{�j��Z����, @�����7D��!͌��x`�8T�p�������R낫�g�Z�Xsj�:ǖ�5�+�a�ʳ���ސwSk�^7���\��9��l�|�l�Yx���Jf3{��$��+8��!J�5H�=Ifl�h�l�����;�&�B `Z�-T�L�n�X��C=��x=�\�W̶��LĶV<���g���DuF�4W���v*�`%���T7"�m�v�xm��ɻV�Dv�Z���iƘ�	ϒ�F_lc1  �1��B�eB�P��M���U㱛����[UUU���/O��*ʀ�t�V� ��~o2��mU]�D�\6��6��D	�U˻-UmUV�^�x.!��<�ܚ�فj��%�a. 
�ն�6��"ۖ֐�8$p��5�ˆU�5P�<�j]�����aK�5\�ñ�3��تtpUP{P�:�6]]�{v�59�V����`'�T�����qOm=qR�/;M6��N�e�t勷��̃�JK��n͒��dӐ[	}0�#��k�����5#��w�6����;FǷ=���7Z�T�fK���+��m]�9��E/[r�Lvm��7bݲ	�]�Z����{;��cF���Q��n�A���v�=Rq�4JU�8=:��k���֧��7y���I\�@��@��`{5�sn�6�7"�-cBn�v��n�4��V��0Sɔ�U�US���Gr����\��X��\Kh��`L�i\]����چ��Ix-�VӶ�pVح��V���qE��q��T���H��TJ��b ��D\�,��vgEUc�a�\UUAE����I��"7o$�sxj�dU�KX���b��v[rKTj�+q�0R	`�I�%,�B8y*Wd&R�ɞ��q;+Vl(�]���(,]pvwP�89㜵n�M�z&ns�<�h��͸�°��pa`�W�T����jkV�X�6QX�7�85�4Jr[�es5prk�]!���j��$��<�p(@��lD<�V�U�6��ڷ=�Y6�OOe�*�ZM�}�#ʴk�:.��ԩŖ[�	ČKU��n���8P�b��T)�f����*�W!k�.,%�7��YVk���a��֭�cfU.�^IiaG���m�f8H�Hʫld�,���MR�u\&��P�Qғl;m�l�- 88�n2m͵��D#�fN	`�ۋzygJ�l㴛q�X����-`&*@+��):Сj�.,;D8���'�\Ә�U棂� *���YQ��؛�h��*"S[]I���:9 ��S���d3���{A�^����Mlݠ�y@���g��uVz{��ڤ�*k�EZ��.�G���\e(�.�X�A�պW[x�DmH�1 P[n��l�֐�u7bx�ZE����1U�\�6f�zۘR�F��eMeь��v�R *�ۆ�d�8�Prp�:�OWA9^��As�!p��V]&'������Իl�v淮�0-�d+m���칌X{m�N�Fܦ��kvpu�V6 �\u�HlC(�Tf�*�We ;6xҶ��qW"��C�gv�9�\D��[p6M$�¹of[P�:���VNd�/��1�b�F�7M�+9�٭�z�;b��
����F"�U&i�� ���t�-PK�L�=�K�&Tc��cj� ��Q��9ʻ:��!����%�'�P���^�9y%k(6�U����i�����,ԩ(-�n!���h�T�v���+h *�Rh���C3:X���ctx�=�8I귭�+h�b�����CM��|�\x@&ҭ�����f:��#�v��:����붰� YmmTk4�������i�)e��J+����
M
��-��X��FE*�;Gpj15V0��&F�7b�p�ଡA��!��5��u�Q��Z�g�:��.���D�"qj�I%�:���)ѷ;EN�S��;�v��S��B�)�����mf�7Y��c�n�#.�$�iEljVmcC�כ�CAEV4�6��H_c����rM(>������Q�76�VGΛc��U��,�W[u(h����.�U��6j���j�z�(�n,UU���:zڕ`�)f8�Z�c(�1�w^�g���j�h���jB8�:H@t=me��n*uN-���x8�""��*W�h
�YݒU�]�m�UU]*ѩ�v�&.��ѮJ��lԥsA�/U�O���Xx�����ڭ���x�B�&�s��V�+�uQd�:�ud"��V�0�� ��Z���6�=�j��
����������
��P���m��Ukevg��³Ή�j��c�m�v�W�:�ڪ�IǉWl]K�mUU*ԫ�W*ۂ9&I�0��&��[ T+�Ғ�uMXF���vثj��e��U���
Rv2��UA�n\pl5@�mUUUUr�UJL��UUW���.��@UUURL��h�V������UUUUU��������URBv��+Za��݈
ꮪ��jZ��j�
�ԫ]UT�AD�=i]�%()^j���꺫�@#h�Leb[AUWOx�퇷m�	�嶪�u5r�1t�f�V��U�u�J�m��Ԫ��[Uq�#mR��֪��8�L0��[lT{ن֠
�+r��[cPŵV���`��j�V���52<n'nq�n˦�O2p0KU@R�S�D�5OV�R������*��*�V�� RS`-���cUWS�3lwˠ 0�k۵��s]�I;��j�����퓊nl/`�r��k���R��4X��p�k.��Sh�᭩V�6��rxV�$:6��;�v��;+�-l ��R�ݧ�k�*��rښy����۪�ST1ְ�	�%���[|h:ڬb��V#vR96b�Pv���˰���%k�M��Ĕ6�2�|�Z�$�V5����f��>Ɠ=Zͅj�3�1�F��IX쪱���M��b�v�y�����D��UT2ݙ�ۥ�j+��x ��c�!l��mN��6�k3Ʊn�-ۢj��ؔ�������N�:�np4n��i�@�k�v2 �m��V�W��U�Y�R�(7!X��������EϞ�B ����;A[!;JI����na���N)��CI��˶66��)�ڪ��m�tt��eCs��˵S�울G8�5�Unשꎸs�A���877LQU�P-Vv*V]��*���uU@*�UW,�O^�/-��T[�R�*1/-R�UUM�Y��\T+˻/��v�Q���T�����/U��P����U�*֨����ę��TpGV����SpG�N!�j��nv�q-�uB����lM m�iI���1R�^8� ຩ�26��XZ��ڨ7S+���U]UA�WV;��I�MT��f�j��!�%���Ƹ&�ͦ�Uck��t�]-���3a��Gc( �f�U�Z��f�����ۭ�a�ò�U@U��]p��*�b����v�\��t!M�Y
��
Y`�\����1p:sUUvl�Q�G���[WUR�QU�*5R�L-�+j�ꪔ���z(�[���[�x�� �͜�MU�mUUEqG����5B	HQ��UVԀ+PV�r�UUR��hᠨ(*��U*�Z�1�ڕv�������U*JT�mUb�*��ch�^ˆ�T��a}�� �� ��j�fם��ʴUP�ӕ�ۜ\,T*��$��ە�^]��ږ�v`�8% UF���V+�=�UV�l,�&�mu��W�n���MU]T*�UUTjx
�����h
����b��+mU��E�5W/-\�@e�R�C��0��om�
���IdiV���UT@*� ���*��<�>�P%K�T *��ň;!i�����ɇ��l�J��UUUUJ�UUUUUUUJ�UUUUUUUP *���PPUD�Z���UV���h
�����j��^Z��������*�`)�FyM�UT說�
�۔�y����
���U�LWm�T��0W-[UuUUUUUUTґ��Ë�f���5@\쪶�U�U|����7:�D���`*ڪ�U"Z �AUTTUj����V�Q�[UUEUUUb���mT [Vآ�����8 �-< ��X�`y��6�)B떫j�j��)Y�����o^�٪�Z[��S��y�iV��uR�6�Z�j�Z�����
��
�����L�p=��9�tu�T ���J��
������y\kf�+j��#�����b�9�\gP�T#Z�R��^r��<̼�6�]�l+ͩ��|�Q�m�%�U[ek��sj�i�yg�M���va(螄ȇY�a��֔U��D��Ih����Ԫ�U��sU]�J��һ�j����tʪ�&�:�4�<��P��3]5�z�9ܕn�U
�w�����p�
�rb�z��u���wS�{�J��1�r�8�u����T��F�V�
�Im1-x��b�.@P� -��UlZQ��� �ع^�H��1n�Y������Ś��S�L7am��j�ܰ���V5�dL�1Ce�X�Z.��� U*#�
�lT
�a�(��"?� � �� �`����GH��b$�@�p� SZB�: �P؀��>	U�=Q ����"&�1����6�D8���J5D�! x'�T$@pWh�&�����)B�G ��
x��_6��π6��	�_�*�+�+�@���� ���訞����W�F!πS����)!�<@؊mU ���_Av���Whx� �|����AM�8�
��*z�����`;P@���E5�"C@�1G�Sj�A�P�pt�l@�<t�|���|�R��� � �Շ�T���PX�XȄ��H�b����4�
�a�@aV �X��)
� ����P�B,���Dv����ʩ�bx�DKY$�F0���#"Ā`Đ$�"����"�_D
��"����#�'���]$�0b�$��(�
F,��E�V��i6�zmP�"� � z�b�a��F� ؅���!)l�Zȅ��`1���H�RR���J�4�8C�D�=F�FAB,U RRH����@<t(�P�~PSj����*�T8	��@ _���1Z�-k�	J�"�jD�B+JF#�aH���q
��+�V�}�k33UN�ҳ��ݗVMkjn�:��M�+i`��p���u�Ms5�:{�F����f U��X�݅�SHI�l�h$%(;<M(p�� �W.o=�*����Ů��H#�N���,+��Cnm���xKbm�&�cp���,�\��{��	�lsB�2�RYcKq4��dݷIɁ˓� �8{�ɠyy\�;M�1���J̖X� 乄+�f+ܡ�1�g�0�Z���+�s�4�����ui2X�8��0nŰ	��ö;Vy2�V���ԧ8�U� �4�"6�^{(&�{(���8�p�F�ؙ�-X5�VZ���o����e�&5�j�7��ۍ"�er���;a��{F�s�4nʫ����y�2����;Yz�����C׶%�"�R�S F�dfb�J�5�ME�P;��c��}=a]�8��ucn٥�-P��l8Ncmp�/GW9N5�����Ŗ��V�,�.nt-��r�.q�$��vS��c��^Ch��5v��1��B��+u��B�l�]��ve3��K��l��n��8�m8��2��[ę馦�s�h����Ö���9��A��ZJ��9�F(9�&-�m�p��E�⁩�p#la��`δ��ÚLէҕ,T�k{�s����e�Z)�Ɛ��͒5��8�!�Ǳ��;�&�۱��jM��3c���Xo/��N�L�b$�v�����\���7a���Syx��(l0����7Lm�#�31̀����P�wZF�S�����a�`Ldg����Z]õ�Fp�;����y��8���<��s�������ΙvUU�G:�7KlY9v�N�0ff����U�Um*� ��V���YP�`9�(dPR��t0��݁��]#T�L��v+�J`tv�gk����գ"`}=��zsOl��zҤ���'X�6�f�v��i��iN�r;�N���rE��b�ɻ5��P�1�F�%�Ή�F�A�(!��Q⫱N�~E���'0>A� ��q@� b�Tl����f`7�5x�wn�B%�n�utnZ�G�lzw:ۑ�8u��^�IWXj�6c��	I����*��؞�c�ss��'W<����P�g gd�.<�pݍ�9�ȼ�'�G�jG#�G&�9��q��k^,Ș��p��荄k-�,�2�q�U0�J7�;q��=�xT���7r��@s��p�N�!r4��fͰ��
jt��{���M(��f[��$˙e)l�	BYDܠ��C��;>�;s���c�X�k�2�v��}�޾�Ù���������3��4]��-v��ڴ�f��WK���<�Ah�M�ڴ�f�k�ZWˇ]X�c"����4_j�m���h�M�K�dqIQLNE��4]��-����h����1��Yjq�ݴ!�B�\��L1ܰ����kZٮ�2얠h�˂�k�uX9~�?xZ�S@��� �٠}�@��a�Cp�H-�)�f`����	�!�@����%� ��s��3�̐�w����@��-�o��6�#X9�U�zm�^��ݛ��ovn�m�>ra=�R�LM'�[l�-v�@�ڴ
�k��{�W��bMHۓ@��-�j�*��@-�h�f^�[�)�[�Ra������`�;Is,B��ޮ�X[��I�h`sTU0ٱn�m����h^נ�4]��:�\:�ŋM���*��@-�h�E�~���nb�w���e,��mZ�lܒw��$����w<P� �"@c	F A�Ũ����&�_��7$���om�@�I�rh��h�M�k�m��T	)����E2-�j�*�� �٠Z�[�)��\6��d�m]��L�2m��3���;>���\���XW��%mD�ȴ
��@-�h��h�V��U�o)#șkIǠ�7��s3=����=��-�k��w��H�ĉ"nM�r��j�ٙ����6����o����J;,r�W2-�j�*�� �١y��Ü�
5���z�]�9|��>�2(8��ŠUmzm�@�ܫ@�ڴ��#"q<���)'����zn��uB�l5R�RhKP��zw1d5�5�\��b�%2cS�7#��{�@�ܫ@���΍黳���v'"|�H�u�S�M�r��)�Z�Zm�@��%2�a1��S"�-���կP=�����է}���.H�l�0��3����������k�V�m��?*���8(I����m���Z�ՠZ�Z��.��n$n�+��t�9��������Yi��ٲ#���MX�̖� �%�B�k����˂��a���Z	{�V���M;�� eؐa��j�h�q����.�D��h�LB+�S�kfi*����)�J�l�I�%tlkC^
�b[(���SR1�T3BZYM6�՛q���z8k�n@���q��78��
�i��ZK�n�u.�Y��h����N�ƾ0)6�� ѰH���j������ֶ�C�Sq\�b�Q��K�B��ǭ�/�?�����-���ՠu[^��Vv� ��J�EeT�o�z���ŋ��Ӎ���=�r��>��,dPq7��k�hVנZ�U�v�V�o���k�����2Zq�I%�������yh�S@�ڴ���M&�rAH�]ʴ�)�Z�ZU����33��} S	�)$s+״��E�8��v���u��؊�Bݬ��8��$�Ly��2/�_zx�-v����5,X�7�5i����H��V�7	!�Z�[y����{�8`a�J��Z��X�RW4�JS�qd%$	�hCt�f�@����B) �"?:}�[�u���yh�S@��η�)&(�����:��@�ܫ@�����^��<�����,�q�ıf#v{<��O�ՠu[^��Vv�"J)������e4_j�:��@�ܫ@���1�h��2!Q�(Z�	�K@�"�M�U�u��
ʝ���N$$2(��C@�ڴ�k�-w*�;l��m��$�71���NE�u[^�1#�~�-��Ɓk�hw�*z6&�$�@�ܫ@�鹰�1��D�UY��5�ܒ��z�T$���%"�L�@��ՠu[^�k�V����=�M'	!�Z�ZU����h�S@��F��dƌnd"Q�v�]�� ����/;�oa瓷WF��d�͛
��\�����:��@�ܫ@��ՠ~�!*��ō�#�@�ܫ}��H���{��ZU��UglS$��<�dZk�h�V��mz��ZF|�C"�A�Z�ՠu[^�k�V���}�\���O� ���r�I���%���L�C+rӍ��{Ӎ�Y�n�Zu����-v����0r4��$�Bb0���M7�l#����΋@�d�r������,:x�S�i6(�I ������@�v��j�:��@��ŗr,	Ƣ��dZk�h�V��mz��Z���y�'�I8�9�k�hVנZ�U�v�V��U�o,M��H�18��k�-w*�;]�@�ڴ/�Ņi8�.,n9z��Zk�h�V��mz�8s��gN���U2Pl�ͷb�Q��օA�V\�u�Q#�`!E��U
�%J�i��8n��U��܄<��P������)�n�i���;]���ZT���ڳ��C�W,Е�5h�l�t��B�a���/�4�ۯY�h���<�V���'> ����U�v�]�M2m���� *���c��/nz�e����qc5��;���Ӊ'FgԳ�)��ҁ���9x7V�K�ɞ)�F�Hڐ�W*��W;s��I��M��|��Z�ZU����h�v�	���7#�@�ڴ�k�-w*�;]�@���H�8���ȴ�k�-w*�;]�@�ڴ�t��؛D$�R=�r��ڴ]�@궽�K]ɋ��DE2-�ڴ]�@궽�r� �>�}U�,e�a3u�V�%��LTS2E%��hڸ!�L�9��EΚ*7a%� I�k�hVנZ�U���s3F��t�o��zE4�N�,l���}��k~/� 0�(#D+ �s����3�u�U�_��@�ڴ��LV$☸��rh��h�V�k�h�����(�mȱ'�̋@�ڴ]�@-�h��hF|�k���Z�ՠ�4]ʴ]�@�9��,<��R\,��\]�pv�&��×�:����mƘ��&�)�|��<@\�٣�m��zh��h�V�k�ht�S���B'�7&�k�V�3�H����ovn�m�{޼Ԗ��x�2�c�L�@����]�O������s!�n����f$�X$ Y���\��#O5����WG8���Fś_9�3�0F��F�T�x�����᫨a���U�'�=��փ9�͋�n�ޗ���f-��y����<�&@�v��́���0�p�!+d3{���!�|ai���Z��-_�%�s����)�7*��kr�B���l­מ^2xfh���3^Fq�|�B�I	+l�� '<ֈ��f3G>�,�8g_�������'������#�/���HLq�0�e��ks~���0�;�6!�X,!��X����C�*T�`�+Y�)�s�0���l]�l�5�S�������͜�[�h4�� S�y�(��S��<<T>H����F�5R1H�@�#M���	�
ASH�P�4��T" AG�&���nI���ܓ�{�nd�d1G $�@�ڴ�f�k����,čۺq����ͱ�TYe��'�[l�-w*�-v��j�>}=OA��<����xEM*qΚ�Y��b��X1��j���Di�q@ӏ��&�k�V�k�h�W�����{�@��/���"r,I�s"�-v��j�m���[��Ċ��{��4�H�F�qh����[l�-w*�-v����&4A)�P�@-�h�E�Z�Z=�{�9�p�,�<Z�j`x���s�����=����B('�rh�E�~�ffg��?�;��\����`��)�%jX�;�܂�o�J��n#e�{d�A`x�2[suǮ�Q���;��-�ڴ�f�k�V����y�$"Y r-�j�m���Z�ՠ����R
8����m���Z�ՠZ�Z~�7�Ĝ�\L��&�k�V�k�h�V�[l�:��ؤ�L�ŉL�dZ�S@�{��_�=�zh��]�=�H�F��bJd!���NQT�����R���O<V÷Vnt��[��@G�08�L@��ll�1��J�]H�<�퍐��V�.R�IK[����]�Θrjb�u���̑�P��ʑGcu��K�*l�q�1��h��C%��In߼{7z�P9��W��6^�mٰD�0�����lG^Zk�p271��g�٬�b�;T����m�T�!(�mB���$��%���|�9����RfP��Q��҈��K[���N��[-�#�һ��݄8���Nu��@-�h��h�M���	� ��"�m��ՠ[e4]�@�s�َ
@�PRb�M�j�-���ՠ�4����rb��1��R-�j�-v� �٠Z�Z�����q�D�I�9�k�h��s1{������Z�Zoj��8�R$��"M �c�{�U]6(P.�෱�rmv��m�N���Ni�8�rF����m��ՠZ�^X��΍��Ӎ��z8��Z�0�[k�@�ڷ��3���3���HW�����m����I`?/m,,N�D;!�{ޞ4�ڴ�f����q|��&�G��Nz�Zm�@��M�)�w��z�(���ȴ�f�����S@�]�@��$����٭�VVZ�a�m ��;n:l�g��	pn�����fh�FpX���K��k$s$�}��@�ڴ�ڴ�f���1rRb��18��S�$Z����4���?[[x�&La4�ڴ�f�~�9s�#@�!�#P���D�$�a�dd!-��؅���D!$� @�白�rO{������=cV:Y-##%8ޠ�ݺ}��@��h{�����v����&.&9$rh[)�{33������Zm�@��s9{�o�������� ��g�,t�P%��6FY�WM4,e"� ƈ��_�I�&���ȱ(�q|����4��Zm����~A���\]X{�4�8c�D�}�j���g3�������h���h�M�39�q#����	A)�؜��m���6����8�X����}���N |��lj++h�[*r�ށ��OK�N ��}�����	>P��E��A�ࣱN���s��9m���
�sEtj�X;l� =�sϽ �K�N����@��/ ٙ�_���dj�Jª�G��n��Iº׆1n��Onvf���Y��O��\x-�� ������m����{ ��{�}�K�����ހ{E9TuJ�%�%' ���;�b������ �~��ހ}'�'6H��"5���9m��� =�o {���MROI�' wv��x^�u·c�e�^ ���ހ|Ox� {޽��(On���>�U�B�X씕��I�I�V$�n���� �����o��[o� ��" ���-� �t8vW�\Վ��a��-�[���� j�qfM��^!v���RS �дfXM�3-����]'��x0nB�1s!��x���d���`���F5���:��vTK�Z��jAȼ����r4�ۅ�ɋ��n��k	fQ;`�]VR�䧭��lQ��ղg���u�ۊ���f�:ܚ��u�!�펪դ�M]�v+:wO�:O/��Ŧ�bj�Vo�x����7���di��k�I�3Ў�UP,bQp�f�ՙ���~�� }�[���<���������v�Ⲷ�ղ�-�� }�[���<������ {���@>�ͣ/FU%������<������ {���@�z� ��#}�9amn�e}��bJz��8 ��� ��x��Rn�u���h��r�	B9	d� {���@7$��`��|��{�p ���-jR֣��fJeեsU����q���2�8B�tv�loΥ�N#��#�G-�[�� ݷ���y��I�I��wv���٪�Z�(�Ye����<��/fw=����$��ZA�)��c�$a#$���!IT�`�Hr���U^���˜���m����>���� z|=��T,�;%%}���N ��^�ՙ�F{v^ ��}���RNP"
:�DKI�5fb�n����ݗ���y��jId�����/oj�+jh�[*r[ހ3�z^ �K�b���?� �~�N0��׽ �}��*��e��-v�e�k�.�vy����a��l�1�Gi6����s�6���O.J�-��﹯� �OzN ������� ݷ������
��j��e}�������$��~���z ��� =����%$<x�N�j��#��N �����oQ�"U`�%�"Q�"�A��<�;�?~��Nr�zO~��3��r'�I0�[m��q,�{v� ����=�8�Vd�w�{�h�j�%E���Ym��}�>�R�[�'@w�{� �޷�~�'�$�PUQ*%t�%��l� W<t���^#��GZ�o�:CƮ�����r�R����7d� {�z����n�Y� ��5����$�HuVGd� {�z����H�m���k�@>�ޓ��d�=�:���F��9-�@۶� ���z~ŋ噖ݓ��8 �o�ހ}�&���5[R�A�m��,Rn����I�' ���s�� >"�J�G�"�q.�K�s�[������ʙd��[����=�8 ~X��%~���~����<�� ��֔rR*��:�n�d�m�2f*������M��ZÛ6<�$�� �	S�ZJ�HK'@w�{� �޷���<�,_��I�' �܉�mv�L#��m�@�z�jř�Iw��ހzM�8 �޽�I �l�BJ�����o �s_z�=�p5$�)!��� {v� O�򩺫�r�R�ށ�Y�,˷�������� }�[�?bK�X�[��w�ހl��I�	$(�R6ZN ���z�,I~X�V���� �]�s���Ͼ��m�>�ō�(0�*�����!�@��W!�)J�.S ������5�@�7���YB��.nB �R\�L2�t���V��Ƅ(_$!7yi�RZ��������D1����#��ƒB�HcB�B�[<-!$���*�@HD̇��n�@!#	$����k}JJn�%%hA��
�2�jS|��H�}eR0�ٸ���3$��IBE�P���uHK�������Д�\֋��0�6R�{���p]o|#$K�U}�q1�*E�)&�L�����9h��"�����ֳ0�F@�JM\�M�s�l�F�<+/���H�.��&�ӥRX]u$�ܺL��e��:�R�bz@�	5߾O�~�q�[Խ��h~������*�N�r��tU��s]��t� 
�z��m�@/V'�;����dq;���R����� ��n�uHLl����e)i��e�f�R,�9a�WsXᓋ`N0e -���!;vpg����Ƙ��\�91�A���em*m�d\1o0nz��qAiv�dԢ�j�`�lBT���7?1���2�N;s�!�rf�<�ݲiu!��(�%�ch]�5�Lv���m��Yi����q�jG�͎٘@��
QY�]r9�숦�ò�Rv��
�d�Ҍ�&�8��j��ɹ;g&�N�8���N!2��-��P�hMhT��#�Gob����n���ۣ �&��9�+pd'`u�p����.G�<s����]+"��@^7\�'�u��:ʜbwR:tv�ΩLVA��)
�ocx1��U��x���x����B�s	(]%K�W�TQL�,��$�bFXz�]�W�F�;[�FX����9�4��!�8[�#;���λ`l��c�����Kv�ڊ	Z��Jt��ŸeZ�鵀��K���4�UT��Wt15h���l-��R.��s`��Zsɛt����uԶvr��ʜ�^zg=�	;v��r��O�� vl�)�.+�˫�s��V�kN���-k1�ћ#����U^{ur���5%P���iiYk[�5tsm��]�]@M��:{s�J�u�;͎��][��,/�����vc�#b�vF�:�PH�[d�c4e:����0ac���7h7�����]�qƵ���k�%Zxn�W^x!m�4n0�P
��������X`t��]d^1oW[�B�*��C�R� fCe֔uj�qۙ���LMWUU�HK�]���5)�ы1�j��z�N��l&�v���7�~(|i�9·�wi��!WDnK��F���Lk���LW5���2�ڄf;B*�98yw��ct���f��ӫM��
�K�kqcʴ�
�-�t[J����w�������x�*Q�_Ez���� ���}U� �t�4���z���5�!Qp�5\]&v���}xˉˡTw�x����H�&�+��7jI��LK��ظ\� n�^U��4cs���Š�I� zs�8�3KGQ�m�=�;x�Z�s�2a�Y棲0 ��.��Ub�J�D��B�b�b�g!��]k"ks��^-�dqّ۞�Z�!��e��.�5ݠ���U�㺱o.�G�بB�IJ�Svfr���I?wt���ai���SR`6�i4��7�x�
Ļ^�RhU�X�f�GA~I::{Oc�Z6Gi+n�w@��� ���z�=�j��� 7}�� ��hʸ�u��[o z����$��l��I� ��^t`Ͻ�y�b� }��0�%���-;�I�' ��׽?%��Y������ �߮�;ч�ނ�%T��k��JN�b�&�����x {�sϽs)�wI���������m�����o ĳﻯ����' ��ם �D�ѵ"���I��Ǜ��|�)v�íd͐��XC2�\,�0_�N���=���#�m��s_z����`����Y��3�P~�����F�U�Yd��������$
"�Eib��	$$!(���D B"
,�75m�~�� }�o {�y���IOj�pv9U�`�I� ���� >���jı��K��������VD�97�' �Ms��%o�4z��ڴ?��g�K��o��߿jh�ˊ�q��[x۷�����w��_�=���@����l۫,e���st;,�͚��"�9i-����9�rGGbm�t����za�n�d�H~�~��{f�w���s9����Y���o㍿~��S���)ik#��`[�7ٜ�bAo�4�|���o�9�Ďڠ4z
'��7&�[�M$�����N ����w�ܒy߿� ?{e��WT�KW9|�wN��N�3���_���@-�g��������^"d"�7"��>]�^s3��ퟀ;�zh�S@3���C`��I-��:���k�"\<c٤h��ˡB:��Jd{WT�ޝ�ah���ǜ]���_M �m����g39�U����^RV)�Q������޼�ı${�x�:����پ�33/��ٰ	ƢQ!�4y�-�mz{3��H����[�M�ڞ���B�$	"����s9�����������١��"���$G$�>�E��K1I�����߿~�)�[d���= ���s����s���>����@����>����ͬy�Ո����pz �H���.a��OQ�h�˖�fm�4s���s�i�M��,C�Hܟ�-�����V���ŋF߷�x�~���v���\�k�[���s���9��= �����w���9��$�K�Fq�#�@������i�g3��o�4.�=��X
Ur�����$���m���@��ס�fs1u��z�*ȗ�����$�@;�f����?��������=������4	��p�3/�Ա,N�[������J�pjuKv#��؞ܕ�\U��ҭ�������i]�;^�t�zs�`��y.]��!�V5r����.�ӆSM�ʓ`�&�L%%	E�xh�����(�V�b�%�%�٠4*�������v�T����������&+�FHj��
������f�e�(�:%_-�����ë13l���CX�\���>��6��d�Tv!�:��c�����;��8ͶZD�H�wfd��768��$9'@�^���;�j��l�fg? ;�zh������B�$��zz�Z~���h}�����$w��3G$mcd�dn- �o��}m�{���_;�Z��}ޕ���C��IoՉ �wo~�Z���fg���|�_b�� �5#�M�����fs�ٙ�{�������٠u
��jF�&u���b_7s����Ƹ��,!H���.vյ���f��F!q�#��^�z�l��l�g9������h��"6���W%��ܒ{��k{  �8=�'��u�'}���I��߳��d�Ӵ�cy5�GG&�z�M�ڴ�g3����zh��.��Ȑ��fb����:����١��3�v��@���z'���bY#�Z����٠�@�v����<qƙV�Cs�=��<�j�L�@g;�8��՘�t�8�Gi���t��b�
�A����zh{l�-v�g33��u{�z}T��Bb�9$�I��}�K0��8����������Y��~�/{#K�E�H�@�<h+k�`&	�HH$@(@$H���>*�A4��@yg��u�!����w�H�&H�Q�rCC��s3����@-���}�f����s}��uz�?4�A�NDĤz��4g39��}����Ɓ��@���[�ђ��pkv��SH�:79�Vu(:f�ѵ�6@-v`wG6NKH��rtU����zh[)�|�k��fg? -����\1s�LYĤDRM�e7ٜ�Ď��= �ޚ�m������3������z&�FLE )�= �m�{9�Ď�zh�������G$��ƞI"��{��ĭ���v��@��M�`(@��ﹹ'{۩3'un����#�I�v٠}l����@;�f���s9��-��	���ѱ�7Q�g���K���x쐅�#��٣�,�ߤ��X�H451C"�G'�_���huڴ��{��~@v��@/O%�#	�$ҏp�>�o��Ă�zho�4��|��%���#����k�[�����M ���=�Ļ�Ok����_�R*(+e���7��{v���<hWj��٠}z��b�$rrh[)�{9��Oy~ �ޚ��4��n3p*������A�mF$*5��2���UqaJ�̍dmhMqVn��)�M �ԥiTqt�ד��KY	�m)���`�f�*��&�P�F"D96�it�����F6�E)X[O-�����4�-����{k3�/��c�b�Ǯ�U��ps;�p��<���y��Z6�����+Z�E)(�@�4[��2�X�!.�b��:I�'����m�j�cU.D���8������渋�<�)Q�]�]��ߺIC���h���
C�?�����٠v���3���Ɓ�|����6I	"��پ�fbA��M���}�j�-����&,c�8���m���i��3���}��i�)�Ԓ94=�fqw��U���w���,X�%��{~�m����uJPv+4�mz���b��;}�~��?���DI�1�hRC�l��1���m&�E�x�-t�̈= 	ź��Y&)9��}���l�?v���s�ѿ�wg~��]�RV)��[o��}�[��')�#4 n*��t6Јvbi��)L�������MT�`�|���y����&���������9���H���bɃ�$�&��'�w]��r��ٹ�(!�W2}����=�M����6�)�) Ԇ��[^�}�٠�l��s9��b��|hz���5 ��6I"�������3�������x�?+k�?}��xH�GA%�#�mG��1�Y�)6��Y2���P����k�_����޴��5�\8_��M�l���[_�g3������@=����F��O ԎI4ݲ��mz�{f�w���3?������?��"c�$G�8h_���@>�l�bř0�Q%�H�x��#��!���&���2%�222��Þ0����%KBRB)-� X\vs��K7A�3�ؑ�z^d�O|v>�6J��F53Ә�� H��qϨ4�IMZm#�	t��Oh�s2!JF#ā"��V�a$� Aʤ+
0� �(��	��a!���0��d֒�ӹ���me֎|OKh6F4����H2�J�d�Ã��{�'�dY�P���t���ićxU��%��!���)�"JV�fa�r����1�Y �"K�AHB0$BB0&R��<�!�14ɶ��i)m�fbY���b��53�Q!�4P��F!���4�aB�"B,�F$#��r���&�t(��'���QS`��z��*z)��4? DM�G����A&�0:��&���ܓ��]��r��˟L�(�'"bR=s9�Ļo��[}4�v���:�Vcx���I&�w��@�s�Ϭ���>^�����k�>�����:4�r�U��6���������N�W�GA�hd�$�=.�z�d�<�0rO�}_������{_�1,��fF����m�ߑY$���Y[�Š~Vנw�h{�4�v��s��z���ԑlm�"��m����i�����9�7�?��u=����!1q��ɡ�s��J��|���$���rp@�Qd	"��y����j��92G�jG$���^��s9����� v�M �m��9�}g���K+`�9�p�� r%�	f��v�&�J���t$t%�6�$�_:�z����Be��*���z�{f�w��fg9������h���IȘ��@>�l��٠��@�[^���Ď��'���X�m����������ǩbA�@-���;��͘dĜ#@ܚ����s�}����h��- �{f�w���(&���b�C@��V���s������> �������M�9��9��_~��.������7pι�r���˥vFj����m)�[-�P���:� hK���1F�0�1Kn hc9���+��N��B��Z��%�xT���������^lz˪�O�2	n�� ) ��^0��\X,��e�ljP����[א%�Qbd�.�a��ҵ�FQs��0Ka��#�Jm.�D���c+׈@���>
�!��C·j�:K���$�|�L�9�Y�2b�	m���Nl��nطAρM��i�R7
u���������(
�w�m�������4��hWj�-�ɍ��H����7ٙď���@�����1 �T~jG��	8�@�ޞ4��i�fs���s������{���@�u*D�#x䆁�v� �{f�w��s�����U�o�F�a"`�Z���٘����>�����Z�W�r5ɈI��ƤeHCjV��]K_���<`���Yfa,��Z6e�Y�Lx���$�I'�}�~�S@��W�9��o���e�g�نD)�35��9���o	�X��
�3��s9��37�|��@�l��@���򸸲8��>�ՠw�����ċ}�}�O׵��9&6�r2H�>�fq۾ ���?u�s��-Z�dƚ�A��$hNf�w������ڴ��s@��u����u�6�u ��,-$x`�b�68�:�XJY���;{�!�WF�"����<hWj�:�����~@[�M��5�1��9!�}]�@��k��٠~�S}��:�V�ԑ�b��0R- ��h{l��s�9����	# �HB0b1�V����s�͝��|���Ly&&�I$RI��@�l���v�fs�[}4�.���,��&�7&���Mٙ��Oy~ ��h{l�./���b�i/Z�Ѵ&�����4�]�4{X9�E�:�\QՖ�.6��t`��Wj���h{l�3���s9��O�@���m�"BMɌ�- �{f����H-�����<hWj�-�ɍ5H���Hӓ@;�f���M=��s����x�lm�<cN8���_;��nI�s���O}��nH�! s��s86��j�X�,��o��>�ՠ{9�s+������?[)�����]u.��j��al�FȚ�"��7u��b�mɰ�l�^k�S�����1�Ș)�*��@;�f���O�f$�7��Ӎ����)%uA�Kh[N }�f�����g1����Ɓ|�����_j��'O�8/��}���f����/�����4��Z�}�@>�@���4���#Ǔ"��9��=�v��v١���3������h��m�H!&��I��_j�?�����O�}_��=Ͼ��l~�b$H�l��E1	�"��ܟA��=:������A"CYqc��謅��w\�^ݝۍ��J'�g9��<��T��j�9�2�]�ۚ���hv�ZL�R�7\]	�kY!������.�.���]�N8U���/.��za����]]gL"Xj�R���D�M��hU�f�~Ξ�-�Z����v4�e枅Y't�<y[e�ޅS�U�	���\��5��Il2h�֮�����&��%�WU�5%R0dĲ��ڛ2�N��hj8���v���9������%�W#q��������ՠ}�j�>]�z�׎��nqb"q�&���վ��$wf���ǽ������������+�(F���~��>]�z��4ݲ�˽n��$���8	š�g1u����@��)��s9�g3���;����@��K�=MBcCC��$Z�m���M�V��_j�?Q��i�s�#���]a`��a�������k�t���,���*"��I^..H�¡Q�d�޶����@��ՠ}�ڿ���s?��f|�������i4r�a4��Z���4����s߮䓞���$���}F��|��	$���G�v����?��K���U�y��:�܍G��I���?��bW���>��ZU��{9�.�|�ݯ�x܆<dN8��?uڴ��39�?{��V��������ji��uԜ`�y'wr\GU��-���NJ�L�&�l͉�wu]�_;M�)7"����|����f���ՠ|����HܜQ�MǠ|�����H���6��7N6�=�Nn%����jj�G#��zh��ZL��G�F,X�@�K� �P(d`D`�I$Q,d�	 ��^n�{��z��w�ܭ�E1�Dq��94?�3������*�����V�v�4��%��I�`�ZU���g3���~ ������ՠ�l��Ym���,�3Z��#Y`2�-5{4�gq�#he�r�dӵ�I�xP'���]���|��5�z��4�v�������%R���%�� ~����䓺��N�����y{��W������r�I4��������3�333�ߗ����{���@��Z.D�#m���9��qW��U����Cy����H�~��Z��ܓ�繟kY��Ւ�,���6�=���%�f,�J~����y{��^נ}�݌�y! h�d^^unr��d��k��AJm=�#��pi���L4I�G����ڴ
�k�s39�~A���\�|�O��TBX&Kx����9�1,H��4/_= �o�39Ď��Di�=�aj-$�~7vq��O�q�IbXۻx��{[|�dQcBo!�@����mz��h{3��U�y��³ɨ�xH�1����ڴ'�߾��>�=��Iئ���a2[d�ɭ�U�=d�v��a�B�B,�@��B1������"BA���!),	p4��#IJB�]��K�`l26]���$�Nx��)(I���MY]p�2��,���٣,��Ą�"�x������i>�7�1��$0t��2I1!�@!I�||�O~K�p@�D�#09@� b|8bA��3m,�R���SX_M�ѹ��1�D�k��6�B�Y�[w�r�P��������=��g���M�S����]��m��]���JJ���@���:�-�Z�tIV�/	������r�68���}��/Ŗ����4oLQ�!u�r�m�'�4Oh.L!�E�E�[�:]��6��qF�#��p�7�.v����K�Ee�[cO<T:[����a��IW%�}���n ��d�ڶ�F�s�.�L�F}Z��5eB���c��\MM^���۱z�:Ŵ6@�퉞�n�(�/]�Mt�"�vW��}�z��k0��H옴քJ�f4�]1I��f	�����[���h-����M�*;V��Mڗ�����79���0�D��I�8���	�<m�z�mpp�ۅ�l�唺7�4m�8���8�KiNvG&[u��	��!G0�vq�@��z#c�v�F��s�Xd`-+l�ĊvIzڸ�n���˻��6śg-�8 (�Ð��0n�tj�l�+{!��5�$,:b֠j�݄#�',�L���\S��X@yT��Dh@k�<z^<�h[f1�ɚ傥UZ��P��s���,1�-lrnN�s�*u��r���&<��2
v`�ˬtWT�b�L:Bi�X]u���B���qd��r{a�:��؄�:`���P�5�u[ý�ZڮA�m�v�N���^^ڃκ݌d#���;�F�LŰ0I�Q�M�;���[�)�j�N3=����!�8踄8��p8ڨ����gcD��d�X�Ҏ��6N[� -��*��O8 ��M����Wk�jE�&�=�r����ۆ۩�l�Ru��5�A@%��P�mۮC;p�8��i4��mm�S7�UU����Q!����jl�'$�U]�)*�qc#j7.UA�0���U�jd�癎\Sm� &��M��R�p ��.!�]v��&q9s��ը�@�7+T�V$�����i(Xñ�3��iY&�iu�ζ����f�N��E7�z���W��Sh� 3ӻ��wIgN�&  z i�O��	�)�Hx ��S�Pد���鈺(��0��I�Md�
%̤V�ê�s��Ga.�$�]��X�\�n��64MJ��7Z����eo0����(Ua4	X�x��l�-d�H���1�&N�2��y[���fS4�ݪ�9�[ f�!,��J]�b�m��;�βzu�ΌOX�mu;E��,H�ݧ�V4h�N��	3Dka��D!�iG6[FĔ�ݠ3cfѫ}�{���'�O�|�ˮ�TW4%쮳0��Jl��,,�bM	tQ#qZhV�m7ޝ9� +�k�D����uvנu[_�g?��������@���l?�$�c��܎-����ڴ��h�տ����fs*���9$�N(�$��<������v��ڴ�����*�J�F�q�{���識���-���=�s�U��z˕y6�	��I$��;_j�:��@�}�@�v��/nL1�<[P7k��@�q�;g��uGb����uۢ���8��ŏ�8A>eiڊ��o���V���_���3��|������n��v��������;�$�L"!��y3����=�}۹'��z�vbt�ȣINE�v�V���V��f%U���|�U[,m���6�@�}�@��@�}�CRH�n�����"z���-��N7=���o�bX�(��}۴�Kı=���r%�bX�g~�m9ı,Om��9\r�&��T�N����ՓR��@CRZ�K4T�4��4t�fd�h�������r%�bX�w_v�9ı,O{��v��bX�'�߻���șı;���6��bX�'~��r[�T�����.�C�<C��Ә���E�DȖ's�fӑ,K��~���r%�bX�w_v�9 lK���x�$�u8K -9����zw��ӑ,K��;�siȖ8+�Bj(PRV(z|��Ț�˴�Kı>���r%�bX�{��1���*Uw�>)ҝ�S��߻�ND�,K���ݧ"X�%��u�nӑ,K�2'u���iȖ%�oO�߿��)�B4T�O���5�b}�}۴�Kı���ݧ"X�%��w��ӑ,K��=�siȖ%�)����O��
�\�fc n�Gh�$܃qV��9ɞMɭ�����u�`r[$D���f�.kWiȖ%�b{�}۴�Kı>����r%�bX�g��mC�,K����nӑ,K��;{�;�̲H�t�[Nb��<C�<^��9��bX�%��{��ӑ,K����nӑ,K��;�siȖ%�b{�N���Fū���å:S�:{�o:|ı,O����9�lK���ͧ"X�%��u�ݧ"X�%���gs4��^	�/Mzk���Y���~�v��bX�'����iȖ%�b}�w�iȖ%��N�XIFR6�,��P�D)T�(B�pЊ�L�"�
��$d�7[(8�@D
%��!�D�� ؍G�>�����m9ı,O���uA�-�-�1u�!��~�m9ı,O����9ı,O���6��bX�'��{v��bX�+��h�U��c�+*�D��&Q{&`hR"�M.��с����G'��Oo z��f�e�Zͧ"X�%��u�ݧ"X�%��{��ӑ,K����nӑ,K��;�siȖ%�b{��%�,톡�V�k5���Kı>�{��rX�%��u�ݧ"X�%��u�nӑ,K�����iȖ%�by���Ó-��p��Kg1u�!�/m���֖%�b{�}۴�KlK���ݧ"X�%��{��ӑ,K���]ɗJY$U��S�����}�0�Kı>���r%�bX�g��m9ı �>���r%�bX�gov?����F쫼���N��N��>�]�"X�%��{��ӑ,K�����iȖ%�b{�����Kı ��t���I��ڣSlG����0(�]q0���uU��� ��ܓ��ݲ�A�qBQhLT+��n��#�c	e �9y�<��av��Ö��4.��1�]Xb�tz�݃��K,��@��E��˭ƻHQ�M����,y�5��6�P�ݷ���2#ڠ�#f��h���X�fX�d;Ws>�]�+�9�h"�&����һ[�vl棋�z�Whd����������ϧბ���їl�<�u����D�Hm+�
�������,��El�k5v�D�,K�}�m9ı,O���v��bX�'�߻�ʐP�&D�,N��]�"X�%����\����Փ4�e�ֶ��bX�'��ݻND�,K���ͧ"X�%��u�nӑ,K�����ND�����,N��S�XJ:7%�[9����z~�ٴ�Kı>���r%�-����pI����ԐI����faL$�$��n	 b}�}۴�Kı>���ӑ,K��;�siȖ%�b{�����Kı=��ݷ��][���]�"X�%����6��bX�	�w��ӑ,K��;�siȖ%�b{o��.�C�<C�}�m�BJ�r���\jGT+-��$1(���s�����n1�%���UV�%h��^!�!���i�9ı,Os�w6��bX�'��ݻ�,K�����ND�,K��w&R�"�����׈x��x���8�� 	�~��<P�Cm�Ȗ'w���9ı,N�~�m9ı,O���v���&DȖ'�����SbָOt�zk�^������{�"X�%��}��ӑ,K����nӑ,K��;��ӑ,K����{�b⼹h*�t�zk�_�gB������r%�bX���߮ӑ,K��;��ӑ,K����nӑ,K��=�&�-tn\,��]x��x���wN'"X�%��w�ͧ"X�%��u�ݧ"X�%��}��ӑ,K�����.
J���F3i�۳����4�b�Kjdf�鮙����Vx��Q�pst��f��O"X�%������9ı,O���v��bX�'s��6�"X�%���l�.�C�<C�����N���ke�5v��bX�'��ݻNC�9"X����fӑ,K��~���r%�bX��]��r'�c�2%���)-�Kը;�>^��צ�?~=���X�'�߻�ND����)�d� IA �`�@��H�@LV�#	 ���i	����KRG�:O���=������r%�bX��_�v��f!�/��$GGa`�K2Kg1u�X%��w��ӑ,K����nӑ,K�����iȖ%��VdO���ٶ|�5�Mz_���߲���7@�Ȗ%�bw�w�iȖ%�`�w_v�9ı,N���m9ı,O���v��bX�'�{�æ��.]j�̈U��\bF����q��j�a8�s���kk]�뫌�r�Ο��N�����nӑ,K��{��ӑ,K�����br%�bX��_v�9ı,O{�����"
g-�å:S�:o{��r%�bX�w_v�9ı,N���v��bX�'��ݻN@lK��}���Z�ܸX������_v�9ı,N���v��bX�'��ݻND�,K��{�ND�,K�=���X��&[Nb��<Cć��k�ݧ"X�%��u�nӑ,K��{��ӑ,KB�,B�E�DK"�bC�0 ��r&���[ND�,KϏ�s392�D�Ѣ��WiȖ%�b}�}۴�Kİ�������yı,K�����"X�%��u�nӑ,K���~mq��Қ����	��v�6��Z״c�x�nr���"4��^�D��Gf�ӑ,K��=�siȖ%�b_��u��Kı=��ڜ�bX�'��ݻW^!�!����H��R�A,�-�Ñ,KĿw��iȖ%�b{�}۴�Kı>���r%�bX�g��m�/O�,��^����}�)�e�n&f���Kı>����ND�,K�뽻ND�,K���ͧ"X�%�}�������ݒi �n�C5�]�"X�	b}�w�iȖ%�bw=�siȖ%�b_���iȖ%�������9����{�Ғ�k5�35��v��bX�'s��6��bX��/u���i�Kı?w]�v��bX�'��{.ӑ,K���	 �@����0�H���+?1�O�i9li��D�0g��[��.�4���ʛ�h�ܯ$���;X�]I-�P�mna�`����tGz8�����VK����6F�(�=��ӕp:0::�v!�1�
�y��dពAC,�=�����<��d=my��;X}f��i���k+�0d��Ӑs2�h#ʹ*�� ���C��G��`7�+9�f����|
������i�.Ż%�`�V�˵�O
��a�[�k#x�s�f�tj�m�ZҮ��ӥ:Q,Os�߳iȖ%�bw�}۴�Kı>��v��bX�'s��6��bS�:{��K�>�6΃�y��ҝ,K�k�ݧ!��DȖ'k����Kı?g߿fӑ,K��;�si׈x��x���I��n�P2Әr%�bX�w_t�ND�,K��{�ND�,K���ͧ"X�%��u�n�|:S�:S��g�[|��"�]T�ND�,K���ͧ"X�%�����ӑ,K�����iȖ%�bw>��y��ҝ)ҝ>����S䢐���.m9ı,N��w6��bX�'��ݻND�,K��ݙ��Kı>�{�����N��N�����]����津�"A��c(2���]�5��b���t��!�C\��nr���O�Jt�Jt���۴�Kı;��ٛND�,K���ͧ"X�%�����ӑ,K��;�M$D�']!-�1u�!�-�}ٛNC�ClE!�/6��'"dK��>ͧ"X�%��}�siȖ%�bw�}۴�Oɕ2%���_����������|�5�Mz~?�ߏt�Rı,N��w6��bX�'~�ݻND�,K��ݙ��Kı<�~'u�YP�Q��b��<C�<[=��֖%�bw�}۴�Kı;��ٛND�,�2'�}��m9ı,O�~�����$�;-��׈x��x���v��bX����}��6�D�,K�}��m9ı,N��w6��bX�z~��>�]��"�,5q�3q�Н�u�*#a5x4��fR]+Hl�!���@Rh�54[.�x�D�,K�������bX�'s��6��bX�'sﻛșı?w_�]�"X�%��N�m��#PF����ҝ)ҝ?���ͧ"X�%�ߵ�nӑ,K�����iȖ%�b^��f���bX�'���m)�He�y��ҝ)ҝ?�~��r%�bX�Ͼ�m9Ƌ�|�%X�!z˄�||��N�A	I�<�%��b�6C!I��2�12�b����0R1Ӓ�ܘ�1	v�
��2Swv�3	IYXYIi'���a(��ޖ��BF�]t^d@FH0R7�B�F
!���8@'�ӭi5q\@��%�=ѓYZi�FR$%aX��!(K�I.kHa+)(���W��)��
BK�n�MЖ7�y�p ;���6�	I�L�$(�
�!$,�bC�p�3	�(\K��It0�aV��������Bd���㠉l##Yik]Jqd͖k�g4�%�Yqx%:1���JEH�%�n�ki*D��(aͦ��f�e�D�!$acYee����-e��BnHB��7
��4�,����$2��T��\k�F$V��.�X$���}�$��wX����>xl4o�<t�I h$%��a0�m8���S���T#!mpQ��TM'�$�@�(�����(���?
�RMD�%��kiȖ%�bw>����Kı>��䙗��]c5��]f�ӑ,K?
@ȟ���ͧ"X�%�}��[ND�,K��{�ND�,K�k�ݧ"X�%��w��ۘ�������]x��x��߽��bX�%����ͧ"X�%�ߵ�nӑ,K�����iȖ%�bw>��\ߏS&�#9�08��$�gp�n��.[���"X�(�-1C͊�5�zr�mm9ı,N��m9ı,N���v��bX�'~�ݻND�,K�߻:|:S�:S����l�f[W�iW6��bX�'~�ݻNC����,O��]�"X�%�}�����bX�'s��6��bX�'~���˚5�fk	u�]�"X�%�ߵ�nӑ,KĽ���r%�bX��{��r%�bX��_v�9ı,O~>���h�Mf�e��Y��Kı;��w6��bX�'s��6��bX�'}�ݻND�,@�F,!�T�&*�q;�w���Kı<��e��톡54kV��m9ı,N���m9ı,N���v��bX�'sﻛND�,K���siȖ%�b~\��kS�0�Q�4��bv��{Z.�N�P�۝�k%�&m@���/A�9�-?^６%�b~�]�v��bX�'sﻛND�,K���siȖ%�bw=�siǈx��x�����6�Y��,�1v%�bX�Ͼ�m9ı,N�ͧ"X�%����ͧ"X�%��u�n����wHn��O����Afҵ�]k6��bX�'�����r%�bX��{��r%�bX��_v�9ı,N罳�������B\�U$��Y��K��2'�}��m9ı,O�k��ӑ,K��}�siȖ%����~���s^!�!��n��J��kn���m9ı,N���v��bX�'sﻛND�,K���siȖ%�bw=�siȖ%�bz��Y�8P��K!d� A�P��GL\H!	e�u ���E��{~m!���c���W�w��aҏ!�������<�W)#f.��!s�7q���bص9�G�B<�y9��۴��K87`��O5ۚt�:�$4T#��	s���[i��g�k�ҨA���>�QM��qy�;��p�N/(<q��p�s��dU�v&��m��VE���&u���wq\i7�m��ms�c��ι��Lm�p4�,u����'I�t�!���e�c.��mK��x)FXF�J]5���ڔ�%���l��6\��#t���Z���,K��=����Kı;��w6��bX�'s��6�y"X�'���iȖ%�b}��O�9��ԆkVIsY��Kı;��w6��bX�'s��6��bX�'}�ݻND�,K��{�ND��S"X�t�ɾ��l�c\E�O���5�O��ߏt�ı,N���v��c�B"~���m9ı,K���Kı;�vE؆Z�+��g1u�!�Cſk�ݧ"X�%�����ӑ,KĽ���r%�bX��{��r%�bX�}�(�6Qe��S������w6��bX�%��ӑ,K��{��ӑ,K����iȖ%�b_����A]a��0�$З��������D����`�Ǟ:����ι��+���˭kY��Kı/}��bX�'s��6��bX�'}�ݻʬ�&D�,O���ͧ"X�%���ӹ�ٗZ�SFfMkkiȖ%�bw=�si�b��D!��
bHZ1�� D!(āw2H�$���)Qjh��@�<�bs��iȖ%�bw=����Kı/}��χJt�Jt���?�c�J/ZҮ�D�,K���ݧ"X�%����ͧ"X�%�{��u��Kı;�w��]x��x��}��tP�W�L��ND�,�)"~�~ͧ"X�%�}�����bX�'s��6��bX�'}�ݻND�,K߾���R�d�kVIsY��Kı/}��bX��#�]��6�D�,K�����Kı;�}��r%�bX��o�4K���, ʦX���]��Q4jخ	R9q��۰�l��ml�m(1
 �/�>,K��{��ӑ,K����iȖ%�bw>����Kı/}��!�-��A�Ю9\�K9��ı;���r%�bX�Ͼ�m9ı,K�~;��"X�%����ͧ&!�!����Cef[+e9��,K��}�siȖ%�bw=��m9ǂ�*H	�7q;�o���Kı=�_v�9ı,O3��4�KF"�B�g1u�!�-�ynm9ı,N��m9ı,N���v��bX�dO���ٴ�Kı?C���֙l4`H����צ�5����ͧ"X�%��V?��]��,K�����6��bX�'sߎ�ӑ,A�-��dD�@���!K/���l<���<���6�vɸ�n9�#^����[Kt��kM���Y��%�bX���]�"X�%����ͧ"X�%���㹴�Kı;�w���Kı;�m��S.i�f���]�"X�%����ͧ"X�%���㹴�Kı;�w���Kı;���r'�9S"X�w��~�R�d�f���iȖ%�b~Ϻ~ͧ"X�%����ͧ"X�%��u�nӑ,K��}��ӑ,K����e��[m�]���׈x��x�{vq9ı,N���v��bX�'s��6��bX_�C���	U������*�ĚUK\��YJ�m��R��l�
���`8*����"_9��m9ı,O��a�K���L������r%�bX����iȖ%�bw>����Kı;��w6��bX�'s��6��bX�'������
uyk	lu�t=�602s��79���ɹ5�Y$�z�ǁI�&8�3g����{�bX�'�뿮ӑ,K��{���r%�bX��{��r%�bX����iȃ�<C��4��;c]$�Ә��X�%�{��u��Kı>�{��r%�bX����iȖ%�bw�}۴�H/�0I����,̄�-̹4��H'���ٱ$D��~�n	"~�ߵ�ݧ"X�%�{�ݚ�r%�bX���ݒU$����l�.�C�<Cž���r%�bX��_v�9ı,K�~��ӑ,K��{��ӑ,K�ﳶ�tP�W��Yy����o���9ı,K�~��ӑ,K��}��ӑ,K���w�ND�,K`#���ٴ��v��)��\U(&�f�5JRր�LK*Ձ;sv���܍M�;���qļ�x*qѳu�h�:�vu�<�vd�:�mȝ�"�Xm�S��c:j�t��9p�g2Ҏ�6��.���ȼr���s�,��ka�pnce�f�Еy�e����� ��;��.���&%^wcSD�0qtҺ��РҤ�`��H��4]Z�N��U�[�3mpv�U��ۅ3q٧5��QDʲ��hm�ˬ�ƋaIWa���	`nȖ����Kı/{�f���bX�'s��6��bX�'~�ݻND�,K��{�N)ҝ)����K��(��5���r%�bX�ϻ��r%�bX��_v�9ı,K�{�m9ı,K�{�[����k�)�����4�*�0���m9ı,O��]�"X�%�{�{��"X��Dȗ�߿�r%�bX����Nb��<C�<^���=��I���f�ӑ,K?)"g�����"X�%�}��"X�%����ͧ"X�%�����ӑ,K��;{�;���s��5��kiȖ%�b^�ޚ�r%�bX�ϻ��r%�bX��_v�9ı,K߻�m9ı,O;��l�ə��J�B�ͩR�`�{SB����n6�;X�:�����Y���X�2�T�"�}���bX�'��{v��bX�'sﻛND�,K����ӑ,KĽ��5��e:S�:{���3l2��m�|���ı,N��w6��P>U�i�KĽ�|�ӑ,Kľ{ޚ�r%�bX�w]��r%�bX��v��.K�2a�j��k6��bX�%�ﻭ�"X�%�{�zkiȖ?��DȞ����iȖ%�b~���m9ı,O{����4B�E���]k[ND�,K����ӑ,K���nӑ,K��}�siȖ%�b_����r%�bX��}l����e��^b��<C�<_�wM�"X�%�����ӑ,K����iȖ%�b^�ޚ�r%�bX����;Eimu�s�4A�� BJ\�#K�uf��&�%/��sjz��%���f�ӑ,K��}�siȖ%�b}����Kı/}�Mm9ı,O;wNb��<C�<^�x�zR�E��Y�ͧ"X�%���w�ӑ,KĽ��5��Kı<�۴�Kı6{�9����O#�ʛ+����iȖ%�b^�ޚ�r%�bX�w]��r%�_HČ	2zSѮ�#0����)H��B�QѰ'��|=������m9ı,N���6��bX�'L�����)LEX����^����^������9ı,O���ͧ"X�%���w�ӑ,K��{ޙ��Kı<���J���ی�Zs^!�!��ﻛND�,K���"X�%����3iȖ%�by�w�iȖ%�bw��~}\� �WK��#ۊ�y��A��Y^s�8�ՓZӴ��:�X����ff��ND�,K߾��"X�%����3iȖ%�by��۴�Kı;�}��r%�bX���d�3XaI�5����ND�,K��zfӐ�	��,N�߿fӑ,K������r%�bX�����r'�*dK��Y.ퟋkh�q����צ�5����~=�"X�%�����ӑ,ı=����Kı/}�Mm9ı,O~�n.�l+�v`K9����l��6��bX�'���6��bX�%�t�ӑ,K\$v���2���@�!N���cȝϷ��r%x��x�o��� �[j�Y�]x�K���w�ӑ,KĽ��5��Kı;�����Kı;�}��r2�)ҝ>��'���\��0�$j�-i09�0��*,�\n7j�m�71�H���%���+�$�s^!�!�7��y��,K��{��ӑ,K��}�skȖ%�bw��iȖ%�bt�ϲN�\�)��t�zk�^���>�=ӑ,K��}�siȖ%�bw��iȖ%�b^�ޚ�r X�%����z�Uی���b��<C�<[=�ND�,K�}�ND�,K����ӑ,K��{��ӑ,K�ﳴ��9k�)��[9����o��[ND�,K����ӑ,K��{��ӑ,K,N��w6��bX�'�}e�>e�X3�e�t�t�Jt�K��zkiȖ%�bw=�siȖ%�bw>����Kı=����Kı6wo�����4��;H;\�_�&P�Ҧ��yTؔ l�'<�3R�!�'�%�]��'��&�
�U.,�v7i\�sNjkR�K�	�Ȝ��W ��f�����W&C��2�[0�&A2��VH�"��t]oL��Ø�	���X�I�5�%eݸ���Ȅ`�Chl�������&�&�a�\	rP�`I!��tGno��<��.�e�}���$Hx�)0J:<��q0	��=�e�|�s�Q�Nh��\�K'9 ��A!��2<xȐѧde�i��������})==�����ϗ�K�o�<|��$���g�l�P�ޒM���F��L�Y��Zk�@|E܌	�D]y8K�%�HJK�.�5�a4Ѡ����"fK��3&R82p���FB$g�|�"ko=4f�A�I�b��ؑ�H\RSp�0�˗�X�sشL��f�A.����ɒ�D�Bh�����@�D�wv����>�v���q-[AK�1��8������tΎql�\iM��O^�
{%g&�[r�z���M[M�݊�Z��
in`��/:�͵��]��a�\�Y�v-��q� ���	F��"8��c4�N��(v8�@�ۘ62/d���v��}��p�}�W�gu�v4B�|�*�㧓9�9ux�0�v�'��[F��Z�"=�($�vp��u�l���)�b�	�뵝�4Q��	�\85s�Ʒ^�Y�v;pY
��6� 6WQ���m\��^�g(9��0��'[rNl{ZӤ�B���]�շO���a.m�Ob��N�g���S5Zp�E��o*2�F�j��x�FWB�ָ1��M���R\a;+vN��vF�:�pA��)�`���,5���m{�e��s� .�[)�R
��OJC��a��۩��*ݹ�s� ��>���t�����2P���M��#)��{U��ze]��z���H��V��v�/$q0�!���:]��z6���`��r�R�[���������2rF��M�(MB��l�[��)<4�V1�S�YiUV��gLmK4mG����:,kD�!�pn���2��O��ׯe�1�p�g"���l�랱�3@gp�n�kx���%`^=�M��su��ˤ״�����P��ˊ�W�Զ�m�-]�Jрf�[)U�̹�	����T)d�uGDoe;
J�X��B4Y�(]q�L0r�۞��;��nm� C�t��.��[�g8ě�u��M�8��֮�2��8w���P���Y^y�u�a���]�(�l��n���dnn3�AZȋ��$;N�FܻeM���r��h8�s�`ۆ�h�V���g!A�N(-��j�ڪR�UU^;"��H:�U�<f9��:�L�U୛/n�g=(1j�ծ{t�$pͯ�$d��bWVb^�J�.�ۃ6Nw�n������5ݎ2�R5]�3b�]��on�
Ͷi�҅f������L2�tkD�jM�D�D���N��;7��~�8"�V�� ��HD �X�F�� �|PNQ|DL@�Uנ}	������D��e�i�Frs���ۥ��W�aù����❶��Za389-���)<e`XT�c`r�`i�۴
q�0����l��gv�<�ۚw,�m���ge�u��T;b�Áa�9ktnړi}��� �ݖ7���Ҭ�vn[���ڔn�� c��\j�#�#�)�׌�������5x�4;k`h.ηI�%����IޝЇ��Rh��bu�Kfl��k-6�t��)0�wV�4e�Ԫ�`:-N6/��������ı,O��w6��bX�'sﻛND�,K������&D�,K��ߕ�.�C�<C����8�5m+�vasY��Kı;�}��r%�bX�����r%�bX�������bX�'g۳�����z}�!�EH"���m9ı,N��xm9ı,K�{�[ND�,K��{�ND�,K1l��s^!�!����U2�s33Fӑ,KĽ��5��Kı>�{��r%�bX�Ͼ�m9İlO{�xm9ı,N���I�W5�2e�Z֍m9ı,O���6��bX��c�]���yı,O���ND�,K����ӑ,K��.�^��U�a�����8�X��q(�yH�sr=�:�5�g�4���cʘ�Ů�{�?^�"X�%������Kı=����Kı/}�Ml?
�"dK��{���]x��x����������A̕<֮ӑ,K���w�Ӑ�LOA���K��t�ӑ,K��}�siȖ%�bw�}۴�Kı=��U�lB�;e��s^!�!�7��[ND�,K���ͧ"X�%�ߵ�nӑ,K���w�ӑ,K����_��m���>)ҝ)����ͧ"X�%�ߵ�nӑ,K���w�ӑ,KĽ��5��Kı=��EF��eE�	g1u�!�-����r%�bX~P�߻��i�Kı/�~5��Kı>�{��r%�b����jr�*��J*Z�D���KM�hlF4q��Y����6�Gk�(���zݚְ��]�"X�%��{�ND�,K����ӑ,K��>�sa��DȖ%������Kı=�����T��$��s2捧"X�%�{�zkiȖ%�b}�w���Kı;����r%�bX�����ı:gg�N�Kj$p��U�.�C�<Cų۳��ı,N���v��c@ڑ"/�b��O�Tّ9��6��bX�%��kiȖ%�b}��n��ձz�ܧ�|�5��:�^�������?���� �}�_Z��R�x�>H5#�/{w4�nM��z]�z��[m�nq��So:�ю�}w�769h�Z)2��]�l.�������iɚ~�&����@���@���hw�9[A�8�s&�������g<���;��� �v�@�����K��q���h^��=�H�o��U��w�օEx��LQŠv��h���U�zb�,\X�$_�q��x=P� ���� �v�@꽯@�}�@����=��k���,&.ͩ��\hb��ŧ7x���v��Ɋ�9m=���4�G	�u^נ^�ՠv��h�����Nb��I�@�=��� ��~�Y�u^׾�$z�J?c9�$"�����U�z�����ŕ=x���s�h��f��{^�~}�C��bW��@�<1���N$�I�u^נ_�j��٠�����K��"Cc��T8�d'���`�Y�N�%��cnru��nx4ܼ#��,7[��m�`|��3����6� X*��g	���wb.0���	���Jd�=��e-Í�t���ix�.+�m�������!H0΢�L�$i�e�c�m�c��Y�%���[�N?�i|�m}Z6�,�`hh�E��n��%t"H��Ն����ıհ�a.˺� س��sJMZ�ݛ%�0b���ۇ0�`��1c����̭�"Ŗ&&m4�����2$�>&���v�� �w,�:�k�;�օ�E�D�ԓ$qhol��i4����ڷ�#��V��m��$�h�|M������ ���Eй�1��8M������ ��h���~:ES��!�pP#�@�}�@-�~�&�U�z�������%&Lj@Ǧ-����\�;n�q��.v��X��:�oR�
W#�J�B���9i�����6��h^נU�נw�X����e20����ޏ�Id�t$;�Ab�$T�ccC��&��*��@�����٠}ވJQ&H�R@��^�z�V��G���v�����^	)��>$��/_j��l��i4�����в��F��c�ۋ@;{f�_�I�u^נ^�ՠ���$F%�&@���ù��ɢkW2[�޹�!���j+e�l�8�"R	�&4�M �v�@꽯@�}�@;{f�qQgr�,�!��8M������ ��_v�@��V�)Y'8�
����٦�O�M�JA�+ ����9���>�.�=��z��)q��0��zol�*��^�Wֽ��^��z�a^��'�`ܚ_w+�*�נU�k��٠|�ۓQ1�`�T���6��u��(j�b�ʣ���Tv�0]���Q���b��z_v� ��_v�@�ڞ-��"l��8�
����A�� �������g;�c�E�1�&)�8���h}�=��z]�z��ĜC���I4
���Wֽ������s�fs3x��I�4��.VGI��=��z_v� ����נ~�J�M��&�j5��#6-���(�b�Z���[q)�s�Y�'�t�1ģs�,����������٠}_]��g? ���S�)�f7� Y"M����h}ܯ@��^�Wݯ@��X��RȆE0RM����}k�*����l�>�D%0���$�����
���}����4�ܳ@����A(�Ȟ8�ӏ@��נ[f�_��h]���s/,��Toi��/J)�!kGP�Ru���v�ºN5�h�A���,p&���B�5qf��%��b2�03��'������pB�H]��f�J�/u��7v��Qz��`H^MI�j� d��]�o�{=��\E����զ
,"64g
;Md7���C����#͞�Х�٤�����f�,�]���@rZ������������9u;����&�=<�5"͖'�n����VGy�H���c�&�5!�m[l٬F����Ek$����������4����������=��נ�Ɠ��nM �\�@��@���@>��}��saE�=���0I�$�*��
����bG}}4��zh��%\�"�$�P�@���@>��@/�,�:����IK���`!�=��� �\�@�[^�W{��������iF�����+L��V�X�p٬�/�㝜�ݛE���h��cq������
���������T�d�18ҙ&����*T��H"0T������f>s��D�k�>_Z��r��1#�|<Y��q�98ӏ@��@��@/�,�>Vנw����$rb���Cٙ�U�y��s�@�[^�Wݯ@��U����<�Ǡ�����
��zWmz�3�^��p�5��'�0����WU�����[x�1����.�4cH��E2O�u{�z_v���� �w,�;Gԕs$$2L��
��zWmz~�Y�|��@�
�q��Ld"jG�uvנ��,|̙��s�_ v��rK�a.i)7~��%	L%�%0��rJD���[��p�)��	���|Rp��P��',�����F���B)!:`Rh2�¤,!��Э�(�2 kk�~�<$��B0]��	@<��K| 5��$$FCm�='��K�5e!Ҳ�ہ.�Id����B�>By�)DaIo��| D�ۺoTN KI�0�:!!�+J��B��P&B]0�ȑSx�T�����|��PԚ	6�RxN�x &*��h@t�#�x�"�B����"�x��
	�U��
� <������>���nI��Z�������@/��4���}���������h2c�q��M�mzU�zWmzonM���2ڹ��n��֌O���`�1ve�N�ve�5� \���Sѻ[�:1�y�)ǠU{^���^�[ۓٙ��������;�'��d�nDL�Š[f�9�H=��W�z��h�J�\R)�ɂ�7&�[ۓ@��@��� ��4�X��r7y�4���_j���As;��ǋ�d EEmm�C��o3�ܚ��K�d���@r=�ڴff.�ޟ�=��Wmzϭٍ#����d{mh����� �iO)�-e�rAaةv���������4�ܚWmz��h}Ղ� �Y$��{ro�g3<���y�- ��o�9��$v���3��M̚����k�Z{���H����{��4��-QE���q�^נ�� ��&�Wmz�v0N��$p�0�= ��h��7$���ٹ'��~��<�#,FD
�jHI@!Od�������Csծ�)Π꘶ f���7Tn�Ga�R�n�\A� LX�X�����T��ơ�����All˷�ҕ&<a�����).����)̥f�[���J�щ��0Gx�aa�jF:݇�`�ΞL��媲Țf�[-.u�i��oܶ76�C��h (r^���1�We�[U+��ݣi��ddyDS�!/n5$�����y7;4�	�����4�1�
�m	��4ZAaBa͔�:����Z��E��1'3���&�WmzW����hʱt.F�BO#�&�WmzW����h��4�}IW2A�8��z��h[w4�ܚWmz�u�1�0�|p$���ff.�����_d�:�k�-즁��X"���ґI�@-�ɠuvנ[�M ��4�_lR(8a #qՁ�����"��=x�V[�g�
��-R4�S�C�q��M�����h���s����M���ǩ"kP�kZѬ�f�}�Q��N
��hm���&���^��݌����I�$p���@-�ɧ��U}�{�x�?"��r8D70N&���9��%�_d�<�������f�\:.�8����ɠU�^�~����h�nM �ާpq�'���h�e ��5�M{K�NZ��ts�H]�]�%�.��b��P˼߾�� }m�{ۓ@��@�N�\f@�XȢ����}��s9��z�d�*���/�S}���$w�`�=������@=o�h]�����p�áq!!pI� ! BIHI"F)�!� pU�3��d�������6���L���"Aģ�4=��1W}�{��4�l��ܚ�ǏRA!�E$�n=�e4�l��ܚWmz˽��71�j���.Rz�!�.���Zݎ�k�G^�m+rH�-�#�2�w���l��ܚWmzW���UJ�H���4�ܛ�ffq"��=���@��}��f$��y�������{�@�������ۏ@���W2A�8��z�/?_=�'�w�ܓ����6�|�D"0*a�E*A] �d#YB*T 0\(CEđE�J����ٹ'<�ٯ��\�I)���@;�f�^���>VנU��@�~���X��Ă6�T�F�),��ϡ[�8����C�{ �Hݭ��Dpt�X7\�I���4���}k��٠w�K+M�8�X��4���}k��٠��4״x�$ �#�F��*�נv٧�3�ď[�U����݌��ě�&G�v٠��4�mz�33�}�|�/%�#�0n`�iɠ��4s��s��9$�����'����$�?*�#$���H�?����B�`궲�,�˱nG5-PK��z�Z�[Zln4{T�y�&�g�#`I�OKvPī2�l89Ņg�S�;q�u*b��:9{xʕ��5���nz�^˭P>̽gAaMc&�)�R�V1պ���XG�I�`�s�˲	�1�t�i:�Q�[�4f�:�ZJF˥�%cz��0�*<Q!���1��h�-���\��ؚ#��pK5�ͪfN���I��C��j��JQ\��$�Mh^[pǥ�ۦ=�.�y�Fh�nc�z:{]�"!'�ɓ�yw��^נv����s���_d�=�Яܐs�QG�U��}�s��v��@=o�h.����%���ŀ�8���l��ܚ˶���z�˰�2cȤnI���4�mzW���٠}ޥ����Rb�s&���^�U�z��h��4��y8�s��n{C��r�S�`.g���Xuwi�遖�@�T�J�E�� yc�#�@��� ��4�ܚWmz�v0XXH�4ܙ0�= ��7���>a�Ϲ����&�U�zW���s���<���Ps�'#rh�}�@��@��� ��4�Yׅ�I@�E&M�������l��9��K޾ɠ{����H9Ǔ�r=����l�{rq����8��Y����%DUJ�Wm4Z�C���h�/���(�])Uw0k�EvHY��!�<rD�B&��;�zh��4�����Uڠ}Չeܑ�FNI�7$���p����:�k���@��HQV�'	1E���@��@꽯d� �*�1R�� ;Y����?}ܯ�!����=��� ��honMs39������`�~�G��$H��٠{3���'�<�������Uڀ^��x{%��8�q�9FleJ�v�	��@Z���t(p9 +Y��lM|���4
�k�:�k��f�\�:�)D	�$ɠU�^��{^�^�4��&����$^.���IǓi9�W���^�4��&�Wmz��
^,m�A�!�Z{l���[�}}��ܝPl`hC�>A1'�O-�jĳۑA�'$��@;{rhvנv�ՠ���E�(�v
�1iP������D�-bBm3�-�u�+X����{W��|�~����ڴ����fs���&��}�y�MǒH��ڴ�l��ܚWmz�U0X;�&�s�Z��honM�������*�+Y&p�ɠ��4����ڴ�l��g^�@�L�Wmzk�Z�����&�<6
�����XџZB2�����̬@�V��y�I)qOX洙���e%#il�����kK�5��3ZK���i- �f�N��7��	��ָW��B$P>�$i a`��0SSD
�!�"3�J���`Bd:�������d�a	kBDXE�K���� B�_E��T�5�9䤩,G���1]�6h)!�wv�!��=�B/���FG�����&)�veO�e�V�t��M��	7����p%�I��G�|���w�܉̀�!	*I�bA� �	�����H����6�@����4z���i��\���L���C�<ל�\�osXk����74]�x�`!ŋ}H��1	�����y�����>30�4����� ��RАcČ٥�E[~Y���m��.A[r��
u6��akdG��.\�)K����lS=����| );��⧳���6,K6p� ��Zl5����E Lk+r<�pg5-�<b8Es��5���%W"�56ґ�Q[V�E�;�=���"2�B�B06ԊJL��Q�	`jm�xe��srW%4),�C���/R)�H�`+�cv��a�����ԥ��ۀ��qP�C�ܲ�Pat+e�
H&)L��-H�s��*��1�/e��w�t(�%-���˖�]�����v:����:ǌc��u����K5��˪���Gv�W N'tf��Ά#�U��#!8��;��c���mqڣc;��3{	���9�P�	kTW�����R�����*l��L?��&y�t55�R�.�9���!�i��h��@��l�[�η%�S�nGd�=p�e�6ۅ)K���!)�	���mp��k�U����
�^m�M�]Hzl�;��@�Z;v�`�V݉�a�cۆ��y�@�2�
�^�뛍tj� &�`PfZ6�/P�(�p�XOo>�Gv*��3	k�H![��U++T��m���6�0Ru��Q��SMb'��_k\!c6���Ŭ�+E�gbơ���[N\�G�lv0H�\Tk�>:Ć�N���6n���X�7M �B-�r�Z1��fwt��a^���.ׂ�p��N��6�f;A����n 0:��1�2�LE��SF6˛�h�]��<b���`�9���wny�L�h3
�Y���
Y�a@�c]m ���M��\'mX�}��U�`c����H����T\<�DB�3�cn4dP�	� �e.m��*v8�u�]]/Aq�v���!��f�g�9�h�AU�UԪ��l��ъ��*N֘m��[Uv�#�v��@��m�t��$��3��l%)��g��Y@F&rQe�!t�R�h�6�(��5��^d�Mbu-Y^�B<V�8�Us�l/0�8��Ŭ���\��0���"Zc4um��L ��/AClE(���0D8�@�U�4P��D�*m5�"nnM{��X��e4x��x�<�ܲb�VV[�N땩}��n{��!����yE�ˁΆ�0
6[u�\�݁l�Y����k d:�����p��v1�bY������e��j)MM�e��-CX�#0��R�R���U�-1f(qC[YfM2 �n%� ���H�^�[s	=�3T�gn�Xl%����tר22�r��y���f��8�#}�10-n�����oD��z��q�Y�Lc����9!�l�$'9!'LQ�$��mz�ۓ@궽�z�/9"A���hVנ��4�����s�,�}��VV\�R�go��ɠuvנv�ՠ|�k�>�R�EP�bY�4�mzk�Z˶� ��ɠ~�h�f$�  nL�G�v�S@�vנ�M��^��v�Q���mX��)FF����Ն�Ȯ,r����ݶ���l]>��ާ�b�M���@-�ɠ|�k�-즁�
�<�'�[ۓL���g:@�A��|N�TxjM�ﹰ>�g���^�9����+��R&�<��h^���oe4����I�\G�]��pǓj9�oe4����I��g3����-�T)�,q�>HC@��@-���ڴ�hξ�
19����J�; n��M׫�Xͫ$�r`�yn4nk��I ���lFNI#�@/m&����[�1.�����o��6X�F�%rX�2M ��7ٜ�9�$z�yh_y���7��$}o��1%0HnH9&���ܓ���f�u� ��T� l(�	�V����o'y��ܒ}�}4�uL�G�6I�����^�^�����@�;V��\�,I�L��IǠ��4f.�ޟ��}<hVנ~���i31Ha2ch�1r\l����\D�\!h���ki�	�����Gf*6�My�4�٠_����mz{ۓ@�����E�&(�$��ڴ�k��ܚ�l�?^�K��� ��	ZU���nM �h�j�;�V%�I��dQ�����}�[�O���rO�Ͼ��>RUc�G���s�rN{��]�h�ǉ��@;m��ڴ�k��ܚ~;+�@p�'	JD��FbZ��u�X	W�6m �B6�tt�nf���&$�rA�4�hVנ��4�٠}ީ�yĞ91�"�:��}�fg1#��c��zh^נ~ŗ:�i)�`����
�n= �k՘�$o�q��wgo���y��Z�q�1�m�@�������ܚ����pǓb�M����k�{rhm�@�9��p����?JPZnȑŪ#$��l�zW�[Y-&��azm��׶=�p�D=@&��!�J�03�BѪ�K �H�q��Sq>���gb\a�o�R��p9޵��dj�a�o�C����ɛ*l�d�F���Ge`9�%���������%KR�`�q�v�M(<-�n��s���+�!1r���(g�]�Ʈ�dGq��kG`լpﳺC���N���ʧ�Re���H�bE�Yu5sc�������K�-��z{E��n�W��&�͚��>W�����4�٠U{^�ߺ�,�H�#&"L"q���7��fq~���ޛ�m�{ޜ�I }�4T�ǑEq�nd��zh^נu[^�[ۓ@�{q��(%8�JF9&�U�zU����4=���J�ޚmS܍�O��#�:��@-�ɠ��������\|�� ����ceiP4tvR!�o%�YCFP�9�"�#���b�"x�2G��q���@;m�W��Vנ
u�(ڄ`�QI�@;m�9��~�g*��� ��&�x�o$1�DmI�U�zU�����H���h��Z��)x���8�ԏ@궽 ��&���ZW����K�'��rL"q���4fg2�{��^�zU�������i[+�,�q2iV�ha�C!a!e�6�^{rFۉ4Fغ�=$���ɠv�V�U�zU������_d�>��<ѣ"&!1ɍȴ
�k�:��@-�ɠv�V��z��G�y$�G��mzonM79˅���BDBR��-�B�](�_k>��I����@���Qbx<�#Ĝ����ܚk�h�ա��+��-��~��d`6E&M���_j�;]�@-�ɠ{��I�N4�b#Q��洶&e��9�������ks�:[}/�a�H<�Ȉڒ=�ڴ�j�{rhVנ~�ĥ�<d��Zk�o�3z�&�W��Z�V�on,Kf8�2$��Z�ۓ@궽����ڴ��Lw�"�$���ɡ��s�����/���;]�C����X��B0��9��%��h}h�F�����&G�w�)�v�V�}nY�u[^���|�L�0��g8��*�x,"��݌�YF�BɃ�[͘��	�"�xr[t�%\��/����r�����ڴȹ�X�&H�'"n- �ܳ@궽�v��ڷ���bG���b����G�h{�zz�ZVנ[�h��K�HǐyM�#�;�j�*�� ��Mg39�����>�
{�9�Ldㄎ-�k��nM�~��=�>��I��$�%"�!	!�i<��� 5ĭj5�tP������)q3,,IGB��րR3Y.�桉ol�eN��.�Ac��.Wp��w0�۞�8Nr]YB��rQ�Gݫ�'d9��m�P�8�Q��B�÷]sK��Ґ!hS\�*
�#�)rb�-���$�[�낱��i�{$+��t�gP�����v..��7�����-u�9-��q�g��� 6պ�.��}�I:~�ӻ�|���n�h��Ćl%����n y.���1v80;��痌�mX5u��pW:Y�I�#q� �}rh�V�߬��U����1�<��ӏs&�k�h��h[^�}{rh�h�py���h��h�� ����-v��vb`���&���p�m���ɠZ�Z~���^��H��G�q(���nM�j�;���m���U�
A��2Ƅ0��g2	rRk�te�f<] �t�j���r-5���0�d����vt��� ~��ɠ}��%r��,nI.�������	��D�F ��v�4
�n=�j���G֡Oq'2I��p�C@=�zh+ۏ@�ڴ�e4{q!l�F̂L�nM�{q��V�߬����K����{P
g��$m���=�j�:����� ������ć��Nb�G�N�y�g��A�����\rW=���8�vi�4&�S\I��Y�Ȧ
E��٠�4�ۓ@�ڴ�ى�Ն<RN5$�m���ɠv�V�w�f�~�G\"r(�1'nM ����;s����Lm�Ŋx$|7���K����1q!.� ;
C���>�S�\ٸ�ޮ<P�'(�K%�1)�N�.|)�e����k�͆����.�O8��P�|�sDMK>ѵ�/�� ���榍I���yA��Y�H"(x�BF�	��O%�|�
p s�e%<Ҳ�T���2l��P��[8k�Ff��0l�:"��R�26�>9K ���Tu��/		�!)�C�X
c�s�c�4���Ry�Ν+�%�Y%0$Y�~��k3Z�sY� �w�3��JHb\I�ޓdǧ{{l�k5�W����(A��=��@!u����z*��r$&^h _�wXn0ַ�����Q>�UlP�A'�Ļ	s��'��7u��۴O�H"	 �p����|}����	�P�4�hM��	��|��fE!P�W�Ĕ�'<ѱ���r�H�h6 W�@x+�x*'��B���M �B*'�� ��@�$"�bD�� � �B� H���'���z �Pڂ ���y��ܒy�k`U޷[�bq� �I2h�ՠ�٠��s��sﯲhԕ�D7�YNI"�:���m�@>��4�j�>��O"yE�B2(��q�13��̖݅K� ���3�۶5mO�ͅ0�
5&"rA��v�4�ۓ@�v�%�ѿn�6����U��#��n�}{rh�V�w�f�[l�bE�@(�q�c#qdnd�=��- ��� �٠^ܚ�jy���c�<�@;��@-�h׷&�Ǚ�>�{7�qZ�֡��rTT4P@�v�I�g�.d��CEo�nI��4�ۓ@�ڴ����ެK�7F����j9q�!SE���2#u�&Z�m����2�+Ճt�u���V�NEF�r&��|�h�V����5f,���ݼm��M�*;,�"��Z�վ�s��w�z�{�@���ZQ�	w+C|�#��$ZWֽ �٠^��Z�ՠ~�B��EX��0r-g���_;�Z�ՠv�ՠ[ۂų!2$$�����k�h��h[^�9��f_���acE��e�M�Ede��1J�mu!p��\-�x �14*�
v�#�9�zÂki�u�Ĳ�l`f�q50GX�ܽ��WY���M`S4���u)�Ѯ��[�F�W �u�؄�� �ݡ�M\Wy_^�!m���G���c�<"��K�c��t4�rn]��h<;�h:-���mTe�77�S"�`ұ�	Ka[ڰ���I>I���S��
��B���fR����M*`%cr�bB]rJ�#q0�;L�������8�!���?yh��h[^���qh���IDD1��E�v�ՠUmzk�ŠZ�[��Ďڦ�,X��LmH�/{�@�}��]�@�}�@��vō9#yI�7���qh�V���V�U���z�n"8ڋ��ŠZ�Zk�ZVנZ�qhv�X�ƘN%X���4S11,ލ�W�(@Ûti4@�J�1ԛ�nn�`�L��6�~�w�@���_n-�j�?w�R�G�9&E�Um{���Ԥ@ � ĕ�_�g$�{.��>��I�ϵh��=!2$$����Z�ՠZ�V�U��}V��&Lm(�9�@�ڴ_j�*���h���ũ""&���E�Z�V�U���E�Z�Z�s9������i���Q^��5���6���M5�X�����Rg���±t_�����]��-v��ڴʇlm(���n=�h�]�@����k�;���ڌ�)	�R@�ڴ_j�s=���s�̄h���ب��
Py����{�{��ZQ�	w+BfEr8�_j�m���h�V���ĥ�qG2rL�@-�h�9�Ox_�����_j�;��q<�3[Q��B��#��<�D�y�g8�\kDm��6.)���YtZ�D1�U�}��-�j�-}�@-�h}V���1���5 �]�@��� �٠Z�����=ID�mcQ<�@��� �٠Z��k�hV����ȁ�ɑ'�[l�-v�@���ܞ�@���$�RYH#H��	"ED�g2fr]r��B�Q��(!'"nM�h�]�@��� �٠{3'}���mLM5�F�cG�B��c����z4b	���;if�-�ۀ�ۦiI��O"�_�����
�k�m��33�y���*3�W<Й�A�܎-����f�k�Z�վ�s3>�
{IH��1��{���-v�@�ڴ
�k�-��!�Ԅrh�E�Z�ZW������� LOrF��k�h^נ�4]��?s3g)�8����【�	gq��)g�Ev{$��ּ���%������`=�m��$��g�t=��$�b/k�mcn�E9����̽��/Q�nsV�-�e� ����Y�D&�3)*l���p]�8�c�;]�f�#�q��Ӽr�sܯ��p�"�r���u(	�7�ތ��+,$��Ch]k�Y6�]V#��\��g���� �S�a,�jp�\��k��f���]V�$�;�$�!:I9oψ�L��p�a�Yн֍���kc��(H�͠����4(��q%Q�ҍ`�]˽��m���h�V��k�x���$&A8��f�k�Z�ՠU{^�g�¶
D��Dܚ��h�V�U�zm�@�+�cj9)	�R@�ڴ
�k�m���hF|�R2(27�@��� �٠Z��k�hٜˏ�~F:��0ь�l���֋��3Şı��u�D����c�!� ��U�u�kO�m��~����h�V�U�z��$<�]�䪾��K�^�K��H,�=0C"�����g�]�*��@-�h}P$�Xyq��Z�ZW�����h�׵���B��y�ȴ
�k�m���h�V��k�x���$&A8��f�k�Z�ՠU{^����Oc�˨W��+Apn`�͚�2b�`�E�f��̳۷w�7��b���nM�h�]�@��� �٠w뱸ܓ#�	�R@�ڴ
�k�m���h_.�E���@��� �٧���8g3���sg399��9E�[e4�;�TL�D��$Cr= �٠Z��m��*��@��ć��xDAɄ�h�E�[e4
�k�m��33ݾ_�ɢ6��l��0��C�0�Իv�óv�h�p딅{Q���4F�][kd����zx�*��@-�h�E�}�U�I�6Ǒ�$��U�zm�@�v�@��hu���,2,$�!�Ǡ�4�h�l���{^�g��
МC1!ț�@�v�@���'��~��x�=��X5K(Laf!*���W#�2X�f�ff<�fsv��h�k���p�' �l���{^�[l�;]��	��}���1��!(��
Q����2����2�yv�gtai{8��ҡ��賉��4����f�����s��{ޞ4�űH9�HLnG��7��3/��-���u^נ}m`��� AɄ�h�E�[e4
�k�m��U�� ��$RCٜ��Oyh�Zm�@��-絛��6Ǒ��@���t���גN�:MI=�=��I� U�p W�� ��� V� *�� U�  
���*����DA����@
�P��A`*"��� *H
��"*X
���@X
�Q��
���E
�H��H
�H
�
���@��F��"������A��@��D��@��B"�#�(F�(�
���"���A�"��Ȋ&  *��  U� �� V� *�  _�  ��� W�� *�� U�  
��  ��  ��ъ
�2��:��P))�����9�>���@(����
  %��* QL��� ٞ��:  �)(H�D�%%��G| �@Рh�P ��$ m�4
  6`   ��� �4:�t@ѡ�iZ��� 4x    �S�[  =^ d4���x��1��t� `n0n`X:n�
�d�����| ���v���%���.cB���w0:o��Ao#N�g gc��0t���� �}  t�� ^ eM7��͞mi޽�kU�{��颤�꾲w�W�{z����q�G������@� $�u��
����@(�zލ�� I�;3�7������wx��>�{����Xr�{�w��x�=B� ��� 7�ҕ��z=�Cvn���O��ώ�-���a�;�w@��&װ7a�@ ���zn��B�G@�t<����Z����B�f�G�'��pO@ �!TP H@  ,`H�	:s��� �s�)���ڠW 6Q@�Ҁ���>��)OGtK�o=)6 P{�Ӧ��)�����빦����%�OM.YѠ��F�4ܳ���u�4�'gJP}޹�4��(� =,�:i�  �@  W�� (�K�<�M��@�  w3K����n�k��f�y�� ; Xs=y�  �9���0��ټ�v�Gw�Nv���/��.���� ɽ����қjRUA���hb'�T�Q��T   j���ԪB= 	� mSĪ��A�!���T�5RTi� �ԥ4� h�OQ?���k���?���$�}���~ßJ
����_�(*��AES��*����*��QV�������Є��_�!��#ayBC4l�Ժٞ1����Se��������Sp�-�\�^yk�7���ߡ�ɗ伎��3~�%��)(K��������I�g���dه�<��SV�[q����j�9s/7�}�V��
�Tb/��*���/�Ǽ)n�L��4CZ�%Z˅e.Y��o��,���B$rĖn������·|��/�5���`\5�G�R4�����$(��0�=�pѷ����o��!L!�d燚��˳��{
.�����{����+&s6xÜ�7͐���͐�xl�1�ٜ�͞n��I�˨_3�Ka��2��"@�Y3E�1�a��7|!��M��1�|6����!sD������xh�X��be1!r�I,�q,��M<	f8�_&|�%���L��*B�%͑�����C�jJ��`BR�sD���0 D�8B��X�a�h@��1
!dH$ @��d*FI�!�,cf�9tm�y,���<�s�y�#�����y�P����j���a᳞xp&i6M�u��S))rW,HB���j�.fo^��</����!���Q��g�$W{��J��'�^:�c�W�G_j���5����_o�;u�~�O��U�/��RP����GO���*�wO@����kXK�qˢ\eeIK��m�q�&^y�rsÁ�ٙ�!��_HHoL���	��k���5t͜�W�o3,!�e���g�g}כ�6aV)�|�nGZ��'�W��I�"�������~��MM�6y6���T�$5	�i�
$X�$�$��.0i��J`A�
{�G�;��uE-���y�c�=;t:�tW~O�ڻ�ζ������\;���s�џW�(K����xoTԓ9���G���G��Y���xg���dJF��Z���A��HD���9���k��a�Ӂ/��S���A�i��ϗٵ�,����K}�>c�+�:�uڻ��~�>���
}�[�=e޷�7��o���ˎo����k��" C�ǀp�	�un:�Q۵�J�4�[ܧ��{�<OJHHb�d�oޞ��G��Gæ���������qdV�����:[�����eo�jꨥv��>�;��Ů���U¨*��g���ߧ��ꢹҊ�\�s[�8��!~���OdabUB�.��CB�C��� �����|7|��E��C�<��oz"�7h�٣f�h`W�F��8q�f���m�c�ܻ�h�v��\5M���M;�w���Շ��������l��d Ҙ7�Mɰ�<�u6s'�7��׈z)��9��F�&���hϷ��o7o�8>
�g�_.�n��)��T��&�}���{��0�y�Z���6�SDZ�(Myo�L�Ϗ�q�B\6ũ"�i"VB	R��$�L2n3���Ʃ�$��F�\O��!��=7ϱ�9�L��C66$"FH B-I#r	\a$#! Km�2o��p!��FOvj0��kdʗ�VQ�[%��Wdѻ,�IB0%�B����s|H[ጻ���g�7�2_5���#�xq!#(�D���5�$��
�X����
j#q�H�<!}�����ㇼ�ҳR�����͘z;�T<<ߤ�B���&�}5�������i
cuØS��L SXp�40�țg�d*bD�Z��(0���'�S˯�h�B$����M�)I=�ܳ~a����P�����&��Do�)4os����s���0�B�ϻ��J��
��P�+��<�ۮ
����{�_a�|�1�W���w�Y�U+�}��/=���������s��S5�ߙ������o;,5��[%�%&�i��y�4��]8����M�	�hKй5@�4���4��´]�����_�>}�|��Y�)U[�����w�Q��ݽ�K���ڕ|���Ͼ�_��߾8���Ѕax�$�!�O2�s1�����J��/shX'�F���߹.�h��4�LCK��E``Q��4leq+��J�� l`� 1 �JF��(E�#���$-"%t
�K$R0c�4��9&�Z,B���9|<�=&�|��~��z�R��G	��>�ͤ s�������+��<�Ls1�j� �p����ͅ���>Bg�4@i7k�6`D�6U��]�ү��*�r�ﯮ����wJ�������-����x�K��g���a��F�_.5�x�Cgf=ѿ8G�<�6���٣o�/�<����n���mGTR�]:u����{��=�\�y�>�#���B]��p��l��sq�kd���(B.�0�huй�K�<\���#!�pq�B��s8c�t��w�/����@� l*VWF1�b@4��Ĩ��HK	�����e��D��"������E��SF�Y�uwc�}g��$�s���!x@̹wÚ��u��h��H1��Y]xgʨ���~���9	xa�6s[������ۄ�4]0��;y��n��.�M?�����a�6�`Kt����>By�1�HD0!s˲2�f�&s2�p�C�W���g9��z���h.�%H��u F�?����'����u����3	b]:<�B[!�(a��C�l	c	Yf2��!���q�MH2�aP� P)�B�l�15�\�q��Jbiw!� �U��H{��M���3��=�}�7�y�b�	�@��B���ٛ�ނy�������e�FƄ0�&��^l��u�� ���1�Rg3�y�Ofa���Y��9�~~$OJK��9�7��Cw ͜גi$��IHP��f��2�p�i�%�
KIi�)���0�i��+�
J��$"@�kH��J+�J�/7z��B��6�lW��W��x·2��l��[+��8��4�!���.�\��y���A<�R]��A�p����[3y�{�J]�wl������j�����֮���*��[���Ks��u�����S��.�q��v�����1۽o�)������\�U�U2��ܺf����e}�U������<���SY���u���B1�40�B�S5U�*K6���ai���!�!�4XT�d,���/���jA!�{	���$#	�w���9�owI�q��a��|�y�-�������ny͔���r����J��ĒB���|�35��<X1�)���Է�0��	v5!#��bFX��$+��,.X\�R4�.:�3R�ٲ\���u��f�������*�uҾ��T<��W���o�7Ì��������Jc
��R]�Hp�$�5$I�l!	sz�9�7�4ns�s\&��^\�W�l���{֌Rq;�SZ�j�����B��q���nn]��_5��l���fm���}�L�kgf����}�zf��\�[!5t�83[�zIRT�%V���ė��z3k��s���O	3^�א<�&g���-��)���ܔ����6j�C94d,�S)(ċ��@���5LAa%��H#R,]!s[%eIYR�b��V4 ċH�T����T4m�%x1�x�A��Y�=®͑��%�S�@�I��!9�|�y��g�"`T8�\tR�7	��$�"\IdI�m sM"o9��d�f��y�4I�>�!sI}����t��^4����]i)����Mq�/KM?�6oQ���n�T�2�G o��Bn��{�+|{���q|��盏2Y�]���!)+��.d2x�b�������s䙽���ߎ�8@�@�ɼ��</��]��=hM K�3A�5)�
�cp�4jӫ�މ��q�|}9����1r�7[]�d-!H\e0�T�`����P�!B5�$�!RT��2�J��&$�5q�\	RV\�+cD�4��4P��@��˒D���#\e���%�L��}<��������{{ʡ[/+��������� �7��n�ު�+y�}�����jw�J���陣o�.kcf�&f$,),���>��T����J�(�&]�P��R���.VZ���muRϻ]��ќ����+�B�B��m}�=�����`0٨Зi�)���[��k/5c���҆V���;��Z��+s���s{�͚2��1!���H�\��p�v��Av@���!q�$�%��5J���(�,#!$ FL֍�s������g{2R�N�+ig�gu��(B��Ve��m��i��������2>�l�u�&��@�.kdb��	B�$Hm�8"A( R�&��af:C ��M�u)�������y�l�wO�|�����B%��S�f���֐��2]y�y��:oR�J�)��Pٽ9<�~���a�~�x}�|8����D��a
��D,�h���B�:\ILH��,t�M�%<ɾ�|�4����,�	����8d6��$�����̥�xH���=}��{/X[�����(�}�7���C����0$t�o&m<v�)���p�5�ᴯ�����u�ֻEWԳ��
(y��6�]����yO�4��_?����j�q]�௵x��_�+�8>�]�b�:����%tl��P�D����!�`�6��!��̖�����<���n��Wv�(C�m�]V�/{�]��{�\��I��4���͐�R�e�s����aq��u�$cnY�E4i�3ҳ���ܛ»�}�2BS[��H�����̈́��
�+�<��*�;�[���aT_.������ו|E%��������k+��B�W�_|��y�=xs��G�����W���;=�Nn�f�5�o^s���=��2J�Õ~�_.��gχi�}e>e��ƞ��`H��u��"D �ЈG^���0���Ӛ��O=eϵ�g�a[�:�ZT|������cy]��Fo��Nʶ)�r��.�9Z�6��U_Uܸc����.��ki�m�R]פ�|E�	����qt���[��ڪ�w���;z�ͷ�Y��g�m�0��57ᣌ��y8�Ͼ��yRK�]��+�+ÛER
��¨��:�+)}�p�V<�����������R�%v����n�UmO��c�t�<gi}y>ei�+ee}�����IU}կ����S���߶O�4Wi֫��Rx��[u����Y� *�_�}K>�QO⯋��t�.��sk�G;U|mw�4�f_~.�Q�e:y�hs>>ʓ8D��3죽��}	p���P�����=�{����4�y�k�}&������ޒ�5Ȑ6� [��>�fnh)�ߚ �2��KX�5�D�=rv��m��m��mUUUUUU*�J�UT�UU]T�h1N2<���;i�)�v94�X����T����G�rS�]�T����v9�۲G<�ٶ5K+V.�UY��zO*uc��nݳP�;VX�z��]����[u�������3^�]̆�SNUvx7�_|���N2�/��줻�HPOd��+b�̳�/UV۶�eT�cS�2��
Z�����wc�&Goo(qsJ��u<Qs���i^G3��$��A�gb0���,���۲//>KWhB�Z���m�AT�K��T���}�FS<5�7Cc��d���R�!����!�H�j#h[n�` �kA��ꔂ���n�X��ekX��%m��yZ�vw�9�*�:�+/[U.�j�Ir�ٹ��R�ԨUU/U�J�cSV��½�[s
c)k%�`�z]�'t`E��R�B���V�ѹT=�R��v��9i��ag�m���Uȼ���AKnj��S��(
��^Z�8ڹ3;-�5�ƹ�怱U�nu�h)cXC�+�k�Zn���VmF���շX�N�mW2�l5S�r�6ʭ�����y���6��I�x���	oKaN���K�v)B����8�!s�d�Hq��oB����ղމ���cjղ��v�vuy�;=:���U�K[��1n��^{��G0P�9�;�e\���մ�CU-R��ͻ���.�]�l�@�Ml<f�6��G�n��E�r�[Nt��M��궅�x��N�vڪmF�0�@)<m9J0m=�,�!��e*�U���T�:{HͶ1]m�]������}�����һ��z�x �]�uƺ�q.0�ڪ��,���	����	UWg���U`)V���H]V�j�(]����	
Wh&�G�5"Mk�.��@�JK�j��;�U���X��5U-Eu�:_DU�V]�n�L�n�nBj����K\�,h�Q�]������g�j
��a�����b���s*l-���r��爚��W��2��UT�ŴQ�UKɄ�O,m�]J�u�����n�bpl��]4m��5�ʫq��EJ�G�����\��g��B��4��M�ӫ��*���bvVz��Z�,�M��p �UOq�m�j�!Ǜ<.��,S�Z�"s�䆪U^]���Q��'�� ��K�T�UT�W��mdڭ��{"�wTZ(�U�KUUPUX�*�ܶ�xj9���$�L�\y.V�RR��@�j�ڗ�r�H�-H!t�@mR�7.ĢZ.ń����a�\K@P[]=8���8ڶ��6���Ķ&����ˁ�\�!fs�2�[��Jv�4�5���T[����pձ�@ePD��5�T�*]���T�&iV�8�ki�+�u�J��AUPPqg�U�2[Uv�v�u*�@UJ�.֧��֭G9j]�`KeUUUUUUX�����&��v���*���`Rм�=l����S.͌O$UmV�v��c��ʡ��b���6��
غ�����uU*��*�UR�mV�t��j��LUJ�H@�UU�R�Ԧ5C-��� kf۶��]p2�����UUUb���ή�j�6t=��,��6�.�5*�\��6�	
�U@[c��h��hز��Q���%Ue`*�*��v��� 
���`U��X�AA�U@n�V�ݩ[Qj��P.���*UU����[�"ݡ�US:N�
��,���TӞE]�^f8����cWp�6A�tʵc��d6�����Uڪꪪ�Wm�[TUP���W���ʿUUUT�!l�PUUJ��7[P𭆪����
���٪�
��������T��U�Q���%.��l=HMUUUUUV�P��Vį ��V�]J��W�W��V����yj�U����c�,�{8����ef�b�Y�!+�̪��l�UUP�Km�-yX���UU^��mUuS�ҽ@�e¾"����*ڪ�P8���VU��ꫥX8�	��T��j�gEW\&�Z������A��&��[]TJ�J\�T]]m�yZ�)`:�P�+rPm��j�AAUU1V���m�UG�U,'ʵT����TJ���uVҭb�Ugh�M�|�}y�V�G�%j`*�l�T� u��W0�	���;���0赊�P��U6mʪ�Mh��WRɅ͐��,�)N�v���,��F�����+r��q��c��UU9�8���n8 ��e�yO.�:+h�@1m<p���#�g˴�cY� �X���Kʣ�ǭ�Q7+m�5
�3�یn�������U����ݷZ��j�59Gi��7��K�Q2�c��2�
���%[$j�"^y̕:⮶�M�T��a��n����]�Cds|}�*�T�Խ�Uvt�#l+��6�g��!���P
��1����a -��㥩�N�h0�[�ƍO84�P4l��`(�� U[V�k���`�Q���[��U@�����e\l�"�[��bB�u��K �&3SO$�=�h1J�I�i�e����
P
�(���t�;-R�n��L�و�ۊ�jN8�Z�y�d�-���wf�!�n]�㌦��8��HN�2�m�ѯ[7mV �c{W9�lm�j8�T�� ���v�㞡@��ݏ@xv�����K�(\F�*�Y�+q,�`���ox9ڨ
�*+j(�:6�)ͅu��ѡ�=���Q"�(�Ɨ���Q-)5V�Ե*���[[�����\EUR�pJ�BMͮ6�l�Ϸ)���QAdڮ���f��AW*�|\-���U��W��ݴه$�n�j�y7N��X���kk�݅��7)#��-%.�[U�
�ݨ ӭ��UT��u�%��Ú�ڻm�M@:ۉyG�c+rQm�dr��J������y˃mn%;��6�lD�$UP'x�`;l�` �2*�-\Ͳ���5��j����m�;(�����Bȱ�)���ѵr�kfʑs�$��羧J���g����N�F$�:�Bѫe^�� �X��z��&��Wv��[ת۪U�(F����.���-9�Z������mUm+�o3�,�PUuQnU5q��/�PUUU��Ꝛ�uz/MB���]a�7X�g�����IUv�j�����Z��v�PUUV��W4�QEm*�A�M��6��V|P/UT�3*�M�*�����m��Tu�$G�����jT�j�x�B���֩�6j�e�ln%[��SѺ��s��u*�Y0!�b�` 5�f��(�����A���`�+�A"n:u���(b�ccrM�ǵ����5����c2�v�5�T/2UUI�i|�*��.v`������UVmy���}�)k�c�8`*���}��]�ȻN�c�+�����H_��<�ɐ�D��-u�*���9Ł .^�ں!
���jyeCmV{��(���� /<�F���2�v�Iqz]+W��v�$v+vI�����,v�lQE[R�G��Yx�f9�UY]�j��7`딖�;�m�����J+*�-��NٓO�vC���W��Un�}Utj���r$=r�������A`�	��ԥ-U��S�+���C`�B����ihZ�\�a�d��S�F�ik��n1�ɍ�:^��>�� U�]9����팼V"�핸V�);5UUU,��c����4����UQӲud�n�8�^��X�ڥM��1\�`�Z�P�.��V*���r�w*�UUU[C��g�c��(j�����U[)*��m�7n0t�2��AJ���R�UBGFA��.�Vڠ*��j��کV�e.UڪBjڪ�Ht\��\,UAU�]�AUUUE��A�����a	�m�Z������jꪪ�檺�]���j�����f�mت�5U�%[���V�Ukr����_+�Pm����
���U���������j� 	V����������j���^�қMm�,Ym� ��UK��yWfꪪ��
��T�J@�X�*����U٪�#�UUUT�R�8��J�UU �,�#%�UUi��@Y�Ҧ�gA�v�8��V*�TUUUUVڵV�T�UU��V�U.�UUUUmU�UU+(�[UU�UUUUUUJ�������UU�m� UǕ��7%AK�\�H�An������n����˲�V�]�JD�*��]�SeX
�\�v2R���X�WeZ���cȱ��=���V�vI�㪺�j��T��۪��UUUUU@]T�UUU�V�c�PY-��m\-j�t*�5C��T�UUUJ�UXt��f�Z�(��&*�"0��\[m�ғ+�sf�n�9gJ�H<�j��R�|�UV�J�UUUUUUb��ʺN�j���UUv�"�
��NUAP��R�Uj�Z�V���i:�W��҅��[+�1C1\�N,�WT�L��p*�uKʀ��VݷE�m���IvaP
����Uu��lP�N��b�e�������2�WEV괎6l��m0C �@��	UX�l��N�J8
�S4�l&�Ri�nS�WPF$뭫A���V��k��M�f6&���eh���k�\+ҷ�	�sa�UUU����am�[K�v[mU[5�SQm� R���M��'�3�e�����Tv�W�m����.n�n����ć]�h���ױ����Y�`x��m��b��0�`}���D��)I���v��t4�p�:�_Y~��Om�m�L�&_v�u�x&pCki�J�+:�Qt�zp�-�%հWd;�mA�Uv��iT�#YI�,0�W&��Җ]�<�W��uR���5�!;U*�UUU�YP&��b�l�fI��ELE\�F��B�tD�� ?��?��CHT]� �U6�� DLU�(!��A�*Q(+��E��U�GJh�P8��#�P�M�*�P�$�DB�E�Ev����b�� �j��&RB  �J��> ��D�+�6�|D�Q@�Q}A)� pU��a"����ҧ�򇀈� z"?X�6� |�>�� b(���P7�>	� ��@������H����>P�Q/ʃ�DA|" mPW06���hR��% |@��OP� �f'��N>�3�@��b�!���XAU���  B � HH�B �H�0�0 �$�4P��(�
�d�T���M�裱x>�z�E�P؀q Q�� �OR"$���FD�"FBER!	$BHAI�a#!$	@�$ H��bH���@����C�Av���8|��"�!,"qR�E�hFFHHBV E�	�$V[j���H%��^��1RA`�����@���_L�XĄ@�$7�F�R� � ��RX|����	�zH20brπ=(��B�Dh���s�@� �pEQWj>�tB'�J�b�	4����t:n�������W]�=�K��1���1�-�b��X�0�.�hM�cU�l�X��ɟ>8��v�'\i�sa�T��y�� �0gu�V�5�u��X�¸D\Ķ6/gq5Gm��݂��a:�\Zb��7g�U���d���ݚP��N��T��"(c��^�#�e�ˌ�%1�L�N��b��u��axr���J&�r�:nם��1e�װ�Gu&4-��j:���D�MQK"�U�
*�
�R˓�G$Y�5��Ǘ�]�[���\�Xvչ�x89yx�@nӼ�y�Wn�L���g:�XW͡P�:���k���x줊4��Y<�.:�X���KV���Z�)UVM�[-�:}e�j�uҖm�0������p�H5�4e7&��g[lDn�^8����n9�[PW-G&�7]GF�e]ӆ@wUv�+�@�hؔܗk���#��8�FK�\q��Sk�ޠ*]&��a-�\v����R����F¡�h\pAm�DR����;[0P-�ܠ�+�SKgk=�r���ph�C�v�U"[��͍����8�`χ��6vr1/��t�N@[j��8���T��<�-�<q�r��m[�D�Ÿ�K�Blj������.�p'��h�<���v��X�&�֔wN^�sʖ��m���v-�bF[��wmqA��U�z5��;kg�^[��.�Vd�5���L�s{m�8�����.����Z���2e��<8]� �a^S�mȼu�n�Gy�s��j4���t�)Sΰ��3�+��Um��J�4m����$%	M�=j���Xvj���1�^A�i�NM�b���`�G���6i�-d��흲�v66:#�sr�P�UZ�PT�)��.Yt�[x��\��d��e!ԩ���N�����t��-�����+�p%���oPۡ�%Z���ful���e؂����Ln��d�)����g'Z%�����2�\�됅�R�k�2,������6�f�F�&��f�蹖\Ъ�� �M�@t��� �9�����|��B (�X�˓17���P͠��:C����q؜{q̠��l�Ej;"��+�ۮy�d�f��j��:�T�v1���� �Y1�Ћ��sKCwD���`�6ےv��6��hd�a\[�m�-��9kb�@�7a�c�N��5�����<��]�s��;%jZ�r�e�p��e�^�Z���V�z��޻�@z��ϹW�P6	�jz����� `��pyN������\`��v㲯p8��W6+���庘{�����9ϐn�e`�/ ���vӾ+I� �엀�<��+ ��D��t�]$��&��� n���L��8`]��	�L�������ն��L��8`]��vG�od�V��n�:M�� ��6^ n���X���ԓ��K�*���X���ne,d5�ڌ@�J��9�v�m�6nő(�<��!�'m��������ɕ�v\� 6j�V�]��N��[w��<��s��B @��R��E��ZR�k�YIH1�ihŃ�d}E��Q}�o~�ܓ�3��un������BV�&�[M�{&V��X{���zz�{�x]����IQlNݡ۬eȰ��x$� �ɕ�%(�;j�Ӷ����I��+ ��X�\^�'<�*IkN�i��"�Iu�ɛAj�M�14-.��F�0�MiXj0��+w���<{&V%Ȱ���	�&���v�Ӷ���+ ��XT�x$�=\�7}�*�Jڶ�O��kZ7$�s���y~�����'+�*�]��ɓ�vl��>ۓ��c�Չ	�k �ݗ�dx�&V6�X�T�mR���N��[w�dx�&V6�XV����tӪ+I���s�#5ht�R[���ggL@��f�8ĽLѭ��쨌p�Zf
�e~���r�	�"�:�e��e���T[�hv� �r,�\�H�'� ==�od��	�D
���w�i�XT�x6G��ʤ���X��� ݒ�YWI���MZ�x6G�ove`O�Ͼ��>���E 16�(�U�2�^��vUv;J�i����+ �r,�l� �#��.�O�佗h/gu]ezzm��{3��iMIc#�c�N8X� x,ᆒw3W|ۑ`Se�d� �d��>�'�-ݵhHm� �ݗ��<�ٕ�n܋ 6E)�ʻ��e:ujۼ ��n̬v�X�v^ l4���ċ`ۧi����r���{��$�y`-�xݑ�v]�R�IQn�n�M�ݎ�]�= l�����������ҕcQ�e�:�#-`�n�c���!&�ݺY�n�ѥXN//8�;Lc��m��q������7NG��Ȗ���
���Z�m���sW����<Fs��xp�ƪ$�Y	��ێ���K�F���]���uJW�K��U�B:y��<���P<�'k�1T �P�4q&��p;x�W�NE��	�r;��5�np�6�[�&�9v��;��ӧ���$3�b���GF'lʹ��uc���[r�4o�ٯ*u���06�ק��Ӷ���׀���+ �܋ ݐ�eПI�V� ;�<�ʪ�H��e`#�uM��N�vUv;J�j�od��;�2��������KI�n�ݕn�u���^��������G�od��>����o��Ё�� �/ >���+ ����=��Uv@G��B�l`��AB� �<x�r�vyk���:vA#�1�מ�4��]�l��շ v{� �ve`ݙ^�W+�d��	����;�Al�r�Ͽy<�>�ޝ�яB��#M.F"B$IIFI
�9��b�ԁ	5CD��1���> �v >�3=�f䓞}�l� �����ݥE�J��m��ٕ�nǀl� �����$N;i_Vف��9UT�}<�o���̬�\0셣*�:���Rwj��� �ɕ�vk� vlx��~?T�Tx�w1MAq]^�Ŕ���wt�e+���(�O��ۧHm*���ٕ�vk� }6< ����e%�j�m�۫-ݷXf�`�c�� ����>���Wm�ؘ jـM� 7�<*�|9UT��\�\�v�9�s1\̬�$Q�m+.��bUi����ٕ�vk� }6< �B剪��ۦ���7�e`��� odx�:�����T�Qt5��dn��L0S��-ϣm������p�)*���j��aY�߾�� ��x���l�X�(	DS�6+�m������9I�y�}��\3�H��-`�ZIЩ;�m��y�ݙXf�`�c�'c�*�)���	��x�fV�\0���ܜ_!��/��(?C�7�<vJIe*nۻ�V[�n���{��R履��� ����7nQI~N��6�䥱�E����@�N5nk[Xɂ^.��G�q�!��-�rx���fǀ}�2���`ȣ*�V]4�*���	6<�ٕ�I{ }� IP�bj��ݤ�Yv��ٕ�I{ }6< �c�"캔�HWV�%mU�u�I{ }6< �c�>ݙX �%N�د��m`۱������$�� uU_�;�����q|�]��^yMM���;\�3�e�iY�׮� n��� ۵$Nh2���U��)����k1��;ǅ9&0g	m�G��������F]�e�D�0�k��LV�ط����J�M��b�6�GcWccG2�wt�^�]h(j�KMV�3C��1�[�����:p����8x؅�m��˻6F��Ӡ���Kr���Ӽ�$���&���M�x�u�@nt�gZ��JK���z�e1���� ��Ql�j8+�c-��շ�vy�ݙX��`�c�'c�*�V��T����7�2�	/b��ǀlx{���[�ݺv�ݷX��`�c�	6<{�+ ��aV�ݰn�C�����ǀlx�L�KذMQ�m]��v�ӻo $���X��`fǍ����ȥ�lv�P�-��V������}�4U�:��\�a5n�)�05Jؚ��hf�n��o �ɕ�I{ vl��U�flm����o�=���(Ievզ^şo
�s���������< ���ٕ�ĥ&�&�|M�m`۱������$�� ���Yi&��:�Iݫo $���fV%�X��x�N�_%2ӵJ���{�+ �{ }6< �H�UUUw��k�q2��d�`�u��m���9�֐��*]���KP��=��	���en�K�X���vG�}�2��L*�Zmب|�X��y�W) ��� �=��M��=�s���q�U�1*v1�o =���7�2�ڹEp��#HC�T��0���@��.��4����H� �H�2,� d�BSH�>Y	�e�'�x��"E5_�[�I�vː7�����C�͆Pq B@� �`�)�4�) ��`�5�.f$����c���׾��ą����w�<<<]A������̄&c,!����5�qאp\I�O5������\-����m�kjJd)	�C��P�G)�L��Ȭ&h�m	x�p�8\&V����͙�D�raߴc6��/���7݋�n�ޞ�B�@�o�K�e��˜[�ܹ�����捔��Ia@"<�➸����p_@�D^ @]"z	 ��@�@�,�DS�P�A�V*!����)<�<Ͼ��r��ٹJ����t[�����ove`ob�>Se�z��I{}�yo��V�h��һv��`ob�>[���#�>�wKM���vw%vH"����B*��	�7lZ�G�yd�Gi�f�9Tg���ͧ�!1U��M��/ >�<{�+��+�\��&�֒���Z�V�5j���G�}�e`��`[���\�${|���y�n�Iݻo �����ذ��x�����K-+Vݵt�[��`��`Se��G��ꪪU|�
���a*��'P������$��n��T>��l��RK�7�2��рoV�t���k�9�8���A�;Z8��!�lݱ���i.������+"�֭Uȝ���Ͷ�{�x�fV�{�/ $�Z�I�Н��Jշ�ove`��`)��vG�E�u*���զ�ۺm��&�ŀ|����<wfV M%�Zbl�)����$� ���ݙX�ذ	�-%Y`Պ�%I�V� 'dx�fV6�,�6^���%``�̕Ąp�-�̿N�)rC�ۚ�f��z��5�F7TN8K�,nP�ێ�d�G�bո���wYen!W���v���f�\4�b�CM��R4,�F�F1�m���	���X��jСu*F�����u�&@��!Msq<(OJv��^��A��*�w�q��7Z6陉 ��I��	�9i	���H2�:�r��2�%�5f5��1�e��ùw���]f�afe�����u��ɜ���u��a}�*����5L&!���Y�%�pʒ���ET�`�u�m�DYl�������&��/ 'dx{����v�Z�v�ݷX�p�>Qlx;#�'ve`l�U�,n�b��jـ|���vG�N���&� I.S�V0E��i��lxݙX��|����(�Tݤ'n����Mٕ�~�s����x��/y������h�'Kb���L��6a����u�c�h0�wa���5�[2�ٰd��t�u�I��) I����Ur���� ���yZV�X��l�>Z�yڮVs�[\����0#�x�L������f`?sހ-F�T�R� =��vl��$��G�NĚ��
m�����xf̬Mp�>Z�x����%%J��iZ�Yi�u�l��G�j�/ �ٕ�z�9�I= -�ȫ�X��Dܮ��%�qځcj�ZR`M�-�W67bȵ����k�Vπ��x���͙X�p���[O��4*.�V�x���	�2���|����(�Ul,�n�V� ��+ ٮ|R�U�u�r��,J��WH@H�20%W%W9]���W/jG��<V˻D��J�4���m��\0�R< ٱ�R���� ��.�`;e�I�m�����7������2��t�g��zm�Zl�s�xWl`x�9݋�c�7H���<93�Mn�W��C�v��Rj�m������Xd�^�W�:�{� ��My'e	�)Rv6��ɕ�������߲�Q~��d�=ʤ��I$�!��e�շX����}-l�=�RD���l�V�d���T�m!��;u����x��x�̬uCD��
#�� �	�;�;��_���vӫ�i�� wdx�\�l���=��ke縑����?!g�l9��ws��8�����=��Rhچъ;D�W2�� ڙ��q��gI<|���[�%m�������-��V�Z��s�������<)���t�U�Eۺ��`z������;����o�w����ݛ�*A=�]z�v+uvRRǙ_�jz�R��?��s�Uʻ���V=��W��	'�Ҭ�h�:&�M�ܤ�{�>�Gw���6{�X{��r���{1{����'�ПnʺN����R���V�����~��߲��nI=�ﵹ"�I,�,$ ��ߟѦ[�aT0���&��jذKڶ<���1]�����Fc$�S�Xީ��'�ثؑ7��q��$ȋu����gr<�{&J����ۣJct��-�LT*��5�>[X�_�/���,��k]������ӌ�*����.��Y�����+	�nc^%��;����"�X6�Kg���-�#���j��
K��Aaxq�9�ǇZ�Ι�;{��t9�o0�o�2���K�Rђe�L���K*[�{9z�k�^+���󻕸0��e����6��O�X�������~�|���e}_ ��ظYj�m��Ui۬�jz�Կ���{��o�~��;$����H$���o�m:�am�M� I�<wfV�R[�{+ �O^ nօ�*�m��������W�����O߿e`m�����R{� �z����V˫�v6� �+ �cS�����>�2���t}҅%�бQH�GP�ӓK�*s�n���;6���7]��l2r�FL�����v���vG�}6e`�� ��J��tZuj�E�� 7dy��,�HBBU� �%+XGT����!D4}c�U{�Tꪪ��}��{u��>�[/ ��V�Hv�I�M��ɕ�vG���x�#�>씐 �e����6� �ݵ��d� �l��>ݘ�ucl�v�Zm��ke��W����{+ �0�Г�!��kwL&v�����<���+fHm�Oj\W3�Ur'e��n� ��٦��{۠&���6G�jK���;TS�T�����n̬H�}-Ix$� ձ]Z%&��uv�n�	&���s�}����0B�Q �\���Uu\l�#�;$���U԰h.ݎ��v��jK�	$xݙX�� ٲ�*ʺj�Z��i��	$xݙX�� �Z�����CEZ�h�i[M01�a��7�/,��7��H�J�,�N��s�<AI�R��ĳ_7fV$p�>��� �G�}�)!*1�n��ջm�$p�;-Ix$� �&V��`�)�Z�J�6��ԗ�H��*�����{�� I���;Wt�l����y�����>��}7' �F
�<���ϽՀj�h��m��ҷx�2���9����~:�_�� �Ix�j�VK(5�xI-R�V����M��՛��1GQ!EFR㶌~IMh��&U�GT�u����ar,)%��_ ��� ��y��av��!�v�ar,�s���/{׀I�e`G�W*�$���e]�N�Rh.��<��^��+Ur�/{���\��6D�Z���j�t�۶�?s����s�~��v�߿?�4���\K�����P� ��wn��X�� ��r�����{���߿<��4�#�w|R�,%����B	%%�ID�� �2r7E��!aD"BF�B�����>�"����Y�I�!#1��xL� 2WVg�ӹ���;m���t%�Ė\%1!q����%�K��#.$����y���Q�𔕗-��+�0&Jc�^y9� ��8��}=��{R�u�U�=��7�d���$!#ZXIHA���P(V4%H�H��.�������HHHIGl�2�=�|׺�5�Y��f�k�]���KZ%B�eˁEbA�1�Ē>o�U52��j�i��"��,H�A+�,��J��"RHI����B$�F`a�$�CL���Y5e�xSߞ-����� ��l����L�2��\!�*a�)|��p%��Ȇ�k)+�;e9�Hz0����M�u���Y��T�R��c)��	�.��T�&.��$��mU\����&7���������\a�r;m9m=d��p��fg �f��8cd�s:NzĈ�7>]�g�������nF훥d�	�Cև*yj8���ي�%��w��曨ҍ�-�u���p���t��v�ZH�n�Vk���BH��m6<O-�!�����c+��`+g�9-� ��f��@l�\��b�]�-�v�Ԑ�k���J+(kmƹ�g��q�ۛ��a���k���g�島6-��n�E�:*�[dTr%ɠ��qB��qv��X��PQ��9��t�Q����9�jڱ��m�n*�r�"��;�wIcn���۩Gu�RU]��e��SF{p�MLk��X�jj]�
�D�-]&��2�B�t]o
``ݐU3c&�ՙwj�6�VҜ}�ֳ����2��!�k�`�J�-�7�Q8��X38�q��v�n�ms֍�T�R�#�C�q��f�����
��p�u���F7�՗���֞�9��d�sta�[e8��Z�#	sEؖ��wظ��0!��v�3�"�g��<�lf�KiD�C���MQE[T���-��5��R]��J�s�㛥Ñ3��,�>َu��ֽL��v��^�3�,�gBa���`�6 }b�'\�!�����c�ƅ8�V	��;v.�s�l�c�\�O[�˛F�Dp�Om1����I�u��ҥ�&ՍA-�)T'�<� )��As�Xܺ�F��N��X�����u��5lFr�6h � �]���m�OM����݂�MJfmض��zqͭ�e��ٶ�P�gh�VOR�D��*K�	ӓj�)jJ�z+&�L�r��Jk��6�.śca��ڤꥪ���$��bZY�skrX;jΎl�m�2�p�8s�yq��<r�(��K��xÜ�]� Ր���M����y�ǵl�A׷L���ɇ�́�l\�
�g��8�V8 ��Ckn�l"a�BQ�<b��0Y\�n)H�%vkl�g�FDvR�-�̗5�b�'��Ut �P�!� � �|~���(�������J��5�ȷjpX�<%�iʈ,n�esvƽOm������{.�"buq�:2�&�gvu�W,�-�#N��*�m�sp�<�Q�c���5љ����d�2�r荽m�aEIP�=�����.�k��]��6٬���B�,�͹������K 6�v�p�6����	���+F^�xۀ@K�nSť�,�ns���3���qm���[uI�L�,�� ��'9����&��'R�[::�n5gn^A�,�ù{p���vC��_$�����.�c]���~�/�� I#�>�2�\��{�~0}-z��]4��$�-��H��T�����=�?�r,�W	*��&�[b�-[x�{+ �8a�ʪ��U߼O�4�}���|����*�VE,�ܪ����� ��y`�<W+�}�}X!��$�[��;n��r,ܪ�^���}�e`I��M�K+�\<3p!���	�Z��E-n�h�*��K���XapC��f=kR4iEEETG
��{�xd�X�e~�U~�s�ֿ~�߿%�-S�[�L�N��xd�Y|Ca E "�!��F	����)��?~ٹ'����nI�����32G���bc�)-�i���}��;���=��)//{ך�G�짉$��Sbc��+���e[��Jw�Z�h{��s�����l��������ޜ�>��ʺ���Ƃ�塠 �;۽�{H���v {����λz ����L�YE�"-�Z慹ɜ��'lh�L��kc��d9��c+��wM�yGS6+����RH����$��>��I-�q_ʫ�@�Z�����\������0�qKT��] �{���,JHwԾ��$�=���$l�O=�r���[W��&��;Kj��=�_C@�w�{9�ڭ: ���{ݙ�m�{�xs��=�֬qtT�����bY�>Ė+o;����m���fn�o���r���C]��n�s��7�IUqB۽�>r�RI}UR��F��w�%��,I$��� 'SQvQQ�!Z���c�F9�j�7<C�4V�uu�dʐ�GTy�Γ�<��]�fK"�Il���^{�x��h 7���g�����@�y{bc��+���%{�x��k�$��~�w����@�s]{ߖd�9;Z6ⰱ����X�Iv{��I-��%��U���{ �]� z�Ґc�	k"��o`}�|�J��}n���mo`㷥ݷ�bBDvJA8#���ľX����}7� ���V:�+�Z�;m�I%���}�Iz�U�C3�|�Iv{�{ s�� ����I#��r�,m�,lc���g�nBӣT!c�Z��F�Y�UlV�,Ņ�Қ��'%�m�[W�����$��#��Kv7�r��]��O}_|�F��4䎊��'F塠 �;۽��,�,���}n���mo`㷡�,X���x�ܒUEE��w� �}^$����}��+�Ww ��ĒK����$��z�=Yb	,�W%��b̓��/�I)�F$�_I�$�U�]��7�$����]��]�CM��$���#A����b�Ͼ���}n�s����5�I&�s��0?I?��e��e��)�X�wj3s��u�#t�!mӀ�;��q ǅ�@,�lplj���K��ۍ6�#��-�I*�B@tS�=��l��竭��n�	t�k��nҊM�6T-�tx��xĄ���=�\�5Ŕt�nka���2��^���z�;�����J)B�޶���)-@CmA��ۇBU:���,�c�`J�P
����wtw��d���0����6Z�gr�s���N����^#Qc���|���!h{�����;-�F����������;f�ݟW�\���R،I$�������R�D�-��ӝ�_�I�ﶷ���hz ����ؒ����U*�W���۫ĒRO}_|�[���K��*��}�]��}�4 ��Q'%�m�6��^�r�3�#I.��|�][2�=�I��ߖ� ��H�䎡P�N�ɫ7m����9m���k��3�m��qo`��� �S���%Q�'6 �3�Pu���SG����I�ÄGMR8}�� �JK]Q��Yo��;�)�wg���%�9��W>�I.��|�Z��F9e�$�)IeS@9��ofb��1~^��5�]rk��v�o����-����3�X���9��m�D�[Z�&�-{��?،I%��/\��S�W�$����rr�Z7] r�J=�'��z��$�Oe^$��{�$�Uʹ��� ���:�� ��(�����LI%��/�I-��F$�����%�"X��lH��ċ*�L�(�k&���ގc�����X]	�e�wq��y���M2շv���JG<��$�G1�K�_���w��6{)�I%!�X't]��Qm��8��k�JH��齀>w�W@9y�{�f,� ��H֣��P�N��C@��zo`�;�t��Y�
 T�� 8��<�y��y�z��h ����A�"��7�KܮW9V����$��y}�IM�bK�ؒI[�}��{ ���Q�ZW$�R�eW@9y�{ �X�=׭x6 ~���� ���] ,��ےȶ�i�nc����M-���>�a��1�mq��	��v�!�I%x���TF;e?~ �]� \���$�ٔ�r�U_]��s��K�����tl%�4 �{w�fb�-{)�I)��䒚7�ܪ��UU6����êW�"$��`��J�]ױ}��+�w~�~KI.�y��I%c�nU\R�(Z���b���|o`^�k]�v�o=��s�� ����C�z�?no�W@�>��+r[P��i��JB�$�_l��H�2�$���m�'wwM�~��l���Õ�r7 g�ϧwX�ܠ�-�����#X
GQ��-�؞W
�c�N��Y� 9ﾻ��;�t�K��/r���Iz،I%��K�r�pd-���;�u��R@�o|oi%�{01$�ײ^~����*����E��wwm:�m�x����&�ea�q.��^ I�<�U��M�H����=\�/C����{׀�<v�,w\���*�Ī�u�|���{�����	.y`I2��A�9\(���j@�tvPq�2�TV�
T,�f��w��.�:��n2ց����q���Wj��7��S\��<T�.ݭq�k������Ʋ��d��j��J#��R�:��ɶ���a��������V�p�m�����6�����k�c����ˊ���gkN� �:���NXFx�q.0�vZ���6�ڌ=�R�\�u�l���p��O{���t>���X�r�,�D �m���xy��tb�-�+�m�\��nnU����_w����~ �{��7ob�&�ez���T�� �����ݴ�V�[N��;��g��T��{�XT�� ;�<��$Y�L-�ut&�� ������x~�9T���x��`d�历!ҡ��u��r��۞��g���`~��s��K'�������>�UDJP�
����G�{��9Ųy���V�܋ ����/鳊m�na5Y����n�y��B�<n1I�άHsX��h볙$X�jݻ��ǀn�2��8z�\���7ny`�~�*�Lv0Uj��xzI�gʇ␨z#�H{IM���U���P�Il-����
�%��T�� O�<��7$���, �����*��$o����N���AsY34nI�{���<�=��~ ��!˳���H~���T#�;BI]���V���� 7v<�$���W*��qv{<`��%wn�6+��+m� ��x���r��O{���?{{��}҅%��QQH����tu�q.���4A�������"��*D)�r�IbX���Ԍ��n��M6�t�����X{{�����@l�x�.��Wn�J�*�X�r,��� ;�ޒeg��~��1H�����V�0���m���]�'����4��<k/�`@@�YJB,�!m�� e1�����hu$�5׍=�xf3��2*I�Ef��1$`�h%�k\��Z%��
��JBaq%s(B"�Vf%RM�"H�O�so��$�RY�2i�0I�HB)0W{1ѻ�����\��f�I��6^�`���eՈZJed�0� 8D�R�A��2!$x"s|�3�	N��H��q�KK�<`xQ&���c �9�r1	�a� �������p4Ofr�p�a45��"A�#`D��kD�E�Ag!B)X��GaD�E�FBC����K	���p��<5�>�m��+i"@��)
FK`Y@�!�"��� �������C�|�D4�x�qAе ����><@؁ל�U}��w+ ݹ�uIP-[n�Vӫb����W*��<��{+ �I/ ���`H�QM���
�i�xzl��=U��;~���7ny`�ǀE�_��Am�����c�m�qc��[��`s=-�qŬ[��,�]tCv��ӧ>y��1E+v+u�^�� �ob�ݏ�9\��Ė~���ﴴ�|�Oꨪ "�)� �ob�ݏ �I2������Uq#�޻�J��t��k $�xzI���W9U��\�]�����_�, ��ߦ��3VhX�|d�t�~���xT�� �ob��\�r��{'� ;6��[���J��[��^�W9ʭ�<� �<��ٕ�~�������tݳn\E�$��an4�q���7���ϕ�^�5�B�ϱf,Nh549-��
�,��e���ݏ �I2�\����w�~0Sǀ�n��m;����ޒe`H�M��9\�$w�~�j�v1"�۶������p��U\��#�O<��-1�tN�![�[��\��UUU{��ߌ������BL�)R���	$��]ZV�n�`��_�\������7���V���+G9��Ғ��QYl����!�H:Zщ
�i��b;my�*�n�e6ae�q�\���Nr+�C���A�ܱ�P�:ݶ���2���ɞ�'�ë�-�Y�ۜ�b�`9�ݮ�r�7=�b�׉�"��9N��n^�W�R�p����W1����ʙz`�a���z�0�v��:P���Kl�<����ⷴ���k��_q��Ozw�|�FwN�|����@ʹ�0��xl�q��â^�\�Ol����I9׮��&�߾��?}<�ٻt6��t�ݺ�w���>��X�r,n̬ ݩr��[�ڶ]
�m�BL��9�$uOz���V wv<�r� ��~��$�]*n���^ٳ+�W�s�vO{��7���X�JcC��E�M$���2����i&V���n{׀j�<��X��c�`wc�=�Uv���S޼l�X7�����J�H'B#��$�K�ٝr��.�����j���g�S�&������*��xa&V��/ ��+��|��<�Se>N�!۲���^YE����\W���?~��V n���>��XR�(5WI$����n�	�2�vG��\K�=�W���>R\C��N�ں�&]���{�������{�Xv�a+�K�gՀ���]Zlv�eЩ�o �I2���vl��� }�m�v�/�5E��ͥVmW]rs��tu�P0FY����.���Qo�:>m�Q�5&������xf̬ ݑ���|�����O%�i���uhM[0͙X�#�>�L��8g��RF���;�J�m;&�rI���$��nT���$!0Đ!#�Q�E���b@��C����~0����'H�14���Ъ�����+ �d�X�r�)=�n��Uo���t����XeȰs���{�W�{� �e`ov��M�Ҵ�i��-j�FU".U*<a���ylo�Ϊ�R2��Q�P,a)�����Zl7dxt�+�s����Wl'���`�~��ut�v��&����z��W6�V��y`�e`v�ʺ��i�N�*j��;��Xdp���r�Io�� ��x�]�!�E����X��{���=�{�rI�}��m�	@�*���r��gՀ}�'r������&��`I2�W9\�R{��6�Xv8`��[LI[�ӡ��m�^� �R%�!ƙ�%#��f�hM	J��pc�;����e���`���=�wM�Xv�_�\�}�e`�{+j�+h�i���+=ʪ�ܮr����׀o�߲�vG������s�vI��Տ��`�;�
�`~�����X����fV IR��1�I&�%b��=\�8��{��	'��6e`{���]����޿!:j�[��LM&� ���ܮV�{�$�w��ܓ�����Aq	�T��@��X�0	R
P��	�;U��*蝐%�JX�l3CM��T���4+�%ȲS���un������;�2�9NܔH�Ӷ���S7d�N��Z�����(�hjP(Xf\�+�R��yi���[	Iuv����N [vtZ�c[)�r�*�{v��h�4ٹu��`�L���#c�,���N*���ê��N��}���u��Y�\�y��]�X�!�5�>�����N��05���8GR�괔�u�=��>)�m�s!�r�:�Xq�C���������y���wISM��=�+ �G����d��$Ӣ�J������s����?$��7M�Y�UU${|�v���:�W`�jـw�~0wc�;�̬�r, �aT�e���`�0=ʮRRO<d^��>RK���"���w��䟾���asWsVK�-;o ��X�d��������V;�k�� �U*)e���4�,!S4x6����j=�����.^-���{��~�^�۰���bV�o���}5� ;��9ř�bK�o�����o���� �335w$���齠�z��]jOu�x�)��}�"�UUq"/z�z�Ӻv;��&�f l�xwT���q.����G� 7j\��m��t�x��UKd^���?�\0=��q-�� '�w^M��-0�n��p�?r����g��$�xwS� vD�����eL�Z�딄w0���X	V��c���`Q�hDv�6�;��?!��:�˂г�;��`�ǀwu8`H�M����Ҵݻ6� ����UUI"~0������s�T��'��&��+h.Ӷ��?�8a\8s�AVB FB@����da$F1QH�� ��8{����W9�c~0�<��\[F!�M�[���$�K��zx����ݏ ��p�"�*Yiۤ��J�m`Kذr������6D�`K�`i�	ڴ�E�+i'�j��&I�͸�6���n�.֚�ms��Q_d�!�dcN즋�M�n���O<�k����Xݩr��n�eӺJ�m��fV~����ʮW.����0��, ���v]�V�t�`]��>�� �I/s��9ĉ'�����'z �Y"��#
�+�~IbK���Ԓ}����{=�f��+��P�SWc�`f��RM�jݴ0�� n�x��9��\�W9<{�k�o���}.CM�~�����Ej�8A1���9�� ����(��@z��;���rb�l�x�\�&]�m��fV���^�+�\��$��7c�V:aB��vX�7X�8g����q#��y`�� �2��Ē����;J��-��)���Oy`��a��ʮU%����;����%�R�vĮ�ۡ��x�`�fV���\�9K�~�����][m4˧t�NـwM�X��X�Ix��z��6�B���BB@��@�aH@�@כ�H����VG�!p���<w4R������ń��w�BHM!,�%���p�b�%f�xM�b���Kr�8Kt��BT8��$4f�0�c��c ���XȄX20�Iag�,7	��u$Hh��8�d4ZRe)u�8+ͧ �J[$!.��)��6��[�9l!lJ�f��<�o�j�aT��I)�A	%rCK#B3Z�a	!	 @pq8�8�!�BN����PUY�㪮�e�m�1�B���N�����7�DnFݖ���r�c8�G��DkY����'�l��3�W6�97���d�w���D;\�5�	�w�ôXȎjF���60s8��B���,r�P��u��� �3i�(a�^��s�;�3���d���Me�:SM�n0�u��`W:�f.uV�7gi�u�d ���*<6�qK	�j��q��{KXy6��	u��T�2�]����`x;Z7W�qrlϷ/YA1l�km.�Jn7�`��"j�����m��2r�9�t��<�k��1���@:�3��+�����%M�Z
f�m�u��5 ��5*��"�q5.��m�ih6-�`��U�rl5]���u��M�t�����v.Cv@U�Z���((g�i�p<�������T�M����ؘ�����u�Al�m]f���&����c)��WX3]2�tR���ⴂpq6�TT��Y��n��sɲ�ny�ƶTt(,%fm�7%!�H�۲���LM�-[����l<Whgh�@}�6yp�Z��=9�`�']d�1�.���\hшѴ�����W��ǡ݂�#��v�ݙR1�d����Xb��m�6Q�n,�&��j_ntfs��s�F':pDp�^ݭ�t��<K�ێ���#�2`PM��kk�Aջ;���b��uQ�a��.P�jK47[�8��к��4ڕ �V)ח�(��K��k�[�8d�CK�--�Gj�U����4-�m�ٞB1��4"e�&tW�UU,N�M� %n�1C�H�5�$����JV�FM��d������eP.p���-u��)�7[V�X0��[F����l�NP8X��\OY,�IE��72��6秜���4X��0�X)����W�m��`���T ��x��&���I�i6�9%5T��*X��p�oI�s@a�6���h^.s����ɢ,)�v���XF� v�/5،絃�d63�5`���-����!'AV�p�}�DP�B����"�;��z"?qЀ/��*hB�x��Oa-�rsSVX�����I:�G0n�a`�u�Ta(��+�C��j7=\�uؕˇ���M`�n��:���m��Cf���L�k�qp�=_
��'�u1Ūom��p�D�p�!��em��� Ks�'M�v8��"�d�t/:���=�C-��s���ۻa.�#�n�؉�1�K%=Θ5�e��W;"w[q���'Y;z�r���c�K�\7�wI�����
m�e0W-�c8����<���;��%�h�
�$u�8�g8�;�(UmAh��v��s� �I/ ��r�ʯ�l'��o�H�!X���ؘ�f�^��+ �2��p���+�s�Uv��]~E��c-7x���Xtٕ�}#��^��eZ��MP�պ��W+�a=�`����$�s����V�?Zm�
��b&� �\� �l��n���7M�X۴�,��J�-X���^Ǜu�y/ۦ7e��]��D���\��T�h��[�p>X�S̬�����Wm�V+k�j��׀n���7M�_�_ ��X�z�R�l��3Z�5sY�'���������~P��-����y`-���R�]6ݴ��&�u�n�2��Ȱ�W*��y`G� ;��*m+�aMP]��>�� �nE�n����R�V��K/��N��WI�6`mȰ\�Ur��x��X�8`�AiJX�9tz�꫘�t#7�e�8�����gV:u�خZZ�AA8E���~��7M�X�8{�U��?}��2�i4�aN�tٕ���RG}�� �y`��g�r�"H�i��]	M`����y`mȰ��[��\����z(|y��}w$�����"���Sn��v�J�m`z�ű�� ���n�e`�"�>R+�
݅��wb��n�����}_��y`[�����V��t4­R��.������4fЖj���f��q��t ��ј*��]6ݴ�	�5v���2�ˑ`[���W�$��}w�M�|,)�
�`��=�U$j�׀I�� �I2��q#��K.�J�Ҥ��cM��O^�0��R]��e`�?ݕp:t����V��9T��x�;R{+rO>�_M��>�H�XB0,!@���k�b�D�5�,b$��F�q1��05F�A�c�5TuD�$$)maH���V`R� �qMJ����|�m���o�srN��wSR��v�L���l�>�ٕ�vG�/ ݎ]�mܰCwI��9dh����)�#�9�u%�Pt&��V`�0�ֵ5 ��"�L�m��z�鷳v^�r,�6e`Y��[.�&��e�0��y��RD��,����;.E�uH��+l��ƚn�ۑ`i�+r���_���O^ wj\���۷WIݦ���}�̬��X�l�r�JG�, �� ���
j��0ˑ`Kذۑ`i�I��1���}�.f\�e��5#G�fm�h��]Z�N�ó]���NP�;��g3��zΞ]c^��Xp�y�\���8s�! <d5KE`�%�5����UD�2=��i�]����d^v6XѣP�s
�׬��ٛB�g�J&�f�Vř������֒��WBa�;���nn�l��6����vV�َT�g�N
Tڪ��Z&��e��¨���{�&����F��7��̕'5��b�8퀬gY�gv����ORj4���J�WI��Z��,v�X�k�ꪯ�U]��������BM�۱��X�Ȱ���8`Kس�r�Y�,����V����;���o�~�dp�s�ulLۑ`[�T+.į��V0�9T�&C �y`�� �Kذ	,�)CM��e�0��x�UR{<|as� �܋ 7kd%b;Z�ʋ�����^7 ;������vW�L���f�;8f�2�;6�E?`���/b�;�"�U|���׀/C���mB,�$�M���tы�����4Q>}P�����w$���r�៹\��U�~����
����ST��E�߯ ��� ���^ŀ}$F[��RHt�m�߫��{��'�?��/b�;#� }�#��t��C��v�X�\�<�}�� ��:i��Φ�.�mb���i�$	���]��V[P�E�9!hh;f �v`mf�nb�i�˦�Xн� ���^�W�$�y`��n��:Cm`�"���=�<�	/�Xн�=UU�f)�G�>�[,ev����v{�M�}Ͼ�� ~�J����10�h��@�$*�l�HBHS�4
�5���n�w=�܇T���[`�4鎕��?r����X|\��;#��s��� l��M6�t�;���0�{�������n� ��R�uv�[���,���Uu� �Ʈ��f��Ƹ�ng7�OLoj:n퀪�(��j�����N�v8{�ϐo��X}�#�N�$:i��v8`�� �/b�;#�{�Ie{̫�lT���Cl�$��v�`�� ��Г�$]۴	�N�0=\��y`�?���r`��%�ăQh��`��*�2?��}��RE�lN�h�
��;#��W����$��v��X �����UT�:ӡU�[i
�=<�˶Sc�]B��<�;�UkAM�C��׫��M��0�p�7c�ڗ�{�_ �y��5Oy��[`�7e7B�`�� �/b�;#�;3�*��9Wa=_��I��n�'v��f?�� �;0�2��ˌ)U�QB�T�����?y`�?�X�\�r���� 崙�Z*�ӡt�v�;r,�U����߻]~<�eȰ���|FH~� �U �
�b$��1��I��A�z"�(�l��5���2�9��Ll�����i�p3��i�%frײ�ŷ%�=r)d6�e�{k����&9���e��V ���v�d�t��-�p��"k��tn��mVهH�b���Դv$���%嶳:��F{�px۞n��2Y{X��v�F��ٕ)s�ԨF�c��	���%M���x��Ӷ�m��0#`W��J�aO���Ozy8���i~f�۫�鶒ޗ'�z:=�(��P�I���q���.g�7WT�m4:-��{w�Xa�eȿs� �߼�����Wv�P��ݺ�;p���URF���{o�X�Y��I����-�bv0C�`�?�Ȱ�{�W�o��`Y���V���m�l�'nE�nɕ�v�������z�N�[t2�|n����2��\0��N܋ �WP�d���[���d��Z�^��$m�2���Th��z��,�/�Ǚ��vs�v��>�#�vGv�X�XSe�%�HB���O ���~�|���@ �����My�v�I�~���v៹\H淪0�]:t"��v���~��;�ea���-��}~��>A�%�ut�m�N�m`�e`�̬��X�����L��`_�߰`%wn�)�� �6e`�\��o��>�~��7d��=U���=lC�|-�ӫUv�.��U&�Ѕ�d�B�n5W?��|o��^m���wfP$���[u�{����Ȱ�2���_ ��X�d�[lwwI�ݳ ��~�$I�e`�{+ �T��m�T��t]��nɳrO>���s��a1$u��B0'��='�`���vE�H�ne�"��O3�tX���6*�
I)5�����A�YB!Lsm�a��J�I���".`���HU�!���P�H�5�ܾc�=�35�ܺ��*���6�u��c��B�r�"k7�Pї��Sxy�8y��]j�H��e�`x�xzH���3{3�7��h&�2L�R3�5�S"4r�f4#�d�Di�+�k!	Ĝ�����<žRV�~�S��4	Q����	+�
f2����Sؠf34MabK@i�X��9�:6�J��M��!#)Im#ZB�A��e	V%��D@<Q��"@$! B1��$X.�C��P48��Q����6�����/��r�s��TUsz�=0�ذ� �ն�+����i�$�}��?}�i�߾�<v�X�X]��_���T��Xdp�=^��/�����;�X�{�C�P��Q9BGUuJ��K�n�broCbs	�&r��ݮa�F0�N��ـN܋ ݓ+ �6ez����� ����YJ��X�:-��nɕ��\�$o��}~��'nE��#��{+��Be4�`�{+ �;r,vL�v�����݌�۬R�?y`����&Vk��Es�dTa��D8�T�7,���&�*Pݖ����v��'nE�nɕ�v2�ˑ`�U�$���j�vmq��$�m��59���I�:ܨ@�[������Z&�)kt��brS�o���-�l��;.E�N܋ ;�%&4ݵWt�M[u�v2��T����{o�X�Y���H+}���+ -��n����v�X~�r�����7��V�دE]:�IӶ�0?r����X��Vڛ2�=�ܪ�g��~0J���YJ��X�:-��nɕ�v�̬��}7$����'���
}D2`)}�I$PBI��%��:�'�bo�G�mF\jfk&�C��W��b���̷�-�J��3En\�����Щ��Wl��:����	�2WC�aW�)�(=��;��g�Jt8�ǝ��8t�'[pS���r�KM��X�6�q��0!Xܝ�i�H)��i�9��\v�h�\u�)v�9I�����qb�7N�4�������קp���jR˒��XX��;�;�����˞�h5��=`�g�E��I�Ԋ�\Q����Z�bs�����Y�-�Jbj��v�O�Xdp�7�"��	=��{ܻ��lWi���`�� �܋�U�	=�k��X�[R�v&��h��l�7�"�7d����R[�{+ �y��:�����CLO��kR��V�l��;#�;r, �ʔ�n�cI5v��ٕ�v\� ���0�*e��I��3$��kX���:����nyeٷ���G:n�:���V�
��J�v� �;r,v8{��*���{+ 崙�|WN����v�;3�]�9��

����
��a$�>T�_<�q��>�&V�r,v�J�R�m[���0��v2��RJ\� �����%e�Į�;�`z�o�� �_��	��n��r�&�Wi�u�v\� �9UU��x�	<�`�̬���%��$�u�"�(ɴHFc�i�+���Z�i6aY�P��0�pU�f�*�n�US������0�;�X��uH���T�v2�+f68e�Ga�+ ���p��R��Mۤ�M$��0�fVI>��}71 �$E�	�}���	��آ�
��cT�v� �0	��M���[�{��;��y|J�ҡ���ـN���*�'���o���8`�Aj]�wV�C�V�;�ͣ�c��*1�0{th�'=�ٻ���C����Cl�7c��I��vG�A68`�˵W�퍱5tݳ �$��;#�68`��=\����U�,v�Whh��`�?��n���+ 6R�wi�U����`c��0�L7'½D{��[E�H���؅��V�B���l���z����=�ܓ��i��֩Mj�Z�իf�0�L��8`c��wI���_~K]�l{P�QN���ƌ%�bVf�t� e',R�ј�O]=´����>|{�Xv�,lp�>��آ�V�(�5I
�`[��	�� >��I����9ʻ6y5Į�8*��i��~�����7r����m���E��Ҷ� wdxa&Vղ^R��XkvYJ���n�Ճm���XV�xۑ`vG�_8W9UR�D(F�wN�_G%+��p���:4t��]��I�$5��!/0z��=�r�eXsX�u G��ō����[M(g�RE�r��sn��l�8���i��
@�u����'E�z�v�5�=pX�MI��{�b�f"To`�c31=p�ݼ�����'t:ʺ�¯�W�(��'es��뎎6�/$��$���U���F�u�^����fm%��L�M�-��i����Nt�n6cc]�L�8��IM��[�M`��*�h���whh��|�r,mȰ�#�;	2�a�vZm;�M�m`nE���I��wnE����{��!Z[E��m�w޺m�e`ۑ`nE���i�t���*j���W+�|���v���� �r, ����P����j���;�"�&� ����L�iu�:�*a]���ʉ!$���\�݊N������Hc�%�;m�<�<v]q��]9m`c� wdxa&Vղ^6�N	��[I�`vG�s�]��9�s��Wy_|c'r��r,lp�>�ȭU��n�ؚ�m���+ �܋W+��.�<�`���mȭU�[����L��;�"�&� ����L� �mB�t�E%j�n�X������;�"�=ʮ�S�j��� Lq1���:F����2ms�#9��ۛk4�̱�2s������F��g��ȦVݹ$p��D��ݺ�Zi*j��;"�Xv�X�� ;�<�$آ�U�MYMRI[��^$p�9ꪠ���.]q�a �Ip@(�@:Qג���>��M��R��⤩:wi���*�{����xdS+ ��/ ���DU�C-���0�#�;"p�:�K�$�e���m�M}�v<�r�k����΄p���0����6�Ǻ5��K�vU��uwbj���ȦVղ^$p�� �n)e[un�]հ�5n��ȳ��W�Wg��� '�� ����gN���Oޘp9��ڮ�|�������;�"�>SK��)���ګ�V� ���ȦV���f䉩H|���$��	!B�`���R�����rI7iT�t����Tշ�vE2����	#� wdxWAJ�[j˾6U��	A#H�6��U�X(�.�������Ƭ�E��i�Wm���$���:�K�$�ݑ��L�l@�.��$*;-��I0�#�;"�Xv�X�N2R���-���0�#�;"�Xv�X�� ��	˫�c�V&�o�K|{�V���M��%��xe�zʶ��Z��aL��;�"�&� ����8`����utcr�f\��Fc���d�`�!��QV��B�5�%!!#��+JD��$$)�*�)>�,�!Lc�0)� ���3({�w��[�x�~�9�T5Y���戛Ì��Ƙ��J�Ԕ%1�	�pf�G�] ��I��珊����u�o[�Hc�
80�}�5�Зe�fYT�Si�4	D�t�W���[���.��UרL׸���C^�,�c�@�a|�a��zF1�����^�]�&�KJC��m,���>)����X�*J,���ƒ�)��
�B,"��U��3i<��M>oz!&�9�L����H� XXX5%�� ��$��G�B0���݈g����!$F1P�T�	�M�Y0��'��d$��D�$D!!7)f�:�k����	��3��@+���	�IEt�J�2�B�A���g�n|b>%�\II��Mee�Hh%%�2�nݣ���K�}5��pY�e��^;�5tˌ�K�D��rX0�q�e��:C��:Cϟ�(*�����Y��u�.�駶#X4�[��u�D!��h��P�5��Ga�W6Й :�&�0]gXq�2Nn�R��u�!p�n��9b����rYǃ��0��3�Ƙ��cnhȩ�В��b8�l�Q�4n��4���НF[0�%�(��s��;6�Z�j@�J1F�rӴ�I�6���!6�m�N��u�}�A�+u�"�^n,�a|�Gb}v.�a�RQ*��f�� :d�	�܁8]Z-�ں��G�ڈ��a����0�[��p���:�l�Gr`݌$�d6�h�����k>�,"@�ڂ���&�D���a�݂˕���m�E^�nSq[f��VH��<ALT���&��(z�.���bԯ�� �.vD�=�n��bGEx8�-�@����[m!�	h��v�5�рt�tq��9nhu2r�u5�$b�e���9	�� +�1A���3\�A�ۨx^��"�p�L�2��[c�a��|����'O6��j��ŏtE�۳��U��E�s��.4�=�0�����nSf݄.�kJ�F0o 4��Z� �ѵ,
�Z�b�'[3�s�x�{V�5�G�R�,k���f�B�D.�9N��fD;�����$k	h��ې����GYw����F���*Ogg�ԅ�b�=���*�՝�W�]�b�p�l5Yu�����p����阁�-V�z��1�l:����.��.���"����ơ���s�H�Ϛ�CӢ��a�� ���C�T&�����Ng(U��ED'�:�����U.��ڒ:M�{3�[Ur�K+
��r��r�W8$�,���rv^��(t��Z�����Ԗ�����1՞݌��M6n˛[xp��]�ɩL�q��e*띹WT��
�����gZ�0��m�x�C�ꎃ6g]��g��`��{\�Ѐru�\��Br�e:i\񗛁�)�ãf뫚�]hlWA�!��2�R2�mF8�l��Y��z~�;wt�@��p�"mt��D�A�PB�X�ATM
��C���
x�b�� ���:�-�a��8(]�Ը�t���q�e�M�YT�Q�g\m�W���sp���,��L�v�m��v(�,٭��A�fk��=�>}�q܆����-��uq�Ru��t�L�m5�]���E��v[���['RTkv&�&�Q�m-ԫbWZ�u�g�t���\8e�b���ݺ�Gf�3�p(p��if��7,��.�1W��$��i$�̮��7�[�,u�ʹe�Ny9Y�&��r��aU����C�j�.�;�R�����ݑ��p�UW>A���u{��bC[N�]%l�� �#�ݹ68`vR�V�;v��Щ�o �#�ݹ68`vG�آ�U���tĄـul��M�ݑ�].�O� ���*�ƅEӻM�68`vG�ve`[%��QtKjĮ��V������n����omטg�.5��wb�hN��7Q���-���0�#�;	2����	�� ��	˫��V�&X6��I�b xq��WZ���ٹ'�{���vG�}����j��`0v� ��/ �0�#�;	2�a��:�*ӻMݶ�2�ِ���I��wnE�|�. �1Ֆ�1�V� ���Uo�{����,lp�>U�8�԰$�U+�d��-DU6R7RS�n��9���yH�K-c%�y�:��l��+o �$��;�"�&�UW����
�#ޥWc�@U���;�"�&� ����L�lA2�WO����e��	�� ;�<%Ur����UA��@oY���7$���rO�'�ǔպ&A�S����qӻo������K������ӑ,K���w�iȖ%����s��r%�bX��~��0�5s2�L�Zֶ��bX�'����"X�%����nӑ,K����fӑ,Kľ���iȖ%�by���Z,-s�u�B�Om���/9z����Ť��aZ7L�V�e�jS3v�n�[M�{�ı,O~�{v��bX�'~��6��bX�%���[ND�,K�������N��N����CWRj�U�|ND�,K�k��NC�"�șĿw��m9ı,O�O߸m9ı,O~�{v��bX�'���:M�Fe��]�ӑ,Kľ���iȖ%�b{����r%��!�2'����iȖ%�b~����ND�,K��Jt�Y��k4Jj浴�Kı=��xm9ı,O~�{v��bX�'~�{v��bX��}�}]��9��iȖ%�bS�l��0�$�5-�4m9ı,O~�{v��bX�'~�{v��bX�%���[ND�,K�����m�!�#��*����mAV��byP�V�I�0Vv��lM�fX� �X��3�yJ4�|���N��N��}��9ı,K���bX�'�{�ND�,K���ͧ"X�%����{`B�W+u�X������iȖ%�bzw���Kı=ϻ��r%�bX�}���9�S"X�����Dm;`�Kn�m�!�.�߿p�r%�bX��{��r%�bX�}���9ı,K���bX�'��}ڙ�7e49�t�t�Jt�O{���9ı,O��{v��bX�%���[ND�,�ȟ~��xm9�!�>����Wk�`[e��m�%�ߵ�ݧ"X�%�~���ӑ,K������Kı=�۴�K:S�:~��yǳ-l]P�2�a�R����\�e����˰0�emc1�S5�1�ݙ�F�bi����EU�[���-*k��	��[���F�]�#��m�nH�B��	V�!+tA�۴�s:Km�ہŐ��c+�]�5�6�^9�x�m�s���E�)s�0�\�NJ��qQ�V҆�=��8ݸ7.25�@�����j�w^�J]L���=q���[���������1��F��d�c�&�d�y.�u�5�Jq��'t8ƛ�Ϯ�ur�\�_ؖ%�b_߾���"X�%��g{�iȖ%�b{�w�iȖ%�bw�w�iȖ%�b_~�{&h�������m9ı,O{;�ND�,Kߵ�ݧ"X�%�ߵ�ݧ"X�%�}���ӑ,Kħ���)�h�$)�l��iȖ%�b{��۴�Kı;��۴�Kı/�w��r%�bX��w�6��bX�'~�'x[��֥�Y���r%�bX��]��r%�bX�߻�m9ı,O{;�ND�,Kߵ�ݧ"X�%�߉׼�2]\53Rj\��r%�bX���m9ı,O��ND�,K��{�ND�,K�~�fӑ,K�� �g�~�3?25��scs��W
�"�m�f���C�Q���֔�1Vl��ۈd*�j`U��Ȗ%�bz~��ND�,K���ͧ"X�%���o�iȖ%�b_~�u�|:S�:S��ϻرT\0`�x��bX�'��{�NCJ��R
�$H)�@���:x�ؖ&����ND�,Kϵ�nӑ,K�����'�>)ҝ)�����\�j:����r%�bX�{��6��bX�'�k��ND��C"dOO���iȖ%�b}���6��bX�'��fvD�[�usWF�Z�ND�,Kߵ�ݧ"X�%��߻�iȖ%�b{�w���Kı>���m9ı,K��/L�3Z.���.��]�"X�%��߻�iȖ%�b{��۴�Kı>����r%�bX�����9ı,O���Z��Ο�w7c�d8 @���t���;6�F(m��rd����"�R��hU�%Zŷ�ibX�����9ı,O���6��bX�'�k��ND�,Kÿw�ӑ)ҝ)��������(h�-�å�bX�{�xm9ı,O��{v��bX�'�~��"X�%��w�ͧ"S�:S����xz�&A*�:|:X�%����nӑ,K������K��+� )R1b0(� ,t>TaAND�&�_�fӑ,K������Kı<=;����ԷS5.�v��bX�'�~�6��bX�'���6��bX�'���ND�,K��ݧ"X�%����{3Z�W>t�t�Jt�O���6��bX�'���ND�,K��ݧ"X�%��߻ͧ"X�%��~G��`�b�
�j�ڒ�ŏ�I�~���[�1�qcu��7l(i�ZD�g��eֵ�O"X�%�߻��iȖ%�b}��۴�Kı<����r%�bX��{��r%�bX�g{�wR�f�[���5��iȖ%�b}�wٴ� �IÿwI�$�{��nБI�=�I��N��N���g�a�A��Q�<��Kı<;�y��Kı=�۴�Kı>����r%�bX�}��m9ı,Jy��ܓ3F�IMJ[��r%�bX��]��r%�bX�{�xm9ı,O���6��bX�����M��m9ı,O~��	ɖ.[$ѫ3Z�ND�,K�~��"X�%����fӑ,K������Kı=�۴�Kı<�W�e��sX`RE�жai,���t���H웍���#ɬiH�eڹl��F3Wa2	Vy��ҝ,K﻾ͧ"X�%��߻�iȖ%�b{�w�a��DȖ%�߻��ӇJt�Jt�?z��2�uL�O:|�bX�'�~��"X�%��u�ݧ"X�%���w�ӑ,K����i��N��N��>�cTc-�2��qȖ%�b{�w�iȖ%�b}����Kı>����r%�bX��w�7��ҝ)ҝ/���JݑM3���r%�bX�����r%�bX����m9ı,O};�ND�,K����ŷ�x��x�Nt���)]
JUdѴ�Kı=����r%�bX��w�6��bX�'��{�ND�,K�{�ND�,K��Ioٓ:j�JK��V0;{f�k,�@"v9�3J�p������Ԙ'��l���{��K����S���T2�:<V.3���i��		6�l��µ�lnpm�ôw4!h��MǳN*�Nv�"�[Hn�l%�X�8��`_nKƹ�RW\h �6�H呢CY[e�
�=k�|���(�4��]i�k���I�$0���\F��k0Vo.,N�#��b�,L�z,r����,2"(�h�כ�m为$붺[]I��"���C:0х���Y)%�q�!�.���ֱn%�bX����m9ı,O��xl?�O"dK�����m9ı,J{�����4a$.�l�ND�,K���ͧ"X�%����fӑ,K����iȖ%�b{�gxm9�2%�����d@TA��-�ŷ�x��x�����ND�,K߻�ͧ"X�R"}����ӑ,K��;��m9ĳ�:~����cJԨ%��O�Jt�'�w}�ND�,K�{;�iȖ%�b{�w���Kı>����r%�gJt��g���5��4\�t�t�Jqb{�gxm9ı,Os��6��bX�'��}�ND�,K߻�ͧ"X�t�O��-��a*�F;iN��3i1�4��&�ܹ�[u��֨0�+���t�T���5&�ֵ6��bX�'��{�ND�,K���ͧ"X�%����nӑ,K����m9ı,K�g��fXkSSZ�5�fӑ,K��o�i�|���	x/��D�K�k��ND�,K�g{�iȖ%�b{�w���O�S"X����ź�jj٬�h�kSiȖ%�b}���6��bX�'��w�ӑ,K��>�siȖ%�bw߷ٴ�Kı/�t�p֦V�Д��b��<C��.|���[�bX�'��߳iȖ%�bw߷ٴ�Kı=����r%�bX����&�Li�l��iȖ%�b{�w���Kı;����r%�bX�����9ı,O;>�fӑ,K���GL��WM���X�t���ύ�S�\�`vf��/���������)��BS���,K��o�iȖ%�b{��۴�Kı<��}�ND�,Kߵ�ݳ�ҝ)ҝ=�x��h5*	ryӑ,K���w�iȖ%�by���6��bX�'�k��ND�,K���ͫo��~\^�la),��*Zk"X�%��g���r%�bX�����9�!�4�1$J��I#,z�z��Ф�XX ,�qu�(i0�HH��Mj�c	5��Zwyސ�ŬHU��t����kX$H��1]��؜�F	<�y�e5)�]��1����rHB2)��-(��bː�ۮ�B�Xs���R�A!���0p B��pnBF	B0��,(T��(B1��!!AwCq�<۪j��ٶ$	�<g�f`K	����"oP�d.l&��D�S4�o-� Z��J%�L�*K1�0(Bb"/��(&�|T�H�M����U�� `��x/N�ȟo[��9ı,N�_v�9ı)�����i��F�<���N�Kߵ�ݧ"X�%�ߵ�ݧ"X�%����nӑ,K������r%�N���{{����gg��å:X�'~�{v��bX�'�k��ND�,Kӽ�fӑ,K��>�siȖ ����"B)S��:����Çz�����l���#I�qڧ&lF���u�ճY��s5v��bX�'�k��ND�,Kӽ�fӑ,K��>�sa�'�2%�bw����9ı,K���fA��3no�>)ҝ)����;6���9"X�g~ͧ"X�%������Kı=�]��r%�bS��}��@�(C�KJ��>)ҝ,Os��6��bX�'~�{v��bX�'�k��ND�,K���iȖ%��O�{t��,e4��w�>)҉bw;�siȖ%�b{��۴�Kı>��}�ND�,!�!��Aa`QO: �;�~��ND���/���qȝ+VYf�m�"X�'�k��ND�,K����~�O"X�%��w���r%�bX�����O�Jt�Jt�����+ekf#�X-��K،;N�\.VJ�	��q�@e��uՌ�0 ���QR�X���|��=b�Kı=ϻ��r%�bX�����r%�bX�����9ı,O}�s�iM5%�A���t�t�Jt�O�������r&D�?g��ͧ"X�%��u���r%�bX�v}�ͧ"~2�E�Ǐ�+�B�cd�X���?g��ͧ"X�%����nӑ,
�2&D�����ND�,K���ٴ��<C�<_��O B���UKf�n%�bX�����9ı,O�>�fӑ,K��>�siȖ%�bw;�si��N��N���g�[����no�r%�bX�v}�ͧ"X�%��w�ͧ"X�%����ݧ"X�%����nӑ,K�����
�����1���Ѐ�_'�Ʈfj�n���yFX&�7�r����M�tS��m	���f���M(P_'�v�� rq89��ڶ�{��g<���2�W��Oa�y&��=�F�1n'�C��ۂ�r���:��ݮg�NQw&��nw7	Ok��,�g��mZ�Mp�s�5����˶�N�1��%�H���wn�x�R�CT�29�8�6��*��5����t�0�|E�l0U����8q�1�Fq��5�u�ݘ�+��,������2�Ĵ�y�ӥ:S������ND�,K��ݻND�,K��ݧ"X�%��g���r%�bX�}�n�JhɄ�F�]k6��bX�'{��v��bX�'�k��ND�,K�Ϸٴ�Kı=�����K�S�����ߗ@[c��å:S���ݧ"X�%��g���r%�bX��{��r%�bX����r%�f!����j

�ZU��b��<C�(�2'N���r%�bX�g~ͧ"X�%����ݧ"X�%����fӓ�:S�:}���M�L�T�Ȗ%�b{��siȖ%�bw���iȖ%�b}�wٴ�Kı>��}�O�Jt�Jt�߿�U3+̀JnknN�D�X����Z�'[��9���"�j)u�\�:|:S�:S�����'"X�%����fӑ,K�����l?"O"dK��?~��ND�,K����5k�l�T�m�!�}��m9)���"���&�>�fӑ,K���w�iȖ%�bw���iȖ%�b_~�{��jGh���O�Jt�Jt����O:|:Q,K���ݧ"X�%����ݧ"X�%����fӑ,Kħݿ^��kR�B�]jm9ĳ�2'߷��iȖ%�b~����ND�,K�{�ͧ"X�%��g���r%�bX�}��K��׶��f���ҝ)ҝ=���iȖ%�b}�۴�Kı>��}�ND�,K���ͧ"X�%�~��4=í��3CjlF4��5�X��z�0h��k���*NV�V4ءP�HD;AUm��r%�bX�{���9ı,O�>�fӑ,K��;�sa�	�L�bX�}}�[x��x�����6B!;K�֮ӑ,K�����m9Ȫr&D�>���m9ı,Oߵ��iȖ%�by��۴�O�TȖ'�j~����.����O�Jt�Jt����ͧ"X�%����ݧ"X��D#$���Č!	%*N�0�M�ϵ���r%�bX�~����K�C��㧐�TB��-5�o��2'�����Kı;��~�ND�,K�Ϸٴ�Kı=���r%:S�:o}�а��eپt�qbX�'�뽻ND�,K�Ϸٴ�Kı=���r%�bX����rb!�/�.��_5K�*��!�.����YG�/9vA��6�Vvؓ���uHS��FJ�n�Ue���/���{��}6��bX�'��ݻND�,K��ݻND�,K�u�ݧ"X�%�O�O��6d�R��O�Jt�Jt���nӐ�(�"dK��w��r%�bX��_�]�"X�%��߷ٴ�O�S"X����Rs$�7&�\���r%�bX�����ND�,K�u�ݧ"X�%��߷ٴ�Kı=����r%x��x������"��U[e5�o��@Ȟ��]�"X�%�����iȖ%�b{�}��r%�`l��ސee�����B1YI%aEĂ$��0)�7�K�o�}>)ҝ)����m����Vhվ'"X�%��~��"X�%�����iȖ%�b}�}۴�Kı>����O�Jt�Jt�������fq3 ���f�с��0�CK�Y���o]s�	�z~��5sv�F�k���6s>t�:S�:S������r%�bX�w_v�9ı,O���6��bX�'���6��bX�'s���j�TAQ��ŷ�x��x���ݧ"X�%����fӑ,K���w�ӑ,K�����iȖ%�by�wե�F&������ҝ)ҝ?}�}�ND�,K���6��c�dL���w��r%�bX��k��ӑ,KN�����e�PV���<���N�K���6��bX�'��ݻND�,K��ݻND�,�̉߷���r%�bX���;���Z�uL�捧"X�%��u�nӑ,K��߷��i�Kı;��~�ND�,K���ND�,K��� �,��Ą!�"E���?~$��Xf%��2�g��e� �م����!ocWl옪�C\�v�&�u˞�N�v�̜�����Ͳi��k����]�#7F�Rb�� ���wŇgcrf�t�t��0�n۫��˺�ݕ�!eɳ`�6��䅢8Pv���9�n�&�f��t�	*�r�iE�A�qa���2h���(jVWn�ar���n�E�4�����m�\�����1�4Hh�.V6mf�̱j��i��\�D��mݩ����Q�M����ı?�����9ı,O��{v��bX�'���6� '�2%�b}�]�u�o��{����F��V�M�"X�%����nӐ��r&D�?~��ND�,K�����Kı;��ŷ�x��x������XX���r%�bX�����Kı=���r%�bX����r%�bX�r�Ʊm�!�#�<E�B��:�k4m9ı,O{��v��bX�'s�w6��bX�'�k��ND�,K���ND�,K���κ����ɗZ�ND�,K���ͧ"X�%����nӑ,K���w�ӑ,K��9圯�R9H�#����I�ʶ�Ia�� ]��qAK�ևlF�Q0J��wN�袪2�eI�2���å:S�8��w�iȖ%�b}߻�iȖ%�b{�}۴�Kı>����r%�bX��|�Ȓ�9k��))�[x��x��w���r�q�MD�=���ӑ,K��=����Kı>�]��r'�G*dK��^�0�kRL�Xanh�r%�bX�~��m9ı,O��w6��bX�'�뽻ND�,K����t�t�Jt�O�߽�/�\��hү�Ȗ%�bw;�siȖ%�b}�۴�Kı;߻�iȖ%�� �����ӑ,K�����g�fY�Zhֵ��ND�,K�u�ݧ"X�%����ND�,K���m9ı,N�~�m9ı,O�g�~�f~�r�YVc[�
@��iH�=ep\�4cu͵��J���@�8��(X�Zo�x��'����iȖ%�b{߻ͧ"X�%����͇�`�'���M�${��t�6����t	�:~��鸝�bX�Ͼ�m9ı,O���6��bX�'}��6��bX�'rw�:%J3%��_:|:S�:S����w�>D�,K�{�ͧ"X�>0" �O@��M���6��bX�'���ͧ"X�%��w��亚�0�5�Z�fӑ,K����iȖ%�bw��iȖ%�b{�����K�� 2'�w��iȖ%�b_{���L�A�1�r��å:S�:{��=<���ı,?��~���yı,O���ͧ"X�%����fӑ,K����j��F�p�En�g3��Y��Iesl2A4�eBb����c��燫d�y1jm9ı,Os�w6��bX�'s�w6��bX�'��}�ND�,K��}�ND�,K�ge�.h��fY��5�ND�,K�߻�ND�,K�{�ͧ"X�%����ͧ"X�%��w��ӑ?*�TȖ'�d�̆զ�f�Y��Kı;����ND�,K��}�ND�,K���ͧ"X�%����ͧ"X�%���ݷ��h����պ��r%�bX�����r%�bX��~�m9ı,N�~�m9İ?x0�_^��ߑ3^~�v����x�����y�ei������X�%��w��ӑ,K��w��ӑ,K���w�iȖ%�bw�o�iǈx��x�ޯF�&�	�ePC����<�nWf��-r7��y���\�Y�H��T*Q�,q��:|:S�:S�����8�Kı<�]��r%�bX�����~E�DȖ%��u��iȖ%�b{�}$�H�V�娶�ŷ�x��x��wٴ�Kı;�wٴ�Kı=���r%�bX��]��r%�bX���C٥�q��\�<���N��N�����r%�bX��_v�9ı,N����9ı,O>��6��bX� ��{�"WG���b��<C�<=�_v�9ı,N���m9ı,O���6��bX�'~��6��bX�+���h��D8:BY�[x��x��ϻ��r%�bX�}��m9ı,N���m9ı,OsﻛND�,K��3u<I��\3��D�H�!I$Y�RR4"F�`F,�I#FBHA�	P;��'�'C����q�T��3~�H)�4@��4	`�&e�%�P �bp�y����8���\�h��^rO�$Y;!���*U̡� d�)2RH>KX@�D��j�i
$X���"�$a$$ahRao03D��`PC4A�a	h�����B+1�p�Q+D�u@�)�`�ă1#��$$HF1��1��,#*BCv�KHA��q86"���%ˡ����!�Dk-�X�)Y����vIB�gӉBN4��Z��,)�Ke���R�o,�b[�'�[��Pd$t�0*E�6)X��n��z8�8���v^s�cn5�I��ٺW�P�	����}Ū�ѭYc,6�	y�)9��U�����=U�.8���M۷cc�Vm��G<[�n��I��-40��X���lYse�ÆY�DqVSG.5�Pۍllu×Z#V�(�1O$�ˌ��.ܜ
s��m�#��k��p\
��Y��tQ)�B�B�u��ۭ��A�������P;�e���4b�ِ�
���	��s��=��n�}�\���ǵt�U�jxa�p����$��n�d���64����2�@Y�6�3�5Γ.�m�	(t���ybД�%k{q���S�+WeӺg3kk�ϲ�<�(��a4n���ѭ��.	�*M[0ջ(�JO(���F�-�y�<�렄�����g
F|&�$uG	7u/jՖ�E�[��܏c$��
p�@pqe���ۓthxi��t9���f��E'��7b8���Xjv������v��Ȏ�N1#��c9��B��U�i�����s��\0/u��&g�E�&�m�7�����n����;80n�ڳ�&�ț�k%%ӞZ]$���F�-c�.�.T���dGU*]5JK
�� 0ja����V.�i$�4�Aآ]��Rc-�륄���"ٌ[�ݩ�è��n6+�e���K@ghܡv�m��]��[�(�n
[��,�%�Ⱥ޻s3��4lôr��<Ocy�c�>��N9q9CvG=�6�K��d7	�N�2`�[6P����]�͞����j��H�t���;�����U�c�9�ȶ�QEM���6�+4��;/M�T���WN�cx�$91Q*��Plo�;;(}.�=�`�^T6����n۹]A�渲���\��5&�x4\�M6Ki5��n��Tch,*Cb"���]A9s 5ah�2([2n��v��1�:�j�@�G]�3���R��܀�47�H󾳇e�qӹ,B��܅����c�,v�-��9p��۔�I�jkW5����浊�� =D��ਟPA�T�D�Db'�x�� ��_�@���?���.1��(�^ܰ��U����7�dl�*��vۅ��.z������A�5!�۵ìp����M�!�9K������f�I��l�˓c�n��fr7LC]��
ގ7����m�<��fuЬ#��SS�{s�T��6�;R��ؕ�˦���K�͜R!YTֱ�E��L�t;�a4�L"�4 ֢��305+�sgq��]���{��B�g��{�rx�vku��UA
2�A��L��%�4�
S$���N�S�Eh*��ϱ|�,K�����Kı;�wٴ�Kı=Ͼ�m9ı,N���m9�C�<\\�n�2P*v���oı;�wٴ�Kı=Ͼ�m9ı,N����9ı,O>�{v���K1Cx��羄��ei�r�r����bX�'���ͧ"X�%�ߵ�ݧ"X�%����nӑ,K����f�m�!�#���X�AU++��ͧ"X�%�ߵ�ݧ"X�%����nӑ,K����fӑ,K��>�sΟ��N�����m���B�W6��bX�'�k��ND�,K�w}�ND�,K���ͧ"X�%���{5�o��w������*��m�3JT��qz�fX��zۮ�dkz����-��j�:|:S�:S��}��iȖ%�b{�w���Kı>�����Kı=�]��r%�bX�����D��+�-zŷ�x��x�;�fӐ�b�`�^��D�K3]�m9ı,O}�{v��bX�'���6���\��,O��[,�Թa2M\��m9ı,N�~ͧ"X�%����nӑ,K����fӑ,K��>�siȖ%�b}�;��%̅5�M��]�"X�%����nӑ,K����fӑ,K��>�siȖ%�������iȖ%�bz}����a��V]WZ�ND�,K��}�ND�,K���ͧ"X�%����fӑ,K���w�iȖ%�b}���ٳVF�1����;]��V6���E=�8��jQA;���r�	bv؄⪎׬[�bX�'��{�ND�,K��ݧ"X�%����f����&D�,O�~���Kı/Oݟ����kX[35�ND�,K��ݧ!�A�DȖ'����iȖ%�b}���M�"X�%��}��ӑ,K��>�\�I��Va.f�f����Kı=����r%�bX�����r%��Ő�N(*�hD���@�XD@���Ҩ,M��;��m9ı,O�k��iȖ%�b_{��s&�au��3Zֵ��ND�,K�w}�ND�,K���ͧ"X�%�ߵ�ݧ"X�%����fӑ,Kħ�����ԙKu2˭M�"X�%��}��ӑ,K������v�D�,K�����Kı;�wٴ�Kı;���'n�S!s4�f�%ͽ\8�b.	%�[����\sS۱1����s�)8������bX�'~�{v��bX�'�w}�ND�,K�w}�ND�,K���ͧ#)ҝ)���}�Cke�lcr�:|:X�%����fӐ�G"dK�o��r%�bX�g~ͧ"X�%�߻�ͧ��N���>�}>+��+��Ô�R9H�����5I��7c��� �e���ڡӦ�M��+�nO^�}�vnI�~��rI�F�N �&�C >����
t黤����� �c��0��x�v��ƴ{^UǦw=��Q˻a�k��� �E�D�T��d��V�@K-zm�p�;#�ջ/ �0f���hv�[vݳ �3��r����O^=~��>���D�*�l-P��&��v^%Ȱ�s�\�%��� ���n�)*0N�X�5m��"�/ �c�68`[��	(�U,�R�ҧN�w�}�� �V�V������8�!	�O�/�UuѦy�\��mY�{JtL�X���[�o0
~���wk��;������٭5s�`ٺq$���CZV[��`�g��8��m����k;��*��X|��'[ 5�4y��<Lq�Y�{fs�����0jxLq�4$�&DVB�fල��F]�lX��-��jr�����Hj����k�bd��)9�fz�<Cc7t2�9����i:H�0�p����ǉQh�[/;T��I�;jTn�;�"]sa�b�6��l���`[��[%�zo���I�(Kꪎ�׀j�מ�s�Oz��?v8g��%�����nc3�J��>���|�+ ���v^����MHV�[m`l�Xv8`[%�z�T�9��m���x������ڴ����Ixv�X�X��ی���)��,�]��b0vζE�Ӵ�"\0����H^v�ۘ�㖶N�;���^ݹ�&V�0إ%X�cL�&�7xdp��W8��&V���Ixv�J���E1�t��0�X�ᇫ�KT�� ����v]�T+hN�۬�8`[%��� �ɕ�l��V�m*:h��0���s�����6{�Xv?ǀ����ĵ8���L7K�
���]uv��gB#�N��I����s
jt�$]��:�K�7d��;����O�>�}�x���w��Ѧ��#�x�X�p�:���ul����v'bC��:bm��0�%����h��Z�!		 FPe� /�CG{�Ͼ��9��lܒ�(�ۡ���ـuM��j�/ �ɕ�vGv(�Yt0�vI�V� ղ^�ɕ�vG�v^ o��r�R֪�I#"�Q9k�)(]/c9�Fٞp@ջ��s���VZޯ"61U��+ �v�/s�_�����ig���m��;#�ݽ� ݎ�&V }�wr��Ʃ��t�l�;��`�� �d��&� ښJv����m
�kܪ�/Og��w�7$���܊�	!Ab/�9{2|������;�e��vـ}�e`#�ݽ� �0�Ԗì.1�G;`Sn(�.;lt/m����
NNS&���%\�,���Lh*��0��X��}�e`lPR�V�wt�fݽ� �r,�+ �3�\�G����,-���v�=~��>�2��� �ݗ�n�w/����:wm��L�dp�:����s�JOg�k}��LWm	��u�vG�v^�0�L� �����?F�iX�(���#5���]��Fxo#����)���Xd�Kn�5]n�-�9v�5�} =X인W��"�RB��96�/X|�����i����96֭#�q�ds����y�G74�N�H�9���ݔ*+�wf�q�x�<�^J&1ی\��Ϯ�'<�՜�����!Q��:`�;)����cLch�Z���}�˃��u��s�Y������_�c�sy���ט��t����P���g�������q�Μ6nőa��by����4[=x�p�>�2���SbN�S�E�"ۼv8`l�Xdp�:�e���)RwM��;୬�+ �0��x[%��
4���v��m�68`[���K�>�2���-��wvZl�:�e����}�e`�� ا�x�����RҎ0,��1�Գ y!3;:�4�m@.I��b�S[�h���I�V����߻�X�]01ov��jj��]�L�N�m�ݙY9�r�tD�D @y�M��}7$��߳ &���Uʤ������e1]�'M[u�zy��>Se�nE�od��>�e����]Z-6��l�mȰ�L�/Og�#�Ȳ��N�hE�x[%�l�Xv8`[���o�*:��Z��K!br�U]����Y;:b�����%�%K�o:�l=1a7n��L�v8`[���%��)�ch���lM��7c��6^ vH��X[��R��t:)��Zl�:�����mQ�(�GB�0#�0�0!`F
,�O���'%%ICN.��a8zkd�%��/��#�ωp��.�����D1j)	��G����n���'�`��߶�kp�d�T\��5]$�H��A��q�� {JD��3=P�FH�B6UA�$ �����*b�"�&��{�t1�>�̷F�7
2f��o,��C�H	B	oRJW��ͫ�
����w	�fzyD3*>S/�h�l1°!�-,��}!  ���0���D��K���i4�B(h��O�4ki7��ԺP��$
9s$�����C0�z��7�_�_�|��D�iHM��qP��U��qSH�����0S=ĪUD5�! �"21!�0�"(HBF*���!$H�A�����= >E��G��8'�k5̬�\0�-!`'V[Rjջ��q)�y�}�dp��9\������6W�^J�e�j��x�L�v8`Se�d� >컥jYi�9�4qֱӽ�;n�yݙ�x.x��\n���t$��)e���5Ud�eT��6��޽�6^ vH�\�s�}����[V�i;�WE�vـuM��$x�L�dp�s�G���[��t�݈�� '��od��6G��^ vP����N�n�ݷ�w�e`G�Ͼ�ɛ^ � ��d%,.d�K�%��J@��!�5Y�3����ww��������{1h�Tțu�I0��x$� �d��<�g��{j��7Gc(��rR��-�bn _`8&�D����a�+�7L��ڻ$�P+����޼ �G�w�ez���O?��Y��"�
�Wv� &��ܪ�RFｕ�l��uvK�&�����TƩ��m��Xv8`]���#�6-]��)�M	�M���W8�{<`�޼ ����L��!�펚N���t6ـuvK�� �d��;#�uUU\���$@��[Z�]5�SF�� [�(���n�p7pmY;�s��Hʜ��dܚv턶
�q��m�t�ͳ�Z5Z��B}�kUi�
+[�p���:^��G�.�'�.Y���-A�q���2���C�w@v����J��t�'��0�;�5�ֺj�V'�/O����!��:um��{��P��8l[.&J�m�0cn�3��:Ku��ԖP:���7�,��a��Q)�s���/�x����㖹��y�[�u6�{B��ƌ)�h+� �?<��+ ����^ IJ�FS��i��Nݷ�w�e`G��^ I#���馩;��lM��$�Wd� �G�}�2����j��wvـuwe��<��+ �0�JV*.�YlI��w�$x{&V�0����ȓ*k���܄�kpѻh���d<�gl�n�<�Ӯ�� ��<v���kGB�}��ɕ�wc�ջ/ ;�<��j�o)�юVx����ϝ:q���^
d� ��fKs]��'�w�ܓ�>�+ �J�v�t�wN������l� ����Xv8`jUڷB.�4�[w����+ ���l� ��HwWm46�۶��Xv8`Se�vG�z����o���kHO]ɹ�xN-�Sv;gс멭cs�4�ؖj�s�]8��K;VІ�e�n� ���un���<�+ +�K�X[�j���ـun���<�+ �0	������.��t��n�d� �d���UΔ��(��R��	�$�$ RC�
�Ep�w���'/�w7$��g�3-1�j��x�&Vݓ+ �ݗ���l�wW��v�C��u�wd��=�UUm���}�<�+ �r��^կ9.��
�(7nM��cTvq�ĜA�,�W
(�))eP)TN'l�M��v^ vH��L�vL� ڛJU��E��n��G�}�e`�e`[��JU���]$�Cn����ɕ�nɕ�un��� }!WIݠv���n���n܋ �}��^0�! $EaN���$	ࢁ�!��;�w��z���5CWj�ـM��$�l�X�p�=\��z��l��n��̉ѵ'���iِ^��z�.�-��v�u�Ƈh�EMUCr�"�e6���z`d��7d��9U�K���E���@�鴩ڻn�	�e`�2�	�"�:�K�UW8��{֮��Wv�&۬g���M�ղ^�&V��12ۢ�ӫ��n�`�"�:�K�;$��;�e`�JU��EӠt�+k 6H��2��X�Ȱ	\��������ˌ���6in�ۻ<��!,�����6IC����)��2s�نV �̀��mV[1S$9��AN��Z$̯V�ݵ-�ejd`�%Hd(�5��m&���[�6Ť��rc��ܛ�נ6�����՞����]��bzM/(��.W��/��\��!��g�o]���[���.5���L�∥���ˡ��j�Eݳ�f)]6�3Z�2������PC�C@ ����93��K�UѼ�z�Y��m��MX��l�3�6I�C��E�J���t&�t�m���+ �&V�0l� $�+�&���V�Qv� �&V�0l� �&V VĢ%+�tՖ]]��&� �#�&ɕ�M�+ �)J0.�(�J�7i� &��	�e`d��&܋ ��pR.��N�6�6L��&V6�Xݑ�����	_��:��ڕ�u)Bm��p�`�nYp�e�ؘ$�0Q��P��Bu��V�|ﯞ6�Xݑ��e`vT�˺uj����]kSrO}Ͼ��ؤ�tm1�$	A�@Y�F�H�� ����x�}��n� �e��t"��t0V� vH��2���n܋ 7iVԫwt�N�n��o �+ ݎ�Ȱ�G�Aؚ�m�.�`#��r, �#�;$��>�IK��nժ�l@� �8�q�әD��c!䍶��#a��yyxtۘ#\<�V���ـn܋ 6H��2��� ݈��*颋t��v� �#�;$��&�v�X�D�,Uh�v!ݫm�d��&�')�S��s�*����|�"�	���%X�V����u�M�ۑ`�6L��1U��Ul�4�0	�"�	�<l�Xdp�=\�)�y�Y�����@pPv	6��4��b�w^cQ�r\�$�<j.R63יہ��$��6L��8`nE�V�J��i�mշm�d��;#�6�X�#�	 �:��@���0	�"��6L� �Ģ(һ�	&�UR�~��	=�nI��}�r_S��%�ȥ,Da+H�L�B4�%
Z�����"VYt��N�Rnݵ��<�L��8`�"��R��v��z�܏"�#mχ��V��ʜCFِ�p@ֺ��q�'��
FF�p���6�w�����n܋��9ϐ=�w��J���
�Cm��;��=�URD��, ��<�L��&*b�uv�jĄ�f�r, ����2��p�	5JV���>[������ �ɕ�wc���/ $��J��6�۶��L�{��7���@��&��򂨫��EQW�"����eQV�*���ATU�*
����E_���*��@V$ `$E b����uQW��*��Uj���ࠪ*��QW�(*���ATU�*
���PU����₨����e5�ivP6v���?����������@@ h P(�"R� �@+�b P���V�>�>��    AB�*)H �P�EP    )
�)� H� *@�J����  ���0    �`4�����i��� �n�!݁!�A� `�:�ԪH#��v	����C&#M� � ��F��4� Ӹ    b`p�waѐ� ;��:���i�Լ���<W�͓������C�� ;�3���&��n���N]۽��×]�꽷 7�    �q���w[�ݝz9�so{t�ΆY�<�9v��u�]�;�����<�l�u���s�W����{��2̠�zn·v;�������\ zw�     �^�6H�Ed� ������gT���noOO{���A�ݞ�� pwz{�9/u�Os�z��Y�G��v�7� ��  ��`�2t�����=�҂��\�JS K0h�;� 3� ��+p��=h{�u@ S&�S��\��ww m`zw��p �P�@hwwU
�R��� �      v򞔧�~�� �S�@ ��  i�$�*F	�` 44` �z����"L�1 �`"{JI�2��� ���  ?I�b����6�  �`@� D�@RH�d�i4�$�	���O)�f)��>����䟟���?Mw������DDC���8UTC�Q���?�C
""2)X������P��$�Aُ0"* �$AQa	�Z�Y�{#>n��k��ܽ0�.w�A#0ʚ�0I m@̐Ȩ��P�`�Iő�g�X��`�I /K#�c D�
 .��K*s�P @Q$���!  ^Yd�� 耞�� �����*�耞��� �z z ��z �� '� �� �� �b !����� ��� ��� �� �*���z �z*�� � �'��� ��z � �
z ������	耩� z*���
����J!?��
/ԟ����!��zϣ���/L}�,�0iN*nO�k'88MdrݩI���
B�8��#%�v��cj����	.����D�#D@���0U��3��d���eD�����D1LԀN.��(R@hnc�e�EV���Y�ɞ��kZ��
aQ�ʹ	 ]S*���/,�(�($
�	�Ql��
�PJ�J�+��3	��)!0#7�e%b��ꩾ����&2d@�v\#�׆2H)����I�2�fN�^�ր& $	)Y�*����R 0D��bGn�h�9W�{w-HDN�o9�	�K�"�a������j��"�Kt�&����ǜ�Lݧ�+��	a��ԋ��1PU��
r�lk
�g�Y����@�A�@���e+L�pQ�{y$�6bnT�McL�B�2�@�B��( D�D�z�q�t�h�6*,dA:N��ܤ)`C0i��-���X�gE������!B4PB8��V$+��(����YXJn�ā
00�c0ԗ��Qj��%<ͷ��j�4^HK�
�)`�6��;*�ˤg2h*G
Jh�;�� ��`�A�H�t�,�Ճ*��U��,�&��(��f�pY�&hY�lT0ڵDշ@c۷�T,���EU�z��,s��#X/3V`d�Qε�q���U�R��4����� İ�cN*��0Yw#(�B��B-��U�i���"��r0�
�NhI���J��10�! ITjVcY�gT�v	5���联#C��QP�)e��$i��

 �B1e$h�Qd(�+(!QhX�D"A)�2��J0Xe��c�M�l��f��!�����$�V�<��f`����^<S8e��;�&�ĵ���EbbF0�`�8��p�1�B%8�K��YU��d	@�$�&J�h��"�N�e+���2�!C��o$&	�X0FM̹ɒg��������nf���H0%I�B��F�`�sV
��f4��`��S�5Lˬ5�a�@Ҫy��q+��3� ʛ�S3gkD�"I���\а���%UI�:Qݠ�ԓKY�����a��dP�U�MAl@$K ʃ*���ʨ���+J�0��D��+��oZ�I*�PJ	E�d��2�B�#R�R@�#(�0�4��(���0�aQ�e$�$)p�
0�s2c���j��$�A�h��"@b
'	�T��'JW���LI �˹�0-T��J��v�!RjC�`�P%2��Xɔ��UJ�+D�@�����E�*̚�E�TD!%�\��W`ԅO7K�s�E�b$P���ɖ��F�
�v��s{ @��[�8�[�!X�*���䡵�.��$�Z�̰�vuCy�oF.�Y�4h�@��ۓF�lٶ�#@Dac �
�@�� b�0G�3�ݖ��ҥZ�(��BI��{kX��3�p�޴)֎���X��^R7*x�-�KXP�� yx�0f4
41�!C(!Jz�,�� ��0p�
@"��A�B�!
pJ,͓Y,roT않lɧz��%�B,e�˖�V��R@����F�p٠���a.��8rjo%��.9�I!���&]stt�z	Xɣ,
�yX��e]���m�pe]�%X��25
�d�!p�����
%l71!�v�-Ƀ�#NS�:	�����Ȓ]I �I:o@:%!v����M%Q(�R_8�A�����!	H�&j]��j�p�3�-[�˩���!�d ��5N���vm�@vX���|LD�I�& ��nT�H�$�f� 8�0��˚�e�4S%��3���E��&�4���z(j�p��ٳ)�Y���`���2��u��"����Z�I�(���r%V��i4��r������)u�fofBB;Ko��N��V2S��' ʃ����QPB��޻�8� �4 ����0$ʛ��9�o�h��^��R­$��x�f�2�"�U�5'@���;[z ���'+sdPk.��2��	7Qb�6�]0����RHB�D(���1L`I��LQ��Ce�Ix��C%�#�D��T(��,"�U��JY![�ʹq�F+�Bˊ��5����H�	s�/�����ʡ�6��xލ��v���`��"A5À 2`�D/�Ą�AL�, $*[��vQ�Q�fg5C�\rQ	�İ�ģW�**��ڧ�(ͧ"�L�\�f�r�5�	*�2��؅����1��n���m�+�4fۙ�H�]j�
;]�4p � ʀt.0i �#E��0ƺd*[��W�	�1�,1*&h �7;Z̓!K
��no)�:"{N٫��6o����u`3T��gi란6�ڜg�; RΝ�f��`�%.u��j�� �0 ���#R�`�T��S����w"qPb$'*���'4N������'�2,]n�j��4;���`�PD+A�H�$ȻtD�� F�\�TⰄ�Ͳ0dp����b�HN4��Lٶ�y��p7�K�wy�1p*�TSU
V+�U	�\���"ev��+����4vp��Q(�d��c��8C�ƣ4�L�c��х�0��H�=!#
(:�^3}`K��0D�u4��(�)�4S�����^lј���00�(:
fm��#P	g	�vC����bՙ�tF�\�eK�1�9VH�F�ŵb�a97B�ح �Dl�h��&U��i(ɳY��.�2��tC��&�()���ܚ��/V�o�j_9��s��1%(^)���x��wr��X2�]�,��f�ͣy����aq�+�Pa
�+jQL��Ĭ2�0�(pE�PJ+�Sx�odـ�b��p���F&aI���`���0(°�B�°ƃ4I ��1(�ą0�ā!+w�e]���'T�V�]4��U�E`��e�����PM���D�/{ Fn���@�S����!�+R&cF%8�4�,��QU��� �J`���횃2�B�t��� �D�%'j�b����=��S3�B�A%���bsL���1�b%�0��B�bQ�(!+zeg!��Q�%b�)�� ��b5��)*��2d�f�pY2L�K�a D0�JKp�5�HVȸ6�$ՑѪ]2��:�@�N]ڝ�%�Q��T�Neqt|�R��	CU�B,I�F5.�V���Uۄ�òk�^!!Atb�vT	$m Pp`�䌦T�%`�.��,�P0H$
�A��	Q��
�B@�4�0���A F�\�J@`�c$i�LF	�2i�P���b�8��[�cW�01�ݎܯ�O�����w@�z���b��v[
�vL1�i`��T"�x���N��*�P�QYXLb	�(:(c����8T��0Y5F�X�ʃ
�u�4�rlh�@1(0	"�l+�̮N&nA�,�$�e`ۭȁ"	M�X%�*AĨ4��J$"����1BL V
E�K�x!L!,Ġ��(d1E,*�y�jca��9�U;4�1��5���U��tpl��u�<]�kV6��Y�����t�.�;k8X��RRu�]��j��d0�q+�^�����l>^�lh����e��v2[���Z�l5{�������9�%D?��O���i�S6����00&��������w�N�΀��.������  8H-� �  ���  �Lh�`                                             �!�                                                                             z@                                                                            �z                                         ��s���'u���;��r=�c���������w0�dgvh���b�`V�j�UwD��p[���J�m���s��B0��n�����`�W"�%5��Uv���y�v��uʠw��_'ݪ��Br�e�J�A��E��s�u�ۮ��h��d7 �!���[�GJ<!%�Z{���Ohq�V4��gtu=���:b��+�gt'=����2��Va���k1l�0�ꎪm�x�;��K���k�}�}���Zn�8v�Z��V�[����+B���' 5P`7���7A�]5$q�c(���Zt5+��8H��ʵ���V�Ь�ְ'E��9h�:�VK��zV��S�d0��JU K� ��;*�WU�����;۶�vbe�[�Ǘ�S��Νo\'A�A��z�=u��ێ��%�h;ǢN�Pۖ�^4�x�&�ީ�/2����� �m� [��H�&����Bj���vS�5AzI(�YР�ޡfL7��=-��m��mmʹ�pi��D�G�⌬���]�j���,�J�$ �r��m��m �L$ �qV�U�^Z�����ݭ��2�n�l��m"T�Ā��kNF��iltZ���է�Wf��V�"�5�i(���@X��-;��`8y�n�h�-���H�^�m�e۱�<f��粜;!(u-"3ˁ)W#n�9Ƚ�_�J��Bk���U<�Y[�1 l
�]UQ���n�j#��Wr�Ƹx�@����t����K�麎'm˹�S���^.��oWo-y��Jm���g5/-cJ�/��ۢ���s���p�θK$MS�����Cu���E2�e�IÃ/p�f�;�f��1���\M���S1�N8*�)�{rTI�$�[��-�` k�����\��<D�K�Kl�ћ �seV!���F����q��XQ�6�
��i%����K���/$�:j�f͂��y���#�����g_�`1�Wk@p�󶳚�r�ԙeU��B��6����D�m�M�E�7n��[v�;q�v�bu��-�W&�e���� S��l6m� 8N�+
�5���%.�N0��]lj������UPJ��\/7[m�*�J{0t;��j���Y)�)/V���s��}�WUVq5��g��?|�U�n��fͷf��` 2r�(λu�F���х;m�!��lq��U��c�\�oEi�J�N	8m��-�Q�ɴ�f���g�K�k��I�rt��Ҽ\�V������YZ��KEp,U���m;V-�Ϯex;/,�	}�����*�h7�Plu.s;<e��<Խ��X�4��t�8�Q�Up��c��-�8vT���F�ݐ�6{�a��x�p�R��E��u��/@���5v�Wv磲 ��R�q���k4ߐ�;?p7O���Ww:�q�v�����we���3��l��ySĲ�I����@m���ōvӜ��x7g0n�
��^���ٝnmGL�\�p��j�St��:أRە^��U��[Fk��=�{b:L�n���Yx�;�����k=�"ЂMr��T�6��`��, ��G)�Cc�V�[��r�/�!��h���,]]vBv�Ȫ�VX�Z�S�UU�y�+�rh��^�ßsmP��8|�ؽ��T��i�tGn5Z7�����M � �ۦ�r��y@�2[̙�8�n��v�ז)wfq�̜�l��a��'h��籶r��q;tb�q�ZU`�ۉu�d7;����A����Gl����-F�Ǝ�x�'���l��X��l�� ��;0toSr���c�g~G[�|�OV�>�/l�U\�oL�Kҹ�G*am�V���
��*F��{d0�\��Dٗ��SrM��+�Yy�_�����P%�4��~�z���$ I��d�V�Ë�V��n轄�Ḷ�%eN�kn��SL�Y@�l�l���"@���\�[PwmMV�%��-�$ŶU��t����6vV
Y�Z�-�sm�mE�mR��0����n�P*��,��g�lm���I�m��׭ d�ݤ$v�4�'K�i0xr�ܵm��[/(���`���������$l$z@m m� qA@T�ϱ��ݻ:�&�]v1>g�[P9h-Ƨs��ز�ق�Y`���B����9l����p8Լ��� &���̂ĭ���V�ڪڷ��[ m m� 'Y{i��l�@m�ۀ�Ӧ��:<s&ٰv�l�[M� r�I%� �`�%�%��l鬝�-9m�tEUu3�V��2�`���� 	Wm@A�C�$HYF�[��Kk�6�b� $ݶ9:; 9m:��1,�I��H-�h ��a�V6�mn��F�I��[G���`:	�Y̭;�*�i��g �@UUUq�ȹ�vA��imK��Hvݭ�7��4�'<� 6�m  ��L�jj���m@]r��q&d[�r�4�Б�-�6� -��nE�b@3J����,R����'-��2���mTa�[jU���{iT����ҭWU �U��7;!]�v�W�U`��֬��ѳ�`��6[U�`[F�ۧL��4�J:��veZ�5ק�{��]���ڻ_o��"��6�n�q�������<��^3�������*��R$u�6ە�
�y��\a��(vZ,�=c&�3v*���� 6x٨b�U.��ä��c,�O@U�����m ���%���.��UG�P���J<$n:�r��l�S��������s�7\�6d��h26형�  'T�/�:����wam� m��"GA�M%f9m�[@��[5��E�%e��������ec� p]��J����^n�T:�^��	l�q�Ļsh�ۭ��`r�
�^�eeuK֩"��;R����ey��^�k��W��*� �6��!��6� ,��qt� s�&�խ�� 	JI�`��` d�Jڶ�C���l -�@  m�$h86���h���6ͷc�h 6Z ���0��,�R�U\Xqӝ����Cu�8<檪4$�&۰l�b@ШVZ�"j�ciV��%Z����ܠ[HLUU5a����r�=r����l�x�)������f���Z�g���n��a�?�����5Ք��IS�}Ks�8���Dg�$�t�:Ű�ht9��c.�*OU.*\�_����|,��D���)�X�"��PA��$�E��a���C�y					 ���������������������   9 @@@@�4>�adA���	# I�0 h�B �`�) F!:��J��.0��*�
�®0��*�
�®0��*�
�®0��*�
�®0��*�
�®0��*�
�®0��*�8p��c��8q�8 6�0��*�
�Ռc�c��} ~
'�-�'�U�G��o�	d�`����D��<�Q2��R�\��� ��F�(.ꔥ��X�T6���Hȡ�R�[ �@-S "�T�\!�h@6��"��#�6@�
�R����ր6�^(a ��P: � �z�+�A�����ݯ�t��t�N�`�Q��&^ �CN�����&���']�T\� ��9�pD8��C��b)j(J
)�
P4/ 'U61T�]D�K��*
�[A.�z��X��z*Ѕc�� ^�X��"	�0����� F@(% �E�#�[�
Tv��؃����"�H�c$#`�8@��hD6(�@�Æ��$H3"�h���h�S*؇S��N'�3* IEj����S�Q���"��e$	R�T%%�*�j�",V*�$N6fT0R�uAKG#H' �	�E!�؏A�D0�X	��� " ��C����\���$�I$�I$� >�����b�C4"�"���ZBj���)�  @� ��˕X�`.b���G�q�����x�c�۳<�@24��b�5sl���Jh�l���        �`              �               �`       ���:N�O�m��g]a�F�xt�s�n݇mՌl�zl�۳`l�;����Nt���v���̛=��mԹ���V�k���l^�Qٓr��vn�R6����q۵n��ܯ�E��;�3	�UJ�@�9+eIݽ�q�p孮ϓ���,l���;��fr�n��k��g:+����s��9�@������d��һt��@c�՞����g�mO�ṄX��Y��	��N�@F=8լS�qh;Y��fݍ�c�$�q�y	�^Ǯ|rq�RQs��qo�'vyik=�{��ŷnk{-��藎j��7�.ҽ��ã��T4��*;����k�қ�헚�=��qp�6nz6[�80
.��lV�(�Q�u���;sW��[�n�=;����v��=�oti^�L��A����˝�g��ܱ	���m��h�d���;���"�l�$�ru��D��S�NF�zکڰ�T��Ԯ�I�� @��TJM�r+�l�UԖvE�5��WU	N�<M=��QK#d�1Zw��L�Mq�N���W��V�vԶ�!�g���s�]�;�El���k�6���;����sضvʘ����U؆۞5��ˌ�YY�Z���I�B����r(@�ۑ����R�l�1c=���V82�;[�X�ջ[;�i7[D/\��Ρ9�����ٶ�F����wx����!�t�`�Q">G�eH�tT��_!�6 �-��U0�p �ǚ�^�Wwwwwwx�0  l  l �k5cR��Y���Ib]��dpͦ�;�!@A-u杷(�3h	\�ۄ8�K<j���rrW.�3����5;;�&;n��b��U� ]s�r�q��J�Mtr����p<�\��	�TN�82\�
�R�q�]`��.���F���J������'���{��8;<v]����}�+~�^r��@�"�����2�䲐m�.*���y��O1��N77ÃD��T�e�Ӛ��+u�:�S���7qh-)A�[R��y���}�U��7I�[����C���_s��D���,E�~ 	䳲tZ�b���e!��S�:�J ;.�FSR�I�e�4�sb��X��q��y��H12����}�Y&�D!�.�vg�=�r��-���]�I�(�l
��6�X�y�1���<N��L&ZMP���}�U�Ev�2�%'%��m8��b��X��q� g���� ��։-�I�4�d��u�twXI䇧k�f2%�4SRԩL�j�o ���qW��f��)��hJL
��6�\U�1W�z @#=�8�-�2ٙt=����q�`Ez�d�9�5��û�JJS��e�}�]��k{�:��5!�)&Rt35 �5�^늾�=ߛ� �V�I�ug�ie-�%���'R](��WK��@ a�!�幔D����cou�_sx�xs:L��L&ZMP����D#w�cw�"�5���2�䲓�⯸8�8�� ��������r䴥��d��/����f4&���`�Ai��39p,%)��jRL
��*�X��y��@<�Ͷ�m�2�2L�,II�nb���vV�
{T��
&GL�r�LlI��ʎ�=Ŋ�C�@R/��x�pR���,̷~�9:���c�5�=}ǚ�ؙE�������C���fs���d&\��2��DD o��;;�U����ÜN��L6KI7Q���81w�ٮp�p~fڀ        ԍ�b��N�ŵ]�^:n;>�Ջ�!���5Qi��Ǫ�۩��;�� �ںz��e7L�N�O�^;U�[�t�1��k=Uw<�ܦ��)���Ɲ,qcӻ\���,�\9A]Z�Z�ض�g!��Zk뻻�w��= �Ω���1[OWi$ڱgZolk�3�[!�r�d�6��<����U���ך�sxr-��-)nT���z G�<]�{̑W�c3V�Ҕ�e�JS�y���}�U�Fv�����$ؓ���so6�;���O4��n�R���,i�_s�����Ǭ�?{�;����߸ ;����c�\��V�ӷ8�q�s��
C��@Z-����2����	�X�f�DD/}���j�	�(�����r��!(`JJi�0Y@HH]� c�$��ʪj3�pQ",un;=�ǣ3XdV��<�RbS-��g����]��k��Q�%'%�N\� �o}�39 ��,W�C�����[Q�e���
��b�����Ɖ>~| v��]����2�O[&�=v�.b�8C��e�J[�Ԥ���b�5�gsz��Ѥ��a��ɗC;��gsz�w���FP��)˙�⳹��Pd@ 舌��+�\u��Ȇ��LI�����+�\Vw8��BeJ,"�c�E���s��sz�����m��S%08�u����Չ�[aA:�][����}|g�D�zu-��g��
��2�X�<���f\���	�Li��@���gs��wgÄ�[Q�e���w��vk���75h-)a��)0+;���pk7�I�@�P��X�r��3��L�^$�ʫ�eб��<""��4/9W�b���m��;�]����u�WE�����L�r���*Δ%&�r�e���b�P}�Wf���+�	�%0e6(^r�u�����+I�rh��-��s��+7������RLKr�j�����6�]�r*�%�˒��!&�N+7���`^w72u�>s�y�߾y��M�         ���j�b��x�x��+���v,�lƻ%�θ5�;���&��Zd�N��"�y\�U������^�.��/Hxp�yjûe�]K��mIm���Սd$�nݻ��0�q��]��%��k�[��ܖeYM��^�m�5o������{ݺ>~���g�wi��$��gOG&�Ώ���o��9O]<���neJfe���^�����nj�ZR�.[FS��ޡ&����@vѤ�`���dˡ���Vo?�f�/=�x�N�BRa��̷��6�W��vk��ҹ�)K%Jn�f�^�ۮ+7�7��| �����E�E��� �δb����x�`�o�܄!8E����c75�f���D=�P$g9�I�n[MP�w;�*p����`A��9�v��x뜱y�̹)&�R�i�f�
����c;5�����-��)��C�P{�gf���Lnj�Zi6K�є���c75�f�x��D`�3ܹ��m��@&ܙ
D�c���]�۞��[�cp�1x���mI|���G:�Iw������f���}�_L��
L4ә����m��������{��!2R�J��o .�^���$�Km��m��ww�QLH��� �p�A��(T�������N��&��V�%5��T.�2dbZe�G5̆�y�h�3,�LP�Mb�C,��0�() g���Q����&q�Ȟ>@��4��3�l��2�F	�A�$D����l+ʚe;�u��BH�,�<b��%���`F	M����=�}3�x#�A�y��V�� h7YUQ�Q(LX��HN��v� �7D"U3�@�oJņB�	Wx1��L��(��q��\��������~���AM] �B$ �dA~��PH"ڤA�Q�uD2#H�٥-��s�����5�L�e�)6�s����<�� ��G�%K	�  �M�߻�/{Ŋ�@;���%Ͷ۫�����5̃�qXU����%t�/#���딚2Ri����+qA5}��(g��ww��D��A32�_j�u��������˃��be���`f��/s]s|�n /�F�Z%�&[&S����Q}�b�0���@�I�|��4�] 6 ����'��I��re������P��x���^m��m�"AR��&_��)�غ�L7f.$�pr�5�$�2��2oZvI�v�������*���^��_�!�BQ����*�X�s��f�+\�a�[MP��qY��f������JI4B��Nguw�}�B�-q��84HA8-�Aн��{�f��o8��1����1~���Iӯv���ϵ�}`       UU�vt�zǛ�::5 G1\�v9�.�v�ob�:�IH��뎱�x5��݃:��4؞�_�\�����f8�f����Sg�Wb��:���!�;`�6�J�D�=�7�ݡ����デJ�R�^Y���j�pJ���A�e9RP�p��K��p �@������ʄ�5M�WD�%�b;sá��l���t�s,�-��$�%�2��y�b�5�7����{8p.T��l�u��+7����^{�x�I��I���2�Vo���_k}�:�J�Bd��R���"�O��y�����ߜV��!2�bQ���y�  ���5�����m��m�[)m��	�]뛈��&�] nfq��8�][�7]%����}�V��#��y�ޟ���cn*��s����߅(�c��/�����#����IN
2���s_��qy�1���r�L%�2���fw8��1�g�@mo�2�-�ˠs=�}�V��5�� ��S�m��wtnm����쵸99�twD8�\.�����s�ibe���1[�Vkf��gi\�L�e�A'B��W�C3��^����&SwSX�>C�����;��ċm)L�G�A�,0��"��Ej�B,$&z� 3��}��|�������h��3>�y�V�A�o1���.T�.�M8��1���`�o:���GD�?/�m��ff\���QF�ns�cH�����0�LHl���@QI�B�3+����f����y�b����JY,9sEX{|��S�s����~^湌E!����r��m$�.�XEw�����Ɉ�o1�'B$�e���7��/���,�~�<'E"��ҊxP�!�M~�G��ǚh9)�)&�_ro5���y� �O.m��m��)4ҐKI���q����m��e�f�3ʞ�Nzi2{���������Y��iJM��m������/y��c3'�\�I��M8��b�PY�U���ÃP�N&L��_rE^�.�X�DA��1�˃I)	��2���1^� ���s����"�N��������         	�n�I�!�X����7C��� ��v3]	p����h5�0�Ӷ� vx�.�l���0�z����W�r���i��'\��P�n�s�X��N�n�����77c���;v������q��O<U���cC֠��i�Z��k�מy��w�q��� <�0m!�l�+YBUqO.93�:iv�P�Fp�����[�hﰟ�7}�B���X�'B	l�(L�}�V��5����x�����i$��}�D��Vr}͑W�qz3\�mIS)��" ��1���<�?D@�3ޠ3��C	'%KM��s�E�z�� +ٮ+ۭ��m�!#!�I9?BY���8��E�Ta]��8�uk���Yܐͷ~~�~�}�Y�3=�;{���A6DəT5������I��9��)��!T@�Fc2 ( � E�Ulg��qW�? v�$�0×3,�y���8y�1y��h�Z�(0�̺� g����{�3��w�Ý=%����̠���菄f��7�z���j+3�M��m�ɖ���\��Ydt9�u�q˃.�o�������3*��~���^���~� ��y���ri���M�^�~'7�^{�U�+N�q��I�*ST=��⯹��D�@ `0<��� F����`�7?jל�^O�!����m== ������k�o\u���Aۑ2e���� 
��Gټ����75��,�K��2r/<ʨܓY�nٸ�l&[��ww�>�5)).L�s2��"�ޡټ�}� 
���g�el̺���/;�^j���@ ��OI@�,72fS����x�} 9�y����_q�m$�̐�t< ���y�^k����@�HU,�lT�q����9��l2��M��o1� ��q��@�y�m��m�e�-�.O�4�k@uB����7��d��N���  �p��@�\ʔ��{�{���!�� @�����ʔ䲛m�y��DD7���o1��|  ����A6�$f]
�����" >����+3[JJY2��ˏ�@WΞ�g��[�|��|>*)��!ϝ���#(0�s2��y�� G� Dn�鱛˻���㿥޻�w��/��m�� l�1VW�"IBGh\�>�T(0� d�bQFB��h����C�� L����"Y���Ǧ
�#0����Ą�)UF�P,a	BA��@"I!$�b�h+.�C�l�C��XF�Q\�p^CF��q6[
���`,�p�7L3[�K��3Z��B����%g&GFv�9�B��Q�$)��%�p$ ,��	(��j`���n��HuZ�j0�B�1�1aK%�Rd֪֪�+��BI$�V��&	#7G;���Ԯ�R�J�>k`   �@                                           ]�;nI-Vذ���А`}�Oj��Z�ŸL�^��n��	���綛��r��ϵ/:n:��q�״c�	�B1�A�{l��ֻۤjQy�u+�2�M�Uk�q�Whziy�"��i�Ү��	�IۂҾ�<��
󭮊�.n=�t���ٶ��M�9�r��v�ڌvͽ����t���������68�m�5��6�����[�9�r��$Lo����i� �$x��9���b"�Z��yf3��u.�X���d��+�klA��������v�{��*����{r��0J�8,�O�l.�B,�=�It;j5�/k��a8����Q�ŹEK,˰Onض17m[J���\t���d�8�C�;g����wn���i�6�MۧQ�����nʩ؛f�-��G83c]�(�+���iv�ٌ����6�{9�!��e2��*]�p��1j��3۶�k��y�Ve4nCQ�$)�n�mk[���I�!v�Vv��+�kiI�!64lI��2L�r)۵�@X��Aʋ�p.4��1�y�ݻ!��y��+�#vK��]�����m`��X�g��xM���X�8j��tE�4���v1p��;V�.�GgcFq�}l�Ѳm�W3��Q/��_.�k<���#�v-�Q6��ۛ��ZYld��)�G[��2r:�,%V$�����e�P-�:�Q�:^*�IH)����U4��#�U�8��m^������{9�~�t���        ��~��竽�X��y��qs=�Y�+��[8��z٭�&�'njõ��Ϸj��w)�؈�4��vx�2O&�ۧ�nN���u��M����{K7`S�u�LJ͸ ۓH��y�&�v7�����:�;}ٷiŠ�1Mg.�8^��֬I�6��"�1�gWwwwwwp�`m�q��u�OE�e��.�,s�c��U���w�(����Y�2�}�~b���=��=���m �ܩIм�=��cټ��s�Fp�9%�h%%7}=�2�C�G� 
Y�zX������A�+� �;"}���sx��"�y�͟K�Ri�-��c� D�`z����,f��m��bX)��%2�e�M��&�.��1ۥ�Z��p4R1舀�Ph �r2Տoy�׼Ǉf�|  �o�c��x2Ҕ�1.�>k����HP�I$@�-QAQ�R�c����w��~�z�� #~�x�ҙA�-�ˡ�{�}��� ={�_�T�$Ȗ�ffe8D7��+3�ٽC�� ϻ�o�'�Yrl�Mо��@��3��={������t��*����^.cT�a�G��X���JS���T� ���(�gy���,�羈�� X�r8���4J9M4�g�y� �2}΍��={��" ��r��jKh6�$^{������ ���b�7�j�9�;�å��MT�j���@�7�P���k:  No�t}�^��&�s(�CD@���o;������m���ɐ�̆�+�;ud5�R������D���{����P����;����*�D@�� {P�O)�I�e�3)�^y�""��=��_�_D@�=�=�Yrl�M��ro��"{y�����oB�B�&Xh%-� DO��o�����Y���V�E�6�P�p����;8s�/`���������@���X����b����m�YX�Qd[�.y�ՍY�w��:�^G����{����̹s)�<sy��� ��B���w�<D��h��B�iG��p�{�f��y���{�W	))JX�����b�5� y��&���$��[&Rs3.����E����:" >��3��ye9��S2�U���" �������\~ T �#|'�'�m��m��     
���76��8g��� \�9���a���	Z��{[<h�L��h�e���m6��kOn^uȯkPk�;��5k���SHk��|�G�&5���6�+��U��o[E�e�.����t+�r��ld�������RC�ԖRDIBe!�#` �".�� N�Y�Y���9�xn��v�aqA�J]�w{�$ɠܹ�L���}����~�~� "�G�_�Be0�JS`_�����M�y��C@ zt�qT�a�I�3����| A��{y�^x�\��n\�m�����^sED��"��Q��"Jp�hP����  b _��}ި����3��m��&H�S�R՚95M��L#��D�6v�)&��@T�RR�d��P�V���ި�(nw8����"�aJ��y9����Ӆ:�)�x>*=#����Cw��k��s~^S,)�,�3-�o�b�Tp���vO��h�@�nT�-�j]��^���8 �{�_�Be0�	Jl^���3W���������� Y��N�<���X��6;"�2�N8S4g��D9BL�D�����8��b�P� �^�s}��L��̦�Vg��> ����c���zw{��A�n��c8��ֹ/��+F! � H�
3�x��v(&���>��P���ҙ&e�� ���1}��<Ǡ���{;�r�L0�92�_��x@���y���qB�}���u���K&�y��-�t�԰ ]p��Rp<��B��R˙��y�/1E��D��y�}����K2ۖ����z �oP�o8���D� "Fxyzh��)M�����6�  �o΍� 77Ǥ9Re�D�b�;�}�[�ι���ք����f{�P��˒�NCR�xx����������"7O����m�$�3-���ɹ��ι����V.u5g�v������?7}Ź��m2�o|���b��~ M���I�]T�
9�@{{Ϣ����*��"@�r"dϱ�53)Ä�̩qA��U ^pL���wz�~��2zp���e7)�$�y���MR]�8aK}���P�1$چ���#nf���� ��I�oUM�$� (��8Q���n���@        n�f.W�^���N�pc�����ȩm9y�;E��^�%���*�/ll{c\v��i^�E���]�d����۶��ON���+�e�uI�ι�Vl���[k�����O)͔�y�]:5�㋱TN��7�Nۓ�}��k�������)�{ }_'�ޘ��맭I)�e���"�Y��a���wv.������� ��
�]P}��r)	w�P�=zb��%��\�u�6���^�����`m��hh��#������a}�q�q-�p���U�^�BdL�C�Jf�b"!z�������������2O����I���1@g9�mE\��w/;�^��n|��|��KM���&׶�9ԮN��'8�mK�J�#�&X53)��)hN:j^�ڠ^���3��")�8`wg%,��i̱����&��_��7ꀒ��«�U0�nQ	+ �(�5��(��u��XH+��k�ə&�v˒k��sՎr">Y���ӗ-C����p��r˟H+�E���d��~b�<9��R�S-�]3 D?w�2Nv�Q=3��ɠD}�$����e��s���r#������8e���'�:Ͽ��^���؝�HƳvq�]9q˖���#�T�nWD
i¢�,2ԦݒNo��n=H6ۍ�Dr"�wo"��بL��r	Lѷ3s�x�[� ��O�#���FKfe2eKjRM����$�oU?W$�I-m��m��b���l��dg��$���&IM�љ%Q���V��6ޙB���
d1�&-e�0BQCA:�Ue�ń
4��VH	! �F@(#K�Йb�u�DL�@�#�\�V�g	&shg��UE)Q�*�a!DaEB�b�q��o{P�o{���$�9�ي&�)zf�Rb�Ĩ�f��F6�H1eF�P�D��SQ*@�d>���(�E��t,ԋ	�� ڇ��xiZ�@"5��1(r�=~���6��"9��>b���,s��`�̩p%-	�r#���� z�X~p��[�dܥp-�ƒn�;��9ܺ����I{o*����z �9 ��ݣ��ծc����v�g�u��ގ
�Hm4���2���|`_��	�f�� ��I��2vg|<�)�d��q@}x���� w�0�
�C���q ���r��q�q�/sj����G�. ���é��y�I���Q�dȖjSn��3��d��,2O�Xd� hA�����g���0��猕p�p� ��|���
�����)�����A�����m��m�D�"ZW�:�J�mwS�@�a1��~���Bf؈1w�m���q(�fU z�w��R�0/o(jfSp"Z��yT�d�+�����c��H��JY2�Li�2�ײ��ۆg9�Ko0+�yށ�46E�A0�mQ?D} B���$���'f��� z��W7��[h��q@m��}��'fg�L�[�2O�� ��N�߽���'�%��m@        ��Z���q��tޱ�(6�/%���.��vsM�����[�����97���nF��R�N{�����m��:��V,��lf�v�aV�pm��q+T�����E-m�Om�Q�zv������(�X��7k��3��jw?:8lG����;���~~���ؐ��=��h�s����A�Q��n�����;������S��9�1��������`U�p��[�=��Q,!,2Ԧ�M�J~�H���;�Q@wo*���H�݊�șp� �n����o��9�o""g�f� ^�,�[��KcI8��⿷{�6��r�y]�T0/o(jfS`�D�N(��P��٠;�p��s۞�ԓ����@%�5�Ie:��][��{3�=��Ӊ��zz�t]�t���z�O>����0;��}Ϲ����T�>��4�d�.^3=U�zYt}�l2O�48$�F���#��??�2M{;��$珥m| 
I�9pA�-J�m�$��a�osj�@ } ����9�a�M��Hr���.SB�N���'y2Mb�N�M�jw�4'���m�oe��c-�ۏ�]��@�r9v�[m�ۄ�SZ�����-��-�:6���<�b����}�8n�v	����Ľ�*�{ۊ���f���Ls)KI�4��z��\0=�ʠ����=�H����nfN8q�'9�gک&��\���|�@ ;"A��DX/ξ�D������L�&e���'�>�,ts0=�q����nv�պ���$ۚ����eC���P�e�Q~I�m��ov.HB#��Ѻ�3�ͱ���ku�d�J78yo=:G"m�bE�`wٕ@������f�`���ܹ`Թ��z~ʭ�)';ɒo7�Q'=�?d�wD��C�m��e�^�Ȉ��sە}�N�_={��K�r	L�lD+ܨa9��$߳j��#��"����;��e�s
����|`}�^w�{rI���Owπ ۸Λ���9culذ=��8ۇv'�VG�%o��������v�1{�T��`U���9Ȉ��p�����)�,�!�$��O� ��s�\2��ו[�&O����i&ؓnh�\0;v�߽T�Ɇ}>��q0��6�y�v�����������a�N���6[-�K��(}yT�^͚�n�p���LpL� ؐb �#����<�;Νm��         <˺��gU�����3X#Mm�i��u!њ�-���1N��h�����27Su�/\�[f;=`C{��q�w��I����lƫf���l���f�#�k#�³P�<�B�<�A��3���-c��ڵ�<�i���<y��w�կ�� �f�Zķ\u˧t�	��b�n3t�������~wƹ��ږ� _ߒ����p���U~��CP��S4r�]o#��x�� ���8�ܼ�ҙ"X6�)�X��=����6X�NH���9�S,$lI��Y����^͖}�mI� @� ��Xd�ߟ�ρ(&�X�M����B��%�ێ�]PO��� O']f�K^^$�H���؊9�mڜu�7l�Ȃdh�cbR�I�=�:C9��I�oW� � 1w�&I�]��	�c*���2M���O*�B�s9��?u�l�;�qtD$��!��SS.[�Pj��U��6Y�������|sUL�
[(�-�D� ig|�79�P��������/6)D����wJJ�a�~ ��D���}rI��>�~~M�� :K:�Mv].���II�v�N.BM���$�3)�#��8�S#&4)��{����u@��_�0=�wfT�	q�A{�U�s��f�ݷ�yȈ������cIL: �l�*�˟I����Ȱ�HĀD$B"�ҡ�g�����A��ĥ�&�h;��%nT08;�d��mQ$��2M��	0�����P���#����ٲ���ߞw{�_ '+$n��{.��\�5�k���Q�Յ�%)̥��s���!��T4��1�/sj�;y,Ի��W�*��I'���r�tI7���DG�@��s��y����#/>�CQ2>9�hn�`^��G�  %;�z�w�&I�ͦ�Ri�cB����9�F}U��^ﱙ>�h�ХB�3��'u����6�ٙb�9��Q'��@�n�=ێ��0;����m����I<[��7Y7�)�]V���8�x�np���Z.�R�l�*�����{�3��G)��[���ĥ�&�h�{�G8��f8�A� �j��r"=sy.%�%�m��c�I�uG܎r=�K�n@w���cd��R�(�r����#��W#�^ܨ`n^SBpܦHږ�u�ؖo0;��]۩�����>ԒI$�m��m$�I��>HB0#
%4B��(��pj#	RBF��L��Q���+Ӫ��T��k�+TXf!I���*���(�Efd�!IC�̏�FH,I�BH�0��U�Y�B3-���#@�AjH2I$p<�}��r�LJ��S�������Z�٤'�[�[                                                v�uQ���g�W��\1���c���،5oEÚrg���Hz�����=iHM��N�����;%:d���	�a=���[ ��0�R�gP���d2�,��)��g- 6$뎳�6,ՆSp�^#��ck�a��s�CcO��G5����q��ܴn�Hۺ�v����^B:�e�-֙�s�gss>Kn6�V�N���c��M��Ƒ����`�ۗ�%`�D���vS�a1�:ci����u}	���C�;�� ���kJn���(-��O:��<�rk�{'j0��=@)�9v�n�m�����fܦ����m�x�q�lq��&��.ۏ9��k�m�+�7ۭ	ؒ�.ۂ,�	�@x¦��s��]ÝĨ��{I�����
��d���;����Dg���b{7W3@=�|tWkG	�&ƎUF�yA�km�ki�n ,8ѵ=��=%�3D4��˹g����v.�I�1ۮ��;9�Y�;6�R�0�(�WP��ͲUٓ�mYWcr���	cawJI�yf��B�Wg��'a���|bw�Z�k���sq����7%F�^N�k�Z�9��:�]����rG���Ѣ��]���W,-�ʚ�x��,^+��鐀̀�js����uSevŃn�m��=m�E����]ێm����������!�GP I~s�>�*'x�I� ��}� } �`�Ӂ�W@!�G@�⒀W^e��f�$B���-���        �~����������*I�ݚC��t��D��ϲ[0\��o6��������U�͍��:5��[���\[
݇�H�M֞
�^�K�&5��v¾;�A��Z�.��mB�g�Fv3�����b7�v5=z=�����Jz'[���$&Z*L�� x�!Q�m��m�3yc�����̊���ŋ�qڹ���ul^�-���������.���ksj$^[�}�_���o9�H�KۻM�2܂�4���c	5{�D�{��$��� �#�s�rۖ�JlI�z��婢=�,
�0;��ܛ�.%)��bJ]�!/f��yQT���*#�����t�1�)lIÙ�R�k��0+�u@��'���| �lv���+a#s�6SF�K�(f�J�}�3՚�s�B�f;ܓ�߮]������"9H=�ၑȅy�|�ĦT��@'LY$f���! �� �.ɟ|�����2Nw0�L�ݼ)�8�.$�m�jW�K��|�^�0=�ʠ/ֶ*I\�|NBT���ݸ`w�uA����,�e6�'0ԤЦ(n8`lG��ހ{6Xv���~o���]6��i�ݢ�����{6�}sn����e�R��ʖ�MKq@{ٕ@��]��9vB��};&�%3#�4&�$�ܟ�""����B�9��d�����	G�>��l��CNhn�`Uی���EO(�N��Ư�s��I��>c�̓���8�s0�n(>�+ݨ`{ٕA�{6&Z�8`�5	˙M&��V$]��ZG��y�@{u��o��v�n�������Xv��P�n�:%mq���MJI�ZI�h�oy2}.��Q>��c@���Py�Hj�BTL��q�t��َ�ڠ��)%�mJND�H�8�=��]��H�l�;�p����$����ؓ���#��������.O���%���G�L�R����>T*0JB�Tk�Ϡ���3�u��9��x)��a�&Zu�$�~K�n�{q��ܪJ#�{��m�g�u�Ώ#GK�"��Yq�xnn�OX0��o�_}|��7)&�zuzL�f8`Wv�$��<�>�q}h�d0�JD�łN�F�e��Po����1/]��I�I�Թ���ڠf�>�G#y3���\2��3)��Lˉ�m���\jGrp�A�c�}�T�����ა�3@v�j^�p��*����a�����<�N�:��P         �XDt�>v���u��5\Oku�n�x�:Xή{n0�[ X�9��M��uɑ��������Ϋn|Dvn�nK\\"�c��CZ�\���,U�.s�Xח�LX�m��ӕ�z��U�ѻ�+�!�ڤ-�)5��w�;������ �v�zZ�^#T=���:'�-��f�c���������L�J�^�`wٔ���9�Gd/g}�a$�I�'��� ��K$�-,�}�?��#�/#�RNK,�2���`_��z8����=�eP�9��������x�o׹Q@_�j��r��f��(q-ȒmP��F8`o}yއR�l�1^&���m��m�������nH�:۝�p+�m<o6ذ�w���%.c����U {6X�)�073�˕)&h$ۢI���G�P�>���g�+7RO��T(�y�*�����ɹ�P��h`�%LM{?ݸ`W~��Խ�,�y�Ȝ���sg>���#׻W�����cҀ����rCa)�'}�U�ٚ���I??><I�>��� wd;[m9���m����-$pF��£q�a�]�_m������M�H=��H;�ʠ/��ŵ2ፍ9�I�n��cC�9	�p��*�;{/yL�q��ء�%��n:}�YrL뜬�`��Dd=A�XF%@�#@�RQ"� �C�B���>x{�2~��h2I�;>dL��ZR�Pg�v;@ݖz�0�9�eCs2�jR�p�3-�>H�},
���E��
��Qػs���m�Nq�l��p�"���F�7���{:�Ć�lYR���v�07���\���,�y��L9�L�bFn8t���aT�����Ȅ�m���TL�CbN(^�P�%�^�e�0/ѷ��*$S.	r�)~ ��`W���6�9Ka�I��R�	`A�Ҡ�z��f�'7�Ȱ�E�I�To0>��}���@�������.�W�:Wnis/Jf�Rh竳�	�N2�(Cnhi7#b��/�[qZ�{��eQԅ�ױ��p�=�c!9pۉi���ܪ ��+��ܷ菢d�wi��$��-��/~�RM�f�{�p��*��^ГPKd(RJ���{6����2M_����@9�&I����f[ID�N(n>07������K�6C$ˠ$��@X�EI�B��!b$@�Y������]�        ��S���]�mU,�p=�ۢ��K��Y�k�V�eg�<��@�6�%�n޹��������X��&j�hZӷB�<műb]�����l:Wt�i�Od��: Дp�m�v���y�`�\���F�k��Л�����޻ݻ�w���� [{�:u�s[��mo7Tfm���:w=�JlR��I�ˁ&ĜX�ڠ�K$�k�N���7���FRpSLLˠ��?�����n8`Wv��G��8c�nfbIm���p��ۆwn����#.o$lLj%��p‽�w�5@���yP�=vk!9m�M�P��Po%�^��I=w��ߠT�l��n�s����������N$�xq+y:��L�ვ-��{7]����nܺ�՗���HI�%F1�&7�d΃1D⇇��9=�Y��;��@͗�/3(����Yq@n}�E�fU�H�},�B]�p��-�!8��ʙqX�w�T��`Uۆsb&���^�vM��p���.����?L�� Do�P�I�y�I��j�= D~���� ����%�9Vl��^{Wb���­oj6.n�Lp�lS-�2��@��;v������P���@Z��Y	�%��n(}���Ps"Xv�W�cԦ�)�hQ39��D�R�yQ�����33?�KͶ�I$�S�(�?,G���S���(���T���D�UUFF�ɑ�8�k���\%�V"H�\�]�¥B$���LI�%0��� @�� �!��yL�D�(Pƭ����ŭ��]4m�J%�h��0B^��0Zicc0a��qX*���Fet+��̬LpR�4:�o}��׸�1;�s۶��=�7�e�p-]&0���KK�����A$�H�(�U��$d�)aI
X�B�R@�
B��H� c
Q(IA
0�
eL&+J��2�l� �q���3 ��"��P�ɖj`�R�
�)�BA���`���c���������v}v����}ݸ��v�8���`�F%�L�h)��*�5
�*��*QR��*p<��p��P�+�����W/��Q�� ڿx��G��ס����^0��&~Ϙd��w[jR�a��M�'��8��|K����0+�u@_��%-�E��R�oy�I�7�
$�{����Ϲ$�=��� ���n����ʝi6NW,�"WJr�,�鶤�H�3���+�I�������fU%��v���s}t!8��8�;�ʯ�9H=�,�8`wm���*$S)�R��)t��`.W����r�3�zr�Řbإ�S.���v������8r8	 11 U*��;;��"C	����P�0;ۺ�fK��?��?D_���� <[�α�/e�j��AB���[�3]�Fx���r�\�jc�n��Ps"Xv�Ynwt�NFf[t��`W����?�;�ʯ�#������>8RL���p���R{���e�Ww@�m��ЦJ���{2���������4`_הBM
I.q@{�e}��e�ܜ�p�";�p���U��`�(�Q*V��V!}������ŀ       z��N��s:���� �]pf[�����m�6y���);��Mȅό�v�vyͮ��/:�t k���[[���B�۝�	�a�&[���Z��t�-#{q\�.�7X���E�]��w7$˸���:��p�+��{��Sz��z�=y��Hj�y-�(^�x]V]�裕�n%L��I�M��^�Ԏ����㏣�ȊA�}�@|�MC�je���9���c�}� �d�WnKdHa�aJL�&�s�W�T} bF}������X�*e�4������z�{v]$v�w05_�49r�!9�m�RH��;s��ۨ�;�ʠ?;���� [-��*1:�"ۧEWnEե�O!\]�YS.%��L�>8S	J��;s��vᚗ�r��r9�y+��`lswj"��*��X�̓_;e�7p(���0 c� ȴ0(�Q#)�P($xDB��r��fU z�X鱁컢hP�Ip��}{�ހ{vX5S�L��E휓"I�M
]܎-��颒��L߲����u@j�1�&\�2Ӛ5/,��������tw쨠���O�~|m� wd�8�,�u9jܼR�B�l̒X{:rbR��u���>�~~�e�ڻwT�`R��^�C��@�s���������L
�p��~���R�"ZI��$���f��K(G H�<^fy~��η�fI���J��m(q2L��W��Wnܺ��K��r$�%�2��8~KW����{�y_�M�x�ٻ��m��|,mR��r�z��[��ZF��KbD6��s[�1�9�'׻T��`R��e�`w&丒fA�4Л��K���i�Yn6�dz�{ߒ+���ȉm)�-��@��_R�8`w�ePw%��ۙW�9rJR���
��Ps%��.y1�R��!T���h	D��)a
*�TjUS
QTB�&���UrCݳX��[i6�W�����H.�X���Q�8`}�G9����m�)h��;[��.���nL�l����õ˚5�%īo��,
^,`}���Q@wەX���`NR!�L���Ѵ��p����z��컎$fc�D��J�&�pƕz|0祁^���컢�K��P�eoPݖs0+m��7jR�Cp8J]jA��m#��ҿm�P{�@(�s�_/m��m�       ;]�*���'�[xzV<j66���]�r4�t<uګc�L�6���㵋��ۢtG[f3L�W[���:#F�k��;^�'���]���Z��'3�k&���Զ�櫉n��֢pk�ˀ��.tCa��8.�Q:0�v��0��o\���}�}�@-Ν�tIs�K�L�TN5�d��K�5�h�AR9-��-L��w1���8`{ە@ܘ`uw�*�'���;��i��T��d]�`��9s.P�siyU@j����p���[�%�r�\"S�Ӣ~@��y2M�8`Vۆ�D/���t�@��6Cr34�;�ᚗ��0=�ʠ�K���� �b<�����V᝽s���g�q��:���C�L���c�{wT��`W���wD	�a$�I��fUs�pCd�rd��a�ku�I�Z�J2����uIo	`z��(�8`w���1f���ʗ-���p��fTPR�;@�%4]��|!��f[���ۺ�Խ{����p��r:y�~z i��u-��n��{nc;�����5�\?�}�Je1\˔5,��mPs%�Wn��0>���
T�Ĝ˗�ܖ]�`Vۆ{�U�y�%�$6AFZTI�y�I���<C���rH�d�)$�% JH\�]�>����wwP'4'#�y��o��ڠĽ����ۺ L	%�N({r�������O\�~y���� :O25����u�v뙙:�s�<k��z�u�
��[��-z�`��*��k.������0�Cl�2�&���p��";���nU�3�y?� 7:����!�S	6�w�0;ۺ���%����^�lC���s�{T��`Uۆȸ�f�$J�+�A���x�rMk��*��a>$�\� �d�*��5.�8`/{Vwܓ�|��@�b7-�zX�r&Մ�l�s��򽜒9p9�I�	��;�p����.���{1��ʁ8�J's0;ۺ��K��0=�t@�Ba#bN(Ԯ�k�@{vX�qt������R)RĘХ�}���`w1���0>������j"bD$�T�@w1��n�]V���X��s�n������� ?��������ۘ�Dc0�X�!�$$$Bd��,T��Cأ	~Y���UL�j��lK �0���d%�dP�B۹�� BɒF$�X#�e42�*$cBH�;�`��Fh�9̪�H�"�$ 0%gH\`���D&+�a���SbT�E�haF��P�-%R6��R�fGYHG�q1���0�$��� "T`hcqb�ʈ�W ��
�K�*P2���[�������Ѧ�+1Xq�&��ͣ:j2H�����r�BB�Qx���1'oj�cc�V�	"�Y����9�J�� qX�(��Є� �A�a1��$�H$e0(!D(!L����I@�r.G��I�݃l<v���m�����v[���Ѷ����/C                                                T��7m�.�a�ŮK`զ0T��^��:
���64�Xt8���N!.��P��Zq�n8M\�Q�`�#�{ @��[�=���b��sO ە���������g��z|�6���q���ٹ�n^���s��kN�Q8��x{�㷷k�Q�w[�W���;8���"�s�h`8:��=qΞa�F6��y��a�ۄ�wb�uٴ�m��ñ[&�w)�[v'3d盭�t���͂۰�w�a�g��u�s�ع�bv͎W��vV{:�9��vw!��[�z%Ɔ�ϱ�0�v3���n�%���O �帏l�\��ͱ8S[g����ەv����2A9ۯf6�����F���:u��<ƺ�C��4<�`c�\"dNt��ף��p�"����qK0�It�S�f@ȱ-�;R+��DA�XyA�f��v��yZ�g�m���������Š&�$�u�u��2Lq.��X��ɍR7M�.|�8��2�'��P�����F,�ԥ�ݙ�"c��b�t�q�u����[����q-�p�9��sdq�[i1�Џ�(���X*�Lt,q�N�z11v�LZ�kk.��n'D�n#.����ͩyy1���	�vү�hq�}�y@���g��@��:��3���fݻc���@�Z����`��������{�ߜ����FѶ��j�J:
�R*�@$PWa���W@���D0tb�5}*���        	����궃g^uX�5�7l;G��\Bgtvj����6��uўYϱrq:�03�����&�k�]9���]J�=��Knd[�e:|m����� n�$�N��[e��O`6"���]�yչ�fny"��MFl�@�����������}�UU[�.�!�fM;5u᝶��d�ok�0DF���um�����~��]Q�${vTE.�{6X���H�@�s}�U w2X]�
F[�_��8S2�%5.] w2}H۟R�p��rꀿ[�Ȅ���}ٟn����n�������$�[r6�n�K��ၱ��כ� _�K ��`o9ߞcm��m�9a��8������A��a�L{,�%a
ݗc�u`���ڠ�K*���uw0;���(�m����N��'>�w DEG��/v^$_���ܪaf���
X�I� w2Xj�eq��nU wrX��Ɍ�������n�`Wn�;�,�r��r8�vk�K`:��q�={�@}^�f��=�,���9��۪���Z�%�r�u9}��n;\UIԐ��k��%Ғ�
ZM:$��&I5��>��P�" R_�Q@e��2�&��f�;y,�.�8`wە@ܖ��BN%��̷)*$�s�nT��� �DA����""@Tk�3�{��L�wQY2Hؓ�������$�Y�Gs%�]�*(l��%'2�e˄��w%�Uܰ+-��{r��k[m��l�
M[�����g�R�v,c��9[�-�m����b`Uۍ���o:���`uw��e�[jT����6���9��D�����;�i�>b̷5.b��ݪK۲Ϣ�mn����]Jp�e>Jj\� ��)]�e�`��q�"a���$�k�ZS"[ �)D�Y��Wn�]Ps%�_Ev�m�V�4�C�L�Z<tjk�=X��C���]�+\#�"%�ʠ;����u@%��}�-0/�tpL8��'��*�;�,
]���;�Q_$_ӳ��9Nf\�J] {�+�����r��NI��lC��i�՘�v�����D�y=��� .���-�*fS�$�q��wT��`R������        ����.��̸�wEb&�a(�;s���
��S��9��c�#�v�v5�ƽ9�s!���z���/���"s���K�����'��i��6K.��l.r	�����!�CNpc=���.Y�#k5�C[mx��v6J�k+���[� ��i�':�����GW�h�5 �5�)̥��f[�G-�x�ڠ�K�z��-�/�R�JIO��ˉtVb�W��.�W��W�$e��2�9j�ʠ<�S
Eۆwn���L��������9�@w1��wTVb`W����]�`�č�8�;�ʠ���:���0>�#���:|���xt��D�{g
�F�,�[���i�q��%Ċe�`NS��-
_@=����L
�T�}�Tu-��j��-�Qx̒�����p� H�� �H1���ʼu��ݗ$ַ��I5ܖWnK�9�R2RR�jG�\0;�ʣ�${�|��j`���s27nY@w�eP���˳6��wpp�ܼ�r)�O��˗@ܖ/Zz���ʊ
]��hۺ�m��HK��#jfD�f-t�t�v$Idr\��*�e��:�v���o�������]˪$�嚑������hR�2������G��T�d�7�x�>��7���Ip���6�����8�$$b@��!"2�c! 6�T��#����Y/���79ϕIFZ��i�K�H=���L
�p�������	��Ӊ�����L
�|`Wt���K��r�m��q�6�1��m�F"�L����7P6a���i�e�=8�m���Ѵ��̪ ��� �N$�;qd��nj\�ZG�j�� �)��`g�$��MIK��I�D�{ɒjwe�iV[���@wӁ��CmBmKsX�V�bY&�Xd��ڢpD0�2Og��9�)cR��8`w�u@̖/Zz���<fOͶ�m��8r�4-��K�Q�(��Z8�r�B[KÎ��9obضsq�ߘ/>�������Q�܈�vC�k��;:�Hr�e9hR�5L����`Vی���P�M��cj[nS�PW����eC���P�e�U��ɘlc�)j�/���C׻T߯՘�\\�㙖����W�{�@ݖN�M{e�I1#",`�W6�m��       n�췴��ɛ^�I@9W]vw2�\]�L3S`у�c�_l��7����B��`+v�7g��M��e읐�H\N!�ׅ:�o7m�2tjn9W<����1�%����avm�U������$t3�[,��ύ&tpNL+u���wx�^��@ߊ��m]�:'m�.�������#l��Q=�n9��3K��5l��$��~d���~`���9��ʠ2��2QI�fh������TP��V$ݝ��ȉG�}�Br��
XԪ�\0;ۺ�!#۲�H��L�pL&a��(g�TI7ܙ&�wUoy�I�-h�Ԧ��NZíH/vXR��&o\2x��~z�=�/ߛo�-�&��қqZ��d����[9�D��:�U�j�~�~��m��[�w.��ݖ��y-D�8R�L�wY���}e�]��@Ȩ�q�"+�@ܖ/Z$���jIn j\����@ݖ/Zc��k�׻JX���R�4蟄D�߾��j`W��]�ꀿ[�d�6���W����Ɇ}�T��`}�y����� �u����ʳ�ӎ�c�q��z�p�"��R�
S(J�'�;�o;�� ��K��?$-�	K�e��nU w2X�i�^���n.�m̉˄���K��88��CRI+I$�I$�Ia�I>D�>	"����"8�LY3�D�3���JF���P`�%C�d��!/&�Pr�WX�nTb�CD`BD!�7�H2]��V
p�b�f�A&	�,�a�![��)#-�ʕ*4L
�X$�1��8q!Ɨ � L�Q3�(� �Th�d��$��9�8
�ӆ& P�#��,�Dm8��r��(p@ઘp��MhM�GhD	�2�: ��@p2�[%����TI��9m�T�ܧ4U��]�`W��;�,��MD�8R�JM��n�c�HW�T�d�)z�..�m��l�J��½���Wm�gs�&����ն,?��d��C���.c�O�w����`u^/�9�r�w�p�J�ܯ�J��-K�G����9�嚘�0+�]W�y�J6���Q��vᘗ}�T��aK�n�9&[�d�T%��ۺ��d܈�L�F�?(�����Dl�&�g��fI��o�*�C�K�e��nU����Y��[n��ߟ= �É&�	6��O^��msнu�/�P.G3%��T���p�7@̖|�Vb`wq��m��0�ClC�\˚$��K�D���'�߽vM�Y��| �A��r�W)N%)j���ᒗ{wFG>�3��E���+ޕ��6�5.c:�������)U�a�r!w�`_�5�I�R|��\� ��亯��2N�{��,l�`�!W���m�       ��=k{ӡ�6�&N�W�sF}�w5�l���4r�=&���w
��ttxw%���mط�h�,��ֺ�1�s���4���MuΒÈ�f�&�6�]��.E�7]d�\�]�MQn��ɶ���Ξ-�O�n�w��ة'FÓ%��ˍq5��Z.����{�w��UU_�˾���N��L=�^&<�V��TbYyRI�p��bs6/jp]�`Wr�;�,����p�fX�U��R�2�۲�����۾	�a$�&\P�ePj^ݖT%՘��p�����*[L��I7A��K�l�:��0+m���f!�	��˚�-0>�eE� ��;�| ���dȸέ&��yՏ3��oE�@���yVԅ!�)����M�&�6��o�}� ��L�r���1.b����L�Xp hrL{��'k���0=�&�$�I�S�唀�f:�-0;�p��zꀿ[�a0�RK���">�j`{uä����f:\^V	̡��Rƥt{0/޺��K����v�m�ہ.9�qae�����s��ޓA9x�+>f�ظ�r[-ߛm�ڡ�w2X]�`ow*(������Kn`�c!&�۲?���'ey^&����}u[�Dr7�2|�ؒls)�k50*��7��@@��A! ��"H,$��E B��� �,Z�ʢI�y2I��jCj��n�#�^ݨ`g�*�;�,>]�Z`���jDơ̹�6�7� �����w0+�s���m�b��w<�jٹe:���]q�sm=��NW���%�Pז��@ܖvO-��p�K��*��Ǡ�b[$�'3@u{�#�ĺ����oz�_܈�2�����N��T��߮�����~N �[�	�a$�&\Pj���P�5�Yi�Ȇăb�OH�)�-`�H2I#D����2\�Z�N�1��HKJ] wojG��e%�c�����$�����o��Ȗ���6ĕu�Y+��u�bT���u�Ͳ��Ѱ����ʒz�nu���x��x���p��R�h�1��G��oP��@y^�V�_bcP�\��i������| DJ[���F�w�a�{6\�)H���n] w��@w�bz��c�s��/}��"/��d&	bm��u{b#��=�RM�ﳙ$��v�$��v�/����_��P        �Qh	6n�.�]p��1�z��j���ay�v�Yqh��](�v�g�#�,����幹��V��e�
�q�ƎY�c��C:��e�b-:8��"퇛�cW�M��i��K�q�ˬr[p�;9���[�	���S�a�*������;��w����UUUp!ʓ�Y�������,�2Ӎ]��n!�;�#fҘ�0*�u@���Ȏs�A�z�|�,&HE4Rb�7��? �;��t��0+��ߦ��-̤��%.� ���&�v�0+|]PȜ����S3-�E�+��Y�Kۚ�=���sK��ڣR��nd��� {b��Pyn&��''m��X��/Ngh��)Ҥ��pu֐Ƹ{�v��~��&4ɖ�H�ʪ �^C�;-m W�B�;�/ȅ)�-�D�~�ual�@����t�Nް�>�޻� L��	�l�X�c�>��U@�8`w�]Pv��x�I�K	mJ��艷�R�ڠ}��>�9�/N�`e���aĒ�q@{o*�;�����R�W�2O�z6��m��q2�KQ�����k`mY�:��f.�Hq�78z�-.�V��onk����]�%�VT8�d/q�=�;�r��R��f[�H#ؤ
�`V{j�;��� �7fV�Å�eKT�\9&y�g2!�B ��U�r���d����@w2Vq�dı�˘�=��YčV���<�S�9�]��`_�?��S8�4ܺ ��:b9��T}�|�����$���ߠ�o��q�K�j�GMWX��<��Y��ff\&��$�6��N�`w�����ZA��t^eBN	m$K��A���#�yT��q@ue��"#�x�'8�\�0‽ͪ �f?���q0=�p�����RɔL6%.�&s��s9>�d���(��" (��;� 0`�u�I�����������n����L{0;����c�;�lMעZ�.n�7��<���ù���Û���r�P�)����c�o�T}����$����Nw��!��M1@{o*�=��@ue�{n���"T�D�\�.�;�����L��0;���/��LL�c��tVZ`w���A� ��/2�'��%�J�=�q���yT��]Ֆ�G~��� ʪ������{o{om��!$�	"H�8�bBa� G/#:J���d$�__	��"�@�0Q� #0� �D��	@!�R�"��H#"�"&P��@B�$HA �% RR!	$Bb�!��!�U`H�����Lb� @�^C� ��Z��3D� Ʉ��%���D��%�Ff"C2�,�Fe00;RXNL���(%45U!��%���C�D$!3�MjQD��%2_|�Ψ$�V�U�!�F��*)-�#�F� #�
�Wz�tH�	B��J!&��!טV,g1c��5y�U����
�E��(��tB) 9&r^BPa�Y�tg.��ΙX%a�w	4I�s�9�5�	O�@��Fd�S"f@W1&���ݶ۸5��z�d�S                                                 �N���]&ƲI�4�hݙע5� �zH��,�^3�en:7�;��I�eD�g�.o�w_ �`��-{�����!�Vأ�ܖu����z�8U�am���<�[Aq��/.�cC����0���OGm�8:�h�sӺŸy�����j:w���y�zV���t�㓵��n�I�)Qs����iL=ro<���_p�6.���n��/kvI{]�\[�c��d���P
�:;P�G9r�f޺y]2�;j|�������/mg����q���gXv�u�Y©����Oh�ͬ\׭���]�qK��c{=<��ڤ���s��́�e���nq���6�`8��%�@��n����^�R��v�sWLn���i��`^���xvz8�km �wc+v�m�=��p��I���LЪ���4\c�}vՔ��7
��[���0&�'F��cv]�n�u�/l�������ӆ2�K��Ae��pS���q�u�xk���j;Y��J���	�iuԄ�:�y�I�*�,6�cp�-4��5�-��y���O��8�F5��˹��8�ۛ��&\�UnssY՘mzW$�uܽ��!�jb�F��M׫��n�s�[�����{D��z���/c$�����5��l�t���B�5��,�$sv޼�U�^�n$����j,�$�w�p@�i�	`W�@>#�Ch0b�E�+��<�~y�{��������@        >O��o~���z�ӶYN�9�i���Է;lj3o���|Yunq�X�@�C��\���^7��6z�zx+st�n�jΆڣ{=c�)�u�+<�.�,.G���4:�;e.5�Ob]&�8�uJ�z�;Xr*�j5ǵڣ��ܕ��3����~��ۻ��z��f��n����Zi�:���y�ѫ�q�*u �L8��Lr��6����n�:��0;�p�#�9ƥ�(�lJ\P�u�Yi��ۆs�U��G�'tnSd�e�M����|��8`W޺�1{w_N�G�59�0�D��-Pһ���Pw1�^��;v[!̊F)q@w/*�;�����&{n}��� �ےV��rv��ݜF;Ow�FBV::u��S	)rD���M���u�^̚����TjYx�L���'-���sүb0bO��&�z%*|9�~�EE�ePj^�u����G���
�a�%�e}��8`w/+�SŒ���<�S�n��a$�&\P�ʠ�cޠ�R��r9���)}9�JZR0ؔ� �ۮ��{o�
�]}�d��Ͽ~� M�:[�y�8B7/f��׋k���]p#\�4s2�v59�I��}�d���V��~�r9����@yE���a�
%�I�$���� 	�}�TI9�y�&�`���$}Ȏ/n��NR��e�@���̒k���i�M���֯���2L��`_�5|&[I����v������ۆЮ{���=x�#���t}806;쨠;��@��@y���4�u�ƾt���˶�������E�и��:�$��"X��}�~�����7]��w �K	%�2�KۛT��t�;�����*��3����ܪ��Iҷ���Q*%D�/��1*D���rZf%D��^�u��D�`I�����NQ��R�u�	0T�9�����Q*%D�=��1*%D�����)���Q�:�2����x���SQ*%D���zz�^,�b�c���J�Q+;�Zj%D��]�u��J�Pj&��k)���TFk�M@�L	0$���+m��m��/S(:[�4�v��^�׷;d6�ge��e�׉!��Y��J�Q*&��k)��b%D���}���TJ�Q7����J�Q*%�Pp(��L	"76j|	I�,�-�I���TM���SP��LD�������Q*%D�=��1*%D����u�	0$�����K%"ْ���A���TM��-3�I�����%�bT~(��LD��{YMD���s�k)���TOw��Ufb�s���&�TJ�Q9�e��J�Q*���)���TM���SQ*%D����Zf$�`I�����a�QM��`I�%*��k)���TM���SQ*%D����Zf%D��{�KLĨ��	��X��Dq����M��m��m�     ��ݖo�����և��m*R��7��sF�Y�7�&vg������c�^{<v�ݣ]��T7�+<�L��kjbу���E'��wk�sk��⼍]c��Sl:u�Y�	l]���t��"��aF.K3�۱r�	�3<�2�[�
�N��w{�w����O[� �<8�k�Ij�O;[�u�N#KۢM�.�¥b�i���[���w�oq��J����SQ*%D����Zf%D��{�KĨ��k��Q*%H�>4�I�-��f�`I���1i�}
����Q9�d��L�*'>{��j%D���;�e5⸤ā&���|[A����`I&D�~d��J�Q*&���)���TM�����J�Q*&�~���Q*%D��+��eӡp�&�`g��P5�TJ��{��j&�I��|�KLĨ��+1��LĨ��w���I)2S����`I�&}�]@���TM��-3�TJ���%�bTJ�Q5�wYMD���l�s�]���\�N�;9:��{[��<�]���=�m��Ķ�]]��Q+����_��bTJ�Q5���J�Q*&�9�e5�TJ��w��j%D�5��}*��$Ų�^&SQ*%D���Zf t��\J���Me5�TJ��w��j%D��|�KLĨ��w��I*˲bb�1�2��Q*%D߻�e5�TJ��w��j%G❢�\N�����Q*%D�=��1*%D���}:Ix�VUK�Uw��J�Q*&�w��j%D��|�KLĨ��k}�i���bb%�{*�`I�&����M9
SS):MD���o��i���T>*��=��Q*%D����k)���TM����Y�&�`otכm��s"Hh��b�������L���6Ů#�h�{��x�J�&"b9얙�Q*%D�{�e5�TJ��{��|&�b%D�������Q*%D�{د7F(ŕ%]�MD���o�}���TJ�Q7�{YMD���o��i���TM�-3�T�&�ϭI)2S����`I�&��k)���TM�KL��赁�Z�$ �l�A�!�G"r's̖��Q*%D���e5�TJ0;z�Hh�l�N\�P,��L	03_��`�J�Q7���J�Q*&���)���|I�����j%D���W�e���@�-f�`I���D���k��Q*%D߻�e5�TJ��_��bTJ�Q4�������F]*μt���UH�V���������[�#7l�vC�bce5�TJ��w��j%D��~ﵔ�J�Q+��}-5�TJ���%�bTJ�Q7���Kĺ��]�c/)���TM���SP���LD�������Q*%D�=��1*%D�����)���TN/�����W�]�UV/)���TM��!i���Q*&�ܖ��Q*%D׹�e5�TJ��w��j%D������b�Jĳ�\�j%D������i���TM���S���J�Q9���SQ*%D��)gh����w:��bTJ�Q+���r軅Uٔ�J�Q*&��k)���k��}���TJ�Q9���J�Q*&�ܖ��Q*y�y��|���V�Yx�&\F���s��{iԜ//g�f��w�7���{�������TJ�Q7����J�Q*&�ܖ��Q*%D׹�e5�TJ����%���2��n�Y�&�`f�bTJ�Q7���J�Q*&���)���T���SQ-��^�TO��_h�\��h�"$��L�8�TJ����Q*%D��{YMD���o��i���TN��%Ye��^&1fSQ*%D���}���TJ�Q7�{YMA���o��i���|@	�����J�Q*'~_��%�]YU.�U�SQ*%D�Rs�=���TJ�P��9�����Q*%D�d��J�Q*&�s��j%D����d C $ �i'�)xKm���ۦ�       Z˭��[]:�t�N,�"[,EM�m�qz�q5���ۍu����\���^��ۋ�e�3��\{puٝ�ݺ7��n�/\ �^9n7V��N���=Kn��b�[��w�:�<'#<물�WW7�3�������������]�{z_~��7�Nz�ש:�[��u�Foh����3����e�%4�-9�I���L	0$��ύ�bTJ�Q7���1*%D���;��j"TJ��{��j%D���&9��z���,�c2��Q*%D�=�LĨ��k��Q*D߽�e5�TJ��_��bTJ�M��z�ˢ�x��$D߻�L�$S]�s�$D����0I��v$�H��+Պ�*�w*ꮱsMA$~���$D�=�L�${�ؒ	"g��`�	����X�^+���D�I[��3�M�bH$��s���H&���"H$�t�������%�0�k#���A�����F��A�g&ni��&\��(6�K2и7|�{����s�'�n%D�=�L�$���������LV/"H$��w֙�x* y ��U(o��J��Oo��D�I��3�M�X��so# �p&�$��9�l �&��Zf) ��l�$DϷ�
""���iL��e�B0.%D��֙�H���,I�3㝴�@������$�H�9�_(��*��^SPI�=rX�	"g��b�	�w�Ȓ	"k~��`�	���rU�%��3�QԵ�n�|���A%��b����K�b��.�U�2$�H��}i���k��r$�H�߽�L�$S{햜�PI[��N�c������wJH'=~�D�I[��3�M�X�	$
��F�DZ�	�
a��r�$D���L�${�$�������y$�I$�I%}` �<a��B>��8TC'����`o)����Q�uP�P2b��]�,�T�F1��b��GeR��md�����S6`���sxζe,�Z�6���%��B ���@�\�]����M�J.;S)T�r"I����+l���� ��j�5���Y!$�XKkIp�A ��g�K��r��sA�p���b���5�7kuw�V/$*�E�[��D�XBd��T��&��r�Ƀ(Vd0� �P�f�,�����7w��"��QoYI���V	�bK���\1xҁ�g0��B"�b&�@mT�*e�S���DuCh�(al��28B@�R`�/@]��U�)�����������KL�$~���$RD�;��,�x��U�)�$�s��ĐI=�m3�M{��D��2`f��D@& o���2�`��)1A$D����0MU	]�s�$D���L�$[�$�H9��c�wwwww݋��]vE�tŲs��m�:�0Q!�<��붝�%B�U^SPI߻��I�5�z�$A5��a�H��5�-3�@�O�|i�Zs2ӡ � ��y��$�o}�đI>�m3�M{��H	� �o�S�$�RI�""{��E$L����A5��D�I[��3�I���aWuEܹ�]�A$M{���A5��9A$Mo޴�@��&��.�B��P���  ݳ�}2�b\˔�A�$�o罜� �&��Zf) ��l�$DϹ�L�$�N�{�wwv�:�@�j]�vnnl�I�8
p�e�{\�ʬ�Z�Z%0�M9n�"L@&���Q	o}�ĐI?9����A7���D�I����K+/��x�j	 �笵���Е^�3�N|糑$D��z�0I��I*�\&&/�řA$M{���A5�w9A$Mo�-3�Mo�X�	"o���KĪ���*�)�$�o��r$�H�߽i�$�k}�ĐI>�m3�O	�<i�Zs3)ЀH�L�y�� ���lI�3�v�0I׹��I`("6 ��Fe�M��m��m�  �`�   /�� �n��G[�c�͕$��k:d�;]v	��9:�4۸����k��dv6-����1As㊻Q�lgu髜j3��c=�����clݳ��:9�k��Ƕ�T�t��5Ɣ��.NC�&���a�qY䨫m�.�E9-��V=�ww�{�^�w��ힽ� �]sN��d�L#)���̀/=�e��h6�[2�{��H��ŉ �&{��f) ����"H����֙�H$�js�����\�.̉ �&��KL�$]�s�$D���L�${�����I��|��cR�]b���T%|���I�5�z�0I��e�"�}��f	 ��/ĺ�S\�/WyA$Mo޴�A7��bH$��s���H���w�Ȓ	"/�xxKfRaHL�UȀH���@0I=�m3�M{��D�I[��=N��;�濻� tu�5�v^ѧ�Q4�j��K�a� �QJS_�U@�M�� � ��}c�$�k��+9A$Mo޴�A9�YbH$��s�I*�e�Wr��H&��d���D2�"���l4�	"k;��`��$߬�$D�g;i���x��t�/w+uU�Ȓ	"k~�`�	���A$L����A5�w9A$Ooǧ�]��Y1�^SPI�=e� ���󶙂H&���"H$���֙�H$�js����]K���"H���w֙�H&���"H$���֙�H&��,I`| g��m��m	��2̂�=�x��������)�BB�c��9��+)a��~�{��>|�D�I[��3�P��l�$	�^�p(����)JR�)4弉 �&��Zf	 ��l�$DϹ��$^�s�$D�;��YUvU�W�����z�A$L������x�(B�j��!� +f�������5�=�|��A��h���)1B"0/���I�9��I�5�OZf	 ��K,I�7�t�%Y,���U\�j	 ��}�� ��9�妠�)�z�� ���D@$@�����m�	̙���u�X�#���[���1��
-״�j�@7ܒ	"k~��`�	���ĐI>�{��3pI��|�D�I|��|�QvJ�p��^SPI�=e� �&{��f) ��;�� �&��Zf	 �]����^1rbV.܉ �&��Zf	 ��;����$Mo޴�A7�YbH r/��)�42Z�5��(�"9�UP�	"k~��`����D6bH@I�$��Y�$H� �� ���3�L�$�9�˪�&,��^.��$�H�߽i�$�o},�$DϹ�L�$^�s�!�>'y�?��� �n���;����v}����e���v9�[4f[����� ����H�&{��f	 ����!�A$M��8D`I���x����I�	D����0I�{��I�5�{�MA$���'�TD���ĕd��*�U^S��$�>g9NĨ$��ͦ`�	���A$L����A<'����l�nfS� � ���D@0Mo�X�	"g��`�	�s�Ȓ	"{~��⋲�Œ���j	 �笱$D�y�L�$^�s�$D���L�$��N�JT � @$d�;���w�O$�t��I�        ���+Vm�[z� ur"玝۹by`���a�W\+i��'��K٢�� [z;i�/W�d.W�}����bCJ:�<
E��{q�3s���%wdf�	�dI��Pf�'�t�/n�6Yn��fǎ�sY�-،۞N�N,�1���{�������{���q�ʪ���m�)rC�\��y����j����`��ܦ��Ӵ�����w�D�;��0I�{��I�5����H���1 � �{>��)�)�j��LĨ&��g"H$��{���MЇ9�  ���Q	4f��I$�wWx���D�I[��3�M�X�	��;i�$�{}�r$�H��|x�J�\���F1��A9��bH$��󶙂H&��9A$Mo޴�H��ρiJ`�M�� � ��>i�$�w}霉 ���i�$�k|�ĐI�Q��{�wwwww$��%���y�Ӻ۞��tyY���k���.˚�=vŶ���pI��|�D�I[��3�Mo�ّ$D׻�L�$Ew�+�������U�Ȓ	"k~��a�K> |�M
 BFa@�U: ����Ֆ$�H��}i�&�����r'�%P�'�|�>^
.ʣJ�/)�$�s�,�$D�y�L�$_9��HA����
�$���%��%�b��I^�3�Mw�dI�5�OZf	 j�l�$D�^�ڬ`ŗ1u��SPI߻��IQ*%o޴�K�PMo�X�	"k��`�	����� z����s���ոn4�沷�$��k���Z����M6������
"�w|�ĐI>�m3�N{��D�@&oxx4RM2����HfDv�dȒ	"k�}i�$�w}�r$�	�y�8`}����ZR�.SS)�A$M���L�$��s�$x
q*)K����-3�Ow�X�	"o���J�]�Uw*�)�$�w��r$�H�߽i�$�w��ĐI>�\
""���)4��I�iЀH�L߽i�$���9ܖ$�H���Zf$@�7��D`z �{���m�� �`Ӻ*"�غ�r��/M����!�-��N��U�]�7�Nw�X�<�Q7��`�	�|�r$�H�߽i�$�Ms��.��.K���2$�H��}i�$�w}�r$�H�߽i�$�o|�ĐI m�攠�,�)�P,���z�@�I[��3�Mo�X�>�l���,)IK��L} �}�/5 ������������!�%b�S��J��B��A��
PZL�q�}����-�%	L�T/5 �5���}�{�> 	o�Ļ5M]z$���V���z�a���sp��\ʐ�-)L�����m��C3P����a�J��ˡ��~��y�0r�0�X�;��M&�SfZqW�����:�\u���HlJA�����8&�y�X�qW�qX'4�Ô�8�����=��Ӿ{�X� �g�c?I$��j��P@��x����S���R  �x��l�X��J� Iڤ�0gE�1�`V�E	H1U~ٹ-C9�a�P��&��*��0!Q�Pd�A�G�
���R�(�*���%E����R� (�("p ��X��!�B  䊩B�P1T�T� �ȃPZ�ĂH`0�F�"T�E�Ws1DP@�DdP�J �� ��s�܆k'��MJ'���?����� @~A!>����s�}T?�'���*	��~g���#�EG��2��*��%��XP+�5�@�������`��`�������I             �                p#� �s���G�~���tڠ��.���}�׎S���S�L~����o� ����}G���d�r������DA�����@DA�P(C����J~_�~�?��
��x���U����_���~�O����!"A�!	#$���~��|��m�������|��bg����$�������b&�K��9@C��ꟐI�����!������'`��U%1B��L 1�EREP	D# D �DE	 	$ FDB0P�dBD�VE$@	BDT�AY �%
��@�AV@@U�A�EdRAF!	!B@	d�XAA@�	 $EA$UdBPIIdE�Y�@dF`�(�! �,���$�b��#RFHH@�dda$D$dH0 ~�(����I	D��$@��D��PY����Bcd?�"������4�UC���d?3�������@�o鉷���ϲ������ �Ug����������"O��L-��������Oؖ@������O��F�>��������O�?��l���X��"��H�0$�k�~c��?A��!����?Q�"�DA�2'� " ������ɬ��0\(�	�!���E����B""�O�$�b2���>QhL��(C�ɐ5G���@B�H	A ?Ƞ6	�&�����%@�I�8�@����D(����	�����?�����؋�>����������|?��@��������?������̩����w�O� " ��)�)������?@�����T�O��~K����y��t�xz�Bd��+`?RH1�I��D�K�H���W��z�,��Ҝ�؀��g�p��ϱ��&>�E�⯎F���A 1���bd�?bd��(��>��b� DA�H?�����~ p�����Y�{@�"���e?����T:3�l�?<������Ї������]��B@�& 