BZh91AY&SY\Y2�y_�px����0����a�  4 *( $ 
*@ @J�+�hT$� 	P   (�D��  O��  � 
�@ )J�*�
 D�IP%TQDQ"������@�B*U*��JU *(��   �`� 

    �e �{�9;�7��ע�t�3�w� Q���|-��VY^��������{�s�F;���V�(^f�i�}󇯠{�Xt)�åS�ç��htӝ� � =t���Ss4���6N�+UT%G��   � ��
��/�y=�W�bһn-J�Ϡ�U��UNM}j���}n3T��� ��U�x�W�}PR���j��6UV M�J��޳�/�}�����ʗ�� �}�Y��[�Usj�=�y5^�w��U���|      8� =�O{zW�W�+�T�ۋR� =�U�U,Z����*�oZ{� }ުW6��������{X�Ϸ+�w|���>��)Y=�W6UVm+�si.��Py�L�;U���NMW'.T�y�O|@( � ���{�U���ҽ�����*���,@;�,��y^l��s5=��Jg��zR�n���>z P�^l���ʗ>� �S-���U�)�J� �Rť,��\�^ۛ*^�E
��  
  �� ��ҥ��g�ﻩ�eɥ�s5K��Gz�b�u9e�ӾΫֽ��U�(=�S'sS�_z�	 �<����iV �z;Ԧm���9׌�W6咮����f�}�W�<����w�ꗀ          �O�
o)J��      S��T#F�     hD��R��y�1��0�F�=��(4T��  �  D�	&ʔ���@i��i��L!H@�$�j&�i������`�F��i�
#�����������?Ň���:��u��*�*�����*�ES��**��QU�%P���*��xF **�����@�������mP� jG��j_���@� 	�eD��|��� ���!��?B�}")��(B
}B#��І}�H)��?J�!�}�҈�?B�d��?J#��:�W�C�@�U���@�T�UC�<�E�D~��`U��@�~���@D�P���T�E>��C�AO`C��>��O��C��@�} ����(�BJy@� y �$<��T>�r}+�C����~�;�(��F���Uj��7��{�sݙ�W�d*�� �S���)䢾J#���
}({*Ҡ}(BB�}
?J���B��
}(�҇�#�">�J@��
�H�y" B*�"w ���y
���H@���"���.����}#��r'�/���B}��B���J�+����{��&�#��~�����O�O�~�>��!䇐��䧒'�|J?^�}?I��J���H} }'Ӓҟ_@�'W��/���)������z��Gp*�"?BJ�􈏲!�"�_��������Q(/~����s����P�\"���wz�ƽ~��L��鼙&���#�]�叜}�-��;���_#��\c�:����y���y�i�=�o.sz�&���6��e�u���Ŏrsw�SF�m_=���D���<1q��Rdه�4�-Z4ؕ��,l`�,�>�q��n�V��}!��%	@�	BP�%	�J��)J����^��/�8�ؖ#��5N�ص�2#�a��rh�1.�h�@�1W?
��'sn�$�{���K���uW{�+�3�r��C1ս���+T�]+�Gw�3klz��9^1)a��:9	X��Ls]k"š(H�*�#�8�9t1�}CNa�OR�������u#-�-�w�ܭ�j�ޭ�yvx�a
ht���s8V:�ui��v��5�A��ݕąD,���m���ge��S��hʵ\.�<�r� C��::�WyB7˽y>.Ogc{�5κ�g�9�j��=�А���n�T��o�;lD��piN�5GR2,}������U	et��>6?�wofb�|��Q�8��1�FKWB%�����y�:��$�t\��;�kg��0�aI��C�d%M'Q�m����{]p_w�9�ܬ=X����t�=g�G�T"�7�7V��V�(z�ǧ����L��uWMˡbE��H�����Y��[��H�>�N�ڥ���n�Sx_Kņ���S:6G��|����f^��]�d*�vJ���:c���f�ШtԾ.'1o76�,�%��noke���#�3���k;�:��0�!Щ���!Ž�~�p�7�j�2�t�q^�����&a�bW�����KL"�����go�n�g/�P�w�g:v�u����a�{��.��������:(�|��k��|��N�<��%	�&4o���GN����⒞`�Ƿ'v�0�D�ܙ{Τ��9�=9�pE˱fbFpV�g���j���X���t��UX��%�5f߱�yT7�������t��v֞���ey׫o�𴽮���[|nn��= d��h����צ���횑�T���[�#�<m�f[�L<#N�[�w�NZ�g1�kk);�8��r*J�8p��)j(���2�MP��h�EfN6�NTA��xsCq�3�s�:+8�K2���n����abV��2�n�q�.�.g)x�%f
���5dF^�U�ʊ�Sʫ)��0�B�f`�[˾�2��J8�u�k!(JN&BRbdh �EmEp:�mY��J^i��Y�L!��h�_(d�P�`!�\1%t��6�C��,�˿#�qSU�D�NX��!��K�7�������s��z�!ahd��xGQ��w	���Jq}�äޠ�x=����t�{��Y�{�E��4~����`ŉ�z��J�aT�f��
(�R�R<�8sr�c%��H!Z�{�)α#�K-L�1�u%���U�7����_!�� O/����@HC�Yx:��z[ú�Ll]���1c�ˠn�DL��X��ڤ�I8')R:{�k ��9|b�H�F�EM��4fd=5�f=�)5�o2f��B��K�Nr�/;�&>r�<�7�Ԋ(Hg����Mx��fV8��K�P](��N�]�sݵ�x�L,��!.\ ����͜�
Bdj���F*���r��M�'��x��8+Tp.#+!�� ����|C�t��Ӧ��9j���k7��SN��|�y�7P�떳��3�qf�P���3����1Đ��ц�|�({h�4���^��R���0�S�9`w��#l�[� �tjăVh�I��惍w��;�4m�̐�C���˥��x+�j�]]F5���K�i�g!w��n����@fن�F��67�m��x�9�2�(�١�yy�sC]f!����8�	�`���bUM���U��V�\������eX�����[.!���3�\�:Y��廤���T*j���KA2z�����	�D��7��jwX�]���6�О��ڇ{�C%��*�8�{$Ie]-��V'J�qesr��n!G���*�s'8�P�H5}}|�z�Y���8�{�9=XK��BrM�XK���0���J]�iq�2��'Xp<�	�B�i���ڮ�ye%�D�'da��$"�̾�+�Z�Vww��#�<�wN[�bu�8*m]��qS�k�4E=�'kUr�5���5P�Z�f���SW�&��h��xIF��s�_�`��J�ݹ1k�Ӏ�1n�
EV���k�pC@� ^V�j�s���^��8pȲh$K�2R/gb�!�E;�[}49\�R6]	��r��(U���.��Sh�а�X�@R$6ʨ	`��ǧ�\ִ:=�,�D+�4�O�
���xqċN��j������'I0*������ 1
�P�����g3�fX�sP������2�ո��Z����K����k6�M��S���B$��ӹÓUj���e@h�0,�)�1��c��$gFXkݧeW=�4�՛�#�U3�$Blv<4ÇGJ��⼵��\�����J?[����|'Bi���V(��T���Nw��5.6J�".2�HP�Y�q6{���8���Џ21�J�LԪt���J��{<��g|����zk��6p��;�M�	����*L�]5v>3�o}̒�U�8�&��g�#f*F&3��$--֎/._�-qU	P�BP�'����s9ٙ��U(w�/�r�\��2�Z�^��j�6Z�i7�r,2�k ��8��u���}N�!V)�ּ���WһFR�#��jG�{�_9�}oAy�r�<�0�)^5�喇/�乳E�xmo���2{���B�s��2p��C�D=�4K��������6j�k��&p-��LES����_l� �X] ���a���LL��		�� {K��&���~�����'J`�NYj��u)�d�~�[z�x:CR%	BP�&Bu�	�'!(J��	�J*�;�w���YyE�"��H�E�D@��B�nea���膩"��-�{}%�ҍ����*.�BD�FI�n��9)�MBP���D�:��M��y�!+���*G-VU5L��{���+V�!�h��m�wt�#��{��Zfb�V��L��-�l#�*��Y�+c�M>fq�_:ox�2-�m����f�%�&\��2��h�jR�d��w;f�;�?�c8:D��Y��[2����XX��be�R�w��9��|�z�R�}�u��GM��L^h^�Z%�|���r73�ټ�X�EN��0BjR�������y�/O-��S��7<��g��z��}� �ZW};�1s);8t�&r���X�@�3w�^�Pb j����mj�5��<�9�)vY8��i��i����$BVE&N���4P�P5F�:D��P�d9!�G24�Zn�ss����É�<�}�,X�|�ӚpX�]+�t���O(��N�"2�S�yn^�8��!��a���*�d��ef�榪�R���NIfËW{XoV�j�)WD���V�77zp����ӆ�X��6�{�]�rx{��sǃP2�a�����'vf�7��V�
"������!6����w>V������wள���ɡ�=���f�wx��.�x�{xoN#��N^�u��)xf�	E,̭5r�zY��T]�o7g^ܩ�t��@�Nb�9͍9�xԄv����[Tӆ�[0���d�T���S[@��Ze�p��8x�Nj�D��34���u�����iį�)LՈ��b�d���f��{={�B�P�*�:��7M�B+�6�GR�3n��}�B)�M�9׻w��|j�w�����P�b�t�:ox�Zv��P�˚r��*�o��X!�9���Z$37���/�U"��Q/4�*Ψ��C�����qC��X�W��W���C�߷�8����Hխ�ޮ����c��(��K�br�U�Z�����n�˫GL�E�9�w�����3���V��Ě��rMZ��SM�rڿnox�H��A�;�ˤ�Κ3�L�-z�ףHI,m5�	|��KS��<vEbj��A\Y�{H��T:GQDD,�q�8�l�zfS�C�E2���U{�!<��!5	�NBn�M�EE	d�j{�}���6\��2��vBB�v�|�.JA
�u+���)&�bR����3�f�e��P�3��a�ގ�B�:6N&�Ҏ�,�$�rp4��!)�������!5 ABj\r�3 �ްJ�M��`b�C�	��(J	I.6f�׻��$"�i�\g+k�P�����,�]2��u%��@b7���U�$�ช����C����6��J���c.���ںFC)Ze�Q9�����/�hbjc��T�9��C��ޚ&�1��tډ�%uf��%�饝6q�Ƹ���l�TT����֘8i�杇�j��8w=��&#EEJZ�5FNj����Dy�n����H�L��3�2nU����Q�ޮ����N�r��`:Bj����2���8����Z��#��`�'�pۨ3N^�{�՗1�d1u)p�c�ģ��-E5	�Kq�D�y��N��3�9��t��+]�q^qn�r�^6�
ǰ��*�%$��#o^z�v� �[Wǽ�o[��>w��x��TԊ�fe�E�|���B�:����^'z.uNf�-wS֕>��Z�+l�L�)��$W�3�ڊ��(J��(J��().�5��!�BbI4�Hr.V���8�\D-
��t�eR��z3A�}1�(�"�J=0���d8	Bw��!45F0����C/]��4����`xj;L��B�<:۹���qiԱ9l��3���u���#�<e��Vf�zZdC �]VbQqP?FP�^a�����A���������mRZ�]a���PӡRj�2;����r�'^�e��:$Up��&p=|��ә��J��f��������U2@�9
�"�f%z�4�gv�i�P4[���9����S���pUS�螞��6n��]���"�"�j���(m�J�4�~��N�Y�k���^RpVܝ3��s��[LJ�y���%�i�hu.������D27��}���5;l���q�;��-�
�.��������3y�y!�D9.�%�8�/�i�i��WV�Z�._V,�F1�W����N�i�������B��4N���|�*�
��HUq�kiƖr2�]E�[Q�k ]Z�
�:@"R&]�c���uP��o�%W��2�K3�d�.���Qsۆ����^��J��H�QBTr����t��:��!��+s�RY�fF�	[N=n�4���;����䚈ֶ�g,�9�u���PГ��'{M����@R*L��g_1�X'��xuk	I6����x����6�M�)��l-zNn�[t�ë�3ɼ��o_k��5��C�Ϻ���=�<�9}���&�Ӫ?����>?W��[^K���]�     8�              6�@     9Ì���    :� �m�  9J	7[@   ��8�    R�       �ǅ�        p         ��R���r��J  d �����  �m�m�          )@  �               t ��� H�8�谑����j9a���Cz�/YU6��E9�pu��j�/lSWY�\j��h�� �I���w��yK4�rf檨� %ej���tFN�x�V�@*g۶j�ʾ֗��N�Em<�sƺ��i��:���-�Ke�v랎	�s��N�Oi$���<(M��_O-�R�Y�<��-Z�U�����UT��׮r;[��˜��t��N˴f�G��9GmUV������Y�E�+�v �MskOi�g�>.���H�V9���u����Hv�v���#mY�	YżvX*�#V�b3A���.�*�@�9��Vzcs\(!s����u`�=�MU�!�l��
K����}�C��,��W�V୪��3�!Uaى�9v9���UJo 9���nݷbj�u�]F�m�@�`�8ZmodۖΖ\��%�������Я*�g�C;��g���[X�)���P�g��h��`'lc�a���Gejڻ3�=�)�*��ӽ���\�k���}��4�T��X��&��H3��%���T�۫%Ol���g@�&^�vy�� ���s��<=���<#;<ڷ��(�,J�5�m���/c6e'l���<��A[���ΎL����؂#�eD������v��G����M7�#��';v���hRw2�V8��8*��#q�v�,M�צ��g��H�6V� j�-Af8_UUR��Ҵ����J�j��6��NP�� 6X��	�@u�q� ���v��T�*�R��m�t֝�l;���Q+3��M�4Άp+V�l ��v�kf�����m����� 4⑹{tU�UT�@�R�#�d��4���
��)v[n����gt�@T 9�m���m'kp�6��R�:@4�V�ڮ�.�P n�m�[m� ���۽ BF�z�G0����^��It�k�$[K�l��nC .�;НVK-_U|�;�����u����y��ɥ��U^�:�5���JHm�u�ě���L������!����"���μmCT�T���+*�������2H�^�dZtN5��  v���U]��ݺ�r��ύ���U �������b����g����6^:K� �&R��x��u�o6�
���7�kɸ��3��m�[�r�VG���~ɷg�Ϡ{6q�<�ףTj�0�rv��l�Y�y���Z����`%P � �S�t ������8N��,�[�R�e�-]�ɖ�a�7m�U�n�K���NP�^\��[V;qlT����c���c[ˍ�x� �Ԡl�j���h�J�mPI�V�ǱYG�zyU��^�ʎv���:�iX%v�[-;m۶ݳ�s�N��-+{-��=���lE�b޼m���@t������ r@r��I۞v��y:U��A��m���i �t�s�n��S�� :0�v�\�$l[M�e���[%� H 4kwV�O.�c`V�ڪ������\Evt<�B�6��-�+�n�)V����~�����H������   m��nl�lҤmvv�e�  ��C�[�-saz��ɲ�@����,Zh�V�ཛྷV�@n�$��RW��+b�� QT��9�m]��\�va�M�*D�l�H���e���u\�� ��V������Sa�n���0y��U�x�SMڶ�C��  ��   @��liW  �$�Cm���Z	�̀pp����H$   �v�Z'G�Mb&�*��L�lp է`HB�m�  �n�M�*Kh$�C���!�*�V؆9��ۮ�mt��  Ԥ����Z��S�ԙ�����N����Q˪d&�ڡ#�f� .�����ʷ�6۔�`m�^]�a� �� 
P �$]6��_�}����q²�'KӬ��q�� �[_p�� I oJ�݇  ^��i���۶�u��礹j���B��1R��%�j��Ry�^Su�W<�5\n���F�K�$	;v�Qz@�N����z�K+ju� q��6 �8E�H��x��組Ui�
��(�����|H[m�KJH��������m��5��3m�m� � �tԲ�ﾸ>�b���Ö�&_[1&�UCm���SI&��	 r���Wl��if��IrY�!�m�@ �ٷn �i�]Ɗ����_lҒ��T�W=]�������T��������+�@mPһ�6N�����5\ľg�X��:���]�=�S`���j�{YM�n͌P2��]UU\�U�7��0P��j����;p"i�gFIoP�C�ё�����<D��U!�eS�*�A������VZ�� �<�ty��v뤐ݦإ����۶�ۂs09�΀*���Bv��nO�}��|� 6D��U�j*�j2>���T՗b�laɃQ؅��[mM��-��i�K���p [Hu�6[$mxݷ�%�1��v�HJ親�bs�7�k6�R��Y&*���)�XZ���,�طC�b���M��:�o����5mkfV������ɗ�Vn4�V��E���,�$����t[:f$ �  p� El�ɛjm˛�M;R4PI�4Y9E�W`m�    j�9n� [v��:�m� m�UUU|j2�ۋ��w#� �DʵYv4��ܸ�ז1ugf�F� �Ұۮ]�aNdͺŤ���S�����e�f��c��-Uu-V�Oyn�� �v@Ve�s�����\�[+h��ܗK�냜  l5�:��mUW�{k|*�D]z�sfAp���
�BzM��b�����mGT:��:G[R�K����VAi���[�Zt�r�SG�j��xZ�
vY�A>y�ڂ�a崧n	��CѺy[8p�B��ە�C։����*�K�\�n8Ij
��ٻWT�n�O:�+\�ݖ�^}U��PT���ů����J�h�&�rm4�e�;N�;�V�pҦs�:� P� I���0� �֕٪�����4��wFﾓ`v�<�I�V�f�հA��hr���ek(�������e�3J ��-R�VQ��2�Ͳ�l��Jolb��e����ڵb�,!���S�-�^��nd��c��8�k��l�M,cm�:Gcs��cFH��6����2� v���r�uy����9����:�]�j�^�_>}7�d�il�I�7\L���m20[d�7&͵UV�T����À �s��ͽ&�L��LKvٶ��ص]p 84T�6�`�gSv�7n���ņ۶�����W�� C���M��P
�Bj��t)"	���*��aUN�u@T	תۖ�h���9�5�HL�Ul��Um\��ܓZ�(m��#gP#����D�i$�]�Ҽ۴��U��U��̀�-�m�l	 r��-���P�����rūY��,�Cn�� ����mf��Y( ���Jxx�U��WcU�	RI�Y7�z��E(N��U�%[T��J�MZ�h� ڽ�D��a��P6�;i):��m۶����R�q�V����綝�#q�Uܫy�^@�X[� m�έ:kd�"��z�eZ�]�n�m��[8�pj�ݮض��ٴhIiy�qkUV0 I��F�>,��|��F΀�UmuFFIjړh���i�U���c��V�Hr���[F���{-��Zl7p����,�56ԫR�Y!J5`�X�W�����O�F�ꥍ����6�w�7m=��us���(�n\� w�W��^I�,4p۰�����f:ő;`�m�m����mvTuF2EV�l�*�v�Q�Ҡ�Z��;i;7%UG��9��nQ�ѹ9�u�C���K���T��BP<�
ڪw0��N�Ê��y�݃v*�������0;c�d��e�S( �`����􄜙�#D�9+��n/���� ��9u�W�n -y�kR�t�l�fͲ�힦9�nm4pz�@j*��fa�,�ͧ���O��� Ե6y�[Sm�9$�E彤� �K���$ i�id�I֘ ���6�m�۪��F��8   �ջ5����0�m�i�m$� �� YMh e�� 5���٘6i��am  �kX�-�y��	-��  8v�UvF+��1�+9^���i�ڹKiv�[vu�Tv+B�</�i�M��e��f�lC!ˬ��ք-��8�z�L���j��[���㥟��﾿k�U��ˇ^7mZ�����Z��^��7A�j_-pC3T݀��     hp m�� m    ?�      �Y@8  6ٵk��Ot]l���B�������TUU��뽀(z$�������������j���������������j*(V�)ȧ&jH�'"��� ������2rr"h
fC�����O��������[���; 샲8qÎs&A�8qÎp�8��9� �8��p8�vA�d�vA�?���/~}L�h�0�O�
�ւ��z ;��A%u�)ѥS݄J��!�"z �^ ����Aĭti_x�u��C���x{D1]�*���� ��H��8���A|U:~���đd�ߏA�"v�����t ���EOL�D��@�v�@� �VOPШv*���G�v�@������@|OP��'�#��xqU����
���g�x���S�:H�� �@z�0��'� �I�҈@�ګ�
' M�B@����_PeP�����j'������ҁ�A�YN��P����@M �hQv�Ꞩ���2EC�� ��Y���$ ��i!�($��)���D`�(��2�����A�D� �Q�T➁ي'��UE;Dz��D$T��0{A=�A�U� z�!"�̙L�i�#0��Aؼ|E|T<N��6>�I睻EШ�ȓ*��a! B�D;Ҝ{@aU<@4�f������ zv��(��?�*(������_?�?�������_���m����c?����:
�505=����I%1S �D�JDTTʅ
�I4�0���BA�)H�D��P���3:��;��F��� qݾk�  A6��`]7}'ŷ����Y� �J[@  �l(0 9�  #�  m�/D�awT�;m�j	�Fup>�n囁�Q[��]d�K3i4We!�5�ml�w�I��힭�v�Xgq��\�v8�Fr�8�:�B��[��#���R3ۻ/l�fR0�s-�)�T=3�����QB�9��-��w���:��۩|�{N�Z���lf[���*�cN�6<玚(z���K��T�9/K`c�8�1��p4k�ݘ����<�t�6�m�TZckkt���st����sv��g���v`�B�;ln���p����t��i�/,��"ut״�k����^.N�6:R�<�m�[�ve�t�ۥ�T�-�p;�u�G���ҹy�8�h�gX�I�8�ќ���;��;q"�T�J�7C���U�(k��2q�]X��
����c����9A�{!��9�i�/Qٴ;8��e!I6�(4�F]���ksu���ѱٺ�;�5��Z��=��*d�y��k����u�\�:uڼY;	����]����g&7�p���z{=Z����&�'���)�����s8Z��� É!��HLp]�����,��CP���(5-�l�mVv�%����
Rf�N}��ݶA��vPu�=�ltF�x��U�=��[E�Ei�� ��S�7c�Z�3;��w%q����B�`ޗv����u���8�`m�v�v�cn^��Xଧl��Ƨ�v��tT�
�2�]ڮm]�6	����âa�s�K�uN���ܹՖ�+�YT<�Ơ�#Tҕ*�,�<u�v��Y�+X�����<�5s�=	Sn�A�흣T�ƍ���5�!�g.�	����;r�ܮ�/E=�A�.�rc�k�j!ǧix��fuq��2���ge���u���3J�=�*��ysۛi����s=���u�g!w�&sr�c���u-� m����o����rN׀ނ8�h �����������a���C� N�@��כ�G۴�t��p�i�Yna�n�
�e���)�n���=�y�m��.Ϥ�v�9�v��#J49�G�ܧ(�r]v�{�Җ���K@g�\ꗍ�`��p��O`��� ��n�cEN��:�%=������:%� =ڐ�s��:9�H{K�w4�nwO�0ܵ[V�����}Fz�-ڌ����lv�îu���,Aj�$]�6��
����L�G���=�ܻs�s�y]�۝����q۱�`^��ˇ<9lQm��-{���\�e�������<�`{X�5l9%:��J�{�x�2uRs�|��7�d`�{5(�T��ʔG%����Xǘ��+.��{��2��r�GR�T)QX��+�̺�:��v�~�`{���q&�r���8�;�˫���`}��V|�����mV���RTn�"Bg��t�)�ۜU���u��Ʃ�9�<\�鸕T�QӒW@��m;�?b�;��V}�u`u{Գ�Q!C�ht)s\��s�	v���6��Y:��8�0S��N���Ĝ ��&�� gH��� Ca#!@�Y�8h`sZ	��B�,h!���� �&`�0,'"b0���Ci'2"lFC4���{�^��}�˫���`�0$��NST�&�p�uNԲ0qȎL�):�:�j���1�%"m#�X�eՁ��c�>��+�~�`}�I�UIR��b���{����X����f]YA���Wյ�7i��	GH^��P�@�=msv,�lN�6��.:}����'A)ȩND)@�<�`{��V}�u`ug����*R��T �S������� ��g0��XҎ��șa\7m')F�+=�u`u{��UA� *7@WIF&�}1%��y�K��Q��p��d�������c�;��V�̺�z��Q!B�ht����g����+�f]X��+J =��$�Wv�w �MҖ7l�o$�k��O�۷S�{U�l����}�ζ��E%4�UU$��c�V�̺�;��V�=��;��M��hp����|�F8���I��i�����>TLɍ�T�)�5%X��+��f�s����U��ݺ�༚�	RB��IKx���}1%���ėy�a�v���A@�BA	#*I�f"�t�&m 8��s{�r�|���*j �S�)��?b�=�eՁ�?b�>Y�v{Ѫ�
���D�ˌ�նL6�s���ӽ�EZ�3�Vh�w:�8}I��NJV�̺�;��V�=�k��c�V���DR	�
6I*�X,�;�~�`{�˫ ���8�)Q���V�=��X�2��X}��G�J�4���yU�/�f�=�u`w�ج�{�:x�cl��r+�f]X�+NtĴ� ��T����D�ap��,P}3�y�ի7[ֵ����l��t�}z����Yg<���C=�E���n{Vtu��AcCeG�1�����c��k��tѤr:������[��s\4L-�d21�<������rfd�*@�ۭ�֜l��B񹹛������2����W��k����stuōk��B:y� 9��JX���Q��n�m�8���m�Z�Z��_�&��w�l������^�O\k%�����ٹEz�Z���j�n���|�wɌ�TJ�ӊ��+�}�5]��c�;��V�̺�༩�eJ��TB��J��s������ ]o# ��U`|<�5EJ�8�����+�f]X^�;��`{��X8Ӧܩ �+��%�{�b5��Ë���9��~^b�E �Pq�IU~����=���{.��d��
�U]��J]��˕t�ո��G�\��ې�y8�5�[N���:;+��Nkqt��r4������J���ü��3��9�RTI��|�{�{[ڜ���
*��#(�#&mc{���TIE5-b;Rv� ������L��J�#;0�d����x�\�RU{~ܺ��b��<،�Ԧ�8����;����γ��޴��~�J�#������G#�jI�%-�3����%qj�\�T�IIu�,�ͮr�Y���n쪿{�|��玁鸤rRm�DE��۱���.=+1ǎ���;��`�s��G�c��\d��Y���s���w��崙wN{��N�r�����_fd��Q]�ͺ�ץU��ˮ��� ��G"���J����w��D���J�B�V/]������N���Whn�iA��;�O*���Þ��3��_=�۬��q�q�_�캟fe�n��ý��8��H\��vZNE�|�/e	�tr7d���̫�k�=��ZT�[�#i�I�\�Þ��3���}<�;���^x� �I8�)*���_��r��fkӝ�ͺ�3%mr��}���6Q%D�#J�}���Y���{���w���~�ڎ�qҩN1�V���۬��U~���(u�����$ AiM�ñ}��\9��ـ�N�r
�]{3%V�G9�'���s;ެ��*�IU��D��{Gm9���)y�[	&�����J�\͎2���mT��"8ܑ�$�W�{.�������W}�Xs�;�C,�Dv[�wxwޞ�y	�q��g:�ELR
.��	��%����þ��3���<��x�eG<���[%�k�ް���þ���{�7�!y� 	'E%U��˯{�{�u�����\z���Q1 đ�����YV�5@US��b3�g���n�Csl���t�M��9.�;W%�,Yv-ū��� !{���;9�����ьue[s�m�z�ڶ�:ʐ<%٤1�8:�������A�+��"t'��kg����Ӟ�{����:�޶M����`�0�p�j��׮���n����r9���Gr.���v�4�Z�����nڍ�n����]��V�d-�q\n�-
�UU[�-6�Zs�qq�V@�B���ն,�8Ys���Z�{b4X��vm�
�����������Þ��3������v+�2�r9j������{�;�O*������e�a7W�$�#w�Y�r�3���Wk��I�#�8�F�%U罗^�<9}ｇ=�Xs�;�C,�Dv[I�K�;�R8�Roc��o{Ց�t蠩�.n.6�D:��&���a��Q�N���]��ClU�
j�$���8r��˯�2Uw��o9�Wk3^����֓��8�Þ���ic���0�9�o�7��U�}�u�!�"�H$�U�]���^�<+;�{{ް�<�\u��iʶ��崙g{�a�������~�ڎ�wVK��U�ｇ=�Xo��a��yW�TiTx����Iٞ��Q�����AE;vr��u�z5oe�(ƹ굹㥷��HxZ�M�7w����j�VGz���,���)$��(�Q"IU������UTfkә�n��{�}E#�t�ֆYv�추��+�|�}��Õ_���uh�m4&���:����&�~��x�e���*��Tl;T��of�X��Hh1�'��X$�ê�����Y���n�(UB�r�@���G$2��m�SAe�d	�	�[FЁh\}&��ca�E��g���8&�d�J�A�o��h4.Ú����A�ZyΜ3X.��΅zRH$�L�]�y�(aҺ$5�s@n��4@�y�l��h�t浣Jq%"���:�o�Ie�d��iѤ����B�B���$1(!K�������X�����f�\:��-�*#��/pN�8PX�Rv'
N���3oI��n��Y��t�P� q��J���U��n�w`�Wn���c����C䫎��^k]�$B$HL�V5��K�.��Af��o�MW �p4!	�l4��BI���s,CZ,F�pꐈ	۴v?T��(�BO��"���z����(C�U�) ��D:eP
�M�/���	Є� �,��:��߽��)JO}���R�s�eaBըl��N6�r��������/R���}�)@�w����臒d���ﳊR�={�X��ϵf�f���9���)O>��R����}��ԥ)���┥�����)O��{7�QG
J$�b��\I 3s�5�s�V�[��[''a�v���5�1cG]�l�R���}��ԥ#���┥����O�ܥ)��߸qJR���j��p�|�).�Ӝ���c�V�)C�~���JSϾ>��)JN}�}�j�� E5T{������wnǽkZ�pR��>���ԥ)��}ÊR����pz��=�_}�R����Ͼ�bnBABۻ��t�(?�¹Y�����)JO?}��R����ﳊP��}:
����X�X��°(gR��@~N���~��j
J���?_4Է�ky�f�ݖ��)JR}����R��q&�#�4�#��%|�q|�H�"��3�N�:m�ދ���_�nM�blK����h|B<ln0��Z�7Dp]!7���{ݲ�����JP������R�����)>��~��)J^�şd|ky�{�-f����(~�Ͼ��)Jy����4�'�y����JSߵo�qJR��ӥ�G�8G-�3&f��J���2��)>��~��)Jy��8�)C�~n�s�9AUϵ����Q4�|i��(���=>��)@���8�)C�~}��JS�~��R����l�-Z��[�7���=JR�{���JP�ߟ}��R��߾��i>��~��)J���Ob�,���66 �5�$j\a� �������&��Ү��m ��b�U:d�pR�K�$�M�lnױ`��u�\��<6L��[u��KOCͫ���G}��g�s�;�Lu������3]nz3U�н�.�8n]�#��ˡ��%Hn}����ײD�J'�=�ٻ=�ǹd\ާ�5�)=�y�qN}����AXq��q�n��E��3�A݀�y.b����8ݘ�{E0���j\]q�����k��a*rh�vslv9�=��RY�Ấ�N���J�����[�����3�\C��JP����)O=��R����=��ԥ)���┥'ݞ��Zތ�f�oy�˚���)O=��R����=��ԥ)����4��ߟ}�:s�\���d��j(�$��(8��y�pz��<�_}�R����>���Jy��p┥'y���5�ތ͛��f��R����ﳊR�?w��pz��<��qJ��<��R������e!���cq]sNR9�
��Ͼ��)@$	��ߺ8�)I��~���R���}�qJR��=>�c������7l�`J�Wd�҂�>)a뛏m�'�n�6�`2���]�剉dX[�r�32feV��*����)JR}����R���}�p?(�)C��~��)Jy�VY����f���zf�qJR��<��Q���{�9)��u�qJR��=���ԥ)�}ʾr���K���{4Z�3�(P�	��)O~����(�<��R�%=���R����~��)Jy����r��R�M�����(+���n�Ӝ�S�~���(~��~��)Jy��8s����6�q�7!"Q[r��9�%<��qJR��<��R����ﳀҔ?w��pz��<�����kf�{6���������pW�8��v�[ [�q
�8���պRHԄj�`����'�y���)O=��g�(~��︽JR>{��8�I��{}�������ya���|�)O=��g�(~�Ͼ��)@���p┥'�y���)K�ҵ4�e!�!�7��s~���;Jy��p����h?a1���*� >}{C�;럻��)Jw����RUBE{�u�_
����̙�=@Ҟ{��8�)I��{��JS�u���)J��︽JR���,>�Y�f���zu���)JO��߸=��O�o��┥~��߸�JR�{��8�)C�^�=?_����oY�Z5�nٽq<n���l�G�I���7\�Jt�jLpYӷ�>.�ݧVZ����f�u��Cܥ)����8�)C�~}��JS�~���)>��~�Z�����{�,�ˉ7c�$��IC�ߟ}��R��=��R����=��ԥ)����'ݞ��ތ�Y��ݛ��o���)Jy��p┥'�y���)O=��g�(~�Ͼ��)\��-�N2"5H�U��+|�߸=JR�{���JP�ߟ}��R��[�P|A4�o�;8�)I��_Z�\��h�ܼ+UP�Q�O�yTP4?w��pz��<��qJR��<��R��� �h���U��o-�z�����X��]�Y㶍����u��#�ɽS���iě�#qt�qw���(+����]s�JS�}���)>��~��)Jw�U�p9�
�}�*ѭ�0rR����ԥ)羟p��%)?{�߸=JR�}�߳�R������)N�Ֆ^�nٚ�f��Z��)JO��߸=@ҝ����)O��y����(~��)JRw�{��f�xXn�f���R���}�qJR�����R���{�)B~�O�����ԥ)���p����j͚޵�o8�)C�~}��JSϽ����L�;���R���kﳊR�������P�CABD��Q������?ouowv�ΐ[r ]6_'m;P�`���AYmx�xALt���jzwJ18�����םw���t��J��EZ�\�m�[q�rC���ɸ������6��s�Iv�LP�,�v�1E͌�D�)3�li��5۝�Cqɮ01׭˸�X��Z0�;\i7O]�x(�����)��ZMҚ��Mv�j:v;�X1;��=�W���f�� �)J4ܯ�U~�UN2��tB����ɧs	��K-�p紝vɖ���Ԃ�g)�/�u�q]��2؋�����~����=��)JR}����R���_}�R����>��ԥ)y����lٽ�{��-og�)>��~���%>�_�g�(y����(>��@���w��e�S�[Dn��Z����w_}�R��>�Ͼ��)Jy��p┴���n�Ӝ��(��[N�N!kZ�qJ_�9�=���ԥ)��p┥'�y���)|��g�(s�(H֖��))U�ww\�U��+ۛg�)>��~��J{���d����n�Ӝ��(�i��7����-�P�Ŵ�Q�Du�C��Q�d]��5;y�[A��I!
&��8�ە|�9A��{6�JR���~��R�?w��pz��<��a�BUBEs���9q���'/
�R���}�p��\*K����=�*��Q��0�C�F�)�pLCq�WLR��`	�H:$L!L��Ov����~��P4�����)>��~��)Jw���p����h�f��k[�)JP�ߟ}�Iԥ���ÊS�!�w�~��J}�~�)JUp��.K�����ʭUBUG~��R����=���)J{��8�4$W���aZ����ޏ�!G%�K��y����R��y�pz��?����8�)C��~��#Jy��p┥r���D5C�N�#8>1�(iN%�g���)p"���B��UW�\���}�m�����v�4fo|�)O|��g�(}����)Jy��p�)I�����JR�f�ۉ҃p�n+�(9�
�}[���?$�J{���8�)I�����R���}�q���k2�V_�f�a��\��J�>���)<��~��!�/H'��7)����┥^~���ԥ)ߺ���GٳޜֶqJT)<��~��)Jy��8�)C�}�9'P4�y��p┥'��g�n5oz�����k5�P4����┥*���pz��<��qJR�Ͻ��R����?s��c;,U\��怮w�ӄ|s�&�Ӻ�kt�/�7<ӷ2��9�{�����}�R�lR�m�����(+�Ϸv�9�<��qJR�Ͻ��"�P4��k�*�����ÿ|"\�츥�K.^f����}�*4'����JS�5���iJ{��=H���{�Z�kf��Z�o3Y��R����}��ԥ)���8�?�*�?y���R�������);��o�{6e����h��|�)W�5���)J{�߸�JR�y��8	�/�?BH9&!�b�k4����N��}pz���)~֙%�6�r����g۟pz��?�X=���)JR{�߿pz��<�_}�R���Ϗo��ћݝ�
��O
[k�EW"��|ԪۋK��`u�6�t��(R �n�]s�9D��}�)@�{ߞ���R���}�p?Hd��~���Jϵe��E�dh��浳�R��}�qz��|�_}�R�������ԥ�}ÊR�=�Fc)�)�й$mˮt�(9����r�J{�߸=H~X�S�~��)J�g���\��Ps���]9JA�Jq��qJ_�0d?y����)O}����)<��~��)A�������R�J���~~�%��[2��+UP�W�{�)JQ�Y���~��)Jy�~�)JP����pz��4��ֵ�kY��m�u�����iN�\��u��EK��r�vp���xpЛ�" #1�&�5�{��:�=;I�&`KZH#�9N��\1kU��l�-�.U�pBJ��	�:'�-Y;J�1�"�c���AoNR�%@�mX�IW�L�Ĳ��9���eI���
f0ٳT�P'� U�q=ܨ��S)JT�I(@I	��~l�#����YD̷�%J�4�N�8%H�,�Sn�]�t��@.l��v�:bT	$RV�=&C��9܄uQ�p٭oxf�W5��A�kA�ȹt8Jy�1]m���s��鵆yCD�kXpS� ��p�Lc��[!�ee���W*�B�]B��
&d�9��qZR�Wp ��ͶЩ�5�6g��ц!aJ`I�C	��B�2�8)�:!	��VH3��4�h�"p-���EkXoT����4�tw5A��5f�ߛ�7��   R�[Pm� ����Z  �U��  �  �J�   Yg   �4��N%�㱕���+pS�M0ͤ����c;k��mlQ�������*�u;(��\����fx��:��v^D�f���vA��!�3�=V�˞���x�q�R�1��Ӱ	�����p�9�c�=j|��mZ��+��|V;��qD�vr��T��"�9�ޏ4n��]�$�c@m��3�ٔ`+��N��Q{8-�k��j�X��оtKm	���v�k�̥��[<%.�����um�A�7e��[c��D\7d��g��Y�� 8Q�Xrv3�8����=��8�[������5�8�Ukp��#�ñѩ���©�F��[F�r �Kpn��m�^*�:��]r��&���ܧS�䧞��˵�&� Z�=�+�n�j�ٺ�mv{!ə����A䐥]�u���	H���۝�7m�;rv���( �t
�W)�ȡ��AI���v[-��e-���[�g=�Gv�Vi^c�������x����U�tG;;�4�9n�c�M��9A��6�L'���˞���dÙn42��21�6^l<np��d����]��ԭ�&,E�����ڔN{9m� �V�ݨ�FP��`���X�k2/(��{v8����E6E;R�NܬK6�7m4n���
@h�Dn����V
�nB��=8���j^ẙ�&�h��]*f�{uY�q�H&9�n�i��3��Ɣ#�e��86*��+�������aI�`ݞ��oV��$ͷ<�9��lT���mRQymtg�u��G��͍�b6I�z.�ۢ�vV�ЖnݧON���[$�<qU�h����s`x�q��'[S�X�\6���=���ܽv{[��;xxR�I��A;/G9�p����u*2َ;y�7lu�s�^���-��<G]����u�;BFL��y���V�Gn��c���0�;������\UuU�  ګb�~?���w^�{����~��R�)�t�"J���6� 2~S��1D���������~��n��`)V����vR7������-����.\J����G�&W$S����m���'-�7`mMqǬ=��ű�˘kWi�kn��>{��݉zy���d�l�����w��v�;:�j�$ݻip�[�-��:�c���z�Π�	�2�T�\�Qu$����4cq�$�4l��l��mВ낼�#un�4�;c�"��j��������~���-b6�^uf�n�<q�7R��G&�5K�^v�4��q��+�ݔn�j���kz��)JO������)Jw��8�)C�}�:��<�߸qJR�����Q�w�춈;��j��9����?�%(~��߸=JR����)JRy�������<�ߵj��z�n�5���R�>���pz��<��qJ �Bd������)O}���ĩUUw���ᯉbwm,*�ff���~�# ��{�w���@/�y�|��\�L;�&*��Ww_S���78 �by�=�۫��G$H>!p���4t��p�Ṻ��&��5�����m؛v�=�J6��#Nw�{�4��wo�{ٷ_��������4���)H6)N6�9U�{�:�K�a1���D�Dx��"#�=��F��@��ٟ��RF׫~��l�SM�]�]�@���V_S��f /�y��JdU\]T]�U�`}N7@]v� _4�C�9��qg��ڰ=�7��P�DS��u�0|���<����م����#ի���ɳ�p�@Y'h8ssf9�n=nW��=7�v��b�u���jsT�\� /�y�|���:�{�G"9�G����X�[B�����
D-˾��yZOt�l��o7ܙ;.I��DǮ������`��t��0�?s����r��gs@^^��7�uT�����Ww{����D��l`���:Ӻ��/nol�n�t�)MJQ�%X~J��VF��{�.�y(�q��a���[g;�;q�d�G)�m���	��Z5of�zU�窷<t��-ۙ��&;���3@�O# �I�F@9��� ��n�4ܨ�� �%X�+6�p[��M�Ѓ�o#  ���&n�૲f�n�t��[��M��;��,ff��Q�r�^#i������|��#�3����^�Fԓ����@��I�0�Cb
��g��ʰ��B����9Bqݹw]�ݸ���"c��~πK���M��>����Bvݶ�c��0�2V�f�y�i����N�j��#�}�`������W����'�z�F jm�#@��������6J#h\�6�z��u�U�$���h	{�ROt�#"f>C`]9Q��ܥ�U�}���@�۷V��������n���7h��H�S��Ww��s����`I=�;��09�@w7v���^�nR�nD����G�-��s��"8��� |��f��[��?r��<P ��}>��B��-��m��j��)ι�r���<��F�=sHq��V�����D�W�^���[Ēiz,�����еv:��#nt�]��:�s�Ѩ�鳀�nn�Z�^�[�٣+�S8kk���o�O}�}�gt[93Ŏ�}�佝M�t@���M��=�4q�'���ػ!��Xl���&3��m�C�-�=y#d�tn�f����t��f�==���ݖ}�@UFUn=�h�]�ݭ;hM���`������ۆbVn�y���{[�@<l��{����ﯹ���`�毿[f�� ���>�y�b9ȐM�n�*�m~MT�i�*q�*�����ܥH���0����y A�Р���-Ji�v��@�۷�
=��ޜ��{6��;��}����z��8�aȈ��'�{I� Gͼ���}����c\�(��UIs��{���1������2 넞� �%ȳ"l�.71�7^��
�ݴ��aj�2ٻm���T����}���'O��&�][]f /�y�z�F�I�G4��0��7F)EG)�����@��n��s����g#��^�}�ݯzs���o�T��3+��J(䂜nD��`{��t�n� "8��h	7���3i�n1�G���;�*���� ϓy�!ާ��9ȕ����D��MM����n+ ϳv���u`}���@���U�߽XU�t9�Q2Shm4AF۫�'��J�u�m��J���n��
j�_w���R�ZjSN �r]�@��n��ٽ�y��9@��o�|�	k���S�$�U�`>��G��s�z�Ft� _p�5Ǳn�䍧;�>��Ue^���s��]���x��g���x����u`f��z��*� �5)Fۊ�8z�F��{���Ϋ�� ��g��5*GR�U����mՀW>}O4�M� /��hj�a�D��[��F���f۬kS�_]˭�f��5����wb��tܤ4��r$H�Xo�{�>�71����O# ֓����2����7'z�{�ꪀ+���o�{ٷV�����R��V�Ԛ�N*$���� }^�f�ާ���>}Ot��U�{��	g�)�\���r���}�$��}��K�����U>��=��[�s�P�����-BJ�q��`�n�����@����veu=�`����߿]�o��F,���PO���O\�����7�)�N��Y6�C=��������N���I�.Ir�5��`��o�}�۫�9Tۙ[ށ�7J�R4੩J6�V �M��D�O#��'�ݤ�9�+��ت7R:�qWn9w�>�mՁ�I��r��s���h��aӉ*I�nD���r���3{�<��N�3�ݾ���n��fӃrȤe*t��t�S� �9��o4��F�I���/^�fS�������5f���
ڸ���vլcQb�����/;(4l9A5��o���^t�sۮ��m�к8��9w������]����Y `��:ݍ� ���{��8���� �����g˻rs��Ƹ�o��ݞ�lO �me4q��ز�U�.���E�h�̮����k;;u��c׃�H�MyD1��m����V�ð2Ib��{��{/��������s�V�6ϞM�b����p�qn<g5�Dn�[��9�k���˧tH�m8�8�����o���o# �����F���u�}
`�pqwUru��hu���"8�'�W�]�gٻ}���*{
t�rJ�>i=�;=N�9��7�[�`��c\[#m6��6�z*����]�/�y�u����9Ȏ�9����+��WJF�I�qƜ��*��n�@�r��ב�|�{�R�7X�9�s���<I1�f�ɧd#v8^��v띳��{pX��Q�WG6����s�'s�nK�룦;��o���{# ���@R���G8 ���hޭ{��q��$#�`}����Ns��0���8���kA��a(��Z
6�dM��4\1ͩ�heX�0Ga�/��(���X�ߞh7�����'eG27)�Ӓw�j��`�n�O�\���I��d`zT����qN�����$�&�p|���<���"+�皬���T܉.K���O# 9�s����� �&�@!3���e�)�)��T���9�eg����B�5�J�k������~w{ʘ���;5E����7��i���o?s�#���]Xz�ָ�Ei�R�m����0/�ހ�yi=�s���䉏�]((�PR�dp�?/������VNE�t�m��`�m�o�� �闊��� �6l�89���hq��D����5	��	PD!�7
na;��7���h4B��(k(TC���8
S9�&N�
C�2���$�Z����]	�B�k|!&c10c��TC��cu���.u���Q/A���34��\0�+a�!�d)�u�]��J-��!�J��'�m7�c9&�,t�Cu�����!�LZ#��"�R��^1���Y��#}c�޺�p���$��8�8Tф��f�̭0X���Jwc��XY�I	IAAIL��:03I��Ռ�a�Fć0�&4g-AP��h��PQ��ȇ�������@{{W�O���������ث� UO�N�Ch��� :)���x����v�HwȈ�(����~����y�T� �RJr�QQے�@���wn����@�ͺ�5o�g@2�n��H��$��I��y���@����}�բ��)9J���s���a=U���1�P��62U��rx�pe��w����M\QUwy; �y�����G����k�E�n��@7
��"8�qrG# r������6����3���V +8����H�	r�@�ݺ�7q=���s�G$���0O���giI3.��9%I��9F�����4�5}��o��Ja),��}��G*��{����Fڡ�Nw�nl��9UZo�g@��F �Ot��s��^�z�J
������hͺǳ�v���Ir���9�n&��n˵\*
��E��n��?~���� m'��F�ڷs�(�pE\U�U�s0n]����`��@I�,[��ҹ\իtdrF�I�0 m'�Nف�D[N���0�n���*dnS�$�h?Us������0O��za7��6�� K�*�)Ir!9!`j�͝�r���W#�����{�~���0��G��"���߻����U�ql�mP,UUX�>ņ�R�V�y�㮬v8�Rgc{v��\��.�z�\��@h�q��iݞ���*�)-�r��t77��w�}���^��<�\+��5d�ɾ��.�(Xm���M�m��8����&7��y6�0fyl�:l�n$ �'\sp�n9�`���m��-��ٴv8���g'u���qպ�:^��	 ��ܽ��"ݿ��x?t:��*��mH;��wWQ�,Z����+�7=;cr	������J�����]����8�au5w2Fef[�_�# o��ճKV�l�X���4��9%7����G9��v��Iށ��FDUW �ј1m�q��z�f����#��Sy}ot�3�F9��p�5o�d�f�Ձ�{7����+ٳK+�����r�E�yzM�Ȉ�!���d�jـ��f΁�����
��㈦DNV�Lh�������/v�pSp��M��+GCnH�#��N'*���oz�f���l�*�΁��u`w=�"���k{몼���sG�^/��"A�<0	0�H��*���?�㾷�^��˫wٽ��5�D��ӈC�H^L�i'z$�F9��{�u�f[|<1z�֓W-��əz�GUU^��,���T��G+�W�9RL̸M��%)�w۽�ݚX��6t�۫��>�f��IN�.)���ŋB�2v�7Uƺ펒��Q����0�~w{�먭5J�8�T4�m��ݚX���@I���"8}Ov mC0.��칸���0/�ހ�y}Ot�6���p��۴2TQ����ے�@�ߏ�r���ߺ���T�3,�HR���� �0@��>Pz{��OŁ�f~��V��q�(�pNVl�ݧ�[�F)��u;�9I�����)')��A��rw�{vi`���>�zM�`�=���T�j�tl�te�Qk����9+����nz��[�=�̫$�����ˍt0�I��zM�`�=��DA�Ds��zp=[KP��$�7E\�s�{7n�����=�:����ӽJ�fe�Oi�Ԓ��U��������uXW9�
��͝ٻu`w|-m-#��q��t�DuSs�9��zSy��� ��a�Xj�JHn^�R�w������eiWQƛ�N&�\�z۽��#���ّ��t�nl�f�М�S�6�r�R��'�
�Ӕ�};;[�Jɯj�m^�����u���
�N�"��w.tf�Ձ����Ǻ�Dl�����@z}���..�wvsQq�I=�s�1�$N���==��zSwW\�8}��*)	G ���;�=������:�������\qO�)ʒD!��V�r�j�7g@�n�X���@�9�r��uX�VR�h܉SrfHˬ��:���=ȏ&���'^��_g~����_�����Y# ���ۻ�ϻ߭�c��m�n��UN�U�̫B2r���:�g`�7:˲�,�౥�	��tf"���.���`��׃\�듬>Ns��g�9����T6.AֈJɶ�n���N��=�0�#�z�ls��E������Ҵ�bk6�����w�c�\h�]:���;r}��q�W10�z�q7[�u�1�F�#PM��:ދpp>�<n�s��:B�/�*�0(/�thBcN��V�6�g�������,i6���c��h��Ę�]s\t��Ur��w�V�wJ����r���ǺU78��w�u;f�.�e�w��#�����<���((i~>�{נ'��>��H�"9 ��r:���6(�m8�>Z����=�4��j���c�VW՛�H�D�q���ws�q�~��*��}�����}�r�*Ȩr�����.�6�/���R�I��B�B�$�@�� s�n��l�>M@2ܺj�.�7d�c�[�:��l�n��j�;��M#�6�0����������莸�*���4�np�&�4�l�#c�UU��w�z�y���D�R��r9*�;�����d�T�?���>���/n��M�DDr" >�JmSP���"�;��=�4�7ٛޟ�U%����V����tX�I,[Q�"�$wv`DG9R{�uE78��w�s�ʮ{6iewZ��8��6�������Dz�����~0Ԟ�Vl���M9(��r��"�gl��Op��;q��m[lY�t7��W�+�{���;��!"���*��������0Ԟ�׺���7j*��u8�Tu���3639��'�]78��w�r9 z�mk��HJ��	�}��������^�`%�ddj" bT���I�(d���!)�	�!)�`(*@���%(f!�a �hU� &D��%�% H�*!� ��dH�h�&XIOB�����;��ޤ�����Ė�}v[V�i8D��$�@�9�U{^�5}���f;f�|�����G���*�䒮��V�9�z9�Dq'l�I��Ḿ꯵ei]HpN�R&�i�#M;gM�r�on��N�S�`4��9E�GQ�����_[|�j�"�\��ٳK(734�@�=�t�n��X�Ic�H���QJ��I��9�r"y�r"$N���==��z�v����KX�'`1�ӝ��np?6�OA�r#�"~�F�߷@~���ڨ��:N+UUU�n��^{��9W����uZ���1�$����+� |���_>���l���`����:���=�G'��s�m�>7��5}���}[�qSI����2*�m���G)\[=C�g������ל�-�RN���	*D6��sٽ�ǻ8��wȎh	�`ևwpL����I�nN�c�W���+��A�{���?z20����r9�L�q�\���\9"��UJ�������۫s��7���@�=�`Q��)�D�"��2�d�"S��0 �S�n��M�#��5}���<�$�ƶ�LQI*(�Xާ�U78����M�`��=�U&6�M�m�u4�kA_Z�A��w)�:�$��&��� 1��L�����Gdwۤ0'[sfhޖ�I�`�>ձ��h�.喁
'�Lp���-�2W8�4٭�gK��9qz^q��N����V�O{��,q,,lF
��¢&0��o��o|s������YccY�I��Fh5�Y���-����St�L��u��k{�w\rt�"��)�J��)���bI���$H�Rh��!�s���,#��Z"7F+8˕cc`PY�[x��96f���a8����Tr�K��p�A%a���;�h�����3�8�Db�����F��$aM�aaM�V�2㌘��`�X�׃6e��ae�׼�eUmEF����w.������ @���,�� `�M  -�d �8���\  ��  mK9���$܄�ͫ`퇋�1��[A������q�έ��pqcf�g.}9�V�#�v)��3�w.���k{j�����	�����k�8�>*F^�ݵ��n��n���glk�E�ç��a䴑Y�>ȋ� nw\����\��=bL�m¤a^q�Y5�K��ł�tC�]��3-(ɞ�Os�����U�vp3��`�;v]��7��I�؞���=��tvR�ۣ���b#W��iís�:l>1�a+�������7N��n�P�y6��.y�9ò�l�غyJ����	5ۮ�n��pI����3-��vaS]�/H���&��mاF˹FzN.�`���LC���)���c����pÖ��#�Zqb���=A'�t�UA�sFڞsS�
-n�Iz�b�����٨�\��W��x�� ��Q��kQ-<�.v�4s�ML� �;u��[1�A��a03Ժiôz㌜�N���Ͳ]�ny7\�a3�q���㊫�׊ujy�Fq<�9����дSXㇸ1���WU�nշaϙ��C]beUgfB��+۲NCvk�6���H�-R� &�=u�Ǚg�6yr�:�C���q1
]3���Om��q�v��6�����FD�s˭m�k� W@���\��݇`"y�Q�6�W��Xݝ������\g��;�W[=��� ���s�Rm[�M�x�I��J�FS���ɢ���t�E�c�Mm]���X� e�;vH�:��^Nh�S���=�-�Ybm������<u�hx��'��[m���q�۶�7 =cP.}x �]g�y܂���ț���;�`!p��n�lm�C�|[��.[n�v(�t��z�@[���>S�^��^W�����[(�9(��nE��f�*��7lD솹�-�s�pGa^���g��V}�'=��m�N�e�iC�[�  )�ֿg���w�{���Y=,�,�I�3?���`� m�����"> � &�؈:DO��M�=���#��y��Y��V�.�Z���H�Z�8�J⭕��uk\q��q��p6	�9b,�.^ٻf�A��u�tͦ���v�H;Y9�
0��ͩ��k�R�n顷N��m����q&{t���n�Ӌ�� Q��g l�x�����d����w+��;=Y��Mi��p8ܓ5�Y:9i�[F@� ��0����6����Y ��/b�{ߝ�w����x�|#�e�uN1A�;I��{t�����'�sVM�4��>kf�{�܎�},�F�N$����U���۳�G�v��
 Ҩ������u%���Y���qK��5s�}?u��:���>����M�z8R���t���L�\��q��3/R^���0ު{�%M�����@;[
��)QAȆ7*�+��}���Ǻ���}���9\�{wn����")ICR&ێw�f=�`|�����۫ｻށ�������@R��>"6SGI۬s� El�����&��9`�¼8�ϩu~{��i��k(S�!7"�<���N�/n�����n��u-ך���o�5�#DN4+�o\���Ͼ��=�0'r
�5E��u�v�����\|��^��$��(�9*F�X}����np9�O�l����扙q.�ʀӉ';�3�H��^΁^�۫UU}����6#Z����:N��>������u�q��}�[��np��j�B$�D��m	@�Bd���Fǜ�:�v9��dR�T����r��cTq=O^F`ڬ��o# ���{�5MϢ"#b#�<����_��Ò�%G")7*�����78��[��o#9�D��vIĤ�GM�;�3^�>_{~���ٳbP�� �$�%*B�qA��B�9���w����%�6Y6p܀�q9B��G�ٻ:f�����f��b��,�4-�U"nD"�;��]� "9��O4-��6~��z_W��7RJBR:)5M��(��3�f�N:l掵��X��_�o�v{�� �����*��@�S��
[u�l�ӻ���@�ݺ�>�YKc�BN$��@R۬�9�@?4�@M���u=��ɓ3���ڨ�㡉�`|��N���|��9�ߺ��
[u�8�$�bn���SS�^^��y~�{�2)m����;� 2Q��vd�鴻�"b
0�@ͽ�ր�"H�u�l:��hBaޝ�Xf�j���sF�%B"ʾ����{}k��o����Ò���D!�V���z-n����&�F�DuK�I1Wt�ٲW�z{m�'�F�.��h�ey8��b�ݫ']^�-?�����_}Q���ƔI���� �~�w�&�F��ot���n���)�*r;���gR�*�9?{�z����� 5%K���܊���w:n�Ձ����NUs��[���}���<�$�댑���C�� ���{�)m�����@�r""n������[�"q$�z�����ހ�y�u��y�Ȩ#�s����kh��i�j�mUT9c�{�#�Ġ�Ud�\\����sq�m0��V4`L�����a�O�u@�v�L�3�3�۲��a��|�:9Wn�v0nrU���":^2�wdtT�ێ�iv���Ƞ)�V�#+�u�'o�]�ۍ�3����[73��S���\�j�4;qm��$n��ǶJ�����^`|q�Z�[jZ�Q���,�Q�����j+��w5�]v��8ѻ^w�@h���s����#�n��1���{Q5u�vz��&�0��{�s��p�G9_������^���RTܩƚ���΁I7�����Oۤ����߫@���׿�9<���_�~�F	��8�4�X�7۠v[u��.Zu�$�F��*

�jB����#��Ғ�Kiހ�wV�{��n�#��8���s�N��Go# k��ؖ�`u���R���&�P*QJR)���E�5��n ;�퓯.B7�J�l6������@��}}~ �y]Ot�n�9�@~iށՉ,l�:"rQ#�`n{7���7����DA�Ds9��3>�V���wM�gꪢ����`��K�rH@��۝���V ���	7��5��@]�L�Ș㡉�aU�Pg��`{ٗV�{�<�u�_W�bDu�ƚ��w:M�`Dr�y�v[u���;���f�6K��y�ʁ���}�y&�Z���bl(�R6Z�NV��msóE[MME��=�;-���U�"9�w�.��3٪Q@�(�j����<�]g���&Hn�����ϩ��9ȉ�Uq�E~�S�#����͖fg�{�_|L�f(��Y
x�ڿ�s��w���� ���O��"��jn.fc3//@�s��y}Ot���9U�R[��`�RI�QS����*� �I���r۬ _%xId`g��8�"J �(��R9N���W&��5���#��_j��.�И�a)�F�h�������n�|���YȈ��f��{�ȍi)Ș㢆��2_�o#ϥ�n�6��"#����ت:��"�uێ�@�ݺ�7}�ހn�� Ͻ��>�R�%:L�HnV#���{��x ���9��Ȁ�9�_*��*f}Vٙ�Q�#�8�b��v n�G"b9ȏ�w�6�F�=�ށ�Xi���	�5(E�f�BNTT�n���'kL]�rq;]�F�6�Ji�b�K �{%���u`n{7��r������}�(���)R$��&����͙��@n�WU稪UG_Ͷ}#��n\�f$����m��>i� ۇ��ĭElQ�DE#nN�r������xId`z#����@K���I7˪*�*����x�"9����<׿u�W�}��W��(��#�$x�;�w���~�U�d.���Y�괋k�:�LFש��=1��qѶsKڌmY���<�%��-&m�u�i�u��Ւ�䀗F^{Q��:sn6����*X���:����'T��ې�6�s���q����9Lt8�{h�s�e0��l�Ƚh��k�]����9�,&96�q��Vtxt';�q͸�=vs��8l��X�G��ӧSU�{��=����w���e0�s�gm뮶��r��vR3�Q��dٻN^UE��p��:�Ӯ%�몋�&�ee�=������ �w����{�,��Y�`�E$:��z��'���V w��	B�e�s��;���B(��GTӝ��w�|��	%��2>�{��8d��M��)#��̖feՁ���z9U�j��`}�kr%#�D�]�e����>����� >�+�>�2�R�����l���B�qx����ΔK�B�\�vŠ��\t���������G�f������X��^ �˫
;�BKQ�F�#�9;�5n���� �#ʵ�o�w����n������=�lG撜��:���n� I,�r"w���X�W�j* F�1:u֮�@�ݺ�7�Ǻ �w�舎��u��n���������� �z���r}���@>�w�$�F ����Ț����	���ۍѸ����wB]	fv�c�[��\�&{cx�����w-@�(�*B&��/��������Id{��9!䟷@��x���i�drK���,�s��̺�7���@3we�w�,�[qS�D�㺲 �y����r+����>�UUEMI4BI$O�ϰS��&0b��*�L2�we�Z:o��sL[S4gz�,�]��V�)���N�$�\�e[$^��q�p��%�	iН)Hi ����a���l�{8y�ݹ�FҌ��.��)ReQqH F�t����]�hn�P+�t �|��)���c�KX:5eP7Q۫1 Ճo0�5�,�5:9��A�ldk[3FOZ8u�����k�������K!ɘd)Q�R�	�\-C��2^�h`- @aH�g�DDD�Sbs5���UZ.��A.�Ե��S��s!�IXbM�]�3 ��`6aF&b��٭���69�3Q��a1��%�@21���0�m���!�X�F��Y�n����fV��6�(ѽmv��>���uU_����RI!��?��Xʥj���
��q-k,ܼ��1��M�Q���6���ʊJ��Т!�Z'%�Q�'{�����&���1��H�� ?�� ?� �HD$@	E1*S2%P �E ЄT����4V?��t: �x��T�%�ڋ�>��J��+��=A4p�����,[����*�<u))I�����Dp�DO�~� ~�� ��*�=��Vw�j�QD�DH�M��&� �O#�ց��F��=�>����e�ָ��%���'[U�On��0�n8����r�oP�#��!čmyt�Ӷ��6~J��Y�S�s@n�ӱ;�T�F�16�����۫}���7vXz���nʠ>����I��UW�S� M��6~J���0��P#j1ʒ$�Rw�s�n���}�*��}��z�%��*��UR����~G����]�ID���?%XI�S݃&F�e���������|��]��n1��u<a�t]nrn�K�v���Ouu�uƞ0�Y�Ls������D�$���n���~���Ձ��V�������1�cX�LX�6�
E%�� �Ot�6� _WiVԕ���U$}�D���T��JN(�s�W�z����9ԖF ���@��,eE'���/��]���WV���@�R۬Tnɉ����J*+g.����{	�X��VU{�ɆD"B`�� 1q��h|׻��ֶoxhX
�.�U�L�1g��ގ�N����e�t[)����2m$��y��E�@� �{FooU��k^�=�"���t=G 9Q�^�KF{bg]-/�$�d,�w#SW/���xx���W[��ֹG7��뇍ǈfڡ�ir9����9��%2[�6��@i6��pJ��Z#���7�s�a���0q:N:磒l���{�{��z���n����c3�o��Wb-�
hQSu3�+�ܙ�#���s�T�,#@�HG)��V�ٽ�
[u�l��{do# ��g�ə���!#M�'zZX�u�/{��̺�7���r�9H7�_��T	M��&�>��XWVF9ȉ�$���?V o�YF��T�$�*���@�f��_R7�7�����`uB�9NJ��`������X��V�Ց�v���F�i��F
QTJN)3�\A��������Ua�g��l��3��F��Ԥ�&N�[�������]~�Uu���ށ�4��Ҍ�㡥"�:���s�@��daD�a��r>���w# ��{�'I� ��b�"L�Ct���D�nmՁ��ozW5����`�����d�luq����'��~�g�GWVF߷Q$�8Ԅ�6ԋ�u���u[s�6�F��=�Jn`��嶗l��x��)���wn�񧍸���Nkϒ�d�3��T۔�F�;�̜.�����9�7I����P抋�����K�̝��0ާ�t����+9TG�����䂑P�`>���Np��#�9��EWݥ��f{.��	-��Tu%9 ��z9��Np���.��Dr9��ɔ��G�j"�������?b�?s��7q�hK���P� uT�$������ˋv07��.�ף��]�&��1�xcr�ns�\�]7wJD�H!�eݮ���u�>����Np��� 6;�Qu1I�D�lnU����zUU��V�<�`f{.��9\����%��H�mU��S��}IN�%Ց��';��7�`�!��V�<�`f{,�_y��u�z��d	fhG���J����V����N�9RIEwk@m<� ��޷��I�`}IN���J���i��R�i��H�B�b#��s�.�g�[��-�ڹ� �O��]�>6%hj�U���~o����� ��Jb0��0}�Im-R��)����nl�:�U�uud`$�W9<�(�UU50T�)*�;�n/&O�qn��'1�z��ؒR6���v�nmՁ���zk�V>_f; �b�eF��Ȣ�MW�S�KN� ��*��Y���q Ln��ﷺ5�6j�o5��[N��i��������Nŷ1�k��GV]�5���1�@�/[q�ϑ��8N�t����Kn1ہ��]pqg+�U78ӗø���ܸ7��]�e�){��U�6�u�8�H��[,�c�������A�r;����W�)�<�4��N��󗃺]6K3�X�R4�8��q�nȷ6�u׷c���p�a���K�����9�H���z��u���9�`�!��xP����{�W��[���|g�\(�m�o�5{5�/{���]XQ�{k{��0�GR�n0C������`uud`��d oݔ�H�����$����P�0�[�?DL��;�3]�G����NH)��`����{t>~���U`]Yw��6TU%9 �'z-�v�َ��{.��n���֔Г�'*�z���=quA��ƍ�܃p[=a�3�Z���c�r��C���㡊G`|���g����f�z-�vW�6)p��o.jK�{�3�UQҰ*��]b_n�� 5����LIq󾘒��:x���ssvMW�'� �w��ș�Rn���۫�~�J�`�EB�����@▝`=���# $�@�����F�:��v�p�3sv0u�n�&����੨�*.o]��u�:݇lk�[nB���ݷ�ۍr���!u��z�U�v�
�%#�D�.N���u`o�w� �͖W����=IfE���U�� �I�
Zu�l�������n[��D�N81�ށ�s]����?~�.��"XOB�4?b��~S�=����ʽ�����z�*6��)��#��ʪ�/�'Xi�`�'�)i� �䝕*F�"Ct�����u`~�R�?{w������^�;ՙbC�JtҜS����vmf5��wf���kr�j����.V����=T�Q�:pjA1�V}���[���n����]X���ʊ��bSu{�)i�z"9'e�Հ&�F�z�����8�~����)0r�M�`z���`]Y���z7@N�� ��[����R9K�o�f��X{ط�5���߀;%3*jj�*�)&�2���#Ĵ��y����*����$#QP��`}�f��f��`W�3i��eՁｆ��I�D�n�j[�R��/%���u�σ�r�l�����M9rO0��($�JrJB��5᥁��� ���Ȉ�u=�;�E�;.h�,��*f�p�XWVFߺ��	�j�p�n�F)p���o�f��`��'8�ӻ�6Tv]M�q&7*��*��7}�7�����nk�9^�eՁ�4PtHECq�
9�t��KN���� ��Ot�s�|+�?��z) �����I!i�I"���m���C�/� ��Iԯ�
Є����6�D��B��,��eĩ�ĶoZ�n�6F�ʶٱ��Ai5�T��:�s�*Յ����='Dca����0m�m�8`�HI�w�v����I*SIgY5J�!�(hl��Z�,�P̼�DB+�e3B�v4��1�k�'�Qu�!g{�{Uv��sv˴>0��WU�H�uP!;�����Yvij�yUc'9��C�x/4����0���8�kq�4/����ټŲG��9ve!��T+���w�&K/���nP�5��7��l��ql4���/�rᰪ�:6����M8�R�+��sv�(d9u����BZj�ؚ�Uc!�ܥ�i�n��M�kl[5�S�#ZS�/3Bu�f����Y�Z1�m�g%�KY���;�v�)�{bZ��U@ @
ۨ	e����u��  �R�  �R����8�� mp  jYd�^�ls�kz�lRQnwЮ����J��<$�qn��Zj���sCg=GUr8ډ�g�qʯ���Wh�ĺۡ�p�԰�-2�cv�k����r�O#3��ڌ��3�n��8����1��ϳ��R�w��Ӟ�b^BU���[OKΝ�u��Ӹwg��O7S��\v�=Tkr���/����m��,�#N�\�P�&z�^ 8��9�շlm�Fь
L�4����)��`�����T���<�v��[;SF�wHcUY٭�������U6^gn-�#�#�Id\M��Y��ɷ��7
@b8�(�����ۨ4�u���K�D�.k�a�����������I8�Y��JlKW!4��-捵3֕��]Sq�q,�p�����m��kU�U�;�_(V�Kz3�\����]Z�{\�;mE�V��v�캮8������ö��bx&�eSԣGg�㶡v4�7m�e��̲�G��%�9�C����"]�c>:^�]-�G%�=����]vأ��X$o#o�Z�N� ���ckH�pgs ({]����e���v�� �ٶ��Þ��:E��1h�pq;��u	n�v����K�aa.���$�b��z�N=sp����<�;��)����9um�۶��NA�Q]vR�Ld���:���v.ʝ<�L��pRpN3�S�9@���z�XA�'��[H[u��m��T8���l;��u�).x��1ՓZVC��pp���Öؔ�iݸ��O���nU�;v�g��u��q�mC�����&y{:����qӉ�3�
@c�����,�`h���;u�=��A�h� x��z�tG��Pu�����64���;{t�����d�ڥ��L���n���kpIщ8�٤��q��[Yɬ�θ$-�m����f�3e�}{�x ��j���'�EM����}1AO�ѵWb��0J/�#��)��PHt*��x��~����4i0H-�@.�/&�.]�,��ݝ��㮴��˱�x�C��Ƭ�h�SXq����R�ו�ݜ�存�����']�vNy��첕�7A�S�og����'h.D�y�ex�v�e��� �kcgL��]�nR�ݶ.J����Y�!��ْ	��Hn��kb:������)�`MFp*A�.7B��f6݁.{c��ċm��{���|�9�v�Iv�х@�.��d뷵�Q�d{g�Q�؎w^ƒs��g7�I�ζf�ߣ ��� _ud`����s��DAȏ�~��g���N��%$�"'vt�۫ﺞ�	�s�}�l�#��v%R����B:�9V�{7�5��=�`{=�VۂKx�Tn�9%!9ށ��U���� �����p�{�qqt�*8�iH����W9Y�����g��t����8��J�����n�M�ն�s�p���@62.^�4]׫���;;,ɝ
�:���\��R4�q�-|���V�y�������{Ӏ}+�]Md�m�%���;��ߪ���9Fb�g�x���ڬg������Tt�"��Ѕ*�@n)9�>�78]Y�u=����J���Hj7����3=�V�{7��u� �U}�[�:)H)%��s���6�F��Ot��>�6���n�H���r�NQI�&�O�r]a-Y�}���/I��;"7��}~�7�UY]\`��@n���MϹ!��u`{��/ԏҤu$�';�7^��>�78Id`}��H��a.#JT8���U���ufp=Wʬ�(�A4�Sy�{��uW�k5X^�ڌR	�tB*ge���r�K����O۠7M��OU{ܜ���V��N8���{���u��٥���ܬ���!�rJK;sm�'�k�«'c��;O*��'F��8xیa���R�v*����Јܾ���U��v�%h�>�S� n�wpQvTISuw8��3܉��l�:�����t�j�m�R	� �'vtݚ`w��"&O{޸�:�~0�Q*�:�� �(rB�������u�f�߳��@Qv<G�ϮU׿X,
�R:��RM��7vX͚X̘X{3{�>��f���N��E7�/�� ���ۗv+���n�t�;u	^��[��Q�
�*�v�f��&����t[���ۺ�D�q����h	��`u'���`Nٞ�s����k����#$��c��=������r&S���v�９1uqqaU73%�^�{�����z��~0�h�|�Dr"'�?}��z���.ʉ(����>Nـu+F�z��oe�u^�ײ �s�7R$��FE%X��/b�����uu��\�E�xI�<֋�Ƴ!�h��q�ɍ<.��kh�뗊�	�VC��<��3��z��*��K�nc�s�:���潊֛7��:���Y��n�t�v+��nJ�g.��k:�u�{r�m��{փ�zs��;��|Fm�㳜�c����.-uA�m�ۮ�v'>kH%�v�Mr����ݵ뇦�hV���u���p,�F+X���v�LoVzļގ���=��3���>�ج5D�5�t/E��>�Ot�� �v��ecy%Hԕ�C������� ]v�%h�>h�a�S.�.���*�t�� �]� IZ0�I��{Մ5�)ETq���,�� ���[qX�ۺ�.ɫ�,�b��4��0�I��78{�K�U�}�����N9t�%5��mau��d�k��oL�Q���ѝ��gθݎ�1�t{w�z��V��4�32a`}��)2$���꯾��g'k�a0���UC� �z���$���^$���}��a��J��j9���,�� ����s��꫄�\����sY�h�f��=��� �]�`|��m��7$$�HX}����� t�%h�}�����W��S�t܍ۯ4�����.-�L�3XN-��8�)��$����uX�`	+F�Г���X为,�����p��0�� ���^�2�w`ҐR:U!L}��n�ӕw߾��V��!1L�$"Dp��@yڶ�PK��5X�M,�Η��dc�����>�'�t���`	+F�s��Q)R0���u��٦ ��`}��@Iۨ*&�
�U��gϮS�[p�PO.n�g�^��np�$�!����]����J:�t���XW�i`fd����f��i�u��Vkm�H㐘���@m�3�S��n��E������X�l�Ԑ�9!`g߷�z��`�ـ$��	H:,�.��j�C����X��Jр�=�T�uG�c��7R]��k欸�(����v�&�fL,��x��@ջ���}��T����6'%�N��7�=�	�ch�7�!�k���wV�93xZ�VM�D��S�h�f ��{�9m��ɴXW�/Vq�! Ș�B�o���� �� IZ0�L&�RSN�P�����u���fL,�f���P����!�%� �� IZ0�S��n��EF8�T��΁��K����[���M,�e�P�t2�����Uj��5g;����Sv]�+kfM�:7L�u������`�(å��I���Y�n
�gs0\t�F-�ln�\���e,� Zۋ[��yf�u�m�"$۫nQ�8��c[���Wn��r�hg�t`��z���A�9ܛbF��ˮ^ �ݵ2t)�����-Ҍx�y��e4�����������p��KpN�(YEW�j��X���h�N݅�:K��צ�-:�x�p�2�&�;�����U��F�d�T��2H����n���� ]V���ݳ�Z�3K�0�*FI
I����=�K�����{7�ެ!��j5#T�mŀ.�f��ч���D��?n��z�`^��H'*���l��4�;���@�vi`g�i`w�:YYƤ�e8˚&.�WS��～4���;��,����E5NF� Tc���Q�:��m�z,֞���ݜ�-�� 8���Z�hB�8�,&j�t��`�ـw��`��� �+6�%Ecc(�`g�ik�΃���(��T� ��}/�.�3{�>׺��*���W��i�q��n��~0]Ot��}^��;�u�6�25$$�Ȭ6�ۛ������`g�i`{ޘX����TH���U{�|��V��� _$��߮���~�������w��{\�&�����β=�+��]�1���7[��$�70T������ �m�/n���+7vR	�*���l��4�Г���� ��Q�c��QDܦ�(Ș�,�3{�5nk΋�������l6�e�Jc\η_���U$�j Č!�1i)"�:!�bCKuv�~���2εY�h�Tr���ޏ 6^̻Ɛ�.�
��w�D=�1��y��i6p��qS��!�om�7�l�c��B�u�mGF�7����۰��v��"��7��h����35�+	*<��xLX���/B[�"4�u�"�𝢚9�Ta�9AفT�!Q�e�ØoFȊ,;7[���J:;��!�����CV�j!���^I�|�����ڋ���9D��:
*���@$hó��,��2�x\̲�wJ��f&���+��  ��@|T�;n� {OQ1S^���>�}�L,�shD�"��D	I��N+ i[0�h��'� �Y�q661%UUN��ɥ�����5$�@R��?G8�g����+�� ��q�l�%v��x�h:.1�k�'��6�a�G�m]�I�M��������R��@R��G"#����}#�tM:���*��Wq�jK۾�G929~�`v~,�2���~���TH��
M��
Su�$��@|���5$�@��!��ۨ�����R���X�۫��}��]Vm����B���!�N�%�T�}��g*�w����mAT�&�g@�n�Ձ���/�w��׽8J-���S]��E�OF���q�\ZA����n�u����(��ɚ�
�p�)J��q%)FD�r����	Ss�u+f�K# _5	��������&f�t���s�26����E����ހ{
ݨ�Q���ģ����`$�0�9��Ϳn��{Ӏ�-�RN4�� ����ݺ�;��ށ��U���K
:���ӧ�&⒪��0I=��� I[0�Y>�(�bi!	b���I	�TF`�$F�M#���zw�'s�)!�v�ΐ[r���;�΄䀸9�f�l�8���s�g� un��<ݜ-�@�4�;d��Y�ӻ:�(��K㚡�n�q=O'��8���16 ��l��=������.2��x:�Ñ��R��9y�q�L�y��FKp�OVዙ�J���ӻi�ga,-�c��ݬ���Y΄������۲��ﶮ#��d]X�[{��=�ふ����9�q��=Yu�����p�ێ��uv���Mƥ�uÙy��=I��[�Ui �{�Jـ|���z���!���mP5%+<�U��K#]Ot���$��VM͕dQ���u���j�{�T����X�:^x��)J2$ӕa��UU/�~�@n���i9�>Id`|Ӊ�ڒm�B���u�皪��3.��{�3ΰf�7#R�ʈ���R��9��ɩ����Ɠ��{[���'�����b�'#%G#PlbQ����V}��� ����Ȏr>������>�E��V��ڷ��R]���p�����U�k�Jn��Np�D�&�EZ���SrU���mw�b��g��[�+ۻu`}��T��6:Pn8SL��~�DD�~�`S��$�0]^��6���
B�I��y���3/�sٽ��u�[��hnE)��'!�l�a�n9�le�c�n/;s��˧���n�uU˺��ࢃ�*�r�@�ݺ�;�Ot-��6A�~��>�Q-�3Ww3P]4U\`�����Ds�2z}�V �?���̺��P�3??ԑ�	�I%w�@z}�V �J�`�o#��G"9�m�Ձ���z�V�G*)�cQ�a�KV�8m�`�����V .��u"|n	�"�k�n��Xsٷ�9m� �I���s$0]]�oluݶ:��wFN]����$pmg�	rqZ=�J���$���N��9��I]��?�[u�%]s�$�F�\����E�U]YU{�9m�{�#T�8m�`�g���_{
�MN(�B�G���' I,�WS��n�	's����QW�6�t=�������O۠9m���'�t�`ڌ�H+$�B�,��#h��4����J!����r���{����$茉�ʰ;���@ջ���5X��V}�j�BD�'	ۖOn�]�6���Ƶa�&���h�5�ܯ���2qG)R���lI%'z��vy�3&sٽ�i[���j�Jn���Np�� ���@r۬�f,��t9)�W-tݚX�f�Os��	=>�� j�� �)*�]]]�_.*j�WW�M�r۬�jp=-��`{?$����q���M�ށ�w]���#�ԿN�۶`�n��G<s�̡�.	�3�_��ի6oZ��3p��uP�ct�cM'N��x�f�A�il�=��bm�v��&�Y3e]��Ŝ=�j1�<��n/<Zz�\�۞'��uiub�`�lM]�{{54u�*�1��W\}�:���H��A\m\�a�j:&[�k���aq&w[6ݶ�'X�-6KXvu�b��q��69m��I,R�=�-v�q�d'b����'d�5����t�j���{������u�u��,���Vέ�#�m�0���;�]�^pv-��qk�':P��q6�S��#U8��?b�V�}��s����`��&�K�**�F�N�۶`��`�5X�d��rD��1�X��w@n�����%h�;޺q17Uw�㦁);�7^�7�5X�0�3�f����QJ�F���J7���� IZ0�S��np��T2�6>�4!�&z�l;f���-�:�{;z��J�eF�^���}�}u�s=�v���y�6�����78�'8ɕ��@�G"s��>�o{�}\�����D\���>U�8Jў������O�	�Q7VEU^��{Ӏ.�s�,Ʌ���oz����*%�!P#��]�� �V�WS�D���X���&���+�|�o'@M�0]Ot�u��J���W+ٖ�h�n5|N�ӻn��NK3ش��Y7kr���$^d<8g:R���*Ԁ茊���no��[����Y]A���}���F�$�bI);��p|�����]X�f���e5���(�Q�`g�j�]���#�� Q
����I|��� 31c֢O�J��+��n�Ձ���@N���{��O��g �G�w57wWe_&��0]^�܎r�ޝ�~V�2���_W��ӊ�n	*����j�s��yn���5�4v�$��]���.�{j1���9%)7;�3^�>��V�2������@>��[N"t�*8��N�Id`}��@N���#�ɓ���rE����\End���F��O�5��=�`gՒ��n�Dd����ﺞ�	�s�}�np/��@DH���]	�Ay��s��}��m*�������@�f�>�78R�`}��@}o*$"��
�6��&v��g���Pr�mt��6�8��֝�q���+$������R�!(�V�{���K# ��A����ܺ�S70]�WqP^fN���a��Ot-���=�`uX��jE$�J�>�ٽ�
[u�Gݦ� �V�S	%�4�I'&�zk�V}纬fL,��oz����DB'NT!���{v��u+F��Ot��?��s��j��$JBD�'��/�^Y��S�B8V��t��m`8fiʐ���xk���"��޶h�l�Ǵ��i:�p$s��dP�a����2��t��
�WP5Ь�*M	8t�ob	���Л����ѥG�K��=���"�sf��&m�٘�V��e�����{&�k��e� IN���5LEFQ`y��{7u��ѥ,��􉘉�ۂ&&�6�9��餝��n L��zc:6�͡b��bfo��:G(�2�� �?R8���^5�ȡL%0�+6v��b�T�+����P�Z�N,f�<!y��I!zB��e]\:���:��dO�&�5�9z�Ol�   5��[xYRۭ�n��a� ^�Kh  v���@
P� ��  AS�f5t��eM�`�k���m�TJ��4��n�r�cs�s��ӽ{ػ8{`��㧛�wH���۵u�d�[K���^=&���� ��J]��⪡��a��6����nNN�]����[r�ph#��`��	#��ɷY���;���.X-b�{tn�)Jܴ�(�I��{�b�r�u��i��np��t���g|��Qv�v��']�v6�n.:u�!���U�ڻh����p.����"�/k�&λ���z�Q�D���1d��4c��K�V�3K�kO���:��H ���P�'61�8�Fy��⃶FUNWn �9���s�uN^�⥉���y�;�i�:�V���{nW��'[$x=�<5UrK2ܛ�3�����T��q����C�١n6�;�:�+XC���<��W-���۴�d���;��`�D��@�<t�q��;��b�Y�9��͐m�Y�|����V�ZwY��3��[����v6ۆ�	�D.��^zg��n��n�B\�8�"Z�iz<�P�Bn/i�������-���'X�Za{k�ˮrH�':�i�sUR�a`g0⧲�[�2;�1�۱v���sQZv�%���'BpVnCe��5������Rՙ��Z�8�4f,�v�'Ad��H���R��^ɉ�>Rr�:c�[V̎��MԎ�a���U�Zv7Ht��c�f뗆���mW9�Ks˶�qˁ���j�ɸsO
�!V۳�ېM��;��;(���ب��Py\(=��燜�q�(��lf�������ro���le��s��v�c��Z:��xm�VzgkG��C�=�8׃3F��˳��:�9�<��8��n���A����f{FB.r�\U������U@U��Jp��t]cn�<0hط:����Buݭ�ec<ϫm�4p��6� �Z����	� O� 8hU;E%O��D�lD�v�����(����������UOx��׻�Z���7��(
��)V5�,�L[�E�E���e�u��;^tz�vnhb3�ц����������ص��ݳչU�\�l�y��d��^��N�Ξ�bWv���3:#�k;����KҼ���+�j2�n^�3b7�uɲ��,��$��r�0�c��N��5�d���:��Wv[Nm�9�-�t�4��tcq���Ր]�`غNe���RK<
+�yq��J�[�	`�g�ug�(0g�&�㞻o!�VC������b��J�� P�nGRr�]���;�}�S� �� �z�`�W
��茊���>�ٽ�A�w]����=�0����9U�}��~A$)(�RI7{�9��X�'8R�N���@3kJڒ�$j�i	(�3�5XT�����
[u�ԥS*d���j�*&r�t�����O�|�{Հfd֬���M�pA��a$U�ܮ�7$�:4�絇��g&0�|Q��7�|�g����n5 �n.�������u�纬c�Vf��$��	�I�ށ�~�\�	ؔ0�6*���(< R��ǉ.z{�\�}���m��W�DB'NrDG���~V��+��~�@Ż��3Z�҉S�F�N�	�s�j�{�)m���տN�������Jp�$Vu%����-��i9�:�)����r� ����Ѥ��OD��G�L��k�0���z��s�t�ܔ(�)%�U!Iށ�w]��I�T��A���'qwd]��m�(8���W��\����?w�۰��g��!��>��x��.ˉ����̘��ޜ���2���"9젃0������c:gLh�� 1hN�}o9���\�������T�6�RqFⰣ�ٛހ��X��� ꤧ �pLˢ$�|*J����@R۬܈�>V��	�s���ٛހf�q!)�1S�mR�5�,n�/��xsN\�fz�չ]�C��54�1%"N�䈎;�~�`{�VPoٛށ�w]��݈Hۂ�S�����=�=����{Հok�'�d�2P�S�8�7�Voz-�v~~�`{=0���f�J�)!IER�����ɟDDDK�?V@��`]Y\x�K�Pe�ڊ_�׿{�W��6��	��Q�`w�ج��{.0�Ot-:�>p�8*j.ʋ����׶�]]W�y�cv��n8��<k�j����m(�k���G宁��uaF����A�s]���+���d��b��������=�r9��&Hs���>T��@��۫��Kx��7$���d����=��r&SO#u�n�{�V���'JrDG��?b�=��V�����u�Q���@�F��B�r�@M�����Kn��%1�c��HH1`���6Z��ٺv�.t�������>O�j��mʱ�[u�Н}���,���un��G�%��Ryŋ:�:u�V���lXb��ݴWn��um��Aց�흳�l���8����aɈܜ;�c���&�x:�K6�6�^���܉��6ôs�tlbṸ��ۗ�A�׳��s�c�E�ܝ�Ql��"�ۛ&{n<p]k,psq���68q	�E6��l��V��ݛ6z�؀�#���t������q��ܷ`9C/\��Χ����ޕ�����њ�Kv�뛁�ŵ�dT����۠)i� oe)�+��k���֑$)(�@m9ޔ�5���&O�9u�&�F��=��!ȇ�O�$%I��bJ8������=Ԟƀ��V oA�T����.��̝4�0���
Zu��G9�ꛪ��Y�*��ԄS�7*����
Zu�}�P��:��0�Hpp����x��dj���c��֎�<p���G��vq�ns�,<�Di�f�f�~~n����`�%8WVF ��� �a�ëm�j��1%��y�H]�UP�F ���KN�}��`���*�J��/+'B*W[��ɽ���"&R����Ǻ���VS���P%8P����@�� ����]�`A���"
HRQR�ړ���<�`{=0�7ٻށ���6���FT[���ӓ���<�77�����nK��B��g��Ӄ�*Jq�%FĔq�y�+�� ���G9�G���8�����칻�.K��@�ճ }M'8�Ʌ�]FW�rF�
���I}���^��~�[�G���5ي�
fL1*��������0L,� b��)��;�.U�za`w5$xǰ�7#���5`v�� �����7� ���]\��'D�'���b�=��X���@�y���+�MhnER�)IBR��ي7=9�o�9�c���Ӭ�m;p����_�|T*r��r-���4�7ٻށ��W��=�Vo�em8�8�N�� =���	�s�vR� :�h�;U��i�B�����'zPf��`}�H�"9��F �M�&�qv]9�$ƣ�X~�){6��3vi`~��}�G3#����T��(�C#��U}��s�M�`hf��c�I"*�7l�M78�Z0��{w��)Q�F�P&�)TI'PI�G��,n84�Y-2].̗��{��}���.˾M�Y������ �+F�Ʌ��Ԑc)�j��ds�5���V��Z0 i7���"d:�Q>���*Q9"�E`{vi`W�&T~�f��׺��۱P�ʎ49P�w7l�M�	�s�|����YNr�)�
73w�5��]�`��s܃�ps����B��1d�M�������N�W8�Vy-q��$�p;�"�764b�v^f�1�}�s�ռ��FK3Jݱ�����N��f��"�e��Qzv�y7*<���\NݯJuh��B[�rܬ[�ub�nv���w6�:jH�m�;P�Nc���ogn�{���s���9X);6�ݐY���S����Fyv띳ll󮅎ݚ�V�-�5���PO���S'��cp����6ѹl���d.ڑε�2�v��u�KcR�ڲ�|�9�꣓su57o@��_� �+F ��ZozP�=�RS��r&ƣqXnL/�2>�f �~� �� ��E�]��r]�Nـ}Ԟ��78�f�>FW�H�:�D�)�!a�{�Ѡy���Nف�K��`?L�y����I�)�;�7� �ץ��Ʌ��fozy�mCu�F�h��	�6������]nvv��6���f���2k��a�t��p�('$Q8�����x����݁�~�`}�f�Hr�Q'*.�����g>��%h.�� 	N	��v n���npD+�e�]�\\U�]\�	$�@J�9��� �<�`}�nĥ*�ECiTM���Ɯ��s�j��9�OtuE8�q��'"lj7X��U��y���fozc�V�*��EEH�A����h:r��e��Kɶ�O1�+��2�'#������ I"r宁���`g�7�1�q�����H�RrG"�R{�%I�Ss�j�� ߜ̆2���&䡹ށ��U���U���?+�Ú�ci1��.���آ)�TChj�:��F`���,L`�_j����'�](��Bt& LM���f�Df�Μ�6Z07f%��1��Ɲ� Y�	!�i6����p�/r�pѺ��EEqx�Ѭh��PB�.(���;|�i21�p��&*�	þ�M��2�sy�u��nw%���*!Ouu�h-ɬ��A&�b��Ӥ)�e"��6cZ��؂S�ׄ�"�)13�)��0o �P��3��k�Bh��ĩ��y��:Xe�f���ǁ���$��G�M�<�����*;0�@;4 ��SJH��6pM<<I�)�2�X�)��"`������$�FY�!i���$e� �+�$�  ���x7�׺���3=�ހ}�4ރ��T�'���s�����>t��	GW�C��#��nߧ �~��	ʍD��#�[�Q���`eg�{�3j�5nk�>�z5X!G����\]�#�]�K;n]���p=��#$J�"���t�Jp��BT��������������#d:��~���Ԓ*)A���@�{��չ���b�3=������H76��"jA9c����=>~��IN �W�@J�� ��t)ԩRD���o�{^�3=��uW��ﳕ�6}��.ccV��#`���`XNkF�L�&������A�H)��vfc.�d�olD�i�H&�V��
QUUB���^$���O��q��Yuw8WW�@J�� m;Á��`~��o�0�~M8����Sd�"m:#�F�٠@}��\�a�+6��rF�`�S$!I�(n}����`j��`}�+�r��w7�z������u99"����N��%8]Ot���Zuʂ�r�uK��=�uX�f��f=�`j��`g�%e9q�J��9W8�'�T��Ru�|�)�;ջ�D�b*&��zc�V��xʒ�|����r=�|�<r8?~�ݲB�UN�U��S8[���}�z�j���k��&����x��f�-�Wk��cr��X�������-Mk!���L��G �"�A��v�T/Vc����C�l��t���:u��n3�óh)r�'#�63�.Y]</f�ٔHi/%� �n�_d+D�x1� 띷Yn�ku�c=���{uۡݛFg��\F0̹9.�b����n'm&�ң�9AF~~~�۞[���Y����k;��ng���kO�[u���Q�WW+ٺ�qvX��f˹`~��Xʒ�|������՛C[��J�$D��|�׺��Ot):���?r&O�\'WU��
�Ȭ��~�@ś�����`}�1Xf��)�TP�ܔӝ��� �N��%8��$�@>d��a �T䈒; ����y���ٛށ�7]��c�@�t�QIکH��[y���<v�uݭ���=^��7�J�l��.��(�s/@�� ��=��� =����VJ�r*�(:t�8�=����]��3�5(|�;>^�.�[�Q�͖�����ؔR&��J�i�{�)M� .�^� o��$��Jq��p�iI)�{�,��,���@)M� ��
�.฻��沯+@�� #��[�Jn� ��}1%�E����!r�,whI��s�!��ccdԞ;`p�R8�T&�q�����g��^�7Dj$�R9�?���w�f=�`b���c�V�ԕ�f�B�rB9�T��
{�Xʒ����r9�/h�kBA���R+�{�*���{�r��� ;!1I�
��L�aR0S���#� `��*��z�i��r9��<�۠z=I� �i��U\E�D�Pl�V��M� �[݀�� S�c�3Ւ��!Pt��q�`n�w����9��Z��`*Jp����vsJ��sνu�g:�8���0�,�<�y��s�|��Z؝t6-�(�_��
Su�)�U`*Jp���H�N2:�44���^�;짘��n��b��`b�P�cڍ�N5J��ht�� �[�Jn� Sު�>F<�JQ���H�Vo�{�1f��_g�{�Wb$(@��!@v���^��s�u�ٙY��y���⪯t)������%8}o{@�mHJ�"l�B�)L�#T�����;��3ta�絺�R��(=����	뮎Jd|�Q�`j���V<�`f�w}Ȉ���z�w��6vr��M���:���{���`
{�X�)YN#���88��n��b��g�R^ך�
���`}��R��q������ I��>�]S�|�)��D��߾��k�R�dt'�)$�>Y�vʒ���� �w�>v\#�����,�ύ}�ŭoF����k\9.�U�����xA���]��NW95iӥ�\�$k(�hw6&1[;)k��\&e�5+����N�;nÖsu�HDWN���Սm��P�,\t�^;t��8^\�W\-����/9�vN�YT�=i�ƈ�=�������s�ǃZ;��{a��r�Y�:�m�8����nm�,u����v�[��.u��VN�kq9�w3Z9�4Y�f�Ex#�#-�-f��Ѽ���׌�L���z�]m�Ӆ�A���v�wK!�.��F���r�$I��o�}�����k��(M�����>��7w7d�d]���u�����]U�|�b�>�I7��B��Cs�n��]U�|�)��{��%ML8���"�.
���]U�|�)��{�	n�>��U)�q�R�U�v������ ��xҺ� Q�
Luw�nC�T�p�(e��gc���ޕ[�X�W�r�ʒ�ܢ��N㍎�8�+s��@r���]U�6C�����E�T���I�;�1f�+��W/����� `��S0ł��@ B��C���QC���ى/��+s۽�ecڕ##�844���>��Xʒ������`
TcK6	�N��ar[�e7��}����u�[����6�9R8Ĝ*�� ��=��� �� �RS�}��h�)(�2��n>$�H�n�WkGy�#qr�^;������DX,�-�k���Jn��N+ �RS�w���,MV�*FTe@�;�s]��<�`{���@ś���{6�Jr�Ԧ�w9�uW�kﳕy߾��Vd��@�H���v��}����G����g�%c�i��88�}����u�vZu��D��s�v�蹋������d��n��s]��<�`{���@�\��o�����DeE	)�c)&��<���]�}�)�[�ݹ�+���J���N���Ғ>����v�����3�z��,[Z�͂r��ar[�t��O�~� o޸�;):�>�Œ�F�C�H�l��f��f�<�5�c�V٥$��$���w�������K~��INǎs����Repq|�s0ĴQ,Z �>7���;����sX|�eFTB�K�3]��<�`wٛހfn�+ن�7"�ȔR1���5�zc��msd��;k�t��d��h��N���לܪ��Sj�]�}��U��foz��?Ur���:�7+el�mI)�QWW8�/n���������>O1XW�VѵT�Q��w�b�u�vRu�j�� ޤ�@�R�qW3u�HiG��W=����^�;����fl��ԖlNH�B��@��s�O����}r�=�~�'�Z�_������Y��E\��DPU��`�a��@T @�io\��;@FX@J*���@�`C7�"� �h%U��P?�` ��i!!�d� d��Up��U	�UX�P�@)Q !J`�A(@Y��`R � ��@:W���u�D5��Ҩ*Ъ
�G�{�_�?��;�l���D?�D?�TC�
�y�G�Ԩ����C�e@��!��"&*����D?���*���@�UUUUQUUUUUUUTUU�D?���������
b����_���w�������G���f��}t�*(�����������'��������TQU����?0��lO�����@�������������K�O����*(��������:�������|������Ƴ�gɰ��( �����oJ��4"�$�¢D(�
�1 �2�C
$$"���,����*$��
J� �
H) B�*J�(B)
R"A�H)* A �(�B�2�D��HD
�	�$��A!!		$,)! �H$�J�� H@$�+)!	)!$����������0BI!$�������	 �J����!"�	!"�� B���(BB �!*�# H,��@$��@�	*�@�$*HH�����!	!	 H2$� �B�!��,�"$���������!,���"��(2HB�(2� J������J,"�B���J,���(�B�J 2"	"� �@H�$���H 2�(J��B ���� $��
�B��B@����$ �"�!(���(��� �"H B!2�J# @�� 	 J��(B�@�!0�H�� ���!B
�! H��� 	Qa	�$RP�YQ$� @�B$	 ! $! 	D!!	D!A�$ ��RA�P�R�B$	@�e	Q� 	!d	�!�f�B@�BYP�Q%�$� �a� $Y�%aaB`�b@�F�&A�Bd�%�hBA��A���@����%!eA�Bd�hBHF�`a�$���bQ��Dh@�bh�
@ZA�H�h)D(�I@�	%�A`�	$R%A@3����?����Qi@�#������:���^�������/������ TUt�5�͞ѯ���?�����������濱�eQEW?��YUH>?��?���?�� ���1QEW���'��(**������LsH
����������������P �D� ��g��5�����k���aڨ����������E_��� �w?���l����UU������E_�z����7����������'���p�����s�Ͽ��q��x�(�쿲��Q�xNiПӣ�F�d���������{����E_���?Ԡ�#|;<�TQU�����g����C�6~��I���e5��`�J� �s2}p���*�
            D    T    �J��(	UP��@�H 	U*� E@  R�$R@}d P � �T�E�QIH �� u D�B�  ww �f}����������  �A�������M}����N�AQJ�}�Oz�@7x �<j��0i��� {�&��W&�e�rr�>��!|>�(T	P  � (|}�щ��"4�V6�#M:� zi���ݔ�6R�R#A@��ҝ6 =t ggG�t�4� )��` �`�'@�D�4�3� 1=:��  � HOL@��bPC�$�x�@B  P 9�FA�� �}|Zz��s5T���'n�rԣ�e� t�%2w�꼍xyzk8q=�B� �c:�_{u	��sW� r�/�k�Ϭ��%��W��� )	UI   wX �DŨ1����deW�P�(�oZ]�Fwp�i��w�+'ݔ�7�z 	�x�+>� ��ڨ�j,��3�� �Š�>�ϸ;���	J��x  "*R   f� y�Lo�d����/gTX }8������C�C��` ��Jd�d7�"3�6��}��.� 8	����{�7g!�� Gx�v���a�>����  OPT�ҕ*h  B��   <z�T@  Ob�Rl�� �T��%6�JT���C�
�ڥJS����)��5�/��DJ�������t��t����$�!_���
��U?�U��U�dV"�����?�)����XQ
L%Af/��p�XZՅ�Z�"��R��gdI��h��xS�2���}T��M2'
��Yc�|�d
dLk!)�"Pd��$D���e��:��@�e��165*��˴�%��{����2�]�UA�kb}��C�4�8�!�r���范U{(�kT�>a
,�Їq>5}�o��H�����R;d����W?;�(����.h=�iv&OC���6.+�Ǜ(�A�Rܱ���U	���ݷfY`�b��dŲ���Zr���O�A��/����y���dڝ�{\C6i{��RjQR^c����p�����>j#q�&J���٢�oj1`�6�x"�f*�/����cCQR�3�o��yZh�fi/�����ĒG<tͮ&�c�Hh���5�ч��y�Y�<9M����h}̿T��+`�M��C��)w��#¶�d���Wջ՜�C�pc(���]�ټa־*�^�g,�\�|]m}~ͳ���]y�G5
%����^��+�u�u��I�zQ���r�ʶ6��d�[Q���2�SN5I�GM�J�6�
���8jͰ�A�) � 0)�5�b���g�]�Q�m��,�(��=޺C0���6q�}��Qye�\�n:V�K�ɄTZ��؁���.�,�^8-D	�Z�8cH�V����{__��HYVmIUe�f�]�B�LS�U׋N2|{U����y�W�g���Q����C�e�^PȆ&�F�ӫ�l���}D1�װ�|^#�t�I��Y}��&v���߉��p��A�B&b��#^�m@�ZY�Qf�6ɶ�i��_!���q����:�v�{�_�	3��Ji�j?m
�=1��Z�L�`ʳ�f��ھ^(�����b5�l<�Ջ�i2�^��
�ɤD�q��4(��M:׆x"a ������e�VP1�G��B�6q��Ѵ>�=v�x��U~}��3��:k�V�6�v{�/���/��?�_�cP�g�Ӑ��{8h����bE��� 
�0���^v�n��WGG}_zv��+�ΔΣ��=���|ᆤ�1�U�����d}�q��znb���8R�%�՞��w6�P2|^�QӺ�������}O�*�NQu����@��)�����Wj&�T]ƻ7�=��B
��`�5 )�#�1�f�)�~��v'Tl��e�]i�!V?=�I!�Q�J�S���fd��d���/���u�U_K�n��w�g�ܫ,��p���j����Ǳ�EV}�z���T^j�w{׳��+��)2�m�;>��8v���������Wj�ecQXL�NZu��<�(ʽ�a{�8iW�V{g�u�<�U�w��}�p%Y�f��g��8Y��{7�z��VEJ�7Th��Ex���C��2��"QJ/�(������a
������h����o���<C�!Dw��x����G�<��h Z�����d=d�y�������;ު�8J!g���x��4�4��&�Te��^�d�n;yXm�]n����}���<��Ǵ�<�B���0L���l�:�́l�w�廞R��5'D��t^�ǰ߃�Iʼ&�w*Ԝ*�f�ͯ1�'�Ej� �OQ�2"�J0PV�V�	#�ib�U�1 �ģ$��A
(F&��Qd#�SN���R*�Hn@ ��HI,SC�$#�
�"X�!(����Z!�����H)�� PHB@��QbA #tD�#�,T�j�H�4Ȁ@H��$#�c@�V@�GK�B�$� (mH�	 0��H)�A��R,�QaM$lT��bX@`�R)0M1�� �5D� �" `�B+6� ���b@c]�7�O��%ը�qe�0�]�5r9���2��߆�dea������ŗ�15
Vav���UY0ӕ�jR�/N^�"�Ӭ��4�d(�,����e8P�6v�]�!5W��}=��sw�/�ɱ��Dʳ
���i�Ī��˸����c%U���P�Q�=�K�0M�8R�EDB�2�ѣȉ�A���#���iū��hjU�w�J��62W��M*1²�,�z��W=6�������1�7�e��74u�+s7���Ϸ�g䚃�Ͳ·-߷<	�/Eq�Σɦ9^���yn�"�ۧ{=<�3�n15�F]ǹ�ϸX5F�݅ߵ�˺>�8��(�񼆚e^i���CLt��V��o�^vN�4��E�o�\�{��K�Qg�hp���7/�����\��uNW��u�셝^�	WY����5*��a�k�����D*�5ﰕ��E�2W�g�f��_d��@d*�ټl��˙�2S,�s*V���$9קqx�e�ی�ɚ[������D!Ax+I�e�m?��2�U�w�^ Ƙ@�/6��ӏ����ihZ3�Y�>�����-Si��Ԣ�Ǘ�xL��T��^�~�� d*�̔V�����W�e�:yS��l_��m7�����u}{�m�3���c���B��"�.;���!_e�gC�����]]��z�<*�c|3��˖�I2Q�64�D���WC�[�8�ןS�$]d[�^�8U�Y��J��+�'�˓���'ǹ+�*��7���︂dP�1-/��J����Qg��M���N�g�!�Y����j�j�A��Wj.ܳL>�6��|J=��qvB�˷��V2��{s'��n�m�82�Jwن���J�5�oz���[`2*-��(�&��,��a�f��u"*H�ql���y11��*�yg���WzK���!=e��զ �W�4}�Şg(���G�����,/�QپҨ����&S�-ey^�ME��iG��wk�x"uyT�]�5S`���hW�}�H���u�ڿ�`�U�,�ٸw�-i���Y����h6ҫ�N5Q���
!Y��{��6h԰&X�,4�2RtX�ӳq�C��4�@ �%��F� �&D�J��1�ن���2r�!�6�`�ZN�r��7mGD�'T5LL�5�r�,d���U�+�];8K� �b�B�!�Di��@�GK�!"mB��t�5��CXU�D��F,�}O�w�j�T�a
mf��g��}���)�x�=ٺI�_3׶�r��nt��$�/	�O��ګCzaEU>�&i9X��2��ez�&�<�Qi�Ȳ�v��rF�T�%���N��;ݯ.f��[����ݞ7�g��xAlPCP����}yHq������ �g+@Ȓ`4�-bM�d*̻==�}|P)�-	��xN
�O���}uq��ɒ�������J�6�aW�t�}i��1�Ý\��Q�U��5214Zhi��2�^2�mb4	�۳��5��"[�[�ccwTZ�d��0���
36hˢo��˶�5�`5
e����4�Ęڅa����6�0d)]��LyUF+@�6�at:צC jQk/%l�>U�2�!/-�teë꛹k�d)i��]I\��`Ԣˆ=/$����9E�N�H^�L�idǷ�Uim���x]I�W��m�μ}�Y'���o<n߯��Xcc\+��a���si8Q�mb�n�(���fq��MCcQ����Ӎz�'y�]S���%@�%m���~}�9E�a�,���MB�Uޏ��*�i�~~!�MEQ��}5a��JE^l�J+��rC�vg�Ϲcm��i�,�3Ȉa"e+ʡ�j���9QG�cC�喬���Z�m��˷�Kʳc��T��ZjU��Q���ɞ�R(j*Yۺ�Va�3޿}��<�	���o�6i���jz�%v�t��vx�(�.���qt�C�v����U����W�Q��9��Λ��0s�����_���
-e��|g�q��jZ0LD)8���&2U�5^���*�l�s�r�����?�B��>��8Uc+OW���]Ģ�-4�p��"B
B0�܉������]Q�Z�#D�}
��ЗR����9~��+����Գְ#Ml�t���M��)�@DcH��6�8%_�i���2��a��w,�Hd)w?vb�j��K��ګ��R��T����f��d�NU��8�0�>�t8U՘�ny���O��ڠ�	W���3��ni�W�j�ôҋ��A��T�L�Q5Y+�=��g�~I��/;t��C%Xi�퇳g�Q>��2_���0��v��2#�͟w+,��ơW����N�4J;��x���tY�6�+4�*�Я��r|@d#+=\��m�CEe�Z�<pZ^p�̲��1Q�٠8R���L!W�5T���V�X�1ӕL��4��od�7겪���r��7^��x�+<GVZ>U�ː�}�_��U�dl��˴ܢ���6��O3�<������|2������Ǿ=y��w÷;Z�eJ{y홝�d(�[;�|qX�Q-����4��Uy��o�I�y�7ue/u�������=W>���ww`  m�  $            �    ���  �      ��              @ �                               ?�>  �   	       � �    �ͤٶ�me��#2��j�k8�<�+UҀ��wQ�j�b�j��{<Լ��V�l���H�eQ٦�<�du���U�VuE��X�m�mN�8	ݱ��$���h9���	�5O!ڹ��_f�Yf���$�+	9�f�����n�U�Z�d2��=9��ny8�K����%<���ZkΒSZÎ�g[d�7i6k��[��Kg��Jյ@S�ˮ�ӧnH �[��m��nѷlm�vgK������[R �9��*�Ur�c3�6�%�ʙR��n��l	6^;#�:���N��ʣ�W���k��ԫq�'q�����K,�Sz�$�iT���'f��\��iJf� ���J�48���2�)�ܠK+[���;tJ4v�k��;K��[��t��\5�c����N�nݎ�j��X�v��{��[�*�1��f�� ������:K&�Nu��NN�u\[m�;t���F�j��X -��[Y$5�'��u�b��ک.I��\QM���&����jz�Y2���uç��Lq�\%$ ��j�wI�H�
qR&�d��vh��ƃ|r(���\���j�z��an*�W�uUJkJl��Czp�wl��s�vs7!5p�l�m��Dq���pۣ'��;�G\�u�m��lUu�=�8�,����RU*�S�/CM�n]hlp���Uz�؇{ed5�6��@
�4'Om�c�0؞d޹�kl   H @(۳R�sZ�;MuH��ݓ0�[% �a���s,�۞]�[j�����)�8-�� ���m+��^#m�L�2P	 m��Hv��tQ�Ɖ��� 8��\I�U[F� !I�l5 Z]���� I���[@�� 8�m�H�4�k%���m�amN�� r鴁�[v��{fG-� lF��]@mKRrH]&��Qn ��l��W/P}6�}7k��E��H ���:��� ������A�ݵ�7$'$n^��m��N�n�8H��@m�D9�^�)]���`� WF��m�su�H�U����
�F�۴�)ջ25��H�8  ����6��K�he@ق�UU*�m�۲�����3m��`M��<�wm��㋧<�R���UV�u��i�;e�V��[�;�؀%�k�Z�!��;M�b��k[b��:�	
�UX6��R�s*�[0,K�0�q�j(�U�)kE5�V$0H6ٴ���&�   u���q��씽QpS���qut�Խ]�Yٕ�t!;�*�ʴ�UTU�L����Խ+G*Ѯ@6lGKe*��*h3���*��k Hk56�G[M�lsi9��*Z۶�sm� �RFۜ �f�L�/K�n��Hn�*�Y�l���� 6� I�����p m��� �  8�  �m�   � v�$����=�ƻO
�qҭ�UWJ���Vʙ�x��׶�%���}�o�l��*����j�VyPGAf�]$�,��9�	���L�����V�;)JPM���&���y��c� 6�l�)d��HM��YY@%��{]e�햀pUJ�u�e8v��{q��]��l       @       kX � ���   md�     pͶ �l�` � �   �A�`�6��F�    ���    �� ְ�   �l    -� m�q��m� А$|q�� m�� 8 h� �ͺ���em�ʵ:7J�{X�UWVհ�Wn.w7E�vB���TZm�Hl8� ں� *��3�H/>^����\۴���N��z�/[V���x[@t�m�l$�n��#Ysm�ձ���#�֒d�h l i�H����mb馔H -�    	 8 i"A�`�cm� �m lm�m �`l ��Ha�h�� i66� $�  �kh8   $� �   �m�    I�@ �R@�     	 �P �   �   � 6�5�l�	 l[@m  ��   �`  	�m    �R�l  6�[@   6�@	  ��6�    �  �   ۲�mh8ەV���&yJ��5&s��k��^�A5K�[�����  UJn�q�e���qmJKUs�N�t;7m�ٺ�ѽ���g��sJ�M�A棒���ve��\��)[��Zb[e��R�l �6�|�   �m    �7m�   	�m�  ����ְ�P-�  �[A�À| ��   ��m�kh   E��  �� ��m�  -��$ qoQ$8��݉|-���[jv�v�91��<�ׁ��RZ��YV����mڥie�&�g�n�m   �*��VriB�8�
|����Z&���`�[��/�-E�q�	�U��� � ��UT�/-]Q���VP��V9�{l����j��6�������5\�e\;O���n�Y���s�9�bu�2�+��d��]�	�Z��O����n\5S�;`+-UWf�sOL�+o[J�R��ͤY�݋�mVǘ�n�6������ˇ<z���5���v��p�M�M nxq��b�Gx�a�5��1� *��m1/+$��ga�M��hzn��K:&���|�o�4l��@ �6�I��%��m���UU�m�s�:۞hK �[]-T�j�r7,]���=c��C��\�j���v:�^c���ݭ+x�j-�%Z�݌]���ԮɅ;4͞�T��k��!,���>sǍ���'����rܜ�%s䗪�v�6��(��R��qy��&[���:��d�P�U��U��5���wN�9�wHɳ<����ق۶
�S��ke[�^���T��\��/kH�-���F+��^v-���1�d��ԗ#�3����s<PQr�<wn�;8wv�A�T��n{�Z;q$���u��Tn���d�m���e������*��9��8�ݹ�MvBm/<�fg�Ƒ�5�tC�qC[LVʷ.	�-.�r�5�mQ]���ˎ˼�M�<Fɰ�	+��ct!f9��Y��2,SlLJ�P^2�D����I��n���pjiL��v��:��[��8��m��y�;�����W�/#��d�q$���P�n���`�F���1ůI�l,�UUn��@�*C�l�l��UekP��utWA�t�Ӷ��v��#^ݭ��gK�Y��l�: m�Nuzp-���(d0k\�����Ƅ��n��gi��u�,e@Uv�(�"�`��h�2v�0�����m�^��"͗g�Su<�J�W��TmPW����m�v�M'`M��&�t��ʖ@j��ѧ�g@U ��2nͱ)���c�n����1�0l철-o���rMRkJ�+yD��Ӧݶ���:C���Ӎ+m��%�Uu*��8ݳV�kX�q��:y��](���� 8)�8@����6>;+��B����d���R�=r2�ӕ@Z5��v� q���i��*B�>�F�K/ӳl;~bO��vHz
���e^�z�۴q������Ɯ�/�Tj���W,��̨d�^y���@vӺ%tm�5N뫇�o��@�si��d�lp��gm�^��q���
=B�-�U@WUUY푮�l`)UÞ&�(��몠.�	Iy�i�۶�;�V1�)��4�kX/M�4�$ HH 6��4�[���h8�	Ӧ�X9:���U4q�6�G��Bkk��f���VچN<������_�'E��
)�e��ʶ���U	5a��#�Ug�j�;��YI�=I�:Um!��l�e�yR³E-��6M�5\�'�]�@n�W$@�p���\�����\v�ԸL��78��f��鴝b��˽:ud^갶�������h"9��.���][���ΐ��k2΋[-�mnN��k7\�`���V�ĵm����s��9H���'lL���v��[����!���-x歮˨�8�F�=�ɹ���E�Z���8��vC�;�sΖ��@HM�]>ք��Yd���OJ������ٗYj�����s�KL���Ȯ˱���L5�cg�m��|�b$������^F�ڦ�p�.j�⫳��-U��8�p�x%�%HG��Z�'F��h'n����.ʹ@�+��Z'�������9�x�E���:�`]���^�vtF�qu '��ҦXIV��:m�7�Z�������ά����3��<��6⧖��I�S��g`,v�wh�F�8 �.�9��(�"�QW��Q?�(�?��AO�Q x�h(D�zH�$�"��Tv��Q��T?�'�? �pW�"���#(�N���]��I��y?������X�U���UN�ʿ(��x�xQ�KP�
Z�r@j\ >D֑��UG���z�/��d���O� t�n*P�A~Sb��&�@<=S�A>^��P@�ES�a�H�6#�P^�|/DD6�i�
hV ���� �|�/���D��8�� AW����+_�EM�'�u�='�� �`�1HB�a$"F?�x*�B
/�������)Q�$0#uV�+��ȀO�����t'�&��4 �QEҾ������J�<D8/��H *��@،A�`@)"���R*�P"� +*�h�P�D*����# ��������m-� ��H�   D�     �q!��kh�W��TQ��93vi���V��s��g#�[��Bv5��Ah���Ή2�mr�T����6�wZɝ����Y�Ӱ��e�)��a�'i��7�b�4݂ӝ�֌�Ck�X�17CzB�s��'+�N�^i���=x��9�H�n@�{�[R��7J���k���m�]��m��
UZ�j�Z�[��&ʨ�:�;K�,�e��e䞃W���ù�TecoXiP�@�&��7�X*;A;m��M�u�!vݛ[c�����v�M۷	�9:v|'o9�]��ӧ���^׉3JK�$֠��U(u��Z��ru�N�tu�{���xR2��T�:�{c:��iP���` �dQ6���]�lH[Cm���J�PY�h��i	U6��DU؎Qm3pn)˃�nr��f�ge�ϕ��RH�6j�"U�R��m�8mZۉnC,-���[VԀ6��Ѷ�pK�]5UJ�U�G
�s���
A����6֨ێs�ܐ��k$��-UmUN��.n(��V�յ��$�bU�n�e�l��Gh�HTi��Om</��Pږ���nK����`���]�$9G�N�ZyՌt���@���/���n+�^"8ӥ��۵���ѥ�۱�v��;n��V�}����;!��'���v%�m듵���{WΘ�c��ؼrW���6ݐх��K�
՗5ϵ�y�m�Y�:^8Ѻ
�AL��W.6�����O"�yn����p�9ENv��m�0W����y��<�]��8�ۧ�l�]�;�xǝ�< �.s�v��u\�r��(�rm�)���W1K�.V����ۅu��ܹ�6<v��d�s�D[v��8�nq���\8�Y�;@�3��s���c�S��<�G���wl��.�%�K<9�O8�eힺ��c@�]=�u��i�irZ�5v\��UIc�BIp%~I(x��QҨ.������W��w~�����>�t��P�,F��:��x�2v&|�[w:V�$��/�z�7Zw'\=��d�Ǘ�a9�\N-�r\��a�S�݉��ml!l4E�-�ge�`4��UV�f 6�<m�lu�c&���K��q�#�St�����{�%�{=]�5K�u�ᎋI��p�=�݃] n݄�']�w�5��w]�$�b1iw�Ջ<d#bꋱ�������rF�vS;��"���v\�vs�^1�����cre��������ZX�^�ޢ"?H{_fhK?D��`�G&8��@�t��֩M�s@/[4���Xӆq�(�u�S@�۹�������\����H�67p�>��h�@�빡ȼ�4�J	�A'I�{��;��hz:�ͼX(j���⮤S4U���S�:3��s�&���ㆳ��F�9��OW='��R57�&��z���;�:��]� ��4u0����x�`�q�~﮾�aǅɠ�m;J,�V!6��!	�@�H�P�ZJ#��� ~m��o ~Z����4��D�=ץ4]k����(Q2��,����=�������J��FD�r�^�ץ4�]z^��=N�6Ŏa&)"29�׮�غ�4�)�r�^���߾#p��]����o��Ĳ��#`秶�y�pkqE.�ŕ{n����G]6&�ͷ��~��^��<���:����\R��G#x�ؔ�@�Қ�uz^��9y[4��.	�C!�n�u��m�~�!D-������k�f����J�H��"Fԏ@�Қ/+f�ץ4.��u0ʅ��x�	��r�hzS@��^�ץ4uBGX�x�'1�6���%�ojsB�֫�tUs�ԒgY|�4�9۷4�#$�����94^��.���S@�ˬ�={��9����Ĝz˭z�Jh�u�^����6�'2&Dcr=��4\��?b_�����~zg\���d��Q�@���x��8���ː���

�J����o��O��s��z�D�?���/>�@�^�@�����w�tm��渫U4J��
����өN���u�ۜ������^���]���ps���O� ���<�_�@���#�g�~��Z�W���I �$jG�[Қ#�f���^��^���If�q�����@�{��9{��>W��>VנpV< F��A94��h+k�>Vנr;��:�WV]TUE�.j�p�۬�G����F����8$�/`�BQ%)%�5cͷ`0" �-Pm������X��Q�j�5E�qݿ�}��dڡ�UU��jM����:�[���Vݵݾ+m5��y
�r`�����\[���gV�.��9�!ݸN�rnN�c���qF�8�BͶm�;t������|?�a��)�졳:ݫ�}Ȣ�FЗ;����cOn\u���á���G��Q�'jv7XX�H�����o=�=E�c�)���#�M�6�G:� ��χ�z֭��rf���i�B�g��k"�i�f܎�l��^.^�����I�9�T��궨ܴ|_�~z#����Z������Y����$�#���g��$V���Հ���?y�YE���.���rh��>]k���@�;��;��\�"O��C@�u�O$u��RIy��}�Iu���$��A���F�|�G[�5$���g�$�Y*Z�K�ֿ�I%�S4�7����#�v�G��<�[V�S�i���U���
�V�[���.�8�`�� �g�$�Y*Z�K�ֿٟٞ�I��ɩ ~~v�N9?gH/������_������B��`3J/Ȕ9�%ߟ�$���MI%�wY��%�qk׍4&d�H�kRI|����%��ǩ$���>�$��ZԒV�lm��d�$���|����ο߾ǩ$�-�>�$��ZԒ_;k�䒹n�� �y$�o{5�m�j}����n ��s5{m��Y���$�[��$�S;�G�1�����9�h{ܽ��:��s��y�h�&�t���L�z�3�� _��> ??���K���RI^���K��P�Jc���9�I���-_}�3����?RI~�����I.�ũ$��p#.9F?�wr���z}:�$�O���e�K�����vlZ�K�-_|�\�ʑ��H�1$��Ԓ^gu�|�K��jI/����$��E�$�݅k�9�%�PNO�I%�X�$���|�]\�Ԓ]��������ѯˬp���:�����z��bU�)��ݍ�n�R�Ӗ�k�G�e&d�5$�RI|�W��%k�Z�K�����V�����f6�i9�ۏ�J�(����cm+�����$�?ߣԒ_;�������ڹ���� 䐑�������|�J�cԒ_;���IZ�����W�FӘ��G�q��RO�﮲I&����d����$��1%�"��(@H��F% �`AiQ"H� ���=����%ϱG��a�$�s�=I%�_�$��T�$�c�W��$��=@����9��ls���[t;z;.ˬrP�m��3��x��vn�5%���s�RH�|�V�R�$�=:��I![\Ԓ_;���IU�T��G�$�⼶�����{�ֵm�������w��l��I%�e[�c�sJ<��_|�I[dԒ_;���%k��RIvzu_|�K���7bd���Ԓ_;���IUn�Ԓ]��W�$���h�V�]q�9��6��䒮�f�����c�Ͼ��$�m}�vI�!�Uv����1z�f٥đ���Xps6^�%ӚfC�=E� �Lۥ�l��h�W�#e�	º�6�y���[������8���k�T�u؎Mzl��L��d���zvر�m��q��� ͬ
J$��AoZ:�n6M���z��/�`�㿯�t�4N�,Z�:y��t�(c�g�S��v*�m'��8x���#.��=�o1��{-����0���������n���n:z��WU6f!��q�
�E�&�\����*��oM�:1oGGY,ra�&�O$���~�/�I![\Ԓ_;���I�ɩ$����$Mc�y$�����I%�_�$���MI%���}�Iyv(�!�H�1�NG5$���|�G[�5$�g�U��$.��I%_*ˎDя�I"���In�Ԓ]��W�$���5$���|�Ug#58�D���L��K�Ӫ���������s�^����${��Ԓ^� [ ��'&��w]p��j�,;��l�c���WeK�����ۮ	�.`����������� �z��I#�w&������$�;q�7*��S�uR�$�m}�vƆ�c`�!�B#��/�9�9��&������I!{���K�`��C�M���${���$����$��Y5$�Ϻ��I.�p�X��D�G$5$�z.��I/usRI|����=�rjI/z��E�LM9�o#m���$��jI/��|�G�RjI/wj��?{��~_�ev�ϫD�:�`6�.��n��NS��h��-դ�����󇗅��S�	�'#�$���ߟ�$��K�9W��$/usRIy�Aq�'����K�ݒG޿���@*���_��n�#���Ԓ_?Z���m~y$	ǉE��*�d�O}Oջ�w���9>Lg���II�T�� X�ԺHH�#R51�X��P�h�w�f�/�R�2�'�W�
���Z�J�pҵ��k���i��4���,��N	FRV�C &��j'��T�����=c�{{�qP"�ݱ�0d�dM@V,YRU��5�$�F�Pe�P�BD�"�6Ӊ�4Af��D� �ĔXU�HЋaR%IXQ�aVTeYVQe#D�7�]M���J���\uHu�Xm �!���jP�EB�)JN��U��"�鲒,���	�� �h¤�+@�B5c@� VT�IXT�I�:�4E7��;E�TA��CZ�
�FC��c�DT�+��5���K0�)
���*� ��@�H]�eu��ě�T�(�5��y���K-8�eU�Q{��YF����D41�VЅaA0�x���Ĝ����r�Z7��!�(�O���П������P���/P��ASኣ��kｮ�Ԏ���m�럵�~�F%P�(�~��'_U�������ީ�5��3�D(������_�� �y\���oBS| �~���I�I�$�ӕ|�B�jH?}���m�G��7����خ���ཹ2���)[ظ���l�j:�7*ZYq�pVە�G"bN?y$��?RIwNU��I%�d�$�w��䒹n�-rdA�jI.�ʿ�I!wW5$���|�G��~G߾���T??���� �k��"G��$+9�I|�W��$z�MI%�9W��${,u�ba!c��I�$�{�ݒG;��I'�~�V�֥���?ШH0$�$��Ĉ��v}�w�I:��d�:�t��wwV��$�z��$��Ӫ��J��RI|��� �����P����.Й��h�(���Il
v^m�nkN�[ ���J�"CR6��%#��K�r��I+�MI%�_�$�W���K�e��Y#p�2
5�$�W���K�z��I![\Ԓ]����$�}q�m��B���$Ԓ_;k����I%���I+l��K�"K�$<NFĜ|�I[dԒ\�:��I![\Ԓ_;k��V�5���)&)��MI%���HV�W�I6���ݒI=��y$����@�4�V`#�0! "!#�B(A�E�D"0c ��a Hb1�N���y}���I �P��͸"2����n�\;�0�����܋��zsys��&�$�[<�<\6���+ʖ;v��WXu��sRmk�x���@d�ivCȯm����n2��5�n�X���g�$u��N��R�pS�&����3�]ON�q%�-����.��pWi��A�F�&��w�o���h��d�U.4�: �u�FY�3D轛�G[�+���!y$��3u�)�%�m�T�1ۊ2��d��\�At�t7\�=%GK�mэ��X�IάdJ@ALx���I�~sRI|�k��\�SRI/g�ϾI%s��D��LY&)#��K��_�$��lz�I{=�}�I�sRIW�.Q��I����G�$���5$��{���Z椒�����%˪@'��x��ɉ�椒^�u�|�B�\Ԓ_?Z��$�v��$��]O�R(���''�$���5$��ֿ�I#��@=��4B�GqK&q7l���I���1=������Z^�)i��Ö�2� j���o��~~?`��� <�����~���
��J�I9#q�V׳��bg�� ����|�g(�;��2��L�uVU�N= ���hu�@�zנz�V�޿єM�H#ɏ�@;���ֽ�ڴ��@.z��"x8L$�@�zנz�V��{�������rtq�o! 4�L��&;�(b&��'��k�Ä���f�7[��Y�5^_��#�@�mz��@:�4��z/r@&Tdhcq�G�� ��h/Z�]k�>�R6V�&�͓Wx������L	8��Iz"��/���6Mn�mkURӊ'��i�&����@�ֽ��Y��4Lu�pNG ��@r۬�!-�__�}׀~�7X�����-�9˱]pr\$;v*<����f$�L��cf�E��7�ݒ½��Hq E&�H��<�u�z٠}�)�U�^�޿��&�NAdy)&�_[4�e4
���<�u�s��Lr,N�hz�hwW�y�4�٠^k.T�7���9��*�@���x ���~Qu	b������E�l��4ю1��#�f�_[4�JhwW�~�_�@���x��yN��9�ָ�9�Y͙�<��&�\�h�:�A9�t�e��OHW��_Ͷ�����l}�)�U�^��{��>��Mɑ0����@����W����@/���H���r9�4
������L��� �w��Ʋ�f	�'�8�x}V�_u��Қ}�h���$����dhR- ~�xD(�y��s��7�k�����>�MC���QuNY;\��v�Iv�`3A6�:�"�La�:띇��͚�î�3[�����n��m��6k<v�[��x;v�چ�c�t��mKi��In�{*lp��V�dmZ��\4��i/.�P�	��3��>�LDtmD��{�wg&:�jFۏG�<��ܸ3�|�:"<C�3X��H���d�bk��Nݪ����W��L��l8��{޽�}�����7"�4�ջn����[�Z�Y��[���[m��Zf���<�I�:Rt���C�w� ~���7�k���@�����˦�j��TM]�v`�k��%�DU�� 5�׀~��9��G:�D�qR��f��]]� ��Ӏ����3�O�@=���>��k"�Nc�-Дϵ���}8����K[o� ��ckys��hW�h��4s�4�u�쨖C���	�&���kP�N6J9ս��}6��;��;'8�a C#Ț�A7�}�@�:S@>�@��z���%���yt��j����2��/�PH�I,.�R�@-�bib@�P��@B�Z�"�b�0�E4��������ֽ ������)#&'YsJ�� �k�ϛ�>J"d�>����αǑ�"�hzנ[f�{:S@;����v:��jj�SWwUu��w�rIB�j�O�o�U�^�}�<X�n�0�{hv���]��2Ȣ�V��!Wڸ&R�qu�YpHC�Y1�mɠ^gW��f�W�z��h{��8��N3e�`��J�ӽՀ�׀=���=]���$I �b�M�Z����%�_US��`7׀n��kɲ䫫�f��9$�{�^·Հ��
z����rʙ�uS74��ݕWx�5���ϯ�;�X+���\X�Ocx����Nr�`�f�K��ByOgG��H~���~��"m$DF�D���
�_�@�ֽe뮈_�9�����]E]+���UsvM�`�w�#���� �n���v5pm�7�N8ܚWj�Ѯ��2绫 ;{� �ֲff�f�Ț1A)�y�^�����٤���T�ݦ�hR��?
/����w��Oc��I'�'�J=�����@�e4����-�%$?�"��M�S��\��WhUQ��I\�� ��Ι��������p��5�s�Ⱦ �߿M��s@�ί@���@�0苏 �FG"Iɠ{��h���s�h��@�qs^$)���<�s4����ڴ�٠{��h��,I�0����WX�� ��ۯ�"'����pw��q�,n(�qh��@��ŀ=�]`�[�B�Y��ؒ �Y�eP�$%	H@'xo��_o�~�5�tO�5��+B�4h���@�$�JB�p�wLL��TLi1�.QC�"�����F�T P�H�6ڈ�D�F 5-�U≅[�0�(4M@��j��Iוn�f1��RV1�	H�������l� n� ��%cGuö��A1����8�Ͼ�S/6�T9I�NS(���ƚcLl#0c,&�a M$K*B
���#���(E(�a�LIU�O�O��C�΄bDC��Hwjl���r�H�c����9�9Vch��2#0# wa�a�ʒ����� �{7�i,D"�XI/H27P�!4�(��V��e"@�֊%x)�zK�&��c����>�am-��t H p  ��      !a�m��@گ1�uxs��e�=N: fj`"Te��b&���I1��k���/��W�:֍ܽm���.�t�������wWAu��s�^�s��\��[m˸U��m�l]��Ռ��^q^Px�ݝ���<�K��l�㎚���v����c�Q�����~�6�n��q���f��9 a�Kx��ȬdZ��C��f�ݝ���WŎ4]��Wb��ۧnV��<on59䳞Z*D�\q&��`z��N�A�x��c�gn6n�el'N��ȱ�ZN�:,[��f6��S��n�������H8�vU�x��k��=�i�����vv
<�h�٘v򜽦���Ojl	V���ԁT�*�Xpٯ����m�m�q��� �!5Jh��>j`�8�9��Y��������6� =�2�m]�d�^Z�Bɢ��
�A�
�eZ��D�K�E�mJ�Ԫj�U��n�Hl[���c�m����1���5�+������XֻX�ˇ6��` ��.��t%Y�P�`*ڵ
Ί�N��{&1.�*4�Xwq�s���
G�9��=�̛�.��]�mqV�뷳��۬���rZ]m�E�n^�۝�yخ��]�vl�Rn:m�sv�z7q�ݦY\�*M�v���m�v�pshչ7yq��ۭۢ�����Ƿ�V{5��x����s]��:`}"Ju�6��k����s�L!$slǘ�!ŝ��ї��X::�w@k94�n-�E�(zm�kWQ���@q���˅��؍*�[k��ܙ������cc��@Yy��$m驶7����eѫ���U��V7����R�T���,��Ϗ�Nj�%��]�[����r��u�.n�sE����v}:�����*�[���b�.n8���[=�\�J-v�����ݵ�[C��gb�����:離�#����X��������Tx�  ڴ@�g�>�?+w��}4Md� �m�F��H��Ԁlvn���ùy��n�ݐ�[��՘��v{'!���d�Xܦޕ�Ѷ]��g���Gku(��\��eY�m;z�<l��v�.G+�vvd��(:����;%���� �=�Q���}��|�s�;�[���z�]<���ܦ�� N�ˇÒ ��6y1۞��ٶ�U�䜧I�[�r���n�&u�ȈF5{8����{�Y�l���;B�����:��͎A�,U�l�bu��욑܆n�8z�+`s�k��4����Z��٠}�h�C�)�4�B93@�ί@�zנ���빠}��G�2O��'�!	��|�`�w��(�
gu�,������{��7��������f�����bX�%�s=��v%�bX�}����Kı37=��v%�bX���3\���$)!I	��h��Z������'bX�%������,K����k�ؖ%�bk�f���bX�%�ٛ�v%�bX���E��
oF���jl;\�t��9����ō�G6�Y�x�cU�N���\ҽQ�����7���{���q;ı,O�}���,K��g�\�蚉bX�{?t�v%�b#G�ːwn]T.:*���4�?���\N¨m@5�5��g�\Nı,K｝8��bX�&k�Ր��JB����Wʪ����u��w[��,K����׉ؖ%�b}�ΜNılK5���'bX�%�~�f���bX�'��=�r˫�n��u��o[�Nı,�����Kı3Y��v%�bX�����,K�Q?g3��v%�bX��~��\VzkO2��{���oq���~���5��Kİ[��7��Kı3��^'bX�%���:q;ı,O�ko������5Ӣ�tÖ!��]���"�g�mȀ6y�va_[v������Vb�x{��޸��bX�%�ٛ�v%�bX���^'bX�%���:p?(��&�X�'����\Nı,Kٿߥ��j��SWd�wwy�
HRB�7�d.�Vı,O�����Kı37��v%�bX�����?D�T���'�%]ЋWwtTՙ�
HR%������,K��߮k�ؖ5�D��dMD�fw|Nı,K=�d�v%�bX��wEޮ����F�����;ĳ�Q?~�_��v%�bX�߿~��,K��{�8��bX�'����BE>��n]���U+����P�B^m�, P��"X�%��fw�ؖ%�b{7�f���oq��������W�n���'��ݱ��3p��p�Q<gh����*�mɧx�/�]��MU�U�&�mwy�
HRB�7�8��bX�'���'bX�%��ߵ��v%�bX�����,K�����r�ݚ��޷w.�8��bX�'���'bX�%��}s7��Kı/ٙ�'bX�%���̜Nı,K>��J|L��-}��oq������O���;ı,K�fo�ؖ%�b}�s'�,K���;��Kı?��ww[٩4[�f�w��;ı,K�fo�ؖ%�b}�s'�,K���;��K�聄FDdA�B@�: ���Lׯ3|Nı,K߯��˶˄�����F�F��"}�s'�,K���~�x��,K��n���'bX�%�~���;Ļ�ow���~�����WWE�b�Tt+�Ş˅cn�u������e�K�gpf�2cn�HŽCvo{ަ��8��bX�'�����Kı=��f���bX�%�37��Kı>����ؖ%�bg�a�z�Wv�;��ws��4F��s���k?(��MD�/߿~��,K��g?N'bX�%��o2�;ı,O����GECizAg�w�{��7��������v%�bX�����ؖ%�b{�̼Nı,K�o5��v%�bX���\���*ՓW6������$)!I	�s'�,K����x��bX�'��k5��Kı/ٙ�'bX�%�����M�޵��no[�Nı,K��e�v%�bX��y���,KĿff���bX�'��e�v%�bX��������w��~$���$�˩*�9tu���@zv��YK�z�K�kA���:�����Г��/���G.w�8o=lh�����ݻL����l9�6���C�;7[��6;Z�Z1�m���aĠF76��9lg6�a$��3l�pN��A��'�Z��z��T����u�cv��5�;3�p��1h�������M{L�:�O��W ��[�i9c\_����|�j��p���˪5(̈x�Y'#�h��7/]�F�3�yڇ�3��Z�٭�W[�Nı,K������'bX�%�~���;ı,O{~���g�MD�,Of�~�Nı,K�3���We7D���uu�ֈ�#D�߿^#a�:���&f���v%�bX����x��bX�'��k5��Kı>����$[��X�U�������ow���Nı,K�ff���bX�'��k5��Kı/���'bX�%��3县7ut˕.�r��#Dh�ff���bX�'��k5��Kı/���'bX�%��}���,K�������ċVMM}��oq������y���,Kľ�f���bX�'��f���bX�%�37��Kıxt���Yʛ���D���U`��m�'%��tR�7g�v��ѳ�9$�{T�����kz�D�,K�~��'bX�%��}���,KĿff���bX�&��ud/�)!I
HN���f��]Ю������4F���~�F��$#�{�,K����v%�bX����\Nı,K�37��O�T�K������U�]ԕeʻ�F�F��.g���v%�bX��o5��v%�bX�����,K������,K�w������u���S�������D��w3\Nı,K����v%�bX�k��q;İ?$�L�~��'bX��4}���*mU]�(�����b5�4X�%�37��Kı>�ٚ�v%�bX�׳5��Kı?�����,x��{���~����;�#c�=�\[2H�A�ͯnsl����u��Vl��0#v�N�uݸ任�kDh����߫�%�b{^���,K����3|Nı,K����v%�bX��x9���WL�Wv;��F�F��>��~�F�X�%����f���bX�%�37��Kı>�ٚ�v%�bX�{&�wR���uw*��b5�4F�������6%�bX�=��'bX����M��_fk�ؖ%�bf��k�ؖ%������}�Yk�Ӂ�����7��,K����,K��_fk�ؖ%�bf���'bX�嚉��~��,��ow�?ݦ�t��Z�����%�b}��5��Kı3�̼Nı,K�_\��;ı,K����.��ow�;���?��8w[)�[�㋓OcIsC�ܖn:z�^6�on�%u�����#m]M�ޭ���oz�v%�bX���^'bX�%����f���bX�%�fo�ؖ%�b}��5��Kı>�zS5�K��wv][�w1�#Dh������bX�%��7��Kı>�ٚ�v%�bX�f�/�lK����um�7�MYt�ޮ��'bX�%�}���;ı,O��f���b�%��o2�;ı,O�}s7��Kı37�n��d�軹	Uwx�h��=^���,K��7�x��bX�'�����v%�`b'����9����'bX�%��.nn��]k{�7��ؖ%�b}�̼Nı,K�_\��;ı,K�fo�ؖ%�b}��5��Kı?"��ߧ��nBˢ]nh�ՙ��u���%s]�3��'�]�FF^��������k�x�f6���w�����ok����;ı,K�fo�ؖ%�b}��5�;ı,O�y��ؖ%�HM�gAwuWsWutZ.������"_{3|N�,K��_fk�ؖ%�b}�̼Nı,K�}��'`%�=Oߏ�۵wl��u���kDh�'��ٮ'bX�%��o2�;��,K��f���bX�%��7��Kč_��?QQU��r��wu�ֈ�'ټ���Kı/�ٛ�v%�bX�����,K��_{5��K�7����c��j�Y��;�7���x�/�ٛ�v%�bX�����,K��_{5��Kı>��N'bX�$h�,�K�������q˻���.���Z��F��6����tm���F���=3�ݖ�gK[��9��)u'\���Ǒ���[�]Q�k��r�\��3�&�� �!�(Եۗ/E�é˴�S�&�x��K��O�%������Ń<���-�9��x�y���qt2`�ql�x���孷<e0v���.�ٺ�At���>��GI�Q�ӵfM6��'���{��F64��^]���n�0鸦�r��[!�Q27Y�f)���K�&�4���;����&D�,K��~��,K��_{5��Kı>��N'bX�%�����,K���M��]�W*BJ��F�F��=^��b5�4F�'ٜ���Kı/�ٛ�v%�bX�����,K�̇��77n�.�������Kı>�ΜNı,K�}��'bX�%�}���;ı,O��f���bX�'��a�Y�j�zݓz����Nı,K��f���bX�%��7��Kı>�ٚ�v%�`�MD��߿�'bX�%�����7��[�����l�����Kı/���'bX�%������,K��3:q;ı,K�ٛ�v%�bX����aY��欜�s�gWb��,�k��;����ݵ�u`W��ғӤ9�¯b�������,K�������Kı>�ΜNı,K����;ı,K�fo�ؑ�4F���~**�e�*�wV��bX�'ٙӉ�{�1X���Q �D!�):u��bX�y���;ı,K��?o�ؖ%�bo<�!~!I
HRB�l�EIv����/sz��'bX�%�}�f���bX�%��7��Kı>�gN'bX�%������Kı?�{.��Z��6[�z�����Kı.{3|Nı,K��t�v%�bX��ΜNı,K����;ı,O{y!4f�7w�����o{�v%�bX�g���,K��ft�v%�bX��fo�ؖ%�b\�f���bX�'�2�f�	u&��ڙ1mش�N�q�����bO����B�	��x�����wCz-��qW}��oq���3ٝ8��bX�%�ٛ�v%�bX�=���g�MD�,O~��8��bX�'��?��Z�޷dަ浳�ؖ%�b_}��'bX�%�sٛ�v%�bX�g���,K��ft�v%�Z#G��g����U]\v\��F�F��Ĺ���;ı,O��Ӊؖ0O��tٝ�&Ţ�󦙥�o<LE���,��_�~��<�?J4��=	H�"�
&QU%�Rr�����&�RDp�8��%��i�zPʴ0|&�dL��8�Dȡ.��@6j����zo��$X��,A�	��> G�%����C������T]�mO �T|���P\?�}���g�,KĹ���;ı��w���y���h-ث�w�{��7���t�v%�bX���N'bX�%�}�f���bX�%�fo�ؖ%�:��~��(��Yݘ�h�����d�v%�bX��fo�ؖ%�b\�f���bX�'�����K�q������90��6n�s!�9�l��V���@��7��*��9�(��c�Zu�b�V��w�����ks��ı,K������bX�%�fo�ؖ%�b{=�8��bX�&{9��ؖ%�bx�]Y�5���-ӽM�{�v%�bX�=��'bX�%���t�v%�bX���N'bX�%�}���;ı,O���R.���jR��{�v%�bX���8��bX�&{9��ؖ?������߷��Kı/���|Nı,K=�p��֮��.�q;ı,L�s'�,Kľ���;ı,K����,K�b\����Kı=�7���jӤ��������oq����'bX�%�sٛ�v%�bX��ΜNı,K=����Kı=�w����Eӗl��ka60���F�-9Y+���.���1�&�8ׯRTXzo[��,KĹ���;ı,OfgN'bX�%���d�v%�bX��u�/�)!I
H]F��U��K*˛	��|Nı,KٙӉؖ%�bg��8��bX�%�fo�ؖ%�b\�f���bX�'��Y�j�{���m��q;ı,L�s'�,Kľ���;ı,K����,K�|���_�RB���6uUWW53uv^����'bX�~U��������Kı.g���v%�bX��gN'bX�%��g2q;ı,O�=����k[��%ӽn�{�v%�bX�����,K��*������D�,K߿s��v%�bX�����,K�џ���������~���M��UY�4�&����:J�σktvFM�m�-�=��w9ɃC�<�.�=-��3�3�q/���4������tnN�����ۍ���x����h@��v]�ݺ�1Uч���^Wel�͂�3ьS�-d���Ynv�)z���<�l<��!�w&:�G���nGT�<5��B�΅�մg�����7N;M����rN�ld������q��t���U_B@I$,����pr�ڢ軍�h��٥y�\ t�.���g���Zd�B��q��˶鲝e�)��	.���#Dh�3��N'bX�%��o2�;ı,K�{7��Kı/���'bX�%��C�9�wu!uw�]�l�v%�bX�f�/�lKĹ��|Nı,K�ٛ�v%�bX��gN'bؖ%��a0����o{��ջ���v%�bX�=���,Kľ�f���bؖ&}�Ӊؖ%�b}�̜Nı,K������J�n軻�F�F��/���'bX�%��{:q;ı,O�9��ؖ%�b\�پ'bX�%�����~��x�h�f�����7���xϽ�8��bX�ٜ���Kı.}���,Kľ�f���bX�=��?F�]��\:ւh�]��myѺӡ�eS�,����{3��7d<g���n��z��'bX�%��g2q;ı,K�{7��Kı/���/bX�%��{�,���$)!I	�gQ5UV������޵���Kı/�fo��P4��6 xw�D�K���w��Kı=�ߺq;ı,O�9��ؖ%�b|{5۽:�����u��;ı,K����,K���gN'bX6%���d�v%�bX��fw�ؖ%�b}�͝���#�ㅫ�w�{��6���2}��i�$�ff�pI�;��m9�2%����,K������wRk{��q;ı,L��N'bX�%���gx��bX�%�fo�ؖ%�b}����,K��ԇ٢�u�'���k=[]�IF�ӄ�,뗤�?�}�?�]A��E��i�;\X����V�{�̖%�b}�߻��Kı.{3|Nı,K｝8=�bX�&{3��#Dh�|�/�˪��*�.����%�b\�f���bX�'�{:q;ı,L�gN'bX�%���gx��g���{����ѫ�5ugu5�����K���gN'bX�%���Ӊؖ;�0q`R#B�1�BPUS]�"n%����;ı,K�{7��Kı>�xY���M͛!�l�޶q;ı,L�gN'bX�%�����,KĹ���;ı,O��t�v%�bX��zf�֮�l��ۻ���F�F��'{���kDibX����,K���gN'bX�%���Ӊؖ%�b{��޷uc�u���g�6���iky�'�mk�v�#)
nva�ݺ�by	�쾜�����X�%�s37��Kı>��Ӊؖ%�bfft�� C�&�X�%����/�)!I
H]\
���EMUR�o{��,K���gN'bؖ%���Ӊؖ%�b_�7��Kı.ff���bX�'���zԅ��黭�Nı,KٙӉؖ%�b_�7��K�,K����,K���gN'bX�%���a{)�j�V�h�5�l�v%�`%��3|Nı,K�37��Kı>��Ӊؖ%����$HF$b� �#B	"$�Ȱd� 1�A`.�{3���,K�̞s�޵��[��z7��|Nı,K�37��KıO��t�v%�bX��gN'bX�%�����,K��3�Z�H[uƺK�q�{�qt�ݴ�Q&v����&Y��Fw�{;��6o���qV�u5����ı,O��t�v%�bX��gN'bX�%�����?�j%�b_~��|Mh��4}����WC.�wd��1;ı,O{3����MD�/���|Nı,K�����v%�bX�}�����*!Q
H]_q�U5j�6]�ٽog�,KĿ{���;ı,K�fo�ؖ%�b}�gN'bX�%��ft�v%�bX���k���zַ�K�z�����K�,K�fo�ؖ%�b}����,K���:q;ı�}��'bX�%���R̚ɽ��Ӫ*����#Dh����#Z#Dh�=�gN'bX�%�����,KĹ�f���bX�&��dB"�����~��5i �h��a�譛9M�s�6y�����r���;5ٺ�Nٻe4���������/Z�71Ԃ���>�����:9M]>�S�Zt`�MwM��χ7vԆ���9��1���Kg}]�sڻs�Xh9�#(��uֳ(/��[�v���]�%�=�s�n�=yǞ˻Q�t�۱��۶�	v��pG/�;���.vza�km�&å�y��������{�Ӷ�B���]N��/�c��ዘ�l*�y��֯igv��o#&�����oc��>R�w[8�ı,O�g�Nı,K�g�|Nı,K�ٛ�v%�bX���Ӊؖ%�bfa0��٭��[�.����v%�bX��=��v�5Q,K�߿o�ؖ%�bfg�Nı,K=����A�,K�Ls��{ݺ��7��{��,KĹ�f���bX�&{�Ӊؖ%�bg��8��bX�&k��q;ı,Oj{3W[ަ��u��wo[��,KK=����Kı3ٝ8��bX�&k��q;İD�.ff���bX�&}�,ֳwS{��������ؖ%�bfft�v%�bX�k��q;ı,K���'bX�%��ٝ8��bX�'��{�P�ů=��<�� ���7J���>`�#=st��)�-';}��w�V�e�uصMl޷��ؖ%�b}��5��Kı.ff���bX�'�{:q�Kı33:q;ı,L񙣶o[��w��n����ؖ%�b\���;�0Q֝ı,Og{Ӊؖ%�bfft�v%�bX����q;ı3XJf���ޥ�SZ5�o{�v%�bX�{3��,K������Kı>׳5��Kı.ff���bX�'��F^a�tCS[ݲ�g�,KKٙӉؖ%�b{^���,Kľ���;ıQ�>�ΜNı,K=���Sf��u�������ؖ%�b{^���,K��u�����D�,K߿~���Kı33:q;ı,L�ܙMHY��&�kp�K]J�l�[�mwX�BöFwg�k�X���w}g�%��٫u�z֮����Kı/�3|Nı,K�����Kı33:q;ı,Ofs'�,K��O���ݺ����%�&���;ı,OfgN'b�bX�&g���,K��g2q;ı,K����@�,K>�kD��n�r�{n���ؖ%�bf{:q;ı,Ofs'�,�	�� B"�:9�.s��'bX�%������Kı=��3"T[��5�{���oq���{�?y��ؖ%�b_}��'bX�%������K���5������KĤ'����%�՗t�n.ʻ2����1.}���,K�fgN'bX�%��{:q;ı,Ofs'�,K7���o�?�gi��t5�e�zd�p����#n�\mG2���G������wh�e�SZ5n��'bX�%������Kı3�gN'bX�%���d�v%�bX�>�o�ؖ%�b}�B^a�u$���m����Kı3�gN'a� �&�X������,KĿ�����Kı=�ΜNı,K��?��V]U\�Uܫ1�#Dh�3�8��bX�%Ͻ��v%��%��ft�v%�bX�����,K�w���\uR�R�:�wV��#@%Ͻ��v%�bX��gN'bX�%��{�8��bX��M|�o�.g2q;ı,L��[���S[��令�����bX�'��Ӊؖ%�a� ���Ӊ�ı,O~��Ӊؖ%�b\�پ'bX�%��eg��kn�ڵaZ�)ْ�-�J�ݜ9VwJ������W\�ok/{Ve����}��oq�X�'�{�8��bX�'ٜ���Kı/��o��bX�%������C{��7���7�ˮ��Ә��{��ŉbX���N'a�"	���b\����v%�bX����Nı,K��2q;򩪚�b{��ٻ��F��K�z����,KĹ�߷��Kı=��8��`bX�g���ؖ%�b{3�8��bX�'��N�3[����j�o|Nı,��5?~��q;ı,O~�~�Nı,Kٜ���K�ľ�3|Nı,K�z�s�UH(��I�Y�
HRB���2ı,Kٜ���Kı/����,K��{:q;ı,O��l8�
��!�E����U3����(R�IZ$i���ld�p ��Q*�!��lAv�%H����T!H�	��lHP�D�e��_��w�C;�a��:j=�<����1�Pbp4����*�l�" �b�	FaVR�=�)iHZJ��+(J�Il�I������� �P�$a63N�Bj��Ռ�HB0�����5�&0�WF���%�H_<���ܾ��` <F�$Y�[�FC��!� j<� 겲���^ė�\�D�q!=��:��TL���iڄ.�T�6�4;F4��y��|��N���t�߷������: �$ 8  B�       �����m �a�ʙ���U/
�bW(�l�J��8���P&{r�l�-]a�Tk�ܝm���g�Ԇ�t�h��s�LGke�S=5�s�q��u�n�v�q�OogG[�s�3Mύ3��.������:��}����z[����A�.wN˨�lY�m$��:I.��ㄭٴ�ӗ4�2U㞶"1n�W���
��(Y��G\�Ch ��b�7�86���n���O���ی�@�gIj����p<�gC�v��WL�]�u�^*wz/m���ɲ��ym��m%�];�i)�o^��n�[[#W[@��Ԥl��V�է�.vk�ǵ�؟*R�))�[�;�Q�+��Uk&��66�l�@�ڶ�^����v�v�$�J�$-���'-M��,s�������9�uJ�� ܼ�rێ��F�]U+� 
��ek�VIUh	V��j������$6�"ڶ�`h7`�m6݁��im����pWKRv�Ku�7dv�]m�X	�x���]J�KU]UN��f�l��
� ��*ڵ
Ί�1v�gn�����9%�K<3y6ۗ¦�8��q��r���ɞ�����Npc���y��q��%��g���tr0��q������H�c8z�ݕyy�WWZ瞸�nnZ<�N�nwjմr��C�#=�z�rm��� �׊��k��Z�qAŷ�|���wnݲ��\OXβ��tt.,��ztݽ�%�8rlv����K*�
�4�a��\ѹ�G &����SS�e./b�+���T�eiw>3�n��:�[�-3�õ�Qvֳ�r�ǋ��7K˞I�����Ll��]��2��r<=e����k��3���3on�h�
�v��c\��Nb;q$��0Xe�F�mq��Ʃ˨��jl��t��H�7�]	���:���Ӵm��=����奺��$a�Z���I��M�q<�PO�Q� _/�*�_<��V�pE؃�Cñ~{{��H-�
5�M����\{m��^8�ֹ6���r���c��g��W\�ܥո�ݸ��p�u�+u;��)��sRf��7+Uv���ȯG�C\c>���M�h���8�쮵�Խw��X�6��rvsg��V1�^�m+�[ukr�����nܱ�<ZJ���bw[]�V�`v�n��ry�࢈�EΝL�s��g%���~z}����;4r�tQ=/hJ��+�n�aD�p���^�Z3pj{~���/ݮ;}�%a����8��bX�&}����Kı/����,K��3:p?D�&�X�'�g?N'bX�%���<�%���&��f�u�nq;ı,K�7��Kı>�gN'bX�%��{�8��bX�'��d�v
6%�b{S�[��R��UrK��w�ֈ�#G�}�LFı,K��2q;ı,O}����Kı/����,K�Ϸ����M�w{��n��q;İ ,O�����Kı=�s'�,Kľ�f���bX�'�����Kı?������L���Ew�����oq����d�v%�bX�����,K���:q;ı,K��o�ؖ%�b?~Gc)�̼��y��نX�,V�|a��3��3q��g��MiI�}����/}��nݺ�n����'bX�%�}���;ı,O{3��,Kľ�f���bX�'ٜ���Kı>׌֡�L��SSZ5u��ؖ%�b{3:q;��@A�D� D�~*����9ľ�o�ؖ%�bg�̜Nı,K�37��Kı3ޒI.^�JY���z���Kı/�3|Nı,K�=��v%��bX�ٙ�'bX�%���i�ֈ�'߇��ܺ���Q*��艞��� }�x�x�>��Q2���O���$�łdcĤ�oY�~P�'�ߗ��׀z� ~���Z�@w��k��Nl���9�X$k!N�k���7 ��{�����Qp��C)}������, o]����BK脡z�����o�$��d�7�#������`z� o^,��&M�b�)M�ʫ�tU�ww�ϯ �xdj��P��6(X�Rqt�HDMd�
!H!$��&�޼X��x�ys77J��IqwwWx�Jg���ϱ`z� �x���QD�v�J��UU���ŀrIB��}�;��4޳@��`��I@Ba�ۉ���.�R�`�d7Y�g��\]�M�nc[d� n��5��f�u�4޳@5뾈�
?Hw>ŀw!�	�ʛ�7u%"����w�
!)�|���ذ^�ϡB�7������!*�ԩ���ϯ o^,>Q
"���������rL�8ȱ�&��~�}�����w��؈�B�$���I@�����T���~�$��ku��sf�ɐpN9�׬�z� ��h�ŀ|�O�������E �����ou�n���9��M�W�щ�<�A�"3�u�N�����w�7LՍH��<�p�������m�^���٠}x�a�E��wwWx��Ϣ>J""!U}�b�ﾚ׬�9\���ɋ1�m�4z�`��Ô(Q
�������;� ������s4����� ?6��(P��|���;�ԓ$��jDńNM ��h�٠u빠�@���g���j"i% �$�I5T�:3��� Ӯ�8��gt&����ט�� d�6�y��lz��KXۯ{�c�^���=��q�YX�v6�����p�h�2�+5[l m�[��.�jr���z�s��pp5�e��[C�igt�y�� 7\v{�索�vw[�4�=rr�Y7k����k��xuˡN�01�*�hn-䴹;E�;�4��� ILl�t7+jJ.��F�.!;A���m�\h�-�nFG�gr��;je1C�y����q�W�m�?o�7� {u��""}�D/P}�_��w���d��sWeʩ����Y�D�n����0�n��P�Jd{NI����]�VU�sv�w���`�&M�V��X�ѳS54�UISSE�(J"%�q�����x��o��t�j���.EuSv`�����";_~_���b��ـo���U(�v*�J=u�ݺ\J����#Z�[�] \��Ju�m�x���bf7�'&�{���[��o��菔BJ=@>� rO���LӗV9Uf6��}�! X�%#�}<`kn�=x���Q
�#���5uj�RU��9���x�x��x��ضL�v)R��M�U�
"!N��]��ذ�x��l�?Hۨ�I&���LNI�z۹�~�������>���yz�4/uR<�$�a���-mS�:���Lݴy�9ö�F�xG�{�5�$�	�9$�Nd�8!ɚw]������D/���`<�U�@�8$���wYM�g�$r�I�w>ŀ=׋9%�*���W��WU`UZ%Z��0?w�x��Xj�	)N3"V���w���}ܖ<�Q	�o&������y��s}� �;f�S�Ϯ������L��բn�`u��>P�P����l���^,�ۿ?���:z�[kku�t���Ű�!\�m;Ϻo�WU��j�Hu��i��v�YT�VJ����z��6^���^/�BQ�;]�o/�fn�*U]�sUf�����%2o>ŀv�� �;f}
!%�G���F�NB&7$�;����_t��޲�+l�y�ӱ���
ʲK�X�$�����_�n�aDD,��")��� �/aʫ��i]+���j��m�(P�']�w���s@���\1��&����nLE�=4�3ۡ-3�#��Y㪘:�{@��J;��;�$��ɋ&'!�r�ɠ^빀?;gDD(���|`���'�Qv(��MI&�{��|�Z���:[wy�P��(QC��L�NY`Mujf��󯾜��0��� �^,���T��i\�5Us��B���� 绮�n�X$���� �8�	���PU�$�Y�l���P�Q�JO��/󯾜��f�(���Y6�પ��h�3 �;�v�v5nW��xt��x녭8֍��ֺ�>�mnv��mї/[n1�7@��L;��q��p�3�"���ыm˒�t���]I¹�wg�-���=a��@�� L���@;@�e����s�r�>'^�;ܛ`E�gnv�#cOt��N�	�P�����[i�ɷ��c:^=7o\�ݭ��tj�\��.�h~
�sk[RPݑӲ� 㷩�e��{PU$h^���ڦuݫ9|�gp�'����RE�|��s@�m��;g�Q�A�w]��檺�f��Ȯ���`���В��w���w]���,�"S#�qҪ�\�+�r]�N-��Ɓ��&�����/��@�[��G"�1�MHh��hz�X�7X�BS�� ��QS<��cQdX��M�[��U�^��t����&�� �M��������!�N��k� ��XA����s�Ev����kp�o��w��dz�F��6�π����{�)�r�ɠ}�w4���ҸȞH��]co���ȁ@�^C���)E
���{;w���$��g ���}
��9wE�M]�"���ɪ� s��x�o(IL��u`��|���bJGlrI�w������<�ف�J"�"+����>uɿ�D��FI�G3@��z�?����? 纺��x��-t�w5sjl�����vꍆ�0V��͢×#n��W�YD����#�2r�)U�.i\���UU��7��l�N��x�_�}׀{��&f�j����+��� �n����=�ذ���@��M ��/�X)�<�Qɀ~m�������v�/\"Q$q�4���i��b�Ul,��9���ܨ��T2"�	x/"d1�g��fݴ�*�L)���M4�TJA ˪��ڱ�n&N��]�;_���HH�$H�+$*l�B�)��d���@�YB(l��3&��9e�C��Q�7���^�sw����yG���T�%�%��U�2�A9T�j��pcU`2�7):(`��61��M1<\��Ɲ�� �H����,uI��p ��������!��'�	�����H;$����5���mH6UU1��M��J��f�{A�n�s�o��og�{M�y9u�9$!p���%�B9D ��4��"(��WJt�O'�B�������ׯ ����sw(����V�>���(�����e�w�~m��7�h�e�.iU̓uw�n� �>��_��_����, o]��lr��ҕ6����}���vn҅�t�J�H�z��.�������k���հ�츭am��~���������ۿ�B�!����<��UPL�]�TT�� ��,�)��}x7|`��7������X�Hē�H�1����׀=�f��]����?:q,�(���T�jj��9$���0��׀?7�~���Q��%��n�w����6�1�MHhU�h�ـ�� {���Q	%�L�r��)$��;Qv�o"�c�%�6}l�jv�]i �A�5��t�������x���|��� ��� �m��λ�7vLY,Pq)$N'"��ٿ���?u��˗׀?V�ϔL���e��4��B�� �w������DL����>��?jql&f�]
��&j��D)t�����p��x$���N�;��)1�7rhϪ�?���Ϻ��O� ���xDyi`خ@������,�w=�
zw�чtWi��غu9���eX�Ć����n0��ۖ͝nw.{�Ν�ԱGS݇T�mg`M���_=�x�
���u�:�c,�iXq(mͫ#g�cV�a�S�g�<d�зh���>m��P\���R燗U=�G ;�m�֓�:m�-t ݴݕ����v֮έmy&e�1���!ܱ�/��<������������G(�k	Zc;b�/m��)���������G�L�D�H�1��������]����Z���E�4E��;������N�>�X��u�(_(���&f�j����+����:{����]a�Q>����N ~`�;.ʛ�wj�M�U���k��=;�X��]�����%��G������� 䣶�O��]x����u���s���e�Nm�k]�F����8�e�w!��	�mv=����Ǡw��@����^�@��ՠ}���A%0&1�D��@������6���^rOoپI?��e䓼�Z�9�7l�����4�]��M��S>��X�� �V��dě��'��z޲��[4��w��D�o� �S����WR\���5V`���DD(t�u��|`z�h_'�wn ��o$n�5�S�,A%�����c�ͱ��g���n�4��R8�$�ɠr�vh�)�}�l�D(� {�� =�Һ˺��.h�$�Ǡwt��������@�}c���	L�܊l�(.�nj����7{�`����D@nֻ�wm��CHVʺ����ʺ�X�%3���}u�n�脡%;�ߖ�]�7%L��&$��;�X���h�����hL��)��bL�o�Lh��4l�κ����bv��ю�ݕ�w��\ϯ����w��+��X�2Fӑ���Z޷s@>�������Q�����Ldp����P��wu��������DB�7���L�SwT)�.��� {�� �z���D%2۾0�ذ�kɛ�R5$��I�+�M��4��<����ֈ!�DX�|
"��^�Wu�xF�\���U�EY75wx��0���y��wu�/l�\��d8bi,#y1c���f�v�(���f�sдC�Nݓ=�9���W5quv`�l�ͻ�6^����B�Pwu�`��I�������՘��x��w�n� ~�f4�(IUq�x�cx&�~���=�����@>�l�=�WX��&H��� �׋ ~�f ~z��DK�}w����C"&,pd�4���w�l�wx�XB�"! P�%}��{������?s��Y@Xn�PtX6�u�;��m�.�	�6��ލ�6ușݻqnTK��i�m�]���/v�s�N�H�m��ʽ��Bd���T�l��l]�bw"ruV�:��©�rm�; +�k(u�R<���m�tX��rY��l�z�N�NL{��c;eK�_�v�6w:W[<��'����<���v���y���{�
�p�պ�Tp�<r�l��-�����j!UU�[�׺��7c�b��������]�,f��(~������@�u��/�S@�uԤ���q6G#�@�zɠw����\��k��&C�N�����ʢ�������X�k�>��}��p
�_�h����6H�s�G3C�(�%���p�wӀl�wx��0�a�2��	��qhϪ�9^�h�)�_>�@�h��'�4���������h�o>�31�ȕ�q���,ja	���{�{�]�Ys��F?�o����M��4����y���2��v]ӕwx��z�y�HH x��DM�՟� �S��6|����J�v+��SsW7k �V��?:�8}�D˝���ŀ~��Dӛ���.U]]M\�r_%[o���������`��h��U��	$�Ǡr����D|�#_}��9�}8����>Q��߿�Gjw]��+7cx6�g�� 4�4Pѹ�4m��2bo%E.`�rO��Y��;Ϫ�>^��^�Mڢi�	��8��RC@�����2n����u���ـ~bIl*�U�533uu�{ծp�7w��JҘAe�`	 <�E�~�I���`��Հ~�ՎEv]�]qFԋ@��ɠ}�)�r��@��U�}�WFLs&<s$Ȝs@��S@�!%�%o��7]���uxβ��63���ŸH<^x˛���ul+��;��:�9qۯv���<��j�18�`>n�z�� n�WС~����{�Ƀ�&&c�#�h�����[�W�{z���w��(�2n��ʩ��	��Š���}�f����H����;�����rH�R&�ێ`�7x�n�z���_��X����J:Y��U��7%UPu����1I4޶h���������������:m�8oK�� �%c�Ű��Ԧӿ������љ-�"�4�4�n׍[,Ҧh�n���O� 7�������#�����~�~mL��L�(ڑh��� ?y��n��=��9���GWE�Ly!&H����h���=��h�����Q��@�Q�1�]�DL�}x�>� ����|�g����?+ph?BX�C�M�}V�{����7x���Y�W�{���/��һP�U�%�^�m��6���I�bhF֠J��[�Hh(�k&�	�70r���\������)���pq	�LCb15�0���mU��iIN�V�szB�b4�Cv��Ȇ�V��ۧ���.���A�� Ұ �    ��       Hp����֙�d�)�Q�k�7WI��ƍ�$%��E\���gu�X)�/G��Mq��1��c��k%s�3����ksf��]�>����c��c��4��\�ڸ�g��f*^���v�5�����	��=ln�c��WS�0�ظ��7g=�I�#qط�#��u�<+5��Z�[m9�����h巪S�h�[�m��izy��D^\k�m�z��, �:�3��kZ�e���ѥ� NKt�d�+ ��H�0*��ӎ����v�#7(��<s��U�M6�ٗ��EYWd����u�P
��WY�S+URF�OT���Ӌ���2�N��������D;��5����.�\m�6� R��nն�mKZB� 9�l��А[nٕa�16�:8兹��-V/Z枝�غU��눎7Xe�մ�i�Wd�p�d�PJ��l�Un����j�m��RČ�gHl���^f��U��U�j���.� ��4d���Z�B��i�cqI��oR�u�W�W�!�l	,2�L�R�-�kd$lq�i�=�^��q��r^bZ���sˎ։�+	 ��.�.\�n����;z᧬�gѺ\K����q��[8��z�ݻbPyz/n0�l1��pq�]�R�Gk15nM7Ӳ���u�V�^�p�kύ�9�[q��;�L��	��t�g\��ڣ����@��l����6�T�9�+�$�ۜ���t
-�K�UK;q��u���d����r l��`�'�Ȇ{���<�\Tu�@a���	BY�p=��Ӷ�c���I��ˤ�Mv�+�Ș�s�r�m`۶�g�8��ke*k$�l����^�V��e�n�v���Qዶv�s'Nlc��ݻ���Ǥd3�S�1�'P:��ø �'fy�l��ۮ75�H)ō�P������8!�q.�{j��7q�qs/Z����Jے��C�q�
��ZK�T$x@�_�|J'�Ay��yQA��jo��N�F��S�����t�iV�uΞ�;N�ϓ�cn�ug��tZ�g���ƞS��u-����J�0���Mh��]��8�S�R��������<Z��q�r�l�ƶzj�X(3HjК�gv�8(NŲUv5��5���Lݶ5҇����G�h��r�ճ��9G���;n1NϯC�lg�r��&zjx�<'rr���A����m[8l����p��{{��9[P�
7K�Wd��G=Э�5����u������.S����L��BF�$qx޵� ��� ��_%�n���:~��������.��������� ����k� ����D)E��16�~ɄN9�rM ��~���� ��s@>�f����J�$���;Ϫ���h׬�����{�^�\��We��Z������ �n� �"'��� w>�}Z� �P��~��q����m�u�ќ�=�]�����W#D���3��meD�=v�����O�b�W��\���~� 7����s�Q�~s@�����dC�jb�jI���6���(�0��>�s���?=�g��*����(c�	94��Z����Қ�[4��Vl�S$#��Š�\�>���z١�3�-˿�~�FG�LNF�s@���@=�f��}V�wus@� �=�ݜ΢�+�v��1�q6���L�\e<����:�/W���v��rW���w��@�>�@;���}_U�}K�D�ېBmD��@�>�@;���}_U���f${�����Bp�G*��p��x��<�r�S�%j� S�����
ITu�}x��WU�^g:F�s#����h^��{]���8$�Ъ���x���h��Jb���@=�@�>�@;�\�>�)�TgWI�b��m�6��E��/cI4g�9)C��,=z==OB�~�}󁍴�H� �BRO����r�Yx�Z���u��bȺ��vGQŠr�Y4��Z�u�����$r��ߣ�"AĦ'NI�z��h�k�>��Q>t�p�}w�=s6��*!1�O�z����>�@����5B�Q�$���P��-�V�~�IL��A&��@�Ϫ�*�Y4��� ��f���U�1D�b����g�Ʒ<�z�d��*�K�\�ֶ��9�v=9x�b��bBp��(�_�u�&���W�{��g��=��Z�W��(�d"Q����^�}�@�Ϫ�*����(��}
��|O�f�ʫ�椺����}���Z��B����x�_V��m��d$h#�@�Ϫ�*�wx�����|��{��X����"�S$#�(��*�d�?������߯^�}��	� [��7@]ܩ���l�9]	3Nۭ�ө۞y��+pr��ny�!2������:�g���=�pm-\�-������!��oiv���ZS ,],v��=��گm�a��p��et�y�ϴeX������|�}`,mf*,x�Oi���q�Hnѣ���vr��d��{mb:����
���qnwl�5��nr�h޸��_OW�%ph���s����{շ�>~�6�+<�����]�
8��C���J�#��&;iմq�ȼO�#���q)���P*���^��~�k��G��}w�s�D���U���jG�^�@�{��*�d�>^�����)���(��@�{��,�wxr�3�Ӏ�׀~���dNQ�I�U�&���U��f��������;���#IGY�PnI�}��h�Y�{��9[d�*3���?��y��.|ۣ���尢�S���^͇s��l�^��]su�H���j��Yi��� ?{]����B_�=��p
�Pcm~�L24D����j����MB�9�c~���{=�@;���kM���j8�nM �n� �>�XrJd{�x�}x�7[�rE�7�9#��}V�w����� ���JaZNE$�rO椬 �7xBS�}���?O������z�z���S�m��rk(��D�z-�	Wn\s$iۤ����<n�:m94�u��k��}V�w��ݗ�Q��srhu�o�s���^���}�@�̯m�!B'�G4��� �u�no�fL��b�K����W�9�����*�F�8�n-ى^����u���M��ZW��۰s��")&�W�� ��S@�}V�w����`���g��yS�E�H�/dݜ�Z�9��N��\�d�wRs�ǉ�}��rtĵ��_�<�����8��x��� =��9"�5�I"��}V�$����4������ċ�)�x�ɌmI0$�@?u�4�[4�M�}V���GQq�(�jI�����_��h��M��k��H���Q����f��˄�@��srh�j��}V�w�� ����e��~o��#�I�U���	z���&�������`58ꉟu��moޗ_)�պ�ۜqO��w��wY�z٠{��s�Q��8�C�)�{�� ��� ��T�=��o��H�����Hۘ���$rh���{����� �u��2֛܀9��G#���L��u�����V�V 8��u5v��5�H���� �h/Z�/Z���P�d@IRI$�I5R��pa����E�;ED�s���۷Cv���������zn2����]��;F�o\^{f�f������p�ۙk����ȯE�<u��dl� ���g���x��]Vņ�Qh��5�6#�����'��#�)�9v�l=�I��l��5Y2�vk����F�5��d�d�[�L��U�Yn�H]��ms�N�g%"H $h���*�e˄��sDc3L,�IƕX��wLX��X��n��Au��=�$�Y�cm�?�q��߿M�ּ ~no���_}X�)/�U6��G�M��^�_Z����^�[�h�K�� �$�@/Z� �����(��UG�w׀9}Xt,UQǊ3�8���zoY�yzנ�S@�|�m�d��W%�� 7���Q�C������U�W��^O1,�?����$8����)2;L��q�U�8��a�h.�v5�\ܗe���x��&��9zנy[d�=_U���x�Z�f9ۊF��?����CpdY��l�՟~�Ӏ�� ���ϡ(�����몚�<�,K"��4~w���f���^���&�z�0XWXےO�Z�䢫��׀t���t���ֹ�?n�%i�DH���)&���^���&��}V�_[4�Σ�Oq�EXFՄ��ܑ�D6u�칫CJ����A����}��_X-�m͙�?ͷ����?�}V�_[4^���H�f(�2HB9&��}V�_u�/uz^�-������Ɖ"�#jE��� ������
�%�QjbRd	>�,���C謁'��]�}�W㚪��1�6B�����.���{˩�U$;�˻i�ݶ�Ӥ�� �c$���5.��ۮ"rQ�f�aV��0t��-������J r�)��N�,(
Br��/T��󔓅1�,��A�9H`GD��KHJƚF�HjBI4��5���Ȝ�^mYVjU�2'*��XZ�t��bQ&���@��E�we2&D�dL�]�t�&i��C"�]2KR�h"���������S((��Hp�2R(� �Q3z$q�ӝ臥TQ���������i
g�<(���L�e
��J���2P�N���\�*���e���(A2�"J)9Hd)gzR����
z�
��AA7wgP��G]Zj�x�.WP�hTUvJ���eP:���RXLy�����0�Q�aŀ*TP ? ���F����32}ޝ��}V�{�+X㑴�JI�r�W�w��hW�h~�J��4�~��ޱ� ��q��,Z�M� o����� �(K\\�֬�N��!��N�[lCb����SX�:5��	�ym�=��iF�bx:3T��]Ӏ�w�l��|��9�\�}�ͩ���
SWWWUs��w�D�U���{����v��؉X�FH���'&�˺��e�@��M �k�V��vLښ.h���n��(�{��8��� �k�Q
"�
%9�����>�G�8'!�jB(�X��D%
^���9o� ���N~���3�,]�ۧZ|g<mv�;cu\��+�p+�kl���/\�r����#nL����9{��>����]� ���<Hr4�#G&�w���z��}z�h��4�-x���M�D��>W�zץ4������������O"kɊHށ��M ��� �u�{��@��LM�bi�?��h��h�^���[fn�I�k޼�C���I!�U�.�� � :(%�.�!M�VZ��1&��{�n��Ie B�v����o藢�|�����8�;��n���Y�Zv��`�Ʒny�x�ӻ��gyއv�R��L����n�oMmp Pmd]�n:���48�*�����;^I'��+Ѥ����Rw[�kÇ�]H�%۱kn'�On��݈�]v�.�u�nv�v싐w^�l9�Ɨ�f�-'W]c�g�v�!)x褢���+���v��.��#M�[�sugC��}���ػ�+�`�S�qz�fQ���~����m��X�����l�;;.Ea#���&%$�;�X��Z�޶h��h�D�90r��F��@�zנ��@=z���U�{�J�)��择.�>��wu����5mmZ/Z�뜝F%"��dNM ��4�}V��ֽ ��4��"�j�X�h�s�G78�J���[2�y��A�ɟN�ŷ:�q�^oZ��U�j��8ϛ� �۾� o>� �e��q�D���-��{���bQ	8��Hy�� �k����8��Lm�@C�LĜz�u���iВ��T�p;�XD�M��Yc�6��������=q��@��^�}�f����#�D�I19&��c�^����h�Y�u�u��'�^�m�Jv�۔�9��l���݃���v�G���.9�gq�ì�f�;-�f~�O��ۮ��]�K�� ����U�қ���.�����IDL����=Y=��z�g'q#� �T\�� y��Ѯ��
�����u��Y�{�UF�P��n
G&��3��9u�@>�Y��� ��rD�Ɋ!dn5�˭z�u�����[.�J#h��MpEJ.ˡ������Zϰ��#��<]���v�f9z�did��ɘӏ�[�h��@�ϕz.����+'#�q��@=m��|��9u�@>�@�v\�ܒ��917&���*�]����h�٠}�PEp�%MU������Q�]>��7׀o�䒠tX� F�da�o i�����R,`1�A�)��T���XE 2$`B1c�����p���J���)^8�1LrA��z�u��l�>��^�˭z#/<c�7�����&}pi��^���m�Վ��Fـ��=����G#���ǭ�@�ϕz.����h�eor8�&���ɠ|��z.���l�[f�vx�۲F�b�Y���l�u���Ô%&�u�:έ�$Liآ�ɘӏ@>�f�z�4/q^����wdu47$n��rI�m���E?�����@?y��<�D(��@�]�xQeH]��UU�桧hΈ�Lv'P���8	�x�^>�Z���U�姁��ۮyU����x�ni���c��wGh�ڵZ39�9R[lV4m˲�'\�m3e�\�)��%�:ۈ�{]���δ�	{ M��n��i��㛩��7$u�uw��$[%ݲ���9N�.,�\��]	�gg�S����	����M�*��]/:�
���1�[�(�����ûY�<_�ﳣ�oA�F��m�;R�&w5�������2���U�ۦ,��8�q�RbnO������9[^�}�f�u�h�(b�&G����U3WX�n��2����׀~�Z� ��J�"r$y�jG�z٠���)�y[^�}�ʑ�PX�$�hu�@��JhVנz٠w��+�ɑ�&���:S@� ��� �h�B��h�F��G�l�W������5��gtNR�GvA��[<�T[�b1���o����@>�f�w[4��M�HSRɚ&�ZUUu����,J(��6۽�:S@���1R)1�h�'$��f��)�y[^�}z����NȰ��&$��>�4+k��Y�����T����2ccp�<��@>�f�w[4�����]߇��������ֹ�Xט�d�M�'.�����;-e��+�n�硬S�9���~���w[4qҝ� �j�w
�ŉ�(�6�ܚ�r�}�Ӎ˭z��h�*��&�<�ӃjG�{���<��E����`���+^�g�x��}�oN~�T���(��1HhVנ[f�˭zw��[�A&)24���]��������=:�`���ײ�ՠx�h�:ִ8r:-9^����\�m�M��	5��/&���� Mɠyu�@��S@��^�}z���r6�1�8МI8��%4.��׬�=�ՠw���P�,Jd���yu�@>�f��v���M�r�����ғ$���4��f���r�AID"���E� j�}��$��d��[��IA6�ܚ��M��M ��f�}z���0@ۮ&�L��Ɔ�������;*s�2Y6���0�:��lH�[��tvZRG�`ڀӆ��Ħ�}�@>�f���S@>�7�;��bYD��}�@>��@��w4vt���kc�QH$�&O�z�[4�n��Δ�<���ݐnc�&�	"NM�[��{��4/uz�[4ge��`�bQ��q��=�Қ������}��o{��ޞA�F�xhN':):N�����L�n�@��$ C@B@)B��:���Ґ�KI�$4@�Ќ	G�C4��Gn�@�"FHB��#HSA	#
�"��5��(�/�f3"N��yT���11�i�i��J鎴��I�3F�i�E4��T6j�$�
�a��6�'J���)9Dֆ������������F!)}�89�ci�p1%*��[d/RP�B1 D`�	$#h����CCH��:��T88B�*��&�m0i��K)X�v!8Ri�11���(N*�52N�l���h��bBB3���,O���~Ki�� �@    ��      Ą��m��I���!5�����W##;�z1��q�\�Uf,.UK�ч��c.�nKt�qm�V����gl�؉3��w�ŭ8�{c�a�ʫ�c��v����ƻݸ���q<��iN#a65�๮�R��l�m�z�q�xݳ�%����m���a�s�gX���O&컳�ƪ��n�ρm�R��Q��,9�[��P�h)C�\2ɞ'���ē�϶�&V��<3�!Z]���<cGWkg��v.z:�h�dTk,^=G v����3h6�Kv��s�mp�F�#ŧb�P��Ʊ�B��S��*�	�m�u�T�UR�m�t�R�mٮܱ8fNȢӖ<��rl#)r�q7��m�wc���Hٰ  �Dڶ�t�ݦԐ�����Xd�ۭg	|�vZF�9s�z��6ֱ�Al��p��.G���}�j�3m�ye���~�ꪩID�
��v��mU�����%
�e[��[j����dm��l 
T�ڱv� ��^�~W�}V�\��֐v�9��F��rŮ<�6۩@�	8-�Hu����5Z���Q��*�u�7hY:8��?>�'�R�9�\��h�
Z6�� �	����)�v�72h��M�r�ə�VO$p9 ��U�f��Ն���G�Nbv=-]n=��A��[W�d��G^��:4���c��n4�m��V�k�k��Cq��L+�h�n2���m���7d�㸓�Ǣ���N��S��囱��\r�Du�J���'����#CGjab���]�Xśb�ڻm�m<s��yؼ�q���5O.ɫW&�64]&������y���*���݃��0XL�RtE���n�v�=����,pQ���b�	�8l��k�������&�	�[Ӻ��{.��t	��9�a4�� �f�d�v�nx��NL�cݟ���[P��n'�k����2��`�z1���ٺ��̼h�sk��vSm��]���/�"�Q�T6y�]��`���QS�<��?�����wO����,��͚�c+�v�3mpAte�A�snzuH���X'�۶�2�kg�������L�l�<>5�j�>w��q���㷴Z��8�i�����	ш��[˰< m͈���j�K*n6�e��di�<�qst]�jv���<�"s���c�W[��#�{�Ż=�C�;`�&��5\:ن��7[��:[�z�É�����wV�����099DG\]+59zQ��9lV�c�1c{vRa�ky��6�<;��_<�&7����� ���޷s@�gJh�J��Q�'�= �[4y�X��f��u�B��C͒�9]H����f���Xkm�r���]���?/���>�QT�9�j��Қ��zW��=�)�f��S4�f�$��7f��u�tDGW>��n��6�ـ{S�ݫ	Ud�V��W�,�q����N���f9�Q��]�s�Ĺ�f��\y)�m�~�����nt����^����#q�um��r��������D��8+�|h���*�^�H�\���L��6'#���g�@���@���z�hܡ�Y"��<S&G��@���@���z�h��/r��Y�c�ԋ��*��ץ4r�h�k��O1,� �A��L��x��Q�����.5�$lu�C���.d��pI��8�m$��=�)�[�S@�^�U��vU���H�Lm@rY�6�� ��u�9m��v�舙���)�4���9~���W��rq� ȶA!�K���߳��h�Q�Lx<$���q�[^�|��ܲ�^����5L�������������9%	.k���l����u�6	��SX��Yk�[un׈1���g:��.�X�롕�,�GNІ�6�:���(�?m�?��~o���U�Uֽ��^�}T1*�$��&ի�Uf�V��I)���V n�^�{,������Y�c�)&��*�^�{���YM�Қ�p,����U\��L�]`t(I%>��X5���'��oӒ^(�;�js�^�}��MRE2bj܏@��S@�t��WZ��Z����lȂN#���1��t�a('m�W u5���9��[���ev9��mŞ+}��;�4
�נ|�נ^�)�w�Q�5d���Swf �[��	D��}Հ~��~4wJh��裈y&�J��?N�X��r�Jg[�0��Zg��b�bm�I�q���h��*�^���^�}T1*�$�LS&G��@�t��WZ��Z����Q��SC ����2����Oi� ��mV�	�:8������](�7��C�y�ڱ���=OmZ�hv���.���p��]v���6����M�kk%KK�El��E�-V�&-�]�)���yJG�'�<QˍcQ\y�F��7���Kb66<\`,]�S�#�W�k^3�-�9�y��m��X����u���V�8�Nbn�nu�@l�u�۷HF���%s)�V6�t��S�t�d3�v�!��ȫ�8��]/�ch�8۞���"li�ő8��P�C�~W�z˭z첚��4��Hu����(�MǠ|�נ^�)�{�S@��zv\�e$S&&�����e4wJhu�@�u�@;8+��h1A�qh��hu�@���C�������/_���H$����hu�@���@��ՠ{��@�{�ƿ��ݧ�����;�����uv�����>�-8�,�
[�4z�-eUu�3~ k����npm78�n�Z��s��Q*��vIW1����՜�rES�wV�WZ�s�h�C�BO��jՔ�� ��s�9���&u�t�7?~zުTŊ8�LJ(H��*�^��v���^��v� �vu�"��EI��s�hvZ�s�hu�@��Y����77"��ufۧK�
�Ӝ�ҥ���):��ƻp)��-�v:crAbj���We�@�YMη]
!/�����t���ɛ�1BLq��)�Uֽ��h�k�/U���I �K�'���O���9$t�t+�i�P��V'Y���S@���1��(�"E#�@�Z�[)�Uֽ���j��2BDӆ�y�����*�^���h�A��ol]���`�h�؜���Anny��Cnv|\c.�ד�cI���cS&F����hu��5�gB��������*n��LJ(E!�Uֽ�)�^e�@��h{�MY��Ɣm$��-v��Z�l��U���(1a\����k-z�)�Um|���͕��U�(F�D��aTK ,���=��$��. �Ղ�����/YM�k��s�7Cu�r�� ��MpEIsc	Z���9��*�BԄ�\�qd��r]������r�"n(=��ͷ��������Z���������c�'mLd�)�yڴYk�/YM�k�=��#V�b�!mŠZ�^�z�h[^�yڴ�P��1�<ML�z�)�Umz�j���gu`��頕uvU�]X]Z��� {M� �� �x�)\#{�n�_��,�T9j��T�k�=ϕ[^[o�n8�՟C����b/.�흑��w �����<Z��ƽv��8��x�z���OO=2�ldaJK�ź�ط;ڀ�wn�`V�`�ր���N�'nN`,�m�h���x{t\ϫ�C׸��;s�� ��]��Dm��v�	&b[Di�T9���U\��,����ۜj�N�s<������{��_k+iI�e[�����UN�\�ސ��Mb���C�ŷ/bgt���=���1\�)J6$���?�Z���۹�m��\J&,M�&�$q��k�o kn�-��&����̴�Q��z��h^�@�������emli���"_4�Y�9�� �F��������M��q��fI��*�^�՝^�z�� ��h>���Ǐ��c{�Ov4�j�4�)Kr���B�����G4;g����)�,!M��/�~P�v�{��9{����
71(��248���ʈ��!�]�|�`��X��T�A�H�8���f�WZ������h{�n�c����l�@��zVuz�w4�Y�w��-o��&��G�ugW�^�s@:��]k�>���e���1��{`�r�j��w]^:���u�By�S�dǏ	���q#z�w4�Y�Uֽ�:��YY�	�)�#��z� ��hY����h݈��i�(�2H��@/��]�=��M$B�AT(P��Px�y�zP4z/�e� �1��4�cc��bC
y���_~����RE^X�M���D$�	,
�1�ώ�ݕ�XӜx��I4�>�M�=������q���en���%�tH�1uy＝_�bp��Yr�J� �#�`B�#���*8QC����q�6/\�T7�Ĩ�����c����V:��ӄ9b�u���k4:%4�H����(P�	JZJJJB���(���H�Ī���ă=�����G�U�r����'|��+�2�n�!�7=���(p���ȁ�F���$��$NA6H�rU�b��q1�41�h`���/7��dSxv�XJuA
I��4^}vbĵ$�
,b�M��!k1P�!XB�� Q�B�6�����k�$ �$�=F*��hQz���P���!$$a	$����@�5Dd~�����X����[�����w7EU]�|�)}c��9�ŀz�ؗ���h��pQ$���/u���f�_[4���[�8���ܩ���$���x�@�Z���,(&x:��m�7Q�rN��t ł�m6&�`�w�����u���C������Dq5$�z�Z�s�7� k�y�Q26�I�x8(����I&�c���}�s@:��{����p7^$b�������m� y�r�		<�Д�KKKh�K	VXRJ�FU�%P�%%�"JJA�iHP����%%	h����F0�RRZR �`B1��$#@��![-��)Z��
Ě%b�H�B%VRIHRR�X���Z��4me�Z�,���`B�c!*�Rҥm���-�$����-ahƲ��PУ�3���}�59���'���u�h�l�:��=�)�{:�� ��$"OΊ�!�͗N�t_am������^����['=�q�q4�L�NI���@�S@����[l�>�\�"H����wxi�3�L��|`wu����ܡbsj0D�7޲�m�@=�f�nYMީJ�"4�E�#�Nm�@=�f�nYM޲����@h�&�bNM ���l�`�`�� ��}�*n�� Zlj
�MZ��^�r��voVp;��wPݶw�0�Ǔ��=E�-;Y���r����)�6�Og;Pq���t��/��
�V�T���;oU����c.Ñ��Bfΐ��F�q�@e.ƙ��k�ր�������:ڣ-g�r�z��y=��g3�����9{�+��l+�s�k��칮݇[���Z]g��6�;��=�m�I8�����Oñ�?0�^���Ĺ���'h�Ωڶx:�6l�\�\�@�[�����*^ �_ݷ���t��e4��@=�f�{;�Cu��B"h��=�w4��@=�f�m%4��kpx���������ֽ�Jh������Ӏ�Ƞ�rM ������=z�h�f���R$� ɒDɠ[b�@�빠��޶hL�;o���"v@}[��sI��[`��[�e����n�{��ʜ�)5T5�Ԏ�Ӊ����s@/[4���-�U�{�)VE�#��� �l߿����"a(N")(�-� n���=��h��;�FУ�(ؓ�@����U�z���^�h�J�M<l�6%�rf�U�z���^�4��� �;�$�x8������빠���n�U��9̀�%��׍�;NGBH�gm��k+���pk�Y���$��{VU�<m��n�m�;��>��h^+�;���=ܢ��Ӏ�Ƞ�nM�����zu��{��=�r)#��	ۓ4/GX�x���B	("D�"��E5d�h��/���?{����+�%!I��FG�^�s@/u��w4_*��JU�D�$�DG3@/u�������:y�Xm��6|�ҕA%���SK��v���S�@�U��=�5l<�Ӈ�f�Vs2H�IHA)&�m����z��h�@���h�x�$l16���ʽ�w4�Y�[n�}��ƒn�jDN8ށm��}�h۹�Z���u���F��WDLݬ ~�xm���uX� Q��+#(�s~�I?��'�[p$pq7&�m����z��h׬�/�:����#i&�YUh��#lآ�a�{U���N��r\�7S�h;\	��	��4��z��h׬�-�s@��%��a'� �N7�[n�}�f�m������ď�R��E�"N(�� ���h�f�κ}U�wwb�?I�CWvU�)̉@�M�)�z���-�s@;��ަU���F��՝k m�X�n�ݳ jC�bY ��(�K�Z^����a�ڕ�FCi.�nMJ�K�>ܼq�����,��X+��y7�ؠ���0N�p<ԝL0tn%�6�P�<���փ�N�;v�;F�=���)��ގ:5[#$ɋI1�Es�Wu[��vs��>1َ�ޖ�;�b�t��/C�x�n(�bv7Xm��)�\헶��[c�G|��M�Q���y�ܕd,�UU��q-HD�,��˛6)76�O�τ�����X��r�5��U�����b���vyg��46g�wv, �7x�l�<�e���u� �@!�%&h�l�/YM��@�n���1R�	�c�94�S@�|��/[����@��[�q��54Wʽ��� ������;ݒ�"�L$��r&��;���z٠z�M��@�����m��]u7��dp��k��f�V�ng��Ps`���-�<��F��ۇnf�{����h�����ϐ[nh��/�pkȔ	$�>�,�ѱiY ��RE�d�[J�)�R(��
u�� ��x���?z�VkI�MƖ	b���z���^�4�ڴ��i%c�4#"pq�oY�}�ՠZί@k�M����������Z���w]���O� ���p��9����ʷ	#\������K�GZ��%���\�[j�����o�����Y��oY�vz�]Cl�8�E"�-gW�{��h�f��;V��\��!���D8�{�a�������!p�!�$�$PHE0�)��������>^ί@��P�27l18D�h�f��;V�Uί@�u��9��<�o&F�ԓ@���@��W�{��h�f����a���H�SQ`ۅ��V�b4k�6N[e!yƹ��u6���c)�y'l(Ʋ4ƙ$Ĥ_�~���oY�}Ϫ�������#��Lq�{��[�hy�Z����Ek\m23�G3@-�4����uz�빠w2ǌn`�Gv����"}��p�O� ��x�*hA�]����oN�o쐩V�n��D��-��h{��[�hy�[����o�;؞�87�U!�q�rН�-���t�ݵ���=u�d:��Y�9�ɍ�@��w4޳@�Ϫ���ٟ �N��=�3g����E5auk n�P�Om>��u�~��YД��+�~�8co&A�ӓ@���[�S@���h���U����$UUf(��]�`}ذ�� �즀{;*IX�1���)�s@����ww_��\X�^�Д$�U��U��"�����W�@U]�
���W� ��TIP�T!BAP���U�B*0T"�B)B0EB�P�P�U�T#B0T$�E dB�T$AP�DT!E�T$AP�	BDX�T$@T AP�B�T"�P�B�EB(AP��"AP��B�T 	P�B
T �P�EB
�P���P��T $EB
@T P��EB �T �P�$B"�*�P�,B 0��P�!P�P��P��X����DU��U�tW�U� *�AW��@U_�AU�U�tW�@U_�@U_�W���e5��@�pX �� �s2}p7�@ �QT�B��     @  UR    *٣�  �(�(�"��"T�*  H(   *� ��� (��* $	T(@I	�  @�
��
  n�:w�����R�`2�s��� ;�oYW�þ�U�x�A�PP`;;���>&{�U@���d�������#��Ll��!����{�G��1��o6�k��&���!� _� (�  �l]g��[�8��}���/�
Q΃'�+�b�`���
tpz��;��;�!�}��w���uI���m+���>������n�\�/���n�k����@�� R��T   �� �^�r|��c@�  �l�N �P"4 14i�f� �6S@���Ҕ� �H٠[Pi�6R�@9P��#AM4�4͔
)��� �6)F&�6i�� 4R� ���  � t��)JY`�<��9u�� �2ްrk���ڔ������经��L��zxغqƗx L��ƞ��0o�q� ��gB�42�r� >� $R@  ��qAZ|����oa�����>�z�� p�&�->�.�[��@>�OA���(��p��>���"�7a�}�]�d����3�!��t��p    ��B6��   �M	%*   "x�T�%=@  ��R�y)P  "����ڪJ����d�a!M�*#FA����{����_����M�ggs���{���TAUz��eDWH�����
��EDW��UX�
*�������Ɔ�L��`Ƭ)�5q���.�ن�Wl��k���m"�� �J�:wJa+�����7b���)6@�h�
�X` i�����Y�P�\�D믃]˿
����Yw�{�^�{�O�����m�gg���U�d�پ�|�=��y��*b���;2�]��6�}-w���U��wk�ӗ��Gc��~�+
��`�C�m'�Nͻ�3gm�=�͘�4R��B�L�KR��"���K�h���"pt�hc:M��p4����ٳXP�p"!LtV՗XJ���P�a�[��t�*utɐ���+k
˕�Kl�ZG�Щ�A�'�f��	*ud0�"OU�a�@�p��<ݬ(FU�/�%шv8�cw{7:��f�D�[�����6���kzu�g���B0��,�O+�7�)�|M]��o���	��{]s�w�]x�5�<ay�ɣM���C>��1�^�}'��R,�i�8	J��J��v-�T:�A��$�P��
�X�CNe���JNά�F���Xɛ�{��RW�k�:�<�¤�t�Y0�I�C.T�*5$S����6�j��iӰ�	�d��FHw�l���ngׅ�&z37���9/q��7���,�.���dͫ3�J��@�l[�	�8꺬e���ޯg_.|P�+;_��=��T���6u9�>�]a1��]r�w=�����O�����=30�e��e atA6@� ����J��Vi��N|�Um���nwz�s:ey�v�٥�����:�R*���
4��(L�0�T��i�"|Ɓ�$�032.��E0��N[��lk��	*tH�E����#H� ĊT6�t�.k[��~Ԏ����=��ϭ8���-��R���"ϰ���W��>�yYt�YfUwg����x�pf��M~�2�w;�N����%%�g����<�X
�jfm��wo�0����R��^�����!��:�4�P�	ՙ.#i��dm=�{��pm5 ��>���]aW4A�+����w�;T��g��ڡ�	�a3:x����J���������}K�� [Kf{w�'tr���^�i�B��d�JF�up#"�������5M�_k��?�A��$�a*�ћ^@ E*�C.f��> �;~����#WH�0YE��n�5����ji����ei��:�y��d vHvh��g^tv["��nRIi��0���V-֨Mi��4��2�C�I�JN�*��(E#���w@�5�&r@�H�7(!��CW���N�%K`	��O�����VO�t!��a[ӊ2S�0�}3)��6���!����*T��*^��vI�	�~�#osu{�<�{6N�U��LӎL��������vx�R�a�>u�_��K�3�#w�m��0���`ʹ�]]K��$��ݓ��$/y��z��Gv8{��;�Y�nqIۆou'��{�ގ"�*v�%fo�/{��T2Lzq�Hd3x�=��s��f�4�f�}��D;�7�8�$�c�gw_���+��� ���Fr���> t˙j�:��.}�ݡe�(��{vO$mA��o]����QKoٴ_f���|uy"�;�fu��<���{ks*��6���g�i�����P��ziz#�eT��w$�����!BwR{j�<���{�㺼�<J���aZ"�^nf�j(���Hyu��gBf�}���⳸�B�L��{�L��SW����x�.�L�Ry��Ż;Ѐ�\�o'��YC�{����w�������c��kr ���V>��hN�x{�鱔����v�Zܛ�8�n��4ܘ��Hv#�jѼ��T�%c���M��>/��Ǖ��k7�S�����<�+��~����߾�י�w0��Z��N> !܇i�
�d�Y8�}L�=��s�{��B
;�Jr�ܭ�Tp��1U$�����z����{M<
�I1\3N:����B���3 ��۹�v*v���M�#���!�lXMG�3I�H�V�:GUW�����7�׃mChM^��}����6��e��o'z5YB,{���t��G�R+^[�|���Rt1n��p��
�\��O^��f�R�^m9��������U&[y{�,6�5��vEφp�)!Q)*J�*�R�S,u!�����GqY_L�ϔ�6u	��/e��ۜ���g�'����c�4���	؎77����YH8� 䄓��S	w�母�8ZR�"��/x�u�β���XGHl���0� ��PbhH41L`�� ��¡���ZI��`EH@��J� �Q 1,ZE� ��c	b�5�Ac!bP� E"1ȩ"��F+XE��HR A�R#�E���:	E� Ձ`�!F@"D"ł6, ��V-����	C P"0bA��A�T�Q�U�bG"@R#@C ���"P�L�!D"P�A��HF)A� 0Y$dH��# �$�RF E�
ȊD"�b�r"@���-�R1)�E"�$B�XVAb0�Z�����\Mj1R+�*@���@��D*�J���*b�:6h���٠���#�d0ڄ��2�0�C�xu�Q��ѳ��F75�[X���em�^UC,�Ĩ��x�.���~�IL4� �.I1`ā�ڡ��(A
E:.�V�y�/;�J� �8��	� Ci.$�
���I�5�d��38�u��4�UlSF�=�A;#<o���P*j�)�w�:��R�ӧ����-ҩ�]����C*`�3��z��*�kk0�N�ɂ�rM?�o�`d ĩ��)���_�?Sz>>H ��� P�P ���4�5�ݩ<.^�E;�)��;��6�2����Y~\�;&k�&�me�i�/g�I�E���ޭ|OQ�Y/6��Y�]p�d��=]���"_�i	t�g#�4�_�}������S/Ȭ7��C��
_%�wN��mӥh���:�;����8�����T�����u���쵺d��x�'�����oRR�1o�}���R)�ʿ�7������<h�ē�3��-����2����]��ϒ7�N�i+�b���)�y�g�B'�f��{���Rb��k����|�#�VK[W������1�~T���4��C��`����C��;`��f���2.��T�ʝ�v���V�sR����b�]L2]���u	��Ë��
�`4���������VL���vʎ��R�P�Ǥ�]�_EB���%w��#�8Ē����̱.�|YHc�t�/Պ�uGÒ���W_c��<Ͼ�����r;34\��{�_@gҲW�eFA$%MQLE4P��A�ͻ���']��U���fi�;�$�Ȟ��YP�y]D���˘;8���9��1��O�{��T�f�L��z����\���!$�n�n�{�,��jVn��\��]*BCh:��S8-��&�ܸm-�L��#b��)J�s�&���^�aկL���������>�;��!�~����He�M9����9�%�^�c}��KK��Fw��ċ����4�:�:W�|��΍e\�^�I*�B�10���Ə8�aƎv?o���J�:h�m�ݯ��YVL��~2��P��Y�|i�3x��м�~;�Cԫ�T!�
�l����Ŋ�	H��w�>�\$���L�_�����P�`�ۿ�E&X�L��*HT��
�Y\�J�Rv&\yy��΍Y�V��S��ԝ̥U�B��Qqt�# ��:��R�v��T�J����@WK1{]�@ւ�RA{MU��n����:}vS�P	�����p�srC$S2�U�u!2�Ru`��ੲ.�\�*@�����z�;���*�KU�g����F\��E��HÞ�0,������<ܴg]f�#`�������� B
�X:�|i�5�4��+@�\)p����Z�<��ԝ3)�^�U�R+HpqJ�W0�@���'7�y'��� c,D�.���t��;�;ߟww���ߐ   6�                ���         �         ��          �   � �[@     [@6�                                           �  �                         ��                              m       � �|���`���9P�'�  )[���ľ�۱R�۳HM*���E1�(䊶�IN�Ó3�g.�I-ޮWK�:�I�N��e�$M�*��YW���q\�#�V�e�g-s�(�ͰpH��<m��$-�m	���m��gm�j�206#i����:�-�y�i+�Mֶz�a˸��܅�N� ���,-�Vœ�#Z7:{u��Z��"GG�!��c{]i�m��VU۵ƪۧ���z7b� r�.sYVݱ���v�d�s��m nܖ^dW=%��I��Y�m� �V�8���*{ku�;	  p���좶���.���r�L�7l�;lمɵ(�mגej��m�9����,��m��XW-ml�#����bR�*�WH��VÞ�1��b�^p�޺�YT��/-UWl����E�W5,�9���j��S�����V�[ ܖ��]+����:G-���� m���Y�v�{g�m�u�)iv�qE������<�}��^��m� ���;�`N:�S�l���e��.�kEl���M�$�UP�K�n�&q  :���*в�UP*�T�hϑ�n�j�.�*
���sT�W/:^�W�[J�0۱�yz;<���oN�Ի.�{��a&�d���x��4E֯U�[�����k��ceݢ 7m���u�%��))�j�K��%�`|p�4�M�08TV��)�qj����۳��Hm��P@[z�Z<!v]��x#����'-����$ []�I�<ż��Z nխ�F�Sr�"Cmm�$		��n4Rڽm�H^���ybI.�7j��ְ�ņ��ON��Nsd�m��қ����!˶Y����Wqu�;2��P�U�l�i��;c����oV�c`�N���A��@[z�$6���.�q��\T�P
��MT�][�`��� ��I0�u���Λ�Ӕ瀡0�
����Zڦٶ%s^L-�M�����3f���7�$��{4� ���@s�Hݤ�r��tM���!�$�jt*�����m����W�x(
Y�5��� 	  [@ᶶ�  �m�9]��*���3�h
��õu��:k'A��f�2 �Օ����caT��A,UP!(�@� �����l�O=�m�d-ĩ�Zq��\�ض��v����]�Vv�t�`l� �^�@-���    6�  m&� 9��]6  m�       	   �	     ���� -� �    8  	6�-�  &�l�@��$   6�$� m� ��@�  $      �           [@ �`  �,�ֈ��8m����m�m��Y�(ڶ 9�Y�m�cR�c3��WGj���h�PƖ˶ܭUTI�z�k�����nٶ��H��ѭ֓k�6F�y�
��Nm��l 9m�(��h�v  �az�9ݶ�*�q�6�؈��j֒N� 	��׶�d�� ���$�`m��  �  �����m     �� mh ]4�   ��   �`q���   �	l  $ �	 m      �` ��  i � �-��� m� �H   -�  6�m�   hm��:mm  m� lm��[M��        $   �� m� �i��Jm[@km�,0-�  p�   m�    � 	�i�   �l m�[dm��m�  -����H    [d  ~>�����[% Z��� � -�[vضMV�s�Qm!��m��+u�r�4�uOnܯ(��h>����_�������;5�q�,qa�q����U*�9��Uj���M�m��7m�l��K��뮻k)(UU+\m�xnY刚���H�I�*ҭJ6m��֡25&��m�v����  �ێ�����kX~���@� �M�l  8 m���m�    m H $    �[C� l �  � �`   m�� m�[F�8  � �m�  m 8 � 6���@ h  ��6��@ h� r�� W/I�ll�%C�Wm���n�n��P���T;fUR�(յU�	 �iV:�lA�< ���9�Ŵ��6� ��okwu�W����$�Q�UlY{�
�Σ�m��t����Kv�]�m  �$imhm� �c��ubI'�k��c�\��Ŗ\n�궏N�@��' :�lpu��(+ �������r�'�^�V�8�y���oC�1�c�u��ܜ�۲�k���i=cu�m��f������*�qu�J�@�8�Qʮ�K��nu�!;A���[-�;<��v�AU�G|��U����Qս��;3���{5��j��9��QZ����(1��#���CE]f��+�l�e���U�� ֶ3۱g(覌9�T�����t_����6��t=��jU��7l�LŜUU��>����h�ـ���1�������@�/��@5����#W2�p	�vr`U;�ԫ��/ n�i�&���'!�UH����G(��VV�#�d���UZ�4󛭲����۞ڔ3���ۉg�nS8����v놱��n$S\�^�^�����JU6���*kkv�y`�~�on���Ͼ��OX�9�U("�|['X{v��R�	�$6Z���^&�����h<a��C��5qu�QFi&�:�����AY�`u�>V�m��mnBt�3V����5���iy���uKr�#�7�_bEU����SA���%-v��ώ;ts��ɬ�����m���ޮ�;Y/i� �m��Z�/!d��F��UN�vZ��'b�&��$�xҴ�IͶ �����;]M�cu�7,��Wexϖ�Zywj�6��P�vA��:���J�j��-r��*ø���"#Ϫ���Wm\�SS��c+*����r�@F��Egi��(�-	��-��M����7[u�1e��TٺM� [�Y��*���Vq��|���D�NH�e�!oI}J-ۥy�s�5�� Ի*��` .��[r���/A`�idonH�l���U���K� 5Am �c{T�zZ�F���ma:t�nk۰� �[9�l���e�ܐ H�����Fm��(Ӂ"M��m2�7�t�%��rQl�H�lR�$���=[Bۢ�Ѫ��  ɭ�l�)�4�6�t����%K����:�H��v �gI���l ��6������Gmȳm��o����Ձm-�� N��Ye����$LYB�ޟ8�&�̌!4s]j��u��ѻ�!�-�	��ȶ�*&�� �:s�u��3�rJ�6�O��die8n�$9[� 8y-�Mn��h6�݀H�z�i��=a-�jZ�c��@/'	�m���n��J�]^�7}_t�V 	z�Y��m�����坕�l��]��YM&� ij롚廷$1�����U��V*8G���E��$���N4��F���מ�w{8)�x���l��j�hI%;�z���:����t/}*W}��eD�m�d�dX��`��Z��mq��D�.xGf�����]n�S\���t��q�����@�U\덌�l�r�$`6��K&�T�&� n�Ӏ$�(�ItZ�GHGJ��X$�]m[V�$�tI��N�T� ,�p	8�Վ�:p�ci6   ��ݻI�)��η�@ m�l���  8 7m��%���z�M�� 	����n�h��휜;Uu �K�֥.��', k��:��庶�
U�Z�+�@ ���ޭ6�Y`x�s�&/]nmz5-�ٹ��:E��� ZUU��8�����S$��Or�+�o���=d(�0g�9�:�,�����l[@�c��MjB����m�t$���ް�ӫl�yuu� �U�第��%)]v��j浯�ET���: ��¡�@?��xC� � �/D*��"����]q �PO�����JqD �P��Ҙ"�;BB�
�����۠�*P@9���ۥFqAҽ^��D4lz!��Fs`�	��A�����&�~ʠ����"�P:�/¢qz΀E� �Eȃ�� _�M��� 4�#�(t�*�P�(TH�QC�x*q,�4�B(�A8 �4AW���E�����{�>����$�c $X��a"� EE���(G�*s�ϒ�����m`���DS��~E��8�� �Q ��	����'�!�UDWJ?�~b
0�����X!F H�X �)��Ul��R
�_{���zN������   � m� l �ۤx          8    ��     m�Um(���p녧+�V��+m -o���&���v������Lsr97'j�]�<]�1[X�nv�C�m'':��G�G]��e'n�]sڴŶ{�38g<ط�)\�ƻ^�vwV.V�۷.�˛���a�Ŝ';7�u�!�L�v��'Ds�Y"In���F�S�+���b��n�^��j�m�m�3�0X�	�-�����=p���i�"��ԛ�0�Wg��U�q��4����X;x����ܵ́�F�Þ�[��:Ie[d�� ����EJ�P6�
�,�L I�Y �-��`$V���:��a�f`yN]�ڪB���˵��=�=;Cخ%�eM�T$f�m5���n�iV�l*�U*�Բ���VmUr8���l�UUA�*�u����t� ��l[\�h-�����k�Z�����X��n�n���8z��ɶՑ�剶z������ ��T�vUvv�U���첀�*�	�
u֐ -��nŴ.�2���#T�PY�=.��3��,���,nĩ���ѳ��1�\hƹ�V|�$��l���������k�-b�Iݞ��B��YޣS�[gA+۴/��g�9D��x���� X�Gn72�9�x�V75��Ʉ��`5�`���z�J�J8�v�ى�i����/�ˢ�c�S��g�a���䛛n�.��Mb���j5�vnλS%��Li���e�kI�*]���Ÿ�tY��k�*0rx��SZ����l����fe�k�8|��v,/,���x{X�\��Aq�Zz��^�!��>@��z���gu�0�����aWZ�d�=��.F�/eRˑ�BL��8�J�mR���1,p��7i�.G�B����u�B�r��4��V�\�B3{��ߐ_�a8�b��?���>ࢮ��U$���$���w�$�@���I��l����}�u�X*^�GF����+��X��c����]��,�ָ���d�^-�n
��� ����/g�.�@Ƃ^d�ܵ�ꀶ�Y�/����T��i���N��v�����	�%���N�W=�m����H탟�ۍ��W�f�9Tx5�5�uÈ��>�X�;�q8�p㬐�^�M1�2�d�V�D
��$�Md$�r��@������gc�݃˝�ey�ۜoa�5�.��r�"[�}1%�~�^�{�.��zmg��$�i<q�i���-�����z]k�;GeĢ�N#�I"�/[��{�ՠ^v����@���ō:�4�L�=�j�/;V���Š{��h�}c�ȟ��qhs�h�,Z�Ł��b!nn��SDL��(R#a�jT�g���l�7b�s�V燠�]���u<u2ex�x�jA�������c�������v��{*f�m�q܏]�}�:��!�!M�𔴨BJ``2����meDLr3��r*�j������e:V^Y
��)�!#rf�����ֻ6"#��7[J�����0�&⢦e8̓����^���b�=�w4W�h���D�bx���q��J���q`<�e��-�y���j�F�tk���� \gnXc�lo]�,�l�nep4+��V�e!4�U.��ۋ�S,�mXyN��܉3�cN�`F�E&h�S@�e4^�-�w4�c�@A"��1��)�z��io�3���w4�)�{�x�W�9"m�@��b�-�s@��M���./`%����R8��@�n�}e4
��@�e�@��H-�,B��E�� |m��;CJ��c�a�P��/Vny�=�z�9�t �'�BI$���h[^����m��,�:�LbQrVנu�Š[n�}e4�2�0S$�0n=��-޻����*�^�؏u�F�6���`7���~t���l69̈�AD!�d �
������I��B�ǉ�<xF�L�/���U���9Vx�,���A2���	W&���5����KWg2����ƷV=�������<d�냗����$x�s�(������=�+Z�w4�j�>�F�<U��5�HǠ[ek@���|�ZW��..K�5q�RH�k@���|�ZW��-���{�d+b�dI��$�L�/��@��z�V�z�h���R����)�U��������ۋ�76s��|�$QD���0D�J����]j ����Z@E� H0�w�m�kn��� [A"���*;�ܣ���D�8�rr4�Wb��Y5��"Z���˜q�M�o=n�Ku˵�Ӊ�e�,��jΊ6Zj6���6nY"D4H[H�K\��V�K	ڛ%����7\��q�L�Y�8��a;��Ym��������b����n�ح��k����Sm�c��6�j.�D�(v�=���khKFx�xC+�N�3����n�,�#U�5�On:w��ޛx6�X۝�l���<����J��\(LJ���<��e���z+�w^nl�9�2��C�o �z�o�31#�w�̀n���+�$��	uDR�s4
�k�z��Z�w4�c�<H���29�[�hϮ-޻�}�hu"m㤘�&
I�_>��z�h{���f�WbAn0�"S!%	�#��F�
��Jc/V�3�o$���m\�<�����`�) ��׮�_u�׬�Ȏ�Տbl֢��
�T��EUUUE����u���A$RA`@B�DDr��D�"(	v��k1����X��	��	�@�rh^�@����w4��h�2�Ȥm�r�$Jj�7��Nq�M���ŀu� ��h�`�o!#Q��1�y�X�D/k��׵`b�8���,��tgv��3����e�Vq��E�r<��9�K�[�<�2]nWT�ض�4���^�@:��/uǠu빠\���(ԌL��h^��Ǳ6׷׎��)L�K*�b+�Ӓ�%����I{��LC�
(�l�<�W�yx1.ˌƅ��4���������{����q
�(B��#�f�{����z�n���빠}�:�%$�J~i��:���9�jD���'E�y4햹My�9é-��X��'#��LDD�@�^�@���h�[4�ea�H�,��R����n��9���ŀfnՁ�^�g�H����m<���7��4�n,�n���ly��B擩�a�j'3@=�f��^����ܛ��$D���c�@ B�R�X$R��� P��~6u�٠\�:��&845�H��>W��=�t4�[4Z ??-h��]cS8��jM������A��v��fą�Dz�g���*��m�15=3v����q`yy��:�s`w�Tˌƅ��4���fbF,ݛ�wf�����<̥H*(���$NL�<�k�>Vנ{��h�w4T���Ǌ~P�z���{��@�빠yzנ�VnA�9I8�{��@�빠yzנ|��@_���':��PxܒI$�[B@�.K��ݺDs�i�M&�Ntwm�k�y�����������&=��ݍ�.�7�i���*�ږ#����� �R�tR�/Acb�A�yA�q7���Ֆwt��÷ rvq�v�:��Ռv�����z(u]�ۮl%�6E�p��&�\di����o[�h���Z�$뛱�4Wm��%�����������{����76��ٹ�z�<U�F�
�gq(=��g�N��.��8���K#i�jH�S�<��s@���@�[^��u�hv34�ג5�A�9���Zyڴ{��@�빠\�,e(I�G#�@�;V��u�h�w4/Z���n�$m2`ԉ���t�h�w4/Z��hy�U�\Ōx�RAh�w4���3+ut���z[�`w1���J���2�^N!^���;�qV�V�/�f�0�zy��\��5�DE�TNo9�����ߺ��h����s@��c�Mi��[�7$��w�nȱX0H�����TtP�z���K�빠{��h��a�4�m���;��+�Ł�n���Kj��!�X�x������@�빠w[��w��@�v��>�3i:�k�B�4�w4�j�=]��[w4�w�ߏ��?�n�]���v�x�U�%��t��S�LE�)؇�/%v���w[$�k ә����z�qh��h��h�U���ɑ)N-շ
���s��Fn�ŀ��Ł�-��H�(�;53ʘ*�f�X�n,������mHF�Y���v������ )r���Z&	�;IV4%V��B�
*ƄK���Q�VT1�h���fˣk)1�mV�r�4Fiy�ኄ�:}�*�;;��˔hc�H�	�eIu�!3�k�l3{H�0.S�R��e���\�*�R	YB�%RT$HV3T�F!Rx�wQ�'��5�\4��K����$����e�F��d���0���%Yq��qH[�9�M�aR!F]1���
�B��*���(�-HVRR4%�
4+
�(J�hB�H0�(�ұ� ���B�xB��?~�.�3�.i(R�.�����,�\I�S�0���S4ʐ�*��)�
$	�L1ĥ+2�*B�(ʐ�
��*ʲ���(}��p	�:�R	K���@�i�ŝE:�'���Qڨ9��*���D8 "����*�E��ϳ�]�;��ŠZq�)��L�G&h��h�mX�J�yŏw�`58�N���&��˭z�e�@�[��f7q`lr#��A=)A��TL�L��ОX,;Gn�ݳ�X��ۣ	�WY4I�,#��ۋ�=���-�n����˭z؏+Zm�H�p�H�cwy����1ӥ{��"=�$-�\[SRP��T�X7n,�u��X�w]��c?�$�k ���|�נw;c�=�w47ه�D�Ґ� ! $aa	�3b�s@�����a�n=�ڴgu��=m��>]��{�����N�&ud-��"�}	�6�n��7[��d.��x+��`��bsAk]�M1��w4[w4�Z��j�-3�+�q~S���f��n���^���Z����V	%�o��h.���ՠ{��h�����h�9,�Q���/;V��빠^�s@�u�@��+Zly"��$��h�w��,�nl�ڰs�\�F0�Y�$"�8V�H�1a	 a) @#"DH )�) �$Da�HX)�;��u�jۭM�� ��@�Y����7Y���b��2]��x�`m�>���9c/p�e1�fɹy�6�ϷgV��!�۵�82�W��N���h▧P�`�B���Ck�4��y%Ebw��ti �<�=�/��7�Ʊrۋ<��pv(,�[��O2�;;�v8��[���T_[�8���s��+�z��}���a��G#������1�Ȕ�$���m8ݲ�Fɠ�* [����2NٵC��,�ƣR�P1��6A~QG2�����˭z�ՠ{��h�3�?!�D����h.����@�u��:���:��rF)!0qǠu}V��빠u빠|�נ}Z�Z�	pI����=�w4�w4�Z����-3�+�q~S��ܒf�׮��v���RIwu�>�$����{�6t�mX��R����̇0�E��k0իv�[��66:�ų�5����z�X��+I%����"9�zR[�~�o���??rA������r���p�K3c�I/:v�I%�M����_؆��li��p�LZ�J���w�$�;�i$��ޤ�t��K��k�b��̒L�䒵�ũ$���ޤ�t��K3c�I,�FT�QEF����-I%����I+e�jI.�_��J�w��^�V6�150��I��ƕ<�'�٥�� �e�-l�i����gm�&�����1�� ~~_����>�z�M7q6�K����$���;���L�G�$��~ϾI"۹5$��u_|�V˨ԒV�ڊ�_�2dwrCu���}���{���u�@]A	E@ww�����������}�HoR8�( �ɩ!}gU��%k��RIw���|�J۰ԒK�]F�D�()#S34�Ԓn]´�[ȎCǾ�y$����K�:��I.]�diș�Ȉ�a{r`����a�Dȶ;���c���TF�t�ٻ�������89	&-I%���}�I+n�RI}gU��%k��RI}�c@�,Jdc�g�$���5$�}���IZ��ԒW���|�]�Ό�\��4�D���I�c]�I7.�ZI'�}��$�wa�$��sU�A�$XԍH��$��p�$��>�z�I�tZJ�<��r_�*����+��#1(�G#��$��>�z�I�-$��c]�I<�p�$��~��߿�sc�U�vϭ�Gi�xj�a�gq]�[g�J�I[6}���N��wOp�X:dm�3�I%���J�u_|�W��Z�J�����%喠�m
I�HI�jI.�ƻԒ̗p�$�6��I/7tZI%ܺ��$��$�bN/�I.�w����c�[2�v贒Okuw�%���i4&E��HG1jI.�~ϾI/;u��K�Z��$���Z�K듖4c����DT�Gz�^��KI%��C��^�IZ�����������;�m�պ��`m���^��/\�re��r���(Z��ܯ&�O�g�����7j�m�\ !G;��L�ZPN@5sLp��lI�˵� V��к�R܂�vv����2>ysp�-;��W�[��\�3�g����Xl��:�an��x�����ܶ���:mV�[�ç�H4ܽcB�B���>���<Ƌ�Wn�B+�*���y�һ�.>��f�m��2U���*d�1ns�_���=�dy�7]�u]=n�{]j�XY��߫�]�IfS�ZI,���#ޔ�s�
��ͯ����O$E ?����/��#�T�����RKv��ZI'�mw���~~���܉�M7 �������e;E��3:�uw�%�;p�$��p��tQĢb�T�Gz���{�ZI-��]�Iy˸V�؈����ޤ�-�s(�Ȧ1)$��J�Z��$�]�Z�J�_��K�]F������i�!1I�ˎ�Q�tt��K��6c���Z7p���gD�6����*C?�����$�y��ޤ�e;E��~��z�^�J�m�WdiH܊\6����M�AZERA�P���B�B�R4�	a@B HЄX"� �#L�cb��� �����W��7f���w�������m��'�mZ�;�V�7[o��bX�Iϛ��}�G"fq��+I%��c�I,�gF~.BD�@n���ֿ�I/s��RI^��}�I{��jI+���I)-���\���}�����PW�}���I,{v�Iϱ�z�X�,p�RP�ǌ�񧣲'�"�m)�q�ש��N���c:����nq��uʓ�8�M����;Ԓ�;���N}�{Ԓ�K�V�K�#�;V��RVY%��n��{�ĳ�Qw)l���RK�´�O���Iy��Q#���I�$I%_���I.�w��Vw�{�7[o��1,m������$������K��ũ$����|�^�t5$�~���$��ˍ�� �)
��i$���;Ԓ�wai$����%���Ԓ^�\�q����~�"�ǻHM�t�J�<k��Y_g���2��p�7Aѝ�Ȥ��q�������$���K��ũ$���>�$���������I'��I,�w
�I?7��RK����ĂF(�29'�$�d��i$����I/7v�I<�]�I^hYw"j<mȖ7#��$���}�J��w�7m��ﻮrۂ*�
"/���^QAXd�����}�=����:J�����%�wCRI+�g�$�s��RI_]��$�����$��n,x�,T������.fHF典	ޢc�J�3t�B�I"�M) jI%{����wqjI+�������$�����q�NO�I.�w����O�I/Yu�I^�>�$�Z4ܒ$�H��s��~v��$���-$�y��Ԓ̚bԒ]��rLRI��rC�K�]E��O1�z�Y�LV�I��;ԒȒ23�)����I$�u�|�]�Qcm����n��}>Ʊ��6�EB���CgFvg�~ ���YBP%XЖT��%%e%%%�La�m�$�$� 3{�$��R��j�4JQ�B0��0e����p0e���ؕbC:g~�5w�_�I��}\�D�*@�1ުc�f�]ِ�d��ڱ�)�I�T�+
���� ��2��73$C�Sۤ�JB�����Z�D�������悳8La��$��XkF@��0�*�$E�ʉ�� �,Hc� ��B$�"���B0d�$(B�+[R����`kDL!���d&�g�Ѿ���� Xi��eJVL��������b�T֬�HŀQ��	H��FB$9KS|�7:~
M�j8�*x+~��������6�  h -� m� kn�� 8           !�         m��Ke��ϰ4NX��0�ћ����E���m�֒s���ײ�P����t���%m��D�N���9�';�>NNe�-�J�j�gٳ۱����9؎�.�y.�ݤ9ιj��&�'M��8ΞջSP��qm�l�&$.j���ۖv��!�Gq[��6�s�:^]�k��ϰ������[
f�E�[y���)��T-��b��{��t:Dv�۪K�3�T�m�����.����x�<g_]}Ԇ�A�<�G\�KUU�9����*�`%P)P��Wf��`$ A^2P@��m�p�/���W>�۷�D�hK�;D�������m�G!�޺U��a��P�m���U@*��
��aI������[*���jڪ�[h
T�keZ���I^	g-�#�� ��v� *e����Uk�%C;kt��s��%m�7:�@/(�[�X��E���Ӯ���bUiV��D��R����i�
x�@T�
�յuSk�n:�7;z+ m�����dHWhQ8�G8��r8�����{]F�ٵ˻vِ:��0������յ���Kmv;sa,�c���ݹwl��Ps�,�1�4�P�x�7[k���C=��qoN�����u�p��9-�,��<m�;Wq�76SC�����v�b��<�S�?�?vT�'[���jE;�n��<(7d ѝY6�8���S��Cч�^�.�g�a�k0a��B���P�g��#��;/\�d�Xm�:u]u���jc�X��0�\u۝�� @����*;��ŀ��[pݧb7N���mۨ�G�*��6�W�髤V`�-ؽ�ezܫ�޳�Y��3�NAi7&Ds�
޵�n�N���ꅕ��V�g�iYt�m]�)�I�9)�a�s[�N�/f�V�G$r����]q�W6�<4����{���w~�f"��T@�W�>>O�l��o6�EM&��� e�:ʋ�l����+vK9
�`��n��vح�݌�A�ێ�H75��:�v� ��G�+�U��2,m97V��9R�hZ�(Jniiٜ��UQ���66r��Z[�x�3[���wq��u�û=�����_3��//8n`3��ڠתx�%ג��:�,�6��%�^�3���������|�X{YR��K.��!�ZQ8���W��i^V��-�(�ڭ�m�̐56o�4�'���v�,W�%�v���#:\��*����9���o-��IyӴZI'/��I^hYu�xܑ,nI�$���$���I%]���$���Ԓ^�N,��&L�����$�]����u]�����#�3�kEi$�]�ޤ���ƞ
I�pBmI!�$��W�$��QjI+{i��$��I$����I$�B����z�M�1ZI/�ݷ��I%���ԒVΫ�KϲP�!6Ls�y��m1��:veMF㴡�k�b睬��t���K�m�����Lq��<����_����I$ۺ-$�u�o�)-٭��q8�	����q��-��}�E�uT#UROi��RK6kEi$�y��~�r#�6�8}�U%!D�SU`?�~VyL�a#ۻV���F�M(�P*�U4����uޖ�V �:���DK�ߦ�{�_%I\Jj�$�M�n��B�{]{6yL�;����5R�w/g��j��2�T��f]�T�ؖ��BͶ]u��o�{�u�����&���W@7^Ձ���o)�r"#��#�o�U��o֢Q(�PMT!L����1��8���K �ݫ ~n��������r"2D�F	Ǡ[���@;��=��`�r.�{ڰ�ٰ�9j�dR�*h�Q5TX}Ϣg_�U�7��`y>�B�\^�\�q��@>�p�{���YM��z�ʶg��\�r��Û������)B��m��]lS4Ƕ{n�u-l=��u�rK�F������h�k�wY�\�}pP���j2H���h�k�wY�y^�@����9�r�G��z��4+��w]��c�$I�h�#�@>�@�^�sﻳrd!�`��!&QAJ��~���Ė��`�.ԌRA	������n��ֽ ����j�$G �H�L�H�،/N�"5�m��Y�Cm���v�ь�S�3V[�0����>���/Z���4+��櫪a2(���Rf��ֽ�g#���1�X����w��'4bNF𙄑���h�W�}�w4W��;�]@�N(4cq��W�}�w4���<���(>�,��x�d��z�������|.{6S�6s��d�IUU$��3T [A �6�h�����g���s�Oq0k϶�&m�%�Gb��C��_[�u�*��CGlql��cjZq7�7&N�UU��h���Bd��Z{���v8�p��k]V���ki�J��>Ml�s/E��k6rt�';G\M�5�Ƌ{ Ƿ�3�����v��k��Q<��j�v�vKdN�s�ݴ��I�,<��#Wo��}_2�N�f ��U)��L��)�+�ВQ֋�d�V�f�m)�h�I�H�Q�x�?���^��_��~�� �O�@�c��F��m$m�X^�7��$ykٰ=�ZX�L�=�u591
&�z����e4��<���ܭ��@X)0����e4�Jh^������:�d�H)&F����Қ��� ��4^��9w'dԑ���ۋv�o<<rm�F��l
ZwY.�OIrd�v%'8��HУ�X�o	�ܙ�r��@>�f��YM��s@�����ⅴZwr�$��}2� P(K���Č�w����G60%�T�TTL���h����;�S@���@/u��u�Oɨ�ۆ�|�Z��� y��5fn�,�%����UJ
�R-�ֽ ��h���/��v���l~~A��JN떉ge{(����L��ӷJ�+��ř.����ܵ[<�,L�{��=�)�_;V���� ��*s"��DRM�n�|�Z���Y�{<��A��Xܙ�_;V���^���;1~�r9 ۺ�31�X�(N�J*�(*"UR�<����u`{��Xo#�r�U���ݝ�D)U4R"E3S`1Ձ�[��_;V���^�z�X�p��a6ND�qXѶ^KcC@���4��z�ʅ����$���ruvh������hzנyzנ���ʭ�G�����h޶h�@��S@�1�U�H�L��G�z٠���}V�W�z޷F�M�`��Q�$�*�@����W��J�=YE��ى%�3�V���) �R=�e4
�k�^�@/u����{��?�χ��F�u����y�c*�{H�gm�N��sW�uΘ��N����d��,q��?�= ��4�Y�w��@�^撲	c��S�q��Y�����ZWν�2��nN=����h_:�׬�/�}SrI�ɎH��@�;V��uנy^�@��^��9]pNaL�jE�w�u��Y�r�@�;V�3��ٟ��:�ے$��� -����]���S��:�u�6ѺX儻q����9��:���a�en�g��nF���׉#(pUn��6��m��k�ŷP7I/E1�kG&HU��-�[[���S��UZ���b9B�)��VRE�.�t��ϙ�cM�㗯��:w-��t+H�]�id��o]s�n�6��tkvw��p�n�P�qB�q�
����Ҙ����]R����펹��MK��9���G83�:�#n6�ܜ�[��.�y�I��,��m����4]���j�;�Z��n�6���I�(ܒh]���j�;�Z�׬���l�G���(��@���@�5k�u�@��@.r��9�&H��b�h�z�h]�l>�qc��`8X�%�EJaW*�8��l�<���=�ՠw���߿?��3�8��h�[��(�Iq���k���݉�np]���z�MɄ�"2&�������=�ՠw����٠{�>���A�rE$z�ڵ`��|ĉ$���`Q��סy7�}�7$�w���<���>���������jנ�@��@���@�1�T)$M����{��˺��v��;V���\i4I )�$�<���>�j�;õh]�����V���� �����VYe��m�G:{�,���k<�4ĜI�`힛�*��-�<Kj���s��Pbof�?���q�L��1�ґh�ڴs�.���ڴ��i+?Œ~�n-���˺�g>�!�~��"@��� F���,�LJС�0-��03	���
Z��B��K�!�:@�K����@�D�R�L��!\�M���Ki)q��q]��#��ϸCe�^/`� �*�A����;@*)�\Sk��Db����~B�:�����i��?����˹'L�n�Xްx��� �qh]��s�h�ڴs�~��&�rH9���T�䶬�j��N5`fN5`o??��c��΀N��X�1�\nM���S;i���c��������v5'��g�K19�jE�����s�Ϫ�>�j�=L}�
Gl�1�$�h��hϪ�>�j�:��hWkh�LS$(�4��hs�������-���@>��Z+�<�b��hs��v�Қ*�U�<��ț�j1��qhz�4��4��hs������ n4�Ȇtu�&qݤ&�ѩ�W�j���k"��vt�3�#iI#Pǎ~����4�j�>�j�:۰�9�X<I�dd�1I��hy�Z[v�빠_�v��7#��r7$z�}V�ͻ��Ȅ��X�vl�'eT�MMUH���SJ��G9���;��z������ֽ�;V��c�I2$�5 ������XDDr9����|9��`>}qh�W��L���F�m$�7$��	 m���:{k6��s�:��[����qY���G3Xq�����[@��nvܗ����}�.�t��t��5����
P��Ԏ��Ii�īi���VyM��<��q,���n,u]���Xv��:^:�<S6����uI�k)���8=�^׆q���$�ϭN!��Ӯ�ۙݱ�@�ɮ<��oL��)D.!/��(�(��r��I�ʺMr;8�vj��u�^X���О�%OEs\��_8J��箎&��������/Z��X�z�� ����!@UD�M%U6�77���kiX�o4
�k����_��8�#IF��Zݭ�`{��y	j�ٰ1��2��dnF����Z����Z�d��6!=��V���*`RUT�\��TXy��7������m+1���j��"M����!n�g���|�bK[n��ݎgL�TtJ���g��zk�0�	��������n�+1���:��w���?�W��7$r6'0�h�M�~r",��L}�������6ɵh�>ʔ�"O�QG������uf�-s����f�~��R��)%�T�XdlL����uX�X�\W��4�5��HELs�@��ZWν�����hvu
�m�r��h�z賢�TՌK��g���U����yG�6���|_Dh�M��t�s�`<n��<���5��7V�?�G#ǎ~��=�����X%�`79.ox����E"f(�����U����2��9|#�"@p�����"HT@0U�뛳s�`fn�X�1ʀ�*�Ī�����L�NK���,7�fnՁ���6Aɑ����m�@��נfv��:��Vc�X�ss1R����$L��6�ma6�y��I���ݧ���݊��w6�	���A7�Ǡz۹`�u`f:g��"9zC흟�����"jHKLj��zٿى���+_��=m��ysWQD�LsMUX�ڰ̗VjX�n,3v��˝Q�IQ�C�;_��>ｳrO��{���X�2�"��Ō1��A� �0#B0c�!�?}���I�z��ؔ� 9�%�������������Z]�����=� �Lz�݃��4e������2�d�kp�;v��R�]�����n�[Sw�m�����}�ՠU���=�w4�wV��S
bUUT�M�ܖ��57;V7�}-��#�Dɟ�誕5*�D�B)M+V��V�Ł�Kj��Kj�y+�I$m�bn7#�C�����}���j�;�ڰ�D'-�Ձ�/y*jd$J&*%T��X�����[��4��X�}�$�WUT�U ����]���+Kc��� 6�r^��vۤ�OcEcM��C��]gq����G6볧�,s��fݭ�q��r{m>%ٶ��\2��l�ݧk�IU��J�Wn0�K�X�RQJ���U��5���(�l6Bx��n`��nn�8�h�������s���z�������x�1�<[����y��.�;E� �bYg��]פs�I{�Ӂp^�����Ym+���K�G/v�e�9��І汵�a�`��G�gs�Fz���g�w{_?2ٗj���ͷ�����˹٠{�w4��Z��Υ"R!*�`T����9.o��s��D���q`c��V}-���,�S�S53JQ�	�@�ۚ����;V��U�y��(!�	�s4?�31y��6�wU��'��r9Ř��`gzH	Ģo�rG�}��h�}V����hW�h�u��8����x��oh���l4Ͷ�vJ�$[�Q;�k��9�1�����ѫt����"�|�w�h{�Ł�8��9��z�r�{L�w)����%��ͪT�ڿ��x���j����W��D$k��!UrhJ&&5s4/�������Ϫ�>�Jh�nDb��Ɣ�C��fb�G��q��X�S,6"8���XCNu*�S@�I0*UJ����V�ȏc�>���-�>�@򼝓#NE�	1��ݻN��sN�mN�m���:}��U�B�,S��T�2ݗy-7$.DB]ǩ.����:��;�Ƭ�N5`u�5<��*
�	����2��H�K�`dd�V}����3�7TL
iT�Q*�UTZK���x���<N�� � �	P�$�HF
��Bg��]��s�u�@��]�D8!� �=�߿.ΗU��u���:e���G���vTr4���7'"�>��?ٙ����|���@�yڴ
��/Ѭ0��fX
ZE����&Z%�^��ڻQ���N�_�]�v�I�!n;�jK��?-��^��)�}�)��ݎ6�+�T*���,��W�9ϣ�#����;�����h������@�*l3)�s)�lr!-ͭ,&�lK������-�d�)qb_��}����76���:�\�"���G/̪f��?{�������/�����>�9��������;��,4*�KFM���v�-�$�u,OYq�t����W4nnw�Cͷ��;)��Mo��u`c2�`w1�o"9Πݗ����[p)�h����PMUX̦_��r""d�߮,���Xq���H͕į�X��NHI���nh��O�~ȈH�ݫ�/U�ܷ	)T�T"b�U)����[��X��X�Ƭ>�r"��� x�v��&f�P�))�`�Ձ��e���V�*m`~&?_�$ͬ$�M$aD�a�C�	�c��7v�%��	D`�@4[(k%e<�fi�^6�N�Y������#RT���:�	�P��)61�t�f<6n4��	I3M	cShPL��v�Uf�滈\<i)m!H��LԖ]7�L�hT�-A�CF��+�"�7�`F�B0!H[.���%��e��2����RR\�ӭ�.f�eR�fr�n�l�ۚ	�L�\cBFH�� }h>VU%���w��O�$m�$� m � �  m���                      -��ۖ.�M�Bt�f������bKέ�ۃ'+v�li�/��ȼ`����n�]�,vħ��Q;=e�X�ujB۫�݋&��st˦���9�Q���cQ�^FR"d^���eA�c���fn���K���{X�+<s�O%�֝Mئ2�l ���z� �v�;��3r�nv�{G[�֑�cca�Í��nKrvd��A^g`��N��t�Hj�j�v��"��j�B�#��n9�i��'L�tM]:m&qf�jB�րUmYM���*�YVUUꭨ�r,��
�r�H�� �[@'c�ې<�r"�[m�j3��-�umJ����H��'�j�n�V��lm-� ��F�[y �i4��@�WQ�dS@G���-��ێ�`�̫OhrdV��
���'�%�V�8j��
YP΄	P�z��v붚z�=�-�n��Vr:���:Ζ$8�m����o$��mG;Ҁ�mK�����ؕ �H�u�$V��]mc��\��۱=��]�I������b�S/Fٶ�X�mn��FݱD�8�����*��6��^ܘ�b.#��
J�':�Ou��U�%q�q9�vw��̚N�7A�h�vǄ�4�m��u���k�d�]A��Km޹Ɏ���z�:��]��BZ7���E�M����������.ݱ�e<v�����`�雙���v�qZ��t!�(�v_ϙ��;t 
p�s�e�]�p�Ƹm�(��\��#i��v�I`$c�8�z��+F��%v��٥��z��x��ۀy������cmpڒ��t���n��rk=����=�c������ݰ
���v�]����]Y��GK���+�
ڻI�C�ӷj[�94l�[�Y�H=�cc�u�A��5��`G��RY�w"!�*|� �l��hU�e z�����~��$���o � Z�]��M/-�ݝ�p��i�v#n�z��k��ۇ���^kv�#[Ͷ���件��u� m�%۰Y]�Y�E�J�l�S��c!h��'b�q��\v��h��@��[v3uۤ��{-���k�nm��۝ֻnv����W&��[�f�pd�st�ۖΝ���%�A��sx9�����#cn��q��;�ˏ�X~�����Дݑۀ�����QLgu��@ݣ7n,`��R�m_��wpd����2C''�Գ��/[�`bx�y�#�{�`l,ML(A�Ry$?H�Z��hW��m�_G���P��}���ۃ�-%.�ůf�1�Rj�ǎ��|^��SJ�J�������s��׵`=�ZX��XlG#���ٰ���SD�0D�	ɠuΔ�:���9^�@:��/bAh2%�?�F��s!�a{r���5�dv���g�kF�����������ĝ�O�AcsH�)����s@�z� ���:�Jh��6��LM�s6I���ͨ�������*�A-���5�'|w^��w�wf��n�&��LS8�޳@�2��s���^�X����Yԭ��Z5�\�!.k[ND�,� dOzs�m9ı,O��p�r%�bX�g���r%�`�X��wٴ�Kı<g׷
Y3<\5���3SiȖ%�b{���"X�%���{�ͧ"X�%���}�ND�,K���ӑ,K�������,�F����7��u�Al������Z*�%�,�Jݎ��RNFv��k4m9ı,O���m9ı,Og���r%�bX��w}v��C�L�bX������Kı?��S���?{���oq���~����ӑ,K�ﻻ��Kı=���ӑ,K��=�fӐDlK��o�K������d�\�m9ı,N�]�ͧ"X�%��w�6��ctD�P$��D��ZD[	��)!R H� uّ5��s6��bX�'�׽v��bX�'��'��5�u���5�՚��r%�`(�'��p�r%�bX�g���r%�bX�����Kı;����9ı,N�^�.��diX�w�2�T5CT5G��߯iȖ%�b�=����Kı;���v��bX�'}�p�r%�bX�����?��5Z7�s�/��\�p *Ԯ7]��c�^�^'v�&��
�Vs(��st��fӑ,K���]�"X�%��w~˴�Kı;����9ı,O���6��bX�%���<f����Y$��ӑ,K�﻿e�r(X�%��w�6��bX�'��}�ND�,K��}v���!�2%��go�Yi3?�Y���V�9ı,O{��ӑ,K����iȖ "X�'}���9ı,O{���ӑ,K��C���Vj�\ц���ND�,�X�{�6��bX�'���ٴ�Kı=��ڻND�,E����$I��6���Dy�����x��{�����_���a���?{��,K��{�ͧ"X�%��w~��r%�bX��}�iȖ%�b~�wٴ�Kı?���$���˫l�tC2�֜����R�	L�=`�(�7k`���ӮLj��u�ċ��NA����r��,K������r%�bX����iȖ%�b~�wٴ�Kı;���iȖP�Q��O���ݻ�G$yF�,K���NC�("�2%��{�6��bX�'����6��bX�'���WiȖ%�b{�z��n�MS,�35�4m9ı,O��}v��bX�'��{6��`��X�'���WiȖ%�bw���"X�%�}����s5�.��5sWiȖ%�b}���iȖ%�b{�ߵv��bX�'{�p�r%�`*�����ӑ,KĽ;ۆ�*���*@�UM�:r�G!��{WiȖ%�bw���"X�%����ӑ,K�����iȖ%�bA~��~m��������UTU�UT�!��������N����.�zp&r�z�Y��˷;�^�Ȼ�׶�G\�f��b����N@ �[3��]-��]��Q
Ù&6��$4��*� �v��
n��쭧S�d�%�g�'m���R��pm�oXxț(/���`vT9[Qk�F�M��:��Q5���H�N����Λn66�u�luq��(4*���4��qZq7wuv��ڀ�qS�IU#�N�_L����ng/u	�����q�E.G�j����=�߷(�Kı?{]��r%�bX����l?� ��&D�,O��o�WiȍP�Q�����.ۉGp�%.�Q��ı=����?��L�b}���ͧ"X�%���o�WiȖ%�b}���NADlK���z��֮K�f�k5v��bX�'�｛ND�,K������K,[��&��!ﳾ�RA$Nw�������KsI�$��z'}��WiȖ%�b}�}ͧ"X�%���]�"X�%��>��iȖ%�w����߼��Ԓ�TT}��oq���b}�}ͧ"X�%�"{�w�iȖ%�bw�w�iȖ%�bw�oڻND��oq�������^���ɜ�bWco�0l�!}e{Z,��9�ͥ��,]�<Iq��SY&j�kiȖ%�bw�w�iȖ%�bw�w�iȖ%�bw�{���*)�&D�,O���ͧ"X�%�~��j[��r�p�F�<�UP�Q��ߞQ�~T���,N���ӑ,K���w�iȖ%�bw�w�iȟ��D2&D�/Oz���[�kMY%˭]�"X�%���sSiȖ%�b~����Kı;����Kı;����Kı:g׶L)s=�u�P�]kSiȖ%�+b~����Kı;����Kı;����Kı;���M�"X�%��!��j�u�sF�IsZ�ND�,K�k��ND�,KD���ӑ,K����56��bX�'�k��ND�,K�ڽ�L��A�^:z*�u�Lvs?��i�ɳ�� �h�9Td�#�t��l��0��3����%�bX���v��bX�'~�����Kı?g��ڂ��bX�'~�ߞQ���j���ߛ��.IW!��]�"X�%�߽�jm9�G"dK����m9ı,Ow^��ND�,K�k��ND� "�"X���'��ڳ*3i��������ow�����Ȗ%�bw�w�iȖ?���Dȝ޻��Kı;���M�"X�P��F~?���(]�r^Q�����k��ND�,K�k��ND�,K�﹩��K����{�6��bX�%ￌ���Y��l�K�V�ӑ,K�����ӑ,K�{����ND�,K��}�ND�,K�k��ND�,K�}��MkVY��GOn�lq�<��-�����mr�ݭ����W��!�\N�.�PP��۸�T5C�bw��56��bX�'���6��bX�'��}v �"X�%�ߵ�]�"5CT5G����b��.]ErE�jKı>�wٴ�?�9"X��׿�ӑ,K��u��v��bX�'}�sSiȊ-�bX�d=ٞ��kR��3Zͧ"X�%���~�ND�,K�k޻ND�,K�w���r%�bX�g���r%�bX�=5�B��%�3Vf�6��bX(bw�{�iȖ%�b}����ND�,K��}�ND�,�K"{�ߦӑ,K����~�̓c4L�}��oq�������j�9ı,@ ���ӑ,K��{�M�"X�%�ߵ�]�"X�{���??_��T�]�致�,�8�3[��'n���uV��9 Ǝɖt�r��ˑ�Q���j���������,K��}v��bX�'~׽v��"X�%����j�9ı,O՟~R�ڷ[�H�T5CT5G�߮ӑ,K�����ӑ,K���ߵv��bX�'���6����Q��{��??��sZ)�8�F>�7�ı=�]�"X�%����j�9ı,O����9ı,Ow]��r%�bX����=���u&�).fjm9İA�w~��r%�bX�}��m9ı,O����9İ?�D����v��bX�'L����d����˨jfkWiȖ%�bw�o�iȖ%�a��UN�o��i�%�bX��׿�ӑ,K���ߵv��bX�'�"���?��a"��` �`�J��nySh�6y�l�ڋ�q���&q]\����tY��c�lw<���$@Dv���#:rN-�Ŝ�: Rv� �i*vIP�]��ۭ���5�#-�.pSgT��T�!��^��d\��]��P�v��O;.�^��p���a����Z'c��%�5n[�ûDm����V� ����^{hX�%iH�R2�b��*��]��Q�:�݅����Nz�����˼=�[��j��[���E�qf��nz�M��D�,K�����r%�bX���z�9ı,O���WbȖ%�bw���"X�%���^�,�kY0�2f�f��ND�,K���]�!�(ș�ｿ�]�"X�%��{��ӑ,K��>��iȊ%�bwݻ�Xf�ˉ��ˍ�yF����������,K��m9ı,O��{6��bX�'�k޻ND�,K��'��UrIwv�\�H�T5CT5G�}�L�bX�%��}�fӑ,K���{�iȖ%��bw�ߵv��bX�'�꯭�-F�ۄ#��F�������ͧ"X�%�����ӑ,K��{�j�9ı,N����Kı>��l� ��jv�|X�tku��n�j�Bnv-��s��*^m��S�{������n�]]k6��bX�'�k޻ND�,K������Kı;���ӑ,K���{�iȖ%�b_��}��k&���)-����Kı;��ڻNC��@����QN{`����'=�p�r%�bX�w^��r%�bX���z�9�D\��,O��d�.�����5.kWiȖ%�b{����Kı>�^��r%��b~����Kı;��=v��bX�'rx�[�#���%.F�����?~yF�K���{�iȖ%�bw��z�9İ?�D������iȖ%�bw�_��ƚS���w�{��7����׽v��bX�����3��?D�,K����"X�%���{�iȖ%��{�����zFG\�u[B�Z���)1m���C�;����v��Y1���{��~7\�.)nEr7q��j��j���/��9ı,N����Kı?}�z�?��&D�,O�����9ı,O�j��I��f������7���{�?=�iȉbX�'��]�"X�%���]�"X�%���y��Kı:wVw/��3Vf�fL�ND�,K����ӑ,K�����ӑ,h����f� ���Rø�)$	BT�!-,���o�ܡ$(���ǅ
E$0aa$��$�3e��,JS&Fcf����.Ḻ8�RB�-Q��6U�mU*���7Ԍ����KɅٴ�A&Q�2@%��L��ld��	C�+j�rȩ��o1������뫅�=���r����a����
�r�����3_�iM@�7�\�H���Ra"0"�$��BBT�Z� Hi!%����԰wz�/%[�%�H[LV�׵i���̅�\!r\��%1�D �шh��"ْ�%�bC@T�HE�F1�,�Oõ��@������*~ @���~O	F�Ev&�8��`(�U? ���� \T|H�������r%�bX���iȖ%�b_���ߦ���8
>�7���{��r'�w��v��bX�'�����r%�bX��}�iȖ%�b~�^��r%�UP��|�1�JAKn��5P�%���y��Kİ������i�%�bX�w_��iȖ%�b{=�fӓ�oq��������H�����Ͷ��c��)�e	�m�ñ��^w$Oi�ڕ�x��2�N�r;%�'wQ���j����ߴ�r%�bX��׽v��bX�'���mS�,K��{���r%�bX��}���w��dJ;�Q���j���Oz�9�9"X��׿�ӑ,K�����]�"X�%���NAĪ���?~C��dj5p�#�5P�P�{��ӑ,K��{�j�9ı,O}�p�r%�bX�}�z�9ı�߾y�.[�Iw"�����j��������Kı=���iȖ%�b}����K��4Q4QD5�=�{��r%�bX�g�==u�֍\��5��ֵv��bX�'���m9ı,O�׽v��bX�'����9ı,N����ӑ,K���������v흭�1�8�� ���>)Ə15q͈e�<7N���N�����I�O�ۖ�Z̹�i�%�bX��ӑ,K��u�]�"X�%������r%�bX�����Kı/��O�ִfk&�[u���Kı=�w�i�!bX�'{�sSiȖ%�b{���ӑ,K���{�iȖ%�b^����I��ZY�5v��bX�'{�sSiȖ%�b{���ӑ,�,O�׽v��bX�'��}v��bX�'{5��%��jG	n'$YF����PP��Ͽ~6��bX�'{����Kı=����K��﹩��Kı=��p��4j���Rk3Fӑ,K���{�iȖ%�a������ı,O{����r%�bX�����r%�b]��;�w~��T;e���Wj��X\k���-ڀ�NN��͞�\����-i�ӝcc�mqq�v�����c�Qٝq.��ָ��jA$�ʱ�B�&�+06�B�Y�Fs��D�Q�t$n�wN�{0pbU�K-�g vV�bٶX��<����#1�ݖ�E�Gm�\�$����x7v;r����-f�A�<�cȗb8:�࡫���]]��Ѳ��[\�ۆ�q��#��ڶVX!���p���,���am�w�u}⛝���֮ӑ,K���w�iȖ%�bw��56��bX�'~��6��bX�'�k��j����;��/�QGi��\n�WiȖ%�bw��56��bX�'~��6��bX�'�k޻ND�,K���]�"(E2&D�;�����S5�j�f]k5�f�6��bX�'���M�"X�%��w~�ND��DdL�����v��bX�'}���M�"X�%���Y��bWpw	.�E�j������g�ӑ,K���w�iȖ%�b}�{��ND�,K���6��bX�%�Z�+��B�-9wQ���j������ӑ,K�O��sSiȖ%�bw�ߦӑ,K�﻿M�"X�%�~��|?��50qt�Q�5������P��8��Pݵ��5��1	9;V����Ӆ��sY��Kı>��M�"X�%���~�ND�,K���6��bX�'����ND�,K��v����Y�%�Ȳ�T5CT5G�O�<�Q�A���&*ؖ%��w~�ND�,K���ͧ"X�%����jm9ı,N���K���I�.kWiȖ%�b{�ߦӑ,K�����iȖ�%����jm9ı,N�]��r#T5CT||�ߪG!q[�;�e�q,K�{�ͧ"X�%����jm9ı,N�]��r%�b�X��w��oq�����~��?�=�3�F>�Ȗ%�b}�{��ND�,K��u����~�bX�'����6��bX�'~׽v��bX�'s��;�2j�X�)v���<�ױ"�e,:[[]h�^�J�Q�G�o.=�Z�!)���������d�=�fӑ,K����M�"X�%�ߵ�]��"X�%����jm9Ī���~�}o�!��K�%��j�����M�"X�%�ߵ�]�"X�%����jm9ı,O���m9S{��7����w���[4��m����X�%�ߵ�]�"X�%����jm9���j&�}��iȖ%�b{�ߦӑ,KĿvI�75u���--˚�ND�,T�{���r%�bX�g���r%�bX�����r%�`  L������9ı,Ozk���˫�WR;�e�j��j�_�^Q���ı=����Kı;����Kı;�{��ND�,K�wܲfk.�6W]ײ����bIq2�g�����=�ؾ�������]����1�7�5u.
%w&m?D�,K�����ND�,K�k޻ND�,K�{���r%�bX�g���T5CT5G��}���qF��p��m9ı,N��z�9Fı,N���ӑ,K��=�fӑ,K�����ӑ?�"�L�b}��w��f��r��f�k2�ӑ,K�����56��bX�'���6��`�ؖ'�׽v��bX�'~׽v��bX�'��x���rG�.Ir,�UP�Q�����5%�bX��^��r%�bX��^��r%�`At�(2+���4~��߿��M�"X�%��wVc�#Hwp���yF�����~��G"X�%�~׽v��bX�'{�sSiȖ%�b}��iȖ%�b~�����][q.�S"H����Jn7]�����۫�֞m95F��l�V���bX�'~׽v��bX�'{�sSiȖ%�b}��b�"X�%�߽�m9ı,K�d��l�jKu--˚�ND�,K�﹩��Kı>�wٴ�Kı>���ӑ,K�����ӑ �Q�I���-���R̗3I�$�}}�fĐI���I�$���^��r%�bX��}�M�"X�P��y����\J�K�5P�X�'�{��r%�bX��^��r%�bX��}�M�"X� �'����ND�,KǦ��kY���k&h��m9ı,O�׽v��bX�'{�sSiȖ%�b}����Kı>���ӑ*���@��@[���ߛrHێ7q� �H �˦���A�,T_JҸ�J�ݡ�t÷!֋�%ۣG\�n�n�q'n��mn��� 
���V�Hu�c!�me7�ی ;���f��E�x��{c�=��)ś%��m�tq*��&��w@�Y:ؓ�k/6#mm�6^`���V`1X7=X��T6л��\�\u\��k[&#�:�Sog+����|����@'w�F�i�!\ܣ����۱��]�6�î�j��{��D��uН�(�����7����{���r%�bX�}��m9ı,O��{6��bX�'����ND�,x�������i����������d�>����Kı>Ͻ��r%�bX�g��m9ı,N���ӐA�,Kǵgr�SD.jLѬ̹�iȖ%�b}�{ٴ�Kı?g���r%��C"dO{����r%�bX�￸m5P�P��~W���$��伣�,K?�H��O�����r%�bX�������Kı;�}�iȖ%�b}�{ٴ�Kı/~�w�)��-Դ�\�m9ı,N����ӑ,K�����"X�%��}�fӑ,K����iȖ%�b{�x�3D�-�c�8��.�Wv)Ͳ���bLf�h6t�&�j��m���
2�c��iZ�!,��QȖ%�bw���ӑ,K��>��iȖ%�b~�wٴ�Kı;��ڻND�,K���Jg��f�Ԛ��iȖ%�b}�{ٴ�>E�ਘ�j%�b}�s�iȖ%�bw�ߵv��bX�'~�m9ı,O����)j�$��j����;����r%�bX��w�]�"X�"��"dOw��6��bX�'s��ٴ�K��߾��d�ܴF��۸�T5C�� Ȟ������Kı=�p�r%�bX�g��m9ı,O��}v���P�������"�%�r<�RX�%�߻�ND�,K�)�����?D�,K��{��9ı,N���6��bX�'��}���e�kZ�D�{=��6��VLN�����֢�K�s�sT��vNɤ�v��J���w�����D��_��iȖ%�b~����Kı:w���r%�bX�����K�j���_�J�I�#v7#�5P�Qb~����D�,K�{�M�"X�%����6��bX�'�k޻ND�,K����%�5�[�im����Kı:w���r%�bX��}�iȖ?��*�
E۵�qB��N�k��iȖ%�b~�ӑ,K��_��=u�24K��ND�,� dO{�ߍ�"X�%������ӑ,K���{�iȖ%�bt�w��Kı;���%.x�\Ժ�k4m9ı,O�׽v��bX�����]��%�bx���6��bX�'{�p߻�����ow�����6:11]eӵaS���dx����6n��,��j���̂��G%����(�CT5CTw���m9ı,N���6��bX�'{�p؇"X�%�����ӑ,K��>^P]le�E������oq�߇{�M�"X�%����6��bX�'�k޻ND�,K���M�" ��-P�_����8K����5P�%��{��ӑ,K���{�iȖ X�'�{~�ND�,K�u�]�"5CT5G����w��.�D�;��Q��ı?{^��r%�bX����m9ı,N��}v��bX]Bj�a�H(���N��p�r%�bX�����q&�$���\YF�����w~�ND�,K�u�]�"X�%�߻�ND�,K���M�"X�%����ߦ�۲�]=��x�xJ�UZN��e]n
�B�E��x�n5�ح��瓣�f�ӑ,K���w�iȖ%�b}�}�iȖ%�b~���yı,O�{~�ND�,K�}|J��]M�&f�ӑ,K�����ӑ,K���o�iȖ%�b~����r%�bX�;���9�,K�Jx�x�\պ�W4m9ı,O���6��bX�'ｿM�"X�%�Ӻ�ӑ,K�����ӑ,K��ٯx՚�Թ��Y��6��bY��"}��M�"X�%������r%�bX�}�p�r%�b�'�{~�ND�,K������"M]�%��YF��������Ȗ%�b}���iȖ%�b~����Kı>����r%�bX�1}��:��&�DC2��)WJ��[��)�,��hW���)>��R�ug��h��+B%����VP%#����T�f�ϒ�CfU4QS��oge�-�T��(AHL!�
�e�����bHf�e���������m   ���� �` m�@�        6�             ���ͮ�mN�H��s�G`Wc�v��*֫�6-�.�n쇮�f������f��E�c��L;�kM�5�H]ȸ_6�+k�l�m�:^%;=�xsL	�k�ED�잇��(�Z�y-:�-TKRU%�Y�7������^�.2�
>8���sg�iIvy]�P��v^W\;sڶ�&��ɼU�M�ܹ4;8�+���֣2�qM9��s\arc[S�ےK��ƺ|�	���Ҭ�`q��X�;�pyd�_!nu���Wi��m��[[N�K$�� AU� sVէ���v�@�e�jڪ�U��j�a捀 ]t�u�h��f" v�GrW�n�)�8��.�=T������j�hsm��8q�����A���	6��[M��V� +�U�%g��y��Z�U�h
���@U�e@���V��\�����g����wa��9����0
�ۉ��;�5sf�Q8إ@�m�V�=��T�UmUJ��Lsm�����\��m�&A&����u�\��*��]�bw��$�������m63���ρ[YC۞}m��7;�a��K	����x՛���G[k��oT'+�R�XVt���*rIXb6�<����W�+et��ۂ9y�ۧ
�s�ˌI�slv��T���A�l�����]N�R�
���Z^;d���$�Sk� �s��Gٝc�=������^�skm��q����6�Q�]���*���E�	ڤ���E	8�\���M�Ũ9X�L�\۱�����9	\�`���N�ۍ�.�
&�h�ȹ(6i5�ku�X���me�c]�����i��q��h�v6	ۛ.�okl�S�e�N�n�]���/kgkr6���^�a}Lplh�2������]�4\��։� ���(2�:mm����1�'V��4�ֵ�p���!�>~t!�A�|+� 0*��/�Q����~��~?M�kn��� [A5UT�!ۭ�ݟ,'=v�S]�Z9��t�N�0��ݵ���Nnz�X�^kضi�Z]��CE�MI� $MF�LNx+WnC`�&�s!!t��2aP��$;m�G&5�cn9[��6����1xB8�=uۺ]g��.N.��w��u��=�Cz;,�����t��0qk��ۜ�sf3����lwGg�;Wc��9���I������{T��5S��dƸ���;Kj e3[�\�b��\� �wS�;��竣�F��f���v%�bX����6��bX�'��~�ND�,KｿM��!�L�bX�=�]�"X�%��j�%˂ĉmȲ�T5CT5G}�?-�"X�%���ߦӑ,K����{6��bX�'���6��X�%�t��n�M��.��5P�P�{��6��bX�'���iȖ%�b}���iȖ%�b~���iȖ%�b_�'�L.k&MX[���ND�,K���ٴ�Kı>�w��Kı?{���K�,N���m9ı,O�������jI�ML�k6��bX�'���6��bX�'}�p�r%�bX�����r%�bX�g}��ӑ,K�w�������l𻮼6Gr�]a)ݚ�4j�n9�VB�B�$�r���|d&jk$�Z��r%�bX����iȖ%�bw�o�iȖ%�b}��{[�B~��,K�����r%�bX��f��#�.�"r�n�j����>����9ߴ�lMD�3;�����bX�'~��6��bX�'}�p�r-�5CTw��l�v[�%�$��<�U%�b~��=��"X�%����M�"X�%��w�6��bX�'~׽v���P�z~�~�ĈI%۹re��,K�k��ND�,K��m9ı,N��z�9ılO��g��䡪��?�_~�.$��$Q�q�ı,O{���Kı;����Kı?g����"X�%����]�������_��{)nEj��a��x�T�2$n�ː��a�|�GD�o.ƴZ��s�7q&��C(�CT5CT}�����Kı/�{٭�"X�%����]�"X�%��{�6��bX�%�O{&d���35m%˚�ND�,K���"X�%����]�"X�%��{�6��bX�'~׽v��bX�'�>�%.\�֤1�r�m9ı,O����9ı,O{���K��������R��E�q9�׾�ND�,K���"X�#Tz���+��Jݸ夝��T5C\�Dn��:��V �qVr9���~V����87Lɍ��yڴ޹4W�h���^�6�2�\�=g9����]�e�U��۪˹�K��4�VLdo���f��<�$�4���_����)�w��@�w��0n6�c�L�̚�Jh�h�j�{W�H��C�UT��*JB�,Y�6zq�>�s�H�zU��u��{"��bX��	��R-��� ���d����ܜ"����3�׹������F�6D`�#�<��zץ4/Z�^��W��diȱ����Aϱ�e�)�(2��N���tk"��mњХC%?L܏��?�Ĥ��Қ������X���4�A*U(�RC@���@��@��Q�^����{��w�˿�������.�g]T��S��<���>�q,ͭ,Y�6^F�����H7��t�h���<���ls�DK���`=��_�L�RUMULԫ�t��ݞ��7f��e9VlA͍����U*�Bf���*����p��y�Y!��z}:�1�l6X�6Ѷd���v�z�Lz���΍�������F�uZo;�X��e�J�Y]����/A&B�RQJ�W.�vn��-��^2�&���%x�m��j���d�]�:+n�Hb��:�n|l6��YsnN k���U��u�c�Z�݇tW��u�ڣ�=��v�wEźR68��[��ջn�xm�o���v��0H���:2�J���օ]�\��x�J��\���չ܆�)4��#"JC�U����^�����ۋ �v
�����	�T�^���빠yzנv[�72D񰟄7����=��z�ֽ�y\m����3"����s@���@�zנ�hG�Q"��N5s4/Z��Z�]�M��s@>�P6���	�5���C@V�Z^8N:e4��62x�s���DȜ�FHLrG�|�נr�uV���,ݛ�A-�QA%I%�w/^~��b��� �J������^;����������9�8�������^��v��u�@��D�E�cq&���ֽ��Z.�&���s@=ح�bN$�l�@��M�u�@�빠��@��;&F����0��S��woUOq�����N�v"���j�k�VK��&��$�4]�M���{���e4��C�n�b�2�MUX��/x�fnՁ����Ř�G���J5s4/Z���|�a��EV]�O�Ė���bJ�\���EQLrG������ƁU��h�w4yڴ��!+�$�8���˺ɠwu��=�j�>�SR\�m/|Z�Ժ�˹,�m��,�]�m��q��l�X�^J�3��EϷ-��U��Y]"I##�|��s@���@��M�[&�s�:�7�	�n$ә�|�׿bE��
��4�?��H8�	%"$�i)����?���M�����@>�[�q0o'�&᡼�~}�,������s`��" Q����e4��CN�Ʊ�!����s@��U�}l��}n�@��5�ղ��	K`�;V�P#)v��:>�2G�2�;T�Tv����}�=��g��6�j<���`u�e�������Xw�	�8D�"�#�@����޷a`g��X�Ư��D�B7�T�ț��{��a�w�����Mץ4�� �m"I�C@�YM�Ł��O^��a��S1T)@�HR޷s@��M�]��޲���RRH���4��I$�$��j��%Q발sX��^�p��֞dN��r�ܥ�^3s��^G^��9w��[u�gk]g�!8��u< ��m��5͢�UZ�F����K���Ӟ�Z�"�\���d�M��7t�� �݃����mۚǱv�m熹�Iݗ:7��g���roWNn��Z�ۨ�C�����t��>�n�-��u��b�c���L\��>��Us/H�][���/N���	f	DuɒuW�V��^�ru�`f6y�BII�Rg�w��Ɓ��a�w�����ۋ ��T�5$�)�,̻��Z��s@��M�U��8��R"�MQ`b�s`{1�Y��G#���Wŀ��tXG�sA2Q
��@�u��=�)�{�,Z��zg�I�HD�"�Rf��YM���9F=�Լ_o�`{��� ��E�M���Xۧ��J9D�K�vX��qͬ�����F,�]v�T�m���Šy^�@�[��w�����b�2�&妤��\�\��מ
�t �T����bK��~X����<��ȎBF�݁J��3B���f��ǿۚz�h{��@�^�S�ن,�HRF�����+���h�?��<�W�{��hv[�b�<y?	���t�hW��=�w4�h^���v^	�	�����ڊ�)���yc6Z��@:hĆ��O�ﾼ�-���qUK�b׳`{1�X�mX�S�`yX\�,R,2I���s@�;V��Yb�=_U�ى(��RH�l$s4���h��-79̆rK֔��|��<f��}�swz�����F��B��.![B\	p%%\�\�LO�wI�dwJ��II�'`�]
����;JC�N��j�1��R�'w׽w7\���I�\�-Ŧ�h�:�E�n��,�6Ԏ����+�9O���q�Fccl�J:>��{q�ؼG��]�mb�Ҹ���	ܣu�v�h&@�~��w�x8�8{�R�S.�7�V��]d��v���	u@��@�3����)p�H��8�%�SS�$0ėĘ�p�eė	%%%0���CUs!.R��-8	���It���kL����\.LQH�3�z�;���^-���P�5��ԡ�����%���)�q�w`�t"��.��P'Y!NkA
��Z)�tAQ? ��x��'B�Q@�8��(r[��z���	+�F�����:t�'�l�w�V�5�1E	�$�G"�<�W�^�M��Z�K���ٙ�����F��
v|��Y]�x�M�@ί
������<n�Ө&�Y���
3�B��6߿�������<�KyA�^̀1��A$#�'���j��H��E�r���@�}V�wew�c���q�_X�.��
���.����dBt���hJ(����s�Y-����7$������PJ
�Ȅ���7$�b�ݚP��UU6^�6�9ȏN��@{/jlY�l䦐K��]*��X�[�]v�9�����f�B&{9|��63�O<�LN��S�[n�ڂ�������u}c�9wW�r��@��1$�� ��zs�=�uz/Z������G�P��$qI��1́��͟D%廳`7;�6���qE��Eqh�k�>Vנw;c�;�)�v[0A ��<J�l��l��v��<u����̈́\ �@�#��@� &JbB1#H�bDb*���B 9��Nɭ�Y���n][�\ -����["�ݲ���K�4h���^�����t��D�/;F��Ҝ��*;
pz���&{Z;Z���	 ���M����� D%�I���G,ܫ;�^�s���P������.�t)�vD�<P�0�7<��3��X�t���ʆ�S)�;v��Wn�8�[x���a7���TAn :x��	�YH�=q����ь��p�mQ����ٺg�ӱl����$��ck3��.��G�}�^5��n��A2nR?���z{�4/Z�������6����7#�;�)�yzנ|�W�w>���,9T�&dR,1I�ֽ�z����@�t��r���s$ǃxI������׳`7/jl�S,/76ײ4�X��,�y�zs����M�ֽ�z��uz�F�m�9�5�4�OW]�"63I�S�zA�ny��d"�⭞�U��vMhUra��'���~������x�y@�^����-�I[�q�$q;�\��^s*�P�Tg�Wk�;�X��Jh���0�I �$��>W��;Ϭzf~J�?��_��]�0��7G��������K�����:e���e�������A����M��^��YM��ǠUy; F��#2e✾8y��ؘ�mu�z��7RWm�u�*ui��	cJ7c"�a�������e,���r:��ZXKک&��$&`��US`w2�"#�	%�M��֚�uz��i$�Db�țp�=��=��sM������7�h�S@��:�)$QHc�8��@�빠{�U�w����>������7��"�I���Zz�h��������s��M��J)��(D�Ue;:��^y���w��f��v�t�r����.E�I��^��Ɓ�;c�=�)�w>�@=�]��"_�p0�8h�=�e4��h�)�{,���Q8G�()#�;�S@�}V��Қ��@��"�L���1ņ)!a���D&��3]i`{��M�!� �R5@`D! D�$f1)��	HXBHE�	%"�����Xb�� �b�H�) �Ib@�1C�DKߵ���:}3��S.]�u�<rC@��M�z�@�YM���m������#�w���s��NG�AlBX�p�]��؍���s.:S\&��/�<�7�z�@�YM��4^��>�έ"I$1I ��ץ4��:����G�^|��T�*�b��%4X�L�1�2��G9�K���@���u�4�I"x���ץ4��=�Jh�)��]���i��%"�>V�z����䓽�nI�s���<#�! ������|�amT�l H���Uɱ�n\���H8�7���R���n۵sΕ.5�q�����E��[�2'L�@UZӹ�������x���.�e o��O��vg*����^�ڴ�6�,i���UgT�v�XS��%�r���[�<j��͈��ӓ��u��{��ms��4�>A�q��,�ʗn���M�]7b�:�C�g��c���IѦw�[�����ᑫ�h�մ�U��8�e��\2� N�w[q��_>�kK�m��u�$Ci1�-�7�3Ł�q���`w$1�LX��Xcrw]��$_��������@�Қ�Y��$��8�h_U�|����)�w[��}j2cm�p_�yN-�ۏ@�Қu�����=Y�ZmG&H�RH71�����n�k�+~/\�m/�J�1$�t�cd%��]s��s��v0@��$�<�ֻU��y���g]���Gp�;���-}V��mǠ[Қ�uu���ȤM��-�j�s���d�p��`f7q`�]����q� I���Š[Қu��W��>��.!��d��ƜŠ[Қu��W��<������m5�����;���*x���m���2��B�UH��.������l�����TN�s�'6�q]�' ���!�Z�7=�y+��o�����W��zS��l�֣#@�S�l��z�v(w��w4
�W�z��I"���R@�)�cw(�!DDW"9�-N9�17G�w>x�#�$�I�@�n�U��W��zS@3��i��ȜO#s4
�W�r���-�M�����di�!?)�8�5���ڬ�*�l�'��9��;�b�b�sm8+-�L`ԑ 	#�9^��/�S@�n�W���^Y&��Y#b0r@��M���^��W���0�Hر �����ץ4
������/�S@����4�<"hqa4��lM�l�X�G��"��T�C�j*w���䟽�d���	��nq����/���k�
���*�$q�,�XF8%pq�z��j���ݫ�/ebG��meWgۖ�3#�df'$��/���[�hwW�Um����<�� �H��4W��*�@�m�}e48�tKL"�7�@����h��w4�Y��V��Ɣ� #�9[G�_[��r��@����ye��+�$O�s�}n恋�̀�c��㉰=�Dr& �EO	]�!�%�Flˌ*~t��b�Q��.30��� ��Ĉ�A �	$@�A��A�i��	pn�f�:
��HB:]&:�Գ��"HL�к`�r�2���4���a�0!HV,�+C5	3D�.K�e�p!	��*oD6��H�i0��ˀ+p!$Y�c�\a�Ja����ip�\&�7i�i�hc74��̡�)�i�D�A�� B@�"��"������*~�?�  � l h  �� M�         �           �`hG.ԁ�Y'��]9�e)PBKpv�K��^^���r��[r9��WVF^U�*5���ьո�؊��y��ؙ�3к���gG���=�+����Fr�r�挠��7Wb���nx2��;k�=7f��Ϯؼt�"/��Ux�a���q(�E�/<��0��.��3��o0�Qu�U�{knÙR�Hq���6�HM�p�m��`YcEX�t%��n�\6l�j^`앗����'.M�Z�wcv9s��9��g`���UR�����UT�U�
�m��B5�`�3m��ݴ��Z�	m� ڭ�%2�����<��ڑ�MK$��i����H^;n�Q��yz�(�I�T$���(6�IP fj�� �Y���V�����0��5@[�mK��n�5�H n�$���A�ay����~�����F㭻qv6�]�v�mr��3�hG�8���<��tU:$��R�0lJ�QyV�j�U�@Caum���	�]2�UѲҹ��*h�CD���Ƀ�-��H����C�a�뎳�7/+�@�۬�[uɹ� r��p���K�q�a9N����8g��]��i����_X�4�q��\��m��m��nݛ���7����!�����]�>�nl-zc.�FV�T��/%�ݶ��֜�YT�%�-v�9L��W<�	^��b6�8�:ۯ�ck�x�fvlֳ�]��&�X�-������<}�v���S����3�f�X.hi0��:����P��{bj�i�q����kO�=�3���nz��nX�{n����t^��t�vT;q�d^֎x�V�#nyLFn�g��55��К�[�r!��,�YM�۬�WC�(fͺ$������݅�?n	]���eZk$[k\,��1�jvuu5�ֳZ��uQWˤH<(t����:
	�@�F ���cnIq�J�I$�I-� m�%����.��^�^$5V����Vgq�=�-�ۃ�n�n��nd��|::'�݀��c	���;*�M'h��ʆ�caJ�Q�Z�+
;�?e�)�8�x��A�f���A�R2�۷L�sR�=s�7��tX-��wT
F�K�qn�t�m]�z{��YHi����H��99d�{dK�O��l`�;����-�2�һ����Ҏ�\wd���1��}����S�aN�N��]mj�G<���uubD0��π�V�=���+��}n�s���m�xD���zY�l'�&�~n��:����G8��h�X����17��
��c�/���c�	�ڰ57�`{�1ȉ�����rA9�@��s@>��@����v�@�|�Y���y$PRf�}�f���l���3%�+�����\�T�[V�up��K1O5�,��[-�&��Ƒլ��َՁ�ۙ�s��jhwW�{Ϯ-���}�f�}؛�H�R�T�5S`{�ج��9���9)�X��Xf9�H�Z��J6hER�rUP��ۋ ��6����`UT�ȰRE�s4�[4
���=�h��+1�1��Ĥ�h{��=�h��)���@���#S����<Dn4�5c%`'(�۵˗uU�!��iy��Y٣�U6�phcp#�@��Qh�ՠ��@����g
�r5?,r4��|�Z��z]���]F����)���H��Z��z]�ss�1O	(@X�����f�s��Z�w<+?LX�R&���wW�{�u�h^����	Ja*�U6���`lG9�ܭ��9w���*�@�ۚ���hD�(٣ a96�V��!@q��Z�nz:��RN��jw�d��Ҏ%�&����h^��wW�{��hVaJ�H ))BUJ���s{�H��́��a`_;V�s���m�xD<q9$Z]�����h�h^Qcn�)��TJ�����DG#�3w�`nN괗u��ĕ��`P/����K޵��$�s�Ɯ��_;V��;V�Wuz�n����z�F��
��c����Yʆ�H��;Qw7jW0m��,�zl�<RI#!"yPn-�v����z���/��@8���D�n)Jj���c�؈�Ff�\X���z[Zz�t�q��f,�@������,��DBY���M��	��)EpD���s&h�S@���@���޷74�
�� �%$_�'"�=�mXf9�=����~t�y��r?:O���mj��p [A"��L8K��S������G�r{Q]�ͷ��x������t��'.ය�f�m3���7JC)�j	w�A����-��n�s�8�^b�����Hmj#<�g�S�Eb��.bn�쁠ظ|ݖɶ�Y��mn�v�R�u�kYݥ��]�y��A���=��v2#�}�S�ɮ���qn��W#��B��x7c������w|��WB"�ӵ�&�����w����m�2q�l��ɶ6`v��9�k�*����\�'��o�`{��ŀ�-��t��,m�IX���=�ss@�v�޲�^��y�+�N9�b��2f�|��޲�^��z���=Ϟ+#hqy#Pn�e4
����qqa��[��X!��
�R��RC@��^��[��_t���YM�ը$�X`��hFH7�y�V��*��N�gz9Y�x�ۢ�����@ve����=޷C@��M޲�^���Vw��^AD���4� ��e�ױ́�n����� �%�b��]��uzz���4�>VB9L�9�^����4�w4�(��t�8�(
G�_[��g�]�>�����uz[^���y1���қ�E���!����q�;�X�ּ��9	LPb�bN6���9@��M�w �����G":�u텁�\�ڪ�d�#��p�-빠�f�o]��� �9pV��H��h�}�nI���ɹ�Ȑ��L���-��}q�P��3I&�o]����Jh�@�/,��`�ȅ��@��s@�Қ{��:���9w'dԑ�d�{\N�g9Iv�Qwe-�n������E�.Y+"	&��2�1)3@�Қ{��1�h��Pnn�X���������G ��hm�h��hzS@�ԏ�A�$�#�)&���F�}n�ץ4�Y�ue�#3'�#@��s@�Қ{����H�0�$Y	QZA��$0�}m�4���E!��q���c�e�7��m�,��XȆ�~���6�X�ܳt�Q`���l���mٹ��ٙ����T���ynMT����n��v��w<�X�1ى'�kI&���F�oJhzS@-�4b�ˋ*����#@���ץ4޳@�n�@��9��g��<ɂp�:���[�hm�h���.p�Y	$a0O����[u�w4^�������?�6�i&���$�I *�����I˃��/k<r�ٹMv�z�8��N�<�y��m�������;=$�rI������W��2��kf�{1��I�]�B�X��J�-Ȅs\v�;y�w<9��u&Ni��b͇kn9Z�1�M�>/����o�f���p��K�d8G�Ks�g]��G�uz�kî78�0zy#I�_=��q��Տ9�޽V�����FUPn�]����U.�v:w)8�mb4؄f�0�c��2uƌ�a<���ɗ��g#�<�`����K@���w��oY�z���c��)��o]� ���oY�{���=Ϛ(�nO�c�H�� �[4޳@�v�@���q������m)&�[�h�h�z�h��h�1���͸�0�M�v�@���}�@-�4	�?rvL�9�&F'2�۞ݎ��sl�f�}�q�����眺�Db��u�"q'��R�/Y�~�M �s�oϸZ���7����� �� �ը�W#�!�X�lV<w�+!$S	��rI�z��;E�u빠��@��<�$r,q�mɠ{Ϩ�z�� ����[4y�*M�~`�b�Z�n�{�� ������@�ؐu�,�s�I��
���t���c�$hɮQ�-���^��'V�$��9��-W}�����h�l�>��-޷s@8ʭ$�b�`�rM ������@����z٠Վ�ͼ�6�X�����eܓ���f�w�T� ބ���VO�,%����iK�j�"	,JP!@�ZA��KBA��$��%����}и2B0�RV0# \�����8��W��	��-1���"�ЃG�߷�R�l^с�/t5:�鵂��h�h%7���g8�#��b�T��Dctˉ4�dCgً.��6$�2�*c�cC��f��	K��q>�vD��e�bF	,Wz3�P�)Ěw�^�d@a#,%��d$#�%%eei����>��f�GTƐ��
����������1��%��#ae!���e���� �w�S cF�I��"��;5]��KB��~��5������	���6*=��A� :��W�2H�a$�	!	'szL�� �#g߾���'��4�V�#���31wn�,3v��n�7��)�d��6�鐀�@jL�z٠��@��Qh�����jD2��s��n� $����!;b(�j��*6�m��V9i�BI��ɠ�Y�{Ϩ�����Ds�@fnՁ�ҦeU5I�̎I�{Ϩ��n�{�� ����#��$b�iD)�jHUB��`{7n,/76�c�ޖ�X��"��"kjL�<�k�{��=��K�<h�Qm����!
��"R�������"XJ%V����RF�Z��֛.B�BYI5-)ZF����%�6�"@1�I(JF0����$VXD�!	Q#a%e%��,F�Iem	���ԃ#P�iV�a�1�JJJKKH�@*&*:����rI�z_���c�LCR= ����v��>�����z�G[�ӒB~S#�D�HQ��#*Ƨa<��u�]��c8�Z-�&%sO�jۍc$�h������<�k�{��;Xw�i���Šw��^�F,ݛ �{V�-°=�3�5��~�����ֽ ����v��>����k�$RI�ğ�q���h������=�j�>�#m�an,rLnI�{�u׮��;V���^����ο�6ܐ"�96 �	 mt�/&{)�˹㧜V�v�o�����d�/o<�o6�u��7o���$�&�ƹ���c��M��x��,i��`N�J�YP+���/�Tȶ���.��+)�P������ô�DT�&����d��u���l� MԸ�6�)���x�g;��ɳ6.Nric$f�����rW�ڐ�t�=��mD�\UR�K0��pE�)�q�e�c"�m)��նL�ӌ- ���p���rݰ�X�)�J~b��$4��4yڴ^�����q��Hk�L�=�j�9zנwu�h����Q["N�L@�Z��zw]���[��{�ՠՎ�ͼ�&�X�=���@����=�j�<�k�;Aى��Ę�Hh�����Z��zwW��w��n52r�����ߥw"}̹J�1Ƌl�rc������I[��oZ���]������h^���^��[��\渲E$�i;�-ȱ%Ͼ��>��u[�/�s@�s@��M�R6������=�^��>�@�������@�/g,VcS��(�h���)�|�k�=z���挸���H8���}Қ�ֽ�W��{�)�}�:�%$�1����቎��j�e�YJl���jJʝ��x�Ine�����I�a��>^���^��u��/�S@/V;?�1�8��@���h�]�������@�\�G�2�"�����n�o]�٘��H�����*耰s3wM��{��fv,mѳ2~�ԙ�[Қ�[4[^��[��\渲E$�HO��8h�l�?���=����q`7���Pn���q�����/x�r�r�!�v�pc�^�e�R�u\$�4�ӵlۆ�Z�m�~Z�4z��ޔ�z٠\W
+6)��Gs4z��ޔ�^�@���h��2�$n �f���Z��h�^�޷s@8�+a��L�#�@=z��k��>���ܑ?
�!���O���ܒwՖL@��!�@�Z�4��9Ƭ�76�l^��@�$MqS�\�r�;k\�
�v�=q�u�xNӊ2ݎ�x�	�!�I$��d�F�|u���:��@�zנ{�{��f\Xۣ�"d̘ԙ�u}V��^���h�n/R6�mQUU4$)��+�wf��77jM�����`wR�A�T���	Ǡ{�{�w]�����l�;�c�F)RC@��q`bx��:۫���`g#�̃+�mk�]n h$ U�W]���������`;g������뛫��E���M�Fw*r!q�W�
9	$�������k���x��U.����u�x���8Ѷ�Z-����[p���:ǚ�.˭�zx�G7d����f��o����x9ݱ�,��p�v�1Δs�`�İA��}q��k��}����\W%��+�H&x�	UFfc/H�g��q��e�W;��٭�����X�ɳ^6�l�˯@��d�s�6]՚��<[�l���=��f;� �(��"G��	��}m��݆��빠r�^�_VY1pI� ��@�[��;�w4^��׬�;����d�G!�w��h�k��Y�w[��>�eō:�1�I�/Z���h��4�]���@�&�AF$=�>�~f6��v�#�q�96n��q<gO-t�O`�Z��&�QS5= ���1����c����s��ٰ=�T���UR
�L�!MN�}�wWqǄ�@���1�ل��ic:u��9u�@�^�@�+�Wq�$X�q9��빠r��@�^�@�Š^�.0��?�'&h�k�<�W�wYb�;��hEl��E�`�q��l�;�X�z������ը$�X`��6�4=l>w[t�X쉬,���%k��[;�h���8t$�ƛj<��M�e�@����9{��z٠v.E�W��!BI��[��w�U���@�Yb�>�2�Ɲlb$���9{��~�u����� $���z��s�uٰ.sY�L#S���@=�f�޲Š{��h���=�F�<�G���rh�K��[��{��z٠w�z�F�m���$�"j4(^Ϫ�)��@�Bg����tn����k I�����#�ȴz���}V�{����Š[� \a��NL�=��h�l�;�,Z�]� �(��G���I�G�w��{��@�빠{Ϫ�k+Ȑ�iG�Qɡ�O�+5�Ł�N5`�8��s�q.�4�Qr�ړ$p��H�^����� �[4�K���v@���N���xs����1��2����y���^Wң�.Y+�9�6��mW}���9�6���e:[��u{����L1�"��Ǡ����߳-��-�����ֽ֑��*���$��4�-����ֽ �l�=��댘�D�'"�/[��yzנ��wK�ז@�4EEO*�����<����ȍ��>��]I>���7$�TAU�TAU�U_�UUZ(���ʢ
��
�*��b�*���������P�� "�B����Ab*
�E��@PH
�E��@D��@@ *D *QV�P"�@`*
�AR���AE *Q
�X
�"�D��@E *T
�D"�E��@`* �U��AP`*DH
�E�R"�R� B����A��AX
�D��EH�� �"� *X����D`*���D`*
�R��"� *B�"���
�b��P *Q��A �"���@A��DQ�"�"�H
�T`��A��@F(�H
�U ����AB�`*B(�  *�"*",R��"ŀ�D ��b�� * ����@"���"�* �	O�� ���TAU�QU�*�* ���DW��U_�TAU�QU��DW�UU_�U_ʈ*���PVI��o��2A�` �����]'�(�U)  �@@$�`4 PP "���  
A@(A�  y@�� R
�P�J$�RH���T�
�B��
 ��� �T" �B�P@D��     � @( (��@=����<��sk����.p w���﷥x�����=�z��< ౽ڗ=��   �y4�8죏x ���F����{yG ��{[���}n�4��Q�  �� 
 @X yTݝ�<� �� b�C � �6` ���K�.}�C�j�ո+�BŞ}������e]� 9���{޳g�.��x�]�s��o  �>
 @   Jf �Un[�Լ�v��y��y<��U���Ͼ���{���{u���]�����]p �L��j������;�-K����p >�{jy>쫟n�9�K���jW��9�M�}z���׶^}Χ׋���||  P�
   ��.u.,��������w 
�t� �  iA��� &�)��A�PR�c@h `  4
� �K,� � �  @ D � "  � ��  � � 	V6 N�� � ��/o��R��P8�b��q��m�wl��Ǜ�� =>��}��ީsۗ��P��׶���� ӷ�s�u�/���4���F�� �,���|c%�o..�� z��iR�  ��2���  "x�T�I�i�@��R��R�	� �������J� 4ha!M�)M" <S�O���������?��|�;;�w��9�� ���5������AU?�QU�����
���S�����.��T��A$k��5�$x�6�8 �LMV�sE6*�CD$����
*V�h��w���ֲ8�k�k���|�h�w8�u�8�4E�Ӆ�¦���;5��x�H�4�ǊF�4n�0��#L4of��8N����3L79�!�vBsF�iss�����5���i��$Q��#Hd��I	Ȁ�RN ��jf\U�^;�9��g��%�u��� \4n�)p�m��G�c� 4���R�7���Y�T�̎ew^ZC ���h�^$�rȼ[�=Ȃ�Z���V��A�A��
!�~��2?P-��w�[�&��
4��X�L i=���������4��e�~>���00�A�]�R�ku�C�iE�m���
�����C�z��Bh�SGtor:x���+3[9�_�ƥ3N�i80����CD?$��!�&���6w��2䖐��M{,�B�( ؆��`,�틽��@�y����c}��h�P<�>ػ͏�D C�o�}��0��Ǉ�|ƃU�5>��<��9 ��mn?<�
"��Hx������ؖ��\ Q���^������<
4��'|�$x��Z�:M�:��i	���ӆ�,����
�L�y��%�C��*ʒ��5LMo�9L�]h�,i&U�[����s_�o�f���3?��J�	xߐ��Њ@?b��p���?�]1O������Y��L��F4�t٭<$H���#�}�ֱ�D*�c�x1�ǈ�"�D>�cp5xTiS�]�[m�� �<-��.	�zINS�x0ǎ@�s���.{X��L(,`jǫ�k��:�ĖxbX�`6 !KN�����Ox�B��{ �N�f�ݘ�ϵ��(��0��ccƨ������a�g��K0-g=��^�� B�-����(�q%516�e���k�k��,�nfT
�6�`]�g�|����ξ���yV�$SQ
x�X{ᆓ�G��E��r�u,B3��������7�#k�&!Ł�}����5�H%��M��Q�@���q�i��F��y�2�0�����'��?.h����g37/ �A:���Ē@�6��2h%���Ff�p���:�*I#3�>b���������3Cm(V�x<LL�}���aX=4h!4 ;��3@4FP)����S1�~0�~���+�l���F���H`���D���UU��H�JA���$c2�Fl�3��P�׍,��X�|��������q�mB�)C�\q�0�7���!Lu��!�F¥D�$S�D�:1�͐�j��0!�NЬ�dp����P���V+B�t͚.�!(a����Fڔ0bWL5����Z.��[�ąq-3D7����l���o $Q	ƩS�r� ĖM�+˻c�1'�~ڠi(@A�V=Ko���m4TX����	�i7x+%���h@B14!��Q�V0����hI�bL�E����xT������H�A�
.^I����� ���`��cA�i ���-����4M'(;�����o���H��M;�G�bP�[]HD�M#�H�F�e��"�v�2H	�����3ח���W@����y=</X� �4����yh�ǅ�F�,y�{�ޞ�:�U���$�ݧ��mS��c3�Fx�NAk<=痵*� 伧ᛕ�� ��g�����*�^��$ %�@��`/�<�v��@��.�-+=\�Ĥ\cb@b560�F?�k�$��ƾ։�1ц��.��F��@�B�+$l9���QE����wt<G0++��s�[?��"��R$#Xs��0�#^t
m�2[n�,��G��@C@5�h)6@v�����	3�����XY"���2��UD�<�!QV=���U�3I�OE��k�| A�d<`%�D��ڰP+@�r�T������h\��^���hX3�`���̫ ��3�$��\}���N @��UQEy#TA��¬g���l�:�^N�4����Z�e�`�p^��6�K'��:y��HL(% \�j�*���T�B�� D����+�'(�LG�����r��<��&o"qaH�G�!���]d�P!��<��|ŏeBB�^�����m Q�2��Nf�&	��0X�H9b�d0ʞL� I�rŪ�^�,�RB<Q��-
����¹:��JfΈ��\\)�
T�Ç�4�C{L�$�`��@�4��6?��n�^�����L��F^s׈JX�	�/gףռb�B���1�Η�k�a����[�c ��+iC�&b��JS˹�����d���22A�@�h	0�h�t6.kj�ݰQ-^�ow����{�=x�Fߥ����P�F�J���36���=ݻ�7�u�t��,0d��/OfP',`���k�H9u��-�9o'��!���cp!9����v��C<=&�D!R.Xl�`A��Osw���Qr�	���H9k1���R(�%@ɹ��o�h��^zTF� \����]A(˧cO�eziT \��;��׵@��W!�6<N24����a����`ˎk|?���D=�hڠjE��xM�!%�}�Ԟ���]Q%�Pض )�U�<��,@���o �����<�{l�܄�  ���鯮@�mu�dx6<X�G��pѪ�Ԡi97����U��wu;��v<B`���4�g��*Y�J�/qNC,�Ȗ/R`�~!�!�D tg�mz�	��d�H�5D��@E������B���"��@�(�`��.�5^˯�R�
LA)��/��Br�3��� �����)c2�1`�����<36���^,�
���<�� �4�����uL8B���	L��+!"HRe�!�	�G�<+�XS��&i��2�Ja�>�O��᷊�'�f_�D���������H'�0!
`Ɔ,��ٚ��2�.�
!�n�o�)>=�xQhې�Fc�~IR��=��Nר��L�������' w�7���4< B�Í�ø͠i���|�ւ4ASP2����
��a�#B�b"]	�P4��
� l6}���1ߜ���2gE<�6 )��w�$�F���!��T�05c/_�S}���4�Z���޾���)ۧ`pc\5�������yO��M�Ц.�&�&�pZ�x=��(S�D�x0�8t��.��3[֤>%�[�D�t�Q�"�mtI#+�~B4X!��B0 Ċ�1�R)E�p`�p`�� �� ,H D��p]R$�~.A��h b1)R	q"P��bT��	��6$J����6�j �J�^ �� `�A�D��ł�h�\t䌄$Z8$�
0h`bA(c!����� ~# ���� �P �R+I >+�1`D��##%LB+I���aq"���_����O�Ӱ�~M)h4���D�"TH1��20�@���>��|W:�*b�Z�$$(A�H� ��B�a�d"dR�`�Y	X�8��#�)!���ŢƆ��g�3[s)������H|C*Fk��)��Đ
����kD��|���jzcW\
d�0���M�C�dN!.h�@�ki.Ͽ0��	~HJ��-���Q����[�B~�o�����cj���B��ī�D�_��
�S��X�7�8��t�xӰ-X�v ܠ�}�,�����b�S� ��x2�Oy`� �u�g��Pbj�x^�d��&�W4s��
aw�o.�Ւ4Q��i�/xBk�'��x,"˗�Nxh��ױY-�
�02<;m��(9��=�8'�=Vۖm!�����j`U��2��͈�+���n����X��<7�5X4�j-�4���5�E�Y@����bǅ	�,��[@��y�5�&��`����kg �!`CA��15h�[��L��e�H���l76^�t6m�]���j���rՖ��]6ǯc��Q�S@�$T��	"u�� ���s7d
r����{�Ptx?O��,O�3X˃
E�)�.!�Hf��!S6ǆi��h4\	��|$%�Dd.h#H�$��"�"@��jB������#V�|�.�ւ7M|	�aEs>h��@��?�E��/����ӚՇ���F�"�@��@�dR˓�X)�V�:-��x���'�3����?Q4Bq�[�S��f��p�{�c&s}[@�R���o�Z4�s���]�(�h Ba���f{�׀"�8�򙻄J���$�0�sd�          �`  1#�            �                                 m�@ l    ��   �|                �      8�   @  ��d�g�*_*�"T�9Yj�����J
����٥�� ֲ�"l��*1UUp9e]���������+X���֐۲��R��j��S�T֚��� 4��UJ��yv�J��W��=���WUJʯ' UJ� $A  *��l�1�&nѳ��<$,��ְ  AĄ�PQ�P�����ݼ���8;GHWTz�!�= �[rD�[n�UE�v�Z�dUY��s��l��p/:���m�%`�VU��ee�r�Ԇv���KmZ�j�J�\[m�ӷ=�����n:��܁&�*�a����o.�\�U�;VvVU��U��ê ]�.QY[��(���;miaT̙6�+�/e[����h�Qg�v�\�zzce���h;h1���X):�����V@Wm0 tV�������m�����u�6`*m���cj3�fy�u�@�I�{I�mJ�dը���s�q���e�-U*ҫ�oe��k�j7M�v�3�3mr����UUJ�@`�ymrۓ��,���I�[��	ѥ���Ʃf���I��9WR��R��1�S֪����,v�X�l���6�e���n�-P��uZ��{X�-��]/��+W)��f˞���j˅
�� ��{Git>���׵ѱ����J��Zغ���sKW��BE��L�k�Z9����*51@+��pqvQ]���L�HA÷J�8ݺ���{n�j��v�V�2e���Þ��Đ�L+;t���+`-�=e������*ﺊ������:�ڷ#[m� 3�HG��c%�v;kS��nb��g�*b��\�8� �vd �����P-cU�v�9^���c�yfVKnCF�m�mNcrc6݂@^ЕV��wj��1��s�,����[-�^k��9m�h��p6�	 ^C<
�n�]A��� Wt̊�:�z�j@��&�g^ŽC�i5��I�A�V�9�e�&^k������ږ�$����86����l��+n�� -�l� !�f���6�tE$y�n�Z��n�
ZRZ��ۥ�XC�^� �	 mJ�j�e[�$�kX[A�m���8ճ��NnN����Kr�@@U�����4����kjX6]�7���f�*ݕ@��	I ��$�a%�l �M�Q%\�P]J͍u��k� Kht�հ�L��v�[R��/���[j�e{�g2%(l�US��m�[C���dH��H$$�җF�n��D�fI[��nx�f��V��yWe���P�e�^g�I�ٵ�,� I�-��6�oV�զ�  �] d��/I����kn�p��h���%���xYVj�eR�d��e඀ ��`� pm��m�m��KӖ�m�����\v�6�d���}���%�7n� �/R��a��{�@wm���� X���$�UN�<Y��i[E��Z^YY@T�ٺUU�P�U U     $�m $ 6�� m��� BC��l�4P,� �R�����UUp];9��l��j��5MO)��������J���U�K����wrq��2u�/if�*T"�^� �,\��7m�m�-���  Np	 ��� p    ��� �d��    ��6� �>ۤ��n��SN�2Y\��y3�>�h)[4��i4��2�URһ>
vn��E�@WT6�U���ī@�Ѷ�;vꓯZ״���xY�V�������V��D��`$ 	5�     $ 4���                h ]6�@  ���6�Ç��T�*�y6m������e� �H��ۮ�zJ�3Q���"�# +��8�F�@][[�]�ʡZ��2t��$^�gn]m�kQ��s$��ղ@@ O��   h    6��kz���a�� d�Tc���m����%�m]/�&�Wa�遈jֵ�ϲ�6A���gYe��۱�݃d]��cdN�X`��L�eӶMm|�]��A̅�v�l��(��]�^]�c�\�����ހ���	)�wL���Gi���  $9X�6f��[E���5mT��PTȫ�����UWcOle�yM�{`��:޷�4���-���f�����T�rώR�b�����v�Lm��&��'m�8֤P���Q�S��R�i�*n�r�;`��w�>~����~����-gx,U3���n�w�M#��m�D��ڭ�v�g����Y�˭��Q�Bv^}m�n�`�P���ݍSj�Rq�p��v6˪��,@��d��2���χg�f3����i��#�۱��@R]��nQr��kN���0�D�����$\�W^�j�*����:�Rif�e[U;*�ʕ�B�'%wGܪ��r�mo;�)ӝVnڞع{z�[�x��ij�5[��qظ�?g/REl�8l8�ni8�-ض����}}m[*X�b�q�6����5:� 6�+6�tX�6u�yC��gQ��J�K��5�
�J�Mr��ȥ���(�ag��L�U�Y��z6-�x�[\[�N$���p�T�{+r,�G\�J�v�7v����qS��d�����[h�N��u]�a���q]�X۝bjx�G(+:�0�ۜ5nܦ��Wq�+ڎ
��H[g��oI'� ݤ�zݶ� 8�]T���Ue��*���틗�hr{36X8x
Iǘ�s-0v�y�_B�	[���ژ�t] 	��m�mV�a���κ'v�iހ-��`*�����gq<p�M��;�m��ݦ�b)�����Z��B�a�$˖Ij��VmF�ey� y��	#�Y��*�WF˴pv�;���vvj���e[���*���5�� m��oIn�� �S�ْ��!t>�=��l�UuJ�  m��-�A/(�T�K���nZGi�Wl�6C Hm���mP絉�8��� ݹwI����7n��ﵿ|3k�m�ޠ U�5�4���&g;_i���෨9�v�A kn���[O+*�[JP�m��q=Y�{��]U@JO6�R��Ie�VB�H�袪�d 	 n�6�6�h  �y��&�9��e�zD���4�3 �P�m�F�@�`����:���\7��w��t9j�Ij�j�q!0��U�    �h  mՖ��	�s]m -�   ��i	���yv�8���ٽ�w�v�Ի-l�i^b��-�vخ�[��U�6(	V�a@�UjڠN6�vrY��mr�r�i������s�C�V�����p,����Eup;�6�HO�_�P>��'rLȨm�1I7K&�&�A��k&��6�Sl�c�nε�Λ,��:�+�%�/Z �"���v;f��`Z�Y�l�ocS*�U���������[꺪4+`�y�*�A��}��Z��:�\:*���W���MG/\�7�{8�#s���tg�ףyl�v�ӊ�^������VuwD�f�+�Ye�Rɜ��ƌ�4�ggD�:�g����Ŗ'�� ��Qtkj����&{h%\�PS����r�UT�UR���v�]-� N��lڌ�R�S��J���J�m�n�覶��wY@  87[Vkٰ  �v�$�v�v1 ��Hl�6�ڴ��-���{e$�գ��ą���n��H9����E�J�%3I�\K@ l�o �� �J\p6�b�$�9�jX��\ Z�8 H  �$Hpv�p		l�ISU���S�ڃ�l֡�*��j��� �fT�����W�:���Ј�u�]� Jے!�ܣɱ�VdA��Gm�G����Yt����V����ʻA���jـ���wI# ݶm���m��-		ˬ�����]� �t�Nĉ��@�U���kle�����@9��][@&�n�v�N۶�6wi����U��Z�6 ]J� m�H���Cm�e�eѭT������w4CZ���6�� �	  -���    	 [x   -�@ @�c��          m�        p� �[@   ���[m��m��	 #�l� �[p   m�C��    	        ��   �p  H   ��      �   �m�@  �-�?}��      $   h ��    -�H��  �i� I�l ��m� � $�o����0`� ��`�c�  p�.�       @  8   �nmpm�	����  8   ��[�n�H  Ԁ 5&�u��jۭkY�k�QPAU 
_�< p�W������ (��,� �0��'��<DH(�
m
�� "
�4���D����Q5�#�@�s`k����*�©��, ����@���(+�A����]Gp���@4(hPN���@ ?���+� '"� �B�  8 �B(!�(:U:��@b P����QO�D���b�Dh��� � &*����)a$�H�
��1d,! 1"�a
D�IHA"��0c�^�����?
	�b�T�DQ���"W� ~PS "�?�f�@0W�?��D����0> �D�P������� �X,�R  ��	b,T�E� E"AV�`�X,T��oZֵ���� �     ۶m�B��   ��j�h�R��<�N�R�$�g\�[��T��d�����q�Jt[�����Ú�u��T"��Ǟۍ����y�G]�ms��Wqٻu��dL�L�^z�)�]ۉ5��U�RN�a��͗[۳��H�l��ݣ�y�C��2��]%��5N�-X�mckm��<A���r�8wH�*��+ɹ���e�4Ò���N٥�������:A7���G]���j�X� �Y�ɱ�m�ǝǱ؞����/TC;���Ю��@h�8��v�K�Ҟ-;=�!:U�t��[W�{8ٲ��9�R<��d\FL�b!�j�s�m��:\c�����h�nƶk�Im��x"����@�C���Ҡ�����M#Ƈ��t�&l�m�� 	 @ݶ��"�˷��*L�l�<�g�`��\��UUT�T���As��M�Hgex�Q��5V	6i�(�e�;i��C8ƎW\�ж˽r�mqm�k�mɹ0�:�e3��A�q�І:���v9��;m�v3ܫ�k��y�nC��A��r{�id��Y��vI"m95p�l緈]贋��������v�m�u;GS�\��W��¹����x�X�U%:���X9I�]pm��sl�S%�(%YJ
x�vX���{l�ش96�n�m���sq��QX�W�m�+���,����*���M��[���ͬ=���xv�S�S�v�u�E��;�Xm����=p�e����\]�̻kn�ϓť�p�\�b���-r�KzZd�LC,B�*U8S����٤��Yx��-�Nܚ�g�ٝ��-`GO;u��3�z��sCθ6$��5x� t�ps�8y��)Û�n��)mU!1�K���a��l m��<�����`ڥ�l8(�q����ڑ�I�9��Zv˦��l.�,��is�KUU*�pNd4�j�zR��j��?�`�LA��)��@ ��;��I$�&�pI`��:��hɝ�3��m<DNε1�8�ƒ�ޛ�볧p��z��{\g�:�� 3�i�#���,c�e��ػ�t��;�&$�]������ծv<>1뇇O;Ld�=+�n������S����6ѓ�vީ�h^��qӌ�caӖ��s�=v jS�sۗڪn�W���k��*lEiz4$��/H^L�u������Þ#<����]�O���9��8N��nx��l9��&C����K��P���,���!'s�c��C?o}b�?u���5#e��rY'=�a�=����� ����Q/��Y�Bd���}�V���uh�Y�}�]Zy
����D�$M����@'�u���4���� �K�|K��n(�Z}�h}�V�}�V���uh���~8��x� #NBx��$���\�d�;R��չ�]u��EX���\�B�%$�O���d����$緬Y!}�h��c����n<rE�_wvoI����c2�!�0�S1+H!a2��
.F�RKT���Ƙ��`}�01g�eY"$�L�I���uh�Y���%�f{��ZhR���#s�ȴ���>���������/|�6���9�M���/���>��� ��4y�vg��1<l4v�ӗ3�v���x���څ����+�u��U1�����ɓf8���@/�����;�UB��K2Dۋ@���4��@�uՠ똱�����n(�Z����uՠw���>��� �e��x�@�RB��I�oX�N�zŒs��,�s����Y�#�L�$Z{���di�}2u���4���
r���2ԁpvv\�X�'�#b����$�]�l�\���~�F��ddh�2Ⱦ��� ɓ����I`	9�;��s�ȴ��@����N{zŒ}\�lr!�cqC�I�ti��F��F�I:��
%�P���2c�n-���{�� �l���X��@� p_����Š}�/��D�D�$F8�{�� �٠}���mՠwuߒ5�21Dkd����]���飰�s:���g���۴�c24G�����2bm��@-�hzF�H���� ��_Wv��Q��I�}���mՠ{���m�x�Y�#�L��Z���=�uh��޷V�˘g<̰k#�L��-޷V�[l�=�uh۫@9^��2O�c&6I�_[�,�ߗ�l���H� ��J( �(���1�B	�RP
R��G2��[_��{Ϸ{��������UU��5uGj�eWDX��������������~����Qk���G����k�k��ų>3�r뚯J��ݸ�C��	�����;��Ue�9Ͱ�x���VN���ps�L��yl��C�9�q�v�'\ͭ�����+�w0��Ո��:sf�er#\&^�Z��[m<�՟m���]��a���0�n��nӒ��n�4E�]9	9���ˇ��R�Fq�gp,yP�^�����q^;h�m�ˤ��۝f�h��5�̍0>�0	�:��
9�BQD�-�d����URG�����X�F��(�N_W+�e����0=�0	�:��di�3#L�s0YTdqF���f�����/uՠ{�uh��i���"qG#|�XzF�24���4�'��Y����۝��@Bz���s�K�v��l:����s����m�����;w�w��3#L���='X{#L'�̕�����5�$绬^ jH2I	�#�H$�*�$��T�*��}�`{�`L�@�z��|i�bi��_[4{#L	�`}�`z��W/�8r������Xm%Uy�~L��0>�0���>	D,3&Lq�Š^���IW�o����`}�0�9�~{OM��֒����k�� ^�GX\��c06tѹ��v�l�v���]x��n`}�0	�u���4��#L2]�`���?��������u��@��}b�9��I9�i�X�@��F�z���`L��}K)RU�s�`%��d��`���<��H����=�uh�f���ՠyy�g,1��8d�7"�=�uh�f���ՠ^�V�����7��6���`c#�y��=v�X�����V_Hr3�g[M=^k���3NH���@�[�@��Z��I�����
e�H�O����T�ٻ��n�LI:�$��@�Y�b�����Φ��L�4�$�h���=¹1R8��Xc�c�@���$�`fH�U%�(U+*��`0�`,��$�E	0,*1���:�fgvnH{�1c*"��nfG�[l�;�ՠ[n���Z���1�pX�y�.1l�۞��_Z,�p9����;kI���C]�˜#���c	��C�9rh���-�V��n� �٠z�#��
Hb�����`I#Oj�Uٛ;� ����n���r�S#�yr-פ�u�����4���Q_)��ȱ�rHh���n��uh�l��ϩ���-9R)%�w��,	�4�����L��r$�*�O�[i> �ז�B�k��?s��I��;s�,�UrT�Yf�2�*Vzw#�&d��g�6;]�tvؐi�f��/I-�lzġB��b�;�,{h��JMOe;�n�&�ō�l������[9�����aZݕ��[o\O����s��ݭ�ᬬ�ÞŲqp>��a�mn�	w�^�c��;|����ȳg��AO@Kk`br:v�n��w>��[��`�Q8l�q�p���g�da����z}��kb�Us��jݼ%�n���Z`zg`�'��=#L�K�[����Šz���_[4����uh�DcːYύ���}l�;���/uՠz���{�l�̂2(�x��;���/uՠz���_[4��m�RCy3�h24����Y�����X�`K����y��v�.��Ɍ�l�g@��n��P�1+g��l���5��u��螥�I��Қ}l�;���/uՠxn���q��1jI�O{�^U
U@I
����)���;#L	%ՠz�������a�70y&I4�0&di�靃 ���b�d�><	F�Š^�@��M ��h�uh¹1S'ư�n-fvzN�'�i�3#L��n��������ȸ����>��ӻb� �l;[t��!��&��3T�tnF��]����`OH�fF�3�`��0WE$��������$�]�&���;� ������Ns�$1G�1��{���JiV��羿�60,*D����(J���)(�+(V�I@�H�H��IXP�aP����U9�B9��S���B
�
��
�42s���»9\��7p�Fc�\.�#���K�Mh$˚٭1n�shև8��i
��XU�%aV��(bD`���N��
�B��j�*:60.;���m������\n��I]��nM�F�kt��Cl
�Ѝ�]��y]m��%��4�P�D��SQ6%���%�����k0%YRP��\P�YRQ�cI@�IBѠ���Ŏa)�SY�$�m��\Iqe��Ņ�P�%	@��K���1J[���	�Jc�.2�B������X�Ԍ� ��:��D���B>�O�g��9�:1$%h[)]h�f�Y��Ѧ��i��P��	Ir�.h���P� ��p�H��6퀿���© : ~At($� @ ? '�)%���U$�uRIRvOg������Y��n��R7�-ޔ��f�o]Z^��qb���rC@��^�o]Z�]Z�)�~����ʛ�|b�@r��F��y
iݷ!�cKһ�;MۆQ��m��Ch8$Ǐ�?�~�j�/�ՠ[Қ���T��D|x21���uhg`�=2u�&F�ҥJ���mi��Y1Ʋ8�߬�h�l�-�@��ՠ�3ȡ!3�n��I��0=�`��ERB	�a�D`H�;����8���$��M�׫@��n��t��{�����<�u�:y;s��V9Ŏ���7�}��'����VHX�:���*��c������i��g`�=�`OIƘ�qf\vb��G"�>�Jh��hֽZ�[�@��%�&&(����;р{�:����0>�0>��U�r9&2FfG�M��ՠ}�����M �u���d�>26ۋ@����>��4��h�^��0�	"�aH� �H���� �I"@��$�"�`��`%d��{��=;ѿn�w���r�,a�ܺ��K���ԫfK��[l��&;`岶z-nf
X�q�d�:M��r�rl����X�ۣ!���"v��P�Ȅv�0��<}:�\�=�/B��Kۛpcm���;�r����{m�v����gy���v�%T�Y��<�Ym�	�s�n��6Z�0�7m�ݮ�s'0��i^�؈V���xz�
r��w�ww�??o7J�a^�z��Cb%��ݤ��3{u�-j��˞�	��F��3>E�k#���l�h���;��Œs{�Y$�t��(!�%M8�p��'X�i��H�����zK�X���#�@�uz���V��t��}�@�K���H5L��@��uh�Jh��4��V������۩�R7	$Z{�4�u�z׫@��uh�_���L��&����L7R:3�Uܼoy��F.}�t�rfΘԊ0�|����i���^�޵���dk�U�����t[}�9b-�6fI3@�Z�h�]Z{�4�v����]�|do�@����;�)�{�S@�Z�hx�2!e��"Ɏ4d�@�t���YM�kՠ{����x�X�I3><s34z�Zz׫@��ՠw�S@�����=���'�7n�㭕y'n:�h�&�ڸ�tJ�[��Y�V<�����N�n�m���~:�����Jh�uhir:�a	�ɘ�qh�uh��=z��;ֽZ�Y���7VLN7$Z{;�F��RV�BUR�*]�\�q׫@�[�@�̩�����I ����='`g�4��g`���t�I�������V��|I|�}_@�g�@��uh����<X�vNvy�e��Լey,n�����۪n�W��:���bE"�XJJ4`.3M�d����$�S@�z��;ֽZq�dB�L�����;�)�}�uhz�ՠw����m���$�P�32C@�z��>���@�uՠw�S@=����L�NDۋ@�������Қ������d�x�Ld,F�nE����=��=#L�Ki���;��f�p'g�k��quPF����8�<j�	�g�����~�|�����K��d۽_2wFzF�d���#LYʦ�'2�F�I!�w�ՠ}�sV���V���M��ЦI�X�1�wΦ�%���#L�J��d�	7Z�=��W�3���n-��Z{�4�nh�^���2!eD���FH��Jh�k�;ֽZ��w�o��~e�ʪ����� 0�ͱi�Jv�7f8x���5�3�#vNCrp�8�Z4��1%.N���H�kt��Z�2�k���"ەwl�v�T�㳜L[��F��R�,u��:PH�5ٞ����]��;:y�
�|��Ӑ�~����s�/8���n��u�(kplw<���ng(�B��L!��s�
4�{�{%��,��h(�M��cC���wk�cG&�;����S��:ݺ���j�����pq�s����Js�v�]x�9���]>ZC�0�x>�7���i����ʕ+���� �~M�?��C�I#�N��ؿ��#ۺ�d����j�U��6���/��#Q3r8,��}��$�q��U%����߿=Z^y�s�X|q�9"a�2=�o�8�W6oɁ\?,�	̙�ԉ�$4����w��{��Œsvq�N���e6��4N�u�mƝ�<��t����j��78����6(���'0��I�}kՠu�@��)�v^�@�����X�q�����}߻�
�vR �'���@�R!4�"��1"b�+�"���)I� ��I��Y���Z\����s;�I��8�a�#P`�8ђ-��M��z$�K3��ߞ����h��e���(c�d��u�4ֽZ^���e4�6�o#���/Z�hIUTٿ/�����2d��x$�Id�u��FQpa�;i�g$�8�:zTm8y���\�!X��lK��$:����#L�v&N�&IƘx��Fc�����������f�M�����:�ՠr˅X��M�"�� ��h�z��%�_]Z޲��V�j�4�dP�M��V��#L�v&N�=+r�:��cqhz��>����f�z׫@>�ۿ&4)#�c�|�L�3w`/@��>�N��cs�9��C��9����]d�2E�}�)�z���V�׮� �ͶY������׬�/Z�hz��>������ǘ\#�f94��4z��>���z��#��&cR��Hhdi���� ���-*UU^J�\���h^�Ɂ��Q�	$Z�e4�٠[n�@��V��f��f5��p%�ng�� ��9���b(r%����:K��!6�q��I?N�&H�0324��'`��
\���BfEI4��4w]Z޲�������?����f9ّ��;mRT��=7z�ٺ�0:���P��8ђ-��h޶hz�4w]Z�ͶY�����,� ���׮�@�uՠ^�M$Ɣ"A�A�8F��
J0�B��	YJ[�;�JU�a�aR�$%"P� n.d�aKYIB���PkB��>ѡ�
2�),��(�ԥ�҄00��,�Kd��-![IjK	XMj��5H�lٶ4n��g���1"#*A�@�6�`¬����WQf�kK))+#
��K�W��\������l�����I�F0�3HCL"M�C�M�Q%!FV$������0�j�!!XP�4aV�$XMsXD�	I&� ah�XR��ҡ!��3dj�@�t�HH�B�ل.:d"�@�l*`"D�WX�B0�
1�򄙢I�H0-`j7+ef0�kZ!4��0�	j�[�d3Y�����&��(��d���~߯�ߐ�_��p� �      [v�8$$    $ M�� t3�6�;����X�*��nۓ���Xn�VY�q��@ ��0kK��\{V��vwˌ��d�0�z;�Dd�V��X��^�ͶػFw��/ 2Omv&b�>��f��!v��L۷]�931[p��p�k�l����9�)iU{y݌'�%�X;Pv5�t�{kZ�u)m׬XC���[��Gn��Z��ι���Gm+�`����8���Ubl�l)��"��<GV9�&��LS�0���������^�*&ؑ�+uoJO)�њ�G<��l�t����R����(Iv�ANv�b�v����K�H/��e[�s�I�m�$��{=n����� ����T�xbTK����㔛���*�r�/Y��T�m�� H p���nW[����F�v،���T�:jڪ���
� 5���}_��}�xyX���i�\b;]�%���y��6#i�s�1l��C�NR��7`*�'w:9�M8.��eC��Lɶz�+6�m�uV������m���k�Wr#������^�n����`	���â	)sWY0�۪BhN�s�KKok�vU�l�C���9�JӵCqj:��G�8��펬k�vu���݌i�,�[��	!M��ml�n�O/9ق��t���^̼c4�g�:M�m���cSm�QuѺ��n��b&�&7.�nZ���qӼGi�;<�sM��y]�����n"l�D�:m���c&v:��ˈNN�.�r���n:�s��ŝS�mBۀ�r��U����W-�e��\t'Q�RS!!�9mT�u�[��ٳ�݄��e�Hc�ݙ������)�l�q�^y�c�BqsA]U��W��p���kb:٨���J���7�|m�� �L@s��Vv�6�6����h�km�Ͷ�m�a�����鱵���K$jSk}v�T��� -��h�$s6ٵ-H�۬� Z)�X�+���{����om� t�[�M��:�y�L�q�/nwm��nTی�[��"���q��c�nw�v"Gc���k�j���1
+�<�ɛ�v:j=�
ҥ،����|�n�b>�q5�ܝ�Nݞ�!8,�=rxf�X�5�y�t���i�%�ظ�n7����JW)������z��]��Iw)v�[z,Og�Eɢs-��Q�@��X��:�Ɲ����wrf���m��x�ݏa۠n��;mv%��;`n듫j�Yẩ���@s�sRs��&�}̍0&g`�>�:����x����L�$4w]Z���l�=z�4^�X;�$��{ަ���'Y�UU*J�6k���j�<���~4H<d�7$4�I��Gс���fv`��}���qɠ{��4���٠}�Yɺ�`� �RLsd�)n-{k��LFՇ�fJ��U�Ď��pv�4ƄE�9���;���;�S@��נ{�v�Lϓ�x�1ƌ�h���v�IR�*��Y��8����Y'wz��B��K�|�vDqD��8��I%��|�K�zᖒK۽�1$���I$�ܛi�`�D�9�,Ē�޸e����`�I-�&�_  ���Ē<D�d8�2���!��K7{bIou�6�K7{bIyo\2�Ic�~{�Y3s�\�s�nx��a�Ty �`�)lv6%`(E��ػ���.:YȲm$��!2H3K{�ɴ�Y���%�pϨUP��^��bI|Ѣ>�e�nHM���o`�I/-�ZI,��Ē��m$���]G$@�Te@�pf$����-$�n���UT�޻�m$�n�Ē��@�&�Q�!��K7{bIou�6�K=��1%�kzÉ$��JTlr1�\N0T�1$��I^{pf$�-�ZI,��Ē���㤢l3 #g��]tt"�n8n+s�ñ�V�r�h٫5�u%���h����{{bIyl襤��o`�I-�&�I,���|�)�ZF[�1$��tR�If�`�I-�&�I{w�f$��v7�*��T'�ZI,���%��d�_���}�1$�t�)i$�q��d�� L��$��%�>���m$��}�1$��v��m�|EI FA�!!$N � ��^��9m��e��FA�i$���3K�Z���bI/w�`�I-�&�I,ա�&B	ພ7{;�K���"�^�')ظ���q���"�HLs�I��Ѹa$�R�p{�%���;I%�݃1$��쟅V6���f$�Ϫ|[�H�i���Y��3?P��$_~�vM����`�I/k����6���%F��ƉNI*A��]��d�I-���� m�9�N�I{����KOrv�&3A��JBm%�o����I-�>��I,���/���fi$����o��L�В��%�s�v�K���}��$�w�d�I-���%�P�s��~ :'i��WF����h��J΢'�㇎�5�6z6x�u:���a�-�h��. \�vC��f_\�N�&�-t�d���������3�Z�ۧ����Nn�ěk��+�ݷ�{FM{v+he{']�zk�OG��rv�r��m�Xe�cUEs�$�;��㒺��\�]���F�׏='���v;1�{���f�6͢V,9�KS�js���d3�t�:\���]�$A8�����֓Go9{9-e)�"�X�KI�fs[բ���� ~~���_�%��d�I-���  ��K�Ϣv�I|>)�$��U$p� �I-޻&�M�����%���;I%�����\F�=P5E��i$�w�f$����]���%��d�I/q�#��A	����I-�:'i$���3Kw�ɴ�]��3K�T�؊"�
GNH��������[�vM���w`�I-�:�����z�Y^�)���������]a��mn�ֵpv�q�a15��ѥ��2��1$�z�I%ݽ�1$�\蝤������KOrv�b3A��*Bm$�{�`�U	"�s�v�K7{bIn��7� i/q��
f����I.�>��I.���%��d�I.�vĒ>'c/��Q4$R9��]��3Kw�ɴ�]���%��D�$��"y�x��(�A��[�vM���P�߾���K�Ϣv�K�{b �'��%��"i�0���lu��x	0�ݸ�!���\�;=�y�3gLj���v�#&��I	��]���%��D�$��{bIn��6�K���	`��R�pf$����^���%��d�I-��Ē��9�#���DӒ'i$���f$��]�i 1B�������[�tN�IwiJ�
 �rH�RĒ��m$���bIn��;I}B�߻�Ē\~�;h1� �p!6�K}݃1$�\蝤��o`�I-޻&�Iw���0'�.��y���x�ݎ)�ސ롗���պ�][��-c˕
ˬ�We���I-�:'i$���3Kw�ɴ�[���$|v#�*�%hH�r'i$���f$��]�i$���3KuΉ�I%��.)�8��*(�f$��]�i$���3KuΉ�I,���%����aAE5rHM���o`�I-�:'i$���f$�U���3	��\<H�<�a�YaJQ���[�tN�Ig��f$��]�i$����%�
 oZV��l4���=��BMێX��S�v�vc��;�˹LO\��tQX�"R�T#P�������w��	n��6�K�����[�tN�IwiJ�
 ���RĒ��m$���bIn��;I%�����KOrv�3
B�*Bm$���bIn��;I%�����[�vM��Y�[+�d�ahInĒ�s�v�Kݽ�1$���I%�����GN�zERB�		�D�$���bIou�6�Kw�bI{\蝤��*��  �w2[�I$�2ܐE#�����9qs��8�	�=m�����om���GN��Z�u��Gj���ӓ�A� ��a�P\��
P|�;���`��Ga���u��JJu�;<$�JBn��9�O+һs;QC`{-�Q�64�<o<�+i(��&��{Vp6ڻ[=��f��n�iyΩ�+V�ϹO�Z#��Gu�+H���6�:��@�ݯP�vl�o���	�Kb1+�c*���C���+�$b�2#�y�U6����q��<�.1
�9$�%��]�i$���f$��Ή�I.���%���a�E5nHM�������^�:'i$�{�f$��]�i$�8�6��� �T�1$��tN�Iv�`�I-�&�I{��f$�=��4�-��&��;I%�o`�I-�&�Ig��f$��Ή�I-�)R�D�C ����[�vM���o`�I/k���Y���%���O��a"��vr^1]����cd�m؎֜a킓��`�:��s6��H���lk-�[~����3KS�	�I,��Ē��m$��l�1�ٌ�#M8,�����B�,(B��bD���HTRt�̚�nF��`wadϒB6�RIǠ_uՠz�ՠ_uՠvw\z�ٙ�j�5��-׮��������/���*�����q��$Z�]ZguǠ_uՠz�ՠ{ݙ'[&M]���<;[���\���-���W�b���t1�y'�Lb�E3Zgt�0'�4���֤��ܚ�rWw��p�c�a�Lz�]Z�]Z�]ZguǠ{���ZՓ)$$Q��L�0'�4ά^�%EQUR��e	YRub�"��`�[�u��^����
����6p����АCz��b�B(c0ˆ���.$����a��	�R��B �&h�mKwe��@�D�-��'��]��$M�*0�XB:55Z��L.]�7��+�E�E Bd���Ĥ�e4�(b�ȼ���  �D���!�QL1>�>PGB�*�/�W*��}����&F����<ɏ"3 �Y�-�������/���=z���[��f��H���`e�K�{#LL�0'�4�����
 W�	Y�x0�5rgu��Jľ���'Х͝s���%XDFU���=���#L	�0=y���<�39�MRF�d!�E�{���/���=���}�V�U|ʱ�"Dc�}�{ަ�F���|f��n����k@��r�S5�L������uh���"����Z��+o�E �7#z�������]ZWս �cB��RB��1۫@wݴr���q�\�K�7(b�q��Y���ɘHH���>޺�z��:����ՠw��o&<�2cp̑h�ՠu}[�-�@�z��q[��0nc�$x�Šu}[�-�@�z��-�@8����2)5$q���UW6oɁ��&F�9��`]����L�G�E�}�uh��UU3w��y7�`zdi�U�嫸oʪ��A��;�����g�.^c���&�6ٴ�-��5��v���g�g�gv'�'\���qH>�޷�%ɡ������i͑U�Ƿg��nMɞFup�u�ִ��x���7��B�'�[���n��/-�7mc :C[۞�\b�a�t��{c��عjv��n��v��\u˷;QvM��٭Fd,Y<ݗ%ۢפ�q�˯�{ݽ����w�>CM&�%J�b5��Iۦ��r]�J��S:�*";K�F7d靝4·K���{u�Nd��`}24���0�d�|i�dP����o@��@�z��;���=��V��Q�$���=z��>޺������zz��+Z�f�qho]Zz�ZWս��Zp�����2cp��S2F�9��`zH�鑦xv�`ڄq0�h`�!�3��88[;=�nϗm������dK��]&�a0���ZWս��Z��V��n� ��
LȤԑ��=mխ~J�p�U�U}/f��ݚ�'2s��fgc2���c#�"�>޺��uh_V�[uhz�uq�Dc�$�E�V[u@:����{ݫ@���P����1Šu}[�=$i����2F�خ.r.���-զ]������v�]J���[�Ņk�WSp��G\�Y��K�������0>�`fH�'2s��.��T�h�B@����ՠw[�@����z۫@�]�$y1�fH��vnI�s��nWQF(@�BX�D#��E_�pM���X�N{�ŒNr\�@�M�24[����9���0>�`fH� �f
C"�RGo@��V���ՠw[�@����\�T�8�������egBϫ�
��;5�k���Ě�mEp"�������dy$Z��V��n�Nd�5UU/�3wZ`j��U�w�q��E�w[�@��vh���=
��Z�G�>6���-�٠z۫@����;�ՠ{��<sԏ$�G#z�����ՠ{���@�V�:H��$0�1`�H���B# � 2=T������s�e�pݚ����;�_z�L�07f���&�o8�{{�Y'<־���2܌�ԌL�u��J��ܷ�CR��n�\��a)�ka'P�F##n�-�����z�tY';zŒNj\:@�Q�24[��2s'8��ٺ��5��`L��E"q0�����ՠ}�uh�ՠu}[�]����Y�Iަ���~L�֘9��a���f��˙���ə�$�I�}n�'2s�	�`}�`+��I"�Tt�w~?O���O��U��NReqy�\1�a�����H�w��rm�n��Ug-��u�+)٦9훨��ݕ��[��ؑ�!vq��Ɩ��Y����N�	i�����<q��w�����C]��Ŝ&����e��ɻizh�&�Pzv<['��;�w;[��鎕�ל��iĶ3nO=��;�Ɓ�N�a�]5�	;�Ӷ�;��������Q�/�j�p�V�CҞ4t9�l�����c]8�cn�=f�AX!�m7���͍}�c&&��q~���o@��V�����/�ՠw��Zy	�90�&=�]O����T�8d������L\�|z�R�;��?5�L�H�"#�@�~��@��V��q����;���Y&F�9�t/�L6�U+���02�m�3#L?P�@/o�`�I�K����d�4di����̗�̍0>�0'�i��.��������9:��>m�?����cm\od�o1�����k�w��w{����|��R"rH�>�������V�޷W�(��_w��$�� ��S�C"}�`}24�P�$�	D�_.p��L^�N�>�u�����k�5�Aȣ-�#�H��ߵh��=޷V���ՠ}U��*�x�c�C�I%���|`fn����i��R����076��5�$mȊ�'d�{�Œ�T+w�a'w�Y'�w��N�Z�*0��l4��M��T�Ҿf�qs��23r�/bm���1�	��U.�F-��)180����,z�Z����=�uh���,�6�26�2E�{����>$��c�;�}b�>�u�����=�p�Ha2E25��S.M�0=�bI*�E!$�dV`E�z"~s>�]Z�n� �݅�C�c��9���I^f�Ɂ���ޑ��U%y�c�W3.,���̌����[���UVf���2���ޑ�g.W9� .�V�&�q��V���ON�Ɓg����6���љ:u���{��"~����.���37Z`z�%��H�ޑ�Ù�W�%�Z0B�I������U�?~i�'��0=24�������N8ې"vI�wX�O��b��R[��ՠv[��ޡ�֦`��L}L5*�y��&l֘��|aʤ�G$�|�~�V��.��ɆF����S�#LʿRUS����7����I��q��L4R����r�������X����Lt���YkPzh���	Š{;�=�n�޷W������_ڴ�V~�	&La�G1��{J����֘�Z`z�%���J�"xrK�+��m����w~�Œzdi���J�.M�0=��0"���.t�d�$jI��U��`�N�I24��*I^f�Ɂ�8j���;`q�(c�@�w\z�uh���z�'��Y��H�D�/����hR0�P��sK@�RPZ��w��u���"db�c�!�2B�~.�;�SA�B��`Bt]a�!��#c���4HH%�ByC0�	��a))FՄ	T)�]l�D���{7��M��D���s6�Lv�eI\�v�A*��RYlsY͒��l�%2�!H����p���ԓg?T���7h)�C[�&2������.V�Jh���R[�<G��om��s�L�4c ���v��4`m�H[`��t5P��0��}�'t���o���� �  H      6��8$�   �	6�6�#9���n�pv�;n�Jбm�s�E��J���V^�mG9%�\�g��u�\+W��95�&L�8iv�X��4-g��Y�7��x�ך�Ǔ�V��c���Ι�Z'!|�E��Ӭz����>kF�{]��rl�)��0������ڣA`È癶��c/�[����Mܼi�����:�]l��'o1Z�6&��OLzβsv�)ls��J�Խ��7���W�7C��A��:׋6�&3�n�'���{,[6бq;WE;��u��.;�:tԃ�nS*�Sأ�C�)m�]I�ҜPh�h7<l�]!�][T{bɊZ�3�nN_]�`^�U�����8�F�)v��U�vivy!��1'��*�;����ӱ�j�mj� @�v�x.kc����m��;���nF��� $�j�P���%s��Gb�f����]NB���mq��k��r񰔄b�8SmŮ�9Mf!-7����n��6{u��Ν��g=�����Z���m��C�۷-��OOgn{�wm�m���+��dc���ώ�a@�.y�c9�ʘ]��ּ�x�h��cv�cmJnF�����&��TF���pՃi�]C$����x�qI�9�c`�۬��Y�&P��&/[M�����>�y��.������#�lm3��tb�ò�a�5ԬK]J:�"Ԯ7l7��n&��K��YF||�6���-�L���V��-��7i�Z��v9����4�y�I�u�۶����c�Ҡ� �<�N9�J�������]]#�[J�zl,eL�+�Tƺ�����͝�����6���k=�.�n0�R�um��'nɎ�=N��\ruD�k:���(`d�C�[S��
�\�*ԫ*�UJ0H��V��c��,2D��m���m $ �[UU@������H����Sf ����-� �i�vm�ѭ[u�����E]���!�'UEt�Df��3�Zֵ�ks���qX;�gu���⭦i)ٺ;<j���k%���t�-���O���Y$ηlg^k���lK��T�v;����8�ucnZ��Ύ���$l���@ݹu�md��A��Y��>y%�1������	�p�;�R���p�v�J�dg{[����A	��p�Z�ɧ
tu��-+c;	f����=���6 S��\.v��צ�q�a�-6�C���z�:n�s��xt6ýE�����:��P�RH��"~$��}b�>�u��ԕ$��˓o�	�i���v)2B"8�z�ZoY�{;�=޺��I/�������в<qfH�voX��|`I���#Lǧ$����8�I�����,�o�z��Z`{�4�iRUw�7�	�N�{ �I$��o]Zz�ZoY�>]�� 
�3ď����I$[E=�]i�n��]�2q���f�uv�I�*^��3����U@�K*�A�f�I���� ���>�ꞁo]Z^�*��h�˭k.�Z7$������
���� H/�S{�}��nI�w�7$�uՠr�U�9�09�M�^��	�4�I*���Z`7z����NLY>Hю"8��z�Z{�� �'Xm*T��ɧ5zq>.�]���U�z��F����ٻ߀������~H�`� 5�<M���mCn�v�P�l-ݎˣ\��˯.Zez���F�YZ}l�>�ꞁ}�W�T�W�I���f����kP�5����$�>�z�]Z{�� ��7�_Y��՟��G&7�RH����kL�F��T��*(_]�T	$�[)*A�,�#
@R@��)!��;��	~�� ŗw��l�$f$O��UP{�߼,��}��}δz���
��:�y"�;���`K̜`m%U^��9���03w�Y'�ԣA�e��m�2cE'��E3����;q��"�<��f����˨�g��Ι�I�=�u��/�ՠ}/�/�����-��kR(dP��I0'�i�I%vzMi��kL�$.�
�����,[��H`��d�w|�fF���RJ�9���`~��4��B��1����#�@��V��:��I����ɱC�X��8�j��H#��Py����ܒ~���	�s#����֏@��V�����/uՠw-s#c�a�B|��F8up�6�[��e�<YP�\��9/3�f����UU���6�B4`�G!xI�~�Ő�24����ג`����s�ӗ��:_{���24�*UUWfɭ0=w������*�fJ�F�D7�G�0&di������RW{��0=&��>��*��#�@����:���4��24�U*IR��~L	&���Ƞ���@��V���uh��Y'���M�!UYˋc��I I��Ѻ[7�Y���W��l����;7ne.�:���u헱E���q���[=8yr��ۭ3�.�7b<Pt��+n�ۓvwc�h��.QN���l�wM�fgc���!ٍ�I͍��y�2h��Fʼ�p�!��ݳϊMI� 6�&�n�훞w6]vx��i��Z79��s=��<��e
�&���hIN^�f1.[tj��De��fm��Xve&�f�d�Kd�ɹ��ѥ�ZN
Sp�:�3�v4��QZ�n����ߓfF��Hs�RJ��%IU{�?o���/返1�G�dn-�n���0=$i���i�RT��<n�oz.�(�2F�qh�����������@:۫@r�7���i����*�y2|��֘24���C�(��O6�i��I�s��,���	�~_���24�$�|P��j�Y%�+��l5n�z��:ݭ���-L�\"N�,��������I�"�:�ՠ}~��&F�%J���Z`j�ݾ�e�K��K�k4nI���3
���`zH�&F���I$�8n��mH��B47O@����V�����-�@��h��#2�F��I�2>��*J��n��`~���`}s%�&MZp�+Pƃ#���o]Z�RT��6���Z`Odi���I����o]5�۱�t'��%�O>b�j��r\�<�t�R"��2K�"j�]���B\�|`I���F�%I/�7f���<��ƣ�)$�c�-�V�}Ѧ��`K�/��J��\�j�wz⛅'f8�I��~�d��l�J��/�/\z���
�Utq$O����{��URT�n�{6���#VO�T�{�I�o}a��Q�:0%̗�ꪥJn���7&���; �VT�Rf0$Q�	�&f:Wgs�6;Qۛ�cv�!�x|p�#]�a���������#Ǡu�V�}�V���~_>!C?/�����)|]�!u"�ģ�����&v	s%�#OiU%W���O�`�<p̑h�����@��V�}�V�x�+�dQ�ԍ7!��$�K??��=���h�tܟ  ��?�D�w��ܒ�L��n&J	$�'d����$�@P }�~_�wF�������S��r�r�kv؋Z�͝5\-kr"�S��\�q<\��t�`�t�w�o�������v	y�����R��f�LXjՍnF�x�#mȴ^��.{�=�#L	��RT�RIU.p�7w���!Hd�����c�;���/uՠz���޷�E#OF9�C�ʥT�ɻ�`nMi��;�����p)vP�ԊC
R$���Y'�UP����RS�������d�0?*I%����|�ߪ���A��D�5�)Pms�xr=��v�㋔���v��{[UҾ5��w`{��A����:�a�ς��.Ŝ	�q���;g��N*�-*\K�qgb�u���k"�����8�0pv��y֎���mɥ\��T�ۃ�]�㱱��&�zK�±��qKz��x;5��*�P^�=�ue�p�� �W���n��teK�����.�ETW��Gns�N��W���K�j���c�����U�\�5��t6N-���W~�ߟ����K�2F�U$�}a��� �����LjG���.[q��I/��]֘��0=���URW`�E�sWo�"s2)$�c�:���@��V��n= �ٜ�Zyɒ'$�-zF���0%�/�6�UW�w������bkfF<d���Z��h-��z�Z�����7Aę�q�q�S�)nx�)��H�v�+�"�CO����Z!�m3�(!�ma,D"B�8I�}�������uh���>�Ն�=��.h���'���������UIv���L	't`K̋��J��3Q��3s �I�&8�����޲�~J�]�ɫ��֘�R��p���28�z�h;�z�[�C�%�������$����~�8iX��:0%�E���n��d֘�v����\d_���H���=oE?��O�G>��n�.�Y#8n��-l��KI����r�u;Q2cQɎ'�:�j�/uՠ{Ϯh=jz.ỵM�2"��"�/di�+�*\᳛���~����H�/U���c$��"�;�\�.^���HQ�D!@�FeHV#VcIYIY|��I�$$#
1�2! Ȗ#!���!�L$#7�`^f�\)3F^sZ~�n���5���vu���,˛yN�f"Dc��AR�a�&`��n�����C��H�B7]0�K���XuA�
�YM	w$H�rSY�da�2�\��)��!l��k}�<���u�ow^=4�ݸVZd	L��1!	"ŀrP��i���rw�އ�9����a�ѹ�S4��Fm��oyRB2s29H���J�-@�L&����Sp�����l��&n��z�]���6j$f�P��nSS6j��;EO�7�ܒ`g#ue�bB������
AA6"&)�S��Q�
|��=
�*�̒]�$�wX�Ntp��e��
��?�W� ��d�����$�uՠwt��޵c�&`���$\`}�4��U�7��'t`K����?���
�Ź���M\۞��GY+�\��<)�u�\nVC]��g�Q���&F����E�UK�Oߵh��b����������t�\ȸ���4��#Oj��4�^�ӊFb��̒f��?_��}n�޺�y�� �rm�#	&5���6�W���07f������z��T$�  3 P �;�;$�ִtL'
�d�A��o]Z�>��\�S�3��,���+Y�����I$�L0�7Z�<��.A�����hs��eN��%n���ܷ���[�֎IrE�;/��\�S�>���޺��P�������;���q�*�=�Z`n�i��{��;֬odx8B47O@��0$��5$��y7�������k��au"�A���U@P_}�`�O����.^��$�^�����Q�Mǘ8"�>�����z{��޺���3(l�I" �ܐ$̌#�O;PuA\���RmȉV��s\;=>�gr<9Cxz�:�yjν�;v筠��N���S��n�xF��<vp>�J<쪃#�<r\p�Ԇ�V�{(�j�v�t��+n:&�3�}�-��	�v7om��[��k*�є"9�Bx�[�3!��/9�lv�vo8�{sr�m[�x���]��jVP�����'��Al�-��ɏ\���mT��g<6[;]�����n<n�e��W5��u4�]�����^5�ܙ���m���{#L	24���N0f.rt�5"dƣ������@����v�O.��U� �����.�S����z���i��̜g�%w��W��Z^�Oő5����Z�>+�6oy5q����{#L��eX�ŉƈqǠ\���?|�����}�_ڴ�z�ۙ|��
un�fn4��V��q���M#�"�����(�5��y#CqA��z����r.Ŋ��k3F���vn�n �A�xi�/^���ӌ̍0<�R�y9�b2<p���>��=h���|Y��ڴ�j�v'rFdMB)29�/�`fdi�=�������� �S�&H��2cQ�����V���|�[�~_���0	��>�����ڱ�
�]�	8�7,��ny��9�i�'nV�V�(�_���>����S��w�I�5��$� ����$��Mi��*����k"k	#qȴ�mz}i�`Odi�J���`��_W-w��x�@?w���;���3/���>��}jm�m��Lk�$&����I�&�֘\��?�$�W{��X��,P$ȤYZ�]Zܶ� ���w]Z�c�$k9�f�9��wgm��v�۷kX��}��`L[]��˯.Z�5�P�BB۱"h(��G|��� ���3#L	�0e�K�e@�A"nGd���2���)#��X�O��X�Nk�W�PD��H�Hȗ��s��N�2n�����?*�Uw����?w���<�α����<�8�h�`fs%�	�����U/Ԩ�T��lFU���(~�������4�f��䑸�Zs��I^��߀��i�=������.ۃ��tiLsv�#�'�����8���7�f��1�-^�t�\[]�k}�ߟ��u�=���F��*K����W��co#�1�����]Z�]Z�vzC��J�.pȁox���q�1�h� w��h�����Q�<Y328���심	�0�UI^�ߓ ����,�Md�&f8h�U4{g$�
 JF�
ޚ�lt�I$\嫢�+f.}p.���q�!��c�ۃ�oXy,yGcF9���gFy�i���u�n�Z��s	h�#���|�&�,2���j���39���`-�V�� �ǥ��-�s���#��W���W���JkG�A�9�#�4.����K� ���B�D�Z��:y��U�E.�������n��	�싵�f	ۛMclq�.�i6y�J���K��)ٞMϛv�t#Pɰ=�N�I�r^g�b5}���I�'�5��>�����@��@��M �ꦁ�W�VA� ǒ'$}�`Odi�3;=�u�=#ORI,����i��[��H�r-���h�U4�uh�uh�	���r��a��*K�R����.�?Oߚ`_uՠ^�@�j̯V6I#o8�4�uh�uh����h��⿞�tQ��1��c�[9W׉�qrC�A��m��6�C�����>�}qn!"�����_ڴ�uh{�����ʋ1F�Px�cp���/[��@81>�!�ɝߍnI����@�[�@8�Ǆ�0�9�qh�E��4�ʕRUw2kL�֘Z���`�!�H�qM���K?~��&�֘H� �Ⱥ��x�$,� r) �N��ŒUU�UC�߿yx~�ˬ	�4��UW�{|ZWx�f�ŋ��H�8��1zV��u��h���mp,�	d�@�"��(H�#Q�0��}��$>ުh���;���.:�L�����z��E���U]�7Z`L�ց�n���56�Ǎ�qM	�����>��vn'�4Q �}J�-�_�%_>�����u�3YVA?��H6��;�uh�uh��M�n���Y1��œ��-�F��%_�*�~�˾w���=�������{Z�͛�уb�C�M�m�n n2zE�)��ӝ�q����7k�;#I�E�<qh��M��Zz�_�|��߿~ՠ�_�99�Ԓ�4�4�ɑ�I`2.�ԒI]�����x�D�7"�/��V������R�&�]`zMi�<d�|�r�]Wk��/��S��� �"�����UR�S���$����b�b0�r$�$]`}�`d��ّ��W�����l��7Z��^u��u�m�b[����gq�/i�e,6��eV�!3m=]`}�`L����֤��77WX�~ٓ1?�qH������>�F��XfF��WfŢ�Vw�Ww�#s8�[�V�^�M�uՠ^�b�'ǆ�G	��Dc���U@%��]`{&���#L?%W��`ȵbqG�dxԒ�4��@�n��di�L�u�I_��%W�IAu*��F�9�p�#��M�5�͎$D̪c��\.30����B��q����7R�y�[H1sN&�A��p"F���	#�$'2�A�R"r�#,?K�����!I�ޱ��B .��a`��)�O�I$�lHH        ��vh   �-�j�m�d^�b�֌�.�g�m�Vh66��=��g���&��˺R�+=�2��]�ݺ�)��(�n�q�n-�ìnN�9�.�=��c��\X��J� n�t�v�#��8��m&�h�&^˖���Oc�z�e�[0��E��ݍ��E.K���Ne�z3�v��8��w�g���4��t��vWm�Ʒls��h�g��6�x�n�<�p���Ya��y��y�����ϋ��Ŏ��+c. 6��`4�aɋ�Ł]�xܰ�h3&3�&L�m��N�'V�eA��T(r��x���6g]��K�%��N$��]�:�1�d��s�����y;�8u���ˎgh
r��J�K�v�\\::�9g-�K]<q�s<�`�m��k  �+�A�#�`]��g��w&��=��A�k��UݺU�8�R 6�h�]��wL��;X�=	Ԛ�ٵӶWI0c�;u�Mۜ�.��$y��=mv�vt��s��]��-Xv4:6�e�SB��s����J�;�4�л������!�9�%���kv%�et�9l�s:c��%�]��	�o��D��ص�K���&䳛I2�	�i[g�9����n;�fp��;k
�m�(n�z8��e�n�6�Rv^���d)�&��< 1r�`��6��+�9�5N��Y�f:���vA�h�<Y*����lʪh���p��<❛�f�1�� �h�O7m��t��nC�*�v
�6���u�۝��Ԁ��]�Ȃ{6���8���{^8cM3%2��4�:��9a4ĶM7K�`R$�]�[�Tj����Qv��D����WM��FT4mi�^�:ۅ�&�m	FrqN��izUnuIX'l���ݪ�U�v�8{)��m�l 6PrE����N6�X�ڃ�EŦ�5�	-���S�@����:�z�5��\6�AΡU�[ -�^
��S���^X�꧒�_�҂
�LTz:8�?DX�����|�7��N�~ꪸj�����y�N���r!��ui]�]�>6�˹����6\[�p��E���5��#�����S�6�Z�M�2s�f����*S2�ۃ��gnx{k��e��w;:{pAp���\hR�*8gt�9Tt�K����u��bU��@n��C�n�w3%�=ko*<�avݺ�g/���c]��fU��k7K���붓��2�.�{����{�K8x�[lM�K�"�ŧ>J*�N#W8urm���P�=�i�����#L���3!�Ԓ�������~��n���(8�NAd����$���{#L	�4����f������:]���Z����>��������@��2�cRI���p$��>���d�0>�F�m+��N�2Dk������E�Š^�V���uh��9��I�k_EF(�)��,��yq�2gpC-�b⧎w%�Ok�M��13�����n+��ISn&�I��Y$��d��s_�T��7Z`5K��Ӝ+����u0	���*�%�J��z_�i���ՠ{�uh�r���H�RH9���4��#L{#LfC�,�n���ɍȜ�$Z�uh�]Z{�4��V�|u��=Ʊ��7��S��� ����H�d�0���r�:w�S�x��zv�R;���˟fz�1�#���k�$8���Ne�5�eW�LfC�zF��4���i���2�cRI�ِ#�h���[uh�����4w Yvc0Ɣ�r��S�F��1Ҫ_,BWH��JЂ���]RN��;�ˬ�F���8��s6JJ�q��O�߾�t0��bX����m9ı,O��p�r%�`+2'���ND�,K�:z�?�j\֋�5�6��bX�%�}�[ND�,K�w�6��bX�'���m9ı,N��p�r%�bX����rg�qλ5��k:�&����ܧV�(�랻g���+�*��ƾ�G^b�	����Kı>�}�iȖ%�b}���ӑ,K�������"X�%�~�a��h#C�߭��0\��=kZ6��bX�'��m9ı,N��p�r%�bX��{ƶ��bX�'��p�r%�bX��wԙ�k	��I�d�֍�"X�%���ND�,K���"X�"�C"dO�{��ӑ,K�����m9ı,O9���i�V]335�iȖ%�b^���r%�bX��}�iȖ%�b}�{�ӑ,K�^��Q<"`��=��.��F�4;y�1�&d�Lp�ӑ,K��{�ND�,K�{�6��bX�'��p�r%�bX����m9ı,O}����	�B˄5��Q˺���jr�NO1i�gv.��7��7���r�ƍ�j��kZ�K��iȖ%�b}�{�ӑ,K����ND�,K���"X�%��{�6��bX�'�z��9%���f\Ѵ�Kı=�{�ӑ,KĽ�kiȖ%�b{���"X�%����ND�*dK��?��Y��a5usFӑ,Kľ���"X�%��{�6��c��ș�����Kı?����iȖ!�[��E$r&$���h"� �ȟ����m9ı,N�{��ӑ,K����ND�,�dL���m9ı,O��g�5ul�kXf�Y�ND�,K�w�6��bX�'��p�r%�bX��{ƶ��bX�'��p�r%�bX���̓�ֵ�k]��t鱤T��y��0��s�|tr�6<˻v�ю��\�������N8B�c��|����3�7]����T��d�XV�9�z$�;�ӻ:3Ѻ�vW�j6�¿��|͞��;���v��v�e�P']��������]�E5�{��ǅ�x�Vu�9���ϊ�ad�[��N�l��,9��Y�4cK���=�^�wq�����@�9s�y'P4��]���9�,��/<2�z㣋=s�����^^�o8�;���Ou��=�{�����iȖ%�b_���m9ı,O{���Kı>����Kı<������Ւ�2�Z6��bX�%���kiȖ%�b{���"X�%�����"X�%��w�6��bX�#w���ȓd�J���h#A
'��p�r%�bX�}�p�r%�bX��}�iȖ%�b_�{ƶ��bX�'~��%Ֆ�kZ�K��iȖ%�b}�}�iȖ%�bw���"X�%�}��r%�bX��}�iȖ%�b{��k��-�fk-�ND�,K��m9ı,K��x�ӑ,K���ND�,K��ND�,C{������̘�e��j��K�K�s��+n�ban�&=g��(��*��Y�z(M�XMk34m9ı,K��x�ӑ,K���ND�,K��D�,K��m9ı,K�zx��kZ�֦֋��v��bX�'}�p�r�X��T����'�'����"X�%�����"X�%���{��r%�bX�>��<k5.��Z�f�Y�ND�,K��ND�,K��m9��,O�k�.ӑ,K���ND�,K�Mv���$մѬɬ֍�"X�%��w�6��bX�'��iȖ%�bw���"X�%�����"X�%��>'��f�[tK�5�ND�,K������Kı;���iȖ%�b}�}�iȖ%�b}���ӑ,K���[���L�.d�7��v3��p��r�tl:ރt�KiW׉�.�]�EI�z�]��t7{�[�ou�bw�{�ӑ,K�����ӑ,K�����"X�%��=���Kı=�do�)�.kZ�fh�r%�bX���p�r�G"dK����ND�,K�k���r%�bX��}�iȖ%�b{ǡ,�˜���f�\Ѵ�Kı?{���Kı?w]�v��c ҇�QѸ���w�6��bX�'��m9ı,J}=�z�+�a5��Ѵ�Kı?wޜ�r%�bX�w���Kı?w���Kı?w���Kı/����K�j�ц��fMm9ı,O��p�r%�bX���p�r%�bX���p�r%�bX���Nm9ı,O�zN�t�a�
ʘ�O�K��/T=K������Q�d�EA�}}���0O%'0�߯w�%�bX�{��6��bX�'���6��bX�'��ӛND�,K�{�ND�,K�Mz���$մѬ�\֍�"X�%�����! ��H���M&��	���͡"�'>��M����D�<�����kF[tK�3Z6��bX�'�����r%�bX���p�r%�bX���p�r%�bX���p�r%�b�����)�d��T2�a��h�?w���Kı?w���Kı?w���K��V$"�n%��~˴�Kı=���sF\�kZ��Ѵ�Kı?w���Kı;�}�iȖ%�b}�o�v��bX�'�w�6��bX�'�wy�Z�LִK7*�\�����h��`�ayΩ��v0����Y��n�"1��V�߭�7��bw���ӑ,K���߲�9ı,O��m9ı,O���m9ı,K���c�讵����ND�,K�k���r%�bX���p�r%�bX�����Kı;�{�ӑ,Dh#Aw�~
��8�n�a��%����ND�,K�{�6��bX�'{�p�r%�bX�w^�fӑ,��hp߭�����r4NH.�
%�bw�{�ӑ,K��}�ND�,K�����r%�bX�{���Kı=���)0�dՆ�fMkZ6��bX�'}�p�r%�bX�w^�fӑ,K���ND�,K�{�6���{��7������W���nr����Ǭ�ݳ]��=t�
i�i�pН�ʚ��͠M�����:_,��s�h�8r$�h�v]v8�d^�B��!�s��C�P����g	$;�fzz��G\ c��wbzT�-�)��0�v���윊�Ѣ��v�`�nU�k�@�y��ۄ�:����ڎѻo.WWg�+"G9t�m��6����0�f�[�����D�� n��Sr]e����d�\n]��Ev�\ q��Χ�A�D�[-P��ю�uV���~}ߩ��g�����fӑ,K���ND�,K�{�6��bX�'}�p�r%�eh{y��-�$��Zq����4,K���m9ı,N��p�r%�bX��}�iȖ%�b}�{ٛND�,K����)t\�浪K�6��bX�'~��m9ı,N����K� R"w�����r%�bX�����"X�%��z0�.fr��k2捧"X�%��w�6��bX�'{�{3iȖ%�bw���"X�%��w�6��bX�%�����讵�շZ6��bX�'{�{3iȖ%�a������O�,K�����m9ı,N����Kı?zh�Z��ܚ����K��{�*�B��Ga���8�%P��+�ki��b�nz�JO�߭�7���'}�p�r%�bX��wٴ�Kı;���ӑ,K��}�e�r%�bSC�~���G��q9 �h#A's��m9��� �;���&{���Kı?w��]�"X�%��w�6���&TȖ'�N��d�\�j�F�$�k6��bX�'����iȖ%�bw�߲�9ı,N����Kı;��iȖ%�b^��_g�I���Is5�h�r%�bX���ND�,K��m9ı,N���r%�bX��}�iȖ%�b~�l��R6�q�n5t0�F�4��w�-9ı,N���r%�bX��}�iȖ%�bw���6��bX�'��|����
����@�aۧ���A^.��M����u��q�$�ӝ�����9ı,N���r%�bX��}�iȖ%�bw�߲�9ı,N����Kı=�FY�e�q35�ֵ��r%�bX��}�iȖ%�bw�o�v��bX�'}�p�r%�bX��{ٴ�Kı/�_\��Eu�&��Ѵ�Kı;���ND�,K��m9�!��@� �ƬjJ��ƌ(���(Q���%���9�����\1�ė	�,�Ip�0]l��|�'��)���� P	u{� З^ �<Ā��%T`�J�SD�)�\�d�/6s����~�˪�)$���!$�$�C)����3W�k)tCC�&�5HP!U�X`�#FeIVRW�s���Ŀ0u�U4S��Sp��ގp�5��˦��i�UI��_�z�K�x��K�����P�y��m�8�J$*�bP" 7Ά�WC=�P�.�r�]Ћs�w����v=�}�m,�����cr�8��K�a�QL�
�)W^K�ٶ�)�ʤ�������JB�Rf���,���kD.�h�	V��0�i��%�.S�� i����!�7F��K�"��	�Gt��`�7�L�!�#!�Zi3��L.Ml7����a�Fp��0]6�� ؎�� �A�M ��W��W���؛��}����Kı>��iȖ%�b_���YAC�1$H���A�F�{���Kı;���iȖ%�bw�{�ӑ,K���߲�9ı,O���EQ�!���Ch#A�{ٴ�Kı;���ӑ,K���߲�9ı,N����Kı������~0�CFG	ep��[��Ǜ�ݷA�m�n�
��<JN�,����0�j�F�$��q?D�,K�����Kı;���ND�,K��l?�	�&D�,Og���m9ı,K��Կ?�ц2Sq�.��F�4;g�fm9ı,N����Kı;���iȖ%�bw���"X�%������Zˆ�Rۓ.k3iȖ%�bw���"X�%�����ND�,K���m9ı,N��{3iȖ%�b~�M�Hh��j�sFӑ,K?�`dOk��ٴ�Kı?����m9ı,N�^�fӑ,K�DB� � :�K�����Kı?FY�!�^&f���k6��bX�'��p�r%�bX*��������ı,O����ND�,K���6��bX�'~����/e�V���c�X;%�϶'p�n6��xٺ�=�ي�ք�)�"�.ѷ3�vӑ,K��u�fm9ı,O{���Kı;��iȖ%�b{���"X�%�~�f{!K��5�kFk5���Kı=�{�ӑ,K��{�ͧ"X�%��{�6��bX�'{��n�a��h#CF��j8�.CK3Fӑ,K��}�fӑ,K���ND�,K�����r%�bX����iȖ%�b{'�/�q�ua�Y�k5�ND�,K���m9ı,O�׽���Kı;���ӑ,K��}�fӑ,Kľ<J[�e���.kY�ND�,K�u�fm9ı,N����Kı/~ﵴ�Kı;���ӑ,K�������!D�3"�U,ȰH�F"@�$ ��#�����D�E$b0����ڪ�r���2sI��my��<i����m�=�3��4V�-�a�v��e����cL��rl(�P�[#����Kn�ٷmA�M��sȩ�l�����%n��gZ�ۣ9�ƍ�7i^�W�ϒ��`�,A�R�'���4b��uhf�� ���2�엎:KGB��.���Ǝ����<��2��&ٞ�	;�j琼��v����{g����mL��t�:�\�:�8����٬'e�:쥆�ݶ��jT�p�lϓ�,K������"X�%�{�}��"X�%��w�6��bX�'����r%�bX��#�~�4e��֩5�6��bX�%���[ND�,K��m9ı,O��}���Kı=���ӑ,K��}y��fkZ��kiȖ%�bw���"X�%����6��bX�'���m9ı,K���[ND�,K����$�2h�k�u�6��bX�'�k���r%�bX�w���Kı?g��m9ı,O��p�r%�bX����)u5f�a�h�kY�ND�,K���6��bX�'���ͧ"X�%��}�ND�,K���fm9ı,N�ס��3Y)�۔xan����a�m҄��v2�*�㮭�9z�;����'7DNkYE��w�{��7�����}�ND�,K���6��bX�'�k�����L�bX�����"X�%4?3߿Rh�c"�)�t0�F�4,O��p�r �QLwq,L���ͧ"X�%����ND�,K�}�fӑ,KĿ%-���X�$���h�r%�bX����3iȖ%�b}�{�ӑ,�"}���m9ı,N����ӑ,K�������q��e2ԍ�4���4;�߼.�,K��;���r%�bX�w���Kı?{]�fӑ,K�����&���j�sFӑ,K���{ٴ�Kı>��iȖ%�b}���v��bX�'���m9ı,O���z:�z.�r:�Q�eϜ�fѝl�`��*ƳG�^��g33�����Z��w�x�,K���6��bX�'����iȖ%�b}�{���~��,K����m9ı,K��2���&����[u�iȖ%�b}���v���1ș�����6��bX�'�����r%�bX�w���O�"X����?�RSF�ц��3Z˴�Kı>����"X�%��>��iȖ8"�3������p�r%�bX������9ı��+e�
�"�(ƛ��a��hX���{6��bX�'��m9ı,O���.ӑ,K���{�ӑ,K��߾,&Hf2 ��\��a��R�����"X�%����e�r%�bX���p�r%�bX���{6��bSA�U=���f2M��E��`��7[��]�eI.8l>+��4�Xrk=uvlb��8���&DD��e�F�4;�����Ȗ%�b~��iȖ%�b~Ͻ��r%�bX�w���Kı?zBx�ж�qˎ5t0�F�4��������ș��;���ND�,K����"X�%����e�r'�TȖ'}#�ư�,,ֵl�Ѵ�Kı>��fӑ,K�����"X�%����e�r%�bX���p�r%�bX��.R�35�ZֳiȖ%��*2'{���ӑ,K������iȖ%�b}�{�ӑ,K|~!D�,0��H�D�RL�H� $!1ڒF�bBU%$��V@1�!�C��A��P�
T��L@�����6��bX�%��̹���j�k՚�ND�,K�w~˴�Kı?{���Kı?}�z�9ı,N����Kı=��3&\��V�{'�u4�w�������<�v@��F�[� ��]2'3��]ss�r�~�߽�7���'����6��bX�'���ͧ"X�%�߻�ND�,K�w~˴�Kı:w�fg��]Y�jY�s4m9ı,O�k޻ND�,K��m9ı,O���.ӑ,K���{�ӑ,K��O�����h�L�]j�9ı,N����Kı>���ͧ"X���C"dO����m9ı,O���ٴ�Kı/O�{��T�[e̹�ND�,K�k���r%�bX���p�r%�bX����m9ı,N����Kı?zBz˳�i�Y�3&]k3iȖ%�b~���iȖ%�b~����Kı;���ӑ,K����6��bX�'���b����34���kp�lcj���ftgY��&�n�h5���דSIh:��YN����ۤ�qDp�^2�v�nu�뗇o��}�v�4�ղ�N�Rҫr�^,<���5���2�:E��i̞w1�s�;�=aݵ��F�l���n:������s��Ɠ
�s�<�&�kE�&ٹ]nlֳ���	{�n^Oi�D�뇻2��7Oi����Έ�*�����w^�������>��\;Z�q\Q�+b�{;���q���1��v;�gI�MY$�7[���N�{�ı,O}��6��bX�'{�p�r%�bX�{]�fӑ,K���{�ӑ,K��}x�nK��֌�Ѵ�Kı;���ӑ,K����6��bX�'�{�6��bX�'��ND�,K�ݹ�Io�����5usFӑ,KĿ{޺�r%�bX���p�r%�bX���p�r%�bX��}�iȖ%�b_z��2�Mɣf�5���r%�bX���p�r%�bX���p�r%�bX��}�iȖ%�b_��)t0�F�4�þV���FHQ�7�iȖ%�b~��iȖ%�bw���"X�%�}�{5��Kı?{���Kı;���L�L��f���3;v�4��qv0v�e�7n�����M�F�N�B�Ӗ���~����{���m9ı,K�{٭�"X�%�����"X�%���ND�,K��-�ɞզj�.��m9ı,K�{٭�!⢅r&D�?{��ӑ,K�����iȖ%�bw���"�eL�b}�[.��i�Y�3���ӑ,K������ND�,K�{�6��bX�'{�p�r%�bX����[ND�,K�;&���̖]kT�5��Kı=���iȖ%�bw���"X�%�{�{5��Kı?{��ӑ,K���$%�,�8�5��4m9ı,N����Kı/���[ND�,K���m9ı,O{���Kı;�}�5��h��V�����Y�g��rkˏ"�Q�n%�Ta݈T�Bu���7}��oq����=�f���bX�'�{��r%�bX��}�a� �$����M�$}��ffYMF�5�֮k5�$D�{�&�z%�b{���"X�%����6��bX�%���kiȖ%�bt���M\��ZԳR�kiȖ%�b{���"X�%����6��c�mE⁆�n%���kiȖ%�bw�{�ӑ,K��N���ֲ�ѭL�ִm9ı,N��p�r%�bX��{٭�"X�%�����"X�%��w�6��bX�%����˞զj�.��m9ı,K����ӑ,K�����ӑ,K����ND�,K�w�6��bY�7�������!��#W<���t�gf0Zy��m�t��!F�Y��=Q��1��j��.k5��Kı?{���Kı=���ӑ,K�����"X�%�~ｚ�r%�bX�}!�7�L&d-�֩5�6��bX�'}�p�r%�bX�����Kı/���[ND�,K�w�6��bX�'}�!/��2�35��4m9ı,N��p�r%�bX��{٭�"X�%�����"X�%��w�6��bX�%�s2�}��][�5usFӑ,KĿ{��m9ı,O��m9ı,O{���K��E? ȣ�A���F# b�H�!������ӑ,Kľ����̲�.�k5�\�kiȖ%�b~�}�iȖ%�b{���"X�%�߻�ND�,K��{5��Kı>��;�պ�2I�f�t��g��ݯno�gD=��ٝ6#)�]0-��V���vg�cX��~����{����m9ı,N��p�r%�bX��{٭�"X�%�����"X�%��;�%$՚ˣ533ZѴ�Kı;�}�iȖ%�b_��f���bX�'�w�6��bX�'��p�r%�bX���/����֬��.kFӑ,KĿ{��m9ı,O��m9ı,O{���Kı;�}�iȖ%�b~�C��ru��e�2�[ND�,K���ND�,K��m9ı,N��p�r%�bX��{٭�"X�%�����ԦfR[�j�Y�iȖ%�b{���"X�%�߻�ND�,K��{5��Kı?{���Kı:}��~e�%ȑ$%��	\a�A	rRR��`f��C1� �� N����ǹ9���=�p��8�VYh��9�3>YP� BR���9�c�P��@������&c3\K��D(D���.:	@�1��J�2V��"j-��.���]\!!i�H����aJL��4�e�k	L�p!!$�$����:�*K���5u���$`�!.2�E����P",Q �V*�H�D �R��] �]d*�����I�@ˁ�R�E��f�Z�!K��q�iTӠd�њ���#�u���z�ҽ�ߏ���� �-� $      ݳn�m-�    -��mH�Mo1u��5�:E$i ��js��%�qL�&h`��`y���H��dz4���������c����ֻ����.]�Px�
[����mu9�q�p��l����F�xڧ�xޤ�(�r�z���V.۳�Ʈf{�bs���8��yp�۞��;{�8��tN��L�s��=�5h��8���Ӻxm��r|���;�F�.65��oH�됝�Å�;���':�/�.9�����q��9wMv�cM���� ���\[�����兟gQ.!�Y �v��a2�g;��Ut�VL=��ɷ<��1jLutnDZ�٩\��q�&7s�7N5q����ۭ��0];@S(Yi^Q��Q�I��{@67����sn���f�m�E @ ���l�&��E�i�f���_ �M���C�m�Z��÷W.���#>R�%0q�׃��r��<粆�һg����=r&��۹�݁|�uϥoIl\�8B����;=d���lv��ī���fy�1=onkɔv�v7�["籾�ն��/����fꧢ^M��˷53�v(�݋jj��\N�.f;Ej��<��9^���
J��tu����"�c����nAɆG3�@�yX卾>D�lʵ��n9����12յu��� ���\* mE�4��*���rV%VԽ��W[X�N9Cu�dKr�;p����mF�1D�m��a�%s��}w�L�iS\wc�F�r�	a�nbwv�,���jw:�vx��S2S+�7a�r��pP
hܙ�%R��rL]R3���{q3�:���Y,�ܾ��j�e�H�k�+cI���N�Y��A�	�p�t�&A9ݪ�V	�lvJ�iVU������f�&���h��kYŦ���[m�s��]�����ʴ�=����6�Na�;��U���lF��W�`�Mk2�Q�~6�� ?"QC� ~D� �*�Q��&�~ �c��kZփ�q�I򶫬���N��U�ٵ�,@��L��xM潢��n(� ���8�=r=���l+�5�'��;�	fܙL�r�b�ۣ�dP��]D��<�sn۸��pt[7i�w1�nӍ����v��u������v;:��]Nݭ6���	k��u�����v6�yen�;\����뷶]��*��q/@D�ݑ��[��������x��NU��`ռ��M�u���Ή�k�X�r:۹�j�I�ؒt�Inf��r����bX�'����"X�%�~����r%�bX���p�r%�bX�����Kı/}뙅/���r殮h�r%�bX����[ND�,K���ND�,K�{�6��bX�'~�m9�DC*dK�����St랚�o�߭�7��,O����iȖ%�b{�{�ӑ,�!�2'���ND�,K����5��Dh#A>0|�2��D̉���E�bX���p�r%�bX�����Kı/��f���bX�'�w�6��bX�'rt��)f��]���֍�"X�%�߻�ND�,K�@�{�5��ı,O����iȖ%�b~�}�iȖ%�b~�m�S��L���ֲ�m��vn۞u)ך���6�v��qzq�!�u�ūn�d�kc5�{�[�oq��K�w٭�"X�%�����"X�%�����"X�%�߻�ND�,K�HOKM�u5�[�ff�[ND�,K���NCbT��j%����ND�,K����"X�%�}��5��Kı>�C�w=d��Ku�Rk4m9ı,O��m9ı,N��p�r%�bX��{٭�"X�%�����"X�%��zHK�Ks8�3S.h�r%�bX�����Kı/���[ND�,K���ND�,�	�>���ND�,K�����K�j�3.j��ND�,K��{5��Kı?{���Kı?w���Kı;�}�iȖ%�b}٣��jܳ0�ȝz�D�_HƷ�Y^<��l���v����g�b5BP���랚�o�߭�7��b~�}�iȖ%�b~�}�iȖ%�bw���ӑ,Kľ���m9ı,N��=�g�Y�ɫ�Z��Ѵ�Kı?}�p�r%�bX�����Kı/��f���bX�'�{�6��bX�'rx����VY�S5��ND�,K��m9ı,K��٭�"X���"��@�W��O��p�r%�bX���iȖ%�b^����\��%�\֍�"X�()"g�����r%�bX�{��ӑ,K�����iȖ%�b{���"X�%���'���j��5��m9ı,O{���Kİ�U�����m?D�,K����6��bX�%�}�.��F�45�_7�"&DN%!��x�`�ܝ���
7g��Ŭ�Ƹ+vv.,�K��h�ʝ�����������d��{�ӑ,K����ND�,K���kiȖ%�b{���"X�%��}!�浬�ԙ�6��bX�'��p�r�șĿ���٭�"X�%�����ND�,K���ND�,K�޳2��:��\��u�6��bX�%����ӑ,K����ND�,K���ND�,K��m9�q�������"��1���o�߭�e_ꤩW?~��&~��0$��RJ�+()����[�p�0�$�ՙ$�<��ho]Z�uh�\�-�@��?�Q��&E35�2�������z܇n��E������p�a��s��$�"�-�@-��o]Z��V�r�eY���@fI�@$�ν��Wf��Ll֘H��"�F�~2I��q�4mՠ_ui�J���wZ`f��,��%���Fd��-����uh[\�-�V�.6H��p�@��L$��I`OH�RJ�frp6��{M�)��l��Km�#�cC�մ'r[I�c\x��n룆�hN]��v�>�8�a�4U��9�ΒҖ�^ 6f �!\YNa��u� ݯm�"�n��셰�v�1nz�5)�w��p�����杺	������Y�5�%.��2mG��b��u�;��f�giz-�Ǯ��x4�l ]vYV�,m�4�.����o¥�Ò���ld�َ��ɶ��ی&\z�n����zɫ���(p^�Dm-߭���������-�@�n� �g\90̐�I$s@�n��Y��������V�z�s@��\�ʳ#����@����`�9��`e�Hr�&f&��I�z�Z�������uh+�30x_�a�$�@=2s�	�4�����`�x��vK�m6��oO5��[nn�#ۮ�;zv����'e�:�sjtݶ����T������̍03$i�}�/��.����@�$@��ww�_��<��X�[�@�n��/�y�bY�����#L�I}`L���#L�a�3_����#qh�uɠ^�V���@�n� �θ�xfHG!$ɠ^�V���@�uՠ}�&�G�����>Wp�UF�n�m��،G`�p"��q�V�z�j��n�\��̱��$�w�Y'۽b�'=�� �;���,��������p8�R@��di�}���#LfF�)g<�ǅI��Z��rhz�ZEI)I*���s�'�03�`f%�X�9"Q��R���^��d���Œ}�uh�uɠ{���b�hy$�gz�̍0=�`{%���H��O����6��a��[
ջ"	Þg4�+�E�mӥF�׷�=�J�����}�N�uP�i80���X�I�o)d����Uf[�V�_�y������nG�- ����#LfF�̍0K��Y��JB`�C$R�9��,��ޱg�_3:�ڴ�d�*�U���7I�H�w]Z��� ��4��	�!�aB����	c�U�Z�b�P~��I�w�Ɍ$ʁ��&�#L��ΰ>�`fdi��*?�����U͑���ݶ1���2�<;;�Y'�=m�y�<���]_�ww��~�� 	�|qA���-��s@����;���=�uh�\��$��i�hzF��`fdi�{�s��]���ocjT����{��I�ޱg�P��;�~s@��ߵh�U�]��K2C�ΦfF��Nu����{#L��f,�##M��Z׫���V�}�V���@�Ř��I$�A��;O{�s�!��)}<�H.�nC�Fp1Wj�g�����:�|�v��wA�͔۱ۍ��ml������1�X{�%I�E͈�v�l�y�.Wk�Y7O��4:�54����uea��:v��M�.J�q��:�g�iqn��&�bq��4t�����c�X�9\�G:Lf��l4Vn�����v��W5��&���LDO�7����&�x�-��]�?Ϟ���+�/O\����z�2a�lr�-��v-�����ߚ`Odi���� ɓ�`b�(�h�dyI�ȴ�%�%�^�� ��ΰ>�ʤ��ٶa�U�6�Nd��Z��V�_Z���ՠ}��Vc3�<r- ����di����=��(����D��qK$�oX�O¨P������@:�ɠ5}3���&LO1�K!8�F���%�&m<�)�s����r���v|ꬓ��"rH�,�����O����g�V�{�p�v����eيҙ s�L�F�)$Ҫ\�I����di�}�V�K0/��`�_��#M��Z�6���di�=��{#L2�.q933$���2ho]Z�]Z{�� ��M��~8�y&7"`Odi���� �%������a����ˎ8G�5lnX������-9�8�w;KD�uTu�M���Q��03�`�:��di�=����Xb�(�G��h�Y�}�uh�uhB�x�pS2G0����`}24��di��iЕ�t�V��(J��U!hJ���Y?klf~�K�B74�D���aBa��;�}�
��	�[�PI�Ԩ �$h^���A�?|JJ��q3-e1�t��f�h����:7�o�i�)B� BH��5��y���;6��>�����4�@�H$X!P��%	XЖ�G�����IJ-%`Aމwߎ�|}La��\�55�w��
h��(��1� ?	��$�&c�	2��J��F�0�b��3�3LI����i���0��C!����Д��CR�� J�Q �A � 4J �|xV1�8-�)���B4f�jR�(�o>���>�����٤�f��$R �)C�����? h�$f�II����5&�M�1���	#B�0�m���5�iC0ִ�������� mO��`D�X��$� !�UQ�|*�/��V�{����@u��2I9wΦ�R�lߓd֘{'XL�h�..�S2D��7���@;�f��۫@�z��;�w�f`�-on`��Ȅ q�y���\)�ƝɎ3���(7��b3#FL0x(�m̘���Y�}$i���֪���	&��6\�\�3	(�x��>�uho]Zw]VI;���� 
H����e��DF�R'��077Z`fdi�L���F���9c�̄r-��� ��nI���7!��"B�����!0���HJJ��(B�c
���IF���K-�*A�$B-����m�i6��#+�і�!)KIm�-aBXHFT!IIa!IIJZB3�2d��� �K��h��IR�*��َa� �,�fa,���7�g�������񑄆L��ȴ�Y�}���/�ՠwuՠ~��s5��1�ʴ�2�ts��U�+���n�����gn�S8�v�H�	��Cq��nL$�ﾱd�����Y�{���*��H��uh�uh�@�mՠ{�\]��d��7���V�^�4��Z�uh^���Q8�72c�@-�4��Z�uh�uh�:���HG#nM�V�o]Z��V�[�h���W���C�U��NRm:,F�[�.�����nz9�8T��`���kI���n9����2m�մ;=��mw]�!��7-�xf]�l��t�\����eiR���ܕ�8vEnp\���󷐄�R�ws��\�8t����B�[�۷I�\ݕۆʜ�츢��oX=�P\��M��q�'�:�nըo;������,EʯMx��F����ʗϊ`�^��hL ��&��vr�7um�s>R�v..��en�e���j������i��DF�R'$I���}b�>��� ��h}n��w"�"#q9�/��`{�`2u���i��#L��4�2d̙��"��f�����:�ՠ{�uh��y���3q��@��uhz��=�Y�w����$��qhz��>��� ��h}�V�}�m߄k�E���Ut�[����A���ƵMm֌f۰C�$�5	ȌP�q��N{zŒN�Y�}�]Zz�Zװ��R47n$�v���@V��\ ���b�=�uh}�V�uέ��30�"�F�z���`g�i���4�=2u��l��1���@�[�@�$����s��,��"�	@S���z�{#L�'X{#L�0=����1l���iH�la�x��r]a\��o+�S����3��-[Y-Y��|�S ������=#L�����1�T&7����>����n���@=z���e@bɒI��:��`{�4ϕRMUH��A�#��!"����٠w�ՠw|�,�&D�8�Z�#Lޓ�zF��0�e��9���)�d��wK$�(W�+���/o���޷V��5k�����^��Ы����j�`��� m�PT��5�̑��������@��ՠ{���=�uh�l�*�țkU1���@��ՠ{���z٠{���ʅ$xwB��@�8QG �N��X��l�=�uh�����1;����s2$Z�[4z�Z��V�%� �"�$���:�w\7$����\m�7���=�uh�K߯��߿j��Y�\��n�Lb��d��9��k:�\������.�Rh/&�4��tI]Y��M�R�AE$�7�s��Y'��`�@��ՠw �,��K#��u0>�0�N�=�0>�=����1c��)�c�@;��{�uh}n��ՠ孧`����@����>��Z�[�@=�Bt{�-��<�8܉��s��,���� ��u��di�*���J�B������ʪ�nr�����,ki+��q4kIf+��tX��e;f�C�ȷb��]�zݹN���.�ay��;r���]�o=q�a�q{v�����G��<� �x�$�K�ya�-Ӄbֹ�\Ʀs��ݍv�{/2ov�wg�]�=�R[�zf�m�[3�b�/.�F�Wpu��C��73�<\�j�(��w[tgmc-+.aZ5t2��#�l7����}���>�[<Ɋws��[�<�\#ֻx�q�sڜ�V�����,�=��Z�����m�7cL�������F�C�.�����d̒- ��4{������ՠZ�Ǎ�X��	#���=�0'�4���4�'�u�0(�՗�I#���/���>��Z}�h�]Zr((� ȖG�Z�H� �������F��$�j��B��=N6ȗl��w�ڲv�^7��X:�n�vf꼚Ì�V��sNq�l���I'�u��di�=���UI}a��i�I|�0(���#��%�}��*��T-)cȅ�HB�
�jwwf�;����@��v����#q��`Odi���i�Od�����a�L�q<q9��E�}������=��+P�po������Od�ޑ��F��0���r�vK�{PCn۔9�a�3��3�&��}�E��ݧ�,�6gM۶��nk�9�M޷V�}�V��[�@/���>"�32H�z�Z}�h����+�;&&D�$Ü�`{�4�3�:ƩRT��$���$�U�T���Ld�0��V�S�BF��1Š�f��[�@��@��ՠ�kra� E���n��F��0	�`z��p����1&^ݓ�-��n�����3v3�<�ű@�xsfpcWQN�f��/R���m�?�ϻ@��uh�Y�{�uh�Ó��DI��Z�[�@/����@��@:��ԙ��s#�H���X�F��`}�`IG"��9�Iq�$�~���Y'��Y'=�bɱUT]��d��4yDy�P�#/�L	�0>�F��N�>�F��O����6��a�Mɨ�ݸˮB�"t��u�V����{<,&&�ת��w��s����4�'�u���5��*��r�ՠ�f,`�(�7n- ��7R�����rkL����s�Qc�8����@���@/�����k1<�#n<rE�Odi���4�'�u���4�Ŝ\��!QB���9��I��UP��k����F��s��7$�UU� TU�E_��\�QEW��E_�UU� TU� ��	E�FEDD�"?� TU�UU�TQU� TUj����TQU��QEW��E_�UU�TQU��QEW�*�*��E_��PVI��lo� \���@���Y�d���&?�2�ԀP[H  �   �	R�E$� T����w@ ��@����Mh�W@m�`�
�Ȣ�3@i��eu����ɋ��E�3W&����:I�:��[c^Y ��9@ 30�kMi�Z9��5��{z�pq^�`	�����t�"���)֍N� P�5V.�
(�P�Т�1B��Z�P���RT���t�Ma�e�(@��p�d  �ò�ѧM
;Mi�Z7��	�j�jh�D�'�h�b ����H2i��IJP�0A�i���S��I����4��i�4���2����4 14ɦ���J�&�2<�њ�4�C��"B�*      ����-�N���ӻ-,�l���e���H�g�*G9	A|�3*�8�
��������1�CDaQ6�@A�U�"� �H�3�A�A�����TAd;<g�-?��.#��M���&��a�|�A\��9r���
޷��,;�NB���[�wF��K��S�%3C�a���s�ԓ6y"S�K�a
H^hَH�[���pH4^�\7��)�x�T�h-��RنQ�B�`h6lǙ��Bu��
��t��4���Q�۝�Y䳬:R��)�	J�8�۩{�z�W�9�wF��c��rAH$�c���L&����Ľwtx�����(���'n�4J����kn�)����Zn�{�7�{ I�o#V��	�5֪Y�<�3W;�XHM^h/0�91�e���Q���f�j�E��Y�'�뮒j�4u�E��	S]uu�n��*�ʍjʎ�]]0�4�W*�|�
		���I�C.�w�Y�������fd��WZ�"��@9�h:*����UL��$4n�0����5��-�P��)�U%����*�� ��qT����zS�ܻ�e!����ĩtb�j,���j_I��s\ՙ++Y�@0��R�@��,�f.��aE�&��@�*�(��Eќܹ��
�d��*�BV2��L�'p%��oU�[�j{D2�)��!��p(-�R�{����CSR�$7Õ�λ'e�DN�� %��*�1�)"ı�I�%[����
��wps�1tYFˢ����-�Y*��n�j�&]i�#&�f�.h��c&X`�4��H�7iY!�n�ᆎ7���s�yӡ�F$��[�¤6쐓������R���,agB3�Y˫�IMَ��E�&�wN�$	
"H�4Tp�L���T7k-��{N�20��FY杒Q!D�H0�QeLp�!&���DR2�D)��!��=�ï�,���[���<���T:.�ZB�,���+��b�0]h��Q�h:np��f�Cl��a}�,e>�N�ô*]�Ww#ldw�k ���UB����ȳ�mX�]�K;th�6JV��y�W�w�dI�T	F�vI fʰ���F�ѭ�a�\,��o|�8ʼtG|�s��8w,��*4d| �PY@B���F0!.�,�$!�e��H�S%/s	TIP�y�d+�I�oo�L��J�l��L���L�u��e�P�-9oU�ekVBeKe0m)%#	 P0��PF�B҃�c!�W3��"�1�;ތHS$c(��t�aE��ԝ;����6Ԑ�A�G���CP�F8�	c�+�x��9�i�FE(ц��B����zw�9�Ν+FHS���B+fs�Hى12�u
�+|�$�'H���'ugV��s]�9�ms/	Z7w�uW!*��T�S4U��R�W-ug:��
{]ݬ���ڡJ�tW`�f�R��eA����R�s;]�|K0>�,��J�ܔ,��+�BU�gi+����Gk�jN��������	��^�-�2�ݚbB�1 EfU���!6��HP�ݲJ,,�0R����4ʖc�aa.�ZM"`e���Dl!��"Kj��j0&�ӗD�*!,��\u$�*4J!�)n�ؒi��^����!�n��Q��*��$���s�
$�n�7� �����}��s��������                    �C�                         �=                                                                             A�                                                                        �bjE�u�-�ks6��[��xd�UP&,�t��5�ڶ��m&�a��P�ņMEUcK���:��e챀[Q�0��P@m�]e4Ţav��ˮA��s4����M�r˳Xn�-�mT-!E��E�:[R-��Q"퀺I�M��*����ܧR@���e3lm�gG]� �h ���ׯ@e�l�ݻd�LB�8�n]UjI; � 6ʹ��t�,�k�e�%HZ�j�Vm��h��.���h)���Z6��-��G.��]f�nA��kQ2u�Ȗ�+[v����� Z�V+vZh���#�<΀�gR��/�]�_^�7Y*a�&�Z;�u��m,.�h�v�j d�3H�6$i�U��`m��.HѶ�,��Û/�r�F�z�ACB:b�7K�^k�ق�ò2\R�Yt`
�[Gi��v��'Z�Ť���:/N���Im����8��H ]4�UU��[��Q �]Vmm����n�#R\Z������ж]Βk)�CE��º�c.[�����,(���c.dݛo��5fR�ah����@�[Z  +-M�Ao�����	z�K9�r� 9[[��m	a�4Se^�5Il��]t֜�$-�W�.U�[pY�	*'�:ô����:[n��EdV�U`M�����lj������� f��V��*i��H [B����t�5ͪt٠�v�`*�L۱��j�Mze��n�Y��l��9m#EY�Ҋ*�0$	BV�]l4�'�<�>cyJE�d�k�K�8�cZD4��mc��Ul,���5Ɍa��2���.i��[UU�m�    �iU���m����i�[x�p[M��i!�l�i��Y��N��:�޽5��a�   k��-ꓭ/���]�ٴ��׃;cLL;��&srKE�c�$��m�UV m�f�43�5�+�V�yA]����m�d��IJ.MW
%�;cXb�\�]H��;uʶ.k��-��Iw`.�S���+	��7)�	mՊjed�Du��c��ǅ�Kuˆ�^}x	��L�-��4]`��e�I,ti��cU������6��Im�6�ݒ]Z�t�-̀�[��Gnؕ���ј��.1Z��pp�C���IWSm�9�V�{6��m�H[G$Z�bO-�k%� �h6��kjF�l,$�6�Z�M�m�m�K"@�m�o6�u��D�BQ�Ph�p<vj[��j�j+�k ��F��.]R��ە�X ]R�CI{ZH ���6�嵢�R�D��]�-�6����,�P5�ط�[Hf� �M� � �`�4�l����m��  l������ϋ���UB�Qл:��	 8XlN�T��(���k�V��:�W8����j�p-6��u���Mn֗`{Z���#��V3`f�"R�e�ʁ&b��Ͱm�`� fffffd�����*?��(��;@�������!Ba@��_��(A���@�L�)-U��"(�ah�A��:��TK�[@ڣ��� ���i��h�����B8p�xQ�x ��4� ���<<jqMD�t�t6�"	#|�D�W� �<.��L�U���0 mqH�� �@��Cn���N1C `���ژ�� 4�"��< KTx'^	Դ�8������:�P�+�#Ah��R"! ƥ��|��Ǖǉ8 qV�)#C�_(@���# �B�a@���N'�z���|�C��JN�@�������\�CҀF�z�� Q�?
� �'�@�/�x�$P�Y�⪳333333 m�Hp   l              ��             ٍ�7]Cm�\�\m5��B;mf�t��`h�k-�Z����9Š.��Z�%�DŴ[�ֲ��K-��v����W"��j��+�(�]�]�Ku�jfN^�p�0��WS��pp-�L]��u����u�)��ưSF�R��x+3�Lҍ�-B��D��m,k����k6^�:�ظ�UChfR:��d�q,[�.�-�k5��FV�7fS�f-.�\M5��nts6�������as���Ƅ.R�K��	�B�Ke-r��X�Z#���ڌk���3�&���4���#P������M��y��%v2V͆Uv�E�'�� �P"$s 0�N��8!�'ʇ�>E��@�{�u�y�wy� �  lu��^����mԍf�����3lG0�f]rcR5�[�:��3ffV�6j��K���Fe�˝��=N�_< ����������/��~;�?W������m�v5ё	%����m�|;E�ݳ"�s��Z�2!�v̈�1��nծݳ1�"$������D&�YK�3�)�Y�ё��2jRڷô�i@Q�$�%.Ц 1Kh���Cw�s�\��6��{c�V�;G׾�I�|���GhȆ<Qڶ�ݙ��Y� ���m��7j�;�� �[k��Z��ן4����"�λ�j�ȃ�lȌ�P{^�'v���3�2#%A�i�fD{FD$�y�R�վ��!��dC��K��۫�C�"lT09��J�{��<�lȌ��7�&��n홈�Ǌ;V�۳"=��@����~��������=�Y���) X�k�G$�c�V���>�̈�>���m�uI��RѹЛ,
�5�ާ�ߎ����Cu�ܫv��hȄ��2y)m[��<��fD9+�M�C� +u�Y�Gh���$ݾݳ1�"	#����wK�N����'@      Z�%�֤�nm��f(A�H����5��snBm�nHЁzm����5�U�P�R6�qB�4�Px�r�:D�*��k���%�a��5nr�PN��w��>��K/tl�������:���;�:��wJ�Q��ّF�{z��\�fb;FDd�ڷn�2#�2!$���T�m���ɥ�dX�#p8�����ޣ�!�z̈r.Wn�n�����<*� B���D��"D���cBH��! I D�@s[���S��s�I7o�wl�GhȆ<Qڶ�ݏ ��r���e�Fʻm>����ّ���ѱ1l+In�5�v�
�Q��ّF�n�;��7v�(lG�wQݭ�[�m���@����%�vy)m[��<��fD9+�M�FD9�ّGF�.ﭦ*�^���J�]ث��кV�M��v�=�Y���Ȇ<Qڶ�ݙ��C(�_�=*��v���fDS�L+UFD{fD�F�4��:���YwU����(�w��~���Ϫ��r��W$j��i��Un�۶̈���I,�'��վ� E�{�wP�Wn�n��s��"2��oRM����3�2!�v���fD{FD$�Y%��	���5�      �e��b�l�b0`K�Sb�2��k���j��vmҰ0�+,��m�%ˁ�04q�i3kX�e���*��51E��Kt�"Ҷ-��i���7v̈:�:�V���>�̈�7+yW�����3�2#%Nջvّё	%�dԔuo�h������|���3��@���D��*�n��mёw�d�@��|�ؒn������VE���;�G�]�n�ّё	%�;�r��|;E�ݳ"�Φ��"��"2��#F��m���˶4�13v6c(Q��=�Y���Ȍ�m�m�� ��;���|Ua����K�?GZ�-x��D��	>6`���!�%1>3CH��4�fU����Ы=f�5�u4UQ�wR��@�¬���
2��T��٠C��:蚮��eQ�n�%�]=Z�;�(��m0��b�X�P]�Q#Æm�A�y���N;Lg
*HS(�I)���>��
+����N��� �A��X����?b�I����[�ѯW+�M�Gb�lȌ��ԓv�7v��~���O��z��Ϫ�A��Q�`�@�Bш�0�����W����wB}��;�뽻v���!��d^W*���V��������r�ʽ��٘������B�����mtz�v�� 뷾|��������Uk
a�ZKb��AU�.�ݤ��|2�8�ݳ"��ۦۣ"�lȄۛԓv�w;�&^N�ۻrs�I$���۴�_7vL(YP\���:�C_G�4Ȫ����   ��]K�昻�n�Y�k�-	��j���t��+�SSk��Il�\�h7떻V����<�&�s-�$�I�x���6��n;�7��B��ƿ}>�6K��U贷w;�%�Pv�v��d�<���V�y�ݑ��v����������W��[�m�ũu��7
1$ݿ{��{�@ݎ-�V������Y����w�v�?y����)Φ����Ir��z--���ȆI��wT���[�ںUM�N�XLӺ��nN�I#�Z�[��7vG��ۦۓ���4 #�
H��A����:�n�����e❵mݹ>w7ww ��\m��t��b�t����m� �g���߿|�|��Y���}�\��^�Kgy&e����������p�w%yW][���3� />�]��&�卞l�l��ʺ�h���g�'RMۓ�;�'�-�n܏�ff?_]�i��&f�s��j�|�3񎊩��I瓻�{Y@     �M$�7K�D����e�V	�-(9�F]
L��v�3c����J]���g$囬Y!�Ʋ]�YR�by|�����5��UKr���&t&��Z0��^~�����gjݷ'��wd���]unNrL��r��m�� ��wd���I�rw�fyԗ��wU��I�Í���nr�Q���L�Ƿ�v�rt�(�(D�(!$C�M�v�~��L�u�]N�5&e�{�pZRw�f^mNջnO��wd�U�Ϫ�b���dJ#vo�7t�qѷ��n�<���m�߉����z~{�I7ow��� n����ڶ��$��ww� �s׎��t� �wd�O~��[V�!f�S7��:>W
�n�n�H��v�E������ 9�ܫv��9��/%yW][�w{���`�k^�M��k�����U�s=�߇�޶�i����+�r�]݊B��B�Xj�6�M���7s?/�nܝ䙙�o���|�3e9�µ_�������W�kE���3��~���A����X��v2��eʰ�]_�ߙ�ujՋX��5]�(uWE<ą����Jb��Y�K� @�x�r�D�D(�� � �����%pΆJ
��!Z��0�#�ż�I�8�����	,�`47��H�0��,��!�P�3|�o�{���cL`BPʢ5QJ${+z��                                    'M��k�î��k��`[fe6�6֤M����!�Bjd.��-X�Z�+
422�蘌k��]�nږ4�u���j�Ѯv�S�n�ufnK��-��+LF����hY���a��jۋq�,�M1�rB0LJ������J%1I�!��4J��F�p�;f�l.+YB72��-�e�mPnNՄc���tm���^C�]�K���GG\;:�X�h�j�a-�K�p2��h&�iVX%��X���#��0�HR-cs�8�b���l��������v#]��5���:��r��nl*�6�Kh]�g:A��St���M�*j!&�R^j�U�^|�Q؁�����_� �t�� ���-�y����:      t�k�tMɋ֦N˖c�E��Q8�.��vƩ��a{:3Z��9-�� �(V���)�G8�����z'��rH��ly
�j�'t�j��[�v������W�uչ9�3/��ZnNs�	 ��=sz�n��y&g��nܝ䙚�S��۫���n��-��E�@s��|����?}�{��]Oy~�1��
�;糼�A3�ݵ��n������ڷm��I�<��X����>|��O~�zUW�� J�⭴�+*�n��'9'� �<��I�{�䙛��n��x�$��ǜ~���i����vOJs��j�|�3s�m�ڡ�\Y�bh�d��0�N�L�ͩڷm��I�}��]unNs��^8=t�L�g��4Q"'��D��;5$ݿo���n�B��m���J��J��tBш�6��ן>{����:��'��g��߽\�&��|�wd�_r�E�������$	�nU�ow�<��|��|<��>��&�X      u�z���^�Z��vx��4�ͥ���o�i�b��-9n�ӥ�j]�����i1v�u�.�fv�6nSF[�wwM��V��fR[ʭ5Ԍ/�;��u���~���Ђwy;�����w��x	��$ݽ����>�����xH n�wzI2I�^;�i��| 3��ѿw���	;�պv1ٖ�C5��N�4|�ƿ~�}��#��j�Z[�H#;�;� ��}^�n����$��^J�W][��{����N�_����3]R�6�v��j�l��Uզݯs�c��ow���<�ܴ����x���z&�>�IZ{��J$j���:�V�ۼ�엕�U�iI�;�"��%�ZIb�n���k�L��rw�h��*�V�t��vN�r]6��9���=sGU6� F�ww<H A:�8�-+v�{�3>�T���N�-%G�
`@ Z�;��|<@S���{HO����V�wA s��t ���贷{� �%�V������wvK�W�uչ4�{��<( �P �����l      'E!8�8�Z�I��S��Ќ�Ei�o#_. ;]�[vфw7M�P��]�v�5�dk�d�m��8M3�s��$���޽*��P��r`s���.��s��AO9�6��FwvO\[�Jݹ;�$�$���wm<$����� p�ޮ�&��i$�x[���UR�L�%L�&�a��������n��G>Չ�o�utQ"�|�\)�a*�Q��v{T��)}=S�/-���?(���7Qs�>�m�Q��$
���1Sm��CI�;��>u�}m�ګT���	a��u �?dǛ��}O�qΣ���7s�n��v}�yFD3�����Յ]M?G5S|7��,�m%�IVX~%0� @(�e=I�J��(�l�79X��K5���F�-!��+WP��,dZ�D��(J*�Jczւ�*8�cA�g�L��<_���!��|���h8������9cЈ�)�UE��Ý�?z��z���<E{PΣ���/=Sv���e��$���w�UT��,0�55�ݖ��v�\un���7	 x7Q��]6��q	�Z}ͱ�����4g2�������Z�4�͞7�a��Cw;m��N����$G�'�о�~UZF���!u3�	I�+���j�z�|C�ZH�"���z.��w�ȆP� ��bn���G:�&����Iuջ �!����/��_������'9��S�Q��n���Ͽ��Y@     o&[sK3�$�i?wo\��Bɱ���J�vT��[0�,B�M��J��{��n�fX���&
�HF-�_Ӥ��;�g�U�v�כ���5 �5�u���D���2~���7_֙@~��vҷo�E�I4&!����EI�[wvӳ��(�$�[�H����L+U��3Tw�xg{F��w^.X{�y 9�;�JJ�sͶ�J�j�Ф�hZb�;��Uv�4ݷ�"9�% BJyߪ��/-����A��	J�H���~Ty��9�s��_������@���|��U7l�@+hgQ�C�z�-+v�7QΡ(�=T)��m��1A��Kt��g���|<�5vwP���#��L+U���S�W�����W�z�Ꝍ$D��8 �C�ﳶ�m�{��Q�4
��Ic�vwP�+�wP�{m���m�tT���s�����G�BE�>%�>�EM�G�Z ��;��?\[�Jݾ	έ"�ё	9�iݵv0[�����*��}�ܔµ\;G��v��2 '9��m�����э+� uά���O�����u�y�K��|/� ؏�Boʖ:N��<���b/������kh��n��jD=ͱ����3�wP�Iy�;��K_Iﾤ� �@   D�$8N��뒶,�C\�.�kZ��H����-5��F���;gTi7��Z�I����Y��e*���t�<���f˼���m���腣?�$��>�|�uP�fs�ӻj�ȼ5�u	H�ܔµ\@>!��b�ܴ�l�Dc�{ˌIЧ�b��5�䪦�=�s�J1�6�n��WmSb�Um��]H����M��nN��O,�ƌ�ķ�|���c0n� J�|FE�@4�leջ`n��!�W���>�����|���Ch�H����wm]��>�����>�m����)���J�!����;Ư��j�6�|Cu�Wܴ��$^�Σ�Q�mg~�x����<�X�D�B! �	0|���;N�]����n��;�H��0/��tN��~���C��ʪ�0�X�!L�q�d��<(��t���w{���;i[��"���%�����^v�ڻ2#�>$ ��7Q����0�W 
�u�>s� ��Pʧ��TdC�| ���(}�u���*��&���hXI�m�a1m��m�	Σ+A��䯂�I��Z;Gu	�N�_���<�� W���\��n��Gu��L@yŹi[����u	@f!g�2�&ok�A��񁍡f�6oL*J�4�%b@b1��($�r���dl*SP(�Z5�d�4[헲����k�兗��4B24k(�BY3��t���:w�����y�=������   "A�                                 �&Ӕ�M�k�H�@��%f���IZ\�#v��¹�k���8V��b�I.M��X���e0�i�6T1��ښb�X�Y���+�0�Fk�sF�-vi�,�W{h�#R=t��$#�ZL+sk	G6��׮QcS��5�69�lB�ZX��3X���5��RѶ�esf�ѓXav��PŤU�Y����ǭΦr�f��	v@�W]�E��[��m�*��d�Ͳ8	Mh���t�ve�mfN��[0�]Fm-s��-�r0K�z�Y[)]3�
0��Z�cYvhb4�	��k���g)=p�
�**�M��v�T�԰�}��S�F���/��4p@�a��t>L �mW�����׫      	�!iQ]u���Ѭ��-V^`i�kU��HֵZ�K@űabi]2�)i����lL\M��V��[�v��UL�Z�c��V]L��W�֮�����@���@�E��~�zm0�W��$G1x�< +�_eZ�@{�w���ey���<@ݳ1��EH�J�X�;;�r���~$�>�{���.��42;����.����C�G1Ϭv�ߟ �Vv�"��)���~�Wۺ����9ՠChȄ~Z�]�vwQ��D�}��)�j�v�����FD-ׯ[m�y���t.�s��L�oH�x��<Y�<߱x6ۡ��#�FQ�W�s��\�Yo�N�����h	���r��|�+�9�{��y���[n��i9�;��?:ݾ��mU��mM��6]J��)�������n�Z	���j����C�wP�}C�W�S
�pm �� �#"��ZZl�7�{�?�)�Xf7Q��a�T��HŐp����>�,�����33�#�BP�w�K��۴�۴�P�o�&&svSo�t�+7���~����3}���|���(f!�#����;un�!�!��En�(�-�n��9�%$R!9���WguP!�����w|�t�{�M�     �e�5����4˓�V�v���6��uq*X���FSJ!e�n������,�$���ץ�e��E�M�����~�����j�H��2�)L����������'@�D$�$�F��NI�K�/��}ݺm����ui�3�W���<��6��BD_y�x6��4�����查��Ҫ�?ټ<���& ��a���wV큺�x�������5zZW��>��(_g�MǺ���Z�~�����ϼ�(��f#��ܦ���Ρ���:�r҂ꌈh;guFJ�s͂�Kr���e���*�mL�����2��BDrW��I��_�ޣ����)F�������u�{"�iV�e�L�Ė��/h�UA�#8�{ˌH� ���Źi[������ghȇ�B��USV�(3u�.�nMF#�Wm]��4�#��L+Uô_�Ť�*�ڵ�U�;�wQ�7��m���홈�}�� 0]�9+�u�vdC���>�����m�.��º�vh�k3�V%U�^��>|�g
 ��2��twP���� >��$����#�G�s����Wc�[��bM�Y�#�M�6q ތ�\|^���S���t�i���      C3u6sh��ؕc@�,(L�\�]��bf�u.-�.�:��1�ԕ���L�Fh k�Tְp.��C�O!犪��F͚�#��u`\�3[�}a�#��I�(��v���� hLGhȼI���+����yGu�_y����y�$CĐH����Vۣ��x�����6]���q��x�!�	S9�>$��Ѻ�u���?(�]��{������ّި������µ\;E�x�E{�ȃ���kB�;�w�ȇ� [G��/�|�9�ew�z߿⪵��v�]���^�:a_vwQ�߁ �#��]6���P�P�FD.}c�Vۣ"�>럫��-"v�EBJ�+-3M\��B�bz�^Cn�Ca�Ƣ��+���/4�n5N�FQ�m(�S!	!(��&�I4[�E��Yl
JeB�)A$P�BRH( A�H0dJX45(��B�����I��(�(�����1���^��|��H�i�tih�b���r�/�ԓv�> ���������̈}]�����>�m����B��n1vh!�X��*�_�m	�W�V����2#�o=�m�	Σ(�#ܭ���"<�;GDp[-��w�t����>��G~n��O�s�ջ���`î+����L	����O^n��w�ߏ=m�|#�FQ�^$�疻Wm]��yGu�}*w)�j�<��Ρ���:�N��U=������~[bJ`RB�$�ʞ�^�      D��s6��Y��v�a��M��SJ�]�JS����YhR���6�3��s�@�ګp�6��X������OR�En���lػjذ���m���s��xБ���vwQ��E��=t�|2�8�ku������;�dG(��u$ݾ	��w������OJ�����58ԷwjŪt�n��WfDyFObD}��م]M>�E�1F����F�O;FUd�j�Q���7��m�F홈��W���Ȇ�+�wP���޾���P��P��t3n��eq	�B��;um�2!�#"9Go'RM�����p@��u���]�����<�" Ig�[��V��h���D��wϚ{����Ua��ih�f�a����k{��=y������W n����2�b񡒼:N��<���b9�����eq	���9�9�X�Vۣ���:	�n�6�iMr�q^w˩B��z�~��Gh�!��;Wm]���]46Wr�*fQ���� �u5j�ȇx���ͮ@ݷ�"9�e�#�6Wg[n��     ��	 2����$t�R%��g\g�˃Ymȅۛ��]0����z�tVQ��M�ءXl�с�[Kmª�,���j�gV��:N�j<�5�s����m��<�#��i�X˫m��C�C�^�2��7�&��`'�=�v#�;�c�Gj�"<�"��<����ѱ1X�D1�74k��_9L+UӴ_�G1U��j�Ȁ<@�Y�,�wQ��W47m�H�u|A46��䯂��` ��Q���G9����o�Q�#Č�=�wP�W���mfd����̰@�I�#�V%��C�Gu��y:�n����1�"�k�v�ّP�#��,� +0}hs����Ƙ����H5�u�dA�}:��TdCA��ϼ��ݪ�>m����i���KI�duQ��Ds���E	�_����� C�wP�t��/����<�������X������oT��pNp��	)V,��qQ�fD�v�=�s��9�xU
r6�H��ll�5��̈�Ĉ�w#L[U���#���*���X�7P��C(�W.:��>�fbG�[�䯂�I��C��fS?f��	E�K����[^�MZ^ޅ�D��@��JpP�8(t�+�4t$��:uN1
�:�D��������!Dዀ�sD��B5z*{n�o>{����m�    䃀                                 -�e붺].Z�d��XSY���J]	��8��r9��eK6�M�*V���`�[f��&�I�+��a���-��aL�K0ku��]�[v��u��Lԭ��m���`�+wB�V�ꚽK�q.%�[]��DM5i`-�]v�n�fc4���F֔ƻh�VRW�j��0Rn�S]�-�����e4Ѳ͋�������f˴M1��T�1�Lu��F�L�ݴūnμKKn�կb����u F��SVm��cef��^!�T-*���E!+�]n�v2܈C���:&�e���U�&���pSmEئ� 7�rY
���_1Ivf]IwxVeJ���ʾ*SJ	�[<|����X(u�Ҕ�Q��N_D���3%J���     vfr� 1l�mu�Du1�u�S\�f������M�ckMI`��CVa,ړVh���%�[Gk�ʗA�!�m6$ۮ�
�,�W:�L�oGhq��@?7P毪]7ly��C�7M���G:���c���WfD9@H���}���-����G;cu� ��~m��I6�۠ݦ��������Z>&!'��z�w�߈�(��v�յ���� ��FE�6�,t���yGu�s����m��<�!��`m�;�w�ȎQ]t)z6��Cm�Q"���>m�z7QΣ�s�����̈�f#�wbڮE�X�	��u[:�]�� ׵�;�|+h��w[V��9�w����O~���԰I*��R����9m'guQ�C1�v�t�|��;�7Q��Ժn��w�h"�Q�}sz�n��9�eQ= |\�'8���iّQ��pf�6�l$���y�&����u�^x���BD9U��j���#"9_9�Vy�mp{��V�(z��䯇m��a��h���������}G���g������o�:  }��   &$vnJ�.�Y��mZ�M���j0��,�����z��Y.��ĸL&�]���v,rU�)6sX4���% �k��^2.V��`��U�����n��w�����I�|#�FQ�C����vdG�?n�">ѽƝ�\;E�	�R!ʯn;WuGu��?�X�wm�R�m�n��N%�0ᘂ�\;���w�[���!����ܗ�Yo�Q�"�xtD0�G���w��ۦ��y�$G1Ŵ�n��w�ȎQ��ԓv�$G�/����O���zUT5����\e]صN�M�ݴ�ȏ(Ȇb>�wv�p�/�H�b�g]���"��"�@�D@�"2�ͮcj����٘�ё纓�vdG�dC1�U.��n��u�C#�9ߥO
�Ӵy�7Q�B�z�Cmёs�(�+�=�$���<�u���?�uwm;2#�2!��2��5�mW�����!����UXg4ZGZ'Y��d`O�<�>;WuG�C�G�G(�}\��k�Ds��9��2W���vwQ��3�go�M��(�H���qz�ۣ��z������kՀ     g�ަ�oR.���F%�]�����F�$�Tm���0!���У6����8q�0�� �ء�����2�v��O�������UP�\��W����\K���(�?~����������o~^uwm;>�<�"��&;v�p�/�� �/y�W��wT}�;�dG(�}\��k�D~#ᱟQ�B}T���mB�-2ذ&��s�jg8vdG�dC1�v��m�A�@�D��h{����Xn���;���'RM����2�b�GWvӳ"<�"��{�+����[���b� ���h�Q}w�Ϛ}��߽|��ȇx���ͮFյ�"9Ի�)��n�����/ѣfBb���O(1Hh�QDQ&�c	AO�.�����	A(�QM(m�R2I7)��P� 5R�b!��$c �V8����a�aϜ <%����-�� �v��Z<:�C��]��r��n���gb<�"��3��M��(�H�b�e��Ҫ��?����,5$���n��m��C�Gw�fQ��ēv�7V�@�1�"�k��iّQ��}&;v�p�/�H��7БQ � I �D;U��wTdCNv��2����.�9б� �%`jݵmpH�z����r����ّx�(v��#9;~�m�G�Z ��dB��v���ޣ"9Gד�&��H���;FM?w�N�d�u�z=:��Ҡ
��    e�%!k�WR��5�R�k�!���!��,��m�u6(�v�)2�:��*;l&v�nɳ�n�U2�q���{����"���rM�����K�����f#�91۶��Q|BDsu[:�]����y�R�mpx�9���W�uջ2#�2!����cmWRmB�H-����%[|2�8��� 	qz���� ��l�G1��7�&��H�ux�FD#��Wvӱ��G�wP�AɎݵ\2��#���sͶ�	&ػt�X�ƃh�P�S��枼���9F�x�����x�M�v���2W�c��������z�ש�����c|>��!"�BD\��6��Q���;�~Yw磌A����D���i&��n��Gh�!��:������^=���j�v���� ���*�C��Q���Q���B`�&	�HH� � :��1F�k�b9��/{��=�����"�d�茺�0�;�	�N̈�f#����6���!"9�^-��6��P��Q�}sz�n��9�e�1�GWvӳ"�Gu	��"�=�ۡM��m��    ��9�Y�j[4��`��
mj�k��Z��A��3���0,��ڒ`�.�*KXL���8���&��~�I�_<UVmS �8Ź(�ǉ���U��_���A�l�wTdC�FDr���Ki��"=�2�b=��]un̈�f#����6���!"9�^r�kmV���"jD09�H�[�"�2#�v�u$ݾ	�CH 1��(�W�{�y�ݴ���;�f#�9-^5\2��#�����j�ȇx����������T�QZ�&�v�,-�aX��j���G�Gk(e�yu5n̈�f#����6���+=����# c�ѝB�lv���ޣ" ~ ����n���� L��dBUO��U\mvˇXq�+����n��fDyFD3����U�+�C�Cuē\��ؚ�TwP��G(�}\���NƱ�;�. �֕t� �V����ݟyQ��_v�v6�uuvاwB��Sdv:���/y�>o�"z�]6��;�dG(��u$ݾ	ί
FD#��V�ӳ��(Ȇb>���j�e�$G14t�Y+�KF�
î�I�*����Ӱ�����vD����p�U��)#	K āY)(���>�Q
����!0!�B0�5A�˷�w|�0J�ٶ��5�5;w{}}�_�o�   �                                  ������f̍���)��q�WF��P�D�65k*&1��m���e��\�8�Y][��4��+�Ү�ٗ��*��Zږ�H�X�F�.���g%i�ٺSmCa��e�մ��]��XYBR�Z�iF]I�^'M��Q:U�X�'2[K���T�NZ �Ԃ�0&�c����m�!P�:夭��n�Sv�E���Fa�y��*�k����խ�.��F�bc�jBئ��ql4�6��d�0�]C�c8NvƩ`o<琍ٰD�%����in�3)�Y[�0-��8�R(���.SKp�i�C\-�L�auī��ff��a�|�:|�
m ?��LD
b��(� B,�C[�Rkv�v�m��l    ,��JX�-�r� �#-40��Ɣmiv0�سiv�����fZ�A�fe�3f�����j4�v�
��Ht��t��y��r�2��U�ӵ��V����x��9F�k�ڶ�$G�FQ�_�@���:N��<��V�"�֓v�v�8���!y���mё�����^�U)�Zk����.��u�M��v�$G:����=Qիt�Ȩn(�E!��B�#jEz*�����mW�|Cu�W�SV���w�ȇ��G9+�yt��u����~������UP���TH�97i4�]��Mջ2#�2!���3m&������P�FE��)�^]6��;�4��ccS> �P��{G���$ݾy�2�b�GV�ӳ" 
��$Gܡ\�m��ä���Kf�h�Q|4��w�z6�:�������+U���Ds�v9N�'�伳��}�%�$�P�	"}�%�$ b,�H?�j���bH$��w޺���&��	�(I�7�K�H'�v$�-����Y����7�~�U��(G QbMq�U*��t�t��߻��H'9v$�H��%�$�P�	"}��*�2�I�$�{�k�A�A$Ov���	�$�H��%�$��_j�%ބ�Iޤ�$�n�G�H��.	 ��ؒ	"~�����ʚM�$�(I�5�K�H'�v$�H��%�$U?{��eA$Oz���	�݉ �'�IpI�$�H�L s��ffe�`     
���*����:�t�Rٝa��f;%��I�
�$K{v�IF��I�#�`���i�x \Ɛ ��e����IӽORM����U]C.��Չ�u���P�S��,�l���N�đ;�K�H'�P�	"w���I���̗��$D��.� �$�H�}IpI����%P�&��~����&��	�$�H��%�$�ĐI���$�gg.f^A$Oz���	�]� �'�IpI�A��$�H���UY��M�$�ĐI���$�z�A%����Y������}���+M�l�&��Bш�6N�Ζ���qpI�$�H��%�$��A$O�o���ʚM�$�R��`�D� �';IpI��$D����MT��˫,В	"{ԗ�Nn�Iȱj'�R\A=E	 �'u����WzM�$ ��$D�).	 ����I���$�NvO�2^^��Iޤ�$��ye	 �'�R\A=�$D���s332��-�1-k���،֪�(��pI�$�H��%�$޻�@j	"{ԗ�Mz�v�]�$D��K�H'9v$�H��%�$�P�	"~���U�y��A=�$D�).���?-Ɔ��BU�@��pP��NA7E	 �&�IpI��W�]U�В"~����	�(I�=�K�H'{v$�H�x�=���4��H'��$D��.	 ��ؒ	"w���Hw{�33m���u%�nGVy"��.��BH$��R\A9��$D��.	 ����I�����WzM�$޻A$N���	�(I�;�K�H$�d��K�В	"{ԗ�M�BH���R\A;۱$D�7߮�2�I�$��YBH$��R\A>��I��C���e��C���i.	 ���ۙw���I�R\A9˱$D��.	 ��N�Ζ��s�ջ��ULݢ��]�� 3�wy珛e:{�����ŉ �'yIpI��A$N����	�~�j�%ބ�Iޤ�$�n�A$Oz���	�݉�P�D�������4��H'�P�	"kt��O��A$N����	���̺��	 �'�IpI��ĐIޤ�$�v�A$Nk���]]�7�Oz�I�;�K�H'��$B$D]*� �̥Ѽ��I��m�     ��l6V�f�Ů�[�f�CJ�]K��G
�Z�,�SBݶ����qi�Ny����!ԭ&�s��J�u��$���t�?�K~����"��U�F]u&�e�y2�/�H$�����M�	 �'�.	 ��ؒ	"k���U�y��A=T��5�9�K�H'�]� �'�IpI�_�\˼В	"{ԗ�Nr�I�=�K�H'j��I�wܪ���&��	�]� �'yIpI�P�!�TOz���	����uW��BH$��ԗ�M�	 �'�IpI�nĐIӿ��l��n�mmk�W,^���ʛA�A�R�Bz	"w���MT�ܬ�+BH$��R\8�����+@n	�݉ �'�R\A>���I���s.����H'�v$�H��%�$�P�	"w���I���̗��$D��.	 ����Iޤ�$�w�bH$��w��K�&��	�(I�7�K�H'�d�l�oO�7BΖΏ�V��*�	��D�*�`s���3�������.	 ��3�Iޤ�$�z�A$O��r��/4��H'�}�$�H��%�$�(I�=�K�H'������ff��Iޤ�$�r�G&Ϙ��c ���+�4M)���>�[	Qi�|M9f�X�45Ld%�H��bA#(%*E
8�P���K��+�q��zۢ�M�j�@� D��CJ�����'�����n��HB A�0�Ȓ2���(��U�P��m�:��tҖ�{@���c$"I	:y00:m@6��R��˸��%�$��`�	"{��^fT�n	'�~���I|��$�~��0I� ʉ�ԗ�NT�ݬ�(В	"}�%�$��`�	"{ԗ�OQBH$�	���ڪ[����v�,�o&Ve�ޓpI���Iݤ�$�}E�H5�>����	;���r]�hI�>����	�(I�=�K�H'���>�D��U_d��n	 ���$D��.	 ��~�A$Oz���	���\̼4$�H��%�$��`�	"{ԗ�?.�(*�G��b��
lw�I;��UVe�pI��قH$���\A>����G�d�����UCm���:Í�\:M7i[�������7v��<����6̋�ڮn&� 7P�;gu	@c���j�wl�Ch	�Qu5m�"�$BIgȐjeV�[�M��m��m�   4� y3�D�H��k��MƘ��&qu�g�cm���p�ityf��қXU�e$rM4�T�����~�:{���m�zUZQ�0��dn��-���!�m�qr�tݰ$C����C�}�&��{޳1Q��Gi[�lȏhȄ����k�ڮ����ّr�r�"bnyf����Nײ2���"�lȌ��V��W|�p��@�i��#���M�"=�"K<ɩ(������2 ��v��ȇ{�?>i���w����=�Sl���	K�t.����m$ݾ�{�f!�D#��n��"�$BIgtwe;n�����$R�	C�uB� �{ܳ��*�u5a��dBP�y_n��7vρ�c��U.km�Ҥ���W$Z�K���+�>iꀑ	%�d�J:���8��ّ+�M�D;�ّ	@m��I�|�fbG	,P T	.4&uGi[�lȏhȄ����wu�۫�WN颓�A]��F#Qk�}���߿O�wY���j�u�dBP�z�J�7v��������ջM���h	�Y�O$��|@s�n����)R�n�N�l     ���2]�K�l��Eslғ;!/ �����+F(e��6��΁*��I�e�S����̩�2��|��y����3����З��VY�0���wM�1��wP��oRM����3�D#��n��"�$BIgtwe;n���n��S�L+	�;fD%�5��j��i]�H0��J�]�i�1Wuwn�_�٘��#�wr��3����8�,6@�"`�B��C
�����}��׷RQվ�9�7v̈8�]�n�!��̈JnoRM����3�D;T)��Z���2M1Z���mn��"�$BIgtwe;n���n���;��VPw�o[��+h&G��4]�f_nծ	�Y��ё�m��2#�2!$��@�����t���*�KZ��MH��6G��O8���2 ��v��ȇ{�2#(���I�|�fb;FD#��n��"=�"4��S�� �VYl#H!�I	!��K�i֍�S�����7v̈	����a$��۬v%�nGV���O^z�Y�;�z��Z���~$ (lG�wWM	��-��;����K<�䥵o�ē^�ޡ�z��.Wn�n��M d�;G� �k�RB�	$�I
�QW�p�-���d�-L��F\G���G{
9P��A?����	,�E�P�V�TD���V��*%@ p�����V�҇���UA���c������|} e�r�xZ��C�G]��h���],mG$���W PA���юo��=��R"���E}Xd��a�m��x�c_G��rtq��R"��؞�A,��rlX���QoB����_���� �q4B���G�[�$AP�@ ��
�DX1BP�E�T"@�P�euq�/���[�����Bl����
��2��֎{�qܮaj�k�MF��ǗY��ma��wfa�zU"-�\WgO9�G���ݖ{��}5�e4U�w���l?֕���k�v�/N�H�^�[r��t�c���:�jѫ݋��0��$[�j�}���j�����1+�&X�p$t���=�( �x� ���!�����AY�D�\ Z�t�v.,�2�:�E���hg2�E��6�ː�W��{t��M�<y�D�sd���<]xw���o~�32�Eޗ�<��R"�m�����ߩ��ܼ�x�8���X;fܙ,1e�����o�գ����j���Dz�C`ےh�Twt�M�W��:�v���600�|0X>B�@��t����#���'i�H�F ��Q��SȂ=�zAa.��H�
 �q� 