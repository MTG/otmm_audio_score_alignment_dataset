BZh91AY&SY��\��߀pp��b� ����a{���T�P�)J� ����II" F%�! �@�A@�����P��
R�P   
P   �B���R��
A
�
 ��R
�P	*��      �  ��  �p�Fm־�C�d^�0 ���ɧ}2�ǻy]���}��#��U ��
,*�� v �)C-���J�n}Z]@S6QB�� �-Je�T���P 
  � � 0 ������\�9y���8 z]�-�=��k���n���/H�� n�b� Թ���I �<����`� =,��O.��;r��ɉ{�:=� ;Ƚ�y�گ�a�3���y�q��� �( �( t{�N�e��;�����ê� �swB�9׶=����ގy��t�������<f�-���x���!d�vS�ǓאnNq�� �x��޵W=��ܼ�y�OR��(�>�  Q@�  0� ������\���L�8��� �Y�yܞ#��0t��{���=����{��T�y5;98Wp �w�cV!��<���3���m��=�\����q�3�����@���� 
 (  �`�F�&������\X���� tx�gT�7{u�nS�w���� }��<]�W;r�B$�w]���w��� rf���^����w]�׻x����@i�ԫ3���y����\��w���J        zS��Sm*�B3S4�24�h	���$�J��ji��    "x�T�S�       ��U*S2J� `   B)��SF�J�  h 22  � J�<�#LM5�42CC�O���o������_���{{}�^� W����
*��UET�h�*��Uq ?�"���e�"*�����P(������*����5�9���0��`����� �\5	�&��w��ŕ�J4L��-B��ҥ�6�@tf!r*J��9T�kBPHl���n;�[��XY�r0���pc(ȉʆA���B1����������*D!��=�D �A�a�(�=x}���f����>!%��g����C�'p��{:9	p�î�ո>^J,i�â_c�bLx�iDe����[���v/����F��T���͜É�gQ�8C��,��:w�[�ԱT$�:+��G	�a&���dL2H�Iu!�;���hu	BS�NA�٩5Z�6e�BPBb���3OD�I	%�hٚ�r�Ǣ����8���{�?��q*�p|ݙ2���_bh_)���s�$�5Ÿ��ߝ�6�S\�V�5��b4V-mL&���m�& y !h�r����m�i#��VM��q�F�h�i�kvH�BTbi������4�Fըݻ`��"s�5_�/'�HI�oħVkAQ�ɏ0�`�G��ʳ
�����[���l
K!)���k5�<���:z��`�iL��Lq�&gR�ƙ�:9�EOda��ĉZ)�#	�XN[C���s �)'�r!�C�4[�}��$�,�_m��;+n��#��(����HC�g�嵠�.�g�э&�fsyo����s�p�j�c�f�֌�7���I<z�c��Č�p��nˑ���M� ٺ�N�]�6}>�ww�4��P�Mf��I��k3[c~xOZ7��A��:��N;�
VBPIi�A�2L��a��$��d���l�4e�������Ni��Loz׈1�nd0!	��;�.j��G.�k��H�6,l��!&�s��#��&�r��FٮUZ9w�3Q�20Ә�$��a�N�JC��:��ϒ��>M	���[~��71-�����VD��B,^�q���Z>^�Ը̒}Ϧy�C����\bK�o�ȦLZC�w�2ȶ�m�F�ѩ��Z��g<���bA�i١#�ӴՑ���>�ڷ��%L�AcS��Z(MC�s{�w2����x�T2E(1C:�#�`-SS^-<������1�lN]�+����\>�	�Lʤ�|��	���!�Z�oVƊ�wK�;��ڟ�x[�yM>9���p���R�TF�0k|�ã�p�B��bbI���Cy�����1	��X�Z�pwM��M5S1��Pe��`�%�eκ�8�\��Br�����i2�D�Đ�TNS�|\��8҉T�dA�� b���쵺�8�P�H�ce�zۺb0 X��
C2�A��I�9�:\�!�i��(L�)13i��#r�) �,T%b�P�&DCC���%$0D�pͮ:M	L��xt�6ġ)Č�$�x�F�Ff��6qM�Ģ;�e|�r��[�CC��&W�&���^y����7�ͭſ%F��W%�&�`��jZ(����5h7��n�<�dU�J���i���&�Gz'��ͭE,S*o��5/W�����&
j����Sz`�P77>E�Z0������a����)/��H;�\Fdo"�a���vbG5c���:ܘ�cH�<��H���g�"!5 �Vjp5.:� ��2p'!�y�ѶFa�N1�ViF�!��<�	~�bl���H3�����<���6�9�������ϡz���kg�L��G�E��1s0j�Z֠�N-n��s�s���Ǥa��!�
�k>Pֹ�#�O|��]y��S���0�Bu�q���Իr0������hdbi֮1t�]��br��O�M"͸r�Z-�w�:8�pl��4C���͐hrM1޴�'#�Z��9_�d�&�iA���{v- \� q!��׸�"Dƞ��``Yvj��,�*� �!4!F��Γ��|&�k!:�c��ţ��.|��%�|5G�oX%�05�<z͞��g4�8�:v��o1�;����+���SVK�w�߯��'�ƥz����]�nj�*��W�5�h1	���U��w����R���7z�je[a�S{Ψ��yɘ�|�{��7�>n��G�λ�}���N�����9~�������}�O�/����7�.�kP'���4����!E]6|�����وiK�V�m_|�.��HH�q��"MjL��MA�5�$��##<���M1���8a���Q]zᝩs0T�g>��$���7)~�����w�}���F'�c�[`�c�5�a�j��A��b߽e�L������;��7kx��[�[@����0y;\�\��oog�<�t�gmX1���7�dl5Д%	�έ^�.���&�(��2(bj+�g���.��'}�n*�Ğ14���dQ�ך��a�XIk ��v�o�6泘AWݜ�8h�%�8e!�`i߻Ύ�pt�k|�gA	#���x�;��A8����;='� ��oȎ}���8�oj�ܻ�V��Џ���qpMGd����Y��/7�pN�i-_s��}�\#��"���Ϲ���>9u�����r���_�q($�9	\_s��߽�5`�vj|�U#=۪�~���߾�x���q����w�r>T��N�>��h���I�ߧ7V����{�U���~PX�b��LK��'́k]�����o�����N�m^ӷ��~X<�Z�#HMsfK�f�v8�I�NGp�rb1璃ɆA<�o����?.Y��8>V����gw��ۍo�-�ȁ౴�24C�.
��$� ���_q��G.����.>���]¶b-�2��Ss��nq*%3��$�!)4������Rv�b!�k8F�@d&BT�%ۖ$mI��'�ø��$�:���|�<r�m�g36l��a�{�����	��-�S�N��ڵeD��8�gA��2���(�8NkF�͔'���f	�&��z�<7�<�GS޳��q�I����i��a2��M5���-o�=8�t�����vBS����I��','V�"l���֜�j�&)U[7��{��q	�1�଩#�!&��s�"�qj��qA}��E�[���$��I4ň �5 �$&�T$??'}�s������mk>5�;�}9���(҉��g0M>��#�D�}���I9�ӏ��o��|}9F
E����z5�K�n��81�q�]��O�� �vG��SIw;cF�<����MBy,jq#��=Br]>b`sv&��ڴ�0���.FK�Ya�̓v�G;t�d���_���	�,O؏%25���KⴵD��X�M�\��8�W���o�y�i�F`f�0�N���gˊ	�sc�_s[�6�	6�©���_';�H(�k���>K��}&�(�ȸ��h|�>�y�3n�� �D�1��%L�.4�1���osu&���[�P1Mg$$�L�2��v���<'x`�$�W����4�]T��Z�,�.�4j|K�<�%��&$��l�0Mɦ2�|���%�$���=��p�}���͹��{Qĸ9��k����1eĹ�yw���f��Q���M۠����~���>�o'q�n &�Ux��H�=x����c�sY��D��~Θ���M_!��|�ቘ��{�*�~U���E񑊘n�'N,����?��j���$�g�!�&���C0M��٫Q�ዽ`�u.;�7��qr��}�.�����_�&bq)9�S$Jj�D�U(��EK=�	pY	�x��]ɉ��1������f�z5���v�Y��C��q0�RDL�L��t��Hy8]跆19��:��b���&�c�ۊ.r��g��������+�t��w��s�F�15����E5Q=�"UZw���(�-a}��l�^p�9�W��}�e�ϵ��š~�O�\T.��"�
6�ʡ�����&w=4D�Z��SӅ:��ȧ�y����5�	��'9��9$�>��9����������l�fآ{NI;r*3�3!-Ie�����Ĝ3�1*bd�9��E��v����8f��FXX66XS=�4���9<�ٱ���%�I�	X6��:6q�b�[8pug[�ؘ�h������ظl���}�j��}��eO'��\�oQ���:'&�|�d'>�+k��/ͮ�"5w��:+�^�,^=_��?��ԇd����f�P��>��������v��kq��z��_y����_��.�-i��|�ڹ��'0J��i߷urs���-Ҧ�I���nc�_*5Y�w�T�G�-r���h�[3w[�rk��q
����[�'pJ.D�hM)��`�^t,OS�+I��8�S��=;:�auV$���b��cL��`�de�fڴ�� �h�4��&ХCH���QȪ�Ў|��\�ٲU��c�AG��'��Iϛ�r$q�F޽��.�Lx4*�_��K�%�	e�ל^����Վ���7���X�π���
q�BT�*w#�S�¡5�bkS��Ɋ��"i�5�VR*�
H��.N|J'䍛����KS�r$�c�'k�K�/>=��5C�&��-�5&�D����>w6��{ڟ�dz��N��������#�&���gl;=�[<���1�E�=B��;��;u���6rc��s:`ΰq;����I�Q��6r6u<Ѳ1���e���4d�$Pd�e[�������׊*�iV����]�����w�]��&��ˈ�*\�'�J��EQφb��0�:�)ǩ�~��w���)�}�V�U�+�Zph���Q�3#r��5&`d�c�`a�n��L��'L���8o�"�����odן!G��&�08�|�`1?�ƣ��n1X�&��L�s��S[�����nE�.�E~�$�:C�_%��5?�W��;�^H��6��W�]��'޽��s�-1}��Ѣ�2�v�1�a�0� ���1 ��NBP�&�Ð2��jMC��Η�p9	�8���%�5&��3��{�氀��u	��,d�`O]`����Q��w&�'!��M�0E�HC&	�	�J�#E�'����0���=�k\���Ha��B%A�FA���ְt����~��?3��#��ߕ���~X΀m l     (     6��p\�2�j�    �` 2         ����Tsan���+H�7A ;.Z�\�aeqhN�v��bBv���n����Xy�ˑ�z0��:���^�A� 2�1.�'cO���*���PյC�cFy��Shr�N� q,��$�t�Vy�8*
K��_m�n�sjUڶ�0��`�H8�H+k!��kEY]��S*�UmY�R�����eq�S�����ԠUWH�%Z�V�x��\c�����]�zX(p��ﳻ��ڸq<����o�yC��7VnҨ�vVԒ��3�V��s��s�nq*(n�QU���3χ�x�)�]v"���8�$�wbI  p�`9J86ݶnMzF�Z�6���
;�h�7D�ڬ��$%������Ie �nwD:�4���TjN-�;H[��mmn��rp�$m퍮��+��fԫu�"�֎�T��ū	u�f��4��O��!ZL�nz�!WF�V��,�Gb)yݲ�ی�yG�n���R���켛3ٱz�:7��/���ͻ-��Ms;�]�`�sKscL�p��l�\�W�dzgN���v9�i2�G�D=n�en�x ��T���q���D��I)�knb@j�[/C8�i��6�E��I�c�v����$��Xvl[D�6��nr�jBBE���t���U[r�WJ��̨��6��9V���	�m6��&�&�؎��/V�hm� �6؛[3#v�!oU��Ah m��G�o�m� l�	��Z�\t�6�9�&�	4��� Bkv����|��S��$
79�xq`��t��ZD�qڗ��Kb5�wc�`]�g�t�J<��mtu�f�vv��b�.��6�c
��Z�q�Om��f^k���1�mk�uݳ�OMn.�5:ܴ/��2��uOO��i�2Mr��*躔v�XkY�i:Ζh���B� Wn���^��Wj�!v�r�İ�Fښ� ���6�H6�yn�k�¯#��j��3sf8*��"�, ޕ^�8h�*m�Ʊ�0[��2��ݧVeY�SW��*������K̪�f��0 �l�-�k�5�Ǫ�W�*p��MU� �Ml����]9���)j���A��Bz��6��H�$l↵��pJ\-��l�� �m�p�jٴ�kdk��Hk�Kk�	:ƒ�k��8v�9ԩi!mp[yn��[��� ��z�h�ն��I�h �ζ�K�l2R�  � oQ�aQ l�@ �I���>�"�۶�	���$1-���8/]W�gd�$��Z�}  H[ƶ�e��u�-���k�o[M� [@s����h �mӦ�  -�l8H,b�� Y@  pt�Ygm���m� �cm��6$^�9z�'�/�l�}u�m��  -�-��z���>xJ�X .� �O���k�t6�Zʠ Kh� N��2ӛa����I$� �@6�m  !��m�6�@��D*Čt�6��� �I�[Rdpmth�:�]�Ma!����l �0�5�ז�Pl 8[v�f��[r@  � �mj�p����m  q#m�l�R��z�8��:�  ��l�n.���vP�V��cu=mu�UU� 2$[@�i�� � ZU�UF8��媕@���  m�Hm�    @ ��H^��)@Gm����  �      Ͷ  9+j��m�����WW`6݀p� �L�Arh�ve�`6�"ޠ $ y���lگQ�gL{kx�������  	l ��R��@ ��\�-�@>����K6$ �4�T���m� ;I�q rn�:���6hm��i������o��t[�6�^%�a �m�Ͷ$    m�[@�	 ��� 8�n��t0�X�I6� ����[���%��� ��3�`H� H�6�˦��Q��.[����)6-��  �@�p� ��hH��j�[�4�j�I�����$  ��  ���Bؗn8צ�b�u] UzڥBf�K9�n�k�llh�I ^����ے  ��wim�ˡve᪇+�X ��:rt�6��6�8[�[)��� ���V�x�i�lEUU�+;lvۛ\�m��r��J�[Pu@�37,����؏Uۉ�.4�ՎL�2�Ƅ�n��q�pM<��*��q�l�R�I;UK�v{n���V}��yw\uU�F�k0�]�m:�8C�P]���5St��qTd9m  Ie����!��l�{:l�j�v�yPj��W�� ��T�;IΓ�ڧR�֤��6�1��6�� �D�jk���N����`  I-׵­���`��m& H-�f�  �[\ �m�h ��h��oU��Ie����6̴� $�   m� m� �A�iͳH��UX�(�����&v$p�-����;m�i���I�t�z\  ��<�vF_/Cn��p@8���^zJٜMQ����7[%>+qU�6Y� ���u�kqc�9�4��Z�I�@۴�ݝrP&�T�Wl�����I�嵴�	;�GF��5��Go��{�e�|��1�V]�L���8r��j��'��z�((gE!t��Ͷ h�mj��Z 8i`UR�9v;&�WR�V�pm�X=p�VҭUW\:ϸ	����=v��[+M�f��5��"F��U�������dvv��e�v��Z��@��+m�X}��7��!竅��-��ڧP	ڤ�v�unf5�*nӓs���%��쒙k�2�a�G@]�i�**-^�+`��ֈ��UjB����ɱm+o)��&H��[Q��8pC�ÛE  �ས  m�V��9m [V�m�;�q�����~���  �#n�.�amm�n����  �6��:��m�  ��Svٶ���5U[~*���Bh�	P�2�Վ���T�eȪ	�U�T6:��k4�K:F��eb��5A��I�ќF	��^ۓso ��Y��˛H���l� Ig��Y�]V�K�$:� m����d�HORD�v��h�lsm��@��Nc&˫l�jڶ�e���� l��@[^��sn�[g@�հ�c���qa�"j��4�s�U[*�J�U⓳�\�R��J�5��WE�p� ��㯪��:1� ��Av�ⱉz&�uͳ����$�u��j���GF�FSka�2@l�x7YB8M��9�W��bWcnZ���1�\��]p���\W��.�J�u1�Ɲ���@�k(�+� n
ٶ�R��*�Z.�P*�U7NF.�2�-���t]�u�6�%�(�A�P Im�>ͶGXf�S .��i��VζZ�&؝��K��W�+WF���� m��
�gN�I m�\�m�  �cl��'m%mfrշ کM�ŴK[W.�J�M��Qm�Y^k��ۙ�m�[�oh��I��m�,�o��M��j��m�m@���&�n�$]�ȼ��T����k����gB�UR�<D�Gg3[J��)q���MUVW�d���N��U�7�ҩkUȵWVzӇ6_P�e�m�&�9ʥy瓴��iZڄ]��S�.qH�p��`��8	�!X�Lu�Z��q�V&]�	U(R�ܜ�:[�ܜ�J��������� �tޛm��`6� �]$�@m�	(Y�T�z� ������JK�T�P]\�hX���ڝ  ��m��Z�L�h�m�݀m��bmu�Am H �].ց��ul'l  �m�����H�i�P 6��T�J�UΊ���P'E9�` ��tعg�j�"�MTUQM��m�N�M�� a�db���֦� *�U�f�i�AJ�G�Z*�9c�s�J�� �Kmƍ��r@N*�U*�UTk������+�']����g�G�(�2����s�Wa�]	-9|V�!f�$���g-��n�ޝ9�^��ͳJ���/"��UmO$�uT�UԨ�˟��Z^S���UR�W �h(-�6��m[  `�\����LruWqd�jKd��d@$h  �6ۀ6ش��vۭR�\��� 9@ V�ͶJR�^����p�-��� �m/K���V��YL�A�V�PQ���f{X��-�'A%�v�  	ΒP�2�m���6���oS!��@�I-��lH	$4[%m[? ��V�u�[�$��e� 	 @H�� "�׭m�k5�l �[��ۈ�p��J��UV�m�h	W���PԚi�:mp  �����l��]Da-����6�U* @�]$�[pm͓��2��egd�bڛ��uM�"Bk�kƂ��@!7O��ff��6KO����~_�e<�k8�)�E;��NV�{bP6��R���C��m9��t�g��T�Uz���N�4-��s+&�HH��4�dv�$v��r����w�����������W���?�?������W�������H�����ҿ� HQ��N����Ҡ�* LA�%! BOϰh�PB���X�!�&P��[R���`��n'H��N�� iM(�
�OCf�������x=��a1(D!ب���;8s`IӋ�G����,J�JI�c!(ANzM�K$� � J��OD;@'�)��
B	�t@=y�<G�-(x>�!�1��HJh�P�; �P%De�D;hP�e�<A6�w��+`QPQTA,��a�/��
������M�P�N�^��F �eY���O8�<=��}HS@1B���E2< |!<A �M��P\�N �M:�z�Qtv��  �H���1�8����lb����
U�$�8�C+઻��v������}����D�|�
�,��* T�$��vleE�$*ZHCJt ���(�#��Q!w.pC�@�O4��b��JJ'���&�h�B�SA+24PQ$�@ ������>/���o�ڧn��G==@چՕ�6�hC�q`�$&��;C!RBY4i]����"T�zD!����-I M���E�$��z�x
�C�A��Ⲱ11�,l��331�32�|4�`IQ����ꇲK+`!��1D� �:Dti�V�BDw �B�HD0	�"��4 �1u�i!��i-�`!�XH܇4��I�(pQ�	M���i�S�����C��U_�?�_������?�~����3��f X�"b�
�9�(�5-���P�̆h,m�P"�48�9$D�8�;o�t����m��\V�D�m����g���'_T��ru�nn����$��PX֮�,�V�"�-uj��r�6���c����l�n�k���V��ѵ�����<Ldp۶����{+��.o]�-�\�������ݛ�|�8��é�r���6iy q����X�����A�=�֛y�]�:�;=���vތ�Xi����{t���綷�ݶ�NG���V4��s;*�E��G&փ�]�p�-��:@elKۋpnऀ��K�P�W�%|�6Hw$ag��4��[���	8[sk�[
����m�M��f٫���J��4[���]��K�m��&,&v���k�Ä6:���`�	YT�%q�E�P�ݪR�b5����Wg`+`�\G+������ʽ-�^`# �]6'�ꬬ�����l�em���M&�4��D�P�[;ں�W��"����n{\UI�Y�{v̰���O<�7H�pM�q�n�V�.�v����Sn��8�n��݇��G)x�.4��na������d(2�;M۰�%Bk)�͜��H,I�r�i9��N1��\��4v��#�3�ۇM�:��=:���r:�,��v���v�k�ͪ�e4�M�*�;pv�س���K����F1$n(�8��i9o	�)��=m
d��\(�[d�tS�V]�b��f���s���ќn�b���gnOg��p&���i�mӣt��gs�:CX��os8�ҒNs�Lc���nRD+i���nw�9ԁJ�*D�8$�'���
��b�Y���
��ケ��۱*=�Bqt��[W���Sy�O3ڱ����y���9v"�uԡ�"Ʀtq\S��99p�*�;��f��Ih�<�R۶��=��e������&6��V����s��pQkqRg��Ԣi��dt�:�;Z�iV���i��ʨ�0X���ƀ�-��T:Q��ʷe9c*�6 KTa��qpc��x��ے�`WU\Ոs���~����=��N�~>P�B�|U�@ S�����D���b��*�Gb�=%} N�د]#� �Q�Є���	�eC�X�a�,ts;Xr����m��E<.7M	��N�zs��,��&��.4)���q�y�k�L�8���g���k����]��k��g9d2�:N�q�,������q����c=��ۈ�-�.�U���w�W���u�S�M��e��c\^i���m�����ݵiM��q�u��nqmK�:R��eCjT���7kz���/G�)�\C�ﳻ;�ݸ�'c�p����2H��d�)�H�@P�6�b����h��P5��� ����9��(����l���f���ڴ?���t?��s�诙iS��r����w޺�I��}�p	�Ào���T�hi���4� =�z�w�@�}|hy�;���挓8�Eu�t?��{��4?���tس1f/{�lk�(�7	���oGc[� ��"m׳.��Z��q��%pR!yT����ή�ۻM`c� ��p������}4���h�q��E!f�U�w��g�t)%I�j0t�Ć��]��~������B�O������_}�������@��ߦ��g��T����r۠d}�Q�V�Ѻ��;�F�U`|��s���l���f����Z���;��=���h�$�w���X*�Gi݁&�<m��tCmvꂶu�z������9`��슼����&Ȝ��S�|���@�g��?��}�{V���J���,�P��Y�w��z���>���@�����f,l�?~h�0��T+Ik�>}��ʻ��xr�ē��1\���Ea�3�=�*��{�pt�#=X��SU�ܳ@�������h������}4�﫴P���V���}4�{�@�������h~���qpu�:Emݙm��������=��'6ۮ�㴁��m�	�j�s�\ �����q������h}女�g��T���u���>��$�l��ߵh?{��;��=��Ҡ��J��h{�ՠq���~Y������@��ߦ�ϳ��N���S�*�Z{�{��z{����ԳK1�/{}�@���DQyY(RGl�=��=����=�{V����h^]�q���h�cs�����\��Ÿw�t�	x�'�[�zF�1ćd�B�[,�@��p��W ��J����\�p��?V&�T�ՎY�{�������<��M�����}��֊�UB@�ՠ|�女��zi�$���ߞ��߿j�o����HT�� �\	_U\�%����{�������<���ڥ�����נq������@9���}���R�!b�!E���~r��kEj�jU��]`��ۇr�/\�]U��i
�>�G ���v�P�/;C�h.�ݍ���c�r��`�n�ݺ0v��UP�qū���C�gBk]�w:iwm̙ܽ�\A�q��4�ʷK�C��v�'ev�X���: p�We�T���M���y�q��O��9�����u�gpq�l;��g5��$ө�A���y��M���$�s��71T����[`�֘ѝ�������9A����{6涁ɽ<��,���+��4���bt�k $�����@��4vw�@�s��N����e����@���4vw�@=�z�[=��TH�N�%
8����q��M ��������&�;
m4���_W��틀H����ޞ��9��$=��q�Y%��{�@9�}tz{�@�ݾ4�K;��~�b�M�P�NNF��5�/"S�4ڼ�d�V�r�9;q��0������z��m�}��ջ|;�����,	?~���MƟ��W۠{��{�z@�}�f��+J�E�f��]��M�@9^����W�}��U�~z��?3;�?!R��M�Kk�>}���t�w�@�g��z?
/J��m�'M6��껛#�}��������}4w:+��
�`�v� ����=��=���h��]��+?~W�c�ێ�y85vS,�<tn[�Y�:ܖ-�v����Q1����be�@�h������}4����s����E�
L)X+m��}呂{���w���=�cg�O?X0�q�X����@9���1LB�Ϧ��I,m�Oq�}呂}��x�&8�1�j�3�ڰ7�ZX�̀o�j�=�v���V�"�tw�Ɓ������] �{�w��zDӵʄb�RTz�+]v*à凥��n�wOg���eˣe�Z�7;��e%�i��-4}��@=�z�>���ק �W�*��.�i�զ� o�j�;���V�H�3�V�y�+��	T�I#�@9�}tv{�@�g|������E��u�F�tz{�@�g|������f�@|h���߼�*��G�jӗ�v�i� ���p	UW�#����;��=� ��72dl��]��T	�v�ǓE��on��������R�k��͎)��.Y�If�s���w��{;�q��������8�0r� �{�w��z{���t�w�d"��6�����2��\ ��| �{^��������[i�ܶ�����{޺���@�g|�|�Z�Ҁ5jLN�mp;�����ǀ{�e��<�\��<%QH��¦2&��%�.��5���Zd�8���rGIVCv��lE�F�֭Mt��ݗZk^�N-����}�t��XE��h��Z�-��geL,6^qm0g�/l+pfT��Bnd�q�VE-�Z���Y���é2v�Xw�	����������T��f��D �#�|O'%N��C�Ɇx8���	x�'��G5�QHWl]9���s�r��L4�N�����gؗ،��f%n�n���H��yv�s�*.�i����%��/a[ۘ�ݻ;�Z7&�O �N��ƣ�9%��w��>�w�@��}4�{�@��*��ʺ����d�@���=����8����s���;��@Bc<�`��W�q������w���N��O��=`��r̲K4?���}t����a��g�{����c����s��s��p�}3~�����zF����Uy�����(��/��]=��m���Skx��ຒ�����]�:��UO��m�z=���ۼ����n��}R���[i�۫���ߟ��W�/��x�T&��+���� �ʤ$� H��!�������v�מ{����	�P��YT��߾��9���9��W:����]�vK"�I$�s��s��s��y�}�j��k���U]�u�m�9��ڼ���������ϻ�|�Q���
��g��[wA��\Z5���U�66�i���D���1]@Bc*�<��up����}�ns���9��W��X0�r̲K3~�������s����>��Ջ���?W	�*�qM[��T��{m��o�X��ω�������Xk���X%��Y��i֝9��׳J���F���*�1*�}���1-呂�1�؜���k �3����p��Q�09����{��Fj@�z���% �@]���	ʇ3��������×~��R_N81�
����m���l��cM,q!�$ƄHkSgby~ŝ{�XU�Did��`9�9����(��3������ ���.�Q�t�9������ ��t�X�Cz�1��fּ�Z���Čq���[�1�wK|{�1�a�`]����� >�{|�V��qz�fb����e_P�Xh�͏���D3��
5XRP�@��l�y��$��l@��;M'H��	���z�t�> ���T&a�T9����A�!�!ث�� �*C��PSb2 ��G%:Ϻ�\R����=��ԥ)y��������-�{━I�ߞ���R��<��qJR�����R��<���┥�Oߵ��o3{��3u����)Jw�{���)Jw��pz��.����JR���=�cԥ)w������8�\	*c�n�Igjn���M�ݝ�t���v��{o�����?<k���ٽ�z┥']����)K�=�|R�����~�~	@�R��=����(������RRQ�$����3�}�|QiJN����R��y�k�R��w��pz�JS�#Gٚ>-���y����{��);��߶=JR����)J']����)K�=�|R�����ơ1��E��v�ᘁ,ľ}��R��{��pz��.����JA�	_ث�N ��`PPIq4����q�����ǩJS��~��z���ޝ�o|R����~��ԥ!�0_>���|?{��K3��b�w����
ڦQ���j�m%cmq�cq��'��tx7���G����H��lc�Dq�V�3����JR���}�cԥ)߾��!JRu�}��R����Z�_a������)JN�|��P R����┥'^����)K�}�|S�*�ޥ��!J�h���ݫ8f X�H����qJR������� R�~����)�=�~�8f �_�
?ªE\�ڣ��� �u�}��R���߷�)JN����R��߾��)JRu���}bj�5�I.�ᘃ1{߮� �D~	��~���R���s�R��w��pz��<������f���ۙ��gvk���q]k��vs�>K;�WOl�����N7 ��5��7c;�[���n(�=�U
��3p�7��2ttc=W�.�
� �-����q6�.l������g��{V����M�� r��Ges۞�X�rnݴ�<uV��!=�m)]h�g1�j���v���#�`�O.���l�x��1���73�{9i��ٽ�l�b鈢=���w�����y������u����U���t�C8�gY���L�ͅ��:n�{׾�r]�tv������JR}}����)N��~��):�Ͼ�R��߾��)JRz������o|޹͏R��y�k�4�'^y���)K�}�|R�����~��"R���}��Յ�n��Z���)JN���=JR�~����?�	�y{�߶=JR�g�~��)=��>5���4l��7���z����~���Òy{����)O3�k�P)I�~���JR��]kU|��Sk{��);���=JP�G�}��qJR��>���ԥ)w�o�R���Y��٨�r88��	]��թ��N���*���-���sOf��bf���m�
V�c7wb���y�k�R��{��pz��.����@�);�=��R���j�5�F�ռֲ���[��):�߾���I@�` � q�p8R�=��┥'~����R��=��qOȀ�c3b����_�'d$C�K�8bR��}�|R�����ߴ=HrG%;�}�\R����>��ԥ)���4}IhZ9l�sbI ��_��,ᘉN��~��):�߾��)H�ߞ��)JR|�������oy�s��)N��~��)C�=��R��ߞ��)JRw�{���)O�'�}�s���|p�I�g��l[AP�m���]���Z�5s��#ء�!�{�|o�p�קҳ�'~����JR��~��);�=��=JR����)JR~�ψ�~ޫѺգvo}r���~�
R��3�~��)Jw�{���)Iמ�������Z�_a������)JN��}�Cԥ)�y�����>�p	�"��)��1J$>T�P��:)=�]���R����빈3,�R��~V�M����س�JQ�<��qJR��=��R��ߞ��)@�'~g����R���_F��ن�kFof���R��y��pz��F��~��);�=��R��y�k�b_�f.�G���x�[ad���%ۇ\�lm�
ۛ�zɮ#��mvLb.�v%�ǻ�>����"�r]Y�1��빈�����ߴ=JR���� %)I׶NW�}��VׅP�TK-&��N�|R�����ߴ=G�Y2S����┥'}���R��~� )J��>�Lg�QEk�݋8%���}��qJR��}��!�*J]���╘��~�賆,��;���Uq�
��Z޸�'^����)K�=�|R�����ߴ=JPi�<�B �H���(`������W�D�:��┥'^zG���c�vjѼ��ԥ)w�o�R��߹�hz��;�=�\R����~��љ����ē��dM��1�&�cjYMle�6Nݱtn�qL`T´UF2ˑ��qbI�rH�Z�m���1w����'�S��ߵ�)JN���ԥ*}�~���1��#���o�M�������R��=��pȢH&JRw�߿pz��o>����)I߹��hz�	b��_�
?©�I�[,�����}��R��߾��)O�  S$�����R����ߵ�iJO{|�~���9!$���bI#�{��X����~�cԥ)�{��┏����w[>��In"$8"f�*�jg{�	I��}��R��+
�����)JR��߿pz��.����JR��IbPX�gߏ~�ꖊ*����������K�ݢ �Ԇ����۠�S��z�:,�&sv�q��$�ȋ.���ݻF���n蒌l�5ӌí��.sʇ�5�[��ݼr�:�6�9�A3�4�k��1���F�`�[��9��=b�0Y'0<&��ہ���з���2f[vZ�r6�5���vƷ��� u�n"�e�ݹ�U�,�Ȗ%�KوY�[u�ȝ� o:q��;���Vv��u��-�3�m�lnPy݆�3����UV��ڳ�b�����┥^����)K�}�|03b�����ᘃ1|������":�o�Z޸�)I׾���EiK�}�|R�����~��)Jw����!JRu����4V�Z7���z��.����JR���}�cԂJw�{���)I׾���JR��]kU|�6����J_�vI�(�������R��=����I׾���J D[�����	`,�R;���P�s��ԥ)�y��┥" ={��pz��.����JR��s�~��R�}����'SϷPʺ��Ykm���A֬�m{6��XL�iCNKWY��X���5�a)!�ٽ�z┥'^����
R��~��);�=���ԥ
w�{���*^�t�~+��䄒���3�}�|����j$= v��34-�bY��y�&
�����)I������)J}���\R����~��Ջ$�ˤ_��~%�k��w1��������JS��ߵ�)):�߾��JR�~����)I�ߞ�Z����oy�s��i;�}�\R����~��ԥ#w�o�P4������ᘃ1}�7���":�+Զ۳s)Iמ���J�.y�߷�)P�������)N��~��):��M�o�cs�1���=����yg��e�j.U�v��m��.A	䣖5[�fb(��5$�hݛ��J��{���JR��s�hz��;�=�\ �):�߾��)J^}�j���f����)JRw�{����2�d���ߵ�)JN����R��߾�� 4�~ϟk,�g�,��Q�9�hz��;�^��R����~��ԇ��~��r
 �m�@�eY���1��Z�;D:a�	�������)I�����R��yya���n֌7�{���(A);��~��)J]���┥'^g�}��R�;�}�\R��^��</Ю�G$�۫8f �G����JR�z�<��R��y�k�R����ڳ�b���"�#�)��ݷvz�L�@hW�E��X5�L�n�׶�����T���KB�,��b�����hz��;�}�\R���}���)N#�{����1~���	���(�{��R��y�k�~H\���Ͼ���R�����┥'^g�}��T�;�C���Q�]�Y��3b��{���R���߷�)� '~翿hz��<�_~�)JRu���mѢޣFoZ��Jn����JR��3Ͼ��)Jw��8�	0�DC� �$�,�����	.��!��(R~��<��)J]��ֵ_��K{���)I�y��hz��?#(y���qJR�Ͻ���JR��]�A��~����c%"���Kv���ņ�+��F��==�յ��0���	T�{�-��*m�`n�Ŝ3f/�=��b);��~��)J]����JRu�{��Y�1b�����"j�,�s)I߾���?f)y�߷�)JN�Ͽ~��)Jw��8�R������@j9%��Y�1b>��]�A��:�=��R)Jw��8�)I߾���b��g�@�KH�,��b��BUrN�Ͽ~��)J}���qJR��}��R���L����┥'�}R1$���Uwrσ��-�E�R�~D<��p{��/?~��)JRu�{���)O�x{��>��\h���2���2x�Ϝ���u�f���F��7.>w�@��)�٠́�M7�4�Hy�|9�p�N����k���t&����FA,�l��;��?m3��`�<m�O�r5j�P���ֽ(�I��4f�j6�g=��/�`7�Y8�F�:gNb���T�:ڢZ�O @�;Ѹ��h;�	�:���c'��Y^�;6���z`M)��l�=5�Y�I;�m�m�ڃ �JU���7�Fݏm�\�GdN:ut�We����H�D1��-N�����}�6�\��ܖw�ۙ�����[�d&8��u���.�ݣ^'Wc�: :{P��w�:.l^�vn%۔�v�9��.�<; T���N����'o�۷���<1�q��8�nQp��!���V�Wa�r��ymK<ag�!M�kGc��mTu*�Ge�状���N���gS�n�s�K�9�s)!�����u��ջS��&�k��r�Y�!q��b�]��V�|�kn����;.tc6p4�:DX�mr*m%�j��K���:�^�u��M��3��*뗷$�5�����e槂v]>Ļg��t�N�
��I�D���=��J��vШ�5Z*Cp�M�H V�K���K�� �ۦ�K��X�`)����T��Z~���#��/:-���'[���/l<��T��\��L9��.�՜MVn�K����-��&b�vw��3�v�����N��\�sN}V6N�A���L�k��Vu�v���C���J�s��Ԭ�!��&������nwi8������4�.���^�ǵ\\񹙼���Fqشg��.�nz���۲;x�p�F�{L��e�;&�h��u�6��y�ՒƳ;���0����Z8w:X�;b�n����7D�Ƚ�$��\���K{v����pni�v݌�����.�X�<�k�#v�_Y��s��E�a3D�U�$�;Y5jsF'�J����:�oԄ��n�U'QJ�^���u��q�`C��:3�]=���n��c��|���k�mw9��÷3���a3 ���$���@梭qT�tp�Ы/*WC[v�(
b�ζ��r]�U����Ë���n���8g:9w��ōBu:%m��k�=��R
�Ҥ9Gm��R�2��;sR���j\d����R�(�n����Bm /V��h\Z�{Ψ�a� 2�gc7<�� ���kv��lپ� L? z�z��~:T�/�~�,��������ڝ`�D=1OP;S��}A Ё��At�#��ۿ��	t��3��:ې���<����'�+����/h�،E�M�*���N�D�8^�Fh�e�tv�6��F�x�>�7���ìq�j}���p9�M��nx�v�*slH���n�\���	��ݞ��z�q�0+4�#q�"]h�)ŵ�z��3�����[\�^Ӻś���v��d�m�;�zs�Yk���G� օ{��A�2�sCKY}绿o���������q@Py>�;h��W&TQ��;Vu0m�6�����X�.�6H�����Ń�}r�3f�y���)JN�����JR�Ͼ��):�=�� JR�{����)I׾f_ŷF�z�f���R�����?�a\�������R�����┥'~{���B����Z��f�ͦf��)JRu�{���)O�׿g��H�I�}��ԥ)~����JR�������g�,�zk��4=JP	����┥'~{���)K�>�|R�
N��~�Cԥ)�^E�gֲ�o5�����┥'~{���(D����)JN��~�Cԥ)����┥b�z~��)p b�e��i;�ǝa���6�� (\��!��s1"A*j��J�M6�_a��}D�}A��g�Ȱ��9����=�v`F��$8"f�-r[n���~�9s�F����S1bA����$(G̛��I���������ݞ�����]� ��[3�_М�^��Uws�-�Q`w�٘UU=���� �E�Du#�*ej�+�Y�����8���t|�"�*���p����W(*T:B�v�`���
���ߤX��|������k��I���@� �s�c6�Mƅ׶�ao)��ۋ���E�w{�_^W|Qt��Wi����x��|��3��� v�� ��e�-1LDT�]�]`Ӫ-�ـ��K0{UXG��`�_U�J,�$NЩ�M;��ɘU����^�`�j�A�s^��wV���Ui)Sb.�������;�<v�����zuE��wf�ޓ�|R�Z�!v�@ݤ�|��ٰ�ٷ��Ł��,����5�u���o�hݣ����6؞�B��k��(�n]Ј �N����K0ik�B%��
�WwX�uE��ږ`���fp��W��v��u4LL�45��ك;0ڪ�>��^ �:���^���($S�*�i� Ol| �}'0������L�M�$K,�J�]Qi�;����׀-UŁ��K09���3��)�H-$ M@�� ����`� �Jg_��|�����Do��:�������@�I<3������uX�y+��k����AK�� ��m<�\��h���6۷uv;Y��������c��B��+}���K0媬５�`����X�l��ZI�o0�c�����[/�w��0��M)��TVU��"�M�����7�e�>;�I��#�	3z�K2j&!�"���m���yL�͏��{�9�o�wX���$35�y,�9����u`��ׅ}��9V�xX��R� �X!8T�aB{����5�f�oj��Ț�]�`�5�g"�=��GW�zZ��-�K3�Gw���l�u��m\v��T����N���HuU@efq�'NV5m6p�gZ|98n����\v��;�wb�M�dMZ����Xx7Q�jmh����hѽ����㩐��3v1׮���-�u���� ����O5�.��䳞:��	�޸��L�Ŭ�j4&�GA�n�7��_R�%��ĵ���1�0Gu���ݍr���q��&����^����M�U�\�j5"��:�߀?���`o�^ �:�ـ��Y�Z�2&������]�����`V����0y*� ��^&!SA��WWx����f�/%V��W�(<1f�ݓ�iX�&��*�7�&`���USV��%��Ce�J�EMV`�*�?ٞ���P�M�������Q����Z�D؝j��t$n)ٺ�/:s���ì��A��ȉH"Vn%�kM�Z�
�I�E���{�9�m���;�I�UUV vH�ʯ\�B����O3��9�^��~�p�a�tx���Wv�If n�V��J��ٝ�[$GI��1�5��ـ-U`���}� �N��=�b�yib�Ij���nwxwwx�.� ������|}E}��~�0�~Q:.�C���m�����'����� ���~���~ ��i�kl��C���c����`e�X%v�>�Ń3K�7�{���|��E�A��wx��６`�*��H����3���?er2�,�@��%�������V�ou�gT_�}��_�@T6Yt�$4�`�]���s�:FWy��,c%`��BVI�!ځ��6�g�}�Ւ�{�3 ��+_D�a$MUU���0}���vuE���K0vvs�X��	�%�4TVE�]���,g�vgf��J� ��� ��%x�$��G��i��80g�hn��n�Q� �v�1�Lh�S�緖
La.	���1L1Q3Q�}��� �%V��U��}�`�e��4��?�*!U��`�*�wfw ���7gTX�,�e��f$�~��h6 p��9n�y%׀nΨ�wvw3RY�$��1�<�@N7��:�����	f,���=�����>�|����M���@ժ�^�xa�As�L�T�SQ`f�� �� ��U�gTX���1�C~S�<{N櫎)��'Oj:���vש5�3����P�fӎĽ����'���j�9����=��`{}� ݝQn��f�Y�IZ?�����li���veaUN��,Ԗ`�U|��ó�w3l'$�nh����l���5%�;�=#��ٕ�M�d� �N���i;�W�f�3 ;$|ۻ2�ղ��JV��C�*��� ����n��Ψ�3RY�S;<\333����O�eC�U��Y��ۙ�p�s=y��r�N[�cm���B��-̜�y8{=����c��t����w��NE�pb�v
�����G �#o> ��[��Imӹ��:�UV��V��:<��Wn�V�n��u�]����@�6(9��\��i����ù��A�F�tplN�)�W����zҤ�u��%S���/R����1A{�ߎ�������L�;<8�4��;ٛ�mN�Un�n�mv��'�n��c�3�4����{}[�jhx���7�]��-�Q`f��ٰzG���W(�B���+ ��E�0�,�����V6~3��� LCG=D�M55�{� ��j;�ٕ�M[/�d��K���h�V�w5Y�;���X}�����,9���fx�w�0�K�L$�%UU���V6 ��gTX����%63�6��{e�ݿM�0naW<�hᚧíۺ���]�nw��d�; ���=��[S_7�rUŁ�jY��U����� �B�J:A`�YwN�3�gvL�_�	Q��:a(���ZY����f ����i�*H$ffF��Z $�*�����F�5I
ː�A��]D5�RDL�KȐ�!%I	@QCB,��A#$D�D�@�P�@�T�&P�Dju��� ȅ$�@��b� ���a$���6�(AlКխ�6'A�!� ��P�(J(ihhJ�J�� �� @S������l�{ [��vv�h�e��P�
�i�/�.�{fV��;3A�W����}�LLHuue����X�p�&��+���~�p+���"�iY��|�n�,����x�%6������?��vwSϷPʺ��w����¼���f���Q���R���%jPM�q$��cOSzF�&`�i��������U`o۫�����p�%�	@��J�M�� >IU��{V6������fg�vg��������e����N�|zO�X����Z0�O_3�GЈ�����y�6���ԠR	���f��ֵ�юՌ�E��aӃB�+�(�
ZJp0�jhY�#r]��������"4G^o �FM���mh���썘�E8�3��`�Ә�*D���4i8��gQ�ੴ{2 ����^tu��̩�1����GV��}�$�r٫4�����5���<�jRV��_Xpja��Y1ލlG�]��Ռ�=��x�F��Pe�HY��bgV�N�C;=b�.).+�ۦf4b�4�,���b��6����_q�jQcB�tw��a�~x��÷����И�0�k��N���ӭ�R���lC%��>�u�*R��؆:�]��k�����)ڀl��3�� %	�{OE:�v<=}=����C�04��z�CҢ�M+�*]u��몯~����H�����`�ݼ\Ľ�_Ɓ�I��#���+ ݡT� ��x��"h�1$� vwc�X��6��,��4B"���榈r��:�)���J��km��[v�pv콴���w��h.h���)�X������XK� ��G3�;3@{��0��Q����%49U`n�X���,��f�$��`O'�6��PV+-��=���@�jY�;��z;�l�v6���Ѷ]�1�m���&ɘ�#�����p
�	J	HHC=�^���n�J��v��i'm��� >o{u[`��,�K0wfo.-�I��x��۶۝��M��x�7/�%����e{Fݹ:팈(�~;�7޸O���֘���ݍ�nΨ�>�K� >IU��1�U�UJ�aL�O+ �[/�w�L�� ��L�>��JQ���)�N�}$� ��*�=�+ �[/�n�6�&_Ε䨶�`Q�#��+ �[/�vl��z��m�B������MU���X�0Ε.��]ـ�>��w���%�S�5N�T�W�����[��L2��Av��H����Ųe{c�m�X\�[��V�J�s�.�]h��6�^6ۨڋJn`�l���ۋWis��낪/o/v��^Þ]ۙ���h8��웊��h�؂��9�S&ݸ�'ld�0tܺ'��9�l��A�uպ��8�Q�u�h����[q�U���g\e����.�����(����k��ImnwK��f/��|�UB�X�wi������"�v���:��`�)t&uu�?ؓT��6��呉;.�����|$�0�G�7wfV�Gڑe�e�hc�۾�I�}��>��2�z{�׉	c~�K���kq���k0�X���fgf٠JWE��wv`��D��&&�(����wuc`�lI,����%V�ctd�}*݅0���ظ��}Y$��� ���`ߊQR�H)]�K�w��뵈6�]��S ��������Ȋ���T�� �O벚I��$� ��ݓ+磌 �݋�{jW/�ۚ�޷�U]������ZQg��.p�!�Ң�s���GTz�b��L�=u����e��_Ŧ��K ��Sf�;3;G�%��J����i�?�,�I�up>MbĒ���If }�4�������6 ����+ա��mp�ɘ�#�n���ln��9��xQ�1-3�2͹��c���瞩#��w�:.�Qǘ��ݷ���]�9���X�8��U�H�$�[� w�����R��7gT[��0n���iu���lN�|��e`�e��ɘ�#��}T�J�RH>�S��Z�lvuE���Y�?53�03<����<G�D�S�L�~��W�<ٕ�nЪR��X'�;I� �와$���u,l��vuE��u�)���J����#��ݓ��n���;�&`�j��IU�t��t[�I���1s�$c6��׶�a��{X�ٺ*F�-�Xn�e_:��M��ɕ�n���;�&}��> g��EЋ����ϭ���7gT[���Y�$���wc`��n���jbJ)�����u,�9���Xǵwc`��,�P�D�T�HBI��`U�>��2�ղ�����$��|R�Z�]Z��1'm���c`�۳�,�K0�Xx��Q��.4c�
4�9؟Bq��n1�JMny҇�B6Ӳ.$�I���k(DDն�:���jY�$���� ��l&'�z�Bi�z����$�9�ٙ�����V����7gT_;���	>�t�R�S�KT�f {�����L�ul��I3 �U�P�
�zhr&�¹����%ݍ�yJ�>I,��wfhff�wuX�sD11��2�4Um�nΨ�9����˻�=��ʽ�߾��8?
�X�Fc�:QI<��E`�������K�A50㒹}fr�q�azr�g���Ӵ0Y����s��y�<;B��6��W[��E�+<�N�`2�;�p-C�n��(&H�^��	
H�q����mh�CMͧ�f�Ge���fԜ������1���5��oOe3FƮz�̭�ɍ�b��OW����N�LK���,�������Ų\=�'6�Hp��|kh���Nַo[ݚ7�_��Dp�o�z�j֋rݳ��ۦ��C��v��v^�;��1]��]]�n���e.v|o߽�~~��z6�E�sQ��{˳ >IU��Ա����l>���M�
�$�7��#��|�d��7V���&a���_ވ��V���;��}�c`��,�������76���9�L51X����f |��ggf�����by��j�/�w�;6L�� �l�X���~�����8	�do+�X��N�Shz�˻72댬�4�tN�i�JG�n�dy�5<HTMf |��}�c`��9���ܻ� JY0uT �/MD�X���$ӂ���
��֭��}�w�f vH��	[WB���%VTUm�nΨ�>���9ٝ�wuXj��+ ���KT��ݱ��n����5w���Ս����	R�<�W�M�
�$�I� vH�I�+ ���=��s��<H�����*14=n܅!��خ�CJt7�0�\�t	�|n{W;������V�ڴ6i�o�gd�X�p��3 ;$|*�^�+TPJt|��yX�p��3 ;$|;�e`�)Dn� N��j�8}홀�>_��DETx2���Y������,�#PE�,5<H�3Y������.�lwi����7Umnʰ��u��ݓ+ ���{f`d��M^�+�I|����w��pl\����v���%��V��۳6MN�1�X]CN7��sm���{޿��y,��U�����yW3,�ڴ1�M������>����{��ؒI����~_����Yd�������J��fwv�IW�{� ߮�Hڡ+Ct;i�o�v��<ww�ʻ�Ͼ����$d���fz`+�e|(t�w]���W����y�a���j����wi;�7�{���6���Xe��0CK@D��u�b��t����Ʒn���vҽ{N���y��Y��h���L)SavSV��;�I�ߤ\�ݑ����;��V��TS�/�'�ߤ\�ݑ����;�I����RɃ���j�������=]� �����n���C״X+�������8����;�I���|�ݑ�c�C_]�j��I6p��f�:��>�R������6� 	�}����ׇ�2�g��ZH�d�W�< �RLLW./A<]?�������,��6��bu��v��7ř@�s����a7�����$�u���S>�u剭��	w��Hs���kf������7��6oA��c R���b.f-��t��-Aa�xa_`�J���4t.�+v6� �맔�k��	�v�	5��jK7E�����x>��;;4;q8sK�ν�{-����my���Z�+mr�d��m�H���)V��F�xv�vyvY;��n6=�9
\�j8�؉&�n�,�lZ�rZ��
[�bl��v����u؞�[�ev��9�l'���b#�uE����ou�/h񬑎�ѐ�����m��nf��������l�M���Kq�8Jr5�=��c[���U��'C��ڢ���UPgt�ޜ�._g��=[c�ۀ�v�I��7VG��Mx�{'kP��WF���tN���c��O ��Y�����/J�����jf�(����t�qny��]U�Q�zU#\�̐���iu�Ke�y�Sq�A�t���r��mvZ�^�U�\�m����8u��<�mM�V��VXP&�L�T���δʃ�Z*C!��BLV�K�YUZ���ݕnCI���E����!�;UUzTE�F��1ƺcv���+j�8�;h�G��H���S�Z:ت��;���J�s����VBj^�klzG :I5B�e���{H�j�seg6�2.�Ǟ�gW,�0u���P��tq����6)d�0R��X�7evjꫮ)������F˱WN�ԇ$c���n.�s�η��m��ܺ�m]]:��gkf����
1ۭ��;�rHh�]2��F��m`sr���[�P�l\�)�˓c���y�3Ÿ�Q����͊�c��sڗv]�ݵ� ۀ<gXn0�l����<5�8�;s՝s:��7n�cq�\p��v0Jl����#��✪��r��YS;`�;'$2�I���V[}$�nNy�`[�m��G�J�g�* �u�N�>�.��krkF���m��"�;n8�c����&z�68�Ԝ<��Ct2�5���܇`�4�As��8��4��5u	�ם�tk��^|����][��3����E�\�L���ն�ԩQ�̜�KYC��u��2+�bz�ڠ2��qʉ�O��-�U �������kO�b�ˑ����M�f��.�Y������ٽ� @H,`z���h|�2|���ڤ��}W��]/l-� �������t�)��=8u���om��v�;3���FΊ���Щ�nS�����H��8q�� �^��H��wh�K���i�gkrN8v����K�Zx�f�{-���;[<���S�Nˮ�ݖ�������<�`14]k�w)b�es������8�ꫩ8n��P�=	�T�pqɪ��U�`z����<�lsT�O]�;(k7f�X�nێm/Ce�R��R��}ŝ��f%ᩮT��;��m���f@2��h+�������R{^}�ؼq��A;bw*Է�񱾝Q`|����͐�ݘx�?W�Е��������s �R_ ���`��/�� ����bX`��+.&��t�E��y,�7gTX�$� �{W����)�����f�:��>�R��)E���5�E����-5�����=����>��~� ;�d�H�&㍵j�&D�5���C�.��J���H^7d�:�6%���6�)��]!�����;��;�I��K_0����h��?�dl��#�l������ub�,���]�='������\ �vN`V�	}v�C&���� �����ԯ �N���X��越I&�O0�l\ �vN`�e���f�]x�V����M�`}�^�Q`}�%�ǵM��6�q�.�rvߕ|d錦�hNV}6;v뫚������ڍ��Ϟ�չݵ���o� �N��>���cڧ�� yw^�i�hꦠij������=�%����(��`�w^�-S`}���M���B��Ͼ�4�~��M$���YT�q��;�I�ꭠ���S_:�E�M�}��xеM���Y���ЧWM�y�GGD���]U���-S`��9�m�b�I'0ݨ��M�}��858���3v�fV�f�m{6;�^{/�n�6�}wBBL�K��C6��$��`�6���l�Z��^�:eM,DS���MUf��S��3@.������٘�zKjĕ&�v�6� 3RW�}T������j���Hi�a���������gh���%����<��r�_�*��u{ll,=FP��!o3�V�@pӝP��Dn�ٝ3�U�x�wB�z���fF��\M٘߶. I�9�v���>��6�8�ym~�mV���V��jѓD��l��mN�J�DH�c����j�)q�
�I�*� �������B�6�w�RɃ���h����������4<�]6o.�cuM�|۰�D���\����$��^Z�`��K�}'0	���ݱ�mp9�=ܻ�B]6�� �S`{އڗmwO�m6� �[/�~��꫓{��=�6�j���ݥ�ڂ1��f㴁*;�sW۷.�8�-��:��Y�����2���m�on�(AzS��W�6أ5�v��T�l3lk1nM�GG��"�q��5��z�n�燶��n�n��ʕi�ݼs�8�[\�^n�ۄ��ӵ�;����z��=����<��1l�M�)�/n�N��Ί�x�Rp�!ۊP���X��WhP�����7�t�<��6#vw3�ݽ޻����w/�n;m�;�9)δ�.;e�>}oN�XH�C�[s�Lg׆U��Zm����W�}	)�>KVs8��	J�>M�7?D�OLVuw�}	)�>KV`��,w�^s�4Ѫ:��Z����f���r��67Tٮ��*�>����W��A
(@�t���h?����;rE�3vL�7Um�ꏭ���5�;{�]�K��&`�e�����~L�<��pkD:1v�Bݑ�j�%�nx`/[��E����Ɲz֢FL%@���X�R�7R�}��p>��U�-[T]*�v�0M���&f}U�|U;ۻy��N��5��G�J��%7����@{����a��fj&f� IW�$�	wh��%6�՘�?�����h��h��Ùݙ��6{�� �wt��&`�p��[��2���?��Wu�}����wf�W�$� �X����qB4�FO�1D;b��;c�71T�pci��q��`AEdCb���W��ꘒ)���$���`�e�\�<�$\���v��k�!��ڶ_?;3�3D��V�]�`oږ`��-���>�S��4� �����ȸs���~� �.����Ł���;����6G+������v��Wb�N��.s� �� �와o�Àv��x����Ar�Hc�\{�f��ۛ����p�)JL �8�b-p�^\�۬s�N<�k��v޺��L������*�O0��|�7c�;sb���3 ���J""����h�������亳��]6��f���� ���
��"b�������IM��jY�n�"���x�����)R+_7i���3 ��\����~�U�� ��,A�ꯪ�����4���k�!;�� ��E������9.���OtX����������鷳d[��!�pA�ڜt:7m��Y���k����#�����-�ƚ���ؤ���3(�ظ����&�d�Tٻ��}�~���ɘ��\ �ݜf����!�-�|{�f�� �����%�	������ZN��`~�����X�{� �Ӫ,9��wfw�-]�<:�!��*j*��3|����՜��|���~�*��T�IXB��(�� 
��`�4%�HH1$ט/�#�r�7EAZ(�S��u�Mxl�1��xw);�X�w;�rv#kwc�s�;8'YᲴ9�F�Q��8�ٮz�;&��B��讫v��㝚�;s7'
���ck�;83v�d:�T�{^��AM˂Lq����m��v8���LG6��=Vn��@���N鈳֜g��Wfխv��e�p�\��ҋf��iy^��v�>(�U�f!�	�"|憗{�^� !�P^e�kF���m��1� 0
A���,�Q�wND���u�۟L2�uT6�Tzm������@��٘o� 3}'0��# �I��|�l��l��틀���}����Zb���j�O0߶. f�N`��p�f�U���>�S��M� f�N`��p��f�|�_ 8��/~C���Z��� ��������;~ظ��s ;��H�WAB���'C���a�1v�;�˧p[�d�{Gzt���t_"�N�X���v���g �{f`}��'���R_ �=o�2��7R�^p����TB, FL��$@$�j�� �Q><<���{�Uw��9�ڳ: L��tDEI@�UU`v�^�Ԧ�߽�0ڕXL�aEAE�t�tb��9�z�E�7�٘��'�s �=r7�T�UI'|{�Y�s��F����W^픢��g�����[p��ʞ����p���,�Й�ѹ�\eg��i��X����x�>��^����]�`���l��� �Wf �[�9���������^J�l��ڳ���5wU�|۰2�"f	`������)E������]363�x�:<#��V)�5�@�(�޸���D���І��|�`c	E[7�f���6f���5�����%4��~�y�F��m���Ĉ"���M���]:"���m$�b��Nl�f�����|'pvV�W��އ{��t.tV���iFֿ�Fk����`��y�A���ԁ��tj:�p��ES� P��#�2��Z��n�+l��	Q�>�)�Q���=�.����Z�M:֐:�1N*6��"�Q�6'j!�'��~z��
�u��z�x��>��!ꫂ�}���c�w�s ݎU*��Un�2����gv���� ��V��^�R_ �=u�Q��v�&�$� =�> d���={"��l�v��UiK�7n�8����]-֥4ųz���er��ڝ�A��Ϫ4�q[p5_m����W�z5)�7�j� ��V��CJ���b��ɺ����ewN~;�Aڻ�0g�π=��ߋ���)Rt$������f {R��c`�Jlk�T���T��O0�#�=�+�=��r�=IY��x�J�ŉ]A*@a!�:[5�:Xt��2>"t�@\����꯼��|oe]1�	��2{fV�� ��f`�*�;ޮ�8&\ �fb$��x�[p��S�ۋ��%��=���xٛ��rn7��}�n��+aH�m�	���7�٘�#�=&V��Uc����N��ڳ <�����65)�gvw�;M�O�T�$�UT5���V/%��ljS`o��9���hu�L��D�5UVݽ��ƥ6�ڳ��f�{��Ͻ�Q�@4T�c`���j� �J�^K 7{��mچ�d�iY��n+s�N�\WB3yTS��� 9�ݕ��N�.�q�bco<<݅���ås��8�
�Z��N�x8��On4浸��m��9�񥋲�ك`��

keX�tO
��g�j�n۰p�ˮ7mu�㝅hف{���-������Yj"��	t�e�9+{r��S:��c�]�]It���r��L]� ��g�5� g�;^�Ӎmɪ5��q�	�t8��͵���UcX�K3�bX�ID��c����Í�Nc�mg��3��6��oH�m�/^ӫ;a��v��p��ם�������ڳ <�����fo�.�5>�~�Ք� ���O0�G�2zL�od\}홀H��ꏮ��������6��M����Z�0{��oz�ѕRS�4�Um��4(]�`yj���U��䱰l�4�Jhj�h�j����}�0v�]Հ|�� ��.7oj��M�S���IScE'MQ�A��-��Wmy.�Lks�k�c6/BcG�]^��t$� &��o���%���W�VXzl����O��V��0.�m��Ͼ��΀�"�R,M "�	4�ҦX�{�Bt4�Y0�f"��I���ZGY���x�ЪP3���K;��
/��՘ �*�K��wB����i��^ȸw�3�6䋀f�L�oƨ?�RC�I1Sa����嫾�wt��K ے.��'vST�%n��nH�o���6䋀w}�0v|��J��r�Wnq�mGɹ���]n�픉�H��Z�x;&	����j����{��e`rE�;�٘�%��z��W���."���6䋀w}�0�K���+ ���}jUӻ)1��� �{�]U�����e�!P B�
R^� 1�SY߻��� �=oқ�Щ��	<�6)/�f�L� �#��l�U_ۤ��̴MMTX�K �g��Հyj��ܑp�D��t�|��@������m\u[l�6&z�us]�ں�6�l&|��:e+�]ӧE[M�`rE�;�٘ܑUp�I��m�mA�ZH�Zo�w}�0��p�I���>��*�vST�%n��od\7�e`���w}�0���:��k���-��kD}>J��*�>�j��ғ;C�Z�lHm� ���24:5�(# �Z���d	����j��݅�eT��-o%�����U`}�՘ƥ6�� �geɢს���:�=�]��%���U�Ϋkڎ�Z�s���ۆ�7�В�T��t�1����~�3 =$| ����� �=oқ�И�`�� ���;$� n���홉��ݦE��� �a�ff(�wu�G�(��ۘ�ڦ���a�ԌLCSS�7wx���}�Y�}	)��͜��r'�+t��M�w�3 ����j� �j��fv�ׇwx�hN#100S��ߵkWZ���f��gkX��ƍ��ԧ<|�.y����{V��[z4�m���q�gnv�`MŴ@��UӶ�;��2t��ô���
���y�o* N�� ��a�	{<���Ԙ�2�n�ѹ��e-λ9��0�-:S��òA�Z��ѩ�.{W���,���9�FI��֍���;l�n��5�޺]X��ճ�<�W(�Eq��mR�P]�w��w��w����&��1���C��d:����2�14��<t6�8��ۏ.�O"+�D�U�X��$�������ٳ�����홀m��%���k���$� 3�g0}��w�3 �Ȧ��� �t71�RP4���7Ww�	.��{V`BJl>Z� �f�QLDTA%55UV�����]������� ��|x��>�+v��U�ѩM�g����UX}�� �n���|�q�����OB��� �&��+�^ާ���օƷnCz��s�u�qQ��5U8��u��UX}�� �5)�;>�u*����N�ğ9� ��|�U�T� MH�$?"#�N^����=sb�{�s ���2��]�]3D�M��۫0�R�9��h�{� ۓ����*w��@餙m���&�3�J�F���j��?�L�T���M� g}'0^�\����>�Jlgww~[�7@�4�Q�9:#rk+�1uں��-�od6���F�swd����"
�-{ww�<�~���w߹�>�Jy� ��׀oJf��"*"b������{Va���]�`}]Հz7b�TO_��B�v[-�	<�;{"�W]�����
`��t������0,���[0�6p�6m(��X�J�x��*y�ן�ʼ��u�^�F�)	��G*��4?�1f?����׀y��`{}�0�R�S��O�LE5FU����S`s>�]��zt������)&H& ��瑸ڎ:3��k�i�-�6�嵬��WӍ�f�;�Hr[�n���3 �싀e���n�p�ī���mP:i&�<�;{"�;<3�B�ՀjUŁ����fv�:W#�5S���M��.]X�i����v�b��IWR�V*\�8�8����h���s�|���B$ҋbFD��*c$�2Ld%���~����Wk��Ɉ�I6pw�f�݋�v�6<��_ �ݢ씕��� T�<��m���y�*�:ΧY�w1������.�<���a����m�7�ov.������pw�f�>ZU�R�JӢ�&��9�>���)]�y,�>��6'�u,e��L��xul���LÝ�#ЗM����V�x֑����S�SU}��=�6����gv�'?_ ���_�N���4�-<�;{�p������=��}�߹�i#��Y�{!���F��0�Ýh{�Hp�XC��[�ųKkFj.[�x�<�9���32���'$�!���	��đ��}�9֗� 1�ή��0�j5+yhkc���M��Y��բ�u�H�y���͛��@� !��A7�����˭pC^�� �x��\H�s7�՚��Ȝ��!����sz�б��bFdZC�,o;�Խ'h�JT���[�hHf�H�8��f"]	�O��������㰇df'>�x��M�HH_j�/��U{�Pg\���b*��y-'rh�rU7�z�GQ�<���t<�}��B�36i���N]����Ÿ�q.smx� ��s�|J5��89��M���;H��H/=���m�>��{~  Jv�lq�U��E�ۍ���NW�˹��ks��Þřm��S��!ҡr�n�%�]��*[=�%[=�t//"�/GZM�y��������B���۞���y�5��n��ry^(6Ѯ��l^��Tn]`;!��v�z��s��$���6۰:��a'�z��`3��Pv�5N�9b�m� ��.|^ka�\���k��n]>:�nwd��P���6^ƺ,b��� �q�7l�W1A��.8�a��f���nNHP��yM���h��Z�s Ur�%Slk�*��6�iW:J��nb�/ �J��N(8۳� ,�s�-mf�Ƒ�p��f�r�Apn� ����	��*�Ll�e�$��T+g�b�����کWl�zƺ��Ϋ��A�y�� ��Y�!�m��K`�N;)2sM���p��(��W\�j��s�X!�)T����Gt��k��u4�g8yԍӻ:P6�M��t�M�*	v�kEIukN�W�NhQԶ�ط<�e�ӛ/G+b�Jиnb
E��N)��eZ55�WA�%�7j�mo4��n�{�p;��a�M��ۮ$��Ꙭ:�ݜIf�����:�u]u�:mۋm�C��([��c�x��0�q�.c]�5����5��c.�r��-L���٬�n�g6ď`�u���z8�vx␶1�v�eY]�n 3�gf�ow�Ǯen��/�<R�[�q�Ȝ�#-��I���q�Q�<.n7Q�{N0NX�q�v��%�dr҆�/#�wmL;wG
���!qIc`nR]QZ�-S��9ny8:3��D�܁���r�Z5�.03��WI\g[3�g�Kvy"c`!�$���q6�IFYڈ�^�{S�%���8|q�=[��m���\�h��hL�.Y4u��h�s�4�mg�vRM�t�4q-(
��!n�e�U��m�N�9�BD��UC�b�@�e��χs[�qK;V�����lޮ"��WB�`=m_�tx��v�=PzTG�=ASg`!ۀ�<YF(��t� ) ����v`x,��{3ݾ7��O���:9�e�G�F8��.2�3�����g=��c�&,��E:9�j�p���r�GM�^d�'λd��uv���a#�qi�b��$\v��z��4v�{��ED��&I�q�]e��ŷv+/4�m6�v��t�!\�� �a�$e����t�Z<�ֱÌ�ty��ۊ�][�r�"�X�r�fg�ue�]�{ߏ{���u���|���MW5`k��<�9�l��^���]���l��H�g,�N��ݻ�=zJj/}#�=��{�3 ��E�;��1��S[1swu�{Ӫ,�� ��E�;}��R�eZbMP�5U��Y�}Jl�fx�G����]|C�[AaC�[l��`�H�o�#�;��
���I�V���Urȩ��&bjl��J�wom.�۽ـ}�63?p�n�i���x*����,c�"�v�u�r�aY��s��΁Ņݷ��i;���4P�e�q��j���{ޓ0�ڧ��ٲ���a	�ix�i�tn�����<���d�P�G��\�����|����[T	�V����틀v�$xo� ��&`u�`�R�o���[k�v�$xo� ��&`}����]� T`��]��{T����338>��{�����d� 7��T����X�^��j��Kk���;���6��׍�upmf�yHH�SLBe��e������ �>�|��wg�ѫ���60s��=[h��`}���d� ��b����x�j�Ym[ae������y�����F
��A"WB�T,��aҳ� �U�����a��)�b2*�9ٝ�=:�l[ݘ��U�ۓc�=zm"��I�]5m���3 ;� �ɱ��l\wn��E_>H����ضc0󨴯n,����F�1�^�m�7#��c��N�1|5�Z�v�`}#��6<�틀n�L�6���N�ꪞ�"jl�-U�����Ʈ�-����S`}�Pɢ2 �*�˛���틀n�L�;~�pܒ<�3�J:E��T2�mpݓ0ߤ\�>���^+��1� 9���PC�i�\xۭ�X+��Zo0���ܒ<�틀n와OQ��Lg�b�SkcIv���[�v��7�0�2���9�{K�Pg��m�=��0�}��D�<�틀n와�eO��Q5<�5FT����������'w~~f j����I*�h�Є�4��SISS`%�ـ-U`zJ��j�۲��b�j�:Jݤ� ;6>�G�l{T�s<%��`
D���3U=<8�|�$� ����7d��� Չg߀��UnK� �c�����d8�srvG�6=�,���Y"۷�yduN�nB�vPav5	ɳ:֛g�Hѷ��63�c	3�$mY��J^B�	
Yݫr =rl�<u��Ӧ��%î�IYj��p�&���[F�O!�nyD�g�5!�O.ָ���+\wn���F�Bٻ'g�;8�Sscٜ�d�Y6�ͷF_�˟�A�[s�Wg5Cr�;�����)0 ���&:V�!8"83!P�2[�m�-ۭcv�	37)�gO\|U��7WX �uX�,����=
H��gʔ����T1����L����=	%X����ٝ��Ɏ�%����H���wuX���>w��' ݒf��]Ie�V�v�u`zJ��� ��`%�ـ	j�*}�us���>/|x��p�&`�U`zJ�ffwmn�,h���~��zg��}J� l���*u�t���k�z޻�L�-��T�_t�ˢ�k �~�� ��XBIW37���,K�"Z�r �S��/8���w��dm`$$�A� �@�&5���(������>�}U�����^�와v�+uJ������|�$� ��Qg;3D$�� ;WU���)d�K�`���� �:���Գ �U���#�6k>T�D[-;��4�n와� ��#�'���}f�R��8.a��u�5Զ�-�ԕ�^K���������f��'���v�Όg��5��m�폀v���e�ݓ0B�}u%�M[ti6�nIs�yl���f Ol|'�۫�)[�2�_U�����^{��uՇ�x a&$ID8��R$o6��M���" ���}�|���߿o�6�o�_t����n��d� ���od� �[/�n�%���� ����y�K���+��G�OI��ݓ0����$��6�S��D�b�l���V�����)SAݳ�:�N�;�̕�w��mp��='+�{vL�	� �ER���|�q�<H�̫�۳� �G�2������H[wc-I6p��3 $��od� �\8�x�K�C��t[y�l|����_}���^���� rR�d�Ъ_]l��n��$� ��#�$���f I���Q�J�������\���{h�oe'��]-Ӎm\n�m\v0��m�u�p����'6]���_Ł��f %���� =�Հ(By%��C�uwV4���f褾ےG�n���|��T'I[�O0E%�ܒ<v8pݓ0�lM8zf�zxi"�l9��==�Հ%�Ł��fU�K�ݸ�VZ�_�\wX�Y����c����5%X���
���՚ݽ����h��ɛ�4�u�Ҡ�)�W�{�Hڝ!����M��Ɲ���-�k��."�7H�������� � (�O9�F\�z�;�ݝ���Cn��>ڧvI�]Y�-i��B�=�󓐈�u���ֹ�NnWrfl�+�Z�8�X�ּ�g�v0��K<v�`:�,���]�t��̫rМ�ط3�əl�]���+kf��浽iT�E�T�l�oNe��kp�����d�n`M�fF7M�>�c���盷�m�+��.z1a����m�_�~~f�)E��jJ�iݝ�����;����R���Zo0E%������R��vgf�7�ixn:�������=�� �T�9٢5.��7��,O톄�4�H��uu��n�� �L�=��;~���>B��C�ucL��ɘ�H�o�#�=���}�o���O�e,Un���kl�j%��㎆/���ۗnM�9Nأ>�J��+�i��.�������;�0e�M;��Z��t�mp߶M��>���H�j#�J�`j���<�(��=�-͑,�5��uWX]\X{R�g<�(�;~���j�Z�e�ӺI6p?3�G�w}�oOtXG�*�7U"�_�Qt;�CI�i��=��;~����Գ �wfn]ђDKI,�"8�(L�A:#�&,z^^�V[ ���<M�*��LvSV�U�ۼ׳��n��l��z)/�f��us�t"ݔ�e����Àw�&`�K�|v��<��|���t+���g ��f�~���.D�����MJ��q�Vy<��3w^5D�'\ﻮɬ,���q(_7��٥�{��`/}�U�f�a����Zz�t�Q�E�:$4����5#%��ě�-݉o�Y<���I�3���d�3����W�����1&eo�q��|�����x����)�L� ��Z��*�R��R�r/|��qGp�y���e�Ϸ�v��N��#��	���3x�م���b�u[�.����C�Q:�>��G@8(ס��E��
 ?	pSb�!�W��,B	��� ���چ�� =�@��/3^����R/��K�<CK�31Q5���Bԫ ԩZ�`�j����U���J������ÀI�f�I|{!u,�v��CwI4&���a�dZZ������q�[�q���ڝf��2�~@�p>9����ÀM�3 ؤ�/�G�{v�W��ZwCWJ�8�K3�� ]=�`towV�R,f���n��M&��� ؤ�/�J�5*E��R������D�@�UUQa�;�Հt%�`-Գ����9��L��^~�_��U�o�r/���E�,�|x�ظ�&`�K����{�Z��A���)�m|g��n���Sij��-��*P���a�v���͗�T:��V��l��O)/�K�#�%���=�/��v�;Jݪ�zR��vgxv��{����n������MMC�4K��LETX�Հ%)E���v`���Ld��5��uWXR�Xu,������#�=�L���]�Ӻ�4�MԳ JR�G�U�%)E���;�;����0�)�
l�SϿe��ߌFcbvۋ5uHݻv]Ʊ�,�..˫R%q�<I»n��v^:� C�v���ch�i5�̸����ۣI���5�l�`z�M9����G6�؟������풹9���>����
��r�3حM��v��{/������ܮ�y���ޛl������;��Ғ��'����[����m�Jwkml'�;�N��v��')\-��f./,X���g��=��{	&���J�Ps�qQ�j۷���B�*v�l�Sp0�U��l}�+�,IV ���K0�ix��[�m��K�����K�vL�$R_ ��K�wB-��e����ÀM�3 �[/�K����	�e$�CMD�X~3�r]�`etX
<��崋g��9���"F����}�&����Iٮnɟ��������8�8�RǴ�V��dz�8�.ؕѽ�����QZ�q�S1�}xi���G�U�-���[�g;�;3�|����`v����X%�.ꮰ�J/��ٵ���ݙ��J�� ��S`K���Ԋ����Zwe�j�w�&와z�E�%͑��K���A2����������fh���:7�� �R_ ��f�U/�B�b��+mX�J��J,��`���@-;m�^_������8�ݸ���ۖ�KV��Y�Av�Nۘ�݂OoQ��8�m���� �]�`-Գ �jR� ���cƼ�/	��$*&��[�fs;D�l��� =�U�;D����/#MT�f����Q�a����@_i@�È)꤈=o7��r�߿of o�aMMC�4KS��M�;��N�u`]�`-If�IM��MSLa,���uWX�J�$�`�Jl?~�����_��$Cj*�L��WC�N�AR"X��V����ݺ�غ�������l���jݴ� �와z�E�쓘��	��R����I��y�z5)�w�.� ��V�R��x�!�Y�CMS556��׀Ԫ�f���ـl.�1>��h�*
�����vg���V�ݘ�R��_V�2�o{��s���/]F��V?��V4� �와z䋀�'8�~�t��������ڢ�nm[��7���N:�e��Y����nj����w��r�Y˫�
�+���`�"�vI� ݑ�nɘ=��i�Ϊ�?��:� �RW�Ԫ���Y�zS`g�j�%�Z�{����Ԫ���Y�3Dlwt��w^ ��4j�"(���"�������Y�zS`jJ�9����pKLs44MLԑ5Y�zS`s���wu| �uX�K0fvv�;D�� S BP	�'����e�Ǽ����
���8�1.MF�r�����zq���l�h���;�>�w<��IaW���״{&�얜��\\Z ��+�u�E��l'�н���P������=Y��7�Z��d���^%;m�3�M�\�2p��RK�c@�V�'ZG@�Փ�X\��[�#q�]��q��sd���;��N�m�Fl��5����������t��G�fb�X��Q���D4��B�-��
�:s��+�Nx^�d��l�c͌�ӗ���!S�M��Wm�/����<�����j]�����@lwt�sꀞ���"������ �J����K�0����G���ߑK�c����� �와z䋀v�H���pz�)YR��'V�e���d\��G�z�E�=�&`���ӿ�U�]mp���� �와z�E�7ђ�\N @@pQj��(XڰjP�u�g-�f��פ�D�:��n�Ed'*�bdZ�0�۷ �싀{vL�={"���<z������M�����~�>S�g��9N����f�61zl��*�=��_4A��Zc�h���"j� �]�`v���%�ݓ0oԴ�P)6v�\�$� ��/�n왁��f���,��LOP�D�PPN\���)E���f�)E��$�`��������~���nH4rzfѺ�л���:���C�u��s�.�8x�����׷>�?]ـn�Q`}	%_7�R�|�M�4ڑ���9y�>~�q������|wd� �{q�*�T����W}���}��g/�>T!Lc0 �3,�V��U�p��b�30\�p�)��Ub�W�*�����X��`���s�<G��� �i�Z*f���"*"jj,�K0gf����.�vR�/A����wok\�(����r�ǞD�ά�m{W��Su�]�4�m��5��# 檆o0\�p�$������3 ��J�U(L�v�v��vI�uI|۩f�IM��s�'�a���)���� ��Ł�Գ �jS`$��'��Bc��O�%48��������ʻϾ���_�}��>�<{��Ł�nM02!��")�����Ѫ.ےG�{c� ��3 ����dIO/ Z6Q����J�\zɺ�U��mvGR���y1��(:H��R$�l�>�U�{U"��Գ������6ԣ����h%������=��|��$�� ۟�.ےG�OR*EcV�c��v��pݓ0^ȸnI�!���i�6� �싀v�����7vL�=>��*�&U�vR�mpܒ<�8�ɘ�d�*��ID�^J�d���;7%�}����vk��Ü��B)���CȰNT9�qQ9P��R'E)�k1�x6�x�у�Yb�Y()JJii?<6F�?,C�6t� �!�uSg�,�����$ʝ�y�Q�ۣE����X�X ��V$bUK��LA�a��e���l9��g0��u�n�T��{�}�ޓ�,`H���T�KSI�汷r�ysf±,4ղ�#IAIEX��p�[��r&�t��d�JHTQ<�)�@N>!ƕ�7wwF���@��e�K?}rbi�<B���Rq���gzѰ%Z�~��ĐB��V�0��}�.j�^�n�����}����HT!'5�4�R}�c����,5�#���m��<��0\;Ӭbӳ�c���P���1�u٣~�7��{��>�����C���e��j��y�����FI(�k�H�<=����n���Ѩ�s�;��pa��L�Ǿ��a&`2SP!�� H!Oc�K��zKo~?�l�m�m��e6��A�Yd�!�����S�F^�2�c
d�{X�,.RX�,�:P1]����#Yz�B6^�n�Tyq�kGBE�탶�n�Ո\���ix+v{9Z�6���l������'��l�[����^�k!�[w�6�t=�v��eL��kN�QC�L�ݳ�#��Y���])���x6��H:��,�]ֺ�9�f{�Lv伜�0u�"7u��pkg��4g���8Ӫ[�������2�cԼ-����k��$���}����E��=��c�Mt�Na���Gh��g8m�DV�u*���@������j��l��8���%Αb5�4�Eib�Nlj,��V�Z��ayz  �%�:�#"�7D��]UR-V�kg��ڈ���P���b��Rܶ� ��Ҥ���6�#EI�( [�jͶMwi!������V^n2�i`� b���Ui��!t�F�.7��m�eZr�ܲav�H�p���-��˥s:v�{-��u�!۩�q�n�[mt���;l��������싎��m�5w;���3��Y�֬�JQ!K�m��,�F������������Q�u�lSa6���ORգ�fј��=� ��ga%d�����y��wk��`.��\\����N��F�y3��d�e0�ɍӶ;Y��:l�X��q���Hp��6nX���#6�f�v�b�w<Qe�6
6x9�
�um��d ]�bn3u�sͤ�]�u�tfN���.��W����Z���Qn��:�L���*K�P�=����Q���[1��vx�gp1�09�Z�v'�÷��8OU��nیp��$r-��Jl�17gf}ħh�zv�[l4�+#�g��n2t ��;2I��5K'[f+bĉ<�0e久�.�`�unC�N��� :��B�L��7Q�3�N���]���a�t�UJm��3���2�m��p�	mr�6��UPCr�TtƮ�X�%cn�k�������GV��*̲�4of͛������v������=��WH*~G�;N��<+�zm*�@�v>�A���f-�S�@s��,��(���u�&۫�P�H+�۶^%�3��6m&���0�w[��v"�p�[��󌵺C9�u�RA\��#�Y�]�l��R������m*�4.������^�d��J��M���r�ۦϦx{��x&I���U�͋qpg��6��Y�r�s��s�;���[U�ڱŮ���,V��E���0Hl�XrN�,XR8U.��):���bS1IQ��B@�۱X�0#I�lnWA���R�Y�,�#�q����nA���u�&��n�K�\O� �S��ݓ0^ȸnI����_\�u
�i� ��3 �싀v���%�	SkU+*WB��v2��ײ.ےG�{T��7vL�7HӺA��t@�\�$� �R_ ��3 �� �nܦ��Ub�\����� �R_ ��3 �� ;$��$ڹ
m ���_���>������T�.��\�1����8\�]��jr�e&��۶�wv��N�	'�ـz䋀�N`�K�+�A>@�V����������DJf,�p@	Bcy	��h�"l�4oi�;n�;@�D1
����y�^��wR��gvh�y�Y-�M�1U6��׀{e(�=��`�Jlo��d���4EAM?E�������R�� ��V��]�X��#�/V��;�� �와z�E�;{$x_�~����D�Ƞ��~���P��P㷎���*�n�c������`ݗng�'��k;q@��v2��ײ.��#�={"�L���wf !":�h�j`�
���ԕg3�4@��E��wf�IM�DR��b��Z�����)�+�}�
xHD�%$�.�,�;����M�o��x�H�*m62بM;�ݓ0^ȸݒs ��/�d<A]*	��lM��=���R��)E��Գ ��;��=�ݶ]��G�dt�q��'��u�=X���d=u� vs����ط�����xޔ���jY����17���&[��>7�`�H��d��틀v����ޣ��*�_��i���3 =폀v���ߤ\v������������]V��u`]�}�WBvm1Q�fb��1��A�j�\!�]E�x�	�ff BB41֩�]��nl� �7�&`�l\Ol���]�.��2n4gi��]�7�.#��n�=������jQ�X�8�"�p�v������3 ��b�f��JElC�N�lT6���3�W��]�{?.����xo�.��E/��i�6� =폀vk��ߤ\}�f�|��U(T�mi6�f�/ ��E�7�&`����ⶕک��n�I�|��� �l���vk��Τ?INAE�Dc�8N�~��Z�$�[=�D�L-pv����ݝk��0��lv���V�O'����u۬	��m,s�Gz06���{3�����lp����cs�r��.Cf�ɰ���Z%#�Y�{O��_t�չ���� �ksu��a��
��c�gw^�!��v��y�Μ��Zr��b��u���Cḑ��V�bma5���@]gP��-��-]��:��-1�T:���[�K�q!9P�?�q۵���+�tnܚ�d��U�;6�=d�L��.6����;�����w�����j�崔`B�6�yH�FZ��(����U���]׀z;�l������"c�Z�Z�!ɪ� �.��=	)�7ږ`�U`n���	jkp�����R�7ڳ 7R�ggv��j��;ZFi�He�P6�f�f`쏀��������{��̑�dh!��"���Y{d\����l��ƺ��=،m�Y=^ܨi��M� {� 3}��}8o�f� �(+��m��4� 3}����]흭�홀������ـ���$���R�[e�c�|��G��Y��;�4A���嫯 ���CH��*�]E�p�l� ��> f�g0�8pݫ�DWE_ʝbv�`���wvh�j��ou����Y�l5������,��ӷZ�ZAۯ��+]��Nb��q�'q�����j��j��%m`f�Vs7���h�wx�0h%����� ��[X�%��� 3v>�e{u�-�n�$ەh�~� ��M;�V	$	$!׆m�`l4�=6�^�o�l��p�u�����N�iЛ���S`���Ϸm�9������6�!�_�T�U���n��3��������{��@��:���K��lMݎ��Թ4���If2�c�7C']��=�O��֧BT�֙n�X����NW �zL�{Us;;�d�]V�7b$yxM�2T�X�r��gfx���� �.�>��{�]� �:.��<���`����{m���� �ȘU- �-NC�UU�;��D|�U��Ψ�3��W�����h1��h4��j�U%I$M���N���~�}�����b��[�������==�3 ;폀� 3�*��+���vx�ѭ�͛u�Fz��I%!Z�h�:�w�n��l7�)��
V��ݦ˫b��������틀� ίm��u���
;M�Bo0߶. f�|;� �MY��n�'@Hs�T4�MM�|���ϽZX�՘��S`$�12ɨ��v:��ǀw���3�f`�l\ؒI7��]������`��W�g�V`��Ͳ�� ���zwb����	IP�G�z���o.�{�������#�G�l��h�#R��!��f�n^�oF���m��l�=/�`p�j}��u�	��0DH��ڲ�G)F0�x�ˋ6����i�r|3vǵ]K���L�]�v8ҳ�א�v�ڍ�/S�.2`	%�t�m��2�x�'G\hxݎl {��k�����j��F6�r����;�������6�V��OG<��(�m,��y%��Mk���cpf���ζ�l�ȗ�'=3h�h�99�^�vI�J�7QH	�U��w�w���do��zwc�� >�]��M1�CC�S�Z�k�e���ݾ��3 �싀w�c@b��N��|��=�K��0^ȸ^�.�e{VІZwE��M;��0^ȸ^�.�-����E*����m:y�z�E�2��p�n� �͙�]n�F�g:.;ny���vr�T�v�'^'�����li�ی��lC�޳�;[=5nY���-���^����p߷W ݨT�*�NR�W�vp�~���K!�$ybWjf݃ۖ� �jS`d}�o�ݚ ����)\�ut
�N�}�~��$\/� �����zQ*t[VҚ�В�#�S`{ӻ��{�}��(��n�!"���}ظ�}�J0�˳ �$��>�[FL0>�a΍��u�m�ɶ����n�[�m��m�gq�@�t6W-�l�EV����{���g�V`�������`|�7�XSn�5Wl�N�w���Wg�H�o� ��up�u*�V[��t6� �$����T؝cC恁�fgvL��r¼2�q�%�:Іai�0TH��)+0��8٢0B�1,�Y�J�Z1�2A��c�B7*ݪ������(�!��"'�(`bU�K�**����L�"��j(��0:$�x�w��dxƪ�L!U7 8e�I�l��c�N,1�'��+CuT�H�
C�i)!���
cpu��wq��M�o:I..A�P��aTSA"���ctP�%1�h(�M��C��l3J�"���HQt��%�/��hQ�i
D�֖�/�}֔1L��"�1�I�$A�%e��������uq��|���HM{�Jt+8k5��$�N�i
��\�G|�ӡ��F�0i�_sL1�# ���ӢC���Q쏨	"pn�bSE��&�U�pS
%�<OK���^d��Sw���iH:��	 ���bB���k���p��q���jUv)9h-���C�4%�0�fIY$@`��4٢�����U�U7����\_3�U�T�Z�ib2�M}�Y1��=<ø���J�f��A��� �� �ЮB#x��v��R�;8:z{4> �x�v���(�#���=��Ƅ +���ʾ��f`�R�W�16�J�\/� �{vl^՘���ѳ��`rm��ও�V:Y|��6�E�2{f`��hw��:���do��Z�'3�E��@���àu��N7u��s�6�a���An�Յ*���=�0^ȸ_}'���ݲѩM��1��t�����L�i<�={"���|����2{f`��G��:��Q�l�9���|��.��3 �싀w�-\.�}b�\�
���=����9����]�a�7���Ƃ	%&��*hƠ���(:.q5���PƀH�_���}��:����Y%��46����3 �͋�gW��_wW ��������T��ֺ�Z竎�W�%�:�^׆��\X��g�q�-�c)����]�3TUf�Z��ϧ�,G۳���v��S���P��5RL���yM�<A�����v`��l��(*�[��ư�H�Ol��6-����q�������e�ؙ�>�]��˦����l7�V/�TVU������ �݋�gW��7v�^՘�08�3��t��b��e*�<F�p��rv����9M�v�D2����`ڏ<k��Dn;Rj��u4H��FɘdR5�Ht��:wcl�N��l�h5[�dmM��p�G&��f��Ӻ�YNU7[DuI�v�枈�䝞HK�n2epƢW�2\Zy�R���d��@�
sՅ^��DH�s��:j�Q��}u��_��>���q��6�=aBK�U,��T�U�b��]X��߰C>���E+#�qIGL�%��l���sz�]�̩�4��Ǜ9���ؽF���S���� �ݫ;ڳ��	t��薎#%������0�X��0?{��9����$�6y1w�1~�K"�j�����ـln��3�� ��|6]AU��P'i���y�m���;��| ��|'��g�S���v&&ВMp�z_ 3w_ �6f���h��??�II�ڌBhN��(t�Ź^��}��kn͋��Nہv�g��e���J��3��ܑp��0�ظyz_ ���YH_��_�i7|&����?f	DA���f�s\��M�����g��*�;)/�CHwj� P��=>Q`ln�����%ـ?�'r�'S�m�4vw��<��K��BJl�.�hc�	jkp*���:;�l[�0	)�3��f$�]����&��T!1PD�O�4���> .9a�v�7\y-��{.]��;��ɺ�jX���&��?;�?3 P���ذ6�up�uWH Rv���o0	rE�;�v���7d��]�}�9N�Q�T�In�����?{�Of/�tNC�������~��~��uX��ɉ��DUT�E4�u� ��f vH�un� ���YHO�4��U`-Գ �w������������?юc�4�?V�v>6�#��ocu0{pm-.��Z�9v1i�\�vz�e%��ii� I#��| ��|M�0M�;)�*�[�R���| ��|M�0I �M�VH�y%��¢�� J��,���ݞ��<���1z�,C
[4�,���};�a�f�bhgf������a��15ׂ!خ?���.�m֊�Q�NӶ�m� IX���IN �%6n��;�{W��'r�m��m�:@��ks��m�vu���e��!�[�l��@v{#��sɊ�~ �$����ٰ;u,�� ���m+��.�m�V�e�\�p	�&`IU��n��3;<A�	@�K�&��b�"�l�.� I*���#���$��������X��Uc+r������wU��n���6v�� ݍE@�?�U��*m��~�\owW ɻ3
�߾�ʾ���1�20"%'�H0��~-.;���1ݭrͬ�[�A�n^�GZ�N�}Wc;W����pkE0F1�=�r+4nP#�����P\�9��t^�H������L�ۘ���F��W]g���n��s�f�,���	��_�í�jݝ�E���m\nPl��`�u����6۷n����M;϶J�ز�m����4Dẫ�8�qv���r��z	�lV'Vn����rBԒ�T�9M��*�������]	�^�xֵ�gs�n7n�nCn�:9"uf���j�䖦���p�]6-՘I[p�z.�W)"��5i�,4��r]�I[X�cwf��P���D��N۶�� �NW ����{��zl���Jr��VէJҡ�\#|����ٰ3�V`	*E���hH�����_�%� �M��D�F�M�������aS�<01Q۬vy:lA�s��nEI��[c�T�rmp�=\\lң�n��붆4���wOـI8^�.����evT��?�S�G/8�߯�_򘺞$'��O�q�i<a��������T-�b��'vffh��o��P��;uf n���.8�Ȣ�S@��MϾ��1n���E���$��y%������F�6/j�j�XyM��?�W�MZj��`�k�d���&�����ݛ����K�0K:��q�����S�;����s�m��ۡ{N��!l�V�wwI�����?O���2��߷W �홀w�iNRt��n��N�8_} ����=�0	�ÀO}�P�*鶓��&�	{"�=�2�?HQN;0�e~����WY�M�~�B����VGl�9��~� Z�������ݛɓC"�$b�5c�O0	�r�_} ����=���ؗ�~��ӃdfQ��Zm%n�&l�<��׉��ek��t h�s�ǌr�	θ�w"�[W ����@��4w߹��m`f�X<����]]� -J����mf �+k#�)�6��R5]���;M���3 �'+��K׳��d|6^���K��6��6�`�����������A�K��ĔĄ �
q�h ���\g$1B1����g�߿u�]��Rlt��Jҧi�/������1{V`U"��v�yD
'���p֞ ��M�5]%�Gi�s��b�ֹv7=�O���:*t6�b�]�k���πd���&���E�;������WN�j۫�f �R,����7۵`cy4���
_:j�v�`c� ����u��٘�#)�Uo�J�L��x�}�6 �*�3��0��`f���$�5�Ws�R�9��]�U���7W3���*�������Y��@"*��PEU������"
����w""��$*�)�X���*�	 (���j{���p���_��?����ο���_�{�������������u����W���o�?��~��O-�n���������-����������?�AW��������֏��l�6�;������ӳ��?���:������?����_����O=7��,����,/����G��K��;���C
$����B
B(�
$�*$*$��@(��H�
,��H,(������0�B*$0
Hʉ
$$(�2�B��H����J
@2�J2�@��JB�
0�B����J��)
$
$��� �
$�J�(��H�)"��@�B2���3!( @�J���J�
$(R��)�
@@!
�2�H�@�J$)D
̄����J0�J,�"4�J)*$ ��H��B�
"������"�
��@��)! JB�*�� J#�!
̄(+���A2���
�
J�ʉ
(�� ��J�*(�0�J�J�)*$�(�0�@2�J���������
@2�H�������
$�(�J$��@)((ʉ"�)" ʉ**�HB0�����*@@�!!
�H� �H�!(,��,��! HB�K+			!,��D�!HL�BA!),! � HB� , ��!
�(�H���HB���@B� ����! )"
!
,$�0�H�!�J�2���#!)!	,!	!!# B2$� @	�� ��� B
HJ)! ���$� @�I!! I!��)!!��22�(�@�*,� 		 �@H�����*(HJ��0�BD2��,H���J���" D!H��A(��� d�B��"4�B@��)ʉ "J���(�
$ʉ,�@)#
%
$2�L��J�2"L�*$J�$������o��"�������Ƴ�c��K���?���W���3�������^�?�����[���ʂ*���O���������k�Ă"��5AW��q��w��EU���<�zA��ί�r+����u|�OW�Σ�k[����gڹ��PEU�������O��PEU���������g��q��G��# DU_����PEU���������Ɇ���_�C�s����M�G���z�ڿ��V���s1���������4?ӣ��_ǜ����c�%AW�O������U\/���[�����7������)���V9����8( ���0���%@BA��¨*��$@T))@$RI�HBB�  
�Q) �!���JT��D��(�Q 
ET @Q  ��� !B��(*���A
HR�}�B�@�x          V ������<�%�ˤ�z :Y���C����܀�|�4p	�ׯ�s\yQCq�g�y[˅�F���2�"�pqz�z<�^�N����09v�#N{y��Gޠ 
  P 4<��x���`t
q h��  =,S��\g@���(
bh�4�:h�D�1 tӍ�4�JJ�Ҏv ��Nzk0JY�Ҕ�ҊR�4ѝ��7 �M)s�����QJ3e)E�iҎJ)y�  
 
 ���@GJ[�}�z�ɥ���=*����쫍�69�����L����}@�}�NvJ��@���o\�����w���`�6�/� _o����.m8�����꫾��R/|    � � ��/����˾���v��t s�f��uC��@��Ĭ ��w�2}9\�sʀwY������3>�39�����r�Ǫ�����5\��}�R吾�@�� P    v� >|���i8î9��x�����MR��6�6���e;������Ϟ0���T@��}�/3�}�n�z;�>�.aݗ9�{��zk� O�m�}�EŇ�s4��     ��)�R�  �)�����  "x�T�S��i���R��IP  "���Jm���A�F��R�" <S�N��?��?���n�jN���;��_슪*�.�������AT�tUQW�Ȫ���
���TO���)���ů��&��@�q%� j��\DbPX�g���bŝ�
	a1hD}-��۪5����9��?�s%D��f	�ʜx�"�5R)^B�u�x��HB�F抴@HV�`&�^��s���e��rLi,l������H���2��|Z�{�84�8iʻ�/6s��������|}P������w_W�H	�;�׽���ϣ�O�����u�Nvs��;�M�����5��qD��Czܩ���I3�>|�����\�ċ/�r��C�XɌF�Y�2SV�F���΀����[S��o���\=ᣘ!�����<�6�,�'_�;9��a�Gf�Cؒ�)�]���Mg�e�/�5v�#� 0�a��5��!.8���j�9�`��a݈�!��1Mn�r<LB7':����x�k���=�g;�u�98精�oR����<��`���-O��9��'�I�ѐ�n�02w?!��Z�wM\���v�B���<���� ���P3��OЧ"��������ظoP��U��{`��K{�ޜC��s~uNj������N��^Ҡqw��������ק�&�?��䖟uh�@�����J4ì,H�`
�ph�
i�L%p���-�aM��Okh��!�%P�j-u�$�*�aBq`�+k6�E-�7ؚ�v�ciz�5�kB=9�>^b�&�q�,om��̦=5��Iq��u�]�1n�ꆒD���i5�H�h`)
����˟F�*J¤���o#',C�]�$s[�贶F���|��*ϳ��lOn�fG��X�$�p�n�L8�]4焰Go��0�_���K�q�4J�CB��H�����(n#G,BX���W܉X$r$$��.��t2F$c^<pgg&;�&�#_����;h�p#���m�� �!L��/�'�ŉ>��b��x��#n�~vp�m6`�5BR!@�
��ӣd̈́�6Ҕ���e�֡	�oc�b�#B!SZf�#D�I�H�dR��h�**���N����9���գ�q�,�ƻ�g�&��]��Q�/���0�g3�M_�IC)�t}'�1@��	���HA�6
����B�����J�i�`�(�B��"�B%q4&���t��C���#�����,�'x"�tYH�_�d�4���^)\H��ĠA�Ĩ@�S*T�4���Nbs4]��"�ť�t�bc)�)�d$0ٯ���RVvB��HP"HH�#n�/�~'Z%�'!����V VHF	Cr=�˻bid\̩b$ w\���7fhԤ
D�A�
$i���0��M�j`h�L `A���
��M+�i��LX�f��������*5����.Bg@C!H����0b�L�h��܌�ňC!t�M�stHN޾w���,X�e��CŘ�.N�x�{�oW�|�o�F�M��w�N����x�zm�>���g��',����H��~�;��H{z��}�������.biY��<N�\Ė����or���=���=����|������IA8�+�q|�hu�l �( X�Ee5�
��^��0��S�1"`T��J`J���@���C���+����+����L@�6k��{�{&!��!G��8I)��ց""�+���HC! �2,�H�6����%[$jU�1�B1��;�i�$�o}ë~׸��>>���{���8��!���A�9��f��.�n����$�`��7�vo���䝧R���oA�y��qU�7��y�x�'q2bAD�d�Ǐb�o|1	���O."�6���T�DD=�<,��P,d(�,��
1��
\��Ēe�c�M<	�K�=,#5N0�$�6U�@�Q�(�i
a,���e�3�7�HҤ%	X�^f�-9�c�!CfT��o��!0���48�07���:pB&<@0`�d������F!B5)���M�ne$�$f��4�i"�ql
�4�L<���>E�W"dx�5���>��z_�q����KU�O�c�=ހ����P�BP04�ā��@<�B�!�K���n���n'�����9Hs2RS���
0�B.0�5�(��~����G
�!b��@��8@L���+�6���V.�'w��Z3�
����]�/5�q�)X��W��-X�!(x����ԗ3��!	�fyv>o%}�y�sV\c1���=5!v�p�#��,<�8q��I���r�s9ý4If,���o)p��=�bZܳ�'{�r5?}�!K�d)%xY&�� �A�p�g@�H@�
a�o2��s�!I��x�m^���K\9ƪ�O8��F��x��.̂=8=T�]]j�9��K�}β�^i���sy�b�VR���ܸ�,�
K��m�Q�y�=zc��{�ǂU����.!q2b�Q�G�X�<��.]3Q��\HϾ�l��(A�|[T�N�:|B��;9��Юl>����Nv*5���TL�Nw���Z��>����#?!�FN
���&B����Y��\!\�H��@�$��$T�sv=�פ?{е߽g��\�87tgVl�O������*�ޜw�8abB:7��NȬ������u�ֻ�oƽ��.�G�������Y�,,��3�D!	 B�E��`	�� R�"�61) a8Mܘ`:YCp*�!���;ܙ��=I�E�Db�j�M����P���қ�a�� d)�;�X�M�X�ѾCm:{:}�1'�ףּ}��c�&ܧ�s�����w���H0M�mӇ�d.��Ϗ�~�f~�D��aFJ��	!F��R�~����+�0"4� W�����H�F�2�w�w�;o7Y������*�G������GzNr�w��=�ˏ��OP�7��\�!�����K.���CCp�������@�
B��]�DYp�np;��)�:\�`�c������9M�s֑��-.���G�ԓ"�����,o�"�8��~���;���C-��ňrHSr�$��IG\8�r��o񣞽�~����s���x�x����Wj��Ѱb��&���}����S4��#�6�!L�y����c2���Ҟ7)�
e�c !��dR�+[��x�3#��)�æ��d������}^GP�C�$|�=}�M;�^K�iK�<���u���O���{�缧��G���Ky� ����^���W!܈ ��5ww�z�oS1izb���h�+����p��	�g~�@�t�w����7�u���,T������W��x_w��48;zn�sd��w�b�Ǐ{؆@����$�w�\������}����q`�=�SE��=��"c��f��������],-�[�2���ݝmzM�m�:����M~�m+6���P	m��;�_W������6)�K��7����z,r�;ˊ��\�^�n�o�������t��%�9�J��;���Q���3Rz"C";mc����vip�b�'����;�ηƲI�6
Jy4�M��˼\�����>z��nU��a\�4��)�M,�$a���2�٥F,(K��X��3Z(����	
�x��p�j�<r��3�Y�I�I�t�E,�.m�i�lJh�H��$�b�̴�M<?�&�Ouĵfg4i�~X�	�0��@��]����%��
d��A2^��ŏ��C�]@��(�BK|W�l���l�^�����6����⑪Ɫ`|b��R�d�Q�#BI5`�tA��j$��(�6����R���nj�Mך��>�˼���w��C)��^�����Qn�Nu��{<{�ŋs.����y��9w���/s��Ř��)�<�
]�W:�J=]���o�'y���a��^�y�R��n��U�:���%�f��f�Ѭ��L��W�:&�r�ao�#�K���$L�@Ř�!�.�W��l�v^r�҇,�����BI
�\BȝIS�,p��$!�X���2�y'gyD�,�d�d��e��ßf��I#���"��+��! "��E�4����w��{���66����1�V�$X.�d �`�@ �hVH�"F36Jht@�]���=��F!72���:t�(!��玱	�����ɔޤ��5�gc����^~���&B�����v���L�g;P��:s�pf��y�q��n'۲On���;���sh�:A��7�5�>���L�
4�[װ�����eź��k��7{_y�jIX#��6n�	1xGU>��_��S)
��(K���\����o'�9DFo7�֙�s�^}�x�i���b��	VhІ�C CX�����O�u!BS|atl�]�1�LX�$
& ��!�b@h�K����R�`��<��@E�	�LF30�!Z���]�����4��}�[<COk�y�{��rH��]��GI�.�q�^�۔r曁p�@����b)�.�R�m��  � 6��m��              ��H�n�^mmźg��!��Mh��W �]HW[��ei��\�Zl[C�K�o-��k��*�R��X��X݋� ��lM-�EY�l����Wi�B��-���@�F;2��㖭�����.�`�`X�PV�*�Y*� �Gr*j���	Yw���w8�m��A:x8�]WUT��	[**�]m��\@Um*�ʵ
�i)K 	l�]������X	vK,��0 d&��fI�%�H�H�8���i�8ڴ�v�!�Q�����w-a#�۰v���O%6ީ�k`8{q��x|�[f�صnpv��g�!���t�$ڐ�FK>�W���6��Uu�A\�Z����*�_W=�?+��yBM�Ӭ6�[�m� @�� ְ[] I�Ҳf���ר6�7Q�md�S��B@m�.�h���Y(�\*�uJ��p�5�:%�R��l�f�V���b^⹪j�nU�j���syY�ȁUoou	3;2� �9�s�.DQ&�%��]xX^�4��lJ�Z�S�����S)յl�Λd �a�ܒv���K` ݥtp�]U^50&�Fn2vNbp�"Αb
���n��کV���,�!0�Z���=�V��-0q��:}���}��p]5�nu��j@]ZH{i ����v�h�o7/�/���ܩep,�p ���m�[�]�����n7�r5݀��,�u
����������)�� %�ٰ���g4�t�i7l�v��� �` p-����.�:l	 u�gH/��������� [��/^��m  -��Cb�t�1�Z��ր� 'qc�m[a�-� 8�m��H8c�46�uUm@u*5�Un�@ m��M��I5��f�� BM�bl��HF��km�i .�8Gv&��H[5u/���7m��my�nm�W%e�G$ mr��.e�JM}||�ʮ��U*�&ЛKj� �����Ҏln� �ڐ�n�kЖ�[%� 8��I�v��&�l�\��q�:�T�^�L��j{E�u.�k�r	ͮ�U�M�81�nm���[x  �^�:�3l�m��� �-�HM���<�.� �Z��5� �AR��7^�6�ojQ%����I�m� �l� /Z [Nm�:$������֥��[��
�D���*�p ��H�m�U���d`���J�^��H4��6$�@q���Ö�� ٶm����çezm@5@J������6����5��J��U=vⶺQL�p�Kq�v�l]���lf�ɲ�O��OK��4�P@�0���l�T����kkcU���]��o����l�\�AR�V��Ϭ�[sWS����Ah����t���.;�� �;;��-UR����e�y��n�}�  	&�&ٸ�v�I����-�� Å�<�X�b���$�9 -u�H �bYP*�Nv���� d�$ M��Νam/�uk@�Hܷ�`�:�m&�	�
�U�����UR0����\-�$K�sk�-�E��U@r�+��8� �i0ZkmdhM톪U�Vڀ����6)I�$��[u� �>  8���` [@��Gn�K��YR�"bM,�m��   ���3$��M�Hת�Z	�ܙ6̲�� �7Z΃v6��aSh7ew���e�k��6T��\u*�m��Ӽ�ʬ���6�OO��]ʚ�%An\Wb�9�7z��2WO+V˘��X��m�-����G4ܱ��NC�s�L�g�nw�ȃҡ����P� �iح�u���Ȼl�0i�8CnC�Bj�U�n��U,\�J��Z"R�5 ��)`uN�T��= ��/K ��pp���������}��n��l���H2!"l�����  [׀6�-�t4Pii�N,2�n-�,�Lb�t����   H�re�I��Tp�@��T�������ms�m�m �G:Ŷ��:����l�`�im H2��%��j�cj����UU�f�ef��J��tt�Kh�-�� �6l���n���-�h H8	-�8H-7e���.�v� 6�D�-�m�� �t�$ � m�h ^��I Hl��2rtm��!:Ԙ�`[@-�v��(A��p ���m&�[ 8 �����kXN� �Xa"�6�m� -���$�@m��_ZLW��l�6����ʹ� ��Żl	 �`m�@  H m�mmհ���h۶[�� M,�[��0��A���KJ��R��m ��ܶ�[�� 5�n��'ϧ�|h�$�$$��Y ���m�m�A��޻mt��m��7n�4ځ��f�$�M��l$ lH'N�sX��͖���@Tq�ʻU ڪꅷ&��$��а� l�!�ܐm� ��8�mt��kd` :Y�iXi  p	 �2���K�6ͳn<��5UP@�hC U�m�v����m=Ү1�m�6�1���r�Ҭ�e�j}T��l�q���N˵@$nYwH�۪M�Z���e��#��8�i,c��>r��۲J��i۶���@;�Tc���z�ýӶ��4�ɝ��O���c\�O@]0�7gM�!��痖Q�x۶j[A�PnG�[���O��3\�(lV��=h5�{:����]��V̪���[��;��r[>�:���kv��9�8-��l 9t�����9=��ݩ\��^\&�p��� ��p m��;  8�(��6�B�;��ZP�t²�U�m�n��bKk� H��G���>Kd�'&�%�zYH�6Y\�պ�S� �v��˦ͭ��j�J��+�*�T [@ �׭�m��U�],�;�.j����`{U��wL�d�����e�|}�����,uK�٫[w���i�
��ɶ� �vf�$�t�u]����ِ�s%��v�����^��Szt��T�nRU�&��)����@���Vx�jj�v-���/Z[Rm���T�P�s��Ch6����yn�v��d�W��3��s郥|�cR���3^���T8���ձup# 9Ň�k�%��M�)lǯm�oe�ذ�ĉgY�.�N Y�eZ��\z]u�Zax�צ���[NRCv��{Y�n��qζy�m�v�u��+lR�k��J���8�\+UU]]�D�h�Kڋ!K�A8-��<Um@W;` 6�m��5��5�Uà�� � M�ݙ�B[y}�hm�	�V4�=$sm&��� ��ػ��l�I��l�h�6ۓ�m ��"-�lӛP�(8�M��u�-�[A��pմ�  浭�@5�e� x|>�Y��i���vV���Z����`2qK�ܓ��Y.H*	e�	��j͛khs+*����YV�Yy��rf�ʱ���j�m� �m     %�	 h � ���ݨ
���u��� lO��}{L�R��ƻ%� 	h 6�� k�v;T�g*^�j�s6�H -��ztv����@Y�e��W�W]�n�q�o�Z�%m ��ԫ�]�=r��L�!;�8�!�j��2��9Xs�l��e���nH /t��8����6�e�����b�ƞoE<ݏ���휈m�9�X�1s��� xD,ѩ�j6�8�7+Q�D�� 6U�=��i���,��2�WZ��̹Zp�7k����� M)�ܵU��=J��s؊���5Q�e�c�mtq"@�zn
�,��p	/o�ka����ܕiN0�4�K��nu�\tie��P�\��R���cXv:�!�F�V��\�5Plt�ge�;e�Q4�*�ěl�(� ⬡��y���w`+���Mv;k�d#fZ��l  � lUT�����Kf��{Mm�V�#�93=\W
�'��9uI0=�ɝX�6��Wmt���vt��,�����\=��XzWͼ���nNw�7(h�,�R�	)���5[q����wmպ���f��^޲�K

C<�ɺ6l�$�"'uIc�C^�zKzZH+I!�HV��[GW+r�[�L��h�M����[@85TJ� �\���ڥ�bzm�{Z��fڐN  ;H��^�$�wY.�  �`�p-��i���敺Z��W�q�]A�:׶��:-� ��AoV��amm��mm��Im�W������(��$ ��mnl UR�UR�1s�2vܬ���n�6��  t��jE�T���+��l6�-����m��8kn�i@6�$�l:ޡ�뭈-[����H@��c�n��� C��^Z�]�땥V��N� �9��H  8m��t�׊�F�o� A��h8	  4�D��[@ t� �6��m� l��RB� 8  6�H lY�z�N�m��m����v 9���M�
��ڐ�4];jm����H�$��صIe���ONk0u]��ݜ�c흏٢�v�E�G9C{n[��5��j�kJFm��o9��G/WgK��p%�Z^�n�
/��x��N�m�[���e��9H�� ff`ff��^**4?���
늁W�"Aa	$���	���b�����Z��
��)�F��0j#�Ģ�
��v"^��h!�A����SWN�UH�"��8��<�$b��q@>� �WI�D(%��>#B D\D�b�i�����x����@�����$��+$d �i: ��H��~@��ʡ���Bd$ G��W�@
��?��#��|+`� , ��$: |σ`
pԑ�m+V4!����*	����}��T���Q4��?*�Ё��$b(�Q���D)�~4p�,�J �Qh"~�!��} O�@?"����~D�'���\6 �`�*��BH�H+^�iUx�L] i+Q]��O��pS�|�G�^��%Qz`�R/@?
Fʴ�?*t���)�N� ����5@H:�FHB@�$��$��N"8� � U8���H�:q҇�Tʉ���	@�D�J�X��8��U?,EBO¯Ew��+�A6�Ų�H��XU Ȭ�HU`F$!�!II$XO��"���5H��#V,�Pz`�ֈAE�b�d�� �����P{BHA�A��I!��PЉ7W�F��D�H�B"Q4�8�tUQW����<I�)i���!���X*��b�d���׽��~�ߏ��Ŵ  .�QN��oo]s �Q��2�kv6鳰��h1d���-g��֭�C���vg�Ԯ��7W)܎�C�x;R1�<�7�Q�7S{y�ە�7A�,ma�J���/XT��Nw!��M�U�Q�'I:�ݻJC�ۧ��TL��8�P<�$��x�:��u\��hH�^�*�[��nD��]�:v�h)��pt�vy�z1��Ա.�"���2힬X�r�v�\��Qi�RvI�˶�@���>�.��Bm�Ռ�J����\���{n��F�w6H�un:١��ݲ�]tb�^�fI����9ݸV��n�m�y�A�����d�C�tnU�s�z��M	x�9��շ<�䶹�*���gS��3�2���Mrr�D��I�����Q�v�c���.�0`WSw;7d�&�d��;XB�
�+p�A�ڳ��]lN�-��&�rQ̛d�h�mNs]�i)�ݑ�9ԫ^%Zm��Z^!�AޮKmJʫ+H<��S��t�κ�f�����(t��L��c�8MΆT��p��y�;��7܏8��n����1��[�ƺwOmM�1<,�e���$_60b�Wjw7J����Һ'�H��󎪐�`�y/b+�:ݓi������GE��ݍA�Џ���z��kk�\�X�ԇ0�1����Ͱ[՞gC&�V��9ԡӴp���X�e�<AG:S������z�L��Z��mV�DLn�#�jK��1�&�p�q��U�¦��0����M�4/�mU@I�Dl���.U����:5�6���\�dű�4��{g��
�����:rE�౮��h�\��r�fx�3(��� x��m��d����gI}1zrh�X��5�<]qq��9Α�,s���K��z"kRl�v�f6�k�e�[6�b�,KL���AQ4��c^�����g�;&�l�̩-�a[��2R�@Xr��n�:nU:���te�6��m�4�^�ݫ��1��f��jjL���CB?Ȏ���)������4~QC�Qئ�N
`�Q?B��~A8?���� �F�b�ݦ�.]��f1m��Ѯ�cH�]�3;Y^��`�m��y���퓟b^e�`�;�s�8��s����b��춱�r6�j�gk�q���ۗ8"�T�äPܬl����J��WA8qb�രn��8��L	�㍻���azb�kr�nm�vr٘1nY�l�ۅny��]�l͈��a�!9�D�x�"\@wFݥ����0P�y�YlyfB�.�0���ˎ9L��+��>�@�8�Wx�=m��ͫ�ʊ �ŕ� 3w��բ]���&H7�8���n���[V� �u��l�>��bI��1(�(���]��u��l�>�����cىcc	?�i�&���W����u���U���=��iI�L���iŠ���u��*�٠}��h�����~��p�������I����v,ny�g��i1�;�y9���(�����9>�nhZ��>���٠|�.j��6�473@��f�5���Cf�ma<�@�=w�f�/�@���h�|̲� �����٠������٠|���LK+�!�I4޳bG^�˗uXt̥��V-�Q
���L����=��hUl�u�@�{��陈��R�O�hr�7N�'J�L��L�{5�t'/i:(�P�Mf��&�<�	{$���CqF�2I&|��~�4�h]�@�u��=�fɂ���cM:��3]��3]��n�X��j�&"R=�����"��N�����������u��POԡ���RZ�`@�Q�s��]nI�����>�D�N��Ɂ�'��[��if���^��mz��sW$�$�)�`�� �f���^��mz�n�<w�����sˤ4u�t�T]ꒆ"^A�Vw1��B��n^�{u;���"�̚�uz������ �j����&%�B�8S�>[��f%#��q`�ʬ,�v/6��PL�L�D��>�w4�[4����ؗ+=�߿=�;�u�)Y2I&XlfՁ噮�Ź��b6I�H� �H�s���o�7$���ܛ։q���y$�<���9^�@�����Y�_teC��������gtrJ��\�s��ζ\z����m�yj7aOE�\����'����<�W�}��h^,阏�b��`{�Rm��P:
��:z�n�w�Y�y{��<�W��\۹q%1L��hz���^�3�.�v�z���f"�U.)T��J��âf!y��1v�>�mŀw�Y��,9�"���	#�<�W`}�ۋ �lmX/f��b>ʌ!j�ڴ���-mg]��1<��.cc�Z�te�7g��[�����8��wBH�u�ݢf�;���@dv�c��8�y��rU���۵��L��h�>*�ʻ�����x���v��\Eh1�<au�nŻr�lr���΍�k��=��М��Ӻu�Z��j�������vrYZ�;;�nB���}?|b����w{�������\N������w8��m�3���/�;k�>�y�a����9��P6�ո�]XtP��m��_ۚ޹f���W�y^�@����X�IH�ɒ93@;�,�?�<��z/���>�]��9\{&#<�)2M��@�^����hz��am�4���Un��L�D,}��u����h/uz֨�i� 8�N=�u����4������&"}�T(K��$�H�v���{N�Ir+�Y��4$�c�v����)+b�ē�!������h/uz�澈����z����E�]
��*���krN_�w7�����DVf�I��B��Q������I@ԙ�(��_ʸb���|���ŀflm_LĤ��@���S�����{6��366����ԗS�֡�R���lԿ��@-������W�y[^��Wؓ��	H�ɒ93@:����@��u��/r��D�ȰDx�d�Wk����yV��(�nm83�8z1v�F�W�C̓����8I�|���Vנ}֖h��vcJL2d��Ǡy[^���S@:���>�@��cwa1�{�4�,ٳ	�P��:��S�����w$�zנ�ͻ�GQ�Hh�+�>��+k�>�Jhgr!T�p�ɄP��hy�Z���{�4�,�=�bˏ<qɑ�܉�sPv(x��73�۵��M��KgGRh�M�g�N�0�?�Y�'��mz��M �}V��<]d1L�L�E#�>�V���n�uXǼ�y��G=��2��:B��������V����@��)�w�Wɂ��x��
HM�>�@���@��)���1f<��C3٘<3/���5%�|?���[���n��=�`tL��6��]�����S@���@��X�2A�&�/S����V�����ci<�b�����&�M��f$�b?�qh{�4+�z��M ����\۹$q�!����z��}���l�>�JhgrT�p��E	S@��)�z٠}��^�h����b��,�y��}�f���S@=z��}��=独�&)�	�8ܚ��M�������u�$���[�q萀0!�! "	#Fԕm�����s��A��)��	�����l~߾��>��z���yrd,�':C+I�N�H����M��T`�Kх�\u��eE�H���',d��\�fV'O8��=�Wgҁ�I���wlU��F����s���-�lJ��s3���w�u����n2�X�=e	�]���SɢG=e�\״�⭹q�U8�[ �/U��fix�e7�q�:ˆ�f�/�H+Ew�f�)9��5�q�|�����,z�usv��>I�KoQ����ѱ��,v�t���m�m�����M�t��}�f���S@��7���x��
HM�t��}�f���S@=�4z�1���ɓۆ�}�f���S@=�4�Қ�Q�۸@�2b0�@��)��\��}E�$�޶}�I�6�$Q�!��jI%�u���%�r�RI/�l����ZԒ^�\+�f!�QD��u��BpF�V���M����]n���WO7)7%V"��R��K�z�m�}y����ֿ�136�Y��}�I�A���
�O[m�w�9�h1��lĵZ@,�b(�0@e��_�ߣ��o�����K�z�Kޘ��dDɑB)��KϥkRI/z�}�I{��Ԓ_;���I{+����&'�d�Ƶ$��ZO�I/s�Z�K�z��I%�-I%��7�Ĳ4Be���m��ߛ��~3���m�+iZI%������O��!G:L��>�"FNm5j�s ����dc���:�s�K64p�%�X.��� �������^�bԒK�rϾI/t�-I%��[m��	�&#�N?�I%�-I%��_�$���R��7�����n�m�TyQ�RE�$��O��K�%KS�g�:6�Y�0ϑ����m��sw��}�bk�.��f&��H7��<3�����pNt[ð�D���2���fZCXY��9��Mu^�ί�#$�8@���g8F	;��C>(na`���;��}����}�SXئLf��s0fa��&�w0��r�.
�駎��*@$X]}��_~���$Y A������&&C4R�캚B��!�T���E����)�� X�f$%�Jf��1�xrVRBW���~I��`0X�B�� �23�Ǽ�����Z�NO������)���:`����J�)�Nwz&bK7Am��K���|���µ&7:xGo|��Jhs�n��]�kL��8t3��{�`�'�c�dp��o���ǶsD�cx���`��1FJ���Є�SR[���&q7�\���bi�=�/&f3=�4)��> ?u6:�8�b'���� 	��z�>U� ��E~�D�#�Z(`�A�I�ֳ~�s�ڻ����^���s��3$�FI��%�ԭ$��濾I%쭥i/��]W~��}�I.8T~P�1%HqMЬI/=�|�]6���!-�:��$���+I#�����?#�jGJ^��ы]�C=[��6tm�<��'���=s[s~���gF��N'�I#��MI$��g�$���/��DG�󤖿����Il~u	�̧	��ꕤ�Y�m}�D�6�mW%i$���6������$�������L��F���$�]p�$��濾]3�6��I%_�~|�]�ٍL�S&<n
�]33�v���3k�������%���� ���VY-P�� ��X��Lh�D�Us~���ZI-��+mtH�:|�K�]�ݶ޿ȉ� �s��ﭷ��K�m��s�I.��k��a��"rD��Mų��}�
��cd7:����Fֱ�@rۛ�=�w�Į�F�D�,�|�I_�?O�I/s�V�K�s_DG��K6����Y��u.�dU	UU2��$��֊�%��>�|�K6����Y�m}���1UH�EA�8Ll�T+I%��~|�K�[J��ڿ��}�Iu��Z�K煶�� �����K�;�i$���_|�^ʭJ�]�Wo?�I,�P��)�MU!P:n�ZI,{���I/�11�{�%�Z�w��ɶ���z�m�F!!�I%���7M�	5e�E�v�oLM;)�t�'�Y:��*��w!��{��]��*�u���^'+ƴ��y�7 ���t��C��+Ϟ��X�ٞyxj���u�d�6�8*�b�S�ݛYl7ݳ\�r�l	�u�-��y�9��!�]���ΰW&��jX���*��s��ַ/�2j�We���M�R���s��z�]	�b�BiJ����;�	,�w�籤�,��4Y�k��o�����l77y3E���;������.~��N�P����$���%i$��5��I/em.���IW����$���n�jdȒ�1��q+I%繯�fif�R��Z�N|�^ʭJ�&i{�+mpR**�'O�If�R��X�|��?�&b����%i$��~�?�I#�Fݒ81DL��I��&f[��9����ު��������_�";�i$�n�|�j�dU	UU2��$���R��_�f?D�����IoW�V�K�⿾I/ftB�dE�f22<g�Ў���v�6,��)�W�v�l�X4ݫ�%��w6X(�![�ʪ��I%����$��VҴ�X����Fe$���%i$�j��TJ��:���9��}����\�������j�f�~�r�~���wm���{���&�����s?�.MZ)�P:n�ZI.�����%畭ZN:f&j�_w?�I%�]J�I{�-��T
)���s��(����eݶ����-�{+iZK�f!��]��Kw�]�5U	TT8n���X�u��ItL���_$�����$��kv�K�L�O��$�C�O�gS���MW:�g/u��e2�e���;�Ƞ@�����'�N��]\oa���$��~�i$�in��I/7��LL��K_w?�I,ZRo����H�!�j�In��}����7i$��s����֯������3��U��QO���_��km�O��s��� 2	"Na�CQ
����J�b�2aKBUV�-��L0W��̬�}Xդ��R�|�F
(�)���7i.��ok���$�=�j�In��|�艈yU�ݤ�ݨ;�����:|�^yZդ�鉞�]��I,oy�I%�w_�$�鉈�p���BqRyc���"V-�N���A��s'f�j�gk������w��r�X�[R�� ��_�?�I/7�ݤ�ǻ��fc�i,{\֤��*���0Y���q��Iy�����5T�?߿?�I-}_���[��_9� 2H���Wid�T�,IF�[Ic����%畭Z]31�����K�n�If�	��b��U�U?�ItL̼��j�IwW>|�^o5;�>�$
U�)d��HU�� ,��f"�&jc�fbw|��)7�T�b�U�U;u��`t�Dy���]����]��&f=.6�.A�ʴ�n`]�j�����C��N���bK<�����w���7�9�QI~���z��h/f����s����4���BcuN�����&fL��f-����������k������uP�QP��N������z���"f?DDD7��~v�?��h�cl�x�H��H�z�"Wus�`f=�`{^��3�&"V��=���c�0Y���q����11�b7����-����^��f'0K�0'�|����X�nJ�w>�u��웶��\;�n�x^A��n��靷�C�N�n���\q'f	�5v���:��0#�X�<����;��Xbɐv5;�\�ó�=`��/��;�]nڷX�Z�籖��1aau��n.kpk;N�(�Ckj�o���t��ܓ�x9ݔ��1��#�$�k�����}��mH�lQљ�p��<p�0���f �y�J;GG"J��:9%}��[s��;ζ\uی�7m��g¯��{�n&�jD����Ɯ^����@�zנn�z�"b~A������P��LiЉJ�X/n�舘H�|����X׺��"bR3���U7�ATBT��ϝ����gLLD%�����w��]��ϕ�jE��]�Y���33��2+/�����Ͽ+f�����]�ϝ��h*�%��ƪ���{��鉘�[���ϟ;廮��u*b֩<[�٧x-����]s�^v���Vn�+%<�KL�}��{��՞��1h�����V�׮��n�陙��g>�`~�f&��<y!PnM�]z��d)�V�!$��Un �P0��P2�DKt 
�"��p �ɫ�~��?{=�$�ﻫ陈�H�5t;��"���m�N����`{^곦f%#wz�滝���V�SeE	TS��v1���X��X�����������r�	�:*��B%*�`��`t�LDwV��������`f���#l(�0���Y��:�ނ(�ʹ��v�2M�]���n���총�7Ҥ:�������s��˻���y���LD���ޫ ��O��TUI�UN��,�w�"#��D6g�ߕ�ow�7^m;蘈H�49��L�Z�P���缬ٛV~��LD�|Q�fC"�(%L"!1�$AH���G�g���z����{��&)�
B8�:"f=�vsާ`|�u�t�J�U����i����dIdɑ��_X�������]��,�v�!S��b��8�b�lpƗd�-��Eγ���/hbN{�����?Wlu���n���yos�>[��,�}? �{��΅]Pӊ�2�:�`|�5���1٫��?/�����f뾉�H��6�~���?���9[��^�i�&f?LL7��~v/�����ڦ☨JT�:bbW>ު�<���-��ɱN�lH�I�����e�8C
�Z��f䓾�s��J��Ymԗ��jK�03?����?���5n=�=�k\UBC���#E�����l�/���ݨa3Cv��cqgN�󌶟�̱T���GF;l�KϷ��{3j�ո��&f>A����p~�j�(�U�嚒]����� �E�~��V.���-�w�""e#�j|��2��7U`r�}V�7]�	b��`��`{�-�uP
*Z�i�UX~�������`b�ߝ�{3j��L�舙���~��;B��:
2�:�`|�5��b"?D�D���^�����R\~��#����ng�L��ςU�o>K"~\��(�ϐEO@�b�~'m����y����D.�MgX�1%� FBk�k�;aN�tü9���e:k�<����ٴ�}�����ۘLJb.ܸC[�$�cm��ʏN����%���ج9w��� '��B�)���X�6̌c�6R���޻�:�y��G�6���Lz1BJJFBHZ������H�20��YI-�i.`o�!62FB�"��u��\�Zj�sZ��nm� ��I9�N/�����2Qp,����u���$H����,�[��;�%�;�qлj̊۲g��͸6�5��S���jûp�l����Ӏz��d������U�y}.��kL�םU���6į7q�ny�kt{>Ѹ��x�.ͺW��W[R�cv�F�uuv[���[UF"���^������bs���tql:�v��-����D����<p�|� e�\K�G��s�Ů_������A֑�Tr�My�v�"V��ĢPi@ɽ��,���H��;s��;e
9�i����/Kuu�$d�[<J���Ԋ!�v�F�m$��:=�q�X�n�6�m�u&-�q�G%m�+]���UTW��l�g�{:�^w/R(i]��6غ�y����N\̃��Zɗc�R�(Ӎ��n��H:��of��/'���=v�ﯴ�!�״u���� q��z���5tO��G&��C����˴�J��qgb�l���\�����]�f��5=��t�GWSp	�R�v�jq�K�̈́C�|�֥Ikb�M�[>V���yi�8���^�*�������:#G&�l��s�^�ۮ���.����;��V@�`T��EpM-T��O;k��;.��9j�\��9�n��s�٥�jQ�g��.�;$��=�m���[��l��l+�y6�k���T����Ȭ5]�ˇn�g��l�q�۲Uɶ{�J9�bV��ٷk%&�6�6�ݵr��F�l�l8s���+��2À55P��e%��"���R�1:�<��\�]�����6���%&#���UFq���<��R�V�ӊ���:� y.Ks�1����3���NբU��W&vY�2�ynh6SF��H��Y����њE9ж�{�(]�9���k�V�'nWN1ɺ��'V�ܑ�ӾHF�k���t\0c9θ��8�<�ۓd�Y����R�z%�HR+��.�z�H�X�h�M`̆0�)��:�y=�nz���5��jҠ�N�x|���	�/����O�/�?*>E���N�-C��� >P�^��D�;-��.���u5mlDZ.�M��hQW���ؖE���8m��&v���\䊗���1�s��7Y��&G4��y���b�ڤ�L�ѭ���z7l(&N�祶�c$��S���M��6�w@��Y�����=g�MvӺ�u�zb�:�S�wg8��[
˳��˕u�{Yݞ��n�7.in{��;s�����Cu��f�Eŵ��33Yf��pS�*���n[)�j�g����n���
v�4���kv���K�z{>��z>�{��>yq��Ȱoa����߿U��u�X,�}�]��h�ުn)���B�UU�����D���l�߿;W�ߝ�{3j�fe ��O��UM'N�*�t�-�v��:"b3w���˺�a���B`�B�UNæfV�w+ �ޫV�ڰ阅��@��H,��LJ28���h�"g�.��-�vk�V`�mA�J�ؗ��]C�=r=e�bܽ5�9�q!�v��K;M���������iv.�[��c�.�:c�{��|L"a�ޮ�q�P�?�dKĽ�����Kı;���g5�Ji�I�.\ֶ��bX�'�｛NC�XP�-$�!D���Ldu�0H�B(F#"��E6�"r%����fӑ,KĽ���ӑ,K��<���>"bQ0��Lnr/�):
2�L��fӑ,K��w�ͧ"X�%�~�}��"X#bX�g����"X�"&<������&0���V�E&�հ�3Y��K�[���[ND�,K������Kı?g}��r%�`)r'�����ND�,K�M[��l+nP�v�Ë�k����~���bX����m9ı,Og}��r%�bX�����r%�bX�>�o��wf�,�gt�[��3m�ֹ��9���ngv���m�K�q�{������4��uu��fӑ,K�����iȖ%�b{;�fӑ,KĿw����X
~��,K�ڿ�ٴ�Kı=���rd.I!�E.���r%�bX���ٴ�lKĿw��ӑ,K��ھ�m9ı,O��{6���bX�'{�}���:Q��+�nX5�X5���{[ND�,K�j�ٴ�K��)t("dO����ND�,K���6��bX�'���g��d�F���V�[ND�,�D"	�;�����ND�,K����m9ı,Og}��r%�`D  ���{�&�8}���&�&��ĩ$r�0H�,9ﻤ�A���6��bX�'�ﹴ�Kı>����ND�,K��?q������qn�a�ͦk�9Ͳ�4i�ۑ������]�g�����������m�Y5�L�ֳiȖ%�b{;�fӑ,K��{�m9ı,O���f��Kı?g���r%�bX�{�xfB�SWW3V���fӑ,K��{�m9Bı,O���fӑ,K�����iȖ%�b{;�fӑ�,K��V��i���2]k[ND�,K�j�ٴ�Kı?g���r%��b{>��iȖ%�bw��6��bX�%ﻒ~v"ҩ-�;\�p���� � �O�����ND�,K�;���ND�,K�ﹴ�K����E ���!"�]*E� ���������bX�'����C%�$3Y)sZͧ"X�%����ͧ"X�%��$3������X�%������ӑ,K�����iȖ%�b{ڷ�d���oDPuZ^��q�{Uxs�;��5<q��G\�3�ěs�>��Ѻ}�/:�֢��Kı/{�kiȖ%�b}������bX�'����P9ı,O<�w1�0��L"c�m�Ȧ�TRJ��3Z�r%�bX�g�}��"�bX����m9ı,Og��m9ı,K����r(X�%�ߧ���K���MY�.���"X�%��=�fӑ,K��}�fӑ,�,K����r%�bX�g�}��"X�%�߽f��W5&��.�I�Z�m9İ��}�fӑ,KĽ�}��"X�%��z���r%�b���=�fӑ,K������5us5l-��m9ı,K����r%�bX"��������Kı>�����r%�bX�Ͻ��r%�bX�Ml����T)@k)>�wmߧ��I��'F�q@�x7MmӦ:��B��=��w*ZN���m�%d������� Okms�7t���>A5�Zu:�<�M�����R��M��2�G.��x���/f!G\d�pn��pcuZ5kk<g\`��kk�uƛ�����7a�_]N�S�	gt�r[�[�X�J��>�n$MK�a�pB��r[�c.�����FFЭkbiX�W%����ᙁ��2���@#�j�u�Թ+=7=�G�N��2q�F�����2���6���GI�%ֵ��Kı?g����ӑ,K�����iȖ%�b{>��a�"�&D�,K����r%�bX����z�%T��l�W-�8�k�k��~��X�%����ͧ"X�%�{�}��"X�%��z���r %�bw�Og�10)Pۄ�;���D�&1�;��Ȗ%�b^��kiȖ
%��z���r%�bX����m9ı,N������(�U��7,��0�������bX�'���kiȖ%�b~�{ٴ�K�F��}�fӑ,K��i�t�QBT
������L"aD�ڽ�m9ı,?������ͧ�%�bg��iȖ%�b^�����a�Dƾ:�T�	*I*�E49 �Ga�����ZzF�cQ�Ɏy��n{]�>��@�{�޾�s�v,��`Fg�w�����og���m9ı,Og��m9ı,K���ڨ�%�bX�{]�fӑ,K0k����KeV[$J;l�8�k��}�fӐ���2	�CHEM
���Ľ�}��"X�%���{=�ND�,K�{�ͧ"�@C"dK���3%��k%֬!nf�iȖ%�b_{���r%�bX�{]�fӑ,D[�����iȖ%�b~����8�k�kx����
��t0�Z�ӑ,K>抎�g���ٴ�Kı>�����r%�bX��w��r%�`+b^���ӑ,K��{��]EU*v�#�K7,��ó���p�Kı/�ﵴ�Kı/{�kiȖ%�b}�w=�ND�,K�ue�߆���훎�:^.�utlu�mw3t�Sb:ح�j�U��̟w��}�~�Gh�f�iȖ%�b_}�kiȖ%�b^���ӑ,K����{6*�bX�'g�ߦ�ŃX5�X{����5J6Z�.���"X�%�{��[NC�"�"X��׳�6��bX�'�����ND�,K���[NAı,O{����Y�����[�q`�`��~���Ȗ%�b~�{ٴ�K "� 0bA*�ԂF`)��� @8�L�}��[ND�,K��}��"X�%�ߧ���K���5-˚�fӑ,KB�����iȖ%�b_}�kiȖ%�b^���ӑ,KV����{6��bX�'~����k(겻7m��`�`�{��p�KıE/{�kiȖ%�b}�w=�ND�,K�{�ͧ"X�%���������3�v�u��a�u�Y,9x��Eqns�m�a��L��:�yS���is5�'�%�b_{���r%�bX�{]�fӑ,K����h�Ȗ%�����w,��þ+~�B�).�	u�m9ı,O���i�%�b~Ͻ��r%�bX��w��r%�bX���m9�P" dL�by��?O�ֺ�UK,���oq�����w��6��bX�%������b�X�%���[ND�,K�k���r%�bX���=��\��-��\�m9İ@,K��m9ı,K������bX�'��sٴ�K����
b�b~Ͻ��r%�bX���۞Գ�Ce-n۸q`�`�����8�k����{6��bX�'��}�ND�,K���[ND�,K����.��>�A7 �'vH�n����&���;7]��G%�������������٭�lNk[O�,K�����ٴ�Kı?g���r%�bX��w�ڪ�bX�%������bX�'����kD���5�����ֶ��bX�'���ͧ �6%�b_}�kiȖ%�b_�ﵴ�Kı>�w=��" �2&D��5�ԶQ�evm�7,��,K��kiȖ%�b_�ﵴ�K,K��s��r%�bX���{6��I�L"c���6��RI� uW1�1bX�%�~���ӑ,K����{6��bX�'���ͧ"X�%�}�}��ŃX5�Xw����*N�P���ND�,K�k���r%�bX���{6��bX�%������bX�%���[ND�,K���r����%��\=�F����8��j�]�¡v�uua��tnьѶ<�Gok�.�8�#�:�O5�5ㅸ��6�A���	�W�9�����t���ҙ�Lgl]��� �vu��Ռ'E�:s�I�JΆ7YӢW���ke�6���-�ŷSƖ�Gkomh�.�c�z^��f��q�#�X1�D��N������2�d`�6[d��d�f](tn5�]�1����p%�s;�ᶛ�Ia�l�]1��Ê��Jq�O绽������u��ZZ��Ȗ%�b{=���r%�bX��{��r%�bX���m@9ı,O��}��r%�bX���{�\ճ-ˆfk6��bX�%�}�m9ı,K������bX�'�k��m9ı,O����ND�2�D�>���պ���i�Z�Z�ӑ,KĽ￵��Kı>���fӑ,P���{ٴ�Kı/��kiȖ%�b{�ݹ���I-Cu'd�p���0��==����X�%��>��iȖ%�b^���ӑ,K�Ab�3������bX�a������$�2¦�۸q`�ab~Ͻ��r%�bX"����ӑ,KĿ}�kiȖ%�b}�w�ͧ"X����������I��9-؎�$�{[S��sr�q	�u�؃�y��ܷ>}	��n-f��$�Z�m9ı,K����r%�bX���ٴ�Kı>���f�ND�,K�{�ͧ"X�%���w�f\����!��m9ı,N�{��r�����da ���p���I,�4ʐ���!�ҕ($#Q�D\mK�q�V����0�
���b9��,�/�R	�S�H���k��ͧ"X�%�����m9ı,K����r ��bX�|j��Z��J)B%-��`�a����n�bX�'����ND��D��"_�{�[ND�,K��fӑ,K�E��EMSUN�t��|L"a'����ND�,K������bX�'s��m9ıU,O���Y��K����+����7,�ı/��kiȖ%�`�w;�fӑ,K���ﵛND�,K�{�ͧ#���ow���|���[�᮷�3 ���p�띵���8������������c�tt���m�8�k�k���m9ı,O���iȖ%�b~��ٰ�Kı/�ﵴ�KĲc�m'Ε0n�*
mӹ���L"a}�w=�ND�,K�w�ͧ"X�%�}�}��"X�%��w�ͧ" 1,"��=������FXT�R�59ı,O���ٴ�Kı/�ﵴ�K�$!1�Ő�	�`5�gH�\�A9�R��#��c)"��Hb�H�MkD�K���:����+u3!�r�@ƍ0`{L��4���[F'��J~�f��4!������#�#qfA�b����w5�ԕ�a^ p�i`Bvk?�0Z� �c�RD���B�WT����ù�"ej�E8�����1�j�w�Y��ê��ӡ�\-(�sA�E?_�Ƹ#̷��a�h}Չ��&T��7s9�LX�`���>���mE��J�曆hq��ٰ57�v�]~���&o�\\U�o�1hi�A� R�cI	�)BT��!rT̩a	�a�2�0��3F�E�.��t��Q����B � ��W�N����z�t"<@�Z�'1P�(�F��,L���>ͧ"X�%������>&0��Lnr/�*�B��%M
浛ND�,,K��m9ı,O���m9ı,O���iȖ%�I�=�w1�0��L"c���6.��J�5!.f���Kı>��ٴ�KİD���{6��bX�'�｛ND��Dȗ����ӑ,K���|R���g��:���3]�kTn�:�*���v�rK0��-q=���k{��T�#�v�Ñ,K?����fӑ,K��=���ND�,K���[�B���,K��fӑ,K��u���&��k.����fk6��bX�'�｛ND�,K���[ND�,K��}�ND�,K��s��r %�bw��{�k5&[��n��ND�,K��}�ND�,K���6��c��Aș�?����r%�bX�g���m9ı,O��/}��%�tf��f�iȖ%��'s��m9ı,Og���ӑ,K�����iȖ%�~� ��RA���%�wٴ�Kı=��=���34۩5��ͧ"X�%���s��r%�bX��=�fӑ,K��=�fӑ,K��w�ͧ"X�%������1�{Z�&	::�Ϯ8u�����㪋Q�l�E��`Y{M��e^�{�����\���u����Kı>�����r%�bX�g���r%�bX���ٴD�,K����c�a�D��"����*)�KVۭk6��bX�'���6��bX�'s��m9ı,Og���ӑ,K�����i�bX�'�z��}����N�\�m9ı,N�{��r%�bX��w=��"X	bX����m9ı,O���m9ı,O�5o}��5&�e�d�Zͧ"X� X��w=��"X�%��=�fӑ,K��=�fӑ,K��w�ͧ"X�%��|����5��l�[%��`�a����q`�X��{�ͧ"X�%���}�ND�,K��絴�Kı?��}��~���'V��^&ç�볅��nJ�{����t���N��N��}�u��oN��r
kg��'�t�/W7vc���ѧ�@;P�G�6\,�q�W��a���jg�SsX
�\v*��j�u��܏Wn�C2鹸�����+v��#���<Q�!A��6����c���i^����f�Z���Оۦ�v�S�'Tu�/,E��f��i���L�eΪ��L�	�Ғ�麛�Y�����N��w[s�3�۵ =l����m<'Uߝ�qu�~�i�-��k6��X�%��?���6��bX�'s��m9ı,Og���ӑ,K�����iȖ%�b~�E����E�L�]fk6��bX�'s��m9 ,K��{��m9ı,O��{6��bX�'���6���%�b{��n{5u�fi�Rk35�ND�,K��絴�Kı?g���r%���"dN����iȖ%�b{=���r%�bX����JEj%�	��p�����;��iȖ%�b}��iȖ%�b~��ٴ�K�K��絴�Kĳ��{���:���ZrY�q`�`�}��iȖ%�b��;�fӑ,K��{��m9ı,O���6��bU�X{�|�L���G[m���e��^c��l�8�t;��EM���[�A<��ĺӠ�Zͧ"X�%��;�fӑ,K��{��m9ı,O���6��%�bX�g���r%�bX��{�]a�5�.�$��m9ı,Og���Ӑ�yC�DY#�.� �x�9ı>�{���Kı?g{��r%�bX����m9ı����OҲ��+��w,��O���6��bX�'���6��`(�%��;�fӑ,K���}ͧ"X�`�||'���ʫN�7,��P�>�}��A?^�ٱ$D�~��n	"*�~ϻ��r%�Va��h��c��T���,�8�k���wٴ�Kı=��siȖ%�b~ϻ��r%�bX�g���r%�I�L~���̃�S�U�[qP�����V�\�6+�;g[O[x�]q�<����M������~�����o������q�����?����r%�bX����6��bX�'���6
�"X�%��>�iȖ%�b}���R�Z�m�%U۸q`�`����6��bX�'���6��bX�'���ͧ"X�%��v��NA�,F��߇��,��ʛu�훇`�X�g���r%�bX�g��m9��M��� � P8�"dL�w=��"X�%��;�fӑ,K�����-U�T�[��nX5�X5���}�ND�,K��絴�Kı?g��m9ı[��}�ND�,K0��o�U��GB$훇`�a��s��r%�bX)�>��iȖ%�b}��iȖ%�b}�wٴ�K�k߅���V�݈D�,i7Gb-�Xgsm�Cjw��'Pq�Ս}b�c��⽄��Թer�-�X5�X5���~��`�X�g���r%�bX�g��l^D�,K��絴�Kı;Ӥ��55�j�d�\�fӑ,K��=�fӐı>ϻ��r%�bX��w=�����L�bX�g���iȖ%�bw�/�kM�X���,�8�k�k���7D�,K�������~�`�%��{�6��bX�'���6��bX�'���?�e�ŵ,���oq���x��������Kı?g���r%�bX����m9İ;�\5Y�}�ND���?}����V�[`�[��Ë�ı?g���r%�bX��}�ND�,K��}�ND�,K���Z�r%�bX�c���{YIluf���I�竦jíɘ�1�ܕ<������s�2��{�������IR:w1�0��L"cϷ��"X�%����ͧ"X�%���}�l?�~��,K����m9ı,������Un�T��	�7,��ù�}�NC�  DȖ'�{�Z�r%�bX�g���iȖ%�b~�wٴ�O�X�DȖ'�5o���ta�4%ֳiȖ%�bg�����"X�%��=�fӑ,K����iȖ%�bw>�w1�0��L"cH�s�Sn�'U�ֶ��bY��B���o��ٴ�Kı;���m9ı,K߻�m9İ?��?����kiȖ%�b{ޒ+?UU%��;���D�&1���iȖ%�a�
��}����%�bg�����"X�%��=�fӑ,K�����Teh�Y
�D�B�X?ߵ1��Z��u�UrK
qq�;q=?���}�sGgj�ն�(f��Z͜���Fz<h�F���C�D5/"9.+�&�1rvP�4�mD��SXl��cQm����Y��@�=�� q3nn�*�먩��@��;�E��/����z��okN#)�n�`�1�RY�ÊR��<��)����r�46f�[�v�ʊ�U[W���$�K�X�W@�C��lӒ��ٖ�f�5�WEՔ��S�>���s��l��ͫ�U�ӈ�ؓ����|�]�u�³�������d�������bX�'������Kı?g���r%�bX����m9ı)1��	>t�@�"��c�a��=�ﵭ� ��bX����m9ı,O���6��bX�%�������#X5���~�)���"V�p����,O���6��bX�'��}�ND�,K��}��"X�%���}�m9��D�gE��I�QN�*b�N�>&,K�?g���r%�bX��{�m9ı,Og��kiȖ%�� $"ew~w1�0��L"c~_��)*��UQ.k6��bX�%���[ND�,K���Z�r%�bX����m9ı,cϷ��|L"a��xw:n�h��6��L��i���g�kg���8w�Dn��uY9u��4��6��(J�۸q`�%���}�m9ı,O���6��bX�'��}��B	�&D�,K��������{��7����?����ʳ5|��bX�'��}�NCi��~EҢ�Wl�bX���iȖ%�b^��kiȖ%�b{=�k[N@lK��tgUU$'	U;���D�&1���6��bX�%������c���"dO�������Kı>�fӑ,K&1۷��UK�'I�N�>&0��W"g}��m9ı,O�������Kı?g}��r%�`"}��fӑ,K�������ˢfM4їY�m9ı,Og��kiȖ%�a������~�bX�'�����r%�bX����s�D�&;z�%¤0B�)���G5��y��)[�n��-u�݇I�5/k�gۛr��|��)+��֒��m�8�k�kϽ��r%�bX����m9ı,K�{�m9ı,Og��kiȖ%�b{����n�UeI���Ë�k��{�ͧ"ؖ%�~�}��"X�%���}�m9ı,O��{6��bX�'�~�j�ڥJ�!	�7,������[ND�,K���Z�r%���$���@j�(����`�,ND�s�6��bX�'���ٴ�F�k������-J�#��XX� 2'�����m9ı,O���ٴ�Kı?g���r%�bX����p�����==���u*�����[ND�,K�w�ͧ"X�%��=�fӑ,KĿw��ӑ,K��{�ֶ��bX�'���jfWW3[����,�s�u���6�Kǈ��{�n��U����w�J�U[kiF�ݳp�����;?}��r%�bX�����r%�bX��w������dK��{��6��bX�'���?�jt�ED�vK7,�����{[NC�DȖ'������r%�bX��fӑ,K����iȟ��1`������QH�B�v۸q`�%������6��bX�'��{6��c� ���>�{�6��bX�%￿��q`�`�{��qRWYl��%���r%�b؟g}��r%�bX����m9ı,K�}�m9İ/B0��Ƣh��M�'��rD�k~�p�����?}��։�VYRn�ND�,K�w�ͧ"X�%��￿���ı,O�������Kı>��ٴ�Kı;�^�s�d5��fF\tS�1d�<���n�xM�]��ټ��um¯BUh[�f�v�3������,K�}�m9ı,Og��kiȖ%�b}��kȖ%�b~�wٴ�K�þ+~��+N�#��X5��b~���ͧ %�b}��iȖ%�b~��ٴ�Kı/����r'������w�������O����sR�9ı,N���ND�,K�w�ͧ"X�b_�����Kı?{^�w1�0��L"c�4|QUT�4�$��ND�,K�w�ͧ"X�%����ͧ"X�%�����6��bX��v󹏉�L"a�qΪ����<�fӑ,K��}�fӑ,K���{ٛND�,K��}�ND�,K�w�ͧ"X�%���ߒIad(���	`��ՈHX��s� ��:���I=�P���ROx*Q
���	�*o>�a�ZX�# ��,�����!"I ��@B��#H��s�/z�d�s1�����h� ��%�!*D�� D�������\ٵ�B��@#(7�?K�)��ujLB���iiA{D�$"B-�X1��`1J� 	!5&�Yx�$9�@1g�$m
f,lM��ix!z?/�BF6�  �!3r2Yb�I;'f��:�WuZ{�Z#csث��1�٤������m�؍q���w8�6�[���:j�m%]m3H5�uvΞ�eeMM�{l�6����lX���OS�S]�ڸٽ���g��j�x��H���Z�i��nA;8v�}P
J����%�u,��6�ږ*���v�&y����0��s�p��[>5K8͇��.���M %�6%��nx=m ;�Zr �5�z �I:^��k�Y�J놔���v�`�m���+�]$v�ɤ���]��g�'/9-��Y�X�^uv�N��t[�#{:�w�J݊��-���E:�1�6����e-]-9��EUl�nv˺틑�^�{H�[�8˵��)�v�hw��_K�@�2x�爙��B����h���n��q1�j��mۏ[������V9QT{Z�v��n@敭����m+`�\�$k��ŭNP+�]!&a�Jxs�V�֪�tT9�e���A�V�S9D��n�;R
�fצ�u��㯘�h ��7h�Dwa(�1�ģ�Q����T�9G0V��@�*<K;�;=R�pP�c>�VQ�1�U�Jl]���^K,��A�X�O8�3�e)i�tl����u���{F�U�sxg"�RB��֑.`��#��m�a�ۧ���@4{[�g�ڃA���v�'kH��('�{,n3���c��PqÚŎf:#���0�
�C����^Yi؄N��zK�F�h�m��r���������s�3\�vv��M����x�a��{u>�ɞ���8ݟfy�[�N6	vy�l5�c��q���ݶdfn�L�;^��E:x%jVW.3���{�#�wk��rP#�u�^��s�XC�2�C�:![�덎xgۆ��:�N�6��4�d ���r�.癇Z����s��힬�]��/.�Y�܇Mö[�I��wbZ�$�J]��m�r�\�`�t8v��b%�H+�%�jfjS[T`�SHQHhS�O�"=:q ~㨁�A�DT�m�J��T>:���UG\���HZ_�-j��uET�);N �]u��I��%��Hۓ��p�vZ�@��n�\�iÙ�٤�L>�\�z^l��z+[0k9�]k.�ƻ]�qk�s�5v�@`����u������&�7X�٤g8z�%�7�v�v��6������Γ�b� 	m�2���)�Fv��l��s����������Tݚ�ǂH��{<��m/�u�;v�������a�� m�Y�9���<�'v`v��)n�ma�&��v�ݭ�/�w����Kv]�������,K���{ٛND�,K��}�ND�,K�w�͇���"X�'�����>&0��Lv����2�UIt޳6��bX�'���6��bX�'��}�ND�,K����ND�,K���fm9�2�D�=����.�j��I-њ�fӑ,K��=���r%�bX�Ͻ��r%�bX���{3iȖ%�b}��iȖ%�b}�]�Z��f��3Z!	sY��Kı;�{ٴ�Kı?{^�fӑ,K��=�fӑ,K����iȖ%�b~�ս���4K��d��ͧ"X�%�����6��bX�����ٴ�ı,O���ͧ"X�%����ͧ"X�%��ç�%��8q��՝����8�%����m%{v��W#�]qΔ;v�����M'5/��D�,K��}�ND�,K�w�ͧ"X�%����͇��O�2%�b}��~n�>&0��Ltoo�C�T��e���r%�bX����m9�t2��
�q,K����ND�,K�k���r%�bX�g���r%�bX�}����v��Rr�%��`�a���ͧ"X�%�����6��bX�'���6��bX�'��}�ND�,K﨟ߚ�QH��Ke�p�����?{^�fӑ,K��=�fӑ,K����iȖ%�bw>��iȖ%�f{��qRB�[kiId�nX5�X"co;���D�&���5gs�>�kz���jQ�y�&Hܘ)�����ٵOq(8�zZڳFr_Om���Ҝ�L�8��>]���k�>�V����� ������]TU7P�T@�;�]��D�${�sv.�v�3]����n" �O�iǠ}]��W�զ� �`S�*߽�ԗ_��ԗW��UqL�
I�$o@�^�������a��]���S�EP��Ĝz˺������o@�^�@���&�cs�!�<1Ό��5��z�mv���+��

x��a�c���7�58�q����Wkz��z˺��ຢ9�#"nM��})]��-�v�fՁ��[j��5�B$7��.���uz~H����������ɂ�$x	LqӰ鈕���=��`}�u���(����e2�}�h�34k��H\=0���0�aB2cL�!#!�T�	`HIx���-���.��߭V�WRv�X'�}�f��v��|���>]��o����q~y��]�k�[M���T�;*�V,n�)��y�0s��svc[a��iI4�����^���@>�@���)�!I#x��.���G��;>H��U��}���S�-�NSĜz˺� �����o@�wW�wt��Ě��M��?%�M����>Y���f�1��QN�Ɉ�j94����fy�������}��`9��pD̙@ڢ�MR��wfG���vd����B��\�#ιJ�#&-��0�w9�i-�]��I�l�h�\y�k"�v�q�؏d��]Q����(ֻ[�V"�; ��`稟(흞*���8���.�ؤ�C�Q��:�2WmN��:�vछnۜ��{;k���B$6��6А�7oeg��v{nH�;oL�i`YٛVyٝ×���\R��ȰC�^`��cq�u�:ǣ6#�u��6�m���n���頮�S�ɭ�]<N)����!��k@��@�wW�wY�}l�h��S�d�����@�wW�wY�}]��.�����$f�*�E*QP'N�=��`}�u�=2���@|�5�#2a"��n ow)�z٠|������<��*��dHRH�9#z�u�˺� �����o@��W�&�Ʒ�ju�cq����cq�ov���E�(��6�x����dm('�8��uz�u���ށ��@���1��5�fk7$�~�������U[g��[�<����f�蘉�H����n	�DC�ɠ{�����mz˺� ��4��uLnd����z13+ϻ�����33j��^�vz��f,� �8��>]��vmXk�n��n�:&=�h������u�/IM�5n#��rm��7]A�1�k���ɭ�� ���m��۰��m�~~����ށ�mz˺��ƕ�#� L*a�N��^�w�11	���V�z.��^�U�2,JG�$y�'��{��r��ss��~p.fT
�W"̪����Y �"��2�0H�� ;l��=���{���)�F�NZ�N���ί@��^��v���;���-���6LI�'n=˭z��ց�ֽ��^��1s0v?�pxn[Ɉ��b��-r�@ǲN��;����/�Q�x��9{C�18��R?�����Z�Z��uz�Z���*���	7�h]k����^��ֽ�ek@�o��G� S��.��.��[+Z�Z�uR�D�2``�z�Z����˭zg��A �+@�'�@�A��]������BI��t����������;�7]����td�n��Ŏ���U��0���������W[]�8}c���9��a&.�
e妴.��.��.��[+Zg�Ʋ���	�=��^��ֽ�ek@��^����1����qF��<�נ}l�h]k�>]����UU	�E0�UNå{����;噮Ô�3=�v�B�U	��p�,n'�<�נ|���<��ܓ�rO���+����"�HFAI����uX5�3�I6���#	��y��N;I�������%�iQl]1�G��nK1��ŷQtE�)�tm������*<�tn��&8�vt{U�L���Y'1��E����S`y�x��6=�x�cL=�ku��H��Yn�48��Ձ���'� ;f���Ǌ
+�����=:H�t�mv�e���,�����[s0sع���&��K.Mas.m*�"16{��o䝃����b�f�7694�#�,m�S٧����T|��rڻf���ع��|���<�נ}l�hVנ{��B'�8	���8�]k�>�V�+k�>]���5]���Hl��ӏ@��Z�<��@�wW�r�^����U\S"Ĝq<nF�+k�>]���נ}l�h��Ĳ��$$����@�ֽ�ek@�m����y7��	1�P]9J�<f;I����3�v�En�K&�N��lH��%�p1	�ۏ@�ֽ�ek@���^��xs�R9����E#�>�*���@�!$��$X����+\
���o�ܓ�����>����U185�%���Z��h]�����>�V��]$�r#"`
2I4�uz/uz��ր}z��T�<����``�z/f��f'���|�ޫ噮����?����J�it��[j����s���ٝv;;���!v�:���G������5T����XۛV�3_L�|�Vo=��~k�dX��(�H���o�BF��v���A�}����Шh�M@T$НU��3]��ٮ�L��#N��d�H\���	KX���l	��! "�%Hѕ`m$`<�>�2�C�!?kH�AV��OߕX\H�%A��aV��D��`$�-e�H�H%X�A�B�cL�1�\��ł�;ʱ�f욒�f>
��5�D%e�L���
��`���)! �ey��q�F9M�i�0�N[�겷����ǜf�B}E���t x�*�	 n��`�L�V˚"-�ݤ2FD�O���lpYɉs8�kt�HD�-ئ��� $Wa����8@���!���0�G6�"�����%e��҄EHM� C�j�#1J�"�E>D0�h���W�;�_������(A����@>�Y�{�1X�Ʀ$�$�ǡ���o~v~�_� �fՁ�3]����Gs��d�Ǡ}l��_u�.��
�����(�x��&���hY#������O��N]�Λ�u�첼�y�@t�'���I�%�����˺��uz��h�I��FD�J�UX�5��ba#�o;��ŀo���U,�N��2``�z^������@��^����vL��,���ԏ@��M ��4]��x?�$�0H�1#`BTj+�Y���@1��ݚs0檊dXۊ)��h�Y�r�@�빠}l����1�0 �֕��,\�ulw11�f�n@��	ٺ�a@�s��r)�@�)5HM��Y����h�Y�{υcS�����7�}�s@��M ��4]��D��$g8]���B�R)'Q`{����mX�5��ێ��nt*�P��2D���4�_�@��^�}��â%{���77������L T�T�.����h�Y�O�:���A���0�c�,�b!,
:,�!)�Z�ֱ��H�Kjw���ӧXO�t28��Z=#m��c�nvu٤v�����gd��5��39䓴-v�Y8��췸3��;0J�L7���|,���p�i���� �koc<�HۅW�^x��-��2�\/\���Gcv�UKvP��]�ή7jż�ݴ8��ڷ1�/v9.��'�֛�q�&�[��_X��qv(��ېI
9�$�\�]�� ̸�ɱ���Y�
_u���'U.�N�x�������9�.I��k�^��s"��&)���/[��}l��o�k�&#��y��z�8�j�QL��G3@��M ��4]���w4y�V��dLO#�nC@/��f�:ff!%��G�{���220*#[P�Bm'Ua�+^�;�z���vS@/���|+���9�8�q��w4���/�U�r�@�r����=��-��s<�-�ئ���d��ɏ[�n'+IVE�������f�����������<�`b���1���s�W*��P�(n����<�nfff�L!F@��a���UIT�c A�\HELIt�Q0�V�&G�;Q�����}�w4���;�t�?���0�LRG�r�@�u��>�S@�^�@��}��JVQڒBr�K�a��}�������h+�����=�����'���>�S@�[^�˺��������ڬ�13��"���d�s:gnݺ��z�6<���d�r9����m���H����Q�h+k�9wW�wu��>�S@����ѕ���O�����;��h[)�|��@��eq��L���f���}�����媀�f F��X��4���srN_����+fI"��"Nf�������]���w4��*��Md�T�7I�`|�u�:�y���Ł����Xn5�m�<�c��T�{H��4Z�t����ۓ�^�J��/���do�z.����h+k�>�UlȜȲb�0N=���������]��xu��F�E����s4���>Vנr�@�빠{�ʙTS�<�!��w]��3]���qa�~�(q)D1DD(#(6�@�"��HJ��/����C����.\�1�?1�&'�H�]k�;�n,n֖�w]�����t���sN�=�Hеƌ�3u�6������<�u����G��6�6Ɯm���z�M�mz.��ܫ�#�LR	�'3@������]k�;��_�=ٻШp�Jbn(.�z��@=�v��>���]&O� do#���נ{��h�ՠ|�נ}�ّ9�dRa�
G�{��h׺��n�n��"	����Vp�a��?�(�X�r�S�s�6ѹ�-&�������m�<uױ�Ѱ�p����1�v��ۇ:�N�.����S��tC�#<&�^�:�qq�"��Xb�%�Fz��]n�oserr�]k�Η$�
�͑�#���+}Od˱��B�(��K���VݔZSk�;����`�l�F*�{j���/q�7YQ�=&l�r,�v<6x�)�� Քc� �(ʑ$v$��g�;��X��rV�[�;6�E��=�^�/�����=GDO�#�@���|�נr�^��빠}�Q2��S�D�$Z˭z.����o�3�1"���b
��ӧ`j��`{3n,Wj�>]k�=jLi�m��â""af�}s�V�7]��7]�}�]�$� �s4Wj�>Y��Y��fmŁٜ[i�b��}lG=I!nl���eY#�g����2-&�յ��>�x����W���������9u�@�u��=]�@�u�d��a�2I5��k7$��������,L\DH�fmŁ�=�`|�u�{u��i̋&)0�#�=�w4Wj���fB^[��[����m��*e(�T�Nf���Z˭z.��U����D�ʚ"�%1����^�˭v�6�����`t��F�A��Ҩi��tb�1��ö��'[��N���W;�ӓR��N:�Y#���ё�œ�U����ۋ��WD|��{����P��8�����@�u��=]�@�u�@�ֽ �ʻ2650a2$�h����r����(?TŅ� j�0`��@�*��a�Z�Ћ��R-����׿nh��bq��c��qH�:"f%y�s�5os�=����=�eEJ����S�v,�vLf�}�߬�h.��L�B˱0q��rt��Վj�d�����k��&��yѬySc�t�M�1�2,����@�u��=zS@�u�@��^��6�ȣ"ȉ0S��=�Z_LLD�$yos�5gs�=���	�I���
�%L�j��<���@��^��빠z���݇#&����Oq��k�=�w4^���
h�� �P��JIe��*�+��!y�w��'��+��6�7$z����Қ˭z/Z�ዙ�X��ƃpZ�N�r�[^v�8�:V�5Zt�:n�t�K�Rkb��8����2`�dI���g�@�u�@��^��빠w\R��Ɠ"q��������5gs�=���+K��I��9�G�1)��ֽ��qgD���Ł�����Z���E(�Ra�
G�{��h�)�|�ס�3?���v��m��)��J�
u�+M�ֽ��z���0����0�p�5�|փ:��o����'��X�.�Gn
d$�j�`� �bKS5�!��I�T���dB���e����}���PYBd�	e�J���1���0�NC�m #��R�:�B��qLH����1�l�!BPM<��֟�k_���}�f^b�'�@�Œ��B0K?~�Iv��ڄ# �no���o���v�(A�5~�!bL���7������X�-��޼hL\0HGEöN->Z��;[x��FŔ06�C �ΰ`G�9�5's��q�'	!�<�_>ۊ������q;V ]�?oxH�w��G�^�����3�?1Z�ʂEJ�����x�B�5�߮�&�Q'�	���F2˄̫��E�V�&9
�e�
��LC3g���ڕ��  ���8in'�m5�d-�'=��=%3��huz:]�Ok-ѽ�f�Qm��<Vwr����Ӷu��9��	]����ܜ�"gu]���c��mٔ-\������4l��+�������򡷶6�q�Z�:.XMz]���1�ط`9�ٚ��[�z��:X��PUu�)��6�1v��{Mf�X�)��-v���'Z��u�4�nѭ�IvIqt9wPg��'�1m���u#��0k���q�؄�<�PH��v�P�Α�:Z�;aM����ݙ^g��kk8��mn{W&ChЎ��f{��{xvۗ�^ڈA6wXѐ��>g0�V���7[]�)Y�AN�:���.��W�4���Ѳ�$<39M�v��S��u����;r�ɱ��m��9a-fء�k&��1N^a :��ݍv�l	�6��@�@(�g=;9�rj�%�Y��	� aq�w����UV���ND��&��ͧ"�n�bG[�S�K�R�U�ڪ�o,�!͎�M��Y�� Rҭm��0pN��`�o���=�n��۲�3�F]gb�c;Y�7�!�����Z��P�Uܥ�6��\��W
�AU�Xq�띜Ì�*�tV7@/�[ܞ��M����'���Tf\�-��)�\��k���]F�D�6���Uޚ���{sĵv��Ncu�s��M(�+h��v�&�^������L����pE�z�ɴ�f���s����=+��xx^h�͞�9�֣
'A�A�V�*�ۮ�h&���=l�I��ޙL��i�s�e�[t�M����j��\�����r����4��dڥA�wY�I�NX�4Ít;K����8�r>9tv�l�θ���Bgm�'[V���7m�x,ї�M1�v�ʝ�m�V��bty�g�,�y�b���Ԧ�T����S�U�h��^Z�O�@a�d�l�fY��	�l��p��p���qg�����Ҁm�ځ��?�T6w�
~ a@^���"��&�1���=G�@���C��Eٔ�/�hӧHk^����:�e���_9�q���X�خ��N.6�k`�yD����+�V���&&��#7\Mv�h�aA�2�\q#�6��e	MwA�y�x���˳�u����6m�Q��=�{zu�����F3j�31о�g�Ն[��t)�í.�t:�t;G<;�xz�g�����f�s�J*�h��dKF�Ў٠��H��0�0���7Ic�F�Ν��l����L�ier���c;��g�-�\:�u䚆I��LL���B����W�v/n�ٛq�? ����݃Q@?��idI<rG�r��@�u��=zS@�u�@�=�U0ss����͸�=�ZY�1	yos�5gs��kאo2adI��=zS@�u�@��^�^�f��\R��Ɠ"q��7E����`t�F����q`{r���Q�����-�tk�55n�[4<���w:�tQ��3�Z�E��l`�6��\tÀT�S�Y��fmŁ��Ӧf'�[���殡�QJ*)�T�g�ٿ����d�w[��r����r��@��x�HȘ���9��Jh.���k�=�w4ϖ6ʢ	J"dR˭z/Z�w]�ץ4�9�X�D��$z/n��j$�����G��mq`|�u�P��ɿ5�w	s���]*�v��f;I����&���qN�NnFę�$X�.�p�UN��f�Xܭ,�n������v�?� �
d��'3@��M�ֽ��z����qK�i2'M�t��7]��ۮ͘�"$�& `��#��"߻��7$����.y{�T��a�n٩~��>���o��ץ4�Z�zֶcNdY28��H�w]�ץ4�Z�^��J�X�l�#r9�D�$+�M��E�f�ܾ3�*D��w;�N6��Yʯ7I�c��G3@��M�ֽ��z���y���TA!�DL�C@�f뾈����Y����ە���" ����x�@��^��빠z�����^��{���1�n'%;ٛq`{r��>Y��="&r"d�32�a�w횒\]}
��""Nf��Қ˭z/Z�w]�ߟ����n|��it���'�o��r��t��6�����Or� :yCG8HΆm�Q��<���@���@�u��=�)�}�]���LY<��^����#����w~���ֽ�h�!9�d��#�=�w4z�h.��^��qco��2$��L�=�)�|�u�^�v�w��(�è	J"D�����^���@�u��>�֖1?f
Ѩ�!��	��8u8�ԛ���=�nn�vf
ݭk�z�����c��vv���d���żmdKۨ����.�lv�<�:4�J��.s6��g]���m��T�Y.���g���܉�V�픸��v`��ۋnh {h�ƺq��l�7'l�ȫ���gc�����M�bЏ;m���� ^�ƫ;R�����1�U�
;�m��`���wvz��>�Y�+�5�-,�뭏;�̔޹���v[�:-��nͧ��`���� �x��|��z���������^��^�Ǔ��Lj'$z�������>Y��/f��1	�\��4�&h�9����h.��^��w]���15�8����ֽ��^��빠}�)�}�W�O� dx�JG�y{��=�w4�kK噮�艙��Z�|�j����;e��e�'qӲ�/Y�퍤VO���W���Bsɒ##�[�s@��R��fk韐b��`f�M�}EEU��[V��߯�w�Ռ0X`�����F`R�J@ D!!�D�TK���K7]����`{2��<���!�DH���>]k�<����	f�q`{:��3 �JjZb��H�/uz���������^�޷SX�<�����)��빠}�)�|�נy{��-�1��ǀ���N��d�n8!��[��+�C�4�t\X��dİ�H�M9�"Nf�������^���@�u��;�GbQ#"`�����^���@�u��>���>�ԧ�dXA�
E�y{�П���74`/�U7RB�G0��!!ȋ�?(��Q�j��1vs�7ۣ�B�����H�w]��>�@�u�@�{��>�ıXL�)��9��}V���^���W�{��h�Yث��6�/5�.���N��:�:-b�ݝ�خNRBz�M�F�Y	&A���-�ֽ��@�u��>���9E�S���<rG�|���bGu� �Ϫ�>]��z!�9��q���=z�h{�4�Z���� �=��nA� �s4����ֽ��C�33<�0a�'��I}��~�8�Q+lp�>]k�>^��w]��t��}�#�#�bxL��G����2pSm���oG=��E[��n�I���ytv��MU;���`{3n,��WD�|��{�����=�Rd� ����}V���^���W�}ō�v#�أ��}��h.��/uz���}�l6(*(m��IUR�處������`{3n,��U��SP�T��5c�=��@�u��>���n�""4���N��-�*j�*���LgV������~dvZ�N������k��MΞ���,s:3әֳrVhMڹ�u�v;I�4lJfl:���{T&y��mrJb6	uk\�>�wfv�k]&���I;\t�-E�b�b֭�@8:�lݗ�sD>ݝȻa�%��8��9�Y��7n�.��ѳd8:� �8�:��׷9/J���'f�혴N|f:7���d�0�0f��lL���=n�V�uXKh���z��mC��l=�D�豴��C��ɞ���3�������Xy�囯������7��x28�7 �4D���>�@�u�@�{���ۋ鈙��ފ}HMR*�Lt�-�v�ٮΉ��w�,c�V�f��Je((r*j��/f�ٗs@�Ϫ�>]k�/Z=�NS$,JG�{��hy�Z˭z��^��v,X��x!�@ɋ$C��t��z�au��GX�;�j���`v:ܤ<�]7����>�h.��^��w]� �ղ��6���-�ֽ�0���1X!E�������W�u�s@��ՠwaѬUO�������@�u��>�h,�v�L��Y%N���a�30�w���������`y{5��z4ѷ �4D���;V���^����`{3n,����-���h�T
�NcX�l	�@�u����cwNR��+�qK��W�O��p� %"�+���<����ۋ�=�`}�k-T���ȩ����@�u��>���>]k�/��'��d��޲��s]���Y���I>#�!���3L�kO1�ђ�ѭ�7�/�M���ۋ�6�b��p)���a�l���]0��1u�B�|�k�.i���;d�;˴��~H[��g��8Dn��� ��'�d���T�1�aox��6 m�� .C��n�0��]9�'6��)3[BGd��	�U+L	L7�lMmڳfFF��)
�/�y5y
Ǌ����*�D���� i���A"��4��A\"? F
�㢡T��D�)�W|��;���}	�TӇ�TS�J�
uw���>]k�<�k�=�w4�Vʈ �#��>]k�<�k�=�w4z�h�b�Li��cɍ��hcp��[���n�I��l�4�1���!�����p�X�����9#�<�k�=�w4{kN���;�Pć	tЕ:�N���͸���H�������`y{u�ǲ�m�)s4z�h.��^�����7ЦI�����^���^��빠����A8�¤�HB��F�2LL����3M�Z�n)AC�SUN����@��@������^��e�~}�`�u�:,Q�Vo�3����p�*⎔�Nq�]��,h�\�^�`��<���=�)�|�נyzנ}�F�7�QN�
��v�����DD$yos�1gs�<�5�DDL�寚L*(M�b�*�����`y{u�Җ-�vgWdMB�Rܐ�U;�ۯ@��@������^��gLb��W!�G$N=˺�޲�˭z���7$�aP$ R�RB4(Þ���h�U��h���T�OH@����9�L�v[�g�ƭ��h�݇�ۏ6�Z��!���3n�&�'0��ٳ�˰�/u�OCv5�yL���ڴ��f���A|����N nF]qg0�8ͭ�]u��닫sh�n���A6��z���ݙ�3�hvz,��'h��:qn���9o��@�,��mu��KԒ����3{����{����r}����wͷ<�[<�lY�v9��}�-1�1����;��]l�X�Q-b���F�����>]k�<�k�<���=���I<�ЦI�����^���^���^��;V��Y�7�a�Q9���^���^��;V���^����t�QP�PEM	U;����;���@�u�@���@���<n��&�ؔ�@�[^���^�˺�˺���5�����8(�d�0i�+����'"�v��)��p]����n��d��ڦ*T������`b��`yfk虉���w;v��r�nHt��;������"E
�Y����䟗�z˺��,�,O
̂Q��@�wW�|��@�wW�r�@��٦��*��©�v1ϻ������˺���^��.GbM���U;�y��ř���{u�-�}3������ߤ�v��� �����r���t��f�VnT��Ҝ'K���v��Y�@���@�zנ|��@��U�^�b&H7 d��R=��^�����.�vc�V,�w�3)�����*�L%T�.�v��U��	'�$�b�!! �!2$��2ȉ�Dt�PIm��z�~���֓	�M��R;��Y���[����]����`gaѬUO���jb"�9wW�|�k�>Vנ{Ϫ�=li�1��o?���mt�5�,�O`�1�;�Z�z9�3��ܙ��c6�8�X�
A$�G�|�k�>Vנ{Ϫ�9wW�U����H���H�;廮�fa#1�+V�;���}2��tS�I����)TU;1�+�uz�ֽ�mz�uf���E����a�+^�;�;�����r< ��IBĨ�A?k_uhܯbɍH?���@�zנ|��@��U�r�@���C�j6c�Cw`��$H��Q�Kc���N3�\W1]�o]nC<G,��5�.�b��������m�>�@��^����@>��i0����G�{Ϫ�9wW�|�k�>V�3 �j��䆪:�`b��`|���虔�����yX��!Bpk2	'$r=��^���Jh~����w���9qN��T�*��`|�u�11۷��j��`j��>�>�D������u'L�k+&��6S̝E�\�����EȻlzr�cnvl��2�Nͻ{O�8��7XU��g2t���2Ý��%�sn�H��^O�7;�tC��,�N��u�����ns�-�ĤdY"e���s�N�8::՜ݓ�F�ig9�v��A��[cQl�`<[��g�{/Y��̰����X�Fp�۴m�v�n6�س2ŗ�0����CrG`ܑ f��7v8hv}�inz�	k�a��>���Ќ�;��]��-9In�p���5К���~�u~,���;�DLL��˻���7��R�R���L�E��3]�DJG,�v�w;s+Kč݋wHN�j@���z^��+k�/t��˺���4��EC'�
G�|��@��U�r�@�zנ�ĠHcl�QE�{Ϫ�9wW�|�k�>�ՠ}�;." �ȓ� �m�盭�w�ӥ�w �ώ�ͷ]K�n�]'��%��S9�˺���^�|�Z������x�����@�z׿���FQ�"r]�;w$���m��3]�D�G(�ˈ��T��St��ܬy�Vf����`{�dCɃDȦD�Z��������]�DLD.��V�އeKqJ)CF,�ŠU�^����@�v��}V��1��|�t�j���p�) ڧ.[�pGn��ۛg��[9��v��]�xj1��C�F�H2	H�˿~z�h�꽟 ���^�4��EC'�
G�w��~�r�^����@>/;ǒ�T*�UJ���j�5fk�v ��&&HI�H�%!h���B$Hp�""�-������3(F�R��UR�5fk�>^�v�n�����/�[�Fc���̘�8�q�/]vLDLLs����yX�u�����*m��k.qm����6���^�z�d�:iR�ʒ:�9uN43I�!�z]k�=��hu�@�zנ}��fD<�4L�d�@��U�Uֽ���`j��}11)�z�-�(����`r��`|���Y��y�����N1��N=��^��7]��<�a�sB�����蘈���;��m����&��T�Y��y�Z]k�>^��,�J�x`�XVt��r�2�|K�lD�����g\�Rd�Gp	�9�!�<�S#����
��>^�}13 ���݃hg5R����
�X�u�$ygs�9os�=��h�LcǏ.2bX�Ǡ|�k�*�^��>�@��zY�U2FH��S	�@/[4y�Z]k�>^��qrY�&"�Ēh��Y����]�{wj��b~�?N�@o, ���@���X5�bBw����^��{0NO��8}���q2\�_��p0Ni�0���ļ�8�&qtz���W���1f,��<	ˉ�0F���h�UF��	���1�⾃�tt�;�����0�O��tî��'�y��
?���H0��MC��4~T�w!��V�ՃV,t�\ISfG29��W�9�n_G۷�g\�@�0���M�{�+����y�7/��Fr?��LD�z����k����3$uϞ��$R"D�#[d;t�ZaP�2b��o{ڨ@����(Fl���8h��VRY`U���5�� c�3�C��8ɂY�8p.R���tK�S�ޕ�@F !shhWY�*Д�)(C�n������tCU��,�#mїF�����Ԭ$$`�ҥ��B*��?��	   6�v&zn����
�Quqׁ��@�[^z+�sI�;�A.[���P�k2�+��WÔ���]3��&>i]g�a�sJ���I����r�.��،�nf���=�;F��ח7 ������[M�(���)Մ�9���v,�[b�}�c�{6��t�{t���v�m���_ �6������7ppk�gnqg�s0�m��CYh��ˠy�T�kY��v.���.4˗s+̒8P�����zy�����"H�=�[��T K���J]uu��k6.=/fx�ŋ�����Z��Ƚ]k��x."���M����{sc t����9�ݽ^�2F����.n�n���dv�P�T��$8���͋���b�~��q��lr�ݎ� v�;���ByU��F3�\�q��|�m����hM�d�[n��
�izt{45v�;m�wC���0�l�pv����<ȍ���h�m����m�ۘg,� ����YF�-�(
X%��� rQ�ڄ���6�v���d"�	]��-<f����$m2���mm����;xi���y�a�I�����{���/1;p���t��[
�V�u��-k.'��f�+PkX�P:�R�I��څc�M7m�k<;�m��r^l%�i�r�=�:�(�n�ƣ�Oe�o;=�sb��\�v�[��Űnb�s�A����Ѳ�W<�La�#��]������^.�dv[Dn�BƤ֓�V8ȀGZYC�՞pպT3�軘,���R���sp{(#n׀���?F͸��ms�v���m��&+�q��^���v�=��b�ۘ8��q���u�N��N�ؓ�GH�leN2�,�OXZ�%J�m�ۻt�.7�3�zU{��*�Aνi{X�6pN0�+�ՆV7�F��'<�1��[�z�]r�hNjZt���ts�S��;���*	� �+9N�6$�
�/S;�m��C�8e Ѣ�3j�,l�D���<MDg��;����v��n��u�Y���Z�G��Gb����QR` ����DC�|+�h���Q�uO����ᄞ^ll}�Q�R�bvV2�
5�.�{M�Q��I��t��d܇�u���q�A�PRv9�r��q[�i���8�� ��n�84f��۞:�.�d8�F��\c��ɻ�,���ۏm�`]n�g�������i��n0��[-����vԙ�mu�8fzc�Ka�;��'�	�j�u\Ӫ{,��瞞]����ty�e�o8�����\q<����x�w���6\�m����;]j�3����2����JG�0��s�t�^�a��9��cB�^���z�ֽ ��h��ݕ�B��1�A'����@=��`{�5X�u��H�:�NAL��T���������<�`b��`|�k�>^v%�CpiE�@��U�r�^����@���ejJr�**�`b��`ty�s�]��y�Z�bˎ		� )!��i]v��Om�nK�D�l�n��$z: xgv�a�<�Ɍ��8�q�/Z�+k�=��h�נU�US$d�<0�8�׽�og�b�1�S0�FcKL �bȒ,F@����ʘ�H�r�>]����]��DD${O�?L��`�2)�$zs���˭z�{�����`t�M�qN)CIAI��>����{���}�����a�1��_�@�n~{���d��z�v����y�Z.��q�qb˱瓐�nqֹ�uگgul��쏘!ݵ��\�x�í�X�y�N���}����v��U��7_LL�D�������s�UQ:T�U;�y��fba#V�;����廮�b%#v����NX����V��v�{�Θ�� �"`D���F� @R0���阗1G'|�Ǽ�ͦ1Ç�1,q���>�hVנ{Ϫ�9u�@�<��H�x
a��<��@��U�r�^����@�ԍ��'v$x�cX�`lu��搓�=�ސ���p���<4�����]������������yڴVנ}�\zLoyD�8�Vנ}�j�9[^��>�@��^�"L2@a�MǠ}�j�9[^��>�@�mz����2&�bR-�����]�sr~VR��T�l%�.`ax`.�>�jK��~�F�j#���)��>�@�mz�ֽ����~v�q�W+��n�e!�����uF6ݹcp�ŹH�ܘ���֌�[��ٓ��>q�0R-���/Z�Vנ{Ϫ�76�����JuT���]�LĤU��zs�����zY�U2F8�URt�[��y�:R������ߞ��%�M��`I��>�@��^����@�}V��q�11G�"qh{��>^��W�i'���n�5�*�	(����[�W]���.�!�gi̠�.y�Gk�.g3��xҤ�-�m�kc .]î:���n+H�&u�g��j�8l�\!��Z���1���n�œ8ػu�ە��w6ӂ*�� �3Ak�M�Z�/�ݑY���Η�X���I��5�;iӊ����:q�z�����3���n5�ۧ/3V�-��-�፰F<R��50�e�®�,�pԶ����[�9�l�r%�;\��؛t����,gav�9mq��VN���/?��hϪ�=��h�Y�^,m6l*e&���V���3)�yXf�Xy�鈈��X.}IEU�P�LrE�w;�h�@��ՠ_;V�݇A�����L`�Z{��>��V��������[����c�~�D,i�&����@�v��}V�^�4xiVbV��3Q��X�9�R�:��zr�Ǣy�v���מ����j��mn�rE�Y2(����~Z��� ��hyڴqrY��(�AH�y櫈&&#b$@�6���U��ۮ������ڏ""�Z{��>^�v~����gs�3�325�P���A�2$���ֽ�Z�y�Z{��/6��Q�5��#�*��@虜��_ v�U����23tV�ݹ��r����q����,����W�g[]���@r��3������~��>�@/u��v��Z��E�X3��NZEC�+ �ޫ�=�`j��@���h�1��.2!cM97$���n䝿��܈j���v���JȨ�+ Dd��DDL���{�Z��}��`j��i۟�Y1G!�U�^������ՇLL������k�uP�U����H���- ��4�Jh�k�>]�o�~�z�[1�=�pPsI�`��Aw>qh^�u\ձ</S��؝<є��n�N��nmX�,^�}3? �u~K@����L�H5�D)&���M阉��Y��wW%`�ڰ7��u���f1�h�k�>�T�׬�;�)�yx\�K$�ԃX�I�LL�B�u�V��V{+K�GJ����$B@CD�/7��`n���~j�9i��ۛV{�4^��[*Z��#�"�o9�sp�Wk�7gOcAD�x�Q'h5Gpmt��2A�Gc���4�Jh�k�>�T�׬�*��j�܆!d����ֽ�eK@=z�=�������U	�P�I��S�=�\��{sj��<�`b��7�wn<��$q- ��h��h�u�t��L��u�V��;*QPUA���V�Dk����J�=��[�|DlR�	 �Ͽ���sF��!z�>�ݢǮ=[;�,�9�w,��Ż-�=�qN�W�C[h�c/n�%�O$��l��Xv
�{t�r/q�a��1� ��U�^��qʚKj��b۱W��[��^�����:�p���::�]<g���9���X�̮ʶ�
1�1v�&�ήA�rŋ̲V���5��t��kcel�թb"�E�8�����0F�q���H|�0]�����Pt;������wf�$A��G����e2�Ɣ/]�[�y~����������Қ���bY$�Fc�$Z�ʖ�z�4�Jh�ՠ{�X�j6cH�����z�4�Jh�ՠ}l�h�1��aq�$49&���M�ڴ��- ��ha�dS�bLQ�h�ՠ}l�h�f���M�����x4��9��Ra�pE�7_���w��ħ;�X���4���O;Y2���V��MLQ�x��% =��hy� ���@���&&�pJ 	K@;���H(q�]d���M�>��znIϾ�7��ck��~���(�Q���n�z�Ɓ����ʖ�wu���n�1��?��4���>�T�36�:"V�����RQUCJ�԰uE���Ԭ���_ٵŁ���Ϳ����8�y��Xj�hV *;<�ڭ!��Y��Z箂cu�G���S����&0n%����Қ����� ����Z[�ư��"��h��=l����������-Y�$x��r���>�T��2�<��z��Ǆ�A̪93>3_,J�
�0Rh�p9�p��B���`H��p\80m��#7��/9��DeeIh���p3&%��a��~(��fz_ ʍ�0X�0�F������?�X%b`�x"�w�~��v����8�|�)�vbF���3�X�-�f�,ڂ��at+���d�~0u��a)��H0��6Nb3�"j7N�����dL��Ɣ,���0��c1g�0�#���\��c����}q`Ձ3������Bv)���f��W�~1E���k{�o>��D�Ş1��dfx�0�ڤâ��y��\�F#E��EBO�Ο|ϯӝ��֮���9��c�~��D!���+.��MkC)B!`����p��^WJ���b�O�P@���C���~�:z�����D�:��
| ���C�8�A&f�c�����Ł��B�8�*�L�T����X�uX皬:b"egu�`{�]��L�J*�K@;��{�4[)�}l�h����f{$�b�}I���ui��zr6��[(n����t:t�:�s#�s�5�Ĝ�@�t���e4��/ٙ����w���E6��5QA,n�۵�����������˅[�� �mO�
C@��R�u�@�>�@�YM��Ʋ�?�kL`�K@=��`g��蟐f�qa�LY<D�1) �X�c���)�1 �m!2G"��� +�Zl0��������ư�c"X��@�t���e4��- �[4�f[�ki~�4�z�1�w:{t�L7]�����Z����g6�:��Ĭ�p�E��9뉭��?n,�kR�f�t����sk�0خ�9-m���jK���^�3 �����4�~4u��>�+�f$ƘHa�G"�u�@�t��zϫԗ{���F�EK���_�0��]�h_��@�Yb�u�@�TM��F52����v��e�@=�j��ei`G��	"I��K�(Zح����S��,�z�
:�j����b0�T��F|5�z�v����g,\	�^�i��n�v9� �Nֶ5�s��ƞM\�Ľq��ݝs��	P����1��ڭX�(\�sj�i%�7L�V�Ӣ���YY�/G3�I��ߡ���zč���#���vc/p��Ŭ=���X��y����ds������2���[bV��P3s0�Z���(!q�5�ė6t��u�ܒ�S�ݸ��љ�]��x�paķnIgs���m�����ٻV{+O�|�5�+2̎j��k�NE��f���M��Z{ki_DD̤f�1�Â���4�~4u��-�Z�u�@���ȞF���Ģ��=�ՠ_YR�u�@�}V����&ɒ$�F(�Z��- �[4��h�)�u��Љ��G��C$���L\ؠ'q��f˘�#<��K�����y��\Gj���h�٠_>�@�YM�ʖ��\�I��0�X��@�}V��$+�2	 :*o'k������ٻVf�M��
bU�?��Z��h��h�٠_t���R�_��r�Hh��h���>����h�p����cM`D<iƾ �M�>�@������kVL�L�t�
:L��-j]m8-�gng�j^��JA9I��������a�X0rO��;�hwJh^�� ��f��=��1<�(�&(G���S@��T��u��}V�G�rf�&ɒ$�1F�}�*Z���:����?P��<Tx"���f!7��r�7?W����[�cL*��F�Z��{���}V���S@��T�z⺦"d�dq,17&���W`~��f�����fՁ����F�{;:pX�<I��*��d|�B�N����{���m� �F� ^��g����ߛ@��T��u���^��乫���Q��Hhzʖ�}�@�{��>�Jh�>�W�5�!<iƴ�u���^���S@���h�S���E�	$�>^���Қ�eWrl0aHE�6V�$0�	 ��b� � �'�m:������K��~�tV��(�r�A����?DLNg_%��z���]���{����)���P�q�����mm�-��#���X��}g8㣧�,�֣�l�U��D�&(�>�����}�@�z��33��?u�{1,la&�Z��j���5X{+K�mjW�132��~�tj�T��!�n�����.w�K9/gW%`��35Rm�����ja'Jæ"W�o����X��V�}V��sW�9Q�Hhzʖ�{ٵ`}皬������HD͔)���T��ܿ�&�3Z5����+KV� ���� �dX�v(ݰ�̓>.�;v�0���1�f�p@u�[g6�i�c�`��k<鋴!g4d�(����D��g`֖�1 ϷVK<%�\ui�݇��/Nv�[u�j��7Y�l��L�LX���l�;"��s��v�R�Ӷ��N�nk��ʝ��༜rGm��ۭ&D�[˹Mc��L�\1`�t��Z������w��V+I �wn͛�8s��knN�Ǔe��L�swS�rǜ�a#29� �<�x���}��hz�hzʖ��g��w��ɬ"��I4s����������h��h�ȶ<S	�ɊŠ}�)�}�*Z����>�@����	8!E1F�}�*Z�u��}V��t���p�=��60���G�>̭,��U��ei`j�ګ�&b������a�#�}�D���*�\9��qt\�-.��A��^��4�]v���I�|�;�hu��W����4n�M��
*ja'J��3n.�<�%*ZCW-��&�M[���O� !(/�?��ߵ��?k�p�Y�|�*���A(��`����M�Қ��4�]�����0n,@�q�4����h^��W���������dx4��h׬�>�w4
�Y4��h��D�;�����v��g���z�:�kn�V�K��8�Q��1�F�GK�ih�]�r�ǀ�����U�&�w�� ������$�d��s�f�U�&�w�� ���׮��p�=��60�����V�ͫ �sj͍�d"$��r�3���7�~��ms@����9�1̟�7�}z���s@-����^��TM��L��	ɠ}z�h�k��]�}��`~�������\qm��޷-���M�k�p���u��Nb������@rۛ�.���]ge�����u`b�k��6��6��́�2��� M8�/Z����@�빠�s@��4ЖV57z��4^��T�z���f���+c�0� �D�rh�w4�\ܒ}�����K�Z8JS���J��0�
A.B��
H[ �aE���n����$��.�I8bQ�RI�m�hz٠n�X�ۋ�Lc�:�T�PEػ2�<���6�m��]ϐ��2v���'`��8��&$ƘI�����~���h�w4�\�>�Wc��EI�� �wj�b3��,��Հ}���Q6Ӹ@y2``'&��빠��}�� ��4*�j��
�hn�âb��u`����@���h�>fW1��X��X�ݫ�D��wW��� ��ua?�UQW��UQW��TU��TU�����
����*�*��*�҈����� �DH*
�A��`�DX*��H*�� B
��� �EX* @��Pb�D �@@��H*
� �A*V
�T��`�@H*X*B
�V
�
��� "�@X
�Q��* �� *���D`�E �D �@��F
�T`*A��B
�`�DB
�`�E@��
�H��*@ �D ��B
�E`�AV� R*�B
�DF
�D�� �A *A`�D��X*  *U��*���� �D@��
�TH
�H* �@T���@�� H* ��DB
�U��`*
�T�� `*R
�@����E*X*
�B
���E �EH*F� �AX�� �@Q��EA`�A*�T"�EE * �DH
�
�@��D �F�����E����D`�D *H*H
�B"���  *`�E *"�D *`*H*
�"*�� *� �H����B
� *"�*��F�
���D?���*��*�*��QUE_"�����*⊪*������H����"����*�*�Ъ���Ȫ���UQW���e5�E�� ]�� �s2}p�� �'��k�R � =����  t��'\���=8y�u1 �  �&�� yj�h@ZP(  P_GC�V�4���4Ц�eA&Z �h(5�45S`5� � kMP     6U
;a�  (րN/v����9��w����@;/�U��'�����r �`<�ꕤ�>�����vH�!����0��c趾����X|�����w�R��o����g�W��b��s{��]j���]T�������u��P��B�mO�{W�s諾k���=U�۫ڞ{���y<��xz=�s���,w���Ͻ�=��廯��׾��  #}�t=<����^=�|�}�}�t}���=��n�v}u�C����} �}�  m�2Vf�8��-��C}gBy����� ��pPR�f��Z��� �r� v�h(�{��=(;�H�(=�� =��4(�ҙ���CI� {r�%�� �� =;:h����馇G���h��N����:t��`�K�)J� iGЯN�耢�Э�m���:��{Ψj�PG��Ҕ^�z���Ӟ�y��jf�������`����NO��$�w�< #�w0�|}���������C�4��gOT4���t.�C k��i��}��`�� ��� 8�;M�o�w>A�}����n�=�y��;�Y��9 �z�L�����gl�o{���J�7�L�{>�v�G�[>A��C=��>�wx>�������9>����p ��M)��)H  '�T�H4 @��*j��T @��TSmT�@ i��I3T�!� D�6T�H���O����?α��g�5�Y����K��w_�AU�k/��] �"���
��_�P@U`
�*�z?ġ������'��Yə�� B�+�bh#\��.X�ۡ�l�XS۵�-L?ь@�jo�7NB�q�Zެ����S	�f�Р������秧Y��,��������v�1YW��UiRyvϻ����M��.�g739����K����E�V�
E[�w����ݼ�W-�a�v���>�uڣ����v}���D�h-}���]��xV��ﶕ�)��+�-��}�p�u}��w�Y]����.�>������o�uuG
.�or��m�����UEqR�}>��|���������\�
���c�;}��}��QNڬ��W����(���_mw�v�+h(��
�-�>���{�*�y���},���7n�����-���PP^����\��4�)�v~����!:�h�E�CA�:� �T���B��۬����ǅ+��#���S��7X��x�kyʗ�,���~ Bf�}�Կ8h֏������U*����W.��uv����)\|)_(ʬ�����}�}O{*��D>��h6��a�5�B%��\�q��77��$�O�?}�ڜ���l�C��k >�>��[���ϸ3{[Δ�����Ҿ���}uћx��k��{�����(�s�e��E��ͬ�HK&�����CĬ��-�P�S���k��эb�O�0���~tB��Ƅ��on����I��ː�_s�|mam�ﳭj��WyE*�
�q�=׽����>�\����|���+�B)a�B^���#P�|��FB���o>��ٙ�5�u�]�����
�Q�ﶴ�M[@�����{����;Y�Ӭ�����i����3��������o*���ϙ�g�M��0�]�WE��E+��뿅�2���?��U&U������x+���v��ޛ�3�E+{��ջ�.��}y���+e_}�fVWz�մ럏��Ə���0ѷp�o\���II��b>�Ϲ����v-ʽ���a�wM?�k8'y_;�+ݼ�>��������ksi�]ݐ�9��Lu/�~����3���o(V���wUw�}�qW��M}���]�t�Pm^�Ǯ��j���7��p�͑�I�:��������$�_���u&�4���#(����=��)�8kvog+/����5�ļuM�ܝ%N���4k��1����H;x��ԋ!H�c@@�np�I lcSW��\$C@;�8ư`l����d)�d6k����!LH�	\����CW�?�Ha����F�	BE�2J���@VB�vkz�����bE��#@�	�4����tu-0����)��Hƚ&�p���� A��Pܺ�|����
a�f�5_�N���|)p���k�߶��6�yG-��go5u+��\8kuaս_f|���
]���|;�}�-�>]߹���|���+c����<�nU.�
�����_ʺt�e]?��.�3���ܯ��7�Ϗ��]=�b�*�}ʵ[�F�����*��Ӭ�I�Ɩ���W�j�&�EOJ�;V7�{�'�����u�\���C��g)���O#f���x�|�M
~�j�ؕ8������LET���hX�]��'�ngX�����ԭ�xR�n�v���%����;_?��������������}����]��z�ҳ4��r��nŶ�;Q:�2���,F�y��.L���;��M�[��+`�W�֯*���^k�on��{J�����O�������6�Wk�v��xY>����/M�)����S.����Y���%�7��]l)�!L�xa�L+1)\�C"@ ���*�W%`�J�CO�&��T����Q���bTp
4Ʊ�E�q��4+l !LH��\X\�Ƒѹ$�=�I{q`���|_N��Vyؚ�,Il�c�O#>k�9�~���#r���(3?��򟯾i���Qɢ�'&��ߊh�0p�5�I����
J���Z_�Gό��'߯��c
�,���q��˔��#[�h٣W\%���8e����M�������g>�s��>w��>���Ӌ��ű�\�+��{��|,��y:i�38̽Ĳ��(J��(K0����X��\!L!HU�[!H�]�HJ��F��vZ�3�ɽn]�&��L4@ @�2�.�X�`E��~����B$�4L���7�K�־���q��/׆��7�0�f)��Q Ih�(��X�J�I���M�R	�5H�h� �F���[7����M�Y�~>c��}_�p�m�w��֌�m�5��}�Xt�dj�����BD��>M��n7� 0M;���@`bh�ō@m)čL&��q���S8O�A��6o��T�Z`hѳ���q�dpMÁ����$+\)����|�#Lm��a�4U>XW
�ۣ��o��������0��>k��ā%"B$@�(ĩ���5
*��b���*�"���p�c�.��N~�����6��7�z����\��������������>���YV��nw��Vѧ{�����
��h![���f�(F���%s�s�������sG⹼l��3HM�~־�ß��W� P1H0#X�?J�F׬~;3�Jwl�8~�����0���5���|ݽ7_f6�u#��O����|��Y@�K�ʶ-�_7�g��I#,!���kfؙNh%ɠ����8�~���H氎�Ƹ~A���8���8���6B�u�_���TQJً��<ֻ�uuuÊ��2�������O�*����}��v�� �f}���}�_;̪)c�����m���W
\��-����i[,��H����Y��۷���ܻһ;�o�S��=�+��}�ky�*�Kn�Yk]��ޝ�)Ry�Q�gr��x�EKd�w哯��U��K~I=���WG33�_f�����cJ�d�#M6^�2 CtK��ĉv|,n)��tSICEK�K�7�O K�Mzfu�=`$뱅p�Hs73R氥�A�I�t.7`�%�a.�q�Ї�����|�_��1.��@��?��RRsM�SJ���%t�J�jJ�lRq F0`A"b�C�B����3�;)O�q��M4౨�J~23t�*�"�4XFvK��k�g�w�{|$i�
B&!�o�����F���]HfAc4��.|�B�X����snIr`@�B�HJ2���*@�
²�M�����BE,
b����L$��� "���T�R4�����:�?~������]��!t�W��>Y��:�9�>�Wo����k厦�eK��}S�)r��W�ҧr�mO��xe-��c��kϾ���T+�N�������tP;1�f�V괔���v�����Y�U���n���/��}W{Q��O��Sற徝ŕ���)�N�5�Of�r�K	!��=#�=�����33s��j�}{|W���7�
�����߻�eQÖ��/��#���}ߺ_p3�����×�2�����5u�f}�l��f��^s&���!�)�H�eB%HY�7�!�y��7+�o�ќ���3LԺ5
B�Iv�'�����|J!�T!par�Oߍ�>c�Y��Y.�'6k>���~�BB�	��9d��䩭�e>�zs{B2ć���,�K4�l��s����;C�C���|�c���Ś����!?B����Щf�^��~S�s�C�ɺ^O��;�Xj�&��,�&�69�n�g�~�,�	�˾^$�J�jh������\�l�����h���0�!2#$� @�	D
0jP�h�"1c�ZiF-Hk0D�/�t3%���^џ��_'��]�����s8|�ʠ�Y���i�� \s<.��7�O0C��X���KWL���>_^�#���U����ۋ��an�K�4����_U�T���ޕ���O��Q�+�$�����>�ְ�M�6�~˻9$X\٭�Mo��D��,#�����=ٶf��&n�o[�%*�v�vٕ��f>��|2�+���%�k�U�]Z����'ϩU��}��5l��S�!�w�F���bB���JB@�I���	d�1$�Du*Ҍ(X�@���B@��Қd�cX�a0!��V52,V��5��3|5���ǜ�4������x����
t��ߵ���d�6��O��	f!�m#BbH�$F
�(�aL	 T B�@�+B8��2%h��f�ri(�қ>�q�M�3|ʹg9�ѳ����:���1��H����4n%��.kl�6K���o�����<��%��n1���.H蕗�1���h��4�*J0���!q%̈́�MP��~��>	T3C
�H�$�R�� ���E
���h�,� �D���������t�n��l��k�Eљ����l�#�$�}w��o�JsKJ�c�RA�Ϙ��fS,ME@����U(@�@�4�1�)�6S��0�G{2Є �d��c��$4|ZA��c1 ��HHńHD
02/Q�����[:fN�0�C9��Ŭ(.,�%�`CF$F�
�, B#��E+���h��	���.h�`�BA�&@��0�c�w i�R�Q4a��Ll3F�dǚ8~�,�>#	sD���~~��1�lɜ�?���4e}ך��_ ���˿��u����
S)��_�a���)���0H�D�F(T!Nk�9��>��|lꐪF��(b���/���sZ���?}��ݭ�5�wi�4��܊���Jwۯ�^�"�<v�E�UՉқn�E
n��u�O�S�e�^r������Yy������%�&[�\6��1"CMw)�d�Y2�F���$*A �!{qt�9��tֻE�x��0�X$�#VYx�&�1�tD�)��o���w{����r!�	$�a��0`�҆��(b荍$��3���t~��UUUUV��IjU��������UPUUUUUUUUUU�
�
���������������*���
��Z�����tUUPUUT�P 7nJ��uʰQ�k��#������.��
c]�_�8�Wg%��h�GC�L�dt����v�sc�37ۦ����8 �%u���:��'<��Xx8�jK0m�P��&ܷc�*��ӻ��`u	�v j�ڸ)m�ns�
�U�*�!k�ؗ�h��^Y_��T�+q�\Ke[/	�����!�+�Z����cj�*�7��U U�*�� ���`;*�4�  ѡ)����	�b�j�@��X������C�B0uU�P�r��L�KmUAVڪ���1� P��nSi�sR�Ұ檪�j��
�n�b������R�V�UmU*�UUU�[@U*�x<:Kf�U�������f��C��Z�@��K9����b��j��j�ڸs*�*�UUUUUUT������n���U UUj����	]���*�������	ejyZ�*��YZ����r�R�=��V���{.�QU[U*�J�T9iV�������j^عjWf��j���z��V @(c"��啥Xs�KU��J��Ի�ŬM�UUUT�J��tU[UGUQ�=�8)jU� �ڥZ��U �>ڪ���WU@UUUmUUP9�UU�U^����m��U�UT�UWUUU�'+h��J��uު�����UV*�WPb���
��UCV�(	Z�U}�C�_���J�ʵU@UUu]R���x$]����j��n��v���&������R��R�U@mUT�bv�r��UTuUWMڪ�( �F�j�����-�s��VR��5UUJ��|>~�$����@Ul�Uت�v�T󽝭��MU��Ku6�TU�
�����ձ[uԪ�.������-�v�.�k�j�g��U��z4
t�Dt���!ª �A�$�S�=*�SZ])ǯ��0Dæ{Fq��nɥ��UU��-2��\��P���	V��ьc�8�Ap8p��*�UP��wE�jU�*��"����^yvH��]�Y�L�O6���u�+��J�d�����=�㬴nlZs��b*��*�� ��+�=I�L���Q����P�v�sɳ����U:L�z*UX*��k�[V�����yeve[��j��l�Tp�Tt n�q�ԫUGN�[csU��n�W^�Šj�y'k���T��UUPUn�+3��m5<q��0�Z��b��J�F(���S��F�J�Uj��m��<s�����*�5UUT��J�a�$��2�JlUV�muUU@UU! UUUU@[@��mj�*��.�ҺF���Z��8-�Tt�UWl�UUP�c�nMW�y�[PN��vy��
��㦪���X
Z61�b� ��@ 
����uUm�T�T��!���n���'�N�%�UU�m@J�UP[UUUUUU@'�{SE��8�������U�tU[ ��h޳ث���&n'�	��U/�Їr�䇃�w�tq�	�M�`�<�k�F'����l�+V(�̜x-�c�K46*��hY�ԔB����%nڂ�V���mƶ8���明��5���U)@��s��u�mWM6y�,g�lj��-�m�n�/R�S��UvtK�5*�oU�k+���,��'�A�M��'c���[��˄ϳR�Wm�#AK��ڪ�S*����v�۬v��<�@�>W�������UT�mU��UU���A����k�f݌�Y����D�qv%��� �U怨8����UZ�����r��]�V,DiB��ڪ���UU�H�*��ڨ���U�UUUUUUUb����\ƪ�����[!�ɬ	�aM0 �����U�e��j�gj�tT�WUWT�*�UUUUK��Q9v6�������O�a�"��e^��R�lUG�(�˷[+�Lv�UUJ����*����Wf]�� �iJ�'si��$ΆFH:n�냊��Z����d�;��}5Uq��촤�UT�p��E�l�!�%����U^�c��F����*�ܲ�Xҵ+9�ueU�� ���*K��&��l]6�(BS"��6��WPv�:��#�CXڎh{v����.fڨ
��RM�@��W"\�R�W6[n�P6j�DH#V\�V"؆��w&}]0t��ny�˲�r�Z�8���L#sķ,-�x�rR#�0U
-���f24��q�T�N��q+���r���Z�IkP=��up�PֱIL౗6�\�6AU�*�8���5ئx�F�J��S��n�sOJ욹<E���U�<�J����I�UUUU��A�UT9Vj��U�-���uUU*ԫmmU�T��NX����@ ŀ��4���X�J�+UUUUV5�ԫ���|<|�J�UUTon�)j ������AUUUUV��j��D��6���������l9��ꫳ؆�+cj�
�UUU}U�UV�UUUUUP媪UUUUUUAv�pf(ޤ*Wk�^{�
�X«��ޮ���
��
��Vص[b ����5c:��Z�����55F4�mZJR��@b�*��TUUm*�UUUU�UUUUUUUUUP�UR�R����V��+Z�v�6�uT�(皪8ت�*�P(�%V��5��W[�)� UJ�R��P��a���U�U��ꫠ+��������UU����������UUY��Ub��J]�Ԧg�A]�ꮕzکV�eU�%ƶ��`b�UAM�����	UUU(*���������� �T��h����W�W�}l�֝����ms��K��681���ڤ��z�̣TqJ��Tm�͕��8V۩��.X���!W;eXA��܎�v�Ę���٘�Tr=4�q�9��jIWj��)u	QD0���̺�4�qf��[,2�Q)�	�mf���<H�`v{V�l�9�l"�)e��h5·�.q\c����6⪧��E�J���w%�L�9�c��2��]@uWI�sZ	�v�mY7$��Ej��;��nM�,)�Z�c���b۶<��j�ofV��/�'� �mW�_UW�$�U�N8H�r���b���gk��nQ�R��p]UV�CUU I{s�5̻p�J�*��	6�ԵUUUUU�[T5Uj���V���k�Z����Um�v�n,9^V�������� 傐j�(�A��)	��UUPUUUU/*��j��6ayB��i��wW����UUڻ*����(M�ݠݐh�]-Tl�uS@��0�em�k\/W*�TUUPlU���	:��B꧜=���UUT��\͹�q����ڪU�6U�*����$�n�U�UU�4*�
�;�����UP秮�U�]���.��j��iV���u������5�	�[*��UUUUUUR�UUV� X���������[���;�8XB	����������*�����%��V�
��v㉠��j��ƙ�V�V�y-�����������U�d.Ғ���b�Uo&���U.��bF�Z�� *��W�����j�*X튪vH��)d���9�Z�UR�}W��UX�m��PTVeVQ����{��rNI��t2������V�RUR�J�K&�ݙ��3P�M���X���]BQ�A�*�%�T
�� ��ݒ�_����㚅��ٙEUU[T%0��]����j�6��[zc��mƚ�*��JY�'ϱ�2��][4����l^�A(��q���q��مr+��mX�_���b��Z��m��U5mƁUUx"��� 'k�2����ǭ6�,UAGl邦�UUSj�P׌�XV��pёCmn�í��P0�����k�m�ԭuU]A�C�5�'d��UL�	K�yF�8��;��gex&�W����*vt�<�Ei	��<UUU��[#���=��Ңp��$̝��3f��[	������	�13�E�a�l$d���Rʙz*8���vn��g�q6T��2�F�K@���BƎ���Ѭ3e��a�D��I%( �Wb��F2 x�X����d݋�`/����9�Zdi��exA�Ȯ�+�V�[V� UKFۇe��j�઀�V�����v���ʳ�U���}@@UU@�0URګUUU���J�ԫZ��=���3>�:��F�$�UmPV��u�WT�5]UFP	�z�,�.��j��l�R�5@UUUed7a���UZ�hT��1�lT�J�ڪ�U�]���V��EZ�b���X�4�h��m�j��UY�UUO+M��*U�����;UT���^`*��K�UVX$��0���V@s*�UUT�UU*�T����UV��}�l}@UU@x�Ǡ�UF���z<Mʻ^��U�
�w���9�����w�}U ds�1"u+9�j� ��ݝ����ZN;L��֝�����o����a���؝u;�6KЪ����oM�ƉwU.69:X�b܋�q6��]T������W��*���5�-RD�UUUU��J;E ���IP5[m��Uz�*��������X��U �cll�Z`*������*�m��3I#�q
�6]�ɔ.L�ا�-��f:�v��Pu�݊f��r�	�s٥����jĐ��ڐ���!.1��UmB<������sp�MsI-Vay����2!sv8�UK��ԧ�emU*��<����^A��ڪ��
��Z��5UR��UUմQUuUUPUSiP�����:��Ņ�j������� *�mM
�`�A4*5�"	�T�*��B H�F+�l���b�J'�lqG��5 %0 ���C�i? �D�J�`(�*�U( hA� M�M� �$�+�S�b�"0�l@�H"�:@�BhAڴGI�Hb+�~U�X�AN"~ �� �`0�	�V*�iW���~t�| FpȐ���	�������O�ʉ�`�O������H��b=P�Pv�V$A������b?��"�L@P�� !�;]��:��"-U��� ��~1T�=Q�v�"�Uҡ�#�C�D:�@�X�B(ā"�H!�t(��bQ��b�~Et�����E�k�Q�
Eҏ�!B@IFEN�#	�0 �	h�*TC�*0�>P
�8���C��@O��RB4@��!$a�?�LEB���F��Oʇ@W��B$IHR@$	@1]��С(0A ���
u�i���-�BVXD�BXB%cB�,�))%[e�YI�$	XT�0���V��%YH�lG�%��F!�Z� ��bE�* h��⦄U:!�uE��)� �� jT&�����T_�>?� DF(%���b)Q��$	E�c*6�Z�`U!j [Ӊ:K;�,���U[j�Қ���*XN��ô�}���eF���Z��k��5"ktx	�7n��&��:�c�5��Z:�C�\���*�D.�8���Ā�WUU\;�X���70�Y����+X�U:y�ړV�,h��F�ŕ�F�=mty#`�d�b�X`L�ha�g���l̵��ꡐ�F�K��]!�a�8�eNv_au�d\%���ᨱ��	sf�bX��,� ��7����p�n.<m �lU7�WuҊ�\���Ep<�c7�nN|&�[�V�#��n�Zt=K��[�\u8Bl��Pє�)ZJ!*KB�'��������`3HV�+�[�&pf\��6�����k� �w0QsZnkln_v� ̒R�Zy�����·�k9���cI�j(���E�q ��E��݆զ�-Q�LE�j�GOr�s�4N�uڌ���e#������5ƍ>�����m�◙�3��-�k3v����;e�@���o`h	U�1�z)U�l�
X:ͣf�@U^u��3�,4p��pXy(�lsCۖ{B���#Q�n�Aq��n�<��t�Rp:�5sm��y��kEۢ�p�y�-p3"N:���b�2'l����+�f:۝�P#H�@��:�z���q��v�����΋$�#��T���۲�n݁�a����&�X3�궝J��gn6�9�Lv�TxU��h��29�N1�ؔ���BQA��V��u��6�0b�g��SX�V(�M���[�.���Q	�T.>��s��ZW[6b��0R-e�J���Ӈr�ƦV�`�J%3�)�)��cc5$xa6�vy[0!��cZ���F�9�r���"�aI�2�r��͑ �� �]����=`�΅Pwv4n�1�j0aE��mFE��\Ppr�\�X��@s��$���ԻZ|й��M]mlp[5��l�]�H�H�˦(�ֹUc��̲w���;���w.�"��h�p@�"ȯ����E���]��t!�QM(������f\�:fkR�f�����v�@�ٙ�&� ���e3���+��n�J;\Ԗ;�f����a%�]ZSA�L�Wkf�����Z�q��\.䭮NӞw;&IN����U8w[Jw[�L����X\iK�����p]e���t]�p�g�3;�m
ؼ5��Wu�K��
�f^fs6m����k1qb�<h�I�=���Iv%�LLś7�}�${�����y���kN�,o-c Q��-b�`X�������iV��+�h�_]����ذ���~ק���^�������uk��Lm`���D���;6e`u� �4D�j�ue7�]��	��}6e`u� �֢�>R�����Ӣ���l�>�2�	��n�Q`N#�� �nD;T����LV� ���;0�̬��s��n�]z�\sl�	�
�;;���rg�m���0n��\�\X�
-���[��+R�9� �5�N��+ �{ޑ�[��К]5k[���?�	�8�,��!! ΪD"`hA�G�*��W*�g�X��X���2��bJ�ݳ �l��&�ŀn�Q`k� T숶Yun�M:����$�� �֢�$��6^�����ծ;��0��n�Q`k��/ ��,���Uz��-]�<خa3��E�v�f��#`뇝�l�&��oc���j�2�K�j��Y�������`)��	/b�7u�X�RQKCun��n�JـuM��E6^��E�I��r����~�!ڤ�tP�:n�Y�'���ܓ��j��~G�#AB�@"I$���`�� �U�fI���5we�n�Et;i�e:T�w�wu��	5� �vK�"�/ ޒ�W�un諥ui���$���/ �l���E�IVIo�n��oiug1�Y��f�n�C�>-�pG�vnz+iU��ەsA�3H��'�|�߿o ��^�֢�&� N�*���&�]�n��%竜�q"H�k ���6^����*uw�vR�
����Z�&��Uq-[�^���Q����VU��v�`u� �왹'o��7'G��`;D�uA�n}���RZ����WE7M�l�:�%�vK�;��n�`n��&�x+nj�'r�b�X,j�r�[sݷ����/��t�h+9�/=N��v�jY����z��k ����UU�^�� ��^���L��ҧn����Z�&��6^d��%8���wE*WV�n�7\0����*���z�	#��d��Z(v"��@�ف�W)m�z�-�� ��-`u� &˕i���&�]�n��%��q�n�`Se�R��ڵbW5i�-X]KT�ks-#3`M���e�Q�:���X�7f�2����C��h6S�6��k/R��2�[�*ᶮCM���__Bӈ%	��k�ݣn��]6�/	æ\M rq:�<�P�Zs��!ڹC���W0"�v�e��v�a1u�v+��m�©M(�v4̤ƞs�,�5���A��f�rl��*�b��t�\��Iѝ%�<�R��,�8^RظZ�U[���C6k��eՊ����[��ʆ�;��0Wn��?5�M��l�.�xTh�KT˫*��v��&�~�VW.�[�^�7׀n�gx��)&����WE7M�l�:�%�vK�7uư	��w�*!Z��:(m�ڷx�)z�޼H��7\0��x_wT�mYuc�NӶ��q�n�`]��	ۑ`�+�����6S��⺷$�%�I��n�7�:⭻<�hnD�%��\\�c�1xYq�6j?����/ ���ʮU|�l~k �����P청��[�`]�y�s���$#��%��B2�� 8i�x	e-�HH��MMt��a�&�@�B�.~W���>�v�V�c�X�p��r�������n�	ۑ`�q�n�`]�x�⺔;��0�l��9U�6g��=#�}�ذ	��j��@���g-�N�X�p�>��X�^�g�������aI��wl��YB����Z��̪ɥ��1��Yw�E�3I���1�[����wm�ݽ� ����7\0���.մݲ�n�7m`�� ����	��}�ذ��%�;j���J�ҷX��w�M�vnlb�HB"|���t�w7��}�2�	S\��v�j�WV4�w�M���ŀNɕ�N��x�1��P첝1�[�`v�,vL�v�;�&�݁St]�t�]"�iA���V��ef�j/`��ձ��2�M��ѕ-���T�um�k ��+ ����	��}�ذ�j�]�w�vR���v�;�s�ďH�`۞X�X���	j�vr�ěw�vk��ob�7�e`�����iaJ˕t1�I�f�ob�6l��'oc��ʥ\�V�W
�8�܆���Eڱ��E�J����2�r�����=���ŀ|���1���v��]i���	OiЋ�e�lV�h�k��&�d�2Y���Q�Uj�t��V��=�<� ٮݽ� ٳ+ �5�|VX좕Ս6��5� ���`6e`����&7V�N��:��i�0�{�fV;{�5� 7dat��۵N�Vݶ��2���f�`Kذ�5p.��v�S۬f�k ٮ;�v�I�~���4'�B"	�Z ��*H*�a �b;�u����~�0��%e��ц0�J���.sل���k�K��i��l\ob�1s�ܼ����9�YbMe]	����p�B\Bb��s��
k�q�Վ1tn��'T��BL�J��&I�5In�W\qŸ�/NP�Yrf=e��P�qp�+\�[��!,tsy=���Fزb��񌵢��mS��&fI��JU�m=���y����䗧v�Mǉ]�5�
�^�7��C������]��^5ٛ�rN����3�+j�vr�V]�]�G� �^ŀlٕ�l�-`K,)R�Et�vـ}/b�6l��6k����N��Eڱ���*�m`6e`5�X�p�>��`w��m&�Z�*���6k����}/b��M�X��G�ʷewVSM��6k���� ٳ+ ٮZ�>�W��M�;X3�b2=�OMu�v��{hm�[��Nl�l��̀�Cm�Xh�ѺTξ[}����6e`5�_�\�|�z?���]3c4��-�=������N�pN�'҄l��l�j��5��?Z�>��}/b�>ڎ������T����r�ٮ��,{0UK�Z�]�cUe۵�vk���� ��f�k �X����O�.�N�0��Xդp�6k��	��z�KuW���M�wN�n�4�y�T��;!�S���a�f�v����l���b��cm0-�Un��m�� ٮZ�&���� +��]�6骱��wn����=#�w�<�=���z����w�wrƹ�ō��<���o�}/bõ����]w�t;|�
�$����{�ɮm�~|���������y[�&���ȱ!��n����o��}��������������~�K��#%��d{�$ǿ=��.}�_ˆUѺ.s�-����0Y�.��j�>�.�>e�ىi�
�G��~�'���T���:2�λ����}��J�}�����-����Q���?��w��+�B�,�].Qw�/�H����e}z�ؒ����5Ԍ��"`H2�����S0�Xe!C�
~�����o�7nè,
F�H*��H��"��Q#@#L���4m5��o�߷��Y;����$.�!V%e%�cM�?o�s0��˽��L��B,Ա�Mj���]:��$H��SLcJ��EbnS 0����e�6��
���r��X�gh�t}W�:��B�8J�I��d�+!� �f��	G��B��9����֝���K���jo.�f�vl:����v�a��t�d�����&:�Ǜf���?�,cow�'~�-��fl �������&既 i �bD����+��Dv#���1HE�  �����#�T6�G�1A�C@+A8(�
�U�(�Up������x�k ٳ��N��:��[�`Kذ�%�5�X���/I�0}�0�t������ݶ��%�k��	��N�ŀv~�G��U&��p�J�õ�=�l"dѠ�W�c��Ѯj�X�Z+6`R��;�$�-`u� �����U|��}��<�ʽtz�;V�ƪ˷k ����X]��	5�X�R��|tӻl�'ob�"엀I�Z�&� N����cm2��V;k ��^w�k�w$��k�ra��(� A��4!h��D,j�X+mD�V�9U�/�� Wf��cwb�n��&�k ��ʮW=3��{ny`�������XX�ٖ��a%����V�K���6�q�3r�	��bz�(�
W�Y�ۮ��M��7�p�'ob�"엀I�Z�6l��!:�T��AnـN�ŀE�/ $؞7\0�#N�մS��۶�d� �bx�p�'ob�>�t������%v� �b��&�;{d�*���Rӵj�j���`u� �s�������{ٹ'{�n��? |1�a���GM�u��U Ԅ�,a������l^��ĂC�v;9�O]��8:�Ya�ĕ.�5��ˌF+@Ĩhw[\1�.+Ml��ְ�skd����)q�K�;4��N���1���l�/��2�>��O_����\h��ԗ��.q�f�"���|F7'k�:�uf�J�Glȓ,Z�ӄ�z�MԜ��5����kXK��ggO���F��d�@�ar�j�c4t�כ���P�뭒k[��P6���*`�È&�vS��y`vK�$ز�	��ڈ��v�)7J�v�d�M�+ ����X]��۱U���M�+ ����X�Ȱ�z��L�Vwg�� ��~�^۞X���&ŕ�lٍ�C��0��i�0���r�o���{��+ ����[��Y�CA�n4��I5fbj�ű2�
�1�+�qJ���)M��/1�]ZM��7�� �E��vk��U�-�� �?:I�����*ݳ �E��\����Uo*��� �����I���;XN�D��nƞ[w�ۀN܋ �ɕ�I"��>�-,*[j�hi;l��qz�޼o���I"���qo�x�<�^G�X�I7WM�w�od��=^������G� ��^��]����=�e�J�ͱ���%��<�m������kaȅJP�
XV1��By�͛U���n��߿,��\0�%���}�z���L�����;�� ���G��׀M���	$YX�K�ac�ZaIҴ�]���Xmr����iXB(TlBFD˓�Pj��ʨ�)Kd��
Bb/�\��~���=<�`썊������w��)��Հ{����;5���R��xey��:W|v7J�v�`H��UW7�<|��׀lٕ�~�r�v}�DE�A�ĎL���yt4v��O���8ձ��ˮvA���7��>��i�&4��Ӯ����.�x͙^�W>A�{�+ �/R�|����v����.�y����ʻ=�߲�߿~YX�p�Us�^�#֬V锓utڷx��V$�+r��%=��}��
�a.�M�-��V�ܪ�/{�_V=�.ɛ����Q��$#U-B�gQ��9������j�������;��bI-�����9�9�d������[o{٭�v��Ox߭��VVg���G8��-%�P��Sj�.�C�͵&�t���v!��$�]�Vҥծ��Ӷn�����Il��}�II�{�ϔ����� |��U�V���پ[m��w�9�
'�֯����ɻm������/������۠�������ޚ�7m���}���O�CZ��=�/�������@>~�Ԅ�5[��v��;$����o��u~�� }�～�m�U?�u���9������?���4d�bwm�|�Q^�x�K�UUW��s��w�_�~Q�$�܇�$��9�AG
*�$PȒ����fe��f\����f���1J�S��Ws�80l�L�@�M��"��cu�&�s�{ea5��1��+�@D�)*�ٜ�j���Y��pM`�LB����R�X!,f��\�w:�k��[�gi�61��;{u�^4�ێ!ԙ�3Vb��;iF��r�%T�����K\'!W�+`{O��\c�"�R뭞î��n�]�ia�.��vQ�I'OzE��ѡ6e�C.�\��ceڼ5x�'FwSY��|\{G:�T��	�YB�$����m4�p� ���?�~�$���1$����s�U��K���I%]ؽv�m:\��6}�II�g������ߧ9m���]n�ow}��T���۫��3��t� ��;}�����d�����;}����K��}����(��)��>[���4;��"?����m�����9m����7m�*�E��{���{�Z�I��g]�����9�m��������~�崿~�]��������e�CG�vq�]�MRU����<c�9�u��V+v���ӧwG+2��w�ct�E۾�$�<�I%?~�������NNz�u�޾�׽R��˲�j���ĒSw!���s��F"PrfSk.0� �`P�I�M`�bi0L�3I�4 ��(~��?s^�ݶ�g{��-��}�����NEC��>�:�,r]�_} ��v� ��}��$�����%� ��y��~�O 0Ci����"g��������ɻm����s��"Nq;���� �߾:�61-t�9s��%6<�I{�\��I���$�G��I?�|��������n�f[j��&���]	Ut�.V�ė$p�n]B�@����;�2��2��T��>I%�3��$�5��I)}���r��]�<�I%!=�C#�A��O�-����>{���m��>�����w��7m��}��s«���;ݪ�Mʹa�w�_���~�[&�v#C����@F��HȚ�2(\Pq��U�6 ��y��{Ӝ�����kr�yӻ3�V\�Y5����g9m������I%�3��$���X��+�Uw����A��&�cq�_ �~�����~���$�^�y��IMs�$��/�۝q�Ұ�c�b*8ԚZ��3"�,A,͵��)e���9$�a�x�L1�Ӥ��;Ԓ^��bI%;#�䒚�#���~���} ��g���!��j�1$������\������Ē^�<}������I}�����k������$���Jn�>�~����\��m~��f$��Oߟ�$��ԧ�;�T�t�%�s�\���x��==��$������Lρ|~�Q�� �$KAP��,bD$#	$@�_.��P{�~��ݶ�w���Rd�Me.��-�>�$��)�I/ܮU~������u$�z�e,I%7r|�RUŔݤ]�nSy��u��<��A>��M�lr�u��5g����I!�x��I��Bi�%����$�ۙKIM܇�����I��o ������y��e���~~�Y��r��������H��SĒJM��{$�$T��FX�U���·����9�m���5�| �f_{��9m��{�x z����a���˵��?��?ʀ�?��������k������wm�@?Ӝ��o����������@tBkMsF�m���w\�� ���������������Nr�g~��n�n���"�"�s2%��?~e�e���B�]�c2�3:P��}�CY���������I�͜���l�hR0���B���mv�TR�tw/��v�y��I��\|������p���wL����(Fl��Z+WX���+��v�ϻ����9�_I���Cy�ѳ�0U�F!9ɭ��p#JKa�៮�F��&Nd��$�	B~ĸ���0�#Q�NO�A�V��r&h C������W� ���N[F�3ΞI'�>2y�~��Um��U@U@mR��C�v�8���a0X)v���S���\��u�f��l�۶�C��Yg<Jc�L�[�5
C��2A�%������U	�l�Τs��	Z��U;>�� �,�Au����]���28�ϛU%^v� )��Q�3]Nl �X�Ѩl,9�m��R��-���с�T=����V��Pu�nW�������#"��]�ٺlr�;�K/9�;e�{C���N��"�B���yk�C�@�IJ��\�-�V]��V ����,6�JV����Y�C�l�-���2i킍�\n�G3��|�j�l�n�A(����]u��9�=�@�q��Ť�e ���\&HY�L�R�$���,h�S��F0D�b��(�]E-�`ץ��:و/�U������H؛k\,m�p91҉Dgd9��N�H�#�Ml4p���+[����������-�\,��N԰v^��v	5tZx��<Z������`�p��"J�횴O��]b�����H�Ѫ:	�b��U���R�*d����ۆ�ְ��mN��U-�F���#gkf4�f�zܱmR�8v���糭@N�))��Z�G�Mf!J�Z�]E-�1a�ۮs�1��)J�`m�g�Mکk���5 X[m�Y�P3�)ob�#,��j� Bm"��SVx�]\) �r n)��6&ZLp#��v���2�6�m{��d�h��!Z�N�;Dݶ\v���V���Ϡ�� @�朗�h�h�4�lpuT������,7Yѭ��V6]�lI�ځɜ퀘�Q9�㤄�g=�lQ2�k�]��EN��ѩ�E
V��*i[	����L�	��x�n	����n��v�t�rgs��aئ)L��eAr�N�BJNuL��,�հ�*cr��J��5m����!LZ�.�(�����vѢ�ϰ��70 �����j��"-�Ұ�76�Jn#�6��x�+P�K�m��텗�Y�tr�`��R���Q"�?(��C�(��O"���?�E?*!U~T?�PD�r�#�>?��o�f��BYKY�B�iK=�C������t�:mD�'��M�=\-t
�b�HJv��v[Y�kv�֦9,�Ok`�p��!�p�Ǩ���Z9�2T�֎�(�*�����5ݻx�VZmIu�f�LcH<W'6��p!^QvJ1���Е�T�Z:��� �L�K��M��"�p�a���6&�4�m�yt�,�M[��,�S5���[ਧ�oF���~%<3;!]b�6[�E�m�j\������X�I�,�k��1�ww3�<��!�Fڶ�K߯�RĒRnC�H�2��ʮz������v;��Wq�gHCĒRnCￜ��U�6��߲�$�_����Gߟ����$�����gg��B���$��짉$����ܪ�6�z�e,I����}� ����5��k6�6�xȆg��������v�{����-�U�߻�� ��񷭪�Ch�UϾ�Sne,I%�UW���z�G���$��������	���`�Jlf�
��[L�[�Y�Mcg�V-n�m7�;�n����ln#���߾��@/߷�x����?��C�m��l��������iQ��O�-����>=4��B A$B#(J@+B��� �ҡ%`�#%���lw���w�|��߿y����rEN��<-
:`.��6�������	�2�%�s����<��$�G��I%]�ɴc�ЛaϾ���#߷}���<��$���ė�r�r���?{���I{�g�n]�GXm%6�������@;�NW�{�|�K����䒛s)bI,��f�l��uc��`x��Ŷ�FE��S�WNC�U��J1#=�t����.��m6�RKc�#G�l�mȿs��~��'�o~{�<�����3X)6��3����yꪮRG���M��N���W$����%��Ch�Qϖ��~�����n���
��� C5���7V�^&�tU�Z�vR���\��T�w~���w��7$�������r��<0:�K�����ˤ�V��X�]0'*����6_�M�y`�ذ�UG?��v���6
�'�pV��Gd�g����=�9��5�d��o�O(Ynf���-ݺ��O^6�,{{�\�W�'������7J�VէJ�j��/b�r���&���'�����y�r����0v��J�P�X۞X͙X{��%վ���<�]���+�:V�k�+�U��UW�����5O߯ �{۹?��H$�"�(���1H, ��*Ίq�g�~������n�]�v���E�n��d��r�����~�ߗ@���`$��>�E��,j�`«ƀH!���0\�8��,{A][�V��z���x6� ��a.���������ŀl�+��|���׀M���W����@�n��7��g�s��\��߿~��5~���6\�=\�$uz���ߩ;WI��+��	�{+ �M�����S��,m�,m� HV餇n��u��s�������,��������� ��=M�o�զ��v� �0ܮW?s��3ߗ@��߲��d��\��,
���lҀB�ԕ���̮�e�u�\��i���E�B��4�K��L^�u�!|U)�Fmc��2@���j��b6aI�m]FT�5�`u���؁m�v.��c�������&3݅��%L�2ؐm,�n�iM��,K�ہ�?~�z�&���10�Y1��l�L]�I�]�1�lb���s(2�.V��6]B�@aH�	�	aL5�`!�1�3����wAk�,INmJ�o.�]�8�4�%h#W`�v��75�@Nͦr�"��t�;��)��J��(v_�,d�X˲]{�UϐOy��"�y��+���ӥm6�	6e`.�x��w��g���$vy��:���Se��v�`[�^&�a��*�ݹ兽�{������|�d�te*��{9+���x�7ny`I���W*�v�޼��+��-q݈���f��ŀ9\�?W9\�߿~�tS���$��%$��&Qhau)��KJ��^��׋�;9���[m�c5���$�zoS��&k��������/ �8{�U\���, �ׯ�b�CCV�I7X˲^g9O�D�"����M�;�����{��t��;�������f^gJ�'��~����Us�Ľ�{+ ��z�Կ��a�Y�nd<������{|�����d�W*�����M�y�|Wm1P���V�$�XWd�K�`�Ȱ�Z�[�m��e;I�"�卍Ce��-҄e+�͚�B��q��M]�t_>
�ʱ��B��|��� ��X{r/r��_ ������^�.�-ҡn�	.E���r��]�_�,��߲�O�|�9��������K���-�}��ܓ��vnQ@b��	$i���#�E�;@ �9��=��{��]�9z_�,�\�����{��rC��}�[���Ir,s��U-�<��|_�b�CCV�I7X˲^�UU{��_�~��$�+ �\�{\��:|T�4�[�֮V��q�΃�,R]�]	cpdՎ�����7I�X�j�۷�_��	��I&W�s����,k�=c��wWM+uE���ឪ�URG��e`�<�'{����!��9����������I�FKv���߲���a�UUR^��� ����>~���lL)�+<{������'���ܓ����Ɉi����{ٵ�OD�^������P���	/b�$�M�XSe���z�.�ꃥ�X:6�G611�'V��w<�@r�p�je�1�o�$��I��!��mt߼��2����r�� ��y`^���vz�Vun� ��+=UIl��}��{��]�;ߵٿ�A?�s'���_���lV����׀Ir,=\�%�G� ���`}���&�bt����{��^����׀I0���Խ�:wu`�uCm`�%��r���x�^��K�`�U�[��`ؿJm�*KcYv(X��0a���C��Tq��9M�ٸ.h�M1feѨ�Y5t��f*5���k�8ܷcWmq��+GRE��v6x�=7���ړ�OH��g�-;bN�V����@8�<\7��]vw0�2��Qn+nxybौX��e���`�-!��l�a�6gjFU��i��=�-h��aH�m�@ �QjX�]��9��<�=�l0%&9�F��Dpu5�B�p��[R��&��B�`[�m��w�{��������~���l�K�z��_ �}��;�?&�U�V[�
ݳ �/=\�RG�~��"�z�	#�*����v/]]�SM:(B�x�~��5vK��+����?��x��R�\wV����%�}�f����$������D_�J�߳��j�K���i4��j��$����[���z��uvK�6k��p�ɓf����;.�ƘP!6q��Y����zڬ��*�¶�^y���v��> ���%Ȱ���\��{�~0���7I��N���o ��Y*�]䌤7�BD��SSO�CH!��)� h�$"��F,$#M2�
�2F$  ,���i�kA�2
Ȅ! $)
�BB�"R$"�"�XC
X@R(�@��N��%W�s�φ��׀O��0����r�6�s�n�mYWL�T6��}��$�~�9���*��?~x�����7�c�|N�b��Wc�x�� ;�%Ȱ=�����޾[���Ђ�WF�G:�m�� �+�^����j�z�	#���x���(̆c���QT��2�e,X��R�6�F�Cd�kJ��t�>��w��i�E+��޿y`]��	#��\�W��y��/
�Z㺴�e�m`]��	#� w�<K�g��+����U���~���lV|n�߿?� w�����ϊB� C0���a�Gz��wZw�~���K�p��2Lɋ������n�YIbo{���G��E5�C�3C�6JL�֎ol�u�����3h��0��C��$���ߟ�o
��J����~�F}����s�d�{�f��Mn0$`@�xB�ˍ�:q�����;\�q�x���$������!p-�`�,�B��B�_~w�߯�'���#2�eĊ����q�$!2���M�7�z�5�.ݘ��K�gn�l�"!����C��ɕ��
��ֱP�.�+	�fٽ��0$�Ò�80�Ɵ���� `�0vi��bF#�����������2�ҊD�h�$Q6��N�� �]`'D� ~z)�z��Q��Tj!� ��A��\Q���w���rO��{7$�'�w�D������\��}�{��,��^$p���St��-Ӻ.۶�	.E�{����z����� �i���2����H�h���rή��ؘuԃqtB2���k����a��uCm|��������� ;�����t�~�>�޶����|��n��
��	#� w�<K�`]���Uďm��t�]��uc�[�`vy�G?UUU~�r�T���?~��݉إ���4Ӣ��m�{�K��x�:�z�	&�7'�&��L��o�ܓ�},��uiP�i� �we��W����vy�G�+�����W�l��v���r��g�5���m�]�k�Є�r�ɓV����*Ѻ�]��m����`���	#��U�������<�
�cI��0��x�� �we�G�+�O)�n�uE�wEݶ��y��>]�x{�I{�~0�<��H+��S-�ف�Wog� ���`���	#�6LL|N�b�IաۼH�~�U���Ϡ~���0�v^���wp��B�WJ��Vʻ�aM\�S]�F�L�h:�s�n�1�.�Q�L2�v6ف�B���i�M(n�;*�;��b��l.�+(�Z܏C�VL�jͣ�Ή�	Վ[F#]���UM%kŰ0�vوњ`ى1WE��5̘�f9�s�K�p3�d�p�(]D˵��L�M4TЫ���	q��v����Aq����76�Rib�F���I=;�D�TڐD]K���.RU�1���u`��H���"���c@v����<����E��Э� ����	#�ջ/ �8`v'b�WwT�N�*ݷ�I3�ʤ�Rz�O?��y��@��:v��9������m��������\�]����~����&�җV;-����$��c� }$x����qK�׀uQR��IX4Ҷ	&� �H�r����x����c�x�>���z������#t��+mIU]\LA2Bȃcn��X�h6Pab��5F,�%;��շ��~0[��	���*�_ ;�y���t��V*e���0_}������JB����V�	`. q�_"��y���I�M�ݘ����j�'V�n�	�� >�<W+�T/O?Rz�	5�n�+���V:�f< �����{�צ���RuP���;�N�뫻�i�Ei��M���x��I�ڍ]AYl�s��{v|a�y��	F�ǚґ�ٚ6p��T��S{�N�3X�y�:b�f�����c� }$~�9Uϐzy��=.RT����_�I��&� �H�	�� ջ/=\�U$uQR��IX4Ҷ	&� ��M�N���p�W��D�ʀ�����>���ܒrM�MҷT[�t]ڶ�	�"�5n��&�r�T�}�<#�𮓶��L�T6��v^�r�����}�<k�ǖߧ����]p7crW*K-�(x�\�e8s3
��u�ֺV-x��)�ut6��ٕ��ǀoob�I'����{�����s-�h]-� w�{��$M���y�M�X{B�Ww�'n�*�o ٮ�w��\���߲�vy�ʊ���q݈i�`z�\K��<z{+ ;ݏUS��Ws�0	��R�ƭ2��|m�6e`�r����	��`ݑ��_� �1�ʔ����i��+<3���<-�nӶ�9Z��L� �����'��A�+v���_ n�<f�`{#�\��|�z{+ 4�~��6p�˥wj��6k�{�\�~����	?~x�{�V w�??�;��wN��}����V�h���< ���lٕ�� ٮݘ��C��'WM6�{��W.z{��{� ٮ�\���r��Oߞ���~T�ݕe�(t
۬ �dx�UW9S�<|��<f̬�U�Ê��\9Ċ��lb�$0
��I{��|n�#���!B5�WZ�pe�E����c֭Z�;�šhҖ���F�#XRِ؟gh��u�p�Y������n�4 Lg�
l�&^ƌ��V�f��>Oc�d�ķi���Iv��;U��� �+�!�Q��.A��4#0 �X�8D�e�ZWLT����%D\s@i*Muq+4��L)]��:�Z�t3l�l�M^Zqʹ��^I9�O���i��Qֳ�:��y���ب9�1+�c(	
](+u��};��k�@9�e�W�{��� ;�&̬ �dx$EC��v*��0�����G�=�����$��URF��_��jӵW����{��X���	5� ;� V�֊�n��+`�����%�<�z?�dx�W*�s��{�k !=��l�v��v�o �\0���	6e`wc�:����Ywm��XK����Ge��:�ϜAj���MC�έ�D=�2��]�m��C-�$��g��	6e`wc��r�_���߼����+���%ц����>��ٺ����;W{����$���G��W=/�ʕ;���E�[u�'��fV���IuOz�	���5Т����Ewm�~�)OO}XT�� ٳ+�ĶO< ��ʇj�v]Zv� �l��~�OO}_ l�x͙X�J��L����-��9k5�8�M���\�<:�uq��)3C�ӟ7�x�7WY�d� ����< ��x�2���x[[Z+�mP�J�+�u�ݏ=\��z{+ ���l��URA����n�.�m���nI����ϓd���BKF�B��X�,B	Xg+��\�j����X�o��awI����T����UKo}��=�{+ ;�$�Xݘ���e��	ձ7x�e`�R����{��V��/ ޖ��pJ�������,!3���RT�*�9GK��k)Ogw���K��<0�]|��<I2���x�e`鮅]���­6�	$���U��vE?~���߲�����*��j�vX�Zv� �엀I&V�U�U~�r쟽���~���j�K��էj������q{���'�ﵹ'{��ܕC�A�H$��"SZ�}�$����2w5I�Z-��n��c�?s�����~���k���<I2��{t�qҦ�նҶ%h;/�X]����e�b9�����-��8������l�V��v���$�+ 7�<I2�ʯ���uyOt�j��un�+u��z�ď{������$ٕ���8���M5�TЦ����o{�|� ����\���� ��<KڗJ��V:|	6� ;6<M�X���=�/z{��6�/5V��M��V�M�X���	6e`wc�
�2��n[i) �e��u��M��#$Q��aBH$���X6J��R0-�	e'$ܮP��n��.��s\"H D �}�I�vs'�oz_�	ˣ-SF h�������Tb9��А�(���DA?~�w9LGw�t�M�F��	e�dX)��3z�Ψ��3gs0��T��駱ֵ�j�����ڪ�j����,a��1#B-���q��$�!q�^ʘ�2֓Q!T� �;�����UȦ��s;���� ,�쮎�:	y�rS���;F�\���;(�UC�N�4�
&��Z������YN�D���M�У
[���M�yVnm�P��m�ge��\l�B�e�7KNW�H��-�9����U�-�@q��^6��l�e����/em�͛`���Z�'J�!ƹN�A��Wmn�R� ;�cbSj�Q۔Mst�6���hyO>�E��j�B��ql��wsu�Р��R������܃��:66V��3�=vx�\\t�2j�f�c�	V�N�U�Ħ@,�:��ÞB.���;�l{cT%z�"�+@Ӣ���u��+#Vœ)ll�ؽ$91QCk������un���	���3���b�YZ@DF��,,�T5��E�]7y6��[B�.ǮZ]��۬�F5�Ί�I������6-k��jXsF�{Gg�![��U�j nӜ�K nG=�ûa�xv�
[���Gcl,Mt���>�L��f�x����)Mvq�-�g�Sk�ɫm����&�
��v,4c�0�Ø]ac�)��⦚hY��ז9#���ܝd܂��m�v��-4󓫒�)��m�nē�.��q��V��#iqRq��N��2{In��l�J�M���#���U��Lݽ�i�Ꮅܚ����m۶�*t@m�WhM�r�#�C���K[*M� R�#+�Z�),t,�l,�=`�n�q�	B��0���0j�	�-P�-��6�:��܃�{\T�F^�!������6,cȡ�ne$�`0�P�MīWlp\%�F�nm H2�]�Yb�&U��,hA���@%�$��퉝��kk\���q��˲,��jX�v:�lr�!�/T��mJ��Z�i�,�.�.�Ȗ�W;��luu���v�t�Bv�ݺ�L�]a4���qu�£QH��(uj�z 'Q~A6l��@Qп�:
��;EZ
�@ئ�	!9$���O�s����A����r��i`�-���b5.�v���WL��q�ϸz\m��ʩu�h�WN�E��4�0sʠ��X�l�K�\�]hwk�{N�Q�g���m�qY��A�HL�Z�˭�*,�[��nBM��i�ޕ���f*.I@{/olڻ8�,J�� �=ػu�Ř�WMZ�\�''�iMSt��c���b,�akı�J��OӜ�3�ol���h�8�K��-m�v͓��N9�ֶv��(�0�9J�
�P�S.�iU��@o��	�2������W�W;a�~���yJ���N���6�	�2�����e`>�u���3$:t��?�T�d�%˚6=�� ��+ >�7fV tꑎ�e�N˵v���/o��`g��	�2�=UIl�xW��]�m�V�-�]۬ �dxݙX���	�2�����n�Zh�cSa0��V]`k�K*��9Jf&�Sl�.�1�����6��7U�ҡ���{+ ;�;&W��|������N�>��u���EDv
��;����'���n̬�5�;�W�&��v�;&V }�<n̬ ��x;)TT;\wbiU��`�#�&����ǀNɕ�j�K��������xݙXI�����r%�bX�����Kı/����r%�bX���x�	u���7��B����W/5��[�U��l6s�C��,�1e�՘ٔ-Dt���^B��~�}��"X�%���ND�,K�ｭ��?DȖ%���p�r2�)ҝ/�����H1��e��,K���NC�P�L�b_�����"X�%�����ND�,K���[ND�,K��=s�j�eԺ��iȖ%�b_�����Kı;���ӑ,t�H� Ρ�!�Ȝ�{��[ND�,K���ND�,Jt���=�Hmv�%e���>)ҜX����iȖ%�b_�ﵴ�Kı;�{�ӑ,K��3��kiȖt�Jt�{�����ؘc��<���D�,K������bX�'}�p�r%�bX�������bX�'}�p�r%�)ҝ=����������a���ER�4�Z
�<��V��lQD����\�F����֍0˭kiȖ%�bw���"X�%�}�kiȖ%�bw���"X�%�~���ӑ,KĽ��OSW#��ui��Ѵ�Kı/��m9�9"X������Kı/{��m9ı,N����Kı>ϋ��72Wc5u�m9ı,N����Kı/�w��r%�bX����iȖ%�b_�{��r%�bX��ӳ]]Il�$��Ѵ�K��D����[ND�,K�����Kı/�{��r%�`i�_�BH1!�$� �i)p��m4��𙌠�0�RD�\h��qC|� m'��<��B�{�N}����'Jt�Jt��������̛Z��>D�,K��m9ı,K������bX�'}�p�r%�bX���m9y�^B�|��ׯ]��J�Q��;m�(5�$J�������Rl7��N{�ǚ���J�ng�>)ҝ)���ﯝ>D�,K��m9ı,K���m9İ?�D����ND�,K�o�j2�M�I�k[ND�,K��m9ı,K���m9ı,N����Kı?g}��r%�bX��z;xanY�O�Jt�Jt�~��D�,K��m9��,O��{6��bX�'��p�r%�bX�ws�X\�j]h��ֶ��bX�'��p�r%�bX����m9ı,O{���K�,K�{�m9ı,K���z7�:�g3Ο��N����{��D�,K��m9ı,K�{�m9ı,O{���Kı ���I���m��1~aF$�u���42������`�0a8w/9���b��j�i47Cz��b+ڋ	��GBݗ��3]X�%�������M���K��Y©�=���m�U�q6R4��6j�X�dti���R Ū�[Xe�����\�7kA�T{&x��bȶ[���f4�8���<����a!�`�%���j\���3��w�����ŧv1�;;��U�ٔ���" �e� �d�P��pݱ.����n���Z�m?D�,K�ﹴ�Kı/�ﵴ�Kı=����D�,K�w�ͧ"X�%�{'{=uu%�f�f���bX�%���[ND�,K��m9ı,O����ND�,K�ﹴ�O�b!�2%�~���SD֥�h֥��kiȖ%�b{��ӑ,K���{ٴ�K,[�ﴛ�H����[RA$N���Ɇd3-��4��H��'���ͧ"X�%��w��r%�bX���m9ı,O{���t�Jt�O���Ck�R��"X�%��w��r%�bX�߾����Kı=���ӑ,K�����|:S�:S����q��]nm��#�2�(�W�к:\��kE��\����t�b<MfC&�3E��m9ı,K������bX�'��p�r%�bX�w]��<�bX�'��siȖ%�b~;���R�CV�F�j�Z�r%�bX��}�i�iO�؃��.���K5���9ı,O{���Kı/����r'�("dK�{��?��Y��!��Ѵ�Kı;�{��9ı,O{���Kı/����r%�bX��}�iȖ%�b}�7��MI������r%�g��������ӑ,KĿ{��[ND�,K��m9ı,O����9ı,K�w�����d�����iȖ%�b_�����K�ʙ����6��bX�'}�]�"X�%��w�6��bX�'�M��.k�#�<t<��w�v�ch��n�0���k�K͔�tHl�QF
ReM��O㥉bX������Kı;�w�iȖ%�b{���"X�%�{��ӑ)ҝ)������Em�;2[��O�Kı;�w�i�� �L�b{��ӑ,KĿ{��[ND�,K��'�>)ҝ)�������`x`���r%�bX��}�iȖ%�b_�����K!���B)V��e%K[H�""~�R�aX �D
'ȼ>��N}�iȖ%�b~�^��ND�,K���̆Mf�n��iȖ%�b_�����Kı=�{�ӑ,K����ӑ,K��?����ND�,K�����T��չ�XCZ�kiȖ%�b{���"X�%��u�]�"X�%��{�6��bX�%��{[ND�,K�Ξ�Պh�n��D��}�ʼA�� �̈́��e�U�UZܻHQ��֡"-���O��ı,O����9ı,O{���Kı/����r%�bX����iȔ�N����K���1��qj�:|:Q,K���m9ı,K������bX�'��p�r%�bX�g{��r%�bX���aO\���3	r捧"X�%�w��ӑ,K����ND�,K��}�ND�,K���m9Δ�N�߶�Ǩ�JE]B��å�bX����iȖ%�b}��iȖ%�b{���"X�F)B@!#�(�D���7�{����^B����N�f�#��@��r%�bX�g{��r%�bX
�����O�,KĿ{��[ND�,K���m9ı,O{^�]]j�Jd�*�qt���Gl�<��X�ű�bTn�1�䭬F[��lb���å:S����m9ı,K������bX�'��p�r%�bX�g{��r%�c)�������&���g�>)ҝ,K������bX�'��p�r%�bX�g{��r%�bX����iȖ%�^O�߼�b*M(�s����B����{�6��bX�'���6��bX�'��p�r%�bX��}�m9ı��;��C�Y2���O9=���/!��}�ND�,K���m9ı,K������bX�l�Q?����6��bX�'��_�g�4j㩌�Zͧ"X�%��{�6��bX�%��{[ND�,K���m9ı,O���m9ı,N�b�c�I �QI�F;'�$-�rѬ�+�<�i-�	/���<�l���g��0(]��S]Ԋ4l�j%5&P*�1c��T���XKElJ��4�-8�J�t{���u�$ոI��Ý�Ά1Ȝ�iv���m�ovL�č)Y� ��M!ZL�%��.p�	h���ԥc�Jo�������M���6z����@#�6]���c�hk��8���լ��O"h 	���k�3Y�)uac�ncWl�k�V�d2�F��ms�	��]v�`��cu�.���>�)ҝ,K߻�m9ı,O{���Kı>��ٴ�Kı=�{�ӑ,K�=����+q*����O�Jt�'��p�r�G"dK��fӑ,K�������Kı/����r%�)ҝ/��On4T�v+&�<���D�,O���m9ı,O{���Kı/����r%�bX����iȖt�Jt�������4+��O�J%�b{���"X�%�w��ӑ,K����ND�,K��}�ND�,K�=�:324i�%�֍�"X�%�w��ӑ,K����ND�,K��}�ND�,K���m9���������m#[[�jXCj��=nXB�X��іu�u�]5�g�ƎT�2j�5��ӑ,K���ND�,K��}�ND�,K���m9ı,K������bX�%�޳-����f�9��ND�,K��}�NC�p�����0��@H�Hɢ�b�! O��	�>����,N��p�r%�bX��{ٴ�Kı;�{�ӑ,K��uK}zh��Sn��ND�,K���m9ı,O���6��bX�'}�p�r%�bX���{6��bX�%�;�S��$�$̹�iȖ%�b}�wٴ�Kı;�{�ӑ,K���{ٴ�Kı;�{�ӑ,K��ڷ�ښ&������sY��Kı;���ӑ,K��c�����O�,K������"X�%��}�fӑ,K��Rq���}ե�c\$�!�˞`���Rˑ�n�r+�gb�'�(6�!�nu�f�G�Kı>�ӑ,K����ND�,K���͇��"X�'����m9ı,N�k�_�]RIr�L�k3WiȖ%�b{���"X�%��}�fӑ,K����ND�,K����6��bX�'�{�24i�%�֍�"X�%��｛ND�,K��m9Ƌ�&���l��Ød������Mϛ�3��>N!�Bꐴ�.�%+��j��"��2h--!�i�f�)`�k�Bf3y�f�M�����Qfj��I	�*´-L�X̗��<ax�Ke�����<�6'���,��T�Ap4i��;H��� �����#L V��U*�e1�3	r�r|x�H�\2z>|:j�q�>y#��&p~�d��ٽY�����YBRP 3)@B��V]-l��n��@���&�SZ�ǘ $��c1	�$�,,
��m
@ @4"P��FЀ%bB��
�K���XPG�!!5���E|�F�bIbl���iD��|S� ��>�8#�D�+�c�LB"��O�9�w��ND�,K�{�6��c�^Oݽ�H�4��\����*Y��"{���Kı;�fm9ı,O{���Kı;���l������;��C�Y2��O9=�bX�'�k���r%�bX��}�iȖ%�bw;�fӑ,K����O�Jt�Jt��}�&b�f�X�	��
��Q�3�X0��&�P������{pd!��WLd��fӑ,K����ND�,K��{6��bX�'��p�r%�bX�}�{3iȖ%�b^���N�qnZ#����B����?w���?�c�2%�����ND�,K����fӑ,K��{�ND�,K:{�==�0Q�UL�w�>)ҝ(�����Kı>�^�fӑ,K��{�ND�,K��{6��bX����Y��r�I�����B�������6��bX�'��p�r%�bX���ٴ�K���E�! �� A��  F! �$"H�"m[�����{�6��N��N�޾���X]�!����O�%�b{���"X�%���}�ND�,K���m9ı,O�k���rt�Jt�O����̪ݒ�b��buY�h)�Zf%�ZF�v��֑1[:61��p�2h�4KsZ6��bX�'s��m9ı,Ow���Kı?}��fӑ,K��}�ND�,K���$�e�4L̚��ֳiȖ%�b{���"X�%���v�6��bX�'��p�r%�bX����m9� 2�D�/���T?�Y2��]����B�����ݿٴ�Kı=�{�ӑ,K����iȖ%�b{����DȖ%���R��C'��c���.�iȖ%�bp�r%�bX����m9ı,O{���K��dN�~���r%�bX���O�jɫp�nf��"X�%��;�fӑ,K����ND�,K���m9ı,O{���Kı>W?A�*J��+HvB���8��ėHson�G�2Ӻ�V��Fib@�K����ҳ[�W��S�#ٍۍ��;��xx�^t�.����f�XG-5a�N ��7&ζWDq�n��iZ�Jb��Q���+��f�me7bnv����R4L3[yٷHjB���ɣJDn5c�K��۝�����7��\���u��]x�:�P��- A\%,�
4 R�s�0�	��p�(��~�����ӏz��=�YH����2�0`�>�`��JY�k�D�#n��+T�p8M�Z�u/LԹ��;ı,N��p�r%�bX�}��fӑ,K����� ��dK��;���r%�bX�����妵�\�at�h�r%�bX�}��fӑ,K����ND�,K�}�fӑ,K����ND�,K���_f�6嚐�j�Y��Kı=���ӑ,K����iȖ%�g���~6��X�%������ND�,K���K��4�浣iȖ%�b~��ٴ�Kı=���ӑ,K���w=�ND�,K��m9ı,N��� �[�V�+��'�����/'{�}�'"X�%��ڽ�m9ı,O{���Kı?g��m9ı,O|OO������]��Du�Xpƪ�F�w92��L�G7-�L��=b����9�m9ı,O���iȖ%�b{���"X�%��>�a� O�2%�b{��ӑ,K����/�&O�uq�X�sY��Kı=���Ӑ��B$Xդ�nK�L
�H�	�GA!!		,0I�D� �A�~q&�@HB1�F��t*?��Ȗ'��~ͧ"X�%���ND�,K�{��r%�bX��}�S�.��V�ۚ6��bX�'���ͧ"X�%��w�6��bX�'�j�ٴ�Kı=����|:S�:S�������j9�\��,K?���?�����r%�bX��iȖ%�b{���"X�%��>�iȖ%�b_wޗ%5�B��ֳFӑ,K���w=�ND�,K��m9ı,O��{6��bX�'��p�r%�bX��K�\��nr�4�7K���c�n�l���C�kQ�pك���၍"%���9Ϝ��B�,O{���Kı?g}��r%�bX��}�iȖ%�b~�]�fӑ,Jt�O�}?{������g�>)�ı?g}��r%�bX��}�iȖ%�b~�]�fӑ,K����ND��^O���e�1[�SP��9=���bX��}�iȖ%�b~�]�fӑ,x�mc �F1HAX �����}�iȖ%�bw=�r{y�^B���!ڬ�p��iȖ%�b~�]�fӑ,K����ND�,K�w�ͧ"X�%��{ܞt�t�Jt�O~���:�ZqvsiȖ%�b{���"X�%��!�����~�bX�'����m9ı,O�k���r%�bX����e�\�f�ќbȺz:�z���ۈѭ��[�߈W�S���8�lBa04��O��^K��=���ND�,K���m9ı,O�k���r%�bX����iȖ2�)��C����j9F��t�t�%�}��[ND�,K���{6��bX�'��p�r%�bX����m9�B����#�,7
�y���*X�'���m9ı,O{���Kı/~����Kı/��kiȔ�N����o����kP���w�>,K!����ND�,K��{[ND�,K������bX_����B�E�%()
����K�!,f	��4
��(9�0y� >>���zk�^������ �cՒ�kFӑ,K����6��bX�%���m9ı,O�k���r%�bX����iȖ%�b*�{�_�&kS.��M�`�niNb���t��9�[�-��� $L15�%�y
Իe����N���������r%�bX��׳ٴ�Kı=�{��r&D�,N��siȖ0���;�J��e�ʻo9=���"X�����ND�,K���m9ı,O}�siȖ%�b{=�fӑ ���	"{����ɖ�Y�M�$����fĐI���&��'�Og���r%�bX�����ND�,K����˫lոh�sFӑ,K����6��bX�'���m9ı,O}��]�"X�%��{�6��bX�'}'g��v��L��>)ҝ)��ﾾt�ı,O}��]�"X�%��{�6��bX�'�������ı8�@D�$<w���왆!��\�1�X�J���ku��.6�h�.9�>�H]��D8oufղ�wi���³f�R�+/
jX��HQ���u�5��Fn��wr���:�Q��C	��8�\�s �1��ѷ�kM4m�ݴ<
3�N:��"�ۇd.Ms�Iػm\���&��C;9۴j`k#N4��s)�Ony�+�ৱ��6U�����R��'Ot���� �!�3�٬m�LCp̩��\�#n��IЅm*����f�n,ț:����}:S�:S����w�iȖ%�b{���"X�%�}����"X�%�}�{[ND�,K�{|��d�Z�i���å:S�:~���iȖ%�b_}�kiȖ%�b^���ӑ,K������r'�S"S�����iv1x`\�Ο��N�%�������bX�%��m9ı,O}��]�"X�%��{�6��bX��w�����j��]�������(�ș����m9ı,O��w��9ı,N����Kı/������������K��I�*�����bX�����ND�,K���m9ı,K��m9ı,K�{��p�N��N�Ͼ��V��#H��:����
sX�f[v�C�>��m�IAΨ��9�d�Y5u5n:ՆK�WiȖ%�bw���"X�%�}����"X�%�{�{[ND�,K�ww�iȖ%�bw'oi:G%.h�����B����w�i�h��Pv��n%�{�}��"X�%�ﻻ��Kı;�{����N��N�߽��XUַ(_8�Kı/}�kiȖ%�b{����9��XdL�����ND�,K�Oߞr�9H�#��R�<������C�fk[ND�,K�ww�iȖ%�bw���"X�%�}����"X�%�{�{[ND�,K�z�/��Y��I0�kWWiȖ%�bw���"X�%�}����"X�%�{�{[ND�,K�ww�iȖ%�b ���~�3Z�0�1A�'vL�3�y��f�S6�YFp���WfH+�"��RŬ��?:|�4KĿ����ӑ,KĽ����"X�%�ﻻ��g�ı=����iȖ%�b{��m-�h�u)���ӑ,KĽ����"X�%�ﻻ��Kı;�{�ӑ,Kľ���ӑ,K��޳v��5����ֵ��Kı=�w}v��bX�'}�p�r%�A>��hB=s&R)�#.�	��E��� �R� &��+A���Ȝ�}���ӑ,KĽ�}��"X�!y>��C����h����^B��X����m9ı,K����m9ı,K߽�m9ı,O}��]�#�^B�~o���#��a�t�ږ%�b_}�kiȖ%�b^��kiȖ%�b{����r%�bX�{����/!y�ߴ�7�]L����bc�r�e�Tkz7T��H�5�	j���йՅ]kr�����ҝ)ҝ/������%�b{����r%�bX�{���Kı/�ﵴ�Kı/~��f�sYG�WΟ��N�����{��9�X�L�bw���6��bX�%������Kı/~����O�C*dJt�{����#���W_:|:S�:X�����"X�%�}��[ND�,K��{[ND�,K����iȖ%��O�y��6�"�,�å:Q,K����r%�bX��{��r%�bX��w�ND�,������I	���V 2��� T��HJ/U�;���ӑ,K��޾8�[��r�S3Z�ӑ,KĽｭ�"X�%���~˴�Kı>���iȖ%�b_w��ӑ,K�?�������e*J�CpR.:M��vL��F�69t�KI�rh	�9��˭kiȖ%�b{�߲�9ı,O���m9ı,K����r%�bX��ﵴ�Kı;٢�d��5n5)���9ı,O���m9ı,K����r%�bX��ﵴ�Kı=���v��bX�'�^�z����k5&k3Fӑ,Kľ�}��"X�%�{��[ND�,K����iȖ%�b~���iȖ%�b}���tK�V�e�å:R�@�~���O�X�%���~˴�Kı?{���K�� �?���m9ı,K���4[��<_:|:S�:S���y�ND�,K���ND�,K������bX�%�{�m9ı,L>? ы,y,��.�Mk2nY�F]�T?��˪v���2�J��Y���f��cp�>LQśc �Q��	͟�k�I���S5���`e��rK�	�}��9y���.��(Hr������&ȠA�Wa���Sfs��&��[����*���
�t��k��ʺ��j�k)���IN2�� �D�B�K�(Fp$�i��t�����J>?z�A���H ��`"	 �?=�������@?��#$���XR��:[k��~`;Y�4HB�'rf@��Q�4��2H��;��N�b������ؗ�� h	@[��`�������RS��ç	�Vh��f̲p&�a���҆2㰒jV,�S�! B	�f�o4����L���K�n���a�5rS.᮷�H�f�ւT"��!������Q�vn���.�'�b:Kr`�b0#��))+(Do��7�Ms3\�ȐV�r A�!��Ƨ5͡T�B$�<|�U��U5j�
� �YV[f9Ѯ�J紋[*�'�T�α��"�(�՚�i]�n���L&.�[��[�%����R���
���±�^���5��N��O���s�H�n�v���ň��t5�CZEEvV�ױ�%kua��M�S�C�֤�`:θ�$�G��t=�m��]c��l��1h�&ԫrm`�P�m\���B��Z�w���z�m�g�Tz[�B@.|�ʅ+��+8C�F�p��z����T��4��%�Y�*2�4���ve���+�ˀ�O@׎C����:vR/n5<ctN5��ڮ�ݗ/e7�z��,&�����+�Qe���]�]�7���<�j8C�ON[��]�J=tgav�l���JHު�N����fn�KC#V���19��Z�UH�̰�m��R�Y�@����9�2r�Gf��4��M� 
�L�`猝8�+ŸnӶ�v����Q�����y4�solEs"��y��B�Y����g,KM)��j� �j�]�	�k� s��� *���;`7!+61�!��,��h�+�y�v{g��˺�TDl��RY��yqq���DƬp`��\��d��&:Q�q v��N�*�� 4�eyXk��ڬYz�#B�����utYu��
�ɠll���5��Tl=��W.�ti�,oJK���QT�1�z6�+���5 ����(h��,�0�X��4�6D���v� ���h�l@�m���'�v;sH8��]9�Ѻ%�������K��VUR�iM�B����g"�學qV�3��R�A�v3��:�Ǜ��ta�1���]�e97	�u�����e��۷()�y[n�(�jm��A��5O<������2��;=��,d+ͪ�dm��zbs��Q��pt�q;�1����NI�(��y�U�)b����mR�طme�-�	0�-	����=(@��E� v��થPN����6ע;@R�PPؑtO�D��D1@&�~P���j�Q��k2K�L�˔�~Z3	H�MJ)eZC-�[XD�@�!�e�a3De�4ʥX��v`��H��	v,vt��]m�$$����	����2�Վ6z6��ڣ:��Q�m�8�0�F����gm�`A�Z�� �Y������\�!�1LL�t��t�=9+=/m8����zw.EgiG�B�Μ�BS���;5�\�78�Q�Q�ԡ!��2��n{K�A.zI>t�����k\�Ӎ'��B�=NZ�Ǝ�M����M��"j.D(�v�����@4ʺ���҉bX��}�iȖ%�b_w��ӑ,KĽ�}�����"X�'����gå:S�:~�{��c�+�<ND�,K������bX�%�{�m9ı,Ow��]�"X�%���ND�,K�w�8�K�љu)��kiȖ%�b_w��ӑ,K��{�e�r%����?����iȖ%�b_�{�[ND�,K������]L�]3.���"X�%���~˴�Kı=���iȖ%�b_w��ӑ,Kľ�{����������u��p1���k.ӑ,K�����"X�%��!������ı,K��kiȖ%�b{�߲�9ı,O�@����Y������ֆ�d$�f�5��)�� �ʛ&�vZ��C��1�M�-߼~�bX�%������Kı/��kiȖ%�b{�߲�?�~��,K����6��bX�'��r�kW	sY.���&f���Kı/��ki�uQ��P��;���'���˴�Kı=���ӑ,K��{�ͧ"X��N����LY�3YZ@r���ҝ,K�{~˴�Kı=���iȖ%�bw=�fӑ,Kľ�}��"X�t�O�P��1� �*��O�Kı=���iȖ%�b_w��ӑ,Kľ�}��"X�%���~˴�Jt�Jt���7�͵�b���g�>X�%�}��[ND�,K�C�
�������%�b}�o�.ӑ,K�����"X�%�����L��fMk�ı8�j�ZG8�ֱ^��Fi��6#X+\�u�1^,+#6�f����ҝ)ҝ/��{[ND�,K����iȖ%�b{�{�����dKĿ������bX�'���������3Y�m9ı,Ow��]�"X�%���ND�,K������bX�%�}�m9ı,���u��u�Q��'�����=���ӑ,Kľ�}��"X�60���P��a$D��Cj<Q:��D��涜�bX�'����iȖ%�b}���SZ�,&�ѭfh�r%�g�
2&{���r%�bX������r%�a}���w$�{��B�m]
݉����vG�M�-`ve`ݏ 6J����4�A͇j�bcP+���{.�6y�=T�Wɝdy���k.DZ������e�n̬ ���� �"	��N�k�][m��&�����Ur� ��x�O<n�k ���]ڱ�t�	6� �/ $���j,I2��E�P�O�.�-��	$x�۹'{��܈~O�" �}����'b��Z�i�+����E�I&V�/ $��Av�9��+V�	E�'n"[g����9�\jV6��ձ�BQ���jj�Q1���ɀ|���	$x��ݴTUnЊӦպ�>Se��<wZ� �L��U$uz�g�bj�6����$j,I2�wc�	�i�[N�E�x�j,I2�wc��UR^������:V��\*��i�I2�wc�	$x�j,�ߩ�ԩ*��i�O�<`�1-�X�ᲖҐ��4��*%GY�n:�vY�笏0�`��e�`cE�ReVg����i-f ��G�ڭ��2�vz<�ƴ!��Ʊ�T֜"�3X����dA�J��n��JE�C&x�]�{:<�])ڭr��J�:�=D�ioVqy�w�Nc��5�A�jg"ȶ�7m�X�ȱm2k.�8D��'t���3�1���R��Y���m�
܁�Qu��+`�έ*�c��Tu�qvn��x$� ��Z�$�+ ��J��j��M� �c�&떰�2�nǟ���q"o�5�*��j�|Wv���`6e`ݏ 6lx�(Z"��V�*b�k ٳ+ �v^ l��	���fݢ��v�P�յn��e�͏ ��Z�7��y<����N�^�ɘm�1fڠźm �Gk�Ԥf��$�z2�Հ�@<N����͎�+v&���n� ��x��f̬.� �ȋH�;wN�Ez����v���c0=d��� �IjQ#�"P# ���*�\Q��y��7$������ݏ �E��Z��⫫��Xf̬.�=\�����=��k �ɖ���մ7I�+n����{#�$�-`�2��T��$�[TՎ���G�I�Z�;6e`we�(�`t��!k�q��jጤP��&�@�s5a/���g�=v�Ggt�^��I�Z�;6e`we��G�wmI"N�T�n�ٳ+ ��/ >�;K �fݢ��M*@�յz7$���srIϻ�na�qI!���XĂX$��$"$%C��:*��Uj�9[��������:�K��t��-��B�x���	��XwfVv^ oa*�-��um4��'c�`ݙX]�x��������&����4�&9�v���<>k��b�h�@`��k1Q�uf�(��6V� ����Vv^ }�<v8�;&[��V��'@���"���Id��q,��L�:��-'�h������G�N��;�2�����Q�Z�j�|E�x�q,�&Vv^��*�33��[�}�,����j�-�TҶ�ݓ+ ��/ ;�<vo��o������(ۙu�BT���KX�D�[}�+샷j�U�b'�9��7G5��;un���O\��� �K�UU|�g���j�<��Ҷ�[M��m`wc�7c���L�e�X�%+lm�:������X�&V��X����,���[e1Uն�X�����z������nɖ���մ7I�&�`/b��O<O?Z�>�e`�\��jȩYU�9��ӳ�j�Q�����ʐ��5�v3��LF3jB�Ņ���R��Z�Ԫ�"^����5�2OPcqF�Ҙ9�:8�MU�V��#p)�Q
�+n�Q�������ӧDnq�&���-��4��@^�5�/ۭg��.
�0�\K��l���A*VB�-�\I��4�u�jx�������X)�;�Oi�[�d�ɚ�h� D{������g+�:m\�5��l�BN&�$ܑԕ�rĴ�I�t�=��ڄ�5%j�����7�����_�ʪ��yl���T�^EZCWm�Zm���,vL�.� ���UIZ$��;��q���o���Eݗ�v<�]ŀoj֠��ݢ�;t�۬.� ���u��	�2����ݷIۻM[`]��v<n�;&V N�x\�.�v�t�]S�Rt��b�D�Z�5��grpLhe�����j��[��V�@�x�j,wfV N�x;����X���m��WVۺ��w��ٿ���,B@` H�"$H��(�
�`I�< ��x�j,�W9I#���Z�m�t$۬ ��< ���	��wfV�ݕ���hmSV&���W��x�~��Nɕ�E�/ ����������&떰	�2�nǀv<��9ʯT�{��@�f�j��8��B.�#����	��i؍dE]h�LhjkB�%WB%ο ����	� M��	��{V�EM���۬ ���ݏ ��Z�'d��:�"nۤ�ݦ��o &�x�r�W�Ug8r��2�T;�	C�# �]	�e$�%�6NҘf]kaj��+�����C\��W�)���^a�%bH��~�_��3�3�������c�&�U�R悐�l�L����y`Gp,ַ��j�>kb���
Z��>?;��K�	O���A��h ��cB0>�m?~7�����0P�@�C��p :pQ>A���@f (`�^��N ��(~E��(TP�)�ﻯ�7$�}�u�6���ٖ���:����=#��wfV M��wc�;["X'Jպ�����v�	�2�nǀv<n�k ��NhFB!�һ26M�[۳�84��`��F��M��s��Ja���� �v^ M��	��W9�o���mOx��Wn��5bn�nǞ��G�~��{}�-�x�T2�*���R�m�u�X�X[��nǞH���z�bm��n������e�ݏ�J+�(���9��#J�B"%�[RW���<�R��J��+ʆ�	��n����nǀI�Z�'d��Ww��Cx�\j2`f�U�!��p4��Kv��N4nm���m�Z)�&5)x����x��vL�.� ���[��V�@�x���U�W=��V�׀dy��*�%Ox˧tYn����6�X����E�/r�ď{�x���;�.'eҵm��J۬.� �c�&�Q`l��>����Ym�j����7Z�	>��ٹ'oﻛ�q�R�R$�(Oߩ�UiO��4հZ���(\�6�'m�.�����`�m�ku��v�H���h^�A�.�,F��i+�]H<d#���1P�߾�؊[]+e��0�f�+��(`.*�
�X:�vZ�*
���9(�#��P�.�Ռ͌6�b��t@68	�f���|eͥ�.G+�eQ��0	���d���;���ˈ۞�\wjhYD��3V������o{5,5y�`L�Zu��O�];���{p�1��YfJ��	x��ְr�+�o@�c^X͙X]�x�c�7m R�c���i�f̬.� ٱ�u��ҭj$��&�ڷX]�x�c�&�Q`6e`)������w����%=<�Hז�fVv^ od�Eӷt���m�n�ٳ+ ��/ 7�<m�c�;`J�mr�.���U��FkI�JDˣYf�0���I7lE����Ŗ��j��m5�vl��"���웼���'����t����;ۢʎ�\֍�;}��@��� �rw|�	�j,�fV�#��&���ڦ�M� odx�j,�fVv^�؆A*���픭[x�W���o������{#�7mA,)�m�)��Xf̬.� ���	��>;=-����5�j�)�ƌ��Yn�����v��M�m��s.n���Se�P�փI1�N�6���׀�7Z� �ٕ�|��n��Cwi�]���G��r�����6Oe`we竕Ăo�v��n�Տ�M��5�?}�vns�#@$2)# |�;:4y���޷$�ｭ�?wT���Z�VPˤ�M`{����=�`�y��#�&�Q`v����]�Zi:m� N�x���	��XwfV�oU�r�m&��ZN�Z ]of��n�ݔ#S�Fz0� �����ݳ��1��Z�M� �dx�j,��+ 'v<k��Ui]�)m�u����RF�� ��< �dy�s��%���We2�)��X�{+ 'v< ��x�j,�U튈�ӡ�7v�ܮU%�x�y�u��5֍d��VI@�	U���`�H7m�V�i:E�x���	��X�&V N�xT�R�p���	Zx����m�1���PûG4ƹ[b��S5v�S���6νk�&�Q`l�X;��wc�;�R�e��2�.�m5�}�2�wc��c�&�Q`��t]���:m� N�x��xz��T��k� ���>��QRM+�j�6���n������9UĽ�� ���ׄ��iZ�q[w�M֢�=\�;'���=�}��9~���'ς�1@a � �b A�}�K�nf�k-+�2��rYss�S�Fv��m��dVH�����F���F��T�6B�g}����q��j�Jl�)Ξl�D%���qĶp*��b�SN�V�EҒ��̮.s`�e��.ѻEp\��^;t��E�+ifLCV�k`V�Arp[�Z�󥮞N��q�·n��u՛�ΐ�n`K�8�-)�M�C�[A�vw$7:ɱn^iU��wHtﳧ���<7 �m�5Iu�G��	��e�T�y��r�\�g=d����6�J�]��1Zk@���+ 'v<�6_�s�ʯ�zF�����*<������� N�y�s�I^���5�ove`)R��t��i�N����6^&��ٕ�v< ��ˡ�v텏���x��{�+ 'v<�6^��#��n�E�I��`ݙX;��)��	5�X�T���F1��]Ԍ�n�P0a�.F6h���h:VX�ft���@���I�:�� 'v<�6^&�k ����;[r��1XƘ�Un��>Se�j����*���r�,�>��&ɕ��{��/g����`G^ϖ������{�+ 'v<�6^ݴBZ�)�����7�2�wc�>Se�{�UT�鞵�wJ��Q�&�Lvպ�	ݏ �M��I�Z�7�2�r���s������3mj0����Scb���1�VA�^lB��q!'\�v^uZg��Y.Em�W�� �\��ovev�@M��'d��n��ac㤭�������� �M��ob���[�Qe�۵�ove`�ǁ��r���W9AB�` `�UC5���������p:��D+����M:-[u�v<�6^7\���r���}XԿW�	��4�vU���/ �r��1y|�� ���	(�e���'VЛ)���Bj�nG�\��x1�ui�+�;<�:9�7t"�iZ�q[w�M֢�7�2�wc�>Se���B�_v��i�{�+ 'v<�6^7\���W)#�U�</![�*�u��� �M��M�-`ݙX{r�-�����Yv��ܙx�r��ٕ���8�~^����޷$���d�kZ���0|t���&떰�̬ ���)�����}�t���۱)����-Dy�C�6�F�nϚSN�Nt y��!e܍�E]��v��̬ ����c�9�����}��[~C��1bd5ң��7c��ǀM�-`n̬��R���cL�eZm��#�&떰�̬ ���]���i4�[)m�u�XwfV M������B�_���n��ٕ�v< �dx�r��9\Õ��
�%I
D�/y�k)NCH @�))+iX��7��JH�+�ﴚ�&������Kws7�.3&�� �F��C���!$�8C7�?L?k�ٓ��������������������]����'�UZ���/��v��	��� �R!�	�%�X>A�H3�G�w�w��Ny����4�����g�\�@"�9|s��PC�P�"M��*�|��~��By�Bqt,�}��P��y�mfp����3�;.����r�d*_��M!w]��b1`dA����tQ7�5β�|���~�_Ne����s��+�bu��(uIQ������	5ϰ�߽��
g%�p���d5�e�������h$%�$��S�)>IG�=�{��w�kl��5��~c�dd�RP�O�ʩ�_"� ��Ѽ1�*,*f������~BȄ
a�FǇ�4��~c��R1A�3Z&&\[��L�]�N�}����U�_����B��I�U6��	�6��p=���J�UF����b��V�"������ۘ,�ع�ˀ΀��W���Ve��,5H�l�ֺT�d��wl�[R��U0T�K�J�F�{U���V���;j�W�3��ƥ�}�����<�����c�(s�x�4!K@�=K��W��@r�v1�ivbm3ێ�s�8�I%��^�V��B�t$\pml��Xݚ:)�Ta�������u#��$Ţ�)� Ԅ 5@�0��mڳzg�e��`��#���WFB��G�qYy�U����G;3/�
E�E�0<��ی�7fG��ab�vq͜ OF���[)q�5Ŵ !H����\��.l79��k")BKl*�9�%ұ��]Ύ ]�p���"���ClD�V��FRy� ���jq�uT��e�D�A&-�U�6u��h6��7\���	�]�l�[��ݦ��nJsu�Y]qI�[����f ]�`���i���P���]��������`wT�)v8xڡ�`T�t��g��Ӻ����P%���R�2��Z��v�@tR�WY-�3FL"Ͷ�T�0��C�v'�x���.�F��;�'���2��j ⽮#ՙ�#(��c�&��mΡ�Zh[,�mb��oz�ɮ�X�;�
⨬�THk����-N��lpu�%}����C�m�6�Ye������'���Ύ�lMLm�l �<���?�B�{\U��S�N�"^ (1F��Sb,Պgq-�CS[�C��Z!�J��:cV�z%�wY�h�ݭ�#H�ik��rB��T-�U��������d�Q�<-�;Ҧ��u�uX��,\;#�XkS3��InD�GZ�ɭp����1JW�}Q���YU�	��*67��;�N�r��Jd���:�V�Ik\���+NvG�bUPvp\&ͱ�g@��r��c[��]��'(�Y3ԁ�]LA&��v֭��T��/m#�`4�N$Ty�rft�\�^��V��4v�I��L���!(kZ�m֦�f��> N #�bQ_"��TН ߕP����O����	U�����vw\�¶�99�Ѥ�27m�xᮃ����x���EJC�t�c6��S�=�x�]7mR��n+h̹N��W��Q�!���k�����h�k��,��m��mH`�7]S7]GB�mlЄ�	q�-�م���j\Z��1.l�T��-(6����v���\��\ls
�m6����#���4Z��L��ml�� I���Ӂ�f�I������R��2���od�����N�}˥sZ�sf�5�*� ��� ��� }�<n�k ����;ەm�$�J��˶���u�XwfV M���9Ig����[L*����zG�XwfV M����얖eZ�VQWt6ݬ��+ &�x���	ے��l[��ڴ�Av�`ݏ >�;rR�;����o��}I�%f������L� ��Z�Zѩ"�ê̖�)�2�ka����
�i��M� �dx��K ����	���Iˡ�Jղ�v�;s��� @���P��0��� �(
듞�6nI=ﻭ�'6G��s�ĉ-<]+��O�[t���X7c��G�Nܔ��V�
P�`�Lm�u�v< �dx��K��ql�����y���vݪ.���G�Nܔ��̬ ���O�/��6�ƚ��l� �J�梞��79��q؜�+���0�ޠ����Ͱx�V�;rR�>ݙX7c�W9���<��z���V�
.軷K �veg��U$�� &�<v䥞��s��k��wWam[�tm� zO< ���nxT��@�HI�H��Az��M����.�{�ٹ'�>�%Ժ���;*�o 7�;rR�ԗ}=���� ����Ui4�[)Zm��%,�+ &�x���	[RRy����m�Ri�5�͙I\�D#��
���±��2,))�Lsp�� �l��	� }�;rR�;ڴER��MLm�u�v< �v<v䥀}�2���Gi��ݥCae�x���	ے��ٕ�v< ����h+�!3η/��N�����|	�����'~��ܚ�Υ�B2�6'�U��铯 ���VU�vQE�
���>�2�nǀݏ ��)`j���Y��̖�D�v,�z۵lRN�ym��#9�U��,����$D2�n�nǀݏ ��)`M�XV�W(V][Cj��� ov<�9UI���`��V M����N]%V�Jղ�m�v䥀}�ᇫ�H��x�<��EH���ڧƭ�Xݎ7c��c�'nJX{V��XջhBm4��7c��c�'nJXݎ�*�R���x�ut���_���|�iS���ʰA�6�Z�;@imQ^(�iB7c�������:��	�3�>��ba������Fr�N't�1כYum��6s���[�4b�ː��-p���f�����B1T+.��J�WJ��ծpIIX��r�f��I��ґ֩t�t�nf�8FŲ�i
�U8Ga��S��n��n3u9�QO�PpXQ{���W9�j�%Ӭ�՜����N�%��+Z�hY�]��{'5K� ��m*�`�����������rR�>�Ȱnǀ숺v�m��%,���;�<��y�[��﷝���~�jyF�se��v�ݹ�v< ��;{�w�jTe�ҫwn��%m`ݏ >�ǀN��`{�ʪ�.�X�^��V*���'�M� ��;{�}�ذnǀmH��m]�B�wN�e�.�ۗԝ�Ig����n��cL�a���N2����!Z�R���'o`��{ M����x�,/�ջ�Ʈذ�{9O��Q]�s�L����N��`�]-*[J�hBm5m� ���{��������<,�~��;ە��e�N�Yv� w�;{�}�ذnǀ숺v�!�;J��'o`�r���_ zO< ��6�[۵�1��pl�i�n"7>MuƄ����"�W�\�$ݱN4��ZN�1`v�, ������	��,��J�]Ъ��T�j�7c�	ݏ ����'u� �ڊ$������Ui���;{��̠��T�ʂB��$$# H}D,�t49U�+�W�{��`�<�	5!ˤ��iZ�R���'o`�	�p�	���+���y�Z9�X.;V��b�'u� &�x;����X�$IZ/�#4m��0�3h��{4��&�*Rz]s/lu���e�t��c3[�ݏ 'dx���\���=#�n߫�ݱ	�,N�"� ��窹�q#�s��=#�v< �H���ݱ�Wt�M�v� ��ٱ�� �d�avU�v�����Ł�r��T�&x����	���*�p��dR`E�O��?������6X�Wt+-�����0�c������6l��;��iF�-�TݒQ��#�..iwIy{V���c��o<*Z�d�� c8u�f�]l�_ >�������fV vlx����Ui4�]1+�����fV vlx�c����G���^�qڷt���==��� l��������+���HM�wn��c����*��Iӥ���~O ��{=s��e�c�o 6lx�䥀lٕ���b��0X��,�m����rY$��~�Z��V��1t��K�8�A��[{���<m��t��)�4�6Pl9�MQ��/���.c\�z%Xۘ�6���-���5ͬBV1.��9U�s���n�cj\hَ�q�cc���S�C5b�`�..�.�b�M����bGh�)h*J���Ģ���(K+�f�=�A)cl5(U���e�2���8�i0 ;r��?�;��;������*�\-%pnXq�uz��)�J]+�P+�0e̦V�;pQ�Ͷۦ�]�n���K ٳ+ ;6< ٱ��e��Wm5J��J���6l��͏ 6lx�䥀}-)wB��j�[u�� l�����fVݎ�+[E��T���6<{{�I�+ ;6<f���J�&+.���x�� �fV vlx&ǀ:�T�T��&�M���LF0��1r�2ԵLм`���+	����Ŕ��U�j��ty�%��ߘ�|�������_tX�WKJ��n��6���7$���u�<��8�x?~{��mI&V9\����y۶!7E�ӥj��	=�oo`��2��c�숺m��E�6�o ���`�e`fǁꪤ������˫���j�%t��,�L� ���vG�oo`��Y%�	������6�1���%�oe��9�6N���PfgJ�·�V�lIX+-���6�`fǀ�<{{�vl��;-IlI�����![o 7�<I��,�fV M���I4T��V"��S�o �{�'��ݛ��t�X�aqe�af��IXXr��9��.}�\��ٮ׼�̹M�.�/�\�ݺ�b���ϥ��:�JJ�s9�x�̀MSs2RZ��L5���f���~)32���f�ک�E~�w�`w����y;�־�{3}���рG�jE��j|F�`�9F!p%2��q!v��a'cG�>��o�㳚Ͽ)�����f��>�y���]w3w��)���vR��J�X:@븽�;MwK�BU�����]&'H��@c�J;����:wi�~��Ƥ*j
�hƅL++/�W�W��!5��ؿ0�f�f\��Bh��}��m�����N�H���3P�!�?)0�B�Ņ7��M���/����*����qZ�����i$��&�� ��	R7	pA%e�)J�K�s�k'Cd�W	'��	�����(��^i�Ed�q4�I��0VAD���~�L���	������\�����t��/WH'Q
�~���� �Ub���GF�BI| t�/ʜ�ڬ:�ý�����,�������X��H�����ݱ`M�X����c��r�ʥ�9�`�t�W~-��6��u�� ov<�{�}6eao����f�i����ة�����]9�n9�f֞K"�t&l�Pݗ�f,b�"t�m��c�>��X�fW��UUW�	'� Wg�����lE�0V� �^�`M�X���ݙX{�V]]�um�t�Э�`M�X���ݙX�� �mHЕ���j��� 7v<{�+���煁�U|s���Ȏb
1fTV�k�4@����)JH:T��8&��T��߿��rOY��k%������"�ove`K�,�+ 7v<�9ʞ�����:I��9�n�z���&�t!(s�g��h;sWmGe�GD�M�+�EҦX���w�<,�+ ;���U_ �=��yD���q1[�|��ٕ��s��) �<�	��X�{�w�t���[�`;cwn����ݙX�{�}6e`��\����i�M[x�UqM���˞;�+ ;� W�D]�m�˺`�����`�2�����2��w����LQ�""�:͍Ԕ$����`�2.�����=��0�˰k.�0k1�iXCMe@F��u�i�Y�u���[��U,e�ވ�n����Z�9��̦�[0F[��8̫B��<!���TlBº��a�*n���E�2�us��FCնb���1aIB�s,&�۷G1�#�B�t�@\�2H���:�[�WY��C������94�qQM_�i�I󻻏������c��GbU52��kg7�W;vy�`MӤwF8��t�`g]�5��WE�b�?{�������2��� �mH�+B��j�[u�ݏ �ٕ�}��X�̬�s��U$j��lI����:�[o ��e`m�;�+ ;�&���Wt��L�۬��'ve`wc�'ve`j\��������wfV }�;�+ �oj,n�qYn�mݔ���T�i)4؟]��;k'V�i�}i���� �%v]e�e]�݃�-ݺ��y��2�����'ve`[���MZtU���浹$�ﻭ��U�P�!!�H�%bш��: ���ٳ�rOl�V }����Ǫ��v�;Wt�V��v\�,wfV }� N�x{���쫫l��]n��'ve`۱��ǀ}���ֽ��E��T�jۯ�;'� N������&�����������J�iqxZ��bd�uKf+(��ՠ���x幦�ɈCG]�)
���X�����x�{Q`ve`۱�h�˥wH��T�j��>�ڋ ��+ >ݏ 'dxZ�"���1�wt�7fV }��^�F'�!�Q���\B������nC}r�,���Ү�n���V��`۱�� �oj,n̬��R�i5i�V�շ��<�W9U5���I� �lxU��!�I��t�5�I�v0���H�v�ױ�-���	�1������L�0+��v�]��?��w��}�X���fǀwv]��՗V�t]7n��6l���ǀ6<����>��h*�V�T�j۬ �lx�c�;��,f̬ ��R�][E6:�[o 6lxw]ŀlٕ��+"B@$#	�I# HIH���" �������;߅N]+.�v�1+�����L� ���d� �s��+ޤ�'HWH���t-%����R���� �jB1��4q+�F��h� r�5]&�m���|�[N͏ ;�?W*�A�?5�w�t�W~-���*ݺ�͏ ;�<��5�wd��W9��)#�}^��C��V�շ�=�wuư�Xٱ�IRU��wt7iSn���5�vI����d��$�WV][tU�WN��2��c�5l��wuƷ$���
�X@`2A�V�8�t�_ſ���mF�M�1U�<�G..��1G��+$u����S��k`3 (筛tjK�R�x�4���^t9X����Z�����MOb�=�8��+,Kh�LY��O�=�ڞ���	���U5im��3`r�K1^c 7����8M��rrc�;`��*��i��mrt�iԥ��*�Y�:{T��y���v�t�XTX�c[4����+��>Γ�=�I����E��j����D�����n��Vx�H�*��(�ۮ�'�9�ki�WWe�j��u���d���5�vI�����l��,Um���m�)�^���;$��͏ ��S�J˪j�Lۼ��5�vI����d�-K���;�i���m`�e`Se��K�;��XҮ��w˦�Sv� �/ ղ^���;$��=U\��_���n�u��qM˹ѫ+Zwd%q0ca�W[��BW�G-�E �8u��U\��=������6L� ����jJ�Wj��vw�}��o��8@���)�&fiXf`�h�14X��W9U�{��X&��I/ �I1U���t�ӻm�I2��c�"�^���>�ܷE��c�@��͏ �l���5�I�+ *ně�.���:�[o �l���5�I�+ ;6<�5-�j�:*�uc�D)���x�ivL�ͅA�X�˴�s�1mV#f��t�4Z�0Wn���&̬�l�)���T�R�;�i���m`l��:���"�/ ��`K�Wpl�tS�7v� �/ �l����#�P���	w~Ӎ`�2��r��;i�v���xw\k �fV�6^ W�RU�n��*v����q�M�XT�xSe��*�s�Ъ�T��hg�ᰜ$*L`�4�[6�t��	9DNF/\]�KM��c�c96Ƕ߻�|�P�/ �{���>�9n�E؆5N����:���6^ŀwuư�2���I����ӫJۼe�X�k���2������QSE�;��k ��-`6e`SfnM~C��G��aJ�c��R���2��
J�m$˙
K�D�02�Mc�<��+����� �:#jZ�]YM�n��fV�6^�\0�r��i;B�Ot�m��v�T�8]4z{n�!�ͼV@yCk�ڋ�wXᚶ�`��V���kwn�W�� ��w\����{+ �߼�i�E�6�����$I�`���l� ���X6��U�*v&�w\��N��l�n�`�&*�]ջ���զ�����U/o����׀M�w\��}59n�E؆5N�]� �/ ~�Us�}��$�s�u$��k�'������� ���򠀪�W�@Q��* AW��W�T_��UYdB@T#P��P���@T �P��EBP� �/�T_�� *�𠀪�AU�
�W��_�P@U�AU��W�T_�����@U�b��L���v���9� � �'����`����T|}``�-l���p�ۮb��Oz�f�ڎ�|��       � @   9��8|P($�gx A��;��i%.zn^�J:g�t�j��/ZoS���ޚ�l���ͦZ������ PP|��z����Mtfq���ӭY��+�w�u2��oc{�n<�u���w==�^�ɯv]�|  �{ޛ���Z�7q��8��ͯC�=���2��x,��{����:Ѽt����֎G����� ��z}q�ڬ= = Z�����r ��X ��|���G�6|�[zУ��C<�k�����)B���c��֞�coUq��z���;>��4�>>�}5��}z�o����o�K�=�OO�P
   � �$�HѢi�� �!�da��R�Sʍ4 �M2dhd  �4�IJT�A��F��i�T�R��i�`� L� �"" ��F�a��6�M6L�ɵA T���L�!�	�އ�����z�z{1��<@q���AT`��!�
*�������3��?؞!d��Sb��0�� ���`"�;��c ��C�޿{[Նy���ν\}9�����������ݽ��#�����wwwwwwwwwwwwwws؎��}��ݜ;�������������";�����������������s����������������}��ݝ�����www}�������=��]��=]��ֻ�O�����{���$�" � 誾�� #� \@_EW� En '� z*��>�� ��z z /b �@�@�UJ� %@@� }=�O{��rg����0C������û��݆fp���wS�v�q��sɋ��.��Um(���ve�y`XNP)�$�F�B p�L2��vn �	����bm4�gBa"Hn]�3TP1x/ �h`F����hy�ٲ��Cu�t:�Z�K5�`cA���6a��!�6�
maE����q;F�$69��f5��(����TS[��K�p�0��bHI��I822�#H4�m2�xz�@ �D"j�tXv�(��
����{� `
D���1ڝ�-��19y�Jk�9�&�\�by����PB��1z䲡�2�)�0B0YS"r0�m���u&�H��L)���ү֌���/a���^� q=�کł2L	��@cc�����7B\@Џ�rFu�o �ʻ�����4�Ċ�*I�ǐXQe�*�*3��3
�Ce�r���+Hԫ˦V��&֕�� Sx�+(�֙0d�$)ִ�-ÕѨ�̛l*D�)���*�Xv!	�P,6Pl��V�*UhK%X���m�A��n�q�8�MDd���F��g��8�����&)`S�,��-0�"�$X�%�ڌ��U��X�[� �ZM&�%UF��N#V[
mH��#Dh� �&��:vf�����t��B����6D�)ı�1�8�E1�P��(��w��\@�c��q�RQ�M4�o*i��ve��Wu8wi��8�x�ũ�������U�$BsAQON!%:#@YxN˘�ŤwB�i6�C�e5�f�.՘a RY�f�Ufe�����eH$B���P�v9�p�^8xVK ��F�d���J SN�L(��Vy�Fx�6u�y7KdN2�6�$Ċ4�blą�n�)�'��#'0'8H�(y �� 9B6�H&#!��N�0c-���X$4�8��A��;�4l�$2��$����	�����El�!�Xr"�P�2Hj$aȓI&�1���'(hd�!!(�I�0�d��� �!�Ł�4,�i�'p�E����0��4��.�T�)����e����2U2�F.a!{I�#Оcc̅�����-h��2�EM�Q@�"����Hu����ϊK�I^�7Լ0��D�Љ��MSj$bA"��U"cS*���ډ9��z{zR2�1�i�������b΢�*���n���.sQ�wx'�Ɓ7*7��n�\�}�K<}{��BHFOc(�I<�N��`#�8�a4�(�D �q:IP��v�ed&�PNE'9h��WB�M u5a؍�z�pcST$�jJ�n��!ō��T����Ŏba���-x�&:�XMb-�
�6E��<TQ��*�$���W��4�.��\o���鋝Y����mm�Ȇ��r���ɞJ����A*���H��- �b���B��8ư��RX����"�"�Z��@Q| &j��l��.V�ꭵ�m"�C��@�LG��])7��!#��A�xظL(�F�[����m�)L��l��R�-)`�����R�HV�E���}rD@jgj$7�x����;�v	&HD	���)fU^I&�W��J�r��!�u$��M�iY��dC��=O����>�K��q�1�Pn���/7�"��LR���W������^�AhQ����}:�	�2����$޸��|\�>\�Co����H$��l$"늰ƌ��n`c��(�#��(���#x.���Ά�i���� � ����Kiv��9dԒ��4�1(���v����T��F�RT޴{��]�%uqm��2�Fjr�SCZ���( �p�BJaV
�!�Vn��K�ۊ`��!o��ҝښ�u{3�K
1һ��8٘�v��.����l�6Db���p���/]��Y�h�!+�n-��6I����4sk��3]A���s͔�n��K�d��K�Vf�u��Bˁ�Y������E��}'a�:s�u��<}������Ϳ����3���[�?oV�m��m��m�ڮ�������������������z�j��j�����������u_UUUUUUUUUU�c�:�k�rʵ��Z�)�ی���Qk��N�����2[�,�����5Y`j��קs��;Q�9�6����V�
��CL�h�%�a����w:��U�UU�V�]U�:Z�@eZ���y7=�S���,�UUU})r�UUU@T��5R���P�J��J�U�S����V������eܛxV�@PT�UUUUUYF�n�vm��Z��U�������iIi��UKʵOh���ꪕej�4WP��[usϹN�K�M*�a��V�UR�G+�U+8�@����T�ҭ@]P,UUUR���R�R�U)9�ـ���j������[e
��f �x������3�V�R���mU�*�KuU:*����4�U�UTU@U�*�K�]zܙZ��
��Ғ�O]u� �KT��-U][U*�[Uj�f�
�V�eZ� -�l$�y,�4��I��hlP�UUUUl�����[Y�UT��m���!Yܺz�T@ ޻vfb:^��NS�CT��b	lnuS�v�jqhu�=<�ǁ���8�l�E �t�.3����W䍘m���,�@+�Li�V�e�;Z"���T]�)�a����h تXmL���P*��g]�=5u�UUJ��K���K:  ������M�H��9v�p�cT�UUP5fN��`�6iV��m4�Gbm�@ڕh8�� Ib%n���ն͌pv�� ,vIz�����s�T���uU]YYc`��T�\٪��k��Bw�j����TuPUmm!5UU��\�u�$v#�� ivB��V�V�uV�T�uѴKƺ�:�������������'�Tn�����a�k�u2�u�x�f��_�O�~$�[��?use��ƌy&R�tUU�]���T��T���i綂�����j��hv�{M�1�F-������j�֥&��.a
���m �{t����9����Tr�@*��UWr�-MSKJ�X�ٝl�ԙ9��*��]�����b�����݄!*�Ips�jKjP8�f����q�5 �φ6���]��cV<��� u X63$"�ݺ;MGD֌�6z���W+���j�k��B���T��֍��|��UU�[en�C��m���˸��ZڦŶ#-�`WBv� ��U�-�ۭs����mu[qT��`�ڼ@ږ;�)M�)��-�fp�۵���`��6]uWll��:��UUr�UUN�4C�,�U���UV�$*��]�-��LD�mM5�̅�pDsZ8T�
��[]Pl@T�U[S���ٓ	���n�t�;&wgz��j���%eZꪥZ��H6�T�Uӗ+�lln�v�4J�UUUr�[��n�'�Z�V������*"w)�k�qL��v�fPkki�5V�T�c9�7KV�A���m���i�+d��Elm���-u��e:�����R�Z�-ay�4Rv����`�j�)j��^j�����5Z��(�X)�/��UUJ�UUUUV�U[ �-T�m@t��N�����J�6�M�M`��M�x�F�8����ƩEkF8����);7����6�Hgٱn[���$�^��ЗcO}�z ~�\��kXDLt��������΍���UUUqtUmm��UUUt�T[vz�anw��W(�����^�q��\r-��NndЀ�3�j����*-e-�j�������Z�VuHUUr���FJy��*�09�V���͔���n��f�z�U�Vz�W��c��HB��h,�j�`#��c�EPz�+��ЗU<�=pVpv�$҇[���p�+uUUUv�*�nm5�l��{ti�Z�=rc��Y�=���1��=FmYj��Y�نhٻ�ss�ۇ�QAT�ˍ "(>1E�>d=��N>*~~�3331UUUUU*��������UUU   ����	�1%��az��az��c0�f ـ24#�4#B�ܮM��ܮx�献x�献x��3�+�2��+�2��+��
g�3���нZZ�b�8mհ�[հ�[>��?'���zV�N��5� �)c1�J5PPG�2���i(J)iJ����p���4'b<��|C���:]#�9�@M$�t�����H گ�	2.
@ɥZ70���mS��=2�w*��e:��¼s��`��E�&E18t���
����z��E�DJ��(�$:
_��&W�2�W(�G��4E�`G��0��S���ĳ�d��6e\	Z���� h�N �W�:���#�@ע�� �0��t &���`v'$���""��4�W�Z�&2��^���QQH�
gjZ��#��G��96l�d0�]�g��":�xvB09�xЉ�H/Uce!�;d��#�6�B�c&�a��ؼ�(� @B�D�I$0)��2�Ā��j(bҬG������VA2��u���R�6�ĠF;������2ȄȎb<�s��-I1�Y�AuJ]�'AN���1DPZ@69�F$��� �Z$0��+��H� ��lH��p�.M��%l�;���	jE:�ͨ���Nv�N�SG�z�C1%�X��X��0������ � ��0�)����d����ދ�USU+��B4�@�� �'XwY:;9����]�UJ�UJʦ^/X���q'<y�Mm;��Yi��g���&r2�&y�X�vY��g��2�a<�bJ��P7)�6(|����d����!*\�r6���jwm��xF{�4�h�8�\Ok̈́����*5�e�y3E��wlI�Ke�u�6��l�m�6��X�p+'S։-���= Z�1Y�G(����8M��5�r�p���Ľ�O+�8p�ښ7����=�zэW.�Nъ�Od����1��n�X&�����ٺ��
Giۮ��x�� Ktj�2�r�@���k�O\�7-�V��]YM������-ہ�QɷN�b�I;8x�8��b�ݵJ�=��
�!�`&A�H6�.�G.�IE^%�e�!�"02���dO�O*)�=<�s����<�c@��xqs
�x$ ޕ�⫘��Kgwb4�a���cmF�'[;n�a�xS�b�n}q� �&�4�`Y���fLmwAB����r��Ŋ��l��8�;��bzu�jN�e�}8�`ʳ:+RR˲]e�T$��F�z�.s_�s�_se/.�˿z��8�{����2�32��s�N��[��8���ϸIj,fB*�e�*j�2�r�����w�o��,�>1�`9�h��}�4J����2k.��_hM���̋��L@�;5�w����|�Up%v19i�Rd!."e�\�]G���k2�.�}Z<���I ���n��ܩ�5�v��8DKޛ�yϰ��g�
�Z����l��R�VbN�*-����{�~o�N�wfE�n�����݌�MÙ��ڃ0�˸ʄ�,ʬ�b����L%%1�J�+*��Tț`�V
w���2�[��l���]
V�_�v'��%;��y�;�d��((ݽ۹ ����Z��"w"���+]h!m�[*�#��hr+���V��c�ň�]nsV�D�C:$�l�I�s�̓D�ۢk��vm3e�!:����wMg]u*�vy.����p���U�����{�{���7���r�H�����ͭ�� �ֻ� �UYqm@����W��W>������u8�[0Bv[e��R�{w������c9�1A8X;FI�ܜ "Fr^�P��~��E��r�f<v�w3�[m��m�z��`L�P�����P�J˒�[��>��e���r�^�n�\�t�6�|A�|� w_EO�Ŀz�vӮ�T��4Ͽ^�Xo�~�����tu�3H��\`E%4������	�٫˼޾��f'��odd�HNJ�s.��(�(8P ;���\8{޾����s.C���+�M���e��!sZ̻w=�w���ӻ*f!�Ue��v��v�x�ȹˇ1195�w� »�q��ּ���.���b���ֆ8�����s,1���s��\	��^ڠ�d�tr)$��v�m����[��ත��D礧�j��`�~Ig1�̫U�ak��[Zr��dUPj���S���������W.,�U�xF�h���W>����jn��{��^��Y��w�߲��
�p����F8"��
�m��.�?$�s�o�{���P�`�:��Q"c�׵6��	����s3;�b�Q3�u����m�r�V]�$J�k�=0�X����Q�$�v�(+	���fd]d\�3n�Fg� ��Ǆľ�=��7m����k����O��M&�5I�</�^/�X�Œ�V*2	��k8�����)�H���%Y(�0Sr@�,�,ӳTc$��!���oӵ 2���uH JIDe�P�&��Y�`1f*�����$��%83C��f��1���00[�ܚ1&��7���_���5�@���d�� �m��`c�":á@
C��Gaa���CH�0?�hMqP]�= 0 	%  M�[��Gҥ,�kp������ L?y��ٔ0��\)�̸��:⃳9�Y4]YJ+��&y���3{�D��� �g��`�"v6�9
����AQ�;4za�^mQ;�X�/��� ��U"��H.�:QElD@��c���R&���� �I���2{j������w�)�����ۄ�Ct�Q��BKs1Bb]�fsސA#6'?�s��,"u���j&7=R��1^=�5>%�n�7�.ba�ظu�36��T�Ju�?�����v�� ��>��]6emu�u�L�I��%nv#K��&���h�C[Ve�|�A�P���P_Zx��u�Ovܾ`q.��i͂�lM���
��ţ�,�h,̪�fl�b������䂐�h��ST�r����{��� wg���p��f�� sY~��,��Z�?*�
�myʾg���d@}�o	��	�y�g�;��T�w�jIo�/��g���O��:�v�.:؝�9Y��X�*Mi2k3��{�%�7�SX�\�
���y��G��g��� �R�߹����r��_{��~@,=�s��D�ƒ]mR���A#v=�>�p��0E��z���n���֘5�V�.ph{6D�15R�����#�gu�[	�v���9�'-xlÑ4F�x� >"@|���% �`~�����w��6G~������乁1;`���g9��YԖm��O�v�%��JP��P"�!�.��-��}��T��bK�g�Qn�߆ ΂;�	��{�"V}��T_{{�:���UYyENDu�s
Q� �*x� ���*�"���}��Y�ڿ���s�G���C��うz�K��0�nLja�ǽ��%S.a���s*	2=�=�(q�����C��t" �~�1X�I�q��G:�;S '{���k���1��}� e>�I#3�V�"�;�V�;O1� }�|����⿃b�Ұ��Mv�r3���eV���]�/��`&��X����W ��kN���F�^���Ϟ���.�5ݮ;S\��ciݴfU�]ıO3ѹ��,m�Q(�-�����B'�bV�u^�K_�����s nv�:�7{�c$���G�b]���3����9��.R��O{[�ޤ�Oz�3�Ԯ�%�}ř��9�w���;������Uer���(=b�ūtj�T_ys)�{�N�o{c\�L��{� 0h"A��D�-?(n��	��� ����mȊ �W �	;��lp�k $wU� �Hw+o��` ;�q.rbĖ?{�;{�����	ʢ�U�I����e�ؒO�ճ{VY>�߽��"sæ[������wI3<����ֿ�S���)Ku_k�c�118 �'�5����T`s,�����������B|�F�,�F�8�
B��⩷"(�ê�����a��q�}9�q I3^�Kp#ޫ� ���S��\�D��u���?�(������
&?L��~�rW�}���{��|���C��P�6��vL���gB�>��s�.a8{�����{�x�bc������շ׍�L���Y�^�����^ja���@0/����^�"#&ffg���Π���<���XF�$c�G�<�G��o�'����M�P�/U� U����SVF �EP�a
�*7���E�>���eZ\8�a���0&@s,$���t��M%�޵��E`"T�yi��oĞ�%8�8 KXX��/e�g�k����8���Y+[���0�pSϤ��0tj�5Z�ەU{vL�:�<�ؕ�K:�:�9�^�cVNU{Tp2�[�����Pc��=�R6��� V]����dų�MN�� l����*�<�qǦ�@��o1�vہ��~�]��³a-��(v��j�vy�m�-���eJ�:j݃�@D�*l�<Y5�[�j��u��<����p��X�l�
�1т�5^웞x��N�s]�ջTP��89�U�X!�s[b�a�1�G�g�����������n��g��7^ّ��������z6F����2�H�x�¶G�9�Y��mU[*�8�K�uFpq����P$������\\ڊnڠ�p�R�zR�ě:3���rQ���"3O[.�x��ޜ�����񪪪������������������I8�?ɴI�q`Z=D(0`>��U�F�FD� :�qQ��K`l�8���t�x ����z�+VUQ�*�*�UV�+c���o�*}���)�Q�m�k�x�&�Ǯ�7$e��[A�;f�r��H[�{=�y�1��I�LE��*#!(EGUO�K�W���mt��C��ۙs8���& F`�����r?	��������}�8��L���_v�fu��>ٝۻ���Y,=�o��~��am���TQ�*�0N��&������y�����o�B���|E�>���n���g?��q{������W.bD�vd�|tut|&���k���N[��:7e)cb�W���Kn@��!n�^1K�����5m?�9��g�]7]!���.a8��b�V1��y��}�X;79��֩��]�q(gS�����6;H0>�m�4��zᗝ���^Mz5�lr�"��F���j��n��fi�{�vng��CW"�c=uꐭߥ9��)w=Y�yz��d�"rʕ)P���Oa��	�D����煘��x�4�����1�^��;����/������oOr������n�w>(Mt�c\�L#�3upwY��{޼n!���3C<�s�\�����m�7]����aȊ<��@�2{�Y�ޫ���lgQ�0���c
@�P���h�~�Lb�5��ݻd⨮����֣M�n��%3���uv�`x��V6�.1�P������u�ǛH%�-�q�
�蛨�����ĽVbF��f��h�dz�����{��"��?������~C���2�C���u��u��ғ��͡�W��k9t�%��T<��$�u��E�LL����H����y�[�ٷU,��J��y	� 2�$���3|��$�����礫*�=��@_������MG�1��I}��Kr"����r
����ƒ-ۏҜ�C�t ��7!�1��ϗ���/zg1o�u�{����[**���v"�m��94�|'�����cu��-�s(��y��=�{�4 ���^/#��fwG�#A�$� ��3��?���QqaP���1K�V�s�I�	��x
�{��? I���}Qc2�Kj����O؄DMKr#�!xǼ蒆�b�=Js=�]A�J��վ�=� �g�=�7%����z����M�HM�����zv��|� M�z}��׫ﱋ��ͥ��~��z/���mH�A:P�4�,���ѧKmy��]���gB?oU�����&��s_�@y�p>�4���eA�^}-Ȋ��o�b�+� R������{�×�vS���O�|n!�z����%]�B��%8rVT����t�']A��e�)���^�h^b-�ݮȽ7+�k�yrl��zj^[A�n�M�����.�e�M��/O���OW�s[�����c	v����?w�H_���f��\�N6ޏ�Db���mj>�@�����s(�5O��p��7�s"&����g��������m�����o�y�{�f(���x�X�F���j��p����<F�￷�Oz��)�5�b��y}����?D (�BBHĕ�U�E,(� �G����_DJ�����@vt�>#�%��y
S^��$*H���3�p �'oG�D���	)��6Y��u��U�*�����*�er�. 3.�L�DY�]1��J�o��KJ<��������Ē�,������zf����m��0��i]B�pdtx��՘�Ĉ@�:���E���_eX� ����%��D��KXc��
ᆪ�iB����Y)�-�	(�ʕd�4�`��9D�'s��3���N�/v�*�!�M�Y&�wa��3�ojp�x����@6�|.v�f����	L4 ���4�(�� %��]�l�L@lP ����s����[�t,\�6S�X�~�[B\��pV�a��/˼��9��L{.5{�(%�i+��bBt=�b��s�lh�S��;����>a�A��ߥL8[c���s�������}F?V�+�\~��,K\��xq:���K]�"����TD0�9o 	�Rn����g� ��녌7@��ͣܘ�؀�ng��!
<�[�%�3�ĩ}�nbн�2���7�x�b�L��m�[���(� �}�w�|T������V8�&�-u�i {[p��!'X|GOl���s<����#Q�91�e���W;����k:�L������g%4(Tqd����!�O����&�ܼtY��\]pU��L����'�[�?�g���wۏ8L�E�Y����b�s����9�R�#��V1��@��3������B��f��G1��a�N�t1�y�Es;�5���}G.5`�GSrG��:�-�Q�Y��]���Oӽ�SU�ؘ����� ySǀ�� �	���{�8�m�{�p�s���!�lAGu��z>
 ^�>*|�#~b���<�3y�7_!��� ���k��6�M1�Д֯΃����>�l�� �����B���[y�u+���T��ܷP���>@@ N�9Y�1�^�r"��r�w:H��*{�Ks�8e���Σ����Tr���|g�L�����`q,w13[-�x ���!���V�>�y�f"(�3O�H��;�o��ndL�w�^��c�((���$b{5�(v��4�������������,�uDܒ�)@���tӀ��3H�~$G�s;ۿKH�>^ y��Ǽ�o
�O�ҥ�Hw1�pWt
Z��|�TKT>$�$i���3�kA��1Z�|>
&O�ǈ�}�;��O� ���>J���^%�4UK1����5�;p�^��F�ļq������4�q�m�we��L�ZA�3�U�+�aM�6ϝiC���ajݱ�<�;vm��َ����䑡��H�M�$��Ң�]@ҭM{?�7�@��� ��ǽ�N�33��.�!�ί��^��n!*����<�k���|�$��ͣ�p> ���C{7�nDQ�����U�Ý���l��PfZ[R�J�@r��n\��.%�y������@�'�����D�X����H� ����Bz ��8O6����ш$z_-�tW�\D��Y?t+������	����{����.bY��"���z#�'�Ǟc�.f��F�Ɔՙ�eh]��=O������Ƚ�u��jg�������!���U���x��_��r�2'T�����.K�G�&% �����y�	��\��4�ٛ�μ�&$��찴���Zv�7@h��ia\$�R������Ig�;����#��G��X�Lw?!�> ��Ƨ33���c	^���?w��p�޷[��5�-S`��_#@|p�!��1���_�(I������5{�N3{��ׇ���j-vM�iN�`�%OY��]��r*��?+󽃺gu�+_!]y�D�C�x�6y�>����A��!��s�-
��*S�k.���3���y{_�� 5m�!^���'��p��u|F2$���1�4�
L�f�Rr�L� �
PG@��C����C:X.А	�K�*�f�%����U��Vl�J���*%�f�/e��~���cH�Y�7�5���2 ���(���=I�hvY�H�^���(�ocΩ�yB��j���j��U���u�n�a�8L�m�ZT��{tlm��(�4����:�%��,��F�'��Z -Qءsg�$�X0Z�%ݜ<��X9U&�s��1�8̃�]��e�ۨ{s�����>]��n"k�-�W.�<��q����1�����[�ű�N/N�ɷYм�A*�rFG ��YWT���5rX��⸠L��k��[678�vC��Ț'�[�L�6;\����s��\=�㓥�<tKs;�8�/:���rc�t&��!7�ml� ɞP�ΑY�����+�����0�C>�p�J3g3�D����b�ֳ��[k����Ĺ4�Z��E2�!�m�9��0GB����ɐ��Wu	�n5�gf�{�0�e�R�-�a�ذ�Z�ٽ�����>�0�FLE�y� �N�6y��Rh'>Jy	���N������D�з�?�1��xN�E�)T*���[��)�{O��5t��<�7m[u	�"XMAB���
;Ƃ�4s�3A��;:-��٧5nF%������.�y�m�&��@ ����F[S
"e9�3�lb�)0y޼M�T;��gQ̘�o�Bp%���ͣ�1���_�܈� �ձ���e�����7�}�y��<ۗ!�s(9�;�H��v�Wg7G����^��}*�p���*��c9���~��O��Cȯߠ}O�q�J[�kQ�t���c:�[�*a�&��;��}�V������μ�"�W���Z۵�� WnKZ-�N�:Y[��L��y��g�/y��vKE ׯ �3�ĩz#�.�(�h��p�������o���%ଝ���?.C�w1��q�}�>+�cvg�/o��[ac��� V�d�-u��]E�O5����.B�y�?�U���<�����Sp��x�B������ObcYς���O�G�Q�"�A�����<G��K��~�*�^^�����FfW?����*�2�[�k���ݚw����o|��>���\&$E�мgQ�z
�l7*=��b>��Ƕ�p�r���.F�1����c���ba�<$����<��s?�Y�ͼX�w��u�8�Tm�o
]�����nݲ%ڑ0����pj뒩.n�K`v����9�u��d�3x�h�u�mn�1�,ca�X[]���f�Znɢ�E+����rr:��N[$����[�<���s?��zg��Z=��k��=y�܈���7��yZ�}O�p ;��c�{�y�"DE�g:�c���{k�m�e����j�n!�!�\EJi�y�X����1>��T�����ҝB��]�������3�f�^*ay��{���~޼m�*I���1��x�=F>�߮\�=D��/�ot��o}�!���5am��G���+��-�Un��{���L�fu,�B?WZr����X�s:���|��$:��d~����B�?��~�>�X��︺�oݦ��c1����\�GQ����݁��PVZ{�o:��BN��L#���;��ٵm�(T7Y�x����@1^�D�$�!��#� �c7Y}-�QGQ�cu�vH�@� ���b���ܣ��x��������QL7!�B��+�3 �vD��K$4��γ+W.�>�C��M��{��3��s1>Z�a�GW��c���{�8��C��3[���}g�T�F��u.�4}�5�7�=���>��	�o뺪1*b�L\A�i��*j���u����l����Rfn|��"�:�4q%v�o3��n�ێ،%ƞ�/�"$J��]6�܉�Y�Г��wi�3xa�B����`�2�18I�������n���ߥ�GPJ���s�8"<%�;�M���#<5ː�n��Mǐ�8����t8~�g�f��c=������67lh���5�(���Q����9��鶻ؾ��R�;��FITPD�T>EN��{�vߐŉ)�\cB"�c� ���3��9p���m�7Y���nQ�~o����߼-'�ß�i��٥������AJ�`�]�<��\��~Fu�����\It/�!��!�w?��D?�7&}��5���3����'   ��@V�\a�r��P� �3,���n�m	�XM����a��o��	$#1��C8?�wz4i�C2�%�D0�"�c6܎��h�����É.M�h�f���ծ9���z�Z@�� ���/�k7�'�by�@�[o��!P������m��	��yS�<�K4KHI�)�3������3BR�p0AYa?'�N���ߘ��l{��Oh�� y���p	���!���	�G*�J�������Z��;G7O�Χkض��/#�Ǽ��?mܧ�t��8����p��V2XJ�vȇT�q�ĵP�f��ZICu�
��D�I��i��c79}-��:�[��1
pGJ�(�&���f�� ��e� �����v�Gz�>�gL^�ߩ���v?>2��}9����`۝@��6�ǈ4K�i���!h%�1��mypj%:;��]�i�{#LK�}�.��~CQ�����w3V�C��C������K�����=��r��-���%y���$y-n"MEm��"��d�.�L��ޠ��v;\۶Np^T�n8*
�QNzmI��#�Js=���ks��n�&��9]{�y��,Igش���!l��7+ *����X�r����n/�<�u�U�>J$J/{�����*6sZ��7Y����	V��>�>La�/�g���f2�k�-��02��!��7��~Y�X.���gt�zҖ��z-�g{�ؒW<��_�ƈ�Oz�Q�%E�GV�-��c�(B��W��P�9���{�w3�������<�X���b��bng{��7���ۑ�씱 �CV�aeA[t��+��������3�9ȼ�V��6-n�!��?.�g�WLLCty�f���0ncY�c�j���G���}ݒu�uħ	P�g�C��9F~?NA)z�d����Nn�gP�$��f����u��{���:�su����� �B=�M���#>׊�T�����捽н��d�;8ĮΖ��l�X�Z=�n����+R�K������Zx�{Se�c�!VƏz!�>�BX�L�!�����dX~�W��1#}�5lR�9�#�С&{�J��c��Cs;f&$M�:���{���0	����>�m��i��J @�P��tx�m�$�õ�WR�����F������i�m��c%+��鶗]u�r���Wm�+�޶\B��I#'�o<�6lJ�l4.�
0�1Ì����k��Ws?~Q~}yy����C���u�� !���Cg�1�}�7S3?-�N[��r[�F?#�1���\�(�ދz��L��W� |�6	�8�@�2�d,)`��{�|�c�V�=\�ܹ)�j* �y�#>��v��e����� � ?y�y�R�|%K�C����jk�*bb+s�Y�{���Q��0�S�.�3�'�0k�]�~����>��	����A�Fm��s.4 ��\LL#|��؎&AX�� q?"e<�wx�1���x��d�<��y�/�4L50wY�wX�!9����Uۓ#uc eN�á�faLG��c���!K��!�G�|Ay���>F:sҦ&"��9l�9��W�LHL�A
[�U�A{�w�P��<9d�u��[]��__n+��Z'.o+X8���{�oS;�av���ؖ�:�.��B�#��3�?	����m���=�s��\��^G1��<@��T�?���16�-��6}����HD�^<}�L��Zր��Z �ٙ3iFO��?�ߔ&s="H&	S������N6{�$;��L`#�B6k��M³C(CI#7��T���,��j@��wq�w!
B�63%)�@9A��!�Ƭ�A�!-��L0�"Ϧ3��0��0�7i��Xv��>��Z�����UU1������ж̓!�J�g{kInJٝ���f��� ��epWB��Q�2�YK��"T��7����D��`�ɶ.1r�
�eÑ4Yp@bs��7 ٵ�MV�m��ӫ��ٰ�m�.��^���!�r��r&t��Z��T�K]��B�[i$S��wc�)-�ӃY펴d��5Nwj�NV�N:H�h(6�p�-����n�gv����p���q8����ν�;R;��ƕ�pp����ȷh����+=����cƁў,L>8���'
�+XW�2�n$��Qu�Ä{\@�d���v=��(�J\�U�󲚴v{���pګ�#�Bqjࠇ�3l�]z:+)���$Ln���n��cCv����f�c��-�Rpp7nћ�������Q�T��)���4�޸�*tO Iz#�^�B����p�k`&����  $8 'i�P�8R��p�w����ft����mI�T"c D&it�Xk�WS��W<v���䣆��ss�z�Q�I�K�J�k���Y(�ʥ���:��X������pv�:�#^v�m��7U���3)ʘ��������/�]��g�L�L���;�f33�͆�9��
��]��;��������>�L�1� -FfwbS��n����3��^�\��s�im��e����B�A�(�Z��}3O=�$�����︬K//eb=�+�b�w3��J��!���;�|����JU%��L��^�BK9;��
�����B�5{�w3�W1�*�*\�ܪ'TR�P��e �=g�]E��x!��g�"v"&\#�16��g��u䫹Y;�s���"q<#�Q�i�y�%[Vq��:�̉�P�A;۱$D�Z�Jŗ��E'e	"\J���\A;۵$D��.	 �0L�~�h0[�7��`�n�JJY��b�L� �'{IpIޮĐI���$�NJA$Ls>���U�5�N��~D�A$N���	=(I�;�K��POW��.�J2$�H��%�$h���H��%�$��A$Lgӝ��J�j	 ����Iz��$�w�bH�@6�G �������i�$�{�Ǯ���f�����1�M��I�1���	9(I�0s��x���0�u ϫ�g��eJ��>�~7$�w�q�$D�).	 �҄�.%D�i.	 �}�q*ʼ�1BTN����	1(I�;�K�H�9v'��݉"V��ŗ��A'�	 �&�IpI��đI���$�	��>��2$�H���$z�A$N�����k���*	"|��b�YMA$޻RA$nR\A'e	 �'9IpI�+�p~�͔��U��t!s�-���u�c�m�ƀ�G\�"���#p�Z�F⎰���p(���R��KF,��t�Y]6���v̲�����_?��sv��;[(L*sy����^�b�����I�=�K�H'9v$�H�ϧ;x��YMA$RvR��D��.	 ��ؒ	"w���@�PO��9ux��Ȓ	"{ԗ�L��I��{ԗ�I�JH$�����ĹYMA$��A$Ml��$�N�A$Nr���	=�v�W��"H����\E��nP�	"{�Zb	 ���kx�����:C����D�,�-륬0�e���:�}��H��%�$޻����IpI�羐��2$�H�}).�E����BX@�\�A$On��	9(I�1���r�w��A;۱$D��.�*	=(I�:v���)��%��/"H$��R\A&�	 �'{IpI�.ĐI�s�R�/)���N�A$M���	ޗbH$��R\A�?��[nUn��+a(�����sux��В	"{ԗ�.&w�A$Oz���	3ʱ$D绾UK�.������nĐIy��$�N�A$Nr���	=�vb��^D�I���$�MJF.U�*$�ٙ܀�	��y���K�MP��,I�9�s��`�SQ1���A$M���	�ݧ"TD��\A8�ԣ�8�L� �'{).	"�:�,I�=�K�6�k��6�7��}�E%,��9rؤ�5],��T�X��&�.�)�9�K�H'j��I���$�n���VD�I���E�� ����К�H�ϧ;uX��MA$�BH���R\A;۱$D�).	 ��q���K�� �'{IpI٫�$D�i.	 q ��l(
y09�jĐI9߻Ux��SPI�ĐI\��$�N�A$Nr���	��3�oc�6b� k��-50��K���q��\A&uV$�H��%�$<�0$�H����]���A'�	 �&�IpI��ĐI���$�c3���s"H$���\A3��$D�i.	 ��$D�9��w�����|$C�ŉ �'yIpI��$�yVTOz���	���%�$�� �'�IpI��$�H��%�$��A$L����]�y��ݠv��t��:��\�e4�{s�f�<	�N0���mĜ��@��.�QD�-�ۆ�Eٻj�M1]mD��)�]�;��;��t,�C�-�f�u��RΟ.�]T���A&�BH$��R\b��qa���'{IpI�|�,��x�dI�=�K�H&uv$�H��%�$rP� 
�$N}�p�x���5�N�]� �&�Ip��$��$D�i.	 �Wu�u/"H?@��}Iq=����Q*	"b�i�$�w�bH$����.��j	 ����I[��$�w�ct�>=):��{��E�������
��3SLy:�D�i.	 ��ؒ	"w���I�BH$�x童�*�H'{v�P����.��'����	1(I�=�K�H'k��*�R�$�H��%�$jP�>D�Q=�K�H'{v$�H�Χ;uX���O��BH$���K�H'�v$�H��1�O����b�dI�;�K�H&�v$�H��%�$rP�	"|.������]�`�TEPe�F��U��+I�$�{�bH$����I�BH$��v�I����*�^D�5�{ԗ��+r��I�dB$Et��
`D��n��e��!D@  ��ى\Q>4�L�&�Ma}AD��!>	VJB�n%]�*iŔY�`#Fy�;M��[�BDhT�@�@���A�I�#q�H0z==oi�n�#�U%4P������TB�I����T����r·8os1��Sd�!�&5P��������|%��������W�gH� dw�䀝�{`0R�+{�;��+G11E���+�gq��D�����Σ�ǣ���64η`e�n��Km2K���KL�H�H��ܧT����c���� ��DL8G���1w3��Nۈ�n��5��Oq$PWs���##^��<�b7�5�q8/�5Z]6*��3��ۡ��wü��lc���!�A� �zϼ�#��H����|�w^�N���y�G���bGۭ�n��t��9�Y��b�����N�*`�	��i�Xfˊu�۷a �Y\�3����I�7��e���+w���6�vvE󵮗���p��Td����m����K䖖��W-�r��o	P ��+B�7�[�Ͼ�Ǜ���2���H�Icu�G��.�N�Ak4����g��B��C����1�������C��+����<fr�6� ܻ����Ƽg���'2�8݃XίH� o1���8���� xR-�Z�B�f"!�:����1�p�"T(x.�2��gQ�����s$��fss:�k�?�v�"q�%��J���e��`��K���3[�K�Ty|�c���4ޏ��q�h�h�PN/ ��H���8�ߩ�D9�C�f���1�+�j$6wY���\�L���Q2��.:�uPpiK�PH`DJmJty��s9�}�9a�;�M���.C=}��DÚ��3��嵰��
��8�s��b�4(��GQ�cu��>���p�a(ZD2�ڛN��}�Y&�ZECϾb��A�f5�h��7Y�gQ�c1��Ben��wX�fE�Z0'GQ�c�tB�����b&#�1�VA�L�0I�!(Ht��?$�N�߅Va3��]�]ֱ�qgK;v�y��K,6�T����*�m��b+���MG	�떻k������zl�:�4��5�eq�\w��8�� �\��7
�������j�������|Ӏ�!��#��c�Y:�*:�[�w3�ĩ{�LG���wY�b3�\9n��5��9�@��3�M��v.B8֘�n������=�n�#<�����_0
 ��0;�c�V"&#���;�5��N�8nR���5�Gu�k�i�
�4���� 
��0�Hm��XB�������N�jj��y�}6�S��T<�b���t�<��:�WU���;�b*��#D��0��Q*�D����[��>��G9Z�*�&}ꂑ�c�N��\47G����-�׽���[�\���u'$A@���{���L���]�W�jfų��?/k�i�p{��{��g�޸Cre�s�9<�t�])�O@ԫ��ߘ�gu�#;�TL���v�xM��}j��.X~��Y�gW��n��N&���-���������F�:u���%4wX�gu�F�����:�ݳ��0��ǲI�   F�o2\�_�I���H�J�$�؂H�V�+@�P�*D5z�?m���+&ՠ������0��>CK��Ґ"
B%�'
������{p��U"��T�����"ʟ�
�CΓ�'����aYKƣ�9���7m������TUV�UUT���]�pv�֔�X��fZ�v��T	%�aWn�YC�Xr�Q(���
кy]��r��.�b��#���@Ye&@� �m��V��|�v�ٝ7E���y�d��5+3�S]�7-��`��]�i�
�@v�6L��Z� ;����	��\ǳ8�.����GeX�sL�z�2�v��=����B�Y�tS�1���9�9�$v!�v5�{�p�G:�[Gy����&yzEwm�:^�R�T#�Bݻbv)��m�i��p\q��]HO#�V�]#����{s�;i�@HG���`�ڒ��+���s�݅k�'g���v4���7��C�E��:�I�4��ջ@5K��sv�T,�\N�2�71�
u�����ъ:��@KGca����a�Z�>Tȋ��;A��)4�����]��g�ҁ���*E��(ؓ��{�}�>�֩�����u�ճi��LQt�(����/��c�z��/e9[�9�0�����`.j̤�����^���8;V���ɞ�%v���-��SK$u�B"��-��k�y�b�&z�}NbF���o��IV�	P�#�Ŋg��B�V�֢S���c:�c1�T������.reW|��m���22��J7�J�	�U%חQw�9�w��*��.����R�@.(h
���P3\�*�6��Jw�&ˡ��Xg��c�ka8� ��m�7Y���Ja�:�[��1 ϣ\J��Hl*J&7̲�9*��!<�bޙ�g��z�Jt7_�%�#����C���˼O�A�d�9 �d��0':��O�&��7Ln�s%�.\���LU���#����f̷:`l;J�-�x�P�V�/��ǽ[:�c=��[���H�e^�3
��V��9�����B;�]3��� %�!<��ɌGZ���W1W���;�����{��9�ͅ�n�&���P���IĴ��6���07Y��8&����lw3����pܹM�.��g�V�8�P��n��o&e���iv��>�1�"����v^	�m�eCJ�t�T␣�1[�8�o��7[fI��	p[i���]ε>�V�ӊm��\X]T]5K�l��n:y���g��� �\P�7j!a�j��g03��Ȅw_�c=�PJ��&��>%E�?+�|����	Ĵ����vX������tx#t��9�}����L@��*&h��%˔��b���W+���t;���< 8�$s2�s>���(���<��5r;W�d�ty�3Y�fg�UBg{�8�ޙ�Z��G��K��	f�\pnaC)��7W����{{�sŕ�D)��i�3�����T9�Y�5X+�6dr빦�E��.[����gu�k;�툈��PΘng^s�6��ە[h	��0�
9���FB��fi�{��.�g7���P����cϐ[�8w���{��g����3�|"&!P��z�<�t�H$���&!�H��@�&�y�]_�Cg��#��c=U�?1]�h��v�`�謜��tu�7Y�b3�\�.�b���q�ۇ*(n�vΣ��s�i�ptk4�� �9w�zT'_!�|#v���Z��Y��sr~�\������U@)э	g��F�j��w����{��I���D)=e,5���L���^b:WWk�\jn[���ў�
�U(�gQb��C��j�Q�E�C--W"r�Du��U�U��ҿ��?���@A�bw����C�� �6��q��q�����8�c0/���F��f���r�`�]L�fm��-�{���H�7+(�r!B�B ZB��u扝yHo9Ɯ�1� � ��G��o����� ���#Hw1�1�[��B.B��>+Q��'���C�� ��<�����ٺ�\������Z�q!9����6�� ��27^��TyCu��"��-7.��U���6�    �RM'���-�<���
��D�"li�]�R%ⴊH���$(��l�6�v��AX�cd&��0���L,0����$0K#f�4����6F���o�6ŕ� �	�D��B���nI]$7e/yƃ��v�a#��F��I�g�����7؛'m��ސbV!Y����c��|%R�v��n��pl�#!	�Ä�W��C��*Rm�2`��� /�0�iL�>���2���v�!� gϭ�-A�f��*��ꟕRk�0,�Vхܵ����T::�!��I�3��GP��c59�"]�gԐ�)\�Nf���幎��v�rR40�vi��gP���tu��k9���*�Q�U�\Vu��bι{a*[��B���'��1�L�ϐ��G�3��R�΃h����J\������z�&\GP�a��m0��G�"�%Odٔ�Ȗ�D�</[P�m�lj��"��b�b޺yb z�'1�B�6��ZM�M�s8g�sC��\vv�r���t-��7 ��Q��,\K3�K5���_��N��v/P�>9�j��r"%�38�/3��[�ܩM��iB��$�����tsY�:Y�bo�.[��L�1�X�z�D˫]��Gz;��aj�ˬz�s(.P���P�Qۖ��3H�a����J�G5�>TژS�{�{�9�ޱ���^i�fш�?�B�Cu��uB������_c�ε�L��,����֖�`�@I�����Ka������Gz'��!]�W���8�S9��7�Qn"D����Ö	i!��	��{yy6t! 3�Gp�+٪��ʸw�7B��`])E����@���b~��2�6;Y�O=�v]��UCЎ!�g�q��;%���t#�T;��9��8�ۤ$=��ĸ����(� �3�ќz�x*�WE՘�[3��Ǟ����c�֜��DUS,�7J�-�]��ɝy���9��/ �0����o���R�>F��^�i�3닕"P� �U���`Z�皣��+'{O�5oc�F��LEg+};l���Ү�!T���p݃]C�2�J����.=���qeB��Qq�M�ͅ-��mtu+�c�\�j<ېsz�"(q
c:�����q�:���Y�-��hk��X�k�T���3\�#�U����BtuCu���U�b2[�B��ͣޝ�2�n�8Σz���m�P�V�5�L��b�i>�D$����VUU�)$p��lT�l�y���oqo���Eq�?�����}�X0<�oT~��E��~�n��ΣhT;�g03H�1���}m���s�g5�	�篦�j�k��T@�R�Sg8��L�.�*��f���m�L����j8��ڈ����H` h^ {�@:��/����P�#Hn��Ϯ9]�]L�&m�r�_����F:� ���'q�K'��,�8��Zz�Ϟq���K@�rf�q��6���N���hnݻ�w-ˏ�{�@��! ,��>_N��Dˏm��g���2\�����G\��$����m�]ק�LK��ٗ�ە0#*�.�/��D���o���;���aﺯc3������DתJ�j�T1�`�*�����}� �)�g:֓��8�>��!����B
H��qQA� uL��@D�[���E@� ��E�b����a�aD�D�Cb�jCP�� ԌN"$�Ċ`J�@re�^����#�1y	0P��b` �8�!H�(
w�C`0K�"��w ���xE		^�B�~$��4�����P��������~���PO�Q?��'��	���T���E�(��q ��@�"��;���t�k�@�?�PKo��
���~?�@�UUUUUUUUUUUUUUT�UTP��PNA�ߗ����{��X9�CGM�$6�%��(��f7�P���ϙ��?����O�����?X���s��#�O��v|��ɉ��r��P�}��|M�������~$	BP�0D�%}ʠ�=�����:C��Hy\�����?���CSS��W��?GO�Si�z�y�=����$x�ޙ�����=���(�2#�%*-( �
P�
R��*���(�*�J�P�H4�*�B"�4� )B�*�B��"!J�-B�4��)C89�,&���H***�b�bJ�T�P�(�
�Ji��$�iV�F� �	IM%@PD��H$@)�AE)EM%MIL�K+��@Ҥ�ts�D�#��}�Hy�o-��:��,���|?�S����J ��|��>��|��B���C�v����p?��>�?�H�o���l�O`{BU����t&վ������e=�m�Oi��b������6>!����8�>��������a����A@};�!�=<���������v<�g럁�0��PjB�(�>��(G�p�|K׃���]�u�|J}jw���񨎣�#�����ET��zy�&�rk��P��DP����a�p�����o@�W#郩Ȩ(�>���O0�
����@{���� �����P���C�5� v+��Xd{^���J�����o�}Pب(�W�+�>��
����P����g��u�xw��G����r�ppHlBO�zf$�]��~n=�������a?F���8:zǠ�(�g_5;����#ԇ�H3��W���5�Dz@*i>Z�`l8��������x�! Pɀ�A���P=a_Z�'��zv� E���3H|��ó�9q}:F����>���P�*vk�z�rE8P���s#