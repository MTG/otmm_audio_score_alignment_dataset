BZh91AY&SY���
�_�px����0����a��    ��   �P(  P � hU  )��� 4  "P 4�     � P>}�0� *  UDBT�*E
!"� B�QJU QD�B!*��DT	(	 �T��HP�w���    &� P      sx����>�=ts��� s9w��D��=71ܼ� ���Ӽ�à�H8��bj�, %a�ӛCNv���3jW�p �a��@���:�i���M��
���w�    ���-�����s۫ͯ{�^���U� W��\�����t��]�j�[�J������T�w˶�yj��!�xں��]ʗ� =ꕛw�R����W�J�}��M� y�W;+�׭9e{��z����Wπ      P����|%��Z\���K�ruU� >����������ŧ s���W�� �>}R�����ipE'�.��4�rt�{�>}*��}��Mu��k���^�_y�ͪU�Z�����^Uw�U
�{�    �  �u :y��3���*��u=�N���r�s���ŧ6��U�*����K>��|��G�@Pa��R�����>�}>}*��ʹۧ�O6��{�Ҫ��ܩY�C|a����v�8  >�    @  �� y�,��w�.�qer��T� }���vҹ�}iɥ�qd;��O�J����w��x���7W�J��ZU� <����w֪��u��6��ܲ�� 
wJVm�jrgf�4���3J�           ����R��!��4�24�Ja"jQR��      "x�UEQ��i��F�0�2a��R���d      ��!�)QF# @a �L��B�5%�&
m0�F�hzI���)��S��?S�~������6�����}׿�����j��QWB ��~�EQW�Up	D�������U�
�������:�E]�_�v  �}�?h����O�C����#�BrW�rC� � <��'$9 r䜐C�J' �� �/!�/$��ܩ�M����' �(r 䜔9 Jr�*rPy ��Hr䜅9r��E�<���'���y �Aܡ����!����$H�U�$9��<��<�@�������9��	�y(�S� Q�
r^H��H��5(�MB��<�^J>�r����ry!����<�@/ ^O$��@�rT�'!������Qy��<�9 y �9 �]I���y<�9' y!�S����	�N@�� y �P����� @����'$��������%_y��7(� �.�y ryr�������#��$K����W��@�@��y
�W��NB%@r@�$�!^O$^@��9r���^JrG��9	� � y�C�@�^Hr���9(�C�%9*���H�y ��'%9$J��9� ��C�<���G�<�9#�y
��$9�NB��9�����+������ �rT��G������./vl��eL�{�n[�<4�B��������f��3�!��X����W4x�1,��BjAܹt��k� ��(L�s)�k�s��6@�yr�����&1��~��{>ij/�v�dH�}@�5����hJ�u��[�܆���I����甿�J�����U6�2��Bn%���.*�w;�č�t�	1�[^���6�=�ܨ�On�
���������R�z�vy� �@�:��3���3���8c��|(�h��C��rq4�#�M{�
�s�uc[04Cx��ܢXɊ�u���,�PI��^f�Y{���s2"�_����˓u'�oaM:5k�b�y�Hצʱ|�]-ݚy�,q�����)�^7�_(\O5��3Y�{��͈":�C�W����&p�8��Z�Q<Z� �1��>�����ϩϙ��/8�}�s��r,�j���2c@�g��ӟr�HQ_�����h�Q�a��Y��;�r�6�>Z�^a^<R��`8�b�!�X�q�	�.�ѡ���C��;�3�{@M<��J��r'!�#�HK,K�#�s�;���e��f��FAIqK�I�y����]�n�'a{״Ir{���K�{��q���S�jQj"���W.+P�79tHH��&'���dx���k#$HM¬J2���0#,L,޾>o¾d�&ww�}��H�a��I_'m�Մ�� �!��WZ�5��,_u�ݜЗ-ʱR&v�5a��P�c�,�zgv��h��Ɣʤ ��!r�,!��8��ƐR��K�ϟ--��w��mC����l�<�,c��'+@����[�W��� ��'���x�w=��s�5ҵO���Bϧa�x��>�Hs�a."@���e���XI���(K|��g��q���Jnt&���w�V��2]}0�"r�}�5#�ōcX�s�}O�тf	12�mwv��ҏ���UB�u�p��(�;q\�,���E��V�F��)�1k��9������sF��}S���p�������f�G�NM��c�I��{���NY�/7�S#���{��v�<"B��c�/#LG�5�~DQ���y1�g�!���6F3Kt�4�S�˚����#�x��9�d���.c$o�b���h!�9��ͺ<�q�nsJk!s��~P+.�F��<��:"TqZ&��yĩ�sT>BYF�"��ӨpxJ�b��qjm����(S��L��g���˿>1ۉ����1���Rr���`��)8v8�|.��r%�j�9�ͿԧӜX�Q��u�W�^���I�&U�(jN�AT�bH�ph�G�ޒ��ތ5T0��l�X�5�K}�sr7��Ac$ē�C&!��@��1:�1��N��ޮ�!UD:	ҹq;��b��I8}��Q�lB]��Q8�D�&(�&C@�=�d�rм��=���Kӂ�y4i߻�mK�j�&U��f�s:�VJ�[�gt��̔A�0�U��þ�u��|����,}T�N�9���Cp�����!��$���1�g��4ֵ\�_ib76_������G;��r8�k���Ge�ѧ]\)u�1>_�-���5H�s֬IKB���^V�yxy���b<��^>\�z|�<Č_ p�C&'j�MF��KE�w�{���Ϡ���o.�;ý��EdD$�hoߪr��5K��l�����r�gW꽴[��|u<�7������}[t��fR,��>""6P�Ԧ-�w���;�L�"�w�154@h��P�3���H訪y�taD�����Ո_��|s$�7�1]��TX�,����!%�'�uW�4氂��y�,i�	P<������,pȇ(�v�dS���',����M=���4|�#
�$D��!�I�WW/wg8f����I2=�#�c0X�<I����*�`�qTJ�:��n�:�C9�g���#{�@�A>|;�����C�ESz�|�*M�;�܉�RΩ:,��@�ǭw�Z��i��=kj�ru`,F�2�ġiฆ��y��d��g{�;�^z���w�6�
��o�>I�qN��I̺ty��B�iB��Q YV8:T�Z�*#��4�PC֮���lv���C�y�k��;��o��{�B������~�t�<�2-�������o1�S�%S�~���x7�������8�XQ|���U7-��.�E����e������k����:�����A	|�ӣ$��C��>ιN��ESr^�]X�����q}���}�*(�
]���ōP�r�b�(���E�J#lя_{�L�r_s��F��.���#��h¢��o�h�x��=�p�wrJҕ;�9�O+>��$	�ț_/�|ڊ�9�o˝���P҂x$�T�La�����#&��8,��i7�;��n���>��9uI�����a�tMoF�6'���
���}��p^��?�W�Wbx�w��n�'ly�N.�;ۦ�&'8�
$"wMv�j�>�"����
�3����7�y1������{}H�I�	R��C*K3��_{�Կ��C(d�$()�>�R�x�
�8�Y\b��I>w���8]���K��qSȷ�\Ns���c14�p�j�>�X���j�`�z�f�2�q�h��iO2�Z/eg19Ճ��ɘ�'pd�I^"Q�2"ޣ��ɼb^�S���:S�G�%r�$��o��߄WK��z��Fv��L}�q~rw��w�����Co����f]��	���!q�X\���7{��ݏ��W�Nw���K��q�z
no� ��Եn1�B���T<P��CD-�q}÷Nwyɏ���q���Ic��u��9�~���!�>m�~�Μ;�9󇤖����{�[�k�:�sq%���F���0���h�@����f2�&t�	H���Ή�.��=O1v}��$cȁ�4��� ����n���ѷ��+9���7߾�|#���9�K1-���ދSӢ�yv{���P����\����J�7@��tF�hr����Z'
�>C%¡�N�Ɠ��Ŵ�T��7ӕ��A2!�6N�I��L��k�O5A �㉛�i�L)9-eY�螂�c���btFXd��S�4dӼR�g��3��l1&����,a�A�'˃52��#��E���Xukio~��������O"��qb/��S�sx|5V5ʰd+@����y�,Wx'n�5�(��9���g>�&�%8�������u�t��	����7�A_�;�ճ�	`G����l�JR:��Ϲ��_��q������e�%7�*��#�$���9�ʱ��Y_�!&��S�y߄9���ע��U�������UY���y@X4c)�(2,�>���&0F�0��t�(�N�T�E�(�E�u�5#���g�E�x��}�.)�Lx=R�"s����X�7q绦�l�b�i���T�qsn
bIA!���RP�gW��S�z�;3A�A�h�e:`�K���Z!'1���gE������3F=���p ��L#��0��BǍ ����i�U�.C	�q���f1�BQ�d�	�C���Mj6d��BY��@�����yޣs]�_B��V���q&���4�cc�o�y%_$��{��W1 C���O ��7H�LY������XK�X�5P'�`|����v&mˢBd���Cr�d�,��>Uƺ	,���b)~�/�|u�P�"�,I��n藮�۸��ٻ�\bqwD�|�Nd��&�'*h�b�)��nh�
&O���"4CX�Nԟn�����}��C��CdhÏ��?�j���j���}u)ޟw���s�Yu��o��n$�;������%����jaun��v���D�e7P���0h_*����Ύ�Z�^;�ҹ�ƜP�ݥ�����w��־�z��W��g\�u�ޮغ�Ȫw�|]�[��4��q{3�$᳐��۝�q����]�X����;2�N�s��%*�	�L��y.
)�s%�t�s_�s\���5��7��Ӽ��8tw.!�h{��'�� �E1#��&'߇0\�w�Ƶ�����#T>�hw��>�����|Dg�x���4:�"���"5�Y���X�GѐIs"�A¬x$�R�yNs�����P�6�@y֏���h��>GY�:ր��ر�c���F���v�2H�W:Vƻ/��������Q���hv�|{�	w�xC��yĐ!�8���2T���ph.VF�;��	ܩ�5QQ�lbH,�:��,>���Ab�iE������3vP�*����B���Ǆ �,>x4"4e�@D��1�T�n��p��:��7�𸤩�A�tōs��� ��;�D���=n���VPD�pX�������%I��)��+���p��T}�Q$T�ƙL���o'}P����#y����>�uu:����W�MN���_�ȡh��|s�3��_z^�Q�X�{�O��ʑ�v��(D99�J"ˊ]Ϲ.�{�w�}{�罀тF	a����Է��D4��Mg.��I���=|w������qq*��u�� �&�i��W.�n����O�I�Las��r��z�>dCV�g^��Q�u	W�V�U7�km�<��T���Ώ��#�;�K���<��E����}P�]�Xs��:}ǘ�e:��T��Gb^�#ĩ������)A�P��ˍ<B,9�I�s؞�M�;.O���f���Ic<�����ύ�߻�	�Lģ��O�c����,����d�狀^q=�*�][���˻:�9����M��g���"e�o:s�b�7�u��9D]8��o�MN?���SN��o�d��'Y��_=�'8Nw`o�8u��D����<��)����"W7��2�8S��Sq;������R\�^��D��Q�̉�����Ϥ���0Hɋ����bK���s�����1�ӉB���i��w(ʆB��S�g�Bn�1cS~�W�����X�C�"#���o��F�>�&n2 ��w��@i��d(�����(D08���Uq�|�<�vh��"Ky���keg5�ߚ�'}�t���ξ#xkB�9V��r]��y������	^-GI���'�۽��8���w}���ݯ��q1J���
dX�!��2\�t4��E���jE�5��	BP�fw�t]�~�ޥ5�Ϸ��pN�8T<��_:���U�w�k������c_5��/3�
�޿�;�h��Ƽ�������S��w�q�Q1����>{�D�1bI>_�.K�r\��Î-K��;r�ߛ�����vw�&��Nk��<��(,�R	���cs���x�v�F�(�H}�����ß[�n�����	���ÁC"��ER��йr��~�	��7sg{�Y�cLc��T�}�2�$���w�WW�o���}�����9u+���y��������v=�{|���S��B�K��;p�qČ{c�"y����=ϔ���b�I�_w<MZ1!q��A}�m�q�∗���蹕����B��E�~�¦:�]VaP0C@1��"9]W4��B2''����������]Ɵ��e�6�Ǌ#�J�",���W�dR<u�ƺ��؊�ۮ��=��c���mj���7a���:N��ݧmg"W*JN�U�����FC����n`9�;oF���Ɖ]��^�wc%�k�v�W�~{����?s�>��ɷJ�I?�$�$�$�I3�@�  k �m#l �`�6Ͱ (0 -���]6   l��  �@   [A�	     l*  ��K�����4+����;;e��
�Uu@:#�щ���!&�g���
�v�m�[\�h�r� qT���\U]T��{qg�@@k=��a�٩V�U��0�O:��ae[r[f�[�Gg�+/fb�ˢieZ�H�
��6��Y��r�z�8a��۶6��b�݀���f� �h�W5�G�ב����H�q"�m��3�ƥyM�Q�Av�m��#y�e5�U��<�m!ɤ|˓&�]�@S4죗kq���j@���v�V�s���6N��=�5��i�rB�Y���鐘5�\ܔ�P<>֊I���3�ƐX*�R����h�'m�ݕ�GL8��M+����ē5;�G\q��S���l`�����>�8�ۀ��d�ٕ9�msT�Rv��L(�#b��鲎�īҽ*���vFs��jzn�gl�說9pv� 4��SE$rBY)�b]vƵ�Q�݁z����)Nf�^R@��umw[��[p� A�-�&��̃�Ζtj��t�e8��`�ַE	T�sM� �T�$�԰'g`�m=UU@z^�(!��K�b� 嵸�F���9��ޝ��F���9��SJ\�n�A�b��0^���烀*�i8��T�ʪ�.�8{U���ʜq���A�23;O2�JͥZڠP��=(�J�]T��/�P�⪩qg�i%���n��,��6�_5R�mU+�l�<;-Uj����]���΢�S�Q�V��	a:xkp6�ѐ�PV�QR���D9TUݹlһuok�� �qy�Qv׉Pa�\��En���V1j1�`)Nu�*1�ڤ	]c���9B���v}Rtر���ʆǾY��I���i�t��f��i�i�\#�.s��'L���G��K��,�v�#���8�4��6q���DSeW�^W���3��r��0i	���j�[����U�lup�mq q�I�X�-����Fy� 96��vېm�kM��pK(kmCۨ����v�p,'��lp2��WϪ�V�yh8�LG��Ug*��X�� �u���eYU�@PR�8 �ݶ�&��:idn��������ݻR@5�Dsh��};�	����n����݀$'����ɛ�����Qm�;r�PGUUd��
Q����E��]HB;?x_>,��odwk�n��s�������\fAS���럁��e��k7j�mbTr�t�;��
���w%n[u��\�e�m>�~(/�����d�;u����˦��҄�=��d)�`�ۮ�l��T��6��#nE�M��z�� �S�&d�T���4�!#3K4�r[%"ZHGYΐ�n���MWm�'�E{X���G��ڔWf��W;;R2Ikeʎ����Ԏ�ѫE����s��R���>��#/�RW�,ge�ٱD1F��#樇��lGI��ڀ2�k/';N�UzX�P�-�UP)-*�J ㍺lۮ���]��7��UT��n{�2�e_e$�j����U�7j����j�Ļ1t�&�0� �m�Y�c�F�s�i��3J���� [%�����fq��i0v�;`��}���\^A�m5�d2���`^2)V�n�����Kʚh��H;Zvݓj�6Y+Z��mi�]KiV^^�[���l;I�*�)m�n�6�Q���h�R��E�:wYpR��nZ�h{Lj���#UpluPغL�l�K��2��U���ώ'mFm(N�9�u�ݍ���a5�ˢU��;h669wVx�ra�g4���Ѽ�D���u�zz�<�܅��vy6ݖٮ�F�oH�1���8�=n�����:Ӱ�tƝ ɛ����]vڽ,s��9�g�������f��G(]��½]c�ch%�n��ڭ=��ݮ�6�Ŕ����"mIq5Р���g46zx\�F/ŷ���6��=�`��[a��*�^k8�i�klS�ק���xל���Uf����a�F�W/k��Ǎ�m�M=lo5W��X"^)ʔ��,MKˍ��sh�<][�/c�ʪ�Ռ�6W���`;F��G�]U!OmR�vl�ٕ�yj���*nQ��݆���̐��9�����ٕ�0 [Ww��	��4PP=%�V��S�]�l���{(媨��௫�u�\��*�QF��/(� 8�v�Kf nsj!�9mm�ԫַK]M������I���m���p�N���ۖ�8�I�n���g$��M
V��b|϶��r�[�N�u�����MR��p��S`⪪�7v@���nX����m�`���d9&�^Ѻ��5�Rܭ�����Wj�ݶ�+ u�]�����^Cg	���@��Wf�.�I�o[�H�l����կ\F�v뮭�a���kc���8�s�CnUm��'��t���e;s��ܫ�
(����� ��NZ�R�*�nܫm�t�CmRݳBL:ٳ�VԮ͵]@Zup!D���d��ҍ�K:��ij�j8(
�x�G@��X�V�9D�'eT�f�h��ȃsn���*h	V�� �e�W���Z�^�7f�����Z�q(�k���N�J/U���mm�M&��8 �]!�j�J6��Y�C�	�u�#��I��;[RP��c�4�-H61��:��F�1��UU�VQ�;S�[�h`+�ٓr����ȃ ��J�ڧhࠪE�i�{;�8Źo���o�۩�P�{����+l��i*/&�ٹ���$sr6�@)��=�Fe���y�j��S÷c3��[�r�.�J���8N�kU�.���{IV��u�p[B۪��6,xީ�j�"ƥvz	�͋�A���d�m��j�b�(���[G6m�H�T�L3��Ȑ$-i4�6Zl8��T��M�a�^PZyZ��稝�Ӻ�p�/N�l�Umc(�{`�vR���,���Ƕj@H8l��]m6ut������ڪUٌu�U��riq�C`�!f���^Z��Y��Y����E�[tͳͳUm���OUʪ��.�[�U�VYnI�f�Hmy�:z.��e��Z�l� ��R�xn����S��y�������ۂuU*�EZ����'E\�=Tg1V��n�5�:�y�@[M�~~>���a��m��˥j��v��3��4�UUTgPX�]c������<��I��,��*��]c禚����C���������"�lYv�q��t��m�$r�n��\	z��<񅝖�Mt;;t�hhH�f��a�v�.x���ڀ���7�+��`6�� 9'WJK5 ��d�j�ceT�l��6 ]&��	;vͱ#Z�n�[Pp]Kp[�T��m&��eU�Z�����햮U�Z
�kB�n��v�H5���L�5T�Q���m�յ��WR��$ �1e�1n�"H��܆��ܕF.^��m6��z��Z��(c#m�ݷt��UUm�S���e%���sC�#���V�9���d ���#�	  �mm�^�f۲p�:QF��iYZڪV���[���$ ׯ^x8Sb�[�6�����K�«�d��k���{�~v6���J�V0�]�mYIAv��g��㮺5:�N��j�*�	�A-,��l5u���p��f�`��cs�p�l��;q#�1%��	��P�K�[!�YG�n�8%�˱U�er�Cq�v���k��.��;��C$bK ��RP*�&��\ҩ�{vh�  �%��*�"%YZ�A����%�����A�9N����+��E�CXc&��`znp5Uv�u	湼�4�ln;#�NlIoM��Om�;j��2G	��'BR%6��8�ؙ{��S�rEZs㭸9��a6@�ڋv��lln	��]T��'4���(���mSUj�2YV�m�ݦ��� Gm,��k�	@���gퟷ�6{*��tn���S�v�Yڞ�omAI$��]�[��vS�՛��3�5;/���|U�]��<OncE�=v���NZ�3N�]UP�������%�"We�3�rAW�[+v1�E�_f7[���-��.0 շ'd-;��Ė�jͱ�V��]��[�T��jUs��ԫV�ͥ8 ��򪭻n��j^W(�h�*�0��5��l ��C�Iv���d9Kan��m&	C��l �ݻm�vZ۶I�ȡ[�W:�yh
�6⌛/I6����m���E �m���6��t��tĊP �a�n�926�b3����I����ֳi6	����$�=��
�#&��P@U�#d���LHLV���n�ZI-[[0*	��R�l������6԰6vP	�o.�ڞ����v;WW��0��.a4+�N��T�Ԫ�UIe��V����[j	:M�v�Y�V�ٚ��P�+�+<�6ݥn͋9�{N��7]���ek��s��!ԭ�˶J����J���lJ�hs�MJ���n��Q��n�Ip2�+� �*�6��^�$��[y���D��knٵ6�P��$����Ԝ�n}%Y�kX(
+j�j�8�k4�U�J\�ʻUʄ3��v�]5U*�l�U@U[�Ŷ@ $�GW;-����^8���J�����%he�Xw5=�L�CXEi�rΠA�p�����0�[#�j���T�� F�m�l �i���N;J�}��(	��UuT�ͪ����`,�v2��8ƻ�}!l԰FC.i8�m�vx��*ԃjR2�KK�+�|0�33����U�����PO��A� �����(��(��(��(��(��(������J�(����������_���J�1� ~ST� T�0@d#�CDPL-)A1�m�۽�^=��~߯��q�\aWU�q�\aWU�q�\aWU�q�\aWU�q�\aWU�q�\aWU�q�\aWp�Ç;�`aÎ��p�1�\aWU�q����/��wW�����D�O���d�Z��ڠ`~�# =�lH�#B�_":�|4 �$ǳ�
�� ]���@|S\O�����~t�z|T�P~H t�h��O���t�:Sh&!�"�9��� <BP��H нm]�:A�(�*�����"q�H�� P���BA�P�G��SH���1>=��||U����	��hC��=_d��;:z@�&�к{U���;U~{�� �m=d>)�� �U_{D�"	����J�$z��������Ѓ��>����)�T0P��G�PU���͢���H#�(h؝�����Lä�t#��T�:(ǽ
�� (�
����t�:(�E~�`	�@�=W�� �@HC�W�∿�B=�2���	��"'����"AJ,	��#��(t �稊x��h�!
&�"�d�bZj�
P
U��(&�R�`$$H�"R%)��bPh����)V"
eү`��!;~"�� |>(���|@���F �B���(�)�PR*�$
�� �dQ�<6�>D��1�JP�l�@�ôj'�|�D C�pz�J��"�B���c��4B�(��!��@� C��IDU�Kx��@��i:US�  �@�;1N�w�M�BA������_�����:�������G��=����	$�I$�I#�����u uA�0�,���CA!&�0�G15.�Wzv.a�Ib��)!D61-�H� �a`��k+��M��TB$ę�q1<Tu�^cLhB�P`���}��{��b�ݨe�*��6-�s�O7kt���hk\h��rf�*�|u��E��ځ��v���xڻ<�������O׎#a�wT��'R�)��l��`�I�=�O#r�c���`�;OJx1��،��u��A����ݺ��Bkpk���d۶��:�N� e�5Phʬ��LR���jLX67'c��Y�ܝ�� �/C�(��:v]���ٷ@Fs�i9�M���8l؍-����sm�l�ؓ��X6�s���#۳���ۋG1�+�<݃=b�I���*[��A�,M�P6¼��L��riK��� �eS��`M�v�gE,�3m�1M;U���k��]ʹ!���C�j�۵fz����7c��ƍ�VWc��N��D7ub�mk��Z!��6vG������b$��s�%'NNwNq��]��6m�D�8�r�=k��
Gv�{\���u� �l�I���a�P��S�l��ֹ㆛X����<�;Z�\�[��ss�9���=�цdy���f��[u�<cRt�V^c�s@����Dm�\c�O(\�/C���ۃ�ޱ�+'m����[��@���v�&�>���=�n�٠qt�D.jcu�{.�9n��su�=#�f{;�����u=��8�C����'�L�ʽ,1p�-��9�&�����nDÎ�c<�FuZ	�9���`��̓Hӳm9pgfȌ&ݎ�nw[:F�U�Nɵ��M:D��t ���!N��!���i�n\�gŔ�)ڬmǇ�P=kfMɶ�Nܹ�-�;���mی�V�Zy�y�������b�ر1sjcc��A"q��7@��8���G�[��^6��������3�L�ۛS�6{u�^��1̡���d���Ç����(z��M�vR��l�n;i�@�jwd�^pF��r�ӛA�Y�b�by�n;J����f���P��s7k׎��Y�Cf��\=�j��v�ڶ�¬��<d�\�Ʃ��m��[6x��S�����>���N�U�@�N��!�&�OE$}>�j� ��N�t�[ߣ���� S/I�&�ا�q�I��f��r�3���-�f��C��^���\�p�/=���뭫v%�v��nٶw��؎��`�Ͷ���ɟ��q���U�6C8��zMm��p�N�t*�k�۳�ػn�Iv�a���`�0nR���n���7𣖎^ʢX8:�9��9���Ǔ��ٓ�� \�ͦ���]ruSF�GIl�������i�;�iȱ��A��Q�$��ƈ$L�I��ܞ9�g����g�eq9
�q��w�p�}u����sf���o\M�(�RA�V�̖{캰;�0�9ט�c��#Q}IQ�/=컫�B̘+Aμ�V��K�+����T�HS�U��Ʌ�μ�`�d�;�eՁ���ıJB��j'�y��=��~H��]����T�^2&۟"/�T�՜�g�4����<�����7gs��;;.�T�n��5"�{2X����d���^b�9�S)'���J�rX�{��߂G��C"˝03�~���R]��V�fB���ڠt̤�$m������~�`�d�9�eՀ{+���28P���s�1^�Ԑfn��ͺ���I�ޖf��Dc��S�	8��̖;캰3�0�9��V�_V��IW(�q9�l������g�[/A�XV�c<�r�9��Aƭ4�]�N�t9G>r�@���;�۫���~�`�d�8��K�R1�B� �J�>Jрoݴ`z���VF8�r&G)�H�(�����d��=��dx��b2+�,�,�*�,�#KC�|�~�uW�}߷@w�<�q5%H�i� ��%�;�]��]s�x}~
Ř&�r2R������9�����ޡϾ�����D�x������F��[\4�<K�䆴;�9�O�gC���� �IRV�q[$�KC�}�i��<��}�i�������FIr����U��9Ȃ>I�������R�K�5B��.Z)\�[C�}��]�z�� ]��~Ӻ�Wם(�d�(JJ�˯w�%W=�{Nu��^�a�#�����g�����l�Umß}�i�?��}�i�~�uw�T$J�*6�Q��G �Z�!H�iٷ���nN��I;[���i����g�y�����]���ʐ��;��G\�:V'#I�>ｏ.��x}��e�{�"��f"�#r2R����q��=�����ǧ��ݺ��&�7�M2F�RB��G�o#�N�>�%��*GR
*jiTK\Bq[�{��s���Nw��>�����<|ğ�-n�Wh�\��On�]YX"5�:d��l/@���zO����ѭ\��E�:2����D��㰜�k�z�py�{4�j�g�66��L\b��;���U����u.����H�qٯm��m�$�G:�7/C��v�ە�Z�����Z��=]r��ݧ��Nm��'%��#8}=`�C�a�x�W��{��=Q�1���Ku��3�L*~/{������Q˜;<��rOI��/�w~5����=��-�7<[�r�,&+[�iU����;���f]w������XJr!�����.��u�ꢞw7y\���{�uδ�?��(�T��>��;�z�}��ӽ����4��g�IX)Un]?f`�yGZO#~T�wRY����j����nj��w�,��JË�,�������G;�����FZA��:A�Ԛ�U���÷U[݂��ח]�[I빧��I�g�\�:�U�w��$.��7�H|�#�CM�"sM�	�#hmI��̽�τ�����LȂ�&4d*�AQs�&f`r��>���u���j���4޶�Ϝh���^��>��e�{���̺�r�OB���pQƫkﾣ}��Y�����ˮ�Ǩo�B��JҲZ�w���w�����ޡ�=�i��S�2H�TLu5vk]�n�P� v�펛vWq�Uy����dy�׷nԐ�%*�c-E����i��<��{�ӝǅC;�����#�H��^�<>�fe�;����u�E/<m�qQ6���K#~T��DTA�F�u+YuR9��*ϔi�$%(��\�<>�{2����w3.�3Ɍ�8��SJH}��ˮ�����i��yg�w�!�p�I�9&<�,Yf���3D�<�N�y,���Kz8uԝN�Yoi;ba��E$��W�2���w���=����ܠM��8J�Dԋ��f^�=����ۯ{�"ҹ�����L�$p�]x�u�ԖG�*GRY�LOj�I˨�VY�����淪?}�{�3�ǅ>30�`���/w�7[~J��B�]�t��Or8Ӗ�>�<�RY);2��yS~M��'N;c���݁����Ꚉ�Z����	j�;ml��W�>������/�ٙuޯb��Խ��$p��nK�uf/��f]w�ؾ�s2�11���J�����.���_{=�uά�A�z���(�B�h���]��/�=�uά��g�39Gr�#*&���p�3ٗ\��_fg�4��z�O�{�g�7j���J��7��s6G	C=d�+[KT&n%�m c��絠�
4e���sb^$�Va�/[=�Mu���j-kō��f:�q�{l�Ӽ��u��mڹ��ln	�]c�r�}o�w��|�ҽAضD��/T�Ľ�s����2\�ٲɑKɖ(^_Q�0wOn_'�-n��N�3�^�z݄��q����:��D�m۫�5�aN���a���V�����J����]���>��L�n�gN�����Ůc��-bJ��J�$�I�����33.���_ffe�z��y��D|�#�ٙ�u�����f]s�1}��H^��TC����|��=��^�g�2�1���!9Lq6��{3.�՘��fe�{��+�y
$NI!R����Q���fe�{�*�ٙp�?�۶����4l�e��[��<�{b�'8-�X�1K3�kљ;b����rZ�r��%U��%Ց��\B�%{��9͏�2�s{��O��[Vֆ�w��9á��5 �&�� ��As�ۮ�f{2�;�)# ��D�p�]K#�uW�Y�R9���Q5d���#r�sٙ�u�����̺�RJ�y��O��I��ff]w���33.�w1����O�J ���ek���H;��MΞcv��ڷk[t�q�'a�vg{Y��Ckn�:r����eVff]]�ffe�<�K�P"r��nO�f<�߾���������w���慠�ג1���9!*	˯�g��}��������o�I$�I#m�{��O�$S�>GM����Q��l��;O�!�8���a��;������.�|��>��������1	DI)0yP�H1"�&.�L�����bdYfo=χH>GZ��%�"X �$!:�l� �0'���0I3��p�� lR��	zѲ7yS3^(p>k�=�1��,�N��t���C�O}�sk�HP؅(��jX!{�0B<���̫�Np�]`i��Ç<��Icp�<x�9��84��(��>[���:P��B)���A	S�BJOe�$�	�&P׮!�$��ji( �'V�ڻ�@L��;���"qkC��Z�fN^a�6AiLI�C�X���s���܁�`DGO����ӱQS�����ߨ��"b*=��T��J衙�)���'l ��x��C�;U�?@-�Hm�%9��)JY�Ϝ��C�R��s�j���7�Z7�������(y��Cܧ��39�k�)JNy�s:�(?A �湜����3�~�$2O宕GlF�n��ܥ)�=�5Ҕ�'<�9�'r�����JR�<��s��R���s��>�`�pn۷]X���S��\7l�=�Dv{=��֭mrk��=��-^�Q��{��~[�I�o��{��<�}�S��(y�y�t�F�)J{�y�])JRy�"ßk[��ś��Z���)O3�y���(y�y·�J�{�k�)JNs�s��R���Q�5�:-�k[��5�t�)C�s��{��>g��R�)9�s�r�����M�����6��gꄫ��^�����J>g��R����:�)O3�y���$? ��	��1�n�U��$J�B�'^���!ǳ�C���]�=�R���?.kY��of�o[ѽ��)I�s��{��$>�)�9�`�~����^��ݨ��z[ayn61�Q��p�nw�ι�sq�����U�<�-�5�v�q��.��5b�緙��?a�L��=���JR��=�:�)O��t�)I�{�t=�R�˜�Q��VG!Y����3��~��q`��yκR��'9�s��R��=��`%�$g}��NOֺU��&���)J|�9�JR����C܀����JR�<��Cܥ)�8f�u��{-���[��R�M�'9�9��)C�|׾�])JP��r�������D��缄��7*��u��j�8�)�{�5Ҕ�I~�8}�����<���])JRs��r���=>���c0F0�F��liXӭ�$�9#,r�r�D�E�s�8bWM)�h{8`��>�����tH�n��֒�b
�ώs�^u�AH�۵�S;���=e�!�k�c���f�k��r�'tN�t��͝M��J1��-f�C��:ۓ�ko`��5�WKn����A���\���E�^^�����Ԗ�pZ�ͬ����n�;&�L����ҬZu���+�ԅVR��330�0��v	c�2R$��X��D�LCE�A��v����r&�1�e�D�$I�d��c$)c�}�%�$g����η'r���k�Δ�i9��s��R��}�R���=̳�0��y���}k�ﮇ�O��g9�]JRs��:�)Os�y���) �9�t=�ҟ=e%�`�	%!ƣ��U���G�P}_���r��3������d2����Cܥ)�>��Ҕ�'>Uy��nսlգvk}p7���׼�JR�<���Cܥ)��o�JP4����Cܥ)|��kM8�U����Y��Y�F~��~�8�
訩>s�_n��)>���އ�J��{�5Ҕ�'/���&e�h�3��]�7ZN�*��Q��N묎�N:���a�8�YLVjM�=���,fɻ�g`�a��o�JR����Cܥ)�s��A���J��߽r��߿~�4fu��{3f������)JNy�s��?P>���!��ꈮv�Jfo��t�)C��>��{��=�7˥?%)��A'	'�E"n]}��>��~����)C�}�:�;W%=�s��JR��9�t=�R������En��f��o])@�<��s��R��=�5Ҕ�'<�9��)C�<�9�t�)I�~mz�J�څ�fۺg`������Ҕ�9�9��)Jy����JR����{��>��s�DY���̳{=��k�����9L��9��mk\����yc�<�����W7 q�⿾����������JR�s^�:R����:C�JS���r���{������.j�*,����)��s�tJP��s\�{��=�9�t�)I��s�p��s�k5Y�oY�oZ7��7��R����{��=�9�t�?�u�J��̤��e0���&���p&XC0,q�F�p,)]!�~#I������)J}����Ҕ��=�fj�7m�ް�Z�]k��R���s��JR����{��>y�s:R�(y�9·�JS�������RGjVٹ�Y�X~��ߴ{���s|�R��^{�9��)Jy�{�t�)I���Q繙�p�>�U��wd(Gg�s�h�f趮;] �Ή����'l�د�[��U��vʤ�gV`�'����:R����r���k�gH%)I�9�t=�{����Xg9�
�a�٭[޺R����:�꒫����}Δ�)>��߽Ϙ�)�k�Ε@K0K��k�o�U����wL��)O<׼ֺR����:�V���s�t�)I�y���)O3�3��zޫZ�Zޭ�z�J)9�9·�JS���JR�����!�R��}�zLJ)��R�X� ����� >�]w���)>�W�����oZ�Z5f���)Jy�{��JR�{�o��)J{����JR����{��?_��}5�u���Zњ�-��z-v���l��k��]t��Zt��5gn�����ǽ�ݹڤiͩ�m+*N׹�Fu`�������)O=�9�)JRs�s�"�K0���繂Y�Fw�~q9�V�	ck}ur����΅ZR����{��<���JR����=)�{g��#rR2Z���`�`�����3�JS�k�Δ��J�I��~��=�W�V���_�P}����F=I�B�R-h�Cܥ
y�{��<�%)9�s|��JS�5�gJP�H$�Ͽ~�=�R����Ͽwa[�5�[ַ�)JRs�s|��K��P����t�)I��~��{��<��t�)I�ӤT������sfg��n����ۄ���^����l=�YWt�p%����vɺ��v���m�`�i���u�m[!� Ӷ�`�{[{<ni�5���v8�;q���ᇛ.�U���;vn�$�ëd?����b�l�T���7<uw+�8��='�^�x��2��u@�� e��ȇ��t���c�v�]�׵�l�T�v#�{as���ζi�ʈ��<`C%||v-����8���w��^�Z{an.�<��u��8.m�Z�Q�W�͕��{UYk����u�)����Δ�)9�9ˡ�R����Ҵ�'=��=�R��Y�o[ս�z�7�f��)JRs�s�r4��=��R�����r���}�.�)J����Q$� 鉒��}A��w3��JR�y�9�C܁J|��t])������Cܥ){s�Z5��Z�����y���)@��>������JS�s�GJR�����Cܥ�Is�s��R��󜾖�Z��f�޷�35����JS��)JN{�s��R��{�7Ҕ�'=�7�{��<�9�Q��n֥]�z�-�}�r�u��<u7l��90�np���rItI�R�[�{�5�%��~�s��R�$�=���JR������D��ߴ��,�,9�!{����v�Z���)K��}���O�(i��C�N�r�!mւ�
(DG%)>��{��)O3߼�Ҕ�'<�9��J|�Ea���9����[��Ҕ�'=���=�R�=��)H�s�s�r����y������iz�H�T�Uv��ga��5�::R����:�)K��JP����o��)J{��g��oV�[�7�ݭ�)JRs�s�r����y���,���|��'P��~�:R�����ZHUH�t�$�P#(7ݔ�ls�՘�۶�9Yڎ�h��^���t�K{K�5f���)B~6y�}�J]b�'�}����)Jy�{��JR����{��*�����I��EQ$俾����svl=�R�=�9�)JRs�s�r�����w0K0H�{��r~�ܲV��݇�JS��0�JR����{����?aQ�*��$$�� �0��>�Ͼy���+���d�W�>���wca��5����'Cܙ RsÜ��R����o�)JN{�o��)BnO��Δ�)>{���+K+r؜�g`�`���]�)J��|��w&J{��t�)I�y�:�)O�k���Sj��{�af��ٳ�=�^�ۖC�g1��l�<;���v..P�=���D��c�V�e��%�%�~���!�R���s�Ҕ�'<�9Чr���=��R����g�a�q�5�޳{�]Cܥ)��3�?!rR������R���ϻ�JR��{���SR=QA���W��}A�o�v�ߘ�){�u����)
d�}�����JS���ܺS%);�\�\�o7�淬-��o��R�o9�7Ҕ���{���)O�k�Δ�? ��H �. Bħ���(&����'���sL����_��iG����J�ە�R����|��J�!���:R����>��{��/9�7Ҕ�'į�����'Pq��M&�
�[r0��;w��%��y���k�W[8�������;���ַ�fog]Cܥ)��JR����s��R��s�o�������=�%�~��W	�E&X��Ii��Y�Xs��p ���=��R������=�R���tt*�)I��r��z����Vk}r�;�<��JR��|�^��iO|�::R����s�r��S��Xg8۳y[�������/�aG$������)Js߻�t�)Iߜ�:~b�U�s�~����)>�Ɨ�6
�d��f�qaŘ%�{����)J>��}��z�����}�J%�%������,�,�������d�I>��m��d��i�~���4F$B� �:�l��*`�� ��I�j,ndacz��(�z��"�T J��-D�[;:�L��,)��F��:L* �O��H��6Q]|�����/����h���֠���:�n�f��؆����|l0��oAC)`�v.8�TM��=�;>g����N�W�Ԧ�c@l�V���,V8`g9cx�M�i�:��,������5.kIN�$��ލ*Zn�#z;�2s�sn����z����������h��&��&�+������Q�����L7�7A,À�ӊ���4P#��o�"�2���2�X:���ɔ�8X�'�D�v���.(P:�&����[��[T�v!ڀ�I�U��-�H8_]]5%�ʜi[$;$I5�F\�<C�ŷ4�bS)����l��:���':�n��s�!A�4:K�+����!��� ӊ�vvT60�+�q٭H����z���ՉwS�7e�Ò�2�����
"8��97nb��=��ϵ�c����Ɣi!����us��8#r�wٲ5��\��g�� ���ˮ�n������v�mAT��M�N�V����ˉ;s3�n��&�/-�n_!muy�I�c��#l��Qq��T��v{u������j�������ɇ{���*�m�"n������q�1Ŷ�Y-�l����험�!&�;;p]�'"�i�`�v5л-�۲#���ܻvf���ۆn�S��ڕjf���(��9������]�R�hA׆��m���vd��z�'�n���ѭ.v�=�Zi{kB�յz�)�;l坡��r����ڭrK���M�����X^�zJ�ZZfv!`�(�-��!�X�8�z{7;b��2�a��I�����S`���d0�e�3}]����\˝c�6�\tM�Iܓ��#m�vɺ;F���&m؇@�;�¹�8:��(�/nԳw+�`�-���p�i��a���얟#��tP��8$��e�˰8bG\�Ձ8�̵�ն囎�W���%�l-����`wA�k\f�^�C����&��Q��ݱ�S.ܺ�)W,]���G` ��n������ne��ɍ�gjǭu���.��L��l��ơq�]��2��4�W�����V`�÷��8�q���z&H15k�Z$.4�t��ڜ*h�k�lϞby�Q�;��O/:��㳭����m�]�7f �����˵&��u'QS4�3�u���ײ�RN]��u�bcu�{�f�OY�6�Ë���A�h����m����9���*��.�V�M�[bvV�<�t��ݣ4��ff�n��������_���TOC�>(�G�����}�DOD1AT@~ ��= �`�ȯ�WIerJܤhP��NF݅�zɒy6ܖÍ��M���<l�'J���buP��7��l�F�*��j�XE��5�[�q��`]U��;v��gj���,6������\���`-��#�ڭs�Bs�ݔ�a�i!�s\�V��φ\]��j���&!9e|1�g5�2e����lU�)z�Z�Og=Qv�m���Мj�+ѹ��?�@� f�$�|��ǃ����R�6�s/�5и�ٳ�U��;�44��\�܏}�_="ڪjZڒI*��,�,?��翺gr���׼Δ�)<��{�C�JS�l�����>�tk�QG����)O9�y���d�����;����۠9���@m�1k	��§��R�s�.�s8{�������z�� 33]l�T�G���]�k�}�{��jm��I��i΀�����Ҙ�c��`s7w����5X̙��g�iv���ʭ$QH�	��W�Ѯ�ۃ=m�4�2<�;��1�������HFD�i�� {�5X��� �<����Fć����:�"b}����������Us�s�]��xGX�)2 ��HD�4B��QC��];�y�=�>t���p�'#�	�E��܍I9g �{�X�ݮsWԏ7���L,y�^f8��"Cm�EaP4��:�9�>Jс�B�8���%�H����ך�ﻘ��;�%8I�6C�< �����L�v즫�ewld�n�����zZ
ݶ�앣��m�K��STQ�Z���+���޾Z�ߩ)��\����r �r#���p��E'M�EO���K� ��u_�UU��� :�9�>J�����J �Y7%2T��$�+wۼ��y�����9�ڈt�	��{��\�^s:��|����[����Z�}��*����wϹ�	�fߩ)���9��&���&�JR�"�8����UUUw��, ]M��I��H��vr��&h���;u��&{lۢݮ����UT�j+$�E$V!V�p����[`�����Àg��56�@��9�qL�B�H�;�$�қ�����V���}���ٓ�~�u����34$�N0t���:Np�V�9�p;�mM�� ^�Z��Gn7����ovu_R%7l�U� �m��D~DDlr��
~	
8���W�	����:��翎�lt��O�i\8{&����_Us�~���;�~��Z0�,�T�\�X�l�q�wkC��^�8�!��J����y,-��j�d�0�q�u[�����I~��߸�!�� ���r9� w��0]_�,I��%�]�D�7���0k���0�l�<�{�r#��A�" �)#���d���}0��������
��V�����}J)�p�"U� i��vg���DAԭ��/6��F�p���`nf�8��Ds����:ݳ �ݴ`��T!��'���̂���{������c1~���:h9�������u����0Fc�F:�9H�ͭ#�ܺ�X�S�P6Ɗj�,[t$Jn�`�@n�<)�:�l��cF����I�h�3�\(�)���ا���t�]g];�p'Nz��a�s�ֻ(�'Z+Ӑ��ɺ��c�[����.�=v;OO.ƌg���8���Z�k���E��v��X{3.n'����'��w �À�M�(څ"IT�I�[��ձ��2�:�@z���km*HQT%��E��1�*$��r��0T����6�;�X����D ���t�6QS.����T���U� ��Y�ot�&��=����7�PQ�ˇ ��m� ���9���s�}�hó*�L,���
r6����o�w���5^$}^�O
�+�w���(�)}(�܉��:Np����t��Ռ�?f��wM�[��%$4�����s-���h2v�ȝ��2�\���܋r�۾�������hDqH�V}�2+�y����Up�Y��%����|Jq�!ʾy�\�� ��W�؝W�u���u|��z���_-��f����DӲ~��;e�75s�y{�������;�h�7�1X��m����`���p
��}):�;�h�7��8��[{�@f�mH�Ӧێ���a`s�ج��ۻ�廮���ǻ
��d�U�0��u���sp��v��y��I�8]���/BN�����16�_�|�C��y���6�@�Ru��9�;�h�3䠐U�]�B�����7=��_U|Y���&<������9�(X""�I{ﺾg��]U���]g�@zP! �U�=���9��^��.��hT�\���L��9�G9R�`�����`a�_��jK��o�	����,q�S@�Rs���m���� IZ0��}Z�h�P�\�"�Jr�D�,l�p)W\�wI]ͱu��ԓ�6y5�aY�	���.���=�{۠}):���Y��_W�=酖�{�V����8�S��;)���" �T�~���[w��K諭A�?/Ʌ~��'�ӒX��}�Jt"9y4�H�'X ����2|F�.�﫸�U����}��=��� �QS�t*z��!�{8X�B"�Q2�*HȜV~�k���u�o�Yo��8�"#��fn������NS�sMm��Y�V6��{��q�G�vY������V����2h�dπ���7�0���9�����BBͨ*	Dq5v3�ue}���WT�u=�>��Y�r �G$<�̺�OYu2M�ƞ�N���5�Ot�����v7v�����d��rQw75s�����0OS�WVF�~�`o�Q�=�}�H�Pns�u{`9���q�o��8]OtȈ����b!�{s�f�-�[�f��b�֑�D��ӗ�ζz��m�t/��,�]\�S�9	3½[�Cŧ����܁G���R�q�獦����Xm�>t�m��7�;��t��jYֻ]b�eӓnSN�]H]�-�k�^��cZ�s�U������7'p�����7;l�%n�B4b�6�͋��#�ػ*�XSb*z�x\�95I&�o$�K�m�#Xp����S_-@ݑ�Q�R�u��k\�������۞m.�+�CY�;�����k��j��L�GM7�5�.�y������W��+�ٮ�3٬hz%Ly��fG#�>�=�r9�e?V�٥�URG�UD�R�mJ	27�<���ғ�r8}�h�;�m���"""�I�p
�����,�-~�܎AȈ���{tꉙ�~�*	Dq���>�������L,�n���K�_}���S����F�ݭ�n��a��9��\�u��=<�m�\�!4 ���S�H���V�ot�y�G ��р.�2Lv�R���Gez����~�?��0�y�7��I��zS�	�L5ã����
b�1޴/ɑX;<` �?�ﮤ�߯�jK��y�f`K��T#t��RHЩ��p�ݖ}�۫� ��g�׼Ϊ��Ͽ{�������Y,v
9n�a��z�jK����������9�u;��:
���]�RU�ݤ� "9�s�i7��f�
;�1X���E[t�(����v���G�W��5V��}=�F�=�-�'Z1ٮUW�}�QF踚a>L��`~�����S��UZ�DDG0����P�S��DJG��
,�vq�+����Sw��ȉ��9'D��0�� ��t�����9��V:�����s��m��l�[m�{�A�X�bH��S�(C}l�'L�Q��Bl��$n0��(p�0�?�*��wu��}�`�&���.�%2	C7�؈$���N�)06F�f�ߕ�oȚ��ϐBP�F�>=���U٘=���d�d�yM`gF'V�
(
���c4���v�;#��g6��3��
h{E�5���R|�:��vK$BBX�,�Jw��3.�4��լ��B�q�"b�;ww&ua�|4j`�pʨ��SW��	,ɜ:�h��؛N�X>�>��O��Iہ��'�=��>��Q�7����VG�\|QګaҠ��o�&ރh`&��D�}�tO�� Q���.I*�E]���΁�Ds�I� ����I��i)�3���)�1�8�7ٻ�_U}���`��VPs�ج�3V�ʫ]r��1q�k��Sm�$���V3�;g�[6���m�%��~=�{������ZU�;��@}���IN ��~��؈�D�����K(��e�2�n8�G$v|�' ]� }M��29�eg9�G |���("5|����M,}��w}AU/��ߺ�=��uWϏ�o�� &���dnU}U�Q�ٻ����Ϊ���� ��	%�R������zX��׃Y�H�Q�I�����s��s��U)���F �O�$��������V�q'�Ғ9WW���s�g)�Jf�g`�1���NԛmB30�56
2�(%G��X͚X�L,�M�G9�4�NphD�#��**�n�l�>jـ>��@]���C�F����;�J��ТQS�����p�Np#��D�`�������' ����p
���<�`{�0�+�酁���p��X��Nȣ�����V�܈��C�{���й��uWO� ���������+-�nh+v�����x�[7B��m�A�c��k]K��ۋ78��E϶��4}*�"Շgl����=�nw��xd�z:�0N֮��}����fywXû�I� �ۄ����{�N]�]��w���cs�c�۞��ƒ���.��|�t�>�3ڦȜq���Bu�!8Sѝ�+��&u[s�1��g�BV�a�jQ�\u(��.a�2�a��p��7A&�����ݏ�u�n���v��W���g=sZ<%rn����e��q�BD��@���d`��@}�� ]V�p�܀�P S���V��p��}M� �x��<����@�sWSwI*�159�3�uX�?�}_UR<���<��n���f	qW�������������:���>�otr!v����mD�1')�!�;��V\�!�7��'8�|�# ]��R�H�9�V�.G�W�ƺ�7����o���*�3..7\ԩ�ҁQ%Qϓ�D�nU��������$�=Ñ�s@}V���z���(�d��I~�����?��0k\dc?��|�
>����ޘ'��2fG
z��DEH(����))'NT��`{vi`g}0�~����"|߽��?N .�A5TU9"�q�K�YO�����Y���f(U溜��vO��S�#p�7����ۙ�>�s�r��# �Dq,~�߮�+�����x
�q��v�9���=�`F'M����G]����:|l�=]y�>�s�u��F�;hȀM�h�%F1�� )���d���z# M7��'9�p]!A.�f$������4�y &��#�">�Gz���dDS�:P��4o�=�M,x����Rt�#I�nU���=�i9�U�0�Dj����FS�����D'9�3�5XW�}֩�/��0�����J^�D��R[��+��]��o4��3��3�}s��qےq{i��t��\jBnG"��ߟ����7�Y[ob9ȍ�I� |ԸI���H�%�;��W��U���{�	:�>�a��z�EEa%\򮨺�����I�s���G>�X���`r��:�����"��pr9�e'X�Z0�VF��DDEw�U��~�/�5��o�� �JB%#�:��0G9������M���� ��{(k�8Rn�O��7B"4rk&k��c�n�;U� ����X��IVC���e�4��J��\��w2i`n�w��3_���76i`eh�U�:#T�jB��{��Drc��䝖�X�a��!
9\��p���ff�f�Z����~��Z0�ٴ`m�� ��_
�%%%T�q�}��7&{酁���DO#���V uz}�U��*n���4������{����:գ��b'nǀ!� IX�1 �<��3?#V����dN�Mv��+N�<���O�z���\�g�K>7e���k
�v���)�8�nyn.^�Ƭ(���\֚q�M�;5�g��y���6۵Nwk)���Bvےӝ�(>��oi4X��������JMq���1gh�ru��uj�;���xv����K2�u�y�G ��.�K�p��.}A�{n��6��V�åe�i#eySqնJ�1��0�� u��hn;aL�I�ooZZ�.�8V6}�������0S-��tq+�d���%:��hC���X���8W�]�ܘX�aZ���7&�F�8���9 u�F�vрu��H�%V6����Ґ�8�5bɅ���a`{w4� ��5��Z郭�Ģ�V٠w�ف[ot���@~�9�s�9K?l���V�%Y�E:#I�!`{�=�;3٦� �V��h�B|#d�۴/�����b����m�\��z�.��w6�bbO�eJ=��7(��R]�K�u��u�F�ݴ{���#d��n�w��p�.l��������:�)��#��"9�"���#�Cy~2 ߼����� ��[I���Q�2]����K1�{��9=��V �M��v���˺���������"��{�h���`u��?|�����Q�g�u��Ԩ��������=���:z�� wͽ��m���?S��ɶ�9��a�5sbeK`6��r�\bG��Q����X;��{=�"�;�O1X��wy�:���f�lm@e%)I9"��d�����O[�%h�8B*fc����B4�q�`n��8Vf�?�T���|W������V�}��������U���
�"I�j����_������;��Y�}�m�ot��y.f��⨓���Ʌ��w��X������`s蝹�כ
����5"�'�SϮ=m�7�/=p�\fx�Ѹ�y�[�0�㟽����.�,��4Ip��M,���
�[�s���6���A�eTUWUsUf��߾�"��IR���v��������_�����Ԥ���9�<����V�9�}�mm��:�$���#J�]�oSY�`��Y�.��i�W9�s���>�Aؓ$��+.*��$���ε�_u�^�=0L)�O8TU��٠.���~G"'��G=�{��|�xJр�"�H&Jv�n$�m�n�׷� ��!��a��y�;jB���1����M�9���m �w�vm���wxT��#��>��# �{h����6�):M�p��/���UH��0��06���#�����1'����TF�7^��{�.�+�ۻ��w6��w1h7I�j�4K���ym�� ��x�	RS�}0dn����wu�8�͖��V��V��}�Ym��m�$�[l�I&�� �Ab�`d�[-I7�8y���{;�N����C��(P��:�ߐ1)�Cߚ�7�?}DC�a�`"Da��F���]gcX!4�i3���҇0�V�O���h�~���6p����@��y�^�!ze�}I1V��bah$V F�R�z:�����s0 ����u#
'�!����MQZ��LL dgì�� {1�b�RB,�+_*�8f`���m�[�̘eG��>Y�^yM�4VUwI;�Y���$��m!�P��[C� �뭱W�*\�g��v�㢺�C��,��9���L���u�]�ez3m��;D����n'����|.�]ȰO�Lس��r�a��r.���U���������R⬕v'"n�(�%�<����$x����1�8�%���ۍ6��Ev�͉ �c�ay9�=1�`3q�%����e��iE��� u۫!��u�G�eɹ��p'kuڮE5 �F�\nC��\d9�`P��n�]�z��.��l/�9!6�������sۍ1���;��q��[��m-��Տs�>�n�{$��o`�tm�b��U�3����r�� ��A�)����id���c�m���^tOF�:�um�=����'��8�"(���"'�6n�fT2q�&7"X��v�K�dvܹ���5㐨�k�u���N|���s��V�gB&h��a۰�uE�q���:l3#�I��m�2�[l����0=�����-��PX�m�b܉(a_g�]Y�����ó��5��cY/Gg[���y9ɬn�s�.�<�<���[���(���WN�;����Ҳ�&�g\�Sv��ҷ:�s�u�S��A�n����v*c�<��v�L��ғ��;�XN6�#ۨ;i3���v�ւ�Z8R��;7^.x��nK8);4b���lk�#�땝���,��pa�{e���I��,Ph6���0����i�*��I�:���ܾ[M5�1�5"�-��w;�����d{[<�l�Qz�
�wX�[V��Fu����m]e�8�V��0��2ut:�]s���l���d� 1��i�,�l�v6�n���u�m���v����#�Zᷛ��kd۞:�%��+T��� �����/k�b
�*,�oT�ֹ�S�-�m�(%���lb�۫��ĠݪoRu��3n΂��z�G
���C�F�,� ��@R����t�x�[fν6��m��w�������d���H�0��2���_�T>�*����P ?D�׵U����E<;�DOAv�� b������f	)���V���岩+M�k��-"T.�]�$�N^�܂U��u�e��q�:u��طA;�*\����ZګsN��R"o'l�!I�˱��ڕ�d��aP]en'����z^ѲHd{a��慰�%�����é.'�k�Y5\��eά���Ge��Z,[�.۴��[���*C�<rC�O���SBBd�(hƲF�p�帱]+�[�<@f�y�8�ԩƆ�6�I,����"w^�f��t�����I��nQ^��[�7w�}u$����ܾ ~��.��y����YގF�H6����$�Ez��L��\�� �58~���M�}��=�1Lã�̜�������~��M����S�}����+)���U���� wse��0�9�eՁ������m��&&��
����f��O# Iy�م
Z�ؐ3�]�� �grY�&o=g�(�����)�=�8��̧�b�a��G�qj���h�7�Y$��G#��C�ߝ�}�V~��Q�J�p�&�WJ�Àw=�.��(Kx���9���������w`n����fc�N�&�:R4�n$�� �'xNрo{h�FJ�i7�$�� ;����م��za`g�w��L�V����i�0��F ��� ��x����s̑����x&��ضȒ�������gmq��9�.Βsh�d����u݊�O��ـj�{�4��͐iߌHĐ�+i�ƢI�!`s=�����W��?O������=�L,g�OQQ�������@>i� �����ȏuDA8���	�v� ������U{�>�8ߵmkT�*)QQ����i`w��0 ߒq�����`S�TT�I �"�p��dӼAܙ��[���E���{G�%m�$��%3�S���7 +��J3��0�:O���6ݝ��h��Wg�r�H���g �s�W:����l���}0�;^Գh��:���Ns�uu�������;�l�7佺\PI3�DQ�P�dq��M,t��¾9��� ���7 U��G����ܔ�x˙>�~�;-���Dw���� `!J}0th_�`�f�s$[(���)��� �XTQ��X�kx��A������+�+��7�n���,�Ç��# �nD�{3��幮�fM,w��_{M-r��%D�H%2�^xl{�Ses��Cr�0<��,�f����v;.�{�?}�N�D�RHG��Q���3&��酤�ff�:�����jR���*I"�*���JV��Lr9#i�a��L�����~����{"��jTp���.�6�F�'�z9���=>~������dt���JtH���w3N��	�?V@NрDr8�VF�F*p�����q��� ���aG諾���}�GV�;��{�/��x�B9Ϻ=�I�,��t��3ALF;e������ECf��ă�8LKtC�F��`{1�
�풓u�v7F	��/Y�.w2urޓ���� +ؔ��w5q��Ν-�쐖n�����:ی��5�{rsf��E��י�lɛZ���A+�[R����T��hyr��=�t�x�������ۡi�������m��n��䬭J�,� �����1_8�A�]��u�x��K�;���g�7/D�=�wXvٺ!�Ե7tU�$���,ԗ�;�.�``�W��""#�=+ެ�R�Yʉ��*����0���u\��Uy����TEr�.Y���7�F�۩����� o�e��伳T=캰;�CM6����}U�J���s�4�FL�I=���?Ύ��V*�_O~z��Ý��o�=����	�����'2��Pgs9;u�]�z����l�mSgJ��xF��7'V�M�(I-��ͺ�;��� ���r" �np�WQQ\S7h�v�R]���ßߌ���:�0;�:P�W{��}��5�~�U|��~!����=ʨ���"����� ��� ^{���}�Vw=��� �Y�D�H$�I��_纬��u�A���p
���=��*��*��t�\�������|���}�� m]9�#{B��5�R3��mvSu熞��Kķ�@ph�5��\+R�1�����N��l�w�.���n��nb# ��Y�!,�R��cL$�>p��/�W�U�NԞF����'�� �x�>��)��i�`z������]Y��{��$`�(�1КBEӢѥ	48`A#)���� �B0��|���������e�ww'[I�Q�BIn._}^�ב�}ާ�֝�zz�ޜCwRTL5�N'%X���8�U��;�uX���Gs0[T�Ҏ�%H)Ӕlr�׃��t�]�i<{h]sa���M�/:�[�n��/�iG8W�]���`W{�]U|}�� �+6�Q$��BH��=�g��¬�ټ�^�w��_�=H��iR�MA����mՁ�{7��ۮ��=�XՉbc�d�F��mʰ�搜{ټ�^�v^ɶ�y��O��X`�	%8��D�R����TBE΁���r{�������%�H��I�9�:���꯻�5X�{.�{ټ���R�A�DC�IT�6g[�{Eky΀+F�ms����-�y�nێ�=aۈ����4�w@g�j�;�eՇ�xɼ����n� ��0N���)�ȸz�F���}�� ]��=��Ls�*ݍ��)�'p�ۛ�� �e��{���}�Vp�6*NJEA%��^��������}Ց��r"#�{sw�~�j�_�D��I`g��ps�9��`��t�i���#}qG  ��F � ��`!�� �#�vݷ����߹P����`�M�����P�:v��Ӻu�8q��6q.����ݓs��֔k)h6rj�{D�x�s��y�؊��n�];���jy�	�<f�GiƷ\�r[���낙�:����zȌ��(^�7l0���:^��.Dmk�'p�m�v���sl��9��6�δ����ɱu�r��Y]�n�g�A�r5�=.���u����T�I7�*UJ��a�w0�f�8`]���H�Ef8�VF85/O n�Mn��g�s���y�q�kk���s˞69�UJ�5���7�����{7��w]�U������f&��R�ۂQ:��z'��;>�� ���;ެ������2F�LiF'$�p��v�78{Ց�.�=��:@�b��r1�I��纬{�u`g����V� �׫Z6��R"	��\36� ]�{�}-��i��>��U930*u�<��;nݝd�m`���/=����0������f��L�kI��&5+�KMI{��t��w�w�np�������ӨL��Kk���Iu���ˈ�F�D�/J>���uZ޹��ב�w�Ow��"d�H�^�ՁDۊ(�~_�+��]X}G�����u{u���@�j/�Jt�� ��n���������9=��N3�tꊇE�M�U�7UW�	�W�Hs��s���V��z���}�VF ��/����W.i���G��e�Jׅ`w=�V�iк��۞�A���?/�:*\�:M�D7$��埿;���� �R��9 >���;�~'�5quTӍ�i����V�캰3��\�^�v���h�R�$DHd� ��{+�?��lr9�^~s���ffg�UT��ꪵ�kZֶ<?�����##,�$#3����Hf�uw�f�nB�{��[;Z;z ���da$�&��tl+ѠN��LMWQQ4E�voR=F����@F�<^�D�Ԏ��=��9GDl���͙�b������c�]�ħ���Dw
��_�||�X	u�SP���A]}���30 {�Z��L�a�D�Uљ��I]��t������!�ӡ�&؄!��Ł��=a�`nH��,J�!�Վ��Y��"�^kK�2�d̘|LL~���	�z��������H(����2&ӫ^-#�7����Zg�o�,'`mﾷ݌��Z�x�Dh!�c(�A�1�B��3M���cM��;01�,2��2�?�_ �C다?T�UП��?EC�:PC�@�T;@_�+��G���f�/�=ɩ����$|{�iU<�	�*殪�0?f ��?N���V �KU�w��`r�Q�=��F�H�s�})���)� }ޫ��Ot�r۶���&�n@�S�;dòHݴ�b��[q��^�)�'�d�nbv16�$��|�U�w��aFwټ�P͹`v��R��B*Rd���pٛ/�RC�~�����i9�f~�J���/�$n	H�wټ�Y��io��{�,�h�{)ؔCrNp��wW<�9�U|��w�[�qU:Ϡ`f�Q[�T~"���������s�l9�pq�N6��6��U�w��`g���՛���}U�^V��
��I2Sd8���vvۨۍrj:��ƃ���CĚ鵟%�?M]F��dC��8ո������{5s�uf�=�qX�0A�i*)��MU���=�>��`:np�>�U��U${
��?�2:�>�%� ����;�uU�{��`{��� �F�X���&fn�ʻ�Dr{��� N� �z�����{ެxQ!>�M�E�[�: �w�{��@�[u�.�f�Dq��	!z@���2ĊD�@�m�3zE��`!���	��+l��mu�NSu���:���siz2^D$މ�n28����ǶK����xn�;Q���	�&2uv7/h�+`2ۡ����f�ѧ��	4����;ڞ��dSL��5��&nٹs{t�4�x���N1{ut��W�,mPOn��,�h�r:]��ql���Ʋ�y�+�y�����4��� ��Z��]��:�#���$�HHԘ񁹁�� ۵A�7%�2�����r��{5���{�mq�8��qsۥ5��o[����RO��7��w]���O�}�����~��?��pM���s�v[ujـ�U�	u9���K��r'5"j�n;wf�{%��������� �����z��R��QL/,� I;��{��۬�l�;YFcwQ����#��,(��o8Rn�ճ >�U�
#�@!�ɰ�����iݗ��ϝ��J�AD� ����C�E
TZF�����NQ>q�#���7G`6��@ޫ�G"#d�����z(<&�&�����;7&���5URHf A`8b�c	�`;U��6A����{�})��;qķ6QE��m�I��]Ot��L���`����;��/`:J$�Ia���g�?������'���z� ��
Y�I$l%7$� ���`v�f��{*X��y�=�:��%C�66�#�����:��+�z�c%�bJ�*��OfS�)HڢS�$qm�`w6m�{%��{7��7]�gkԍ�Bq	�ɻ',��� ��Ot�7X�X�X�Jk���(��g�o8U|湜�V�RA��9��u/w�,a[�ͦ�RJK�#����`�ـw��=�D����=yR_�Q$����f��
��U|�n���� �w�u�uu7W�ݠ�8�v�/L�z�t����Ln ��]vv�n6��S���5J*t�. �ݖ���pwvXݚX]i
��7"i)$������u�6XݚU�ffK�U_$_��o�i�I"�7$�@=�z���`I^��=�:�M����G$��wf���,{3{�_=	L@�)S!hE��GtJ���zQأ�}�ϛ꫞����&�#�\����`{7^�m���ـz9�DD.����L��TwW:���w�y�:n�k�����Oo\]Ù�FO���j&�D�E�7���8Vnɀ��L��� �zC�rV]�|����� M��>�`RW����{�~s��Q��3誚�	����:���fO�ث7��t��� q�|�	���,��46� ��=�ۼ�ɥ��B�:�0��%$�]�{�L�m�\�jT� ԕ�� �f��?g�ʹ%�?Kk����U��\6���u���8���nl ]�J�66�(�;��.���ck�֑2u6�rl�.x�L��8��n����W��Ʈ�e�u�¼�u����\
�n6X�%/#u0[�D�0I��cnkM�٨���>��ԃ��M�������&��u����Z��e ;V9+���27l�J��u��b�NWab:ʜI�jG�e�֏xù���{)UJ�m���2x�������;��\�M�hr��bNvh���v''Q�T�Op}�,�M,ٙ,{٫�۔�{)8&9T��:�l� �J��Sݹ�M��s�ɐ���'n�\7����`���=ș���:���|+�&�US$�Uq7%��UUU.�7�x������ف�r"b[n�����V]�4M��^�m�u[0�+�7���(�8H�O�
�"����|�^;��v���Z�])���5�J�<���n�.��&��@�w� J��W�@n���m-�j���d�8��-}U^�s���9�ø��>�x�[0��*��D��NI%���� +wv��""&{�~0�� �݂e�]MItH\]���m� |�3 ���Xr!w�6�|A��Q6�[NR&�	�`u�F�ԫ�u=�L�<�����մ�
J���J"�6H)C��<����st�M�sP�e�Uw���Oɝ�G�6lZ������z��S� �[�X��^c���D����y�{vX�M,��;�=�L�*P�țJ8�� =��`w�4������_y3
#���h/������s]��������t��R��`{��z���;=n� ߺ��޷x�~6��j�Qӥ#�� ���?w���| ��xz����3e�&��b^��r�a��ݹ֌��v۟Rq3�:�G�����Q�D���)��9��� n�.{Ռ�;=J���|����任�����r#�"N�`��X�g�s�}_${R�&�'c��HrK'~0�� ߒ���v[� _u�$�R$�"�+�yx�V;���W�s��:� 3�Й�!x�aL���V��|��I�IՖ�e��o�=����;�l�����5�/��׹TŠ;n��pb���e���q��klM]���.u�cN��c5�9�e�۠�w�w�ـ}?%Y3&���D�=�QRSrK�}Y�����`s����{vXߍ�Z����jU�@vz�d�$�OrdK޼�w���F!W�R$m%NH��g�p�n�����Lv��`�	�W���N�$�$�'8�n��ɥ����t��~���$���?�F$|��m���I$�kZֵ�k[B!�$fY��H"f�)���H?I��@S�8I}s!�V$�b ����)�d��HI$(f m�.慣IRd6�&Y�eaosDKLPQLC��ӯ��;� �i�,I��'M�M4�|�BJsO�f���0M�&LX��m�)I��
��O2��f@�ֱ����Z��A�k}&�ݽ��@A�W��v�a��3;,�C◌!�~�/F��!��M΃dA3��!2��֥� �*������o���&W�]l�bu�)f(�d�"ם�͉᠖F���6@GQiV���"����� ����C0�[2{#���" ���Ԏ�n��`�B���Z��ie|��XK��L8k4@h$�4�Hp���	�� 5c!ABcDx]�բ���ͪ�<����UV��0H��L$��h�n̒	�E��,�&�V%��n��f��s�=����m��&�NI�����LI����EjꪃQ�[�	��$�m��@9�]4�!�E�/]��N�y0��v+m��\�;�NY�5�c���J��cθ�:��#��cr�l"H9���61d����5����g�������[N��Q�.�`��Nt3����s[H�y�u�]�v�Bǝ�8��862��i�N&�%�n=��+5��<kq�wv�z7�<!��l�^5#�Q8�]Wc�cy3��Ƣ�K��59=)]@{��l�xq�i�Z��v�m�e��ny�\�96Z���N�3 �/Oqǎ�oFv�6�[2s�S��v�6�n�D�|�0ӏV�[��A6�&��u�kv��/��oL�l�6��k��u���:�C�d���Y���N^^z�Ξ\>ļ�Ѳ��t�^zg>"�̯=�`:.�h�ٝV��\onջ.�`�D���X�+���`��Gb����g��������u{ub�;g3�x�S�h���hr]�["^�RC+�o��]�]i�Y;BX2]���-��a̲�k����m�NL�Y*]h��"ʲ#6+	%��ݗ&�6n:�b��ᤸ'�!��e�ca�hם"Ⱥt�G53V�r��۬��x���:�y��Wn��Օi�^�m���2�cVSn���J!�J�4�m�l>4��z�\�鄇]�<��[����.�lX"�l��a�����^���9�jꓶbؘ���v���	9��6�F�0qX��M/6�5h��6���gmC���|'F�g��������k���y^�u�ɹ�m���<�Σ=��	��"����8���cj��-�]P�p�zŵڎ�i���v�;�<q�+���y#���26�l�z�!@�R
� �[�R�pU���8�6�Z�ܙ�;�;�f��x��yݑ�������O:؛a΅�yk�`�]�Ы^;mqۘ�氥�j�nCoQAQ`0-��-�m�u��=�뭤nνcI�=mx�mY�]��'ud��Ya(�D�`�0��s�`��=O���m؇��(����e	�dFD�LRW��@L~"v����P߀�-���S�DU���H�3d������6cld˙�:�!/���^)'H�X�$�;gv#6��a�9s�-
�nDyM�x85ʜb]Ɏ��4k���6��)�9�j�g�M����������^�u۠�ѳ��⭋������M���� �m��5ڮ�c��`�ٱ�i�g�-Vq� u,q�ɨ� v5��M8��ʺsu&U�}�>���{��ܳ3�cM��Q�J�
�a��G9�w�n��^#���ǬMڷnۋ/OLV��R�� ������,,w3y��e�{}��)(d��dWg ��u�o�=����r��0;u*�7E(�J9���o8�n���M,��;0�6
�HF����p-Oz���l�>���z��D�����Є��9%�G�v�`O�Q�7]��o۠u��=�=3^���Quɢ��9��s��w\q4�y�Z���v|�v-d��n�ߗt�cUQ0�RK�@ś���f�qw۳�u��4�;^i
��"Fģ�o[�E]��{��H6�ب��^f�]�������P��ַ� 5J"I'8�n�
=����c�;�f�W�iD��㎣�8�I`{�l�>��� ߒ{�u���s���R�Jq��m��<����}_wۿ�Ҁ�~�,{&�}^�uHBlq1���m�m@��ˈ�N.'۶��x83�x�Ob��F|���[��IT���v;���}�� �S��l�g���z&B�*��f.�j�@:��:���>T��Է�>��[t�HJJNI`{3n���UZ�w�Dd8�G#������ ���ߍ�+YU5$|�ꪪ^�7�%7�� ]N��<��}3$��IwTL��j�p�'� ����F�����6��ʠ���u)�At����A#��[��n�JER%�
��'��dsr��)�$���l�9�U��~�`s����m(�؜rS�D�	�`{�ٞ�s��D����߷@�N�8��elDMJ$��dWg ��aG>I��DL�?^ ���ȋ�U�]��]��Խ� ���I�`}��'J���At�wߞgU{�˚�j��D�8���{6X��V1���fo8׷P�]LhqК������\uA�E��m����P�÷JC����q��Jn����ܖ�6���?V+�������l�7�K+i���IƁ�Np�Otu;��*fz"*��HK��liO�qX����{6X�M,-s�xX�ѣߤQD6�$�s��l�=�X�L,?.�j���殺~�Ї�F�I$J�NK�V�~� ߒ{�u;�"/�G8���ߪ���8gC<6��Z�g<1�]�_;���������pc���ǉ {k����9��i��t�(Er�[.˽�t�:�'h��RL������EO:8�T�u@��d�r�F�H�n��p��O�q�Wn�L��ms;kd�v��]�� -�s�8F4v�`@�����m�����,�5�cP�тw�l�:Vb�wIWS�+q�쉖�(�LW���T�\Ck=N�u[����m����v�D�ѵ�E�<�;��Fy�s���o��nk�j���@Iߌz���S��:�� �>1Tf9L)��9P�9��� ��k��36��w��RGt����I�@%B]M^���XZw��oݴ`�s�iZ�HG*4�7�v{&�>� ���@�z�`��ŖIe�U��V�5u=�>��XJ�ԗ�������Ї$�Ѫ��r�m��݇�X�M�s���n�-��m����c."�liO���;�o�p�f��ɩ��A�<�aG���癩&�"$��}���y�5ށ%
��S��O"9�,�v�﫪p]Ot�
$���RF�	8��d���_�a�rg柷H�~� }�݅���wDrB+�\�y���w�<���vfb�X���K��
qF�����o4��� q%L�#~� ��IU؂����Yu�N3�7-���'3���.��f�뵮4cOew.th�n�P�~?o�z�`	'��oݴ`}?$�t�}��K�$%(�"q��q#3�K����ԓ�i9�DL���\z(��������4:~�ROtؘ�8�� ��
F���"�U�(�l��XB� I�Ͽu�3��~�?q#ؒ�Q�1O����=���XI�`��9 $���"t�	$��W�]�Y��N�g������8/�Z�T>"tۢ��(��2�z�/g[n1�V��ڜ)sٸ�z���t�&�jBHҨێ�����y�����+�j��館�n7)�����A�y9�2.����X�\X;�T�t�DNH��n�j�붑�ɥ��ɉX�LC�¤D�B���I�D���k iߌv��G��G�_U}1�p��n� JHq�$� I[0��Rot=n� �8�����<�V#�{Z˳\��B��i��z/i�L��g�����3�k�x�u��z�l��� ԛ��[����䐅�Q�T��qXR\��������m�`g��X�7�H�H������[� ��;� �]S�jKy�=��8��IUq�ꥹ��0�9�5GW�@s�� {'w2�$iȝD�Pn<�`s=���{�R^�ߍ5%�0���{lrJ�TnM���F�Y4W7W')v[���������yɊD,`���z���v�yAi�l�M����p�3��.��ѭ����A73hkZ�<qۺ��s-���!�G�:��K[� ��n��?7vJ��
\;j�<=�U�)��U*��u\�NUӵ��.r[�=�{)�{>�sΜú�A��їl�vf(ꣃ��?f ��$�ޱ'Z$�j��n�=6�u��������*�����ޤ^�<�/d�bB�.j��z�����7X�~�����q��V~��9B���� }�� !|���uN�����*O"�-� �Н*q����~,�uN�3�^���^���&8��b��N.C�n<�`s����{��{&�~^Đ�2Tm�T�ÐW@o�=�i��;�l�k�p�fP�̶�wIq��'[=��Լ;����Z�p�����k������bN���4�B������'�`��8����q7)�qJYe�X)%���������+ I�RAdF���#��-���z��z�g�#�2�Q[��))�nE*+� ����9��� �=�dKٓKՇ���!�����r �����{Ӏu�f �^�`w
��D���QҎs�o�갣ۓK<����s7�<�TuN�����\rSۻ=.í���in�6�+��nsݦp�uN���CI�S�JrE`�)��uN@|���i��%èJ����� �y���7�|�U���i`Đ���t�)��V;�������u�+I.��m��m��OL��Ni�5����	F ��2B�41)�q�PT��ӣ-	�F1�Q_>ܮHDD�d$�JA-2�-Ȯ<q$��D�/1ڐ�<4�d�h(S����Z0��i�d�j=��raބ2H�	���%&(� ��F��#MF�����"�-ٴn���%����Y�A��3�&�S��I=r�X.�
&���*	B`�&i�-F����3*(+,æ�0��:74�3n��f���22��$�������z�Q��3$p�2�&������	�7�Bk4�ᕘ=:ӹ$��!PĉMˉa�A+��.ǣ��kE�M�6��6�;-̴a$�	Ҡ`���<�:Uؾ#�U�؃)�v�0��'`��'�<	UI=O�������[�gUy��u� K7�q�"E$� ���v��K<����s7��ڍ%�I#���ێ�=�{��H��U��n�8�n���Ҋ)"$�qЩ�*%"[�����������e�A��Tk,��D�Q���Z��ܥ���]��hRs����z�~DF�n��\H�iFą�P �"rEaGs�۾��L���V ���uN@/L%�}#�����fM,��?b�9����Eb��UlTԑIs�O��I�l`���Խ�#�؎F���b4�@H0���>��9\���`r�{���?R%�Uq�4�9�7�=�i��:���7��A�i�!G$j�J���3��N�C�98չ�3��a��λ��ƌ`�m�yx��\�Ԟ� �M�ԞF �]S�'��k�EN�(	��|�U����3_�0j���ޥ�܈����]I'�NB�#��n+3]]�g����_TG"g�?n��^��}����욻���9�5I��$�t=n�=���o*����"�"
�P�����~�z�`�y.�T�q�#�B�K��0AA�}�\�[��e��z6�;,���U؋/P$�r�73a2�j���g�e8Ӷw+�ݸ�&�iӹ��؅N�f0����뛠�,����۶�˂Ό\m�N�km��̆K ����[�Ճ�~ɛ� ���kh��a��^�2i
_8i�r�:��\�*�>�٠\�=��������r'pF��Ԇ�[]�h5ͼB%��kq�]E���I� ��˷S��dJ�����5u�n�9��v��-��.ӳ9m��ݲ�qy�A����8�Q���?ߗx��6�`g��X�f�u���(�t��.n�p���uN�I�����Ē͢�j*���\q�
9��� �=�`{3n�1����MM��\�~Ds���~�@�z� �O# �?b�3p��QIR��|�V �y�uN�'��'���#�{v��Q�1۷g*h��z���wZ;u��v���O܄L����Rv�),��J�%�����.�T��{��9HyW�8�B���Ijd��Z�Ӊ��������#>D�X����� �yЀ��	�j�H��R�3��� ���`o�n���+�4ͨ�s�N1�R�C���s��^�`^�G� ��� ]��{̬T��Q
C�I�X�۫v�� ]�{�>�s�(hs4�(�|��ۄs9�m�R��%�����G ��qnO<��k �nҲ�EYF�8�����jd]�{�9M� >�q�l�$�Ԋ���8���x�������?c��X�q��.�T㈎r&G�8'����VHI7w��{Ӏ|���ˁ9� T1����Q��z��uW9�~����h[B�*m�㨛��?|����U�۶`�W�@�����,����H��p݆���o8Pn��`w7n��o�ur�M���2O�b6�YM��ַ!ɸ���V���B�]�������S���B�l���@�O۠9m�@&�0̩���4ͨ��>�)G9���Y��r9*S�d`۶`ޯn�9�$j+U%�� �u!$v�]X�рoz����`��`N.b�(������G9>���8�?n����>�^c��0sDc���i�7�ʰ:��4d#LMJ���罛�[u�&�J�N ����n2��$!I��P��D�e�)x�tG��h�m�Z���;t�&��})�9�Ԝ�[�Xnف����J���'RC�(EMȣ�ۉ��ۇ��=&@{37�V� �t3QD�(D�8Gp�v��:�{�{��DDL�|{Ӂ����;Xu�R�4�,fg�p�˜�v�r9��`�G�b�S@�A�M��> �{�����[�/�6�R^�w�Dr#���Yr�Kөi9N��ڌtiR<r���@ӎc����1�#�i�Knݎɰv�dd�{KX�u�m<�loKmvyn8ݔF��Þp�L�i�vnx��Ŭtz,猊��������P�k�Fv���h�4N�)	��KFN �}���w��lM�q<��XwŞ"�9t�M���� ���9�qlWGc�vn'����[������q��B�p*_��� wݽ����ی]��7&�1����[q۰2�y��T��9��覄&%'�N��E�7L,Jр|���G"9��=��� ]�~��"�������l�L�m�tz���36iu@qfRHC��F�&�D�t]Ot��V�%p�[�Ҙ�����v��7ri`fd����o8sj��)PM�GM7'�ləV�w��t�����5�ª6�aN|ۈ�#l����ݳ���QZ5zcs4랫���_k�a��u�/�;f ���t-���L�;Xm�hC�Ӑ�3���2�Uq�o9y.i��U� ���=��s�2o�ڟ�B�)�R�Sl���~���,v�%h�z��
E3-�ɒj`�����̴��V�w���{ެ���ދ�\$]�V�6�]Ot-�2A�l�=�G"W[*'v�T����h�:,�i����O�������m��q���c=Z�]�o��Oۡ�n���g`��Xېiϗ��Np�����XܘX��� �mD���$����i���s���}�~�_ ��
&%@��� H��� ����@����&
��9�wik��Nr �����������&���l��f�
Ru���#��D��<`�榩�I%]�5v`	u{ts���Z�������s����R(����jTE k�p�{\dݬ��#i7\��������^���y���GlUuSW���`�`��>�'"�-�mR�F'���,%h�>����)I�z#�����̙�\��"�'p�;�_�z����� �zi`uw)$!��)Q8X�7�@)I�]]�h}�"#`�8DGت`k�OSH;�y˺����\�����4��
Y��g��3&37y�<�+V���:������Q+�Ļ׷�vu������=����
A�;��=6�WDݗ<&n� K��R�`�{航�[���w05��HF�F�$�4��`|��JN���0�,M<Qr8�)!`w����3]��l���d�����(u��q)�F�^�
Ru�}�l�R�`}��@RV-{$hCTF����iV3&{�Ӝf��R���$�[m��zֵ�k[��!�����*�*Jo�+��3��h�2p��5�a�;tbɚ�*@��P�3���]��k0��L�!�d�Ku8u+�RD�D=���տ���I�
v�����E1�QVۮ����=�Uټ��f�耊�������(\������MU��N��ET��gY�bQ��5S�&)�ժ�a�]��ϙ��ș��-[����lL2й�,DEC��Vl���C�m�6Z�	|/�[p�r�ȣ -�jH�蔈�.��R�ɰO�;�{vES�4�$e����f�+0�")�Uw�R�j�ݎ�&�!���H0L1C7nJ�aD�5F�刺R�; �Cr��)C��330΄�ߡ�� �.fD'�8�m�/���$� �;�W��!����-�㋫�A� ՜/��E���w��-A۞P�;���\��uR�=�}�o��>ȝ���Z��*�t���ӹ�k�e���Փ,HѮ9�{g��%d;V��]N%�t[��ج�����'�۱6˻d�֝�QĆ�qt<�X��i*���;�r��Pg��c��[$�1ɝ�cn�a�� ν��nP���lV2�l��G�l�'c�Ub:���6��E�is����m��m����Yl�w5����Cg�t�1��� i^�	u�E��܄`͝�3@�ʜ�xwX�	�y%zKq6Ƕ�<�8��v�av�x�#s���:-�����u[�^�lc�ewW���u��Փ��:���q(��L�h�Vψ��JhVX� �5���E���:lN��4fKw�s5s��:��Ԟ���Gg�%��٣��#z�q길�,���qv����e���o[���mp��a�'p �ؘ�w'R�4km��3{�8��n�mK�H���Q���`[ql{c�;c������n˻=la��NAԫA�ۭ�&n�&8�m���f�0�-r��3�u����c�XӜQ�;�v/&%x-����-������1Vd-��-������o��2b�=o=/ZNSkq�Z��~
��%����FI�J_C[n�s�dQ��Q�,���Mlu�;B�[U�a;a`���KM N4:奅�`��lks�8-]g�K�M��[!��}���c��j�L$�>����3�-���ā!�t��h3d ��;F��&vOisl�Ӥ�u��S�6��&�6��trx�xݳ��Z����m�K�o<q�W����؎qɞ�=&kl��yy�`�QΊ8��[cv�q��Z�L���WN9��8�O\er�s<cz�h�[��K��sŚ܂[�ͩ�@����Lp�	�S������]qfJ��sp��v^��m��:�'lp�ӡ#8pFӜ�m�Uwg��A���e7$gl�!כ7�v��~ݽ�6�ۺc`�"��7g6gc�^R����͟��oF�NT�@=����/�?�) hP�>�~
�b�����d�gL�fV`}�#�ۤ�"KV��u"<v�2��Z0�n�iT�E�.۱�c=mΧ��j6&�mY��L�f0ے
�m���ګ��vq�Qpkj�KpN֢wq��iXM�t��w��o���q�]��_=*��Z��X������s����9��=�񍕪�ۦݭ9��{9Ό��"ʆt����!��vu�J9�lV�!�]�I��3�e���7��+���8�qC�v��kz�X�^*x3ԋ6��d8뭴g�׳٨�5���ـoퟋ�;����5�͚YA�ܤ���@��*'.p��{�9m��]� ԭ�'�~�_���BP
G'+�j����f�3&��6�sj� ܃T%#���i`w�0�;��� ř��7��3\�)(�Tm��8wf�{�{�)I��]� ���� $�ɀ���4ӻ�(�=:^�8�v�[��h��8�ϞbU��T�qDR�2�r�����'Q�}�l�5+F �㬊�74X2��/8���{����@fb��\�q$!	Ѥ����/�v|뻺�������g�s�����Կ~��&�(�bq����jV�� ������`��\�T�f.˩�4=�����z��4):��DDD�{<F�뉙uQt]*bR���;�g�pY���٥��Ʌ���5j[*5U���R���(���eV8�=�λ/-յ��{n�հ�B^}�8��A�% ���b�֭sfs&�DF�w���;�b_��*�ʉ�f��g���Drd��fޯ{t)k��$�}�kh���۔��dw�w�ꯟ<���z�� ^�r@�Dr".#�Dpʖ�Q�5�F߀�ST����e4�,����f��٥���d�����m5�$H�s�JN�r"#��l�>nـ}�|�@����s߬�[����2�\tq�˞�����\]����y�vj�\Z
��KQ5u�o]� ԭ ��O7@N��V��#5R�Y��K��o8��,(�i`�Iy�XEBR�n.n�ﺞ�I�u�0J�`w6���'HjF��~����߻�y�����}߷U���0|���;��u������}�_y�Y�Č�D�nAҤ���k�ק �+F�I�!'X���L�5D7+�^z��y-X��v{nK��;5�l�b9;��쏪)�\v�n��(�'p�݌͙'�=����[0��TJ�Uɚ��*j��7�=�G9�DDL�o׀f��U��Ʌ���ߍ%6�d$U�$��?%l�܈���]� �/{��LĶE�A�nK��Ih#R�`$��I�ބ8�¬�"f.˩�4��f޶�@N��7��Z씈%�_ c]f�2+�jŹ�庸.�����sۦ�S���̬�`^�6�)���N�'�]��f��wX��m�<v�́c��s�^�6ٸ�t���ɹ� sl��3X��aۗj�ݹGC����J��Mʼ\�G-M�۱�N^p��*[�lR���B��v2�c�����%�d�����x�����f�!͆���Q��'����F�N©iUc�� �"Iﭻ�X�+�����;�A[:�����3nK��딻��ƀ���`.'h�	{�t$� ��F�Z0�0��UA8�C8�8��/��}T��߭�T���0���}ȎL�G;���S�)*II,(���K������ ffˠ�V�J�m�I�w�v��m���$��{���%w��tK[�S�l�����~��
36XݘX̘XQ��T��NQN����퍌�qݵ�&����ѣA�������:c���j*J(�Ns����۶�RXWS�>Q@����S*ڜ��K߽-�32``�"]��G��f���`w�^��4�HF�f��v����D������`G�FT��M
TR�߷� �͖o��3&siP��Ӏ	YUW� �w�'�f�Z0�����Rm5QF�qJ�����V��5��.�Ysӻk=ѶX��l����D����2'�f��рuu=����꤃߰ԇ���n���;� �������@N�ճ ��S2���l�������p�fˣ�J.��ozd58O����o��=��X]<�KQ$q N1�� fc��v�R�`zRo�hq@�A)0j9ܗ@{vi`s2a`{��� �36X�ku�]�&���J(M�mg:-�mk��Rm��Jq�7�Ŏ[�gu�ۮ�EN@�E�8wvi`g�7��fl��L,�#ͣ*SH�#�U,�Z{�	'y ?�� ԭ���E'OTi����flUh7�0�;�0�3ۛ�ݠz�К��LL�]�z9�D���`7l�|��_=`Y=~�a�I	0�����qN_�`��?|=%'H'�p�l�i�$���рoД�D�s��:9Ƿo2�#OkoBs���&Lӎ���[�WGO=	���^��f>���4�@N��h�5+F �T��pT'�s���������d�����s��|��I�	DDr�r]���p�y�� �w�uv%��"nj������ $�� I;��9�G'�y�N�t<��\T�uS7p]ـRbo��=���{�,�;�������S�U\ٙ�-�޲��\X���J�VX猈B\WE�s۴n�[hX$��l��۴�A�sm7*�g����ڲWm�+�z�&ռ.�1����mEY�����gW��8 �����v^q�v6�������s۶,�9߷��|�nŨ�9�/i�f�\��\'Lq��k5�y�lx0�R����B�!��ܖ�[^��֞��4p�K���3l[�	9$��j,��ִd� s�nn���8�&��\[ry�]����X�)���P$�p��%��Ʌ����] ���p�-oA�� �fj�@iZ0��'��@:Ӽ�H3�H���! ���8{f�f�w� ����za`{�D�����5sDMUŘm=��� +F듞��������H��u$㨜� <Ӽ��~V�u��BM����fc�p�gn���z�T��ey��tm�v�]O\Oke(�g��+�k!�����=<X�˳����?��*�Cw�����_�`ffgp�|I��>|ﺋ�{��W9��u�~�䌥��m��JH)s/۠v[u�jрu+F�a��t��P�H�8���aFn�,,Ņ��Y��~� ��?ߔI�Ғ �6�V��D&�|��n���X���+p����"��ZIF�#����N�7C�4�ޫ�lr�}��y���:���Y�&� }���
[s^��~�g-�lkg���/��7y�n�;�0�=�X�1����u$�q�pۻ,��,�����ZI%��$�I$�J��G�d@7&z,�����-t�B�q$�0r�2,Cm��������@*�0��ȓ�;N���[��;Л6:��G�۵v>���I�|�31
�a`�:!���g���L,3F/hq�#ůi��R���ڝEG��Eֳ��6����5�Y�5fDP�K���J��:�ă�Iy��E�`���@���^�;՘�*t�c��nj7�����y��֭�K﫯z��L�TU�L��a��h"���M��>�/<���<�ދj�gOz�;�0��o{�<�l���=֊�utt���/�	�Bo�MM�ŉ��H3Iػ��sꝘaН!|%C�U�<�3�:/��%���z@b����Zyq�DM�玘�,Cڎg�AQ1�aI�=���8��``��~w�Qڂp�A�^�1E8/B�HDǋ�i^
;;{Qvv���hD_=A&���@�?v�C��o/f�`sٻ�^ܨd%?����sWxjрw�рu6�C���s��^��X�P*_��2��8E�3f��ot���V��$\D�S�������]sη�����.�`��գkt��t�4�QƇ"N�u�u�}�	j��DN�y ׈�:h�`�� 3۲������{&�wy��U${(���$�R �J��y�0��U� ﺞ�[w��Eg�u�d�$�;� �٥���w��{�s}W�=a	hf5��F6zkF��'�Ύ�`����,T�N�[��t�;W��}�ʰ9[Z�65��L������ n�nـu+F�Dq�R���b�#�xU�������B�{;�e�ۀ�-;c���qvc�ĸ䌅������n�޼歘R�z""6Au?n��S�㈟'H��,�M/�}�}T��ݳ _'��ۼ��8���"n��.n�p�v���{�	�^�٥�`a�`J��r
B��}U�I�}� ��^��R�`
�zJl%d�s���͚;A���uW���;�"�BEy.�}���f���05�v7g��`V�dD�Bv�E�q�ׇ�V�A��v^ݚݰ-cb8u��\�':v����t����
B�y�7Sr�2fM����p�rX�����O�^��ݔZ�ir���Y����rs㭴v���\+�IN��j��݈��g������7.��Ϙy��-��8zcn]q�Ѯ��Y�E���m9z"1�8{d���X�n
�;#y���a�e��|V�J(6)H,uQA:�%\���e��!�p�$��%c���y�-Ó�r�հ�����0�h����}!��x������*r8�IK���Eh9���&���/#=�����qQN�$�� ��0>�I��n�u�x�<�;ܘX��m:[BP*A�99�n�3��V������ ﶠl�deN5�����������p�=�����1��鍸��J�"c=�q:8�h�L��*��j�je*B�!D��HYU%�\�]�h	;f���M��ͺ��4���4�JB��}�5�}#�$H����:���e�Q�mՁ��[,(�n�k��	�U��$���y�V�~I�wz���8�M�,�͕`W~X��{�i� o\�5`�q&��\=�K���pۛ,u<���9�Gɲ�M��*��UE12�ۥ��ӓ��'K;-긪���w��sI����ȉ���R(P܇@�~��� 3se�W�mՁ����73@H��
�r� �w�}��0��2 ߒ{�G"d��5���������`{ٷV��?��>С;UPUz@0NDF���� ��x�v%Ê���.��*�c@M[0��� ��x��d`bHƖLiH)�9��� ��~��@;������7�˸���#" ^��C�Y�;r�F݇)qmFn��[.|��S�>��ӥ(C�� �͖�6d`]�S���}��n����J$�H�)SrK�ͺ�=��XQ��w� �͖��ZR�$�q���� M[0��{�̉�xSY1��d�%#��^$w�{� f��������H�"��)B%*Fdh����%M�'@��PC�=��n���xe�k�d�\UY3W� �w�{���j�`s����i~��ණ�"�O�)��9�5�;rl�Q��s�l5������q<L:�<��ܦ�!�����f�������R�������V��
'�諚(.������v�~I�')�ާ������H7RF����8D��q�s�} &�=�D���F ��`G�N�M�������T������o��酁���� �5I�D�M�x~O# �� ߓ{�	�x� M|,K�O�6���KR��-��	��j�"�G�V�5�6�Ñ[.�oXx�Pm�6��;0��v�;�Ӑ;8�%��\nЏlC�jK�����د]���į�{�m3a�ƺ'T��6qh�OdyN�^gf���|]���Q��v��*�(��i�4��p�%���ܨ���W`1��v��Im�u�YG�1Ĺ�%�I,qV��}��=��3fe�t���$6����r�x��Z-�9���v�ϏKL��ݏ\�v
�Σv��m
ȢIGi)u�7�O��4�@N��<�aB�������,Is��� f���ͺ�=��X���C����R�%(�8����y=]�`|���@Jd�9�"�G�9�۫�酁ϻ���nl�9�R�ߜ�8�\5\3 ����e4�@ߓ��?9������Ӡ�C���5I���^��t8:`�ڶ%��g�	wk=��i8��.N�5f��|�� �w�o��4ճ �w~�Q6E�Ӝ\@f�˺�|����>��B�d2 i"4��:S�U3.k�Ό������}ș"�~�������������~��>Jрo�Otɑ-�z�nL����(�T�R�{vi�}��� I��7��075$�D��HX���n͖D��۫�酁�a�T�N�(��D���tz�lj���v:��^��
N�0xuF�]qy�\�8'�%(�8��,w6�`w2a`w����`-�DU�B7%�WVn�ht�`w��$��2u(�x"����Ɋ����~0������P8���T��s��ey�u`y�XDF�j������8��,�6���d����!-آl�sTQSw� �w�z;����0���p�}[��r�)&ی(���"i��3��V����$��a�Ëh��y��ӎݶ�$�4JT�p�����;�0�9�ۼ�f�nji
��R9#I�p�l�7���M����`�
H��#S�(NBZwwy���`w��V|̘X��7O`��(�$B�{�	7x�'��|����/Q3��'���,� a`H��E�˚�"C�J)�>�������D�E8F�=�۫��~M�$��q�陏Aɹ�L�r�$�\���k]���l�A��Y�z�&��^�0m�v�#Ǆ�8țQ�S���3����9��� 37e��ͺ�=K�,%!D�U!5f��{�L����8��>Jр{r���Q�Ec�� �ݩ`w3n��L,{ۼ��f��I�".&*h���DD��l`	�f���� �ݖ��M!-��#m%.��m��9���O���U��Ց�W?��x����QQW?�*"��gO���(2��m�[�":U�@R�A2��`E(AR�TZQT�jTBP��DJQC� �@ �P@0!��D �RYM���* ,
"�*"�

D#Q(
�D�.�Pp�@(�T�AR�U%!DbARdU&ER�)@�X ��eS @ZDA�D{EP���mu~�*(�H �G�k�������eC�5A?�?�'�*	�"��(����*��'��L��_��	��D��?O��UUUUUUUUUUUUUUUUUUUUUUUUUUUUT45UU�A?������A'��A?���}O��@����f���/������G�"�����?�������QQW���QQV�����=���C�o���?O����~����C5RCSTSU�袢�����������o����|���������?����5��?T��ኪ�?�k����'Z:��!Q%HQ%FTIBI`�THaD�`�Q%H!D�P���D�Q$�RYQ!	Q eD��BE�&I!D�Q$�R�TIaD�HVTHQ�TI�Q�AaD�eD�IVIA�Q�T%D��T�I%�R	Q"TI%D�I	!D�Q&TH�Q&@$�Q eD�`�%D��FHYQ$	Q!	Q%dD�I$RTIQ%%D�FHA�P�BTI&H�&B�����(��Bd$ %��!!B		A$ PIQ		D!%V$!Y	BD��`!!!��D������B I����`%d$	BR!$������F��d @�HHU��BQB��E !IXB	 !BP%%%	 ��IA��a%$	RBBP��dFBA$$Bd	d$ $!P		DB		VU��U��T�%��Bd	��Y	T$TIHUB$TT��DI	DV@�����P�	`IBBRB@����HBE`$�! ` !	��BRP�$`ID!!  H	DXBFYABAHQ�!` e! (HB�JB�)B $�$� ���!a���F�X	 �$ed�(A!!	HA�$P�B		�K�
�(@$� �@0��,	"H��J�� �� J���H���� HBB1(CCA � 4 ��"̪L��)��#�"���*$�*$��e��������~���B�(�*�\��h>G�?SY���=p����������TTU���3Z���~�����à�_���7���s��?X B����u���(��*����TU�������QW�;������mTU��?O6v/�9���<�ʪ���3���?>N����à��|c#?��C�?���EE_�?��	�o�9���D��}pTTU�=�H������ 	��[/����1��3����O�������}ӟ��=_�B�������ֽ?Zt'������ ���Ϧ|��ǟ����ʢ����|?Ԫ����G�ϊ�����#���w����������b��L���"�L�� � ���fO� �
� }e�4J�vul�U���]�6 ���]���@ K 6M^�0@�ew`�v������@ = j�5[j��
 �� 4 �   hP�h @  @@ @ (�T �    �@��e@�Ps����=���sjWms�B��B�Z�j��p��޷T�緪����o��A�� @�w�����Y@=��I�=�9�^v��AA�6���{�{˞ޏ}   =��J
��e 
�$�s����}� {�t��: ����7,�(���ҁu�R���P�J)���N��V��4�8� tv�� ��(�k4� ɹJ �4PR��J�0���t �AI�)@���;:PR�w����)A��[P���� ����(
����o��a�������uA^׀s�a��}<�@1�}^�<��{  !�����8����	������a�=n�j0����=70��@v{h��*� (��g %xOA�a��tȡƤ+� ��`s��r;1@� �9!��P ��as9��T=d����:��m���6���u�;�z�{w�z  �! �ր �@
nn��c���/^������Cos�'o@�=��w��`z ��-o@�0@= 8{�;oop����� ������';��(�8ow�=�tw�8� 0     �S�&��)J@  =��*M��  0��U`S�j�b�SM�ɐ�S�j�d�H���jR��@G�z����_�?��������3��>��k�@U~��dQWJ��dQW�PE_*�PU?_Ϯ?�r\$ ��@�K��)2�����-7l����I!�#"�1��B��&�4ZT���]g����s<&j�!n70!L
�����I,xm��Ը�zK�rM�B���,t��5�r��.��p�+!q�l���E9����]�ˮ���u��4d�C��3a�[�l���*h�n�A~}��J3⇠��\�v�Oo�<��K��'\V�(�V��Z�N��
(:^!�S�ϗ,��G�`a�����e�a���cI�X��a�����z3��J�w7z��d9a�/y�O��3�;��u=�kڜ؜�	Rq H�bG5 ��\��o�=���xa���3q'���h��h�#�)���b��a�o�s�fG{N��R�w+�S�mwwKu��J(��8ˇ�Ip߻�Jc=׆��B��)n�$%(z���ѧ�a����� ��j7̄%+��X\42&���/��޷�{{��{�.�+��w���-�E��>r��沝mQGn�]�{�j7 ���5�����/�z��(p��}ܫ����fw-.�9ZW��ߌ���$4�캗Z$�K!`Z�had��!��
F�Ʋ�%1�
č����aB3Dj�Ů�Ͳ�R6��##@��0#HL"5����l.0�0�)�l
ԁ ������!�HHatl8xzR=H�$4$\(lx�H��0��7���Hpӽ���#C`�,K�Ѽ8��64����L��,D��XS�4P���6_<	s[�����!Ltp��tF;�%q5ĂA�;�^������ZJi���/�^����gkٺl��k�����>M�'�f��[y�]s��GsM�g��Ѹ�^l��=e2���I�\���0
]���k;�Sˬ�o7�ֹH��~Vo�Á��p������3�Õ��KwC�ʷkMBt��vs�k/�G/��W9	K�|�gK����%����&��9�e�7w7���x�5����Le�B�	L�0�0�BHR����p��(���zR�?��X;�(����s����5��HG�����9��<�)0��'�ai���=e	��$g��<,�.�<zJf�L!q�!XV]�!��<��C4�㩛!��JfDth��XZ�}e0!Lee&Q�v�g�$�津g��s�*��'�q�/���f~y�� ����=��mv�|*�c;���rΟ:�:)X���r��c����?JJNCt�뾢_;�5Nv�[� R�]�EY��TR�h��-�[p�HR0�Ȑ!�¤`F�1N$��aA�o/�a\$M���~��120��:}x��>�ۅ=>��!sz�<���ZġN(Ua���[*�\}L:����;�^���kw�ݭ��O>���J�Nt�oM�WҺǖs�}y��zm�U"�+�͝�ڨuc�Ц�2�s�j�y������>�V�����{c�}�@y/����%�����'����c��e��g7�:�����}�k̈́i
��`B$	t2�&�r�vn���f|��%�&�E����i"�$�z�՜�T}��]T��2�ffwn���{K�Ffc��;ρ��R�'��:Tp!X�\aq��%ɜ����)%�,s���=g��xR��>��=��No9���3�^�~�6��S~�V]��ʼ�ٻ�^r�u�3�����r�V�k��z�����G{E+ξ����s��P��k�υq��\�_{Z����"�������;E��V��7�Hz��o{|w\Ut����U���U+�����º�ǭIi줻=���.P�FH�a�Ns�7/)��SAU�h`B�}�5������hysz�9��Ѳ	b�R�_=�u�ޯ8aB�7�9�h�Jk�GzIg�9tO9O!CL.a�KN�˩�����d�68VP�+
����� j�77=J���8��!@�"̓0�ȗ=��s���º_Dφ����Bu�*�{W�Ï����|�8Y�93��>��Y���).NQ�t�{������W=�-�<���2N	�����ƺ���e�{}j���Q����%n+��2��ʬ�7���Գ{�1��Jd���B�[���-/.��ڕ]���K�"��rAJ�;p����F�(>tsvp���Z|>�Uw����ی]u�U���'Z��]��o>|�N���as�	c	y	cB������SL�|��w���^h��x���
bB�HP�!sU��B�	�$�!K� @� �c4��LH0$XT�2���0!BI!$1X��	 �,<1��6�6�o9x����!Xz�N�$5�{�9���/8m���g���L4��Ѭ�R^s^N00�D�_���ܪ�sS�	����YIo���w�׋���N�/��ev�(�ܭ�U���$CÚ�e�w����4�d�>b>�r�֪������s+���y����}l��.om�0��g�9�9��r��K�@��fkl�Fs|����f�-�.�q��^��ėD�0�t��a;�f�l��9�9�-}�����c�)_(8�HE�X�8���2\�~8m�G����G�Y�ߟcǏ�_��{y�s͐xV�u�qr}<��K�%0~��Ƃٺ���
�%9)��p������q�q�=���Y�)d-o4g��d�돑���ᙻ��f�9y0��0�9�{�톎s>5�,p4jq� �0a�+��n�&�Q�=C�?%,������Jș�U�uWb���w�t�ǖl��噷�k����R_*w��;���x���o%�N���{}��j�wwIZ���zӔ�d��ߟNw-L�m�|JU���"^o3�����=�d0�.i{�8��.$��J�B	���˒�3��H���y͞湔�5�1������㥿|&�KdϒSWRa�'6߽�8��rH����.o�	9��B�/���o�D�e�Jx3F�u�g��Ю��X2�1&#��)|.|,��ց���0�ʪ�m���+��QUx�q>����]5l�q��>�~{����f�l��K�x��kw���>@�ns�{����hߺ<��fOu�~��n�R������f��
�%0fh&��a$e"XR�
bb������0��ņ,
(¸�acV�*�$hD�
�
ˉ(D�-4���0�d�@��H!Gg���`i���M���"�h�-�����Z��,7�����7I�0�����Y�8f�6W���4U���xxH�M��B��R�"@(�"@#
�+(��Z�2�/����w�}��]���ss!�|��]O�6�w��\�uFٻ�*�@ Ю�#����|�x�߮�Y����1�<�˫�I��Osfi��e����m���gf���֟,�JN��':=�7df��{������e���κ�O����|������JA�3�����%(�G5鰗5���XR7�\��hd
d������e�D�� B��XR�`L�XVVP�&L7r��7Ŝ3FC��&�i�[ߢ�@��w�.�{��
�y'�KXV�ЗRp7�5.����X��	<��E|�b�:j�6��jϏ4��g�������n!'{��%7%�װ����%;�K���;+��9T��(UBҰ_-X�V��V�Bv�/T�2��������uͱm"B4�<��BbC�ѹ����|P���>%�|��\���+����>���[�s�L�y����s5̇�ālіm�����Y���{l4d�m�璘h%�A�C��b����=ϡ��N��(ɋ�n��n���U�T�ݮЖm�Nc��B��>�ow9ھ���I�B�/vs�]J��y�nmo�о���'8v��wj4u�B��)]�R� ��u�]|���h���*+�Ӽ��q���ߎWh�yE��ݾ�ނUBYx�9���]��ܾ���39]��}���v�Svw���ʛ�WI|R�)�t���%|*����3�Ը�i�R�mu5Y�];ڻ��ݮVя3�>��X�+�[eѴ�"��sD�>��ng��<�6g���.�
�	c.�j���9����9��	�$�	BP�%aX�S	Le��q�p�<��4�X\�a	璑��H��x�oWp��7��យ��w����ō�C�	LbRsr^ZGWQ��ߨX��c	��m=��ۗ��B�r��EVѝox�>зy�TV�řK�]�lo
z���|�����[������{���Eڽ3s~ܢ�WG޵|{��eq�{����^wz��Ͷ���~;	s�󚔓~���|��ݔ��}+��!FY���7mHZMo��6,p�WhBỞ����ˣ[�\���$�L��e�Å�����N<RS|��$�'������|���S"A=8NY.�u�Ng8��$c�J�jl)]n#asL(B0�Z2�Hp�$��d���5X&�B�F,E��)�+����y��$�~�^k��d)(C5�p9ͻ�o��9�5	�.�˄��4MbJJ2��3Ϡy�v�w~�!|�	�ry��{%�}�5�)��L�3���Q���u��޽X����W��Ъ��J��c�\��<)�7�f������a�3d�.j�3�.�ƄR��2�K�
K�M����<�6y��z�(�~�Φ��̔��K�[�J�%	p"MB�s���Na�rB�ҳ��x]�-�ƶ���ݏ؇8�>,�[�(�m�"�E��N�U.�\%��	q�c��\e��%��SZ�5�l�i��$�-"��Q�6x�᠅!v�J�BF�	�"��SI������z��
ጒ!�g E�A���e���Y�����y�Jf���o<��vx��BB�LӾ���.���<��͙�2��K&I#�)�MɁ\�߾�.���8��$,,a.I��t�W�f��A��R�t��))k)�go}�)!�	V/�|ݾB��&��d;�HF�|?{�}�{�[In�`�k����2�&$..XL��y�[�+��w�K~��qVV[�bK�[*�e۝���Y�o�~�>��ϖh���ګ���Ϟ��sV�eo�8{��2�0e&aX{�j�����w������.|�zIa~p���3��ĹtL���i�}�6��~�׏��p���r��s�2�*����
�X������F���
����0���-��8�\�U�`l �e��L����Y1��8%	k-ą�$Ѯn�ه6f�r4��H@$HP�d$�R+絚e��Vs3ox]*���hYKs�)1U��i�u}��������}�u�g���e:���Ⳡ�s/h:���o.k�|�V%�`F\��F�!Yw����-��p��F,ׯɚ�dHY�#�=��Ep�HQ��A�M7�!���9��lѲ$�O8�b��E�2��s�W���H���Q�|Ѹf��o�����ɹ��Ӈ�l,#)��<|8i��i�s��<%�G�cr!V G4F0�Ӱ���	P�"ͺ�/9��X�������*������������
�UU�h�@j+�:��je�Q!Rlїl�1t�1Tی9�a��I]���Ul�;�\�5sF�����Ďzt>Zy�U��W��á�Ʈ�����(��"����[W�;#E}�#zSv�SU^N.�e��z�eX}W��$�:7�LH�Ov�M�j��fU"���s���\��Y�N�wf�m�!Ƨ+t �A�lqF�x����U���(����;g21��Y��Z5P���8��vG�)��Y	� ��D�����Bɣ<۬j���]�N5�sJ����l��̥��l�ꗫX,�N��n4e;�Ue���j�l�
�U��G�;�x�*�A�.R�^5��[La6睷"�b�;�n�V���^�UJ�J�J��p����&0�z}�Α�Wh��-[\�l�ۣ�� �ܛ/��UUW!��!WMj�`�h��c�a�����UG�j��&r�����eAH*��v�;���^ݐ�������U��,)ձ�*�:���L[������a�*�����[WT9ϧ�֩%�&�*�9V*ڬP��*{f��(v����\�6�X���E^i�v������'�u� .���U[P�%u	Z|��,۬S�Xz��N����m\�q;,�UVS3E1��<UQ�േahwn�OCU�y27S���e�ڄ�e;*�2�M��88֎AX�W�."�^K��n�q��֚����K`c4��Ȯ,�XDZX*�2cMeػpPr;��[��x2)Ӻ�.����m�֋���J��vj�k�ۖɎ��5�ƃ�z������T�?
;ʼͩ�4X�Q���������*� �!Sݲ�9�O3m��[l��
��e�5s+7:8��Ud.���&�-$r�Bf`Z�B�lP�����vv�0[�F��M��mOc@4��e�Li��ƈiT���"��V��z1�q��"i�*�U�Yq�,�J��]m)��=t��Ϫ��g�z�T
�mV���֗cS�G�j��.��D�,LJ���hchm)�R��W��O��˒$k	)WK[B�F�UU[K^M��A��*�X�\�۱��/��v�����F�jL�z��يҲ�vJ��l=�˔�OC���#gX�O��WT�m)'lۍ��TS����۪5���e:.�0���"��MT�m">�2h�Ǯ
�<��C�x��mT�mc����Cjv��6^j\E�5+�X�*pl�n�ZLܗ(<j�מ�策�l<���;����}���6�*V�K�n67OJ�t��Ī�@,��u��ݘ9�R�֩ȵuS��=ĩ���z���$��]UG%)�J��]u�@V��UUmU�(�������b�.ĳ�Ht���lm����SIVĥ�x\�Y^4Kb*�-�ܨt5Hmգu�q����:Lݢ[6��f
��Ӏ�`'�]�����8���J��Q�mҠ9F����Zp��.W�ZڪW�>���~�h�:��^;g2�UP:8+Jk�v��]@93+PV���­�+�~^�G�z�[�86���*����,�*��p3��q��u�e櫦�΍�vW���ҭK��QH�b{ꠛqΞn�N�8�>�ͧ\[	j������1+�08���[4��;h���A���5�U��ݫC�Я��Mn9xN�h��Ujګ�JF�vB��+ҁyT*g.��K���ms�6/��G�7T�vͦ���u>��)�	6��;K'��En�k8�P�@絠� f hŔ��γ�lm4�kviݺ��Y��n�"�6��%���j�����n��x�!�Q6,�ͱv���k5s��3�K��'n��y����^(E�����N�u�9۝e<<t�tO�J}�x�(
�`)Un�J��7溠"x[j�ښ��Egp�ud�����#�zy��q7�S�!���ۧ(@q�yw�t�e%]Pa�ͦ�ͨ*�ej���8#:�W*�U�P�תm��	�R�e�4�[Q�nҰl R��pUUch�P�R[�[UUJ�����<j�,�P���mTm*�U@=�cWO*��%y����a!@�L��:����n
�{��N��V�Fv��ch�uհ[��6�&��e��v�F4fd��^�	l�s,�5
���U����J�gz���g���L�]�:^.f�v�5�p+*�WUJ�W]%vD�J�$�=��� \]_U|`�u����^_U�<�Q̨�U���ͅ`yZ�ꯪ����f�R�UUUpV쭗����f���W�lp��S�&E�[�� +�P�UUlpUc
�UUR�C���mϊ�㸀���*��(Hw-����U��uN궪-����U%�T�@�1=���w/]�����c�=���<T�� �@tp@[mUUUJ	(�v�kn���R[�T�u)-J��]�U�yy��[���K�ҭUW�c�8�Uj �����K�1�`6 N;o.82`Z����@q��Bj�U��Z�����Vu��\�byd��9�':(,�Uur�: *�H��.��BD
�ua�;U,f\5A��P��VT1�BK*��Qj�T���ڪU[:��^Z�`*�U����^ڰmh��[�U]!5uUUme��
��
����RUPm�Ʈ�e^��P��tU�� �-��+<���U������R��5N˳U*�l]v)�gI�m@]W@�(
�����fUV�m���� �m��r���]UUU��B6KY	U��Y���Y^���WYc��j(�uV�T�������MV�WT�*�����XA]��ʺ��`�J�U<E��Ԫ��ۭ�֨�U�Q�
���*�j�'d-�=K��������YV�*�UU��nI'=n�򍱴X����q����#&�mWmZ5P���;U&B�]UU]UT������u��
����@UK@R�PյU����-l]c��k.9R(.��20
����f���V�++���UcPQ�ܮi��j�W�v庪�V����'T��UUU@UU*�UU�UUU*��UUx��*����sX,�ەV*���H�h:jRkU���5^U��T
R&^j�ڪ��jU���A�ٺ��������^Z�cb�z� UUR�U\�U�@=7YF�U�e ��%\
c�m�]�t��w|`>�u\���Uf�ݛ��e9A %Z�j���"���o v�V�/.үR�UU[.s�e8�e���n�%UX���q��Bmҍ����~C��UU*�VҮ�U[*ԦQ�te:n�TWZx^�ٟM�[�ҭǃ���ڗ�R�U�ڴ[Wb����j��j�k�kRU@R��Uv�UP)-�U�UWUJ�URpJ4�U6��K�ꨢ�����Z�]�U]�bu eb���V���ٸЪ���1�EF��@S�Pyz.!-ۅ�T�j�Ne[���U��Ucd��յ՞.��_�o���;�;�[@T��%����v�5�����T���*4uJ���4� I�2,O+U*��Z��ۣn�6�W�y�p�v٥]�e�U���f�g�r�	�Lqn�֫��Q�6��ۖ6{-�h���W 5V�p\>؛������0�:#v+�3�m�x��Y�ڥ.�����]շsU-�v��ʷV�VВ���b��7�����$�u������(��>	�T	V�rY�p���^�j��eUA�P�3��7*��+���HM`N���?*�:S.���CY\usWR��g�yi���/.�6;U�U
����U�OӲ�O�L�'+�8���ڸ
��e.Z�5mO;L�U��L��8���q�*�@�X�����m��U+��VXb�j�ڪ����J��*���mj/\�v&��n,����UT6+特N�l��RGTn�g���� �vtWl�
�j�ЫUFu�v�V�]n��'�����U[u*��z��v[�Q��8{A�N����&�	R�6�9b���㞺�9�:ꭩYܨ"Ѭ�n��
�jFݷUU�`1\7�	��b���J�R�q��=@��j���Z��l�(mO�9ݻ�[�:���U�����*���n:�\r�ꗎuR��꫕j�UM�]f�a�ѥ&V��ST:
��jX��bwK�n�U��n\j]C2乜��pҒʵ��7c� 3NM\R����}����X0#Su�8D9�
s&8�Z��%K��-�Vў�^�U��]����F��&ئ�;<�ִ��m���,&�q�dU8��'��0՛����6�ֻ�r���#څ4�L�-�m�����I�v�1��rc����n=�*v見��C*������u�ѐaT��t�v�,�J�7S���.	s�૶�
��k�������ލ=d�lB�@�]��mu��l^2m&�a7d`�`�lm�h�X���ӸE�j���`!�Z���-�G��-֓S�|;e�@ݎ���*�֗�"���*��N��;'7-n5c
�T�y�[r6�W���l�� ,\l��l�n�[���LA�� *�V�݀�%J�8��iv���m� f��Y��U��h�&�����V�m<�ګ�y'd)j�m��27mT��+��-�g����1T;��7^������[���UAKC��d�n����n�Uu�vm5V�J� U[UU�j�j��j݇�f�
G5]WR�UJ��+��F��\�8���sM[]U[*@�͵\�(�*��������UUU���*\E�;m<�D<�&m��~��"��T�@�6���
�~O����
��`�`����iG�;�,H)�CF�J�8���Ҡ���D9��E�A=Q=M �Qp�G��Sa t�\ )"b�p<F����$�������8�XCj �Q����O�@���S�+� �>�`#��"|�����)� �����Q"�q~�S��� T~�����>�� �*$أ��.ߏAx�/��"�).�h+����b��<<h.�hx"ES������ '���=PN ��@�R$�1E DS���(>�D<E|G��� |��
��xf����HBBc�$I�	 I I	,� �"� 2I�$`II!&�
�=��/�⊀i�u�-��dB�!m-(ZE$�) H�"JR�ƩbA�$�	DS]
<�B �$}><��TR�H���$`��R�6�Km+�IJ��㤀"�A�$�k������	UT8+�ApkD>�����
�����a`j�
�@��E����!Q�Xc�ݷ�{��/��]/0�i���\����;Wg����=c�6Ç�㝗�u��j4��a%�v����Emҕх��`%LgAɴ�1�5����sw]�0agu8��۲"l�^dwDSݶ��a�T;n�qu�t���݃���Sƪb��S/�^|F]��ۑ��\��vS�mb�l:��,�l���msV;#�-�G��wg��Γ��K����ٰ��q�R��UEж*7\��nB�z9pl�w.�kS
����s�eqn\������d�'`8	�t�؞�6����P�:"�kv\;��t��D�A]��O\�y���Gls9�!(,muItɢ��U&r�����$Ɬl�p�hㄨ�!I�3�5nc,�(��Q�Z�-a
\�ƴY��+2[Y���X��Ep�=ewg�[ڂ1��ӎ7pn�䨞{A�;e�vq�:ͺ�b�vQS�n;%5�LT�8X�Lho3F��k�%�Q�6�2Ҵ\Ս�uA�Sb�F�Q6��@Ҹ��s��Tk.�saݵ�RZx���xmlt�֎�Y:Ù�&�l��6�2gN��i�ډW.6P��\R6vٌ�S�`b����CY-ŕ.��2�c2��1�{	 j[�E�#�99���"k{k]��`�B�
 U4�f8�-mUJD��q���H	�톬Oq��>�R�n��t5u.D�WB�8��]�cv[6a�aƏsn����񛸎T�=�v &N�9ˀQ$�îX8�y|W���1m����,�֎5i�8��^��ݥD{Ai���<\q۳��:[�4����v+.���w��@+0���l%34˩̰�:�ٓ���t��N�v3���\��׵);�U)� ���e�:�Y���O&�����ٴ��U�#�CŘ��ѣ�Wl��j�pQ��6ك��\����6�[m8�長���=vٺB�2N��ڦ�|q���n�*�]����Цm��p�hr�v*�M�Xm���Ի;�y'��� �q�pCb �Q�.�O�qD>G�S�SN
�D�$眇'9=���7�5�f ��v���l�I���b ɘ\�Z�ySA� ͖��;S����JrM�I�<��.��ہ��m��@Y�Wcc8窥���c�t���.x	%�k��5�W��M�$�d�E�u�8m�f�����Y�WN�7a�S'u\{aܹ93ԛ���y���;&\�wN�n��͞L���=3v�|n�N�K��[.f����D4�6ks	���9=���q��s��ݰ��r�^{*��|�һ���&�3f̬ ��7o�����5I��	��B60wM�n۬�d���${��,T��I2�MC�hnݤ�uj��w�Ir,�v^$�X�x�����]]�n���ջ/ �L��d�K�`+�X��J��wi�n�	$��8�K�$�� �ݗ�z��z��[-4�C��٭�h�!7mt�a��۴u����u�Y��v�EЭ��?��n�T�� ��,�v^��+ ��R�!����mݻ�>�����>B�(BK, Hra�1=E6�%�\�3rNy��7$�엀rF�+`�t�2�ݶ��ݗ�od��8�%��� ݽ����N�v�
���e`]����uwe�vJH��N�m���/ �Wv^�&Vꯪz�
��2�V��m�.f�JMW)���S��A��{6��6�3-�2���Rh�\��?�o����/ ݓ+ �엀vk� 6��.��ucl�:�%��e`]������� ��J��<��)ں�Z�nI�����<�}�nx*Q��b'�Z� �7�}��7$�we�j6�B��ֆ�`]��$�d�s�%�r+Ē[�r�Ē��Y}K)S\l�3t ~�޽�����lI%�'+�I-[2�I*�ңU�wiU��kq��\�^i=�W�����T��<�Yx��t�vF��4�ao}�~7��In���KV̫Ē]�!�$��4�u�v�����=���I9&؊{*�$���˜I.��^$�]�*c�6[-�۶s�%�fU�I-�b������}� =�޾���Y�*��i�V[V��$�Ǳs�%�r+Ē[7$�-�HE��Db�b�*0Bi'9����� {�S_b,\�¶�8�]W"�I%�r�Ijٕx�Kc�}���z�Vf�6�V�pXmy��b˭EEd�z5�8�Ց�-�l��]�V�LI���Il܇8�Z�e^$���/}U��KU���$��"R��^������9Ēճ*�$�Ǳs�%�r+Ē[7!�$�v��aBn�bۻ�W�$�=��I.��^%뻛���$�S�W�����R��h휝�Ӝ䜗���x�Jo��8�Z�e^$��{8�<�>��L�L���������W�$���$�Tp�I%�Uw���o&�p�Qj���r��u�5֗�}M�3�2q�r�
϶p/ײ&ഞ@7tcSu���ϧ��v��Rb�	f���.!��=�<댻=�gx{t�e..��7�ɐˢwnxt�G"Ď%�۫��-�F.b4�`;�;&��i�G)� P��rq�4�u�у����
�;�s����%��r�8��h��ns�v���S��9$�cKNӼ���ҋl+ss���1&��!��z��j�v�m�Cvm��I��ab�ɘ9��-����ڼI%��.q$����I-��s�%�g���[V��� �|���s�mkW��ĒS}�9Ēճ*�$�dʲSV���n�m�q$����I-��s�%�fU�I.Ǳs�$)�vR����Ze�K�s}��IE=�x�K��\���ۺ =��j��s��s{�$�lʼI%��.q$����I-��s�I��>������ʛ]Iu&㖘�.��L��aa�m��zMi�@sqv�'�.P5eٛ�ϟ~;����K{2������IE=�x�Jzb�6�I����9;����~��''��p�!@��	+�,����*: �J)k%YcSF���$�Z��q@�"�m���'9m�_��7m�ϵ�}�y���^i��A#i�t y��s�%�fU�I.Ǳs�%�r+ĒK���R#�W72�S��������~�n�Io���K��W�$��E�$��I���Fa�L����:����{�$��ȹĒճ*�$��Ҕq]��rD9ӗ+����q��GM�5I��Ŗ���@������j���Z�-��ȯIo\��I-[2�IvnC�I!MH��wH��W�$��E�$���W�$�7!�$�UȯIK�[E����e�ݳ�B[{2�I%ٹqf|"� �!1@���s3>�� ���o}�~��=kPلu6]�1$�f�9Ē�ܗx�K{2�Im��z <���9�c�����?m�x�K{2�Im��1$�f�9Ē��Գ��d�˖�ny.�M���p����P�E]4��L��i6�7,�m���[ِ�$��̳��܇8�]W�� ?y��R%[AeW7��<6e^{꯮�-���Ij�y^$��̇8��z	}�4e�rfn���׷��K��W�$��!�$���W�$�,�˲��Ֆ��$�UȯIofC���o�l��tE(��\�}����%"@]�����;j�I-��s�%꯾�����g�q	v�K�I���t����s]�¦�ƂL�.�Vfm�\ ;�@e�1jl�;h���7[�p+v�q$��e��K�r��ܗx�G�����`���u2:桲����܆q$��Ex�K{2�ճ*�$�=���у,y��ao}�?�M���q$��e��K��\�In���Wt��a�Pɺ <��^޻ ��ަ�v=��I.���I.�%$�M���t���$��̳Iv=��I.��w�+}���9�m��VhՆ��L,C����u���Xa������Y�(���l� Ta,�`ێN�\dY�=�� ���qX6��K:�cō���Ė�������ݳ��zz��Vq�C֗NX�s�v�nG]Dv�����e���b�ɟ%C{u\�W�֙�q��e���5��z�;ln��01����k��%�95yf�xD.��sh�|��Ӝ�w�Λ˔2�[���xt����vEOS`�տ[����"RѩM��4e�rg^�������r]�I-��s�%��,Đ�d� 4��vR�ue�s�%�r+�$��!�$��̳IvnC�I$��E+�T��@���$��̆q#ofVٮ6�X[Kh-%r��hB�l�;�2��p�9�"�7�� �`��ջwv��v�۬�\0mȰ�p�;�2�ϰ��wkq�H���b���6U;�5��P�\�J>3��u=	�N�g�:��m;��ـsve`��sve>������ �G� ݞ�t��&�wu`��$�ϵ��O
�|@� }����=��,�0v)I:1�t:t�l�;�2��ذlp�7�� �D(��I��e�n��ذlp�7�� �ɕ�e�Pһ�Յ��k �܋ ���&Vٮ��Ͽ���C��t�eefe1�d�u/��8�C��Kl9��L�xb�ŉ�XnP̍�C���?v8`��wnE�E����W,�۱	�fݎ�H�G� �~��7��=��I�	��v�m�]������ݹ�ȫ�X:�h���a��f]��醒}�)�UҒ�@��kЏ����х0z��Y��ד�0�Ɏ��d\�o4l��ރR��İ�|�X�a	)�NHs���!�0V'�����������9�{�n\�=ߺ}�|f�x�E�([��5�y����yaHYp׌bB�^{���1�
$w�#�M�pP����J{��;Ͼ���L�C��BrE�jk.\ʱX��鿈�[p��ғ��K�Z�ui� �uě�\�*�>�B�5LI�Č�8���tw��{�{7Xa�>+��q�Nv0���]^K���6��[�K�|�Y�6Mm+���&��y�!u����u,�h��ꆐ�8� 	�H?x���"�r	Qo A�$c$$X0��h���(�E-�0@M�'ʠ}UT��_WՇd}0ݙX�.�*�B��wv�0�Ȱ�p�;�2�?rrN_?{��@��_�)��6�P�0�p�;�2��p�9�� ޛW޲h�f��$6V�f�]�<(�p�e�5k�*�
���qP�e�#�3F�f�ٕ�l��=��}����<�z��baMҲ�۬f�`ۑ`5� �ɕ�KD���0j��l�:�K�6k�ݓ+ ٮ�_�gͻ�����,�~�f���o����R��X#d,`G@hVg��, �����n���ݓ+ ��zg����j����)&��Vs��`H	'g�w%�Ɓ9.5��+�ntt{%g�\�j�K��̤�f�s:�|}0�Ȱ��`�2��&UӥN�]�[�N��:�K�6k��ٕ�l�� �u��,�v�j�v� ٮ�̬e�X%Ȱv)C�@���l�7ve`/b�9.E�l�-%(��BvSj�j�`/b�=�w��\z?�̬�����'xY�N���i4Y�j@��O�C�c�;h�8�X�u�u����v�j����#�@�7K��fu����vN^Ұ�öʽ8��q�퍚��;�A��s�����;n�O�hȜ�������:!�yvc��T����Ed�o������A[4
��g�j���;�Iavւz�ƚ�2�5�Ϝ]��㓅 ]��he��
�^:�I�s��'i�S��̭q�ql�Ǽ�f�2�����/33^��I%��Y�6$�hQ��ucmp���l�vL�e�X�]@MU�ci;k ٮ�X�ذˑ`m-��Au*�E�ݳ ݓ+ �{�r,f�`[�>eӶ��;m[�f�`�� ٮ�Xf�*�;)�ݤـvG�UU}S�<p	=�f�`+�]��ݰ���N� A�a��ɋv�p��0[n�)F��=8k\�]6՗b�%l�6k���+ ٮ�諭�������cMX��5�֦����7�(U��9�߾׆�0�ឯ���#��䆛WWtҲڷX�~0lp�6k��ٕ�KD���mڵj��l�9�� ٮwfV��,TԀWP)5v�6�m`5� ����6^ŀw��ӫo��䟼e>�B*�f�s��=Z' �vrX�X����U̼�Ry�88���huM��n��6Oe`/b�9�"�6k��ڗw>eӱ��m��X�ذmȰ��wve`uL���`��n�;k �܋ ٮ�T/Ca#��A���0	%�01����@��a�#��$+������e`�"�;����M�]Ҥm`E=3��{+ �{�n{׀E=~���V'@��ـwve`����{׀oc������{�
}�&lc�����uuڰ���<dleQ���\�z�a����~��hqӴen�����8���oc����I� �z��4��+�ue�`[%窒&���6Oe`�ឪH��"���
�m[�ջ�&���;�2��p�8�K�"�[@Z-��X��`ݙY$��u�ܓ���]��!�� �1Q�����r����!���h���wn��p�9�"�7�e`ݙX��/�e����� ��8�Kn���NSBh��J���r�z��.��J��vv�n�&��~��7�e`ݙXf�`ݙN��+�AwJ�]��od��RF��}��r,V˔�۶*t��n��̬�\0�%�~��&��XP���I:wV�fٮ���X~_������~0	��&ZU��N���w��n��9'+����r�����G� �ꢏ�>�����G��Ch2�6�STr���)����an�`���٦Eͮ�렲��
����Ka9x��;���* ��g������;s���lBl� f���Oܥ�p��G(�\c\���8���Cig�s��İq�p�4h�CLv���`���G(�K�]�9���WB���D�1	h<���&��j�Jm�Vb#�6��\��it>)�*�
���z�j����������Wݑ��tg<g���l���'����i�\��zsp2��n���w��7e����v�۾�y�0T�<p�?����{���҉@Z��g͢��ـl��z�#����=���RSc񜤎��w걉�Iղ�l�9�w�<p��^��q��`���*h�����M��/��W�uz���������]��['�N����*E�w�M����3� ��qI/ ��p���;6�k�˕�Øʚk�\u��ACq�gk���0V�LL����we�j����n��G� ���Ix�8`V�*M+�j�i�[M�f�e}�}��0)�T�"H�I`x�FLF	B�,�!$4�-M���k��,��� �ٕ���7��̶Л�WH����y`�ᇩ)'���~0SR(�"��e�N���g��$�V��U.߽��J%Y���MҴ��0ݙXw\0)%�ۑ`JJ���t�T|�$mٻ\-	M/;mPL���	3G��0���n���4��5v�ۮ���d����� �=��O{ה�����cwbl�8�K�}I����{+ �u�=�i翿v8�5`+4�s��7�ס<�߶ni�E4*"��l
(!|@]"�9{���������<�{���r�X�g-��}T�Or���,�d�}T��y`U�T�WtՉ��ڷXe�X����z�����ٕ��R�\,.a���gr�r�^���G�+���4t�sg��ܒs��æ쀶�S�oT�� ��ŀwvez������^T�n�hV�V� ��Ş��䍓�X}s� �^{���
��QV��h)�i5m`Oe`��a�����W�z�~�x��� ��.�v˲ݶ�X���]�XT�� ����ⶾ��Fb��@4
u ����v}�ݓN�VJj�3WrN_~�7$�����~]{߲�Kذ	**&1S�f��nykl*�������<����=;;\a1պ^�lG�9$�ؤq����7;��s� ����/UW����x'��"��1�gd����_o_I������{׀oob�UU}IU�y*Wt;I��ݶ`��,�d�=�W�IM��l��rG��wl.�&��Cmd��O�k��f��;��I�k�?ʫ�Z�3 2	�ۢ��i5�'�g�]�?(���s��I����'����Ӈ�n�@��M{�@�&o�6�(FA!%!��q'ku������ �ĉ2,�&!��*HJƄB! D��B$��̓Hr!H��mm-��o��RVl��#%%�ff��.$��Rx2�l͚�kg4�sW�3z�kA���כI���!�B1B$�����|֎p!8�nP�p ����#)*A�`A�%�ܫ=�C������0vI�aKe!�1�q�#	O[���.h#���H����Fb���҃!Ĥ(��c�8�0/��f�0����
d��y$bI�{�q�0sE�VKI[X�Ki	5/$a�$a$� {�fy�<sG9v��l�vCf�6
k�T3y/�d�#@���I $�D��3��Pէ��!�1D���H"�0�����D�$�0��$d�BH��$B`�9�l[�)#$I";�����}�����C���+<�d����R�����{�5c�L�13EY�g�
�)�d���k�v+��}}���jbz���2�7�1��5Hnܛ�X�"�V�k��&{QF�x�S<:�pf6�jƪ�B٪)�.��c	tq�t�ƥQQq��x:��s�;%�ڌ��m�ț6���v�*�ô�(J�������U�.Z��;e�{/y�zr�E"�t�=�[u�0-�8{YE.`�c8D�@\봮��:���,�+�dpv��X���"�I�7s��]͠�Pmh�<��m�F]�s�i,ۡ���X��v`@k��p�˝�4Vx7#m�ٙ����c�0�$��ғ�ݲ�Gi��h{<ּ����v⸀��;7;�*�]R1�.��6�yf& Ŷj��Ʉ;3"�bh��7m�S��影险��n��A�P9��]p8�(��N�n=��p�Lt-��`(���m�S[k�ް����d�pwl[3M��p�(�+1%k,.��+!����������-3�A�ʴ��A	�m�6s�`��< ��U���*���l�:3V���i�m��3qbh�;��J�5��z.��z�]�1������"���&rN칰a	a��&6��ȼڧ*P��Q�7XQ�l���+5φ9x�F�!siڜ���4�!5KLe���Z��H�U�C8^Lu¹dۥ����)���3V�v�/M�gj�u��kj��M(��6`g[��m�dÍ,Ag��zgd�ٻqS�bd`ż�Ƌ�^g�A�(ָCY��u��� N��=���spf�KG ��ݤ:��I�n���'b�r�A������(f#��7�<Lb�H��C.��e'(�x ����7	`9�p����k6 '`��qP�Y]n��T�(��b�����֡����]�:��=�qp�$]+Wn��12d���ݥh;K`1�����f�b��ӧG�����������Q�-وB��m�P:�겖6W��v�b�Y�`U�*ۦ�n�r���'>�$"�@�*��:*s�_�W�Qh)ꊀx(���C[3�MK��������kZ�0���[�Ot�grۢ���8'3DbK��i�ohIM��e�/0qWc
�[s�M]'X��Y��^F`���S�r�8uMzB8;<sȹork`�&��4�x�5�$׎��`m"��;`8�+d�2ʄ(�.jF�(�a�6�Wl�9�Nכ\�<G�4��q��cl#ĺ�E6�-G[t�h��ض5��__���rr������Y(q�7M�^����ѓ	u����ã��sFb�ٮv����"��0v��u�V�����t�ذ�%�����	��,-�_�B�A���-�����_Ns�	����iȖ%�b}�۴�Kı>����r"�%�b}���)4�Yl��[njm9ı,Os��m9ı,O��{v��c�*dL������Kı>����ND�,K���5�k&]3Y���fk6��bXX�{��m9ı,O���6��bX�'��}�ND�,,Os��m9ı,K�ݽ-�ֵn��0�kZ�ND�,K﻾ͧ"X�%����}�ND�,K��{�ND�,K�{�ͧ"X�%��~�5L�b4ʒ���`�Rʰ�@ؤ-f�S) ��������現����Zy�Z�ND�,K���ͧ"X�%��w�ͧ"X�%����f��"dK��o��r%�bX�~��?�.��5u�,�jm9ı,Os��m9�B�+$Q)	Ya�M�X�@�`B-� �H��E$Mı5�wٴ�Kı>����r%�bX����m9ı>���Ҩe�YL�듻�^B���>���r%�bX�}���9�ı=����r%�bX��k��ND�,K���7�jGZ.N�|9)�I$�8}��۴�Kı=����r%�bX��k��ND�,ʄ r'~���i��^B����?��i��՛eru��Kı=����r%�bX�����9ı,O���6��bX�'�k��rwy�^B�~�_��;�$[2�R�ts��M�kcA;R(��d�{!�����'��rH�tJ�pR& �듻�^B�;��{v��bX�'�w}�ND�,K��݇�('�2%�b}�w��>��%9<����3�y\���oxr%�bX�}��m9Fı,O��{v��bX�'�k�ݧ"X�%�߻���r�bX�%��ޖ�,��֡�ֵ���Kı=�]��r%�bX��_v�9ơ�(P@�PdK���fӑ,K����iȖ%�b_��e:[3Mjk�f���bY�b�dO�o��ӑ,K�����ӑ,K����iȖ%���c<��N�$���{������0��	 �'��~�n	"�{���m;ı,O~�y��Kı=���r%�o!y>�6�{%�65��C��5e��]��u����(��x��x+::��������+�s5�˖[u���Kı>����r%�bX����iȖ%�b{�}۱ �Kı;��{v��bX�%;�>a0��զ��WZ�ND�,K��m9ı,O{��v��bX�'~��siȖ%�b}�۴�ĳ���>�⚊�D�g�N�!y�^�_v�9ı,N���siȖ�b}�۴�Kı=���ӑ,K�����Ri�4�W-���ND�,�C"~��g��r%�bX��_�]�"X�%����6��bX?�@Q�] �BD��~��9ı,O���L���W#-���'Ò���'���ݧ"X�%��`�}���v�D�,K�����Kı;���ͧ"Y�^B�{=��1M��l��$���]�oB���>1�Q����M!o�������#�pe��gd듻�^B���_�:ND�,K���ݧ"X�%�ߵ��6 "X�%�����iȖ%�b_o���cRe�g)�'w����/'���ݧ!� "�L�b~�~�m9ı,N����ND�,Kϵ�ݧ ��^B�}��p�:�Vj�2�N�;�,K����u�ND�,K�u�nӑ, ���w�iȖ%�by�}۾N�!y�^O7�l_�!��Q˶��bX'�뽻ND�,Kϵ�ݧ"X�%��u�nӑ,K K�k��m9ı,K��~a3��5�l�֮ӑ,K���w�iȖ%�a� }�}�v�D�,K�u���iȖ%�b}�۴�Kı<�7w)��<��cs�#�7x�Ҙ�TYƔq�Iq��k5��k�����l��mpk�h�.��R����y��b�8�ݰ�6+Q��p��$�ݙ|9�M��[Ζj]L�q�.���n��2�[�:٤hs�Z��Gt��x��l��\M�Wc&�v!��:�y�M�a%�S(�@44�^���;;ou�D�.�]���<���I$�9�K^�˥��^�n�j�t�n'kn�I��b�8�p�;c7nv�7��8m/M�m.sFm���'Ò��%������r%�bX��]�iȖ%�b}�۱C�,K���w�iȖ%�b}���)4氖k.e�56��bX�'~�{��r%�bX�{���9ı,O>�{v��bX�'��}�N@��������vԎ�<� *u�Ȗ%�b}���r%�bX�}���9�Bı<����r%�bX��]�\��B�����|}0�Ͷ[�WSiȖ%�����nӑ,K���o�iȖ%�bw�w�ͧ"X�"؟{���9ı,K���N�r�n]jS5���r%�bX����m9ı,?��E�w���i�Kı>�]�v��bX�'�k��ND�,K��,�ۋ�+���Q.��:���#�T�(������7�^y�A�\X��s��\:�s-S2�Z�O"X�%�����Y��Kı=�_v�9ı,O>�{vȖ%�b~�rwy�^B�y�����S,�rf�Zͧ"X�%����i�hZ��\�bX�}���9ı,O}��6��bX�'~�{��r'�D��"[���(aD�P��'w����"w?~��ND�,K���ͧ"X�X�'�k��m9ı,O��}�ND�-�/'��>�!��(�m��;����<����r%�bX�}��Y��Kı>����r%�`�X�g{��wy�^B�{����+��&\�3z��Kı<�]�iȖ%�b}����Kı>�����Kı<����;���/!y'�]/εҙ�����ʴ�F�j�ls:����N'�����j������r��3
���u���/!xX�{�xm9ı,O���m9ı,O;��6���bX�'�k��m9�B���m�u�ȳ�N�!Rı>�����Rı,O;��6��bX�'�k��m9ı,O���6��$��y�^C���>��P��&�ͧ"X�%��~�fӑ,K���w�ͧ"X��HE"EIGJ�UЀ��b}����Kı>����r%�bX�w]�t�[&h�Z�ԓ5���K�lO>�{��r%�bX�{�xm9ı,O���m9ıA[���ͧ"X�%��w���L��\��rwy�^B�{����KİDO���m9ı,O;��6��bX�'�k��m9ı���S��#�PZ���M��r�e���۝6j8���wCW*����0b�����$�֍�"X�%��w�ͧ"X�%��~�fӑ,K���w�̀Ȗ%�b}����Kı<�K�wS&f��tK��5�ND�,K���ͧ  ؖ%����uv��bX�'���ND�,K��{�ND��D@ș��_��d��ڙ��f����/!y,O{��v��bX�'���6��`�bX�g{��r%�bX����m9�/!y?y�_h#4�+��S�N�!R�F�����ӑ,K��;��ӑ,K���o�iȖ%��< HE~M�����5v��bX�%�������0��e�듻�^B�����fӑ,K���o�iȖ%�by�w�]�"X�%�����"X�%��Y���	g��I��xL��⌭O<*�g�#�`�Xv�歛yu��>o�w�����p$j᫙��yı,O�w�ӑ,K���ﺻND�,K�{�9ı,O���m9ı,O{��;����5��Y3Z�ND�,Kϻ���9ı>����Kı>�����Kı=����r'�V�L�bw}��R;E��
�rwy�^B��߿p�r%�bX�g{��r%��%��~�fӑ,K���w�ͧ"X�!y�{���F�2WZ+:���������nӑ,K�����iȖ%�by���fӑ,K�����ӑ,e9)��y/���l��cf����D�,O{��v��bX� �k��m9ı,O��xm9ı,O����9ı,LGD ���{n�L�,˓F��C��m�#�W��uX�k5��L�`�+*A���[����n����ؾ��J�JV`���"VY�0�i=k3���e�����jZ.�9x;��^�M��(B�\vn'���v�s�n�����.�8*�
����Z1�z��i7V�iTh���N��byy8�۝��4u��F:ˌl.�hzz�������^���*ߤ����z��:7`���$e�S`]�����ۥn-vG�B�����*�f��ܓ����G -P�:������������ND�,K���"X�%��u�݂��bX�'��{v��bX�'�����f	�J]�'w����/'�}�NEı,O����9ı,O;���9ı,O>�{��r%�bS�����j�("���JrS�����nӑ,K���nӑ,@[���w�ͧ"X�%���w�ӑ,ay�{|=�`�@�&��������X�w��m9ı,O>�{��r%�bX�{�xm9İ?�ȝ��߳iȖ%�b{�_����̺̦�f���M�"X�%����u�ND�,K�߻�iȖ%�b}��siȖ%�by߷ٴ�Kı/�vL��:@S�������D�L��vؽ��BDVz�؍�v]q9ݦ�:�R�
���c5O�9ı,O���6��bX�'��{v��bX�'��}�PD�Kı<������%9)�~��B~AڍK�Ѵ�Kı=�۴�9�)����"%!���7K&��SL�Q؆�A4U%pԬ�$5AlL"�	 /��= $K����ӑ,K�����fӑ,K��߻�i��X�%��|^̝e։5���35v��bX�'��}�ND�,Kϵ�u�ND��� DU ș�~��iȖ%�b}�_�]�wy�^B�{����#��-���r%�bX�}����r%�bX�{���r%�bX��]��r%�`�X����m9ı,O=���jh֍[���-�kY��Kı>����r%�bX� ��w�iȖ%�b{�}۴�Kı<�]�iȖ%�by�4}/rF+ô�i�iݏnp�`���|�R���;;F�8�#D��d��'��5��L�����ND�,K�뽻ND�,K���ݧ"X�%����u�A �Kı>����r%�bX����ܶ��\���k35v��bX�'��}�ND�,Kϵ��6��bX�'��}�ND�,K�뽻ND� Ar&D�/�����]v�١��'Ò���'����6��bX�'��}�ND��sG��~P� �`�$�I!�yy���$�f�ć
�J	�B�@�A�
,RD�XFI#N�$�c�E��@�O��a
[B[bZ��Co�y�4�%���
��k�]rR������Z�Gjf���P&���o� 1���0a$�&s�b��!NÄ9!8xLXP~.����;<�C�H�BKne) �`���r�0�̈́'9�brD�f������,
�l����#�xx�{nr��-�2Y���7���F� c�a��D��=��}b@d$,h��FB,,��4�l���$.ffc�k��t%�H�lf%cJa�j�Q�Dt*=(	�h���|�B�*��v�� 5��A*l\Q��"X��\��9ı,O=�}�ND�,K��块Z&�s5��Y��k6��bX�%����fӑ,K����nӑ,K���o�iȖ%�by���fӑ,Kħ����u�e�\�e���r%�bX�w]��r%�bX�����m9ı,O>�{��r%�bX�{��v��bX�'}�KI��hV���%��au�V��B۔�Yc
�3\�	��v�L��7��I;YSv�9�kr��]�"X�%��~�fӑ,K���w�ͧ"X�%�����a�D(�DȖ%������9ı,N�_��p�fĹ7�N�!y�^O�k��m9ı,O��ݻND�,K�뽻ND�,K���ͧ"�ؖ!y?y�_a#6���%.듻�^B������iȖ%�b}�w�iȖ?�"��L������r%�bX��_�k7���/!y�}���l�ź.SiȖ%��X�w]��r%�bX����m9ı,O>�{��r%�`T:)H�"�QO2����nӑ��/!y���XEDc�N�;�bX�'��}�ND�,K��w�ͧ"X�%����nӑ,K����nӑ,K���}��$��5���0f�K���B.�7�-�±y��
�fm�t eI�|����z]�]mԕ�N�}9)�D�=�~�m9ı,O��{v��bX�'��{v
�bX�'��}�ND�����>��_�b7h�%�]�'w��bX�{���9ı,O����9ı,O{��6��bX�'�k��m9ı/����u�sW.Yn�v��bX�'��{v��bX�'��}�ND�A�,O>�{��r%�bX�}�����rS���������G#�.��]�"X� ���o�iȖ%�by���iȖ%�by����r%�bX��]��r%�bX�����5�DպԷ56��bX�'}���iȖ%�a�������i�Kı?~���iȖ%�b}����r%�bX��Ou'����L@@"�ZP�6!k��,w3�J���9��CIk���+*KcM^:ck���YdF�S���*c��o[�ɗ':.{kdK��m�Λ7���¸��gR5M%�5ۢ��v��)�NMn��T�<�۷P�6�p(��,�&5G[g�(�ܐ;tPX����S�u̽��K�]0>^�yP64b�=�^��6 ��k5ٚ4%��+4̱�K*��o$�$����+�5��mX�;Oc\��
\s��ݡ�nmۇ�X�k���=\�͗Bh���:�Ȗ%�b}�����r%�bX��۴�Kı>���m9ı,N���.�;���/!y~���͕��L�ND�,K��{v��6%�b}����r%�bX����]�"X�%��u��\��9!y�^C�������Z��fj�9ı,O��}�ND�,K��}˴�KlK���ݧ"X�%��뽻ND�,K��'s�fYrK5��5�M�"X�%��u��m9ı,O;��v��bX�'{���9İ��߷ٴ�Kı/}�Y�u�K�u�2�Z�fӑ,K��o�iȖ%�`�{���9ı,O��}�ND�,K����r%�bX��d{�M{BR���c��A�b����	l� er�Fi�lӻh�x;sXA!�{�"X�%��뽻ND�,K��fӑ,K���r�C�,K���n�;���/!y?o!���p��,vM�"X�%���o�i�P<' "���v��@�,K}�����Kı>�_v�9ı,N�]��'w����/'�_~��3GV��/IȖ%�by�w�]�"X�%�����iȖ ؖ'���6��bX�'�}�m9ı,O;��.���f�)���֮ӑ,K B��ﻤ�A>��sbH$��}�I�$�����uv��/!y�}���1�S`�.��'u,K��;��ӑ,K��w�ND�,Kϻ���9ı,O��ݻNNB������ݦ�X��yX���
���[l["�Y[)���"�S��gB8�:�-7�s���l�2���;��NJrS���߿|�r%�bX�}��WiȖ%�bw߻�h�bX�'���6��bX�%��߷��iQbg�N�!y�^O~~��ND�,K���ND�,K��{�ND�,K���m9,KĽ��_�Q��5Vrwy�^B�}����Kı>�����K� +�C�E_@^)�dK�����Kı<�_~.ӑ,Kľ{�)Ι0�e��n��iȖ%�bw;��ӑ,K���}۴�Kı;�w��r%�`���~�fӑ,Kľz�~ƨ������'Ò���'�k�ݧ"X�%����9ı,O;��6��bX�'s��m9ı,g�%��㹕���r�a�R�K����[X�G`,^��h�fs+e�����a��I���r%�bX����9ı,O;��6��bX�'s��6!Ȗ%�b}���r%�bX�w����k.��Bf�]�"X�%���fӑFı,N���m9ı,O}�{v��bX�'��z]�"X�%��w���3Z�k&[0��jm9ı,O���6��bX�'�뽻ND��,O{���ND�,K�{�ͧ"X�%�~���6���!��'w�����!y<���iȖ%�b{�w��r%�bX����m9İ=�"�j's{�m9�B����߾Si�B�c�u���"X�'��z]�"X�%����}�ND�,K���ͧ"X�%���nӇ%9)�NO���=����e3)5������3Ţ��]��������/-gf:����-��U��%§\��B����y��6��bX�'��{�ND�,K�u�݇�By"X�'�~��]�"X�2���B�m�5���w���NJ%��}��Ӑ��S"dK����r%�bX����v��bX�'��}�ND��D��,K��~�?d˓F�L˙��r%�bX�}�߮ӑ,K���ﺻND�,K�{�ͧ"X�%��}��ӑ,K�����)�f�kWVk5v��bX�by�w�]�"X�%���fӑ,K��>�siȖ%��*�O����iȖ%�b{�]�uCY�Ma�ۚ��r<�DȖ'��}�ND�,K����w�m<�bX�'�k���Kı<���ӑ,K����!�b`!(��X�w�vf3r��^������ͻf�9�s��A
8̷Ya�(�f%��Q͍�x��a7�^�b�v�����`�xj靋�+�r���1�x-�ݝ	e��q���`�.�
1%`N��^��1$ٙg۝�-�1XL�]���l��vMC's��d�(�[�L���4���ٽd�tu�8��]�`К�e�`�+	�2�Tv�w^���{���C��8�Yw�Fn��HM��<<[a�$�M�9��f\ڻ7a�w�9;׽��#
�i�ʝ��rS��������6��bX�'�뽻ND�,K�{���9ı,O}��6��bX�%�����*1�4C;�N�!y�^O=�{v���%�by߷�]�"X�%���fӑ,K��}��ӑ �,ay>�����pXZ�;'\��B����o��ND�,K�{�ͧ"X�%����ͧ"X�%���nӑ,K^C�=����j[�:���������"X�%����ͧ"X�%���nӑ,K� �C"{������Kı/�t�I��K�ц��ִm9ı,N���m9ı,N���v��bX�'��}��r%�bX�����r%�bX��|[������/W�����&	R|a��g��rA��;gF��>���+�㟝�u`2?{�7��bX��_v�9ı,O;�����Kı;����~QF"�"X�'���ٴ�Kı:~��𦋚��j��f�ӑ,K��o��NCA(8��"X�'}�}�ND�,K��{�ND�,K���ݧ �bX�'�}�ė"i�S)�'w����/'�k��ND�,K��{�ND�����?w]�v��bX�'���ڻND�,ay>��MT���b���'w���,N���m9ı,N���v��bX�'��}��r%�bbw�w�i������李�V��n�.듻�ı,N���v��bX����߼��yı,O�k���Kı>�����Kı/���~��.�\5���]j��˚�a��m�I�u�Vcځ���n��rp��N��.������|9)�NKϻ�jm9ı,O;���9ı,O���m9ı,O��ݻND�,B�xz�"[�L%��N�!y
�'��{v���bX�g��m9ı,O��ݻND�,K�{�jm9K�^B�~��Igݮ3����'\��%�b}�w���Kı>�_v�9�b���F�$ B@�$d`�
D0�H@�1
1ljA� @O�q@�"r'y����r%�bX����]�"X�%�{�>��)�s ��'\��B�s�/'޾�v��bX�'}����r%�bX��]��r%�bX�{���9ı,O����%r�Q+��N�!y�^O�����9ı,;�۴�Kı<�]��r%�bX��_v�9ı,C��K��6��1xm0ejFÒN�LkE��wB[n�A1.�W*�CF��p��S g.�0�]f����Kı>�]��r%�bX�{���9ı,O{��v��bX�'~���m9ı,K���L��\��%�f����r%�bX�{��m9�1Qș������9ı,O��k6��bX�'���ͧ"X�%�}<�+�GP�&o\��B����y��v��bX�'~�{��r%��(Dȟ���M�"X�%��o��r%�o!y>����!���;'\��B�T,N���Y��Kı;����r%�bX�}��m9İ<�H ŀ�A�j��N�_v�9ı,K�ǡ1�]�D�(��rwy�^B��o�iȖ%�a�
'����i�Kı?}���ND�,K�k��m9^B���/��}6�+�f@��;C9�r��溗e��-���"���wY�i�Z�j��Lִm9ı,O����9ı,N���v��bX�'�k��lyı,N���6��bX�'s���ɪ5�'y>��%9?x���9 Rı,O>�{��r%�bX����m9ı,O���m9�2r������Һ9���'w���K����]�"X�%��~�fӑ,����fӑ,K����iȖ��������B�g"8�*u���,K���ͧ"X�%��{�ͧ"X�%��u�nӑ,KlO>������/!y�y��Bk�Lf 1vN�9ı,O���m9ı,N���v��bX�'�w}��r%�bX��]��r%�bX�.�����T� �\a��)L��I�.$c!���J��+P�ݏ�20�`�B8r�6�v����p�M�e(H��HA �(@��A�1�$�i�"H�)aI!$��<�����CQ��p�	��y����*��d��!6D!!L��i| �H� �$#�ń$�HINo�Nl������l-aiHa	�c�9j�	B��@! �B��9rg�M�rI8���+i/�Y�B����f���k��Rfw����&Nb�\�n\kN���GĥpJ���;z��.����Z��3@�H��<"�ك�3��2d�!ZYve(�pMA�8cy6<.�Z�i�*B6�C���u	���;u� �mke�SbC$3`*QM�u�p�uO>���<���`Pyö	yNz{sۜ��Uc{pVc�C��[Iκ��Nx�R�c����_,ɘ�-ˊ]la�����X�BFi���j�ҍc�-jl���� �j�.�jwh9�Gu�<��y��3�w6ţI����ҐGi�Q5]��H�k-V�,B�a���eR�a �\X��O4�o'��ek�F��3j�V�f��a68����S�����&{0pM�Ӗ�G'h�p��؅���4�U�v�;Y�MT�+�-�,H�����枚4�s�&�;z�5���vԙ	;)g<���e�0���@���I�=��85�sY�렀{�m��҆a'x�(�^�ŷ'a�ٴ㕐��mke]���`�nG[�cvɃ�IY�X��ۖ����ViӍ��pT��rn��ev�V�ˀ��ۑۜ�q��'���q�q�v����3���{8uu�j��j�(d���,�
Ƨc����k����l����t�Q�5s�=���v$�V���*�vf�� P�P�a�� �0�[�SLv�΍N��u����V�e¥�7n���d�M[s��k�Q`Mv�Ԇ��@f��Bv7D�9�,+�@��$�8�Σc���u\i��3�ny-�c!����FQc�H��]��g����1ͤ�ݎ0��:nZp0�7-�Ņb�¶)\�;&:�iSvt`�[��Ds�'N:�=��<�g���qhZ�n<�X�h�XD-��*GWd��#�륦�e!�0%�

;�̩�'�X���H�����3�x7d��p�%����p�,;s^āDv�(�¡���֣�]�jU� Lq��)Ř;tp���/&rch-�9,n¥vfSA��ֳ5sfh�Ѯ ��(W�~P��T�� �����}PH@P�����u�rw��i����dc`�*T���[*��	fD�;l]&��݉ r��֐.v��g A�Nv��\���Q��wF�]!d����	��A�S%T��g8/,v�N����<{j)���19�l)۲�b}�b�n��Sss�0��#շ� �=,J�v�u��+���7E����.��[S6�\���nG5�[u�8�/[�zE/j��'~{����,%�˜8M3�����Z�;`���\կY�[t»��K�C����]马��r%�bX�}���9ı,O>�����Kı;�۰�"dK�����6��bX�'��~���f�j��Rk4k5���Kı<���ӑ,K����nӑ,K����fӑ,K����nӑ? �șĿ��������
,�[gZ�D]u2�ND�,K��}�ND�,K�k��ND�,Kϻ���9ı,O���Bw&[�5�L����K�,O���m9ı,N����9ı,O>�����Kı;��۴�Kı;����� f���'w����/'~�{v��bX�'��}��r%�bX��]��r%�bX�}���9ı,e���}���]�da�M��%�oGv\��笱��-�٬�.�t\�s�xn#F�ֵv��bX�'����l9d�����=/�_������w�~���+��l�B��6�,_W�U���ꪦ
\� �r,�8� rIJ�Vʷm$���f%Ȱ	ۑ`�#�n�`���4%t�uh�n�v�X%�� ��K�`�Q\e�MRl�v�ݵ�r\��Mp�$���� 9��e����6}<�pD�7E�i@��.��k�$�3���k[�)�఑�ۼ�\0	.E�oob���q}~�H���Yb�k��+v�K�g�睊#�s� ��w�N�ŀuv�� 6�E��V�;{�r;�}N��>#B$A��GS��9�ܓ��ŀmM�*�wM�Lhv��w��w�{ny`\�����y�拥I��e��x��X�"�'ob�>{�����i��j.ˁ̓4�`�o&]F;"�U%]�;D�)�1[;�sW�W��I:n�K�`ob�9.Gx�ȰWV�mSt�t��X�ذK��;r,K�`�Q\e�]���N���w�N܋ ��X�ذuD�(�V�]�`�y�:�^����I��{w$����:"|�d`1��y�8�@�FFG)!��$�Iб�K��H9d��Ac ���jh�FDt�I�"RV�)
Kk0�b��|<hϫ�;�=ؒ��Yb��E�V��K�`ob�9.Gx]���� ���t+@	X$C�2�\�efU�J�� ���A���fb��mu�5B�\�7�{�ذK��d�K�`RE�t+[tSV�m`�#��I[�^�_��	��`��i+���i��ۼ.�x�"��Iz_�����x�%*�.�ݻ�I]4��%ȰMp�9.Gx��/g� =Z�טZwlt�t��X&�`�#�Wv^%ȲI��#����e�Բ�.��֢��K���祰^�Ks��]fM��u�ON�۲\q&�Ȕ�2�Xabb4�1ñ��n.���,���f@�Do4ą�rmA�۰�J;7X��읽A�&�#����lm��Jyw�s�m�������B�#��y�|l*l������w=̽�J�^�=�;#��,�%�2J�%�GM#����!9��jֺU��{���9��;�����cl��6RV�iƆ��i��a��&�Ԃ��6mQ�:�@����;g ݿy���/ ��^���;��`�y/%uv]���Am��j���"�^ɮ%��?}_U}���쟼%J��2��R��?/߿^ɮO�K�K���,���YwawWt�a�S���;�?5�N�ŀE$�jBe]ZV�դ�0H�X��� ���x�`���m۠����<̓�ð�t�SE��f	^:�9ģI�n���G4���V���=��$�{���;�?5���+�Ӳ�t��xRKľ����}�ʫ�o\0�8� rly����v��U��M[M�]4������9#�`&ǀE$��p��[��[�ݺjف��}��X�{� �Ix�`�7cj�����[m`� ������H�`�ư	�4*Y�ҧK�J�
c�`��͸�8$�h_I�z[Q{h��㵗E��|;o �Ixf�`�ƽ��� մ��̧N�Ӧ�n��៫�;�?5��� �Iy��#Q<y�իBhm]؛0���`�s?Dl"$I!D"�$�
B�l	��F�-"�`�D���#$�"T�,H���b�v���;���rG)���Llt�m��{}�y{޼n�`~���w��5��zˤ]Zv1�];�k ������g��y��v8`I�X&骴�Ӵ��Ł��apK63�3�6������g���v����;T��ݦ65t����~0	#�`���}_q}~��=��_��M����tճ �8�;0K�`u����������AS�R6� e�0Kذ��I��s�*N�E'v�R���7���$ٽM��"��`0�"�"�� �_�����{}/�'�jh[;�ـl�����~���=�>���{o�veJ��9�#lT%���UT�6�1��L0 �:�l�����Z���զ�M�� ٱ�����	��`�~���L��nЄ�0{#�95� ��M����Ԑl���E��MZ����;��`��I��j엀���S���t��`��I��j엁諭���L�{o¿]�l@���bl�$ٌ�=_}T��� ��lٕ�O���(���� B"1��S����! $+"�T�,E��ۖe3���7Z�.��t�,q����9�f��a�9����ռ�[�wX�E�)v�[q2vM�B/;���D��'�y�-ۤ�	苠Wq#m�78�{����6��ݴ�N]�Q��x���5�411��!jw;��i�D(�,7�+3.��f��h\��\h���W��,6���3���d�7Y4:5�1�4��h�m�����rlu�rg둍M����r�w�7��%�1v��qe&��>F�f:��L
F�.�m`���95� ٳ+ �\k �b*)�mR*�	��rk�z�=��ޏ�`k���Z��]��WN�m��2�	5ư	/b�'u� �6�զ���V� ٮ5�I{;��2���U�V�ɖ�+m`�"�'ve`ve`5�um�{�}�&,�m#��@]�.�����èQs�Gf�2]��.�a�P��n�J��I6�	ݙXݙX�q� �c�J�U)�����um�`l�� x����g�ޮ䓟{���8g���"m�_��t��n�f�y�� �c�9#�&̬ ت(ݷe۴�Zm� �c�9#�&�`{��{<���*TS�6�E�>o �����zg��y��/|�t�Nr�z[}���m�6��*F�4bgU
�"m���(����2�C[5Kc4(�M]XX�]'t�V��G� �8�&�{���;�?�x��?�t�զ�H�X��rGMp�$�}`��.�Ѕm�v�X$pɞ�|q)!m0)B2�XFP�e%%%d01�E�!=�"K���eH�R�&�e�U���<�m�ƍ��ꉑa�Qjb��!��B�I��`	H�F�\�;����]��܄�)�씜��9�o{��K��s@�`��I^�q��I+m�	�����-,7�6)CZ�e�s3�C�ȼ���@��H`ci&@(B�-%#B�6H�����P�Cf��Kw��	L1F�`$�FZe�z�:T9 L��B!#M�>�tWS<5y⥡��	��`S�+��)@�� �IBEҡ��>Q�@�����}D^"�ȯ� U�g��nI���]�'�Iv/��un�բ��0=U�.��� ���$q�f�`&�d�L6;N���f�`G�6k��0����R�N�MB������7�6k�D���{388����m��X�U�L,�t&��g ���� l��H�l�T*+�خ�h�;m� �c�����G}�� ���Ik �u
�4����H�V��0��Ik 6lxWij�R���V����`5� �8� l��*�W��U�1b�!PUo�����yg�O�a�۠wN��n�	#�`͏ ��fV�kjZ�tR�O�t:-�j��V2��*��m�k��.Ch���8�.\�Ѳ�m���򻤄+mpzy��"�6l��$�5��˵H�Wn�N��ـr\� ٳ+ �8�&�g������S`�v�j�[���Oe`G���r,�z]��褆�M�v��/{����x%Ȱ=Kd�^+���N��]$�-���#�9.E�wu� �8�+���(��=�(P����R6T�1 `�
���Ue@�2B��9�AYp���%�	]*p
�&��ۈ�1�(׈i[)a�H�PɃ\gZ3�Nѳ���n�^�Y��K��6`���%���pu�)��,�ۡ�쎍o	�13���M�vf�[��c�:����i"۰��r�k��-
E�"a����,�,�F��W���q��3θ)�ѽJ����˱�f8:�2:�@�f�iQZKYv2�b,��s�Nr6]z(V07�ZPͷ��$��$��U���1�"�3ez��Ӳ�cWAI[xe�Xw\0	.G~��� '���Q
��4�i�iݵ�l�K�� odx%ȰF�:�t����wbl�$��͏ ��\0	�Ɨ�+�HE�w�6<��X�p�$��{�YH�]�j�]*j��9.E�I��#� ٱ�[ Q�]5vK�o+�i�V�Қ�\�d�Y�&��ӷM�y��.[��0��J����y%�� ٮ��꯸���y`����)eR�̬�������9:KũB�$`XE
�$�b�!!_}O���1� �nE�l�+ �
��m4�Ut��m��6G��X�2�	.Gx��ZAr��郺@�فﾯ�|��o��K���0�*�M���;����2�	/c�v8`���!q'v:���K�E�����T�x[�,v�n[�:�Q��1Yc.I]cft}���V�x%�Xd�X��L]�Cm� ݑ���`�e`k�`+�>V�4۷N�*��r^ŀl�+W�|�}����\k 6H�H2SC���t�[���&V&�� vH�=K�s� �K�6�1RlWn��X��X�諭���� �y`�e`����բ�Ţ۷lJ��<<�a.ћ��M�ϗr������SM�cJ�b3�[Ll�ʺ��mpK���{6L�K�� �oU�>�퉺E��0Kذ	$��$��$��,Rڴ��黻k �L�Mq�dp�9/b�	R�t�Ҷ�;�we۬Mq���+ �j�ԯ(B�Bd�,#,$������Z�)���R��l���$,���!���@�>�vnIٯ�/�6�˰���X;0Kذ�fV&����꯾��:G��Dv-�F'��z�p�Y	�5�hs�uڧ��	׹��c�cj.������V�߶e`^�xd����T�[��un��ٕ�Ir;�8���9/bͪ���e+�-]�ZWt���;�8����}ՀN���5B
⶚��t��v��Se���`ݙX�����V�Jui�6"�����`ݙX�q���^�}��}�E�Yۿ���Ȼ�yK�"�ǝ��0�.���,9���n˄�Y+��GR���:N{ol�gD)q۲*k����Q�,A�3yPl��),��	X�!
�a���@-�hj���I��a���c��f��=��<�V�W)c�d�<-BT+c������4�����nM�s<r�3�vWx����R�͂(�u��ڜ�N
j]����&����3@
%��OJ9Vۮv�޴���uѦ�"B����3��#�����+m�4��7�e`$�`]��	��[[*j�ZZ�.�`$�`[��	��sve`�2�|�tڴZC��Wv^;0M�X͘� �wg�զ��Ҥn�=_}_|��<`�{+ ٳ�w�"�94d��`�lwN�V���+ ٳ�w�"�'ob��m�J�I殈M�:�	V��00q��)@��wW;^yָA�l�8H�ks*�j�S2��|���;�2�	ۑ`�XP����V٥��������s������� ��+ �&3 �oU�D�Rwm[Hv۬v8`�e`$�`ve`;F�\�W+m1����X�1�ݙX�p��[*�bT'e۬d�����p�;�;:�����s.�lJ�l$��/Gn5��yp8�f��h�Es/:R�;���v�i	�`��`�� �+ �&3 9]��i7n��� M�;0�2��c0[%�H�֪1]�	Zn��m� �+ �Lf�}�� A�J�!]H�0��`�c6�&�f_��ܓ�;���?~��{f��f�:���}�ݷ�H��x%Ȱ�X˨�˴:��*J�.�0��r\� ٳ+ �Lf:o��+�h+�T	9`���A�&�j�3j�� }�j,M��C��JͰ�f�r,vL�I1�@N���ZYr�]����wv�7fVz��]�����=<�r\�=��|�J��:��7t�	ح��Oc0K�`��nɕ�vI�U��]7m!�f vH�Mp�7d��_3ꯨ�*H�U�$��LQG�־�~��9�g��m�]]*I��rk�ݓ+ �f3 7dx�-�*���䋍�8�c�;<.��U�1�W.�p��(N�7Vjۚ(�(]T�F*��<���g@�f3 7debKذ��K��I�i����7���G�r^ŀlٕ�l��\�C����Wt��0fǀr^ŀod��7u�0�괨�1;���n�K�`�e`��]�xiie�i}j�m7wm`�2��r�v�,��X�����  cɌ��\Rk1���i O9���p��3�MJK�ᴗZ��K�0"� B"�J��lHI$g����� �)	b�i]�!!8� B&a.��!L6�XR���Ád��j\�.2��qXB�ȗ�T�WB�����s/g;ަ������yk+�q���+LV�ϭrr��8�9��\�&��V)$��k�}�F0!5e�"cB� Bda%���&B�
�4�
a	EdBI�� >�HY!a!>�\��^�*Ҟ c#�@��cm�$8T��(���"� �(ơ+
#YY��FFnj�C4D��3#I4�L� �8J��Ͱ��vn�p���$4a���S|�6K���ӂF�l|�Og��t~�Y��ڧl�����}�bo�e��y�' �h�� ���f���)�d	$���<]\С���HB1I� Ԕ�aIX�!0�HA�FXA4)��	B�{`!�>	P"�s�7�D`Ba��!�Ѱ�߀Z��8J��H3�k<1�T�]*Z�{6���{p�u�H�CP�Fm��L��0�0l�k�En��X͒�5bE���e&i�LVs��Mݹ�v�w.�k��Y�s��6!kHp��)�*���&6�^�/<�^)�x���ǋӦB���y9�՜`���]�7K;����i1bGU��	KF��t%�%`�B$����\4#,431�o,�Q��=��+��:8��A`�:�T�%��̫����6�w.Ӏ4㷘�+���l��u5��s#�������"�]��@�ͪĖБ��i��\�=0�gOR�e��]�mO����� ¹ ���V�L,�hR�4c����H�˭)v 6힁y6|��Am+]��3Ult�O��g��U��.U�9��$�ϋ�m>'l\p�6wm�K�z��	DŢ��ӎ���!ˮ�����o6�Kۀhj�Cl5S[��3&B���|�+T�/cV�M��;B���gE-�"J�tf-������*�WT˄9s��u@��dʫ�[�:;�C�j�Jfv�FU�w]s�'R
&��`�'b�m�͹.Z��oS�.t7X&�Aq�܈�o��	�\g�mOgWAq2G
���I�l�R�5'5��5��� ���1e���<���!�t�ӕY)"��'[C�jCc.H&�^�[^%"�8���N��^[Wi�2�9jj�.Ԝ��-��n���aȸӳOa�ح�Ȉ9ϡhj]-��R�ԲMt.L<q�L�y۶
�C�-ֺ�h#�A��8Չ �-ګ�cY�&��T�c�vx�w3�:�,.��r] �#��i�v1�K�F;u�[����y�\�����)l@��8�v$�A�\�ͦ��ܤh6�Q���v������m��\�h�A].R�e$&��K�k!4ʄ�6����Y�H��nL�8�pP�E��5��&q�G;	�w�ݗ]hا/�;����y�������z]!����A-z�t6�1v��;�v8��U�v���U�Ԥ�ֺ�1=P*�xxD@~W�#�4PO�G��`���(�S��W�4P�G�ryC�Ӟ0���l�7V!3k]w��ܦZC�����7$c;Wq�eh�R�M0�lZ�A�YYRh.����XY�-�R�Uy�Gn�<��IΧ	��GZ�]����[d%N98f����øڭ5Vr�b�8�l��وoF�F�]�P�I�أa#n�m��=:���Ƚ �G��u��}�mpL�w' ����D��hL+M�I'$$�9U��vJ.�7G��@��v�S^����x7V�H�5�VnX, Q����9F;{�r/�W�q�{+ �{�G֛Wm��Cn�n�`�"�$�+ ��(�n��+eZ���;�`�� �&V��(�5I/ �Tav�:�t�ـl�+ ��`�R�{���1]4�M�Cuv�`�r��_|��� �y`�e`���@�UҿSui��ptA�zw��[=4l�n��+qC�ǘ��ZV��:�v�Wt��8'��Kذ�2�\A$~� �qZT{�j�N�&K�f��>���Q|i[5=��ٰ9��ۑ`]����,�[M��X�e`���� � mHGWE��TЮ�[�KwrQ�I0K�`I��vI�U���i�-Pۣ �8`�"�$�+ ��!�=�o%�o`��8ģv�4�hkPc��Z�`ˉ�tm��-rX�c��ٖ��᫫�;n�H�l�+ ��(�}�����V�F��.݌�c��f�L�w\� 7�<�8`�Gwi�E7j�ui��7u�0{#�*{ّ�d@�B.�}਱��s]0o�V���.�V��
K����%7�x}~��;6e`��� s��D��	�ACm��"�6I��n��Xٱ�� ؝]����%�P�U��fu]���v[E�\���yܗb��6[*b�՛f櫳z���g@�Ͳ� ov<��X+�GM��V����n���K=�}U����w��,�fV/�#v)��'lM��m��ݏ �����{+ ���X��$���*ut�+o ��6L�n{�w'
�]
	<��krO}�jg�Z�Lj�V�f͓+ �{)`�ǀN���B��;�J���VJw��C��W [�F"E���A�t�!��Dx�cwv�[�7lN�n��~� 7�;0M�X�DW)�'e'�Wt��0{���H��� 鱗�	�r�����/����.�k
����נrk�;{)`�c�8���)c���i�n���]�W��ǁ꯾^�<�ka�M�;baj��fvU��c�'ob�95� rSEmg5�p�k���r`
����[cfC�:n0v�&�vN|�9�� i��V�u�٬B�Q�@T)-�M�r��L�]�vRt���#4p��K*jM�D��b���]vі�j���"v��6ܧ��<a ;8�P;́�۶ԁ�n���X�k��K5�֧k ``2v�X��HN��s@�	q(@tY`m]�X�����c��5�S�m�LF.�s(q�a�kG4Z[v��G%ԑI�52������v�j�u} ��<v8`��N��X��$��[�WJ��x�f�wfe`����x6S.��*m�[m�;&V;�Q��;�;�����n���$�`�������rI��ItEr��vS����mрݏ ���fV6�R�?U}_}_lq$]xsv'q\ex��:�c��`s����n��Z6��s�uR&�`�*C`����=�<�M�X��ϫ��� ��_5��6霚��z�|������@c
�$E� 15O���ﾺ��|�K�*�vG�N�ŀ�tجi�CWv��vU�7c�'ob�9�2�	ئ�C-�-�M���c�'u� �ٕ�N��X��!2���:h�x�ȰM�X��K 7v< ڂ�.˺v��8�����\g=m��v��wi�+
u�-u�\3G��c"ہ�1U:�}���{�Q�ݏ ��;���[���n�n�	�����	��rl��$��c�����wWmрݏ}���nS�4��B����$ *�O�(�1P���ٹ'{�`:jTGn�&]*E��rk�ɳ+ ��`�c�8�wIT�];�ڶ`�X��J8Wv^�{ C@J�.	؝�M�TXμY��r:^s+�: ܭ�93q[hl��n��ެ�:hN��[�{{)`]�x%�X;&Vݩ0
J��M2�n�,��/6�;.vL�����g:��;cT�`�C�x6�,��+ ��`]�x6S.nƬN�un�X;&V��(�:���>���UU_e/���X{���[��6���	��7��Wv^�{ɳ+ �����j׎l�R�r�Mg�u��Wkt���x02Z�;�0�1��Tu����X| �<�KذM�^����	�=K ����۲�4�"���9/b�96e`��K 7�ʹ��
�2�v�6ݵ�rl��7��� ov<��,�$���v*�@��u�ooe,Wv^�{�ɕ�wjL���M�6�۫�;/b�9/b�7�e`����ZoK���6�Ϊ�������]�f
�۱���q�o\�zh��V�Xv=�-�&)�zƎ���:C�=]��yz{>����5�R���f�����g`�)l;B<k�Ӄ8P�v�(�G���ݳ%n���	#.�aݳŠ�:����sWe��i��18�t�1n�\\�"I��-7v���j�=�܇�N��\l�29<�����9���
p�x�"�xٻB�}��J(�O:�C�O8C�R�znT��׎�vϲ��w��,vL�w\���}�q�{׀wo�_�5cV'v:�m�vL�w\� �^�r,���:�b�m����� ���:���rk��&V���v�մ�+wE�F�$��\0�2��FūDj2�cE &� ��f̬{�Q�j�/ �
ߑ�FU�G�M2�N�m�\l�1�` 0��n���h9�ۢ@Dj�v�&�l�6l��7�����KذhlυJ�]�V��v� �����(�`�"Pb	`"l�R��=�}�nI���rO>��ꑲ������m4�[=x%�X&̬w\� 9���튛���ۼ}UT���,���n�`���.Ϯ�XՉݎ��k ��v�R�5we��"�=�-�.�����S�aw:ۂ�@���ƲF�œ.םM۶)���:�ه�H*�^j߀Is԰]�x%ȰMp�6]X��'Lj���v�`���K�`��n��XWV�.��4!m��0Hყ�:��>T�%-"͹�e#l	���1�a�`H��P��L��FB$0dS	B`Ȥ��-*�;I����b^���46.��K	yYm94��ƇQn���+"B�:����iRHR��ah�d�	FVZ�l[,gZ�_ן��7s� �i��c0����y�H��3� � ő0IB��$�d<B�Q*��!W�!$$�5�	2���0r��\��a�u B�i�iRR� �	�w"�l��#KH�*��n, � ��$tQ��RF2��Bi%a	��L¸�1v�  �A~4 � >D|��a�t����Q�D= =Q~�i*��<�|.�_=�7$�o�e�ϩHc�m���8`�r�V��\0��L��v�V�!6`�r�V���,�8`q�YIl�H-��σ8�Xэ�{\g`F�v�LT�Г[���EhG� �\֬:��x%�X$p��_q��F l'��+[�_�ۼ��,�W�$w�~0	.z� n�xg�
n�j�5c�v��9#��{)`�ǀr\� ��=���j�nWES�y���t�}�[�s���4��X F@� �*�H�����a�[�o5�s�D�6�+5I��ۣ ;��{͎�\� ���B���� Wt��!�sx�[V{N��Ϧ�u���6��5-��2�3\�W�{�y����N�`wc�9�����aLun�l�9��=_}�G�?Q�'�;�ꪯ�#v��*��E�Sm$�0l~� ;��������;<�`��)|�Vē�li�0�����sc�;�Q���]�U��I�.��'u� ��n�F wv<$��|`���&��Y�������ɗ���DP�غ���(!��&�-(����,͛!Y�L]e��3f��j��<g�8ՠ��`L���#�0�8Q9����v^^S/l������}���9��nuB�.s��W��q��^�Bظ��QgLne�9'�8�0#K,؍��c]���ZJ��Dn�Օ77+�
�-�j��t�u�kvQ��=�:v�������e"[{<����e ��Iq�.�:�3�}�}�~�ɘ�ϛX���V:��:�?�F�v^�r,M�)��Cm�6۫m��F��/ �ɮ�	we۫��ջt�]�x%ȰMp�7��WUjEϕ;��x��|��y��7����x6��Z!t����8`�r�V���,J�)w����n�g]���U�:�,TkR�0�#�h5��QZ�9��W<�8ىV�T�}�����w@佋�}U��~0�=��;`�j�5u�nI��߳~��@��.Os>���p�7���ؒ�튭պM]��9/b�9�� ��`[��-�\�1Ӷ�un�X���]����Fջ/ 佋 �bʷN�mRm��ـou�0����,�}}:�`i�5��-�t]x�j��yq�6���ݴF���t�O9h;[��mS&[��M��Wv^ɮ;0�F���"�2��n��w�rk�o�
[<���ܓ�~�I�'��~��E*;-)H�x�uwm� ���o}����d�H���# ���a#	!� HBB/�T��P����;��`�l��۫n݃m�������ٞ� �'� ���0�l�_?��*v�����:�e��� ��V��"5JT�46}s��7B�q��닚��fSfa�ms`Y�(����2�ln������ے8`��jݕxWv^��
n#L�39o@�I9�Z{}���-����Y��H��YV鶝۶+mӶ�)=W�j���9.E�rk��ȣN�v���7tݺ�){;��y��n���}7 � x0�X����@�p�@��.l����H��������m��r,�\0[�� �ݗ�h�Kai�K�]�Ζ��i/�V;y]��v�����nQ%��6��6V�m��p�5nʼWv^�r,{[.���Vպm�� ջ*�{���"�95� �ָ/�2݈i[-7W�ݏ �������`I� ��B)����-���r\� �c��vU�{���ݞx���o���۫um��v8`���'���<�K�`���b"�$�hMӦ,�G*d]\��&Ŋ鍹Px0X�X�����WK�s�d0o]��� �8�,`��3��\M��އSkY��6܇9J����P�j;|�����mwm:*���v�v�8��sx��뵔�l�����H7=p�:�P4�̨�c�3X]�T#��a��@��H�[17.ŉd �;
�c��y��<��ym�h_h9��uY�p������{�=��������<�߿������%�e��B��fN�۱8�\�!���	ssD6�Wm�m���~���c�9.E�������y��������2�sE�9�@�Ǟ���#�~��;��,m쥀ҵ"��v���J�m��"�9ۑ`oe, �v<�-m]Z'�ڶӤ���v�X]�� ;ݏ �{����5m�v�[�+f;rR��c�&�ŀs�� 9�*�5M;t�Θ[�t�+X.�İ����Ԁh��{V�%�5�vR)3�6�\���|���{��v䥀�R�i&�m ��m�Y+k믾�Ͷ�Nܕz���wrI�Zy������d���;���'nJXv^v^��e[��WN�V�ـN�`]�x]�x����ݙ� ����5N۵e�M�-�0.�.���m��:��$����}a p��m��{Ku��Pcp���3A���F�<�[�^���v;���X�������X��K��[�-m]Z'ͻ�I&��������^�6^d�v�^Pն7v�;�`oe,��/��� "� ��Av�V�%��`�9t��Ҳ�v�m��8����%��`z��������T�m��t�ա[�.�x����� ���X;{�
��.֙�i��h��F$p�I��Ό�k��"�is��%�E���5r��s��`oe,��� ��^����V�wt�Z���k �{)`��X]��v�,�W�}_${�yz�����)�t��Xv�d���� �{)`7�\�0t�������/_��	<�>�ܓ�ߋ�?( ��/z�I9��=[|���hEs���;������ŀE6^��˽+5o ���%V�����q9h��$ms�Kt����z��tOv��U�p1�I{)`��XSe����Wl6y�0~��.�61]]'n��,�v^�x68`^�Xٲ�)�t�n����w�E6^͎{���z��O^͹
��V:M�Ӷ����M�����x]��	ݕ�n��N�J�j���	����ݗ�E�/rNy����xm� �^�q���d���$!:�s����d���ggu�D�N�m�P��$�IϹ��d�1�0 �		���HDX#P�����0��H�U�˥ٲYHR]�ke���!P�Ғ��Ylh֛MBC�!����r�洚fM��b����$B$a $B�93)v���[$�� ��#D1P�l�	d����aF4�����a�$�B2E�$ J[ f h!s_9�����9�w���5�(���X�! �<�B��R$ �XR`@�"ԌD#D��BHHdR��I!!&CA�abZ�a!6�l&m���f��l���,���YRQ��F��nE�7���{��f��тܣ�rA�0`V�e5)��l��0��R��d�!!B!#�c�Rɦ-!$c0#	0	�h��V%�$X!��':I�_�o�i������n%[zZ�p��.;6O.�A���ёN�ʢ�a�6�X��S[�V�c&]P�4�� �R���[Z�ԭI`S: MWe�t���`[[6f#@���1�:��#�)�d�rm����;J���ã�ZƟT
��6�N�;:驜��m�m���f;C���" �8yŷ4��ڮObn��<�'k�0�d�
W��V������O�^��wR�ǆwS� �������ҙ5Ъ�Ҳ�v�\�s�rd�ۉ����>��B�9dV�g��r�n�Um&�nRS�ư��_h�E��Lo��q�r�5�7&سp��Ξ��H4�4��ڣvݮE�^�e��<d��v�v���tE�!�F��ѭ�Baбv�.u nlӞ6����߿���4n�uΧQ��l����3��n�3���Uo���Tz�(�uk�����f����B;b���$NS�k ����nR�̻��Jt�`V���7FԶ��̜n��ؤ���岖�a���JCw1㣢��hc�}���u�Њ�[��z�,WOaA���u�E-�\�]�
�EU؄����%8�L�LɎCy�[E��x뮱�2q�;l�]�0�rؑ�;�i��{bN�a{�&\��XA狵��V�A�5!J�\N�s�v�2�Q l��%�{�a�m;5<���g�*����8�u�[��)�;7n}v(9���p�nv(ڹ*���
)V1.U*��.��ၒ��zr�f�ѩ�RPؠn\f���S�MD��b�T����nk)ڐ{6�pgq峻FQS^�u<�pv��@X{:��f�M3�h���������V���N|�"���W�D7<�/&�Y�����O;c�����異���9��>�]sW�ɇ�a٬:���#,L^�z�+��v�٩`������n's����`���붉�lv��`���4s��CiQM�Ҳ��O+��7Z1ubyI\�ɰ����ȆN)�J�,ͮ�*ɲۯ$�~���$��I���?"��1Sj?"A~O\>P5ழz��]��ݑ�[+�!��]��-��.ܮ$���Q��S!�A����^Ė�Ө�v��T�����y� ��j�F/�2����;�:�S˱Z����	�5%ܳ#%i��li9��n%���n�����=��6�q���\rTn�Ձٍ��q]h�/a��qu��h4�Χ�q�����:�����9�������HNNL�`�v�fv֩�lj��a��b��.�ؗ4�-�b�f(k����s��ލ!�[�����t�_���"엀s�� �{)`6�E�ct:WV-��"엀s�� �{)`]�y�����96<�[�\_�0�%�]�<���:��K ����"엀oke��C����JـM�����x]��=���x�7}^ʺ��N�;v6�`[���%���M���T���R�3X�]IvWu8�ƪ:���n������ύ81�Z²�3��ZF�%cMͳ���^͎��K �ݗ�snB�)R�ʚ�]�>y��ߒI��8N5 <Ch;Tj�2~��M�?_z��%�ꪯ�=�Օn��jګ�ڡ[0H�Fջ/ ��^͎����)���0?|����[�^͎����zL��PV��c�tU���vK�9�"�&�`[���Z(+Te[@��5E�A��F9.&7�[l�һm*�^	��`{tHo�h�I�x6�X�r��v_ܒI�oǟ}������:᢬ʙ�� ��Q����着�5I��<�޼�N�䖞y�~�з)j�j��_~�nI��߳s�C��D	FBP u
;�f�ٹ'��]&��ﾒ�պc�����x[��lp�'nJXV��lI��60M���sc���U�wc�;/b���T���k,7.i�Pa�Sl���jE#n	K���YN���I:�p���,i�X����x����ذlp�7n%/�-�S���n� ;��{͹��U���ZQ�Yhm�t[o 콋 �܋U%��x�y��[b��w_0��������償_{�7$�{��ܛT��*}�>�����v�4ݦ]ۼ.�W�~['� �׀qI/ �$X컱6y�U����N��)z-��u���e�C�i�6.!L�v*9s7@<��^���Ix]�� +d���歃�.��"ݗ������#����[�U��ǟ� 戮�S��۴��� ���vK1~�ꯩ#d��<���H���m�wm2���d�-���e�l��M����I�t��ۼ ��x�\���=��"웠|��<Ƿ[�=K�HP���X]JA�`�,-��p��ɖV�+��z����nj�u�J!m03b�M�-#����M\�وrj���gnیl�.���fkX��Ƭ� :� �d����gm�R��|č�8���	�NQ�5lujn�t��D7clns/Evǳ�@&1�������}���(�E��h�l0L�iK[�YV:,A�l��9��F��L�)-��5���˗5�э��phc��'6dr�y�w<>��G�� �V��n�m�Rz�mȰ�%�wc�9���i!]D|­+n�lp���}��˳�^ O{��"ݗ����ڋ�R-�m]۱�6`[�^ wv<-�x68`�S,V���Lvݻ��ǀE�/ �������z����_��[wn��o ��/ �]�x���H�;����ӹS]�kl��.M��nʄ���O�����}�dܫ%�Q2�5`Ewv����z.��v^v^$�)��y�rK������y��'����{�]�x�x���i:�wwV���ݗ�Eݗ����.��� ������`�һ�6� ��/ �c�v^�ݗ�smm��V�D|­&���p�=_}U������Eݗ�I[IE��v$����C�E�eA�0t��s=�+���ٶk�݂�$v���C��l�"����ǀEݗ�sc�٣��E�v[�n����we��� ��� +d��h��mݺ��v�,�Ix�g�R��R�(P� H2,Hb�*���}�W���S���< ��'n�j�ݶ�)%�������,ޞYM���m�jڤ��;������`RK�9[E�-���%�u��8��l[	
J����]�-G�����sm<C����ǀN��$�w\0�5]Ҕ酅���n�g�#�O^����c�9��˴+����[l�8���"엀ݏ �����Jcc"�Sl��'$������|���$��u�ܞy��T�D�BE�M"���}��{��kX�+�m[v� 7�7\0.�x��}�[{=n�oX�x��3�(��^j&lf[�1��L�Z�\��M�R��ǣ4��m�e�x�`RK�"ݗ�� rlAt4ջ��t�v���� �v^�ݗ�N���URG�<��[��nڧv��׀uwe���s��`\J&�'uj���xv^;�;{���������Wt�����[w�N��܋ ��/ ����;Y�Ԋ�����k��͋,m�m�@K6*�-x����w�v�� .J$�A��Z��j�����ږ�n�Ҡ��H�'n:�=fvN���v�獜cԮ-��d-��܃n��ni_i퓾�f9�b�)�����J-���Z�����@YJy���Q�s�%ێ��lp��!q�{n���ȱT���p��۵7����;`��u&q���+�dE�e��$�}��zt��)�/g�n���<1��P�]i���nzt�·nQ%]���ov�=�zt]�xWv^;�{Z���i;t�4�.���^;�{r,���_*wL,�+�w�uvK�'u� �nE�M� ���_4]:��o�v� ��{r,n�`]��wT���Cm� �ob�&���/ �����JYq:N�D�74m����-��LR��8 �]��6�n��m�2��pl-�1��7)����������7������7o�A�t�T���&�SrN_>�7�@���D�����UUI�Kذ	5� &֫�V�JiYiZ��k���ŀI{��/ �m-��H�J}O䭶`��XSe�]�x��w��I+wj��6��"�/ ����$���� 9�*��wi��l���n�ۊ�[��p^������hy�ٕ�֞hIRv��Ս&���ݗ�I�;{�x\�|�l����wn�	5� �ob�"�/ ����	�P.�t�(v������ �v^����b)¸@�a=4���lע3��;"ը]Y ����� �b�# �����V-H���55���&��kB�i��D��!��1~����4��uO�H�,`0Bl���p�3e�frk�h��n!"V�C�珞�o[�g�O-�$(KL�˓2�5��fM�,h縩��&��Y,�K�I�Mu����=��K�!.�{��ng�`�FE�B1X�2Ɣ��$������"��o��)��DO� �_m�evȁ,�*�B ��H3F��l���G&kie��fZ�!�(T4��Is(aY�2|BŦg�4��%�1)r�7p���5��'ca{����,t7�w�a����(|�征��i�ӆ�)��SA	4���^q	kx5�f��<%�0����B|�O�6E# � H�Hd$�]�����ԏ�CC�<AhyT	& K=<(�0��ED�A�P����E���G`��QGJ�(|c}qT��h���# 20�BF C�� L �W��Q =@2����	#�6B��v�-�m�[k �v^��/ �������[�y`��/+�WLJ�X�w�qvK�'c���ŀE�/ ��V����v�H|s���\�㉷[��J�����V!V
k���+T��!�h���x�p�;�ذ�e�靖:�޼�iJ����ﬧ�M�`��X[��.�x�p�;��u��-�Ӱ�M6�7\0.�x��`��X���Г��v	� �엀I{��Ł}J����D$�t1`�@]��9�{������?�6Z��gt	/b�;�ذ	5� �엀{��_���-Uv�+V�!ƺ<2(*b���v�&�-�B�=�4���7T[g��H�[g ����$���/�W�Uq������n۷i[��T�M���}�RGV�^���s��`\M+�t�J�,� ����'c���ŀM� ݭWt��-+�*�6� ��;{6�,��/ �m-��H��Yc�&�0w\0�� ����{���$�$�|�OY��&���l �4Y�MWSl;r�qQ�z���f�V�z^�����a�9�ѭcv�nH�]�smoi+l�,�m�s7$DM�lP��fLl�2�Ď��E�ݲ��b�̰��:�ps6�k��ٙ:�X��Q�����I�6=���ˤ�)�k��폎�C��3�(4ۊq��1��[I�����	�tH�Tu�ن4-�Z�P8��4��nk$�RHI�m˃�O�ga���`���A�aN\:�Huqv萻`�V���V�m������/ ݎ;{�G�S��Кv���ql��n܋ ��ŀv^ş���x�c�۷j���&߼�m�Xf̬�d� ݊RC�2ݫC�m`[%��2�����Ȱ	$�ʷv��v�����2�����Ȱۑ`�(��*�cun�����r�n�P�]n��!�;(��t`����Jꕩte�nj�t��=�{r,{r,�fV N֫�A��d�k7$��u��C��� E"���4�? ������I�}׌�l�m��wIs�,$�onE�l��l�e�X�E1T�]�i�m`/b�:���6^ŀonE�vh�t�X�0M5v��l�e�X��X�ذU}UU^�0����,f:e[i4P�3��Jŕ6�r�B���*psl.�I���̱��0�w�'�y`��X�p�8�%��%cm����m`��X�p�8�%�/b�;�u�ڴ�ݷwLv��\0.�x_�����|W�)	(B@xQ�%),��,��� ���5mR�t�v�m�d�e�X{{�\0mj��DӥeՉn���`���u�.=���^��Q��E�U� P�Y�"\K���®籷dOA�M�/ؚ&�mG��%�^�����绫o�\0.�x�ذ�E1�MջwI[�� ٮd�T�x{{٣��ui'EӶ�ݵ�qvK�5M��w��`5� 7����;)�ۼT�x{r,f�`z��R � 1H���b0�G  {����!�P�6�4ݍ6� �엀l���^�l��_|���W^tӦ��{p٬���^��S17#������X�f�2��!k�]��c�h������uvK�5M���︃V�׀{���U��YvՖ6���^�l���^�\3����$ډX���T��� m��� �엀l���^6�ڻ����E?�M��:�%�/b�:�%����;�J,�&�-Zb�wn���`]��Se�]��	#�E���@�V��\2\��ŧt�G(�ݻ�x5q��A��CiAμ��6n�gK���]S���/������T�ힶ��X[o=GG1<�O���s���m�0�Mi]��=�ղ��v��Okr�?Y��eM%�Ц3B$
R0,�*Z��;%$�c��4��$���#��8Iʽ�V�b<ݸ���"Jn�v���K���q���
�H�lk�'1]uD�𦛤�kY=__PC�E�<��qr����ܜ�ח��t47��td�9Q�ld�fQi�xK:u�&���ef?6:��^��^��/ 콋 7v�[�m�0�w�j엀uvK�;/b�:�%��%cmSM��2ۼ��^�{�KV�׀M�y`����7n�;lUm[���,��^���ݗ�M�"�}i;(�i�����/ �܋ ����;/b�6%e�$��"�+�R�*;v��&ʘ+g���N��-:���0�����ۑ`]�xe�Xd�m���[nO�6�kWrO/���؝H=9I$���ĒHB$$����U�UU`G�.� �܋ �u(����mnۼ�fV��/ �܋ ����6h�];)�`�wv���6^����^ٳ+ ջ�h�J����������^�{�6^�6�Yn�]��ݮ:��V�0�C�rX�`^/�{ViK-!�s�*n�1��7N�v�\-�� 콋 �/ �܋ �"u�`��*�����,�l�{r,Wd�lt����Wvݖ[k �/ ���t�H
�����rN}�}w$�xz��wwmX��ۼv8`�%��"�:���'m-�bIYT�Jݺ�5vK�;.E�uM��n���?}_}���w��L�fY�f��0:Ѝ=[z�la�O��-�,��Hۥn�G<��v�w��,�l�wfV��^�ӫ�ӱ�������$I=��E����"�5n���-Һn����7�2�]��K�`Se��%ccn��շX���>��I���f��������\m�B���+�Ia#1�Z�
�"�E�u����;ؓ�hnݡ1ժ�����X�x�̬Wv^ mv�4�PmƬ��hq)UڼI��hZ�A\X���#�l�M�����ٴ�Uf2ށ��� �ٕ�j���9/b��b�+�˿�v�[w�oveg���"-�����qM��N�[J����}O�n�]�x%�X�x�2�mE/(j���v��{ﾥ�9�uzz�	6e`�%���WC�������着����@7޶��V��QW��E_����DD�����
��� U�����QW������ �T )B(T"�B0T �BT �B
�P���AP��(�P��B$�0T"�T �0T"�AP��B �T"+B
�T"+B"�T AP�!B(��T"*�P�B"���P���AP��T �U�@T"��B(�T  AP��T"��B*�P��T B"�B �U �T"(�T"�0T  ��,*,�$EB(���T" AP�,�AP��B"�P� AP��T ��P�,�EP��(�T (�P� AP��AP���T �$� AP������(T  B(�P�� ," $B
��U��"0T" �P��P�AP�+B*B�T")B(�
AP���B*�P����P��P��T $,�B+BP��P��T"0T ��)P�,�@T"B��B @T $+P���B�T �(@T"�UP���AP���P��T B �T"�B �T #P�B�B($EB*����T"$BU�@T E@��*���@U����QV�*��@E_*��QW��*���TU�(
��� �*� �+~�PVI��bm�?�d�` �����aOW�����
��U`b� �e��AMf���Y���E(B=hU�AI�֠�C���� [��� wj ��gw4H
���]��ۧC�MR��@9� t9�@ :u�ͨ����4�t��    ��
[j ( h���:^����}��y���צ�����:[�|�Ν���������Uh�uNZ8� �\Ǝ[�n�����ѻm�m�����Z���w��t��z�����>>�{�w��=������[�� ���*l�}�s`.�� ��@���W��|f��oOm_>��[٨p��mv�P,�������}އ���}����ptf���5\ �{��}�{;��[��.g�n��>A��۪<O'm{�7w=��o}���t}`����-��ѩ��Z ,<{{�>��]�i��ws��{�zz {����Gw��K΀sҝ7�Mf��)kN�׽�l��t��t   �� ��� �Ξ�4��� ҝ�N���� x�Ѽ� 6��I�yJSI�秠��nSЦ�;�=4��tӠ  �Ƈ@�U
�ׄ=j^�Ҕ��]� >��݇��3`3�]k��(s۾���:�s�����SKg7���c�= ��`�����{�蛾y�o0���`�g����B���}���<�y��}���4p<�7���h���P4�{j<��o��t=�3���i�o�]����/Oy�{��|7���|���8�� ���N�����y5�B�w��q�w��w��>�⏣'���@��97}���  D�&��R�� �=��Ti?Ҧ��Lʢ�z�SL 5=��)�*�4�� ���I��J� h ���ʕ'�j@�������X�����������{���;��UTU�k/������UAT������ꪢ��*���UTO���������;�'0�i�l��_��g~�4}#K*5���Tp��}�?���\�mQ���o�։�̷��O���%Wxl�\�F��.$*F�@(�E�i�Ȇ�	RHb5!Q&��W�n�0�\!M�Nѳㅄ`Q�k|8CI�ۢS�J.���'7�����T�HSz�N��x��D��cp�7����~G��L��~�9��h�1�L�)�H�HU�DaBR%c!!�U��Fj����J�p�?��%���&d�.c%���3a�p�a��0�������3!��W���������d޷7HVFׅ>^�~��jB��E;��^}���>w�^V���B{�Y�y�s��������{�ŕ��~5��W0�g���/�P��3��+3/�WnR����K<����f�m�^h�)��`B��(K�]��M���~&���^B$����8O��ri瞏���w߳�+����1|�(��)U�k/~��W�v�����Wt������ov��J���E;�w�:*�ޮ[�p\�)s��w��rg7����4�`JČ(D�*Ji���#`S��r����彧Y]ܼ�_>�r�VU	[�]�V[�WZ�v��WMWk�w/�gs����=��5=U�}�ՙ���}Y���N���'�w	϶N5����¡)���lʹ��k!c
²�f���f�^Y,������_lW��Q�v29���s6B��?��\(O�}ջ�i�Ue*T�+�W�'s�*w�;ϖn�|�¸v���߳��P��{O�%�Щ.�p��	YbF&�0�qc܍1�\%�͜�Y�����j�0�ßw;��~.ψ�n�����焔Ϸ��^Ͽ&����y�\H3\>%#d~zh��HP���������~�6��tB	w���&��?kF*U�s]h�|>�t�����ҫUJ���Â1믡r�me��W[�����w�_WI���|\8����_�k6we>3�f���ދ�>���Sg	�����{[;���h��TP*�O*��{������F�!����Ϲ��~��/�!�n^N�A_}}���p�
�QG*��)[YW�ݛe���le1�4n���P)��6k�?v?��r�]�G�Ǽ��K��9�?P�'�GͿ�6�O�pwFw��������_�����
���-�J�D�yY���9���WG�c���tQ�p�J�6v�!=q��)�=����1�i�+�cBk����f�nq���'쳗Ë�ڥ��UJ���;��Ӵ����:�wVT� F��N��R��˨�]u�}��*�T��}���:봊K(�.s��44d���?	���Y���KϦ�+QM}ھ��f�Y�e;��P�+�8P���U���M��������_4.���2�b��}\-��}������.�k�θN7�^��K������.esI3l�	����5��~>aaIq%2SB,c �E%�?ew�T������|���B|B���!� a�7.���u��og38fŁH�J�K��n~	�t�HT`�,	)T�L\S�C%Ԛ���:�}��fv�����_u�U���>�n��ԻX.��E�*���x|��EY�B�XU�)ۡ[�[�f�]�O����|��ǜ�6�r}K�7�\ޙ|P�_$S{Kﳵb��妵?��{���]~���޹C��#�5�?B���0!L����J[�\S�#9O����&�"~�f<?@��Ĺ��+ă�4l͒���>���xv�}���k����j�����2�b�f�s+��yGm�@���(����CV�sQ��%��N��o�)��ɨ��-:JbB�ibAP��#T�S�ό�����C3|���l&�|\4;x~'�$������kws�Wa���KWT��G�Y�N+8����������W�.�����/�q.�ԡ��0�&Zgϵ�e�ZS��Q����������,	sa��\4B��J��H�vʹ�i+��[$	
�+�LH�-�<Ɇxn�a�w��O%�ga��咰|��g���/�����p��RY!B˟��gk�)_k�"�e�+����U�Gw��{Ϋ����tu�ܯ��ﳧN�[�g�>%�C[���#�ܷ����}���&����߾�:�^atW�]e}���Ю���VQ�N ���}���ݯ�ԟs������)����׻�^��݅���ML9���$!�.~7�xp�����B��$*B�F�0�	H\���%1�\��!Bq#L#B	LU�X�@���4��#aL�1�1%�R_ߵ��nϠ�B$5�F����/��M���cy�����_*����V�>u�w}�����}�O�-��%ndd�S,�\ ��	C����7i.�\�J�e��fs!��䳗�JJ}����ފ�qǇ��er4���!��қ^	�PȓHJ���RnGWߊ��	��\G��+�~�>��U�E�f����2�4�p#X�����3Fߣ���vg>v��\4K�3|�K�IVw�8p�А/!H�0��BĄ*B���A�F�W�V.�՚SG�tux��Q�o+���}]���÷���_׹��M�EUaK�_;�΋���X����ݐ�F��$�5�f�IvB�Hj8B�D�!(@aѸ�"`�pt��+$c��iٷL(c�f�9���� 3N�s���h7�I����F��7���$>%0��o���x����� �Lu�����|O�*q�ˤ�9�~�y�nb����S��r���7�
㡅��4�,��ۨ�������t���N¥�)ًm	��|���,��	.&�B�
b|Is����"B���]|~#_�.�o{)8s��B��9�/%|�{�y��a
���.S�83>��4�k�ۛ8]��	?s�F`S5����j�N���8�/+���}�>�}�V�sL��5��2p������1�5�5�j�[~̌7���G���.i�����ۇ��/\{؍ό�[7�q.tK���g0��yM��⟡���W!��kޝf����(��g����_4	����+��3j�����p���w���|w��=wT��>�u�fw�W�|��yɬM���ɟ�f��2�6�.2�`B��!q������~�^Y��쟏��X�{^s�����n�9�6e��:+���+:Ք��>��ޢ�*Ք��(}��a�I��ߤɟ�~�ן�P��V�����
��-�w�k�ϟ{FG��������Ot��[Y�WH������D�����sd��f��M�L�T*�W�..����޺��'�ggw��9�
���z���ծ����w噎u}EQG2��uj}�K{��et�y��/!�D�Y�f�f��͘\��	�W�Que:+��{�]���6��V�h��oL;�j���>�Ϩ�O�[E��:W��ﾡ_�n��+u�JYy����f��ѝ��li�~���h�H�;e�]
�y���c+�ן
�}���]��X�gz�)<�)Vq��1�ݘ�ov�,is?u�5���	��t�[%����7�^��B�TW��R����ҭ���т�/��+w��첎��J���nS���{�sv��}��X����sg��%vS������dsn|t�]}A|U�x>�����W�����\�2���.o�,$ ��Ry���w���?k��\~:B�, F�j4�7S�Ը:��oO�5�����M�p"����$�y��}��YU��6�Uۢ�>�|�+��|���v�*��^�T�/����ƺ�w>�m}ޡ��{���;���-�m׊��K(c�f����R�J�[TRy�2�J�Sޕ���嶖��̺���'}M]���Uu�÷��o)��>�
}��>������G-,���}U� Ϻ�z��^1��:���s����
���)<�+�������	U��>s{�ֱ��
���H����euw,�e���%�w?K9�5�^W~+�_�B�e�W�O����w���Z��)F��3�d����a�^o�LK��Hv/n�Nn4���.$�e�\e�c�:��0Д�c�J�}C�t�n:f��ߵ�)QTu
���		�.n�uZj;֗�9���h��.L��T�Q� F���9����e!ġ�i�!W�
�&i�ScD�!Yi+b@��'�Ϟ�����M����F���_w���w��-g��}���]�޹4��l$�!����4�#���V
�p�1���NlѮ��`w�X9��������+�+\)�M�9�O�c���j�Լ>|�U���]����N|���_[�mg�î	,8��PB���c3Y3��$(A�B:�͜�V?���Ik���k���̼�������쬷M!�F�鷏?�e	f����R�wu�ނ�.�r�o1���Id-�]� �T�P� X�LB�h0�� �Ѱ�q�!aI[�����>��WJ8+gW��{Uw����oD��_m���g����Y'�>­|�]��2p_*��k��H�^}w�s7tNgp�$������������1k���iy�����[�Wv��}�����~�՗8Μ�@�<#�YÄ([H0���!>'.�#ŀT"�A�+(D�G�w��3G醈\���%�ѽS�����F�I���~������:W�
�V�-U[���]�!9up��w9
���7~�{xw�l����7��Ʉj3U%�F$�Yh��	K$�V�瀄ڙ�#wY�zޡ�%\������!���4��1�E�!!*@�,�BK�ʴ��F��%%�ؔ��F°,�dB�����F!���Ma
A���)(�����G��0�%a,��%�������{�4	{�)��c�IR0�@���� S:���t���0�!�'�w|�9�M��?�Ň��6|�?~�������n��HG��eIe	H\4o��$ٽ�2@�8.%0�yMo p�`5�!H�0'5�sd�����d>���|��.2��:�ff�܉���h�?�&���)�Ir[�7���~x�njs{+�j`�N�������߾�
�S���m��_U|��'��-��}��Y�q-�>�����,��1R�O�U��V_��͵����p�k�ňĖ4ɯ�?�k��l��;ƚ��j6�!� 5��P0#r޷��r��k��|b|ˏ�_g���<��;���0�^��?�a��xk~6����K@�Yr�2�>���Jyw���ўO�3��~����;����'h�B��"CbBH��*��)�
��Jb �$I�,`� �,$�(�����J�!8H$�1c0�c�!�D �j`肔1б�3[���_�'!w����4�F�hه�?��t���/8������:��s�UӢ��!7w1ӷ>7���s�C�9���]�6۳f]���h?G5�r\��#��F1�~X�������0)�4Y�jn��\՘@��`F7A��K����K�e���7&�דp��ô��UU�����������UV�������
����������U���
��Z�������ܵ\�ҡ�[�'���\��譋�V�ڨ�y@���)Z����e���T���e_�U��vҒ�UR�kE;$��ԶNXȵ@]*ʵ@+�;j��A�Z�p�`�	5���5U[r۵uP*��.�C*
�FgA�W�_Ps��l��ƍ�6zn�Э؛�U�X	0���UJ�+�=nX �I35U@(n�W�C�Cv8��bp�J>�'���71�]֥�W6�,�@���u�-tk�V+V�ϕg#Z(+u� �k�|�}[��\��9��lP8	i�ĭ�M�P;09�؎�9��is���f���{Y���=a��b<��<�㞗��^�v�;T��-v�<��!6�{m�{6"�|�=�m�N��l�y�˶�q�p�ꍴh�	}���U�V�K�k��nEd����2�۰+��v����*�P-�Ӎ1�P�%N����b@�cv�l+q�ɱX��p��v��J����WPqJ�����Uڗ��FZ�e@{:s-�U�jޞ`e񚶪�Ϊ0�Pe� mu����UAUP��W���S�Ɍ;QXHq�Iu�K����K���E�,�!4pH��k���j��yXԻu++J&�j���c�gc�T��*�����ul��,��jr!ĭU[7&�O0�ц;oeX��8�z8⥂^v�lYn���j��n#�������1�%��ɧ ��Dq�wX�A ��I����	�,\���-9f��蚓u�`%L�d�yY�dc-`gkWh���֬vm��7bݲ	�]�Z����{;��cF���Q��n�A���v�=Rq�4JU�8=:��&�rD����y��xX9ض֙ ]�qY�\y�i����Ȳ]��u �U�"�Z4��V��0SɔەcWZژ�0��P��U�1s��V�-��A`1�S.��4��K�Al8ʶ��#���luJ�UVÊ(qYmd�Cd0� ��H��iV�
��t�UUD\�,��vgEU9�ٍ�N��qUVը	�����3�e�!niG���"�^l�1y�����iQA��:5�n
�vL����d;��͚�r��/%J��\�3��N'ejͅ�q���������<s��Щ��A�­�n|v�^-U�XV ;,����UFӭ&�`�M�(�z��i�mQ�NC+sl�f�B�p��5֛�R �䗶��N7�m���J�J��ջV��&�q��쳥Z�I����`9V�p�E�\�8��s#x��j�B�<Mհ2�
V�J�<��U@X8�D���)���o6ԖU���l=��@�zձ�lʥ�+�-,(�6סP.�y�
��V��Y�wi��-R�u\&�ۍ������t��w;�m-�M�����h�q���,[p�H	P*�.�5�,n��X�Yk1P� AYl��p�P�b���A���.i�
�[*�Q�lPRR���mlMǴAӕ)������h��pqR���`2�d��=��/WTKZ��n�p��u� �[��s:�+�w�}�mO�1Uj�v��x����vR�+��U��m�X��3QR4�@V����ݠ�k,�58�۸�ZE��,eS;��n���7cX�-Ik�1�f*f\`�Ƥ@Uշ�,ɲq.����vu����r��΂�&B�e���LO#E/=Eѩv�0
��o\�`.[v�V�W+��s��� ��6��M��Agm�
� p.9b�6��f+F�*�We ;6xҶ��qW"��C�gv�9�\D��[p6M$�¹of[P�:���VNd�/��1�b�F�7M�+9�٭�z�;b��/e��z�WUOKE*���]����&`ظcY֪�`�0LmP��˘���Zط�|_}��v�{��T!���W��^@� '*9��q*��H�@�����@B�ԩ(-�n!��{T�J�J���� b�4en�V]cfQ� )GC���'�޶���`�;l�Y�5S.}�y��ɠ�h�MU]��1՗9���-�E��O`7>̮�kj�X`Y���}7���g;��.�٫����\�&�uc�U,gӣ"�R���85���n�#V��C�PpVP��[�g�Mb�]A �CFj��T`�:��.���D�"qj�I%�:���)ѷ;EN�S��;�v��S��[8n�2ҍ4�%4#�(���`��r[E��ڣ�����{9�	�x�6{SUs��e�^�c�wJn�I���t^���ŭu����VGΔ,�kUU���L�X�]��$p.K'd��V�X8٨k`v����p�oa��L��(q�tAvٶ��)f8{pL��Y�v����g���j�h���jB8�:H@t=me��n*uN-���x8�""��q���u��%[�۶�UUҭ��j�b���{v�JP�4R�[�pAb���L\g�wV�j�q��ж����U�
�]T�㮲�uU��0�� ��UU]y\����mUUUT�UUV�@UUUUjUPM��
�l����Vy�!ԭUR�Lrm��U*�U�UQ�8�*틩y-���Z�v��[pG$�<�����=�d
�v�R[n���UU[n� �mUT�<���U���e���lܸ��j�@ڪ��U�
��DUU^UFԻ/]UUUI2�m�%[�
����������*���������L��(��L��e*�UUƥ��V���mJ��U@]tKS֕�R��� *�����+�̺D����U����=�lpM�-�Uk���q��خ�s5 mU[V6T�Ŋ���V�\k�T�4������7��F��n[��Km��G��6� V![� �m�[J;j�/G�/+UJ�T���q;s��v]5y���
Z����8
%Y�z����UwGI�ݥ.X�f��W�D lpmHM��g���U]N�ͱ�S.� å�n�S��wq$�]��
Z�N)��+�[[�(6��Z�C�����E��
�6�"��L�6�Nڕjv�WrxV�$:6��;�v��;+�-l ���@����Ͷ!k5��se��T+v��c�aJ1�O��[x���ፅ���[���@i�dj��.�.8�ѧ��0y���v��V��ֶ�<�@�Gdh�٭�:ϱ��F�h��5!�6 h�xAi+�V2���m��5��ig��z	[tJ�[UU@S-ٝ��^XƢ���� ���;�Zv��K�n*V�s<k�@8��ݺ&��=�L�JZ���ꃩV���F�i^j��`��c H��1i����m�*�T�U�juӑ�
�`�힠��wfb.|��U�\���
�	�RNPN-��9��4jL��lF�STUT��GKD�5]��d��9��R5�Un�ꎸs�A�Ó�st�]U���˳\UUSn��Xપ�z��ym����j�@�Q�yj�j��m�^+��ywe�޷.� *5;@]j�Dt���q��U��v���Z� յUʙ��TpGV���ڊ��2��V�ڠ��k7l�]P��q�@.�,��v����H�O)��q5mյPnFU@�������@���O:�J�[�uZ�i��:�J�sҔUUV �7��@ۭ��K;4�g:�ے����6������*��j4��#�f?�j��ګ@UPma��\��IP��O�z�c`U���,[`�@�mT��.��[q[[M�hb8�t檪��
�����U�UR�QU�*5R�L-�+j�ꪔ���z(�[���[�x�� �͜�MU�mUUEqG�0n���Uvʪ��^cj�V��+PV�r�UR���hᠨ(*��U*�UYJ .�
���RUT��+jڪ�T6U�VT�ch�^ˆ�T����� �T ��uGd2��UUUUUUUUUU]V�U�Z��ki����.��
��v|� ��� �-��UP�v^8*U��UT]W���UU�k�iɶ[]l%UƠƁ۪��SUWUJ�UUU��������Ub����X�X��n�
�����e�V��FNj���F�m��4�@�c����U kl`
�kn�W�T���[��^Z�����	vz{����\�x0,��T�JUUUUT�UUUUUUUT�UUUUUUUUUUW*ʵ*�++UT��UUJ��UU[@UWPUT�UmR�ʪ���Ul�*��X����b��AV!�+i\mUmuQFq*�T��0W-[UuUUUUUUTґ��Ë�f���5@\쪶�U�U}����ж��%��[V�T����Um�Z��Z�Z����
��Z�GUmUU�UUR�Um�ڨ ��n\�����8 �-<�U��^������� ��3��A���J\�[T�UUJ��'��&z�.�U*��\J�6���J�mk��@��*�[U*�USj�U@UU@UUUUT���۬lZ�j
ۖ�6A�=K�+UPTUUUUT���@V�]G-UVQ�ꭦv'2l[u�P�Vܵ�W�DI��^[îݶ������^�(�ƶ�Ȫ����+��WlJlW}]�i��� =���L�sH[��(��*�Y�[F.�.�j�����Uv�*�[J�6Ե||���qUUtl��F[y
��r�t֛����n��
�a\oaC�b�� ��v���w�ǵ��yapz��*:��vh��Me㤷JU���ظ1����J5U�s �=p���`c�Km��LR����@�PQ`�gl�o%�"Gb�8z�%�@S���ڲ&k�!��긯��{ʠ�QF���B�������(���?� ��qb�H0QpD� ���D�`��8� �V��PP�b� 6��� Q�J.	�D����6!��H.�x�S`PޕIF��P �	ڃ��"`�����! �#�1O��0+��6tjP6�
��~~�� ��	�S�N��tTN����W��B�LS�lR� �H|6"�@C��H��uN*��ژ�!�h~�����W��8"Cb	�Chu�*|!�D`t�E� Sz�"�74	Pz
mB 8�:"
!��h ��ࣥ�)ŋ�'@:(�`�C`�|
����8�'R����%��H�D�F)�*#A���d`@`
D@����6�*��B,��4 �OʧUS�	��P����I�a#!FE�  �� I$E0ȉ�"���DOȡ�EW���*l�I$`�	I Q��$Y!$�@� D�m �ڡ
A� �	�O��LV;-��6!B$!!J[+��!e%Xda *��������� N��4O���P�HT��&�0�?���AУEC��M� 4�t�/>C����������_�+Te�`� �)T�Q�H�hEiH��`�� B��0B�+�gڶ絩V�
vV��N�캲k[St�ԯ5Jl�[K��,����k��1�؞�j4�1���][�*�8��nƐ ��F�HJPvx�P����W.o=�*����Ů��H#�N���,+��Cn��ѫ��k]e���#]ui\�됶�p�=�� �0t-3.�%�4�B,�7m�r`r��E�*NĠrh�^F�=��q�ie��4��e�BK�B���������{�š�n��>SO@m�]q>�P�Q��%���y����[ �9;c�Eg�/n]%sJqĨZ�p������粂n����ۃ�: 7��P<\��ͦs�]��7�x�𠵘��.�1�{W%	���i+��w�`vx��5�I�p�U\�'E����ٕ��ey���gF7b��.a�B���6�#3V����Ze�8�'����f]��[S�E����me�4���;�T��ݱ�:��G#�Kyc`^
]-2v�-���^Ch��5v���r�<i
��������w;u�Y�κ.;	��=�J�4�0�X�� ���lg���A�DE�;;�b��zm)Z�{v�\��1�s��Ps�JL[e6�ødi"�p��p#la��`δ��ÚLէҕ,T�k{�s����e�Z)�Ɛ��͒5��84�6�5�x�{rscMW`���9�mn,7�}<2sv�d�:��p���d5�7ilnî�yM1��6؝��&�'	�-<�n����ɵl�E��G<�x��Csڀ�I����a��C��ŵ�Fp�;����y��;��Z���<��s�������ΙvUU�G:�{�.N]������n;p��uU[J�H*�ձ�A0I����fE �A��C-m�j���f�8�J��ĦGl�v� yH��Z2�����fU��=�TE)8���p�(�!�f�L�R�l��mz�wN���٠�{0f�ͥ��8�m�3����Mh�i��<(����x��Sȟ�0Q�tR& �U: ~?(D���|t�m�<aW�β�jc�e�4�*U�/L!5��\$9���ڇ����<F=�a)1kn٢ sIrD-хp����瞖�4\Jl�읲EǓN��99��1D���h��H�z����'=��6X�kř8�0ى3,F���C]�[5!q`�v���=�W�Nn0+mcq`�)�4\C�-�9;b$�3R��4�.e����V����̷fI�2�RَJIJ�`�C@�$!`K�m.���Yt�S��&6S66�~��7oF�����+� �� W} =hM��H���x�"�$�)`\� $����;�v��˷N�X��0	.E�H�	.E�j��*UcN��n�K�`�<K�`G(�&�R���E���� �G�Ir,H��"�=7���͆�e���hC4�d( �n��n�wR��a[3+��[���k�tZ-����� �9F��I��	'Q�4Zi��m`G(ϫ�(�B���eHDc�$� ~r���*��f}x;#�$���wW��t�ݖ�1;t����H��s�{��,޿z��K�+�j��iZV� $��\� �䥀E$� ����m��+M��x�"�$�)`I/ $���UM���M��l�m�0�SZfl�B0R����2$x���N�u��7�vj.��"l�-���K�=RK�	$x�"�5upۊ�*��v�mۥ�E$� �G�Ir,K�^��NKO���\�4�
��� ����$�s����4@�$0�`,Z��]���nI�߻��~�{�wF]����7E��	.E�I� �Ix$� �b����V�t6�X�%,)%��<K�`+��uA�M�9�4+�Ѐ&C���zGg�q�q�Z�R׬��c!/=,<J�d��XRK�	$x�"�$�)`(�n��5c�iZV� $�竜�U${��,޿z����v������Cm]��Ir,K����%��� ��z����G8ț1�z�%,)%��<	ʜ��
����:�w�f�w$��Y�v�)�Iݶ�v�`I/ $��\� �䥀���j���o����d���ʻ Qqr�Y�kZy��.��A�r�6�L]iЛ�V��{�x�"�$�)~���>�}��}��C�m�^��$r�K�`�<��N���t;M�H��"�ԑ���}���<�ݴӻ.�\�V�+���������%Ȱ	#�`(�n�4퉍�J�m`�<K�`\��	.E�]s�h��J�4T�]�ä��g�p݌�s�]e�rkfȌ��6b:	`���,J�Xm�02���vy�v�^�ժ�6�N�9��v$��h��4v�LǣXb擭�[���)18�liN��r�{C��åG�H��=�rc�ֲ�˯X�-��d�v�ಸ�'�g�px�8�p���y��n@���:.�~�\w�=���ۑw����4����'9	'$�^�0)6�ʕ%lR�a�fen�ͭ����]`.�$�睠43E����/����-��\� ��X�%����6'v��˷N�X�����W=������$�]��*��v�m7F%ȰRK�$��䥀I ,m���6oC�$�����n�����9F%Ȱ�.���v0wM؛�K�`#�`\� �$��9�'���`��UR�6���h�R�HMCs:�a`��)��uЄv�!1+�!�ͷ:];un�k�'��F%ȰRK����������o����OH���Dܓ�����a����HBBB1���V��d)��0���BR@�.��7$34�  	�"�A�#�糧�ٹ'�ϼ���0�U�um�v햬V��Ix�"�6G(�$� T�ҡٝ��\���ߤ�9�C<���$��Ix��cM��t�˷N�X���"�5I/ �����M��V&��9+���kS�KӲ���yD�Pv�ۮ�t��m0`Γ�m��� ��X�%�\� �� �@XҷWn�:t]��j�^z�#޿y`�~� ��XwUEx]�춆��� ��X��eQ�B*D?(��+5��v�I�����;؄�2��uhn�i��l�Q�Ir,T��	.E�}�.��eյe��I�0	.E�j�^%Ȱ��:��}WSga��f#k��q��� ћ"Pb5�o)���dlK�&#6=�A��m3kV+k �$�K�`#�`\� *wi	KN�*�vݻ�$�z��"{��`��� �$�TU��M��42�Ӷ��䥀Ir,T��	.E�DWCc@�cN�۷K ��X�%�\��*��T�K����	�B 9��8]�;߻%���L��]+�m`���z�ʯy���'�ޥ�{����<�x��.�3

�sx�4�y�nz'����q�n9t��j^��[9�g#k�����7bn�޿y`.JX�"�5I/ �bJ�L��Zi��m`.JX�"�5I/ ��X۲��WLE��N�,K�`���Ir,e�K �E[wQ���v+.��5I/ ��X˒�%Ȱ�v�Ҷ�*Uv�w�Ir,e�K ��X�%��.��WˋM	X޷��ch��+��4�t�*b��#�ʉ��4����)έӧJ�l��7k�*֊s
nBv݌D�����xˆƔ���SܯiBQ���b
�ب�U�֑Ū�!,���F�d�ejK6���G^�cv���m��l�T�s�����GuÉ*��[1vy=52m��;X7c8P_lt�E^��\��b�Ijf,��{���Nd��)R�S![�3��r�<n����L^r]�v�[O8��4�iv�m'TS44Yn�?~ǻ~�,K�`���Ir,"�v�ۻm����$��Ix�"�6\��	6P�j��I�ݰ�k �$�5)w%�$�����%.�� ��^�۵6�*��]�۽׉$�9)}�IK�.�$�ܒ��	nĈG�Ì�2��� �׽���t݊�$�ܒ��$���I-��F�Zp�e�16q���KR��mf��j�v_aԛ8��f����4V�հV�s} ��x ~��w��t�����$��`;�������}��es�MvM� w��ϖ�����H	��1T�k5{s}��m��������{st ���ju�!6\�����7�IH���%ȯI)$|�B��1v�7f9M�޽�=���u�I%$��J]�w�$���H�Wj��Uه��wn�o ��_} ��� ;׽���}9�	���
�WKg��ݸ�MnJa�͝v��jvF��2k�(iL�4�m�7���y��IEr+ĒR9)}�IEr+Ē]��齺]�jf�\���t���s�l|��=��}� ��}��'6�{�������Sx }���������x�Ǵ���B���$:[����J^�$�,,���~�?sDi�Z�I��5ts�	�tlY��͙��l�daJ�Iǌٻ��o]C\���V��������l_ٻ����j8Q��HZs����4������g�U��ad�BV�f�u�HCf�<�����Z��Z�H���;��S�ܪ����,��6����?���B�@�����HH�ќl��d��a$���na�����;���h|Q���;�s{�����x�R�e�!0H?�l 2S5!1���m�{٭���4}��t�C�l C �$XB�X��Ӧ�d8T�H��V��Sd��0���l]�l�5�S�����������C�
~b)��!ш����@X��#�$	 �0 Dڈ? =H*i���EB"~˿���m��ݹ�m���駬[�l���@:n�� 
I|�R�K�Iz������ޥ��$o�]�39��go ��_} ���I%#���$�W"�I%�I�Ɠ��J1�&^�V�7�NHj1�[�X�J�SY�&�B��¹���]HM�9}���M�޽�=���M�$�݀>��} ���ȹ�e��� �^��ȯI)$|�Q\���UWv���>��� �ʻ0������ ;���҇v�v� �^�z��e7�f+A�fݓx �z��v�v�;׽.�m������#h"YbР��H�S �Q�?s���f���g�]���kQ4�_} ��� =窪����z��w�+ĒKwo1	ow2�T�YY�K3��18�6��Q�x�i5��4qc�FEa3��Yt���&c/�`�u$���R�䒗r]�HJI�$�W%ߔ���zŻT"�0����W�$��?�I(�Ex�JG%/�I%�v�`�s�MvM� w���7zo ��a�7zo �ߦ��u!����7zo ��a�7zo ��_} �I���X�5َSx w�������� ����@����ݶ���|)�F��ba5�^M��y�i�-`�ˑ.�����v��Β�Kr�u��������P�Lf�"�]+����m�:H��[����띈�m`�n55%�A�jJ%�b�sM3cjD)ڪ�k���C�֋+���RTS@��wj^�4!��7�M{������x�v��T�G�$��Mu�D��B�n�gc�ڤ�M)�l�t���6A;��I$�䜾�i���"q���Ŧ6h��=l�e:^��Oa�ƒ���6�� Y�V�`���e����� ��}�ȯII2Q��%��c��Zuv�m^$�RH��$���I)&J>���M������3E���a��䒊�W�$��(�䒊�W�$��?} ���Ï���0p�� �^�|�Q\��$��G��%ȯI}6]i�3�����@:n�� 㜜��{�}�Iy_��IH���$��T�9(i�C�3T4�H�lP�]u�oc�ɵ�bG,Fزt ���wLRX~I$����IEr+ĒR9)z��W9���|o�7������n�5ʹ}�-�����
;U>w���s}'9m���M� w���NI9�)�;�8t�Sn�ر$����|�Z�Ex�II#����i��o�^���#�eq�}�Ij��I%$��Ke�,I%$�/��~;�M�FQ�fݓx ��Ke�,I%$�G�$���^$��rI;��~Ș����]P�Knf���G7])0��-�AMXQ�E	,�2��F�p���� w��O ��a��ޛ� �{��@?~��Vb��.E�$��(���.�E~�I$��y��Il�i��{ݭ�L�sr� f_} ��{sv�o{�뜿�����!�"�BRR��������
F#bBVY��f l ���[�z]�m��߉�[m��I�u���5�7�}6�}�Ͼ�w��,I%$�G�$�ʹo�W�$��Yt}k�R�\�����< >�O���Qޤ�W�+ĒJI�$���+�j,��J�	u�2[n���J�5Z�Cde��M.����'�㯭��C�i���%����G�$���^$�RH�ʪ�{i(����~%���`�n˱�}�Uȯ?W+�r��m��~����Iy_���$��|���$�9ͱӿJo5������I%�{��KUȯUUr����F���@���q4r�fa��}�I~��ٹ'��x��~�w��I:�#��0"�)����|s�f{� ��R�t�麷I��$�Q�{o����{� 7dx��;d�{iwX[�T�P	� �m擅u�b���ٝKVܣj��o�K�Zꄭ��"�����< ݑ��A�y���=���a�sn�gt�}�������=�ߞ������Iy��*��.���v� I�<H�z���{t�����祥���s��I� �^ I#���W))=�J�X}�B�]�r���}���>��o��k�I���ܓ��M�6�B	�9I��<�m����pvW�+��q����nʦ�`�]�\qř7�x�ۯDEp��d���f�2�X��8���G��� �:�2��h�.Rj�4�n��^�[t�z;*%ڭp�5 �^E��ٹ\�� cM�s5����n^^�e*nJ�WlQ���ɘ
���u��@\�3@�Z,�]d*6i؀lj�-��+���*t�I�y�|��M���6 ����)<�������Zj��@��Q���
˄�6�]�B�po�� 7dx��0�%���Yt�+�t[o 7dx��0�%��<��K�K�����[o �9F�$� �G��<�%�eէE�M�m%n��r��߽��{�x�#����^���`��Wx[E�ڶ��ݻ�	$x�����{�~� �^���M�m6LT�A�% ��ҹ��Q̷<n�/l�݀�� au�};��iz����U���|�dr��I~��{� '�z�L�خ�e�v�H�S�\+y���9¸rA$N���M�Sȑ#	$�We���
H�C 2C���
���N^sٹ$����$�}޾}9��?�}tA��T̾[�� $����8�'��{��`]ڽ���%f�)��Ns�>��-���� �9F������^%Oc�.�tR���E�x�#�?s���W����/߿^ I���/c:j�%I�c.�ۍ�����A��Bf;�q.��c���imr�5ﻠ�)q�:8��n�-���~� �^ I�����Oy��밼��$�ۦ�J�T���?UU]��������巽��_>�}��o�b����I=��[�O��u���"U`�%�"Q�"�A���ʯܪ�?߼�Q�j�?^ٮ�F��.���m�r��I�<ޏ�`RK��9�����m���o��0uSe�_(I�Q�z��~���zy�� �d�
l�\�����Ji���@�x�m��j�q��u�{o�t����F�W9-��n����z�M� 7d~�W>A�G�0[*�����&�V�[� �c�s�ĂOy��~� �^z��H����M���t]��{� �\�����¹����ٹ$�����$�߈W��fL�L�C��9/�{ߡ�<�}��{�u�4p�@�J�$������$��n�x�>����v�V��T���ʯ�\����ߟ@=�ߞ��������TK�h��"���d�m�2f*����4���i]�DS&KrI ����[��m[ڻw��<�vG�I�Q�W+��^�� �Gt]/1�ut���m��=\�s�I�~� ��z�����_>����o~'���Se���=��F�r,=UUʤ�zy��|�/��g���k��Vܒs�"����w$��������nO��A���������m��m�Fg!sz�G�~��U~�UU_�����_�R�;.E�0�w��$��)�(���(0�*�i���!�@�d�CbR�>H\�A1�)6	w�kP��o(G2�%e�.nB �R\�L2�t���V��Ƅ(_����4˩-`�FA�A��r�~>���c��~i$ ��	��V4!X�!ie��i@�$�l �V�BB Fd:L&�A�0�O�%�~��Ĥ�f�2RV�a
��c.�07��YziO̪F�74C?C2I84��$Ye	�T���YH��~	L%�h��h� �	ce-,)7��i���7�2D�5W�'R�]h��.��HB�B�B&+o8CZ��	)4s�A7�������4?����\J@4)w�,��N�Iau��.��ɪV\La�Мb���d�)�����Kv`V:�U��s]��t� 
�z��m�@/V'�;����dq;���R�����4������م��e(bo��0�T���rC�l5�8��Pr��AZ���gq8 �n�i��u�#��Tn���VҦضE���^��hsdƭl���؄�-方��3;jR�h���ʐ��fף���,C;JQH(J.��лk� ���f��ba�ZDm�-���)8�%4��·n�X�sZ� ���Ȋn|;.�'j��-����-��Fm�dZ�E8L�M`cQ�6�!	��@�Beu�[If�������#�Go�� UI���t�v�FKJbMK��A�KMk�� D$n�������x��Jȼ<P��!�ㄝj鎲��Ԃi��zR�Ku�8�hE����a&�7�kUmi	��ƼBKh�!s���.���+�I�(�n�Q�M/X��n�VYkyF�;[�FX����9�4��!�8[�#;���λ`l��c�����Kv�ڊ	Z��Jt��ŸeZ�鵀��K���4�UT��Wt15h���l-��R.��s`��Zsɛt����uԶvr���e�s� �,��J��6g�Ёٲ��$�aב����#���d���<ρz���^��u%�R� �,33�5�m��[cn�F&�J�&N����q���Q�J�Zs���P,�	e�h88�l)`�����lQŲ��VԨM�)*̻<`b�p�Oc
97h7���!�]�qƵ��v��J��ݲ����+m٣q�lڀT�U嵍�!*t�n�9����!���a�R�U[H{)x-�R.����V����%��R`�j����B] ������9Ø�Px�=M�P�6@�N���~P����m�+�n�p��U����!���͗S�ĸDe�Kq���:�-��<��c��<;��okt�=,��1�.�8iā���M
]Izۈ�QS��5u������ ���� ?)D��+���C��*����	�C�gob��Jpɝ�e�N{P�(W b�燚��tM�Zt{<X2�N�rb]ݞ��"��u��R�]vv4Ȝ{{�+s��Μ�tt����{�Kە��:�L:k<�vFk��g	��k�v�Nz���؇qع��oh�Z����Z�nک�f�mǠ�l9w',Ä]�koh-t9�n;���G����C�3۪���\�����'������H�gl3<�I�6�b7i�Hs�<���U���CY�YWQ�P�i�&/�N���m�[�4m�� z{��$���ˑz��W�zy�}�%�ӱ�f�f�W�{���{�'�I9vO����߽���=U��F�޻�V�m+m'n���y`����'96>���~���/@�{��ۘ�"����X��q/zy����$�(��99/�?}z�{P��t��*����Us��L���y`��?v��l�m�qC,�3�73���ɳ%����Ɩ2+uu��p}$���k�j������G�0ˑ`��W9���'��߿= �������k��V�~�w�x��A �-dV�) A�@��BB��+m DB"!b��P�u'��kp�y�k�g�W��+�dS�w��C�V�B����~x�#��ʮ%�\�^����@��卾̴6�2���o{�krO{��7$���n��T�3?~��Oޢ�?VS��lv$[o �\� �s����������)n�v;�3Tf�#�x���d0�3VJ�,H5���&�L:0�h���O<�ڇ�Ɇ��jM����� I����UUW��Us������z����ݹ]��T�f�M�=U�U${� ���Xeȳ�\�RFȘZ<���E�mݷ�{� ���K��N ����oٹ$������}�U�3�v\��~䓜��9ʫ���~� ���׀lx�W*�Ws޴����hF�+�����s�\�&����x��[[.Z-�a$�z����ȉp�cv�zNN��֕�V0��i�N�0�&�h1�"V��zy�� �\��\���5Oz�J��^��*��e��m�vG��*�I�~� �=��	6<�9UT�=(�^�`:�ӱ"�x�s԰�%��r�#ޞx'����m�ε̽�N~��z���t��~z}�{�Ɂ��~��Dq�A�i^�~PO��������w���L��k[Y�Tn������?Ns�����}���߯ߩ`RK�;�dƓ�Ƌ����>�����"�rx����h4a�*���@ە��rI8��viz�Zg+�� {��=�oe,�I~�r�_ '�� O*^�'HX�۲�/@�����9'?s��&Ƿ��׀��� 7dy�r�\H$<���)��m�v�`��^ l���+��H��x���un�w8��V�ջbV�ܪ�R^�� $��v��Ur�m�޼eEM/U�5V��l��vG�~��?W*���~/�{����	�T�s���;�{�@��A�e�jf�h�uz�x����Gc3�=�+Ը�� �b���v�م�щv�Os].ޜ��a��g�K�z��lՍ\�g_�3�<�������l�ҭ:��n6�Wf�dM�gs(\ڨ���-!,&� 84T��KaHɊmi,]�CiG��v��m���19���RQ�)���ey\Y�vU(l�J�]�j����q�#˜�6�@ӻ���ܾY��� y�,x��Cq9Q�YX���̆�X��r��2�A��9${�/;:�͚դ[o@����x�Ȱwc�UW>@y��=Ͼ��k�fع�X��E�� vH���/=\�RF�z՘[n�U��)�� {g� vH��*�����X��,����qt�m�շ���U%���=s԰���=U\Jzy��=I�bWm۶������Us��������~����G�yO�}�5]b��2�B�;9
�ٵ�Նf	`R.�"B3��n��N�/�y]eb5wm�n�/������< ���U�z[߷�C�o㽻o�]��3���O���{E��� �R�׽��=�{�ܓ�����/�d���j��0�2�v4��Oߞ�䥇��T���^ O{� ٴR���t���"�x�UR�~�,T�� 6H�=\�q-���;�y^
��:��7m$���:���$x�#�6\���e��݈v����\�t��#�� ���`�jՇe��.:6���t�x���B�(9=��߽��<K����Uϐj��x�&�#-2�U��{�ߧ$�->�{԰^�� $�竜�r�	�KާiV[[M�9z�|��������94��HH$@(@$H���?�v��D�<�����$��{[ ��{o�H1m�+a�������=��	=���U�r����0^��}��c,�Ks�����$䥳����V�x������t�q��۫�M"����YƤ-t̤�Z Tn��[m)nk�51:)Y�}�ݞ��;#�`[%��UW>@I�<}!/>���+MU��}}�~��KMS޼ ��xݑ��W?r�\�7߿��,v1SM�&��"��׀�<=\�RF�y��?Q�wv]�am��WV���n�=�URR{� 6{� �Q���^����߳rO{�RfOj�MZm�M� �����V�x��@��Nr_�=��0`�qK�n�cfn�F�e�;K����0X�⤱�(33F��N;�,���N���?~��;�"���\�����	����C�ҵv�7n��r,�s��I�< ��<������s����Mw�lSfr
��{�����[�?Q�l�ye�����t�$�Y�r�[�$����o��F�r, ݑ����Ҧ
�am��9F��V����	=��<9|�QG
������	�� ��K6��[�V�HS
�La���ə� 0����	BSX�)�J�S;�2oH��g���!4�Tqm�-���U�7E��f�D�r4ml��G2��8�.b1�:)J��yRPŔ���`f�!�;^ZJ��^ݝt�X����r+]`��s[8@����c���I��gB
&���7gځ�&���Ƥ�.�+-�
/��N�<kﭵ
�f!L��ggiǷT簥�5�^���ݝ:	�AF�q�=���^
��;���tt޹�`� ;�?W9_ �y��d���m��J�v�k 7dy�UU$=�o��Fݹ&�W�:V[j�m�vG�vG(���U%�{׀{� 6*[�iY��*��}�I���w�t/�z�vG���Ur�Us��������/�@:��E�Iۣ ��/ �+��['��=�}��0����V[mP��[���o]�."�V��{k�0I��/2��ź�95ήm֬�Ks�����nǀ}��?��s��W���'�*~�Uv�mf/@<��^���9'=�N��Ԅh�� 7Gf:�hD
�14�t�&���P��`&�*	 ��v�C�����`�=x���ܪ�URF� ��*t+�������`)%���Ur��9\�9˲{ߞ {����ʼݪN��m�i�0�������ǁ���$��~�����m:j�Ɨa�]�ݏ �W9��)'��vy���$�-��~gyWZ:����J���	e�0�ئe��256��a]�4��>�Nw7���:V[jڶ� �y�lr��$���I�'���~z��>߫���v\���9F�^ wv< ����UW��'6�?[�h�m��t/���ܒ~���sD��@:"H��#D�IEc,�M�1M��24y��{�쌉tL���!����䔰$�hJHA�%����~�ĳtC?D�C���a�>��~l�n�jg�1	@�$	2�#���m%5i��h%��c	?��s2!JF#ā"��V�a$� Aʤ+
0� �(��	��a!���0��2kI�i��HA���G:O�%�#B��Q�l�m�Ja��0�~I��!�����7j�3�N�8��J5,#B���SD�� �����n)c��\D�#���`H��`L���~�!�14ɶ��i)m��1,�ł�ƱHe����(��Ě(XA#�ϑF�أ�j"|�6ʧ�t~ �:'�4���/bT��PJ��
�4��9�r�|�� �����Z�[�����lJ��{��U%�y��� �nJX�Ix��NYWulN�ۦ���wc�=\�s��Ծ����[������hh蔕�[E�Kv���������N�)�ҭ,t,�I�2�|�ѕ]5vm�e�԰������ʮ~������~z���.���NX�4��������ǀ}�%,�s�I����Zm��eݻ�������U_��s�{�������׀M����X�J��M�o��+���� ��^I9{��������E������'���tCeʾ[}?w�ym������޿�6O< ݑ��������el'<��dD�y� l���$�	P}�qЕ�XC<���Hu�oF���U�7W�"����wc��������S�5H]ߓv۰n���x���vG�I)�RK�r�������U貺U�6^�{��= ���c��9%Z��^ I<���%c��%nՁm���W�s������`����wc����LWv�X�@�0mрv\� �ʯ��/����{��}#�`������m�:}!�Ղ4�fCN��r���˥vFj�� C��S��[.�3ru�@Ж���Fd�%�4��{2W1ĝ �q�d��K��5Ž�;e+��=x�)7~�m`~��wm[�U$W�;�c�;�8YҁF"V�&�8�	U�:2����QoB�ts4��40Sq�e6�l�A�N8ɕ�7@�9鷯t���QKnӤ��ΒN�>)�,�[+1�LX�-���	͖6���9�)�=�t�QXSۏ�{�_|�}�����Q�o�����Q�v\� �U:�\C.�]��V� n���UĎ���`��� n�y��) �P�ZnںwM����x}��0ˑa���9���]���< ��~xV�%�um1���t`�"�ݏ 7dx��}�����n�un�+k 7v<����y����XzE/m�j���rUŻvS�&��H;�
��,��8�l̅��u�1f[�2]�X�e� ��y�H�eȿW9�I�o�P��c��l�o �G(˯�VWr�P��,�PWJu?�7�{�7�܆�� 7dx{)2���[\T�0mрv\� ��=\�H��x}��0͗wX[n�ա]��k��r�L��$������Wc�`EN�Z�2�Rm�����Q�v\� ��=������ٹ���MZ6(	�p��qB�G�
�-���h�M�hb�s���]��N��m۶����eȰ[��\��'����kɪ)մ�ۧmрv\� ջ/ 7dx�9Fz��H�*]��n��;�v�[X$�����nkC���(�0��!#P����z��׉�'޹�vh�cV]7J�t�o 7dx�9F�r,W+�I<��J��:T��-��}#�`�s���/�$�x�#�%.�˶*n���a�`�f�[�e+���r��@A��+�j�����iX��*v�6��;.E�� n��Us�s���o������wX]&4��۱��wc�Us�H$���y����X��իPj�	6۵m�� �G(�ܮW)-��� $�x�i��g�f�s����r_��w�t��� 7v<J��*�
7��W����R�T�Ս�ۧmрv\� �*�ʗ'��	=�}#�`ml�"anE)�[c]v5FȚ�"��7t�kcn��-��ֺ��7��vZ����v�[_�� ݑ�H��UU_P���נy���zݑ��\�6o@;�<�+��ܪ��}��� ��ߖݽ�?T���&ǿ������X���Z�@����v�Xv�, ����i;V���q�[�����W��,e�, ���?W9�������X��]�at��	]�cm`�ذ��)l���v_�K �����6����H�D���bTE  ���S箰���R�w-�eŎ������s{vwn4.��(�m�����S���\�8��v�nk�;m�5/o<j74�ƭ�p���c2ā[�@m��]�84�V�+4�t�i釴VC�8�uu���a�C\hp�x��D�m�hl/T�����VMB�J�[,�螅Y'r�.<���hU<%X��u�"b�u�Mcr�,ֵr�.�:���97&�	rA�kIT�1,���p���nc[�ɮɰ�R6�jA������mz�qj�u��{��>ے�ݹջ/ 7����K��r�/��n�}$�z��j�׀�<�9T����G�T�մ�m�mрo��XV� ݑ�lr��v�[�cl����m`z�T�������>��ʮs���U\��?~X��+�i���cC���#�>��v�Xv�,�Y#�V�۞L�Z&�u���`U�9(�<�]]-�Kz�pă��&�mI��%L������0�Ȱ��_���r�Us��'�~x���ZV��e;�|�0�ȱ(�� &�3���rIϻ�nIϳ�.�\H�=wu��l�V��M�x˞X�G����z����$,6��;N��J���))�y���R�5O}���_7������v�)4ڹm�x�rR�?s��+��{������z�m��:Swer�h0��(u<����9.#���]��NIq\@W<h��w���7�T��I�Nۥ�^�� �ݗ�H��䥀un����ۻn�;t���[����U$���;/ޥ�j�^{���}���k1qsQ3�����ϒN}��w4��G�#,d H%�Ĉ B(�0"0H��(��
H��6�/1_�x��,v��ذN���j�m�~�W9K��԰��^ݽ� 6H��i&���q��[����j�^�W9\������>ے� n�l��{D@7D�h�jP�e�ʫY5٤�;�q�6�\!�X�-K��;��̠O)���l-6���=x�c�>ے��l�B���C��l�v� 6ly��\�~�9�W.�/��W�y~���5M���uq���e��v�m�T�W�j�/��~�*�\��/��x�����R�)��[Lm�ݺ�UW*��/�׀E��������| E �,u���3`uwn�wlmݷJ��Wn�Se����s��+�W���>���ߪ����;�1*�-[n��р	�*�PK���a�6�=/��s��-�\ؐ!������ջ�	6<K�K �l�W9��9�/O^*T��W��N���P�x����%����nI���7$�w����M�I���)��M]�X^�� ��,?W+��$O{� ��z���w|�)��v+�;n�	/b�:���I{)`}$�%�{�۠y��>���\��7 �^%쥀j�/ ��, �s�MS���fҰ��#%�Kl��Oī6q������a�`}B�BB"BB@�	xkP���%��2�I%)%w���h��dl�9!I����R P�����6���6e]�����sFX?���Ą�"�~IXXBP��NƇ��a I!���Bda!$!�z�kS�*�BBHB$Y�� ���$ϳ1��"��
B�9
a�76[�:c���=ޚ쪠.�l��G����=��g���M�S����]��m��]���JJ���@���:�-�Z�tIV�/	����a�1�C[�ĵ��E�8�v,�0�(䷁�zb�6y�P���m�8�Pp5�mf��h!Q�����l��n(�Du���&�����9��u��Kli犀�gKvp��]��>#��I*�������bL�[V���ny��闦��-���(
��U�V���b`ke�3R�6�n��s�����)ͣ#�S]mH�݀�U� _m4yt2��6	��Љ[,ƃr˦)1Al�3v2R���ys{@�hZv��uq�t��ժ��v��<v;#p��y�"��8��=k�n@HZ��M��tW�m`Cp���l�唺7�4m�8���8�KiNvG&[u��	��!G0�vq�@�����ƍ����crN�P�Hp�����Vb��ؐ
P*d1�.���sV�\!�A&`���Silv��!��5�$,:b֢��`e�(���2��}qN�Ia�S����t����B�1�L�,*���mp��h�c�v�`��9kc��rv��YS�ۗ�ֹ1��Q�S�VJ��׬.�
�X@�.1�7&�0I�qd��r{a�:��
�Y�0@IL(͚���Q�>�-mW
 �6�;r'C��//mA�]n�2�G�v��r�b�`������Ԗ+c�j
�6䕥�#�Y�\B@θmQ��4�MF���FY ^����LcS� =�z��/!�[-S�5ڑsɵ�c�4:e��q[;���kp�B;��P�U]��.�Fv���)�.�B�<����)�˪��[[Ũ��Ciy�6P�j�����P8����9�f�íT�Y�i�Lr�h0Y5�h�n֒�]t@-�K�|h1�)J����ƸlQjF�7X[r+ ���ڄ�8!/��P#IR=\�T.l�� 0��eXiMu�Yv%��jK(l ���P��E@��A1 ����u ���!ǂ�mU:� > D�O�E��G`�g9,g������3;�*R⫉E����+qk`���F:��cc�*t���"h�3P٬�V��gL�B�	�E,�ԥҶـ�-d�H���1�&N�2��y[���fS4�ݪ�9�Y�f4��s��h�ˊ� �����'���ΌH�]lҋ76PX"i�n�F뙍4�vV I�[��ö���ٜ�Mmt��/Z�-i���Ν,{���=ǺQLj�쥍%��MY��Pm@3E��a�M	tW;7n+
fXm����� m��n۷z��԰[%����N~�N�{�~�z����m�L�U�n��d�eȰˑ`.JY��O�s�c�����V�Yc�nw@�����ˑ`.JX����IK�$f��ƵwC�rN_>~��~�}/@�$�Us�R��^*T^Ww�T:*�m`/`�RK�6\� �r/-����F�\.�j�ebh(�:�l�Ψ�C�v9��R�y�(B�$���w�fR������%9)�NO~~��r%�bX�����I�&D�,Ok���9ı,N��٘re֮d�-���kY��Kı;�{�i�lZ�� t����k޻ND�,K�k��iȖ%�bw=�f���^B���׾C}]�uEl2�rr%�bX�����Kı;�w��9���w�ͧ"X�%��k޾t��צ�5��}��*dA��Kı;�w��9ı,N�}��r%�bX�����K�K�?|y���/!y����� 6�G+�֥�r%�bX���ٴ�KİW�׽v��bX�'��}v��bX�'s��ͧ"X�%��k���52f]\�K6���VY�b�S���45%���Y�-��c��2(��a�	�OoMzkŉ�k޻ND�,K�k��ND�,K���f�� ~��,K�����{y�^B�}����������D�,K��}v���"�"dK����ND�,K�����r%�bX�����T�,K�N�ffre&��5�ۚ�ND�,K���fӑ,K��{�ͧ"X�)�Bj(PRV��vj'"k��.ӑ,K���]�"X�%��y2O:�jf�u�L�r%�b���}�ND�,K�׽v��bX�'}���9İ?��=��L�r%�bX�{�٘reӂ��*y���^��ק���o:{x�,K;�w�iȖ%�bw=�L�r%�bX�Ͻ��r%�bX���Դδl�pMXF[SK�
da�̭�&�5!�[bi��b����Kd��l�8h��"X�%����]�"X�%���}3iȖ%�bw>��j�bX�'}��y���^��ק���/�����r%�bX��{�6��6%�bw>��iȖ%�bw��ӑ,K��}�ۼ��%9)�NO>O�>LTlZ��kZ�iȖ%�bw>��iȖ%�bw��ӑ,ı>�wٴ�Kĳ��?}O9=���/!y?�?m�ʸ*��[�ͧ"X�*�2'�����Kı;���ͧ"X�%��kޗiȖ%��*p]|�J2���e����!HB�	B���V@*`�D�XVVI#'���(�AĀ2 Q?�O���G�v'u��ٴ�Kı>�m����Md���eֵv��bX�'���6��bX�'}�z]�"X�%����ͧ"X�%��k��ND�,K��]����jk���M�`�/�r�����K����f4`�!g�К9 ���X.��<��Kı;�{��9ı,N���m9ı,N�]��r%�bX�g���p�%9)���{)�"L�����Ȗ%�bw>��i�-�bX�����Kı>����Kı;�w����^B�����m=�SkK�7eͧ"X�%��k��ND�,K�k��ND�Bı;�w��r%�bX���}����������O-��;l�a�]�"X�%����]�"X�%��k�.ӑ,K��}�fӑ,Klg����Ξޚ�צ�?��~@@%h浭kY��Kı;�w��r%�bX�Ͻ��r%�bX�����Kı>�wٴ�Kı �*?I��*56�x]u���FXb�1�0�2b\�kP�lìC77l�t�C�V^.�ڍ�vDac,a*m@���b��jI���m��\@v�.�1v�1f!o+�,��@��J��4��[�Q���km�q�J���6�P�ݷ��d^gY$l����]�̱�H;5��a�b�zZ�!Rs�[q��ػ;Z�{>���s���$��'t=<�hb㣳�.ٶy�.뭐]��^��Whr�;m�#K*ٴ�*���.W(��t��X�%�����r%�bX�����Kı>�wٰ�R(�dK�����/y?�JrS���z��~�(�̹q��ӑ,K���]�"X�%��{�ͧ"X�%��k�.ӑ,K����6�����L��,O{�[��nj�Y355��ֳiȖ%�bw?���ND�,K��|]�"X�b؝���n	"��jH$�����30�&\�n	 ��w��Kı;��ͧ"X�%���}�ND�,K��}�ND�,K�R[��CP�L�5���9ı,N��siȖ%�`=�wٴ�Kı>�wٴ�Kı;�w��'�����/!��������uj��uB��I�C�Iy��hp�sH��Wx@"e\�乚�Y��"X�%��k��ND�,K��}�ND�,K��|]�Ȗ%�bw�{�ND�,K�v�L�����Ժ�K����Kı>�{ٴ�<h H'D�@���Cm�Ȗ'��p�ND�,K���6��bX�'}���9�&DȖ'���?���\	����O㒜��'ߟߋ�O�ı,N�}��r%�bX�����Kı>�{ٴ�Kı>�_kW%�Ū�ʗ���%9)����'�߿n��Kı=��]�"X�%��{�ͧ"X�%��kޗiȖ%�b}�x���j[�e���'�����/'~{��r%�bX/��{6��bX�'}�z]�"X�%��｛ND�,K�N߿�j�!M�Jdt�C-VO6x?M|v��I��1��ӗD1g���0W7N���f��O�,K������ӑ,K���iȖ%�b{;�f��Kı;��iȖ%�b}ӷٙ��$�55�2˭]�"X�%��k�.Ӑ�JG"dK�=���ND�,K�����r%�bX����O�`dL�bw�)-�/��2f̽��9)�NJr~�~��Ñ,K��{�ͧ"X��W���$�BH1�B�2%#Ē&�H�Hd!#F�A�d"2@`BԞЊt��O�s_]�"X�%�����9:k�^���}��{�d$<��K�,N���r%�bX����Kı;�w��r%�`"̉���~���9)�NJr{���k����,ٚͧ"X�%���޻ND�,K��iȖ%�b{;�fӑ,K���]�"X�%�����xәe˭CX�m�e���*�#5]��5H��,�i�R�M)�6�AɌ���9Wy���^���;�w��r%�bX�Ͻ��r%�bX����yı,Ow]��r%�g%9<�?_�q��AZܲ����%�b{>��iȖ%�bw��ӑ,K��u�]�"X�%��k�.ӑ[9�^O�����-Ks�3����,K��}v��bX�'����9ı,N�]�v��bX�'��{6��o!y����m�36��T���bX���뾻ND�,K��|]�"X�%����ͧ"X�4+�b� HX�H�b�R@(| & D��D׹�kiȖ%�c?�:}���J��3@��'�����*w��Kİ�B+�w��6��X�%�}���m9ı,O����9�B���~����͵��N;�@�b�Yif���#���a1s�4��n�H����0�L�5���9ı,N���m9ı,K�w��r%�bX�{]�ؼ�bX�'}���ND�,K�{��,�uus)�5�f��ND�,K������bX�'��}v��bX�'}���ND�,K����ND��"X����5�Wmr\�/y?�JrS����~�v��bX�'}�z]�"X�%����ͧ"X�%�{��[ND�,K�{�`�K�j������Md�z~����9ı,Og��m9ı,K�w��r%�` ȟ�߿�ӑ,K9)������v�H�[�^���,Og��m9ı,?�)�{�6��X�%���{��9ı,N�]��r%�bX����HR`�X�D � A��"E��:��,���O�K�?@n��c.3��-�˙�g��[��M8���6�Ͷ[[̠��D�� [e��1̸̫���,Es�8�[��m�-s���E�ɬl�FQ�{;�*�"t`tu��ݺ��6��ѭ^�J�'��
KIn�-��Jmͯq(�DͻKP��$��a�R+��K��G�lC\'�L�C���^���0c(�[v�Te��NNN����t�on����.3.l�e�8պ��p��XGk���9�P�i��ڔ��m�3Y.k>Nı,K����m9ı,Ow]��r%�bX����yı,Og��m9ı,N��e��h� A*)�OoMzk�^�~��o:{�R9"X��׿�ӑ,K����fӑ,K��{�ͧ �%�b}�����VU+1L�r{y�^B�w��ӑ,K��}�fӑ,K��{�ͧ"X�%����]�"X�%��N�۶�CP֌Ѭ���r%�bX�Ͻ��r%�bX���ٴ�Kı>����Kű=�{ٴ�Kı?w�m�}�[���l��Oo!y�^Og{��r%�bX�{]��r%�bX�Ͻ��r%�bX�Ͻ��r%�bX���O��٩j�kJYr$M��A�f7@�f���a�f8�3`����}��d~`��E5���r%�bX�{]��r%�bX�Ͻ��r%�bX�Ͻ��r%�bX���ٴ�Kı?g������[I��f�Z֮ӑ,K��}�fӐ���C��P�� �_�2%�����ӑ,K����iȖ%�b{���?�O�漘�'����ɵ�G8�]�fӑ,K����fӑ,K��w�ͧ"X�%��뾻ND�,K���o9=���/!y?������l�f�iȖ%�b{;�fӑ,K��u�]�"X�%����ͧ"X��L����fӑ,K������rLѬ3�Mf��ND�,K��}v��bX���]��ͧ�%�bg��iȖ%�b{;�fӑ,K��~�ܾ�U����4!��it'l]mʈ��M^-ut7/SgH])���*�;]�.L5�~�bX�%�������bX�'��{6��bX�'���l?�'�ı?�����Kı;�Զ�Ě���D��kiȖ%�b{;�fӑ,K��u�]�"X�%��뾻ND�,K��{[ND�,K����,况2Y�kFf��ND�,K��}v��bX�'���m9Ƌ�>����eЦ#��ЕbЅ�\$ 0`���ӫ��$���,�CѲ�
O��8JLˌ0��HC���b�L�H�NJ�r`JD0�%�d+��mM�۔�%%eae%�7�U��f���$�i�J`jK(�Ȁ� �`�n���.C��8@'�iִ���. D[��hɬ�4Ќ#)
���i
k�%Ѥ�5�0���ISl+�	���Fl~����b�1!MW3N���j\�$�.q7M�Rf6ĉ
$d� �K.�v^fYY��B��	L�a&­[���	a���.�	IJ�A�FF��^�7N,���c��$��%��CKR���#(K�	���T�IHPÛM���n�� BH�2Ʋ��)ckZ���ܐ��nI�i
YIYi��$2��T�L\k�F$V�ް�����t�J���]G	��`����F2�PpQ��TM/�~I�Q>~z�<�	�z�hR�D�%���[ND�,K���6��bX�'{�䙗٪]a5��]f�ӑ,K?� dO�{�ٴ�Kı/�����Kı=�{ٴ�Kı=�w�iȖ%�b~�{3=Bv�� ��OoMzk�^����>qȖ%�b{>��iȖ%�b{��ӑ,K��u�]�"X�%�����8��]ta��J�Q�6w��[��9zDK(b��7\A6+����k[ND�,K����ND�,K��}v��bX�'����9ı,K���'�����/'���~َ�a���ͧ"X�%��뾻NC�A�DȖ'�����Kı/�}���"X�%����ͧ"X�%����}�e��0�d�֮ӑ,K��u�]�"X�%�}�}��"X�%����ͧ"X�%���]�"X�%��N�fg4e&���ɖ��m9ı,Og��m9ı,Og��m9ı,O}���9İ>�D ��O�)�LU��{Z��iȖ%�b~��e�������F�ֳiȖ%�b{;�fӑ,K����ӑ,K��w�ͧ"X�%����ͧ"X�%��&w����4L�	F$Ӭr��/Y�h�.�:�CPcgq���lBL1�2��!4v˴A`)�O�ŉbX��׿�ӑ,K��w�ͧ"X�%����ͧ"X�%����ͧ#�^B�w�|�l6�ΰry���bX�'���m9ı,Og��m9ı,Og��m9ı,O}���9�s�kɎJry�~�~�L��"�esiȖ%�bg}��ND�,K����ND�,K�k��ND�,K���󧷦�5�O���>���F ̎m9ĳ��]��ͧ"X�%���{��9ı,Og{��r%�`3OϿ~���9)�NJry��?l�f[V\�d���r%�bX��]��r%�bX���ٴ�Kı=�wٴ�Kı=�{ٴ�Kı>LS���8P��K!d� A�P�4GL\H!	e�u ���E.%��j�u->�&q�u��V�:Q�5�]cS�q'�5r�6b�kb�<�w�z�[�!ۨᘈG�'8]�;v�6<�g��	�sN�'Q�����q��.x3��m<t!�L�mauzU83W�ڊ)���vw]��<�^P8x�m��[j����.z[���wQZFc:�#��wuθ�n)���F�mD8t]�"Vll��Ga6$�NHs�p�>�J��ql�8r����+	b[JSD���mGt�e�Z��[��	���n�^g֯�ؖ%�bw>�iȖ%�b{>�iȖ%�b{;�f��'�ı?��]�"X�%��zR\��Rf�Y$�k6��bX�'���6��bX�'���m9ı,O}���9ı,Og}��r'�eL�bwǭ�M���֍W5��"X�%�����ͧ"X�%���]�"X�C"dO����iȖ%�b_���[ND�,K���d(��t�w���B�r���~<ND�,K���6��bX�%������bX�'��{6��bX�'~��6>�E� ����^B������ND�,K���[ND�,K����ND�,K�k��ND�,K�'��UM)T���l%��Ί])�r%�6�n�	瞤�]`�v�9Beay�Z�jͧ"X�%�}�}��"X�%����ͧ"X�%���]��?DȖ%�����m9ı,O�?���ٗZ�SFfj�f���Kı=�{ٴ�1 z�F>l�AX��m+J1 ]̒3	(�fJB�Z�DJ����%��k�]�"X�%����ͧ"X�%�}�}��"Y�^���?m����0%�y���D�,O}���9ı,Og}��r%�bX��w��r%�bX���ٴ�Ky�^O��_���ct�u<���,���?�����r%�bX�����ӑ,K��w�ͧ"X�%���]�"X�%��{+=����3Y��f��ND�,K���[ND�,K�H�k��ٴ�ı,O����iȖ%�b{;�fӑ,K��={�D���2��ʦX���]��Q4j7,��	6��]	E�.bK�1BJMiCD(�X��{��rS�������ͧ"X�%���]�"X�%���}�ND�,K���[ND�,K�~>�аPnD�S;�Oo!y�T���ӑ,K��w�ͧ"X�%�}�}��"X�%����ͧ"X�%����&�d���ry���/!y
���ٴ�Kı=�wٴ�K��E":(ḛ�����ND�,K�뾻ND�,K�z�3�Xf�e.����ֵ�ND�,K��}�ND�,K����ND�,K�k��ND�,���^��ͧ"X�%��g�����u�e4ff���m9ı,Og}��r%�bX�����v��X�%�����ͧ"X�%����ͧ"X�%��{~����
��R&�}�\['|�G�q�U�;d�O<p�d�A���-�մ�K���3Y��ı,O����iȖ%�b{;�fӑ,K��}�fӑ,K��w�ͧ"X�%������2�a�.�ֵv��bX�'���m9ı,Og��m9ı,Og}��r%�bX��]��r'�*dK������ZL�3Z̓5��r%�bX���fӑ,K��w�ͧ"X�%���]�"X�%��｛ND�,KY6zK5$�Mnk6��bX�'���m9ı,O}���9ı,Og}��r%�`A�|�J���%�%!P��$ҪZ嶒�V[m$���Ke(P�d���D�؟�%������9)�NJr~�����ek�f�й��r%�bX����ӑ,K��w�ͧ"X�%����ͧ"X�%����ͧ"X�%������p���\�kNea-��n��F�Nw"#��4-!
�Zm��uL�2AM�ޟ���5�O��{��9ı,Og��m9ı,Og��m9ı,O}�siȖ%�b~Ϸ�~MT�f���Ξޚ�צ�7�ﵴ�Kı;�{ٴ�Kı=�}ͧ"X�%��뾻ND���H�����,̄�-�.i7�O����ؒ	"w���n	"D�u�]�"X�%�}�}��"X�%��t�f��ՖkF\ԗ5�ND�,K�w��r%�bX����Kı/�ﵴ�Kı=�{ٴ�Kı=��}��\ѩ�f]���"X�%���޻ND�,K���[ND�,K��{6��bX�'�ﹴ�Kı6 >�'��f��
g�&�qX�NK��i� �h	4Ĳ�XX:�^�;�����gp���8����l"[�զ
�PB�����n2��m[a[�Ȥ���U��[l�y-Q�I��Vs-(��j�b�m�� �ً�>�d����Zs5��	Y�sn��1+gXsȇ<���y�ug�`U�v54JM�[vK%ФUZ!mmf�m#��N���Y�O6�k6�e�V���ع��u�,�kEY�m�BP5f3]
E�X�6��:��ܞ��%9/��kiȖ%�b{;�fӑ,K����ӑ,K��w�ͧ"X�%���K�o�D�5W���%9)�N��ٴ�Kı=�w�iȖ%�b_��kiȖ%�b_}�kiȟ�S"Y�����BʸM�M��O㒜��?��]�"X�%�}�{[ND���Dȗ�����r%�bX������r%�c)����6�Tes{��rS�����3�����r%�bX������r%�bX���ٴ�Kı=��i��^��ק���/Ɇ���8E�,Kľ���ӑ,K��w�ͧ"X�%��뾻ND�,K������5�Mz~|�}�РJ%+1s6�K	���Mk��5�3��v�:���v9�t�mTƹ^���%9<�����Kı=��iȖ%�b^���ӑ,Kľ���ӑ,K��ڽ�ٛj¬�@��'�����/'۽�m9"t@~GI�q,K�~���"X�%�}�kiȖ%�b~�����Mzk����o�qp��ΞԱ,K������bX�%������c�$2&D��_��iȖ%�bg���ND�,K�v��s�!I���35��"X�%�}����"X�%�����ӑ,K��w�ͧ"X�%�{�����^B���gB��R6�,�u��"X�%�����ӑ,K��w�ͧ"X�%����6��bX�%������^B�������(�� �h�!%.R���:܆��^�l�U$��UсL�b�<��������;�fӑ,K��{�ND�,K��{[ND�,K���]�"X�%������F�M����r{y�^B�w���"X�%�}����"X�%�����ӑ,K��w�ͧ"X�%������і戈3Ξޚ�צ�/�����Kı?{^��r%��C�HČ	2�a��L��FBH�
R,6�ƀ�tl�H�>�������ND�,K�{��ӓ��5�O������)L6���ؖ%��2'�����ND�,K�=���r%�bX��}�iȖ%�b{>���Oo!y�^O�ǿS3mXU�gj�9ı,Og{��r%�bX��}�iȖ%�b{>��iȖ%�b~������^B������X���`@��v�d{qW/6v�;=�+�x�NՕ,�ڞƞ��-)	�8O:{zk�^������"X�%����ͧ"X�%�����ӑ,K��w�ͧ"X�%��{�4%fX8�<����������ͧ!�	��,Og��iȖ%�bg���ND�,K�w�6�����y1�NO~��{I� �L�����ı,Og��iȖ%�b{;�fӑ,ı>�}�iȖ%�b_}�ki��^B���~���tȗ@��,K��}�fӑ,K�����"X�%�}�}��"X��H�Q�B0e�1��BxTMǑ=�߳iȖ%�b{=ۅ����R浘k3Y��Kı=���ӑ,Kľ���ӑ,K��}�fӑ,K��w�ͧ"X�%����,��Վa6H��-i09�0��*,kj�,�,�.K���ZM�����m�2�3Ξޚ��,K��m9ı,Og��m9ı,Og{���%�bX��}�iȖ%�5��>���&\�)�U_:{zk�D�=�{ٴ�Kı=��iȖ%�b{���"X�%�}����"��%9=���s6�E��l���K��w�ͧ"X�%����6��bX�%������bX�'��{6��gMzk����o�qE�!0�	�OoMRı=���ӑ,Kľ���ӑ,K��}�fӑ,K,Og{��r!y�^O����f�����Ooı/�����Kı=�{ٴ�Kı=��iȖ%�b}���ӑ,K�٧��(��#U���*m?l���.̈́/p&P�Ҧ��~�*lJ6h���ԡ�u�	�	p�`�I�h�v�f��S���4��A��55�@�%��dN~�&�U�$c�G�12�rd?/,9��l�T��6!X @�+��yu�2��1��	�)���Dk(J˻q��3�"�q��&B3sH�(�u��p%�B�$�c3��;s}ڜ#�\"�\�IX"D���H��Q��\C��`� �����C�%� 4�f�y��Y9�?I�s�d:��"CF���a�:r�˚g3f�s[&7sL6ow4r:�9��ޜ�%�`mS?~�B�5�$$��91��%$�$�G���@"�F�	�".�N�p���%��Z��M,��a2\�i�2��9���X�"2�#>�&�A���Fi4��&.	-��p���%1��3	��yU��>�D�-�k�*h�΁�y2PH�ry������(��Q]1{{�Kp�L���UƐT�m��됧�Vr`_�^h�&ȭ���\�RkZ<AM-��B��R�mc�`��՚ؘ�*1��(�#�E��Q���#��4�S����&�=v����93�ݸ:�`x�8_c�������	N%���$5+vr���a��=�Np'Z��[��D{�PI�.�M���0�r��SDŢi�k;h�9����*�f��lybܳZK�T=q�)�����j�\�uB��9A�Wla��Q:ےp�`+�֝'2dt*�ƭ�"x��֓	sm�{�2t[<h�6Z�J6;[a���]��z�p��[P����2� �޵��mrlt�����k	�[�t>��0&�׌��z�N�Mԕ.R�;D)4����sU���)Kͧ�!���am��d�n����tJß���:ru���m(s�v&����l���w=����=؁��A慫su�a��8�g��z���bRm�A�ch��6݂�۲"��=�X��3s&NH�5I�	�UR-��s�E'��j�9�`��-*��>l鍩f����|�:��E��h��< n�5&W����쾦:����[ ڝ͓=s�9h���֍ݴy3�X6��n� �1�36G��A������ϗ�/m�4[���y�P�� �C6�J�p�v�h�v�ŝH�����e;
M�$�s/Y�.ˌ<�>�^�`^4s�gr:��v9 �����v&ꩉu�[�)H�ha��^�]B�f=ey��5�@��+�%M���Z.6譮F��9����VxZ��v.����vʛn'k&�a��q(8k7�@U�jޛ#ul�(;	��rM]U[UJP*���dZ����q�jYJ�Q M�ѡ,e�"b�c�\��]9'	3k�{	��X�,Ľ��L][��	���m�sН�^�S]��!���-�*��Kb��5@��A��'J8�s�nL�`�۲ٙ�SZ�zQ>?(���|�}ڧ�Tz�R"�W�(��R!V-Q� ���PN@"&"|
�O��"�9����=GA�ќ���u��t9$��p�x{m{�8x�m�x֘@L�Kj��OG9��E��l���mL*@{L�փn�%,���%��em���ge�u��T;b�Áa�9ktnړi}�4)B�d�Ĥ�\,��͍�z���n��X����Q��=�ظ�y�#�ܸ�i��s�;��I�wHC�
B2�V7�[6���e4ڄ� �٬un��=e�؀�AE�
�̶��'�%9)�D�{�ͧ"X�%���}�ND�,K�w�6��L�bX������r%�^B�w���OK��@����^%���}�ND�,K��m9ı,K��m9ı,Og��m9��������B�$LC.���r{y
�%����6��bX�%������bX�'��{6��bX�'���m9�B���|c�c(�*��r{y�%�}����"X�%����ͧ"X�%���}�ND�,�w�6��oMzk��}K~��)�U_:{zX�%����ͧ"X�%����f��Kı?���ND�,K��{[��9)�NJr~��z_�&�-��.`[ڣh�]bwģ����,�B6!��f�h��6K55���Ƭ��	�O��^��׏�k��iȖ%�b}���ӑ,Kľ�����V~��,K�����r%�NJr~��ow錍ښ\���'��NK�����!�0(�����%�y�m9ı,Og{��r%�bX����Kı>�iO^k
Rh�h�˚Ѵ�Kı/�����Kı;�{ٴ�Kı=�w�iȖ%�b}���ӑ,K����K��$��4f�n���"X�%����ͧ"X�%��뾻ND�,K�w�6��bX�%������bX�'��r�Y��t]e�fӑ,K��u�]�%��C����������%����uv骷V��!�-y얥e��c8�l,�004�Z	e�%�qD��9<��w��ym��<V�~�Us��<��%�^j�6e��M� N��[%�ob�=��{;���~=��;+.ƫ^��｛�w���r	�"D_�Ő(�
��W9�Y.}��nǀoM��&6St+h�w������s� ����	�d�t�8�.��at��7fV N���%�n���%������� \κ�4c��]��͎Z0�&������(���cs�,�W\���<Wd�-�xf̬���.�0�V�$��5vK�W9\�$yI��7��X;��݊�%I���uuj����`�2��*�=�� ��׀n���'t���N��6l��	ݏ �6^��Uer��Iu�XTJZ�&���-6۷X;�����'ob�6l��'omD;��ӶU��;N���`NNj�C�-9�+®�</]�b�xM2:vV]�V^����w@���� ٳ+ 'v<tѨ��ce7B��n�	�ذfǀ��l��8��y'~�,-�M������ 'v<T�x��X�U��T�؝Z��wc�5M��N�Ł�r�)��l��Yv-��%m����'ob�� N�x���s-��بq��Os]`�1��k2�FKѠ���뇴�@!\͡�!�f68��]����vό�0`�w]�'O�݈��Rbtp&j��r�)���W���;7K�4Vl�hC�a�SX��s����8�dMbB٦N`����1�E��[����<�~��N�mN��RQ^�A���6E�M�v�gs��@�[6�m�-�%�c"��ef�� d.@tݞ�մ�r�cm%��fV��3*c3P谶�tf�g��߯@6lx;�����7om
�j�im�[��fǀ��l�v�^���_���6��Κ����=�����'ob��)AhJi�e�-7C��Se���`� N�x�Ѩ��ce7B��n�	�ذM� 'v<)��r���<��]rV��ű5���뗀'm׎2������$�mF�
�QH!����0�����zy��ǀE6^v^���{wt�.J˲�����9&��!�$,"EI10>���ʧ�XD�^�ݗ�lxwD$������$��.�x��X{��� =�� �]eВl���WI[�v�, ���wc�5M��n��D�7j�n�]�X�c�	ݏ �6^;{ }D��m��t��Yf,&p��j�Z�L�A���y��nr��6Ô	�m&�wmզ��x;�����'ob��)AVԫv�6�n�'m����'ob��v^:kJ]�M����+w�Eݗ�l���'DM�JA�+~�Uʪ9�U\�R�/ ��^4�'*�V:S���x&ǀEݗ�E�/ ��/ ��D�IP:���]��Eݗ�E�/ ��/ &�xQ6S�;q�#V5IX�ca�U:ޭ[$���c���](�	�CJ�b���[zvK�"���	�v^�"�X	;j��]%n����RA�-�vn�y�~����{[3���W;��� ��/ ��^v^��4���n�l���"���"엀E߻���р!��־�$�{)Ӹ;j�an���"엀Eݗ�v<.����wE�V��c[�}7�o�f9���s]��ۉ@8J�4v��80;�I��7B����׀v<.���W>A�����O�e]Ӡ;i�w�v<.�.�x]�xwU*%�@��nӢ�.�.�x]�x7c�;�!'D�7V�J��vK�"���͏ 'v<�"�X	;j���WV��v^ vH�wc�5l��ms�9�LvZF��M!xm(�\��l[����t�![�t�k���ڣ��,p&���B�5qa��n��3IYh���csG�^�/T�٬�D�N��Չ�4WV`�����2�0$/&��5c 2`ˮ˷��=��\E����Q����D����mcs,���V�p<����l�\��N��Y(ٵ���lY��u@s��y���KY� �[��;���M��ԋ5%Ѐ�wC�������l�t��]��u����_cI8Lv���i�M�@>���vG�j�/�9U_ �׀uy/Z�.�ZV�	�ݷ��<V�x[���c�rNrZC��g����\����>�`n����F�y���x�z��鶚��탷x[���c�	���^4�'*ʻ�@*vӻw�j�/ 'dxT���e������iF�����.\�T7X�p٬�/�㝜�ngE���s��X7&d�3�� �^�V�x�WD��!�Z3E�5��?^����T��H"0T��&�P07{/ �엀�<�8��<]*�N����:�n�)=x���vG�v�ﻠy����K��W;����˞���y�RK�"���>Q)j2�؋n�����ǀuI/ ��/ ղ^ꪥ�/_��ح؇J����\sx��<Wa� V�F�JF\�gh�����!�gGZ9���o���[z~���K�	ݏ �^���ll��탷x]�x���wc�:���M�*ʻ�@*v�V� ղ^ N��nR\�\��JZ�φI���;aqӹ%�0�4�����%	L%�%0��rJD���[��p�)��	���~)8]�jsD�D�eu�EѠ$m���HA����0�FCmk�+d
2������ę��F�8A� H퐸���$	 @y.��y'a�K|1�k��E������K���Y% �f�BWA�Ě%����X[���!on�Q8-&L�X脆�(J
$6L!@�	t�7"EL8~��T�C��B��Ba�]j�A&ӊO��� 'C��> u�<�qĂh v���@?"'T����
�UUWdQ���e��S(bEҶ�c�x;��RK�"���5l��wt@�(�:�[����:���j�/ ղ^ I��v9n���Mt�F�b}lvl�p��y�n;vN^�l�`uE=RWfhD�$����w�ޝ����K�	6?W9UU�^�� ݎ�_��Sb�ctյ��<�s��{�� �{׀I{�KR�m:V�
����	6<V�x��`d� %EJ��;�l�'n���[%�^ŒI���'�N�:)H�B[[Fqzh�9��rOvgm��Se�6l��$�� �UR�{��zy��K�%vLuh�M�Į�T�,��k�G#th~�� v<o���ٺ����ɬ�)h�f	M6h�� y��= ��=p[%�^ŀw��B�C�n�-��ly���IS޼޹�g�~�����{�B��b2fZ��S޼Kذ�W9ďOy��<��e],M5Bcc�V� �l� �#�	6<-���]��wJ���ۼ �#�	6<-�����:T�H�����RD���o��K��47=Z�r���;s����'O1���v�;vt��a*2�[�r �ҧm	���n�[2�%[=�.�h��b��`�XN67�1r]GO����m���3]U�� ��,;-H�[��l����ɈV����&��iZ\��,��цN���'T[rgm���֬�nU�@�Qeq3����}dLt���Cd�%��[$����y�yB��
�p���Ԗ�H�B�;%�&�l�i�,�V�G*4�E��)���۾�x[%�M��M�+ %EKBS�v�Bv�[o �d�)��	�e`��^���l��uj�6� ��,�L� �c�5l��}C�eZ�E��Bl��������ޞx���	5� �uP�yI��m��lx���	5� ;$x��=j��7�0��s�FՁ�x�&�b�B�8Ts8��Ɲ�3f���[%�k� vH�\��zy��z��@�I��V� �\2W9\�W9�s��s��ʬ� ;$x����]��wJ��6�f vH�M�r��{׀{���>DQ)m�.�	�]��ꪮR^���<��x�p�	�< �h��jݱ�;t���E�^;0�G�v< ���QnR�앍�R	H���ZV��V����ЄD�Ri��W#t1�Ĩţ�6�yi;0�G�v<V�x��9VQm����l��{��s��H='��� ����)#v*��LH�m�M�� zO<V�xz�¨�H�B$!�! �XHI$!$��FH��E#B? �@9����rI�{�ܓﾴ��]�-�N���s��.{׀{|�`d� &�xݒ��@�I4��ջ�'c� vH�nǀj�/ �?~�ًn�3���[-�%�mۡ]QK���{&������$e�a���	W%, ��ݏ ղ^�xȊ%-����Л.� �c�r���Oz�/O^�d��W9T�z����Ƅ�n�^�� �l�V�xSe�s]�6[庵lw��qz��f䓽���'o~�nB�zD�D`4TѩE*A] �d#YB*T 0\(CE���U��/ ���ʰ�T
������ &�xT���%�.�"�����h0��-�%�8�+p'�h�]5�"f-�
��M�37k)\6�nǀuI/ ��^ n���J�嫺+bt�;o �^d� ݑ�ݏ �l.�@���V� ��^ wdxz�U\H��x��^��W.�1�Wm�-��� &�xV�x�*���}��:�/%�n��n��j��	��W+n{����rI���[�x��# "�%�Ͼ���IVW
��˵�jZ��")�V��^(Zln4{T�y�8���/[�Bi��KAv4�������Y�T�N�v��J��9N�4	sI�m95m��[��e֨f^������9�HLb�cD����ɴK��u =;�>]�O9�k�5�t��C��{t��vNnOv��Z�5��pb6h��8����.SFۦsy�k4.��#��99��p�;v��mWY��j.<���	��هr%��Ԇ΂%B�3.�F�A���-Xe|����)���#�ʮs��ޞx��%����n��x]����9I�y����:�K�>���]]ۥAt�v� ;�< ���[%�vK�;�D�c�E;��;�� M����������ԨNZ���n��I�x������� I���<�Me5̪�[����@�eVdgL�Y�RbK��2�j�0��tʹ4B�m:j��M���< �c�5l��w�����Wm�w��<��1`��.����nI�߻��v������i����~�L�d*������j�/ �l� ����n�Bm��7Bm��K�"�/ ;$x�*�I{�� ����l��uwm��"�/ ;$x&ǀj�/ �r������z���Th�n����_��Q��D�(��f�sz�v�5 ���#�'��y���d���E�0;�T�L���t��x��`uwv�Se�d� ��Bj]�:��S�orO���nI�����	�$U�b�S�� ]O���rI߻�nI����IL[i�V� �6^ M��͏ܪ�U/\�� ��t*/̧uwv�n�l� �W���)�^�o������H���K��;9m5���*��^�&ܺܢ9�nn����6�[��fǀE�^�l� �#�	QV���Ɓ7I6��K�5M��dx�c�r�\��Š��cM��]��n��=x6G�6<-���P�⫻t����;k &��fǀE�^�r��U\�T�_��)�Os^��s����5u2�F��2�x�c�"�/ �{ M���O|��w0U���cJ�`-cR�K�(���bH���7F���c�@;		�j�N�-����`���Uϐ�� ���u��V�
��t�w�l�� ;$x�c�5l��w�:8�һ�li���< ٱ��K�6^ŀ|��J2�6[lwm�͏ ղ^��, ����n�C���;t&��d�e�XT��	�~�$�]��8fM(!�V/>acFr����/IL��%`K/!���IK�u�kI�A�ZVRR1!��+iV��SP�	J!c5�Թ+	����m����{߰��Ƶ¼t�"�ف@�V�V	{�
jh�B�!$Fu!R��!$X� �`�d!,!BZБn�-�"B��5���Ȣ^{Z��`���?JJ��y�:��3f�����dd4��ak�%�5���רLS������j���	��a&�RR�]��i3����>&s�ۑ9�D! �I ��H1`@A>W?}͟)���#��m��@���Yk���as{4�YsA.j^�_k�gB�޾�'��`�{Kꯨᕛ���8�o�_���� _��Q���A�3!sK�X��������F$>�����q-[;+J�ɐ��akdG��.\�)K����lS=����| );��⧳���6,K6]i�f�
�e���ջ�܏#\�Km����cn!f�
欱��H�j�DlI�iL6̉V�v�jE%&Q�(卄�L���ݺ�QbT�����G����ܛ�,n��0��X݆��cd��(�Au(�*� kn`����Fٴ4W(0���օ$��T,Z �7P�5U�,b0b(�G+���D�)lp�x�n\���E��=vhϔ����^��D��<c�����gY��V]T\E�8ö*�q;�5hD�t1Z���	�FY�8�c�k��ܵq��LeLp�ϕ�ڄ�KZ�B�t�k��s�Lw6\�Qr7���[��|�{&A�p�oF�]�M��G/R0�#g����u�,2��r;%P�놋-��(�J\'v�v���F�\)-Z�2 ��f�[>���ڡ=��v��6�%f���F�Զ�P�;<���\r<�q `Qu�@u�ƺ5[
�`PfZ6�/P�(�p�Xw�����χS�Is�[����UR��N�1f�(�mc �PQ@Q4���@������V\v�s�S#��6-e�Z.{;5����r�
<�c��	k��q��X�݉�>�&�ٽ�����E�R�F�.j���@,�)cE��Cu.�i�Xr壥oa��v��C9,��ƙɭc\ч����GB��)뭂���g��.΢�QHkF:֬nX��P���ݫ�%��ή���o:��Ӱ1��[B��v����0������ۍ:�xZ�H/0s)sm�S��먨�Z��z+D�Pe�mu���*����4e����U�ʶ]�i����t�n7jګ�y��D��sl�;��']&N^��s�^8����wI�7I���9�H�*��cl�^�k�-�4�!����^�B3*�;t�W*�xqB�����������öS<�w�Y�fkS?

|
�&�
�A|
������(|�D�
m5�ț��_k5u�m4�M9����,����ôS��j_m�[��e�F��v9�Qfr�t�b����cl70-��r.�v��vC��=on75��l�y�K��1R�Z��@�+������Ye��SR#�p�a���4�|���p�8D��F\*3 ]kK-� �Ogm��=��ۘKuypqMS���rQ[K��8�)v9Q鹞z�,�8>�8�!|ρ�L[��m;��2�&%�Ț8�VZb�:�J�]QnHewd��
�庻m+n�˞X�%�͏ �$���'8��i];hv��Ix�c�5l��l��?UW7b����Ċt�Н�x=<�[%�/b�:�K�;��	��J؝*wm�[%�/b�:�K����.��I�����4��5� ��/ $�������qM�;�,ZE�+"kc]Kq���@s�.ǆ��@���Gp+���<]dj��m�?w��	6<�d�Mp�>�"4�٬%�j��nI;߻������F0�@�O
Tx��w��nI��k�r_��{��rH�>'t�GaLT��_ ��z�	#��d� �G�JGP�q��V��v��$����I�\�R�?y`���V�*��Bl�5l��H�ˑ`nE�~���aXTPmb�a�^}7^�c6��)Ƀ�]�c93^Qs�C��R�u�7n�l� �^6�^�s�_ �{׀I��X:V��Rm� ����9�$z_����x6G��q#�x��I&�B�M6;o ��y`�K�?  �*��� V�R���UV3ٞx;�<��t*.q����զ��d� ���d� ���*���+I�T&�V� &�x��o����?�%�T���+���ecT�hfkB��4Nu���Nv��qطf����;;Gf$�	��*�`�#�'c��Ix7c�%#�Rq�MU��lV��'nE�j�^ M��d� �j�V]�AN�����j�^ M��d� ����IT����7I;n�=�r���x=�<$���n�Ω*��È��t������$	�ʰt��I�x�G�N܋ �$� ����\�m���A�jP�%�ݽ���;uv�)�m���v�$���)*fi��+��|���v,T��nǀ$xwS����%umݦ��Iy�W*�IRz�{�xSe�R�Z���5Bm��xSe�����r�����{޼ �MWN�6�ۻM� l���x�%��8�
N6[*�]�+n��x�%�� l�����8C�����[Q�5ղڢ2N���q�u���i������{c��$F�-465�F馤bFE%Lܤ#�ͪ��ܑ��uĦ�}k���7����ns���Ľoj�۲5xط�C����ɛ*l�d�F���Ge`9�=���3O���$#���e+��4�0���T�L�;�į �@��øP�6;n
56���m�0�v0�/ӺO:I��K'K*�P��uu� �E�!MF�V8�����3k��ێcOb�ͳ�.<�o���)ն�۸T���M� 6IO �l�{����j��St4���9U\��{ާ�yzz�Rwy�$�/��%�7��39|����S�"�/ �$� �c�>�*�bt���iۧ�E6^�Ix&ǡ�'9�o�}�z��X`�q�[�\-��Ix&ǀ$��E6^��I��v"��`e[��� �tt�����W=v�9D���^X��M����K�x$� 6IO �Ix�%��pIݦ;�M� �%<|�W>�W.ȣ��|���lx��)8�l�j�m6�����5I/UURG�<�	���`MBs���!ն�ۼT��M� �rR�"�/ �ꢏ�n���Wt�|��I9=���|��� �$�zk���i��$ƐҥCX�ɠ�*[���B�BˇhU&�lդ��@�KhųDD� ���������M��j�_�\�����;����M��6����"�/ �$� �c�6\���E��C�.�c�x����$�~�6)аR�B��@*@�Y���"�4���[�䥀v^ŀ}JV�5eӦ��� I��.JX��`z��y�� ��/����M��x�%^%�Xˑ`� T�W(�ݖG�4�N�nkKb`v[a�����ڈ��Ý*b�ɰ۫=f��~ؒ�,eȰM� �$��>�I9ʨ�a�msz��}��I-���E�z� ��,M��,um]��I�m� ٱ���x�ذ�"�?��ћ��3�[���9ûﾛrN�;�'����O�*@�Pa�!�#�"&����ܓ���a���%c�������l� vH�RJ��\��V�E�j�D��L��ǭ����`���6b�0<�M��6q�2;�e�۴�_=~����IW�n܋ ���՗N��J�Wm`d� �$��7nE�l�{�\����|b�T�l����M�7nE�E$� ����-�;.�m[��W�n܋ �Ix�#��rNK����{�+�-�Va�h�������� �܋ �g9�I>�H�HBI�vN�n��5�P�J�6�\�����쉶���̰�%
B�ZH�H[
��@��%c	��B�c(\�����a۷=6p�亲��8�<�ڎ-�W,N�s�C����q��3 ��[�n�wJ����@��MsĨ+-�V��l�0��[����ECK�x���3�n7vu��d;M%sv�Ed�ɂ�X�ဋ,�C@�8bn]u*���?;�������N���??][���R���4�J�nu��]�lKz��ZB�e���]�h\�]��}%�K ��)%��@'W9tݧv�S�o �䥀oc����c�>������wM�;�K �� �G��%�K �5Ұ�q�%i�i�0I vlx�%,{0�4�lm:�wB�����c�$�)`��H��ڇ�(�M3�LS3]a444�s�v��v��ҵ�dk+<"����[Cmm������L ��`ou��u%*��V�m�X�8g���*�_(�O� ������[�v����$�)g��GdB~�V�V:�Л0����6^%�K ��M�����LJ�e�����	.JX�8`{�Ľ�y�b:�*�ݧI�n�	.JX��x$� ;6< ��z�.��������].��`�`L�kF4��BIsd�5����Y��FZۥ�� I#�͏ �䥀v�]�*�V�ui��H��c�6\��{#��K�ƭ��ؕ�Wm�fǀl�)a߫�uWdo��S�1�����XT��ɉI����8́�ö�w�˛7���g�Rr��1)�N�.|�ˇޒ�^6����M<�̡��sDMK;�k/�ۀb}�榍I��F~�� �Y�H"(�9��Q�`�F'9S���F89�2�����?�bFM���< e�ㆹ$fl�#�#�*.�!H o���X��;�
����!?�~(H����������JN����^�R�$��>����ַ��pC0��hw��.�\���͎����3\5y��\���$Z�s��Ҭ���!2�A�7u��k�ߚ�>$�tYU�B�%�K�	r}`Kw]��v�ؒ�H=�K�Y�
A�?��B�? �	֝�d�b�F����Ȥ *
�~IJ�%B@�_¢~�0C���� O�iA!�HEXĉ @	A��!$@�d���`| �bp?\��#/��{��n�˺+v&[m�.JX������r���������v|�h�3��-��%�� vlx˒�ݽ�H�"GK��ֺZ��Ə8���]V���@�,�׶Kݮ`�a��ƺ��m�H��c�6\���s� �}��'��!c�;�����m�fǀIrR�� $��ĉ� ���ӲݧJ��x�~�, ���I vlx�Eu��44]��ۥ�� I#�͏�z��������J���h��&�����������`ƺWb#)һ�n��x$� ;6<K����^��W|��J6�-��c2�سP�cs��ʢ�%�@�Kc�)��st �V�4L�е��X�%,Wd�W9\��{��w��h���J�O-���a�Ӝ�RD[�^ {���;/b�5�-�h��N��m�K ��/ $��ob����a���(���HV9���~�=~�� ���IrR�6^ŀI��K1ݔ�탶� �{%�K �{��\��T�=���T��L�V������F�\V�J�]h��&�]���G��Ȁ�s��l����Z�Vh]��5�K@��ͬ*�� ��Wh"k�7;��hLgA������znu״+]F]�؄�� �ݡ�M\Wy_^�!m���o)��uG�/]��3ሸ��]ӣ��β˵E�t�;w-ʃL0��maeJ�ҽs�����O{�ww]|�x���:˗A��3)Yt`�&���J�"B]]�8fhZ�)&6���E];-4��V�@�oޥ�l�� �Ix�ذ���.�Mv�bv�`/b�"�^��,K��~�KO=���>[,��v�z���e�X�%,e�X�ƪն��I[ۼe�X�%,e�XRK�6�ێ�ۻM1[b��	.JX�ذ���I{ݎ��-X<�͖���+6�K�/bL��켣�Y�P�+��M���8�q������۾XRK�$�� �䥀}������Xh�h��]�;{�����C�P��H�D��tTW��e|;�X�䥀I{&�+���l�x��`\��	/b�"�^��B�S�WcN�ڶ�	.JX��`I/ ��X�K�bHhj��V����$���	.E�IrR�?UW*�\�����ekd���q�e���X4�����`2��2����WK\��l�
{m��﷖��w�%�K ��X��v�i�hJ����\� �䥀Ir,)%�Jm�v����b�M6�	.JX����S��	(�����@�	����޻�ٹ'�Ͻw!���mKB��wm�ݺX�"�	$x�"�$�)`ݤ�⶝��t���X$� �+�����{��R�'��o@�y����јjڍZ���֋�Q��/3�� qˍf��{�e�;�����)��6[o ��X�%,K�`�<���;':�un�k �䥀Ir, �G�Ir,��I4��V��'n�%ȰI%Ȱ	.JX�֥t��[v6���H�	.E�IrR�ڥʪ8Ur�ȩ,����`H���*'��hwy���?^�ө�[i����x�"�$�)`I/ $�����j:���Uդ�MR�n����-�hDX;B&�C�5��,���ps�j�Z�1�������T��I�ʪ��~��"+D�zЬ���m�n���I%Ȱ����<���@��ҏеQ4&w����	.E�IrR�"�^&�.�'t�e��	.E�IrR�"�^ I#�;بC�SJ�V�6�	.JXRK�	$x�"����h�K2@�$(1�:���Pxl���ak^K�˞�'���49��u��x��m�E��=�-�ͳ����t�[�m���̽��.��Q[t-�e� ��m���X��fRTٕ��q��)�v�:�&;G��k9�x�:����g�+����m am�I��gaN�	��M�/lj��N�.Sr\k��k����*�T���l.8S�%�JX��\W�����/���;�I:C��w���E�`D�K0W�u��[c��(H�r�Ռ�LvJ��c�2�Q!�7�[�� �G�Ir,K������D�5E���n�I%Ȱ	.JXRK�
�V�.�6��E����$�%�K �Ix$� �Sn;���b�M6�	.JXRK�	$x�"�5�[Q!YM;�m��K �Ix$� ��X�%,��������Ze�.��1�G��+�4W�����q�{qΤ4��D2��P�qڵb*�7M[��~����$�%�K �Ix�(H�ĝ���+m�_{v��T�A �$���<��W*��.䥀E6^ I#�;؁$�0];un�k �䥀E$� �G�Ir,��HN��LN�,)%��<K�`\�����%1�-�6+w�H�	.E�IrR�"�^�Hʔ��۴	�ܱH�Mj����KF�F�`E�V2��z����X�k`5`�Wt�m���	.E�IrR�"�^ I#�6�ێ�ݶ����M�K����I%Ȱ]\�+)�wm�ۧ�E$� ����?���R���u��ܓ�9F�6��t�i2�&�w�H�	.E�I� �Ixd�$]bN�hwM�m�K�`G(�"�^ I#�?r�����Iڧl)ZN��0��C�0��e��bі�Q��Ґ���^Dv��	:l�t6�_�y��)%��<K�`�R����;�-�bMрE$� �G�l�$r���De5Cm�i[� �G�l�$r�T����-
ڵIڻo �r,H��%�*�}���p+�e	� L�%W�pj�sK��� �����!�����۶;c�&�$r�T��I��X[�J���f���;c)�%=�e�8��j���\Xf���.�k�U_-�����	$xˑz����=�?Q�I�Ա��m*���w�H��\�D��� ���F�Ixd�
��;�0wM�m�K�`G(�"�^ I#�;�l)Y�FV�>�������z��H�	.E�w�K���t�ݖ�1;t�	.E�/r���{�}޿I����ܓ�UTU��UTU��UU*� W�� _�UU�UU�@T�� �P�B �T B@T 0�EBB"@T"�B)P�@T �)P��T �P���B,EB,B$BP�DT"@T @T �T �T"�T �EB!P�P�P�DT"�T"DX@T"DT AQ"A�T"EaP��`1DX0DYDI��UQW�ꪢ������UUh ��UTU��UQW��UE_�UU�UTU��UQW�  U  *������)����cV��8( ���0�/�@
}  ����P V�B��}� �d�h
� v�]����;hQI*;���J P�A�c@ d��� ( ���@�*��  ( 	: �hh �4(6�4PV�"� *|    �]���(�u���m�<{t��{�-�x��ãs����F�xzY�;�{���������ww}��>  �oC�o���B���>�41C �[���6�}�lǴ�UV���^�t�����U�n�����4 �= }MMk� Z;�n�mm��>��n��׾�^my������U�Ϫ�����n�����^�p=w���y�w���m�(��/ @}�C����������{��7�p���z�`ӝ��Wҏ���o���!���� 7z@�B�R�a�t �<��έ��7�����q���`x}�}�Dkh�g�>�y������}�%���z;7�3��h� a���k�p8}U-� ͝s �`�|����7���;�}�}<�@0 t ��lh 2�P)Z8���w>ۻ�'}��4��t��sgA@��jE��tR�q觥7������;�M7 m� {��F���z ��ƀ���(^zR��<�J6tP��E)yg��l�:�E � ���@���S���=)F��   �t��(u��P
-:�k^�i����� ���Y�J.�(Y�va�n���ϰ����Y����  C g��`����w�������}����C�<�p��x��}��=�^��|D�&��R�� �=��IG��4  5?SʪT�<�H �Oi��O��J� h ���M��SM�ɐ�"B��� )�'�������q�����}>�_|?aϿ�EQW�֯�E]�����E_�U�"��QAT��k?������_	rS4h��<a�B�:a�[<�|<By���j�=���k^��
�t�og�iRĩ9t�n�Y�\v]�Q�R��eл�Щ�MM�4��4h�e7ɽh��A �B�R^j�G�5)��I��0ˉI�SPԤ��4������jk6���9��-�<�!$��IOu���yK�eވ{F6��$��h��=�[3�65���l�s�0����n�B��k�VO|6���n79ﹿC=�.!�yMf�$8K��LRP�IM�3Al3�7��n�y�<ɳ
y���-H��)]l��|�����6�[|���_{TU�
;x_{�z���S4ƳִIV�2�YF�K�m!����vK<���fF9kY�Gq��K������5ۚߞ��kď�iS%0,)LHP!SP`^{R�o��߳�B�B'��5#�g���\���\�G	<8VL�l�9�o�!��!L��$ca�9#�<��~�%�P�g���%�e��D� �f�6c��g�n�CP��3�cv�l!sS{�B扁��<3��!���$�ͺ��bB�&�SI���F�fke�)��&�a�T��K�#�Si�� ԕ�.r����2�q)�`@�p�`�"�2bЁ!b$B0"ȐH@�	$�T��1�B+bX��zr����Y%߲y���~Gg5)7��P�7���%����g<��L�l���v�RR�X��OO|��\�޽��2x_P=��B�}�����\H���3����O:��_c�W�G_j���5����_os�|�ָ^L�4nVXYij r:N�W��N����іkR���]�+*H�]�co���2��s��en�͙p���BCxd͖XO.S\xG|�]y��l焺��y�ia-��s<�8���<I�
�)L����ɨS#�׻Ѳ�^��f���߷xC��SC��M�)*D� �	BF�a�!�)�(bK�`Db��hq:u�N��]QK~>��tX�ON��]ߓ����󭣃����W������o�2P�A
g��ީ�&r;�.�yo���$�=٦��9M�Ȕ�#H�1!�	��}�s�y��׻�Ç�_M�<
�o���	�WO>�}�Y������{O��
�N��v��uߏ�#�JW9U��K����2�}��\s~OwMe��_?9�><�HH�h۫qԚ�ݮ�T�����<���9�zRBC�&c~�ݖs��Gæ���������qdV�����:[�����eo�jꨥv��>�;��Ů���U¨*��g���ߧ���>B�nk|���/ܜi�,J��U�ԐhbhC�`�w�P���ѽ�7�o��<��[(p�rM�DX��{4l�7�
�hߔ�4�ܼy��s[�|4M����K���xyɧxn�y8z��5��]��=ۭ�,�SF�ɣY6����d�F�ߚ�@�=4x�5�h��ѴU:����o7o�8>
�g�_.�n��9�\�z���w��t]�p�ۭx�^p�p�)��-r&��ϦOg��8!.bԑ\4�+!�)
aBL&7�������T�H��p�.��S�q����ɜ֦CA!�#$�!����0���%��7��8���#'�5l�W5�eKɉ+(᭒�䫲hݖM$��!XYIN9�$-��]�u	]�͛љ/��R��I�8��	�d"Nq�f܁rh�w,o�|�5��¤g������_q��y�Y��z{��f�=��o�L!u�z�xX>���f�s�w�X��1���)��&)�8K�\�M��21"V-d`�Yto�ɩ���4j!`X[�Ȕ����Y�0����(at{�Ó[٢7Ŕ�7���~s�9�HI�)[ϻ��J��
��P�+��<�ۮ
����{�_a�|�1�W���w�Y�U+�}��ڨ�)k���so﷕E*�ӿ��zHy��0�] HJ�Y�R��o~na��a����ĉ����������c��!�Y		 1�I��O|פީ��|�9Ú���B����m>�zUn}������=�W�	]�������f��}~�hB��BB�k���:�c;ߵ݊���^�"аO.�|�z{�K��'��; S��b��Xp"M\CJ�`�� �@c!HHbA�ґ�F#
`���!G��H�]�ĉ��!B$F�� F@V���g_9�I�_9=߿k^���z��y鼡���i���na�4J�;�7S�e�ڰ�,=��rsa}��ϐ��MC�Z�M�&���ju"�Ε|W)U�}}u�__[�F��˚�����rZ�]%�Ԏ���l0�#d/�	�ټ	�3��ߜ#�B�xjzlѷǗ�H����sZ)]��h!RC6������*�Oﯭ�h��Ums��QR�_#���g�����[%/�!Bti�#p�4Đ��e�B᫁��Y$XЕ.�t3F�kWZ�xK�][9$�¥a5tcV$I��J�(d���y���f%�Я�Ee�/+8�;���V�����&�k�y��N��9y���˗|9��'߂�h��H1��Y]xgʨ���~1��r�Ül淳��3�7sg�	�h�	��n�C2�9N���t���q��c�_tۘ����)�G��|���B�0��.yvF_���fC^�H{
��y��<�yOXa�aw$d�0� ���@4�8���߹�7�^{�s\��&h�5.	N�-С��y	�
L%�%e��3<�xbHY�Xe5 �	�B0�@�!��P��s��g�)��܆p�aT61!�&�7o<��e��R\�5灋�&5	
�V:3foSz	�k�È�	�`I�,t��my����Ô���4�IHy��9�=����X^g]�U9W��9(*�[[J������
ˀf�k�4�fp$�(KB3��y�S4�%�����э\R4���P�	%HP� V5�$P�yK.��w�??��yqK��߸]ޤ�Ӳ���*A����k,�;�ka,ˤ�'�^r�Æq�O1��d.u�%/09)���o��T�f��+;����Z�m%<au����J��V��R��Gg]w����T��˺�&���������ϴI����Ye�o�L�n������7���c�+�
�������[9�_@��o9���zg�{��`�"Ɛ��Uw
���&�XZb3��s���¤�!e���Z�\��R	3��H_P��!M��6��k{�Nk��s���Ym4o�߯��s�l�=�×�� zP=�$��՛甙��������Ml�楾��' K��DeC2����!\�qar���82�)�	q�)����͒�����V������*�uҾ��T<��s��V��|8��ᬾ��0�
� %�D�RH�RD����7�C��y�F�9�5�k����y�},��pl��S3�ka�7��:ѕ��o�R��V�U�W�Ϲ��÷�o2�<�y�!� �����4�MO��V���j����P��QE}U�o�%IRP�!Zo�.�\no���9�v!�o�y<$�{�^@�$.����XR��p�E���o�e2�3�FB�%2��H�.n���j���T�t�!��P�ؔ�B5"��Ѳ5��!BVT��!H�,�ecBH�!�1�H��!H�CF�ЂW����049�3���*���[�8$!$������N6y!�&C�p��E l�p�IrHB%đ�D����4�&�m�M�6j@�'��D���4��y�Nl��OykE�撞p�M?��5�,^KM?Bl�Q����:���*8|W��t4;��[����O=a盗��fSF�2�Ie%x\��C G��/��a�i���nkd��~��v��
��M�fy�}�2��y�Bh��\	��LHVk���P֝]f�Oxn������\������B�{!i
B�)�H��+��2�i
�h$Ha
� ¤(�!�T�I1&����J���![$���D	���e�\�%p��MH@��,��.jf�n�Ni�A@[�齽�P����w��y�~�kU��t7i�UP���>�k{}�5;�&˞�[�_�f�M����������,%.������Y��JS�C���˽���*^?�%��Q���-��Y�Ol�3��_R%|HWS5�����xB�y��5� ��15����X��jFt���0����ֶ��ݺ6����4e��bC|N<5
�������9(����	�(B�.IK�)�j0�!F-HQ�X F"BH ���;�s+~���;ْ��u�[K>k;��B�2�-��o�{O��tgΟ^Wّ�~d����M�ԁ\��ţ�L,�+:H��p"D�Q�>8@�MEb��t$
�4A!�v�S���K���z���3&���'����08K�����79�!
d��Z�g�tޥ��SF��z6ry�f�c��F���8�+�q%$# �C�%��Y�Ѷ5��pt������X�6�4Jx�|	B��9.i�]2�FS! I���q�@�c!��!x���ݬ���-�M�<(��]``P]ok/좑�P�RÐ��37%
`H���L�x�S5���__��i_kEo�:뿭v���g��TP��xm
��e|��i���}�Y��?����_j��t.��WTp}����x����Jq�Jr�Q��\{�3l0f�X$69��_c_4y�Zm%�E���ݺ���WU����Wu9�{��nZMf����l�5�s.3�%�<�8s��Ӭ�hq �r��)�NI���f�g����=���y��߮�@����l'0%(��qrǂ��Q�pkqؾ�*����������l���������y2��ߤ�k�<���'��(z��5.�=M�G���͜v{���%��8k�޼��?&l�갭|9Q��u����|�v��˧�w�L�/̦4��8�Dהۭ�)!�B:�-�y��>��_2y�-��׳
ܩ��ң售����w�3~�vU�MӔ1v�י�fP�3%�\�H\!p��[MCn��%e�ơ�NjkF�A�;Nˤ�������Ws�Uw���նm��	>�o��|�$aBnj>n�G�}>����Ѻ/*It�Uep�xsh�AB�;8U1GUEe/��Jǟ�>Y��v����T$��7�w~�ü
����Qp�|�UUUUUUUUUUj�U��j��V����Z�b�d..y;�v�-,S<�ri�c��˲�}S��]��mN�v|iR�,6���P�Ì=vrrT��b�UU�1�7��r�V=��v��5��5e�g�U�ؽe�X�
�����KS5���lu4ဵWg�}��ʿ+^�T�*B����K�T��Hꢶ*�:���Um�n�vP%N&5;�.��P��ڝr�z�����5++U��W5�Һ�Lc��wc��b0����V�(8������ܪg��AOf�kŴ�v�փ`���V�q\Rݲ��9n�Cm��yZ�vwŵ�V^�*
�]P�<��͕�*�v�@j��x�B��V���\>�7/h�,6���-�!ۢ�z�txe��nU���d㦜n�t�	�^��{���V�[�PUT��Tq���w�mS`+����a�]��ڍMP�n�]����{���SK��s��vd�
��	��ͻ,�,��� �z*����OG.V���agm�%y�;=:���-n}�ؼ��c�g���8�zƎ��W<����6�Q�F4��w>��\��wl�@�Ml<f�6��G�n��E�r�[Nt��M���1#��7UJu˶�Sj7Pi�I�i�Q�k�82ɺ��y��^���gOi ٶ�lP*��UP@��k�]/�@�ݝ�]+�r컮5�;��.
�
��g��$ۊ�[ƍl���V�n$.�^5U.��og�+�O<��KjLj+n�͍õU@v)�`9l�9ô�_DU�V]�n�<wa� d]�R�wLV��Y��]]>=w�7t���1#j&MG�
���SA̩���v��>�"k�i_(�˲�UUS��F�U/&�5<��Qu*�hwrN&���w�qP�Fڮ1�[L���TT�tq}}�������y ;D-mcO� t��:�j���6'eg������r�ݍWUT��ݦ���y����*��9��b'8�Hj�U��ܡ��;"xI�
^���5KUUJ�x���VM����g�.�uD�%�\�UUUU��Y�6l���0���2�p�Z�HUJ�ea��j_-�� 7� ����J�ܻ�h����]�Aq-@Umt��k��d�kjڪT���;n�k�������� ���v�q������;����A�Qn��ja�V� u�AJ�ׂ:��X7N�*�t�*�wn�A�J�*�z�������$d�*������U����z]�O�EUvE�Ls�5UUUUUUj��"�wMU*�U��j��0�ݪ7i�� ���@�Ѧ]��H�*ڭ"�ժ�E��C���,������b�mj�ժ�V�R�UU*�F�ms�e}&*�U$ j��کyjS���P0���]Pjy �UUUUUj����UER�1�l����\��Tڀ�
�Ԫ�s��<$*�Tm�J�Ţ�m�b�sF����U�������ڪ�� *�U����m��ꂂ�U m���R���Uʠ]UU@T��U�����-��j�d��c���K&i��4�Wj���*������z��{]2�X��������v������U���*��������~��~����VB٪�*���evn���[UU]UPUu+�UPUmUuUUS��yj���SutJ]��8�z����������%n	���^ 9��������es�U���s����Uav�AA��Xƥ5^�&���YY�ت��u�u�UUN�㪪������;m��\�UUU��Վ�T�O/J��
�~�-��C�[UUB�[VU�n����V'�j�U'iZ�Y�U�	���g��x�PG����W�umuP*�)r�Quu����j��i��C���٭���j�AAUU1\�5��ꪣ�A�����Z�VvU{f��UR庫iV�g*��P&Ǿ�>�<�+rU#ے�50j�`*U ��MV��s��A��[H�u��Pj�b�������i��-Uu,�\�핵ȥ8�ڠF{`��li�������9�[a�S5UT��Z�m���]���<�\譢� `Ŵ��� <�	�(O#qsZǜ0e��^UF=m����sW+i�1��J�r�l�tS*�UU�nۂ�RյE���������j��
��s��r�t�@VS�����5h/<�J�qW[P&�*j��傉�7UU�[.����9�����c�uj^˪�:o���n�����N�\c��d���ΰ��l�����qS4
n-��cF���T�(6�v���-� VՀkZť�T�=��\�W!`:�5GMm�mU�9k���HUn���`���ji䙧� �)P�;M6 ,��[��J]�:�w�ge�XA�Ѹ��{1�qU�I�KPo9익��<�.���3�˰�q��{I	�TP��5�f㭪� �cOj�<��-�MG�*�Z�v��|s�(������<�_��y��Յ^�6�`�%�L�@UWQm��;UTEmEF�`%9����Z4#�G�C]J$[����X�%� F��A ږ�V��+kt��;������Bv�	V�I���ҭ�`y��1�^ڊ(,�U�ׁ�����*�@�/��e�0��[*��0܏K7v�4��뼛�'H۬V�k5��n��w����uR��a���{n� ���j��V`�ݒ�Y��mm]�ڦ�mļ�ű��(��ֲ9ET%Y`�K�U�<������z�n�"^����n0�xˍ�0m�\ڪ݂����rY�mQ�~����^��Z!�\v�sx9)�R��=��ѵyV���fʑs�$������ҳ�3��vx0�N�F$a��b�[*�㍘j�8�a�/Rtd�s���/[תR��{�&�C&��L����QIu�#�[���V-�ꭥs`��q��������U�s6�xZAUUTAX��s��zj��]	�@�c�J
�
�:�%Uڭ���jڧ��j��W����j����)��1����Uڂu�F�W�
�T��>(��W��U��A�UUW��[���#��TF���M������+ʮ�j���f�vYV��U������=�I݇9�7]�
�d��=�U� �u�j����R[��{-�������r�d	�:C�#�lh�<@�l�4uU[��T:V������@���2m/�eW=�D��U�`���ך���►�V0��
��%bmD�2.Ӣמ��<��xB�����}��۲�˝�$媪�u���Ġl�pJ�j��DjyeCmV{��(t��lQy�7(���W��)./K�j��V�Ӷ!#�[�O$H��a�Y�v,����(�:�����6*���+��UTw�9��/��m��8s��c.!�-��NٓO�vC���p�vqU����U���kuȐ��Dt�������7S�J Z���_����-�a�.6�s�GUEu(Nt'`{퀃$t�U��5[K]lR�֗<=c�i2ct�����O��m���k�,s��ܺD�ӛ�utl+V���������1Ԫ�jN-��&v��� VLN�UGN�Ւպ�C�z��ccj�6#d�rHM��j�@j������U������ꪪ���hrԬ�qUTy����嫙�QCUUUT���V��������֠�)m��j9U.UT$ptdy�m��	V�����h�R�]��&���Ov�̩J֪��۫�U������5UUT�!5m�T�UUUUUU,ڣ<��Z��tUUTUm�m<�]UUR���R�A�8�jꪣU���b�(�V��n$2S[UU�ʷWϭ|��A��.��*���T
��������U�� %Z�������ڠA�T��^�J]��X�Z��r�UR��ʠڪ���YF�S� �T�W U6� ��'PPUUUJ��TY��������q�-��j��VX%�FK��ӡڀ�i�M�΃j�P4p��WT�TUUUUVڪ�*�V��m����]�����ګ���VP����%Z����������������b�� UǕ��7%AK�\�H�AmwuU UT�UU0��U�Wm[�E:*R%�V*�*�U*�����U��KU�N���?e{������2���Uu*�UT�UU�US���������V���j���%ؠ�[s�ڸZ���U^j�(z�)z����j���˶�J�\QW@Vԫ*ԝ �Q�T���2�3L`d�I �Q��IH�������*Wf�*��*���������8@
���UU��ETUS����*�[5UZ�V�U���X�v��m([L����8ٺ�a8�PU]R�2�q��U�/*�U[v�B��m���IvaP
����Uu��lP�N��b�e�������B
� h�K��Q<��wJ�0�5 Q�d^R:��@�+�������3M6�f��M=���b��Ă�uU�cc7UW*�Umx��Y���Rr/v�'���md�W�o��p�*������������j��b�MME��J�]8��n0�6�8�1��-}��|�}Ӱ��B�<F*==��6�ݑ���ćm�m&�i5��1�m%/b����<ˬ�3�1Un�f^3�� ����w��@`�<J\��A磴c���5����jAik��_�l��D5[y7���]�]m	���wR�JαT]:��,�v�ul���PlUZe���&5���[v���֗�v,��^
9�J:VX|�iU�����U����f�`a�,-��o{o*L��h�*��D��?��W�п
����@J����P� ؠ�(�E�h"��j���N��6(qWG�	��=Z����"!8"�X"�Tjxl =QC�>�.�>����@�J��>P�P�<D�+��M���=TP<D_SWC�p 4��A�F>�l4���/�������)̀`�#��"��8)C~��� 	�$`�j����H����>T�Q/ʃ�AQ|" mW0n�"'�PJ��J��UG��h���4P=Aى�1N>�3�D�����!�"��SFC�T8����2"F F H��BH1*�)$�"�*@�=�$!
!B�EYAdU(��0M�衱q���� T=A6�_G��L�""H h
�dHB$`�! ��U"��B@�$��HF2@��B��F$���*�j�0�pDA؏��ة�F0�����U Z�Z��Q�`Dd��!a%`X��Ee����D�TE:G���c$	��&9�� ���l�$��BV1!�#	�ѣ��!����B),>Q��P�=$19g� ���t�#@� �T� ����*��Q��"!�W1j0*���ȳ;�kRk-ֲ§�	q��40�f4e�7U۴t%��)WP��y}�#�\�
�Kl���uփ%p�M��9�sդ�@�X7;jΪ�:��ܖ�F�X��زnG0V;CY6(A](��T����T�:��<[�ύq�i��\Ƚ���X���r�ˇgy(�{�A�����,k����>79�P]ʚ�,-�,e�3���К0�cț��G$Y�5��Ǘ�XR3t�n�
2������ q;�7��q���!�f{�X�%���^�׫n��Gv���;H.������P�aa�4�m-u�ҕUd�Ņ��}��{Z^�	�9��4�,�\,f�M�ɡ������W�,`��j���Qɀv��QѵYWt��]�A��9�6%7%��l���sÎ2���vv���7�
�I�*��K`W���4T�lj(Ѱ�Fb��ն� �����+��p	n�2�;+p���,!,�g��,y���u�)T�nN'66k�`��>����ľ:)�9m��3t�Pc!R�\�t����͛�m[�fb�T%�i�˵ڮ';s�,pK��	�#jD���K��n[�;��J;���^�s�KpƶڠRC��ŰlH�`{i���⃭���l�FO�r�k�J�0�=���n��<��E��� "�x��-�̽q�<��$��e��\.�k��)�6���<vH�6�
�i 6�V��a�9T��۝�9#�prp��C�U@�ܢ��4m����$%	M�=j���Xvi9ʅ+���1�^A�i�NM�b���`�G���6i7Z��-�;e��lltGd��L�UUZ�@Gh�5�ĵ��*�B�9A�f��P�e��JW���)#��ogK>yp"�H)m���Y�hu�Cn�ȕk[�rљճ���k�ˡ����aY:ݥ24U��t�㫩L�r۪1��mێh�䩰�:�d�p�Q�N;0�r6i5�S5�E̲� �/TA4�T��T?"TH<@q�� x�\Q��1�&fY���`�B;+�	��f�:*��KMu� 5��g���h��S����g�:݌j���i&VLn4"�������8pn���0��=ɉhpb؆ݭ�S�p�a���z����5�kK�o1ɧXa��#�u��pjZ���h@�=e�U��rH�[��!��e�^�Z���V�z��޻�8��3����T�mGZ�ޤ��fL�2�C`��pyN���8��ˌ�)�,6�[�����C�W���� ���;���ʪ����V hD��V�N��&��� 7dx{&V�0���])WI:�I�.����ɕ�vG�� ��O�Z��ն��L��8`Gdx�#�7�	V+VҶ�wI��`�"�:���� �ɕ�}'�{ߨʻ<�a�[m2�dԓ��������k���Wh��lt<�d�d^�ĊN�_������ɕ�v\� 7��F���|��[o 7dy||a	d� Ё$mT���e%V��ZŲ�RBe�A1`�`T�>TC�N�nV�܋ �7c���arЕ���V�o �ɕ�l���Z�O< ���QF�D��؝��۬eȰ�[ I#�'d���hTWm�w�i�XT[ I#�'d��$��W��_���(m�vV�D��{��w0mE6b�1%�tD5	�1 �v]'E�Щ5i[ {���'d��$��ǀM�5(|Wc�J�i�o ��+ ��XT[ I#�W+���U���m���m�� ���XW�ߵ��< @x���_s[�y��e`l��v��V$Rv��:���l� �d��&܋ 7��\T��vS�բ�x6G�}�e`nE�uy��?~i_Mn�Wi2^,�V����Kw���l�똁���`q�z����s5�yt�5�ue������&܋ �ձ����Bۉ%E�;e��Xۑg��RF��� z{� ��+  D
��]�e��m`Qlx6G��ʤ���V�~��6jI:�S��E�jҶ�l� �ٕ�M�r�Q��WH�&��Q��_~����vUv:��v�m��e`nE�uE��� }ݻ�cN��i>j�/=Νr�<xo"���c&��mڞˉ�!n��.nU�9Y�=�{�������G�}$��>�s(v�n�T$6ـuj���G�}6e`�"��j˅]�[��Z�����ٕ�n܋ �j��k��j]��t�6�=\�Uqw��V%�� �j���#�5u!V�I*-�M��`��{�ۊy���x�X�W;��e*ƣ��vn65�jsq��c[3`K�V�Y\t�1��6�
j���?s=�����89��ҁS\+V�@�@�nj��'��qq��D��+!<�{q���Ip��|ފ\K�@�]�n��#QW�Dt�S6yoo.1�FC�� bӢ�h�}�+�v�m���r/O4�z� �!�}��4�h]�v�	apU��s�rrp��.�� �]�:@f	Md���.zۗA�7�����yS�^^� {c�B5��L~�o��<��#�'d��;�"�6h��8��MZV� wdy����H���X��`Qlx�we\(�c�;Wm�vL���+ �c��G�w���zkW.�bg+:N3��}���/)�l� ��+ �l�RM�7c�)M��ǀl� ��+ �｝�9�~�п@fH�q��j8�8�������fF��:%�H�Lu��.y͑wI��0�i��g���̬��+�\���y��)V�uh-�6�޳Zܓ�{�ͧ ����4�����#	!$��$�B��ѱtj@������b���Gb�3�vnI9��������iu.Ң�%mX[u�wve`�lx���	ݙX� $o%ڷi_Vف�UUr�.��x7�x�̬�\0�Hut�ZIЩ;�[x����e`���ǀ{�ޞ�*<4��@�P\W6/��ݺ��&�ۇ$��F��u���Ңi$�+�m�wfVٮ�6< ����JK*�6ۻl�-ݷXf�`���{#�'ve`n�e]�t7baH�`���{#«�ÕUA�+�[�Uv�9UU��fV�� �m�q+.���*�6�{#�'ve`��Cc��آ�Al�ۦ���'d��;5� ;� 7�<v:�c��8ya���J�mB���ql0���v���9��3�vv���\0�lx���I2��h%��v�د�ն`t����W	���=��Vٮ�$OA!�/U��
��E��}�N���;5� >�ǀN�vU�S-;	��x�̬߽��rIϧ�krq!��/��*�)W>�����RK)Sv��eYn��6k��s�K�'���� ����<�{Rw�у\��6��\���s��^�Q� �䗋�:����n,���ڜ�"����M� 6lx۳+ �{ n�e\Jˡݻ�J��o $���fV%�X�nǀZ-�EE�l�7V]��ove`^ŀT��M� �����B���+wt[u�I{ }Sc�	6<�ٕ���,�hW�i���ݏ $���f��>�=��I�"�k�\�w���#�º��!<��-�'J�Y�f��T��sA�5�����s�Ԇ��ѵ��������3��£�փ�ێ���<\[�rִF[�����l[��NxZu�K&��1qm���t�(�݌�}����gV�Z5�=v#uK���u��W��7 ��r���S�獈[6َl���a�k�yӣ(�M��+jKI�ڠT7&ˆ�u�m�5	R6ݴ3��ָ1҃��*lz���v��Exdݒ�8��+�c-��\��>���@����`^ŀT��	-iW�ʴ�TRv�o ����$�� >�����줲�V�o�ջ�� ��, ��ǀlx�fV�d�ʷl�SGv� }Sc�	6<{&V%�X:m�q]��v����x&ǀod��$�� ;Sc�6A+lCuO����-ٖ����}�4TWv��Q���\�hI�j���J!��f6^���}��^ŀ�����W9�|����媤4�0��ڬ�����O=�r�[$��UW+���G�wc�;�2�V�-��l�7i��V�x&ǀ}�2�	/b�$�$�%Z�V�;�V� I��n̬Kذ�ݏ ��U|��N�E'm�x�fV6�, ��ǀI��UW|��U�wN���CO/a��m٫�Hk�̙i;s�w%�y���\*�pa\���g���w��C� N���fV��ŕi�7b��� ��c�r�ă��<l�V6�,�9�$�Ny���S����x����ٕ���߹O�uO�wTH���xCZ!�$#HCYS5l�<��@��.��4����H� �H�2,� d�BSH�>Y	�e�'�x��"E5_i[�I�vː7�����C�͆Pq B@� �`�)�4�) ��`�5�.f$����c���׾��ą����w�<<<]A������̄&c,!����5�qאp\I�O5������\-����m�kjJd)	�C��P�G)�L��Ȭ&h�m	x�p�8\&V����͙�D�raߴc6��/���7݋�n��v$!B$�3ݗE3D3Z�bܾ��n���/4l����"Hh��(���T�DWH��@8F+U�@�,����V*!����	�<�>��I���< ��-∺-ڤ�X��wfV6�,�ǁ�r�/o���T�tyV�Wm�m�6�,�c��� �l��>]�*ۻ*�:v�*N��	�7lZ�G�yd�G�	ä3z�U�wp.�s�)ô���v�X�VǀI;�'�rz[���ym�� 7�b3L� �H���X��XV��=\�)#�.*�y�n�*);�m�����n�ŀ� }$x{%%���n��Nջm��{ M���#��^��0��2!`@C�J�,N3�䛒G�wߧ@�߽�f˅Ń � ���R�^;�+ ݽ�t����9�8���A�;Z8��!�lݱ�z���4��� ���"��Ѻ˶� ���N���7ob�	ݏ 6�Kj���;L�Jշ�N���7ob�	ݏ 'dx���U|�ui�vۡ�X�ذvG��<n̬ ���K��)��� ���� �ٕ�M�� �$�;�T�*N˶�vG�N���&�ŀ�z��� aBV	�\H@�2Kq^��;��;[��$(��s���	pō��x�H�L@����n�,��5~��b\;�;r�����x���H�ٶ�p�����$9J��2F��b�M�[n�td�sD)�n'�	�N�p�{�#�t;�8���֍���� ��Du��r!	���f������4����'X-��Z&���$K���Z����]f�afe���QD�.�L�k����UgMYTj.�LC7b��Kf�hVT�����T�a���r�}镀M� ���vG�w�RT�.ݫ�)ڷv�`u� 'v< ����2��N,���*h�ճ 'v< ����2�	��VՑ�"�[m��7fV&�`� 6���Q�Bv����Mٕ�~�s����x���< �c�=/B���B\gE2`�SCh7B%��9R���c�h0�q�.�\][!�f�����X���< �c�9\�r���� ���z�[V&��0{#��Y\��*�����^��+ �^�>���_��:ߌA���W�m��� �ٕ�I�����8Smڢ���xf̬Mp�� �6^�d��VYm+WL�Ӷ� ٮ������;6e`�M��i�:��7��Itn8Ӽ�c��H��\e��z
��f�Y�����~�	���5M��vl��6k� n����M
��m����&���6k� N��kh[Up,���J��{��7$��u���
PM
�"����PpJ�	!��@��ﵸ� թ$m]JUi�vۡ�X�p�	� l��?��}� $R����]����`{#�=Jo����e`�e`��\������v��eǶ�N����ؽ�=t)�;x���&a�i��k��´��a��'B���@=�ߞ�ɕ�vI��U|�����k�;(M�TRv6��ɕ�������߲�Oߞ l��T����$��15t�-�n�	�{+ ��/�9Wv�����%�~�X�K�����qPJY�3�@�M��'�[}���9m�{�l���B4N@�?(�4�tG�;���-����sZs5Y���ʧ����_} ����{A%�����$�떳ܻ��Us��_~-&��{���YƎ.�>��kG=m��%�wi�t���lb�g$��B������r���?g�eݽ33߻���>�r�S��6�w�} ��I٧Й��X� ����9�fe�}��ݶ�9�����w�쥞��.�% *��WN��O���Wz�R���I%꽞��W�ڪ�6���+x w�߽�s��{�u�Q��6u�v�&f{�{�s�3/��ٛ�����r���9&���}��x }����Q�s�,5�k���3��xf��T�>��ޞ�m����]�m�����-��$���� @s�=���2�sZ��qv�;�0�P\qՄn��a�7jz+�3p���{&�8N6w�ęn���,�G�Od�Q�7[tiLn���	��S�ư��k��%��P=�mf�-�xrу�Eab����Dru)�9T����3Ǝmc��{��w2�wr(Fb+��+ۉl�;>%��v'K�:�).��fxq�^�����gL������>�NO|�͡�FcŖ�@�Ü��h�2��=
����Zj�8���M��?I6�
���u�Vn�����} �u�c�I-���+����{*����]�x��Z��`�&�} ���<�m�'�������߼���{�g����`���X���؛v�$���|�Sne,Kܪ��������_�� O�N��.\VZe��K�+������KIO߿}_|�[z�I}9��~�������	��ʴXbI.�>��I/G3־II�<�$�.e ��VSD�AJ����R��C]n�Y7�X��gkc�9wK"lr�t��>�$���X�In���$�.d< ?��;}���m�f ͗.��}��s�� ��`����$%X�BR��wAI�*��CG @�*�D4 �w��l��������%��ZĒ[��U���1Rv�o�K�L�Ē]�!��%��ZĒG��޾��w�--�7;$�QY� ]�!��%��ZĒKd��K��RĒ=��g��j�Ƙ&���������.{�}�IyOe^$��2|�Z���ۦC\�#�͕0���9�r��3�1��ʩՋq�}u�)^���J�I-�?�I(�e^$��2|�R��^ ���ؖwbqYq��@:��I%$�}�IK�-bI%$��Kn�IJ �]]��m��I)&C�J^��v�P}��!H(�PN(eW1�G��%�L�ĒKjR���.���wl�䒗�ZĒJI�$�[2��{�;}����^�Fb�rĒJI�$�[2�II2|�R�˽���<�9V�6�i[M01��t�7�/,��7��$���DC�I��p�<Yz��;�m��IE�*�$��!��%/_q� w����{��6gd�g-��I)&C�J\r�$�RH��$���o {���mb�`�V��tr�$�RH��{�Ww��e^$����>� ;��xf�m�9��m��|��[�����m����-�� F=���|���-ݶ����a{����ui[��I(�ʼI%���?~����Ԓ���w{��:β�XE%ᶮ���H��7j��KY�n'/�V�b�	��R�$�](�y4���aa���y���	�bI)rK�*��I{�쥉$��T��nљ�Gf��z�>��&�>�{���%��x�JI���Ur���"B���3a�_ ��}���w�M�^��U����|�S�،I%�I��h�f#t����rrs�9�����7��߳���%��F$�U˻�����%�ޡRE�pv�&�Y� ;�����99�s��~�:�I~�����6L��$�����}W)��[+�;�o��@�)p
�S��!����$�JJ�i��"ƉI���"!#E!H��`D�V]]��,�������g<c����޸|wx���\���Q�ى
�����$.2��Rd�	s\deĐCW\q=�4:[�3����B\%sF�LpK�'3@�q� v/��s���jBՎ�*�@���F�̞�B2�$cK	"I!�

Ƅ����#���ٽ!��2I ��(����en��^pw�#���@����e���J�!˗�ăc�$|߬�jd!	|�R�$-`E�#X�)<�V%"Y+ �m�D���� 3 �I0�� �!I&��+0!�>�j�>�<[���s�
A���m��Le�%0�C T�\6R��?2�K�ӑ��RW�bv�s� �$�ag��63@����A�r'|}�+j�ͷ+b��/���q�����[ k�=�Gm�-�ǢL��t��t,���*���e�ts<�\ه�e8n�v�+ �D�Hv���Wm��	<-/g��5˹����}�"Db�t{�v�ZHxyuY�\�HI��ǉ�$1�<�V��a�u��ll�Kk�#�rsg�F�����1��f[^��!:�>7�VP�ۍs��7��5�780�;E�q]� b��l�
%eiQc���V��rh �q�P���]���.k�y1�E�v�+Tj`-�N|���f�jG���\�ȹ�N�e�X�ۤy�����U=Uk�ǨQQ)�n[MMŐR8�)�AP��J��l	C+t ZwE���S62n]Yv �h��^����GR�E�C�b�B)V�Ŷ���!�5g5�Э�M�zѵʝJ[Dvz �^�����
��%���vF7�՗���֞�9��Զ.��z�q�{u�%�-��]͋���L�h�=2+�|s�f�l1P��c����0��!�H�۴J1x��i쒣�x��p�L�K">쐨�/]���Ha��`g:X7Z�<��#s�mBB�Ɖ�Yu��VB��T���r���	��;v.�s�l�c�\��D���,��l�G���t��v�2}��珞ѹau֎ ژ�U	�;���"�7-�ӵ��F��N��tDbr�|g`B������� rx:����m�OLv�x���hn�D&�36�Ye�"�����2��fl�]�X3��T�I[ud�*�K�¤��96�������m���G���JS\h�Y� p�v,��'d��'U-UU�y'&����#��[���Vtf��e�ۻ���#��v-�9�/0Q;Z���9Xe%@���X8���"��ݫd��d�Ut�������ع-aV,���Y�m�1����یٙi� ��K�[ٵ ���t���N��9K�I�tMfh�d�5�b�'�Ut �ء�� � |~^#��
�P<z|��hg''��ق�Ԭ5θ�uS����=����:{)�#�+v�\-��&;��竖x㑧IÕh��9�f
E����Қ����[Rv�ps9tF޶n;t�Ŷ��\zu����u��Yf�5O�xÁؖ���N�VM��q�:��Inl`(��y���)Q\F��a��;p	u��x�M,�d|!�\:�6Ờʄ�\�3Mu���/$���$��O��}���Hb��T5WgH�E��2�,���ۅ���q����������w���4�0���/������_�{�~����}���@�~�yt`�A;v�X�II#��s�v��e<I%�{<}������ɶ�?��kC�5.2����y ��v���$��8�ߗ�x �~������콚M3M4]p����~���������������9&>��c� v};�C�M����ޯC��I7�}���~��#�����} ��S���4��K��۝uԊE�=˫GTPA�����D���~�[H3O���6\z }�Ͼ�^��G�$����ʪ�\�i/�����$����S���n����@/{�#�$�%�䰊 E�C�(�A�B ����_������%.?ֱ$E$���~�U]�~�B��_�;�N�������X�p���R^^�� ='��څb.�v�Wb*ӷX�q{�<`^�� $��?s�m��g�ϟ>�������Y�7t�f M���U/zy�����I������/��!k��&r<bܝ��A3gE���:b6��T1����Nk�;J[WEݷ��<�	�e`k���rI��9?`?���@���c�4��X��x�2���RG��� z{� ;6<�rr��}=ږ�YE�΁�?�N{�����j�TS5��w7$�߻�rI��ܘ}M]K�3Z���?��U����E�߯ ������r�~���ǥ�;��lM+�W�~� I=�����	��`�#��EԤ˵]�5����q�<�q��8�7�9���n:'�����rw��-���Ι�i�o�{��}�� >��Uϐl��wޯ��)�-]���f���9�H;=�l��wu�=ʤ�lO͠.����v� ;=�un����%�?g���y<��Oe�#n������'7��f�w��nI�~��r~U$$G`A���hS�/�{�߳rN�쟪��]&][tݫn��̬ܮUv{<|��<�v^��%%[Wj��L��r��;/�0f|��-"����n�%ƻ�֬��NrJ�WZj�����`�#�:�e���|�d�V tԼ]��5Md��sZ��N{����G�>����'��+ �c�{�\H�����wn��.��v��g� �ٕ�������X��z���Jz�Kt��&˺rqI=�`�{+ >�<UU-������6#�C�Vt�����?�I'�W*���ϠE=��ݙXUg
���w����ݷ�(�B�Rj���t�6r�8ø*��c��m6865
��rޥ7�q1��$
b�2��X�H�x��v��ܐ��h=̞1�>���;�qFU�V��tx��xĄ���qg��;����@�au�ܘ�ۗV�D:.���r&J���P"��?��[},��KP�PE�- a�``ک������M��7m���M3�GYw9?s���{Cf�4�gYk��e-�". !��7p8z��o�}��C���=���,}u����t�x����ŀn���s� ���X*D]]#Ԓ�lWE�o �ob�꤉'��ｕ�I~�q#QU�����V�6�ۼI���+Ur�;�y���}���_&��2��gC�N-��V w���>[%�{�JI� 7ʞ�c�ck,vg@?��נ��O��k����=�~��;�2�vQcuz��͈��sòv��{�h�^1�zȶ<]�Y莃�&�jjvl�1evr����׀n���;�2�Uϐ����z���k,�f���f�rO}�훂�����xc����y�-���9\�W��]���ꬥvSl����M���e`)%��W���G� ��X��I;�X�qv��^�=��7ob��9T�O}X*D]]z�I]6+�J��-���ذ�̬�$��!:�$'gB��0dɂ�햲`:/Lz9��;8ڮ�ۤQ��ӓ�D�6�Ҧ�b����<��̬�$�W+����< �}/�/�ee�m[�?y��ߤ�J��{׀���7ob�r�\�A�H�eשSIҡҶ������#Õ�Uq @�C��訞s�gݻ�w|�`�h˴�E��V������%7�x�<��p��U_���������/��?س-M��3�/@��締z�������:��^ odx��&�-z�DcM���w>;�4�;w`�MÙ���� �V�7X�
�0��n6�0�E������o����>RK���W9ϐIs� ��,t�E��P%cm���竜�$}�Is� ����U~�UU�z��]_�Ē�m+�wm���� ��Ň�\������y�F�l.U�eշM�6�=�R��=� �dxU\�T�	�O���s��rI��:a��a�֊�m`/b��G�6<�{��䓟����fL<�ۉu����y������]����Sq�F[�[V?���q�!ҡ�m��o�~x����ؽʪ��{+ ����ݶ�i	ݦ� ody�s����������y������}�����+̹�k����|�;$���\�]S޼ ��x�eVR�m61"�&�W+�}�}XW�����{;�c�;��RUcM��^�s�R{��$��vI��_
C��'��ݭ����m0�0�mbhKQ���R��-h�o1Ɔ�u]��L۠k�]SYe��S��X�\k�+rp!zEq����,=��҈�����)�m�pq�g��n�����+hܮ]�v;����d���Ʊ��羾\W&��k;]�'C
;k�@nV4睡�4n��q�8C�1K��m��{n�6�;z�**�������b�M�������5����a4@���n��hƕ�و�h����KB�a2�.�s���Fi�a$��J��[� o�����`�ezNs���}������պe�G.ݽ�=Uʤ�����uOz��#��q ��%��Ӷ��M;f����>[%����RF�y�#�� ��C�P�]���9\���z���xw_�r~Q?*}���ܓ����7����(�n����9�ql��{+ ��{�����c�]���&�6P�z�7V��c!x���);�:�l�5�.���9�Qv�յn��wc�;�2��8z�\���<�{�����;2�p��͜��sϾپ+O��!P�0�@�
H��h��"���Ī����Kah��7,GPP004(D���5� 5>;ߟ� ��y`�Ǟ�W+��F�yce'HT�R���`������ܠ�" �N����'�~��rI���2_�	%uc��� �ob�ݏ ��e`z��\�8�=�0Q(����6+��ݻm`wc�=�r�ʪ���W�vy��?~�{z�����atl�Zњdn�Y�ј�]ƈ<]� ����4��v��7���rNL�;�Y�]4�]
�m�w���>ۑ`��^�UUU|��<��*=j��ZT�P�]��>ۑ`��X����&O?NO�rs�k�����vL��)�ﳿ���}�[�y��O�D�Y�HGA��&!�1���� !Ed e)�@��R2D�}������6	�+0���JK�3�Y$�"�dh�0\4�5�P�-�P�e	p%!0����!t+3� ��ё$@���9��l	�),ٙ4�$�$!�	+������ACP.WB3a$���/�0LH�H�2��-%2�Q�@�"j�X� �Bp9 �!���Js���aH���x��M6��A�s�b�Æ��iy1,14�h�&����hk- D�F(���։(8��"�$*B�R���������1'����eݎ�cxk~}B�! V�D�	BS@��t�(x�/����)�~���i<� (
�Q�5C� 6<� :> |P�/UJ���w+ ݹ�uIP-[n��ulV���9��R['�ݞ��>RK�>��X�J����cb�N��>�̬�\�s��z�v� n�x[B�7w/�Xy-0�<�س��k�9��˸�k���&4m�������(FZF4!�[�����x{{ n����?W*������V z�G��*t�We:��V� �ob�ݏ ��e`)%竜��GTH��*lWMӶ�O<�ɕ��?�g���ٹ'�g]�'���2f|L����SM�UUW)w}� �����X�\��r��d��bTK�r�J�*%n���x�\�*�\��d��>�̬�9U�O2۶���1�S�%i[�<n;iFú��s���L��X�7i�����<�I�vݢГ�}e���ݏ ��ez�UU_ ��`��v�݂���+m`�ǀ}�2��p�=��ӿs�������7b����͜���e`Hᇪ��IzG� $�x����R2��3�NrO�I&�~��� ��?� n�x�X�����$��:�����p�?W+��\������?O߲��8`�\���+�&�j�B�gMݜ�[!��+�]���2�%B4�t��l����c�rV�Y9Ȯ�Sc\]#r�8lM@`�v�TtF�˃G�&{`�XZ�j�!SB�Bheŕ�k��[r&	Z�1���GbS�j[���we��6�1��֬�7t�&T���]����Rm�lb�(p�ȥ�yD��{pV�齢L�?���N��w��R��zС�Ú&h�H�o+�շ�p�8㝱�D���ٞ�ø��s�]��9���No1]���h�h�>�;��� ��+ �nE�Mٕ�����\��eЩ��;&V{��:��x�{+ ;�z�T�O%�w�I*�T:J�`S޼�fV�W�s�vO{��=?~��$6cC��E�M$���2�����2�=�U.��� �<xmڰV���7X���Ur���W�uOz�	�e`�(���V�i].���Y̼�K(��=ͻ�,;vv�T���[=����˱��Uv�l�X�d�n̯Us���w}��O���;N�F䜿}�o
���T1 #�UT�+��ʧ���ﲰwߞ;&V mm-"���WL�]�w�Mٕ��<=��^�{+ ��z���E�ҩV�][�۬ת���l	��VݽJ�R���`�R��y�ƭ�B���{&V�0͙X�#����c����8��P�f�u�'<�l�j���R�h%ѩ��j���%�%ǒ��	X����vl�������&��X�{��E۲��&��`�2�vG�od��;#�{�\H�<xv�X+j�`�� ��x�L���UWp8r$!0Đ!#�Q�E���b@�5@�C�*�]�c�`����N�U��j��B���m�{&V�0�2�=U\�����<�����5c�u�v\� �s�����|'���2�����l�Se���͠񘁤K�	�!��Z@�����B��[t8��&��d}��+ 7dx�_��_���+�����/��i��C:�%��:����NNq"O{+ �_���2�j-��������Tշ�nɕ�vG=�Us������	=��Ԣ�WJ�I[�W9�U-�������vG��(��D�#�=���rN}>�|j幬��i�f��+ �9\�R��$�g@�篧@<���ْ�4`�2�mʆ ��D��8i��R1n�l�l�𢄵�ٮ>�9�#�²�M�Э�cn� ��<wfVݹ�W>A�{�X���2ںJ�eզ��7veg�UU����vE����7���X�#�ܪ�ܪ���'�,���L)�wtպ�"����I2�wc�7ve`�����e�՚ۋ���I$���� $�x�̬r�UK��x�5E��������n�ـ����I=�rI�{���9���nI��,D|U($P �"@T��D�	{��.�(���R�attj��:��Y�Nq��v��8A��q̸콍I+����c����S�-ֳ�2q;J\�ɍ���nhI�:;qŻ���vv��;q�Iz�{�qӈa.����^5�\�ӓVLcM��\���h��.��Չ�eH�`�Yu�2zLP�8.WnT��X�v��+�p��=mY�3mE�Ֆ8D�S\�C�'s��;��߮t�\�����0��K���]�q̆��t�40㈇f+\��{���%�?QWN�*i��7}�+ �G����bU�V�H�T:Wn��p�s�\H���O<��+=�URG�D�/]�un��4ճ ��`�ǀn���>�"���M6]	��`�0=U�RRO<l�V�^��s�~@s����'�e7��[��\�e�7�ove`-����`wc�>������&�jƲ�ʸ4N;v,�^�b��L��a�:ݍ�A���$�oc�B(v�v�o���}5� ;����?W9�����~�ym�O���&m�rN}� 1���GZ��{��$�l��>ۑg��W"���N����t���0d��7�2���K���w������i�ZѺ:[�C��I%��}�`�~0��`z��ĶO< �J�*�"�-:�n��p�?s��9�L���� �� vD��&ݖ��1�̈́ư�&%�1-h��mx���Kq��0?��9Č�-bJ�6]�1�g�w���ݏ ����ڸ�N�*�ݻ6� ����ʪ�����;�?�\3��*�#�OZ�n�Ҷ�2�Ӷ�	���>�� ���s�s�Ⰲ  B2���$�##	"1��D�~HN��UVd��`�y���e:aB��˵C�`~�r��}��w���ݏ �� mmm���HV�v����>��`��*����&�� �\� �H�Y�-���smxMCr�bd�p�e)=<�Bu����.+"E������}��wFT�V˷ I<��p�>�� �\� 6�ں��hj��%M6�ݙY��ʪ��s��ٿ�?������ lJ�\E���v� �G�$�=\�r��$�x��X��8+�t�cV�s�\�qv��^ I<�ݙX���P}A�My���ܒy��}aj�+D2ހy瞽�$��9�I+����@�ߟ� �\� ��jR��cTĉ)����G6R���M� ݳ���&�u@玭rm���[��4���<��{:�8`K�{��W9U�I�n�c�B���#Vt�}};�''99i���� I<�ݙY��\�H%J�G�ui�m��m`��� ݽ���9\�JI���y`Z��C�bWv��l�w�n���+ �\��\��.��� %yJ��6��wI4��̬�r,�$�w\0�sj�)U.:�b�B����)0�X�����������&)"B�C�x�h����'�%�HM\�h��2��`B���2��U$��	�U�]��[	n]�	n�q��hJ�$��цL~�ld���F),,�%��15���[��JB̥.�' ey��IKd�%���4���4��c��-�-�YL�G���Z*��i#% Y��!!�Hib�c!8��8B���_���UVWǺ���w{�0ps��@;u9�n�Z���0�cE�`�n+!�.����v� {�:�ȯX�Zȥ+��۳�a򵌘��ù�D&S;BV:�ns�^q5�v�l�=�� �|�m�G���6ۉ��z<��M�z4]��Қm;q�K����u^Ú�5��B掩Q���n{Yp�ۖ����m�g��	ɺ� e�&�y�����v�n����ٟn^�۩P�D�ģ�%%t�d��-m�Gf'nt��m]-*:��<�&6� �!ը�\�y]Ev�By�,��j۫�5ʻm+�UA�^dԪb���M<�e�Z�i�&tUj���V�mc�x�hV��E	�!� *�-mht��3�ƴ�CFCU��R*[���ru�c��Ob�^�*��A]��Iɵ���;�����j����9��l�2x� ���t��y^����`��ɲ�ny��8��6��\��}cvz7^ݻ �ɮ$��-���h9�y���v�v�d��g�ծ ��Ӝ�QBu�N����8m�ƍ�NLK�x��z�#��t=�4��[tkD�7Z���XD0{�^E�tS�<{B���K��"���t�J:�#�Hk&�K+R�W����H/Gn:�H�x� ��PM��kk�Aջ;��b��uQ�a��K�<Z�,�l�����`�ljkH1�5*AJ9b��\#t+���B)r�:�	t5\��kt��qQk;'<9�@w8��@<(���
�q���aWEq�m�EUR��`D�2V�<D�CNܭU�i$����JV�FM��d������eP.q�Bp��2�Y�B�cu�El���Pإ�h�����$����������(���B��f�����\`a��S�Y����\ۍ����bu@�;��L�&���I�i6�9%5]m�;D��:;��[�u��vM���g��#������3����>n���3�@�^8k���P�lg�5`���-ϳ��U��<A(>��"�;��z(�()�H�8��
��==�����R���� -��F��,H�a�$]�f� U,�f�uؕˇ���M`�n��:���m��Cf���L�k�qp�=_
�ۺs�Mۢ��j72��#H�����+(�-1]\9%v�6�[��J��g�;r�[��Ns�7C8ݝa%����s!qf��+HYNGL���y�\����9�F�Kšv�*j�1,u ��k��rNM$�4{h���\63�ιN��;��E��V���T�����
?NI$�Z��v��l�@���� �I/ ��s�\��I=��{�H�!X���ؘ�f�^��+ �ٕ�}#�~�9_���U�o��u�6M۱������wfV��Ix�K,�TՉ�ҡ�u��s��$�Հw�~0���=�UU)'��d��ڱP�,v"�n��Ȱ��x�̬��+ �v������w�i���n�O%�t��v�����ź��ni�Iڄ;�{ޒu��tY��η7�_����<ݙXwfW����� �=�V햮�kVkR�rO}���Gɂ@OE��Ux7���;�����/ 6�ں��hwc�I��`ݙX��Xz�ʤ�/�X���Ĵ�Ti_
h.�`H�}�"�7u���r��� �x����f��*5N������,�ܓ�I����{+ �G���%;h����]uU�d�����2�5,�E�[uZ�YM�奬ѤUp���<��Ӡwve`H���W�;<�`��e�`;I�+ wm`ݙY���$w�~0����{~�9IO,v;WBE�ִnI�s���s��빰q��������'Ǟy���rO��훒Og�|	�˚�����>�����נ{/�XvL���X�E�
兢�wc���v8`�s�{�W�o��XV���&U��Cl*�$+�e��{���.7g�3`�-�׉����F`xz�hwbbM]� �d��;.E�un��W>A'�� �K�
�Ҿ�
�`��=U�H�'� �����+?W;�˦һt�%t��f��׀n�?W8�g���o��`vU�@��I��e�w����'���=��vG�qC���0*��`XB�-	�4�H0"��kZX�IP�2�,c$`j8����4j���JHHR�#)4���`"A*�0���)	/E��Sj�~߾����ɐ��bM2�m� �ve`�� �n��7c�h[ �j�j�妓-������)�#�:(M�],�#�kt�X��s��|�N�	_��|����ݗ�n܋ ����5��El�n��wl�f�/=\�$I~��&�e`�"�:�ۡ+�����M��r,{�+UW�_���O^ mE�u�v:��v�V��ٕ�v\� �M���W8�~��	��4�
h-� ���� ݹ��9���U��9?��]��Մ��7X��1�mUu�ó]���NP��:��22!��I�G�g��3^bW66����HR�QX��i�@q�3�UQ2E��kau�a�a)�](��..��`����w�k,=Ე��̛�8�g��nx͓�<7t�K�Ĵ��
�'�9]�Ɓ�1r��ی+]�7pr�f�g�N&q��:ƍ[�u�՘��9}�9��}���:=;v�T��ы����f�����=�Gs�&�=m:�x�vց%�� ݹ���\��Wl'���`���Ё�n݌.��7nE�ou� ���,�\�W?s�Wf���U�VS��P�6��=<�dp�s�ulLۑ`��Yv+���cs���2}s� ݎ��,Q�-�&��J黶]� �M��{�U'���M��wnE���lJ�1*����̼n@v7)=qv�
��L�x�����"�wi"�Qlcv&� ��{{ݹ���^�� ��R�&�nˬ�e���ܓ�3߮�H����h�*sy��w��Ȱ��Xv8g�W?s�v�%_�U�@Z)�m�/~�x��Xv8`��`HL��Ҥ���X�W*�L��O~�v�,�8`�R:.�N����E�X�Ȱr��s��7�~0	�ذ�(��M�e����6�,��JŹ����#�.�@��yH^]��0]B�[�=��Xdp�'ob�r�A%�� ������vq�)�k �~��H����$�y`��g���W9Wg�8��ɻv'Cj�V��_�,v�Xw���U��T�"��1b�"F-�h���Z�P�x���w��ܓ��>����if�Ʊj�������m�,�8`~�9�/k�X+��m�.�ݦ�ـN�ŀ~������{ny`�� >��n��1�����<]�P\rj��jp� �\��q�{�p��ڧiX
���H������N�v8{�ϐz\��;��ĩӰI�i� ���p�&�ŀvG�߹%�����4�P��*t}��M�� ��p�>��x�"�ݠL�vف����X���;�r`��%�ăQh�4H��fG�0�@�E�lN�4q�k ���^�g������{ V�`�rηh.��*=<�˶Sc�]B��.�E��*���ۡ�gϫ��\����7�� ݎe�^�W�7�~0^�]*�0j����]� ݎ�ذ��N��ʪ��U�z�Կ&�n˫wi��`�~��ˑ`�� ݓ+ *E���(�q�m�W��� ����7d�����+��&x�;�	բ��N�!�M�X�ȰUW���~��I����'�g��nI�d��"R �"H��*����6��I�L���2c�����N��GH.�.�*z�E�
O/z�Ɲg����k8,�ᵞ;5��"N���[lJr�n�x�qlۄ�H!^�\l��� ܓ�c�;p�jZ;Qh��|��b�Y��c\�s�ڰ��FK/k����
j^��Z+�.�B7k���g���P�1�Q�1k�������R��S�rNr{��BsW�t�f��-M6�J����D�(�w=C��]8 �݁�b��3��խ؛�,4�n�+ ��e˗������wO{Wv�P��ݺ�&�~�+�I����m�� �L��\��o���m��LN�����	ۑ`��{�����t)��OFeFm�U�v�X�2�	�����ǳ��)WJ�ΆSO�ؕ��M�+ ��a0	ۑ`*����][��J��d��Z�^��$m�2�c����ph۔�2͐_���7Wg�ڷ,��}~:�H�N܋ �&V T�l)U�QBp�f�7$���>�� $�A�|��s�^�W�o�X�{+ ����Ď�ð�]z���ݧm�����L�?UU%��}~�^��,���C��'E��	$��&���;.\����U�~���~��+�v��c�u�Mٕ�~�*����_��{o�X�e`�O�}ߨ,a�1�ͩe��S#���ɭZ&Kt!5���bʽ_�o��7+ʹ������f�;)�)�u�{��w�X�Ȱ	$��W*P��~�����|3*3m*��z�ȳ�q#����I��;� �ն$\`�4�݉[X�e`vea~���]5��H		e2�@�$�N.đ�B�����	�xV na)d^�&��P�awr7���?y��i8�1�b�҄���A�YB!Lsm�a��J�I���".`���HU�!���P�H�5�ܾc���6]ҶBo$���q��NRP������;�Y����<B������j�W5�D�8[-�+��@����ٞ���kA4�fґ�a�����1�S$� CN�\#YH�$�dt��!�-�ಒ�`�[���f�J�e�e0I\S1�p����Z��0���kZH\��F��HѰ�RT�Bm$!�JKi��@��z��iDe"Ȅ�"@$! B1��$X/C0:����hq�#�}@8m�����F�|�޳۹&��X4�Q�nƮ��շX�*��������'���,v�X�e`H�����e$]��;#��W����=�{+ ��+ >�(�'m�-�v:z�XmIv���NM�lA�h�{���q��z���'E��ӡ�;i�X�Ȱ	$��&���s�����m_�������t[k �L��\�$zOe`����	ۑg�H�i=����v!2�v� ����;.\�v�X�e`�p�-�7e0E;n�=K|�~��~��$�f��G�
�*0�E�D��ӓ�����?S��=q�v�W9�;r,I2�	�2�˗/ �ʟ����B�lL�(�InIf�ѫ�ލ��[��I�:ܨ@��6̪���|h����h�݉[]��߲�	�2�˗/ �� M�dM�AwM$շXݙY�H�yߖ�y`I���\����,)Y� [)"����,v�X~�r�����{+ �A2�WR��Rt�m`~�q{_��{���;6e`{��U8�߾�� ��_�����IX���$�+ �ٕ�vGq`ۑ`���9L�	
0	����(!$����i'i��%3�K�k&Fl\��M�6. ��+\����L��=P��s�KGkhT��+�]ЋV�Y�֙+�!簫��l)Ì�Lַp:g�!��<�yçd�:�c����<��A�ڶ_\bӲ�7f�р�
���kM�Aq,������8��1����K�c���j�86v uł����I�M����hܗ�Mί�:�4t۞�4/��T
	��ˢ�Z����j���g�E��I�Ԋ�\�ϜX"��C�*'VX~m��o��lM]Xݺ�w����vGq`ۑ~���e`��2��ڦ�17Xdw���������o���Gkj'bm��h��m�{r,M�X{��%�=��o���թV�������>�%̬n̬�8�;r, ������hcIZ�f7fV�r;�'nE�I�ݕ�v�vI3$��kX���:����nyt�6��z�a���F�u n�Xe�� ��&�{��*����X}�2���J�Rt�n�	�Ꮚ{���@� D�$(V*땼�+y\�I�z`�Xe�� ��R����IX��ـI�ݙXv�%.Gx�p�;]6b`����V6ف�/I� �_�� ����}�s.�&�Wj�M7Xe�� �+�U��x�z?ݙXwi@Ya�^1��ql�1������l<*WG;Z՞[�r�Uq՝���D�l.j�>��� �\0	�2�	��XV���*m;v]�0	5�.�&���'c��	����wQ7n��IZ�f7fV69kʪ���U\�����*���0	���A]K ,j�v� ���N�Mp��\�������wĮ�J�R�v�m`�� �9ʮ{�<|��V�k �mj:&tņY����[sS�ӎ�*1�4��::ܜ�v�����8�:1�@:v�U�	5� �&V�h� �0�eګ�v�ؚ�6ـM�+ �5�M��ឮRGg�Yh�ۡ]�8ݺ�7�~k �0	5� �&V mv����l�WWm�m�lp��}�}��lܟ/P����%m�!"*K�Kb�![i>G��@o��y{�O�JkWZҫEݳ �\0	�e`�ư	�à}�99�y����kDX�P�QNWZFcF�1+3\�P���4�9b�n�Ǆ痢����i5vπ������w�M�f�`B*к�aE!��XV�o �0�c�&ɕ���9ʻ7Ů%�(���ݰ=/�X��`owr���o �D����V&���fǀM�+ ���T���ݖR��n��5i&��&ɕ�ul��nE�6<�W��r�ֈP��j�Y�b�A6;���8��]FcFlI�3�>�θ�<�V��k�nۯa�utrR��xٻu$Y�+�mW6��zͣ�y^6�� � \�[��"tZWX�]4a��9��(������vBy��3uݝX�]D�5pG4�Y����"�$Å^�5p'G ����ۮ:8�`��PҔF�!V��f�P�P�2aDhM�NN{$�<Ҍ�]���K-Z{t�A��f61����3�hIM��[�L�kp�u3s��N.g��o}w@��� 6lx�2�k��vZm;M�m�6�X�c�&ɕ�wnGy�9���l'm�!T���������2���� �r, �֢�Mۤ���J���=U��/���`K���nE�6< �E�]��cT%n���� �0fǀM�+ �\���N:X�a�6̴6��n�'P�n�Ϙ�G1���W��4�Wv�c�֑��lp��6L��do �D���I10t�f l���Wk��}UUU+��W���Xݹ�c��݊�],��݉�I6�6L��r;�ܮr��~�~0{|��L�V�n�����۬�r;�&� ٱ�d���֑'I�RV�vۼlp��$�Xv�w�{�]֧�愪@��R�mR��8Y�cɵ�O����l�kF�iәcXMǫ�:��L�� ��x�e`ۑ�$p��E�ݺ���ISV�$�Xv�w�I0fǗĂ��Wq4Qe5@�����$�eW�������d�� Q�y3Z�!�k�H�VZ�T�'N�6��ʥ�{<`���$�+ ���$�q�n�LL&ـ6<H�ul��G{p.�[j�C/�.])�ָx^��G���r���#��k�=�n[)&xt�]ؚ��m�I��ul��G ٱ�l&mպ�j�a�v� �܎���U�]���� ��<I2��\�������VmWew@��l��	$��;�#���vTE1մ�Uh��`͏ �L��do �HBC��0����$d�I
�=D]
T�����I>���'nĮ��Uj��$�+ ���$��c�:�
F��;*�hI.xwOn5�put��3˸�s�3�Bo��瘷YWE]�>ST
�`[#x�� 6lx�e`{˥s�
�N�m�$p��$�Xv�w�ID�%+M]&�I�`͏ �L��r;�$�kt����:�mZV�����}X����c��IOO<�ǰ�n�ի�n�`ۑ�68`͏ �0UmZ��r�����L�r�9��˄H�с��9�r-OGQ��ɼ�8D� BFdD	Z�
X�P����X@ ZR�)@���P�������1����/4C�\̡��߇�n��E��P�5g'�w�"l2�K�bB�+KRP��\&e��a�t3='��>*h7�׉�o�!�(�°�
f��B]�	�sFk[��v����s��z��湞
��Bf���|7��g�B������1���o�<���J�\&� �c�Ґ仆��o���r7\�����@�IRQe�H�V4�aH��hP�a�B�5��I�ri�{�	4a�g�7w�bD�����-o��`@!$�EB?2�$���C<<��`\a	"1���ʤ�H�Jh-b���f�<u#!$d��� !"!		�K6`�1փ_X�8p�g�M�9�ނ]��hM�J(c�RP���ͧ�#<Cs���.�JM��k+,"CA).�ٔv���r\3鬗Â���-�"��ѫ�\eǓ}[UW����u�u�.�駶#X4�[�ސ��ݗ�� �X%8�kQ�ۋ�5%�cj���S/k�`�l�V���0jD���؜f7l�ս4e`���c*Ԗ�����S
U��z���ɂQ��Qjɶ�c]Z4M�J$М]��&��� �A���pg]��!������қsIGq�ei,�6,+E�Lvba۶�l'0Sr�uh�kj�/j#O%��^.�T�)nCm�<0A�ι+�6ܘ7c	f����b�:�ϭK�;6������.��'Cm�`��r�ꃸ�C�QDת۔�Vٶ8U�/F��C�19�v	�&��CK�<�ص+�`�;���9�h��,��F^-�p(6�v�V�Hv�Z'p��b4`8�`Ћf�+���'��#Z�4�h�L:�p t�N��㘝���,m���e�2*�d�+A���96ݱ��I �^��t�lV�ܼX�DX-�=�˅]��t[w0�b�H۳ m]q�9���6m�B���c�KY0T����G`��]ڮ�LݠgM��2^ծ�tQ�Lg���^��#Y�n�`��(,�ە����c�׷88;Wh���q�r���H�.�{A�8��qۦT�;c;=��-��N�UP�J���B#�[��9��u�����p����t�R�kx����g�����K�d�.���"����ƺD�A�bw�U�F��E���Ej':,5�DA�ը{*���<�v.M��r�^8:�TBq����]6�� �XlRyf�$t�p�g&���d�V-�3��Ì�۴��K{Gc9;/Fv�E:
[R�UVځD�jKn�硺��.��1��<L66����Ƹ��5)��8��,�]s�*���U�#�E�nW��r^�!�S�:ٝt:\6����P�"��50�D�f���e;���vn
pv�;\�96kn�r�]���8D6��Qkuè-t�5��<P�F��x�p�*mUt��D�A�TB�X�ETM"/�C�N��I���I=�䓾~�s�l�5�g�+�C�E�ۢ�t�u�L���F8Խ-狛�_1gŊfӶ�n�;���Gif�h���:�0�],���ω7l���w�p]\p���mn���[Mn�dz�y�B44*�:(�%��,�Ck2��n�m�4�b^s
kk��g�n�8��3-�]DVwA�L����!A��z��d�CS�7B�].��S��s���������]^(��͈f�AW,�)�'#�6dԽp�U�v�[���48ܺ�÷eZuv��m�@�� ٱ�c���W>A���xT��bC[N�+��f l��	�� �܎�	�� 7�V�t��I�Z��	�� �܎�	�� 6lxP�h��S�*�M�V��68`͏�M���$�U�4*.��m�lp��6L��do 7���I���Ƙ�V]RlK���R���ۯ0�]!���v.6��`Ֆ�iun��UN�yl�XV��68`��r��c��e�&��nI��}�h+���]j%�7�vk� l���e�Wv�)�u�ul��c� l��	�e`�t�t;vU�Wi����*SfC 6lx�2���� �l���V[����ـ6<�U#��R+�Q�����i�Kı>�~�m9ı,N���m9ı,Op헧fk2a�3P.�5��lBh�IOA����5vr��z�����%�,�[���_9=���/!�w�6��bX�'�k��m9ı,N���l?,�&D�,K�����"X�%�O�~�L���$0Ԗ捧"X�%����u�ND�,K�w}�ND�,K�߻��"X�%�߻�ND���'��q��qKewy?�Jp�,N���m9ı,K�~�c��O���� ��ț����6��bX�'���m9ı,N�N���.�V�MZ��r%�g�=�CQ5�����"X�%����p�r%�bX����Y��K��L�����m9���/'g�_��C؛gb�U|���X�%�߻�ND�,Kߵ��6��bX�'~��6��bX�%��w[NF�������>-�uu��0m t�`r��]n��ӻ�p�\�"v�jkŲ�*FgD�\��kY�iȖ%�b{���fӑ,K����fӑ,KĿw��iȖ%�bw���ӑ,KĿ�'n�rنW+�����������p�?���,K�����"X�%����p�r%�bX����Y��Kĳ��w�>����L�6����^B�/����r%�bX�����K�C"dO��ߵ�ND�,K�o��r%��%9/�B{>erjaf�{��rQ,K�w�6��bX�'�k��m9ı,N����9İ>�}�} ��9��iȖ%�bS�;:L3��!MInh�r%�bX����Y��Kı;��۴�Kı/����r%�bX�����Kı/��	��uէ��򡀭���2`&��I�.�2�9��� *C���ҼR��2��9ı,N����9ı,K�~�bX�'��xm9ı,Os��Z�'�����/'{/���0�6��x��bX�%��w[ND�,K���6��bX�'��{�m9ı,O��{v�����,O��~i��5��Y&M]k[ND�,K�߿p�r%�bX��{�kiȖ%�b}��۴�Kı/�w��Oo!y�^O����s�Seŕ��ND�,K���m9ı,O��{v��bX�%�~�bX�	�?w���"X�%�t���55���%�ֳZ�m9ı,N����9ı,K���m9ı,N����r%�bX��]�iȖ%�b|/�m�3Z����R�jX�i��D0�T!�����!�����M�������%	�5m���U�Mr�a8�qq�W�^�N���Ɯc�uv��!n�9v�gI�����3v-n��lq��N���ʺ<�"f�]��9�a�E��]. e�]{X{JG>]��Cg�O;��� u~}j��tU�ףK֦]�{í��r��e��B�rL�Jw�]̈́H݈�H1�ny[u�[[g����{Y�q��$:\iTc��2Ř �d���^B���/��~�ӑ,K�����"X�%��u��6��bX�'~�{v��bX�r_|���+�`9����'��NJrX�����Kı=�]�iȖ%�bw�w�iȖ%�b_��u��Kı)�;�L3��!MInh�r%�bX����Y��Kı;��۴�Kı/����r%�bX�����K��﬽����D�]�'�����bw�w�iȖ%�b_��u��Kı;�{�iȖ%�b{���fӑ,K9��e��zQ4mi��'����K��w[ND�,K���ND�,K��{�m9ı,O��}�ND�-�/'�䜓�}��~��fif�85¡Ȱ[nل�����y�ݬ��蹅D��p/�f���[��$ֵ�'�,K���p�r%�bX����Kı>���m9ı,K�~�bX�'�v��
���G3���%9)�NO7�|���mS^4
AV$�:
�
`u<}��K^�M�"X�%�����iȖ%�by߻�iȖ%�b_�}��\�j8��y?�JrS������6��bX�'��ݻND��C"dOw��"X�%��w��kiȖ%�g'������!��.o���B����u�nӑ,K��w�ӑ,K��>�u��"X�%���o�iȖ%�^C��{>���v�r{y�^'���6��bX�'�k��m9ı,O���6��bX�'��ݻND�,�'�}>���60�\6�L��3�� �}�ӧ�.a�q�s�&�\��c���SRۚ6��bX�'�k��m9ı,O���6��bX�'��ݻND�,K���ND�,K����L��Z�L5fkZͧ"X�%���w�ӑ,K��u�nӑ,K��w�ӑ,K��;��[ND�,K��s�fK��պ�R�Fӑ,K��u�nӑ,K��w�ӑ,`�E$*F,F E#���*�ȞD�k��kiȖ%�b~����r%�bX��u���5�fj]j�9ı,O;�y��Kı=����ӑ,K��߻�iȖ%�bw��ǜ��B�������zՌ�䶣��r%�bX��{�kiȖ%�b}����Kı;�}۴�Kı<���ӑ,K������5$�9�cJ�Hm�b{����;+�����XƝh�M�
li�j�[��c�W�O��^B���w�ӑ,K��u�nӑ,K��w�ND�,K��{�m9ı,O����@�� �Y�'�����/���m9lD�wI�$�{��u�BE$O|��&�v%�b_�>/f�f��5sDə��ND�,K���m9ı,O{��Y��Kı>����r%�bX�����r%�bX��>�I��D$���5��Kı=��fӑ,K��߻�iȖ%�bw�o�iȖ%���#Ρ�D�o�ND�,K9<��æ��]hi����9)�NK�~��"X�%����ͧ"X�%��~��"X�%���w�iȖ%�NO�7�}[�5�+"�-	��.J��в\��ѱ�����5	�ʤ��Fۮ�%�V�MK�ND�,K﻾ͧ"X�%��~��"X�%���w�a�y"X�'~��ND�,K���ԓ�h�֮]55��ND�,K���ND�,K���m9ı,O���6��bX�'{��6��bX�'�v���V0�ڎg���B����w���bX�'���ND�,K��}�ND�,K�{�ND�,K��엷dSF�R��y?�JrS���y��өȖ%�b}߷ٴ�Kı=����Kı=ϻ��ӑ,K��>���3PL�g���B������>�ND�,K�{�ND�,K����m9ı,O}�xm9ı,OЉ�v7ѢXX�kh�#h�`�s鋱�1F�d�8ӹݞq=d��ݴ�\�\"����*����q��v�3M�wHI�d�.���cs�����;��l�&�٧s';c�K��7X��D����@���x�:v�����:k�WGbƍ����k����qfR@l.�㵈�g��x���qwRqn�L8!�煞�j�9'?ܜ��.+��O<<�Z��u����欬k�`!�Q�ʰKck������т���6o�'���bX�~���"X�%��}��bX�'���6�'�2%�bw����ND�,K��o�L3񄐺���iȖ%�b{�w;��"X�%����fӑ,K����fӑ,K���w�ӑ?9S"X���)����r�&�\��kiȖ%�bw���6��bX�'���6��c�HdL������Kı>�����r%�bX�t�f�L�]Y�u&��M�"X�%��{�ͧ"X�%��~��"X�%��}��bX�'��}�ND�,K��\��ֵ�kY���Kı=����Kı=ϻ��ӑ,K����iȖ%�b}��iȖ%�b{���t��-�Ҽx��5�w���w=P�q�+vZ��^a@��.Z� �-�V����/!xX�����iȖ%�bw߷ٴ�Kı>�۴�Kı;����r%�g%9/��~v��M@\���9)�bX����m9�� ,"D�x�
�y�,N�]��r%�bX�����r%�bX�����iȟ�2�^B��ԟ@��j���r{y�bX����ӑ,K��w�ӑ,K��>�w[ND�,K���ͧ"X�rS����}��e��vN��K?@ȟ����"X�%��w�~�ӑ,K��o�iȖ%�b}��iȖ%�bS���&�Li�-�ND�,K����m9ı,N���6��bX�'��{v��bX�'}�}�ND�%9)���>�˔6f�Yf��r����gP��)�S` ��x�vb9:�X�v6��$�5r�5��"X�%��~�fӑ,K����nӑ,K��o�iȖ%�b{���ͧ"X�%�߉�w�L�j�[�5.jm9ı,O����9ı,N���6��bX�'�k���r%�bX����m9ı,O����ɜ��)�'�����/'�����ؖ%�b{���ͧ"X�4���~�%}�$��i�Z�	`�II!$�����4�A$$X@&�J����N����O7�]��ʉ���%�MNK�yFa�j��F0I�3�k)�M����َ�Nf�pC�B�H�_<�iF0d�\"e���aI	R��JMR�R�A!���0p B��pnBF	B0��,(T��(B1��!!AwCq�<۪j��ٶ$	�<g�f`K	����"oP�d.l&��D�S4�o-� Z��J%�J> /�.�0M  *Z$B&�lC�O�!���| � �x#�zv&D�z��iȖ%�bw���iȖ%9)��߯���f��2N���,O~�s���Kı;��۴�Kı>�۴�Kı;�wٴ�KNJr{�=��:8�vt�����X�'~�{v��bX�'��{v��bX�'���6��bX�'��s��r%���/!��w�n"r����&,8w���Ϙf�O8�ȃ&�ke�j����a��SV�f��˚�ND�,K�뽻ND�,K��}�ND�,K����l?
$�&D�,N�_�]�"X�%�{��?\����D�r{y�^B����6���9"X�gg�m9ı,N�_�]�"X�%��u�ݧ"X�%�N�ߤ�gu!jKu���Kı=ϻ��ӑ,K����nӑ,K����nӑ,K����fӑ,K���e��fM�u��ӑ,K��w��ӑ,K����nӑ,K��~�fӑ,K� B)�����'U�'w���[ND�,K�O��&L�h��Ѭ�k6��bX�'��{v��bX��#��y�m<�bX�'����[ND�,K�߻���������_��锂$���mX-��K،;N�\.VJ�ɻ8+-�\A�{����EF��"�r{y�^B�}�|�m9ı,Os��u��Kı;�����Kı>�۴�Kı=����ɦ��d�S���%9)�NO7���i�~F9"X���fӑ,K���~�v��bX�'{��6�����y�����H����i�����*X�'���ٴ�Kı>�۴�Kȋ��?~��M�"X�%��w�~ל��B������;��(�����Kı>�۴�Kı;߷ٴ�Kı=ϻ��ӑ,K��w﷜��B����{:|�k3����Kı;߷ٴ�Kı=��;��"X�%����ݧ"X�%��뽻ND�,K�H��Tk`BDVA����h@\~����d�̱2�c���@���c=7M�N^��&�EӻNpK�=�~_w�;o���ĝ��|���8��Ӭ#����X����</$޶紨چ!���yZ�pP�Y�ֻL�%�[�Ò�yL��������������������Y]u�@�1�Qj�
������X�A�*�v�ӕG���*d"q�
a��Zl,وi��rO�w�����P�H�q��ٍ��8�ȴ�&��K�ͅ��i&�ۗS5"k��(,B�;��%�b3�g�[ND�,K��ݻND�,K��{v��bX�'{��6�9)�NJr~����>��7W/y9ı,N�_v�9ı,N�]��r%�bX�����r%�bX��{�����/!y��gп��*T#��r%�bX��۴�Kı;߷ٴ�Kı=��;��"X�%�����9=���/!y?�{�}����k4\ͧ"X�H�����r%�bX�go���r%�bX����r%�bX�����r%�bX����3��Ln5asZ��r%�bX��o{��"X�%����ݧ"X�%�߻�ͧ"X�%����ͧ"X�%�N��e�]�5I�^6kp�X�ru"&x�ĄO��z��9���̈́`��.R�j�+m�r{y�D�;�}۴�Kı;�wٴ�Kı;߷ٰ�)<��,K��~�ӓ����%��߂��(U�����bX�'~��6���(�D7q,L����r%�bX�{���ӑ,K��u�nӑ,Kľ��\�n�vN���%9>���m9ı,O{��siȖ%�bw���iȖ%�bw��iȖ%�bS����u!�-�Z�ND�,�*������ͧ"X�%������9ı,N���m9ı,N���m9ı,O>���޹��F���fӑ,K��u�nӑ,K����iȖ%�bw�o�iȖ%�b{��w[ND���%�ϡ�Ңg���kqӉ�.utm��`f��f�(���В����Kp����V�5�f�ӑ,K���nӑ,K��~�fӑ,K��;~���DȖ%������9ı,O��~��.�ɩ���WZ�ND�,K��}�NC�����,O������Kı?~�]�"X�%��u�ݧ"~D2�NB�w��?OT��i�Xeo���B�,O������Kı;�}۴�K�H�d�B��G��������~�ND�,K�����K����}
�f�w���B��2'�����Kı?}�߮ӑ,K��~�fӑ,K����w6��^B���t;i.�F�v���'���bX��]��r%�bX�����r%�bX��W��ӑ,K��u�nӓ����/'�I�~)��Q�33a�i�8���y�.E�ˑ�=B�=�P��OI9�53�#�2{��y�^B�~����ӑ,K����w6��bX�'{��v��bX�'}�{v��bX�%;'��6>@�I�T�'��NJrS�ϛ�si�~#�2%������9ı,O�k���Kı>����r'�r�D�=��i7�g��dѫ�3Z�r%�bX�����ND�,K���ݧ"X�%��~�fӑ,K��;~�b������)��E#��'���,�������v��bX�'w��"X�%��}~�bX9�C�aVYJZJQh�#��V�\H!rIPq�S~D���v��bX�'N��y��d�ɬ��5u���Kı>����Kı=�W��ӑ,K�����iȖ%�bw��iȖ%�b{߷�2��5��KuSrݮ������aܽY����Z�������"j͉�mI����5K6s=�����/!y>���ٴ�Kı>���r%�bX�����r%�bX�w���r%�bXϵ�}~lt.�X�9=���/!S���ݧ"X�%��{�ͧ"X�%��~��"X�%��u~�m9ı-���wb�i�n��X9<������'}��6��bX�'{�xm9��(�"dO�k��6��bX�'�����JrS�������s�9�d�'��ı,N����r%�bX��_gsiȖ%�bw���iȖ%��	�?}���ND�,K����.�$2�e�ND�,K����m9ı,? ���}�v�D�,K�����Kı>����Kı/䀽B QdP��F$!$H	,{|>|�����͊ݺ��<-���ݺ�Q�$��q�{�/6&zo6��LX��Nmd{L`f�4��5�ËVVK����v)1C� ��ó��3v:l:lw:W�g5j�)��k���;D�]��m�n����nFY�{u�x���j��2�d�T�չ��C�PB��\����d��PA��05�b�_]�VEh���=�cl>J��Ͻ�{�����j�suӞ�g������`.}�k�b���
���)!ͣhPpg�J4i�k=O�X�%���_��iȖ%�bw�}۴�Kı>���� ��&D�,O�j��m9ı,N��Y��.j�]Zhֵ��ND�,K�뽻NC��"dK�����Kı>���ٴ�Kı;�}۴�Kı==�m�̓f]e5�V�WiȖ%�bw�w�ӑ,K����;�ND�,K��ݻND�,K���ݧ"X�%�}���֭�&KsR�f�Fӑ,K����;�ND�,K�߻�ND�,K���ݧ"X�%��~��"X�%��O{:�n`���;�Oo!y�^N���,K����iȖ%�b}߻�iȖ%�b{����ӑ,K���>���Cb*�,5@3A��97���xK�hv�i%�춌!���J��V���k3fӑ,K����iȖ%�b}߻�iȖ%�b{�}�ͧ"X�%��w﷜��B������_���K��r�j�9ı,O��xm9�ǂ8�&�X����6��bX�'���ͧ"X�%�ߵ�nӑ?(S"X��O�ap��&K�0�4m9ı,O�w�siȖ%�b}�����Kı;����r%�bX�����Kı<��Yw��[�j�Yu��r%�bX�����r%�bX��_v�9ı,N����r%�`~T��ӿ��r%�bX��~���5�u�W'���B������v��bX�'{�xm9ı,O{>�6��bX�'s�w6��bX�'�g$����p�"�f��[V�HlJ�g�'����cF7\��[�*�46%�=	k5�V�W��Kı?~��ND�,K�ϻͧ"X�%����͇�`���Ͼy:N@���|Y���b��`�4lI�<�{��q;ı;�}��r%�bX�����r%�bX�������%9>ǟD�F(YY�{�Ȗ%�bw>����Kı;�wٴ�K���D����n&����ND�,K����m9ı,���/�K��M,2���'��NJrX�����r%�bX�����r%�bX��~��iȖ%��@dO��fӓ����/!����[�+6c3�s|��%�bX�����r%�bX~��������,K������r%�bX����m9ı,O~��Z���u�+���#'{����c�0nc��Cj�LV��3�Ci��CY]5*���9)�NJry��u��"X�%����ͧ"X�%�߾�fӑ,K��~�fӑ,K���{K�7��B�2�r{y�^B�w;�siȖ%�bw�ٴ�Kı;߷ٴ�Kı=���kiȟ�W*k�^O�Oǟ�	�k#�y���/������r%�bX�����r%�bX��~�Kı;�����K9�^N���{��a�J1<���,K��}�ND�,K���ֶ��bX�'s�w6��bX�	*��T�"f����Kı/��K��$)ve�ʝ��9)�NJry��;��"X�%����ͧ"X�%��u�nӑ,K��~�fӑ,K�����{*P�Ն�[u���/nWf��-r7,����1sf�"b�����u�ͧ"X�%����ͧ"X�%��u�nӑ,K��~�f���&D�,O���ٴ�Kı=����5��)3Z.����Kı;�wٴ�Kı;�wٴ�Kı=��ͧ"X�%�ߵ�ݧ"X�%�|��L.h�L�jL�kWY���Kı;�wٴ�Kı=��ͧ"X�%�ߵ�ݧ"X�%��{�ͧ"X�%�N����ՙKu2˭M�"X�%��ڿw6��bX�'s��6��bX�'}��6��bX�'~��6��bX�'ݓ�M�;!p�,�˚ֶ��bX�'s��6��bX�'��}�ND�,K�w}�ND�,K����m9ı,O����@�ϡP�*bLD2�^$HČ"$�bE�	e%#B$a� Fb��1d$�����v��<	|��J �#7�Ă��D
xC@��f\P�e  A� ��ߛM3�0�<u���`�5�$�a2E�Ӱ�
(`r�\��Np"�#!%!D�䵄�H@a�F��E�aA�� HF BBF�!v�4JkV3DV��	�"�#�
��OGT��,H0`1�0�JBD�c�� ���0"�$7id���G�b(Mo�\�]�M�F��@ E�2�Fda$^.jKd��`��4��Z��,)�_y�AV�<�v�]�����إcZ0������7��fhq�BOn���s�l�����Du�%�e�U�UH@��{��l��83�=Q���T1�q�8{:u�;���gmÐz���kcc����IF��y'E��_KnN9�X4\s)�qg���P��%�`9B�u�)sB!W�g��O'g�@�+Z��ε-ـ0t�rn�nx�A�T�n�ۇ��`�=�:q�].mZ�{\< <:	�%Jj��q.�jn1�@�h8���w&��e��s%n����,Z�ĭcn1<��jr�`ʂ�i���ş
C��x�m�Ѻ���F�N�t�&��5l�V�=)<��s�X��l󫮂NV���,	�)�Б�$h�AԼE�VZ�mn+;r=��N8)í�Ŗ�wnMѡ᧷��n�1���BbK`�Q �q�9�wqH#�-�dGj���c�1��x_!YW���4�[�gfcs9�ϭ�ܻAt�⮲����7�����n����;80n�ڳ�&�ț�k%%ӞZ]$���F�-c�.�.T���dI+jRXT���Ja���2�U�ۮ�I�i惱2.�q�c<Ѻ�8݌USڌ���b��:�L���Z�lW>�U+����7(]�b��W;Z݌���<�v0"�nK��u�v�2g��4lô>�B�\/;�y�c�>��Q�S�^��ݮ���:Sj���n���:��1�[UG=0j�xx�P�$ݑ.��ګ��\m�D��[��l�+��VՏ`�B["�UuuUV7S�]���K�����UAKJ=�t��7��C���<��}A�������l�;���yP�j����n�uW�^�񫓓��/��)��m&�|0m��*��h��aP�cun��	˞���l�-�7]�;e�����N�wJ���i��y1������n@G�G���;/���r[��Qìv�n|Zs��1l{E��e���.�[r�i�P�p�Z�B����(b�������x �"1�|B���������<�K�'�&���zs�1�+��<
s�l� ܻ���Y��w]�9�0{v�t�*N^�N�T�s�����%!`Tu��p��Դ�)�[��!��C��)�Q��zB�6���fuЬ#���&M�ƻq�T��6�;R���ؚ�vy..��\g��9d�e+*��1��������rEu ֢��f6�X0�J����ؽ�a^.����F{��[�r�s��6`�Vzl��r��۱#)v�`�c��ܟ�!y�^O���v��bX�'~��6��bX�'�����r%�bX�ϻ��r%�bX����=�iFU����^B�����fӑ,K��>�;��"X�%�ߵ�ݧ"X�%��u�nӑ?�TȔ�}�/�c��0�ʝ��9)�NK��s����bX�'~�{v��bX�'��ݻND�,K�w}�ND�,ay��~h�fe���r{y�D�;��۴�Kı=�۴�Kı;�wٴ�Kı=ϯ{��"X��'��}�:8гe�����%8X�'��{v��bX�'~��6��bX�'���u��Kı;��siȖr���w�'Σ�Bk˙�F��I��͎{ֳ��%Su3oY}\�W@'6]Z5�ԙ���֮ӑ,K����fӑ,K��>�u��"X�%��w�ͧ"X�%��u�nӑ,KħI��/n��-���jm9ı,Os��Z�r�@���v�&�X���siȖ%�b{���r%�bX�w���r'�r�D�?~��Y�?j\��&�]kZ�r%�bX�����ND�,K���ݧ"X�%��{�ͧ"X�%�����%9)�NO}��>�&��&�kWiȖ%�b}�}۴�Kı=�wٴ�Kı=ϻ�kiȖ%��dN��]�"X�%�����y��Z-֋.���]�"X�%��{�ͧ"X�%��}{�m9ı,O���6��bX�'��{v��bX�'��>;%ֲ<ܡ�9�+�@!`��)Gv6���E=�8�k�(���"�h���.�ip����D�,Os���iȖ%�b}��۴�Kı=�wٰ���&D�,O�~��{y�^B�N��%�,f��K��ND�,K��ݧ!�DA�DȖ'߿o��r%�bX�~���iȖ%�b{�^�[ND�,K���w$�a�0�fkFkZ�ND�,K��}�ND�,K��}�ND��� �d$�*�hD���@�XD@���Ҩ,M��;~�ӑ,K�����v��bX�%����ɬ�][��lnٜ��R9H�"�=�>T^��&܋ �P"ں���&ZfժG�~��G�/��y��&���֪3@3V���U���t��[��m���^9���Lr.6ug�;��5i6�	�"�;#�68`Z�x�.r�L�M*tն��ឤ�O?���M����cn��V�	�NـvG�Vǀn��0�F1[�C�N�i�`{��[r_�'�����*�9\��s�{9+}�@?��w�u����V��7c����8`[� C���vi��y���M��l���ͬr��$��M�rAmN�Q�C��tg�x���dp�:�n<dp�|��8�r�r�'@��_N��''"F�/� ��y`Mp�
����wZ�5hM�V�ǀIr,=��s�Ļ��`�~0��T0�;�b�մ��"�/ �Glp�:�lx�\��X�t�T��n��p�;#��nǀj�/ �(�W
�QEmֈP��z3��{3��$,�#XWc\!ni��S�o�ϛ��;������٭5s�`ٺq$���CZV[��`�g��8��m���TBzu�[����)h�F�6⹧�i�:�6�l�cq#��`���znK���1��nf��X����&:p�S�ڱ�NSz�[u�-V�լp�`5�12	v�ݹRs���^x��d��ң�x����������b'�4:
1��	Qh�[/�j]&�ڕ[������l�d�bXU��k������:���[%�A���ĶD�M�n��:CM� �I��q")�^���~��ӿI�-��k�u��ft%��6_���L��0�v<庮�;T�t�V�[m`l�Xv8`F��=�r�ű�� '�=hh�N۴�v�u�wc��� �܋ ��}��~��oe�ڍ,����{Y��`����a�ûQ����!{&�۬�m�0�Bj�6`QH��Ȱ	�e`�� �m%MQ�v*MZM��8c�+�H�&V���)ݫR�**ݪCT�ݶ`�e`#��q-Q{� ����wH��*�Bt6�`�� ��#�7c��&V }�)M��T:t��fժG�{�R?y|����;�� 7�N�1�x�ؘ�K����v�I@�m�{u�D�Pd�A�/���7]tX�#_m�cd�l�Xv8z���^^��:���wt�t��e;n�	�e`�� �G�ul���j�v$;jӡ�۬�8`QH��}\+��*�+�pZ�!!$��2�Gԡ�����f+���&V T4U�Yq��wvZl�:���[%��e`�� �j;�[��MZV��d��&V�0�[ }ݥu)2�n�ܫ��1�C�F�[���#7�g]ټ�`z����Jն�လ\�*F*��o��|��0��|�K�����3�ۤ'Cm��0��n��&V }ؔ��cT�t�M6��ke��� �I��M���)ۻ�S�E�R���W9�^��}�ea'�}���U�I ���nϯ ��K�J��vZ��vـ}$��6G�ke�#��Q%�b�t����ۊ8��[�a퉈;1��27]hz�\jŚ�]u6�J��{0��l��L� �h�lUr�`'wI6`�[/ �r,�&V�8g���=�!S��-���j����,�&V�8`Z�<v��|H-ڤ5N��f;&V�8`Qlx�+�Og�kg���e1]�Bt6�`�� �ݸ���}6d�����w���+��ԅ�%�lhle��2�{b����9�e����%�G.� �b@Ϥ����
�VjHV��&�Y��84^�m0c�;'&�դu�����+}=�%vl�5&�����B��P�4�ͻ�����c��Ϧnzۢ���և T%�=6�Th��t��vS�[���Ƙ��*�==�u�>�^� ��gF��c9&D����������\R�+l���*.�V�����\�����s��m�|��f�YV,O7]pZm��S� ݎ�L��8`�v�b)Ӣ�)�x�p�>�e`�� �ݸ�T۔�;��h�V��ٕ�M�V�ǀE�^ }�6Ҍv���@�۬lp�:�n<-���̬ �A#@�t:)��i� �ձ����}$��7�_N�g��~��O�:
�5kL[]@����2����yj��2RC�F ZZ4�.�I�J����`o�ܬ{���w^ݭMR=˶*E�v�o ����T��|PQ�97�5�|��< �#�UW*�6�y+�FSۤ'M[u�zy��>Qlxۑ`�e`I���uut�M� �c�&܋ �I������Dl�e�N��H���"�/ �I��wc�@�|�z�߃�V_e٫]&����Jw$n�����Ύ�\N1/9*^sמ�'#d��;i��7n���X�p�:�lxT���u�.�6X�m��0��< ���e`v*�W�tU��Zl�:����G��>��`� ܰ(D�$��P�S1��� F` �0"˹����䤩(i�ټL'Ml����e��Du9�.�ִq3xȂf-E!"Ә�����m���L��[���nL�*��������I�h0�y�"}�iH���g�j��	B!Fʨ2�rW �%LY$Td����t��2�����&�CF@��m��`��� HA#�jB)J�y�u�U��R�n� @4l�O(�eG�e��̀�8V=%��ϡc$ ZC�����~c� ��p�<�!�A��)�ƍm&�Ớ�J�d�G.d*ɋ����>��;�Z��:D|D_A����%R���TI@	��F1�	 �BB1VD�!	"FBH@�$!�P!��pT� '��o�}�rO>�� ٩!0R���ի��=\J{�x�{+ �0=�r�ŷ�~x��k�i]�T���m��2���uE��d� >��Ա�J�v�T���X�ގB��d�����6x��m���IG���sv��LWn��4۬v8`Qlx�#�9\��=��V�{µ�&��uuh�� �c��<vL�dp�s�F��V�]0�V"�o '��Nɕ�l�Q� J�(�wN�huv���+ �8`Gdy&t!��(��!)as �\�-�%RGP��a��i$�����������K���-��"m�$p�:���I�ɕ�~�����{+6�Hk��Yr��X���	���'cӰ�a�e=�&4I�v^�g��Wv	��5�< �G�w�e{������z�+R-��5e�x6G���U$n��X�?Q�6��ueӺ���m��Xv8`Gdxݑ�����էHN�m���ų�� �o���#�;�2����fSI�:��P�f�vG���ɕ�vG�UU\���'�+T�6ɴҭ��U
��u0mY;�s����,�Mɧn�K`�w���'J��8��U�d'۶�V�p���Og	���S������D���4�xŨ2�4���Q��X(w��a���ii6=�Bl�֌9��O�[�HgwN����^瞞9�x{\�l`��蜻L<BZF�T�61���n^�5��9W3��٭d��4kRY@��"l������.����<q~3�O��vZ�]��PwXR��q�5���F�V���ퟞ�ɕ�wc���#������j��;v�����$�WT� $���J"�&�;��V�۬H�uv\x$� �ve`v��h\��twam�Wv��	$x�fV�8`(�j��V[Rj�� �#�7�2���uM���o}�V�n��!7n7m���C�v϶�t�"U��`Ml ��<v���F�һ���ٕ�wc�ջq�vG�n�-]��)�Mt�Xv8gܪ�	�5
d��!�-�gu�$�{� �ٕ�}%D��SI�:��P�f�67��7fVݎGkiEn�]1�4�xݑ�ve`��uM���[�uv�T6�۶�	�2��p�:����#�>��I>�|�3�1fY��6�g�vЅ�x{�j&C]����Y�]K�]8��N6]��ݻ��_=�� �ݍ��ٳ+ +�aq];��ڢ�0��� l���2��� ����]N]Ӣ�5j�x�G�vl��s���a_XF)HRT#�@��H5|*�=DQ�_}����䜾}���.J��I��5wm��fVݓ+ �ݍ�vG�oM�����ӱ�m�ݓ+ �+�U�'��}�<�fV���&|���t6��+4��&�`R��8�⧔9e�]s��8K�V�N��7n���� vH�͙X�X��6�n�]1�4�x�#�;6e`�e`[�� �+�W.��i�t�6�͙X�XV�o ;$x��m���n��]n���nܗxT��7�ÅT"@d��"!	Ք$�# �TP=9��}7$���0Ȯ��j�X�0	�%��$�M�]�=}:ӟz3�|�0��Nl�	ѵ'���iِ^��z��	 SN1�HyM�+��ut��WI�v��W���$ٕ�nɕꪯ�z_�w�zQ~=e�*�*v�ۼM�XvL�m�w�ul��䓖�x}��M�[�qFUY�<��0	�%�ղ^�fV���&�]Z(n�`�%�ղ^�fVݓ+ 'hڅ�t�n� 6H��2��X��/ �\�B���:Y�(��fPB��1Ά�q�m-ɲH�܎�c��̜����p۵�e�V�sv�ĭ]ԅɖ�xeu*�r���Yq*C!E����GX�,In�F�k ��Yff,Ҽ@�dV���͍c����K�e=E���9}�r���*��S�7��v��w	7l��ֶ2I2K�"�`{�'��g�SwCj�m�ff�m2����������I�97$K�����N%�U2z�Y��m��MX��l�2�p��D�!�k�,�ܴX��T6���;��V6L�v5 M���hQC���*.�`d��7cQ`�$�XZ��u�vYtQv� �� &��	$��&ɕ�IF���"�t��v�k &��	$��&ɕ�M����.
XRE���ݦ��$�+ �ɕ�M�.��#�?W=��~e6�U�J�:��6��v�6ۚ�%��n�A�3p��1���:���V�V{m�w���	�� ����e`vT,YN�*ɥ��S�y�����g9��N[$82� H2H<�	>���� �ﲰ����t"������ ;$x�2���n�R��WjU˺I���Vݷ�l�+ ݎ��/ ;$x6�n��m�n�n��� ݸ����L��t��V��J�)7H.��`��i̢Rw1��F�hY�d��yy�M��5Һeӵj�(M���/ 6H��e`#��6�:����+�ݻN�d� �&V68`��v�b�*�[�ն�	$��&�0�"|��<�5��f��}�[�}6$���ղ�0�۬lp�&�R�l� �L�퐫2��ګe�E4�0	�� �#�$�+ �[~��;���9�xع�%
[d��Tűv;�1Z#��%̡�OC�s�Fƺ|�`	Zw����$�+ �ۊ^ mu��t�Mn��o �L��8`n)x�#�	��
��m�n���M���� �L� ���[Av��I��T��� $���L�����uT,L�R�$F��T̤#IbP�F�)����ܓߤ��L/�%�2��v��� �&V�0�$��y��֣Ř���ՠMˠ�j����[۰��[x�d���r��{;S�p�ݑ�[o �+ ��_�ʪ��=�w��J���
؝��n��p�W9�H��z�g���2���Y�n�ՍZBm��^ wdxd�Xv8`鴢v
��MU�E���#�7�e`��u���P��;��4�����+ ^������I=���I'�{�$��*��TU���*��TU�
���U�"���/�(*���U�� 
�0"�1`���*���U�"���TU�
�� EQW�*���TU� ����U�"����E_E_�b��L���u��]� � ���{λ`����g ���%iZ�5�ً�Q'@5a��UF�Wݸ`d� ���    �( IUP   P       Q���I@ 	�|(�� "�     ;�px}�罜���:��� �e�wo^���0
`�'��(�g�Y���7���2`��=�y���  p    }s�W��/��ʖM9�縕�Vt]��NM}��e�ܝt��
���2�����=^�N�� ���OO{F@vg�{� �zK,��=��������     ��}C&�vuFCy���9��S-��;�W �� �{��+�m�z3�p }/q���9�)�ٜ�#FA�܀� �7gC!��3Ҳ� �    ��l��}�=w03 ���;����m�8 �K�20|���r����ٝ{c�N^������dz=�����     <� y�w7����״/0�� �@N� �:(;�:f �0]����  ��`��s�S 6a���>���f�8�]��s �UK�yT�   �	����2a4j��1�f��ڞ&OR4�T���0   `D�ު�I)24��d@��=��(ȥ   4�@ S�F�)R��      	5L�*�OD��@d`�#�Ow~��㯖9�iӧC�t�ӏMPQni�`�E��E�Ez���g�jHQk�5�/�?��~̷da�1M�
,4��gL�(�⭰���0o�����՞�\$Z����e��t�_��ӧ?�����,H���	��#������U]n�q��ȡu9���bd����@`X=��׼�X�ؕ���\-�|�K:L� ,*ѱ5{$��H���	A^��ϰy�˞Ӧj�YB@:�:��Y���PqW@�od1�B�� ��f�z�o�)�)ͬ}|M`��g����Qq�-���
�2�4�����pe:`T��(}��ݜ]|W�G{���� YQ)����EC*�U��^j �P%��6ƌ��	T4\�,�W�j�p�1*�RǗ��$%1 Pqs0���<��B �Y��$����	��$��]�'{/x�@�)���ۉ��u�|���_#2&ĎݾѰr�`��Z�����s|��B��+Ղ�"w(����Զ��)�*��C% fp&q�b�7i�J�D�BXh�u"��T�uvB�����lu�*8R�Qt(�4#�L���v���e�(ֽ��r17*B�U�l���EƬB�
PȗD�D�z�q�t�h�6*,dA:�E�5�K��ˆJ�\�����F��4Xġ�� ���(�2ۅU��U�*"!BH����U�%D�F7)s;�E����6�q�8�uy!,t*����O,쫃.��ɠ�-))�U���V��0`�W@�B��X2���eQ�n��y�ijB��4���VG�E+![DM,.nh*ۤ1���*[@i"�ʽZ ���H�ʳ4�"�����g���*�r�8�uq϶Y���e`4ܺ����34X%�%�2�W�0�w�"��r0�
�NhI���,��hE�6Ճ{��o[������</\�j(�aBQQ(��*F�Xʃ*2�X ��25P�%%�q(�(��	l	
�d���o�h�S|��r'$�s[��\����(HTr+CY�30D΂��ů�0@����0�G.ܑ�*4U���uc*ZPY�e�Y�"��T*Z# ˔��U�����S$�1*�U���`�:��n�L�tS��������H>�
Em�j5�85̚ldF��4"+R���N��c4*�i�
�Z�j��Xk*�F��T�' �V�,�Y�u1�,��ǟA�����╩�QTD�Di"�]ܧ@T��5\"�ب��	ة 7;.~�I�2�ʢ%:2�(&(QBTa��h^XU��Ǜ��-Q�����@��(�%4A�4TH���#J����(�Qq*)�H��%I`�X�g/E� �u��z6%*�XT�������
��f�f	ҕ���@'2�lL�A�OҮ�4�c��5N��1�ՃQ�^O�z5����j�`�ADh��D�F�ٚ�\��՚����u!S����\��7��H#!Ł�P�`Q,ܳ+�AcW�5>6�s�54�0�?Hja �x&��[�r���EKx�f�\1'gQU9a J3���ٳ�B�dɣf��Ñ*h�`0��@H�FPʀ\B�	 �3��>��
�j��^�0I:�Omk�q�[օ:���qRK���F�@/�6q	@"6(��JXa�P Q�2�%�!@� Vn�"\@1cK�a��0e�j�6`�}*Xц�w�	���������mɭ*2$��0�553[�s��|F��y��J77��`��2�p��%�ɣo4`s���Su��M���Ϲ�j�l�B�f�b%^Aj����y�Y���ī٠�J��&kX �ZJ�q��&�996"d-�I)T��L5�ı;5�$�6�P�tހl �����BP�BU.}�5�/�B*�
LԻ���z�!gh0Z�[�SA&B5 �H,1^j��0-B����{�����$��LBs�-�\3줯���*30�˚�e�h�K�)g/3`�OV
L%�is��P�p���fS.�A������dQ4*�41vE��)�"�"��&Q3&�J�W�
�p...����"b.��P��-���5W񭜫�M��j�*�*��P5@�CY���H��)�n�6�PD�ܦ�m[���&l��eT��E	*��-��ȽE�MI�$#@a׵�ʹ�@br�6E Av��# H[`�u-clE� �*N	� ���&�"Hj4]F ���T����l��h1њ��(B��U%%PdFJ���F�T���w���+VM���U�i����	+R���о��gTG'*�����z6X��B+{�����N��ej�M�2���L-ЂR;(�r05S"}�3E��)�R�.�[�j�PcT�E��ZI�˚�30
��Md���ّ��8QՌ�k&�pddR��b��f��	��j�
;]�>:"d�f�� �O�7��f:d*[��W�	�1�,1*&h �7;Z̓!K
��no)�:"{N٫��6o����u`3T��gi란��mF3,7�S#M�E�ĕ�����o�����F��+�wqYM(����bT�!G�Z3tW/F��UE�9�t����L��8��b�wP�/k������9�`���(�2.�)�@���3�8�!;3l�DcGH�^"��T^H2�hXs�}}�=�ݣ�}��v>��o��YTCj.�!#���_D���:�T�bP�U9�U���;PĘ0�`L���V�{�KB�_���b���%��]��"E:�cs�V��)�Y`�N/6h�N]�s�36�쑃�(���;!��@�1j��:#g.M	K���9VH�F�ŵb�a97B�ح �Dl�h��&U��i(ɳY��.�2��tC��&�()���ܚ��/V�o�j_9��s��1%(^)���x��wr��Z!�f�KVJF��A�>_:!x�%�Ԍ�)"%\j�SEF���m\j����D���J���������*ЖB��0���.�5QJ�J(�" �J#*	W�2����*q*\aB�TJ%�(��Se78��� �%EE�!:wX0hYFf�f�D��%��n�������c��m
J�>01�����(�T�eB�*P4UY�4�T�U��횃2�B�t��� �D�%'j�b����=��S3�B�A%����\��l�>8wm��DE�J���,Jk��kA���e�j�ڕ�awl�B���l�-1�i�ť�j�Y��!g!c����\,�j�x3g�-4汱��.����:��u��i�j�Tb�3YwN�JۓuWF�h�ZDd`�c)ʃVʂ��Vd�*]���FZ)A�^G0� � � ��/41�҈ՙ5,dD2)q�,RR*�K"P�A"W��Q���ȩQ���RD�F20eFD�"A(Ѹ�*7(��R��Z^�rĲ0A�.�Z��0��(j�ʫƬ3Fl��cs�D�3@n!���"M�R���o/�	��U�@��++	�A "IN��$�w�&��
	�V�+F��Y|�eƢV�ʭf�Nώ?D��
�mM�fW(��E�"U���n�"�%7Tq`�`��ғE(��wHc��10�aX),J��.����.�a��"U^k7����I6������Z�)?����,��J����fd�3�w?o��������y�μ    $�  �[h �   l��-�                                              ��                                                                             t                                                                             ��                                        ���Á��a�����Oj<�F����T��	��omڕ�<�E͢�It�`+:ݡ����J�E�Jk����C�p��8��@�:�>�U����/�T*��眜���VT��d. �!b�0�.�z�lf'{���Ohq�V4��gtu=���:b��+�gt'=����2��Va���k1l�0�ꎪm�x�;��K���k�}�}����t`����w(��XKc���\^��ez����0��pv��定� �˱�M�j�:��Ĝ$l`eZ�T�+ahV����v����t��Y.���Z�]N�m�«�)T.��lp�U]V��6����n�ى��n�^8�F���V�V���n�^��]m�ܙǢN�Pۖ�^4�x�&�ީ�/2����˖@ n�-� @�5��MIgnl�Օ���fh���b��ݨ����R��ս:n��V� ���ݫl�`����	u�Yçʻ@�ɲk ��cX%� 6������٫`	-�����isgv�+�0\��YZy%��6�0� �� �ۺcK�VpgE��.Zp�v`*��mR/s\�J7��v�5rKNĦ�zۥ�+�l�&�6G,���m�.݌�6�n�=�ਙ�	@8��i�R�)W#n�9Ƚ�_�%�U!5�C�b��r�ݱ�`Uj�G3���wQ�nQ-]�'��� �cS)!�Y��we`�ۍt�G���"��P��v��.�ݶ�^CZ�J�h�QVqs[z,zkWa}U�^����mqu���p�˵l���GIb���c�6c"=����7�
W��4=��'����+��4yݛ4����inbn�EWaݸ���S1�N8*�)�w=��r6�n�-@�=jj���W��T"�UR�\��<D�K�Kl�6����ۛ*�ag��[]j�S.��%�caF���p;v�îĺ�mMlkvKq�Z���M�ں��i���Ǯyj��-�M�\��0[�r��*�v�L�����v{k��
{@�j��Phm�[p�4^v��շa���lq������\��9�V��c�.�;��fؒs��b���ZM�j�%.�N0��]lj���]�;X}TR�������n&yVc%=�:�͍�5WF��˒����k��g?�w�uUg	\�����=����X�Ay�W�
mMUUUd���t�h����eei�C����lq��U��c�\�oX�.�mWeː�@��j������e�l�<M��v�n=�\S\��NӚ���d
m��
����Sݍ��m���T�Z+�����v�p�P�Y��Ȫfӵb^�6#ug�2����·
m�-��k
�Z�m��lu.s;dwc�cO5/ks���O�K�8��uT�E�� �h��R���vCp@��݆r��8\%T�j	�bv�����Ъ�=�m�lq�T8��ɵ�o�{�����>։\8eܳ�r]�1����]�n�7)3��l��ySĲ�I����@m�6�,k�������8�v�U�@*�5UԮ��s�(�k�n�m]Jn�yg[j@;r����J���h�cR>n���&gv�;���nȴ �\�u� ��X.zl�Q��ڱ�Cc�V�[��r�/�!��h���,]]vBv�Ȫ�檥��Z���[
qJ��/2�yM�t��;Xs�m��Ӗ���8|�ؽ��T��i�tGn5Z7����H�D�	� ��n�A�-M���!ռɞS��v�Wm�ѽya��vg�����N0v[rv��n{g(�F!�t�����T�nwi_:.��1͵���\![u�Z�Y�&��lOEWn�ʱ��٨3�;Hv`�$ަ坍���������6���}�^�j��<ޙؗ�sx�0T��
��L845UTN�X�����[SVQ��d6e�T܅�n�*��^@|�����?�T	Fgvz�����U��H���+�ir�0�5�wt27(��.���Z1n|���s&1UUU)-Ԫ������P�BCw2D�ݻ&��0�f��j�@�#��6�������&��U���
����U]�N�IY��w@$�t5\�hm�Kh-�ж�77@vI�@bF]l�VL���vj�\��-[m,����nX'X5PW-PEi�� ��#�� 7J��Vm((
��l�Ŕ�*��� 8�j�`�Q�Sj���	�M�Nl�  �xĞdF%mU�ʵV�@[���V���m ���q�\����j�^���fKkdq��ՠ���P�UUR�lV�V�UUR�UU��%e�&ݬM`�����tUU��[�(�݃J�� $M]�UU�$6h��ۻD���l���%�hl��� ��L�@n�"��s�v�UUVԪ25�nZ ���r1$�ڥق������
nӰ�,�V���ڕk��ʳ�[�*����8�w6��W6�V���꭫���ͫ�[h��26$�$�mn� $ -�V�즩Ynp&��*��'3hz#S�v��h
��h ��	�.#l��Z�Tv6�ŀJR�v�;;D�ŷP8{m��6�mJ��P�m*�p���њU��ʲ[&�d+�����ʬTZՔ5�6|�0��Ĥn����{vn�#Iģ�ݗfU�S]zy�{E�-�]������)ICmq&�L=@}.���}!5�8��\���y���"G\�m�[�����p�����تǻ �d��;f���T��
W�V݌��=VZ:ꮭ���S\�ld,d��GiUyB� 5(<�����=�N�����e�Hl�ms�ٓ��@UM����@�kv�7w	2�Ċ ��"FAXK&�j���`U�UT05��+][[W]U/+����`�U��F��uJ��2��hKe��(�%ۛEV�n�]��HT����s++�^�I�Qڕh7���+��J�\�u����V�*VV�	l�m� 	����6�@1 [h[���@ 	M$��H[h jM�V��$1! H����@  [r��E����]g��J��]@U -n� [m�7y�ٷ6ĵ@�����Z[r�m�`�m$ X�B��IV�cJ�]n1*��m��V� B�Bb���� @ue��땥�V�g]K�9Mʹ�Ht֛7P�:�S<�T�p�9��v�|�q���oRJ���[�p�y�MÛ���Ͷ�!���Hf�2۫�v�f]�w�Y���Y��! �'�P��-�G��X��W��8�u��S�:�Ի��ՙ(ֆk�I��U�I�Z�SD�����qIj����I�Hd ��$�����e��+`�0mSYj�SEZ�2ЇN�!��VėM!��9EZ���}%l�NO��  M��@�v$��셄	�@�,$�$�I���am+p�S�>\�\¶j}n@����'�4� d j����$�H	&� Xt	����8Tt#�JmJJa�7�H[�r�'J�,e�*1�&�	&�r@�D'd�C��$��|$4'��B��8���X�X�a��e��-iUbW9ʷ�'6(Ы��� q�)��F'�LYXb�E���K  	'>��$��$��$�C��,K$IB����a$��`�@�C����>�FJi)AYITj���R��T$A�X�"��B�
��|$ �2FI���p�%5��'J)��K�-��t,��7';	��H(����b�m�뮋��@1�J�`�'́r�(��E���%�,���0h`0�g&d�g9��9���-�/#h        �              m�              �       $X��&���/��ya�۰���/M�c;vl-��vT���Μx�Y�^��Y�g�Z���8��÷msu�m��j;2c�vn�R6����q۵n��ܯ�E��;�3	�UJ�@�9+eIݽ�q�p孮ϓ��x6�H˱��ٜ��:�x��ݜg:+�]qzLrB9�(�j��Ez�3tl��͐Lٲz��]�i��N��/Vx���g­���[���X�O:ϷM��c�#���wR:��gh�E�Ͳ��z'vny�\��u������q��q)E�qJ��^)���;Z�5�Ƚ���b۷oe�==\�Wv9��v�xv��B}Px����Bn�Jln��5z{+@�ᨸ�y��nx�.E�]-��ej 2N�>r��v*:�;Ʒ\�dzwgs'��{6z-�<��ҽ��ے�E�5ճ�;��Ue�bk[��n��!���zw7]�E��@I��5�'#r�mT�XY�v	YjWC���� YF*%&�9�f6x*�K;"��a@t�����g�&���(���m��;�^w&g��݇���Of�h+�T�s�j[[�ݳ���9ܮ�۝ۢ�z��Y�um�pݹ�fW�ų��k��%�v#[Zq��!�*�Dۮ��2�n7W	�� P�M�#Qڥn�,b�{9B�pj�ƺ�;un����M���6���Njy����ي�fV�4I0���O� ~5I�[�v��9S(��tF�u���%I&@�O�w�effff`��  ��  ������sp�.�Ć��#�m6A��9
%t�n�Ժ�9��	\���C�t��xI����rrW.�2�%5;;�&;n��b��U� ]s�i�3iW����Y#Z�@vN����s�ت'FSu��S�����o!%r�z�w��%U^q��{�a�Mʛ��9y�(pvx�' �-��uLW��^r�ځE{5���e����Rm���~7���o1��q��%�-��)�j���ך⯹��ZJPa�Ԥ���co5�_sx������L6D:]�����R}��\Gz '&̩���U�d�-��э�:�D�����2����2ӊ��.� �5���}ǚ���be'C3P��L�"���	9p��p�=�Mo�ɾ��̣"\D��v�[{�~H�����I�h$�	��T=��*������2�3*\�Rm�⯹��@>�c�5Ǡ����UUXB��gn�/n�=�q7[7Gt,�CӵȪĹA�r\��JfZ�����z�\U�1��AiJd�ڔ���m渫�b��D@#=�8�-�2ٙt=���` [%@�2N�J���s[�i�Х%(�SL�N*������:�\u�jBdJA����@=�c�u�]��=�}��ƬBK�5Y[����dج8�J�.2�IH,4�C��Q����m�b�q:�I&-&�vw?D@E��f��X��3.fT�,��i�_sx�� �������\�.KJY��o�Xg���a�$I��HI�}�����K-�I�]���k���*�f<�<� Mbl��f�vm�i��5��n��Z8)�Q!�$XE ��3-��C�y�_sx���E{y��
RR�%9fe���1W�٬u���<ԄșE����@=�c�u�_s���R�(����� �y���~�.� ����a2�j�gs���.� �5�0s9%-��m��       �̦��5�H2`�t�v}�%�C�+tq�Y����"����ޥ��;�1:�������uM;� �<�F��^;U�[�t�1��k=Uw<�&��)���Ɲ,qcӻ\���6�f�r�������ml�wH��r}��wn�y������Ŵ�������$�V,������U�j���݄�B�ߟ|λ��>��}y�77�IrKd���j���Wo1��qW�c3V�Ҕ�e�)0+����qW��^ /�F�%�f[3.�����/=�*� ����
RR�%9fZqW��� f�ך��/w�M��m���׫5�H����c\t���9��l���9#=�Rsnn�N�o �^�~"���_\�,��j�\�s�E��"B�Jò) D �f}�.ш�Z�UJc��I�M�_fN���{��&�~�<�R���m��y�gsz�w��^s2�eK�ԧ.[� �y��@;��^�q��:K�[Q�e���w��vk�y��{��f�͵�.M�z��kc��u�\ŧ	"R,2��-��jR`Vw1[�⳹�����V�r5�C�}����j�P�X㻨��d�.f[���.�A �@d	�@�L�_�k�}�������&B`�N�g �]�⳹�h�iʔXE&���b�u�gsz�����m�����7[�Q����6�l('X�][�lw���q�u(�ķ-��g��+;�����2�&Qr�$�i�gs��@V{��f�����Ôe�j�� �]�⳹��ZJ[%�jR`Vw1[��y�8Hd	�$a	�wa����k�Y�.������P��_����m��m�]���Ѫ8�7E����V��#�T[��8xV%9s2�Vo1W�
��+�\u��Ȅ2SSt/9W��vk����5�h��-��s��+7���a��ZE&%�m5C{y�f�x���b�9�re.BM6�Vo1��
��3�\h@ w�I~         ە��p��������H��ۚ]سA��:67\�/m�f�-n�Xִ�s�O}���O].�tQ����򷗭ˀ-�%��-Xw`�+�b�^��-�y;65��Żv�tR����Y�C�^.n;]��w7%�VDny�2I��w��Ng�g&7����Ļ���]���t�rv�λYw�]�ȸ盝]6�32�{�W��{5�f���L�R�.[FS�����m���i"X,12�2�oo8���@^{��̝��LJi��qY�co}�gf���+�2R���vj�u�����^d�m��V�k�N-c<^��I��F(P����F�:����E����c75�f�� P������Ԥķ-��o��Ƙ���\�"���؀��b�9�rR	���qY��� *�X��q��:K�[s*S3.�f�*�X��qY���Ԥ�.[FS�����m��~���m���1�ˣ���������[�cp�1x�%�R��z�j!��k��Vo5���_k\fF�(�LJi��qY��� *�X��~�{=�y�%)aKn���{�|?0�dB	};�vn�4#Yf��`��ˠ�UM>��=�J`:��$�#��0��h8��V���:p�Q�+!���p�/��T���5mX4^�1\NO��h�O!L+53&x_�&�X#�Q(3K��/[�hvT��:�$��L8nK��dMwN�1|7ECys����� �Թ�`�$Uue�o2q1l���Qy
6Y���t#
����̼�" �e����5T�������U��k����]�H�����h�"�Ԅ����d�`MB��B@�
�'o�s'9�qZ3Z@���(����V測�c�  /��ztxt�JXM�i�����W�\λ��w�� f��m�mݺ��s<�Ng
��0���[�nF]���r�˪W:�ߙ׸����������.IM��feP��^�ٮ+7���\%�I0\��SK7�j�5�W��W�)^^�@�j!��C��T^oz����?G� A�Ȁ��FC����Hw���8������*��n*�~��@����b�^f/6�m��n���\i�f�;^�7f.-����d6ř�֛?;�d��H��f��5����A�ި�y�i�%M�y��^늼ޡ{�
ӃF̴���m5B��^wP����2�y�I�
ZM8�����Ƴy��s����.I'���{���z��y�s�{D�	]J�ǯE>��ff`        nn��rX�7���r�Ѩ9�N;�`�b���t�q%#�Ȝ\���y3�s��7���8��O�'$�|r�ٸ,ٶ8�ϵ6x�v-n�<^(B��	k ��T��ސCv��7'K;�g\tn�p�JFz�х�H�༘W��O�ٟ��s3�ﾀ��6�Ի+l����F��=z�S�R�vs-��mf��Y��f~w��{稬���� //F��Ia��ɗB�y�^oP��^kwd�@�NJr��qW��/yW��_k��ҹ�%&����{�
��*�\U��E��i�m�FS`^�1� ��Q{���@Uf�m��m�Բ۞�:���]A78�lݮ�738�M8�]Xӛ�-��fw8���܇�"�y�͟	sue�K���ɮs����!'�%B�~�2��]@�;{���
JpQi�� f�3���}�ܸKR�`�-������*��C��07w�ҙa���e���8���܀��c�"/��m�Wtnm�	�${e���s����qظZ ;^�=�NT���qy���@]f�w��x�D ʖ\��:܀��b��^�T^��,�ܕ2�3y���A	�� ��*B�BπIC"\��2+�$�*,� 
�����3�@V��KE0�-6�f{�U���Q�9��nl�K�()p��i�^�xF{���.��>���m��l�˓*�&�n=p<F��ɫ��%�����U���?7}����Ɩ����kk�^wz�{��YIK%�.fX����D	���f��P��= ��8��e2d�3.���w��{���<wd�@�E��-�o��C���7ϰ���C�A�N�$:HG5�t}�q�IM9H��_r/5���({�C�7��Ͷ�m�E&�Gm-�=#R�fy�g�-�i�ٻ�v����I������{�*��B��N��%��	�T/;��/;ޡ���k�>�J	��M8�������b���f���$�d�n�� .�X��c� y���������.\̰2���  fwT^w�B��q���~��/�h         H%���u�����Ct8�@� ,�ac5�{)rv��\cB�2��N�l�N�<�(g�u��Ͱa�Z���F�_m�[���6y�딝�٭��czkz��{9�	U<0�nn�a�v�ч�#78.���Y���1T=j3�s,VK����{ܷ��UU{\���]��y��f:qɒN�]�8��~�+�%��A�-������{�B��Y�qݓ����2&S���}���.�\u���bJi���B��Y�]��������4ڒ�Sq����y���{���=����d�)9*ZmP��8�^oz�{�
�����m�ڐ��夜��.�<^��Iڢ�d�=v	�ĉH�_�Ӗ&�J	��M8����@U��P��8���A6D�i:ݳ_I8P�A�Ͱ�/���*!�
�
�D�c) �T`��c=��=���yxK))4��CJ���nk\�{��,�JW��A̙A�[3.� 3�����^r��y���($���̧���G�7��/���w�u矯� p٬e�mFY�̮9�:�ڸ�3%'%w�%]��bJi��O��3X��D E���ü�4�AL����~�y����/5 �㣸�r
YKuyz=�}�\�{��@�D"B�2 ���$��� �7�}aל�^O�C�2[!&�Lt@�ow�P����: ��Goxx5܉��t/9���=��+3�Q���m��IH��ۨǛ�E��m�n;�.u�	�%߿ww�>��¥��s2���1���7� �����H�"ٙt=���/w�C7���� �t��
�Xnḑ�ޡy�>��DNwy������=-�Ē��E7C�	ϻ�����>���01$���@>	& }Đ浞�S�;�/��S`^�1� > oz�;���@\U�&��̨��6��1�uB�z&��_�}^���E�%�)�2�5����+3z���� $v�����K2��,��m�no�興sy��ǯ5� D��B	�!"�t3y���DD }��/��Cw�Is7wX���U�� ~$������ɯ���> } oz���x��2��3.�ٽ�����	9������Ú��P��<S�h��(�b]�
�nL�����V,DA��)�IAp��Ȋ�F �FQ�I^�NpZ���VH�Tc?U�Rb-�2�)RTs� ^AHA
Q]�,��¬̌`}s(�`%�4 �A,�����8dJ�5p��2\%�j��Il�5[�|��UưkVE�6k��hR�h��#D�Q���`8�����wQ7�C�%Z��L�����#����E�h��$��jD,�{����%mŶ����   ��                                           �]A$��ړ^yz�v��]��{un<h�n۵pBb���y��ܹ�;s�K΃��4\mu��n��ck�ƛ(C�����wR�/a�d��V�v�����*�6��*�К��-+����p�:�譛'7ݹ���7��h�wT��<_V��ڼc�c�u<�l�źB���ɰEφ�YM�K���݆���=/O3�����Vl�7�W�ʹ�1'<h���{0�H�j����'L�n�xn,vN�wJ�uM��#I\�wJ���nz�{l�c�6�lԯgk��yc�%e�����]�`At�M�Ǳ�#n�mF���w��"�n�1�Ź���2���cv�J����q�ºw/�q�`�8�(p^�&ݺ�c	�dx�u7n�F^����*�bm���C=�͍tn�t��*#�ͥ�6�f2�K��6�p�L��E�����9�Ue�ݴ[\ ���)�r��!MKv�kZ�E4�L`�r�����\�[JN9	��bL�prgk�NݮZ �ķ�T^��q���ю�Ȅ�����U�\Y�\Z�>�718�,�o	��6Zk�\�Ж�l���X�Lr�C�]����8�⌾�Q��6�j����h����d����{D@�;�v;[suu�K e�ۭx��\{�,ۭp�K�%Vef��p$>��Bx'd�P��&�]�pv��ا:(�}H$�	 ���WV�j�33        e�]r\��3\�FF�fȯC�l�O��f� ����ۚ�X��6	�۵Xv<nCY0�K��}Z'E�1�y5�I����nڹ<g^t�\nP�'��Cvqκ�&%f� mɤ{r<�u�;�����c�s�ݚqh5LSY˼�����.��ߞ����3�뾻 �7jd�����wZ9���g�x+�cs1�y����b�@��椠T��fL�q�ﾡy���=��=���m$ٖRt/5 ��ǳy�n{�� ���ia������1����G�@s���7��zpn�.AA�*ST8��{���P�� ��76}.Dʖ���M���u  Fo06���渱��Ͷ�m�`�Uv͟FM��:l7n���.��p�.^�߿w�����O�j9E&�f�+5�^k� >�"$g��{�/�Ʈ����ʬ��s$15��
��
��E2��I�PB����;7ޡW����"G���KJe&�n"�7��U nw:=���3|���2M�j�D��S�̧D�@����:7�075��^�/����P�߃��!�C%�@_kL%����P����3v6�m��CDˇ-�.�sѪZ0�#�ìLA�F��{��{���t�d�w�d��ڢI��?� } �߼�`��D')�%ʠ3��W��%��3��oZ|��}n�`h�-�m�$��Ή7��: D�	$�����37ʓ�*\��&[tO� � @[��2O��2M��TN� ��&I�y�K2��ne
$ޠ�r_$�sn�=��/9�l��mշt��8秥�e}�1۫!�:��쯯6G�%o߻��7�f!��n"�3����@^s^������03�� DL9�"] no�x L��0�=��$߳j���>���!�C%�@g�����}������������L�mP~D�$����1_����]�����"!	BI)M��� � ��p�}O�ޙIA�.SB�9�uQ'�  �����'���$�y�N��@j[Z��ȷ\u˴�R:s��/S�ut��k�������o��Ոq۰��/y�f���T纨�����)7D��a� | D�w�d�߽TI7��Dd��~�̥)K[�B�=�a�ksj�DD@�9��@f���=��6�CT���=޺ ��:�a�K���L���"L�iK.fS�I��:$�} o}b���L
��T|��ﱯ���m��l      ����M͸�N�v{f 8�z{��d�uG%j��Y�m\�.�5��gvt�U[��Dy۝:�I�S:�W��5ָ�V#gY0���gr�4�VLk�%َa��v�����Gjc[	�MW�l���]
��5q�i�����&��]�x�ǻ��������d�e��5�.�Ud������v�aq[�n��~��rZ��5��M]�O}�L�i�_�k�/����@��9�2Z�LĶ��i�[�Ty���a� 2rO�ғ,9i4(���U ^w:=����4���y�����q۠��(��y��i�Y�0例�����J K��D���i�� ��3�b�9�z��o>�D���۪���Y�Y$�]$)�rĢ1��E��䱌��o�9���������`gy�nmP���4�����d����5@s��S�؁�TK~�No�d��a� �D �ߗ�ρ3)ʖ\̷D����@^sL�����0/��@z7�ɸ��nZI�'�'7�'s�d��mQ=�3��@��9�2Z�LĶ��i�[�T{���i�w�[m��m�fJ�olJuZf�uI��'y��qq���������0Cb�2�X��P�s�/9�/�_Tg4���"�����q۠�s���  ����I���I��j�" ����
P�!/� �@f��޴��-��%��+0̕�(�[��t���Q$���{y��L�2��O�DO��&�z��w7Ή�� Q��L�|&Ii��pCT�z������No�d��a�hZ�km��wF�����\��M�t�԰]p��R���.؉q0����/9�����P��=�Ĩd6�Ķ��i�D�=��$߷��'s|��"#� ��߇��A�)�D����[�Txo~to�`�i	���˕A�%s����߻�һ�p����I=.{�'w�*.T�ӐԦ�N�����sZ`Wf�����'�Ͷ�n�X*�^ܛ���\�Z��ΠƬ�v�n�������82�������ٵ䒸���w��f�N\DJ�;y��	T�wZU���i]�g�!!�@�{��&fj"\�����sy������2O��2M��L�&ReK.f[�w�Dv��@f�����f�ѽ��5�lp�t�4���.ޥ@_�O|��ԓy��9��=�        
��1C��/8��:��c���-�/<Gh��\�g��9�:��J�/llm�㵝��j�f�q7=�`��4=la��X,��9�0Wf�&��s:�&��bt���G-e�vA��se �q<�5�㋱TN��7���?|�.X_�w��;����U���d���T�/8�@Q�],��0�� �j�4S�Sc�N}�2MnmP��~_+���L7�!9���\���U�� ;{΀��L�i���SC��9�%�@�΀�����Dv�L��P��Jˁ92�� No�2Oo0�5�ڢ � %���@~���@�`��r�!���`{����`��@^sL����m��͕y��\<�G:���<�\�յ.�+�ˮr�B���������@_k^��J�;y��zb9̲!�"����t�B%V�I�&4"ւ �u*P�s�$��$���7�$ߵ�I�ͪ� �>�����jSۢN{�d��a���� ���P�ߝ _.��	��D�6���0/sj�77��_}��F{�0�8��L�Y-&�s��D�@�""{{��9��O|��$���@�ۚ�KI��M&y��tPh�u�s[\p����w{�/�~Л��$������i���y$�J�/��@n��(LS-@�!�t�4��֘MvmQ$��:�"�D@H�����)���~i�{�TJmJ>
�(�����9Xr�pGCS�ҵF��Wۮ��3qH���B���`�H愻�����J�S*�BT���W2A�  �bP�@ʑ�����M���QP��ro����WZ����TT�1!eTK�PĢ����>����Q
�9�A!�P~氺������U��z��3%�H��(i*@F�P�)�(x�Bn@2B�NIP| wp����=�@9 {8jI]����	��0�h�I�������<�7��w����h��5A�%�o��@��@_kL�i�];1�fY����<��=Ԩߘ�w��u$��ϯ@��q��c�-իA�d�F;a�� �����c�|j.nX�`g��f���f��_���7���/��D2\���m�w�`^�� ow�o���$�q�!ʖ��ZM
}ު ��t~K��}3�����0?n�TKD�a��6螁3��:$繆�9��4(�$$�_>ޕ��R��2�B�@_kL$���T{z��|��/���6�m�ӂa
Xp����y�!������ P���뿯w������6�DCX���nmP��~����f��v�&fD�����P��/9�I���@'<�L�%$��.f[�wy���<��Dn�L��P���ܹ2�a'-�'菠[�Xd��0�+�mP��t|�zD�Kn	�m�w�`~��[��`�ߝ}�0?%���|����۠        %�j�Ӹ�q:oX�d�����؅�bc;dscF�Vx��rܽ���M�ɹ�iۃ�8��T]�n��o\vknkvgQ��Ş��ݎ�Yl*р� m8��@�Yb����݁�����=;U�]�yG�ƎA�]�i��������	���wo����~���ؐt:P���Stn�>�vGYe����}�{�����rკr������y����Z`v橢!�P�Ķ��y׾_D�i���0+ٵ]��D��J�P9&Zn�9�a�o5�$Dz 	g��I���@v��9�	dCD5@f�L
�ڠ��A�ћ�L��L�6�P��<�Q��vo�`^kL
��� $卆I�֮�,�L�p�g�{s]����8��h&e�q� ^o:�Z`^k^��P��=�y7p�0ᷥw߰�/@���2�b�	�/� �~���y�i��� ��: �]= �p�&!���i�{�T{�A��t{�d�z7fCI�i��4(� -���3{΀��!�}�I�۾SDCP��9�m�������Z`U��y���˫NEܓw.nMdNX*[ztmS��y^����R�}�9r݁��L�i�w�%poy���1̐K�r�"U��0.�j�/7�}�?%woP�f%�H����U ^o:�&$��&���{�{W�wW}���A1."�Cty�t�4��֘y/�3�t��&��l�p۠/y��Y�J���U ^o�۰���Un��Dv�jN9��71���ku�d�J78y�"�G$6���0*�j�/7����Ho�4�7�ވM�#lK�@^~�/�7���4��֘��4D5	��.[ty���i�I(��i�y�s|�D�B�A�gz�7�`_�j�o����&�k΀�ަ8��pD�7�`y}��v��}I;��$��}� I���r�ˋ��&��X�=��8ۇv'�VG�%o�{���*5�Ղ�Ͷ��Ty���k��|���i�~���A.&�!� ��:�I}�)�y���&�ͪ��	���7,L�l�8m���0/5��ͪ ��tl�)� ��XCmP{�{Ԙ��@��D� �-��$2)��.S�@g��?}��`g�����P@��	@��FD�&��`         �ی�eEX&���7P�Y��p���&��R��-��J���Y�c�%�mz��=�:�W=u�/\�Vُf��orsN=n��~�F�l�[1�٫v��!D�����D�尬���/��[��v[���k����l�vֽ�e�y����9�������%�n�뗴�Nic�.��0�@+���?�w���q!j|��΀�֘���6���P9�A�D�M�&�X~�'7�d���Q�|��}�A��Sq�R���@oy��mP�����w�312�Kfe�'�9���$���o9�O������/)�JML��e�$�����i�y�0/�j����m��m�n=vn:�s�붻7b(睷jq��:�߻��}��"%��p۰3|��Z`W�k��|�} D��|��^�$�����b�9��舀0
���I��tI�������%�!ĹT{�Ty�����#7�03y��6j ��$nn��J#7�:7�0/5��Q~޺$���Is	-7D��a�~ �ޥ@_���/7΀�'���m�(�Ȱ���,�|�����Cj�_Fz�[��u}}@�t1���4��ͪ ��:�Z`n���R�%��I�ު�DL���tI�s�y�>� �7���S)'3,���ү>�J�a��bČ8��(Ɇ�L�1��"#b ��\�$ﻪ�>��x2�3)�!�n����=Ԙ����T{�tI�[�&8��M�D��a�}#;z�;���i�Y�[m��m���4�sc�Nd��rܶ��R�;���IC������6G�\�}ު ��t����֘���L�2�E�m�$���_�����0;�����z ��ʠq���r�=���;�/�IL���P��:$�oSs(',�eɔ(�����Pj�wZU��{4�$� �!PÝ&�=Nfb[D��P��@~��!o���N��'3Xd���m��]Ѻ�jJ���뛬��N�����q2����\�28�"] ^�:�Z`fk^�����3��@z=��ch��Ȇ�t���"&N�0�9��I��:�@d�.�I�L ��T��`^���_|�����4�3Vl	�Y0�K�@f{��/w�{�0���w�0=���!����m������3Z`U�֕���?�npc�FDBt������%K2`�K��Y���E�r5B--̓.��st�ʠJ��fƮ��0*(��iÎ�8QZt4�B��:'�T����DI�J�r��u2A����c@��IP"��������˻[̺��m��V�                                               
�Z��BwM�s�̫��������clF�����93�nt�=u��YM���&�e���q�������2u��n�۰��kdjTl��8�l�_�ۅ:�Lᥠĝq�vFŃ����n���wX؃]�]���y ��yWG'V:�.9�yU�v�r��m�c��ڶ���w���:�e۔ͺ�;�qkX���ϗ=m��];9ӵ�Ns�.�#��C��o\���bK���� ����jv�0��5�lC� ۲X��\���\Zv1��@��nݍ��xrn5���.�cm��^���h0��=r���ڌ+F����n��v�0�۔�4��5��㱑�i��a�g�{b��ƺfЁ�»sp]�Н�-r�}�"� ���*k�w:z��9�J����q�j�����KJ�s�:`�4Fx�!�v'�us1�ڧ�Ev�p�rlh�Tj�6v�۰��ÍS��ASђ^�S4CO컖xz�ىb�D�����Os����h5+�b�uq�)��!E]�9�ѥ�v7+��+��6t����mm�*Uvx��v�-׬.��U�s<;�n74=f��c���Mt����[���nkr�#�z�V��]L4��Itj�,��Ya�ł��u�=2��t��G�]�`۪[d�[sf�v�`)^���$�B	9Æ�C��@�Ѓx�.'3�V�Nr��jV�
Ip��@� o�W��ffff        -�Z��ɩ$M�r���m�������Kf�+��"��m�/Ouv���{l���oc����.6���d�����g���f�m=�����Đl�D�V:NA����΂�N�]������-=��X�l�S�:ܮ�x'&������8�w� M����-�sX�^�9��h��'j�x�WV�IJLzC��Is	1%�f[|I�y�I��&��_�G�����Ή;��Ss)Kr�P���v��y���� >>�~%)�T�fX�N��U ^�:��`fkL��5LD̃LpD�|�Foy��i�y�0例�u��x�m��@^�L�i�W�Ty������m��M��S��붖-�Ss��e4k�tEb�8���ަ�����ڰ7���v��|�$���4�3��@�Y0��.��3z�����D��tI���y�?�OݽN���n%�@��@_sL�����3�T��T>�C��-����Z`]���Q��@g��n%D9N&!���i��;��3{΀��$��_@#)�[��.�.�uo4-��=�c>��O\H��ԓ-9��l&"�3;��/7�}�~_$�\���`g���S1 �n�&��u����2s�a�oy�I���~�(�;�T�Lmse�=���  �@�#�ַ�D���蓺��l���s1�A��oz�3���|��i�^�È.fC�r���=�ћ�v{�0/5�~�m��nN"�txX�v��h��݆ tJ�㇩��6�-H�e�@�΀���ג��uP��P8�`�%�t�4���i�y� ��:����QH�#j���{�G���3��w��h�
���O�"s~��$���o��X,��(%*�AYVx��HD�@�E�W��!���p�.��11����|��i���X�u���ԓ�>�� 8n��V�F�u����e��ṻ==`�����_-֮ڐ&��������Ty���ޑ�0�M)�آNo0�$w}�I��Έ_sL�d71!ĹTguP���Dg��7�`{wiÈ����s۠��/������sz��CL��n���������N���RN��g9�ٿw�        Z+h��x��гN���.���v��hw�zu��A��뭀,gc�sc2�5ɹz�<���G��p��b�z�'f���u�� >p�9��t5���.J��*ܗ9��,k�Φ,v��ri���fv*��݋j��E-��d�{����?/� 1�fNZsw7xL��m�xnڸ�9���vl&8z�)�Q`r�M��0*�j�/7��ߖHo������DC��!�!�sUM��Oj��7��� ��9��>
eL�6L� ���@v���Fl�/:����$�%%32�d�O-�d��0�e窀/7΀ܞ�#桹"!��3y��7��3{΀�ކ�ͦ�n��.��z�����:۝Ѳ�����m���}����I��X����@v��7�d�wu9s)JL"�M�$���b�$�`|Y'8�׷��a��}�$�$}����0�Z%4�w���7����� ^o:{�!�!�P��A�����i���U ^o�@^��z�!��L6D5@^wU���;:|9'~zē��}� I�P˻���]�[��p��;��@F�A�
��.�Ø\��~������Z��y�;�S-1�8s1[t���/�A��0/=�@��^��G�/|�fa�S	6�{�0�5}�-""�"�XE=@�D�"1� �""
� в2�I(�!Y��w��$��:̒S��P~�3}���/y��	�����,�R�ZI�D�y�t��R�3y�_��[�|�m�ڂ�Er�F|Y�xm�Vv�hЃ��r<�b�U�8ӬC%�t�4��֘}�� ��:���9D9NeC�@f�L
�ڠ��@^�O�D��DCS, l�j�����77�{�075�t욤��j!�Q��y����Za�5�11�e4a1V��iP1 ]��$�s�Xe�[��i�D��i��/�䷽j�������݇Ϊ��b��b��������s�'8�v������>9j%���i�W�Ty���;�0�9�Zm�pܪ��Ty���i�y�?�~S'�{��3؇1-� ���@^�L�������T����D�I.[��ޤ���&��TO� 	����'���Ze������0=�f�ـ����i�r-Ř�f����3*���"E1��-v��^f         ��f4�ܖ��������j�賱R��Vm���u[�ە�-�Lm��ێ6�%��n.�6q�4;�����7) `�pA�x}kN�\�ň9tv����:t����ɕ�4tA�(����;Y��q֮J��w�m����M�ww~��9̙�޻� I��ɛsn.�������ኌͶ<��:ID��dLKQ��DCdCZv���y����P���=')"f�r�D� ��:��Qw�`f�L
�mW����4�(n&f\���4��֘~ڠ��@v�􍐘�KS-�@f�L
�ڠ��A�;Ԙv��-�hpܪ��Ty���i�y�N��~ 3Svڙv�R���/b�S^M۵���N$�(��T�����6�s{Έ^�L�i�W�T�Q>!��I9y�Ww�L�9 t���|��� �o��/7ο}w��(�-��5@oy�^�Q��f��@gy��=PCS l�j���U ^o:��a�|���Iϗ��FR�&Zre:$����'�"3ޡD��a�n��D��"7��ꪪ���f�����+E��f�U;y�U��F�eo���%ˉ�-�~i�y�0.�m{7�����dKS-�@f�L�ڠ��@_sL�d!�K`8nU��Ty���_�?%�KjTh��p�S�������(�EF���(�#[&IxȌ�bEh2-[�Ƭ\�nHP��**T-vA��q��� Č�$R(���ꌉPJdH�4QY��W�W�bK�ܣ�,�Q��䭕 �B��i�����DA$������1���
��c����bɻ�%L�%^VZV%��U����R�d��&X5cV9����
4!(��(hh(�#@�+�J�T��cKL2cH�D��2т�
��Q`4X%F�����Ui���Y 2��7�]A�E\�|�j�qWJGJF� dG �F=�a�z��I�ݦЙ���9�m�{��Fo����`VkL
�mP��DD?��%�t�4��֘}�@�΀�'���m�F�U�U�]Z�]��^k�kmb�WD�g�ʕ����7aKj���{�@�΀����AL&�l�j�����/����3���Z`W�d�$LÂ5.�/7�{�0/5�_mP�@����˙n�����ﶨ3>�/R�8J� ~��7�ҽ���cJ�sL6�{�0=��v��:���~�<�޾ ��͌��[�5�At)�;��� �0�b�l�9����r��z������Z`v��r�f�̶������Z`U��y%�A��� b!��I-�@gy�f��(�ǵ@�΀��r�m��&JF��03;��/7΃�(�?��C�RKQP����@_Oϰ�P���A$�I"�"��Ĉ P��[��H��Τ��        #D�f�eɧ\V���@)�\��-��[�0�-��N��;;rnK�{�nv�vL�1v�\F�/:��:5�]R�����dP�v�q�n�t	��9�gk.-Ӓ�����p���qbP"uȻk�����wv���2��6��}�s.s:M�z ��$�zW1�T����˽@���s��9]��csy����Z��|�@^{���{Ǡch�r�e�n�����������s|Әjbe��4��ݪ=�Qo�����+p�B��@�T纨�����Z`tnl8C���f[ty����Y�N��޺�N���7w�����$�[�94Uv�]Z]O!R�r���v:݋�j��^�
�i�W�^�|��7�t��R�j �D�@^�O� !|c��id � �d�X�,j[ "jBkO5��J����+{<07whQMI-D5@^wU ^w:�z���vMRL����A�����2;���֘~ڠ:;��6�2��˙n��ކ��^�*��Ty�tl��m��m)dĶ�N;v^�-�<R�H�2Ia�8�����u��c���L
�ڠ��@\oC ��Ys�ʠ/;��/;�q�
�i�ѹ��b[9�m��s�.7��N�2!� fr��+���i_��taC�6'Km����֘}�@�΀��9DCj!K�P���|��u�o����`TnN��m�{\��K�h{���\[��ZF��KbD6��n�JIj!�������֘Ӳj�fA��K���@\oC�Z`U��z �{ǠRډ�.&\�tGz����Ty����r䘉q@^�L
�ڠ��A��])�������z
�*�% �Ԣ������j�%h�H�5DO5r�'/O3 �-9��(�uP�s�/g�f����/�I����UUHg�hl����e���W�ɚ�=s�V#]�v�In�a�s2۰�y����Z`U�����	�@؜2[n�����ﶨ�֯��h��&	�D��4����*�]{<07whD0�KQP��@�΀�����vv&"IdC��@�΀����ﶨ_%�߷�m��        ��M�j76ؘLst���x�lm[<���i6�\�٫n9%��aS7&�v�{x�n�k�M7��i拁��Wj4j-�y;^�'���]���Z��'3�k&��	�g5\Kvx�^��]�\.�s�sv{f��^;cR�Lf��ww:t 6n�L��$l�2n2Y���Ԏ����]b��dXٔ͵[jӹ'|ē�=cﶨ���1�4����{�0.�j�/;�}�0
�5��.e��@fwU ^w:��`Vk�ӹ�Y2�K��)�D�g7�tC=�����T�D'1bp�m���`VkL�ڠ��@t}� �y3b9���n�w6��5�g��ձ��B㇮uH��Ӂ�ȉT�4��ݪ ��t�4��ݡ�I-D5@^wU}� E��/��'3�d��a�o�����4Ƣ%���/�����������f%��-���`^kL
�ڠ��@dgL�||�%��mP���v�����~��m�U[K���,�y�ۘ�� �l/;Ӷ,?��d��r�\��V�Ty���i�Y�0;wja�LL?�˗@�΀����ﶨ�|�NT@؉"[t�4��֙��@��'����(1VFE!�
����/�:j�3=�@wwR!4��F���Fw�03;��/=΀����"C	%�������@_sI'^zē����'*.͵��nκ�n9p�v9�5��6:�R�p����~�Ӡ/��f�������m-D9���i�/y�g������ ����G̉�L$�I���w�Ty�t�4�+p�B�6@�TguP�s�/����U}�#�
DtD
!޵��n�iK&T�q2�r������Z`]��ku�UUWkOA��n���rn��A��g9!��+�s��!�	"[t�4��֘}�@�΀��BjY08CT�4��ݪ ��t�4��ݡ�H����Ty���i�Y�0+�gTIȆ8"]�������L
�i�w��w�D�%̷@_sL
�i�w�Ty��_ķ~I
$0B��U��-��H��1�Ȝ���I �'.�X�bNa�#���U*�
a��pH��A"$��9wX2�2f7�b�ѡc� �Ȑ��*Q�S1��AaD�E�F,vUf��3 �@E�5��� �����`'��u����Ӳ%;��Y�hd�B�q���A�B��շ,���" Xa.�6o�\��nv�^��"j�j�p7y¤h���q(.���.�]�#�/�!�b�b�﷏�
)CL�I��E��r�
�p�W[������ֵ�0��� \���3��X S@���p��`Td�Rj!@�%TJ��RUP�{��wc��w����HOJ�ښ�                                               	���lՍ�-r[�0��������8��UŞq���á�G��qyw���f��c�#q�j犎�Q�����q��ި�8��O ە���������g��z|�6���q���ٹ�n^���9�n5�t(�vB�=�q���:���1n����epv�1�7k��M[�;mC�9mۑ+�9q\�Ӱcbcvnw�,1ٹ�=�]:���m��vv(�F�Ǳ����5�a�n��l��z�'YwJ����݇h�;ذ�`{]��<����=��P����.��o�����;�s`��7d�K���bTa��k��wa.�wZy <���l�\�\I���l�\Nܫ��
l����$�ۯf6��Oc�TN�:�ўc]]!��n�s���1�.2':c�������ӑK�����h��u���3 dX�ݝ��[" �<��m�3�v�d{ ��[�i^vi��VSt��K�@:��:�c&	8��	�a,N��dƩ��>Lu�b�v��s�Wv��u�r�R�n��1�i1]�Y��:�wl�n-��m�8��8M�깲8ۭ�����(���X*�Lt,pӧ��L]���r���ˮz盂��;�ۈ˄�4�!��sj^^Lj�m�xݴ���vh^P#��mjN����yd:ٷn��d�P7��80ݶ�:6
W��������w�d���t&��d��>�$�B�t*�L�	�U���Gy��9��s�˟fs�s���         �հZ��ke
K��6�j8ϰg�:��;���W�^z|��5q֞2Ƹ�rpO�(�< �P��7A�َ�������{k���.ȷ<�t��!��\�7f�X'��w���}��a����6�ͻ3s��b�̓���w{�{�#着�݂�Nb;�F��.z���p��Z7��
"�3#b��d�2�\�4��ݪ ����;��/��B�n�r��uP�s��f���ͩ�30��q.] ^w: ��`VkL�ڠ75�!�A�d6��3ޖ�4���� ^{���J j\�F�fh�i���3��7�t}����fw��I�$�6��q��g\�OM)�!09쳞�L6D�b!�&�l�j�����/;� ^��*������Cm�C��%�$�{�X� "!�_rd��a�n�j���@�QK	s-��K�Z`]�� ^w:#6Nb���ԓ.h�i�W�Ty�����Vᬄ9�lʠ/;����3}�`ީ'^zē�<_�57m��M�]q�,��
+ۮ�;\UIթ9�#�KaR�K7�m��~�N�/zX�גKꀼ�U��ȆLB��2n�/zX��������ԡCR��f[���/y���i�6A����E�p���w� ^t�7whD0�ԍ�P{��ѻ�] f�΀/�X���vv	�s.f\�.�/;� _t�+5��mT��.�� ���a&����LW7�ԃ㝋X��"fZQp)�A�\�t}���֘}�@�΀�͓�!�m�LKj��柾I$����y��� ��Ys2��r�����G�FG��i��ͩ�30��q.] ^{�n{��k5�L�D1o�(�������d6�q�
�i�w�U$���Τ�y/� 	6lX]�ջ��'�� �uǫ�����R��%ӆҟm�?�Ԙ{�@�΀��������!�3�������֟����C�s2娉t��:���ﶨ���m9pK�n���f����}����67��d1L�&"%�{�0*�j�/;�q�jI�d�{@        ���i��s.'��FX���M��,���C\�gq(n����ø|��r��`�b��N�{Q/����.ѻ����Nr��%�`�nj�t˂ƴ��%���\�P=�q��Ct����{qg!�c��ΜXj�k�d��]9��T 8�&\X���枎����=J ݱ��IC���iZ���X��P�s�.7��Y�0;sj\�&f�eˠ.3�h��`VkL
�گ� ���C&!9p�ۚ#�
�i�W��;����
%���9��/y�^�P�4��07whD0�ԍ�P��@�΀�ކ�=bI��fs��ܞ�����$����q�x��Y���=���np��I+1���l�y����֘}�@twF5y�]�f��}���\ ��b@@T�I	>	!�'f������j�/;���'&C̲b"\P���v���o����0
�'T!��hN%ʠ/=�@�΀�ކf���ͩr���L9�.�/;�q�'^zē��������� n��9l6� Y�n�'U=���;]acc��+b�uG*��q�
�i�W�Ty����P�����c����`U�� ^w:�z���C	%�������M �d����sd��0���OCs�`^���$9�3.\.�/��q�
�i�W�TGq�6����ķ@\oC�Z`U�� _o:�=}@2��6"Ssr[��V��P\ܬ�UN�v9(%\�ܧ$D��/9�^�P��.7��V�'Tf[Bq.Uy�U� 3�X���� vfT���L9�.�/w�q�
�i�w�T��Dt�BmD����`U�L�ڠľ�|�ě��tv�(NA�j%�&(�i�w�T}����`{������[��Sr7.��b��:���gz�Q�a椙�I-D5`f��@�΀�ޟD$�s��\�J2�IKNL�@��@\oC�Z`U����r����ۘ����`U�L
�ڠ��@��2$M�rDK�Fo�0/;��/�΀��Z�cP9�m	ĹTguP��.;��W�0�Z�K�         K�en嚗�N˱@r����e̸�D�l����v�W�6�v�)�g��<�/g��3�l�xn�1q�ܽv^��	����C]���gR���@N�B��*玬T�4��tS݌.Ͷ*�]#�{`�a�H8�6�l�^#>4�Y��90�׻�������UUT�z��ܬ�9ٽ�����#l��Q=��s��T��%�\� �o�q�
�k��}P���{�_�!�i��D���zz���T}����%{��(NBZpD�����{�G(�=�tG��{�!5$���� ��t�t0+q�t���%�3���;y����Ƙ}�@�3<�m��pD6�^���m��Z�]̗�ų�dD��:�U�F��n���n4���� o�΀3�ՔU�u��fV��~��	�$�� s�D&@3M}��J�����z耾�@�Im	ĹTo�T}����`U�L�ژh����Ér�<�����:#�
�i�W�s_DC&�q�m����֘}�@�΀���I�z[m��i�*0u�=��GkgӇ%�1ĸՍvz=s��%�#d��3|��v������`nk߈jRK�e���y����֘ӫS����Z�n�/��q�k�|v���c�F�Z�`w��
L���Ic	}�x:аH�Dj5
��H1�PX�
O���1�a.���e]_c!��"��9�R.`5ueK�m2@5��[���p+�]���j4�L���V�X�X��|wϝ�m����;m�/G/}�g �S(h#�(hF2�&���5*\ahQ*ؖY`T���Н��(N��p(�ET���bo�q�\B��|P'a	p(܆����+�y��Gq��Ķ�ķ@\oC�Z`U�� _o: �އ
$MD�S�P���v��y����[�M��݉W�XW�'��
��wI���=�m����$��Ē��r��z��y���/���&�d��j|���R�4�o�μ�J ��C�`U�j����d����D����`U�L
�ڠ��@owR��l��d��y�0*�j�w߻�]��d�$@D����X�)�T��D<g3Պ��g�X�5$�&Z�3;���g�������W�N�=���p�IvJ��.��;��۶��^�ڗ�(Y��Jی]��ֳt�I;�ߝI;��`U�L�ڠ:;�P6�����t�t?/�Q�4���U _��y$�� 3��a&�a���o�`]����3��@d{��+vcP8��N%ʠ/=�@�΀�ކ^����qȘ��L9�.�/��q�
�i��{�RG<�s���g����        U�o���OYxٷ+^q��#pچ��3G,��ƹ�.ٝ�^����ù:�XG���n(��W�u�c��-۬iٍ�u �֒È�f�&�6�]��.E�+Z�:�j�u�nM�g�.t�m�x6����k�RN��&K��@.���ڭ{�����~~���u�Gpu����'���Q*���ӝK���nfY��tw��W�0*�j�/����J�e�32�3�4��ݪ ��t��075��5$�$�T�uP���Q�0/9�yh�Ԧ�.\̷D� L���D��t�J�i�~ͪ������!�f[�.;a���P����3v6�uV틊�͡�f�vx��άxy���蹈�b9ZNȚ�Z��‼���@�������C ��@�Hc��\�=�U�|�!%�Ԓ����~[�>�tG�
�i����Ș��L9n] _o:�z��6��}%6�Id6���������LٛT���ψNIr9"X�b�����@�ϩ'{ﺒu����w���͆l�V۝�:���h��n����%oߙ��.-��[�6߿���@�΀�݆^����Z�Ķ��D7@�ο/��}�A���i��ͪ� �����I��f[-)M�'c�
�i����G�|� �X
�D��0RDU�� ��\ �y�Q$�Ή&���Cp�R��K�/��Fo�0;7��/�΀�͆[�	Đ�	̹Tf�P��.3a�W�0+1�6�m���ӹ�;VͲȾ�P�v����{iԜ�k��K�(_L6ܺ ��t�l0*��vmP��"J��%��t�t?%�J ��&��TI7��^�'���!��2��LP�i�{�T~�t�l075��5$�$�T��z�=�t�mb� ��	�Օ	6[�"�E
�B�Y���b���|cv��KDK���@\v��Z`_g�u$�˿| '&l����W5��I*��9+��u�bT���p��
1��B�}��?_�m��֘ٵ@�΀/��&��1.(�i�[�T}����`����2�9�*��ު ��ty|�����~�o�`e�8��bdjHpܺ ��΀�Ά^���_}�_������a*[$�Cm����K��f�Ձ���D�o:$��dD�O����        f��ݺ�Y3m�p��19���U��k�C���B�tY�]T�\�Q�g��cdx䵚�n[�+[�-cU�U�[c�r͋�R�n�,+i��0m�l<���:mnM����|��%�C��g���a2� �t�<1e\�gv���{��w{Z�ꪪ��'&�	ԓ�n��
1q�Y�e��=r*�Cc��#fҟ�����][�T����I+���C�� ��a�I�$߷�� D~ H���:$�����֘�ujd�s!,q.�/��q�
�i�]�T��Æ�\L̷@\gC�Z`Wf��3��@=�C�MB�3�y�0/sj�/�~u$�~�RO<��@c�I�:nu�I�Ev,���Z@g��2��RۡŢ�]�������@\vǪ�`n�?H�˖ӢI�o:�� � \vn{��v��I�ͪ�@�'���e��l���۠2=���֘�ڠ��@v��4Kn&(<�f��;z����<��(��C�� ��5$�&Z�3��@�΀��^���K�յ>uUU�=��E�=�7;H4��:��f.�Hq�78z�L�2�"%�{����`U�X�;[�Op��h��nfe� ���4��Ϊ ��u� ��Q�5
\�^V�������ZP��L�h�������`�1��I	��-��z��y����_|��076�D�#RC����y�K�tP��$���z�I;����7x� �J��M��駷�.'O�p��ʫq��g6*��~��z��6��y��ԡCD����y�?� �ު �w�q���/��|��Ԓ�j��w��/��q��i�]:��ɘ%6DK�������޴��I)��?!' ��� b��mo�{�j[M���q��i�}�T}��ݿMT�^lxg�P�����U������c����r�&�G1���0/sj�/����}��d{��gq=q$&�L����P�s�.;a�w�032H�&\C����s�.;a�w�0/�j�����T�I,�-����֘ٵ@�΀��
%��%�&(�i�{�T}����`	')�BSEUDZ'�7ڌ" �`��-I�ƽὃ�2P 貎D XFF"@A"���|��+⤅�KdA��"A� �J$JhFcL���`�a��M#!Vy.�
$$A�H���)�-%F2EA��}�����n�.��`���H�؆�j��F�`��P(�E'$�@^�(�J�R��(��sTFW��:�����#�z���WW	 w8%�*�d�A��D  1�*�����a�H�)��8�țߢU��	�r�Q��"աM�h�3&�d @ևZ3@�\�Gg(֦ݙ�Ƭj�5�]�a5�Z�xJ�v�{���0~۽uն��J                                                	5�D�%��$�F<��kHv�v=��h́׌�[�������l�Q.��K�����?A6�d�^��Gb�4v�oU��(�7%�k���/[b�
�l-�v��`+h#.7p��E�plhc?};}��p����[#E۞��-��V@lA�����lg��z\7����n��g���m�M���R8��8̳z{
a��y������|��<8M���n=�8�C�mn2��ك�-�1،�]�������Gjh�'.X73m����.��U��1����=/l^����nxy����#��p��d��S���ڳ�-ٵع�[Gg�6$�F�;��`���y`���s����헓s9��N����L�Kā���m.37�����ۮj���S8��>0vy��;/�G�m����en�m�g�0����>����]�[&��vϮڲ�0f�[�rs��D��Ij�^�i�QIY[�en�; ��7��kX�$�T��	��v��3���UV-Y�p�Z��Î���e
����&KM!3�eKF�B�h=�S�ű5�;�osr�F��N8v��Ms�U���gVa��.��\=�zJڛ�B��61ɺ�%�:�\�iE�@��k*��Ӕ*^�I;v,%�;=�k]�n�[mAԛ��kg7m���\���I1�m����m���l�l���RKT��"�p�j�Pu�ۉng���#�         �1l�[��n���ve�j[��5�����˫s�J�q'��<���X;
�B��=�[nuq�7.���m�7�z�pJp�j
� ����x��؝�{�5A�軨BP���I�ÑQv�q��3��*�g�v7	�����ww��UUU�2E�
zrt��q=`��<���ă�]��}}�=s�$�_������@\gC�Z`_N��Ĳf	M���������&�6��"&Nx/x���Q��RۢNF�z���T}��_oC�MB�3�����@�΀�Ά{����H�"Z�/���/���|�RN���$��} v\I�����e�xokM;����bk�ێza����S}�/��q��i�]�T澈�.cM�Yy�Wu��l�dH�����#D	���n����TI7��^�2}��(P�)�%�f(�4��ͪ �w:�:z�5,$�$�T��Q$�w:$��K'�'3�2Nyp�-9�	M�������ڈ"��v{�RN����ٌ��Vd�i�Wa����kŵ��y��.�c�cY�m��ԓ�/�$�I�]�^�}�� g��@=ǜ�cR�I�$�s� D &M��Q$�Ή7����|���qs.D�@g��@;���;���N��oy���`�9y.vI��e�i�'�����aL)�>�90�o�ѐ�
aL)���w�m�0�ÿw^���-����Cl)�0��<�4S
O�9��d6S
a������	ϻΠY�&�`j>��m��l4Sp[�=���;�h�.��S��v���qˮu\qv]q�k-�6S
aϽ�!�S���P�
aL)�s��jaL)�0���!�S�赅��ym���S
aL9��z��S
aL+��P�
aL)�>�90�o�ѐ�
aL)�=�;����1���6S
a\�}���S
aL9�y�i�0��|�S
aL7﻽Cl)�0��{�����e&Ԧ��`I���>�90�s�h�i�0���������v@u!7	>��_�w5��W}��e�P�x]��m�0�ß{FCL)�0���ޡ�S{�ޡ�S}�rfl�l�l�y�}�� &D�nn�ոpWm�e훎v
�mhذ��ݤ݆�ߛ�0�Þ﷨m�0�Þ﷨m�0�ßg���S
aL7���i�0�L͚�JL�e9m:�f�`I�=�oP�~-���w?90�s�h�i�0�������w���Ubݹ�7��y�m�0�ßg���S
aL7���i�3�l-�?w��6S
a��~ޡ�Sw��Eae�RV5��aL)�0��ѐ�
aL)���w�m�0�Þ﷨m�0�ßg���S
aL;�u�k���ۼ5��s�����s�����s���
aL)�9�0�T�͞�����        	�6�b~�^��N�<v�iR��ɞ�sF�Y�7��N�OkssS�,�X�]�{<<v�7h�k�&6yn��l�#�07���`�=dRy-gv�76��+���;q M�6�ta�[ldx%a��B��Q�:�݋���	�3<�e1.����$���I@�W�������][d��Hڳ���j��[�H���Ѕ¥b�i���1���?0�=���6S
aϳ�CL)�0��td4S
a�}��aL)�0�~��//)�����5��s���	$e���｣!�S~﷨m�0�ß���a�IuaL+��e��CV�uw���S�����S
aL7߻�Cl)�0���oP�
aL)�>�90�W;��I�m[���P�
aL)�=�oP�
aL)�=�oP�
aL)�>�90������l�`I�&��?Z�JL��9m:�f
aL)�?{��6S
aϳ�CL)�0��td4S
a�}��aL͜͜�3ﺿ�n�"��,����8kg%�<�]���=�`-�]�{�7���0���!�S�2aL)�0߾����s�����{�ך+���5��aL)�0��ѐ�`ЁSc
a����6S
a����aL)�0���!�S��tZ�0m���Cl)�0��}�Cl)�0��}�Cl)���[�����S
aL9��d4S
a��Ӣ�XU9�Vf��S~﷨m�0�ßg���S
aL7���i�0��~���6S
a����^^R�^]U�jaL)�0���!�R{�!*w��d8S
a������s���Cl)�0�w��f`�1`�u&��q�ܹ���[�����t�شG��E]�ո]]�m�0��｣!�S���P�
aL)�=�oA�x��S
a�s��
aL)�}�]yL�輕Y���S~﷨m�0�Þ���m�0�ßg���S
aFgPp(��L	076}jI)2[���桶S{�ޡ�S}�raL�$CD��T �P:0 K>a���0���`I�&��^���Rْ����6S
aϳ�CL)�0��td4S
a�}��aL)�m�߽����S
aL?{��4VyU�8�[�m�0�ß{FCL)�0���ޡ�S{�ޡ�S}�rfl�l�l�w�����"��l�uv�V䔊ѵjh��x�x�V`�틫���w����7��S{�ޡ�S{�ޡ�S}�raL)�0�;�!�S{:t\�+
�1���6S
a�w��6���al)����CL)�0���2aL)�0�﻽Cl)�0��������Zs3)�0$��L���S�2aL)�0߾����s�����Q�u�wCV�uw���� D-����!�S{�ޡ�S~﷨m�0�<I� �A��Pa��k�5�q�i�0�¾�>�#�Q��Y���S{�ޡ�S{�ޡ�S}�raL)�0��`I�&���m��b\ʔ^1�ݧf�E����rg�n(��N��x�x��e���/5��s�����s���
aL)�9�0�o�wz��S
aL;�u�i�n�ʫ����6S
aϳ�CL)�0��td4S
a�}��aL)�0���a�@�P����k�F[v�e5��aL)�0�h�i�0��}���6S
a������s���
aL)�y�tZ�.�-��P�
aL)�=�oP�
aL)�=�oP�
aL)�>�90����a��ِ�
aL)�߳ǅ�r��s��Cl)�0���oP�
aL)?A�w_���S
aL>��2aL)�0�﻽Cl)�0��@���@?t��������fg@       IM����f�d��)��P�kE�U��Q�D]5��-�q�b�v�.�
���<�]mw@�۫+�=�؀N�C9(u�v�坊N:#ڀ뛶��6�[�խ�ŹxٝsԶ�:6.[Ÿ��Gq�3���r3�q���ɦ����q"ޓ1D�/i��w���y�g9��{� NM�Q3sIeI�.��/*3{D�l�82P`�u��fv� ����oq���Sw?90�s��CL)�0���ޡ�S{�ޡ�S
竵�+.�����Cl)�0�}�d4S
a����aL)�0���aL)�0���!�;O{H�f%Vf�)�=�d4�R�{�R���i �9��R��z��7ymeVU��H){�ֈ)���d4�R�s)���rH)�_�̴Ja�N\�B"0/=����9��R{��4�R�{�\�I̙����� I��E�vFH��6�=�ۣ\u��3�\���v�z�����?��3�}�&���C����d4�R�s���uym�h��Xo��CI�I :�I:��㚪ҫ������ ����!����;�R{�-s�ƫ5��=�kD��|��H)s�a �׾�CI!�ץ^^Z9yUYy�
Aa�{�$�9�0��Xk�w!�����9��ވ)��W���CY�WWy�m �>��a ��~�CI!�wU�����
""��Ͷ�m�X��c�4�G',7a\��c PIqvT�����W��)���d4�R�{�R���i �9������^��M�aYU�yz��
C����
Aa�{�$�9�0��Xk�w!���nk�`�I�-ЀH�L�y��  fs@&,ͼE�KJ���f��ֆF`� ��(=;$��egJ��3P���h(H�L�;$@�[��8�UT�"�1�U��8UH��$�c����PǗ���0���Bm ���D@�nPE1�̆�g�$��7���@J~��#���Ү�_n]��H&聽諼Uʸd����I��|��pr�֡2jj��%C*0*!BT�J��d�Y��Е��ɚ%�65�ts�S���d�����;x5f�-SVa�2��F	�,AO�9�d!@�H<�%;��� U�~����K�܀v����` ��c{�XI3�M�vA$: �'} n�2ɇR-%�f1)�X�L�uWIQrI�n�M�C�m�o�d4�R�{�R���¬̺+��6�R}�0��Xk�w!���߾�A`~�@aϿ~�i �=�g��3��n�� ����!����~�AH,7�{!����;�\�I������ 95���nU՝�Z$�uv۪� �RQE���f���NcU���
C�ﵢ
Aa�{�$���0?H$����솒
C�^���/1����� ��?{!����;�R{��4�R�{��UX~����YX�K���桴���a���]��$��w�� ��=솒
A�i��C�Tf8�� ��}��AHo��AH,7�{!����$6N��na	=! &�|0��X{�W�����+*��/P�AHs���R���i �9����^��$���3������ &͙��6�Sk]pݯ'Kgm�8
F�/s�*�D�;7Yf+��w�0�߿d4�R�p�
Aa��w� ;H)~���
Aa�����
��ұ��Ci!���$��) �߻솒
C���h��Xo����AHw�΋Xf����
Aa�w�$���u�
Aa�{�$���0���{yr �D6D:�X�@�Y��R�R���i �7����^��$���^�yy���UU�)���d4�R�p�
Aa�}܆�
C~��� ��Nw�Vߪ�3330   ��  UnmA3v�pX�ۥ������@;mgL�a5�`��;���I[ԯv����kcn��b�á3;i��)]�ѝצ�w����u>�03��7l�kN����Ƕ�T�t��5Ɣ��.NC��МFqY䨫m�.�%��W^�����y��s��k�� b6kj��ط�'�-*Eq\.ǃ2 �@�9#=�3͹;V��w�w�n�ﻆRw��4�R��u�
Aa�{�$����j�2��q��4AH,7��!����{�h��Xo��CI!�w!�!TAa�v�S�k*����߿~ֈ)���d4�R�p�
Aa�}܆�
C�}�*�������R���i �9����^��$����D�ÿwǩpk0�/��6�R}�0��Xk�w!���߻�h��Xo��CS9�g3���� �Ͳ���[��:�L�;$�[v29[�7l\ݑ��}��ݷ����CI!���h��Xo��CI!�w ���:-`�VcU���
C�ﵩ7 �N� jF�;!	pjm ��o�$�>�AH&v�D@$@���&�.e73)Ѐ�罐�AHo��)���rH)���D�����e�x�W�wy�m �9���
Aa��܆�
C~��� ��=솒
A�i��C�UyN5y��)���d4�R��ֈ)���d4�R�p�
Aa��g�~�? ݕ�Sr9S��]�yokKn���zv�����y�*f\�2R�%�r��DD�彩
Aa�{�$�9�0��Xk�w Q	77�e�JS�Ӗ�@$@&���i �9����^��$����D�ÿwǩp��*�Ʋ����{ ����i���葢6\T]I��J�UÖ&߷�Z ��߲H)����[x9W���
Aa�w�$���u�
Aa�{�$���0��Xs�t赃�Y�VjH){�ֈ)?B3�~���AHs�a���_��CI	3���� �ٷ����sq�!�!�OZ��s׋k��d녔�pZ,$�e̦�e:		�y�84�R�p�
Aa�}܆�
C~��� ��=��t^#M���jH)}�0��Xk�w!���߾�AH	�y�8DD}'zd9&J2� ��}��AHo�wZ �罐�AHo��)����OZ.��ʼ�Ci!�w�� ��=솒
C|�A`Q�TB�@T#	0fB��f�r����H�����R�a��r���|��H)s�a �׾�CI��� � �@����m��l4sƟ��i�^��c\DZ��N^��<���т�����Ă��a���]��$��w��~�D��Xs�߲H)}����^U�xh��Xo�}��AHo��AH,7�{!����;�� 
��wǅ�0��j�P�AH}���h��Xo��CI!�w �����H��=�%&�.e73)ЀH��|��H)�a �׾�CI!�}�h��X{���/����Ci!Ͻ�Rw��4�R��ֈ)���d4�R'"=�T����9�2fd��d�dė�       UUY*͸��oR �D\�Ӡ�w,O,STp�׊�x[M��;@��v�,nY�㛶ݺ;k��=]�&�\��=q�v��ix�<
E��{q�3s���%wd;5�nȓ���͎"Nb�@^ݠl��cp���\�t�v#6瓴Vl	�0��ϻ����9���9��/[�`d��ccb�{^�I�nb)�;���- _��S}�v������ ������AHo��AH,7���i �9������^��U٘�yW��m �9�{Z �罐�AHs��)���rH)����ww�7yyY� �罐�AHs��)���rH)s�ֈ)�~�S��^5M�Wz��
CﻆRw��4�R�{�R���i ��>�)��4Rb�D`_��
C��u�
Aa�{�$�9�s$�d���3;�~~~ ���m�q]���;��vq:<��K��=6K��]�v����������h��Xo��CI!�}�Q �����H��=�%&�,�nf[� ��=솓����vPD��,n@(�Hx��C׼0��Xs}�CI!��wZ ���.�Ī/��P�AHs�a���]��$���u�
Aa�{�$����j��Ŷ�0� �߻솒
C}��� ��=솒
C|�AH,>���{E]��7�yz��
C�ﵢ
Aa�{�$���0��g3��~s:�̓9���� ��5�+�&�e�g%Ɩ#\�V�����rqV�.��7��H,7�{!����>�)���rH)��u�
Aa߻���5Y�Ux�^�������)���rH)���D��|��H)��˺��˪�4AH,7��!������Ag�!�$d��Il>�{!����{�Rw��s�1��Ci!�{�� ��=솒
C�}�Q �����H��;��M&Y�����)���d4�R��a �׾�CI!�}�h��X }�z�fffeU�v
�i�M�1q�Wn3q��ukZHZ����u4^%]�U]��Ă����)���rH)���� ��=솒
@މ�R��%�  ��p(��y��D��|��H)s�0�"06���AJ	�S��@�  {}�h��Xo��CI!�}�Q׾���-	IK��i��ϼ���X�T�EU 4=U�uQ.Қ�X%H]$�0J�$���wqݚ:K�[s*S2��@=�c�u�_s;�|� M�.m]K�6N%ú51q�Wl#uCq�qp��2�&JS��&v�{�*��P��{xp&Xl�-��C��� /=�35 ��ǁ��Ri2̴̦⯹��@>�c�u�_q�&D��I��w���z�\U��V	�R�)�FS`W~��=�}�Ͻfkv� ���*"�جs332Ȃ�M/� ���5���_��>�i�5c�7ipv�>ݚ\�׿���e0 T ����D�X¢Z��	���{5e꤄��������ܿ7*�6rky�Ă��,��N�寮o�~�����F>��lǍ���խ?��L�d6j@3��?sfM|
/�]�C��~�{#���Q~v]*����xh����<?�¼q������w�j{�
./ڞ�O���ir�����<�����.U�5��W���y�rq�w>�_F1�4�q�eO���v���Vq�+D)Xa
CV@{��/t���їn4��V���g%�3������$]oJ�e�����_���b��v|��:.wn��{���U�>_��&R
/6M��e�__�_��{��V�Ɣ�l�W��5;O�q_���VgY�s� ���x3��s�e���y�᳏���޲=`�/,�АQ7����|�^�4i��!٬s���h/I���贪
-���c���w_��E���7�Z�r��dl-�Y�/���!�i𴶈(�3���b�(�o���.é}���;�����5_{�����ѣn��{�|	���^�ކ�g�u�=���k� ��ѱ�_O�p�t|�#��L�V���5��z�L�Ŧ}^+د/>�n^�z��6��vD]���67����w����o=��c�'i��W�l��)���^�S�5�j�v��.�}�64wly��-ܝq�H�r���2�>-�cϥ7���)���S�