BZh91AY&SY��� N߀Px��g������`�-à��e
U�	0�f�~T�L�����S�S �M�����@*h0&�# � hɉ�	���0 �`�0��E'����hhdb2 � d �
$l���&	�44M0��h24I��b�MLS�j4Ѡ ��7k�u�� �@L�WH��3��O��"
�aP?�O�*.1�a""�TG�7_��Dc�v���Aρ���"85�kh��?�{�I��� =2$UM.(_
���(�a���fK�Р�!� "䂓�p�t9�0���6�6�3���S=T�)�b~�h���ɿs5�x�84X@W�][�$�E��Y9r��oU5�X�X<�p�_����gN!��xX�r�ě\Mb!ܗ��)���"�������9��}�E]rC�M�g~�1��9{55Z�C��(T��9O�T��D�N�(�A�(y��S�s9�I�� �)�I4�K�v�[j��jvA��8�.�BŃ' *d�E�E�"�I�%���RW��k�r�+m�5�Z����4X�.�5�E���M5�e�Ik�(E�(�d��)ňmas�����D;�ms�S��bBwqR��λ8'�a�ҵ:"�tr�n:<�ܫg��sI�*�jD�d3�+RK[8�[���'+��Cu��MZ)��@�v�fF[��tr����W*nu�Y��C(NF�d��R��Ȋ;�9�)�WӅ^����Nq��tI$��#E���}� �}^C)-�^� �U ��Th�['��B,J�h�DW�	T �\ƽפ.@�>�g](��ϝĆ�[��`0�>b���u#��
�k��r��X~��Q5z!0�,q�F��'���W5�Վ0����;M��!T��׎K:E�ˊ3�@wD���w�������<MpJOȮZ�GS�!�����;e����	.<,����~�4�APP�<��gR�:Ч�,l���K�l���_$��U��̈�8u�p��lj���1I~�=F�Q ��#-�dc�k��L�:F���ų_kn����B�C��z�E�m��J���&_Q�$oف�� O��]�Ҳ6S~�
:5���AEu�x��-�,��O3����R������8��?e05P�d}����ܮ�0��m��&2".�(Vu��B�i-$3]��96q�&K�źT7L�PF������Ҥ�oA/1���HN`?�=Ӈ���ڞ�yk�m�u�6����s1){U�dߐ<H#�t��ln{�w��b�P]�^BYaǌ����בe,��UD=&��d��j)���Kә����F;�G/)�eE���8��+�m70�B$؏1+���A$Q����d�c�ƃ�|�O���(h?N����@uQ�2��ܑN$:��� 