BZh91AY&SY�s��ß߀pp��b� ����a^��`h%� 2I$�       @ �       ��y(  �     D!     R)J�@��(���EB� �@ 
8  1�
�)T
��@���O�Žrj�,��}�)�� �oZ\XSݝW�{=Q� �r2z��� !����  6`�A����
���Z����ͩ@b ��3B�    �� �@�(  F��� 	ﯖ\۬�m+����\� z����Z�Y}�^��x�r�� 7*w��+�ݼ5��ʹ��� �RŽ�9e�\ڥc��������n.��;�uun.���ڸ�} )D�*I   @ >��W6�����Թe׭��{�V� ��՗]W+�r�ͥ}9r��}n�[{۩z��w���ݫ��U�x �J���[��t�ʾ��ޕp n��x�:��������/]�ޕx� �$ PJ� 
2 {�_NZu.M}z�uNMR� ;�,�r���W6]z�>�/�� ]����5<��  ��ӫnMr�� �J��ϼz����}�O^�p u,Z�ɯ^�^U�}��_ .�� ($ (Pq ���㻬��on��]nmڳ� f�ɥ2�\����o�p �{��]��{�W�/  ���o�{� =�K�z���������'�{���R���w��M�4��w:o�     	D=D�y�R�=2���4�@h�hb~�hE?�	��U &�L &aǪ�JS�L � 4� D�*�)�%F�d14�� 2O�$2�*��4�   ����U&&)����h  z�i�O��?��?����?��p���_}���EEW����ETUv��*����*�舨��@�DTUo��`�����̿�U]�ǺTUo����o�����R�3/���������h�����<5&u8�?Y��xǚѰ�N��-��>�~ݿ ۸{u7}Ƿ;�=7]�c��)�����w9\<����|es�p��y�捶�ŻF��,��# ���cV\�$q��(H41�	C�hy&&lJqr�Ő�8:\���a��L,,<��o�p��&���ܰ"��f<��4��ֵ�3+�.^�q��ax��x�֏7�[֨����0��j+4<��$�~���2	�A�w���	BP���dc��v6G��h#'a�$��'P��8Fj���0�5AkP���h�:�ܙ�z���V�U����(���P4蠦q��8YĤ�9Z���9�5��s|��A�kF�����ԖP�I�F�4D�FF8��kO������_��_0��r���*��*�%��]����T�\���%v�5�Ӂ�S���5��7�(�u��k=�wٞ�n��7ݸ�}�7���껏v3۶�8�9�^��Z�Ni�0�hJ�2qh�4�ّ��I������Ñ���wl����!�5�0�f8����t�8�!��� �4KF��D��(j��4~�F�޷��7���he�X�f���,�������a���)$%�l5hĞkD8%`��%b�F:e��d%	��B��&!P�a����8霒58kS�}��5BV�%�t�A�P��L���`h��M�Da5I$b�a)6�5Kp'*����>W���J0�Q_9��6�]�ϻȸ}>v���*���tvs�(篂p�yy�\5�5����$����X'�v�Є������4�e}X�\U��Y��ϲ��P|�⺟]�un�$�\��>���>)η�ӲԞ&qч����A��p,��*Ōt��{�k#1�R��$E��D�}�+�C�)S��m�|�YχTY
�<����:w�\�J[-^��,�y�2�֊[F�r�5���O�~��m��N���rq##{�ϕ2����j��H�
��sݡ��*���N"TD�>��t�I�Pٚh-ic0ċ'2Lc-�ы�:H�0r�`�4j�iq�t��c��12��� ����)0١��I�U����!)q�%!�bk4Ð�2qrt�5&&ZM���-!��bO�����r�i+hd8���L,8�%��i5�88������I��nC9�$3 �Y�'c�Bs4%�#a�J1�sp�����2�k����8���m�%���q�A���Ø%	BRbj0�
�*M���%:v��iۨJ�ӨJC7��,Bn��ւ%ƍBRI����7���3S&�jC2t�8ubA��.�K�@h�Jt��x�p�t����L4�d�C'K���=�N'O$���6��Q��!33V�vZ]i6��l ͜3Fא�f���M�qֳHe�Y,j��&�Y&�j�kL<���Y���`�r�߰�ٸ���Dr��Lǖ,d���F��nI�6pL�(p3�) ����c�F�2�F��ĩ�'�ZuC��`�)0�,�C�&�'%Ӑ�2Cz�c!)�֝�#�ܒQ���Á	�4�@a�sZ��[5�+I8�֒�[9gY�fB\�.N6��4e�:��"���ӎkX����d�-�Y���f��)�#���58�9	�}7��#��w��_�,C0s[<�H�[���H�������>PG�9I�e�1'�[9i߳���O٣x�kB|f#�I5�̢s4Q���?N盏�����~�x~_��c��q�LM�ag��#N���$�I��m�[8d��;��y��7�����9ʜ�B�]Uv��S���2����,H2ă'$�Þ~�7��ay���[u&1�?KQ�֣���!��c,)��ڌLM����p��xp0����	-A�����d�:?A��	���~���hقq+�!���X���Q��{.¸Mc�5HfL�^�>#z7�������;��k,�U�x:�:�]j\=�%���T���S�Ɂ���5	hJq�jLM��ۃ�8bb�P�e�P�Ě�	Z���h``Ѱ�{8��ylJ�J4��0	s!(Nf.���(JD�Xh��	�JWc������!BP�B{���r�X��$1���#7n'a>k6Ó�5j�������O9	K��lὓ��k�h0�%�ن��1���	OR�<�u�Q�9&-fL�x��?[ϱ�������Z�����e���BD�a�9�/������6�:OO'ѳ��S�)`$�5����~���y�xPH���!����=�� �����d!F�bi2�^�A��^^j�������d��%'�fF�n4d�sA�r�m5&��7�|<�I���	Hk$Ѿk~{��s���Lw�;H�Ų���/3/Cc���e'�L���M泿w�V}ˎ,���&%2G�`�B���4'�h<RI�bL�i� � 0�'��L'�Mrp����&�-	�#���܄��������m�x~�{!���c���^���ԡ���Y��dm8��Pl~�4�O�G�p?F�~�������/����m��'$<Հs�1>�a�0F���M�~�4O��.�с�0�l:�۝$~�������>�N���4����sZ��# ްtA�ǻ��~Y�6���Gޚ	���߁�BL����O�*����)�N��J�g�l�TgW�afn���X�kI��򍙹��6F�&�N�&,��HAL����Li(��.9BR��49&%��L� 0���S����c!`����������J���)J4F8��IS��	HfA��&Y�.BP�d8�!�`�ZI[$e�nBF�0�?~��f�I�%	FP���%$�A�,80I�`��Jq# ��8?������4��BX:�4c�t�`Bo1�8l�N��r��ې�9��%ӑ�2�c	I..o0J 0��I����jtoq�L��K�v�ƝlJBX%	F�I��L��LL��A���:�4������xoBS�w��x�5f�����xi�a�z�M6���ٺ�`�N�Nh�P8��h-?�49��'���٬����fF�F���%Æ� ��j5��/������.Nk1�k��É��f��� �i�ְ�G���l��l����a�kHe�p�`	BPk[�����(y��9���4l7�f�|1�j��F̓ZC2�s��i3I��ǐ2K�FkNT�U]EyS�J�)����ة�9uL�����,5웵��]D�I$.��2\r���# �4ề�)�X�����XN:6s=��hߛ缣��?����}�NA��lJ���d%b;2t�5��X�F�S��6<���e���&0i����i��\1�A���$�|'!Cǚ�Z3K-$!&X�O��F���i�!8j0�A��P�u���������Z� ��I�1[C0�[3���p6p��v�pR�3w�� ���#K�A���x�z���֧!4��y���yn3��-�a���_6hq#	Ǒ��c0,�Әh'4٬��̃WV���0�Jq�#�?1������	�8�h�Ǉ0�Vk�Y��<mZ6���\r����-f}( 0JB
Y1
�
M&K�I	��b�W��f`��� �Ʉ�0�l����8�4��FL`h�h6�5��sfkz��ϴbqi!�,>�ٸ0��B$b����ӳD��Q�CNP���l׿�5�5�6q�BS.�&C�7��2�i����I0������l۩�F�Y &��		��q�C2\і8��A��K��êY�S��J�\ �2#0J1ѿ�&����_�X�Fs��I����^��8~��20U#�]2��x�>󴫞�_�˨X��Z���Z޳�ֵy��X�?3�^-��?ި�❋y�W���U5�������e   �JR����` J4��m��l�֖���C�� �]h��ņ�ӫ�Wf|���n�+u��;^�t�-�vz�6v�:��J�ٶ$	�����j��mGm[^'[�,��vєW:�m�����/Ke-��  6��� �j�  $�� ����d��Hr��n�-��-��  �  l���b۶�p:� ���  �     ��6�#� H��6�lڶ���   8� 8    � m� [\���Xim �( x�$h�8m+�7m�ض�$  �e�Ā!mH   �� �ڳlֵ��B�	�mqmH VԦݰp6ض��m	     [@8Hm���l����kn��U�@  N8  �m����]�m�ٵW,8���b���v�Δ�	�����A6�� <m�ۦ�6�!�� �@�  -����oU��jB�CZݶ��H  �`�-�j�oV�p 6�  �� � I�� �m�8 [[l�$� m���-�L�`  [@ h  �� pY�  ��[BF�  6�g6�ݤ�Z���-��@ �qm��m"� l,� m������B�rN�kֹ�V�[@������� ��l[B�Ԏh  $  -�hA� @ p $m p  8 H!    [@�[C�	m��n�l. m�  u�[{~��ρm   �nHn�m�m ��H[\5��m�@��EӶ ��ᶶ�� 2m�Iź�m h�m$[rm�   ��      �6�-�     ���  $   �m  �-��6�� @�   �lm������@6ٶͶ��ci6H    6� 4PCm� ��@�� � �m���s��n�(���[vض��0�̖N��uql�Kkm�mml  �$l �6�   �mm�  �i�	�-� E  � �$  � �������m$ *�)U@�W��km"�6�8���!m 6ؐ�>mm�� �`7m��-�IQGJ�[;+@HMt�5آ�XH�V��*�U@R�++lն��]�v�n����W���mW�$� �hp�L���p@   �E��m� �g� �i� $l�UUU�F�  +[�[��UU��@Mێ3�@B^9݈�� ���)������G*lM.:�+nċh,���gF��I-hm��@�`K([\ m� ����� �}EmB����  ��9� �, ���kskZ8���H�#��t��Hp-�km��8m��HkY;k��[m�Z� ��e�	I.�� H	l  �l-��&� a�H�[N��S�u�	 �HÀ$6݀�l� l	 8@ -�A�m�  l   4� �	$6�f��I��ke0h��   ��[ն�m�8   m&v�+j�p	l��q�� ��9!��m�8i0��$ 6�ڶ 6� $,� Ѷ�m  m���9�8	   ��gJ�� �$d8 &�@ �K��  rC���lI ����m��[@ 8 6� H m� [�� �� ��ݷ�8 ��n�@�m    ���-��m��6��>��ޓ6��ڪ�[p8t�[@  6ض��Ā |km��[p ���9�   Z7Mm�%�t 	R��6[�E��`s���WT	�O.�mU��mH ���v��[v,��j��Ƚ�� yӦ��-T�(>�V��{����f�u��ﾎ�����
�U[h��0 ,K�^m�ާro	�7T.n�;@U[Z�	UIU٪���ږ�@NT��� �8M�-�������Z��[�UTl�� m��n��	�ݹvv�<�9bʯ0msmW�&նH�� 6�imm&5�  �HR���mk  �� 8��_Bێ	��Ҁ��[Cu����$�h ll�   ���   �Ͷ k�6�'$  l�4P$6�/Z�   -�[@qi��J��Uhf�)j�}�@J�    6�	�  � 	 �� ��-m�[\u�  ���m��[V�  � ppѶ� �a��A��r�l�"�[��m��y�UJ�lWJ�1O)F����� �m e� H l�h�  �    h �� -�  ��   >�� [@  -�mHm�d��  ��� ��	  p   q��h   ��m�^��c���X��/  U*�YM����W��8m:I�Y�hs��[h�`�lݰ H �Hm��m�$� �  -���� �  l 	 6-s���6۰ n�M�� ���b��6�����j��]e���� �  ۶�` Wd(�\bU���a��� Hu����kd�*�!v�hm��񸡕��Y���w�� 6�i6pi%�&Ҥ� �N�Ė��l�VK�˜,5��85��βX)�n�エs�J�*�#(9%�JX�J�D/]�,��V[u�� m�����pn�P�#�-��X;ns3�%]���ꅹ�6�"u h  	���m�UR�q�; F�Ť疭�8��=����Km�1�F��А$䀗�WU@K�A�*�^P�صnͫc� �h�7Zh�l��UW8�* 6���Im
�j@ �����8K�V��@ ղY��P��� �5�^�p��[F�v��m$[@$�`I�Ƚi��T� ����| m��H  [�� �ki�jBv�ت4uB�e�U� 6� $	 � �I���)Cm�ۀ m�l�m�q%� #N����n�ꪀ\_mkm	>��  $  �   m�۶׭ ��CA�W:*�c� *��i6Zl  �Im��$�P ׶�lB��	� մ  mm�l��I6�J�ks�n����+�4������V��   6�@�m�  �l m��  l �`   m  h ��H  	�@���$ ��h��   m �i6 p��YYV��¿}U\�t�4��J��H�C� ��<�Z8-� ��,b�n�,�p ���l q, �X��V��� TX��m��n�&���k�� mm	 p����Ŵ�M�$"I�t�]��l�N�&l6� 	z�m���m�   � ���g� ඀ ��8 	Cm��m�$  Hl6�   p	 �  ��m	     m� [Kh   q� ����6��n �  6�۵l[@m�.�  �l8�B�j   $ m�h $��_Z p�m䞶Je���n��-�e�lඃ�� %y�`��۠�*�&�ۓ�ݪ�u H�� �σm&�ml [@   m�  -�    6ض�$ imm� �o��[@h h��A"G�H �� 6�-���� � h    ���  -���[p�m�� I� ]$ؒA�� m�n�jH�J�
�j�8�nvRN�@sm�Y�U�`��-��	 �h  ��p$  m��l   �h $$� lpH �m � /^��D�H��ٶ ��l�Z�-��J��a�m�W[KN̴  ��~�m�۾ 6ہ���ޭ�� �h���ċ�  ��m��6��mpm�}���V�0 YKKn� �J    mְ-�6��   �u�&Ô��P
�m�]$�[J���ƻ&��KL�U�kL�����`��@N?���-�����_�
**����UEW\�����������4�>����EFS�� ��=?�W���/�@��T6����Ԟ��P��D�
�PM��� �ਐx���t���Av����~� �>���� � ������0U|<��Q}�������?�����<y慐����� M��'�q=A�o���,����| Q8*�,	�4�B���+�3i�$x;S` ?����'��UO��P�O�E\�"q}!��� J�A~W�0�$"���?"�M���ӈ��!�*hGE���T�4+��}D�߄�0Dy��
��6��E4	�6��,��^
�x�?��m��HO��������y�?�����������	"�m������ǽ�������M���:��Ҏ49\Dnɷ1��ɞ�y��]5��,Ԛ�1�Ў��[8K;s�� �,
�U����`8^Ӭ1EWUF�zm�ͪ�ij�
�6�vQ�Mu����}I�'T����ź��WBq�O�mu�n�v�*�� 3��a�`�nN�8]YCb˶}������R�I.�Uuv��,����]+���M.҉��	���;N�ۀ(&Y�c���4=��N��[Y��k�J�tѭ-R��+���)s��k�e�A���T�-͐ 1��<�+J]��������^z�	�%�Z��ta����NO7!��<�����SXS�VU۱F�����m79���[�a�4�V�ɳ���UUA��j����lSF�\
�z�2��N�:/���W[���/; +/0UtqUm�R�9����i��6���;ioT��t�5R�����uN+@4'@s,!�*�ugrcC�'vܴ���M��l��g��V�MHn�ݑ�l�V:)*s!��)�������m��.����A�m6+l�ܼ	_I�a��U��Ť�;�
܉ڶ$$8-��sVƪ�:[(s9��@]N$��ۇ5bȺ�X-�bgtmP;����6�d��I�I�$�řhr�[����v�۝`��G���u�n,��ٶ���F�Vѩ J�t�t<��qI�p˱hB��]:F��!+u��B�L@R�i�c\j���US��q$t�Գi\�H�}:]Ij8\�2[�T�]�	�=�vvT�;M�mA�A���І�Fƹ�O+��*Ý�V�TQ[R]�8� : 8uEICbg��Hj�2C�5t��No*��R�� v�<I��NV�	�r�7.�N
ݙI�VXZ�)�T��75#���t���������A�8ӵ�����9�}OI�s$m�;��m�azɦM�OX�$��4��^�:��l�nK��4�:Cb���%����	L=�kv���f��\�T��xB槃�� O�����Sa\�GB2���7�ճ[�k[�h�v�<'8�uA2�:'t���ٸ78���@KT�;24�\wnۖt���L��x,=p���l���':���ݝњ�@w^|^9��;���n�sҽp��5��j6
P���`4]��OGn��4���4c��vq�mÝ��GlZ�)����j�uIU�T۰l��;:�筹Z^�."{o,k��t{��{��绞����������\+�v\��*�vrq��Ǳ�`��9^RmS)6SM�-�C����`r>��_��wgwg���(n�J��m&4�(�,.���RA�͖|�U��������&�q(�#n; ^�x���Z0�r�ގ��Ԣ�$m����}0�3��X]�v��K��e*-�DB4ӑȬ�`>J�{���r� ��*�z�#^�n�+c\]>��ݓ�4�v�ZS�+��)��]��Fхjj��g�V �ܫ �����h�;ág�m��H�]�;��_}� D���� 窈���Fz�K�酁����:uy#TI*q�4�v{�;酛Ij��5{5�z�"�m$IQ$7;�O��O�V �� ��)YpSm&4�(�,]�v.��������a`�dj9J�)#aN4��*m�������Wh�#����u�xsL�g���a�̉6��(⃑���v{�;酁�����|�Ԣ�$m���]֌{��%X�%X�""d�f訶)(�M:����ɥ�����G��)�U�/u� ��FD�Bm��Is������za`g�0���Ϣ�q�����`	u� ^�F �r� �t����Y��6��ɗ�ٍ)J�;U� >�ɰ�x:��yæ�Ŭ����2a~�%֌{��ʰ>�XޘR���IE*4��`g}0��Hչ�����`fza`�6d%�6�r���ʰ>�X]h��р)\C�D�MĔqA��]�;=酁��w����G��AҢm=U��x��~��TD������L,�`
|�`
}ʰQԬ.��.j�؛�nVX�C�kk(o39%��f��QJt�.�N)�ۦ���*!ER1T�w�O��O��wZ0pB_dL\�MƤ��}�����`g}0�3ޘXL�g�i��#q�����`�р)�*�=� �"�R�Q��q�m}�R�e�`nd����c�1w1�:��
�4�%F��,���fvgwS���Q�M�g�� ^/�!�A��h1օ�C��8��6d9��{ewn�j��[8�ncsոKFͲ�"�j. �V�Ѧ:f݁J �yd��֖̼;v,�M	�y��wly�iO������Y]vɷ$[�PM;M�̮�� X�m���y��m��0 l�c������;lO ��n7kbs���%�qe�j6��=����4�[�W�l���+*5Q�W��L�9�U5�'�t�t�v6�0���w�>�K�ٺv!��j�G6�r�![���k{붷.�l�֫���ֶ��+pM��?���*��р.�F �qO*JM��Q���v.�;;酁������c�=�}p
��Q�uu�/u� ]�# S� S� ��T��Jt�2I=캰1w1������|��Ҩ�ۄ�9uq�)�U�)�U�.�F ��F������wf��\�k�%+����ʧ��-I�4F۪�0���ز���Ѳ�����<�`�р.呀)�U�;�THC��i���������q>k���������ʾ�َ�;�F`TI��*4��`g��V�%X�%X�`e��КrD���6��k��5{u��L,����Ş)�II�܍������ q��,f��y�%X.��?M�nx�B�G���e�vfA�'�a�c��Q���ps�E�ՠ��R$�u�{��pܲ0�%X�%X�*0WO�%
U$�X�e���UUW�$u{u��������f}t�$�PnBG*���c�1w1ٵ�ʪ���_R���`nf�X����聴���� ��V�W)�r��6|�`�@���u7�޿b�3�˫�������`s3�BDRR�)�'[��:�ns�z�9U�z��R�O&���i�C�Aj���5"�3�˫�������`w�ج<y�A�#HM�7wϒ� ^J�z�N ��F:��H���%(�rI$m'�o�f�W)�r��6|�`СeL�5*!INK�~�`g��Vs�� �, z���s[�|�񞢱]/��)Td�E`g��Vs�gs%�޿b�3�4fTD�!GF[�m4�uV��y2X!:��'S�k#�^i�wA�	��"���nRrU����`��`w�ج����<w�eD��e�]� /%x�ﾈ�;�9�O# ��c���YED�N���q���,w,�g�V ��V {�Au-T�Ҧ�V{�u`qw1�w2X��+ �u��ct�%$�����3����_��=�O��x��5)ɝ��8���0	��&��f<2On�S�ҺK`G�"�Emi��-8�Z1��۶�8\і%��[$a-���w��͠� AڬV�����Љ�OfCv+knҽ���尬�� J�m�D�Ŷig�5vS�W`Y_&,����ݽ��2kH&��axH<\�<(���n�'.tQs������;e�gǠ6��ǲ��L�#r���>�����Pp�FD7j
N��+Pgh�qaƵ�\pr���s��j���u�ċU2�~}����W����=�W��]{Օ��J�R	'!��w�d.�q�%�/%dyA*'뙛"���!w+��y,�y+�w�dwA	I�	5�䪾�2���O��{.���U�^��d@�i�D俳����}��}�{�����U}�e�w�K#i��*!��})-slg�:g����Xn�u��9���]�]�V0B��E'EJi���=��{%U���_}U�ܭ=���yQ����%MIu��J�T��0L���<�Ͼ�þ��9�e���:�mQ1�r��U_|�B<�}�ܲr����q7SUwe]�SW��%_n�,�ܮ#=�;�|�ə�b�I���j���吻��g��B<�|�+��{R�q&ܔ08I&�{�-��+�.
��4ܛ�H������ܗ�E�]�^�I�F{�d#�W۽�#�JJ� �Q��NJ��s.��c�����=�]��S�)�i����?��{.}!� b�9G�A+�#��B�N��5杈�3�%R������(iQ��l��@� J��P��O�)��~Ar ��	0��M(��+��E$C`���Ɨ��P^3�t�#��S�����)?}���|��/�s��:F�#4F�f��qJ�����JS�}�R����{����s��\R�����{Nf�Z7��5�s�%)N��xqJR��}�x>JR��~)C���w��)�*>��Z�/6��v\T.tf���x2Y����#vm��'�㭷=s���s=p��9Y��{�)I����p|��;���┥����%)N��xqJR��{������f��l��f���|��;���┥����%)N��xqJR��{�x>JS�fV��E
�Bc�R;���������|��;����)JO=����)Jw=�u�)JO�#���3q�z��s���)Jw�ÊR��{߻��R��{��P�@���ם������g�݁ݱ�r��[��&I�L�ԥ)I���%(		�w`�����W�g}������YLM��O�� P�9(8��vv�ݚ�lVC�n��E����Kf��kYk[�y���JS�����(~���|��;����)<�����){{�fY�7��6k5��R�?�}�x>JR����R��{�{��R��{�u�)J�^�w�e�,ѽ�9����)Jw߻�)JRy���JS�����(~���|��.����k,�kXkZލ�{┥'����|��;���qJR�����JS���qJR��{����f�����5�5���JS�����(~���|��;����)<�����)�>����ֵ�����/m9�#����x�ֻ+1v6�X��n�'	��;6P��3e�O:#��;x�4�M�%45��Fݕ{l�`�l(5Z6]�3�����mV�-=�e�r
��d<x�Y���`��U�-����k	׶���M��A�X�y���j�.l<�s��;"�5[�p"�y�`�T��uul�����6�zs{��wm�n2�ۻ����=��>�u@#7��3�&&E�y��z�<��y8���SYE(^ȷ=D���0��W������{���R��w��)<�����)����R��􏳦;��ڭ��9�s��)�~�)JRy���JS�����(~���|��=>;܎j�Y��7�Z��)JRy���JS�����(~���|��{����)JO~��Dtռ�k-kyo5��|��;���┥��}�/���~��8�I���%)K���2Α����Y�o\R�������R��	�����������%)N�w\F���ܣE�d$�"�N2$���(Y��T1uË�s�� �m%Y�p����ctֵo{�kz�8>JR=���┥'����|�)N�w\�@e�J}�������}���ћֵ��f��Z��)JP{�{��:	!�����qJR������R��w��F%)?g����rH')4���>�������R���~��匔����8�(�f�S=���ɕG�b ���������k�R�?�{��|��;����)JO߽�x>@�s߻�)JRx{�>Θ�37�-��9���-)�~�)JR~��{�<��;���qJR���{�)�)�g�_����Z7���[�2����v.�hmod�Jw6�T!-����ƛ�Mі��ճzٽf���)JC�~����)J]����
߾��%)N��xp���>��tG�f�Y���[߃�R������ )J߾��%)N��xqJR��}�x>JR�׸}��-�kYe�ֵ��JR�����J�}�R��jh���;����߻��JR����}��ޭj����o\��JS�}�R����{�����{��JR�����J�{�t�m&Ԓ�%_�P}���{v��JP�($�����┥������)߾�)JR���ټ�l�3y�K̆]v���7<2��훣ˮSu�uq��3�������]\Hա�F�w����o%������)C��{��4�~��8�)I���%iO�:n��df[�Y��Y�o{┥���x>JR����┥'����|��.���R��􏳦;����z�����Jw�ÊR����{��R���{�)JP������)��ޙpѺ�Z٭��k{8�)I���%)K���┥����|��ꞩ�$�w�~8�)I�5hW�d�M�IDRK��}��Q�ݜR����{��4�~��8�)I�nm��>����bߛ�ԃ�q�D"]yHcK�=J.�P�&�l�.X����88zt<���X["�fk0͙�k{┥����|��;����)JO}����)@��v_�P}�}�m���ȕ�%�}�߾�)JR{�~��JR����)C����%)N�{��f�޵���o7Z��)JR{�~��JR����)C����%)N��xqJR��{pfԔ�N29������P}�����)C��{����~��8�	�@���c��$��;�����މ����JR�����%)N��xqJR��}�x>JR�}�w�)JOG�Xg���]idOV�n�v�臵k�<�lh7l�F���G[���v�T�!Qg8ӎKj���&Ʋ!e#v=H�`�L;b��}�[f*rMZgM,WK�y��c7#��۵�q�:����e�3�[�ۮ��㵴����L:��n�����q���ӫpH��^��#�`M�zwN�32v��q\��7ʥ��A�E��
J��ԁ7着�j}Ww�`���n���q2Ʋ�s�Mo��Ib�u�z!T�/e����f\��.= X�y���)O��ÊR����{��R���{�)JP������)��ޙsU��Z٭��k{8�)I���%)K���┥���x>JR����┥'ﯳ�:j�V��ku�����R���{�)JP������)߾�)JR{���JR����Dn�՛�fkZ���)C��{����~��8�)I���%)K���┥�m�JHD��.��}A�չ�ujR����{��R���{�)JP����}��>����R4�%*4�'P,�^-���&�%[\�v����kpۈ�ur�^�d��m��$C���>�����6��%)w��|R����{����~��8�)I����{3z�n��7�7��|��.���~�)�����?�(~���x>JR������)=��w��)�ƺ�v�3-�7�ݽ�7��JR�����%)N��xqJ�X������R�������)<?t���;��ݛ�����p|��;����)JOw��|��.���R�>�����)Jz�v�
蔓�N'%_�P}����o�J�s�����J������R��w��)=���p�kfo[�5�5���)��"�Wl�qh�xܨ�i����;ѵŖ�$¥2R��N�E$����P}����)J߾�x>JR����┥'}�ۯ�}��Q�ʌ5T�m��┥���x>G�)���qJR������)J]���R�>��`=��MIM�ܒ����}[��W��)I���$1_@$?
�7)w]���)C��{����p��Wue�kY��7�Z��)JR{���JR����)C��{����~��8�)I�����,�[��������)w��|R�������JS�}�R����{��������]�f�33as��S���{�4��
���l�`B�v���r=hM����}�v��m����x>JR����┥'����|��.��w�)JOzG���fn٣\��p|��;����)JO}����)J]���R�?�w���)Jz}�l,�n�5�ݬ����┥'����|��.��w�)������>JR��w���)?}}�Q�V��hټ����R������(~�{��R��w��6	����$�?/@�_���ۯ��g�݄݁l0����A9�k3Z���)J߻��|��?� �����)>��������~���-ս�F�)� )DQ��$��[��^��Z[iӖ&�vE%�4u��7����I��ټ�of�k�������}��8�)I���%)K����ZR�����%�U��!F�m)RU���P}^�����J]���R�?�w���)Jw߻Ê4�'���Wwl���,���-o|%)K����JR����� B��w��)=�����)�ڻZEI�p�'%���UPW����}�)߾�)JR{���J%�z�����0�	����U>���R���w��)��{�����{��JR�����%)M*"}pH�="Y��
JKs(7����F`h^��c8���ky����ap�(	�	�ff��1a�h���Ė+XdR�NIfH�"�fI�A�1
Bтd��-b$���X64RUba�RPME&&�% feB��֤�
p��<��UQfE���f�3	��S�e����,qM��(JX�rT-������`�$.by�'%�vD!�a��6��5.HD��HC����+��v��4ᬳI	c�ƌL���Af9�2�̳��5�%()���'�;�QM���3LI�t�3)�Hh!�(N�=IS!֑��RD������Ha#D`AZ�/�УBR!PIV������X p4���H$�@��W-h� �qs�ǐ@2̡$�	pf�L��!(�ʲ"�(\L,ɰ&�R$L���(����3+>����4�7��6Q�����������I4�H�2�3)	�`��y%Οv�w7�o{޴h��oO���CMq���{Jx�Mu;\�^��tFՒ����8������ms5j�UV����J��α��l�C�dKyl���Ru-PR�A�[b��Ɇ���	�[�&z�h���#l����s.5Ͷ'h�'D����nS�ۨ9�36�]�#ָǶO�}l�t9jW��kf�լm��P6mS��,Q��nvi�b�)�ɕeZ�H��݄�,�F�p]�T�%lS`�Ӳ�E���l�gi��v�覰B�V^i�-+lsS�G�-Nܵt��+�ԹS���d�\Z��r�\���K2�ݫZ�@��k8��!�l��&R�]�;�m��h0ʚ��UJ�D��$��r�,+T�!��\�r�!xΘu��4�]� ���� ���H� -i�m	4�Q4�Jم�ݖ^1 �+h�r��NjN�ksh�-g�5\6C�MC�Q�Մ��n����CƻZ5�8��;qt��]3�h�9��iW6�еq�@:.Y��rU*pwm;ۙq��L8��N�kG�����n蕊^�j��{nɰ���mxӷGNր/����+UUr������@J�ʆ̡�������-�{=s�u�!�X�F�Vjt�@lm��4�8-W�5N29 Kb�����Wgg͌L9c��U���!���n��d�����3������ؗc�]m�v�Q>�~.���ݧ8�#R����t�\�9��V�b���&���m*�WV��#y�<�Ϩ��*�"�+	���Nd@��SM�J��-@g;�l�Z���U@N��nÍl�"�s+Ŗ�ں�����S�s��˷Z�U���Q��,�Ku�c��W�lD��%��Ҫ�Z�g)���6�l�'��0��a��8+�t��W@��0� �݌fZ�<����[J��8v:�C3�l�d�7i9i#GIt����-��p۞[v1����b�a9T[1�[ X�D�8�׬;�v�H,��4~>��w���6.�G�?( ��9fy���]h�(����ɫY������r��2�"ք-�����&�� �m\Sl����w*f�¡ѝ�´��sOc`�t�OY�G�ζ��''n�vm��v�Y�\魈U0�V�ȏm���m���Y	�[�<1�(��z�����>�/�Զ��۠%NQո�-H��s2�i{���r]#n7��۝Y�V9���w�/ww|��>��5�z\a��ZՅБ�6��Ӷ��u�t��k���7��w����;@e���淳�R�������JR����)C��{�"y)Jw�ÊR����Ϩ�yFj�l�k{��)J]��� �S%(}������)���p┥'����|�)K��/��[�V��5��|R�������JS�}�R����{�����{��JR��~��],�k7�V��������~��8�)I���%)K�������x>JR����]�a��kY�7�Z��qJR��}�x>JR�}�w�)J߻��|��;����(K�ݾ���ދ{̺B�H�=6��wL헮vp�aY"��n�D�	B�jF99���y��I�`����p˛�&K$$�I`���3�W�{�C^����Į�%��x�c.a�<������"�}UV%��f%v �/P�$���fh��u��(n)%X��y�����O4���5
PC�.B*������@7x�i��y{����%���n�ڥP��R}��s��@u�YJ`����휵1���v�j*&�*�� 7�<�O# �s{���`���cNܗw�73i��� X���w�5D�y*I���ے��~�� o�e�Y�}��}v$���O# �T8�,������.�t��`���sy��n���3kH�(U�R8��̘y,�ϛ���X��UN.nj�;l]���I�m���'j�[q�ƴU���M@#
j������(��r����0�ot��`����L�.�D*nJ�IV���p-�v������Ձ�1`V�"�)���-:�y����0�ot��*�T_t�(n; �wv�{v����{�<���)BO�0@�T.}��?��n��(���$���۫�����X�6�@螇N�n.ʘ3��0j(�@�v�����ݡP�f�[���g�B�1�qI��	ʒIV���h-:�y����0jUC���'��bg��޻!j��wx���������8��-QDP�H8�y����0�ot��`М�R�$�R��w|=�u`{��� ���`��� ���Qt�!SrSN9ww7�KN��m怚y���~o�[a�5]�u:���0R�;���1�]u�2Do٬���:F��qFa�]�n�wh�WL�ϛ�Wk��L�!G,�&Я�aҨtz��ϵC�.(����;�v��8�MɈe��*���Fo��y����i��u;z1��\�m��=�av�޸,���h�\v{r=)�'fA ���8ZvL`6n\�n�ݎ�m�`󝋯Sw����rJ��3������ ��^��]k��ն�ۡ)�r�;u΍�嬕n���M }�J�Z��ݙݮw{��3]*�ʋ�4�e�`���?S;3��SP�����h��a�L(�$�NԒ�f��X���F-�v����<�[�!&�`�#�U����:Np���4�0jUV�ТjF&�Npך��}��=�����]X�����jH�i�PF���Q�<�,H���9�n^^���˔��!������T�RN8�����	���w4�@N��z9�n'뙏Ly�.��U`j�M\�����	.���4��*�wvhx9�����$O����0����
Zu��{ͼ�N����)o� �5 ԓ��nk�y��i�`}A���#�Dâ��M%Cq�{�����V���p[��պcz�I*O���I�"�Y���`ld;C�˞.��[��u�}���Yj�t(�IJS�$����V������#�=��h�T�f���nʫ�����"" �� =��h��W��{qc���FԕQG'8g~�U��{�ym�?0�4"d����?�\�����]��&��z!���y��M }�J�Z���J�9ݙٚ��2�:<����Ly�.��U`&�F���X�6�@ղ���2�;m,N�����=Hq��civ&2ev+-9�^K�z0�1U�����X�6�@M<��b���P�8�jI��s]�{�怹����� �Dâ.~&�I���� =��h���;���:Zu������H4�I.�{v������yW�߻�W����b:��w�� f*���I6� 䒬{ۼ��M }�J�ĩ�wwwf|ĺ�<#G�+�u�ڌ��^r��h]9ۯi�;0�[Up�(�M�FБ7~�
�`���syw7�&f�E
�D�p��;�ݾ�ݺ�31+�2��vg�2�4��#�i���UX{���J��g����@��߯�mfh��pI5	$m�*���;���:Zu��o4��`B����69"jI��y��+��o�n%M@nbW`G=3�p4tpy��3�K�Yz��0��'=��ڭ�kui�lF��]N�21���#SHL����ݻny;_}�o����3��F-�W ]��'+մ0[�7Fm�@��C]�2�(�(<8�ƺW���ڼg�jTt4sa�Սٛ�;/!�,�(:�ô2�.��d�.<#�S[!ol\���Vӭ�
�k�ˍ��Fwg�#m�h�Fzc�gN�Vϼ@�l�����3v��`Ԁ�z�睫��oAk�ѷ9��O$\߮,�ҫeE�LDe6��~�/�g�n0��ƁΓ� �@���͕vT�M]�h��� s{�s�� <�v��U��4�m�IH)$�=��pt�����@\�F�J��PLm8D�Q����� �wv�nmՇ���y�3��Q*�BRSN+ ��X�U5��]��uE���������o�4�fm��-��L=u������\N� Y��%"�K��f�?�su���>�#�i��=UV���f%v����P{���6�4T]8�MBI�J��������YU� ���;8��怹����� !J�tXL&���s�{^j��wo�ꪪ�����������]�a�,2��$��g�@3|��q*j3��ٟ�k�V�``:�JRnԒ�g���wwf�Ī��:��>�%V���S)�!�p��-GMlۮzL�#]^�����X$�hf�?��w����B�:U���J�33��pk�V����*����gw�����H��蘟��M����9�y����0�ot����=���"|*�BRSN+ �wv�W���9h��!J$<E�
�N�lB���6�5am1���%p`CJs���[�r��Ō�_�̮�56f(�%-�)�!J	J-*�~����ؿ�c�$�����	Mt>UWB���6;T6 �R`*~ީ�t?�v��M���;�����]���_~>��D��IF�-;��Y�۫���8�� �wv��f���CP�J����;���>�t�����sy����hnP�D��8�!ȇ[N^gj���
	���KU�7�fyk��x��|�c�br	I/�{^j��wo�g�n�Q�[���v�R�t��x�h#�3>� ��y�.o# ���@�I�@rA(4:��rK��ݺ�=�n�����`��߯�{S��tۥ$E��`A���Γ� ��y�}��i��YN��9n(�� ���`�6�@\�F����Au�f�+�ճ*���[q�&Χ�[��]oJ$"mms�mҤ;���"|*�DnRn+ �Zy�.o# �s{�s�� ^���qQs17StN���h���;����5`��� ���Qt�HiE#RI*��s{�'I��4�@M<�aBT�dI���''8�o鿕�{߷�����;����!�d�UIUU� {�<�O# �s{�'I�?"&b��MP�X8k�w�����e6�ݦ�̀L�de�����5����Z���8;Vɸ&݀� <�%�1v���1��W�7U�v��ǟ��;��h�IV��(c\"��l��[lq�lXn]ю6�H۷����#�Հ@�YbrX ���vq�;;�2��vv�l�����lj��M�������ƺ@�����=��e�3Sc����7���hT۰c��=�.����z>��V���BOM3p\%��j�u�]�r��Ѹ��8�R96���Q��ڷ%��������s{�'I� {�<���wd�UEM5q3wq�w��ߠ�9�y��nmՁ�3o�Д���9�3i9�y��i�`�ot����E$H(�����;�;��u`{��� �y����f�%:�R�F�-�w�O# �s{�'I� {�<���_��(�z�i��
�דi���Wl��p�V��qN�Z�<V;\�K�못���'8�4�@\�F��̤k *n������ך���U^whx39uX���}�]�a�#)"�骒&���� ��y�.o# �s{�=�5X��YOhEF	�R]�����,�7��S`��h�c��t�r��U���w�5� �w6�nmՁ��6T�'��6�]Ra'�Wrcp�k�c���4��S�nqn����a���Д��I9�3^j��so@M<�������䉒��������y��i�`�ot�9�>�f�Ju��\��� �ͺ�=�J�w�fkq�:�1��t���.��Y�J��E5(���V���p�9�=�ƀ�y�GD\LUE]]T�]'8����O# ��w�}����q9)�l�(�#����Ŋ����u�SL��Q�@k�9h����E�IUDM�UW:����O# �s|�P�5Xp�YKhEF	��.����;����ȝ'8w'����eD6馓r�$����8k�V����O# �)��*&f�n������:Npy���&�F�菾�~��� �{Z8�)!�Q�(�+���4!4�0�ot�9�=�*�}H��vPۋGT<):0�A",s�ڵ�`�^t�\�6�gv���z�4�Ŋ��5j��31+�5N��{����k�o�Ԩ�q$SNRn7%X��y�3^9�y��i�`�	D���
���������� =��h	���ws{�3�詴?����_��� M<����:Np�S
%��]YUYWw��&�F��'8�w��`#�.�@>�5	.���>���k��F�[��r��]���������'�TÞ�u����$��Ndi��e<���ov��X���n�l)�B�yv�u��sl���[��a� v3�]
e�����q�q���-���KT���a�=Kl��_�������˭@:�kv[h��݋�'kiá�0�$��䑟Ul�p�Rv�BOnu�
1���c���	���mM�#=Κlɩ5Ig$��:�q�n���<�AلX�n���p��S�Z�Ӓ�t�mH&���߹�3^j��wo�f��X�ʳ~��br)=v������V���f%v�c�����Er�qX{���1���ws{�'I� ��.��d��IQ5U`j�M@fbW`j�QA���U%�~�����ߩQt��br�q�*����@N�� ��y�&�F��TP~�^]NҊ\ue��6�x�;uȱ�c\��cm��
C�Bc���?c|�]����	�s��o4�����A%��`P�����.y�g�@|���ݘ����RL�����y�����xk�V�1VR�J�ݹ%� M<����:Np�m�.�t�M�i��rU��{w�5� �w6��u`{LU����"�I.��:����]_ �u5�bW`������F:���搐��8���(WX�W�5�u>g�Gl�U,P��?u�w٨ �j�*�� =�h	���w����݁��oҝD��\��� �ͺ����X�4�@p���"�fF*r���V���p[���
?���(wgw�v����ʰ;�*j�[4�Hހi�Irs�V-�v�����۫wvw��������?�Ȓ<�3�y��i�`���
Zu����u]^�6i;�3ݝ�\���\�Khܼ�
C�^�4`O�}��m�;6毳@M<����KN��m�.�ײ�I1�� ے�{ۼ���5~�΀3;��Z��FCjrX"<��>������ =��i��i�`���ǵ��$�N�p��aUUA����U�����}�|�H��hD�E��Aԥ�'�{��5ʻ��ß�/�#��Qꪰ�M@��٘�hZu��O4p��\UE�w�Y��Rv�X�D����d��$h��;q���=m�Չ�1��8�Q)ĩ4�Q9$�`{��� �i� {ͼ��������=
:.$�rG$RNp[�������������w���)���� �&&�k�@|�U���jfgvv3�J�T��l6�&��������Ù�;�[P��vS�(����c����D�4���6����8��vU��~�<����9W˳�L�_f!�[
"�Y��jInm�v+	��E�:�����P8I%�w@�5�O߰�F�"&����O�� 9�ռ����������;x��Ԟ���ݸX춀����q۶�//n�ll9<���
��(+`��l��e#h�Z�T��c<$�6E�����aKe�^ ��4uR��=Ф�.|����ó�k�J��Ύ{M��'E+���e��;T��ѻnK� ��<d6���l��dQ 6$����Z���جz{a�Be�jYW����6��l��$�ݶ�p4Qu�	N�=�]N�kk]t�����q��͠-�����er���<�๗�8m�n�T;V�E��i/�H맛��uL(��9nm-.��U��z��vb�]�c˭OJ�*U�u�ۑV���pˬ�N����i���^��]%����V���M���R��Ă< =lhӞ�G�:����4��}�Vn�T�ؾ�H�	S�P5���k<��j�6f�ɭ�6k�BV�gf�ON�!�9=�Ҥ'^^��Ӂ���Շ��a�l�su�����v�Gq�s�-V�,��:u�l�m	 ����Mc������M9yְq�.�1��!y��k�::kkv6�k�nrL	.�J�UF@YX��NȨJF�ix��z��O=C��GcM�i��P e��;�[��٠*�Υ�-����lN�OVp[�ˢR��u�\���'`�'\N�[v�;��ٳ�[Hf,���p�%�r��`^:1���q�6����a�n�<��J�[$�;9fe���ګkE�ݎ8��P�%�dr�*8[c<�q�-��j�i�e{f�]b�=����n�	ހ4�&͒+��s�R����
�t�Kk���(J-bCaV�V^��\q�x��g���*��v�����j �+J�Ur��n\mL��:n�$��e�畻<��x��ҫS�����n�+E�T�s)l�m�]\J�p�v�j]��U<��7+=�a�X�r���aێ��j�&ݘ�4�����R�R�l[.n�[�f�Z��f��z���_�P6� ��^���D~Nx���޳el�v�p�8ϐ�m۱ٺ:M�6Ć���B^vg���'I�nv'��ϱp���-� �;�{k]��ՙ�p�9F��X�ց��ѲѻU�F�!1ǌ��g��ۉQ��uI�q&���kg]n;h�-�>qu9�+tk	���Iə�l#�8v ��ecn�Og��8��B�e�D���0�=��� v�c��`m���%�Pι��zW&�;[Q��qk ���mg��N:u&�2Vږ��={_�{��w�tu�1���E_~�ߩi� {�<�O#"#��;���	Vֵ$I$�A!Ɠ��;�;��u@gؕ�
��a���bK��3�LE�{�Vr�j>Į�P�M w��|+7iQl�M*jA�$�
��;���Zu��o4�����=
:�[H�rG$RNp[���������ws{��5�컠.����ș`��=3�}�u����L��v�>̦l�}_*���P��Jm8�������`���Zu�B�_K�똫�5�k{�9�]����_P8	, 	��ޝ�k��U݀�j� ��X�C�D�4�ڌM�V���p[��>�so�n��X�f��))Q!I���X�i��y{��f�Z�$�R���I�`��� ��������'X�*�M�s5uQEr[m��v#�����8�Vz�CP/�Û�X�$l�FM���.��v��ϱ+�n��v{f�39uX	w@U1S�'$RU���w��U_$~[���{߷������++�b�D�M7$�U��4�����+�""#�>������Vw7y�
��-�/�b�)4�y����0�ot�� <�0���1VTUe]�f���� ;�����`��� �f��)P���E�
W�c:����
�V�n�A<ٲQ$�A�]���i����j1'%p���� �N��m����0|H��2D���M��]��I� {ͼ�7��ws�s�U��������m$��(L�'%�fwuX���7w����P��*0�RmJk������Ձ�{w� ��w|�P�D���.�X 9R����|�����@+�
�qH�H�f%v �W��U`,J���m�w�o��x[��6�vgU�C]b�vv�:���Ô��mj`�x�c����WX���]�������^ {ͼ�7��ws{�
��-�/�bQNK �wv��謁��j-�7w����P�l6�&�.⢫*��4��`���I� w��| �-ke�F�cNJ�=�ot�� =��h���9�L�d$R�)�#���l��so�o�i����Y�2yh~�$y�L�'��v���P�]�[BR������d�.�m��ԩ�Hn���V���u��^�qf��Y���۔SsH\k`�l�Eݠ�m\P0l��77c�]+�nÓ���ʭO&� ;Y������\i��h�clBcl�6ܜ���uέ�X_it%��82[,��hcP�8e�ڃ���K�m�o;�*D�+��W%t��D5���"���F	6u/mu��.]�4l�dOJ N�k��~�������0�7��hI��B�7 7��������%M]nou�%ް�so���}�7~@+�
��ImO5���`uz�w�>Z�@,J����^2��SM��n�
����X7so@|�F���@#��qd�M7ASWx�4�@�>���y{�� i9`ow�(m��䊡Q�G$D�.΃P�X�A��t�8�ʌ�R��UD�\��>��t���U��*j>Į���3��;�@���| ��[?:%�&8Ɯ�`{�J�]��A{W���ML��{k�f��)���l����i�`�ot�n��ffn�j�n�j���=�h���w����w6X��)J*$� �-�����0��Ӽ ���@n�5.��6k���uv�"5���CM#��\�٠�]�a##�,�eЛb�K�B�����Ӽ ��y�F��yk+�b�D�MI$rI'8��,��U`%���ϱ+�fgwvf�Hd��z!�&"=!1>� fr��MG;K;<�=��s��n� �X�>��`ݿ{�VZ����B�4������l��F�ۍ�ܕ`{��� �Ӭ ��y�(by}	�]�U�)7lh�N]<q�pcnp�� <cf�\^����Ѻ
�T�$�s�j�׀�O4���;���	2�E�D�
H�RH������H��]X����V����)ED�$�w|��0�7���`�'�M�
�$�#)A�VFwۼ��5�������>&����ʿ�K��@�7$�s�j��`�{���7۷V���p��-����Ф��5�j��`���5���F�z)k�C2��y���?��$��Q�NK �w6��v���s{�@ �w��Jt\��5�wy���0�7� �w��O4�����tJ��m��NJ�=�n�'x�4�@|�F��qAvUM%�Uu{�}I� {�<�7���_WԳ���xo�~u��RG*)$�y�����0�7� �w�(��������	κ�J�4��mL�w�{7Y"G�W^�m�Z	tJN�8��i"���ٸ|��2=�W��Avzp��2��۞�pm��c<��+ؓ=f��O[��8�n��h#Gl�j����"9�U&=�i�V7g'k.�]#�G9��.3���{g���m�(쏗( ��q
B��SemR��÷<1N�x{q��ln�����f���{�i_���2�:)�^G�hp�wk��f�#��'$���Ҏڀ����[qv�V_���fx���;���I�DD {�<���uI����IV���s��;;D%ޠ�]Vĩ�݀������D�ӒI$�s����;�;�ݺ�=�n�uW��Kh�T�� i�@|��bT�f%v��uz�>B��>���*k&��4��`���s6X{���=^f=pjA��'&��aU$�rtN�F��ġ��pb�����j���Wm��ۍ���`{��� N��m�����%T�쪖$H9� 73e���_}T���׭��������8y7TL����]��]� {ͼ�7����w7� ��`gp3QJQQ$�|�.�o�n��J�n�Ps3�fwuX	w41L"#	��{ۼ��������ް��bT�;oji#�2���1Ҋ\u#:�l�kt=�g�]�uki3�Mĩ� Ɏ�~�S�E��D�ӒI#�_@?k�� ��y�>o# ���@��*�%��Sd@Ӓ�;�ݾ}�o�n�{ۼ��l����+X}H��9.��SP���������44��)�!���;�333,�b'�#)Їg"��!�U�jك�ш,�/0
�
�C�^�޷�u(ka�	����LR�4�$61DTS�%M%	T�f"d/��MB���#J�sE8� z~?�U���x�i|@�A�C� /�ȼ}�@o�]߻�W���o��ٮ�Q1���I�VUU���4������y4*�DcI)#���l�?�����{����?g��V���p�1mI�In:�2�� -�7#�2�mS1�%ڎgtp�Xh�s����*J9 �E$������T�f%n���`uz�ߴ�,4y����f�/@|�F���4��]��¾����3v�N�P������ i;�=>mހ>n�Fz�Ŵ������rNp����s6]_��{��U�{��*@Ax@��[��yW���	J�6D9,���@|��ot�� :S����6i=��9')��O\�'e-�p�%�A�kxlݙ�� ���[�Q��Z��Te����� ]��4���6���k�TLbC�'%X��y«��"�N�O�w�>o# �R�F�����pY������U�U@>o# ���@��8]Q36]Y7�ޚw����X���f%v�;��$�6X���E)ED�mN9w8ĩ�vf}����K�@}$�`c��������m�H�7p7E�+sfƦ�^['�#�۝�&He�+;:��W[�ET��F��мͳ���9�*m^$�s�I<Hu��һ\qw`�1��v �G�H�n�:�c�$�dܚfw=���+oW�l`�ۇ���
I�iOHul�E��o�v8��n������9i� =C������8��p%��=c^ݍ��"s�+T�۾����/�ogRv�Xu�gzSAюHљ랍�c��Y��0�Bٷ�����O��.�mN�}�]�-����%�vo�;�SP�(�_�TI2F��9���`uwwe���j3��wxfgh2)�#��2zb}�#;��Z������߷�����A"Jm��\�;��%����Į�����%� [�ֺ�#M%�7%X��y�>��չ��������u`w���d`F�m�\���jz ��r&�ٶ��I��r�!�!P �Hc��4�)�A��8��v��K�Z����w{��K���zD�)q�9#�:���������ԽU�Q}��"4z�# ~m�&��ГTR�TBjF��s�f��X��y�+��͖Wwvp��T[��J��
����� M;�=>mށ�ɧu`v��V-�Q$ƣ��$� 3se��͓���\����Į�3T������'+s"eI%"���>[��Y�H���]�3ݘس*l]���Z�m��6�@M<���؍ M;�!J
��cM\�� �ͺ�����8��,��������֒T��:�0�ot4��QEWM�w�&������lbRG9�>�����}�z�վE<f�w�]�=-�P�mʎI`uw7g �_o�� �g���nl�7�c��E8�J���q�a��u�rgHt�J���/+YqӺ��)��{�T�@)EJI�F����76�����i���n�	��2�䚛����0w7�}�|i��\��sn��W���+W�ULj9rNp�?��=+��"" O# �&�@��M��DIӐ�;����3sn��?}���~�8(�$�jU}�o��Xx�������J��5j��fw��*�Z�@}��`s���������:�cp7 MP��X���cŞ�=V�DtpvHW�<ņ���������g�o����˰Z�@}����33�t���`o�4�Dbm�)#��i���N����7ɽ�DD�}���6:hN�n��f���P�s9�f�=����T����9&e����5s{�Ӽ���J��mf�*-�Bj��%$����p�w�yW'Zi�`�}�x�,�����#�Մ#����U��]�z�V.�)��uY94�<�[ʲ*<��
s��q���գ��\:�|��3��.2�j&ݙ��3%�av�V�eݢ�v��nC�Q^BG7A��
܅���(�l͢��VGp�k�i�=��f�bۗjv���ȇ
�<
���b���Η�n��B�G*C�$�c`�����\���8�d�������C�kf�$b�٧N�:�u�<�+����¹����7h��p~n���������z�ߚ@M��<���4�0\���J�kX�I���;�ٯ�f��X\��i�DG�����A�,�����+ީ�5j��/q+����˽@f��π[��i!l�R��?}UN㳳3�|���yw��sT��SP�`��I��R�9�nl�;+��4�0\��	�.������E�.���#[b]�K��]c���q����Ҟڞ���{���r�w�=�tl�X�rw�.o# ���sN��7��TBj(��˹�3۷W߫��z��">���9k��4� ��N�	����Bj�%,g�y�nl�8�ٳ�g�i`v��+�I��"�?]�3;�3333F��PGow���Pb=��p��:U�蔁J� NK�b^�9ٙ��ffv[�� �W]�b�,�b�F�9#��RD�0�r��Ƹ,h�dBٚۮ���mɬ�NtX����w�NI��*J2����ـ.��@9�x�vp+qеQSdR�ۅ����O���N���ހ��`	�YQ��rNp76X[�����kG��*/ �����������kZ��(R��I`l�n�ճ ]��&���72
QD�Ґs��� �ɥ�����U��3-����ޠ.%�T�%x�D��.�S��"Ɯ,�rt������5�m�7l㔎���ʉ�*0�M(�	����{�	�x���ﾈ�@M[0Gt�ߢ�rEs� �͖�vp[�P����JZ�X�@L��HD������V����nbW`���3َ������r\��;r�����ʯ��w��P>P@׫n�p+qеQ1��n{��@RӬ����V��BwaMk�M#��Ya��;�q�ۄ�V��nYj���X:�N�獷g;Z�^�a������X��w�&���D}D ���1�-QTE
T@��I,�����/q@nbW`�z������:�]� �Jm)JNܗ:����3��� 3se�վݜk7Ul"4���P~3�����.��,K��3��6�M,׼�ߥ*i7#Q�9���@|��V��%v���A݆rJX����L�}�/)"J"�����	dځ5����'A��hJ�G���EU%�%�#��*
!�p�#��gY�	0g��-)��`P��x�9�	�0CZCT �uG�q(!P��Wb�� �@� ������{����h 1S5�^W��vC�!.i"͒���m6�Z�$ut��N�m�ȫN���rE
���zfK�Ȩn���R��qc\��u5UeH����8:)y1 TKC��4+*�ݰm*`��'T��Gi�i'I2$m��)�BO1�pضb��F�W�5H;���z�R��'q�[E�M��y�8�Z�unq�X=w'E�P ��UU��[��m�j��*d�� ڜ�Ml�tk�^$H�IBi�N�k���vv���̩�x+��<�v�C�rl�j���N�����^�;3�v.-�Ñ�
��[�:[�CIK�[;u�=��g�L3�ڌ���Y۬6�-t��cl�'h;\���
캮A���\�k*B��[UU��N���^v@oe���3�W�,��yul$D��E� �\C;.!݅��!�&��;6�vlh�v7Yr�fb�V�G��	6p�\m��ۺ�����v�X+s��bO����k��R*�9�ۤ�6���+n�%�[�����1��Yť�I���#DK�I�U٥gg[J�q�7��]�e��ͺkn����ssd�X��2��@�`aBh�/ �]���)'l�me����n�I6�<�M��H[m���vYlR�8��ɺ�q�Mv�p.�۞���ED���1��#
�-��P3��^��-^�\Π[k.�m��qqٷ="���Í0p۳���0Zj�^wV�I�8d�G.:I�v�"/9گn�i����mSʫ@/cqMf׈2���t(��5J�+YN`-��d\�u�uж����^�Wj4�����V���kRR�̫�me�\�U)u���V��D뢶畑�-L`;n��0mԵJ�:J�:�q�,���+,�\����9��V�ĤPn���
�)6�l��PI�Wj�j�=@��e��):l�K�^MȆ�2��c��\��^���=��� 4��y���
0���m��i�JV�/׮�_��a�� ��D�ES����9�l�k[7���F۴�w �7
���Hmom{tk��cq�Кd�8N5I���$'a��ێ�����vI��9�n��i�%��,k�%9��g��e�	��\bC��n�ܑ"�%@�`KWmmB uٲf�+3`�ѻh�S���m���M���ċl9s�&��݆�e�3S`�]�]�r�p,m�9N H.���{ӽ�w��,��ƝW���ː��7[m�!-�qge�����a1�UJQҩN�H�F	ɠw�����ob>���� M;��T�"ɒ�*�'.�ճ ]��&�������������t-BLnDڪ�0���i��\�h	�f��Y�tIq�p?}�%����t�t�	o�@�����%v즅��(R��$���n���K=��p76X��ڑ��q���Q�Sl:6�ȅs��Z�����.�ڐ �ٷnڿ�z�:���J*!��)%�o�f����Į�5j�33�3�t�t���a�B!SN!9�����9��H7����<���ܚ_�����T-�R���j;�� M;�<듭s�`���<���VӢR��rX����3��j��@���w���!�E�%�UN^eh�� ���sN�*���?W��!��pjF�
��M��vru�I�.ݪ���Ziq���t��j���{�>��|�1�j�p�;���8�͖q�u������?��F�ThmФ�{�)M��\�hݳ ���@��j��"�*(��)��~�|۳n_�r��� ��d ���������`op�h������M�<j��ū���Ԧ����ݣ������tU��TӔ��8X�c��7X���@��|��wOU�(S��Q�8���8���6��`����N�Z�pX�^��PS~?oț�esw�rv�˛��	TL8tJ@��R;�=�8�f�sۼ�Y��}��aPU�����3W�@}������h��ް�t��#M�$mSnsۼ�Y���q/Xk6;�3�Nʪ(M�	�D46�)���Y������͚X�n��kj9J��m�RGr��1i�ev�Y�cZ�KṠOlE<�;ڑg3�SE
T�5R;�}�8�f�{ۼ�Y�����J(�⍹9rW���P�����BĽ|��ԑ�o�E[�M9I�ۅ���߹�25)��ݙ�2�z���q@cc�1P5#JI9�1f�:�۳�{6i`w=���Y��m:% n�Gq�F�^�9�ٛW-�#uM{�ߟ������/\�G@<F�vs�d�]n�z�eE�ܫm��:�ؙd���ȸa�/;>)6��1��p��3l�n�/(��v;W2Ul�#h+5��x���N�9˱ٞ�l	�l)�܏j�203kӰ
�*�v�.���u����h�w�gF�Ά��l�Cn������R����[X�'9)���4�Oav�c(ù.3���`;a�ƆB5�Eu��X'�k��e���Ē`E�������Z6 �v��]nF�ѣ�{w��c�C�������� ���@�I��\�hs]%���i�tۅ����8�'X�su�y;f �q*�L��U7d���ғ�ʹ��<���<�w�3tV�����Q8���k�<������:Ru�/!�������������<������:Ru�w_�_ �W�U|�񿤨�Dq*�*�H��,�k��q���8�箻v��T���ZҶ,�]�D
���RW �g���Y����k��۫���Tm2R��r5'�����3�;�4A��6jT�wۼ�U��V�	@&J�%#�;��ցɼ�{���7X �*�Y1utLQYy��ro# ^��@�mՁ�~�| ��Ih"4�nH�7%X���-��<듭&�0�'5n����vV	�ũ�^-Ӝ"]˛k2vu��CU�2�����LV���-��<듭&�0�ot��Ԕ�B���G��~�|3v� ]���۬y��\U��U���T��SP�����wwf�wj���5����i��I222F��w7�Kn�:��@I�0Gv
��)TM�"�I�囮��n���0����;������J.r�&���GSz睘��S�t��CA.�1��ŘT�Ja(�QĤvu�u�f�`���:Su���!�E�wS1Ee�V���3`��\�`)��<��_꯫�� �k��M�$J�p�7;�����)Ħ��^E���{I$�j@M�p
���w]��~�~U���nW�"!U $aMw��y�34�dt�B���G��~�|'l�s{�t�� ^b��\��=t��!n�lu�S��e:x�s�\^��kpI3]7����G�ti9fV�|}Znـ.��@R۬ι:�;��J�����,�y�1n�<듭7lȈ� ��L(����������Kn�:��@���=� �X*�a(BnSq)��~�|uy��]����	)���a��Y1wu3V^eh	;f �����vu�5����J��HېT�c^BS�rpv���mr�ہ@V��9	xLIP.ɠ��������F�����ύ`��5����g:�r���/i��t���V��4J��.S�[��0{+���P$7j�Z#n;d�2Ƽ��1b��1���7.���D�Cr��uxW;hx���4@*˷k)D��ln��6�l���c��܀��p���z5����w���n��pWo73�#��3�i�<Yў���O��mѻPZW���O���x;�Di	ԍ&9+�~��9�<�u����_U}�=��Vm`��$�m���	���۬ι:�9���/s{�r�U��*dbQE#�;�ٯ�{wm���ٝ�f�]��wM�i��=!����������9���/s{�)M��~�|<Z
�NS���;���gfgq�Ԯ�3�WM��*j;Zk{RD9(�F(&����#U0�lNL;=�e���+�Ln�aG�[Uz������Ww7Ww���`u�ցͼ�{��uW�
��J��JG`w_�_=G�X>2���|����ʳq+�65)�fvv��K�/� ����k�S`oOtP�%vs�B��4t��| �k��i
*I�M*I�a���o����h�橰1JQ@$i)�$�t�9����u�����=�uX�n�{r����'R� 1�u-Xu�Y1'ZA�p�Y�e�6캘�Bg_*EW�)Q�E���?f��{� ��7X���n�,�.�oo2�t������� �N��3�������8	�`s=�����\����O�= �d!�Y�H!�'����tHҚ��-4SFA:P�Z5�Lt�$Į���u��D��ȍ�����X�8�8�84��	��dy�X�X#3�L��NPF!J����UKAD@8�"J�X�� J$�&��ܦ	��kY��beQ�XeUN$��!�b3�;"@��I�l�y�h'���Y�60TLH̠���IAI$FM`�ؔ�d D���E��A�(L��H��mH`�����m��ă2���qD|�_���`��
		0Պ�h ^A��(L>@x��8Ǌ>�8���"z�G���»O� }�������uX�z�Ŵ�J�q�$��7X�ru�s��\��U傭�ڔ�JG`w�_ 򔢀�Į��Ԧ���%�1�F:u��
n�g�tp��',׮�7��۫qq"�7�wt��%	N��]�����ʀ߱+�65)�fh���`2��B���)�I8��y�1n�;�ٯ�f��`n�,f�Ht��	�� ��X�ru��nـ/s{�rcVD�*�J9v��^�3>��~����П�>�m��7�Oꉸ"��z}�UM��*j��ou|������c1=���')��&�	M��wF\Ό���A���v�g�x�9{vl�Ȃ�rprU����8-�vu�5��۫��QX��4�rD���	)�a�3�WM�����߱+�j�H�Z*�N�HN"S�8�~y�� M��{��Kn�rU8��ffˊ�+/2�M��{��Kn���k��F��JiRrU���W`s�3)��3�WM��*j���Q_ʂ�& 8�e�Xg��[�2&��:|'%��i�i:��N��0��"8P�p�$L�VQ\z8��h���X2��'��p����PWG��ݞ�X�؛ݩvWg6[���p��esҽp��Oq�u*��d���t�H;YؤҐ�s&۷�]�!�fhޫ����������[�&[����u9�"�B���q�l����ps�v�����wvq�ul���`�2�H���>�m��M�g��ܰ���C=�=�Ґ1�d�$�C��I�ށ�w�:��@�o#">{���d�(_%*4�q8���k�ݚX�n�b�k�3�n��J*"�9.� �V�{��" �u�y�'Z�hih*!' 7�`g}���ۮ��f��ɥ�����[H�q�$���� ���y:�9�f ���o�!l�16����pc�:U�F����b���6v����[)�@vi.�`䔌��r;�����&�wۼ����=�譧�IG�˷�=��T;���c�3Hnj��61)�>S�M�x��4�'RSJ�p�3��� �Ħ��vgfh����7���5>F�&�huI79�*����`w_�_ �����{w�ٺ+C��JTbMG#�<뛭��`����u�{�T���Fn@{kN��v[bS��B��u�a'g%H�A2MK�N�~=��}��Ӗ"��=^�M��|�s�c�vg{�Ν�s���KL���@nbW|������#���-�)���*Ŵ��mI��9�1{u�[��e�36������z�n� l��hT�T�rF�NGa��^�3���3����]��� \�A*"买����+@�I� B�o4<�`u�ց������?o�P]��ũ���r{S�j����RG�g�R��h�8ŭ��[������u���)Ħ��;���<,��	$�J(�ns�b��ι��9�s�.��@�l���'�R�j9��~�|��U����8,�vwߝ)EDT�S�[�~�Y��n�]���M�����vox��q��U�P=N}�w��yW����\-�IJPj
E`g����7]��~�|��U���l�۩%)RD4�������y��\E�S���u�.R��93g���H��ԑ���n�������=��p���Kiĩ$�8�� �n�t������u��tV��%I(t�r[�ך��y��B���t���"[�j�����<����u�yW7Z:Nlҽ�[@�m��(M�p^�v�8���TPn%v�k���^#���dc�+ڲ��m[0�6���,����]�+\A���F�vH���=A��q<l�vJm;=(���(��&�P���k��$��Ylө�E��S�;����g��N0*9�U�j��Ϊ�{�89�b���9�F��A�l���n��n�ӌ*�9����A:�m��B�p��p溓6�7m��<�ݜ�Jݦ��Х�q�G12��+`Ƨ[;s/M�GBH۩�}\jN!(=ef�f�v*$"i�����Z:Np.ot<�`�D≸"䊰������9�s�ys{�)����?n��5��RR�qX\��
y��<����'8��Kim��RI��ۮ��?n��y���{w� �z�R�q*T��I#��*��@�I�����������\�^x��>�$ \;:���1C�8%ǭ��,]qo���s���r�+@�I�����ʹ������6IM*M���{w���J��.y��9�N�jـ6G*%�$�m��s��]��~�|ۓK���pf�`�*J8�J(�vUsu�s�� ]����H�P�Rq>Io�{ri`g����ۮ��n� wL�B:���(;p��<�$8�����pxz;s�\��q��t��0��U(�!JpI�`g����ۮ��n���Ś�����Sn4ܫ�� �U`j�%Z:Npܞ�{�Q��*T�q�������=�79 ��$�
hT7�������7]�gs��	"��1ܖ�)��j�c��f����6�~�¤�6�M*I�`g����ۮ��n�����jq��Q�J(.ai1j`	o^�B�����L�F"��N�B�9��m�P$�4�%$� ���`s_7Z5l�s{�rV≫	����������<뛭5l�s{�)i���|������(���������`����� �n�p�PNAB��2���{w������9�ټ�N����(�6�1�&b}麺����� �n�ճ ]�� Ņo�e4�G%	�9M�IPݜp�i&Ⱥ���*�T%iTqڍ�6����Gnn7$Q��]�v��=��p[��=�譧�I����� �ɥ����O7X�7X�)�d��q��7=��p^�v���酁��cKhM��r��s�b����u�yu� ]���[�&�&%9R6��G`j��;��X�f�}����X���R$Ɉ	�l �]J�t�m$��Ɖ2J&��Մ�R&C����o{F��6��8E�����2 �2���A��B@��`B̲0	+0$0����0C����
2
@��1	 @J�1i]/��9���%	�o�O����Q)S��vn��ª�����*I)��6ؙ"fL�k��v��e�Vs�g�kkH춸$����b&�6��h��v��(Z�����vxp�L�����S`�F�e��ﯟ�5U*�^��3\M�&���ˆP�r�P�u���76SB��V(x	W�ηF��4�ڕ@RN��M��s�k�������m��+l�Lm��p��X��Ձ�� 6���!��R\���:��UUꪪɜ턳��qm��V$�:����r�d�i��k��[D��<d �V�S5j��Uv���"�d��J:���۵�Q�TeywDp:
����@�j�jv�g��Z�rsۊ�W9�핗˗f�g�d��u��f��p@���n�F�
G/*���l�UUg;�a�� �ѬM���Sv��-���j%���P�/!��ko 2�d�5�L�*�ܹq��p�3ī�T�s�ؐ'��GL�a�f�c��s�Vx��cF�k�|�e���Xۋ4u�PmΚ�m��K�'D�6t�Yx�5Iq�`�'F۴��ӗ1at�!#)R�u.�=��k�+��5�ӸXܼ⚕Ӳ�ڨ
�m�ZH�P
�lu����v�]TE�����Jf��]�V��&����(c<v\�ql��7CAT1��ɔ1p�8�
�*}f8�7�ۆ!ܞ�l��v���s�^F
ot��|%Fx:]=�i�LS�+�#n�%�q��d�d�K3��nͶΫtj�rT�Hh���9��g��[���ì)�9-�RY3P��F����˞��li�՞E��a���%���t�C,3Z��&m�N�ԧK�2ɹw"CT��Gl�F�������yY^MLW]���� ,�ݴ�#v!�V\b<hy��6N���*��U{<����V��A��Nʲ��&�A���n0��ϲ����yb���R@��&�[�9�"��ˡ_\��[mf�l�����`g$Gn�f��������h;�k��f��_���qE�"�U��GI��W��W�b�D-���湙�l�Z�����k�����u�g�OVc���:39�����*��hXjP�b�n�����"Zn���r�p���Ŭk`�9t�vv�v��ҋ�<t�\���M�Ŭ*�]��h�b���7�X��̭ɺɰ�<Q�k�-�i��7��9z'�D��B�/. �x��g�������6�V8NT(��[z��Լe㟜P$#��u�U_V}K�-�$�B�V�c)��uۧ�����.�(^s�Z쨶ܼ&�CDS�(���)H����7�M0ܞ�
y���u�o�	�.f&n&.�*��r{�)�� s�������,H�Q(��cq�9�1{T�
1)��gg�žE �{��1�#i�QN(�	$v���酁��o8/n� ��:+i�H�T��o�b�"��wvw[����4�Jh����~�7v�s<@¹j�\���	�W����g@ZUã����~ܿ`�'*US15Vh'���n�<�`]h�3~�imI��nP������{�f}�w�O�h�=�����ݢS߆9(U�F�Q���?~vs�w/���u�rR'D]�w[u��sV�w'��n�<�`�c@��RDA�`g����ۮ����`w=�V{�ֶ�%9(���=F�Ru��69{=�\�q۴�E�6�#��{R i��R��cq�9�1{u����<�d`�=�:%⋘"�nOx���bS\����b�M@-��1{u�{1�[O�%$�&�|��xr��������,�����.���u�h�Κ �o�b ��L�\ԑ5V`����ϛ�˭oٍ-�I��7 (�8/n����;��žE�����A�����560�m�q����`�Ō�i4��<X�HN���2n���@P�(�H�~�g�� ��F ���O7X��.��R�J9�n� ����UUU}T����s�j�ߝ�owe���b@���(�%U�U��ot<�`�w��O�b0a�Z�����q�p?W�|���΀;{�@}��(!ݙӰ��Ϭ�䗻8��h�S�R���; �n�ʹN ���O7X䉗tU]E]�=�:�^�2R�t�%��2��,ۮ�y��v�tkr�����E]?�������pk�V�Ot<�`�� <G�$�.�*f=DO����W|��� ���kB<߱X��Ƶ��m6999�1y)��z�vvgg�žE �W]�����JJ��$R2)�o�e�����]���r�.+�����/r�/@歘�ot<�`�w�{�}���߮?at�[J���Gm����t��:�e��������� lN���AGM�n]�&��dl������`͂�,ͬ<�fvmշmV��lݼ�=Ҷ�[�,��]#<���\-mu6�FM�5�5ճOX8�d�������-Z�=��dF����U������9H��;U\�7Um�a�p�oHY�g���pw97;$F�uߎ��g|/�p��=1���Ӊ�N��|���a�����s�l;���F	�p������]�owb��w=0�9^񂥿�nJm�$� ���`���֌w7�� ���������'#����X�L,��o8-�v�̧F���77q��7&��ot-:��� 8�$I3sDT���D�Y�.��@RӬ ~n��L,��3e8E"�*(%*!D)�n��m�{/�m]���c4��g�6ݝ�P��I�������5��vX�L,��y�=�522"�jGDn; ~n�.=}���^���X���O�T�%�n� �ɥ����8-�v�ݖ+���*!%	I�]Y�.��@RӬ ~n�]h�;^񂥿�nJm�$� Ź��7����za`g�����%�4��>�Qg��mfB+;m��ͬT3��v���Wkt'h̃��AJtDP�Dq9�owe���Ҁ�Į��Z�� ���4�x��Lצk���(�J���h}�,�L�i(�M4�
M���{w�aj�����w��{����Vy�f&� �m6')&�8-�v�ݘ.�`���9;sE��rU�U��U� ?7x.�`����u�w�c{RD�N��A��$s�㴻.k�iғvz��&�m6m����S�o\{\�������`����u�����bAl*!D�M�,��y�1y���� ��F���q5Swuww{�)�� ��˭�otǫ-�DE	ģ���?�UT��~����r�5;;��0��P� D̐1�Q�i*YB$T!	P�!&D�� �$����Id��H��b�PRČ/��翿���s߰t~�A�Hn�w8��~Į��Ħ�ڽ@s3�;��ކ���f���VBya�Km��q.B)@ϓ��9G�k��IN+���u'��	ہ��~~n���� ^n�*�8q�^ȁ&�lNRM�p^�v�͖s�;��pf�L�%Q	�BwX ���]h�s{�)�� ^�	�q?dM���V^��[0ܞ����}�,W���WED"5)�� ]��� |��]h�t#�({���t�lݽ�zֱ�6n���W�ba�4m�M�X(�T�Q��� ��*��q�5���f��L`�+�a�pjRm�f��e��<��SE���ɺ8�� $��۔ۣn`��v�%�M*��l�w9X�f�eŝ��$�H���6��gm����}�ݻ�n�iu\h�v�����۬��i�;v&�r<e��;b\6�����{ߗ{��s�{������*�]��n���]��wg�"����5�\eK 0H��������q��`��]�>n�.�`�=�:D��.H*������ |��]h�r{�~�γ����h����6�Cw��=�4�s{�)�� �� ����f�b�b= �3������{���z����/Ki�~�J1�9I79�1bS@~<vwz�žE�������fM����jtVѺ�����]S7M�uK] ��v��Ry�:�v����րy��7�|`�Y�t�*��B�f���Z�y�o^U�~�nqD蠳;�;�z��ơ{~W`(IM �䦀����
�R�Ԧ�wۼ����]�vs�u`v�������;�����u�9�u�yr��s{�=X�k"�ࣉ��{�,�F ���O7X �8����.⠝ۊ���l�����f�����hۃ��cn�(�a�P�R���I7��N�ɥ����O7X ����
T����MM�IUf ���� ~N�.�,�1��JSN���s��]�w���/�;H1:v	�0��e� �3)��&h��	54@E�@03%��@xu����J~JBr �C�M	��PRSLB4 �4P��@J��������y$KJ9TP� tH-
�R��-@���p$�)T��=�A5��"���L�T�4ґ%%H���
�%��I+����4�����"�>)>zN>����� �j(Yi�%\�H���"C%BR�LQDT�,r���,��P�J�e��J�#F��,{�XՐi		��I��΀n�}()�����
�dW�-��b����p�:�P�P�B�Ç�;N���_x�� k8 ��l����,�Q@oڕ��bD�R���N	'����{KۓK;����ۮ��k+7�K�S���ܜ��`���
y���� 5��;f��nؘ۳��kl���73��K7Uًۧ����l\�n�J<����ޛ�f�{��O7X ���l�5l�=M
_��N88�rNp^�v�ݖ۞Ҁ�q+�wx��YKGHh"'�7W5wX ��^�֌W~=��� =�h��D�q�������V;�{�}����I�G��Hb)�?}��UQ�rX5@�t�Q4RrF�_�t-:��w�r呀{ܘ�.�i�]���Rb��O^����.]����m�:�/1�ި�9����L����h>��76�����]��7����:�n1�Bn; �we��ͦ�/�J���k�� �ne��<�]�U{Uwz���7���`{6X��)P�� *9IG$����p-:��w�r呀lt!}.�iB8��Np[���͖��u`s�w�yW���Ο�s��oz�f�Cs��X�N3ɱ���[��vL���q�C���it�[.�Y���G_�_o��E&��t����5�/<�2�t��6D�,��x$A7<p���ö]Bn{��iR��*����۱oc:��-�Ɏ�[v�u���1�c���n^]����Et�R��K�(��dU��n���u4�K�'�m��v�o;x�H\�W��{������ۿ?�sWa.G����y�����6l��o]�����ι�d��xqs��j�S��o�[�76�����]���M ,�K	��$�hn�8nmՁ���8-�v��� ��̠Q�m��)9*��{�)i� w���,�4"�]�I4�ۜ��5���,g����sw�5�f��TM���8�����d`�ot-:���)���.٬e1�V去t�4���srb��qF�J5���&2<�z㶹��
נ&�F�&�@RӬ �7xǹR�]A9MG$����s����EoԀ�: �m:������\���o�~�߮�׫�~�!5�I9�1{u�y��<�d`���
�]r�Iv\��`y;�<�d`�����{�:6��$��۹�=��V�ot<�`�w�~G�}��l�eٸ+v�͝ҹ����:5l�kՍg�ٴ��������q)�Dn�������c� ߵz��si�Zl�oz�J$�����ۮ�7����{.���yΤf���:�n!9JG�w�{�U���×�A�P\"�fs{��w]���Vo� J�&78���	�f ���KN����6=�@+������q���{w�� ����酁��u��	NB(�RvӘ4�q��'a��Gom=9�Ƚ������ڥG��J"P��rNp^�v�ݖs�=��pǫ-eJT�jH�n����<�р.��@S�� {ެt���$�Q5qܜۓK=��p^�v�ݖӡ��i�����@nbW`lbS@�A�N��� lU |*�����W����7�� ۜ����{�,�{ۼ�~H��l��R:#I��b�t�A���kPstp�e���&�m���jv���$�J�4�I�QH�{�,�wۼ����v��J%*D���r^��<�w7��n����6;�]
�H5����y�1{u��vX�eՁ��ٟj�ԊG�n���� ~n�.Y�ot��t��&������7����za`nbW`lbS@w͍�C�L)������m����R�l\�7,�5�-�9V ��/w���ʑ��� tt�6��h���N�ݢ��;�`��5�0sr��@s�V��Jʚ���ڰ��lQ��S����hN:tD�J�V�Li�Ѭ8�� �':��͉��ݛ��}����$���vك]p9��'rr�&M��]<1�!�5d��5;$���d9�.���nz��:�Z���j�߀OP~ؠ�_��l�6'v���� &&�r&ۮ��P�ӓL�xl�m��۵��������@��M\w' ��O�`g����ۮ�7���:t3�m69"U���{w��ٮ�7����_�X�X��P�`�n
���=<�`�w�o��������Sߤ��n�Q8�{�,�r�{�����ޅ�\qw3EU�U]��Np�otO'X ��,u�m�JQ��䡀�&�*�Ӗ�I����5��B��%�n�'g��wC�b��*�"E"�3��� ��k��l�}�U}���V�>����ԑ�#�sʿg�w\�U@���re�����ds�� �u� ^��@�TL��A����v��������w��ٮ�=�`��D�aN۷�;�����=<�`|�`��"n�m�"Tㅁ���8W�]������}0�7+�͔��S�H�	4�=��vݭ��7:v��t����{Oni$�4�݈�6�m'(m�p�f�Ws]���a`g}��ոSߤ��n8�R;ϓ�ޮS�/s{�zy��;С�	DIH�����=皬�y�����(:A肠m�޻���W�~���*�{�J�tD*!�#�X�~�p�n�Ww]�޿b�9^��V��M9�uw{�zy:����7��p���o�������Q��v����)�����:kg����P5�ɴ&"j -�=�ѳm�#�����ߝ�οb�3����^�v�z�i�m�M;w �j�s{�zy:��:�<)RE�U6ԑ*jE`g}�����`j�k�9��V�c���6ؚm�#s��U}�d��:1t����'�Y��[��)}5�����S�ȓi��r;ϓ�ޮS�/s{�zy��=�S��]p*h!�WM��.h��ғl����h��0	C�l��^��Ѩ$g�2uE�bW`}��;\F.�����WD�M�7"�3����^�v���~�`v����A�nI������ s�� ���������o�m��8�]�v:�����w��ٮ�=�,H�J�h��MM��N��+��f�f��<���U�w�s0?�QU��������?���E��y�sq�QTJ k�F"�&����5���� EEV���?�����������gߟ�������������߯�?���4?��[�ٝ�ݝ�������o�����O�@����/���(��B ����a��������3���**���������������m?������/��3m�ѿ����ޖggxgD�QU���Q&b"d�I�� Rb`�dReH��Dd�%�d�P�iP`��F�D��A�U�QhQ�QU"TH�BDHd�TIQ 	Q$Q Q$Q BTIQ�RVHQ$�!Q( ���B� FBU��BA	 	$"B����BF �	 d%P$!PBBV �$ $&@�Id
��
B%!
�P�BU�!�$@`$A Q!	UA�%	QTHBU���$e	% �B%�"@		���$XBIB@� d	af ���@���%aIP�@��!�!�%�!e � A� Qd	R@�F�%BP �XBDdP�%Y�e�!da� �!�aaF�a� �%�eE�!QaPRP�dE� UV��aP� �aP�!A�aQ!	A�	aAP!@� EXF  �BQ�$e	%I@�eQ�A�X@d�aaYFI�b�eda�h@��e�``X$IIF	@�F��R	Q&TH�S?�6������EEV>����3�w������袢��_�����5�?���s�w���~�������\��>������MQ���TU�QU�S��s��EEW���\��<ڢ�����G?��Fh�������������_�=�~DTUf���o�����EEW��?�C?��i�����DTU���EGww�����5����~�c�>o���DW��O����j��j���������kb?��Դ���n����w��_�?���5��TUr�_����hd���1AY&SY��a��ـpP��3'� ah��@ �  }     �m�    �   ���    �R�J�))RJ� $�B"���EJ(
QJ
��P    �  (�  J (  � ��9����һ���^O���|Χ�>t��I}�}��������^  D��02L@  �=w�u*�jX tnR�n�}�y:�qgW��j�  �� P ��T��#�R��� � �   �  ��` -� 4  	��� @� � �  b '� b����8  @ D @ {  �$ 
   B�  @̺vk��޷�}ެ��� }���ԫ�R�L�˓���Ku)��y�y��{�_>�_o����.>��U�wתyol������j^� �*�t��n���ť;�Ԯ�}�H   � 1 4^��e㻵m�5�����s��[}��}�U�}�9��w�s��]�>�}�g=�{���k�  ^����e^��ү��{�O-��O-J�����{��� �s�۽�Jnξ�v���n=�灠x>  �  HL� z��;u�޷_|sɥ{�:ˀ�==9:�s���׋.���m����y|n�:��Y�  6��>����_{� sҙn�:��z�͔�ri^�G���m\�垞Mzӓ�fw۽�� ��*{iJ�4  )�����J�  �=U*��L��"{J�i5Tz�&@ ��#%)P  �R�(�C�6&�����ҿ��?i`�*j;n��P�"+л��*��ES��E_��E_�U`*(*���<������l�V*R�����iv��Ǆ$.��3� @㷆3�Y�l��B%k�����H��M�*T�_��'�k����~X%2����|�Y��a�54�/!�렃&;� ����X��@��@#���2:Ѻ��j�`@�x~����s��p�6����K�qH�Ą���5��%P ����Z�!R[�������j�(p¤��0�j�y���A�kIr誻PJ����������*�"݄)��9��sZ�8h�%����Ň	�^2�e2NMe�#	0�&P�JKp��!L��,�5�5h��]S���Krk[�B\µ���D	�f����X?,��13Pvq�i��@`D�B�u�}��#	��0S䬳1���p���� C S�-0X�H����,p�p!LHič4�f�L��+�5*F�!S�����R��sC
Ƅ�5!,0e�b����j�X�mh��8�1#C S`� B�3 \ɚ��m�4�;�m����=��݌�������#S#�l.�\э!�,�0�cp���"a�D.RSY�l!pvl�Sܙ�l%04#��i��7L��m��FG
`�d�k5����´�"n�]na�p��2�5���!�,�5�4h��o\��~H,~� 5aYC �$�@�X5 �1 XB`��<�\RHRD#�"R9l�� a$J���Y B!F& I5$�kc
��A 22�A.��R�"HKi��U�&���b���?2��E��у����#,J�|��{0�$%0� �\�0�p�����c��B������%1+�Y�~!��?S�"F�-�MO��j�f��]!%�HRa@2�t�m�rvQ��:���AP���]��?I
�5�s�@���rCHm��uf�RM�!qb@�4n�tf�~���?~8��&�Y#`BSL
�a�b�d*B�b1���s_��>�����o�&�߉M��F�M�h�pJ�"E
�Z~~�0#4�$�[����75��럂D��l

l�",H$ #L!\I6�|���dn����f���a�Q�O��Ѐ ��Ј1"#!b�~`ARHB
"�D1�`$ 1H�K��T ЀUҲ����aK*,
��$M�%����!��H�bY�i��q�a��PM�t��K%����`@ ���!RVF!AebL$�YVÈ@*B$jca$���V*D�D�EP�Z0
�H��k������.h�h�i�t#&A)P ��`#S�,U��B�X��$hALX���V!!����d!LI��SX��	��}�����\�l3d�� � h����\�6B�˭CoӢ��r�P)�)`����
`K�4B��E2�qц���Le���&��?O���2�Z9���ԅ�E�p/w��:c
bJkz���\� ɖQ�!	3eѶoC��ZMᄬ)0��u��(K�e���E�t��7�B�T�ùc��8u_�$/��(bB�K��
��I�0���.B���	-1$���`C���(Jm��S	��se$�z�Ea�hJ�~���"Fi����ut�����Y��� HXY��c	������0�)��~��qI�,����k�~����\!f�Ѹ�t�?~���h����$.�S�S3�56GN:�?NH�x��C-�$��?m���8h��#s�n�)��)�#Dƚ�%���2晼8B�E�� �vK��6d1�Ѹ\4]��[����8]�!�Ѱ�¤)r�i�S�ix��J��?a�L�h�S���)-eIme-类񓮲^Z�5s{z���{�q��+�]
��[%�*�ub���պ��>+��WS�%�w���]�R�NJ3�س+Uyx����/of�iZ>�{�e9�l�j����y��?�?J��W��R]�N��ԓ����/�'V��}/��̮�o(T����eQ=��g?}��~���Z(P4��q�y��!�E��.~$'�ƀ��)��b@�!΄Rr����0��k�$��n�݄�:�E�0"�<�H���rYi�Ʒ���0�0Y���+�1�J2�]��o��� �V%~.�@�Ln������ޛ�#K���!M��2 H��.h%B\�։�.ss_���?/`�(HE�%l��Fa�)oz|c�_��aG����.dB��hf�Úe�@�~��9̚���)�4���>�f���/?�8kk
rO߿&��d6ƑÌ�����'�pQ̥]yg�y}���9߆r�JT�fs�'�9�Lќ���s\eĜ�\�se�"D�c"0!$�I@��HĐa�AJ�!Tѯ�!nH-B\��qi������֍���
�ь)��%+iLtl�HR i4):Մ,�kt!i���)��)	���V8F� R¤0%&h�leѶo �H�C"�a\{���H��\t���C�1�P`Q �LtMd2�1Xa�[�"0S�1҆����)��4d.04h�R
$�"�ЃX��HF����I�`Ё���
�楎ht$Z�֧�]*�b��A�5Yy�<��p� 8�`GG�Ja�T��!����F�揍��Sj�fi��i�۶$Is[��n�ѹ��H�4h����!s����B�џ�h�<�ѭ�����֟�݈p6�0��������u��\��r�6	L���H@����oGo�{�$%�X0�fJe��aLC$p�A�r��n�у^sl�i!sZ	sZv°��7�2�5��r����t,��˦h��#�l�;at@��V�(B�!���~Ip԰7ϟ��x��O����8f��fP��
\�%��������;ۇ��p�,)M�Ғ�A�i��vp�HRC4��W[�?h,-�?F 0$'Y4|����]�!K���.�Y���fݔ�!1��?l殮�8:XQ1�sxs)�.�yQp��(�f�3S8p�4(B��Ϲ�����sD)�N�aċL�O�{��yt)��Һ�@��8o��A!��E#�	�I�.��ف�@@B�B	���ϙ`���R�Is$+)?sW����@�2��vJ��~0���?Mn�2�H�c� ���E~4P"$M1bX(E`iB	���:v�A�P�R�h �q"��XB�+�SM?�\4WhE�0X�@�R�
�.U R�h�����I�6C�1�b@�O����H��h��2��B4ٖ忥3�ncj�n���&���d0��)��,cB#1���L��M�%���>B�95���%�����D�iU�E��WȄQ�pH��� Ud�$�@�		��$�f��6��r�� ��G�Ab�"��ąb��)0����`A�
�������t�l�@���f��e�L��3Vr�Q9>��k+0A5pNd�dK���WCY�p�.�DJSF���R@�a0����`f�2�g1"D��<v���f6^!1�	M?�S��$l)��,4��
�CF4��CD)�)��0d"D�eXT#�H��B�K�}���Z�Zր     m� ��[@  6� UT��(���������1Ĝyҹ�ݤ��5�;2<"����\b�nέ���;6�r��7��w��&�⓷��e<ыq�&[�n����H,���s2�>UV��j�U�6m+�u_���}�l"�m�M�� a��6��c   ���S��m��m�[\     �� =�l�t���r�Im @    ��2      �   �n�cHI$0`�ㅴ� p  m  p�  ��� h�D��n m�@  ��m $��� H   p  6����  ݶ��z� ���m���H    [@ -�.�X�u�� h   �� �|     ��  m���C���	  H�I�l   �����k��#m�6\�@     6�    ,0m�ޠ������ 	�$�� ��  -�۶ ��  �I�`-�K����h  [@  �t��p��cc�zq#l4kgE��۶��  �pi6�m����m�UT�P U �m<�m��� 6� ݴ�רڶ��`p�F���Z�����ym��llG�4�K��@  /[�� �` �[me��mn�ඁ���u.H4P �N�i��l6Z   ��][��-� [C�(  �`i0˥���H : �\� H��`VjZ�*����Qv���6ϯ|�M���J��kd˭�jεrk��f�,�k˛P9n���6�rޤ��m� f��*ڇ�N��3�u'���P H�.���M�rU	��J�Pr
UU[P  ն����[F�Rid��ᴒ^H�:�N �u�[hA�m�M��'[��L�l�pR��Wtn��T�U����U�SWWKˇ]m*�q&�Zzt�f�8!�+i��l5ʵU)� Yj���n�e���$qĀ����� ��`���ib;v��6��	�t�=R��3�q@h�� .�m sm�Z��m���� z� -�Ӧ�gm>�O��P
�*�W5m �����	 	�V�^p���X[M��K�+�UUR�알ttA:�qUG%Rk6� N��a��ڪ�c�6]�
��T��A5�X�-T �UUаăj��R�6�iлmʻ=�T���UTt�N.T�Y:�]�`m�#mm�@��J�{A�^�*����5S�fҩj�Z�s�7�l� R��d]�[{/��O�}a��֝Z��C5_��}@��evj�3�9�`6���	uԵԵЩv��C��[٠��&�-ֲ6�$  9wM��"�[�i:  m� � �L $I�oK@	  ,�` �ml�$$m�7  ,%�tۯH�h��6�6����ր  �       �@K����;���&�k�,劶�    h��   ��@ H   � � %�[d�o'GH�G-�M\�� � :<� 7mmÜ���`z�e��`��f�[6����XsDd�f���z�ڗ)v��ݕj���Q�:�x�lswh���Oe��9����j�Ͷ^����Y��LY�� ��v�;qG|o���ꞡDԻ,��{j�]�x��Uv�ʺ��S����-��G�UUR���&�J���l ��6Z�J��Im �m�n�!,�^�a� $�d��l�%�5��� m�nٶ�sM��r@ �qp�ti��6�`	9��m�q�6�����dp��u��r�8 [5�	�6�x���-t[�n������pg��kj��1q͔z�m���Ur@ MU$�@q�2p�)�     hm�N��㦭�W\$v�q#�E����`9�-+=�qJ��A\�U�t���Ul�VQ��!=z��+����8�7Th�m�oeU.���
������l���КJ��ۅ������i4b�oI�ɥZ���j���7_����@@V��f�aY��T�~������&�%��J�B��ְPbu [g�5/WVͤ�٣�����j�tUg��j��Zګ��8q��4vt���(@4�:�5y�H�7WN�m��"���	g&����� ��]x����qN��� I}, q�[f��aF��:m��Zܧ7/��� �L�K�u�q����KeX����\.ۥSHmm�(�#t*.�A{����ha�h
u��-N.���"�<m�� m�UU[\��ۜ�L��l�['K4�&�ܐ$��pM۝л)���CP nû��̭�h3�ħz�W��dgP�aWg�ر�񙈶���P�U��!UZ��tJ�VV@��,�m2B�s@]^�kj��Cd�Vy���L��m��S�c�M�x�JH$[%�۰�] H9�Y$�   �	��"��K�șрl-��p      �%V�6m�(�l˳l��WK�
6 ;gVf��4P-��  ��n� 8�n��[l����m��Cm�H�x$  m� h  � $iz�Q,ݜ:E� p�[��P���qPH-�m����%�Pm��vKd�А�m� pH�5�@P#<��^����iV�m�MN�  $�i ��5�6ٶp��&�����*�&D
m�+,E�]5�d���h�m�Hk�gB���5*��I�I������qm�m�ٶͶ -��Y[U[mUp"��6�2�@�V��ݵ��h���[%�!���Y����ԍ^�23��^����U*ҭ@Um,qT�	t@x$h8�  ���e�d�I�s�m ��$,]�A�^Ѷ���RͫIZ�t��I�84�ݜl�!��V�6�� @ Wl�uոŞF�*��e����u�9��mc��f�n�gm�����U)-J�@mu��--������n� 4�ͮ �vq�t�6 �b{PS��v�2�a�l����5UVSd�� ��   i��@f�d��� }��U�UO+E���m  ��[Cm���A��Iζ��ݶ  m�m�8p��h �    p�C�����U\�=+\��â��ܡì�$H���@ � 6� �lH    շ���Jlpp[%  ��p �fݰ$kM����A&�g 6�&�� 	 m���Vj��Z܇�.n
�9�5�:]�z��(�	-�ִPm[  �� �`��d�h  	�-�[��` m� M+h�$ �$8j]=�;���H�9,�9[�Ā�� ���ۀq[$�}X  �P���O��K/�.X����?7�|�W+�ٶ����n�[t�yӵv՛d��C�� �A��RԯJ�r P $t�:�[Pm�f���� �n  -��m� 6�� �"�����[�$�h��m���`  ax�d�m�m���JP m�݅��p H-� �Cm�6�%��     � ���m�� �m��֛n�HĜ �b�	�m�[@m�a�6ۀm�l�77��m��[D�HlՖ$�6�D�l�AV�hH��@�9wI67m�  N�Ӌ3Pm�9m� ��q'nӘt� u�	��&�kӦ�������v$��p -�&	  $      ���ܫp�j8 �  H  �8 �-�$  ��-� � ��mKm	-�4@m�$ ���� I���[m����m  ���m�i ��,����mH ���� �lzJ ����t�h���m�%��-�mN��m� ��c���6Z���H�����Wm��*�x6��9���y�9F�a챌Q�*��/l�\�U�UJ�';���F�Foj�#��,� t��d��  k�I.v�$���  � �m�          �      [@6�      �`@����N�ě`     �     �m�  -� 6�   m�    �H � ��l  p �`    ���Z릖v���Ͷ  ��	V�
���.�*�����m u��	eId�d�`  7Nu�5��>�}z���Q��u��-�zm��i�0�0ֲ�����(��E�H�"�S��"'������#�@�^(��:f*F$"�U���A�D4��Gu��p1
�^(��A�DMl
mQ؛Q:��Ѐ� ��z�~
�z�?��Dj�vm�� O�"#S��T�#���U~b�Ă� "�$A�؉8 �'�b��V��Ez�+�G�t'�ɴ��ĀU�>��TL��*i"F��$ F,`� B(� H �
�� ���1L�P6�.ǂ(A �~@_ʃ�D�����:�&��(�2�=S኏�� (�8��N
������"t`����(��1[��N�EB?���a6�A�Z�,��x ��A�"��=C��p!�Tx��O���X$]#���*���� �F ~w{�߿=���UP����p%�ڽ���ۄzu�/KvzՄYʽ�W4b�b��!5UmmѺ�g(J�f�WE[*���]uR���;j��ZU8�CM�jj�n�\i��rG[5]��ir��옶��6՛.�b��,�
�T����l#Z�L����h�*{\�dtrYp�0�5�#�IE�6ń��Tn�]Y��8;y�2�B�nqb�w��@
��ܚ����ͅulV�b�s�%��V|/lFZ�k�8�����h���]��<�I�wZ� ��V浱���;M�q͖�#6��i��ާIn؈�y�ћ�n����-Cݻ8-Ի;=RZ�S!���$ f��M�efF��S*d3.���.y��4sf��q)���غC���+j7\�n�����Y�XN�n�ڌ�U<;^/�!C����)�k��gŰh�������N�u���AH���"g�u�:\�ݨ�L#nm�[5l�����#��*�*24��mZ��:%Pa9��R��v���s/6�[e:^C(̝��pZ�,�]y��xN����T�D��̗ H�Q��p��[l��4�Id���=t���Ft�X������nm0ns��S<��=dPp�G6!,��{9M�l�7�t������h��С* ��q��N���u�;m�j�1=9k��SOh�K��Y�)�'z	��ge��b�v8���.n)�`6��+:�nݹej4*U��[��s����v�[<�٬��fD6�L)�mXh�sV�y��.�[$e$7b7����]Iz��q*Ɲ%�\���Y"�g;����U\P�ͧa]����h@.�K�5WC���A>ۃ=��km�@�3ʚ6�eUj:{\gap���t��m�L�J��Ғ��.7Q`F�9m�^6^8W�p�5@UJ��U@mUU �\
�Ҭ��UTpT����Q�s��;6��Ѳ��������SD� ?�D� �ѣQ")?�M@��ȈB�q�(�k�'-�fY���絝f��pF[=@�z�3M�h���k�]YZ晏mʆĞH��F��	ճ�6���Z9:8��;���c���x/g!�Gd 8P��2Gn���%]�Dg<pv��ml�rM�A�me룎U\ӣ\q��;R��r[Ac&��d��+��:{>,������A>�y���m���vk�=y�m�Bq�f���{��w�{�����](�sWd���0�e�e������\c>So/.ɻ.v�`N��;��s�~ꎷ�_9�=�j��������~�����6S|\�\���$*�p6�g(P�$j��KV����<�`w���a"��J0BnU���vX�����Vw6�����Tn�Q�h�+I�x�:8� ��- �O��[�n�WV^f��9h�*@>2K@b��7�6��IH�Q��"j@�Z##�s̼X a����=NS��m[��8��!�EB�#�����X��n���U�s4�$u%��I*�>�3���� ��Q �T>�"����M���3�5X�۫�R���s�4��@;rb�9h�*@>2K@qhiZ��ptܦH�vq��W��z�����Y�����$⦫4�ݴI %��1�y���yF�R�@�Rn�t�)ӈ��cH�(�I�'mvi4�B:db-v7I�q)��`���:=�`b��`wj�;��Vh���uҌDqX�L@s�-��H�Ih�Ĩ�*B�!7��y�����X���@�� H��\@�����ܓ囮��f�N�	�d��NG��ͺ@>2K@;�1��� r�h�w�����@>2K@;�1��wv���M��H�ȔM��[Z(�M�����z��v-����rԄ\���#j(���N+n���U��ݺ�3��V����7M�d�G`{k\�BS&�v,�]Ӏl�u�zV�)7N"�;��Vt{��ś���<�`w���a"���!'k ���:�`��8�$���t�B+��(�?m��V��ZQQ�$ҌDqX�f 9㖀�"��$� ��w��[v͗;L{h�W���_h��W�,�
I���5�I%ze��p��.������-�EH�IhnL@t�\W��[�iF}�����"���- �ɖu�(9����(D����`:���L@t�-��H�c��4�(��b�X����M,�۫+�uXXV�(�7)�)�Z� �	(����[O� s��	>��� $�PX�bB!�,X0`[77��d�sGl�qM������K|nx �Ϝ�A��þ��9PTpBR�Pڷ,
ն:��vu�Q֪l�b.�rN�r���ɱ���m�m�5��k�w-�<�uW	��<���.���lFɩx��u���:k��t�Ƕ�gAV�@q�n��� 3�9v6Wy!�Ŏ�3��!!�MqN^�]��ݷKG3�mC��S�U�kg
�]�	2�:��˝���~��kY[L��=k�S���e���+��),p�h�	s�Ċ�)7	M�"�=���c����b��u=��n���J0I7*����V����U���u`qf�J*9)&�`�)"�5vL@zc����H]�ZG>1]m��n�[V^f��9h�T�u�%�5wu���m�DT�"���qX��`�M� ����Z� �.\���)���.:`InK�KDp�`�m�l65��+q��j�4mC�؋��-w�����@K�1��n*@t�>�^ˬ�F�4�2�WrN���o��AĈV�z!(Q�;����=��`�VV�kJ7M�d�G`wj�#qR�Z_I��nw�uy�j�$*�p9B�o�,�]Ӏ9�u�wj�;��U��JRR�Mʰ3�78%
:��~]>��^,�Z���1sȤ�]ZS؃T,���/��5Gll��Ij႗��6D��K`BvY����b�9h	�*@:������rU�݊ԓWu�yֹ�Q�"d�}� kz���]`��l�ڻ�TU�\���`��dDCKa)�	$�q�FT��X����nC.j��ܽ�,�3v�� %��+{�u`whx�Z(Ҕ��!�J�%��Zs��� MPK�����QSl'1m�ђ�8�ug�,�)�;b�t�m�%��s�g�9㖀���EH	|� :�H�H�6�����X�v��s�u�{k\�%
�=��]e�ڛ�7Awy�H�ߕ %��Zs��f�hrP���4'*��R����5��������'�5(���=.�V���ڢT�$u)	���ʹ� `���b71n����ϖ7/m/Og&��1�;��knP��f�i7'=]��\q��J�8�w���'���EH�� %��Z��o*�SqR"��`��3�%'N��5�ͺ�;�<`�q�)G>C74@K�1��� *@r��kF�ptܦH�vq�{�t�|H�/��]7(�v���2�9��ͺ�=�{ܮ����Iw&~���������6�+T�̣S&q!���3�cpV�.f��c�<`j36�g�l�7W3�tά�9�ӭ��x���:,k	5$7	۶�4G�������[��`����4���}��Iv\Ặ[��{vƗe�L�������d�%ۀ貌X�"΁�c�\;;��@@��ZS�È�,vڞ ���ɘx��ˬݧD��6�v#�;/���y�{������n�.\�g<h�rS/w�|���4Ƽ:x\>��	���){ہ��EĔ��q�K�{�+�I-Y4v�K�3W8�[�m�K��� ��T�@���$���;I%̙��I-ɶ�I%�3y\�Inm�)ۉ)$qԤ) �$�2f�q$�&�-/�|��7ܮq$��xv�K��-�E8H�9\�InM�ZI,���ĒՓGi$��5s�$��"�dPL�DP܈��Y]��s�%�����=��$��\�InM�ZI%�ϝk�������ӥ��&�:�=g�sN���=�R�t�-fy�;���Y�\��r��KVM������$���E�����\�I%�Z5��L�8;I%͙��tE�#@� $D���7�������m��_v�����2�Iq���	(85BC�s�%�6�i$��3W8�Z�h�$�6f�q$��%V�E)8(�$�E�����\�Ijɣ��\ٚ�Ēܛh��\ʹmF�*j N���KVM������$����ݶߏ������(�ޞ��f\�W	Z�I��qF�F]��AkM�����.����I4�
�z�g� �ɾ\�InM�ZI,���ĒՓGi$����(DS�������Krm��Iew7��$���;Iz��|�ĒK7�n%��@܈��Y]��s�%�&���h 	EV��EH��_V�@�����!.�p�����
R/�	�t?j.������A4�h²�!�S { h������M�XŃ�
ʡ���P D�F��8��� 0�xx N�?� 8��$���罙��I/l���In�G�8�Ȧ�q%������I.�o�8�[�m��S{Y��s�$��x<H�%6�"D��$�6f�q$�U�qI%���W8�Z�h�$����aY����Tr���:w4�ms]�n����zz��Z�<��۫t�l��3ÔBPpj��"�RK�=h��Y]��s�%�&��Iw�|�Ē�[*�	��Q�I��I%���W9�����~^��i$�����$���E���m��TF�*j N�r�Ē��S��\ٚ�Ēܛh��Y]��s�%�4
w"�8�R�;I%͙��I-�5+I%���W8��ܯ�����CJr�]���m��׼P�Ƣ������KrMJ�Ig���s�%��i$����$�<o:�юx��`8��:�Z����d[�ѻYl\�p٣��-V3,]z6V���?���KS�N�Isfj�KvMJ�In�G�8�Ȧ�9Ē��S��\ٚ�ĒݓR��Y]�ӜI$�4�IJJJRr'i$��5s�%�6�i$����8�Z��v�K��4"��j��"�Kvm��Iew/Nq$�=��$�6f�q$��*���Sq(�$�E�����\�Ij{��I.l�\�InʹZI/�������/a�K���#��]�A����
�b��q��۞�{x`H�1����P�[h�@ɂ��1�#�p�-�W7`�ዐ#]&�t�]��Ӵ��\�m�\�h��h��8xv������t���nJ��6��[$�7;��<,�R�Q����Z�����!z.*������7jw�4�����Wt�cV�w(:7%�>+$fѮR  �:yیv������׼���}v#fs�r��]�+��a�����O�iœ]�ɛ���y띚իD;I�ݥ���H�Ԓ�~�v�K�3W8�[�m�K:L��$���)܈Q��HM��$�2f�q$�f�-$�t���I-Ou;I%�ߖ�E)����#��I-ٶ�I%�&��KS�N�Iw&j�I,�J�n(�}7"-$�t�ӜI-Ou;I%ܙ��I-ٶ�I%�-pm��2ÜI-O5;I%ܙ��I-ɶ�I%�6��KP�m%R) ԧ)��G��Ι��yyתgj�֫��N.�:��Fxg��"�St)R���I%ܙ��I-ɶ�I%�6��}��Uw�%��ZI,u���EJP��\�InM�\���Y�oNq$�dԭ$�rf�q$��%Vԑ�n� i7i$����8�[�jV���������&zo�8�^����Is6�m*#p�@�%!�$���դ�����$���E����ޜ�In���IH㎢)���]ٚ�Ēܛh��Y]�ӜI-y5�I%��{�|��"i	Gֺ�]�PpωeĽ��,)h��ˇҬ����o��QJCqGC����RK�=h��Y]����Z�h�$�vf�q$�_'����Lh�D�K�$�_�q$�<��$�rf�q$��+I%�Tr4��55�����ݹ�m���ݼ�Tڵ���}r��+I%�6��K=a��MХJ�Q��$�rf�q	n=�V�K:m��$�����̭�I�**�p��8(P�'�g���Հ{^j�;ܕ��B"�RmҐ�N"4�7&�Y��Hp�ݒ�%H]7��;%v7I������2�3m ���s��@o^j�9�)m*$�� m
B���1���r���@I�
�%%�J���vq�z�U��7n�]�vw~[j)Hn(�9V�r��EH	|� �����S��r�f��6��DȬ���Xۘ���-;$�T�-nU�{�t(]������������زI�9����v�;��&�@m��Vye���m�~�s��'d��u�*@>�D2��(���4���ZvIh\�s&�nVԎ
F�IBC�X�%�s�������T�F�� �n+:f�X�4�9�5X{���;�����$�M�@�m #{�9h	�%�*@J�~~�ϖǇD9ӹҎj7�۶�P�C͔�u��
���*X���s��� n+N�VްA�l��X�cyM÷$���v8Fnz�N7W�r[ N��i"h�7���d�Q�5���{#�=r�{L>-��t�=F9���i��7
wM�ǧ�9��k�˲tW�.�rF;Gi���K�(���ݛ`��puZ귉�����&n��o�w{۽��$��Kꃲ�z��L{O$�6�\�WV�݀l�sl��l�nS��3�Uɺk�o�����K@>T����kn9Hn(�t�qX׺��u`nd���<�`�h��m�>��X� #{�9h	�%�:Q�([���rU��ɥ��y��޼�`gL۫;C�Ek%6��"z <��@N�- �qR7�@;�w쀖�Z�n{r%�;Y�D�u��Τ���K2SXµ��Y`�=u6�.���v��K@>T���x�=��~*&A*��Vtݺ��UQ��Ȅ��b*d�a� 듚�d����Z�m��Lݢ��h��&�`�l�=��p�"L������Ձ��
z�(�rJH��,��H	��*@N{�­m�mX�QP���7�5X�=�W �l�`wj�6�������"(���)K���Ѡ[G<���ke��l�
�g���vlfX8E�@܊��ۇ�� �l�`wj�7�5X�:Ƅ�7>�#������
&Mt�p�}8�v��J7(~TxjSdMJd����{�`oq�E���U_f6MBs� :�����mn�vn耝�Z�"�簰;�4�9�[�����M�`>$T������M� =1�@u9W��e.y��P/�&h�uu�8�7����<�S��=�]���l�r�j@6�o`���- ��Rɴ��Q$䔑M�X̚X׺��u`nd��I��J�FT�*��� �Wt�⛜>I}]��OŁ��v�8E�CNEa殺�}Ӏ6�۶��*Q
* I"�H"bX�(@R���G�?:��Ӏ{�S�O�RMXU\A�E`fd���Uf���������77h��"��&�H�4�1�����Q�s�3�O���-l��9�-�����o��6DԦB8p׾V5�:=���Uu�����
��?(��*J��8�M�t%#һ� m����t}T��u�|TN*I�0bn+p~�7vه�B����N�W�N���H	QM�H�=_R���`w^�X�np:K��N ����vUt�,���?mk�菡B���O��} ���rA:��0R,B '�$K���:
�'��H�k	�(Tj�-H�e�%����Д�c�Qec5��xa�@B�6/��(�i)
B��,
+� A � ���.+����)!�j@�D ��!�
H���H-�a��T �b�`D!��[��!A�!0d�(��"��J'ЁԜ#4�9���!o|w��`���R@�mHԄI%Te%#d!1AB���Z�Z�i᠌�:# ��Dc��$�xA�BffP�T�X�� `�"D�?-"��$bB&|ə!�sP�BX�"�LU>H@��BIZ�"1H2�)O����~@H[x{M�]&��%�S���=s\ȳ����sW/V��SvBJ*��k����D5*�*Å�[����)U�e��UJ*��pT�BX�j@&���$ F��n$n�\��۶���ڣ)i���l\MӚe[Kr�	�+�S[��,��*�qԵ"ܐ�I-�*�ڎ;\2r�]n�Dӳ���Ʈ�@��8��w.��+���im9�ؖV��0:�bv���-��Fn{q�8TTu#�Y��d�k��\�f�q14���.��,`7�pt��c[�]M����v7�q<���ݱ��v�����G9��[u:�=�n�<p�Ko�  -���i'���[@�ʷvz�t4jkU$�d��A86'�b�=�u��b۞��M���@2�ӗ���s�H��y0�K<�\q֮��䄡ۣAݻ[�u�cc8����Ӄ�P�*�6]�P]��2�I�6AaN�mt�|�����,�ݶ�=�1�] �JƬ+��s���=��+��(SaW��]َ8���R���f���۫0q�og7Ivz�ն�=���q���6+P!�m]�X�u)�I�CF��қys�m��˩v��r���]T�m,&ɟX��ֳ�L$��b��C�g��Ӻ;f�ĝ�kq�md����[�䅮H�UR8�H�[F�\Q�7fM��7f��鶘�H6j ����\��8u���d^��:m�4ml�WI����`[H1�i)��`z6��6�-'0��m����є'u�g�-KYZ�g�)@�=�;����㉦k��ҹ%[<Şt/]f�Y5�m��So��m&M;��Ү���U ��Km�T8Yf�[&�&�Y&$�jt�6�X:��4��o7dW�m�P���
Vڶ�`U���%w�}�0At*=��U�mժi@S�۞(�<��x�4�*���` �����m�Z� -�v��I�V�e���*��
��[v�hX�ꃖ��pZ�d��δ�X�����h�tJ�r����P������A\P�J&�uQ�D�">ұkT��i"��.�.��i\>.nOk�n-{�;#>;�E�qӶx[��j�����%�T�hd'g9�0]��qs���'��	��=�ڹ�j���v�3�'�7ADj�3m���5��[s{;��!��.�@jӋQ�.������H����t�3Z�`��kg�4�6M�Hօ�[��˥��w�~�v}~�/���<��i�j��
��{'&�tp.�!]��WGw�����$��kUsv|u�Ӏo��`�wВ�!�g�����J!M7"�3���D}	*�����W}8�79�ɼ���I����d��۾�s&�}�EV�_}83�`ȧ(eM�SsSqJ��9B�v�p�}8�oB����`���p�%Jn��r+z���ӻ�����mk����;�w��l�n]�5��i�9�F�.lnץח!�z�����b�'d>�r%�bX�����"X�%�}��[ND�,K�u�]�"X�%���]�"X�%���ܞ���h����fh�r%�bX��ﵴ�>{H�P�y�,N�_~�ND�,K�k޻ND�,K�N��ӑ?�*dK���l���֤���WZֶ��bX�'�׿�ӑ,K�����ӑ,K��Ӿ��Kı/�ﵴ�Kı>��K�F�*8��qH_���Gԏ�W��}v��bX�'~���"X�%�}�}��"X��2'��?�ӑ,K���пܹ�&kE�2�fkWiȖ%�bw��p�r%�bX��w��r%�bX����m9ı,O}���9ĳ�oq������G�(���v�ƫ�^�4mkW'nŞ}p֛(�Y�j�s�]��cfi�ɚѴ�Kı/�ﵴ�Kı?w]��r%�bX��]��r%�bX��w�6��bX�'~5}	�Fd�˧55�ͧ"X�%����ӑ,K����ӑ,K��ݾ��Kı=�wٴ�O� r�D�)���Y�f�h�%��j�9ı,O����iȖ%�bw��p�r%�C��R�ș��iȖ%�b~���Kı?wG�MK�kX]d�mֶ��bX�'~���"X�%���}�ND�,K�u�]�"X�BX����n!"�ur8E�w$��B����(@�'��&��	ϳ�ݧ�X�%���m9ı,N�;�ND�,K��ߵl.4�F�'M�:)�.�b2,R�<=n��L��z����O|f{V��cuS�r%�bX�����9ı,O}�siȖ%�bw��p�r%�bX���ٴ�Kı>���殲�P�j�h�k5v��bX�'�����Kı;��m9ı,Og{��r%�bX�����9ı,O��/�sRMa�C,&k5��Kı;��m9ı,Og{��r%�bX�����9ı,O}�siȖ%�b}�k�'�Z̹�34�ɚѴ�Kı=��iȖ%�b~���Kı=��ͧ"X�ȜH(������{�iȖ%�b}��OI�2�f]7R�Y��Kı?w]��r%�bX1�������Kı?��?�m9ı,Og{��r%�bX�������7�:�қ/:w6��q66�]�����q��*�un�������nk�^�L֮ӑ,K���{�iȖ%�b{ݞ��Kı;��iȖ%�b����_�RB����w"ɱU�.�����r%�bX��g�m9�R9"X���fӑ,K�����v��bX�'�׽v��bX�'�k��&����K�
e��iȖ%�b{;�fӑ,K��u�]�"X�%���]�"X�%��v{�ӑ,K��}���Z��kY�kY��Kı=�w�iȖ%�b{�{�iȖ%�b{ݞ��Kı=��iȖ%�b{��߮��SS5�ՆkY���Kı=����Kı=��p�r%�bX���ٴ�Kı=�w�iȖ%�bs����WK��u�u�lI$;s�Sq��j�Oc���z�t�l�[�۵�t<��b}ۭ��[���v��!��n��&����Nx�.��u�ݏgFqu/H�s-�s{c\K�g�s����u/Fp9嶔���=`�R}���nv��,�s�yīۚ��Q�6X��w/�݌gM���Ż:k:�x�>.����V���ܖx�;�K����w��|�Ӳ=l��ꗭuD/sk�V��O�s:7k-��]�U�����k�v}��߻�{��,N�vp�r%�bX���ٴ�Kı=�w�a� ���Q,K�����ND�,K��k�٭f\љ�sWSZ6��bX�'���m9�Pc�2%���{��9ı,O�����9ı,O{��6��bX�'~Ծ���іk2麗Zͧ"X�%��뾻ND�,K�k޻ND�,K����"X�%���}�ND�,K�|w�Y�\ֲf�f�v��bX�'�׽v��bX�'���ND�,K���6��bX�'����9ı,O���R��&�L�3WiȖ%�b{ݞ��Kİ�#��{�6��X�%���{��9ı,O}�z�9ı,N�����&Ν�ʯb鑸�V]����}�)�V�.�%a�C��JB;9tm�: �V�u�fw�Kı?���ͧ"X�%��뾻ND�,K�k޻ND�,K����"X�%��{l��Z�35�,ֵ��r%�bX����4��ș�����ӑ,K���=�iȖ%�b{;�fӑ?�Dʙ����/�.������3Z�]�"X�%���]�"X�%��v{�ӑ,K��w�ͧ"X�%��뾻ND�,K���r�.j܄�fkWiȖ%��2'�����iȖ%�bg���ND�,K��}v��bX�3"w��iȖ%�bw���I���Fh�4�]Mh�r%�bX���ٴ�Kı=�w�iȖ%�b{�{�iȖ%�b{ݞ��Kı=����`�	������rՋ��9Rq��c:NdGn�N�t�v�xö��ғu.��ND�,K��}v��bX�'�׽v��bX�'���ND�,K���6��bX�%>��ڗYLֵ3$���]�"X�%���]�!�)"dK�����ӑ,K���{�6��bX�'����9ı,N���ԳXMjL�fj�9ı,N�;�ND�,K���6��c��� #]D�O��}v��bX�'��}v��bX�'�k��&���][��fh�r%�bX���ٴ�Kı?w]��r%�bX��^��r%�`*0Ȟ����i����$/�����T�ҕE��d.D�,K�u�]�"X�%���]�"X�%�߻}�iȖ%�b{;�fӑ,Kľ�﬚�)3RIn�W5uB�c�z4��
��GZ��Fu*К���xWp�9Pq�)��p���#�G����r%�bX�};�ND�,K���6<�bX�'﻿M�"X�%���o�sP�5�!1����r%�bX�}��N@lK��w�ͧ"X�%���ߦӑ,K�����ӑ?��9"X��&��f�њ%�2Y�Ѵ�Kı?���ͧ"X�%�����iȖbX��^��r%�bX�}��ND�,K�j_I=fɫ��n�ֳiȖ%�b~�w��Kı=����Kı>���6��bX�S�Q"��\����fӑ,Kħ���u3&�%���6��bX�'�׽v��bX�'�v��ӑ,K��w�ͧ"X�%���ߦӑ,K��Z�����_HDP*M��N|������է:�<���m(�un��%v7�:r��Г%���O�,K��}�m9ı,Og{��r%�bX����m9ı,O}�z�9ı,O��I�CZ։r�d�.\Ѵ�Kı=��iȖ%�b}�w��Kı?{^��r%�bX����6����TȖ'���$3�$֤˭aL�ֵ�ND�,K����ӑ,K���{�iȖ?ȩ��?����iȖ%�b{=���r%�bX���/�us4j]d4Y�]jm9ı,O�׽v��bX�'����"X�%���}�ND�,K�w~�ND�,K���r�s5s)1˚��r%�bX��w�6��bX�'s��m9ı,N���m9ı,O}��m9ı,Ni��}���ؒ^�G��ۑΠ7X3J�`�������:���3Je���$�YGJ��7Wgt
���[�c�����q8�P;W�
�I���F	��g͹��6G�r�m�<�$gk�:o&�wo[qɂ�F�!q�]@zJ�6k��^��v��m���αòtK2v�컛^u�M��<�YV:�[s6¼���l�y�N��v����`+��sM���}���Ge]����mip��h�n�H�	m�s�۵n4���jB�+����a��3]���d�,K�����r%�bX�����r%�bX�����r%�bX��w�6��bX�'~5|C�h�M\�jR�Y��Kı;�w��Kı=�����2%�bv{��ӑ,K���{�6��bX�%;Ӿu�WV�֤�MkSiȖ%�b{�o�iȖ%�b{��p�r%�bX���ٴ�Kı;�w��Kı;��C�R�a5�2YsSiȖ%�b{��p�r%�bX���ٴ�Kı;�w��Kı=����Kı?w^'�f�K��$�ff��"X�%���}�ND�,K�w~�ND�,K�k��ND�,K�v��ӑ,K�� ;��������f���k��|��X+�R\ލu��9��R���#:ti'gd��ݻ@ߏw�{��Y�;�o�m9ı,O}���9ı,O}��ND�,K��}�ND�,iVg�/qD� �*"�$/���#�BX��^��r�b%uQ,L�w�6��bX�'���m9ı,O�w~�ND�,K���.�Y�jj�a35���Kı>�w�6��bX�'���m9ı,O�w~�ND�,K�k��ND�,K�&���jau%��kZ6��bX�'���6��bX�'﻿M�"X�%���]�"X�%��Ӿ��Kı;���F�j�kP��Zͧ"X�%�����iȖ%�b{�{�iȖ%�b}��m9ı,Og{��r%�bX�����j[e���i7����j�x��ٹs�����@�uF�jFR�Yc�պtB���+}��oq���=����Kı>�w�6��bX�'���l?� '�ı>��6��bX�'���!�u,�Z�%���ND�,K�w��Kı=��iȖ%�b~����r%�bX��^��r4��R>��hyQQ8��&�!W"X�%���}�ND�,K��ߦӑ,`�~�	�B�$��A#!O��O� I�I h��$�F$ ���$H��0E�B������2����?��v���$H@ �T2$$�$!X�F2#h_��q"D���X3��P�)�b�n�~���4���(�V"���?`(�� ∛_��N�_v�9ı,G��2����$.��r�Uut�ɭkY��Kı?}��m9ı,O}�z�9ı,O��ߦӑ,K��w�ͧ"X�%��ޥ�5�4kVk!��֦ӑ,K�����ӑ,K�����m9ı,Og{��r%��2&D�����r%�bX�����L��Y�cDg-�F�u�+�K�k�<����ܷv"�+q��j�C�.K��tؿ{��g�����p�r%�bX���ٴ�Kı?w���r%�bX��^��r%�bX��5�%��R\�Iuu�iȖ%�b{��ӑ,K�����iȖ%�b{�{�iȖ%�b}�o�m9ı,N�j���Ѭ�����]k6��bX�'��~�ND�,K�k޻ND��dL����p�r%�bX���fӑ,K����ɭe�u�,2�SiȖ%�b{�{�iȖ%�b}�o�m9ı,Og{��r%�`VH����m9ı,O����f�i3RL�3WiȖ%�b}�o�m9ı,Og{��r%�bX����m9ı,O}�z�9ı,N����.��tj��]����sin)|َ��Mϣ%om�*�m�t������'��Dn�����{��7����ͧ"X�%���ߦӑ,K�����ӑ,K����p�r%�bX�Ӿ��5&�Y�0ɭkY��Kı?}��m9ı,O}�z�9ı,O����"X�%���}�ND�,K�z���\֡�YXdֵ6��bX�'�׽v��bX�'�v��iȖ%�b{;�fӑ,K�����iȖ%�b}����֋5�I�\&f�v��bY��2'{����Kı?���ͧ"X�%���ߦӑ,K�����ӑ,K��/��.������M�"X�%���}�ND�,K�{�M�"X�%���]�"X�%��ݻ��r%�bX�#��`PT�֢�1
TB���UZ$�J�MMR�흫��mŔj 9z,b:I��1�c�r\�ѷ]f܅]qۮ{�gcs�0�6`zw��Np�J���l�Ÿ�5,m��m��m��]m<e$ؓ%[���ވ��ݸ�;[������K�ò��A�NÝ�WO��/?�����۶��t�:�ͱ�v{��M�u��h䪇3�S�3�Jo"C�]]+�UT�:	�}�w���>���qڃ���j�^B��c�L����c�	9F�j�ṋ[����L5���Ժ�u=ı,Oｿ��Kı=����Kı>��~�ND�,K���6��bX�'��h�Mk.[�Ia�Z�ND�,K�k޻ND�,K�w��Kı=��iȖ%�b~�w��Kı?wG}!��B�3RKnf�ӑ,K�����m9ı,Og{��r%�bX����m9ı,O}�z�9ı,O��d�&����.�K�.�6��bX�'���m9ı,O���6��bX�'�׽v��bX�'�v��iȖ%�b_N�غʲ�n�*.��!~!I
HRB�y�'"X�%���]�"X�%��ݻ��r%�bX���ٴ�Kı=�n�_�@�yc4#Ѹ竩b�ޛ�GX.�����+���um G#[��ѹթ��Kı=����Kı>�w~�ND�,K���6��bX�'﻿M�"X�%����s�Z,ֵ&�p����r%�bX�}ۿM�!@�ʃ�D�K�=���r%�bX���ߦӑ,K�����ӑ,K����p���3Ff�R�ֶ��bX�'���m9ı,O�w~�ND�,K�k޻ND�,K�}ͧ"X�%�߉�Rzj��5���Ժ�m9Ĳ���}��A=�{�bH$�����M�$OD�w�ͧ"X�%��=�=5���e֤��֦ӑ,K�����ӑ,K����siȖ%�b{;�fӑ,K���w��Kı/����-�u�Dn�v�3i���n�������K�]�ܹkՠ���q��m�ۓf� �����oq�����siȖ%�b{;�fӑ,K���w��Kı=����Kı��j<���GJ0M���}H���#����6��bX�'﻿M�"X�%���]�"X�%��Ӿ�ӑ,KƗ��Ez�QӦI#���ԏ�R��ߦӑ,K�����ӑ,`�� �(PѸ������iȖ%�b}��iȖ%�bw�R��˚5�.�X�3WiȖ%�b{�{�iȖ%�bw����r%�bX���ٴ�Kı>���Kı>��,�f�]\�5Md����r%�bX����6��bX�'���m9ı,O��z�9ı,O}��m9ı,G��ݽ������[�W���:Q�]���&�zH�b-��{k���FjJ�k�ا��34d���~�bX�'���m9ı,O��z�9ı,O}��m9ı,N�{~�ND�,K�^���՘k3Y,պ�m9ı,O��z�9ı,O}��m9ı,N�{~��'�ı?���ͧ"X�%������ ���_���Gԏ�W����9ı,N�{~�ND�,K���6��bX�'�׽v��bX�'���.���eՓ-����Kı;���m9ı,Og{��r%�bX�w^��r%�`q���"k9�]�"X����n�Q�I����/���#�ı=��iȖ%�b}�{�iȖ%�b{�{�iȖ%�bw����r%��{����� yB�)�@�ny��9�mNa��k��8��Y.ݸ���H��e_RSZ���0ɭkY��Kı>���Kı=����Kı;��p��"X�'�{�ٴ�Kı=��_�k.k&��CV:���r%�bX���z�9��L�b{����ӑ,K��{�ٴ�Kı>���Kı3=�C�r��1�"���ԏ�R>;��p�r%�bX���ٴ�Kı>���Kı?{^��r%�bX�����XL�342f�m9ı,N�{��r%�bX�w^��r%�bX���z�9ı,N�{�6��bX�'�&�I�[��k3Y�u��r%�bX�w^��r%�bX���z�9ı,N�{�6��bX�'s��m9ı,L xb#�IX����߶�a�۝��3&r�:݀����kh����;Q�٭f|�8�zz▵��{ax����G�6с*�J���YgN���!O����d#Ud���t��Q�ζ]p��R��ˎM�y8�'k:L������>�l0�{{d�베�R��5��}�qFq�h��'���CH�t�ٸ�5غ'@U�UcS����+�{��'^~.��q�T��N�͡#$�jN�c^�����)Ah�hڭ�]qs�Y\��������,K������Kı;��p�r%�bX���ٴ�Kı>���Kı?��I.���eՙ.f�ӑ,K��g��i�����,O����iȖ%�bw����ND�,K�k޻ND�,K��e�&����&�%�34m9ı,Og{��r%�bX�w^��r%�bX��^��r%�bX����m9ı,K��V�R��֮��MkZͧ"X�%��u�]�"X�%���]�"X�%���{�ӑ,K��w�ͧ"X�%�߽K�k.k&��SY���r%�bX���z�9ı,O���ND�,K���6��bX�'{�z�9ı,Ow�̶Od�i�%D�A��Q��َ���@�Ƚ(6-�(�7�G�e.�#G�����oq��{�ӑ,K��w�ͧ"X�%���޻��&D�,O����v��bX�'�I�a/��L�.h3.Mh�r%�bX���ٴ�< �DJ�&�X��o�iȖ%�b~����Kı>��6��bX�'�&�I�[��k3Y�u��r%�bX����Kı=����Kı>���m9ı,Og{��r%�bX�þ0�֦ap֤�WZ��r%�bX��^��r%�bX�{��6��bX�'���m9ı,N�^��r%�bX��;�I3X�!�Vd���ND�,K�xߦӑ,K��������~�bX�'�����Kı=����Kı:w�{R�2CF�\���mmV\�t�:�]��:��l�v��Vmst;O��õla��{�[�o%���}�ND�,K�׽v��bX�'�׽v��bX�'��M�"X�%�};�_jf���uL2kZ�m9ı,N�^��r%�bX��^��r%�bX�{��6��bX�'���m9ı,O��/�������Mds3WiȖ%�b{�{�iȖ%�b}���r%��` �MD��{�6��bX�'����v��bX�'�y���h�tfSY	��]�"X�%���o�iȖ%�b{;�fӑ,K��u�]�"X���L����M�"X�%���k�K��&h����56��bX�'���m9ı,N�^��r%�bX��^��r%�bX�{��6��bX�'����9��K8�-��\�\�Q�J�&A�oe��z�6k�a�0��	ډG��Ŋͧ"X�%���޻ND�,K�k޻ND�,K��o�iȖ%�b{;�fӑ,K��񇮵.K��%��֮ӑ,K�����Ӑı>��6��bX�'���m9ı,N�^��r%�bX��;�I5�5-&jL�3WiȖ%�b}�M�m9ı,Og{��r%�X�'�׽v��bX�'�׽v��bX�'����j��5��d�fLѴ�K�lOg{��r%�bX�w^��r%�bX��^��r%�`i8(�G�A(U���\���iȖ%�b_��Wڙ���k)��ֵ�ND�,K��޻ND�,K}����Kı>���6��bX�+������$)!I
YϨ(������<�
�XY��,��ֶ�5���	�%h�[p)�I���s�>�~����x�=����Kı>���6��bX�'���l9ı,O��z�9ı,O��}ˬՆk%��3Z�ND�,K�zo�i�(��bX���ٴ�Kı>���Kı=����Kı;�5�%��Lԗ4��56��bX�'���m9ı,O��z�9������ӑ,K���7��Kı;�5�OkY��k2麗Zͧ"X�*)"w����ND�,K�����ND�,K��ߦӑ,K���6��bX�'��O\�sW4f�&��]�"X�%���]�"X�%��|o�iȖ%�b{;�fӑ,K�����ӑ,K��h�80!���ȑ �/�~�"�9�@11v0��!��� ��	��1aFFI� ��D�b�"B0 F+	$`�r�ᅅ�e%�q�C���-%D�ā$�2S�� � A��
�F A�)",�6�z�8#A�U ҥu'w�k@��m��U��f�����uOcw=]�ag*G��Z���A��Ǳ�rն�[lp)2�UJ�*��P ���W��Qnhr���T�����UU��`H �9�M��&�(6�jQm <�k[I��� d��*�OU8�1k�<��]v��nۇ��J:Y�UFVs�ϥ�qȲ�u�<l�6�]��%n��ێ�1��3gb���쳣dk��p�{�X^���z^�Pe�s�����k��d;#�\AvC�l��kB�kE��9���3�Xc�+���A�g�qe7e��Ur@��uY^�Чndyu���s��}Zk[��l�9̊���P���ړ9��9���m ��m�h�Rx��M�e{l�F\�����<�M��V���ջy�n����-�ɎW$	Lz9��-'=]zݎƜ��*�j��9k�18W��Jv��7e�+��q�;gi8B�6طIt�1�9y���<c.; �]�ʽ�j��Q�v㰜mt\��*��vy@�a���E�D�=�h�%�<���q��m� xn�h��kn��'T�<���n^�5��:��
�.x×��k�u�fs7^]���U*��*%�>��l�KYɮ�X�#pzAmm��7e`���P�d٢�i�;��v��v4a��i&e�k��
��݇C.�iZ��ђ���J(�ӎ]��uN���6Ú�����׎m9�[5Pkr��[�X6��nY]+��$��X�/�mGjt��S.v�"]J��L5���*����מۛ��C�{]iډ��mi0л�d�S�s�viV����Xq)�ur�����G�4�u�6�	oluGT�&������t�j��jBF����L�-O ֒U�TLl!D�OU�T��
`C��RB�pۣ��J��֕`(v�T�T�<�H ���5�Vl�l]�T� *�ez�]�Z�g���\B�x�KA�j̹�5�L4L��v�=WK��.� +�?�m��^vk)uùs@��n��bB��OYn�(0y{��I���e�Au����s�L�S�B�Ж9��<�n����E����U��u�$C�&[��a$���7b�m����ܤ=�y�N��8������#=gnr/f�b��l�i�Ѯٶ�-٘���X�ܻp=9�q�������ۧ�Ⱥ؉���sn��u�.�  �v��J�t����)���%
j�z�
�qך��[d�N���TQ�5p�)�nI�a�l��,���O�X�%��xߦӑ,K��w�ͧ"X�%��u�]���L�bX�;���_�RB���݋�t��\܅�Ѵ�Kı=��iȖ%�bw=�fӑ,K�����ӑ,K��{�ӑUlKľ��\񚚺ֲ�Y�kY��Kı;��iȖ%�b{�{�iȖ%�bw�=�iȖ%�b{;�fӑ,K����}�L4kY5�k#n��ND�,lO}�z�9ı,N���m9ı,Og{��r%�`����}�ND�,K���r�5a��a�$�֮ӑ,K��{�ӑ,K��w�ͧ"X�%���}�ND�,K�k޻ND�,K����?�h�)�c���g<Z:\=�[Vl&�tAX�&w\d+Yn*���{�Gk�q9n�5�i�%�bX���fӑ,K��{�ͧ"X�%���]�"X�%��t��"X�%�߉�R{5�sf]7R�Y��Kı>��� �:@�mQ���&�X��˴�Kı>���6��bX�'���m9���,O�=��\�sW4f�&��]�"X�%���]�"X�%��|o�iȖbX���ٴ�Kı>���Kı?wޒkXj[&jK.f�ӑ,K���7��Kı=��iȖ%�b}�{�iȖ%�b{�{�iȖ����Tu$��(�	ԅ���`{���.�~�;�M,n�T|�Ҕl��W���-�2U�90V�F���6�5���h��/�"�5N�$���=�`o[s�y���B������`���st8ԅFS��޽���H�x�,-�;��U��ߖڎ|���FP܊�~�gvnI������h���(�Wsr�� ���9E��WU5V����X��7Հ9�Հ?;f��u`ghz��M�mO���Ź��}����>ŀ9�u�=��B��D���u��IO\$z2i���B]���L�����u�������T��oΛ�*@Knb�s�� ��]�hYy�hT������ ��>�JL���r��L����j�`-�`/]aЦ{z��>ŀn��`���t�$vq�{�f䟾�vnO�"	���~�,�)z�%
B�)��`ovi`{[ŀu��� �Ir��I
�d�X���m�����[��n���Q�Xۜ1v��͘�]!�fg�t��t�~$��R ��@s�-:l�wF��WU5V����X �]�(�
&Mu�6s�K�������`ghz��m��"U����np�l��}|`7׀j���)� � �E`ovi`w&� F��1�rQ[��]�hYw� {��w��RJ��M	�,R(=��� �S�u������E��;�V���Nn��.���;^����k�wj�cD�2��ɷ���\����6H�S��nr ��+�pC )��)[ib-�Vn/m��+����s����a�R�'�y��k�7��X'��yM���St�նu�tb]<����w%��R�[�'GF�!:����f��m�x9�Fg�X*Vz���{�����w�G�r$A�	;>XK�ۨ�����vc(�zt:7l;GGM���a��m��e���9~�}O� 8�Sd�R6�(���Ź��UURG��Ł����73e��#�◭E)8��H|�� ??��@8�{���h�L@{2�	Е��]��U�n{���<�`ovi`fQ���:#iJ�Q�+ ��%������������}ձ��0��/o*6������i^�'��vëvJPM�\�K�A��-z���>n��l�<���P�J^�?{ߥ��W�0��(rA:D�G`ovi�2y�ŀu����9BIL�R�r*G
T��BN{g�Vf�w]��٥��䥪����`��,9(�������V ����0M�_l$���N�$���=�`z��Gog���� �u� ��t�K��S[^XË���u�������f8nû/��+���i%)8�R�Mϣ*�`ovi`{]� s��Q�C]wN�ܤ���RpQ�sf���vq���3��_B�UF�t��-R���+WUV`OwՀ{i���(W
���,wv��΃�F�N�j|�v�%��� ��� ��� s�� r���"D�St�I��{����}��r���{��6���j��$��Ϯ�f���{���䴗��@#[�.C�n�'n1�)(�D�Nqp�z��ՙ���=���� �?yX피�*�	AFMU��묅���L��p����,�
Ъ�����]�7uR�IwwX����'d���"��� 8U�D��NEI�n+UR�OyX��Հ�u��(JQj�ڶ� �jG�v����\������,�}}�W�~�+z�U�f�[D��m1"���U���m�WkP��@6̇c��Ξ�f���T8F
!ʩQ�*�ՙ���=�`o^��f��V�?:=m8&�3n�q����r*@Knb�}�W�W��ʽ��� �7T�I��_� ����z[�����?)Z��THT�!7���r�-�;w]��(I)���7]��E�VMқ��j�`w]`.����>u�Ӏy�ŀbK��B���@뺛�E31u6X�0ljٖ,����g&ڝ����=H�QǙ�;Œ��s���U�uJ�ǎ��1X\A��4��Zsa6�e;����4iu�h��7�1�r��˭����2e6�sOn�l9E�<���볘�%�<�[	�y\ik2�\L�P'7c�[x��<;����	������X`��U�:mlE�L�@,F6�������wJ�}M���E�۫�s1���K�
M��/[���n�j�۱0�����	U�n�����V �M����:[��77�'h��"�
I�`s^���}2>}� r�V�s�$�Ow);.IM9�����Y����V5������4F��R�rU���� �ֹ�?:np9%
|��,���6�r���ǚ�k�V3f�,�vV�TS�*(�J�I�g�u�Ӓ{�q�u9�mq��9�c�fI�h�c�>���v�Ԩ��Jb$�>�?yX=��s㘀�]9(�ܭ�.�R[s5w$��wf�� �N�� ��Հ~t���D��ڞ�Ywjn���Uk r�V���%�Ϻ�� �o���_l*H(��H�G`bz� ���5�Ł�J">��Eu�}X�ߊN�TSqQ
I�`s^�?|�C�~�}X����7�WM*]דa��Z���]���n:�y���:-�I���s����{̳��-���;��o�@Knb�Ih	�%�<�bh�'*�F�,Y���_}�$f�yX��/�A������G�Q�	��Y7u�{i�����TB[+�H�`h��ȡ)�J@�(4	����m(�u J*~�Ȅb0�H�����fZHVK%,m�,-�aSD�1�	�`	D,X1�d$4�LI"�#q�.h	* �+�	m�Uj�8 ��Ȣ�QH"W�`nBP�b"!���0�k���@���.��ws��P�)���5��9��`wj�9J�v����	�����%�}}�W�������>�~������yv�܀���\q3������o��8�m���F���Gl�C�H��%(�	�p-�;�z�Wﾪ������ޥ��B4Jt�$v��X�78��`w]g%��7=�C�E)P�TTq���+7$ۘ�w�����Ы��
�Uw8���8�:[��6^��H ���������IΓ�MwI�19U)��`j��`b��`o^�3ri`+�／	W	�B�j�x�r]u֨��h^'���q�m���;�Z��?��U},t\J2JMϜ��y~��`orK@8�	m�@K�0%�mѹ{XIwuu�?Ss�
&G���:[��6^�ϡ)��S�B��W"�	&�� |���>IDL���;k�p=�&�jJ$�!9�UU����3_t����|�Q:�8�;��+.��Qj��wu�{i��>JQ�}��}~,Y��U{�ɾ�6:�G%%*eY�L����\��1>��..���Ϡ<kj����k=F|��ݕGh<r��ܶkt�Z��rNW����ZBc<j��X����ўٵ`v��}��s�e���ik�=��+l7gb��d����S��ݷm�X+�Ҝ��m��=��؜WKӵ��u��'m맚D*��<h�����V��p�^�p)�Ѷz�j�g�u�-ak7��غ5g[�^�[�q�*�Fn^[����w��}�E�V!YeUπ���N�v��믒\A����＊��E!
�����]� s�� ��s�?Ss��СE6{h�~��	�T�F�`~^��`b��`~�Oyp��t�4�"JUV������!D)u�Հv�t�z�`�5��5��QP���H�v����BP�＼���`>n���~&�6����793;i�J��۪���`��m�D7�絛�K�F��/3m��H	m�@;�1;$�s%�q�n%!7*�ՙ��RT��>�(EC�"os/��nI�g���mՀi�K�IR6Jt�$vϛ����:"B��}� �o� ��5��8QP��v����u�9�u�В��u�Հ{�I�wa77d*R�Vw&��=�>�=�`o^�6�Jۊ�J(�8�Tb�mԘz��p´ڻA�ڹ�3���]-�k�����EH�,Y��]�v�(P�Ho;� zԎ
�]���E����I�	�%�:=�<r���ꯒ<�|��T@���H�v������fJ���8ϛ��B��"�	&���!D�<� �O� ���a����{����H�F��F^n���@;�1;$�G�A<*��������5e�e̴Ѭ�����f��L6wd��y5ʹ�q�eF��Lܷb����y3q�$�%:C�.�忿;z�U��ɥ���U���T֢��NT)7��M�t%
d�w�ΟN�s�%�Fg�Hw%JC�B��Vw�Ł�Z��S:�����8�T̢��Z]�����<r���@N�-_�b�Q �D� ⫿����ރ���	��H���V������}|`k\�k\�Wb\�p�^��:���*��Y��	+�7(U��X�@�ú^��bn1������9�<�ـ=�s�DB^��}X��������Bn+��Kq�g�� �M�8�������"��*i@� ׾VWq@3�1X��,M�_mBJ��S�9"�;�5X׻8�v�P�)�o� {�"�*iJ'4��o7m;$��� #�-�3U���%��	H�MӢ4Ҧ8ۑKku�eU�3���U���+�7u�t�#u������
��˱�m�����l�u�����;c�s�+f�V�A��X�1Eq�\E�v䭇��Lf�z���$��%y_^6Ⴡm�.Y��j�1�K��^
�Ծ��1�&wF�����V�GaͯX6��2�;�����ڕ!����Z��L� �`+��2=\����~���58��\���^� x���;8l���Sc�]��b���{�ݏ��?W\f�sa��l������<r��K@gq�lC�NU#p�7j�;�\������3�(J&G�]H�MD��8����{�`o^��UU}�%���`{^�X�5��Q�RH���G���߳� ���0��8����7h�C"M�`s6i`nֹ�=��pΛ��}2�K��;iȑ��{<����6rl\;���N[8�k�^$;M��{���q7�b.Ӱ'!�=�����<�`o^�9��V��*Ѓ����!���y��ڪ���P�%vvW~�ϻ ����nEq�B�NT�Ȭ��,f�Ձ��U��y���w~N�Hr(P�rC舄��!D%[�}�}��N�s�ʪZ�i`gq�lC�NU#����p�D(��D(���O����n���F����(6�s�$s�=zA�9�ڭ�8N��6��P�-˫�l'kf����ٷ{���Zt� <�T���Uf��* RA$qXݚ_�IDD��݋ �O� �ֹ�?)Z��DI��BN3v���y��_}�W�� �	���� t҃�'�B^�]wӀ>w�~{jF3wSt�p,�ͤx�9㖀�69.�M�ZQ	%:C�+��U���Т">~���}� {Z� ~��x�8tnX�v�y��]n��.ѭv�\���FG�8����&�x��ͻt�]� ���o ���D(��C]?+3��;��!�EI�3v��{Z� �ֹ���>P�S#�$�첦�f�!]���7�����8}�D�秋��]X����)҃S�E$���8��0��,�
!$��
!r�IE�~ΜҟR:�	��I��@>����1�@s�- ����� ���}q4�������j�Ϝt�M���׫tQr3��ۊ�������O�<��`��8����$�_�=��l�e#�"��!7*��}[�|��}8�Z� ���ϔ%	D���S�n%%:MI�������`s7n���Vwuq�B�8QQ�"��Q�Ӏy�b�7ծp>��J"sf�X��RT!��9��H��9㖀��-uuU_z�ﮗ�#A�H0W�Et�X1H��0�YP@�SH�w��r�B�����IL�\�������Ml7U6�b��8�H.�X :��g�����ɿ?�۳n�$N�����ש��9��CՍ���`�v�cvm�8�ݍ푇�ն���\*�nf�X
�[�M�*Ҽ �RF�ndV8)^,�F��k�b� Hs-;$�Iۅr�����3l�Jk�+;[1R�,ʁC�J��"��x���cn�1�ϕ�sq�SUUr3�o'B:[�����:ɛe�^�=;V�vm�Kq���6G��9��H�q�d�;g�piσPv|���2�R��6Hs�]��g�DHD{n��҈�@n�<������Cv���!�͔�^�a]�����w/IWg[u�m�9U��c&�z0��P�.�2<� �@e��z��fz�䋒� ��we��H�-�ջn���r�Z v��z���qۢϳ�v�Rz���3.9��&�g�������]�*%ǡÞۍ�4�P�N�����70c����@�6'�V��
Sn��݀x����8�G���gH<
h�\<��\��K�@�݄Ur�ڮ����v���ō�-����-�<<[��r����Aq�"���E��<-�p��Nӻm�NT�p��g�i��
b9�--֬i�s���z�kC���`�.��Z��� @$�7�Ű�i��1� U�����cj�D
�Bv����d�ےY'�͓�:bAj �7k1;v�T��t� ���v2��7;��(��I���!��.����ck`f�lq*&x�i�\�R��Z��Km+��U��'�S�ᠸ:vmts(��Ge�)	D��v}a�68k��!Uӹ�.��:�nۻ9�����;�vU�ԯ�u�3Os,������U���ԛB⺛6屔�ݷD�Wg������hK6vw8�x�fRW���T:�(T��V���v7�H��e�d��](N9�4�BZ��	�++deXv�TR���@-��Z͊fͱJ��� T�� � 5�܇Ӹ����%�&i�Zֵi�u�k��ү�q�mo��@ �EO��,DTv�Q��@�5>�4af��5�K��K��v��;� ]@�y�g@kp�ڳ[q�9����6v��rt(�0H��[���y���m[*�y�ݲE���0�.ڞ��<�[C9N'n��GT�*���jܤm��wIWU�bmv��m��B�.]��8� �9��呆:���:t����Fӻg����UuK%�[�)z�G�6��)��ےk�`���������{���?��t�8x�Om���W��㶢����$i�ΔҤ�.��,�I$J4��*G%X��Vq����(�Q�Cϻ��9GZ�6T�Q��hx�=1�@yȩ ������H���rA#���� <�T�}�Z�9hUԒ��ͻUT]%]���O�w�=�Ӏ{k\�J_(I$�{����jzQeՓu&�W���}�Z�9hLr�r.�m���/���#u��U�ڌ�m9@��\qWh�v��Fu��r�/�j��������_�|Q�Q:��5$\5�y���7��P�%�A�>��t�.��	�������@zc���UWن9 �-��U������#3}�v�ISc��9VOߕ c���Z���e��"Q��QR9*�μ�`wj�9��p:!$�|��,W*r�
�Jl���7wP��@g��~����5������Q��aR��S`�R�l�Ԛ<�gc���Wa����z�d�*�,v?��{�����o���!�.����+��u`�����׾ViW��*G����H9 �j�9hLr������zQ�D�Jq�0bnU�no���y۹�  0K��ݻ�s��f�qn�U"mԧJG$�;�5X��8�o�D$�IEW>��}"�h�r*T�r+��U��ݺ��l�;�5X���麔�I�"��R7o�]�"�[x�ɨ�TG6��Y�NK�j��q��7�jD�68�C���;��Հgse��y����`gq�NU#���5���9h9/�Wc���Q�r�(5>tI%�������g仾�Հno����]IH؂]\��k���� 7���P�(ȏ���+��wh��Q�E`s6*@��<r���%_<���.�x쨦��k�K��*�����|�v�rr�]-��Tvˢ�/B�6�&�g~$��@s�-�Z�EH\�K����)ґ�,��W�#�{�`w{�`�]�%	)��r�,�w3%�
UT����}8�o�������X�o�ڐ)0qP�#���l��9�x�=1�@>vXfٹ3V�������9D$������]�9�{�rM� E s_N������f��s0�x�0�7�u�gn+p��:�.�ڀ�9�����S����l�,b���p�k��^`,@�J��I-�ڣnq�o��'*ｽ�^����Ծ^���e:�lףDp�3=lEج%�N޷�!!֭�]�ں�y6�H�Sc�,�=6���.9z.X7m�ZB�6i�8#M�g�l�Ŧ�h�IU���(p���֡nƐ.��dv���J�Zڶ�x�e���;�V�5�R�&��%(��I0׾V5�h9 �j]9�M���7v�7sm�Z�EH��Z��wh�uPq�E`s7n�;�,��V5��z��8�ay�H��Z�����[��EGRSL��H�q�������5 3�\(��+~/F�vy��ŠY��^z�uy��z�֗�;Y*̙�yh�	:D��D��M�"�9�5Xr*@��<r��}x�w�2��D�wW8�oZP��Q*�����xu���U����J�'*��7i >sP��@zc���R�i�XF
&�҉$�;�5Xך�9 �j ���n�f�������-�"���9㖀o���ʹ����=��KN�]��j�؁�%m��5Z��
�^�8tF�3L�7m�"���9㖀��-νTGD����`����H�{�`w^�X�۫�u�����r�8����<�`sj�S����_?�u�۫ �f�;�HwN�H(�t���<��@yȩ y��x�;��'jJbt�TS��`s7n���,��V1�+0����9R�|u�&��L=v�R�W-�D�Y�*�!(��C�$�r��FJ�'*���V�͖q���U��ͺ�;[O�JMO�E$�9�5^��3��������U����$�ҍ��H؂G��{����������-�rV���殊����}�{�������_v�O�(�Q�T�Q���EF������Z�ܓ���:Qr�����`��`sj�9�5X�۫�W՞�Tx��q�#n.�]{>�H�1C�fC�.�w<sl�fF���T�}��Z��dMS���$�|��Xx�<�T�<���*�U���W�VaW�����-��H��@sǪ�_}UI�x�ړ�&���;��*@nj�9h<r��a��EF� �f���U��y����}��|x��{%�-�˧F��P��@y㖀�R �sP��?`_�<�ڴ�v<`z����ewm-�b&��l�s���h��j�4C��nm��t�I��\�0�՚r��C��ȴ�\�X�t��Z��lӮ��%���u�}���cf�ۇ�7��>9ﱭ��##�M����<��C:�s��nχ��c]su4���tպ�9���x`#6�g�Q��q�:6�]j������iA��v�  �Zy�q���{����q���٬]g	��îܭ�mYgq�x�w��V9@�a��\�s�v�1�����ΟN� ~�w�P���w�viV��B:%"8��"�;��V��9㖀��-�ssk6R���`��`sj��U�����o|��X�~��8�Q����
nR�{�<r���@y�� yɨ�RV*V�UwT��*�pmk��	DGВ����^ ����=��p�/
�Ub���gv^�6� �v��X��Jq�	���Z�sk�lCN�OM��ۮ�����R �sP��@y㖀�ae\Ѭ�4�f�nI9�����q�h⦑	[������B��>���;��pf����ꯒ2�OUbQ
6�Ң�X�������|��`�����;��M]�Q!wW8��IV�wӀo}�, �k��Z� ��6�e�Zͳ,��@yȩ >sP��@zc�`fj@Vӫ��1��RD�(y%�È}4R��n{hy�n'	��AC�A�����}�q�rR�������;�5Xך�f�ՁŚ��*7T����I`s�-�Z�EH�}U_]��ԇl%�M�r+�{�`s7n�6sn���)!�$XD�X$H�� B�d�B¬�Q(1"�б�,R$�bH,���`F(�������\"D���!HP��˄��aR��X�
AFI��hE]�)	QN0B�� F*�0��( ��T�c(`@a$E�I #HFH���n&�a H�Ef"x�̈́�zp�!S�KBe%�����"EDR4�H?
�"~�&�aYqHē#	0���!(&
������~bP�R��bT��f(ƤZ�jB��@�$�����`��� $?C
R�H��0���#BQ�Hij$A�48���lNĨ	@W�p!��A����A�|���ǹ���^j�;��ԟ	�5MG�[ŀ�w�{k\�tDD�����Q�D��r���`��`wj�?:�8�o�D(���\�M%S3��it�=A4n�$�9;%�ś�yx۵Gj��[�ss|�5Dj��H��Q$�5ͭs�~��|�G������:��*wwp��ʹ�9h9 �j��V)V���PG��V3v��7��IL�Ӏ{�������Wv���j�`|�DL�}x�}85��˙�ʰ:�R�EF� r�wuwx����腿g}>{�`�vX�[q�EI��DpjS��H�9�"���_f�-z �����!մx��v��2�3v���<�T�9�ǚ���C�'�86��rH�f��tB��z��t�pε�}���L�։Q�NU$��s},c�V5���u`v��*5�)B��J$��(�;}8��N�u�����
��e(��8�k�V��y��� =}x�s�	BKK�D��*b-�V�5!���w<w����U������[9�i^`u�`7v�^�l
sڝ8��8kE[Q=��˲�ӹ�H���m���nО��F�Y��^!�6�n�e��sS�����m#�L��m�Gm�!�l��,�z����6�{e65g���+֮?�-�rv�T�T jvK9��e�����.��/1��y��Xm�s���̇Z��x94i3=R������~���r��ST	I��#�V��j�{��q��b�0�rt�%��mn'Y�N�Di%��RU����X��x�s����q|����zx#�T����9V ��@y㖀��-���˹tTn(�#�Xǚ�k�V{ﾪ�.����77����턨�pt��ݴ�9h9 ��Z�t�ڑ�D)�rH�f�Ձ�ﾭɾ\5�y��3q=Pn����-�1Z8B:u��o]A�� )�\[�'B�B�*4'*�q�V.��9hLr�r*@uJ�tL.�j]dӢkZ�䟾ϻw�E� "~�+��gN�݋ ?n�������$R�8�9�5X�۫?���U�Gw},׾V)Vn�* #�hr+�!(�>�� <�^�s�~��8��
Ў9RJ#&�X36Xǚ�c�V3v����6*I��R�B�6v����呶xo&�t�vrvm�S�ub�b諭��P��8�QL��p׾��ֹ�?n�_$�~�<�^ ��J��q��c���<�~������k <�^�s�$�ɽ�"�n�Sw%��U���o�`�n�	%�"#�o��:�U����h��R�]���S>}׀y���=��pۯ�v��*5��5>����<�`~��o��o�`�n��Q��]HEv]���ŵ�8I�f�}��8�w��sصl4u�L�(��z��qdY�l�~��d�h9 95��U�J4N�ڔ��V3v��}Iwޖk�+��U���(�9R@����<���9h�UUۙ?Z������TN!�S�9,=��ߕ������sﻳrGJ��T� b5*# D���P(oy�w��9���������9��y���UU��r������y������c��"IF�����Ć����;Ln�h{T���ҩ�����x�'
�*%QG �ﮬ�&�<��@s{�L�+6�0�ڭ��ݤ�&�=�%�9����H���Q�P��J��`s�uX̶a��M�ذ{� �e9�YS5uvXn���� ;�T�<���$���ݢ
JH��IB��sn�O�u��]Ӏ{vـ|��"!-��*=���@g�����.�;fM<nx ��`y�I�nm��t���K�nЛ��1��J �q�E�ڎ۰��]{+�C0��ɸ='�׶��V0�vxj:�����{o��ok������u�ú+uو6�
4۝3�5��e�G��ݕP��7:�Y��.mk)"g�V�-v�;�3�d��#�˦�q�����ٸu���n2	%SZf��\�^=�{�~g���v�eA������2�=����^�׵�����˝r3��EH��$i/K���O����?�{o���O~��}� ��'�*'��)�ܖ:�U�U$g��X�� �����{�R�(�����h��;�T�I�vIh4�"�����#���sn�;�,ަ��N����b;$�&�U�u����<���$�<r��*@w������N4�!ӈaC˓bMs���z��ƛHN��L���:��8�I����n�=�%�9㖀�qW諾`t���V��F��D ��`wj�V��*@���$�U�J4��T�Q�E`s7n���,�URY�|�׾V;���r��F$��a���~��2~�<r�r*@z�.TrP��)��q���U��ݺ�f�;�R�D�����ª��Z%�o��t�:ĳs�n�]ɠ��;d�����.�JQ9�C��f��9��V�ݛ\A��n�Fڎ6�Sj�!�ʹ7����<r���_����7h+}h�&ەR�rU�w}�`wݻ�U∐�@X��@W��}UI9�V�|��*��0��˸�]]���8�k�����%���~�_��W�(�S��H�;��<�T�I�x�'=�ɻ�!O$��L%�T�s, ^��e��Mۆc����L3�e�;Z�X�8�pf��<�T�I�x�:c���M%�G���r���/��ԑ�����{�`s7n�,�iEG%��S7P��@s�-�"��&�z�pu*R�Ϛ�V���l�+��lܒs��[��WpJ�O�
a���qX����cj�!��9��V�&�9㖀�Z�eE�f� ��uŰ���BF�c.�Iv{u۰�r�`t@�uf�V2Wd�F�U�����������mk��Z���>�X���G��8ڟJ �;�5_�׾Vw޺��,�5Q��j���G�s�~��a�P�F���t�l��v�))A�A!ȬfmՀ:�5�Z�9htЅ����F`Yw�H�I�<r�1�@y��ܓ���H� �V1�V-	P� D+JăB$BI#
A,�ZBP�T �`#&���2�� �B)�4��B,��#�!�)�UK�Z�FES�E��κ����Z����G� �F2�0�	B�H� �H�b� �B �(@�ă�� @�a �`�*B B!]���
�>(&�\,�a���ֵ�kV�k0�]��S���neH�5�]�Gk�T�i�h�-����!���D�յ������U@�UtTj��<�ղ�9�ͺ}5 �TpT����imm[Pm�h :C���ĚN�2��t�xض��7dz�ݴ�gA��L�=�г5�[�;@G�.�}uZ�W���7�ʵg2)�Z	�fN�:��h�����@�� �7��vyu�N$L�l�pu�����k���	s�6{l&��s�p� �9ux��N#������ے���+g�:�uԛn�6"c�tp<ڻk)��v,�&{k,��n���[��v�NSgv�S�)�;ѴuA��i��e@t[UN�Yed�t��۹@��A��X؉�����T��ӈn��\.�4s�O=�i/m�7ۥiL#�u��ݳW]*J�ڳ[uIl�!��l�mh����i�\�Y��h�uOc����o=P2j�:��'[����6�
����;q��NQǋ����m��09��RKʹ��q��u�Eu��!7f�fM�@�x���t(���]`���	GA܀��V(�G�U�p��Uv����w֗-b���ەp!���.ހ-�%]P�ݻq�vs� �2�3 m�TlX�V�"��i��|i��1 [T�C��r`"��c·A�m()��ۆ�nVI�`A�p�bT%�;�t�R�Pl�h�Q r2�U�71�l4l�e�pp�f&&�K�6X�v�����^Ob�c�B��6eԖs 4���S��i�p�#�����]]s��(]�g��ѧmR�����Ͷԫ��,�q�y�\ݍI�<Ԫ��)�6�Rn�Gl�{�l]�Z���R�Ր��;���G\mJK���]S`.,�4���3Ӆ��&w�0`����lf�
���뮋3���;�ݺ[�&nm���m�m�oP	-��q�ֆ՛f��[J 
�P������C&������U�n�F�d5�����D( �G��PB$U�U�� h�@ý�q������w����N
Q��VL�uƐݎI�rpP�%��;R�r�u�l�fGͱ�vՌ�����O���cq��n�:��T��i������֎�=��v.�u�=�8������A9 �Gl�nc#lu��=��,cm���rk������qv7[�<a�h�~e���m�{['���� �v��vsH��s��2ˬݮ�-���1��-��� ���w��uY�v��Ҹ�Ӯ��[�kP�I�v��Gt��v9j+��x�����3��nJ9E2JNO�{�+��U��ͺ����;��pu*T�DAʹLr�n*@�5�Z�_}_RG��=n9I�&�R�+��]X�n��(��g]>�]>�u(y$Dm9U*7%Xtݖq���V��|��, ��\���
����YWx����J�}?���ŀ�`nf�A"'PB����n ۀ�0�]K���!b]�ꂙ!���;�;W;v����@s�-�"� ��c�Vii�D��6F$9��ݺ��BJ=�
���x�}8�k���#���䨤��!7*�6�ޖ<r�1�@yȩ 8\(���XԥLpNK�T�f�X�V3v���wvX��R������E`t�-�"����<r��ř�һ�㌗���FAc<-����9���,��*�tM����6����#�sL|������<r�}^�s'�@IF�=j$�iʩQ�*��ջ,��V<r�r*@R������ߴ&�Zܓ���n䟻�v�`�E �����R�Jju�Xɭ� '�P�M�R�W$�]\�}�T���p�ŀl�n�mk��Sm
�J��ؐ�V3v���K��� �{�`w^j�35#��i&cMH��I�y%��/�%;��th�{VАP�Po�.���2���&�pF{���<�`w^j�9��Vh�����5)SpnKg��}��7���ϱ`'��{�"�D��R|"�q�ך��m՟�-F{��՞�9��S�)�q
*�5ww8D�>��;=׀l���Ȉ_US��ڪ�������Q%NUJ�7i ��5��Lr�r*@O����${�/<��[�kUNד]��2�wl�m���fn��cm��;N:�R���u��Lr�r*@;:M@����j���T����`s7n�Gwe��y��|��������Jrw8�v,d�w�В�S<���3�|����B8�'!7*��wf�#�Lr�ȩ�p�Q[��Y��u��f�9�@t�-�����U��:�Ku�7�q	8h �]�[�u*���m�K��*�ӽv#8gA�GH���\�N@1s!���ް���������;��ь��E�ٞ-t�>���i L�ם	���bx��[�������;6v(���<�g�������vѺP�jtql ����7sl�mևc��2n�Q�v�5J�Du���q!\�@ �U��"�=+~��������Ga��l��l�r�!���Μ�2�gO^$F�fxnĲ��ōI2�|�4�{_�X��V#����٥��ݢ��R��QQ)��77mg�drou����<�\����ؔM9U*7%X���sf�u�sv��;[K�R���@#���6��#�R��j ��Dڍ�RTE$9��U���u`b;�,͚XU����!�&�h*I�U,����a8�<e�I�g�5֎���e��qQ9J�d��ȸ�޺�1ݖ��,��V�jUmF���FMʰ6O7yIBQ�
!Uݳ ��\�wn�,�iEG%jR��ܖ��1�@G"������[w�[��V^h��Z9 �&�76i`swiS�*A��U�qX�*@;:M@G6��r�^�� �:6�{����]�j�>��\�8n�y�3S\⣢��]s�͎�I�y���f�Z�����g�%2}Kʏ�U)������Ł�y���EHgI�et�,ݭ��ʻ0:�8��`�DrQ
"%TB��t��׀~}l�<�6�dթ[�me���T�t���l�4�7�R�jJJ%!7*�2�������ȩ �܅���D;�W/VⱵX�XӚ.z�(�ҵc�6��:��-�X�n��!s�r��h����ȩ :�5 ��ŭDD���M8XܚX��V���`nl����v�DT�⦇������P͂�9h�%��ҙ���J��]�IB�k{� ���'��ݻ�� F
��,X��1	���ađ�@��0�,��$)Ec�!$V� �R!HH#0�O,�V��(BHȅzb|�ݙ�`/)�C���M�qhWWx�l�<�\�[ŀ��9BP�:���w��B����Z콣5�t�2ۗV�q��h]�Nf]vX�����3����wg�}]��[ŀ���e��U����Jl���ݺ�Ě��l��@Hͪ�Vn�����Uk 7�w�=v�:g]>��z�����TrQMԥNF9,͚ 9㖀�EH�&�8X��v�.�7������@G"� ��PN��vnI���*���۾浬u�	:�L�jQ���^6���@�[Vqqn]������p6,�ݱA����6�8�6qs��/5����7��r�['E��+��W7��ͷa$�	м�'c�$�����Vۛ�;	���Ρ��(.�#v���m��m��'Qg�Y���F-v1�+��{�.�[g<ٷJ���;�ͮ�JlnͰu歺dӡ�q7[���nkWZ��K������?g�}$�\$h	a��F�V����%\�7��ʽN�jݖ�	�7F��;>i�������H�&�#�<r��%�6:�MʥM�*�3��76i`wj�77n��RA��k��"SJO�rX��� 9㖀�EH�&�9�utT�V��2]ف�J��o� �݋ 5y���
!O>�0�ςɫ�uH�JB�� z�,�JZ���>�,��V�3mQ�T���T���9�t�Q��ea����;�m����7)#�Fq+��GpS��!7+���s���]� ��]XYFS~�6�N��ܖ���TBIdZP�"Tyֹ�<��������$no�W�&�p��r+����r*@�M@s�-$���R$��#���n�Xtݖq���U�w#��nU:��V ��P��@s�-�"�t�o����$�!��ki�^������nN�c�K��n��M�RpWa{O�'^�[7P��@s�-�"� ��P3]#MTr��8���V3v��3��;�5XU��⨘F*�p��, �����0�����B@����H��%J�)) ����@b�d�BH�F�,�:X	�$JF0*D��@� J�*�1BH4*��R�Bm�Y�b]п)�� X|J>HE�� 1X�T���@#��[@���p���O�!̀~ �K��D�h�Q͠@��	)R1�4B�0�@HF! EFA0QtD�ol0!)`F�0�3� -�+�X	�I	�����oF���� F,�FD�`Y ��C�!��!�1��*�j,qF�u@~E0T�?:�@���8|���T6���@u���n��{����*�䤢Q�r�?�Q�^�׀k�Ӏ{k\���X��-(���Jt�c���<�`wj�9��V.��`w�"}$H���=1�q^cDOs�d��,��A!fv��F!��CBp�r+��U��ݺ�1uf�}��|���=j�%F�ϳw6�r*@;�sP��@y㖽��V֪=#��ܪTے�X����Z�����R��*���̽�CowP��@y㖀�R}G�,����<������krI��ΏH6A�r�H�9�5X�۫Vl�;�5X�{	$QH�7`ι�gg��0[7��'����X�4i���XEG
EJ�"E`s7n�]Y���<�`sj�9�J��9(PQ�����w��9㖀��-�"���:���EG%Ҕ�8Ԓ��{�`y㖀�R�[��|�f,3p����,�7m�Z�EH}nj��7jJB��T?��+��u�l�u���� ���pJ!*A�@�O��l��2h�\i��5\�l�]��+Ze���l;��ܻGE�;]���}���L��-��Z�ɣ1��k�z엧h;s@�W!�U�JU���;s�<����mӳ�ۉ��)��^�cK&�͋8�'m�&:��ۨ��v�^&���60ԉ���k.�!�Xӹ�6�l��Zt���t:�٤ZFRؖቌ�UmUTd@�Q]�����w~����l�7.�M�@�x!.;]�f7b�8���@GR-c],Ա����MD&�RCNJ��������`s^j�;��Vki�]*R��O�I`;�1�Z����sPp!F�6A�r�"��ך��m՟ĵb�KV{����)*P�9����sP�L@zc���f�l%5���`b;�,]�v5���u`v�iMT&�*R��J[�n�ݎ�XX�N���흎�Z��T��)z)�ab�$���)�q�%������<Ԁ������1`n���t\.�Y�'��ݻ�hh�
iT4@K�������`}=׀l���5��'�H�P�r8��mՁ��l�1wu�ך�+uQ�:��R���6��sP�L@zc��������MT/
��#S��pY�;��Z�����P��7M��,���0��6�"�	��M��f�y�%���(��r��H�vu������P�L@u�p۽۬��2��7m��H�I�}& :<�{�$fi*�)Mģ&�XW{�nI�����pt��@] )�ռ�畁��]XY�Ҋ�JMҔ�M�����1�@tqR u�j;�!�	�qQHM�`w^j�;� �&����|�,�̭�·6�3;���p-ҝ�f��;�ǳb���C$���8��)��G��ͺ�Ě�w�b�9hԗFM�ڻ�ګ�/7i >$�����@t{u`v��*���#S�D�.��9h�*@�5�L�0�tͫ7ow��@tqR |I�*��BDw7�s7$��玲֭fVV��h�*@�5 ��q��V�eyʉ6)���G����D��٪���qY;=���R��6L�H8�7�����ޖ.���U��ͺ�8�E�$���)�P�L@s�-��H�&�=);A Rn*)	����Vw6��RF��KV{���n�v��N$�f�m�:8� :�5 ��Lr�V��u)F�SCRJ�����X�k�ͼX��B��IBc��A<���u�r�+��1�v���������×�jo=kh{h�mv�o�}i�r�u��tg�(+�έ�v�c��Ҏ{K=;[6��psY�.糵�����t<��z�]���[�b�б���M�iZ��]Gv�c�v�If:n"F�����չ�Wc;a�r�);���ǚ�q�s�S��s��틆���[l�ѫ��%�un�����TN���' W���]e��s��L5��*�U�����bTv�Ί�2�g������j}(�����y�ך���ՀewvX_��pl�������~�I ]&��1�Q�fn�U*W@HU��m��^n�舯�վ�3�|���Ul$R��F�ͤ ���& :c���"�1�ZQQ�I4�%7%��7]��nZ�����PԸ��2��3t�9���ڍ������rݺ��Pm%q]�d D��N*$
nEJ������`y�� 5y�興� ��V���\չ	�kY��'���7"��hD��m�TH�	U`������׀l���=��pSrd�IUjIV.��`b��`wj�;��Vki�h�C�����ۓ��@t�R�\����ҍu ��"E#�;�5X�۫V�1f�?W���'ʃR�(���s�sMS��_}�2�	9�rΩL�s�[Z:vkp&�N)7N��t���V.��`b��;�5X�d��H�7�,�ͤ��5 �Ɉx�:H�����T�P�#�ܖ,�v�s���*�q��,N�����Ձ�W�X��'j�S��T�	��x�:H� :�5 �ɈI,2ܟ	ęC�#�����XWwe��7]��y��7���7N$�N�Jt���-Ō��II�;g��FH�j�狄���.*q�T��45$� ���1f�;�5X�۫���P�J"(���uw�l�u���*�z�� ��ŀl�nXZQ�6�#�H�vu��������5 �Ɉ��w�u�At�]�D$��w~X�{� ����T@�
�$�Ic�w���j�	��Q�r�][��ś���<�`wwn����U
 q��M�"����b�z�5tlЉi$�ft�2I�^�����
Tn�Q�q�%��7]��y��y���Q�A��u��D�Ij��U՗����Z�������&X��ܩ�a"�S��`wwn���5 �Ɉx�8@7wkj����/wi �M@;rb�9h�]X�����(ȣ��9,Y��䖼}>�Z�=?�v��P�"B���*����*���*�EQW��E_�U��*���@�XAP�T$BEd�T �P #P�B,B
DT"�AP�
@T"(B
�*�B(�P�+P���BEBB, ��?�*����*����*�TU���� EQW�E_�U�TU��EQW��E_�U*�������)��t�;��8( ���0���  �0   ��   t �P�   &� ����      � � $E�D
�J��
�T�� �(�jT�&�� E�@�

I
�PR��a�  9Ҩt  �PP33��Q��E�B#C�� f����7{��짧s�	;>����oX�����:�z��;�� jV ��@����  gҊ  �f( Q��U�}B��%�3�}7`T[�Cϰs ����P}����6������w{���{ȇ�f:�9n`u ψ�@h@P�v���z.� S�� f�@�P�� M��)(@�� i�4�@KX �� w,�`5!e�s@���R�� )wp�������P �  � n�t  �@)J B�5E:p:P6e ���ǧ��j��"�70	��g;h���u6�j]o��  �0	�� ftT�[��T
�l�r{�s� =�
(���  ��C�Y��t��� Ҋ,-lk���vQ���f�>���� �X>�� ������F�M��d�=��An�9��w`u��p   '芟��)P  "x�T�M   '�T��T @���MM�U*   ��T���F�  DHSeJ��ѐh�>D��?������_�����t���u��E^����TUҨ�*��**��TU�tAQV (���S��a ��� �ƿ�7BcX���C��H���($U����K� 7p�!p�����'6).Ml�� ~]�k����!p�@��&o��!���m1e�Wd*ⰹ�$�i��K�Q���w���DN|IsJm�x���\ѵ�X5HWP�%F4�I.8��+�!q@��������F�0X\�_���/���y��R$���42�F�B)+`[��
e7
bT�(@�����SO0�HJA�Ѵ S4Cd�1X�c��J���٫�H���0�&|�1��@�X�FL�)���	�59����1#|�����
C3&2�q�(B���!q��2�"��� �D��aI�@��`0u��4� ��0�Sp���h	�܂�37��� ���3�F��(J\�g0t#F%H~0*;�E�B Q"�%AĂ`$���G	;�?l�����x���F�;��+��!�Hh��.�,%d%%�8K'!��v}��3�$�/�o��B*�7���;n�Y�	f��LII�Ě3I���cr�1�e��%u���N�j��q�p��%�T�Ӷ5�N|�bE!F$bA���bC��\��-�2�>�g2}������ߡL\XGf�L5b��4�aX����0X#��u�s�뙠��kf���W0a�!w�o5ȕ�0"Tcg���i)��0��B��\N���%�KS.fɓPoE8��a��޲nF,I'#�f��:?~�.o�v�1�XO߱�$t�cL ��H�)�Fs\&_�s|�2i��!.R)��,�n�#
K!$��hv�c��D��+�5�?'T�WC ��%��4��b�
(8�d�F]NO��7�D��H�S����S��.M�᠍Ms�|���I ��XB �B$P8�
���50H5Ht'�:�!i�"��H;8r�-qQ 1p!���^s���^&�k
f��?@Ʌ�����)��4�m~0�̑��2�����������?.R0� Da�hd�B����cG��H$k/�8ƙ��� ��F�-0�?��0�豀P�Q"���� �a�ũ���@�� P��%CCq�.6
��@�b����E�U�P�P�AH�����$)��k	��D �$A�E��@�ƴF�#G�q�a��J�*T�RX�aF @��0��r�.�B��)(�P��*aXP�sD+���.oRw?l��Mh���N��\�}�3q�9�6u>h��y�׿D���>Y��~N�6��e��YB/-~t���<�WOz��<g#֗�߿~�[[��(���}�N�����m"1��HR��gy��������&���5�i�I�*F$+*�ō&j��5,JG�ޯ���}HU�N��\�#�7�Im��6dݟ���Ģa�\"CC��Q�B- �bCP���X�(0je�M5�?��"6��Id�,�ʐ-0$�)BR0�ЃB�c  E�20�H0?(l��Ƨ�������
�a���B�*p��a)�+)0��?����m�	IT�ap%�\�\���E�Q��+(B��
��d���lxb�Y�B�IbH�LelɌ�
��c.$a����4��I�Z@���B�Ѷ\4���5?$/�?s�����o���h��?�g�~S57��h&]�1�e��.���hK�A.f�B�����jl���0�Ä�%�c
2�&�9����V��ۢ&�cB7	n&T�a�l)�0�dHF20�
�#IH1d�4vh 4�Y���ц$)�a34��D��D��00��B\�!��aqқ!����tʹ��lM9���ik���6�^B�КB�I4��d�h`vD��c�@�F�̄���e����,�A)����т���	 ����WW5�V���wp0�a�J��na�,���*B��c`����#[K��K�ݰ��:6D�B,	����7MBa�7����@�����)�H$*~b�`f8Q�㥍�l�4���[B��*B�"� c��7����ߠHU#H�p>p��>o�c�t��N�ϯ|��I�ܷe&M�iE�B�ʼ&�	�ze�[������M���Y����z#HV����G�����A1�ƙ,��aX��܄��(D���e�P�����j���S�6������-��}ۆ�2w�߽�N�}�t��B]�%�ě%B5%¿�ua�
��5�JHF�H�r�J]c�F��Ŗ`K2f$Z�C�oW(�KXl2����bB�0!.�.!	,r�f',ӑ#� WG3Z�)���fD�
@i!
�Cbi��?g�|���,��!P�HGS��{�N�)�dr�T�f9.� �~Hv!J~�}�v�
E�0�\k��B0��
ĂB:I
S������Xa��߈o�	��K�Y��� ���!R4�1!����B���(F�Mf(���M I�2\d�"B!\�6fCLq�����&��� a��²��I�6Lf��Cd���p��'�c9ŁW&�m�4Lj⑪H�a4@�F�Ē
����Ȕ$#_�$!F$)�ѯ�&ha,)����lM�*rS4�a�m"@�'�R:HQ����\%F	p�:4�㓕�Ѡ"T04}�ٴ�Cl9��4���t�!7b�ń��B1�Ʊ4���0��GD,��P�!�F�1��```�
B�	d�3P���
����7�f�Jxc
r������vB);C��@�݌��fͰ�J[޾���vf�Y4��aB$H�"!���[�I��4��s~�~?D�.L���Կ�q�e��)
�"B$�.ٮk�ϸ���M	5�?hvhFbP�8M�\�!.,$5�h!�c��}�>�����~%���~%~HO�d������d%�^N�FB]���wN�,�p�#	�6�g�\����'�\[�ʄ)]
��?)^�t/*����~��v������<Cx�y����&�N`J��]4d7��B~!u�,I�.i���p��
`hH�>��?Gp'XY��>��3wu���Ms��� �x �d)I*�`ĄK�ٛۤ���(K�bB�U�HҚdacm�R�~��D�ć̦��5�����I �A�\��J\R(P�����5��HF!R����F�顾�̄)���j�+��D	��Ǉ�,!�vO�Ě�)	I�H�#����F�����Bt���� �H��c��7Ɏa�!2�!5�"E�q!���2$�-�5��]7���$��4�i5�R�]Rs�s,R"F��M3�]�i�ׄИ�:Nϝ?~���*B���d�v�H����[���ƙ�#R�Y��F����.�%X1��Z���hH]��yL��xp���8��hڇ?]BJc���$%�{#���g���.�� ��!n�&Mc)����5��sI.h��%��h���j��@��c��1cp	L�c�URl���lIϰ��&0�R@�3!P�5����'��Mm�[*RR԰0��a��9�oy0�rf�kfl8����k �S��ת'�~��i��:����޲n~�mz�l)���>8:>�䐆�~g���5�B�@Jf���>%��4����?ǿz��  ���    �^�Vm��RlG!�T«=�	���aN�ne�tU�q8qE,�U@�`Z/V� ��ޠ��8-�vm��g �ڋ��u� -��  h �d�n�a�� �ӫ6��  շ� %H          ��6�/l�� ��[_�>�6݄�l��36 h��[@  o���H�fݛd�     ����	 		     ���m  ��۰     ��ۤ�m� 	�$      �kj@�m�����`m�        [G� ���� -6p[@��m��`  [x� mH 6�m�[@ ���   �� �`���   p���� %��8/Khp� ���l�d���h m�m���`  �p$$ڐm �h   8 ��     6�l    �� �À >rM�� �Ͷ �r�l�햀$�۫`    m�[Amm[;m� �n�����U�jNH � p -��-�-̈́�p  H m��  km��a  ����  ��  h����[\ IbF��h[V� �u�\m[ � ��zI@6� �I,6�cm��m�l!m[A��kv� 6�V�m'@�m�u��-m�Σ��U.�Jp5�K[E\�ʯ2Jjg����h\�6[%<��\����e��^��` �� m�m� m�6�kh�[A:Y���-�       �    ���V�&Ӧ�� 'A�$�h Ą�	 ���mm�8@    6� $  I�   ��t�C� m[A^j��e�vr���^�l�a�� [@�� 6��� ��m �m��L� �9 m&��$-�-�փ����)�ěi1��4����l$)@��cm��l$   6�t��� 		l���c���:�zPqm-�� 6���l�l�8 h�����  ж�� �� 6Z	�  6�\�m�u��֒�k~_��m���� d�sUP�V�K��UU���S��n��tο��7�U` ��tu��Gp ��w�-�6�Y�n��I9 ����TYU^ ���@KԧUA�ɱ.��ɨuK���L�[Ԏ[��ki��v�k�!5,���[`T+GEV쳨VX�W��)X�����b�z��tۢN����� $�d�n@�=Y��UQ-چ	b�g��U�lE���Z� 굚�ih*�ei�ۻ �[NH�6� %�����Zl ���eKz�l�m��|p
t�ne�𥷤���>�u�ݶ�$p�� �'&�2���U@UԨ3�U(Ռ.׫ E�C[��[l�6͜.�Pe�6�`�aoY�9�[\ -�6ݚ̙�]%\ m���V�  ����gizϹ���m��^����uT�R�m� $u$�m�ζJ�Y�l�y�S�I������mW�pUU[K%«Ui�Ul�w-��׮�pm�$ٻ)���� 	ղ�v��^YWj�ge[���5�D�m��F�S�m�UVZ]6 �+��z�$��չ�d���M�G�|�����l��m�U�8А6���yZ�U���,�m�۠ ��F-���-� :�L�U[t��k�*ҕ H['��	�p $t��H^��e�-�@    �%�m����&�  h�tI�l ӎ\�Ѷ��H9\�	�� H���@��lHs����/+*���Wl  9 ���UWP��o�|7ʻRWm��[m�@� 'Ki���%.-� $pۤ�u��۬ײ@  ����w%�.6� 	l ��Z��D�H*�WI��YV��C�-�$�i� �֓m��
�گJ��+oj�.Z
�[{�  �Cm8��n�UJ�U�JJrD�n�6�H�  ���m� x6�j�
j����2=�&�"۵۲� �ܵVz�^h���K(�[;��-�pݵT�� �.�:��B�m�gG`v�-���v���T��6ڀ�V�q��Ȏ����
��SRp �d�@�E�#m�����V�
t�,�WSv�w7e���j�\ĉ$ :�]�D�M,�L   ��[gN�� -�h  �l��ɀ	 �m�m��Hm؛Ip� ����$�^�sB��[q���v����d�t6 �m�&��m� $Yx֔���`�K+� �]��8�p�m��M��I�HNf���t�sm�٬j�7.�]�
����#y��e�8m� �.�6�0     ��s"�	k�l�U�������������ڬv��U����ZE�5r�M^.���^P[cΎ�ܶ��� �Uj��p�g�N-�p"�Tmm��XqvS��I�P��v�6�j�  ����[y# �!r^���sn�kn@p$H ��Y[v�Y���� ^5�C2�)m�.ԫ��6��k-�\l�t�PTŹm��1T�4H[d� @krޒ����)�8�oU�nIWy�kD=�d��1��*@�6��$�M$�֐j�e�v�*�)�\�S�-(*���A��U.x�X�*LU]�K���۷Bڨ8q��H;j��7P�Z�f��p�-W(�Y囎�n�=M��i6�@ �?��v��t� �mt�3L��MSeVQbF��R�,�rגn�:�ph\��W,��*��V�ȧ]m�\���)�![ں�-� �8���v�O�F� WI*M�	ι;SUur�G;9�)�b]�j��*�.�U].�=��*����7���ͷI���%ěj�Sfӎs��f�����yVڪ�)]<��U�l* �� ���m�n��h9	YV��W�SU��������l*Bpj�P%r� h�F�T���Y�-���:	@
��C�ɴUF�U�^���;��c� *���CtQmV�m�	.5�՞��� Y.)V��U�@S�r�]�e��/U*յU*��eB�p�]�V]���[i@豶��۶kX�6�  �ۭ�@�ݶ��dP�j�8iIw<#h���  ������d���lv	3$� �p�`�I6$
<�l�m�� Hm��l{b@%�m���$X�Sh��6 	9:� AWV.԰UUu1E��5�#v�6�mA�WiV�Bk��  ��I�j��s]0 $6�-iWUURD����b�yVNh��   �c�i( ˷m&�8� �Rl��Lֵ���6�n$�a��-�� [B� l���-��^���'� ��`U]A���f�R%�
X *������@\�lg 8H[% MW�w�M�[,��*��Z� ��   �Jۛf�b\��W8c�� $H     h T/  �疶y[��Rr�۶ -�� 8�  m���j���H L��&�v��v�۶�m9$�V���[[m.�vv� -UUUR����[*�r�HU%��m��L����m���ڶ�e�u�zi�E�!�� lHm��   �g9���HYZ.l��������0  H@Usq��٠�<�WR�[h�N�����z��n �b�r���tr���HT����2sUT�4���I8 Xa� �I� �ؔ��RN7a�ej��Z��#�YYL���uR���Ԭ���j���FG��'}�_,�@�gZ`N�+���m������@<�k�n�y�V��[ui1�m��Φ9m-�u�I���$8h�ۀ9!%��klۮ ۥ�.��E�uu��$�$ -6kz�ޡ#��m� ձn��� h ���I]�e9���%�m�U�W�U��ցm����[M�8 �    m�  �ѢH�m [C��t��m����Ln8� ���*��r�9k������w<�[�嶔8 6�p4�-3lj�V5�F���UH�Uz�^V�����[*j���t��R� Uf���mU��m������b^�Qm-�#�� �^�_�����2js<��*ZlVঀ�B�	�� ��mS��h�O6l��!�@�Jk�#m�� �-�eZWX϶�d�vβ��E�eT�0���P�dp�k��[p6�[[l "� @;o- 0�e�n�tP6�k��N4��RmT!��Ė�Y�4ֵ&�j�Hh����
�QU?�Dv~D�a�ES ?�T� ��PvD � k�J����C���A��`F�TN� 6��q_�~z!�:��z| �A:��n?t@�!�4(�>� ����H��G� �
� ��/�E~P��� �D�����*�Ƞ�8�i�H	����H� "�$$&�L^���v�@ ���? ?�((qW��#N�+�h@P����A^��~X
wa��A6���R,"�b��B��EڬO�.�DD�
/�@�*!�O��h!b�P���(��Q� :������0@ $?"`'�QE\Q�e� ��(��������A�ز\^���s��'m=�(�.ٺA����L��{Y��/K�9��IpZ��+.�J�K"�UV�V*�Z[��7I�:��i<����DjU��m���m��\���o^ �j�Q�g�6�MJ�U���m����Ĥ% �e�vP�^-��I�%T;�Ftlv��꣗��<T`+`٣5. P�Q�\��UK�S�r�kDaz(,�Ŵ`O-����ў��L�5n�9A�ٖ�FkZ�Q�h/m�t/N[m�wh *e�]%V���AAn*��;�W���]<.ۛ�����צ�e�q�v2�W[;��$l�A�Z��8i�`�l���j�ɂ���Y^;
6C2@���X-���'O%
f�Q�,�N�y�j�������[-3i���gg��T��LR�n7l����Z���Vǵ�v{
�k"[��&�/����&+���;\�C�2:<��Ѫ�v�r��AV��K �<aʜF�t-h�b3h�)��pM�X�V{�r���p�[���RX�6LD���v`;{9w8&/UUPbT6{\]J\�
��\mcA۳W6����g.$P-�6 70W]*!s���c@�]��p��6y������om�V\SJ�/�BZ{$@*c��I�����n��ٞM���6`ݹ�E� �րW[�"C&� 4���v	��n4M�ga����m�\�]�ݍrc��Ì�-���mX�c���1�s�nˊ�R�XL*����*w#"J���99�3�4D̔8����A�V��s�@vWIvX6�E�A�!�m�sL���3�z���jH�/`k��-�]$����4ks���-Ԛ:7q���ݪ��:�;a�re�ÒY-m�k�HI�II6[���h�l�By�ʣf�q)v�M��5��4�36�ĶD(F��!컬�nz�qe�:T��X ��؄��T��ڱET�Ȍ�TB���O�M  ((b�� ��Irp��98O�Sm;\ʺ#r�-b�5u�-� L@
5I.�k�ǇxY��2q���,9� �T���.SQō9狯n������1�9��_;i۱ծ�țM`��umcY�լ�[��c�]sK�m��I(ᭅ�xnmT�Xj݉��qM�ڪ\���9���{XR�F5�
j�x��pa�Egf4�;���S33Z%�&�֋�*���1M����	��S<;�
��|<�*G*��ˇ��=��I���R�MvU��2�F�?k�_������_�l��0��i��;���Bj��ty�U$ts�l��0�&V�5Ҁ�����V��;x���.�+ �gG�t���h�n���`�\0�&V��G�o>� +�J@�V2��+.��?I2���<��X�u8K��3mu�֭����\0R]�Q.��r���F}��&ff;a�5nV�ߞgG�w>� ���~�e`��,�\��Y5�Y���>�>��Ӫ����H���
����zW�W����wL�y���L�.�eU�o@���à|��;:�<��Xu>��]�����Wf�I��z�:?�� �ϖ�.�i��7t����xs��p�?I2���c-v�^0r��e���1�%�s�ĬZ�Z!��YIc��uՀM��,j����o�^���X�+ �r7�Mb��E�t���`�E�~�2��#x�����@�Uc�~��?I2�$��w���q��~������]�5�X�8�P'@��I&ۺ�7����E�vˆ�L����ך�-��o �r,�\0�e`�F��J��,wce�N��;2����qz�Ƽ�4����	J�q�c������m�wwv�v��p�6I��o9�;�� ���Qc�cWf�L�y����Xl�`:A�Rt����b�`�F��"�;e� �&V�5Ҁ��컥V��v���Xl�`$��+��z��DBE� �B�3�����>�_J<6�mһ��;e� �&V��Xs�`V�|R��mZ�n��S:m`�(	��� ˸�n�{��[̄9�2��-�&s����?���:��E�w9�.Ӝv��J줓m�`�G�w9Ӯ�2�ӣ�*ך����ݼ�Ȱ�p�6I��r���L�E�i��wh��k ��d�`�G�w9Ҝ��5j�+Z�0�e`Ȃw=�g$��{�rO���7$�| ��~c��������A���?|���,e�*͚[�5J؀��x4G�:�]�	Bk���f�Λ���'c�a9�������PSѰ��ngH�ۭ�a��f�Ro�!��+R3-b��YX�&k�� Z8J�&ʑ�4�[�^!HKs���B�#g�v��Ey�ܘP�mMZ{d,�AK���tm����Q�z��m*v������V�V�)k�\ɍR��;3����j�s�ڬ�X�Wi�.�ek�H�j�qX����]<"˪��<���C������;�� ��d�X��J���t���ݼ�Ȱ�p�6I��r�5�J<6�mһ��:t��6I��r���X�[�	5V[�T6]�`$��9N� �r,�L� �;T
��WI6���txs�`:e`$��.���� �����F!��\��K���F�a8[�n����G]p+z9�S���]��Ȱ�2��e`�E�>xy�c��Z@sz��>9��Lv|m`��LrO�Ȱ�"�7��D��TX��0���e`�E�w9�&V C�b7v]պC���{�]/�#��oI��l�+ 향���v��V����w9�t�>?�}�V��X�<�xF���X,S6�7��kk�Z��g���@lfqJf��v�u��
�wk ޗd�X�`�E�E[�	5VZv!���d�Y����ꤎ��#��oK� t]�t
쫤�n� �r,�Ȱ=]���{�To�ԯ�^N�X�#y橤�m[
v��"�7�E�l�+ ޻N$��y�����ģ�_u�,d�X�r,�Ȱ��2�/&���OW9�S�L�R��֥:�6�N9�:|��7������	�L[�>��X�r,��X�� �黲���`�Ȱ��`Ϣ�>y睝����Z~�_=�6�����ށ#�,y�X�&V�H�	�RQ�ˠ�]��`� �&V�w��4��(DiACW{�w�rNU:����n���l�+ �$xs�`� ��Ѭ-�j�VӧuhC�-�=�l�\6Ɏh�g��]1Һ��me�+���+͌�m��/�����E�tr,d�X�Fg����l<����E���UURD�ϖ�}�V��X�I�t]��m��(-��7�E�l�+ ��E�w9�>��;j���L-ݬd�X�r,�Ȱ�"�t�CT�;����`�E�}QϾ���� �&V �T���?���@�
;q�P��q��c n9m��L鲁��%���f��D��AA��;q�?�j���VI��y����u���HY:Ԙc�,�Ȥv�5�1B���Y�+b��+8�ݷ��v�"\���9��Gl�X��,��a6讂��J�.I�Z�L�Z�Z��
��!��xn#��5�{=��s��$��a�[ŖjL-��h�]]B�yWJ��GN�%tU,�rXb����h̎�a`��L[��0O['D˺��sӶ�5��.����x�`$��7�� ��%���I]�v��"�6I��r�ˤx�[)�!;^��T�ݬd�X)#�9t� ��X��mR�[�WI6���H�]#�:9�L�{���Tē����ݼ�H��{��T���~������g���$[v�4����A�YyV9�0)vz�%�,H�������.�+�̢�wh�ӷ�tr,d�X)#�9t� �r�@�V]��wk �&VeA "�IH) X�=T��^���$xS��:9 C�:N컥b�`�� ��<��`$��65ҀmwmQWv]��9t� �}�L��96���[�ZB�j��Ϣ�6I��~�"�9t� ���U[+�'v��V�������#�d��+�.�������k]��jͦd�7�d�cf������>~r,�H���`t�ڤ+���[m�`�ȳ�H�}��:9��6I��or��kΒnՠ�Wk ��<$��w�s�I�GJ�@����$�U��` ����R���߳4� �h��"�D&��H֣H� ( �lv�R� �ES �lC��DK�'E��!��������7$�޻�s���`�6�ݻ�Qi������s�w�}��r�<��9�� ���_$;MӶ���[�XΙXި�������Ⱥ��䜿{�=m���6���)���UŒ�$�F��k�����r�d��g������t�E�ց����x-����~A�}�V�5>�E��TU�6���G�RD�ϖ�}�V�ty���?���a�Ѵ��������>�睝���$�v�Ė���s��m9�L����]#���+�=���$���9;��/@'�</�Vu�.�]`�Ȱ�r,yȰ3h���Xr�
f0N�J4k�)]C��u��C��Js�ϭ��n*凯'��۶.��H��2��e`�E�~��)�m;����i��7���6I��o9ˤxp�
�m�v���Wu�w�}������9t� ޓ+ !�4�����V!���tx.��:e`$��?F�P���Wtӷ�r���V�L������{֨�L�Ĉ��Di$���ñz�Z�@
��9�V6��`F���+m�$��P����]\\���j��0[u>:�@��N��	��G&�͈�Cb��%A�(����G8vA�[[7�;R7��,f!)�����8�5��^=��SX��m�`9Ë��I��9ۗ���G��I<N�n�XK��l��C��"R�%ab�j���'$��{�R麻A}$��Bi�ՐR�4*&���&�YX��dC�tה�茱l��� �}2��e`Ϣ�9t� ��S�IUڦݥM���2�[#�9l� ��+ +�(�B�l�bm;����[#�6t��6t��?w)Y��&�Z'v�[#�6t��6t��7�E�mt�Hv�N��?]��I��l镀o>� �< ���Q��n�YshU��t��q�.���aA$�)�m�u9嘧��鱳̓����V�dx-��z���}��X�>���:N�v+wu�r��dx�2��2��t���v����i��9l� �.}�?Q����V��~�V��E�˫HM]��6K���Vˤx-���td�*�T���1;0�2�]#�9l� �<|:��f�{5nj�.xIV˵��#�n(����sN�Wh᪍zOY��b�cUlM�u���<�����l�+ ���}_�ם$ݫA����"�|���N�+ �Ϣ�?T��4�wv�����N�+����N�ު�UT��Ȱ�G�~�}E�j��n�U�ـN�+ �Ϣ�"�	o{(p *���H8��rf��r���33�g���� v���{n��/n9$��'�8I"4�c�]2�\�q��t8�K	��gx�LWn�ӍO�$�8� �׺�d��������G ���bKR@���G��d��������G 
�k� �:�#$1������{n���r��}��}�(p 3��kO�'0s7@>� +�t��C�}�s�st �K���ip�X��8 W�^��r����uʎ uaZ)�.,<�Aٳ��'F���V�s�[�W��F;
��\A�!�I�5�U����|�߿�Q�������G 
�k� �uʄ��2<H��G �w7@>� +�t�Qζ��򴁣	#p"�ɛ�uʎ �׺�\��{n��Yۋm�$Xc������@;\��{۹��s� ���,Q9�$�t��a�������� �����{߷�&���`�[��®�0�gC���)M��VՍ�y �5S�gxƄƫc���c޷�˴�v�wc;�v��-1�}�Z�=�:�;3Ƙ�]��v�F����ȯX��s���g;���v�r�]v��a���5d�·�^��i��㕗�l�Ec;Ǝ�-���c%�fR�5�w�=���D�ݔA��Ke#���j�r�%0�5�����I9��I6�/zM�h��(Zf�dR�mk����jٳ�̞?����/2�rQ��8X�;f�h��������> �׺��0� u^����F�`6�n�tv��}��v�C���z\���H���9����@;]� /m�� �� �n�x������t��b�{n��Gh� W�^���F)x�fLO �. ��n�tv��}��v��\ �-hq����<&I �*��7!Nf����F+6�gn���tv�B�N�ё�H&�rf�k� +�t��p ��st���X�r2E�����v�{�w��Pp��(��ö�b�~�st�ʎ �!jKNEH��m��������31�|烀�����w������%������(p �����x. U�Љ�D�hCnf�l�8 W�^�l� �w7@:����I1C7���e��=u�
�ոG�<Mׇ��
:�dXݜ��`�G p ����� _Op\ /m�� 풇 �j��<ljc��G� �w�s߿f~�m�}�nn�_9�p ��t�r�H4ڂ��70���st�ʎ�f~�߱}��v��8 W��FF� ��7@;\����^�k�À�����R�ۑ��o"�#�_m{��� [w7@>���^Qb��!T0��`�Q�ZM,c�lXEX�4�Za���CA:5]�h���%?� ��� [w7@>�������
c���Ħ4�À��v�b�_m{�u�a� �ޗ?(�im�� ��s 
�k� ��� ��t �/�&�5%�G1p ������0�{-�嶠�<*a	�DkF�k��Y*(XE��9�|޿a�m����>s:b�囅�{�u�a��}y�|OO'����@>�%�d1�����	�'�9�Ocaγ�(�o=SN�����;	�hpP���p�*~&F�G0�{-7@>�À}��}�y� 
���h���X����0�a�}����8 ^�M�f6���$N~��G0��}��]�f6�g�n�_9�p ��RYrA��FH�@��}�n. ��7@;\����ߥ���L~~� Hco�ԓ �i���}9�h�}��g1p �f/ߖaD��!��'߇��0 ��X�"HH�#^Ն�Z3@P��QC~F�(TaB�JƬ �H�
����!	[�� �@F1\d�Ŋ�$B 	 � �"(@"H#!��F!��䁭�a �B�H��VB0�% ������aFF$�R�DF���[%H�%��T#A�Q��-�Q�`@�'MK�wd�h���@�@���)!JA�J�)�R��J�A([%eb~�LB���"�hJ�KB�"D�P�a4� `W��!��"��;u��(J4Ҧ���?\y����0��R� �"hD�`BD�q���1!B�6RS*��"�P�E%"��*BR�XFcu�2��+"���q��8��o���R�U8
�U��=^*ur���[f�f�ʐf�T� :i���ny�U��]���J���UV쬺*�6%Q���#'m���%�����;1���.����'��*�dBWS�h�@4Q�J�8���Z��Tc��'[V&� ��.u�$]6%9��0#*��,�vr�r��6�W gg�������n8�JP�`���2��R��	�	�$c/&��$1n�[U걼l��$g��욹ݝ�p��*ƸB\`�e��׷1(� ����n\x�-��$מ�ǰ�Q'cBL6۲���ϟ�h�my�ת�o-�4\�nD�X�	��ه�pv4k�@����l�حU���]�y��9Kb��Ҫkuv��*�C6�"U0�hj����dڣmS���B*�x秏n8y���O<n+n1��0���0��#�K��ۭ��wd���Q�ۚ�����kkr����qtJnIk�`����9�&69%6�P�v�tBA��ቁ
b�����;l�\�C�@kP�N�`���Ԫ��ڶ�bȮ�e[9�ܗ[]���� r�uj{E��R��.��Q�D�g3"�6)��Qim����ї�[˻�i=ld�`�ɱy˺7 �#��s���,b`�ୖ�q�7Iv��^9Xd9	n�:��f���8�i��)Y��-F�j3р�v }�#`�R'/��{]�x�j�N�@:�ʳ��u�	8WmQ���� Q�nԙ�v�L�\�N�!�<� @�k+���@Ӹ����<���@8��]���3��q\�<v��tI�a��B���ܭUV>~���wl��>��zr��I4f���sa\�ZI�v�@�;/�s�>~�b�#�꡴.ծI��M0ƴ�Lb9�n�N��+��s��N�r�d��	ӓ�h{(�������l�cn�� ���M+�s+Nm�lW[����!�TchԪ]\��]�A�k�N������
���7U̝=����ɘ]ff�CZ��|]�!�I#�NN�I���Q[*��YM���q���i�;cv�Y4�2�L�c��d�����u�h�^8���P�5e�*d�PA���(6��EƴO�zy�r�a�j�x�#��:k��MCum�N��t)Hm�"��������Ô�ְ�*�p$+ �jͬ16���fy�趼���UVä��7T��&�8�[����k���;]�kG)�www��p��'�nI�j�y�la0]�vu�`$ڋD~^憲�ڳ!���98L��?"D������?��_m{��s��k`z�x� =�܋�be�A�wbĒQ�����U��]����� ?������G 7-�����rc���:I��N}�_����_�)����+���i��v7V��Ծ�>XO���"�˧�~��S視1նX]�7v��p�>��}���}��W���InS:T��$�'� �8�k�ً�ˠ�강�M�z����<lv�H깑��m]��iՖ��"�ӦV9�XN�`��԰*�5v:)�wo �������E�t�����I���HI+�˿]+.��>�|��p�"�Ӯ	ī�»$��XN�`l� ��s�����&ն��ݘ[#�:u� ��,�\0կ��7m�۴&���g��=��sun\Tm�Z�<C.���d�D�t��;t�v���J��:�N}�m�q%O�|Ioz+$lja"x��s��2��G�oK�}���I*�}C��Jڰ��n�`>�+ �dxuo�UU�o�^��`��
�Wc�ZulWu�r��.��`u)�u5%�M]�v���;_�{� ��-����`�I�/�^���/O]%
���E� Xt�X�D^[�W\�[j�*G'@�E�t��dxN�`T�U�W�;󤛷k ޓ+ �<z\0���"��P��&�W�u�r��.��`�e`�(g��i���~�x��`E�oI��#��@� �w��'�黎j��c�T��ـl}�&V�dx��`펊��-���M%N豵6"�d"���A�岫��-d�{Hm�nX�r�Aؐ1Ҷ�.��v��2�[#�7�� ��, ��%V�����lWu�r�}U��GO�� ��`�e`����P���j����l}�&V�dx��Ē�L��Ҳ��c��2�[#�7�� ���B��nݬzL�����p�6>� ������+R�v㍋�\YC���S�u*UrZHfS)Ơ���]��A�ƪp��k����a��6sµ��z.�q����M�ee��#�`����d��<�c#�g=B�ۦG��[S��M�K��b0���(9s7ٶ)M��#�1�C�G;a�ةy�	�Wv�l�j��i���\w�.G�y��s%��K=�R6V�f�I4�Ը�6դ���W%�7\��u�5(Pr��̥&��bhJ��WvP��-��n�@�N����O�ϻ�	�O��lܓ�'}v�`ӻ���]�z\3��W�;�>X_{�ėO�|Inw�e���H,2��`�e`�G�oK�t�4t��o�wk ޓ+ �<z\0����HRUi]��m��wX-����l}�&V N����'�h��eޝ��M��q�0�������7�F�%:zn��H56�.��`�e`�G�Mq8�Wj���L�f��XW��PoI��r��.��ު��|�����������k ���X-����l} BIe.���u����>��c�>��]>��`J'�<��V��U�j����l}�&N������>_���M�5��S0f���s�J��q�"����6ݵ�ue�7nt%�8z�;m;N��J�]���`�e`�G�oK�t�:T�J���v��2�[#�7���6>� �K�Ui;�~��j�[#�7���=U^���>� ��+ �:�.��w@j���&V��X��XU{�T��x��_[^]��w@����6>� �+ �<d�X�r�tզU���h�@����N��Yx���.5�;Nwm��]\Ė�6R���߼�r��&V��X	%� �T[�U�u�r��L�c��2��H�Q>Y�n����W᫷�O��X��`:e`�G�mJ�R۶�����Ӻ�6>� ��+ �<"  ��~�E����;O��Zc�e���]��L�����2t�o�^��''99>�|�eT�9�q�*�`b�!rF���2^)��+CP٭\Ej��ۜ<nY�/�}�����`E�t镀~�b�G�N�Ӣ��ݼ�L�c��2�[#ϫԑ����ׅWj��_�.��ϖӦVz�(��>�e`���cw`!�v��2�[#�:t��6>� *IB�V��ꭻ� ���2����:t��=�^*�{{���j�r7(c8-��l�������܅q��L�$��l��ȏ�{s�q۫�'u��(�i���äm�j�S�v�˘��L;�s��}8ܻD�5W�C���͝xA��	��90؅��E�m���t��2�7	�A�:�m����'��<���'f��;f;C�1ľ]j�t�\Dw)�rB0�v*�ٔ�T�gI8u�s��s�ۂ�4�$�X\[�����ѣ����6K�^�r[�{8H��Z4�6�+���kU����g@�����:e`l��mJ�R۶'i��)SN� ��,�L�ꪯ�"�x�}����������Lv��2�[#�:t��6>� �K�Ui;c�&X�� �<�L�c��2�	�RQ���v�ջj��:e`E�t镀r��������)�M���jB���\V��1nc�Q��ɴ��I��z�v�d!����b٪<�V}�����:t��9l� ��+ 8��(+1��Sg7�~����d�!9	$����s��ӦV��XRH�ZN�uV�� v�xN�X��`:e`����;wv�~i]�ӦV��XN�X�%�R�Էv�v�wE*i�`E�t镀�^���q$�\����G�xLrF�eanf��fVK4��N[^������Z�1\�:�V�Lv��2��K�:t����W��|�� ��_]!U��5~c�� ���2����:t��'1IG�.�V�� ��+ ��,>��*>$� �_�$c3II I�c08M��4�,�T��֨X��?&5B�F ��@�|���d! �d�#Lt@�)P�"�v�"(Z��!%4J��C0�$��8�lÑI�r"�A�I#�TR���H"!�x��E0Q�> � �?
C�M��_�s�7$�{��rO�vj�G��j�;)��� ��,��V v�x�&V q9��WLm��۵�wt���/ �$��6>� ��b� ���rX[�˒�h���5�k��^�	�{/@
1��n�ѡn.���/ �$��6>� �镀N���+t���e��wx��+ ��,��V v�xT�����N�n�M;�c�ޙX}꤉�}x�>��	�����Һt�Wk �镀�^�t��6>� �K�%m;M_��v��K�?N�X��`�2���[��a�0ԚͣL����h�,"��,�ĳj���l9��]���J쒻��镀l}��+ ;d�z��J��;n�.����;ze`l��~�2���O�cL�!�v�ޙX�%���X��`v� �[n��RWu�����׀o�}��l}��+ �GE�J�n��/�+��?I2����;�e`l��?Ut��H*Pl��#�k�K��rsrr�/����5ܢ�x�V/��1��po��ml��j�(�&�m�:�&��� �g���Kq�:۱�f��K�.)�)9g���B(�X1���@���Ѷ���(8�͡��nլ<EF���j^������E�'.Jd`��sk��&�{��c�Δ�q6y$�<��c\� cs!��������� K�z��8R���Y���%^�5��X���I�7Iנ$�m�u��WT�6b���)2DˇJL�v'uE�M�"u�S]�M�V����J�wX���`�2��K�?I2�tr�I��Ҷv��X�%��L�c�]�VӴ��*�n� ;d��I��l}��<s�y�t�[������L�c�]��l��oBԳ�S�[���wX��`����/ ��e`��];۴2���כv�N�s�\%����;Y��=OK: ��Rb���rW�WLJ��Cv�~��< ���&V��X_�DP��mݎ�v��K�_�ꫪ���~����|�]�����U��j�һ���+ ��,�tx�%�R��wm��m�wX�N�X����vwvV ws�&:�J�2�v�]���/ �$��'>� ��Wʢ��v]����7��_f��7n�W;kQH�Y��k6X�-��b���w�{��?I2�	Ϣ�9wG�w1IG��+�cWw�~�2�	Ϣ�7_E�E�<��C�S�*�l��`�E�~��v�""n��(�([#�:I���9��"��Bv�`��X[#�?l�X��`t����[�i�RN�-����V9�X��
��때�wwv�ӻ(ٶg�G�����`��hX �	��cI��9��'���$&H��߻y�I^�Հ~޸`l� ���M�bw`��u�N}��+ &�{��ﲰO������WC(Wk �镀d���+ ��,�E.�+n���B���`�/ �$��'>�k�U�*�UG��t��;���v	+�Zv���&V#��X'K�?~�妷f�if"�  ][��o(�9��%(A`�B�ؖ3�b�^�����c�u[wX���7�e`�/ ��e`Wp�W���k �&V I���2�	E�;����1������ ����E�H�,d�Xutu�J��e�ջ��Ȱ	E�l镀t��J�*��mU�l&�	E�l镀t���V �����CH�����L׵�
;9ȉ�v��\лE��q��M�YMSY�[�#�p�<��`�n��=X����r�QK�gkBg�'��Ӧ���+��藚CGn�uv̀�k���\ڵ����! ;h1�]q�T�<@��D.pSkn�\�D�����D
̰	f�񣃱�JtlÛoF��N��أV�U�W.y��e�!��C1umMm[(��vNNu�Н@t�\l�v&x3B,5�b撕c4�\W�CL�F�5�&�m��.4�kB��y｝ �t���V#��r�Bn���2�� $�y��$I��X�9��6I��w1t5w@���v���2�	E�l�+ $�x�5!䩗V�Z.�wX���6t��	:^�&Vwy
�&��M۵�l镀:^�&V��X:�Iv&!�n���H�9���<�k1�]��)�)$$���u��	U��yo]L�����?x��2����6t��'TP�b�M�]�M[��;d������*���G�`:e`N��mJ�*��mZwv����Ȱ�2����vɕ�l�Sŉ���`7f;�V t��	�e`%� �9K�	�M�V���� t����}����	���M镀}�������n�k�cumؔ}�rWیY%�9�}Q���1��K��v�a��>��;wx�2��E�N�+ :Ix�ԇ��][�h���XG�`$��9N� ��wy
�w��f���{�rO�~�nhDG�@C$����|��r�H.���Qn� :t���G�`}UU�O�V���[�ӻV�w�v�� ��,�镀:^��.���Z��Ӡ���M���%vē�9�I�6C&f�8��ti�b7T�9�vi�أ����O�y��ۀl镀:^�.�#�(E��m��XΙY���}>�w��t}�r�Bm�ʴc�� ����p������ϖ�O��ӪӁ�O�ګ���>���;���'�|���~���C� �	 ��1�����rOݙ{��d֦Vj���:>� ��U��~�����eày�O�C�g4�X��,ͻ[r���I�%4��Y�F����N�LNo�l�ci�v�	�2��K�&ˇު�~A>s���}�餝���`N��Uz�T��}�ϖ;�V:�:�E�M;.�RV��	��t}z��R]��+ '���6�N�[J��ݵAwf��U�>���;��V t�xO�E��o�rI��g�K5f�3.L%�XΙXӥ���t} W� )�q�1#$H�!aA'�� ��d�yVh �B�8U ��Iv\���%�ere��!�,�0�#$����2$��h��@�C`D� A D�a)%mSLp20��a@�X$�L@��c	A��6$V F(Dph�QhO���V̬��l�� HB7�s%0!C$ �	N�<ꭵU%v1��c3;i�L[�����7t�qa��tD�WUR�%�
E�6�[mC�n��ZL� [P[v�6�m�&�Yimv˺�D�#z�s���3U$��U83)��]l��PQ-YG��U�eJ�%�);UUt��P�e@�56]�1*�vZ�si���R� ;ci],WF�lԄv���	���d6�Y��K+UGY#i�EZ L�l��\F��se�@ưtp��U�����.�P�:ɠр��)�s�T|U8�Ɓ��e�[���hbu�5ػWGm�nIw�<vrÞ�D�Kc�>*�����4k�jMv������(2�n��#���.zˈ��f� Ѓg�6ݢ*���\��v�v�W��]6��<�.^��!5l�6����ݧ���]� ��$b�� �aU�N��kr�[JnλX��X�N�g�D���i���g�݊�7��>�Ҕu5P��E�<�a%��`#1��C$j��;Z0e��� �#`��P�xy�����C�m�煱��[2�UGn0��(��\m�f�m�(f�)f|s��y�n���we��v��鈮58Ek�e�(���[����r�@=�� f��n�9ۅ;X]���N���]��)����tW/�Zݐ}�"�6�q[�n=a����u�����\�0��!�5wgsR/e{=gm�"l9=nnS�{UFځX�U�fT�P"TY�r5уB�E��=�ʼ�tu���T]CbI�Y wLv�8�4���F抻�#�6�;�U�-8uҎP�îW��on�NB1P�����^���`)���Y�V]�;s'oU�eу��A���;��N0� 8���jy�4)c��a���v��"�]sņ�]�fM-�X𡣂�vp�ٟU����a��'E�P�M���u�[n�󝚪�ӆ�\`0W7<���Wq�Χ�a��v�Bk%��y�l�aW:ܗj�i9s�2�VW�j�\:��-��h�ֶ��Y猒^I�v�1^��1M�~���{
S��坶x��õ�b�[)%D�r�휝��u�1d���]�)n#TLk��{t�i4�L��Nzy�`X�Yz�p�Jm�aƇ{m�82��`;2ͣp`�V�H.���cV��α��u��!6��wL�{x�����Y�����P=��HU����"8Ѷ� ��u*֕ݹ,b��CŁ�IHX�V<n�D"0�6s3�N���ʭ�t8E���oFz���,bCBf%m�P��A��ʞ��9��	n�d������}xl�`E�W�U�~A�O���U��zӤ[,����.G�`�e`N��z��ԑ�k�L�;I]�ـO��`�e`N��M�*���e[m�v�>��y}'߫ '���&ˆޯR�\�`t���AtГ��-�`N��M���	�2�	$���N�i\K�R69���*+m��U�GX]ɴ�D����y�q�t쥅p�7-r��޾��};�V t�x�I��ڻwzդ��M�>�}ۿ�@��`�W�!�>���}xl�`�)<���N��B�XΙXӥ������`�>X��]�M;*��Z����/ ���>]���a�ԏR=>���އ�DJ��O�%9)�NN���m9ı,N�]��r%�bX�{���Kı/}�kiȖ%�b{��|��#muC4�.v�
�e��:H��fx��J�	��A%XCA�X�H[ss�*�56��bX�'}���9ı,O��p�r%�bX��ﵰ�'�ı=���M�"X�%����3���kP�̹���r%�bX�}�p�r�r&D�/�����"X�%������9ı,N�]��r%�bX���<�5f�Y+f�Fӑ,KĽ�}��"X�%���]�"X�*�R+Qb�b(`8dL��k��ND�,K�w�6��bX�'�w�q��Fj�F6�MkiȖ%�b{�{�iȖ%�bw��ӑ,K��{�ND�,K��OkiȖ%�b}�{~���U� +{���%9)�篞��|�bX�'��p�r%�bX��z{[ND�,K�w~�ND�,K���d�"m1��\���\f���S������sv�F�f�&�����<s7n\7(�G�Ȗ%�b{���ӑ,KĽ����r%�bX�����r%�bX�����O�%9)�NO��OXK[�I��U�ND�,K��OkiȖ%�b{���iȖ%�bw��ӑ,K�����" �eL�b}��w?�uq�ɨd���m9ı,O���iȖ%�bw��ӑ,�!�2'�}��iȖ%�b_w�kiȖ%�b|wSބ�段���MkSiȖ%�bw��ӑ,K�����ӑ,KĽ����r%�`hU?��TZ�D? lS|��}���Kı?����6]HM����f�ӑ,K�����ӑ,KĽ����r%�bX�����r%�bX�����Kı?� ������Y��mWh���ўY�&y��F�*1�Հ7V�tXy;^���r��c�F��R�\Ϝ�NKı/��?���Kı;�w��Kı;�w�iȖ%�b~�}�iȖ%�b{�}�Ktf�5q��k[ND�,K�w~�NC�Q�L�b{�^��ND��2&D����6��bX�2��������NJrS�����ֱڵZ�Iu���Kı;�w�iȖ%�b~�}�iȖ!bX��z{[ND�,K�w~�ND�,K�{���34e�).�v��bX�'�w�6��bX�%�ޞ�ӑ,K���ߦӑ,K�;�w�iȖ%�b~�^����u�CX段�iȖ%�b^���m9ı,N���m9ı,N�]��r%�bX���p�r%�bX�_� �w��~:V�&���ѽ���Dd ���m �6�r�3�W+�	�6�0�f����wH�9�RXa&�����ݣ�TA�Q�lk�s��9�d��#������l0��΅;o`i,c��c0��Ֆ;R9�Ͷ�彍u��#*#m�9}uI��/6�)���q�d6�.���!��ks�6շ1%9.FCR�b8�9�fsB��'�sY�K��3[)>�l[Szv�=1�^2ʤԆx\�E֥L�cs7D�$�Ƚ��rX�%�߻�m9ı,N�]��r%�bX���p�'"X�%�{�����e9)�NO�������ʣ��|9,K���]�!�(�"dK�����Kı/��?���Kı=�}ͧ"��bX�ý��RFK�˚�]�"X�%���ND�,K��OkiȖ4X�'�ﴛ�H�}��ڒ	"s�m��rJٙ��A�/~�����bX�'�ﹴ�Kı;�w�iȖ%�b{���ӑ,K��N�6���fk2�MkiȖ%�b{���ND�,KW���6��bX�'��m9ı,K߽=��"X�rS����j|m��ֳPeK#f+	�P��#�gc�A3�U<\m��/���])3�\�ӑ,K�﻿M�"X�%���ND�,K��Oka�"�PW�L�bX�����ӑ,KĽ?�������.ZMf�ӑ,K�����!Qc"X�%�ޞ�ӑ,K�����ӑ,K�﻿M�"�%�NOߟOXJ몤w3U���rS���%�ޞ�ӑ,K�����ӑ,K�﻿M�"X�%����ND�,Jr}��۽�7G[��^�|9)�Np ,N��z�9ı,N����r%�bX�{���Kı/~�����NJrS���=�nkb�M��O�%ı;���iȖ%�`��m9ı,K߽=��"X�%�ߵ�]���NJrS�����ͷm��3�l��DF��ƍn�kԲ���1,tn��CD�WF�3%��kT����%9)������"X�%�{�����Kı;���yı,N����Kı)�|y�j�Ժ�4Y�iȖ%�b^���m9ı,N��z�9ı,N����Kı>�}�iȟ�2s�c������_���WbkQv��bX�'�����Kı;�o�iȖ0�%2&D����"X�%�}��kiȖ%�b}�{g�tk2��5a&����K�A�;�o�iȖ%�b}���ӑ,KĽ淋��Kı;����Kı/ǽ��Z��əi356��bX�'��m9ı,Qo{��m9ı,N��z�9ı,N����r%�bX���z����^C���/g��V�A�R�v�՘��7�m���e�+Wn$Jc��}��o%�b^����r%�bX��^��r%�bX�����,K�������NJrS���t���䘹���bX�'~׽v����D+���b{���ӑ,K�����m9ı,K��{[N@Kı>=��F�5uLԚ����r%�bX�����Kı>�}�iȖ%�b^����r%�bX��^��r%�bX�ӽ��RCZ˩&k5���K��w�6��bX�%�}=��"X�%�ߵ�]�"X�V���;�o�iȖ%�bS���n����h��Ѵ�Kı/{��m9ı,�k޻ND�,K���6��bX�'��m9ı,��7���˶sU��d4�G;�����*1-�5�s���2uӭ�z3һ��^N��S��u5��"X�%�ߵ�]�"X�%��{~�ND�,K�w�6!Ȗ%�b^����r%�bX�x���]jff�3Z��kZ�ND�,K�׽v��bX�'��m9ı,K��{[ND�,K�{~�ND�@�"X�����&CR]jf\��5v��bX�'���iȖ%�b^����r%�bX�����r%�bX�����Kı>�^=a-�����w���NJNINK��{[ND�,K�{~�ND�,K�׽v��bX��̉��~6��c)�NO<������rJU��Jp�,N���m9ı,?������v��X�%���p�r%�bX�������bX�'��`����[��Yu�f���g���@li�^7d# \��"�ܻ�\��#�=��l�� �sn^T��ֻQ9�@�ʛ��ǌ�õ�LÝ��p8���kC�xc��d�kn9B�Զ�yI�Ӹ6dG[[a�����n|e
� r���ý��C�̒�WZK�lQ
��p��)@�
헫��:��f��k&�.g�X��
��D5���{r:�j�&�0�`6�n��g���/��x]�2�\O�oj�\Z���WT�I����r%�bX�k���9ı,O��p�r%�bX�����Ȗ%�bw�o�iȖ%�b_N�g��Iˢf��]�"X�%����NC� H�L�b_{�kiȖ%�b{����ND�,K�׽v��6%�bS�zy�D��u��.�Fӑ,KĽ淋��Kı;����Kı;�{�iȖ%�b{���"X�%���{���`�*�Mj/y>��%8{�o�iȖ%�bw���ӑ,K��{�ND�,Ľ淋��Kħ'�!�g�̻;e-���'Ò���;�{�iȖ%�b{���"X�%�{�OkiȖ%�b{�o�iȖ%��%��g��f�7P��]�Ee���ݳ��V1�c��	�Z�F�$%^�)]k.L��5v��bX�'��p�r%�bX�������bX�'���6��bX�'}��m9ı,O�ק�K-�f���Xk5�iȖ%�b^����rSqE 0EDș���ߦӑ,K���{�iȖ%�b{���""�L�bw�۷?�5�ԙ2�Yu��m9ı,O��o�m9ı,N�^��r%���b}���ӑ,KĽ淋��Kı?|{sڍ�j�Z�.�jm9ı,N�^��r%�bX��}�iȖ%�b^����r%�`"+����M�"X�%���7����pe[�O�%9)�NO|�ߓiȖ%�a��,s�����~�bX�'���6��bX�'}�z�9ı)�}�Y�\.Èr�
a��oX�W�nH�VQ�����ġk��s�v/N��6�Fi�Y�iȖ%�b^����r%�bX�����r%�bX�����Kı=���ӑ,K�������L�kS�SZ�r%�bX�����r-�bX�����Kı=���ӑ,KĽ淋��Kı>���˳r��
���rS�������oy>D�,K��m9Ƌ�|1��"��?PS��U"��8���AY1i���T!���A�=�M&B�g *@ ?#["15�	��-�@�@���h9�v� *P��/� "� �*@�
�"��P���Q.w�����bX�'~��6��bX�'ǽ�FXjK�e3-&f�ӑ,KP�=���ӑ,KĽ淋��Kı=����Kı;�o�iȖ%�b}��=�Yn�4\u��h�r%�bX�������bX��Q�����O�,K������ӑ,K��{�ND�,K��zn5h+d#rgԕ�6!��=aqn&7�OY|m�Ӌ�^d����H�q5��"X�%�ｿM�"X�%��{~�ND�,K��lT�,KĽ淋��Kı?|wsڍ�j�Y�K���ND�,K�׽v��bX�'��p�r%�bX�������bX�'���m9 T,Kľ�����5�%�kWiȖ%�b{���"X�%�{�OkiȖ%�b{�ߦӑ,K���]�"X�%�N��ͺ%�[�d�&�Fӑ,K,K��{[ND�,K���6��bX�'��z�9İ:�����w�6��bX�'~'}x�Md�f�1ˬ5��"X�%��w~�ND�,K�׽v��bX�'��p�r%�bX����m9���'�9��/����s���қ��nãusll��Ǟ�.9��u��wzw��6��ia����rS���O��]�"X�%��w�6��bX�%��{[ND�,K���6��bX�'ǽ�FXh�Y�j�%�]�"X�%��w�6��X�%�}��ӑ,K�﻿M�"X�%��k޻ND���'��OXR�fW��;���ľ��kiȖ%�bw�ߦӑ,ı;�{�iȖ%�bw���JrS����'���6�l��'Ȗ%�� 2'�����Kı=�����Kı;���ӑ,K T�/}���r%�bX��=��F�5a��%��M�"X�%��k޻ND�,K�#��~6��X�%�����ٴ�Kı;���iȖ%�b{�_r�Sf�n�#�b��v�k5¦ɗ�{MW!t�T%j�}n�Z����nN4�Nu��@��`:�r6�
)A�a蘝����I]�S�q�,�����M&1r	��9-msmE�`�ѫtփt�A2�,��j�����S���i3�����R���f�(�"��kZ]VP�R�W�X�P�Mv(J��ΐ�"�X�u����g�͓seT�^Ņ��{W3��ݻsd f�@k��N�*Ƭ��X�kshtps�ɦ>�$�)���*fhl��'Ò���bw���"X�%��麟iȖ%�bw�ߦ��~��,K��_��iȖ%9)�g����-asU3%ٝ��rS�ı=���m9ı,N����r%�bX�����Kı;���ӑ?�R"��2%���׍��3Y�1�u5�ND�,K�����r%�bX�����Kĳ�����O�,K����ۼ�JrS��������f�U[I�Z�ND�,�׽v��bX�'��p�r%�bX�������bX�'���m9ı,O�ｌ�h�Y�e�K��ND�,K��m9ı,?�
��������%�b{�iȖ%�b{�ߦӑ,Kľ��kV-&bn��YН4�$͇,�٥��,b�KS6�tۚ��ĬF�ۦ�iȖ%�b_{ǵ��Kı=����Kı=�o�iȖ%�b{��'y>��%9?~O7�*5�f:�r%�bX�����r��U
� Ҡ%�b{�ߦӑ,K��}�ND�,K��=��"X�%��㻞5L�u�������Kı=�o�iȖ%�b{���"X��b_{ޚ�r%�bX�����r%9)�NK���{�Tj�)�O�%ı=���ӑ,Kľ��5��Kı=����K��;���iȖ%�bS�zy�D�u�֦�34m9ı,K�{�[ND�,K�H�w���i�%�bX�����"X�%����JrS�������a\:�M�S-�,�ێ����s��5��UD���du���#G\<��ٛ��/y>��%9<���6��bX�'}�p�r%�bX�{��G�,KĽ��kiȖ%�c?{{=Ͳ�[`*w���NJrQ;�{�ӑ,K�����"X�%�{��ӑ,K�����ӐVı������l��6!�w���NJ%����ND�,K��=��"X�"{�߮ӑ,K���NFS�������������ܳ��K�lK�x����bX�'~׽v��bX�'}�p�r%�`#2'����'Ò���'�'���Yb��1v��bX�'~׽v��bX�'}�p�r%�bX�{���Kı/{�缟JrS����|�w��k��F���^L,7J�5;E��i�w�� �s~M�״HS����'Ӓ���'�����"X�%����6��bX�%�}=��"X�%���]�"X�%�}�۞l��h�fY���iȖ%�b{���"ؖ%�{�OkiȖ%�b{�{�iȖ%�bw���"�Ur�D�)�ͺ,�jk&6fh�r%�bX������r%�bX��^��r%�X�'}�p�r%�bX��}�iȖ%�b{�Ӆ��Fk3F3.��iȖ%�b{�{�iȖ%�bw���"X�%����ND�,/�(��Pj Wv'�����ND�,K�����+6˜�������NJrS��}��S�,K�~�}�iȖ%�bw=�ٴ�Kı;����Kı/���cu��X�Ô��m�1�ҭm��Ȗ�����$\eK�'\R�9��۳_{�ı,O��p�r%�bX��x�m9ı,N��z�?���ı=���ͧ"X�%����g��k35�NjW5�iȖ%�bw=�ٴ�Kı;����Kı;�{�ND�,K�w�6����$��ǽ��B�e�f�pI���]� �'��t��H�����ND�,K�׏]�"X��'�ޝ�	
a�ٽ��rS��bw��6��bX�'��m9ı,N�^=v��bX�؝�^��r%�bX��w3<�L&��˖涜�bX�'��m9ı,N�۞�ND�,K�k޻ND�,K�����K�Jr|���8>���g\�uvv[4�#{V@C��vL�`���#�<����Υ�;(�H�=)J����ss�4�F�`]GL������,n��L`�6�]$�X�ۘF�vy�mq��ۓ�^�Ͱ<'96� �,݇��d5g{Q&��`�M����E��s�y������s<�^�qs��6�v����\\DN�6Ń��+m)�ڶ�j�f�4Ҋ��F`*�K^�a8cq��]��<�nG�܂8�١�֬��	e8`Z�a��ߞ�������0.f���,K���nz�9ı,N��z�9ı,N����Kı>�}�iȖ%�b{�Ӆ��Fk3F3WSWiȖ%�bw�{�iȖ%�bw��ӑ,K�����"X�%�߽���Bı,O�z��ִ]��v������NJrS��_=���rX�%����ND��"{�ۿ�iȖ%�b{����ND�,K�}���5sA�U���rS���p�������m9ı,Ow�w��9ı,N��z�9ı,N����r%��%9?~}7�Gl��H,�'Ò�,K�{w�iȖ%�b{�{�iȖ%�bw�ߦӑ,K��{�ND�������<g�9���b�*K\�w��� g�2�T';52���V�M��~I$�w�8,��r:���NJrS����?��iȖ%�bw�ߦӑ,K��{�ND�,K���ӑ,K���f�����!����JrS���{�}�NB"+,K��{�ND�,K���ӑ,K���ߦӑ,KĿ��[��iֳ.f����Kı=���ӑ,K�﻿[��Kı=����Kı;�o�iȖ%�bS�zy�M�j\1�3Fӑ,K?�T�*dO{���9ı,O�����9ı,N����K��3"^��6��bX�'�v�p����k4c5u�v��bX�'�׽v��bX���}�����~�bX�'�����Kı;����9ı,O����Й�Ԍ�mk4��7��3��76��qo$�4Tz�um��,�:�\+bd�WiȖ%�bw���"X�%�����"X�%�߽�e�r%�bX��]��r%�bX��׼[
a5��L�I�h�r%�bX���p�r(�X�%�߽���Kı;����Kı;���ӑ,K���zg��Y���C5	nkFӑ,K���߲�9ı,N����9�h��QE�DM�:P �7���M�"X�%����p�r%�bX�d��5f�j榲��9ı,N����9ı,N����r%�bX���p�r%�bX��۾�ND�,K��7�5IfMj�3Y��ND�,K���6��bX�� T�����~�bX�'����v��bX�'~�}v��bX�'��sY�����ru�,kQ�6Gk����h��^���z���uu���$q�S��Kı?{���Kı;��}v��bX�'~�}v*�"X�%��k��ND�,K�{�ͺe��3-��4m9ı,O{���ND�,K�k��ND�,K��}v��bX�'�w�6���
.TȖ'�z�N6���k4c5u�v��bX�'��]�"X�%��k޻ND������ӑ,K����[��Kı=��g����f��5i%�]�"X�%��k޻ND�,K���ND�,K���nӑ,K

K�k��ND�,K���Za3Y5��Mf�ӑ,K�����ӑ,K����[��Kı;����Kı=�o�iȖ%�NK���C���Bkm5�Ƌ˹��M�����m[Q�͓�wV�D�ı+5&Icl��nkFӑ,K������Kı;����Kı=���b��%�bX���p�r%�bX�d��5f����\ջND�,K�'��]��%�bo�m9ı,O��m9ı,O{���NE Kı?{�~�з
#˝��O�%9)�NO}�ND�,K���ND�,K���ӑ,K����ӑ,KĿ��_dm0�f���֦ӑ,K?���~6��bX�'����nӑ,K����ӑ,KlO{���r%�bX�Ӿ�6�m֤��f\Ѵ�Kı=��z�9ı,N����9ı,O{���Kı?{���Kı8l@{�G�HP��S��@��<�$B!ږ��Xd	e�i�X�����~b~~Hd$�"i
FH�7c�sHp B T`���D�C���l�C@2�|8';���Vڪ��-�cj�1�S9�W%M�����ƶۮ��:C�� mٽ�����K-��sv�6݀<�ctam�Հ2�0PU
��5m�;i�AQ0�Tk�h
��8�CF�f+ n��@R�J�UR�@[*]���:ꪗ1Ҷ,�+lv�V
�L2�U�9x[v�T���(s���i]\/a�F���|�7c�]G��c WP9�Z�8*�:��V�ɔ��ڮۗ�Cq�ẕ��3��i�,r֐��D'9mtg��>�sӳ�K��(i:��wfx��;V̀�����{� <�]X��1�9֑r�WEm��'�Cz��Nae"&wm8��4�8�'��K����۹6z����s�<P��L�wX5AW7)��X�EEÇ�ll󤎡�N�j�J�S�ˢ�C%�mv�5эM�UYX�D��sJq�6��$v68�W2;L�;\vܹK�8G;Zf:�)��܉-8g(�M�3�s�12΅��ͻ��ׇ�r y�:���P�7%e�Y�T:��
���V!� �l�HJ�r֗6h���;�tb���VM��;s�q����.��qj�K�R���xZn[h �7E/nݻ�\�vw$a8�p�s�tv�ܸd����Cͦ�
�e(H����A禮t[B9@�S���ֱ�(/8w9�N;n����#h<;^M�A0���`�u=�179����R��9�U�Tr�*kRtʯ$4v�m�An�CP����	��7g��<���s�8��G��Tq�y{6�k�hn����{g<1��m�͛��!��͝�pUl[\��ӳΤ��qP� Bc�H��H� 8pVV�U-m�O\�pOI�Ƨp�!R�pL��흲�rp.�ʶd���u��x͓�X�O9g�D5�-mpʱ����/Xn���V�d��#���gG�!�gg(�s���\Y3�r�pl�{N��pg۬������3Ukm�*%]m�F��䟾i,@�|��G��DMAP�#�GH�}��\����h���̲SaV.�I����B�c`]"�m��]rb�����̯b��7%������kRZ@�j�5vWn�����/Ni�Ր�]&%T��[y��Cd��h0j�IAɒ�� ���]��a68Lj7-�a%�D;�v'n]r�S�l�����8�[�!f.0�8�[j[�v�����o=wfjn8R�����(A:�ۘz��{��z^;[{$ީ�F��uD9*�L\-[\	���v���'q�k���ֳF3WZ���Kı;����Kı=�{�ӑ,K������D�,K���nӑ,K��}.�֋������\��r%�bX����iȖ%�b~�}�iȖ%�bw�߭�r%�bX��]��r*
%�c=�}��43����'Ò���~�}�iȖ%�bw�߭�r%�bX��]��r%�bX����iȖ%�NOߙ��0�H�-�;���%?�D����nӑ,K��u���Kı;�{�ӑ,K� T�����iȖ%�b^�=��asF�٫���[��Kı;����Kı;�{�ӑ,K�����"X�%��w~�iȖ%�b_��뚷V�Z�s�F��n�
�m���� ;M��d� ��3E��IVvrI'7S���nG�7'y>�K���ND�,K���ND�,K���n��AB~��,K�����|9)�NJr_?���9l�x73.M�"X�%�����!P2%�bw�߭�r%�bX�����r%�bX����i�(��bX�Ӿ�6�m�HfK�3Fӑ,K�﻿[��Kı>�]��r%�bX����iȖ%�b~����Kı=ӷӍ��Lֵ���֭�r%�bX�}�z�9ı,N����Kı>����K��;����9ı,O{���ִL�5���K�]�"X�%��{�6��bX�'�{�6��bX�'}��ݧ"X�%�����ӑ,K��U�zY�7��e��vu���`fG.�k���kq��'oT���h��r���$�g���8ql�ZѴ�ı,N����ӑ,K�﻿[��Kı>�^��,�"X�'����m9ı,O���?��Y���MM6�5�iȖ%�bw�߭�r%�bX�}�z�9ı,N����Kı>�����,K��ތ�.i�K����[��Kı>�^��r%�bX����iȖ?�p2H��V����k���K~��X��2�I����v���L�vL��K��?��z����ɟ�� '���g��E�Yt�wX�X�-`�E�t� �J��4բ���3�95i�[2s���'i�V��t<�:�s�闏<�]$�]2�cw_�������,�\0�&V:�C<�+c�wN��v��"�:u� ݓ+ ���Y��W�+�\��V�=���~�2���y-�[�`��:��I �e�t���&V�����"��
���ݛ�s�Γ.�3Y�5tۧwX�-`��t�+ ݓ+ <��)V�\��%�Y�7R���UB�̔	viF�J<� ����.�v�����zq]�k ݗ�L�gL��Kq`�`$�ue�;�� ��+>���}��l��� ���U�y ߣ>g��E��ƛwX}>��?t�z���%;���'�� ��e%WI'WWE�'u�~�n,�\0�2��2�	���[ۺuE۵�vˆ���ޟO�W�;��V����Uz��]�4;��f�I� �t���D�3c[���Nq�lε�kSLh/��KY�lͰ�9�T�]�%�Z���;��)j��6X�3��h�eS'f�^������:��uȣHV���h�X�NR�hnk�42�Q�.�]L4�.� IJ�B�+k|{[S�l�K���C��`�Nr��=,��n����7%�*l�%�k�Z��%�f� �vm�bӑ��\OW������-p��y��=.��.�����Y�=��΁���vt�-ŀvɕ�N�r�@:n�WWH.��2��-ŀvˆӦV$}������9��ګ:�=w��~��� ��+ ��+ �ԇ��]��-:�n��.N�XΙX���?N��YIU�Wj���ـt镀l镀~�r��.�	�Ӕ:J�\@�bfk0�e
���VgXG�]͘���%���mKX�
h�&�ft�~�|�r��.Ip���*�]$��D��sF�����1 �'���́�\0�2�	���]7wwN�wv��2���nɕ�~�%���p�v�ݫ�w�u�t��ɕ�~�%�w�V6��IQN��e��v`�L��9-��2���xx_����ib�vmtrl%=e��z��Q�<�]b��U�ͳ��WUۙ�+E[��������ޙXI2��&V9��v"��ջx�L���`�\0�x�-)VRUe�W~���:K��e���^�^Ky��&V M]R�t
�4�ـ~�2��n,w�V�\0��U��I:�T���r���+ ��,�ɕ�rt�;�I�����۴��<tލ.p�8v�����ԡ�ru�kk��V5;�efʳH*߀~�｝���� ݓ+ ��;�W
Whm�wn�
��:9m}^lﾺ�'}5�n���'9%��g����K��2�[�?�ﲰ�j,v\0���5T��:mY�鳖t=���$�����^����ܓ������|S�("�0 �1 �@"�+���f9��v"�춭`�E�t��&V�-E�r�8�;�����0kקѷ&+�O���#h�	������[��$��obKb1�rߠ{���X�Xl���X�xE�+�,m�� ݓ+ 햢�7\� �&V}���	�S-]	����bwX�Z�`�E�t�vL�mtu��E�v���-�X�`%� ݓ+�U{ޥ'ؾX����mӻ���`� ݓ+ �7w�^�s�}��m�Y�V�bi��v�sʝ�Õb�����\�:�G	N,���g+̴�%�i�T����`@u�R#]�˒��2�7KU0��l�l����t��AFh��4w�W����Ts����.���ظ��즩� 1�30��#T���:���=���ԕղd�h��.gڮX���l�;wN+hp��LS��j�l\��Z���d�rBcW4��3�X�f厅��X�/LV誜/n�͹�h�	�e]�ɘ6
�1������;����p�������}������a�����9g@������p�:9�&VԔP7N쫢��mZ�7e� ��,?�{����y�?�������Hҕ
J���WH�-ـt}�&V�-E�n� Cz��t
�ʶ�ݬvL�����{��^�W����Z���`E�~�+-��8��s!6G�ϑ1�]b������	ϭ�ּ�a�n���X]����ft�-E�n���X�X���)¬��z߻�/|�d'���4�P����o�ٹ'���7$��uܻ�d�9i���}%[v�+q-�{ｘ�X}U�Jw��Xs��M��*hVa����NI$��{���<���X�`$��	�J�	]]Yn��wXl����XI2��2������(U(�K��0�x]�&6��+[�عU�tI:�(g5��'ǰᴪX��v��;��,��X�X}egV��VE2B`�D�]���2��q�uȳ����ĕ��t
�ʶջXw�e`��X]J��m8�j�) h� �F���
1(I���D�E"�W��;�c 0B0�T�� �m2�BRRS?~���'�L%
Z�	�� r�b8�i#!8��(������
�*A)+0(R� @�J��$�@�4n!�I��$c���@ޘ,�)HN�`�AК#lF��q��(�Ba\H$Q"A A�@#1$Y�XE��@�2�D��``��A���	a# ��6�p5 ZjZ�2X��XD`H�"�!.�e�@L�eW�RJ���8,]q�`BюbĄ��JX�ki�!rL0\!���#� �ʠ����9��H򤬸Ą�#	���	�"I���e��i!X!��9�1M��Ex��7�
�(����ު����j�;�E�Je�t�N�lLn� ��7_E�t}��[�}����β��-�v�x-�X�����?l�Xt���ꭩ3{)��y�����V��4�j7��u>Č+C�mi�׮;O��9�����'�|��&V�.5����Uk	�� ��ֿ�P�t팺�@�� ��e`��X���e`i%�HWactݻ��;eư��a���%>��{ﲰ����]�EZ�-�X�^�R���'�}��~�2�
�l��#Q�Ueӵt��;XI2��V��~��N��k �}���ݤ�l��ӓ����S�^�)����c������L<;��!+.kxR<�H�vg�>���΁�eư��`$����v��4�ʶ&7u�v�Qg��UU6H��X����X�+?��>�:�B��eۥත`�|��e`�L������m��wi����UT��}�����;�Q����$�JT4�Z����wX�+ ��UT�����ϖ�wf��g� �h� �"U98I�_7��|�S6�-�� ��2��������i"�nu�����j�<m!�(80 ��>M�˶qÎ�sh��;N�a,��a�v{6��\�\ٍ�]v�0��;Q���3�y
�8�r�N3�(8���ns<]�s33��ЧQ�Ɨ;!��%�s�kBz�K����3t�N4�n|��]F63(���2Mc��\3HWd�>3gv!�x�o{��r��X4�2v�կ*:y�u��)t;9��Ӭ,�
�u�C;m:7e1[H�-V�9��x�`$��*�����>]_|һ�j��v��"�6I��nɕ�o�tj2��Y~wt�bv��e`�ea�UR]�� �|��tV�"���ʶ�wX�X�.�`$����X�I��iSn� �%� ��]������e`~��g@�/���Uv\.������dı�KΘ,�\㡻i.v�-nh6���'q������Ҫv��"�6I��nɕ�o�l�W;lM[�O�ݬ	�����H��-�}�lܓ��k�rM�"�'K%*N�ZeӤ��2��\0�=�Uz��|��ﲰ���Ӥ't[N��wX�UT�g����`$��7d��"��@ӻ.��ue�0�"�6I��nɕ�o��'��x�3�͘�ah��q�r���	K-��hM�3��8��M�2�d��wk�������-���}>��7d��?q.����C��﷠{g�oq�H�1"궰�2��z�^��6_����`E�ު�H�|�E�t�Ս*m�`�� �r,.�U^U^*�U���`�e`����*-�WwJ�-ف�^��|��ϖ�&V��"�6@�!�cjӴ�	��6>� ��Uw}�������7\� ��{�K�U�?�+.�ݭB�&��������NV٥�=k+{	�;9::���2�[�]�4�V���}��8r,uȰ���"�JN�N��t����?q.���$w?�X|�� ݓ+ ��� ӧl��J����7\� ��,?��w}�V���0�-Gh��]�!Zv�>�{������`ed��N�rH�`�L�  :��o{��ܓ���팮��b��ݻx�X�.�`������x���݇�����s[-�9�D�uخ��,�eb��z�u�U���Tۺ�7Ip�7\� ս�&V$��y�I���P'k �r,V�x�+ �� ށpC��;��N��z<�ɕ����K�|��>X�*R����]�ݼ�ɕ�n�E�n�� ս�P�cI�E�I[��tr,u�X�������ܓI������Լ�L.���\�m�8h��*��m����V�Inhͷ3�痟A���M���i�6jX;r��i��B٢ǇDW.%��t;��fPF�d[�a0��M,�6�0�`3%۞�jŵ�d���s���T\a�؛u��;��;:t�0r�&�p�m�]�a���	v��e�ݚBR'o������B�:4_����l��)M�6�b5��䠙�� ��@��:5��ݱ��Մ��]��%�,5q�3 �L�0k��}�^����t��{ﲰ�\0�Z��Qm]!�M[v���`�L���u�Y�W[��t����.�`�L���u�X���2U�lc�X�cwXi.����`�L�{���T����h�7k �}��,�ɕ�v�E�E��P���ZL���\ëa��g�ko,�5\���:sx�HPR�؛6��\ށ������L��r,u�X�*R'Wm1�n�`�L����D��X����`i%	�4��V���;G"�7_E�o>� ��e`�u ӧWE����7_E�o>� ��e`��`��.�(���ƭ�X���&V�9��,���0o!�lyYMH����#m�n�v��ZS�x���e��W6�W4�x���ށ�d��?s��u�]_�j��2x��Ʈ�I1���>J����,k��&V��Vy�����xI��}۹'߳���)@
0�,bV Q@ ����vnI��ze��;j�(��v�� ��e`�\kꪥ�s�}���1:�i�`�wf�d��?t����,��%%5t ��n�t�Ƭ�9�t����%vNnR��J�6�Fۜ͆�ЛcI�Ul)Z���K�`���;z�~�2����uv�]��v���,���+ ���X�(�`P�Z)Ս[v�޸`�L��K�`���"���z�˪��ݘ�+ ��F���`����=[*�@"E;�y�$��fg�n.�*�&7u�~�x���`�N΁���mՍ����!u���.��mvщ�s\l����JV��� ���z�e�P6�����;��~�2��� ބY@�ڶ��`�pϒ7��+ ��_<u�XId��lc����?l�X�qG�n�� �� MRP����j�R�wX�qG�n�� ���d��"�(iӶU�j춭`���;�E�~�ݛ�s����I���"����B�
 ?PP�i8�CgAq�Z��u.�+Kd�7�/HBu ��1� 4��H	��e ���a��"Ab�RD��$)(B�X��@R%#+m����
��!a
V�bQ�A�� �@���BB6��$HR��)mH4%B,6�R�)+
	��qX�8�jB�E�HA� � @�ʰ!HȰh��xH),��� �C"� FTH�"HV��,H� JR�%aI`@���t�}��E��ݹzr�)m�جB�i����m<	��\��m��kW���X������qͮ����UW�g�V�;0� 5Um�P*��NS��_��e��P+�[ 	u� 7L.�iU��窪50)�#���-� Nk�^��'E�m���Sb��nnتT�T�C�dck����H	��a5�b�c�UO8�ln�X������e X������*j��\�*�}]e]�D`x�v�ml2������A����Dl���"�d8���UGV�N��cȆv�.^ջ\�FĄ�X�
�N�%��2Z�Y�<8^��EGC���m-��fl�+�V�%vt�x�8�1�Q�X-�k�q;r��w���DKv���
;Wgl&63�%'8��'�����K5��ή4"c�$���6�"�-�C����n�ڝ���'A�\��c5͹�b���pW�2�SJK�m%gfYI�1��Kۺz��3qɑ��cPI�E�\dtF��`gS,݅��tgU��c�����AQ`�}��>�֖ˆW���������ۂ���R�8�g��vuǱ�\s�b��uD@čgJI�m�%�u���HĎ��n���Ҝ��F�v۷=�ӂr,�c�n{'-3�ۭ�s�vۅ�����m�ȍ��]��nC=�?|o�G;��J�TaJL�ٍ����v��MO�`����
�l2��瘷fUY6�kE�쥂ug*#�Xڻ{=���u����.�W���������2�/�<�-�ha*�Ѻ;$v[bрT7U��@l9�\Zq��g� ��C�[��W
��P����
�Aڍ��i���r�nN6�`�Rqj�7:N�W��إ����6=�qģm�m�cnӝ�!�U.[�i[����Z�p�UJ�Ԩ����2��Ұg*�tS{	Ϣg���[c�s�1��p^v����:�1�9��"��ZfK����n��K&�+�@��Cʠ�@�#�?*��W�F� ��'���@誤�a�e�g1�s�ƚ�[�쉤��2;�/[���#rmф�k]�#���
!�wK���f7 N���l��ָ�i���񺑉�H�M�Ͳ��L����rRKH4�в�@Yp�b��u��2罻�ˠM����´�Ѯ��%F-)s$����,[��qb�&�w�
:v^Y��#=�V].�i���ǜ�I#��{�9�t�ժf�A�DԚ�`�ȻZ%��&>n�M�M�+
�
֘Wf��7���ɕ�oKQ`���"��) ��5ue;.�`�L�zZ� �}��X$i�	:bw뤘���-E�n������JG�� ����tfy�M�j��P&�`���;�� ��e`��X�"�m�vմP'k �r,������W�:?�� �s��<���u��T4�s��Y��k�B��s�:ͣ�Z��Kz��pP�N�u����6�`�e`�(��"�;�� &�(I4ݲ�`�ڻ�y�o{���/z���1`�E�nɕ�{�Z{O}k���+]�?~��zs�`�e`�(��(�`P�ZXշk �r,vL�y���XU�� X&��;.�`�e`��X�`�E�oIX[vʱ��R�q=Yb"'-ngu��5�Y��#6�)Cq�� [h������������~� �r,�Ȱ�2��љ�6]�Wa@���n���X�X���e��;j�(��}�w�rN~�vnpzJ�T��#���k��,��yU�Ӷ2����?l�X�7_E�w>�+�n hy��BL�K{aN$��U�z���~G>X�+ ��qU�L�É`\�r���33�3u#[r.��n�N���2E�v4P��.pF��ށ��,��X�+ ���X�9 �Z�`�+cv���gު�URF��e`>���7_E�E]�R(Ut7wk��v��&V��ư��`�����<��߮�cwXW�Kg��Xs�,��X�ު���Q�d��7�3<�&�j��P'm`���;_E�~�2��.5�~�q��I;B`�7\��>�.�]p`�G`��,ei��o;Zw^���ځ�ˠM����
�`���?l�X��7_E�t�'�X�;v��Hn�`�L��K�`���;_E�T�$���wj����?t����,>��z�(�|����:9Nuwv­;��`���9t� ��e`���	)� �ںt]��ݬ���d��7���������[���5�\9���w;<t�v�eˣ�VH�
[�)�CZ�=ce �i���k���d���Mq�t�03ƆH�M]����ڍ�&q9�JmGk�c\m��<l�u�r��)�hr��"�:�n�.���X^�Dd�����|�C��]{m�ZE�<�[,�R�1i�jƃ\$���;zB�BX
b��Yrj\cl�xm.�.O�w�����[�J�U�#NN��ԛr;�U�����5k9��;��c�,�;�d���2����q2�߀����k �gG�n�� ��G�ъy	��)$���tx��ˤx�+ ����I�ڷv�x��ˤx�+ �gG�v�	�6�ݴP7k ��G�~�2��H���`��V'Nݦ��m��?l�X�$x��]#����sX�r��v�կ&�����U�ggT<�һmt�v��	v�m��+E�]�o2G�n�� ��<�ɕ�t}[�	��Ѝ�3�߻����C�s���H��X�:<Jj@(v�ή�ln��t� ��e`�����`WG)+���S�v��&V�Ώ �}��� 7���BtƮҤ1��y���,�9�d��?u�C�I��m/][F�Z��ɲe:��]c�E����!�T����v����էn�;x����X�+ �gG��W�6C����wv��`�,�ɕ�o3��7_E�~�T�E����.�n��d��7��ᾪ�^��{�z�,yȰ�RP+Iһ�V����7������?s�`�L���r�)�wv��;C��n�� ��E�~�2��tx�ԜNK�u�m��V��abgV�`����L<I��%u�N��t7of/=F�����X�+ �gG�n�� ��KB�n�1Ywk ��e`�����`�Ȱz8��'�J�C��7������?s�`�L���fz�'M���(��}^����6?�w$���f�A����`"�B#�!�H�|�
cŃ��b�D��l! bb�HG�W�	��>�M�Z��h�n���� �:e`�����`W��z������h�F��+V�\VQ`t�M\�����J׳�ym��Ã3ǫX^���ԥ� ۵��}��o3��;_E�~�"�	�J�t��V��� �gG�w>� ��G�~�e`S��;�AV����;�E�~]#�?I2��tx�k�xwJ�쫶7k ��G�~�e`�����`WIb(N�ZvX����?I2��txs�����'�s���~����su�Jm'�E$҄c��)S)ɥ�R��	G���$�e4BpԺ�QL�4��+I�r�۲�Ma؞�ѭ�n1Z�,f�h�lZ�9�Fy"�t��Z�0j�� V1-��є��K��Sc8ۈ�m��͙���_��=�� �Gw�.�tl���륭��Ș����{��7h�Ӻb��ku�1�6$�z�	�W�C�.�4eճ2eֲ��SV�f�봏\ȗ�MTN�,-��[fi�.�؉i��I�R�j�������,�>����ﲰ��3֩�حڲ�o �}��,��+ �����J��]ݦ��`��X�&V����Ϣ�?G*Ri�-�t$[�XUU-��V���w>��UU/�>{z���`f����:������`��X�&Vt�r��;XX���5��:���%��0�ڊf�e��\\E�.f@&�+B77W|�E`g缰��Vk�� ���4桚ə��'?gݻ��b�d�d��7�(���`T�R(N�ZvX��k �$��?s���,��� 7���h�n� �ϔxs���,��+ ݑ���i�nզP&��Ϣ�?k��L��>��%J��C�"r&�bxE��v��`�^�z�q��V0�mp�ј���ř��(��~��`�L��>Q�ϴ�Kk�\�dQ�����K{o3�~��<y�X�} ~$��un�CWu�~�tx�谝�_�{�Ao�?χC�z �c�?<	��<? � �:���Z�6*P�V"̕��#�;��CBI�q5j7����B�� �$"�`B Ā�a2�d��$�e,�K$�P�H��1��#+�Y"�$ $H�,��� 	X� �	��2?����FR0���H�i�&��!�&ݬ�$صb�`E�@`��I��l�֠��y@�O�si���^��j�&T��6�����HBL!B"R���#(^)�"E��� *���R+� �GP�;T��(��](|'� Њ�%�ٿ����vnI�s��G��wj�Ӵ;xz����s�ls�~�2��Ώ �Mt���W�e;cv���,�I��~�tx����y�*
�i��������Zڞ��\�q�1���$\�\�B�rX��k �$��?s$xs���`tqZ�'�Vҫ����Ώ �}��E�~�eg��RGw�5��M*n�mv�	�`��X�&V��#�?qҲ��b��i���X���L��3�����G�P��R�D	��R�J�b߽�}w}�r�-���]] �v��L��3��;�E�~��`�QD5t �mI��[1��������2s�c&�ڏ+gq���g&E`f����:�����Ϣ�?s��L�.�
<�;�T��;xs���,��+ ������G�MO���WNҧv7k ��� �$��?s:<��XU��E	�E[�T�ݬ��+ ������`��X�V�I�U���i���3��7�E�~��`�L��z�Q�zrBrBI'9��z�5t�[]Bcgfv��$��C���KY��fyz�K�w3ڻA���"��n�.�n7�pSՆ,�rr9���M(m���a�"�����e��۝	8ٳ�Kh1��s����a�;:�nYv�:�	�ˍ{\m��`$%�#Ga)]EձeGJJmr	L��6�&f@��
���3nTY4�[��V:�x�n�s�4m]��G��C��ަ�۫]�Z\�]JW���.4�.���74l垊�;4m��ʗ��3�m��o ���,y�X�+ �̑���Y@����@��y�X�+ �̑�Ϣ�6J�E6Yv]] �v��L��2G�w>� �} MRP&����vC���2G�w>� �}�I��tr�(�t��Zv���w>� �}�I��~�H�ʢЫe��ڡ�����m�z���nBn^�U��kA[���X��RWWCa��+�iSvݯ�ts�~�e`����,*��"�ˢ�ݪLn���{�|D��T�5�M�7G"�?s��8�P'⭥WCM�`����,�>� ��e`:7����j�P!��7�E�~��`�L��3��?���~�v�N�wh�N��69��?t�X�gG�o>� ���õ!f2j9�t������\)&���$I��3�s�ܜ���u�k�*t����?t�X�d� �}��, ���M'Wwv�����2G�o>� �}����P�
<�;�T����Ϣ�7�����{y�!���ｳrO}����>�Ʈ@�v��Ҧ�X�`�L�y�<y�XU��E
��-ݪLwk ��e`̑�Ϣ�7�� ޓ7\ܕ�j��恧��D�]h�(�mČn�m0M�%1��yl���#�n��.� �d� �}��X�+ �:7����j���"��Ϣ�7�� �$��7����zVP[m'bwh�Wk ��E�~�2��tx���O�*Uj����L-�X�+ �d�nI����rE|�"`��wY�]�r���t�������`̑�Ϣ�7�� ��e`�.�u�n�w���dm�Y݌�ֹ5�R2�p�6R*���/���!ͦV�nh����{z�r,�I��o2G�t��x�V�iSvݬyȰ�&V����,*��"�e�;/�˻0�&V��W���� ���`tqZ�O�[*ؚn� �d� �}�.�&V�to=käի��E��;�E�oK�����7�#�;�ꪥ#U.�p��]��':�� q4k� �͵��sIIؕ�$y�$Xe�UY\�5�Z�]v�sOb�y���lM�k�^��o������G�V���!�5I)���v�L��0�E4t����X���ȶx���K	��N[�"���Z�	����Z�6C)���r6UIwd�,��u�
F�ܺve���N<�6n��`�%����d��Mk2�Z�?���A<rO���L}���f���KE��ۅ�80���Nu�9��]�`��q�]ͶҠ���(ڀ}���~�e`̑�ϴ�K���S�BLx҃��-��0�H���`��T�	��ݵwIwu�o2G�w>� ޗ��+ ����ӻ�Aj�E��;�E�oK��I��o2G�l���ںNۦ�X��`��X�$x%޾Ӊ-���#x��1��,qI=��Gj�7m%���f!ǉ�Yl������S6f,��2��YV�&]���}��o2G�o>�����O�� $���P'�Ս&���O�d�sw�`��YZ�� ����
1Z5%{��=_�Uz���� ���`�L����zׇI�V�o �}�.�+ �d� �]� -���wv�v��p�?t�X�$x���}�EZun�]�X�+ �d� �}��X�.���E�m0q�;Vզ^ x���t^�AH�	���6��n+��s��0.�L�Y�uY��c�w@�}��X�+ ������۠�v"��Ϣ�7�� ��e`̑�:����v�7m��7��	9�{�s@qD�O�����-y���Ns�E[�P��YwW�c�X�&V����,yȰ�8�P'��M&ۺ�7�#�;�E�o9�I��~�+�P��.�ɣX��;8hɔuZTe�1������m��V�v��ך���.���,yȰ�L�y�<�wL �m7j���`�E�~�e`̑�Ϣ�7��AQj��un�]�X�&V����,yȰj��4�;���B�`Uz�ԺY�� �ϖ�仓4���b����ܓ���C0��t��]���X�`��X�������K����J��EfT�u�U�km�9nx���5A&�t�WL�E"�)�\���in�m��7�� ��e`̑�z�_�ts���&YWn�.��?t�X�$x���p���@�We$�N� �d� �Ϣ�7�� ��2�ӣy�^hNڶ�x�}�.�镀o3��6�L@]�۷wv�v��.����{��I�;�ԓ����rO��**���**����� *��**� ���"����"
����
��򢪧��#� ��E��  *R�`*b*AX
��U��E ��DV�P��D��AF"�`*X
�F�"���E��D`*H��P��@H",B���A
�  *��AP��DQ�"�D *��A ��E
�@@�"�A"*
�P���E "��
�EH
�X�,���D@�"��`*","*��F� ��@ *X", `*P"��
�V� "*AB���@b��P�  ����AR���EA"��X
�P�"�Q�,@ *@P�"�E� b��",EH
�@"��R
T��
���D�TU� ��QE^(�����
���**�� ��������
���PTU�(**���d�Md�����f�A@��̟\���@ 
DP H��� �@�
($ �UE�έ�  �T�P��TP��3X�Zd
E"�ZJD �TE!i�@ U PQ@��J�J�  b�(�  �   0 rd�
�B�ms�P7πy:��F�\�;�=4��l�����{�eA����# �05���b��\ ,�=��� ����>��o`y�y���  .>�}`��GT�� z��ʸ�En-Uzב�^:}t{�Un��UJ��G�����[��t�{��y�@��f���w{�g`;�@��$ `zn`� �����*�� �{ہ|��s��9[{��{z�I*�@��9vt�V�Тp��V�p�!�wX�ԅ' �ށ�Xl9���n�P=�>���t�]�� Ā4 7& ������Y��R��S�;�J
)
}nziJ\�ҝ70���KX��Ol4�s:(6t    ��� �K)A�w2�R��@�����k 
Z��� M��6R�z;�Ҁ-`�   ��$}d�  �s�@����8� �Q�M��|���\\]�>�݁���}��.����  C=����v�J��x����fy��]���m� ���&ã��|  �DmRR�  D��T�  Ob�T��"@ h �?d��J�4�� �Ѫ�f�J� h ���ʔ���)������k�����2N��]��w� ���j���*�TO�U��*�¢��AT����_�2Y���L�bs�܇74�ĕ%b�˘�fH��Y��r����KgY�-|;�Mg�N��Gͽ;S�#"Y�K���"�C�	.��q"B�`K�P�H�di�!LI�� ��K��$��$!$���F�M);��q`i�$"�b`2Bcq$% aBe� !�L
,�����bԆ�H�I�P+v���B�0��Xh4�HƸ1�ĴĂ��1��aHYU>O���U!@!�D&��4$Ϸ�F�A�k��)B
,��H�*�c��	�C���_gۓY�i� }&�Hء(�:�� �B10 �@�I�����i�H��S�A��4�XaBa�08B�,/!���M�������O8|!wO��|��5�sn8s��9���������޷��_���O����bC�,4�B�2�H���L�riy�~���cl��,N��B��a��hu�EY�va,���#���o9͟^m��8��E��H�'�]~M?�H�� �R�� �4�&F�IL!p�%�YdH�e	L�$r,�s��6쐥�l��V��0&�q�;bCi���O8y��5a�k��8ۛ��%	FP�4B!Hck�)�(Fҟ���P�a�r%�%���XK 듥�O4�FX\�ŀT� �Da!H�B���p�2@�pc����lA��W�e;RZ�H�D�XY�9�oy��󙭤y�ԳxS>��T��SMHY"\ԛ7fkx1�@�Y$l�#���K�M����&�́BX�P�q7��f�!+�*Zh�@��$����xW��E����IIi/�5)��Ml'������$��0�.�ۇ#Y��C�͛�70Ѡ��щ6G�M�ro��Kۑ؁v��L�Y���'�<�^���<���|�>o����=+�i��5�?m���>7ϰ�&o���fkd��.�q����k|!
`�aani��D��>���BV.P��{��꭯QZ�=���AWE&�f��
al�ӟj0�� H|�hĐ�u.��`���Ͱ$p���0`� N2H@�0��T��spd�k�dJ�8Ct>*y��hBBC�V�B��.�JD��j�!H��MJ0Á�A`H:٬���L4h�oKr���!��`B즥�G,*B�t�+��CN8�0�V4HD�:�	u�1 �i���e!��!�H2��7͑9�M�
fo��?����H^Bk/Y!\	q�))IK
�"���w�2��OYY�ua#.WNͫ|�n�S�0�h��F�(B�f�A#�(E�
Mk\jA)L���!���I��¥5�kS2`h��4XO�H�v����HF�&�mX�14�]�8#C�M� �@Ӳ�*S�,�?I>���w�ߙsF�B F��i��7��4S6�����!�y�37�'��'���㉼pa1,&����J�{K�*Ɛ��)�.dނ氲$�Hƌ	0!f!��� ơ��\����a��- HN
�xql�	l�$&bP�� �(Ƶ���e�Kn&���!puu�t�.H,��#��&:����
R���~�N2�SZ"c��+ *,��K��)�X��&� h?�6�$�rC��w���O�Y��hȕ���{���	����p�c"B"B�$d͕c2@�)F4"FZa���F�;Xsx�f�eR�1������3z��.@��D%���C6Kg=l���b]�K�;4��C�dG��vF0
&0 ��K�
R	HSj�! i��I
bN$K��O'����]����$�[fP���&�0\>��ݚa��.�a�M�7�n"H���ŁV�@B ���1�B��7$/:CZcY�̺��Թ�c�`K��w���(�HS�	w��h�!`s�/�S+������S$�)/8q����s[8|�R|��1a��xv&��c���%�H'J�����C/p�sA.�r�p���%�����2�"U��I�BLY	����!�:�3��u�iC[�y>�����<O;B\�$.�+�����X0�.�̈́����y��).����7\�)�[�f2�@.;�ė[�-��w�;����F��l:!�F���c��p�L$X����A�K�\��	�}��"FV�B�+;�����U:�_����tVw2��r?�B���H\��������Ń\I��	.���8�&��v���$#�ą]+��U�V�!8��|�L�-����͜6S�C
���4�;j��F�H0�[J�\�,�'�~p0���ɖ�v�R
�v�#%SD��]fI:%ѣe��I,ь����v<�^��<��g��.x��G���B�,�r��/�������@�<$�� �C��o�����K���4�a��HbK��3����#ݤ��A�&�#�<�4ˁ�r�aBSL.�Is���B�7��as!��_����C��q�ٛ�B��&��w=�!|�C���?����&��E"1�X�
���g�o��g��B@��.`J�$�(IB
Ro'��k�CN���ϰ�	}�z�c�A�t��i�����\�IFW=�Z�ko�;·��>t:Q�R��q��~�����;.f{�՘QF�s5�re���q�bČq�Ё$�D��u��+�\�.�ϵ���&`pt�Rq!���Y�G�i`Hst��K�.0�	5�lLqo������tnY&󡆸g]��s�o����U�;���N��}���9&���4C1�����]ms��ﯚ�����o]���R�����59�/�>8��)�1������͜�&��$.V�!��J80Y4�(0t��s]�.^kL���D���
a���a�f$H�(Jbơ�2p�-6lӜ����.��k��Ys[xK�[	��0�\	�\8}� �>9�A�љ3����N2�.}�]`Ma�O�vq`K�ܟ��hG�!
`B��s�&~!����ncp������a�"Sk�@���0J���}�w��B;���F��4H`��H�%T��%HR0 �X!V$`1##,�!VRc
1�l0�!d1�!��B�hA0�! B��E�0��"8@�0cX���,��H�+X��4H�#LX\� a�XL��X`J@�A��"�L�n4��i�8maLR0�(Mc�Eq4�6K��k ӀB����Z�hA�:�8�ǊIp��8���K�0�1�F,�����0������J:ep�n4���/u����<	l�3���3Жe�.h�aJ1�(�Tx��&SN(�`|A�!�Ej	
!�XĠ�`�a#�h�@h�j�Z*��˷�Ј�pP�p����S$t�!��BS����u������]�> ���n�F�6d��2�v�6GA� .�H]/��#��A���æ�C�q����e��ׯfHN'�t\�����Km4�`t	%�0�DX?;��`U�A��H�jSX\7�&DX��_�n:�)��,aFB���v$��|�4�����5�D������f���e�!I"I3d)�)�@�0�2�&kWhDcĦ4�IsE6�H��HĮ7[��NgK� �3�0�x\H!!���H]n�� CLR�$tl��A�@��>��n�HHI��FI�P��c��$d)
ā��0�$��A`0`�##B$!�+ D�$~�(�Ƅ��J�J�!�B��)-�}��?)7��|  m �h    �` -�$ �`     m� m�5��$}��l�d�I�P��d.��]m쌄X]m�"�:�m�-5�� -$��m�ۖ� �     �jA����p  �  �Ŵ     ���i!�9�ր8 ��\ H�4�����$ 	�q 	 &���m� [H��6�T�J�U+�ڸ8	
Vհ�l�� �C��6�H m�i��Ӄm�m� �� 6��TZ�����).QJsI�u�$��%5����c-s�t���1v��pR�7�~�1��]��9񊛰j*���m�$m�ܐ۶  mKE���֛>��l�ZV�s�@* Hq�����yWvZ���Nk�Đ��ڐ�9m��  m�� 6�q� ���`  �e�/���2�P���j�9.�]UuT9n�����IVY؉訵���I0 �l�v�]3�m��(%��5�E��R��y��p�hxO.��U�/UM�{
\����	��ۭ��G��t�#�F���ȴ0�q�ێ��uq[ Pu�-�.�fE��� V�&^��jv�vCwj����m�u���Se�$s���jI.���-*��1�[�U]�m���_���:	:@l����^��/�����uP
��XԲ��Z�5��kGM'i�Vݭ�NbÄ͛�gD�j�� @\�j�Y��{]�`�Z� ઠ.֔X�(�/�s��8$H�ٵ�� %�0�+�K��j�  h��faE@��s�
��`���z4��2 $��)t��f�t�I�[�(z��Nc�w�z쑖9��
��F�q�^%Mk#[�[q"Nqm-��x�`޶z¦ss�˭�J�H	��yzn�-�e�tJ�`� ��` ,1����u;q�u�:[($IZ�nl:@�����E���f�H�m�M��WF �  �6��z5����`U�k��-��h���P���jh��Uu@���$p��5��^f�U͵!�\8�U�/kם��`�A��:�lդ�[H0�ۀ��[%�i-d�]�Uz�^zV���c��oWNi��uؑ�m�p�#�g@[%-��mmZ���Up	]���l��<��-󃓧����������%�sʷ'��c�%	��֎nֺi����T��
���R{��#�� 5,Y��c�ns���R�z�v����(��z��z�*���ej�ڻ�j��m��\�7� r%���2�v�W��s��]���h$m�l9l�þ{���-��K�Sу��,ŧ�R8S;UT  [M�[Rm��7�K�ܶ�F�$�t� *ʡɞ���U�/]uWE{Tu�$��$86���;&��m�^��Ŵګ��YɬH�J�K3� U+�2�-V5��k�j�Ғ��UV�R�v�Am��Â��%r�k,L�m��k���m[�#��p[BB鸒 [%���    8�z9�m�:8U�^�B���v�(X��P ���� �    �m�`�յ%�I�N��ڶؽ9�  5Z8 ���m2n]n흝�be��G���%�6�-�m[v�,I�����	Jݶۤ�[tNH�[IM�v�lR�̪�I��T�l��Dk�v��Y-�lu��l�i1 m��Ͷ�m�|�5Ul����^�Aɧf�j�겍֜H N�[D�$�Un�QuK�u��`���P��%��E�����A���ͤ�6ؒk�o̼��׋z�$t�L��-z�]r�����*Ղv҃�mPUs�Ӱc��2���5^V��_W;`�MB�8p[$�T񀺄UTv�m�4�h�J�z� HP3�{/ma�"��V��K��͡���t��3�����,���[s�*�+d�N�q!��K��7�-�/lD��Mu�<���-�M���@�D-��Rn&��VH6`WVi���X)�[��uޞ�RU[�u�]ʭa�� �ɶsmz-�k�$�֖k�A�����7n+0��ZN-�m�!{�qj�;B�^t�p�[: 8lj鲳�w���/9�U@���4HN�\
bי6 i�@��6ۀ   7kmŚ.�!%�;<fW n��¬׭�-6�`V�M�nK�ٯ�l�@[�m��m%�0�Vu�nH�88��E�[@��`��l��8-�hm� �g5�m� n���m�>�v�N�C������]x�b�h�� E-� m��O@-�5��M^ �m�vͶĄ�P$' .4��yg�*œ��n��y���q[m�l���
��78�*��U�+�ÀHh���lմ��(s��-���mlp��[xm�i� ���  $  �-Hm����H &�Lvݰ  p i[mf�V�   m& �m� 	- �t��ں��Vyj����m5�mju�U�8�&�[�    $-�	   �I���$  sZm����u��[�� $�������l֪��t�n�l�$� :G6\��f�t� ��6� [@lm�eZ�^��ꪕ`*�"Y@�e��c�$�$6Ͱ $ l  	g�}��|��[�-�  8�כl86���@ Sl�-�햁��$� $ �����^��I��%� -�$��%���}��-�� I����`��9mq  �` �6��hi��2ԫA�t�vZ��U���V��hY� Z� itہ�iW�/u�����m"�dƜ��n�]f6��m�� 6�   �v��7mx���T8�%�i��&�H -�  qm���l=#j݀��R�!���	�� Rښ����U��'���y�e���kՍ�L�   vܷ���M�㵬�vͶ9Mn����UWKU/2��x6؀��P-�m��:X� �K�  �&@�}l�|H          ��IÍ�]����j
�檪�]�U�M�L6�z�$ݶp:�ʨ
�U���, R�\]��m��ڶ� u���m ��m�X�R���S�����m��`fL� �$
�A���UҬpUmu�Wd��x'����c��v�[�"]��V.0����Kh/D�sm�%�6���m�  
�u;7Sj�0�lm i$�il��  ����MΆX*�])rk����9�ZU-;e��& �nڝz�
�����Y��-4�����Rʑ���=uˢ��8sJ��  sj���y�, � 7mm�\ @	6ؐ�6��&֛` ��n�!jۀ  p$l-�Jٷ- �   {�� m�k5�i�in� [@�u�Im�3u�m i�'8ͶH k���6�m�kn		  �v�I� pm� $Ci��n�o�||pXք��k���m�6ٶ�    	m k��4:�&�HE���$m��<$�o  [@�	$ �e�j�N��V�m��@�� m۵(-�֚���ԺyA�4�fl5��T �9�
����V�6��v��j%��6� d�ݻd���m� �� #e��9�W8t�)�b�,�P�(m[[n�\�"[B�����093%̰m�R�r��S�UVQ��L���ὲ���j��#�����㝪��Һ�v�UV��ڪ�Βmֹm6i[����a��ye`.����aZ�K�")��qJ�b��آ���uN�ل	n��v&F�d�-�� kYmHV�Eq� �l�l   �uͮ�s��   ��	��b�l�C��o�Sl�	m��@   �  �M�9���K.�5�4_[:nV����� -�m��	  �A�� ִ���vI � [A����m  ˓m�vě`���ۇ 8m��m� � �  '��m�$m[d�� m�m r���!��,��g[@�m� m�!��H[Kh�M�t鄽(m6��I��ަ�-n�R�ZV�@9��M��n�v��d��bE�d�J���UA[-�b�j�"�PlYV�5�É 9Ͷ��pm��l$���av�8	e��ݶ �G3Kl  ��� H6��W�'�m�[B@mmÖ� [K�� �m��cm�6��- rO -�@8      � ���  h� �� �l���� �`��� ڐhl 	h���h� l i����l� I��kZֵ�3�QAPU4*���C�T Ћ�t"(/�����TqA�ł+�V"8*&�"1((b�?�"A�Qچ���� 0�T����`8_��ڀ!�UC��� `(uT_�P��� �@X
���N 4�	E�j@��tO�!���A1>B�U?������a""$`�H$ $���` ĉ�@� !��d$ 1�=E� ? �Q����*mD?	�'�+�J���\@�� ��AC�U���z�E�%b� �4 ��k�G��кjuT"
b�t_��B/�Z	 �u�
�@~C��=E� )T��E��)��"�*���pQW�>H����a�I �I��`��*�vMN�6�tݳ�L�09rsBm����F{͵Bܘ�y@����ק���v�I�=V�UcPs��:4OI��D9p�C=� jm��HKi���:+X.�J�L]�<�͐3=w��+!��۲�R���L�AFd{r�hM��ɳ��we��&���/k���g���JR�T�<�)F��.#�m�q=3�g��.�5�C�h�vYntݮ�MJ��X��\� ���kA�
�ut1s�Z^Dôv���!��V�KC�;A�u��i������70Z��'VUH��W���V̖뉻:p��ڛ�����gb�q㊫Nt�͖����E�t$�kUA�Pr�0q���4^�I[��iv;rEv���O�X�8�y����P%�A1�,��s5)�fE�]f�n�&ShLe�Lp�5lM��y�ts6�5�m�D�Waűlp�@N��9n-����3UIv��<s��N����:�2�"�[r�c/�O*��A+s*��vvƱ�a��ݖN{70�m��$��gE+n��WoFʧR��냊�`構/,m�a���KR� )i�`%Aȅ���mT�g(��鞶8ݧ���S�2��-�BW��,s�:������ Tu)ib�ڱ�iKrc,�v�-���[-sOff�-E��7,[���� �f�BX��Z1hC3�F�uGOVԻaԌ1y�3o3WL�P�p6����˞7��;�[F���ZP6�5�q�I�6���-�nlqJǴ+�-!v�� ��m�Hls6mp6�]q�c�8�-�PPccV�� ��bQ0��K�3%W$&8�wN�u7nz`����g����w�($ͳ�avj�5���n��tpm*t�&�x��aƂ�'D�Ę4���pҵ\�W9����k��L *�&u���e-�)��d,�z�����i� ƶ�[&�4�R��@J��r���a�x�mkp��ww{�{�_�	�Tj�� A 
 ���*b�~��X��k�0��@��j��Sj�v�(`o	�ș���6�c��b�7���v��R(u֝���l
m v�R�+c
s�&6L�l�i�݈xG���i��
�k��6⋢O[`;bQX:]͂Znv��[
�v�/;�I�d���$�\\��< ؑ,p��Q�l\F��ԝm��WN|k�V�W����tf6 r�-�K�.�3@�b��EԖ� a�kbD��XE[YX%���Ԉ�@�1KRѡ�E�������w^�u�W�W9ʪ��>X����v���][n��=�pϫ��)#��� �|��nT�9V�,�ҡ]	�0��X|�X}���wm������|WBN��{�m� ��� �ŀE5�Rn�S�e&�`��0��0��xu�X�xJ��-�[,�e����`XRa@n�=m��Ұ�f�L�Q���Dj8YX�;���t��� ��� ;헀w^ŀw�b�6=�B�]YN���$���u� �"DV ʪ�r�UU��Ur���,|�,��V�"SV�7cM	���ױ`�ذ��0��x�����>4Z.�wv���Xwn�l���,tq���X�;�n���ۆ w�/  �ŀo�]65mڰ9�v�,�c��9�HZ# �ˮ�����]�H�3�k-e�'�?��|��,�{�ۆ�����ն�/�wxu�X|�,�� �^)Mb���i-����w�p�N~�����`�"@V$X$�`�(9���rO߳���~��ԥ4�vR�]]ـwv����;�b�;�`�$�]��Lwf w�/  ���ۆ��SL�M�����5k�b���?N�kc`g#��N�=��
փ\�ۖȘww}�ϖ�r,�� ��x�����>�i;�X�Ȱ��0�%�ױ`��(�]Ҵ�;�Jݬ�� ��xu�X�Ȱ�m'*ڤ;��J�6��l��w^��I���n�ڟ����@DJ���P<�����7$罬��d��je|/�wxu�X�Ȱ�ڋ =�> ~��Oɮ��4��ҍn�����DF��hb��#bvz5G'\eӺ�\2M���I�X�Ȱ�ڋ =�/ �ŀj7iJmջHtݬ����l��w�b�<�G�l{���e�Ք�լ ��x|�,�dxwn5�E���7cM	����ذ-��ݸ� {d��c�.����]���`[#�>�W9�1|�I?w����?v�I��
4��F�m �"ȩ�������!�t������>��T�&����Zc&���HE��ͨr��: 4n���7UA�Aj�!V�ـ�ؔ�����2��M���.���R�j���L�ܺy�;�5q�.Z�7R��@��Y�Yq��n�n�{=ld��
��F�,ҍ%#Mڋ$��p�f�x� vgu�6��4�]�q R�m���#����YM��YJ���h�B�@z�t���m�,��J�[/e�ή�#=���h��h��&Knm"�#w	�$���c����Zփ����m����� =�^�=� ����D��q]�T��m�X����X����ڋ �[%&��v4�_����X���ݵ zIx[�Q�6��N�����j�պG��^�=� �=��6�]�t
ݼ�t� =$��{�dxf�Q��n���,hZ'=s���kt��ǒ�н<Ԟ���)i'N�B�%��ul����;V[�I/ �ŀj�պG�EJRb/���Bn��Iϳ�n�1�hD?  b��-��i zIxV�J]5O��
Չ���5l� ��#�M��w�b�;�[cl�wJ�V�xV� zl��{��<�ډe���+�l��M��~�s�s��"߾x��^��R�N��ucWamV�&�/5�*=��cV���V52������2�6wt�(�����X�H���� ��x[�Q�6��N�����j�>�9�r���>� ߧ׀w�b�:�m)M��j�
��x��^ zl��� *(~U��ٮ��?_��n^�"5wcWWVS��e�����X[#�����SLe������=� �dx��^�v��qZ�,�ae5�n'Xd2gnG�͵�����p�b+Ș��x�N}����;�X[#����G�w�b�="�8��+�E��m�����G�w�b�"�}\�UU$ylG�Ye��	��w�|��<�{�����Il�����4�.������� �O�x��^\��s�����:��ݽ�x{�NE�hX��.������ ���{�?�ٿZ��n�v�ccl��N��Id���4����e�3���h���h��
�V��wIx��x|�,�v<���Un�ۺe:v���ݗ�s�\�G�ϖ�'� �݉�@��i���4Н���{ջջ�:�c�<�:R�|.�+,N���� �݉�^�����ح�1:wV[�Wwo ;��^�����/lx|=)6�t�&'u|���s�];�r�)GT+sW�b�i�	����mt˩�^ֺ��@����^�x����ʇ2�*�fm�Z0hJō^X�m��T3me;, <���9֩Te��*���=j��e��"�^^K�J��g��*���k�|ٔ.	s=-ƣўۉpj��0���v�v�1F�M��юB�	�a4�ʠ�A���:Fw=�N�<|�n��L�K�
��h�nRw��͋��Jz:�7\��b��ڢ��H�&�^�|���x��x�د �m����4�.�;x�l��v< ��/ �������[���{ wt���U%�>���}x��B��]ڥI]"��������}��kذƫiT��n���Yw�ul� ��ʮ/l���>X��/ ٩"2���t�f��W	V"��+��PB娴��H5�W�puڒ�'
���&Z���}��kذ}��ղ<�c�.k7-Dr��}�_?I�,�	�E��A�L������^��nI>��u�n�m8��e�Yn�+�X���ղ<��<��,�ډWiڥWE�/�;w�ul� �� ��� 7v;�$�dC)4�+|W@����<��, ��� ���*���r�_~���{���5ep�u�� ^�lO����.j{Pf�ö�ˋ�	s��r���ϖ n�w�ul� �� 4=�)MUݪT�����5n�y�G���yo�<��,���Uv��"��k7$����䜿w���|�ȇ�x��#�p�ASAJ���#	��]9���a�`FX�t�Z��.h��B,�12Ɩ�LeJ34��ġ �"�[��j�`f0�(.�$A	��AP�'��@�	��x����	C����rO��q�H(��;
v�hn�������[�:�G�z8�˦�����+���ynǀn������'���7$����O���3DӬ���v��ñ�����aU�u]Ŷ�hI\ާ۱jy%GlLj��.�ջ��$s�xV��/H�-���j%]�i�t����xV���$j߾x��<wnZϒ>���I�j�(������� �ۖ��H�^�)M���0�Sn��� �ۖ��H���P�J	3;�ܒ��e�&Me��7v�ײ���`^���5��������"mD��2d��n�m��("�x�R��Ӌ����c}���x��[�E>'wk�yl��^��[���e�)M��մ����yzG�ynǀn�q�[#�;t��L)�IYb��x��x��ղ<��<v[i�&5n�wV�ݼu� �������D��� ����hN�ղ<�dx��x�Ur��a`�b��]X��A�lE��&Ѻ�u���f�s����;1�v���Z��h�'F��9�T:1h�����Gɫd��Mie�"�T4ل��z�ݣ&g�,��u���9�`7&���4UyI�gv�/nhي֍6��س����{��K9��m�p�8�ڭ~��go����RQ6+�������f��e�]� *���f��-�Y�,���>��YTA�Ve��F:�(¸��Okb�Q�,���\��̷hMRiڴ�.�;~W���<�c�7M�`[#�<�X�6&����M�x��xղ<��< ���F�j�W@�����0���[#�<�c�;��PN����)���:�G�ul� �ݏ �z��"�Q$�+b-$��ݼ��<�v<u� ���	K.�M�tuKX�ƌ�e���G!SC`C�[.�aѬV��!����q6%u��Wx�����׮<�d�\�-��I����n�v[��j���7^���Up:�G�uzG�ynǟRG��}V]�(.���ݼ�}��:�#��W+�j��H����	�MYvĨ���^��[���e��dx�k����[)�o �ݏ �r[�:�G�j���x?�������V��֫@cl��wM���Ǉj�\��[��Gn��vtʊW@����KxV��^��[���VҨ'n���S���:�G�yl� �ݏ �$��"�A)�J��hn���<�v</Ӝ����W/��*��d��5nǀz=lpJ�-]
����<�c�7I2����[#�7\m��tӲ�]�V���I��}��s�}����<�v< ��sC&&.�1���.u7
jPˮd� ��6�sy�	Vc��]j����Mwu�ul� ����`�"Hv��IQt	��:�G�ynǀ{Y#�:�G�un�F4�.�E��v�-��k$xV��-��o�
0e�TR�wo ��G�ul� �����<��PWwbv:E�o ���dx��x��ݷ�y�v�vԭt�Q234L͒f)��|��f�R*B��26�gE�h��j��(+�ZI���}-��ynǀ{eư���lpJ�-]
�R��x��x�\k ����<tq�N�컫�j���=�c0����#�<�c�:��"�]�J�E��0����#�<�c�=�c0�$�LV[�N���<�v<�&3 ���\�T��-�۴�ڱ���X��;34��y��0\nz��XȓW���1C��e3���F��} ��8Sp/l�7:%�&j�K��lVĤ��hҫ����`�<�_;��3iru��"�Pr���4���TaA����u&��(BM�UYLe�h��1c��z�.�);��mGJ컃�G����7id�ٛ��
�q�;F�`�%�`�d��wwH�g�����4��(b�Ф�����P��t�k��'<�ڵ�7 36e�3Qr�6+���s�Ol���dx�H��څ2ݪ)]���{dYXV��^��[���h�v)������G���'� �_}��E �!�[i6�wv�>Z��<T�<�Re`|���<Wѡ�%O��
Պ���[����`[#�<�G�lз��	����77%\^��
[�a,���ؖ`D[,b�=���}��|��b��V��@���0���[#������R/�v������Eջ0���rU��0a+����oٹ'�����r,|�J�)�Wm"��N��<�v<۶��:�G�j�b�iݱ2�e6��[��ױ��dx��x[�B���)]���{^������`[���h~xh��n�p���' �cE�{p]�^ҷv���+^�]285�nl�j��dx��X��x��o �AA&�|n��M���=�"��r��H�'� �����dx�R�*|.�V�N����r7�����W������_�;���-�E6�������:�G�j� �ݏ �����wV	]&���m`[#�5zG�ynǀ{eư/j��t6˫i]N.�n(���ݞֹ �����<J����lW�m
��v؊.�;x�H�-��l��ջ��b�iݱ2�e6��[���q��v<W�x[���W`
�ݼ�.5�unǀj� �ݏ �kD�+N���N��� �ݏ ��ջ�+���, Ab��(P $����1A4L�VY��Ru�x�q;��rp�D.k��-�x�H����l���v< ��P�y�s���f���s� �E�����;���4�$ƥz�u{	�V"�]��v<�&3 �ݏ��s�"߾x���ciݡ��5n���1�V��^��[��^�һ�ut"�5t]ݳ ����<�v<�&3 Ꚓ�q�b(����#�<�c�=�c0���/k�˻ce�m��:�c�=��XV�x��{��i��ڲ�D"FA���U�BI0#1H�d��cL�>�XÀ�E��j��H��J4h��\apaR##F1�R!	�9���qM���
4�5,�
(�q �a$$"��
H0�%ĕ�2I(HUXljJ����)*�R,# F$�*� J�B2*�-W�.�ЄBSZ6����EW� H��A�9�M�Ɩ�
P��(D኎�>�BH!��"B V�b�#�d#((��JP`Z�|���A�ER/�J��xE���#�cB�rB%+P�#HF�+)m
R���7ςX%-�
K�,�H`B���� ��Z�0JE"��
�� �!��X�n?`0��a��e�da#�"�B�m�$P�Qa���$R��bFĀl��N'���� 
�1�eUTe5�r͗Y6������[h�+����.�Ԩ���T�m<�Qu``��bm�e�����bqZ����vFPZgfV�5-�Q�3�ܝ���S��x��ۣ]4�n��]�Kr�֕�A �4�,I3F��GA��b��Q��#�-ĭ&��f�25@t�  ��m��Q�Z+�Ŷ���"Fy��Ψ�`0�b��&�X��L!�D��q�tn�U�p���vA�hM6n l���ZP�"Ę��͇m��E#lq���kn�K���5n9:�r���[���e��uX�۾@�������qi���t9m6�쉗-^�zd\d�vN��U��U&vٲXRddۢ���uRp� N�����:�RZ�:�l�[:��>���6{CV2t/S��՝$�ˡ�h*K��viJ
�&����P!c�2�uI��bUl����<t��$�+�UR(T�II�`�rti+�ֻ*U]3�-���w��+���d�S�`�5�4�ʓ����C�)e}sj���+n���tP\�xŜ�z36ȸ*N:v�"�ZE1�/"�UJ����v�5�+X�8y�]cc;�#D��\t�������|��|)CUڌ®�QJ$�A��6��wg��\��jn��jӋB�p��8نn���� 4�n���Z����1�	v��l�c�5>v�	܁��'�D��M���:���{bN:�-�B�����N�cSJ+��Y"���Y�
�I�����b�R2B�v���!6�YUW�kZ`���e8]��![Q�[��瘴���v�=Y��8�kPgv�Y�z��AeE�s1��5貨ֻUR��؛�e�ړ�%�eٚԛFӒ�D�	����@�-ϔ���`9v�E��g�'�]-��i���Wv���T]<�n�+�U�J��D���8[���(͕�m�cq��	ӻ�wN;J TDq �/��G`}���]0���l5���+G@�0p��i@��񰰄�îX��5)ZL栅0�ly4n7S3 �+f��6�VU`�X\u���A��jԲ贯3�K3�a.њ�k4 �Fe��Ƶ�l�g	S�1���9�Wv�7�K�ڣq�@�SF%r]�,�fS1[Xv�"�5�� W�8�ﭛ	��<���<�Ǒ�mʤ���c��!�w��xN�6�3M���<��'E����OtFr�џ]y�<�ܦ��o��<���02���޿�p���^��[���h�*��T�Z�:�c��W+�Ĉ��<�O�햢�.9QJ.�N�6�v�� )�8��}���Ey󏇰��|�����n��M.56�݀.���Ԓ��D�$�^�}�Idw� �����ma�h����y��NĒ�ݏ�I!zGx�K�v>�$�ڈ�.�;N�r�g<u���>#��˄�[�z��]UF�q�=�����d�K!�$��c�RH^��$��ݏ�I-�1��Ǘ�D�����KG>xO�㼪�)`�]{���%6f4�$�^�}��uԊ�y�}��l��\n�̟>�$�LX�I%׻z�G���$��V�)�v�����RKd3Iu��ޤ��"�I%ݽ��I/&�@A�ĵ�����}������ݏ�I-��I%=�uWn��z(9����^{��u�v1l�Ci�.�l`��&��ʸ*��>x<��v�.�$�C01$�^�}�I
F�r��t��v�� ���< ����n$��ݏ�I!zGy�9UU��Sh����*�1�����v� x��<=��W9\9Ƙ���$�v�.�$��,���ۙ[���^����>|���� <�{�� �_u����� ��!��p��KG>xO} rI�����>~�`�����VRs�ƚ�F[��vX�ɚ�[^悗�� �L�<δ��j����]I���ݍ˛�� ��w�ޤ��1�Iu���s��I~��$�9xr_��l[M-��� =㸏u�m��'ϽI#_�+Ē]��w�Uq��5�I���In���� ~yϟ< ���_s��I��IO���ĒQʊP��WP\�� �D}��v ~���|���k�svމ� �UM}�߾s�_< �?1�J	Yu�v��I.�r�I}��|�Τ�����RH��������H�K�n1nщ�u��iB���&�(5��F�2��U����GCx�Xm��b����}�;o`��q������@��w�����l�ٛE����?���?���EK����n���RJK��$������b�>@��z�G���$�}��$��������tA�-�6+��	wې�RJK��$�����$/H� ��}��Y�-���k����{K��z�G���$�}��$��\^���,�˹��(�D:�7��^;��f���nK�n�j�z4�+lS�v��� \��M���KI-&R�:h"7�5�)��Y��'<(���W��0�4e�d.2�\b+ӛջV�G�4l��uѻ &�[�9cm+)1`�f���������'V�N�p�DϣNR���ïWq�;�JM��;?�}�I�+kEt���8�k[�6�6�s��t�M;��,��^�d=U�mC7Ľ6,r��Q���ͷ#�4���k��,;a��;qL�I%���RH�^$��!���=�����{ >y>>��j��\�� G����r����K�3�I/���3Iu��< �xǚPH:ˮ��7`}��$���K��z�G���$�Lra�-�v���<{�`����ޤ���$��!ޤ�҅�^]l5��� x���� �s=���!ޤ��L��$�B��uv�5���v��Ly�)ˀ�NF��*�������\�#5�"�f�WKM�< =y��$�}��$�je<I%�폽I#�t�v4[.lg������N����]�q���$����ԒZ䷟r��6�Ns��Dnض�Z;x���q������$��oIwױw�%�ւ�3k���������g��y��v��*9�{y���o����������.s���`���<��ǔ�$�_�>�$�!���T�wE+���ud9lL�Q�:���{6�mҙ-�B�P���Tji��iF��ۆ��=�~���Ē�ǔ�$�_�>�$����$���J̺[F#�<��x���=�>�$�߾�Ē]��]�Im(Z#���An�.�`��x�� ~�6�%s�Y�So����I/Io)bI.�JT����]-6|� ?s�v y�{�� 9�g�v�u��oy����>�u�!E��ww�$��ػԒ���bI.�l|� =�6� <���mJך�`�J��u������9�5�#�؍���1Y���R�����V��KGc� 9��ܽ�?l}�I%�]�I.��.�$���U�f�j�
�/`��x�� {�m�o�{!&V�J]�'i��nݼ ��x|�,tٕ�u{c�	�t�И��E�+���;�`�V䜿~�nN� P ��Q3?k%��F7)U��wM;�X�+ ��ǀ�/ �ŀ}�s���������ӓ]�j��`X�jݰ���X3�0;j��A�;=2݁��Z��Ϟ {�^�=� ����JT��lo��+�����w�b�7v<����ۤ�&U��E�m���ذݏ+��������߾� ��Dc㻴�:�����`^��ޒ���XTZ
�'WeX�u�u{c�zK�;�`�3f�X�D����d��l�ˣS'.z�V�u�I�Ϝ�f�ۜ�I�# �cE�&��۠�"6�&6�����I�&,p{.I�793�׃�t[e�d?��6~�ԡ��w7l1V���;p������]v�� x��7n�M큭��B�"�8�;#��3%�OP9��]cfČ��/i�N�V��:�.z&���N�o:�n[��Yn���uζ8
w4�v�+sP�/y�՞Z��������5������J��^�(M��Y���&`J�����;V[I�v�l����X�Ǖ�u{c�	�ӗCt�Յ�+���;�`�<��� o��|���+�H�N���#��:����K�;�`��;n�I����n� ��ǀ�/ �ŀn���JT�∺k��+���/ �ŀM���lx��UW6]C�]��"��.�
\�p��f�9J�l���[J<��u�Cu�D�l�@���v���ן,wc��:����%�n�`�v�W@���=�Vm|���>r��,�3���^�=� �AB��n�U��]`^��ޒ���X�b��"�)B���Ym&����K�;�`��+ ��ǀ��:��L��'ww�w�b�=*L��� {d�dt0t�5e�+�e���#7[+R�+ZJ�#s]��O]��9.-#�K�U���n��=��+ ��ǀ�/�ru�S����}{��g�Z��Ы�[��� wd��ۆ�2��JTۥMp�v��%���0��P_�	�?~V#� �	�M���mGLx�4*v8�]�(�!4,�1KFP�R	"B��Z�ĊD� ��L�F,0�� F$$��BA���&+�08�ݡ���A8�1�	�O�4ԊFD4(;8"��#�� ��]��UD1*�A8 ��LTTi��t�����\�Vq.�7+ �$x�n���I�E�wx���E��uzG��/ +wP�
v� �	]ـzlYXW�x�Ix����Q8��@��tuƐ���؜�6�V��"� ����+�\U�q��s�
���%
f��>_���}%���0M�+ �`�"պ�t�۷����w�p�=+fV�� ;5�u)��+�Չ�����0Jٕ�u{c����o�m�j��HwM7v`��+ ��ǀ�/��?=�`��r�VZ(L�5M�`^��}%���0Jٕ�z~����\a�����M����&C�5Z�K+x��f.�Txh��<j2ʹ��5�[x����n�l��:�����%)3��E�wx}�Ҷe`^��}%�n�aNݠ�Wv`��+ ��ǀ�/ ��uj�(�1;���T�wu���Ϟ M���;�`�L�-��J��ڷb�7n� {�^�{f|t�|����w7$p��R�T�(�TB@k(4��w��f���u���Й	�na��lk���e:�+N:;15#�Ȭ�-�Em�[&��6-�a��훝��x�X�z��;Nv�C'�բ��Q���ۓocg��YUx;j]��
�*KJ�m�6s�K�rr�)��ٻ`��2�)��r�d: [H�N��j��N�6q[�c����t�9;<�Mյv��&|��&y�:4P�P�r�Oz�I$z�ڀƫ��n�8�g��I�$ƛp�nܼ�v���u���QvѮ���l���W�>�}0M�+ ��ǀ���o���m]۶�N����b��:���}%���0�DԻ;
-�6���lx�Ix}��b��:�)So�r��]�x�Ix}��b��:���ݴ)M���2��&���n�ŕ�u{c��K�5z�}�j����ޡ1��pt�]�z�Bg�(�ۗ[�<�d�K�HL�Ե��@.�U<�b��:���}%���0�Z��%6)!��4�����=�?�$����=B�}xϯ� �ز����*�Sm[��ջx�Ix��,�b��:�#�H�:�i�]��'ww�)n�,M�+ ;��;�x�+cQ�vՠn�n���e`^��^���ذ�j-��
qU������k�λAZ��{*w3���5�r��.�T��'m��WXW�xV��y�X��+ 4�5���$�]�xV��y�X��+ �� ��B�؆[E�I�x��,�E���E� �"�A ־���ܒ}ݗ���JQNݠ�'v�IV�� wd��{իP�
�
�Xj� �� ;�^�=� �=������B���6fG\e�.�ɺ��/a�*5]ƍjB�
*EaFj���ΛwwH�nݼ 祿�{�e`^���t�N�]�V'ww�{�b�=6,���< 祿}��˻j�7t7wk �ز��H������X�*]�:�	�cm���� w�^�=�*�Us�^�,���@���K��+���/ �ŀzH���lx��*����WF�Rx�o�ծ���C�Z�%[���"S�NG�gk��M�3[.�n�~}�ݷ��e`^���%�n�$J)۴t	ݬ�E��u{c�엀w�b�:�j��2�T��u�u{c�엀w�b�=$YX[QR�j��t�����엀w^ŀzH�����dhu8>5vX�ݼ��,�b��:�c�:�#�*���ʣ�s�:I����w���B;?�i�'mk�0T��4�9��[u	+�W�mҜ�h�qr�ٝ�Ъ̩u�u2N�tɘl���tDN�����1G�����`BQ[1�q]uʥ=�U<B1<)�+he��][P�U;.�<o��#��{@��(ܽ�6&L�ybMG:q;���y�f�'7&^]*��Y�����=�R)��1�,�H=�evA�L���t��o-���hh�c��9u���\MQ���rd[,q�h��g������-Нݯ߾�e`[��^��ױ`��v�;
V��WXV�y���UI[�� �s�zlYXT"�%�����o ��  �ز����n����+�Qt�n��{�e`[��}%��hU(e�T����e`[��}%�ױ`z��R%�ۻ�ҥWe��'un���X"�Y5�5{
�8�/�}����GK$X�Vʥ`;W]�O� w�^�{�e`mD�I���"�v�����s��*��!kذM�+ �ݏ &��S��hj�����ذM�+ �ݏ ;�/ ���Ҕ�ݖ���;�X�ŕ�unǀ���w^ŀ�R�ګwJ�ձ���ջ����@�s�zlYX�K����!r�vyx����9U��E�Ӡ.n��k�J9��C&�]Ѯ=��g ��  ��e`[���t���Ҵ2��I�xwn��+ �ݏ ;�^ {v�R�[�@+�Wv`�,��v<*�\��s����~�� ���uj�H���]3���WXV�xݒ���0>�qo�|�X�|R��ڶ��t�M����/ ��� ��e`[����eИ�t+��ᙅ�l՛d�!1ҩ�ݰ�ٌ�А������gv�Չ���I��+ ��ǀul� �1)J��t���7v`�,���<�|�)�� ��Ќ�]���5lm5u�u{c�:�� ��l�e`P��9uV��Wo����<�/� �"��)A��@��)�\���<��MJLM"�]ZI��;�`UO��]�g� �$x�F��̥gSӁ�XC�����&���J��L�@tõV�P��&sa��VT���e`^��Sc��Π����<�JH�t�.��`YwXW�<��~��6E���l���L�-�*�m[MۺC����I/ ���ʪ���e`[>x&�r�Lm[�ww��� _�w~��w�}�rN_�w7'�����&��%�+weҦ��ـl��XW�< ٲ��n�T>$�U�	bl,X�m?tҁ��aC��J1�D%�H&���`�N0�8	�B�&�B�!$���$.��0�]~�Q�8�F�"H{�G�mJ0c#,)
TKE��ڿ"|���!�!�A�t1"c0H`�F1>LMBRU �	� �D�H@9$�8��`�"B0L��N:F�_̀q�b⨽a!���!d��U���sY�sZ����L�� $6��vni��Ҝ��nr୚���v㍊�N}5�Vѭ��=�`YBj@啚�����kh�uۜrXi��(����JsɸR���r_,ד�bY&iKwL��B�kx�#Z�ax�@qc�ں��D���8T�'mK� %��4F	�[h2��St=X�b6-�ɷ;%�ۓhi�:iR����#H٢"&,�]P�k�c�㴃�����ڝaS�ٴ�<�!R�\C�ې�-�ĥ�ڹ^��i��6���l\n7:ci�t#ٷ%���Q�K���m��`^e�l����ѱ�]���
Vw5�P��]���T���0�g�qe��RqU$\�F���P�F����nq�St�Z�8,�0E>#q;�I�WI��J%Y�Ga��f�p��r49�G;�:���bC�$͞�t�sk�n���Ft7/,]�Sx�6�r��k��ȓQ����y%xW�T`���D�v��΀��'3�t����^���V$�K%6ښ���n�v8�m��H#�m=�N56m[6�padl�� �F��$�%�Q��ѣ�d� �c���b�F�m�,����S�y�\��Ku�m��N��c� ��A��H ���:��&�U��h�����t��l[s��ʱ�!\.X�d���˦��6Ν�aŷ$� �u�P�E�<�\�Gk�3���tSi�e����1Ҙ2s9�c��$�`hhT��$Į��[r�]���H���C)���b]��yUy%8�V�T{4:���B�(�[Tnc!Pn���d�+��h<�+.���Rj�gX0J����v��s�Ɓ�tk:l�FJ�l�.m\w���I�.�BYzT��3�0ܻʫ�+&ϵt�1�N��Ͳ�	���ڢ�*�I�/cj9��b
�K^��heG	ѭ`��.9y�*�K;q�&��^�\�EUU]uH �BvN�9j:�35&�L̚��^�F��B(���*��4	x��*Q��@��#�R��e�AqQa��01�õ�Ǯit[P�`]��k���]���;IK�N�+�ey!��)����\���ە��6S3Y�a�XT.�iyD��6Q�4nƔ���h%Rk�5x%Yk"tl���݅�a�r-6L��&���� ]��4�e�8��rı����h�nb
��3��؁밤��.�x�:0ucWm�P�kN�ɞ�q�]<�ԍ�knx�j��Gc�C`�f��dr��ogwI0y�\����V~-�< ��x|�/����u�|��/��R_,M���+��uM� �ŀlز��ly�s����%�_!��.�E؄���>X�V�� �< ��Jt�
�ݘW+�J}�˵�yl��RG��9�/lό�T���N���+˺�:���RG�w�p�6Be`��]���Hwm�q6�f�A�p�����s�hҗ*���Z�6�n�vB�\�,g�mۺC����~�����0�&V�� zk�,tҷ3WR�kZܓ�k�}ډ�|�͞�� �>���� �1)BlT��t6��eI��uzG��J/�����0t#%�nݠM[���H�Sc�;�`|��>�`_R���X��Wo �6<�ۆ��e`^�ǻo���yzY�����i�4.�e�y��\���G���ҩ͜����3m�ܑ��L��Bv���0��+ �ݏ�ʮ�������>��N�P��]ـl��XV�x���ݸ`^Z
���ؙ�`S�����lx]Up�<��"�@�"`��Q\�.��p�;�+ �aJ'hl�@�v�d��w�p�6T�XW�< ��JX�t�lV�M���m� �Re`^��d��l��I��?�=��z1��$l��-pL^�FLKu�3��r�jʎ�����ز��]����L��{ l���\0k`Էi�]	�i�N� ��ŀ$��s�rO�;ݛ�����=�L�fVh��WrI�{�ܓ�g{w<�����lܓuϖ�m�QSt��C�&����w$��{�rO��ݻ�|ԕG��������K}��fXV�|�+ ����/  ���UW��*}���\�-�M4Mi��[h��ogR�8p�7�Sʣ��J7:�	���%]�@ݗ��/  ���"�R�I�-�:�Wf {d���ʪ��M��� ����{n&�rƓ�+b�bwwx|�X�&Vr�ݗ�>��	��%(M��ڷCwv�M�+ ���uzG�����, ڟ}t��:�i�n� ���j��nIϳ���}ӽٹ&ת��� �t!�}���j�6��
�X��XKF9l.��Č���q��jR�q�Jm-pX� W[��nv�xr�ΜX��s��5����;:��͸[����n�)�ֳ�V	L�s��̣���km�.�s�C��m��e,ՏU�d3cn��Ȍ�	��j-��$��<ł�km�����
���ҙ�`'y ꡴�{j�睌�O"��b�Sm:��{�����M�[�@�h�:U4ʐ�BK�y�M��'ؼ��*ԃ�箣,����^k��W��w�E�zT�_s����G�lSF��U�v�?<���']Hߧ�e`��0[#���q �D/��.�ҡ]wk ߫ﲰ{nNq(�V|�XW�Z*m���������R��!�E>���`�&V
N��o�iـ�^�W9U�]~����=�`�$�)'�-]QV��+!;���V���"u�[iD�����:���)4R�+V'ww�w�E�zH��{o��T_��$�}����vg�[����v���ݬ�E��\�)#�ۆ�6>�~yÿ��u$}����9��dT���/� ���9�"��<=��y���^���{���Ru�>����� ��e`��`�]
Rct��C�Bv��\0�\�*}�˵�7e�`d��E�5�E�v]�m;�����XŬ��n[�;��9��G�Z��ݺ������
�ݘ͋+ ����/�Ur��=�_�� �l.�[\,j� ����/ �� �"�� ���?����������kW,�������a�UQ���9�U3fE��nˆ l����O�����v�>�W����'�|��{nT����MJ6[v]�ۻ0���Un���_}��;�"�=6�1���bۥ,R�l��a�K�b�0<�qp4L�q�fq�Sh�[m�iݷ��w/`uM� ����u��e`_R��ڵe$�]%n��ly���ďo��O��rO�����O�L��zh���3t����l��}!��{�p�͗�dcn�����ӻ��UT�����7e�`f���\9\��U�U5��-Z��n�,�� ��� ��U����o�^����'�,~{?n����M�<sr���]�j�,4!�5��3c��Y��\DU���l�z�f vl� 祿}!��9\��ݗ�O�?�j��lV�M�� w�^����=�`Sc��\�9_�\�l�?[i��6Ҵ컢��� �}���{n~�����< �����Ɣ��w��wm4�u���UŻ3� ��|����?W+�u����������sR[�e�O ��*�r���~�~�����=�`��K�>�}����m���U�gN��^S���.��`htR��#"���I���0��X�ۦ��j�#!��S�Ă�#]�&87���jA6^�$�kpԈ�Gg1ێ���.�k9+tW+Vw4]V���G�8���r57mrԏ]$��ٛ��[d�sv�m�j��m���
+����0e�3s��6�����8ϩ�mz�@`��M��	eZ6kW؛Rv���q)��hۮWK���h��SA��ҳ̥����}x�ee`��?r�Π��|����m��@+��wx�eeg��9UI��0/�� ;�/?W+�H��|6
ݠ�`����/� � w�^��YX[�WI����;0���}%�핕��r�Ż3� >���%WL-��!�v��Ȱ����=�`Sc�=������M�[)l[��c�C+�W�6��X��q	�,tr\���Kvg�uԙ�(���F:Q�[y�>���{�p�7�E�w�E�y{Rn*�wA�ֵ�-�F�}�]��5�E �L��o�rO�g}w$���l���_R���ڲ�eI[� ���`�ذ��r��ߧՕ�{e�`�.�M1��C�����{鲲��n�!� {�����O�{�.\�.i�]M��=6VV����lώ�5���;���~�-�/7Yfp&4�%�31�%�Q�ڙNA��v�I�&sMMw��W�S����Iӗ�0��[wN�`՗^g���7�E�w�b�=$2��D7lv�]�iـo��>�UUq#��� ���+ ��T#ht[��m��;�`��ݛ�]l��C( ����"1�1T��^	��Q A�AA$��P�1Fi�5SHLS
 bNm*H�����} ����SM� �"m話~ ����u� �{=-�Ԧ��]*�t'n����UR��˵�{e�`�"�;�`^ԛ����t[�6ں�;�`��U~�*��_L��x��� �Ȳ��K���$��[#v���<V�S�aAԥqZ����͔h�cp6���Lu�ݮ	� �9�=� �Ȳ��Ur����/� ����.�T;�i��;�`�X}�|�Y�W*�I)>����t	�X���V�m� �9�9��A��݊�Av��	���w~��w�{�rN}��w$ȯ�UR$���	�2!;v۱q�v���Ȱ�ȰM���{�p�?Ur��g���e��V�U�6K��/b�Y�\���jR�n���k��;�5���5�Ӵ�m���� ��X���H�	�m��5n�V����`�Y�9��F쿌��x|�,Vě��w��Ӵ1�� ��uIUW8��ϖ'�X��P���Ui����ف���r���|�k�,vC+�s����l���4�N�C�Bv���X�s�RO���=��0�"��t{�>�e��K\j�橸�&ӂ��t�`Ɓ�K��۴��WJS��U�Nwf0��.ò)�6�HU�k���\S�i�9B���g�S1&*�]���jBm6�%f8����tp.ҡ�Z��fMn���Xt킮�{8⢫`��ΐ6,>q��nT75$Ϣ3��('[9��v���j[�JL3ke2a�k[X�x�{KU��f�=��ă���OP��@{05<�wl��Ў�L2���Sg����x��6�.x
�6o������;�p�;� ��� ��6�6"�U$n��z\0�"�=�"�7vVV~�s��ܮs���~�۷w`R��;0��~X��X����=�p�	#]1�������s��/m���&ϫ+ ���v=� �ٍ��+wt*�t'wk �l����9\�ٟ�9��;�"�;4-����]���֝X՚7<����s��y�N�:�j��dU�uCp`\l;��8��v�߽ܽ�|�b�;�"�7�++ ꄥ��j��	��f���~��M�	�u�����VV�m� �m]D4�N�C�I]��r,}��������Kv_���,-�F:bw��'v�ݕ��{�p�;��Ur��{o�娔|:-;T�]���=�`���ϗ@���X�ee`��]���J�+�M@�"�Ws�y˼��i�P�cS��l��f����i�\�	QnO�{�{|�r,}�����*���7e�`�|}WE��؝�4ݬ�r,wee`��0�"Ϫ��T��O��իn�	5t'wk �}YX��;�r���E�w�E�j�qYn�T�E������-ٟ�s�w�E���UR�>�����/�]�-+aE�MـuM�  �l���ۆ�9ʩ.�!����Y`�)L,e�;j�.��������K�[��G�Ӻ�'��q���j��>��,}���{ncذ�Y��
�'v�ݕ��r�#v_���,�r,�\�W)#V����i������7e�`�E�w�E�n쬬 �D6�ݻ��iـv9ϳ���~������߄	 ȩ�I��yi�]�e�ڴ�n��9����{nT��KI�t>
u���NJ7\�֥��s\�1���]R��\�.�T����;c�o�����=�`RG�9\�����X[��Yn�!&��I���m� �<�r,weed�?Sf���m��n�/���[�������{���u)1�� ��9����{nW8����|���t�v
�X����=�`RG�w�E�>N���w���~�YJ�^C]C1�Վ�\E�̌un��ML���9��`�mq�q��]� ���Qv�����#��R�����;v,�<��מx�6�xH����\nu�s����P�nC9��s���<K�Gb���K3yZS��n-t]pFҧ@Z.�zYm��:�X,��i�������.8����t�j��	�*[����{��}ᧃ���_Crg��ܯ�$9n��8��ɴ)6IaV��gs��2��	�]tl���H��Ȱݕ��E�DCj�۰)Yv��T���`�++ ���Us���>����v�-&۷�{_�,weea��U\�%�/� ����mZ���CwBwv�?r����Wk ݗ�uI�9��QYnВmM'WX���H��Ȱݕ��j���{8l��`F3d��x�M�v|��*)�{:"H��!i���Nk�_�T��n�t/����`�++ ���{��q�Ze*� ���~�}�:Od�9M�O�+ ݗ�uI�5)S�+
N�`�++ ���uI�9�5� �Wc�������*��s�\r}������  �l��-�4ի�`Re�v`Sc�?s�U���Usf~���}���{n�߸ }�y��t��h�6ئ4m�*����"Qg�"^�<6f� u�s�3��&U����� ��YX���H�M��jն�����n쬬��Us���0/����`�Q[�R�Һbuu�{��uM���s+�9B��"�0�Q"��!�z��ܪ�s;-��������;�����+aE�V��:�� ��� ��YX�.��u��V�WHWo �����?�G�E}�I;��M�9{��~�����&R۵QH�4�WZ�i�c�+���c1B�ͥ����n�����p�������z\0�#��ʪ���|�֣�wM:��۫�ޗ�H�yȰݕ�����U$E"U�i��ݰ�uv����|�yȰ�\���}YX�������7v+V�m��=�"�7vVV�K� (@�?k��䟽�o32�:�����n쬬�ۆ vIx|�X}QJ�t�l-�*�V]�k�"]��,f\�a���p�u�ҍe�gg�8�@쫷i
��t�uu�{�p��/s��o�T哽�}���ڹ�][��Jݘ�%��`핕�{��=�t�Z~��3�k��\z�|u���7�++ ��� ;6^�4J��XRwk�r�����v��ٲ�?s��r����� �j3�L���N���uu�{�p�͗�w�E�~��M��!�؄1(n�~ ��ڛa4���`@��p)Qރ0��(H{��g渎�qq`B1)�"`ASj;�1��!
T@����J�+			`e16���(�@�)��)@�?8QN+�����~5�z�n� l�K��x�I8��×ճU]�ݧ`��W�h�¦Q��(����ez	�[[q��iF��7��Ŧֳ�Em�q&(��6�\<i@;���n��R�p��4�I��Wv�s6ַ]k�q�� ����kG�k� ��hR�݁S����g[.�k;sB�J�^\h��]�ؓ0V:z���NY��ݸ�e��ڰ@l	1�$�����\�nD#T]�N5��n; 4a�q�l��x2�j����õ�Û�\5[�&L6��,&���m׮�z���wk�z��\ڑ�d�WBP-�@���LZ
�b,-��!�V�(�i[=��P6�)�Fl�]�å2�UI���[n�9��
��N�;:�ٸ�%W��$������%�](qnm*E˙�u07k��v��O[8nM�{+����ۮ��4�a��gۮ]�]eB���cS��kt�A��t���-0��t�a�����H�ʘ��z�ۢ�9�v���R�]�m)iSn5݉�����w�x�M�I[�����	0�41���%�\C9�eԘ+i啧D@�k��E�L�Mj�U��4.2�n��E�٣7=q�m�wG	([���ŬY^v��� �b��:i��T:iNyN�\�k`���;=X��ƚ����Z�ն|"��uJ�1�Z����ӱM��keS+JYvq�ҁ�W1�U&v�R�v�cUh��*�Q�w\�=����u��C�L�]��v���,�&PUq�]�q���g�S��DlJF���n�j-��m�]�ChMMkp)F���I��$E����js]ŗ�
�*��Q�X�ʹΓ����� 5����6���*;-,K*����ŕGR��6����e�Il�*�7Rʵ�h��F�N���$UNH�ؗ�9���bGMѻKb����<خ*������Ţ�`�aX��U]uH 9b�pmV�P��-�U�:O��w�;�Ӕ���0���� �� �T�
���DL��;��kN+�ɶ	�5�EDL�4T�Ƭ6]�B�:bǙq�s��V0\>��E��i6�f{vPMv��q���<�a�<��K'�u���Of�y3;�a�nv��p!�Q�;���ˋ��w�FHm<u�wl�2s�DUF��e��mP�M��9=7][-�]@]��Ļ�#l����=sN�G9s�g�5	��Mw:�5�6��	pT>���{i�6��c9�ۯfUؓ�n�)��a�Յ�;�E�У�vUm���]����N΀{v^�9��Y_s��9UΠݗ�|��c�;hM���r,}���{nT����+��q#~�cm�Hl�����I>���ۆ�$x|�X����aA���3��N������O �����9�w�r �7���}�h��W|E�AE�V��:��  ��YX��iiT����t�&ڻzB騖��nٝ�^2untl"1�փ�A� ��$�7lӲ�]2�B�|�����n����=�~��9]@{ﾼ�������'v�ݕ��ʮ${�p�zK�;�"��UʮRG�j��r۫���]���7e�`d��w�E�n쬬 ��Tm;�Wv�iـ�^�9����>�*���f|`�*���U�I�Bn���Ȱݕ��{�p�͗�~�+�[>>C�Ӧ��i���1�n�\�X3)ZC!tF�M�l`�̸]bJ�O���/�m�u�b�H\��������{�p�͗�w�E�j�Ī�ڤ��t��� ����/  �����y�I�-?�����)Z-v���w�ܓ�g{w*��H�� 2*� 1#D�R�����f�������r%�bX����=��̵�W�WΟ��N����{�iȖ%�bw�|p�r%�bX��w~�ND�,�A �3������ҝ)ҝ?����j���o�>D�,K���ӑ,K������r%�bX��{��r%�bX�~׽v���N��g�����<�8�G�[v�a��GMvqh�-�.@&�n����Djy's<��&��E�,��6��bX�'��ߦӑ,KĿ{��ӑ,K������Kı;����Kı/��g�\�[�dG'�>)ҝ)��{�kiȖ%�b}�{�iȖ%�bw���iȖ%�b~�w���,K���o`Z��s�vWΟ��N���u�]�"X�%�����"X�(�ș����ӑ,KĿ������K�B�9�>�Tȵ
�e��S��/E�bw���iȖ%�b~���m9ı,O���m9İ>�D����ӑ,K��:Og���jRSR�ɘh�r%�bX��w~�ND�,K����ND�,K����ӑ,K��{�ӑ,K��d�̦{.�jh���7n�+�̙�C�1�V55�730HY��*��	nIq�*��1փ-ry��ҝ)���=�fӑ,K������Kı;����Kı?~��6��bX������U-p���t�t�Jqb}�^��r%�bX��|p�r%�bX��w~�ND�,K����ND�A{^��N����[����B\�Ο,K����p�r%�bX��w~�ND��"~��fӑ,K���]�"X�%���׶z�S\�Z�Fӑ,K������r%�bX�g���r%�bX�~׽v��bX�'w��y��ҝ)ҝ/����뙲�L��jm9ı,O���m9ı,?� ������>�bX�'���ӑ,K������r%�bX�q�0*D`�"��'m��f�`p֒����>�����(M��-`J�[��b�(��T�i` ��4��d�ջx��K�̶��i2e%�`&R[�U�i�u�&M42K.#ai��V+�$�<�ص���T��m�����������o-dri1�g<�v�Yj����K1�N�s�&f�2�\�i���R�����[-����Cŷk�7�J�:�s��>�T��nH�S�2��l�*��<����f2�+�0�����#Xz�gSl��ON��N�������r%�bX���6��bX�'��~�ND�,K��}�ND�,K���*�!���;�yz���^�=�ND�,K�{�M�"X�%��{�ͧ"X�%��u�]�"��2%�>�����%��Y�ўt�t�Jt�;�o�m9ı,O���m9ı,O��z�9ı,N��8m9ı����B��ᣭWd�å:S�����ND�,K��޻ND�,K��ND�,K�{�M�"X�t�O�x���Z�+)Wy��ҝ,K��޻ND�,K���ӑ,K������r%�bX�g���r%�N��}�?�l�J�r�T5�{hݳaa�=��<��^�6�6�Μ�tu�Y�Ip\�t�3R5���Kı;��8m9ı,O߻�M�"X�%��{�ͧ"X�%���{�iȖ%�b~3��=]f��5�4m9ı,O߻�M�!�	���K�o�ͧ"X�%���{�iȖ%�bw�|p�r%�bX�ݧ�۫G�2-��O�Jt�Jt���iȖ%�b}�]��r%�bX���6��bX�'߻�M�"X�%�}��o��PΦ�;Ο��N����]��r%�bX���6��bX�'߻�M�"X�%��{�ͧ"X�%���v�}F�lJ9�}O/P�B������iȖ%�b}����r%�bX�g���r%�bX�~�}v��bX�t���y����B+���u�'-����D[�Ұuδ�ݛ�y��l�4����j]3ND�,K��ߦӑ,K��=�fӑ,K������Kı;��8m9ı,O�׉}��3E��f�u��ND�,K��}�ND�,K���ӑ,K������Kı>���m9ı,N�����rf�u�K�˭fӑ,K������Kı;��8m9��G�2%���ߦӑ,K������r%�bS����[��3�*l�:|:S�:X����r%�bX�~��6��bX�'���6��bX�'ߵ�]�"X�%:}��?C�;F]5��å:S������iȖ%�b}��iȖ%�b}�]��r%�bX���siȖ%�gO�Z~�%�U�qs�d�c0���������IG��=d�W j͘9�����L�3�Mj��%�b~��fӑ,K������Kı;���ӑ,K���w��Kı/�O_I2��a3V��ֳiȖ%�b}�]��r�	"w���pI��u�$RD�wI��⢣�S"X����fe�2�2SZ�%�kWiȖ%�b{���ӑ,K������r%�bX�g���r%�bX�~׽v��bX�'���z\�֩,�5�&f���bY�(�C"w����r%�bX����ٴ�Kı>��z�9İ +�(!"��R)�a�"�H�Q�������"X�%����_W �.�e�O:|:S�:S�����iȖ%�b}�^��r%�bX���p�r%�bX��w~�ND�,K�	??��١���IX��4a�E��u�<m�8��RN��s��6�q�m�׾t��y�y.1�n�I��]k6�D�,K�u��v��bX�'w�6��bX�'��ߦӑ,K��=�fӑ,K��w�-�S5�Iu!��]�"X�%�����"X�%���w��Kı>�wٴ�Kı>��z�9 @�,K��=\՗�kY�iȖ%�b~���m9ı,O���m9ı,O�k޻ND�,K���ND�,K��vK�c0L�ry��ҝ)ҝ?����t�ı,O�k޻ND�,K���ND�,B������r%�bX�ާ���t3i���å:S�:}}��r%�bX���p�r%�bX��w~�ND�,K��}�ND�,K��~~��g\���1���Jx{!N<�v�\�뎌v��=�wl�m&)��k�X��c��tps;�0���H�0��
�Y�i���V�6ݐ��͕�<�Ʃ콬�8���<��r���'k�#�h�Jө;S�eJW9cE� \F� ���"�l�(�3l8qV��:3���R��B�s%�*,7%�շm��b-�M�V�����v5����{���� y{<�Ml�E�&��ϧ<�^��ƕnuݢ�7#X��TK�D5Ga����ս�%�b{����Kı>���m9ı,O���m ND�,K������N��N�ߚ{��*��0�3��Kı>���m9ı,O���m9ı,O�k޻ND�,K������N��N�޾��9.+-rm9ı,O���m9ı,O�k޻ND��
�DȞ￸m9ı,N����ND�,K����.L���d�Y,��m9ı,O�k޻ND�,K���ND�,K�{�M�"X�%��{�ͧ"X�%���L��.�k$%ԅ�j�9ı,N��m9ı,?� �}�M��,K�����ͧ"X�%��u�]�"X�%��;9���cUڛW3���TH�;i�E�םs�FYk�ؠ�v�=���xv��"X�%���ߦӑ,K��?{ٴ�Kı>���Kı?~�y��ҝ)ҝ/���/�j�����r%�bX�g��6���Wq�8�y*�RD�%��k��ND�,K����"X�%���ߦӑ?��&�1ҝ/��g���enXf�g;��Kı?{_��iȖ%�b}���ӑ,�"w����r%�bX����ͧ"X�%����e�d���f��%�f�ӑ,K�>�}�iȖ%�b~�w��Kı>��ٴ�Kı>���Kı;�Y�������Y5�&f��"X�%���ߦӑ,K��;�fӑ,K�����ӑ,K�����ӑ,K��~��e̖L���v3l�qbn98���c����v�oGE.�����=��j��.����<�,K��;�fӑ,K�����ӑ,K�����ӑ,K�����l���/P�N{���$]���\���bX�'�׽v��bX�'���6��bX�'��~�ND�,K��}�NDı,Og�e��u3Y!.�.kWiȖ%�b}���ӑ,K�����iȖ1a�J�d�	 �#P��
���H��L�A)B��`���(0(�Z
T0&q�F��X�t�#HF@e�0��:�G�a�i$`��) �d�� BB� ��*����
����b�� h�vUڛ�(���"FE�%-��H�Ԉ�!B$F�� V���J&|B֥�l����"|�4�$����%�<���aBRP�m�!s�qd�r����R&a�``a�J���	s��+
¬�jJ��.��X��lt�\� E����\�@�)T$�Ȍd�p�����@��xA�F0v@�"
��bJ8D�P��Q�� ���"� �,� �"A�#@6���1�LBUbT�F%%�����b�e ���E(E� Db!"J�@�Q|���&�?�P"�����n&���ٴ�Kı>��z�9ı,Oߦ�f��֭���h�r%�bX����m9ı,O���m9ı,O��z�9ıP�>�}�iȖ%�b_vå��]d̐�MMf�ӑ,K��;�fӑ,K�����ӑ,K�����"X�%���ߦӑ,K��Q=��m�Ϳh�m�FN&�u�v���;Do�Q<&j^7s�:I�t�[p���2�,0۳���҉bX������Kı>�}�iȖ%�b~�w��`)�L�bX�������t�Jt�O��|�o�.��El.V�9ı,O��p�r%�bX����m9ı,O���m9ı,O��z���ҝ)ҝ?~i�=�3IP��6��bX�'��~�ND�,K����ND�,K��޻ND�,K��m9ı,O��-��4Mk,�%�u����K�������iȖ%�b~����ӑ,KĽ�}��"X��?w���r%�bX��z۬ٚ���t�t�Jt�O�Ͼ��,K�D��}��"X�%���ߦӑ,K��=�fӑ,K��~�����M�[��M����bd�Gm&6��4�F�Q���F����V��B\�]�"X�%�{��[ND�,K��~�ND�,K��}�ND�,K�뾻ND�,K����z�ոIr[�k[ND�,K��~�N@D�,K��}�ND�,K�뾻ND�,K��}��"X�%�}�å�ՓFd�jjk56��bX�'���6��bX�'��}v��bX�%���[ND�,K��~�ND�,K�����E��h�5nff�iȖ%����u�]�"X�%�{���ӑ,K���ߦӑ,K��=�fӑ,K����33�.e�Y�j��WiȖ%�b^�ﵴ�Kİ�Dc�����}ı,O�����r%�bX�w]��r%�bX� `�B AG�)  E@�@C�;��F�XCHb�I�
�6�̖M��b�v����#�B�u{C�`^<�z�4Ѓ�����L"j���^ۂ�$A�u���d�g�8��!��u�9{u��(��\�st�׬)Χl��=�����d�lztx�nG�3�8�3N�z���Yt�Qƍ�Dї�-�����8/ZѪj$u�3�����'����Z�aC�N�����x�u]ps��H:ێ���C"�1�ZݤӰ��[mP���6�pܘe˕��Ȗ%�b~���6��bX�'���6��bX�'��}v �%�bX����y��ҝ)ҝ>�ޖ���Դ�evfӑ,K��=�fӑ,K����ӑ,KĽ��kiȖ%�b}��ǝ>)ҝ)������is2���Y��Kı>���Kı/w��r%�-�b}���iȖ%�b}���iȖ%�b{=�/�d��$�R3WiȖ%�b^���ӑ,K���ߦӑ,K��=�fӑ,K��\�g+�)�r�ʛ16j�'@����m9ı,O���m9ı,D���m9ı,O����9ı,K����r%�bX��'Ose�����-R�q�X��s�5��`<��b��̙��++W4�V�jL���å:S�����ND�,K�뾻ND�,K������&D�,O����ӑ,K�/��g���!Z�S[�]�O�Jt�'��}v�� 	  �TL L���%����r%�bX����m9ı,O���m9ı,O~���{�64´.V���ҝ)ҝ/{�kiȖ%�b}���iȖ?� C"dO�����ND�,K�����K�)�����2��Y���å8�QlO���m9ı,O���m9ı,O����9ı,K����r2�)ҝ>�����H�VWd��,K��=�fӑ,K����ӑ,KĽ�}��"X�%��{�M�'Jt�Jt����eR4�9ƗU(�ifZ����͗snn{E* ��,bF���m@o�'t����Z�mknw�>)ҝ)���}v��bX�'{��m9ı,O���l?��L�bX�����6��bS�:��ٯ�Y�6P�f���ҝ,K���6�����ș���o�m9ı,O�����ND�,K�뾻ND�b �"X��r��]M\$̓Z֦ӑ,K���o�m9ı,O���m9�S��4F�5�����Kı=�o�m9ı,K��O��Yef�ȎO:|:S�:S����6��bX�'��}v��bX�'w~�ND�,K��~�ND�,K��}�l֘͠��{�yz���^�����9ı,AG���ND�,K��~�ND�,K��}�ND�,K�{�>���5m�L�jkX\\�a�Gk\��;tp.
y��n�W�1���,��Z[��V��ߝ?���N�����O�,K���ߦӑ,K��=�fӑ,K����ӑ,K�����z�̶:�U<���N��N�߿y��?�	�2%��=���ND�,K�����Kı?w���r'��L:S��X���(����<���N�%��=���ND�,K�뾻ND�,K����iȖ%�b}���iȖ%:S����Uh��5�w�>)ş�T������r%�bX���6��bX�'���6��bX] @R1Cd�@�� *!�����ٴ�Kı=���3W5���B�j�9ı,O߻�M�"X�%��������%�bX����ٴ�Kı>���Kı)��ǅ#��+�;J4	uE�e�r�i�tV6ۖй?���O��Ӫ�u��.��.��Si�Kı?{���ND�,K���fӑ,K����ӑ,K������r%�bX�߬��E.���MMf�ӑ,K��?{ٴ�Kı>���Kı?~��6��bX�'���6��bX�%���d��s	�,չ�5�ND�,K�뾻ND�,K����iȖ?�r&D��o�m9ı,O�����r%�bX����\���0�ZՒ浫��Kı?~��6��bX�'���6��bX�'���ͧ"X��3"~���v��bX�'��[�k��S8�SΟ��N�������t�ı,G���fӑ,K����ӑ,K������r%�bX��r3�ӻ�,����)��79]��m�Δ�s���?���}\E�	���(� ��mr�7Y�T4��D8�h:Ȓ�l�=Cs���J�eyLDl5+콴�u��Yư�aN�ż/n���
�#=����"��Y��V��vzܦh}����ۜ0��!gJ�B����Վ�49�Qղ!sI�G���43�պW ���\
��liX,���P��S�Қ��=�R��wx�^Nd����vn;�Tۙ��'����2u&��v�T���
�z�7PƋ��N��X�%������ND�,K���]�"X�%���w��Kı>�w��Kı;�]'��sZ�5�Mn�Y��Kı>���Fı,O߻�M�"X�%��{�M�"X�%��{�ͧ"X�%���L�)���$�R3WiȖ%�bw�ߦӑ,K���ߦӑ,K��=�fӑ,K����ӑ,K��w�)}Mk5.f5�M�"X�%��{�M�"X�%��{�ͧ"X�%��u�]�"X�bw�w��Kı/�Y�/��f��f���SiȖ%�b}��iȖ%�b}�w�iȖ%�bw�w��Kı>�w��Kı>�L��\4L֑��^���u��lڒ'��|��r�Ɨ3p�y,��
�Y�	�`akn��:|:S��b}�w�iȖ%�b~���m9ı,O���m9ı,O����ND�)ҝ=������aZ+|���N,K����i�D8��"dK����r%�bX����m9ı,O������ҝ)ҝ?~m��vG7YL��iȖ%�b}���ND�,K���fӑ,Rı>���Kı?w���O�Jt�Jt�������[u��˴�K�������iȖ%�b~���v��bX�'{��m9İ?������ӑ,K��u�Y33Z�Y�Mnf�iȖ%�b}�w�iȖ%�b~�w��Kı>�}ͧ"X�%��w�ͧ"X�%�}�����3.��!#�6����K+7�Σ���8���x��'Tru�yq<����k�5wYP�f���ҝ,K�{�M�"X�%��{�m9ı,O���l8��>�}��A?_ߵ���VY��\���N���߿��D�K��;�fӑ,K���w�iȖ%�b~�w��@�,K������S\"+�O�Jt�Jt�߽�yӑ,K���w�iȖ<��@#��"�G�j	�Ax���5���iȖ%�bw�ߦ���N��N�w�ٯ��q��ew�Ȗ%�bw����Kı?w���r%�bX�{���r%�`*�����~y���G)�r�K����j�VK�֮ӑ,K�����iȖ%�b}���iȖ%�b}���iȖ%�b}�w�iȖ%�bwݓxL�s�a��@�f��t�Q�|$�	�� ��� �ꫦ�Z�� �X��8�o�߶��ou��{�M�"X�%��w�ͧ"X�%��u�]�"X�%���ߦӑ,K�>�a���H��eevO:|:S�8�>��ٴ��,K�뾻ND�,K�{�ND�,K��~�ND�)ҝ?}C�ej���:|:S��b}�w�iȖ%�b~�}�iȖ%�b}���iȖ%�b}��iȖ%�b{=�/��SZƗR3WiȖ%����{�ND�,K��~�ND�,K��}�ND�,� 5�j	�������r%�bX�g�����h�K�n�4m9ı,O���m9ı,O���m9ı,O����9ı,O��p�r%�bX�{W��a��ʖ�j-%Ԍ�
�Ŭە�f
�c�����lM^g���XW2��&Dryӑ,K��;�fӑ,K����ӑ,K�������&D�,O����ӑ,K��S/���MKunf�Y��Kı>���Kı>�}�iȖ%�b}���iȖ%�g+�O�r�r��G)���m��4�wd��j�9ı,O��p�r%�bX�w���r%���b}��iȖ%�b}�w�iȖ%�bw���=�j���ۚ�ff��"X�%��{�M�"X�%��w�ͧ"X�%��u�]�"X�%��{�ND�,K�M=���SRܥ�u����Kı>��ٴ�Kı>���Kı>�}�iȖ%�b}���iȖ%�bt�"cE�hJQkRT��"Q��
`QqhFؑ���hV�!E�	%Q�C�1m�
ň���kR0P��c*X	)JFZZB	��V�%%!!#�d$���V0 D�A�H�%%��"@#8 �ѡ�B
U�H�# �F%�	FH16�Q6`I	a�n�!����$�v��~�BE#�F$�"BHBc		#��<�j��%h6�(If�����(�B�b@�D�R+�EH$ �R41B0� ��"1�X@�$R2���;��w�O���U�eU�B�]s��bHJv��j�n���N�<�UJ��6�e�qtL���3�Y�m�$�eE@)tBV�S �^p���f���4On��JnyA��.�(���.�{��F�G���� m��n�vHY�Gn,�7$m�������R�.&%]`�'�B�t��G4�v7.����vS4��Wc��u��Eq�ySҺE�8�����-R��\=b0�Մ֬�h4�V�-�V����>Nwdz�N��3�m�v�Z��e&�Ī!IV5t)����[fT���P�`�T��F+*:;���C�H�;��++�P�f�k��L��<I���Ԯ2�j-�_�\!�,�DcY�����8�Kl�1���5^՞�,Ն���f�X��*P5iT�µȀX�ؖ��1H뱽pL�3�6�L�\&�ܖv��r����7��|ڒ�5	��H��R����n�t ����l��n&�Y�p������ù�sx���ք��T�B�"ev�Y�[���sK�aL�9H�9qi��$3I�[���2�4��S��ѫ�eC�QK�6��sS�]�B�J��[@Zv�\0��w	�B�J�Ur����[,�5J�0S�@�C�����PGl�^B�`�@(.���	�h؊�룄�"�l5K�&��z�v=/mK�K<n 6�xQث�e*4�TuӑY�4�N�l :^j�9��˚ ���]���띷)�T�\�h��\���V�h�c��:�7��䉎��u��5X��lt2����+�][�r�Kŉh�pڟn�A���q��[���3h�6�V��'tL�M�
yM8m;m�.wnD�z��[pqɜ�v�(�4:�����8���Lr����4*��ԋ��X
�F�Q�1����J��Q_<\�la.P�9�j{�R��lP(��:6�`��.KER\Q�n�xƔ�Am��M�h���"�TT�̋7I{v m�y��i��wniVUl�i�P�Q��U	j��o{���G���Ab�P�(���!�G��t �T�.vf���������i�E���T����%�����	{x���Ɨ�lm�rE'gA���)\YYb�D%(&�y�a݋�n�X��3X��Nܹ��i���g��˷I��ԩ�XI$ $�i決З]k�l� v���+ָ8\�b�5.;qp/u�8��,�v:�:�Z	��I�r��ݵ��d7s-�`,#`�:���5/�/�Y����**��֔n��$c�	p��q:�qu�8u�(�w��N��P�,h3[�y�ӥ:X�'�����r%�bX�w���Kı>�w��Kı>��ٴ�Kı=���ɩ�cK�����Kı?w���Kı>�w��Kı>��ٴ�Kı>���@�B������hF�t���X�%��{�M�"X�%��w�ͧ"X���C"dO�׿�ӑ,K�ｿ��O�Jt�Jt����/�fu�%DsSiȖ%�b}���iȖ%�b}�w�iȖ%�b~�w��K�U��~�ND�,K�{���!��MKr��kY��Kı>���Kİ�=���6�D�,K�����Kı>��ٴ�Kı/���,�U��eF��2Y�n;]��z؎��O7q����I�\�%RvM���j>�~��ou�b~�w��Kı>�w��Kı>��ٴ�Kı>���K�)����E�KnquSΟ��ı>�w�� *E��dL�b~��ٴ�Kı>���Kı?~��6����TȖ'|h����4jj[��.�56��bX�'����m9ı,O����9ı,O߻�M�"X�%��{�M�"X�%����ORf\Ԛ�dі�k6��bX�؟w]��r%�bX��w~�ND�,K��~�ND�,K����ӑ,K��Ot�ə��cK�����Kı?w���r%�bX�w���r%�bX�w]��r%�bX�w]��r%�bX���t�3Z�^H��5��{=9�y#�T`ˈ*�>3�l1\kc'D�-���$7}����ı,O���m9ı,O����9ı,O����?� }"X�'�{��Ο��N��߯��f3����r%�bX�g{��r%�bX�w]��r%�bX�w���Kı>�w��O�Jt�Jt�����)�-���Y��Kı>���Kı?w���K(�P"4	Q?w{��r%�bX����m9ı����S�ԵL����<�B��{�ND�,K��~�ND�,K�｛ND�,K�뾻ND�,e:~���裆RۜSfy��ҝ(�'���6��bX��$k��ٴ�%�bX���]�"X�%�����#�/P�N>��A,ME�hK��t�ve�ma�.� j���h�m�g�x��[F۴����O�Jt�Jt�߽�yӑ,K����ӑ,K�����ӑ,K���ߦӑ,K���t���ю��˼���N��N�ߟ��8�?�B9"X����ND�,K~�?���'� �J_1�-YJ��&�`ݙXwnV�xu�XV�BP�n�E��m�`~�s��g��'� 9ʪ�;\�q������B��t] �e���:�c�;�b�;�2���0��Jq,��wtq7iR�r֣مū03b��]2fC��1'L7����/Lvu�V�"�M&���;�b�;�2���0����[mFjݠN���ٕ�wv�ul�  �i)e�BI؆���0����W)/G>X��V�a!c�Л�t��0���ױ`ݙXwn��P�uv1�M�Xu�X�fV�ۆղ<p�r��{K��a	z�f�lu����N�*�ț*^1�<�`�jܔ`6�>�8�����(�ܔ=�.7.R��պ,�A�p[q��C�K&��δv2�`��.���1�r���;�R�Cecp�d�@9��70S�L�b	�E͗kfv�'Z���v4S�9v�d5Z�ɨU�S7lM���6�M�C���+o&@ν�4���m���?�N�۟<���UIvK���gE����q����[w;#We��vnF�)Zp�qr5%�	vo�}���'�wv�ul�  ��hJV�`էu�wv�ul�  ����	媅J�Ђ��[� ���{�ٕ�wv�yH�d���J�M&���ױ`ݙXwn�C�Ͼ{����S���L����n̬���H��ذz�f[�/Wh#cr�,�.��0<��Y�2ݕۯ[h���\n'v:c��i���[���ۆ�$xu�X�fV�a��
5�2��>_�o7I;��Lůb�7ve`ݸ`��"����e*�i'o  �ٕ�wv�uI)M��7e�)R��ݬwfV�ۆ�$xu�X�ք��W�[V���ۆ�$xu�X���x����/�u��of�+j��CB���I�-���S�JWF�]+�Vf�i�R��B
VYn��H��ذ�̬��T���EV���M���w^ŀo�e`ݸ`Sc�'���MRt�V�wv��̬��=\��s�x�J���xE҇�/n����`֒�v+�I!�N� ��� ��{�ٕ�{Xl�j��-�ҺM�0���ױ`�Xwn�����bI�մ��t��I�4i���N�G:볋�c!�5R� ��P�uv�]4���o�ŀo�e`�p�:�ǀDM��7We��X!�X�fVٷ��<|�, �m
�IYj���V�͸`^���`ݙX���(�+���J�-ف��|�	�|�n̬H�Ur��/�� �$bHc�R�@����9{�e:Bhպ������o�ŀ{ve`�2�����'RI�}~��Q�$��Uv���+�B�M���/�4�5�E�鎹��͵J��:M�v���]d�+ �ۆղ<|�,u��Gce��lCwXf�0�`�`ݙX��eX˲��t��n���X��X�fVٷ|�i��\Ut�n��{�ٕ�vm��qz_�,�})/���i
�c��{ve`�p�;�E�o�ŀmJ��UW!7�wv�l�et^���֩,7�VBm�͵e�d���F�˅���)���0g3ܽ"�\'$[h��vɇ<i��v������)cm�i��:��]aWj��,�-��d�'�+x�X�`��حs�Ц��ζ�"�j�msV�x�8�n��\�{���k�t��7L
��v�=u:.�>Z2�&4���	q���:2W���cj�N��I�#�Z3ƈ�W���<t�v�cYcGC,���
j�ܒ��e_��O%<�P�ڠ�i����ﾾ�����{�ٕ��[B�Xա+,�f�r,|�,۳+ �ۆ�"��Ҷ�$�wwk �=� ����;6�w\� ��m4�
t�i�n���UW��k ���0�`}\뮤9���v�q���#�UӺ�p�;�E�o�ŀ{ve`S�3���ʖ�ٳ���=���$�if��l{�{,�W`m�7j�:��^.��<�V��� �������lۃ`m�3�`\� �����Y:N��%1�ݙX��0���i)MղЂ���`ݙXf�0����`�AC�UՍ�m�n� �ۆ�r,|�,۳+ 7Զ��l��
VYn���X��X�fV�=ܽ�|���j1�(�ܣ].�ut=;4�:�
�k��;a��j��x���ŵ�v�l��i;�k �=� ����;6�w^ŀOm��R�t�[��XwfVٳ+  �=� �4���Z|V�7u�vl��;�b�z�(��$�G�HE�2E���+� �R,
�F$$*��BI ��*���h� ��J�D��+BR$�8�儛��XЅB?!A>B!7ςYX��ȥB^U�1!�� X�2� Ĭ$8��JA�D�$! F�)@�4B� �qH�-b���[��w}�C�� D�JI>6i��S����4�
��n.�����t�!�Nl��M)m!eO� �@K���iB|.� �X�C�녴�
!m\�� s��H�aq�D� ��J�[H���Oՠ�!��h��ΰP@�~Dմ��U)�,
�4$b�Q���8��$�(�D���t�E(� @�#�����)�������u^ &�V���UV-o"�;6e`P%KV[,n����`}\�������>�>XwfV=�+ �nZT��-Z�WBN�<�,��+ �ۆ�{ o�0ϕ��n�mu�û�𬞢&M��Z��,�ųD�2�gL�Y�p4�6�7�;�2�	�`ױ`�b��P����M�J��`�p�;�b�'�ŀwvegܮq �JQ�V���
vU۳ �s�O=� ����'��yH���]'VЭ'v�`�b�;�2�I߿k�rw�T�#�@$BQ�v����rN���.[�e��5f���;�2�͸`ױ`�`_y�s*��J�]n�;j�ۖ��t�2Y��t'U���=pT9m���t�t�LCwXf�0�ذ�ذ�̬��j�vq1�Ҷ��;�bϒ&���='�Xf�3�H��ZH��;-p��'k ��� ����;6�w^ŀDM��7V���i�XwfVٷ��,|�, ��U
j��t�4���ٷ��,|�,���<�Q���
�`�@���}�i�D��;V�u%Pɑ�(9vjal� Y�h�l6�6�/<�m�kr��㳬�1P۞�@A��mv�X
�;<��4e��X�ռ��ɭ����vM�CiH��ĬR��&�@i-rY�6����J��,�ݖ)�<b�z�ga4c\n-$��[!�����j���=�#v�h���莦��v.%c6v�F��i���$���kZ�Nɘ�u؞Ϳ�M:��S:%�/=fҺ�SU%��t�+Z..	��@����,|�,��+ �ۆ H�)Bv�IZN���7�b�;�2�͸`ױ`�m��M��cwv��̬�n+�Ľ�`\�`ᨈ���*�����ٳ+  �=� ����JR��[�Ʃ�ҷwXu�X��XwfVٳ+ ��ӑFUn������.�W@	�P���4&3-���:���݅�nW�ڡ'k �=� ��� �ٕ�w^ŀDM��7V������;�p�^�s�Y@h	����P2o{�����,|�X��J�]��i]ݘ��0�ذ�`ݸ`I�'WWM�;,�f�r,|�X�n��0E�M�]%i;���o�� ��� �ۆ�r, �*�g(�YH���Z�k�,W;�Oft'i)��<�CnD�H��p�՜�k ��� �ۆ�r,|�X��Dv]2���N��=6�w\� �9�ٕ�yMJUڴ���at�v`�"�7�E��\+�ʮ\���� �ۆ&ۈ��h�i]�x�Ȱn�0M�`[#�"&�R��Һ��v�n�0M�`[#����;��O���Sn���j��k��\s�+ї(�/9煰$�ݮn�6������lE�ـzm� ��r,۷) Є�.�
vYn���X�Ȱn̬�n"��vZ���۵�o�� ����=6�w^ŀO=m��][M۵�wve`�p�;�b�UU�v��UT�^ŀo��#��ua�lCwXf�0�ذ�ذ�̬/j#I�5P�\��k�F����ݕ�@�,�΂���tu�H7P��mb�כn]�xϻ�X��XwfVٷM�I��v�(�v��ذ�̬�nV�xD�JSv:WE�7k ����;6��\�^R|�	�|�wP�J�lEۺ�;6�unǀo�ŀwve`M���Zi"���v`[���`ݙXf�0r��������+��1���C�Z�g����]s)r�n�í�)�Z�U�Ĺ���]�֮��ʇV��Fk��A҅�m+��&�6�0��.d�Y��	�W]h���A�(u� �76'�Z�48����<D�v��|���QGn�(�{	sݚ��r��2V�#klL[��k���ã�f�{b�݈�V���j��8�V-����h�$��wI�t�|�N���m>b�"�s�i��1z'ss7 ��3�v��n!7�,�y�:�,��hV��v��~XwfVٷ��,y�m�Đ���cwv��ذ͸`ױ`�`ᨈ�բ�wb.�`�p�;�b��9��*���� �s�uM��һJ��t�v`ױ`�`ױ`�p�$�d�i�e��.����{�{ٷ��,/P�aJ��i+��j�b��&nE�'ljZ$ s^�G76'-SM���3�I]7c��E����;�b�;6�w\���	�|�l������WI���ܓ�������;F($�jR�@b�X� Č-Q(,"@$0J�b�D���_�,y�� ��� ����m����ݘV���ذkذ͸`�$JNݡ6�7wo �=� ��� �ۆ�r,y�m�ēE+-1��X��Xf�0�`�;����{�*�wX1Kb�=u
Zhe��gZ�J	�'�JWfC�jy0F�"8E;�v�͸`�"�7�b�=�b�:��YcJ�*M%t�v`�"�7�b�=�b�;6�I����j��EBN��{�{��9ʭ�+��s�ʪ�fl���6=� ��IJv�ƇE����=�b�=�p�;�E�{�E��J
��t�n�`��`�"�=�"�=�b�7M�
�����J������[s�%$��4�Q���@n�
0jUKJUU���꧀|�"�=�"�=�b�=�p�"�H�����j��۵�{�E�������� ���0�ذ󍶣�R�����w^ŀ{��w^ŀ{�E�o��x�&��t��;��:��}���t=�`�`.r�«���{�4R�VZ����ݘu�X��Xu�X�.��QEJ�+wN��x�����$웲T���p��IF3@+T3f����m���v��EBWk ���  ����s��G>XR1}I��halCv�{n�.|�,�r, �m*��;�*�6&���=�p�;�`�`��0	�!
���ue:M]�|�,�r,�ۆ�K��H�);v�n��;���{�E�_�~�=>�~�zjI�g߮��
����
���Ȩ�*���*�QW��E_�TU�U�AT��@"�P��DX�E�E�@DX�"1DX�"�E��A`�0DX�,Q �E��A`(E`#E�Q(�DX�DX �DX�DX���Ab#E�E��E�E�(Eb �B#E��Ab�A`�AP�0DXQ T"P��`0DX�B(A`T 	E��P�Q*!E��B	E�AP�P�G��QW�
����**��Uh
���QTU��EQW�
���� ����*�Ң����E_�E_��PVI��y����6` �����[#�   P      �          �  <�   %U"PU%����*�%J���*���*HU P ����  ( �I��H ��   � �   �Af �)@1��� g����  �)c:�k�w^���K��t�p>�s�K���=�5� ����Ϸ)p :ܥ���95������K �r���ꛋ���gO|��7��  <   @ P �� z��[�9;��x��ri�� �^���gJ��ܻ淼�W� �����{J�wl WUX�R� /=*������{�����Ҿ� ��qwi��:U�e�r�Up ��@ )@ (d w�Vf+���e��+��T�@S����0뫾�W&Ub�Tr�>�>�x��w}Wݽ��z��@=����^��R�{�}�u}��� y�^��*�x����ۥ=�]�U�  =  ( (
c` {�>���s�m9w�]�< >��/�ӛ:ӓ��;x�v�p v[q��e<{;� u�|ܩnΕ}����m�'�������o;x�:�� ����唻��ͯ}�={}��ϼ��  � �(  	(*��E�U1�}om㻷��&���
 ��  R 
 �  Q 6       � ` 6�)J$

6e(   Z���� iH@ D�t ����*T  �������T��� �"x�T�"l�da'�U$zITOB B*�J=�R�  �!M�)D��#�6'��O�����Q�۟�-T���t��P����p�DU����UWT��*����*���ª"�TPS������a��X�JLt��`J��d$3{?Ԑ�	���"?�	 l6���i�kg N@���A��!)���|a$$BW�0�����[	$B$aA���`�*H6���M!]��t�c��\ol�q��k���(�h�ȄBS�kSP+�i��%$q�J�f��p�����V+/�A�H�7dZd��P։#��e�sF�bC �@�H��8�H@�F!Xd�qO�
I �GA��}�6��(B�f��oVo�G��cN3Q֩�p!3[��1(`|�Ӏ@"`CƘCY��a��$u�	����Jad��6��#$�l$�B7u"B��6.M`K��̺���]���aM$��,+��5��0�%�(���5a��BJ^`C��5YO��䁣�#�4~�����`���9bH���5���f`K&jqtJL�HY��G	y�!�+5���Fٰ�&��0�	)AB�@�# `�)��a?F$��p��		��	Mư��%��6�o�ka���Md��6�~�k��~�^)ZE�pE�PMP�%)
EM��!�!��Z�bC#L�Vf��`��JI.�T�8B�|�FJH!w�\�.��d5!�I~��e�]ka.���\f�6q�0��T��
p�?�3����c6�T�Z1����,7���zHcLc%��C&8��,�p75+��p�Ɂ����ku!J9 &�k�ӌ
�(��@ �!�#*h�T F,B1`:`A�� DԄ���)�N��`px���hӵ�t%�|l�0���̲'��\����5��oZy?h	d	��!��&g��[?$�sY�~��3���)��4�bE��$t�"95�	�S_��B��i����t��*q�����?d6�, `ʐ�
��l	�C.��kt# �p� �CC|��&�.�o���MM�D���|N���MK��I3N\�w|�yL/柒��4K�o��񻄙���� v�y��n�[sR��F\��;'Į��!
`��9��)����@)�M#��
`���5
����Ì�+��K����|B��B�a���f|^n��/�
� �:�
�k�+�lę�nP��XT�tM�dZKv�d���0�q�r��*hp���	&��g�]s8��j�@F*H�o�������\H�A�x��
!\t�s�,��5�����5�#Wh@���|X�5��~�L�]�"K��޹�z#	�f�P0#74KKLYC	p�!�ٹ!pѩ���E�ƌB�$B:v�ŊCF������a��2Y�ָq)��Ą!�]�����p�M���R<aL4�X;8q�#pѳ�"�0\	L����0%f���aM���9�9Њ�e���J�)�	���m/��޵��SCxK�8~��>y�y�)#��\ϯu�n1�0������V�" � 	��XH(@`�b$BQ0�0��Oε��~3>���ٮkm7��?~�K8����i�D�8�)�.@"��L$%1�Lso�_��q�/̬H�,d�6ns��	S$��~���?<�	Ëk��� �B�����FN,�AGxo|K7�n�㹵��Ou�wu�,/wonx�q"B�&5�R���f�a��S
jP�C7�xh���3sC�+��B�o!������4�~�Z$��s7F�T���Db��h�棳A�4n4��N~�1���!]�.Ną������$��7�s9��).�~.m����?��P�HQ��1 \P�̘m��-��\$��"��B@�C!��)�
���k2`B�0�k[�.h�q��!�*�0��d&ɬ�I�h#s5v���ѓ��d.kdt&a�L�H$5�޴kf��I��B�/&�.i����:v1�F�Q�� D�^k5?���|�M͜g5�r^]l�4˭S'|�k_�ɭ���p�x��fB�! R�+�&��<��o�1&�r:�)���w��A?��FԉV������"%"A��e>�F0`�N�`���8��$)�+�%)��~��Z������)�I��K0!avf�RB�s5K/�e�~a(Hf���c7�J6���o�X]��&�!��&l��c�p&�q��*K�3�)� Ƥ�F��Ȑ�
5sfa��5�f�M�k leMmȑ�IP�Ӷ#A
�ˈK�Jc+72�!�"Bqp W�[�4nk��5�jBK�_��y	{�~�)-~�b��� ���D���L%��\���6XN�fC[y��
�!BM�L	I��C,��Fb)�1�����{>!fjܬ�9�f�u��|��4�n��<�rBX�!�g�W�0���$&q��~���52��?c�Ț8��o��[�OВLG��?p����?^8o�F���܄��5	.s_��\����l%T�v�� �?�hlHLGK�h$k\4�*�i��1��HXcB8����G``?��\tf������k�B����8!��7����;5]����Ѿ_��C�|���'ف)��7��:a��R? ~q!p�l��6�A.&�F�����z�������P��CJSZe��_��v�l	����Le6i��\�/)Ĳ�-����z��l�9�FH�Xf$.,! �ČH� ���ka.�@#-h��A��s���T1a��''ณ�!o���'㟹�7v�ؑ���y�o	����|l��&�n�c-ѫ���8�H�T�i2d�MA���
B�&[��6�5�x��7�@�HLލ�lۃ)�e���a�I.��٦ꕤ��q.�8�#$]5y��f�l��9�cH$)3z%$JFRx�p?k~H%a c �*�a��y�!1�8�BF��4�(BD�"�
�	0��o�K5���D�)I�1%+��HE�F��!\i�Y��~e�l��1��F�VL�K�ke��0�����s\0
V����S~��]�&\%j�$#�6�E٣6����4�4k�hB��˚�qp?��d�ACf���\�m6�a�� ��nr�韌��4b��;�ˎ���c��Ha�N�����'�(����ӵK��?�:M��a���h!S��o��0�~�����dd��)�f�a��~\a��~��h�1c�HF��L�K�b�?K�P���`B�?��@�j�!�6k��h&�V�c]���t,[�f��SKkL\�	f�:XU!r�����Oߍù�a%�%!a	�<�;8�/h�3��I��MP�DM���8~��~�����6ː`��GA8a)�G�j���@ј��&0�A��Ԥ�Ӹ��W@b�d��a`qE kY�Nl�6~Pt��Bj`lhF A�u7���%)&�4ֆ7n�ؕ�p��>�o�Ԗ@�]l�bK�p�	$�D�~t�Z��������.����?&�1!���F�JV�����l�k2[V��9��A�F��!x�y����B��f�WҐ
$(E(����k�0�@�@��럿@�$
��P�� �A���C��1�Ё`V d�1�݋����b�D�%/����E!!�i7RHU�nl��9��!r�� �Zj�\�4%CaĊ�5p�kL4������	M2�	��0$	C&G�k�jE�g�w$�i��6BD)2ST�� �Q $q�A�
A�)�Rg@Ç?]�'�h86#B��H�,jJf�Nh����j�s7o�I�A>Hc�$&3`R$Lu6ea�n��#5��L�0�5��3+5��H��	LasLk
m�H�h�	�4��L�B�(:&�e�Ra���k\��ˁ�f��ͤ��1%�$5�	fh7��3C)%�+�h�L��-�.A��F^�Z�`�R^�|pX�4`H�|�A��$CS0�� %$_�*]��i�!�w^I
�{����2#d�u��O�J@	<��N;[���"��4�_HI��~����� m��m��   [E���O�WRi�2���ؠ6홉y�]: lh���r�  $	��(iϦ�}��p[@M���m�K����F� ))%� �I۳-�6�bOHĀڶ�M�v�l���(������   � ��m�U��$ m4�Kn ���%�>o��� -��	  �     �7m���s��SP!�A -:M�p �l�6Ͱ<G  M�m r��` �     �p  6� �q�� 	 6�k���@hn�9 6� �a�q{Vlu���I�s� 8�oQˢБ!�Ͷ<��cm��zƨ�m��n�  ɴ�Cm� 6Ȳ H  m$�۫i � $ 6�wYm�'cm��	Z\�b�H�nEG(O�٪��U��]����e:�]�C�Vʕ�h�w=%����'o�m�XӪ���;,��-ʀ��n��]6��� IJ1���R���R^� �@��� J�u�K�u�u[J����-@UUVҭT�����/Z ݮ���׵�]{F�  &�i@�I]cH�i���P�Ԣ���{*�KR
��UQb�����Pv�` �׶���I�tn@
%����M�8p��*�� @V����j������yvh�(�)g��]�Uc'��յà�v��]0�];^[i�n�% l8jnH�Ê�M��ʵA%	oh���bBn�u�U�aܗ5��T��y���7#nbR��/f���V�ݳlp5��mE�N�	�)sk�\��205����n@����q�z�gj�6�&� H�!:C^�:rn6�f�kn pp���@�P  �
�K��2ò���l�@@��q#n�@-��Ŵn�δ	l ��	ے[ �v���[Ci6�h�%� ����-�H8��wf�[�_9>R�:t` #�^���%��I 	 828ĵ���V��� �[�e���h� �ٍv�N�I7cn�VM׎M+2�J�� �f�,�t��	ȶ�A&9#K��ƚPx��$ۙ@h
�a�:69-�cKD���yc7I��U]�8ږ��V��3�� <�� ���>Z��N�mv�m�֕e�gXl 7I�L${%8�Z]��0EꠍMJ봘 薒��54͚�G;�m��4�6i���j|R�\YZU�A�m�#*��TmY{���K���rCj�6p[�^��t�)z)�,�vX�^�;V��%�Pj���$m��v�����ˬh��a�� �[zv#Om����b��n�R^Nݦo6�h�l  ��(�B�Ȑsm:�6��܊ �R�K/[�I�����[(�D���jyP*�����nx���1eP]=k�*ҭ��n����g:@!1�!s'��sUuQT9-0�\:�iI-�v�VT���ʩ*�q�檪7C�:M��;-�ڛWYM��s+p[�ۜ	��-�v�Zm������2
�ҍ�m,��Um^�Åӑ%����T lje�iUZ����-��O��RY�4���ۻ_�9;k��v���h*�+m�j�V��@Cv+o-8�ܺ�Ü	 �l����l�j�r�U�īT�@�U]��`M�`sd�� -�ӛ����[UJ�RҜ��l; Z��gNi�m]�=�+[#	[v��	�uf�m�I���ޒ�6� ���u�]Pݳ����}�m%��`��m��v,�e^ϟ+� Um�����7kmm�-���
N�gM�lnԫ6���z�j�:F@��2��6���Z����$�&���:B�g�j��E�@]1�t��v�mA���ky�$4��$����|A�wI�pSm���km�
ye�6z�� ���UCă'[ζ��Xv���,�d܌�����UGg�0RU:v����o �Zkm��x��>/��J��Uu�T�޸$�-;Y` m�p�5��L ���p��TpF��vFۖ�c��.!��m�+�f��e�p ���3׭U�cP2�UUUīT�C*햨���˰A���įnE%N6:��r��;���@�����bX)Q��
�j���H33/"ަ� M��5��Z/i�I�l��8�h
8:�ۍ�U@��m6m��:��s��k��� 
�V�R���[jؕ��9d6�ڂ�Z)�8�:-� "ҩ���y6�^�m��m��f�Hm���bՌ�1ms�   ZpZ]M����@[A�j� ky�m��U^�e]�cv���*��EU���ZKH
��@Kki�X:��*�j�gbM��6�  ru@B+UT�����mpUl��9v�~F�3��%�1ͻkhH  ��Ͼ����i6�$	�m�o ��%��I�b�S� ��*�U[HA��٠ �,6n	��'dm�� �vj��pn)j�qm� t�I-g)ƫ�0��H �n� m��  Hv�3l m�8h�`86�6$�#t��m���I ְ$4�,�k��&�`�&�m�۶@�a� d�qm@m��i �k2ۖ�B��D�TJ�Tupm�!�[p	M���N�8ΎX\�%�e�]6Xal�   5�Ŵ�m���wG  � �m���� �[IZ͖� ��xm�� q��wc ����[nBJٴ�J���Ʒ -�@��f� c$N�+Lkl����oZ�]u�p��UPZ2ʰ�m +uu���2�TX�[�����QV��mJ�[���G�@ �.���ibg<�+�!X
�M����|m��  ��Lpi"�  �@8�m��v�am5� m 6ݖ�@����/P��d�	�m��.��鵿}�  ��v�UT&��i��U*�-EJ�۵KQ���ko�} ��	6��  "D�H �v�"�n�`��[Rmٵ�:m   WN��jˎhsl��N��r�j��uj�aɛiZ��v�dK*ʳ�&^6v�Q�U[�6]�	�lZ�j�6Ͱ-��g��F�pq�W!5�IZy�*� ��ZL�U�����5�J� �2�X��0$�JV�AH�P촺X��WbZ�-Mr�f�=r\h6��	@��k��b���{GmJ��l�&*�u]*�J;F�B�f���p&ucf��;1N��S�5�j�j�I�&U�R%�6݄�  :�n��  ��L�$�    �6�� -����I�fI,��-6�ݳl  u��  Y��sm�m��-�� 8�km������&��}nؐ$ ֤�BBڂN��h 9�( �5���d�e�m�r�]��l5�k���V�������-�d> [d+Tځ́r�$6�^Z� ��m�N���` 7hֻl8dqm�i) �e� ���nH6�I��:G:K2e�@ 6�NZH����i$��-񓔒�0�Kz�Sd���7k�fض�����`� m�ڳn�U�� u�6��:�8�� �rP�m�f�kW[�ZmK��� �eTpUW*Ғ�ThYvx�` �i���v� ܐ-�[n�-�6A�=kv�5�G��,���iV�S-�Z���#+��[<����B��u�km�sV�K�pj�V�������[h-؀U� *��z��Ry��Z����mI	K]��m��	8i7�   $ ��h��@ .��p�+UU�Uus�Vv�䃆�j�m��&�� ����'�  m�s��V�m�m�N�L8K4�:m�16�Y@s�[I�kV�tͰ	9Í��n���&�!��n�Wn��$8 �Ӧ�'Tv�t�M��-Ok����M�,=�C�ڜp8�t�jͭ��9$�OU���n@m$�]$�)IMR�ʧ9�[.�g��ZΖ��  �U& U@HK�ʏf���ej��
W�I�*�` ^�5�m�umU �mx  m���c��߾��v�e(5��h �	e��b��	 @	 :��}km��� =6�6ݖ� $6�6�fݵ��� m�HsV��q �� �� �`   �-�[,� �� �'n� ��Im 	 �� �  m�� *����6�/(�4��lG � �ZN٭��i��� 6C Z���`8 ��Y�I6�l�p �X��M�      m� �m���m�H [@P�g P�j�rư���U��� �fݱ�ݰ��[�$�`Yf�V�?m~������Ӗ�fm���Ƙ�j��n�i�@im9�!K�Qګ(�T!s(
��.t��@�I�[M�6� $  �L6C 6��m��kP` 9��@� [@���-�3-�]XCY��j� �h�F���?�P�@�?*��R��tڀ��_�@`b�*�9PX!�(q����( ���A�A*��]��P�q��D@₇�TN��p�|+"l�q@��*��� ��B�Q�Q�X
��"`|�x��?�h������Z(D@�A�����Ҩ@(!E��q? �P��51�@01��a @AD�`@��1X�#�HB0�@�t���pP�@�� )��S4��_� �4��b5� `
A�l oE~G�Qڡ�B0R0 ��Q
��S�PD�M�8�E6�
?��Q:��Q~P芧�O�G���-
  lP b�"A^#�  �P
���#��*������?F�������� �eg���� ܼ��@�l�ɀ�`�ZB��lr6�tLP(k�N:Ɛ��n[
��UK�<������Mz�j�qp8�{T�)�j����Wjޘ\���Rn�GYM��{Ute�H�t�N;p��I�Z��υ'h��t�ݗWv�������ӏn�����L:�qs���hwUqŜ��Ͷ���+NKc�6*6�<�g/b`���e9��$�q];t[8D�u&v��'�_.�&����P�[���q%��Bƣ;�v<O=�$��U�+sP�Y/6��#\N�&+&�ħT���&�Ӷ�7����ivS��	D�\�g�t�[tX�]Ḯv�f#%t��g[E�mm����93��`f'H���޻.��f3��V������SkXعer Xkx��Ѹ�U�6�Vi-d�L\l��C�J5�n��9���q6- / ��N��Ԇ�m�N����ϋ��ѱ�-$�39Ύ�ӹ��8�i�-��*�I�����۵�����FSdpXp��xخwd:�x/f4*Ifܫlk5�m�;�
���m�2�-pIN���=�a`��=�� n�ü�	��`� ��왺��L-��vK�(�����uϚ�qE�M�ըUV�aa�r�W@:Ki\s.��f�E-m�n�	���=���qu�����\�]����<c���9���2`U%-b������RY[��x�f����
i8�썵[Z;A��sT��v�9�vH�p]^�Wq���s�r��`t[*��@�w;nIsqΖz�-�]NȄ�DY��xJEӷ8,�#�Q���l��.����3���Π�0-��l�Vm��LY�ZZ���m\�9ɼ�ty��FMnyLF^:��gN��k�����@B69�V�vM�ꪨ�]��^��TjUh]�)��'(f9�-ҀܴUJp-U�[����h����I����x�m�H:�"^��������{��@O�H	X, <���P�LG�G�~7�R�Mk@Y�$��rE��P�k��S�u컨�S� v�|���vvx����ꉰ�r�k�غ�^1�v%u�U����ָۜs��7AU��.MM.;&����y�x�w�6��d���</�/�㵷9w�؛{hև�hx�c�dl�S��֣��Ø�`:.n��:2i��j�ZD�nup��������{���>��.M��,���KB�e�Ǎ��� �;��&xL��e�
fK�&X��?#��zpO��ɢ� �&���&��	��ϲ��h*ODȖ%�����r%�bX�w�6ˣ�X'ձ������ow�����rU9"X��粦�X�%�����r%�bX��{�*n%�bY����~�u"�R/=ߛ�oq��O���"n%�bX�~���r%�bX��zl���%�bs���iȖ%�w���~��孇�7C;��{��7������ӑ,K����eMı,K��ݻND�,K���ț�bX���w��F���{�7���{���zl���%�bs���iȖ%�b}�gr��X�%���ͧ"X�%�������g5�2�W{ N.4Ի7�q���8:ݻX�k�l�ݱ�sl/W&扜���5�*n%�bX����r%�bX�g�ܩ��%�b}���iȖ%�b~�鲦�X�%����f�jkZ�5t\�f�ӑ,K��>��M ���@��EP��Eۨ��bg���iȖ%�b}�鲦�X�%����ݧ"X�%����BI ��)��5�4���������_3�bX�'�ޛ*n%�bX����r%�bX�g�ܩ��%�b}���s,��.k$���ND�,K�oM�7ı,Nw_v�9ı,O���T�Kı>��xm9ı,O��f�S%ԷY.�kF���bX�';��v��bX�'��w*n%�bX�~��6��bX�'�ޛ*n%�bX���}ｮ��D�-v"/ V�����y|Y���]n{7�f\�C0��P�#Gb�x�]�"X�%��}�ʛ�bX�'߾��"X�%����ʛ�bX�';��v��bX�'s���iu�YsR�!��eMı,K��w�ӑ,K����eMı,K��ݻND�,K��Z��~�~�~�~��:Țn3 ��#Y�ND�,K�oM�7ı,Nw_v�9� �@H�"!�DdF��Q2's�����%�b}����Kı/��?y7,jM�����{��7��9�}۴�Kı>ϻ����%�b}����r%�bX��zl���%�g��������� ��,|�~oq���>ϳ�Sq,K������Kı?v��Sq,K��u�nӑ,K�w��w�9�	�T2�b���(붖w]
���/k�O3��R�ՎK���k5tdֵ�7ı,O�}�ND�,K�oM�7ı,Nw_v�9ı,O���"n%�bX�v}��a��.k$���ND�,K�oM�7ı,Nw_v�9ı,O���"n%�bX�~��6��bX�'��ͳ4S&j[��W5�EMı,K��ݻND�,K���ț�bX�'߾��"X�%����ʛ�bX�'?k���Z˚�%ֲ�Y���Kı>ϻ����%�b}����r%�bX��zl���%��Ȍ����:��sq.~�.ӑ,K��}�릗Z՗5.���T�Kı>��xm9ı,N�zl���%�bs���iȖ%�bw>��Mı,K��t��[oE����\��KgQ/D��]	�%��%G&�,=�&��-T#�[���]���B��^���?:�8�k���Q�A��s@>�B3#$�DI$���].�'J�zz���+��{w�Fӊbq��
������}�p�<���:�ŲF�Bn8�28��^0/O\]�0*�u�)=ww6,D��J����?m�`
"�_t��_V���y,�@�@(�� b"
���D���}�{��?�#U��[���a9�OiؽK�n��]�OWgY�F�'\ĉ[T{q��ȉp��R�2췷qݛ�Ȟ:��u�X�w`3 �g:�A�Ϋ�����]��v�.��gs6u�unѱO�]�}ǣF���f�"u���l����2!����7����_$�ʝ��ʹ�Z�٪��(���n�O�������ۙ!Ӗ�n,�m�{kk[<\%Zxg�ݹ��֤��=f�K �����wg����ģ[�n�ٍ��'���������
�]`I+�����է��|@R4�(��*�����ċoۚ�g�hWj�:��x�8�'�8�	%x��V�ژu��>��!�2E�8��4�t4+�h{k�;��h��̎)"��{����W[�	%x��\x���������˥8y�DI��zy�m���m�.xU��u<��Nv�F���h�e18�^��zw]��\��<�ՠu�\�Ȅ�d����;��j��~T������9ə����?~���
������y�1!D�h�ǌ�ژu���W��+�j�U�7D�]݆DDO��� ��Հwu��/�t4펧��hR4�)W8�k���m������M�m���_�F�u�,I�ݐJ�!v�k��q�y�kj�{j�����nBa�i���yo��$��`���Wuz�:Ȇ�k ��!I3@���ΈQ	L����_V�� =Z��E"CQ�@�V�W�^�S�"�^����{7$�ﻹ7$��E$Q��bq��
��������v������
Hԙ�����W�Ұ`}v�����m�}��Κ��7,�l<��c�}���}�I*m7V�5��T�� �.y�E5�3[�-[����ǌ�ژt���W�m˿��1�
9$��Z�k�w^,���>��������˹�<JH��Z˯�@�빠_m�hWj�=�Z<A�8(̉ǡ�%��� ��1`�78�������T�/TSR��f䓝�wZ��F\�r$�I3@�ۨ�<�ՠU�W�wu��<��du��c���r��(��c%L\Cr<��;;�s�7f�⡹�Մ�<ֹ�����f��v��z����}���;�.��6�Ɯ�-ϵ�tB�IL��ŀv��Λ������(��dq��w4�˹�y]�@���ފ�� ��A!yo��z�x���T�XJ��w�Y0c	��y&hWj�*��I^0/\�8*=@��^�u���aݶs<l��dQܽ	=���c��:/^�L[y%Ҕ7=$<�ݼ�מix���o1�l�N��[;۶�g4 ۇF;H6�3�02����� ;D�S%��⯕�Mƃ3�3��(ͮر�T��+m���gsG)הh�7˾gm^����z��8�H�rOnKvSk�����۱�Tݹ�Lm�l�cHA�j؋��{�ww{��g�p�u�U���V8�ڋ��Da��C6ċce�	m��.�Y%��"�<����+�=���}�w4+�hV�呎��ȷ���W��+��mL
���<�Y�inD�)&hۗs@���Q=-�`�ŀV�.�wwd����I��ڴ
�נwu��/YR�;�.�	�F�Ɯ�-�m��Q���λ��?:npu���ڋ��f粄s�uY|��θ	�K��c{%nϰ�v,1�rO@U4:e�$�m�`}v������˶e�csLԺ��rN����.�H��V,R<DZ���n䜿w�@�빠yn]��D�b�)1h]�0*�u�$�l������ȞH6���*�נwu��/>��+�h֭�Ɋ
3"����`���o���]Ӏ9�u��}��q���6?B|�=yqvרɲ��%��)�.ǩ:�n�ݹ��]�.�u�y{j4��H�X���W~Šy]�@��^���s@/���r j"8��ڷ��:w���b���`��\�eȤjLi���*�נwu����3'����1$�S�������42�e)0�ϵ��W��A�F�*oZ@p
h �pB���.�E����P�P6; @""1��b8���@�$		$�
J�^�j��Q(٤O�'�����AN��P�D����3�A�;��߾�y��z�A�lll~�|^f��֦����5�͈<����{�p؃� � � � ���,؃� � � � �����A�A�A�A�}�f�A�������t�3M�\�֍�<������r͈<�����k޻yK}~�� m�,�J"#��qQ4]+�Mҹ��(��%,�cl�ո��Z��$�[	.e/M����}�jy0���@����@��^���s@��C@��+Y�	$��� s��>Q
dm�,���V���5����cy1d�,�G�[~��/u��<�ՠU�@<�Yo�l�%�I���ڴ
���<�|r+�Sj8�=�Ow}� ��XO��H���䁠yv���vT��W�	���j�ۛ������O&�WI��A�Z��ۍͰ��X�:6�=9׍+<�* ��k��I?R�u�$�J����S����G�I$��Ǡwu��/u��<�ՠU�@���b���!�4�4g���mL
�]`I+��穛�L&(�q���Z^�zw]�ޕ��T�a$� �A4��@�����`[+с��S�?����s��8mcB����`�������CIŅ���1�n�h�]�D�Jc��(=m�c	�W��ݨ�]nL�A'5>n�vɱ9͆w����;��nۓ�M�M�by����.ܳ��n���.��k0OF8۠����s�����뙑���^�;�])�(d8{t�E�b�C�i���ڍZ��z9���ƌ�C%,�*k�c�:�N!9=����k6P�U�3�<Ƕ-�/Y��I}��%�'BM�h3S���#gŲ�'tS���o�ez0>�j`U�� ���Ȓ/��(�4z�4+�h{���w4��a?7!	�QI�}v�������`[+с$���	q9�n-�z����}�Q�y]�@���G��I$�����W�ִ0>�j`U�� ��?x���\dj�;��#�n�ům�4�ڃrsvu�zt�ʵ�~Z��nK˺�21K�ϲ��� s�u�%�A�ذ��#�y0��NFhWj��331"��XJ�l�F�ua�z4�IҎ-�z����g�ľ����=����:�h�(LE�H�J�l�F�mL
�]`X��r,QLr$�I3@��f��v��mzw]�����ӓR1F�k���mu��G[q�ˬ�:8�k�z[�oZy4a���,�Q9�y]�@��^���s@��f���v(BG�[��&]n�$���^��ژ޸��<�#�ƙzw]��������~hɭ�;w$�u�@����1���dm�&hۺ0>�j`U�����z��naUE���M�р~�npP�����[��m�����."x��[a�ۨ�(g��N6��E�����3R�rS.둣XI#K�Ҏ-�mz��s@��f��;V��j��S&�Ƚ�`t���^��ژu��<���s"�L�$�I3@��f��v��mzw]� ��XO�8�0�"'#4+�h{k�;��h~��u�weء	iH�)�@��V���s@��f��v��zc�eds+k���hTvNK���%�:��%��;;����(��Ƭr\LOV��������~v�m����Z��Z��OѴdc#n)3@���@�V�}}V���s@�rS$��S��3@�S�ʘJ�l�F���������14��@���@�빠_m�hWj�=�Z?�1I�j6��-I^0/m�`}v������,�����.ꇪ� �]%]#����������kup0���r�n,\�mJ��{-�y�₼�nq�.�$��]�q��Z;yۛ�%�س�9��)t,˝��p\�c2;��M��`��n.���$�˷'��]ьp���PjMNv�.�T\�`!�iz�kv91WR3���!A#���Ϟ��m�c��!�Û;�[�6Y*�Bf����5g�GY���̶�"ج]�SmcR]��"�U������vV��T�܌Tk�z��8���o����&�mL�*`I+�S%����I���Ԙ�+�h{���w4��@���$q��1H�Z].�$���ˉ���S�����#�q51�G�wu��/��-��Z^�z��9���4�ۊL�/O\]�0*�u�$�T\W��7\݉��\�NrVE�4�βt�uRzGB4����n)�^�S헋������mL
�]`I+����}uaDf
F6�qh{��~���~��a
�P��Q0�ǋ ����?:npk�P� ��EY�@�빠_y�a�L���p�}X�컹-]�v�4�)&hޗ��Z^�z~��V߼��j���̒9�Q�@��WK�	%x��+�e�tN4��U�GK��{�&kxu�ۗ��3�ح���u��z����s1�S6�N�XJ�zV�ژe����]Y5r]�]]`��gB�J&N����W�^�oEq��4�۹�X��� ����D(��
f}���8�Ǔ	�9&L�<�j`U��I^0/K�K�<�1O�q��Z^���y]�@����iDc�!�D��rr�A�vJ޲g���Gl�$�Ug:ɝ�)�)�LQ5�8��y]�@�ޯ@<���"C��#Ib�c�����S��XJ���Ց�2F�DG&L�<�ՠU�W�wu��/�ss@��]jG	&H�ĥ�\�}���x���01FDRH4�H�#�]��0a�@"#��B�B�K�����kS�]қ.j�(��XJ�e��ژu�����}�Mgf�Eў�V?��>\�6r�����9pV�.���p�r)q��A�����}�,�� s���B_�}� �˲*�IE���UYk ��������`Yh�����۾�"q��Z^���y]�@�e#LS$��Q�G�t���S��mL
�]`X�����D�%�I������Z^�X�X��f��D�B�"""BR)`�ЅjZ֐��i1).�2@0���̤˥r��P%����Xb��	0F ���� @����"@�Z�$)oc�b�`@HX��m�l#�$��apj�0
�(H�5�\/ "2�ChF�(Z%HV��� �s`���
�JƤhR�XL��-��dA�BXѕ�FRR+R�#��n�,bE�c�P��l���H 6Gd�P�)8	@���4[ �0�+%*U"�h���iJ~@B��p8f�V�����6	U�h����J0�+
�� ?;H͏eDJI��,�]����N������
Č̡��o�>��矁|��M��ܻ�@�UTiz�:ps�3�v7�"���k�փ2@UR�);L� ���\K+Uҗ<��(ٮѷc��hŃ^m�7�M	 A������μ9rhQ�[s�m�M�btWF�[�.Ɍ6�md�6ͪ��\z�9�g���;�V�d9���w����ѫxx�SB<.ć=����kq��S�逶X�F���s�z�z:�20�f�T���WK�Y�]��q��q��uۊ����.���,�@��w:nfe���z8�����VSx�g��F.zȹ�;g�M���t'N��`�n�Qɥ�P�����tr2�ƻ2��mjݠ���A0Z3���v�vJ�=��ͼ����\��.:��\���w9S�C��ԝ�HQ�r�0y���BۓڇY���<���a�AK-�����wn�d�Kq��bu�fj`&��]�d�p�(+�ɤ䛍�Q9x�u�K	��s]�]�, ��,%�H��͖0��7= �jz�T�O.{�=*jt��@���a��Q� ��j�����`��V�Y�h�[+ ەns��֋V�[2 	V�n�=Ӟ�=-�_!>lq�|�C�5vݲ�Ӊ�-���$�@u]\.B<� t�X�=vB�t������k�^�%�gU����G�?܎ö�Wǵ�I�	P�/\�d���Xq��z%{uc��ݱhMW#`���᣷;���/`툖��#e��"\��2�pU�Jʀ�[����jNؑ�]'ڷu�MՌ��0t��W��GZ����Vp�lq�Qe;)��l�/A�x�pi���vB.�=���m����|��n
��X�4%:��el���g3�5��^|XMkq`�<n��O�D$�D܇F��ݹ�y�dЁ(���o�>s�~vf�9��q���9gp��y�D��&ٶ�t��ML�� s�<3�5e�:�6Č�<�]Q��(�c9N(%��ӴƳ��V'F�*7l�+�6U�rS5!�]]M5���D���1Q�"uC�?
|o鯦Iu�N���b_�v�w
Zy֗J��3�q�2�n6x�n;[m��֛�8���d8x�.��Ьp����3G<��K͋�om�nY���[jgl�}�.x�O\�X]�B���8q����Kڰv[���qh��ʯ6��r�^ګ��ݱu@�ܨtW.�k��n�cq�V4��s���{b������mQ&eT^���.��w{�Ǧ�un�-�=pZ'��N�z��녗��ȯ`ݛ�f���[�5�'1���Q8�P/���
����w4m[����N9��,�������ϒI%26���8�+�hި�F�@�2Ld���q`[1a�3���:w����Ȫ��0�����\��<�ՠU�@�빠_n]����a0���d�붦]n�$���q�밫������<q�%v����s�T�X�i�6����g']�mL�4ζ��6׶���W�%`��������2I�E�8���f~����H=��0�78�79�"�{���ڗ�RD�)&h[����v���Zw]���VFd�j`�Dr@�?:np�np�x�9%<�~y���RF�#�r8��h�w4�t4+�hu��m����)�糳=f��PU7l�˸���7�]g��z�,Zr�Dq7�q�c$�@�빠^뛚�ڴ
����U#L��	M�ﱁd����S��XJ���
��x���9�Yp��kF��?{=�9�u��IDD��C�����,�YZ����QŠU�@�빠_z�hv/l���#�)�D(�-^[�`wOg��tx��m��WK���n���Ϝ�./F�b��ӝ�=\�����^6���fԤE֧�<;j9���8�c��]�0*�u�$�]]Y1�E"CQI3@�V�W�^���s@����=��[���&$�~L
�]`I+��^0>�j`Kj5��<��c�$�@�빠_m��?:npDP$$�P��*+u� ��Q6㑠q��h�w4+�hwW�wu��/����q<S�L�%�Kk�s�3�ۍ�dtXZۮ��}�cR2�������q��M8�(ۓ<ߟ�-������β���Ġ7�R�p;���
&F�b�;{�`�78{eq�$$���MF��;��h޻��ڴ^���u�4~��$�{����`}v�������`yZ��$�b��I��ڴ>n��x���`��Z�5jtMzp���e1���v8�����K,u��4��sKmi�s�ln�M�6-:�.�c�ݶ�tW89�շL9h8���g�ùŎx�ݔ�Ug�/���i��ɡNõ��J��i�ʮ�Y]��m� �S<�]V�y�b��[F����Ϭ�`�>gl�s�m�[��ҷ ]b⋭��GZ�1�	
3��-�[r�6�na^Uۧt�nN�V�_�{��{��G�y]O,����i���;��	֓ o1�\���:6�6E)Յ�#�i51F91'#��>W���x�=x��	G�uwN���WUJ�Wuu4]]`��g(I)�y�,�]��9{k�-|�&(��#@���:����S.�XJ�z�y��N$��I$���Z/mzw]���s@�l�dȰs���QŠE��I^0:����S�g�������V��Ps�>B���y*9�I}�[�r5�)Zku�ϧ\i�Ig�Ē�`u��붦R�`R_y<X��9"K�4o]͙��g�+�h�����rJ!L���rQwwv���/{��~�ߓ.�XJ��]���u��Q�D'�@��@�׋ �׋�DO��� ��L���Q�⑦G���s@����<�ՠr�נ}��q��	��rdɓ1,!�F.Ղ���*ή��l�ӛ�ݮЈ�~ϓ>f��4I� �ۚ��Z/mz��s@�ܻ����&��f��Ss�B���u`�b�<�������!9�MLM(��9{k�=?��31f~^޻���Z�����R�UM�]`�x�=x��M�(��}��@=��H�,s��$�&h�^0>�j`E��I^0$����g���J鋡OO&.�!7kx��.i3��-�<���ڼ�]��I�f�(w�O�ژu���W���`Y2�-	��
F��9{k�=4�����%�K�Ԓ^�Tx�LN�F�7���%&׉����������Iv�߯��ߴ}`'��ٚn>��{�>���s�����ٻm���{���WB��y����m��Ӽ2k35��5��g��K��CI%����$��^&�K��9�m�(%=&�[�5���Ѭ�35k3j�ku�='����mg��v�&.ֻt�u��ȱ)��6�q$������Iw;��$�����%�Q�$��k��MI&�7W�}�|�Rmx�I.���|�]}ZI.�Z��$��Y�s29K������<�$���5/��������J���Ԓ^X�X�I1D)$�<I/l�$��Z��$���4�]e�>�$��t�&&5"��jI.�Z��$��v]�m�߻Ü����wf�� �������y���B�TDj�çe���fQ�ɚx�[���;Ʋr���m�7T�3�f���ϋ���CvcA����n@v���z��R�1K�[��_�]��۔9�i�-yݴ�����ٷhnm"m�y[�2s��!�d�Y�Vu������+��fb*�<n�9��!)��ݒH竮�k1�HX�/m$ZT����Tlg����{v>u��'p'\�G6ͻn��&sѱ�ڬ��n����V*%�+�b+,���?o牤��/���K�׉����W�$�Wq%G$�$rH�I%���x�]v�M$�w�_|����4�W�>�=��n4����<I/l��I%���%���Ԓ^�o��K�͋�)��&�s�����o�/<I+gڍI%���x���������������}p�ʗ	-�|�Rz�1$���>�$���4�]�ns����wD�xe�M]SE֥ԗ]R=:.�􎷯Sj�bb9����ih�F���<̎F��$��I.��<�$���5$���_�$�s��RI/)�����ue�kG9m������)��A&3MJlw~�$���4�]���|�UL�	��D'��$�~���$���M$�Y~ϾI.��i$�J����o�y{=���o�$��^&�K�߳�K�l5$���_�$�Y�%G�H�I%�o���%ֶ$�o[�|�Rm|| Ϧ��q�n�un���gsx�d�G'\m����'z7Hf�V��&�mz�3� �q��Ē�˨Ԓ^�-^x�]��PP�e�������n�kV�֭�h�/o��Iwz���%&׉�����Ē�˨Ԓ]n֡�� D���ng9m�}��wm�����9q��$B	�eM��)0����9 ��
ZJU��g�8�FqM�F0��Ft#�$� 0H���*F(H`���6�F2A$]IĐ(��`4" ;W�P���H$I�~ �H2A�AF1D� FjH21 @� ��B��]  ��D�
iR����>D_�S�UD? � �<@O� k�~�v]�m���s��IS��xH~�F��$ũ$���3�K��CI%����!)=ZI%�&���$nj!9&y�I{]�jI/_��<I)6�M$�u�g�!"����KR^�{�0��Y�`�3��V8n�� .x�6��N�����է	��WM����>�?)=ZI.�~����IO���i$�����N�dm��$�t��I%���x����5$���_�$�Y�(Ӎ�`o����4�]���|�]}ZI.޷~�$���Z�J�i�����)���g�$�_V��K��߾I)6�M$g����x�]�nn�q14��Ԓ^�m߾I)6�M$�u�g�$�_V��JȾwލ�d�L��@
j����l�-vޫ]���[��Y����Vm�uv��On�~�$���4�]���|�]}ZI.~���$��YXH~�F��$ũ$��~ϾI.��$�o[�|�Rmx�I/�Nv~rLn$�BrL�Ē�˨Ԓ^�[�|�Rmx�I.�~ϾI*�V{E���ĜR����k�Ē�wQ�$���3�K�f�IwuG���pS#{����II������~��ܒS��<I_������qA��T ,�Uh��@�������Y�fj��]��&�q���x��m�s[�GWnk7d׮�,�[.��o��\���"ݥL\�q���*krW+/Zv���������5g�:� �pۮT�q���s< ���4��[t��M�V�S��ڶN�V�u���XRe62��28���`]랬R9�68��ȸ��/�u�������v�'="'3]����@x��ͳ�a��}��uo��O�."D$4]uT�>���,劗�f�d��Y�x+t=:�8n�OdR�/#��L_$��_�3�K�wpԒ^�m~x�]��5$��������s}��%���\��`I��u��]?<��II���^���Z�۹�{m��9u���HF�-^���$�S�׌��`wm���Y�C��cFE�{��׌�0$�S�*�'����{�M��[�j6�Rļ���&����{6�4�Ue�����7'�$��MD'$��n��ՠw;V���h�lmLq�h�5u�rO߳�����Q #�T���N �݋ �o��LWj��.׳۾��0$�S��mx�����F��$��
9$Z��܀u�����wl��:��7ۋwCئG$s4m��/mzs�h޻���.4�dA��y�a֭ml�vr�.8�[���voFu�`��빭ۜk#�R^�0"�u�&ژex��n���G���bj7���ZY^0:��[��%��������T����<���<�ņF(�Y	@� �B ��o��7$���n䜳������5��4m��/mzs�h޻�{-i����ĜRc.�Xm���W���`\�����ƶlFwj�ע2"�� �,��/�1��ˡ'$���b.%�Xm���W�����
�������ϡ�FL�-��s@�۹�r�נw;V�}��CPM���G$�c��u���mL��`IU��mI�lM%&h����ՠy�Ł�XB��*��,g͗pUȤ���zs�h޻��������X
�_�?6��5�
q�Nv���؇�)��h���"kH�77n��م�)~���	"�=�w4m��/mzs�h"���I!#�RI��׌��`I��Y^02�Z��b�ܘ��L�9{k�;��@����=��h�Tn86�LQL����;����W���`E��Y�Ysǖ���
9$Z����s@��B}�w�rL�@��U��:^�m�<^C��m��cl�K�]=ۆ� 8݊���;f�Rv�#v8�ku�� ^��N[Y�,�hǃ���1��<����B��v2G�۞�|�π��|�f3�@�^ccs��[\�-b��#�/Q63E5�}����:.��f�^�M�Қ�;�Mo	���z����bmWC�Z�{g�NJ��5m�璃��N��^��v���1n�{8����Z��|�{������ג��ٳzɅ�Wt�6%,������pj�^?>|�3qdM<&D)$�8���9{k�;��@����;��~q6��D�4��`>n�舅27]Ӏo>ŀy��@�u���$Ȥ���zs�h޻��������N�&�k�����`u����u���mZ��;1��H��%#��{m��"�u�&ژex��.�j�����7�t[qŨ��ű�u�����☔7V�U5=���e1r��6������	6���+�[^0:J���uo�nnʩ���7i���
(QTm[ŀ{m��9{k�:�k.2cY1�B�I���+�[^0"�u�&ژ�70���LP�L�=��h�k�;��@�s@��&�90��iM��=:�`�$��O�5�b�<���m����a~�sg'[�=@�-�h� �� ൹����l�\��X�nr~�џS�h��Q�����@����=��h���*u�D��H�XI��[���ɽ݋ �}Հn�s��L����T)pCS$��w�}��z��E���~��ms�h��h쵬i�'�ɓ7sv�:)�������7[Ł�(�]��y��~F��8�Fڑ����$�}ߗ�7��`��`�M���v�h��\n���.[v��������<u;�j�5�]|����7����k��M����ŀy�� ��� ݦ� ~�d�RL�E��.�`m���(_%	U~���;�� �o��଺�"��i)3@�[^���Z}����[�ۚ}�ۚz�pƚ�"�@j'�(P�����X�x�2"�I0`~U? 	n���䟯��D8������-����������3�9}��@�v���3X�XLQL'U՛��v<�S�h�m��y�ks��8��{IpN�"<Q&G&18����$��n��m��M�BQ��ŀ�uJ����*n���ݬ�۬�}
"��￿�4�l�<���Ș���#LRV�M���,9BQ	L��׀l�uhz55��(�h~����}�����=-���BP�����hJ`L�R)&h���=Vנo���7[ŀ8�P�!��JH`$?��E:?��P�>`�$6������IE�T�����%� �F D)��|8!���f�42�\���Fd�Ni_�D�a��	�$!#"Prq$c��XFƭ!BH��D�D�J��6�A�5531� D� ��R��9��@��`Ȓ$bly�L"�&1�CC�X~b<E"8�+D�$!4<`�#����$�A��� ��D��,��0	�"@���ј 4@D6�:��@t1`��$��t#w���əu�fj�u�L����`��f�:qώ'˷u������;5��3J�����ۭ'L��m���#]��E@p�g�
@ z�:�-BI�=�yd狄�uvMڶ���n��7h:����E	$�B�k#It�4�ʨm#��^U|�d��2N�"�D��K�]�RZ�k[:�h�ȹ\�^��]:��ä8�� ��oh7�`Ӵ��y ck��	�=��cMu��C=�NK:K*��$��$�u��Y�M�:��Q;����4�؋#˻X8�o8�Qղ�hz��:�|hj��x��!�x'S���'!��Ej��v�����c`�tNv��c K<��;v��涵�皀���ڭ9��n��q	��ز�7
�#Y�Ig�8��-]ul�)Vʢ��Ez����e�;��vC���^՞q�^P�j�!a�u��8	��q�;O<w9X�ηpf�k�x͋�'������cpD�x�+c.^61g�j{*Q�@v\�$�7��n]MH�uݢg^�)���.��m�wV�{a׹6���O[ʴ���L�9r�gVݶwgN�(�y�ս!{�s���Wl6�K\ZUC�7Qw`���Ni�B�npHck���8D�c��l�n��d7�j����g����tٱ��l���;�_HNN�A`�mֶGI�#�U �]m�cu ���]�;1���	�s��e�˪�P���]vL�Y�[m%�P[R�G'm�=PP;���7S�e��sq�����P���SEm����a�"r��@����s�v��&���b�	�n
��Ci��:��2M��WV�-�l��=c�&��&�������Z�qe]�#T��m�r:��86�4����,�ݥ�9�m���y�A4p�;nF��&�웞gs�]�+Okd���5�]e��;M���+`���0��mNѰZ���xU6:�3�WT�O:����n����On�wa%�v�3�ik��Vڛ�i5sSFjMִd�ՠ�؄PD�Pz �j� ��Ң��w|���2&?��˲���O<�f,p�u��k}5ҲU�v=zN13jL��I��j�o�nyWVi7#���ָ\�p��i��7HOm��='G;g ���nF�hf+"I+����z���=evq�s�ۈ`����*��s%�ns���K�ęj��v��ۧ���t���R�b9���'hn���ƹ4.�5mr�ţ��l�;���T���BpX��^��c�N���d6.[����Ҳ�����w{���|���c��׀s�� ݦ� �o(��@�� ����cMI����@�v���X�����gB������ܕs7_�q���-߾��m�@=���ڴ�[&1����$���~[�ߖ ow^�M�(R�w��sIF�22LJE&h�٠w;V���,ͼX�gN@L��왺���sQ��GnN�����b�����n*�kՏ�{�f�&70q��jI�|�����n��s@=����Q
b����7[ś	�$�$�";0��ذ��x�79�BJd�}�*UL�jKE)���X�v, �n��np��h�]2F�$�H�4����f��M���,�{���}=`��jʟ%�R^�&�j`Ik�[^0:�@�ޘU؂C&'�S���=m`�;�t�p��f��t�ZvɚTf%�\ܒ���u�X�x�7l�"ޠ���������14�I��$��k�[�0$�SK^02�Ixr�I�H���e4�j�s����18!�$%4�D%��x���`���sj��E]U��������� �����=��h�)�[n���ncS��{�L	-x��k�[�0$�S�oϿ��ɒn�b;�Ekcr7`��k��ע���j�8ke��t��h8�4�]����c��o���mL	-y�wUt�<I9�<M%&h�)�n�s�n�� �o|�DL�/��UMYSs6$ݘu�8�x�舄��}�ۚ}���<T�"Id$h���� �o��,��0.!r���p*� ��w��w$��}�i��
FLH�f��s@��M�ڴ��`�$���(�5S6�-UT�ͪ��\���h�u�G/��9�@ðݻsF����G�.�����H�"s=�O�@�v�����n��]"���7�p�7i�Ϣ"">UGw�b��}� �v��+9�̑�8�h��h��a�3��� �wN ��&d���S6��E$��n��s�h}�������B��S3V��QSv�7l�7i��7[ŀy�ŀ\G�Q�
�t�㟣!	�:��f�b�v�:��TH��D�2<my�c	{<��s�J筢�c��of!�-�;Y�fa:��Gk��6��ϧ�R^-�4n���9����vl�nk$�V�wc�r�ɰcǤe�D������ׯ0P���s�l����)z��h���0/�ku�/j4�-��u�s�m��xk��P�q�X�sZ���JR\r���f��f��$K��n�1�T�;p�X��O�P*�`�w6�p���7X��"WF�`�o�������7[ŀy��������9�ꯊ����%Z�]����ϔDL�ϱ`�|`�ns�J&C�w]�&�6��S%ݬ{�����b&v[��׋ <�B�j)QJh�V�!O�7�`w�������t+<��o�-����U��7i��9BQ�����v,�m��-�RB	8�rcrF���?-��m��=���uY��x+v�ճ���.I���kW%]]���7_b�<�ŀ~�x��
_Ģ#���Ӏw��L��K��m�����y��7D*���b�?m78��rQ	L��3|
�fUZ��EM��7��`I����`u���wi��ɔ]�2MفД(���8}ذ>����h��ǑƗ� �b�H���`������|`�np�9SR�h�Hdx8�"'����C��b<��n�;�l0W��c�i�i������wk �׋ �v�}M�BP��~�s@>���%#Y2D'��{l���� �׋ �׋>P�BK��Qo��Ȧ2H��(����-���&"DD$�����<ݳ o^T�]��Z��������R��� �}� �l���b�>�hu�R��)���ݬ�^,�=ݜ~�wN���}���kHG#���k���m�GC�;����^��7aۋ�Vd+neۚ�<c�f�岚z�Zw]ϳ�x���nh.��?�Ė1!Hh�g�)��ذ�ذΛ�䒄��T9��wtLU�ʵ(���;��X�����Zz�Z�-���L���J�X�N��� �Wt�>n�%������/��vZ�Lq��$Bq���78BN��� �v,�^, ��}QYyJc9:-���e�匂����[v5�7&�ѣ�6ݖD�����ֈkQU7s�l���7[ŀy��В�!�]��>���2dǍ�q7$zu����X�78ϛ�����BUGϾĘ�"S�h������Z(���s�Հ7݋ m�ӑU���UҢ��`|�"w��p;�X�x�>Q�N��� �}]pUW3(��d���6|�`�G�w}���wذ:nsm���w���������:Γ�J���1�Y�\���OE��u�מ�;�v�sVٍA�m�4Q�*��`��x�5Ę4�6x����Iq�a��7U�֍�.�o'��+\c�w���^����2j�^0����YR���.��Ŷ[O&���c%�SD]&������9۳�k�Gb��uƥ�q��:�1��<��,�c+4��W�����ζ�����b���Q�+;��lt�+���vN��:_�6���H7]jzy��IOU�Δ뎊�o��ŀy�ŀy�s��� ��j��RZ���2]��<��ϡBJdޮ���u`��ϡB��滪nh��P#Bq��|��h�����h޻���t�2D�&ԋ@�� �o�D(�޾��;�eM��Q7$zu������v���� ���G�L���#�Loknz�6��q���#h� ���u8"�X��[������x�dm���9������=�ՠr�נw[��[Tu�dP�ǌ�f��?w;ۿ�B�H(�z!B�.w����`z�g�B�:_W_�I�dQ�ŠU�|��w4���Ļ����?�Z�����F�LJ����`z�`t��}	B_$�W[������EU�-\�Z�.�`z�`D$�z���w����`�i�#��o����g��$^:��&��J������b����z�u� Kb4�o�}�?o�Ɂ[�	-x��+���t�2a �&F܋@��~���&F��`ϱ`t���ʚ.�S5j�K����u�X��Xz#ЕD$�(mbDаR@Ї�ZU��j�X#]��"�	!A$b�H1�P�Fʪ1N`� u�6�S�<tiq)��C�bŢ�WD6`�Q�J%���P`�/^	�T:(8~T@�,]��S�O����]�9{�s ~�r*�,���U�eլ����}�h���r�נw[��[Tu�w7Juk �� �/�$�[�����,�^,��aT�.�]U�M�-�c��#�%�����Amru�Fg�A5���n9?�LJ
!�8�^����\�D~��Wt�/���ݪ�Eѧ�g���	%x��+��mL��ΈQ
d=�u�L܊ຫS%ݬy�x���[�	%x�,�u[�Z��j�`t(I)�_t�w�����7$����z
��?�~��Ѩ�!26�Z/mzw]��^,�� �!'�9����E���u��G��GkJu��O-<��6�ݹ�F��Gi��������{�����nL71�j�o��������`}v��������G�j��wSsuk �׋9D$�ɽ��W}��;���;�u��"��hb�k �� ��u�D$�e��X��Z][���6�H�-���߳}�X}ذ=x�>��Q;��8���wtJ��ԫ���7[ŀ|��Ky�����g���BZ�Zk�MEۄs�Lj���!ˣ���؀�t�4Y�@t$��= v�ecTy�l�ctn]�nI�M�,�v;�ے޷�˸��:'bܹ����I��Y� 'g;�Z��}H��֣ n;BY��j.���Q����X�GN��Т�[:��nilf���� LAիb����p�rXk9����;�j1�b�:7T�F���ۮې�
l[I����'�p�k����+m��5bkюu���U��7�]y��+�0N��{����6O�D@�71"I������<�ՠr�נwu��*�(�Y?)�!o�}��ژu���W����=���w{ܻ������+]-[���{� �׋ �o��f �ySE]M�7%�U��(��[}�`�ذ-��9u�@�����Q4D
�`m��9%��? ��V���zP츓��a����$�����峄Ŏ��ٴ��p�y�ve�Qv���GKj4K���������W����*��F&I1�F�B��9u�n5^ ��	��{�ٹ'~��nI��z�Uc���21�E#�;��hm�áB�3��������w4��F�$I3@�۹�y]�@�ֽ��)m��t��r]M���D��Z�?:np�>��o�`m��=���޴�5�vd������[X���ζƻN�穸S;^�:b9)J�J��:�`��`m��(�!���>�ﵦ`70���#�;��h�q`�78�79�
d�vr�����"(���w�}��y]�Og��sv�����e�c��Ț���S����t���`|�N��� ��7�����#I�8��ڴ�2�ߗ�7�b�?:np��-׈��iV6��G��G���������,��z�z�*�<L�l����ŏ��8N����߿����`|�������%����QeՄ�Wk �׋:"������t���gД(�k���j�L�Ԣj�`��}M�DL���_�4{���H�mHL�9�޻V�}�vnI��wf����AC����M���O��s�dD�I����o>������7����2�[�&\���"�/�{g:��1ㆸ����������&8I�"b�m(��pRf��빠~��`�n~_%���`�}�J�O$����9�����ڴ=x��GB����x�h�UMU`Y��&���>�0?+n�9J���md�&,$�@�빠{z�h*�`r��{}Ӏzz_]���QeՄ�^�0:����vژJ���j��g{0÷D��3.�&k5qۤX�8���G;I:��=��R:0������&���I��ݹ�lq���`�'Z��n��#�o'Y�ʞv�F籹;m�1�.�P�O�q4��;���dU�:�"7F��&�#ѷn�yY��`6���OV�뭮 ��s�,c[�uj�o;;�r��܇�nt�{�ݺ�����ʤ�
,*���Tk���q	����O���En6�sM�&�G��=�j��X�ÕP0�z�5�U�!�o�����?��ґ�NG3�;���@�]�@�s@�۹�y�MM)"J8�r-��8�x�6�`t��B��d���+2	�4H�h����sO�ٙ��~K�|�_�-�и���j2)5eլJ>Q	%O�����Ӏn�s�w[��w[�Y"y$�9X���u�SM�0$����/��v�\��@Y�,�d�t[�WHZ�y��L��
���[����w���3�ny�E���|���`Ik�[^0:��Y"Y ɋ	"�;����3�\�Q
�w݋ ޮ��7i��?K�w?69��p$��{m��=�ՠw;V��n��ܱ���"F�8���DD}����}����Ӏn�� �ws@󺆸��(�dmȴ�j�>��	/�!BK�＼��`t�������k�[��V���~�`��d�Z��=����g#<�S��xk&����~x��+�]�0"�u�zB��%���'�h޻����~������U�|��w4�v!#�IX���{]�@�]�G���33 ���AQ�O
�
�K=���,�}� s���J�T��ꑨ��0'm��%�ex�붦��dD��y ɋ"����h�!$�ДDC��������6|�`�q�їvέ�Nn��{���I�^^�۷C��q�kf���@-��[C�L�8�-���^,Λ�g��%	D~�o�U��?�8�N�L�=�ՠr�� �o��,�(��O7��s5j��n�WUWs�9}Հn���D%;�ۚ|��h�X�?7 �#rG�n�� �o�M��J!%J!$��$�\����Ҫd��7%M�Y{�`u���ژKu�%�w����9y�uP۳n����O<�/%��*�qt�d��1�7#g�ڴMc����J)���y�s�l�u�n����K���ۚ����8��)��8�]m`���<�ŀy�s��DD)���="$���LY�@��4m���ڴ]k�<Uu��`�d�C�0>I(���� ޮ��6u���BP�So�y�W���D�q80N)3@��g ��� �o��,�$�B�'��B�T�b�kgm��H� Z�@�
����C�4$�kHm�B��)@E��CF��R��B	!��bF�H-"�"��F�icL�"�N^#�"�$x�*�2<x!�Da!Q(B�@�Q�D�T�����r��V,4듵h���2��j���a��p����Um%��̼-����*�)ut��G�2`��R�T�U&L⹞��t]v="㍁SG#���Rk��w;\F�^x�tY����.t�3K۰c'b�.ôj���Mؠ������c$n�ᖞ[���e�N^���9v���fn$�Ў[��$9��I[���H�i�n݂�NFJ���\c�5λg-�m���[��Zu�l�mQ[�¤	��v�evÄ	���l-;Jf}!�������O⨰�ڞra;i��"���/Kb�=kT�0<�̷X�Y�eZ�v2$�K��&���:����Վ�0��@3��!G,�Ũ��Y�g��v#=; ��hJۀeP�;X��PR�[�ge�e਱21�
�v�j`��ƨx�C$%%�݆�C�AۄG��֠�c9^1����u��M��wnAܾ;g�ѧ`=�'�mo$WV�v�=
8�:����7<�x�;�+[q4\;ns�{{SC�9
�'�����&m��7mc8�J�+�j��+RP�h��w��m'-�9�P&�U	[n'��[n���H��`��9"�cy��s��$ ��m�>@zS�۵��Ömy�lHc�.��m�J�@��6lp�sV���+�Q;�yU�Ğ�r!Zr��'t�;ݐ��.�s��l�n8�-�lk�1���eU�e�7#���6L��l��]v�r���Š���ns��ܺF���۶R�*6в���b�95Aĳ��] �&w��ۧg'7-�]�ݞ�5�9FO�m���s'�ج��A��lrn^��m�TХ�l���/�웴�չ��vE�tJ�q[Ӭ���8��KZ#�(XS�rŬvQ��­5<���n�S�[�nn���c���tn5�z�t&熳׌�a�,�ЏPQ�u��-j�YV�В�ģZ`��VIu�F����5܋�U�Ŵ8Xh]N)n1qr��9��\��9;�!;:YZMd4�ML�e֮� �Qh��P㈿�DtPO�x(��"��#�uO�Qvo���I�j�,�"��,lrY��MyԞ<l;���ո��Kj�K�ݎ"�g�f�{�)d�VyGb��+m��r��x�λWX�7i3��;wk�쇎����3��Y��[��F��.��c[T`��`ë�i��n��{p�r�]��נ�
��CAʹ�l^;ۓg��t�����j�q iŲZ۞�x|�Y���1�C8��ͳ���w{�=(�9͛��������A×���m��%����Ga�xh��ՙv��r(�R.�����h�w>��""�!�]Ӏwu������������7[ŀy�� �� ���:"",H���E�D�!��#��w�}��{]�@�ֽ����׸�F㉥*�Lݬ�DB�����u�X(P�%<��,��WJ����mMI��`U-���`Yk�]�0>�v���q���V�J[Gl�h�+Ή���;n'�1n�تU��]��s�������f�Һ(�*�� �v,�x�k�|�Q�K����wH�J��&J�X��dB��D)������ ���?�?f~��_���G����I�_��`U-�K^0,���|��&8H894
�נ{��h����Q	D���u�T��U�ԗuWwL��`Yk�M�0*���Y�/���i��MtW.�u��Q>�FNɁ�k�zn��N���,��|����w�??7Ó��ђ'�p����nh���u�@����;�{�LQ�6����ֽηX��X�l΅�������*mvM�������V��,."Ј@�Ei�U!`����f䜭�@�uVDH4̈�őH��q`]� �����Т+�ﾬg�}�'��s29!ɚ�)�z��@��zu��{ե��7n~J^x��]��4[x�kY�77�3ۮ�,�v�߽كٛ5Q����;���@��zu���)�y�U��Q�8��ԋ@��zu���)�{]�~��~�|�4���M7z�}��{]��%3�]Ӏ9}Հ~{c�+D܄DQ8G3@��M��Z.��_��{���rO{�͔��)��]fQ-��붦R�`Ik�[�0/��0�xz^Ζ�a��|u��Ʈ��{R���d��ڸ���!�6�e��vk�o�M�0$����]�0<��D�M��1a$Zw]����#{���]Ӏn�s��DL����q4����ə��X�_�M��%2���[�ۚ{:��'2A�@N)1��mL	6���׌��`}Ҧ��HHԘڑh�ՠ}��3��}ÒO��lܓ�s���
��H��ܓ���ə5�rԳ2�5�n2gg���q]�gn)�.�������c�b�p���v��d�6�tݛN�E��Mk��zyu�g��_�=�ɟ����[�6;b���ĝ�����)�lq����l��$C�m�n6p��fd������G=��>�<e���WO<u�玗q:8�7)u[��|���:�m�3&E��r1����u��w��GG,�bK:��$���M�]׶��&N�3��p��_>.����55G�����x��k�]�0$�S��V�(���'�h�w4k�h�ՠw[��wZ�!�s&�Ĥ�۶��j`Ik�[^0*�mZ�J	H&&���;��@�s@��M��Z��ȇ��1a$Z��`u���ژm��$�$�C�k\\ɫ7o�k�.�X�vo�{n��>3Eל���(�5q��� 5�6:�Q��mL	6���׌̗7(��vQsa5sV`t��%�
!$�;V�o]��e4=�6�HԘڑh�ՠw[��{l���v����!�26F�h��hg��붦�0/Oa�b�"J(�#��{zS@�[^�޻V��n�zP��$k�$�F�((��z�wU�-��*8�z��m�Rfyȷb��[ٻh�4^��]�0'm��%�vU�U�:�M(% ���Ǡw�տؑ��4���z�נy],�y�.l�(���=���<ݳX������z���k��[&!�q~�@H�{o���-��j`t�� ��19��q8h�j�;��@�s@��R�<��B��1LLJسN���:n��X1r�t7<���P��v�qD�n`9"�cJE�w�ՠw[��{l�h�j�-�<�D�L�����7[Ş_Ī���z�� �W���߿g�ċ�B�
"$���9�����$�붦�0$��Ku��d`�f�����D}��������'�w�7'T@�O��	 `	UQ��$SV�[�rNߪu4�PJA14)�v����ͼ� �v��[�]EP�d�:51�mr�7<��wa�xm�=qGc�Ƙg�����7���|k�NzQ�:�G�m����|�[��ژ���>���n���Iɚ�ʖ��;V�޻V��orP�L�4�U
�ի������I�.�������k�[��ji�0$�I����;�j�=�w47ng�DDN��0�sʑW���F�h����ʖ��YM�v� ����`̂�̍�ċp9����u��kn��l��f�[�F�;w��9te7qk����F(�YLN3�����<6��Lk<��6�;��C�s�l�8���r��M�!GS�I���e]��4��e[8w'Pr\�����=�z�Φ��oEm��bw6q!����hu�j9�s�O]&��GfA5��)��ΑG��j����q/S����G+m�Q�Z�rݬT��ظ;t�W��mֆt0�]\����[h��կ�ou��������Q	~�߾�s@���?'#Bi��;��vژmx��}R`Ujڵn�ɛ�h���� �Ss�y��ℾQ�U?���;����۫�T�jjʚ/����o�L	��`N�S ��d�Ҏ/�H$��4m�-�D$��
\����9��N����w}�B7k�4γĒ<��b�������z������6�V|����|�.�X����+�[��U����܊L�G�޻V����?d �@ �P8&+�T���v,���8ϛ��BQ2w;�T�?L����$Z}~��=�T��������-�aV���I�(I)�����V��� �׋ ��ƛȌ�	��K@��@�]�@����=�T���ks"������v3# E��ت�+%7 ���~����G���r������~L��`u��0"�u��۾�n����&,$�@����=�T�^���ڷ��H=����S$Y$��rZ�7��g ��u���P��"�,H�"�-hD�>��Y@�D$ED"�$Q"T�s>�d%K����C�'VT�!HQ���a�	��2`B:\%7��H`@�IR�!bVVY��q�G���i��(�Uq���"�Sm�! Ѷ�U��"@�#�!H�!��X�h� ��H�,`���!J�HBq�cR�D�,��t��F�h B$`��H4"�1a!Q�B�Rb0�V�1�$fc���A�kh��
�࿖�X%XՊT#@ ���Ype �_�� � GQ,B��$UE�DWH��]��:�S�Cj)�o��+�+E?��f�5�-�z�h���q<�H�o��&]n�'m��d�~�S���-��#ZI�ɸԙ�=����X��3�9�u�|�%;��3WDM�:Գ9�����ϧ�E�n�ny9�4+ۭ��n�]��+!r֊.{7�����m�߿��X��3�9�u�D/��:���;��a����4m�-�mzz�Z�U�0Kf(��us8�7X���:g��X�_L��'Si�IL��j7����ي���s}� �jp.�^n��7WJ�&乩UhE�� ��X|���)�O���@�]�@=�����C���m�џ˫CU�p���'^��l��4]]5P$MȲI1&ܙ�{_\Z]k�;�j�/[�����m��JF	��:�g(S#���v,ε��?^�׉9�R�5zz�Z�w4k�Z]k�-�X�s��ș�w8�������' s�����@��Ն<K @"#�L�=��h(��}����8��`�0�J��D�6
"Q ������Lw�l2LN!bQI�}���B�e�&:���t=O���8��8�v^�
���ۯb-�6?<���;��^��wnJE�WS͵v�:B�^�i\�hy!۶���IшF.5�c5��<����q�m��" gۃcRv���R��TɺZ8�{6y�,v�`�F�����n{;=�uy������tW��'�CX�m�Y�4{0n9�Ӕ�{��w{M��x����C�ͺq��=nm��:�$:F�!地���{V&+[��F��'@��u�o�������G��U���������6�q��hZ��m�n�9Kwۛ�����V�]��[ŀy�d����}��/?�Z��	r,�LI�&hv�0*��vژJ�u-����pZ^������}oۚ��-�Z+q1���x;c�̴6�:ʆ�O�6�v�����۳F̅gx�ƜNG�q��h��h�h�
�����x82d�,�f�w$��wf�:X*� "*J!�K�If븜��� �Ss�u���% �&h{e�@����J!D��>���X���a3t)�&���(��=[�X�>��]��l�h�'SDL��j75�ݲ���`}��]n�/R��[گG��̅ێ�=�N����9x؞l ۳��K�ٮN�}��wg�|�^m;�B.���,���`|�}��s�- ���B
8"I1&䙠{[d�%�L�;�X���^,�J1 ����pZ]��@�Ss��TB�I
*��ŀy�d����օ$X܎���;�j�=�w4k�Z/mz�+a2GwWs�y�ŀrI$�����9���7���B��d�Rh�V����Wuj�����K<��Hrtk].u��zw\�=�����#�x��"$�L������r�נw�ՠ{z�huV1,��B��	�6|�g�"!%2=���7�b�<�t
�'SDL����zz�ZY^0:�T�u���*���ļ�UhE���DG�(���}�?���p���7'�)� %B� B(:4Cs�k�r{��)&"I1$䙠{l�hߒ�[�_�{]Ӏy�ŀo�䫚���AIq�=y��Ke��&1��:ۣ�ֺ�ˮ3q�.#����~]��<�j�ga�K�*��kvژex��kC��H�8�H��@�]�@����=��4^��zV<L�2Gr�� �׋ �o$���BU]/� �_��_l*�%0Ȃb�I3@����[���`u�� ���<�J�ԖsUw&��� ��N������ ����P�S
1$����5m�h�2�j�.�sW+t�
D5���]��4rk��;u���d�Cvb0޺�!�c�����z�g�g:����e��"�-�ͧ$��hw���5�ݼvNn{I��\��tZ������y�>`DM��Dr�*��zI�ܦ�g����+ף�Y�ɧH�+ִn#ڼc��M��ut����;�8v5�;gn4d�Q5�8�����dζ���q��u��y����_h�[i��r9�1	��l�6nY�RH⵸�PÌ�%��%�����k�׌��09Yu��U}��niM�eZ��`��g�(P�M��F�����9{k�)�F�'?BI1%�{���}R`r��.�X�x�/g\x�$��q�q8���^�ަ� �7��Q���8��YUr��LR9�%#�;�j�;�w4m�-�z��S�D�̊`Ԏa�y�v�!�<���oB�s�\kOn�3���s�>_w��{9!��M�"��}��{m�h�־�I~�{]Ӏse��JfЮB���ݬ�ۙ�X�"��o�`����o3@;��ɉ`��@Q4�U���7Xt%/{�`��N �vi�
�Z�WVUM�]`�
]ou`{�`�h�U��WUc��lQ$�}�	ּ`u�D��e�]n�$��|�ѭqu;Vn�d1��3���z;v�T.��.��u1�m�������_)Nޙ0JI3�;����=^��^���{l�{:�c	$k`��a�z�� ��ݜ�o�ѝ'��YTY7j��]��� ��� ��ŃJ�P��)�P ! A`&�P6"�9w��M��{����x<sd�&�h�^,ͼ� �����B�!*�}8�q?�1��� ��rL�=��4W���0:��qB�I{پ�F�D�HV��ܚ��]6��g�#٭��8���-�C&%�SD܈�9{k�;�j�=�w4m����ш2BA�UM�]`�ns�DL�ϱ`��&��^��Y1�D�ȠaZ���[ZKu�;mL�[�n�^��wV�������{�����X�;۹?�^*H�E?+�pG}�����/���I�	��4]k�'m���W���`vY��un�-�{��MI*%��D��:x^Ga��t��N.cd�^֛������o������ͼX���!/�_u`���Ec�$���@����=�t4WZ��ڴx�i�aLR)&h{m�[�:��^�t���`uV�51N9����^�޻V��[��{m�hun�XDI�=��`N�S��mh`r���Gg�E��l��SA\H%�J�!
�A  8�$#da0�0�K(HD-�X��(Ь!
�R�0B"Kj�Vτ�)�#���֌L�]p���HEi���J�#(B�+)!iHД%-����J!	X�"�eaXV YB�B�RVR1�HA#	B��(6��8���l1 "@
�-P�X��"H%!R����X)R*0%#��W� `�bD�T"8�	�4*S��D"�!,�a%
QK*R�`��9���+��څ�8��eW�<�q��-d�v�v�Z�T9��Ȭ�`�U(U�()�`�5�a�R�T���?�>Oͩ�m`C'mt5�Qv��MT8Tms���k��3�ny�v��=��\k��]���]<ؑ���ܸP�7[l��l�\x��d�s���8���܌��[�(�K����ʝ�Uzvͬ[��s���W=6rN\#�tglmۮ7<�4�ZcQe��ծ¶�u۵v2
�;r���۹�.E�c�6��;b�OϜWEc��T����tN�3�c�x��_���&V5\Z�<S!���&]nu��t�Jʻ.m�E .=��`�[��r��@x�h�bL{Rr\��g�o�����@�r�N7���R�l�e�h3���g��Ct�pS�oi¯/L�%��ע���Cm�5��'N�9�2ݲ��Ѻ�0󭳬�v��p���d�6����;v�ܳ��vǶ��us������l	�C��n�2<lg�#f�T�� ���@�r�K�klf������l�<��;w.��nٺ��XN2(=m7:�Qew�ƷuӎZ��Y͉	͹V%v��r�tB�\�*򀻌N4i+�EK�؞Q̰i6���@���:�CKak3���V�;q�����n���RCb��Ӷ�MG<���v���nޮ���\eƄ�������2�$�Nї\�6�{��Cl��-��{ 
gO]����sH�s�5��a�n�� \ �YM4Jn�m����bvvSZZ��vj��ɗ�w�a'�ҮM�җ�hl��6�3,H��M���Y�X@��8Ք9���8H���af����u���j��y��5��"u�`:��<�[�E;��cZ_[��DM���6�u�m��8�'P�v� K&��P�}�Xz��v�Դ*����^!�pŵ�l[HkN�eZS����,s�%�[��w)m.��mI��n�m��,�Lۖ�j�lq� %P�X�z��hֵ� qU��1E]��PN������F	��+@?~ܓFp�Ia�P�u�5��c&q��y�,<�Rvk<Y�9�kۇ��m�߿����w>=s���V���xm(.�UyK's�v��:^�#��XֶU�{:^iԽ4���yyy3t�y����n6iU�j\b�tVlt���n��<͎ծ�0���sn��6� �ѹk���YӅ�sk.wZ\p�����67gv6n�-�ɶCa�vY~������'��5n���Ok���NN������#�،i�{b�m � W�����#�r���y#������Q�z�נw�ՠR�X��"�`�$���I�zu��7�����g(�J&C�_���r7�<��h��=�v�ĔDL��ŀo>��?y�*�eݖ�s	q��h�����nhd%
"v�u`���EU�任�����=��`(�ϗ��K�}M����>�k[0�rV�f�m�b�8n�<�8z7��nan�x���sg�s\Q��0:ˏ)n�'m���W����X���
'$�ֽ�?o��x��<��f������f䟻����߿$|���X$�q�F��/o�Ɂ�׌��)n�9Z���wRU+�]\�}	$������|��ֽ�v� ���
~�70H�����)n�"�u��׌ϻ����ף.b�����A�D��nr�z�����3x9���smٝ��˹��{M]]� ��u�l���=���/��}���}�)2G�H�@���׌��)n�-��n��任���� ��� ��h�ay"?$�"`CZ����9w��'o�Y�c���I3C�����~Šr�|�^��z�� ��$���	���S�zu��>P���W�5�b�=��-�y�&���0�� �G���\�ژ���T�����D��տ�����1`L�	ƙ��*�z�������9u�@�[\��R$G�@ȝ��}
Jd�w���ug�I
bX�Ͻ��r%�bX��z{Z��W)���%��Ѵ�Kı>�w�m9ı,N�}��r%�ؖ's�{6��bX�'���m9ı,K��L5����	sY�iȖ%��02'�����r%�bX���fӑ,K�����"X�� 6U�#�����iȖ%�bw�z^au5�Z�u��ˬ�m9ı,N���m9ı,S���6��bX�'���M�"X�%��w�ͧ"X�%�~��}�sZ�jkVfhĜ�(W]�T���� @�v7NOt��ЛK�%�ĩ�a��T�������{��7�����6��bX�'���M�"X�%��u�]�"X�%����ͧ"X�%��ww�%\���]j�Z6��bX�'���M�"X�%��u�]�"X�%����ͧ"X�%��}�ND,KĽﯵ5ekT����f���Kı>���Kı;�{ٴ�K�E�Dȝ����"X�%���o��ND��oq�߯����=��a����w��,K����ND�,K���6��bX�'���M�"X�%��u�]�"X�%�}�{WW-��a��\�m9ı,O��p�r%�bX����M�"X�%�����ӑ,K��}�fӑ,K��Є}�_3�a�hp����Q<c����&楡Sr�x��l)�vG:m��F�{)1�A����[�Qq�'D�8�Y_�u���ݝ�;���l�������ȕqB)�n�$4r9wa䞩�]d�v�]�gnwa�v�+�c [O<�ϛ�E�!�ۇ�W-����8ֱ��;D���T\�{m7G
��Fie�+O-��]z�,�Y���{�Ͻ�/��.��ˋ��`z^M��Z(ݎNN��u��!ˑ��#���&LjSW)���-�5���Kı?{��r%�bX���z�9ı,N���m9ı,O��p�r%�bX��=�5���.��5��6��bX�'��޻ND�,K����ND�,K���6��bX�'��ND�,K��~<,��p���w���oq��_��iȖ%�b}���ӑ,K�����iȖ%�b~���Kı=���p�4]Y�kY�5�fӑ,K�����"X�%����ӑ,K���{�iȖ%�bw>��iȖ%�b{����CW.h�Z��ND�,K�w��"X�%�����ӑ,K�����ӑ,K�����"X�%�����KËF梽���y0�q�o0M����ͮ�0�j�j�Vȷ���[�F֍ND�,K�u�]�"X�%�ߵ�]�"X�%��{�ND�,K�w��"X�%����֌�!�5�sV��]�"X�%�ߵ�]�!E6�\r&�X����iȖ%�bw���iȖ%�b~���Kı/{�k32[3F�jBk5v��bX�'��m9ı,O��6��bX�'��޻ND�,K�k޻ND�,K��OkZ�k2�Y���sZ6��bX�'��ND�,K�u�]�"X�%�ߵ�]�"X�%��{�ND�,K���1�.f��˅�kND�,K�u�]�"X�%�ߵ�]�"X�%��}�ND�,K�w��"X�%����GR+�/K���H;st�]��m��7W[Fsj؜��	䮖�s�ֳWiȖ%�bw�{�iȖ%�b}���ӑ,K�����iȖ%�b~���Kı=���p�4]Y�kY���]�"X�%��{�ND�,K�wܓiȖ%�b~���Kı;����Kı=���䡬��0�u��h�r%�bX�{ޜ6��bX�'�׽v��c��#�$q��4���:�9�����r%�bX����6��bX�'{��I�Pֲ�V\���6��bX�'�׽v��bX�'~׽v��bX�'���m9ı,O���6��b�ow��������#������7���u�]�"X�%��}�ND�,K�x��"X�%��u�]�"Y�7������w�جk7����B�";�u��q�A�$��Ga�vn�:�̘i:	�ôa���	���r%�bX�w���Kı>��p�r%�bX�w^��r%�bX����Kı/�������.���-�ZѴ�Kı>��p�r%�bX�w^��r%�bX����Kı>��iȖ%�b_t��7��Ve�橭ND�,K��޻ND�,K�׽v��bX�'���m9ı,O���6��bX�'�w���-��=ߛ�oq���}�~��=܉bX�'���m9ı,O���6��bX�"0�|�Z�H#����	"��B`D"@��V,"�U�"���X�E�@!ĒB(��R&��z�9ı,O����	t���f�3WZ�ND�,K���6��bX�'���ND�,K��޻ND�,K�׽v��bX�'�������?ݻ6��9���s�ω;N��1v��ـ/N뛓M6v��[����|u��v8�]kF��%�b{���ӑ,K�����ӑ,K��u�]�"X�%��}�ND�,K���$�+����˗0֍�"X�%��u�]�"X�%���޻ND�,K���6��bX�'���ND�,K����2kV5�u��.�WiȖ%�bw���ӑ,K�����"X�%���{�ӑ,K�����ӑ,KĽ�}����]�ZՄ�j�9ı,O��p�r%�bX�{Ǹm9ı,O��z�9ı,N�^��r%�bX��z{Z��5�R�f�mִm9ı,O��NND�,K��޻ND�,K����ND�,K���6��bX�%B�TQ�1A{��n[7�\�e֮jkZ�L�M-Q-��ճ�w,p;�ksq�M;��;���df'�Rn�t&-���d���nL���s��K�p&x;���v3kz��/"�z�� ����u�������\�e8��I��2o#�^6l��9�XS�7<�2��$v�����n�p�Y�n}Wa�:r��t��6��;�w����Go*�[���]\։,&h���5g�|����}�?/�Ѓ<�f煛Ovv��-Z[y2m����h�ۮ���/n[jy��U�f�5u4m;ı,O�k���9ı,N��siȖ%�b}�{�ӑ,K������Kı?}�Nf:�ՙ��h��k5v��bX�'~����Kı>��iȖ%�b}�zp�r%�bX�w^��r%�bX��}ɘ[�.��k35�kiȖ%�b}�{�ӑ,K������Kı>���Kı;��ͧ"X�%��ww��j33Y%.MkZ6��bY�
@ȝ������"X�%���]�"X�%�߽�m9İ?�FdO{����Kı;����h�ֲܺ�5s54m9ı,O��z�9ı,^��siȖ%�bw���"X�%�����iȖ%�bG����q����CΖ#����kb�ͤ��Ah�wF��]���h�s���ב�M4��^	 �'~����H'�w�6$�H?���&�z%�b}���iȖ%�b^�����s4L�WV涜�bX�'{�p�rA\T���D�K�{ӆӑ,K��}�fӑ,K��}�fӑı/������k5L�Z%�ZѴ�Kı>��8m9ı,O��z�9ı,N���m9ı,N����Kı=�=�&[��ՙp����iȖ%�b}�{�iȖ%�bw>��iȖ%�bw���"X�%�����iȖ%�b}��s3R�k&�5���f�ӑ,K��}�fӑ,K�{���ӑ,K������Kı?{^��r%�bX���{YL3SX7$�Uv�4�s����u�خ��ñ������c\C�/��X䬼NIj��?����ŉb{����Kı>��8m9ı,O�׽v��bX�'s�{6��bX�'���S5���0�5�Ѵ�Kı>��8m9ı,O�׽v��bX�'s�{6��bX�'{�p�rؖ%��}7�4K�k2�ԙ����iȖ%�b~����Kı;�{ٴ�K�O��X����P����<� 1�W�$���I�i�BXP��YV+Ρ��%"5p# Ԍ�T����1���	�h%�?}��֐���~��o��08�x/�$D>!w�`9Is|�$`���B��H�`� (�"H����	�@�I���Ьk�B�Ƥ�P#1�"����4�ǯ"�-!�G���i����RT�Jա�u%e��!�b ρ��U!��B$�`��@ `LO���B��JU-)~���p�@�� �@�����
$�I!
@�-*¤k�
�i(�c*D��@�
�CdX����p �� v�b�)�ܑj�gP��H�aSa�H�U����~E��~62R+D~D�6�iU? ��>����6��bX�'���iȖ%�bw�{�YMM75�u��.�WiȖ%��+"{]��ͧ"X�%��{��ӑ,K�����iȖ%�b~����Kı/{�]f[�4]M�Xj�iȖ%�bw���"X�%����ND�,K���]�"X�%����ͧ"X�%��{�l�;F�Eb[bzLvh=���sƱ��&�]a��zn�ɋg˪���0�|�~D�,K�w��"X�%�����ӑ,K��}�fӑ,K��{�ND�,K�Ӿ4f[3F�&\.kXh�r%�bX���z�9ı,N���m9ı,N����Kı?{�8m9�D�.DȖ'{��s0պ�MjkZ33Z�]�"X�%��￳iȖ%�bw���"X�%�����iȖ%�b~����Kı=���0��I��Z�eɭk6��bX�'{�p�r%�bX�{�8m9ı,O�׽v��bX���+� X��)RB0�D��Ng��fӑ,K���ۿ�&���ѣ
j捧"X�%�����iȖ%�`"�����Kı;�{ٴ�Kı;���ӑ,K�����O)�[���ugF+1f���Z��x�m�q6�B�J-Ƣ�smv#�q�ѣiȖ%�b~����Kı;�{ٴ�Kı;���ӑ,K�����iȖ%�b~��MMdɭj��u��ND�,K����NA@�,K��m9ı,O��6��bX�'�k޻ND���,K�����\��ѬՆ�k6��bX�'���ND�,K�w��"X�%�����ӑ,K��}�fӑ,Kľ���ֲٚ�2kZ-�5�iȖ%�b}����Kı?{^��r%�bX�Ͻ��r%�b�bw���"X�%����3.kYu�j�sZ�Fӑ,K���{�iȖ%�bw>��iȖ%�bw���"X�%����I��Kı?�?D W�:{?�5u�ne�fe��YsxL�O;���F|ciu�NXv�x�u+�-x㞤sq^�zvJ�v��c.��a�G\��;AV��Q�3�=�횡�k�On�7Z��ɦ�nnɤL��笔��K*Ek������ݱbT�� \�*�cgX[���1��Z�k�5ݣ�y�{j��b{r��IwN,��	U)	������ �ζ�������asdf�$Y�Y�q�GnX���O'"�g��j�4��uY&r�Ѓ��j�=ı,O����fӑ,K��{�ND�,K�wܓiȖ%�b~����Kı=����.�&�.��eɬ�m9ı,N����Q�,K���I��Kı?{^��r%�bX�ϻ��r%�bX��w}rk	3)�F�e�ND�,K���I��Kı?{^��r%�� �2&D�w�ٴ�Kı=�p�r%�bX���I�]R�2�IusZԛND�,K���]�"X�%����ͧ"X�%����6��bXb~�}�6��bX�'��޹���L�֮h̷Y���Kı;�wٴ�Kı;���ӑ,K���{�m9ı,O�׽v��bX�'���g�r�\Qb�G>�<��u��+�S��#�vHˇ��=z7Wf�N맢7E?�,K��{�ND�,K���I��Kı?{^��r%�bX�ϻ��r%�bX�����l�j9�h�]kFӑ,K�����m9�D� uP���?D�5�~�v��bX�'���m9ı,N������oq�߯�����R3�\4�|�Ȗ%�b~����Kı;�wٴ�Kı;���ӑ,K�����w���oq���߿��6�Z�V����bX�'s��6��bX�'{�p�r%�bX���6��bX�'�k޿=ߛ�oq���~�����䭥*��;ND�,K��m9ı,O��ND�,K���]�"X�%����ͧ"X�%��=�m��5��0֮k2���f�7WF�z��L�s���;�6��d�\�t)5���ѣE2捧"X�%����Y��Kı?{^��r%�bX�Ͻ��r%�bX��}�iȖ%�b}�M�MS	���˫��Y��Kı?{^��r%�bX�ϻ��r%�bX�����Kı?{��ND�,K�����\�Cr���w���oq��_���r%�bX�����KAX���MD���Y��Kı>�]��r%�bX�����d�4h�5ua��ͧ"X�%�߻�ND�,K�{ܳiȖ%�b~����Kı;�{ٿw���oq�����iA���pi��r%�bX�{��ND�,K���]�"X�%����ͧ"X�%�߻�ND�,K��a�����5�K�[�:��uJ&{fH�-�ݎ������";���	H��p���{��7�������Kı;�{ٴ�Kı;�}�iȖ%�b}�{�m9ı,N�����cS1S�X�����{��7��}�fӑ,K��{�ND�,K�{ܳiȖ%�b~����Kı?~����jj��?=ߛ�oq���w���"X�%����Y��Kı>����Kı;�{ٴ�Kı;���\��fa�F���6��bX�'���fӑ,K�����ӑ,K��}�fӑ,K(D��ESV'��|m9ı,N��~�E�����˫��Y��Kı>����Kİ�������~�bX�'����iȖ%�b}�{�m9ı,O����Þ�\t�@D�64sl�^\)[.#=�v� ��e�]ڶ��\�Cr��ӑ,K��}�fӑ,K��}�ND�,K�{ܳiȖ%�b}�{�iȖ%�bw;�\ɒ\֤�5ua��ͧ"X�%����6��bX�'���fӑ,K�����ӑ,K��}�fӑ,Kľ�����sNj�kE��m9ı,O��rͧ"X�%����]�"X� C"dOg��iȖ%�b{���6��bX�'��|j���fk$�ՙ�֬�r%�bX�{^��r%�bX�Ͻ��r%�bX���iȖ%���ȝ����fӑ,K�������֦֭�������r%�bX�Ͻ��r%�bX�����Kı>���6��bX�'�k��ND�,K�D�=�߮[y��ٚW`Kv6^ړi��u�<�U����/[�Ӯ�k�J՟�B>�ݳ��84��q�ֱĸ�Qvqn8÷�n'�n��<4om��ke�{;�6�J����'n%
iP6t�ζ�r��W[Z���ru�/�|�'�s�),<s��Y�!W1�m�ݳ��``:6ӹ���S�a��8ns�K�S6��4z�e��A��ݭԲYsWR]]dЯ�!�Dw������Z�,lu��.�]���>�>;E�f.�M�'tԝ7l1�¬ᜓ��j4��kY�v%�bX�w��6��bX�'���fӑ,K���w�a���L�bX���fӑ,K�������u��4h�3Fӑ,K����,�r%�bX�����9ı,N���m9ı,N��p�r%�bX�ﯸMY�2]Ku���kVm9ı,O��}v��bX�'s��6��c� ���=�p�r%�bX�rͧ"X�%���{[,��q1�������ow���ٴ�Kı;�}�iȖ%�b~���6��bX�'�k��ND�,K��z�C�j��WV���r%�bX�����Kı>���6��bX�'�k��ND�,K����ND�,K��po�Ϝ�\^�ֺ0=O��F�޲q;9'v���!˒麉������pi�iȖ%�b}�{�m9ı,O��}v��bX�'s�{6���2%�b{����Kı/��fMk.k$�ՙ�֬�r%�bX�����9�' �? ��QA(�+T*;���'s^�m9ı,O���m9ı,O��rͧ"X�%��1i�k4�>{�7���{�����fӑ,K�����"X�%����Y��Kı?{]��r%�bX������٨4�9�?=ߛ�oq���}����Kı>���6��bX�'�k��ND�,K����ND�,K����a]I34h��捧"X�%����Y��Kı?{^��r%�bX�Ͻ��r%�bX��}�iȖ%�b~��������AnxeQ�\��-�ݫ�H&/k9!$=J�.�MW:G7�MZ]\�MND�,K���]�"X�%����ͧ"X�%����6��bX�'����"X�%�����e5��5m�j̗Y���Kı;�wٴ�Kı;���ӑ,K���zp�r%�bX���z�9ı,N�}�.��3]Xj�Y��Kı;���ӑ,K���zp�r%��Ƞ� �]�Ț޽��Kı?g{��r%��{��?�����[�����{��%������Kı?{^��r%�bX�ϻ��r%�bX��}�iȆ��oq��￼�Ԭ�	���=ߙ,K���{�iȖ%�bw>�iȖ%�bw���"X�%��������oq��Ϸ���V,�W�:\7js�Rs\��;;[e���6���NP���6-UꜲ��w���oq��_�����%�bX��}�iȖ%�b~��8m9ı,O�׽v��bX�'���Lֵl�kZ�L��fӑ,K��{�NC� �L�b}���8m9ı,O����v��bX�'s��6��bX�'};���!�&f�]\Ѵ�Kı?{ޜ6��bX�'�k޻ND��@dL��￳iȖ%�b{����Kı;���I�X��ˬ�W3SFӑ,K?���>�����r%�bX����6��bX�'{�p�r%�`TV�~2%�|p�r%�bX���z�SZ˙�n��0��]�"X�%����ͧ"X�%�����r%�bX���6��bX�'�k޻ND�,K��Z֮֬��tg�]�m<q����ܵm�/[]r�Kt�L4�H��yka��O�w��bX�'{�siȖ%�b~�|p�r%�bX���z�?���dK��w�ٴ�Kı/����Z̶i�nj�.���"X�%�����iȖ%�b~����Kı;�wٴ�Kı;���O��7���{���}����Rh���|ND�,K���]�"X�%����ͧ"X�%�����r%�bX���7����{��7������z�T\����Kı;�wٴ�Kı;���ND�,K���ӑ,K���{�~���7���{�~���ئ4�9�?�,K��{�m9ı, ȑ1�w�� P����-�k�P�D�TE_������TE_�"���DU��UW��TE_�"�������""�AX�0",�� �@�H��H� B �@ 
�X�� 
�@"
�`
�U�,@�H�� 
�R" ��DU�������"��TEZ��*�EQ�UDU��DT,�DU�qUW�TE_�EQ"��������)��a��&��8( ���0���      4@M � �  h       ���

  P   )@P
�A�

*T%J@(HR�@� �
P�))!E �R� <   �� (   
1 
��19:r�.��� @fi��w��=o3B���5� �h�������     �  d   P z   0  ( C��^���SӐ^��� `1��j{=Jx�4  �� � H  � �Jfޚ��[� ��z
��nZ�%=����΃ 4,΁�� �:2��w�b �z�y�`z��ݪ���WU�wy5��)B�   ��4ުL��\F�ru;n�:�� z�6$�ԣ�[�Ҏ� n��=�f���Uv��C 4�����U,MNۛTXJ94��W�\�.�6�p<�    E�ޥL�Jf��^&T�	{� �A�A��bq�n`k iK���8  ��1V3I� ���a��Y9�^g#�� �e;���<l�i�`���< �JP     ����ɥ1�֮`t��,  6,�q]�`=<�t�  9�mNN@l= W����K�9��� �c}���7�})�����S2R���Ojh�T�M h2 D��R�h  !تT�)%  !��BT��)*Pa2 �5%"D 4f�������t������{�C!)�Og�=���cw�EEz�r��U؊

��*����U���*+(�����;g���?���~���1Df�k���Yh�����I�W�h�DŚ0��ؘ9�b��C��8���$�	0 ����0#��[x�l����0%��Q�	y�灪�Z5���1E�k|��p,�f�m�#�f�1�a���n�^[�M�1���-���ZH������<�<�K[$�Y�I�O1ӻzc3���g7�8���s9�Ƃ �O|0&�F8{����y�U�|2s�6x����F1�č��S����{�\V�LtlE����J9��ci$�Ѩ��+4|E,��2��ID�HBI���;�M&є� 1C�KR��}�E�	�S���* �t`�I8k���ֶ|q�1`�?yk�3{�|`�\ַ�}o��цϷ}�<>���'��!��c DA!���T�K8�I�N͏(�ı#Ѿ0AѦ�4�j4l�s#	p����i;�����Ʋͦ�`�aa��٭�F:6q��[�$a����ѳ�e}j�o�6�'<4���5���$�x1��kLkF��ݬL�61����������p48���a��mx��	/ ��'#A��Z�90@��>�8��6�h6�4n1��p�3_y���0PRQ�����٭�N�1L^�ky��qtmq1$�D2SD%��F��0��F	�V��# �Ha�����K0�2�I��BP���P&�������u��<��b� J�,��b�:'`�Q�l>OG������_�W|�����	�p�#���8�
(YX�f�f���K9ϯ��\����F�3M��������,�;�d�%#E��xC`@��y&&�`�IK�k�K��������R�&!�kbG���p�Ѵ8��8x���d!���iޟ1��!֍orG�8`��oX�����0��#���I����6�;�0ѽ�h14f�}C$G~��WyO1�s{T�.�U��|-�ƹ���s���:f�4sg�̳9h0Na����Q����#0��r*�-��捄��>'>,�f����<Gӛ>l�<7�{�|�p� � ���$�lhQ��'�&k ��u��,��O�xt��-�m��c`:%�����'�j��A�Df�ݞ��gɠ�,H�>��6b�	����&:6<0��1ta���!�H$�~4o��	1�獆���|w�k�f�LM����5��4�만xkZ��s5�~6���a�8�Y�ӷ���==5��& 9�ag�K��5�`��Fl���)S��o5�7u��{K8��^�o�1��R4�Df�Č����ؑ���M3g��LXZ]� K�a���i���m:�o�Q����f�!ÆE����w��.�}�]��|�������.fk|�%CЅdf~<,�f�k1����a��cX{��.�*)QT��V۬����k8�n�T��c��h���X�p����k|l4�1�gi	����N�ӿ �[���zz,SC�]��q�7����ٳc�û�����*I�!�#g�>6Xhv���U���M�zÓ����sq�\����2^o��[mo��5�xl|xk��r�е᏾y�����[�Vo_i�{O���H�������cG����ag�Xkd�h6�s��s�n5�6�6h�Y�l,y�F��ap�N�3[+�#�3�h#2�1��k,�o|x����������i	,�A�E�24@Adi������ݮ6�$1�ֲ���sF�����a�f��Y��F�7���s��opV%�f�m3�)瞗����8j6�Ʒ����f���B�0�$�xn0�� �F���08�8�/=><_LZm�Y��s5�p�F1���Af�1t�țC��PD�A�	�$�έ&t%�jA�C8i�`FKFќg��Xo|֭sg0	���9��(���Q���a��'�a��������m�]���{}�����W���}�n=�n��N1�a��h#caF���4��5��H#6��[ܚ��Ѡ�H"$�$��1� �4:#D�,�&f��1��
LX�̴n8�АiX޲��4�I�'(!�t�:��^�����aĜB\1�@@�9���b�DsX!z�Zހ°��7�[9�'=0}8�3K�30$�m&���٢0�p�20Ѿ$%%b:�=,�!��p�|���14��Y���I����6m#�L�'o�Y�[����`hjI�c�´�[����(�#2,3L��I�u#����i�`��$!&�ѳg�$��e�o �����F8d�:��6�E���h7�HIR�8A��J&+#!3�y,O�Α�b�[�0�#$�j"�If��fm7��;�4y�h>�C�Lc�Fs\(��-��� �0ٰ��J`r�mYx�g)
�73�C�m%�Z�̵5�2�������ma�[6�&!�pta�c[6�'�'f#�e�x�.eG4X�X$��0&$�	m�Y�y�3q4�42�L0Lxm$�!#8|����2�8N��R�A��PY���q� � �E�>6�X�0��F�
�I1�,,"���/R0���$%�Z�<8��{kD�p�Á#�2��� ٣Lf�A@��DD��N�n�-d�G��M�8ƚ�,,�XZم80,+��Jb��!��>2�:l׆����Ö��|q8oݶkf�3��aae�0a�[5�x6kia���q�'N��PC&��<��c1Ѿ6�~�I������#a���<�x�{=9��鞖S@CbNg0$���8h#kz��y�f�db�#3Lb�I���<�{��1g7�E,��ӛ8;sIaf�� �N9��M�3^��6Y��Df���s~��}���1���d�����$8VM#�� �A���i��<����3.����f��k�y�oF��k�c#
��_a�<�Z=$��B=�6�	��8���O���{34�o�9�6����4H`Y�I�a�Fm���i��-���`��	 ��n�scD�}�|�c5�f�g7�h,С��=��s5f�moi�g<9�}�����ǀ���H1�o���Ho7�[<7k_h'Ϸ�X���f��E�����7�&uXm���y���9���q��4��1d����'l�fkg����Ϗ�4�x�ϩ����ad`A�f�� ��jL��m�Da�>u��������Fh�FIœ1�᭖h���G�#Zb���Ͻ����>�!�#5������ ��t����ց���Ζi��4Y��<�[�df�\��s�;�w�;�q � 0�����r 2(0�9	�3�2�)"�H�qpLL	�t��|t<`��l!`���b���3��n*q�������8�(�	))�	1�b�z����bqp<_|-�����x��.	�� 1Ӊ����c�o�ăt��$�҉8��I!���x��<=�5A�pL14��������'F;������� �$I��B1Yp4`i�ЌSF;�4I$`i ��Ӆh ������ߞ����	���ݭs�H�Z�X�*�ψ��q�������1G�x'��Ǣ~,y�������X�qR������^Wz�ھ�<�\���>�5{^���w���j[�՞�m��m�� ���@ �c�  h   ]"�{m�8[m�ul�v��m �����[@�d:l�w 8��m�m�'7���OB+ϯ(�įZvԼ<��Fj����v �힔���| ��oe6��<,X��*�;m����[ٖV�]k��^�;F� ��1�c��T�
���z)m��n�����l�8��F�!o\�4���?h��I��Z�k��%�K�h���P�`�M�6ZC���� ��u�� ��m��1m9UU��uUI�@T��` X`��[m��E �l��-�kf\   �  j�   l���    j�SUUJ����UYE�������i��  �| �� 5��v�hlh9m-6  �%�� h�ؗ� 	e-�o��l �$ �  mH   -�  ��m�[M� H   �[v؃ �#��� m�  #��    	  8I#j�-�n��˪�-� 6�� [@ $�l   �Y0v��i,�����m�� +}��� �Q���[VʴX�����8�-���H�`�`         H�� $m��` 6�b@ ������� m�-4��� m�pE�m6�$p  $p ���m�l ��_�� �   �,�l�m-� H ��m&Y�� -6��H����L�p����p��   �cm�l� m��h �   d  ��m�   $  t�     �p6�e�m9m�`��`�Mm�	6Ͱ n��	;e�vti��  8� @�� ��nͱm^�m����l�t�I��@մ5�M�� 	�l�� �lҴ��m�R%����C�sid��(� I�m�[�V-�p@U�� {8�-�� 9y�ڕ皜�(P�U�N;i	 �[�kn�@-��. H �m�Koړ��e�m�V�R�r��/����۳��O��m�-��	8pH����-�ۛ.�J�UuTR�q�.�a,saɺUݣ.�  ���6���E�D�� ԍ���m����^�6 ����{ �$h	K����[ �$�"ڶ��)m6��������m�P �3��
8⪪�� [@/Y(6ݹ��2'���m�� �}vu��s���l��J��  k��^sr�� 	�Hp� ��b�88m����tҰ	�f�[P��-�O-�*�pX�UJ��b��j����omtb]Ƚ��}�۴ﻷ��[����{;;sbȝ�3��c$�Zcx�d��(S��B��k2��bk�TWd+�۟0V�Ҳ�H�$���si���<[�;V� mMyp �����Ͷ�m�ml6x�g�l�Bu�@[VPb�%�n�b�vQ�c�0Ոe��ț4���KUUF��)j�r�v�v��*�m��!-��u\uml�v�KU/Tt�Yx]  �t�I���I�n:��V�$�M*�n႘�UJu�5W5@d��mURƮ6�ep��e�� 
�N1ċ�pSn�˒-�d]��EQA��@qen�q-Usj�:��2���n�j۪u�48u ]����*�][L�Zګm�6�Z�%���l���9�f�u۷1��q� ��i%o`Ή��%��[��M� 6��J�g[U�S���p[T�p[�.K:l�5�&F�p �GQ���f$-�+j��e
Z
Pp  H h�ݦ�������{l�F�[�ٸ�j�!�Z�+1���r��rz�H�Ӯ7�m �m �a�M�j�lm�`rn�l��Lm[  ��\�Jq�+%�q��R@ $jV��8��A�m�: �`8( �2h�M��'$�J�N�� �6��pm����M���`�́UY�c�V]�HjC��m��f�D��m�ȑ����@�i������Y$�m@�3UTb�k�[�m���H.���-��[�r�Y*6��%�$�W�}���۟���]��am[ղwrFݮQ��P9�;k�˻De�Ft-ֹ�^I��m� ��2/Y��l $	2'A�bu�9����������\��T�0���UWY؟p�n�-��*�*͞	������:�G5��t�� m������_/�1uA�5�$ �[An�&� �h�t$��A����]�v[i3���l�M�� ��m���/��m�&� t�6�.�m�[$��  ���"I��zM��ޠ� d�� 8m�KCe�v�� ��N���I���0$&�rtѿ���t�&�$P
�uS�
�8*��������� Ժ� r���l ��&�mmͧ%�8  6�m� m&    6�t�� m�)p  d	�g@  ��m�  Nm�h׮�� m��c�W-	j+��m��cm��	�b@	��n�h� �8�ԒG:�m-�� 6j�M&�l�%�z�k�kk��������c��U7`@��ԅ�}��#I������E6�:�� ��km�.�$ޒc��I�����3���Kyc$!�$�H�|�ʿX�����m�������9�[&�"Z�	)ֹګ {m�tUG[�k�C�m�F)Wm������۔�7Sct�n�N�VT��lq�̻-[J�;��c�i�i	M���m��5l m��m��Y��&��[��^0�S�*����zM�iZ�R�'�� N�N۶�{v���  #C�N�E��v�z�m� 4�n�h�)M��m �e��ZI��`&Q�]F�O*�UUt�9vZU�H9�[m��Ŵ  6�H9bD�֤� �� �m6��W�%��%�m�886�p���3gMm���y��`�`6���m��U�*-�n��)�uUTU.�;6Qt�f*����N	%�6 ���U���[eg�ԁ  Am$�6�   mm-��o#�_����[z��� h  x$�ntZ�h�5$  .���ɉ�- il��  'F�\��HI�   [d.��isZz�V���]K��Q�, z� �( e6 -y��B@  �[���mC&����km��-��SB�@m� -6��ӯ�m�lۮ�\���p �ͰM��� �.�A���]�۰$��%��۰p�eU+sR���G!Nʵ���5� �v�.�� �[C��$�T��*�VҭWO$� � � -�� k3ݱ�нrI���ci$�&� ���m� 8m��`8U��k������)d64��lm� ��   �        [���$d���K(��Cm�Ś��!�6��!,�*[3�Kz�-��  $K��ҭu*�R�P��\��� $�v�   � 	21���Є�=UP �T�m�eY[˚i	��  ��m-�ŵR�K��xPj�Cq��2 sUW]V�M� �4l6�[N8H6�[q�m���   'F�9,�m�n]�k��nջ[{f��v� �sm�Y�&�9Cu����۵�H6� �	e ��M�H���j���m�WjE�F1��\��u�~���*��u��3M�-�m hֳl��$�v�Kۋu�6R�	2�%I˵�9ۢZ�p��L�Y)�k,d�V��C��-@K[( m[ �m�$�`u�		  m�m �jݪ���vXYV�)V��y���  $�Md��:� !�-�p �|�GX�ml�r�k�-�-h 	
P5��n� N��m'l 	6��K)m�[%�ܛ  m�bK�I�����u��\�l5:w"��UNج�+��-��,�iz,m����kx�T�۴�^Ė�e5[��L	  6ܶ��hn�Z�vR}�&�3����n-Vl$��5q� T�n�p�cl�*�Jv̆��*=t�QĦp�+kJ -� ���KteM#�Ť���[GRڝ8p�]n�[�6 ���U*�

���]�e�[@ H Ŷ�m�d�@m�      8 @$2	 $���m��nƵ�m�mf`$ 	  -�o       ᵶ� mm���'@�cm��ݳ�v��H"�������{�������(	�Qd?�_�OQӴ� ��O�����h�T�	���*���ǉ�
��sB�f�A���Ң��@v�8� ��ب!�����1: ����x��h�E||A�^�+�=�P�_A�$�>D~�eXBP�F@HH�8�����D �b&*uUҮ ����N��ꉥ> 4)� U�Q��:P�U�Th:^0�-0�C%*�3)K2(�HLA�)J�ڝx�[G�S� ǂ��z*�_��|(��hQ@�& �:Qq >E��S�Q~��/��{ �!"B�)0H=D����>�#$@��W�'��s��G�yU���D|OAW߀���$���i@�>*��tT>�$�!D&�\���U؏���(␁=/��BJ[ v��vԮ6��F�,Y�]G+uv�]	������x��(�����Q�wn�	+g�,�s����Pw6�'e�������r�z�D�ڦ����)-v�UX�k�n]�ӱ���N�A�m\��7*�JP�;a�#�8��8*�^Z֡�Ӹ��ul;���\�JqE�x�M6N��`7i_J�!�Zڷ&�$�[(��8J������NR�q{��t�簵Hyݸ:6��蛞�-.x8�N7m!���������t]�qݽ+[&�y��&���Y^{��v�N��-�:�7E@Iiv;6q[O,lT��k�x�)�Be�\�[h����|DƮ�qn^lWn�^-�
-9��*s�uq��'gO�R@��Z�+���n�]��a��-����kѦ���ɚ3�{8����q���F����h�1�1����zR�=�Ο*#rmv�v�O<Y�bѩ�I�x��cI�d6�70j�������̠̆U�%�C:,Gmv�kaX4���ˈ8��{k��Ë�CE`����ڞimp1N�kr%tc��[��ڳJ��Uc cK��[t �@�Y�^ֵ���sv�<t�j���v[��{c���#�pA���	����3n�Ao`jNS"
&i��V[N��eT��va�u^���v4���.�q�<�����^�l�EpD�� 6��]�WU����&L� ���e��v��ۃ]�`��8ާh�K/`�_�'��^��U��5!�zu*�9�QP�ڪ��	�f]��]�!S&�tѤ�TV�.�;]��{8�A#ƞ���'�����i��na:ݽ6����W[���9��N�\�k���Dj{.�ӗk�j2e!^3�3I�m����	��{S	%�+�,EK�����-ӣ���|b��L��v��g��,[3-���x.����؉�����놭��mP����j�Z�ٓ�e�=U !�W@8#!*�� �C�`�A~�~EHFS�־=�]���Ń0)��vyUn�b9�Sd0jg�L�O^̷��Ssс���[�Q���'	�˥�+�]v�Ű��j�F͆�9nS�=���
�Y@7d����=y�C{9ţ5
l�����vgu.[ �ga=����3Lr��]&Ы�	I]�gc�f|����r��O;��iyɔ���b䎪��F�H��'Eļ����J.�؎�[z+2�Zc,�Fg��Gý���ʣ�sț��ē I<hbO�,�z��hy�`����D�DL|�v�U���Q���T�����7s]�&b#*�����w�{Ϫ��:�
a�x��h�h��@��S@-�4��Tcnc�	rM��h�)�����4}��<$m�9"�;�U�����4]�@��9L�?:)�s�i�,�������$��Sg����z�-�ْ���l9�ؚe��4��h��@�}V�{��0�F�X)rh�lٞ_<�3�1BeE�`�F@� ���\��r�{��9U������LB�2B94_U�w>�@-�4��h��H�M�&������� ��v��vW�hޘ�\��9�y��N/�}~���4_U�w>�@3�w�+Q�D5��.�+����N�<7̥��OXɛn8���nX�"�d���LXǋ )&�~����hϪ�z� �ԋ�Nc�7RM��hϪ�z� �m���D��NF��9��>�J�߻�\%eX	FJ� �t�٠~���?/N�b1��b�G�[�h�h��@�}V��:�C$Q<X)rh�h��@��U�Uz� �s��"F��tF�F\r/l�t�:���Q�T�[;W	O3vp��&!Iᄂ�h��@��U�Uz� ����]cR1DԂJ))�������sj�9���̮�-|5B	�c̈́bq~�����h��@��U��uo��Lǋ$	�������+����D�D�"$�#)*����ꊃ����������X�Plҧ$ҦԒM��h��
�W�~]k�=;���ɟ�ۋ��<7']=�yv�M���H�
Y��u�b�gs�芇5��b�r6�oy�
O~ϻ��JS�߻�)JRy}��y)Jw����)J>ό��,խ�3z���JR����qJR�ϻݏ%)O����R������<��=����Z�{Ѽх���o\R�����c�JS�����)=�>�%*f�q����b�0�b��ӕb��<��;��qJR�߳���R������(|����R��{��t����Y�ٙ��z�qJR�߳���R���N~���┥���c�JS�k��)JP	+�T0�A		3fb�)3P� ̡�Jb������,5o#6e�V`�ob��'c�ٓ���ja��Ko����M�k�c���2�7�cl�퍮�œ�I��\\��m����1�iz�9���j�[q�^
��c<<d���i�g�6m7Q�q�[8Y�V�#���4s����V��rշdǩ�q��j���v,u����L�;p��pg������H�����lMܛ\��i�����w|�����r�]M�=��cv��:8�ʃ�l�c���^�K�ض��\pƺl�����=�Y���)J_o�R�>w���R��u���)=�>�%)O3���ћ��f�F�5��JR�ϻݏ#�T��Oߵ��qJR���`�R���{�)JP��eu�kf�3v������%)N����R������<��.���R�>}��y)J}�������7���ٽoy�)JO~ϻ��JR�~���)C���ǒ��{���R�������3V��0��{��y)J]����(|����R������)JO~ϻ���`y�=G�4V$��f	4<]n�'E�}�k�]��5�$��j�E��C���Ԗ�E���[��(|����R������)JO~ϻ��JR����)^e���j)��AI3�<��2��<��qz���|u)I�����JR�{��JR�ϻݏ%�*�jSvX��v��).r��w���<��.���R�>}��y)S1��⹘	�	��Ь��U8���T���� Bg�����JR������)�����)=�>�%)KϏ��Fo{ц�n����)J>�v<��? �����8�)I�s��y)J���y��{�Jd�LY��񨮹�M���:��A�nF��,܋ĈtE�734���5f�n��kz��{��R��u�s�R����w�������JR�ϻݏ	�	��:�ULm�BT��j�`&`�߳���? �d���o�R�>���%)N�_w8�)C��j֎ᙨ��V���[��)w�w|R�����c�}:������k��3�R����w����_w���ދz"��z���)J>�v<��;�}�┥'�g���)w�w|R���]`7����RL�O<��̵�Z�)I���py)J]����(|�c��ff;̄XBjҥE4P�/Y��M;&�m� �Z�Ks©��F�]r뷽[�k[�e��z�qJR�߳���R��߻�)JP��{��)�u�s�D��b�c�*r�-Ҥ�����	������JR�ϻݏ%)O���8�)I���py'� 9)�~;�v�޷��h�vf��)JP��߶<��>��┥'�g���)}��|R��{�HȡS�
��t�M�0Lf￳�R���w�%)K����J�!J@���E4�*��s��ɲff9�x*�m5E*l�j�`&JO�ϻ��JR��w|R����ǒ������)JR|||�3���oy��m���wn.a��#�.r^,b��8霘�Ȑ���IY�y��u�8�)C�{ݏ%)O���8�)I�.�<��0<�=�]�0��)#�j����v<��$�Jw��~�)JRw���<��/���R��w>��Z݅���[ݛ�ǒ����{�R������<��/���R�>w�����������N�k�����������<��/���R�>w��򙀙��f+������]b~*��E��Y���)J_�~��)JP���c�JS��{�R������<��>��w5���"`�q�x�u��;qpb;�?\G���H3�d�0�pN-��f8�\�=�^�b۪Z�7e����nq۰���,v:(zV�q������¼�붶ԛc��@�8�B)�v���!���[\��͝�Ml�`��-MQ1�u����I/Lћs�����A����.j�H'v�H�w����ݧhۇ\�
���M���roF�޵k{����PA9�'9[�o���ݶG���1m�찎�؎{*NFV�-��ǫ��jܥm��i�'N玶��ݷ���~��R��u���)>�>�%)K��w�)J��e�Y�۳Z��޷��)���)JR}�}�JR�{��R�>w���R�����Ӽ��Y�Y�����R������<��.�����X��߿ly)J~��߳�R��^����+5�fZ���o������┥�w�JR���┥'�g���)�o���j���z���7��R�>}��y)@~D'�����R������<��.����-�~~v�����*ֶ��#s[��=���1�����v�[fv����d�p[7�oC�JS��{�R������<��.����)<��t<��>��]d��7&%����<���3�]Vy�y��P�dj�7)w��|R�������R��u���);��I7^N��E�E*j'�ff��s%)I��{��)���)JR{�}�JR�g~���[��h�u����)I���C�JS��{�R������<��.����(~���Mfkf�Z��o[��R��u���)>�>�%)K��w�)JO.��JR������;X�������m���-4sؙ�X�9�\W��X�ѣj�a�Ѷ�/��mf�����)JRw���<��.����)<���y)Jw��s�R�>z�eH21��Şi�y�����Ӓ�����C�JS��~��R����U�i�y�ӫ�0���I5JR����C�JS��{�R���?,.���{���@X���!1�� �X���2���h�[]�ث��c�q$D�cI%�Kb��XoX�����a�da��Sb��3,r�h�1	���i�چ�М� 0�,C�,rt�Dl]�1��2� I���6.�րФ���|�ئ�HOD6��<?(*8Q�<S$_�S�C^
���T��p���{��)w���)K��u]`'��1�	�H��<��2�]�qJR���ǒ�����┠y��k�4��<�E��FF������R��}�v<��.�����BP�%	Bf`�%	BP���ߴpJ��(O3�(J��J��(L���(J!(J��?~����P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'�)����4yf��y��f�\���7h�p�Xq�6��f�H1;��#�Bj�g�z�-w��w�n�m�B{�%	BP�$BP�%	Bf`�%	BP�	BP�%	�������(J��"��(J3�(J��J��(L���(J�����	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'����<�J��(H��(J���(J��"��(J3�(J��{���(J��0J��(H��(J���(J��"��(J�~��-跬޳7Y����(J��J��(L���(J!(J��30J��(Os���8%	BP�'��S���%	BD%	BP�&��(J��J��(O���g�	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP��~���(J��<���(J!(J��30J��(H��(J��߿~ߞ	BP�%	�%	BP0�X%	BP�$BP�%	Bf`�%	BP�g��W��l�akV���z8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP������<��(J!(J��30J��(H��(J���(J��;����(J��<���(J!(J��30J��(H��(J��߿~ߞ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP���ߴpJ��(O3�(J��J��(L���(J!(J���Wk�gȻ�,�����%\���	BD%	BP�&f	BP�%	�%	BP��%	BP�'{��8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP�������(J��"��(J3�(J��J��(L���(J�����	BP�%	�`�%	BP�	BP�%	��P�%*� �^��
�ꈤb/���%	BP�'�9��P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B^�w/ٕ����k{�k|��(J��(J��(J��(L���(J��(J��߿~ߞ	BP�%	BP�%	Bf`�%	BP�%	BP�&f	HJ�*����>@�@����~�?}�v �ӦY}�j�{�a�5��U�J�n5�d��ڍ����۳3�%�.�N[�l޷���l͕f������(J��(J��(L���(J��(J���(J��=�߿k�P�%	By�%	BP�%	BP�%	��P�%	BP�%	BP��o����(J��(J��(L���(J��(J���(J��;����(J��0J��(J��(J3�(J��(J��3��߷�P�%	BP�%	BP��%	BP�%	BP�%	��P�%	Bw��~�Y����ضo7�pJ��(O3�(J��(J��30J��(J��(J�����x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'{����%	BP�f	BP�%	BP�%	Bf`�%	BP�%	BP�&~�����J��(J��(J3�(J��(J��30J��(Os�����%	BP�f	BP�%	BP�%	Bf`�%	BP�=�{��v��۽ߎ�����"��w�x%	BP�%	BP�%	��P�%	BP�%	BP��%	BRI���~���(J��0J��(J��(J3�(J��(J��3����~x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'����pJ��(O3�(J��(J��30J��(J��(J�����x%	BP�%	BP�%	��P�%	BP�%	BP��%	C��:�������&&J��0J��(J��(J3�(J��(J��3��߷�P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B{��~��(J��0J��(J��(J3�(J��(J��?~����P�%	BP�%	BP��%	BP�%	BP�%	��P�%	Bw���	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	B{�ݿe����a�F�5����%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP���~��(J��0J��(J��(J3�(J��)�!(J������P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B~������(J��(J��(J��(L���(J��(J��߿~ߞ	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	�tgt��������J^�g��)����srmiô��vk���N��+�	�X��<����2�]m�dq�WY-,��w2V�ue����:s��Mq�#p�m�N�p<�nv��ò����7*�[�l���꽜ۮKw�m���Nn���5NN�հdmnq���qn�\s趉����y���ԍu�����[�mB���w~{��]����4w-�ݎզ���+��$�5o���p�}I]p6�͛f�����o7�og�P�%	B}�%	BP�$BP�%	Bf`�%	BP�	BP�%	����g�	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP��p��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bg�߿o��(J��J��(L���(J!(J��30J��(K�߿l��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bz}���}�QB�����v��۽�w�n�n��(J���(J��"��(J3�(J�������(J��(J��"��(J3�(J��J��)L�������%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	~����	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'����<�J��(H��(J���(J��"��(J3�(J���.���Y�ޭ�kz��(J��<���(J!(J��30J��(H��(J���߷�)J߿~��R��u���);��d��s�Z( cC�	��w2R�=�{��)���)JRw��ǒ�����┥'�g{��o0���l���%)N�]�qJR���v<��.����);w���R��ui��c�	�F(��@��q��gz8B��5,�EEÛ�	�����tַ�R���{ݏ%)K��w�)JN��t��y)J~��߳�R������@_.�cv�s9Is����U'\P�%);w���R���s�R�1���l�ْ%1Ÿl'P6�DTT2�o|R���w��%)N�]�qJ��?w��%)K�߿o�R���
2(Tႁ�6�:��ff3+1\�JRw��ǒ�����┥'n���O<������F�F�dM�4�[�JRw��ǒ�����┥'n��JR��wۊR���{�]�hլ��V�.�vf:�7���6K2��\L���6d�)�A��3jn��{ݥ/߿~��);w���R��{��R���{ݏ%)O�߮��+T[���3{��{�JR�����%)N����)JN����R����|R�����4��T0��M�M�01�Y��b���{ݏ$/_UA�@�'J�㹘	�	��Q6L�L�Q���moF���a�oz�qJR���v<��.����);w���R��u����Hz�h��lcn������RH��)G�R_�~��)J~��߳�R��}��y)JG��k��z�ٺ�v؞����}��l�^��vym�v;U��7��Ul�h��͙hѺ�o|R����{��)�����)>����R��߻�)JR{}��MZ���V�oY�oC�JS����)JR}�{��)w�w|R�������R�����h޳{��Z������R�����y)J]����)=��t<��;�}�┥��v1�� ��S��ff�㹘	JOo��%)N�_w8�	��I���c�JS����j�elۆoy��|R�������R��u���)=����R����|R����;��,��۷7�`��lֺ9W�[�v/^�ݖ^����=rFk�z۵��{��v��~~~]��)I���ǒ�����┥9�ּ�O<����[X䍼mĖG#��R�����y)J]�{�)JP���d��fVb��	���c:T�������%)K��w�)J~�v<��;�w��)JO~�v<��/;��5���7��F�5��JR�߻ݏ%)N�]�qJR�߻ݏ%(?2��ۮ�`&`&:f�����)��q7)Jw��s�R�����y)J]�{�)JP��{��)���3��5�X��0�1!����FrOH�n�D�d�;[T:M�mνv�쵝�A���c��t���Q��]'[��p�b�ґ������F�A���a�&Z�x��n4����g�'��mv�Xݚ�F�X�u=Re�ɓU�y�;����ڹ{c.	�]n�t#rm�e���n�lM��g�մ�]Z�eZõ�f�l�U�I�z8��;T=�����{�68w�c�g#�Ӻ��1���s0+�2���u�n.���Z��f��������v��m������﷒��߻�)JP��{��)���)JR}����Y���a��z�ǒ��߻��JR�߻ݏ%)N���8�)I���ǒ��~�����ٖ��f�����)J~�v<��;���┥'�w�JR�~�w�)JO��wyk[�VY�t[7�oC�J�'~�;qJR���ݏ%)K�w�┥'��ff8�̢�uUT�P�˙��)=����R��	����|R������JR�����)JO��˸f�Z�ǖ�����n�:�Q�r��..���z�{<�xN�������wy>����������m�����)JR{}��y)Jw���K���w��%)K�ݿ����-7Z���)JOo��#�Op�F�D��fП o����J~���qJR���~��R���z�f6f!)�	����QT��&�y)J~�����)I���ǒ�FJ_�����)I��ߴ<��<��;���5�浣Y��7��R�����c�JR�����)I��{��)߻��R�����;l�i�n�[����%)K�w�┥�뿿h|��?w��\R�����c�JR����k.�6kv�n�qЅ��r�v�s�9�6W��GA����C��H�"ǁ1& R)$�<���3ӭx�R��{��R�����c�JR�m��y��u]b�iby	�8��JR��wۀ~D'%)>���JR�����)JR{}��y)J{�{�Z���hֵ��7���qJR�߻ݏ%)K�����CJ����j�������{��\����Rt�J���ڵ��y)J]����)=��t<��;߷ۊR�����y)J^w�kU��6e�F�7��JR����C�JS��}��)I���ǒ������J��ow��7���F����PI��׹[nҧ[�T^�f�d:"ꂛ�I�M󾋦�Kz٭�3{��)J~�����)I���ǒ������JR�۽����yY"C�F�"��y��w[3�<JR�~���)I���C�JS��}��)I��g�m��6��kz޵��)w�w|R����{��)���R�����c�JS�}ӛ��-pM�M��Α�黵d��n��\�)I���ǒ�tJh KB&��20��@>.�~滙����ޭ֊n*�
���鸛%)N���┥�~���%)K�����(}����R��7��구����:�W9�Fg�\�"jl��8f�ܘ��$k�������9�^C����m����ly)J]����(}���^JR��w�)JR~�����z�5�U��-o{JR�{�w�?�������ly)J~���8�)I���ǒ~B���w�kU��6e�F�7��JR������)���R��@d�w��%)K�����)=�Ӷ�Zֶn��[���ǒ��XO߻�ÊR��w��%)K����'��j����򙀙����H��uT�����L�'�w�JP�g?~���JR������)���R������<"tCDa�!DG���f�j$�貌 BC�y�S�$e�&&8,�$���e�(pP���ģ0���X���@mO�W�Jg���l]C|�|!�d�$"�]l��fc�
��c#�[��i#���<09!zC��c��0�ad��`�$8��d��+$�����%d��4�� ��Lp�-i�����➩�7�O�iXe��!`Ls(gj���ab�0xm��&#[h����|Cr#�&�H�L!�4�� ������Gg�+��0xl"�4�� �&�W7�) ����#))(@B����J�g�a����H
D��I$�@���\A��n��+����\���v���ݼ�q�[k�D�cn.��b����rlv�ʆݍf���)��H�$Ht�,'6��z�����V��I*c) 
Ҫ�p&�UpqH[��)�T�-cn�j$�kl ��7&�΃mMT��.�w�j��s� jiW�ÄBi��Lx�6�&�;��J�mW`�j���Z9Jl��m�5Um]�+Xx�%,�-{�W�����@mm�n�g�n�9L�n3���W�mv{U�i��v�iA�c�]GEey�!n�+��u�� �}�?|^"��s�N�������8�nrǚ�Nl,����,�ӷ!ۚ5�Z a�3ËjA;z��k�<͎��W�-�s�V��O������':un7U�cF�O�s��61���ɭ�v�*�a��5��A����"v#+7b�!;h��Z����Ɍ͝��'-vh��mE��$Θv���
�s������9��]�<Yx�8N�M���`$��e�gk\\��U��6�l�R��25r�F©�`.��]��&�H��vN�HH	�N�Փ�l��v��&��ݵ���#H [O�N��{�!{��k/ ۲Ys��e`�=�:�����.2c�8ō籬�&EJ'�";<cb�u���f�����Rnt�R�W�brkmZ�fc5��u��͜cK�hg (�^@��7bYm��(N��{��|�A0���c2m�j�۶v�B��e_U�w�:K��5��δl�	�H���Ǳ]S���7:08M�qUmUUQ�x�'oO��js�l�j�g�t�Wc���Í�v���nQM�p�jd�OJ����{�lo
\v�&�һ��ݵ�뮴�mW���u[]]��	����Xh�:(�(���&ͣ�7H�u�lb:\Y�TqjH,�v�we]�y@�۞������&[1�7m����sm]Pvp��'���mUVǜ�tH>�c����p2m4(����?(tw�7���J�N�u����]m׵ԋlq�Y.�<��cj�tl�\����n�\Ձp�*t�sN���]�h������6�5�<&�#�W#d�.e�	ny�C5l�qv�8K��
�G�Yݶ�d�z�^�4��mk��_Ǐ��-�nu�d�q��J����q&ݗ:��5�ڒⲹu��(��\���ӷ2�3{n�q<lݢ���{�����|s�>��5gL8��$;v��&҉�]N�KɁ��\ZX�q�{�Ow��۫s5G{�{�J_���|R�����c�JS���8��%)>�~���JS�{���El�F�3{��{┥�w�G�+�!�O����8�)I������JR�~��33	L�Lf�֊n*�
���鸛�?~��R�����py!������;��������M�01�s�I6����[�޷���),'��߰y)J_�w���)C���ǒ��~��"�`&`&7n�N�*�DT[h�ډ���/߻�|R��� ���l|��?~��R�����py)J}��cܳ��^Mݗ��l�`�a�dg�p�r拢[�=v�랴V�)��E�V�T�TT0T��00=����)���R�����py)K��f���`y���"m��k�c�JS���8C�<N�)>�y�%)K����JR�߻ݏ$�B=
&��̯���m'QUM��\��I������JR�~���)C���ǒ��{�xqJR���>;l�h�{�o[����J�	��w���)C�~��R��~�)BY'��߰y)J~�l["�&�$	�黙�����sO%)N���┥'�g{��JR�z���<���p+��b�Ҙ�Eq��RȂ5�<1st��s�,�n}s]�)55�Zs4�z�ǒ��{�xqJR�߳���)w�w|R�����c�J���{ե$i������o�`y���g{��JR�~���)C���ǒ��{�xqOʠ�)C��w�oz�7�m�ލk{��R����o�R�>���y!!ꨘd�{�p┥'�g{��JSΟv��fk5�V�F����)J~�v<��;߻ÊR�����t<������-�<�<�W�܄Ƈ��/�{��|�>���R�����(~���O<��̾{�WS��	�D�a�[�>X���%;�8����ۦ��V:�V]��Ir�ַ��kV��[��)JR{�w]��R��~�8�)C�{ݏ%)N���┥'׶|v�Z�V��޷���<��;߻�)JP���c�JS���8�)I���wC�JS�}ӛ��{3*�Z�o�R�?w���R��~�)JR{�w]��R��~�8�)I߳�ս�3F赻z�ǒ���~���R�����_�<��;߻�)B|)��aa F! M� �p�{ݏ%)Or���3{ݚ�f�y��[8�)I���wC�JR�~���)C�{ݏ%)N���┥'{T}�Qnٽۮ���!`��h���`�9���sa��'s�����4�ݨ�e�=�����o{���~��~�R�?w���R��~�)JR{�Z��<��3�Πމ�ci<����)I���C��BC%?~��P&`&;�n�M�00fw́��N1Ӑ�X��JG�[�s@�����f�궽��E�N%��f��5k�z��mz�w4^���1��8�R= ���=Vנ[�s@����癙��S�!�hld�0��S�홱ez�Ñ�]m*��s��Aj��4��^�^;^������i+��<����R\Í�RU:�s��������� kt�_c��u����p��w]�ę���n�r��8��-Z\�pS[�6zү^g4B���g���0����똣��x�{%[�܈:u]�ŵ���U��xgʒ�_�w}�;�����l�F.r�\�ٲ��n�����	",�N�7m��ٸ�����]�G'U��޻��կ�<�? 7s]��YF�:�R�K���u`fw./f&fb;��j�7s]�s3��w�T��x�����h�V� ����$���Ė��`6~��u�n� ��v��vgr�����[�`sc4*�*)��*n�9�����ߣ�:���@-�4��r�"Q��!;�-�v�(��ٺ�ґ�q�hD�瑶߾�l�a�ɌhpjI���nh� ��=�����#u�BT�%J��9���g�fg��f�~��޻���33Ċ�W> cxE$�7�}��h[f�m����@��=ǀL$b@�Qɠm���h�Y�a����7k"����!*dT#�@����jנ�4�l�=�Zz�	��C�B�0m��B�m/+��Rн9��u˜J��i��	���8���jנ�4�l�-�s@�gV4�3�r�-BUN� ��w鄃7u���;YYV2;�U�L�DRy94��@���'�ffnd�=�]z�[4�|���d�485$�3;�:Vb���ؘ�K����_/�Ēr$�j1I��;V�[l�m�@����|cm��701l���W���v��nt�h��Έ.fe�Y�2V�y~6$��#�@-�4�l�-빠{õh��&�)rh�٠[�s@��w4޳~�Hݬ��I�D$ܐS7`n��X��s@-�4��h��ڒ	��QNf��w4޳@?[f��<t>�z�;�9�ʽ�~��3z���kr�-B3���`fc�3;�:}�ܫ�@D�ӯd٭�eY�3z닜�{=��{0�w\�g��gz6�ɞ=3s�՞\�Q�,����=�女o]��:S@-�4��9sƇ���v,t���3;��>��{0������ĜbQ���gƀ[�i�x���}4��nh�e2x�1��9 ����٠[�s@����/Z=�L$�Qɠ��@����)���xa�a���ՕV�7Wn����ӧm�U�-b1�҈� q�<�m�i���˶��87���,k<<H�H�6�#�j�N����c�1����1��Zݺ;o��z	TKX9���k��+�����yYPa{&��
�턌væ�v�`�s��ȋآ���+Z�k���E����i�8�)�lăX�9���p]Rv
����mv�v{k�B1��Ƚ���L��vצPa�͋�g��nd:6c�#�98��4x�M ����@�˪jH&��4�8���u�`������v�mŁ��U�G���<׈��>��4�l�-빠{N��?e��o5A)��h�٠[�s@��)����w)NA����rM޻���M ��; �f;�31ڌ�
��T��Ɓ化�q�C���խ�e�s��q�Gyd�"DM5q�F�ds?�|h�f�_m��w4
�e2x�5�z��ow*�߻���pFֲ����]��t��z��0�a �X�Qɠ�f�o]��t��[�h����6c���94z�hӥ4޳@/���.�� �M��#���=�,ZoY���޻���T�әS&#�������G"g��վ�\`���[�]>�\��eb����NS�P�6��o��g{����\~����v�]X��aUE�$�P�6��Y�[�s@�����f����(}�<lp�@�����}c�yڥ�3�=C���9��A�`8�8�MR��K74a z��^�Yi���,�INh4	f �Mp�FH�ec�L����BAv^��z�p�H6����! �$� pO���M	�`@A^�b�sjF#6��+e����T�R|^x+Έ�����A{(�AM�� �WB��'����T@|����]���*���T1'0yQ���=��zoY���޻�^���<oS�H�޳@/u��w4oK�q����a+:nw`Li���W��Ϭ�ٲ���As����P��k5��������@/u��w4oK�[�h�q֖G���x�"rh۹�{z�4�f�^�4\����i91�#���=�vm�@/�f�m��˝X�M��S���&�> ��v��[w430��Š{����	S�d$��Y�u�s@��Šm�{Jf�Q�m�Ȣx�F�!׌h:�;�ae[� ��q��r�Em/;V�^p$�@�n�ץ�@:�4��h֪j�$��S�4�,Z�٠޳@�n�W��L�6���rE�m�}�4�w4�,Z����&)��"�M�1/��4��s@��Šz���:����d�$�ɠu빠}~��_�/��]���c�BI�� D�B�m����D��nNp��w��۴� ����Q��L���bmn�f���oGH����&�5�K��Hc\� \հ:S���m�=�#�Y祫c �]m��E�O���a�\G����}[<���X3��.u���t!j�kG`�.{cG���Ӈ�z{({l^c�.2�6�X�d�v�J���C�:�3����Ur�0<VC�zm�(]]��{��}6Ƀ�u���s�q]gOQr]�+ �����a�smv[�(J��\��ͷ�����u�4�l�:���=^�C����u��5$���,'d{��ʼ =&Fn�v�����|eА�x �=�ze^ �k[�=�nW��:��WVҶ��=2� OMkt '�x ��tv�Y) �J�ݎ�۫��Mkt '�x �=�I�x z�^�WE�-��a�ݦ98��#8�޹6�Mr���K-�f�㎵md��˳�t�Q�� �� I��@!&U��23t�'�Z�N�ՈCc�� �v���Ur�s��Un��e^ ��� 	#x K�¢���>&��{��*� ��� 	#x �=�	pp�m���j�M��W�o.�,� �7���� <{�W�o��Ս_����
.�;� ��� ���BL��c�w�=�R3��Yv��������8�v7
���z;^��s��9�vܖ�����o@���te^ ��� �7�ܨ�h�էEմ�ote^ ��� �7�=#� GT�%$�v�X�^ ��� �7�|�Qʪ\���s��P	�<�E5�w����33��yW�^��|�JӫN�m�� 	#x H�@!&U����t�'YV�S��()6;m� I#� ��W����t $��w[) G��0���nŴ����X���tVq�h�ײt���ق�Ss!�yڻm���?���*�l~��@=� OH�@!%э���h��۵����tKx	��=2� _�D���|.���� ��� OH�@!&U���;� �]�J�@�ˡ!�� '�{��*�%���^��4-	B���}�*�:}]ݚ��&&�94]����=� �l�?eH�Rō�Lr'0���Zy٢��b�� \�^i��9���uqVT�`�h#&4��?W�=�mzz���~AU��~����df)$�=�mzz٠r�^������&\f224�(�����Z�ץ�@�[^�}}����G�H��9u�@�_X�U���f��֍�117,�7��������~�wʾϾ�V�
A	"ȫ�<��T�Ci��b�a� �ɆL�P�y����BI�x�f�ٻ[IN[3�v}ayW��`��5�;c��}�g�����ud������G-�9ke�G���ͱmwm��9U��Rx�šӒ��`��n�	��9&�"uu�7!؁����6���.���5*�j��ۖ��5��Wb;c��9���ly�e��Ǉ�{n9�v�&c~����m�P�C�k׳[&��j�7cn\�,��]�f:b�[��Z��7��86ߧ����ؽl�9wW�~��z#��ڀ���@�� ��;�LD̤b�ڰ9���@���@��P�Ncj#8
I�r�@�_X������@��5p�h �q���=�mzm�@�ֽ �N����f9$r=�mzm�@�ֽ�vǠ{���n��͠���[6��Y�"Y��v{za��[hE�s�\�ӧ��L��33���ʰ>��u��V�Ձ�����w�V�N���{�W�w����*����Ǡz��@-�oؑ~�捑11U2��6�n�j���ʳ�)��@-���:D���x�j����W����`�c�؈]ݽj��b�aP�F�)�[�h�31[���;����3*�&9��2t4��p�n�]�us���m])c���Vҙ�.��s�ۏ��{3C`���C9? [~��݆��[^�_m��������2)�$۰;���٘H��ڰ���~�3����x���$NC@�?~��Uw��|�����w��_��޹2� �H����3	ow]�ff������V�Ձ�?����<dOń��4���?�����־�wj�3;��� �aT�?k�qۊ�vFr��9M:�E��0�u���sx�rB���w�~�}C��2��m����b�?+k�z� ��4��dn<�7N��jm��qn�_陏�A����}���@��@�z��PFF�&��3���;��f%,��u`qn�X���6��Crh}�g�[~�Wk���y��u�Ҙ��+/�U�s��9C��Ĕ��I��8���Y�����V�����`�q���O��p�7��Y#�;\�-3�i���M��iv�M�q�b̗V�m��ۛ��#������٠�gٙ矐_��G�u�&}�dd �G�_s�"'�3T��`o��u`|�2�묭�#�F�XI�@;�����͉���K�wj�7����fR-�B�T�4C�T݇�f&ef��V�Հg3��b"ba,��`��T�?7I�֬JH���_m���h]��ʽ(|p��3 �@��q�d�~����7� e�d���� F�| ��Dv��kC-	0l�H��=U�0M'��T��L�t҇�b0�J�\�"e�����Jxp�p�5}��!Y$4��C@|�)�$$��D��j>p��!~'hx�mF� 	G`�����K�	�Jc M�����C� �y������I� I�;e���H];N���
3pj�"֜(Ԏ:5k��h���-V9<sS�g�㰇h����Yv �k�!�I��8U��(��ٖ�<tfT����f����-�JPf�I�u���tp��Z"..�6�d����� Ҟ:��W[vi^[R����� UF���:ب�,�q5˖��r���5���ρ�6�{ U)����m����f=v'�`�n'��v&�s�An7�:vv$�<:{r]m��Gi���t��F���;r�[h�$k�E\��Z$(�eԛ��`����3s��q�����:�c���6^�i�;��o-K�px���S*nSs��v	�ۓ=v���d�7l\i���C',cnp�q��kx���=��;�;kv�ϖ�N�ڧ�c^ŝ3�;		�Џf�l&�)wD���5܃B�.�7�{N�@�p"�h,�i޽y�:K�6}v�<q��qvH��H�fqٖՎ��CF3��W]aZ�9���;v��;�,n�.�s϶�8�����w.�tӜqZ���M*�U#�r$�:�-�%���Yr��;��ʩ��1���TIc����ۈ�n�0��Z� ڗ	��5Yi��g[�s�plN�s���\��e3r1�i%�fǌ{�l8�6���mM�1��)s��l�=�r�l�Xvvr�k����t�l۠���>�� 3����Pn�ջ�շNS�#�^[ 0&�v��)]�s�Jk��ȉ4�����yV�V�Y��ѷI9oP�b�Yg�����2�����C��XbڲXP�h�ʵ-Ld��D�R��iJd��.��s%k��x��T�\c!8n���a�;7M�W*܊�'�!)��m��3Q� ��}U�J,9��X��P�@�u�����G>�q��'{Iq�� ^�+��zڷj�.�v����U��rg����m�H��zͭ�4�.o~����oH
��Ux 6��>��p���њ���g]x����8���sŲv�ѹ����d��yӲ�P*Ҙ����fN�k8�Ϧ<W=zy-v_m[c�ۂ��g���&��̛���M4�c�Ɠ�&M�.ѹ�a�T붷�ۮu��q�eW�u���%��I�vۓ��Kzv�\vL�M���a��x��8ا��=�x%w4�Gm�nJ{j9�%	��{u�7����wn�\\�N���m��^��x���3�S;����������sm}��FF�) {o�@;����?�bfb#�[�V7��T�8T�47&�wu�׫��mzzٿy�L�BF��[@%N):j�m�76���[^�^�hwY�/S��f��mӰؘ��\�ݫ �� �{��b&e,��vr�� ��u 6��@/�� ��4��h���{���I:�"���ndq>E��k0��Ѻ��qM�-����=s����w�x����9'�o�@:�s@���@/�f��֍�1cMdidq�4�W�i�F��过�/3��5ʯ߿~�*;���x�w}���y����Z�8��9{�`����Ffk���v��k"�q�26�H���hwY�z�������=����dC�nK �{���ך��8�v�9�v23������I�<�����3���Sb�&]�#ձ�z�Gr�3ٴ�2���ۦ�`w+����feXfc�1�P��`��Q4�m��X,̫�̤���33]��Vc��F,�Ax�Ezz٠�f��y��0�1$PĄRVrKJ����X�����]����8�	$rhwY�~��z�mzz٠u��=�<i�SnM�}c�?�}������f�}��-�i̙$�Ʌݹ�ݩ�c��L�W��O������3o5�QsÛ�i��Í)�Z�)#�_���@-�hwY�~������q�26�GV����$������噕ɘ�<�#���	�2!�D)&�[~��Y��و�Uu{ޫ ���`}��c CdC��M�.k�u`qn�Xfw|�Á2��b/�� ��|������x�LȈ��G#�?+k�s�w��`}����٘�暒��i��a����7d��Z�>�ؔ�v��%dt���N��8��2dfG�H����}���@�]�����֮V׋��I6�7`�q��LL����ug�������hmi7�k�G�@�WqՁ��ʳ����33]��s/#$�8��<�X������= �l��C�{��G����j<FF�)�^�hwY�~��z�mz���Y����ݭoZ޷�0�`{�T�v��Ⳗ�=#��۶��,te�h1����+�t��ۧ�v{>�	bxG����2f�7��[ ^����\�9����.�Ѷ�� s!NFv6qA3ô�;�}p�Ρ:uI�������^C�=�[(۲ �,ЇXn؎�9����؞�֙�1���g3�m�v�m�n+� t[�R���7�r{���[��{ju�-��1v�Aa�Ʒn�ʽv39J�tu%=Em��n��ќ�7���`}��u`|�2�&~@nn�߾��!��%$�?Wl{��"!#�wj�7w]�w��~����634�x��0�I���[l��f$wW �]���\�0ƌ~6�P>�3�J�f�w_��U��궽��emx�4 $�I����333���W�un�Xfc��$ �ʂċu�Y��$�(n��ʽB�1�ki<�bÞ��K�)"�f)�M94
���U��w1�b&g�1�w�vo�p�c��9U
t��:�v�LD�A��v��;{�_��31Tjմz*���6�H���������=�mz�܃��dC��M�����3�[��<�|U�ř�`����1�m@�Ȥ���T݁�;�X3=���>�呂w[4�j�I⨘)�f�q���#`$8�޹6����N�bdUhz�1�x�L�6��궽 ��`�c٘�����*�ܥ��l:� �9#�m��l�*�G�qfe_�b""#�35G����JT2�! �t݀n���ŝ¬么���m�����hmk\�4�F"8�3��4��wj�33��!,��`fV�t3��)͸N�_ջ�`~��[�����`b��Vrq&	,�}�����;���xy��%ɸTn��G�{$��9�v�'\��kқ�6������`�s��VVW�&>Aջ�`s������j!�4�ٿ��<ċ����[�V��;و���L�Q�y������(��@������궽 ��hu�@({h�13$I�C�3=ݫ ��v��;�&f%������+�@��cfr8����= �l�6bVf���[�`qfeXw ߛ0��vn����mU���\X����vݻgH]�mq!I�.���zv�Z�m����`w)w*����ٟ���`f�Ҷ��5���9&��k��=Vנ��`�c�DLDǢ&*�[�7I���Nm��$�|�߿U�g;���3	������@�˝Cq1"y@�z�<̄����37]��R�U��fev�v�lkU��6P�E&�M�{������D�ַ��1{ޫ �w�鈙�l���e�i:qy2iy��5��,a�d�|x�����]99yy6^�%�#+vv6���3���h�}x��z,k�:�+<�ƞ-�f9�ZTl�xQS��FGrԵ���I�u��b����6��m�V�,�kc�؈�XSM�e���g3֎��n7'���f�9��*�����yÉ�(6š��bu�;�[h�Y:���y��>�� j܏�9���֛���i����J��+8\�#C���jg��u$�4Ҧ�v��XY�V��?D��������߄a�ő<$�)�ř�~����H7���37]��R�U�33�;�g�X<"��@>����f������k�-j�Mxd)��I4�٠~��z���6&&a-�k�3um:)R���M���נz��@/u��l�=�����rQ<�����7�9��7.mg]A����RY�n߽�{��ﾤ��}n����%~�W�����Y�����נr=�a�H�F�)�_z���&�%a@�;��b��n��`wk+j��fe_鉄�lc��uM��1��$�~�h�ν?�<�3���= ���h��x2C�QD�v�]���3*�3����13興������x7c�A
����n�XY�V�baow_�������X3����d���,�Bskf�<���*���e`�'g�aË�S��-�����{�n�t�g��?@?�����f�Wuz����\�����I4�ٿfdLJF�ͫ�wj�3����d,�UI!��4��I�U�^�궽?y�a�!�4���A�*�BD)`���ɃHɀ�a�f�$�����D8H���'4��f !��S2hB_K2p��@0���0�"��Ǭ��e���LZ̳�("h^��v�|B��C䌘��"bbr3"��n�;��8�1����Cqc��t���DDDB�{ޫ �����@��������D�6�7V��v興����En� ���z�mz����r̌��^�'c�O+��j��ɞ68+m��-ێR�r6���t܃&&���M ��4
���?+ml�D���������R���4ҒhwW�~Vנ�� ��7���&R��ƥ*i��uUMՁŻ�`�� ��4
����:4a�#���n�6f"!-��`�����ʺ�U��(LS��{�r��_k��'�A%�$nM ��4
������w��D�v�ջ
r *!A�ta���r��o��np%��mr��{>Zi�?������Hi�(�z���@�[^�^�4�٠~W��d�l2L�b�G+�:�v��1�nf� ��v.fU������H�FД�@/u��k�fba-]ݫ�[���9�:[����)4Sn�舙�K3u���V2���""��v3^�P����T݁���`zfb{�u|�����w���w~�~~��uC��q
��8���s.0Z�rg���v:ٓ�;k��a����6��K���ۺ����mm6�x�N�^�Ý�6��a$��]��[m�[#�u��|�'G)�O�M���lѶw=˯j)�!c�K1�w����nvq�nDu�Z��s:(�nS�U7E�Y\�hΜ�Fu��*���6m��I�+]�LAu��󳫞W���\��-��]�#�q�v��g��m�znT��A��2��3�H��CU	6�6�z��`���1�#���Vv�T�#a�X�E�I�^�hu�@��Z2���DO�""j�mmz
�!��m��w�vef+�Y��33��q]Q��ӏ�q�4>����}���w�[�hu�@�m�,��I8M:���[�����D-���f��-}V�{. ��Nb@�Q�%�g��Cc.�:�����7��:����/7.e�i��m	H��l��f�y�Z�ڴ׈��܆8j"94���>SD.��'@��?*��_�k���?�Z}�h��Y"�Q�Ҧ��w�̬�f��L�F�k��}4.^ʱ�	�RD�Z�ڴ;����v31+q���#�#��I"�����+~�~���h�j���P�uG�ő�7sC�_ps/;=u��G:���E�� ��~���H��l�/;V��Vb�D������vn��I�T*)�CQG$�/;V��v� ��hu�v&"fR8���P�~P�Yp�uM|z����Y��3<H�Y�_]�@�{���m$���$ڰ�L��[���37]��ǅ��]׺�n�êl�aE(�$��f�}���ڴ�Y�߾�����~��?�+��Dq˥5��<9��U���պ�m���[��!OU�_﻽��~c�8Q''�_��h�j��f�w[4��*�7'�I��=��W�)�k���`g1�~��������ϲ8ǉE�I�}o�@;�;=2��^�v�U����AU$&�� ۪n�;��`g+1X��VL��� BF�<� U�s_����=��WEb��j(��ڴLw^��s5�{���� s��	��YSl��3�÷����5���/�f�lt��1S��jIY#3�$�qj�����- �����Ɉ��G(=��+af�1�m"3"hJE��� �h�j�=��W���U����"��f�;���>��Y�~�����(�94��U������ĭ��\�b�D<Q	Šz��@3��`�q��ܫ�".& &	�����w����7f��E�
A�N�q*�g��1��<��7-������g.�r�bvn�q�����9�OWv����tk�ŵ4b��m�L����	�h+�:�f�w 2Kq�׶y��9{B����ܳ�;4ma{<n����5��.m�u�rԻ��zl�a�>�'m��Cm�M$/uN�]&�c�^+�ӵ�
�띜�b�ư��y������o���[�g����s��/m9�y�.�r�Gu>:�!&F}���/���LY��_����h{������;�~��A$NM ��4
�������Y�g��E��_h�lLq�5nMWwj��feY虘�����`������bLtG�qe´�:�=3?�f"����z����@;���mz#����LdM������f�W�^���^����M'1Ȱ��q��c�ܛ�x�]'��e^�p�Q��ej���6߾������ 
'$��:���*���=]k��Y�~��do0&
8�NM�w*�931;2ً~��{����zC�ʱ	��x�m��WZ���h�l�*���.s��yr8�I5����DL�bb*���`��1s��*�ez���߆(�ƐI�@9��`zf&=3y���}��q���\X�fCm��nD<�i���ԯ,u-��{g���k��%�6�[��lJ���Ƣ�I�U�W�z�נ޳�����f���Yp�'N��7j�Fg��}��~�h{���y���P� t��3��`�c�bf&?LAD0�;I3O_�7�����*�����?^#W"r�D�h�l�*���=]k��Y�~���k0��J��1s�V�"g�1�}�����h�l�=�\�x*ɂ���7\���O��M��N�STf��@�y�+`�E�X☞6�z��z}�4��{1 ��j�62�R�a�T�QdNE�r���z٠~���=�j�DD��FeelRBi����T��;����+�����%ܭ�`b�mX̅�%�� �9&����@���@����+� J�
�w�����{����f��7��_����h{�h;�������N$�Fjwd������Mٕ��q�A����;�]r��m,�q�����'�*���z٠~��^����r�U�����j����I4޶h��yڴ��7��3��#��/�o0��I4~w�{�ՠr���z٠=�,�)�� ܋C������>�h[��z����L���`leh�l:h�&�'"�9wW���@�]�@���B���Д�4C�Q���:�O� O x�_�!��@xy�N�I�Б�ڼJ��\�D4�Ͱ���	�� ��S17	��ا�� R�pC�$&�8'��6���C[�9�\P��� ��B諘`L5�6�M�5���zݼ��k]V��&vZL�==�q0 �B9���9.];�;�����GI�j�3*rN�t�[[E���[z�%�M��	�`KM2I��'����B�l��YT�əX.��+�8�Mp[����B�0R��<��6��@�<���T���gq�j�㍊��K��P�N���J�g��$����&��jV�����6e��G��6�6��*���ݰ�n8�"=v�7N�/���ۘ��9�6w�R��ڏ\[�5�k�.��y78�Q�]S��@�ɩ���t��Y�HQ�������u9'c���=ð����$t]��H�����:^k���d�s�T�q��{cqͦ�y6�8ä���v���4P���lm��5�� ̶8㝹v��[C[-dM�����{mú],"�U�k�;Y�m���������Z��.�IU�Z,bP�S�6��&N5Ԥ�.ۈ�v���v��c�L���=h���iwaʖ�V���S�F��u��Fu�Wi=���=[�#q��K�8�8	X�8�ѻ.�Hr\�=��v դ�̢�*�T�'X���Pu�sC.�6�s̮�����ր�x�L����n-��[�s;pNC\�^XF�d�\���v��B7I�c�,B��a#�������k�v��v\�mBaϐ(p�ڀ�r������0Eb�Z�6�i�J�)2�m�WD+�l�w#)�v��YԹ�f��m�[. ��U�8�dս���魌�D#K.^�@&b��T ��I�A�Nk=�ۭ����*4h���ݦx����]uX)�+V2�:�� Wlm�ۣ+��+K���9f������GM��Ѹ���bk�@�зd3�1�N�\�PT7N����ѣR�h1�*��+�����QIH�tλJ��v�J�z�,�Wu <�c�����p���˃9�9=["cvUP(
��z�T���`�N����n���_DSk�:�6*H � x�&"�� t�*���վ�G���^9�:K�p&m�v������]���v�A�M�lsc�k����^I�-�d���l�[3����pމӏ&����5�q�������ǫv��\s��X�׋���R����v�Ύ-�IхI�;�3�K�oX:���֭�(lm��k5C��@�:�f�
٫Qv���}8�v�b�*Dz-q[nIg=�t&N���� Pۻ��^����Q���n�7d��i�'-T����+m
k����Է0o��An= ��h��h�f/G�""&yA�w�`g�֒j��L�H���Z��Z.����;ؙ���H�wj�7D~n.Э�S_�^�:�ܫ �s��Vb�:�v��#mDN-�y����~�hef+�31��uX�-���#����@=�f���V��;V�˺� ��^e���C"~?r/�7[�����.W�bK��hn��~�����E��/0��I?���;V�˻+�? ;���4;�(ӅP6U8�yڵy�fbG.��޶h��o�bbf62�P�64RP�6�V��޶h��h�hϝ��DDq��޶h��h�hl��D��ͫ��ۤ�T�&�F�94�ڴyڴ]���l�?�33� ʾ��dhXE�
8��L<�6���V�l��s���S������������y�����
�U5�7���:�ܫ �s���?�ZGW��œDN-�w*�9��`}���v�����H�`�}�9�`���z�女��V�0=%B�@�A��F�<�+���9U���LIC�^$�y����� #$�@�]�@���@��^��ff}15Y��{QM8U�r-�v��uz�[4�ڴ7��?��}��b���c郱ν�O���R�2��;y�u�v��u��߽���Y7n���'"�V��޶h{k�=]k�/>w�Y1���z٠U�ʰ8��V.�*�ba#���hi�l$lt݁���`|�ܫ=2��ͫ ���@��Wq�F�ę��F�����V.�*��s�V���fg�DK���XrU�LdMq�wW�~^�z�ڴ�ޯ@3�v\2�ć�0��u��z5��s�f^��;���C7�v�n3���6	�NG���4
����;��? ՙ�`sq�T�
Ҧ�\̫�0���ڰ5fmX.�*�"f"=A��xP
)�
�n����w�`b�r��D�%��ڰ5wv��|?�#���Y��wW�~^�z^���ޯ@����D"�Gu`|�ܫbb'k���]ͫ{�eh�� ������u�=v�C:W��#��@��l͈��q���<�i�MF�s�F��a��g��C���gS�����m�nN6��F�W^�8//:��u���G/@e@��޺�p5v�q�qlgcg��8x�g��:�V3���5S�����9�������@�Y��ˎ)�n]��Z�GU��%ac�c/S:�vz��o;X�Pd�`�8/cj֟	�1�3�Lv.����d�L�u�6N�M7g���NՏ	�8�W�{��wW�~^�z�Kwdo�L�ģQ��W_��W{�`|�ܫ3*�3�բ�[�'�q�+~z��W�U�@����/��W"r&�9���˺��mz��^�Wuz�e�<X�a��Ǡ_]�@����*�@����=Y�bM$��cR6�o�!'8���(��Օ[d�]%�@�Os�,�����ls���ӑh�uz]���uz^��x�~/&GI(��=��WQ2��&	��TR�r�]̫���X�;�~%�kn=��@��V��wW�U�^���T�0�<&H��*�נ~]��wW�~]���-�ND�9������[��*�@?wY�U�@�s��cMLP��v�Qs��>�vt/VJ7�ln��.����s��M�F�Hؠc�@�z]���uz�ڴ˺����NF�m��$�@����/���?.���Y�l�Fʺ�L(j�2��Jv�1%���y�gy䅷f��wW�}-	A��F��@�����f��wW�_]�@����	���J(�@/u���^�}v��>�@3��aP��v��eq��^L�鸳��;=uˋn�t+nHz��v�V�}�X�R��o�����h��Z{��:�r���H$q��j�q#�t����Χ虉��H��eç)��&�ӯ��W��9�v˹�`b�r�������)���V����^��/�o�w�}��x���8*,�,)B(�D$TdLQ%@�͊Y��ʻ���������M��^�}}V����`��==��E�)b�M0��qƮݞ�Np��e��^ӷNkX1iJzh'�fb���Ȗ,���'�W���=��h���?s�h_N��!�Ǐ$iȴ{�4��h�ڴ����3ď���0ɑ��J)��}��~�j�/���=��/>w�JM��"rh�ڴ��{�,6"&R��6�ƪLA���6ց}}V��t��_z��;V�{��_�7]W�Ɇ#;X�
B��l��njz���5�йv"����:���u���y��ɲ�R8מ�q-��V�z釮�1��xF��q\�Q\e�<v;�����˴ܿu����Sj�	&8��<��ݝ�q����bf�R8]v�7�S�c:�lQȴ"��S�-O2n��<\i yc��K���%g�R|�5)��{�������0��e�f�uOi���.G������y��֙�\F��a���	�9��i�QH��>����@/�]��k1&f'���V#j2�[Pӂ��17 ����v������M��5r7#���I&����@�WqY�"&=335Y��X�|��,i`�A#"$�@���@��S@/�f����@)��C��Hӑh�^�f#�35��>ݯyX��m����pu��7��f��s�y�v6���㱹�糫>:�s�l�XyۮX@QH�4��h�ڴ��{�4ϝƞy�$NM�;V��;!�RX�
z�����������^�{�K ���b"!#�KcU& ��pH�����ڰ9μ,ى����h���~���̘����"'����f&kw�~,۾v˙�`b�eX�W7\Yr(��4�Y�~^��
��������2�F�sɓ���<���8�9=u�{fIN�9�%��C��Fz����fTkr7#���9'�=]��@��^�ﯪ��f���j�cs `�Dԏ@��^�ﯪ��f��{k߳��*�����x�F܏@��g*����,>�_q0A¡�e�	L�2`��d�[��ٰ�X"���� xXF,8`J�A$`B`��#�&�̘_��y�p#,03,,��0lK�&lK1�'2IqBq	�'� �$�q�� �K<C~��r�ͯ �곇��tT�#�����I�#ĉ=ٽ13�|��=��ؖQp}��,,|�s�Ժ4N�7���=��eĒRa"Vo��y��5���	C��k	hŲ��6HS��VĄ0�_P|6b�x�!	Z�Bh �"b�f�� �@�@a�)�&$2�#f@�DL�)�U$^�äa2D8H�xiK,BsI`����OT'i�|��C�6��祒LaAccca��E�#e��KC�oov	����i	�l��+ȉ�v5�����~��+��aO�=_Q=@u@ҩژ�fg�)|��j��k1X�x*���M$��ȴ��@������C���]���__��B6)�h����h��� �l�?��{�v��c�bxܢ�a����Ř<���F�/m\��RڱS٧[�K�,m�48m����V9]�`�Ǳ���V{�`f~p�*wbCt鯀�������נ{]�@����qdp1ȣ���f��{k��33��-�_����\���<1��a�&fbW+��`wkuX\�U��1�yء_�M��5�A��2)�&�zv�����Ǜ����v˙�`fl��=��]����kX`6�>�c��vax�^�SWBó�1�m@1,�iL�#�h�z� �l�?/mz�j�/YD�LmLhQ��zzٿfy���Ձ�[���:�DBGV�ªD:�ǁ�D�������@���h�f��j�MA<s	�H�?����j�;��V��v˙�`s�<p��T�7M|{Y����7_�qwk�w�w�ʿu$^���H��
tOW0��&��a��5e�h�h�U��U#S��"��(����G<z5��n]%���= ��8�U���n��������uuc���K%ɞ|�):�����l�Nū#nW���u�/��t�f蝯$�Ǝև=_�Q�:ny�_a�q��p+�n�[8LFk���	�ܦ�(�U��A ���̐��������P���v.���Q�uPvS������>�����p��;��Z��)��89y�m�筭�HA����9F۶��j�"�����@�����W��3�]~z�T1G$�jrh����h�z� �l�?W��271�E1A7�yڴ��z}��_���~Z�V��,�LX�F��@��W���z���h�J'�2cjcĢ�ȴ�Y�}�y��7�������9������zd�I��/M����K͓I6�n��Y�]]3�T����&ё��<R&��;��h�j�?+���@��r���=�n���*��s��qBw����ߪ�73]��WqXtǂny�vĆ��_ͬ�`�q��&bR��j�=����W:F�r(ĜZ��1Wo�@�w�~�ՠ~^��������<�9�ﯪ�?Wj�?/mz.�����L�Y!�<Ǌ]�:qSkvv�F[b�k$�lqq��X������_k40Ra����_�����@��h����33? �w��[��H�
�ʦՁ�+1^��D�BF,ͫ��Չ-�!��s��S����������l���`s��VLD�݈���;V�ǆ��FG���1Ȝ�C���wK��;���@��h�נuj�MA)8R0m��Y���L�:�W�b�ڰ9��+�� Ŵ�AH����Ĝuv�v�3yvї(�WN)ĭ�R��@��mi��&�s`�#�/@�����wu����@��V�Z�؛�p1�I8�;�w�b%#���`okuXr��}�*�RH���@���h�j�?z�Z]������#mI
���1鈚�_���{�����Xl<�i	�G�nX��O��s3��r���u��Ն��0�#NE�~�ڴ������ύ����:c�
�PrbČ���	-�u�W�E�ԦM�;���m�l�RZ][��������)<�E��_���)�__U�~�ڴU뉴dxɌ<p�Ǡ{�Jh��h�v��z��W*jӅ#
l�3��V˙�g�"c�1^Y��3_���MÊ����CM�_�?�Z^�z����}}V�k�t��<�9#i'�W�^���guߏ�~�]����u��*���,)�
|}=�{�S�����ٌ�Ñ�����ɇ�q�O!��]1#)��^�\Dke��q��8�slc���R��I.Ŵ�ugN�:5˝�]��S�c����ħ5�zڶ�\+���^z��06v���'9cwi+v�xw\�ݯi:�mح�3�1��9�4���E����{n:r��A��5�5ǯ��:	��w�6f�'\��;�b�z��}v�+�ޜ�0u�χ��3�k2�b�,&���=����+��)E����L$�������/���7�!�(w��%��\�!�B-��9]��b9��V��Ձ�u�`�m��Y"hHӑh�v��z��zS@���@�z�'��cj<��`b�r�s�9]�a�+�{�����h��x��@�ޔ�/���?z�Z^�z�
�*�OE<m�q�!՗����ey��O.D�!�K�L�jdMA6L^��}}V���j�1s�[? �q�`sۄ�8�*����횒���u�Tڃ�x��o�ĕ��Z�9�AH�rF�N-�zՁ�WqY�K{Y���kuXΧ��ۏx�1I���3t�-�w�~^��
���?WY@�����Z�ڴ��^�Wuz���@�g���4\S�i�g!����ϵ���BKK��1�i�la�Q����׳�L����wj���ʰ9��.G�1f&yܴ<a�#Q�YnG�r�P?yh]�@��W�fbG.��FG�<P��\��k���w�w��>� IH�$4mN���ٮ��U����{�gJ��l�� I�}v��^�W{�a艏D����T�p�*wi")_��w�=���}}V�}v��r��h�&��a��<SЉ�.͊8.�v�\��q^Α#�:��曛�/R���S�@����_U�_]�@�����R�
D�$�bn=�_U��bG����=]��@��z��(y��rb�-�h����������T՞�5��#r=�<^���}���\��u�s���i��>���o߷~z�j0ɑ���=������������;=F�o®��m�Hs��y7S��Ύv�K�b4�vr��i�r7e7�wo�~�y]�`b�eX,�W�f>A�7j�����5�1x@�-������
�נw���=�]C���NlI8��.�Ձ���g�fe.��U��7j���<vE���$M$��*�^�ﯪ�*�^��{k�/��b#�x6�&Ǡ{���ՠ~^��
�נ|h6I��6�!2Xbc��NBc%�P=��j,�BAA��A�g����̋kz6!:WM�7��A0[VB`(�vIA$BL-.!��!�(B�@ca�1Cd2�	*@1C"I�#I�4��D�8�!��C`H���#����x�l /$#%�M@��� M�`AM�G;�+��F�U��{�N<�AF�;L����eлu�0�P��f�GV7V5��N���ܙْ�Ő.A�3է]6r��mw��L�'W��Yle'\���neLK2�\�\�mj������A���u��jZ�]��\��,��3х���Gi�8�>��e�n0u��*uWl�M5Wi<�&CN�G+�[�m-�M����i�*y<Y &���L�27l�q۰�l<À��L�0uhN�њ�Fv�;[�E��wN��Uu��v��]����T9FX��ݻ-� ::�\`�/؆\n*��:t�g�$M�j��H�rr��N����Su���3�wj�2pjG*��T���k�b��$�ɝv�olF�����@�xnɗ�-����[�ȩ���NK��Ӡ�YU�:��Dam� ̜�����:�;kV�7;9��B"5�u��([� �n�wn�c��k��hf�y��kF��g����õ�.��[Aθ;i��`Z�~y���y�s�����:��:�m����۶�4�l �TY�6��yYxWk�@����d�������tL�cV9��i�+�xN�9�쮔 �]���-����m��ݪ�y�-�:���k��u�X�ܳ�Nr=�Ź��ss��I�i�s�E���	�!¹�L;Tpvv܆�\�[g1�� �`#���e�3n�v�m��)�n`xֹ%3��n�qnyN5nӵ�Q��3U����Vv�a�.XҨZ� v(�5x�k��`9�ˉ�<1����ʠ;pq�]�+�re7)�p�mUUR��z6!0rqYg�q<��tL� ˅KvNҽ�����v�����i�ͦ۝���12U.���'gi�ٱ����'��=�8m��-b��X|�l�	7e������|�aA�VM�L�=��p�6�X��͑'�pDu�̦ �5\q����e7[⃙#6�PRvvfN$T
�$n�۲��$�	�����Y��0�{�����SH��*TTO�*�x��OߐH�l�LPA/6癭�19��L�6Y�ۆDu9�<���N�x��'V�W�v�c��9��:�m��rD9���5���3�[�[x���퍢��lOh�Ўڃ��:�s�ۮ<�^�(�7�1�ry�,���Y-mt�T�Ų����x��D�حN�=:#fM�(Uql��v����)����5ͲWl@F�J�oUK�s�<�<���s�~{��~�}��$���G�kC�q�L�xL󮅰�u�b*GC�Ʀ�*�{��3C�b#���^�~�-��נUֽ�_U�rꚳ��&���Ձ��eX��V9]�`gk1^�D����'�2dj4�rG�|��=������D%�[�����X\̂���3#������h���L�����ڰ3ilj��T8R0m�;Y���D�_�7j��+��n .�)����$p^l�</�a>�r�uMRX�⃈����;4f��7�R8����z]k�=��Z�j�W6Y!�EN=���y�����&fc�13cu����V˙���$}�C�&7�m"`�zs�-��Z�z������(A����Sp�5a虘��{����ڰ1w�Vz����5fR&��1���^�@�ֽ�}V��v��{D�`�,�!f���T\�wn�n�`zs�UpWd;g]>�Iu��:;I i�������X�w��Vbو��s�������!Cf(F��=��Z��Z�]�@;���W*j1�x@�.U�u��*��w��Gӡ@ �y!vY�{��i�P�G��6$����D��?yX��9��+;Y�����dX8�ICp�����DN�e�_�[�����;��+ ��F�����I��l�]gYq���s��ODM�Ԍ�E y�6-�rcX6� 7'�;��h��@������u� ����91G�yڷ��33=�ƀ}~�h����ѫ�44Hӑh���z٠{���ՠw�*OKj1%�CC�������;�����k��V �T�O�~��yr�W�A�B�8�<R'$�=��Z�j�?{e4��@2��Qej&�-�V��(V��sd뫆F��۴�������f�H�Ț�x�$�@��Z�l��^�h����u�9�i͉"&鯀�u�~���su��f��Y�@�NL�,j$�!�h[f��+��ى��K6�U��������Lkزrh�����h����٠~����7&8��:��`}�xXs1��w�qL���ñ�䳊�܈�u��#��ۦ�����Ӹx�V��\:�����N��#�f�cbL�v�s�72㠠s�v�s�.�׍� �ctm�닐���][<]�vd�U�`��OV�3��9B��bRkn�wg���/Z���m�X������8��(`��9Uk�1F�g�F�h���r痣�U�9ۜ7j�;���ڞ\�����{��H!^�뮸�R0���^8���67*�.k��z�3�Z(&d�ӃR`5"x�9�Ƚ�O� �l�=��ZWj�;ޕ'�Q��
9�����}}V��ڴ��M�mԓ�Qdo�$�@���h]�@���9[^�ի�5�d�"$�@�ڴ��M�k�=��ZS����{�$E#�����@-�4}}V�k�{�ێC>���8|�p[W]g�������u�܉v̰ݜ��u�I�2�Y9"Ȳx䉡�~ ����=��Z���?{e4��X��<1�,������_��g�����@��)����k(cncƢnL�ŠZ����S@-�4}}V��w���1ȴ��M �٠{���ՠw�w�&2c�9$�@�mv�ך�6�U���eX#���
K~s9�{%�ꌓ�A�[Q��l텈��f�utÒ� �g6�x��=�qj����?�Vr����el|������KcU&,$�"�/��{k�9[^�ﯪ�:��(4�đ#�/�{�~��U�w��/�l���$ ����>O�=��ן��{�������+ �O�bN=��������h|�}��@��} 7�ቤ�`�z���@��Z��@�mz���܏�mvٽ���c���6v.A�]nۘn���/�X�]l��nF���K��ڴ��^�u�h�����w���cr-��נm����@��Z{�q<yLdǄq��u�h�����h����m7F(�G�
E$�g�b��_���r�3��\�d�a�*%
!!	$C0`��+����|���>ʚ�b��DI��ڴ��^�w3��WqX11<�[D�����;��p��n{{fo/kN��4詮�%�U�F�d�?�{�$H��9_��m����@��ZW��q��Fd��N= �l�=��ZWj�?/mzg�,��G�6���@���h_U�~^���Y�~V�/�9�"xԙ�@�����נz��_U�{�]Ɯ0r6��1���{k��g*��}��_w_w9W���� �o����+Кyxwa�W;�0�"7oNI�{rrh�v�h���c1��u��g���dC+w�-s�ۛ`fs�k��=�㫩qvv�^g�C�$[&�&��5�D7`�o�wݯ�Ƶ��j�Z��f��v[��'\j��w;������s!維��;�x�1��MJ��[8-��3N�[hPޒ���ya��ܭ%7%����*ӐB���N��[��6gQ�!�P?�g=�h�Yg��k��u����unM�)�4v����w/7=ۭ�D�$����u�i��ݶ�����}}V���Z��@��M�ъ<J`�Qɠ{�����?/mz׬�:�r�İ�DI���Z��@:�����@�0�a��B���_���z�7u��w��L̬׺��p��mU0���J�X[f�ﯪ�:�V��{k�&,���Ϳ"�6ӽ�z�{p��lI�zӡe�m�h���:��)]�����a������� ��r�?.� =��~]Y|y��7�5�ٽkyʾ����@�<���^�wu����@��]Ɯ0r6�I�nE�~^����@���h]�@�z�'�"I����I"����_U�uv���ՠ{��h�% "�M�_U�uv���ՠm��������8��s\�.;�<�n����ޢ�]Us��vp����Rx	"�:�V���j����_U�uvXA'�RY#�/�{�u�4}}V���Z^��D���(����f�ﯪ���#?fd�!�f4�|a0���&8��l_B���Y�~�ǝ�M���#�0c	\ZW�8u�!���xTQ\t����|�y�{И W�77�g��Kfk� � 7͟�����3D�i4�N8��fy��&�6�Ҟ[�@����|Y �y�#�TD�� ȒC$�J4�$x2J\���=��ଔ��:���)���1.��vOP����&�b`��T���3p�|G��=������1!�f���]��Fa��fh�15����qB�i��=@��x#������= Ch|�<BA�'�$%t�����T��&'�'�3s�O���=��+!fjp&:�%7a��ך���V޻V�u�4��e�1�x�&F��:�V���j����_U�~Y݈ɟ��ꗆ��ԓ��W�ngT=�	7S�p��i�芇-�۳J 7-+�Vb��c�9��-�mn�;���<"ɏ�-�������Y������bff;���A	�'P �$�@�w�uv���ՠr���V�8�4�&aH�_U�y���]����{�1	����\�C �$�8(q3\���]��R&/�{5%�I"����h^�@���h��@�ܸ��&I��)۷3�1z^e���Y��ׄ����Wdb��ubp$M��$M	ŠUmz���@�ڴ޻V�qwU0P��%���=��Z���?z�ZW��?.�e�1�x�&F��-}V���j�*�^�ﯪ�?{n�rx9��7���j�*�^�ﯪ�-}V��ޭ<~�c�I$�@��z���@����U��s�	�B�U&R��ow�����1��,��Nvٞ:�s8���D�6 nyrv��ve�aI^.^ĚxxGC�h�}�$�bh�r��g���	�z�hH�9�$���n�Ѻx��inC�����q�[��e�6Lv��^I�&�r�mt�����%�ƍ�Y*�w]�]m�c�	��F]�|nd�U�F��lI���m���秗���t$v̫Z�dՖ}ls.�
wO{�����;|n��	��Wm�s�$�n��çoN�v��s�M!j�&q� ��v �ۉ�{m�T�@�׿+2�������Y�Vr��N%�D��$Z�ՠ~�ڴ
��@���h�G\���=�%����v�U��3*��1�{Y��ݭ�`[�˒&�2H��@���}}V�k�h�v���`��L�@���h�V���j�*��۔�l"b��1�<Q�r$�Y<��0<���p�adX�]m�v�(����1c^V�.�F��-v���ՠUmz���@��w����cqh�v����m��/TJ/�^g��\��u�h�V����LfLo�I��3*��+����Vܬ�`}�ȴ0�F� �#�@���h�V��ՠ�4Z�Iİ"< I��Y���+1Xfc�9��Vs!���"��Z�a���2%�L��}�9�e䲈\gI�u�].?�}�"����+ ��v9Y��̬�`fu�ya�x䉡8��f�ﯪ�-}V���j�./z���x6�Y0R=��u�s�w����@ 	>Hh?� �T4���y�������W�v��ۘ�d��@��Z�]�@��z���@��w����i'�Z�]�@��z���@��Z���-q�j:�Z�E�ɷ`l&�،.�<����}8�z�c��:��v��Z�W��=��Z���?z�Z��5G�1 �#�@���h�V���j�*���V�8�'�$Z�ՠ~�ڴ
��@���h��H�����(��~�|�
��@��}��mD��w��s�w߶f����rD�'�[l�=�ڴ]�@��j�?������#0X7�#�Y����g'n� Wd�5�Ι9�H�a2vԓ֕��C����k�h��Zm�@?Z*�m�n$�&F��-v��]�@-�h��Z��F��n6�I�7��ՠ��}��%���h|��@��%��2"$�Š����V�k�}v���MC�Q�L@)�h��Z���=�ڴ޳@3��ffy�g��m'bCɑ���e���<em	�wT�������f���u�;.Z9y�t	������]�ek'7������Np۷`�ygِƮ�]�k"�㝅��X]��tѰ��]���6{��ǇF�U>-�-\v����$z�ׂWlf� �TIuTL����c�� ����99�Ej(�H��<�:.qt��ĶY�F�+�s8�jQ�Uz*�D��Ҵf{a���T[P\�]KŐ&�0V��i�)�Il�f���0vMu�tj��߿����=�ڴ޳@��j�9UZ�#ɽ��I�;��- ���=�ڴ_U�[�˒&�c����z����g�ffa-��V{[���w���<�d��=�ڴ_U�{�h���uۘ�CD��@�ڴ}v� �٠{�h�j��М箺��ݫZ�9u<�M�̜�1�5��z��v�&���-{,�9c�9Y��33��Vb؏�n����Uu���f$��<�U_9T�U�i�	`	 ahrFpc00R��d�Ed&pq����8�Zr�ߞ�������hެ�xB& �94���]�@�}V�[l�-j�'ƒ�02d�=�j�;�U����mz*��H��Of�J)$_��ߖ�[l�?+k�-v����zg�y�b�LO!1��]u��vNrGG`��V�)q7\.5�vj9Z����l������h����V���� ��S�d�cŐ�@���@�ڴ��h���uۘ�CD���k�hϪ��y��g�
*�O �/߼�|������W���7'�q��N1����h����j�?,�tBdhq���m��mz�ՠw>�@?e�Ӎ�:����gW��k�Aƈd���d�,A��Ӳ�.�v��Q1��-6��@���@�ڴ��h��֭q,i) 2d�=�j��y癉���wu�,̫�id7B����J)$_����@-�h�Z�]�@����䉹��BcN-��<�ľ��`qf�X��V3�&b*"'�v<�1K�|����x(G�1��
I�~]k�-}V��>�@-�4���p#��k�{����5�v:�(X�5�� 	l�dG�X�]l͘܍̈-?m�+��v���3;��3�,ݫ�����R6ؓ�r-�}V��}��h���@��Z�ܒ�1	�&�I#�@-�4˭z���=��h��Cj1 �Qɠ�٠Z���}V�[�h_;�q,i) 2BSvew�{3ܼ��ͦ|�_*�QQ_��QQ_�ETTW�aTTWQQ_�UEE�*����*���Ȉ�*���""+�aTTW��TTW�����TTWQQ_QQ_�
����EE�U���*+��TTW�EQQ_�UEE~UEE��
�2�Ʌ��n�����9�>�L��ր          ��>�� @ ��+cC�T�* �� *�    Q@$B�(��  �EPU@(P�*��EPB�R       �@  U� S�'.�&�N��q^�� �гo3W3�ON��ﳡp ��;��<7]�۷����y�� Lw ��  3`  1�����p�燣��C�}c�ݯO|��{� �}B�   @ }��s������S��G�o O��
�� ;� R��P%��= p ���  �bhU%  � ��3��'@.��J���% @�f(( 
 �t P   
b2�= bh�J�  �׮� w|�\�]���y����N�_x>�>>S'��j���w�����}w�{��z�m{��l.��֯���_}{S����{n3�ڹ:�o<\.qڮ���    A� ��K��L�ug'\NI���Ϡ�}�w��o���>�ۏ@�%����w[� c��}<�ɹ�� �}��C�_lw����GU`����r�ri��f ��U @ (*��p xt���z{���^M/���{��O>C�J�ۯ#�w|�`׻���|+�{!� �,Wg.#� �}|_{�����>�=S�} }>�=���>�ǰ\ �AOMJ�40��!O
���  <z�U!�  تT�)*  U?�	OOU)U4��""CRRD@G�|	������������|;��G�����AQ^���AQ\EAS��AQ_�*����
��QD?�����_����<4˻�|���"'��|��Nf��}��yV�Ț�|ҁχe�6���㹬��]�zg3���)))�s����I�^i��<�9�!6�T��(�0�l64�r�2�q���DJg�MV�o3>��VI�T�7�`���4�C���n���<�-�)�~�+���
2O�MV�uw�M�>���=>��� �f ���!q!�D���
B�F����`$H1�OJ�LM�#����2��M�!p�f���T�q%���ʒ�x�d���k�����XS-Y%Ip!L�C# ��\20bA�t9�:q1�5`�H�bD#�
d��!�CbT�S4P�&$��XЙ�	Т��`%
at���5�o5�@���\"�_1x�ͼ*����Ѕ�y���!��}3ۤ!.%[�	LՈS0�F0�d!q�X,�2�A�	%	X� F,!`RD�4 �bT�z��,4�m��}��#<�"�ȱ$B,1��X(P�676i
�¸��0��P�"��H�D�̅���34���=�T�%����%�!q�SX�X,)R����.BK���,R64!N˸�6{�5�HV�!F$0%́%c�<$	|�#m|��R���\4a��J�S\!,IY3���!r˗���9�a/��.k
�k�RVai��8���ϗ�#�v��11��}�0�!�� 0`�� �L2S#$�Cn�0-��1��\	�as}&����4�Ä�VQ�Nl��O�&B�W�<�i}e�<З��F����e<��vP������rzz�2M𓁙�3�=ԅ�O��`iN(Y�n5��t%�\�.�C���h���)��1�u��l��`@"��2�2�B�R���KLcP0(@!
Q��si-���e�nzH�a���H��F��J!$�E��H!j�E�@"��!�""@� �����!��4�щL#LH�0 QH�# �H�0!!��J�L�\4#�6h�D�@5`��l��,C�`��"ȅXR��(p�F1bxG`b@ӏ�
���ݬ��bB#�k �R	1�HՍ\x�b��!!�A7����۪F9H\$�Q��FD�@"D���k>$k�B��p��15�0�,hĮ�L\#�.�i1� ���p$V$F$%0�	dH0�!	p��,$1aVaR`R#Q �����̄%0q��F�0�#	q�Za&XI)%���<���׆����C�
��3M%�)$��Hh¬fB����n��j�h80)`A+Bj`F��ŀ�� �,R� ��"T��T��"�1`J�N���!WT�Tȕ�0H�0���a��J���CHW�q%b8���A���H"PcS\$��5%0�H�10e04vS46X����4J�*E)8P���*�"����(B�)�Ҟ��]�B����+��˼����`\�X� fz���D�}����CS+���]9���'7�#O|��o#1�T��Ӛ��s�B���$*B�6�sv�O3v��0"��$�o�������L0�.P��R�0�%XT�q�@��HP�ńH\1&YYHF�HV�lnI720��H�1�H�&�@���`� Wzk��Ƙ�
$)��	F��5�L8z�bj�bT�Q�0��k\7(@�B�jq&H���+����IOx����A������9�<H�%=З4��p���
�o<��KL��
m���}�yCs|=y�X�dd�$�r$�!��a�F�#@� �!HA� J��F0*F�/\�HHQ�#	'�2#Z>�)Oε���W�p��͡'�>�S_5�G�Q�LW��*Nr�E9�d#�E�~���>�S��_�ec�J��8�5P���p�����P����~�C�C"�e�����]:iů�y����J�(�6Vq�}�m����Q4�_�M ��y�9p��p�f�9$
I2�b�Q�zT�O�Bj�Ц5D�JW�J`��<]�7?5H�hs��WPQ2�*H�����]��T�R�W�d#�%�C��7����e��>>Qt}V� ��%�΢���__��r�C��C���I}�1�0��8�\�=ϾX�qn���
�U4���QW*>��8��B��_G�]d��쯑4� |�,�T�>!'�lc�a ��H��b�1J����Ǎ#@���	�hR(D�1!����m!B5�JBv���8�e4�
��x��aw��(B�<e���Ӂ�B��È�����0Zf�7�卥h\lۛ�����	L�p��HJ+s.����Z
�iCB2��X1�!B�q�\�@�XP�KJo<�&_9�U�H��ʇ	=��}���cM����9��A�$�X�愦e���}�^8��OO%�G�� a�K�w�.:@�9�@��%�F!�b��AŊ1 Q P5����e3^%|<~=H\u8��X%!�*JS�Sˬ. �HQ�"��ۛ�����y���'�B�d��2^C̣����&,������!Ji���D��h��|g�/�`cUyyK��}��!�!J�JP� �X|C9��j�����^>>$k�"0*1���@�C�<�3^'��	j�"�h���cL>/�@�Jc��|S7��F%#n��WՂ��F��
�>=����p#+����c���H��}XZ�Y˞��ﾩC���<�+�Db��B��)5y��i`R@́XՉ �Pq%��|e�|�x��y~0��>|}�af��+� 	��ӄ��:F��)�v$4�!q�| P�B5 ȕ<B1Ӂ�⌦p$|\�x0
�<"�9�����O�B�#	��q�y����w���xB(�����o\�qׇ�b�c��%�:��}��\7�
ĩP����]�H(jB�`Q��8t:��cfo�=�%�z�B�Aw1�X�w��x(iA �!"�З$4`H�`B#SԳ���A`A�� A�y���8��'�S9��
��ƱHhE�ѩ���7�c>=����߳��hH�A"D�c0X�� F$�Ej���#���`BP��2�2k,�z�4&�39Č�������`��D�E0h�&x�H@hfG�(R8�0�ĩ�)�R
��y�����ÆxC�=x���x��8˞���aOr�Ԕ�����V�-�HP��8cb�aʼ/LO����8Xa��/��<�$��}So�w��Þ���9#��͖�)V���BH���+>�C��R�B�p!U�)D�T�`��v�aIp.O!�F�&�@��i�i
#HSXU2$	YZR��F��!)��(��JJeŊQ��ŪĠ*DhA�B���$*0H�)B%��ą`�5cBtBF�	f��.@�fj!D�K�Y���LK<'R�Q��ު#P���t��H֨�����撘i
Ĺ)�a0q�5p������D�P�t�"���}��7�وʿ�)�B�,P�"%"'�Q�B�����(`��B���of́%%e���0�݄ې�"���#B$�D$YBP��?FMB����CS�����C~^�Y�s	(BVY!$�!� ��,!J������!5��z�d����ٟd��j��ח*���[� B�0%&Cy��  	  2��!瀶��	�\<(k��i�n�v�Zu�/�)<�PY�A�����.T�͸�1��A�e�8���%��m��n�h�H��%
�6ݘ�΂y�\ݎm�;������:�}"�6���J�����N���H��7=���]�7^����6��t��]@VvE!�[��`���۳-�/�=����c�%����U�9$��c^E���|�|����G�=��ڨ���n��AS=��K�5i�}r �Z2���q�-�9�]<�m��S� �{a! ^9Y�ӵ˶�:v�7oOP[���6"��hv��r;�P6��M��W��me��k�r�k[��J8sԸې
�a܊�`.ܛH��.�!=��d�]���v䶌�1��I���R�O�lsU���=#�J�/J�]��ݹ�Ī�5�=gk�Q��(ˮ�$�`[vձ��:������Dy��[ǶH"ޤ�����T�  ���rݷj-�9�-����9��0 � Y���LiNKm�����I��  �Amm���������	8l�  ���BM��[`m��i�kh����� m� � 	��F 4�-��"F�8N� � kɚ=.ջ8mphܳ���M� hp�&��n�t�bvM��ٯg�C� ��tۉ��MQŸhn�Z �
ѭ��u�
��ʩhŶ�K�z�D��	ĉ4�:p�-����lV�#  ����Yj��/��J��ڗv� r��U[TH�  �H[f�K.��nA�U[U�KS�H4巎�  	   v�<zn�d����ΥI� ���  �`p�Mۀ�KonE��Wk���z�  6�$�$�[�����ׯ�;m���݀�l[C����5�J	 ���*@[��j�f�A�����0� &����UV�+��Rޠ��l�+`A�����N��U6����jUط�N���	�vͶ-����l-�"�}��� �@+lKk��@  i-�E�-�  �$5�u�.���  �N���@$��m�%�m�i0 8p6� ���l��n�E� �8�H�[FۧM�� �8m�m�}ﾭ�� "t 㭡�Z�רH�m�m[[�`�� �M���  �-l�pm��lm�m  R���K�v�rPM�i��� �$[m� [C[m�m�   �Amo0	 ۶$��CZ�-����)klp�m�m� � p�m��A�j�    H��I �  [A  ��   l�  ��t�-�Imxݳl�  $$H plt����Hm � v� �ݰ�M���lH �-�
Q���;m����v �	6� �� ���u�|�zI6h6�n�-��pm�bN6�Z�5��-��q�-&�n-��     mm�� $m�p�+ʮ1*hZ��jt%��  � m��    �Ӝk�֍� *����; y�X�M���"N �Z�����\���`-��h��U�;o��P  	��8dH h���l�6۝� �C�j� �	6�i	e�f��tۭN�; U�M�^�6��9U�
_l�s���V:�z��ǃf�Y���ʓ��[e���k    H���rQ��� ���n�-�F���g���XP���V���+j�u�6Lj�\��F�*-&۩�kn���{*�0mt�Ov���̡!Vm�&����$X�y��X'v��u��	5�t��� �"EQ����V�w�]�A���6.�jUU��j��bW�: o]m�Mm @,��z��d]-^�]jԬ��!KU�mI{ZH[@9 �f�8�-��` [V��ZM�J n�N�q��Vrc �N�&�p ��i�l8Kz�8�,��6�2%��pN�� m&�K鴄�[�[Rh� p�Qt��8]3���^ty]�'�0-�J��q�N�e�j�Ω�6՗,�
^$sj�@icZ�׭�m�_��I��I>�YdΚͷ8$H֊$p���m� ��i�u�Y�� R��*�UO+UT�:[�pm�n�6꭛m �kĀ��?h|  m�a�p �6�  �m:m�m�klP�� 8 I 8 �  �: ����j��q���kn�u-�m�m�m�@ � � �j�lz]�� lm $t��knm���@qmm�Ӹ���	$��l�Ãi6� $uu��l�m�����  	�=&�l6��X��u��@6�	7E [� �� u�o����;kz�4�F۴�H��'PH �K�\�ר�d��*ڶ� ����Mf��MT�t	�4��Um��	Xٶ �9$�-��[U�6��D ���y:��,�
�⪔��] s�ڕm�cR;���Cb���U�e�0��Ӷ`u]Ö��� km��{���8��e\�t�4Idm�bezT�U�ڥ%��N�n��� �6ݒ��Uk�e[iV�l�  ��o�� ��SI�]�4�L̀��[NQ4�8  �     I���  �  [@�`$ p$ ��-�Jۻl�}w�]�\����!�3k�hA��d^�i6H\�*�mҹi�Z:���mݶ$�\�on���i5��4� �kh  ���8  h�H   [@   $ ��(�$l�@���j�&�[u
�-f�' [R��jy"ۖ�iVRy��ە2���K 'G�K�H�ZZ�`���5V1J�E@oSm�mm�m���A���H   �   l�  �lH   �6�Kh$�tےl��Ԑ-��.�*�m�Khs 9۴�l:�mz�Z��{�z����Ls-j�v�#{Y�פ�:ŵ��@ H��Kq���ٶp���[gNm���������5W*�K�5t�m!��[m��u^ڕ���nl�t!mZ� ������ms�ܚt� d`m�%�V��%�dm��v�h��� (O+��C d��]+��u�		�{\���t�	0@���1�+��b@�6*�ttWn���i:^u�V�i�D�*��j�lLǬ�Jt�qU��&�e�%+m&�   ��j�Z��ɱTs�j�SK���tR�m$.�V
�+ɮL�� T����m�ש�$�������&m���N�� m-�z@m� H�d�*�m��^�#���s�j]�j�ۗ��P�p��Á� ����m���m��$m����JZlR�@��u� 6� ���@A��T�+F��* z�6������d�   N��  H�l�eZ�vx�`*7SN�����m$�� ���HP*��V�:*;L�`H[@[]!m�m-��M&-��  I�u�P���;&۶A25)����� 6��m�2�N��2�`��-��[@�  
�UT,,���< *�T  $l�fl�nI;rʵ@v׶U��'l$-����&�a�	�k  h�m*�	:�6 8In��-�M�6����$�sU�6ey��@��v�q��	-��� l��6���	$R����cRƣm��mm�-�D�V{m�)k$r;r\�n� b)m�*��|�V�*�V�N��r]V���᪍;���Ao\��$j� k4�]�oO+�*ʜ5mԪ*�r� ��B�`.�[`,7 8l�Y06텴�  8]Wpm�0]$�-�@�m&��I��i�/]3$-������     �  8  �|Hm�[[l��n��� H  �H d��(���� $Hp6�$ $��nZf� ٶ[d�$ m��[A��  �        I[U���� � �6�m�ۧ��"�m�h ���ݶ �A� ��[zJ[Ŷ5�` ���dݶζ�m��r��� H   	   �   l�������u��I-�����-�e  	   �    � Գ���w���@ [[l �8 � 6�  	 �m�ӿ���@�ֲN�6�v]�m����#����TQD  ��04��A�"��
�ZoVg�� @�8����=���>PR ����(��>t�C�#ቪ¸�����1U�OS@4���W��+�~NZ�i��tG����^z�Ə�A&����E`�Pӟ"	���Tp)�����Q}�MX �S�:�<CT�!�@�U`)�s�(>���AA�	����H�Dp р$b&	ê�ਇ���ZT����P8*@#�G: �@y�
�F����A����uU} pP0>`	�1 ��+�Q9�Ǣ)�J�=z�'�2��b�'~U_C� �EMN���pSׯ��$��ł���`A�IЖ��[e���2��ьX�R����.����P׀-Q��s�T���M qUC�꠨�� ��  E ��� ��̶�ƍk%���6��nl
C�Y�֐��� ,2OF;>���]n�0�8�!��lˬ�������3�'#n�����c��La׎wSmlt�s�˷�r-��S��:�ݠ�_-�gl�j�S���vg5�[Z���fEv����,�`N�n�醭��s�e�X���vؠ �<�T���	�v��gN��ŝ7��=��95��F��s�N����۷=�[��W<9��w����p�k��Vɮ��;3��m�K�Y���:���㤗jl��B�Ԣ�]UVX�r�ᡎ{Mar��I��UP�RI�2[l�	̏9W�ҭ$*�@Ptɪ9,�5$l��K�	�֤�ekv�cN]����:2���7�l��ᶩC�ٞ���Q��*g�k�=��F3գ���=ql4]G�KeW���"�;v�xb�,.θ�3�h��Wcl,t�u������	W��9ݒ]�1��L���4�T�S������,)<�k]m.����9�`ە۞z�9U^3�Bؗl��^v��O]���kv�.;b(��E�wE��Ů��P�|\7�S�[D;��o&�7�v�N��v@�iV����P�4ӕWSl6"�����)l�k6+4�U�2nL����e��fiT�g������ܲ�JC�������	x�S��p�:$��\���Л%�v�6�jx�CqVۋf����v��t���WCD���7<�'a�GL�&n;K؍�`�z��0O�cW&�"���LX8��"�b\�e�vSb{�T��=eUW1�M�!n���U� fyKd9���P��׶�WnL��2tul�v����3�Ov�a��l�(�L��<���j��[�:�T:nJ��FIKwN��D%�4�WKJ�z`UUi{<@�OX�}�ʳ]m�r�]n  $v�C�n�U�Quہx����3�]��ˤɷ0W��	E0_��������DL}�F��" {ݞi��a0˻&M�32��-pӥ.6�0콞{K�%q���$���۵X��ݞ�v�b+�S Ԥ�MU�'�\=p����b�j�B;��s��[؛�=���]�6$+�XCc`z��v����shweݫZ�dIu�a��G>��yz�qd1��6���F��=�;��7�v��O]ֺ�"�<U�tk�:�����h ���Pj�#��;d�r�a�]���<��<��3�태�y��L9�� mC�s0�׹�@]��d���y/{�0/���/����K�B&f(�j�;���w[4]k�>�z*�cb�QD��Zu���f�˭zs�h{=���S"Q8hu�@�ֽ�ڴ�)�{�J���$�̑�#rh�נw;V��e4�٠U�(�I��d2G��5���în��$kFìj��v����M&�H�FF7��;��@�v� �h�נ\W�&��12L��O}����)*� >�"�D=��
�����I=��zs�hò�vm�x��@.�f��{�G&�#������g���!��RM�Z��j�;��@;����쩩0�M@rG�w;V���Z�l�9u�@�yr�e�W5�V\��ù���'Nj$�U�Q��[�f%��E�C8x�DX��j��f�˭zs�h�ѱ;�<P���Š���Z���t�n���l����Hp�Tԑ
�j�G;ٰ3'v,��4�Kk1H��h��4{�V�[�F��q��ՠwYM �h�נ\Wɶ���L$�@�l�9u�@�v� ��B�H9#�g]V2j�
wmu9aA9�(0����\���.�A[��9�ɉ��Q�����w[4]k�;��@�G���!�����v+���fdw:3�� ��h�������H��j�.�t��fgt��(�d�q08NE#qh�ՠ���Z�7�P?�: �/��@U�TmW:yc�n5C���Kq.�;��.���ՠw;V�u^x�y	ո�`kv(��'Cr��[�2]0(Z��t湝�Bh �7S����r�^���Zs�hu�@���i5��j1�7���Zs�hu�@�ֽ�I�P$HE��h�ՠ���Z��j��eN6B"r���e�w�����wF���Zs�h�²@r���34�݊�������΀.�j��Hi�&ąQ�l��*��������5��Jv�u��q��1��ٺ�$R���ԁ�����u��hu���ؚ�&VFH�[�;[�b�s��n͍`�շ���&Y#�=�Tkq����[n�lK�B��>%�9�W���k]v����՝��jKa콨|���:�U���u�1pl��L����8�hh��
�s�Iͷ)�Г<X���ƅ�Bw=��m:����{޻�����dh���e�j�f{B�]L8��4N1���q"��r��x�N��4�9#�y����)����Z�q�q��QQ8��)���l3;��ǝ�@]��2�sƦ�)��i�@;��.���ՠwYM��T������7&�˭zs�h�S@;����I��ɍ�JǠw;V��e4����v(��5q(Bs3$9�M��g&�f�q��޸e];�-k�s�p����l���M�Rm�	(�/���Oƀw[4w��{�����(���r��TXf�_1	����6���Ē�M���$�/�
����O{f֖�G����o#iI4]k�;��@�l��/aY&E&�)�����y���Ξ(�vhw��q誑��B(�(�Zu��9�wO�c��.�u����ʘ:xFCk�����p��V�f���+qm�$Y#i���"�'1��a D�p��f�˭zs�h�S@�xU,opCT�R�U3U`df��[i��r{ذ9�������U���i�����̝ذ36��^���M�I����ֽ�I�P$H4��H��)����Z��j�
��1��L���4�٠r�^���Zu��*�iq��F�N,�#�L�Z�hb����p�7���o2%��n��3���RM�Z��j�;���w[4��VI���n�=�ڨ��(�vhw����6n,�'�DD��=������Z��j�=ǔi;�<X�DD�p��ڰ23vl�݋	��B�i6��8= @������I�ݗ���C"Id�jb&hw�{�ٓ��<�~Z.���Pv<r(�D�ibk:.՚��l��#
ݐ��IU7rbi��sn�-��S#O$Ơ�zs�h�ՠr�^�˭z�|�n�H4��H���u�^^^lǝ�@c��.�u�ˍܘ��	�H�]k�9u�@�v��ڴ�aq�̉�cR=�Z��j�;�����Z���+$�$�$zs�h��:����t�݊�מ�m2�Ѱs��ώ:ǧ�������o�N�Ls�g���r������l#�9�[�N�x�{I����kܦ�L$�7�{&�ݶh��9,�e�Q�0�wI�mĐ�'b6��q۳ӎƻ\�n�p��k�>�y�[h�g��vl�)��͡��u�ۉq�z�vq�)����Ȥ<i�,�����-����v��&trirO�|G��\ͦ��l.ܻ�z2��
��ڢxzPq��׳TgW/n�1@!"��'�5�8���~4�j�9u�@�v��yF���ŎdDJ'�ڴ]k�;��@��X��X�dɑF�Z.���ՠwYM�ڴ{�V�[����('���Zu��;��Cؼ�u�T6����-��h�$��Y���wEw���fF�!�5+��ƽZ^Z���*��i��l�ƐK�ԁ�.�6���x.��[��q��w��n��^��3:x���ST4�%T��E����z�m���P�ձ�ƛI���b��r��3&ՠ\^²L!"M�RG�w;V��e4�j�9u�@���o$k"qh�S@�v��Z��j�>�yF��O9�(�4�j�-��Pq����(I.Z���S���Q��6KA�A��f�Q�sAqW9y��ף1T��r���]1��O���@�v���h�ՠ{�J�ǹ-�P�q1@]���fgOdw-�Z���u@�xI������;�f�P!�9���$5�tT�(��!���H�I!4S�=Bҩ	+��Ԍb�r���)�ST�8`���?P�=��f0��� ��*1h�K���A�F�D�(
��6�܇��p撈�j�?xt�RR�ZZJV22��e������U����z�ڀ0㇨�D@4 �Q��)�*�~�]�w: е�#T�p9�L�&J�㜮�,G;ٰ3'v,<���}���*/��D��'��h�נ~�fOs�Ξ(��t���vP4�#-�����lU�#�v۳l\#)kk�Sp>+f�sP����Ÿk$�&�$|�ދ3kK2wc���������p��P�ŠwYM�ڴ]k�.�u��/�r�0�~�2K%�q&�k���˭zs�h�S@���mDRmB�*T���(;�#;��̎�@fmiak�7�����ZM)�������!��'��('���ZgYM��h����漞Cr\�s��b3�ɐ�lIÒ9�����ĝV�K�^�������Oj������~���h�נw;V�P�w&D�ڄ��4�)�r�^���Zu��/<^ʉ"�O$	!�r�^���Zu��;���^����s�9��y���Ξ(��(]k�=Ǣ�D��	DQ8��)�wYM�Z��j�����H��?+/�ݞ-�5��
N��}v�q��+�`g�üg�x�ms�u���0]Z<)���[���;n�a���$ych�z�'��ɇ($j�!�L�7��Oi���ƀ�86n��󽎖s�nɎ-ґ���	rb����=m�]��p���/a۝�j���I���c�]��v��.�=���t������[��&�sf"���ϛy'77L��͘.����o)vx����/�s�������[�땺DZ�&2bQ�����p�-��r�^���Zu��=�%R��ǒȣn.���ՠwYM��(�oa��p�8�9LP��'���� � � � ���~�|�����~���� � � � ��~��|�����>�ff~�[2�f�7v�A�666?}��� �`�`�`��߹�pA�666?g߿g �`�`�`��������lllo�>?d�ƛrne٥���� � � � ���~�|���������� � � � ����x ����ӂ�A�A�AFfu
-��N&G!m���G�ܷ6��n]֛���V��%�q���M�4ś6\7d���� � � � ��~��|�����o�ׂ�A�A�A�A����8 �
A`��A�A�A���8 ���I��p�f�4���>A�������ȏ@_j!�A� � �������lll{������lll~Ͽ~�>@S���A� � ���˟۹��n�̳n���� � � � �����|�����~���� � � � ��~��|�����o�ׂ�A�A�A�A��o2����&�nfl���lll~��?N>A����������lll~�~�|�����~���� � � � ������	Lٶn˷3g �`�`�`��}��pA�666?}��^>A����s����lll~��?N>A����D��߻��<�n�	�Ӳ���7W7�"��7ag�9kW,Z�L軝s��ss�� � � � ����x ����ӂ�A�A�A�A����8 ���߳��A�A�A�A�������d��5�&��`�`�`�`���s�pA�666?}��� �`�`�`��}��pA�666?}��^>A����I����i�&�]�\ݜ|�����~���� � � � ��~��|��8�>�B�A�<O¿(�}A� ��|�x ���?N>A�����d��34ۆ䛻8 ���߳��A�A�A�A�����A�666?}��� �`�`�`��߹�pA�6667���~�w	�vK�L�����lll~�~�|����1W����pA�666=��?� �`�`�`��}��pA���G�����lvY�u\e��,|�]U�,栋�S��w�1,YkuS�jU�M����h�S@�ֽ�ڴ��Q��ɓ$&�4�)�r�^���Zu��=�%R����p�9u�@�v���h�S@���i�r$�b�#�;��@��������kIڧ˻ٰ5G6	�Աby�a$Z�e4�)�r�^���Z��^71�&1̑'��ո�S��em�[���L��:��F^�`����26�L���e4]k�;��@X{=Y!��Hh�נw;V��e4�)�^�ڋ���H��j�;����e4]k�=ǢvD��"�ƈ�ZvΔ�Δ�͊^y����\�o�ɓ$&�4�)�r�W�w=�@}{:P��x���d�����m�fbֆc��w#����2\��'�-���eb���ۑ�flE��������X�i�rq۴v�W)��̦�wOfvɓlѻI������Gk%i�!6��s�<��=�Sq�k��5��@�%���q�84OQ��i;Q'e2C�B��T<hx���Bڣ=�qဝK��\�>���� �BbY�2��L�囶�L����5y�=�쑫q����D���Xe��S�8d�$t�%����HN�ibջWm�G��p/_�@�v�u��=�%[x�"x���zs�hu��;���˽^�quCn�ŉ�FE��hu��;���˽^���Z�Ŭ�R��.�D̔���:��<�=�ڴ��ha������Hh�נw;V��e4�)�\����Ƥ��2I��!!��)N���)�N51�n��.�LN-,�,��I���Zu��;���˭z��VH�x�Q���@�$� Ȱ��b@~�����w��^���ՠ{ǔi:��@���(��(w�w�̎�@^t�@g�*�kq�s	�	��r�W�w;V��YM��h�
���D��)��H��j�>�)�wYM�z���.nD���䘖�7 Lf8a�.�s �/o\��nmζ�m��n&�&V���đhu��;���˽^���Za�S�R�!�D̔�Ε�y&�y�dw:��Ҁ֌�TL�DK��RTX�6d�ŉ$�&�g��jK�S9�:P�:P��{�mǃd�$zs�h�S@.����X�m�D����Zu��;���˭zs�hy���#�xFe�z�:�ۅ�b�J�d��i�XiK˂l�HAs����ڶЭ�����n�b�����_0����5�8�J!D�T���I@[�خ�fdw:��wYM����W��7#x�H�छ���,�kK<�K�L���X�M�޲"54Ӆ)��3.����:��9��K#9�a���v�hbbBd�  � `?� MW���5����`rW�z�S2��U"��3kK�?6����v}�>ͭ,?;��6Zgm,�BLl��n�1U�5{j�x^oY�j�] �~>�w_�'݄�+B�	�>oEw����t��%�Ξ(�z>�m7	�R���w���{�l�����‷{�\��M�r��8�bq�dn-��?u�����&��tP���W��q�8S(�\�IA�������ǝ�@]����/y�uq@f�}!҈S(�29q4X͛�M4�oތ���`fml�~��ꑄ�� R�u	�aH�%%c), ��F ��y����BH�b�BJZYZ��Vba�آEH����#b��$!F1�u`�0�H,!�d��Z"��h�S��%HX0XQ-��*@�!�,�0H#+�$!��X+�Ą�`f"HX�1\0�
F!!&,Qi �1�1 �@�2��P�"� %"� ��A��E���!� !e@�� D#!��e��H�@�Y�<8���>A/}̶�32ͦl�>����齲5+K���ͳ������;���`�ǰb�%I-�86�C]ێX��춇Jj�9#��zzxݢ���Iz�`�LE�ۦ��qӲ��&x^����6U;",<E�pGne��ъ��S�E{X���6[r�z�gK�=����y6�ۘc��+<m7#��nɪϦ��x�:i��:�|��NWWJ#�x�r�ڱ^m�sw8W����1.�lk	-n6�۵8���빕⍜&���)���.�:�]%-B���y취N��::Dݻ��aV�V�9��r����U�p���a�;;$�zgM�ҥpƥT����k.[�wge��nl^c��.Ċڅ���h'u�ܵڭ;q�n�c�lD�՗���ŃQ�N78q��9�ї�k���K�ݷF[���.�.6�u����;m��z�r�M����_5�͋�
l͑X�)*�jז��8yщ�u�i�/�Gl�:�18]WJ�riJ�Bɹ<�x8@j�8�Uxv�U��ҬcP�N%�=w&��kn��m�hܷ"�ls���&v���As�C�[�z˓�l�C8Ӭ#���n;	���nxR�X1Ʋ�z����U���f�F�e0ru!���m@c$�%�l�&��Ο1�-���	��`$ ᪥Z��f3���P��l�Aͱ�����]4�u\* 7����x9ퟟc�keٸ ��=�Ӱ.�2����y9�u�aS.���ۮ�t\<V�T���\�����[������*v�rI@�#���d 4t�D�J ������f�OW"��F0i��L.�yE�Yu�0i��۵�b<�Q����V Ȳ��� �F�v4���<5l�ڱ���Ӟ����W|��ۜf�r�E"me���j�z������Ɗ����I>��-����clm<��pv�R�N�m�m� �L�D�I�fݗM�k2�މe� �Ͷ�UMgL����va��ʌ�����l��gs������%O-�E�*��? A~ xy��3�7wL��ܛ�z�m�jY��K�k��v:��23��jCv�I�N�z]�+�����H�70-����</<J���ݺ����t뎛u�ő76�'���n���S6�d��E�)���O,Y�jX3�rP�V��ջjh��/c�����Im�1ǳ��w�hYV�)��Õ�V�z�GY���]�Xp"��{V�������{���{������?9X��$8i�g\�-�%��t'V�_mn��������wz���܍�� ����������YM��r^I|�oE��1�r��
T�3.���t�^�I�3��oEw���K͜�W'�,q	�
e2P�<X͛?M���������X�8j���r�L̔�O#7��̎�@}{:Pr����;���s0�A*&&(��ty+ή>3�����m������F�Y��e����^:�yt��V����M���t�:��>�w�_��Җ*h�S5���,ͭ,�ݟ5����h��#I���I���Šw]������Q�3f�{��ϳ��2wb��O�!ޝ�LL�L���TD�Ĕ���(��tw�̎�@ft�@f�ÅJbI.YDLPs̞�@fGs�.�t�瑛�@ry�q�6B��Lˠ>��t,ή>oEw�������x�ZH�촃y#��T��v��6�v�q��t9�b������Q���I��|��~4]���j�>�j�
�q�9�<�$��˽^���s��Ł���,ͭ/ɷ���s�;��X��d�z���Z��Z\��M���[m�V�t�9�́����*�&h�S5^m9�߽�Łn�b��/z2{���t�n:�e!-�D��0�7���c�;#��\n��,�y1��`ɐm�ƞ(E z�����4Eқ��N7�]b�l��_}��s'VҦG"O�ǝ�@]��.�u�_0�~��үɧ���p�!����k��l̎�@ft�@[�خ�g'���&�B��Lˠ3#��{:Q�7�7��̎�@kZ�̱�'*%�q2�<��������`fN�XV��M5�Jm�^�{Ͻ�����f�D�������l�K۷�F͟z,�)�^�c�B�I9&�<y?�PN�u��`'�Y�Jl�L]��-�3�����4Lq�����hs�h�S�|�����/���5"M�dn-�v��6ך�7}^,���̝ؿ��i��{�;��/�Wj�	b�}���bX�}���Ȗ%�b}�wr'"X�a�2'�o�׉�Kİ~�߮�"X�%�~>�w.e��4�n˗3gȖ%��D����ND�,K�����%�bX>�{u9İ?3"}��?N'�,K���~�r��s�n�vf�D�Kı=�{���%�bX~`}��]O"X�%��߹�q<�bX�'��w*r%�bX�:�t�;2fm̹.���v���j���z�ۢr�Ѯ���'v���.ᓦ�ѠҮ[��]�:.��F���v�V���;s)���vf�:m8�dN[Qt��0�z��6쥷8�Ƈc�ܔ�����qna7C�0t�����Q�Ȑ͆��s���ג�h�䎝�s��77.g�w��1�th}�(����(D��zF�=�W���耉{<V��7v1�f��[R��Q�2p��3�VW6m2ܜѰ�rf�m&��S�%�`�;��r%�bX���vq<�bX�'��w(����*��j�kދk����W�UU��K��3v�r%�bX���vq<��ș��w?eND�,K�����%�bX>�{u9�ʙĿ��vJ�D�*�U!UE���@�l�~ʜ�bX�'��{x�D����~�߮�"X�%��߹�q<�bX�%���{�i[�-�f��ND�,��������<�bX������Kı=����yİ?	2'w��*r%�bX��w���Ɇ]�s6Ss6�<�bX�	���5cP5P/6��p�}�-�D�,K�~��Ȗ%�b{�������oq����m�i�j[u=C8^R��+q��\_�s��o�����7m��rֵs����r�I3rD�H�
����k�j�kw���O"X�%��}�ʜ�bX�'��{x�{"X������Kı/N�~˙w0�&�������%�bX�g�ܩ�C����u�ND�7����<�bX�s���"X�%���gȟ���;��,O���r�Æ��ݒ��ܩȖ%�bw���x�D�,K��n�"X�UXdL��߹�q<�bX�'s��*r%�bX�3��.t�\�r�����%�g�U��~�߮�"X�%��߹�q<�bX�'��w*r%�`)�݉����x�D�,K����]٦\�r��۩Ȗ%�b{�y���%�bX�g�ܩȖ%�b{�����Kİ}���r%�bX�}�/|��˛&�6�v�7g+�+�͜OA&����h�����:�L���?{���}�����&f�pܓwg��Kı;���S�,K����oȖ%�`�������"dK�����8�D�,K�K�f�V��f���S�,K����o�~Q�DȖ�����Kı>��?N'�,K��>��ND�&TȖ'�����7���l��m�yı,���Ȗ%�b{�y���%�� �P�����&D�w?eND�,K���׉�Kı>>�rfw&a�M�6��۩Ȗ%���y�q<�bX�'s��*r%�bX�����yİ?�S����MND�,x����w��K��"��w�{��2X�g�ܩȖ%�b{�����Kİ}��jr%�bX���vq<�bX���m��su��&�5�����Ju��TKU��(��&�9"�:!]t�ݷd�37*r%�bX�����yıP'�ZSV5P5Y�zZ]FH�D�;���S�,K��g߬�?˒�Ct��x�D�,K��f�!�9"X�}���Ȗ%�bw;���"X�%����'�?�?��ؖ'����TR*�MQMX�@�n��[_D�,K��;�9ı,O}���<�bX����ND�,K�O���sd��n�n��yĳ�"w{���"X�%������yı,{����bXQM���u�O�<�������%�bX�����m�w6�iww*r%�bX�����yı,{����bX�'����O"X�%��}�ʜ�bX�'��x~�sv�3ss32�a�]�Dynf-Yk5$��ėm�P�lD����~���r�R�K������`����"X�%���gȖ%�b}�gr��DȖ%������yĻ�ow�~��r�tD^ﷸ����ͽ-����#R5[;=�jƬK������<�bX����ND�_��M�b_����-˷�lݗ.f�'�,K�����*r%�bX�����y���"d���Ȗ%�bfuq^_L�g�<�V�qRs
%!vfnT�K��"}�?~�O"X�%��~�u9ı,O}�;8�D�,K��;�9ı,N��l�:S.Iu�&n�'�,K��;۩Ȗ%�a����?N'�,K��w?eND�,K�w��O"X�%����}�$�h؞�@��ɆF�^33�\����Ȝ��C�v�'e���L��:8��GHh�:m[��Gl(��<�J�J�{Y֖ة�u����nT��	ֶ��x-+����9+�N�6�9��u�.�}���2�/d^Y��[S3����ȃ������w5�8��v:�&X�[^��963��u�re�Db��p���Sbh�v��z����[���}����⥕��L�J���&���Z�NJЅz$�>bV"�$k���w��=�t3
�U�@�@�{����%�bX�g�ܩȖ%�b{�������Ȗ%��~�u9ı,O�N���p�3M�nI����Kı>ϳ�S����,O��߯�}��,K���59ı,O���Ӊ�Kı=�}e��.�ۙ�l���9ı,O}���<�bX����ND��Q�Dȟ}���Ȗ%�bw;���"X�%����[{��͛73f����KSlJD���MX�@�s�����X�%��}�ʜ�bX��	v'{����yı,O��7-���nݶnf�ND�,K�{��'�,K��{���SȖ%�b}���x�D�,K��n�"X�%���.���nY'j��0-�T�veŦ)m�OTmd�Pz=��+t�]�-#�9�5a��w���K��w?eND�,K��{�O"X�%��w�C��DȖ%��߹�q<�bX�'�fa�&a�m�ݙ��9ı,K���<��
$��NR�U�by��y��r%�bX��w��Ȗ%�b}�gr�"~2�D�?��K��m�]w2]��yı,���Ȗ%�b{�y���%��� SblO��?��"X�%�{����yı,N�}�37d�.�]�]ݺ��bX�'����O"X�%��}�ʜ�bX�%���x�D�,�,�<��)������5od�T�j��TMݜO"X�%��}�ʜ�bX���5߾��x�D�,K���S�,J5Y�z[_@�@�9��.&j��v�P�r���f�I!5\�\��I�'vy���i��������Z��+�j�����ı/�~��O"X�%��w�S�,K�������ȩ~��,K���a������ۈ��D�4*��,���yı,s����bX�'����O"X�%��}�ʜ�bX�%���x�D�W�7bX��Kw-���nݶnf�ND�,K�����yı,O���T�K�t�o���B1��R$@!�	!0��|ŉ�"���"$B"�"?
� �i\M@�EA!b�*D�H�$�`@�	F��r�_H����)��A�HA"@IL��f��0��.��u��0���O$g�� ��adX�gތ�� � �����I��#�{�H#!A"2�A��'����_T�(bu0]A_����	����MU^��ê�h�~�}���yı,O���jƠj�j8��f$�$�*
�r�l�yĳ�"w{���"X�%�~����yı,s����bX�'����O"X�%��N��̜.a���.��ʜ�bX�%���x�D�,K�0>�߮��,K�����8�D�,K��;�9ı,O~zw�p���΀��-ԋ�����.�l9�#��EO[<6������}�����C�wK����Kİ~�߮�"X�%���gȖ%�b}�gr���_blK�F�}V��P5P5�=<�&�&	�����S�,K�����Kı>ϳ�S�,Kľ��w��Kİ}���r'�ʙ������737e�t��8�D�,K����9ı(�fsj��j䟛�CT'��E5cP%�b}��N'�,K���ovit���*������JF���յ��İ~�߮�"X�%���gȖ%��Y2'��w*r%�bX��}�{�n˛��,���yı,s����bX�'����O"X�%��}�ʜ�bX�%�߻�O"X�%��M"~cMۧ��F�ϮhDۉ�c��KIb�ա15gd�j�Lv�p�����S�,K�����Kı>ϳ�S�,Kľ��w��Kİ}���ﷸ��{��?�����sgV�X�Ӊ�Kı/�gv�"X�%�}���Ȗ%�`�����Kı<����yı,N�v�fd�sͻfa���9ı,O}��O"X�%��w�S�,K�����Kı/�gv�"X�%�����L6�)�M�8�D�,�H���59ı,O~��Ӊ�Kı/�gv�"X�%�}���Ȗ%�bw$���ܒٺe�K��S�,K�����Kı/�gv�"X�%�}���Ȗ%�`�����Kı8+� @����/~D&t�� Ź[���\Gn{9(6���x�qf��g@�����7u�ų=��۳��q`��l���Rc�������k�3�������Mq������Mb#nz��..gY�q��ṳ���:�$
 ������;qե��.o9�,Ӳ��n��lӫ\m�]v3KŊ��_��^W|���c�x��������Nڨ��͛&�I9"���t�w9����t6�s�V/Gmɸi��\7I����Kı/�����Kı/����yı,{����bX�'����O"X�%��3�����ݙrm&��ND�,K����'�,K���٩Ȗ%�by�y���%�bX�ﳻS�,K��ܗ��p��ۛ2���'�,K���٩Ȗ%�by�y���%�bX�ﳻS�,Kľ��w��Kı>�[�nw%�7f�i��59ı,O=�;8�D�,K��wjr%�bX��~��<�bX����ND�,K�}��\��&��n�33gȖ%�b_���ND�,K����'�,K���٩Ȗ%�by�y���%�bX�̓��)�t$�<���;��\m�Voh.�'��;f{�c�l�^�X%]p���/KG��%�b{����yı,{����bX�'����O"X�%�~�;�9ı,O�����0ۦܦ�74�yı,{���������br%��y�Ӊ�Kı/���S�,K��߻���%�bX�3�3rKf�e.f�r%�bX�{�vq<�bX�%�����Kı=���q<�bX��ۦ�j�j�Q�͒����A�MݜO"X�@ X�}{`�	�͵i�Ms��	�kF�ͽ-��X�%��3�����n�6�wv�"X�%��wÉ�Kİ}�y�Ȗ%�by�y���%�bX�ﳻS�.��ow������F��)E��`������H.�s)��,N��;j��%ea���͚m�8�D�,K�����bX�'����O"X�%�~�;�9ı,K�wx�D�,K糧��rfa�2�M��ND�,K�{��'�,KĿ}�ڜ�bX�%�߻�O"X�%��{�ND�,K�}��\��M7dݖff�'�,KĿ}�ڜ�bX�%�߻�O"X�A9QO^�ND����ND�,K����O#���ow���]�˛���{��bX�%�߻�O"X�%��w�S�,K�����Kı/�gv�"X�%����3�t۔��ww��Kİ}��jr%�bX�{�vq<�bX�%�����Kı/����y��{��������jf"��ӆ�@h,uj
[�ֶ�[M�U�7.�V�m[-�[7r]�\ݚ��bX�'����O"X�%�~�;�9ı,K�wx�H�@�;])������j�ɹ�K�Zn�wgȖ%�b_���ND�,K����'�,K���٩Ȗ%�by�y���%�bX��>-��.�����2��ND�,K����'�,K���٩Ȗ%�by�y���%�bX�ﳻS�,K��ܗ��p�7nf�sw��Kİ}��jr%�bX�{�vq<��S"fTϾ��O<��3(y�#
�L�Ng�w7��LOs��{�?0|���z�tt������2�D��s��<��S"fTϾ��O<��3*dK����'�3*dL�>����yS"fTș�����Mݻ�!�,.�/B]�|�3<r��5�e�[�]zNrEL����H�N���`�����=��9S>�;�<�D̩�.{�sx�D̩�3(��vh~P'��ؙ�2'��?[�w�{��;ܧ���~���p���/K�S�*dLʙ�w7��?ݩ�3(������Tș�2'��?[��&eL��S>�;�<��S"t������n�rI��8�D̩�3(������Tș�2'�s����Lʙ2�}�wjy�L��S"g�w͜O"fTș�;�25�$��k����{��;����m�y2�D̩�}�ڞyS"fTș���gș�2&e{��O<���;�;{���
��ڠ����婑3*g�gv��Tș�2%�~�oș�2&e{��O<��3*dO~�;oș�2&eU7�Qh*�b����|��YYܙ�ۓp��as68ڭ�q���	�p�욬�3�Mn�"j�c�wD�<2�����3�eV�oq�a��B:���y�y�< ���q����h!\��T�v��6��(�9�[s�{v'����Q��w\����ݦ	���d�=�/X�94�67hC��Hh��%l�G����w�[���8�S��k:���N����揟�!#-�u�۷=��6�'m�z�K�����p��d�%���v�
�"��T{��Tș�2%ϻ�7��Lʙ2���f��Tș�2'�s����Lʙ2�}�wjy�L��S"{Ӝ���0�7nf�wvq<��S"fQ�����ʙ2�D��s��<��S"fTϾ��O<��3*dL������Lʙ2��Ky��rfa�2�M�٩�2&eL����m�y2�D̩�}�ڞyS"fTȗ=���O"fTș�}�;5<�D̩�/{��̝umt
������{��Q3ﳻS�*dLʙ�w7��Lʙ2���f��Tș�?�lO�短����S��r�����*������:[jy�L��S"\����<��S"fQ�����ʙ2�D��s��<��S"fT�~��O<��3*dN��~��$�M�����m��nX�R�
=I��<gs�u9ybf�^h�nz#N�쵾�7�Os2���f��Tș�2'�s����Lʙ2���w(~{�M��S"g�������S��r���o�ܭl�e�ûu<�D̩�=���O!�D�DN����3*n�=ʞyS"fTș�{��'�3*dL�>�{u<�D̩�.I��rnK�-7I���<��S"fTϾ��O<��3*dL������L����ݣ���u<�D̩�>�9��'�3*dLʙ=���6�sw%��̻�S�*dLʙ�w7��Lʙ2����O<��3*dO~�;oș�2&eL�����ʙ2�D��9m�˓n�2��w77��Lʙ2����O<��2%��F?w�~�ObX�%�{���9ı,Os߻�O"X�%�}�8����2nX��k�ĵ��=p��Xxg�>�v�kZ��4ጭ�::���bX�'��{x�D�,K��wjr%�bX��w8�D�,K��n�"X�%�ޝ��.Lܦ�i�ۙ�x�D�,K��wjr%�bX�ϻ��yı,s����bX�'�oݼO"�TȖ'���������v˓s7jr%�bX�����O"X�%��w�S�,�ł�z��D�O���x�D�,K�����"X�%���ݶfxi���Ci37x�D�,�BA�~���bX�'����O"X�%�~�;�9İ?�fD�{���<�b�ow���,�e��E��{��,O~߻x�D�,K��{����,Kľ����yı,s����#�����v����8s���;����z+V�[���7��,=>�9��d�-q~����ힾɹ�[��7I����%�bX����S�,K��=����%�bX>�{t?��2%�b{���x�D�,Kϥ�~�pӆe*=�oq�����?����<��?��M�`�?���"X�%��w���<�bX�%�����Kı<�[{�䙻Ksl���O"X�%��w�S�,K����oȖ?�XdL�{���9ı,O����'�,x��{���4���[Btt1{���x����Ȟ��߯Ȗ%�b^�?mND�,K����Ȗ%����@���7����Kı;���2���nɦ�nfm�yı,K��ݩȖ%�a�Ec������%�bX?g��S�,K����oȖ%�b_����`U.��������[%�ʃF�@ZwX(�;l��!�6��^kgNn��Kı=�~�q<�bX����ND�,K�w���
ObdKĽ�~ڜ�bX�'N���3�v]&k����Ȗ%�`�����?��@
�M�b}����O"X�%�~��Ȗ%�b{����y�r�D�?v��w$˚\͘\ݺ��bX�'�o�׉�Kı/�gv�"X� ��"dO����'�,K��?~���bX�'rO��f��s6�7I����K�偑3���S�,Kľ����yı,s����bX�ȟw��x���7���{�����\4�J�w"X�%�|���'�,K��;۩Ȗ%�b{�����%�bX�ﳻS�,K��o9އ��@di*�"�x��8�$�
T��e%)+@�PB�X���a�XE�`���3�uR@[i�sL� W��'�9��hH�#@#�>��	$���?�.��E�(�n���x^�����:ܘ� �ܸ��yM�wm���۞N;vq�B��$�6��2	N<$=��2��;�D��n�x��v��a��λA;&L��`8z������ǎ"�ܩ�ɦ,��(���fuMRd�� ��v��w:�i6�l����{n:�c���k����g�KJ;Pu�;�8z����@����hS8j982^v���h�ټ��:�hq����8i�zҹ��`�su�:�"Q���F^���/R�5�-�3U5m0��mͻ/)�u���9��I��c��UQ�8���HP.��b�.i���t��q�R���Ued9�r1�Zr��
���v��c�ʋkm�CvK
��MW[="��ڔ��<j���A�����u!��4<Ģ>Y��:��U��'#�&��W\v�k83���V�T�j�
�ࢩ�P�M�b��dɜ����FN:�TGnONj� ��1��I[8�1�Z�vviUxvR�m�@���lݓV4l9�[sm t�6�[[c����G�X:g\�:�l����=�sc*{!�KcW�]ێ1�(�2���aRmVc�b�,�(�Ѯy@�[�� q��5Х�v�f;�v:�� ��A\�A�In��e�ЯW��%�F���;�Q*ƺiIn�
�X�v�:'��h��1
���� scK�:0u�=�cJ�Sel�Zq��h.Is�E�{;l���p�(�3Usi䫝)���2��em�E�i�\�t���^���!�[ ؝�h�^���ur-S�d�x��t��88\��lp���96��Ꜫ�N��d1��l�v.�0�ۣn����@[����<k�a�h�^U.��ז�7\e��N�q��ۍ<G=l�U@UU*m�+�ch+�˹��K�U*�{L�H�"،k�si��UÐ�Wk����\�����)l�!w�]�n���-˳s3aoA�5�*�z0� �H�|'�� ���Bm�K2�,��˗3-͗�=`�zv	��p�=��ڮ�q�l�67��u��R�W]��hT��3�\�"Y9��t��g/[�Z���ĕ7T�'D���ֳ���`���d;f6�9�ƺ�g^s���'%��D�9��lM<.�h�Td1�y��'&��,��r:�-��"�0p{]��OU[������V���6ckkh�������H�v�X���63P=h6�n;���bfZ����w��|0;4p0E_��ı,K�~�u9ı,O~߻x�D�,K��wh~D�DȖ%��}����%�bX�;f���Lɸm�m6��ND�,K�w��O"X�%�~�;�9ı,Os߻�O"X�%��݊jƼ�^M&�Z����z>��k)�M4�s3oȖ%�b_߳�jr%�bX��w8�D�,K��n�"X�%����'�,K���ne.p�ݛ�d��ڜ�bY�T��>߻�8�D�,K����r%�bX�{���yİ? ̉��~ڜ�bX�'N��.g�lܓv�.�q<�bX����ND�,K�w��O"X�%�~�;�9ı,Os߻�O"X�%�����C�K#��E������6��D���m���W���[i�����{����>vF�m��۩�Kı=�~�O"X�%�~�;�9ı,Os߻���L�bQ>O{Ս@�@�d5oT��D�R-�n��yı,K��ݩ�b/���P�+C�My"X��w�q<�bX������Kı<�{���%��oq�x�b�dY���}���bX��w8�D�,K��n�"X�HdL������yı,K���Ȗ%�bwٿ[�ۘLݥ��]��'�,K��;۩Ȗ%�by�����Kı/�gv�"X��������Kı:v�ə���p۴�mͺ��bX�'��{x�D�,K�s���Ȗ%�b}�w�q<�bX����ND�,K�M��t�Mɶl�.m��Z�)��+*��p�˭�e�N�JV��U<$s'�t������oq�����U9ı,Os߻�O"X�%��w�C�g�2%�b{���x�D�,K���G?v^kgKG���7���{��߻�O!�E#�2%��~�u9ı,O~�߯Ȗ%�b_���ND�ʙ�������͛�i�s%��'�,K��?~���bX�'��{x�D���D"Ռ��'"dKϳ�S�,K��=�s��Kı?9�����#p�xh��oq�����O~��׉�Kı/{���"X�%��{�s��Kİ}���r%�bX��>;ٛ��3nSt��x�D�,K��wjr%�bX��w8�D�,K��f�"X�%����'�,K���69�MS���T7.�Cڵ��Uه^�$Ө�]y# sC�T�p�q1q2�]ݩȖ%�b{����yı,{����bX�'��{x��L�bX����S�,K������6�7inm�ss��Kİ}��jr��2%������yı,K���Ȗ%�b{����y�C*dK�l�˟��nv�M�٩Ȗ%�b{���x�D�,K��wjr%��2&D�>���yı,�o�Ȗ%�bw���eɛ���w&۹�x�D�,���3���S�,K��>���yı,{����bX���� ��O�FHD�_O�D��}x�D�,K����\��f��%���S�,K��=����%�bX>�{59ı,O=���<�bX�%�����Kı?� ���~?nf����f���������"��@6ڸ�>�2'mѰ�+l�!��s9K��6nI��̗w=O�X�%�������bX�'��{x�D�,K��wjr%�bX��w8�D�,K�^��!�4�͔��59ı,O=���<��"�r&D�/{���"X�C"dO����'�,K�������bX�'rO��ͦ�3nSt��x�D�,K��wjr%�bX��w8�D��R5"|�t��j�j���ŵ��oq��������.&A�J�w��@�d�6m���j�O6����v���[M��R��o"ĜB�M������N�Xf�X͛���0}Q�!�{��B�,���l�Y���k�װ9�P,���n�dk�o9{[ۻp��\��G�$�
J�a�j�=98�@�bb��n��۲t ���.��ݧhSh�+r�ռ��c����9yY9�*�l���6��OY@���[���Fvѳ�*N$85,�ӭ:��fԝ���ԯ|�ǷKx�ҕ 1��
b)ぜ�7���=�_��e5v���2��尉�{QJ�]����������<D��s�<�,!��z��Xf�X͟y��Ł�x�\ēPәD��1��vk����lǛ�@ft�@}q����Q���H�Q*\��4
����;�����.� �����ܦ��b�DDHrI;��(�����٠r�W�yVӸcMLmKDL�����%��t�<ފ�ҚmƋ�&��(ゃ�[1$�����s)�=�1�y�ŕ�ft´g�+[��UQ`f�X͛3���M6��O$9��E�s�:��QJ*�H���j���y�H��$�˼�(��t���y���jd��؏MDʚ��15T��O�}�ՠu�@�ޯ@�yFӨ�S�$�IA�I�Os���-w��;�)�[J��8�'2%��.�f��$�3z>3����@?ߝ��r�]	 f�m�lm9t����E��GmG�{BOM���ȷ+��sjb&hw��Δ�������4��X��p�$$�@�;�`��`dg6oɴ�^nd��f'�SҘU����Ͻ��Vy5�&��S�w�����5�=�A�K��Q3.��I���1��P{:Ps�h��Y9 �r5$�9vlP�,ή>�;� ]����b5�7F!(b��(� �n��՜R[ulh��=�Nsۚ१HL/3<�bg�.�t�>��tw�=�/�c��7����*U)UB(��,�wb��M(���oEw��~^I���u�X�Ȕn- ��~�.�zu��>�j�;��F��m�Ĳ7&����of��;],�wb�P��1&��fz�4gz�M�8�nd#���{:P��y=����-�lP^"�ˇ�*	�`�R��m]je�gc��b�m��K�dՁ��6ԣv��㧳2P\n� �͚���yy{��<P#W'�H8�p��&e��l��6ٵ���N�_�^m��C�G`��G1��iɠU���YM�v� �����*�o"ĜB�=��j3���r{ذ�mXy��q���tKm��<��E��hs�hmy��S��V����f֖?��
� ��~�&���,۲ff[3f�0Z�j.�q�w;\�u��l�V#�;knpS��F=��[�OX�#��;��@�;n��ax�ŋh-�����jj�K3u��d�UtI$��3�I���6�#���n��QA��x�d�bѴ�s]1$�-��WI��f�<�m�n,���(��������gcn�NU��:�6�/+�g9e��ۮ�{���4T�t�����nMJO.Z�m���m����Omu�I%j���9���:	c����ޚ�������$���/#���_Cp�DB�DH5134�͊�����y��y΀.�f�{���lջ�DE'���z{��hs�hu�@�ޯ@���i�1��,�!�}�u�����6(9{�I�uq@�_�~��Md�I�w[4]���)�}�ՠ^b��L�r$��.y��VT#��:���]`ڝ�Vֲf�]�n�������j7a�8�jI�^����e4�ڴ��h�䫉�$�$�.��$�{���PE8"���	�䚹+f����#9�~mD��D�&T�S"��"J�;� ]����~^�����?�ʵ�H�RdI�Q`�ڰ23�6ٵ���^mO6���/����&�x���.�z�I��o��g'�� Y��`u��gb#�^\N�n��n�pP���ڥ�<z�/t]��v�������z������ᒑ�����>�j��h��������C���"d�>��u�I&�fwM�7����Ҁ5�=�A�K��Q3.�����6(�{qm���hV�d���)a!YFQ�!%
Є%������
 /�@	@�1>ܑ�
R��,,[j[h[�e��(�&N��ۍ�x����8U+Y|�T�b`H��@LmU&32�A�b����J.@# )�A���L�����~�<t�e��R�ebЁIx����B���WӢ�"�qOP=1�C�F/�> �t�/�i'�[j�i?�ګ,�݋ �#�j�P����9�����FoE����>�j��h\~U���HbN����3kK�6��I4���F +��˽^��h���Ei8�8�׮�k��;������[�Ջ,)��&egQb�s	2c��p����hwz�������ay���˝DB��9R�	n"%��͚�y�oEy������%�f鯠pR�p�D�o�3@c��>��(�7] +�٠1fkN"�KĦ8��b�����:��/#���$=���$ T�)P-����,�.,�jb��r��Z �9�`dg6l�kKɥ��f{D��m��f.�7X����L������s�bӷ^t���V
l������ݞ����)�٣�2���r�W�}�S@���@/�&ʉQ.!C�����w����y��y΀�l�j�{1��F�X�&(�gJ��G{�K͋3�hy�Y�5*T)�KQ%�$���: Y��@[�ؠ������‴�6��Fb�28�ۋ@3�٠���O����9��`}��ؓtĜq��~=�t�]ҼVW���\��R�Mzvs�M��.�-�N�]��:�kR�L�v������[���P=<u��vAz��^��#;a�Y3��L7H�%�!���<��3��&9���Y������9ug�Y�wJ	�՛��zW2r�/>ظ�s��-)���v����#�K�3d�`�4��
M��]���T��{���/�Uؔ�Ɔ	����:�FZ6*LZ�m�{vw���m����{1�V���m<��I(��/_�@��Ҁ��u����^oM�w���NX���R=�����;V�g��4����&כm̝P���*���
�RP�������ooEy�� j1j{"��&!��Dˠ����W��@yz�z��M�v� �/"�e)��D�U���ٰ=����6}����f�s����q�5�bM�Ƴ[�&&��i6�-���"�Oڢ�l�2�I�q�w�4�ڴ;�g����a�7���m�Dʕ
dR�D�`g'��v!�i'6�$BI�2�RҦ�o�$X)�����f������Q��#22dq!��gvl��6(�y�Ξ(��ta�`�T�)Q2�����~K�y�f�P�<P\n��M���5n�QI���C���w����Y��� Y��@[��@��
���$n4��,�Ɛ�`�rv���E7��uŪ��'zX�j�GS�d���th�L����Z����Z�ٟ ��x�F.O�R�D�52��t ��g@�ֽs�h�y
�`�JSQR�&����ٰ>ͭ,BM��ՠ�z����r'�E�1H��>��(�7] +�٠���FoEi`'�	2c��p�>�j�?f/&�7��1��P^Δ�<5���k;ti��3c���b�^3�[\�kR;q�z��u�S����^��u��V?�m��_�@�ޯ@�����;V���*��q�&A/��.�z�e4�ڨ]��~�M��y����O���b���※��G�ř�4<�SX
�Ǒc��I���;��@3��hOo�w9'W�̔ �?~@�|�z7�>G,O�R�D�52��t ��f���ޏ������u��^O�����a���l���1��så��n�;J��"%����T�u�ss�����{6����̝��I?4�@\�z���B�dlQ�5"J8��Jht�ŀ/�v�������ս��S*(�7�y΀ّ |���連��#o.Fd�2(�ۋ@3�h�6(��(9/y�Os�3V����5&A/��.�zw�4�ڴ>�f������R�&Ү�'V��Ry�l=ZqD���[� ��3�GBs��!ĩ��.w�����[^h�E�{T�g�P�{m�����9���5��FY�%����ҵ�T�[�����\02��6�S�-8]�l����ۣ�K36:
��ݧI�X�詷�t��Ū��ͺ��R.r��Ѹs�&8\]7J+�4j��ku��i��v04���M�����W+$�����6��8�.�aw���Q�h����w������HdPR?}�~4�ڴ>�f�˽^��Y�+�&Dɍ�I�v� _^���v(��+����9�.O�R�C��"e��ޚ����������̎�@m���&Iq.#��U�Si?&�jv�ޛ���`fN�h}޳@����ء"nD���^N��n� _^���v(������޴��i2؜�=�\�N�qWl%E+qx7Wgqx�EgCڎ*6�����\}���f�=FE��p���h}���Z��Jh��yr3#��$6�������o]M6�U$�w�`s�],�݋��U7�p�L$�_�94]k�:�t��o2;� +��1fk�"���
�TQSa��k�$�Jw{���>�h}���7��b��\�2'�)TXd�Ł��M/&�iJ��ՀU��wzS@=}�.Fے8E� �E;��6���nt�R.1n�cW�� �SN�����LM��I��h}޳@�ֽ������Z��W9�8����-��Wyyyy��g�2;� /�6h\~B�$��	$z��M�s���<TE��)����Ȁ{�~���9�~�Vd�F�eJ�%�j"$�;��@3���.��w�4gx��Z�ET�** ��� _g6�4�Kɦ��ޜ���`fN�Xl��� K��
�z���]/�d��a��XƳgC�W[�Zur\�ݡ��E_m���ٰ>ͭ,�ݎ��� \�{V��pDRq1"�#���gJ��6fGs���4�݊��ɬC���SpL"fJ2;� +�٣�^I�y�gO����S�s�DL� _^�X�6g+KM��C}M�����@?xT_������@�ֽ�Қs�h}���r����+Y�l���Y��x5n�֭��W�h�mӜ��vib�1t��p��O�o���Δ�n� _^������y�,��`�2L�"��4�j��h�v(��+��K͚�I���`S(�D��Z���4]k�>�)�w;���X��ⓗ22��33A��O#;�`g6�X��M6��Y��X�&7�����	Ǡ}ޔ�;��@כ4�͊��Hm�Mi�
�	#H�:g��F#!Q 1"��}�ŉ*"QA5 � ���C	a��[�̄əHHL����JB���$��J��Ie����X���BD�c��'��	�#:���
J��J��BE���b�%8�L4�(�f��c9����&k.i�ݎ&�d�
�Bm�j�c��<]����V��Gl�\���\a��=�t��؉�I�a��i{{<��e�5g;��9�q1O=b�76ګO6m�d	Z뵞�&���G�>[�n�:�hh�/Kf����������^]l�nX;k���v��;[�oF���s5���l�Dv�����e������n����0��,օ/[7�n��ʠn���j��I��c3��P�26��Z7�un��N�n��Kd���Ĵ�=;sj�8.���mC�؎Ħ���&D��5�P6���Ev�����+(-�v���d�R���2������yj�8��	V�&��A�u5�U�t�-�J�cۦ�xm�4�Mv8��W-��Xܖ��[Z�;^ˇ[q��� =����.!,��{\b5�ضuS.�x��J;;��K``�Zs��kcq�9�f`�A�����.�KM��g&N�r�K�4��:��v�D,��#P��kt�9���4d٢�F�mVii�\G`1֝K��탦�b�;���Y!�G�WTm��V�%�Ȋ'b��E����]���Ĳn3׷j9�e[�Xm��W��Fu/k�8�Q�Z��7�R[�r��iշm6�B��;�[�.cl�Dʪ�tҒ�\� ���t�R7n�yS�ck$KU�nu��nݺ��l!e�J�nm�&뎌&����'�i�؅4�tM��[/N���v��U5�U��˒��eh�H�j[���m���ySj��@YbuիqL�R����QD�u�F��6T�hs%�e��N�u�ZQ6�J�ym�^��Ƭ��ƭ�1��Nuv�M��v�81W;�/<���틝������q��ڢqv�rD�oK�F�h�
�	
��rYB�!r8WnjU���|f�`"T���!����1�V��[d�xbU皥.zu)!ꫠ.7*8-�ٞ���T:>��j��D~DU��QV1�G����rs�;�5��p�\�$A-ۊ�6-�g�	Xϳh8�\��]�d��e�]O��`4˵�O"���ª
�{I��0�ӆ�v\h��\kPr�l1�bE�h����nb�UI��x��e���Pa�G.I������N��(��7<��^�pv�P)�W]m�����/\��%��s:��)�=�c�8h+&x���{���>���:dB����6MZ��Rۓn˸�5v�Et�&5``G��)�$�F��Hhs�h�7j���l���o�sk���]Q�!17Y&E��[4]���N�����/yy��ON�$2�"[x9&���ߞ���M�ڴ>�f����+��8�	��G�wzS@��@
�vh;�I{�#;��՛!ȉ%L�jZ��(��t�5��?�;���e4�*��I���2	�1����4�a�(�X�m�������q��O�����r�m��fI��H���{߿M�Z���?//{�/�fGs�3V�m8��̒(���ɠr�^��fc�gK)�{њ�]��~�^I�V�8")8NfH�	Ǡ{ߧ�@�v� ��f�˭zŝ��rA<��	!�w;V�g^���v(9{�y�\P�'�INc$�ȴ;��.�zu��>�j�?����ߵ��&A9C�����MYP��s�u�]��A|�w��- s���\���v����
L����RN�����)�}�u�^�K����F��I�$�N"BG��e4�ڴ;��.�{��^l՛!șR�T�-C�t�w: Y��`�mC���́�;�`g"�aj�D�.�DD����I���4<�́�;�aԒi/6��~�X���B��QL��k�'&�˽^���Z��Z����y&�IL��D�$�q�pP�Z[�CӰ��jq������5��P,���=}����"���8���-�ڴ;��.��v%r�bn!���:�7]~�`�;��ǝ�@]���M��'�IN"`�e2�fwMn�b��^^o3��2;����TD�9��椚.���S@�v��ƚ�וR�w�`s�uGf���*�L�UH��)�w;V�gu�@�ޯ@��̘��sD���(�׮����ݎm��/۾��`֞U�1ڥĬ�!�X�����͸|y���;��.�zu��;��yr9����;����G���������u�/%���_6ȥ�LK���f�Ǜ�@]��G{�^n�;��g����=��M���)LN
G�wYM�v� ��f�˽^�qg$�jp8Q0D�"d�>��t{�ɬ���y��Δ/yyl#^-h$��3=�=s���z�A�8=f�2@j���;=�^�r�պ�&8�S71�;G8�M'4���5�f�dh�$��ݸ���,�^���s�c�R�ʷ-KuqM�1�����iGp���;'>JLJ� �V�`L9�X�����X�Ν�m��+�v�$d9g�'�t�j휗�7����c��,��p�*ƃ;`�������ph�.���6�[����y���c���;^���&�l�lu�ָ[��	"��~�4]���)�}�ՠTy\n ���M�RM�z���hs�hw[7���ø�8�ǊDہ#�@��OƁ�;V�gw��9w��=��I�#��C"��4�ڴ;�f�˽^��YM��Q�r#dMD��Z�޳@�ޯ@�������9%�y�;\t(��r�d����PnY���n�K��m�[v���V���K��9�)��_�I>����>�)�}�ՠ��4g�Si�7�5��H�$���g18�D�T��nO~�v�}�Y�r�W�\Y�+�4����hs�hw[4]���)�Tˊ�&&�&��H�;��.�zu��>�j��<�`���M�RM�z���hs�hwz϶ߝ�?�w���'V��o��$V�������5]��nOД��ظ�.x�X8���hs�h}޳@�ޯ@�=��<�$2,m�@���@3�h���ޔ�;��w"1�y$��fj,}��`dg6l�m�Җ�^�^n�'J.3]�c���\��dk��M�Z��Jh�ՠ�l�=��M���(H`��zu��;��@3�h�נ}�$ǊH�b��kC)�m[.pV�ӈ����:h�%�㬒�yۦ)2bBy1�Oc�!�w;V�g�l�9u�@����Pv\V1752��t ��٬_��^�36x�<�}w�F�<�^ٛ�f鹛s	���y{���ޔ�>�j������F��
���
����^I����,l�^I!���@�A@��B Lm!jiQw6��"'QR�J�F6�}�ՠ�z��z�����|x��M0N$����x�c��+�ܙi5�k&n[B�W������|��F��ۋ��_�@�ޯ@��)�}�ՠ{Ǖ��dd�_Ēh��(�'J��@�͚�yy6j����q��A������v� ϻ�h���ŞB�q�X<�I���>�݋ _f�X͛��Q�m��9��O�R�A0)�Lˠ���n�^���M�v���Qe�'��G����=������c,vm��l����n�w76c��&�ˋb�����Bꧪ�[up2��%�K7DQ^+a9e.����x�ؒ���)noO[�$��X�8��k��j�u��n�%ݹ�3�l�T���������������8�ɹt�M�ݬ���[��4q�&%w���n$��=�;$z� A��D����]��{�j�z�K�6]� Q&�z.�[H�\�s��v�6��R��	��ٮ���d�W�r9��3����N�~���s}�=��G��)MUJ&U)���;�)�}�ՠ�[4]��Ǡ��*���L��;�`�ݫ<�Iy4�s;�M����`qs�1��SRۋ@3���.�z��M�v��<�&�$O&9��$�9w��M�ךM6����͟z,}�ڽ�������9�.���nb�t6Vj����hÚ���l�ZwZj&��D(ܶL݅#�>�Jhs�h}޳@�ޯ@��m��
&PL�&J��O��|�Eh��ƫ���/�A����1��P^N���y&Ñ���	��3$�H�;���9w���%޳�w���@��ʡ�L����ܚMy4�S�����׋�ذ�sf����UĦI"����@��)�}�ՠ�z��z��/�tƱ8¶n�{/6�lj�b*)[�M�x��m�Oj8�H���j��"f�T���D�����t ��٠-�lP^N�,�qT�Ǔۋ@3���.�z��J��]�yy&��_Cp�D8R�e�說�9�́�r�����h���߾�|�UaV1���R%L���`$H:���@E% q�Bp��D�$`�J�jā[YL �@���B,D�F,da
6(� 		d$A�FEK�`D 1 �j��V����!�F0 � �FOrB�����x��MD7ʂ1��ĩ�=�om�9F7ߑ_���hM>}	YFRR��2	1����'���꾞x?"�A�!���tE+��|*�p>P8܌�@/6hY��DR���'Ñ�����@}q��}y�A�^�I�f�P���\�CD�	�D�@}q��}޳@�ޯ@��)��/QH��8J]ܵ �^�nJ��M1o9eHz6��^�5�$:SN�H��Ls�b�S�L$�@3���.�́�r��i�4��l��`s�zz	�	&D�o�nM�Z��Қs�h}޳@���*�S$�`�LrG�}y:Pq���/6+��1�tW���l�#��S*Ij"$��{�2{� +��X͛��CI�m_+s���ݨ�W	���c�#qh}޳@�g�����?��Z\y�19dM(�W<��	��ԡْ� �d�:����X���M���Ӏ�B1I&�˽^��zS@���@3����ީ6�"�0sBj���9Z_�m��9=�X�oj���خIy&�Mjo�)P�2
e2P���}y�@[�ؠ>��(Q���b�)�&E��z��z������;V������'�rh�6(I%y���^Gs���� }�a J�	�
�s1TtG����?8��ڕ��;m�m^�=j�jv쩚�@rg�Nm��9�c;�oon����y\��nx��}�������6��#���:�ۗn	w	�NӺ�#q�`B�Xy�iv�1&��C���'M���Yٶ��:��n��b1�3��>�ƀ~X����+N[s�Nw�|��'-FN�����:5ӋU��ͥ��ݓ��f{\�wtX2:nb���N�ul�λlg���i���F��0��Wf�S#Ȝnd�,���=l�hs�h}޳@�ޯ@�=��)��Ɯ4�ڴ>�Y�r�W�}ޔ�=�Ѷ��Ǆ�F����f�˽^��zS@���@�g�i5��y1Ȅb�M�z��Қ��Z�u�@�{�&��X�8�(7���M�ڴ>�Y�r�W�P�/�1HFK2��;4n�knra�M�J���3m��Y�����qa��&5��D'!�}�ՠ�z��z�����P{��LQ��f��{�w��D��-��� �zS@���@>��q�y �o��������G��$����@
��������Y188��Қ��Z�w��9w��/�A7qG�a2D���v� ϻ�h���w�4�U�d�rI#"O�i�g[�ɭ1ò���9��6�؅�	�vEs[��J�k�@� ��Z�w��9u�@��)����3#���_CQ�p�L����n�b��Iyy��g�2;� /�,��-��or$L�$(7�޳�fN�Ym$��.�T��߫�`ln�lMf��T�Բ}2��(9/$�d�: ���4]k�>�Jhaq��5�`�Z�w��9u�@��)�w;V���?��q���q����Q�N��/�wsm��4 �I�E�nJ�4�[]]��A����^���w�4�j���f������'���$zד�sfdw: W��@[�خI���&�"<r	H�4�{����[4�7�;������LD=	PL�d�Ɉ�A���M�oM�;����t�^I��AUhb��-:�਄_�MTw7|��y���S3���#k�h�נ}ޔ�;��@>�[������P<�n�
�ꝓjܚ[�Fz�[u�;���q��\�˗Eej9�V�u"Ġ�z��M�ڴ���.��Ş�N�Ă@��r��Z�z��z�����Pv���R	%�2��͚�����w�<P�����{� G�&���9w�P^N����������5s���l�	�rG�}ޔ�>�j���h�6(~9{��G65.���"fk�8ɮQ�U��Z��F�1ub�^)��\/Q���ݶ�L���4�TOk<�d9�v�V��ٱ��tf�e9�ŋf�U.u��;:��KГ��I$5� �9�̥?��˾��w;F�@3�3a!��A�xh�=
�;]r�Ņ��<��=v�؎�C�L�9��*��/�)6ɱ]�ru�y\��c=(7nϿ��_{=�m�i����H��z�EX8"3�+럀9�ΛY̹&.ee-,b�ƞh
�>z?��@^l��6?�����ձ��a1��D�A�������#����;��Z��Z{<�X��I㐍�RI�r�W�}��hs�h��4��I���$��q�s�Z��Z�z��z�س�iܘ�HE�}�ՠu�@�ޯ@�~�@8��AD9#��L�,LId�;�Q�:�W��G�M��wi&��S&:�/Gg��fX�"��٠r�W�w?U�}�ՠ��+�@�$M�ɠr�W��g�yG�1����t���w�e�\�[��"��@�;�hs�h��4]����M�G��F��>�j���h�ס��z_�@�ʣo�DH��@>�Y�r�W�}��hs�h=�exڌ�D�Q� 7������.�&�5���.��C��!,���X����dqF�)$�9w��>���ڽ� ;��.{�6��i��"J	Ǡ|���?yh�l�9w��=�=X�LH���	"�>�j���h��;(H���"=TO<���I=�>�@�;��L��8�'"���h�v(�3]{��{��WA!0�a��������ד���;� }޳@�s^���r)�k$o�,`��Jj����I��X8�Ou�v8f�u��<��$Bpr94�����V�}޳@>���z	����7��?W@^l�ۻ4����I�ys�����0�"Pn- �_�@>���~�@����;�K�I�&��$�Fń�O6,�݋	�MB��9iyy7y�4+�n")9p�L�nG3��V���Z�z��z�����nj[%\��:ڶ���KK���F�Bz�nò�f�8r7\�i�Q��7] }{�@[���a�΀��Qޕ1�LK"e�׻5͘�z(y��@���@�ײ���7���@�ޯ@�~�@���@>�f����*q���N�=����v� ���.�z�=�Dx��6��>�j���h���s�Z��H�)P�ԙ*?�R/�{�"�`1HF�F+����Y,$Q# ����� �- Ё �d!$d ��!@�т#	BXVBBQ%�B,YBVw"~��Ķ��^�q�ZF���`�9��K�o9xB��BRۄa�e*�U���	��m�,�"�(j�W��o���1c��!@�$$ E��ߝ_]�4O�߲L�7&nC3M̳s��X:���]��Ae��#����m�C�n�D˷9�P��vM�4��-�e���lw<ú���f����
� ���v�
h��mm�:[A�λ�&ێ��Wnb�@㠝g[�>[˧i�CG�3��\��v �l��-�V�8d� �V�=��{}�`̕�[��3�:I��RnА�i'mFGLa��-��0���iL�*%w�7jیq����4H�i�j�|/>���m�����g���'�#�F6�DC���
�v��<�Ɪ�P�68�Y�/�j��]����ᡇnū
�W�uKʖ|��LL�T��.��ʼ��p@PSd��4�KQT(�g�w-Z�%Y�۲�s�Ppq������YTֶ��<�(�N\6���;I�ι9�;kuGNh�DL\";H���D�j�ܞvU�9PݷCR���.1�>v\��.y��l�d��]x�Va���u�Ż��p=ɹL�`��NZ�]��+��\�=m-��Ԇ6T"��֐�(�]n��V�]��b�N{�Nr�a;.�WKoSj�Ea�a5�f9���j����NWmYÃ��(���RF�v^^�c0=�z.ٺ</8�UYV�`-��Jep19B-��`�R�:��B�K[[�-��U������8�۶+�QGc��z�&UU7#T�t3Ő	��mkn�l�[�t�x���InwB�c�<hܛϛOȝm�u�^5���pnT���/�gY8�I7��;z�������-�\�_�fd��Y�3��tC��p��x�vM��/+;������6(�+Z��E��n�BPv�0OK�4�-vT3spj���o��\�AdQ�~��K�J4Kݬ9u�m.7�ۈ��]Ƕ�N8:}<��ۮ��:qc�9r5Y��mV=�h�7%-�m� ���;vBZLl@Q`\cx�V ̛Z�Ɋ���4��m,���%j��� �˵Qu79(�9�S:i��f���Kv�Sv���#��=Q���P����'ʉQ�w�����@(��R*�"G ��J!����/`�����Iuۣ��˱`��\�p]��ٞ������(�5׹k��0�g˶$3�1�D7@slc<�E��Lz������y�{k��"1���=��U2��M`��/e��v�ٴ
Z��zH��n0'J��4ChRݕ٣��&�	��c��uY�-��]j�96��t�J�{�߾�ww}֧�Msm�a���0�힧��X�][��ECHA��ڋ%<3Es	��	(7�=߿M�Z�����ڴ{�T�=��rD�X��@�ֽ�~�@�v� ��f�s�D��Q<�$IAH�����7]��l�ޚwE����C$b#�H��j���h�נ}��h��������r- ��f����#;��/#y�q���{�ێJ�]���:������u��Z��5�m��d�<ī�L�떶[K���m�k�>���j���h{��)��e͓7w9$�����z�TqԒI��W�sj���l�[M�s�X&�"<n"8,�Šw���@>�Y�r�W�}��h{<�n�?�xFAB"] }y�@[�ؠ>��t�y=΀���7�po�4�)$�9w��>���ڴ������c�E24�����V&f�����koN��׻���9�4]��	ۘ�y!#J	Ǡ}��hs��כ<��1�tP��"#��dL6L"f]w���$���1�tPs�Zp������Z�zՁ���`�v�mI�nRnL��Ł�?U�}Y�܀�#y�94]k�>���j���h{��)H8������@s���̎��z���l�.z�Ѧ8�q6�n���j�5]�,��Ʌ���.E�6ܯjZ�y��Dx��,�Šw;V�}޳@;����V��Q�p��<# ��]�خ����a��4�o:�7V��y*�Ǹ7�d�IG����~�@�v� �[4��&���əm�s3A�O6{��΀/7f�� @�/��]����'�>����ƚ��<$�@�v� �[4]k�;�ՠyvy'��ۄ�ic�!���X��b��R!�3i�mu�I�t:r[O��7\Ljb��H��l�9u�@�;V���Z՞ˍ��7��NI�r�\��y�6;��΀/7f��b��N�qǠw��@�v�?fbI6f�M fwM��G��Ne
VD��;��@;�� �h�j�=��t'��(7�w���v���Ł�;�`[m%�|T���B���;N�6]�6�6\Ptu�������r��㱶�n�3w7l\ݽ;&����=�A��n�Iv�1!�ꛄ�߾���{-�gh�LO%q�@]eT����9��H�x����N��ֲ���Obnm�&ބ%�U3��1�>5�m�y8��G�}�d�v�7n��8a��ݝ�/ca����(q�议|���������<Q3��|ɲ���&今�yٶ�ֲ�>^ff8�&�Xn,�㵁���4M$���9�1&D���~�yڴ�j���@�ޢm�(�Lr	d���/#u��&���t��4w�5�{͜��Q�T8sɄLˠ3#��z٠����Zp�Ʉb���H��l��f��v��ؽ����������F�6��@;��yڴ�j���@�_�c��%G		�SmҜ�ݮͷ&���+/b0�=�tV�L==�u�	5�������@�v� �[4�٠}��&�ȪEJ�UQ`fN�Zoi�	���9w��;�ՠ{;�mП�L���q��vhw�w�͎�@^Gs�;��I���9�1&D��9w��;�ՠ}�ՠ�f�s�RMnH�L���b����@w�'����4�ݍ�vW��!#�'NDD�����͜�b:H�u�hgM�
�V��f27\�R`�Zs�hz٠��� ��:���j9G)D��02�7�h�٠w��@�v� ���q��ID*���� �ݫ9;�gk4�����R�NRMq��M�Xo6������pɍ��rh�j�;��@;�� �hx�I���I�yD��>�j���@�ޯ@�;V��Y�~U�Kv��p�<V��Ѭ79�Q�:�V3WCG�V��SpiC��$Yhz٠r�W�w��@���@���RB)�"rh����j�>�j����ީ&�y29�AH�yڴ�ڴ��@;�f�qv2"5Jn%�e2�9//y;��t���`�ڰڦ��Bi�$4!��H�I���� �!B,c� 1�� �"",",`��b)"�a�zi�% �È"��\���$��='�;����I�u�hw��=�j�>��t%䗷�y4@�B	S2���C���7�j�÷R:�]ru�2[��%)�"dC�2d�YRI��M�v���h\~ʜr	�&7Qɠ{��@����u����7��G�X�����<�"qh����� ���s�h�x�vD�8D�H�P����6(��t��y�Ɓ�U�b{���d�M�z�2wb��6���ڰ>T���lI%��o̶e�W0��\[p�*�	��KI:T�K�#��X܏n���I�<bki&W����mtmv�e:9��!�4�,l�n���N�Sb���[o�sGE
�5�Yf`�9�o];���Ar�q��З*� 7=���ʗ�^�B`3���VnүR�\�mN5%�v4\��+�4gA��;��*
�q��p�d�n�r��%����P~s=�T�n�Sb�:�gsy7l5��[u�3�M���:�rJ�M��-��79�jTŁ��s�>��(�v|�oE���i�ɍ8�jL�@���@;��.�zs�h��\w&
b��	"��f�˽^���Z��Z�G���L�(�FҒhw��;��@��u�w��y��@��:%�
S��M�ڴ�ڴ�٠޳C]�����ߝ�-�vŕƍ�4V��������V�E��]s=2��&qܮ+��Y�������������Z,�G���2C�Ɉ�@{�R��%�-E8�"�	d�����y�w��O=v���S{���$��&�wz��ڴ�ڴ�٠{�V�[�29�dRM�ڴ�ڴ����Y�\^�w&4�!�0r-�v� �l��f��;V�gx�O"$�Ӻ���u;��8����i^[����ϳv�)��s��2`�#2L$�@:�4�٠{�ՠw;V�}Q쩩�#�'����l�;�ՠw;V�w��x^ʜsjpjI4�l��s���qQ���>q �(��j����!^&(lU�� A�D-(��TS�����
��$a(Ĥĩ�����B*������*�)� ��D�A$�D�d(�$��a����
X0HDd���� @bD"�FA�L�
,��(�(��:ă1�a�*G� ��A�B�P��dcYp"P�ێ�5 4La�q54x�!Ճ��#�"� F{'�B�"E�:L�.LV�����B0���Q�u~F �D�UD*���b:'}E}b+�����%E@��_<�N�9/����[4�z"���I�yD���ff<��t��4w�4dn�,Ʉ�ȔHE�����@�ֽ�v��ڴ��ŕ�j2C)Rn
a�o`�nJ����u�Ѩ3k����gt��bܧ1��4�5$�9u�@���@�{�����;�nI0�NeG3dn��7] ^��n�b�$��g'�Ȉ�)�Rȉ�Dˠ3#���@�ޯ@���@.��`
"3&Bf] ^��n�b�̍�Aػ�B ,>G�+�	s����$��z~ML�Q<��$��Y�{�ՠ}�ՠm���.k_�6�S�H�x�۵n�c0���q\Eь魸@�eb˵\���bC�NI'�Z�~Z��Z{�<���`fwMxl��S�)S51���u���a��4��4dn�����f��nHQ*\�."] gwM �h�h�ՠw�*cOq��4�5$��f��;V��;V�u�h�դ�㍓�,�I�{��Xd�ŀf�j���l�m$�	����޻�����j@k\U�m(��d���,w<\�d��mX�R��V���+n����q=C�n3�����Z8��睇�|An���c��1bn�P	q��]a����4��[cLm�[F��#��`��]n'1��ۇ�A���M�b�--�zJ��4$�t�OH�[��Z� u����pi�gE��8���p�V��v���[t��nYL�nK��
�� y��%���T�F��靟[Wa�.`��*�s�n�70�tu��m�#7p�V�f�Oj���џ� ^��n�b�ˍ�@�F�����$Z��h����j�;���^K�P�L�(�F�rh�נ{��@�v� �h�^ʚ���zs�h�ՠ���Z�q��&��dyD��;��@;�f�˭z��Z�?<,sק��e,N7N��H��[�O1T�d�E�JLL�z�Z��7DX�lw[4��h�ՠ}�ՠw�*cSjfUQU1�f��39�r�O!�[B�
A]��s����'�g�גC�٠{�V�[�6LRȤ�s�hs�hu�@;�f�q_!�rb@��$Z��Z�l��Y�]��?��� L`�3/���Xf�X��d�Ł֛k�����#j]���6�ix��'/KTvz��j��J�ڷHmAQ�Fka�^�*� fwMw�����@{�@c�SRbY"I����;��@�v� �hu�@���bll��D��3'v,3v��L$�&�4���$�IG��_�%�tP���œ
#f[��H(��@;��.���ՠw;V���=��HH�Xۓ@�ֽ�ڴ�ڴ�٠yTee�Uͪ���ԔJɎk=\�79�-�m���i�����u�"�������?�hs�hu�@;�f�q_!�rb@��$Z��Z�l��Y�w;V�P{�����H��٠޳@�v��v� �����	̍�m)&�wz��ڴ�jИ �j �>��{��O��쩩1(A'��@�v��v� �hw��?�ߑ�<m�S��ԊE��W��؊�M���Cel���*�-9{ui�����9�"Ȝ_��- �hw��;��@�����Ƙ��$Mˠ�٠�٠.�u�\n��/y�֋�=���H��7&�{���;�룽���w: �����'.�q"�h�ՠw;V�w[4�٠\W�mܘ��AE�w;V�fnՀfnՁ�;�`jocM!r:�~p�,hs�<����75��ແ�1���	\�:�/KrG�oN��9�S��@ v�{j�o���������gO� ��J�����q�K*8H�M��t�Ã[�sn�nv��G�E��We�����^�e�9���^�gh	�*F8���ʜ����\T;�ݼ�GN�w8��*p �۰c��-�C�*v��s�N� A���-�,7r\���T�ȩ�+�����˙��a�Q�ӎ���L�{=P�	�{V��)!)�b���k���g�|o�M ���s�hs�h何@Ndo#iI4]���j�>�j��f�^���ĲD���@�v��v� �h���{=N1�H��Y�@���@;��.�zs�h��ln�LL���@;��.�zs�hs�ho�����#�'iĪ��f�X���ϖ
�h.*�d�n�1�X+�܍��ᩈ��-�lPq���7_�{��g~��_�mn(�Ȕc����ծ�#h�څ
qE?�S$�������4]�����&D5&E�}�S@;��.�zs�h����Q�i��w[4/Z��j�>�j�/5�rs"yĤ�.�zs�hs�hu�@�w��_����`)�������yQ�v۵����^���TYt��XH�%r�t�l�?ߖ��;V�w[4]������ؤJ8��@���@;��.�zs�h��ln�LN!L������ڰ23�6C��i%��ߟSM���IW׳�b���;8r6c��R1,�ɠr�W�w;V��;V�w[4x�1�䐍�#�;��@���@;��.�z�2��?n;<V��6�q��3n�+QSDQ�	9�E�xE+��Mr�f2��:2WfE������f�˽^���Zp�\N�i��H��٠r�W�w;V��;V��g����D�7�I4]���j�>�j��f�}SŮ���ĄLLPr���̞�@_'�� �ݫ
I$���M�����uQ
';���䓽;���ə.ͻv�7��;V�w[4]k�;��@��n��~j�L�f�yEN�P�x�����N��ԃZ)���n��6uĹnGb�q% ]��n�b�����%�ft�4j_���y!#FF��9u�@�v���hu�@��*��O$dm8'���Zu���f�˭z�|�݀�&&I��h�S@;��.���ՠˉ��LBq2P�����K�';��ݎ�$�Ϸ��'��
����
���*����*���T��PTW�UAQ_��AQ_�_��AQX�����T��T��PTW�*+UAQ_PTW�AQ_�UE�T��PTW��AQ_�UE}UE�1AY&SY�>8S�Y�pP��3'� ah�                        ��
EU%!@�P��T�DJ"�P$�U�
T 

T�  �� P�$��DE@J� 8  hP  
 (P ��=�/������g�9=;���>�p =��}�^�=9wo��ON�x�ON iv���s���|{��s4p 3�ӽ�m��>��     z� >����O}����r���7J<  �@  E(� @Wz��{^�M)�w8�k �u=;��vu���u��>�/ :�U�U3��� �}�_O{:<zW�;�zSɮ��!g�=g����9����}��*�[�{�� y@  @
  �h���o6�������,��x�xx� X  
�4�P @  � E   @	 �� $P  � �@"� � @  � 
 P   � 0 � ��   Ю�}���g�8��3��>� ���w�9q;���  >����S�ݩ}� 8r�u�q�����=t���s�Kũӛu���Ε�w)�  � ( T
(  �����gA�ݾ��Yy��t��
Y������˳qe�o�{�3�����  �w��^�^����4���\^��o��ϱ�m�Ϧ���2��zy5�㴽n.�/ C�7��J� h�HM�JJ�0 �O��&�� �ت��Ғ�  T�Д{T�* �"$5%"D 4f�����������������w����w��������*+��*��*+�A@TW� �@DAS���?�����$��@��Hk�g9����s�����cd1 Jc
A,�4�	<�g��s��/		D�ї��f2��P�6�ny�O�V4\XT$p�3|<� K��
B��n˺]�%�y���ˌ��������x˅f�l��l�X�x��
�y, J��_�r�sR]72���LA� �`D�bSp��ya�LcLYbxŌH���u�ÇF,	��Q�$ F,B&�!���@��ݞ���,��F8��k�=���<�{�B�	�X�0��<fs�<43\����8˜=�$ᒘˁ��
��(��0�
��$�3(L��d+�Č.FJ�24��ÚK��=��y=��l�	fhJJ3t�fp��$B��M/	 �(jqR5e���p�c�,�B{�Ǔ^ė��J5��F�ILԅ3@����[�f��
hXV@��d���a�,J�a)��0!��Ѕ14�0��Vno2\Á%H� ��x��d5�g�@��B`B�!
�!��m��fdݧ!C�����8`@�'-��!LH\оϵ�����.�=�>��=%ĄVaR\����y�8�c�)�<��O}�7�)���o�3�L��YO1��Ӟ����l�� x�;7|����.��^�ݽ��f�����x�$+�{>W�ۧ�[^�<w��qyJ����fw��yHT�>+;k{=�]W��M:zVQ��t/m�/%k�/���/�7����2��bį�-ʕ^�Yuř��җ�~���{������^o������9��
�$��C�|���GF5M/�=�g�S	% b@�3g4ep!L!L4���0�)�0��� �rn`J��5�qe9m�Ӑ�!�w���³�$����`F��
`KL����1 ˜፱��B$��|,9���L�Y0k,Jn�3 K�Nn%hF��F77��ĉ��4�!B�W���F�'�cd-BaMeX\�O<3]<8����`:!�p�@CXH@"�X��b�
�4�4�B#b�"��"a1H0��c�J`��k(�l"�H�)�X��01ԍr[}�������	�k�	���vI�Y�2c%��!xc/��In�'I�����	���
B�a�4�3w��))��$�Hf2�	+
B�B�.`K�.BK�K�	(B���K�́,2IO9�H^�>���OvӇ|�=�r����,7�x���Zi74�81a�Is8��Ҙa7���$�� ��@�hJb\0����=����y��W��RR$cR!L2g���Þs	Gg9���v�$��e)Jd��}�	p�	��400�2��bLɁ��Ji�%6D�|��y�
����n�ۧ���.{�&����k�H#b���f�q�<=~��ϐۡ-����ۇ7��ŀ� B"A*�$��(����TL
>��c��4�o�f��#�8x�6Kw��f��h`D�5����a�9|��7���!�FJc�̸��T��I!Kb�(�o�*����R��B�(B�)�9�d��H�2�aF,���s��U� ���M�ɗ�D�@�1�F#��Q�4\�<��c$Ņ`F0
Qx!��� ����MB$�P��g8f��B�s.�<��d������4��e I}��T�b��1��f�������Q�X0�1��b�,X��
Hƛ��� @`p8�`�<�k�־C���fR�8i:!NxlOV,V$a�Yd1!D2�2��
f0�4ӎ�
P`a��)�B���I0��,2nq�>"?8�]w�_OJx��)Wy��z�� �� ���f���XR�&�G����a��h珌="�'� +�F�BL�7tK��(
cl͜<=6�!L�9��ߏ�����s7�OO$��#�zj`E��x�7����c��5����+�����~�r���@���!O7�|'>9�l�$+,�OHs6pb�$%�S4b��H0�P3		��&8K�S��7�͜%�I�BB����+ �B|3ҏ���� XOS�BBģ�Ƙ�P G���Ni��8`�݌!!C5����=��0Ӈ���v@��)�������SXH�0��c��pӁ�J�F�d�ǀa�L8xz1�:����1)�4�8xz1��i�� �����at�8�$k�s1�����M�8��
a���3˲J�4�燩)��|=�#	*8�R4)���V!�XGy��i�	 @� Ab@8�B1�4���CԔ��_�s�����/ۇ�crs�vK�<���E��!7.��}c=��u����Ӈ��+X��e���i�Øa9�	p4�
�ל�y�^b�M�%�H� B�Yf�!�3aM�i��ˌ����3yK�����!��la2B�02�y��93�������Hɘq�ZX�(z�	�.Z���J�����SD������s_sc�aLe�HV� �#��\t�X�HXȄ���P��Zd)2�8x@�(�=<=1!R�\���F��<'��>�ݴf9$�B�g�x�9YO,<�4�Ěf��f�)33Os�0��3��$��C������0��!2�3 F65�̌!XX�i�)���#�!��9����4%Є6n���sc B]1%��bCf�c.d!)�g��r{�xZy���H�̐�X`K�zL�HB���y�Y��<��\!�*J�6��0�32"FFSI�%	fd�y�$gR���,A+�.����)�@��)��D�)+
�"B�.d�2 ��@���Xd����0� B0���B�c\!L�!HIX%��XS2	%����X�{�3&������\ԇsct�9�Xs�G�7^x�p�Ff��C9|�Jy�t��ﮐ$��)vnY=+LKt�����i!�N�x�F$.��a:���8i�;�SϽ�}��>N���~�Oz�a$�hF�R�)�F��
��!
&R�B,��@XZ��)��"�1i �bE�a��M����H-D�D ��@ 
�L хR	 $P� p$�#�X�"@"4`�L��eld!
a*0+��,R8	  D�DHEb�c"�k ��
�,�`�0HQ�A��  �*$jX�H�P��A�#��D���a�#�!�
�����c��cP�D$@��!p�a�\&�@āT�Ab��ha�s����bǐ�	f�,	a���1Ս�!^7$�cP��ȱa����2gS���d0ἣ$�f�)���apL�k�d�m3-�ӓssP����(�f��Y��!p�&:i��F�8A��9�Ô��¦�%1cĄ�wZ2S�8��+	M6�$bBm�����T�ܼ	M"I����dIsN(B���6$��Ï�4%�;�x�0��0�0���0�!l�o#�
�CP�Y��X`��LI9�sv��$&X���a
P�[͆ܩ���LN�z�ݹ�)�I.$c0��B7<�<�����R1!H���]�C�(B�K��~����~�P���$)�$�9�w�A���e�/�=<��=�B@��0K)�}��=$甆��(����{�f吏�0W�{"B�w�g�B�
�2��Х�����!L�0�"BBo󍙑�������{�鰦i7���Ԇ$�a����ϏaB_�f�}��R��e�2�2\�����RX��!�r^By��d
s��U���\�I�=!s�
��
��/��p���a�����q�.�#����قse�$�6ܐ     ���l ��  ���I*�. ᫌ�sg��n+�Ô�n.��VR�z��	q���{�;l�z�<ӡ����]tjLcb��\fh�N�AG
��v�ra�Z�uO\�l��S�1a��B�
�^zt��$�mb�����d�T��v㶠�Q�H�n���=�vl��%  
RCm���E�ֹ���}��m�����A��- �pf8���Q�m���*��]�i]p `�q"�L�*����u�AK����)D��i���~�-����͌�@��Cvj�R�������ga�5	 ��n�m���p�p8TQP&�;2�KR�AAKA*үUU�a�C �i�� 8��ll�5l��5�ʪ�u�l�s*�>���jr��/Z�;�`.�-� �JHh��` ���j�.  m�� 	$ kXm���*���i	�V��B��6�` $-5�&�mf���l�m�� 	&�ʑi�ln[m�-��   s�o-�Mm�I�F�n� ����[%  [_�����ڶ��`4�F�   $,3f�����ݶkm����YN�m�� p-��f�m��%����m�I� �m����T��Z `����wm�"��r�I٫`���W+��̬��UUt��ʵp!��� �m�v�`m�6b�/Z>7�|�v�v �am��lp8N��pR�@+��-�c=t�Tm� ��f�}v�}�(��I'^�@���m&��b�o[p	�Ib�Yv��$q��'�
�X�)���pKi:uv�[A���7i'�>���m�t�(��mUU��͸�;����7E��Ff n���ٴ4Pm���8l�]կױ{�e�b�     p 6���t�n��� mzn̺嵠$/Z���l m$h���lk�[{m�M��Ø��8-�+�Ԏ ɛq��N,_K�
T��*�l�2�^q�ڪ��0��(-�]��n���q��r2��mǂ^���`�{e��
v�kl�� -�sm�� ����C�I �k�f�� �,�*�J��
a%�OU�T身�vj�s�
�K�6�.�*@�v'N�,�@�39� V��uUrܘZ]�7�����٫�`*�1Hn� �[�TN˶�5�a!�� :�,�.���`�x�-��P$ �,�mi"ړ��@�m&˥bմ88HHv�-�z�Zi�bm�����m[grA��~6��Zi:� [vZ�۪��H���)hm%�� �Ԯ	�K7 &E	#K*�s�e�֥mUR�Ф�u���V��-��<��V8��0S��ny�rꆪ�㝖3t�5S˳�
Vp%@U*�����(����.�pl-7�Ab��Ŵp�P!�)��I{N��nR�'ev��!�{v�Vyj���|��lpY�.Y(�m�o��un�]�6���`܀�v�rg.�=j�d��*��k�Ci6�v[9�6ݎH[� H k�~+}� 6�����#ձev��ㇴ�[��t��m���8 V���nN��;m���  [CZ��l�I�h'm� H mZ5��4����a�d��-���!� �*ʵ�k7/A���ie�v�ON2bYw����sn�ml�-�l-�������iVU��� $m[q��sM/]��'*�ŵ��@�Z8e���^7SWU>3�m��n�q�b���-�坕�=���-c6�Ym 5�5�i $m���%�s�+��N�#������[+�|�ҝN��m�@Y`���A@[WZ�[u�v͖�]�Uuk�6Z��u/ ��S���\��Ϛ���<��UV��+�!+V�Җж�� $dM����zi3�����D�*@ ۶m�� h�|$[d�:P�1uY#]���n�i�V�#���4�n��n	%�/V�¬kk��E%t�   ��@�-T[(��8�
e�g�ŕ7�4�ř���ڀ6ٴ�ۤ�$��/Sb��K/Z�w�
f�
�Jn�#B��@@m|��Am�P � � m�@G @���  ��    �h �I�춁�P-�B��l�n�ٰ6ۤ���RY���л,�J�[ci�ɲ�u� ��t�VӁ��մ��nd 	 88�m�Ql�84P z�:Ns�3��%�5�ԪҠ0��a���0�۶�$l���ƹz8�j�9�MY�Km -�ܔ�	�ܹ�cx�\T���+���*�    �mh$ ۶ �� �` �   �	�m�   � lH  ��  �"� m��8$         	   H�    	6�vm�Ën� � ����'6Z �d����XȝiI��n�{��t�.�I.HR�nQ�eZ�=��clWT���V��#m�$ �$��V�c����oUr�I-��l M��v���D� �Y��  �I �X:'���	Z����Ɏ	'A �u�lX`-�h��-��e�ط��j���W�bu6CĀ &����\=�iU�[@�gT���-�<b��[)/UAד�`�ڑ:H�� �� �-�  ���m�@    ��6��-� �kh   � 8N�� � H m��� 6� h@   Hm   �  � ��� m��p   mp 	 l H[@%�[G-r��u�tؐp��[���� �u��6ʭ��l 8 �6�@�G���Ү-��l��S��'��!&� nN	ж�v� �[�h  m�-� Y%���� ��NYQ����
�hٮ��>/���um��k��6�ܶ�	���!�8�X-��`��IKn#�»5K����UUPWY��i����-���;�l�
����%Q�@W@-�-� $���$� [F�  H�  �` � �  � mm����-���       �x� [@-�  �jF����}��l -��	   6�m� �  8  <����9m�S�d���Pl��l6ʹ��l�,��AͶ"ZK�e��]�ȶ�jء��Cn�nͤ�m��  l�i��Ͷ    �5!<ly�t�$પ��e�ְ$  88^��p۳)��a�mp�gltY@�n � 8͒Y-;-��x�,�6q=o`)�V��R�+m�i$���m� m�ڶ  \��5�v�H H���I����� m-6���  H  Hm��6�p  �k���s`[y�����VVypf:t[J˳VtMU�[/*��: h46Hpm�i6 �`[[l �a��8 U\�l��[���vy��]B�  m  @)WE��i&�.i �`宷zYvݲ�W6��*��E��ݱm�`�Ci��@p:��m�M�:� [��}��H�K4m��# ��L�l�m���Vm��z�v@-� 6�   	:� N�BF�r�h� H  ���Wj�v(������bN�U�y�m��Z�ݥSm][u�)T �Z(u��:ۂ�:�0�m�j�*vQz����-�$X����]r�@ p�     �f�3z�q�ٶvk�W2�[�l�C2��\�*�j 0��i��]&��Hו�  ^�Խ5���NuI�-�֫��'t�L�VQU���J�ۛO*�J�@);!�k��˫j�@����;)�Ēt�کjE�k���Pj%e�Ԅ��mUP-�۲B�]�,�?����	 8Z�N���4�:]� �om�m   �H�� ��-���gH�8�kX�� 6�` ��[�  sn��z�v�I�m�6�����i0kn  6��[����� �*]n��8z�v�wea���f�p۬ג$7l۱��I6ۜ�m�v.�7nj��E���jW��B�Hr���-W[�*���5n�%Yr��.l��Hm��&� 8� ͖���V�j���EE�I�m� �Y��v���UT�V��!<�Ԅ���W(H�5�1=�%�:� &�l���#n� [N�I�m�M��F�` �9���az��60��9�n���յT=�Wn�p@iT�m��X��m��  Ž@ >�      H  m���l��` [@�:�h@'8�k��6�+��:hI��4K5h�������*P�)	���#���&� 8�#�� D�"(W�~5 �1D�D�A[�z@5@~��"�� �D8�S�#�{@C������Ȭ�� !�Q�ED��N�E�@�/©�(:b���"�	�D� T��
�� Y�;���@L8��� �M_E_H x�	�$BH@ �B1@DH�`@ BX�T�P��|!�U#��</�TT�@��C��~ �> �|!E\Q8�tEZ*x|��o��}�M��+��b!ྂ���~T:���EV�z"��~�P�z|)ǩ��qO��YJYV2�Ym���X���"!�����LP�Ȯ4LXP<���
��(
������X�! @<ɗ�T�u��wm�q��8rn|�9�&�
[>�<���I8�t˦R���u#�qpUհPNH�Y.[���ݤ�A��筇����u�F��袩�E���
��vjƲg.�d���L��%Ue4ѮS\4�ݣE����yx��sl�]��O�qUiy���l�Z�v�@��*,�'\�����=�>����y�v��q��j��D��d䝻q��c*�D�+n�9�Jy6�aqv�i^�;����	�xL�쫎ѣ�{u��gM�<��v:�u���{��[�:�.�<�wi�+݂ˬq�s�X�{BQ���r��m�^p��1������.s�Y�P�th&�cA@s0�@Uq
����˳�]����z�"��v�sf�w99󮅬�=*�>յM���r5�<-�8��vM<�>Ƭ��u�Š#{�nѹ����d�}������.D�5�c	��c�h���
[Q;6Nѻ:�]�!�r��r��k��4�.pi��vۑ�jU�8i��5*�j樰�l�Y16� ���)ck��H��]Z���h8�R����[H�Y�ۜEZtZ�M�r���v�2C���Z�6�
Cm�4�jjʂ�[F�4�4�*ͬ�H��U���F�ƍ�gcsdkqj×g\8�`��ײq��r����ʹZ�{�=��b���@��R��<l5U\�Ix+��� ��e��RR{<�n�g3n���լ+�mO5���ƪ��-�,,M���9�\�h���T��v*'��n[<κe�3/3�0r�t���c���kp�k����B܊�����Z�ۆ�S�qqy��n
K#%Y�Q�Լ�C�8>'�[r�֜��G�ٲcr�ը����6*����6�Rؚ�d�js�ӳr�.�q��qѲ*k\ͻt�زN۶��ts�t�U�X�UZ�|ʍ��z�X3�� 6A��[�j�o4�0�;��ww��{�����`�!� �D�_���x��ꢦ���'�+� � g�70���&ͳ,ͺ2%,����Ҹ�s��!���t7.8��m�ӎ�{���G��.۷]�q�m��:����wt$��&���ȹ�u�gq�:��GI����i�.v�7	�n�Y�n+u�����d�޴�e-xe6�&�q��`��u�m�:3Ӈt�Ѫ��`F��k/�1��{ur��T��7-�.�\�Q~�k������^��m��㲃����PN6�x�g�{l�8Uܦ�)+�QK�
�"r^�>w����33<Ay���;��{���,h�Y���\���Ui�էZR��D�OH�nI�z�7���^�N�4�IIJ�Y�M�I$�@�Қ+���٠z��\��ǎE䆁��z:L��7��e��ϭ��6�s�+�\s,�B�9�)	1����S��yd�2G1�d�I�H���h�3@��.���%fR���.��R���I=���H����������}����4�솁Iz9��<Y�`��&�ĖLIɠ_zS@�G/@#s4���zH���
�U��^Թ^����� \�h�)�u�ޏ�9?4c�)�^�4�Y�_l����z��*nBI�"{ d�\�����n:�������pr��,AB@<�ԍ|�~�~�6ӦC@j9z��wZ���b�Ϯ�#�G�_l����z]���W�bG|>�<q���C@���Н�}���Lb��c#��Tpn�r��ҚS��c�NAdY��Dܽ�qh�C@j9z\[FȚ��I���Z��h�W�U�^���]��O�d��;;��T
M��թvwVܼga�c[�\x�JUk�Ә�p2&�Z��h�W�U�^���Z�Ճ�iaX)�r�q1C���	�u�/�#@��oFڊ)#Ic�)�WuzW�h�)�r�^��tM\x��*���[�@�2Q����U|��{��*�:=�Qܽ�3�O��J�LY&1�F�@��M���
���:��@3��0��\�FM��j�t�����o8ܩ,K�؝6IY��s�n\�����CdqFFG!�}~z]��_U�_l����t1�ȅ�Ȥz]��_U�_l����{;�LjD�RF�#�@�@�e4W��*�^���{Ӭ`c���/D�OY�*mހ����b4m��6�o��JC@�[^��鉉v���$�ƀ�b4�110*��>�a|�2R�fi[!��f�u���.�:�Gd�.���=Hu)��M��+��!�K�l=�ʆ���J���lpP�c=z�!� ��4���n��&��������=�=k1���'	c�=q:7cq�ʍ�΋�d�@���v-V�F3!�:PɃ���lh[�%fb4s�u4']srgNL�=�jFoj�Zg���D��5����ϝ��0Sp�b�m5��"n�㷫�&���q��]P]�39�Si�	������;
o̓���^�ܛZ��9I/@��Z�%K#1Ȝzu����/�S@��@����Zĭm`I�q�C@�&ց�$�&�������q$�Q���h+k�/>�@�}V�}�����c�j'2dR=u��ҭ|�Ԓ��3� ��5��ݸ�:-ˠ��vh�K�7XsK���I:N�C���Vq�Ri���H�G���~Z��9I/@��Z�u<m��`8R-�e7���ٙvc���UUV�U�f�j�/@�r-�qh[V5�`��)Ĥ4���U�wt��}���S�m(��B"�2�/A�M5�ր��h��?RU��D�i(��"O�Šw���/�S@�^�@����;�(��I.����h蓠⋌�A�D�2�Tc���m�$�"B�7�7�"�/�S@�G/@��z]%��6��W�Fa��hR�z�bf"&*��:�sw�_l�����MƔs4��-���I>���ɕ�}IQEg;���mz.�pq�#SN-�r��C@�^�ȴ*�uwP p2!H��S@�^�@��Z/z� �9+aA�<�	��Ζ3]Pj���v#�݃i��<j&$4�f�)�t0liH�%!�x�W�^v���^�z�hڞkiLCr(�$R=W%z�j���h<f��|�눈������IL�	I�Ȥzs�-���<^��
�נw� ]E�G�Ǆb�4�C@�r^���}�|���1tPi�o��������,�4͘fy����W�8�i��K�.X�ͷ���}�u2��8z���]3�:V6��]��6���	HjG���CR�vx2:.Sm��+~zs���<Vנr�cmc�$��D����o���115C��:�w�*�W�~���Vb����p�/�S@�[^�WuzwJh�^=�i�#X����^�r��h�C@��hڻ���Q�Iz]��gw���w��@�{k�~^�Z��UO��L��h%n��)_]�\ާzދb��=����ܼ�ǒ��m�J�l5�*6�=9F�L�Wk�6��ŹK89��6�c�l�5c�*���t/<dg:P�r��v1v�nb��:9iNN��R�:w�2���˵���eers���/m���p�����Uy�4ka���n��[����s:��]p�WF��T�m����~{�{��޸��5M���zT�wg{[�c���J�8; ���Ƹۈ�7Q��2�(b�'�8���Z��h�mz��h�HQ��"�/�S@��;qh�C@�%J�� �B9�ֽ�����u��@����r�n$�ӏ@������	�!��'%�71Yv��3.�*�2�������|����_�z��h{P;	�cm<��Ȇ�gAv�h��͚�
Z���d��̑M�\�c�����e4Z�Ϫ��g�:��}�|��H����Q`���y~�s��� |�w��^Hu����h֦����$dr)��Gn-��h�C@�r^����i
cM��q��Jh�)�x�נU�^���aΤ!�R~'�4	�!�J�/@��z7�������&��;;�ֻon�Eu��K6����ч�k!ӱ��m�o3����4'%�7/@����<Ʈ�$����q�wW�{�)�_l����^��ޱ��0�71L�߾��I;�w��י� ��
�O@N��,�D�b��[;U�~�0!+$n ����b���qS �}'Ř� �'����� �� �z	\913\��g}�4�@�Iށ���资�E�fAww���|��ԛ�Wr���ߍ���rhk�,I�@�rW�8v���rX�|��bff��	��̮�C��n yʗOGOJ��kt�(z�0�lZ'�sO����O�Ț�6,��?������C@�2������F�iD8�{�7����͟��/����Wuz�՜�hB�9�gֳt�hNK�"n^��ͭ�_�dS#s�nC@�u�@���rI��w�$����1� 7����R���$ړ�cN=��3�6�	�!�ysX��`�����Qзn��{)H���2��=p��b���M�͘��bm�"Ǒ�L��MH�=빠_m��=]k�/>�@�g�ԑ��ra��3+@�&ց��zv��9ɵ�_ml��(�&�bĜ�������W~Zw]��n��jkP���j,n=����/��h+k�;�7[H�X�DŠw>�@�۹�x��@�����ˍ��<MLS��\�6Xѳk+��+��i�Zb��F� l��M�9�\�Z�+���:��k/f�eC�Τ�|8q�pn�ݧ��`�;1l8${I��Fͷ=���\dc�vM�e�W����|����1��+��� ��ݠOVݭ�mK�N���J@nG/)f���cv�^��e� v��7Hh��������wm�t����1hͳl�����w���[��M���i3�%2�-&�8�ګ��ar��
��M�նj��9i�[&d��q���ۚ���Ϫ�9wW�{B��G�&90�������Š4ܽt�hcSlJ��/-9�&��*�@��^�}�����^��I�JAI��=�uzeS��>���
����:9ee�%�G�67�}�����
���z٠uꆍr"5cl��b�<gmY�b.��H�pi�8�.r�l�gzݦZT�a�rr^�r����ꪯ ��������ɍ���H��/>�_Ԑ;�4	�!�rr^���H�e��Pk� n- ���@��M��f&�����n������+(ˢ�ʼY��G&ց��zv��97/@�����bq) ۙ�x�נ^�U�}]���[����� xfڎyw�䔗ea��ke����Di)l��r;^J��Hc��-ە�ͷ���������n���^��쯯��9AI�)�uw�_m��<]k�/>�@�ggY��N-�n��y~�s���qDQ�[�{�N@��Z{ս�I�6F�$�h.��G��y�Zp��Y��Kj7#�@������ٟ�2ۿw����'���s�,ll��o���%\��U�-ܻ�-�R�9������@����i����R�-��� i���lll~����Ȁؠ� � �������lll}�߿g �`�`�`��������lll}�����mٗeɺd�� �`�`�`�߻�Â�A�A�A�A�;��pA�666>��?N>A������� �`�`�`������6fK�f˻�34���lll}����|�������ӂ�A�A�A�A������ � � � �������lll}�;y���]�ni�fnpA�666>��?N>A������� �`�`�`�߻�Â�A�A�P��A��߳��A�A�A�A�}��ə�3t˹�nnl���lll~�y�pA�666=���8 �s��g �`�`�`������� � � � �~���d���i�f2�B��r۫)Ӝ��%͌�n���-�0t�qU��5^ҳ���͞>�����xpA�666>���x �o^>A���߻�ӂ�A�A�A�A�����v��K�nZ[�pA�666>���^>A������ׂ�A�A�A�A�������lll{�xpA��0r9���<��6��M۹�wo �`�`�`������� � � � ��y�pA�666=���8 �~�߯ �`�`�`������30ܚL������� � � � ��y�pA�666=���8 �~�߯ �`�`��������x ����2����ݗ&�vpA�666=���8 �~�߯ �`�`�`������� � � � ��y�pA�6668(����02n�i�^�M
Ֆ�'W�e���
���)u���t\�vyHd�k1��+>[͒]˲T뭞7X�ӻ]v�e����p�d޺��Y����X�f�\v���c�t緗�&��

���m�At�ݓm�J��6�gl��=�v�f�,s���p�e�r���x�L�-�Z�CUu)�v4n��i/y�{&G9гCʤ�`"a�~�rDɒsg��r�y���7nk�Z��=����dijj���JORm�0�V��d�͙��D`�`�`�`�������A�A�A�A�������lll~���8 ����|����������3wmٚi��x �o^>A�����Â�A�A�A�A������ � � � ����x ��߿33.nܙ��n]��� � � � ��y�pA�666=���8 �"b&�����ӭ�iց�p�/3���9&h~/_���ߖ���M��>�h���F���bNf��Šz<�����ͭu[�y@�:�nͽ��$v�bγvwge�wP��f�N�KO��8�Rc�����C@�\�@|�ց��zo.Ԣ�˷i&ͷn��߳��� "�	2g�L~���Xo��>�n�˱�ㆫ��Ll��-��M�ֽ?Չ{��W��@��!#po0�99/@�y�ȴ�!�s�"s�cƜz��4y�Z{Қ��z���+��#H��໳!�9��P�L+��fMm״��CD���%�6��G�<�8hfgY���/Y�z����~��@�gS�q��K���;��o�&f&=vu?z������������D��I��<]k�?.�i��$DA137�_*�?r[u+�"dM��E�ǠyzS@�U�wܶ4}m��9,��W9pa�%�0����ͭ�Iz��|�}�����\�nc�P�<jל[��٧�$1&�ua+gus�n��|��g�(���?8������mz��4��hԣ�"�I���m{�G�c4�:�;�[��{Q�fY�ew��|�3@�U��"}3m?nh�������u$ڎ7yp�s34�'Z��4Ԓ��1�LdDQ�@�(P?x*�)���<������)0pO�4��;޻��z&{=�_�w�x�;��h�����T)�zR�Ӵu��Dp��:���l;\�]��=OtG3Q{���������n���۽�U�wZU舏DD�`��ƀ����PO�4c�F�q�^�߿g�Ą���'��}I+�TrYWN
����ʜ���4���;��h�"j��w�{��/Qì�I�#jc�-�L�.Z���z�؍�7Zn�-�\\^E\x]�Ԓ��LG�k? ��Z}؍"�%L�H���@�) �I"��� ��p�S8 z�
��BF2�(��HH25م>d%�\eP��pĹ3.e�`�����A�Q��B�B%
Z��+
BI!,,��j@�F��$�)�4�W!o�@"$�s��b��`T�F2�ZE��H�$�	!!�S�C�#F%H�%!E��āhB��(J�����
�X���*V��#�D��HR�I
x]�BSR,e�B����J�#
++K	(�(Ɛ(KF��a!d	X0"ڿ!0�PXA�*�b$H�, �P#X"�BR!A���,HA#RT
T�+)J��"J�IP%bD�"@�e�m*B1bA�	$	 �$Yĉ"@�H�$"B$H�� �1��ܼ���ڪ��"�u�����v�pP��[�)�5�i��;AE�����v�6��nո�˹y�F��G��g��F۬�!�Vճ�O��>7)IF�]��(�8��SĨ��W0�D�xmu6�'rv���B�=#��[aۀ��Nd_]��9��T�PsN�����7*�g�c����K08�\-���ƴpO-��,�J��룅v����[���U���7��*�^ȝ�@lOLƶv����NL�6��<�;|����n�ԫBp��S��<IM'F_m�Bԭ�N��Y�Z q��{!k�����r�+k��;�gu᧟c3(��JR�^�ɓT��As]��r���NՁ�������"�ؔ����-$��3����v�{�n98ͮ��`�H��壛�t7"m]�[;�(;�t]b5pJ�vg3�;��<�G�D��@ZM�Xq�`��� ���,�\�{��mk�z����܊�nڏa�/C��Cj݋]����H�d�OR��[Fٶ&�M�\ U@)-lF��F�ʻlZdӯ��PK$Lg�U��E��cJJ\�B�9�Ƕ��I�2s�gUgS-�6��T�����P6�Ԫ��|��>*��ƶڶ���I�\�С�*�$�-�%qm�uװ���6�͓�R@�Κ����>���mÖA�ø�5m��9���z:��K�5@p2�=��u,L3��l�E�;���sŀۮ��ʻ3�t�ñK���u��s2���2��f��N��k�d�T�m�|�SV���dV6���EsUVݴ�mb��n�³� ��B��i� *ѥ��I�i��ٴ�-�rij�kjAn$��.�'<ѱ���Qs���n�j�	vTņ��4m�s�&m.&�
�0&�]+3��T��I�)������m-��܉�����u.^��������R�:�Ӓ㮒s�j���ͳ*�K�m*�!5x.������W�P�#��Hj������p*�;5��i�6e���wr��=�n�)
^tn�ݐ�����~|y�cs�����R͹�v�N�A���Gs���9x�7+;y�'k5�ΰu�c�ђ�-qm�ч�=�av��)V���z�ꓷn�XX���rmf�2 ���8��.�h����%�=N���l���=�+LΓpUqu�ڴK)�y�Ч�tF�CED�K;,��M�;����ww�Q�dF4������*a�HZ��g]�k��o���4<a��Mi�����M��&�"E��y|y�@��&Pu&�@���1��r8�8�{�տ�����cO<h
��z�|�\D�Q�G+�eE�W�e�eh�3@��+�ޙ����V���ՠw�J�ȣ#.3/���A�Mu��@��u�}\��9�\��j	�&�r(�R=�����Zn� �c4����݁t,̼�{b���;f|X��۫]<&A��r��<���T�{���>p��O��?6ߧ����<�������s��qU���W	��f9���'����؍@	e�k�=�ՠz�נ[R��cƜɏ/��@����Z ܙ�>y�r!bpn0�	�8�+�\���b4=3]m��$��.��2�G6�Z.���Jh�k�<�����v��8��Iǌ#���͗�p3��ܚ�Z1ۇ��E�L��)���]�ȉ#�;ޔ�=Vנy_U�ffg�-�|h��a$f50�A�R��z�|�@�iV��v#\�LDU5N�J!�$j)������է��fff.})�r���蚬m���.B���t��z��:�+�诒܀w,u�I�j!�Ǡ{������wJh�k�.*�n�G$k$��M��b�u+�9��f�9�uݷ�3]�gs��T�	��0�2G�4Vנy_U�r����M�ȕBLML"��N=�����h�Jh��@��DO#RGF�Z�ՠw�)�Umz��Z�=�)�O�v����4���z[�C��Q_W��������]hط̲.����0�$�@s1�����u�w݈����ߠ��K:��T�e���ځN�+\*��r�7(�0$qn�$�ci�i�G�y_U�Z�Z{ҚVנ{�J�k�ő~�E!�Uz��1"������<�)�{�`�)dRI�w�)�Uz��Қ׬�-�)`��HG�4W��<�)�z���M�q��eAquyz�؍��Rm��,f�����?~�/��>֑7m�E����:�u+���;6��8�l��s�u�LrD�{=V�+�:�!�{a�V�����Sv��qr�N�we�t�pix��܎�ێ�&�&-N�f�J���T@�끀�öW.��E[�XXW��fd&����N�E{�[hxsb�B�6�k�-q���k���N��٧�x��+,�o�{��wY�&��$zl\�S�v�,�뫶��5ቷa��s���u��e:G-e�0� ���@��u$��0A11��߬��=Yկ��L"x,�r=��Ms3C���5��$�@��-��?%0q�X���U��^��*����M��^����i�F����!�E$���hI/@��Z\q`%�Ԏ- �٠}����x��z��Z�g&�F�I�e�:��&y���,�IN�^�]\�t�Y0+V�8�H"�M��M�k�<�����ڒ�`��28K�4������DDG�>v�h��@��F�b&#�7c���f]�afTw��w�ޭ �%�8���3@T�� 㭉<NE$q6�Zg���/���@m����D��b���V���x2#iD�Y1I&��Қ���+�h�נy�PѮDdq�by		3{V.k�e�LE�:��Wt]:2\��~�|�}�s �j9�p�_}��<�ՠw;W߿g�-��@���RQ��6�M����}舻�z��x�>����Dв��	D��E�w;V�����@��o{����{y$�{��E"�y��;�S@=���C�114�?Ѡ6��wE�ff'0�f�y�@�ڴ}v��w4=����B#�@�h��nPĹ	���]�ӻ]1/^;k(��^�3x�A]k5�crh�V��ՠ[n�{�@==챡�H㉤��=^��m��}�h�V���#՝Y�J<x�$�Z�}��{�@�ڴW�����F���N51�����^�;��o$���v�O�Z�w���j�RQ����nG�k�h�؍��Ɓ��+���1m�.�2����j��Ny)vx���ۗX���&����-�:�H�"hX���A��^��@mͭ�9z�ȴ���U��efb�u��+@mͭ�9z�ȴ�o}��ww��O���k~Ӯ���蘭����?+J�����.Oc@I=����&q�Wj�:�����s@�z� �XІ�rD�qh��h����Tӽ�@ș��߿w��K9�2L�FF���\�.���9B^$���bN�����8���A�i�Yۑ��[6�Ϯ�;V�Jj����m���K{=��l;���O]�/L5��NeB�la�[(�$�J.@�q�GY��۴���}�k�llC�l����"s79�n\Y�nH�c��=��K4��o.���vC���n{bv�����1��I$h� �\j�k��������sZ�<<�km!�׵`��q��!S����ֳH��JDӋ�����9^�@�W߼A~w�^>�F�9�5ɏ̍�r�sT|��D��~�z����<�[�JE�24ۊG�y]�@��Zf%m�s@��zwFб���+2�
���sI=f��{Ԓ�Dg�������
����x'2FӃ�hܶ43?[n���@��W�zbb#�bϳ�>��7qE�Ls���0���j�y��=�{m�;u��`ۊe�k1��9	$s=�����<�ՠw���3��-�nh�|��I�ő�ɠy]�bDO�_ɹ��~���/o�Z�籠�Y�fg䂗���j��qh�u�wr���蘋�^~��~�h�>�\#M�x�$�Zw]��z��A�E.��@\7���wYYY��.Y�9���u���hܶ7m�����p)Nƞ�ڽ���;[<�k`�� =n��h�؛Iz��]��~�o�������2�3�;n���V���c�1311����?f��˺*.�U�w�U�-���sk@=$���[��#�*���!���-�nh��y4�N�A�T#�$�"��RH�BYHĉo�O��F$���d%#k���'E��Z�2B�MB1�#��B2FDHBi�D�ɠ�B	�T�`�$�!	B|u>tRXB18�)_�SF#�y��H��F,�B	N "tCU"��^"����q�!�8��.�1;$L���+���x�.��Yu�Efw���y*�m���@��M����:5@DɐȰlNM�@r��~$�4�Q�o4�W��^�P�ݍ/���1�1�N�@8�^�X�3����ﾕ+gU�*ܿ��M��h	'���X��Xw�ޭ�_���L&B4G���s@<����Z/z��"�������S&L�̍ ����iV���U�ހ�{[[ׂ! �mȤ��ڴ\�������?����ho.�wW3$p�7"�9{���w4��hWj�/���"S#��	'�d�ɻh����soC��n��7'[��I������I4��ԏ�-�nh�٠y]�@�}V�o(ۨ�(�ML�G3@<�f��r-�qh���z��2lNM��ZwJh�w4�l�9u�D��!X�qh+n�h߷4�l�<�ՠx�ޱ�&	���@�빠[f��v�$�ﷳ�J���j�JU(+U"P�P{�aO|03r���цԑ�z���V�h�L]BMs�	�yz'�
�*�vs�bS�b�J���J��v΍�=�78�t�MҒ�\�+�K��4Lnٶ�J�Vcݽ�@Q&��^�8�iF�gg�+\��O�ɰ o�aýZ�L�+���˹���I��"�c1�<Ƨ��7h�@�,\6��Y�e����mu�s ב��z�'K�V�۝���;��m�g��s3q�u鑸��W�_��}3vz�;vRY� ?������Zo!�6�ց�Xb&B���hWj�-�M���[�h�Cx�dRD̃r-ޔ�;��h�f��v� �Ҵ�8
B9�9���s@:���ڴ���-�j��8��+��h�f��r-�qh������~��]EV�M�.�.�jBݎˡ�W+$u����:ﾩeM�Ν��ҦY,"Ȗ�ʼ��|��:���ܶ=�����V�$j,�G�'�����X��,mͭ �4K�hU�e�V5 �(�Zw]� ��4+�h�S@�Kt�����bRf�ĺK�=.E�w[0?&��h����QJ"nH�$�@�V�y�Zw]� ��4=�H�Ԙ�#�m=[��ڂ<�qn#Z��y+t�s���Z����|Q&��E2D�7"���=���_m�g�=����x���`�FH�6�znmh�3@���r��U$~�ToߦI��D㙠w�M��Zld�E�31I�L~ۤ����h��X�R%A&���<�ՠr�@�屠�b*�m怫�ʻ�2�32�*�+@��W�8�����>m��ZK@������1$�i�F�L�r9�;s�qg::��ء4WGgn1�r&�tSsS$#�5	�4��;��ym��ڜL��V�h��̻2Ƞ̂2*�#@?$�\DU;n����D~�I=������D�8�q�&��v���i����� ��h�m��)�7�nE�u��w]� �l�����^�uh�g2�FҐ��Cp�;��h�o?��@\�����MY��h,lڛq&���Dj�u��X��9vݞ��?W-����ή\��I'�7��iV��үL�~�I=��cǉ)���i94+�o�bE�ߖ�m�s@:����H����D$��J�h���@mͭ q��=.E�yg�����☣R-�+o�f�_�y�~V�h9�O�pޑ�q�E��U��,�=����	�u�wwxrI�`%=C��Ap� ~��=�~Z^JKfk��T��m��Ō���C�L�l���	�b�.�W[���2jr�;EQvG�Ɲ��۵�MS�V�:S���2��ls�7:5��t�iu6�6��mi�b�ɤ՜�{@�_k�5 �wR��ų/S;�{3Ֆc`��W��x�[y��+xv�m�>I����{4z��D���rv@���4	]�bY�n���ww�L��K1!��cNu[E<�;�Ŵf�Ρ�S۵k�`8�I���Z�b�$i�#��p������ۛZ 䙠6��H��,˸ʻ��2��*�3T$�ƀ6�hWj߳3x���X�j!�1��[~��m��ڴ�S@��b�3������q11T�y�|��,F��b}36��Ѡ/=XVfe����rhWj�/;V���s@/[4
��0��'���C��ܓ�ʅ��.^�8��+�Ɏxt�|�^/CO�ww���G:FJ2�+2� շZIlh��L�A�������FE7Ě�h���DL�D��
ĳ@T�^���V�����c���*���2*�#@7��v�������(�Q��̼/34�|��$�@�屠�f��ѱ!XH���G"�*�F���?{$�_����$�]�w�$��7_2/��S]�6���v�2n�7�-=�'bb��m�/���i�lUR�p��j4��Y~�I&��$��3�I.���RIKn�<I*�!e����2I���^[3�I.���RI7�/y$�spԒ^����qȔ�����Ē��[Ԓ]ӻ|��P�76������o��~�<�ޏ�ݬ���e� ~�߿O����jI%�&{�/���}V�?~�Ԓ]t���FLDnI����Ē]�a�$��l��K��Ԓ\���I.��m�"���8��j���wm�n���q9]���N^��}��/����v끭� ������K��ԒO���I$��5$��G�%�(�S%_������?�ʇן�/y$���I$�9��I91X���$��!$��I.��<�$�u�j_~m���<�$���oRI/=1s�䈍��9<I}����!�$�}~�x�^�kz��_GD���D�s��Ǟ[os䅗42BD)�H�5$����x�_߿������]�I/�����I$��5$���?���J������s�P����ݬv�%+����=�����s�r�g���Ē�.�$����I77�UUz�$����%�w�$6��	6��z�K��U���1��M�pڪ����~�UU��W{���*�߿Q��uƖ�3�� }���RI//Y��?fco����$�}~~x�K���(D�d��r�Iyz�<I/[��I%��_�$����7o�CRI_���q�ٍ��G�y�Izݭ�H\����,��,���'&0�$�	���!b�)E�b0b���@���#<q�{e%�R�0$��#(Q�#$i(��������DO��# �
(��@X���a�`DHD"F@ ,H,XF@#) E�B@ ��bń`0c"�b��!֥� �0#!�[5HJ���98���'jъH��f�Б$!I� FI��I;�~g�� [\^�_gZUw[��F�F�jv�og��2s�_��,T�բjt�:����Nm5��{9���؈�V��֠��m��ڬ#BKd��IN8��+`�8�3L��R�`p��Rw\�p�ְ&p�<
�<��!j1D��v�=�7J�$˺�b��	��Y\�m��盐�V���9��f�رh���,��UR���j\�s���[X�Iӭr%��u�A�8�wB:�r��/�+su�c\�b�x����	�'�s���b�v�Es�]`�Mg��u�ݝ��8����@�3�){W\E8|KͲ�էH\n;b�ޘ�cl*%�rPGP��Tkd�[�V9\�v�U`�seZ�(mpͬg�d3�b�c��L;z�Ls�=gyu	C���,� f��y�uGan��۷�=�E�gxH�Qp�N�R��c\��K:T�-��ۏ5�
�(*�� �Cc'sc��v���\90*KT9���s�؝۳dn˜�ƴq�RKs��ڠ��&؛`�I�lI��gYヷWEOŧ5�ګ�ĽNή ��fɮ[����,����{nͬ�n�U$Ģ@x`Cg������  ԩF�[J�kr� �@�m���Vv\�O0�c�H烧��dݍq��m�T��t�� �77Y����*ԻN���
VM��e��-�ڛVS��R�R���]�]��zw�݇Xk�0�N�v���ĕ�NzX��e��� � ��=5I�Km�2L	�r�ͪ�+��3*��Eb�A�nU���*��q���r�VܫƼ�*��ar�
�n'D����e���l�&F6�XVu�sJ�/#�rg�c[n��F葧�h�� \����CkO.�оβ��1Ú��CQEP	����B��OU�������7)�7`%h5(��]�9�8:�����<�#�*n�õ2�֭��Ҫ��*�:��ۦɘ�ٛ'� 5D袿� �B���W�9��C����#�ݗ1D6�֔�CT��l��P�SN ���q�:�SV�M�N�!2����p��6��et�^������:b&:2B>�$Cf�vЇ,�ؑKtس�w�E-n�)]v-��t[�h�N�]����v���B��;s0R����T@�m���6Έ8F]i�<����w>�omI��`[����%�`+o����6�F���VVc�:��B7h쩓E�ͥ�i����/P?]���Ջ[nFق�!$���_�z�� �r�?�:���>���c*�⊪̌�̽ �4���r�/@����TݞE�9��eFY���������>��zwJh��4)خ��9$�$�ʼ�]|��	'��|�h�h�ԉ4��&�4�zwJht��rf�ˤ��'H���V�v�<׍�rR�����a �q]���]��
�4�-�ݑ� "y$ěp��呂x���Iz7��łH��[���O>�w�<XE�)�[��z%���K7�Tsc��˼l��I#�94]��@��SO�ﾚ���u�1km̍�
rG�sy �4�L�9t��y��*V��̬��f�yɚ.��y�Ze����ɍ�� �$U9F�Ůq%�`���̐л����k���f�{^��D9��h�mz�ҟ߳�w�M�\_n#�H�I�����W�ff��ƀw7�W�^��}j>�i�Fx�q���nh��4���'�m���I;{�s�O)߻��<�bnI����ڴW����s@</P�<4�cĜ��h�K�:9���f�9�P���!ṅO�n�Վ���=��c�pH.��ތݬ�g��T��	:ʎ�zi����^���4�L��/@rEkn��/��D����S@=�٠U�@�{k��ٙ���8G�傍�B� ��<��Y������w�5iց}c�)Y#RM ��4^��$���o$��<Aw�@��pG�D}�����I����3e����neW��5�^���������{��������W�,ge����B��g�6�J��1�\ ��B�.���:���`i��<m8����@=�f�_m�/mz�=�$�BJ'$ěp�oY�~̈���柦*�sw�5iր~ ̎%�x��@/�����?�������4m+��q`�2'�@k��7�Z}H���#�]���}HKĽ���9ı,O{�ܴ�&:Y�ۛ��O"X�%��n�T�Kı/�����%�bX�ﻻ�,K��=�s��Kı ��⋻}�����瓶&�mZ�Uͳ�uJ܆{@]��,�"v]�����wl����tŒ_5�y^:I��Ny���)�[��3˻n�u����u�\���(獪�]��J, �M���5qsԚ�-�m�&�`�S;����'ɬ�hq�I4�]g�^w;w�JdA���M%;WR9��d��b���k0�.7%�E˗��D6�x��:���-�-�g����c`댉�[vѹQ'�\�&Ijr[�h�6�]̶ٺ�ݕ<�bX�'߻��'�,KĿw��9ı,O���8��2%�bw��ҧ"X�%����L�����n����'�,KĿw��9�9"X�Ͽ~�'�,K��뿥ND�,K���q<��.TȖ'������
-ow��7���{����8�D�,K���Ȗ4X�'�����H���݊H$�ϧ��YrYp�e�NA$��N���*r%�bX�~��8�D�,K�����Kı>�{��yı,}�wwf�l���-�͕9ı,O{�|�yı,?
�����Ȗ%�bw>��8�D�,K���Ȗ%�b_~���ۻ9:��E�F|����/V�cm�'0��!��s��N��T���4��ͷ ��w���oq����v'"X�%��{��Ȗ%�b}۽�?�� /�6%�bw���q<�bX����ܙn��f��ݻ��,K��=�s��>�Zș����Ȗ%�b_}�w��Kı/���ND��2%��߿\���d2�nn�q<�bX�']�*r%�bX��{��yı,K�{��,K��=�s��Kİl��-�2�n����"X�~ dL��߷��Kı/~݉Ȗ%�b{�����%�bX�w���,K���gf��M�����yı,K�{��,K��G�����{ı,N��͑9ı,K���<�bX�%��^��3n՝f�gGHuv/H��۝.(����w�������sv䩬���feZ����7�ı>Ͽ~�'�,K����Ȝ�bX�%���x�D�,K�����Kı<�����̒i�l�̹���%�bX�w���,Kľ���Ȗ%�b_��؜�bX�'��{�O"���2%�N��۶m������n��,KĿ}���<�bX�%��݉Ȗ?�Lx��<��9�~��O"X�%����9ı,K���M�ɲ���-��'�,KĿw��9ı,Os��8�D�,K���Ȗ%�b_}�w��Kİ~���wd�6����؜�bX�'��{�O"X�%����Ȗ%�b_}�w��Kı/{�؜�bX�'�}�e�n�lF��i��*���]�NJc�E�L��ҵ=�2j��<�Ħ�u�8��5?=ߛ�o%����Ȗ%�b_}�w��Kı/{�؜�bX�'��{�O"X�%�g�ϳ��nm�f�ʜ�bX�%���x�C�� ��ؖ%�߷br%�bX�g߿gȖ%�bvg{q9��L�b~�v���ݥ�����O"X�%�~���,K��=�s��Kı;3����bX�%���~{�7���{���>�O�0�%D�Q9ı,Os��8�D�,K���"X�%�}���'�,K�)��H��wv'"X�%���t�70�����˛�O"X�%�g~��r%�bX��{��yı,K߻��,K��=�s��Kı;��^��4��e��;�g�����H�6"{F�ݬ�˻�m\���`�ڛs:���狀�u�b_}�w��Kİo~�jr%�bX���q<�bX�'r����Kı/��76eܓ6e4�wx�D�,K���"X�%��{��Ȗ%�bvgݸ��bX�%���x�D�(��;�n���|�Wa6�Ίow��2X�'������%�bX����'"X� �Dȗ�~�'�,K���~�ND�,K�����5�$�6����yı,N�s��"X�%�}���'�,K���sS�,K� L������yı,;,�~��p�.�7vT�Kı/�����%�bX7��jr%�bX�g��q<�bX�'{��S�,K��D�
3��ɇrɾH�v��E6CJ�9�-��ۭ��ֱ�V�h�R��=�\МOmh��lY������x
'�t�6���i�=/K��'K�������	�m<�p
�v$v�B��ZE-�GF�v譭Ȼ�q�6�ZP�����S+҉�x�F7@�.�Y��p{#E[��j��O���)eL�h:G���6�6&wf���\����޾w���hk
ڡ9���g-Ξvcv�X�@jq+�K�m�{V��Vp'[e�\�ۻ�'�,K�����Ȗ%�b}�����%�bX���r�"X�%�}���'�,K���s'd0ə��ۻ�����bX�'��{�O!�c�2%��?g�Ȗ%�b_�w��<�bX��{���bX�'���M͘a4Ͷnf\��yı,N�s�S�,Kľ���Ȗ%�`�����Kı=�{��yı,{���m�rnil�ܩȖ%�b_}�w��Kİo~�jr%�bX���q<�bX�'s��T�Kı/��76e�m�0����yı,߻���bX�'��{�O"X�%���;�9ı,K���<�bX�'ӽ�,���]�v�q�<�6a��>s���j��{�����]��5�uI8��)�9����oq����{��Ȗ%�bw>��ND�,K��{�O"X�%�{�sS�,K����e��݆a����7w8�D�,K��w*rLQ+�2%�}���'�,K�����Ȗ%�b{�����%�bX�϶�3��ۅ�wr��ND�,K��{�O"X�%�{�sS�,K��=�s��Kı;�wr'"X�%��gז��w7p��ݻ���%�bX7�w59ı,O���8�D�,K��w"r%�bX�����y��{���>�wݔ^.j*Y��7�ı,O���8�D�,K�!���<�bX�%��oȖ%�`�����Kı?g���I�f���ٻ��Z�쭆���hq�c:����պjGU��ۮ`ң?���{��7�����9ı,K�~��<�bX�s��ND�,K����'�,K�����Y�sKwwH��bX�%��wx�C�V9"X������Kı;�~���{"X�'���9ı,K����-�n���sw��Kı/o��ND�,K����'�,h��>�8'����Ut>5PJz\���[-�9���M�3���Tbd$()� A R&��\#9
$(B�%<n�a����D�}~@� �: �PG��OU��X�Ԣ"!ON�'"w�g��bX�%�wx�D�,K����m�-ٹfn��ݩȖ%��������gȖ%�b~��*r%�bX�����yı,K߳�S�,K�����<�[vL���sss��Kı;��mND�,K��@������>�bX�%����S�,K��=�s��Kı��޲/��3@U�O=sI�]�q����:"ұq�1���^i��
�K.I꺭�ܻ�S�,Kľ���Ȗ%�b^��ڜ�bX�'��{��=��,K�w?eND�,K�}{r��k���f����'�,KĽ�;�9ı,O���8�D�,K��w*r%�bX�����y��L�b}�n����v��]�wv�"X�%������yı,K߳�S�,Kľ���Ȗ%�b^��ڜ�bX�'���M͙�M3m���78�D�,�"�������"X�%�~�����%�bX��wv'"X�T�U�� `�bw~�s��Kİi߻����̖niK��S�,Kľ���'�,KĽ���9ı,O���8�D�,K�����Kı<��nY�ݰ��%�͍v�\ݟ�y� rI����˸�q�sIt�s���Y�8n�K7e�����=�bX�%��۱9ı,O���8�D�,K�����Kı/��w��Kĳ���}~���٫5ow��7���'��{�O!�Dc�2%�_߷�,KĿ~��x�D�,K��݉Ȗ%�bw���Y�i�]ܷw78�D�,K����Ȗ%�b_{��Ȗ?�B"_߿n��Kı;���8Gؙİ{����l��3m4����Ȗ%�$��~��x�D�,K���؜�bX�'��{�O"X��+2&~�����bX�'���忶d&�6��ۛ�O"X�%�{�wbr%�bXG��߳��Kı/��ۉȖ%�b_{��Ȗ%�bUg�C��=I�n�ܕtU��bѝ�_g�<]
#��<Z�t�3��˄����q��1��䗠���.և�+�ʳ�qz�׋����t��B��+m�Z��*Jaz3�X�,�Tl��L�r9�loP�[.��ɲʀ�f�J��ȼf�.F��qSAU��[��	�M�;����O;f�4W�s=�'����]qN�"Y��{�������|�k�̑�W!�eg[e�Pr��7n���SRK��C�ڰ��3���l��p�H������o'������%�bX����'"X�%�}�{��g�2%�b_�~݉Ȗ%�b}�~9�f�a&����˛�O"X�%�~���r%�bX������%�bX����ND�,K����'�? �n&İi��?�Mɶ�M�)n��r%�bX���oȖ%�b_��ڜ�c����~�'�,KĽ��n'"X�%�|��黹i�.�-��'�,K?�D����S�,K��>��8�D�,K�����Kı/����yı,^��3�ff�7L��e�ڜ�bX�'��{�O"X�%��H�~݉�Kı/�w��<�bX�%��ݩȖ%�bw���6�i�����p�anwc���p&�J�B�Z�kh��磵U%	�#p搦~{�"X�%�~�;�9ı,K�wx�D�,K�����I�L�bX��߿gȖ%�`���/��)6f����Kı/�}��yz�$ z��PJ^��șĻ�wjr%�bX�g~�q<�bX�%��ݩȖ%�bw=�闻,��M���ww��Kı/~��ND�,K����'�,KĽ�;�9ı,K��wx�D�.�����af��H�{�oq���@Ȟ�~�'�,KĿ����"X�%�}���Ȗ%�b^��ڜ�bX�'ݟ����m����˛�O"X�%�{�wjr%�bX��~��<�bX�%��ݩȖ%�by�����%�bX�wK����i�$�p�nKi6o4�M��� @7K�͞�c�1
�5k�������9ı,K�wx�D�,K�����Kı<�{��yı,K߳�S�,KľN�t�ܔݛ�᥹���%�bX��gv�"X�%��{��Ȗ%�b^߻���bX�%�߻�O"X�%�߯s��.f��Yn任S�,K��=�s��Kı/o{���c菁�b\���Ȗ%�b_{�ڜ�bX�'{�s<̗an������Ȗ%�b^��q9ı,K�wx�D�,K���T�Kı<�{��yı,r�ܙ77$�\����Kı/����yı,?1����T�%�bX��߿gȖ%�b^��q9ı,O�-ϵ+�|��n���"c�M&�#��x��s��5�s`J��c���=v��,n�Xٳ�������,K�����ʜ�bX�'��{�O"X�%�{{���Kı/����yı,O{.��.�ܹ�����ʜ�bX�'��{�O!�1șĿ��ۉȖ%�b_����yı,N�s�S�?�*dK�ӧ?nK��&�s2��Ȗ%�b_�����Kı/����y���Dȟ��~ʜ�bX�'������%�bX4�s��m�2I��-��ND�,K����'�,K��n�T�Kı<�{��yİ ��������	̉r�����bX�%�}��vɹ730����yı,N���9ı,?���~��ObX�%�_߷�,Kľ���Ȗ%�b ��p����[��;v�e�ػk��v-����6��A;u�[��F��i�N�95��wl-�nmO"X�%��}��q<�bX�%��w�,Kľ����	���ı?���*r%�bX������P��̡L��~oq����}���r%�bX��{��yı,N���9ı,Os��8�D��A3�~���,n$.\��I�}���I�>��`�'���q<�bX�%��w�,K��{a{�e&l6������yı,N���9ı,Os��8�D�,K����Ȗ%��U&DϾ���yı,O�K���pݗw7&K��9ı,K���<�bX�%�s�S�,Kľ��w��Kı;��T�Kı0@�>��M�]Ch�f��\����t<u�\g]eK8�l[�3�C�i궱�F�΢�Wn�h�a�eͫ��us��`�����
�4�`�f�x�A�n�����d˭*�l��ڲ2�H.�y7m��u����,B�v���D��F0��\�mm:��v,�v:��\l�Ǥ���h�!'0�r�{Amc`�I��@�9��6�-ܗ~ww.���^H��-���th���Y�4tq�(v� �Q�:��R��������qC��H�~���q���X���۱9ı,K�wx�D�,K���T�Kı/�����%�bX4�s��m�2I��.��ND�,K����'�,K��w;�9ı,K���<�bX�%�{��?"��2%�}��~7,�7&�f\��'�,K����nD�Kı/�w���%��2&D��~݉Ȗ%�b_�����%�bX���r�2���e�.nD�K�ʿ�*�؛�����yı,K�����,Kľ��w��Kı;�wr'"X�%��~��3-�B�̻��nn�<�bX�%�{��,Kľ��w��Kı;���ND�,K��{�O"X�%��w��d��f��ݯ`��N݋a�ҷ 6�][w�ɣ�Bݳ�6�7��w{������cK�r�D�%�bX���oȖ%�b^���9ı,K����<�bX�%�{���7���{��������$AZV�'�,KĽ�wbrS��<�Ȗ%��߷��Kı/߿n��Kı/�}��yı,O�/yw��fl�3-�؜�bX�%���<�bX�%�{��,KĿ}�w��Kı/���ND�,K�ώwKrf��K�v�f�Ȗ%����6&���݉Ȗ%�b_߿oȖ%�b_���ND�,dL�����%�bX4����p�$�җ7v'"X�%�~���Ȗ%�a��#��#]���v'�,KĿoȖ%�b_{�؜�bX�%�߬�ݚ�Cw!f�R&�{\��n��l�f�n���&=�{
M�:E�f֚l�v����4���O"X�%�~���9ı,K�{��yı,K�{��,KĿ}�w��Kı{�q��٧.�k{�oq����~}��x�C�r&D�/����,KĽ�oȖ%�b_��؜�bX����ߣ�&���L��w���d�/���ND�,K����'�,t  ET|��`��@�T��QT�<�w��؜�bX�%����'�,K��/���ݹ&nep̹��,Kľ��w��Kı/{�؜�bX�%���x�D�,K���D�Kı;��^��f]��fnn�<�bX�%�{��,K��ES�ER������Kı?���r'"X�%�}���Ȗ%�b_N���f�T�b���de5��.�յ�ݣe��q��ȗ�Vp����1�Z���D�,K���<�bX�'s�܉Ȗ%�b_}���� )=��,K���v'"X�%���ә�.aswm�wl���yı,N�{���c�2%�~�����Kı/�߷br%�bX��{��y�TȖ;�3�n̘R��-���9ı,K����O"X�%�{����K�THdL�}����yı,O����ND�,K�=>�ݻw7wL-��'�,KĽ�wbr%�bX��{��yı,N�{��,K�A�T��Dw�7��x�D�,K��fs7&[�m�f幻�,Kľ{��Ȗ%�b}���ND�,K��{�O"X�%�~�wbr%�bX�}�I�y���.l�Y�f����Ŷ��n�7��1��F�c>Itd��"!��t9F��{�7���{���~��'"X�%�}���'�,K���ݰ?��șı/~��x�D�,K쿡s�͆����2��ND�,K�f}�����Kı;��nD�Kı/�����%�bX�g{��?�DC*dK�����6���tۙ��O"X�%����r'"X�%�~���'�,K��;�Ȝ�bX�%��wx�D�,K���6�˛I�v̷7mND�,K��{�O"X�%��w��9ı,K�~��<�bX�RdN����9ı,N��9��Y�i�&��37x�D�,K��w"r%�bX�����yı,O���S�,KĿ{��Ȗ%�bx}��sW�'�� x	�/�P=�S�oI!Y3��]9�[)%��!�}��X����X�T��@�I0�l"��"�����'�#(H#8�K���A��P��8Ð(�!��H�g��n�����d�����{u���x���/=n�&���/����ij��˜H֝=��;N4��t�ѹ��Y�@`��\8�Y�� ݟ5�����YW	��@��c���b�M1�[F;;4��j�J�g�*wm	룩�����ٕKrƲv�3ݲgmq�,�7E�D�0�t��a��I-;q촣�m�iw7cp���UU�.)��<��n�F��p�I�C�ojJ[�����Y��F����#r��M�W/Q���6��rb�#�7km�q�\�(�%&�]��x���I�[�d7
�HA8|����s]��G����{��\�ȗ8f	��t��!*�� �JbKv�=���4��eH��g��CPgln��@6��B2�k*�\����ݎt�6�v-AY�IvC��qiy`���h�x�s�ٰ.���o\p�s�{F�ӥ��e�6�vv��l��Ƨ(p��ǚ���&[��`
'��ݎpTIؔ%�R$�N+����묒��kIg��8ؖ�@���<Ҧ`ͮ�+f� pd�kz��Z��V�u	��f��!��$�K^'� a��)*�z�n�JXc���F���cUl�AbQ#�Tj�5�-���&vZ�
���r�1 �WZ�.�3m�nU���<�ݽ�۵��-�����;;��<ۓb
69uk��8�AV�L\+&��}����*�yY�g���Z�9ۍ!�u�.�us�gm�kф�ڸ���%m��ʺi^N*'xT5ó�>{�jV	��W�����g7�<nø@��h.�pv�Z0Wm���� ��h�\�ڬ��]�������nM]�� �;x�:��kb��TvE�v��< �6-Z[,v��Ş���r8���k��J-�]K�NPf+��ـyh����.��mk��uƸ��`㭛j�=�ŐkGjN���]�jZ�l�6��cv��Y�v�>�˺�`��]���6A�۫��:ts�������}���F"*t ��cTVA� �����>��ͷ]v�B3Y�8IM�L��h�6���VC,Y7P�:�/���U嵍���ƫn�����[r�z�ڋYڻm�x.r�᱈�n7\����'[�mť
�ucQ�� �l�f۶ݶ��.γ9�ZkC�\���M�uSdq���p���
�ͥ֗��V)Sk���
�Ir�ۅ��a�y��ՙ��L�7����$n�9�sJ]���z�qK���I3�(��gt�8�k�R������ni�0���[7w"{ı,K߾��<�bX�%��ݩȖ%�b_��w��	�"���ı?g���ND�,K�:~�6]����t��n�<�bX�'s�ܩȖ%�b_��w��Kı;���ND�,K���x�D�(��L�b���3�����nR�wr�"X�%�������%�bX���r'"X�%�}�{�O"X�%���w*r%�bX�w����ri2ܹ�.n��Ȗ%����g�Ȗ%�b_�~��O"X�%���w*r%�`c��]��~���yı,��?90�.�37719ı,K����<�bX������T�%�bX�����O"X�%�ܽ�br%�bX��r�_홫��x)�&�!`�7\���s4��g0l=��+vi��}���y ��+v-��ss7}O�X�%������9ı,K�~��<�bX�'r������<��,K����'�,K����۶�ɛw&L�ܩȖ%�b_;�w��Kı;���ND�,K����'�,K��w;�9� *dK��Ng�ɶi��ۙ��O"X�%��?g�Ȗ%�b_�����%�bX���r'"X�%�|���'�,K��N�s4ٸB��-���9ı,K��wx�D�,K���Ȗ%�b_;�w��K���ȟ��~ʜ�bX�%�w��l͆�wf����yı,N�{�'"X�%�|���'�,K��w��9ı,K��wx�D�,x��������ɿ*R��b{sm�H�t۰(S��<�78�N�n��=b�S�����_��ܷL�R]&f؞ı,K����x�D�,K��݉Ȗ%�b_�������Ȗ%������,Kǿ��?;$#�"$k��{��7��{����Kı/����yı,N�{��,Kľw��ȟ®TȖ�{��0ܺd!r��ND�,K����'�,K��w�br%�D� �GD�K�wx�D�,K�����Kı;��^�3snS$�w7ww��K�� dO߹�lND�,K������Kı;���ND�,�#v&�����yı,N�M��M�n�f�ɓ37"r%�bX�����yı,K��v�"X�%�~���Ȗ%�bw;�ʜ�bX�%���mP�k��#v+X�L�i�.J8L㴣�1�ͺ����j�5?��[|���te��w<ObX�%��?g�Ȗ%�b_{�w��Kı;���ND�,K����'�,K��N�s4�vCr�f��ND�,K�߻�O"X�%���w*r%�bX�g��q<�bX�'s�ܩȟ���,K�����͆컳4��n�<�bX�'�����"X�%��{��Ȗ%�b_��ڜ�bX�%��wx�D�,K���sw2�M,�e�ʜ�bX�'��{�O"X�%�~�wjr%�bX�����yİ=�����L���T�Kı>���%�C&ܤ��n���Ȗ%�b^�;�9ı,K�~��<�bX�'s�ܩȖ%�b_;�w��Kı=�ق���6��E�tܾ���N��]lJs��X���;����tf ��Qn[�v[Aۈ�ND�,K����'�,K��w;�9ı,K�~��<�bX�%�s�S�,K���i{{�v̘Kwswwx�D�,K���D�?��2%�}�����%�bX�����9ı,K��wx�D� S"X�~����3was%����,Kľ����yı,K�s�S�,
C"dK߻�x�D�,K����ND�,K����2��ndْ���<�bX�%��ݩȖ%�b_�����%�bX�w{�'"X��	�3����O"X�%�{����6f�Y��73v�"X�%�~���Ȗ%�a�H��?m��Kı/���x�D�,K�����Kƈ';���{��~۾��~���]��J��-ʗ4R7e'u�=Pj:!xz��˖M��š�=�%�/km��g,V�$��;� Os���D��]7/c��͛j�vM�<=qn�A��E*�6�g��uٳ�*�����L��_RIw,�F�ULl�`1#���zѐ�F({>�]��2��/�������wL��	n91u��79�F��N4׉��]x��ח�yt�nt4�$�=�6�Km�iy��rs�@���?D'��X���>���@<�f�u�4��4s�M�A��4��/Y�z� �m�oY�yz����I�LnM �٠޳@-�h�W�y�T��a���ሎM ��h�����޳@�֖.U�14�Q��@<���r� �K4�,�=Q�8e<3��\���p��1��5������)L���mۣ"[p�8d�k���}?��:�L�� nL�$Yr�Օ�fM�M��I'��w�4D�Q~a׬�m�@�z���:��9���,�I�z� �l�9^�@:�4ø��?D'��X��@:�4W���� ��hgZ��$����@�z� �l��f�u�4�B���O��0�X���g�L��&zf��X��qF��[�1��E#��f�u�4�Y�r�^�ﯞ1��Y�y1�ɠz� q���^�帴�J�D�,��I&�[l�*�^����~��UUN�w��_{�ՠ��n�-|�cbm�4
�W�Z�� ���m�e쎳512��:�V�[�h[f�U��^.�Y&mum���������Ʈ8|�nڄ5�M��nƎx�N����ƛ�(���~���m�@��z�ՠ°��1<�b�ܚm�n$��Z�Z�߳
 ���ۙ���&\4�䙛Z���
�W�	r���Z�ʬ����$����̽3ȷ���@=����}��o$�B*V=  &1Cf�y��y�}���a�e������[�h]�@��z+k�?�?}���3��w��~Pȡ	 ��{d���2\v
 `���c��zo��������`m'jI8�����Uz�����f���CX4�H4��4
�[�:�W�	r��b5��P�(�v~����8�_}��z���h^�@�w;���"9�G�r��b4K��8���mހ|$WЁ���s6��;���U��U���� �Pb�'��J#�lq�Nl�Lաv�ӡ-J�F�����B< 1�Η9a��dG&�lu�Wd�Q�6E�����vzq�myӆ`�Ι��d��0����1�ݼ�q4��J�4N�@[bKcFQ:tA��݉^��v5�N����s�jcc#��ˈ2�<˶mm�����Ş�n綟h�ݗ���۞c|��g-y�����ww����d,OZ�vm�ɉ��ptpu��Q���x��M�t`׍��5�Ȣ�j��:mށ�$�@K=1��O��~LY��LmbQ�"���k�m�u��*�^��>x��D�j�= �l�:۹�ٙ��|��=�����K*�(��&D���9&ցIzRK�����ol�s&�[-��$�����'�"��>�{����h	%��..�Z�̛"���]�-��^:m��]��6�\ÇI񫘲F�cs�H�j#�m�{��-�s@��^����"m+�niM���wﻼ�&�<Q �B��t��<�?p�������f�g�߱ ���0ɍ<�b�ܚ'��|���&"��7z �y�~\�j�3 ʸȢ�"��4�z&bb��~�S��@�ܱ�ʬ�ټ�I�8�R=�ֽ ���;���U���K��)����Lǉ�vMHܸ�;b�})Wod�L#����%k$������u�BbLO$����￦��e4
�W�z��@�֖.��&<CI�4s!�E����G3UURC�_-�HM�#Hp�>__��^�4�� ��Ob�F&�Y�	Z5�)��1$��dR@�AI2,8D��	�D�ST��X���� ��B���#"��X�j$
Vڶ���
��0�V�R��1V" B#�1��(��B=R�Q!�JJ���e%�bB	IBVT� ��@�< @ BI��0������BA�Q�%ŉB��e%H����B	""`0  H�"� ����D!2�'�>*�B(��E�Q �b@�`DbD�F,B!F,$H$bBXD�)�!24�� ȅ2T�S#GkF��D�uO�X頄@]|1Z)��舘UE������Y�.X��vGs���������h�f�~�F����m;�>�V�ʻ���/"�)&�[�h�S@��z}�h��������N�wS��^�̅�f8�+c[�m��ʷ�#N�P�l�#�n{lh��*\�@�g��1���?f�����[s&(�LB��rW����hi怗b4�WeF�auQve�fe��.Y��f�������5�|��#��_B������_$�@\����
�Q}|�@ﮖ.��8�!��{e4��ٟ>���}~�{��3���ҎH�It�ãmqͻ��r�y�������}�s��=�f��4�j~	�"�����|��l� �4��:���+ϖZ0�32����D�&f"���@J���>�m{����=]_�)i$�9�"rh4�@���Z8��Tӽ ��� �tu���<���ܚٙ����@����:٠z��+��&%��#�̽�r��1K���	��Թ^�:�=' 
�h�Ͱ���ݲ�M3FS.m���N�v��62��4��ke`sk���x��-t�8�q\%�x{6�gN��N?�Ǜ�cct\]���<�Dq�N��D)t���n:H��.v�v��qv���r8v�q��#"gv�t����+����h�0p�f�sd�s�q�x�n�B�ö�	箲�]����#�m�=3�WD���F����^�w����o�6f�l=�7,q�6��Kͳ��:۔�ss�� m��tsb�2	�ƣ�E#��}4�Y�޳����U�����_H�bmI��&�u�4��h�W��@�֖.�q4<CM�4��hK���bb�\�hi����������3C�J�w��� ��hwW�N��F�0��<�@ܳ@����i��rw�u.W�*>���W^p�^����g��z��jЛ��rvs5�hE��K&x��
�l�f���W�u.W��I�|(V�)6p�3w�N�{��@ш���bbkM;���%�4�
�7 �1	̒G�Uz� ���fL������N��WeE�aWWqw���Y��蘈�|�hi怫�^�U��9����jL��4޳@/u�W���@�+\��㫶v[^(ENz �f�J���5�@��涻vM�vi����,_i���A��m��y�*\�@垈���i怘7�ńQ�1H�W�߳?bA���	������@����]Y��YE�W����˖is1S$DLN`�}V�������G�Ĕ�1e^fhz"f�4�@m�4���rY���k�F�bnM���?�bU���M�r�}��s2� �ZӘ�:�� ��av��}`q����V�a����@756ߧ�߯��f�u�4�ՠ^�ؙ��ӻ��+2�/@%��&j�4�@i�4W��<��\LLcII��&�r����J���������W�W�M�uw�����p��@U�ބ��{���U�H"�P�$�LD�*&*��f��F�wFQ�Ay��Թ^�虦���	����4��0��$��$D���d�J2�v��Z';u��Lm���a��S����f�9_�� ��<�����z���h�W�x�VɎ)��S'$��H�Q���f�xl�����o&��/S@�z�?�?~������@��@��U�ٙu�T]~NC@�z� �l��f�s���/ulL�6�6�4�����"c���������u.W�|�?D�����������ۖ䙛�&n˛��v�L�������Zn�u(��qf.+��21ٮ7@�	p���|~|eW��u�1v�{����E�r�ü�s�ɱD�.���2���j8��E��q���N�c�q�ʍ�ꠒv���q�΍�j���E<(9q�aplg��t���q�3v�5�� ����;u7j�8���m*6i�X��v��)�y�bzƝ�h흷">L��Q���a�p�����S�N���ZsQ��O����h����M;���ﮪ+�ee�e�W���(Ilk��Mث�נ������7��H���$	�!��V��9z����S�k@=�cw#nm�sq��f�{�@���h}��>��z�_��ǉ)�)R����3@����9t��ɟ6ߧ~���x����VC�y��'�l=�'������)`��k�-Û�������t�+��%96�]%�rg꯼�}��@��Mk$k&~m��=^���]�����f�)̆�#�b�DX� ӑǠ����4�?~K�O����y�q��bi
L�I4=U�<�+n���� \�h�K\���8�nI�\Vנr�^�[l��f���ʏ��$&!�%ɗkm;-�1��q>�9�[�QV��<�@���7�g0/42��#
��ʼπu����f�u�;<AUU��cv6�0�yI^^�sw����Nf���������~�$SS��9&�_�ӒN����$�X�H�
EP*���3/~�rI=�{��O'�ȦD�7��X��@�9�Z��z�%����LE���h���l�03 -�,�ZQ���f�>�4�n6�϶��VU��:��tۤ�s��1����6:�櫮��1��nj�)qA*a$ƤR= ��h{l�;+�U����I�b�I��Y�d�
�hSN��,�L�Q�uQI��0r$��h>��@�^�@:��׬�=�}C"�~��!��hDM+��@O4��4.=�:'T7�hޟcF�A)$�z׬��f��[�@k��˥)3(3�l�nx�˽t�9֖��`�T8�^d�e�s��gUj�K�U.zj�����߷ͷB�U�u|��&#����T%�,�X���,Mɠv+������W�޳@�Mn8���@��W�u.W������y�(���.TŤo��9$q��W�޳@�W��9{k�;�&b��J#�ԙ%��G3@h�f��IzNK�Q8Cx� �	$!�@��!�ӵ��Kl��˶�2�Zfxs�nf4�8�����XD$�@�#
����V $@�$H�0BX E�$�i(RP�@�JQ���[D�HV�(�JV2��` ��ʀ0,Ȍ��(��H��P� ��e����%,J%��HB��� �@��!*@
��)J�!��"H@�T���"D���� �2��""���r򧐛(�/4ш$��B*$"���R���eHA!%BXP���V ��X�1H�)��e%J6�H2��ƅ�IR�(JС"�H@� ��HdX�)lX��ŷ� ��t�t�GI�q�&��C�ם�Ah�13���e���Q[<4�u�gB����}7]VB�{v������a��r��FS��5�Wj\�JIs�Ae9\�Z��h����Y���ʍD;�RZ�ة�:�u������}�"���u��$�Lq����3�$�yE�m&�	e��e��g�"Y*Qۀv�R�[I�ֵ�Fp<�)kt�ϗV�7�g�SN��Ý<�� m�0�Ӈj,v��Om[:�p �����I�s�/<�(�v���k؛���\�va��&80��V����WY�d��$MZ�8,p�Q�a�,.���I�j�:Rͻ�݇y�c٦�TmY��O$ֶ&Sc;�<I��ܺ��v�5�9<��wS�U�v�A���+<m7zs������X�9�r톱�9;=uUm�oVlu��2��[u�F
�:<���CFT!�����]�Œ[���������H���f��%�/�A�շkoM�Hj��:t�Mj�/D�+UU n�iS2�mզ]�A�6�k�Y�çn�=:�n�r�mm6萻a���� mzL^��:�;qֵp�
�q�˹N!��dt�q(�m@ KUU�F�ڥ&P�
����)@ش$��-�&�����/F����/gk� �l=mq�p��y�V-jd�*�ڸ)\V�:6	{EUpr�}�>���t�$IiU) �T�.�/Og;�6^�;8��a�u�M��n�������m�L�C����JL��W�˓�2�SIv��(6��r��?��&�f���Q�G9�`+��r�S�3:�L�2[A�u.�٫���pV�˹5ٴ��:/:u�ŶS��v�m��宰�
z贐��l�-eW�p��X&(##��D�����w���i��ٞ��P-qg�D�p\�ׁ�ʹbd�p���Q	2���h.n���gBu�q�qn�zwk��� pOF%�
�B���4�n��ݲ����P@����z�@���Nz�J�s�&+|_l���,>0��{tՂs{6�H���F8��v��)����^k]GcZ�W�R�[;�mv�鴼]sjX'X����vݸ�v;7g\�d	rFPA]nl�Ś�T�A��Z�p��s����tra�k�]�)�e2,��;�����q)Jl�Z���0g�q����Ͷ�q�ܓx���ul�R�,��ib%�d�⊥4�9͞m���.�.�3[�=� �q�r\�L�x.�e��d�͸:���������-�1F�L�	G$��_�����^�7&hs��{��@fe�b�0���<�K��� ��h�&o���O�"&�;Ǣ��VVa��yyz ߽��r�=1U�6�@��w�}]]v"5�F�<�ɠ�Y�z�l�?W%z���I��>�I�yY�E]�]�Ee�hQ�f�蘙��7�97��u�z�J���QɈɎ	�� ���jÄ�#��V5��od��˺0k��GG0Ě����+k�=�hwY�{�ޯ@�ژ�SD�����@=�,�0��9�m������?RJ��G�bb>�D�`�"�M �女��ՠz��@=���ZX���O&I�rh��Z����l��f����I�R0�-�mz��4�٠v+��{�WTp����Y�%�ÛmC�69���mˎ�kk��x��:��1�����#�2'�u�hnf�����Iz.Neee�E%�Y^f�wr�q1B��f��6�@/u��=�'#�bo#x�G&��}��I<��s����\ ��s<�=�h��4�[[�(Ǔ&$Ԭ����Iz����f�����:ژ�J�,rE#�/Y�v|�s4v�^����,���%��7mˍ�g�ٜu=��"[�u\�c"a��`������j�aƹ����%WͶ��?~��n-�9z�&h֕'
�$q�jG&��Ϫ߳�~�������߾�h{�h������"P��4(��������sk@=а2��"�����q3T�y���B屠L�L���\�@���U�y(�1�RM �z��s@�^�@=�� �jrO�#̙�E�]�ΫH`�Y-�2R����`��d�n�Vܣ�x�)&����h+���٠�Y�{ֶ�E�#��S�-�y^��m�$�h��*���"�K�H���hwY����%qw�=���=��b��6��#�����L���$� ��h֖.�((�$YNM��)�z��@=�f�u�4����[��(�L֙fӗ]8�LRqsTp�݁���^�����89��ȗGi�&�I%W8�e�^�9��� ��wQ4i��U��������C�f�.:��C=r��66`�٣�=H	ڛkю�l �� ���ec����~���: ci��ԯ;jR��]�n�[%۝���s� �m�[G=�>;�Ǵc��ٛ��I�ʱ�ˍ�?]����׾_9߃\�Rt�-T�8Żs�&����"�sq���Z}_%�z��çc	��E�;2Dۂ��z����{��oY�r�[4���� 9�O#q���4���>�!�5�^�_$~_���Ȏ`8"c���_��޵k�9{k�=]��,����8��<JI�w�I^���J���^����h&��ƲB!�N'�'���z��� ���;֭z��&��(7"	�\��b�a�����<k@s��M�s��K6��G4���8�ı��@�wW���#�f�U��w!OE�nnrI;߻��&�@S$��{�䓫ޯ@�wW�{�K3R7G�@h�3@j9z(���3@����ɒFۄ�ɠz�W�r�@:��/k�@:����c#ye�]��1I���U��hK��o��O�m[^� �P��n�n����N-'&��;�Y�y7Q�J�^����=Nd�6������3@j9zM���|���F|ȑ�87�rhw��r�^�˺� ��hu��Qd�X<�Wj�4���rn^���t����U3�DL�D���/ŷ٠}��W�|�U����1��@�wW�z���@��@�ѱ�Ma�//@:9��d4�K��3@��[������̇>�Exؗv�ʭ�gEu����Ӭfݚh��2΍>��4������L��f��u5	Lr(�n�����^�{�@=�f��z�Z�K��k�6F�2���L��f�ԺK��/@���T\fYytd^�zffj���	�w�rI����H� 0�$��	ń�#?4J�$���B`ă!b��B!0`F0���BH�"�@�#���>���"B!� H�}W��z�Y�|ҹ����NM�W,�>���R�z�ܳ@q1111��dߕpLn���Ev�;MH��i���.[j�n��j�RL�OS��,r��xO����� �4QI�^��࣍���#�@/[4��h���/mz��b,!x�F9&�{z��U�@��@/[4����,n�"?��$�=U[4^���f�{z����)���@��@��z{��=E��I<>
@D>'!�;C5���n�hF�6�9�l]2��\��� ��E�<=C� [GFt�C�ߋ|���v�ƶ�u���Psu{s�nz�A�F�VĄ��E(ͫ����cN�6�v2*Q@<f��N��S�[C� 6�hU)�
x����8�,s��x��r<d�بMܦۢ1˞�Y]N5	TvV���7�ݪ�N���Xyg����K�sl���*'�y���rnɮ]���[�������O`g8�\��F6��v�� =�-O�6��ƣy#��>^��@/u�����mz���,x��D$�@#s4�$�.�����ySue�5"o6��=��ZW��9[^�[�h����Ȟ$�)�7��"b���@o4.Y��b"iC�|����ل$N(�q�#��� ���;+�h^�@yސ�݄�r'g�>��ۭ��o=C�םGa,��q�׋fUD8խ
㈝U���~�p�m��� so4	֕蠸\�w.��$�����8���������%�nf�8�h`᪅JB6��H�W��9[^�u�4��Z�K��5�D���R=�%��f��\�@j9z&'u�Ƒ2A���Y�vWj�9^�@�mz�9v2�?(ɘ(�?)��� ��wV�݁ӳ�]dv��y�D'1u�ι�0qF�bnM��V���z+k����hz�����E�7��r��3@s4R�ZG�نH��Q�#��� ��i|���c��)
�_N*��,�@H�1H��N����Cт8x)� ����	deX3ߚpFtB���*A0#`Ъ��ցX$aǞ��+�l犇�T�2x*s�T#I#1��=H�`��HH$H$b@��!��VO ��=ȌX��DL��#��4�4�1��"��D� �YFB#! $�1FDȆ[dRF`E��!@��'�N��4 ���W���} ��L�G�h�:�����W�-�o�@��Ya�aQ�a���陪�h
�ZR�z��4}i<�Oċ#�I�{��ZQ���f�8�h:��S��j�8���=A�L��ہ{3IAG
���&̳�˳h4��uź��������K4�,�:��he(���9�E#��٠r�^��/Y�r�^���sʠ�Rcy2c�M����s4�����ʹ՗��7�Ǡz��4��}�"N����}=�p�΂`��>�|�������Ơ���8�����Y�z��z���Z^�*JG1��y�-�P��J���ts��CwC״t�M̒D6ێb�B'1bpnM ��h��h	ʽ1��|�h,�������	"rh���-U�޳@:��sH+�BrL��q�4Kqh�3@s4s��t �"���!$Z}�4�Y�޳@�}V�ucWHq� ��M }&h�3@����Iz�_���"�A"@ �P ���!�߬�MΖ��j`֗���
�Ԡi�8�9�'S[F�zW���V59�*[;�s��^��&�.����78w=p/$\��v��{h7;]�f燮;�\5�*�.A�u�cl�n�'Q��UZt�Х�88y='ώ�/�EL�Sp
�y��oVYĉ91������Li��];����nw&�[6n��p�sh�7)"��|!��8Y�n�M�6�,+�	Ӵh=�mt5��mF�M�z���eҼ�C���H)�y2b�O�<����\�� ����[4Vu�P��q��bnf��Nf�Ns4�������;����`���ӓ@>����٣�����y�:T�h�]�f]a�yJ��w���� ��h4�h�@��4��LI�,���4��h4�h�3@I�����,7i������`C%�-u�,�v60�w>�;\]�x:��:n8�кf�ͷ����|��r��3@s4��m���	�K�6��$�_{�����
�1311�ؙ�����f�.O4]ֳ@:���y�␎9&�{�@;޳@��u����*�1�$q)YYJ�3@�4	��^�t�4�ɠ����g�'�7��x�c�h�,���ܖh&>����2�
g����;tů,eƂ��i����;L�j[$Xc������~�h��h�f�}uנ[k{$��DŊA�4��4��@���������K*$X<l�I�I'~�w�N�۽����ɂ��y�呂u��w5��q�r9�^f�:,��G&h73@#�4��sZs��I �l�?�~Vߧ�[��/���=�Ֆ8d�F�H���'��jĔl4�uv�q�*l�=N��ul*7Aw�M�}$�����>�K�f�},��_m�]ɧ���S&<NI����YM ��4���=Y�,I� ��Ĝ���M �&hnf�F�hr]�h��+�2�P��r�^�6�h�3A�C����k���o���Ӑ;��둳�&�)��}�hnf���!����]S"�_�ĕػe݃���:q�e��v���ιX)�F����vuI0�F�3˺զ�6�����@u�!��� ��hکwubJ)�$�g�S@/�� ��h�@��e�i�q��N���_j� ]�4qT4�h:ۭ �p)�x��mI&�^�4�Y�\^���l�9w&�Q2Ly�b�M ���%.��t����U����1�~�c*�*f�EtRM��v��szq7T�A'Ss�i�
ꍵ%�)C �렧P�ۚϝ�P����)�nŒs;g�����G6�N�������nݻj�Z��yd�fҪp;���S�;��T!�|@�bCT�m�ٜ�M���e���,	��xy]�ջbJ���vGMc󫶳�e�\b���
���͒��]���3r\��u��P:���t|�{�>7],�̹$��f�6.�ƺ�b�b�m4d#�����2�0>d�nn�d�5#X�7'�vs��h����f�w�f�嵼�DD<mGḴ��hnf�>s4	]r-����.�M����iɠ�� �z�?����_g?�Z���wtm,���7��'&�>s4	]r- ��hnf�ݡWX��#��$��]�@/�f�^�4�Y�{��I�G$k!�Qq�Z�x9�!�nR�_�����_2j�w�&�ۚk��p���1b����w�M ��h�Y鈘�@㭺�e7YW�y���e���wﻼ���E� �Vbc���4ŧZ �K4]�uhʆ�ȅ��4��@�K)����u��:卸�H�,JI�w��hrf�ss4I3@�U��&��qŀ�4�f�w[4�f�x��^*l{"�n&�!A�k<@�"k�۸Fw.���U�6�����,�9Ɯ��l� ܚ�l����e4��@�Ѵ����y��&�9&hE��<���$��к��pNdrh�)�x�ק��?�
�u[&����$�������5c��b�$R��z�h��h�)�y�)��GȜz�h��h�S@�u�ͷ��奄ڶ��
:��<�*t\s�����1����2m#2�R,3I�ۂ������2d4'%�rf���{,x��8�,�ɠ^,����z ܙ�������-]+�^*�hNK��� ��h�)�{֧��JBG��G���?fb��� �h
>X�ɉ�������/'�=ޱ���d��Hԓ@9��s!�y9/@#�4�Wy�Uq���FQ��|K��.Urr�\���d�(5�vi�`�"�զ�m���-��z$�����%J4�FVYw�Z��}3T�� ��h��@���E	��"���f�6�h[�@�^��ři(5X��C���}�-�mzoY�x�����x�LRI�In-���	%�>y�U��U���(
������
��P��@TW�����B��������*+T_�
�������E
��P�DE�(
��Ƞ*+�q@TW�������������d�Md���loef�A@��̟\���(�)@
  :     ��         �� (%R���
)B�IUP"�B� H �P      �I@H �QP   �`  l�  (�Ib ��m.}�������\����{t��>���9o��������w}/��m髀 ���}�|���g_��s����iV >�Җm�m��Ͼn��N��]�������     &�zx��� �  P
� 
�7�� ��ʼ�ziw��Vמ��N����!�wϕ�^�+��v�{{�k{���� �Y�u���|�.�U���|�@�Tž�rg�����u�� ��.Y{g{q�^&�[�{m{@�P  T�@�l ��u���o��Y�\ |^t�6�L���/=��qw*� �Ov^��s�f�Z��}��^ =.�l���]���nf�\N��������u�ܛ��o��w�z�^>�  %$@
�� ���8�r�7v�n�=+�gWm���  f�� 6e ��`� �@    �� M� �P � (�  �6 �� �@   �(  P
V@ E(� �   �� 8�=���gr��=�w�+�;x�{�҆��W�w���.�|�  m<|�w�_w����4��}�/;/x�u�,�7'N� _{��'�n^���ާ��zK�=AM��J�  �Q��T�M h2 D��J���4  =��F�R�  T�Д�*R�  ""CRR) ��jP��~�����]/��ڠcvڇK��j"���ݿ�
���"(����AQ_�AQ_�Eb��
�?��?2�����<����a%���l��"C���=����/){~�H�De�=�8c���\�Ͻ>�
@����%�k�O��g����q�7�}��
B��yﱒ�=�.$�I�B���(y��!I������!\�+.1&L�<����|8���X�����п_�o	�ޞ�����5�ٞ�5��]9���a�˘��͞6��.��4��0�0 ��>��
TL�+T}�tQB���%+Y���K�����4��� QU
�秧f�8�����d7������9�}��JbK�.C5)T#��~���jթ0$*�ߔ�S7a�=asI�yBS��7�`Ov�	|�i}��I}��й瞌=�ɼ±�MnR7~>�D�
��]�g�������#7�%��f���<0���|�|�2as3�xG�{�~	r�=�i�ny������y>����=0��a���<��
��rs�N|�	p���}o�8����=�3!��32i��zq�=|=��	sU�&{�aʐ&n��zx@���2f����J1�3N{��l!h�����f��X8�3y�Ō!s�}�|B���<��+�.o<��#Ll�ɚ��m+�5$�3M�B&�=>�D!
j�ϼd�Ha���{�{�}�<1��#3y��aa�,.�}O%�-��
f0�0�0�d�\O|3ݿ2��������.���C���8|�)��{���Ke%��d���`;�����z��F>44�B#@�L) fiSRL`1ؐ0!q��4x��#��8�~�y�{㞅	n��МT���ÅaY�M3XR�ōW4#\5��ơ�E�1�D!���Ly��R  ���)�t	a�)ԕ�^s�q��H����IXFL!���K�K�i0!�����oĆ�F��ˑ�,sB]"B,B$#6�p���G��^LX0�r�3+�!��St�42���	���I1�B���F�����	�y>���(t��mQu��*-c�uW����=e����HbA��@!���,	(B�d�L� ��g��I��L"o���yd�$SX�Ғ������
��p._<!B_~�!�)�d.2�
c�=}o�=Sy7П�v5�Ԅ.��D�+�C�W���Ç F1��`���8j@�����@� �	r/Ǉ���)�I��Ȑb� �5�Ir�233����.O=��L�&� c����^$�(B%�H�2��,H1HH(Į+<�q0=�!R%"_�t>CR�B Nzp��$Ф��4�L)�����t<�fBp�G#IJZH�l*@�x�"h�d� �����&�������b`zp��̆'�Sr$�aHA���B��0��62�3��s��0e�B�X`K!f0�HJ��R��VV'�_���:/�է�b�V�TYYXs��xs��B�L��rG�����34�	�H�)6E`$B��Ћ E��%H!�!D H�"c"E�	@���j���R+	F$a5���!�i�I� ����� �>�<���p�@��0��hA*���B��1
�$hE#B#H J0`a��0�-#q!Ǟ0+�5�P��$(D�O
����x��F�y]�Sl�hk�!��.�
�0��
]�f�NV��0��Ռ�|]VU�@H�q4���B���J�0Њ@ P���chc�CdЍ0epb��jE�U���G�Ca���R4�n���B!�n�!��X�1"��ik1H�5��$$�!Lq P����) Q�$b�S\ 1�b�B@��H�Ha�
`@��,�A!)��ň@0V	��Ƙ����@(��B���X�(D`E Gc�XJ`¸�g=�k.f��l���9R�C���2�Ҟq�o;3����o�<�e�ێ��N�e�e^���l�<����<�L$��C<�|o��M<�u�=�9��{33�
�J��ڶ��o
������U���>�����k��}B���O_��FS���~Ov�����/����_������V�~�����c�����dۛp��^��S�ߤS8E}�R���
`��}p��4�xN��Z�}��f	 �Yr�BF`��7
A(dV�)��7�\7�peĉ	���&L��a`���ɛ��K�Ɍ+c0!�%0afr� �ǃM��\a&:I��Ě�1��F�._��HXR�ЈV���ԍ�<<!~��!C�'�B�0��2�rR�^+�Jf�`<��P�!HH�F�XG�xP�M-���"֛p��/*FlF� � �V+�&�
,�D.C0�B兲g���hB�
�ŋ A���HH��,�@R��>İIf��\b�Sac%8��
aJ`KA)H��%�#\\RK���%LB&�$(K@�6���CE�	�LHG-:#T�FA��B1B!Pz)
�/ :�@�	-��BX�"@ b �	e1%)ЧĔ�9tЁE D*�$R0)�.A���
�R�=�z1�0aL#�C!I�jT!X�X��`@L�`�X@��p !X"�p�P��$�JP�B"H�+$�H�)�l��K�B�8! $��JB!"��A��	��
�)��H�"�$���[���4� FHY��`�A��@�,Z�P�V�����`AO�Ԃq^% �#	����q��BD0M8��&�J�і�`s�ͺD�hb�	��b�0
��@�D�����+��(�
J�kĀ@�P���6B0э1�0�Pč�����C	 P	H�Hg!���0���_�5��i�#C�I�C��-U�� �� �q��K��1̸�n0�1d���2񄤒y�ɳ2g8�B��s�!-rq�RF��e�B# ���5D�RFB.�}@�?	�z���8��$�
�P�҄+ə4�7�d�X���^7�U����,q�e4�x���a�</���+���¡�:o'�k	 pӔ�|�Sf�5�7�Oхso��H�7
��m������;!l�P��
WR,���m�5�㉱�a̐�0�ǅ��9vM<'�����b:Y#k�JS�"�ݓ�s7�y�r]i�4�\XH�|7�.�	�p(�`c �`dn�
$
hc�.la�(�� 
�
$X��¬�$i���:MIL|�iP�\"����E���14k�[�2���6L51�a�h`�3w��aJ��)�!LW@"Y��,-�i��I	 �%�9�9�8��a.$$�C4Ӆ�����A#B�i��bC1����na
a��M�FR�ӓG�(Ʀ�Y
HB��Xf��P���7#L���P"B��p5�2hư ă.0Ȅ�ɼ��c�jG��N�:��wN��~�| �P�� �� -����  h  �M,�Z�I(��ʒݵ]��vZ��j�:<���$݇���f�2�[��ca�B�rr�۵K�4;r�����u�TХr܄;������7?x�Pַ=�79����4�ҡp�8)�[=�[\X��.��l��Tܦ���߀������l�@��    6�u�P�x��3v�kKh p-4ę#� �:��۶��k��I$�ޤ��E� p	�k[mӖA�I�3�$Hf�q� ��  )M��azI��n� �r@�u�B@�Ն���`�!m$���8մ-��\  �  ��.��.���` 	 	  Ko ��[Kh  6���UZ�b��ɛ+$��kn$H�( $:�h[A�j� H  8 � 	 rv�G�'�6�n�ݶ5��H�������
g(W*�rd
۲h&Wl�U*�uUu������� m��[sR��fRWf���Cm��.�$ ݚ�]@:�b�]�GW�lSǭ�g`�U΅`9Z�cd��Nٵ
�l$nD��&������M���F��&ᰶ�z͸�iv���ds�X����+B f���x����Y媦��lX܍@V1OcLIo,�6���O[�,�&ܷ[I���-�m�⊉�c��2c�%��Z�u��ض��m �Wv�m����c�tm@�=�˱���� ������j��y�a̧Yؗ�-�
���� ��)��MU=zmc�[%�g �[��۲u��H.��� ��m�J ��X=f$�lճ���a��+���'Z�-�ݵ�-�  $۵�d�lD���@"N������'gi�B�G:�>������Pm�Ζwmƥh��^U띠[�;l3J���QE�U])�*�W!J
�F�[�Q���pm�#��8�ˡ+]�Im�h �*�ݗ�l\���8����8 ꮀ�m(��H
���W\9W�4�$��5���F�u�dI�i�Z����GD���L�2�xĸ����rl�ԙ	�0I��r@�9H� ����T7`:��l�s`���#��2읩�\a��z� �Z��m5a�Ra��8���u�kZ �vd�m������o�L��U*��V���78Z�l�m�$&�g1�ݤmq��jVH$x��EѨ6�	�\pK�u�pvgcf�Sp]O��m���_@��T��r۵Da]�lN��	dyy���m#�A����I���8wmr��;6�z�Um�[�˻5US��&����Fݶ8  9m$$��m���mG �!��dY.��a  �`mzw�o�����p�<����mU@T�g�+���p   �d�!�h�a i�߃�m�mH8�jڕv�JZEV�jZ\�Iz�%��4�n�mUV�^Y�A���<�Y.�H���i�i;nI`Y�ګ����P�2�m� Hpsm.M�I̐��� ���E��8l�U��m���m��}'W��-���p   sn�6�`Ȗ�6�X��6�!����X��h)�5Z��8�t�w��S�A�� �kC���e�	��u-� A���`���K%6��h�fm�l �˦��H�'��i��tڲ�c�-�� 8��l�6ii0��n�m���mR7m�� m���m��6��a��0Lں�AH�j��vZ����U٪��Ux1��� �/e�i�kH�e�i.kv�鷎�ɲ�r��%���K(m�@�(=UV�z��]���=����M�$ X*�����iU@YV��� Ā 8 pH�� $[S@UUUR�®ԫԫ�h�ͱ$���;Z̜�`� ����-�m��  	�A$�  -��L*WgY����F�U�>>�� 	6�dY���`+iV�U�������'L�����H-�~d�M,��6֢��kz!���� 6�m�'   [I�� 4�M�` l� � 6�8��p	6�  �	 m����b@�6� �h����[l�`��6���}��    8�[���&�a��   
�
���U�����i�d)f�-[6���%�E�@���8��E9��$�l����  ���` hm� H7m�A u�� [F�@N�6�m�]��			n�� �m�� �l ��6�l�$�K/��u隀��U2PԖX���m�X�]6 H �[]	9�m� �I�`#Y�m�� �e�jN�kd�F�K��Z���d8V�%�n �-�*BI ����H  �ZWj�<Bmq�U@Z�Y# .�MY��R�m�<�
ڝr7*�Խ�2L�O��7 -m��$ �ͦ��H�P6زyW"�kM��-�F��북�ć5�i3v7jQ�9#��kh[@� c�$�� H��$  ��l[BB޶�u��P��A��Ya�l�� m�H� l-��v� $ m9�͵�sm� �l�[n�I(Amh	�]��b֪�hp��$��7m���d� �A� �巀���� ��օ� �۶Ͷ HItu��  6�   p  �m� h    � �       �5 p �Hm� %�u[�     �     6�  m���lm�v�||�` ���m�   d� � 	 �� ��d�ڰ��5� [&�`HH{M��aNH h�m� l�m& h�    � �� �߾�   �	��v@,0m�,� m��� É ���%��/]�ۍ��h    [@  M�  ���RBAm	k��m�kd6ͫkh    � �$�M��	��   m��� ��` h �6�  [@ 6�	 p Y)�n��@   �cl�mm (-� ָdݻi8۳�]��� ic-פ����9zu%���^٪��ʴ�DQmk���j�t�U��p �n�yh}���jF��eu�����s� �� 9�oYm�-��K��*���*�(��M$�ݐ�-�����	&�$��k%�pfSSC��Z�����UTUS�d Z��y��:E���� �ݭ�Y'^rړm�� �M��@ ^Idb�<[����d$-4�P���]����ԇ �����  Б���LlH��@mZ�����e����  	�*@ 4k�d����� C[�I�YE���L��n m�I�� H��;m�շvض�R� ��e�ŴHls��ﵲ;8 
畩d����mUR��j�e��S%("�O�� �d� ����m�����0K([[Vm� 5��Ԗ�	�8�u��Y�d�t�k����@�%��3i5�� M��%�wl�l�'  ��h[��ka�[��P n��T[�K��{Eݶ	-��v� -�      -�  �&�Զ&��[:���� Ywg�N6�i8Zl 6ٶZ� $Ӊ :���,�UE#2��tpU�-��U]�=�m��8��+ 7R���,�lp�6�K�[�6�ss�\�$�:X�K�]UUUl��b�h����]v;[p]-A�J��l �`�i�6�]UTT��\aU\��bA [@     ��ulH   ���� 	 �` [E� K+m��Sm�   � $      m�"��ݤ�i�      p   ���   �� �    C���"� ��n�   $ 	
P�  @��6큶�m�   �  �>    ��uI��qn  	    &� �`Z6�� -�h���>� ��I� [@ �l�m ���m�� �
�L�   @�� m    ��f�%  	$��rFٶK(�[� pm�ֶ� �&�[d 'Nd6H p  ڶl  6�   l�i�  6��Z��;qԶӀ-�    !���l�ݧ���^.�jU��Z�a�mp���¤ !(\�ڀU�:%�x�-���m ��v����[Ub�%Cmv��䃶���H�]�����w���w*U�C$ EY�7� x�����<����^V�#��S�U�) C�k� F��A�ᢠ�j��j(���P8�q�|�W�$��O�<G��5��0�נ��U=U�*���� z��DU�bE ):F��� �Az��Z����ɪOA �*o����'�� #��!@� 0���! 1H�0�"^�����S�"�S�:��:�C���>�� ��UEV����������8�A�= ;�P�E�׬1�&��z|�!�����}S�XHI##aal$�~U�US���C(�.��eC@u`�����_*��"�!�i���*+�?��*H�T'�;��{���{�w��� �HSCm���\uͳ��>�m�ڸ«m6����ٕv c�ŊY7m-�ƒ�=����%�ā-7\�$wd&
X)[t%����iUy�^:�����֙�%� ���A���n�n�D��f����t��X�а;;/g��́�x������T(���9�p
���������/j{\f�cK��	��M���3ǧu�`��yc.���θ�pn�����֞7bv�elw�k8�!�Jfl֓m��(�y��9CS)tlF�ڥ{)�R��ke�k������u,k�L��C�R��X�h��[��)zt�u�D�ˋ�[�&Hf��j���9�ڱX��k2u�,�-̓vܗp�������N�F:�g�{!:�svn1m9n��2�����]e,�I�"��c�H����������]]$�.��j�t�ld����6l���m�+�(��=�@�CvFA��n�r�Tc"8�����,OݭDPR�˵�a���-խ��jG-��袠�vy5i��eN��e�H�*Ԡ;!8wf$;Na[v��=]�v��@T�2�*�Jɶ͛`/[Z�h��\��MA$�l� ��q4��l�L��l�J�u+�T�6]�	D�\�ì��;[# ku����-��[�HT�������۵v�؍2�D=�j��;Zz�p�ar�rA�Kb{.�+�*u�6LKӕ�U�ѭ]�.z�;T�i#���cVN���9�@���헣�n����-��.��[�1�\l5M�n�G1ttkd'H��D�:���\y��y�Zȴ�^��Z��WrN�$Itv`8�
T�HR��[V�$im�&� -���	��Uk�jR�j�UV��v� U.��nf�i���k��ӭ�
PK��Т�j�M�͚�@(�D�UU�"�c��yA8=u�m�v���s[��~�t��B	�QB
1P�U��� ������Uz�Q��{�~�{���6�I����ٹ�D딊�l���-М#��u�E�L>�i��N�㧔�ҥch�YbƖ���F�k��IU�����9�L��@�8�v�븁΋��8S�X�x�歞��6P'Z41xX��U�=��A�ch`�s����o��j�]�+�϶��Q��tg\G���M�WZۜݵڙ�w����T|9�0��.fVRe�p�%Ƕ���˹�O���$�M���I�@�֒�u3zX�����\����d���YFT�b.���g��G!D%TV��oQ�v�oKw����'(��o(06a��D����*��*8��,�o; �����Ӌsgk�$�&8�(# �0N�������oD�+���� ��#sq+�]AN�e��V+crmu���'W�4��5]c���H�m�ea�7�����oD�=:&6DYTM�WE���� �m�2��Q	}�y$��{Ò�� y��m�����j*�NTI�XK7��}�o(0=�����]ىeԄ����ޗ������������[��TA�b�Y����o(0=����{���`v�O�e��:�.J;x�m��C;�ۜCչ�bˮ�$N�UJ�L�8/PVѦ�6�������Y� ��L	���;�UաX�/,-$0%��0wD���w(07�A!b�b��ZI�{�o$�������1�X@b�Q��F�~����'l���$����R�Hiԧ�X�8�36q`K7�`� �%�V2�U��!���	f�L�"`M����?]��5�G��l6��Y�6N��qդY1��3�\չ�����L�V��A9�r�����X�8�36q`n�gJ��$�!���wK�
&G���7]�9�����SSX�Vb+$����(0%��LӢ`t�e+��RWV�+!���f �Ӯ���&2�""�I\D(z��)��s�y9$����l۶l�qE����D����P���P8P'De9M��J��(&��ۧ�v	�˷g9�s<F�����X͠�d�� |�� ���}��J!B����`{}�AJ�!�R�Q�`M�o(0%��0N���M���ڢSQ�X�8�9�,�ޖf�,;�6�jJ�NT��䧫e������`�`����$*r�Ӓ�>��`{�RO^q�]�9=�����(IEo~~v��h&Ʈ%���#��
��/k��4,��|���l�7W!��طd��c�8ݩ���Eb�6kl��4��s� �k��\��8��d����;oi�s���ל��M�@��'JJ��.�3�q"Ƌd/\���K�qy�r8�$I���T�Kf�n:�u��8xv�Wf� E��͎o��)nq����6����rh�2�;���]^��ʉ5�Ǝct�5�nD��I1��:i9L%!�`�N,͜X���D��)��.�R0��X��P`K7�`�o(0%�]�Ո��E�L	f�LӢ`M�oGL�U�E��bT
�i&��0&�����z&gG� �H�өN(�;6q`nl���f���zXԻ�G�4Ӊ��u�GG33��tLN�t�q��7��sm<�n.�:�pm�QJR�ڢSQ�|oO�z&��0&� �2a���S4�i����t���=I��W�}��\֘�����w,2��C�HT��M�`v��;6q`nl��:�zXs�I:mJA)ԓ����|`^�x��xn��M%*5J@����Հuf��l��7���P/��F*Ee���ۅv�\ղY��ƣ�;*h콬�r]��8�\i)"(�1���`Y�,�ޖ�P`v�{$Uh�Xb�EM���n�D(��Om>��� }Y�,Ώ�qA4�J�)%��=��'����GӠ���l���y$>��`�ʕGNR��D�qXf��:&�����:L��u��	fU�J�*`N��{z&o(Xf�Ձ����7���*@EHh��� jݎye��W=+p�4e�E�z7F�#�x,2ˬ_,1&��ܒ�ގ��7����������N9,�M������k� ���:"d}�΢i)!�%5"�3{�V���>��`}��X��RDQcq���:!%3�^ {_^����BK�����s3��rI߳���3M��.Չ$��D�������{N�`��$ی#�Ҍ�8�ԨJ7��D�0�I'[�����8��.1TEE�����I���-���� �� �wK ��TTt�ڢS�8���脡D�{G׀���>�78�Ӗ�NJ#n��H�X�oK �;���>�`fo]X���Bdblu*�� �Șܒ��0V�LG�u:MJA)����=�������`�Uo)p�����,qpx�v.�G�\�-��rnt��8��8�<C��4ik��8���B{,��gZθ�yo'LJ�X�̆�"�rܻ[%y�.�!qՕ��:����a:q���w2`�Z���m�O&Jx���f�=�Vۊw^���|~|_�����L�&%��Da�pG���E�*O*APIN&q)A���k/F���{��n[���f�+�W�7C��4z6�k��v�POKӮ���b�Г�š��[A��I��^�D�=�&o(0%�� F�-*`K���t�76q`fo]X��(��R�j�n� >�w�o�ه舅3���WzX�:E�*bN�8������w���&A�"`:]���*�Qj����=�l�:(Qղ�� ��������ݟ���F�h*ntlkg�\cN�ڬ�����;bV�S��k�C�6�NH&�)P�B��zXgt�76q��溜�|��$c�Sn\��{�{��UlQd���~�����&�u(��V
�H��&o(07b�^�D�7dL�JA�r�MH����b`�ے[_H���Y�˲n� }�]��B��>����t���V�R��!�J��
�'Pj���I��3�����t��e㗴l��g����VZ�nS$$�=ޖ������u`a�,͝"�9R*�ԧrXz���}� �쾼 ��x��h���M�D�qX��V��������G������C�K �_��$���.�)'���$ 2	 ��	�E�R'�%�$��#| q��uP��tT�'���� �������y��o$���V��e'$J��H�Xz�el�� ��^�����u�2�� M�&�R�M9,���v����|`}:� �
B�;��|��U9��M�'N�^�k�:q9��{Jr��/�/Wk���ĪK�)]5NP�!N90w��`fl���zz�@f����zy�6��U�䪳 �����
&N��׀���76q`b����nU�/o�`��������YNTڕ	Q)%�}�����Ł���rJt��N��q�����'������YW���I0=�%�%wGL�-�`n�����A
S���A��I�IVձ�&اq���e�9ڻ0�k�ͷ&��_�*&B�e�Q���<X,[��>��`}��X��i���j��$�����LӢ`{rK`v��}�HM�&�R�M9,��O��~�76q`|�oK�u���a(����I0=�%�=�%�={} ���TQ)���t�����&��0=�%�&�-*I��$j���Kc	�@�������%s���݃J[N�s"��nY��4�m��X�^��v۬�<g	�	��{¯`�����.�d���N6���km����m�\�$���۳�AH4�:j�V���櫢q���N�wm����՟\35��Q��a���̑���a�v���)Wj�8k'!�������ww"��4%)1���n���m9���m�+��uXu\^4u�$t���k8P,/1_��럓 ��ܒ�ظ�7����Rڕ	Q)%�f�Kے[������%k/$��)RWi&�$��(0��n����9A2A)��V�ӆ�] ��ܒ��.���Y�uj�K���wD������q`}K��R���&/�AAӍ�ۛ�Q4�+ ��͂�z�rt�I�+vق�g�uv�T^a���`����A�}ս,�[K��DQR#���m��(���f ?� 7u�~S#������)�����zx��޼:+P(���׀v�� ���UMȌ/,.�VȘwD�������}Q9Lm'($$��w�n� ��f ?��"%���pb��p��tF�@��I+b��[�����
\�nd�j��PWk������w��v� ~� ��x)k���2�Q��RC�3ޞ,����,ݜXn�
c��cT�I�vrI;��w�I��wyD�k������A��r��%E�J��ĘwD����P`I1�.��DEHT�Kwg���З����9ou���:��ʪ�@z덞mk�ѕ��z���n!��Z�X8�sp*�pSU+8��T��7hF�ͷ����0	["`�w(06�u��Fe��aw�`�D�;�&�P`}�8�7_S��Ci9A!JI`�w(0="� ��&�(����W�B@�i&�P`zE�c��nۼ i�5W*ʪ-MU$��P`K6D�;�&�P`�Ͽv�m��s�0���t���aF����W�=|~>����]g2���g����V��?Y߿&��0'r�Ӕ��sԔ&�R�CrX���;vq`}�8�9�/=�r"(h��V�`N��(0%�"`�����mJ�I�"i����q`9<���]�~S����	U7%�����!�,� ���A��l���4��s�a%��m�jn�錘Z玸��nh:z6��J �F�P�|u�ϙ�-=��ƭ���Qe9���PW�+�u�Y��n��\�^�����.)9�a�L�OM�:݋���C��s&��3��9I,ȵۘ[D6���t
�ZC���
l��@��n7�]ƩP6l�
i�lC.�����UT�v%&�Mmh˻pޅ*�h֨��ݽ�{���nضo/k�//mv��]rʵ>;M�}�r�V9��*�����f���Iw:mnt�J��>w�=�f��g�:M����%'I�$�BI,ݜXv�,	fȘoD�*T�LH��VL�ـ|�ـ9<���I%"��E	D����>A����{�ӂ�A�A�A�A��v~�\�K�2�Mݻ���A�A�A�A��_߷��A�A�A�A������A�A�A�A�{�ӂ�A�A�A�A��y�pA�666?}���˺[�SM˗7x �߻�x ����8 �w�� �`�`�`��'߿o �`�`�`�ߦ�?L��wK=��n�@�cXy�������6Bv֬���
[S�պ]t�q9G���~N�������� �`�`�`��������lllg������lllo~�����lll~���7&fn�-�&ܹ���A�A�A�A��y�pA�#���$�UCQP���A�A�A�v��x ����o �`�`�`����� �`�`�`������L�6n\ܛ����� � � � �ϯ���� � � � ������ � � � ������ � � � ����8 ��~�f�ܷ4�M�wx �߻�x ���~�|�������ӂ�A�A�P�V�A������� � � � �����Jn�̤ݐݛ��|����~�?N>A��������� � � � �ϯo �`�`�`�{�o �`�`�`�~���337-�XZx��N5�hU�Vq�� ���ytg���쵩Q��\��X]rMo���7{������������� � � � �go�����lllo~�����lll{�y�pA�6667�㿶�iw2�i��vpA�666?�����ȏ�*�� �lo����>A����s�pA�666>��?N>A����v��ar���r���>A�������>A����w�� �b��C�:�:�� �s�<�|�����������lll~����	��������lll{�y�pA�666?��~�|�����������lllo�~�>A���������3.�-���36pA�666?��~�|�����������lllo�~�>A����w�� �`�`�`��w����\�^�N�0q@8�����L�Ʈ��F�s�hl��[���s��&H]3F�������ДH�(�%
g�}x��x�m��wO���C�NP8"I`��tL�]�sw� ?�:&O:��H���($$��������ş�Q�����xϿ^ -M2�;��&��Suv`t%>�`h��}��IRE�UO�)�0E>G�Q����`����UMʛ��M���� �w�~_�+�~�ϯ�|�ـ?����,a��v������vN��������.�e�<j��V�?���>;�"Z�yU�*������7�l�>{l��!(�U��{�X������������m�9B���� �^ o��r������cc���D7=�ŀw�w�B�2=}x�|`-��*��h���&j���3�>� z����0?/�"+wߌ�~�d���
*�U�]� o���"���=����]䓅>"�@�H�0� �`@`D"C+j���aD��B	��HFB, D�)*�,��$��e��B �a���$,�&� �֭��x,�1!	��A E� �l:��jDLd��K���I�[
5$F�� �0F�"���[ H�f�p%����V!H ��/ !�O`�h��'�a �E@���H0�U�H"�B0bDO�g1D#=�Ex�!��P�h��E�Ȑ�-	c#�����;�{޷��$�}ΐH,�]F��u�S۞�
KշIv䋱g�jg��vj	"�R�f���/L��x.���D�2\��Eu�r���E�[+�7F�i;+�l��� T�S��Zɳs�Z��Ŗq���od"wRS[�$��UȸT����ɛ����NM]�󇎨<,��#rx(qj����Z�W)qeڙv4ԭ�9x"v��cF6�lt���K#�5��uB�i[������9�'k�ލ�n�F9�v��`U��Ƀ@���qq�ƍ��\$��B�T��'7N^�h�fH�iʑ��6�	�ے�l����N{�>izu]�9]���]Vz� R�P�9�<1ڝ�,���;)λPc���rk��3��n{�ɃY�������rݹ5�p/e���$.ۈ9���3�a���!��&��8�3�WM�RK p)�5e��RsKc�1�����:_��ݭ�@u�du��l�1�MI�9�]�V2 ��^�$�H�h�e	sl�Z���2	WK��cv��Ӏ1�2Umnms��S�5�����pfݶ�^�[b��{(j��B�m86]�v�h�(�iY[�@��v2�uvI�]�`��Jٶ�@*����U]���j	 H7E������4������8r@U*�*�JD�ڝ�<*�p��@6�Y�$�5�߾ᶗbZ��&�.lm�	cdeA�M�^q�<�ָBʜ�8Ay��1)���&X��!.U��kl�<��}��UUK�!)M]�'OV�b��I�.��m��\N�l9uI��"u�e�e�l4W)��%M%]<��=���g��j�m��M kiwAd{^�؃t�A�A�>2�;��;�v�z������$K��/Z�f�-��P��X
keZ�[h'^�۶�n6i�x���d�m�Gi�$1�ulrm͌@WUUT�f�TI��%8�U8@O-�j��WHK[���|t��\�q����~(��`瀿��	C+�W��E7(QD�t*���8�'!&���5�s9m�wc�^۴�]��{��-I��^�P�<I���A<��n��'����}��ic�N�Zл��.��Ը/Z{���>5��M����qr�5l=�������ʽ)�
&��؋	q1�%�v:��Ă�bU�W <;:���[�oWs���H�D�B�	�N��:l���<c���w����(����s,��ԝ�l���5�	�h�Fqvl����m���f�3� ~�������m� �k�I%����5����]�2i���������?�����߯ 9��x��3���ܬ���)RE!`�ޖ��,���U��{���;����35J�i�R�t�J�QWx�L���0=�`r��;���}�I:D��!Q9,͜X��q�h��}�����-P��n)ԝ�V^�ӲYT���	����tcb��Q����i�m)PI�J!�|{��4�oD���\�,��j�ɛ�r[�9$��}��]@p �<�ܠ���vH��Ix�1$�oD����(0	�t�>淪�D�r���Kwg	�����"`z&]R�]�Y"�Yv������"`�wg՛?uH���m��T�H(T�g�x��F�ڧ)u͖,�7N�C�1�9�9;d�UeժIZC^܉�v�L�P`}�8�35J�i�R�骕i�`�� ��f��f �����Q
ɻO�&�JA)��������qg��%j��9/�����<ݹ�US*�yj�//����� ��u.j�E5Pc��I���wb �o&w(0=9A�t��.�-��-��Äh�ч@u�)s8K�f�e�)Q��g.˺��;�gI�h�I?[�0;�A���	{r&�_JJ�$R�(�(�76qߒ3�<XZ���77���~H+���#��)��0s�0>�w�$�����]�ս���)RE!a�竽,���7�l��R_�J����}��9���M8�t�J�4���`v����O,[������LjTq'M�f�5d����)ѵ�%�'n�\ݰH[g�(,ׂ����+)"��������,[��77���ӓ��R��r�Fb������0މ���]�Ȧ���dbN,[��77���������/��R�I0މ���NP`K���})+K�V�bL�P`zrf �Ӯ�}��bP�!$(��:��p������@]��)sX�>鱱��{tm\+Fn���<�=J�UUͣZ�(64g:�&h��h�v/Uݴq'9Ij�өہ����qaB';#T²�mdr��4����4u���$��D���^p���(�I��m�)kH+�zv0͎��u�sr��ۍ�Dvz���.�	m�O5ȌQz�T
�
�[hq�ڇ���6�Y��nz�U�?ל�x�L�wr[���Q6�>�v�����ݛ�tk���Y����z,�e}au�5��o�����6�gӮ�}���D(����0�oYP��5JT�HXK7��������=�<Xv�,�eu$� 'IT��Ō��`M��(0%�L`n�Hfeо)U��$���NP`r��`�����ԝ:C�)Q��0=9A�/zc ��yA�ݜ}��Y�K�m˴b��f�D�;v�ԕ���8[�ؗuzĒ:��&�lڞs:q5g�t��������В�Cw��y��A�*��(��3;��~��Tv�� ��� ��~_�J*���_���H�r�B9,���,ΜY�ozX�,���O���&�MG!�{�ـ�� =���B�=�8�z�Ц8RR��*T�ٽ,3�`N��P`J��J�}��,��:t��f��ke#N�����%�2;�n�![����%JI�P��TrXgt�3�A��l��7*J�Ŕ��$*)%�����ꤍ�O��K ��oN�颜�	J���`ft��7��
U
.>IE��n��ـl�D��Yx�YE�� ݑ0������ n��U�M�r��U+K쉁;��A�/d���>�7c�׬e'Ѝ;�]��;c�Z-�@����(Z]�3G5]c�r\B�ΐ�`N��P`K�1�nȘwW1tn���iI3�,�x�7xݶg%!�ˬRU�f�J�J�H`����7dL	���݊Ჺ�q��*�ܖKwޖk�0y�0��S�5�"j��`�Ni��:D�E$�;6q`ft�M�쉁�d�Vf+.�"��5s.���������C�8�z%�N���4���ܤ���	J�����ŀvoF�"`M�\�O�A���/�&�LvD���ؠ�W�|���̃n~��pRK ����۶�:!B����� ��~��MY5v\T9DQG%����Ł�������3;��WusTcu�C��X�l�9K������>�`�)����n}����v���Z�7;ȝ15�7/k�h����қ[�q%��_]���Y��ݜC�^��v�ɰ�ZY�� u��s' 4��g��r�Y$�H�=Ff�O0�J-�>{�r
��s&�5=�ěuev͡��u&��UW4���ro�C���Qu�fqQ�����r�<���g۷��=���Z�ny�J�l��s]&�u ��R�����7̈́m�:y���kCm����B�b�۰��{����v�u�L���Ƚz%!B���J�C@7{��37���t�����,i�^BrT�*�ܼ ����;g�%��_����NM�%t������Ӌ3���,3�X�SN��(JTu5V`~���� =}x�7x�}�<X�Ώ~F�dbp���`t(����s�0y�0�BI(����ql��gg$v�q���U��T�r��c�=��d$Y��\f��ylΐ�~@7{� �� ����_H9�Հy�W+&�˹EZ.nn����0P��B�Ir�7:�����y��Jdr�'�1��n!��,�O��,����J�o���7�_� >m4��t���j�C�zc ݑ0=9A�ꪾ������+�NJ�'C�Q����`{�o���n�x�1f�2��q�GF�m���R��V'�ڮ.d!:ѹ�\�H{�\�b�����I��I>7�Ł�;f�����$�~K��^ �����9
����Ӌw; ��gN/ߩ#y���Áӌ�Uf��Հ�w�)p	I		(�E�#	2BH��"D�c���gj�FF	�A`�H8 �O]U��P#�B$�g��<�xF`z"�$�$�H�u��b�r"#DDSMy�j��������Qq�('��Q@S\�ê�x�QO��_��~����Os�M��$9A*)��R[���7}<X�8�1gs�>�Ϫ	�R*���K3��n��|��������5w�R�m�)9���dn��Q�=Y�79@���Ny����JXg�CH4�A7��,ΜX���cwУ�޾0�˒.�EҕSj�]����c ݑ07b�v(0;e�iJ�'C�Q����`ft��U%����վ�;�l�MГ�����A��{&0R���Q07:.b�	J������Ł�d��"`{b�ݐ�P/��Y��dηM)�D.�,R�������-֋�n��p!q����ś��3;���A��$1]�/�ؕ�ic ݑ0=�A������)���$����P�3���`��K�1��n!�Ć�P`n�K`�&�(0IR�Iv��-R�I��vM��{���{�w��Ex	�mB��Q`�L��i�r��s7��^UoMrH�Q� �3�Y��ɪ'<�N�z]&���Fb�}M���6ع�l�Nڵf��ZKq��k:��m`.�t��.�6��Y8Tt6�l�.��Kq<ocGlq���S79zP*
Z�g�� ƀ�Sţ���X� &Ҕ���c���5��h盳A4��瞳�ڬ���7Q�������@�j�s߾�������;^�I�`A���+�� o=+uʭ��<i�6�[��N���[3�߻�`{b���D���]ј ��.�|�`{b��f����`f�\�)
�<�0=�A�n�Lw�`{b�����5ӌ�N��,3zXؠ���L�J�+.Ĩ-$�7z&�(0=�A�n�Lߟ������d�<\@A���B���4c;�������%,<Z��ny��	$����(0މ�n�L���r�j����r�Ӌu�_�(Y	$�(����/ =�� ��ـ���	]�Z�X��D�7z&�(0=�A�6Z���T��(�T��I������(0=�� ���s�%C�M�I��9,���Ӌ �ޖ��,��}Q�)�P�$3�Z͖������F�ݷ,J<�]X���	)�	�(	��(JTtۇ�f�x���`����:q`}���S	Lm8�ň`� ��ؠ���L�J�+.ժ�"�Lw�`{b�8�¥@PS��s���$���yݒRW���YX�
�I��lP`� ��I2�]��)x��C��D�7z&�(=����������E{W=Ku��������\E�6{;]Y����3ٺXݵ^�Ë�I#�މ�n�LlP`{b����brTI:J�nK �ޖ�Ӌ��Ǿ@n�����Z:�Q�I���LlP`n���0މ���p7�R$�:M���7���;{� =�w��$�%BJ���0z���m)Pcq���37��fwK��Ł�Ӌ ���LNJ���eۢZ:Pˠ:Ѩ�5�\k�Fyw[�9�2H��T��)]�UbE���D����v�J>���Ο]j�*��$��������0� ��k�%6TI87!`ft��76&�"`{b� ��YF%�����*I!�n�LvD����P`vr��㎤I��TrXgt�>ζ`�`���	����Dn�3.~�낝9��[u��A��ź����:�c;�36��gԛ��@��mk�_�ÕW��ػ���~k���X��;!�y��<������HC6����l�s�#�5�	#x6�f{l�mf�[!ԙ(:6N�q�	uj��Am&�O�Y���թB����=���6r���mlU�b�(��Ng+v��/��~�{�����ϙv��t���KN�K�U�ړ�ãT����bI����6Ri(�J��ԓ@������ŀnoK �ޖoE���HRIԔ������`�Ӕ압)4J���N��,3�Xv�,ΜXϙ��Q(�"TR; ݑ0=9A��\Ο���'�UJ�V!bLNP`n�ٽ,3�X��{��%*~�J�2��C\�p[�>���C��nv�����������X��Ą�H���n�x���`���%�^Q�j�$��7z'_VU]�쉁��A�6)]N8�D�4J�nK ���Ӌ?)�޾0u����*)]!M�ʫ�����A�n�LvD��躆�B�N�cp�3:q`���3;���Ӌ+G��D�rDDFt��Yvx���i2��Qm�4��K�Ǝ��k.��8	�T�Dbp���`���݊ؠ��&X�]+�j�H�� ݑ0=�A����D���A_�AX��0=9A����@��Lξ� {�x ��sJ�u%��9A�v�L�D��Wߖ{�ŀ{��@I?6�iJ�䅁�:c �0=9A���W:R�_a]�K��C�U�Y�6^�(���N��q���sn�p޺륋�JzA���V�m���D����P`��Lu�R�*���Ee�����݊��`������)
I:��p�3:A�v�LvD����*Veڤa��X^!�v�LvD���1 ���QF��w��O}��;n�Wj�X�i&�"`M��P`���0��P�*BF�J)e;-�g��I���E�m]v���G3�,Bk��v1}�ZAX��0&�v(0	� ���p�:P'(�,�gB��׀�׀|�ـ�R	b��-R��oD�7dLl�X�8�;9J��R$ؔ�6��������;f {�� ײ�(%JRJB��XgN,Μw�[>��7��o��������IE�	 B !$ @�� !@��H@�`B0�I	F1����1"�R F,�!��"�`A�A�C�;��>|����=H��T�0#d	$��x����M�����+}�<H�#%t>C�"@�b���	��)�!�+R��(������x>!Ǻ��H�0�$�!X��#?F�A�T�H1F��~�����Z춋h��Nu�s��猧,�/m���%lV��Y����i0	х��d�K5�-ۄ��������sNS����䭅�Ƙ�vGf8�$ Sn����Ui�-�u��ؓ�{n��Q)K$ݨiiV).{S�v�fʫ����H��������k���&�І{b7=�}�4Y\�s]���\���ْ+���]8�F�i�x��qk6ۗ,q�v�Ι��{8�v�I���֡�\q�[FQ<��jvN��'cc�UՇ�*��[�k�P� �&��9����ld���NC���A������Û��N|�ynx�^Wb+S�gBM�luR�=��u�ejvDnGUk�H���Q�=9������֞j�vLc�.�7\n����qL������ݮ���ftT�� ���c��.m �خ����n��m-F�� :޽�^���N-�B[ڦ�kRqv�P�v\d����gMmO.��t)�vnCs�W����YU� f��P���p���IS�&n�)��T��ܩ��cՍ��I��]Hq][<���t� ��qM��j��lۤ����]�D�6���A�Z�P�` �ݷ9m;m�HUe�Bګn�P1���:�N��<��UK���j�сl��d�L��m���#5��nIjB�p[%��E��Z(d�z��`kj��^z5�����#cD��M#��Ͷ+��H	79ck�m[$�5�]=$�
tV��-�WS9��a9�8�y6I�^ncn��,��OP�1nԁ���\r�7e�E$5�nxvT�5p���d�8j��):�8�m�u<����q���l�v����!n�ثg�{v��15���UWPrA�i�����A@���m-��p�
��EW�{+�sU*�UT�;j�j^�l��SJ���m�B�t���^�Dٵ�P�o;h�Ӏ�Qk�j���[0��!���r��fmll�v��{ݽ����ʞP5���#ɨb*���|ʝy�2��h�J�sz�X857<U�ԐI�i��盷 �m&�q��\��5�q�#Y��̙��On]t��wcs�H��k��ì�h�GGm�0�;%�.��1��l�˶�K;:X�wQ۵h�P4��k�7JȀ�[+��팹�t���2�����RF����kV:Nt؉��mt�G^��6�;L�r,�#i���W�l��t���@Z�g�Z���bVꪩ�d�ww=&i������4�IM�$������7z�ZI%��>�$�l�$�o[|	ҕӌ�N|�Go]KI$�;��$��������K[�>J8�%�H)*ZI%��>�$�l�$�g_|�Go]KI%���J��ԁN���%�g5i$�:���;z�ZI%��>�$�;�iҀ��:�r5i$�:���;z�ZI%��>�$�d�$���ʆ9
%9w���I6K���q�a�����Ǟ�N�8(��M�4� �E@�Q*T��${�u-$���|�Y�rV�K3���I%���m7mɖi�s4�[m�=�s�>
�?u~�R.�ZV�K3o��I#w���U{ʇ�ߧ���.��?����~�������H��i!|���K7�X7I)
�J��p��f�|�Go]KI%�����$�gEi$�z��M��q�����i$�y���$�l�$�f�|�B�] �M�e8�2P��Vr�@l:�K�W*���wf�x�$v���а⨔R� ��i$�y���$�l�$�f����G��R�IgN�DC��#���q��I.��_�~�M��z�}�I�]KI%�����%���R��#��T����m���;<��g~�� qQ��3����YӢ��K{z�D�T��I!��/~k��ZI,{�?�I%�:+I%����$�͔�EI����-$��;��$�ݝ������H��i$����w�s4�����9��rj���i[n��l�kFv��K�@,�秃��V�K=�.��L`n�gGL^Ɍ�y]t�"����Ł�݋ �|�`�7Y�"!L���.SRZ����蚳 �}� �|�a�
��������ռΈ��J)H�RU������w�{�l��
!,P%w
!&�$l�Հ}�ݫ���*��UW4��vȘ������ײc�W���������\��ڎ�`�J���A1�՜ss������7�ل��]Aŵ�c0%����~::`z�L`�&�\�uv�`�V����^,��J&ON�VL�{� �w� }����PQ&4J�nU����`�����[�<X��Ձ����R�$������=�`z�`tO�{� ���2�"�ڤ��`n�gGLO�� �7xDOеlJ���h�jE|��H���=2�����Ĝ��mC�m�;=���ݶ�u�B��Duu�eu�v�[m'2t���X�ɫ����8{�NX�n&��y��x�Xú�-])��S�ض�>�6S��Oj���m cj,��I.�X�鶻X�#;K�rr�u��4�D�M�W-�c�mk�[\$e�n�˙��!��3�m�N"�4����Ѥ�l�*�u�)���&�f^�\���C�9��Ј�s֧�f^�Ibp#��޺�>Y��s�z�U|�w���y�22(�"AIV���?DB��{�x�0=x��P�Fs�J�������q�o�,͜Y߿%�Ҡ,�v�jJ���UV�DO���y�,��u��� 7��Q�E�D�RHX��V�D%�����u���0�P虩��Ǥ��*� nN��õ;Ԍ�=+���nM�n`�IRBI �`�T#r���+ �7x����B�J?B�K��~ŀw���Ҩ�JI9DR+ ��u��~H����׋ �����I~�
��߲��T�
�J��rXޟŁ��u`}��X�t�7z7]M��4�	�a�ߩB���,�]Ӏ�� ��ـl룉Q��E)
J�>�ܬW�Ի}���<X��V�k�j:��Mf��2݉20q��n"�]vD���==�Ms�P��t��AӐ�F�)�8�s�X�l�<��興�CӽՀw���`!^ Ř�`n�gGL^Ɍ�{������'����66Bi��ـ?�������
�{n�f�,�|�N%��T#r�=K�V =���f��e�T��)�Lՠ����w�tn���7�b�>Y���ަ�c�n���� #{�͠��ٻ'VՎ;*]���%$,�;A"�ڤ��`n�gGL^ɟ�`v�����n�M�⦓� �,�x���(�6o���u���3�%�˼���D���%X��v�"`{�A�����H�Y�������x��vȘ�P`l���ꯨI,Q�z�����$��
�j��$��r�gGL_t��"`{aw݉����Gj*�݆���ݱ[�*�n���y;7����u0�=��n�4$06tt���L`�&�����#q(&�R��`|�y��t�>ݶ`z�g$��9��TJ�B�	*�]�`���>ݶa�	DL�>ŀb��>��`�Ґ���)7%��� �׋ �w]`t$�%2����7^��qSI��G;z����}� =���f�at(C�v
բ�q��{O���x�c&^�"�]B'����݂��lul��Y1�Ý�˞׳�����d�j�G�:͵qq�[���� �e.�L
Z��؉�d�m�����V��v�M�*j[*��@�����%���Q�����c��WgrJ�;�Z��h<���C�n��l6#.�����L�b2�6l�ev�O��a�D�:y�u�v��ԛ����'��v�f�r�̄1pS�qu���E�^nO��;dLw(06tt��>�9P�n"���`����vp������1�Ht��*>H�U�1$��r�gGL_t��"`:^ZŔ|%E
�+H`l�����7;������>��m�"PM�Af*`z��0����0;�?>���8���r��s��jzr��	�9�X^jz��Dl�Kh��s�<7��c �0=ܠ������1���ҫ�`�@�+��I����W�����CTU��oxrI����$��{�~H��n��G4�	Dp�7����1�vȘ�P`u�DX�T�w��T�*`z��0	�&��~��������>��n66�)��v�������,��u�tB_�����Z�p��ƍ���:u�91rA5��ϙ�3p�q�q̲.��/�גּ9Ӊ�ٰ�@�_���ŀ};�����m9����J(�$Rn����$b��o�?ϐgt�`����C�R�Y�rI����$�������U�u�'��A(����1\�I��m)m�����%%as2ZKIHK��I��T�8
�ݑ�!G 8���*�� �z��AWEW�^���pEb=
}	%�^��=׋ {��QJ�\Lՠ����3��x��0��`-�vv�ԥ���T����v3 ��I~����6{�V ?7xݹ}!-k�k��v�� �]��Y�8�[0Ɯ�uPz�A,�-�zs�9��6��ŀ};��������w��y��HEPL���`|�y�g;�>ݶ`u�΅	)��O��D�ݑ��n'�{}�`}�8�;w����; �7�A �8ܒ�ߪ��7�`�b�>��X_T$BJ	��QI%u�/ �]U��j���`N�����&Ș�P`J��qs�ݎ�廛&zB�W�ہ&)�0bv��թ��9{K�"������v��_.�s��U�6���l����w���$O�9@�v��/�_�3���9�ŀ};����
n�Wb
��MU��� {�
g��V v�^��:(��D�ah���O7�,��V ?7x�)�}���\�$�(&E�`|�y��_����ޟ���XDD{��T�h�e��.�-�t�sX�=�k<u�v63��Ɯ��;j��H7bv�<�\'\�n���ۮ���=���\]u���ڸaܕM���ur$5��U
�F�S�Ye\�K��&�m��k���[�t�م�n(�)�Vۂ�͑�����	�NL'0m̆���0l��ݱ��
/�r��Y3VHd��ŉ5�$�cO��w��k��pפ�P;�Gb�(`bŭ��c��hs�n�n�ә#������>��ʔ�p��Sq8���ޖ۽u`v���#�K}X �}3!jЮ�V��LwGL	�0=}�މ��+0=��M��($
%I�`w������Ok��7ذ�-UT�ɋ��W7Uk������� �u��>z�X���4
�䜠n; �ޖ���wGL_t����#1Y��$�u�uV:3���v4"��T�/���硇���9E8�RRnK�;u��=;��B�@������*��d�ah���=׋5E
>�Jߡ}����`��`}��V��ԁȑȉW7k �������>�X7ذ��H'*��Sq8�?�UU%�����݋ {���o� �HU�K�X�LwGL	�0=}���`�K�����#i�@���Yـ��V�r%���ϏǮ�;ӵ��l����H(T�^*�����1�M�0;7���C|�/�'N�H��`|�y�	�&oGL	�0;�c±e�����T�� ?7x�^,>�P�^����Ζ��
���E!],I0;dt���ft���`wE�S
jBp I*��{���g�y|�����XDB�ޞ�*�t"�Q4\��vB�	к�d�^��k��C�9(��z���D�Ci��"��<���3�����u`nw]Xk�%D�2��l�, ��x�^,|�,�Z�:!(S!�=� �(�N�rX��s���:[ ��0��"E�@�P�b�T����:[ ��0��f����O�^��V��O�t�#B�R&�X���Ή�����GL�_����G3Aڝn�ݳ9x�۝�hcX�ۋ��W[��8��K�]���c�vF?�~�����l�����b�V��T��+��&oGL�0=3����Ϣ?������T �B��`l���ݜ n�`o{2U�$�j(�RU��=�`����޺��W��;�����yF�2����v�����XͼX����d{wwn��o���묖^wex)Z:�Z��:P6[�=�a8�bE췆�,mm�q�s\���t����&���;:�[�\�KDqe�m��N��܌�Eo�sG#l�j�kawf�T��9�N���))���	;�ev٪z]YV�sFCm1�6r���ۧ��#�$4F�ќ�M��n!�v���sN���2GZ��� 	7v�ɒY�on_�����>�Z�d.z�!�s��[���3:�+���[z�=��7ճ	K��{��o�mu���̍6߿{�`6�`K�X�� ��S�Se*(T�^*`zH��1���3 �kŜ�B��m���T��IV���X��V����DB�z�����'���n���K.i&��$���+U�߯ �߱`���>����m�.�ʌB���`v�t��#��o+ �ޖ����H��B��1�Eoj�y�5�ȭ�H]k�:v:y���\_�{���rܔ6HAQIX����������`no]X�_0�Ti��*T���|�\��DB������X��V��W(ܦB7)��`:&oGL�0=3���eh,��j�������СB��߼��b�>���6g[��mU:�&PU���j��o�(Q�(Q���W�;�����޺�7v~�Q5R!T��:�S�`�oEs��kl鱴��t�-G���l��NE)�GIT��r��o; �ޖ��Ձ��u`no7�(%S�NP7 y�脡D���,�v,�z� �
����Q�WKLގ��p�"��%���ph$�R��I%立���׀}����VZB,J�	*`v���1�N��� ��a��d��ܫ�z� �	$��(Q
�w~�Ͽb�������ϯ}r��JL�����'t���u�7;�_GEk�sK]qԕW5u�u��׋ ~oBIB�/w��w�ä�( Ӏ�N;s^,��X��� �u�~�
dro�*j1�*8����]X.�v%�z[���ŀ��v�� �S*���Z�>�����7��`8�P�T"~ ��߼9$�ݿ�l��wJ��T0	�����0>]���xN�e9IS�*)N(�x��g{P'4v��'6ѣl&�K�`z��`���'_*դ�����0=s�~����W�wzX��SmHA	%X�{�_��Հu��׋?(Q�v��J�!�Jl�ʰ1{����`v�K`zH��˕-#-������� ��x����oDB�UK���=�0RPI�q�%��Z� ��� �^���w�B[	%~"x�Q
��LQ���.���%(P�e RV�Ii,��yNL���`C5�!�
J ��Dn		�$e&A ؒ�zy���m�wm��̚�!���egD��rn|=�ʋ�@����r�UPH#Qt�#3�յR�L��Xs*�\�g������3���!���Ae�쪠Av�v� �m<՜v��Pk�tLQ�mlN���9�N�.��x�ۀ��E�a8����c3��F��u��rn�u��Q��n�ɳ��>���>r�4e�zMt�m�6��\���+�'ֶDخt��VE�t�[��'(�)O�zMY{��2a4����I���������<m�(i�u�`�¢�9��1qg;�,\Hd����)��3�lh6؝یe�SU��3�Fv��SR��uѝl�!�I�4���]Z-m��i-m��ѻ;H�x5ծ�6�m�a�xvMŤ��pR .4�D�k�Nu�n�¤�k m��ft9���,\�p�^�ي��(�uPq��uk���7&���B3cll��	�N���ѻ`�uT�]��ns��O ���ll�[9�v�p�5��ݶ�9�3��yg��t��S�zDE��8�91-�xɭ[�m5i{$��:�j�1���:)u�*=춫�FƮ�j��l�6Ͱ &�rN[Kh	 pI�kKmU�@��tpR;f�UZԻ;4�T�]@@J��s�Z�7-8ԓrʩ��2H��[@ִ�Hp��ڤ�nݸV�weU)����5Ir�Ÿӽ��K3�Nݧ\�m�ؐBշ]<�h�k= �GL�@L
��ҵU�
%�]V�;����֜#Ļ�uKsS�mۡ��U�Rϗ������:�-Xp*�I��痖�v�I�+�nr����z�l=u�͸掶�D�%2���'DĘ�U�K��8��D���%5�MT�
�U��� ��[v�@3]-�v���Mm� �yv٩\��� ��v�9[����pUz\�Gi���o-��2�Jgf��WJg��ݫh3�w[wss}Q*��<��h �C��ɣQH���z�'S������N��L�-ݛv�]�s%�:�A��5��v�m7HXl�m]�q�綜ٹFӝ*GC�F����yk"\ks�p5	�n@ܑoJ��1l�<��D��W�۷���J�[�{\�۬�n��V�����x9P*��Ěv1��TYM�գ�;\]Ι�i�*#������Pq	���ke��zNΫ(�n"��]]�P3�`�Rڮ�{���[�����4�5kJ��;m{a�Q,��urn��b��ی�vn������Zc������ŀ}/]`���!D%��}8 �^NTu���Tr��o; �ޖ����or�ID)����e)W"�e�X��I?&nt������p�
mT��E�r����
"���pwv,�Z��P�J&[}x�z��RC�H�����������wzX�yX.�]�pbt2�Ӯ��rBk��l�P]T�^�+��Wl���S����������"uW\��6�������]���?�(�_Hy�b�<�yr�V�#*�0X��otN}_U}��Scu�� ��ŀ|�\��%
d�k�)�"Pi�pnK������]Xs�V��,{����Q��TR8���Xε� {u�B�P�� ����@�)*�ܫ�{��3w��۝-���WIY��Hŉ�`�2�v�%5�9U�$>z�ѣ�͢߾��~�wn��DT�'(����zX��p��_�}!�Ӏ=��WEJ��դ��:[�GLL�l�z_�~����޸��RC�H��v,�z�%P�Ck]���8�w�Q�H��%8)*���U~Y��V ���7ծp:$�D(U��~��7�)� � �������`n=�`}�0=3��:���]�_!P%K��g�Ӭ�͐4��Ţ��>��2Y�8�*�����v������ܟ�����>缬;zX���JT���SR8���`:�8���k��2��Q�
���Pmʰ3ϼ�[���ܬ������wPh"*"��D�=;���78��,�(�
�}�Vo���O҉�9%������H遳:[ ��:�)eڼ,N��n-׏j�6�{[E� En��Z�n�G�d��Q�$pi�!���V��u`g=�`������+W��(�9e��n��Z�?BS!���k�p������~�H�k�� ����q��׀o��á$�L��b�6y�`�Jʶ�Z.�#1&nIlt���y�����i��:MFS�QIw8ͼX(���}_ 6���79%,M 4`��R��{����a��+��n���FS��(qm�%뎰;���8����]���@v�
��H�	��3�A~?0�p�v�kU���VB.|�ķsl�bG���!:ym��:+lr�����mݖ��Ӳ���C	E\;��Fe�؋���jA�	��ձ��z�3�p5<a	���i�7oA>h��y`]��r�&��,&�Fw6���Z���6��n���A�J��l0��[�(�nt�ǗN�	�9s�����33O��,K��~��S�,KĿ}�w��Kı>�{�'"X�%��{�'�,K�����m�f�K�I��S�,KĿ}�w��Kı>�{�'"X�%��{�'�,K��;�ʜ�bX�'}�;!�&M6I��ws��Kı>�{�'"X�%��{�'�,K��;�ʜ�bX�'sﻜO"X�%��׼�ٗ.��fl�%ͱ9ı,N���q<�bX�'���Ȗ%�bw>����%�bX�}���,KĿ{;ٹ���L̚fM�Ӊ�Kı=��r�"X�%�{���'�,K����؜�bX�'}�|8�D�,K�3����6�[���ȷIf��Pq
[^zճ����fY�m�d�P��bcr����bX�%��߷��Kı>�{�'"X�%�߻�'�,K��;�ʜ�bX�'��釙�m�nl��sw��Kı>�{�'!����]��,Oy��q<�bX�'���T�Kı/�}��yı,K��[���u��wwlND�,K���O"X�%��w;�9ı,K��wx�D�,Kﷻbr%�bX��;sM�d7KM6ff�O"X�%��w;�9ı,K��wx�D�,Kﷻbr%�bX�w���yı,O����ݶ�m�����9ı,K��wx�D�,Kﷻbr%�bX�w���yı,Os�ܩȖ%�bzwz�f�ݺM�̍�+:.���kLN
�6+-u���Zd��H�h��>�~Ou��=�'�ov��Kı<�{���%�bX��s�S�,KĿ}�w��KĻ����]	��3ml1��7���{��w���yı,Os�ܩȖ%�b_�����%�bX�}���,KĿ{;�wM�̙�4�ۙ�Ȗ%�b{���ND�,K����'�,`0TL�ı7>��ND�,K�{�'�,K����/vM̛.�ٓ73r�"X�%���w�'�,K��>��ND�,K���O"X�%��w;�9ı,N��f�Y�.e�7��Kı>ϻ��,K���Ȗ%�b{���ND�,K��O"X�%�~��d˦�\�rn�xx]&S^��f�`�o��6��7��yQ��L����L���Ȗ%�b{���'�,K��;�ʜ�bX�'�}�8�D�,K����9ı,K���n����33N'�,K��;�ʜ���A$N���9�N�?m�H��Ͼ�S�?�@S��D�;��8nYv[��f�nnT�Kı;����Kı>�{�'"X�%�|�{�O"X�%��w;�9ı,O��:l���6M�v���<�bY�_������9ı,K�����<�bX�'���T�K��/�S����0*�$ �Sy����%�bX�N�rM0��e���.m�Ȗ%�b_;��Ȗ%�b{���ND�,K����'�,K����؜�bX�'�9����Ha��)3r3��'M�I:�Y���MDqu�]d:6Nl���Ѕ��w����̮F�Y������{��7���eND�,K����'�,K����؜�bX�%���<�bX�=���������Y=�7���{������'�,K����؜�bX�%���<�bX�'���T�O®TȖ'��?i��n̹�f���'�,K��w�؜�bX�%���<�bX�'���T�Kı/�}��yı,K���θB�i�]���,Kľw��'�,K��;�ʜ�bX�%�ﻼO"X������9ı,K����6d���Mۻ���%�bX��s�S�,KĿ}�w��Kı>�{�'"X�%�|�{�O'���{����)��ԍ�x.s�s���Y*n�2&m,���tT��V F��{�Bs�;c���wMַ:T��8ی�U �v���˴�z��tm�-mN���k��m�n�;HE�;\}�i~u��7�cr��i���b@yܵnWO=y;;���n}^=��M�s�E�ts��Z���\�KT�K*�Rϕ�����z�Kb�"���ܹz�t.�-�73v�g��l�X��[��f�s��T�\P�i�[���ٻC��ı,K����<�bX�'�ov��Kı/��w���&D�,O�n~�9ı,K���з4�4�v]��'�,K����؜�bX�%���<�bX�'���Ȗ%�b]�w��!I
HRB�۠�T]�IV��slND�,K���x�D�,K��v��K�ș����O"X�%����9ı,K���nl��ɗ33wwx�D�,K��w*r%�bX�߾��<�bX�'�ov��Kı/�w���%�bX����.n��e��͹�S�,Kľ��w��Kİ�W�A���m��Kı/߿����Kı=��r�"X�%�������V�9��u��j��O�[S��F":�{���KFa)a�ب�W\����yı,O���Ȗ%�b_;��Ȗ%�b{���ND�,K����'�,KĿ[��.�)�]���,Kľ}���z����P��
PW�X�Q=lL�by���T�Kı/߻�x�D�,Kﷻbr'�eL�b_���lɤ��SM˻���%�bX�g���9ı,K��wx�D��C"dN�m�Ȗ%�b_{���<�bX�'�^�e�n�v�&i&��ND�,���*������x�D�,K�����,Kľ}��Ȗ%�b{���ND�,K���e̙�L�K7f���<�bX�'�ov��Kı/�����%�bX��s�S�,Kľ���ȗ{��7{��ߝ[k����+s�s�[c�X�!���x�<�غ�����{�ώ�a���3I�\�Ȗ%�b^����<�bX�'���T�Kı/�����%�bX�}���,KĽ�t����3-�M̻��O"X�%��w;�9ı,K�~��<�bX�'�ov��Kı/�����'���,O����wJF�Ow��7���{��߿���%�bX�}���,bz��D!¥ Ek(A"�+@��hęJ0!�Z)�) a`p�S"VP%Y$%#@�BT�V%	@�X� �# "ThH0fd1#�²����`ht������1�F4�! 1�����\`�h�@�X��c#ȯ�j�A`D��iRQ��VXBD$U� XT}V����HBC��x�T�Q��X�`�B��0��*J��
# 0}b�qF	�! F|EQ<qS���U}EC����P��809�DT���~�É�Kı>��r�"X�%�~���3K6fd�6fn�<�bX�'�ov��Kı>����yı,Os�ܩȖ%���>�����%�bX���Zg�[�4˻�br%�bX�{��q<�bX�'���T�Kı/~����%�bX�}����7�������hIδ8�mWǟ&ۧkA��65�7N��M�n΍Ek��lf�M7nf�O"X�%��w;�9ı,K߾��<�bX�'�ov��Kı;�{���%�bX�}{�n�]��M�&��ND�,K�ﻼO"X�%���ݱ9ı,N���q<�bX�'���T�Kı/�_�.d�t�if컻�O"X�%���ݱ9ı,N���q<�bX�'���T�Kı/~����'�2%���d�a���3I�\��,K< dO�~����%�bX�g���9ı,K߾��<�bX�'�ov��Kı<ώ�����e�i�73N'�,K��;�ʜ�bX��s�~�'�,K��w�؜�bX�'~�|8�D�,K���Bl9��ܹ��K]�q]������]�#rėK��k0�Q����nXf�"X�%�{�{�O"X�%���ݱ9ı,N���q<�bX�'���T�Kı/��w	r�f���7r��Ȗ%�b}��lNC��k�6%�����É�Kı;����9ı,K߻��y�W*dK���L��t��wwlND�,K�~��yı,Os�ܩȖ%�b_{�w��Kı>�{�'"X�%�{�ݚn�4�6�i�s4�yĳ�`dO��~ʜ�bX�%������%�bX�}���,K����Ȗ%�b}��ɻ�v[�Y7d���9ı,K�{��yı,?��{��byı,N���É�Kı=��r�"X�%�耆Pbp��gge�	o�.�YH[�}Pd�[����&�)�5��ŕ3� ���6���nAv��wO;�F�hw�/�?5D�A��t�N�<g�ã�h8w�����0�ګ�;[d�b�n{�p���of�u�3����D6X�nմ��5����VW��gn����q�'�����E����x����RŻk��`ㆁ��V�[S�qu�ͭk�vs9�ߞ�w�_0���n]Ձٱ;x�t+��l�Z5��\Hd{E�cb����a�[�\Mٹ��'�,K����lND�,K���O"X�%��w;�?�g�2%�b^����yı,N���	�vYfi6˛br%�bX�w��q<�bX�'���T�Kı/{��Ȗ%�b}��lND�,K�������3.d�r]�8�D�,K��w*r%�bX���w��K�2&D�w�؜�bX�'�߿xq<�bX�'�nwI��a��m�f�ܩȖ%�b_���Ȗ%�b}��lND�,K���O"X�%��w;�9ı,K｝�.f�n\ͳvf��<�bX�'�ov��Kİ��G��~��{ı,O��~ʜ�bX�%����<�bX�'��_�`���;�hw7���um������QǇ��{4���e��I+�����֬��,�r%�bX�w���yı,Os�ܩȖ%�b_���Ȗ%�b}��lND�,K�߻7f�4�v�i���q<�bX�'���T�)��1T���QLr&ı/~��O"X�%����9ı,O���q<�bX�'�]:n�]������9ı,K�~��<�bX�'�ov��K�"w�xq<�bX�'��?eND�,K����ᙙ�l�n����yĳ����9ı,N���'�,K��;�ʜ�bX�%��wx�D�,K���L.���6K�br%�bX�w��q<�bX�'���T�Kı/�����%�bX�}��������ow���?t �jv���<��H�����z�e[R���h����k2�w��'9�937wp̹�M�w4�=�bX�'��?eND�,K��wx�D�,Kﷻ`!<��,K�����y�7���ϳ�l7GX[�e���{��,K����y���,N�m�Ȗ%�b~���O"X�%��w;�9�E��,K�ߧ�s4ݹ3&��sw��Kı;���'"X�%��{�'�,pH�T���,ND�~�2�"X�%�w����Kı,���θBݲi�wv��K�����߽8�D�,K�����"X�%�{���'�,K����؜�bX�%�߻wf�4�t��r�i��%�bX��s�S�,K��QB9����ObX�%����9ı,N���q<��oq�����y���"2�ݷ^�F1�vHS75���0y-��-m�f�� m�m&i&��O"X�%�w����Kı>�{�'"X�%��{�'�,K��;�ʜ�bX�%���ap�tٶvf��Ȗ%�b}��lNC�TB9"X����É�Kı>���*r%�bX��}��y�*dK����i��l��l�6��Kı?}���Ȗ%�b{���ND�,K�ﻼO"X�%���ݱ9ı,O3㽙���f\ɦ���8�D�,�VD�g�Ȗ%�b_����yı,O���Ȗ%���*�V���ț����yǍ�7����F*Ʋ7l�������bX��}��yı,?�#���؞D�,K�߿xq<�bX�'���T�Kı?��{�ݷMv�l%˦饫�L�=<��شV����8ynm=][D���{��|��QcR5��~oq��������,K���Ȗ%�b{���ND�,K����'�,Kĳ�ܹ�!�l�e�ݱ9ı,O;��q<�bX�'���T�Kı/�}��yı,O���Ȗ%�b_���wlɤ����33N'�,K��;�ʜ�bX�%�ﻼO"X��/�4؛�����,K�����É�Kı>��ݛ��f�d�&��S�,KĿ}�w��Kı>�{�'"X�%��{�'�,K�Y�>���jr%�bX������2�,�v]��'�,K����؜�bX��~����%�bX�~��jr%�bX����<�bX�'� D��bF @#�l<zn�n��7K��=��CrH�=p�2wKy�t�'H�y��;awg��sr����CN�:3ۮM۱��S�E�jۇ=�5����w^�ꮄ�۷on\e�i��mv8,�LӰs�e �M����T�MMR�*�l=t7T�cg�����$\r+�/ْX8�p�c�ϔ�m���[c��;�|�e9�60��6W�ig=f�k�Xϟ{���|�ŝ�Ѡ��c����^�лx1���j�NkU���e�4���z�F-�>�bX�'{��'�,K�����9ı,K��wx�D�,Kﷱ��7���{���?���4�(������%�bX��s��!��"dK��oȖ%�bw��lND�,K���O %�b{���t�ve�$̛�jr%�bX��}��yı,O���Ȗ%�by��É�Kı=��mND�,K��Ι�v��˙�n���'�,K����؜�bX�'��;8�D�,K��v��K���L���oȖ%�bY��_�l�rɦ]���,K���gȖ%�b{��ڜ�bX�%�ﻼO"X�%���ݱ9ı,N����4ɍ�6�i��ў&�&v���3�������8):��]�I\X�6�MggXu��؟{�'�ı=��mND�,K����'�,K������g�2%�b~��?N'�,K��n��ܴ�6�&i6�ڜ�bX�%��wx�B!��L�b}�s�9ı,N��|8�D�,K��v��Kı/�^����e���wwx�D�,Kﻜ�Ȗ%�bw��É�K�ș�۟�ND�,K��oȖ%�b};��K�]�3K�n�ND�,��߿zq<�bX�'߷?Z��bX�%��wx�D�,�ȝ���'"X�%��t����Kn�ٹ73N'�,K�����9ı,K߾��<�bX�'�w9�,K���Ȗ%�bw;��I�L�#�F]�,�%JƚK;���m��AZ{vqYm��V�(_�{��|.�j�,��.�=���"X�%����'�,K����"r%�bX�����x��=��M�H~�΋�I#m7#NK�����fk�ؖ%��{�'�,K�����9ı,K�~��<��W*dK��uL�h�j��M�YRB�����'�,K��;�ʜ�`
�TB0E`j�:�4�6%��wx�D�,Kﷻbr%�bX������f��I���3N'�,K��;�ʜ�bX�%��wx�D�,Kﷻbr%�`?��b~����Ȗ%�b~�t�����d�ݒn�T�Kı/�����%�bX�y�lO"X�%�߿~��yı,Os�ܩȖ%�b{��ﶘ����-�Ml�N��ͫ&T&�6)V�:��^�ٮZk3Ex}��͋wx�D�,Kﷻbr%�bX�����yı,Os�ܩȖ%�b^��w��Kı>����7a�3K�]��,K����!��,O��~ʜ�bX�%����'�,K����؜���TȖ'����.f�-��f���8�D�,K�����"X�%�{���'�,K����؜�bX�'}�|8�D�,K߶��fͷf\�L͹�S�,K?���3�{�x�D�,K���br%�bX�����yİ?���WÊ��'��?eNG��7�����߇ު�*,jF�{��ŉbX�}���,K���Ȗ%�b{���ND�,K�ﻼO#���oq�~q��F�FX9��ŭ���/3��q�V�e3g<���Q�kk�1�.�e�ݱ9ı,N���q<�bX�'���T�Kı/~����'�2%�bw��lND�,K��s�v��n�&n\�8�D�,K��w*r�șĿ�����%�bX�����,K���Ȗ%�b}��'vI4�%&�wr�"X�%�{���'�,K����؜�c����?~��'�,K��?g�Ȗ%�b_=�u�L�l�,ݗww��Kı>�{�'"X�%����'�,K��;�ʜ�bX�%�~��<�bX�'ӻ�4�M�Y���.�Ȗ%�bw�wÉ�Kı=��r�"X�%�{߻�O"X�%���ݱ9ı,O8���(D#a�XBX0�!X��	HQ�@��� IJH0$@�)��1HB,�`B$�RVV$aډh�%B�J�BP;�E4�1 Ab
�@�,��@P� *8�� Ab0�E��Xb0`P�$B)�,$,	 � �1b�b�0X|O���J_O��˃.4����!�w��#�# �� @@ @b_�-�$A"�`���`LP(�'�@�S�
�$`�`b��$���H�$H�#-eH�! �H �03߽�wth�����ΓX�Ɋ�q׬%��Gn�6������9��[V�v���4��'��uA (V%�]d��s������1��P��^vU��Y���9�:�a�m���c�b;�+-����͂I�Շ��=yճ�>^G�k��̳�N�|�l���6�:�q�Dvbݲ�M.4=q��h�Qs���H�U�;���gd�5	�kd;a5;�]����Nõ��F_4��s�b��]�L%�.7)�8�(.�ݴۭ�<u��en1�����35��p�g��������@V���0��֖K]��'-�s͝�^��WS�Ix��V����%;��	����,H�rjӕ�N�{j׬�s/d�%à=�Ʊ�9�Y�b���6;]�(�Jt��b� j�R���	�� 1�]0�ms����mJ�.z�5�GJ�@�v���fI%��l�ঁ!h�����m���k�N�\v����M�bm��\�)��Js�ǡ�h��c�[�e ���=����=y�I��L�ݸz��\N�E� U5:{n��8,bU���[t��z�Tz⪬�p�7l1������@� ��l�	 p/Qkk��A:-��ˤJyͶ�6�-"��Ŵ�r�C^LK=��$jI+�d�"͂@�ݮ�`6�xճM�Y̆�A�V�\qn��ݞ�N�kt'S�Y`ٴ��qʀ��{e7S�j+R5�y�L�d�U��vC/Z`�fɜ�(�� �s��ڹ�Yy��K�F��ѵ<�3ڶ\>��}צ�\�:�u�'fm%�4�f��� �P��P�ۖ�U&�L�IWGd�y�1�h�6<b��xl觨��hL/_��e�ٕxԚ��j�@
�Hu4*� �UUU`E�e�:�[^]$m�mΒu T@�A�m���R%�����������FE��q#,�p�޲X�W*ݴ���R1���v�nn�wr���?:����
����?!��AT\Ow{�~w��(\�ԝ2�=q�j��z�{F㴜�S;Vk�8�<�l�LYv0&)�V6�qvv-Ƕ_%���qf��W'&q���Ź�K� �o�������B:r���)n�f:��gC�C�6ۆNw�쒹�Un�<�ҽ�,�g �cU���)�zA�Y��Z���F�xa�ǘ{Ok{�j6Ib��@�R�sr�k%9GF2�+s}�wwx�|>��nwb����e{{L�&�ƣ�;�
mѲ0E�z,o��M朻nf�-��f�wO��Kı?g�~ʜ�bX�%�~��<�bX�'�ov��Kı;߻���%�w�����}�: �7l�������,K����yı,O���Ȗ%�bw��É�Kı=��r�"~T����q��?~�U�T[��{��,K��w�؜�bX�'}�|8�D�,K��w*r%�bX��}��yı,K�:t�wLܹrM2��ڜ�bX�'��|8�D�,K��w*r%�bX����<�bX�E&D�y��ND�,K��s�v�4ݸL4ٙ�8�D�,K��w*r%�bX���{�x�ı,K���jr%�bX�w���yı,O���d�͹1���3��s����D��^�sgC�\�T���qst������%�I�狀�u�b_~����%�bX�}��S�,K�����Kı=��r�"X�%�{�s��e�fYf����'�,K����ڜ�������"lK��s�q<�bX�'s�?��"X�%�~���ȟ�TȖ'g����K��4Ͳ�ڜ�bX�'��s��yı,Os�ܩȖ%�b_�����%�bX�}��S�,K�����ff�n�ٻ.l�yĳ�@X�����"X�%�{���'�,K����ڜ�bX�'��;8�D�,K߶���n۳.i&f�ܩȖ%�b_�����%�bX�}��S�,K���gȖ%�b{���ND�,K��{�mͱ#�����ڬ��:'Y.i�� �dV�4ڎ�e�6U�\9��e�����ı,N����,K���gȖ%�bw;���P�DȖ%�{���'�,KĽ��?;�a�K&�.�Ȝ�bX�'��;8�C�B9"X���~ʜ�bX�%����O"X�%����"r%�bX����,�sMۄ�M�����Kı;���ND�,K����'�,~ꮪa"lL��dND�,Kϻ��'�,K���L��ɤ�)7d���9ĳ�@��3����<�bX�'�߹�'"X�%����gȖ%�bw;�ʜ�bX�%�γI�M�awfn��<�bX�'{�l�Ȗ%�a�����'�,K��w;�9ı,K��wx�D��7{�ۗm���<��qs�ׁ3vk-g[Ts�s9rŵ֝z,GＷϏ�[���n�͑<�bX�'��s��yı,N��n'"X�%�~���Ȗ%�bw��Ȝ�bX�'���K�\�m��7e͜O"X�%������?��L�b^�����Kı?~�͑9ı,O;�vq<�bX�'~��nM�n̹�����ND�,K����'�,K��{͑9ı,O;�vq<�bX�'{w��"X�%��{��wM��̹�f����yĳ�!"~��͑9ı,O{���Ȗ%�bw�{*r%�`b �DDm����w��Kı/פ��sft�i���Ȗ%�by�{���%�bX������Kı/����yı,N����,K����=ݹuɛ��2d��j�v���i�v���7c.����\�{u:)��ˉɆi�p�i�34�yı,N��eND�,K����'�,K��{͑9ı,O>�;8�D�,K���٦I�m���n�ʜ�bX�%�ﻼO!��ș����6D�Kı=��~�O"X�%������O쩑,K����XQjʑM�wwy����$.�ˑ9ı,O>�;8�D�,K��ىȖ%�b_~����%�bX�N��Iwar晻�6D�Kı<����yı,N��f'"X�%�}���Ȗ%�b}�y�'"X�%��Ӧ��݆���7e͜O"X�%����br%�bX~�}���'�,K��sdND�,Kϻ��'�,K��_{ݾ��wm�y�;+�Q�-*����@����)�l*Rnsvw���!�u��WV�c�u�.��:�������L�3>�y���,�l�t��.�mW۞�; 5=9���l���{]na$�zPgm�=��BUU٪�(F�mΝ�q�����|mrӯM,a.�Ie���qף:ٷ�K�n���srs�rd�T���^��wt����5&��r�F,�m����R�H�$�;/�(��l��G�.���7l������KĿw����Kı>����,K�����Kı=���ND�,K������s4����Ȗ%�b}�y�'"X�%����gȔ�Ic}��3w��gpt*8:jR	Yk�:`n��6tLؠ�7����r�'R�Mʰ3r��w�{�ف�^�|�ݮ����XJ)Q����v(0;dt���-��o	�l�)&J�Jt�:�N��u�$��3Nr\�ں#l������(-�7��7[(I$�݊�07rK`:&�S(X��a��X��5_/������wӀ���=�l�=�iԥ�Q��J�J�3:q`�����Ł��u`f��s�TpI�Ґ���׀n��}���=�np�s�#��i��$����Ł�g{�W�n�x���`}���$�Jd���+m�0탮U���Lo���f��V��6�.�f�b2��X*�X���H遻v����n�x�䃿����:��7R�M�`wg���'tLؠ��#�w/�%��,�1Q���	�v(3�j��S�
E� E(�jQ��vf��7��8��j�L��A17e]��~���� ��ŀ{����w�f��D���9N"8X��Vc���������+Y��p�fS$�ZO]h޸�+R�u�,=8���Y��"�Ԁ���4�D���1�+ �ؘ�A�6GL�D�@�x�3-b�;�`n��07rK`nt]R9NF��C�9,ΜXws��Ɍ��`��>X���V
�n�����w|��� �����#�"B! H����!#!H� @ �x�A�����!!�C�s�W�(?'㧳��3=�*�*GMԨ6�X��`�]��`kx�P�"#�}���8��$�oin�5]� �VM�VlX:��^^��䶶��@9�î��1ٻf��'��݊t��{&0I�E^*���!bI���05gs���`f�U�)�F��S��l��{&0މ���*AF�:cn!�IV,�v��,ؠ���遽�(��
�w��2�!�n�Lؠ���遻���}*(zJ��_���_��� n�iJQu�:�������Ą:Y�W��.,�v���U�d��g:�
�yE4��-�u���S�WN��:5�rz7n��D4g0 u�1�U&�r�'��v�1��r�����g+�t-j���%�L��� ƂSv��G�s8�q�t)�vJ)���B��܀.�m�U<���יڐ%k�6�2.�B�ϊ݀�Sv�7	�:
�����m�hl���6��q%�k�M�ҎRK:6�����S.���Bk�)R9NF�ܤ�ܜ��Ł�w]X�8���ޖ��=H�8��X����遻�D�݊N���8�GMԨ6�X�8���`v��GL�_]d�WF*�09D������|���興S��ŀg��j�NR�HG$�7:q`{dt���w�`]l�d�VZ�V�9�nCFvd�
�a5��ֶ��V͎�Q�8ise!!']rjNssm��~����ri`����,����R4��v]ӒO{��s�)�C�#
��>��$P`{dt��ː�J�j��P,+`�&lP`n�運����өȣ$Lm�N�`nt���nt���0	%�b̫XX*�X����遷:c ���8�3�����B��ड��JuR	�5���X��"��}��Cgl�GN�6麕ܫo; �ޖ�N,������\� �PI�fk�|��o�z�?�!�
jԄ�ݗWw�=�� �������`@� �0���"B`�$�F��D���1�!1�q�Bz$�F.r':@�V1�@�H$X�#�А�B0�"1[�<
H�G�X��,��
���@�a�@��!1���+
��p�$1`�!V���!#"������O3�N0�U+E����ޜ� 0U�[H��� /"�5E0�*��ʭ E VUe�X4%R%%a@�d	$�
��
$I @�
$(F���#���5@"D��##!A�#(Ap=�: xA��
�����胚�	�?�P�(�"'������_ 3��`wz/���9N"���>���ϫ =�� �;f���R���T�*AIV.�v��ߖ�>��Ł��u`j��P8"��b;3�t���B��hz�[gcZr��ⲯd�Ѕ�7i���L3�m��߿o��A��#���l	�Jĭb�a����&lP`n�遳:[ ݎ�Q2�.�J��7D����� ����ft��"`v�㤰q�n��Pmʰ3����`nt��?�$X��@(�f/��y����e/D�DA)P�H�3�X��P��q��ذ:�8�N�+*����\F���S��6X�n5��/z�LvjI�gN�fv��������A��#���lvD���R���QV�亳 ��ŝ
""dާӀ���7:q����I�MSd��0;�O��7dLؠ�ݑ�{5�B5NPFG�fwKs���,С(��}8o_*���,���^#Lؠ�ݑ�ft��"��_*X���}��)���ٹ��]+ɣstg����\�zI���Q�ݎ���g���Kώ�|t���^�w�`,N���f�%q�e0��6��E-�k�"�]�N�C$�&f�N�V�]&q;s"�ӷm���a��nڤ'T�C�2Q6{p=���lW�7�|���vx���y��J��񎫓{f��v4F�^�}������<K��u�B����u�kp��o�r��.c�m�M��(v�ďD��Kq��'�;s��7��5�Q��ZHq�Q�%5���?�����{��3;���Ӌ ���76麕ܬ���~P�L��u�z��>�x�ݔ�	���T9A$v��,Ό���(��}�ذ�}X��aJfj���bLؠ���遷:c⪿%�ޖw��Jh��c��#���#���vD��\�P/-�ٻ��������fu�.�Sn�d�ًf�X���T���o�����7dLؠ�ݑ�{;%	!e��4�snnrI=���z�Q�
Q� '�T�����NI>�����������$�۔�����쎘s�0� �R+��YB��VZĆ쎘3���s���w�$9"��7R�ە���pВ�����|`�x��:��߮X�[���NA3+����,�h�f�0�3˻Wh��=����'N�vnե~ ���0;b�vGL��������R��bLؠ�ݑ�9�+ ����Sgw���1)Q�9N亳 ��ŀyֹ�\-��������}�;�,�O.�BND�T�JX�1Sft��"`v�쎘�z��F����`����o���n��V.�v��IQ4�IN��t,c��4n7	�vܕ�HqΌ��� (�ќ\���� ��1�)89%��ӋvGL��쉀t��e��a`�.�CvGL��쉁ӗ�wThrEM:n�A�*�՝��7dL���ݑ�{��*�)`��1PbX�7dL���ݑ��RQ
;#�"5B���=����v�	*�D�.˺��<�ـ~P�n�|�����voK�^��tz��Tc��ۺ��yQ:�ƨ����e0��f�Ѕ���bR�Lr�Q8|��u`j��`�����Ł�w�&�jN�)�X{&0N����07���H�C����zX�8�ߪ���]X��vgN� ��1�)8㗀{�ـn�ŀz|�`rJ&}�׀����MGDb	MG!`n�]X��0Iv(0'յ_W(��Z�^]�P��
Q�W�t��� q163�^��u�롕L�I����ֻ�Tݺ����9n�Wb��\L �^��mR�:�=����ƵeU\�ZX��N�}F;\����5Ʃ���ɩ�1��ns�x%
n�NW{m��_�u�6���1��*�3Ss���Gp�9v�	��w��f�/U*�R��ku���C�:��4���(���&z��{�7&��̻�d4�����J9���tvk����{i^����t;9��Ҝ�'!I:T�A7+ �����>��`ntg�%H=}� m�X�R(�*IW`,X�=:&lP`v�t�۝1�zH���(��"�$��ގ��(�3�ϫ =ϯ �w)��f�a��X�ގ�{&0N���'�ޤ�#*4�JRʰ1gs�N����0�*Y��T�ݶ)W�.R�!��ݫj�l�I�l��R�֍���MիPFn�e��m�������v�}�B�Cg{� ���*�U��33K�����{�w�����C�F�DB��çذ�}X�n��]�R���1����7w��Y������t��Iw��J����{&0N����07vt*2��H��ݽ,ΜX��V,�v�n��2����MzmDWX��:q9�8��^s'\�ܽ7ĸ7\P0B��P�I�P�)��������t���1�ztL讥,.Ċ��b�b�06�L`��(05n�*n�*:���`b��`g;�#�$�$�"BH��<��?wb�3_q!Q�PG��>��`nu� ���`~����}X޾��UZ���Ux��Lؠ���t�ٝ-�{w����y�PI:j�H�O�GR��:x�Iږ7
��s�#Y�3��9b��[5�ѥ����z~t�ٝ-�{z&l\X�S�ڎ~JR�*$ܫ9�+�(�"(�}��z��>��X�۲�)�*@U D��zX�8�ߔDDϵ�,z�N }������Q7d�]�rP�D��� ��ŀz^����>N�<��?o$�����m�l2�jň`{z:`læ0oD��m�>�o����K��f��`��K�L[Z�t�^4u�V`�9z7Yl�f*`læ0oD��oGL��ILqPFA�`���܊l��0�آ1U�"��Vb-$��l��0���X��TF ��rԳ{�U����v�oKs��������Uu��y��r�c���N� �y��9$�AQ_�*
���
����
���T��PTW�EAQ_��AQ_�EC��VR"�"��
���������*
���*+����AQ_�E�T��PTW�EAQ_�Eب*+�*+���
�2�����5�
�@���9�>�)�  �     @          P  p�B�P�*�@ �   
  P�	T P         T
HI@  �"�`  �    (�� m��SJbhR����6R�4��R�`�4�}���r}{��eOn}� ������o���/�zy � �K�Ըǡ�t��� �vK�n�i�|P
 b    }�I  �

� 4;��|�@�룎�1�p � ��ӑ���a�`��x�}�k��π�<@$���{tGv�� =� n��A���A�ܻ�^ }� �P  �*�b �}e���H�K;���@R��F��z�jT���϶��|�� �O�C�� j�����W��;�VOG����i{9�>�ʙ�*fkѸ��q��/��A@ ���� 
oz��e\ZR�c����} =v�8����o� l�ϻ�5<O����>�C� =}=���ݔ�t����r��x�p �ceWs�&���{�� ���(H�d :^_iriLm*��&��=9���4
M4i�M (��Ҕ� �Ɣ��JSJ  
)�����)@�K)Ji �h�H�R�ce)J`l�M1JR�iE)�ΔPYf�R� !�4����UC#�����OS  �~=U$�Tɀ  ��U*%Q�� 
����ڕ)P  )%Jh 5<��O���g����?�Qm��n惷n�ATW���Q\UAS������肨��QQX �����?����	 �7���ۇ��9�0u�����G1��*̫�88�K�tgvw��8����<�4���J<<B��:@&�����-�����\�S�`U��K�k�:�xE��ng;��(�C�������Lr�p<�9HA;�2(��|�.z{�,m�!�p����1��;Ry���.$0'A��N���I{9/:�.>G`T�X����j�� s0rێ��]��p�#�˝k7�L�91`g'O��\E8TO:�.p ��.' M> ��Rp ���f>�B�����A�y�9�W�s
�YR�h��@��rC2�4� t ����>X ĉCdh`���"(0.¦�4`���{Y��@X$&3�A�������,tBat���+���a��P�D���`�4�D!���Ii�Ji�0X�b1$4��YB_�}K)��D�0�����6��;YK\�P��]�A��ۙ3�t%E��P��c��C`ƄA���,�*h�X�	c\�����A�C�!�
��*l- �h�0t��%B5����Sa�q0~5��Ɔ!�,+��6F��]���\�oXHH@��$��uӲ�]���²Ąd#!$bI���)p A#BVd���Q`BK��!k�`'�E`	P�D
*E�@()z���C ��8ӏLgrHS4�Ӕ�y�_��M�D�R�,J4�2#U�@M�"@;�`Q��M˚n�i̞���͇���s}�s�ZD��,��x��)�D�6jr�aHy�in��� ��=HDZ��R)x���h�(`Z��j��K��������xN�X������'O�%\nϙg}����E��$8JLH��}א���pX-8h7��f�i�0!@Á)�)������)��[!VM	�i�f�˧2$���ӭ��/7UxE�m>�Ͼ8h�82�i3���i8h#����*��7���[^	x�8�,��ȡP�� K h���&�ƤJ� ��I�t>x��� ��0�h�\80���N]ȴ��Mga��)	L	p!D�!��\�bB�B��.h�0 ��FȔ`U#D�b�jD�l��+�ޒ�"W[*F�4�B}����5ɮ����`X@�+��.i�sSs��R`J�m�'F�w�q���!sN��J̑�yh-�$�0.2e��K���5���_}���1��R@��5���@�.s��(�T��FugJ���,�u7����	���^,��
2B�*Kw�sW|�F�i%H�$�V4]}��>&�a9�����P�̼�xm�g~���t�ŊH��+6��]��X:hA\��چιB����s��
al��!���!1�T�7�e�L�f��������֙7B-H�6�n������Y�,�JJ��&j���B�V�Y͙ĉ
J]p�J,C�^D���!	1RW�1e�ۚar�#�X/MR[��59��a�T)�ni6�I�c��du�ɬ��5��l"a�2R�}�cVBT�2]�@�0$A�+8�,
���)1��5�4p#LX�b��N���M�qHq`S�Q� l �`�K����	�RD�w���m��p�LR)@�T����%2aH�cPeĨD�*B��4��0�%p�	V`4X�(@1"� 	V%L"U� W �T�@"�H�X� �`Ł@�T�S%BE`Q Pc\VH�B#�R-`@ W%@�@#VV	F�A �pM{�jX�F�h�A�@>O�tFb�FB8�c@�j0��`l��=���R�Hi ���!��@�"E)�J��P�#"B�$� B�,!���I�A*1`�b��0�$
� "$R��$�a�$j`�H��jD�@�0ґ�ģ@+�G��2��X�Oe�#�J$p(M�*B����5���� B���@�V����j$
����k@lX�%�-H��D�p�E� ``ģ�*����l�����߽�\5���S�`�SB(bk5Yh�F�VH"Ё�T�F XD!)V�bj� W@D"�#	9&���P$*�hbi�X4��
�M���kv��1�)�t!W2kC�ip��IB[L#H���j�313Q7n@��1�#d#dq�X2�`fP�L֝�j�`@Ԕ4.@ծ$&�pԌ�H&[m��h��j�M!�P��9d����P�I�I�lk��oaM�)��$hб��M�J��4�I!+��@@!��4�n�&4��4ș����k���rKD�B���ۚ7T����ȱV�� �$��3i�pu����5k&�t�h�(f���4i�@�I�w#�����%5��*�i��l	F@��N���B�o7b@��1��Zܘ����"����a��H[J�����X�X0��Z.&�FeɭM������aL7��Z� FF���.�������!�7YjY��R�T,"F@�$C2�ۭk4�ЗD!�@�*iD!Ck��!\T�|
B1I&�z�4�!�Z������@�4bАܠa�ل56Zd�R���L]���!!)��$��P��p���XdY,�e�5���*p���k)������hg��h�!�3>���jܦ�l��9!!.7^�r\���
��&Jp᚜6h%Û&�L�7�\���hB� `@�х��J��]a�6�+�E�<B��(/������ƔE!�RI�P�B��%��0��`Ub�6�f��~)��*����"jZ���
)�BS46�cCF�)���F��H�t���h��R,��r, +hۄj�5���9�����K�oޜ�+�� ��F�[�إq4���Æ��I
b�i����H]�
��B��ˌj��$�l�CidW������ @)�G35�k�ZcLHDa\#sI
1㤅0]$h��hq��CP�L4B᠅0cq��`G ��d$�46�����H�:(���a�jxH�z1(l=w��GV�HA�k�
�f$	��4�@ >G�J� �h� �4 ��D���$	��S+�@�+f��            � m�             $     +tkd��lְ 6�8)Y%�h����UU@��     �Hr�۴�8$]�_5S�	V(�C�*6�WI+m�!#8    �[RM��@ ���m����eZ[�#�	�j��U����@1��È�ݭ��@^�lm*�U��,����� ���������k1N�9�l	 �Gt2l�pkqp�����C UYF�YU��6�@ ��EL\�k��H7]5U��n��]+/p���[r&*�	�a�e25���m�k� � N�W�Z��Z�v�X��J�+���f���蛤)�.�J���b�86�"��T������L�Q&� D�P2�WevPeW�P\v��b8F'f�l�u����SrlɚW����^������mT�nT�Zv� u�u�m&� ��E��ey�X(���x��(�j�s��%�6رv��mH���v�!ʫ@l�ʮ�[uֵ&[բ������� ִ����Y�L#n�^jU�����ϕgQĎ��V��z�$�W�]���d&���RO5ua���.�XM	�5Pe���9���J���	W`(Ԁ�`ݨ�Vմԫ����g+��iY�R�M�i�- �Z���� ��.���Iư�{hs�[N�l<y���U��-oNUy����pv1@Pj6�ѩ񧛜:��D�A���pj����Rph�XR%����J��[9�,A�̹���Ē��[입Ws��U[v1`�+�nn���(iH�9�{/gA4�UV�l�������u*L���h΀C������#uT�]�[u����S���3���U���ķ��ק��m�=$ ��V�w�o}�m�H   �G��� ��M�` ��vͳx�f�x��:�p n��mM���D��m�-�h8$�٢��[�m�     ���  K��ݰ  m�$h�H	��=    �VͶ�i��    m� 6�m�h�d�       m  �i0��N��h��,����V�m�� l 8�!�l�f�ۚ�       ����-��|V�     [d9 l o]��� 9��[G@   �v���       �$     $ m �m����     �ж����Hմ@���%��m�$ 8��p@l  ڶ4Plv�n��鰑�I�m:Ķ�q�Y��V�
�V���IW{M����  t�]��h
�Zh -�oV�M�Ĉ�ڐ@m�v��F� ��m�ޠ ��!:���[����  �� dt��`    ���-��N6�u��� ��4�e`����K.z���m��@ �@��6�&�h��f�@&�Xn�ۭ��zP  �h v�Jm �M� m��um� ]3-I��9���鍶c�b�!m m�@����j����'��   R��  -�l�h  stRD�i�  �$A��,0���U䍹�@j�V2��$�ULn�քNk,m�9t^m�����@�]m :l��a���$ �M4����m����6�.qÃm��� ��%��(��6� 8�K�^ ��2�;   M۴���6A��� NֶsT6݁d�h86��H������D�2̓mÂ�nJ	gM:K��^ѷb@l�l.�i$�޶�ղ�2ջ�#"@p�.��׻i.u� Pت��6�`�T�*����w�8�؆�m����j@F�l=�Z�Bt��غ�v��=�,��t���qKn��������ԫM�\��ꂖ����6s4�*���,�p��U�ぶ�ɶ�@ I ��� p'	�ݔv� 3NY��lI$���ۀm�j8*���:���(�J�� X�H 	 ;m��$h�3�D����H$	-�d������!�-� ���s�A����&�9ש�n�   -���&ٶIf����m�i;u�vC�	� [M�ke��$�GH嵶Ŷ���� t�k&^�9�+(��ʭ,�V�]UP�m�m���lpݶ -�F�S`-�m$�d� m��`8��� �Y-�����Z8m�H{j{}�@ �5�l���[@ $   	�����$ �Y*�  �f�$ ��m��f͛` m� -�p n�۸ �`-�� I���6��a���}� -� $ o ��ۤ� �%6�n��-�hhI� �Rm&�A�m� Xe���    hku�  m u� �   j۶�Ëhm�2��  Y)� [@ 	��%� [V���m�A��	�7m�� � ��     8� $l� 	l �    -��8[@-���� p�6ض��������� $m�  h��x6�m� l ��� ��۶� m��`$� �  �i8�	 ���Ŵ  �� s��  ��8H�l �   $�� l������� @��   lt�� � ��G   ���l-� =_kmo_Kh �mi7d���5� :@ � �[p a��  p8 n��� ���$ ��m۲�mm      [Kh$�m� �` �`�[@�  h �kmm��l p  6��̓��   � �mk ��i�l���n� ��    m�[N  ����[p8 m������mp H�  %.pkX�l�`l m�  6ٶ� �   mi�   l�9%�km�6�`ݶ6�v��	�  �  [@�B� �ۖ��oW��l m   �m�!"A!m6��pp/]~[�v� p �	8ڶ����$�@��qtۀ mċd��-�f�I� 6��.�8۶�l �m�e���q��!�+F��� č��i{]�m�q뢝�ҽ�S/%ո̫K���6ۋ������Z^����X{j|�R�:ۭd����wm: n�u$�+�GV�z�[�k2ۄ�Y=Y�{7_=  KWkn� %�$��ܮ*�݃n�s�q�F�md�v� m�K���YA���@� l)Gn�	zP[\mf�4�ͬ�� �ZRUP*�T�U@m�s�=[/,�U�Uy,s���m��l �$ mm���6���� �6Ͱ 9�� �Se[���(U\]��-Q�K;�{;��}�&�c�P�A�ڬX���%�M{  �m�i�m�kk"I 6� 8��BP�z��j���������E�	 � $�M����]� ��   �n['Ptm��`[I�l [:W[`�  �8 R�6kY�e��L� m 6�  	-��	� 	� �`۷mm�H5P6�H;m�m�  -�իu�ݔH�d�Nۀ   $ ��   G  �    v���bGbI6�m��i06��8Ӕ��`pkz� ��m�m 6Ͱ   �M�`�B�����  pm�m��l��4RY@;m��� �m��L   m�n�.� |V���k�h    6ؓ5^��U��MX���Q�m  �M����6�8 WV1ҭq���yڪ�(Rk]f��f�mm� m�m�A'��^�{ｳ� �AR�]PPH@-��T�m��i���u�n![II%U�J��I�T.fӁ���b�RYUR����y�� �dWgj�U   I�l[V_4�# Ԭ�WT��h��!m ��m���e����ٶF�U6���@%����O}� m��.D���T=�v���Zɗ5�-��֡5�� PT��?���<��?���A�
 	��J�0 1OS_�(�S�K����١���)���E�j�z�&�Fhz �:DM�7��hx�z��E�a！���!���@�|�`!��AN��Q^����PC�A�`�Ax ��o�tb`��ڈ�T�=��{����_(gǃ�+@�\ ��S���@�AQ6�������@�H���~TЈq v
��Q���* |!��P�����%���~ S`�U<��>��>௓� � �b��	�P)"�Sh���zv��8/J�D�Q��C��p�E#��|�~9�RBO�X���$�H�@��,!%����,b/�y:�x5PE�� ��F" � �j�; �Q:�4w�ATW���b���P�0�?��B 73ﵙ��kZֵ�[@� �4ڌF��8ݍ��P*��UZяj��T�<��#w ;�ݣ�y�^c���]�c��X����`'I�օ�Ξ;b�<����Zm��C���0�=.�Fj��7�ԗ-F����ݪ^��nH�]���JEn�wnm�q1�5�e�]81�݃E��b�Pݧ-����YMr��6���fN����p
�ޭ�^��L�L%8Dq,�׮�ij�RP ���V�ksmR��������MіB6�W���]���*�s����3F5UV�&�T���-,��jzNUd�bT��z�{m�'�0@�
M�.��t�h�i�u+@	n��&� �m
ad)&tJ�k��&2Μ � x��"i� \���6��^�U��PH���ѭ��]��Y�nJ[����vۖ�U���	�;XL"��nC�:v���k��Z��<��|0K�:��-���D�6M����1��R�I8Ќ��b�uۨ�a/s]X$�+&�ͻ6� �qˠܡR���Yr�V� {�;`�`�]n����OM��BC��F�S���(�ej�1L��T�tu��y�[HX���-Ht��[Eѷ)-QWK 1�nSP��nF��Q�r�0 &.)Q��U����� 8�V�Gp:��C{ :*�͡�꺨� ��NKl���'
��3R���R0���
��e@��r!А� ��C����v �l&x��^��\��v.;v��l���|��FS�u;�t��'��;M�7*hɶ�[��p@�U�hz`�^.�v.-�H�a� 4]���Q�ڭ�׮�Dfx۱bh��6oE���UyX�b�ڷ*�IZ�Պr6]��T8�<�mŷ�.t�H�2Z� l�j�i:�ı��N�d�2���<p��3J'��Z��i���ط�Ռ +v��lZ"������](�� �j힝�\$Au��5��5�`(�����@�7�	��+  H*$E��AS q v�M �8�N?P =ݷ>ԙua��٫���zV���v������m�ѻN�W;&C��ۊKs���^86m�F�t�mWVݶ�&f�3=���.�-����n��C��0=	٣��U���q��6{6ps�]4P�I�6ݍ�Vwf�Н��AKS�q��GM�iF�49�V�e�&���5�Q��r�	2p�":݋$���I%�d2��	��2�PULU��@� b�Ƅa�E"D�#;ûl��l(&�/n6�n�r��l�{�n������w���{[A$NϻSPI���͇�@���L�bX���oq,Kľ�����e�*��~����{���O�p�
�r&D�;����r%�bX���oq,Kļ���ӑ,K����� �*�ﷸ��{��g��m9ı,ON�x��bX�%������bX�'��ى��%�a��RmWj�d�9f�CD4CI��oq,Kļ���ӑ,K��^�17İ=2'u�s6��bX��7htH�J���l#�%������bX�'��ى��%�b}�wٴ�Kı=;��n%�bX�������ԻH\�����q��O�y[s�=��Om�X��K�\����6�7=j�kZ�}ı,O�}�17ı,O���6��bX�'�}�Mı,K��!�!�}ꛂmn*�t[&�Y���%�b}�wٴ�;���b
1�!��(sb��T{�_�}ľ��X��bX�%��m9ı,Oe�q,K���n�k��PpZնaD4CD4C���bX�%�}�m9ı,Oe�q,K��;�fӑ,K���5�&�\jn�i�h��h��n�#�,K��^�17ı,O���m9ı,K��kq,KĿ}�32hq�ev���D4CD4F�퐍ı,K#���m9ı,K��kq,Kļｭ�"X�%���#�Sk���]k� n-�뭱z��Y{�+�y4��Ia�3�*���%�b}��iȖ%�b_^�X��bX�%�}�m9ı,Oe��CD4CDwn�i�]�WERV��iȖ%�b_^�X��bX�%�}�m9ı,Oe�q,K��;�fӑ02�D�;���p�j�Iu���5�kX��bX�%�}�m9ı,Oe�q,D��@M� B$� ��D=�P7Q=��3iȖ%�b_�}�Mı,F��ѩ78��P�b֭��!�%���bn%�bX�g{��r%�bX�׾�&�X�%�y�{[ND�,C@��'��U'b�+,�b!�"��;�fӑ,Kľ���7ı,K����r%�bX���f&�X�!����������\�N��J�͡�[�V�n��c�*��u9��3���c�;�w��B����൫l�D4CD4C����,Kļｭ�"X�%���bn%�bX�g{��r%�bX��&�36Z�EZ���F"!�!�۷��#�2%��/�f&�X�%����fӑ,Kľ���7ı,K��2I48����p�"!�#c��Mı,K��}�ND�� dL�}{�bn%�bX������K�7��?���9�����{��7���;�fӑ,Kľ���7ı,K����r%�`~v���� ��#�@8)�Oב7��f&�XCD4G{~��j�P��-nK0�"Kľ���7ı,K����r%�bX���f&�X�%��w�ͧ"Y�7����?�ŵ�\�ELN��5����=��Ѐ���Kj+I�B� 82��Ut)mRQm��CD4CD>{v�r%�bX��粦�X�%��w�͇��DȖ%�_~�&�X�%����78��Qb�]��!�!��w=�7ı,O���m9ı,K��kq,KĽ���ӑ,K�}꓂llJӱ[�B1��>�wٴ�Kı/�}�Mı,K�����bX�'��쩸�%�b;�� �Z���֭��!�� ������7ı,K����r%�bX��粦�X�%��w�ͧ"XCD4G��d�e�P��m�b!�,K�����bX���׳�T�Kı;����r%�bX�׾�&�X�%��#!>(e �۽����f^���&�ӹc#�S�Rg����ہ�0�s^���v^:�Yn=��S������]���$6��v�����x��/5���vJ�Е*����9�AvU.�kg���Z���=��#m9�ݙ���Ggb�T�f�Y�9؜s�T�D{k����P�L�<5�OA	0�1.0��+IF�+�
�c��2��O��pfpq9�Ht�bd�̝<��N���nΩZP<��s���g�YDUn
�)U����X�%���~ʛ�bX�'���6��bX�%�﵁�g"dKĹ�ۄq������+N��G3YSq,K��;�fӑ,Kľ���7ı,K����r%�bX��͌�D4CD4Gv�֛Uڅt�ks5�ND�,K�����Kı/;�kiȖ%�b{;�ʛ�bX�'��l�8�h��h�m{E�U]
[c�Ym�b!�!���p�"Z�vbK�}�`Io}���A7�m�
�"�I�U�^�v� ��`�ٛo�q������e0�5���$A���d�l��@������.ݣv�jp�6�`M�1H�W�� ]�0�`v׀w�&��C$���"H��ٝ"~ ��!��ޓR�ė��ى.�{f0  �׽�Y$�c�~np�I�m� ����v� ��0��m�&�R�Ԓ`{�U��V��nـm� �l��AU]���K1%��lė��	  '��� ��� ��^{i��H(�q��Z�����{zw�ӏ3��ЩO<�Gb7J�:�D���9��7 v���0]��[���������5�X�[Y�5C��i�� ����|x����rDI&����>��s��'TE��D��� ����.$�7�$�ޢE5(��K�R<�v� ��0�`�k�;�|n��Gĉ$x۶`�l�5v׀un׀r���\D�E.�����g�}��>~7�mF���v,�̼�{k�� )�I��hЬ��$��}q%WmxV�xwl���i�x� �n9&WmxU���ـ�n~ �]�����n��G%������ݳ 7������Z���WM��%���  I���K���Z��1&��9� ����ē����-
��Yj�������=���j�� .�ܼ67Q��l�d�mmkB�d�n� 0;n�j\��8��.G������i�=�}߯���[��ݳ >�f�����Cr�V%e%xպ�:&""�"�7�, ��� ��^�؛�u)��< ��0�`�k�:�k�7o۱Ȝ�`�� >�f����v� ��0��m�&���jI0�����w�u� ��� ��&c����G��݋�;t8Fw�Z�pY�����C��n�VN���G��[�b{-u�nW�S�e��FUeŗ8��G����n��Յ��C�[=�e����Σ� Kv�n-v�3Н��k��a�.)��	$�U:-�a�>C/nu��ӗVȹ��6�n6�f�ق����Gbq���
�y�rgb��CK�\qYA���L3.Y��-�њ��8�<A���J4�-8t��������ik�q�1<��v�Dv,�fȷQb��R(�~�w�� ��`�l�*� �(��!ȧ��I���ـm� ����v�Qv���s��1�+I`�m`�n���W�o� 7�,vӂO�'��.H�$�5v׀}׵`nـwl�.���u%Ƨ�J�J���w�t�LV�����X���x��w�
7i�E�''eN�Y�qѷn1�u�u�Q�]�����I��r��E"�⑎G��f }�f���s����x��~��E�6
I0���������os���nI���6۶`-�$ۼM	H
6�� ��^�ݯ ;v� �����E F9#�7�ݯ ;v� ���WmxyKơ ��$�R< ��XD��W�ܿ �{� ���xDGw󿟘����DN�x^;Q>x5gj2ڷX�x�+X�a��덪�݇���XqL9�� w}�U�^�ݯ .�%��A7�E�Hŭ[n$��vg�6j���� >� �����K�N9Z�'lė_}�K}� ���w��2������HF�Aȅ�T)�hK��́���}:�
@�F1�_a�d����� ��:�&�7s�`ÀDx &�X��N
~F*?��`��"�?�h��V��םTo4]��QuITTRVZW��&�y����t���uϯ�O���ė�|�}dR�l��H$9���%�}�ρ  Og����  [�k��ϗLDL��DDLz9zʯ!��t=j�Y9�N���v���%͈�-8$�˺f/�7a_�L�)U��www�Tz���x舙�������ߪ�""&)���%�H ��>���Y\�Hܷ�mk���DL���w���F�y`���D�~"����t���ERW��"*�>X��,:j�s��6���Umcq&���RI�vـj｛�}~�rW�<�^�	��~�&����9�'\��LWmx笾_ o�� }���Ԧ���E���������ׄwj�F���t\۴�����nq��N(�� ����nـvـj� ��7��R.$H�#�ݳ >� ��^�ݯ �w�6�lr/ѰRI�yw}��o����x۶`k�	+�M��RI�j� ��׀�f }�f��y"��#��6�� ��׀�f }�f�������E"Q;g��O[3�/;h��<��f��jl��0&�e��-Ѯ�Z�Z	{nKt".�1Ά^��.5�����4�a帠e�Ӻ{뫭N(.ƍptb�a{*�qh8�As�L�C���7+��;ccFu�\µ���Ƹ�r�Լ�pl�-���ŵE�^Ze�vt�ˡ�zr7"��>��49�M�Ӹ����0�4w{��*�@d�][� �g��3���p#���';#��gv:�a��8�P�	H� �_L ���WmxWv�U[X�I��qE'�`ݶ`�k�:���nـ]�����8��J$� ��^�ݯ ;v� ����c���
(�� ��׀v� ������݃|n��"�D�r< ��`ݶ`v׀uwk�>���p�|�fB)E[���6۱fՒ�ٽ!�b���u�-�\I'�#�|���WmxWv���ƒ�w�.�М���IC�;m�|��L�LMP��� ?n��u��e�@�' �n<����Zæf*�o� �{� �n]!".5	 ۋ ;v� ��0]���j�5]u��ۊ7��L ��0����z� >z������i�5��`�w6�|���X1�=�tofKn�s�7I�p��e�9�cW���_��[�<��X۶`�ـ{���	����HF9�o���ݳ 7��Wmx�7��h��(���	'�ﵹ$����;���������;]� �w�1�����h�I��fU��׵`�f���m�&�j@��$�*�^�~����|� ��� om����>y��s��Wc/�� �җY��>�etiGi���[\�4�-�9"�d�$�R$��[|�ݳ >� ��xyGyx�$8�P�	H�ݳ >� ��xWv����n&�Q�NI$��l�*�^�ݯ -�0�A�><q�~J%I`���>��� 7�`}2�/��=����>;��$#$� ��׀v� ���U��]Ӗ>9����rWl�mbܝ�c[ҵkq�'��G8��wF�;al����8�4����ͳ >� �v���^�w�1��I?6�I& }�f��xWv� ۶g�^�M����ҒLU����x�l��l�6��Jr~��D�xWv� ۶`ݶ`t�S�}x���t���]�$U%x�l��l�5]� ��׀}���څ��s�X�q춞�6�m5�>7.��M���f�n����"�9�uu���۳�d���9��vƢ٦��9nή�05��՗p�m��Әы��W���խ�x-@k���v���yܷ<�n^cqd�h��*[H�������.i�x8S<���������K�Ӫ�=�%�7Z!�����9��m��P<��;\t�v7�
Ĕ
-? ��Y&%cv+oLT�'Ru�kg�n��(WK-ul�q�dN ��3$x��m�(�78�@/���5]� ����|���������!�!H�I&��xWv� ۶`ݶg�;���G!$x��x�l��l�5]� ݷ���|�q(�9 m�0��0Wk����x��$�����Ф� >� ���|�V�< ۶`�^����Zn�-�'J�4���t,�L��Nu��Z&g?Ю¿	
�i
��
�|���x�l���0��z:�ڔ��ܳ]}���@�	&e�LL}3|�j�������Q�^5	8�$�R< ۶`ݶa�%W���o��u�'o�EV�ե��m`O]�W���bg�w��,�����T��J�I,i�xWv� ۶`ݶ`7���$���MlV�b �Z�`�zڡf�����e������wOy�,#A�I?o� m�0��0Wk�6ۂ|nE�T��ҲҼ ׭g�b}v��r����:����x��M�@�
I1$��ۉ/=��P��A���������>׼n��m���)$��wϯ ��׀����{� ��=Jr~��D�xWv����|�����x�
NG�C㐱U�m��|ŏ��Ǚ�ch�qG��t�6�{��7��P�Z쩻g�!�@/~߮ �`�`�`�~���؃� � � � �?{�l�lll{���؃� � � � _۫蜮I��e��p �����ߵ��A�A�A�A�~��؃� � � � �;�ٱ�A�A�A�A����؃�� � � ����e3�Y��d&kZ&��lA�lll}���6 �666=���lA�lA�P�������[y�kb �`�` � ��bi��YSV��` A�����~͈<������~��A�����ߵ��A�A�P���>H!��,���"��>D����f�A�������3&f��j��5���f�A������kb �`�`�`~���؃� � � � �?{�lA�lll{���؃� � � � ��q���bB���yWg�^?ﾤ|�n'g;h3۫��Cэ��w}p��ٮ/��E�ֵ��?A�������؃� � � � �?{�lA�lll{�����DH�}�������[y���.f\����u�kb �`�`�`����ٱ�lll{���؃� � � � �~��lA�lllo���[y ���ߵ����sD3Rf�sV�b �`�`�`���f�A������kb �`�� � ߻��� �666>����y�@-��_�J:�B5l��-�yF����kb �`�`�`�~���؃� � � � �?{�lA�ll�}�6 �6667�|~2殳2k&�k5�Y�lA�lllo���[y �~��؃� � � � �;�ٱ�A�A�A�A����؃� � � � ����� |!b���"D�B	Ԉ �W��$d��H�H,%��T:�"��&�����"�1�>bK�h@�q^ ��yyO�$]��#k+8�}	�>��$"�	��{N�]�@��s�$�@�(b�bE���$`����bD��bF$H�bF	 �� �F)-]!qX�B$VDa �����LF(P�),`0#�k��� A�@`�@��r|I!82`D�@	$�R;!��� ��q����BE�F���B�@�g�շZֵ����m�Kh �� ��v�K=T�UV2
>x{4b�'is	�=v�t�W�v
3�;ò�k<����oim�M�ţ_f�4��[ktf��]�ۑ�e��;*kN�x�*7�6NqIOr뮗Em�@R��Ҏ��K!Y��s��GC�b�]�э�����-q�&�:���$��<]6xͬ�s���;H&��\:3ۆ��5�%zݺ��M{m��\��z�Վ�ղ�n�Ye�6:`T*xW������pdQ�< �R�*�m��fr�mt ���`n�p�ڎkٱ���r��)n��nvۭw�|m���r���y
�뮞V���
:�k8�v[C���a6�Il�sv��X���;9�G�R9�A�&��=j�jth��f�`ym�4P����n%�<ERvS�������Fnܖ���l@N"V�4=�.z�V��wP�v�'>v�u	��-��cemTvy�6��i��-.6m��Զݑ�B]׊���=�H�nӮ��.�iuu� ��e�g�n�{3����[�������͵��K�^�����vM
L�9檙�1�zKj�m�"
� u�ڠ ��邪uKl,�Yzt@I��J(�m@��OJ�j|��A�J�[JKHMԨ	��r��Q,gn�^�<�[;puHm �\F� !K���b�V΢j V+����)Tat��ki��-*-�hH+���&�h�[����&��-��W<svq�ܳ�7�wb(\k���#F���e��"�g	A�f����lbp�<ko-�&i��8Fm�AH���q�G\{g����N�(J�v�AmY��Z�͌Ql�� l��t+��YEm �յU��UTx\nD7k-lU������ص�۳ebWݲ�Un�Dڌ.Ƈmb����@�yݶ�l�	���]���4ã\����Ř�*��D��H�!:�ɣ,ˠC��<@�PDґ�.͝U���}$�u4�n�8�kƻk&n�u��mYPkd4ui:O+��x�p7�k/of�ų��ح�PQev����&�z1��͓A6��k������qQ����.q����lt�ح�q�N]';�>���9�bZۄ�˪�Z�tv�5�#��8��]l�v�y���=:�!����[:TvԚ(�Rꈹ#6���P�����F�����ww�;_?YG�Gl���`�`�R��c�-n�:���s4+��5{� �bQ���%�)m
ۄ�$�������ٱ�A�A�A�A�w߳b �`�`�`�}�ߵ��lllo���[y��r˓����K5����f�A�����~͈<���F
A �`�}���[y�kb �`�`�`����ٱ�,ll}���Lə�ZֵeѭY��lA�lllo{�� �6667�����<��?�T� �g���b �`�`�`�����ځ�'���rf~��a�%E$�鈪�{� �{� ���x1Ľo�v�m�&�m���)$�*� ��k�����`ݶ`wn%�ѱ�#2���y�N�.�&)�6�ќI���j�������� g��V�< ۶`ݶ{�o����%V����R��I.�惗����0�mxWv� ��qF�j90��0]��]���ـwix��D�)'	$�*� ��׀v��~K��L�a�?7!�xWv� ��`ݶ`v׀[�J9'8�m
5����S��yr������Q���U�m\��V[��"2D9 ]�0��0
�k�:�����&7P�d� >�k u�w�}_k� {�gDDLEP��m�'�@99RI�yz��]���tH�Kmۉ%���In�]nP0NF�N<��^ [�`ݶ`o{T�����#dN���\ Ϸf��xWv�y�J����E�\<"�pv��F[V�BAvgP�n/<-���c����#�u��k��|��=w�}_k�G����|t]C�d�\JHI&U���Hշ� =ϖ ~���13T}�_]YhE	
ĕ�Z���k������XW>�[xU�څI HJ�J�:f"*��, �{� ���c���1�k��[��.����\+I`�X�=1>^�_�:}����ƺQT8T]_|�/M���A:�d�������T�=9ȡ'>H�����[*���m���������xWv� �l�9���L��=I�.j��UZ���]����z.���, ��,��y�F��IR�)]*�G�����l��yo��[|��	8�q��M���w}�yo����xwl�گ�d�HN5$�]��]���ـvٹ �#B��ޞ���a���$�kFZ���%�m�d+A�U3X����v�{t�H�Y����vQI�7Ie:%�-�W��e�D5X'ۚ8�1n!�8�1���f�nd����6ܛZ��6C��K8iwCə��!�a6�em� <qe�p�tz�u��T1��W��5��V�nm>��N�랦u½����� 2�8j���3�T�r)����ķ]��{��������_��+��v���uv��<��k�6�ԅ�KAw5˵scPn�4��'H�Ь���:�}x �Z��6�3�-��}�`���HrD9 =ֳ�b"*���XV�^�}���|I��q6�'#p��m�]��]����`݀�tO��?HҒLWmxWv� �i0��0l,Q'8>�ډ����xv�`ݶ`v׀}��{���܉!�S�έ�p+=�'Nͱz+���jc����z��jEh�ǀm& }�fWmxWv� ��q(�ě�9	�vُ��o*�^��׀m&{���[��5�5 q�$�<��xWv� �i0��0�b��k��8F9���x�� >���}�_{�'��"���G�m& }�fWmxWv����>ο�}�}��ժ8"Żsv��v-������ln Ł䵩�f�r��[G]-��;���*� ��׀m&���D�9��)$�*�?�$j����0��0]�$�	9�(��]}��I.�급"�!".wv�[����Ԋ&(�$#� >m� ?|��6�n�:b&����s�4�Q�8�MƤ���l�5]� ��׀m& ^Z�J)NN>G�`�g�6�|��-v;q�gb�#A�5��tf�&���/R��q�DԀƤ� �v���^ m���m�ݰ��k��8FI�ݯ 6�L ���U��ߢ*���U�څI HJ�J��p���0�9Ī���5m��;��&7Q�Uj�E�+B��D�f�_���w� ���r|(:W���{��ܓ�����E8��RI�j�^�ݯ 6�\I.wv�K� F��A�*r���#�j�  �kL%��=2ȎՎv��]� !��@'$Q'8I��ID��o� m���m������EQ(�$� ;m& }�f�����^{�������q(�r7"$���0���:fj�����p�u�.���n@�RI�j� ��׀�� >� ��\�F���F)��]�ͱ`�X��� �������?����H�!5�L֎�u�t�gt!�69�m<��uû\�Bܽ�����c��;`��C0��T�����Y�պ���&'7�ƬgW2�g�I��a���u�pͣ�;��s�k\k]���nNI�B�6�귪�ہ�v<n��府I�˳fy9�����#B-\��ڡ�1%�"���q�6����¶�3�@�qQ^\ə3e�r�[��?� ?"<��fyqe�e:��J�H�1n�]c��瘋:��d�vۈ�GNפx��]�9D�,���� >� ��^�ݯ �w�1��4�IrqG	�vـj� ��׀�� ��۩>99#J$������]��3F�p���X�I�r9Q7�ůo� o��`ݶ`�k�;Gh5qD�c�G v�L ���WmxW}�_ȐA>����R8%�m��h�L�Rz]�{>֞���J����-��n�t�Ӂ"R@���0]��]����:��E��r G�L��ٞ��
 ���8��{1$���0��3������j(A�F)��� 5�k����XV�^���s�IBD9 m�� ������=�qk��Z�ĘߑƓ�.N�0��0s�}������\����5ĉ>H��(�#`�N�	����c,��Nu��p	V�a�U�h�����V�^�}��[v�11�~��=��yR��P�*�Uv� �����\��l�*� �؝BQ)�llr< �k��m�.��Dȑ���d6:Pa��S��5��,Eޘ���@с��]h����p\ �"��!a[J����!đ�ȃH�"8�TJ)���(`�u"n
�� ����X)�D�� �u��Dx ��4����lė���Ē���'i��) ��`y.�0-���ݯ 6���u^E��'���2I0
�k�=�o�����m��߿�ߝ̖Nz+n!"��j5�m�0,���v8���yͦ��-��?%��$b����x��0��?�ϐyo���{���R@�(G�ms >� �����^$Z�Ęߑ�ۄ\�#�`wޘ]������x}�9�ovmԟ��#JI0
�׀uwk��\����cvـ}�yb�NNH�!Iǀuwk��\��l�*� ��ȣ�"!�H�����m��|Ŏ�q=���m�qG�$:������j%!��ӑ��\��l�*� ��׀���ě�$i�(��m�]��]��m�`[Kȸ���rFI&WmxWv� �k��m���pN��$b��]��m�`ݶ`v׀nۃ|nr) I#����yw{��:�����w�\l�ē1B������*���������f���X1�Ɉ�`�h���F�ڬ&Wq�z.kI���m�mgr/Kq���
����vΌe�Y9��cTa��K�mzR��m�Wj_��o��W�y��`5ә,mm��/sqc9���eN�9�Fٴ g�x�p e;���ٺꂹq���q�v.tOY5��y�v��gE\��a�JA	��:���{D�Ic�Χ���S	�\? n�����ᬖSY55�MS9S��x���nxO�q���6�Ho���,>�S�x^7�ۄ\�#�x��L�����x��0��m��qD�HҒL�����x��0��0]�% H�!Mǀuwk����vـU�^ݱ:��R6�M9 m�� ��������x{yX�I�H�G��l�*� ��׀ms ���GSLD�@$�5��$$@����p��:�������8z&�iʨ�A-�*��mĖ���Iu�k����vـ}݇�P\����K�f�_��ވ��" mQ�m���{�L����po��E$	��$x��0��0
�k�:�����Ln���8�'�Ļ��*� �wT �^�۩D���JI0�j�:���v�0��0w�}�Q��#\���"��5���{[8-8x��T9���ќ�6��f݋�B�䌎r.D��[|��k��m�׵`��J%8��I1���k��m�׵`]��{��N7(�[d�;,��\��ė�{^(	1����".Da�GϾk�^ v�s �^�8����I&��XWv� ��� }�f�vUAr\r8���xݵ� ���kڰx��S��>)�8��Ck�r�X{��NN+m��݆�.���`��	�l���$��}��I�m�׵`]���x&7Q��s��q� ���kڰ��~���s ��6�(5��RI�m{V�ݯ ;���vـj��(���Rq�D���׷� 6��`ݶ`?�$�&���x��Y�7[�GDI1���k��m�׵`]���~w��~]NF�:���s����Y�ӛN�B���O�>x[�k���ၺ���9�vـm{V�ݯ߹���y� �|��q� $RI0�j�:���v�0��0�a��X�9��"q`��0�k��v�kڰ�po��H��8ܓ ;���wl�6�� ;ݳ 귂cu�I�	�8� }�f��X���ܒ}�{5�'N��8���㻟���r;v�g��nu�C!s��=h냘��<P`8���oX�q�<�׷X;8�6ɰ��s�-,��'�T.3�b�Rt��z����k!����/|]Iq�]]��v���\�nK�nN�b�0�P��	Y�k)��nt丩]=�9��	&u�����L��V�9w�ϥ�]�gF��C��Rf����)��A��kc���/w����q�[�w����HxJgv�:�荂d�7��6Ҏv��"��s�����v�d�J^�w� ;ݳ ;���vـo5��Qb�J+��Iw�۟� 6���9��z`^ՀwlN�(��j1��0�k��m�׵`��0{��N$�$rD��`��0�j���`{�m�����\k�jC�$RI0�j���`v�0������>i� �4�����m�y^5�8��e΄6B�oT��s�Yf|N즠�8��"�|ݾ�ݵ� ��f��X��M���S�I0�v\��A� I�Ľ�ۉ.l�x�\�ـu[�1����Bp�9�wl�6�� >�ـ�\�/;�n���m)$�6�� >�ـ�\���`v��C��R�q� w�f wms >� �����s�^��Jy�:pV�:�^Nv�c3�f@�=C�]2#!nY�9j�m����0��0�j��l���8���G�9�vـm{V w�f wms ;�R�\p�R9"�I�k�u��ְ艅30N�%T�����w�����69ȤX�v������kX5׽׀7݅�]����8��`��`��0
�k���`v�˃q����ɄR��1n�ݽ��ۘ �c�����=�S�����v���#�|ݾ�]��{�`��`��۩D�FҒL�����0V�0��0�UM��#��7 w�f��&�H��� ��y��)X�M�7ĸԓ�QN��, �{� ����*"#f$ �_ @����n$�;��r�-JT�$R�� ~���t�u�u� �|�V�0�Ͱ��%'C�ͭ>���`���eꩣ��\���Ev|�/����\j@	�L�����0V�<i.��$��'��B	-rY�}�gL�EP뻒���`�n��po��H��S��`��`ݭa�311Uս׀����
��ЋJ�� V����EW�ܰ�� ��k�13ﻒ�m�*���UЈWiI&Wmx���l��m��|hW�������%�$$� �G���(+�`�0!�.�EЛ������ �DI�%�q-�qC$��Ăc�D�TJ�!���@a�<��My$�!��F1	�5�e�l�b� 4�Jq�@���Q� � JlF�0&Eg3>մ $���m�h����J�U[�+ <��Wf�K2��wDv 7j-�VY�dQt�!e�B*�ra�P텍Ӹ�n�zǞ��lp��z��Y�M�ڑ�6��0�r��Z�.��ڃ��ckwih��� �9B���¾��xt�{�WtZ1�crvv�v���5ͮ_E.�f�< q+tm�=���{X��,	��s�H��I���ٳ ހ���U/-@cR�`n�[D��Ηn� J�Ȉq�x4G,@m�!*ԁ�Baajt� �nM�I�\3 ��ƙ�2�G9FY6�#�O���,lY'�psI�;z�ڪyZ���luB���������-	�p@h bs��Q���+�of�Ȱ�!*A�s����vʓ��lk`�Jn�xݦ3��ꠘ�M��o1���Kmk	���i\�M�o1]^��6{jc��;�9� 1U��ڑ箛f���26�Y1ve���h7Z��F�aq;���w�K�h��f�Vz�Y';<]!��w77@B��3�����s�K��=�G�<��mjx6]�"X�;I��l�sn�fNH�Q�#��'"����U����U3a@���#YW3�(���ʫK�2pV)�P�Ep��.�R�<�H/����:EQ�by�^�<�[tn9 ��Mk9�2uB^emSUJ��p:����t�ҷmH�u���Ԁ���-(�ڸ�;i{p�ʯ6�Z�i��e�a�8��rO;@Q����>�C���,;5������٩��n6�r9�c&[h�6��f7�gzx<�	�����8)��Od�v-�zk���Y���gjx��56�Y�}R�!l&����Ԓ��,��B�o
�U�uX�ې����j�kih�Mssr�ŕ--��BId��*���-��NS�S�mmɉ5���u.w0�i�bl�9�Z�;M�iUZ^Ѱr��6�5��e2�S�qM
)�2UN��ުqDP�#��)�zT> /�|pi�՚�Z�.����Yc�m*ܔ5�U�<a�ѻ�x�g�uk���{nps�����8��V���cJ�ζ�형�Pp�kv�9�tN�,mY$�w�u���tJm��h���8@��;�n��av0�����9@�شmӝJ�6W0���5:��g�(터��5��l�u�p��N�5�x���֛.�S��ү��MV���([�X�n��T1��v|�۞ͳ��k�ϳn��an֘Kb�B����٣������{��{ݾ~>I��!8�M��{ޘ�l��m��L�D����^ �¿YT��.ՔT7$�5[d��l�*� ;ݳ=�� K�|>��ܴ)l����Iw�}0
�k��l�5[d�5m��\rT]$ �$��陈���k_^��K�b*��,u��:�ܡX�#� ��^��& v�]�����o_�k/kem�ٰ�
Z�=t���-X�lIh9�uۓ��j�{�*�/-�7���/���0�l�*� ��^�o��#�~s�#�`nٙ���C��t /�埮����}}�ٹV�3��/5�	��h�#jI&���5v׀j�ɀ� ;�T�q��H�n<���U�L �m�]���'P�NA�8��#�5[d��ـU�^ }�fwjM>��Z���"S�:�޲v6���:���B ���:K�
�U4�V w�fWmx�m���*��& o������%k�ۉ-}ݙ� ����� /��0��0���L��Yk��I.wv�I{we���O�˄� �����Z��LIo���Qbs�8��`y+�y� ݾ�]��ݶ`��Ln�9'��8��`{�`v׀vـms 7�-i^���ӕ72t<��������1�v��M�<����^콕`D��I�����q���wo8�kf�m���y��[�k��%�[Z�9-��m󻷜m��vK���{��m��m��$$o�}�|�u�X���r��6��o�\m���m��D��o��m��}��mzh�ܭ�kv�e�%��o���q���ܶ�y���r���"�� 8*?����zK���>�Z�kڒV�m��m��m��m󻷜m���%��o���q�
�ܝ�����2SWZ�拚�P��R�x-���b��A�� ��;��SU�/��+�'�rAȤ�u$����>�$���16��}��m���n6�{�jlYERW-����m���\� �kow�לm����q���wo8�z���Z��Ģ�e��m���o8�m�v�o�#��󍶾�}%��z;|�kq��;-��m���q���wo8�kf�$����~�@��������W�����mlݒ�m���o8�m��n6��>ʾ�U�ֵ	5�L3W5�k�ֱ�أ`݇iL�^�mŤ��#�%ɜ�,���Yz�ɣj��Y@��4��4�f㝜]�r�%[�d2F��� \#Ŵ4umٍ��9�m�6��`�ۘ%1�]e������T�nHmb��蒞��<]���x<(
��xX��H��1)���g&�*N�x��Q��J��zu���rVL�!��g��^����w�i�f��3.&�qW'3a�,�Y�װQ�,�z��
L�v,@蕶�B�.'$�I#]�sI.�l��K�d����?������ o���p0U"�R�m���m�?H���n6�}��^q�ߏ��o���*�����9��m��V�߷�q���wo8�$O��m���m�o��쉈�G$���&I���q���~��m���o8�m��n6�wv�A�A�9"�JI��$W���$�$�=�����߷�q���wo8�k�y7�	0f	�
�8�k��s�}����5ns�[��]ѓ��7��9cN��e�@����r�m��ַm���{_�� ��@o���-������W��2zj�q�����L�����q��g�K���{���d�_�|�t;R�Z%�[n6�}��^q���l�m���y��o�ۈ>m]��T�UҲ������3�g7���`� >� �w��8�IRJե����ְ�������wޘ�kx��U�D��j9�\�CfT�(,�a�/Ηm���/l���螭�Ȇ��L��	�$� /m��m�v��DLO�u��>��UyV�����MɀvـZ�o ;ݳ /ͬ���Ǣbn���*�ji��I,޿z� >�Z���f,���舙��V�� 6���	��F��#Ao�5[�� v�, ��k nۻ�|��m�2F~���{l�=��wޟ�?y� �v��n�B6����#@�/b^�ۥ�e�:��TN�ֱL�M��RT�.�Ԝ@���|���{$��ַ�����z`�
y�EMN]UEZK nۻ�艉������K�ݹ� G�퟇�ܮ�k���H� [���� ����kx��^5��q�&�rI0=Ľ������nI�g���:
Db��@W��9���\��c�ȪYk��I.vـZ�o ;ݳ /m����e�q	�8�8��K�;vi98m����u<��u�Kzm���)���{$������0���ϐ�z`ޜ�#r~���7��ـ�� ����n�=13��O����U�VJ�J�X��, ��kDLMWu�]����;lu6��$$�Dܘ�w}�w_u� }���阘�����X�U.��Uڋ�UAi,�n� ���}������ͬϦf6�����Y���in�dN��[ca��yI�Q���֧@9� �}��eN��-�@;��ΐ�Ηfr��]K��t�ql�bj.�+h2l8���ɒ�����ۧqX4ح�r��u��\�و-�u�<��6�J�{`�ɈKrm;���
�i�׳���jد4&5jKc����Na�^ ;ny�,��^�����:#���,Y"Muvxt���j3][�6�Y�O���c���qup]p15�)8���}0�ـv���y���7�=Ƹ�N1�ӎI& ^ֳ�3Tor�;��� >�Z�?}��ƌq�C�E��m������0�ـ�RPs�)�)Ƥ������0�ف��wޘ�����?H�G��l�ݳ >� ��o �9`�%�E�<9�S;�4	km��ơ���q���h���p��%K��6�q��(��|��m��k����m�~Q���FI�]\ֵ�$�����E �AP9�fb?�"3�}w�>��k=TotO�J&�$lK��`�o ;ݳD�U�� }�� {m�U���V�+JĒ� ��k �� ~���艉�D��{;���z.��UұV�$� ?���_or��|� >�Z�;��?{�����։Ȧ�%�tA�3������s�����\=N�s0����r}��0�NG"rN�m���׶< �v� ��0��(9�I�)Ƥ�׭^t��U���� ~���k�1:�?H��x��{�a�ߩ��,$�RP��I��I+I��e)B)j֔�	eal�Dv(@BW�a��E�� �h�T�ƨC� ?.�iqC�� P��X��,		�� �$	!$d��$��"�$$bK
�bBB)
��"1bĄ�`��,�# @�,(F2F$��B��2l� BD�$�I²�D��N�p�� �AP!���M���S:"��B��8+�_'NQ��`�lx�^�M�)"k�qƒ��D�EWk�or�5޵x���ݱ�$8E �rL ����1����gy_��� ?����c����K�)�3��
�"!��:�Lfz��J��x�.�L��$-j\����z���kX �ֺ&b'���,���'�H��$x��{�`�X��U�11A�t]EڧPi�$� .�L ���{e��{��wCbE��B�-rۉ|LD�W�ܰ��V }����\D��3A� �VI���\���K+Q�8ԓ ��b��l��ـu��zwEP�WI_׋#)"�E%Q�C��n�zM���� /���q���N�#���w�a���R��U$�@;���~ְ�ͬ{e� ���	�EM�8��kY�5A��,�.U�}�g�EQ���F��\p�ĢrL �_L{e��s�}�o��Tt���"j�-$�=3O{9V =�X�kX�8���`���JI$qE�`���=1�����`�MV?*�X�=�j[���茸f���L�u��7c���.�\�,��v�I�v}��:j��܆N'�HNYQ�����F����Nݚ�{D��H�5����b�dՍ�w��\�yp��	���3��(��\��hW�w=.��r���Cn�bT�)�Þtv�=��fB{<�vK��!ïo��*�][a�4l��Wm.��x�W>����V���s̓;<skO���k��c��OC������^]�Jx�����}��慹�e$���� >z��4�z'� ��`�{�q�M�rr9�`nـo�5X�6�~ֳ�c�v}�ը�V��T�I,���`����Z����7�
��`�ґB
H��%wޘ���۶`�)�w�{�]�)!Y�j�X�m`1��~��� 7�� ���W"���D��m�� �kL�ٌ0�P9�Q��&��C�-�i���	J&��ݳ ��X��|�������Q7!#i.95��;����}!�$�'!�M*'?�8t=�0����ـ^�A'�9$M�ۑ`{l���=���F�0��, �v���4�㉧�L ����m`��蘘���X7�T\]b�!"ҥi`�6�D>]��w�`�� C�#X��(Uݢܕ�=	��V6�z2�n��\����:��:�D�B#�DrH�� ��X޶�[k�3����X�P]�_���Dq`{l��� �m�׺�����|ݪ�*�YmĒ�{� ;�fKk�`{l�>��TiҊ�BV��]���3[�� }}Հ���_{� �yG�qƚ��4.7�5�u�|��m� �������������Wm1�ꎧ���n�pmGk�9 ��u a��N����u?}�0L�nD����L �l��ـmv� �v���4��qI$��� ����۬ ���zfbb��}���B5H9r`�0�Հ� 6�0��N��9'�`���m`���5;�Lt�1N��T �9����}�D�.~�nO��q`{l��� �m��j�=���g����$ph�v:0��/3�c������Hx�䜙�9Їr<
�ZB-Z����� >���k��&?P���;�?(�S���E��0�l�6�V om��ٝ��"ֹZ\���p�Հ�p��0nـ^�A'�H7"JE��� �l��f�ڰ�iX��I��r)$��ـv�k�`� �~�}I�QE�F���Hse�皹�G��	�	A���-ɹ�!%�K;��^�uc�дavZU�%m�U!�����:�\F�t]fU�Ί�gY�����&c�eΧHr�w:N^�7b���W����9���YgU�j��ہ�r�n���j9]Am����8z�=bTU</At���Tun��nFB��y;An�y���+s���N]а_�w�����w�v��E`nX"y"���k]lWb:��5l	�=��՗��SU��O�ps����Q$#���� ��X{l��� ���Ӽ��6I�ܘ�j��k 5��3T>�YW��ҕWQJ�`or�m�=3G7� �~��;��ětR���9&�"'�1}�y`���v�`���}׮��S���D�nL ��`]� /m��ـw��n4ӄ�F��hk������4�+��$3��>B7�6����+�wJ��H�v	$��~�`� 6�0�ـ^�A'n)v�$��*��kD���D]�.���mv� ��+i79RI0m� ;v�k�`�ـ^튨���+�BBHI,L�zf&.߻� ������ 6��u	�x9%�v%�,]��11����~����X�ְ�m�S�..�����W�;8��s���ʡ�vM[�5��{,�2v-���LNI�Ț�/�.�� 6�۶`^Հw����tN�#�9 kֳ�1A��`��`���>�֬m���H�Q9& v���]�'��4S�� 8b���������z`�7E�HB0\rI�m{V om��l�ݳ ��ƜQ�(��%"�� �?s���""b�����y`�]`��Ҳ���%t���$6HZ���
`6�km�Ԝy{a,]��vg�ٴ���ڪ�m���� |��]뮙�����v���3����I��f��X�6�^�������aWW�\$��J)ZX�}X�6���MP����� ۳�bt"N.D�q`�ـ�}��'�ﵹ:��`�~ %��~�ⷉ��7���I�v� ��0�j�� ��D�!:]�U�9�Σ�4iP�\YK��J��.L�M���Y�+2%õD���~�?���mw��~mt�����or��Qh���Lkڰ{l��f ��۟m}�_�n+c��D���x���L ۶`nـZ�� ��+*-��IBI,DLMWs��,��X������X��]E�IU���I�v�׵`� -ﵹ&ǚ��JF��I)B�Eo��@Բµ��A2H�6�m��i]���:����;A0-�|B��I��6�
����2/v:CH:���4��*� ��mP�w����__^�� ����`-���K(:mjnͶ���]W��D�J�P^x�H�8���	Ŷ�3�h�jx�kn,�KmՌ�ڳal�P�[�c� �Sm�:�X��A��^s� �fۍk����M��t�m�;e��吚��	�w����ykƊ'���[��%-��mvZ����u������+�%v�p��Ծ�ܽ/`%q�q��V��u�i�m=����H�vj���k�` �U@Uk�`�J�[�-�J�Z��UWc�x�[!'I.X*�۩`���tT�l��2�m@�M�|[-6�8�#^<��u��0�wc[�Lm����Ѱ��O ��Vĉa�-Li<m;Kj�-���ś�(`P��`�`�6���W[�Uʶ��瑪Bjx��C��G�[rS�"�T,�sY�8]tNn��i�x�����-1�Cg`��;6z�a�ٸ��l��n<m���G����@l�@��݅��j�ΐ6k�U[���L�f��\=�s�Y�k����4�kֆŎ[V/c����mk0$lԆ�ѭ#��9��d���]�Hr��[��J�n�m��mWjB�����W�[j���ۇETͅW'E�ZW3���c �+�2v�eƝF�V��g�j���()v���f�Z'[z�kt�HP�\a` ��r����P����"Ԫ�8Q�HX[w6�!�R��Н�[��B�vd�R+j�]���/5�ZA��_�X��E��q<N�c�ܶ�.8����&Dϱ��k�3͹�]������#�16���k�Im��p�\N�uW)5k4�%�td��gc���.�@ԑ�g���H��:��&���@6!�ɕ׶��W���bq�r��U�*�]tӄ�pC�+i�v"J+�g ����\l��"����Jt���l�%6É���vKfy\�=	��G]Lc`27#S-���~�߫�>DN]1D_m�)�3�`
��!�v:*E
'ʃ�����ߣ/V]�[�;�z�]�l�jK��9^������b�
�땴�v;����ޞz@�r�z���������n3k�V�0Z��㆛�:�[y ���r"�샜8�e�u۴n�:��XX�^8 �<m�]�ِ��x1�0�;;���tm"����l�k7 �u�ն����jՕ���2p��G��e5�х���%̆�D�I�B۽Ul�W�(�vtl㮁;O;r{I�˭���Ip�<�kgS���%�:��9���|w�����������@s|��pLO�qr&�X{l�v� {�`޺Έ����b�����Z�6GrL ��� ]�0^Հ�����ں-A`��J�%�陉���`��������LL�w>X�+�"�`�$� ��X�����z�`nـ{�ۉ�̊)�1�N>�黥�6.�.+uF�x8nu�{�-��;'k����w�&!&H�'�#��@=�� [�`�Z���~��Հ�����\^�55u�Zֵ�$���l_ʀ�`��`��� ߛY蘈��>o��,�"p�$$��`��`�� 7�� �l��A4�"���Qɀ7z� 7�� 7�`tDD�Uo>X��~���4���� -�0�`޺�=�B�렂��\,���bkv�-m�v�ԸQ�:M�8���'������w��r݅>��156������ >z� ��鈈�@=�X�GRhs�$�i�0�l�-{V o[X ޵����7�]�H�J+����K �Հ�k����H� �&"*?~���0{�`l*#j��r��� ߛX ޵�=k�3����X�x�*-�*T�$���� ��0^Հ�f hw]�ok�<<��$�tA�2�kx��6K���A���筝������k�{Jrq�I���L׵`�ـ���&��RDqNI���j�� -�0�l�7�q.4�4�\��G o[X ޵����|��}X�_lwT�)���� -�0�l�-{V%����۳6�K}�둩B���N7$�ݳ ��X��`���߷�߉x�B��Ig�l+<����/4��z9�х\�x�II�,us���`�V om�m� ;v��¡26�q$�E��f{����� o>Xv�gLD�PC|u���	+T�$����u�:fb*������L��3�NC�B90=Ľo��?y`� -�`{��t$Q$>I�ܘ�Հ{��ޟ {���ܒ{���$�D��@O}���G����mF�ۍ��]�����T���hD��qzx��r�q���8b,�&��s�*VՐ�VȺ��F5��iԯV`��o���F��K��]�J�h�!�k���-�$��.�Sk)F�4!;h�Mmv�S\kNK�����0P3,hܧ�8��m��K�����mlT��0���r��Q@�����v�	u�����sx������Y�Qش9�v�פ0m��A����\F��C�{f�f�LN"�r1�_ z�L �ـv��j�;�tj�㟙QȰ�k �Xw�����EQ���mpdr9Mɀ�� �ڰ�ـ�m��A�D��$�$��j��f [�`ݳ ��X�S�8$�E����޾� z�L׵`�o/�S�@�
!��D�<uu�pܹm�1ׄ��EB�\]jo&ɧs�9Ѝ/d�)���I??����$��m��j��f����E'!���X �Z�31�f!#��X뾘nـ�iѨF��'r`�� /m�nـv�z��Ȥ��iG ^�0ݳ .��j�;���6�N9���� -�0�ـZ�� ��`�߳����gK�f�/`U�f���lRY�iŊ�덵a����ٹ�22L ��`�� /m�nـv��"�II0^՞�o�0޾�wl�-�T&F��$�T�`����X\�?A1<� ���r`��, ��V.89��I�$�nـv�׵`� �v�L�$s��BI0�ـZ�� ��`�f r���"J"n�%v�BD)k Pv�z��c�I9v��v����:�Ji���q�&kڰ�ـ�wl�7�q&7QȤ��iG ^�3�$� .���{��	���	���e1Y]��I-߾��.��j��f{�T��8�
��I`t��EW7� �Հ�� �=I���"�PD�}ϱ�� ۱:��8�bH�I�7z� ͬ oZ��������8�ܠDj'��z:�=�ܞ�[���F��vձ��#��G�����rP-*�_ y�� ְ7z� 9v���qG$rr9& [�`ݳ ��X{l�~�Gm�4�$�r��I��� ��X{l�v� �tN��$H��iɀZ�� 6��k�f*��,�*�.��U$�c�� om�nـv�׵`���Ur%8��S᭞ˣ/n-l�y��5����n� ڳb��̪�,%O/!l���u�m�l-�1���n>�գ4h�Gg7Xkn�*��;�sV�7��R]���[��{y)��i:�A�c�.ZP�p<bAR�c<%D/�k�<�g��n��p�2�FE�u��n��G!:-�\4\T(����U;���w��������OFQmM��N�,�nn1<�D�I��]Lp�NL�Nv�;��)C7�12X��`�k n�����DD�}`y�L��/��jqH6�r'$�ݳ ��X��`�f��u&7�qҲ��I,��X�6���bbf"����� {�� ���L��5"I�� /m�nـu]� ��Xͷ�ʋE��I]Z�i, oZ�=3蘈������_z��X�e:a-K�.�\�D�D)C؈뭂�z�h̢�=���pMՍf&�Hk�ךǲO���^k�`{l�v� �tN�+�Kf�5%�f��w�pU(�MS��h>Jp�k�PP>�gr��, ��Y陘��Ue�QI(�Z��U��X �k���>��{��X���6�N9����ߢ=33w�{� 7����� 7u��b����m��Mɀ[fk�`�ـ�0�����@�N$Bn��cL�6�ONqŬ-t
� @�n��,�2������?C�Y{\���W�m��?��ݳ -�`�l�-{[I�8���rD���ـ�0�`���y�ֽ�}S��nZ��n ww, ���~��6LQUC"��I7���A>�A�$�&$�B �4y$)B��[N#�)�	qBB|D�#�!@H��H���]m �	��b��4)IO��e�C\8�m�)
��B(od�(�D�F��V*�~ +��,M�@W���"|"�ê���� ��$N�$��=׉%���IsޣI�G"\��ɀm� �ڰ�ְ:f"���`�)U�*�QT$Oɹ0]� ;�f [l��l�o�����-��?���zt��]�vq�L;n��ʧYp[�5��{,��3�Of���J)���|��X �k ?n��1���~��=��mz'$��rI��0��0]� >ݳ �تm58�dNDܘ���Շ���H����m�Ԡ�N7�r`D��sO� >o� ?�X3^��}���dN0r1��`۶`��������`o]`G̥Nӕ�*�\�9�B�n�(�dU����q�>�8g+rɜK�3KqY�=�O��f }�fu�X���������U
-$$��}��ވ���}��~���k=3Tv���*�BP�G�z��vـ����^�ؓ��RN(8�q`~�Ļ���o�0��x׵`�oڱ�"�#��& ^�0��׷��=]���n�$�>AR�V! �T��*�#rǇk��v��Z�;q;�Y�׮#��7O�Fݳ^1����m��-Iˬ�pp�o����M��YW-�Q�n�d��<��=<��<V6j]'d�-͎s<sq�Aɨl:��ptM:`�kvYi"h펶����l�<+�m/E�g<�t��>�:�M^y��Ӵ��x�����m>n�.q� ��0�P�H-c���q���U�����\��9��(k�.�M�R  I�uÑ5i��8�"r)$�:���^���6��'��ܰ�U}T��%B�x׵`ݶ`� ��׀]v��"q����iŀvـ��31U��� �o� >�a�Qhjq�$Nq�& ^�0��x׵`ݶ`n�5�bnND�8䄒`����3�>��or��k �t��?D�\��)v瞬ts=&<u�� �m��uX�,6���Á���W]f��.�� >� /m���5m��7}d�0���9^$���@"�E����眰]�x��X�7mXۑC��'#��f�^��9Ľ]��*��^�U6��S�2'$��f&��}x;}X��� ��u�u&'��$Q���^Հj�׀���v�������6y=7t���Ԣ�v��s!����/s���&�]_�w�ݾo�)v)V������>� 6���ߢ#�;}X�㬡*�X�qʔ�bIown| ����z�v�����t��&f&���E�Y��(J���BI`^�^ ���&Dϕ|@��+ �����y�$�~���U]�nV��J-+�陉�i�`���� �]� �lM�q��2��Z�k�w�z&f&�{��>�}x��X�&#�N�����T�Ѕ'Nź�I	:J��L����;��1�O�ɂ�Gn�ڑ�"�#�NG����0����j�5wk�>펨�S�q)�RI�~����1�11v{��XS�^ ?�Y鉉�j���V��*�EAI^��V��^ ^�0�������)%wV�U������E�}��?y`���ܜ~DCJȉ(@D x����x�]��Ī1b��*RG�����_���z��j�׀Ϳ��=tXyM�K���Q���<�!Ë���t;:�4���������|��.9!$����]{V��^ ^�0�lw�Nq(�$$� ���Wv� ��`ݳ �lM�q�pYj�V ��� ͬ=鉉����X��Հ8�pU�5wiR!Z��� ͬ {�`o]`zbf�����qԮ��R����t�X �k �D��O��]�x �m`+�2�" �B"o�He�W+v����������&�"��vv��[\��W��A���c�ɦ���p��1l����R;:��R���x#N����<�9�+h��*�j���$v���}���Sok$.{ �TMAiy��ZųY�g��c	��ZJK`N��ͻ0��v��'2�i�i�(��� ���ɓ�#`�	j��v!^А�P�q���6�Yܥ�踆��Ѫ�,���a��Kf��#`�z9�6T]�x�@�eF�A������?�U��� -�`]U��4���ZUV� tۼ��L݇������u�X���\q��(��x{l�m�׵`[^�v�3��5���RI��0�j�*��s�{}�w�&���'8�S���0�j�*�^ ^�0ݳ �.���$gv����v����š�[�]m�l`��mr��NW��Dy8��0��ۆ{	 ���}x �m`zצ?Ps�ՀtS���m�H��< ��f�6m��ڰ
�ן�5o�8�S�q'8��I, �|������us����w^�F9N!�
90?������ ��׀�X]ϖ�}]eE��P��iȓ� ��xnـ���x��F�Q�@�bH+�(ծu�}Ӗу5�"9��fر7�d�����|��!�$ {�� -�0^ռ�[T���|f(�䋋�Ȝ� 7�����Wk�v��7�$�~�B�J]���}X��𭙈�&B!*��3{�����'��k �؛�up�q�MF�� ����k m`z"}�gz�Ew����|�>G8�� -�0�fkڰ
�� 7�/,MNF������T.�Z�7W5l����v�S�������9��NI��0^ՀUmxnـ}�S�1H��K�90^՝5GWw^ w>X �k n�;*-])�$�܉H�
�� -�0�fkڰ�\q��B8ǁ�ܚ��� ;�� ��d��7�}1%���1;�Ė�mđm� ��XV׀�����6��ث���)f-�;[={b�c� 	���v��:�hXn��u�W�o���X��`z�G�f>�7���9�S|o�p�q�C�� n�nـ[fkڰŷ�mX�#n�9 7�`��æ&"*���`o� w�cW�qN% �i�0�l�-{V n�nـv��I��A���� ��X��`�f }m�I� �xK�������褿�d��rÁ0�4�����"��Ȥ@7	��>W�Lv���T���h�>4l�,�@�cĐ�`����g��N��da��FI$*�d��	
��Ƶ��*�0��y0D�  �"Ń"E A �cbE�@���O��@`OZAz 9U�>��_{����φ�  � 
�V��iW��y^� :r%sM�V06B۶�� ;��_w�댛j�V�%�ć93�Zw8�=V���V�:4�f.L:0��eWub·-�m�a�R&$������Z�k����r�utvE�W��K��`l���@�!ś�W�w���!�*ݳ�g���xzZ3��N�ً��/&�먭�0 �/<v������Ӹ��%ӳ���:�َ�ILm�$�Wim5V*9�����ڥJv�0 5���5���^T�vee@��DeY���h�lwki��n��K��9�ԩ��*pu�2�j�a�k ��ԭ�G�[����=�kK\MB�R���	U)���jU�X��6z��'�'��۶H��l�q���J �!�)-k�==�<���� I[r��b�񩰁��7k��˹�7y�N�n�<��,���fv�%�y	�j0��u.pb�b�{9x���f�k�\tb�f%�S�簯mݻp�G#$��Ӧ�;a:�mƂ�Kgu����u @��[(�(g��u̻.�oRW-�n�����ە�\���SUPb�Uvy��r�6�m!D��91R����U�[\l誉2� :غ�T�ڀ��*�A�c�P��m����@�x�H�nZK:���9��g�*�I���Uʉ��㡄�:^���
2��Pu��U�;Z���ET	!J��8 [Bt$�[�6u�Y6�n������7E^��ܥ�,�j��nA�!�L����N��A�gk��as�`V�Ό�tMX�m �m�*��AZ��٪UId�˒�p�l	��D�{QLS̯#���nsfc�R#�۵a��Fqu�M_mm�kz����V-�	��&��z�ls�/Q\��m�ji���j��\�}�H3���Wm�(�BK���t���m=��ng9�"�#u���guvJ��%��W<������Sh3cC�� �M�a�GBD"�(���'�:8��������v�n|WJ��nݬmE��X�� ԭN.9Z�v^\�N͌��%���6Ӟ�E�+k�n�wf�lhz�&�{v/A;�6j�8��I�qFQ#��OO0�G��Ӷ�'����uKPas��m�\q ��˵ �s�`�h��'g2�U�]�2�[c�50qۭ�0�i�,<j�+P-=��e
�ʒL;j�� >�;�%q��N\32�����g��wi.�V;9 �S�]p f�dJ���$rcȘ�7D��%����_m��{l��� �����x��p��R9$�{l�� ��z��%�{n~ �Amww���XbKi$���X��Xz"b*��, �}0�bM�xD�$��rL׵`�X��������`yU�W("�\v��U�����|� }���-{V }���$��(�����猓�r�[q;:�`3�[K�Fc��j�r=�QD�#�ڎI����`�� 7v� �h���jq)�NI��k#�ʈ���蘉��ߏ+������v������	�i.(��-{V n�nـ[fk��1]ҲҊV�U��陉��m���� >����K�yo����K��"q���v� ��0^Հ�f�ߎ7����e�N�X"y"���F�n��4FLvG�2V��x�l�':%ur�V��͵�7z� 7u�LLL~�;�� ݱ&����D��NI�Z���Uo� w>X�������j
�Dv��U��� 7�`�f"!�Oܟ����Y�^�� �oڪ$6�ue+I`w�&.��������]`�ـ�m�&�q'�L �ڰO4�� 7ܰ�k ��J���.����x����ӻ;u�4�ـ^�=�	v).�{������D&�[�X�l�v� �`����%j)$��� �mg�b&*���`�ޘ׵`v�ĸ�K�� �K ͬ ����MW;}X �r�?n���2�݉U�T�X�����s�Հ��
����V?�X۪��w�'8��'�`^Հ+}���ޘ�l�-`m��%9P8>�]�"qH��n��j�Tskku��Y�F��Qx����N, ݶ`� ;m�׵`m��UD�db�ɀ��z�7����V n���wm�&�q'�L �`^Շ�~��$[�L ��� ���S	�@��� ��� ��0�ـ��뵴�Q��#�$���f�������L�ڰ��ze��.B7����N8��Ɓ�ᓋt�g��ˀدm�Nv,��Sp ���g��{d�""R�:뮪Os%]��mz]�:�w)\�WL��Km���a�s��E�l]\�w>���v:-grs.Q����Lm\me����=pg�����cs3�����?��|}sf��s]n�=A���`\�P��T�,S�tIu�
��6]��H� �@� �q@�*��]��C�
j�4��M�f�m���\vI��y�y���9���%�"\$ �9% ���{l�.�� .��q���� �D�X �mg�Q��V�Q1]O��a1BX�%������bX�'{une��4[3F��֪n%�bX����Kı/o��Mı,K��{[ND�,K���T�Kı>�۹���f�fje�]�"X�%�{}�bn%�bX��{��r%�bX���j��X��dO�߿]�"X�%��g����u�8��'d����h��{�ۄq�X�%�ک��%�b{��ӑ,KĽ���7ı,N�wye�ֲ���6qW�:�z���q���X���px�ͤcʭ�F�)*��~��ı,K�g�Sq,K��u�]�"X�%�{}�bn%�bX��{��r#D4CDwlqk�AZ�֓�Y��,K��}v��C�!�ꡤț�b__��&�X�%�{����Kı/}��Mı,K�׽�nM\��kZ��kV�ӑ,KĽ���7ı,K��m9ı,K�g�Sq,K��u�]�"X�%���E�kV�u���l#��DO����!ı,K���U7ı,Ow]��r%�bX����&�X�%���2�9K��!5�˭k[ND�,K���T�Kİ�c�����%�bX��ߵ���%�b_}�kiȖ%�b{������ؗv)rv���ѻX����n(۝O.���ycG��7&n�j=ۉbX�'����9ı,K��kq,Kľ���ӑ,KĿ{=���h��h�{�� v�-0ITr�#�,KĽ���7ı,K��m9ı,K��ک��%�b{��ӓ�oq���~g�L%������bX�%������bX�%���T�K~�B��[�۸���z���Kı/�ߵ���%�b_��I&�j�ݱ�n�CD5����U7ı,O�׿]�"X�%�{{�bn%�bX��{��r%�bX����YlF�KG���7���{��w�iȖ%�b_^�X��bX�%������bX�%�sک��%�b~�������r�:^CuwE��V�%�HX��:a�[/p������AГU����]�"X�%�}{�bn%�bX��{��r%�bX���j���L�bXG�w�q��7�CbZخ����kX��bX�%�������9"X�����n%�bX���~�ND�,K�����Kı9���d��˚�&�Yu�kiȖ%�b_w=���bX�'��}�ND��!�2%�}�X��bX�%���kiȖ%�bw�V�\񫙢Y�4fkZ���%�ȃ"w]���r%�bX����bn%�bX��{��r%�`~�XBJ��j$��D�dN~��j��X��h�}�����LX���!�K�����Kı/>����Kı/���Mı,K���ͧ"X�%��D����˶�kxkf�5sSSWZ�8[�$��IP�NKU��+�4@���������e�.��.�Z�'bX�%�}����ӑ,Kľ�{U7ı,O���6��bX�%�﵉��%�b^��33<r�mV�m�G���k#X�%��}�fӑ,Kľ���7ı,KϽ�m9ı,N�Yrz䒶�q�Œ�F"!�#��لq%�bX�׾�&�X�%�y����"X�%�}���n%�bX����rW�ڭ��,�8�h��h��v�2%�bX��{��r%�bX���j��X�%��}�fӑ,K��w٢�Zخ���Y-�b!�!�;�p�D�,K���T�Kı>ϻ��r%�bX����&�X�%�P��*�Q���P����ɭI���v�;���ӎѭ��qnT[����Y��y�;tݹ|�Ƶ���v��nU�yVɜ��0%�/V����sc�0`����;]���]Cֹnϑl۪�eJ���[';�;2���ܓ������i�
x��;#�(���;W4g��`���^�_�@�H���uu�u�&�.��p��Z���j儱��n�+"#��?V>��C���U8$��X�,�����F��5��x�u�qlk����s����T����ֵ��Kı/��~�Mı,K��m9ı,K��k�9"X�%���kiȖ%�bw�V�Y�JV���1��﷘G"X�%�{}�bn%�bX��ﵴ�Kı/}��M��ʙ����0v�-0Id��D4CD4C�����%�b^{��ӑ,KĽ�{U7ı,N��siȖ%�bzg�s=�Ye�՗%�f����%��@ș��~�ӑ,Kľ���Sq,K����6��bX�BdL���X��bX�%�h�I�q֭�[��D4CD4C�ک��%�a��}���,Kľ��kq,Kļ�}��"X�%�����5�����ˋ�*�^(�q̗!��V�΂���VDM�zt�����r�Q�%.�Z�H$�߻�&��	>��I�w߻��OD�,K�g�Sq,F�h�����;-��kv\#���q,K��kp�< >�&?#��Ȗ%�;�m9ı,K�sک��%�bw>�iȟ���,O��٦��6+���Ka�h��h�߷�m9ı,K�g�Sq,K��}�fӑ,KĽ���7ı,O����,N�NX��!�!��{U7ı,N���m9ı,K��kq,Kļ�}��"X�%��n��M�Bj�B��F"!�#Ӿ�m9ı,?1�_ߵ�Ȗ%�b_�{����bX�%�ک��%�b}��������������hs�׮5�q�HX�>ޣq��:����Wdax�������Kı/�����Kı/>����Kı/}��Mı,K����#���h���47&�cMZӉ�-��Kı/>����Kı/}��Mı,K���ͧ"X�%�{}�B1��}�I'��lv�lzֵ��Kı/���U7ı,O���6��c@�iw� QS�Ҹ�� FP���L ��X��o�t^�Mo�ƅ~Bbw���&���&c8,B[IxB`��М@$~	ϺJH@��j@������!��"!� $P�(A� qt��GN�"� *@�X�!�!i�����"����bA/�Mh
����bA ��J�E K+FF�,l�Ƥ
Ȥj
@�ejQ$�F6XX Xe�$��A��$Hqb�)I@���e%�H�#c�I&��@�zqU !�%x|*|)��\ցC�t�(�£�

�t ��r%��z��K�4C�}��!�!�;��5�%m�s$��ֱ7ĳ��@ȝ�}�6��bX�%���X��bX�%������bX�%�﵉��%�b{���-ɫ��l�7l�8�h��h�׻a�bX�ȱϻ����D�,K����7ı,O���6��bX�O{7�-�*�z@���Y�7N[mq�xH���z��xb�rH���07c���7KO��%�b^}�kiȖ%�b^��X��bX�'��}�ND�,K�}�bm�����r��a��n�p�D�,K�����Kı>ϻ��r%�bX���kq,Kļ���ӑ?��SX��bz~��ɟƮf�f�h��kq,K��{��m9ı,K������%�b^}�kiȖ%�b_?m�b!�!�;�� sP������m9ı,K������%�b^}�kiȖ%�b^��X��bX�"H�ީ�c�D�Z��m9İ���d�:�uԜN�l#�%������bX��+���br%�bX����m9ı,K��������oq����w�v$�DL�̝.A1v0���pꪙ@��v�����x�͡�[��;j�9m�8�h��h���D4�%����ͧ"X�%�~���7ı,K�w��r%�bX�z�����շ5r�e��bn%�bX�ϻ��r�F9"X����bn%�bX������"X�%�{{�bn%�bX����'q;,�9dv�#���h��}{�q,Kļ�}��"X�%�{{�bn%�bX���ٴ�Kı=���LK[�[r�%��D4CD4C�u��Kı/o}�Mı,K��}�ND�,��F�&�kq,K����L��L֩KsV�Z�ӑ,KĿ^�X��bX�'���6��bX�%�����Kı/;�kiȖ%�b
 �E`�#n���1�պ��L��8y�g`8�^7�:uڟknGI��6&��v�`n;u���c8vH���R���ڲWRj�,q�3�cV�m��v�{��ʆ�xj�tnI�l;����HV�8�i-ЯQ���v�Z7]�3&�u�r\r���kf�����!PGe�������\n6z�K�mqW*�S���t��8@�r�����c�C�� |3����Ed8�r�"X�	�6�ԝ����@�c�J�s�.�׊rN�ͅ+����e�������L#�,KĿ^�X��bX�%�}�m9ı,K�﵉��%�b}��s�����U+l�8�h��h���G� �DȖ%�߿kiȖ%�b~�g쩸�%�b}��iȖ%�bvxVM���U'���CD4CD>{w[ND�,K���T�K��"dN��6��bX�%�}�X��bX���	$�v�mV�m�G�'��쩸�%�b}��iȖ%�b_^�X��bX�L��{��m9�7�����]�,�2",�ﷸ����;�fӑ,Kľ���7ı,K����r%�bX��粦�X��������`\٩���&]Q�\>Y��އ]��v�h\�N.x����Du�Yá����ֵ�Z�m9ı,K��kq,Kļｭ�"X�%���{*n%�bX�g{��r%�bX���h�f�i�L՗4kZֱ7ı,K����rB�x���S�Cț��O�2%��}�eMı,K��~ͧ"X�%�}{�bn%�bX���L��˚�5sV�Z�ӑ,K��w=�7ı,O���m9ı,K��kq,Kļｭ�"X�%���L̙�5�D�ѭd��T�Kı>��ٴ�Kı/�}�Mı,K�����bX�'��쩸�%�b}��s���f�5��5�fӑ,Kľ���7ı,?s�~����,K�����Sq,K��;�fӑ,K��Ο��A�� ����n���Ԣ��s�l�b:!{&˙{�����V��ݫS��d�,K��ߵ��Kı=��eMı,K��}�ND�,K�����!�!�}�$�C��m����Kı=��eMı,K��}�ND�,K�����Kı/;�ki���'���{�3�w�y`0",��X�%����fӑ,Kľ���7�����⡡^D�K���bX�'��~ʛ�bX�'��͉�\U�Uv���!�!���X��bX�%�}�m9ı,Ogs�Sq,K��;�fӑ,K��o�ˇ���������oq��;�kiȖ%�b{;�ʛ�bX�'���6��bX�%�﵉��%�bs�,͹�@At����pD)FL�d�FC;�=�0�ep;T�kd��Fݺ3V浭�"X�%���{*n%�bX���ٴ�Kı/�}�Mı,K|�ۄq��^�H��c�UF���YSq,K��w�ͧ"X�%�}{�bn%�bX������Kİ��H�CD4CD{��@���U�Z�m9ı,K��kq,Kļ����"X�%��ﮓq,K����aD4CD4G��d�c�J��;�ֱ7ı,K�{��r%�bX>���7ı,N�{��r%�``�� #����D�'߮�kq,K���G$�:���[p�"!�X>���7ı,?������ٴ�Kı/����Mı,K������oq��������|i�+j�y�g�����m��KVQQ'�'A� ���L� �xjn*-R�t�"!�#f���%�bX�׾�&�X�%�y�{[ND�,K��]&�X�%��k��&�J�Uv���!�!��m�b%�bX������Kİ}���n%�bX���ٴ�Kı;��јf�آ��[m�b!�!�7v�D�,K��]&�X�!�2'����ND�,K����Mı,K����gQ�P�V��!�!�v{]#X�%���}�ND�,K�����K��$ș��ߵ��Kı==��)�JT[k��1����ͧ"X�%��s���br%�bX��߿kiȖ%�`�;��Kı;�����߆~��-ѲE�V�B�y����������c:ݺv������X8�%J�'YqR��%z%��٬j�wK��-h_a�Q�w��Ok7X�p�ɘy�J��mcleڻ8��<vw�F�#p��cj�Y[G+��ʚj��(W$�z�c%;g˳��;ۈ:���Cݧۤ�ZMͮ��tg�
{SW�9��q��ɗ5�ˬ�	�f�j�!�?
A �  s�J�E�����AG���;Jv��L<v~7l�u��A�;Z�L��q���(��NKY�ZԶp�D4CD4C���&�X�%�y��[ND�,K��]�Q���,K��~ͧ"X�%����+���ݫS��{��7������[ND�,K��]&�X�%����ͧ"X�%�}{�bn%�bX���I��l��dvۄq��;=��Kı>ϻ��r%��D"_�ߵ���%�b_������bX���]asRܚ5��e�]&�X�%��}�fӑ,Kľ���7ı,KϽ�m9ı,g}t��bX���׻������f�CD4�%�﵉��%�a��}�ߵ��%�bX?�߮�q,K��>�iȖ%��{߿�]��6e)�Oƥz��L��m��*���Zײ>x{T�]V�惫5�4kZֱ7ı,KϽ�m9ı,g}t��bX�'��}�ND�,K�����Kı>��&rjkY�]j�kZ�r%�bX���f&�NlM�V�YJ&�]Z؛�b\ｭ�"X�%�}{�bn%�bX���n�CD4C@��9�\�&��+5���bX�%�}�m9ı,K��kq,KĽ�}��"X�%����CD4CDw�� �[��l�e�ӑ,Kľ���7ı,K����r%�bX���f&�X�%��}�L#���h���Ь�l��PV�e�q,Kļ���ӑ,K��^�17ı,O���6��bX�%���CD4CD~�o��ح��-���s�*�<�'Q�C�ƻ74�]e�W���!��N���鬊��3LJU~����7���{����17ı,O���6��bX�%�﵉��%�b^}�kiȖ%�`�xk�9[qQ*�7,�b!�!�;;�fӑ,Kľ���7ı,KϽ�m9ı,Oe�q,K����К�֘�V��0�"!�!�﵉��%�b^}�kiȖ<L� ��|�D?��N����ى��%�b}����iȖ%�bw=}�0�[�Z��e��D4CD4C�wnȖ%�b{/}���bX�'��}�ND�,�dL�}�X��bX�'�~?H���L�ն�D4CD4F��7ı,O���6��bX�%�﵉��%�b^}�kiȖ%�b{��ߋ=\ȓ�ة�۫�0gI�մ�6��v��� k����.~�K���L�r%�bX��{�m9ı,K��kq,Kļｭ�"X�%���B1����I�KeA�kRٴ�Kı/�}�M��Q�L�b_������bX�'��~ʛ�bX���l�8�h��h�-
�&�\u.�Z�&�X�%�y����"X�%���{*n%���Dȝ���m9ı,K����7ı,Kߺffg��W,����!��	@DG�gѦ�X�%���fӑ,Kľ���7İ(��	�h77^������bX��٬.jۓFjfe��T�Kı>ϻ��r%�bX����7ı,KϽ�m9ı,OOM��D4CD4GW�=�� �&�M]�����v-���x F*��yݕ�^2k��(MWkLZ+v��G����&�X�%�y����"X�%���{(_�j%�b{=��6��bX�{����]u�9ji�}����d����ӑ,K��w=�7ı,O���6��bX�'�}�Mı,K�ѩ78��Sv�m�G��{���Kı>ϻ��r%�bX����7ı,KϽ�m9ı,z��������e��D4C_�������m9ı,O���x��bX�%������bX�"~�����K�h�{�r	>q��Z��#���h�Ӿ�&�X�%�7�{�ؒ	"zw�5�N^}�ؒ	"�Q_��Q_�ATW�TATV�
���*���U���
���'���"("(� ���B"�1� ���
�1B"�0A���� `� X� �"�1"(��Tb(� �H� �H"�@�Q_��Q_�"
���QZ(*��DE�*��� �+�TATW�Ȃ����
��� @�E�ATW���e5���v L�� �s2}p���� (PP�*B���@U*B�   Q@\�P
  TI PR�B$
��� *� %@   �@UJ�(�*�R���p  ` P J
�7,GO�=qn��\�/K��>������}_y�*���J��uz�W-J�`��R�bj^��  ���R�x�����P���M*�Z�*�Ԫ�&��` 3URϳ�R���z�a��-�J  p � EPv ;�B��   � P  e����e���X�UQ���U� �룐ub�;�@4p;���,|{*�� r:��yy��n;� w�w`u�j�Yʙe� �    >���;��{�Nm��r��8�Uch^���=f�k�L�ch�p �XϧS�μ��rX���ӽ#���`��s��c�ũV7���ťL�K���� 
 �Q (vt >����)��1�MJ����$���O�����#��ޔ��;)�n�׾��2h_p'�������m_m\�\۞�� GS-U3�}yx���{t����    UJ(R�n��}ٗ'�G3;��6+��ȳ���JdҬ�|��d�Ͼux }9��خL� Mq�F,+��
}<��}����%��85���ސ�u�����vr諀z�$ޒ��� ��� Њ~=T�Ti��	��&B'�T�i��d ���(��IJ� 
BM�)"!����S�O����������o���Y5	K���GX�{=���Ez���Ev*���������E�DU�TPT�?���� ���I��'��t�4��L�A�����%�?��ۆ����ټ�M$h�Ӵ#�N�sV�-Ca��f��i]������Q�FД�1����?�9(����bt�H�K�4�D��Q���������z�J~�����sXi��kEa���TG9k���;X�H�@�b��!	�[F5{
!6Fhٺl�r�j�Z0Y�����Q��B�8 �H�b��	��Ǉ�����һ�y�f@EfF:yc!)f�P0��.F�<�0���������h�q��Z�to7��(�L]�,0������/sL�]x�0��4�0�������Q`�%�5������(���s�61�`ap��:�F���ka�~qCB����a�����0��N)&:����$֍o���t#La���a��AFi�W�a#"�0'd6����h#5�iE� �@�d�q� c� �A�BT�fw����cd~�-$����cL�LLc�����b!�X!�H�`�	p4��0c�n �5�уB`la*�h=H1tW�.2��J�r�? ��N��ؓ��4���rq#:o���e���Y�X�ִ�@�\�8�8����a�)�T�_w�B�PA��y_��8Xi�dd�\��X��}0JC���@�Bc�.@;8��N��`Z�3�bXi��xqߏ��~6`0c&0,mo�kџ]$&:CHFa����	H"k�2}ۆ��zx0b�v�ņ���I����I����0��a@�q��,�Hb���J,��"0xl�Ɂ�%` �P�����8p66x|?=`�Iz���3v]L@�k�A�x��s���q�p ��X�L�)�-���	 BD�k ��y��9��M�$���4/��S򮗨�4@ˁ�g5ae����$0tmc@`N����6$�	�N���A��4n��A��i�L4m���<s��k��CS�:N&���6 A��!�[	&�%V�B��	/�J,�`�i�4b��}c4�aNP�6��>Np)p&-@ 9ȹ`K����)��q�$�9�XSY͗5�5�O�<c��p"��h CFɛ���6q��$DYVL���#4Z�;��Grc@�ѣ�sT�΅�|) C��1����3��N��٬78L��D%�����~4�2k���4f�32B��,��b�E��0ɀ�T6#�iؒD����%$C4#�aId1B�Ю�0W@�Q�J��! �+�� !1	H%�BB�!���с��@�:D�� �jqI2k5�,��j�Ũ	4���4l8�0㥳3Z�m��c���!��������Q�!F�`x�O��h�st�x�a��~Y�a���20t��s��x��#��i���tNj�<�������� � N6*�ᄦ �0�E�mJ�#"'s[ẌH�"H�@Yk4m�) �\MG1� �+[8���h0�*����@Z�[��Ï�I��s2*��a9	�Qek�<�;����t�f,%��;$�yEFh�o�V�Yc5��(�6�6Zٴ�l�B2�0Nq�L�$�c�p������i�qᎫMAoY���D��xkÆ�\����$H��]	��Q�q�`�/(�Q)D�\|(1
c�,yFbGPM(!��6:	X8�İ0X@��^�CbL'v����bjq�t H��bFDB[�s'2��8Ʉ�����a��L�AD4�=Yq HIǆ2C @`���ၬv��^�.oG8D)�� S��r��1�A�F�"z4�n��i���)����HSF,�����F�x�N�����O��cS������6&�B42S%�1�	�M��G��Áz�@@B<3���@@"�0^b\�T���`0b�D��h�x��Ս� BTj�4a&`l���-lᏓ�h�Ç�FFFXi�p��y:v���XhZ��-�#'���L�;x,�g2�������l�c)#�r����\B@�|��'$�99�BH[�Cb�'��OڼX�01�D,�FF�u�	�\5�������1�'X2��)!:GC�\0��(	�&Lp�&�K�?[]�����;]P`i����;xIY��N��{���!�$10t ��4XTCP�l�E^NZ3$hf6e�ؤ�̴#��)�~���:t�Y�c��;Ʌ��ǧ��~"$�(�H&BM�x@b�h�	�$ %#`&�`��%c�n����G),޼���t�	��ff#8���a4�L�F4}�8�m�s�&\����NCĎ)+e����&I@�tnyk�s'Ld[����F�0i�1-c8�`N5��$��3M����#2�xp�0�����Ӱg0ְ�,V����f��4�`sD���e�9�d����Ww��q�N�p&�|3[T�8$,��6pʰ�Jc��u��!6T	�偓���iݫF#��1�Y��4`�0��:\]5�+�'5���&���֭,�n�N����H���`�0��c��������S`���>e��Gs��PN�0qrpAт�j��;T]||��L��w2o�!�rK|�����x�LEn!��r��X�N�U���P��:*cS\���&�wQ\t��eN��9{Z�	��I��	:��B����#�
&����x���3(Y�?/s�.��=������(r�
�y)J,"go�<�p>g�⸖H^'PS��*-�	�Ri�R�v�P��� $�`P0��Զg8!l'U�rP� PA�3#d�1��'h�	iŃ�&:�	hPd��8ř���}m�Ù�[Xڋ���
eS�x�\�RR��@9�2S�1���]��L���=Œ�@�^|3��09��g8�+�7s�F)�}� 	MX�(���
@I�'(� PP�EN@�"�s�04_2��*A3Dmw�)���^^�m�R�b����D'x�QR����O� �xy(�$#��r��}�b��p � r�#�;��ވ�^!�\�+�Qt(x$���л��L��\9w�>gp'Ĝ�0<�s.,����
p48x���C���у��c�ù�w7�<��
���28,�+�
����W.p�>9�fvN��5�ە՜�9���
;����	��VpL|If+�8��/��&� �����"9��x��O��n'Ą�Y��	$� ��1Xxl5An��AibgTU��O�Ɇ��d�8a8@@�K��	Ł�PEŀ�x��\]o��5��6����������Æ��A��������RN3����o���ѳi(21`�CN�U�$@H&Ѓs��#F�̵o���IW4l�[|��F�;g1�I��M�l���|��o��0�%���M�Z�E<= �'@It$[�h<ӆ��)��$c�$��~��Jl8l<a���C=?�ɡ�n	������4�[�c�a�v��c8E�pޱ�98�xq4�Xa!�N��(�� �pg���qX0&1Ib�І�p�l&�e�a(��HKݝ��m��h�m� m�@ 6� �	  $�   8  �  ���9zi:���y\�w-�P 	�u����    [G ڤ�"�q�6��$ �M��� ��F���o�km|?J�J�m���	 [@ �l)A�g���	���`�-2�Uya1�^{*���s�mm+�w�f���E�q��o'I�MVG����tِ������Ã�D>����ǷH)�\�ږ:�t�#���:�^�����+��kW-O��wQ�Ō=n$�$�wez���IҬ�ii�g4I2Z�n��,����]��W�c;�x�1�i��j�n��.����pDO;Iڭ��u�m U�ki���<A�Z����9���\�1�F*r+O[N��]L�9¼8�|�M��*�
@eTV��Pݎ,�y1����q�]�'Q�CiKqu�	˦�.���ic3y'������y�n=��k�f����4������m����ݵ��$q�s��=.nҬ27:4�1\�9�m3�#U�=kC��īdrZ�fZ�1%���r��rd	�y�S�m�ø��̾I@��7,Xtvce���O=�����Bi� E�i6G�,��(�mgl�3ӶB:9M����63B5U� hS[��  ���k�8 l��Ė�Jp��     �h�6ؑ!�� ]6�l�-�e��6�	H n� @  -���!�m&�~�l  ���ݴ��HH  R��  m�E�[@  ڶJsm�`�   n�i3�  �B� H6�6�N�:ĉ$��d�-�� �[���km��ݷg H��� ��iz�U2��p�]�\���\��u��[L���UU[J��6]����8��7m5@6��(Ӌ��Y�[��QͶ��L������X��K���lF�6�m��N�UT��A(RT�pU)�6���[T��I�ש��m&��.�/�h�<�d�::��U����{�K)��כ]��� 8�kz�qm�jD���vn)�b�]�k]=�-�g�P.V�l6�-�酴v�	6�W��Xf�v�L-��$�`�U�pv�L�aͶ���`-��8��n� ݶ[% �� }m � �$ �lj�	87ְ��]� �[%�mHkX  6�e� l8 [R7m�/P��mj��K�g@�J�-����@pm�Xn$6�^Ԛ5�!����/4�5RN˲�   9 [@*U��X.�٨
�� ���2ʰ�h�[p ��� m��-� :�m���M�I&�l  ,W&�հ���m� �` R���,��[�}|�4�̄�� �m�-����&ݳ���W@��nyƺU�T�V�!-ձ�N;H����Hx��K��jZ��-��Uu �*��U�eь"�j�	U���4�Ap�f��S���U��4v6��^�8'b(��j�,����ls���U`6࠴nT[@ �m������o�m�z�����F�9���d�m��8
T�� [@i�6��lE���e�$� 9�:��U�vl!�Hp+UUU�[!	�+@PlT�2�ɐ
��V���T2ښ��m��gg�٥ZN���s���m���	l���t�H����M!�}`$�d�Z��8+�Q�(SY�]PmMt���n���0d�	e ͭ��m�ҷj In�p��ٵ�N�[|�-�kխ���l[E� �` Hk���l #��������!l�����q���m��շU=j�J��-J�mm��j�B�ڪVP jv24�,�-]z#�b�$ր�`�[/kn79eg5Y.�w 0����gm�y]l��"-m�c&%�.���m�m����ڪ�U�[!���� 8�i�����Иn8�S�j-�M���  r�m����P�������[�ր�����S�1�Jv�`[�	f�� ��fDС�A� � 8� g� 6��[B�v�`I&�!��m%�m��LU�A����4]��� �mug�����i$#vt3Z��^��v�[@-N���r�l�- �e�� ְ H  ���` �� �� �A� 2 � ��5��8 �  j�[e�߯UR�*0"ԁ���ے� [A m��T�@[���6Үӫ�m���p@ֱ�i�#]� 8m�` m  $[@p 6�@ � ��ٶp�  [��	ԁ�������[B@� 6� �tV�X6��-���m�p�!v�knؐ8[%{oe��H6 � -�m۲ ؜ l�M� l-�j�Nڶ�H�               l @@$6ٵV�)��n�C�6`+ҭ� P�'�M*�]UJE�;i�  �5T��`��-��Rj�69r�� M� �Yd�8 r�n$n�]���m��-��  �� 8 �@H ���  m   ��mݶ		  ���X[dz�Il���p�[���kWV@	 -� ��)m6��v�[y���4ڀ   s���n�L�!����  �� [@;6�i�m   	l�[@  �p 8�l ��ċh -�l��ې  �m٬CT�i0  l$��  �`�   H �� �`  �          H��6��4���8�  ���)lHŵ:�
l5�VhH����U��4͝ϭ�,�E�۷ ��HͶl��Ue�j�U77\˰u�ݻ5���2ԀH�Y@ ��8e�l�    	6�&� m�e��I� [I 	��i�l 4ڀ�  �̹E�BB@  l    nϞ���� .�r��R�uR��,V�@����6��Y��l ��lݰ�� [�� z��iF� 6���t�i-+
�-��uJ�UT�۵L@  $ $I�����U��$m�M��H ��cm��"Am   -�  �f� �    � ��  ?�=�� p ��    i   	 �������        �  `�  �  8�5d�ST�#�Z��Z�GUU�R����X�ڝ R��iG�gH4�:�ͻ` [@8 �  6��p m�e� -�Edt��	�{5 �T�C[p�� 8)�]UD�l�B�I�ְm��kj� ��R�l��JK[us�nY�e� E�@,3�mcV�jP 	��*�lQe݀�iVU��Ā m��� ��t��z�s��u]@Um�ԉZ%�f$��	���m	      ���   � �  [@ lH�m�[W�M�A�v��m� �/���[$뮶��jB��H�֝�*T �ya�<�V��  k��  ��l��   /v��b���ٶ �\Jku��,��m�����mR��b�-4���۶�m8��R�J����=��$4n� @[A߉g�}U֓��6U�eZ�@�.�� h       �`       �     hM��ٶicHm�n�������4�kXR��n�2ӱ!uZ�V��h���jM����K���L��QQ89bZ��E2����d� -�cm��$}v�����f m��S���t[@֙z��pA�޴gBl�$vU�[�˰�E_��tJ�.
Bu	h*�m� 8	!j��8�`��Z�)j����kem��o�[�~([t�l:������e�@J��@*�<�ʥ�V�Q]��*���C���*+e�`X�Jն1[7 ��m�&�/Jֱz!�]U*����cM�D�m&m����	ѕ��
eej� mq��Tpv��8 %ZVVݍMP�m�6����z�Yp�H��l�o ���7�V���� �\��:���hy��j����zRU��U��ʫD�`(� $   H�^+Z�m�v�R`  -��  �m��a�Ͷ  �M��[�� ��$��  []�m�Z�6б[-Oh�l�v�EG��ث���N����ny4���$��[�{p��9��EU뎥�n$%7nm!���rT�.�UUJ�o{7��Z����
�U��@h� G�>���"��\]hU�G�:z�b pE qFTFR>��Q?~�`4��'��0�h��� �!��Y]����}D�)�����#��y'QS�U8	��=S�"������Ba)QF�a U����EpQ�=�P꿝$�� t��@���TOP x���@Л�SH�
q<$^!��.�#��T��=G��A�ߑ@��6�#��7�����C��v�"!�M.�<�`��|v������_Q}�Y��Q��!ꎄ䜪��ʊ(j&�&X��[,�h
J"J� �a��#,��%��êy�����D�"�0��v�  翉EE��UL�j�DEQ]�����	@) 9��B,���@D ]�u�#�%,��m���n��h�GVh�&6�`���=��eLU��i�L����H�9�N����Ѵ�ʏ����Y�'؁��R��m�s��[��2g�=f���9�-\�����bΗ*�Ó�;i�-�W�y3��N��i���Vm:[m�"��4��km���x�4HsT��U*�t���*��s@6WV��o����;Nh�ձ�#Oc �n��vv�(iQ��m�vػ[�a�����ץ�]U��e���tc<@v�QȤ�X�YU�U�QA��y��{(�gS W
�h�XI�0I���ۉ�[�)M�<�wg6��"�f��\��Ў�����;dǖ�7c`�˫i7V��M��l��K�t�i9�^�#f�:��ړ#=�9��l��(�aS�:ڴ��iЭw=�7M�X,��M�d�t��D7GV��l����a;b��U����!�Qd��;P�y���j��:��"kY����%�T
VW��ѓ�8��j�ֺ�)\����db�P n]��B�:���E�t���(K�sl���  �v�-�Eh�퀡�K��p����)���l0I!�&ݳ��؇O85�Ԛh��(Ԅ��+�·[PWl�cB��$�lm�[@�sК�6�c+��<!n�ښ�����8�Rgi.��څj�ʻ�r
+<%e���ە�I'NR&yt��1KM� ��M��`��EP��
�
���9j�jU�`�b@"Xΐ�4�i�VM�ʜ(
\���`J�]���-��$Ci*���s�N�̮���w6gj��yBc]�y���]�;><�l�� ��9#wZ����i쾀y�G9��ZDnL�tjk����6��S=�Y�V52i:�0fN��#�(h\�\C��z93���g��b+;��<<�ugc�a��I�F�@�ڶ��V�ݳ�I�.��%�1���EcHA �A @��*B�3�2�)���A���Q�QxuҌ"mX  FpP�ҝ	7M��b	2㢫v�c�����{fŞ���5 �]Ж�[A���Z{Y��K���fg˻Y��6g�FJӚ��&�\�=u��s���&�6/�T�gN(+L�e��TO
�-5Gj�]rg0����k�I�dR����+�Ç@�Pt��.;�������<!��'4<6m�9���ن�(gY]uKtm[���EN�!x��o�� >��v��r����=�v\�T]�vQ�v�)��W��C�Y]���� ;�������3<A~w�}�\�(�#r�E��]���\�P��#���>�*��w�U�^��{�g����5��9#����_l��Wuz]��/j���L��nM�e4
���*�lĀ$����\�~��	efZ���*�^�U����@��4����:��#�q��9�:ۜ.θ]�[��͸j��[�\�%�o7e�����w4zS@��z�R�t;S�ڲ�Io�pg	 �$x �D8�"�w|�.U����@-�4�d�F@��q�nI��ڴ
�נ�����Τ�I��A��H��@��{����}o�@����}v���FIR���W��k &be���۬�[�6�����%7I˖�䫱���5�����pb��c�y�����o��"\IIK��V ��� u�� [��ڬ��L��nM�hu�@/u�z٧��=k��A㖨,HUj�]n���aQL��!#H)2�£�0��D ���GK�4�Hd�����g��K{��)uT��Ǡ�f�z����
�נ�,L�bqa"$�@�n�y�Z]���٠fg��g��7,9�m�#L�֞�s[];�,M*Ds�9���nb�v���]���Z]k�������i*�c�t�����Ҭ�[�ؘ��{� ��ۚ�j�.^�Td����(ۏ@/[4��h��@��z��}��WJ*)B�+K�k���i�s��\�!�&�(����>��g�q%׿=�:㖩���j�*�^�^�h���*j1�]��v-������S���[s�v��F�]�c�v��jΎn�ͬ"������k }o#f&&yA��k ���ѹ�B#�0n= �l�/[��^v����ă��&`��D$G&�z����Z]k����c�c'�m"!�&�yڴ
����� ��4�%RF<�ŎL��@��� ��4��j�PxyA��2���*��ٍ��tM�q��\}�?���<��!�9�;����(qk��U��h����<hӇJ�E�k#��ҴR���8�6nݷb�;iH�Ð:+j�v�5��$�B����8����l,�{9�2j�ᓲ�v���
[2��O�Д�s.���5�fm����1��a�],���wn��׷;3�����GsH4�n�%F@ꃀʞF$ƫ�S�lnKb��Y�����9zg��j�����s�ܽD���"���������}�h�S@�ޯ@��_ǒM�Y1̘����MX�y�Z^���l�=]k��Cr
dp�rh�U�U�@/�� ��h��� �Х�Y��Ik��ĉ	�ݠ�$R�}��┥'}�{��JS�{w����M:��K0��! w��D��w����);�w�<��;����31艞�/T��P�E$�!"�3��R�@݃�M��nb�fΙ�))x �H�����k-�{%)K����)I�s���)����({�{��=�Msc�WE�Բ�$$HH���pyt�bT�ܦg})C�{ݏ%)K���┥'v�r����Z,�����#^�f)C�{ݏ%)K���┥'}��!"F�V�(�[c��0��?,���%)N��}�)JRw��q$y���BD����?��X���3{�e�oc�)����)J?����`�)Jw=��qJR����JS��7��'$H��p7g����ظ/nM��hc�{U�����YY� R�ӣ7�޸�)I�s���)�~�u�)J���y)J~���qJR��{�R�0�RĬ��X8�	<�� � 	�J���JR�����)JR7�u����#�yn�K���ݳ�({�{��)�w��S	�� ��+� ����s�8�	<��HH��^ձ�[tWc�ƭ�D��{�HH�����JS���u�)J���y)Jw󮹱�S���u�f$$F��qR���\R����ǒ�����\}�{ݷ{���ɋ(u���m]Y�h��ȲRɷ$� n�g����s�Z�9�\"���Z����#��ل��	���JR�g{�qJR����H�u��Em��U�9%�		}��y)Jy��u�)JN���JS1��]������j��v�%E%z���JS�}��┥'o{�%)#�۳		}�A�HH����Cu�� u�0��?�$��߾��)���k�R�=����R��� J�\Iy��\R���~�J��j��7m��$$H����B����ǒ����{�)JRv���8�	=��A��jZ��B��x+�7X�8z˄��u�nն뙒u���o1jAUlrY���	�ݠ�$$H��{�)JRv����R��;��R���[U�ln�j�A�HH����'׿}��)����)J��v<��;�^泹�v�l�#��0��!"5wv���#�wf�}��JR��{�qJR�Ν�T�'C����`8�	<�va!%({���R��;��R�����!"F�w\�ʭ��$�K0��J��v<��>g����)JO�~�C�JS��{�)JRx����[>w��6F����K�۞?�~�|�q��^��:�հf�3Õ�۵�>��Y���eҨLE��A[��68r'&�z�F�n�P���QL�=]�"o3f�t���� ��j7l�;n���5��*����������*�S��	��'m�A��c���n�l�n�m�!�z�HӴ`�ɗc�����\�]��u�T�V�����}�w�K�����˫`z�r:rͱ�S��A�=�#a�%D>��qQˑ:��hV���Ȑ�#�{��qJR������)�w���(������#ϻ���+T@�qJR������)�w���(w۴D��{�0��! {�lm��j��;-`�$$H��ل��	���y!���N��}�)JR}���"BD�w��҅�U��f$$=����R��;��R���;�J����$$HH��qkn)b浬޷��)�w���(� '�����R��}��┥}�v<������~o����p��S���f�{r�x�-�;i��v{c�%�[��x���-��7`M��{┥'}��������\R����ǒ���{��JR��N�ݩ"tU$
Kd�����#�wf :H�,���J���R�����HH�����HH�����"�ج��#��$$HH��!"B���)JRv����R��;��R��x�E(��	��*҉�33���)JN���JR��{�qJR�}�A�HH����Cu�� ��p�)I���C�J�=�ǻ��k�R�?w�<��/{��R��������u˺���[��v�8��a1v� fۭeᗋ��,�]��N8.�ԙ��C�JS��{�)JP���c�JR�����)I���C�JS�u�{��n�Dk[ݭoz┥}�v<��.���R����t<��;���┐�=�����Q��;-!"B�w�┥'o{�$$>m�Ze�܈��x���?])�3I:8�@���9���]��d�4��H��$��`����rq�%��!0�t���L��5~�D���2U9��p�����j�`wtKYW�bC4�U$��E� 0U�	�������.'(| '�TօG��O�%=����x2�~��I�Ò�u�sY�kn�l�h�o{┾
I���hy)Jw>��q>Qa�J���%���;��o�R�����3Z�ۙ�Xk:���%)N�~�\R������c�){��o�R���w�<D��� ?ߓ�1l�ECr�]=-0�c����d�iۣm�ZV�I-u�:�~s�ת�V�V�T��W���O��(�&`%.���R���w�<��;����$$G���_�:��cv���"BE/����ⓒ��}�}��JS���L$$HH��"BD�vn��;,�WUN[���	��X8�	5���)J����R����|R���{�Z�0����KX8�	5���JR���v<��.����$<�d쇈��G��yo��<��<���UJ����%�BD�����qP���Q����/����|?Y�K���0�J$պ1=vŭ�M�틷�9�*�!��l��5��фgr
�]��JR����)I���C�JS���┥}�v<��;�sY���V�&�R�p��!"7�u����#}��IJP��{��)w��|R����U7#u ��䵃���#}��HR�=���y)J]�{�)JRw��8�	;�x]tW,N�]�Kp��%{��y)J]�{�)JRw��a�)���┥'���o�Y�Zճ[�f�V�������~�|R���{���JS���┥{��y)J~S��̥�'�l�m��0'u�VZm�yw^�s��!'[�UrgC��h��:��8���ͷ.�r�br�N���"����E=�N�j���m�v�ۚ�;\vۜ7dq�v�fɪi�Wkm����g���n�p���ȴ��iÒ�l��<�����L���Q�<�� �Cם����GZ�mY�&'F���о[�%0��D]a�Flu{�[�s�<�AY�l��]�|��kvh�7���]���n�,�EeUIo		#ﾟ q�;���┥{��y)J]���		#��ړ���5lvZ��H�;���┥}�v<��.���R���;�JR���twy���Z��ַ�R����ǒ���{��JR���]����}�{�R�����dZӎX��9,�D��wv�!"JN��vJR����┥}�v<D����u�]�	Br!%�		����<��;��u�)J���y$$H[��		#�~kkjH�;[��ۆ���sیu����&��6�5Z�;k�/��u$�QSr&�MT��[P8�	5�vqJR����JR�}�w��%�H�׷�N01݇B�P�Ք�RIU�8�)C�{ݏ#��QQd5)}�~��)<���JR���{�RD�����؝J��BR�!"�����JR���]����5)�����(~�߶<��?{��6f���[VUS��!"BDo�j!"F�{ÊR�=����R�����(��?jN��4ձ�k!"F�)JP���c�JR�{��JR�|�X8�	> ���_��쮫E�z5ֆ�n�x���u�l>�k���m�6�P�W^�L��U�4�t�h�!"B@��}A�R���{�)JRw��py)Jw���$$G� �ѱ��M�Z	����)J_}߷�)JN���%)N���┥}�v<��?v5�k;��iJr(�HH�����HH���ۊR��  ��g��n��$$H]��!"BDwۢ�$n�ұ�S��q$n���BD���n��R���{�)JRw��py)Jyм.�+�'R��$�		}�A�J�@�����)JR}���J$H��Մ��	�{j�H���D�m�3�5�E%�6΄�M��g�2+3�cW@4��1:$���V���"BD�����);�w�<��;�wۊR�=��!"G{7]�%
+k��m�JR���{��JS�׽�)JP���c�JR�}���)I��=�f�,�K�Im�D����0��! w۴<��.���R���;�JR��l��*֘�Jk�a!"B@�h8�R�}��┥'}�����$	wٳ		ڶ8��t%+rYh8�	��p��!"7�u����s�{�)JP���c�JS���_��Չs�<�0mZӴW1Xg���KZW�5��L�Q,)�Lݹ���.s[��);�w�<��;���qJR����JR�}��┥'�}�5�á�Kv9k!"F���$$HH=����R�����);�u�y(�#���Er����[�a!"B@��ǒ�����|R������R���HH���{��N�%*ա-o{%)K�{���)I�s���)���u�(O�l����ǒ��{���RKSYTNۄ��	�{�D��s����({�{��)w���$$G�uSڔ�5!�2*�t�=kn�v��ygه��ݢ�2N�9�L�LA�״��Y�@����X�7����GO�x������Z�z���k�֐���ǇG�q�+�nQ��m��:In!�(VHN73v.�"�2Y{n�qB��]�nj�qW��t1DW9���� �m,�vdٝ�$]la�:7Z+0^����\������[-<f��+pI�&����mT�қ^�Cs`�]�[
%ꕪ;߭����~��({�{��)w����\������<��>�Y߳{m�̵ ��%�HH��;��"BD����)JRw��py)Jw?{�qJR���vH�IȨI������!o}�	)JN���%)N�^�8�)C�{�D���<�ڢV	ER(�HIr���{��JS�׽�)JP���!"B���$$HH��tT�:��r�"BD���xHH��;��<��.���R�����<��.����/���n+K�lnKi��7i��Ռ�&���0;!���n�Mb^��jt�5���({�{��)w��|R����a�)�����)?^���m�*VP졩m���!}��p� J@��~:��zq�R�]�^C�JS�����({�{��)���ܡ�$�0�V4�HH��횁�IJw����)J���y)J]��$$G|���IH)v�\�D���u�s�R�=����R���{�)B(�'��_C�JSﵝ�7���35"��mxHH��;��"BD���R����a�)�����)?~�᝗���+�z�^0�y:t�N�vV_m��#�Ƙ�������Fȗl�[�ǒ�'�Y���|R����k�y)Jw����)J���y)Jy�]�6�\��#�9n$$F�f�q�	���w�┥���%)K���$$HH������DM����;�{�┥}�v<��Q�Ց͜����o�R��w�}%)G:��p[m��e��^$$�v��������JR���]���L�00����*�ijH���>JR��w��JR���]����v{^$$�v����#�[vF�	OWa�#<��:ї
v,����i�F%��IΝ`p�qҕ�&*���)I�{���JS�׽�)JP���c�JR�}���)I���]��Z����������JS��{���������R�����)JN��vI�D���~v�-��"��exHH��?w�<��.�����?�R}���y)Jk��┥���sV�7�5��o{��R�>��o�R��w�}%)N�]�qJ$$I@`�˭z= ����s��JR�w��?Y\آ�G-�BD���l�%(����~�)JP�߾��R�[�ۄ��	зt1S�:eBZ���ͦըy�g��9#j�$c�9�v&W!,�}��\v��H�j�m@�$}�ߞ)J����R���{������S6L�L{޿8L�L�Y�^���+�F������┥{��y����������)?����%)N�^�8��d�����,m�[�[jj[A�)}��)JRw��a��'�(8jS��_g�(����<��?g��PŊ[X��Zv�$$OĒ
�;��my)J}���8�)C��c�J��>���)JO׽��f�V�n��Z޶���;�w��)J>EB�߶>JR��}���)I�{ݯ%(E<*I� ��Q�ZV�HT�=`��I��:�	�bʬ����)����Z���qO1�)�&Kd�(��#	D�����P�H��)oY	V�$�(H�#L�"`�$ �p1`�`Ą0�+�`�cWd�lc!���$�l�����J�d��&�`�����&��0�D!$&J�1�������{� (D�D��1=�?����&mmJ�fjU����0d�ۤ�j`-�x����z�^Y���	I���$�ttԓ�+�kT[/�1�*��a1�v�|޺����9TU��;(�ǫ�����.��1<
fv�v�k��t�=8-�yշ�(���Tű3��US���sr��u��z��vF�մ��U(ꦨ_:I�4Z�:cLsgc�Q0̜�jB맲�����Bql��gp�n6���廰�PYg�#Jksl��{�`��h���ΐB�A�oX��X����&�+�3�\Y��k\�I��FG2qXv����e�!'��]���Ӳ%��ێ1qɻ�m !�f]D���bJ݀ dn59v�KŸ�����,l�Zv�w �mF�0��M��k;�nm;j꽖�0�v�S�n��l�Wj��h���WU�z�5�΂2����J��N�v.&�(�v�3(��V�3h�k�l╶���]l�P@�ܨ��j��9�C��.�Er�*�P*k���.ͺHz�6��$��Mвp+�U*�UT�����WŴn]�(32�h�
W�<[B���m pke���K>�hH�H��	�yrj��ew`��r�	�-�o���K5h���'l`w`v�==�L�6��U]c
lcl�˧h:�ej���غ���<�ƳTIӷM�m��L�&^��+J�kj�-m�  �� �V����i�G+���Ѣٕ2� �ۗܛ��"i�*�B@4v�V�v
�j����B^+[r��m[*�R��$��\�=��qb@�b����/[�����W>�^��vvݭ� 8�^W�hu�	���[�yӀ��g<�j��р�8-{8��k��&��T �uc�u�H�g��}P"���!Hm±sݎ��L/G�:� �3������*�[�u8��+��_Wr�.E[�:�F%]նH8AB���ju6��Ȋ|g�߯(?�+���y���z�����707GJ5S�gm.�b 0�yc��������k�b�A��v�\�]�����׎m���:��h�N���P������Q�!�;gn�а�&ю	�&�{g�CY������j�(T��ZFUB.a�ڞ[�R�	��t�n��}�m���]MA����b��'7�6x�&��S�M�Øi9ߞ����w����q�'9룭p��t�q�&ۓ]��t�YۘWIe�` �#�1ڐ� �4Ul���R���ly)J]�{�)JRy�{��T�JS����)Jݳ���%]iK*R9A�HH��wn ?��	����R��￶���?�����R��ﶃ���$D�}��>����Z�����)I�����)���)O��I�{�ǒ����}��BD%	BP�&f	BP�%	�%	BP��%	BP�}����$�V䍺#��! B@�	By�%	BP�$BP�%	Bfb�BP�%	�%	BP�}���<��(J!(J��30J��(H��(J���(J��;�~��(J��<���(J!(J��30J��(H��(J�Ͼ�����%	BP�	BP�%	��P�%	BD%	BP�	��P�%	B~��q��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	 G~��|��Y\�Yl���$	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�{�	BP�%	�`�%	BP�	BP�%	��P�%	BD%*P�%	�}����(J��"��(J3�(J��J��(L���(J�����(J��0J��(H��(J���(J��"��(J����P�%	BD%	BP�&f	BP�%	�%	BP��%	BP��w������ffI����G3]��ѹ1:J[����@ ��?xs}́�cz������P�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�}����(J��"��(J3�(J��J��(L���(J�����(J��0J��(H��(J���(J��"��(J����P�%#BD%	BP�&f	BP�%	�%	BP��%	BP�'}��8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP����kfլ��f������J��(H��(J���(J��"��(J3�(J���~��(J��<���� 8X$#�T�!(J!(J��<���(J!(J��7���<�J��(H��(J���(J��"��(J3�(J��߾��(J��<���(J!(J��30J��(H��(J�Ͼ�����%	BP�	BP�%�0�X%	BP�$BP�%	Bf`�H�! G��材1j��천��(J��(J��"��(J3�(J��J��(O���g�	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP���p��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bg�}���J��(H��(J���(J��"��(J3�(J���~��(J��<���(J!(J��30J��(H��$H����ԅ�$El���(J��J��(L���(J%(J��30J��(N�߸pJ��(O3�(J��J��(L���(J!(J��3��~x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B~��q��%	BP�f	BP�%	�%	BP��%	BP�*NBD%	BP�'��?����(J��J��(L���(J!(J��30J��(K߬��_ټ�z�f��z�l��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bg�}���J��(H��(J���(J��"��(J3�(J���~��(J��<���(J!(J��30J��(H��(J�����y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�{�	BP�%	�`�%	BP�	BP�%	��P�%	BD"@��	w���Q%�D��� Q)MHuA=�l[:yi�u�Ƴ��)==pv<-�-�9,�dn5r�p�! B@��"��(J3�(J��J��(L���(J�����(J��0J��(H��(J���(J��"��(J����P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'{߸pJ��(O3�(J��J��(L���(J!(J��3��~x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B}ޟs-�Z�6�Zp�! B@��x%	BP�$BP�%	Bf`�%	BP�	BP�%	������(J��"��(J3�(J��J��(L���(J���8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP���}�<��(J!(J��30J��(H��(J���(J��?}��x%	BP�'��P�%	A���%	BP����(J!(J��=������k������B@��	$BP�%	Bf`�%	BP�	BP�%	��P�%	B}���8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP����~x%	BP�$BP�%	Bf`�%$� ��J��(J��`�%	BP������(J��(J��(J��(L���(J��(J�����y��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	B$����9c�P�[.$P�'��P�%	BP�%	BP��%	BP�%	BP�%	�}����(J��(J��(L���(J��(J���(J��?}��8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	�����P�%	BP�%	BP��%	BP�%	BP��9=�~��q I	 H>~��B(��mi�{� � Ѓ�{݈<���J�������(J��(J��(L���(J��(J���(J��;���	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	Bg�w����%	BP�%	BP�&f	BP�%	BP�%	Bf`�%$ߧ�E�4J���ltE/�N�j9�yكTp[v��ؕ�:���灞)#Ij��e�`! B@��	8�!!(J��(J��30J��(J��(J�߳��(J��(J��30J��(J��(J3�(J��{�8%	BP�'��P�%	BP�%	Id%���|�����ly	Bw��{�փ�&�+mxH������.���P��w�����u�s�|-�|�/�m;����b(K���%	I�{ݏ >X�O��~xH���#! F���6K�L�e����(~�$���ly	B}���pJ��}�Ӑ�@�+b��7�BD���6�c���n5D�����;�{�┥����c�)}�~�		#��I�HH���S��%�Ը+k\/MV���k��(tkJ�tvk��8WaA�d�=]QG#5G��m�v�=���y)J]���)<�{�䤉���!"9�f�S�)jr�޶<��.���|�NJR~��my)J}���qJR����c�JS�~�mX��%b�+-�BD����i8�)N�^�8�)I��{��)w��|HH��]�zӡ�%��[�T"B��u�s�R������R���{�(�!"7�5���#v?k���7o{�qJR����JR�{�w�)JO;�v���;�{�┥&����J��(�������ޭ������;lk��nQVh���tt۶kG����l�Kl��k���==�K��a�3����Ϧa��Mt��76n�]x^u�����I0�����G����6�FT�[��Y�DF�M��ʍ�p.˝�:�Ǝ����6嫢�J����v�s������f�p]��v�)mɬh�a�pH��֣&I�m7�quý�{ϻ���ﾰ�������Q��z�[��[i��ۋgB<)n�)�i��<C���q�c���BD�����BD����a�)�����@ً�JO���D��t�r}-P7\b5�		)I�{���JS�׽�)JRw��È��!n�n$$Gz=�㪷X�o�{����{�{�R���{ݏ%)K���┥'{�vJR�t�.�,��[K,��!"BDn��q)J]���);���R��u�^$$G��h�8�V�-�K(8�)K���┥'{�vJR���p��!"7wh8�	9�vX]��c����8�H��2�h9��.�����6���H(����L�#�~�-�����-�t޳@�{�T)����H�Rf�k굤w�w@-�h^���$}_�蚈�1�2~mŠ^�n�[�h^�����xU2��F~ ���@����/>�@�z�{�D�r��$ӓ@����-}V���� ���<���$М0�"`]v{r�-�=�$���b]ݗnE�ףqu��N��ZS#QD�	��I����;޻�������+�s�GU�w�͈����z���F ����,����$q<y#�oY�y{pb`�|I�d��I{��ė{5m
�&9��rh^�����;޻�������119H�Rf�k�����f��빠\G��S$�:��uj
on�̰����N�w-���F�V_K��25�5�cBd�ۋ@�z�[�h^�����xEj��F�A���������h�w~���#�����D5iɠ{��nh��@�z�[�h�tV4�ɂ�HQ��[��`�� o�`d��?/-��{�J�F��I(�qȴ�ט �Z�8��0ﮰ���������(�����xe�ztŻ;z����mM�(z\jф3�X]��Ë�f癿@�V�ב�:m�ߺ� ��Ơ�Ƈ�"94/Jh^�@�z� �Y�1T}�w{E(�*�(J���kwo ��y��Q�����0
�Ꚉ��d�8��;�w@-�hޔ�-v� �V��$��8D��m���4]�@�m���((Iۡ|V��i	PnևMմ�:wnLۙ�}�6��I��j�|g\�θ�r;nS��	:]�9d�"���e����\S�FC	���7�-l��^��-�DE9y�uß�W���*�9%�
�bع'�8����j#`g�Ӣ^��m�%��k��i���4��O3�:�����y�hg�c�7!��f�gVd�T`�A-��(iI� �4�3';Z��W�A�<�mc�:l`���u�v�ƺ���ֵr�Xs�kd��Q�>|�_U�^�oY�{�EcNH,�7ȤZ���/[�߿~����}_�-ۇJ�F��PDqȴm����s�h��@��ˏ"c��q<l�h�f���Z���=����1A�D�#�#�@�v������ ���>��ٟ����u�f[�[�l���jr��lI����n�Ah;6;0sm�u5R�.-Ƥ�qx����/[�oY�^v������Fjc������ ���<�)�Uz� �V����mEs@-�4/Jh^�@�z�{�Dݒ �?4�ӓ@����U������f�������8H�!�Uz���oY�yzS@�g�;��3�n+K�6��h�����泰V3̜��M�a��Rr�zI26�B��Z��d��>�� }�XS=��ݼߏ���By$q�`�m�@����U���]�<�����#�Vۉ.o�$����� ��@B�,D�0$0���xU�#Sh���7�v��d"J��y�-��b	�j�&@�A@����!���l6��ȍp(�t���D5�·����:@��;�0D^�Ї�8����C�D^��EL� �	d�0pz��mĒ�}�@����)��Ha#�9�Vנ�Y��4/]���M�d�9#����z���sO�/���������|7h�j
�����gM�E)Wn���cy����5g�<�\��i" ^ʪ�v��V�Հk���|���k@��Dݎ$E1 �&�yڴ
����f�^�48�m�O�$��iF ��� ;޵���Q���>�������H�!�'#��@z� �L�#"b"`w�w�8�ln	�0RI���4�ՠU�@/[4=�[i�d��#"���)p'N��U/m��-Ф�5Xoc
8�Nr��6�7XB94/Jh{k�����f�篛�S��H�^����4�Y�yzS@���"bQ��Lcr= �z� �l�/;V�WZ��#��!Li6�q�4��@��Z]k�����v8�Ƥ��j�*�� ���]�{�T�+x&������s����Cp��ܗmhȝ�S����4n��ݞF.��<8���cNuй)��ZO����c"k����#�:;�lm���}�Ev�s�v��v��&�e�m�X�ۚk�7e�V몥�9���;Ѹ86�+W�r�֖�\/'Q�n�0u��rQ����:Άmm�&_o|<"<d5�kY��S�����ߋ�����y�77&�.$�U@���0[�O`χ�p��ӆ��l%-�����N/@��|���@-�h��@��*�8�C��X�@[X �k m�`�w�v7��Qp��.RIpwu`��ӵ����],�&48E�$�@�۹�Umz.���f�篛�S"jn5&h[^�˺� �٠[e4�V�6݆/�H�6�Nֵ�8X��n^u����\���!���7Bb�q����Li�Lcr=�k����)�Uֽ �#��!O�4�q�4������� D�"��s\����= �٠[��nǑ"d���&�m��*�^�[l����:+nA� �G1W�@m���wt�@�nJ�G�5`�X܏@-�h�f�m��*�^��u�x�Oz��E�s�M�/;�t���(���4,�m�v�ɭ����!���wݱ�T��b����,����z� ;޵�w�cAjc�B
I�ym��*�@;�� ��4=|�B��Cy ܊Lڻ���r��}��mM"2�"
4�E,A"���w��|���s@���DL#x�c��wY��f��s@��� ��V��mD�rh�٠ym��/t����mēt��A�,U�,n�-rn�Қ�U�-���6��\�Z^�l(v��{cclV���nG�P'�!�'�ym��-�M ��4޳@�s���#��1�BҌ��`{ְ���c�n�F��d�L�2<�2I ��4���q���7�����ldE�-E\ ���z���X۫L�����p�@�f�Iw�VԬ��m��NI�yl��Wuz��h�٠T~~r���]��u%�k�/����6�/f)���nij+]6O&�1##r�(�w����X���f&9A���`��"`�	�&A9�wu�{��<��h�)�$�>k�F��������h[w4zS@;������4O�DNM�n�}����h�@�s����)�c�4���@/u�����Da�� � ,� k�m���oR82;"J�l�f�᳍WV��$.ťw�vƌ.ʘmۛ��sY7:=�PLS�tr 1��K�i�gOXG�+�m��B��=�[��F�,n;kt��=�y� �TX�6�s����mV�ª���l��V�MV0d� ��i��/��N�٦'����fն�9J�;;\U;Xێd���[8����}����.e�}�{�8��^��K��Z�zZ���Sm�Ӎ�QC��s@�E�Ѯ}f��]�5�H��'$8޿M ��h[)�?�f�n�ldE�-E\ ������<�S@�۹��f���\Dm���r�ܚ��h�w4�٠����5P��i'�q8h�w4����f�岚�+�Ja1�L���� ��4�Y�yl��}빠{��cu�I�� ���I��k��M�[�l�8z�q1wI�h�XL�T�:dh�V,�x�cRM �����h��hwY�[���Pd�2bH�ɠyl������o������Y�w��Xܑ�r1� �4
�������Y�yl��s��T�9�d$z��h�@��M�mz�nl(*.mJ�\ ��`m3 ��^�wu�����_�$J8�E\�ќR�E'z�
��1;m�������9�86Lo��"�M�n�W�����^�4��B��7��W�����^�4l��y���BL�ĜZm�@/u�2fb'�D��{���>�0��*�QdM��5$��f�m��|��l�DUn�^��$�]EšCY�@��h{k�m�{��o���q���f����5���5�]d����%���8�nn�R���'��M�@��^�[l�oY�[e4�{%R�ň�rC@-�h�k m�`�3 ��l(����������Հ6�0���6�F⥡d��I9�h�Mަ`�����r&%��LNegZ�:�n�5��'�[Қ��h���)�_ݝt$ddR,�c���ݶ��]F"�4���m�5��W-؜l�G��q�L#���h۹��4�g�9A��L q�N�iT(������(��Y�Tn�� �զ �y��e�#��G$�-��m3���������Հw�ꦮ��DR.*)�`~���0��`m�L��M}���a�[IZ�P+JҴ`{ְ����F �L��PHFVa�7��Om���F�D�^��0]��\;� ��h%�	��"���� �>@ƏqE�l=S�K�`	� 9"`�3) ��a�"qd%�&�7 XQ �A�J�s'�#1�F[D��1c��$bYaCh�h$f�1��b�#Y�5Eh4ɚ*��ԅ�����D�H�dٸ�	m�`H�#�$p<M.c@c)�a ZQؕ��!�3`��'���D=6r]aD:�J�BP!���&`YJ��HYS��afY1��E4Xe��f;�تh�"5�A���'p�&	Iq11��jl0#��'0�B)@,�( <��j�d��Up�^ݡ�D0d�{o	�:�^��)�!�<k�^�b���v�Exr[J�kuY��ŭ�S�_]<8��n{eD;`��]pvi��[�<Wt�CXs����;Q��ۋ�iǰ'D">8�lhRc`ƺ�b�,�;��`�8;\�ű\p*�-U&YUl�8����@�0Jh���N�TcUTR��,-+�걅���:961s�X"ڞ�2����ۮ�o\@N
�����qCh�ڳ:K#�	m+�AZ���êKetph���Kt�i�Tq�C�3+,P��pW7]]+6R�V;i����B�5m[v4�X��>�6��;�Oڜ���.g��[hv��]�x�b�q��չ���we��ǈ�ޫj	1�]'���:����MCVЇ6�a�A�rŵ��N��U���Nևyqtc&uu�=�˻��)�s�4�.����t�pH�D�ܝ�`v�D��c���Z�Z(Z�m����]l6*�0�*��֡Ֆ\-ˊ6ۂ[(�t:+�%�Up�P�GD��B-˵΋��mm륺����$�[��v��j�\YvW�`�@�h�h(r�*��-��fl�:�㑪����j�u�µrB�7W6*�Zt�tѷ$�N6�8�b�PUpj�*��t�	��hO` �)v ��kW8�D�3g�u�niZ��v�`x�n)溥k��53�.��V�m����6Ͱ��f �C[�-n�;��vϛ���Ve�:�s�lR���a�jNѹlvtN��jV�Oh�ض��[j��հS�4v���''�:��eV�(j���[��ms�������Ų��-j�
�  c�����>����cb��4���:d[�D�ފ7l܎��l�ku����샐�����6
��W!�ٱO�mb�������եZ}m*�\f�5n�P{=ݣ���\��<n�i-o37��-�=�)���@S㐒@��  2��У�����ٓ^���j7�9μgs�m�u�3'b;P �cSu78�;r:�*���f�����e��1ڝ˹���P�����ئ���U�퉜<{f1n��uڳ��%���깧��y 
����k�<Z�A�GM�[��+9ɶ��r�b�r��&�L�*۫j����!�mk�\�9ܽ�Gnݜn�cB�v�D7a�gD�ژ�\W�PF�jݘ�Z�{^��z�T�ev�j��NW�� �e��8�$�����8���:��鉉��m�h�����5�Hc�9&��s@�Қ��h[f����#�կ�y�sqI�����f�u�4l����q�L�MDbn11[�� ;�V �L�و�}�� ���&#1'&�{z��)�u�M �٠�g>��m�m�� ۞e��4t�*�Z�g9��X�n���fOiʥ��I�+*U��eTRI|��� �\��[l�oY�w��X�s�p�y�5�ܫ�����@�@�D��ԃwu`�� m�g�f�p�-���&,�!8���h[f�m��9[^�n���5�F���O ����v�w���Sls%25��S@�ڴ�f�[l�.+��&�4�ۘ��Y�q�{L���U��nݞ*�˱wn�W*���B��pn�ՠ�4�g��n�F���VU()@]Ҳ.�V w�k6ff&�7wV���`�w�s���q4?<pĤ�m�@�۹� AD����Ù�{�K��q%�զ	YR��WWP�%�����0�ߞ�wu�m�@�s����̊1ビ4
�נ�f�[l�<��hm����=����qP��g%�t#���3���d�e��i z ���:q�tr����M�� ��4�f��s@�ڴ��Ȋ�VXX$���Հq۹�Z�� ��4:�lsh��WUi`m�`�u��&&"�m�����y���F�Pl�M�&h|��v��� >m�bb"�LLL�F��>�1)�����JE��f�u��6�0�n�������
�%X�mD�#�=yÓ�a��nNݩ�m��mGg���J1���;�c=��H�k��ߟ���h[w4Vנ�f�nR�~R,�e����Fl���U�v��D�E��ﾚ{��7QǄ�&h��@;�� �l�<��hnJ�����	#��@:�4-��+����왯c֒ H��׫ �o# �>����`3�	�U�F�i�7[7�-i�W`�唟`��A��n���vt��^2�������jѥ���Y����j��,;*(9uGfӱ�Y᳇i��4�U�6�Y�7'Ee�4NTkU���8�emt��g�D8�;f� ng�9�a�X��3��pUutE���q\m�˷c����v�^I�6�=Y��:�>���h1�f��dd�ͬ]8�H�)p'5��=���P@7�ĝ�͈`�qصm.n��u����[w4W���@:����P�H�##M�&h�W�߿f~H-�M �_���s@�}\bSS'�wu�׬��ߒ�̀w;V���I����ě����{m��}����� ��4�R�d`��-$�6�0�����oV ym��֢<X�!&9��q)��T瞸z卸�R��/fɺSq�ā�2�&H.-�`��� ;޵�}k�13��þ��0��z���+�I]��^ w�k*b�8�Xyk�w�13T7���\e�^]UIp�������ޯ@;�ũ$��R����btT�r�q�����g��{7�8�o�RjI%�y�Iz�'B8�0�"Q�hX�o�۳�m��n������}yĒ�ٸjI.�\��B~R�I��k]�.�k�n_Z���	<V�@�uR�����3[���F7�8��$�t�jI%׬�������H����9��^��+PV����'"ԒK�Y�%�pԒ\�w�UUWz���1�IU{���t���[�[o8�{�����ߦ��q���@�)�ũ$����%ݎ'[M�Epra�/��v}���I[>�RI.��<I/m�����sj������xG�$��-I%�c��{�Iw�M�RIs�_�$�s��9�n���	�b���榑��D����F�P<����C>6]�}�|�p=��I�$�����x�^�7I%ϭ����ZI[>�RIs�/�F���)�W\��m���?�@�k{3�8�ov�^6�}���|A G�-�\���Y$�I�(�I%������I.�bԒK�l�Ē�ٸjI/}��!Lp$Ҳ�q��"M���m����^q���p,m�'I@��e���q���nI�A\e�dK^6�}���6��{ﳁq�޻���H]��Kܷ6�7�a���FWW(]O�饉���;�`�hr"s���R�g3��W9�����������s������$m���^q��D�}��NLI�Ɇ����W�$.���|���o���Ē I���֒�+P��Cr�q����\m�����?�$$��\m�{�8�~��8���]]��%k�U�&.�۾\�UWwVA��{;�9���H�n�.6����ꕑ)B�Si�y���������~ ٿ~��m��ߥ��o{��m��#��@d�N�k� o�I����Ėݺ`��\v�{i�!�L��L��Hc����^��]j��1���K�Y7\�mϯ���]a���i�Nvj��*"{tT�v���Ru���K�qN6�=J��sN���,՟�q��*&��԰�J
��^���Л%u��s�HP��6�.n�eӷ
��I��
�Yv]B�ޛ~L|�����3��#n^7�\�ִn*ݺ�W8�s�+�^��a��m���]�v� ����_�wW5$���?�~��}i.�馁y���\+�j���Y舉����=�|h{����٘�u)�Q3qcn= ���@�S@��� ����cS�L��4;�4
���w�`l�MV�Հ6�mZ��H�V�$��*�נwY�޳@�S����~�v��v+�<��=v���0�݈'��g9�۶��Ft���T���yn��;t�	ZJ
�| ��X �m`�S=������{�Pe�yI()$��w����IEB������X��o 9޵��&��wkP+��EER�U��>mi�:����MQ�z�{~���u���F��C@�ޯ@9޵��k�1����<`�ߑB��?GHn= �� ����Қ^�z�g�ٝ�~x��Cs ۅR�������'Y']�I�5ۧ%$
gh�C�˺3Z��)��������hwJh{����h��Y�L��8F��9ަf�]{x�z��z�`ܟ'JA�&'��W�^�y�g/�tz� iIX4�w?y��b�� x����䓆"*h��}�?y��&ҡ���P�����̊��V��-���ō�XN&YdN9����2�K
0#2�Z��ZӚ�2j��,1���̰�7;�� �n�`�v���̲�,�"�k,����(?~�kd	�J���x�x��<WB�� ��z��D��Ԑ������_�{�܂�J�(&�BD�17�y�f�_z���M�z�����bĵ��Wh�I. o^��3�y� ����wY�{z�2A��E&�D1H�`��U�Vp���,lP����vU����1bS ����Қ^����4�Y�x�7Q�~�di��4
���.���Y�y�)�r����1� �&9���@�mz�Қ+k�<��ej#&)���@�mz;�����LFL' �13��ŀyr��?$s	#�<��9^��w�`��x���l�!TSC�s�Jf�O�͞Wu�=sT6\����]J��P��=p�o������;��=W��<��;;�T��HH��ӏ@<�@�^�@�S@��@���1b�fq�&
I<���y�)�r�נwY��
����H��&ӏC�����~4
��= ��4�^��ۺ���!B��V��v�]������� �^���3 � �S�}��j0�V�V�rO�1��ڄ���94n���.��y=����p�jz���i�k�VF�sƺ�t�j] ��˃΍G].�r
��������.��;���n3�1V��s�V��Y(�)#t�0i��v^��m��l[k>�[<o9��qv�^�WJ��p�kQ�3X��Ѷ��ˬd!��;�v��s'R��p��u��6;���n�tΎb�;R.[L��`�4��\�y�X��dv��N�.�]nz��#'�����
���� �>��9ަz"y@����hg�Dd�?!�q��W�y�)�v�w�r��y��<�DyAjj��ըW�wux�;M��=[{|���߸�8�R�q��_�|�߾�h��@�:����Ț��$�@<�� �٠y�Z�ջo���w��xm/Er��.�j���&k�>�W�۱ґ�ɎZǲ<�����q���򼤒����9ޫu�7m� q���={R�*�M�,J�q%�z�y�GA�H�R����]�y����{�U[l�<������Q�I��@��X����F���>m^��w�N(�	�2O�jE�[f�^�hwK��k[��ݲ5+]
.һ�x �ְ�7���mwv���x+���ޚz�A�<�b�4ql�����#��/X�{N��MJg�g�<kWf�l�6���y�,Z]k�=V����~��O��� �G�dNAh��h�k����ۋ@��.���ԓ��7�궽 �l�;�Qhu�@��]�\T`$
.I_�^�y`��VWZ�?��?������Ƣ�L��@�}E�Uֽ�mzzـl���Í�̀H�Quj��H)3�yΒ�z������l�^�#��"�匿��'Ƒ�$F��8��}������f��tuh/y��S��b�@�[^�^�hwGV�WZ���fbA��3>���LnF�z���y�Z%�|�W�|���,�0I�n��9ޫu�:�w�r�w��Dzb&l�@�� ��}>�ė{���;R��h�-�k�<Vנ�4;��v���x���0�qP�:���T�w���~��Ng�2j��[�=��e㤓����u�4%%|�����k �z��L��=^�� ���ȸ���B���W�{� �X�
�נz��{3?�6r���<lpm�E�r�����@;߬�<����1�~q��-���Sn�6fb�o5V�n��E(N�`���=Vנ��@�X�WZ���:a���Y�n	K82�;�ɜ
�!�Gk�Le�7Jl;>km<g=s�fxZ�6���b��2β��n^-]��n���r��cm�s�v�s/[.��v�\/l�
N.�#)��q�����v7N��r�=C���5�T�͎�֮UY�Zg�:=��f��d�s�.�K��P�ٳ���m��лn� Uj���պ:u/:ͽ�ww�ُ��k��n��G�=we%6f�͗͌86��ض���v]���ޚN��s�o7#n?@/��y�,Z���U����X5�p�@�X�U���k��f���f$^��8ƢP$��IV�����k�3T;��@���Z�ݗT�D9�����������E���������5X�����.*r����$� 7wV��5X���͵�~��}�7�5��+��ͳ�F�<��Ϫ�etڕ�ng�[u��0��������Ӓ�1�����wuyV ���6� m`o�B4�Hc���h[^��?f}�&%!�o/ 7wV��5X+��e�<�$F(7�궽 �٠y���
��@;�Yd�1�/�Ez��#�~������x���8��w}�@��B��Hx�NM�uנz"&c�3^���6��� m��:>�?9#�sqz��p�\���mu�@^�1lm�a���M]�/c�N�Fr]tv�.��WZ���h�@����DJ���
K1$��۟Amެ�n�`�n������.�
��Ip[Հr��kٙ�����r�#��4'��T�Ms�]���~X~�4
�J�QT�+�@�w;4
����٠����[ue��+��J��|�����DDGW���۾X+���;�e�!%q��]�F�.�9�Pd�̥��ַ0ۜs3vI.1qj��,3���~~~8 �ְW{ml�(6��x �V�j���4�2Gz{��<]���mx)�y鉚�v�B��e\U�B���7z�_7xzb"�����oV��u�L�L$�qI&�W���k� }m`r"b933N�J�ޥ�|�}�c�H(���q��k��f���h�j�2ڄ�C�Mq�&t��f����D�Y���ȇ�4<%i{"m�(��"�!T�]
�W��|�W{m`�n�DDr�����oMAJ�R��U$
��?���z���k 8�X �ֳ�15G�l�ue��+��J��>���@<�� ��h.�f���i��\$Z,�Wh��DU}�� 5����X���{�� }+j5\(�����94��@�w;4�]� ��9V���&
��Ph:�I8:�Ц?�i�;��a9?�� <�	�Ċ�t�b���m4��`$���02���;x��0АL�a�L ��Y�fa��f&aX@ؘa��E�d���bM�Af66f$QfLNAY�YdņDD�7 �����l� �R�+v�@[T6H�\���o㍫n3����\��W��6J�y�!�ѻɸ�̣���.6�un���,�4JX���u�#�*�qe �݌�'Y2T�;#�[App��ax�Vۭ԰E�B��vF�n:J*��U�!��MU#3���:6z���5���v��i�r�ܔ(�zS���R�1��y�du�nζ���l 5�kO�4�clBx9��n{�p`�(P�n�L]��c�F#�Я<�u��2�WT�m��ymt�T��ó�ؙ�a�܎M^�\�P(�i�d�[Jv�rI�4$$����WJ[/n��f��@���lW�JȞ��\����l���sT礓�mu��'M��nnn�j�r�O3�+���M�&��m��k�l�&��B��vݐ-E`{o��z�pd�xub!6ݭ�rT��h��Jv�l��S�6c��V�@��ڣt�c]9���[N��nmU��P�ā��Nӄ�m����%uc �#uppͪڬ���F����+��ʂ�5[�6� [[�KVY�h%��\EHN}�<.Ͷ��s�6�r�5Um���[���)�
�t�5�^�*�e9Z�usN&xs�ZM�nI�F�qml�T :AY4m�/���`�my%���aj�Y�l�R��v1Ԭ�R� �{<g��i�=+J��%��;S7n�{lֺ�U+�������|K -����l����V\�.'�*�$3�g1�݅ZN��ږDݶ9��눴�ngR���g��v�vVڥ��ml�Kc\�8%l�p�G6{K���̪���jy��WD�8��Q;����s�sʸ�,UV�i+c��4�v7MjK�q=D��:9N:����p5���dO4S�+���
A���p7bL��ru�c�a/nɛ���\/ob0w=l荗��  J�Fٽ1���쒼�(=u�y�4�<��Q�Vz��Gj~�?hM��PC��V6G�U�Oz�� @ �C����qJ�%��]A�m�;�Q��]^�gq@�S��q��q�.�ɴ0��Z7����n8�kDc�/g�G��ZJ)�vn�j]q���C%�kt�
�C��)���;�� �TY��;��'�'m\p�u�mandf�B�ң��gu���
R��J�՘Nǳ[I�Z��۷�{u�]����pfr��S�����s]N������.��,m=��Hb�����; z7��Yk�&bծ�.��5_m����# 8�[�z�`�_���s�ǉ�Grh�)�[f�^�4s�~���1#�s�S��(�z�������٠[јl�����ª���$���&&j����>��V �S02'�DLE��v��O�(�2���$���٠g�<Ӏ}[�x �Z�5贊��Wv���Xۇć]V񛇆�n�x�ט��s�:
����ݾ�_�#�[�E��{o����)�x �Z�����n�`Sw_�V	E�\�bK�wft�� x��9_v��Zfzfbj���MO&,M%�ȣ�@>�}4s�@�e4��ūI	�cLG�94W{m`�3 �6�ff*�����?�dƇRE��)�[f�_m���٠e�����~��1&�KV�V���r���H�pLmLJI��_��b�̥	Z�I\U�� w�������m�LL�r�u�0�?{�qQ�$��4�< ����<]��ޔ�-���#�@Q�d�$�>��V ���11Tq����`+��F��?H�nG&�k��l��@�w;4���)�I�E#�-�@-�h.�f�U����߿���}�u�Z�̄L;��̈́�y�&�۬$�d}��U��u���E.���H��z�����*�^�ⶽ�-ZHL��`��$���٠Umz����f���u�O�jbJ���:m��m��j��Հ}]w��/��TǒBHG��h.��m���m�L�FD+x�X_O�ȸ��.�(U`�%| ��X+��X�S@�u�@<�cx� �%"�ˊ3�Vx*J����P�����a�F��3�
�@Q�b�N@nM��;4]�@�u�@-�h+��F��̍2��ZXm3=3135A��X�����߿g�V��!L�L$�(ㆁ�=���Xl�W��z��Z`S�����-	ZX1U������h�M ��yB�D��J
�,��m�b7w4�Sݼ m��m M�� ��=��^�s�~m<Z��q�;��vt
��#:��73��W9�/c�av]�mۧ���닮���킱mM��h��	��6�H�b�P\->vglG,Ӥ�}���Xū�l������MIػnݪ��fǲڧp�n����k�ԑ� lҵ�3	��K����������k���T.���b���;�u�(�q�;�]��i4-��C��l4�h`[�{)D��E���tzd�y��!:m<�cv�r�X�ʘ��Q�Hܜ����<]k�m���vh=캢Fӊ(�iH�Z��f������ՠu��y�5�rCNG��}��<^�@�ڴZ��X
cS��rB94���-v��ֽ �٠x�7Qf724�ێM�j�<]k�m���vh=MȢq�	7;-��Spzz��H�O1��sj�6Gf�G^�c[��&��)�I�E�h.������;4]�@<�������,rf��r�����2O��� kv���h|��@�u�@�/(XH�I<piɠx��f�oJh.���f���u�LpH���ܚ���:٠����vh;��pM�9#R- �oY�x��f�oJh�s�Ҍ$"�$xМ�1�-E�S���q�]J�6鴝;BN�;^�b����n��`�I�I��_�������)�u�@�{U��52(��rM��ZY蚣]��i�� ?�X+���i��Ƙ�rI�^}V�WZ��y3;�y��Հv�z���n�QJ�ME�hu�@-�4�f�k�ˊ�LPi$Ȥrh�f��������=]k�<^��yg9�c�u���浬�$_�/d�ƗlTӸy�gZ�.�=��5���~������<]k�z��GSU�b�X�Q8ܚ��۟��_|��_�$���/����[��hQ9k��[�@=��M ���<^�@��ZV~�EЪ2)R���i.�bb#�������s�k�|��׽�W�T:ʀ �	� �$[72�K������2F�p�M��;4_U�u�@�X�b&\n��
�]�Wi+P�ʖ��rN���h����6G��+�{eZY��y�����H���m�'�?���y�� ���<^�@�w5q
dn&���H�ζh�f�������߳�_|�DdM#�7&�}��h.�f�k��l�/��,�$�c�94s�@��Z�h}������;���ͬS#m�N6��@��Z�h�f���vh���nG�����=���h�rђ��f�eR6�H�ݹ��(;"ֳ��8����hM��Y�9����.t^�әzC�7,s��/���q�wҳX�H��Ƴ��S̓��AVG+Y���C��"�g+�=<��ݚ����U������vl{��i]���m�:���:EWFD���"����i5�%��:)�l�����5�R��r�� �1:�s
Uv�q�L����U?�}��?Z������RѺ�Ӻ��1�Q#�J9#qp����X+���DDO(7m�`���"��U��m�J9'�w�M����/>�@<����V��d���94u��7}u��bf*��u`�Հr�j�F�P�F�7#�@��Z�h�f���vh.�!LQ��Pq�� 8�X�bb#�13~��|kv��
�W�u��M:�y�E1��V�c�b׵^��f읰��a���5عJ K�F�cqF��z�����*�^�ym��8��P�'rh.�w|��p��4����0AU�F��Q��W��f"b3�v�� =z����������6�L����ҎM��h�٧߱#���z�M�K�"BG�4ےڬ��DL�_W���{|�W{m`��@�����X��q�6�#�x�}��<W����h�j�;�+�'q�K�6ͳ�X�f01l������v.دu�q�������}m9�,��<��M���h���<�án,���#�@���@��V�_z��yٿ~���˫_b�n:E��� ���`��a���LNIç� L6`�;m%� H�f�O�$C$�M�L!2+�
>)����xPRH�x�>/�0��Eo~
/-p�HQBS2D�)�EMƳ"DS�m z�mTz@�
.x��Q��O�?��0xAO��������Ē�^��EDY&E"��Y�x�;4��6&kz�k ����UUV�i,�y٠__U�_]�@/�f��W�����sqϩ�J�L5
&sL我9iI�^�0��v\x#��#)�қW@*\{ok [u����ծ�`_��E�$F'$ȜZ�ڴ��h+���������1b�zE��ZU��Հr�m�=[�{X���o�=]��cNA8�nI��f~^���hs�-��Z�%}�49��F��#q�m���/���?�g�>�x�_�����<�5[��#򐏐mQ�ic��g�i�b6�.뱙+� ��;�u3f�S�(�q�8ԋ@��V�_z��y٠__U��,l�Q�Y"�����g�=v�y`w���޷�ٟ�f$}�H}��rM ��__U�x����Y�{�:�fLM�Y&D�rhb���h�~z{��;�4iuE�G��ܘۋ@���x���\ �� ��� ����
J��C���'nF��7l\�ڎM�J�cI�v�庻��Zm[eyA��0Ʌ�	!��)�&�ݸX�����t��#�<�8�.};js�z����Y9�16˹/-�Oq�!�<�;l{�N�75p5--� ד/�f�֗\e���u����7SGV��k�N�J�`8:YA�9,pF,�/[dk���7{�.ٞx���+�l����ɼ���ήn"�W7jneZ�lP�~ f3�5���T7.�r�꭬ݻp�mVrZuq5�y4�����l����7 � (�q�����@�w;4�������=]���9�1�crh��f�WZ����Y�{]�y�on94
�W�yO��ٚ�wu`��V��n�J)Zn5#�<W��������*�� ���"##x�E$zm� ��z�����}w�s�۔��u]GX(db�h�ٻr�1��*��݁6{d��m�8���9ԑ���Ù��߳��l�*�^��^�^�h񎦲��T���1%�۳0  �TLDG�;3�v�6��u`w��0�����#��ܘ��@�^�@/u�&&����`]ݼ�u�ȸ��H)]YJի�~����=��;�[��:���uz��TQ�8D�JI�{�+��U�@�wW�޳@/��p�U3n��X���pF��|�N�. �E˶�h���d�`�}�{���g�nn��T� ����8ﮰ�ֿL��u� �u���b��$�#�<��߿g��T�Հv��X���z&"bj�{�"27�!$�E�}��@�w;41$���!��g�s\�����ʼ�솮�WI]�i,�����z�]~z��Z}�4s�ST2cO"��,��w�z&&&~����z�x빠e��|�#d��NbO&D�ʳ���6Z7T�7a������b�0��j"N9&��m�����h���=�F ������E�M�*UV�*��ug阉��>�[��k���?����4�y��1'�D�h�Mߪ�s@���>�ߒ���- ���@�j�6�R�B���ؘ�LLD_�o� ��`Ww��x�� C��ID�p	ECP�C S��gs�f��>n��I�5"�/���=�z��u� _]`~n�"�z�b��q��ps�ʻμ%ћv�3�F�e��pne�;��	3$�kV+ ue��$��呂yyY�^}V�W�^��8���	�Iܚ��@����z� ��4r��^16���6��o��_u���LDLE��X ���4���N9&��mŠU�W�����<�D�ַ�`�k��\��¥QVUڵ| �����Lw]o#�}���w?{�r����3}����~������:��Ƴ���B� ��&�\�Z�<��� �{k��ւ�M�9��%V�+`�:�P9qmg�����Y�u�;Cg�sm2�%��s�q��0�v���,�p�G���]���ҧ���� �3Vx�@mn��U�p㳕�g�6[�$E��x���c�u��J�+ccoQw��}���n�A�}l%����V*��Ċ��I#T<&��Dh�:�8��C[[����)��)5�<;k��GmZ��h�&v����r0D�6������}�wN�e�VZR�Q�7}u�?�"&.�S�^ {��|�O#& v�v�QHH�M(ԋ@�ޯ@-�4�����h�WH�M�Hԑ��٠{O�� �w��[}{x�`�³rL�@�^vhwW�U�W��f���Y��یpI�&��7������Jm��$h�z^�s����g�X�JDA���*�@�ޯ@/�ϿL��r0�{�����.˻Quv� �ޯnL����٠yy]�������B��h��Tj��{���i�i���|���.�=�^sv/�4��V�鈉���F��� ���z��u���ӌIBF�@��z^�zoY��Vh֒
����\�&��B���j�A�x�g�e�݀�]�9����޳��f�ڦ7�˯�@-�4��˞ /W /��F��m�E$z��yޮ��*�^�W�^���$^ϾZE��$Ӓa5��߻�o�w;�u��� J�hS��ْ%�^�_m���S��i�!+��� u޻�}�x �Z���bm�k�F��e*�J�컵v� u�W��f���w4
���Op�\jոb\cr\��jZ�岶��W*�З;s۞coXqF��o��6��:L��m����@��]��{��g��
�즸,n�n$��{�? @mk��b�}���@��18!�i��*�@��^�_m�����=]Σ#�AƓ�8�>�ٟ�/�}�����8�O#�L�ʈ.M�����M���_U#��Iq��٠yy]����
���{J�z�!6I�Q,ݦWD�/0m6��cy%�[���Ɏ�P"S�j<��$�
94/+��Z�]��n�3<�7�� ���^�S��m�4
���*�נ�f�yyY�_J���q��ۍG�k�� ͬ6bfbb���z������R��uU����Հ}�4
���*�נy��X)�8d�1��M�y٠U�^�W�� ��4���y�$ת���#���N�8q|�L���΁0"?�e����&?�<3j�X�I$�2��$tB8��0�M'�hM&�v��a��噕�~0dca4������`d�a�A���E�aF0�]�
E(z7�[֍�q=�7�܀zH�H��O�gfX*�j�i��,RYr���*Iz��ԷN���b8gYѕ޳�]fۊ܆�[[�N�vN�6��h�.����$G;b�gp��4l]���C���]Z�l�p!]�g�Jvc���v9'p(t�֒ǔ��Aη�sK�8!]��[��ɠ��FKeJSN��k������m������T�U��8�A��N��`���=�A�:�Vk���MsFs���n3���͹6#-�W&n�	E���G���3���P�`r�Cm��9�+!b;*ٖ1�N��Xs"�.�L��W j�%AI�έ�u��
X#n��K/'1�-�1q���Fv��Ϙ  �!�۶2<E�*분�k`����yŒ�]nqT��ةP�����S������{b�+�n�i�R�V�aY���$2���I0��6i#[\,��N�F���&^
H����M*�ڀxxn��1F決�qR�Og ��v˻J����C�U����N�k
�=K�"�n���Xo/[*n$�ꛈ{qԄ�r�9�T���`#v[l\Yl���Lm��r\����쇤��ܶ�`�B�I+Nޛ�����hh��I햫��5�1�$p�mRW����*�յ*ҭPU�!���q�t<Z�vv��{۽[,�:r�U����Jo�)�@���S*�0�����^c�`;�t���B�*����X֍�l |K �.��R76l��\�r65h �&9fRKaƜ���v��GF�z�j���\<��!�;��]s�-�SP�m%V�$�݊^skHq[P���fUjR�*�aQ�q`��ѫ�m�\�d�;n�m � m%l���<08��NN�4]q[4:���v{*�<���X3�(�ї��^���qc��G�On6�y_d�͞Lm�\7k������V۶n��WV� 	l6��Mڍ\�ۥV�n��G�:�
֢�tf�ʬ���{�w��B�R>UA�+�H�'��#P$H'�\��!]�2�9���=v�fxԤ�f{F�i�e�^N�a�8��.:m��zr3ζ����ڻz����69y�tDOG<��\���mS��]6�%�{!�d�y�U�"�����B�s�bh�1Ű���N�&�6Wm��l�x2;l��=��OU#ɑ{m]+�W�~n�&�����+l��M;t`���m�2q�9���^�čռ�	��κ�u!d��v��Q�y�e:��vt')�g��2S^��w+l?绻��r�g��nD�N(ۊN���=�mz}�h������dbmFd�8���:}w��&f�7�� >ݭX���x�H��/�F��KZ��K���yN��]��{��e�LX<drAG&���w4
���*���؈��������;�Vի�QtU�P�Q�:�]��������u`�]f�{��q�c�lBq���� �������C[V��Y�P�F�aM��!�y�ۓ#qx˯�@/���WY�^}V�r߾�AG��	��w�o��| ������Z��k�|���}��
�W����>b���d�drh���h�U�U�W��f��:[�YIH�+����=335�=�W_��_m�{��=]΢&8�@r7�W�� ��4�l�/>�@�c`1�Y��SO E	�'��Z5�N�f����Mܨ���֩{&�Z4+J�^ ?�X �m`��[311��oo �5�5\)��!+�����f�y�Z]���٠u�ҩE��Brh�U�Uz�'��*���!o6�ygs|���{�U���Y]R8��^%��� ���x��, o�`��X���̀�E�p��.�+��u`�";37��p��-����U�I�7&4��dGX�b6�ڬJ�x6.У{Db�P{��wL�Z�ye(��w	
b���܌���
�W��f�箎��L�Nm��*�@��z}�h���{�FF7�4��8�
�W���3[�r0����ݻ�Y������l�-빠U�^��H>$w.�ė�7^+`�A]V�	%�7ב�lLDLm���Z����@��Щɑ�1�n&�Yt�͛�˹��QXŸ���w\�p�5�Hs���ɱ�)�ɚ]k�*�^�^�h���/�����H��#�$zW���� �^F ��lL�EQ����̀/]�TE]�| ��� o�#������>__����WX�&�y!2�M޻�VנUz� �٠y룸F(ɑ7s4
��@�g���׷��Հ7ב�D�G��QWE�ь�a�z��9�2�8���s�\% ���um���"WC��gK,�D���u����X���3��aЯ9;7i�V����yC����1��9ָ�]�3�F�Z�N���&�`�l+����9K��3�7;aD�:�e�Y��N�7$�L����W�{$7cO ��g=;6����πc���z��6V6����N�.?��.��c�Sb2�dMAjb��f�(�V����3�e헭948օ��L��Z#!��Ƚ�~��������ՠ]h�RD#�H���zj�{���� ���X����I���$��w4]�@��� �٠y�IT�"6�������`��x �kk{���7�nR�W$�	�X��@�ޯ@-�h޻��ՠ�z��?��׬���E1/KOe.u��`�7�4�юj�H�2<)����f7�ci�������h�f�k�hu�@�ꮱLMő�1�M }mb��L�K��LfW�V�����f�޺;���D�r'$�*������� �l�{�J4��T��Ҽ����x�����`��@.�h�RD�H��m����W ����}�xc��Uj��
s
��+@��n�;�	�.3�vv:�2c�ǂ1���I�q�G&�_y���`��G(׫=Twc���1��)1�3@��>4
���޳@����<�]QH�d���`�9Ws���*��{�ZA_@�X�JFe$i��Qٙ112�b{1�7��F;�`?�mr��J�+�T��+�~��{�X��F �h{���U�)��,���G&�}�s@�ڴ
�נ�4/]صM+6�nU�9�����<���:r��K@;Q��m�������ج�CM�Q�7ov�]n��� ��F }�֔�9?7"�*�^�[l�/[��Z�ZjT�4�0i�$�������f*�ov��ݼ��X+��UH��K�D��V��#��}�r��{�r�,�4�0��	PD�,�|E �O��>��K��ߝ�*`�9*��Z�ZVנ�4m��>��ߜ���Y������s �[m��=�nY���T�v�ŝd�4�ԛo�ܯz��uV���U��{׀������� ��𨤭+]���_ 7wV�m���ՠUmz/Uu�bnp�X�i`���7m�����{z��}4�KLI�!��ۙ�Z�ZW��m��w4��҃Cq(�F�4
�W������U���U���Ȭ���u��le�/�>Gyk���y^wU�<'��uw-�r9\��Ncu������Fq�0g���AE�\l_�������wa�z9�IsN3�;i5Rv�J�c�ۉt*�!�2v��9�# (;J��*vi�\f$ڻ`�[�3t#sWmm���^��B��I\$�]ͷ[�,���u{e����7�j�kk�J[Q� 
A��z{̃��*�Z%�踈j�����=μ�5���.�����Lrgk<,��Ē� crG�����z��)�Umz�K���F�m��I, }mg�7ui�mk���Y�}ߝ_G�$m�4��|hwW��4��h���I Мi������Հ�1[��`���¨J���i*����� �[׫�n�� u�]�
>�}��`�$W*2fv"�������&\���V��M�� ��.ë�Zk��z̀wt�@��(��4=|X
��%Q�1%��VB �� L��u�x�ְ�^FlMPu���4'�X�rC@�u������s@��h��b��R`nF��m����m��*���=�]L�P�*UwI`bcwsN���@-�h/Nh��I�H�����F�Qy�\u`ܳ����Jp3�eSq9:zI6��I)3@��hwW��4�l�-�)�(5�cBr��� 6���k n۬ى�5���fRT�Z�J�+���, }�\�x"o�`FL�b��bɁc9R@IPx�x�*�CHkdi����0��D?1��FXHZ�����Br)0��	�c�&SH�@�2 Q���`�&e8�`����!DC�&AN-�	THK$2Y��b�@C!��_��!��{��C~b�x?�1j"4����s��~80�B%�Ldt���z����;@�� B x ����#��R&#݈�����^��r��������)E]��Z��
��ڭoV�{��:���m��ڬ1'26�R%$�+�� ��N�wo��� }�����Zxz�.�l;<�g��!�m��$�vӨF]%܆y�>��p3�L:5�2ѠU�@-�h޻��ՠ^�*�LH��jG��4�]��n�_u�zf"=1v{Ѫ��(V��m4�G&��~���-v��z� �٠_>V<�hlM��s4]�@u�]������`��$�I#�蜘�^\�u�RV�BH.�E$� u�]�113[���o^�`�u�;n�2�N��.���T\R�m� w�%��5�(1G�;:������d)����� �k n۬��w�v+�V
bn$�S�rh޻���33>����>]~zm����}LI̍��s4�|�
���z��n���Q4��AH܋@��� ��`��`o�&o���`~��J�P)�R5#�z��n�m��.{�uʸ
1 �s/��_V�f���`9փ�j�)�(^�m�֔5�n(es���4 m�g��뜜��v��g�J����4��Bt\�l�n�/&���!ō�;��mv�������Yrk��.ݲv�n�m�bm3�fe4��i6z�����;�j�8�c���dӑ:�!��mG$�6"NN���2����u:�c8�v�`֬������%����7NW!cD�����t$���S������䧇TpDQ�mil�c/'S�����;s�ɎF�x���/�ۚ�S@��� �٠_>V<���ƚ��&h��؈��i�� ��X�����E"p�2<��$�hwW����&&b�{���n����WbJ�Z��I*�W�׫ }o# m���3Z���9�}17%�&&G&�o]�޻�Vנ��{eQdSY��.�s���Ԝn�����e��*��_;M�SQ[L-��n�m�����h^�@-�h���{�M&Ӕ��Q�-~�� �:@�H< �@M� ��*x8�_�����}��m��=�
H�,����q����n�m��]k�-Ή�L��H�m�M��s@��h{��������ү���B�<���p�Z`���� n��ב�|7�L0u���,��eYY�}��o���2I�B�A�È�&�cf�ܬM�p�E�p��� m��?��0�������v�]�v��wu`��h۹�U�W��1!g�����,���V� ?�� �Lñ1���*"�D\L�\J���^ n���Z�r$�i���S@�ޯ@-�h���=Gu�(��`��C@�޷�mn�����i��Wû�8�(��Z�g\�n=�@��������B�e����T ꛎ���g�����@�n�z�hu�@��*�1������S@��^�[l�=�>UL��	�mG3@�e4
����@��s@�l�9��cpJ'!�U�@-�4��iJ)�lM�Tw�w�\������ٻUj���wj������ywV���x����[|�EڰEZ���WX�C�ҧ�! �=*���BFv��{&HF&�Ĳd��$���nh���WZ�޳@�{U�F�q$�i����)�Uֽ �٠^�s@��	����NI!�Uֽ ���/[��[Қ��,�b� GV� m`��`�����{��_�>S#	#���94��h�ەw=���W{��!��(��2��9�
���pm�rr���;\�V�gM�R_#�Ӻr���TX��Ѭ0ɝOj�����a��r��k�7Mt瞻�e��i�k��zc�t���e9�^���Q�0NpIf�sґ+�YZ~u���ҷN��XN�^m��7N�K�C�*�8�򽶭�v�d}�(Â�mWl�pe�"�מ�8yA�<�\��yݧr\��p�of�����?Ȩ� ���������L�5g�(q�A\Uq�i5�ƴm�M坸�:�n���[�kq�6|��\��� u޻��_�&y@owf��}g�I��51����hwW������i����j�I]�QV�%V��wu`��0�DDDDMV���@�[��;=t��M�bɓ#�@�۹�[e4
���m��ڬ�6��&��$�h�M����f�}�s@���$Q&9�2B)�=nE�֤ء뵄F�u�N� <���gk �d����D��(���Wuzz٠_[����Z`�HԭE%UAqiik�]���?��B�U�V�����z֘��� |��X�B�IM������hwW���{��HɃ��"�f�yڴ
������n�r��I�Ec�)"�*�@/[4��j�?�ϯ�����f�ɉ9�)�����j����Z5U��Z�[.@�Ț�k��ߡǲG&	�$NG@?���ɠ�f�yڴ
���=�],&4�X��`����@��Z]���f�箖an@�$f$�h��@���<��qO�}�9k�����W�w���Z�p�x�73i8�
�W����w4?�/���}��F�)I'�b�= �l��@�e4
���߿���8�^,�0�B,�X	�.�s.���|�W�)���/r��v�&��踬P����_��}v�����@����+\QshT����3�3ɉ���kw��ެ 6��j8G	"cp���*�@/u�}�""*����7����^m+Wi�J��W�����������~����al�T> ��qY���r����И�QbS"I&�}�s@��V�Wuz{��=�\C�ci���;Fīԓ���I��@�-[�� �lF��i0S���9��ڴ
���޵鈏D�a��d`w[~�"��j�1��Wuz^�z��������71H�ĘL�@�ޯ@�۹�__U�U�^���V��2&H�)Z�������0��z� u�W�w�IT��4�E$�/����b#S{���yެ�LLL�į�b"����TV��DU�EQ_�E�"*�����TW�E @��RA�@��@�@��P�U@DA��+�qTW�""���+�"�����+�"��������"*���DU��TW��EQ_�"����(+$�k0��@2J�0
 ?��d��-�           �     ( �<�I
Q

T(    P ���@��P BQH
TT HPP  PB��	p   Z�Q ((  (� ��s��g���s���{<���
�;���k�ǈw[���p ��K�d< �q.rp;��ި3=�\Y�9� ����������ס�Å�aU� � @�   �P��s�ڏ{�^  �  @z� y�p@ D @ l h� �(@    
z� � 0P)  @ @ l� D @ D   l )@    b� R  0 � f (�, A�%�o�\�^�}�y�� w�m��>� F���������R�}��}9 ��4�ɽ��Ϸ+��a\�(��H    �$��N�z��x���4��/p }x�#�{�}�9+ Mҕ�˓��i�IX�+��@�p��o���rj{n0j� (��Ɉ�oO&���< >�(UH  � ��1 hq�c{���s�W��*�Ɨ�= <�>�s�{���^�� ��{x�x  z�iV-J�x �=Ucn�!��:�`��w�9=!�NMN���� C�7��J� h �@�JT   D��RO�P � =��CH�4� aT�Д{T���!����"$�JR��P�x��������?�?����rv�����w�� U�g/��������dTW����� 
��@EOO��:I$� �Ab`�(a"����@���/��LFZ�Zqe�,Z�aR��XX�62!k�i�B�X�(�D������V!8hp-�l��P�e��K����+��r�ʰ��Bԑ
�
g$9mww �d4�,	ZP�F��VB���-�"ܦ4���"G�9�I�@�	��7���15'ÁbX��;�	Jc�ą���b5�NK�$���M9:L�d�rp�t�IH�0�%Ӈ!��4f�(K�C"���(D�:p������!s3�+����H��I79m�Ni�I	p�V�Ӓ��(B��yBG$�@��#SH�P�P�e!Rc,��&�#9���Ѿ�{��D�@�F���Ąy.GÈH��'�B��$J���"�A�@(, ��T��A`8����(��"�Q(@��F���X�+�����"Ĉaa$ P"0V�A ��*bA�bl(i��!B���B��U(�".!�D+���i$�*!�% ���f��*`;�bKIm�	9J�`BZ��hbdA��1"ŬV����H�[���E���%MT�BZ� !r���i
rB%��␑�qj�n\�-cL�LY�R�����8y��!���D�\׏��
�I	���O#S80d�	. "�X:� ��|�0Ȁj��b-��pt+"�0 �@���o9B�Ֆ��'"�"\5� T`T�A"���Q�6�4�S-+�,�?I!
Y�B�B0"�cD�VaT$��ՋK0�80����m
T�%���
BD*XR��,�@����BIYI�,«��S��Ƹ�8�J$|ILi��y���"�Wo-l����FSiH�!|�G����,o��$ҁ�d0#�F����!$�E�L)�k/��j����顙78����0�h�¤h4�stc���i䑩����/�d��SNk�)�F�	�0��|?B@����HD���*�@a�#H0 Ac���Bk�Y4*+8���x¸b�rX�,�!�HF��0$+ HB&Y�
`�B�d@�I$���20�`����P�"�Ł�i.$BF�M#"5Cj��I�XE$�d�e0��)F!3d!\@�V4#	 ����B�BB�$�1��V�,	 Xa�����
`��!�p%D�FY�!#S���'��x:B�< ����@HĤH/�O�a �_!$�K,F��4�L���Jc�8�!�%)���E�$Û��Ð%�x�B{.���SaL�VK�O$�IFY3�a������C���$��� X���K&�o	"э��\�p�N��S�|��E�y�����{�xs������ῧ	Ȱ�Fo�O��	�2Y �퍄R��bo��6@#�$ha$!?A[!�2X����y���`āRB'�
I�0!`��$��@�H1�Jc��$&�����+2�&
L6@�E���$
 �q�$�"��˼���V��y˸emyh�;jZԩ��T�B	Q"� P�b�r��LT�HF4I�6QbH��I!�[��ZE.I�Fb�LRA$c Y
Hq���!%&\�C�"��$0��l[�@�$ I(C		aR�Yc�2!124�1�bP�(X��*9
��D�
@���h�*H�!i����H� ICCKBP��FI� A��_�@(1H�⚄�@���z�鍸h��)�=��@�Ht^��$�����)�A��B@�
�:�(@�`<��y� x8���G4�
�)!e�B���� ��$$Sy�:[0ѐ��uĂŋD�5ȱPcOXS�}� @p�����3C �MX%q"�թ�B!��px�9V�k���&d���@�B4.cB	����BT�1����ᄷ4�u�p�%�$��c���ׄԄ
aL#LX�p1$&hJ0� C��ydM0�1%�1��&a��C�i�+�
��7H��4��m���33$��`�@�3��	��
���I;�<!�y��С,Q5�8���M�wwH��%���cFa��,�1fj��X�i��Tg�n��B�z�VB̻��eIsK+֢+��*���E*R�/r#Ol��ۂ��qR
v��Fe<+ҌY����7vz�D���A!�4���&�+����/I���Ɉ�M%�IT��j�JV��n�mTR�医�AT�Q�R��6U�<ۿ^8�Us5�Z��5w93m��J2���2"U!]?6�Ş�P)���<L�#�=4�x�����A5e8�Jݿ���:�0X��h�
���ۛ��`j�<dH0�w��hQ�X)�(U�Mr��'���u�*B�����X����ZC8ž�'�#
�nK%�B!f�$�������`X�Y32?�ar0��,�I��m)n�eٓ��h��<	�!��@��H@o�[W���h�xE� ���[�� jF�p:x��?_�J�i��!�E�� �#����hi�6p4�p#�)��.��,K�K�	�/�&� B���� ���%͡&�Na�"�����8��JA�<#��~0e�v.�Sg=�穓$���ّ�IÁ!�����h�⟤������6������TƁ��B��e2�1������g����'Đ�Y���B	!�R+^����%��p��H�W�ju"jƑb��tӕ!#3��H�8�!
�k�JI��.D���� �l�
��ƶB�?Oό,��فns�~=b_1�	����l7M��]��X�!�� X�$d�o�$H餅����4э15&���_���H4�a��ྟ�RSx�@��)ą-�$F�M*����9�!D�]˂��$��o�E
8Q"�XF!A*a��V404x����:���x�(�<o����\4��_��|cdp�x������J'���Ĕ�C�n�IM�����}�J��<�IxBS	 A ��M#\bÞ���L4��qWN����R5`��#WH9��3w�<H_��!]x�?$�	���A�?N���43���)�͜��H�Ã	�/��p!�Y�K�:T��	3y))��`@�����d:j�ZB儓 թɂ�W��B59*��ZD)Z�
�!@444㥳5��Y�\ׄ.Z6��������@�OXHBS$�R,����H����va�zs|�e0!.I�D����"q8H'�Z�k�9!�1�<s���48�F�J]	Ǉ�h�U|P�\_��=�	a���39��(����$	������U   m� �`@ $    ��   h        p8  c��� sl�Ŗm q�#��]5�m[6���Y%�
(�
�*��'b�mUR�0 +�A��a����� m�$�m���[d]��j�ڪ���N�j�r�L�+l���Sj���P�   h   � ����H�Y��n�$�V�m���R2O9E��%���-� �F�
.�s`  �� �a ��M�a�l����V��Xr���UYV�����	��c��j���-!ʹ�X6鴒]�m���j�W��\���-U�%��{eS��@j��pR�U����v�L��,�Ԭt!PU�D@[N8D^f����k��mh6mH�C`�u��U�_=�T�(m�O$����*���v8�����`�ƻn�͕��W������˛�2+t�T�n�⪨���j�Sj ��۵U-�� [@ on���ؐ -��$H崐	��m�k@N m���d�b@��ۛg��e��F�I`���m���M� I"���[u�v-�� m� 6� �  q' Z��'@��[v�� S�m�6/*��;lmmP
KT�[T�� m��m������ 6��� p    6���im	��$ -�� If�"��	���ݻ[d� � m��z@ 8 �6[e����!s��U�)��Pd�*�c7�[��s"�Z�+I��.L��YM���]�e$60�FV�[\dѳd�)BҶ6퀷�m�	 �P�,�$�mKm�t�5�   -�E<��٦v�)8*��������M���`    a��  H�  ��  ��6�ඛl���ky�[\%��nf�b�m m[H��� ��  $[iI mf�p�ͳI�  ��    	 m��@hm   &�$     ��lmt    m���m���H Բ�m�:�0p h$Zlڶ�i���:Ԁ [@    >�	 �     8Y��� 8�` �	     �� �  Hm���H r@  �hۖ�� 6���  յ���%�/]sd���  -� ��v�j� m�ڵ���JI��#*��K�*�8�l�5�ʾn�n�x�ɴ��烐�n�q\dm����x�=[@Y�:	��DE�,r�W6��vF5���:5!V+��n��l���C��^��y�IFֻ��r�4���n�f�����LǶ�\i[�V^����rn`5v8.jv�mlm�d����N���it���-C���7�&	9���чv��ou��q��&`ى+��Q���� m���l�\���T1t�U*�J���-�2O1�,O��U	
8��ʺ���HRL�UA�f�J����WMU�UV�@���yNh�N�� p  ��X6����gR�/@N$h � "ڷ\� �@[E:�ۛi0@nݱml m�lͶ�5l� ���m��6�mm�   � � �m��q&�L$ HXIm�n ��`m�͵� kn-�&�� � �����I�����m��-�W;*�PGD�Q��K(P�
j8����`��h8�
� �(��;m7'\�����e�L�}m_J��@�U+�@��m�m�GU� �����[@H�9��;l� \�A�Zm��mP�$nX�	��88�m��q�N�Z����y햀f��P�%��Ӧ  <5�sV��T�� �v���:Ʋn��6�Cn�{+,��Ҷ	�5�Mlܣ[S�7�V�Aj���o���@7l角t��Amr�m l���k<���$%�6۶�m�[��   ��I"�D��k�]ڪUꀎ�b�W+ �:ح�:���Z��ee:Y`��%l�V�*�Y�� [x$ �M�t��b껎kM� �\��-� 8ڥ�������ӱ�( -���gA۰2	$����[����� m�4�i0 Ir� �ͤͬ�]�*Ę�m�  8�n���*�ٺ�eNRT&���6M���x��
�Y(Ac��o[H2��=$\Զ��I2�pm�kMUUR���4��	 �`�6�I�Seh�G6�S��t�Ԯ҃��<��ܫTR�Қޒ�;m�ղ�	 ��A"md����c� 
U�	V�����m�ݦ	-� Id��M� m�4݃ZŴ�U]0 *�+�]��Ut�����c �� �` ���HZl��i1���Lm����im�cm� 	-��ۭ` m�m����Kh� /Zu�k5�` ڛIp6� &��UlY��۲p8  ��������`�ѶĎn�mm�H  p   9�}�}��m�I�`    ��$Xn ��.���#��$6� 4P�UT8W���6�UCi�6�m@�[��  K(  Am&�k5Ė� � p$l�c9@ �a�E�ց  �M�  ��m�lm�i�i����[��Υ [BM�8qK�lG���UUl�T���m,��M����  �`  �I��@�����ض�  H�X[@�ƃHԫUR��UO.m��((�iUy��n�m��i\��[ǎ H�����L�Uu�*����WT�O[�����uP<B��AUU1�(56�ے��m�Y��vӲ��^u�mm;�%Ѩw*p�UR���c���u�A���zS$ m�~�m���[D�o8[:S�8�m�9�bB�Y��m͒Π�5U�k���		�� t�v�z��g    $[vېK;6۷�l-�
W6�=w[����UT������(����m m���J m���$ ���M��5M������ ��ם�u�n�j�T�����j��Wh��kZ��v�ҫ��;];H &Mk� mUv�ɕ�u_UJ�1����>w���!iKF�yE
���7i,��*.�M�6E�m�@0U��ݙFv�J�qRòb�+�V橳ŷe�������q\&��(6�5W[z� l�N9 	f�k  Am����ma�u�m&[@fN��ض� 4]�[A�S���[t�km��  6� k�&�k[m�&�a!oP�%�Ku� $dm3V��fD� �[N [�-�$ �u� [R��ͤ�I  m��nIV�W��ewf��=5M�MA�p�� U@V�F�Iф�n�kX~��-�p�����6݀�eY;l8�O���u��-��k%��8p ��Ԭ�T�I�(Z��nX[�`�I��I  $pm�F�[@I���́�6�m��� J���[]m����  m%��� �`kB�Y�@j� �E�4��X m���m��h��}mm� 8�� �  l	�����   6��X 2-�e%���( n��kz�6ػn`�Im�I���Y�D�k`�[�a� t��`�_��� ���a�m�e��� �h-����  �˻K��)v�a&�3���   �J�źE�[D�n����`sUH� � �^���[@�Ca"�ok��-�   !c[l�k�L� @*�s[�n0$ Z�e�(�d�� 	� �9�6\10$mT.�B�̖Y��a� -� ����pI�)Gm��PӀ  � �k�[`��^Ӣڐh    �;��.����6y�89������PaЪҼ�N����� ��EUTRJ�9�Ij��r�-$�KC�l� ��� )\�mA��gJ����@L�n��+`-�;v�kX [N�m��4�6�[[l��ݢ8
�6*����ʪ�`�mִ� �C`
Uګ������		�&�++UTJ�*��Z-   6�-�hm��n۰���HV�     6�� .ipp$  ��#F΋�T�R�J�  H�6� | �� imP��8����J�kj���m�-�8 � [@  m�$-�޵�k�඀6�n�-mUU�UrX˕U�V���j���@*���R� ^� m�-m�ln��ٷ37s2����@EJ�)�+?��pT<�e����x�T ��P?�!�> �Q
�AT�G���@u` � ��������"� j	��
�=tQx(��	�)�OUPx����~W�S����W ��%�x������ê>"u��P J�<b
���P:�#��� ����~ �C�@	�@2 ,`H��2"��b:������� \����CpG(��j$�`2 �Oߺ�P�P  �E`D��E�$LE��.�z���}X���: ��¾��/��t � x�� ��L �B�w�=@���c���AS��?�=���b��C�H�C
S��@z�E�x�N��<��5xI8FJ���D��$�a`A���� ���G�"	�(�������N"�E^���+��Erz���z�*~�*�����@`�"~�y����73c��mp�v$�r.�\Rl�l���܁i�IHK�6�X[m���z����U)Z��村�ں���b�Z!E�eV��a�fXӀ6�{u�����=��ٗ[Q�v[!;U�\� ]�S<����X�enX
��Mm�.7,<�`g���%�T��L��K;�X���&�8�x�I]sU�/Z���,�n�)j�p�Ը�9�v�cC])�ya��a���pGK�EPx�ո��x���m�n��1K����$�%#�(5ЁH#* grN5*�f�n��,�\#����d7	e1�h�lR��JQy"(�%P�l��U)x8�w"�T����V���s��^@3��յWV�d�n�ۀʀ�Ӓ_)5�ݥ�$��8p�;#[��a��[Pl�B�i��k�������1���L碷)�������ɲ\�^0����e2�N�vH�#.��G<ٗ���65�c; k��ٞ8ѧڰSö�Wo7J�7����Ӄ���O[u蓮�Cn�N"t���6�Y`��.Ԕ�<�hh
<�^@PC�a^�U��k-f�4:;]z����c/ 3J:�kk qV�*�*��@z��dL5^�[u��j�J
r�Y�n�m��g�̈́ڃG!���%�NW��c��`q!D��*�@9�����)�s/6��p�j���k(93�F7:�nx+ͻA���`�nv��2d����dkWi�B�P!-ɲ�B5�■%w(���89'\�$�v6J��z%�]�����n�A���17F^�\�%�U��UOF<s5#���� A�����1�r�;n�yC��C[�%�j�h�r��� �f��]W��Mp�+���v5!�Wlhr޸��m+ڙ�8�^1�Ͳ:�nW$�WZ$h�D�nWm�m�r��N�UYF:�Wl��CqJ:��ӇP�J�A��z9�R@�T���{��PC�A}� �̫A��2 G��?�/�TB�8~�����6l'��~�kr� ��5N�E�!���l��X4�ol���,m�M;YYG�E��nɓ�ƺ�է:�dZ�3��p[6�M������Pp<��ҧ[s�񷝲j��pBY�E��)�nRZ�����hm�ʍqѫv�t�U�xL<{��,'�|�i���֮5����n0V:�j�9uث��EBP��]�s�i�u����ۻ�������k�����}��
�

cۇdE{dT9��s��!���cf!�x��N~�s�,�Ҡ3ޭ��	��@v�|X�|FM��\�sfL���'}��s�U��7g,Ǖ�4��ҭ�UTb��1�9�n��Š^���ڴ�S@3��HD�Ȣpiȴ�q`{��,ޮ,<�I���uE����$��$�r'��Z�)�y�,Z�)�wX�$jb�&��Ƨ���GN�i�t�oX�D�I���b�7kdqd���'�z�hwK�z�h�j�=���&a!'2H����}����U:��qEz-�i�ߤ���`wN�X�\X�@̿���ԏ'$Z�)�{]�@�e4���U�ȤIbO"X'��Z�)�wW4�S@�Z�L��'pCr-���=��߿~^�h����v��Y]J6I��熃%Ľ��S=2.�U�9�<q�Vw�V�oMӑ���m��?���h�j�/YM ����i̊'&��w4k�h���y�\ٙ��?$w��,Rd�d�"s4'��{y$�{����&(�"��Y��!�B Aj,jI���4��0ެ��;��Xܢ��&Lr2<�Z�S@<�h۹�{]�@�ޯH��`��� ���^h	%��|�*�X��v����l�ڵ���ul�/2�5��-��n:a@���L��K���w��gu꽥H�A��}��nh�j�-���us@���2)Y�93@��V���x� �'y�$�Ɓ�]$U�N!8���h�M 󺹤����[n���ZגX��1��r
' �ޚ�;��X��M:I$kB��"�#�@�7���O;�e�ys"�ŉ��m���ڴl��y�\�=Gv'!1)G2Êڄ�r�6n��nL��F7t���??�b��{���h�)1�2c�9��~}��-����^z&f#�m�h7����̲<�Z�S@<�h۹�{]�@�޻2,a!'2H9�}c�-�s@��V�m��:���I��H�b�G�3�+m�4���-����ǠU�R"2700rf��@m�g�>V�^��[LDF��1g99�6.]��m��s�:R,+�	NA�9�n�7D�'0�XĨ�&�q�q͞[�m�X���Zn�خ#��3�8�q�����XV;ۭK^F��3�k�_}ʂ^t��R"��[��'��H�C��݌�;-��÷^]7� �p<n�6����k$��k��\MÞ��Â-��n�O8H�Ql��ؕ�[��̇���{���=}�j͛m�v�ڣH��Y�<k\<��n���ݜ��ў����"q
D8!�޻��<��=�n�~�ur� ��X��1��r���Ǡ^�s@��)�^���Z$"NdQ8�NG�^�s@��)�^����=�v�b�sɎD�h{e4�S@��ǡ31^���=��e@L�jL#N��V���e��-����ze\r�fdL�]q͵Ƙn�����j��gȻ]�[�9����ps��`n�,~������u����M���=�̮�r�����I;�{Ü�`)���qPO���=��o��O>ϻy�k�w���ȜB����ɚ[)�^��^�f�z���]EfU�yUxTxh9����@u��h���=���%��s�'!�L�W��h#�L�ɿ��x�rž�o�~����;k�5rNneس��뺽;.kpY	ͻUA�l����rh���=��/YM�k�@���%�Lq�&G���M��D�EP��h���r[�(��@H)�i�@�e4
���73�߿
�@:���w�E_DRI�m�e�~���=��H�B��P��#R^�f�z����M���=�5����q�7�z����M���/����y�W�Wg�\t�8���a��:��+��Kcjka^K��=~{������gC�:[�f������/YM��@�n�y��dN!8����h���}uנ^�s@�ޔ߳�$���2cq&�F���y���/[��y�Jh���y���I���͹sm�ss�|�� &}�}�`o}\X�\XZt�&���p�dTQ����rI���e��3sIsl��3@�ޔ�/YM�|��/[��x����/~q�&d��ૅ�;M�[#WU��+���9�[��#E<6�f.-�7���;�ν��������uٍcı'2HԆ�޾u�߿g��b""�i����h�#@]��/�O�D�H�z�w4=�M���<^��w��ʱ�29��{�\X�\X�&��M�ov+<�Q2&LN$���4�S@�{�z�4��F��"b`�`���.���nx܅�[�kF7]s�m���6q9ζ
�����b��d.;NNѺ�s��"�����l��lە�u�k-�Pd��^5�1�]��?u���rwb/U��ݫd�y�v�#lH.E�x�V�/m[��/m,M�uk4Fh�P�H���#y��B��Ⓩaf��Gzۀ
�։q���+�j���D�J��7=ۭ�:�U�(�Y%3�0�L�ٳn����Jt�t��`+�Ԧ�N)zԱ	��b��1��cQ&�F���U����/[��{�Jh���y�Q,H�q4�	4M���j�����;z��2=�M�k�Gg��,Rc�q�3@���3_W&^��{�Y
�/��@�e4�G�^�s@�ޔ�=�Ǎc
ı'2L�Hh/y�8�i�����,F���V�����	�z9�<:[��k�j��m�i�)��W{6#*�{�{']j���̰���h�Қ�)�w���*���a��L�<�)�32l��)�yϪ�/[��uk��&'�؜4�S@�_U��J�����h\�c�ɍě�dp�;��h���<�)�^���D�y"�ʺ����4�lh"&Z��4�^��<^�$1G�$�L#�9K��iE�˝6��V��+�V[\�ܤ2@r�$��Bq�3@�Қ�)�u�E�P^�s@��R�`��"���@�e4�)�^�s@�Қ��f4�#Ĝ�#R^���w4�'�U�U(@>"�J�`��J���NG%�$
@�����!J0��!�{��A.�O�0��IF-P��	] 9Z"V0��~'t��20#�F�$��_�:�O~ �_@<J�PH��ೄ�~Q_������4_����w��T|�}߷�� �}��2�;�͗u�]�h~����i�Ѡ&��"&fP4�~����"�O�h�uD^dTe����8y$��ߧ>e~���y<U�M=���L~���Dy�ڢ��F^L�!YKYU^n��(��;���jB3Ѕ��uٷE\~���s����߿׸7���/�m?������~�L�{�<h~���~�D_�̲���0�/��7�艉��<��?LDLDU{�<h<c���<�r�o~?�&�ٻ�r����9'�@��?{�h�"e���O����m=�G[eTVd]�QW�9���͏�6���*��3@�-�g�芘&#�1G<��T?� �{�o��O�;w��ģ�4�^�����/[��{�L�og��I��H&Ĥ2,Ӎ)u]/7"����*S3��w-p�{�i�� �$�I��:�V�z���Jh����p�&H����'��-�=U�c4�1����h~��m:�/2*2�  ���X�sCO�~�}���oc\DEP.�Qc�2*����@���~��Z9������X���Nno,�.�,�/�4����L����3C�%��s��'������$fL���%�9B�qػv�_k�kc�m��W�noZ��15vݭnC�n�r�;<E۴R�^�V�sx�X��FE�Ηה-�����9��u���w4Nز�O�Χ;g_&�'�+�8�	:-v�����euJ���N��7�؅	�yK��=<�[�}�Ar�
[��]���`�"�1�7f�.L6�#[��������{{���{��w��c��J-!�[:�t�OS����4M�r����;}���iy��F���)m8�R/C��3�f~_����3@����L�LO��3C�D���>��@]m�P���I8�"s7�����[>4����D��Mc4���;��UTU�UyYo��h���ץ4��hzS@�.4�)���5!�u�M���^��/YM��,����d )���^��/YM�Jh�4�O��$n8�h%��Wm����7O���x:,[1��bC:q�y!�F�˱��9v#�3����4�E��ȬȻʹ.��,F�At"�,W2w��ӒO�}�ץ4�r1��1A���u�F��-�DMRk�4��䊠�"��ӊ6�^�s@�Қ�)�u�M��h�)1�N"8�h��.X��b4�lh&&y�`���B�VЂ��C
Ku\3�G<v��lV�vTe�{�U��m�P6%��/0�O�r�F��-��b4�_cLb�I)	25!�u�M���^��/YM�n�K&(��s2���;{�X�\Y^m��j[X�y�f�M�e4W��2�LY�L��u���z�hzS@����}ʱ�Bb������Қ����>�x�}��{�4+:���̘�s�@��-�K=2.�U���v9��v,V�̏4c��b�7 �p�/�ՠym��/t���Қ���d�GN$��@�۹��٦��Қ�ڴs�h�)1�D8��L�/t���Қ�ڴ-����RX��x9���Қ�ڴ-��~����������>��x}�2�����wd�!�_]�@���o���M��M�{��$�&q���5��p�#�OfٽI���]G1ӕ.֛�uί-!��@����/t������}v���4��2b���Rf�{�4��4�h^����,eP��c��������}v�'�K��s@��hqQ��q�4܃#��}v��屠.�F���\��ԛ�����i�I)��빠^�M��M��Z����#6а�DA��Y8	��I�8���3{%�z�T m��v9��m!v���ck���[���9��!5��"0r�,�9d�:N5dS��/j�Vzk�c�H˅J�B��nW.SbV�\zL�-�s�l���i�x�7g�'.h�-s�$tv�m�&3N� p<�ejxM�:\�WjP۷n;-�]i��_}�d�[�Mө��TӫzrK��{�ꏧ:�XіBBr�1m9�nۛq˴nwU��g�h�k�����ϾD���oS��fY��8��}؍}iW�&X|���>���K�rb�#��;ޔ�/�ՠw��h�S@�N��ҐI'2HԆ�}v���s@�Қ��4z�Ȗ<D���d"�-�3��4����4<��U;V����Xʱ�1G?��{�4�S@��V���h���XLR%�x�ش���/MnT����ۧ8�gsų�N��tZ�#o��4�S@��V�����Jhq��9�D��dp�/�տ!��I�� �7�kRIT��������7���I(�e�Q�$N8�yJE�u�s@�Қ8��M�4k�w֑U�ve�<���;�)�u����4>���~��3@��>Ib�pQ��r[)�{zS@�n���M՝G��cU��!;C-�t�ܓ8nQ��-3Y�+�a��Z3�m����k_}����J߭���4��h��:�M޷r%�(̛���2��[�"b�\�O��Қ�����s�p�'�����{��g'�"	z�\��S@�e4]r�dP����x7�����@�����{e4��c��ƢM�28hޔ�:�M���[)���b��q��INv�Z�Z�e�<GkB�뺼[9.f{�\��5�����Ku2��F�p����@�l����hޔ�;�h�)1�D8��f|�S.&�M�4��h�#\���UQY�Yx�y��h	�f����OLϦ.߽�47�4��.��0����˺�4���n��3@^�����!��*H�$X�"��# �$�1  ���~-h�q!Ub��)���?����'��p�Lnd���a����|�#@s
&ba���[���/�ՠ^�0�F�B�5ٶ�^�WBOe���n���u����[sv�.����؅�Վa�9�$�<�gƁ�e4��^������`���z���ea�Y�w�p]�w,F�""&=1g��ՠ/{<h��&&*�!Q��.���0¯+@}mց�%����Q1v��M�w�w�uK$28�i�I)����\���X��|�C�虉�-��Z�?���I��!�<���/t���bg�'_�}mց�%��l\D�&&"E1��E�)'�E�5P��@@�#$Fb�X2@�Bd$Y�@bB@�AXA"A�D �,G@萑`|�@�"4H)#H�RaFH�{ ��	$d#�HA�,0R�!!E���!HH�BȐ	��������b ���H� E�@�đ�
�
�O��q*<�A��%,B-"�%�%hP�!s@�)�,6F~�Y��ƘE.�bK����͐�.��m�A�2��=�u�eHD(�h%ҕ�+H����� D�� 	��F(��,_H�L<'�<W�@ax�c��_����m��h��r�mI��[;<�8<�mbR�GZ�i �U�������n�!UR�����ykm��mY��]��&�k��U:К�z�m�YTga�k��c�y�sZ��j1���ͤtJ^��l��m�LqGV�����ۈ�3��溪�s'�+A�U�^y�x�mXq]�˫]�1nݔ.p)�-������a���u.��6�7l���F��pa'�%�����ҭJ����<7릇G���� �J���.�Q�T�ƨ���L���K��\�lP���"E����ێ7q�5ڭng��%X��d��tP��/3j���+ъ����{�����j��2m]�P]Ԫ��kW%2�DQ#���T�)�J���N����hW�n�Ctdg9Q�ņ�6�f8�aײ�8�genǵ][:��[l;a�Bs�`�G]�ҫ>`����e���e�6�N����2d��7M���\�#gݱ���ݸx���ێ�&�v�����/��(�=�o:�K֨�����[D�6]i��٢n%�m���j�;0᪍՘Zݥ�<���>j�*s5��$�HXm�z�*]��r[\@WT�����c�.�D��Z&�Z�����2�;_'����Il3ͭ�m'X���ۜ\�4e9.R��mA�u�l�8G��Uo`zv 9�E���V�^`9ͧ<��e����Q.[���'Wm�w8k�ǰ��m�2�n� 賟hR٤$V|L�/E����!�"8��ݷ'��^�V�s�Ug\��oD������J���nW���G	 UrY᪤S(sU�@�Kv۪�0P������\��ӧ����lU$t�N�df��vw]|��<|�Q��0�?}m�� ��\�j� �=�ש@��X���S�i�nh.�ݛ�����J���Z����5VT�c��^3�72�]��s� Ao��*�6�0����+���w��w�����&��G�8(�x��N@}AE<U��ŗ��3a	۝\$�'NIwN��i۹���s��]+�\lKq-�=v�fUmbM�V�7a!����.Z���G<��Ȳla��8�]`{G����8d��8��X�d��!y}�v�����軜�#�iSs��v;vt�Y��7b�F^�[U�����/<���M�mu�8(�ܫ��;a�-��v.�-*���y�y(����SvzSGO3�����T���<���V��c#r'5su�*�WGU�>[na�Db�����I�I��9��_���/�ՠw��8���@��hp��QuU�UU�fd^��I;�;���Qx����>���I?��f��U�&&����UE�fM^U����h���v#G3\�:�[u�[RD*�s�6����g�_[�;N��b4DR��F��8ued�p��9$��o$�#�TF!�g�7��w����U�,.�ȚmN9�حL�t��lЇU�r�Rݮ�U�c����Y�ǿ�ƢNH�'�w�|h�w4��h�U�w�uK$28����ff�I;�����
�=H��$O�����߫@�v#}��ߊX�������>����=��i�{�113v�ۭ��ƀ�V"�Ȭ̌�'#��;�U�{zS@�۹�����{���=���,i)�s$��Z��4-��{e4y�Z�t��l�V��X�ѳ��5R�f�c�9Q)�LUoj�a�D���a�Oɑ��G��[��^�M�}W����<A[�hjH�Y b�~i`���Jh���h�-�s3C���Y��fYyw�+N���Z(}�3��=����ң�1���(�Z�ڴ:���Jh{��Hzը��(�yJE�w> �g���hl��}v���T�s�����ԋ�\�ۗ8ٶ�+��b�(T1�x���I��!�9��}l��/YM>���1��w�_ �`�`�`��~�ӂ�A�A�A�A�ݷ�KI�]ݻ���n�>A�����ϧ 
X � � �������lll~��xpA�666?w��pA� %����Ϲ�Jd����ٹ�wg �`�`�`����ׂ�A�A�A�A��}��� ؂� � ������ � � � �߹����lll{߾��rB�&��wso �`�b�� �}������lll���ӂ�A�A�A�A��s��� � �(j' ~p^A���^>A�����m�'�ݐ���K�pA�666?w��pA�666($?����pA��������lll~��xpA�666?}$߳>�]6nI���qG*�̅�8zgZ������X�2�ٷC\W�}�9L�M�n���&f�>A�����ϧ �`�`�`����ׂ�A�A�A�A��}��� � � � ������ � � � ��}>�݆i�m������� � � � �������G�PH�dr6?�xpA�666?�}���� � � � �߹����lll{�߾�݆n�̸m���>A������� �`�`�`��{ϧ �`�`�`��~�ӂ�A�A�A�A������ � � � ����iwIrnL�3v�|�������>�|�������N>A����w� �`�b+`��~�Â�A�A�A�A�ӷ�KI�]ݻ���n�>A�����ϧ �`�`�b}������lll~��xpA�666?w��pA�666?ʊ��Tb&=�,��/�p��l�����^H'on���r��n�c�h�9W(`�rr���U��:t��mv[��q�%�S<�;������Au���72p���.�f��<��+OglL�ϡsmwkJ��[;S��<�^J帻nv��Y'N�tֺN���g����]h$�{h�"cR�F��\�q�]��˺$D��)4<���M����с��ո�������{��{��ܖm�:��v���C�l]WC���Ȯ���"%R\���ၺ������q�]�nnmۙwg� � � � ��o� �`�`�`��~�Â�A�A�A�A���Ӏ�� ?A �`�`����?� �`�`�`�~���L����ɻ������ � � � �߾����G�"����s�pA�666?�s�pA�666?{�}x �[{�l����sY2\�8 ���}8 ���>�|�������~�>A������� �`�`�`��>�>�6���ɛ�L͜|���`����O }mր�-���h6:"��Ⱥ�����@_,F��!��G�X����<��W�&6�C��d��L/d&�t��Cϥ���>�xs�u�����[�v�7&a�n����,O���§"X�%��}�gȖ%�bvw{0>�L�bX�����<�bX������.ٛ�4�Ȗ%�by���y�c�2%���~���bX�'��ϧȖ%�bw��*r'��L�bw��ϥ��.�ݶ��n�'�,K��}�LND�,K����'�,K��oxT�Kı;���yı,O��ϮNP�ZT�����{��7����vq<�bX�'{{§"X�%��}�gȖ%��̉���LND�,K��g�.d.l.e��v��'�,K��oxT�Kı;���yı,N��f'"X�%����gȖ%�w��m����-���S,��N%�{lq�v#Z�ZA��\�8�<c0�շ����S�,K����Kı;;����bX�'w��O"X�%����Ȗ%�bw;�;2mݲ����&f�'�,K����br"�ș��߹��yı,O��p�Ȗ%�bw�y���%�bX�{��f�4�&���76br%�bX���|8�D�,K���S�,p]��U!Ȝ��y��'�,K���{19ı,Om�l3\ݛ�pۙ��Ȗ%�bw��*r%�bX���;8�D�,K��ىȖ%�b~���yı,���K�Jf�ܷ7niS�,K���y���%�bX����ND�,K����'�,K��oxT�Kı�������t�j��ҳ5b�8�b�y�u�v+Z6\Rẞx�T.��l��q1��ݜO"X�%������Kı;����yı,N���ND�,K����'�,K����s-2ۻ-���ܻ��,K�����Kı;��9ı,N��;8�D�,K��ىȟeL�b_~��s!s�\˻��ݜO"X�%����9ı,N��;8�D�,K���S�,K�����Kı;콶��ݐ��2\�*r%�g��ȟw�}8�D�,K�߮�"X�%����gȖ%����]U�r'�_�9ı,O3�ٓi�Mܙ������%�bX����ND�,K�}�Ȗ%�bw��*r%�bX���;8�D�,�����v�~o���n��j9.��&b���C����[r�d��=w	������͘��nm�3sf'�,K��߹��yı,N���ND�,K����'�,K����br%�bX�����n��72��n�O"X�%����Ȗ%�bw�y���%�bX����ND�,K�}�ȟ
9S"X>��KK�Jn�ܷ7n�Ȗ%�bw߹��yı,s��ND��XdL����É�Kı=��ҧ"X�%����ge��.�ݶ��n�'�,K��=���Kı?w��q<�bX�'���Ȗ%�b{����yı,O���2�-��ۚn�Mͺ��bX�'���'�,K��۽�9ı,Ow��O"X�%��{۩Ȗ%�bATy���tø0�cI���,Q)�6�,�$d0�v-�ch��+֓�u	�u�;=Q��7T��MC�-���wh��8��^�\�f�\x��Cn�8��M���H:�JtG ���hO�lnu�xg
��ԙ�pq�z9H���i�9�@2��u����t��v�����ֵ�H�]��S������ۚ���[�ŞtS�܆D���7v�eݺ�o��/?�?����g(�%sl�3(���=��Ԅ�:�����ۙ��m��z��{�7��bX�v�eND�,K����'�,K��=���Kı;����yı,N��;m���4���K�T�Kı;���yı,N��f'��2%�b}���q<�bX�'�]�T�Kı;����6���ɛ�L͜O"X�%������Kı;����yı,N���ND�,K����'�,Kĳ���6�Y76����,K�����Kı;��9ı,N��;8�D�,K��ىȖ%�b{��{a����ˆ�w6q<�bX�'{{§"X�%��}�gȖ%�bvw{19ı,N��;8�D�,K�Q��n}�6]�fnm�vL�6���z�wl��2��;[�������[jf֗t���v�ݹ�O�,K����N'�,K����br%�bX���|8�D�,K���S�,K�����m��.�ٶf�n�'�,K����br�"dK�y�'�,K��n�T�Kı=��vq<�bX�'���}q�­ʥg����oq�~���yı,N���ND�,K���gȖ%�bvw{19ı,K�o���\�-˹����Ȗ%�bw�{*r%�bX���;8�D�,K��ىȖ%�b~���yı,O{/e�9m3H]�r�͕9ı,Ow��O"X�%������Kı?w��q<�bX�'{{§"X�%��������譙e�M{��S�jxBN�m�v#8z�+8ضv)�������9�	����Kı;;����bX�'���'�,K��oxP�Ug�2%�bw߹��yı,O���Xf�4�&����ىȖ%�b~���yı,N���ND�,K���gȖ%�bvw{19�2�D�;�߾��svne�nfn�O"X�%����9ı,Ow��O"X�0H����!"� b��� Ux p�'�V�~���zD�C�c��ԡ���$�&�`Db�!W�B�"@��������c��i1��bxĀ����k�&���N)�����w����3]Ux�@�M`�� H��DG �Q)�E � ��a؞��y��ND�,K���O"X�%��;�iwILܛ����*r%�bX���;8�D�,K��ىȖ%�bw�y���%�bX���
��bX�'���v�]��m�L�����%�bX����ND�,K����'�,K��oxT�Kı;���yı,Or��;�\��b��s3��!�&�na�m#�*N��S���딠�aV�R���{�K�����Kı;��9ı,N��;8�D�,K��ىȖ%�b_ݾ̹���[�sa�wgȖ%�bw��*r%�bX���vq<�bX�'gw��,K�����Kı=�����\�&n�%�*r%�bX���vq<�bX�'gw��,~!�2'��ϧȖ%�b}���ND�,K��N�&�6M�3e&f�'�,K����br%�bX���vq<�bX�'{{§"X��2'}���'�,K��_s���2ɹ�s76br%�bX���vq<�bX�'{{§"X�%��}�gȖ%�bvw{19ı,K�N�gp�홓K���b�jyJs/i�:,��Z��dB䣐l�ڧ5R���n���v�͜O"X�%����Ȗ%�bw�y���%�bX����ND�,K����'�,K�������]�sv�ʜ�bX�'}���O"X�%������Kı;����yı,N���ND�,K��o;m.�w6ɦn���yı,N��f'"X�%����gȖ%�bw��*r%�bX���vq<�bX�'���t�aV�R���{��7������}��}8�D�,K��*r%�bX���vq<�bX�'gw��,KĿ�}�s!s��.��v��'�,K��oxT�Kı;���yı,N��f'"X�%����gȖ%�bTQ�g�,Y(U�ΚYg�`8��)m����qY�h#kQ�)� *\1OI��������+�,ܑ�X�E���A
gB쪽y���M�웃��c���טή�v��i�w0��gWt�p�X�i�
dt�3V��F@��I���t�<�mr�pgn͠�v���4f;y�jD�ljx=ͧ�P���rm�պ`3���ɛ�n�6Q�:�n�ݝ�;�p��������j��l���kv�x^I	���Ί3��f�ݝ�pf�7d�v�sJf�]ҧbX�%��s���%�bX����ND�,K����'�,K��oxT�Kı;���2m3dݳ6Rfl�yı,N��f'"X�%����gȖ%�bw��*r%�bX���vq<�bX�'r�;a��,��w3sf'"X�%����gȖ%�bw��*r%�bX�w�vq<�bX�'gw��,K����{i�����7m����%�bX���
��bX�'����O"X�%������Kı=��;8�D�,K����\�nsr�ݹ�ND�,K����'�,K����br%�bX�����O"X�%����Ȗ%�by����Q�!uuS�.�NnA���}p��qA��+��TIe���ާVY����%�bX����ND�,K����Kı;��9ı,O;�;8�D�,K��y�n[.칙�ff]ىȖ%�b{��vq<��TG�+������O"X�}|�S�,K������%�bX����ND�,K��s�.2�r�l7noȖ%�bw��*r%�bX�w�vq<�bX�'gw��,K������Kı=���vkwHf�]ҧ"X�@ X�w��r	 ����A$O�~�S�I�;��9ı,K��v�6��nܻnK�8�D�,K��ىȖ%�b{�����%�bX���
��bX�'����O"X�%�Hv]$�Ik��i{8�k��S�����f_
@������V��srm1,�ND�,K����'�,K��oxT�Kı<���yı,N��f'"X�%��?^��u�۹�nۻ�O"X�%����Ȗ%�by�y���%�bX����ND�,K����'��{��7���/�8n&F����}�X�%��}�gȖ%�bvw{19ǁP$T*��({��ؙ��vq<�bX�'���Ȗ%�b{�m�m��.��4ɻ�8�D�,K��ىȖ%�b{��vq<�bX�'{{§"X�%��}�gȖ%�����Ϩ �aV�R���{��2X�����O"X�%����Ȗ%�by�y���%�bX����ND�,���߽�n��r�+��\����-�\5�"�ك�+v�����:nۅ�M��v�ٻwgȖ%�bw��*r%�bX�w�vq<�bX�'gw��,K������yı,O{�;%�5��ɻ��4�Ȗ%�by�y���%�bX����ND�,K����Kı;��9ı,N�};L�L�7n]�%͜O"X�%������Kı=��;8�D�,K���S�,K����Kı;���rm3L�nn�f��ND�,K����Kı;��9ı,O;�;8�D�,*���"vg����bX�'s���n��w3�w6q<�bX�'{{§"X�%��}�gȖ%�bvw{19ı,O{��'�,K��풻c��<�j���g���.u7n�g�m�A�U�3�ݸ�ub�F��dh�w�,K����Kı;;����bX�'���g埢dK����
��bX�'~���\��m�L�����Kı;;����bX�'���gȖ%�bw��*r%�bX�w�v}��oq������~}@�3�[�J���bX�'���gȖ%�bw��*r%�bX�w�vq<�bX�'gw��,KĿ��;��n2훷v��'�,K��oxT�Kı<���yı,N��f'"X�%���y���%�bX��}�/f�t�7v2�9ı,O;�;8�D�,K��ىȖ%�b{��vq<�bX�'{{§"X�%���DX�~����w�d����ӂ�f2�v��Ž��PU�XKi��@5��WnܗnՓF��÷3�x�[���rqf�Ƥ��6�n��!��	���8n��s�n|턎�yMdj�ӳ��.��u�{r�×�Zq֞�Ao']���>�S��j����H���X:�,pF�f�x�����Ş���h.��]f1m7u�,��?i�=r������ll��+Y"u!7r.^d.�f���Z��e�["����B�����&�6Mۗm�sgS�%�bvw�'"X�%����oȖ%�bw��*r%�bX��{��'�,K��^�lɴ�&sn�nl��Kı=��;8�C��DȖ'�_�T�Kı?}�}8�D�,K��ىȖ%�b~�׽��wv�f��l�yı,N���ND�,K����'�,K����br%�bX�����O"X�%��w{m.i�t��nn�ҧ"X�%��}�gȖ%�bvw{19ı,O{��'�,K��oxT�Kı=����sn�rn��'�,K����br%�bX�~�{x�D�,K���S�,K������yı,O�����q�v�:�)�kcj���jk��]D��2�ծ"yNk�p��t4#8U�s.���%�bX��߾�O"X�%����Ȗ%�b~��;8�D�,K��ىȖ%�b_�{��r��.ٻrfm�yı,N���NC�D��6%��s���Kı;;����bX�'���gȖ%�bze�L����f�mff�9ı,O;�;8�D�,K��ىȖ?2&D�����yı,O��p�Ȗ%�by���2m3d͹�i36q<�bX�'gw��,K�������Kı;��9ı,O=���O"X�%�g��6��a77s�ىȖ%�by�����%�bX���
��bX�'����'�,K����br%�bX�~��ɗs-��l�l�3�&'�&�b�K�\�^����:s�Y^����i^��}��oq��%����Ȗ%�bw�y���%�bX����ND�,K����'�,K��;���4ۺ\ݷ7niS�,K����Kı;;����bX�'��{x�D�,K���S�,K�����K�]ͳl��ݜO"X�%������Kı;����y�O�H����>��§"X�%�������%�bX���n۶���s34�̻��,K�������Kı;��9ı,O=���O"X��ȟO����Kı/N��e�aq��ݹ36�<�bX�'{{§"X�%����Kı;;����bX�'�ｼO"X�%��$��3�M����2�Oe4�i��	����(p���)gO%�V��%�M���-ǻ��7��,O=���O"X�%������Kı;����yı,N���ND�,K����ͦl��3m&f�'�,K����br%�bX���vq<�bX�'{{§"X�%��}�gȖ%�bY�{fM��M���7vbr%�bX���vq<�bX�'{{§"X�%��}�gȖ%�bvw{19ı,Os�����n���v�͜O"X�%����Ȗ%�bw�y���%�bX����ND�, ���=z���ؙ��Kİ{�������sJ��bX�'}���O"X�%����}Ϧ'�,K��߹��yı,N���ND�,K�}�˿-�*%`���������m��V�l�C�T;q���V�%�qQ �S��Kı;;����bX�'w��O"X�%������"dK����Ӊ�Kı=��n۶���s34�̻��,K�����>9"X�}~�S�,K����Ӊ�Kı;;����bX�%���ܷ,�v�ۻwgȖ%�bw��*r%�bX���vq<�c�2&D�}�LND�,K�w�^'�,K��%�K{5���n]��ҧ"X�2'��ϧȖ%�b}>ߦ'"X�%���oȖ%��L����
��bX�%��O��i�&m��I����Kı;;����bX�'�ｼO"X�%����Ȗ%�by���yı,J,CF*�"H�p=�b�B$E�  �`�"�"&�tX� #<	TH�d@��TD�H�H*UCT�8@*�	�P�GT5�/8�W�� ��7؇�@�^CH:p�� ���j�(1�S������{ xЁ�?%���<8�`ĀA)� ë�"�$�S�= ���}����l��m �����9Uzn�Th8�edJ�61-I1�E j�^GUӆ�oKF�SE��Y�9��t���h]˱�,q�ȸ�xv���	f{r��������P�N��W�N�լ;�����j�n�NWh۲�WR
َk���y` 
�EР-N�ۭthø6zۦ��hB`7���n��J*KT�bݕثv,9�X�&��`ֱ�+j�SIUm.ݶ̭@H��Tt��չ��N� ���̺%��d��������	vXr�+r�O �kpIv��R���NIַ@]�^W���Lu����ɮ0b䈑�V�r�筦x]q��y�lcf��Wm�j���M���T�����s���H!��:�g�rn<���]��@�Ӹ]l�/<�:���Cgm��ۚ�T7n��{i�nks1�7[ ��Q���ΝĝK�]�t����N�6"��7;'U�]�(��5��DH픨���rt�)l��ǣ��� *���#cs¾T���j�]���\S��#�����*멸��S+[�r���vh�e��l���n��Wu	]n�y\�4Ѳ�WT�Z�Pe�jyvs͛�ê'SK��gj��z
z#	�V	7[ɶ�n�Ț�wls�<�!��.��X��l	ԂT�y6]1��*�c(�v�p�Xb��cl�5�#8�����R��â1;`�u,t"���8�խ�t\a7\) S��Xڞ�t��N�e0Lq�qU�&t�l�R�aV����u�`�m��{a$��x�8��c�)m`
^��V��:;5�.�yv�+"8��@�V@�ʯ/F�+N�%m[e��WG��utr�vmv��=�]k�Tu�j;i��r�U$��55\d�%����]�䗪5�64��yP%���ٱ����UU&a��˰�̧m����@hu�۴I9yRɖۖK�v�, 0J���PS��"�����<�L�3e���̜�fs֍��8"�m�F^����3ŕ���c^�讽��z��kQ�B�Z��N��s�6�;�(�M�j3�泋{K�DXM֒�9#GKN�+�wjm��ع��vً!�,r�EW[��vSdjW����Nώ8<=�7\�<��6e���9��':��I:���`�r�Fۢ�%�[p��ٍ���ݶ-��`�[lN��ٮ.�����]��v��κBp�4	+S�/6w�3�nݢ���n3�b����{��}|gGQ0����n���%�bX�����<�bX�'{{§"X�%������2%�b}>ߦ'"X�%�����M�7f�\6۹���Kı;��9ı,N��;8�D�,K��ىȖ%�bw�y���'�"�L�`��[K�wK��&�f�9ı,O��}8�D�,K��ىȖ%�bw�y���%�bX���
��bX�'���v�]���r�����%�gʂ@ȟO����Kı>��}8�D�,K���S�,K����ϧ�����ow�����g
�*���bX�'w��O"X�%����Ȗ%�bw�y���%�bX����{��7���{��~��. �y�rҩ,��ճḽ�����Ւ����Kn����W9��r�ˬ��v���Kı>��§"X�%��}�gȖ%�bvw{19ı,N��;8�D�,K�=�e��fi�����ҧ"X�%��}�g�(�*T9��0_�X�ؖ'���&'"X�%�����q<�bX�'{{§""eL�b}�w�fM�왹��I����Kı>�o��,K�����K�HdL����9ı,O��}8�D�,K�{�2m7d�nn����,K�����Kı;��9ı,N��;8�D�,��>�s�Ȗ%�bw=���u�ٹ���l�yı,N���ND�,K��{�Ӊ�%�bX�O��Ȗ%�bw�y���%�bX>�w/�t�ʩc�2U�c!k�2v��;��{-�'{\70պ�J[�\���w�,K����Kı;;����bX�'w���?��6%�b_�9ı,O��ן���wvᙻwgȖ%�bvw{19�9"X�{�>�O"X�%����9ı,N��;8�D�ʙ��ﹻnۗ4˗7ffeݘ��bX�'��ϧȖ%�bw��*r%�D?�T �τ�r'"o{ϧȖ%�`����r%�bX��}��[�n]e�v�����%�g�+"{��§"X�%��{ϧȖ%�`����r%�bX���vq<�bX�'rw	ov͙�f]�e�*r%�bX���vq<�bX�'gw��,K�����Kı;��4���������2��Ўi�&DpO���u=�N�w2l� ���Gn-��͂X6M�왹��I����Kİ}�{u9ı,N��;8�D�,K�oxT�Kı;���yı,O�}�ٓn�.��ff���Kı;����yı,Oݽ�S�,K����Kİ}�{u9쩑,K����t�7w32�m����%�bX��~�S�,K����K�F"}>ߦ'"X�%���s���%�bX?����t�ݙweܹ�ND�,K����'�,K��=���Kı;����yİ8/�T炋|����9ı,O�����wM̙��vq<�bX�'gw��,K�����Kı;��9ı,N��;8�D�,K�P;��}%�m�6ۻ]K6;l�8�$e���P��$�i4�ۘ����p�����V}߭�7���x�߹��yı,N���ND�,K����'�,K����br%�bX��}��[0�u���ݻ���Kı;��9�Dc�2%��{ϧȖ%�b}>ߦ'"X�%����gȖ%�b{��2�lٻ2ff�2�9ı,N��;8�D�,K��ىȖ%�bw�y���%�bX���
��bX�%�}�f�vL��ܤ����%�bX����ND�,K����'�,K��oxT�Kı;���y�q���~'��͊Nϻ��"X�'w��O"X�%����Ȗ%�bw�y���%�bX����ND�,K�Uz0��3&y��s]�J��nF����A�;Ex��iݶ�#ūt<m:�*��J�Q�����[\d����'G	ɖNV�ZDGF�۶�I����ַl�qR�����t�F1���W瓍a�u]��u�tG�TXz��k�M�l�c�ظA�٧9�dk���g�v�,�E���.�pZ���;�-�P�;#�W�%�y�q�4�������ڟ�:�Y�g�6.��)YY;O�u�h:����!��kZd�
�E�v���p�n��'�,K��oyS�,K����Kı;;����bX�'w��O"X�%����iwM�ٗ4��ͩȖ%�bw�y���*1ș��}�LND�,K�~�Ӊ�Kı;��T�Kı;�o;m.�wt�ə�wgȖ%�bvw{19ı,N��;8�D��ű;�؛����qI�<��ɒܲ�p�̹S`�'bw�y���%�bX���*r%�bX���vq<�bX�'gw��,Kľ{���f�Ypݻ�vq<�bX�'{{ʜ�bX�'}���O"X�%������Kı;����y=���ow��N?&m%(cV��J;s]�y_I�&�S�88[U�6۱�f(��\˻���9ı,N��;8�D�,K��ىȖ%�bw�y��� ��dK����*r%�bX����f�vL���I����Kİ}�{u9,K�����Kı?v��Li1D�L.�F�q>����{2�2��)"Mȴ��?�ηs@�Қ�)�wT�O�$#i�IG�3ɿѠ4������w֑U��Ye�V]^F�����i�? ���^�s@�zْH4'�&L���'4&�t��ۤ�Wжf�iۨ��"��:�D�)1I2'���4y�Z��hu��g��}l��=���H���ncm��e4��h�S@�e7�2f"=7a���*�(����3+2��ߖ�ݮ,�I+���)M��%�}�U����@������E��#�9�߲�Z������.Kc@�Ta��ywyu����z��5�ۚ���_��2'����m�j.q�8[h�̺u�ަĐrY��#�Y��I<�ȱ7�e4��h�S�������Y'���$����-����U,f���h��1�׽UP_��+.��˻��<�x�/YM��Z�w4펉bs�2�*�/0�q��h���%��� C�P���<���NI;߷�l���®��.��0�֕h�����igƁz�h{�(�1Hcq��M�1;���vȳ5�L�DX��tv�i�0�*�J!E?4�#�@�n�{�4�S��������_DH���q�i�`gmq`v�q`o�z,��W��i��M��^�E�Qy���Օxh~�}|�ODDMSM�h5����TY� �Ȥ�p�����K��>�}��y{�鉉��i�4�n�3&�3*��2��2��lh}1��|��Ɓ�_��� �y(��t��0�0ۓoV�/Es�l�Jgm��F�o2%m���땸J;D�۬Kh�`���i^�[U�v��7	/`Yvx�lZ�l��3�1�u�[��y�*���F+p��}n��1�Xmv�\qd��t۶�����<�3p�{f+7n�'>�ç�t�d���i�&�Ђ��s�TH���5��MYG��+M�DQF앹�v���}�L\�#�ӊ۲�u���av˘F��y�-��U��-��-ƭ8����n�8��h�#@ﯕz&'�M��K��o�,Nd�c�&I!�%]���M4���v�}�}_\�|f~%�T���iV�F��I����?��J�u�K��O<I*�jI%�[#J!E?�G�$���5$����x�U�Zԗ߳3����%����)"�Mō8�I%��$�vV�$�{:�<I+e�jI+B�l�A�B�m��G���.���ipq��XxD��(�:�fM?��yk�kE ��������b�"#}[љ�]p~4�k&b#�u�fBH]~HdR	<�H�7Ԓ]���4�F���~�~圶���~<�$������I{�|�I��6�D��y�I}��Q�$�������?6�w��$��~^x�]Ήa��Gdi�jI//m<�$����$���y�K�?f~̟��z�I%���$�9�8G12I<I%Ϭz�K��ߗ���}>�jI//m<�$��w�������u�B�<.+tC!
�WE��[����uӎ�V�:�cj�����6�&��bQ��I%��/<I/l��I%��$���=I$��\i@QO�p��y_�UU|�m阏DNfUw��������cԒ]���$��pI�$Qcm���r�o����ym��������8�Q�B)"�Y"`Ă �"0#�`F), `��2H�~S�@!W�����`j�`��[)
2�BD��$������am�l�1f.s.d��
�k�		�Ic�!	"c��߃X�d`�bD�]A�W�j����4��? �����h��,Ah�;����$��u�I[�"8��nD���/����~�RI^���%�Q�$����Ē�R�'�9nH�*�ﳕ~�UU蘟/~��}UU]�?~���������������d�\f�3�&'��t���9����0W�v>p���v�:��Cm�I)���}>�jI//m<�$�>��x�J��/<I%��'�&L�&�#q�K��O<�cm*���I+����$���5$����,Nd�A2I<I%Ϭz$�{:�<I/k��RIy{i�%�8ۙM�lJ8���/�@��E���ń��'���x��S�������Ɣ�I2���}V���M���/mz�g�Zh��w;;RSvu��4�a�ic��n��D�UjyT�'�������Ƣ9�t���~~g��Y�x���W�h��"8��n4��Uz���@��Z�������C"�$�'"��z�ԯ@��+��w,f��ӽ ��UQ�7�F�YI��������wY�z�W���^���~�LR%M&)��v#@�L�D�[N� �ӭ��d��� +ݓ,���74ܒ햄x#U���m���n�rєr��n�T��3��`.��W&�x����/0Vy4{]����QE���M�{F��v��gwc\�����Y�մ�֓z���Y\L�ts��&�ܛ=qlm�.�ݛUـ�s!��k6X��Γ�-�B�cF��J�c��2�MG��sζ�]m���R��93���m��X73��n^�{�ƴ�scV�qW!K��S�z
S�ٶۍZɲ��:��s�\�o��p�ͦê��*���������>k�&��JcR9&66�zz������Қ��{�� ���,����&C//+@U�ށ�v#OUu4�@]iցz�B$C��M�n=�Қ��zz����� ��"8��neYW���.W�?CZ�_ �{נ~]���[n�HF�2bɌ�"��d�V��k�y��dI��X����1b���A�����q���^��/Jh����ږI�䑶�D��h�����8i�4��$�ʭ�,��zz���z�`�&L�&��@�����^�bW��hw�=β��9�Ȅ�$���~\��=�-������~4��h
%1��y��w�ʴL̫���5��?R�zm�;����E]Z�(LW�t\3+ջ<���:�@���{-�C�9u�8�C�"���GZ/z��Қ��zz�����H�L�M�r=�Қ��zz����^�~H>��H��nD��z��=�}V���/z��Қ�Z��@y�bn=�^���rw�~]���E}m;����̛�#M��%"�9{��^��<W��;��h~��33���#X�L��4�]�Y�����w$���w���@��n������}n������D�{��#��LN>�����<W��;��h���9�%��nD'�$4����H���@���@�����3/��D�5#�ccnG�^w�u}����W�c4��z�������?<�QŠr���<�)�x�W������C�&
�����I�ﷶٚ�L�M�r=�Қ�~�_�����h���=eXۭ) &����v��]]����v�$ CV'8k��[�&�Y��k:R!5�18h+����^�߳?x����@�~�!�B!�NE����h���Ϫ�<W����A��x�I�ڀr���=^�j�y��j�<W��12c�m18�Ϫ�<W��/�ՠr���9qV�p�$��#�@�^�@��V���^�y�Z���D.a�6:�@�%���e�5nX�r;v��V����P��i�����sԘ�@Ғ��X�dӺxy�r-^h����L�0nt�N��`- <F#�����L�{�v����@eD�r�+�:%NgX�*���];W\#�����K�Jvnu�d.�<�k\��,���2�d�$S��t3nCi�oOnM�ٛ�n��c�v��)}O��s��a�W@P\�����Z�b���F;���H�\b#<�z�;�}��b䦮\�G@����9{k�/>�@�^�@<�\b&(��6B(��9{k�/>�@�^�@��V��1#��Ȅ�6����̽�N��r�=311O���*�z^ҬdR!5�����~�蘵�~�����:�J��ʴ��$2(D8'��z�ڴ^��Ϫ�=W��L���km������
])�i�eF���p.͞�{]O��/�{�?}�d��9���$���*�z��h����j�/eFbdd�i�K�_*��1""��z�@}mց��O@�,��C�$�h��h�j�9{k�/>�@�n�PS��Ȼ.�2�=3>����z�I��Ϫ�<���/W��F`G������^�虏D�y��|z߫@_ZU�[��5#�$�7�!�D�Y"ê�e�m͕ct�ᛮW'
�c���\"�6�Ƶnm�nG�^}V��}V�}v���^�W���N6��8�+�阪[u�*��@]|�@��*�̬*	�&���X��c��g�M4���#�8��Pz
.�8,zg��^�h��Z��UFd�^F]��RJE�r���/>�@�@��V�y{*0�H8���@����������_�~�h_%z�����E�U��x�:J�kY+ ��K\���JD&3f�i�k����-�3�,�&�I�~o��t��ZW�[����Zu�&ޅV
cR9&<lr-��Z�����9ڷ��A���Y1E?y��@�iր��V�������Z�n���	H�L�m��-��9�y$���o$�A� 0^ ���~�Z����!�N6��8�9ڴ�h��Ϫ�/�_�i.����IMˡ�g�X
o�^ ���A��mt:��Fl$r1�����~�_*�ZT�fg��ۭ �TfK�26�D��h���ՠy�ՠ^v���g�ă=��%����lmŠ}_�-�v��h��9ڒ��rd�&H���������|hu�L���X�h	'�Ued]f\�69�yڴy�Z�j�<���I8k�ȐbHFB���S��A�`UEq��4G�QH!�!$B����)��$�K$�s���x25�*zH�T�%����#���%"P���!d� E|�h~ �J��y�����d H��p�s�V�]N�8�RK=,֧Jy�������J������z׉=�d�e��m9�ƌS�a��c�k7&̶^�4��I�:J6�ͬ��\�z�P��9x�	]�ݞ�K;rʛ+R�tgQ(9�M�Z�[����:;Z�V��v8hv��Zyje9:LE�6nq���n��ge�tv��ȵ�Ҷ��$�J����Ex�K&k5���A�������m�eh
N�nMv��1{!��m�� h��%ඦ�j���L�*�[WXrԬ���.��Y��=�����k$���x�V]��)�%Ki9.l�m�oI/Q (P�FTۖf6�*t��� ����l;Oms�9J@d �3*�ѭ���S�] %�㭶�q��q�n7u:ūv9-���;��8�]�=U�&�6Q�걪KYF��;n���p��w ��Bt�0�lR���K��b���&�l��gm;0mi�@����V��y�H���Zq��ҽQ.]��<\��`<�j֑p�9ɓDQ2�-m0�mv�ڗqt���tD�ŔM5l�j�<DK���%u:�U��tjب�ڍM@K�<�4� ���g)"�����NB6�['Ha�	�����j��T�����!���GH�� ���xw=wZ���b�n���T�;=L���]�dT.�okk��v�pF��zB=�˛v���h�d�Z�n��*���9�6���Li�3�Pl]��A��ͺ�=[��p�v�q�@1���nP	&3=:{0���ݶ���Yݺ��\�hvƤ%��Wf�����$ ���WYI��7euE+�m+;�F�R��vmP[�l���#�W�����vIcr�^��5���x`ث������������n�*�c7'S�����uļi _��]*�Nm�8r�UJ��<��%b���r��:�2��67���:8U�d��ٷs3�OC�(�p�E4x��@���Q�`
��]��C��頂j��Oŗ���g�ܐ��ܤͼh��Yk l��p&Q^M�X(Q�8�u7W	\�m�ʇ-ͻd��s4��vI�^ز�����瓧h���S����w]O\F�u�rx�:�Ș��3�9�p��C%�&�UKv�7)�������k�&��B���<	�n^��N��v�y�÷�u�A��LݻlE�-�O;�z�[�r��{��������^�:�EF�i�f%�B�mb'���͜��qr���#����h:�W�=h���	_*�ZU�~�J��LD~�i�Ɓ��}�5" ���q�$Z�j�?u�Z��>��Z�""j��a�	���)��|��S@��U�^}V�WR�ȡ��kqhg艧�Y�r��@]|�C�15���@�ߒ͟�&D�ȱ(�{Ϫ�?���_��{_�-�}V��>���n	�p ����ڍ�[��kr�5�A�U��5vȅ�L�{����?w��\Z�W+�����u�~�J���z"#�+N���UQ3L�4��f���I<�;��߾E��%��1�<y��?+N��ʷ�T$��LS��1�c�hw��@��U�^}V��;V�y�D�b$�����;�`f��X��4�Q���t�����?6�)"�<��hu�Z��W�}�ʴLO�{wuL235`l�M��#�9cj��36N�{/R��F:+��n��_��v�o����+ga��۝�ՠ~��z�|��?�>V�h�>I�B!�8�6��=��Z����]�@����H=��O͓"i�ASS`oO}�w�ĩ��Fl�E���W����LP��66��<��hs�hs�>�ˬ�-�w�d�&G19$�@�@�U�{Ϫ�<��h�dn�M&∑�Ha���v�=b���3�����ɉ�qF�ӫ��5���dC$�69�{]�h��9�Z��Z��� ����2'�����k�zS@��H�9��cn=��h��i�����>4
���2,�	�ƜZ�w���������XsK�i����@�u*L�	Ʊ��oJh��_U�y�ՠy�\�dMD9&���f|B�bx��G=F��}\v-w����<�����d���D�Ȕn�ߖ�k�9ڴzS@<��I�8˺�����U�����mր��hs�U�,�&LR`�#�@�@ﯕh�"b���Z�ӭ���A2b��1�c�h��^��+�h��h��\�&B~j'���W�8�����u�v�h�ʴ�0@"  w�t����vKv������1:�-�XCr��U�=5on�{6ɵ�
ua�fl���vM��L�`äy�̬q4�x��䭕L鎋F�oF[O��uKͮs�Ξ�m��Fn�c����7/n��ӵ�]��ܬ�I���r�Zv�:M0�.�q	�u���F�6Up�6wm%<A�ӈ�=a�g��\=�?�s��ﳚ�;g]f���wulf�;,D�6��n�X�g-��G975�1U��]�t�ssP05" ���q�������=���;�U�r�נx��"�0��&
E�{_U�w>�@��@�V���T�H	Ʊ������v���Z��� ��FI�ȔM<�%"�<�j�<�ՠ{Ϫ�-�����LP��&��z�ՠ~����K��]�h����;O$q�e^��lWb�Wlí��,�s�k�����.z�F��̒d�&�H�k�l����^�k�hm�<��rL�2f�䓽��s�|E������Ǡy��}V��=�ȖL�$8�N-�����Z��Z�S@���$C�ێ1��k�h��h�M����x(ȲL$c���h��h�M����j�Ah��̂ڟ�k�Q�K��*��/3Ƨ��[�@'E�%�u:GV͇��Z�S@��@�ڴk�޵'�"Q4�%����^�k�h��h�M ��Ta&(F�"bH���{���N�Yk��n�bBI�5�5�%K3���>���3��s$��9#�@���@��h����V�o@(L���,x��Z�S@��@�ڴk�Y������\mh�RsEu�+նy`ܵ��<�4v��w�"[y���݇7+}�����j�=���-��[v�s�n8��z�վ��>W� ��Ɓ��S�33?$U�eI�c�I���H���h�M����j�:��*�ʌ����"���LǢf��~���}{����w���I�?��TP����C��9�����5����b��@��@��Z��Zz������ح�� 6��#��Nm�,����ǒ�NR�.�c��g[�M	�������S�������$��7�b������@���@�_U��U�|�
���@�bd�Š{_U�[Қ/mz���DD�EP�zFEf^fE��y��7gƁ��^�k�k���Ɏ%�c���4^��]�@���A��D�6��m�fQe���^Yv��-v�����)�r�נ������O��0n�hb|]�Rm�x�T�Z�nݬ񍪺�w6Z�y�z��YYv4��8�h�. ;U���N�1�؋�:��ZH�;LlkDlV+�r�m��Ѯ��یt�ݵ<�,�\�U�-�͉I����v��;�<q�/Q'hL����"ͻi?��� �����'0���c�Y8�ݰ�����PB%�{���Xܬ�7"�l�gN�����Ĥ�͇f��;���u=����-�3��s6�^[��P(�E��	1��)�w������:�J�31���n��m�F`H�CN-���9{k�/;V��}V��Z���ȔM<��/mz�J��D�bbbf�z߫@��x�ˢ�	1B7�b����@���@��Zz�Z+D�;�HLX�V��U�z&=1~���/z��ՠUܐ�������)�7��&*��i��W����4Ș�ѣ�Ck�]dklm[�1�c�h���޻V�yڴk�U�#K&8�㘢R/m{��%8 �,��( '���"�����גO�g~��w��hm�"D1����q���@�_*��1M<f����R�UeE�fE�]�fV���LL�E�k�h~�/mz�j�;ҕk�$	�HiŠ^��/mz�j�=����������v��.�,�N�'�-��N��v\1�-��n����������J9$�<���^v�������/eFb��!4�#�/;V��U�.X���\��U
�*����@�b�$qh�-����0�~̐�f4(�����B$b�1�,\}!��L���Fvܡced�!	�9@Љp��%P�+�A�6� �$c��Ax��Q��Y_ �����
*#��� ��:!��A�:Uq` � �C�9��;���}V�����nLx��E�^X���@]iV����x�hM;�,����sJC@��@��Z��Z�)�e��<rI$x��nH�;s7-<���) ��2se%��b��-v�ȑ"���q������h��h�#�?�sw�:i�eF`fE�l�@���@�e4^���ՠr�R���D8�6��/YM��^�bj���@�iր}�Q�y�YwWUWxhz��w�5mց�U��Dd�ߝrՠ��%��x��M�#�ZU�?D�/k�|��ՠu|������LVu��ڐ��i5�����z����V�.32��X��k��tHf歪㚜Z��Z�j�9{k�/;V��˂XI���1�c�h����~�ϒ��@�z����LLUM;�+�@7���@������@���@��Zs�b���q`ۏC�33*�o4v�h�*�:�J���Pș&79&��}V���33>�N�~�9$����I?*����b&�	�}���-s���e�۶�Yf�k3�qÐ��m���]�uq�Zx і���퀽�:�9�͔kqs������_�Oȭ`�\�I���v�]vw-q5�Ƨ�[Y�m�g�!�N1s�	[����j�.�&�m�9;[gI�m��x�m���et��гf���
��`*:�;s�wH[�r��km�r��ǜdu'n�igE��{���$��y�f�ni�&a���Gfs7�]���Fmg
t3�u+��mtZ- H���_������� �l�g�߼A�;��:��?I���bIŠr�נ����Z�j�=�%��x��M1H���@���O�3�_W��@�����Ԗ�s�4k��ՠr�נ��[.	a&
F�ǉ�E�z���>���}���o�M�����,{�"���=��M�A�rtV�I�\�V���jy�B=�%��8 ɀ��@��@<�f��}V���@�|�,C�܏i33s�I����
��hS~O�Y�}7�XG}���|��$	1���4k�Wuz&fj�sw�&�@�����ʌ�̢�.�+C�1]i;�sw��,�>���=�*͟��F�ȰIŠr�נ�������Z��&�j���6�Mw2T�0;r��z;)��W�k��m�.��������o�vm������$�h+�Z�үO�\��8��ȼ�̊2�3@�_*�133Ts��@U�ހw%���31v4�/�Ve�d]��Z��ՠu|��虉����_$�i$�ϲ�����,w]�P�@@70���>�߿b�����女�}V�yڴm�"D2C�^Qwyz�J�D�L����[u�r�נg�>@����#q�2A�,r<�1v��fڞntXu�1�Ae��H��1ōH��w�^��/mz�j�9z�J(��$C�cn-r�k�L�M��{נy߽Z��V�e#�>Y��Cy$�4
�y�Z:�v�h<f�G�/�Ȭ���/A�O�"f/�}�������?(AF �,b��P
)�3��ş�m�z�T�c��nJ�>WʴDĴ���U�ހ�ҭ����/��5��v���q
�Wj���I�nzD�nu�8�N��O���w}v]��r/ ���Z/mz�)�{_U�{z�b�	`70���^���ՠ{_U�^v���H�9��Cn=�h��i����fc�?��|����=�ؐȡ�2��@�_*�ZU�u|��zff���@\}�Z��0�5��Z�j�?�3?+���[u�|��hL?�����&*���$�e�)g�m˻vܒ��t1u����s�źj«kQQ��]s�H�Q<n��`��L	��m���=m��Iͺ��qXN�Z�:�[d�n�3�k��Jz���������3uv�z�;��*���/<ֲ�[�ܜ.�1@�r��J۞^��On.�����P�!Wm�F�������ώy�*+�m�vw�����W��ӚӶ[�3.��K.i��M�$A�+2B]�W5Kv��X,ψV��7O<A�լ�m�ÿ��[�����N�kGW�����/����/;V��}V�yڴ<�� ��Q�6�z�j���~�ؑ�;��>��>�@�GjK2I9�7"�<�j�/;V���^�yڴ}f	pR9&6`�"�/;V���W�.��A�LW<N�i�YQ��sQŠr�נ^v�����h ao⹃Ƣ�8��FLL��A�f��F��T9�5[P��Gy�ա�j3���Dn=�h��h�����<AW}��;���!�B#$d1'��}V�L�͖��@�ֽ�h�jZ�d�"j	8��ՠ{Ϫ�옚����>V�h�Ȍ��ʬ������4?�f&+�'ZV�h�ҭ1��oƀg��� p� �qh�V��;V�m��=��hv	\��)ḋV[����
;��2s�G�0��(�
������������h�m�u���-������Z� �Z(�$���Zs���Z[)�y�տ~�Ď���� 8 ndPrNI;}��䓽��rx
�	BI��i&�$�d��Ł��Ł��`��rG�@��h��h	,F��c�6�{נ?_��E�Xe�P��4k�l����^�m��ð�F�(@�S�#EN����y������Vq�ہ:��t��&��ٓpHiŠ[e4^��l���}V��qVl�$J6�E�������L�P��h�:�X� ��%UAxdsb���m��=���-��/mz��%���$�����쉊�ր��h_%z�����&fT�EDLc���}`P6V^�d^E�[e4^��l���}V��;���.��]uZAԍ�zt\3+ͳ� ���g�&�m�����i�m[+qb���@Ib4��3陉�����������D1��H�#q��M��W�[e4����ȡ̻�u�%����DDU:�ށ��O��-KTL��M�&��@��h{k�-����h��Y'� �i�I��mz�S@���I;��g$�}}R"D���Y �"��H��F$�X1�B �H'�����cW��"� �T�E`'H5f�T��G� ��(t�� ��%H�`�"�"��,
%+C�ٹ(F9�M$�	X���C�]ۻ���p�1��W�ɛ������`����"\*���JX��+~@�9DG���=���OOu�������~�[x�mUTu\;��v��� ���:�݊�e�2���8������&q��x���F��X��t��r`��L'���^+eA��*�[@�����m8��F����褧I��	�}� W����	g�����[UE��W7.�b\���/5mU\�6�YL��S*�m�ݵ�ݸ{F�뭪�ײD�$�b#����d jT��l����&1�hH���Œ���r ۵R�QV�k9,�튳6��z��d����Z՜��iV�]j���Q��B։M����K�����7Ж�}g��v9]A�5�<6��h�j�s�j���ں��37��]Q6����yܳKhU�ta�y�����O�s=��ʘ��`�F�;f+{���3�g]�6�z���^(�8z4�8��L�=sm �'
C���N��z[�q�MR��FX�[��y���tC��C��XGh�=�#��&�hs;^��Ɓ�n�w6��v�+�D�zwi��dm`
5H��d}�m�X�3mU[X�nڪ��8��#�ΐ^"f����+gE ��id�'O����6����m88��%7!�ٶ���H I�k����\�f��H䅆�dy#E-�v8��Ƃ][=�����ù�e��������sCNN�d1�k�O$A�0U���yՑ�4; 	C�;���������aN�%N�K�}Z�v��� V��U����.ն�	�W;�x��vj,�X��М�ɤ-��ե�ki0���#�^t/E<�1��vb(�JT]�1���{UVኘ�^��2��mJKN�v�qQ�&��ӷ,��Jɹ�*�Jd�k��+#T@,�n[u貶�Ś2�ƶ_Gt�e�.�ث����K�&�[�(�8���E�Si��Leh۱�R��.�˅�UU�-�!J�+UH@�*�H�qT9�9�C�9V�B�gt
�v�B4mɓz�4X��N���W���z��ŋ�QG���[��=3
hY��ۘJ��{&�6ٻ[��cY܉�.�]�v)�o8�.�n�dn�ڻ=h8{���<dD5<=�����(��kr�8:5��.&�Wk�D��\����!�Ͱg�ph�m�y���I0CX�S�(�	����vf�u�X��1����]��F�D�s��b�䦦��WeѦġ���"�ủ�ir�3�e��ƭC��m���j�����{����������c�%�⶞x����]����a����4�zl��B/������f���#��LR?������/>�@��h{k�=�v��s$�#�����[���������sw�$�鈙������l��32.�,���x���OESo�s��@�rܲ�0(32����@��+�X��|�C�334��h��U^y��e�^���h����x���@��U![R�K�i���{]Oac�z�����pզ��pJ�X3���K-������Z/mz��h�j\�risnf�f\��'{���/ >"a���"b"'߿^��,�|��o�$u��6~r
6�E�����[e4k�l��y� p��(�ʫ�̽11艉��{߼h��Zs�y��@�:Q,�$&������Z��Ǡyl��Wv<��v�P�6V��u�$0�/�ӝ3-ͤ�vI{.H��T$�G*��v���$��|���#�艈����-�}����	"�C@��X�l���}V�m��-�ZX�
j�MD�UT��\X�ދ3SV�i��1fg�+�M�}c�*��J��ˬ(.��s5�����>���m��9z�J(�Bq'��ZK����i�����>Wʴ������n�n�r�])�e����-���D���Hܗ2����E�ĭ��6��]�=�)�{_U�[e4�mI�G1F(��5�[e7�!�N��3@\�٠}�P^Ff`U�e�a�%|�@Ib4���4��h}���<����s�"�-X�r�u�$���3�:߳V�}�lb�	"�C@�eu�ze���v�h	,F��eZ����
ܐr�q�ܴ�j��qz���jݱŸ�k��j��c6�c���S@��Z�S@�ek@���2)X�P@�4_U�[e4�V�l���#�+�"Iı����h�+�=5M�f�ݧZ��Y��(�y&�4�V�l��k�l��y�,2I�1E//.��#@�x�~���,WZI� &���w綾쑇�RRL�̷-V�(��*㞶H����q�-��}C�U���az-X��5���J9������X^�dZ��[۝^�5�.i<9#,�Ҹ5�W�fy��y������e�ܡ���\nV"�Sf@�l�l�����P�lA���v���v��5��r�&�ٶ՜A�b !sr�'=��m�l[[���6�M�v�=��{�����w{��!f���\�,�k%8{r'W'k�*���4����qp�n ����n"9!@���|�l��z�ցm��<��5�7�4�Z�S}COր��h	_*�>\� � �(��4y��@��h��h�M�u���I�&����M����)�{Ϭz]�!�8��5�@���@��h���m��<��q�ZI�1̊y,���n.&��`�sP�
A�ݧtaz\���"d��N%����S@��X��S@���@=�*�?7�F�p�=��S$�oI|�j����,���`^��綤�p�"#I�#�/YM������=��=��(�dRbn"9!�{_U�^����Ǡ^����.X�#��ӑh�#@s<�<��4���V��u��]*˅��`������jv+�ˬɲ+U��in���6愍��$i,�!���b�/YM������-�F��1�1�Ԓ=���=���/YM�}c�*�R�,q� &h�=ӽoWC_4��Cd*R������f>�����c��v#@���+����cn-���=��=���=���m�Y'��#�&�{�,Z�)�{_U�^�����*�hC[.wf�C-�v���GMa��1N6��Z\#���Kr4�M��z�h��h����t�h�%�����r)������=�-���<�x �cP�cxcNE�^����Ǡ^����Z�۳@�IQ��3?b�/��_�Ɓ��５�+���M,���E���]���c��$z�e4U�r�hu����LCc����,d���dJ�r�'�j��u���R��a�:(d������]�h����>�������h�L��N%���y�Z��Ǡy�S@���~���O���N4����ߣ�/YM����}V�yz�`�B&�I�#�<�)�{_U�{Ϫ�=��=�J%��Ț�r)����}V��>��u��.1GU���a=,�v]�,��+{����c0%�W�3�l��`0i#�{WЭ��@أa��cv�箛0����s̻BۑQ�]���f�	�u����5ō�:뱞���u�5҈飵��� s+Aj�q�;���9�ݶ�`�����6�ε�=�9���sĥ{Po`�"��26ݻ*�@���	�,��?�3�[��$�mh�Ϟ���\C�T
'�&��燗���n[�i�m��kJW1-�v���d�]��"v]Z3�8��M4�]��#P�cxcNE@���Z��Ǡy�S���-��a�	"�Š{Ϭz�e4k�y�Z��~X�?9&8��G�y�S@���@��U�{Ϭz��HdN!c�<�����Z�|����/o��^k�ȱ�Iı���>�@��X�:�h��h=��
B�՛q�@�[�V)����WTyz��s�}�o����9˺y���#Y(���p����P=~��7fܹ�37s�O=��s�P1T	I�I&������t����N�X�ާ���[>�L�LM�9���;��=��h����YM�	��s6��@��U�{Ϭz�e4k�}�fE�#E#�Š{Ϯ^�������iց�_*����C���m5%ղpu �3]�ޣL�=P猍;�8�Q×Vl�|׊���~�~���4k�y�Z��Ǡx�T�E"K$�`�@���@��U�{Ϭz�e7�߿$^k��2,��Xۋ@��,l�T��b���&6�'�4|FF�$�$dE�
� B�,�!@��"!$`PH4�4BD�D���P"FF QF������F��	 �I �! �Ą�(Ĥ��B�X�Ă@�
@�A��*B� � /?��b� HD�#�AdY"��@��RBB02H"B@�B$$�I�"�Y HA�<� �c8��4V$#!	 �O�x`0H�X�a0�Q������H�[)+��.)�q:*C�����K���)`@���-��+�f������������õ�,IVQ#@���0���E�Ek���"@���*@x���ӂ�	�^�	�ݦ�I����[UŁ�;�`���?71�#JE�������-߾���Z�S@3�mI`���pm�^���h���x�~���>�ŕ�z��\�!	QN!BHf��sll7��ɪ�Q���cT�`�]��r)����)�{�,_� ��Ɓ��AĤ�NE�[e4��eh	,F��U�&'�1v%�^���`���A�h��Z�S@���@��h��F?�OēM9"�X��|�@Ib4>���٘����h{�!�H���L0n��Z���m�?����X��3�~v���jԚlt7N�Q!u<�WO�(�����;���sv�[bL��::�69���o�}��/@Ib4�� ��Id���ӑ6�{Ϭ{����bCo�s��@Ib7�T�7UP^�Q86�z�}>4k�l���>���e�L�LM�9���}k@Ib4��e�9����������@��d��I�6��@��h�M���Ł�;�`~$�k�HI!�ȯ}���|i��C>nfI�a�Y��]�i�ۏf�Nk��r�Yx݉�2���v��C��ӗ�L��u���dz��AmY�Ĭp5�O[���9ի��FG�j���ş���w����R�dh�wb��݌��[z8q����g��[��f5�ٝض��'K����V0��qlm)8L�yWw&Ʒ��������iG���!�z)j!3��33\�.;����<7Ʌ�rf��n�cFu#pޛ$ȷdxu�°�|��6����}fD�"��s$������@��h_U�[e4z2��~$���e�^���o�&b�Nӭ���>�lz]�!�H���L0nW�h	,F�Ɉ���V�^���h}t�S"�0pn&6��-����@�b4=31I�u����̌̚���*��@�����M��l��w?��m@�1*i��,��Ř��E}wW�x����'?���#i���vl�D6[2� ��h��h	,F��ZYz�;RXI�I���"��:��{��������E &*!�U��P8�&���V}=�M���Ł�'H�� �Ra��"�-����@��h_U�{�BE�`����4y��m��:��@��h��F?�Ođ�j9�m��>�~���}���=�lz�p�R(ۑ&���-q���z3=��=Y��)�]���n��K��6���D�G2a�p�:��@��h�=�)�{�W*dY&���Z�)�{����S@�����A��Y'�&D4�I�h_�G�^��ɀx!bZ���;y$��)���%���(�pnH��S@������=�lzz�RdN	��q�����oǀu}�z�h^I&������%��,t�U�:��G���.�θ�0�Ɇ4�pmd���B�h����;c�/YM��}��FM̑�!�{����S@������-�ː��$jr=���:��@�e4y��U�ȤIds&7zw��������uM�JI�Z�k�g��
����5�S"�0pn&6��,F�����{�e���Ɓ��V���?{�lq�����Z�.R�U.��􃶝��iǅ�u%vHn�ts�9�WFF쪻�����r�h��9���9����,GQD�ܑ������Z�)�{������Ď�}�����r)���@��U��b]_�G�{~����H.HH���
E�.X�����f)<N����&a!72FԆ��;c�?�fLCOY��:�,F��LOv*�N�ѷ ��]c-�v��n�7`��Nz�6�_`�7mb��˸.�rZ�T�3��(v[�Ark��[��N�2��8�Mc ֢5��c��K���)s��6��^�ݸ-���ց�����6���]F�v��x���<���v��Y.�`ݴ�,Ig����e���.�m�c���[f�'�fL�������v�u�͊����z���A?xd�r~ש��/jr���Z�qT�X�j��5Ǳ*˥=K9�zSuc~���v3@�|�@\�ɉ������M!�H���L0nW�h����;c�/YM�g���;���2&LN�YwyZ+N������335_'��/������G21�2`ԋ@����u��:��@�e4��	�9�pnH��S@���?f_��xW~Z��Šz��d!c��E�]T������ȝNű��pr4��V$..3��7��$s��C@���@��U�{�,Z�e4;�Ar8�Ŗ]��'�s��(��N �<D!�l�hl���}V�ﶽ"��s$Dqh�K��YM>�߳���~ZW~Z^�̹	?F��9"�<�)�{_U�^����ŠUz�2(Db�&'������=�-���?���L4��C�$�+��������Q��P=M��E��;�u���߿~�պ&D��q1��}�?���b�/YM����$�_�̌iɂ���t�h����}V�z�hyz�`�7!N9�z�h����xk� �B�OZ)��?�ʫ�5Q����ӒO�}��y!��ԒRd�qE!�{_U�^��ز�=M=f���P32�"L1
E�^����Š^����Z{���I��H&� �ppC�Uĺ���+��{"�Z����2�s��w{���0���#jC�:��Z�)�{_U�^��^�̿���#��rE�.X��D����:�x���YZW�C"�%�̘`�4k��#GU�c��x���H�2�(���*˻��s31興��?~�&��y$���I�b� ��h��s�g����/�%���dcNdě���t�h����}V�z�hs�o~ D��ն[���j`vp9�Ӷ�+v����資]ds[���7D6F��\���V��bLLǦ""c����h_��$��$��ND�{_U�^����Š^�����@\���0�)�z�h�K�z�h��h��fD�#&�Hڐ���~ȉ�K^V���h+�Z������@�XϿI?�,NH��S@_b��s�_�O���$����o$�� �+��TW�� U�tTV�
���*��� �+��TW��TA?�PB,E `�@�@�T�E a@�PAPDE a@�E b�E b `�E b��AP D@��'� ����
���*�� *��TW� U��TW��Q_�@E� U��TW� 
���Q_��PVI��[߹B�K�` �����Z�          OA�  �      ���T '��B��H�U@J�I��BR P ��R�  "(  �  H �  ��   � �(P(�@ O=>��]C���^�As� �=��e�������k��&�� r��ϯO�3� 79q R�8d<�ru�ʬ >��,o}��y3��ys���p  8   H�����m�}�]���퇐o�8��>���� � Y�  �������\ =9�{���Y�c��\@�s� x�_K�>C���Ł� n�9��F��N���x �E   	I"�� �>�{�9�w����7���� ���ל�N�&� ����t�� 4��@ 3J(�l�Y�f�E14��AFF���`j�`����@R��JR�)JPq@(  
(�� I� R��AF (�Af� )� 1(Ҿq}t9:{�y��� ���/=�j��n� ����]�W{�=���y�y�Ϛ]��N��zo{�i�2��8�����9Y۴x��  
I"P� {�m�==�^^�ɮz�<we� n�2u޳��{wo]���Gp ���7�;��� ]���ݼ��OW�Ӟ��݃�^����yƗ� z}�_m<��wG���������=���)�R�@ 4 ��B�iR�  �'�UJU=M2#LЉ�U*EQ�0� *����کJ� 4ha�� b<S�N�����q����w����{��@"��B���EQ\QAS��EQ_�E�U��(*��I"$�G�t�D.[MB57H1`�!#�k��	-��In�i�R�Ha7�����-k]��z�<e���HB+Q0�@�z<iC�I
kN�|������aF0Ľ$��9�Y�.D�~ɮg���fr��3&��f4�5%āF"!H�Xb�0Ѕ�cP"�00�
��b@`�奈Y�W҆��H���C�@�!��Be�p%%�4�����}���f>�!"R.���<��1�4HU�4�B!@�O$��p�V�*H�����@��<��������2 A��,�"L�x$�8s>׎L(��4#B4cC��3t�L�H�˰xW �0��q!N0��l��L7&�̴��e�x���zC�N<s�ɦ{x��$r��HLI�˙����2�1)���yD
	RPb�R2!>�jQ"�Q���|�
Of��J�r$O_�f���r�l	��~;�8!��	F$HB�@�@��Hh
��`@ �`F!�ŀ���D":J�� �V� "b�H j�P�����`i��S ��h@�(�j1(�b��1��#h(i��"\_ЉGrы �x�`x�Q��������J��$� �c�*�Z� �A��!�SA���$)������� HX2\]Nj�B�	�� �`��#�`e(hbD���@�D��E"�&���
�BDsym�\��5�� ��Ia05��4(jĮ:;�V50�`BP�CC�)
[�F�i�B����0J:�*hqMO-�&k�p�� @�C����D�jD�$,vaD��"RaJ)���i/3�8�>S�Nz�]{,b1#�$lR��!�{�0 bD���H h!
L,#U���2\�fI<�+���M��O$c���ȑ�;[ǖb¶�6�fdZщF$��b�B�+	�w����xF��@$jpQ�	 b��b�F��c@��B��=5�
�3NS����s8�mM���l��$�y �80�r���7t���!B5�ׇᰩ��%eH �O$Rx�²�D��q�0�	�`�4�x���r�p��5#`��56,|`V10��e�����ߥt���.$
�R4(a��d$`$%7R&�`��d
(nݻ`E�_��O2�Z1#���v$��/��80J����@���yOO_]bH�G4�����f�;m�8�B䎐��l#fk0���B@��ttO���0���_��y&\[\ʤ���4��_}/XD�N}0>����q�]� �(`��B�=V#N	ȒI�Ș.?1�#B�C �Cx�8��>B'��e���@�Ą�!����y����{M�NsI��s��Ç4��N)��/�^yxT>By}�ͷ��!��OI�K�=	t�ᐸ˧!��3�K�������%H�$rF���-&�i�)�7�y�1Ѕ�_�m�ͅ4#L5cvL!p�\&�Ks=�g��s}|<���N'2zL����Z�K�$*/��\�g����g�?_Hz��-%�ԗM(\��j�Ć&��ӈ���<��<�n�NfF��"L�\�%P��
1�+-�B�@�r��ݳ�׸��.�����{�m�)aYJ��������#�-1��(JR�ԋZ�є�-���1�+!s+R�	R��+iXT!T��-K+%V0-�C]7����}��E�}=76}<g�#sf�tۚ���d8Ce�zK�y=K���	�=0�Iއ�,��w\��<��C���8�,SO|@��\~F$�˛� �͆i��4�=����|xh�^�cXH@̌(A�pcLL�B`B	U�$��p���"U�L3F�\�H�d3��4�.�B���4�N:���B�aRnCn����<�mˤ.*�B�F��HI�y�f�4��B�Җf��|XF�^$+����a�'�X�ą)1}$H��dd"Q�!\�hA�@�����錄B@d�� (��hdJ�	��)��eXѕ!B���^S^�p�Ë.*��L�6qk$�R�r�$u$����i��8��k�1	���H�	��x1��@���FF��(c��Kp�.�A$���h�`��$�	/.@2%�C���L]C����<ld-1��7�<>#\5yhy,�K�\j^�11a����	�Q!��2��,g94-XT<u��e��/9|���|�/�B�LЇ�.;��g�hp�)0�䌹��K��3Ra�,+hA��`%xƘ�`B䒘0`���B�k�yey�	��B9��B6L4�^4�Y]�.L��$J���9R��t����0�7(�����c@�!QbS��9����������ۣ Bz�,Q���`��_A0��Y�4��X�XZ�\&i�T��,+ R��@�R:�ki2�d�s�Ń�V)d#�*��`��~J����	(ڰ��򇒘45�.j�i�`ƌ�.$#�d�l�y���<1`WY'�.�	R0�\�q�~6�2\Isd.ɉu~5.����
i��K6,���9s^P�zSM�N:d�>�i��3�CU9��3� Ɂ��L�����	r6CF�� IV�A>bU�_�6�=6��.�'��A��t#������|f��XX_<�{)��xJa��+)�\	S	p%aCS�x�=RF!�3y���i-��t5�{��"||������'�����<'���<�"}B���Ŝ��!�}����||xiÌ(a��o��S7�k'=�`�缼%���y��o<�����M�S�x_�.���|��\5�C�s�7���|�`��	��M?1����������ǥЗ�Y��$M���a��K	����9�7�%1�N��a�Q���L<�3͹���Ͼ�
�q�~��e�B���
`|�r7��pǆ����_3Y�o���i��OM�y풏��'=
n��4��}��8l,<瞲�.�>1�='�'�����p��=���1��3
�v��D�Ӈ����0�����>5���7�^p8[�d���=�r�p���}8p���}z"����$jb���HS�����&�8'��F���0�Scg&so��3�Of��ǞzlF�)�A��7Rf0��!^	�NG��#P0%����S�i���a\6֬bg��k ��E���2%#!B͗7�<eӃ8�!�=C�������JT���1��*$8�pF1c!F�Ҭ�Q�S��yĔ�8�0�xًS���q}0NM=���d%͗�Y<�!�� W9�'�pՅ�Ͼ$�H��V5�Os�#L�Ç��Q�+�������<ԅ0�xz.y�1=�g5�������       �       �  �    � $  UP�a5�%Bjn��Kr�l�E�-��K�����c�?���`^T'�]�����t��V��d������A�^`UWU*�
e!���:�` -��+X��r�ɱ� � -�(m�P�m0 M� ���5P- ����ն�p �5�� �H5(�ڶ   ��  H$�� �[@4]���mh��	 �a��l�0 �h  ��  -�h  �l�\�]��ٯc����=v�H�KŌOϙ�phZ�T��m���wmSeX�m�  Jyi��IPm����X����^k4����dҳ>�U�UR� 2��ݥ8 m�b�&�����h��"C [@ ��kղUE�D����$���I!ŵ�5_۳� H	���E �e���$�غ�#m� m��d䷉t���� ��Z�*��6�H�<l�\�@芝m��p��d� $����$�mエ�ѻ5)2K[U=�.�D�;������ �Itp6��(��b��ᶫؓͅ�z��-�9u2��]v���M��9઀�Rê�m��5�r�m�4��d  [sG_Tݰ� [%[!��W���!PUQEC��p�K�iq��[�䉥�UK�R y�tҬ�������kS``s����׳��lr�,Iɺ*���Ҏ�&�)ҫ[^���n..k8$����[uN*�X m�[��5�U�gZ�l�	lˎq��Yr�ʺ��m+U��u�n�[[I|�,m���*�ն�p������P�Z�V�yP$�,�q�mn��m�@T����x��!z���Lp MRkӥ��� s2�AKVԩe�U�u�N.��$�i6���鶷�KZ�l�@#�7�[������q �u-��� N�Y՛]��*��-���G�L�d$m�`m��HJ��$qmr۶�#E[���;v�r�+��*�UU*�J�U@l�U_l����	����[����J��kh,����XEr�v�mm�@}r���@�^j��sҷ.us�ljz�?_|��K�;jY]����)`sm�]/(�"f]��ꪮ�U�.Z�xUU�N[&�Sm� m�   �-�$�Fi*��k�S(�p*-�i^`#�f@�,5�5U���v������&���E,���8��m�P e c���UUs�m�� �[n�h�;��Vspd���lF�+UI�8H��TV���v�lU�YN�P+jWf�j�V�k��GлQ@qtͱ������v��n 9�o��V�l����V��4��+J�YYj�Xɤ*�ڠ%'�6�ٶĂ�ι������'�(��U���E��S�ڥN�����؍m��l6 �d2mpm[FG��-�9&6��U�yZ�ųr�QuS�.���V�v�W����U9^k-���ҭZ��V�2-US�U��@� #�jΣA�H��j���t��`�2y�m#��.� #����RI�� �   	l�m���.�H�%   -�
��@��^@�h�Upr�P���ub��$���wi��p6���K,j�iM�,�����%h"��t���Rl�qsz��B7<X�aj�A.i��%�&�@v���n�%@�v횴�p����	�U�h3�� �]I��=����{,�U��c��vnZ 8�F�v�"���M��Z��[t��rMj�V$ l�-���'6�Y�[ ��)R�6�m�!�1��I ������'��XH  �   �  d�	�m�{h0	7n�������l-;mm۴����� [@�V��S!+�g��g]��pn��` m��h  �|���H�U��Z֕�� BC[@P9�]��@����28$ ۲Ś6���� � l�V� 8����ր  K��p�NP �"۴��$-���kh&����I�޳:ˀ�-��K ���m�L  8�lHR��
U��Pa��^'��T���+b�Im ����  ��P��Nڸ	e�a6���JۺL�it�`4^6��&��F� 0���H��Sf[l�mz�+��ܥ��� �6���kX��P! URM����UXNG�l�2n��$�'+�[#2�mI.9{27$����Bإ��U��1Q��]��O���@AJ-6��I��#]v �l�z�`�h��n��p�8�p� �I�[~ݶ-�%� ��m��-6�v 	���k��H0[ �_}A��VtM�Qz�� �M�݀ 6�
]�6m�k��
yZ��J�]ۢ��Ь�g�f͜��� �J�`  t�"Jmz���\�m H[@9��fՒ��u� ֲBM�:�,� ���8�!�.ݤ[n�v�m��m'ɵ�	ӭ�n��[S#Gn���m��h hp9�  $i��l����m�H�`��gm�X��K,�����JY.�a��;\[@ ����m�m  H�  �i     D�@  ��-� [Cm������ �g mݰ-�        m Hm�ڕ�  �@��� �ӆձ 6�E���h����mm�[';  lUY!
����bT��;&�ʶ�]uU�Ӱ	�O���֠���-WT�L�]�e����$-�H8	z�����E�f�U�V���Uj��M�GG��l��@�$  p  ����     �   $� � p ?�H�m� �  H          @ `��       � �     8m����m�M�[A��m� n����mH  ڶ6� Y�-��F�d H  z�$�h���$ �.�q �ᵚ��l�IzeP9v\�uUR�]uR�� ri�IVܷ�m��6
��"m�v[�J�Ҩ� ��$-�l8 5� lu�l-����$�C��gl��h    $p  �amH �� 	 m��@      -��[@ �   8$      @l   � -��[@����@$    �8  	 �d�$l��6m�m� � >>�� vհ�$�X  H���� �`mm��]��	5��J�x`�[j���� Z��2�]R�Um km�9@.ʜe�N��8lM���H��[��e�m� -������  l   [@  �am   �    l�  -��   $   s���  $q�{` [A :���gI��m���t6�6�'m��� -�m� .�4��������>t\;l	C�j˻���U5�5UHM*���$��z�l-�h�p�    -��5��5m� m�@X-cj���U*��W *ʴ��UUUW)k��ܫN�)ۯ^�V�&��S��9��6����\��Pݭ�!��ݰ i6��:$���	Oj���m̅�6��oI'4Vݶt��.面I���s�cni���e�ݗ�6�Ƈ��)[��ɋ��d��:�B �U탩j�ܪ���dZ�����"��J��NL�e�T�n��Ђ�m�$��m)[l 6�   Ař0Hp�d�H�t  �z�7m�p6�kf���	 � im�v��:GH  m� m�`   �M�M����n�m�m���Hp8�]k[@�n��l�٦Ŭ��6� m� 9&ݳm�hl��6��]�I3m� 6�cE	   m  k,f�۸�H ��մ����[p   $ڴ�մ�@ݻ{6��aJ*����<@'T퀶� $�Z�������]����h�6�:�7j�  ~|�tp$` �l ��u8Y�m��Ā���C�Z��\P����ej��jX%v�a��$$���du�(kn�m�� ��tV�l'MN�S�6y��l�A�l�f@�#��ݤ�E�imp�P����Z����9Zv� t�趱�$m[����q�$��n���m���
�
��R,A��A � �D	�`��z��Q �?�!D�@V�b�)��Dת�P�D��D�J��(`'��"�>��E"@|8�*�`z+�`���pP����&�"'|�~_QP�S��0���:����#N�N�DX��'���!��}Tđ@ I�B�j�Q �"UE^��z�����
`>�<@�# A�HH
�D�t0} 
��U< uš�@�&���=�E ���|"���⫪� 1b�}T��C�}E
��T��%=O|zD���OT�QO�O@�QC��
`	���C���E>��@}OL� ��G�+�#�� �(#� ���E���{��A>�: E8
|4�a��C�A��_�M=x�ʸ�������z�|a���Pӡ��Ex#���@�AE�b�?��@m�� H�i�f6KX�Ǌ�R5���Ӣ�iIa#gmB�: ��J���#1y@��BSj�M��q�v�9fVڥ3u�v��p�gJ��:�����,l�8�g��XӻU�5��e������6��ݱ��m�^NR�l:yIƪ���@m�kl�@ �Ѳ"���\X}�\'.ۭ���[��Od�c+�Vlhl��	(�ҷ��U����&�z�YH�Nݗ]=G n�v�z]�E�.���9m�E��&�y]c2Ʉ�c�6��u&��&��5�n<�Cֺ��٬��܉
�M���='�LH��*Vuu�l9E�+v4�I-4j�<v��&h���*Pmؤ���v,q����e����[\�mI�!Y�;;zX0nz�禠��K�#3����U�[��[�^KkS�ݞy���&u͞�G��`��9��V�G�����N��$�&���I9VWCp6���svݻ+����.�S�B�ִ>�0]��d����lN㱊7S���Ki)�M�<�H�9�nXp�ku/ucYӝi͝��{s�vY@Ll�s<�ۙQ��b���r�S(��d�˗:����ðf�r�h	��PO<<��£[u3�m:�Z��F��%���m�N�I��v�h 	�I�j�Rvm��n;u-�J�;=1�-����N��ʳ�m����gvY��u]z��[���M�`�b�a#�I��z�W�KL��q��2���+T��<�a ��E:-%�m�
U��%�� m��""�&Nt�O=���{8�7c�GK+UV��$�\s�0�J���א�4;��p1����@)��hM��28n��s���Ue�5E��v�P�X�a�0�D�n�-���s��U�%UP�.e���C�O�*l���q�p��a�S�v�P(�=N�r�e�7V4\U:u���M3�X{M=��;v�b��?§� h��D����b��@
�
���Q8���J��@���f\2}��Кc[��
P�6�L[\ם�E^|�s*�ޟ9n�؋[�=�v�@�T��[	�nX�v��Y`��[�<�/um�V���l�;�e���)�=z\#˹����j6�^ ��S�cs��"
�R��'pp�Wg����vp��7�5r���Ԧ�z�`ЛtfW�s�n�.d*��aIҽ��;]����wy��{��<�m� �G���e���|�ppr�wg��q�vP��oc���U�C�z���P����G�mLr870Ȝz�v���bX�z�$����}���:����~g���Nb�4�Z}l�=��hwW�}�j���+�DI'F�UVd�V[�l��6�{�I빠}zc�$���&�Z]��yڴ�٠{Ϫ�>��WdDx�E
Ksa���b��\�t�ce��h�wH���s�Ĕ����$_������@/����������*q�"s.3s�I�{��!�ơ�� ܟx��@�����^��`�*�ɀ�U**���̝j�i�6rX��l�����¨OS�"�ƤZVנ|�k�m���� �=շ1���E0Ȥz�ֽٟحvh��
��@�W���ư�PĆ���K]��6���ܨvlGm�퍹R�q9��h��2)�nG��4y�ZVנ|�k���+�Q	`�d�h��
��@�zנ�5�ff$}lǖI�Aa�&�ZW��>W���LD�VR����B��@�9;����{��o ^鎍ĤY$�������@-�h��
��@���ǍD�'�8��f��}V�U��+��������{w���W�nnb�����r��z7g!��h.g��[���oh�{��6�{Ld���r|�-�k�>W��z����T'��8dĜZW��D$b��`Ϫ�ܝj��n����JH��U�8��{8����s&$���w_ ׾����}�ΧDꮡʪ� o]X��X=s`DG�����x_� >�[��g$�����85� 8��������/Z�޳@�=l��&�0p$�S3�ι�7<��.����@�˱�q���͓��w�-��d���,MȾ���y���uވ��7e�;]D�UDA9?��=�;V�[�h��
�W�}]xQ��&Ԋ'�8�޳@��U�Uz��;V��cW
�Ƀ�99$�Y�ؽ��h^�@��ՠ�����T'��8�bR-��l��6���Ϫ�̝j���j!@P� �����%�"F,�cB����9y:\�(�\<�p-ҍP�f�rz��T�rGM�v]�8=m��}��*�Y�E����pv�G��Ͱu
t��җm�d	y볣c�q^����#���r����m�cc�Lm�u�w;��V�1�yvܛ��Rv�r���A�	�j��[]�uH����Dc7k���m��mT��Ki�=��j��齶0���X��v���)��~��}ؾ�8mNT�Ɍ�šB����]����»��/Zu�)�n��Y�L����s��h�f��>����ϐUez��U��"A!1��zoY�{Ϫ�*�^��^�u�T��B� (���ֽ�����h�f���Y&5,Q�ƣ�@��z��ZoY��ϭz����"RO��@�>�@-�8��{8_}��bĻ;��[X�+�[�㇮��5g�<�n��0m)�#;`˔pd�8̎DRY��(Ԓ�����??{٠Uz�����Ʈ�0d�H�7wy$���� (~��꫖e���`k����V�Б�o�Ц��*��i9�U��s�޳@�u�@=�է1���	%#�������w>��̀��6#Rٕ-�TZ�nZ�����5%��,������W�{�U�{l���#a$M�@�F�Vtѧ[8���3MX�t6	��V��9�H�L�M�ֽ�����h�f������d���i��D$k���;�U���������D��n8�s�޻��q"'�Q�� �y��g ��w�{ΰ�ǉ��8,mŠ��˭zW��=Ϫ�;�+��L"� ��@�u�@��z��Zm�@�\J�$�(ۙ&	��M�D��i�tm�Y�t�������[�ٱ'�����������	��Ei9�Uz���� �٠|�נgZ�1���	%#�3gZ�۫2u����G���ԶG5��U�&寀���y����u[^����@-]E!BD��d��7�Ŋ��������g ���_D)�| � �gw��I>���;�T�*
�(S5J�i�6{6���߿M�}V��q�jDy1����������x[�o�c �1��c���y[��/6nDC"q�7��- �٠{Ϫ�*����5�1�L1��6�_�{��L���X�zl�[Vp�p�)�$�qɠ{Ϫ�*�^����@-�4��¨OS�R(cĜZW��>�h�f�����N�@=�kc�dp�N=�;V�w���<�������=ŋ7Ħ#x��ݻ��=����Xy�u0욠�hgDt�s�]c��]N9�˜�)�W]���J�x�u��Z�[�cs���\i�e=gv���=���Hv,獛ո��#�on�xsź��lM�ZHv���%��J��8u�kH�m�Uge2��\E�/FY��xp�ە#n�
�M�GO�6�a�-0]���5�y�X��qa�?��wu������y���t�9�мfۮ�7n�����L��i݂�-n:�g��TcG�y?�߿:�3'Z�z���%�`�H5IH&I&��>�@��z�v� ������[Y �IH5Nj���nl�[V~�z!#��X��h�1ѹ�K$��)#�>�h�f��>�@��z�ׅkc$ТjiXz���z#v�/��Ϧ���ՠw{$N�
B$��0n8svdܜ�&���8�m�:Z������<K��$�P�HA�&��>�@��z�v� �����%P����Pǉ8�����"�B$B��;��m��{Ϫ���mF�G"`%56�-� o]E����d�VMנ|�%SL��'2cƜ�@-�3@��U�Uz��;V�Z�U&V:�m��y����jŋf���y��| �}�\RX��V���d�F�V��Ͷ�	N�w[��ukg��:.���ˮm��a$�Y2c ��|���z�v� ���3�P{Ϫ�/t�F��FH�UzUMM��Kj��䃹�E��/��U����*q�h�&��z��'��ݼ��E	�I�WSc%�=�K	��IbP�!a�ĈFI�H:����)C�
�	$FD,V�_E�'hf_��'��I	�!HL!D����G~�"�OσĊ���,�R!ġ�F_�҄(U������*/E>��|��*'AU1QEa�C���(x��}Qz>O@8�� �|��=�ė���|�����覨�WQm�%���?}���5�vjX�0�ٺ�~Ēl����=�Dޱ�8�lT��b$��׽��Ēl�ٺ�~Kf�v�ﳺ�,_�|�%��
�}X�tҌ���2ೞ�R��,�ڡ���zeI�LpHs!gق�U�p3�����7�����?$�wj�����z��8��O�z޸��D�UE��w�W>�����oχ�X������{7^���0�P�����m\�f?}���?%�f���y��|76n���<ݰ6���Sqb�����ݜՙ���^I<�����I��'�'�:����~�=�������cQǠ}�j�=���@��W�r�P����䝴�`eUz�d���7�V^��;6�ݐ��Z�H��68�D�X�"H qŠ���>�{ݟ�׽��so�f��􆨶�9-c�I'�^U�����1�{ݜ���ԗ��v���މ�c���H�NI�~_��{�U����u�@;��T�C#��kq���h�fh�l�*�^��r\��rE-*j9k�k{�ڸ�wn�a�{���?{{��|�k*hw[��!"(Y�#F(ĥ̠�X0�%A�o m����J��=�u��p`�S�\:7k&DW��r2�]fd(BM�bc�7b�s�.�l��훂��[�yv���{Xpue� ��n�6m�KfkT���:9�d���X|
d;\8��.)�\,G
���A*�j��s��N�޴�g�j��i�F�Lsv�n+[�2]H����wc�q}h��c�r�J���;ׄ�Kv�*r1�pF �kN�g��/�n͛-���m���I7��^�{�R_�{��|�1&�{�p7l���i
�y��f����gu�X�07{�p?c~wv��j�;UE��ۑ�g6!#\�V�����>��t��7ٰ5�K%v�K+��w�W <�uX=s`�Ӯ�+��0��L�I"�j�á,}�`r��� �/��n�jԿ0�3�b��j"E"�N�u/#ӻuwV�Y�iw	ΚU�s��:�is�݄�\��*A�o�{7�8����Sf�v� y�۹���p�جi�g �����%�X���$�H}�U�>����_�k����KrC�u�����Wjr����\ ��{x|�b�o^�g ��~4+S��j!d�Q�G&h�٠Uz���s@-�3@�����4�jH��*�^��}V�[�f�}���fu&/��F�����g4�c@���tg��'+��3��6�96�k�[��fc#�&L�)'�RG�]��޳4�hzנ{ΰ�Ɓ����@/u��y{��*��@��ՠ{�\�VE�p�	��y{��;}���� qX B �A" �j�:�fo���I'}�t���
�lM�P��H�=���ʾ��yڴ�����^�[��1B(<������޾��X���_�����@��^������	�"@�M�]�[�l�Ő�nlG�ݷ�v�"�f����2B7"NdȤ�@/���<���{��>�h�'S��BD�8�$��y{��fbENנ}�j����>�0�F�M9�%$z^��yڴ�Y�����LtRd��ry)���Հ=�Q`b�sa��FB�w�͜�&��)K-�"Y_ �Q`LG�s\�[�l�[V��ǿ!Y`{BI��3�&ލ����.'0cn�h��6�n�s�k�yl����,�6X��d����$�lM�P��H�
�k�>�h�4/uzoT� �X�Q��z�-� y���Ś��k5́��9k,#d�Lxӑh�Y������67���k�ME*BETS%93@�Ϫ�*�W�}���4�����c��m���9��X��i�3�Ў�wUθ6�r�������\=���mV�e{:�����.!�Hgslt����l{b=pO���ٶ�;C�X7��]�֌�b�.���V8�[�|���s�Ξi�n�.r׌��ʵN�m�����d��ǘK��<��Q�g�9�u��l�][�ר�˃JN�ɝ�e��uW׋	4&�������O���L��TM5;q<��nn����q� j���-)�dY�Rt8��KG�o����́�m2�k���f��`su�MD�)r$�z��M ��3@�Ϫ�*�W�}ΰJưrH�jC@k��>�֬�\�f�,��l'D,o$0�ɚ�}V�W�� ��f�_[3@��Ĩ-��B	
E�5���>�u`��>�֬��~P���7�NI�7]jۛ�NS`%�P͗ms�xݖ͇�b�K�p���u�}l��>�@�����s��l�TԲ�������3ǃ̈`� A�=ȧ��D�_O�+�>� �5Ձ��eME)@ը�B�W �����u��g�X�l�_�@?w��4�U+$k"b��dNR��s`5���7Qa���O�������dB$i���q�{���fhϪ�*�@�����&������>�1��d��׍��Y6����qNzX粩��`9$�b�G����/�U�U�^�W��خ\n���X9&j�,��_G����lZ�l�$v�%����"���T�M��N�~�rO�H%�����t��s� {�z�:��N�cN[8�g�������V�]-���NepUF�����8�=�\s7�����vh{��p��l��8�jE1L���7u;�u;�:��J�閳BG*��v�X��o����D�b�0��I3�?s���WuzY�{�k��Q˪Q�EU*"��+��7='-}6Ϻ��y:��f��M$�����#������|�j��_I�f���w��?{P�lh&����T�M�B]��l�V[�l��^A~ �r�!��7�����5?W�Me ��,���'�X�Nz~��� x�E���[.�wD-m�D�Z[Xz�ݵN�˭���s�z*�	�a�����_x-���=h �������~{����j�_%�~�������[ 7l��e��罜�f,�% }��\ߦ��_����l��=��[�:�;,���W ���_�%�g�ߜ���5�~��ﯥ�WMZ�d-�p71?6�_ �����=��|�Y'ۿU�>�3���4�k�,���;��5%��v~ ��j��=��L_,^<���C��*BE�	I�b`���X�
���� b�`�� ���
`1���,���Q��F��@�# ��- �+�ˆ���HK��)����^X� 4�X	�EH-D�!�b��0|�X��Uc�U�%KX�)@��
�$ A#���X�"�+��!�&4c1"�`�1��	0#
d"��FB�quH���1 @���� �F$��D�X�0a�$�H@a0"@�+�x0�1��+��.,3+� ��(�����)�!��� p����}�R����z2䙐f7�V1�
�zǢ�T�A�YH���	Kh���4�"ȍ�bk�HP�	�����w;�w���?F�� 6�I @���%��E�.-�q�z������n�ڹ.��Cm��꺨��ڲ�P��uf#s�P�&H�Fn�9�׆i]$Gh��ҥ�.�y�z�C��k;R7nO6�qPb��{	l���<4� 3V���9�Qq]۶e^�V��V�v��]���,�A1�Ȍ�1�QnT3\E�q��m��qnmFn �Jq�(��Q�N���ᴙ���2�'Ap&�]���I�zκN����	�rgjl]�)�'d�b�nքk�F+ا�"��n��k}�n���.��t�T���Z݋d����=fιs`+Kv��"�I���ÒNfժ��Y�$�Ku=����J����(�I�.v:��]`��k6���]�ժ�P6�k�r%)sێ`7@�+�c�V�ZU���Z�*B )�A5Q@��q����Q
���!��R@Ҳ��7ewFѸ"{<J�;�X�"ԇ�X���,��� ;��@=��5�v��b�"�v��������h쇴^ 4���݋z=h�<�U>@&A���q�m���u��ᜲ��l���U-���� =�x
���8
��UUl��-2��Im��.΀X����O��v�����<�,�Mv�3��&Ե�*�R%�N��w��B�p &�U &��Zں����S�(/l��ؖ���^���wFh݀��qrJmm��@8k[�-��a�m�3m��I�N�u����v����k�\�����)���8;\۽�Cl�M�h$�$ ����d�:l�Ӄq3y�G<������Ҽ�1��N�܉���iL�V���ڦ�+rmu���;]��4�ӜUt)��«d�SPxj�*Lt�Ntum�����+]��/c�-˒��#�g�X�+Y��&iOK�g��))��9uI�qX�=bj�+���T���v�%�)�(�芕b((~J����z*�� ��)�~�F[���n�f�n�W �5�sh8�S9څ�^�i�w:
�ZMz��bq��Zx'Nd��8�Ͷɝe��Z�Ë���vng��80k��m�����?�ݾ��Y�v�A�_+�z��p+G�ܘ��MN{fɴ�L��({лI��3�#T�^s"��ؐ��Nv�s�Z��O#j]�Ea¨v�<�GA���$[�����~�������cs�5�A��}�۪8S������%��m�cn�d��a����b�U8KJ��̍�:��Ӏu�X9ֺ">A�{��Ε�%�("[m�;-� ���bQ%�Zz�ߧ ���Ӏz������z�I��h���ڸ�;��u���$��&��Ӏn��h����lS�	H�
�k�5f����Xt,�|��k�q52�,i�g ���g ��Jof��6wV�U����M�E�<db�##����Z6l�k�[���Hv��n5,u��Ĩ�T� ����q��fhW�hz�}��_���:�^�*��j�[!e��O;�v�T�H  �*-b=�G��iۛ� o]E�ܡ� �D���ZW��9{������H�Y���Z�Ltr$
?�SU6��6 ޺��:Շ{��]7�8����D-�ڛ�� w����}V�U���]�����"����r&���9Y�s�&W�OJ�
q�:WX4y��@G���b��oLN�c��~���z����q��ޏ�Ө�o�x-�b$��ĤZW��;�w4��\�g�|Ԓl�ף�DB�cMʛ�� o]E������<V��+������RL$k$jcȤ� ���������}���@<��dS&DH���}ψٟ�Ϻ=׮�[�f��.%u!̘�dd!��,�7nwi�n�X��Z�����v����[�șR4E�L��a�@����]� �ٚ��Z�Ltr0H$���빠�3@���@������x2H��73@-�f��}V��J�+�;�w4�r�(4�7�����:Հ�nlͦXDz}�А�	2w�}���\��&���UJ�i�6=w�����u�6������#Nnh77��' :�S�x�Ѩu%�!�mͶ</i�8��d�LJG�}�j�m��{Ϫ�g�*�^��>,m������'"�z��=��h[^����@����LX�B�293@��U�Uz��;V�[�f��x�cA"m���#�hzנ}�)��3@��U�[��Đ���8��>���=��fh�괓���rI���Q�B�(�_�;p��onxs�נ�6�Z�vj+�3�'6Lfcl5&�^3�|��n��G�.�v5�ێ� tWg����^����d#�n{/Js�rj�mP��^�Jq.����Yy �p�<��;�@��4�"ë\ru�V�Y�� ���H� ұ��U��7B��k��m�uъ��g�D�GL��P�hL�J�dtf�(���.�ْ���D\U��.�7sv{Yn�ʮuV���)��rحԾm�=�I�6�w\n㮮&ܲv�
�l��t�7�d�VO\��{� ͞�`d.�ԩL!L�Q�UE��:���9s�3g�h�fh��W�Fds1 R-��l�[VbCn�,�֬�jb��@��cN[8�%�{w_%���c����pA�666?}��x ��������lll}��~���7r��t͹�x �����pA�666?}��x ��������lll}�~�|��,bı�ǫ�'�Jɍ�B��P	p�אc��
�'!�Ά�q����3��<R�Zv�0��\ے���� � � � �������lllg�߳��A�A�A�A����� ��� �`�`�~��8 �iOۅ�vۻ7iw7o �`�`�`��?~��|��'�@1�A� � ���yx ������ �`�`�`����ׂ��DAbY�c%�o�S��Q��3ss��A�A�A�A����x �����pA�666?}��x ��������lll}���/���M����f��>A��������|�����o^>A����~��8 �~�߯ �`�`�`�韎��nܱ����st���lll~�{��A�666(E_�����>�����������lllo�߿i�� � �!�X�x���mm8�+VY-u�K��۵wN����v��h5rGi2�����i2[��|��������pA�666>���^>A��������|������g �`�`�`��Y���f�vnn���pA�666>���^>D���A �`��������lll{����|��������pA�666>�{?nfl��Mܺf�ݼ|��������8 �����>A��?���:��� ������ � � � �w�^>A�������se�2f价&f��� � � � ��w�pA�666?������ � � � ����x ��`9����ӂ�A�A�A�A��K�?�&�vn����>A����~��8 �~�߯ �`�`�`�~��N>A���������A�A�A�A�w�����	��jf�h^��c���퓇�n�sq�dݞx5��Sͪ�q�
9���>A���߷���� � � � �߿~ӂ�A�A�A�A�>�����ll��͛�8�,�$��͚�{+�[j��	��`��0��5̀��6�v��W;�<`��<rf���@�����Zm�4w�+�z�$)��>�S���N�g�> w���
��'��g$�|�����cP�E�H���Z+]��y{������lM�FDa2<I�����ZN�\hAs�n^_&�kcn�g��\�}���m���$�Q9����4/uz ���f�r�7��QSB�%UJUJI���1f���������V �u�3���ϟ�&��-i�l��}�������%���!��}W ���8}�S�qd�7m`�A�/�-ZoY���� �٠}]Ǖ���G&8��fh^���f����@y�1/���%};�������۴(��E4���'��l�H��N��q�3�W��n������WRv)�2�����x^�vN43���M�N6�L�Z��)���{D��Ӳ<�q½��lF��`�������b����G[�*�)ݤ��:�)9�5��x¸�;u�V���6�vu��b�J�#��t[7T3nhd�&6ꮉnB�E��}��w����y�p�m�����nn��͹�vs����.↚g�փ!��9�9�u�wc�h�AI�&���yzנ�4�e4�fh��W�F��"��@-��a#�t� o]E��5́��֒��cP�D���>����fi��r����߿M���s#�(���[l���^�^�4�]�����A6Ғ%"crf��^�^�4����|�j��X�ݵKm,r�;4��jwn%��%��FE{kn��MY"�:M��k���5lx�D����? ~��4�]� ��f��^�z�tn(F�#�N9o ��{��Ē�1)}ݫ�z���@/u���y[��I$rbM���fh+���@�u��=���b�)#�ܙ�����z^���w ���Nt�%>���UM���s]ŀ<n���=s`b�{���sU0u8��h�ݹ�����3<��͵�M촒��@7;��GM�����7Q`|���G�9ot��3�Q��Ĝ��&h�fh+��^�@�u��bGWud�	��I�e�ӒO/~�rI���98�i�H`� | ��"04l��@�C�@�`B$�d�$:�@`��;��F�GS����@��cA�	�Rl� G� �����
A���<SH�j8�%B@�	Fa#! B@�C���x�B��.�D�x	W 4j#~T��@0S�x�(uD>pC�>�����}O�_ ����)��U���=�k�>���z��<����c�qB7"�3R=�YM ��f���@��z�����	��n;n��i�{j}�^���ɴ�X���9]g͛c�<i���O����4޳4/uzW�_٨>���=��c�G�$s$�9&h^��
�W�}�)����{��\�m�I`�zW\�c�Xz�,Y�l�Ħ��#�b�=�YM ��f���d�(h�G{��s�O=ϲ���m$�7���[�f���@��z޲��߿�c���3k��q3��1l���N���Ѯ�;sB���R����P�'&h^��
�W�}�)����}GEd� HH�)#�*��@�u���fh+���c�qB4�������M ����z��uz����D�MI��- ��3@��W����;V��+�,�l
&��UTX�\�����6{�$����9$�!"qbT�� �N�ɥnfit˜�n�j��X[���/>��l���=�y�w`�.�Gs4�	fDiV�Ȗb��t�V�ղlUg���mی�v�g���u��sJ�������8A�N-��Bg;�b�)�l�l���VΩ� f�ű*�vL��[��-�9�51��_v���^t��c�n�Ք]�S�x#��m�8̨�\ڵ�I��j�;��{�w���p��ݛ��J#f�1a���m[.�K�+�v:�pЙ5�u1�{(�o"K#�����v� ��f���@�r�'��jȱI����@/u��y{��*��@��U���9�ĤZ{����^�W�z�v���Y�7�)"PBrf���@�ֽ�;V�^�3@��b�b�dc��Ĥ�@�ֽ�;V�^�3@��W�}r�ԅ	�$�$F�_wݍ���;��t�Ccw�klm��o&ys�su�A���7"C�MI>��~Z{����^�W�z����rE&8���ڹ��f/�B<X�-K�㏻��=w�=�;V��+r�F��
I3@Ś��7V�-� {�����AlM�6�`�z�����@=�y �}�z���I=��A$QI�}�ڰ��,Y�l�u``h��h*�.��¥<�ؽ m`�v�5[��3t:N�-�]rhW���۰�]�>�=�Q`b�s`��Ձ�cZ����r$��rf���@;���;V�z���}j�Y1a1G�Ĝ��$���y$���o"PX��b) *��	g���p/uzz�tn,�7"M��hyڴ׬���^�w������q�&8�׬���^�w���v��aqW�D�O��L.j9�f{mɕ�d�&�nУm�g�M:�]u!�"�$��y{���f����@/u��{��POSLm9�<n��[V �]E��5́��LI��bD�DI&����@/u��y{���f���T��%�	��)��b����p_������X�x������-Z�α�����PB�f��5̀=n��[V ����8I����޺ngv.-�����Gmlƛ#p��w<��9�� �����7:�S��u`}�ڰ��w�A�_M�ϪḲD܉4bjI�}�j����=��h����
���I��- �ٚ��� �l�>�hb�r�E�1H��G&h�h���v� �ٚw,�<M��1��[l�=�j�m��{�ՠgwﻷww���ߌ��uVب �gBN���޵��׃ +Wn`S�{y�X�9��t;�9]�9��"�b����5��\'ہ����	�v������.���^V����k�FɷiO].ͬ��h�	Ѯv
,B\v��7���n�6�UY�˳A�ݭ3�,t�����9����6��^��m��c����m���㔪q.�L�[�.mW�X��;�����w����F�nh77b�����N�A��cu$�TA�V�#�	��<��ڢ3U�7<Հ6�E��-� m��>��c���E���{�j�ؖbM�t�+ ��wi����f�*��*�������ZoY�wt��u�3@��DA"8�A6������4��4��h�1Ѹ�A9#��&��Қm�4��h���~�?b����E�<��꬇O;{r��s.4��Hs�vu���.��v�ϴ�UUE*�> �>rڰḿ�Қ�\��18��ɚ�ڹ C�O�F�b��e��>�����]E��2�M�����1�����yڴ��4yڴ��*$�1<	"���@��M �l���Z+k�>�ª���'0���@�n��;V����yڴ瑊�D?䱩�c�����u�����w�O�C/=�K�x�9��뎳r@I3@��U�r���;V�׮��u��%��'mŠr�^��;V�׮��>�@�Y��Œ	�*%T��d��z�,��G�ve�����>��ʜ��$������2u�Snl;��D,��VlOD�LȞ	d�8㙠{Ϫ�9[^���M����{��ybX�x�E�)���˙��N�v�������n@X:�Z�7a�ba��@ȜZ+k�;�)�u�s@���@���D��'�$S��yڬm�X��X�s`d-�^J�LJE�u�s@��U�r���ҚW�cx�D���$��}]��O�{�����I
A�`!�È8����{���w��gm
D�J�I������:۹�}]�@���9d�5%���cA�y8ݮ/A��� \q�c�knLk���XjP����:۹�}]�@�mz����I��䆁�����Z+k�;�SbGv?�����ɨ�3��5=s`nm2���Ł�17�9�8*
�_V,�M�wo m�z�,����k�Jn!HETS���)�[�s@��V�U��I����$�xY	�K���1���`�6#��1YB$e�r�K$��*	D)�(ĄAxC�n�0�VHH0(	
� ��d(��E���U]��1HBJ FH0��H� ఃā\"�$����f$$7F8ah����bE�A�T*y�� 218+
ʤ��B�Hh�H�d!S�7��aB �l�V��`�0��S���H�,kԶ֣�N@�^�D�"� �	������3+�A�D�0���\1iF@lg��3�n��@I�Ɗuk"�RU!8�!�������!�-�ӳ�kl�b��g�X�
��K�\�P2j�bF4Y�u;4X���լ���/Hh�����f=�YTHV�U�������om��u�㤗��:���n���ص�Џ$
U�y#Z�%�.N}�]���Jql��˹�f`vq��*Ke-8�QoA:yF���0dO.��N]��W��E�,�l���P��{n��5�N��㚩 GE�^���]q"�\�Qr��@�i64�BO`ŗaԣ�#;��h\;����+��n��)tF�����E�t�Z:�7<<�p�B�U���A���2��i�yճ@��l�'\pιp��=v*u��v��j�7n�WH��gA۷L�`�#(�gx��B��;G�+Un�X�{km����W�QzA�y�֮�A4ͪȆ����V]ج����-&gm���8���ݕ�'���9�ix)�^��e��gpfW����m�M`���@��.Uj�&�SpWN�S�"�a�6��Tl��v��V&�b� ����u�@��������
�d�1#�� ��f���{l6[K��%�%9����l3�3�T��J��sJ�jD��km�H[N ��!��6̴��[=�é�`�{ec�mݻI� �N�3������Ei)R���λB�ۆ�l���J�m��-�U��j�v�@|ga@]r"[s�jxش��8ۧ��yk�������z��v۰H	��۶ -���F����ڒ�Eqd�/
v�{dv��K�ӌ��J�ն1�N1�nyA�S���me�8ι�M!����vB�jS+;f���l�)%����z��6&�96�nvԫ�lug�BiW��-��(����T`t�:ó��:�`���=ش�k�]{n�iS�f�u�����<�7vm.e�P������=8h*y甆�
	�?":C�L@!���ݷ�͔��K��
���Q��\�]vQ�`.�o�n��:�y�<n��4�䇞Ԧ�N���v4�����]�mHf�����r�b��VL����`srY����y7b�	v��8��0.��F�vcM��-[�P�6�P�r`3s�͞!E�7k`[���b�v�n&�l�=��n:�	˱t)���Kخ�2�^��ٛ�\��#��ڳ��n�m	u<��w�kF���+�z6+�� ���nә����Ł�Հ��=�|��\X����20�F8`����ZVנwt��m���T����"r&�ZW��;�S@�����Z�Sqd�rF���@��M޻���ZW��>��ʜ�9$�䆁o]���ZoY�wt����fvwض���r�Gl-��ܥf�^�죓f]��.%SA�`k��Nz�<�H���3�=���@-�4�Jh���>�1*��<I�q�@-�9� ��N�诊 P��g:��9�>rھ��Б�ܸߑ4�I"�@��Ɓo]���ZoY�}�9+I���	�[�s@��V�[�h�)�rʭ�&Fē��hWj�z���4z�h,-�c�B4Ә���H����ǒ��.��4��R�<�.$�����*jULҰ�Ձ����w�{�0�f����k��h�FӖ[�=ݦ_{Б����Η���V�\LT��������-빠}_U������+����C"�����o$���Ӏy�Qv���v�,������u>V���ͦXz���	T'��M8��E�Uz��;V�[�h�h.,V$̘�0�S���+kQ��� `�村2�]��С�Hc�9���$��z��ZoY�{ӽ��5�vp]�6\lC%
�+�z��!#v{��˟M��-���Hmkݣ*�*����=�n���{8nb_b���|������N��A5L$�F��*�^��;V�^�hO�@q�C�C���{������O�6l��6�7zwJh�f��v����p�ffy=Bض��;ʄ
�ԏ��>����cc��v�N�Z7nt��\�����n��Y�K]��[O >߾��g�|��z{�4{ǎĠФRA'' ���_>Y���ؔ��~�p�ߎ w�f��g*��4%"��@��z��,��G>�3��>�4�M�5�I����Jh�f��}V��X�wvpS]�6\lC%E���u��>s�Xn��76�`_��������c�;�D�b)v�*������˫g�v
�j�˕n�M�60g��:��V�x�xأ�����9�<W���-�`� �,��{v��]��ޫ�vJ
�f�Azқ�B��>Y�C����V'[L�(4�%�ᇲ��{eZ�es�1܏i�ޢ.�p�Wz6�g�-�z�`�3ք<nՈ����,�o-�v��9뒐ul�=��{��{��?_� �Tt�L�9�F��nM��Y6�9"v(jY{z��ֶ�D�N1DG�y$�rP?~��@����ޟb_$����׀}��?�B�ж�e��u��g>�����{t���x��z���I�wl5ڭM[]��%UM��� ���b֨�\���z�Ƥ���
�7����<ٺ�
�W�wt�����x�J
E$�U��Ձޏz#��O�6� ol�<�����`��	E�F���nB�:�XAJ��lqF��!�n���Ɇe\��u����ޜ �}��1,��bIyߦ����?��c%�+bvY�=�]�ߣ�䁽u`fN�`4�����*eL�b|a�ٛ��	fl���bX�%����'�,K���ݱ9ı,O��w8�D�,K��xbr%�bX��~�K4��]��sw��K�Ȭ���~��,KĽ�����%�bX�O���,KĿw��Ȗ%�`�����i7d�ܻ��'"X�%�~���'�,K�����5<�bX�%�߿oȖ%�b}��lND�,K�<�Sw$���'��c�W�7V=M�wf7gl��oa;y2�zP]��Hp�~�߽�7���߷���Kı/�����%�bX�}��C��DȖ%�~�����%�f&,٪-��(��::�..��ı/�����%�bX�}��S�,Kľ���Ȗ%�`�����O��n&ı>�����[n��ٗ7x�D�,K����S�,Kľ���Ȗ8�� ��D�<����Kı/�����%�bX���e�\�]�̰ۛjr%�g� ��3����O"X�%����59ı,K����<�bX�'�nv��Kı<��v˞��7m���O"X�%��w�S�,K��(�=�����%�bX�����,Kľ��w��K�7�߾��w�ۡ����n������h1[�A�ܽ!��us�>��ү������is6jr%�bX�ϻ��yı,O���Ȗ%�b_~����*�ؙ�LY��..������h��eM]�K�����O"X�%���ݱ9�9"X�����<�bX�߷���Kı/�w���'� �Q7LLY�|?�h�ж�e���18�%������%�bX>�{59ı,K����<�bX�'�ov��Kı=�xgfl�.��n����'�,K?����~���bX�%���oȖ%�b}��lND�,
������(s�7���x�D�,K�|a�3p�f�ܻ.�٩Ȗ%�b_>�w��Kİ�������=�bX�%������%�bX>�{59ı,O~'C��T���q�xJ�فnc��2�k&�"grCEd2X���o0����)�e�'�,K����؜�bX�%�ﻼO"X�%��w�C�O"dK�?;�y�񉘙������M��mݱ9ı,K��wx�D�,K��f�"X�%�~���'�,K����؜����*n&ı>�g��.x3.�&��Ȗ%�`����"X�%�~���'�,�!�2'{����Kı>����O"X�%��w3s[ai��.f�ND�,�Q��3�~��O"X�%����9ı,Os�w8�D�,�T����59ı)��i�u¦���m�Ky�񉘙�����؜�bX��G�R������}ı,�o���Kı/�����%�bX�#��@H�
����}Ӹ��qV�gre�Nf�n�=Y�8u�m�mY�;�`�����{z
�^X�{tr�Dͥ�
��YեH���yY�I/+��a�5��%�6���í��mu����;v;"����;qV�W�­OP�sFZ.,4sQ�.�ˎq��Lyc�C�њ²�=nG�xBûb���h�s�n-�]OQ*l�m��n��i��f�m4�� i�.�d�a)��]��غvWٽn�Xݱ�U����+�X�|r�%���*����I�{���{��7������yı,{����bX�%���x��bdK��w�؜�bX�b�w�i)jl������b�bf&bp}��jr%�bX�ϻ��yı,O���Ȗ%�b_~����'���&,٪-��v��딸�bf&ab_{���<�bX�'�ov��Kı/�}��yı,{����bX�'����&����ə���%�bX�}���,Kľ��w��Kİ}��jr%�`~dL���oȖ#13���㍷k���Y��&bq,K��wx�D�,K��f�"X�%�|���'�,K����؜�bY�7��������� �V7V�mny�.v��vXt���6�;\F6���T�;�.�̹77x�D�,K��f�"X�%�|�{�O"X�%���ݰ?��L�bX�����yı,Jw��nkl-3Y��٩Ȗ%�b_;���z��@X�`A@�S��?��O"X��m�Ȗ%�b_����yı,{�����*�S"Y��iݱ¦�]N�#���13����9ı,K����<�bX����ND�,K���x�D�,Kܝ�����f�wm�ݱ9ı,K��wx�D�,K��f�"X�%�|�{�O"X����O߼���,S13�����e��[N[o1~11,K��f�"X�%��1�~��ObX�%����9ı,K��wx�LL��LŻ�S����SiҨE,���n�z��̽V�ݕ��Rh���PbC��,��E�+�,���d�����L��O߾���%�b}��lND�,K����Ȗ%�`�����Kı<�ޘ^�7-����n��<�bX�'�ov��?���M�bg�����%�bX=���Ȗ%�b^���Ȗ%�b{׮1�H��]���131v{��'�,K��;۩Ȗ4_	�3���A�������@�HA� �B�B�-"��0�� ��JI�'�b��T �"!0�hŊA=M����o��Cb��H����I<��Įk����B�� B+��<1��z ��b�血�ʔQ�	�~Dv�p h��br%��{�O"X�%���v��Kı<���<pܻ�]��'�,K?���~�߮�"X�%�~����<�bX�'�ov��Kı>ϻ��yı,J}�fnkl-3Y���S�,KĽ���'�,K��P?�����؞ı,K�?gȖ%�`�����K�f.�(�{Jɍ��$9PDʮ޹u�х0=��̊[�&��]S��#�Ll��sw��Kı>�{�'"X�%��}��Ȗ%�`������ș�L�����_�L��LY�5���*i.[��br%�bX�g��q<�bX����ND�,K���x�D�,S1{��f.�G���{��ZR��s6Y�����%�bX?g��S�,KĽ���'�,K����؜�bX�'s��8�D�,K���m�m7B���\18�CRBV�W{�y��2�D�o�S�3*dLʝ߻��{�L��CP|W�?	�?(���*s �ＳS�3*dLʞ�s���ܶ��%����ڙ2�D�7�r�"fTș�;�w���ڙ2�A�{�592�D̩����'��ș�2'���zߞ��{�^x���C<�e�����F�n�C�u�f�V�5m˳�s�?���F�b�s#�ǋ��1H�}w�1y��S*d���S�3*dLʙ�����ڙ2�D�7�r�"fTș�<���=����ws��2&eL����jr���M��S?~��x��S"fTȝ���*r&eL��S���8��S"fTȘgݙ�����f��٩ș�2&eL�{��{�L��S"}�ݹS�3+��T�kŷwg1y��R<PYۼe��{��;ܧ������Ŧ�-q=��D̿�$����S�3*dT��ݜ��1H�Ag��e���ߒX�ǋ�}�ט���)(,p������ҙhOw�ܧ���=ߗ�{�O}��3*d?���jy2�1H�n��9��(b��/e�q��2�D̩�A�$QP=��n�ס�Ln�+ ř"�nݠ�R�,�p�hƣt��lc�e`(j �2Ɂ��1;U�O��Ia��!�n�痋et�e����x�1�O��h�)�;;,��m�\MŨ�"ëSm�vE��Ī��e��)6UK�J��`zч�ꨍ�µ.��ѳkۛ)PŬ�����k9�Iu:tz.!��涚�2Б-�IZ �<n�d�:�GӸMs��=��������g�ZѪ�+jK,���R<PY�s�qp�%L��S�O}��3*dO�{�(O"n�ș�?o�߳��2&eL��t{�6z�!���or��{��~~w��'��ș�2'ٽە92�D̩��{�O}��3*d��I�ȟ��NsS�3*w�?�/��rܦ��r��'��ș�2'���S�3*dLʙ����{�L��S ��rMND̩�3..���9��(b��'��s�8R��v�ND̩��v������=��D̩�{���S�3*dLʝ�|��{�L��S"}�ݹS�3*dLʞ|���'%��)m���1H�Ag��$��Lʙ2��=���Ӊ��2&eL����r�"fTș�>�����ڎ�)�w���?+H/i�mI�F�i���cG��9�q����f�`�6�\�\����4�I��jr&eL��S�O}��3*dO�{�*r&eL��S���8��S"fT�?w��S�3*dLʟ+ӳ���K*v�ܧ1y��R<P����ʜ�;�
��������ș�<�߿g�jdLʙ���592�D̩�{�g�jdL��wxw�~]��A�S-	��{��dLʟo{��{�L��S ��rMND̯�!�7jw��?N'��ș�2'[�	��{��;ܧ�����5kF�X�f���jdLʙ��jr&eL��S����'��ș�2'ٽە92�@�($ݩ�~��8��S"fT�?�]��g��ڂk���)�w�Ow���2&eL��ov�ND̩�3*}��s��2&eL��y�592�or�������ߐ�tS��Fa�tvJ՜��۲����%�)�{��qg+���N�wv\˛8��S"fTȟf�nT�Lʙ2����8��S"fT�?w��C�ț�2&eN������ڙı/���.p��ݛn9wr'"X�%��w��'�,K����Ȗ%�b}���Kı>ϻ��? ��0��^nk�s�2[e,R�9�񉘙�����59ı,O��vq<�bX�'��w"r%�bX�g{��yı,O���75������S�,K?(�"w���8�D�,K���Ȝ�bX�'���8�D�,������\1313T�f�,��[r�O"X�%��}�Ȝ�bX�'���8�D�,K߻�S�,K�����Kı?*��%�ۦ\�r\�rf�i�ۍ6� �	"gF;�90vӲ���&/󻕛���I��曙ff�D�%�bX������yı,~�ND�,K���'�,K��>��ND�,Jb���.�R2�䭩,�������~�NC�
�"dK���Ӊ�Kı>��܉Ȗ%�b{��s��O�fdx���7lr��ܔvJ�.D�,K���Ӊ�Kı=ϻ��,��Dȟg�߳��Kİ~��\\1313�+��F�e36q<�bX�'��w"r%�bX��{��yı,~�ND�,,��uD����O��=�O"X���]�lc�RIKG �l1p��LK���q<�bX��@��xjyı,N��?N'�,K��>��NLL��L����{誖IB�v�m-����nڶ(s�0+h9�6�ɍ�k�1�kvm��i����%�bX>����bX�'�w��O"X�%��}��ʯ��؛ı;����Ȗ%�b~3����m�S4�	sMND�,K���'�,K��>��ND�,K���q<�bX��w��"A `�'V�����Hۗ�/_v�b�'�}�� �'�>����bX�'���9�񉘙����ڈ���U�s7r'"X�%��{�8�D�,K߻�S�,K�����K���"���\1313���m)�-�Lۛ��%�bX>����bX�'�w��O"X�%��}�Ȝ�bX�'�w�q<�bX�'�����2��
�\�)�3*�[��r]�^�K�v��ˍq���ۋ�j�㘆MZ`���۬u�]c��a�%�7ak����Lض헳�ڞzH`Gsi���3��҆_kgdűp���l�Xh��R[R�^�sɵ��t���K�;Wz�=UД�rË@Vi�L򴰇�'�d�s᳘�����,�Pl��:�[	�����:sw�/n��GI�7f�n��q�͏+�;y�[q�:q��n�<��sڿ��v�����M�˛���5=�bX�'~��Ӊ�Kı=ϻ��,K��>�s��Kİ}��59ı,O};̳��ٖ���L����%�bX���܉Ȗ%�b{�w���%�bX>����bX�'�w��O"~Eʙ���r�5G\C����131{;�9��,K������K�a�2'���Ӊ�Kı>��܉Ȗ%�by�����L���)���O"X�~@C���{���S�,K����N'�,K��>��ND�,K����'�,K��ϻ3s[e�ݒa.i�Ȗ%�b{�y���%�bX���܉Ȗ%�b{�w���%�bX>����b]�7���1��A��SZ��Rg�N"6g�&���j���Uv��}t�
�}��|���ٛ��inl�=�bX�'��ۑ9ı,Os��8�D�,K߻�S�,K�����Kİo�v�I��M7f[���9ı,Os��8�C�h���,����bX�'���Ӊ�Kı=ϻ��,K���ye)����,�������~�ND�,K߻��'�,�"}����,K��;��q<�bX�{�v\٤���wI��jr%�g�O�
�����O"X�%������,K��>�s��Kİ}��59ı,O=��Y���3)�������Kı=ϻ��,K��@�P+�~���'�,K������bX�'����<�bX�'{){��ۛI�����]:���f7!�϶i9Pj����Q�X��]^d�"�û�w��oq��O���8�D�,K߻�S�,K�����'�,K��>��ND�,K�_�d�6fnn�L���yı,~�NC�+��,O�o�׉�Kı>��܉Ȗ%�b}�w���%�bX��r�kl���L%�59ı,O{���yı,Os��D�K	���A�"� 
�'�?������Kİ���jr%�bX�T���Z:�,�ʉ+�/�&bf&'��w"r%�bX�g��q<�bX��w��"X�%��w��O"X�%�?C��F"�괍�l1p��L��>ϻ��yı,?�O��zj{ı,N�o���yı,Os��D���L��]��}��ƭ��˄)er�}{����6���bKj�ɜժ�p�V�BY��3ss��Kİ}��59ı,O{���yı,Os��@��<��&bf.���b�bf&bb�ڦ�R�n��͗34��Kı=�����?��L�b}����,K��w���yı,~�ND���S"X�}'�G��H����|����L��^��9ı,O���8�D���D�?w�ND�,K�����yı,N�1��!]��bቘ�����w���%�bX>����bX�'����<�bX�*AP� sȝ��a��&bf&b�7��P%��XK��O"X�%����Ȗ%�bw��oȖ%�b{�wr'"X�%���������L��^��ô����lI̻no\YN R�IC%�sr:��1��=*���eLm�JC�\\1313}���yı,Os��D�Kı;�w����ؙİ~����bX�'sM�Gc���$������������9ı,N���q<�bX��w��"X�%�߷��O"~ʙ�C^��#��7%���13��;��q<�bX��w��"X�%�߷��O"X�%��}�Ȝ�bX�b��]���#��),������	d���S�,K�������%�bX���ܩȖ%��ȟ��߳��K���v����%�H��Uqp��N%�߷��'�,K��>��ND�,K��{�O"X�%����Ȗ%�bhj�C�*����(�
���!����hJ�B+��5Z��՝y���,�1���Q<b�(���B�#�b� $����@4F�_U�Y��*AB�Y�(X�\���3͓wvۻ���!� q����m*Kv��%@��%�ہդ ��|jٜb�O%3�V
ZU���5�k��کV�nS1�\L���D�V�ٵΚh7g�j�D�˩�s�����vĦ�#-ٙ��nN'�j��<��6��.�V��x�;���>�ׄV!+Bvۭ6�j���xm�إ�κ�FG���8�r<dJ��� -<��jÇ��4�g���n��ɹu�4\�/��NѤ����:��f���K<qۭy�sNs�v��O�y�lJ`�,��Q�<�R�Pٱ=sy84��I��$�,�B�\�i5�m�L[��A�-�wY;]6ݍWR��n�����n9�c����s��\��!�RU8�3AE�Uy�K��Nm�z��L����<a�x!�[Q���@y㳩�j[�:�`�&��2ʰm �]��a�- Yj����^z����'��� M�8A�'3J8(2٬�';v'l�q<�p�e��n6\�>j㕸������[����n�	�q��St��A���!Z7���U�O0��:�W�F�y��rv�\.���Q���! 4W��<t�Z��k"�d%V��*�V��kn�v�h ����⋩�h�H9�;F���y��`�6�Z�F�i�,jBـ�v�e@�H[@ -��B�+6�eZ��e9����j��µn�N��`J�� ���稂w6s��)��� �M��f�v�ޠ[ԒFEV�Tdv�=5):xm��m�F�r=���u��F���9��ݒ-$�8hE�R�ԫ!��/֧\��] �YS;��[Բ�U\��7'
=�^%ܧ��0ʜ���]��A��yg ��q��8�&��ל�S`؀�xp[$���-Uq�7I�UTU*�_mu.Y��J�[7n5Q�H�[��Y��Ob�Z��@Q����u@�p�6 �`&۱T�F�]%E�xN�3�������|�� �O��8�P�U5U�Q��C�������S�Ps���n���7&nA3ZU��anܤY�t��j:u�N������u�(l5�\��u��a����#��˪1�6ɴ��mlcn�q��Cv�a�b����c6�U���q������qke�<���;+ΰkg\��uX8&Pno#�*��3t�*�ݧT�I�tΖóY�:zx�ꃴb�Zq�mjg�<�q.�c�TT��K���x�;Un��w���n�����_��o794�]x���.cv��ڰq�r��$�/X�U��&��^�KeݼO�X�%��w;�9ı,N��q<�bX��w���'�2#13��g1~1313�lc��{$�	sr�"X�%�����'�,K������Kı;����yı,Os��T�OS"X���~�͛$��͛d���'�,K����jr%�bX��{��yı,Os��T�Kı;�}��yı,O���w4����l�]٩Ȗ%��	"~߿~�'�,K��;���"X�%�����Ȗ%����?w���"X�%��~�^�d+��)-����������w*r%�bX��w�q=�bX����S�,K��{�s��Kı?b�=�D����������ob-�e2��砯k��b0���{�-��vҗ.[���=�bX�'�w��q<�bX���n�"X�%������{"S1{;6<\1313�����7d���˻�O"X�%��}۩�x�|FE�*|
���q�<�b~�?}�O"X�%����ʜ�bX�'s߻�����fG���v����2�ث�6�r%�bX�����'�,K��>��ND�,K����'�,K��>���Kı>�N�gsK�)�n�n��Ȗ%�b{�gr�"X�%�����Ȗ%�`��v�r%�`~ �����_�L��LŹ���!]�%�Ȝ�bX�'s��8�D�,K���S�,K����oȖ%�b{�wr'"X�%��������l)��Wm� Ɖ�.GN�A��c�+gjI3�29.rlnx��=��V�Z�4��Z~����D�{����"X�%�߷��'�,K��>���y"X�'�����yı,N���w4����l�nm��Kı;�����%�bX���܉Ȗ%�bw=�s��Kİ}ϻu9ı,Os����]�2m�f˛���Kı=ϻ��,K��{��Ȗ>!  ��"�"�F0�����>�ݺ��bX�'����+񉘙������h,��#r[9ı,N��q<�bX��of�"X�%��~�gȖ%�������L��Lž��6R��� �v�Ȗ%�`���jr%�bX���vq<�bX�'��w"r%�bX��~�q<�bX�'~�\��ݹ�-ܺl��h�A=q����gnư��H�9����[����Lۛ����ݚ��bX�'~߻x�D�,K����9ı,N��q<�bX��of�"X�%���t�v�M2f������%�bX���܉Ȗ%�bw=�s��Kİ}�{59ı,N��w8�D�,K�ۖ\�K���nR]܉Ȗ%�b^���Ȗ%�`���jr%�� �Dȟ����'�,K��;�r'"X�%�ߙއ�+d�JU$���13y��S�,K��{�s��Kı=ϻ��,K"�Q��3�w��yı,O���w4����l�]٩Ȗ%�bw=����%�bX���܉Ȗ%�b^��w��Kİ}��59�31uyD��+&6����FIS"#[z�)֗F��=��H��&ˎ��Cњs���sm�f����yı,Os��D�Kı/}����%�bX>����bX�'s߻�O"X�%�{;�wf��˦f[���9ı,K�~��<��QH�L�`���59ı,O��gȖ%�b{�wr'"~P��,O�w�6R��u� �v�b�bf&bb�{���"X�%��w��'�,*C"dO���"r%�bX�����'�,K���˟̱s5p�׻��7���x@��?}�?N'�,K��;�r'"X�%�����Ȗ%�`��xjr%�bX�{'Ngn�fR�͓wwgȖ%�b{�wr'"X�%��#�~���{ı,����"X�%�����Ȗ%�bp ����.nJeAT �� �K�W����{F�ظ��P�
S������a�C���z�O����{'V��+��'g�v���6�d9�Α��˨n2����RW�J�lN��n&B�&�n^;F�c��,�f�|�v�1���ڥUgg�4�] n�F�ӗ?��~�\�j�d;Xyv�t;+9�t݄^��=�疧+�f�t��q������*�6c�v�d�a�I��+��}�O]��m;� ��7YŸ�0um�c{;ș���F�m1~1313���a�Kİ}��59ı,N�w8�D�,K��wbr%�bX��������7I���O"X�%����Ȗ%�bw>����%�bX�߻��,K��{��Ȗ%�b|g�˹��sm�	sMND�,K����'�,Kľ��؜�bX�'s��8�D�,K߻�S�,K���3��v��m�6fn�Ȗ%�b_~��ND�,K��{�O"X�%����Ȗ%�bw>����%�bX7���vm���˙�37v'"X�%�����'�,K�� }���D�,K�w����Kı/�wv'"X�%��{'s�ᖆv&����-�SɎ�z���\c=�\JN�i����w)O���Kİ}��59ı,N��w8�D�,K��wbr%�bX��{��y=���n�����X����V����bX�'~߻x�C�� �*��D�,K�n��Kı?g߿gȖ%�`��xjr%�bX�{'NN��9%-�1~1313����,K��{��Ȗ%�`��xjr%�bX��~��yı,N�nY�Z�8�-�.��������s"X�%����Ȗ%�`w����h���r7	������h�U�{��*��@�.%lC\<��; ��Z^�[Ŏ�v@Ӎ�nax��صn�W��]���u�6(�=��ߟ��V�}�@��z�빠r�a2*S4���U�k��H�Ϧ��}q�[ҚV���$I��rM��w9$�߻Ó���^������h���/�Ǖ�cYE1���>�]�ޔ���h^�@�َ�ɊG"�	�3@��4�u�W��>�]���,BpxƜ�1H���tvK��ۮPv�A=
�\Z��4��Wg�"&&&�䆀}�@��z�빠z�M��u�ō��M<�@խ��$f���Xٳ]�$n��rr,r`��@�~���z�M ��f�˭zb��HN!c�9��?wy� ��ݜ��{8	bIfw1��Q47���I>�N���6��&9�p�>^��]k�>�]�����5,O�P�mQ�89r�*vQȐ��������E�wU��cm�rF��&/���|P�RD�lnG�?/����>��[)�|����O+�Ƃ(�f7z�:Ձ��,�k�V�7������SnE�-�~����@�ֽ�>�@���uDE�p27���խ́�N�a���ou�`z�?�����ڐ`�z.��y�Z���>^��ˇ%�#�����j��b��9���zq�tx��{	zwGom�ð��yݹ���l]��s��c�$�KZ1�66d�)cpɵ�d[������]�D�3���ض�^^y$��1fx�d�&�j˓��'���o[�o����N$�KW��^Gl(��{r�n;SЫp)66xm׍��v�;\٧�u��b�L�gr1��uƮ���O{���w��>��}���sU=�2�=�u�%�'g;��쥉3uu���p��+��X��UN�/����,�k���DFy^�����G��-��"���ڴ����Z�����;��@��Q%|��������>Y��K3��oπw��πu����h�ei���˭z�}V���Z��^����p�0�������U�|���bY��s~~���N�����~=�c�:苶�<ӂ��r�������4kiո�lɺv#�C�ݓevl�J��:Ձ����Ս́�-�0nv�S-���so$��{��<x�X�E=O�P=Q0x�bW1j�K1�u��g �gu�;=��ر,l��&�ejA�� Ig �����ڳ�����|�[�6�4>Q2Zյ7-�K�Y�����>�M��X�����5ĝ$������h���<�k�9zנ{�ա������:��X�螁8�ۙ���⵽j��n��]]>�v�x�����~�~u�	���9w��@��^��;V���� �Τ�C!I����́�-��V,no��H|�&:��������8����<����O��H��R �c>C��Q�������V�,Ȅ&cp�#4*��2З�x)F(|x�j�O_����&s�c�'=��-	��4��e(R�"�y00`A@)$�1��N2�7�����.��@`!��ؔ"@�A�!B%l�q��!g��z
g�(t0>S�Aj���P�'AA��xu>Q�@�x���|��_����'U��[1Ѹ�8�$pR8�W�X���5=sa��DBݮ�`=��Q�ĞE"�<�k�9^�@�����{��>�X�獵�����\qԂ��,m ������oA=�3�5�;)�m]�j�+FG&�܃��
�_�@��������{���5ot�|�!]��TI�9��;V���z��z+���Q+��
E1��$Z+��X��ޏDBMs�7g�X��.J�T�EUJ��p>Y�b~�wg ����y;��&n'�1/�y����f������J����p�ff{������z��Z�ؕ԰Y#ALqF���xH�@2*�O-�"2*���#n�p�V��=7X0ɒ�ԏ�;���@����v����[1Ѹ�8�"�RH������Ė3Œ����5��N瓽|�g}VB��X��8����9^�@���@�z�݀�:��
Bё��%�bO�{��{��|��k�=�j�>��T-�!ȡ&<NG�fKj��{�~v{����6�"/  +��9���=�e�,���HIs�Jb�`�;It��i�u���>K�1w\G�)u�N��y)m�b`��k��M��A�%��E�x$k��tA�v����q��v��]�I])�4������lcD�Kg��T*�WA���J�
���S����^�m��:g�+�ӱ3���j�yX�s�u��cb�],?�\O��!<^�eʇ"�M�z�:2V�;���v".���9�͒ۻ7%�L��f�Q��/E�\m[���6���n1ѷl���p]y
H�Ǆ�p�z��Z+���fb����gu�_u����8�UJ���yڴW��=��h�W�k�8d�m	��W��=��i�,���������=}���UD+D�1�#�=�j�:���=�j�9^�@���'�H�6��:���ވ��7k�|\�l�mXd��ô���������ge��P@+nʱuuU�w]Yޢkw�t錏C�������~+���hzS@�`;���3.if\��'׿w9�%=� �����V�,�mX��Ю(D�(��Jj��̖Ձ��=	n�r�9~�����IY����ذ�-�z#О��`n�r�1=s`fKj�͒��&	�2c��h�h�W�{�ՠu��r�X0X�&$��+iG�w[���gϷ][��ى��d�����rÎP��-�H9+�^��瓽|���|���=�n���ql��� �mH�yڴ��h�h.���,K=ݪi%i��Z@�W�:�ݜ�'z�w/ر|��$���z��8���w�����7`�z�1n�r�1wt��ڰ5n��7H%�r���J���~}�g �f%�u�����<�w��|����[X��ʭAˋ�ж3�{^���k��/^�;��vy�;��,'�B�9I1br?���-�uz��Z�h�Q+0����`5���{�	�ܬ��Vd�VV�\$�d���yڴ�j�=�j�*�@:�*pFԑ6�%|�}�O�Ͼ|����~���� �z4D*��W�0T�nU�|���̀�XH3����>����{����͞�`<�Հ�[.����k��S�'����$�lv��2��1�;�u��c��[���?}s�X�Ƶnyh�m�7�`}�ڰKj�̝j�x�M��n&�H���Z�j�=��h[^��0wqdbbs������<����,�R|����=����=��[d��&&9��;V�U��yڴ_U�r=�52���UR�z���{ѻ]����3%��"�S�	��I���[�urN0�J5B��م���wMg�$�&��z4&F�:�7kCc�a�ƺ'sQ#ui���<vm��+��dYտߧ���'n�����˧rv6�u'@��n�۠lk�S��pn�V%�9-���z�ۚ1��v����I7HN[)/8Ы,n�Q��;�d2X��\e�̔G���g�(�Qsv�g�Rl�N�թ 睃�!T����lۅ��L7$���<Vqל�B��s�{jd���v��Fi���a �&8Ԏ���>�@��^��;V��z� �̩�aRD�I��X���"=	�ܬ\�l�mX�'�L�ѓ$k����=�j�<��@���@�ֽ��tn,S�C&F�X�s`fKj�խ͇{��k�X��~sh�D�G��;V�˺��v��ֽ ������<o��E`�^rSƗ{^Ӎ���gl�̼{&(9�lރ���GF&718�.����Z�����f�r�������U!5U6d�W���Ȋ���k�&��;�@��^���T��,$sH#�@�ۛ�՟��$��v_+v@~è�R"�c�p>Ib~{w_ ��vh��+��ZʜD�i7��ֽ�}V��z��;V��{??+����ڳ4�F�5��Յ5�f��l	�$�*n�����E��t�}]vv�Z_�G�w;�h���>�}� �j�zَ�Ŋd!��h��~{���ۛ2u��$n�T�ʡ(&��,�{7_ ����bȒ1$�!A_�:	���9y$����$�{	�qd����ֽ�}V�����}��,�d�����=���|�e���	���3'Z�?{:�/�͞�`j�s�U��18L��H<1)xHs��X�N̮򅸍��t�k\�g��ɚ���4qhW�hyڴ^��y�Zy��e�Ad�LQ��������u���-��� ����6�6�qh���������ZW�L�<&(E�ԑ�~���ﷺ��;��~�w����Kx�3��K��4�o&�pwj�IZw�,x܋@�^�@��ՠr�W�{�޾���]�r�BISI�hۘ�vK�]s���!��g+�!^-q�L=��r�*�jIAUS`}�ڰ5f��3'Z��G�3�u��"j{+�܈�#��_��p/uz�����Z���`�q�j�B���1f��>rڳ��y,��VV�z��F�Aa#�ز'�����v��uz�uzy��e�Ad�LPN��Z.��.��'���rI�Q���7�@4����*D:�W�LS$�£$ ��@�V%����K�O��z���4@�U�)P�ZT�(p >*�Ȭڤ�⡱yH�V#4�"R��D���A�cBT���t��;���o�׻ۻ���p�l$�#e��f�U-�쎓T��$C�t��Aem\�H	�؜lm6����ZN�2δ;qR�*ܦn.&�n0$X�El��t��1���%V��*�먻�a���ٮy��q��M�ղ�푦C�ݨ����<�3��`�5k2�8neNM����Dn�3�u��u���kpR1��M�Zq�6�g��	���&�-���}�(]��F�g��n�-�1�`��F�kN��U���eG�F�<t筶�.q۞{p׶�;����˗R���}�mkOL0�=\u�n�ؓmĸyF��uڱ��籺#h���.t��O��G*�&����a�f�qkAnN�� �Z�9_A��Mo�-}Ԩ6�Ĭ=��OWU�83�vH���4�n�lq�T����4V44��yGj���y0��{s�0A�eX
�H�/bSl�!��j���zSh��Aj�d<�lD�m����$��F^��:mP놓GYNI�N���F7[yr�&K1�'��Q��r��X�snHɵl��\�&3�x��j�rյ�vs��VMT8���ByS����A;�����Hv�JUA�jx�e�v�]���X
q����Ҡn����[@�����:̙	6�F6W�j��]���8ێ�b�!�ֹ��@m@E�)�kn�:A�� $-�$ mHv���ȹj��9J���T�k�;����ۮ�"Ap[�Qmml9xβ�٦��r�/Zm[�;m��G �z�'%.z�����X�m׫g):f�-6�)�v�qCm6C��-�@T��[Ae�� m�KE�km���n�ml��gl@�J���U.1�ݮ{Ku��a�<�[B���=^v]_[�*��+W��z�����R�.��P mT��Z�:H��1��N�ULj�J�ȴ`z�Sɒ��Y1�K���u�ӝ����s�*���p�q�\�b����ge�Nv���3-߁_�u ��!>�1�b�ȁ��	�� ��b)Ꭓ�ә�7$�6�ɹ�wb�����Il3�����dZ�۰�e'kq�n�\��(�ol��ڳ���eK���%ĺ�����c����ݶTvطG\ ���6xi���l�p��^�d�=��[��[(9�k���5��Y�z�9�Hn�3
��)�8͗.^!��U��������6�]i$�N��w3���&Й�+wB�l�0�P�=7���w���7c���r��p�HqcF{l�甗tKe�"s����t�EI1����};�Y17J4����������^��YM�v���L�<"�G�ԑ��\��#�������=��պ��G��I��ڦ�V�b�֢v��<}ݜ�՟��DBZ��5>�>�u)5	�H���=�ՠr�@��g�I?&���&����Ȋ�TҰ5n��?G�/�~>�6[_m������kf�l��T3�-�n���gnsէ�e7,�q�5�z|Ɋ�t�X�G��mz��zs�h���gu���cb�z˺����?b	�@a�� ,������v�~�@�^��`%�r(�I�����j�>]��W��>]���eR*��F�nJ�$��X�X��w��:�߿�@��U�w��@���ɓ	��5$z�����Zyڴ�uz��ey�,����C��d�#�[]�/N�Ǎ�;a���r�.ʜ�\i�y����Q7,�����|������jY�bK�^�g ����\N*����|�Ձ��s`bz���gZ�Б��zJ�,mJ�9_ ��vp}���ą�@ �Dz��,TJU
%G��G�v�g$��}��'�������ji�gs�K3)���8U��zyڴ��zԷ��Rd�ET���\���C��_�{���z� ����ld�1Ǌ5!yq�ng���n�s��n-3��t�]mӠG��������L܊%"Ja������>^���h^���2�� N�&�>X���Hݞ�`j��`fKj���h�dƂA��G��;V��ىbM���|�gu�;ڧG(�L��$����I�=ݜ�f��y=���� �.��~|��o��'����;�e�a%��'z��������ܬ�76��9��SH@�YT��.���g �n#�e�ݵ-b m��dHFa&(���6���Š{Ϫ�=�j�>^���h{8U��Md�$�qh�hyڴyڴy�\�X���Q��-�k�{�K2[Vd�Vc�X$�R��IL$r��Z���޲�ץ4�2�� N�&��;ε`tG�7z���\X�ڰ.=���T�Ӿۏ��Xm��t�m�2�	D�*02���	L�^��91Ѷ����v�4�Vg�����(y~p��b�Y�H���h��ظ��m�ٍ��]`����c���k'��NOG'<⎹�nщ7S�� �`�b�ٰ��t ��젛�s�k�G&���rG �ɛ�Y�`VKYm��b똓 2�P�W��V�.ܴ.n�Y���fl�7p��p�8	_;�����wR������׶����듌ns��۝�=m�¨-׋�SM�NՎ�T�/�o��\X��`fKj�ܖՁ��tN�#$�`ӆ������3?�;��Xg�X��`f�UL�&���'��;V��v�޲����qWdMa0"qh�j�=�L�1εa����v�����K�JTH�I����YM��z��Z˺��w�!`�F6Lj2DQ��k��{jUu�l�Ru��n4�cN�8�+sȸ�C@�zנ{�ՠy{��=�)�|�K�W"iI�Lq���;V� ?�� �P����Nd����p���4��z�u�Dx��Jf���5́��~��%�{��ݞ��<�e*�-"�#��ى,~����ս�`fKj�ṓ��KW�țx$�yzנ{�ՠyzנ{�ՠ}�\U�I���ǉ���\\S�����]J��Իq�.wI�[�#�����J�&	��2[V,nl�m~���ĳ<��߾�tD�?�iWm��]���2[V,nl�mXF�ضd�$����h^��3�?����"+X�'WD���+n{��ú�a˙UD���U#-���Y�������=�n����v����7r&��SjG�{��`j�����q`bz��4Bn��>�<��α&.��}�����r�m�n�`�������p�O��������k]�����l�w,nl�[V=��0xH<�����=��<�k�>�h^��[1�I�?���0RC@�%�`}�ڳ���D%�{���uŁ���,rGd�-��1���|�����'������"$ ��**{�
p�o��rI�Й��6��m�ͳJ�ṓ���76�-�����<w���8碵�{Q��#��ݘ=[��E��cb�����;���=��z{fq��$n(�I����=�v��;V���^���]mI#�)"�E#�<�k�=�j�<�k�<�k�<�\�v	����&��+2[V-nl��BZ��t��~4�u' ��)0����]k�<�k�=_U�{�ՠu�¸L#�j8�/Z�u��=�m���{��xb��<���4�vnni�ɚ�����O]��;Y\���n�<�v%��f捈�y�iJL��)|v�N���qٶ������۴o�М�v0[v.C���km�5s����Ș��Y玱�]vQ��f�v��0��^G�UVۏl��Q$����wj��ƥln��,��T[y���ko`�5�lX�]�}8t�7�a���ϩI�������������ݹ��m��6sh����!�rOM�d�{�p'�l`��\��
y�(�Y%V��g�x����<�w��z���^���:�8�mF�<$�@̖��"=�z!!��V�M����䇤кiz�T�R�Ұ5ot��נyzנ{�ՠ{�V'���7n�8%�bO�����{��y��_s����=z�l��b������'Z�?F�w/�Ž�`b����q�B��ܯk<u��u�jV�ܲiwny�8�؎�M���ڹЃVТ��4���� ��s�>]��ޜh��=�.�7%���'���8���H!2
:	wg���9$�ﷳ�O}�ՠ}z0����/棏@���@�t���;V���^���I$�=�Қ��Z˭z��z���6��Hp�=�j�:2w�~V�M����x��t�fWW��
��]�"��ѶAyuj����vM�\y����x��"��qh.��^����h�hvp��C�h����1f��1f��>�mX,no�=z�l�[Z������{t�{�����C�P��E���p�\1��1��d��-�� ��P��V�R"��T)�&^4 ����!��	-��1�D#�" B1#1D�R D�`B��� y��`c��*�H�� #��D		&���+�Lb�����T/PՄ}H���� W����T$H;�b�	�:b�.$�+geX1&$�3�4��!�0��<M=�U�1�<����:�B��{��E��%u��('�C�N)�@�>g�=;���'o��rC�z��N���aS���%��n����lY�lX����)�I	UD�rW�<~w��|��g���_���}�j�9l���(��#�I$pۉ�7;:�C���m��4��t�s"��v�]�L�"�j8�/uz��Z�v��ֽ�f:7�F�"����X�ڰ1cs`b���G��=����C�X���B(�|��|����p/Z�{�4񃸕�A�Hډ:V��76f�,3���=�<1HD �dT �`Ե���Ǟ+=���{գ��d���iX���?DG�z����Vd�V�w�����j�t� s[��99n��iؗ�َ*m��g��4�t��N���jNA+��z޲���Z����ֽ�yV�wK"�cjHh�o���č�|�[�6�����$�����@��U�yzנ}�)�{�ՠ}la\&	G�&�Z������8���p>Kس�y�>߾�|7��8�=�YM�ֽ�~�����1bϱ1-�[��*r��Z�2�N&�n�W�����Fp�]�R�C�1o�,l�X{f��F�q� �^��ظ�Tf	���[b��.�s����5��n�,�۷6�F�#�8�ݒ�l\���nѥw`�%t�C�\]����n�:kn����)*���v����:�+!u.%�/��h,0�v{�,���_i�q�Dk,�m����gj\ь�6�&i+�W��9�6ˆ��i{���hٹ7\;ۯF�;fj�w�Z���+��5$�s&<M����=��h^��z�h��V��D�`fN��Dy#V��7����cs`}��U�`�$l�"�<���w]�?��ot���3dn�fUQJ�*��U6����2u�ޅ�����r��o�(�E�Ԑ�>^����/uz�v� ��+dbicsC��qsR�k�gN�N�ê�b�n�h�Š'H�D�m<��Eg����?�y{��>W��>^��^�+��LWp���y$���s� hOPH������{}ތ��y�`4�M��:Ձ��tn(̍���$��+��/Z���/uz��<�Ƅ�r�����zy�Z����z��`�%a��H�)��}V���9���������z�q+`�H��ݕ�QL���^ڊ�n��ۍt���CK��]]���	<R	��<���<���+��/Z���s-��$Y"&8����=s`|���7'Z�1f���G���m���(E1�$z�~�����5����	C���g ���g =�gD�0NlmǠw�U�y{��>W��>^��^�,����`ܥ`b�s`w�y��-�ru����~=�C�]5��3(Zʝ;�[&��ܙƉ�a�,c��p�����e��+Q�z��z�ֽ�����^�|;�*q�m��ǃq�/Z���X��'�o� ��������R
G�^w��<���+��/Z�����	��<���<�k�>���'��w9'���Ng|���I�ý�Ke��]uJ��g�|�K>]�o��7�~|��{8��\��hqB�΋
�'�N3m�N��+��7���[-rj�=md����m�1C#�L�-��zy�Z/Z����:'��q����}V��ֽ�����g71��큶�(�H�h���:��z��Z������c�qFdjI�qǠ}_U�y^�@�>�C���{�8�MQk�H�,�E��x޹�?z2w�~��2u����G��������!�ߖl���Yڥd�f��]9Ϭ���]�6v��۞��74�`ټ�{�A�v坶8�p�9�J�5�V��c֖K)����oR����ߍ���#!g���ڽs�c��m��6�dN������pA0����d� ,��IΨ��	��ؓ`���V7�hU��9��2s��ے0���EWR�u�M�Y7M��2�n̗h �W����o��?T6حeRc,l�u�t�/��c"�����L�s��x�:i9��B��@kw��Ս́�:����G�5s�z��f�&#���z/Z��֬O\�,no�	��S3UU1k�:��gu�}���Y�$��w��@��~z�˛m�P��7�����́��3i��d������ӏ@�zנ�+�ߟ�w;�hW��/��+�`���ic��}��&#y�u�blv݉��Wv��S������6I�<&FD����
���{�)�x��g�$�~a��vp��4��U$������I=����q�Tv ���ȏ\G�"�%}�lM��5f��3"n<+�5�Q�X����^����O�X����8����=�D�o�W	K$��>^������Jh+��w`%qlI�#p�I���^��>�@�^�@�zנv{r���.��(I�`�'S�2�g�Uj[T<ШwN��ݤ?���7s^��$R)1E#��-�z���^���^��r��w1L�`��h+��/Z�^��/uz�����)D�q�/Z���������x���-�����_���}z0�L1�22%�����k��6�'{��}��q)mI�Ǡy{��<�W�|�k�9zנ}�\U�I�ȘLCV��'��=8�t���m4����q��V�����n�熸�X�ł��/���>^���k�<�����,�Äm�q�,no�����$5��`j��`bz�@��+���(I�ȴ^��'�l�DD%��M��_+V×2�*�R�:���I/�b���~����rI����I� ���� ��{����x��6��P�2)��E�y^�@�zנr��@��U�*1u�@����2A..��=���-���ڭ��s�O@�p�q=��bNliǠw�U�r��@���gرg��������څH�X7"�9{��>W��>W��;Ϫ�:َ����5����+��+����h���\wT��n�����bJ{~ߧ ����_��p>I�7�8}5=���Im�e�ru��=�_N��-nl�ȈEQ_�������"��� "��TE�U��TW��ATW��P��TV������ATW��TW�@EQ_�TV�
���"��� ����*����+� "��� ����*��*���b��L����Yn��� � ���fO� ��>    4             ( C� T� H���P JU"� P !J%    P *�
P)T
 � �     J(� ��s�y�qz�1���-���8�;��ng�g�}�׋�;��B�q�nM��v| n{�{w�A� �/^Z�o��ǸV}�C� �|�,��-ۏwh�   <   �!@�F� /��������|�]m����w#�� ��|m�;��g�V�|  b  �� ����5��L�oO.�.}�׾� }�[�r�W���]�[��G�_eϻ�ѽ��o���w}V����� ����� � ��U��K�n}��r�m���������W�=� Š0�n�����5��W�Ng���}���  �J��U�`$)�ư ��|��x�ǹ�n�7uoO.��x� �  H���q �}e���ʽ�����{9;���P)|'���4�zΚh��� M(B���@ �Y�h)c(4Q�t
S���J �ݹ�QM�4Ў@
t�� �h4щJ ��tҀ	� 
  �� � i��A��iJ�B�N����ҁ� J(�� �շ�om{��x Q���>�v�}�>  |�n����Ε�� {g���}�W�����y9O� z7{c�`��c�o|��_ 4�T�)R�  T���M�T�M h2 E?�U%�(4�ت�m*)A�� S�BS=J�(2 h��"�&RTM$G�u�~��_�?��.h��kRz{���s��
��3/�� �� 
 ���AQ_�QE�D��*w�Π~���E������4�F��)�Xl�)�aMB��%���y�^:̿�}���WA����o0�ą])��]��aR�>�al�|���]?}��(`F�Jn]��������aO��eцc��~_��
B4!D�c��>���6��~��>́�$�Ɖ�}7��XQ�Ǘd�0�TÁ
���
�4�(m �4�Z`����eIn�4e���)���*F�u��{���<޹�\�р�z��u���_���o:Kݩ��Jq&��ώ,��	~���l�a�6M}���w����y�}��.p9�������B$��cMK�>5��W�
�tbJk%4+��Q�
Vi����f�}߷���4[����T�7����m*��E��"E>i�u�ן}αm�>#}���;u�޳)P֥�Y7G,W��R/H)_:��Hc!٢Rޜ6�qi������9.�&��6����5�Qe4�`ƚ�MB���-4d.�M��SD.���.p���>0��.��RgYtL��]��X��BRR|D�٣�z�a�.�]MM8��) ��Ė^/&�R$!HCD�l9�6P��Rt�K���41��]MsKx�g��τߦ�Cنn���;�a���e�u�����x<:�
�:���y�[8Js7�[8�3�SY�]ko�A���]��lh; A��!��s�Ԑb�4��Iu�(h��I����a��0��ۏ�L+3N��G���)�4i��K�Қ�7�&��k9��f�oG9�r�{���I.����.�� P���$I�s���u��8��e��f�f��*;4t�)�6�>V5�{�5��eHie#)V�+bF:��`@��k�f�: �SK�)�7	
V2	�&���$�FH1$"�P�`��]k�R%V)H`�jjU�X[�VF!�@"��c �B!GA!&�P��0��Hb��2kA(q"�C�`��S��B� Iu�)�}CD|��#��&�H���P��{����X04�@�
�"i�X7��hF�bB�(�@ B�D��q��d���J}Ѐ�"@�V�.,.��e�ɭ�����b���rzI]B�G	u� �b"A�bĂF� B$�!H�!u
��F!tb�L�$M�p�$@�,D
DjVflC:Js��P���7���Z��a�t}�c����G���XB�D������!
i��h0S&�0�B$I��XQҸ$�
�%$H�¦���0�@��"B�-$ $aj���5sa%�b�BT�b�!MF�&�D�g9i �  ��, ���lLx�hh0�n�7��}Irjk��@vD�X�R�t��hhbP4���1T�X�P���d0�� }�w�C���!����e�p��H�$���2D�P�
�06�i�H��Z��.MCy`�E�
�SC��*��1! Ē�!�[Ld"� E8'V#���	F��f���F`�*Hp������) �H$�R
Պ ĉ�
X�"�H �#"� 	�,Ta`, + `1$ A �ŉ P� �`�BD EH%VH��F�$E �"�B
�"��� �@"�HA��N:!t�"�	"F#X�Y �"đH��2YB2BR15�(�P�F-"$�#�� �H��A�d�$H���T�Z����
*�H `0.��fo��jk#��l���!Vd��lѸ��%��m�j�D���h���
��(�X$��"��!�7Ł0���@���h�Łm(E���� CYM�gat�8��"�XT� `q-�1��BJ���0eCXs���*�4f��"���ąCF��+�{bB
ؑxD�ih�'h�*l`�WM��º0�E Q�BR�M�[*�m1���ф.�SA����h� S6��p6S�1���-��	,HT���
�.�5�5�Mh�f�6F4����j��BWQF0�(�IZ%4������~�6`��(�
����Id�h22E�4C%2W [B�tGb�ٙ"�bj��H�����X�3�d�q����D>F,'-���tn��	S�@,"�
��Z�(*���&B�`��ڐ40�X��@��x$]!H�BC��aMT�+-�I˘/$at$���E��I	RY5�pvP���P$��0��XD�`l�n��].�)��o!��IM,԰�0���P��Bh��`D�M	�9ٳ,a}�|�٤�hJ�R<
���vK��CI����[��]�5��$B*r�Ho�`k��cR5%T�%��'fj$�B0b��`2�XKI��B�B��� H2[��4��Qڽ�DѦ:w��N�sZ�6��e4B�p��پ�͑��54nSn�Uӭ]�i#��A4h�4jp4��ܻ¬6i�SDMN.��Z3`l$�
}���BPt�$H�
��I���@�B`��xE��<1eGF8l
d�JhƎ���C��h�3r$a�j:H�4B�H��d���@�RQ�0"D��>�`HSFA{kB	)�I\�*���Ub ��D�>�]5���V°���י��v��.l��5
�[�F��2�	�	����	hԋ
i42���e9t���u�<M��m"�*��JU�e3:�G�~��/ډ���	M}�yvh"���2 �Z�Ѣ�Z�X��s�:�-ْ���w�s6&���Y�����3_j��^s����M*B�X4��w�Y��Nd����@���S���|Y���bM��q܁Ά(�0(h0v�̿a��Hm!td.�a�xO��K��!^�$k������>%�p�SK�cCXoY�LY� DH�M1�h�ώ�p튐xF���B��	M$���cXA�4B�cX4aBa�%5��`F� �H�#H0��
,0�B�`B�)��a�F��!$����#�T��4����"S0�7�k������|�=6MI��K�\�4��Ŋl8�������o��r�jk���>���@��u�)Ȱ�0 G��(L9��e兿d�͛�9�.f���r��u� i�v�����` m�   $ ���� ,e��S�hm�m�h���Di����#T�ܬ/3�l46�wk��hM\:8�e�N�e���Y5h�JN-�I,sh9 ]+a��"K���t���n��8��@'6�M��ړn�[�p  	 �  M�Ln�&m^�5�P
�e�� -��q6� 6�@��<5P�v�ٸ
���v�BQ�V�q����'Om��k^���[Khٮ�u[[e�l���^��,0��ݰnݳ|Aӆ-��Aö���u����pp �	6����l��b[��l�l�nݳl�0�f��l�]z�t�/6�a���v��[NH ��V��h  �` � Y-R���ڻk��\�̖��-�m�� ��6��i5��I�ݰ �  )@�l$� -��`�^�nk��eV�/+��v6�dڋh &� 6�c���h�e%�h�u�Vʲ�]U���T�0
�u�p�յWJ���oR�$ݤ�=%��'$ ��Y;^�N�����^�t�w:�c�/K����^�vأ֫�Yg�@Ӧ�F�    � ��G��~WΪ���7ٕ]Rr��C���S;{>�[Zu��� iS��4�J��V�U�(�U��m Im�e�[���f����5ur�J���-$;�v�RM,�k��k���$��d���v�U��E[VV{h��n*Wg�����.y%�Gm�8� Ӕl��8ං��zu X`�d���@keZ��.�@v� $H��͖�� �pHd�T׶�  ���h������i�m���̜[vڔrA[���hrKݴ���h �����	� 䃜���l z�@m�sE��6�3l[\$��V��Xપ��U�X8�m&��ә�[pt�m�k��-�[%�G%����m� �[�9l &�rY;�3Ze��hHI��ph�%�,� 6ݑ-i�  m�e�j�q4V�05@A�E�V��K��l�W*�Rԃ�9�@�f�9��l�&������@۶3l�$v��$���@m'N���Y'c�m�q����u�I���4і�s� 	%�n�Yқ[@m���cv����m����|�P+<D�,�HŶQ��]�:}�c��Kn�L� �m좭U*�5T�b&
��P�ۚ�+��e�$��f�� [%l�r��A�\9m�5��5����dn۳ f�f�5Q�ϕ����v��eZ�!�/ʾɥv����փ��LH.�i�:�Ns��m�`�aCn��'E�'a!m -��[wn�*9�R�GZ�X6 ��;,����K/��H�^�m  �:�;m,�k��l�K$��d�m��-sc��v�S�1.��R�UKh Hm��l� ����\�`��֟8H�y�_�؟Z���  ��vMd�C�Ee� UV�'��������ˍ�,�۷LYd5��8�:@���k���@n�m��� �([��� �0� -��2�K0L�BJ�UUU�ڕꪪ�  U���[նÁ��[m�Y6�$�i���mt�hh8m�}$��ۭ`h�՛l$8   -�[%� m���t&�լ:�/Zm�m�  ��  l �kX<Mu$�m��l� :$�ҥ-�u@�e��#mƦ�����.ٶm�R�� 	%�!���v� ��l�@��I� ړn��mm�m�շm��� � �u���� mm��`�` m�h	6�[E�i�� N���Xm��!pv�5��H �8    ���l��y��z��m���[v�fZ u�� �ж���l���M�]URl  �����ml��ڦ�f�6j�V�඀ �\�a�"{i=AU�NԶT�8���Uj�]�	m�`����+[v�\`	v+��J����T��a���i�N�6� s���[S��m�  -��ޠ Z�	-�]��  m��8-J�I�UJ�S�j��TZ�U�l$�z��@8�iM6�[sj�n)V�%�n�b�����)�q!m��gQ#� m[�j�6e� �m   ��  @ m�      �8 m�5� -���am �a�a�NP����	Ӕ�V�BU3��q�댣J�u[JKmuJ���KUm�q���I8��&�H7mzΙ�m 8 A��U*�]JʁP    I �  ���  �`  -�-��      � �      �    [A�� ��q��l@���D� �  	� �  �     �`  ��[m��l9��hvkmV��o���H 6�$�iXm����qtj�$�@	�@����  �m �kM�    Δ�һs�][���U�ڧlm���@   z�@l�Ĳ��6��� �      m�  $  h� � �x    �  $   ��   �   H    	 m�-� ���  �d`     �� m[m�p�h   oկI�H �m�R��6�'f� �b�1   n��� �!��  ��  �m�[mT�:w<@[@K(8�i���n n��@�q24߯Y<���mKN-�i3m��ɛl�m'��    H   [@     ��    m�6�   �b�@ � h�   hH  A �	���n 6�m�G m�  m���s����I�M��E18kh6Z�.�I�۝4�kX�m,��m� p $�#�����Hm�tD萨*��{.ô�:vf�-�	�K$���I�J�$��!�pc���X������WSJ�m  ۮ��zڊ���]�����D�UE�h ���v�4P� H���7�.�q=�y�;u��m�pn�h1�-��U��vv@W�wI(�]��t�@ �ۖ�' Xm�mmZlմݳl���  7];m��lk&�� 
�8pK*�R�B^��@m�[@   X��H 5��V��ZmAI�겛prpK��6[@ ��඀   H���6�E�Mn�m[l ڒ�mm-ioP2�[AoQ  ��D�m�ְ4��7m$�<����q�j�
�'���m�m�`�K��l-������R��q�M�jV���    �M�VJ��]���4r�T��m�d� $���l�I}}�m��@ l-��     B���l 0�imH�C��*��( �z���j �G6��B@�H$۳o�JqJ�8`�ۄ�p�m8[[v�[d�-��M�I��@-�m � 8 ����H���l�T�Kҭ +�R������� ͮ�9%�6ض�$�mm l����kmm�����i���� ��e�$�&e������Ii�@���-������޸  J�������7m�Ii�O{��Y-��v��[@ h���[m���\m�lHS��nm1��i�� ImHz�v� m���b�J�����mm$ 6�u\ lsM��[Cm�m���f��H$ � �RvN��`�b�n�xpm�bAn���l���8 8    6� 4Yi� m�-�$ [E�*�����j��Z�\� ��m m�!z�m��b�ڤ��r_���R�V�A���Hu\|����S m�� 4V�M��$��gHq�M��XL6�[B@l���# -�v�԰6�Im����ܽ.�Y�I p r���l��={zm�r[׀�,p�m��$H8�mo\nI��[vE�e�R��⮥�v@��6�6ݦF�T�9% ��A�pŷmS`m�u	��ۚ��4����45��l�m�hj��)mi�fNR�T̬��r*��H�mE��RKԢ�\6L�2�*��&��8�mnH�jǵ&��6gm��J���l�S'/Zl��4��6ٍܰ��YM�j���ۦ  m�{��oml �cI�[�� �`�a�����l�l ���Z�� QM���1R)	��C�����!�?�T ?�j�V�]���D�O�� 	� P�!�CJ���AU�P+���ؚGå.�1O�
N< S�)z(��Q8
�;P���U4#�Р�0�PU:(ox	�"B0H$X�b�B��lP<��P��
|(��U�(�˴��ʢu�E#�C`�sM$<�� ~�P �`��" �%QL�W��P`���D��4��B�P@^"��v��Ё��<�!���� ڢ8��O"�PC�AO�¦�*U=��2!D`C�C`��:" �1∯TH!��O"x;`� �Q:�Pt��4&f�C�z��@�*/Q@�xT�@Ċ�Q?�QE~Qڧ��U���W��GlpRM��q�wv6�u�u�{�G5�񍝎�s�7��B�]��t�>d��N�2�,4�[8��Ӻ�e˴�+Ɖ�v����X�Q��1�ݨgOfF��:��X�[˳B�"f�+E&��˻[GX1S�\n1��Ym�M�n��v�e���M͆{Y�)�=qH�@�"�&�70M���ot�֌^�X��j�]�9��K�a�X�X��cuիiэհ�Y����F�2�T�5��KV��<;���0f����.6��8���dA�ێ����9�ZXA:K�ˠr7���ps;��M��z�덚0F=�c"��;wҥb�Y�_g�"sm�ӗ���3M�b5]:)�9U���]y<���i^+@�v�G�ͅb6�ܲ�!7��JP$�.���F���Lbw�]�2�#�����m��䨸�@��F��ˉ� ��в@uP�u!��U�mv� Xke2hx��۳�D��XЈ���UB����R��V��[@�ۇ�`�[�9	[k`(�
r��7I���n���*���
�ڸ��FqҐAPP����� $���V�in��j�`�j�]f��et�!=J�7NNZ"�3fC�Y\a��9�bޥ��c�&�
+bBe]ڃb|�	���vzj�j69�O&�K�gY��qq6#C�8�Loh�����kr�9E���qGGm��ԫ���s$�QI�W��v1�ѐ#&�9����؁u���ַj��^P�mƨե�6f�1!2�!��ƝX�V5KX�ش.��K�c=�ݴ��M�7%怺�v�%�U��Gm�;vEK����N������tY��Y�H]l��9P�ڞks��v+��	Ҝ\�f��gj��<��`�d-���V	��<����K��Z�(�#Y�ɝڱ�jvft;��I�6f�w>��`���s�mzլ4(>@�xU��� D�)��'@CcM'?���9��}�߅��wm��]pױ�cq�t2��d��p�7���e�N˱z�\�=j"��Mk�
��{:U�k�b�Q�;Ta�.ݧN�ݹ��jۜ�� 6�[��W`�5���ٱ�id�-�	-���c)�/��(hڴ�M����׵����YѶ�<T�烶q�1�=��Y��-rs)A��L`�[U�:��.��B
�;QӼݚ���&�f��4۫5�p�v<

l<���gd&S�����yܯ���o��o�{Ճ?c��P��ټ�o9:��麕T�l�m��z_BQ�L����_zh�l�9����4����$���p���J�z:p�ֵ�F�l���$� �־ �W�{�Ӏ�������,׉�&�M���ގ��Ӏ>����>���ٻuTaj-c
�N�v���6Ӌ]K3u�-�롗b��N:m��r�&�z:pWN �־ ���d{�RۧQ.�m�X���Q`!�� WDI!
��&�T�Yh@A�t�}&�ϳrI�Ҿގ��%�5��q4-�� ���`��Ι�޵`v���̩�Hf�jx�m�i7�Z�	�{8+� }e|ҽ*Ʊ���Y�٩7�OK��Y]8�+�[_���������C���F�xc����sкq�8wm��ЭM�X���Rȩm�n��-�� }e|�+�'���%���䤆,sp��l�^٠OK��OWN�����X�,M7`��`{ٶ�q	&���� $E�#`$1 $�D�~�znI$���)Q����ch�Z��=�{8	���z��J�	���i��M~֞6����p޵���ޛj��I(�s;\ܹ���rT���K��[%òu�˝^��{�o��{z������m�F�X�R ����{�4s�s@����e�3Z5<f6޽M���ޗ�������|ҽ*Ʊ��X�u�&��K��_WN �־ �W�{*-I1jM��By���/��M�'>��rI��ٹ�Q�QP�lM�S��� >���7$�f�{5����ћ��I���|d������/,���mI"B)q��qR�H�W]��w�%�AT''G3	�k���ƭՉ��i4� Y+�=�{8���/������yJm��4���=�{8������=e|��+)#P����w�S@9�f�r����s@�*�G�H��� Ґ��3���;y���=�K=S��d��8m�sM��5��;�/�ns��=��`5	J��%��h*h��G��q	������65k٥"N\�Ju��j��hݰH�Ǝ����˺�m��hŵ��4p���V�v�2uc;����2�8�kv�Ɍv������9�v����qV�p�2�Q>��W�Wj������>7+�Ώf��r�`�#��J@�OI�>kۑ9'	:kVw^�Ɠ�ז@x�V�S��nD�L�v�x2�r�+�b����Iݬ�Y2N��z]��y��17YSOM��7��NI�-��4��h9l�Y_쨵$ĵ��c�m�=]/�S!���;����4��R�)!�$��4��h-�@�-��$�����Չ��i4� z��z��J������yM��ԋ�S4��9�w4��h9l�n�:I.U�G&�[��T�.�B�;k�g=Qg�zs0�)�:��1%�`�]>�j#�8c�d�L�}<h9l�[f��[��^t�ǊH��c�iI7$�}�f����(������~|����Ӏ�[.!����1���o�=m|�og%t�z��}�^G$X�)ܚ�]��٠[��@>�@9m�2�����6�Sj��ץ��O��� ��v��s@�]1W1��Ȥ#�$��Fv��nێ��6��;kuzݦ-�qٓb�M:V٠�$��z����ޗ����p�dwF�<C׭&��[]�BJ&L��V�>,��]�����)�nf�2Ԫ�n���mX���TBIL(���N=v��vG�z�,lf&��O8	+�����������/:J��$Qı�4�4�-|�+�=�{8	���O
a��#"ݳNF�l����Wc9�n�V��3c��� nu��oMH�Ͷ�}��|ޗ�������W��J��-N
	l�m��m�興�79�`��`��}	L��usm�9p��Tڰ,�� }�_ z��z^�QZԶ�K���e�D%3��v���z^��33/�Rt�=����Hx��ZM7���ޗ����������n�Q�Y~���"�A��[Y�.��Z��VzI4�[�Ь��n��܋���ŭ�ޗ�������|�+�2=��)cnb�cn��3�������w; ��v��j����:Rۖܘ��g }�_ z��z^�z�p-��m����z�7���ޗ�������|�h�b���[56�z^�z�p޵���`\%�"���Z�4��6)��M٧\��l�T�l3Ff�6��xNqkeЙ����Ү�h8��ݗ�ќ+��=�F��=�pt��s�-�V	v�h�%��20��n���;�n5���٠�]qW���T{l	f�Ps�n��=DC&��i�����q{�I�:�Qf���rfW��g�N4�0u�B���ֻ��Nܙ����L�z�!��k���J��y�����w����;�������#<=�\��a!F{R���ޫ�Pr�gDd�L�.��j��u��mX�����v��v�/g(�k[ŭ'��$� �־ �����p�Ӏ�엃Q��`�֛�Y_�og=]8��h�>��#�M��@ԓ@�s����%��=e|��;�jz��t�Sj��k���!D��?�����s@�K�19LHs$Q��Ͳ$�v�4��ձ��;h��'�6�g�E$F9���w�� ��-���� ���s�_c ���?7"�ɠ��d(�D\M����ץ�fn�z�U�<x�jm���p�Ӏ%������V��&�6�jo8	������W�Kog�;cRcQ��cn�l�=��)����޵`g��`tD%�ɞ�P�,f�n�a���[Y�јi�솊��,ok�9�M,�����v����m����%������,���yM���N��Թ
�݁��j���s����ۚ�G��*�:Lt�j�;���rI�wٹê!�ARD�<|ºV�b�M����j :LM�i��P �4hk/�ECAr�2����X��� ��A� B��@���&Z��J@�%kJB�$�X,��H�!!	,��b���"������1�`@�"Aa�8B$R!D��G�Et;YegQT�sx�|��l��T:D/
�
��8�����v��Tt��A:)�*�X��|�����SY�5���ط[8Y_ z��	m��'���}�����f$޴��Y_,��z�f�3s]��Gw\�êt�eP��].{bq���*���ڣ�\k8�r�l�V]�FG����rO����4��� ���Y_**��k[��1����yK�-��>��Y{8qZַ�^���k{����+�%�������2��Q��P<n�[v��vnm�=�K	_��!�C�T~�?f�=���5�4�����	e��=�^� �����s�ŝi�h<�?�9��P�F�!�v�������Ӷn�ǧ;u�/P�47n;3�bLCo>J�� ����������9���1I2H4�4��p���������p��qԓ�ى7�S|�k�=e��$��=k�'�WV=b��kf���/g%t�	�_ z��TU[lCx���y���$��=k�[_�͵`d(�"Ė�(���墪hE21g�uЛ��a�6G���^�[�r7
�6G���v�{���n�#$^Źۛ��'-�������h������v4�2<a�m<�b�t���A0zy[u�6� 7&�=b�hCHl��v6X]\�TuU*���;j��{uWi�h(V�,� 7�0�6u�5O�I�7WΗ:����yasՍ/eԃ8b�ш�`�뮟}+o���a�l<]\�Ն4�u�|�P�8T�n$�� g%�K�EsnjJ���I2 }�� z��Y{8	-��>ɖ����٨ku����Y{8	�{8Y_��sq6ĵ�כ�[|��p��p�� ����on	��$�6��� �W���Y{8�WZY�5���ط[8Y_ z��	e��$����v���5��J�뜌:vd�۵�W��n���.��"z��uǴ71µ�p��&����K/g%t�����}}4�G��(5 �,R�4���?~��3�I]8Y_ z��	U�Zl��4�mKmX�����gD$�L�����޵`n��uM�R鄃i$� �W���Y{8	+��w-�&br$�)"NM �h����Ӏ%��l�cM��4ޱ�a��-`)��
l�{�i�;]�W\��8i�u��o^n&ؖ�Z���	e��$��,��=m|������[1�1��$��,��=m|��px���LNF�	) ���l��D*5�@  @Q�t
K�Q
���Ձ�k����sU9S3M���޴��[_,���Ӏ%��ի��kb���ē|��p
!F�_�7���{w]�Хa�P��<��1��tgGc�Ժ{�Ͷ�Mc�P��q�1S8Ig�\5߀[��@;m��l�;m��-�lI�Y�0���$� �����[{8	+��oi�blk��S|�k�%�����p�����&�K�zS|��pWN �١�r�4gK^�I"�$$�J�������Kogt���]���� Iue�Kd�9�1PI���m?��۾^=5W̑��jm���h唟���4�٠v۹�w�S@��c3wSf�57�6����Kog%���٠w�:�EH�ŊA�'-���Ӏ%������Z�֍M�ƛ�M�%t�	m|�k�%�����&�h��OL�&�W z��	m��$��f}{�������#ٴ�G9�k��R*uo�u�������qlA�ZpPt�Nݷ<�m�����^����F.���l�b�,�D:��gX8�clKj��>2Ʊ���q�j��]�ۖ�Wey����ᝂ��c�.��h6V�Ȳ �68l��Ջ������<Uc�z8�vy�Ô����gt���l�U��Ba�{��\�Ӷ�v ���|0j�L�����z�+^�N�鋎]X���s�;��́��0�M�nJ�m�����	e��$���*�=���bm�X�נ�7�K/g%t�&�W z���ī�����X٣o8	+�6ʸ���K/g�z���z�m�=5��%������^��v��5��bI�(br(��k�%����[��Z�	���YD�\]���SӞ�&7g.�(�:1�zm�ֱ\0W@�=�S�++_6���{8	��}�����EkoZ32�Y�e�.f�w����
�X���'t���Q	-׽��'�z���s@���1��`��iŠ{e��=m|������=�-�5�c�O^�����z[��I]4?��.��=��<ǎ23#j i��z[��I]8l�p���������Z^-r;]��l�k�3��An���S��qv�n"���N��+��L�cU��Ӏ��W z��K{8����(�rLdɊ8�.����?$���;}���v��5��bI�(bq�t��=����nڲd(���ݛ˶���SȠԍ,1H6��9�w8J��{e��=-|��޴���o�����[��Z����z[��z*`�V=I~m��Z-ѷ	�c����hH:�X�҆(9�"cU�-r-m�h�����W zZ�K{8uڴgr�Bf&���ӏ@9�_�og���-\���,M�נ�7�z[��z+w���W zZ��%]�jM5��6��W�rO�}�nI>｛�hx8!EU7�/3@�^����8"dĤ4)j�K_�og�]8���o޹�[ٮ����r�y�<�8�E��B�X��z Ԗ�+E�k���m������nڰ=���(�!���`vWWSȠԍ,1H6��9�w4v�h�j�K_"���66��-o56�f�,Nn՜���7���֬	EkI�[�=F�hI��Z����z[��zWN�2��Q���=���k�=-|����t�=���l�@�`H�&���k&�D�E153@�K���!	��`�� EHg:��F!�'�������$�B\�ut�"���B�F�v�T� m`�	��A�$b�H�!
0"B��4�@��Iu.����I)���5j<`�#,D�F#��Ea jBc0c�/���~�h� `�M"@6�d5􆁒�� �b�1��4�H!R��F� �"J��"�"! B�@��"$@����H"�h�B�.�4CH�@��	j�j��F�D�A�F���54��%$�
�*J�+]+���4����@�$j�c� �V4�Į��M��$%5�0$�I��Ԡ�� ��S�$**A[	CQ�X�MEI ���c�,�JCL	��]kP��T�	XЈ�!.`h�P4����aJT�P4F�n2�蚀A6!�ݩ��"Ќ bi��!���?�n�r_���J	V�-,��K���Ʒ�v6+on���rt�a����^{F���ŖC�w�xL���f�|
ٖ��۶�.�� �S��PCS�,�lf�m R����$h�klN3Z�cn<,�t�r�ۃ��n��UQ�_�8O���ݵ�Pk�8t$/f�ɥ56����;^���v76Ұ�0˝�l8V	�+V�N6B�R������SF���$��i�p�$�b��z�c`q�d���wU��J�u=�����ݶ��zv�]�0; q[uy���1=G:]���s\���9�C�ҋW ��#]�����V�ҙBY䕧���;n[n���m����
d�t��j��j��1�n1�N��6�j3WNp 4�2Kmd�i^3í�ݷa�eUlkH�9ea��vB8��|��5?:���r�M#���X�+�f���S�f`:6�<*�O[h�r똝���ժ�j���G��dwmZ� ��r0L�U*�UP��U���}=���Y�����mf��e�.��� �� -��e&VWE��Uml�e9�(;�ys����VW`�A[t�R��怨
ځ	Z��hj��eU�V�]UJ\�Se�,z�{�9KβZ�ݩK*�T�٬<�N����0h6m��U�$z���q�lj^kZD��vB�}���(��5=d��ѷ�	���Y�<96Q4�O]��v]�)�d���.��yR9��kHȄd�]
�y�Uƞ�l*ֱ�!��l�n��;u���[��U��p80�Gn5@VT6Bw,<��ln�2�aV�ڱh�J�P��v�]��v�dvpQ�� ��t�ZY�I����^�"tY�t
\&�3b �<AN�V6�ٖm���Q�aD�OU3M<ݓ-T����5C�)�J�i��ɽzu�l���IQ[��bv�i(��a���.\J�HE�ʛ�2s�`(B�m�i�T���{��{��� ׅh�l�(��ww���?�ɆaZ&8��)�xsd�/@���?~[�eN3�0�9�\�oO$_:}-���^>�tY�o�RV�8�]LBCdf���v�'5�,lu�0AⳲ������%u�=�*�쳝�&�h�z�KF���m�is�!�g�Cm�]t�j�5c�{���a�@��n�buvd�ݽ]f��+�ӭ��.��Ftl�\P�Gntت݄[��u��u��SDҼ^��.3	�r��c�;Fε��p�Т,��c��袈rx�������Z����\�*�3q7�5��6Ձ�ץ�	DDDɓ��`����m��>�Y[x�r9L������]�{7]��)���Vo>,z�Ҝ�i4���y�5������Һh]�����EH%�)ܚ����t�=�����g�½��Ύ՜�X�$8�c�x�2���f6l���]A[8͝)��J��{e��=-|�������U9�U:*�`zsv��D������PHŃ�(Ya��v�6Ձ�ץ�D$�L��&�i�2,qD���zh�;e4.��g,�x���QNM��Ձ�ץ���ڰ�
"&s{�����b�"N<�D�4v�h]��;l�9�w4�Qql�$x��H�c-�d���; �klu�3���`�a�۲�Y�Ri�koxl�p���zn��
?Hf����w�K�t�2��֚���������R�햮��ؑ�����b��nM��s@�R�g߱%�����EkoZO*[rږڰ�Q9�zlN�U�~�١qv��h�ɍ&�b��Z� �H�I{8E.�b���B]sw7cP�W[Y��
���/.���p�jY��6�s���b��>���^�E.�����=�X���z��-M���p)w�'�|���ī��Ci���D�p)w�'�|�����pg��,Ե1����	-|�����p�
#WL��́�Gu:R�9LI�z����������K�%�@��5r9$2c�ЁHħH�@�M*���	�k5*��[��<��3�a�3[M���p)w�$�����X�m�I�l��ko8	���
&Cw�������W���x��T�4���ƤZo�4�l���1.����-w�@�B�Bcm91,r�a�)�ws�3��X��6
gw��Y���M˪N\�
�n���ڰ>������w�; ������BH�J�Q�����F�2�[��5��kR��^�eӮ�H���x�5�d�XZ�i�ع�!���ק��^և��.*�͋�j�kTm9&��s�T��,�l�[���R g�c����n�gl��C���]�k��o@����g\�Rm���OK��w���!�j�����7r���\jl8k�;l�GA7ZKK�qi�݉�c�bwf�Um�ڒV4��^I��o������.�������|>9�e1�,N1�ß���L�:�Mlֿm
u�}g]uE��u}�� ��v�w_�_�3��Xß:�*��������|�d=��v�ۚz�V��2�(�qd�^���k�=-��$R� zZ�	WP��l���OM���p)w�=-|���+[z�`��"[N�Vef́�
s{��ws�=�w4��v�����L"�D���˭�d_-�94�#`�=4um��K��v�--r.�x���K_ }m|����]�&Ky-LI4�bM������L��Vef̀fn��Jd��}E'"��QD94��Ɓ޾ՠ�@>����ը��MB!�@�K�%��>��ֺpx���qf���F���� ���Z��H��g�<[sSoD7�[z�<vYu�2[�{nb%v��n��볶�v�6���n�٭&��o^���k�=k�"�xK_"������᚞$��=����ɻ[�`���?n뾈�����D��O#lRb���h{u�P��˒N���`{��`n��uM��q��1���g����s���9k����"�������uL�R�A*����������]�	-|��鹘��L��I��K�k��y�m�i�r���
���Df�s���r3�=+�"�x���[_g��� � � ��sV���5�\�e��M�<�������v �6667���6 �6667�߿f�A�����o�؃� � � � ����Z)��.�4e��v �6667���6 �6667�߿f�A��������A�A�A�A��߮�A�����=�!���e5��˫�͈<����$Q5w���6 �666>�����A�A�A�A��߮�A��CƔS`���߳b �`�`�`��g�~��L5�m!u���͈<����g��b �`�`�`��g�]�<������~͈<�������ٱ�A�A�A�A�M?�w�c����ZW���҃�k��Kԥ�9�a��dݸm���c�.L�A�Ը�/��`�`�`���~��y�~��y��߳b �`�`�`�����؃� � � � ��g���ej-;���������r���~͈<�������ٱ�A�A�A�A�����A�lll}����A�A�A�A�����k%�\�$��SZ�؃� � � � ߿~��y��߮�A���:�����~��y����lA�lllt��f��f[�3Yr���؃� � � � ��~�v �666>�{�؃� � � � �{��؃� � � � ߿~��y��j�5�殮L�ˬ�y{=��A�lllo���lA�lllo߿~͈<����g��b �`�`�`��x"	>�?|O�jkYLՙ�۟V��S�#q�[���ȍ��n��=��3Y5�>Ւt����b7/P�ҩ�+������7Z���b�q���ŗ�"r�m���^%�bn�%��۪thq�]���a��"�2�P(�U����A�zx�{�c�j����㩱Ӟ��8B)s���%X#�<�I�j��C��6e:��g�'錜�gv�N����ӟ���7B=�i�����V^��Hsٻ11/,.�χ�u�鶹<��['mff_?A�������lA�lllo߿~͈<����g��b �`�`�`��g�]�<�����eb7���t�UM754ݨJ?
������ٱ�A�A�A�A�����A�lll}����A�A�A�A���ٱ�A�A�A�A����52�k2�B�kY�y��߮�A�����~�y�~��y��߳b �`�`�`�����f[�Y&��j\��˱�A�A�A�A��߮�A����߿f�A����߳r������{���"M��ȴ��X��v��f�ٰ̬9D$����X���h�c =Og4u�b�킶��]c���]��il	[�fr������ݛ2�g��@��vn��sJ��t�]9Ni��[�dD(_�"�Q*)�H�J�����7{��~����H�/�%��$y���-w��37]�B_%Tg�|����l�5�K7$ś�{�Z��k�=]�C��[/����/��)x�r&�v�w]�г�t�v���37]����`�H�Q�űr��3�Jh�ݍ:�19WKe��\Ʈ��r�ϙ��4n�ʪo���6ef̀fn��!B�#�}������s.[
M�Rڙ�6u�� �m���h�վ���?z7"rD�s�h�����M˟��#_I�Ґ�0aII(�a����]�0�ڏ&$��0�M*��������18���$�HE" ���H�X~p�,E��j0���I����]H�t!Q\ڡ�3D�RW��? b�AU�Q��L ��E���j b
|����Pf!B�I~Q
!��Qo.�f�ή�=�ݍ�!HbHq�ɡ���s���;����$R� Ik�,�W=X�֓i'2'&��e4~�e���zh�٠\\�.9��x�1�LP$N)��x��h�Ke9�#��0ܒΎ�����1)#��7���- �m���{��gs�����)T��R):s`�f�}m�-��;�ڷߒ:���9-ӥU4���v��v�^�|�D/����l��S�P�4驔)��M��Ӏ�K�%���������Z����m�kL�$R� fn� ���������f��s��s�	�c�������1kV\����k9������]��ؿ��~����>��ֺp)w���y��ZI3wDГ|����Ӏ�K�%���e\�bck[I7�[|�t�'���Z��+�'�y��OZqG�n��_- �ޚ���t�=��ksqbL{�Z������~~��X�͛R����@�F �P`����Ri��-�n�LY�2���m8��a�Wf�U��=�](�q]n�;j��?���|\v|�|^1Z녥�2q7%�\M��-��p��Зk���lP#�x�W�h �n�7nף��:��^M[<k�u�� [�̲,�n�T�M������	Xx���'H\�p�u;+!�7A&�lYld7�s;���A�c	���n�{b�M�\I}�����;|��\?��8E������6�ty�D�����tؓ>����GZ�e�.8�q�iȚrPs��@岚x�w�$��-�C�x�7p�lI��s�S@�j�v٠^ٿ�#�~���HbRcn�Z��4��4[)�[��7&4��4�ƤZ��4��4[)��W��h��lnF�8�D�nM �����{||�Z��4��7r&'1 �n��D��q��a�����ډ.s҄2DQZ:K#�<p��rdRM��h��\%��>��x���4��6��f��rN����?�A(�D����a��; ���=���<��t#7��2H���h׶i��O�Z0�,qH��ӑ4���uWoS;�z�a�9���̩�({�{��jx�o�����xK_ }e|�G��li$ر`�a�<�M8�s΋f�uoKƧau�d��<65��׭f�y�3��R� Ik��l�9l��k-�I�G �sqp�� ���Z��O)w��Is��cr6'#$crh=}4[)�Ń �F��P�N�`S	d(�I{����`��`nbڷ4���m$�=m��Ӏ�R� Ik���ˏ��@�/�%��L$y��w��h���z|����e4v����r��kW<�@D$6�<l�`�%m��\�MZ�"�7k�;viN9�{=:���@�^נr�O�������@����X���9NM�{^�3;��-��- �m�:�FE��,18�#�9]�@�j�߳�E���8�z��ݪji�2Z�mLӛ�DB�"!Wm��`�|�ӹ�a脢�!(R�(��Z�́��u�mT�73S4�Ks`����P�����3��l�v��-D�L��b��,�8�{O�sr�9QZW��r��<�"����{�����iD��nO�9��r�V��>ՠZ�&U�V&6���x���z�پJ"ɹ[�`���?nk��P��z_lK#15�'�zw�� ����ڴg-��,x�
���tBIL��; �o;�[�a�f~W��h�z,qH�c��&�}e|��x	�.���31L?fq���߿{���NV����fn{4�j�v�I%{cf���Y n�7:tm�Ӡ�3�!��(lXSmt�;θٵ��Wlѻ^m$�H�R	New���^:�h�x�^h���v�v��86�L��q��36�"�I�12��m���d�ι1���$vN�l�.5�v�a[qC�B87C0��A��p6�"�-����n:k2fS%tk����~ڨ���s��3�k�cg��D��FJG��ѻ#�E�ؠ9 -ŗ�g�����GN�A��H�z�����h{l�^٠}{*O�������@�,���}A����7����ݛ�IBG��zE&5�s#p�}����[��t�=2�i6��ޏF�náBQ3�����=�K�|�D*��v���l�Ln��T����Un��Ӏ$�����������O�>]����E�93Cc�^9]�lS.3k�B�Ŀ��}���-���I�>���`���=���DBQ����-�����,x���JC@37]�P�KbZJ�c�vmf́�ץ�DəA��S���SsSM���π�V�=]8K_�Wn��t��UM��v�s�t������a�
"g;y���*�������jf����K�w�� ��v+�h�ڱcdrby$ő�L��˭��yu�;�\FE��[�;e���h�fu��������&E�s�n [�M ��+�x	������m'��{��o�=���D)�:���՝֬3u�(R�v����F�mI�I4���@�s�ٹ��E`�HE$ �g��u�����%绍!�I&��r�Y��X�s�nk��D)�}�`b�뢉T��R)��i� ��vЧ;y�:������V/95?x�e�%D��]s�̖��s�흮��uŶ�[q/Ǝ���o�����M6��ԁ?���=U��L���%���+�$�:C`*����[�/��9o�Z�{��h/l�>�{F�7�q�p��6/nڰ��g%2go;:��@�����) �N~m�C߳�V��@3����ץ�DR��$��P��BY��~k':pļ�m'����&�ۚ��K��߾���9o���3-�U�F@O�ƚ#��m	�㮗`���;m0�dÛj�d�����������o�����WN ������ ;��^�����2nW��}
"d7{��go;ۯK�(����ｭ�X�4��}���g�"�w>,Yϋޠ�r��n�UJ�&[vDB���vw>,^ץ��(�3���mt�Rr�!�Sci�ֺp=og Ik�Y_��LG� 0��) |�)�J�Y*8��	���>
� �F���@�4���b��*mB�X�Y�� �ŀ�°�A�I ��P�1"D�BA$��HĀ�"U�E�q"B<҆0�Cf��w���$4�xBu%�RF1��bPV@�HP�E�#@e%!@�@T!AcB	P!HV<4�uI#^�������{��߿�V���š�����8���v�׋�r���4��+d:d��r�1�-�1�^�ݵ0;,���4�������*P���m5A�'��@M�kr�H��Ķ�*F3��U�kv��[��7:�Ӵ�`"8���&GZ�uvvq^���Ӭ�;I�#��f�WZ�抗�*�6�eXp.v�1ӭɁ�F����m�Ɲ����4��e�n��قڃ��˽��@%u�[Ie��ٳUM�% mg0m��Sײv佺5��!��Wl�r�TL�1��+�KeP
ڨ�k�>K�{K<���G3�������[����]yI�n5J��S��g�8
ֹN]��x���T-�vLj`1��mG���2����j�mEb�Z�"��Ki
�W�W��BY�մ�9I�7i���l�4�5l� �:�3�
�mh�p<Y���PI��6��[�F"6s�)��r;4�U*�F���R�

��:�Z��R9����ڃUΒ����n���UP��T����j���`+�U4�)��:�;������i��]�F��/,N4���@U�@R��UR�@R�@�VL�m��%e����J��mU<pJ�Z]�E�z�(�g"H-WJ��lA@,2B�s�q�lk�s�uK�9�{ �ъ�մ�$*m�3Ȏ���8��	�vl6�e�m��m����L�+��&M�r<�m˹|�MI��D`�]��K4�mx��+�&��cl�6wf�u�Umj���E�
�[)AHĠ,������7j����a��Ŷآ���m�n��[=(��ݬ�6��*�l�;��<k��B��K���j:Uؕ���+���L� ��P�Q�J��qV�m)���V�Ъ�wm��[-�.WiT�&�[��,7���k^u�tbPA�ێ�>�@V�niZ�G0=�:wf�n���[7/$��sD��4��w{�(�>N���Z�< (�E�
ySG'zM�C��ݱ��.uOl�:��w	�.;i�-[9yXz�m����^@W����xa��#�+[���v�l��m���s�=V�m����X�l�b܏\q��m`����)�@��:�I�Cs�`s<����V+b.��\lt��ҷ�=�m÷V�Ê&B�N�7k��m��\�/�/E�\Gb���%�նG���XP�b���-��,O�w>��9Lp��8n�RwH7Fy�G�9o���M��f���2^�v�������x�8IĜp�{=�nh{l�ۚ�(��C;�u���m��S��y�Z��+�=k�3��w(P�MӺ�U:cnT����7`���z�Ng�� Ik�,���X��ꥴ�a�
';��VoZ�ͳC߱.z�h��Ĳ2G��"�,^�ٰ��`�5��zXDG;���%hG��c<�#]H�j2t/�(����c�2��������ۦ���d�L�-�����~��`{u�`b�f��alX�D�!�I4��6��_�%0�G+���Ł啽6���DZ��X6$��o�����>է�-���s��@�����BL53Rg3�Ӏ$���W�z�N�R�i�M�^��L�	-|�=}>���w9�M�mJ&�'�b�YI,���Y�����t�gY����\��qs�(Ձ�b���ű_6�������S@�s�������=n/lo���Z�=m��Ӏ����Z��+�'�y��Ckf=4I��L�ܒw��ny]E�RQp=p�$���`n����Y;t"B��(�J�l�䒅Uw}���v��h�vS@�[8�RD�F%$��������GN ���O���N(ы�r��JA�ݭs�1�f�(���ڠ������::盶�Kv�^�/c��37_~�=����^���8G&	�7���h{l��l�9]��"�t�m�PT�2�7{��~��g(P�)����l�w��5#��œi�4��mń����q	t
�/Т��!�^&�G�5��f���/���ȣn6�Ȥ�+�h�vS@37]�~��`}
#�f�IM:m�R�2:�튇�HƩy[��je9�W�Z��YnYI9_(ݹ��n�Rc�I�>����	-|������,��f	2��SM����������v���@�s��8ö���i,lJI�^٠r�V��ى\�4�zh�-k"�0s��ɠr�V�������aДL�����=�MJ[ƓL�Ox	���%��>���}�{�rLZ��֡I{��&�)4]��kq�Za�b��4#"��r�)Qqҗp�kz2X�o
<���1�7ib�rm�v�gK5Ӓ	��κ�)CЉ�����r�}k�u�e!|m���b�h6N:5���Z�P0R:A��vN)��0�&�n2{q��x�ܾ����gu�mb�{p�-��6��%wQ�X��4����9���p$��:�MՎ-��{���v[ۏ�5НZ�����3�=�;8�«��ͭ�����j	�Vl1OP�#��� ��; ����������J#���Ł����[�Kd�T�j��ۚ��J!L���6��ŀfn��J!EQ�r���*n]SuT�r۰7����&z:q?~�%��}e|��Z-�� ���%
q{/K ��v�s^���Z�Evb��0�'!�����(S���ή�1{�����/���]���[\snS��=�8_j+������S��Vj�1�l��*��s]��ٰ1{�D(�(���;����}�Jr����ct݁�ٽ��	(UF����ٺ�����~H�/_	�y$$�)�Zλ�Z��+�=U��J)u��֞�&�T�6�BQ3���ݼ�mn�3�]�$+�ki�٠�5�7��5��Js��j�|Xf�>���z�ڭ�n��0Zi��g0�e�ru� l�9���s�C���iY�-��[�`b�=,3u�I(� {����s�T��mâI�6/c�����`��`{kvo�D(_(JQ�q?[%U9$R��,�~��nE@�X ;Ј' ���~�w$��=,z�5���4�UD�n��"gݼ����6l>�����vm�)ʖ��RM67M��zX%�v_/�-���}{f�s��TIi�<�bχ�'	��ke�E�<p��O&�hn�d�%d��8&!䐎�M�@�q�� ��v�s_D(�����7�ޖ��!̷-̀fn��(Q2��`gs����͛舅�QTw?�Ktɦ��ST݀g��=��V/Vl�����S��7.���m9m�rQ9�ߕ��+zl��v��
��%�%
~y����۪��n��6K�Ձ�՛6(INgs���v�6Ձ�߼}���X��e��69F�=	�����+m<7g:j��������[����J���{u���v�6�(I~���|�u��1�r	dbRM ���ۛj���͛'۵(�	}�U�}�Jr���T�M��v��Z�1z�fϡBS;9�V��v�;�MI��[D�KmX|�Jucޛg;��?nk��$��o~V�N�7T'4�-�Ks`d�v�J!|�%Y�|���Z�1{�В��	$��)|��R��EYU�Y6�p6v��(ƺ��iΫ�Sr8��U��nw��]v6}����w-�^݇����I[b�f%�^k`�hF��:ې{qu����x�[A�l�=�����;�{VU��gZԩY�a�gE�*�6Ƴ��=2-���t�=����!����\q��Z�5�4���+��F�c��k�ƍѺ�;���S1o�����8А�x���L3��wPN[��1imF�Lݶ���[;���خ6���� ~��`{smX�Y��_���z�^��9nFܙ�@��������MY[�`���?nk��)�Vw]R��G��D�4�w�@;�f�}e|�������E��n7���� �n� ������ڰ�"ucޛ�a}qF��Y��@>��@����&yK�=k�%.�r���H4.g��I��3��[*��ҝM��x���h%����e�C�-6T̔�N��v�g3�]�	�_ }e|ٶSQ��k&���d��nI��w�q:���R��Tb"5T� ܓ;��nI>������ڿ�DɽS�M���d�-̀nw; ���ϡ$��v��VV���u�ma��Y��ԛ�����͵`b�f͇�$��*�߾v��~��9nFܙ�@����?��\�_ nw; ������[*�)�����]�Õ�f��n%69C����0^�'���7#q�{����uR�9t�LtH�^��}6��h׶��w�ۚ��!�mJ���{u���{�����j����Z�a�qF��,�JI�^�ܓ�w�7:�HI"VU�FD��!�Da3#U�!�r4!�N}D4F.���Y1Bi� 	��(i�V"��  �!�P� $H�eGQf�P�TJi��:�$�!�A��J/�UT�S��~�C���e3Y��$���nI�u�١ʖ�(��l�M�|�I}	V��yX������h׶hb�ʘ܋)�Ӗ�t��6l�B��������v����fʕT�R�bm�0�.]m�g����-�v�v-3�7��M�:qHق�)?5"��٠^٠r�S���w�@�==����c�I���:p<�� ���L���M�I�I4���z�Ng���־�g�廍6��h��,:'V����`~�ݫJpG���߯��ܓ�����]M\�Sŉ7�=k�>�j�=c�2)V�����r�U��	f8Ӑq�Ǎ.���Kv&��`x�Xv�"6�ٷ6r�׿:�I�/8�R4�F�������r�S@�u������uTȱL��������~H�]��*�����ܥ�6��׏kf��dR�7֮=�q{�z}g��v�0R'����P�w;�����=����uY|���ѩ(��8�rh+k�>�Jv��յ�6��vD(��������ppm��:,�������	wE�e�Mvë�04nW3�UӀy��A[�{m��:�Z;
<�ZP���e�Ӂ���Ӫ���X�[�t;;g�;�:Nى`8]vZ�s:EW�&��m���Q:Q���5�ݱۯF��g�1n*M�-
0�g�WdmtM�f�pu��(<u�[hN9��X�SΝ;�P��Z����y�������SeЭ	��u����r�r�a�ـ�c�I��3yP�B[��K͙��g�m����� ���־�g�廍6�i膙�L�]�	�_��W��M�Ďg}���!���h��π>���:p$t�>�^�{�[[���� ���X��L��@;�f�κ�dY�6�90�=�:p�WNo�\�֮ �&o&G�7J����˸�z���S��ɶ]��vudi����E�.[�8m-�`�r�h\��\��g�w��4ַ��T9�`9n�X�n��-���1����В?=�w_��vtp�Ƥx���,pmǠqrנs����!L���';����;n�S*fH��qǠs�S@�qڴ.Z�=
'+;��՛�S)�uU�#sL�<��Z�u����y���:�u���J=�Kl��b5i^�F�Y|ڂ���	i���|��^����-���I�;7��疏͌����ڰ=�z"~�ŕ�69���sRcH� ������ ��w&���r�>�$��+[����iv�/&E���90�?�I#���Ԓ\�KW�'����m��V�$�-|�K��BH�72b���5%����s��/�I*��Z�K����I��߿5�{욒K�/y�1���I�)�$�_ekRIq����$r�ɩ$�����I/~���('2)�hա�`H���j�r��t�7W׮\��f��fn�ljG�9�Ŏ��IW���$��w&���rZ��$��+Z�J���ѶD���N8��$�[�7ʹ�����䒮�5�$��k����߳?6����.�W�cQ]| ?{���?? ?_��|K����I#�RjI+��|�O��iLX܋�K����$��k��9n��o�~>'�yD0>����^rԽ�Ŏ
EJF�$�-|�G-ܚ�K��j����jI/~����?�V#&���>&ǧ[v���S^UL��6٬j���t�	ٮ�?�����ٛ����{ל����_ʩ�j��w��s�����S#Z�ͪ�� ��}�}�Iu�V�$�-|�G-ܛ���̒%]�k���ƛ[�%]�kRIq�u$���ɩ$�����I.�rƤx���,pmƵ$�-|�G-ܚ�K��j�䗱�w�jI/[�D�1�7�?�I#��5$�3����%��G�$�ܿo��{��߿uv�E�6�s�gs[
l\ծ7H]���6�κ�����{M�!�/Ki�.�z������� �MF�lq������wd�^,�+,9���s��)� ����ut���9��j6(�U��0X�+���/�s�Wu�ݺ��1a���+��ٱi5͎-������ks��h�D\�#[&�nΌ�iׯ4�u���o4_w}����7CYy���بza�j���������l.�i[�5u��9h:i_C:���Is9;W�$�We��_r���$�n�RIw9j���9�H�ōȾ�$��(�$���π9m�3��o�~Ď��OE��n�d��e��=���?nk��J&s:{g��e�"��bk!n��gݼ�Y[�`g��`���	�K�m��i��1����t�'������Y_���+kƞ⺁}L\����l�9㎚��;]�9׉�����P�YN床R�	�p�3����>�*������.�
V�5�M�5�Z�M�9}�k{P����г�M�_����r���&�8�rE#��l�;�}�O�įl�qz������m���H�����D(�[}����,ӹ�`�5�^ݺ�SAN%���U76{����������w����͛t�S4V����vm����ۅ��{��6�%k��;���ۮ:�����9�o�o���׀>��g��$t�=h��N7��(����}��䋝�Ɓm�4��zx�T$���1��G&�t���'{����@pA�VJRJ�,I(�,�K��7��`f��H�<R�I�G�m����}m|�GNxR�����LJ�`~�ͫ�B�(����,̾�o�s����vh�]!� �k�㭜�ًn)C:��3=s���R��h:N�E"kRm�k�>��g��$t��ٟ ����;������r'&���=,f=,ӹ�`�u��!%&a�lk��51c�m�4��z|�D���v��Ł�ڇ�U9t�t!�u��>�� �Z�	����I��	�P��o�ܓ����C�&ƒ�M����k�&z:p�Ӏ>��g����ֵ6,K[͙3��A1��K�������4<����ൻkǬm�4���1��3�Ӏ��s_DB��@��;x��m�	lz���8H��Y_ }-|�c��J&M·�M6�Ӂ5N��������k�&z:p�Ӏ��:Ĉ�M4FG�C�3�b\���.v���B�Q3��va[]"t�UC�hoS|�GN�:p�W�K^�t`m4�!J��]���`�X��
���(̈́��N#K�� WHP��fÁ��ǐ5Ӣ�h�@+��x �"@�9)Q�"F���H! qX)X�B��� �4��W�����?�-$����.�ꪛs2ڙoZ�&�l=��8�f��^��M6G$e��=�6:�#���DkZ�Q�@7mےg���q"�4cj��^���Bz��em)<��i��#��%�&�A�\8خG,�\.�/��^���m��Kp���Юȃ\�FN�.+��k;v��nA�|4�ƫn_5Hm<�'Jr����Mσ!��]��E�q1^Q̺:���܆��C���ʹ���i�u���;k]nbѵ��qX��i���pg�k�	^��c\�Cք�vm��CWS��j\#��βmq��vr��rա9N'\��v6m�`�/-J���m�*��-	�ZV��<�6ֈ��z�O4r�4��E�!nQ���l�g��Z�}V��Z������չ��Kr��ԫl��j�5@�X +���l5H�j��Yk		�j�0ul��㱬v]�����ɭ�/=�%�@�f�y.U���<,g�٨�`-�j���K�ª*��6����Y�<�0-D����z�m��M��[p �[p��f�:(���6���9��)W�E��d36��*�K����L�X�W�����kV� �[M��
��(:U+b��<�<���C&膑�ŻY��*K3�Z!�]�xn��@�YR Xbޫ��`ְm��#�i-΢�J��yi3�'�m[�񝫫��M����n9v��r�.n�[],�0L��i�R�SZ[6��+Qd���0E_i�p�r��W�,`Xt�%�n��v�8�.����Au�ܲ��&�HRZ,�YmC��k�{k��Znǝ��.��*�v��I=6ٱ�����NLI[�l��T�g[.%�+����ڗ���X��i���IH�V���+T;[����l����S�H�U@78Ē���$yn8�:n�����y6�{h۷hW�3l6�YvQ��=�F�#6á�6�����+�MRQdhɆ��pt�
�©�� � ��Q��T��0��p��5�v\�[5k����{t�{i�i�X����˫��x�1%q=mĖ!n��67e�:ڲ抶U4H���L�\O^:�sn9�ͤ�Og����l��^���v�iě�k���jڗey5l��&.�ŗ��&G7��U�,/T���<p��[ϊ�����9�Ia�<	[RuDq�
�3�	;��쉙��W:�7)[+����&Ln�5}�뻻��:��f�/S/n���4CҔ���nNCV�zc)�e�a4!�뮅1Rp䳔ꚕM��n���?nk�ٺ�P���!%���,����S�M�E��� ����k�&z:p�ӿ�~��Ď�{�"��Q1�����>����zGN �־����޷R�%1�n��Q
"qf�n�,���BIL�{���Wt��T�4э�L�$��������L�t�
�D�l��9�% N;.�ƻR%���vĄ��#v��F���{:�H�gN*�UL���v�w]�����#��-�Ɓ�垃dmF'��I�N{�́�\��G{�9��ܓ��4�ۚ��J&Lç�UV�SM�9����〒:p�W�[_��[�'������pGN �����P�Vm�`{���U9t�tP��p�W�[_3�Ӏ�:p%
"=�t�%4�Tȥ��) �L݃�[u��4�M�9���4��M�G#v�n��֧�4V店4U67M�>��`b�=,�t������.���D���1��3�Ӏ�:p�W�[_(���6�M፳L�$�����~�����]�w~�nI��M�;�kSX6�3q1$� ����k�&z:pGN���Z��Ěz���������Ӏ>��{���-�l��ҝr��Ra�x��afw�\FN�<�Va�ضᡮ�D�=8	���Y_ }e|��v5���F��)$4���?$���z�h�e4\�K8��LmF����l��l���3��Ɓ{g��e�dN)"���rh׶h�zX�zXlB��B�$��y��܎�ƞ�M����	���OGN ����+��]�Bi7���ܸc.�[��>���{9zL:K6�\�n9�m�z�h��4��OGN ����+�$�����Mc��1bcn��o�~H9��[g����DD(�7��T:�tKj�Ӗ݀{�����K9BS;���ws�=��5ni�4���v�%;�|X���ۺ�:Q3ټ�b�R���'USMU:j��c���>����y���nI�`�Tb?a��Zɫ5��簒f�	b\z�ύ�wl�ɀvu�ݖ؁/hѳ*��C��k�l�t��WlQ�gQ����˖;Y19U������X�2�=���n6eN�݀���Ͳ�ṗ64�n���	��eSn���v�C���m�!�j�;u���\cu]i�*yT֒Ӭ+�k0�K++�x yIٓ&��Y/W5I3�kZY�>��ˤ���J�di'�f�]ps%�x���(Ts�g��M�q�gL��9��V4-�l�> �����p�Ӏ�WjX���M����W�OK��_GN ���	���y�==m���p�Ӏ>�� �W�J+u���m��4�p�Ӏ>�� �W�I/gh�kSX6�3q1$� ����_$���t���~����0�	��QkP�i�].:nr��;h�nd:]�ӮĎk(���5�ܺLZ������>I{8���[_�n��4�=M��$���%�?%��zX���}��x���ԚX�Z�$���:p���־�^��{�Z���̶X��v��v�3+���$) �=۞�7ı,N�=}�sY���Mk2e�ͧ"X�%�}�fD�Kı>�}�iȖ%�b{�=*n%�bX����iȖ%�bvMt�֦��Y�t��7J/YS��9���%�m���ŠJ�L����q1�fk{�oq��K���6��bX�'�sҦ�X�%�y�{6��bX�%�}�q,K��L�f�Mk3EsX]fND�,Kݹ�Sp�D�K��߳iȖ%�b_���q,K�����"I
HRBЬ�SN��`�S*��
�V%�b^w�ͧ"X�%�}�fD�K(;�P`P`*a����{�6��bX�'}sҦ�X�%�ߎ��ˡ5�d�k��{��7���~�"n%�bX�w���Kı=랕7ı,K�{ٴ�Kİ~�����UI�:-����$)!ff�W�,K���zT�Kı/;�fӑ,K������Kı=��u��j	�mJ�F8�ZW�Q��6�d�Q�׬L����_N7c����<��e�Q�f��w�,K�����Sq,Kļ｛ND�,K���q,K�����RB��<�=r�����f[&�bX�%�}��r�$���C�I���͡"�'~���?� �S[�ow߷���� �|�~oq��%��ߵ���bX�'��m9ı,Ov�Mı,K��m9Ĥ)!fm�,m�l&����d+!I
OȈ��N�߾6��bX�'�\�*n%�bX����iȖ%��<�A"����g�"n%�bX�����B�2�e��a��Kı=۞�7ı,K��ٴ�Kı/��ț�bX�'��m9�7��������7C��T��v��F�^�r���ˌ�SgX���NwFm5��|��䌓0�
k&���>�bX�%�����r%�bX���dMı,K���6��bX�'�sҦ�X�%�ߎ�^5��ոk2�Y��fm9ı,K��2&�X�%��{�ND�,Kݹ�Sq,Kļ｛ND�.�j%�������UI�:6B����$,����~�bX�'�sҦ�X�%�y�{6��bX�%�}�q,K�������ֳZ3Zְ���iȖ%�b{�=*n%�bX����iȖ%�b_wّ7İ?MD����iȖ%�`��G,�S�B�������oq�����r%�bX���dMı,K��m9ı,Ov�Mı,K�;��c}��,�ccsF���ϝ����]�b�v�f��4흫��6w]s�X��z�c#��c�i��a��n�9���b��W��q�5�т2M��.�66� `G��4냬�����.������U+n)�[�q���8�(v�1ݗv�N�3�wm�n�]����>e��[W�v�w���j��z�ۛl�j��v�Nt��3W34�2�5r�B���C,ٲ�[�[X�q��N���Nlzv�ݥ�����'`g��nf]\����h:kS_�w��bX�%��ّ7ı,N����Kı=۞�?�r&�X�%���w�
HRB��Zr�ܺrS	)���q,K��{�ND�,K���Sq,Kļ���ND�,K��l�d)!I
H[���mQT�H'MMfND�,K���Sq,Kļ���ND��
'� ș���2&�X�%�����ND�,K�k��]f��YiMdֵ���X�%�y�{6��bX�%��̉��%�bw���"X�%�������%�bw�;�S.��Z�j�˙�ND�,K��fD�Kİ��E�����ӱ,K��������%�b^{�ͧ"X�%������\�ˬ#v��Ιx�R�q �5�m)��0je:�]@�pF�B���kY�7ı,N����Kı=۞�7ı,K�{ٴ�Kı/�����$)!I����R���'ST�7�6��bX�'�sҦ��`k��#`|�T� ���%�s���ӑ,KĽ��ț�bX�'{�p�r'�(��j%��I����T�m�N�e�aY
HRB������B�,K��̉��?�Tj&�{���iȖ%�b~��Ҧ�X�%���v�\�h��-3Y�3Y�ND�,�TX�����q,K�����ӑ,K��nzT�Kı/;�fӑ,JB�f�r�ܵMSD�i�l�d)!X�'��m9ı,N��Mı,K��m9ı,K���q,C{����}��c킢x+rsM/-�a!F���2��֗u]M�Ӝ�v��M2�����|���55���au�q>�bX�'�s����%�b^w�ͧ"X�%�~��"n%�bX�}�p�r%�bX��]�j�4M�Jk&���7ı,KϽ��r%�bX��{2&�X�%���ߦӑ,K��nzT�O���j%�ޙ���К唊k��{��7������2&�X�%���ߦӑ,b�N�1"�R�(2��E!(�
*H��JB��Z*RД""�H4� �@�de �	$��% �#T��iV�RRHP-"�V�Ow�u�6!T��)��
B3A��±�+))F���������1U�D��jE��U���%���� D�`�4MP���y N(� �G�)�����@�"�yz����O�sҦ�X�%�}��6��bX����N�]t�i�6B����$/{/KND�,K���Sq,Kļ��ͧ"X��D������q,K�����3T��]B��5��iȖ%�bw�=*n%�bX��{ٴ�Kı/��dMı,K��ND�,K�	w�ҩ���T�!6�%SCCnS'a�Sm1�KӧU�:ۗj��u`6kr�՚��j��S�,KĿw���r%�bX��{2&�X�%�������U/bdK��������%�b{����d�]�Z*�����{��7��}�[��X�%�����"X�%�������%�b^}�fӑ,K��}�.�E5M-�����$)!{3+ND�,K���Sq,+D�K��߳iȖ%�b^���q,K�����fj�f�氺�6��bY��D���J��bX�%���ٴ�Kı/��dMı,< -Ȟ���p���$)!x+5�Ӡ�܊SeUd���%�b^{�ͧ"X�%��*�w��Ȝ�bX�'���6��bR��%�0��$)!IpyUU�:R�8�AB�E�\��`yjۂ��y��z�nih8�-á5�)W�w���ou�~��"n%�bX��}�iȖ%�bw�=*n%�bX����iȖ%�n��}��ғ�Lk��������D����!�����\��,O߮J��bX�%�����r%�bX��{2&�X�%����s5K�e�-�3Y�6��bX�'{sҦ�X�%�y���ND�������fD�KıY�ߕ��B���Q�lT��۪)֭̕7ĳ�D j&���ٴ�Kı/~̉��%�b}�}�iȖ%�bw�=*n%�bX�w۶�殝S�"�lr۸_�RB���ۭ���ı,?������%�bX���Ҧ�X�%�y���ND�,K(�Qp��Q���\?ư��䰆�d�u��2���)ۣ�����ڻt���1�;n���gջ,�3�Ս�b��fLp�����m[U:|�<[�nέ"m�ĝ�4Ne���\%����Τ��d:5����P�R:A��l�M!�q��&�o*�k>Mۃe�77\�"=�\�{�����jtI�>�����fj�L���-��N�-ƞ�������A04<�vIvDfr..-���`�ڋ�N%-��RwB*l��i�̉�Kı>�p�r%�bX���J��bX�%���l?	>����$)���VB����ڟt��UM�\��a��Kı;۞�7ı,KϽ��r%�bX��{2&�X�%�����"X�%��5�f��SVfXS2kZ�Sq,Kļ��ͧ"X�%�~��"n%�� a�������"X�%��\�*n%�bX�|gu��sR5M�S�黅��$)?����Y��Mı,K���ND�,K���Sq,Kļ｛ND�,K���T�U.�:r4�!Y
HRB��7��Kİ�QH���ND�,K��߳iȖ%�b_��ț�bX�=�������+�*%ݮlt���b���ܜ/(j�T�S�˵��2uv�튓��pQ���iȖ%�bw�=*n%�bX����iȖ%�b_�����MD�$����\/�)!I
E���N]��Y�[�*n%�bX����i�`&��<U�q9ľ��ț�bX�'~��iȖ%�bw�=*n*HRB�n�N����-����n�~ı,K���q,K�����"X�*�MD��~�7ı,K��s�_�RB����X�)t�3-���q,K?*�Ȣ�Ȟ����ӑ,K��������%�b^w�ͧ"X�%�~��"n%�bX�����CZ��\�Y�ӑ,K��nzT�Kı/;�fӑ,KĿ{ّ7ı,O��p�r%�bX��t�JkZ	�6�j�Ӻa�.��kv�P'ԝ��c�v���7l�����������FrE�Y[	Ȗ%�b_���m9ı,K���q,K�������&�X�'�s�=�7���{��������Bk�V)�iȖ%�b_��ț�� ��j%��{��"X�%��\�*n%�bX����iȟ�����g����kW5	��0ˬț�bX�'}��6��bX�'{sҦ�X��@~Qtn&�]o�ͧ"X�%�~��"n%�bX�~���R�Yus��ND�,K���Sq,Kļ｛ND�,K��fD�Kı>�}�iȖ%�E���NZt�M���Ʌd)!I
D�｛ND�,K�*��~̉Ȗ%�bw���iȖ%�bw�=*n$���$/������N���0����L݃���;��#m�nuY��&���6���t�Kn[lR���B�
HRB��vdMı,K���6��bX�'{sҦ�X�%�y�{6��bX�'{�I鸛��WS[��{��7������m9�H�&�X���Ҧ�X�%�~��ٴ�Kı/��dMı,K�3���f��fh�k��iȖ%�bw�=*n%�bX����iȖ%�b_��ț�bX�'��m9Ļ�n��?�dg$[qՕ������� �DF�D����ͧ"X�%�}���q,K�����"X�@^�QN�G�U6.�M�%��J���oq��z���К敊k��x�,K��fD�Kı>�w��Kı;۞�7ı,K��ٴ�T���$,��p0������rˢ^V��<lr �gq�.vjB���=Xi�n������T�T���Ӛl�����$-����r%�bX���J��bX�%�}��r%�bX��{2&�X�%���{��.��P�Y332m9ı,N��Mı,K��m9ı,K���q,K���ߦӑ,K��d��sͺ�
ǻ���oq����߶ӑ,KĿ{ّ7��	�4ș߿o�m9ı,O߮J��d)!I3nM���t�bt�書_�Sı/��dMı,K��~�ND�,K���Sq,Kļ｛ND��oq�߿�Ԟ�帻u5��7�ı,O���m9ı,?��D+������Kı/fӑ,KĿ{ّ7ı,J��J�(�"dB S���&�����&��j܍F�m	�-�&�ͺ9�V]��9�9��v�A���es�wu9�N�:D���1"�k���ե�����"I,$�*������-Y��1�{p�\3��ٲ��<��nB*�Mx�K�*��I�d�F�q��<��^�6{��V��@P���;Yl�H*��ĝl[ٞϱҭ������;���˗����r��]Lww�{���\|��\V�dy�˭��a�M�����+ָq�݇\�����kY�+���Y>O�,K��nJ��bX�%�}��r%�bX��k�C�g"j%�bw����Kİ|k߳WX]��dֵ���X�%�y�{6���:���%��~ʛ�bX�'}���ND�,K���Sq,K���~?yt=9�b������{��7��}}�7ı,O���m9ı,N��Mı,K��m9ı,��n�:�t!ӑ�-��d)!I
H^̽�ND�,K���Sq,Kļ｛ND�,K��{*n%�bX�~���R�Yus�̛ND�,K���Sq,Kļ｛ND�,K��{*n%�bX�w���r%�bX������7R>H�`�٥�\N�`m��\M*=��j���;�Nj���4���̜.��7ı,K��ٴ�Kı/�ײ��X�%��{�M�"X�%�������$)!I3nM��n�6�����r%�bX��k�Sp�`]D�K����r%�bX�v�Mı,K��m9ı,N�=��3Y�Z�5%��ffT�Kı>�}ͧ"X�%�������%�b^w�ͧ"X�%�~���7ı,Ot��.f�Mfa\�Y�ND�,��{��Mı,K��߳iȖ%�b_��eMı,K����r%�bX=5�f���YiLɭk%Mı,K��m9ı,K��쩸�%�b}���ND�,K���Sq,K����?~�e�Xed�
3 -ruJ=2pnv�j݄��͍u�{�W/k�n����±M~{���d�,K����7ı,O��siȖ%�bw�=(m6	"s��&��*��RuR�C�#N[r���{���OD�,N��Mı,K��m9ı,K��쩸�%�bu���K�eԶ�%��m9ı,N��Mı,K��m9�~ �+�6H��{�{*n%�bX�{�������{��7���7ߝe�h�+T�Kı/>��iȖ%�b_��eMı,K﻿M�"X��Bݛ�aY
HRB�o\�I��tjk3&]fm9ı,K��쩸�%�b}�w��Kı;۞�7ı,KϽ��r%�bX��]-Ԛ�׋�n�8�ẑ}	�O���֊M�\6Hؠ۪:m�����"#`n��w��7��b}�w��Kı;۞�7ı,KϽ��r%�bX��k�Sq,K=��}����iNj��-�{�7���%�������%�b^}�fӑ,KĿ{^ʛ�bX�'�w~�ND�.����߲6�uel{�oq��K��{6��bX�%���T�Kı>����r%�bX���J��bX�'��w�٫�5u��k.f�6��bY�@�Mw��eMı,K���M�"X�%�������%����T|$5������ND�,Kӿ��њ��Bf��2�eMı,K﻿M�"X�%�������%�b^}�fӑ,KĿ{^ʛ�bX�'�>���%izEmc��.X��":s���mf�OkW�X�����=�N8Yx�V�����%�bw�=*n%�bX��{ٴ�Kı/�ײ��9Q,K���M�#���ow��k�YgMЅc��x�,K��{6��bX�%���T�Kı>����r%�bX���J�������ۓi2��N���w�%�b_��eMı,K﻿M�"X�a����\�*n%�bX�����{�{��7����߿=-8�܍�P��bX�'�w~�ND�,K���Sq,Kļ��ͧ"X�%�~�����{��7�����~�)�\u���ӑ,K��nzT�Kı/>��iȖ%�b_��eMı,K﻿M�"X�%��;�FW�#�`�H��X���$B0H�	"@�%��wM���	Yg�>cH�FE(����h"���*u����P6��0������(j	4��]��le	P� X���"7Ph�+tЌ��a�HG��<��)";�}~~�� ����{Lplgq�mS�LFɴnZsO5U�&Y.��X�^��=QK�;��A,!L�9�N�Ѹ:�r��X�UUM��66UCm�ι�3f�W��[8�ˣ�j.ebg��Z^� ���*�wN�Fz=��T��$m�8�d��$5���u�Rn����÷s��q�4K�p�p7�M����|��Ή�n���h��kj����ݶ6\�۴�u�V���
��V��m��Q�B��vL�G�����%�[�,vQ�nѯm�z�;�z{v��p�.P�Jo��|��y�z�Utۄ��k���!�eDu�I�e�4�ɷe��g3�\��%O;������r���lVtݵ��67���:%3�3+P �k�R�h;Q�Ѕ*n�����;��R��ԫv� ��q66��)�n'F�[�]��R�T������κ������Yȳq�Ö�p�gs�S��R�&C��E��*�ʵUF�����4;�HX`�Q�������Z]���Uj��T��AX۪6 ����
7B�st���y	6���' H�w 耶�rt��𶅴��u�p H�)]�HUK�J���e�a��Aa����h�+J�Ya3�D�PS��m��6�ˤ �[���ώ�E��i��\���ɚ�ge�騯ӎ̹�.��unm��È���"x���<nMظJ�pr[3f+[9�2�ʅ+n2�ij^[�H��*CH�}�]ʪ<a�l�۔�k-�ι�\c*�բ����@�Π�C��ӱ.�,�cp��jRX�I��t(�83�v�%���Sj���av)'�Z��%;�A	�vY�vmQm�䏟|G?2��X#F�[wK������l�[��V��r�2�&�"�m=� �D��砤�fu��|���Z��V-�0��0a6�n; oVt�^��5BIOF�νl����ɹ�9]	��XK,��L�5�" �� �N#�? �6
�CH��J����lJ��_ ���B?���]s�=d�ƭt���q���9�'Xmmf-t�:p�ϛ����t`��<\#���v��.8^�v��l��X�23e�vAub�{t�<q�O�Z��2Ѡ�����b���\8dt%��scc�6�d���㪙�m���A����8� �i6Ϯ���Q�ggT$q����.vQr=vy9=5����m��Q�m�;������L�鶑�vr��	���ϳ��C�W��v�ʼ�d�Mo�������SL*i�R��UL�_��$)!Oݿfӑ,KĿ{^ʛ�bX�'�w~�ND�,K���Sq,K����ϼ7C2�5�������oq���ʛ�bX�'�w~�ND�,K���Sq,Kļ��ͧ"�T�Lҙ
E}����ЇNF������bX����M�"X�%�������%�b^}�fӑ,KĿ{^ʛ�bX�'_���Z�k&�s%�fM�"X�%�������%�b^}�fӑ,KĿ{^ʛ�bX�@��������{��7���������*y�
ǻq,Kļ��ͧ"X�%�~���7ı,O���6��bX�'{sҥ���$)!g���T�XT���������:O5��X�gr��=�ƂB䢸:��OY�g�ա�����7���{����{�ı,O���6��bX�'{sҦ�X�%�y���ND�,K���3C�n�ST�i�����$)!{�z\����PO
*������?�Mı,K���ٴ�Kı/���VB�������6������ju��ND�,K���Sq,Kļ��ͧ"X�%�~��"n%�bX�}����B���Q��]KpU9t�6UVJ��bY�T�����m9ı,K�߳"n%�bX�}��m9İ?�&�{��Mı,K�Oo�n�֦�ֵ�3Y�ND�,K��fD�Kı>����r%�bX���J��bX�%���m9ı,O���:�`��an��3�NcZ��[RqgK]�lXe�y̰��󊗦��c]ow��2X�'�w~�ND�,K���Sq,Kļ��͇�O�j%�b^���q,K���n�)u�֋��j]fd�r%�bX���J���GQ5Ŀw���r%�bX���fD�Kı>����~!I
HRB���N��[�SsS/%Mı,K��{6��bX�%��̉��8�i�HDSjP�(�P(U!��Q7����ND�,K������%�b}�nM��r�:TSlsM�/�)!I�!}�=���q,K������ND�,K���Sq,Kļ｛ND��7�����OKL�x����{��ı>�w��Kİ�#�]��9ı,K��~ͧ"X�%�~��"|��{��7�����>�D�=��4�+�qHr����c�9��pK]v����4OϾɯ�-9�A�nVߞ����oq��~�����%�b^w�ͧ"X�%�~��"n%�bX�w���r%�bX��^�%{,O=Y[��oq�����~�NC���j%�{�dMı,K���M�"X�%�������%�bt��~}�Ac4�S_=ߛ�oq���}�q,K���ߦӑ,���j'�\�*n%�bX��~��ND�,K"=�uT�9)m�Ht�
�RB��Q;�s��r%�bX��s����%�b^{�ͧ"X��8��yD�D潼ț�bX�'�ww�.���sZ�K��6��bX�'�sҦ�X�%��}����}ı,K�߳"n%�bX��w��Kı=�}.����]m]�[��n˪�0��mV6�3����9�Z�<X3m�sn��E��{�o%�b^{�ͧ"X�%�~��"n%�bX��w��Kı;۞�77���{�~��b)�sV��{�2X�%�~��"nȁD�K���M�"X�%��\�*n%�bX���w��	DT¢��z�t�S���E��3Y�7ı,N���6��bX�'{sҦ�X�"�Q5��߳iȔ�$)!Nw6B����$/h�6��5s-2kkY6��bX�'{sҦ�X�%�y�{6��bX�%��̉��%�b}���iȖ%�bvM{٫�I�e֍�Z�J��bX�%�}��r%�bX w��Ȝ�bX�'}���ND�,K���Sq,KĊ{�>���ۅ�p��ݦ;XÌ
��<��i޷l95��кk��pI�Ք|��ƌ�syrkr�lsqۮnV�\��=�nɰ��M��2Sq7Y�k�T�Y�1��%�pnm��i�S��+��f�X
:����k1�����݇��V��m�y�7m�4��ev�ܦ@;����=k��C&�G�Ί���{9ZeZKj �n��u�7/N���wwoV�+�ݧi��ƭp-u<u��x�ۧ�M�諭7������p ��R)����{��7����ț�bX�'���6��bX�'{sҦ�X�%�y�{6��bX���߿�AQ���w��7���'���6����"\��,O߮J��bX�%�����r%�bX��k�Sq,K���w|R�Y�\���s3&ӑ,K��nzT�Kı/=�fӑ,KĿ{^ʛ�bX�'{��m8B�������SCn��ۙl�Wı,K�{ٴ�Kı/�ײ��X�%���~�ND�,��Id.���0��$)!I�����楱jkY�5�ͧ"X�%�~���7ı,N����r%�bX���J��bX�%���r%�bX�;�ɬ��K���+ng��br.�HJ[�lj.uJ�^��J�ێ��ѹ����s�~�O�Ϻı;���iȖ%�bw�=*n%�bX����iȖ%�b_��eMı�7����d�qI�nV�=ߛ�o%������b"�xC� ��Mı/w��m9ı,K����7ı,N����r%�bX��^�j�kYu�Fdֵ���X�%�y�{6��bX�%���T�Kı;���iȖ%�bw�=*n%�bX�>;���k,ֳZ�r�fӑ,K? �D�k�T�Kı=�o��r%�bX���J��bX�%�}��r%�bX�{�ִf�ۖ�e�2�eMı,K��~�ND�,K���Sq,Kļ｛ND�,K��{*n%�bX����K-�-T������lY��ɶxCV�Z��/FM'�6_\p��J�V���!I
H��zX��v�s_(���C6��a呹���I"N�m�����Ӏ����kj�kխ�����7`�5��zY�+Q�Z���~3>�wΜ���բ�i����3M6۰�%;�|X���ۺ���4Ѯ��i��B2Lm�@�������W�I8���{Cz�:�u�×[Z��Dg��S�%8�c�ݴ>��o�{���ϒWdey���������3�{�/,{��u'�M-z���Y_$t�'�)�[f������dJBcȤ�f=,�=,�)�������~�{ssu�1-l��8	#� }m}$��}������F0�!��4�+3���c٪SM�)mә�p���Y_�8	����ىG�#o���`�cE1����U5���pvӬ��FygZkUո�;�ﾕ}�y*�ب��7M�>��K=�K �Z�	��V4ŭ���lm��zGM�즀}�f�}{f�~Ď�j��m�0F9��h�x��l��3?$s��@�Ɓގ�Ԙ4�X�p����>��ގ��t�=���n�I4$�ׯ[|����Ӏ�c��?nk�1d(�(�(P�M"���]��Wf�n��,��l�
ܻ'0���e���1��v��0��h��T��]9�f�q�F�m�1�Z���[���ђ��u�N]V(v� ev�ɶ�n�i]�箶�c���Pt�A���G7o��n�����2 �g��v۩^��q�kms9�+r�J���`�g�ݵ�-;��Ț���cp���u���r"A� �%�\D$����W����o�1�qen1@�D�'����f�K+��eЗh�K��[�<�U�������8	���Y_ }e|�z=����U-�M���c���	D�{���{����ǥ�B�9n��UM�H�nf����π>��z:pGNE��2\Զ*&��T݇СD(Jgݼ��|X�zXr��o;s�I�t6Q*e��n��c���$�v����z��hp�.�4�5&)��cg��l%��sкq�8�T�8�/Wa���FV���k1<ԙ�*0���>�0=��8xR���4���$�s��n�<*#�>FnL����{�S@�{)������Y�I��c��M� �w;=�K3��s]���Ků��c��$t�$����h�٠s�UǉH�6��$e���K��>�������zXo���jl��ǣTչ6bK��[�[;�+K��m7noU�s)�]\��n�R�u��>�� ���	#�$t�=�!��kf#Si�� }m|����ǥ�~��|�L���&�9	S-��v�,�zY��B���ZDJE	[����i��4����I�5� h�����:��mVNy����B%�F,"H���F0�!���8 mD� H N
��P$ �h� @�$$���c�  ����
�
�(��hD�B�h+
$B�
hhƐHE�0�J�
	U-	U� 8(��,	U��h�%t���D,ĀI����I����`�H�%HU X0#H"mJ E�+(@b0 FI-J��4��#"���BV$5��t�+�x�nhM@��G�����W�
<"�Ғ!@�����<�  ʇ,ޭ|=k�&TJ���&�5�$���;�|X�����vf=,��I�N5����}m��~��{��-�Ɓ��S@ⶡ	̉�c\-D ��R#����%	�q���<ڕ*�81ɉ4䍹qE$���@�q�`fc���@�w;0�T�*��i��o��:pGN ����k�Q�
Q����2���j[l�=�O�@>�� ��4�����l3[�jKu��>�� ���	#�r��B�$�A�HD D�"D�"A�Ҕ�!h`.�4E��A�AH�b�@""[	l/Ϊ��3j{J-�m�Km�����@����m�m�4�l�?�%Ć���L��QNd�}9�F�e��d�9:��]���-=t�77[M����Ӏ>�� ���	���n���F'�&pGN�(�2��`��`fc�����[�jkq,OL����>��H��I8	���n�M��z�O[|�s]���K=�K�3��va�\�7�u�Bǭ�H��OGN ��ܒs��nI��X!E`�����w�����Y��+��v�6.�[T���i	rk�D�:�Q� ��i�S��Լ^rF��*��;rj9$�2qtU�."�`���3�Fnt�s��T�:a�C�ڕ;wj�f���+�,�G[n�1�팖���۵��,]Ra�v��A�"����w�|ݷv�|������֭-Y��ݲ� q�Rvd��$���c2�.�)�����BI/%J�M���,�5u����c�k�Tힲء"���:����g����$�拞[(�Uo������ }m|���GN�S��2d�y$R��o��bA�_M���z:p�e�3[z��km4��ۚ��zY�"IL�k��=����UmX�6�In�6��$���t����>��eD�k�oq/��I��t����>����m��q���v������n#;f��q#��.�ڣ���9ۡ,Ɔd��N�vݞ4��K_ }�_�8z:p=���Z�i&�&�M�޵�߲f~� <��]K����>���$�m�8Uu����q�"�h�e4	���K_ }e|��R��I��$�6��OGN ����+�$��.v�S&I�A�!�[f�}e|�Ӏ�������V-�׸8E��9r6�Ғs\�m�ӹ\ۊ�v�]:l�N��**�2������\�Ӏ������ʭ��ִ�wu���$t�'�� }m|���*%I�����x�g=��N{��� ��X�P:4��߻������H+Z��	�1�OL����>��H��OGNg3��M<�%ܒ94��4ff~���/l�v٠\�&��&LY�NIɵ3��Ƴ)s ��e��v+�˔��4�F%��mn7��OSBǭ��:p�Ӏ>�� ���<
\�I4�!'����:p���Ҿ�:p�)��x���6����K_ _J�H��_GN�l��ko[x�m��� ����Ӏ���~��fB`�*��Ny ~�z��rN{^կ#�m�
A�&���S@���n������^v��f*��I��9�(��F��ڹq��S�\ه/Sô�6�cC�Ǎ6�ƿ9��h�����@9{g����@���ȌoƓ8�k�%|�Ӏ����dw7V�m4���J�	#��ye4�l�9��ֲL���,o��:p�Ӏ>�� �W�{��K��&���m���������k�31�`zV��D/%�R)?]�W=aE#-�u�/$�g'<f�Zy�3�N �;W/k�&s��Z�s��s�f�2Pv�nL��xl�[-uhX�̭I`��������v� ���A.�[K:���8�3Ou�uR��&�^2�����
h��m��Ý��uڶ���t�*u�T��sj�<����V�.-���[r4�>C��7U�d5���\�>z*q6rJr��κڌ7[��$�&s�v�׷Eq�F��R�4���G���r�6���y��k�31��(�����3jw��޶��M&��W�I8	�)�[f��X��<���Ф�X���3����D$�Ows���`J-�&�n���OL�'�� }m|}k�$���k[ź�1,OL����/�|�Ӏ�:q���~��v-�����jn�z�����t�*�ng�V�m�̃sCHv�5mB��`��`fc���ǧ%�@�w;.�M��St�:n��ǥ�P�"�P�$�b.����{u��5���R��M�Ǻ٭�p�Ӏ>�� �W�I8I����ǯ�h[�������H��_WN�l��ko[l�m��� �W�zGN��p���\�銳Z�؝ӵ���.�M$��e��\�80���ժ!�{7�`�Ʊ��ă[m��Ӏ���������[*M`�k���I��t����,���S@�vƤ�)$X��m�@>�I'��s|�E����g&���3��ի{�I6�o�/�|�t�/�� }-|��/��i6���zGN�:p�����6߿�x﨏���꧝��ZW�"��ܛg��;d��5;]'9�^���������gdt����/�|�t�;Ϋ�,QHӋcJC@>�}������vn�,�zXʜ�C%�M�N��4݀o�]��ǥ��B���ƀr��@�,eyG#X�)v	%��Łۯ� ����R�^Q�%
���ҧ6�YS5C
<I3��:p���־�:p�o��������:6��bN��p��u�1X�e��)�q���m��I\�I�7US,�n� �f�ُN��C�_�Z�L�)���T�t݀nf��J�3u�`vs��?f�<��h��I�аI��:pWN �Z��_?{#�bm�c5�6��Y]8�k�%|�t�=鷛��޺�tT�e�~��`OD(Uۼ�mt�'y��ܓ�D���*+�Т
���D�����(����
���

���(��(���U��(*+�*+�* ���PTV����AQ_�QE�D��TW�TAQ_�QE�D�D���d�Mg�ѣ��f�A@��̟\���      �        ƀ    �D�	
PR@*��
  � 	*� ���( P� $��E	� $()RH0    
  @Ud5A� � �C@� ��p  � D;���oK��ۦ�>�yz\v�m�������R���s�2�S������t��J� ����������T��  � 
$(   ��ϩ}�o��W|�:]��^����� {ʯ������L�sq�]}�M�80      _{�U� ��m�K�/��ˬﳥ{� t�[�)��OT�jF;��� x} (�J�E �V@�>�W3�׳�׭9=u������Δ���ӓ����{�r��٦ j�����޺���n�_]��]�} zz\[�oy�y�f���޽�� �s�9>����woV�ܪ���P B�  �@N}�[�;���:ӓN���4w�M����۵i�Ξ�o�OK��/��_m�����w�����������x ��m��s�9�]�>�׶Ͼ O���������js����׶��<>� (���
	� 4�魯3��m��y{�z}�x� �r��w�<� ��@ Q@1h@   }`P@ � :;�JX��JP�� ��dQ�'M D ��R� ��=�R�5 h�T��56T�T�@h2d1Ǫ�*��!�b�=��Q�*��db41?�%�)T� ��&Ҕ��2�☔-�_���_���(����t���[;[z�kkq�@����D�D?�
���D�uTV 
 ����Ʀ
��	����"�0O���<�x���ÄT�ۓIxQ Д���	��K��.n���������c����0�4�\e�Bn2����r��7BV��e��%�i���5H0 ��FD���t�]F��O�K���f��\�ƾ<%ͼa!L#L��p�K��K�0(f�H1+X��RN��ML�(:�P[s�_� ��zy��<�9�=�&)��OD W��'�5!Hc��99�����D�3���s`H�E�����\��z���� Ĉ�!bK��X1�F$!p��~Oe�u8xxH��.�l�0�1J�] �xJiOH��6�%�
���i��u\.JB�b¸i��T8��4<M��(>�^Jbx�aG8�B���Y)�ӟ�?$8z�8xBHA3! �E!p�	$S(���H�$.D� "4�2H��5�s$X�F���I$ A��@��)�,��#RS5�a�Mfyuċ$�˙9�T[��s���P� _wջ�~�\��? x1h�J*@�t�������|�)fs�@�@���k��L.��0�M(B;y�xC�U0���3|�xT��4�OΞ�Xz�4�������[�$n�)Ļ�����<LhB�CC`XP�K�\�'��~!��~Ҟ�bF�!��~=/	Q��%9�e�JKo��D�^s@!�p9���+ą0֤F����}�����|�~����S5�B$p�cZa�s� ����c����t��_XY�8V7R]p�X�4�yObąRzᐱ�J���`S�$#P�pʘX���
�Fe�b�,!$���z^va�?~��i������U#W�"v40<N! ĽG���I�ƕF-�	FR���!,��#,U`хj2F���,�B�@J$���*�,!%;�N�lFE� ������?߱ku�i}�۠6�rl��7yr�w{5z�T���V�-��z�����]��o�w��^H��=	����X@lg���K����Ll-�R�)H�n疆�$B��L	%H��bA���xĠ`�*�&1�Ċ����H�R�J�1h�j��01t-�P��qcC4 �LF�	T08B�!LB�@"�M9�d���Ja��B�F"P���cLV|cS-M��ҕ�(B���Ą�$��2�HJ��0HF��	#���!
F��2�#M�s�7�2/�8SXi�A�p���
>O�)��,吩��0�pӁ �����p�$)\�F����Ȳ>�Ó%�aZ92Y���e�h��p�៦f�0�x�� �*�o	���l�?B~jB� Ӟp��!&A��G�������|I��O&C2XT�p#\!L�%<�2!H1"�`�5!�YaV���y��9��CY�=2���+�G � "�D`�B�K*��,��I#�Y-���FOh@��-!C1��Sd��r&�-�	i-�����V��XR�lI.m��l	0���!F4��!Lr�NI�Ȓqu9B�mc �a �r�HM���$� xFɁ�������H�%q��R[P�dБ4J�!J�*��Q,�cS6�R�aH�S �e��I �đ<����)���m�D�J`�@8�*� 0
��<�pX1����C��k�
]�A ��<�d�5��x��빼<c	5)}������`��1�$�S�!*A�� �D!��H�0� �IBDMV#B-T @ ��A QpS�<	k��Bo!d�&T�7�#
F����$dΞf��<w��C�����^8�aD �Ƌ
^<�8<��aP�B�'� BSH��Pp 4�y�3��/�d��ǆ�g�(�c��J�����4�g�
B2���&q��@��ܾy�i��$�i�!_�G쉨�G�c_��_�9�`S!��`�2,������� ����°�`�� �! �G^P�L0MB6^�8>!
����0�U�<B!P��v�,l#�� H���U��"W�Zf���lk�$J�֑1`%�%�hd+��+��B�]i���JƘHHA��$H"HB�� �"���H�2�!�,
,+�p��I0 �a�hU>ni,.	�%1�5N3��� o��03�<�~�)XFgB������4���I%�����o��p>�R�"0)&���`z ~6�\|�t�{��W���HWW"B,�O |�B4p�|�_��S��\8鯄�
�ZH0P�(�*�bJ5y�מ[B�=��x�:m���a�P��	G�
v�(��8�����p��F��y�9���a�J~-�{
���BD�����졇�Sy�hSOB��9�O!s�=���!��+�~U����
�bR
�h'y�W<Y����.�+]�������(\�)�L�F�&�g$�*��s��q?�����vČX-�<I�:C��$O��̦�"@����54�=����1xm*�Z��?F�矋��$�
HL5�{kfԛC|�'D4<_'�\����CE���O���1�!��xv�K�P���pd�2@�p�2M�)�2�9�Ya2\q$�3�i"pGO	dxH?��CbBB�a�]n@�����ș��ݜ�B{�5�?D�k��I)��qJ!�eƄKC>/`�<�?��b�HE����0�!Q�cd�O<�e�"��|��:y�y���"�2fq���Ђqh�3��ce�N9�inQ�$2��'��i�@ �O�����	 �%| c\5�͒\`�X�H�Z�	��c���
�?�CB�xC�,�,�w�l��Bm�9���aX%)�����)W�<)e�^��S	%3�VAH��cC�7,.f��!!�1�1cK4�c�d0dn�Ŧi��C�!d���q�<��8�"8�&��Bƾ1Zc)��6��&�)Z�Z�B���"��X�M	BT�%j���Xxs������H1
�!�5 S1���� ���Z�R-#�j��k�A*d�������q��o�Y# H�	$bc#�R)XE=|P��?-��c ��?1*@�d)��jd$�H�)B����0bE�D�HH1"E�*D�c�lH0I�H${�;�ӻ�����  � 8  vɺv�&��ۇ�lX��K�v{Tgn���<v2X�T��[�Z�*	īj���sl�^-�!�`:mw	km��%�8��2�*�����Q�ʪ���Be(l��2KJ�P���������Fv+�;0*�D�WWR��*�TY�Ԡ.$�L�֑Pu5�H\�&hM��s��U@\Q@�F���e�$�i��L���ҬUR9���2iV���U+UJ��v�V�j��Fh,u5M�*�1����v H�v�[Khs�h2p-�\�;RA�Z�S'=��ڪ2+��m��nu�g$ �@�H�j�v�mo���|     8Ԇ٤ٶɝ@      	      XI��  �  �   �-� �e�']��v�i�q���Ens�j���f0�Oi�Q*���� mJ �T�v�`s�֘ � ַ�����V��h��$�i���l
���m���5W*�*�+`�ִ  ��l��6���*�kX8�m�+��;.�*�W����n  m�    ,ݫ$Z�B�:��$ٔ�oP	�V�A���E��D�mm�E�落o���\^��U���We�bcl��   ���c�3m��B�k�l��l�kq1TxA�P��[N�q�0T�.Y���ךL:�[�:b�������� -�u�f��a�J-�X��֤�9յAmĆ���T�[[m��G��}V��l8��1 �[���p�H$˦�mS�`mn흀[Kn�7���v�m�7n^Wx��Uz�0�[7Y��` ��[;K�P#;;l�5UF�g�+�����e��m�� -�g� Z+e�eZ�m���5m�[%� ���`�� H���Աv�  6��np-�ȑ*��[Q�jzu�VQ���6�`��b�V� W���ue9{[m��-n�V��Cv흶v�� m��H:�� ��Ѷ��[Am-���@ m�Z��u[�m�� -�l� �c��R[vݪU5% ���Y��kzn���)� id���m�v�	 �om��     rC�Y�l�m�kI���`� ���   $H �m����6�c�Fδ$$ -����u�&� m&�k  �   ��e9 ��}�m� �m���i$�85���p��j@ ;n^�[NO�����l�`kpG}����+sv�]����`[@H �,���� ��n�4��
��l�u@+,��@UJN3*�< Ur�`Լ�԰mpW,��R�3p�[WJ���S�7l����9@-�֋��[l �i&���6��^��� �e��  6�cm�e�sUj4���Fl��.   ݭ��i0���� 4���� 	Km�m��    }o�| [@  � ����5\���[p�  lE�6Ƶ���i6H�`�J �[II�	D�hK$���˦����`����x����'\��])�˱*Ҭ�p���  �����_Iz��mz�M���$��@�mT@�'g���Z�R�ʐ�  e���^h
�]�l]�[o6�l䄇�m   
Y  mX�	 �c��`��������}�m�6�6��Sa%���$����P�5� �N� �6݁���  �m�m  ���L���  m���I�m�����T[i�4���U�WTۭ����]�Um����� �b�)�m�BD��	e l��`�[���J�!� ��om��H  %��҉��M�`���Kif��-��-�8 m� 6�m�@� 8          h-�@m�   8       $ ��p  6�  ��l YxB��Z�`b��Z�V��c���j�����0�I���-�[d���۶඄�-� ��m�wm%ٶ �  @v�%m嵮�3Nݵ���� $l�jN�K,��  �8$T��nt�$� 5��m��M�� �`  6� �6��4P �(n͚.��wZŲQ 8-�H�� ���S�m��D�Z��j�zU.�^c$�U�ibke�@ 8�n�r�� 2[m���[G8ݶ $H֤�m��m&ͷa#� �H���4ۘ Hڶ"�*=�� ݶ6�  6Ͱ	����[pH     $       ������z�k3+�[�moQ [xl�pUv[�͖� �Z[[l������2���Z��/êX�  �k%�CI��khl �|   h  6�-�  �`     $  l� l m��� m&   �� [@ �cm���xp؉v���u��)<֣n�S��鳍��6��m[�k-� Iz�"�m -����H-� v�$ ��� �		   m�  ��8  -��H�k m��gp��[4RM�2�mN�@[&�0�4P 5V ������	5�$ �`[\q��� $-�l���ynm�8����(�R�m�c����i�ޮgB@w�,�m��`�  �۰  $�������pp �V�Ԫ6FZ�������X *�N'v^B6��l��66���*6
���е<�R���Jy��sh1r�pϳ�l�qs�J�<�YI�r�˙����ݮ[%�ۢm�� p[@�I�m��a��&�ۀ6ؐ�[B�  �ںȓ}��om� pm�8 ��$ ��� l�a�  ���]�@A��^l  �8 m� ��m��!�-��iю��"h[������B���Sd��M�q.���`H����[E�@ $L�\	.�v������n�Iͥ\m� ��mZKn 7n�� m���IU��	�/=�f�����wn�9�� Z��nu�[��!�m� ��[C��!�  ���u����u� [oZ������ Xe��6�Hs���e�Ў�X�m�n  �U�Cm�7]�8I9t9&�mmZ��T�@ꪲB��/�@�.���HM*�[AÉ 6�m���Yf2@��t�� ;j�W����W@TG]
� ���mW �ll/m��   ii l�iY%m�&�i�|�_uUK�=,U�w�Q�   v�  ��}I�F��kK��-�h�-`   �	    ��  �m�`   8 �UUJd��;-]Y�{C3kn 
[��vN�� H$�,�9�6�gC[@mF�m�Z��ԟg�>��*�ȡ�%�$^��    m�m��    ��N��u��L�%��`*�g� X��-V��-M�T�V0��we��vŘ���UW�m$/T�I�r��6�k��5۔�O0�5�9�D�*H[0Rʲ��խ�k���tkB! /6��2���ҭ*��RCO+���8�m�i��j�$m��&�Kh����t�T���jiklv6,�K�*l��-��j�wՇu����CK�g͌��m1�VV�K���	��W�
����U��J��A�
�:�f���U��m! :1iN*UU��UAVůK�KS-�l  @ �L m� � -�m�I�l�V��m�[@� 	�ݮ H۶�I�n��l�x ݳ[F��Fl�lڵ�bt�  ���a�ր�ZY[6۷#�m��!�̒  ��� � @m�6�� i6 ղ޲+cI����/N�nč� O�����-�-�m���8��8p�%lvն  ��?�9�|���X�2���KD��EUʙ��Y� +k���6ؘ̋��n��f�,4����߾m� lMmv�m�4Zڍ	0^��iT�
�U� ڪ�l �a[Q El  �J   �V��fٶH  �aoP �zvٲ@��n�YR 	 8ͮmT��pĳj50WF� �:� �nH� �` p�kh5�f�Fej�r��O-�+ʬ��l  6�b��*@UpqQ��;5UuZ��ΐ6��U%��T��vH8       �Ͷ 8�d=OUVʵP��媫���l��VAb)��j��m���@m���� pI�lq�-�n���aJ    �l6�m�Č	�IKoG˾������ww�������!�YH1D>����� ��_�(p���*��h�D'ȡ��� 	�櫤@��C�@G�����|#�( f�C�D0QS�(� :(@���4^q=�� �_�)g���P�@��=��C������� ~@'F���	���	$ dDB�@C�T8~U}H�$
�E_�0 � dG�CJ�<}"�A�V0L��T�
<�v :�h����8�8�h*�^���
'� ��|L@;� tU�d^���ǵ_ɠ��F�Ԑ
�U=E�
�'UT��+��0�/��#�)�"������I�T�������A E���p+V�@N� ��P�U(uTP��(�|A��eTW��A�	R(TQ�>ύ�n��6]�팻s-0�A4S���:b�R�"8f»Wm���ьm�ME����:�fj�����6���Ď��[s`	-�Zl��6Ͳǝ���$���+;�����eB�JJh�6�m@Tx�\f�Cg�S<�m���3�Kmklf�.�md֣���A�,/�[]'nGÍQU:��n�)�x��۞u�!��'i����ClV��*�n�'mv�J�pSGk���������nj�3�2@�R��c�݆�z�U��d�):�e: �g�,��=Z�;vs�i�vݸbL�@tlh����5����t���鶼rn56�՚g&'H&�U���w��(p�
�Ш�y!��U��s'��vT��Tq�Įg��<=\U۷#�v��v8U�"<��吃km� �l@z첨�;[t�e$���i�WL�!r���ܒc:����EPe���ڀ�[�[t�J�ln�F��(�lV��w�ʩ-ӯvp�U]].`�]���U���m�b��*һ\�U*��.��R�<��Tnom!9�q�F�Wk��wh8�j�j�Pㆁ.�B�\v�+X�0� �]�9ڗ`���Z�NE��ӱ�۵
>�h�ȉp˫����OL���"�ZT9ܑ]D�kn��7O&���LV,G;�86�yGU�u�H`GY�!�T�[�JF{(/k�둮�"�[k��ޛ�@nY��꛴���[i:�{l� 2�κ���Bڑ���I��C``L1Ҭ��`oi��,��+5&���l�{Q����/�=�d��=��8حj�͸y�R1c:�m7��2%T�v%^�9'��V��E{N����#���ٔ��W��kf�cm ��[#7hր�1V�6G[.k^K+��Ҵ*M�3�ґ��vn7(	��s9}�v掗YV�Ӧ`���m�=m��	�wY�gxwm�3.�s0�須*�T�\x0��R�Q�[�~�_wwn�����9gl���<���6;.�*��/f�jT�:cVV�*2-�\)s��(W�f������7I��T��Q�,I���̣�%݆�!mn9حN��\9�J���-DI+��Χk�rh�[clo>�i�n�1�;9
r�y\�6�}�%��^T崮Z�j:�ct�&�	��1�q8\�WQp���k�i _C� �O2e�e�r�g�l�y�d�81�<&v��P��ö˻�@;;a{����@���i�I�����$�I����}"X�'���8�D�,Kܗ��m�m����ۚD�Kı;�����* {]��,K>���Ȗ%�b}߾��Kı;���!2!2�fK	�슄�Ԏ�n"X�%�g{���Kı;�{�Ȗ%�bw��9ı,N��q<�bX�'�{r�M0�L�ܛ����bX�'}�|�yı,N���'"X�%�����'�,Kĳ���r%�bX��Oy�sK�Kl��ww��Kı;��9ı,N��q<�bX�%��wS�,K���O"�oq���~~?8`X�sM���d[����n:�I�����ųڠs��f���L+I�\����4�Ȗ%�bw=�s��Kı,�{���bX�'}�|�yı,N���'"X�%�ｲ�;0���30�ə��O"X�%�g{���((P菌�%�_C��'�'������%�bX����'"X�%�����'�,K�����v�i�L͹swu9ı,N���q<�bX�'{{§"X�%�����'�,Kĳ���r%�bX�d��;s32]!w�vq<�bX�'{{§!�r&D�?w�}8�D�,KϾ�u9ı,O����'�,K����2[ov��rnnf�9ı,O=�;8�D�,K����Ȗ%�b~��vq<�bX�'{{§"X�%����ge\��6�fvq�,U�8�i##�$&�KN�z��9��c.��]�8\��q̅'�,Kĳ���r%�bX�����O"X�%����Ȗ%�by�����Kı=�ې��t�%���7wu9ı,O����'�,K��oxT�Kı<����yı,K;��²!2!n\���.Zm�TUM�D�,K���S�,K����oȖ1S��D�b	 �`(z5p؛��Ȗ%�b~��vq<�b]�7���~o�V��MQMǻ��7��by�����Kı,�{���bX�'�}�gȖ%�bw��*r%�bX��^gf]��v��.n�'�,Kĳ���r%�bX�����O"X�%����Ȗ%�by�����Kı>��幜2f��l.�i�z�=v��N5mi�v깅�F��7��a��]�Xffݹ���D�,K���N'�,K��oxT�Kı<����yı,K;��"X�%��Oos�33%�p�wgȖ%�bw��*rr&D�?w~��<�bX�%�}��r%�bX�����O"X�%��%�d���)�ss4�Ȗ%�by�����Kı,�{���c�ș����Kı;��9ı,K�{ܗ,�݅�3r����%�bX�w��ND�,K����Kı;��9İ>~D?<*+��|����w�����x�D�,K�=���L2Y���wwS�,K�����yı,N���ND�,K�w��O"X�%�g{���Kĳ����~�,Y�`�V��G]A%�N�9]x�
�궨�֓g�t�S:��w{ͷ�=�܉�f�����~�bX�'{{§"X�%����'�,Kĳ���|�,�&D�,O{�}8�D�,K�ܹ�.m�fe��wsJ��bX�'��{x�D�,K����Ȗ%�b~��vq<�bX�'{{§"X�%���e�w.f��ۘn乻x�D�,K����Ȗ%�b~��vq<�bX�'{{§"X�%����'�,K�����:nY�ss.n�"X�}��Cb{���q<�bX�'�^�Ȗ%�by�����Kı,�{���bX�'�cݧ-̷@:�#�.�!2!n��Ȗ%�a����^'�%�bY��n�"X�%���y���%�bX�v~��ő���plp�5� �&b V�F�.��bAVRF�v0B��!��+����q�:yEe�ۃ	l�MXN�c�d�f���m�@q+l��Pfx���kp-��F�/a��C��$��v� &C�ܳmmr^�p�xm�m�G%vۊ���N�q��γ�n�ݮz�eE�k<g�����ڷm��Y���M��8:�*F�\��]���Wm�X?=�tæ������uv6�&������Q�@n9���B��x�fؗ 6�:e��~��ı;�����%�bX�w��ND�,K����	�&D�,N���'"X�%�zO{��;���72��'�,Kĳ���r�r&D�=�y��yı,O��8D�Kı<�{���%�bX����^�4�%���7wu9ı,O����'�,K��{�"r%�bX�{���yı,K���'"X�%�{�ӷt�����ssgȖ%�bw��9ı,O=���<�bX�%��w�,KP�������%�bX���.m˛fr�ݛsH��bX�'��{x�D�,K����Ȗ%�b~��;8�D�,K��p�Ȗ%�b|��'�g��zk��ۛBL������^�m����l6�.�`L�j�0�JY�aV�����,K�~�q9ı,O����'�,K��{�"r%�bX�{���yı,{m��0�w2�ff��r%�bX�����O!�WAO~k�����#�S�؝�bn�p�Ȗ%�b{����yı,K���'"`"S"X�d���̷2ݒ��˻8�D�,K���S�,K�����Kı/o{���bX�'�}�gȖ%�b~�{�,��䬗f��iS�,K>RD�߼�q<�bX�%����r%�bX�����O"X�%����Ȗ%�b^���2N�6��]���%�bX����ND�,K�
����q=�bX�'�^�Ȗ%�by�y���%�bX�=�se��tٹl�u��B�s�cO�c]Y�BpӮ�Pv��vv.���;�V�8�DT����{��2~��vq<�bX�'{{§"X�%���gȖ%�b^��q9ı,K�d�����B����͜O"X�%�����|�$r&D�?w�}8�D�&Bd'Ϻ�����ei`n�Nu�qiG�f��u���������Xz|
ނ�C���7��'���4y
:6�R4ۍ��� �l�<����� 9˻ٟ�L����{����s� #�R����y���ۄQ8�d#����7[�,f��nj�`�(mז)3�:��];[�������Ҋ��.���N��T��8� G&�=�Jh#�bf5�$���<�����ouXͮ,��W�$�F�Ğ<�o#M�@>�}4=�M��������=\bT��d�(���D'��zX����͵a	CQ � N�T��{��w�=�n�3"m:�&��svՁ�D{7�/���`y�Jh�9؛�rc��92/��c]�1��vn�H���.�K�q��2p�
¶0��sj�wi�qR �M@{��z���B��8��i��h�ھP��B��=�\X��������T�T��􌑍�4=�M�������������m�J��@G"���rj��_���C@�[+1�P�73@�S@77j���ZX���J��B�V����z��]ѹ�=F��\�vd逈Mq����p�M:d^���B��mّ�+�u;�&�جm�T'9�6��9��e幸�N��[\ji#j�\v�ƫ�._�]@o[fT��-�kl:3��B<67mU<��Q��qt�,�v%�̱H�klw\n� '��5�5�����L�vƽ78띏G0��ml�����Gqm����#��w������>�5j�(EӻyF��ۭ��q=�)����/\�M����PxF�7�fB"nL��w��<�@G"��� �[(��fPY��m����ȩ����~�Ă���16bY���w,ٛjϔB����V�k�VeL�m�m4G1I&h{�s@/[4=�M������8�ڍ��� �ݫ�J=�|~��Ձ��ZX����~H�u���=��l�[OX�|�\T�]z\�Y-�z�w�(n�.�W7u�{r*@{�� G&���i�2�HM�#�,��WK�(�yu~HZ���@{����,.n5�Y#�9�����^�h{Қ�w4�Ղo
̆G�������ȩ�{��e��e*��:��?{+K�$�.������z٠}�w?�$Rdyqtu�;H��;`j������6�f(1O����XP5�9���BG �����)�������s�7Sn���n� =�`�#�P�@G"����2dmF�nz٠y�JrxS�����HYe%eQ�b�~ ����:D�%��Gћ�'��BR��O�&�k��`$;jHi��a	HFD#���d ��d�q$"�B�]2b�F�d|-	B�D@�0 `@$����CR"��)�D��Qڨ��A�C�EJ���t"�<Pz >b�u/� "�b��Z�sm~�ók�7�t�T�T:eL��U�C�m�`v�Z�?{+K ��4G+bi�)�&���4���no�	6?f���(����=�\t(�������~��:��dQ��۱��k�c���[t�f.ɞ5�\�����_�c*�]�S���^�J!&����?BQ	>����k��-(P�w�Z���D$���nd>�P�UK���;{���K�P�)�7�����7�}��ٵ�(Q�k���3(STS�����o��P�v�~_��mqg(I6v�U�v5=4�dc)�tC��?��j���,sv�Jz"{`���x�/��P�O;�@�=���n�Mɚ����q�@{�� ��h��c�̽�\صp���##i܋�!�f�v6�����;	�����с���Ң������@{�����@s�w�/i�diFےh{Қ�w4=�M �l�9���ئnN�U =�`�#�P�@z�3�m5�L�4�h{Қz٠y�Jh����V'���7�����s� #�R��	_��~��R+{v�����,��wG`���58Z�ưSf��MU��+��lp�i�u�B�qڷH�
gX�D�[����L�(��_c}�L����j�c&�i�����L��7J�v��ⱛe�::�NVY�'z�ݸ�Wm=7pL�&@���e�j�֎m�`���|.��H�����Z�f�V�ɐ��ط+u��^�'�k,�}P\�;臲]��O�v�p�֋���O:m��1����;e�7���"�z{gƁz���zS@/[4�c�clB	!#��\���@��s� %s��y�cCn5$�L�<��4��@�ޔ�/[��[ȍ�P���#m7 �M@{�����@s���LdiFےh{Қ�w4=�M �l�:�X�jB8&�F�I�n;�p���X����������}������(��D��<��ۚ����^�}�{6��<��æ�JM�L�+�������v�U��6��77mX�֓���1��&���������	$�}�֬f�5�L��"9������z���zS@/[4�`���E!��zEHs� ����O��g���74�.ݭ��pS��Gm�ɰV�ĥ0��l=<l��,-redjk�ͷ9�95�{r*@H���%q
26�p����zS@�n��)�{�J:EsN&�rM$�����'}�xr~8�H"�'�O�UT�T��{���O����'��lM6�1,n$��^�s@�ޔ����zS@�[H�E&	�R6�X������>����k�sv�@����o�F7 ��!��$^��L�kI.�c���t.<u�Sd��m/OiA�P~��ݼ�<���@{�����)�r�WN��	b�94=�M9 =�`�#�P��E�+�ͽ�s4@G"���rj��4��:ۓq7$�f��)�ɨs� ��r�T��ٹ�����J4ۆ�^�h{Қ�w4=�M�Qq�dG��C��p�>�tX���m�3a^�.��ʱ�'�
�!f(�M������z���zS@/[4�v��lS��Ln�v��@ɨs� =c��a7H���#nf��)�������z�� �Z�t��~$i�@/[�@G"�U��.��/>-A%�HD��<��/[��y�)���`lB�ũl�34*m�Rd�'�z۵�R2�W]�3�c+6YA��X-���B몧����N���kgX�՞j۴���2�N&:�!]��1����S6�hvz�連l��-X���� ���������;<��.�cl���ѷ�������݋+��һ��Q��<r/۞�gs�ɘLv1]=k��#��Z����n"�'D+�
Y �n�*6���GV��G\�8�48+ݸa�5D�"�T�\����4�b�dn������M ��~��ύ�?�qLI��dRf��t��^�4;�4����U����Q�7 ��<��:EH7�@7.�rz��d�������Ɓ�}���t��^�4s��4�Dı����:EH7�@ɨ7�@ut��T]��]g�㥜�He�!'[��LS�c��u�	��m�CU�^)[���{���{� 	D�s4�ͱ�7w.l�w�{������W��~�UM����*@{�� ��f�,RB)&��)�_m����{�|h��4�cl��	E!��:EHs� ��W��_�����������SM�I1�3@�S@/9�7�@N�R:1�+��.�J�ݸl)\��h��+4��rc�+un�l��H�q!H���$����~���@�۹�y�Jh���D����L�f����/�!���Ձ����/u����&�h&,j&ۆ�}�q������U���im�@w=��մ�$�bI�F����M ��hwJh�w4�kU�� ~���75��	�*@y��w��Z
��l6^���:m�z�cr��d��ו
M�:��N�^�lWi61V�u��	�*@y�� ��@��6ʌx")�4��Қ{��<��/�����	5�dR���2���ڳ�o۵Ł��j��i�
EM�$p��f��t���ݵa�J$B������������q��F����4;�4�g���g�{�|h�@��Zkj4�kE$�{��x��vw�s�����&�ۖ)3v;+Y5�mo��݉��"5m��?�����)�����D/��oWŁ��[>���M̪��4�������S!�w�`f�|X��WЛGt����5UUNh���?{+K>�P��3����7���Ƽ����6�U�Ô?f�gu��������U�v52��J,��73D� >�ǀ>��@{���I0�?+�(�F���f���
PҜ@��w�è���b0����H$BƤ,��$H�,�! d	8�MF1q��{�N��\ �b\	<�Q�S��e���� 2�B$Q��`M���X�X�IA���H H'�"9�B@PbHȲ$�8�8b8���FE����DT��`FBI$$$V`HDBH�dH�I0$!@�!$$#!d$$�	��0�I		YI!#� j��*ES�C�(����B����"Ĉ�+�V��0�F�.0 ¹���Ak0ـb@��V,H��"��F%aXUuW'<�ݓwI%,��gSl��q���I\U���n��g�8ݝ���Kv'�nQM��u�����ݮ k��tOn��붴cmoT_ [@d8&�^ek<��#�{E>�2�8�n�q ���kH�5b��۩m��
�ۖ��ANo;���۱U`��f;	���,k����.^^TY���v��j�h���Ckb��K�;V�ͽ��%^�Z�nJA-vh��j�Z�/pC�+ԯ����(�
H4�U�L�j���YN�Ȇ8ɩ�a��K-�#�T*e6+��'�9��c��V�]=��*�
��BJ9�"j3K��@�x#�:q\�(4��\��,�ض��;$�q$�v:�
��L�v�������Yf��$9`�]l*��eSm�#W�2U<��U UOC�8�E+��p�.�\mKGF��6�ڷf�d�� �`H ��[WD;�#3�.m��uqWTp
� N�j����u�k��ѺU����v�/uɱf��&1nN�mհ]����.�gi�T�-�rn��^6n.�J�n�WZ���µUUl�-U*��<3J_/�r�*�q۪%�q�ح�6֥�Wm�⮩Iy��ę��
i�����y9ʫ�;AK��j
�.w:&�k�Yy���8����V�`��ܦ�L�u92(��}��*ɮ��tp�� �5�r��lEv���vr�@9c�6�`�
��1g㯾�0��m�!۝��\l���4��E�g��n
��r�A�v�@r�K�=��**�
���x`(6�1�32�ݰ���^v��[��U��N;qnihL)hx2�g�g,=����w�|�۠(-��\eͳv 6yL�UDa�n;�N�U:1�V�ӞN��L�<����D+v�V�6
���H��cj�э�O �W[PA��CQ�jS%�\*�9[n����t�ζ��K�9�T3����Pu�:1��vU�.� 29,���j�UB"�x��8���q������j
q�_]E�DN|���W��a%˝�%�m�cBk]4�	$�G��.�d��:NX�j\�-ͭ�ȋIZ� Y�X��*bo��}|����r퍶�2�.PQ���z�×�)��W����
�km�6I��2�I�oG
����T��.��b�möG�]�&k�<v�[�e��Z�:��}���ę�{vu���V��NKm����(cݮ���{���o��mU��s]|l�⻶M�6��%�'�G�e�;�tN-�6����s�2�,\q)$Rg�_��h�@�ޔ�3�w�nh�#$)I&�p�L�ݵ�$�(�"d����>߾�`~�V��4u�4������@����/����oٵŀv�U��D�Ӗܲ�d�s34Xt'���X��V��V��w�@�_�X��D�m㑷3@�޻H�������� 'H��Ż�i�l��ӻyF��m֗]�ڙХɢf��iwG�&D��WM��\�I���~I'�'ڀ�=�t���Xs�*@K�2���nYisv���I<���r���|F+#(AH0H�H$ H+���$��	��!B]���Ձ��j�73j�Q	&ð9��<
P�uEL�`vwZ�?{6Հ^�4=�M���LI5$n�X��j�73j���,9D$�;�-��o�"�$܎I�{��=�`��"���H_��������n���F�՛<���v砚�xzۯ0�:{[!�H�@���51D�mɠy�Jh��V�f��K��z��Ou9d�"Hj&ۆ�}�s@�S@/u��қ�g�H�_�X��F��Hۙ�z�� ��:�U��~�Ũ@N�R �Z:HH�9$R{��<��4���� ��x	Ѝ	br){���c4�� =T�#sPW���5X���Z��n6q<�
���m��	i��I#;]����Ӳr�m�Ek3D� =�`�#sP�@J��u6BbȤmI�����^�4=�M�n���U�8	&ܓ&f�75�{� =�`��AGG$4�m�4>�ߗ�w�@���X����J4�	rB����X�Q:��a�D�p�/��h{Қ{��<��4z�rH�dpM�E���1����&��R��"��:�{s�r������#0i�F�� �߷4�Y�y�)�_m����*�'1~X�U9�`��6{6��;;�X�6Հq�<�F���RM��M�b����nj ��2�e]ѻ��h��"����nj��=��M����)Rf��u��ٵ`~̭,��B"	�""!,@� �! H y�K?S}c��[:d%��Ix�^P̔ݕ,�$�^�p�-���m�u��B��������u��y�n\�pT�"�m:��&8��������8���d��cq�ps��Z�I؄ ��s�LZ���:*�7k�7�6u��k�tv�j���89Gy��\��d#�v\�նQ�\͍�6���&�=n8`����w,��g"��+4g������yYS�h�]sC͋�+���=D��g��ô3ɲ���z�A�[�"g�5#q	&��s= ���<7۶�����3��V���~&��ANGS33U`~̭/�Q���j���Z��f�~H��%�67�����vwZ�?fm�9��z�n���2Ʃ1�i1Hۙ��/m�����hfV��gw�`��_:N�p��QY��#sPt���|��R������i�sϪ����v���/�;h�WG&�� �0��Z5���O~�M��ٻ��߄� =�*��`}'ڀ;�l��4�7T9�,���L���V�ޫ�������:���LԶUM�+7��`��gC~ͮ,��4�,j���,I���� ��V�ei`o�mX}����V���~%Ĥ�M�ܚ������}�����s@/u��UcB��	&�S$��Ì]���L.ً���ۑ�O=f۝�1���w�d>��67������w�nh{�s@/u������:��T�4��m��=�*_�vI��9��@N�R �Hbx�9���$q���f��t�����_m��=��h��O.6���su��	�*@y�������@pU�F�bQGn�����M ��hwJhnW�N$��"mn���е�u�ǵ����T���1#����8�OQ�d��3@�S@/u��Қ������	#K����� F�<��:EH7�_~�G_�G��D�#m7&���@�۹�y�)�����Ԟ7��%ә��âQ�;�+۵ŀnfՆ(Q*K�V~���nL�vU)�K�7s3i�Z ��@y��t��������_�������r�3e
�n7\���Mr��c��7��)�5�t�v����Y$��x��M��M�n��>�@8��tBXێ9&��t��}�j�����}�W��֛:�����3E�ٽj���ZY�I��z�m���:�&)��E"�f��{9�@y��s���n\�㐘(ԓp��Y�y�)�_z��'�����p8�"�����I�n�;f֎�q�`�r��i��ܭJ�+z\�A��v�i%5��s��)��n�mj1� �)����h�W��4�-������3HmQϯX�؍�6���������;�;U�����ķ9Cx�3����x=:��b�&�B
�>�:�=.����g�϶2�Fd6�� �s6i�S�b۶���C��<��d͛���ݳ2I�&ϋ)R͂fui�v7j��g5����&���MF�ܚ����/�w4;�?�~`voU���t盖K)
]9��,�m��l��Z���?fV��մ�s�$�#Nf��u���Y�%߷k��zՀj7Behjj���a��f�Xݮ,�(J�(������ � ؈� ��~����lllog����L�%������|�������N>A����{�� �`�`�`����Â�A�A�A�A�{߷��A�A�A����(���}M�4U�eP*��#�#�D�8-�n�i�yd�܊]W����b��Iƶ�ݛ����lll���� �`�`�`����Â�A�A�A�A�{߷��A�A�A�A������ � � � ����}��I6n�ٹ� �`�`�`����Â�U�<A�A�A��>�>A������N>A����{��"�`�`�`��O���.���]˻����� � � � ߽���� � � � ��y����lPll~��xpA�666?��}8 ���K��avnɗ.�L�����lllw��pA�666?{߼8 ���>�|��������|������[ϳd�e�C.��͜|�������>A����{ϧ �`�`�`�~��o �`�`�`����ӂ�A�A�A�A�}߼��ٹ�&��0"�x�8�c�;[7Z��+x[`���(��%�����̼ɗ94�-�.�\ӂ�A�A�A�A������ � � � ߽���� � � � ��y����S�r66?���Â�A�A�A�A�����0�?��wff�>A�����~�>A����{ϧ �`�`�`���}��� � � � ��y����?�����}�73���-33sswx �~��ӂ�A�A�A�A�߾����lA��ф�� �$'B�:b ?�D<��h:�IL �<?�Ā����vy� 8	,A��dHň@�BB! �B1F)0�1H0�9�T�G6@�LQ��h��U��FE�03����BF�`��b�� E�"�u��
 ����x��&�����MDSD@8�7�*��_ �`������� � � � �~�����lllo���}�.��sv���>A��F��~�Â�A�A�A�A���ׂ�A�A�A�A��߷��A�A�A�A������ � � � �����2̗I6n��wN>A����{ϧ �`�`�b#~�~�>A����{ϧ �`�`�`���}��� � � � �݅�3ww.a�wM�B��p؂�$ל�]����	Vu���V�Ne�]v;wf���n�ss��A�A�A�A��߷��A�A�A�A������ � � � �߾�������������� � � � ������0�4�.[�s3w��A�A�A���>�I>��4uz{��/Q)d���a�D�p�/��h.���ď��h�>4Qʱ�b#ē������ ��@y����t���$���Uu��^� ���� 'H��}^�}��5!&L&7� ~nc��$�鬱�[�E�!yУ��������q>2�3777u��	�*@zۘ�#st��V�i		Ȝp�/��h[snj�����/J���soLݤ���75��	�*�;�j��d��'$�q�}�/��h&� 'H��nb�܆U鵸�Q��&��t��}�s@�wW��{��TqV#C���e{sv�˙v9�u;(pf�@�W]�7-UJ�K+]�9�5��h]����:y3-U�I����2�ۮ;'gB	�c����I(T�.psnA���݋^#ATm*���)s���H	���g;=I�c����ގЎJ��Q�c�����ܩЕÝmq+��1q������$�Хrm�'h:p�u���	Q�m�A�z�y��b���;�޾}�mP�.������}������f��'���i�n������8��Q���y�bƢm�|�nh.���Y�y�)�z�U�;1G�&)s4uz���{� 	D��U�@����/wnj���T����@8���&�!�rM��Mt���� ��8L��.˲�v�sD� =m�@��7��;׊�7$�1ŎL�����"]�-F�؍��z�fNY�:|��8�l3�qv����7i�nb ��@y��t����Ad��'$�q��f��T���Dyg��~��~�߸rI��@�QѨL��Q��&��t�t���� ��p�ٚe��)����د]���� �y�7�g����I��ND����Z ��@y��t��s�{w/6��VNV����7\�<ݳ��Ґ�fβN�Or�:�� a��`�Df,rD�~ }o�@�{� =m�@o?^M��0�����@y��s���� 	�n�_@�$Ą��n8h޻��3fɘ�J�!B�����V{kK|Jҋ��8�$���^�_z���M��s@�q��		���377�5��	�*@zۘ���_~�_��1��UY���zv�ѹ5���Smŗ]�s�����RA��Ů�R0�����	�*@zۘ�'9��JW�x�,j&ۆ�}빠x����Y�y�)�z�U�;1G�m�ܼ�@zۘ�'9�7�@NqR �n�F�l�9*�����
M�oU��o�s��*���Q�"�3��6�q����Қ�����@/�f�k�� ��#��"���B\+�4V���S�.iv�Ngc���Z�k		&���BMI"������@/�g߼A��@����X���	&h�� 	�j���T�}Yr�
�b�= ����Қ�����@�jth�d�ډ���7�@N�R�������>���/�ĒOōD�p�/��h.��s6�ٕ��q	&��f1�n�K���ӧ;�#�y�vf�t`뮺�K�O)�6��m��<�Z�5�;,%�6�g��wXN�3p�s8-�r��n��C���}���*��kVԨ[s�H�wX��N�s��,�:0AI�h�Cl@���E�Bi����$�I�.�w��{[ �N�3�gy:��&�ӊ�ۘgn����)v�y1��J�`v�ٛ^2+�+�ɒ�����y�N���V�p&crkf�WE�HE�N�M�����y�����D�ˈ�rA��_���@/u��Қ��� �Z&���A8��Y�/�"d����>߾�`~y�7�a���?�M�Ĝj)&���@����<]���f�\�+��!!�,:}�ߕ���`��aС'���@��,��	�L�<]���f��t��o]���`�QD�sC͋�;M�T&8��<;i�M��z�
�lģ�?~�ٛ�h��sq�1��w�U���ZX���DG�y�6�1��m�L�w2fn�$�~�{9��@:�:͵`~~͛ �n��I����lBC�1cQ4�4��s@�{�����}��=�>4ʱ�f(�nD�V(I?NoM�v�U���ZXt$�{�f�}��M'��f<rD�zz٠~��]����nh/z�޻nA8�ɺ��M��C�;p�d쎬�5�n�jǪlv�e�#��ɦ��l�m������r*@z��@ɨ	]Yl���]�H�p�/[��$z������@�ޔ߿$}B��PpI��E&h��6��VJP�B�*�z�gu��V5Eq4��9�8�?�����=�>,��VD(���9�6�1��J�JcMF��������[�����= ��4X[�B8$��HL_�L�J[���9^!
z9+�j�ɷ�y��D?�����t��N\���X��f�7۵`y�Jh#�i��Q�$܉I���k��&C���3z�,��V��$x�Qf,nB8��l�<����K�~��=V���y�U�M�ĤdNKQ۷Ł۽j���6li(z�؈��L�mX���%L�ni�P�s6Ձ�������V�+K?�����gT)�6��$��\�۶�r�e����k9�Zy��4��vJ6²U��H[��5��>����>��H��E�"jbj8�ӏ@/�����I�7k��zՁ�����!&��c��pS&D�lnI�u��@��sO���!�=� ��w��1���Ժr�h��>���������X|�'��������BNH)3@�u�@7۵`{2��73mX��	��(�2)D�CC�R	B�$���zG�R� ���v$d��ZaX7O� ��H1H��X$B$&�m�`'䊑�����	B!, D#�EbH�m눧��X,h%`$��61�"R,�1 �w�H�� �R�VFaHB#	*R%$("D�� ��b �S)�dI D���JSKD�H��R`�������vM��2fe-���Y��ڱ�P�Y�^74m��3#�r2W�e�6�WdTМH�f���:�3v�<���	��퀶m��7 m 	�[*c=����ۮ5=<��2�`մY��,�m�m��3m@U���^V��CFN���TY%9��v�f�g<���0�+���-��VFJ�6���Ҋ�p��C>剈�TČZ�������aJ���\򶩝�<2���Ci���j34���*@���l�� rjn2)�d�����b:h3��ɉ�eY���;�#�1�U�=	օb1�t��p�9��U�ؠ�[��!%��M'9ٳ�=CZ�^k��
^��*�L�w@YD��V��kj�v�q���t�G��GNd�$6�4VN���ζܳ�%@�<r��\�&m٭�ԶKh ��[@�lֻk1/`Ir�ۜù.�\��
ԅͥc���s��.��U6��-�r��Ϧչ���S�/�ձ��vN�i&��;M:6� �.��[	�[a˴�8
�u�����M����kw\Ԥ��*����9Pr6漡qbZ���UmJK͕�%�n�]35ڕ���8+ѧ��ͬ��j���zUr���h]�c�1�;�x��OM/gY�d��p4��q3���vj�v9���y.L�X���Cp����*��V��2�n�@��g�Vݨ����X���m�n����k+�W�R�IŴ9ʧ`���%L���A�UR��Q��c;c+*>19e�K���R�_�n�`�ѩx�b��m����g����v�����y��T+��������n�� �h*��۬KêuحR�Ĝ����58�g[��"��kE��+�[X��)2�`Ĩh��J:�S�G(F)r� �7K�Z�l��\�Ȭ���6�.�e�5s��%�f��X -�u�`Cu�0�.7P4@Rm���z���@���
�=8�����*T�<UO��gp��ޓ����e��驪��(�z�ΦS1�%�X:�u��T����&�;�֊�%'Q�vc���B�n����um._gl��΂֚VH��e�ncnx�nO�*V�Sq�b��'kI�tۊq�<�n��F�Le2v��-G[D�`lO&��-��8��������8�x����l���rIa",�Jn^�K�������:s԰ܻ�\䭣�n7\��yvn����W:�5���g<ި��"r> ��h�Jh�����=�R��|�&�bD��@���9 <�K@ɫ�����V_�ё�$�$Q���ۚ��Zz٠{�)�{p��Si�ܑɚ�������fV�������}�s�9�qh�f��t����j����������I��*6h�=�->�9�ˊ�K6
�#��m-�d�:���W%�ޡk�pS&D�lnI���^�s@�@/[4xJ��,l&#.ܹ�9$��z���?.�����6�{~��fV��$���Ιr����rB9�����m�~K��X�֬Q�I2N�4���\Ӱ	$�7�@H��Ihu�?\�&�bD��@��S@����;V�[�hZD�N$��f�-��h���cpp��P�n8�5�dz-L(Ć�$r�w4+�h�g����|h|��	4�RI��mi|���ޫ3��w6Ձ�#(Ѩۙ�nA��޳@��)����A"��B�)�U�9�~��'�?��;څdȢ��I4>���BO3���zՁ�N��ڰ=�ک�K&%��6�[�s@��j�z��l����ˮ7���H�4�qx���<�X��}4��)��������U���\J4�#x����3@��j�z��Қ�w4�:�:E��Q���	�G�@H������]����} �@�I�I4�Ɓm��}�	(I���v��VyK�ji̒7)H8�4m��=�ڴ�f�߿~_�C��2���� #9�{���A���	���ړ4}}V�[l�<��h���.+��r�"o!%�����
�9a.{�v�,v.x'�����']'2��5s!I�'�[�h{e4z�h�����Q�qFH(�j������"M��֬��̝�`}~�u��K&%���p�-�ݎZ ��@{�� z�f^���IH����_U�����M޻�p��<yY������z��6	T���- �~�UW��~����$�L�\�)&�m$���n�إ��+�����K6bc���J76k<��5���0�MUlt���F{GV(݂j0(��u�Z�D�Q)������Z�D�"ǩmڻf`���*@tq�<nX���o@�����7hj�ٽ�v��0cOi�/=tSF��9^yx���ƮNv���u�ut��3Ό��%��L���k[1��s��!��$�]{�mm梧Z��cIP	C�f��<4lvAdo��M�@�Ȥ������o]��_U���g��8�`�sw/t@H�s� 	��l��E$M<��䙠{��޳K��^�޻���8Oؓ˼� o��=�`���H�r��tS��69$�<��h���=��ZoY�~����#N&��n���}�BM�Q/'G^l,9�M���7U��Y�&1��'X�0��Q93�>����{��޳@��)�x�kuƤ#i%#���嬫���@wM�G/���4|�Ģ�'�}��h{e4z�h����{��"i&E*�?�����zՁ�Nk��ڰ1{���ҒC@����t�/ >��4=����W#�NL�qc�G�:���n��]�4B�ٵ�]�quE��^ͷ`x�pRA��$���h��� ���<��}� ����݃�>s!M�36��j�6	T���-UDDG�'o�u?ӥ4��Ӓj��߫��'{�xrz/D@������=�h����RU=Icd�qD�49'ݽ�X���}�V'����2���5$M�)$��{������ﾞ�}��{���tu�H(I�Z�v۔[�n�\=)Mӂg�K�<������]��(�<y�������@��mX���(K���v��0��9l*��kw7P� '8�ݎZ ��������/��7fY0�]ܛ�p���v9hs���H�c�) 6�$q�&h}��~��/�@>���?{vՆ�Т"'��o~V��P�sJJ�s5D�; �fՁ������ۚ���@���S$n(�#P�$���b�������y��hv�n���z� :�ZLM��2H�crM�m��/�w4}}��B���ٽVo6�Ͷ��Hd�9���T���- NsP�_�_����{���o����*�L��m�?���6��Q	7�����޵`��*t��uS53N��M��U����:EH�r�Q�*�yv���U���ZX$��K���/�=��ڰ>�IG3\��.t�[d�P���]��	n�j�7V�[�8�k�6��-��c\;[�)0Vc*vFvD��5�Ԧ�\"�u���5�� �$λg��B(M r�i��3Â
î�N�_nݥ�2l8s����>1�vnW���g;�o=�
�ܷ:}^Lqل݁U��6q�7�5�v��trJ�m����uNZX�P-�˹�A��ky^e+7﻾z�o�u�x&����N���@ks�������#u�[l�ƲLy1�G20,jFI@��U�{ٵ`���I/�=�\X�;<)2cm�q�$����o����}o�@�uq`o�m_Д6f)|��4��*go/7P�}�t� 'H� w9�}�R�j�"��I4=���� ��jÒI7۽Vo6��1��j�6��4@N�R �sPnj��M��.9�DG���� 1&���K���^sd�Ȩv�j7Bl�Q�>�����]J�rF�jH�Ng���4�Y�y��/��h��cC�Y�H���}��U4D�@>Ur{Ϸ����V�f��%	6��O�S��6M���uq`o�mY�%�37��>��v{�qd#�Ƥd��/��X��V��V/�Q9�~��>�'���d��c�)� �޳@/u���M�n���_|��R&�l��O��@������7\�&�V��&��\;�u�n�I�w�J����)*J��.j��w�`~�@N�R��t��me�n�3NI���?{kK�脢&O��X��; ��h�IT�%��7M�@�ݵ`{Ӛ�،H���P��4�B9���0#IP(�	X@F@פ<6�|��y��$!	 ��HD�HD� ��!!H�FA��bD�@���H� A0�`���0Y"U�!��b����C@P�U=��Vx���
#�������`*��<?���M����}������nH�mBI#�������%;��; ���?{kK}�j�5�)Nt����u3N�73j��GТ#/��Ǡ_����_U�[Uؓ�N8�M�p\�l�{[����8FsvM��h�Ni����I�H�RdM BN94=���vՁ�Nk�
?0;w��Պ^�R:hX��4����@/u���M���ؑ�����d��x��3@o'րsP�@zH��Yr�(Ԅ���cqh}����4{��y���$��H���A����oo$��!K1����LrI�y��<�ڰ=��v��V������*��6k\{p�mնtG��g�h�-��^�V��s�ݱu�����qˬB-�[o����� ;��@��t� =gL˛��F�Pq�&h����1 ��4{��ym�������bn5�@;���lM��� �o*�ֹlm74S�������������5�f%��}4��S��ؒC�28hM���$���M�Ug�+��ٿv����8�[�lpۊ��3���j�&{5뤛�]]��k��ٹmВlusZ���<��);n�c��q��6Iֽ��y5Ls֎6-J��R������ex�T��gg�I؄U6Η�L�6v;l��Z���͗8��r̠��
�k��6]���;0(�<�z����ܽ5v�����[kqųU�#�s�j8�[#'��*K��������~�������6��f��6���N�n.4�8b�X��64�dO������i�9�8�w�hfmX���п0�wZ�3�\6�j�Q�����@��)�ym��=��[�g���~B���L�om�&����I ;��@���vE��!1F�p��1}�}�h����Y�y��<G�����k#��)ݎZ꿜�|?��9�Hq���\3�=K���j�%v���:�����˳p�I�+��u�V�N3�Gp�Nm����l�U�U��}h���}0S!9NM�l���L���VB�	%��oe�6{��ne�g��1F��jFI�n��Nk��gf�Xή,����4�m1I�f��.�~Z�_���SC��~�4�3�%����cqh�5�\�_�>T���-�&+&BG�Ŏ�z�R���v��s��`��=��Ԥ�"Ҝ�1(F*��]Xs*�����@NqR���ް>s�@I�v|�<si��p�/�w4}}V�_z��l�������}s#i��G���Z �棪�l�T�"7dd���&��Ӛv�f�Xή,�m��D'�[�����R&NE�@��)�}��y����@/�j��Oq3<���t�9t2�$�V��+�z�h9.�ȑ!u�qt��V!��]���r�bě��C�?��ۚ���@/�f��S@�u�ȓLRE#��{���M�f�Xή,�m���1OI���Dq	Šu�h{e4��ľ������@�څ,��&D�y��t� '8�ݎZ	���W���i_�(�K�D�ޫ�ͺ��SLs3S���s��ߛ����>��l���߯�~��^�uE�j��`��}Rʚ��c�af��&坣u��u)�р��ʧR�d�; �fՁ��ZtD/�zC��4���'���f&�Q8���h{kK}�j���5��rS!�ޔ��^f����@{�ց�g;@s������j$�&�d��/�w4}y��73jÒ~ξ,�^��h$���v�siݎZ ��@{��:EV���bj������*RT���8�X���2
�:���ԉ���p�WX�;�78���m��4��FGb�l�'�C��b:��Bv����38A
�3t����:�0mV��ːQ����N����m��n_+�M<�)�;���q�f�p玐�s�	�� �n ����k���Z��f0�!u�HɁ�(�������B��PS��V��z�ts�q�"�@�s�F�q�뭇ki��:ۂ�V�GO���}�T�.����}�t� 'H�ݎZ�Y{fI�$��nI4=������Iw;��$���y�߳1���H݌X��9���3T��gw���m�N�v��B������$���Z�K�z��r��J�����o�>Q	Wu����������߶X�$���3�HXZ��Q��QD�-I$�u�x�K�,Z�J�o��%���ԒVԕ��dBE c�nB�v�K�\c��a	��M��P@��wwsv�x�`� Cn8����K��E�$����x�]��-I$�u�x�]���h���ɻ�ym����<��"��w���$���<�$��X�$��#��ؤ�G3�K��ũ$���I{e�RI_m�<�$���S#q%"l�!8���$�f{w����y�����w����.�w���څ��&L��6��m�ki�m��B�D/��f6�t�i�m�{��Ē�z��	q6�I���=��֤akr���f�Jz��s<�h��f0j���M��nE�I/���<I.�w��W��<I%�-I%�=J�4�1����y�Iw;���?f6�_[��Ē����I%}���Ē�6'C1F���\��{��<�����^[�(E�U�/�P��_�;�9���<����ũ$��{��)���NO<I/]��I%}���Ē�wqjI%{��Ē�x��!91IԒW�|�<I/���%�y?6�w}_�6ߧke�m�N7�_�una����ӌ��l�O0�g�e��%�b{�6�ƶG]6ܩ����?�%���ԒJ�Y�%벵�fx�K���3�J�_ۍ)bs�-I$�u�x�^�+Z�J�o��%���Ԓ�څH1Fܒh����w4�"�޵`��`g�l���4�fk��@N�R�nj	U���ߗ�BD�]oM����uL�4�e��Lͤ� ���9�	�*@ymo`�$$��7��1��m����|������W�kƎ�m��6�&[n7C���@��\s�U��߫�ϖha���`� Br(ܚ��z�vՁ�͵`��}	�SZ��%���MJsU6gu�=�j�7ٵ`x�W�^���m�I�f��fDC�����z��sf�脔'ٽ�X�m|cn��'0Nf�_z�Ź�`o�mX��V)�+ވI\�DJ5�H��x!	���`?��aaM@�T� �H�B0��ȉ��K��f 8!�^$1�"0Agy��7wm˅�ۛn�@��]�;� ���������մ٣����T�K+�)Z8
Z��"�-Զ���[e� �� ���,�[�+9z[ת%J��l������c�aȼ��z^��m��H��/[���ۍkj�$æ�[��VM�1s�w!lm��wn��0�tN9��x�;=</�rޡ�A �p�j�Ѕ\r�96zә�O<��Yf6*��2�ې�`l�5
��C�V�US6�f�vŶu2͜�['��f,qBVۋe\Pq;�y�Wk�4�^4
p�uAʚJi�ջt]�^�Ӥ:fD	�H��a�3ˎц�페�ڥ��a:4T�d��8�]:�j���p�{j���p[Df�0���R�U;�U����[n.�3�GYgZ�P��l��Ӭ���5�]� d]�� �n����*&�L�r;`�7jT�Ws�4�ԋۍ��z� 
U�Q͡^kH��}3m�4����s��[�V����8�-�]bH��8�ݼ��N�c�\���l��ݫ`.U��H�6�-��eV-����E��l7,����L�c^��P��G�bݠ���8\�����3�X�@*�*�MPL8ÎxM�iܦ��b��G��.�cfP젼����iwh6����橇v<���ۄ��-"�u;�R�me��q�;ȅ��5V��#n����8z]�z�<r�'UV�lsn(���9�K[QEۉ�@�GH�UUV�U� ��^v��v��հ�#8mm �Y-�XG3����)��F�i�S��t6M�.Yv�<\/!�����,c��Z�nՓq�َh�hKv%m������	�n6�թ��)ڱ�L���v(����i	�Xα -ۯE�:�b�@9-�^v��we�hӎԄ��ѭ��1��Wmm�6Ѷү]V0��kO#ù	7���q�sZ�a�z�� 4�O������(~9�QSG���+D@� �!��x�;W�(��C�� �r_}�v�Me6��M��>KU CY]vG�,�,�<BڛnK@0qU�cs��Iv�B��m�.��n�4˱7��+q�+=�2(������Ç��Gd36�ɔ�ې����t��rt#�!��^��c���6۲'6l�U;v'n�ہru��N��p�\m�+���=oE��YH�Ƹ��k�<�g���k+�q'mH�l7*գ1���w��]�7_��W+d�k:4��^8ɬ���C��t���*�*�]�I��g�`�f���k�ٰ7۶��m��B_DD(^�>���߆���jT��.�356� 8� F�=q�_W����γ��}"Nmcr��/_�4�Y�x��@�۹��x���Ʊ�)�a�B���U����`o�mX|�D;��3@;���NE�@򾶀�"�� ���ږf�zV��4�`�v!.Sg��`��u٬�]���5v�um�n������,��\n�g���gu�=�j�73k�Q�>ޛ�%�ʪ���:�uSJ��fڵ��BN!BB!J�Q��û�V?oM���s�~���z���6�9bs�h�}�\s�T�|�t�� ��@26�@�^�@�۹�w�mXrP��ޫs��ꑩSCd�r�7P�T�|���=�����~�:����t�Fκ�ہ���|���n;Dc-�B�wS�F;/��o�����c}	�M҉��T����V��V�sk�#���V��Q)��&!L�N�X�mX����"��/�t9�m��l�T��=��`o�mY�)-N��A�B���Z��mX�Ǆ�c����̷UVD>�����޵`��a���ϻ�>�%��S2���U4��a& G5 䊐���^��:�Ӡ����hlc&�F�b��n��ûu���VRܭ�L��m�_�9���@8�� ;���S �@Jx���/Y�u빠w�w4������,x�n!����j��fڳ��7�&��}�6G
�r8�m,nB9�{�s@��1�b?�U����,�}H�yC������ugW�x�W�u빠w�w4ֵ�r	�O#RdS�,��+�\�1�G�%�}9Cr�M:��u�^$Ț@��q=�z��]��빠ugW�v,��f
b1'��8�}vG>T��a>��9����#���JF�s4���՝^�fb^���@������mQ���H��iXt%	$��ޛϷ���͵a�~�z��h�
<�LY (�'�z�9�	T�|��9����@$"����e-���n��BiیZ���KYk�M�e.-<���-uu���AGks�,k�����\�cd��%�D�q={8�a���6�����b3�M[J�NR��y(Y̲��`K�m2s��ӭ�}����w^�Kx�WKN���.�ըP^�Y�Ob���Q�9��b��L92������h�;�+�9����$��
�6KrL�33*��.��\j�`�um�q�p�X-H;d�-(����|��ӣun���q�6��3s�s���|��b��Grwr!��5$r{�s@��<W��;ޔ�r׃����m���1�bG 8� {���#bA�H�$z��Z� 8�&b��yD�/jʻlr-޻������|���<���>���|����"����2~nc��`ͷ��n�綦sT3H�7W,�b�k���m6(�rL�����uz��Z�w4��j�n�DӘG3@��^�+B�KR���J��Nk�3۶��n�％W��"x1Ǡy_U�H�� $��@y˻"�2��I&�qh���;޻����+�
�9�qɉ��52G3@�z�@I�����-#���X��al�6�M��W9+��s���=0謪�79z��귎�P�'�Ēq�cp�L�-g\@zc����H�*@GL��[��bn��*������BP�ݽj�ܿnh���;w<,�LF$8��V�m�=�j�U�
�BW{�U΁��ZzR�o�G$���H	0s��$qR���h�F�M9�s4Y��W�h���;޻�]��<��LS~tMt�;utn+��ݲ�r<;Ә����Ys�V֬��	7�<Lq�W�h���;޻����:����8�MD&��$qR�]�ͭL��3~����]�s������9�}~��-gW�y_U�w��h��Ēu���R��
!$�u�`{�y���V�W��j1�P �f�v��fDБ�H�$z��Z{vՁ�͵`{d͛�;{���-�Y3m�p��낢6�Z�6:,s1�63x6����F��bN6���֬��V�6{�t�;p	M<Q�ܙ�wu��<���+�h�]��|��ԉ�9��b�$�� qR�e�BFP#����v��빠wu��<���:��؇�HL�NK@>qR� =0s�%�9���`|c��8$,ZR*�X��S�0U�y�Beo.[��h�T�=��Eu�n���kA[����@7:�m�՟<��Gx�}�Ӝi	y)Y �q`nc��~�'���-2�U��\�o�K���'v�ң�����1�����ާlE�gk�p�.�ݩ��]�Hd�k<v^���!	�mD�=nY4�u�!�%ײ<��&�� �C�9�9�vmۓwZ�����s^`ض�ޗ��y)L�S!�8�c�d��!�cRF�h߷4+:���Z{�s@��$������ͤ�b�$�� qf�v��fD� ĤQ=��Z{v՟(P����:M�1�Ƀi��^�嗛h�*@6�L��ڴ�kp�X�G�f���j���u��t�;=�j�ֳ'c�����9ۍ��m��t�\%u�õ��n�8��8�(�1m%ݧi�1�Z��T�}����6�x���<���ؿ~����Q���"0|@x"�
��|�=���'����~�O{��"!��;wL�*i���:�v�u�=�jΈ�I��7���N�5�;Gɍ���"s4>W��f��2��+�����ZؒV%�`ԙ��郘���- �EH�*@FC��V����v�֩q�4lv����%��qqU���C����<WB`�(Mn =1�@>�R�0s�Y�b1(�B�h�{�s@����<���;�,�BdMc�N����͵`{d͛������
"a+J�+d�1�a�Դ����@b6P����H��3'0��^04%a�S�u!�bF'xI�5Uv �`�G�%"o� �=@@�V�"��OE����Qj��_����~�o�{ր�qR��!v�����9���^��}V��۪��C����o��It�L�R��X���- �EH�*@t��@~��~�?p��,������G�Ɲ�2h����_f^��.e�I[PF�<����i�߾�`g�mX�3g��^�ϧ��������8�F4��9�{�s@郘���- �EH�L���t.�S�V�Lٰ?l�:!D7��k@����ry�"hHĤQ=�~��v�u�36Մ�j~Q	W��W�U����Hİ�4��;�w,�"�����&���w]��e-�
�][�1�����m��Jӵ�Z���tj�T}m����������T�郘���- �EH�;ɷnݹ�r\�\ӒO���s� ʪL��������V{6��	����x�RɊ6�x���=����;�w4��^��T�[���B�-��{�ߕ���j��ɛ6��`Tp�s�$�#Nf���s@���l�;���nڰ&5BS	,�DB��ĎU��fS̻&̳7-�-2�eol���Y]v9u�il����̓��1m��up�����r�KuN&�ٳzu�p�*u��n ��kkU���9�bh���@[�e�]���݅���0Y�l�����8ݝ��m7`ӷ �(#��3v�����v �n��4'���V�XD^3��v�4ۯu��Ɠ�x�^�N��Ѭ��@�.V�Z�@B�v��w���{��ʿ:gM�/Om��m��Rj��MD콶�[l=�u[K�w:ʸ�v��]�}'�6��`g�mDB��0�޵`���b�DH�+�h�*@6�L��v�&ѸYV�T�sN��nڰ33mY�(P�t��`{���w��+�ǊH�s4�@t��@zd��}"�f&ݹ�sNd������ɛ6(I/uw?�^�����4Wg+�qF�K��ᘺY�"K�k]�H�m,��1R�g��� ��Ʀ(�(�1Ǡy]�@�m��;�S@����<꒫b<q`��]ݼ�{�����D����|�f{����@����+�h+ISJF�ә�`fei`{d͛?�(o���h��s@��!,����)�(y�oM���`g�mX�ZXa�<V`���D�@�V��۹�wt���gW�ZX�j@o�2���`��3m�h[��[]�rS��y-��4�Sxm�L�ۖ��nܹ��'}�`fei`{d͟����=���	�]5JeKR�j�jiX�����ٝ&����v{v���l�$��m�I4�I��Vt��`~��v5	jZ(IBI�B��J���ڰ33mX�c��U$�N�]9Rɩ��'��`nwZ�3��h�uz�RW^)��p�����Jn�~_�Γzl�;���DDFm=S�:���.�IJ�D6���9��A��h��K�7:�zɓ<o��W�ݵ�)��1'������nh�uz�h�]��ZؒYa�N9��&l��IBM������Vfm� �;�'AL!)D�@<���빠wu��<���Yˌj��BI�L�XDB�B�I)�Ｌ��Ձ�f{��^% ~
��<��@�וɉ�c�$MI�w]��Q�7������m�}��T\�q*v�hHlm+;�[<��vĜ��'�?w������O��i�]��y��;�'؀=$�� qR��K2F51F�G��= ��4���n*@z`� <��ŕ{FVm]��K���3۶���Vr�Q�Γzt߾�hS�I��BN's4n*@t��@�j��L��A$�R9�`{d͛�%��wW�7;�X����(_���Bj!!�"0!R+�|Ks>�2�fL����C�ɚ�Kv#\��Y�:2��NѰe��;5��nQsDضT�Lq�j��s�cs�l�KMl8<�q�'u�UBi�[N��L89��(�K�nݻV�hG���퇋�o�J�8��ٸ^���Dv�SYy��K`�,eWa��8�[�1�j��â�LXEk'V��B�S�@�q��/9��{���w�Ϲ"̫�g�͛L1�s��*�ezR3�����r�X�Wl�LS�JE#�{��h�w]��ί@8��5Q�K"�7&��ݵ/�
���Z�7�;�ۻW��Ǖɍ�c�$MI�w]��ί@<����s@��ĤQ6USniX�9��?n�X��V
b���h~��Rc�Q�Q����I5 ��H�T���r���%i�Kz��I:uJ����/X6b��*��? !�]z�, S���pb��͍��Vfm�ڧ5�	(���wU�̿'�A�bN's4���߱��d���5 �EHY&avU�?]�*�sJ����v�wj΅��u�wzՁ�{%9D�bu4RuN��!B�߻����Vfm�ڧ5���ZJb1,$�ܚ{n���s@����l�=�J5	�M��n���77i�ڻt/����Ӟ�x(�8������X��[�lX�I�g�[~��=��� ��<�u� �9�)DM�#�ͤ:�hm������}Ul��>�N�*��Ne53N�=��`g�mY1j��B�w�[j��S��٭)^�!1FӒh�w]�ڧ5�}�S9��U��;�?MMS�LI��Nf���s@����l�;޻���]m28�M<�8��c�]�ͻ�NIe��F�8�C��\�8��q�����n�y����r����|�w]��w<OA��&'�ym��$^�nh߷4.>��
ULo�щa&&��/_�4�U�[f�ރ�+��ǒ8ۓ4>�{�ߕ��S����ՅB���!	(P��dLD%{U�V�$��*]PK�����i�X�G5 ��H�.�I�g�����$yiƝ<%�LL�bn���kYn=m�zJ���b�"�̽{�u���=�� 8���~����hߒ_k�1'���6��@�z�@>�Rұ�@���ɛ��iH�ӚniX��V�S���g}~�����-lB�"�7�lNbұ�@�� H� �<X���##p��Z��4��恞ݵ`~�9��!/(IYZ&"@��2Oo"@b�`E␱�A���#�m��*%`���}`���ya���x�zkV�r% ^ ?�
)Z��� F1I � �-�K#��qRA��
s�&. CD�X�q�W�{�&��a.�ۄ�7.1��Ơ#c�Ɓ{EKnE����̩n��D��^X��e�K ���Y�f���Y��<�}���CK��AͶ�g��v�c���In�uF��֖���p�J�D7���n7Vv�Z��1��!�����OP0&�C��QV˷П�wX'e�Q��hm�;s5���l��Q�w^��V͹�A e�S@����朜��5���Q�۵�GJSֹ]u���pVL�n����Ep9Ef� �U�[b� �GM�Hul��n��QEr\[	�U<��ŝ�[�+3�cP9r�Aۚ�dڲ:21�l��9�-���X��z���s�Z�F|sVZ^���Z�n�t�]�ק����p����ZA�9݁`AQ���X6 �D8w��-u�郎��+/ӣ��Q�U����I�� l� 4�P.�Ml�!�d�&�@��F6ɖ����0�P���( ��Ѫ^k(��M���i8s�}?o�!���Dm�m@�M.� :ۧ[u�Y�瓌�+A�!����UJ�U�z�g�Z�*�T���2RR�#��q�	Ѷ�A4�&��;�=9<�3�jsn��<v�۬�CT�)�]��'�@x�y���t�k�ک0T@70�ҡ�(�TxL�r��˓��6��b� ���s�s��S�U*��L�Ir��Rkb���lj�Y�b���'I��+�)��j�-�Ʈy��OnMut�c[�5\�t
�E+R�U F�u���w[m����]�[�b٠)V��
c�)�,;�k���x�m Q������Y2;���G�A��W���w3�UR���4tY�$J[Ɏ���-���ql�|���c��֘��u�E�@*�t�Y�D��d-�Ŏ�e^��HtK�W^�Q��+m��/\ǘ��hw!�(	�����y�8!f�V훵l Hz�M3�{ 6�T���-��푴�?(E� ������PT?(���������,:����~���YLݛu��I.ݓMߕ_],4]�:`"vnayv��v���4��0����nΪ�р�ֶbƞ�P��Q�9÷{=�^��VU66�&Ԭ���Lv޻�*G-��\*���6�m�dv�-�jI�l�x{�ڪx<��ؕ��\�t��x�5��ݸ���d/�7.��Ӏ�7v��T��v����epp\���vQ�-��#��w�Я�&+�l�nrOm�u8tWs�λs��N��8�vz�ٍd/�ww������c���}��� ��HJ�- zI����x�I�y�93@�빠yq�Z�wj��fڿ�P��BP�N�N���u@�qH�s4�����-�O�J��s@����wT*�QLsLQ����ۻV{6Ձ��j��!��o;��o�%7iӑ�˚��3ٶ��F���������l�<��F�"��-��|8.��=,���>J�vP�5ga�ȗ ݒ!D�RF�1'�9�w]�ˏ��-�@�z�h"��%H�D̕#�V�S��W�rI/�DG��U��`wo֬��V0̔�'Ii��h��m zI��*@6��c����J�cM��9���I�o~V��s@����l�;�u�n4�<y������m�HJ�- zI��,�*�U�RFFC$�0�,i����YJ����e�l�	乡�b&���eGVə�����ұ�@�j������s@��/��)�c��cr= �������j���`jy�6h�-Q���e�n�#�R􊐿W�`UBE7)"���@��� H�#XLA�a���{��O=�4ָ��sI�"Nf�߿g���;�+���nmX���3vdczSLt*�&iX�ń���� �����n�}�(�!&D&��wo-j2�m�!V�c��+k1��º��F�	!����F���x�}��/[��nEH	V�� ζTͭ�*��Nf���ݵ(l��`r{�6�ݚ�|�O<��ܙ�w[��jy�6|�fwuX�֬�q�Թ*���q���..���٠^�sC@����#�'��I;�^�%�1̑�q�nG��f�����������qu�@�~��P��F��I3n��V4�×M|^hrC�t�n�t܍NՎ��x��m9&�z�������^�{m���\q8���Ĝ�3v���9=� ��sv���g��21�)�:M4�O{��=��g�	&�{�X�֬a�Bt��1�&G��f�z�������^�q��$	�brM���nw~_����lۛVID��
�����r]��R�IE!�Pl����,��V��h���յm�'�3���:8q�[G:ڵ�Pר"9�+��I�g�k��n����ӡ�JV�B����s��HM��,k���MĹ:;[�ⱝ��q����M�aö�c�gk�}=��D�:Ƀ�s�tsٴ{e���7�s�k	���S��ٙ��a�-�9��s�sSd�;w��׶�_�k�i����H�D!�!��V�b��6ݜN��_`m��w[+��<����~m����*ܘ�:9��T�|c��.JT��Ӛ�f�������"!��ޫ��Ձ�ݵ�ٻ�}6:�&���Q�nG���h���;�w4��z�U`�-�m9&�z��3vՁ����|�BI���<���4�RI������s@��נ�f�z����Z�'!�q���m��Е	�c�Zv0���U�l��5�q�X����..���٠^�s@�s@��Ӯ,C�#�I����?�_�� s�>����>�~�`jy�65�֦�(D�����T�nEH	V���M@n䭙�nT�USS3T�9B��{�ߖ��+��@/[4��h����HLM�܃s4��z�/��O ����z����u�ME�"�&7�G���p��st9����c�"��2
�2s��al[�4��3r����?%��w�,K���Ȗ%�bw��(  O"dK�����q<���2%��?����x]�]������bX�'���'�,K��oxT�Kı:g��q<�bX�%��w�,K��'���ffdܖ\���4�yı,N���ND�,K�{��Ȗ<���> ?_by�w���Kı>�߼8�D�,Kܗ���{v�Y����*r%�g������yı,K>�۩Ȗ%�bw��É�Kı;��
��bX�'�'��ɗ�w�.n��Ȗ%�bY�{���bX�'}�|8�D�,K��8D�Kı:g��q<�bX�'N��l�ٹ��y�VKvwn����umd�kc��B�s����qYk�uo�{�����-��gE٪O"X�%��~�É�Kı;�s�ND�,K�{��Ȗ%�bY�{���bX�'}�}ù���I��nfn�O"X�%��{�"r%�bX�3��8�D�,K�����Kı;�{�}��7���{����k�i[+KXb'"X�%��=�s��Kı,��ND��"}߾��yı,O��p�Ȗ%�b{�l��%�ɚn�d��3w8�D�,�D��~�ND�,K����Ȗ%�bw����bX�A�H0BHC������~�'�,K��v�~��^i��.f�"X�%��{�'�,K���9ı,N��q<�bX�%����Ȗ%�b|���s�����a+�un��k7�x�ض��t���g��A��o�w����
��I�˚z��bX�'���g��bX�'s��8�D�,K�����Kı;�{���%�bX��̔�����7v�9ı,N��q<�bX�%����Ȗ%�bw��É�Kı;�m8VBd&Bd,�̗27���75R��Ȗ%�b^��q9ı,N���q<�c��"dO��p�Ȗ%�b}����yı,Op��;L�0�%��nn�r%�bX�����yı,N���ND�,K��{�O"X�%�{{���Kı;���ܷ2L6���Ӊ�Kı;��9ı,N��q<�bX�%��w�,K���Ȗ%�bT #���㻿��;������^Ńև�Ui����܍J,��D�Rc�sd����M��-���ۣ7X�l8��䱮{nz�Hl�m�7Iwe�v���)��;���eXܼ��3@<����J��J���;s�vyv��y����x ��Zv�ܐ�q���p��t��d1Nv�rlo��n�Q���r'ZBW[�!;I=��ȸ�!a��n�w3=���P?��{�g��M0,Y���P�`X�[�;�&��y)8���nQ9��\�èiu���ٙ�Nı,K�{���O"X�%�����,K���Ȗ%�bw��*r%�bX���/sə����fm̹��O"X�%������Ac�2%��~�É�Kı>��§"X�%�����'�?�G*dK�����j�S4�SU
�L��L����Zyı,N���ND�,K��{�O"X�%�����,K��'���s3%�l��v�O"X�(�@ȟ}~�Ȗ%�b}����yı,N�����bX$ȟw�O"X�%��K�d��n�[��ۚD�Kı;�����%�bX
~�}�'�,K���}���%�bX��s�ND��oq���ߟ��}��bb��Sd��1�mZ�k�Y�g	�j�;�z�E���b-��m�d��仹��	"v{ڛ�V{2ըA	��J�!i	��g7f��%�bX����v���L��\���Kı;�{���AP���\r&ı;�s�ND�,K����Ȗ%�bY�{����(9S"X�vM�fn[�&wr����%�bX�v�§"X�%�����'�,Kĳ��u9ı,N���q<�bX�'}���:끩�n=�oq�������?'�,Kĳ��u9ı,N���q<�bX�'}��S�,K���d��K��vn�f�˛���%�bX�w��"X�%�ʊ���}��~�bX�'ݿp�Ȗ%�bw=�s��KǍ���~l}�9�X8�n��ۧ��Պ#�R�8ʹL˰�/IN����}�}�"����s�r�n�yı,O���O"X�%��oxT�Kı;�����%�bX�w��"X�%��Ogs�32�m�v��t�yı,N�{§"X�%�����'�,KĽ��q9ı,N���q<���+�2%�ܗ��K~ݬ�)���T�Kı>���q<�bX�%����Ȗ4����aR�!U�.!���P4����"���PxrQ� @�0	%�!�"�����ZM��x�G��1b��%"I*a�!�+���H A��$Q�R:��{�7�+ BV$cD�H�H�RH���
��(��hD�$�!2�i�hA�H�D��"Bʡ,	F$@�
F+
B�ba�	BD�����\��V@��
���@<����,�+��X)��dX�� �D`ŋ�#�`14�$�e� �BTeT�H��R�0��DH1� ��,HF��$,@������AZ@�x(`����	�?�E¼U߄zv'bg}�É�Kı?{{§"X�%��I�p�v�2Ysr]��yĳ�PX'��u9ı,O���O"X�%��oxT�Kı;�����%�bX����N��a&Kse����Kı;�{���%�bX
���
�D�,K���gȖ%�bY��u9ı,�~�?_e��ͫDz���u�"���sI���&�e�9ggŇ��A�{I��,���Sst�yı,N���ND�,K��{�O"X�%�g{���Kı;�{���%�bX�����˓M2���ۙ�ND�,K��{�O"X�%�g{���Kı;�{���%�bX���
��� n&ı;�����+%jVY���oq����o���^�X�%����Ȗ%�bw��*r%�bX��}�q<�bX�'gm�w��.,�ۗ7wS�,K����É�Kı;��9ı,N�{��yİ:tU�]E���L�y���Kı<���;nfYvYv�4�yı,N���ND�,K�����g�Kı,��S�,K��{�'�,K���w9�rnmɹ2�-��ss�]q�9��<�c�p��#wo)Z���q�3lK�
�`N�n=�oq�������s��Kı,�{���bX�'{��p?��ı>��§"X�%�zN�.>�p�e�ɹ���%�bX�w��NC�U#�2%���}���%�bX�}~�S�,K��w��'�,K��nBw.�	2\ͷswS�,K��{�'�,K��oxT�Kı;��s��Kı,�{���bX�'{'�÷4˖K&�ۻ�Ȗ%�bw��*r%�bX������%�bX�w��ND�,��.���������oq������k�4������T�Kı;��s��Kı,�{���bX�'{��q<�bX�'{���,K��C�`Q"!￿��~�� �Ʒga�]+A-a���\S)p˰vz#s��C�e7g֥���k���3�-���r�`�-��)�9l��n���(��WO^�4�[L:[\�y�:QJ��m#$��vc�97g�[kh+Eۻrh�+��N���÷}��$�l���i9V��]:�m��9o7"u�(e���n�Ġ�SgX�r�TR�Ѱa�e�����ANӞ�&���+�ݽVn2n:n�����nطn���J��͊�0�fJԬ)S�������D���S�,K��{�'�,K��{�"r%�bX������%�bX�����[��l�3n\��ND�,K��|8�C�X�L�b}���'"X�%��}����%�bX�w��ND�,K̟�s���)�݆e�8�D�,K��p�Ȗ%�bw;��Ȗ?�*���,��S�,K�����yı,O�/s%��me�Mݹ�ND�,K���8�D�,K����Ȗ%�bw��Ȗ%�bw��VBd&Bd'�̗:�jf�H椩��<�bX�%��wS�,K��{�'�,K��oxT�Kı;��s��Kı;�nf^l�wn�&f�i�{nhr�+��t�!*[-㚌skj�<��%�wm��p�%��w7u9ı,N����yı,N���ND�,K����<�bX�%��wS�,K��d��v�r�I������%�bX���
���r
�z��:��ߟb{������yı,K>�۩Ȗ%�bw��É�Kı;��\ܙ�vL��svfiS�,K��}�gȖ%�bY��u9ı,N���q<�bX����Ӆd&Bd&B�k�"j]QU9�s7wgȖ%�bY��u9ı,N���q<�bX�'{{§"X�)���z\/�&Bd&B�[n���ʢ�͹swu9ı,N��|8�D�,K����
�D�,K�~�Ӊ�K��	��U
�L��L��X���fh�E��.����C�cv�<Q*r���V��r�l�+\�&Lt�V�����q�ı>��§"X�%����gȖ%�bY��u9ı,N��|8�D�,K�K��l�ܬ�d���*r%�bX���vq<�bX�%��wS�,K���É�Kı;��9�*dK���,ϳr�$�sr�l�yı,K>����Kı;���yǥ���CND�Nv��ND�,K����O"X�%��܄�i�	,��n��"X�%��}�Ȗ%�bw��*r%�bX���vq<�bX�%��wS�,K��{�;wf\�Y7v��8�D�,K���S�	���������.�	��	�}�T�bX�'}��O"X�%�O}��͆�]n��ɽ�Fm�`b�7mJ˩O� L�+A�,e�ul����{��bX�'w��O"X�%�g{���Kı;���yı,N���NOq������|�l�Z��j�{�Ȗ%�bY��u9ı,N��|8�D�,K���S�,K������~���q�߽� �ok�����W�D�,K���'�,K��oxT�Kı;����yı,K;��"X�%��Oos��e��i�33N'�,K��oxT�Kı;����yı,K;��"X����j����s"^'�,K����2[ov�[2n�f�9ı,N��;8�D�,K�O��u<�bX�'���O"X�%����Ȗ%��]�7�:�UJ�2�:U""fiUr���v^2��T�Z̽1�����]#+=�32m������~�bX�%�}��r%�bX����yı,N���ND�,K����O"X�%��܅���\ݳswS�,K��}�Ȗ%�bw��*r%�bX����yĲ!3wj�Y�p���]��+�Q.Y,��nn�O"X�%����9ı,N��vq<�bX�%��wS�,K��}�Ȗ%�bw����36M32n���ҧ"X�%�����'�,Kĳ���r%�bX����yı,N���ND�,K�ݲ�;&�����͹�����Kı,�{���b2ݽ�p�Bd&Bd.�֜+!1,K����'�,K���B���!�s���v{@��e"�X��P�I����f���oe��9�:�4�<���N���1�u���UC���y$wY��׳��{���v	�*��ԽB�6�9���=/��9M���m��s�ܦ-��]<���Ů��bE����c�o�n]���y��(F�n�vz�)m��g��WAĕu��&)�ܷ:�B����o���sKL�sI��S�G��«��=�tʹ�&:������E��F�O;���"��^�j�6�ut= ���XE�����%�b}߼8�D�,K���Ȗ%�bw�y���~��,Kϻ��r%�bX��v��[�������8�D�,K���Ȗ%�bw���Kı,�{���bX�'{�|8�D�,K�K��m��Ylɻ��T�Kı;�y���%�bX�w��ND���Dȟ}߼8�D�,K�}i²!2!<G�Y.^̴SNjv��'�,Kĳ���r%�bX����yı,N���ND�,K��{x�D�,K�=���fae�7l����Kı;�{���%�bX�����O"X�%���߯Ȗ%�bY��u9ı,O��s;�7eۺn�=��t�������V��ږF��<<�4R�K�mݙr�ٛ�����%�bX���
��bX�'s��8�D�,K�����șı>��xq<�bX�{����0�]r��-ǻ��7���'s��8�C�W�*�� ��Ư�<�bY��n�"X�%���}���%�bX���
��bX�'��ˮ�����8Ӓ=���������Kı;��É�Kı;��9ı,N�{��yı,{m��ٚd�3n\��ND�,K��|8�D�,K���S�,K��w��'�,Kĳ���r%�bX�d�{����Sr�fe�8�D�,K���S�,K��{��Ȗ%�bY�{���bX�'}�|8�D�,K���|S4�Ea���fs��c���	�m�3Y��]�Rt�㛸-c/��}. �c��n<~�bX�'�}���O"X�%�g}��r%�bX�����yı,N�{ª�L��L����r�e�T�uSpyı,K;�wS�,K���Ȗ%�bw��9ı,N��q��{��7����ߡܿ��8�N��r%�bX�����yı,N�{§"X�?�P�C��@O���'�9����'�,Kĳ��۩Ȗ%�bw�=���.R[3v]�8�D�,K���Ȗ%�bw=�s��Kı,��ND�,�>��~8�D�,K�ϧ3nfi��ww.�9ı,N��q<�bX�%��wS�,K���Ȗ%�bw��*r%�b��?����
Ij��r-v�]*������ݭ��]v�'+�;�1?�_|c����\��s7s��ı,K>����Kı;�{���%�bX���
��bX�'s��8�D�,K��w�m�sL�.ne����Kı;�{����ș����
��bX�'�߾�'�,Kĳ���r%�bX�d��;s3�2ݦe�8�D�,K���S�,K��{��Ȗ?*�2&D���ND�,K����Ȗ%�b~�{�-��k)r��f�9ĳ�C���?����q<�bX�%���۩Ȗ%�bw��É�K���v��
͉���9ı,K�wن\�fSm&nK��O"X�%�g{���Kı;�{�Ȗ%�bw��*r%�bX��{��yı,N��NY��3]sϪ	�wb.��\�uk%���]�Od�/;Bf�.�nGp��e�M^ﷸ��%��{�8�D�,K��p�Ȗ%�bw=�s��O�2%�bY��n�"X�%��d�0�4����ݷwx�D�,K��p��|+��,O��}�O"X�%�g�}���bX�'}�|�yı,N�vs6�a��2�ݹwH��bX�'s��8�D�,K����Ȗ%�bw���'�,K��{�"r!������~���"�2-?{���ı,K;��"X�%��{�8�D�,K��p�Ȗ%��ȟo~�8�Oq��������qf�+(�{��,K���O"X�%���߳�	 �'���NA$O}�tI��TW���TW��D��D� ��������
���"
���"����!� Ȣ�2����� �* ��("�0 �"�1� �DUG��TW�uTW�AQ_�AQZ"
��(����
��ʈ*+�� ���(����
���TW�*+���
�2��`n@�Vn�����9�>�A�e 	T(J��R�$�*QT�*��D*  )U@ ��= PT��% �*JI
E(PA�TQT*J�J�$�PRH!*�QA@ 
   
p   � � �)��_|�y��#C&�g;�x  �б��R�l�(�&�U���%)N&�R�YJR@
RݹJQW,�R� ��!e��)e��)��)R�)JS �r��14IJbiJR�)JR�)JP  �   
@� �r��>�t��,�$�Ye)B��JR� zw)JSE)LM(�����>�w :OA�� 91�(Qr�
(P�>��(Q�'�d:r^�A׸����W�X�&�u>ۛ+�x w��@
    	� ;}���e�����T� n���kk�*��9_m�j}k� �T������x�v��uUp �[��.m��������8��T�ϣ˓_&����}����y|5   � P�� �}>�=��6���5L���@+���z� }}Ņ`��)\��F��U�y1�p >����OG�_Z��u=�_1�X ��4ɯZ�i,m#�y�J @@ R�pK�W3ӣ�j�iV1����p�������{ ��4�� y��t�-�����O��Y�/��O[�ps� ����7��a��ɥ�ː������UC#���D$�M� Љ��R� CA� ��U*��UC#�������JT @Eڤ�H����~�����w���VL��f�7��@������**+�D?���**+�ਨ�AAS| ~O��'����{HD�G���i��L��noZ�c�t���⽾(����dɐp��T4B�!���N<_����s�i���|4�5�a�ƞ��d��G�6\3`�ɓ27S�lnx�Q�hP20���6P��J�
�(;-��s�t�xq�0���S�������g�Y�r����r��2r�{�9�vt�d��R��9���ȅ�P��xk��p}Vp*!�tclJPL�3�1-�j���i�}�`���M�u�w�wxt�r㌗'.SB��������h 8�'2��qΝ=��C04�G�K�����9�]�x|�c�$�N^�¤�|�|�H44��Ӵ����D��.��ד,����ܱϏ����`Ȑ��"H�Pq��|��;��rcN]��}�n8������BƁ��$�P�M}�u���;��~�Ã bB�`� ɠ�A#H��w��!�l!]0��'{z��z�M��)��&%�"o~�yG(�
�z��N%|�jh�N1����e4F;���]1�6�����H�U�9�T�P���6®��:��[H��Ռx2�|x�
e��&2�L|�\F=�:x4g�|w>w��Δ�Lr�!���n�kG�n�P�Rl��Ռ��ks������>&Dü[�n��!u�ĉ �XH�u��t�l�� �r5d��#I}�I!���5�>��R��bc�CJ*?)S��(��
�щ��`"A�*@�D��qJ5.N�=#�ҧ1�B�����59��{���x���k�y������}�\���q��e�.���~�1z��#��5
8T�S�(�P�g�w9ӣ�s�x@rh�<�������Yp��%��:5IJ�v©��J��yy�|�<NT��X?yw��Ĝ��x8h���Uby?z�C��!�� E�HP�T�a.���æ\�V��pk�2^�4)8̝N%�9}����:w���G|π��0僗�s��{����H7#�w�^n��mڜ\�Γ��4�_~��N7�'��y�9��WN|e��Qѡ�4hb$	�X�"	�@H�4��E��R+��5 h4j7I���b��˃!RB���Mp6��0`�2*oNtyYFA��A�CI�0+ �D�#������y8��4�k��|�kz��>�0k��Ns�r�r�2q��S4r��58�x�����Ⳝ���{�ݕC�׉�q���*����5�dYR!A�IX�� C@m*L�2��!����������tf��aQ3Ȇ�{��k��'y���58� ����^}�l�>�j�"Ͳ�aXЁ���U4��y�tޮJa��
FƄ����b�b�E�!H�b��rk�O�>qoX7:���Q��!��i
�E�: �>ﻜ�$SP�uR[��aIt�.�T64�băқv7&G��]�q�3�+�8p� B�
"A*� �c]l��2n�I<�p�L��8�B��^ؑ�ß��:B�!�١!�_$D�D H� LD�ќ���+Sq�Z��Cd\-{T��0c�n���T��m�"�m�&zr���p��ȗ2���z�����I��*�P"��x�7:q�s�__E09F�'N�Q§*P�1a'#%�b�M'+���UB�`�m0�s���˓��ݟwo�������9���S����2	�c%�:=d�����N��!��NbB�(Ah:g�-4c�c���/6;���tL]�����Qâ1�D��wPL�T��5®#�;���1>�d)��!P�V���<]%ɉ�9Ӝ���B=�I
g�JD��&U6�L�:9rdk�P�⭧S�40� c����X�$�T��2SPe+^'9�Ev:M @��4i)��E�5���C���DzN!
h�Û���(�����&���hp�0�aO�/N&�I�]��EL��ɍ˦
����!�w���6pI�&nT�ǯ�r�B��'(�O����I����v�ڏ\��jJ"*&3]�����|������::F�%%
i�T�.�K����6�"�]ih�Ƒ����)t�)�f�m9n��a
�.�
�2M��.�C��U�m+������/xsǩ��L8dԣ�p��p��4S�9�c�����#!��T����o����S���a�(�\MF��@r�k��]V#��K6��*B��42Pr�J�
�Q4D�A8n�Hp����3%024�A� �"������d�V@4��@%�`���@��2�`5"FH��Gk1b58���T�$ �c�;P�"^H��$(I#��v����pp$i��C��@q�5SP��R.�IaR$l
��I�0�Y)�s]���}ξ�geNs���'��o���/[p3rnz�y�7���9s��=��}.�������fg:n���s�W�u4#_�!
�JRM2B��s	N� A(�J
B���	f��M4jZ�B��B���"H!
hH5�;���)�N�! 0�D$��!X@�V	H�C�$��������~zI���~�����o�9�<����C%�����wΆy5��{�C!L�%�z���������c"g����ёy����Ӡ�/9��T�h�5s*��Ύ]IW|=k�:����c8&Gw��yn���g��Ww;�~A�<Ó��7�pZ&xcEPA|����7�:P���B��(i
�yļ��G������X@d-��L���!�����V�rʜ�&�!��8tw��w�{�˂�v��90�d��N�hd�-D� ҵ�F|�L�D
a�)�7���N�j*�e8>�؛�x���/RPib@�$��޷;��|pbBbŀ�4�
�F�` ���t�t*1J�(��,H�,���g�peX8K�71�i. ��]a��12�a�铇�\8&Lq(1²��pbbd���xWN�&J���y���p������<��U�A���t�CK��B^+��A��� jT��pO4�:[�� LQ�4��*�����>�0�k�����	��|�F��%ɔ[S�z��g���qQ��)�ȼ�p��H�+�dC��4�
Jig�M<�-���ȀƈgO�9�O��/! #h%RT�� 6�&P�;�xo�����N.@s�Ȼ�{IA߹q�{GZSc���N������3���%��ׄ�����=�({w��������Tsra����%��{��/eo�'�rb�X�^T2g{��^�.��N��y��9��/o�ގ]�^;��a����ǣ.����5 �q�FFFK�cd�_� T�B[��B0 P @#$`bX, B��D�c*�� J@��R��`�]Ӻ�i��H�S��]=Xۇ�k�cD��`1(�҆Ҭ)M;P�Ѵ�Z���Hl��D��[���0�M	��C@��B�m_�"R�.(�U a����N�k��M1+��DhD�wDFx�'w{�k�k �"��b���E �E���� Q"��A���R�5�A�M�
��� �XN�J��a��a���� ,�DXjU�%�>��C8�:�5GDJ+�!ua.���N��Л���P*iX�e��R,j�WN�4ºa]1��d�r�(ѵ�Fd�}NC�H��t�!P����D�?x����6
y�3��m��m��` h m�� m�  ��l ��[z�:��f��T�����eBۦ疨m{E+W^�B^�~��[�öY:��u[��q&��ؑ k��%X�5��1o��}�ο2q������	 K) �t3l����� �wb�@�L6���\�*�ҭPPtj�`���ڠ.�uاJ\�M�Am��K��    m��ݦ���f�r��G  [��m �-H 6�� ��  2� ;m�lnۙ�tWmUUPR��^�ZW i69z�ck�/��t��[Kh[@� m��n��ڴ�� 7:�-��oN_I]6� ���v�7�Vƛ#��kڪ�h�n�ֽ�Gj���p�V�Q�n�@ �X�a@��:� �\9�j�v�i�@p qͶ�%[��n�M>|��$$��0*Պ
�v���j�������)��ۆ;%+E�m�H  �l�6� m�ͷd-YԀ�P*ɦ�,�m��䁶�p9�ڷ��"�vlP���7'2�U@]m*��˵R���mSi�^�Z�l�H:� uT��J�q����-��� H -� -�l       -�      $  �v $ �O��䀶���ۀm��@��{N�f�n�5�  [B۲�*�UT�+tdތ��J���j�v�$Q��m�\ݖ�\pm��$�4_:K�[WJ�T��,;e���٪;S*յJ�eU������ꐐ ��۰ 8m�[% m     $	     8    �     �l6�� 6�  ���	$i �m��  ѵ����m�%��n�ron�m��hr��ɚ���obƧ`6�ҡǪ�� H 	e'N:ε��jVV�����ڸ|���Ŵ�]�Q{t�o,�մ ��G�}��-�h [Rն� p�cm�R�q k���Im�hԳi˚�&%[V���0G]�.�$P#��� Ǎ�gX�l�X�ە��m�}�_��3	  	욽W�9�sm� l� �` (�
����S%/)K�v -�ӛln�,^Gk3�����媮����vU���h����9ֲ�7I.ؐ[G  h륝�^�TW' ���ۣ��v�J7mX� �㱷����� -׫tK�&��[VK%e��6�Vۀ�g&�t{H����!�\�ĵu�U���fЖ�e�rl���h���7k@��k�7��4���U�Wy�����:[�.�u7J�Ô' &xxYW�d܆]�3�m�g�ڭ���Ch M�����X�����U�0Xx်�W5�Q�N��F�)�d�kT�F�l�㛶�����;j�k��Co8O\�I0E�v���;c��� v�ەd6�r�5KWW��l�����_m��Y2ۀ s��d� ΝM�q�gE.�[�k�yj@cW�K kX |	��6��Z-�\v�M���������  8N��v^�}��m8^âj�8��8j�,ud�[��lH��m��JçN�M��&�YƑ�7��-�z��A�ͻb�	8�m�� �$8	ݲ�;m���A��V���W@+��m����	ܰp�m�ų<ts�X%N:j��Z���0��Sn#a궫��&U�V��r�)  ���m�$��ޓ6H $��L�d� $���H��:`�`8Hm� �
P�&m�m���$ �m�e�]�i\�Ւs���0qW, ��.�UM��:$���Xg4kw H��ZM�����[p��v��')l�o96�mM��
�^1nA��ka1����n`HH�[S:K�	F�uW]!m��6�kjB�$5� H�mm	ft�,�`x6�&3k�-�-�lI����s���H��z����GR�-� i�(s����:�����Zn�6�az�([@h�6v�F--�kg[[4� �`���
tW
��A��7.�$-��G.��5V�݃m�8  	�6�qn��[�� ZmΥ@Uj��]PE�?NͶ�v �zJd��p��U�vJҁ��^_���ȑ $C^�\lכZ-�f�z�m���h���q��H�9���.�@����cu�!�"��]����+�Sq��EU�.���gEt�D�М������
��HvM��m��
�UnZ�8��e����Ҳ�^� sm�te�v�X��[U�c �@6[��^�{� nm%Ûk���=�L�˲p2�[VR�\,;7�WR�U;�=)b�"4�N�3��@m�_W����cIS�����}�hp��ڎ��,���h�Ԅ>��@�ܰv,5׀y6�M�t�m�(��j���n�K+��(�f�76k(Ʉ 6旗�V��v�6��[�B��Yy��B@�� [E�i5�F�m�ѵ�p�h��̀��bE��}�� $�u�E�mK%�-���y%�۩UyeZ�ۊ�����st�U�wdȢ��$�b@��m��H�s�����'�[�mt��� 8 Y�$�Q���.�  �L� ���=
�Z�H�p�i6��\m��v�� �a��F���R��uU*ҭ�wca��U������ꪶ���  M�ܛm�ě}�ﾶ�l�-	0H9�f�
�[v}�F�����p���ڵ�	6� �m� p��BS#sd mv�U*T���XU�
�˳@UA� 9%�BE�pwm�l]mUUU_������ʽ$��^��*��vŷ���u� 9:-����޴�[@      ���[q��  6ٶͳm��cC�rƵ�u��We�
�e]������'Ch���[Ӥ��Z�H   H�@n�Y]���X��[`m�z�HMS�Px��1���se��+e���S+T�*�(�if���kpknݶ��$�-��V�
jU��Pl^�U*@����Ѷ��� �$��I���m� s�$,�fݭ�k��M-]>]�ڥ�s<r�����+�v�Z��U�j��h{-ӠqAҭTp�wsh�v�ˢ0bڀ�L�v�HVLdc��mp��O-p$�l������M�R�m �   j�m�x��I-�n�wj�Z�g��������$8g+��j�yW���X` m��?���[FҨ
�U]El)��l�1�m�M�75�;�z��T�F��@ImpH�'@�iB��U[�7X#H�l�oUT�8�Ҷ�  M��nQ��� �l� �-*p6�c�z� �5[n��6�a �#m,�  m[�KV^.�*���`uͳА� 2��PA\�q�*�[\m� "@�����86�l�	�$�L9�n������   ��   $  m�`f�m�uT��UR�۝��Љl��-�  �`km���� ��\���l �ړ� �`  ��- �h%�	�kh �    ��%�J6�hp  H �`-�G p  pIm6�jSjڀVV�U��j���qÀ 8ڶ  H�-����c\�  �[V�M�i��`���l��In�d�&�'�^� m� �   �Z����| ��e��`q��\�$	�&�m��H�බ^��    o M� ⶢޢ���S�Z$�m m������v���)�ݲ�    �V�R�a�P �j�VU�(-��]���6�   ���m��6�6�9[ $�-�����h9 �� �.M��[  �6m�n�:��u���m� �m� [\�� i��$��j��.@ � ��m��d�6��^۶ z��6{&�[@�%��    �Aa& $-��޻l�v��	m�   -�3��2֝Ki�+�5��	�m2�(����㭽J��($�mj�vV�(�����ԗ�҆�[�g]�nč�b�m�@ ��������!m   -�� m���m��/����mpml	    �|   �`     qmm�h��m���m���8>m�[x  HCm&�E�Üm�` H6�m�� ���L    �i6    m   @�Ć�Ll( 6�h.�m���ҭP ��[umAI  m�	m��l� �l�@-��v�-�Ӊ9�Z�6���N ��` 
j������� ���d���9o$��EoUWU*�T�Ǩ�e+5M�M��( ���D�r� qG]��¨b �Q?�g�h+�Ƞ!�
��P�A��B�P٥4�t)�@
>_Ah��bl� QD���Qۆ�b ;'��8TS����&��DW�����
�E XQ�B1RB
B`������� p�M&��<<At����ʈ�����WH
�U/@�@I۰��s�/��Q{��UҊp1�SR�1T�A6B )�/E*/>Mm�*���R,�iRP	��qu�'���@
��� lCO�������yAF�S �UX"w@ �E�X�� @���EEv#����+A�3z֏oO-U[e ���j�%�l֞��C<[i�W
ىw��v2���,�y�MIUlb�|L����Z�Kv7����;����ێ�;=�C�]ikgv�V*gN ���l��x��ڸ�C]N�6N��,`����!<�i���).'�iz��4/	�K!�XKF�cm�#�m��$��-��	9U��L�!�p,\�gF[����rJ�����E�:�oGm�<v磛�І�՞��{0���P�;sl�;�e2v��.�M�1��u�D;K,�n-sj5o�����)�7�v��[n��U��N`��9A1����]ÛRV�2�L��+�OgdiH�g�:���l.	U��Qr���b�9��1(��`,��{u���c��#�F���9��`x^�)��L�N�,;n�f��u=]N�t��q�+f��[ \�+C��;k"ht�Ή�jN��35�3ԍv�����y�t��L�u����ln<l��֌<<�h�"���.;Kٺ'nz�|�V{(`4��n�ue�k��Nĵ�P�C�����ڇ6T5f�!;r$�h��H�y0��,�Nۗ,�r��6���탏l��:Ȳ�;p�9�F�x�6�<,ѤG�Y&��ayX*Y���<��n�mO(���ƥ8���̑ V;F�	�v"�땺��v����D�v��.3\u��k�W(r��4lʽRT��Gv�&K{%��h�==�û�*��g	��v�M���rgj�U�e��$�nIA�z�NJ�эΦn�]����*��6%��+N��\k�	p�UTQe�[�R���-EX(�v�v��y̭[�Ll$�9�:����ɱ[n��@Tv��Y�SU������P�*�ٳ�!���������ɋfK�۫jM���k��Z��t ��6S�m�u������d
%Zm��X6�]���an�Fu �ldRk�6��s����!Ā�
П��'ȃ���Q�N�|��G�,>֩��.�s�Oc�>���&�iܹ�k/ '�"�v���v�1�xq����ĺe�q�68�*\�'\���r��1��6�;jo6�6�Wh)F\�����°�/=<�����Sv塱�2��U��# �*��� ��]ʔ<:+�:�rFp{d͖��M�vZG���V�ؔl=�]ls���n��&�k��B��qը$*����[�R�GX�+p�����6<�<'�S��x�
��	�B��1j�y��S@;�/ ���DL���I����p���.��ʫ�@>\��1T5iր���)�~T���m)"�E�����;���oJh��4zPj1��x@�ŠwYMޔ�oRhv*�U�~�Ʒ�$7"m8h���{z�@��Zu��?{��}��p-����	�j7N\(�!��=W�x����`�)���P�N�*��oRh��@�)�r<���h��R�.{�����9D��x���b�@R
QT ����ﳒL�o'$���&��g��I�4�Zu��-�M �ۓ@��Z��+c�2*�,̼�.�k�m�h�u�w[��^�ErG�8�X��ޤ�-}V��n�oJh�Tv4��Tc�����I6��j5��zd������1lg�v%��N��j��o���h��h���{z�@��1��(���@�s@��4�Ԛ���?Z���QĆ�n]���#4و���蛚�]�^��?ew*Oy!jI!�ޤ�-}V��e4zS@�����2�8M��h�S@��4�Ԛ�YRx�i/��O���l;%�l#q��{Wg�e�d�We�R��ȗg��a�6G�-�|h���{z�@��Z��u��&I�d����T�3@nӭ�b4ʲ�aopXƈ' �ۓ@��Zu��-�M�sn�b��y��ZWʴ���F����L�l�1�D �*���� ����Z�}(8��c�"qh�S@��4k��k�� ���+�ïY�q=�3̗9�:�pka��s�>�-��6S���ع&��m�����~�ۋ@��Zu��?b�*m<�B$ԒC@�[q���@�)��w���H�2'1����)�[Қ����e�M\$�l�-��h���{z�@��Z��V�2FD<I!�%؍���4��k�w,F�J����H�(��!��]	�F�1"&��XE#aJ�@�Eb�i
�HDI�����ɶe��\n���.��rQۑ��Ia�NY�Z�H)֡�����{[6�v!�{P]��z���N3�8�X�X ��,nv��oF')��ek���ڬܶ���v4 ��u�5�t�=AYv��r�w�۳�m؃�Y�v��e� i�́��yU�833�Lu%�b�<keu��uqJ�Fa��m�n���u����]D&&��l�רN[�]��Rt�vO鼟}��ѭE�˂���	��u�z�)�wYMޔ�?+�7f�Ӎ�M�	�[Қu��-�M ��&�oK���qx@�ŠwYMޔ�=W��_U�~���Z���6�4zS@�^��-}V��e4�:��`���RI�z�@��Zu��-�M��
�5	�<f8A3Z�.ۧ;K՞�w��]7^��F��َ��G�`�2D�H?�}�-��h����G�~YxI�O�a�6G�ܱӱ3_LL����+�F�rH���hڑ.�R	<I!�[Қ��M��h�S@�VGa��c"Ng�}o��>����S@��4���كq4�y�Bh	_*�LL����mc4w#4��������&Azw]��[���W�=u`ᑻw#u)x0VY�����'���Z�)�[Қ{�4_U�~��-cqĆ�n�)�g�y�fU4����M�&(��1���b�#G�9��[��=%�m�G#E�b_g�o�ؖ%�`潗iȖ8P�Q1P �؜���Nı,K=��ND�,K��.��5&�����\�ֈ�#�ߦG#E�bg��8��bX�{y6��bX�%�{&���bX�'�٢]atJl2�^�dq�4F����s��u�4X�{y6��bX�&k�ɮ'bX�%���]�"X�%��e��kT���6/=ljLOnDk���W`�|O%�;{Π��]Sg�)��J7n�>#��4F/�y6��bX�'s~�k�ؖ%�`�^˴�Kı3��N'bX�%�����B�L��#��4F���k5��?1�MD�sY��9ı,O���Ӊؖ%�`��ɴ�O����h�_G?_ٽ���M���u�4X�f�M�"X�%��g2q;ı,�y6��bX�'s~�k�ؖ%h�^����4t��7��#��O�5������Kİ}��ӑ,K��o5��v%�`s�TH��Mro��ND�,K��'�}�]t������u�4F���o&ӑ,K�﷚�q;ı,{y6��bX�'�����Kı)�~~y�u�v׹�r��:�B5�:�7������f�;WSmŃ4Y��JlV�*�6��bX�'u��o�ؖ%�`潗iȖ%�bf{�8��bX�&Oo�Qƈ�#D���m��׳�gf�[��,K��{.Ӑ�(��MD�?~�~�Nı,K����ND�,H������u�4F��纲K�p�]jo[�ND�,K3����Kı2{y4��bX�'u����,K��{.ӑ,K��e/0�[���nٶ|GZ#Dh�?wΣ��4X���\Nı,K5�ND�,H���s��u�4F������2�Y���'"X�%��ߵ��v%�bX~���ӱ,K�����8��bX�&Oo&��,K��_2仆�v�x��x�]X��a�m#�.�b%r���Jv���>��9�l�v�m�9ޛ�!�M^3؀:x�lf��$s8������N�Uts�x�:�N݌�`6�6ƨ�t=���� �Ӹ��;���۱�CWz����8�f��b�iSj��*N���gm{k�gl�c�0���:�F�:m�Wo`�s��@!=����ǭ�m�~�B	�ݜ��O��nXZ�7jޥW��uH�� ��j�
����%$9mt�2�Қ9u��|�#Db����h����g2q;ı,L��M'"X�"4w����h��1}��wG,��ZLޗL�4F��>��|���F������r%�bX���Y�'bX�%���]�"X�%��e��gu.���ͣ�����F��>~�G#E�b{^�Mq;��5Pk?]�"X�%��߹�q;ı,O�]��֬rR�Ie�gQƈ�#G��~w��Kİs^˴�Kı>��N'bX�%���ɤ�Kı.|eֵ���g�ν.w��Dh�����#�%�a�������Kı?L���Kı3^�Mq;ı,L�G���ؖ9*n��6�u��'��ώ���:q�g*kj��sN����Ⱥk��Kı3�̜Nı,K'��IȖ%�bf���v%�bX9�d��Dh��Ͼ���˝�I���i��Kı2{y4��N����H�1:�i�ND�3^�Mq;ı,k2�9ı,L�s'�#Dh�^�5�=-q�:��:�4X�%����k�ؖ%�`潗iȖ%�bg��8��bX�&Oo&��#Dh��9>f��k�4�l�֋İs^˴�Kı>��N'bX�%���ɤ�Kı=�{&���#Db����;�����.�h�,K�����Kı2{y4��bX�'��d��,K��{.ӑ#Dh���G����n⽴�[.���Y�y6�=�o*�g�åևM��LH����%�W.����۟Q�Dh������ND�,K���k�ؖ%�`潗iȖ%�b}�̜Nı,K�sY>�7%.3��yh��4{�{&����#���`��~�ND�,K߿s��v%�bX9���r%�bV����ύd��g�z\�ֈ�,ײ�9ı,O�9��ؖ5����b]St&���M1���!�2&�v���"��魪�"͛T�H��@�X�$HA��(�D*L��&��I*���@R,����m�oZAc�l�)���!@�P*�.���	���	���:!#aHTt�t �
���Љ�_�h$	�;�1�4�ڡ�l��@�HǍ([BV�"voby��τ w�
Z<>�T/ʆ 'Q`�Aш#��
�Q�������3y6��bX�&k?~��v%�bX�z�c��1�e�]28�#��j'�~����Kİ}���"X�%��{�5��K����~�ND�#Dh�������[\�nmv|GZ#E�`���iȖ%�a�c���5��%�bX9��v��bX�'ٜ���J�#G�>�>O��9tĲK$�D��wc���B�yŮ�Cд���҉���wm�nCK\x�Bg62<h��4~��;��Kİ}�e�r%�bX�fs'�O�j%�`���ND�,K�z?����I���]��GZ#Dh�^�r�9������&s�q;ı,����Kı=�{&���bX���^#��b�W��#��4F��9��ؖ%�`���iȖ%�b{^�Mq;ı,k�v��bX�'~��%��ˮ!v4�c��Dh����ND�,K�{�5��Kİ}�e�r%�`T("r)�ʆ��"o�ߎ'bX�%��K�L�)i�l�W��#��4F�/�|^#��4��@��I�$�}��N	 �}��6#�]�?n���n�p$�����4��K�ǲݢ;֋d���N˛���=Of��F'�mc�b�4F�����28�,K�g2q;ı,�9��Kı/��7��Kı3����F�hò׮�h��4y����h�%���m9ı,K���;ı,ײ�9ı,O�,��֍kR�74�>#��4F/>��h��D���^'bX�%��{.ӑ,K�y����h��1{��e��<k!7.���Kı=���ؖ%�`�^˴�Kı3�̜Nı,K��G#Dh��?m>�ݜ�Li-�޸��bX���ND�,K��d�v%�bX?fsiȖ%�b}��>�GZ#Dh� K��̖�Kn�[�\��WA�J���pS�K)����E��B`�Y�-��v;/5���=C�73vb���y�֫k�����jiyvȯ6Hv:Mҋ���ut�7\;��6pWn+����s�:�f���n(�u��-ͬuح��w��v-�mCb��N|ݸ��d�;�p���͍����������c�7��s1!71-�HmQ��_^p����Xe������1���+��ʑڟ71q��K�(q�/	=�ٴ:+��ͳ����dx�#Dh��ߺqh����3�ӑ,K��_zf���bX�����#��4F�>��%rt�\B�keψ�Dh��Ͼ�ƈ�$O���k�ؖ%�`�^˴�Kĭ��|���F��<������p�팎4F��<�z��GZ#Dh�}�e�r%�bX��s'�,K1y��28�#Dh����e�g�wX��^#��4F/o�L�4F��"w3�8��bX�ٜ6��bX�'���k�ؖ%�bg�۫���Ѳj�Sz��r%�bX���N'bX�%��g�"X�%���d�Nı,K���ƈ�#G���ݕ�ۍ��v�u��7���z��%�\�=sf�ޚ���U�W��[�imra���qh��1y��iȖ%�bg��K��Kİ}�e��ؚ�bX��y��;ı#ߴ����cY	����Dh��>߲^'a�V:�����ND�,K�߲�;ı,�8m9ĭ����W~�Mt����:�,K��]�"X�%��߲�;�P�MA�3�ӑ,K����q;č��~�q�٣�%z�.�h�%��o�x��bX�ٜ6��bX�'u��k�ؖ%�`�^˴�K4F�>���t�\B�knӈ�Dh�,�8m9ı,K߽3|Nı,K��]�"X�%��o�x��bF��� ��d?um��ی�I�5���v��p�F�nR�s�e2�rh
yKz_K�˥�p�팎�F��?_~��֋İ}�e�r%�bX���/�,K��3�ӑ,K��9�{����ɞ��CK��<h��1}~�28�bX�&{~���Kİ~���Kı3_{&���bX�&�,�S���t��Dh���w�N#�%�`���iȖ4Q�C��6n'"s7�f���bX��̻ND�,Dh�I9�z����q�t�:�#K��ND�,K5��\Nı,K��]�"X�%��o�x��bX��ߴ�2k]��!3�h��4Ϸ�Nı,K�!7��ӱ,K�������Kİ~���K7�������/���	�ѧ������g�溉c��h &�ֵ�:���Q7Zi��qh��1{}�dq�4F�&}�e�v%�bX?fp�r%�bF����8��F�����W-�:bW���ƈ�#G�o~�GZ#Dh�~���Kı3��/�,K1{}�dq�4F���O�d�-�F�ƶ�8��F�����h��DϷ�Nı,K��]�"X�%����ӈ�Dh������,)q�.�c#��4F����8��F���^˴�Kı3��/�,KX��p��Dh���_�)���=��&����Kİ}�e�r%�bX�����ؖ%�`���iȖ%�b}|���u�4F��<�R�d�v����/jIr-�-�V;F�2μ�@�Zа�J���%��)�e�]28�#DhϷ�Nı,K��ND�,K5��\Nı,K��]�"X�%��~s�����Ɇ����u�4F���g�"X�%��o�x��bX���ND�,K>߲�;ı,Oe��Mm���L9��ƈ�#G�or�;ı,k�v��bX�&}�e�v%�bX?fp�r%�bX�k'�oÛMn��]��:�#Db����Ȗ%�bg��^'bX�%��g�"X�%��o�x��bX���F���bW���ƈ�#G�o~�GbX�%��g�"X�%��o�x��bX���ND�,K���SN?���Gn����`���c����33R������Vg6Z�f�sS��ڳ��ԯ���d�m�Y��r�sv�w,�6���v�\=��,�m���m���Olz�pF����݈ƺ�v[��R�kr݊�B�nޜ�æ�`�:�W���%v��K�Z��B��<ͧ�/��=�m�;XV��
Ƕ���nzt¶�L͓�Χ#^���\{I����]�Ÿ�w-�c6:#��:��Ҽ�Vi�6S��nb�]ضݧ���4F�����6��bX�&}�e�v%�bX>ײ�?�ؚ�bX����x��bX�'�����,)��.�c#��4F��߲�;ı,OM{.��,K�Ϸ�Nı,K��ND�,Kޞ��Zޚ7u��^#��4F�]�]'"X�%��o�x��bX�ٜ6��bX�&k�f���bX�&M�_�Bò�]*8�#Dh���^'bX�%��g�"X�%���ٮ'bX�%��e�r%�bX��Js��ť�ǭӈ�Dh��Ͼ��Kı3_{5��Kı=5�ND�,K>߲�;ı,Okį୮8�IY���ջNݛ^�>Xޫs٬�tGkn`rp��$kQ3и����u��%�bX�����v%�bX���]'"X�%��߲�;ı,�8m9#Dh�����m�3M�׈�Kı=5�NC�ڐ��*ث�E��֌�&⩀�Obv%���x��bX�{8m9ı#G�Ͼ�GZ#Dh�S�~��rkcį]%ң��4F�>��8��F��`糆ӑ,(CQ55�ߵ��Kı?Mg��Kı;��5KzkX�;�e�N#��4F/���G#K������,K��{.ӑ,K��7�Nı,K髆�oT�)��.�c#��4F�o�}x��F�%��^ˤ�Kı>��/�,K��g�"X�%�߷.f髹�:D�Ʋ�%�(��뭥�<ܘ�#����r��e\a���6d��w����X��~���Iؖ%�b{����v%�bX9���Kı=��5��K#G���_�B6��J�4F�%��o�x���#���`���6��bX�&k߿k�ؖ%�bdײ�h��4y��?�����a���q;ı,�p�r%�bX��ٚ�v%���M��L��]'"X�%h��ߧֈ�#�Mg�K�������r%�bX��ٚ�v%�bX�5�ND�,K�߲�;ı,���#��4F�/��_���ͫ4����ؖ%�bdײ�9ı,O�~���Kİs��iȖ%�bz��׈�Dh���1������vN�6��ǭ�%;��h�u�c�]I������z���qf���+��]*8�#Dh���/�,K��g�"X�%��}��'bX�%��^ˤ�Kı;����Ζ���ŗl���F����8m9ı,Ok��q;ı,ײ�9ı,O�����Kı>��߫t�Bm��ƈ�#G���q;ı,ײ�9��D�O~�~�Nı,K�~��Kı3�Oc�;�F��k�u�4F����]�"X�%��o�x��bX�{8m9İ!�!�j��䜉����ֈ�#D�O���B�Z��iȖ%�b}��^'bX�%����?t�v%�bX��~��'bX�%���L�4F��;}���e6!�n�L׵����=I�Ξͭ��9�g1�{ε��rW�7���5Ď��-Ө�4F�����6��bX�'��f���bX�&M{.���o�7ı3����,K���5��K���i628�#Dh����'a���j%��Y��9ı,O~�~�Nı,K=�6����MD�'޸��I6-�2�mu�:�#Dh�5����,K��7�Nı��MA���m9ı,L׿~��,K�}����&�<J�4�J�4F��"�{�w��v%�bX?���"X�%��}��'bX�䚉�o?]'"X��<����I��]زݧ։İs��iȖ%�a���s?����Kı?��]'"X�%��o�x��bX�$B+��H |��iYYa+l����q�:!�+ ����"Sc��";A�� ��Z0��Q��	YQ�#�;&���� XAt����5�}`��P�D ��*J�"F���z$��(�T��(�$`A���>��oڪl�1�c�z�	� �Чx�t����E��8���E�BW஠K
Ƥ
�Z�!8�۵���{���,X#@�&�t!;~��YK�Ա��M*@~�K�"���//�wlmin���V���Yn]]�.n��e�Ng+��1ب�0�tt�\5D8ʩv�R�n�F�l[V)�����l��!T����ޅ�n��6c WL.��+��v���ؓb�m��d{z�q�Ƕ���2۶�����iZ��^�lɞ
\F�tĔ8��:ޖ���e.$l	 $M����d9��7;M�u��?<���R�3nM+&�B%�sh��[�D�0ڮ�fz�u��WWU&b��Zq'H��0��6Ș�pv��E��W�	;/]i��1�k��������|�r��5�:���ם�v��N6h5��]���.���\\J�,�5�O8-�z��v�M��\��p)�t �kp��s����ltZTqʳ8JƬp[�\�� 9�!�zD�S�"������v	�Hѳ��dwC��s	e�ŗ�ڐ��\�Rs̅�klk�p��v�	����t���Xv7�`�5[Y��P ���V���n���7g\�n������3cfX9m�6XU2���\<��k8M����D�Yڪ�A���Ύ0�Ǥ8�QN5���
;X��q	ⶣ%3H����@E�g�W���Ok�ӷd�vJ�8�}��w�_�D���PV��Dkg�7QX��+0�lq�EY.6�A;;�y
r����^^w�m�ӵ=y�n/4��1����h�ݶӤҴ�d�����)��a���e�hVz����wd8���qwD�)r�����������T�Bz�e�]9�[�����d�=5�Kl�4'^�焞�t���fZ�EJB�.�:˔�-�`*����p5UU�F���l�?+<�Z�M�tX�2�،����m�+ʚu��K�n4pZ��B�`}���#]�g����c����f�i�6��ڛ6P	j�*ݪ���@4p�����ni�
$�6����]
����:sv���y�`���5�9��>�� �TM)D��x�����:-��F��x�[��^�i�C��sZ�G5;]i95i��z���;8�ö��	�clZ�g�)�PZ�;��g�V��j�ye\�g�5:��(;0\
�8�*�9(L�Irh֭�qչޙNͻ����x�6���3�3Pú���彴��l���r��S�ؐ���a��m:T�'!(�N�J��E����jU[�������y!#�J�8���»[�����A�y����p��k:@�]M��\T?qͦ-�q�g�.�c#ƈ�#Ok?����Kı2k�t��bX�&{~���>���%��?p�r%�bV��z}�d�Mt��^#��4H�5�NC�D�K�o?^'bX�%��?p�r%�bX���5��Oɪ��4}c���6e.�Tq�4X�'��~�Nı,K=�6��c����n'����\Nı,K�k���r$h���~�Yݶ�GI�����u�ı,�p�r%�bX���5��Kı2k�t��bX�&{~���H�#�Mg�K\��M&�G$K��}��'bX�%��^ˤ�Kı3��^'bX�%���ND��G��3�
�S!#�����pݹ�ʛh�<�W �`դ"��Z��.]�v+�j�M�׈�Dh���}�Tq�4X�&{~���Kİs��iȖ%h�_>��h��4}��wMlx�9M%ң��4F����8��ί�D�K;�6��bX�'���\Nı,K&��Iȟ���'ْ~)�e��;�m�N#��4F/�~��Kı3_fk�ؖ%�bdײ�9ı,L����ؖ%�b}0�����6y��28�#Dh����'bX�%��^ˤ�Kı3��^'bX��Fj���iȖ%�>�{��k$�h;�4��h����{.ӑ,K��o�x��bX�{8m9ı,L�ٚ�v%�bX����pn9L=q���ڔw9�;l�W��X]���:w���^܌g����ۛ�M�wiȖ%�b}��^'bX�%���ND�,K��3\�>���$b�~�28�#Dh��П�����1%�ַx��bX�{8m9ı,Ok��q;ı,L��]'"X�%h���ӈ�G������Y��k&4�&�c#��4F���߯ֈ�"X�5�ND��u�D�L����ؖ%�`�g�"X�%�s�{0�ŻVRk.�:�#Dh��~��bX�&{~���Kİs��iȖ%��&}���BE3��kf�ݱ�\�4�J!���<�#�Ci��L�bX�&}��'bX�%��^�*8�#Dh�����l�v%ƛ3��n��"6	Ŏ<cvn�[���:#��1##7M&)��cg.ƶ�8��F����8m9ı,L�3�Nı,K&��IȖ%�bg��Nı,K�k���٦���28�#Dh�ϳ�N����j%��k?]'"X�%����׉ؖ%�`糆ӑ?)���b?|?�?ٻ4ҹ����Dh����~�ND�,K�߲�;���Q5�~��Kı3߿w�ؖ%�`������c{��]*8�#�Q=����;ı,���ӑ,K��ٝ�v%�`y�	�� )B $Qa#ń��~T�"~��ۤ�Kč~��u�9&�[�ֈ�,�p�r%�bX~9�~��'�,K��5����,K��7�Nı�7����>HŜ�[����.��k�a�og�7Q�ae��M�����c���f�p��ldu�4F�������u�D�,L��]'"X�%��o�x��5İg�ND�,K�韷%��v���]x��F��>wߥG�/�]��K?����;ı,����ND�,K��3\N�����b~�ܓX�kcƹ�i.�h��4{�}�q;ı,��m9ı,Ok��q;ı,L��]'"X�%��z�)�e�ƗSKv�GZ#Dh�_{�y9ı,Ok��q;ı,ײ�9ı,O�~���Kı>�.���Y^�gK��dq�4F��>�߷�,K��f]�"X�%��o�x��bX�k2�9ı,N�ޙ�L�In���i���S��l�����9L��;훾���ԷQ���� \n�s��m�N����c�汅�vHZd�U�4Rs����]uB�n	����d�7n ��b,��R�uzݖm��Q�V᱂�r�n�2
���L��͸^�3��\���n�l�8\�	H۝���]IGьr,��b۳��1�.��F�l��i�%�RH˴���v77=���z�m0jێ�i��<��y�W���^���ni�s;��u4F��?;����E�bX�����ؖ%�`�.�������KĿ�����Kİ}~�����2�]t��Dh���7�N�� GQ5���߮ӑ,KĿ�����Kı2k2�9ı#G�{'Ӻ룒��-ӈ�Dh�f�m9ı,Ok=��v%�bX�5�t��bX�'�~���KČ^�#7����t��l�8�#D��g�\Nı,K&�.��,K��o�x��bX�f�m9ı,G��{�n\k�e&���u�4F�ѓY�IȖ%�b}��^'bX�%����ND�,K��f���bX�'�o��l��v]�����SѶ�o���Y��nɌ��#U��<'�譛�C��a7n�t��bX�'�~���Kİs7�iȖ%�b{Y���,K��߾�h��4w�d���1�.��'bX�%����NCH�GQ5������,K�ɬˤ�Kı>��/�?
!���b{��w_���M6-{K�G#Dh���~�Nı,K&�.��,K����^'bX�%����ND�,K=�xk�d�M+�ݮۈ�Dh��
�O߶��,K������v%�bX9�ɴ�Kı/��o�ؖ%�`����Z��v\�ڣ��4F����q�bX�����6��bX�%�g��;ı,K�3zND�,K3�}�)ۋ��;[z�!s�8ռ\��fAs�6z��5����6�
��*li���,K���M�"X�%���f���bX�&Mf]'"X�%���}8��F����G�����)	��m9ı,L�{5��?$uQ,O�_�]'"X�%������v%�bX9���q�4F���~?oÛ�YI�����Kı2k2�9ı,L����ؖ=@7�Ț���M�"X�%��}��'bX�%����[&�tt�]*8�#Dh���ӈ�DsLQ�#@��+�q4�7Z�UW�n6��5�G"�:�M�mzWj�/>�@���%! &C"Ĥ]<O�r;4�7=�U��Gd�<iS"��
yKrLy#�$$����~�@��Z/z������@��1��4D�����Z�&�U�ހ��h��5�>�c񹀓�z]~z[)��Y�r���Z����En=���׬�9[^�fy��o��x��ߤy���b��I �z��������S@��w�����>����2�a�c�Gjx�;��������m�.�I2��ݢ�d�Η#v��r~���h����S@/�f�ws��DO��8'�W�^���h���9[^��$u��5%<R�'#�/�O� ��h��@��^��ޯVH��Rcd��@=�f����^���S@��c��b��I4Vנr�נu������� K�I��Cߤ���6e��J�,�(�v67�����ݓl/���3X���۱Ħ6Q� Y�7Jn��%��y�֥�5�.����-mk�z�lp��3�f��fsv�]ly��1ͽ�=��xt��4�Q����g �X
���8�4�X��q�3[�:��Ӯ9���6���J��s��iV47s�RK�H=+���nj X�|����}�����闏.���e�e��G9��-��]�5��v���V���&ng`,��K���~V���S@=�f����}:�n6����(�q�l��{z��3? ��z]��@���dy1�����f����
���l�����pND�<LNM���{k�-��{����tI�H��q�{k�-��{��*��������������D�d��;%���8z��.��l=:|p8�9NjK�����f8���}����f�U��{k�=���D�dN�' ��j<Ȓf&f�"(T��W�^��b4�SX��iD�M���{k�:�M ��h�1QA�Ә4�F��*�נu��}�4Vנw���F��(�q�l��_z����{���p]SoLx<&D��n���zՇ���kV����ۃX�O3��$kPE�̏&<x����u����@U�+���DD~�M�4G
�U���a�6��=�j�*���=�)�U�W�ˁ�PO$h�=�z��f�rp��v�	(JH�ZH5m!��&�����]���8E;�$����!�H+���&��X��B�@B
T ��%I ��LX���$`�,���"�ZZѬRkC�� ��FD�$�<u��!"HH"E����X�$�"�B��*�J���!# ��jt<
�N
z�B��^ E�
AT4�EC� <UM�=�*⫀��(b�$��-��a�5F�`Fc����)�u}V�궽���������7d��@����ֽ����.�O��b�豩�f5��A���Fj�ջCq=���+8zNe�"���sǑ��CQ�qŠz�נr�^��YM����ǋ��
�޹$��k�~�������������?o?^=������^=��F Q�����^֒�h<�ֵ�pA�lll}���pA�llls������ ؃�DAPA�����{�����=���b���r���������u����k�~�����ٿ߯����5�?k�`�`�`�D�����������I���M�d&�k��(�
1�A�o����A�A�A�A�~����� � � � �?~���A�A�A�A���ׂ`�`��@�/߾�?;�����G3ܹG<F�Srj�/gv	�F^�Z�V.H��H��M%6v[�ӂ� Q�b`�������A�A�A�A�~�ӂ`�`�`�`���������ٿ߯���F ^|�߇;d��X].ׂ`�`�`�`���������?g?N=�������k�`�`�`�`�������A�A�A�A����v�Zkt��68 ]b�F l{y��A�lll}���\{��~��������N=���F _�{�O��L�+֖l� �66/�Q5����pA�lllk���� �666>�ߺpA�llls�s���� � � � ��r�~ԅsf���u��u�b�`�������A�A�A�C��������A�A�A�A����ӂ`�`�`�`��g����� � � � �0".��y�%����Y1�嬍��]+·f���Ųf����X�LgQ:�)	�����8t!
�[n1�0�.z�]�)�v�P�f�N	���n��ƣƖ4��{\���IP[��pi�.�$זW���s������}\��]�t��h�Y�����.���|_$��D�RD��Z9�<UQ�������,��s6%Ⅹ�i%�m�m���$V�����[X�u��Ht!��m��u2\Z�l�b-ێ;j໲f�b���;Z���w� �`�`�`�����{���8 �6667?~��=����k�~�����3����{��1+sMq��(�
1�@������A�A�A�A�����A�llls_��� �666?�~�ӂ`�`�`�F _V��_��4��Bk6|.��������� �666>����=�����߿t��� � � � ���� �666?�f?Y�)��ҭ6�.��@�(���?k�`�`�`�`�����8 �6669���\{������'�&~'4i6�8&���z�}����zm�@�z��-�7#D$18��-��T�3{��+WSY�j��n�
⡮��C�m�)3@�z� �٠r�^�m����<����&F�G�Z�nG��LLՂ������:�+�;��
�1�B$�@�mz��h��@-�h�W6I �5���b��@9[^�ws�z�����$jcɉ�$s4�ՠ�4Vנ[e4��/��LR?�q����l��<lیh���˻7�ƭ˻Zan5]HNܘ6��G�$������r���)�uv���Ǖ<����@�mz�S@�ֽ �٠~��kG��d�7�&��-��.��*M� l��ꂆ�I��� ~]���Ζ�NF�$hq8h������z��)�^m")��2G�[l�9^�@��h�W�L��.��� S	(���;����Ep��b��,�Y�X9�5���R,B������z��)�u�O~�o4bq�yyp^a�wyzK�r�U�	%�?P*iހ�ʹ�#b��"I���f���z�S@��xF"d���	"����r�%���"&b,������������������]�%�e$�9^�@��h_U��4�;��ࡶJ�D�o���5m�mgv��;C�`��LH�b��<&�І����M���g��__���g�lx�NF��D8�ZW�o��}��*���]�@�>hU��S"c�- �٠r�^�k����;��U<X�!�d�rh�������Z.�h9�����ٹ�yp\0�M��l��ץ4�f���5�&�v�@@�҇���H�w�(C���cd� ���5���ҷ6W)̘#�؎��2�D�ی��=,�-]Q��9�%9J�a�X�{4F�r�F�����8bT�s�R��πv}��%	u��Ջ�	D�WO����;[Mg�1���hvz6'>�.^nv�z�l-�t:�d�2A���b�Ӓ�h0��<:�V�Z�ɳ]��ݕݡ�v�W���.͛�6�i[b���6&�:��0�vwGnM�bY�v�œ������r6Lq��$������m�+���M�{��"d���!�	%��11>��ן�@����b7���<�$O�bmdRM���@������f���qjH�9e^e�9�m�Ѡ'iր$�h}������{>�c�"q�8��L�:�+����r�%��=�����W�4��ۮ�qB��l��uΏX{�e�"s8�g+/����P�� �t;2�� ����:�+�X���;_-��'�Ĥ1���M�����D�DD]��i�|��hIf����w��>�H����iǠ}���@���@-�h����Y�2c�l(��4L��5������A����ߍ�~�)��$x�A�hIf��|�����>]����V~!�\+�h˩K<s�nݏ��]n�;&1縛��Ѳp�9�;���u�:]�I�
�m��=�)��4֫��Y&@S	#�-���$w?�Z �y�}_%zꏺ7+3�/�˫ʼ4�n�$�M���$�LzI����ڭn���4���UuYU�veXfehz*�o4�n��#C�1�.���@�w�x�
L2)��=^��l���ՠUmz�Um�+۰��R<��7p�&=v�<#��v�x���R�3w����K#�v����������V�[l�}�h�yȡ�yvff�ZU��L]��{נ	{�h�M�{ΉL�)#ŉȜZ����%�8���3@��@�WU(̬�3˳
̽]����rI��̼�j?`�� <�3��$�f\�2d
b2I&�m��?��<̲�����ՠ}_%z���YYq��3�ܲ�wc�vy�n��4�U��J�w<F�\�2�<Y$rA�85#n'��@�ҭ��+s?�x��(V:,�2*/̭+J����Q��ހ��h��[��y�$[T��O1I������%���33U�mրݷZ�����]f��a�4�����@"~����ۭ+J�=3]|��	:�dP����E�{�h[^���3\�fk2�I��}$BH�@$(�ˠM2#%|`V��HH������R�(�`Ji
IP�&��C!B<H���/δ��Q�%֎A[	�6��ki�G�D�4h������F�P`�qJ!��ۭMV���頑 BF2�	��	��7@��`B,@��B�x	�c�4�i�{k!!��T�mx�0` �"	"&���$�}�w�m���mW�NJ�ʫA�5��Div��Vt�a;4`ɇ���ꋞ�N��pҫ�VL�HR�c�b�X���)�:ɶ��D���n�n���@��V��.�
v��NƸ.$ �����l;<�����k:��� ��Z��h,��\k֚��Ya��K��i�3�][�������ej�j���V��e[���.��!:����O���a�n�Wi�F4�m�'��3���j3�������WUV�:[��;%��dC�R���4jr.x��G)��`ۍY��یqӹu�����㱚\ji��ĳ��e�63Y��&�sa"чlk�V �荌g#ݰ��8c�'6)r��d)G�8iv��L��y�ۮ{As�l+WR���`-�od\�c2�d�ݶ어�QQ0p��ζ4�6��6�6������sɭK����%<g����!��O\�E��l*�4�����w;N�Onyv���n{V�9뙐��3�c�^�;��K=�r�vQ�K�m�[3��t
��<g�����vi��gH�X�!`��1�%7#<�k!������l���1R��5eyg;�mFѭ�n�m�g����.q�)z����&��Z�ݳ�8�I��G0p���Wd�\[\#He�m[���^��vz�ҙ2�b�7b���۴�'k�q[A�]I�E͹��$X0Y�a�1ʩvlc�q��������h�Z�ۥ��mn5sRem�3��ut�bp���+���t���	�U�t�n˻U�h֭�o�@�l�x*�����jhs(lJ�K�uZ���ך�q�*�U\Q�3Ӻ����gEn2���y)y5�j@�#a��,7mh*-�n�`Ͷl�*�V�Us��-"10T9NRm�!���}������K%����G.�8��75��-�m�9fv��4>[!�Ad�f�6��b�5���`�*��mFH�=PVx�usr���pT���C�DP�G��������u�i,���ͱ�P�F�2rqA���+�Vރ�,�-��[��t��naqx�7��lh\�l��u������D&�%�hШ����m���@�ָ	�{�	�hG�cq{q۞i��l.9�c9����V� Ǘd�|k6�{<���u\皺{p���Q��ٱ�#�t��kn|�ʐ�����L�b[�3�S��2��`m���Уj��1���r]pH�6�\�4��N�)�L�)8��~�����&4�mHK��z��}��}_%zV�8���A�mրC�_�"l��H�W���)�{�h[^�����W؃pɐ�����x��*�$�@��J��e˱�1�I�Hۉ�C����>�h&��W�^���m�4�V:2�+12&E�Umz���)�{�h���덠lN����rb�6�\ڷ5!�w1]���g���'��v x����S#q���4l���ՠUmzR�\ID�&M���-���i1+&"bI��{�W������+7�"ߗ���2(�2I����$�OU���{�_uB�#*�2<X��ŠUmz���)�{�h�䉲Hdl�I�z����M�]�@-�h���E<�)�.�x����l�VN����z�y�p�2r4L���d"Ħ$�@��h�iV�$�z"c�X*^�����³"�����̫�@��J��@�y�usw�[e4Y�u�E12&E#������f��z-�H��,3�fxնi�r�@��1X�ř�]�h9��^����Ɓ�|�����c�$��M4��-����^�[l�=^��W�.��ͮ{u֐��#>�*������Y�@mmǴ'����G%�Q�u:'�uV�������|m�@�{k�-���Գ�<�RI��8��f�����-�������<�ă��Y_�l�"�h�w�$�8���^��@=�{4�T��PL�X���q��M�mz���I?��D�!\[7��k�O|g�'!28��'�mzm�@�ֽ�)�}��������MG��r��]���$2�N��] ���>�[�į�PB�$�	��<�G������9u�@��h�k�;�LN���I���3@��}3����x�蚥^��@>�女}*�Đ���"i��m��>���隡��@T���T�*22(��$��=Vנ�4]k�q1M�f�}�Jaq�VfdTU]^^�$�h\��	,F��$�@ɕ3���O�N�Y!��a����;	.���z��ݧ��&�T�)�S)��V��.f�Yx�����.�tͣ�>�a���$5�GpmƼ(s=��4��l%�KnDOgɝ۬��b�ٺ뇝��9��c�zW�&��۞6̖Q60��'.�gu�^�ح�\R���nb�l�Y�v2��i�@�nodtN{\�c�
�[׳*���zm��["d�1	~^^s���a���:����n3�Z[�c����B=v�ܽ���2��c#p���.�����I��X��I_�31?X���G��A2bSǠ[e7�31#��;�������D��Q�E�qeaY���H�4_}��m�w�$u�m��94ŏHm�y��%m�@�_�z�S@�[^���bu*�� ���/3@��@s13��~��|��f��*9D���f.�C��U��8��k�m۶	9��Ӝn�������7�`D�R=�)�z��@��~���D��}`��נ7�˨�e�fU��,D������<�<�k�?.��o��>~@�������M�bir�M��:�+�X��I^� ~�_�e�l�n�k�� D�����oﾟ���
��@�Ө���YU�ee��	,F��&f'���t۽�Z�
�ꯊH8b�4�G�lQr�Խ��Bn�ī�����h��+���+�X��!�8h�k�*���Z��Ɉ���f���V\eYvff^��%zW%zK�}I+�L�L��&ff�i�E��(��#+#2��O޽�)���<��Vנz��@�p�j�����������s��hM��Umz��*��=�~Z�L�$�.(��4�%z�&a�n� �7z�S@�=�T�H�73��P�m��H��Z�d�6陇�������ƭ[��
��8q	,�tv�#�bĢq����=�Z�l��g������k�4�&B7��\���J�.Ǐ�u6�@T��q鈙���+���2���{����
��@�ֽ���\�Y�Y��fU��f&��w�:mށ���rN���� ��o�M��QJ(��&�L�G�Umz���V���6�Ԓ�"�\U�)�!w9un���!��&��}���W5�W�'<Q�1ᄘdRɠr�^���hRJ�������@�ç[U0�a�4ԏ@��h�k�m�������DO�&bb���[u���w�ff�{נ	%�z*�&�@�oύ�����=v�$�����LU6�h
�w�$����mހ3-x}�M�d#dRM �hy�y��31>��x�^��@K4LL�~&"=���*E����3�[�Mq��z��I���uv���k\֚���;vЈ�6�n��5�Jm�|��;��n��[�c	�`�a	��St[�v4X��ҝb�ꮜ�\\�sg�/J��]�Cu�ɛ�Xd��l��p��m�v9��R����&'��]�Ր�$�O0�{%;\��*�I�az�{��R��I,V�K�6���zP��k���d���{b#.���;�[��y���iq���lq3rS�L�D,��)�q��Қ���$��3?�&�@��պ����Ȫ�.�2� �%�興���Rn��#}311T:�uu]U�e^Vff�6�h\��	,F�}�f��_rX��$�"��M�ֽ�j��,�q31M���e�2(˃ ȚiǠZ�� ��� ���=]���B��1�Lۏ �pU̻^7=gKSǯK����āsV!�{�����䶜s#�dn/�z��= ���=]����@=�\aq�D�Lx�n= �پp~`���O�"�sW��mց��+�DLMP2��E�e�]�Y����%���311U�&�@o4��PmeEVHfff���h���RJ�=>��������\��cO#RLJA�"p�?.�����m��RN��#@s̡��[U7�'��m׹9�Aq/n1Iui�;��ޘ�U�cږ���w{ɳ���v�us����{޽��W�$���@�cٷ�6����߯?���@���ƀs��@K4ˠřYe��7uuu�rI����'o�5����GÆ�HB0���i��6��ͬ�-]��J�p�Z�WT)*HA�2��m"I$@�,5BiIZ`�#�����↴kH��!
�Q�Bс$F0
�&� j�P�3-a$$f�(���@ J7�|�M�#�|����.	D�#��E}�J
>E̞�6h������q��xc$���G�&"o��נ����ܯ@Ib4�E�DG$ŉF��m��y�1��_�{����@����-ees����M������9��ZzvLc��
�7]nF���Od\�����9^���h�K����o4��dħ�RG�[e4�[4�f���~�<�=��퉸�$"NF�4���@-�h��h�MP.%U�e]Y��y���b"���@����I33y9"�҄AE�����;���\x`�Rɠz�����@?rY�	%��"g��חtX����m�J{[��ύ:ܼhcDL&N�B���uŴM6��!;G���z���.�6�������l�m�����uY�3./#/.�/2��%��&j���@�o�@�ڴ}P�"H��Lmɠ	%��ܯG33M�u�}I��
g��\l�"�hy�y�x������@�\��z"""���@\&mP�L�X���H�_U�y��|� 6�hWr��JC������3ʌ��磞�"��.���c*��j�X�[���lF�n������ɧnƎGk�-pd4�����Q�"gvq�n���d���=�\�ptM��\{lq����ջ������ծ×�N�=���+g[�6�=���Xyp��2u�=q�u¤7V��gkn:5��讔�cZ��L����pݫ���/.7F�"���m*g�+k/O.Nٝs�t݉���'si9���;Zl���=����??	�b���+�:��z �,�>��~�@ݧZX}O>QM26dr= ���=]��	_*�?W%z�&&c�3v6[.(�<0sGrh}���-}V��������_�����Bɐ�iǡ鉉���:�>���\�@�������jdx�G��Z�ֽ�?�<�������M���*�?.�řV]�vv|�l�`�����ۺ���#�H�$�⸴Z*r�Vx����~~~~_`�wW�Z�Z�ֽ �����dٚ׵ۍ�'��y�xi�$1�1������z �,���aHY2bS��@��Z�ֽ>��33�H����9[��;�שƙ�m8�˭zz٠z�����3<�1}g�-����L"i���4��@�rO? շZ��� ��*�Ue�u�]r��\u��,5j5��q�`Ɠ���+v'��MI����R
I��Y�.��@?rY蘈���M��YU1�Y2m94�ՠ~]k��� ������3<H���5���dQጎE�z��= �٤H�����Z7��{�ŻI���j�׍�@�'�߿m �h	ZU�陉��7z �\\[�&�!��)&�{�f�k�h�[z �Y�9����uL������˻��#�+6�㮫GT�g���b�Q���k5d�;����n�!,��)�RG�����h�Z��f���@��ש��"y��^V���+�1T*mށԓ������$H�F�?��&�[5��N6*mށ�ܯOD�Rv�hͼ�;��T�A�)�#q��]��]�@����N�Q�A �`@X�E��"��]g߻�rI��j~-��6U���h�*�=3_6��
�w��f��թ��G�0�)�"26�[B�,c��Xe6:�՝}_���X��,��9Q��NU�~ ���RJ���L�D�}`�����*���1��H�)�rh��@r���Z�ҭ�2�&n���xō��� >��{ψ~}�@�w|��KH�	L�X���I�uuV����@�I^�����������j8D�q���/�ՠr�� ��h]�@����<�ĲԢj&`�2̈pOM���=��|: �!�81��Uv܆��w%qls��5㤞T9��T�g�ִ�nv�m�����nc,�A�p@��nkOl�:�E�q�p�=�"�٭6��v2�y($��g#^/M��EF#gf�����3�<�n��QlGR�a綄a�yşd��j��%�6�sPY�`|2����7kD���1������k+�Í�ĸ��3ny����ua�W���s<��R*��H���|�
���:�V�}v���K#ǀ������*�@�iV����@�I^����>N���PT\`eU����	�u�/�*��1T����~���y�dY&G�š�LǦ&&���ƀ��נ�f��ҭ �=�271��ŉHh��@/u�Wj�/�S@��/�q`�&&�c�� �Y�J�u�vF:|y��r�a-��]�#+7��g��bDFı�HA�#�����Wj�/�S@�mz����	��IF��q����1�� _�9�~~Z��z{��=�mZ�F8���m8��h��@/u�Wj�-b\�i�#M��$�C��3�<O��^�y�f��ҭ�iv-���^��Qa��yw��*�W�z&&}/������-�����U��j3�i��*�<��gv.3b�wM��㎍��]�3tƜ��X�I���Wj�/�ՠr�� ��h�U湑d�`2^eh
�J���LU
�w�:Iށ��Z�{�dNcr9�ɠr��/�����0# ��1J*�b�EI�"~O�A�=�w��I����@)�����z]��]�@��^����}:�j!�W���+J�LLD�&b"=�޿��= ��h�:��51,1��y�n*D�z��������U�-���W]`��ܒ1�8)#n-�mzz٠�c�����[u�7B�wV^eU�]ڊG���{��/;V�}v�������ߟ���lٷ��m��$�=�ڪ�]�W��阙���v���UU4�~��^��f8,<��i�2jI.�i��ۚ�f��m�ٙ��ۊ
�U~C�$�������O�}���k3mڤ���%[��I$��?~I"۹5$�[���$�θjI���Pר�ؔ$KOV�mmָ�l����65j�N�-�'P��J:3���(��I+��OߒH��MI%�j=33}uT�ۻڪ������Pl����I�����I+�����IV�oRI.��߿��3�3�ڴ�`j!$�$�&���}��$�n��$��~��U[��$������pRdo>�I� Ao�����I>�����'��^I?��E����Ͻ�O߫�_����ˤ����I%�l��$��q�I/m�~��W5��r�nϑp)-�"�:>�o<4/"�����Ց�JA�diR�E����-Jh��m t�J�1��d7OO#g~OW@"R ���jh40����@7���m�$����"[��떲�U�n�N����6��ԕ :y��i�2u�qs)+R�
��ܹ%쵰f�g͎���v���<�0qK��
\��ݺ�f��^Ç���G�I�kd�٥nͲ�	���F	���� u��.۶{^E{e�btbj�Qc$�ٶ�C<u2�*�v�m���l�:2�)k$�a��LK���� l����q�vj�k������\����O�t��^�TcY�,ƦI�u�i6��]�.�ո����K
���a����K��i��9�}g0�7&<4nۍ"0�����$�I%�9�z��3>{/*`��D�q��h�J�ۘ*^#RL9s�:M�|���1����csM��L�c�+��yl�yk.eņ�W�/H�q�,���m*�@S��!�t2�>�n��(�N��|
Y���B3��vx6bx��q���ܝ�n���DƹYK�G�����Q�a펤y��;Fq�̱�]��vwl�{bQ��N��֦ҒNv��c�}�z�Ƈ1�v�e�3��m)��{9(t�xd�n�;����qWnGn�&�kL�I��q�����R�IVK �q���؊6CcT�t=��C���5h'�t�B�ZZH�vH�B�[�v'�� ƁY]�f��f���1�`S�L�eq��]�m�;;lQ\��&�:n���Q�����C`�x���z��D-<���5ʵ���l7[�Y�^�Is���<��O8㮺g��;l�*��;��$�u� ����*��5ں�S"�9:-�D�5\�BF��{nRZ�WU��b� �ó�7Q���UUpR��9�b��5Q�^MM��r���U��6]e�u��՞�C6ٲ�Z��-<�e�ZNjR�.3�Ѐ�uӲ��N���Y��M�q��牝�QZ����*�����g��!V�Bt[V�m�Y%U�+�L8q�۝�*�����	�ُ�驉�@I\8d.%�P�&t�<�TL<�/�$��O'�ke�����y�k�n�kW=��a��ʶD��j����γ\p��a�]�����*��ylc �WmOo,A�mm�-��[{h6�.�1�.�".����bkO�𵱧��mHn&{m����ז��Kш��c�,oLk��E	ּ.��P� 8RwO !��@��������L<عis�5��������[��{���#�)��kKm�ԗI����V��γ������ç�����𛮻S_@���\�۞�e�m�5��k�U�@�{�/￿���%�<��x�!��ǩ$�KW��%[��I$�[?~I*��{�fg�cm/z���Lr5 ������oRI+��ߒJ�w���-_�$��>��'#s,Q��$��l��$��r����bU��U8���y���UUSR�5��E�ܛ�$��Y�$�KW��%S�=I$�[?~I/SK�A<����UɃE�4廜�Mv�D\�r{t�\n�s��[R}�y���[L&B$�I�$��}���$��=I$�[?��<�=���_}��$�ο#��Rc�6���$�vǸq5�[sٛ�m���\�۞�e���T���~���O�����~��U[��$��j��$����$��j�G��$0�D���$�V�=I%zZ�~��V�]mU8���i��9�]E���̆5�4�h��@��zz٠^�s@�����0	00cQc���\�`����Aq�m>:F���I���V!��{�/�����ˬ �/2������f��-�O�W��@��0�&��cŊ8�rY�$�ƀ�ҭRJ��@�T��x܉��nM�>4�դ��� �B��T��� �1!$����^�%�4�d
��LdIL�4�ՠ~Vנ���g�b��Ɓx�3�1���F�Z�mzz٠wt��yڴއ��Ga޺�lYN��;q�[A۔i.�Q����5�lS��bZ�<Nsk�*~ �l�;�S@��Z�mzb���x4@�"�I4��/;V��u�@/[4��l��d2&4�4֕h������P�y�rX���u8a9x#�h�Z���@����阙ɉ��ܭ_�@\�D�s$�cł�h�f��t��yڴ��Z������LNL��~Mq��%�\��:�=Y�Nݸx�6.���6�k&4��D�nM��M�h�ڴ��@�K�
�a�%0p�ZU�"��[u�7��؍s>y���K6s�9qh���@%�8����䱚V�h�Q��ڊ!��nE����Қ�j��3��|����i`�	JI�{�)�^v��;V�^�h3�3$�G~��6�W��M6�̍����]a\�^vV�:��Q���p�Sv�3��ϐ�����/m�m��w��\8��m:�g���\�zyu�<'Oʽ$␗���I��;n��hƳ<�qT�#���q�s�<��K��,s��I�f]s��Py�&����RЌ�=su��U�:M����x(�K�.x#0����v�b�BvWjb�b��s0������lmyS�Y`�6�u��1f�u^]�YQR�z�V�q̻��o������4��Zz٠{�)�~���#�#� dr-�;V�^�h�Jh��@���Lm�I<PmǠ���Қ�j�?.���e��� �7#�@��S@����;V�_m�ފ�T�̈SƜ4Ϫ�=1,n� >o4���8U>zrt��vXQ۞�eȴ滚�Qì����������GMg���7/WR�������h�٠{zS@����<J�d�Gu�۴�m���nA#̗��P��6���/>�@�]�@���m h�0�AI4oJh�U�r�נ�f������CA1%!�^}V�~�� ��4��?{�א$�� Dn- ����@��4Ϫ�ފ�Ӎ�2I���	��cmHxn�մ�;d7M�v�����=1�\�d̐h�q��194�l�-�M��޳@(w%A�!$F�rh���yڴ޳@/[4�K�4�c"��h�f�&y��������Y^��������[&'�9��N+��u�@�Қ�)�~��*����m�"�*�^�ץ4�S@�����u�n3&4���h�[6�nj8�]�6w=< ����^�SV��#�L�G�u�M���:��@���޳��1d~�bJC@��obE]T�k�;���33�1#�uH؇�PHh|��@�ڴ�)�[e4h�d�FG4@n-�j�:���m������`� ��X�$P�y�瑹*������ �$�@�؍%��9_*���@r�A���m�6��sn�IT�q˫G4�2g���a��rHZ7 j��Bs�:1y�o�r�U�*I^�˱K6s9 �p�:��@����)�[e4�]�S����@����)�[e4W��;ӦXŃD"�$q�zS@��hK��S���t*�yraV]Va�[e4W��*�^�ץ4�������H�ͥa5Slx�8�v�d�I�\��8f�
'�j98ƞi6:��$��Y���ն�����*q�4���)�8{M��۠y�[�����k��tm�>n�i��x�O��8�J�ų�om����'m�YX̚�Q���$����g!���{z�;	R3a4ߤ�{K>I:���S���h�slf�p����Q�+ϻ��{���ܙ��烧jCI�@A��q���b�ű�jiz�.��9��#�D�Lq�E�Hz����*�@�؏��@��h�n�ȫ�#� ӏ@��z^��/YM�����5pq̎A�z^��,F�򈙉�DE���V��~���.FV�<��<i�@�e4���*�^�ץ4ݝZY�x㘱ɑ��4WʴLLO�=�޿�~y�@\�4�mR(�H(�c�xƼ���$A��.�`;'=��;k�s̽�Ń�C2'#�;!k�qȴ
��@�Қ�S@����:e��B,!!�^��fxdL�ٙ�Qg>7?=�;N�$����H���2�	i�һ&ύ�ߛ��9_*��MP�y�&����Q[Yf]�a�f^F��"���@o4�)�[n��T9��G4@n- �٠u�M�w4���:��?1l�����
^��m��	�k��#�� �e��ku���6X?{���%�f���8����Y�[n���Zm�@/�r2����B�4�[n���zm�@�қ�f${�~̈́�£2�#@TӽRJ�����L��}� ~��!!!@�&�8��|@����څ��!�Z�HߒR�P���>~bC�����()))������j1H h�������ob1zq���Z��XAې4la�!�1��#�d-e)i�#���~��S�Y"�I>j�@v��`@}�>%,+Z�B������!i*F,��Ȅ�"ƃ0t���w�
��ba#U��[������}�>!P��q�&����!�
�k��@F+�l���"��#Āf q(YxKޞH8V�XR"IO�Q���6�T� #hN��J0�J�'a	MG�!�5dV]Ɉ���X	���G�@4�(�#���MJo�Ɔ����L�<��p�B9�� �� HZ�JJ[[HҶR�E����)���M#�*F)�1J)��(B)�(�"*B�V�R�>�Έ Q��i �(:AzȧPE�AD<?(�y���NI=���G��ˢ��ȫʻ����6�@�؍$�4?�i[N�ʲIqQ5�&H��:���m��+��If�鈘�̧N��Ȭ'+2�s*�7C��칣/l��&�^8$Ύ���^�j���fu�y��2�0�m�hK��Ic�L�`��Ɓ�����3/ ��
3/#@�z� �٠u�M�w4xv��� ӏ@-�hzSO�����*����sj����D�hz&bf"�Z���4����f"&L��� �U�C���2�ɺ�4����%矯�{���b4^����qEH�t�ٮ��b�Cg��^�&z�ōl7�6XD�t��뙶9�Jf���zm�@�Қ��h���q�J"m�#�m��$_���oc@�|�}5B�X̚��0���94����h_U�Umz�yO�d�FҐ�-�s@����k�:������F�I2ALH�h_U�Umz^��-�s@��bE@%Z(A[AA @�E�*��wMe�����Y�	�:+;"��ўw�ml�ϖ8[���v��v���S�"ڹ<껕�wb��y��F�d�m�=�68��OS��O�h�Mη=�n��֭v�Λ{S5����ڐ�yݕ��#bM��Z������uXzW��g��51�򕚭��r[��m��CW�I{l�h��qt���lqc��ƣ��kl�j�4�m&긻@+��ۋ��iwa��%�dݣ�Z�I�uk���3C��#;a��vm	X�`.� �z.�h	%��%|�@.w6�I�A�dR)�oJh۹�Z���k���ŕ5�"��w4_U�Umz�)�~�:�cܘ〱�Rf�k�
��@��4m��?Q��Y#B�9�@���zS@�����ho��?�ǋ�`���4*U=���+a��6P-̡��j�ǢT�5��dk^��6�oJh۹�Z���k�?{T��!����6|m���p�BK	�/<�\�@��^�oJh���q��0#��Z���k��3�<�<I���oc@>⒋ʸ���Ⱥ2�ZVנ[Қ��h��@.w1�I�GY�G�[Қ��h��@����⮦��6��	�ܦ�:K#:��vs��6�:��]��z}��R!�FdD�Jx���z����hrV�""?P6���	�Q{��Qy�e�F���q13C����f�����<ď~k�)�,��D܎E�}u���3��Ȃt#���Oʜ����4�w�{�^�y�YLqš�6��M�h��h�*�?Wu�RK��0���4��h_U�^vց˱���P�3��de�#��O�to(Y�в=�cn�z�R^'��WU��YDjj$�� �s?~w�[e4�)�[n�{��8�8�� 7���k���5��oc@�|�\�P}�����qő7Z�ύ�v4uI�u�7mր/��)YE�UVM���b&&)��F���z+J�(�.���	'��Ђ�A�I�B9~��>6���;h�b뜎�������ՠu�M���7��?��܌�-���u�x���!���jOO�x֎wS�k�-Q�#k�sdЪ�=��hzS@�n���z���Ǒ<qE�d�I4�)�u�s@�z� �l�?.�V�x��	K0�9%��u.W������=�{4�?���V�G1�L8�h_U�	%�.�hzf)��F�r)2��3"�������К�~��4���=�&.	T�r8�'M����cmւrܘ��etх��t= ��vr��!�6��|m���\�u���
m�m��΍Ħ��]p�R�;o�IS����KG]��O����A� vl��[�Os�r����!��!�4˻�$�5�OiԹ�krh�͜�11��ū:�Zk��R����`��s�tj�����]Y��6�{{��g:�أCK��mv�nݸY��9޳-Վ�=�K��q�s�v#�f�3���	�f��[+�Z �Y����*̈q$��8h۹�u}V�[l�:������xn<q�br693@��� �٠u�M�w4իX�	cɏ"m�"�m�^��-�sC�_��h��Bcb�,�$�@�Қ��h�W��4��?��?����mŝS�r�\��qC���6�s��[!�-�Z�%��[�9d���6��@��h�W��>�����@���Z�)���9^�nO<��<���f��ڴl����u�q<���J8���hzS@��h�W�ׂ��9�"�94]��X��r�M�� �E������)��4l����zm�@�Қ��:����� �^\]^�w5az��mў;k��E@`^-D���<_H;�O�X�����}~zm�@�җ? �� �K(( ���M�$z�u�w�ƀ�b4����P���l�P��@�Y�^��g�cЈ	":N�����$������,n��<�F�R�)�yf�.K4=���Ɓ��j�
���+0$��u�4��@�Қ�)��]�������k;OH"B�·����8��Α.�g��W\�V�sk��Va�a(�rh�f�ץ4�S@:��}\�Q"I�I�I�^�߼�CO�*iހ.K4}�v �	�7�)�r�^�[l�:������kq<rAbr67�U�~� m��9v#C��q4D�3D�L�����u�/ (���)���@-�hzS@��h�W������u,8�ׂ�Ω�6�ݺd�����Dh�0��B��v�
T�<�P��yz.�h	,F�Թ_�f?P:mށ�걿�$d�m�!�[e7�ċM;����b4�rڼ����2����@�\�@T��=135I�f���O� ���q4�pJ8�
��@�Қ�S@�z� ���Q�&D�q�zS@��h^�@��e䓧Pw�>���hl�(,(X#Xlښ�"����a"Iu�A�$Wu�6��)8�p��YVT� ��Y#	i�GI0
B1A
���R�c��L9�4���5[�O������D"��D�*#;	$�*�EX��F0 �5>Y>�ZFУlc$��bu00�nz8��m��U[j����&��m�	�&hycm,�[��v|�h��[�n�m��T�i@�U�V�.��$�e����]�V�E՛����)�5у��\rtH��j�C ݰd-�)��,b�{[k.\�b���m�wN�l�kX �[p�n�_L&6x�R[��h6�)�u�'���&Ū�@W�Wn��	 l�x:�ז��b��1!<��4]VqJ ��/}�����2��m����݁@�뙍L��=c���󧴡�	T90sWD��̕�V.��g��c�q��zgX;V�u����	����g"ηF�n�-]�G�wn�;<S�m�8�3��X�,H�.ˇ��x��U���F	U�ղᶮs�\�q�z���ҵk�T�Ӗ��:��RD�ݮ�]��xI�h��=��[�D#����l7b78v6��ڗȖ5��;j2I���,�$�ٛ����4�&YJ͈���Hy��Zy��$�ڲ 9Pt[d��D��vOH*����%�����V�'*������t,U���d�su����k1Ի���u���/�CF��<�����pf��5Uڀ�]l��[(���z�ص۷�Ҍp�p �S�"2v�����<�u��ڝ���W���7Pib�Q���\�;\h*��E�g6f���'h���oYn��t�N$N�m�}� ��Km#݁�c��髪S�Sɬ���V�K�N�Q��Yg��Uuu�=�\�.�=��� /E,��h����g���q�T�T�\!�[\�
�	q���mPPm�&Lm�����+F�	�/�[�bیUT���{�����\�˳�+��ձf�B� )�cJ��vv�+`�ض���t@�M�$���J�l9����E�Z�1��c�y�l��#۳�g�fkXv5Ri6�-�Y@HHԐ���V��ݐ)^eXv��m��dz�C��IR���ڤ�l���o5C'hѣ{��)�q4��0D�)Q9Я��ҠD"���9�3+���Pwf�{r�ۢ&��b�)��jl��԰/2�3�N7k�u���7c�&6���hg��[`�i���j��¦v7!^��r�om<<p�G��?����dޞ��a�Zz���R��z{v"8���;�(j��ɻR�ȸ���<���mp�{]X�����&��A�u	\�/�v�$:�T��p�dk��VLK�Ãѷ�O�@�8='�i�\�snu��#�xi'��D{Fn�/��Q]s�n#�� B��)[�m�]�9s��߱�˖h	ZU�r�F���R���$'#cp��f�k�hz#@Ib7�"#�31g?Vz����,2�����=���@�؍=1T��h��4}ίrI�Q8�,#�@�؍%��:�+����D�;mށ�2�|D%� D�JC@��h�g�b����n�]��;몮Yud]A�;�զu<[Y�w>�C'�h��3�'w����ִ�a$N`�x�C��/��Umz^��-���
�q68�p�Z�[�$�s3\����(�����?���ƀu�4�%]�D�I�9z^��-��׬�*�� _u���#"�(.n�334��h��4
��@�Қ=�x���ln׬�*���Jh�M ����F"E1���d�<��p�+m���37]�N�mˍ�=6�LP�7Dn�ylrI�Umz^��-��fy�~�M�*�<x≨�Ȝz^��/YM ��hu�@��>p��L�H�R�S@:��<���y��y���{�=�@�e4��Z�4�.̬�30�uI�������^���
�q<O#�	6��@����13
b	����g�x� ��h׀u��d�C"�!I�.�ԉ��6�7-�n[2�k�srY�X?�~�� <��2'#���>4�S@�z������0� �� ~4�^�阈�4�@t���b4ܢ�^������N+��u�@�Қ�)�~�K��1�xA��A�L�Ӵ��	�f��b4*f&&Fy��>�*�;�#�ǏQ�Ȥz.�hi�? ��Z�J��������M9�-vX&2�;'b<�щ�#�q!���ݻ���N�\q[h�V�b���:��@��z^��?{�k�M��$��k���<ď���}���)�ؐu�`�i�qA'��V��7z]���13T��h�u��;�C��"r8�zS@�e4_U�Uֽ��%^1�@��h���k�
�נ[Ҿ6�$!�kg����z�����:xe5�a��zz��n�/cCw���v��1;��p�,=�NT���ܔl:5�}s�ΰ��p��g��9G�C]M]��P\k��&��ӷn��<z�Pw:ª�n3�.��c��ȵ۵��Ȓ$Q�6���a��(뎎�.�Ó66ce]r���m�8��2��m�D�+�B�[t�}�y�|��2U��.���u�t��K-��]��'eF��Ŭ�ӷM�d���rܹ�!����z��@��z�)�^���;@S����Z]k�-�M���-}V���n�<qLP��R=ޔ�/YM��hu�@��;�e�b� F)���-}V�WZ�zS@����7���$��k�
�נ[Қ�)�\��_��n�Ȓ�2�%�f΋�9�{u�N��B��t�nY�F�ܒ.��=�? �7z]��,F��� _\�4��nL����-}V���3�H�f����*�^�޾U�A1�@�8��S@��Z]k�-}V���+��68��(҉�@��Z]k�-}V�z�h��Q)�C����@��z���/YM��h�uMd!�d�УɎ��K�A�V����8�[��i��\މRU�/n��#y�@��Z�)�Z��������x�Շ�5��Ŋ@"��-����-}V�WZ�_U�{�GX�#�Ffa�%|�@U�^��a��������鍘���}Z�v3@>⒂��ؤ ����
�נZ�����-}V�_L\�4��7D�q���@�e4_U�Uֽ򸫩���>���N<v�����\���gk����:�l���aps$ppi�&<��bqh���oJhu�@��Z��c�s�(�4zS@��z���/YM�ʒ��<P��Hhu�@��Z�)�[Қw)��c��Ȭ2�2�/A��x�h<f��b���:�"�(��$B�#�!V�d@�TBQ�>���߰��r�Cٷe�]4��%؍W%�%|�@s1	߿7���<HG��!m{=!c��y%�кG%����z�ŵ�ճ�I��+�,��ݞq��C�}gƁW[�@��Z�)�����D�DL��W[�@��Z�)�[Қ}'r$����'#��_U�^���)�U���;��Tm�&<���qh���oJhu��_U�~��k7�19�6(�4zS@��ǠZ��	�����J�S�K�ɫ6]j�9���o29�nD�^{{�+K+֕	h������g�%.�m�$��h��ؓt������rnZAwR;��qˮҭ����m��.�T����g;��9�Z���+�p�:A��Z���hN�<8�\d��L�]ێ���X�h�.�wM�(�e�묦!z���L>�䲍u��X���f��:��[~w�HII �N>�B7+ѻ3�Z��m�
gr�R4.�O�x��5�l)nؐd��	c��,nI!�|���k��S�? ��>4GC>�<qDEȤǠZ�����-�M����e�7q�Œ�dqh���-�M���k�z��Bd�&0�H�h	v#@U�E�	_*�s1M7�4���&���D�8hu��_U�^�s@��怳��������%�-���,V��;�hJ�����L�K��� �s"JH��"r9���@;�����@9{ݏ@�����a1��2����%��31��1�%�c@���=��h��q��ONcQ���[�s@��ǠZ�������P�%�#ȱ�#��U���-}V�z��޻�.��;��P�E&=��h���-빠U�G�^|���:�V9�J�-Q�䮝��M�������\�EJ���y�����WnE�-����w4
���_U�{�dt$�La����-빠U�G�Z������T��MDd�0Y��*�E�	_*ӈ�!T��19�a�{�ZC����b��!t�#��ҡ��N�; �ST�C{���|jl�D��ݐ��tM���J�B�i&�z��g�>�6�H�����1���S���<C��*:�M=���I�aH%#qP���RI!��C&�:cD J�4J4�a��ZU HD��RH)�@�����G�hJ� 	6�/�4��|��lH4em��!����:1+߂��fn�S��*l<,hJ!	���,�^`�lHx����dL�2bR��ѩ��0f(!p��h�b 6��� 4��6? *�C�v ��8�x :�,^���|��I=���$�>��k5
��.��*�3�s3M�u�4�Ɓo]���=�}����cɋ&!��z��޻�]�z�)�wѷ��0�.s<j5�u�S{X��K�[@u��s���ǔ��"l�S�\�p��"�L�-빠U�G�Z�������\x%�HcrG3@���@��V��-�.[�f"&j�\���7
(�<���|��@�e4z�hwQ��\��ǋI�4�Z��屠*�E�}1�Lˈ �PT��BD��A`�I�F
R%	��#)I��ZK%�l%�Kh0 �X��"�hb7�g���>~���]��E�Y��h���/>��-}V�z�h�pVݎ��J���u������{V�<�����ʺ��\��7R��*N���W}���>��-}V�z��޻�}\�܀�Cq�M��Z������w4Ϩ�����"LY18���h���/>��-}V��8��7���iE&h���*��-}V�z���2��,y&nH�4]Ƚ+�Z�4�lh��& {��~�ˬ��Gu�g#u���\`�&�n��<�d�6T6u]7D�cP[M��::퐶�F�Ѭ��ob�Pph�z�oZF�&۱�샇?���s�t��ZNF�xm���+� 3��s-��j�&���^�2��R��lB�,�X�U�D-m��[��5��u�1p<�ؕv�StqF�<����4���]�4]���J�����k��w�{��q!�}jU��礭����mD<v��Ϟ�C������iM�8�ӥ2���Z��Cg�;�r[\�4�ȭ�G�w,Y&�dqh����#�ۚ�߅�Z��ޫ#�6G0��$��o]���-��h���{յqDۍ�s	��4
���_U�.X�M��4�+�xAW�U��UI �_U�wYM޻����k�Z�(&?$ ��26y&1�]lT����Wuͱ�sa���B�b���aS\=s�N-��h���oRh��@����7���iD�[�s}��0Sk���}�>��M�I���א;�����VX�L ܑ��oRh��@�)�r����<D�#�D��_U�wYMޔ�=W���=�v,�i�8���kY���zWʴ��W?�v�u�ڳ�f�l�w�J�:�]�s.���.>�r�d��[���\�ƪ��ٵ��>�Ƚ+�Zr�h�T���LQ
`�4U�=ޔ�;���oJo������2bq�M�&�$��Y��I�f�rtM�@��qQ1��L�~ױ�*M�w��]M�S&<���Zu��-빠z�Q���@���Ǜ����iD��屠LzVy��������Ѷ{��X=�2rb��-etr=�萎�qm���'��Bv�ON�ب��������f��G�Z����h���9{�ھG��B<q'	�Z����4�lhˑ��j����2���lR�O�޻���Mޔ�=�dw��La��C@���O��7�&g���T>E ����<����@:��|%��D)��4���މ��� ߳ƀ�-���R�N��(�l(<ܯ-�g4������-�/:�RC�5۱:]�r��ޔ�;���o]� ��&�޾����c�LDnu��-�M ��&�oJo�g���/�F�x�7Q8h}gƀ{z�@��4�)�~��T<BLyrI ��&��b4���6����wNr�/#����3@K��!'��k�?>���i$�x����I5��f{[vMO.�ϭ�U����ñ�:�\�ڌ�:�gGR�v��vNSB Wg��iy���³&������y&�4Nq�6݉l]t�{R5�9�<v��`q�TY�n�%��J��Y`�<*��T�
��ּxw����Ͱ>�gq����[��v,+o�a�k�~��}9�����؞
.�V�Y���'�aBd{<�{��ȯ�T07���}�]Ke�ލ0��-��ƞ���G�av���2qpY���]^����2<1d�cM������h���{z�@��Z����G0��$��oJh��4_U�wYM ��r�A���8h��4o�i�311T��h�f���W\+8��ȣ�@��Zu��-빠ޤ�;��1Vb��G���ŠwYMޔ�oRh��@具ζiA�vM�=,v��vs��g����êۉ�Q��\�N�!��K���f���13��'��>��~���1M-�l��~}��s�%���� �Q��B�P`H
PV�Z��0F�V"V&��0DI�;N��3@K�W�ͫ�xd#�D��_U�w[��[Қ����z\�ŋ$�l�-���ޔ�=W��_U�{jR��I���ޔ�oRh��@�s@�����3w�h��+#^p�v1��v�=�Y�ٰR�.���3�ș��H(�S����@��Zu���)�~U.y^ �ȣ�@��Zu���)�ޤ�-�A���1�""qh�S@����i���"Gj�k�?w�h|��@���Y�LrH��(�4��.Fh	_*�����@�Ʊ61&8&����M��h�S@��4F���(9�X7�X��b�˹���٭���E��=�	�[��k�˥��0�G�$�4_U�wYMޔ�oRh�apwLY&�dr���335Ck��3@J�V��J����1�9��)�ޤ�-}V��n������&����31U�34�:�;����*% ?� �k;�rI��f�~�5���rBh��@�s@��4�Ԛ�qWS���L�H�M3�T+v͉�z:ܬ\sq����Oaxm��$b��G��Zu���)�ަz"?P7iց�7C��.�3*�,�����F�����晚v�h�lh��LOHy1�5$��oRh��@�s@��4Y˲�&1̄x�N@��Zu����h��4˰�;�&,�i�8��w4q3��| �/ ���"fbe���J�*+��**+AQQ_�EE�����O��QQX"�
����**+� ����TTV����QQ_�EE��pTTW�QQ_�EE�**+�**+���e5�]�E�E;�� �s2}p��   D
 

�
 �� @�@*J
$@���}H�    @@��!U(�PTIR(�PJE(�QJ%����AB�	P���"��%@B��   s��   J	b kN|�]�w�*�e֜����osW� ������ݽt�j��y��� ��������7���S� ��\Z�ɯ���t�R�������xw��Zrj{noN��  ��     i�*���';.mrӛK�{�ԯp ���4��VC_i�5JbʕK@:���U8�� �Y��U��U �TP b    
 � 4  
 
 @  Ԫ�R�� gU*�ԩU�uR��;����*� ��     ��ΥUci*�-I*��JU��U, j��f�T�Љ�v�^���W��וy{� w]�ޯ�����x �=[^m��O;�kv��zy��[� ��nN�V�ח�yn��y�]/��  (  P0��}m�zÕ2S#A��}K�f�\Y�\ۥ�ׯ:V��
9�m���t���  ]w��5s�w��χ���ݞ�}�.[���Ϭ�������R��Թ�>�y4��ﻩ^ � P   ��� �>�q��\�=���i]͗I��{�X�:\���M=���.�=�n��/-���sg�  \�{�o.����� �E�-�t<�'\۶�7�����������^�y����{On��tx�B��%H�� Њ����ʔ�   �=U*iF�  '�T�Oi5(A����2RR� 4 B������ h�O�?����S����n����:���ǲ�g������ �+��ɗ�����PT�� �+�tTW�QX@EN{����#-fV��MK�&# � �X	?�Re���а��f6b�A���"+���4V�,�3
���)ĵ h?�Ip���G�D���z�pM2��|�Pك��Y���f�o�����M�ԭQ�d�NFN&`C�O	�'�R0A!�	%�$µ��B�!=T�i�4F�=HI���0cC	����Q�k�m��m#t��24�釙���C��`X^��`FZ24���$&16q�再y&��47�6j_N$f����Ӡ�y���o�C�_G������ ��6�֘���A��f ��lf�m�&�݋�l�{8�ᤌSK��7�s[8&כ��qӱ�ÊH�̴A��ɍ�|4zym��z`N8h�q��8��.ki��9^xN�����9L�sXY�4���ǉ��Kk���l6��A������>�h��5�� ��~�,���H��`��������EL��]D�4[C�Q<lqP�S%ua.���DI���Kdt�/�D�PUy;�E�����^���Fގ��:�*�='�d�l��Xk0�xi|ILz��1�4&�6��Gc�,8xi�8i�7<Cq���s|04z��OM��p�o�|/5��4��5����{�{��狎�bJ'N��w)}Ċ��,���0e��.f�g[�($�@Y����a��߾'���`�<|&7��׺��OP�q�$H>[ȣ��q�8x�iه �F;#80�`�������1���x�`h�<$e��JB��M&����xc�j����6zo����0�0����<1ߧ�捯������Ѱ��x�f��Y�{��<e14z6�`����q�����H#�祙�6y��A���X�!$�k�$0�Q3lƧ,"0��Y�������H�/�IS� R��y�q�h�����=�����`��	��9������6����%pи�%�F"��sx�q�N������8���EW��X$R>�+�q}0�FTp��U��f$��ƅ��\o�Ux��i��L�|��V�I��9�ax���$ǉDL�)�͌c#��$$ܩ+�6��@@����>4l8��8C�J`H�h���ȼ�x�kzEb�n�MT-"�4*��ą��o���5APRW	'M�|�"c���L��*Wʈ	t�Hq��X�4�����6�ZM�dal�,6g3�"�,�\���5t�P�v�������kE�4.�X��C[��ؚ6���W����<
��aa���Ig:����p �86l�8�w��9��F$�h���3��|����C�����w�ϵ�R��K��`�a�8���q	��UR$ͯ�����lbrǎ�S�p4@ఁ����v����0|�f4�A8h<r0�[Y �3Aj3g�����#5�c�f��SCg<Ֆ�X�F%s�xY�/����o5��$f�郤O�%��BY}N3�!�&�c�����2�i��}��> ��߲�	!�I�w��{��L�����jȕ1#�J\�%�
R�H�ø���}��q�	�	
h!��B �!�4�B�. iE�  RҲ!��.��� �%$ŕ!`0d�\e�A����x̔@��6��J#K�88>/�)�f<}=L4�x��x0�h6����֬4�����H14�Ќ���1N���0�t1	����p֋Gǽ�z{�1/�\x��Z����T��Ըȩ;��̲��c�"U,�Q��2��ˬ�JR,#3lf�2q! �  ��g�L��r�2;]��+:���t�!gܸ�"�Vg�b�m�{�sZ]�|=#4n9毂�	#g��7��X�3|ߞ���%�Q3���,��B��2;v��F�0'G�o�Ϧ�M<=,�&��XzA�1����.�>�n=�dh��p�t[ּ����6�y�����nIM1����yx�&,c�VhĀ��XC2gcDi�o�Y�������3�AoI;#���7�\q�i��f��-��0#0�h ӳ|L5�5�5htol���Ѡ0�6�I!a�i�ͻ�n�A�D�0��fHb�i�󁭒NN�'�bx�a�r*4)��b��(a�7���Ѿa��1,WFl��x�h�b�!���h�a��K�CL	�=ᨓh@H���8����A�q���ѵoP�C�BSvA!�0'�#�I �_�2�cĩ���(Г����+�f81��L���Yu8��_O`g\�l�:D�k#�hp�D�&I&�)��'�|�AlH$�fXb0&_(�Y-v<9M��®0����AKЂ'+�M��<�V��r#�b2���L�LB�"Vqg>D�>��
6E�!��M�jٰÇ����C;�̌��>sz8���Ѓ$���%/���%F�rϺ(������.�$V	R*�-EE�������]��+X�.>�W~a��Q
��˜�LO�[�z2���ݞ�DG�2XG�HH�l�������k�����5�ь�o��7�&B#��|Fj�#*b.�z����7���8se��<��Ѥ�@A���&� �'N��f�o��{瑚�#���Z��s߼6|3�`����i.3���l4�'�t��%/���9���s��R�%��=3F��=�#4�`���V���J/���)gӍ'S>Շ�N%��3��/>\�]%R��*41�5�ChѶ#3pV`Ů��^��Ϸ�=���<0# �XX�3��c�1GJ]}Vo:�ࢵ����z��6�i�Pf��A�Xq��䏍�l��9���'Ќ#I>.y��}�>���0��q�������OO�7���A&���|�"��#<\6;'LSl���ؾdH���/�_�}��X�*�|���h~Q�h	�}�y��a��k;��F�s�xi"  RVA��B��I�2�	�iL��Б�D�C���f�3���I�BH=�]�@`��Sa�e��|O9
�
�ȱ #�AA^,H|Ć1\|1���`qbe0HL3	Oz��5,IT�ь�,LG��5�0�$dZ�e��!�N�0��E�gEN�8i�\��F8t|:#	�M��	a�A��p-G�H#Գ���LLf��Da�\_�c�q6'/�*A>��b�+3��N�-
Uس�����Ϫ��8Ăg$:ݢ� ���#ddh3[�>��q=bs[�fz����3�D��G��Q����J��c�T��!��E�]�;��qlR�m�B����Ue�U�X�2�ゅZK��fz��341����F��#0ͱ�'z�Y������N.�I��F�^�h�	�7��0�cDa���jʍh�j���ܙ�f�NhcA���sF��Vq��f�#8�PV��ChR�`��ѕLBc���J��$�kf�m���8��h&$$'(Ī�+�+*�#� �CZ�p�4�i��DŚ4h�̵�$�Fc��ը5��ֈ�4�h�3F���f���4٭ot�Á^�<�a���h�WLUI�(�RIU@�ۤR�Cڮw��{�{˵\|���*�y\�N�s�un��9���W�G�IdUd��T
ěw�+�Q(�.^.�g�(�%+H��!F(đ��������   �  $��-�  �c��  [@  �� ���`      ���N='es�u�.��+[���tGk��|I��	 ����ʷ�e+GlWl�K�F��B�#
�pUD�Y� ��m �Nؽh6�m�[��o9m�m��@ ��*��WL2�֦  �Ԁsn��[@��8 �۵�3Pl��t��ݶ  �D��c����ɫ����b�1m $	k�Hj� -08�[G)zԲ�l�� �   -��$�"�-���  �!�m�m -��m�����  �� [@  "Al��l [v��m�` -���    8	i� qmI'm�p�� ㍶�i;  6� �   8 �         �@ �b�-�Hsm� ��8 �    $  �l���� �i�b�lp�� � m�      ���tm� |m�8$�m!mq ���@ lHm���rNְ�m�!mp  �  [\ � @ 6��  m�� ���� 8 ����o��$8�($�� m��$Hm��m�       � -�p�ݶ�h� m����jn� $ �N������ �[mUTd��&�vԫ�R���o�6���+m����       8   -�Ͷ[@ �m�m� -�F�H���m	$�6��  $ m  �6 6�� �zJ��H���-f�e�*�m�v-��mmlF�H [@-�me
��
ڀ�8��ݘkfݛH[@ [xHͶ !m`����$�mt:��l�� ���(��Ts��������B�8��YZ���l��=e����Ԭ�2��ykj��s*D�-]@ �B� �v�:ً��U�[��� 	 �8�v�l�;m&pl�N����ԝ m[9�� m  m��!&��*����%Ul�
T  �M�4��۵�s� ��N	  6� $�l��kn�܆�$�'8  	 ��&��Uŉ(�Ʈe���%�� p!4dZ��,���[v�� 5����ƻl�t�Ӂ��M�J��̗�6�Im��;ey[5FUUmդXj3[NC�<V��l��/mڭݰ  l  	 ;��n�Gh����n� �8$��[rh�� ���� r�������W�55�L� �������UUJ�q��t�'��m ڵ�r�(��#�c��w;Q���&��5U\*Ҫ�m*�J��`��$:Az�J��s��4�5F�� �U�ݣ��ڀ���
�zx�欓ܤ�R��$ݲ���A����>6��nN��jr*͗��ƒ` -��$m��[�\�����.�+I��ڪgA�x��M��Ck��ۮ���K��9��;,�\ rb:5=rriB��v��);s��Ӹg��+�ն�U*�Y���8�'��һ����bgh �69���u����O�l� q�(lUJ��8�w&v��-�;I��ڷ�si�7S@P �Ȼkh 6Ȳ� �$�uIm6��n�d��lI  m&����鐁n�d�v�96uUUR��R�A܅�kkln_f�B�Il� $�hX^�ܓ^�-�h�ةx���	��-���4u 	9>�}��v�6���j����Ս�!�R���[U�V�C	��݀ ��7F>}>��։�H�k��9����z���v�6�؝e䄉 $)W�b�%�2�^ �jn��$֦sH�km�q$�1"H[Xd�j�<��h�h �lv�$�s6�΅ƅ�xz��j�!��	��]&^����� v�`H��M��S�۶�h �m�  � � �z�ybwK���m���h-� p M:��[k�mPq)rչO����T�$[@��m�鱱&��m�-6 $ �m�� � �'���&���@Hm�  n�F�5�	)�y�[���a�)��"�NSq8x�i��ٍ�r5�[�A%4�i�Mӭ�Q��V�p�*�v궴ޞ�UuWUH�Ui}�l��p p��Hu�vGAzմ8m���ֻ@�cۭ�����'��vUeUZڔw`�v�nrKn  ŶCm&n�X��l����S[v�6�C�ln�wt�UV� ����$���ǒ`m=;d��H�V�M��v�n��	�냀p�,�l�`�l�i�l�$��PS#Ѷ�۔��հ��f�=/^&�ͳ6�p6� �ɯ~���^�}��td�۵��N�-��Pv,#UuV�Ni�U5]���C��������,�������(��V��8`�mR�5\�ʛi	8-ѳk @8�t]$MͶ���u����=��	0[@ ��i�`y!J�i����M��Vݴ�lg][TkʫE�25I�m� ri���ur��$��b�(���u�i0� ����OUg8k,Y78�m��z�ݮ 	��VN�I��	�WV];`m���Yd�U9�  ���d<�év[��Bdvy�������e�mlHl 6��a�  4��e2UP
��ݢ]���R˶��J����e[j��^j��ٻ7*T�hp�*�O/5l1Ͷv�<7ceo#��@UTC�3wm�h�L�&� ��K��B�*�9�hc��ۧ&^��Z��4�N��ͪ�PEԤ�m��-�����R� �����-K�e&n�MQ�R�4�](	���퀑�h�Y@ $�X�Y�� �d�]m��@ R��ԣ��ckķ�pJ�T��ˌUP��8q�v8*�C���*�3�Ku� %� [d���M���8���J��Pl��t��!0		��[e�oP  p��\�S��6��v�`��Ug����a�m�ݷ	a���d�>���+�\�'���ݪ��F�m [@m$����vm��l N�wc��m���� 8�7��`�"T���m���IKjBF۴�  F�����Bm���'@M�Y���`8���O��k�,sH�:�9{M�  í�-�:	Ԓ�  6ٖ^e�FԪ�T�UmP�m'k�k�   �n��� h 	�m-�6���AT�qΪ�	vYUS6�S˸�sR������++Z�sm���  9mH6Ӥ��8��m 6݀�Vݙ6� � 8[&�����+l<J�u![[@KӖx��c���Q� �`  �(6�)���U`�gn�v�d�m�KI$g���9m۶ ���m{M� �@H�Ŷ�+j��[Rm�'@�u�I��U��^�4;
�P/,��[��Ί�
.��B�V$���&�H/b]�Ǝ��d���8-��m�I0$6�-��,^�Dk�xְ�����<�v���/ʙ�� [�@		�č�[��Im8Ho�[�,˿O���#�Mu�y�P ]c�J���q6��y��R� �  ��8��m�2�Wm�/#Y"dU��vm�/
p*��橮ڔ���7Y�m��2��]��fZVZ��?_?}��<t��J�2(s9;UP NY�[WM�^�       �Jm��h�K��m� ]�n�$RC�����ۛ6���$%��` = l��M��fݰ��۲X5�#]� h����-�-+`�G�#��-  ��Hl(
��J�V1W �M�im u�m�l�5�psm��� u�   ��um�o  ��[�l ���� �J  Im�v���-�ɤ�-�/P  [�l� '5�l�$	$�[ur�Y� 8���jTz%؀�����%�y��t!5*�<�
��lֱ�t�٢�(�r�4U����⼐� �h�&�4�C���8@ p l   $� �@�]�����      �`�z� -�    m� ��    �-�-� �  �	  v�3�: �m�  �   -��6��L-� �l5���͝j��0��U�2�IDʮ�n��Z�cu�jĲ���9m  Ht����     h$[M����
�U/Nyf6��7�ߙ�"]� �[hpڶݶ-�i,0 �Hll$H�t�'%��(�-��5�A����eAL��Yv����<�xՊ�.��J��UYw?�I��m��m��@���?���B�=��x���Sb��v��\E�Gzb�<_T_�À<Q�%`e㊡� |8���F�@�|����`� z"����^
��)�)���t�v]C�b�s�@��1O���@<����:?D � 
� ~C��FPO�'������A
�P��VQP�$/EP�E� :� �A=R�:��T��@1T���	 }=DU�^ ���i&P���ZI�`t�A( q@U��UECb���u<����tEz��&W�">:fT6
. ���A|�S�8:���!��O�Z!%�P:(�������t6� b �S��є�T��8i���Ej� � Ǫ�{U�G�b��M������|�'����*H��#���Q]����B1Q0� ��������� �J��m��ݚ޸H�k.�Ħ�iU3]c��;d����$ĺ�b.�	�����L]����R�Kj��BSk2���Y�D��vZ�[���v̹��ҭV�@,˦���6ۄ42���+��Uuv(�l��gf1�j�*�pU®�	���0i-UV�.ێ(�h�xʌ�-�`[��Hdq�4�6r��69c;˼	^��Mt�d�2vM��0㳹%�j��\pgL�^�n��p����BPJ�tv:����p+M����S�x�r��֝;%�I�f�)mtnq�B8i���lS:���9ܻmV���k�C���=���/"�)-�j��V��h��ax��6^����%-��ë�n��Ru�`8��tD��������G]�� IW�WX����dpq̷��ٜ�'<<E�z&��)��;
�=�w&ʖ�C9���Z�g������ ���b��Z2�K��ra�������{b63�O��n:N��E2Lm����M���
�ܻ�D���\Y�c�b��W=�:7��#Ż6�&6r-���lb�tl����˸�U���=�{c��X�96*�������r���v���s��Kv �/�0W7kF�6�;x�"M$]�8�����k��c���#��v�6x�NA���;<)z؛����6lDn��e�T��mɶS=��j�a0�]-b�n�,�]��\!5\j@�
�����q�Rۻ8�9v�-�-m�W���:������9��&�ru/#��tAq�T�%I��%H�[�Ώ6�`ɗ�l�� ��\��dUм;7d�J�� 餉.�ڽ
OK̶#��aW��٫)�P5�)����Iym �@����Ƥ.7d�Z#�Ju�V��vm�Yq���An���)se�� 
��UV5��rS�	-�4�t�s�*�u����m�9�*K-�ĳ�[�%�I-Y�5�Y�ޭ�Q�|��
���aBF��"�����*��'@dW����ۏٜ���pq�dGA
�k"�st��i�F��Wь�y�60ٶ�mux�����o�F�V�٦M���T'7�)�n+����u�՝i�c�\d��G��o,�g����g<�����mݟ:�q�js[$��+*5tn���3�[ܰ]�!��Ԍ�V���Fu	�Q��j�;$�pm����\Be��o{��wxx;(��|�U�3Eej�R�p�w(��vx�;�AC;�s�9��x�1�Z����v���X����ɴ�O���, ��⪬$B��Ww�};�Y�jC�'ր�j ��$�����U�{fQ���	��nj ��=rG`g~͵���t7`��. n鹿NsP�& 'c��|:�Yw�enї���'9�\���@���Y��%(�������I�' 8;!�Z[��9���$���ܑ)1	��+/���\���@��s���䥣R�E
�(i8���W6����X@Xz�#�W�8UUT��~��T�=�j���^mAB�*D����ͺ��l�8�5�ך� Տi)K��Q�)% �j������ ;�Z�=1�۔"�T�P����U���H�l��L ���fPi�,�b�pg��y��QODq�;v��U�8Z��J)6%�rG`s^j�3��V ��@z㘀}RZ��Z^�bͿ�R |�=rL@zc������fט DL��'*�77�����r�a@�aR�|����w�ޫ{�u`s2a �HQ�Fff��$��9��T�9�md�mJB�U!CJG`qnk�33n�;�,-�v��帼4�~4���\� li���Qu[��t���<]�s�;k#�%Jt�IPL���B����nﮬ�<���9�	0.�J�۠2�l��ݤ ��@rj��7Xf������H9%�s7e��b>�r|� G>��%#woh�ƒ�m)%�Ź���f�Xw6XJ����A��LTO�� ^i4��z�/ ���3��Y%T�X\�� ��R |�95��1�]?��㿃�U�0���ֆR6�q�����}�ޝo79��m�/[=��t��ŝ=�2��^ }���>�ݯʹ��;��Xs`�	
n���ے�9����였���梃Ҟ��ܻ/�ٺPf����b���s��<��b7���)b*]�`y6�w}���ڀ<������o%]�ђJ�I.�`9ݼɴ��������ʽ����^�ߩT��qh%!3�VT�H��E�5��萟;��]���F�U vM��mA�ַN�R����8CK���G���]�x���ɟS�X�\�Y큁�p۳e:ڰq�uXӝ�MWY⠛ǡ�v�S�]n�h�:q����Y�]r�q/na�K;[m?�ܿcn|���=�ImZ�B:-zݍ�q�\�
�I���.�/+:�+���⤃\�	Ii����:�k| �n�U'�읊�Y5���b�R+�Ń��nv|ܚms<Yd[��qշgwX�����7 �5%n��#�ScDCiI,.���u`�l�f�3����\m4�37<��H��@rj��b���J���NU�w���9������;��V;�{NEM�m�Dy����@z�L@y�� w9�~���aƢX�y��g]۔g��H3��znB��^�%�����Hc��ݳU�_I�7 �5 y��tI
%��؊�wX����ORo�����K���4��w��7v��7k �bKV�GLT�BJIV��� �sP��n*@�y2�6�����$��_|�w},�����ͺ��6X�ST� �M��RK������U9ǀ�j �P��_�0ԃƼny�_92�V��*O'c�@.�m�&۳z*�	����\m4�*) ��� w9��M@z�L@wt�awB�Qt��ـ�v��i������ ��y�̚X�A�97Dm�D��ʯ>���^g��i| �v�;�M��w6X��Z� _
�(�X��n*@�j �sP�HA4�"��	I��ͺ��6X3vX;�,����D��r�Ҧ����-ۀ9grWB�n�[��>��S]tX%(�J��II*�9��`��`�l�;�4�
��=i�E �RI`rj �9�o`�=�j��~��웴��L�6�:��$���X̚ s��<���Nf/�K��/rU����7��� s�����x|�]a1����k��|��h��r��.�(6�D�sP���=�j��K��I���>�$��(�L}ɬ�]n��Vsj]k؝���v��5�nh��m�������@�5��ݛ,md�d�/�RI,�͗�i�!�������ݬ ][�P�T�JB�G%���K �se�����9��`f1%��Q�'���������@F��Sˉ�E �R 9������.��pk�+��������MBIJ��J5��0m��Wd�fk6�+9�Sa�Lk�m���s�[<�m�Es�T&�E�v�c ���vj,E��u7g#�<��;KG<�\[����s;�\�s\��8hwN��:��紝���Ng=�~��l!����n�����̶3�����(��g��n�Q����+��n���՞�g�k���9w%�٠*V�~���{�Ͻ�w{��]�(q�3�uܙ�	�re���-����n��!-�v�f�]���*t�Si9:��K��U����`��`sJ3_�.؛cN�
I�;�|��s���=�j��wtUƪ:	VWs]�s3e����H�{����9ה�����F���75 {���9h�{1�Oja�rbWu�sv�6�O�{���|�]�va������i�e���U;�:�6[tu���[�s]&W�Z�*�Y�p��T�JB�I%���U����`j������Ku�-Mz��:N#33[�U�{�u΀mP&a )$�J	IX".�o>�uʯ��w�7�
��f����H �v�و�&�#�-��b�ٛ���ӧR�H�v���q�����՛���f�ϗhI�Ӳ%$���L�i��w��w}x�7o �I5��������Sq�۷X��1q�q�s�vø[ԙ�w=X{E�[7����6ĝ=�[~۟b ��t����-�z=�"�荹(q����/Ԑw=�`w_���� ��:�H�!�.� >���v��/�Iq��4�5뷪��b�E��R ă���GЙa�v�k�5��$s�	l�SN�4�2���aiD�����"淭�H�)���s0u��w�DH�
��W����
���@1_ �DGr�z���$T ���y���W߻�|��7t��HJ���KUU.�ߋo��s3e���K��KQ似�o�BJ8X]�v�wwӀ�zX�oL�I��[�TYD�Q*袙eτ�OT�y��L�ny��CŮ�tg^�q��` ,*�t7s�'ڀ=�j��]�vw5��������9���7!���vw}X�n�y�s������li��p���X{�,]�v���z�	 �URӝ��6sv��wo�ĸ�m��U���ߞv�]�۵�Z��r�v�s7�L@:�s������Ic�����DE)�F�-�\`�=��Ʋiy����7;�[��Ўu�LX��Y�Q���=�j7�@z��@K��`�SM�%JB�I%���u`z��@K�1 {��X;y.�3��Fm�w����󘀗�b �9���XnR�I@R��"�5wu���@F����e������a�����=�j7 =��%��`�mn耧�V���Q.��vq�Mj�����(����k�<�@VwC&�r�����v� ��7)�ml�L�`�<����;�ؤ���K��t��9u���W��^6����:��[Sf0f�k��h�����f�U8�r�2���g�8l�#�Ӷ�<�Ҽ����C
][��-�E��OF����L1��z��.�����J��{���x��T��6�V��)ھ=TRprcTk��[<��<�:tt'L曡z�}��U�6������� =��%���=�jpS��*T�n���B��^j�5wu�;�,̚X�A�N��%���<���sPo`��c��#�dT��C�I,�͖3&�:�U�s3e�hn�M1��)
&����r����=�jܿ~~g[cД�n�T�gcGO�u���1���:��hN��G]6܎���l�a��- y�������~�U��~g�[���RJE`��|��UU~���sP����-}Wd�߲7�m�pI�`���9�4��U���|����2���������7���- y����=�O4HUh�($qX��V�͖�����U���������5#L��Z�ݜ��6��,�XNz�f۷E��R5R�)*N:�.��wvX�5X��V��z�Ο�T��6�3w<��9h�r��k��wJ��$�HP)$�7j���_w9hLz (��S�����Հs����+6τ�JE`s��@K�7P��@y㖀+�V��!WaR]� ���x�I�9���׾V:�U��1V����9��Z1�M���.�=QhJ�l�c�;v�랪���҉��r��s����<�`s�5X36��̬Z~q��q��6�w|L�ZݎZ �r� {��:�D��U%�+�y��՛�X;�,f�,w#U����F�Pf��[�u {���� u3��v�k��슐�Hr��X;�s`���--ɺ�'\2�3&R�lY��nx���v�fs�aN���7.:�n�69%�p6��nؚ�m���_�ݎZ[�u {�����e���M���^j�5f������K �iK5
$!R��"�5d���&�<��ݎZ�e��̥�i9R�9��`s6i`w�5Xs6��̣5y����u ��������--ɺ�=�jߪ���8��.ܳ� ��t�{��^�lr`p����)���qlH�n=!���D⚃���9�c�ܫ��uls���=c[:��ӥ(�km\�dR�ys��ܲ�%�:�㵬�vw��6��<�h�v������lW��⿿;}��m�o�B6n�,NGB콍KҦwQ��<r�;�A#Eg�:v��YxHtr��:��.�;Eڳt���������﯏�;�%�smݧԑ�a��cv�{h����|o���m�Dtt�l�U �DM�RPG!�w_�+ �wU��ݿ��_@���`��E�.){��A�������&�<�����`]�OdT�)!�$�`��@yȩ��b ��j r�
/o.ʻ�(/7u�"����������)�kh�aN1$���b ��j �9�9 
�(����f�%�8N�H#�q���Eu�K�[��ϛ���2h�@qճ�~�nnV�s���R��b�e�ͪ��D*®�� >�v�6���& ����˟w������w>ݒ��Q��8�`8�N���w}�������^[�I`���9Ѫ�D�U%nU����`j��,�͖��w}�U����y�RUd�8�	nM���}���*@�5 C�;�~s�V	�V�G4�ݺT���tEnG�u�jw�x]v����.��y��7c��f������>�R �sPܛ��!Z�"]�*�� �����6��37����zK �we���Z��G��%]� ����6wv��3���F,�,��ՀsR�5�!R�����&� �9�9 s����J�48��K �se��ݺ�w6Xs6����TҚK�n!�{ny��_96R�u=�s8y����l�ݹ�e�k�ڡ��q����N���f��Հs���9�ږ������t�&ҧ 76���@�+P��@{�T��Ģ�EITm�Q#rX;�R�9�j���sP�2�n�]�E�mf�� �9�s����A����X=�ГbL��'��'��%������:(R�,w"��sP������R�ʗ��<�u�M�St�ֱn�`��!rxی�θ���ֆ�i�Ȣ��)��bQ�V�����ۼ���~m��s��X�H��J�*T�9%����_ꤎ��;����w6_�#+5(z4%
hp�f�:���#��Wg9��s�6���#�#m:������Y��ʰ���w6���ﾦ�~�h�{�R�J$T�U� �;��y4��w��*��߷ʼ����Z6��<L$ ���*N������00�C,I)EQ$3U�1�k�l�<6b��� ��|�1��B�D�(K J��L���.����TIxc�TD�#���#��U��$�	@2��	�3-�to�Y�dI@�Y`d�� ���)���#&@�0p0��14o^����X�)Sd�IÑLBL�o|t``I)�`��0^ؒaAb8A���`@a���r6��B�w��>>5��ŒT�T�α�`X���c�zo5���\�!,,�V��(01q���� 2FJ#VV�	�120�1I	 ��ӺN����π[%ྲྀm�=P��Ue�4�嬠���Z�Tk���6�����T�wd"�8x�9�����UM�����m�s)Ӂ��j�sB��S��gn�9=��۰H ���eI��n�l�Z`��Z��S��g��d�IU�]��A�
�@.��#��-U�@Ul�MWn����A�����A �ٵ�+���)ŵ�]нj�R�\'$��짯���$ړq�G=>�6%έ�������@)
��ªO.R�Ⱥt�/�T,�6ڡ�uSr=��9��Ovx�������m�IIJ�A@R����R��,ct�&u\�sh���9�w
����@r1��M|-ﶱvY8��;l�ݰ
��7%��AM��FLqil�-���)����\�T䱵X����.U��1���[X�Lv۳��,��b��y�<�������n��\��J
1��B���=}HӸ�.�YS��u[ZRk�i����r�/G�uˢ	7n�^7WV���'|}���ѠV������숁<;st��nێ7Pgs�63<aB�0�r���5�g:]�nŚp�!�������V�ˌ뺴�{kg�y%��m�nv��p{���Ee7�Q�n޷�56x�!�[F{>c��u�-�b�n�m�q�d�P�Ntm)�pƗa�ɲc����;(�n���-v�����cjSu�R�]l�n�Mt\p�-���j����'H�-U�2@an4An-plR��, ��N���̭T�Xu`ǉ�������!��Y^݃L�]#�L���{�4�擟�m8���tpq @vv�s�����g�&��^��� �m,�wFz���V���ܠ:+e$Y��Bm�m�s��:�hT�m�F���s�6�`^3c��"5s�a�&sB�誠Ű6�u�O+Ug�U�rqWJ��綪�	�;7],! �uU�KU����5Qd���v�d�e��f����w�<~����� �N����=�����߯�����M�J� Ƭ�(7d��rW�d�7`+W[�I���GB��h�&���Y�N��y����X^�e�v��w �܀�1�Z�ڗ�ˮw=��l���]yֈ������X�x���p�5O�c:��;u=�b�񙰢 A�����>��+l�F7���;n-��q��rV�\�`�-&䙔�t����䭂�u=S�Xf��v�;���ǻ�}�뷾
��	�%ɓ���nzݡ�sD��ؐ���6K��1��.~�k�����ږ�̓�}�Z�=�j�⯫�s�@�>�^��EV���^ }����o�UFo�]X�KWsd�RFy���q��R�,秋 �se�K�w�Xsޖ}��ji5E9C���;�؀;��@�5���,��.��6�3wPs���&�=�`�;��`s�kUt�N&(��$�*|�Ղy�
�vlM�!�m,��m۵�7�z���0E48F�����٥�w���;�ږ6����兑��D)' �z�`�'��_4�Xw�����x�7o?�nC�*-�R�ʩ+A.� �wڀ���@z㘀�M��ޙ3n�T�dtHܖ�͒����`s�4��l����*�NQC�K�9�t� �j[su �%ݬ���"5��Nժ�h5�d���%nݲl�jNʇ�Z�ڦ�2TR�(r��
B�����sU �j_9����1 �Y&�e�*s��%Xw6X��%����`}��,�I% w�z\$
�j"�� ���� �sv���m��ӻ������`v��CcB_(:��nI`qww� ;��U�s3@���[��Ydm�R����ʀs��X������3��Ӣ���DhN��}&�Wn�ܻ��&Mխk\y�e��n�7����g�F^V�nm ;��/��@z�L@s��Vw��
�l���������_I�s���`��yDͿ�Y�Q���_I�s���`����,��{C��!)
"�;�.���w�~0����Ri.��؛@�Bj�M�����;6N�uTE[+sv��`���n�=}& =�*@�G��� N1������K�nsh�s��#�bc���Z�F����ڌt`�z�3sD�su��1�qR���q(lhJ��9�X]�w���UU��|��o�_9������nʵn�i�8s}u`s�4�5w6K �we�΍Vh:Q'BN�r��@K�7P��@{�� ��^�%B��#�jB�ՙ�X;�,woL���q$�v�O��fiJ����Mm�o������Vp;mJ������4�I�)�`�� +�+�hҤ��q��z$���u�V��W��G�5u��s�=u�v7 �ⵋW=:�@��	oլf嬢�Fy����oc�/;9Ӥٻu���۪��B�Kmt^&
�a����X�ׯ �*�Im�[۞��HN
�`���8R�U���ijߝ���E���i��Ӯ�:\襱���8|��F3���s�^�s��f��m�ݸ��� �}�t� ;������z���,��=�N���G������MHw�~0mo���7k ��7Km�C�I*��ri`n<��.��ݺ���n�TB@�JMG<sq��1��-������t媞�D�Ɏ�8���]�v��Y��ˠf�~,�͎��
�m��S� �+q��Dx~�(891�#���yθ��n�rGf��O�.�����V�mԃn<|��������ՙ�~�� ;��`f5Kk�)4ؤ�h.�`s��ci�%Tzn�� ;���soL�	6�6��o�����Ut�)���I`�l��T�s�Ł����3q'B�P*r��Xz�.��X�O;�K��~����K�����U��Awwx��� ��|�珀�������5��PĪ24���'*V]<�i"��K�9���F�x��Fu�:��*�D���9�p�͞,Y�%�s�����O*��!TI$&JMGVf����M����`f����ɥ��#���OD�L��R���0N�Հ}��X[M7���ڻ���`^���9�j��wvTM6�A� �{�U}��%)N��w{�'����O�6�ڊo�h�URJV�7��R��}��%)N��w{┥'��wC�JS�{��R�����]�ֺ�����=<t�96�@����Đ�����v�6^��8�����{`���)Jw>����)<���JR�{��┥'�}���JR��fh����l�[���)J>��JR�{��┥'�}���JS�k��\R���j;��R�$�U]�x6���6�┥'�}���JS�k��\R�����h]�&�uT��
�K��R�R���_��)�����R�>}�v<���@����ݘ��5�H��Y!
�jT��>JR��_wz┥'��wC�JS�u���)<��vJR��TO{o��p��u���t0��랪l+Il��p�v��Ϯ:��n���}���bw�z�)I�����������)JC_w��x6������6��}ӻ/�*�"�R���R���mk��zbK������y)J~�����)JO/��'�_͡86�ڋ޲�%T�%+Aus�R�����%)N��w{�� `2On�������k��┥'���V��"�J��Iv'�h?	�V��)I�����R���w��)JO>�h��m��H�`!U�T��Ɣ�'��wC�JS�u���)<��vJR��_wz┥&"!�6�&��D���D��՗E�R��u��B���֝X#BvG�En�;tc�t�\�0�J�a��nU��#,��9���[����ӃId��S�/F��3^|�[�vgf��z4�"__����t�
�c�y����[u��!�0n ��푶`4�ú��݉k�m�9�9`���@�F�ZMĄ��b/76؆�eӫ�+�b"��,�I�:�ǣs¬]>#�-VT�;מq�1�}b���c�^��ٷf���#O{�o{����mo�6��}�։������X��6�����mh�޹UPQU�\����5�{Z'�h[���c_ɇ%(}�ly)J{��~�)JP��#vY �R�.]X��mok�u�R�>}�v<��<�]�qJR�ϻZ'�h_.vE{r]EAE+Ur��JR�Ͼ�ǒ�����)JRy�kD�mkg{�x��5�we�e^dW*UR�u%]����;^���6�$>nׄ�@�����6��|w�I����I��w�<��UB%ջ�*�H�3�-��l�v�c/:;���Y�}�s�QӧL��o;Bv#Ij�R�W8��5�z�	�����n��k��k�6���6����6��w��""�J��Iv'�h��}�w��~C�!���~��JO�������~����)JO>�]���6���7�%"W�!E*Љww�)JOn���������)O�	�8����C�JR����JR�"�T���EJ���mk�V���)I��k��R������(O�d����mh������TUl�.�)JRy���<��? O����\R����hy)Jy��┥/�O�~=u�5=8���%�v��-�W^+4�O[��7<<��{Ӿ8��`�^�M�p�)J}�~�k�R��_}�%)O=�{����ԥ'߿k�Jk�}%����TTT�QR�mh�����R���w��)JO>�]���mrst�m~R6����_�U�Er�T�Qr���mk�_�Lmh����Ex>�J�!/�S��|��7�g8����<6R- H�|'5�F{��&)c��3�����ID�,�@_�9$$@�(��3��!,�1��J�QJ��4���F�(#��C�dG��|)e��p{��G�ʈ� �YT=P6��"/�	�D�+� ]*�" |��¡��G�@z�'D 'ު�"|{)�w�m_ov�����Bݲ蒪�IJ�]\��6�����<@�9��)JRy����R���w��)Jk��j,�E�WH*]�����n�┥'�}ݏ%)O=�{�R��0k����mkѝ^<�\����U��o��7�jR�g�kb/��ڄ糓^��m��]4�{:�Da��Y�n��)<���y)Jy��┥'�}ݯ%)K�{�|R@�v�%�"�]�����mk�u���)>���y)J^���┨�{���m�mmTRDU�\���)>���y)J^�����@IA�{}i���;^���6�>��vY$��Z�]�x6��s���hRy߻��)��s�P�I��ݷ�h_.�mT�����(�vV6�JO;�v<��<�]�qJR��~�׃h\��+@���mU*�%ͧ��r��\�ɲ�WMێa0�ӓ�ձ�v��u�ū���]Er�T�PJ��mk�V��)JO���^JR���)JRy��O�6��m�d���Z���JRy����R��=�mqJR�Ͼ�O�6��n�mh�;�E���J�J��mk���ch@�����R���w��)JO>��^JR��vR*��Z*]YX��Ġ�7ly)J{��~�)JRy����R����X��5��tD����EUՏ%)O=�{�R���ﻵ�)�{��┥'�}ݏ%)HJ0������t��`� ?�~�?Qӱ1�:`��ݦ���6�l�'�iN���){��&ݗv���a�7��g���^[��!�}B\�wnXY����7-��kr�s�M5IQ�oq7a��GYl�-��i���=�f����f�1؊OV�8�^C:�1�56�����X�������Ց]s�ۅ�.��)�m��.�W<����v���c������=���댇g�t6�=An�`��N���7g9���}Y�N.��"�꠪I������6������R��=�mqJR�Ͼ�ǒ�������6�>���$W$"�V�K�o%)Os����)<���y)Jy@���v������6�]JEVT�+@���v�����[��)JO>��^JR���)JR�ΛR��W*J�j�U��h_r�f4�)<���y)J^���┥'�}ݏ�y�%	BP�$BP�%	Bf`�%	BP�	BP�Mk��Ǭ�P�R�J�]����$�(J!(J��30J��(H��(J���(J��=�q��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bg�~�o��(J��J��(L���(J!(J��30J��(O{��8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP���߳��(J��J��(L���(J!(J��30J�۽�w�����/��ygI�p��6Eg��>U&�=�ʓm<k'V��y�8n�1�Y�z+Y����(J��(J��"��(J3�(J��J��(L��߭���%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�{���(J��0J��(H��(J���(J��"��(J߷��y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�{���(J��0J��(H��(J���(J��"��(J;���5���kef��~x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B{����(J��<��T?���(��*^BP�%	BP�%	�`�%	BP�%	BP�'o����(J��(J��(L���(J��(J���(J��;���8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	�}���<��(J��(J���(J��(J��(L��@��&�<OxD��%�]]^&P�%	By�%	BP�%	BP�%	��P�%	BP�%	BP���߳��(J��(J��30J��(J��(J3�(J����ÂP�%	By�%	BP�%	BP�%	��P�%	BP�%	BP��߿[��(J��(J��(L���(J��(J���(J��=�s�P�%	By�%	BP�%	BP�%	��P�%	BP�%	BRk���z�
�"*�.]ϾMh@%	BP�%	Bf`�%	BP���J&B���<����߭�hhA�ﻱ� �	���(J������x%	BP�%	BP�%	��P�%	BP�%	BP�D�&�4	�M&��!R�5���	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	Bg�~�o��(J��(J��30J��(J��(J3�(J�����	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	B{��~�<��(J��(J���(J��(J��(L���(J���	BP�%	�`�%	BP�%	BP�&f	BP�%	BP���&��T_*��r�r�Q% ��O<�ղ�m��0y{F��nݯ7�=ls�)9���kY�ݿ<��(J��(J���(J��(J��(L���(J���8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	����<�J��(J��(J3�(J��(J��30J��(O{��8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	�}���<��(J��(J���(J��(J��(I"h@��&��}U�r+���Qf��(J��<���(J��(J���(J��(J��(O~����P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B{����(J��<���(J��(J���(J��(J��(L��߭���%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP�����(J��<���(J��(J���(J��(J��&���U�V�*U����&�2��(J��(J3�(J��(J��30J��(O{��8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	�}���<��(J��(J���(JL�
ȩ Hآ�
�NBP�	BP�%	��(J��>�����(J��(J��"��(J3�(J��J��(O{�߳��(J��J��(L���(J!(J��30J��(W{�K�,�RJ��*U�Mh@�By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�}���<��(J!(J��30J��(H��(J���(J��=�p��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	B{��~�<��(J!(J��30J��(H��(J���(J��=�q��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bf�&��� ��AWV_�&�4	�L�"��(J3�(J��J��(L���(J���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'�o����(J��"��(J3�(J��J��(L���(J���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�&}�����J��(H��(J���(J��"��(J3�(J���w�� ?M�	Ĉ�3��%A;\`1����U�m�j^��P��]e\�Aa�b^0u����g�P�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	����<�J��(H��(J���(J��"��(J3�(J����ǂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�}���<��(���H��(J��`�%	BP�	BP�%	��P�%	B}���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'�����{֭Xa���k7���(J��"��(J3�(J��J��(L���(J���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�&}�����J��(H��(J���(J��$�����)����8�)K��4���V�K�o�6�st�mJO>��JR�{��8�)I��wk�����6�]JEVR]���o���<@��kޘ��5�{��JPtG�%V��)�/���6���ݪ�����XJ��mO=�{�R���ﻵ�){�{o�Ch���O�6�źE�]"��B�m�mї���Y����]���mFN��c�;u�x�a�⫢�
�D�@]���6���ݶ�R������)JO>��JR�{��ch@�9إj,�D�. �V�����)JRy����R���w��)JO>��^JR�ݬ��k�Y�h*����6���ݴ�mk�V���R�Ͼ�ג����)JRv�7DK�BEv"�������[�D�'�}ݯ%)K�{�|R���ﻴ�mkf�t���(��d��1���}�v���/}�m�JR�Ͼ�ǒ����}��)I���	�0Q4���|�5�Z��Y��[teݮIڃnMh6�B��vV�)��&k^ӣ9q�lrܼx6ۄQ�&H�e7<O��}w�ʝ�N��5�NذL��s�y#+j
��=t+b��m��1�s�z��W	m��^�M�fxNw`f6�k78�nݘF�m@[��I/��^�yݳG]>4w���<��+pmCu˶��՜�]����I�:^ܚ�b����{��s��1��j,�c<%�id)ջ&��E�=v�n��l�����#�<�Gkc�^��o{_�)K�����)JO>��JR�{��┥'�}ݯ%)Oo�wuR\�H�ªK���k��m<��)�߷�┥'���%)K�n���m]�wj��Ep*�n�Zx)Jy��┥'�}ݯ%)K�{���k��m<@����V�pR�*�h
����5�{���m��x�)I��wc�J����~�)J���b��Y�QqJ��mh�;�|R���ﻱ�)��s�R�����x6�������}h��
�]�f�p�݆�����N!;a�v�Kѹ�6�^�y�H)ʪ�"�h.�����kw���R���w��)JO{��)y)������6��'�"\�H+�Y��%)O=�{��pR~A�����^JR��}�|R�����O�6�j7IuP�
U��]�m������R������)��d��z����v�鍠mz�E�"�(��%K�o�6�9�V6��w��JR�{��8�)I�{ݯ%)O�6�]JE+TT�+@����JP��~����)>���ג�����X��5֗AwaTw,)��3�y�A�ɍU����:5�]Z;��ۣ��&��uwWQ\
�Z�Ui������@�'��v���=�����)>����mk�Q�m*�Iv���@�I�{ݯ%)Os�w5�)JO��v<@���zch@�{�Jй$QxV�[^JR�����)JR}�{���T�("h�J{�����)I�����h]�WJ۸�)e�*��j�����c�JS�{��R�����ג��	s����┥'����E.P�؉R�<@���zch@�{��y)J^�����)I���ǒ��՚���kMPF@���i��֩(���w<P'�ل9����mƎ����}�����eU՟6��w����hG7�/�)>����R�����)zp�tE�QUXJ�v��m��I~rR����c�JS߿o��)JW7v������{R]JE+UR����)I���ǒ����}��?����}�[x6��w��x��5�v���+�%R�r����i��w��D�'߿~��R������J��0�x tP>�I�o�JSk���MWUU�.�mh���x6�%������kw޴�mk�m鍠m]���Y!r�Ԫ)����7e3ۃg�8�ۇ�6���I�m�zl���E.˒IQqJ��mh��e�JR��ݏ%)O=��p?*��-]��m����T�^��"�\Eɭ渥)I���Ǒ������>����)JRw���k�JS����qO�1Jkǉ��(R
�D�v��ms��R�����גʢ��g���qh@��i����F�%��mkz��)�R��߿my)J}���5�)JO��v<���Q%����m~�Ǣ,"���T���iJ{����)JR}�{��)��s�R������R���Ԗ@�P����|�*M��D��~ 	�� �8/6R6<��" �|E�M�`�	�H��oA�J�0B�ؠ�頒H&`��ij!	�*A����'|� t�� ~����6� �ϒ�ԒCD�R�D�L�!�4xI2h5��L|HC���R�4���	�@D`�8�,�66��xr�Y�f������N�I66��v�YC9u���kMCZn뫮E+�R3�tjm*[!���ώ4lK�d���\��l.�p�6�5SNHsXK�S[UK8Ŭ�R���]*�mU*�I4Ƈj�Z��T���fe�邪�$%�W{<�p�M��h	Tr����@t�iC��ڠ.�2�%x�ՃȽm�`���;6��ܼ͍T�DX�� t���;#P���v�r걌a����<r��ʛ]1yb5̤:�^�Xp�R_Z�˰�L�T�qb���g�ل�ח�G=ls��	�1�����`)y!�.�:��.�ṷC�!ȸ+���m���+��bgS�Ǉ�p�ܙ{ykiy�܂x�[���yY��U��\��àUcL]p�<�<�4%���Gn��c�.2�T�4�BLi�1���Eр�ͱ )�n�u�8���x�x�ρ)֋P����9�+��Bn��Yuf�����-Rn�ܮ��^��٩�3&Irn�qٝ�cgE���oV북��(�\Xȯ�)�`�49���+Z�1��mѰ=+��s���WF��`�Ξe��ܻm�Y��tЖy��KbŶ�9��w;�-���:�c��)3����\i�[o�1�R��u�Յ�DΆxʯm���g$WW�RPgts;�4�Zz�9�Y��tjC��`�j[�|c)òj��r����ۜs���6�\��C��OhAC�v�U�D ��(^�㍃��[����yMfl��z�)e���:ݗ�(غe��g���E7�6��<�+Yr�T�'�����@�ꊳv	L�vӸIڔ�
/7QoV�a�Ib���M�]�cj6�J�� ���D�g;;ml�Oj�eP1�����힌��Ӎ�m������K��6�uҫ��]�EV�⮕y����T����Z�J���PWR�ݻf�\Ke��g���Q.�J�qB�K��ē�6�>4(T`_�S���E�:u+i'�Nh�㈗D�j˻��Q�#�Dڙ�Q��=���.�@���$��fW�:�q�Ncrٖ��rm��N��q�wZ�`�ٶ͓h[�ֱs��[qnSt�ݹa7O=�E&둛���LY�w p;g۠��<�����#�nP����+b�K��Ǹ�v��ݣ�� ���N�l\�.����@x�vY�Z�F��gg �gN�F��X��==;��X3����K���mX��;m��\u6y����{�޹�|��g�s;�uJR��߿ly)Jy��┥'��v?� �JS���ٮ)JRoC}WחJ%R�wWv��h\�{��)=�{��)�w�渥)C�wm<��I$'�{S�O+�UU�us@���z����M����)C���ǒ����}��)I���5�!$�(���[x6�ɦ�S��M�JR����c�JS�{��R��#L�]��m����T�^��"�\A���|R�����c�JS�{��R�\��o�6�ov^6��	�&�E?c�:�=d��5tx�J�.��[�>�qŚ��m�#�u��{��/�b���l-����~��R������R����mh�wm<@�;��	taf������R��}��y>(x��O���������(w��<@���zck�H��'�DXEU�����mh����O��i��)�߷�┥'{��ג����b��%�
V������6�>n�%)O=��qJR��ݯ%(?3s��K��6���=�����Q*�*�[���JS߿o��)J?�{�߶�JR�߻�7�)J{��y)J{�Lr݉/U=�y���l;9�s͓����mՋ����voGK��C� B�l����)I���ג���w|R�������������w��1��k����!fU���Z�ג���w|�g%>�޴�mk�����6����_��[�m��\p�+����hT=���ǒ����}��0�����%03�I�wݯ�6�s�x��5ä�.Q	؂U]��h??�5����@�����%)K�~���)C�{ݏ%)K�MЗAJ)*�*]�mh���y)@~������({���%)O=�ٍ�m|8�hˢՑJ,-ErN
�]wNt@Tv�24�V�q����Ob�E�UXK�v��m�v�����y)Jy��┥'��v����b���H����*�@���{��)��s�R��w���R�G9ݼm~M&�m\�ޫ��ˋ%��v����������qJR����^H d�����)JP����JCk����K$�U%���6��ww�^JR�����JR����JPq°�P<D^ �}�_�g��k��
ې$�\B�V��m���R�?w���R���w��)Hk��m��גI?S:�yU˺��Vqg�S�]y�T�mt�8����K�]�N�Ä�Qj��0#�]]�͠m{�z���)��s�R��w���R����m\:M�%�
A]�%U�x6�O=�{��*������ג$��������O}�Zx6��wI��)E%[%K���m]��o�4�=��┥��v<��<�]�qJmz�M6"���%˻o�6�=��┥��v<��<�]�qJ�D�����ms�د�#�J��
+5�qJR��w�JR�{��8�)I߻ݯ%)Os߻�)JRB�?(��ChiS}�Z(��J���i@8�B�ܮ[gqOQ��vw�q'6;��6!�6*P��9l�����v���Y��9"�k���2�#{j�����m�Y7t3�$�D�:��6�!�$���f�=#���������lu:g��5���&E�Wrp�zy{l��xh ��d�v���4R95!Ld�4��䛚�! �=b���ջ���s�D�|�\�>�l��p� /C7V����ӳձ�v�e�jؚ��G�r��&�o{e)O����)JRw��k�JS������.JP����JR�}���R�**Uv���mh���x/�FC%>ϻ�\R����߶<��>��ck�I����(W�@�	e�T�my)J}�w���)C߻ݏ$!F��ݴ����m������J�M/"0~����c�JS߿~��)=�v����Nwk@��dT)#{��k{JR�{��R�~AI�������gwՍ�m}��h��n�������p��g�$��Xwn ����Ͷ��n�V���6����յ;<p7����)I�{ݯ%)Os߻�)JP��{��PO��e)O����)JR�ZO��$"���]�x6�����cD��)C߻ݏ%)O=��8�)I߻ݯ$�_�Dpu)���7���-Ғ��EJ���6�?�����������)JN���y)Jy���qJR���mK�������*VUݧ���4������8�)I���my)J^{�w��	�wm<@��*i�R�P�UXV���R������R�� �����┥�����)�w��)????�MO5�,Eӓ��8�&�a�;elO�wi�m�M�N�6s����6��5��)y����({�{��)�w��
˒�����ג��x�U�B�Auwx��'�ݴ�l�<���┥'~�v���/=���₏��JP�����V��t���k{JR�w��)JRw��k�_�� ��K�<���)C�~�ǒ��;��	t������ch�m�(5����@�9���h@��v������ō�mz&�d�UWYk{��R�����R�~UB���c�)���ÊR������R��3�;h�5��}>`���O/S�7��YS�[��F�k��O[�d8�������	�v���ŀowqy$����K��������۫�PrN��b���r�{ s������m���mU�?����R��
�X�~�� =�j �M@{�T��IV-۰�uq%Z��I'';�� ��׀}����<!=UÂ)������t��0�b���>�ݬͤ��gޯ�R �9��ѵ�{WF�+rZ�	��҄i�.�A�KқJޯB9�AD�����"B�����sn��m����y���'�Հ�{�.��y���ݤ� =|� =q�@{�U��m��4Ӫ�~?DY$�U�*�� �}��\s�_���R9�pGKڑK��*�u���Ҝ�o� �>T�|����U_c�b�K���nT�T�����u������_ɶ�����;7߫ �ov�ɤ�cmi�sV��VJ���v+
�pV*��{@� �t`�gg��\��-m��}�r���]��n�ӽ;m�u&v"^2J��[E��z�r��p����t	�u���{<�:�99{]a�S�٥����G�^(�"�oW3v�����ѫ	�Y���%	�C/m�q���[N��[�x�x�(�r��!Y؍7f4<x��̏pF�����%�盳%o~��}�|t%�m9s�9�n������n[��eSu�="���7��-$H�i�� �V��]X]�v&�k�i/�s��X��(e� ����*���v��i$����� �wذ��,��NC|��S�2AK�.���ڀ�8����s�n~73?eY�P^f���r*@z��A�R{}��G��RGV�uv��T�=�j �M@{�T�wҰ��I��5n0.u�ǋu\�6d5��nS����m�3�`���w{�q��㵃��m��9������H	�`����{R)r�%XUIWx���i[Ld$eFS���W�_w��X�o� }����jC�6x����d�۫��$���u`nl�����#����������=�$ӡ�$�soL �������4��i�w߸��ߩ �H�8��9V�����I9����9��,{������=j���Zf_dv�j��1���zh���e�Ǜ�cm��W�կɴ�j��e��K���Wu�����s��͂��b r����e0D�nK�ͺ���ꪪl����`b�~v��,��t��>T�>rU��{�ܫ������ʇ	!^ TDAR�m�D�C�'�އ��2���jSzѢ؆�"b8X�z�����A A�i�qsb@��p�4
mR0���H�	� e��Ҟ�`*h<�d�u���@�0A4�N��A<P �Ux �Q�����.}��_}�x�z@�b,����uf�m�Wg؀>��@{�T��6�l˺�TU�*� 7���?6���k��ܮ��OŁ���`ni��le�*G.�����~{Pprcr�m���I�0��'n�;`��Y$���n����f��Ձ�٥�����_U}\@{}�`g�:^�M0��ݤs`���#�P��4�rＨ˲"AWr]�'g؀#�P� #��]�&��	uqU��y�����^��`��+}W6H�C�ڦ�}V��e�Wt��M�@�
�9�H	�`�=�j ��@�W�ߪ}�����d8ӝw�23��n��dX���h���c'I�zT��QqZ��6��,��C�
�^f�p����sPnj��� i�$�UXB���>���y�һ��P�ʐ�T���Lٗu{��U\(�WX�ݼ�wqa��jOo��`uf��Y����q��ӫ��$�&�S���,��b�>����i�'�ޖ/k�� I�JIV��Ձ����w}_ {}��>�w��[bIw��o��)���]��'n��:r�{)v]��A ��(��h8[ZH��n;kd<�&�e� �e{�{:@z������9Q�\��{O�s�+��=��b�i��:ܒ��l��h&EN�ktf-��	�e9��Z%���+��⍆�1j�gײq�ս���F�E���i�92��J��ݥ��lܺ���\\܄g��佑�ke��?}ݻ�޷��� ,�$�Í��p݄�q�fqշn��=9m:x����M�#����$�r
��#�����j�~v���s��ȩ �s	�Yv^��y��95�qR9 s���~M�I�Tߏ~d�R"b	Uw�w}�R9#���[�b �}��
p�7q�*�*����s��|�N� 7����sn�z �U$�)C�U���1�UW꿧�o��>T��EH�Eb�B[)c%/��I�:�6���]B�Q;���ɦ�x�ml�㩳�ώ�!Ļ2�q G&�=�*@G"��sPY�����pm4���8s}u}�����@`N�ߗ�?~�ʮ����77e�ո��$ۡ�@9*��EH������ϧ�j��R�m2� �8��9V�Iw7��=���s���M�=����z�P�D����%�nn��W���+�{}<X;�,�4B�*�D�IQ}C��wh�@��tb��#��޲�������
�]�����8�� s�����@=�����x.��*�*���l��@ɨs�����U]��A�ʈ�J���$� �o��nn�2��.�۫sf�~�a5�J6���U��NOo�x;�ŀov����U�]���=[��Q�]�6�ut���|�� s��#�P���S�>���vZ����\�Paێ�P�pi�FTe������� �ގ�����ww�3��6{5�lݦ���o� s��#�P� :m"l �:�����s���UI�}x;�ŀo6���I�o�'��
	
8��X�},w6���I{=<Xs},�L��H��NI`s��X�oL �����x��M.&Đ�J�ǂ	��߹������޴��eU]�y�� ���w���}x����?6����P+�E�"���K��K�g�9��V�O�%K��n6�Y]t�6�v���Bp�s},s6X�m׾��~I�P~����5hx��"�����J�@��s���� {���~���l�{�F��i
�66��~��3�ܖ������Z���t7 &� 'M� �9�75�ꪫ�>� ;�}<�*'Q���w6X�m�s�� �n��)$�!�v�@k��=���N�m��ݍ;u�K\�O��41n-�u�#(���v8�nqn�`�f�b��x�l�DJD��َ�Q��n+dӫ���M�5�[c��ܕ�n|����l\��\WU��چ��َ�OGR����Ԙs���d��[���Oc(��[f�;`d�V[�N[�[��]Z㉽Y���F�t� ��4�3�������:�D��,0�۫�\nҧ%ɯ/���汰��Lv��]=�z��Q��R�����& {7���sU 'H� {��RT�^f]�w�P^����� s��#sWԒj@[���B�R��Uv�w�ŀs�x&�JC۾���b����AJ�B��`y��&�J�{�Հ���P� 'H���͆]m�Qu��y��#sP� 'H���2���W�K~n�I"O�PSg�2pK� /D.���=�{[L^��mۮ�t�[_����_n�o�p�c��LnL}�������X]�v��,��ը�$ӡ�@I*��n��.��m�M���fg� =���>�mՁ��D�!**'Q�r�.�:M@{�T���H	a&��T����I����u_����;��� ��HU�=��)�@/3.˻�(%U��;��ͤ�_�I$�{�~8V����
��Y�F�i(�LۋLd��p-i\�98,v��zϫЂt�-ZQ�%E9𣒬̚X]�v�ݖ;�u`�/�@��I�!����g�m4�w޼��b�7��0WC"��D�*�!$���9��9|�i_�Q���I�C���@@�����E_}����r��{�73J���p�ت����w7�H����1 N�P}p�f��eR%������6�o�$�}����߽�X�mՁ��M��V�t7
v��<�,��n)�2:)@�#�OS�n�^�ֹc�����HX]�v��v9���i����y@����)e��7q.9�s��=���b���i�|{�%T�E.�T�u�s��X�oL?$�JN�� ����n��Q� >rU���K����չ��(�M	���������W�V�	�8�`w�5X�l@{�T����!X����*��Ev�	��cS�V.^����[Q�:m���x��ǘ&�j�N�RD�N+ �͖;�u�n���I4�����`[�]_�Պ�]6G' ����W ��x�8���w�y��m%!�ؽ�%�*��.�v���*@z��@9�s��:�v�H�r��.J������w}X�o� ���X�m�����`P=�=A#��i���$sP� $qR��w\�*�W$ v ���� D�H�K!��hD�ʸ�E6@8��W�
bǻ%)�P%p���/����B�g��lI$��l��@:0X��İ^���$�GOΞ�Ξ��� �Nt��m���k:ۺ���;vee�cL�.��z�	��ѕ�'8{ٍ�.��aЮ0�wC�⪕����ۣ�6!q�f��Y�GbV�v��V�j���Q�k���V��eA�;3.�UU( ����\�p9p�j�� r�v�]][M����`����;eRɴ���YԻr�ۀ9�ԥ�d�MTkn��v���xm�G;]-�7��vv�y�d�A��G>t��\��%XŁ��c`z�:���k2�s���v)Wn0�ٲ��F�q��κ
c�=�2��	���)u����A.��{E�eNd;.kGO	��3>��<gmh-/lu�'Tds�, Y#�wd򉽻\���L����V[t4� ��J�ev�p.fUڷvr�sI��v�mI-4��oo9�;�m��[����V9�ʼXpt@����
��\cvN�Jm����Wd�ݶ�ٮc�d��'�`�U�P{W�:ѹ�@�5m�(ꓴ�4�\��L�N�qΔ�:�3rZ�d�{p �^�"���J�c�D�=�������d�f��rp-��˰��+�̮��d���"ùz��-����$��{ܚ�i��a� �\���k�Bp�6x���v�rng�G�\����^�y�0��UQ���.�W)(t\�#ʛ���2Z^2�\�]֌V���	���u\֐�2mn�+�0�z�=��2����X�+v�j�u�؁V�nK8�zB9Q�u�K 9jt'��ۨg����L�&v9�O��6�W��r\��SF3hܫͲ��n�V4t���e�[h���A A��<��f�!gR�l7g)XS� ��cvY�ŶR�ۭ�%t�l�V�	�G;{=��.^�*'l�ٖV�]���q�*��1f}�����y�՘�آ�G'E��u��S�L��f�U����]kjk6��=�J��m���5U��t�[(��WV���)���v�ߝ��M/6��b� �f ���Q�Pq������w�p֮LkY}���Nv,��r���&ʜ�tH�E�C/q�@�ٰ���څm�R��m�Z�q
g����n�x���z�$E�f�v�Ӻ�q7�M���Ncm��r�7=���.�힂���,��+��G�;Z�紪k�mV%3��p��w)���qd�%�`�>�^�a�D�c>��nء�Åh�÷lj�ꎶ�a"�߯{������|ֹ/<V��@2��!�Jۮm���GC<����#��nl��v�Pe��� $qR��g߿SM?����o�x�t�!U�]]�G s��$sP�/�U~����=�Q[�"HT�9%Xs},{&�=�*@F�~�{r�6��wd�U���JOw޼���o{��)~�����������jO�!Q�UӦ)���~�� s�P�5 �@������]뵲�zڱ�Ng��ӚԦ��;Hvl��f�Y����������-���hWwg�{wذ�ݼ �n��m4�������m"?R��u) �n�ki.4�$�T[��s�z`�ޙ�$����Q�	��c��� �}�@s�o`�9ɨ˹�r��J��@s�o`�9ɨ>��R{����AO�r�B�r��bI-̽/�$���i$��vs�%�f�`c��ww��?����I�VMX�=���_^Aْ�ާZ��-4t��;v�N��:���w�Hv�	I �8��I#���-$����q$�������K۷�I#�E�2$�TQ	'#��K{�9ĒųZ��[�zs�$cݎ�W�M���⸧��
m����]�9$����XI&����H4��ؚIbIJ���/	$���Ϥ���Km@mҒ��Aؗ�W��w�/�$��묒I7����O4�ɫ����Y$�z�o�!**'Q���Icݎ�I-�l�K�������$�kI+i��e�2����]�1���kY�u�Z�t��yu��]a��R�U:v�`�)R��I#�I%��Nq$�l��I.n^��I,{��I%���%!@ܓ�I,[4v�K���8�K�v�Igsg9����/�
�]��ued�N{}���$��۬��I7M����KW��i$��TV�D%E75$�q$�=��$����q$�=��)�I�m���+��/��Ahz�E�@�(����I%�ݜ�Ib{��I.�o+�I%�v;I%��54�����}�9�������N&^	���	��n97\���C�)�\�ت���1$�����I.�o+�I%�v;I$����I,x��8�6�'��;I%���s����K_���[�z��I;+vVy4۪�;�P��\uNW8�K_���Y���/UW�WͽO�N�Ig�ܮq$��M-�RI R9$v��osޜ�Ij~�v�K����Icݎ�I,6�A(�E%!A$��I,Ou;I%꯫��v�ԒZ���$����<����T $RPu��gu�S�:�Wo5ضu��[l���]u�e`LV�a�{v�}�b�v�l]�ۓm����8ؕZ��_����A؎�6a愶�x��5�8�����[���<���N�X琶�������Y�[��r�nun���;V�ہ1���u/[�TԹ{5� lf!=t�$p�խ�	/m�h������ua!�{U�z�X�:^����RD�{�WvL��w�9�ָ�Sum\H=���i�l�v��]���<�Zآ�
"R'�$��{��$�ǻ��Y���$�'����[�Q��!*)�	�ݤ�Ih�5�$��������8�4*�!$���`uf�=$T��Z�
W�-��3�eay��Ͼ�����K@����Eӈi���$v7v���Y�ޟ n� ���`m�[��E���#n=���q[�q�=�8K�G5vS�����z:^��)���i�t9\5���3������`ssn�a����$����w0���F�ԓhM$�Qٹ��z8��$�Hy���A����& =T��Z |�%]M�&�HQ���۫��U�gse�ՙ��+t���!*)�	�% <�K@���� =$T�!Gn�������@u��q�L����+০�W[�kg�M�n|Y�c�ƈ�0��Pm�@9"��Ih�*��rT�2I8-�;7v���ri`����f�-��4�S�V��ŀs��0ŉ�I$$�U���`b��`n��{H)|Ө�"r����j��b� ��f�]��ٺP^��P��H�������JJ���(��͔:[�����d�eƯf9r�Q�ܵ��t������h���(2�w�u����*@w=� �ݖR���â�
"�;7wqz��׋ �{׀}9��&�r���IQM�MI*���<Xf�8�5��۫ ��f��B	F���M%�U{߿^��߫ �����&�ʧȐ# �`�
�4b�Q��bM�rU�w��%�eڲQY�]a���:��b����� 6��ʹ��}�Uw)\�v�$IJ�Z1��c��;;� �#k�n8��.dE�@��qYT�-7�WH�,ڦ�
jG�o���Ձ�ɥ�ff��s]��߈��R��Q�D�Xܐ@��\s�*_U~��B��A!	
B�7w�����`swn��M,kV��Q�BD�rK��������_���jU��7��B�������XܚX{ݼ������sFj��GJ�']j�0���ȥ��l���JGh�������$H�;lc�:��z9��[!���t�m�k���-i���ͮ	3�&Z�&�4���5G @R�W�X�м*����ag�Sv�D�7�.y�6���k�n^no�����»�
�M��N���vz{f�B�/Ԧ�:]"�ݧ�Ft�6��λ=���hٜ�����=u�=�rPݛXK��J�3�#����m�[����Փ
k�x���c�.jI]�饀ff��s_ﾪ���޺����I�RhA H�,1�@z㘀��R�� 9tf{j�eH�EU��r{ެ��Ň�i��������?�{��9��WN M�i����@zH�ݒZ nM@u�����V�T� �V�r�f�4�_�I���~��~���� �vjFu��U�3���&��e7U���)#�1v�%��N�Ɣ(TH|���3$�_I��*@wd��%K�+oq��r�� ���`ڍ�_4���&�!���ʃ��{�,��z`N�k?4�RQ{��e!b.U�`��,�V��ɤ����`�|��JZj�P���&��a��UU�_�րw��؀�nb��H����pC�R�N+�3]�ՙ���f�XǺ���iRLRD�u;n{�.%x݃��!��zLh�R���g^�!�g��{�Tv�o����t1�@��~v35R�$�����e
�l�ٙ�Y����qR�$������/������.W���W\�X6��y�}�r���GP!�A���I��hN���\�cAbX��dX�e�q���ǜ-�Fe�!	�XؐDᵷ&�vf�����sXc6�xq�; �DT��J�C�e���0H3ݚ5&��L���I��F	�<��!��0p�G��p�@7D�M���X��D�1�c�2Kz&e$B!���bd!�eA����M0)0�+1�L�|���$��|C�$5��$��,�Nڇ	s���^h�a�*A���=���w�<d'8�� a��@eiB�,d���RR���BbXYI��`�����  ��I������ 1��'�	�+�*|�z����)��(z O��lI_Si�{���`owΝڊ
�*$>RE`qfk�:�5��۬6��߽0�'�T���.�m�@y���Z�������������Iċ��C���F�;�9ۀ8k�qٝ���<6C�ǫЂt�:���v�[�7u���,����>��גo�I�Pl��; �~)~�JJ�njIV1������ <�T�����^fn^ �@�8�,�vVf�=�UR]��Ձ�~��Y�*M�rA2�i���M'6�߫ ��`r�f6�J}]�vwuա�6�SR;��u`y/��}���p�{�`�����eS+��G
�X�ܜ�G3����x7<��$v�L]p;u���Gb�frN����.w�O����� :��@y�� ��l��QK�˻�ӽ��ɯ�6�Q�}����]X��W��x^�Ҋ�$(����v�؀�qRݒZ���Qn�]R��.�����m�n��q��Z �sP|� 
p��(�*�24�RJ�wvX��wwӀb��9�w�*�
	�4�QGP��2 g@�t�'uw4�[�Ʊh^@6��h��8+q����s���6H�t��lK�lQ(�؞��탳��-s�5���iǣ�E��ɻwD�:oL������5�&z��9��m�|���z��c�Sy�۷n� ��I{f��η8��롯l,�x8�&-�dCg�şnq�������*g�z�X�=L�r%�Ͷ!���e:��`*�6��;��Y�.��0�C�ݤ8f�j]�-��3��Aź�b����.�M�����@������Ws]��ͺ�������Kp��'�rA1X6���;s�@y�� {����:I��Ȁo��
jG`s3n��ݖ~���;��`b��3�=��#��"r��&�=m�@u��qR�����		$�8�5����2o� �ﮬ�ݖsu��ƥ1Ԕ���KNn�c��t�k�{GYG'X/.��<��bbN	(��R��'#�;ך�fmՀs������`m*��&�P�"��y����(G���s��������;ך��JZD��7*J�wk >���N�k��iI���`��,����T���(��\��ɿ�W�'؀v�؀�{�P�2���lCLVi��1f���۫ �we�ř��9�/��H9$i'�vwi�N����x��b��띮-.ˍ���I,�������V�Ct��TR>��]X;�xӽ��M4�����`ݲ�`�%�\�X�7o<�i$�97}XgwՀ}��,��I)�B�r�"B�V]��������é�m$��ir��ɥ�w���7R�Ԕ(�R��o7q�[�>�I��&�=m�@m*�ؓT�H� ���̚X�M7�߽>�wՀs�ݘ��K��:��@�Z�;]E�cn-��:��ދ�ʹ�u�ܒK']���<�k�ێY&߬���nb���� =����tR�$�8�5�ꪪ��ǾVwg��{��Λ����lCLVi��1f��̚Y���w����;�ٴ�pD�U+u.��6��m���� ���� �w�X�T�LI$1�.jM�b @�*��q�\I��i�r�+ �;d+U����R:�U����wπb��9�4�3�Ͷ�ܡ�#�&Su��n��ļ��tv�,��[���9bOC���s��ww�D�}!u:R9"�[�vWs]��ɥ�ν�`un��
*)!HQ��]���� =�%�=m�@J��m�]]
�E˻�����>�n�?4���t�{ߝ��}���4�P:)Sq�ڙ�ݒZ���_9�7�@z�nS�Ӎ�)T�qXY��WՏ7��ݿܭـ?�$6��!7!U�(�yM�TRJTS*8���Ņà�ɰi�v ��&��D!뒌�3W&뵜��5�����I�+�|�:t�6�f竝�v[�ۡ�Bҡ����ݕ�۞����2���z� R,�v���[]�]��u��lf��4�no,s�ѻm�%l�unե�A�_k ͺ�74�;q��k�N0g��3؉gu�]����&+f���B].����7a��y�s�m�}s���_����|X�7C8�����6c�v�u�U�����5��#��r3��O�������|xy�ր��1 ܹ��Ͳ�i7S�v3&���T��~�:�|���ą܂�
T��tHX���� :��@y������:
�>�E`qfk�:���fM,=K�=�`b��~B��$�(����so`��d����1 93
-?2�t�Nۯ/u��Z���7E��Ƨ�j;y��@q*��t��e*�I��ɥ�ν�`qfk�q,�;QG��J�QR����]Y�}�ݙ��M�J��ͼn���K����	��)T�ʹ��:��G�W}&� 9��Z:n��rq��"����UR׾��ɿvIh��@7.e+3l�̫̭����7�@{�K@rj���0�T+S
��R��_bPIH�{y#��:Z�:��V�n���z��＿|���q���ot��� yɨ��=^�琀gL	�"t�H|��9�p.gk ��z`�ݬ�N@������؂����� �{za�I�Lci0P��_D>9�g��U��l�6�n�)P/�(�Ȭ�M,�7k >���~I��$�w=�`�_�_�Sb�MƓj8X��V�ݖWs]��ͺ�:*+4�2�C����v�̡v0�	��^�����wl����l�s��&�LR��9�����k�;��Vw]��7]98�M�-��RN���g�ې��`��� >����R�^t]8�M�n��H���Ձ���`��`uw5����#q�\�X�iNW}��o�x';��i��$";=GB�>��|r��}[�[�a�����n� 95��b���]�v��,A��A$mIUM%��{�9�yK��rd�Ԩ:Ag'm�v[��x���4�������1��H_I��UU�wޖ�W��& �I��ȩ��- y���s�$�WX�N��&Ԓ�u� �f�=_}T�,�����]X_wF���*pN$��:�L@y��ݒZ�&W󓍔�2������v36����w�ʯ>���^���R�U4�x��c.8a�I����e�I32p$`���Ā �'1l1�#0l��1��31���
1l,��G�=S䴎�x���)�:C[M��H�� ��
���T� ��d�Ba$�#6��& �	 �%)%1�"l8��lڸ�0���I! �L0�%�Bȋg$�J0a�$���"��IS,���Y���"`b��2d�E���Q����_���ޝ=�~w�I N���*m�:o[�K�[�lN:�Mڡ��]s�b��=�u�9˳�:Gm�n��q���إۀ[��V�vl�`H:Ll�ʪ�â��mT����2�ҩ��U�ڪU��@�k��z���^ݙ�g������+p�2 Y9��Z�h�T�Uy��.�U���UmP.ۃ�(�J��(���[w��R����j�4kn��eoc����y훴�^U�-$��I�i�����F��"�pm����*���r�;^9sh�����(=�v�Ե�Z��Vg����ۅ �ɪ�8�%�ˍ���⭪�e֑��Z���r(7����:�8���ێF�=������[s�W8@
�rq�� �+�s�:�eV}�����V��ֵW�g8�]��W7X��o+��h��7eG�n�;Z��m�vv���f��y6����z²oC�I�g�8;��6��]m2���P;rq� [V�`�b[%7�r��kn��w�5�!��V��4=�9,s�<t�zk���s���G!����8%ݦ���mŞf�ίn:��fa�m��;͚Klew1ն�܏-	M�{G:�Dؗy��v��x"���������4==iH�jlqջ@9�%ts�7V3\vy�N 0�5c:��>b�@�k�l�i�y��� �Zv������&bT6�h�Ռ�J��&pL�ۧҠ���EٜnF���d���������pG8re)m�g����5ٶ/�ﾦ��,�:��;E���뱞N�k�z�c<j�3U[)dm�����h&-׵��\�0�Ѱ�knu(j��I�܃t�� ��t�×4KP�0�<k
�6�����C��v�,�=���,�T��j:[��ll$N�`)N>��O\�!Z�2�uUr�0W6H�h2m�m�}��}�p��0�7Z�U��s�D��ѻ[K�+UA�  fƛcn6m�=k�V�än��~�{����A ���PS�T�� �@~"x@UH��nߟf9�u��vzͭ�N�.Ō�f�e`�*aM�T����H����������#^ �Z����rHrEn�Ix��N�C��ύx=�˸���	��[ƽ7#�<����ݏb-uf�'@���d['BDkv�#�s�۫b�k�Fp��9��ԣ�����fx��6.6�u%�c<���e�����\]t��1]�^B�nL����{��y��]ْ�n���\�����v_NV��\-'~��Wۉ�n���/[_�}U�ێ��I�M�dr?�f��u`w�K@nj����u������ܠ�ͤvIh�M@u������I7!��K�.��.�ww0���_I��*��U�I�y�ր#&d�GCR�,����u`uwv�?$�rs}��<���rT�wb.]]`�w���k��|��� ���f�w�~~������/;T�ֹ���<��:(6�F;wz�aMu��Sqˎy�^e�� :�L@rj���7 94�کjFEVJ����y�i$ji/�6Һ6fz���������n��'1�e�JI�5o����dT���1 y���e
�l�̫��dr;着����r�Y�; �f��s]��ȕ=�P��wq y���� <�T���r�Y��+�\���玖獲��K�m��K\r&.۠k�Q�T��D��D��H���,M���{���k�;�V {I��.�IHPG$�:�����H�ﮬ����s7e���wbM"�!DRG`w�Õy�����&�� ��*(ډ!&�j&��Ϸ+ ���`��M��7M�%X~��u��Y�4_9��*@ķ�2���u�J��;9�X��Q1.���;��,������֓HU#�T��:��q+��^��s`�����S��k�ݺ�n!�e�����st�t?���Y�vw6�����1wu��Z+�I�M�dn;��k?4�r��� ��z�N�k ���U�(HDM@"��,�v.��������X�T��"c��!�r;$�������V��q`ci&�ɤ��u�v���7CR%$vVd�����& 󘀕 \U��F��on;��|;-�qٝ�=�������� �ԥJ��&�B
��'#�9��V�Ɉ|� :ۘ�s
������+3p˽ݤ�Ɉ|� :��@z9u�a�ͩI|R���`j��99ݬ?6�rs��X'}��>�f����Lm���8�,�;��u`qwu�����-ӈ��&�27�����>�ݬ����99ݬ�n�M��!�9��V����*캠,Nv��NK����%�nCM� yHez��ڼ��O���/N ����x�r��c��Dl����<q�I�u��]����Z��/���'ltݖ��9�y���`�0]��Ex�xná�^v����v��Ƭ��7�T��:��uc>���9�l��k���P�uhƩ$o)K:��$�$U�.�$�t�f?]�ww���}��OUc�m�ܡ�z6#�ݦ�,��7[Û�	K-I���mg���cb��]��.}1 ��_9��*@>wW��
�����]�vWs]��ͺ�8����Ki���	G���b������L@J��m��IQRE$vw6�����1wu�,y�v��Zz�F*t�cJIV�����|� :8�-�~,X��emۧlGf8ؙ6�76��ɹ.�O]Wv��:����=����?`w�b���G =}& <������EU
`S�w_���f6�M��^���Rܟb�I��p�Y�U�U�ha����*@z�L@;�1�ٮ���*{LGI�RU��u����b����*@y���n�EٺPn���I��� :8�囮��խ\N9HL������jٮ�`82�!Ѕ��#��8c�=�^�s��q:�\�R$�vVf���u`qf��q����U$~�_�~�4�H�B�����ߕ <�K@rj����U�%]UR��*K�Xܭـwv���|I � �	��'�����皰7�� ��c�Ԥ�)S��qX����1��HvIh7p�/w�Lm����JI�1f���۫�{��9����`��r�$��M�(Ge�LF�r�Ti�t�W(��^ʛk�{2�r�}��ß��!�m���|7}u`s�uX3vX]�vfS�`�A7 jJ�;�K@rj���7 =ίe
���+ �n�����%����;��V൒�lt��nK���w}Xw}� ���0-��I�~�dp�H�Iġ+4�JRD0QL4A4Ȕ0�A����~���|��v$�)|�B�����f�X��Vwk ��v�&�Inߩ׊,	a*]ɯGN����e�� Ў�%�Ӣ���.��&���^r)(JTؘ7ҒW �?yXX� :��@y�� W�L�ڻ�U�he�m�=m�@u��qRݒZ��O�'&�)�ӡ� ś�`wT��d����1 �.X�6�/�Э��@sqRݒZ���_9��"��ĩ(�p���{�����`�����q`���4�hI#����x���,\��:.}�"���U��������q�8�$`7,����"=t���&������`�ݡ|�ɺN�H�a�Sl��L�^�vEN�]2u�ک�) ���R� ^��+�n�]�{��ޝ�{=��C��e�����<��Z�=&��×�vō�!��P,0��'�z�r�J�,���U�;&ԕδU.�IWr��W�ߒm%I7�����vaFZwa�����rkK�Ģ�[�=�]�i�R�H���^ۭ��&�$����:��@sqRݒZњBI8P6�:����ԑ����;��V�ݖҭǩ� A!DNG`sqRݒZ���_9�	0��j���WEIwkͷ9���ɻ��99ݬ4����� OM�UK�qEZw�h[s|� <�T��d��u��5�:FPB!T��J����SFku�t�;s=�u�ݸ����dw���7:�cN< �~p�f:��Z�q����hqn�u*'��ɥ��RD��
mPع{��uʽϾ�W������=e%ID۩BRU���ր��1��b��Hs��W�u�Wvn����<��_9�7 <���n5��rK����������&`�C�ն������Gc2�t^��va-���v�ZݙU)��IQ&���9��ͺ�8�L@nj����U�%]f�y�]�����b �sP|� <�U�� >���T�GUaD�� ��
�>���ݠn��<Y���a���: ��	F�� ��F&��5��fx��mGr���kc�z�SK�ꮵ� ��pM0� � %�{�t�H���J�ѷF���>!�6e��K��H�GtЧ�h8� �{����`)�kȈ��a1�$N,ĸ �x)�c�fIQ`A�2�,$� `WjF�zD�@�͋)�Y��Bd�~emB�@C.����0�ɂ:&�d���kd�����q �~`M�,��0"�i��/m���*|)�"0�|�.��� <@ChpEvB���O��@:	��A�ʹ�̕�ŀ����٧�w�)R��]6����}UUK_�~vw}u`��`��`niKlBCp)����ŀ6�����7}x'7k �v(B߃�Z��({b�N�;	���Ô�ޝoP;��۵z:^�x-��bU�������P�����3��zä�R��Ϫ�T�	)
$rK �f������f��;;ݬ�i/ͦ��^-~�� �U����w����7 �1 y����6�Q!R�	I��ͺ�1}�uʯ>���z��_�H��K,��[ �خջ���py�����J�7ҒU��3]��������'���>�w i�!wBg�t���X�'eX5�:�%k0���I/i�lmy��l�>,���smb�������@z䘀�qW�W�%�� %I�_���J��b�������g�I9n��w��9����74�����
k7'ʐۘ�<���I�p�ek�� JJ�1fk�fl�>��X�nsw�,��u�.�D�좷sq y��\�n*@;nb+����H�B�������<���M�m��ݐY\�����Hu������{���������sA�y�ty �6�8qu����r�)�nk��ƻt�!e�r2����ִi@Ne^ֆkt�]Qũ�ݛ�l��<������#,˘Gu�+��?���7� E��l�ӭ�.��$.�L���֌L6N�h�c+;36أj��4֮���{����}��c�o��!2����Cݼ)j�q��`��JW):��[n`u���DB T�A$�����v36��ř��9����,3j%$�(�wu�}��,�m9��� �� �n�2��Ci��hj1�$�f� �f�?����������]���B�R�
G`��`qn�9�4���jmn��[�����%!R�U%������� ��M@{�9�d��Z��׍�����2�e�P�v�"�]�O���۳z:��׫p���[nFX���;���&�:�L@wt�h$��T�A%ـ����6�RLi���j��� 0���}���Y�;��K��=�"�������M@u������M@zS�SQ�T�G����`w2i`��8�u�մ�{��
�R5$|7g��}�c�y��������`~�����D�%%)D%MJn�Ir/X�v0s)�+�N0lvz��u��Փ��6��N܃Q�(��1g����,����K ���B�R� ��9������`�oL�������/{�K��BR`UIw�~�����$�$�cm8�M�_��f{Հ�x�J[`���M8��M,�� �n������A�Z�$TN��K4@u�����ꪾ�}����@s{v�mUҟB8D�Bj22�SD�u�C�i]]��0:9���&/m]�q�XR�N�+v37q yɨ������b��-mF �T�9����`nd� ���`9�Y�ې�<{�����{���߄_I�	}& :�L�:�=Dm��cJ8X]�vs��\�����+@�i�H���ɦ�TV�� t���J�$�(��*���ݬ���6����\��� �we���E�&6��7l�h��+�����M��i7m��Dqd��ۯV��}������X�7s7<��؀��t����]��+v�D&�7��̚Xt��<��_I����a���.쨝G@���f{��9���ꤱg����;���e7@���%�s3o ���`w���mI��׀sղz��AB�
$�Ww]����~8��׀w�xV��ABF�)Tt���Wm�����^�vN�Y�8 �,ͧ�498 �ji�����ܹ�@ly匪=Z��g�LGPM��mDҬ.f�N��EK�$��.WYǴ��Xu;N��^^ʳ���ǁZ�L�cۣc�v�t�AE�s�3�1�"�r��� 2�[�t���j�]�&ᵲas��2IB���~/���1�N�굤�k�m�ݘ؋����=>U���W�@����[5�N�S����g��[�9�;-�qٝ�q�m��<��n��V��QR���	���#�͟� �7o >�v��o���� �zOOB1���cJ8X{�,��,����K �����R�`nj���}U����I�������J�`���Y�;��K �se�s3e���6ТL������s��<�����n��6��tnm�������s�mÐ��٤��\�E�]�����N�h]]�V��s�������U_�a�o���J�S%ˈ�Uu�w�x�Q��Y!��WS!10��FӃM7��1�T��� �v�`]�v7"5�)�P�B��%����@y��������ܭ�۱$�B�����d����k�fl�8���F��Q�h$i%,��� �sP��o`���d�4�f(=�m;cu�vؙ;V+W۞ny-'\m��|���*bM��*)S�G`̚������{_9����^���M��t�rp�����ɥ����`��`g~ʹ(���!���ɷ*�=��峇�Q%?�����7��5{��t��)"4�J����b �sP�����_I~,�ƽ�?��*n; �f���bt��|� >�]�>��ۻ��-�Y,��a 8Q��7�y֎K;�淉=�^�s%DӥR�E
�(jH�V{���"�_9�	m�@;%�Z^�uvU؉Uw0��,�I&�=;���}��7�5X�KҌ_44�rU�����6wv��I9=��L��b�6v���	�� ����M4�}��=�w�r�����p���uN�9�W=�_������.QI�(�CR>����#�R_9�	nL@F2���>� @������'��챔���[�:}����۳5k�=Q��=���1���~�{� ���`N���i��v�� �B���	Tn���ʰ5w5�Y����Vs6�����A�����ے���1;�����5���4�4�HPԑ�ך�fmՀose�ř���jͨ(R����7"�9��V�}U��o�@7�p��+� �+�� �+��"����'�����Q_� E� U�� U��AC��TVTQ��*�� U��TW� �+���� �+���� 
����*��� �+�H��� 
���
�������)��F�5�Ԭ�8( ���0���         ���     J   8!	 ��   R�  �J��P(�U IJ�(�I PP  $AP   ��   �BJ    �)Ll i���[������m����M�� �J}ž�:��޺y=/g�j\ ]׶ۓ����k�����>�^��a��nu��϶��:�`0 �w�5;oK�[��qnϮ�p  ��BE  � Ud ޥW���_6�Y���oz܅�W�^/,�b���{����u��Ѳ]�w�N=���ǹF']�� X���|�z�����>�  `   ��=���{��{�z��������PT�Q@  P%�4��,OsS�]��at�Ȯ� 7*Vg�V�ޞֹ�:h��蠣��  :h�4  �
z"�� �( D 1��%)�@:i �  t�@u��P"P 8�!P(  ( b 3���H�Ms: @� e zgY@�D��E/�緋�Ϡ����;��Sɮ  {��d��x �m�'���ەU��ϛ{�r���� 8���u)��{�]�r�n=��>���P � 
 b�@}_m�wJ���ɥ���]���,]�:{������ۙ�w�>��U2{�q�s� �}��m�Ү��o=Q��;���r���q�Ѻ^��^��g{iﳩ���^ C�=��J� h�DL�J����O���OH� hت�m$� O�%M�R�� ��	��� њ��������p���g�ug��׼:��������7��DTTWJ�(*�**+�DTTW�訨�TAAS�����F!o�M\�6J1�2��t�¸š"B:at˛e�LX�
a)[�3E������|��$0"MoE��k�h��G9�%�����/�*P�A֏�6��~5Ô3��!�9���²�Iw6�X�����
q��������
b�vW�@�v}���g�_��D�cd�:F�40۲\t���F%��\�v!��x�HS 4�v���Mm�
�hv8?�)�u%�,�Z8�����}�$Z,
`po��nw[8&Յ)�>�R�I��|˭�v@�{������M����wÓ�(x�`T/�k�پ�f�]����JP�oNs)���@�:���3Z7������|��/[��6x� C��P�J�����{�4J��l��x�0��}�$���a�p!Hb�0����!�g	߮}B6Y�p!~��� �4�@��`���Z�w�4P$bѨ@��cNh��eÇЇa!\7rS2�KAu4ȗ��RX05�!C�Q��z�X�H�T"�@6$
�C��]��F T��4~h@�~t���XL4lf�2\�a%ޘl���5!!&ą�R� �$$ >k�HS(B��%�(e�if���R����"$T� �#�2C�^�	��cL��\4�˟Y6t�ޮ��R�tr���٨I��oZ��IR%pt��	 ��uvg,/k)iF4��1�Ѓ��C��&�HHF/p�e��		k�$ �HZ�b���WWS�C�>���\\�L�󠜻��6nJf�[4I8�/��{�i؁7��������R�$IS$��kz3 ��"1HŌT�����~H���A�@����d�X��aYp�l��k>��i�;�0�`X-0
@�Sf�u%0�m�|]�h�\��z\�&�hF���o�k
�:��>3���h-�W|��`B�i���a�e���Xm����Wѽ�kK>I~�.k|>9�	\�͜~��0�C
hћ8F@����cC>0-�]���tl��T���7�fݵ"P>6`�(�h��w�F�@��Sg����ѾO�Xf�O�;�bm�J�B�i4m�ɤ��h�	�JC#Yv|l�L��o�ۉ��C!77a>�kP�>a�1b��\c`T�p`F`R1�"55�8�4n��pѵ��;]nA޵�����nf�Cl+!"��.��B���+0�D��!�\ɚt�my�0�s���ψ��F40 G���04횺�d.|������A�F8Nk��gu�7Ѕ��\��6!��s�������g��}>��y`�BT��H��bQ�%D�C�B%Ff�2H�l�.Y�)ǐ5�6V��T��%�~
D)	A� ~4l��ԉ8E���%pe0�#B6XRMl�j854������SP�h!BcT�Ճ$��ו6Q��(�Q�x lr0HH�2c+F�H}��\Ѿb[��B�$�Վ��p���p8��`O�����#��/_�j����ڡ'W�����)3z���锕*P�l��c"G �cGD0I�����7e K).Bh�f�s�M�kP���&����9�G�%�9�>���0j��B�)*>�k)Xą�M��R_<�3F�*�x����"u>8������ef�e>�����T��]���<߂���>n�!@�HX��������h]��kD�۠4�3��k\M��"T�F��r����Cf��>4p�.kZ��&�Ev��q�]�d��w5&�Xs�5���a��)���h7�.�4��ˬ١�0��XBO��sf�le1��i���8kA��0��)��5�q���0�5
hܒ@�i�i��ލ�.P�m��~);u�5U�l���Y����X��5o����@�X�O������8
mx0ȱ�� E�\���f�o\���#q�n<��19rNp�&����\5
��-�bhH\֨m��������4��q"� Y�9�`E��h�\`A��ֆ�$���h�R\HSf��XB0��FF�"�`��aBd!FBX1"�0��d5�i���KjIW��"�q4O���
�@��
9��"K��w���l���!\O��l�cR_�50�	RMaD�bU��lÛ>��1�x&D�a�d*86��$����e0Ҙl�e�to2�`E�gМ���`��
G1L�0u��F�l%3F����^��,�Hk�CW�D`u��Y��4)�Q�&�m��4.�$FX�-��&�`s@�㩭H�0����%X5�Ə�i�^��3x}q�����IZA���V) �`� �N AbĦk�B�
m��!sN�W ��"E�p�ÇsA
˾q���l)��)S P#X�y<xt� ;!7�\5��jha�
)��]l�M�	π0i��$Qp�t��߉[��ut��!�W42�͑�CV��|�_F�͝a1�b@1 �  @��1��l�Z%R �\H��D^#�*���(�
�F,M�d�*�� h"@�Ӂ��a���O��P6�!�"U��j�LX@ū��\k����pT�� �@�U��P�-� �A�-%T�AH"E"�X-X�  `ă`0�V0�`Tb�cXB�����Q�U�)5�\D�!H�1�B7$��IZ@����V\0̥-Æ�v���2 D��T�����u"���7�����앯m�N���mnz����&2��q�+y�O�\�7�&���59��s	����L){W¡ފ�[wC{�m�n�wYO>������eS���Z��^�~(�z������U�jW��-KW�]ޣ���o#mz�`�6��6��G�߅w��>��m��-�,�Y�����g�Ǭ&���f��e�jk����w�P%ͳNMs���dѴ�3I�,B&�=�}���8t������>�@�_$j0�E�R(EH�F#"0RŉP!f��C#!b�$
�Ym7L����Jc0��!%%��p�0��������H�
�ơlltɵ�&�b@w��E�����K�ly
DLCN���@@��F+"1�1�0Ӳ	k,)0aXH@P�� XN�HU��)sBm`�}��!�#�E*K�"H �"b�p��C1cL�"l6���0ɑ��0��r/N|h�.k m T�I�ש���:08�`|4	
�SF�����4l�?5�JcMsg�!\4m��� I)�]:3g��D�5�|���d�!�f�mӇ �04�n�B$HPƚ����|h�75��&�БW�sm����6H� ��X0Z���X���ɯ���$�"Hp A�aB(�`�q�B �B]}��77��4��:�3}G�Ci/s�~c&�!�(D�= �H94KW�+�Ro$wN����I'y�N�{���`$  H    �       l���n$�.����v ��6��Y+kX9�Iוy�mp	ӃK�[p��m��U�mFQ|���f�E��B�����f�m���-� Am�l     ��|� �c��%�k j�!�  i]p-k��GPp�Z�
�J���zLQ����f�]'5�l�#Aw���Q�ut�X���A� 'n���djGN�2�D�9%���E���p7D�K��
s��-誮6t�g��㓶��ۡ��8ڎ2��1q]s�fC3ۀ�6Ԭ�;K]�v;dܷnz憸l��vz���i�{i�mUm����a� 8 �骪�+�������@�9p;uT�n�WLc��vWIͷU�]*� ���ڶ�pg:� $;]5�j3m��  $l  �:� �l ���m�MtÍ�  6�[@j�	 ��6��*j��ْ �j���]���[x��� �@ ��m	6�6�m����`�q�� 86�m�nܛ�m� p  p    ��g6�$H$   ��   @ ��88[@ H ��m��w �6V���ԩ˭�N�a���}�|$� �J � m�D��a,�Ѵ�@�  �m    �H� ��jU��Uڠ ����i $   -�   � i 6�  �   p�M� ��  -�l     $	�  m�   h �  8  � �a�   $�m�  $�[D�  :�&�-�o����@[V�ZҴ�Zm�,�[��:〷[m�(�H$l m p$ �޺��e� �`�`h��4�Z�` M���     D�   m� m��ڶ� -���m�m�          ��   �}�ϭ�m�      	�-�    6�   � [@��m� -���m�����m� 	8�����HW� ���m7R�EP���-��CM� �V��86���WT �6v�P������m����7m�  ��   m��[p m�m �[A��@   8�ޠ6ͭ�I<J\���gݳi;`  h��m�n�d�v�@�m�� m�崶�l9m [�u�I��aa����`m���[@����m����6� H   �.�H8���-����c���[B�8-�h[WU�m	:v�s !����D�] ����i>��[r ܴ �a������+��k��Xv'��*��R^V4�=I6���E�-���#6��Fݳ���[d���s����"��$   [|p� �ִ�J\ [�6Z���3�����ޭ��oku�bF6�m�mt��� �`��)�h�v��Փj\'E�@r�����öy��\m�� ��@9��/?���d�n�8H�rkz۸$H�6�[\8Yl4��M����   �Zζ�'R�l�Imp f��A!#m� N����6��&��T�Tj���i{e���*�\AÛ����`�&��+][�uh��YlK� �`�`�"(JJ�u���Z��n�\���3A�:S���v{!Ÿ���i���6�.�V�WK�-*����b 
�U+@[D��Z����� $�z��*�:�6��kX�!��"B�$�B�9z�� �T�cv��W �[r  �㎒�	��9��f�,m��3<�m@]��{ r�c�ؖ�����[USʀ��Cؖ�����@ 8 5�!:[ZE����h9��R� ��f,�U�Y:鱌b�1�d��kb�m6݃�[x�݀␴��@T��@c@T��R�`ةV��ڪ�	Rͯj�vs_k��� 5���-�M�n��k��o� �H[A6����)"]���6��/[H�A�l�h�7fٚl���i�ݶ  ⵛ$ ���{+��� [[lf���k5�s� 	I&���!�z�8��R���m[@&۳m��:��]�\��OkZ��m���#�i5�۶m�u�m�	 �m��Es�v��$`  4T�$[%�e�!��ʻ)-UUc���]p�%��;vGk���ICa  �%-��d��	�D�6[ԍ� �j��V����m�1�z�l�N88vC��p�����-v�UU! Е��$�7l-�gIsm��l��I6~��ﾪ�UU��V��]�	%�g55M�Ulޣl˴���*�R��um.�I����ֳ����8K)m$9��` ���\tm�Ɗ�m_v鳀�L� �m���[�$6�`�pH��4kq�p��g���<�tm�[@�� ��m� -� �A ��nmwD��nZU����ul�N���[u�1CnջWJ�UKC�-�(9���^�-���l�p����	��
�
�˴�Zm���6� �Yv�&D�{k�j �@�H�C�U�x�@�U Y�� �)��'J��K9k�V��&N�F�[&���[@5��
P�6�6.�[%���̟[,�|�c[@u��"�n�h�6ޓ=��7h���x)V��Tz�خ�CX� ���Kd�I;m؞�ݶ�t��⦫eX������P�Z��L�.�Ř��譨6A�P�e*�����Tzph��/�-��m��T�u��
�J��mWP�j��������P/;a�9@���s��G�)k�:����r��\	���kh�� ��jI��[�g]��p'A�Z�+���T^� �Kt�Im���
�.�:��@ � �r�c��6��̱��m� 9Ē[@m�m�u� �`-������u�rB���nYk���-���H[@���P6�� A�s��U��۶�u��k�v�ӭ� p&��|�>/��U�@U��6�nE�o� m��gR[ӃE    ����5�h  $i2�8q"��H�p  mm[@�e�j��K]�@j� m��/-����p �9����}�Æ۰�� ;m���p l��l4�   Ç[x�       >�|     [@��h��\si6 -�@ �J�v䅶A���m��%��	Cvw[�8Hm[i@m�8 � [@$��6Z h$[v�'	m m��-�VÍ��H�����	 ��8   ��        /Zm�H � "�:�ݻi8���6춉6� �U�A�]���Te[e�کVB�U��ioPz�C�rCn�Z�����x$I�v�]� ��i����Y;&w�4�����6j8��i�2PV�]F�hL�1kVݵ�j�HMu.`�n�C����8��T��E���p-� �n�k"j���yښ�x��5�Qi�m��p�e��M�8m��	V�[���ܳE�m��	@xm�[�{ m�Im  	$p� �[�]f�`$     5��3$ ����m�,�k��	�AF�\t���`��9J^,[�5��I΋.��:�l�C�p5T<�jݓsJ��[Hؚ�0T��kt\�UN6��p�[��O��o�$ 6��)����׮eJ䲇 ��GH�� }>��m 8E����M-�7n�n� 	  	� $�`#Z��h � �`  @���m 7Z�Hm�       � @  � ��   l m� h�kט�� 8  m l    -�[\Z�vVÀ �  ��t -�   l Am $ ���56�[   �M&� �hޠmƎ�am     -� -��  � u�����w��E���l m�8  u�� m[9lt5մ�.X�\�(��3�m�Z����W,�	�� �ÀlI����m9 [v�|�m�m��Km�6�l�y� m��[yU	53�P�uڛ6�GF�٭8�a�I��u�ץ�$�L�[��l,RN0$ pm�n�-�L�9�Y��� [%  K���֭�� �N��6�a�����((*lE��'��@8�P!�W���?Ӈ�^pA\J�_��Ep�/�P�x��X�@��ބ� >H�F��B��T8� �1B����>t�7����"G�*b t�<`(�@��|�G�p�tt��R��. �p �8��� ~W��h� ��_�'<"(>8���4�@B�S���"< �x�TV�XQ���Dh�_"�E*�'�8�:EL�<`G��@ڈ���� �E�|!T�!���A�Ґ �6|�U>��>N��t�q�@�@�(��-*���;���`�t
�80D>@�PS��"uD>H�*v �$�H�@�$c���	�P����8��T�/Ȱ"�l�">�7�X��*"������>-dF�F��	���'>M�A�6T6"�� !�MAG�8�A<��DO ��EV*���</���8��QQQ^"��� �{��~~mWVʵU��D��g�.s��%$g`�Ӆ�wE*�8�)��0B�k�t��,k�'�<M�bݣ��V�x�w&��{-�P�g�C�z��D��M�cJ׶�!nʻu+��V�g���62���`Z�h��l��U�mV�T�����rhݞ�6��a,AV���%����n�cg�ɵ� mzF�]6-��RԠ,@UƬ�Xv�Z������n� ��i��,�F�m��CUTpUT+(�vV�L��k��Jsl��ɹ f��Tĭ�]�VC��j����ƺնt�:tH�Yf	�]r�+s��ѷ;f@�k�����^r��!/\$]��d�r粼`���+컧��;��� O����;���s�,r�.��@7e7ONv;R<���:g��a%k��BH�\���m�q�j�g^9��s,Rd�i�#�f���u��3����j.ϱLI� ����7�K���������� ���+�NtT�#������-N^f�V$��
��2֩Ź5L���]g�CS�͟5�]����1�6�z�]Q�2b
$Sy��r����p� IY�X����꣪4A��G6����pp���n�*;pkWŠ띎�k8�e��[�cv�Dp�!�v�G�͒��fګ5r�5,qme���QE��w�6�	0�U����<��vF�wWr\M�6�݋G����%�v�g�M����f�d�bt7iZ��m�����h�lH Q�*Q;73J<�3�;D1k���ۉ.v��^L����ڷ���ѱ�m�QGd�m]J�k��U]Z4�Ӆv��qe�2�B��|��3;T&��-��mA��$
ul� -u�$-M�Sk�����
3eV�*���p��#<������h	$�-��l���6v9�)��v�u;-X��f������bwNjMhֵ�e��U�Ub@F�T�` �P`��
�
��Rf��5�#�N�����������_��&�&ɘ%BA�<��֛[�v�C�Zpne���x4��*������\�Ѯ�$�dz�C��['M.���޺��N�ܺݎ�X�<�2Q6����g�1s�U��^7	�t���>����}�w\�vF��pl�:�^M�f�j�Y]��/$ta���p>'RyY�u+��l��f�V:��8�Y��=W
�M ��ۤR.�u�n����ۅC9�QDq�����g�.^�dv��	�S¡�AI|��<ݳ ��Vz�W�D�LD���|`G.����J��WP�Y�y=u�1����L]��~X޾0n�h��� �KQA�����@�{����޹l��S����;e� ���tx����ՠr:�5�5��������X�Ȱ��r��ݰVN6�%�e'���>���lI�u��b4��dTt�ó���ME�mV����>���Xl�`�p�=
��V��j˩L���'>�z�� �"�"
�؎�؂�t�+��_S�}�� ��Ȱ����Wx�E6܋@��M�zSO�+_�-�|�Wx�țA$MF�$4}���Hn����y�f 8mRxF�0�G�p�;�����<�]�@��M�zS@���O$���IH�Ztظ��X���y�j�\4�$b�
Q�gW�5ڡؕ;V����Ȱ��o�)�wYM�>������ �.�\0�p�=�E�U�F�ޮ,k$kI���e4�)�@lF.��Eb���$���(s�Y�]�>�u�@����H�'�Hh����r,t�`�p�;jG����m�b�ݘ�Ȱ	��n�� �.o�o��?�O��6�:�''hg�Kx�d�C-F.�]lt
�gZ����c�ʶ��2G�<m��>�O��zS@�e4k�`���X�*��մ�ݘ�\3�%#�_��� ��0�j����E	�@�e4޻V���W����e4�H�0A �8�bp�?z�X��`ݶ`31ICHA u��|�&�k�� ����t4;�i���l�۶�u�0�M��!i��Z��ˣA�X���2��۪���mҜqG`�zn�f�d������zwϟ��Nبp����[0�l�?m6�ff ��� ����)�C�p�u��?s�h%� ��bD���ҡ���iة�f��X�p�7��wK��:7G�dY#�6܋Cs3��4�S@�v���.v��"j�R�� �� 陙�����<�a'���7$�D �
��� HE	� �$F'�o�*�V�fU��:m5͞�;mgۡ���c��;k�/�U��`��-�2���Di��k���Ym�����U�&�w=<s��6�8�^��8��Y�(�티{��ts�ڗ�όո]��{l�=fԛ��XS�����qh��^-�Z�ϕz:���3��y�nG\l�ulʋ�/�nv�V㳤����/+;�w ܼ�፯��ѵ��\[n��7nX�St�B��<�2���%��'�;D�<��	r$��F@�a"���}��r,d�O�� �r�]�c�&'��տٙ;�Ɓ����;���˩r`���8�x7��{�t�`�"�5�YMd�`)"bp�=��;������Cs1{n�@�e�b��0MG�n�f�i��y�f��fҼ��#�y�ٓ-l�U8��ڸ��PM�C��MδD �"�nf��ޅ�����y�f��f�����ǒdY#�6܋@��M��,��ƞ@��@N P���s_����M�;V�$z����������`��{�� �.�HP�ǒ(�ۆ�ٙ���~4k��{l���t����;�Ic�*Y�~�m`1?�{�q�u� ޲�q���oǓ&2)��������I����J�y�-r�'<���tێ���d�%�'Š{l���t���e4s�`�ޖRT�wi�ـn��:&"bR�� ��r�<ݳ ��tڑ�`��D�wYM��էٞp,O&���~PQ��;Ms[�h�)�_rױ,�D�pXۆ��r,d�`�p�;�� �]n]<�"�8��Z��h�Jh�S@��ՠw�W6H�s"��6��PC���ܕ���]�e�ۂo��9)͉ͱ��{����A!jH~���/YM�;V�z�h)ap��ǒ(�ۆ���0�M��`ݶgD�L�{~#� "(��Ln-���h����t��yڴWR����,q8વ��?�k�~� }���6�=32�$ؤ�4֜ ,h�FoK�h���bX�X
H�p�=��/;V����@�e4{�5TjA�v +��%y��c�|�����:Y�c�vM94�˺�,��[��Co�������=�E�N�w�mH�"�w6��X��Z�?z�Y�DL�艪9��[���yڴo
*,�y(���:\0޸`�� ����K�A!jHh�Қ�j�=�E��W�Jt�`�K%�]:�V؛� ��X�Ȱ	��n��@������b��M�1�!�@�l�g�=
b� p��J���Υșd�Q7��Z^JId��g�O7�φA�;��Տ\�������)Z��ug�2��&�g��,�uv"�ݷ.�RcOY����{f�۷%���Y^���\��%��Z6D�_<��J���Iu�3(��#4<�[�cB�(��KvZ(v����N��`�U��b�;������|}����>5�v:ܹ�l謻�unv΃]+.�f��ś�9���ӯZ�GM��Ęݨ�s�X�p�7z�Nr,�R����,q8�n-���=��0	�E�{\�2���EoK)&[t
��R�X�`i���1������|h�֨�rEQȜ4�E�{\� �.��� ��P���R�R�X�Sk 鉙����;���/;V�W�E�&�c2cl��t�XX��9u챮���R�B�C��kAd��ȱG��"�/YM�zS@��Z�]�@�w�u�h$##MI&��^���7�$D "��PE,�_�-�]�@�e4婫�l&<�ۡ�0	�E�{\� ��X�\4�H��(�id�67���j�/9��s�`����bT�U�V����:"gu���]� ��m`31�w(����.�*D]�,�4��Ε��\��T�;J��RF��t�n��N��F�q4������/;V��>�@��Z�u׊G$P�5��@{M��mw,�w,[�8��u=F
O"m8,iŠ~�ڴ�զ�?	��+������=L͏v���&wk�W_0���1�ऊD�dS����R�@���JfĂ�����R�	��@�֕M!֫�� �[P8���F0��	|#�iH6)A~�a�:��J���)��_Ɓ�� 8
�ڈ��@*�"0C��������8��'��߮��[;�)���&�(��Z����}��7]��3�s���D���r�59I���]�E�麼���|gDJB�}���&R��r�9�r舏�>���}�~��mץ�'L��Ю��!��rsjy��M�u�g�ע�	��;�;�b����o���䆻���D{o�~λ�	n����>1WB�V��V�+��=�ܳ��b�ޯ�X~�I���S}]�阤r���*-V��
�X���|�����jo������ܰ:!��
�-�n�N���Wtx�Ȱ2�<�t"X��R)G�W�����j�7Z����Ք&�ݧf��<ծE�{�� �� ��ϋaN��e+��ԗ.�����#�M���nmV0=jz���Z�K"s�N	�#�����s�`�p�5wG�l�\t�Zv��+t�wk �9��Wtx�]�@/�[�L�di�"�?�������k�`�"�%G(Wv
�M�'w�j� ���r, ����R'q
4�1�%#�?sm`��X��x�[M�`
��G������n�m����o��]��GPd�V�!�vUq�2t�e�1m���r,llWR�kz
�PlƷnQ�z%״r7#�ok�Q;��k�il۴��Y. ��v2�+�{(kulp�3��Vw�G��i��wdȗZ��#�ˋض�#��!�J(�"�=(7P��WO���x�i���<tYUzvy��
�gYw��{���{��}��~A�1�W p�콞�7I�ˬ�i�m7X�c����ɚ1�xb�y�ێz70�e�ݿ����O� k}}?�jo��B��y���J*�]Z�V��&Ro� ��WLL�A�]���D�;�X�]r�wWv��R�-]�tLBF���:�]?�z��Z�K��h��硑I䍧ӗYґ�]��[�����������:�x�D�ȱG��"�?s�h���]���"�;yJyj�°Iݜ��hǦt�ʹ-"b`^�N�v���c �u�2
F�DD#��9�{�f���u�~�m}��w,����݅TYWDWx��虙Ɉ���<�`����/ �BӔ���v�RWu�~�6��M�:b'�1Tn��������@��#N<�@��Հn�� ���r,���vRL�ݦݬw����k�`�ڴ���+�����q�@jcB�q�k��wL�jܺ�V�ޔţ��,;>E�(�&��8~��=��ՠ~�j�=��4�2�||�E'�6�NG�7��� �9��Wtx��Mէn�R�M�v�s�`�p��%D���]���^�ٹ'{��ܒx��M<P!Liȴ}�M��^��r,��X��%
��������u��3���:�X����}��w����ɂq�u��c^�W��+7VBu��fJ4����F�h���%v�k�`�"�7z�j� ��"�4+E;N���=�E�n�� ���r,���vRL�ݦݬw����k�`�"�?s��R9"�&㑸�Wuz�\� �9}_V�V��VUVu础M�+�Ȥ�FӉ1��޻V����@���h����WX�D�S��OhnR.�s���t&��] ��+=�k�����dF���'E�<m�����@���h���=�E��'N�]Yn�wo �}��<��X�H�R@�(Ȓ�An�v�'k ���r,ˤx��IV��%h�S�j��x�Ȱ.�������.r~xR~�4+E;N���<�� �}˺<��X��U��V[��a��mi�tp&����Gm˘�쬛��5�9#	�nм�q���l()���2;rmH��a�7[Ck�M���X�n#PsPdP3�L �=�;tMm'e���خ��cnڸ�n����l����ڵe�z�s7F����X�.�X����\�m�p������W@�x�T�s���v-�q�sR8��Ez��ݹ]�kh��Aj������{��~�����S[��ہ䋞�6Y����ka^بB�ЗH��r��C�RD��@�w�r�@��m}��wV�]]P���Հ���]]`�]g${z��<���/k�v�SV���m;I����p�<�� ս˺<g
��N�Z��m�ـyI�z<�tx�\4��bo,��crG�z���]���p�<�� �oLV��C��5�7h���g9��t:8	�m�p��HJ"L01
d�dy	Ǡr�@�ˆ�$x���N�NR�Z�j��Y�'>��7���I
��@Έ&�"��o��\�nI��|�]����PB����~M��<����I���o_�6�bX�A�H�q��z��uz�l���fb����@�����H�	�⺺�5n��:=�ܿ��Հy{]`m����q!u�10��۷L�'	&�Δ��՝�@���5۫���گB�*UwXG����<���/k�V�۝�y�"Ġ�r-��̉��Z�����?z�X ��v���d�FH��=��W�r�G�w�f�S31
&"
��ŀy6� h��aN�[����r� ���$x���Nr�J�h�j�%v�km`�WwW�5k��5n��=�m5B���AU=�E�,2���f�%4Ҧ^m�\<��.�j/]~��_4����E������u`^�X�뮏�=�ܰ:!��IS���Cv�[���9I����u�~H�����H�	��<S}X�Sk�~��]�Հ4���7���Awsj�U��]�L�m�,���ܓ��}����"�E�]�A"�#r'�'�����`�9]|UX��-BVU7v�.��������)?<��_6�7������H�:L��]V�#rI<�pM��e�ц3��������\��v����_V�� ��m}3?D��W}�`"~����]E�u���u�}31���*Z������/k��ba#��u�bV�DU�P��`��X��11M>��57Հj�e�J��V�X��`t�L/S�V���u��D��kϾX��ը�t�բ�� ����:b"v�������w���0�/B C�
�X�D��c�	Z�j{��B�*/��G�ϡ���D٠ځ�m�!�?��&�p6
@��*N�~M]T�k!u
�h��D "��cV��'�$�2�����-�В�(ȑ!�d8K��	I��#>C"lq5��"�����肖FoLH�@��BJ�0���Im�!8|+��)Ia�bF���HBj���Mj���F�F!Hԉ-R�V@�� F$�FW�Gj�n
`S,��B$U`�B!bD�AU`�BL�a�eu@�
�p&�B����b�4�

(xc��+*J0�+��Q4o��oۺ���N���� 	zvH�����e۶X�9������0�X^mm���rN�y#�:ښ�$��RL�(���.{b����i�I�E�VT+�cv���F��J-�8�ٺ(j�c�cC�3��tQ-��"�V��@U�_�g���[l)���vԕL'e��m�,�im����t��ɵ��!���<ԫmP.sj7NY�m�3�4�J�H�
V��e햪h�c���I�-�-�ڐ�;g�H jl[H�3�lٛb納[WJ��-l��m�M��)%����vy�N��D[Q �Ϯ��)�s�J�m9vه+v�,7���C��VC�v`�ڛ>wUV��l$+ɛ�!�H���3�nئ%s�S�2m��&��5mj���F��g�M�ˮ87�gc�' ��X��r��vSs�R�s��{u��`�6�C���4�.��eŕWF�k��v2
�s�j��c��ۂx�v��E9$�Ʒo*lZ�(����T�)��Y{4��sa�2��\��5m*��r�S��b���as��r8�z+�@g�m��Rl��hz�<�l1�mˇ�-���u�A�l:ꛛ�X�����&�;Q9�aō̯�l�r�.�c�P�m�e��7��yhˢ0�k���s��A���jܜrm��� ��h��nn��Gnnڭ��0Jh�[\�H�Pj�[���Wclo��ĭlޗ����l]��ga��5M�t���d��St*�m�����a˰i�Sc�	6�|$e���j�\��E���G��`�G��&Ơ�&:�e��@	3��������n�v��-*���Z��V]�pO9��c�-��̋�,2��D�>�X���彷d"�0��������m���v[jB��+��ڇgf�Z���Ƶ�7m�mVF		zP��V[m�^S	v�6�n�����]�i�n�j�	��p��s-j���2�����8���UH:H n�<�����t\��r��%������T7<��:�.UD��9+�,�L�����m f��#j�������i1�X��޺��FĐư����E��c�:^��;�t6�c.~�6>b�Z��l�e�]mT;�۱��=[<�sP���0h�C�k�z��.�g%ΞmT-Ր�˺Cqs;j�G=��&��B�VR�͊B'm�A)�m-�A������S�����`�#Fdz�6�l�����|b�uC{��4���.�����ױ��$�8n8�����=����~Z�t�O���`g�b �<"m�D�z�]��333�g�y���� ��u`[���&7��ةX���	YUUv�'�X�������y�����VO$d��#��%mk��57Հ~�6�:az�u`���oG�	Ǡz���>�s<<:w/�y>��<���&��W�T+�����%�k\3td�:3Mk+��N��#�&���!�����DF8�Ĥ����-���z<Wtx.�[I4+E;V�.f�䜽��c��uA����=}���o� ��mg�1��C�QJ-Z�(��@�w�z�������?�Z����;��^)$��r5"�=]���"�<�G�n�� ��)����-6�V���=�E�yt� �}����J�A�p�܃r&D��ju��͑u�,d��K�-�v!��t==������%cmݬˤx��]�������ՠ-o+�'�2Dۑ����5wG�{\� ��Wԑ���oG�$��9[��?z�Z\_W�W�꾪������=��Ԥ�-�Z����r,ˤx��7�˺���F8��n-��V}_}�}k ��<��X^����"d!���:�6'�&��==�.�p�n��ݹ&%V��"����IYf����]���"�<�G�v�8�d�4���8h���޻V��u�@���h�]FL"m�D�z�Ȱ.��>��仜ŀj� �\)��vZ��m���yt� �}}{�f�Љ�,@6���fy?z�Z�w7��œ�"m��޸`��'��7��� �����*v�Ol�;�M�Z­U�^؉���]�Q�9鼻��망ƚ��O]��m�cWtx�Ȱ.�����;��{���Q����v��<��1#�~���|h���]�H	��1�j�ݬˤx�\0]���"�=��n�5V�R�Cv�޸`���=�E�yI�8�Wwm:)[�v��9wG�{��\� �<w�4�g�g٘��
m>��%"�F{Vf�nݞ�۱q��:ز���
�0���̺{n%�җ)�I.N7[��7��m)�
�g5�X�ڴ�	��I��t���GO;'���:5�� �M�Rh��;��3Ƈx����F�k݌��z�.m�:��]�x@���t�ۣGH���#�(ճ���s�r+Dܭ�(��S�%k�$b�������[���f�������ﾎ���I���F�]V%P���F73\�hx��,;u�Kc��J~��$��$�O+UUb�Wu�}���`�n�{m�ɘ��*��w�E�����X��"�?&�gL�LBF�0���?z�X ���x�y#����)�r�O|��"�<�� ��#�7J�����n��tx�Ȱ)#�7z�{am��m+E;V�+��{\� �=�zS@��^��ҒG0rd1�0؞L;6Ѹ���lP�Mn&+��K�d��<4�!4�F8��n-��zS �����E�{�].�J�e�����n��+Ԫ��G.��k�`����y��$^��I`(�q�@�O� ���$x�\0߹\J�w�۱Zwo��"�<�� ��M�uz��U� ��X��"�<�� ��t�0]���"�=�9�����ۋg�Iu��9�i3��9-]�浸���dGk�t�N�z����޸`���=�E�yI����YLx���˺��3<H���,W�ߞ���-�M���Z�u�ܓ�g�w$�����t�� 9��n��S@����R`�DF8��UZ�?&�`��0[��:"be{g�-�̿HbP��rD��@�ޔ�9wG�{\� �< 㔌����M�k]���g�M�2+��НI!��3ν�|�d�h$���G4]���"�<�� �����B���iիn���"�<�� ��˺VtJF���t�UVZ�]E%v�.�{�.��s�`�%:t�����C��[�V����ZO��Cb%P�{���=c���c�V��v�f˺<��X���ݶ`13<�(밋��*�R.�Y��7
qm�H��Yp�f�:Fu�v�3%avu;��q�J#QbR?�{_�-��zS@��^�ݏ�0J"#QA7k �<w�.��k�g���<H��/��#0�$��;���5n�âba/mw,˻� �������
ݻ���9wG�{\� �<w�����%w��iիn���"�<�� ��˺<���|UW�|v�o��/nj�ı��tkY�;cj����6��Ӹ;;oZ}��1�m��.�+�٣H+T�7�XS$�h۳Q�������{&S�BX��r�����izݓnݶ��\cd�w%�o	�.��ɠ4sZy�ɶ�n��!^Y�G*h� M�r��MӉ8:w8�B�0��xoj��7@�7h���5�3IA����뚐pq��<���yُ����7��t����Ѯ��H�x����s�9��#�j7<���d��tq������~~ǀn�� ���r, �"d�N�L�8�ܑ��Қ.����y���=_}��.ev�x�<�8�7�tx�Ȱ)#�7��{e��)�����T���=�E�yI���uz��ܘ%�(���@��u�{vـj�u�~�m`1	����.���dm͠���m;I4:��8rka^1X����٢q�\����v�@���_� ���r,�H�s����bi
8�4]���<���  A�`���;��ܓ���7{�����
�cN�[wo �9�$x�\0]��>�2�$ȱ�JE�~Vנ{�Jh���=�E�j�d�N�]]�m�n����tx�Ȱ)#�=[����$��PM۷�u-�#2�N��؞��	u��RLj��
�x��;6߇��?z�X�ۮ�����v�,�ȅ��iZ*�[����r,�H�ޔ�9wW�wc� �DF8��n-�r����>�;빳�+ς�Ր@%ck	��N%�U~F)d;��q $&'T�c�]�$ Aͫ�2D8q�*w�����bH$b1�"�B �KH��HMZ!�TٯjL0��~JLő ��D@��E� 6�>�'�DV�PV~ �0q :��4�:T�00T��1��)�DX!�xuG�
P:*�@t}��~�~���j�?s3��%"k�i'o ��˺<��X�����Z�E1%r'�uz�]�@���O���@����Ȉ��LL<,*�wf�E��6[�E�ƛ��7 �.��j���]��9�i�m�?������wV�m� պ� �uX�]ŪE�i]��H�޸`���=�E�j�r�'N���m�n���V�:%/mw,˻� q�
�Qn��lv`���=�E�yI��{!�oO�s��V�,�I]���X����p�9wG�n�r�j��^u3K�E"8f���3e��/�Xk��9�@���EYȚ71>m��߿\w�.��k�`�t�j�v��wv�v���`���=�E�y[^���u�$Sҍ�#qh���=�E�yI��,v�[�НՔR��uWu����ܰ.�ޭk@��^���z��Ǒb#Ɣ�@��� �}˺<��X�U�}��@�����Aj���Q"^����}�y!��N�`�8���=�x�����;�v���8����0[��5 X�ɔp�@�OmO�T��mQm��;�]]2<Oj�B�3�,]�av0�L�5����,d0�k�sm*�z}��0��[\����\��8�5�vT�=+^���֝��ۙ4#����ݏ]rax�e:^.�L�r���R�*��1G?�o���ƞ~���{�=�|0\��ֺs�b�Xt:i�J��c/\i�k�U�쵌=�m�'��e.xy�iY�??ߖ��,��X����9�Un��lv��`�"�<�� �}��õm*���[� ���$x���`�IV�M�v�X���yI��,��4޻V����8��XH�q����;��{\� �<u�HM�kaP��R�9tl�`L7�r�7��nҽH�ǫvM9005
��k���Kʹ���Ȱ)#�7_E�n�+q�\ѩ�.j]f���'>�z��>Ub����������]Հk��n� �i�U�n�R-�J�`RG�n��%�%4޻V��m\x�<�"r6㷁���Vw\0k����� ��Q&,�&0IŠwt����j�<�� �}�㖅t�k�ؘ�J�Dm\3tf�G3V��f��9�u�r�,���r�Q%�F�G��ՠ~Vנ{����;��#M���&���@�<w�w\0k�`�t�4�k�N=�zS@��M7�<ŋ�v���ec
$4*�}���U�W�~�]k"���#qH�4�`�"�<�� ���k���;�ӱ[�� ���$x�Jh�)�><~�Z�(
G I�L�R%{;WXXX����L���Sz`�zX�g��ޚvi۫T�t�v��#�7z�n��mw,WqT�*EE�ګ�����=��`�l���%1������A�A�A�A�=��lA�lll?��?Y��&k$˚�y���6 �666(E^����؃�lll{����b �`�`�`����f�A����~&���n�������56 �66/�Q2=�����A�A�A�A�~��͈<����}�~�y
XU?D�@� ���}6 �6w����������ޑP��E����� � � � ����6 �666=�{�lA�lll{�o�؃� � � � ��~�v �6664���]kk�Yʀ���7]WK�7M�n�ŋ������nܙ3r�H�2��f�an�� �666=����A�lll~��lA�lll~��~� ?��A �`�`�����؃� � � � �����)���2ɬ�]K�]�<�������M�<��������b �`�`�`��w߳b �`�`�`��k߮�A����t�_�R�L�u�浭M�<��������b �`�`�`��w߳b �`�`�`���f�A�������A��������He�a�Y�2�j�A�lll~���lA�lll{���؃� � � � ��o�؃� � � � ��~�v �666?���\0њ���˭f�A�����~͈<�������M�<��������b �`�`�`��{߳b �`�`�`���"���뾚&\3�fe���6��V5�u��ڢ�U�IM���8h�c1ñ0�1I1�F�;�sd'FcZ���a��\�b��;���hkx'8�5��Blꗴ�v�P����n�>b��m�*u`��m�&�[���\bIC$��	�mp֢��(��+1���ն��4�ڌ�R��k�ءڣ� �e�:�JA�Zp�����������w��6ޢ��ŕV�2�l�=K�Tq��6z��݇u��k3VkE5����%�gD��`�`�`��߷�6 �666?w_�]�<������~͈<����{�~�y����څ�Z��ֳ5356 �666?w_�]�<�����A�����lA�lll}�~��y����y{W��Ys2�Xf�����؃� � � � ����؃� � � � �����A�A�A�A�����A�A�A�A�����A�lll~�_��S35fI3Zշ5�y�}�6 �666?{��6 �666?w_�]�<������~͈<�����������љd�f���Y��BQ(���D�������X�� ����>�L�]��WpR!e�J�����sr�3J���)k����z��a���|;&;�$��5&'$��u��@����=^�z��M۔��Ɯy!A�"�N^�پ��P�gow�ܓ�{^���r,)ԥIӫ�i�m۷�jޏ �u� ����>�8��Un��l���`�"�<���5oG�{e唑v%Wvݍـ{[k �&"=M�~v�,�� ��_uM�5�BYƐ&�^7���Ji��+��gdL̏���7H�F�"���<���5oG�{��{\� ����T�.���N��z<����Z��^��${_��(F0#qE����Sk�����" ����]����= ��9����0rcrHh}�}� �o� �����fa6��ό��bN<��ґh���ٙϧ��$���=�E�{zS˶�J�&)zN�'j���i�5���d4OGa�܈N�F2ф��30{�kq�x�c��ێ?�r����p�=�E�yI>�8��UL`'��қ����f6u��@�����W�^��۲d�ؠ�9�4ަ��6���KV���|`�����1�qh}��b����@��~��;���rUP�"�:��(�@��w$����k)��FI2��Uu�y{]`1-�����X�mz�+X��Q��$���;$\����5;;���v�Ig�{$DP���]������)�~�ڴ����33��9u������91�$4ަ�tD��BG�wV�_V���eB������HV4���$x��Xt��LD$۾0mw,ɲ�:�L �m������3�1s���-��@��m`}13+��Հt�ur.�E�\�	��;��{\� �<V���8��v*��B&�祎E"�>�T�x:~T���H��@@pl�m$��H�vT>D>#�DaF֐��1q ��`�B��3| � ���0��5�-�@ ,���Z�T�#�i����70��3�A �,^$E��>84?��{�_��[B@ �ؗ�R��ێ�;�6���w]lp��D�N%��,�%��]���3�\�JZ����7�	�i�<�[�l��Av��l�# 6�UR��q�4�Q�k�dQ(UT�-Ӵ�:�Z�6����IK�N^���ln�J��j�T.�Y]	lnm7���A�#�ذ���M����4dX��gD�[vԻZE��8x�%Vm�ZA�i�Z��]&�$m������� ��p[;n�2.���%l��+]*ʃ8��vI��h�	�i�܃�#���C�U��j:�c��a�c�2�)5�Ď��;s�y6�B�L�#):H�X����#���.=����<���=��8�\��ʜ�������Ӎ�An�z�ۭb��5�l`9� 9�"5n�۬��!�{q��LN�C/eֹ��8��]oZ�3�P"��j���8�؛�����!�q�T��aYˮn#JvT��2�ts���]U�H�P�c2����u�-�uvI�I���m�����m�C���� ��K��CX^�˘���gx9GjK6����gq�ml�C��X�8E�
c��E�����d�ɱ�@���	����^)Ü\��ko"���;9��u�Ő39�7OX�!n�==��޳�5�F�}p��n0x:69vݹʓ .�Pi���fL�ld���rc;:��;f���{C���KV�T�^�j�`l��psPPIK6�]�l��@m���n!��T	Z���8�.��X�2�l����C�uÎ�:.5���f{q�����u�ц۸_@��Sk��P�����Zf�ݵ[�:����3g�>�:=�%���Ʀ���-�U^�yX
�l�C�ۖ�L�T�m@WTmez����IY���)�m���[.�-�u�$%�Q������ɛ��nL���u��K!�tl��3�]�.r�I�cM�?=�{��{���۳�p�C1�*�<v �\@�*��lCJN95����f�nώ*T�'����s�ĆҴ�l7��i2Ճ�'n�iVS;j�mۊ���-�J����HA\nN��q�v�zֹ�^��+�Z��%:SI��QNl�J�Sx��Ȇ�Tm�>�{u�y�;g��t���sH�<n:�*�[��m�nN�M;�Sk�����f�s�d)�..Ձ�	�fR�u^�F��fJ/��]j�eՄ���c�B�<��A��K:蒠��4����������sf�26(%�F�G�����@���@����陘��Pwu�`���UIZ1���h����f��Қ�)�y�癘��e�H�6�0�$��}׀n� z��۬̭wDZ���ª��蘈�M�� ����6��b"R��x��Q�ҫ� 91�$4�S@���@/[4��������P�5�z��q��]�̚�<Y����;����ѵ��k����z{��͸�,ID�p�_���@/[4��/YM�hگxA�8�qǠ��o������D6��O���_� ߝ�`�n��Hr��"�]E�Z!U���� z�}1)ywu`�女��.ɍAA,r5�8h�� ������L�����r�h��R'!�~]k�>�������|h���w���S$h�i$n�;t<��M����T�]\��^*5��$q`ژ�rD��@/[4y�M�}3�z�W}�`⺾���(wb���=��3鈘H�����Հ����q�Z�D��@rc���~��'/}�܏���` ��?� *b*b �ßu��ј��!*��P����������� >ﾚ����z�h�j�I��㊪������ݳ��s�� ��o@��]QD,$J7�bs0)˛Rt�6�u{u�t�2Lj�����#�hϊh�S@���������v]�+�E]҄�� �v��H����5wu`��3舙�H}Gqp
��j�ګ� ����6����"�����;����Ѯ��J�q�'�궽�)�u����<�@��N q >Q�>����3rN�?��,���$hnM�)�u��*�� ��4��3�]�?��1�M�^r�F]ٰyi;j�h��n$�n��X����I�֨��Ly�z�O�@i�X���|��8��8��J���+�
�� i�Y�11�ow^����h�>4��ĞjA�z�h�L�;���U���>ub������S4�)�4۬����v]�+�E]ҡ�f��e4
��@=���)���O� U�T�Ĺp�~)bX�mUi��;/;,#�Bd��Ÿ��6�;Fж��%�VDS��P*l�:�ǀ�6΀��Gت�%�hLi��n��y�V #�c�����S�yz϶��D��]��)k���Ս���벋6A���׈�vh����.;K���t��J�gE����A��������h�6�f�z�8�bWm1�K.���������/���NSƈe���9[��K��W��vkvy��]Մ��]�L�#QH���w���m�@m�#��b#��_��Q�]Z��\PU�B�� z���11	��>�0�����3ď�W��&F0����t�F ��0��^M��n���I�6��2ٙ�b�v��ߞ�WZ���4�2ס�H�,Q�n��?&�`�u��g�s@�r��(�L�")$x��#�ArW6�1�;IWk*8��,]ӆ��x�N��������7kF`����fb#陘������.���w
.��������3�]U}T����#�oKΙ��H�G�qJ�bQWt�+,�=��������ψ`S����V�V`t��J�wu`���ψ`޸`�t�j�e�۴'u�����/�bb{��Q�}��~m��\wߤ�1��a)��Ƅ��/n����>���=�V�	��`jR��ӹ��*��t�0��f�6�陘��z�4��?�'2jDF���Z��$ywu`Z���љ�3�L��Q�#���BWu�]Qv���ﾬ�z<4�����U]9�`Ϣ�J�x��# ���q�}�fb����8~0k�)#��� 7J����%Wu�n֌�:&&=��~˻����I]*_]4�ВE���6m���)qtI	[۵k�<������7+�o.��kYKu578X���]&�X�%�����ND�,K�ﵐ?*NDȖ%��k���r%�bX�����JhՆj��54��bX�'3��m9�R9"X����D�Kı=�z~�ND�,K���I���D�5�d�&7����
���*�Ъ�&?��,K����Mı,K��g�ӑ,K�����n%�bX��{ٴ�K��{�? ~�C�sث[��{���2'��O�iȖ%�`���4��bX�'3��m9İ" b�Dt �&wߵ���bX�%��zg�	̃##P����1b<�g�����Kİ�?k��f��%�b^���q,K������r%�bX���~����6��������.�ݤ};���'�%�7�祈�z{m�M�=O*թ��%�bs=�fӑ,KĿw��Mı,K�k��a�B}"X�Lk��0�D�&0����	TR���ֵ�ND�,K��kQ7ı,N���M�"X�%��u��7ı,Ng���r'��?�:��K���અVAV�WvLa0��L"c���r%�bX�wY�Sq,�!�2'��߳iȖ%�b^���q,K����眺�R��[����K��BD﷟�Mı,K���ٴ�Kı/���q,K��TI�=��q���L"a�}e��qh��j�U�Sq,K��{�ͧ"X�%���A����Z��Kı?{_���r%�bX�wY�Sq,K��c�_o��p�߭��7Uj}E�=��Wnu�x��b�1�����6���80��ia����;�Bys��[*'dl��HY��F4utnt�\��4��E��],\�����N�;r��z.���]W&�zz���X
�ݱ�
�=;��]�����1u�\s˱Y�s+e��[:��i�[�.5�t�&N^�1�c��S��kP�;��hF�V�������er5�lN:�덥��M��\��Kk*�rd����:#�����S~�����g�ľ��j&�X�%�ߵ���Kı>�և��DȖ%��~���r<oq���}��=��b�-ow��ı,N���M�!�����,N�Y���Kı>����ND�,K��kQ7���,K�l�_�R�L�5��˩���Kı;�g�Sq,K��{�ͧ"X�%�~ﵨ��bX�'~�g�ӑ,K��_n��5��s��j��Kı9��iȖ%�b_��j&�X�%�ߵ���K�� �"w��֦�X�%�~�����!����33Z�m9ı,K�}�D�Kı;��=6��bX�'��z��Kı9��iȖ%�b}=����Ssڵ�KCڳ��2N-0X�eNY��ܓ��vy�������<����O\�2�kZ�Ȗ%�b{���6��bX�'��z��Kı9��a� ϢdKĽ��j&�X�%������Xkf�)n��ӑ,K��}�H��πF���X�P����ND�=���m9ı,K�ߵ���bX�'~�g�ӑ?�2�D�?~5�Z�[4j�5uu��ԉ��%�b}���6��bX�%�}�D�K�"{���6��bX�'�~ޤMı,K��;�踠*��Wu���L"a	�֢n%�bX��]��ND�,K���"n%�`*���]D���fӑ�7����_�t:�=�����7�ı,N���M�"X�%��*G��sR'"X�%��~���r%�bX����q,K��	�����h�欚��9n6z�Mu�H�G4��"q=�Q<Y��Z�=�����)����gf�%������K��?���D�Kı9��iȖ%�b_w��Mı,K�k��iȖ%�bv>�۰���T����q,K��{�ͧ!�!�(��MD�/���j&�X�%����?����DȖ%&9�XLa0��L"atr��	TtYZ�35�fӑ,Kľﵨ��bX�'~�g�ӑ,h�"[4f�i�U��-�p�.�hD7|%�N�� Ȧ�%�0iS@��O�".����,�N���
N��MoJ��"��% DҔT�"��F2F"PHDh���@2��h�6o�E�aԖ���m%$�dK3�4$�(�0� �'���R ���0@M�A��(
�^*. ��i�Av��!��/@�$ND־ޤMı,K��{6��bX�%�/p�L�Mf��f\�kQ7ĳ�A`dOw~��ӑ,K����ԉ��%�bs=�fӑ,Kľﵨ��bX�'�;7�u�5�3Y�S3&�ӑ,K��}�H��bX��?�W�����Nı,K�~�֢n%�bX��]��ND�,x�����)�3unz�
�@���u��aE��YNۨ��g�!��Jplְk�vj��W5�q,K��{�ͧ"X�%�}�kQ7ı,N���M��'�2%�bw��֦�X�%���OL�	��2I�֭��m9ı,K�}�D�?��2%������r%�bX�������%�bs=�fӑ?�Dʙ�w߰�����V�����oq�{���6��bX�'��z��Kı9��iȖ%�b}���&�X�%�b��9����0r25o����#�RD���ԉ��%�b}���6��bX�'���D�K����!T��?)���?dN~���iȖ%�bvo��j桪\��ԉ��%�bs=�fӑ,K��u�X��bX�'~�g�ӑ,K����Z��bX�'����}�f935&������V�Y�
�)�bl��
��-<:�d�k�������7u���CY53Xff���;ı,O~���Mı,K�k��iȖ%�b}�g�Mı,K���6��bX�!�����nzz�Th���oq���w�vzm9����,N�Y���Kı>����ND�,K��ڱ7ı,O��o<���̺��56��bX�'���D�Kı9��iȖ?�R"~��j��Kı=�z~��7���{����z�k�715�n%�g��ȟk��fӑ,K���~Չ��%�bw�vzm9İ?�BdO���H��bX�'��g�Mjk!&kZ��Y��Kı=�{V&�X�%����ߧ��%�bX���z�7ı,Ng���r%�bX��N���{�O��o�����93n��"!�>'��1��&���+�ڛӝ'zRR�)�*���0s�hݱ:r�g\�.�����9J���ղ�vW����q�[mnŞ��ړDF��v�b�;��q.�E�u��O��(�ZN�ñ��燝e�9��rt��z4���ն5J�t��p�It����n�Q���Kn����Y���f����j�JĦl�\�ճ�E�Z��h�[��ӡ�ڼ��""��k������>?#���b�X����bX�'�k���ND�,K���"n%�bX��wٰ� �DȖ%�����{�oq�����?K�vi�SSiȖ%�b{�ޤMı,K���6��bX�'��j��Kı;��=6���Q�X��b~���a��:��0��H��bX�'s���m9ı,Ow^Չ��?�ș�ק��Kı?{��"n%�bX�ǯ�Թ�ɩ��35�fӑ,K?�D���Չ��%�b{���6��bX�'���D�Kı9��iȖ%�`ޝ����kf�2�bn%�bX��]��ND�,K��+����H�D�,K����6��bX�'��j��K7����~]���9�n���e�
������)됋��XR�I��j7�:�l�[�Ԑ�̺��56��bX�'��z��Kı9��iȖ%�b}�{V&�X�%�ߵ�SiȖ%�bx���5-��i����3V��X�%���}�NC��T`R8�Tb��PǑ2%��k��Mı,Kߵ���r%�bX�wY�Sq,K��tC��Mjk!&kZ��Y��Kı>q,K������r%��E!�2'}��jn%�bX�g�~ͧ"X�%��w3ڦ�5��]kY�3V&�X�%�ߵ�SiȖ%�b}�g�Mı,K���6��bX�T����X��bX�y��E5�A��dj�3��#�G�b}�g�Mı,K������O�X�%��k��Mı,K�k��iȗ{��7��~}B�vu� �m��uI����K���mϜ,�d���x�I����7E{V���f�jn%�bX��wٴ�Kı>q,K������(	>��,K��~�7ı,K���3��v��g�����oq��������Mı,K�k��iȖ%�b}�g�Mı,K���6���r�D��~����s��*4ow��7���x�u��m9ı,O������%�bs=�fӑ,K�����Mı,K�vng�S5�.�.�fMM�"X�~��~�7ı,O���fӑ,K�����Mı,�&D�w��m?��oq���~���%�=��+'�q,K��{�ͧ"X�%��u�X��bX�'~�g�ӑ,K��;�ʛ�bX�'�C=������Z�4�k31z����д�ڵA�������yw])Q������e����N��5O�������D��j��Kı;��=6��bX�'���T�Kı9��iȖ%�ow��_���6�K�7����oq�k��i�~�DȖ'�k��Mı,K���ٴ�Kı=�{V&�>����w�����o��Yn��Ikm9ı,O���H��bX�'3��m9��"~��j��Kı�8ɏ��&0��"��w6��FfjD�KϠdO���6��bX�'��j��Kı;���m9İ �����(�����(��P��o���q,KĽ=��e�����a��ֳiȖ%�b{����Kİ�R>����O�X�%��߷�q,K��{�ͧ"X�%��ٲ�5����nl3�˞���
��u{r��ś��ȶ�==2����{��ı;���m9ı,Ow�ԉ��%�bs=�f���Kؚ�bX�߿�q7ı,O~����5�!u�u33T�r%�bX�﷩q,K��{�ͧ"X�%���7q,K���充�H/�3�?�d�r�%̙�0u�O��~͉ �'~���'��]�6��bX�'���D�Kı9�u�Q��H������#�G�{��Mı,K�k��ӑ,K��}�H��bX�&D�_��6��bX�߯����q�*\V�|��{��"w�w��r%�bX�﷩q,K��{�ͧ"X�%���7�<��,��������/�s25o=cĀs�/�!�ʎYF���<�}��gK[®\� ��vk���q�a�yl㫝��ۮۯR^���]�0�,�u+;\.���3� ^���n��3��q���.7"m����:ۖ{�ݍ��V��\�����v	v�ʂ�qr[�2��=s&�(�^�՝<����PZActM%�@焀�V��6d�1���X~5¥a�A�ܨհ����I�)��W'JK.j���N�����o�Ĳ�'f.�����"X�%����z�7ı,Ng���r%�bX�﷩q,K���充�Kı;Of�2�N��e���q,K��{�ͧ"X�%���z�7ı,N����ND�,K���"n'���,K���3��d��a��ֳiȖ%�b~���D�Kı;���m9��A!�2'�~ޤMı,K���ٴ�KİoN۞��F�Y�̺֤Mı,� �45�����ND�,K����"n%�bX��wٴ�Kı=�oR&�X�%����ST�u�u33T�r%�bX�﷩q,K��{�ͧ"X�%���z�7ı,N����ND�,K�{����;�I��a�Oaqs]be��s��L��g�9���/_�{��?/���F�5u��ԉ�Kı;�߿�iȖ%�b{�ޤMı,K�k��ӑ,K��}�H��bX�';�w��k2�!&kZ��Y��Kı=�oR&���Q��c���b{���m9ı,O���H��bX�'3��m9ı,Ogq��7�RF��y�y���#��gZm9ı,Ow�ԉ��?�2&D�?{�m9ı,O���H��bX�%���{WS3F��Z�5��SiȖ%��C����߿�ԉ��%�bw?�fӑ,K��}�H��bXfD��a��Kı;M{E2桫e�nfjD�Kı9��iȖ%�a��ʡ_���jD�%�bX������r%�bX�﷩q,K��d�w���msA��ip��է%s�#ש*�cKW�qp�]tgN�s,��լ�+S�����ı=�oR&�X�%�ߵ�SiȖ%�b{�ޤMı,K���6���oq���~[s��*U����X�%�ߵ�Si�~H�L�b~���D�Kı>����ND�,K���"n%�bX�{��y�5M7Y�S35M�"X�%���z�7ı,Ng���r%���P�	�Ј� �/��ƐZ���x�2'���H��bX�'�����ND�,K������j�5uu��ԉ��%�bs=�fӑ,K��}�H��bX�'~�}M�"X�%���z�7ı,NwDﵐ�e�BLֵmֳiȖ%�b{�ޤMı,K�P�k����M�bX�%����z�7ı,Ng���r%�c��}q�~� �0�ŉ��m�ݺ5Y�r�,9i���u��i��-$���㱭k2\ԉ��%�bw�w��r%�bX�﷩q,K��{�͇�}"X�'�~ޤMı,K���?j�c�fFH�Y�g��G��1e�<�ı,Ng���r%�bX�q,K���充�O�ʙ��c�畎�"6���oq���_�~ͧ"X�%���ڱ7���DȞ���ND�,K��oR&�X�<oq���_���fyZ������d�=�{V&�X�%�ߵ�SiȖ%�b{�ޤMı,�Q�N+�U5ȝ��߳iȖ%�`�ޟ��j�F�Y�̹�X��bX�'~�}M�"X�%���z�7ı,Ng���r%�bX�q,K��u����ۏ�@k�ٍfى츸��K���ڵ�g�x}tL���]�x����=���,K���"n%�bX��wٴ�Kı=�{V�@���,K�׿�����{��7�����óѹ���"n%�bX��wٴ�Kı=�{V&�X�%�ߵ�SiȖ%�b{�ޤM����S"X�{R{��f]d$�kV�k6��bX�'�k��Mı,K�k��ӑ,K��}�H��bX�'3��m9ı,Ogs3��f�Y%ֵ�35bn%�g�a'��~�ӑ,K����ԉ��%�bs=�fӑ,K�I�?{�bn%�bX������Z��E�Q�=���7���'���D�Kı9��iȖ%�b{�ޤMı,K�k��ӑ,KĈD�$`� d��� ��1J*P��4�YϔO)�0�E%�	.�5�!�@���|@7�B �3B�
-���H��EGdf@�n�6R�d,+�XH�$�a
0��|tc���b� |t7�?tS[>�䀶�	kiWI<r��uj�V���&'N�i�;m���sQv�4Î��eu�m�	Mv�oi&��w"2��"OB%���v؀�k�Q+R�[@e�:�)B78�a����T��v6ˢ�tjUjS3`�����yܡ�q۹��4kr@ڶְ��4d�F��i����lX`Wh݀�Nض��KMk�D,k[H�y;�.���W��W��[M�l_-޸lI�k(UT�5UJ�$���[;4�\+��:����v��ԫq-cmmA%���N[c&r�z�ݫ(��V��V	��W2:�vKs�yEx���K���Y9;4j�zp�/WFLL���lڍ�ם�\�c���u�K#`�ͣə˘n��d�۪��uջs��1��(v�w�a6����t��6G]g"�/!�*I���7V4'm��
��ƫ��m���z�H��̕@�uq����3��G5�ǁ�7a[q����l��#�$n׎��m�s/;+��r��v�hc=;n��N�ܼ��RW#ˣ��t�S�k4��6i��mn��{bd��N9��t�T�0;�V�K��)tgaр�õ���TM����j��y���E�����R�Z��x�;�m_(Z.u��b���w���ծ ���8۵k{U��+���s/۬/�S����؄�%M� �+e�v@�ݒ��;s�xj��v��xj�[�����&YXm�D� �.�����,��SC:b]b]��l�<F`���&` E���k�.�nˍep����%��v�6NA�x�t�m@F��3J<�g��^�ү'�p� tΕ��K n�M��z�s��n۵�G��m]	E+��s��Qev���8���)V�������THظв�^Ci8"nPj���rګ��WT;��e�n�6(b�b�9�ݹ�`Z5�;6�Il!r�z�B��1�Fk0�k5n�fjj�t�	�>M�W@8�'��v$ڈi�0@T6�P���'�ч{���w�����?�~��xl��rkW���6�\nJ�"�L[��n���VP��Mb;
� � �;�)%fHs.����He���͙�Yn� N[�5���p���n.)�Xe�$x� =����[m�;��r�3�;WZ�{.�r]�s���V��ȗn4�V^ڲm[(����5�r�cJ[m�N9X��)@�yx<-���; �ihի�=���Y>|_8�6�����..�e��Gӝ;k�����,F���o�ܬt�+H��bX�'3��m9ı,Ow�ԉ��%�bw�w��~F}"X�&9�XLa0��L"atr��%QQv\�a��ֳiȖ%�b{�ޤMı,K�k��ӑ,K��}�H��bX�'3��m9� �S"X7ߧ캓Z�Ma��f\֬Mı,K�׿SiȖ%�b{�ޤMı,K���6��bX�'��j��Kı>�a�j�����2�ff���K��RD���ԉ��%�b}���6��bX�'��j��K��@dOw~�M�"X�{������Xvz715�����D�9��iȖ%�a�����V'"X�%���ߩ��Kı=�oR&�]�7�������Ac�¦�'p�m���g�������Kʚ��z=W��{��{�m��);�f1O�����{��7����7ı,N����ND�,K��� "��2%�b}���6��bX�{�?e_ӕӝ�P������oq��k��Ӑ�+T&�T�'"X����D�Kı;���6��bX�'���D�O�PʙĿt��ں����Mj�Z��6��bX�'�~ޤMı,K���6��bX�'���D�Kı;���m9ı,N�����j��,�r�Mı,K���6��bX�'���D�Kı;���m9İ?"L��߹�q,KĿ����`y�g�����oq��������D�Kı;���m9ı,Ow�ԉ��%�bs=�fӑ,K��S�����6n�
v�����gJ-6X���h�I�-S�g�F;,�����i�|gU�k�e˭jD�%�bX������r%�bX�﷩q,K��{�͇��>��,K��oR&�X�%��އ��5����e����m9ı,Ow�ԉ��%�bs=�fӑ,K��}�H��bX�'~�}M�"TȖ'����Xvz715�����oq�������r%�bX�﷩q,z����Uڦ����]�6��bX��m���D�&?m�ӵ
� 3Y�.��ND�,K���"n%�bX��]�6��bX�'���D�K��EdO��߳iȖ%�bw��3?S.Ʉ.���5"n%�bX��]�6��bX�'���D�Kı9��iȖ%�b{�ޤMı,K����p����>6�55۩Y��'di[��n��Y7"�v�cv��6u�J){�w��X�%���z�7ı,Ng���r%�bX�﷩��L�bX����N�D�&<u`EUڋ� �J�&2%�bX��wٴ�Kı=�oR&�X�%�ߵ�SiȖ%�b{�ޤMı,K����,�kT�a��ֳiȖ%�b{�ޤMı,K�k��ӑ,(C"dO���H��bX�'��߳iȖ%�`���dִSX]k.]kR&�X�%�ߵ�SiȖ%�b{�ޤMı,K���6��bXGb'���]���7ı,N{��r�֊hɬ�S35M�"X�%���z�7ı,Ng���r%�bX�﷩q,K���充�Kı=�oQH�/mmմ��vn��E�@M�43K����fGd�0��;=���7ı,Ng���r%�bX�﷩q,K���充�Kı=�oR&�X�%���粗2k!&k5eֳiȖ%�b{�ޤM��ș�����m9ı,O���H��bX�'3��m9�S"X������ˆ�d��Z�sR&�X�%���ߩ��Kı=�oR&�X�a�2'��߳iȖ%�b~���D�Kı/>/s�e�����{���oq���}���Mı,K���6��bX�'���D�Kı;���m9ı,N��ٹ�j��,�s3V&�X�%���}�ND�,K�{�5"r%�bX����ND�,K�׵bn%�bX�6(1 �� "
�����U�3QA��R��uC1z�n��G*�"�1� �̕��Й�ڵ�6hV�YU���՞�Y^:!���j�%�aihwls�v�c���q]�����tf�u�E��2҅� �/\1�1���6d�(`E�ew'n�l$zk(���=y�ۈlv��eUv-��nkY�mPs:�nz����Gj��B�]�C��q#�v�Ȯ�������f�6�r�����AV�9,Á�^������è�A筮��7nzc��j=ߛ�o%��~ޤMı,K�k��ӑ,K��u�X��bX�'3��m9�q����w}f+��)������rfTȝ��fӑ3*dLʞ������3*dO���ͧ"fTș�=�sR'9S"fTș��L��Jhɬ�S35l�r&eL��S�ߵbs�2&eL��{~���Lʙ2���jD�*dLʙ���l�r&eL��S�ߵ��rL5a����ֵbs�2&eL��{~���Lʙ2���jD�*dLʙ���l�r&eL��Mj��~�R'9S"fT��u�7�6F`8���3��6��y��=�sR'9S"fT�����?[6�D̩�3*~��jD�*dLʙ���3����{��S��p~}�ڤJ���p��������K]:���ݒ'b���r=9��{�����r��{�?5�[6���S"fT�}�H��L��S"}�ߦm92�D̩����9ʙOs������[��J�����*dLʞ﹩��'�b��H�"]Tȝ���3iș�2&eO���H��L��S"w�߭�ND̩�3*v>��HfkT�Yf[���9ʙ2�D�=�L�r&eL��S��5"s�2?�֪j'����m92�D̩�߹���;ܧ����}>?M��3��g绑3*dLʞ﹩���3*dN�[��iș�2&eOw�ԉ�Tș�2'���fӑ3*dL�9�e=��֊]K�e˭jD�*dLʙ���l�r&eL��O�{�ڑ>��D̩�;���fӑ3*dLʞ﹩���3*dO����델���1�
�5m�C�Ӕ�K��]e��Rc�����Wm�fzz:�HY][6���S"fT�}�H��L��S"}�ߦm92�D̩����9ʙ2�D�u�[6���S"fT���j�S5a�����jD�*dLʙ���3i�W{����?�sR'9S"fTȟ�ks�ݧ"fTș�=�sR'9S"fT��{�Gf,M��8� ���y��1�feOw�ԉ�Tș�2'{��ٴ�L��?�0�&�q5�?~�5"s�2&eL�����6���S"fT��s=L�k!��ֳ%�H��L���j'��~�iș�2&eO���H��L��S"}�ߦm92�D̩����9ʙ2��q���~��p�%c����{���=�sR'9S"fTȟg��ND̩�3*{��Nr�D̩�;�o��9��{��S��?>�v�3���+!Nx���*������q�+Y#��]����[�������33Tղ̷35"}�L��S"w?o�ͧ"fTș�=�sR'9S"fTȝ��v���S"fT�}�H��L�����ﾟ>�3��g����S"fT�}�H��"���j%��k��n%�bX���z�7��,Nw]�����������N���8�H�o��IH��$����KT�<I%:d=�OHu�.��Z.����X����"k����rO{�_�rOw��ܝ@��A�B�����R�g��o����<y�(�NC@��� z������f�������q;W!�۪n�jME��s�t�%��WY��t�Dvz�{���|��ӻj���<���`��K z�~A���򵿖D�3
H؜4}�R�/YM�l��z�o�����+��7<Q'�H����|h�e4�S@��`�B<
i�V��Cn�v[0�ـ{�m,���\�8�=����8�$4�S@�ޕ-���=��h��fe�7^LRGQ�c݆�Ӏ�" G1b1��P���0C���5L�:5�hn�bµ��ף�u�탗8�Z�ι8��;0#����-ۛ�����˸�����usɱV�Ӌ���_v6-������rv�y�q�^-cVNC�MV���c�;�������{^lÝ�;^��u�ZR��]v,e�N�c��.���+{4����r&*��mI6W��W�Ys-�Tڶ��lj��M�ڮ��d����yKT����K z���L�D�A��|h�u,o"Ɉ�(6�Z�)�nˆ:\0޸�])��8�EZ�v���=�l��fȈ��f'<nߧ�Z�����=�X�6F`I#J��'K����'K��.]�Ց<�ǂ�6'�zT��ɉ�ff">�|x����`�T�� ��
�H�e@I�mN����� LG�A�D��;k1�K-�)+N�v\0	��n�� ���c�y�m�@����<̙��/*h��`���Tog����rO���g�1��R��W�uuUwfϯ���f�>�0o��@����'$@�)"jHh}�fy���|�����=�l��f 9��cxBb#J6�Z�)�{�)�^���v���f�Q(ɉ6�Cbk���	��T���83���y��]L�]~�����3wǋLC�)��[>4�S@��ՠ^���ƪ�&��	$i]��l�?m6��ـ{vٝ3	+[�dO#1ऍ��@���Z�k�s�Zn�$!���2Q�`��O$Ť��?mV��F�	�H��Lf�++
H:g�u��XD��$ *XB����BF�<ai�����DS�	#$`� ����`�&��X0*D�
�@"E� 0jD�"����,�)��7��M&�,���
�(Ĥ0��
�@�J�KIA��(T�� E%�,9U��q�]����*��H@ �"�����a+.2�f$��܉�,
����>@M�PB����HT yTx���qM�@<�tA����.1���}�p�ޘ�\0֎q������EU��`ݶ`]��"W���^ό��c�y�m�@��S@z��� ��0�bb=F������U�H�.Ӣ�J}�c.��WkV�vF��@�lfr��9�kS��o�����~�m`]��">���W��8�"�IRC@��ՠ^���Қ�)��WSȲb#J6�� ��0n�0阈K�_�w,�#���jT\"�Z�Uv`~������>�0�M��S1ϳ�{��+�*��.�ݥV`]� ��&'{>�x����=�l�?:6����B$"닒����K�i.h�����s�:�ݎ�r�{5���Ԓ��x)#bp�����/YM��M���;ֹ�(7<Q)%UZ��f}2���>�0�V��<�1"�ǟ=q�#Bi�hl�`�� �9:\0Ч"b�,�������0>���ϳ�λ� ��h�Jh�S+�� Y#�2Hh��X�ϳ��kw� ��0D��!�Ȅ
��	�i,�w{��=�{ۻ����֞kd��Ӻw���r����g��6:4��a��!N�#�S.w���4����	�nڣ��mq ]Oۆ9M띮c�g��rf�Z�8�{A��s����6���7��59[sBYk��ù2@]����|'`�� u�S��NP����t����l�r�&���W\�/��h٦Fi��zC�[��t�%i��H���������.��k� ��m=#B%;u�\���`�v�q�u;��m�\��c���3]*�Wk�����=�l��g�f" ��@�>�~�bɓ�D�4��Lt�`�p�'K���j+�'W@U��J��<ݳ ��هDLBM��{�O���$X�Hc�I4�n�� ��.�p�;Z����4I1��4�)�}�g��}��ﾟ�v� ��ռ�&Ȑ	ŉ���[�3H�s�q�\�sWR�=�X�g�����F��p�=��=�S@��ՠwYM���[�<q�nI7$��צ�^ʁ$EqC���w,���m�嬇WEݠVGd��?s�h����y�b]l��>�O�篝Y$Lc��ڑhy�0��q�kw� ��0�M����E���R'!�{�)�^���v����;�.H��x(ēxێ�g^v�H���K�vD]#��g���\V#~����sZ�0I�`8�i8~����?s�`]�陘��5�� ޤ���R����wj�Y�~�mgD�LDBG>�0n|h���g����y��s �8�ڻ0}|`��d��A3RLLݔ�;������u�F�<v`}3���`���=�`]� ��խ�a	8�$4�S@��""<�~�_�m��31���U���{=��n��J4�
v��uB��l�[�����wL��R�������	��ou� �.�|���(�m���e7�3�H�gƁ�}>4}�M���a2cQH�� ��l�<ݳ�R�w� �_��)�U@U��J��陈�f"��~�nI�~��ܓ���7#��0� �,b��@`+q�T:���3��Jh^�ōd����N�����8������0Z}�`9 �=n����Jgh�st�WE�+I2��,�Z$�����=�w�	��Ĳ�gi�����w}�;f ��0�M���"�2G<�x6�{�)�^���v����;���L!#�**����`��X""b>�������/�O�@���\dqbP�6ӑh�Ȱ	��ou� ��X�|⫸(�m��z�hy��n�~�g��rNw=�'�1XD
��c������������jj��-�}�\�v]��7g�L�L�IH�r���0�s%q�@�ٍ�"��GMї��[�v�qˣ;f��y'%�I$Z������X��i���N��חr[�`W&�wF]�zK�%�8��.���Á;����3��`mN
紅�G�8����ا%̭�h�t�%%;�+=2��t�L/�V㳌i(5�j��v@f�`��w�mTQ��;3��*�`���bkmu�<�X�٭pg��V�0=�]��s�.��Eo����Ɓyڴ}�M���?wF��$�0R4�4�տ�y��|h_�Ɓ��)��[�ōd������޸`�� �ˆ9Ȱ֎��ndG#��/YM��S@z�0��`x�vQusv�I�0�`�� �9:\06�ￏ��6�yq[/��h&�sl=��:8Z�����;�D����<�Wk z��� ��:f �O��󌌂P�6Ԑ�?s�og��DTDLQݗ���,��0����H�9m���e4y�Zg�w�O����hG��L��R'!�����o�����m� �v���j��O#�#MŠ{l�����@��� ��uȦH�j(�G���v���q���G�M��-��7"d��<̉���ƲA�H�p�����;�� �}אH�`v�t�X�Ռ#�H�4��>�[e4{�3�;x�vM��ݢ�����<�`{�����X���E%N�D�9���o/|���t�Ŭ��nE�{l�����@�?LS����#�.�IYuuT���=�E�N���X�p�=[*e����\�(��y}���"�N���]e��"8�q����1յ8�"� �.s�	��nˆ%>sb�1�(�NC@��j߳3ď���@��|h�����4Y�&��m��6K��.t�`�E�lu�ȱ��H�p���<]�oƁo��7$�������+u:��g��i�}���72#�H�4�p�7\� �.�`oF���3v:l���;[�Ψ�\H�n����:�8��<�ζ���Kz�!��͏z�X��`�}31�}|`�|1̋$x�ƛ�h�)�{��;����S@���\d��$lR��=�l�7]�����z��7���;=|��F!��p�;��@��p�6K��.Jk�!R��c�j�]��7e� �.�`�E�N�,hs��zo80#��=�@>�ȁ����U44C�!�x�1H�DX��+i,h�����"@#�U�,D��%�⸭P�#��7���� ��)m)����%�Qy��8u�
o)>�=��m60���rzCP�0�~��((��؁�(K�������y�O�W��@H $i��h\�ɹn�
�7���SK�m���n��F���s�q�۬p�7LѦ�����v1�س��nj0��!lm2�Ksq�������n7_8>JsۨH$��e6>+�m:�N�\��h�� �n5;�6�";�n��%U(�B&�P9�n�V��T����lX`4��I�mqJM�Z��Ut���b����n,;7�����ځ�c�>
���bM�&�\z�B��m
cO-l�u���ԹZ�fduUV�$6���琜���A�s��06�ل�&�c�q��ݜ�;����[k%��'n��tZ���Q���sB]Eӱ/E �,���/.�r���e5��v���8��s�V� ]����Yر����N�]�V�U�&fu$�r)�
�MN�ٓn�l�S�h��n�M-�N�t�˝aj�i���s�u�	f8�6�I���׶���ILt�{M�:ѯ-����	-=�V�\n�&��½k��lp�K���;v��)d�i�Q��閦nT�Q�:>r�eC��N��e8��	%�*�|r�g]A�[�r6�a�� n�:��)c ���u+����8�:���9XKˣFvٮ�m�����t��n���9�c��+[���Mmq�u1ӯ.n���P�e%���I�� ]@#��-m�8"����nƺ]�*��pX^�ޚI"k�&���6$S(i�)�(rF^�:fj�3V�.F�������sQ�TP����RBJ��Fn�q������PWk��+H�9���q��Ny۠�9yk:�����'m���u�k�đ����0u���%81;XǦ�w��n��2[���h�z�-d���^��ö��U�-���m�r ++u܆�pV̀����t$�ڗb�j�
U�`0� +��-�q�[L�m�;�����<�WcE#t]���¢�P9�������C �E <	����|�c����P�/�&�(���N�Mh���]3Z�]�=t��$,U��#H��M,�L��K��+�-�u��fK�A��i�����B�v1�{6n�ڍf�v����̝Oc�.���R�E��{^q"�3�����ٍ�Ouv@lEv��y��`��sv�cJu�6�6N�{s�n\�.�-��3�/�к���pb�m�u���hu�r��ݦ�l;U�����mN*�b�������u��|�N'f܆�gf��i32j&6�gN�.n�7(����]�BRk=����?|����N��}?��l����]�u�h֩d2,pxb�6�4}��������`�|`nٟD��BGs�~��9��jE!�Z��h�e0�&"&��� ��� ~d'�J.���t4�`��l�v\0?������[>�h��s"�8�$47l�>�������r�=�l�7��{�[W�h�U�֨�vw8��ڶ��ǰW�MC�X{N̓WX�L��L՘θ`�E�vˆ�\0�|���	�r4��4�j՝癙��Ɉ��bbbm�|`�|`{lϢ%"����)��E$Z���{l���t����Z��׋�!�C�]%V~�3��D�S���v�X]K!�c����N���Ȱt�`%� �u���Ez��Z�{<��ڐE�Ӗs]7^���b���J��i"gP�s�#5)>�~�M���� �vΉ����u�o���G!�!��Z�l����\0�"�6P>����]�v鷭jnI���M�>����^!�O!H�C�D
�Q ��٭��9����WY1�(FF�$4?��<v����;����ـy�f �լ�줮(��TUU��6��b'�Z�?���{�Jhuu�$���,L�`�EӪ��Q:M/c�����g<>�8��]������qE"�/�{��������Z���Y�!�,qH�p�<ݳ>�����n����~�l�*�Y���p�=��;��@��S@��M�x��F��D7�����M�r�<���<ݳ ��
s���P�}�nnI����Y�H�<qh��h�)�{�Jh�ՠU�+�c���9�:	�L%>H����n�rV��*H�qI�b��ȲG�A�$4m��=��4�j�=��j�Sq�N�ul��wf���Ȱl�`%� ���c��1�F�ۆ���Z�l��fy癘�}���;���:��p)���Ewk �ˆ�\0޸`�E�{�:9��LKN18h����)�Ow=�'>��7$ҿ�x	V#kߟ�����D��C�/m��e�U�g*p+I���[�+�ɒf2���c�4�'B���t������A�6�-oOL��VR�m.'�8x���n���/%ѥ3��q�ł6�w�1���o�q�X�;��L.���osͧ�9��>-�p�j�t�����%�7T�� ���\��H��l�k�+mn��PD儶Y
xq5:�Yv4kZ�.��Ԓ���E��$��tԶ� $� ��l���[����>���'c�9BvF����n�l���o�����a�Nr,�.�p�;].�۞8�q���yڴ��M���=��4�V+���C$Bi8�l�`�� ��9Ȱ�2���YRC@�e4}�M�h/{���9_�o�Lx9�MIw��"�=��N����aq�t Fz�)�Jpc5��(��b�C��ѳ�V؋�rYק:�r���"�=��N�w��])p�C5uu��j�IϽ�M��C�"b'���޿��6�۷N���&%�'�4�S@��S@��Z��Y����{��"�=��N����vF��ē��Hh��@�������>4{�4��Zɐi� �QbHS�W"\�f+nGN�J �I�"�%�^^�-덼��$Bi8��e4�S@�����:�Y�RK]�E�Z���T���9��{vـ=���]� ��cu�A��RC@��S@��Zz� �;����|��3;��ߧƁoJhQ����Ibn�s�`�"�'K����.����f8��I����@�e4{�4�ՠw���c�7���ێ��J�V���\:鵥�H�����,Pq�$ı���@�e4{�4�ՠ~�j�=���dX���$M8h�Jh��@��ՠ^��z� �s�N7	!�^v��;V�z�h�Jh��R��7<�	�R�X1+���ϯ�۶�P:XH�!$$D�H�T��1N�b�_�����'���HH�Ǎ�"�/YM��M�6��M�陉�����iEXR���n�˥�iP�b�j��:k1�f{:�.��������@��5$=���4�ՠ~�j�/YM��2��-�&��'9�r,t�`�p�:�u�,S#1��H���Z�)�{�)�^v������LKN1���S@��S@��Z�v��:��E�#ŊH�p�=��.�k �����f�/�蘘&b&C�w�����p�1E��f*�,���N
A�ǳ���%mDX�����[vE泌ca�$
i��2;��:z*"��Q`ˤ��[�ֺK��B݄P�;��Ϯ�n�mr���s���$R����[����������7+:�5�\g)��>�t���M��UE��!)����3�`u����C�]�2�卵 �C�{+�óXL��5���5u��-�_�;?���Vg���(Y٠���5�b:/����i��h����9~Ve��3Wvm�v��,ަ� ��0n�0�QJ����D&�Ӌ@��ՠ^���Қ�j��H�x_���G�<I]��_�m��m`��X����@��5$4?�3����Ɓλ��i����gB|Q�e[i�(�ۆ�yڴ�l������@��S@yԺ�#��P��B��G%���d�f��ָ3��+F�ήL�"dF8��I�=�H{Ӎ���z�������h���n-�צ��A(�*~�4���w���~�mg$oR���4�u��@��Z�v����;ו��H��Hh��@��ՠ{l���t����+�7<�
�)U���k ���?���?�Ͷ�o���s�P;u���j��hs�3d�u`[�íq�z��ӽ���E<ۦۻX�p�7��w9�r-���뉠rF�$4{�5bF�6��M���3�a �;��V�Qv��*� n���i���`�	��XC�X@�Īi�@�: f&�O� B`=T���1h����0 Z�:Ņ�mA�_ �B#`HH���Ā��v��p�@��ֆ�o��,��Q��>��-�)�$���G��t9� �H�����P�����LV
20�ڝb����L�7��f`�����;/�FT	8i A��
�EZ1HT��b01�"Q(u<'�4Ş��;Aj�PQ�L4�UiH:�P4�T>8��4A�z ��T~��w�����O�����⺹!"��j�ڻ���3������|h�Jh��@��K1�MBQV�誵�=v�鈍o8�:�Z�v� ��uȦHڑ�)�I���b���\��8ӝ��i-�ɬ:&�r]#���,�`��D�{�)�^v��;W�f~A��|h�|��q����rI�6��M��`ݶgL�D�3ToZ��QuW7hT�J�`��� �e4{�4�ՠu�����8��Z��h�Jh�ա�`��@	"�(R%E)��#��~��w$�~��g�W,����Wv`ݶ`33-�r��w,�e4��LsQ�D� �Q8L���d�E�w4Ji�K�=�%�n�:j���mSCd�<I�@�v��;V���Қ���H���R)"�?s�gD��G>�0n���k>���k��9���,q8���>�O���M�h�ڴkV�E�IN�۶��6��M����&"+����}^?��	�$��/;V��i��=v�۶���&&`�&��@�	������I��\�kZ�X69�42�n9αut$�T^:�r���d�eɅ˽�F�
�U�a�ۄy9�&�f�n�K��ǿ��t�;��U�����=���[����n��n��Wc�Mó��lUƒ�a构3�Mp�m�a�[][�e�s'V�=��/5pc+�h3���dV�VtkA�zclmX(*vYc�!=���f�k�bA]��B�73"�����[�k.Y�]f��e���j]�qb������D�R؎�Y۳D��p����M!��>����z�h�Jh��@��%)�cY#�6܋@z�����:�X�����뉠ncQ�����t��yڴ�D�^uܰ}|`��.եT]��'�h�ڴ�SC�3�]n�h᯾1""#QH��@��ՠ^���Қ�j�;���J!��d�խ��fKZX���D�7��z]�.록8bɍI1�M	c��7�z�h�Jh��@��ՠ^e�őd�!u�\���'��7���ZJ3ʞ;�N5�L�}��;��-���?.-�����N'	!�^���v����=��?u�,Ojy"Hm�@��ՠ^���Қ�)�_��o�I�d�qUUv�ϯ�����s�� ����6ߟ�����B��i*�q@viWsN���6�-�݂��Ma2�Й�:���&�cQ�����t��z�h�ڴ�S@.UYp�@l�G�8h����i��=v�۶��H|R�!B��QV�]��0:�X�l�����"��(�h ��}�~��~��~���ޖc����n-V�M��M���?s�h�lqdY ��wj�Y�{vـtDG>�?�]� {e4{�4�di��! %2b$�.��fs�V4��[�A4ϱh�P%�.�өn�q8I���?s�h����t����W���H��cN�v����=��/YM�r�*�1���nE�^���Қ�)�~�j�=]��SMs�5$4{�7$�}�M�9�����-}�7�g�9d���*��G 6H�Ĝ4���>����w�}�m���߷��v.	�<V6s$�"�q=uF�p3���n�Q�l��9�Ύ���8�1)������=�S@��S@��];���J��ln��\0��;��������H����"��6�4�|h�S@��ՠ{l���gu�����N'	!�wYM��k �v��&��`��DUҹ�B�EUY�~�m`L��g���u�0�3�&	��P���躵$ن�VQ�;��j;3b1��8L��1Qjx�A��B�J\�R�'��^}�������tZn����{曁�F導Nm�5�|�'<�u�A1��Ҽ�g��v\�@S�4�w<�-ƍ5l���67*��k�k�έ��NT�i�9�ѣ�=���4Uh^!�/\hQ�HVQ��ZA�M�OdzmOLH��<��Q"T?"}~���<�<���i��gP���˯#1�%����u�զ��D�uru<�*�����۶�u�?�1��w,U��&� �hrC@��S@�����L�˨�.�¨�WVU]�uܰ�M�>����K{�������X�X�E$Z�r,d�`�p�;�� ���e����8�cqh�)�g�����-�|h�ڴՊ��H�Si&��@tnxn6#�uS�&�|x��Ε:�hC�����-#��F������|h�S@����y��}���=Yo��	$�p��ܓ��z���+fA@"� �!@-a�A | �\����w!�Y�{�)�~���D�"4;X����t�Z��7���9G�d��H�Ǎ�"�=�S@��S@�v���*�i�rF�wf���\0s�`%� �����S�	A;z�L��U�B5�U�O`�u2c=j�7^��'\?���N��ke�[���O���=�E�l�{����X�A,qE"r�v��e4{�4�)�~����48%�*�*�`nـ{vه�0�IM�6"��W����@K~���7!�?y�c���RFӆ��tf�M���k艅������s$X���Hh�ՠ~�j�=�S@��S@=:��23�8������Vr-v�[8uc��	��t�r/	������wK�[Y�H�q~���h�)�{�)�w;V��7�d��E6��`nٟL�LADD$kw� �w-�;V����6�9�C����v�XtLLz�:�X�_ �C��*��]BUfD����3ݟ|�I����w$��צ�Ъ�v���c�&aDG��~0�N�P�]�EZ�v�ـ{�� �.�\0�"�7�/����v���az뗳mq��B����e��u�2f�<�]-N�&l�%U���0n�0�l�f"'蘉�|����Q~�qcY#X
H�p�=��;��@��ՠ{l��$z����G$PĜNC@����?s�h�)�{�)�~�Uv5�9�PXӋC�<ȕ�}� ��� ���M�r�C���$Ʋ(8��Z��h��������'���RM���ܓ�EEE�EEE�QQQ_��QQZ�����**+��TTW��TTW�Q@C��TTV " ��EEE��tTTW�����**+QQQ_�TTW�訨�������EEE�*����**+����Ȩ����(+$�k!և��1�0
 ?��d��-��    @  �               |z�H@P  P 	�
H�*B�RT��( ��*�*�D @E$U �    U(`   �
 �	$ 
1 �����{�^f�e�gO�ϗ{S{�@��,g�������뷹��K  ��{�}�>����i�o�����+A��R���=o}�_[����{o{:K����O��O.�eͥ�����/� ;�*���(((2 �}�����m��ީ�����m��{�A�2�;��=�j����{}�������o����m�kϷS������ ���������]>�:^�N�w ��+��  �  H;mťW � @  (b ��Vۓ�uͺ��ǹ׮�a�� 
���.�u}�ū�N{^���ԫ �u��r}���f� -\Y�{o}�OUx }9����K}n�]�������eo �t�[�]�����|���y�W��x�
 @ �a�=��������{��{m[�t�� �>�W�NZ}z{�x q(�� �4�v NP  P.� -��  u� D� 1M�  +�#�� �	� h �  (P � �  P� :q� � f
 �{ 1  H�n�}t�� �=+�o{yo}�^� ��Ը�C�� �{����;����)��=Ϊ���y_O'�g��^�w�v���:o ORdm)J@  O�FQ�J�   <z�R��MF��Ob�Ry)�� h�BFJR�  ""CRR(��Fj|	�O�����?�����S���G���Q�d��Q� ?�(����Q���*+ PT��??�`T0�LB�V�?��@� Q�SR&�u!L4M�Mc\t�BA+�Jc������C#������0H�
�	C�ѡ�����aa2����%텣
d)�(Bb� �K����D�)��@��Y!���dn\�'����#LB4qcL�V!qԉS#\��>�#^{�3����������R#E��b�``I� � "�H��ň4�ƄR$B������a4!QĐ��ĩ�@�Mcq&��`0�H�����@�8�J&�ĪA(0�.2� c0((b�#�Ǟzy���s|�������@��T5#\)���=��.o��鞕5 @��º:�[�F	 �)���r寇�
�&X �_RA��
t��g��>FfL62%B�Q�� F� ��L-�C1`AdHH��1�4�!�~�H0P��<�;0�;^��E�S�����<�lI)����i,�f�C���!���+HJ���xƉ��$V�<��SB@b�!u!t�o�,2�o��<7p�s����жa��?�~q|2 V% f�wl)CшH)�0�F�`4fOC�6�bHH� ���$~||�zd3y��F�hK�{�r�iXZ�F�����̆B�%�ڑ)Hc.2��&Y~���g,��\p����e}���c�;wn�$%CJ��1J�B�JB�
��V)�PtX�� @��\)D1`�<������4#D�F5��6�$<�Ot�{��p!s�{�}�o3xp�_=�������.pB< �pX�G�I���s&B��)
�I�7���)
\�%%2��a2`H> >=0!\M)xyYi� B	"���#��ȱ�x)������K��C�����f0�B��
`����#�i��L5��>���.k(K̸p��8`D i�xRRy=�/5��x=��^\�\�p���Ig����H�>|�4��xz��/��V#M<���H�nr��s}��,2>JK'���Sx'��F��b@���!j�k'<<&�	/<a�˙M����<ĉ��
V���ĥ���t�ā<XC�wq��	LS!p�8˄�2�������3V09�K�rf�9���=@��3�NzJ��<��8^g�76]���r��i6xJ��>ny���r�S�**��o��P�{�O�U��v�~�&����᯾Ly��=|B\p"u]n|�*�r��|�N<�k�YT"������\s��:wB��|'y�TQ9X�y�M������{
S	�5�'XS�	]�h��ǡ���:�C�� ��0Ӈ��H����#sNy}��`��0!�#[��zzbB� c�<#L]H�04 Q�F��"����RR\�#HU�X��(D ���V�B�B\�j|0c�PЁP�D���MӞ�8�y���aQ�P��%�y
��i�.r�^d�'��}���ᄤ��$+�T�o$��2sD�1�0�˔p�!W%�S<�L<< T�9�=�I��g١+(��xĜ=�ĈP�AS�T�B@��C\҄)ru�>��Kv528�VO������������.�!�w�7�xOf�B���t�%e��)XGS!W-�'2��<_w����L.� <Yw]��R�\z-
W*��<<!�B�a/�}Ἶ�>�$����<�|�_��T�v-@���!\6�þ��F)H��|���{�9ĈbEX1�E� `b����<繡hK�Ï���eY}�Ynj����E�����d&\�3�[��Z��
IhbT��!aR%T�M�aR�4J��T���\Y���8�)���=�j@��=�>���T�@���c�!R��I��a��=1�=����7��Ē����@���&rb�&�
a���|�p��}���x�朷ZxB�'�!/̲��{�Bc��3!��L���h��00�JR����(a�p"A"e�o�8�<S{9��{s>�.y���:m<cX`L*���F���T4��9��'<��3ЋzŇ����|ǥ0`B5"� P)�����]�C�V$}#�|�!p��`�H���$��!J�L�����F��>"�S0YbƄD��C�OSW�W���0 �3�LeWB<��L���6-l�o<3y�@��0���N:j�X�R�%8z{
f�	�y�����Hd1�$F=��d�>�8{+�X>�
oz�2������g��� �T�;�O�/i!P�s� ��@"1+�A�B��"D������:��x|z��)���d.��'���C�vxK3^�A!���|�N/�Ja��¾�
�w�ݹ��k�x�Bo��ˆ�=�*�jŦ3y眹||(*��HD�1�
<Ha��8>$)��p ��N�E�`�<ɜ�>�`V���yą1�8��O}���^	�_<<�sN)�x��$��}B
��9�o<�>��3}>ዠDa�A��J����`���G�]��������
�0�#>�)�*cÈƘhq�>��8Cn �
0X`B�D!��H:�!B4e)�@Hk�%XhJfL$�``ȑ!����i�&�a�	���Yk�	L�D)�ɗ������1Ѝ��X�ELڒ�qa3��yŅ/0�'3xRHR�S80��"I��0�M���V%�g\�FjB�2�o&�Bg92SJ�#n8L�2./"�va�}�i����2|T�HP )T�Q�u�@�Lܤ�h$K06i)���������!NK,�8bJdݐ�������������
ld)��B,+��ޜ4�����0&�9>`B��_'����+���I*l	����w�᧤
a�#!�@�
0��T�	i�L5	&d4!@�W[l�(�J�h`���E�B AJ��hE�� 1(@��&� @(`k�A"H�A���|�d��ЀU���$�Q>�OP�2"eY�K@�|�b��ji-)�pcׇ ��`W4�0$)�'�����< S?���=_B	CadD� ���.�хq�^1��¬d�Ԇ.�3	�du� ����
��K�$��K��'"@����V{���Ո�X�XW�41�@����4���i�(I!��˃a�aRB�`k�B��5�1ؔ�CW�F�k�"��GX�0��NbG�c���H��z>��aϫ�}�����d�>t$����YVW,vہn��y��D���<����$@�c%���ibէƒw�>'`�8LW�u��x$B�B��D �Ή.c�b�6WM.%:"B�_�(z��X�O<-�`�r�h¬�=�B4d�#C�b�JB��1(8B�LSB���:�Sq	k
XW	s��qIf+��a��#�~!�M8&)-r@���,��S �2l4I7C%�����0du�c	�����F!��X�Y$���Y#L$f`B|�)f��)l+H�0!G+
Ƥ	ňb���/��	�>�{�����!4!y	"�G#db��A��j��cI�t�{������m�� 6�  � m��`L�n�[v$��+;-�eT����mE�lְgj�`�n4��UUT5���	C�m��[F�H Z�4�16���WIi�pkqZ/,H� 9�r�Ojn���й[��v����6��:pq��M����]� rD� m���vZ�j�Ɓ:65���l:�MZ���A��NȵR� �ǜ5U�UT�*�PJ�UU��%]mN�C�������m$��d����9��
  [vݍ�Vԡm�@$6گ���d��     [x [%��oVך�d��8H�KG)gI4PmU/'m�y�9�1��T ��cZ�l�ݻM�o[z����	a�   $�i��/i �f۰m�e��I��}��,kV� jrUM��h2I�n��f� m���ֲ�8 �cl� 	��{i $$&F���� �     ��mrI�-� ۰ m��ˮknZ���  ���J�׭�����$po�~���m� 6�   I�� �$Pf��	-���  մ�m �[� $�k����Zչ�l� l���}�|6�`Am�l �l�oPsm�A�}�Ҩ��t��V�U� �lޠ�n�i��$K.YC�Ę�	 @� ��nݰ�kh  j�!��9�H kn�� �&��.�  $�` �l��#v�Z�  6�tH��	$9��[u��9�$ �Um�Ie����,��Vv�m��� m� ��n6�Jm�� ��[V�p ��m�e�6��6��*�]�P�%
3U�WV7R��@l�t��Ͷ ۶�j� 	-�[dp-��$�o6ݸ	��gI�pͺ�  ��u7U��-�i��mm�j���b���)�4����C=���B�)�#q���\/Zs�ڶ[�kn  �]6�8��d�/'�(�V���UU��+�� ���  6�HN8w ��)�K�%���uN���`���m��� ��	��at�f�G`H/-�,9�ձ�mp	���v!K[77]M����J��#�ki6 m��� �e�mm�p� q�Wj���
KeUb��8J��-c��p����h H�p	�����m6ؐ��_H�ėm�� ��v�/F�/��;F�.��7t���o�#e���� ��v�E��J m��g&װ $/m��F�w�n���*s�۪���Q��豕sԫ$�UU.z9@���6�]5�d� ���^�z[����'d(]d�h���<ݪ�8�',�	zkܱ+�D�4�zj�T�F���TZ6��l�(<ԩR;V�u���P:��3b���R����m�3Uz�q�c��`!oQ�6���8Ӷ*���m�R��v3@a��狕jUƶ.�8�4���1Tuzx�U=!Nl�8
U�����	;]�I0�/I[hF�ʵ�'r[:[,�.cv  Y�᭑�M���V�R�PR�U=���@P��iM�a� $*m���}6�l�v�Hn�)I	n�K�J�mA��s4�WR�P��MmHK(�� 	�������J��R�D���=UTacp�0KU@Ql�9�8�n��� R�N��!À�c���^ѭ��9#'Y�emFݱm����5�[� m���j�2���[�$m�'-���޶v��d��Z�TjU��'�����p6�l�`ֱ�v��-�������g�W\���{�<��V�t�H  �� $�`8HH�6�j���� .:��;�� �M&m��(���a��-� p�$ݶ6�fݒ��L��Mh�@�im8 m� �׫	8U��kj��(  ��H-� ��   p   9m�m�������m1�� �R ���   �` ����UUJ�R �**���  -�� ��M� ����]ɯI�jHm"��-� �t�(���m�bI�%0[�^��~����p�iB��gckb �MhW��܆��{-���nr�Z�/;�3��6���T��l�`���pS��8  A������f  �V��@  �ۭ�oY� @Nؓ�/Kl���  L��U8�Z�ݭ������@ 6�6�' V1@ mV�4�UcU*�JN��.�]�1�W�]����5l[�=�
�h�hxfU�z�q�m��kd�S`��:�� m[Hv۠(݂;�V����M,f�h�  zA$���L[Ce�  8($  �m��uR�m9ldKKu  -�'@�`	 �� $m��  �-������|2��Ja�J��k�M�ڀ�>��� ��9m��A�j�-�Ԫ��U� �e�d�6� !!�$n �ζ�@   �Œ�dX�H[Z��m��\��� p��H � �`�i. l  ��  ���.�m� HHH"Z d��N��]6�I0��lH��� mJ�!��ut9m��R���� $� 6�l6ٷlm&� ��`8�-"ɲV�*��Je5�k !�ըr�Pm:�PS�,�9� �*�^^�I��3
�[q� ��`   ��6�-� �k�m����� � ��ce�i��H�m�: ���j���!Ć�d�\m[�3��m�� �8-����-������_���m��`p�`    H  t]n �v�#�f�Ɗ��m� ��z;8Zl�����[+�5UHMR���m-ִ��m�8H�  ���Lٶ m�m�  �۶�Z��Fx�]��� �,�@5�G�)I���-�g�V�YF�V��ͩW���jk�` ��V��ڃWV����[/Uն�J:�S6ԫ�Un��VU��[k/.ꪪ�`@9��@kX�-�I9mp��č��$�K�[�mImHi�lm��mJN��4�UUԪSb��^���m���:� �l�      m�r�I�  HK(�    m�8pm[X@]���1*�*�UT wm�f�޳�H٢������$�6� �����	:������e8��[j��T�RdX�:�rY[e� �Z��d�%��[�6���[koa:>��j������tZ�KB���� �28&U������m� 5�qUPH�$��Ā�M!���v��M$k��G9K' ��`��7R��` ^���C�X�R�cfp[KM���m�l��#�۷6�*Vj�ꪑ��IoS`�b�I#  �6�m�v�[��Ӌ�,t�T�[q�.ӷg`�C��:o^�^u�%-�e�Lմ�-��{T��� A�I�m��h�$!��3���t]-ת l �v z��v���ۜ�n��m�m�ɵŵ�aŴ Ö�4P6�l  H6�@   � :�l��p ݶ85����Y��� ��� ��i$�-� ���Ԙ[C���ٴ�@ ������ۀ s�H ���vH� �/T��(浀��i�D�       v�V�h2h�c� �     �6�5�(s�m���T�[@r@ 㜶�I�L� h,׳l$�Z8h �@ � iÁ�  .���u� � �䄀�r۶�9# �� a�8m�FݰԖ� H $�@|#�m�[� �v� l�@�F@�6�#�M� H�`[_k�����q"@m��ڐ��`m�   -��m����m�������l�[N��.ٶ�ݢ�  �@ m�-�����$�H	$� m�Ā$��p  �kM�� $  �� kZ� pH�v  ���` 4P �d��8]��4� A������ـ%�7I�����񭙣kj�Y&����8p� ���ڶ���Z.�I f��kk��`  m�Cm�� ��m�BYն�/ZD��j�` [G -�[GUW*�և��ڈ�0[[m����qу͔[/,d"^TЄ4 S�
� [l��������v*��N���E�)T��l-�}rv��\��  l��սڀڶ�z��+R� jU@�����8 6�mkV�� ��  �>�f� 5]nl�,t��5�gY·��www���&��� ��@'A����Z�~@"�HT��_Ȝ�E#�:��"�SĊ`ux��NU��� (��=����
�b���OAz*8��5 � q(�����>/��|)
 u<�A�S�U@���>(�h�!�A���P:��!�� Ep���=> ��+�"}�E����T�Q���O��|(�U���=P>A�RC��@� 	T�xTE>:"�>�4D� ���A=x#O}U*�xb!� �	D� BH`�d!A�]9�A�^(6���`����>PC�'}�(��:�A
��t�8
���|(*=T~���TO��:���X$�� @��P�E�D�`��,V$R1�U>D= �Q}A�D膈C�6*�YE����ʄ�_� �P�LQR(/�p#����$CTA��q:"�>���j"����Z�b&�8�@P�T�=�"��D�Q>��b�������1�*s��.��1m�P�'<��bk��p1�vm��g��uA����Net2�s�L蛒M�+�4�v����q,�`HC�@��ыpn��O���L�Un�u�W[pnv�s�<��`�g�NeL�l��JkшZmWS�+�G�l��nD�Я��jWj�'-\v��PƔ ���s��8�-��^s��Zm�� �#���#�r�n���5�u���B0����n���)D�3�u�zsi��b�G++[g�����5�v�2m���ˊ�<�͞8�m9,ݫ�n�E���mn{����x�!HJq�m��'@.�m�:���Z����T�c��ʲ�شu�t�� H�"D7g@%���:����ő���WJ��bv����C�79��*g:Ps�'Q�<�]��	�T���uZ�U�9^���{d�8���tm@u6�
`0I��2�]nH��� y��k�)ӥ� �ll�8�����koq��
�t��`UU'99�R\P̒g�^Xέ���x�I�Ik��5�2`AWnP�gvƌv�x�2���/���M�����i6In����nJf�v:r���j����wU�,[c m�Cj�"US��n�Hk8�n^��jU���VU�W����kSs��l�TXF�tsu�q��h���L�	�v�v#��sx�Y:v�&�R��A��J���O$�V���Zb�$;c��|2l�/h�'��6̦�,
v��㌹�kMk8�ә��x�^�m�ˋ���
�d�e�e�/�M�v2m��:���W	�$i���*wce��vW7!\�S��6[HJ�烰��T#���2+���@M��)H$QںLCF��Ѷ۵G0��ܨ7)�I4[�ځ�8N���0��'XX��ܬK��G0�RrG-�3Bk�;Eu(�II8�dq�S:�v�\s��Y���ZW�X��;l����`8	$f�m�Lk�qP �����A���	�P5�OG|���?|/���tR��M��%�)s4�vm��"�-��d	����@n\����h����ѷg9L���Nȝ�����&�����D��w�ۭ�-�k�'���ր����nZ�2��L��ns��ۍ:�7�q�N�N莔w��49����$��Ge9��mN�ґ�V^r6���,#�:b%s2��nj��v7i�s���d77v��4AGE�q�,r���9�����v��Ȼ���ݐU����!�h}Q¡�ݺ�w�f?�������f�w���n4�GI*�;���(�S'�wy`f:����j�޽�m)J��q(ܖ��ɥ���u`��9�V��&5 �(�ukފ�	%|`����{j���cY�JRln�(�,�۫ �L������ܐ�9��柗�#v�������ZƎGlm�)��:�(��k���%D75*E�)*�9��`�Sފ�	%|`[���H�	n�����y��y�z(B 1@ ,"	����
"��$�jB��%�~��6�X|�X����"��l��%������ͺ�wvX7vX�֚w@�mLY�P��W��Z�m���EF7u'pq�N��$�`��m���EF��0=� ��w�pX�i���[��,ox�;�9�6��G(�u�Y�#uGB��*�R�Q�,��,�&�fmՀs����=[�Ԅ���Ԙ�T`I+� �L����cY�JRm�ԥ����u`���b	 EDbc������&�t{��TԩRD�� �mL������I_�-��5�-Դ�I�vژ�T`I+� �we��ﲙ�I�߾:��&���W��s�ݾ��ns�N��F*H�^!\���+DRS���#����36��9��`��`w7Zi�q�EJ8X%|`���vژ�T`vZf��ӧQ�J�wvX]�v;�K�ݺ�3�h[JR��*�ƛrX�7���e��7jßD�!AR��8����<��|
��fw���հq	���RD�V;�K�ݺ�w6X]�v�ܭG��i�r��������+����Ļ�����[;׋�\�
9JR��lJ�8p�z��9�u`{�nv���:���|z�'9R���#R�ĸ�;�S��q��EF{�u`f�nա��	���`w�u0;����|`����[�ZY�	JQ���<��~,�z��9��`w�uX��5p�h�((�`w��V�%>ǵ�39�6}���1)xAp��D��?)��`��on���~s����)s�βq]Tu�L�蛭��d�-)��'<h�$ᨱ���jGs	���{��iɏN���|i�X���q����`���s�l�tqkƦ�[f����f�;#�=+g�0N�y9Fcn�dq�
6��^e���_Ѹ�� �B[35�w-�JNrv�m�y�mY�٥1�M��n[K�#X!��k�͞Ḷn+���'%ʠ8�莪")�=Fkn5.���Kqt�!�74��Yzcj������`w-��H�����/1R�%�6�8�u���36x�7vx�wvXǫ`�$�HJj@�kފ�IS �L�X�����!��)D�`���9��`qn�.w/K��v����%G$�Ԙ}*`w-�� �T��ߎ�����M�`v�Dp�3����8��.��n�Zn; Z� �7N�z�2�mKTۏ�u{�v;�K �͖s]��������Tm�5#�9ܚ[�ﾢ�_�FB _��Tz�<}a�w,.Ż��RFn蚸q�	n#V��=�K��X�M,f�Ԧ�iө"Dp���U_/l�k���kފ�	"��o��J���'m�`qn�=�}�����@���`qw5�;�T�[T�R�I8
k�n�3�㬺�q¸w����v�l'kodE�aRRL����9ܚX�4�8���-�v+�D����2��3)��DB�=:���wy`w�4�;Z�ZI���RTr$�,.滒y{��&����P� m���p�7�<X���Z����)��ܶ����	"���u��Jir(�IQ�HԎ��ri`fd����k�8�u�]�e5�RHN��Q�K�(�[l� ��j���ۋ��5[v�k�����;q��H�$p�ܚXY��-�v3&�3tN�Sn4�ԑ"r����{
d���,7ZX�L��ꪪH�~�z��Q�U�6�:��k�*0$���X�r�W34&���R9UV�!*����,�Z\�����I�� 2$`��PB[�r��`�h�� �h��8X�4�=כ���ޖ{�K ��$ִ���k�55��6h�s�td{k������vۆ�tq�]=�p,r]]4o�;��Xm���EF�Q�?^[ǃq9D��6�n�}��l�������`qwu���2�Q��l�(�ފ�	"���u�ܶ��֝����$j5,̚X]�v��ɥ�����܌l$��������[u��EF�T`w�7�����v߯o�wN�5N��r���urtj9���y��9l����k]��cqv��.�b�(���q�2��ك�|�޷c�`���5��D�"���]0��.V�y.a�r�&y�zV�vdCs����b����ph�(�t٭��t���N�Y�c;t΁ӵä�6����m���r�W\4?����(K�n�(M6p�S-��绷��������\�T[�"B7E\:�Ň��8�[j��<�&N�y۶�kQ��qq�q�Ȭ���}~���Q�������F�fhbBH5-`{�Q�=�]v���f�)HA6�D�`g��`v|�,�B��}:��c�,V��$�Tԧ"r!8X]�v��ފ�	����/��5[���Z��Yu���~����e_��$��i�)�l��c�f�f4��a�a���/qm����[��F��q"]�R,S������e2���e���|؈]����,�y�n r&ԍF�����K�}Q*!E%�8zi�X��,{)�stN�SrRc��Dp�8���-�v;�K3&�u�iJU�Q���Z��[u��EF�Q������z�� 1�@r;�ɥ��������=8��e��T(Q>c����'���`L7=��q�[!�l�����l̞�W���<�tb��M:�ͷ�����K��X�T`{�m�ẳ�Jr'"�����~�#���`wvx�3�4�7��j��N��6�8���$�}��rzsЃ�i� �5 4ns3ѡ��� t@�B���JC0@�)�*J@��\(�B�����41��*F�d�M3B I�HJ�@-�\T��.�&J��RT���A��ʀr�T�h�"�6UP#@�4�}�r*@� "N A9���	
�� �4�G���*�
������N*D`z����Q`OO�Q:��W �"Dy{�Ζf��RG}[��DD�#cQ-`z�������X�.�=&�Q���#P����������`��`s2i`~�����8�b�ol7Է<�9*��	����*{&#T*����Ӆ)9�M�D�p�[�v�}�]�֟v~Jg^�ŇT�_"~SJUr���i��w�����f{��g+���~,��?}_W?}M���
�)�H@�Q�&�2}��*�`w$��;eLV6��m
T���ɥ�����I'����0�}@?�4sW������瓒O����,��f�r�3P��Iu��g��dT`{��7��~8�i3+�]\���K���/^�:Z����\ZŴ�˞�=^�zr�mJ��`��dT`OEFrK�mf�N�")*F��%��ɥ��ɥ�ř��9�����V�r��i8�%�`OEFrK��T�슌fm'pn���J'�3]�sse��ɥ��ɥ�޽�j%���Kuk �0;"�z*0;�]`J�����8$G�Ф ���N�4:�mЎ+�:M;���j[�d�]�-����ر��:�1��1�v-��a4�y7T���O���pl�c��4l��mg.7B5�_F���R�t���E�����=�Ma5��m9��ult��-��C��)t��6n'Wl@�f���i�xt��)������H�lE�z����X61�6»K�K.ٚؠ���NC��s&˕���C����-{�8��j�U��dKa���TR*Sq@�P�=饁=�.��S���ņj���.#5	���Iu�vʘ�4�;Z�F�⦥:�ƅ!`qfk`��dT`OEF�.^=7Vj�u���vʘ�Q�=Y��mekI�JP��l�X̚0'���%��*`K�ɜ�8m����(�J65
��U��Z��ɽt��]`�J��백5���So�ߟ�����c�u㯢"";!��K��]I�n�rnm�sg$�_��r!�b����V��X�^�2fsQ;%!G)"8�n; ����d��W�nl�`un���հ�)�8�I(rK�*0'���%��*`w��x*N����`gri`j��`�u`?7j�؅�NMG9�\(PMⲹ����j�!��:s���M�Y�1궺;l��MJp�D)��`��`own��M,�������B7l�T����=$�����i;�J6I,��Ձ�ɥ���S��� �'�����9$�{��$;���nP�m�5�U��ɥ��2� �0/�|`vK�փw�swx�L���c偰�O��t��V{+K�}���z�BH��$��2n�ãx+�Uwaw�����v4�[�7J��	���n����&���	���%v:�l!�P$�9%��ݺ�'���Xl���Ey���[���$,�\`OEF�.��S�mՁ�]�I�MJp�D)Ws]�u����GTr}���9j��Y��Q�V��S�W��ZX���F�N��D��:��Dnu��S����m����{bd4��a��b���k�ZF�J���#`䓀{w�Vw&��� ������G 9d�Dܕ`OEF�[��T��W�d��h��G������`��`nf�XܚX�hZ�EI����T����==.�;�P����b�ĸ-I�}+�z*0.zk�nl�3����7)���1�J�Y�Ѩ.wM����g!�,����!Q���2�Z�ˀ��v랅c;0��:q�lr=�󸺍�J.;V��=Y:ε9��ɤ�l��A�*6�Ex�m�;�Ũ��űu��om�J�S�ݍl��C����̺+=�g�t����ir�[�O���b' �ۭ���B���@���nOg,���;��{��{��&�}q
/�WFV�a�͎^6^��x^��;wV���ˋ�77�6�Q7+�ovx�5w5�76~����f����͞c����G�����z�L���X�mX�X�ڸ7��q�76X�۫;�KWs]���֓����#`䪰�
w�Xi`9�>X^:�;���rq�H�I�Vw&��� ���{�u`԰҆��&���sha�5z�n��a�L���VH��F��l�<���IM��%������9������XܚX״-�)T�Q�H�rI<���tpAa= �LuB~���1J����0.z]`w�r�8��G%��ͺ�3�4��}UIyf��}��;�mII�4�dqD�V{)��c�u��P�q�U���<�ӎ��ऌR��Ի�����Ձ�ɥ��wG�!��Jm�^y,u���&c�&���z�%��i�{k����Q� �H7��q�76XҾ0'����l������H�9$�7��W���76x�<�|���,��$�n6���9*�����s�|���	$�$���U�8��6���f�w�q��H�N���*`_J�����]�2�i���Z���`�����	������9��M��)ē%EMTn\��]68�r�c�G[��� pU�۴$֨J֌�j�ŉpZ��W��T`\���9����b�NRp�m��q7*������*`_J���=�w5o75��=.��S�W�w&�a�m\���q�7X�S,�S,)D5�%AD2D1U��������ߤ�����#Pj�1$��T`OEFsһ �����L���H�!�Ѻ��:үR�f��1c�SgN��\�l^^<�mY��F܉�F�`gri`qw5�76z�����w}I��Jm�q(�,ϱ��~.p3���{_{)��2n?P�Q�ģq��v���������}_������1o�;�z��c�)R8�#��Ի�~,��s]�꯾�T�7��`g���r��nD�p�<�`lB�1�:����e2���<�$�t`5�v@�ER*@�e�"���>�H8J�Xo��>a+�V >5ܢ�#L��
�S
�! <G�����@!G4�XüX����w0"��n0�H`��RP�Bх�-�� �x���E�s!Z/\�qHB�	#�@ ,�FD�F)j,H0! ŘB��+ @� 1	/�@�&u��bƥ��2����M�����R0 D�E�D�z�OQ �
�x�Z� ����� D��z����(f@�:t��g~k�$��Ƚu���Jv5��p�b�pZ����rk�fu�k���#��;�M���CYB��Zi���csCŹ]g��@���U� �-\n�IyJ}b�U�̭�N�Y�ģ�'�St;v��Z��8�r��Wk��f���t���D�%Á&�X4%+���7t�	zY$�,�4�֎	%�KEZ�>���V�v]xeh�؈k��nn�,�ٻM8洝P[uv��1r�ڍ]�;B��7;�Sm#�$�;��������}v��s&N�4J:��k&0Q۳
9s����kf�v��U[oIi��ӗD:p�2^گc��nwnN�㛅��`�2�wn�ډ'��x�Ė�83��L����(��X��n�4��m���e\u�ِ�qB�J���J���TsYݴ�1<�f�����!լ�۷L��(㎳�Y"k�}v�;���Ҩ�l(UmR���e������K�枴����7AGH֤�zI������^g)��'YU;�N���8���p�R����֧U�K��v�6C���jF�N{n˻*�l����b,2�Y��eI]�`�xŷN�̪�e��~]���D�ң���c�aė��'n6�9�	@�W[��mT���G �tA�7a�÷�j�����UeZ��n���Q���$��B���m���cXT'�Z�43��!�tjv���e��,�6� kv���M%���$�:�:q�nB8qi�h�v\�T���f��x���cA
�ns���6�5c���es8�:u��..6��*�E�z�H5O�~2w��p�V0��듦�ձ\�A�N�.��uKN0����{]�CU���0 �n(	��W��U����eۣ���6�\�sp��U��\q��0/����fb��q�m�]+a	�Z��(��lv��8k���dMu�OR�.W��ȧڶ�X��uc�*-��cv�n���zp�º퍤)Y]��]ٺ2tV���������� h��z(�O�LP~
��*�|�C�>���c�8��Q�%ۓ	�Ivt�ɲ��J[��::������Χ��{�[=��A�_n.6�؍��{v��ݹ��	v�8���l'Fq��.��l5��i���ttl]����s@D��L�s,�Ҳ�/3(��q�9/5�7N'b۴�ہ�cw�G����A�� �\���"ea �C��lr;i5�{Y� ykk�J�{���s�Ч���+c	N�:��g����Zv�u�(*ݶ��tp����W�&����:�ƅ!�~^�������*0=b�йx�č@���Z�`d��_�D(�3i`f������X�i;���8�
G`w�4�;�4��%՞�5g�����#�r6�[���Q�ܶ�g���Q���&\RJn��������`b����*0=b��#y�a��Di�:�V�3�*�8/bɇ�7����{�5��(R��F�q��.�;��X��;eL�n^%�5j�ĳrf�rI��og4C�
��{߷��:۫'���"���u�iO(���HԸf��>��vʘ=n�'����5D�5)Ԏ4) ���'����e2�b"s]�`6:���5��Z� �0'��z*0nl�;�)���(�H�PjD�O��7�Đut�mt�����q�,�I6_O-jr�݋(�X�$����	��;e_s��P��X���$�Ir6�Q����2�:�Հu�=���Q	L�{�e�h��NAD�`��X76Y��P�aBU\��X�S,{��j�O"��#I�,=_U%�o����Ł�ɥ�R]�pu��BRi������@{�P`���*`�L���g���*�\2��j��6WY�\�x�Sbd�H�]��ՠ��6���HOEF�*`��dT`{�W1GMJu#�
B�9���9����b�z*0,�=1#P!n�ũ0�S�*0'�� �0;g.�k�	�)%������`nl�`}�w�|� � �$����F����}��$�(H�M�H�`gri`���*`vEFe�w?bXc�^==-�u-�(N�Hv��q���]祼��
���F&Hq���(�,��,�T�슌	������Ŧh����rf�U`x��"!D���K�,��,u��BRi����2*0'���%��*`v/��#wR�ԃ�Q�ܒ� �X̚X�TLQ�R�#�	����>X>׵�<�i`g��`ZJ#�4
� �E��O0�w0�6����sYsbL��Vx{u�m���N�g(:x��#Ļa$��F7.No^�M�q����'<���7�����Q���y:�7F�����#��K���_���ʞ���,���򼦓�)C�W"��[�b��7��kH�V�n7f��Ս���Ӑ/k�"�V�I"vW�l�٢�M�kk8�@8�8�qڻve�e�E��w��x�{���C�MX�+FQ]����Tl��;�����2]�0�u����i�f�Ѹ(��zX̚Xܚ~�︃�w��ﶼ�n�Pp$n(��3&���(�:�������u`{����BF�mȣ���ɥ�Ź���G}����7u*w R7M�'P��׼�kڰ3�L��R�ޖc�K��N'���9����Unm���<X[��h�Ť(N�P�e��0��ů8Ty�sm;���۞9"��l��ﾵ-;�JM8�#����nl�`gri`qnk�}\@w��`w^�R�Q��$��,�M,���꺯������3���9�4��U_$f��5)�8��,��; �����K;�n��	�1j��*`w2�`g��a�S�7��=�o&yˡA�����X�4�=�}_V�ߎ��y�76X��!��aR��JQ4���'$�7ic�]k��P���bz�.t��s��h䐊�nF�,�M,-�v�͖fM,n�T�$e7I�J���z�L��ڰu���;Vu�%�)&D�#�Q�`����ɥ��S���q�������<j�Cj8���i�`fd���ͺ�8�u�z�ꯒ�����~�*8�M�RIF$0-��ܶ� �T��*0;��7�go��}m�b%Ⱓ��+{vkX^A\���[�}����kinU�'.�����[u�[*`I��������HH�Q�V�eL	"�w6�����`n�kI;���H�QH�EF��0;��`ʘ��$"�mD���}�Խ��*����� oX8�
&N"�P�[�K����E>nF���w]�n��3)�mڰ6���X8j�J�ӲIN];9tYֳ��禮�E�n#����ʒ:�M2&�B�> {���32i`n��X[��ǫa��q6��W*����e��M��V�wy`�/�W�����JTqF�������?~��Ձ�m�ϡ%�8}��U����`{�W�N:���⍹V� �ݖf*0-��98[�Ą�w��������e��v��o��P���|NB��-�&]�7e�3�u��\�;Kpm-��;�kZ�v�^ݑ`-�s۶��^�����Õ�8����zM���d����9�]s�z��)�馗�%�xt[ևNz��%�2Ւ��x��6�$����X�[H+�)ۧV�ݞ�a���+����.���A�_}X�ܓz)gk<�;Ug�ڥ���D��f8��7[\�m��'g�aݘ޳ݟMNq���o�����e;�^�xf��}�n��c��:K�Ky�Ԍ;y��sh���ܫ�Pp$n(��~���_�n�mL	v^%�X���3u-�C�_�n�mL	"����I� �O����*����`�Vl�n��7wmX�b%�rx�jՆn�`ژEF��0��s=�����~^�"Q����fM,۵`v[|�۫TD(P�ɫ.!E��4-\QZq�TX��9��w [��{;m浒h�i](�̭���r��I��j���`�_vA�ZX��j�\�7r�Mͻ��rI��{���� D*�X�'�@lTf��;�v�̦X�j�)���rrj���k�yU� �ݫ3)�lBS;���/{����ѡ�%Q�����XܚX�j��|�؈S;��`=��U�"�6�Mț����u`{������{ޖw&��X�J):�"�i&��x��jp�tVGt��{'qt�Gi�u�{���-&\�J����+�u{|�wvX�}�K���}���j'�Oi�Ն-Z�-�0'���_76_��U�6{��~c"�����^�ŀ�v��Q�V�B�!
 ����>�D|	!L�2N�'��13\�8F�#���S� �hR� �ecIR���8&�:�D3��R�p��@I�F���T1"͔�X$T���#���p�h+�ԈR�R�1LW�����b��_��xUG�꺈:#�TLP "����""�^�zT>*��A �!��Ⱟ"[�E^mX��X̧G)W*k��J��*��Ԓ��ޫ ��� m�3�4�;�#�m8�F�#�6�X^:�6"wwk�<u���v��Q�w��w��0��x9��7`��G�7q���=s���i����'3�~��۾��f�$J�r����}V{)�m��	v@��������F�QI,�M,۵`mՀ6�^�29��\�4W�7"n��]X7vY��=�zX�<X�ԙp9�R45%X7u0mL	"�s����|`{�8e@n��j�Ē`ژEF���n�9�-Ф�q$�IQRi.���]�͎8P�mr���.��{u�kZ�9��un�-\ũ0$��m|`�� �ݖs&�ʎ(�uH���0�S ����*0=�-�֜u#M��r���,wvX�4�7sn���.��� �CrXj�3����i`7�Ձ�m��o��8�RK3&����r��wy`��!"�	LDG����ۭ�~�ޑK�Ĳq�v�����ًn��n��b����z�]�'SW������M\���\���+p����m�]=<�œ�4۶u�^8Y`�{t:sG]I�N��k��}�R��2D��ڙi5Pb	 �l�����P�;n�G$n�u]��9�=b�/(����u�-�����ts�����(>�[�d ע As�WU�Y?;���we����=R��.E,h,�V����ۗ�X����:�5�WKh�X������?�w��n�eL	"���w�AbsV��V�0;��`ʘEF��X����1�����l�$��e|`w-���"��un���%�0$��e|`w-��-�0="�ԍZ�wx!-������[u�[*`I=�]�j\E�V�١�.Ҙ����m9/h�ƫ�n������7H�R.���������l���������p|�Hݓe�.f�$�����(�*&�EjQhP�J�%��K76Ձ������.��	n�X�`zEF��0;��`ʘ�KP�wf��^e��ܖ� ����9�GK�����(��r�-�vl��$T`[+���t�n�Xۋ�4n�ٲ�s&&q��{X�ޞh"���h�A�U4�p:��ܦ�����X̦X�lvC��y`n:5IJk�j��j�Z��*0'���-��͗ꤌ׾����M҄�$��߻��$�ϻ���Ȝ\#!����c 
>���g��o$����`w��ڍ��6����s7e�u�3)�/�`d5�%�MQ AGI����,V�ߎ��ŀswe���L�T�A�BcP�48����7A�%[kK<r��<6	"�.;O�����9DMI,̚XܚX7v~�U�~��`{������pmě�n{)�����{��kڰ=�L�:۞:��:q��Rn� ���=_U%��Ł��Ł޽�mJ�1ʓʮXjP�}�j���K=��JA��g��W}��s�O>���&�7uȝG*G%��ɥ��������:��v�͖�����r7Pm���ٜ�c��g*�m��kx�Km&�4��۩n?���_|�%��P�����<XY����,�M,�{Q�(�� ��`vq�^�L���X�i`g��z�ɟz��]5! AGI����K��K;�K�7]���Z5j$��Ny5Ua�N7zXi`vq�Xlϵ�X��#��pmě�nw&��ǻ΀{^Ձ��e�I"!(^!%�AF��D[HIޓͦM�K��]�u��msm'F������>p�V�\�M��[��j��a��u�n�Ab	��}��u���.wm�p떘�5�#����򬋲�pt�Ln=��G]v�[U��s����s�Ū3BX��	�� `���e�E�su�Qŗt�s'ܓ�P����<���.9Ճ���u��c7��7'<�P��&x�'�k�g\/T��?=��w�������m�Ħ�:��ҷ<����q��|����-��9Y���������ى�Ks$@=�����*`zEF�T�;״-�CFSnRNG`��Ͼ�%�D.p{��`k���;8�/b"d�t/S%'$r6)*I%���Ł�ɥ�ś��9����<z����(H�U�K�zX��X^:��"#�I=����7�S�#N:q��A	���P�{���A�6667����|������?N>A����w�� �`�`�`��"��촔���̻�.]�]��kt��كB�;�=�����u�} ����ލ�8eݛ�m��37x ��������lll~�y�pA�666=���8���~�>A������?_.�M�&˹��� �`�`�`��{�ӂ��Ŋ<�=?<D<� �`��������lllo~�����lllo���x �[��ߦ�黛33m�ٹ�8 ���~�|��������|��?�r9�������lll~���ӂ�A�A�A�A����%�7s��n���� � ب� �{���� � � � �w��A�666>���8 �[��~�|�����o�_Ɠ&l˙sI���|������o �`�`�b�� E_�~��pA�666?���ӂ�A�A�A�A������A�A�A�A���N��ܲL���.�qE�\�h�i\b����n�焖\��ʺ�����xd�����d�����A�666>���8 ���~�|��������|������o �`�`�`��w����w3n[6�䛻8 ���~�|�-�������|������o �`�`�`��{�ӂ��A�A�A�����s3p��2]�e͜|��������|������o �bP��AO�@������N>A����w�� �`�`�`�����|-ݛ�m��3wx �[����>A������� �`�`�`�߻�ӂ�A�A�P�T��s�߿���A�A�A�A��?����fi6\̗wx �{�~�|�����߻�ӂ�A�A�A�A������A�A�A�A�������lll~��%̷��-�l��`��Nqs�����.���u���[�l�Ց�7N����y����w6ffۙ�s6pA�666=���8 ��{�x �����>A������� �`�`�`���͙�n�fnLۻ8 ��{�x ���A �`�~����|����߿s�pA�666=���8 ���������c��rX}��3&�{ꪯ�����;��`ori���9#�$�a�!$��ޖ�ZXsXqBJ��	��POC���"l��7�̏Y"Q��DR0�w&�ꯒ�������o�`w2�`w�$h�sƹ�^�ĥaF�I���kX^A��:؊���rר��:Vx��0b��m���u`x���e3b""; �֖F�j�JB@�6�$�nl�������l�z�,{_��W�B�3E���L��Q<�	���֖{)�}
d�{,��K�lqԎ��p����K�zX�ڰ�ua�%
'�ߋ���ME"TӌQHX36X^:�;�L�3�L�;�"���H�HD$��0��Jjj�Z@X��y�q��+!�B#�@�tĿV�ÅHB �4����FU�T-JS��`qF5�$�VT��|�j���I�wqP��� ,# �H��B H� ����b B[TL`ς8®��:��) ��Ç�*�x,I�	��%�(B(ԏ��`�z���8'Q���!�3=��ƨ �C��u1l��I�L/lqXA���<7N�$hٝuۍ\s��B󵷏���dy���sK�hwm/�X��X�m1��f	-[��9SN���#cv���*�F�C&�^`q;2�G�*z�QT��ֳ�����s�g��8�!Īp]�;<�s.Ѵ
� �e�jj{]Α��l��kGbۃ�A��N�,sص��\�K����΋3ؐke�'��V̄k�-�-NȻ$-�Id�Ԗ�yj8�`��V���cl���۠��fx�$D���ݺN���<hZ����Hܼ�쵎[��^�=�7�� ��;n"��n����{h[GX0����ӆ�n��!	�<� �u�4�$�q�#S킒d3b���E����t��l�ܲ=��MƑ'n�gN���x*�\�n&K#�[6Ht*��s<� ]�$)Z��V
L��)t�' k�M��Tk�ܯG��e��m4FJ^�r.��u3p�(=9��s;m$�$t�.�̖�i�N{I�)���`Q��y���G9�s�ay�&R��[�T�'i*���]N���K�j�s�e�۲�2�3�Z��q�:�Ŷ�Λ�2�mT��qR�h�mM�Z��[5�(%Z�li8�t�-����Ö�:6��$^;v�,��S<�d�u�h �Ө�b��B������˦� U����J�I��h�\�ru.N�&������EO$�<L��e�vh��y�ttq�� [��Y��V�<;�S/��O�7O��XV�5>�d��b�C���*��tU
��g�����u�=�b�A�uhV�i{�UY-�9%TQ���eX��Wc2t��7
ID��9�y
\s���M�f��^����he�Y:���A�m���.��e��u]<��J�M��@U�e.N�g(.33��^�=�i��vS�ci��
U��r��l݄���_��g���Z��W��W�O��F�<}辩�54爞=^}a���8�=�ݣ���yHx��Ռc�q�w��G�#��I�M�_��L�՞��A�p�ѝ�p��M�n�S��֮bȸ26n��zM�<ر�"�#qO>�6��M���MW@i9�-\bۤ�,Jt����Z1JG�/c%u�pW==775�R�U�c���{Xy^^����r!V�[��;!�&�ֵ�0��K���zCr޿���ܜ�q��J痮����Fմ)x̮�MS�>�-�q�K������{�}�º�2Ji� �rhw},fM,�S5B�P� y��q�:�R�W+�U�%ĒLȨ�����T�;e���U}_}M��G����6�JHB����� �0�S�*0=&+�m�J1�$LR�ﾯ��鹿w��`w2�a��%/�`b�͛S554����R`��dT`OEF�6X��Y�K̠�#)�M�����o��c�x;U��)ѷj�զ�}�:�e{WF�}�������*�J6)&��O�`gri`��`��`�Z�u#�n$�#p�3�L�";
!bI-��r��`��`s2i���#���ME"TӌQHX�ڰ�ug�ϛ�,���=�-�C"��NSQ�a��K��K��Ł�ɥ��.��X͂�2!��LK�RLȨ���������9��`gqC�t�Ā��*���$��:��r��b0��OW�<���\�ݥ�h�(Y� Iz*0�S �_�߹���h{}?�z?�أ��)��q���{7j��u���e2����j�J(�8�r(��,�M,R�O$� TDa*��-���mY`�ڰ<��753*�A���a���?o���7}?�͖��� ����q&�M���ri`j�k���v��S,�O+��.ɓ�<-b�\%��-`�&��bnwS��L��S�BE%!��o����`���=�T`{�8e��R�i�j9,�ݗ�͞,͞,��/��W��G�`�L�d�5)IQ�,���=�Y�""d��� �nՁ������6�9
$������9���y�{��P �,D5Q���_}����p�=���I�:Q��"b���S �L	��������>���?�x2um���'� 	���\s�S\.�+w"�	�1LսNx�E�s�2���&�T`{�Q�vʘ�)��IA��6��3�4�W�Wߩ�w��`�ߥ�sse�nV��i��r(�`gri`��g�H��������shwC��r%n�͖׎��S,6%�,YƉ�H�S\��պ�&�*`OEF�T`�wy$���
� EB�}�wK�ת��;��96�\x��h��	���Y�NéՅ����\�=���{�=�nllj�[Ssq�㝯8t�Z�Lk[vhp�mX30��&�nu�<1�c�.���-q� �ly��p�O�c��kj���7fP��m�[<v����+S�Ol��[���Tɱ	��=����;��.�����u�p�@d�N�'�����4ڋ�A/6sɆXz�w.n�앴ḓ�z�>�68�m��r��d��v��K'�t4iN�9�$�M��������9���UU�}��wc�!$mҨ�9�,�S/�2׵`׵`g��DU}�FV�^��%)�$LR�o��u�D��J��e2������:M7����|�76X�<XܚX76XҴ�\��m�I`gr�`jQ��:�{V׎�O�;g���ݱt��^L:�E�Z�hN����t�d�Av�oMl�h�dX����o�e2�:�Հu㯢>��=�׵�`f��5q$9�"Q��`��|u�]Q
U:�:e���e��}�6�����q��q��������F�T`��}4�sPjũe)������P��,����u`��`s25��#n��
#����e��(IO��t����S,{��?i���\�0Q�M��:Q⋐��*�NK�41��ٶ��qڋ�ع�e�Q`x��:�Ձ��f�P�d:������t�QJpQƣ��9���}T��:��x�K ��W�BJ#�G8o��pJI�)%����Xܝ��?���*���'�?g=�I'����7+6�u#�7�D�,?}��Kqޖ�{V׎�>P��,f��d@�n��G��sse��睊w���76x�3�4�7�i�M�F
))J�uνsi�Yq1^8W��3қŚ-%K�>��'apĀ���-I�vʘ�Q��ɧ�����K �k<ڢSq)�I$�z*?�3*�`���l���'���>��r�6����0݄�C����T�;eL	���#Ŵ���Ju��B���}Iw��`�����~��I⨞	�"z����;�����j(�8(�Q�`�ڰ6!$�ޝ�,�X�X!�1m�l����[��Վ��p�sע���M�y� \v�ٺv���6�K���g��`g��`m���{V���R8�qF�Q������9���:�Ձ��e��|�#�1���eI����G��g�~��͖~�������������u�jST�@ۊI%��P�ϵ�X�i`g��a�D)�7�`�g��RiG���`s2i`{�_DD-{ߏ f��`x����	C�]�q�ݿ�%y�9��n�=U�t��I'g�t�7<�7,	q�6��\� si��{lѶ��nQ�� �[m���;�ƃ��̦;M��0[t2��ē���!��E9GHZ��[qӎ4f9w��˵�C��g3/@���%kEhN�c�����0�<����[���X�{J���6pv^�l��\�4�h73���vܼk��3�-u�q{�ǽ���co��瑮��#e*f݁��Z�V�Cv�xf��mԷI�;4�/V�m�����ٖ��V׎����u�����N:#)��!`���������ݫ�֖{)��	L���%�MMMsQ�V�Ԙ��&dT`OEF�͖t�6��U�lRK��K=�� �c��
ϵ�X��r��չ��w�P�����T�;eV3&�7I��T�0�5��8�����N�Y8��<�/��:[�1�`j�v"���{����ȇ9�7 ww��9����d��nl�`ec������	��O;�w��OD����N�(���;[^,{ZXs_�S!���:��Q���`wvx�3�4��}�}T���K ����qG�FF�=�@-Cz*0�S �0�s�?r�}UU��=�~,�?~���Jq'$��;����BS�{]�֖{)����~��M�%J��(�C��q�F�9y�b1�ڧ]FX�)�@]��������o�"%8(�Q���},fM,�M,��,�Xm+�Pp"M�I,fM/�J>P�!s���� �ߪ�:�Հ<��qԎ4ۍ�8�`gri`��g�Q:�@�V��)�<E�B� x)+�#Pa䑄m����F�a!_+�H<W�T�$@!�H���(,݌X|j]�'v�QsIP#�U$��b���s	G̈D "��S-F du1*U8��h#��q0#��0>0aЅ1� ��1��z'A��꡵D~@ O1�\?U�z�(����p��K��K���!�ND����c脒\�n�V�o�`w2�`g��`v��������	��͖��(J3w�^�ŀw1Ձ�p(���}��E9ͣq��.�Yz�V�͖�+����)t�:jk����`g��`�u�
v@���1�s�FF�7R,�M,��,��,fM/�}U�RFV��6�t)�Z�H`���;eLȨ������]5R�q���W�UR]���7ZX�XZS���Q��L�>P=�⨾{{���'za[J���lRK��K;�K �c� ��V�	F�)�O&gB*�.���)����.�F6�bs��ؓ]���6�f�*C��U}�ܫ�q�R6ۍ�8��=����vJ�}j`vEFy//�$��Ȕq�X36_���� �{�����`w�4�;״-��M����G%�w�Ձ��e�
!)��ZX�ڰ�1m:��Q�Ȥ����]ݿc�,���>��L�7j��s\خ���R �,�&����wwӀ�ڰ;�L�6B�BQ	$%�h[�=s+v�],���v���\;km�h�F�4!�j��V9G�C/[q9�S]J���.�Mgdv.kr=>2	�f5C`�e'�6+`��$،�9��.�������e�@� �����mH�h�ɻse�1^�ϡ���yoa��圴n�p���u!n{M�\młh�]��<qv�[[qʌ.���9�&�]��d��DM ����I�Y&���e˱s9室�<r7Q��E�,���#�ㆲ<ۘ����{�����n0S�� n{��wvXܚX�M,��]5R�q�Ԙ}j`OEF�l��9������7��ߪ�IA� �b�X�OŁ��e�D��{V�{V �c\�*���q���������;���nl�9�4�9]�ڱ�)�"Q��`�u`jJ�^�@�u����e���g���Qܖke��3rk���#�u){�ܷN9��%���=����7jk��u`w2�`g���B����sX�N�&E�8ے��d��>������>P���ӭ,��X^:�;�Q��P�m�d�G;�K �c�5BJ&Okڰ<�i`yg1>��O�����K����o���ɥ�����nm��;�'t�PR�Qƣ��:�Ձ�(�w�@x�K �c�$����t���nH�B����}����#Ӷn���a۠�1�^�����7k
⮁��K=�� �c�Ĕ.�׵`��S�����mA�;�K �fՀu����؈IL�Y�rJ���9�7 �鹿sse�����|�̚X�4�;״-��M�9D�K��}�j��u����e��
g��X͇����RA7%��ɥ���e�w1Հu�T(x��s�	S�.L��v��.納z��σYQ-�z���V�9�i��W�Zj;�J��L���=����*`��dT`{�g2�w7�}8�,��/�}I}��wg�;�K���}_RGsǕ;�����5U�{^Ձ��e�$���ZX�ڰ;��ڷU�
6)%��ɥ��ɳ�I��wy'˿�)��"'���4�z�矹��O};�7*)iƔp�3�4�?}�U.��p�o���ɥ���{�ަT�6ڦ4̯R
�W#�Q�Y[s��U7�u���9��ۣ7*H4E"nD��À���8�5�ܦl}
#�{_|�O�iJ�T���!-I�ܲ�z*0'�� �9���UM��A*t��m��P͞,�� /;�����;�Q��P�mҩ"������T��Yu�߿~�Z�,�z�M�N��:q�HX36XO,�S,�S,�P��B�E
q�a���YU�{��g]T� WN�����A��m0ml���i;�۶��v�;�D���rr�[��d�f�Ga��YudF�J��"b8�X0��l�8c��uV���v�rX�:��k���]]&�-s���.2�����<�1�j�Fz�i�3�s�u�76-R���c��ͮE�2��b;HF�HvE�g�`t�s���cx�>��:����{�9����k��4���)u��猽�e��-�L&�֧M��'��慪wME*5j98,�;��K;�K �f����ƕG(���KX�Q�=d��ܲ����ف��8�)iƔp�76x�f:��Q	Dϧ^���u������IST�9�7}��~�����K�~v3&�w&�z����*r$5 H�;�]`OEF�T`��a�ݸ	��g���]�lq�.�n^��ޖ��u�n�T_�������\:!�S5o@����T`��rˬ{{�8�t�H��w&�J���}KT(�kڰ=:��{)��s$k��>��pR�͖�?%��Ł��Ł�᪝�QAJ�7�KB���Q�g��X��,�S,�X�_m�4�9DlRK;�K�}���{���~� ��V�ظ���8j7��(fvC�f�	��$�%�t�b���N�N��q�MJ������;�K �0�Sz*0;�Z�j��8��p�nl�}�A�o����Ł�ɥ�޼�m)J��H9,��.I��og&����(�@h�DDB$�P������F�_���=�{��:��NGӒ������� �0�Sދv���V-�jK�S\���e2��G�Ϸ��}�U��ɥ�Wzc[�m��B��#���x��9�7i�/mtPU�0� �;W);��j�bC �0�Sz*}�s��<X�<��5��q(�n:��G���:��:���DB��3\��iTr�(ؤ���w&�~��#��K ���漦=�(�7$	<�Q`g��`x��:�ՃJ!$���*@@���~s�}�䓧~��8�'��͖�ݖw&�fM,,�ؘ��ƜP:�\��B9�*/n�^vѮ��,�iX�S�L!�b��[��X%�0�Sz*0$�O}�UUq�o����<�R�"�� njL	���*0�S �?�Ϫ��͍��(qF���,ݞ,�T�;mL	���&�]7qheEqr�D�BIDL�^Հ{^Ձ��e��"%/�`y���k�SDҮW9Y�R`���T`OEF�*`idL������H �� ������T4dS��"�G�%@4�eq�
�A,��,��;�FԔ�������82��"�H�� �1Tt�a�D0#=��H���`$���H���P%� ���PG��'��*��PY�^B�����슣l�\7�AM�5o'Tl�듒T��t��uOC�<+�1]�=,[4gcy�m�)�����3U��6��$�+�m��"�c���Vr���� ��L�࣊Uv6갶Q�i�a��u5
��VI��k!e�އf� �A�t�@�3ۯ=�V�e9�7�s4�k��g��ؓf��v����c�-�\e���F��B"m=�`y�w]1��stv��/N+j3p����q��V��t���`�\nC^[��۴��Zk�\;�޳a��dΈ]��r[�B�J�j�X��666\C[t�V�������� ��h���jӛ��Ѷ6����C���]��q��c<����ܺx��&���99����%ӛ�4]���eV�:MN�L�˂�vˡ��ٵ;��.�f���GO5s����B�- 秋+uuR�M:�I��kvبA	Ѵ&:@�b��[�����8�u{e^1��룤ˎ6V"�'J\htR��/*9Ά3A�U��k�mNSA��HZ�]������ײ�@�v94z�Je��Uj�ʛ�3���nUWe[iz�\Xv�@��5 �F�']��9T�O%v5��j�ب(��+���b2�;(:�km2�R���8�m����痂�G`㊙�q�g���{aƦHx�4��v�쉝AՔ�)���%[n۪�V�9�HeK'�T��6� p���--c�����m����sm�s�4Ḩl����<;��t��v�s��`��}�zpM�2:N7=J�Y�l��R�y���m�9^b�MV�-��9�H�Y�P/.�i�(p��Bm��(Z;2�1��:SJ���-��!��;m���n�e�5�=����l���qsY���T!sNc{��I�5�%%�՘�(�q�V��훩�@p�)*��F0��je�_6��`q��R��(l&�s	v��� �5t�x�4O�Dp* b��}(�>EuUF!T�C���j�!ꉾOl�>w2晗f�͒A�6�d:5��[Ɖ��<vL��s�}N����v{u�F�Ka��Ž�WeJ�3����&��N�����[��urcmQ4����u�����4��xם��&�I�6�sDr�v�33���Z�^ ��أ�	ϲ"�O������\�8�u���2s�;�M���Zz��Ӹ]n62J*z1\�	F����m0���w��}�<�;t�6,�r�����]�TN�rz�3v�"�qH^�f���ِ�X�~�&X�X^:�%���3�������J�G',�M,��,�X�^����d��T�ks5`�n��{��`���T`Od���r�@jF�D�K��}T�������3�L��DB�>׵`nl<�%&Ej@i�`gri`grh�;eL�T�;&�w�Ú�-B�L\k��Ҭvux2��5���z�{r�\u�]w���}���n�r�m�H�G��ŀu� �n�P��i`b�֩�9\%�p�ͷvrI<���uߑ*�Z����Q����j���e������}T����t�PR��ģ��;�zX�Q�$T`���9Y�s8�pF-�LȨ��*0�S�s朗��`w�YO�%	�G(��3)���V��X̦XB^�/nS����ۮH�z��F�Y8��+̮o%�t��>hv��Z�߯���;�Ϧ�4�,f�<>���l����Q��l��ԍ8���͖3&�w&��͗ꪯ�=�6�Iģg*�g�V��,�S,p�!qyD�2!(J�p h rNw��$������r7�9C�6�DG;�K �c� ��VD%	|�%���ŀ����M��O����s3e�sse��ɥ��ɥ���ZB���CP%&�C'+/nu�㚍�]��ˈƷi��25�-z�}��L��()Q�"#����X̚X�|�B����ыl�reW)f-�I0;"�z*0�S �?�|��=e?T�)�Q�����V}
"d����֖S�%���.o1.V�d��vʘ�Q�b#�	'�vo}����	�(95\�-Z%�0�S�*0'�� �,h�3h�MG��o�>�Dt�Zی'#������g͒�5ˋ*먴��`�jA��0;"�H��;%_s��=��,͍��(qFێF��`fd��(Q2oj�=��`w2�{
!D}�/z�Rm�
}8�R���`��g�K��Ł��Ł��˨ₕuRW*�5(���Ձ��K3)�}UM��X�x��8Ҩ�J4��s)�Д$۽:������) ��@ ��@��I��%�{G>]y��b�gl�ҠU:c�7�m� ����]��@厭�s�s�n���9f������[R̝��A���akHB��Ñz�x:�94�24b:�N��3fN�X���H�:\�6ҋ����N�݇ӵ��km�z����>c���u�1li�Z�ɋ��Jn�m���"���h��1���L��'۽����[z�7QZu�br4�]�']������9��2��i�.��N愥"M�#q�@�l�X36X7v>�� ���`v��E��:rQ��T�;mLȨ��*0=�j%��G#��9����d��U}�[�<Xw},��m:��J69g�Vs)�fS,���6!B����3c~��Q�"�!8X�4�?)�{] ��Ձ��e��B^���v�s�)����<��k�k< <�M��Wk�2<ۘ��i�d���`���oj�:۫��Ϣ!.�6�K7u�]G���`��k����uP�$��]�n�X�2�;����`�ڍ��Q�Ԏ��d���ɥ����H�論��y�ݚ�r��7(��P��*0�S�m�dT`r��E�H�)(�G �f��UUW_���;�<X�4�3���oR\g;��mv���t�\fG���t��^��\s�\��9N(
"P�$q�9,��,Ȩ��*0�S���\�Y�i�)%��ɥ���H����;��`qn�9��9C�6�RD'3'g$�Ͼ��iÊ�*�'�@��2�������`u�
7%>��q)���7�`zww�s)�fS,6�J�I��29,-�v3&�fM,��,�pc֐2TE	SO��\���}o�����a���;�nZ�'N���_��*mF�G(�R�"��OŁ��K �f�z�U��٬�"��I���`nd��_6�pc���μ;Uq?�U��,OO����6��74��sdND�,K������%�bX����ND�,KϾ�gȖ%�bw��Ȝ�bX�'���^�.I�.�ܛ����%�L��_�(s�?�����*dLʙ����8�D̩�3*w��dO<��3(z(�/� P� `��o�<�y��'�3*dLʞ��t�4��w��[�q<�D̩�=ϹٜO"fTș�;���'�Tș�2&{�ws��Lʙ2�f���*dLʙ���~2�I)]7Ksa%�nI�֮�ݧPp�<����m�v�l'k��f���w'�~�vu"�������{��r�����"y�L��S"g��w8�D̩�3*vo{q<�D̩�=ϹٜO")�w�Ow�m�g��u0V����D̩�3����O"fTș�;7���yS"fTȞ����'�3*dLʝ�|��*~A��S"~��ž�vf�3wvnn�ș�2&eO�~��yS"fTȞ����'�3*dLʝ�|��*dLʙ=߻���&eL��S��߯�A�X��w��{��S��w�����y2�D̩��͑<�D̩�3����O"fT��n��9�������r��{�����uE��I6~��Lʙ2�{�6D�ʙ2�D�w��q<��S"fT����y�L��S"{�s�8�D̩�3*�g�C!s�������^�Du�	to-����<��1+Gi۳۱\��iδ�'Y,lk�w7nu�8��ki�Fڍ�����B�g��6Z���kr��F�_�v�Q���j�M�J�+79y{c;��D���"a����f�=�n���5<p�nen.koA9B�^�*�1r�s�HV�эAbێ��b�f��l�Z"�&�t��Ş�r��������wy#��L��<<��<+s��)G%l��Of��Tx�Kt���l�nz���CUēm���=��)�w����s��Lʙ2�{�槞Tș�2'��;3����bn�ș�;��l���6��}[���P�AE##r;��&eL��G=�sS�*dLʙ������&eL��S��ȞyS"fTș����'�3*dLʝ���i���7f\��O<��3*dOs�vgș�2&eO��"y�L��+��Nr�"gw���ș�2&e���jy�L��S"{�}��7gD6j1Y�����=��)�����'�Tș�2&{�ws��Lʙ2�{�槞Tș�2'��;3��Lʎ�)��-��lK&/�
�����&eL������y2�Ḑ��C����O���3*dN��L�y2�D̩���dO<��3*dK�ﲙܲ��'G=�u�A�1����^ӱk�仂���=Q��W\�mk�L���{�'�k��ݵ�=�sS�*dLʙ�߻s��Lʙ2��w͑<�D̩�3��woș�2&eO��yr�7vM�p���O<��3*dOs~��'������"-�O��H��k,���D�D�=C��ܩ�Lʟ~��ȞyS"fTș������&eL��G>�sS�*��7jdK��~�n���ۙ�n[�s��Lʙ2�~�dO<��3*dL�~����&e	��G;��jy�L��S"}���8�D̩�3*t�p��sn�]����*dL�����s���'�3*dL�9�߳S�*dLʙ�߻s��Lʙ2���"y�L�����fo�D��r�R26H����<��3(���jy�L��S"{��s��Kı>�y�'"X�%������y����ow���������&Y՚�r�9���,�n��=�מ�F�����2\�OdY����7���{�����~O"X�%��{͑9ı,O�ߧgȖ%�`߻���Kı<�{s�i2m�3f�Y����%�bX�w���,K����vq<�bX����ND�,K����'�?S"X�d��bY�ڛ����7���{�/��q<�bX����ND��UDub�  �^�,JC� qH��H	,Z)��N����$P�x��ƚH��o�C1�eeX�X�%aB#B�#4��n9��
-BR%aB%ee-��kJBR�ٍ�-��Xa�YIB� ��FYx/O5_qT�)�ۤe`�+/��B>�F�*��/���g�J.d���<��#H�'�rWX�VNЌIYP�/�zB3�R���U���%؁u�)ڗǚD�C���9�X�1@��bD�C�
	 �Uċ$�� ��� ��'�C����D�C�=_AQ��!�'\��|#���O3��q<�bX�'�w�"r%�bX�w�?z�K�Ui������{��7x��sS�,K��;�s��Kı>�y�'"X��dN���Ӊ�Kı>��s��l͓e�33sS�,K��;�s��Kı>�y�'"X�%������yı,�{���bX�'�)���a���f�����M�.�%�ћk�m�;I'cFŗM���Ԟ	W4�]Kq�r���=�bX�'~�Ȝ�bX�'��ӳ��Kİo��h~��M�bX�g����yı,O���
p�n�̛�w.�Ȝ�bX�'��ӳ��Kİo��jr%�bX�g~�q<�bX�'�w�"r%�bX����|�I��3n�M̛8�D�,K���"X�%��w��Ȗ?��Dȝ��l�Ȗ%�bw���8�D�,K��;f]36��3vm����K��FD�w�q<�bX�'{��"r%�bX�{�N�'�,Kx�T6���"X�%���۝sI�.�6n�78�D�,K�͑9ı,?'��|�?��%�`��f�"X�%��{��Ȗ%�bS���ٻ�w3	�����2	%�P�]�t��C\^�蠫�(�v; ܖk��-�ݻ.�Ȗ%�b{��;8�D�,K���"X�%��{��Ȗ%�b}��dND�,K��r�t�۹t�wwf����%�bX7��59��ș��>��8�D�,K��sdND�,K�w����'�2%��+�w88I����gԏ�R>��߿gȖ%�b}��dND���2&D����8�D�,K�����Kı/�v��ۥݷ3dܻ��O"X���߼��,K�����8�D�,K���"X�%��{��Ȗ%�bt�p�6��ɻ�ss6D�Kı=�~��O"X�%��;��jyı,Os�gȖ%�b}��dND�,K��	��J uG��-U��;��3M˻wt�%˛q�)w�$m#�o���|���Ө^a����n�'u�7	����6��8�E�KN�E�`�z����`����[ocv �]����}5#\��e6��e��\a8���&�r���löÒ��$U*�zeuq�\f%Rݫa��y���S��"��L<$�a��k��m�N��ۜ����_�������w|���^L9��2u�E���ݸ\�����M�����p�ڬ���g�s�w&�m>O"X�%�{����Kı<����yı,O��l���&D�,N���N'�,K��;��ri���Y��s3sS�,K��;�s��Kı>�y�'"X�%����i��%�bX7��59ı,O=�.u�&L�]�7$���yı,O��l�Ȗ%�b}���q<�c�a�2��٩Ȗ%�b{���8�D�,Kܝ��v���2Mݻ.�Ȗ%��"w�w�8�D�,K�����Kı<����yı,O��l�Ȗ%�by��LΛ�n�6\�ٹ��yı,�{���bX���w�q=�bX�'~�Ȝ�bX�'��ݧȖ%�b~�7o����=%�ny�!�����z�I�eFósvH��űum�+:鶱<���Ȗ%�by�����%�bX�w���,K������yı,�{���bX�%���0�ۥݷ0�r���yı,O��l��T]Q�F�"�U+�9��7����%�bX7�߳S�,K��;�s��Kı;��rp�.�̛�w73dND�,K�w�Ӊ�Kİo��jr%����=����O"X�%��߹�'"X�%����4�L�6���ͧȖ%��?�B�����٩Ȗ%�b}�߿���Kı>�y�'"X�%����i��%�bX��l�ri���Y��nf�"X�%��w��Ȗ%�b}��dND�,K�w�Ӊ�Kİo��jr%�bX��e�ge�#OU�76	#���^0"XKg-���#͞��Ժ�����������r�;,�ؖ%�bw��l�Ȗ%�b}���q<�bX�����y"X�'_����R>�}H����"iGJ1�$�.�Ȗ%�b}���q<��X�L�`������bX�'������Kı>�y�'""&TȖ'���f~7vݺl���si��%�bX7��f�"X�%��w��Ȗ>�ŊLG�9��͑9ı,N�{�q<�bX�'����L�nl�.ᙛ���bX�'�߻�O"X�%��{͑9ı,O�ߧgȖ%�`߻���Kı/����ݚ]�s7-��'�,K����Ȝ�bX����w�8�ı,K�����Kı<����yı,O�U?_ӟ��)�k�q���0�O7i�L5��r�i5r[�Kw����8����p�J3���w�{��7��;���8�D�,K���"X�%��w��Ȗ%�`�����Kı=����&�	�f�ܛ���yı,�{������,Os�gȖ%�`���jr%�bX�{�v�O"X�{���߶���	3Zow��oq��;�s��Kİ~��59ı,O�ߧgȖ%�`�{���Kı<�{s�M.L�]ܛ�\��yĳ��hl߿�59ı,O����q<�bX����ND�,���P��
3�T�U@�s�!���M����yı,O�5�hBx�����}����ow��ӳ��Kİ� ��~���D�,K������%�bX?}���bY�#��a�T�����	Hc��Sr7[�a��E��n6�:ݖ����v���w6_��v����ɳ��%�bX7�߳S�,K��;�s��Kİ~��59ı,O�߻N'�,K�����s.��&˸ff�"X�%��w��Ȗ%�b}�y�'"X�%������yı,�{���bX�%�߭��ɥݷ0�r���yı,O��6D�Kı>��vO"X�
#�
�bl�����Kı>������%�bX���8i�v�Mܻ�sdND�,K�~�a��%�bX7��59ı,O3�w8�D�,K�͑9ı,O}�d�Y�ɗI�w&��q<�bX����ND�,K��@������O�X�%����6D�Kı>��vO"X�%��]����}�߽��ιNg[:�9u\d�u77`���s���^NM]���-�.�Kd�l�a�ݛ��'H7S֚�C�F�N��a׷l]`���{WY�+f�b�0��Z�u�şOF[X7kv�&��z񳖻s��<ʑ�9���

�ƼT$av.%,���ʸ����ќb;�`0���Q�sM�#V�h��5��;nk�a�;`ܗ&i6M��/򚆉�'$�͓L�m����$�x+��mz�רCN�k�ݝ�7-
7Qi�\: �hY����7��by��~�'�,K����dND�,K�~�a��%�bX7��59ı,O=���K�.�6f䙛�O"X�%����Ȝ��ș�����q<�bX������Kı<����7���{���?u�@��qڡ
��"X�%���s��yı,�{���bX�'�߻�O"X�%����Ȝ�bX�'�7�3��۷M�7v]�q<�bX����ND�,K����'�,K����dND�,�ȝ��~�Ȗ%�bw�'�2鹲l��fnjr%�bX�g~�q<�bX�'�w�"r%�bX�{�;'�,K�����Ȗ%�b|d�ŸK�Cvm�9���e��ے�Oh�y�{�=Ӛ�����82ݙ�4��fn[��O"X�%����Ȝ�bX�'���É�Kİo��h~�DȖ%��~���yı)�{��e�j�`�#Q������#�Q>��vO!�!\��,{�jr%�bX��{��yı,O��6D�Kı=����].L�M��73i��%�bX>����Kı<����y��2&D�sdND�,K�oS��Kı;3�ra�ɶIsf����K�� dOw�gȖ%�bw���'"X�%����i��%�bX>����Kı<�{s�M.Lܖa�	sw��Kı>����,K������yı,{�jr%�bX�����yı,O��~�I��[�aИ��2���Xt�c��v����#�'c�[�ӏ��|g�+&�tR�m��7���%�����'�,K����"X�%�|����A�Iﻃ�I�>2���v���˦�	 ��}��;ı/�����%�bX�}�l�Ȗ%�b}��;8�D�9S"X��?K0��76M�p�wS�,Kľ����yı,O��6D�K�A"2' � �D�O���gȖ%�`�{���Kı/�ϻ�ܚ\�36e��'�,K����dND�,K�~����%�bX7��59İ?���7������%�bX����ٜ�-3rK�7.�Ȝ�bX�'��ó��Kİ���~���D�,K������%�bX�}�l�Ȗ%�b_;oӳ!�
�ptGDM�Ɍ�
V�fG�Ov僸��v�礸�k���b����4=o����ı,�{���bX�'�߻�O"X�%����Ȝ�bX�'��ó��x��{���߶�2\� �hY��o%�by������G"dK��͑9ı,N���Ȗ%�`�{���Kı<�{3�M.L܅�vIws��Kı>����,K��߸vq<�bX����ND�,K���Ͻ���7���{���~��N:)B�ND�,���߻��q<�bX������Kı<����yİ?�T`���M����dND�,K���2�7v�]6]��t���%�bX7��59ı,O3�w8�D�,K�͑9ı,O����Ȗ<oq���\���έ������T������-�ڻ��,['K.�9۴��jL�e�33sS�,K��;�s��Kı>����,K��߹�p?���Ȗ%�~��59ı,K�ӿ���K�fa�廹��%�bX�}�l�Ȗ%�b}��;8�D�,K���"X�%��w��Ȗ%�bw�����nM�3rn]͑9ı,O���gȖ%�`�{���K�0ș������%�bX���l�Ȗ%�b{�{-��ܛ�d��6᳉�Kİo��jr%�bX�g~�q<�bX�'�w�"r%�bX�{��'�,K���Ι.T���L�ﷸ��{���?���Ȗ%�b}�y�'"X�%���s��yı,�{���bX�'P�D�k���,�@H ��!jJ�B1[�z���Ln� �ʴ-"V�P;�M�M�V1���+׊%Ca(%�W��p�42 U|�c��Ƒ���F�r|Ӏ��;$�B
b$0���\IC���'�+��@�WE��ՅbT�"���1	H%�?�d ���O=�s36CM�l�6W)�n�ܕs��(�Q��z��jLf�<:u��kx[��r�\�y�r����kZ���g�q�梜�0��.�f��X���j�n�z���N;r�n���EUR���0�֍J�uFU(�
v�-���u;P�T�:.�N��d��0W&�!.�X�J����T+ ���2� �h��ʍz��I�6��a�2[�N8-�6������?dl��D�G�X���j���p<х�
Ԃ�`n�n�T��-u���m9.��sӎ^C{	\�B���ώZ�'�[��,��H�@�^�b�t�6ﯨ���$l�*>��rx$Q�8+��Hc��	�E�V=�n��h�m�Z��K�O��vy'��p.3�Ű>)��(n&ɴ�։�t��5��NM$R��ٲ�[v�9sR��ݟl;G<�ڷaW99���ڻh
� ��kh���@�yͩw���'c(��ei2񘎻��3�%��Fw��8��W]�[$t�g�� <�[8���*���s3�Z5��N�r�*�Zmg=gf�q¼	DIb��ܽ6�,H�6�	�k��mk��k�$L�a��rt��X�^L];m��l�x3��q1��(]Ŷ U)9�X۳P�+���<��!O<+̭) �<&{A��� �VW�V��p�*�ykf��*���j�]Gq�m]3�m`ٕr)X)��U��U����#r�,Y�H��{N�wQ��!����r�ۇ6��zΎ\w6NZ�W����|�v�|�N�lv��nuN]�>�=e��.���<o)۶m&���EP�Z,dvثɲ�\���
�"@{3wHJ��{4誣l-�J�\v�*���.�;Z�-:��@lPu��[.��	TMoC��V�X��^��m6ʆ�B�^N�nΩuS�S�4�<ge�sWI����΂z[,c �c1g��v�ns�^�:{e���0onXZ��}�c�����.P�m�����������w8*�':����^!����`? ~@q�T�����S�I�!�f�ۛ��&CvfE����!�D���x�ACl�����rֵK�ɇ	,n�:nV���-�;����lw>�{��6��X�[mm�[% ���X�#i�BK(j�7/HЏ'l�:�m�Df�B�`�6���w;p�5�oa�lޝ�������j������۬���Fm�y�zx����5�׭����sǲ3��u�J�7���w�����I/Nq���;j�u��p���ʶ�u]��	��Ez���{������g�l;���%�bX�~�Ȝ�bX�'���É�Kİo��jr%�bX�g~�q<�bX�'����nf��L6��[�"r%�bX�{�;'�,K�����Ȗ%�by�����%�bX�}�l�ȟ�𨛉�,O���r�w.�77v\�q<�bX����jr%�bX�g~�q<�c��ș��͑9ı,N��~�Ȗ%�b}��L9����6\�3759ı,O3�w8�D�,K�͑9ı,O����Ȗ%��
 L��~����bX�'�N����K�t��n[��O"X�%����Ȝ�bX��ǿw���{ı,��٩Ȗ%�by�����%��{��7�����e�=�֗�5�8�᭔���H���P.� �rАf�nI��r�l�Ȗ%�b}���8�D�,K���"X�%��w��Ȗ%�b}�y�'"X�%��{;��InM̲n�sa��%�bX7��59� ��Q_�Dؖ's����yı,O߿��'"X�%���s��y�����q�������r���gS�,K��?w�q<�bX�'�w�"r%�bX�{�;'�,K�����Ȗ%�by���L�\��ɻ$����%�g�?�
���vD�Kı?w�?���%�bX7��59ı,O3�w8�D�,K����3iw&ws-ݑ9ı,O����Ȗ%�`�{���Kı<����yı,O��6D�Kı/����{�&��Ds`�C$���f�<��5�r%�ᘋ�n�=f��î���a.N���=�%�`�{���Kı<����yı,O��6@���<��,K�w����%�bX��?[�se�wd�w����Kı<����y��L�bw���'"X�%�߻���yı,�{���bX�'�ϯe�&�6�wLܷw8�D�,K�͑9ı,O����Ȗ	|b��Q, Hb�P' ����~�ND�,K����Ȗ%�bw�v�᤹��n�ܻ�"r%�g��T(lO����8�D�,K���59ı,O3�w8�D�,K�͑9ı,Nn��$��	""p���}H���"��{���bX�ʤ}����ObX�%����Ȝ�bX�'���É�K��{���e��m9������t��M�����B%7;��'a�ם�k����y~��K�2�I.�ۙ���Kı=����O"X�%����Ȝ�bX�'���É�Kİo��jr%�bX�{���&�&nC2n�.�q<�bX�'�w�"r��G"dK�w����%�bX7�߳S�,K��;�s��Kı=?oۓ,q9�
�����oq�ߞ�ó��Kİo��jr%��ș������%�bX���l�Ȗ%����2�6��T$�	�/���#�G���s�߳S�,K��?w�q<�bX�'�w�"r%�``d*,_�DC6&g��O"X�%��gm�˶鹲m��fnjr%�bX�g~�q<�bX�����"yı,N���Ȗ%�`�{���Kı=��0��m�q�6�kE�-	�dH��i�u����4c�+F�wkMk�8�p��:R���D�,K�͑9ı,O���gȖ%�`�{���Kı<����yı,N����4���]�w.�Ȝ�bX�'��ó��?�c�2%�~��59ı,Os�gȖ%�b}�n�g�����R>�����'l$���O"X�%�~��59ı,O3�w8�D��F"w���'"X�%�߻���yı,N���t�˹$��73wS�,K��;�s��Kı>����,K��߸vq<�bX�%����Ȗ%�by���L�\��373rK��O"X�%����Ȝ�bX��{�|?N'�,Kĳ�߷S�,K��;�s��Kı5��w���v��oۓ-�;nvx{^�i�b10�dC��v�0�W�9m�ض�L<��!��8���N8�{�wQ��y�'���kF��ovf�t�gј�SqkT;���,�)������䫲�A��<6���M`P+��^ƃ��Ō]�xݶ�n�˭��+���yђ;WI�۵`&��Q���&v5�2Wl�i���C����Ӝb�nYd�f37����Ls�<���%�/K�]a�%�:v����[RY���Sbd�I��0�3l�G��P���D�,K���;8�D�,K�{���Kı<����yı,O��6D�Kı<��.N��vf�ٻ�.8�D�,K�{���Kı<����yı,O��6D�Kı>����7���{����ߠ�.�h%�Rr%�bX�g~�q<�bX�'�w�"r%�bX�{�;'�,Kĳ��u9ı,O~��̚\ۥ�ɹ�w8�D�,K�͑9ı,O����Ȗ%�bY�{���bX�L������yı,Oߋ�.p�nnawmܻ�"r%�bX�{�;'�,K�����Ȗ%�by�����%�bX�}�l�Ȗ%�by�Nws,��Yrfm�[2]��/
��wn���=I�Y�ԅ��gM��
N�̆�q��w�{��7���{���Kı<����yı,O��6D�Kı>��vO"X�%�~��~�.VSb�,�ﷸ��{���<|�]��_��!Y
H[��VB�,K߻���yı,�{���bX�'��ntɥɛ�̛�K��O"X�%����Ȝ�bX�'���É�Kİo��jr%�bX�g~�q<�bX�'��ݓL�K�0ۻ�n�Ȗ%�b}���8�D�,K���"X�%��w��Ȗ%�b}�y�'"X�%��~9rt�۳7f���sa��%�bX7��59ı,O3�w8�D�,K�͑9ı,O������������ߡ���fΆϪ�㒇���q;�@QS�䋪cv+"���Հֈ4��6��3759ı,O3�w8�D�,K�͑9ı,O�����{"X������Kı=>��/�4��L�ɹ�w8�D�,K�͑9ı,O����Ȗ%�`�{���Kı<����yı,N��˜4���]�w.�Ȝ�bX�'���É�Kİo��jr%���� �	W���@@@(~DOD�}��9���yı,O~�Ȝ�bX�'�>�O-3r�.iv�É�K��>��59ı,Os�gȖ%�b}�y�'"X�%���s��yı,N����t����nmۙ��Ȗ%�by�����%�bX�}�l�Ȗ%�b}���8�D�,K���"X�%��v���f�Rn릳^Ӕqk�#�l��7��[����Wu�u��w�ys�M.L܆dݒ]��=�bX�'{��"r%�bX�{�;'�,K�����Ȗ%�by�����%�bX��ovM&l.��n�e��'"X�%���s��yı,�{���bX�'�߻�O"X�%����Ȝ�bX�5�ʴͧ"�����¯���#�Gԁ����Ȗ%�by�����%��a�2'{��"r%�bX���?N'�,K���~~��wƋ��	�f�}����X������%�bX���l��'���g$�)�Q`�w��'��CU�R�Jr26�v{�K;���;>o�e�偩BJ��O	\�ԧ��؝�99�F�հ�N8\�i8���zk{�:����~���U���Cq�R%���_��������`w�4�9��N��n�x�,�!������Yu��EF�J��޽�M)JH�≸�-�v���6!L�t��=9����5©1�&�i	�`w�4�3�4��������`s��
Q�����,	��s���e������@H�-�'��s.i��isKȑ����.ٶ$�3��mú͔Ũ7N�H�.ܢ�GU���\������.�����l�î�gI�7S&_������m��O\YR���h�*6[�����˫zWD���c\�"ݘc�p��h�=K/-��H���J�9Z��1�wRc��dL[}]�r���:4����s�.l��[m�r�ӣN��ww���T�4�Oc�ѹ�M&�m���n�=&n9�������\�i�=�W]j�@]��:�r�18W�1g��8�5��M,�M*��ԍ��I%6�8�/�ɘ�K����|����[m)RINFFԎ�������Ҭ.��s]��[�wR��t�Dj8X|��w��=9������aBJs�`wվ�t�Q�	�Q8U����`w,�����z*q���Q�U�f$�i�M��N�=bܵ�(�L�]�sw7S��Ɨ#uOB#��,�6����[�f:��f;�b��Rm)O.�[.nrI�og8���@=�vE��GG�W�`vs,�����<���c��m)sg��8����.�=���Y��-F�!q-3Q�s���e���S��F��R��rSn;�s]�꥘�N��֊�;����#ə�8
���f��`GqnK�=�7=���]�ܳ
��%N�B�TT2�iJR)N)Q�#�;ܚXܚU�s������`fV�ԡ8�-X-Ũ`OEN0����Yu��E��ﾤ�����6�6�9J'P���X���{&":��	D�('"H8H�B9��$ϔ#(> �X�X���}R�VReHЅe���F�]6�"0���D=N�I���22�# ��S�E~萨�9�IJ�La����)'V7���\��a�|����]B�9��y�I�%����J�{�Bbq5%�fo�HFB��<�<�j�O�TS�>,^��x� ڴb@���H��0"}��}�P7���@���F$)`��DO(@:
z�"�TC�C�a���< �QpH���H��"�UC�b��("&!��DuD(�̪�`g��,�4�4��j]E#rX~��ﾥ���36x�3�+K �we�νOi��b��E�v����	㵧@=��`v^>X�w�{}q�s�+بij�"�C�����)��#l���n:m8��ٱ�L��{)2�;����|�%��ZXͨ��H��H�H������������`g��/aDGСDs�����R��r1�,_����M,�J��9��`r��m��$r���nM��e2���L�����K�%b�B$�X- 2Ա�,-,!X��`Ј��#`�Xa}	S�6�^I?~>�ԡ8�)�G����?}U�|������V{�K �K�n*J��q1��Z���ʕ��vX}�X;��7k���,��g!RS��Q��"u �we��{���ri`wrV����)H�u#�M�`g^�W�_$fl�`g�W� �we���;����)6)�$I�`IW��.Q�w֦�ی�eC���C�iHXܕ��s���ν�a��}���}�Ł��u���%E�o�;�S{m���r�H��
"���?p�w1�ˍn|у0/Xt�N���J�WN���V��:n��q��z�Y��m�k�mpr�sl툎]��Ň�y1q��;Cۍ�n��{ $m��H#�kC�n�1�Y�dŬ;<Fa��8��a�q���S4�'�R������z@�6�r�F�1t�l��B�	�H��,�#�gK;�I�];r.����؉�]�nm4����Q�g'<�廐�7I)n[�s'N��J����ﾓ#�\=n�s-1�#:n�`��E*H�#��f?��X�M,�J��9��`s�Y�����r26�v����!BS#n���ݫ��偙[�wR��tH�j8X�+K �wj��"!)�N����u��֛9k���qr�B�9��`qn�;ܚX~���[�u���?P�JRcS�bnK�m��E�0���;�ss~�ۮla��uu��ą"���r��u]��	���W�]�θ\V ��~����	"�}j`w-���L����˷-&n̷vrI��i�ϔ�A�|��P�s�y'9�7�Oo�ߝ������)ֶ��u$d�'P�����[u��EF�r�.�pR��r1�,-�v{�K3%i`��9�Y��"G)��ڑ��S,J!�kN�{7j���`�{������s2�G[��:�'9���Rl�Rwa�3��b�(x���Hڷ��tj�� �0;��`zEK���t�J0�¬��,�o��)�fS�	B�78�:����Tr6��������M,�}�p��`ӇU1 \G<�|�a�$�we��z��%&� �Rq�̚0$��`��r۬��x.bF������J�?~���y�ߧ@����`w2i`�Ě�Ӎ��5$B�h��J�ٮs��Ļ��0�{m�rѻ];U:����I#I¬��,-�v�T`I(����ƌ\Z�n�Zn���[u��E�0�S��?Wԑ��W���G)��ڑ��<XE�0�S�m����h�X	n-[�`I(�;-L�Xo�~�@�	@G��_@�� =�{�����t鶈� ��9����%�	e}���v�,̦X�ɿ@�-t B73]:�"�b�89��LU��u.�̇ vժ�ظ�u'C#���m��T`Ie����=��Ԅ�H	�`w2i`fd��9������~���ֵ��R�Q4���UQ`6�Հw�>�
gӻ��3vx�;��%&⨥G#JJ�f��;-�X̦Xl$�[{�`kٕ��)R@��ܖ��}Y�~8omXq��1G"�P�'�,i:��ruul�ä�n�[��eN���#����N�AQ��')��:cZguu�l�\[V�nh�|xM�rs���r�l����x�{f�=ۓ�z��Rof�Ě�k�+3�yC.�:�m(J˱��Z���Ȣl��nò����u�9Kø��{\[U�n�F�E��n��l�8�ұ\V'�Y ����7 <�e���0�G�Ǡ�T����qF��7b�v^�]�l�����g{[id�d� ������f��ƍ��Hr�`fc�`���"!vCӻ���xN���F�����ͺ�f�8�u�̚_�ꤎ�Ǔ�t�D`)@UR�=ڰ;-�Y�Q	$�q�����]Xה-�)1�TN4ے���u��J��;-L͹Q�cR
@n;��K�V�����,-�v\�bf�*���SDm>��m���\�9��V�}��ٙ=�f��ܼ�v�HR�M�,�۫ �n��w_ꪮ �����|JM�QJ��$Kt�y�{������b�H� ��$a
1 "�B!]�-�X�2���j�x9MZ��I6�crX[���M,�T�����;���9�V�lh�Jq�6�v�T`I+� �0;��`IK���Q��736��9������`w2i`s6��4&H��҃������XE�N�*r��WK�YgP�ek����}�v��l�I+��zX[���M,�۫z򅴥*n"�q��L�X�T`I+� �L͹�q	�H9J@n;�ɥ���ud~�'X�T~AQ��QS�f��X��;��͢Rp�n��NO(�31ڰ���;-�X}���zX�"��BBH��`��;��`{�Q�$���(8��0gC�z��S�Sv���q;�ETO�sV���XR���j��	F�crp�{�����I_}j`v��q�pX�s�W&������BP�S#omX�vX[���&�58��p�31ڰ���T%>��偘�K�֧lq��8�IV�����M���,��������P�Iv!	Bq�\�wVq�iJT�J$�Q�,-�v�J��;�S�ӗ6��f��i�����\�װ\`N�)l���[���sb���R��q	�H9J@n;�ɥ���Հw��С%��?}�,[���iMB�ԥ����u��H;���:��;�ɥ���H�|D97*H9ĸ�=>�0;��`{�Q�$��h7jФ	���`qn�;ܚX��V�K��K��|���'	%rj�`{�L�/T(I��^ Ǽ�.sﳒO�Q��Q��DEE�Q������"���EE�EE�A��  �AP!PP$E b�E `�E `�E�A���Q@�PT��/��Q_�EE�(���EEh�*+�(����Q��DTW�∨��Q_�EEآ*+�*+���
�2��!tp'���@���9�>�a|   � �                 >4TH     P�  DJR��� UIAE( ( E 
�   $   E   ����P� ` ��)6 ����	 " ��(�� }9��>�ﱯ�μ �&�����}�"��y��sw���k��ҙ5Op о�����ɮ��+����� x>�P( U 
 ���}�O}�^;���,�����=9:�q�s���x�t�x ����j\[׀��eV}�#��S�u��qv{zW�ri]� {���w��M\�=��� �    `  
 
*�
)��  �oe9o����n���{��� �zk�WMsi�n��y�ꗼ���\g�ն�� �-{y����� {�jrz=\�U1����,��� ������k֮f��'W��� �   ( 
)� }�����������[�^� ��;WM�sɸ����,�N>���^۝�{:xڼ  ���ۋU[� �t����[�q���]��&����>�y��f����k�+����ԯ�w� P   PR���ϩ}����������]{o=�]�Ӟ�b�iqg���\JP /�()D@ ^�P  R P   ; iI� J 3J" @4h��$�;4 " ��f �  ��MM��*  S�$�3R�� �<z�R%   D�*���� �T�Д�R���!����"Be%$��2hl�B��o�O���b����_L�̧O�ڇ�ǋ��DTW��
"�� ����Q_��"���EE`�

����_��`��|_���Bj��������b��)
�]�%��ܺ�z��N|��e�����HFq2B%W�@�)S!
��cJЩ�Si�4���l"�y�h��4��:u�����4|d0>R5��h�HEv�zh WZ�$X�pt5��"h��a�.�S�>9�\�K�!q%ĕ%0#Y]��l���;W!pى���ӫ�FV��	t�&����0�;w��i�%�(@��Ą((|�(-4:p"SÀ^s�Lѳ��x�]�@�a�c�F��1`�s��o�D�H4 �F��Ƅ"c@�XWD
�SO����\�,yϾ���T��čqӶ�iU��Zc$�l�L::'F S\+�A���i�4|�%�4�)��W��	���>Mé
�6t1`��1ѷ��iCw>����kJl�)*JB�F��`Ј�"$i
�FD`51�XРF�$&���h�A�
�$�)�ST�V� !B5!�/7y�4~A?�c �y����ɺ!�
0� �'�%��6��H�1#]f�Mk��3Y϶K�&��)���4����I@ł��1H����
�i@�!�����[�FI2Bh��%I-L�LIrS#X�	BR0�)�C;���;�%�o_j�9Rd�ɯ���w	]B�(@ D��7�fsv�d�.W}�a��s[��N�H����ѷ��7;P��ya];`��4@aSd.u���y�V5��Ww>�GY�����޳[eH�S��P�͞���!�\hZ;�T��
B��NK�%)�]���-i���2F��u��V�i�K���>>aS���\ֹ�9�pO��l��ī�w�sS2hu�.��r�5�F��@!���ل���p�}���.0���V1�8ov��v��%߭�v;�o�Jc\8ˬ�ˮ쳐�s㻅��\Ѿ\���f��\� �m0�B�LJ�)s4$)��D0��y����ek�x�XЫ
T�j� c�tš��57�qs������4��V�k	sD�6�H��#�'�����¡�HC�x!GW� A`��W���v�C�IL4X�|�:me͒���^�,+��6��7��N:7�٩������9�t��k��&����
f����5��A�]w�L��B1*ƕāT1!\M)�@��s�s|538$hň`�$(u���f��nrl�BB�ַ���I"� QJA�[3Z�3[4�aR"ɲ9��Ro@F�ZH@�1B8c\�1 ��Cla.km����̙Ϳ=�a�	T�	���HD��H���Ǜ��=~�2X����V����� �ġ���aO��)�́C����E�A��(|��(� ���с ��M�����eE���!B��a��܈A�
��-C
 D`��-+`՗揠@���&k[m�ӆp�:.]s��d������	��
�,I��Q�@b�H`5@LM#�5X�dT��~�uC���$��)�R�I��o7C[>*��H�%H�W�
bB�H�Ā�Zb�i�֦�k�޸�!u�Gw�f�wN.��B1Ͳ����5��B\X�L+�֭��p�A!�W6K���_}�p�%YBVa�ič T�4|�bK��|��~����f�V\6�M�R��w9��0��Z|C��7�?\���d�= �� $�w5<��V#"C�B$�"� !���d3V6F#5%tZ>t�8�Go]�|�F0ӷi��Fp46o�-���;%3[TbG(`�rP��S./�ti�N(b44A��J�f�Z)u��I.��ē
ai24ąlI��	$Ϻh�hD�	��� �W,J�:B3|�gM��Iq̗\�'w��� 5�=����p%V.���.��,I��c�e�"T��,(a�����8���!�@�0t�j`iH0Ѷ\u���a���%��(�#0aX6˳M`4���	HS	B^?8kl p�a�7ޖvj�R4��S�3>��TvA�C�>�@��@B��ӿo{����0$G���_�H�^j��.��g��e�FjB�+��K�)
B���� D�)�F��
�浳��9���XSx� B�s�]�L�5��L�A5�P�hѷ1`�V*qѭ��6o7��ݛ�a3F��q�D�D @Ӊ���0�H�BZ`�dJ�V�l����e�nFT��m����B�H�Ѵ���M
�#�i$�����qXA�1ц�b�4��)���ɘK�p!K��D ȱ���{�l���.ހ�yy�B�~�9��ĖϏ�k�M�l�t,�4�c!
`��m4}�fh;M0�f�[��Kb�h�D�2�F�#C&��Ґ��~:����eލ�Ye�����3M4�"C����I��1 �cU�L�$$Z�M��!F$`0z�-���B�:]�1���ѽvd3F�^x�$�	��١cA�C���h�B�615#\�41Gn�]kn����x�����Wv�6F淿x�� ��hڄ�C`ĩ�����*B0�l���{���o:�́!s�>;�B�
0�B��])"I�BK�Ѱ�C@$B�M��ȑ�5
Bcf7\��	���A�B�=e��_l�ގc�S5����X���"�� 1h�F��*ZB� D����%#N�BI�1Һ	\֩�S�ޢ��D,�$�
����@�5�K
kQܮ+"�&�$%���t\4�al0h�@�1:��5��Cw,t,��H�Z�i��i*}��,����|�T)�4l4;O,�`qcLtx��|漀���$LO���!04l��4L`W��4�|`p�@�(@�@���F�H�0!H0�4+����W@F���7.�6B�����>aM0d.$F�����Hm5�@�5�i����H�� �`A�0�!0��ĸ�K�!ew�
@����c
��H[���yu�K�.����4w40H\	N����!q"A��LMB�&h%�$A������1����L2$e0 Q �
hB��mX��R�֭��a���rMp�Y�6_�7 �k{dǺ��B
���:����4�w�+B]kvg%ɮrl�5���� ��D�P�U��T�R�(,�51H�4
	*�:��,c��|�Z$iLt���W��y��;���!�*c�Q `���3F�|��no6�=O�RP�S/M����ӭ��Yts�8u:/���s�Zp>�%ˠ����CZ�����,5�S]&�&�xe�ﶜ�L�32fSCi
a��RYBR\��>��|8Ԕ���̶@�.��ԣ����R�X�P ֓&D�|hb&����d������P������O{;��5E�2���޺>	k_g�;(="��2t�bA��4Y;���3�{���}���;�]y;���   � �   ;Z췅��d�1�g\TRᲷ!lVcW:cm� m������$ m� ]�M�d\ ,0�$����$Z ��m ��m��39�0 �m��n*�R�y[�nn�6f� ke�\  �6�!oH�[�pvm��N�ޠ'�V�����:�T��ϫm�s6�]��U�e2�e�MC����'nUk��)'��j��USWm��j �5�]�����E����z��趲��0U@:�z�&c����7��
wg�79vՒK&��޿ݹ��np k��m m�   -l�鴂@[x-���#�I��t�n���{j�'8�q�@���^U��<ײ�ҭJ�Ҽ�M[tP�k�$ ��۰	4Q��m����m�  I �;gZH�m�m6��H�x��cT�-6� ��h巚���/��� �$��ls�V�   ��m�[^m� �`�ְ[�  � -�� �l��p p jS`�\�����n��mm�ڴ��b@ 	7mfe������$�h����h�v@	�ĉ$ ��m��8 j���|q� pd�E�@�h8v�	8���N-�lms� mn�%�	 m���U� m� [lH�l�M���-�k��  ]6m��  �   N-6m�c�M|mm�rN	��� �[\     h 6�`�@6�p>	>�$6�  H�M�6�m�����hH[dԉf�pH2	-�۱�$$�Zͻ`&۷ ���[M��6݀���
P  �m&Am�  $ ��� � [N[�K/  pm$v�L ��o6�p��h-�hj� А �J��p]�P$UUP$�[���[�ζ޴   >�Y��o�� �k��:�մ:M� �b@�lm�i3m�ݵ��m��㍤�sm��$ �+v5�m��í�� $H�Z��UJ��t	®�V��l��N�F�Z�ٶrE�d�		�m�����vw`%k�� ب�����9�^`���������i�O��}�ݶ�&�VNm��Ͷ��4%�:il�k�wq���pA&Y�	�-� l�I����][`6� �!%��l �` �J ��x ��F���8m�q6��f���	   s��Z��d�MgJ�l�H�vߟ}5�]6� 8�t��$  �u��I#��f���	�6�m� pi0 	 �'[]�lkX�m�]6qm  im�m���l� -��(m��  $ [@ �!	� 8i����&u�J�oK: M�6�����C� ���v�X��I �i�� [dH i�e�m��2-UU�Um+�J�R0T�d�#u�s�5T��V;N^ vp��z�V� �P  � [��V�vS[p�j݀ 8�qS�����2�@J�T��
� ��[WW]��j�������q��TN:mp sm�PhYV�������խ��J��V�8��˲�]P�zm f�`[Kh [:]�v�@��jݱ�-UR���TJ��&�m�-�䲀 	 9��mج�:@֛v�U��+�L��Y��Rey�]3���>����*Ʃ�����j��VV����u�����-��V���X�6�V7`W����n�A;eSQ�ksʗEm�U/,�UR��4S�j�N�r�OF5��@�`�Km������y�JPl@P�*�l��,�pM����t^-��܇V���ѡ��UJ�0�dP{\�@��ەj�`�'I�4�Ӌ�	��Kh qml�If��͹�m�3sL�$Ԁ����[m%�W,z��k	�pH�EF՗M�	[`��u[WT]�@tUɵoI�5[� H	el2l�r   t�wү�y�;��Y;j�vse�ٯi9k [dHH4ڀ 6� -��t.�H��z�۶X��{4� $8.�M����]�	-�V�m�m��gk�+Y�;m�M�@ ۑ�  m���p��I9tM���D�-�ۍ��5��lm���� �   q�m�Ryؤ���P��}w_���c�I�l
�]��S�mUҮQ8k�$-궃�F ��m���>��� �f�ʱ��U��ޤ��r�-��z�P6,��@U�[W\H�m�lnٶ�d�հ/[oP H� p H  -��&�
��	V��%��:���ccl�Wf����$�lA#�I��j�8ͷ`m�@ �u]UR�V����V@%� l�!���n� !m�� [@n�L��Sm�6�ѥ6Z�i6�r^�ր�H%ӯb�À8ZVĀ/���V��vZU��)�Π�-� 6��Y��Zݵ� ��}~��Ƶ�X�i!Ä�kn-� �T�R�e檔���9�ޒ�ٰ�� ڶJJ\/Z�86� ���ŵ5�ZΈ����ڭ��&�ά���9T0�pardِ��]mUUV�2u�yD���ڪ��U���nۛzt�7D��f�l�#�t��*%yj�kP�R%��h6�:��m����` �  )dHHz�@ඝ��@9,�mm��c[��i�$6�ӵ_ lm��/�jF X�$��[d=�)�+j�d�\�J��h m��  H[x �'9mm���.t�.�mͶ����ձ��     �  �X�$6�5-p[Wzk�M#l  �ˤŸ�j����А�UUpA�* � j�uH��n��H�� d�m��:mm�$�&L���mUE&�p�q̥�I�I���"�s�l� 8��[@	e����$�$[@u��QbF�h�6�)��p !���LImp*�؅'����n�u�K� � �p�x�޺_��$ $�: ���K(     0� 	��F���$��9!��m�� m�R+mm�� @mp ( ��ܲ�� H      ��Y@�I�$�m�l�� H ���  �����m��)-T   ��%��-��e��� Ͷ��� �m5���i06Z����
�UR�F����Է��$�H�Zmې�׶4� ���-��     [@>s�o���)l��	-��� $�mڶ����$ �  
Wh�[���lR�/:IZt�_[�����m��m�6ZH��m�k ];��5��崽oe��K�Ԁ(����V�`�H��j�C-�lWUP�Km�������z� �턋W����k����[��B�d�F�-�j�ګn��;guYL�:)�B��X]����� -�Ԡ n�m��`6ٶ��ճm�$�6�q�ݰ�a�ӭ�n�r� u���$ض��8kv˰,v�6 t�t�-'a�)Z�L��ڲ��!�n�M�*@�E��	:9m�`�Z��s�Z6�b۶pv�7Z�p6�%���*v�f��v�I��А���9mn�6�� 8�v٪�V�tyV*U���P��K���6�v�Yb�mM�� 6�X   	�`I���mz��d��f����gZ����M���� -���6ض�Z8h6m� ԲJְm$ص�m��H   m��f�h���f� �H K(�[M��`[v�@[~� p9���6�a!m&�rmp6�Ed�	   9�j��  �m� ��A�|      ���&�l -�e�B@ �  6��`��-���  ��9�Ŵ-�mۀ $kV�t� jͰM�[vޓ  ��6� v��h�[��� [@ $  �[I�� �V0 �'N6�}��}���'lݙo>n�m�q'-s`  k�� m�](t�޼  ��  [m�>w�}��&�&vն  @ڶ�u���%�m6��[W��$��m�P*Ӳ��S-k��u�2�U,�	����,^m��  Ӏ6��n�߾$e�mH-�t�[@  ��p  �5��  m�mIv�ڶ�-� �n���lv�[ C`� ����m�� ��$[�F�����*���yxG
�V�]U*�f��R�k)�Lݥ�8�/+�F�S�y���_�]�����R�"�X ���
;QO���hmC�N*Q���r>D�=(:
M� �
Hl>p�^8'�`��I(�(M�O���ڂ�
�ʆ�S �.���LO����S�������	��<��<��G�|^�A~ uWq�H��? )H��N4"�¡�צ��~M
hP"�P �T<���?*���	  H ����E:��DC�~� ��h�. )���S�H |�t (�}�uda� "1P`��M��L�@|"�6;�y�6"pD��"�T���F|'� �
� ���z��C��</ʋR"�"�(�b�� ������T<���4R*F%�T�����z�����X�b 6tS�j���<����T]j�B��ʴ���DANT� ��Z���R#� ���ADTW���@? �@>�k�ѭkZTvS#��n�M�F�U��eá�1#�Wv��'�'vwa�M���c7Z��ŕv��nv5�%jչ�̼$nG	�u�VȞ� ��x�W���kN�X�#���k[N�^� i
�emlm VλB<�죠�tI�q����E�Z�;X2��L�m�uU�S�L9jL����pUT�/l걇%[��`�m:I�1��9m�j������2:��3�n6 z砳�7V�rEER�gf�����WJ�*u���JuR::C�u�u��,lt읩fx)�]u�tF����h�=��.�Dҭ[;�� �|>]����A4��T;E�g����Sp�G�Ȗ\[��ŕj��P��6�.��Y=��;Z�h�;H�)hW��c㋞�Q��h�rݹ���;Ǔ8��t��:��nz�;v�����l���Vu%��<8�xŲ��R65�ݵ!���K@`��퍠�����3�49r�{[����l S]�rJ*nv�]�����iН@n
�$�0U!=*�Y}��0���cAO7P[dt �f"�Q�`���Hh	�eΓt�lf�n�����z�q[���Ə]�"H�l� �e�Mm��e�Ι�Z�L����)��d��\Z���W92[&t=��/um����\ۍ�yg;m�,C ��`�eV�qt��=�8ભTClp�[�4ʶ�s-[U��6օ��n��B��d�a�����u��%Үt��h�l�x(
����P�[m��6�ܻ��y�L��mV�Jl��:�Ě�k�k���;���G��K0m�L]�����R��x�-۶*��֓$�ڱ�]�q箪�ٵ�ݱ͖ڶ��\ؐNr��9坵�]	wLn�ݖXv� v���Z0�ݍ�B$G����H ]R�+�0T�I^Z�ǥ]��l� t�M8�]T ��7;��V5=I:���{j�(ʲ������r�q�w{���� ?�D�l� *�D�#Es��{ZS�'	�ns-�!�7yv�<�u���Ɲ�������Ƙ�$ �n��m�g����ƷWYCpl��˷;q��=�<�v�6�ͧi����-�8�v.��t璅yk�뎓�ɷm�뒭l�ۉ���[rە��bT�B�u�(U�&N�����]s�JƓ<m��A�:C;I�&�e�Q�9۴�y�d۶�ݘ쌏JN������u���3[��6�e��l�rY]�`�v{� ���8�32I�d��fr�csX������$�H�}{PI����������"X�'~���Kı/|~��)��&���w�{��7��������P�]D�K�߹��"X�%��߳q7ı,Kώ�[ND�,K���O��i]u���=�oq���X�ϻ��r%�bX�{ٸ��bX�%��}��"X�%���{*n%�bX����h��5��5���5��r%�bX�{ٸ��bX�%��}��"X�%���{*n%�bX�ϻ��r%�bX�=�ssR[�k&�.����bX�%��}��"X�%���{*n%�bX�ϻ��r%�bX�{ٸ��bX�=���~?�z�6�"�9�Z*��ֳ�m۫[9<6�q�s��v��sجX��	��ֶ֚��bX�'s�쩸�%�bs>�iȖ%�b}�f�n%�bX������bX�'�te�.h��5�ђ�k*n%�bX�ϻ��rEj� �1N���pH��0 	1pD*,�C4��|)��'"X��sdMı,K�ǽ��"X�%���{*n%�bX���e��a�5���f�iȖ%�b}�fț�bX�%��}��"X�%���{*n%�bX�ϻ��r%�bX��[3&�ѫ�\�7ı,Kώ�[ND�,K��k"n%�bX�ϻ��r%�bX�{ٲ&�X�%�~���W35-�kV�5�ֶ��bX�'s��D�Kİ�~�}��r%�bX�{ٲ&�X�%�y��kiȖ%�b{���֎;����]B=��^G�� ���s����݂�����Wa(��92�3Ow��bX�'3��6��bX�'��l���%�b^|w��r%�bX���Yq,K��Ƕ{RkFk5�kWY.kY��Kı>��dMı,K���ӑ,K��w�ț�bX�'3��6���F�5��~��o,���h��Z"n%�bX��=�[ND�,K��k"n%�5�Ć$��A�`Y�vn&D�;�fӑ,K���͑7ı,O�;���V�շM���ӑ,K��w�ț�bX�'3��m9ı,O���q,Kļ����r%�bX��їĹ���ֳFKsYq,Kļ�}��"X�%����"n%�bX��v{[ND�,K�׵bn%�bX��ǽ��3�k)uN�6�`�.z盂%Y�vW��, ����^�m����f�+Kq[*������{��"w���q,Kļ����r%�bX�q,Kļ�}��"X�%�a�zj�2j�֍\��h���%�b^}��m9ı,N�^Չ��%�b^w��ӑ,K���͑7ı�{���~q�
�j	��������,N�^Չ��%�b^w��ӑ,iZj&�w���q,Kļ��m9=���ow�'��]gV����%�bX��ﵴ�Kı>��dMı,K���kiȖ%��S��P2
R8����v�&�؂'�j&gߵbn%�w�������srS�_{�[�oq���͑7ı,Kϻ=��"X�%���ڱ7ı,Ng{��r%�oq�߷~'�V�n7nڠq�Wv��t���.�;v]�Mt�ƻHs�i%?7}��^�d�MjK�h�Ȗ%�b^}��m9ı,N�^Չ��%�bs;�f��O�dK���ٲ&�X�%��O�L�����SZ�r%�bX�q,K��w�ͧ"X�%����"n%�bX��v{[ND�,KӺ2��4]\���d�թ��%�bs;�fӑ,K���͑7ı,Kϻ=��"X�%���=jn%�bX����~k�in�³�������ݻ���~��"n%�bX���~�ӑ,K��u�X��bX�%�{�m9ı,K��T���F���.f���bX�%�ݞ�ӑ,K��}��ՉȖ%�b_����r%�bX�{ٲ&�X�%��OC�`��H}r!�F1D`��`3U}�Ö��u����A���65+v��lj�)����n6���y�v�n���/:l���] cnu�n��݇����^�p:��{Gc7�ێ���Ƶ����I�H�cM�)2=�Mֶe2l�pu9j[vj݃�n�������!�YY���ǣ)�R���D��whq���u�h��!2\��W��!��Ojt���j�sOfWV���j�H�k��Yl�RT���Ѻ��=�<���/^���ۥ-)&x��]�PMV���{��7������V&�X�%�y��[ND�,K�{6D�Kı/>�����bX�'O���F5�Yժc{���{��7��{�m9��L�bw���q,KĿw�����bX�'{�j��K�q�߯����錴�D�W�����d�>��dMı,K���kiȖ%�bw���Mı,K�����bX�'�I���)0ɬ�ԗZ�q,Kļ����r%�bX�q,Kļ�}��"X�%����"n%�bX�w�{��\��5��SZ�r%�bX�q,Kļ�}��"X�%����"n%�bX��v{[ND�,K�Oڗ-�9sN9���n���N�^ŷk�)�p�Z�כV�f�F���VnK�Z�2]f�%�X��bX�%�����"X�%����"n%�bX��v{[ND�,K�׵bn%�bX���瑩f����33Z�r%�bX�{ٲ&����ƈ�P|".<�Ȗ%��9��"X�%���ڱ7ı,K����r%�bX����s&��kR�K��&�X�%�y�g���Kı;�{V&�X�%�y��[ND�,K�{6D�Kı/{<_�5�e�պ�kZ��ӑ,K?
@Ȟ��j��Kı/���m9ı,O���q,Kļ����r%�bX�2��a7];�Z�7���7���{�����m9ı,?(�����'"X�%�~��m9ı,N�^Չ��%�g������:<t��(2�D�3tj���ivȡm�8�t�8��M�K�]e��kiȖ%�b}�fț�bX�%�ݞ�ӑ,K��u�X��bX�%�{�m9ı,O�ٻd��&�kR]kDMı,K���ki�~T#�2%��k��Mı,K��~�ӑ,K���͑7ı,O���3Y�Y�Yn�u5��"X�%���ڱ7ı,K����r%� Ȃ��������dMı,K���kiȖ%�bzwD��j��K��7ı,K����r%�bX�{ٲ&�X�%�y�g���Kı;�{V&���{������~hW�nXʵ����ı,O���q,Kļ����r%�bX�q,Kļ�}��7���{��?����N;vte�8����(ܗ��θ��nSU��\��`���!͠��kfK�.f���bX�%������Kı;�{V&�X�%�y��[ND�,K�{6D�Kı/{<_�]�PMV��߭�7���{����7���F9"X��{����bX�'~͑7ı,Kϻ=��"~@ʎ�������a7]s����ﷸ�,K��~�ӑ,K���͑7ı,Kϻ=��"X�%��ﵑ7�q�������m\<� ������K?"���߳�Mı,K��O��r%�bX���Yq,K y����":�Mw^�[ND�,KϏf풓�ɭI�ֈ��bX�%�ݞ�ӑ,K��Ǻ��dND�,K��~�ӑ,K���͑7ı,����~*c��j=���Q��M�5��8GN�|�V�S��&��t�X+e[ƺB�s����$b��wvq��#�����������8�!'�}�پH���4������^�k�$�9��nM��s@>�K4.����� ���H�"ycnf�}Η�[%���03dt�7IR�
��"$J9$$�8�k���4v�� ��>X��&�8�m�*��p��:�L:��4nͧ��
�Ov���eHp�v��|�,��/5grg��ݸ�RW���
���T9{Z�F�������r���[ݼs�� ��2]�]�/{l�-����<.s�7�є$�z<�ɝA�u���ti-��v��<J����A��z�Hu�~H��cY���6]�M�'	]�����JgW�((	7w��&Jk4[)�3�cgK�aM��p'ø��\x+Y��qű0���&�.���&Fd$rG ��4v���Ε�]��\��pJD�ȣI��I0:�Il[%���0'һt@�x�ɓ�4�:W�w�է�(S'[�X����K����I��'�[V�l����:`uf����U��c�bq���-��˝+�;�j�z�XL�D���jV����z5�
I��N�:���2v��Sj$6���7�rh��h,�[v�^����'��d=����W%̗3F䜿v{7�*}6��N�h\�z-��ޖ�8�h�F�p�@��@�w���˝+�9�e���&Fd$q����k�3dt���%�3nD��Y.P���'�E��@�m��=����i���vl�1Ձ�
��6t�����T�9�ePu�-�æ����=f����uև�X���GX�x�ɓ�>����;�j�>]�z-��;�sq���L�Sp�7nD���O[}�:`uf����U��c�b��>]�z-���W�
hT|0	�Q?@M�)����؛"8	���J�!�aIB�2VPˇ�s�d�FB\8~��b$E ���"_����C��N�a�A{��a[�8���~���%��A")F~:@"��B�f�I	�|���WdQ���6⡂fJC�Z%��+������#0�j#�oF�6�E*
�Eȑ ���|��0E�C�C��1F�@ N�(?���A4!`�������9d�y�}��A��ۏC˾���-���A%�ɝ��I�`S�8�o"y#��ߓ�s�8�O=��ߒ-~���[�w�����T�~Q�#4��W��ι���F�h;�{A�-����f;8���$i(�x4H�c���=���������s@�]zs��M23!%��|L��o�$o��07n_���r-�bEY�?bR'�E��@ﯷ4�ۖ�ܹ�v[T6[Ut��ddɉɚ8���;�j�>]�z>D4@OEb�T�����x ����rNw�����6h�M/��ܹV\���c�V-������Md�*�ۖ2s{xz����u5��i:-Ľz��ᴦzv�i�[��n0���ջ-��c�e��`n\��kö(�r�&�z/n��>���ڿ� ��C乗�"Cy�$����w��=�E�����q������� ��y27(��q�^�ytRz���Θ�/���ڽ��v�L��H�-��נr��{��;�kj���7f�q	z[I7>�O
�):�E��3��p<��;+����ŷV�7$�k;��%9'gJ:ܜ�$Im�w1"-��Q�r���%F�y��Z���o>�����m�q�ٶ���Y%-g�B��H�����n�:�&!��º��K�&�	k��k�-W�r�<7	Y�\�f��e�g���Ō]�E����5�Hm�]�
�s���.���?\��ζH�7c �_0��rh��ѧT�d���Ԛ�!gr�Iy]g�P�;Xγ�WXQ`��9��
n(��t?ߗ?���h������-�q��{=|��	���193}���j�y[��}!�oj��׿+�f�nA21LIG��E�����o���۹�s������nc#��_�v[&�L�ۖ�ܹօ�5��n!6��9{w4q��7.D��ݖ���J��\*���cS^M��RQ,9ػ��!/�~��״$�;h*,�Cy�bNg�w��=�ú��:�J}!��Հ=�٢xs���֮�&kY�ܓ�g�wT'u���������}u��bEˎ�m,����Z�z/n��ؗz���/_���-�&%"x�Q	��]����-��r&V���[��c#�����s����v���נr��hrפ�2D�4�?$Ԃ������<��;j� �A����4���b�e���i)�QǠw�ՠ|���^���}u���ws!Q�@�ZV�I03/n[v�L	-`�b�A��ۏ@�s@�]z\��|O�>j�'��}w$��}��Ngn2�y�$i73@�]zz�Z˽�@�s@-�LY!�"��G�޻V������;�{s@�]z���޹�K}&,aHII�����f=��g��v��ӭЗ��#�tÒ��P�1�q�_�o���n��>���ڴ;�X&5"x�Q	��[]>�e�ܶ�Ș[����n�	��"b�f��>���ڴ�{^��n���]�1��	G��r&V�I0�j�W�N��l^�?`�!Q�@�Z˽�@\����>���ڴ�{SI��nph	�ۺ6{i�Ī��W��, ��뀩xx�:#���G�G$�z-��8���;�j�>]�z�v�.7�<q�;J��̽�lۑ0:�e�2H�[J��D�"��G�޻V��ݖĖI03/n[k*�R��\8�F�����{^��n��λ4�ڴ;���i��!9��n���S偙Ḿ��:�*#BO�
��`s#�.�zc��6W�i�*����{hا��xL$��5���y�i��5ɹ띞ۚ�4�@���]������R�vV�Q*�G��֍�m�n�h�'\vA5����K���7�y,(���rHnv��m���ma��z�MqV�kG1��fS�L�����S���}�=��]x���pD�S����JN�j�x��³� �P�w{�w��:�����;k�:=���E��dۄ;v�Vw=H��N�M�2H�����x���:�_��޻V���k3Pr۹�s�WBF�iJ���K�H�'�����01fܚ�b��B4����z˽�@�s@��]�Wmz-�'`���$�ӏ@�s@��]�Wmzqۯ@��[.7�<q84�s4.u��ղ[�v[$��Js�+�[/H�MĮ�F��8^���=�{\ַ\:�>.�r�Ԓ=-��T��o�����V�I01f��k*�R\�kVܚˬ�fk7$��}���b^@�ȶ�?:j�R�@`t%��:<�������9u٠uv׵ �n�&4�bqD'#`d��m�3�_RQOz����.Z+��a?8�)&h\�@��`}9��5%9��+0{aʪ�s���.P._8�ղ[�v[$��������4�-PA��f�0�ڻ	��+�1pF�շ����:E�>��~�TdiG1	8����[w4.u٠uvנrقw"M�)14��9mt���e����l��l���*�"x�pi��h\�@��M��Y�$�DJ��Wf�Ձ�nՀ<i�L�x�&�l�94����{^��n����4�1ܸ��&F������l�:`bų�[%�;/n�t��ɤ(��v���Hڠ�ڹ�n�8���]�e��\�Z��ˇV�O�2H運�05l���͖�� ��	��"b�f����4����;^��n����rHbm)���`j�-�՛-��GLX�q�7y���diG1	8��;^��n���{�nO�6�U�@A!�1i }�Sg=s���{�-��Vk4�&&�z-��߸��Wmz˝�@?��W��~D�I	b�F��Z���bY����qܙ/3v�+<T��u����M73�:������^���k����?|����4����LM(�"�h�K~�ꤌ[=l��運�06�˕���&F�����;^��n��c}M_M��= ���&�n6&H	��[w4..٠uvס����|�g����,28��I�l�6��_�ǵ`u�j��}Q�����I� 0�E�(��b�# i1��ĈE`2E�ٰ h%��)%(R Q����-�l
@�[FfЖ�Ҩb`�+,D�� wz��ʰ�j�H���"�Z2�"F	!#��Z |��q'��CC�J"b4L�*�E��#�tR��	�t$mR,Q��tBO�5�/�0R�F�, �Ī�L�1VMEZ@�T�)T�'�`��E��%Ak��Ve/EڤH*o6v�h�B����9�b~�{�ѭkZ��KL0�Q����'[r�XH�v:;r8�T�n���K�rg�p(q�a�7�A�D.�(&
$I+V�smƇ�pg7n%��2Wli6��.��nݸ�jS�5ano����d)V�����六�բ���]�;NY�qr�1'�n�Fj����۲��&�8jV�� R�ԯ+�q[JK[2\�Ɲ�%�G^�l�m[p�9�5��g[�i��QVV���U��s�R�s�m�9�{H�GjF�gm8���@��c1�q&p�w&;X�M��MQ&�#.��їi�9�
��<�u��g�d�y�r�&	-R��t[u��9;���cZ%��Ԗr�1�U��#K��H̡��+΍l�
z�-k�:4�R�RV�cz-��G�E:;vR��x�B��rծ���y���E��y�}�J���x��g����==�ہ��K�O۾~_��8VwF��^��l��9��lp����H��K0�v�c@rl�V���e��n6b^g�ɝ.�u�,3���)�pq������v��I�r�dM���v��k�M9iм�vi�<l�We��3���ϵH��v�y�I�'m��y{]�Η!�����O�$誩C5�h��y����5n�N˭�vv��.c�[��� �UWۚw�]�u-�1��77#���KJ��Qi�9͍7�M�<��z��5U��� f�Ze-���ڨ�P9.ۖU���PcI�g�{q͵�G]W)��m� ۲$Kd���[r[�9��u��%���9�u9�@v��)�i�;�a@��ڲ�aoO>gnvwO���.L"v�s�Y��B�WVX��mb���Ha}d٪�����h�i�t�r��G	5�+*��8H\�t��%a�d��T��UW#'J��~��N���|I����[��T�P�a���`/U6�Z�\���a%ٷL:�e���qU*�NZNsA�7����S�"`^3Z�p�fj�%��?������|����>�t@0^ �B�>=��S�sF\ѫ�e3&��\��Ǉ4�[h��e�7�����sֲZ�"x)7@����6�#^��`�d����J{kۛD0����^{���J�`�X�L�٠�5�t�W�g:ӽ�Wh�F������Mڪ��.�cI��Cu���g��#��N�S=Y͝�[7�yi�
�yu�T�������5���E��mB����j  �w�h�ֆ[���I�LuT���m�Y����Ry�8��l�t�84�]t�V�e6
��o����͖��#�,[8�����Rq�Q�BN=��׿߳?~�;�{s@�⾚Wmzm����q�-_-��GLX�q������1l��*�Vˍ�ORcM73@���z�Z˝�@�s@/mN6G�6)l�I4�ڴ�}����h\]�@��7P2<s8�"#C���c�q��[;���zxz�;Za�d�Mtg�N[��EMŠ|���[w4..٠w�ՠ�n�Q5#c� 7#�9m�{�?A0���(������ܓ��l����!(��V����J)Q��S�r��Oq��r&JK�l�03�nnFےۍ�JI�s�ՠ|���[w4=��1.v�h�cg�8̍._)P���՛-��#����m�}�ߟ�������N
��)^��:��UZ��OC� v�yi|��R���̱�qMMr��v������Ss����u_k�*�y�����M�3@�s���nl�����n��Q�C^��F��i)mG#�-~��>��Zs:�Tɞ׶nI��}��t�=�����<c�7��1s��h����|���.+e 9[��#c� '"�;����]Ͷ�Ș�ؘH��w��W�E�0�ltuv��&�>�;���Z�!wL'�G��tƸ���o��g�"`w/b`f�遙�S�r��6�k�h�hq����� ���@�u���Ҏb�8���d��ߒl�eȘ'���#&)1Šv۹�s�h�ղiW�~@ U�A�*~_f���__-���W�x�)0i�)�w6q�%Ș�ؘH�&�ۇ��2�|���b{V�PX�f���Ώ �����6�rQ��3�桢�E�
��_@���L��L	$uߺ�,�l	��ܮ6ژ'�(�n-�>տٟ�f~H�������@�ڴ���h�����h۹�|���]�@���h-؁a1��P�L���4�"`w/b`l��3T�Ö��ϛq��I4�j�=��������}�|�*T�D-���5�^Ҟ鰻���K2u�{v�t&�t�[�%D�i3��l��^��r�n�Ì�n-t�7vTə�p��]����'����NE�Ю {X"��.� z��	�om[i�Xz�/`�l+8�.�Et����ʭ�GUHgg����GF�h��n�NÀ�N6t�����l�L�֮�1m�k��we˜h�*Z��f�En��ԍ���{��w�����Mg��-�ջ9��� �OOQ����8�f���uv�<���5@' �����n�}������-��	��#�����;[�{
!B���Xkvl�X����U���O�&73@>�l�;]�@���h��h�$I1&�"M���06\��ܽ���GL���	K���&
c�"7��j�=����> �o����Z�ܱ;/�)�!���n�u�`����;�&�uj�"�^y��s�d�����@�s@>�l�;]�@���h�Ev XLdqE�+ ���y�-(��鹰3��lm��~�߱#�/�cLq�͸�B����Ɂܽ��$��Y���ʻ%'�j(��@���h۹�|���=���=�_zbO�Y$�����H�콞���_���ؘ��v{~On;GfK����73@7<�;O����x�붶���n+�~��>��q]��.����`7Ḿ�k�}!��j�-��D��69l�G�Z�[���ߛ1��l{޵`w/b&MS�j��8��O'�Uɰ;��l۵e���DE(Q�ø��r�f�;�T�Jx��D��W96
ww~V�{��nl<�/*�{�<��}|��⣜��qXwg���{ˠd����GL��z�v��JM�����	;�ڗ�B�� �4q�pٞ��s�ZK!!,���W�I?r�L��L�:��Uu)=l	�Jg�'2q��N-�վ��������v�V�"��~�$�@.����Vl�z�)���6����WȞ9�Lnf��~��}���@�W�6ݬsa�P�(��:�/����}��<c�M�H��j�>�c�v�����ԡ(I4�M�X�*�+Tus�^�ʺ����<$�s�<t�t&�:��{���}��|���Q:X��l�~L�:`uf�`l� �!Ó"lL�����h.���ڴ�{^��֗G���b�Rf�}��`c���DyUd�����j���kSI(���Szk�h.�������נw�r�Nd�Q �L��l�:`un�`l�����X �a�z�_��!�T�� �����G��	�n��N��������`C�twa��#vޮ�v�	�����wL;m�*Q��i�#�.7�x�IϷ��ɆU�I]Eխ��.ܽ���!��N�/)���v��.1ui���ݱ��:�9"v�W��	Xh����s]��mX0]�ʻ�@���J�7;����N�5��َ��H��?��{��������~���.�����&�z�L�`;[Y��ۮo
=�s��}�a��c5�_/�o��L��l�"�u)=l���{"x�)0i��˽�}���Z�zm�����ŒF� ��_9l�"`un�g��)�y��z�{�bnbS$���Z��?.;v�����1Շ��*�_�6�{��I���9��n�����/����{^��������zG1$�	�֯E�a��Irj��ۂ�Nz�qƭ�4&�/ђ$��π����;]�@�s��f|�����;��js�lP��Y�'}��އȐ^�B�Z�U1BILB�J�s��X��V��uz�z�\�$�A�5	Šqv���ڳ�y%Y/}V���1�)�eJ�D9���n���k�;]�C��?.>�=��/5�L��Lnf���:�5$��7g�;-�X۵`uO��?�����z�a�]�n����\s�4<��a����^.�:k�?���}?}�[�e���9����6ݬs`cnע�";A��=�?����bnbS$Q�����&�0:�e�6\����5{�,�bN6&9�r-����>]�z,�߇�]'�A�|�+��B	@%#S����	��ԗ`O\�FD8��
ʝ�t���tM���%@�JN�	�Q���$�dp����s�h���M�A HD �e!p�#`�� w��b�"A!AN�-x�}F-KBЛ��hc��eRV+�&Jjf��E��b�M���M�AJ�0A������]�'Μ� O 
�� 8þ������-��-��.��$���Q
{M�X��6Ә��m�VVv�q�G?F�0�ŠZ�Z����v�|���s`yn�t��S?J��a�$��ή�S�]�qsuXॲbw6���Q�c�[��y.>���I݆?{o������m�V�X��
<�h=����~��xq��9��m���}�@�ڴ�{^�qsj�y��4���s`7M͞�S=�����V��,�ț����h�V���k�nՇ��DT�1́�u���UqL�$Q��Z˽�@����ՠZ�������.��2Ra���
qK�P٬�\2v�Չ�1���:Q�t�K�D�0NG�[n��_j�-v���נ_֗G�̒b�Rf��_j�$��v[I02�`:�._>�ع\J��\���6[I07/b�;ǋ�q)�88��C߿~\~�z��nh��Z�ՠs�bN��D��ӏ@����}�@�ڴ���ܓ�!BN�C�&O9�s3Yr�]n�A�������]�gt<��	�d^�'b˞�E����Y�C��Uݵ�k(h����1gt=�Qle�k�\N���E�)��v��vs���8p�B;fշ�����i�L�94�I�=�mٷ0aɥ䗫t��I9N��fEn�8�|�GŎ���^+J]�e�BK�q�^�{GH2�7[N���ҭ�fיnJ�)����_����N������i^���#g]z�*GPt3���'F]�MV;�s���3�eOG
\:b��wʀd�~L	.D��-�$��{ۋ"ț���JH�]�@�^נ[n��>ՠ\��qɍ��L��(��>W��۹�w��h�V��iY��lLs�z��h��Z�ՠ}_j�.v��1�	�Dqqs��՛-�%Ș��0$���o����)��*��\S�y�VNݝ]bFhq}d���e�1�Q���b�2�3�W|��"`v^���GL�ؘ��ܸ��8�f	Š}_j���g��AS��U)FV��n{g�4y��@�ڴv�I�7�C���-�s@�j�-v���V�qsj�dOR`�s4.+�H�ՠus��������Œq��iI�k�hWڴm��:�����~��������W���vylv2������p�V�٣�d��:qn��.��V��	Z����������/�{��ZW�/I�8�jbnE�[n���נZ�Z����${�H��"`��qOO8���,鹲�%i(" ���� �pX�T���;��;o�4gmm�Ē�b����-v��ՠ[n懳徚��sؔ�c) �@���h�}�}� r�M�ڴ���Jd�d�1zK
�]�$^]�ۨ�&��;��M��^_a�t���N
I�&�"��;m��>]�7>^Iv�6��`j�'��&�M*�Lnf���k�~����Z+�Zm����������I��zk�l��͚��{�j�췵`4�Uɍ��O�B(����عe��=�{s@�������T"�R	@���1���g䔵h��TS#��6�SU�M��v�����v�f��+��������c`�� c���ۤ]t�Dd��W@5�#��OB'����5���I1B)3�8���-v��ՠ[n�̶���I?�1L��-v����
�ͭ����j��s^��2<�-j�$XǑ�`�Z+�Z��h���ՠrى:(�h� n-B���ߕ�u���76����ٰ=����E	�R`�s4����mܓ����I�{�7$ڵ�E��wv�������;�b�\�xh�Ħ�/�:<�p]�uT x�i9��SU����j�׈����a�WL��7i�@Rd����s�x���>�j�LrseDt���>��9ڞ^8[��y��k�ʻZf��v�}�nv�7He��c�nD�n.��7	t�suR�+�s+p�.V6@n�iqA\2-������$[���s��zk�V ��_�=�﯃��5���A�̱cSs��v��i�;<������6c��A�/:�����}��K��⵹��?�����ؘH�wvq�*o'�֋��5�SZ�]f���w���(���j�3wܰ���Dɛ[��q��ژ��h����w�h��hu����ˤȘ�RDE���ߢ&z���{Of��+�y$��$�}��h?���oq����q���hm�L�0:�e�?-��h�t�!V8Q�>�����[A�:��۶��9'p�;=�%�(���~z�nn(�xǑ��p���lx�XNc�Dz]��V�l�q���M�DŠv��i���p����+���e�L��O�URD����$ǎ)0i���zk�Z�}�@������PY9i�ܜ����f�맳`c�j�R�3�����d�ۘ�!#$�hu�����~_ u�偎�̀�|�|�Sss�w%av���=v6^'t�9�n7Vm�r�����5���l٢�$q���bnE��Θd���{m�LȠ��IX�R
93@�v��~ċ�|�W|�����~H�{�i�Ē�b�ґi'�g�]�=���"�����f~�����h��ܸ���GE��^��h�ۚ�h~W��h�`���#�Šv��hP�s���i��u�l��T���k>�I�Ӎvp7+hW�4"pu�BC�~���mm����8��{�羍������-߽�)���6^���{f�L$��x�yM27���V����g���?+}��`9�u{
!H�(�BQ"��W�n~ɫ�3F�����Z�؃� � � � �����A�lll}�߸lA�l��߳b �`�`�`������A�A�A�A����u�Z�fe�sY33Z�yB�߽���A����u��؃� � � � ���~�y
���bb�N���C�w�w��A�lll~���̺-�n]jkR�5�b �`�`�`������A�A�A�C� '�����~���������A�lll}�߸lA�lll~�g&���qZ��n8���	;�)��K�ᵏ�m��u��̸n�>g!G���~�x~׿]�<����k߮�A���߽����A�A�A�A�u��؃� � � � ��/���kXd�Y�$�j�A�lll{�^�v �#� ��A�A������A�������v �666>��~�yO�9��~�.K��rk5K����A�A�A�A����yg~͈<����6=��~�y�׿]�<�����M~�3?����2�h؃� � ؿ�
E ������y����v �666=��~�y~��y�߿L���j�5��r]f��A���ߵ��b �`�`�`������A�A�A�A��~��A�A�A�A�u��؃� � � � ��09Sj@�I!02�D�`�O����^ ���Eh-$(.` ִ�M
�?���L�CM E� %7���>W�PH?ҪD1F��O��@��P)�ϟ�(h@�%6Ŏ"@��H p�X����B���J�kn�1h�1��0�I 
�yM�I�	��	��
}�ن��(&0$1% !�"�)��@�!�ȡ�P����!�Yi��{���t����p�I��˛.�-�FQ[%�ʭ�)�I��jV��������Պ�e���S���:\�9ˣ�v.W4��KTnT��r]����`�����C���ڶ�Z�&(�ԪX5;9�v��MUH$�`څ����]K���R.#��B9���;�umv����H\��{/CL9jU��-�djq4�eRZ�"�eتL=g�D.j�$ ��4�۵�Y��6)6.j��QƄGK��On�n{kK!�N��r�2���@��¶jS�ٛ�z��Fo���ur��l�dz.�s��D�Nޑ嵳f̓i�؝��z���F`6�F�'C�#L����E U�8�`���A�N����3�qKϠ�؊���*���XÑm��<`�,+m*�K�����]�!g;���'s�J:}��I��ڡF�ɹ,�����L���.�w-��K:�Ya읳�Pgl�*�L�p��ێ��r�V�4}��yVAs��Kն��bI�J4�.�^Wnz.���>��mu��n�9�i�fh[ մF��5����1/c�w M�3�n�P�6�Mm�l[a���Nݚ��N�f4�˟\��OMixv��qnN�h�7<I��qK(��J����.R�Ǌwh4�M�+��;��$p9��^�%m��n�dvd;vNA��lAv��'o[�d4.m��ې�v�ڶny$��]x6n��H ����vƵg��5U�@���zU�fq���[���gM���f�+���ت�ܽ2�]p��Ƶ�
\���氘9�9\�Oe��`2D��;j\�t�Kё�fՓ�s#�z�I�mV۝d����>{L�,�K
ezn��b��+ �UV��@hg� |�e����q���6�"^��:1�m;���6���Cm�������=��T�N�T藋v�y`�)���6��V�z�K���VG��9�&&d��\���Qu�h���q�4eUƩ�l=q�xiΖ瘇��u��w�߾�C@�q^
pE�%z� �&� �l�_8ɢ�7�d�:ڝ͠ƕ����j��>�γ���m� M�d6y���gW��A�ø�K�k��5��S��9��Y���u� `0���sg�e%�s�ӡ%��){8�����s�
��-.��܀ę��wXw1ԥ�R�ی.�6��;����8��0�\���,�v�����p��u	ԓ+ZC�r��v1�-�^�h�Ӊ�K��{}��EX�Xm!�d9k�x�ՁtiG��խҚ����!:?��{���w7�Zə�Z�\�u�kk�D�lllw_�]�<�����{��<������߮�A���ߵ��b �`�`�`������F���,˚�s5���A�A�A�A�~��A�A�A�A�u��؃� � � � �����A�lll{�^�v ���D� �l{��N]jK�ܺ���Z6 �666?�����A�A�A�A��{�؃� � � � �����A�lll}�߸lA�lllz~��&g	2�u���u���A�A�U[�׿]�<����k߮�A��������A��,}�~�v �666=���u��0�j�3Z�y�׿]�<��������<��Uw�z|���：M��`�B �:�f�Ƿ��N�6��v�������U��{ٙ�wpLB܂#�qp_����v��������u;�dO��.f��;�{�|>� ?
�{Wٰ;��lx�_����յ�W9�#��i�8��|��ڴ����W�ۚ���\��d��S#1��I���Q:��l�mX���y){ǳ`u��Ȥi��ۑh������/��w�@�}�@�ut�7�I,��e���ٖ����[u�x�q;n�'=J�`����$BbmHI�93@�v�����c�(P���o�X}>
�SQ<�yV�8�/b`d����c��ȟ�/Z.{qA�#�"�;�|���f�<�@&�Id�p�(�*S�D<sy����=�>��&��k�G+����a�Q�[��S��~L��02^���[J*��D�nf��;V���V���V��۹�q]vdQ�� �LM��D)�z�uWn�3[$�FK����y�T�����X�|L��02^��ٱ�r�Z��VI�d�nb�E�r�ՠc�j���s`c�s~P�)����r���cnE�__nh�i�ٙ�+�|���-�����Rb�E`gi��1�9�:��j_$BT��� pC5�����o�ܓ����4�(�1�"�;_j�9_j�:�ڰ3���Q��[�Tʕ?r�5ɣ�Cl�nƢ*��v���8(a1;�V�=�c���Ț77�A#�"��~�Zf�L	�"`l�����P��Â��ɒ��`c�j��!L���6�{6��Zqu;��<Q9���^;Se�L�Iz\�`OO:`�Z9tp"y$M1G���V�z�V��۹����yh�Xy�y1����h+��ڰi��1�9�*#�	?�*�O �@
���ȧ�f�)�v���wj�l�re�ն�v�M�`\h�uoۭ*M72����e��a�t5�SD��wm۸�]�z�6-�5qh;�R��C�/=$�ׄ���Wн�͟.���]�ź�rѶ�l�H���,��.�ya�s�`���n��c<��w3��Nx�񍠣b�� tLA�(8v�Ԗ��$KOT�n4��{����������B����֮���C�R�ڵ<�=�+;�]���a�oH��G��Lq�����ۚ�76:�>^P�h=���wg��9$Դ�$���^;V�~��H�w�@�w�@�����ٙ������1cO�SS��=sɁ6�&g�%�r�ˑ013��bƚ��331^�ՠv�nh�ՠv�ՠ}��L��,jBNW&�ǎՁ��"�7g��ٰ>ՠ�~nc�!�q�!,m&����R;\pƹt6M���-�瞧S���ف�Uq|�ń��̀���%����8���������l�&���@�X�څĒIU��lmڰi��f~���������	��nb�E�w�<�6:`n\����&e�.�H��bnE�����د����~��;_j�/_j�;�ך�BbmHI�W8��nlJI=���t�lyw4��FВ,1�Y&'�n90۱���\<��si�������N#�C5�&��|r�⩞rlu�l��lx�lB�>A��y��=�H�����h+ߡL�^ڰ6sv�u�oT(I/(Q	U��W�.�k���������z��f���pD���W]��;�ڴ��V��<Q9���Т�Y�V�{6��6Q��٠�{�Ɍ#d���zk�Z�%�{? �vՀ����s�#B�<����<BN�r������e��킵�����뙍�]4s�vN��/�O��X��ηj�s�u��G���l��IɑE6�r-��s�g�.�=�=����ꄢ"<���wޥ|��6�$���+��v�ՠ^>ՠv��h��Q��i�Q�c�Cٙ�^�����lx�Xb��DBW��U7��ܻ�}�Y��kZ��a�ԁ\����l�����|�=��Z�[�L�6,0����Loq���	��/��X��:����ᱻ^�n��l�����06lt��{e�^����u�-����	�N`��h��lu�l��6<v��BI/B������2c�$CiI�����^>���B�2��r�́��Z�5̐��)$Z��3��e��/��4�ڴ?���W��h���92(��bnI�1�`j���G�易o�}6�w�rO��Db��H�T�$G��ܝ���n�r��x �&�5�G�9�8�#i��e&������u��6�kp9�;7���E�綊xGڂڵ�n��Q��5�uF�vY6y���M��au䫂;a�Iq�-5�/�v� ���ͦ�4U�ۏ���#��sӺ��n�{sJǣg:��#��W%���xs(m뭷*s��3���qn�uPYԛmkK���h�E.��w}����c=���)�a 7H�[�ɷcJ]���c����u�Њdn�PM�	1G&tW���6�c�BP��z�Ձ�el�ʕSQ<��*��M�����BP�L���l�o4�ڷ�?~��"�����8�s������#��ؘ.D�ܰ]
�y�!���w4�ڴ�j����߱{��h\�~B�#�+�0&^���r&�ؘ6:{o���]�{��˧<y4s��gi5F��4睍n��>�~�Э�l��_�{�������՛#��jH������x�V��۹���?|��w�@��,=��Rdf71I"О�;�> �	@D��i(�J���V]=�c��(Q(�ɑE6�r-��s@�x��D(�/i����l���	�!&(�������������L�����=����oYI��e�US\��X����=���ݵ`>�j�޺ё�B��͉)�'���-n�k u��1nö�.�8��m��j��w{��~M�}�I!�q �_��}�w4�ڴu���x.�a8'Š}�ڿz��UG�o��{[�>u�l��n�L�d�sә�w��h����1a�\��<�Ha>�����V8J�ˁJPq`A%&�sI�qLD�D>�M����@tqA�R$0�Z�ـ�F�N�إb�tmSs@ "b�(De�p@�D��Ɗ�	!�Wut�(,x�l# F	�P{��:���D �)��A< 
|�|�|ky��ɹ';n�s;ړ&2cDsmI��ffyBP����M���x�3�ڰ3��l\3��(�Dcs�-��M���ޅ�f��]]o���V9�3�&�%`�/Bl�Hu9ݛdy4�A���畸�Z�i���Ɍ�JZ���� վ�~��Vv�́ܬs�%�u�K���n�mIĤ��w��h��Z�8��n��(Q2f쭒�R��9D�+�`l�����A�ݑ�r�&8�r�rE�y@9��g�˞��B}�߶nI߳�����B �#P��8�����۹'{����WSS5.r�+����遹{6�&f�m���?��p��AŞ�Y����`�V�3m;�]��G	�;s{4�F�4�JIMf�����nMY�	�Ng@����-�}�@�즁�m��e�I��dq�$Z:�f�(S&��^�����JdƆ�1#���h�x�>�f~Ľ��-��-��SrdC�$)��8Xy(I%={�+r�f��V9����w�|h��1���&��I3@�)��<�Dc�����,��V�J;���[���K�\�l��#��>	C���"b����آ�.\G(Yypu���}�n�c�d��Qڰ�99�mb�.z�쫗l�	�t��O:�����mщ귫K;v7@�]�d���ѝ�u��k��]�h��4on�8m�Ս�WJ�]v^���6sv.+]R˭2x;	���]U'u�!)ugQ�vCmayVZc�Z�C8��{�w�{�޾��j�;��A��]�(U��%�td^X��9j�M������?|w���ûH\�-=~���"`wdt�̹2�r�qŀ�2`9��;V��m��;�nl�c��Q�$���D�\��� ��`o�~t�̜�?%��u��@��V�$�S#�&����߱w|�06\�`f\��ݑ� ͭ������&�R:�V����?g{=������YM�*�,m�ӄ��frt���S�\�]�;<V�B���'B�]��1#���h�hv�����ٟ���;]��9�s�Ǒ4����Y�]�9�{f�Y P�����k�-��-�v����J$�$jbRL�9�j�9�ڴ�fg�ؗz��r�ۚmYQ��0�S����V9�;�nl��V�Nfޚz���7X#&�h�hQ׻����r�́���j�T��H�ΩY۵��%�h��c���k:�ϛV�`��Z	�)�@&H�� n-�۪��_`w+��Q�eǹ��U�JD�FG�s4qڴu���v��۹���3�䃷/�d� �M2y\�=����Ϣ8D"!UV7j���ՠs�w�Čnb�E��ġNg7f��ݵ`w���y$���ٰ9�sɩN4��iG"�>��g{=����h�h����U=#q���n�K��넚�*�n��ϝɣ��d���њr3������\�R\w�bK��03ob`f\��ݑ�dU�X/�#Ɣ�@�_j�g��������vՁ��s~I$�L��.M��+�OW96eń�n՞�
&s+vl��-�x.�$Py�D��;�mX�76]c��L$�	BBP1"�P`#�o���>Ig���δ��H��� �Nf��;U��f���NnՁ�nՁ�C�[���Ӱ�H6��c��������N��%�x�T�WA����q1��?����;=n��v�Dy(�u�M����+bLs1��I���^��[��s�ՠr�ռ������~x6��<o�M��03/Nݼ����-��l�$�D��1)&h�h��h\��廚mYQ��<�SR-%�LY%�7$t�̜��UUU���t]J��a�X�LO��z[S�j+Į��dլng���\T��n��Fp�Q��[��+tF�q��5�=ن8э=���z�$k�m�ۮM��Ռ$��Y-��v-q���ݕ�<��6ܑ�Ո,B�Zy0�n-�ݦ-�g��i�j�
�E��\j�������g9��win���e˦�1��բ㐌��7���w��뮿YC�;~����ۢ�:3#��Vc-�Bs�V�=�c��ӌJ"1̍!����\���rGL��02^��ݺ�S�\\�W�`nH遙9Kؘ�G�H����jD�F9�s4��Ɓ�X��$�(���ڰnڰ�n�W?L��F6��h{3����8��=��s@�j�9p�6$�1#�I"`ud����遙��6�&����%&�;��C� �9���k����⳸��I!�QN�TWB��82�f��#�f��ؘˑ05M�-�l�rh�h��hܓﻯM��/���}U��<��`l���ٱ�dU)>%���4�6�4�ڴ��Z%}}��w�ۚx�P�9��8Ҙ
E���B��7f�{�j��qڰ1�s`gi�e�H�8�8��w4s�s@�r&r�LMۗ�_Z���(����+je{F˵ӷ��.��p�j����T��E"S#�bs>����;]�@��ՠv۹��r��d�$ci��`l��$f߼���e�L�\��5��l� ��hqڴ�w6bD?��Xb�a�&!3?M]~��>��Z��*nL�H��.s�L�:`f\����Lˑ0;��ĚH��&(���v���{ˠn߼�$t�0�P�BH�*��]X��n0۱��5�xm�c:�c��5�P&`:;NI<R%���4�6�Zk�h�h��h�h�]I\�mbpJP_8���06H�ܹeȟ��ٙ��-x+�z�x��	"�/��r�L����Ɂ�g���TS�K�I�c�LNf���@�v����C�pA��%CA�f�nI>�hǓ&�H�ӎ-�ڴ.v�����;V���.��Oc:��R�˷;^��G&Ol��h�����!Y����!�L���E�qs����hqڽ��|����@�<�p�Hc�w��6H�ܹeȘ�e�}��*��Hi�1Bb�rf�οyh.D�̽���GL�����}uʙ⪞rl<�D(R���`fSٰ1�kC���߱s��Z�T��A���)��L�ؘ$t��\����LL��`�(�/�"B	��LSB'�D�&0惋�2���&.lֳM�fC�@bD"�ā�0�6����1�\U;��:���4��$T#	�� ��	=�d,A��Ԉ% � T� :�RJ��sBTL]kE�Nxܬ�	��H<R����v��߼�h�fM��de�7!KU����ƜuR��r2��[;�;3������S-�ᝳy�Y^��KTVll;��qcc& A��M�b�W�j�cH��G�3�\��^��T���"0q�%D��r��E�f�%q��VQ5�h3t�*i��zk�ymZl�E���� ��=B�WAU� ΂�ȴ�WG!v��oEN�^����I�U��C�zŇf�Ņ{���Y���g�� [f�A49�6G�Iw$Ny�\M͛�j4��<�Q'^Jz���N�aH���F���i8����n�R�]�q��=qC�#L��cI�	�`��b�\9qͳdyA *
��*����"��AŢ��E�-��Ɍq��b��]�7Y	ʵRZ�,��)!��ۑv����L�ٸ���z����y��q۠��lnC�^{[W���@�cm6�l򫩮�B�'�� *�6CE�n�� c�܄����⬭ΗE<���\*�v���#�(v��@f�c��ʣ��i�l<�+�ڴ�x���1�Pr�O4c�dj��B�rvpUF�I���V�>�i���5��n�]�E��2�";���g8��x�+c�P%S��\����[���:Gn�F/["Gm� �Y�[gU՗c������e̼Զ�=�:C�FBʑ�����F��7JZ +\��l�-U:�X�fÞ��%��ĵmV\l둵*��;e*�s����n0cV�x�w-Ӻ�U(r:ʺ퇎����������9` s'I��g���b�*���^c�z<�_
�V���R�[��2s�d����>M���Br�
d]��c-��79�+	\�VՒ7V�r���sT�2��8�Z��F#����lq��%�l�Z� 9��tQeR�
8���;c��ƢV�zJtGj	��.�u;��������м�Bw��t�s$�ao��E�KY�.=��se,�m��8���y)<�U�ʝi{�w����{�g�Dn���x MT����Qz	��@)Pt|���D���=Q�Ov}܆|d�Y����]n*�����\�mET,1u��΍�O��)��+�5��y��rX�q�-�/mE�v{Eێ�^Mv��7ll��:����-���n�v��u�Ths�J�Kq�v����cy�'��$��x�#�&��z��m�f��v
"!]UA�n-�/=R>0V�	]���1�N�ll%Sӄ�5ݨk�S��f�W��ww_|�'��q۶y��;VSf��j���X�����/��"简�������`I ����;V���_В�D%��}6�ϧ���93K�s���_)�ܹeȘ��06H������3��,���F&��h��Ze�L�:`w.D��D�I�ҵ�$�C�?.�{�@���4qڴ?�33�+��-�w<�y1HĆH9$L�:`w.D��r&e�L_��?�*qv��$��1^Nݶ:�w@�s�=] �4�v��'����u}��d�sh�˗�W@Ϳy06\���{��0�j�.	�\��)��&��Mͥ��Qi/��K���O�`7�Ձ�i����߿f$^�R^��'��h�L�0;�"`l���6�-���B�0#�@����>�h��h{3��ػ�|�
���'��D����r&�ؘ��06lt��U[�v��NO'hu�l���lc��^x	��~�}�}����nzq_�w�����x�{I�Ew|��������{f�L�Ș�w.-�&���H�q���c�r�L��?U}�$d����H9$Z�����M�����d#�ˊ���# H`D�F s�Ϲw$���]�;}�jٔjc�D���4?ع��-��-�}sa��G�%[��U��<yM�.T�|���03.D�ٱ�2r��������4h��ڭU��v�Qƴ�؃.�%&�r\�u�H�][�����VS��<A\��eń���|g��]��=^%Q�F�J7 E�v��n37�Xi���c��˝�U��&FIM9�;��@�_j��?g�K�w�@���4��(�$bm��X���k�cv�(J2Ev�f}w�x�/���li50b�9��{�#�rr�ؘkk��v;c�t�>�]��� sg��l'��t���]�3�'C�b�6uf��mݑ�3c�m�^�ﺃ6����{�1<��&7$���������#��M�ܭٰ>��^�J/%F�����0_�F�rf�|�����Zݷs@�;w4q����iL"�������{����Ն�QOo}6�ļ��Q�ҍ�qhv���?~��ǿ/��Of�}�2��hP��)J"B �{߭����R]MK�ն˄#��`�q�X���KX�'m�sͩ��4(- �zu��ы�X�S��0�&�g�/j*�N9up��ؚ�]�C�%�9����흰`��t�l�ƨ*��+�&�jŞ�s��v׻BG�F����sԩ����c3Q˚.^%njK ��X���U��Ѯp�<.�Y����p�8t�H�u�p�4u>z{�xÁ�[WP�x`���?}׭�:ۈ6�M����uӪ�[o��mX��6�q��
>��ݵ`[���xA�bm�3@�_j�>��Zݷs@����;�r���j`��ds��ܽ��ݑ�=_%�<遲�:��4���c�'$�@���hs�s@�_j��~����U���<��&I$��v�h�޲�|:yn��������a$~�	x�����3)�-���qhL��g�D�T�:�(���E.T�T���5�ٰ>�c��v����s�ۚ��G�!C�)��Zݬsv�yv!/�"2(��onՀ��j��}�@�x�QqF�B�0#�@������?}�%�sɁ�sɁ�TR���&FI����v�h��hq����� �^���H�I��V9�6s�g�77mXw��g��Oe���ܔ=\���2k��ʏ�.��z�盦S��<R	vt���r�&�0;�0&���ͽ�6���c�'$�@��s�cgo��4�?-�>ՠw�<L1�(�Mf�nIϻ훒{��]͚z`$A�A�ū�O�� ��|��s�߶nI�v��瑩�5&h~^��h�Z廚����>V��H6��J`.q0;��0&H����6�&�����/�Ũ����:�vq	�S�4��lb�θ3�շX,k�Ch�n�ɉ��/��2GL��L	��0;��05v�qLq##�����v�m�ceWg�w)��fqs�B�2OIH�Y"�m'3@���hq������v�h�ܨؒj`��dr-g���脕c���~����`�!	.��V�B�B� ���.�Z;Sm�JL���c�E�[�����%�L��L�}YqC�8÷������zs��b�����<�����gqi5ΝX7C?���݆�xv�`]]5��6{���0;��0$�遳U�!bF�4ԙ�Z�V��j�-���>�n��?~���Uy�1F���(/�L۞L	6:`w6:`I{��]E��%�G�on��:�X�9��J�8�l/jvN*䔣#�����v�h�ՠ}�ڴ�w4,�\J�ȅ<mE�)���(�hzӻ �H1��^p�͗D��מq���� �c�<��u�燭����o����K�r��=�ڮA�\N+�uGl����70b0v��#݁U�2Ñ�7mn0I�5�������1c���u�������q��f�lМ� Mݸ�#�{a�R���+ρ�v�uu���f+��8��q��������?"��\{;,��P�of5��!;<U�\:�=�o8��Hb�F�Y�!76����s`}��6�v�?(��c�Z�=���lI50dj29��j�/-��>�n�z�V��:���%&LX�c�I�[�`}�v��(K�!U{k}6:���kX�c�!�L�I�����&����^���#��PI�T��T�T���yX���J;�{?��j�����2��,X�x�qȚ�zϛ�'�������%8�ק&�������_,��{d��͎�o�h��.F܉)1�G��{w5(�bˠ��
A"��H"A��P8��������[�`}��7�
dr�և9%(��nf���nhu��=���:�}���W0��M19����U,��L۞L��L��L�j��5�"5�@���hw�q�I/���}�Iq>��$�l�u r$*���;Ή0Mg`��n�M����gq��5�JM�ﻻ����r������� �έ���l�w�%��+i$��ػԒZ�R����cNLz�K�v��|�\W�[I%���ޤ�-������Ҟ��]��F<�Li�3�K��'�$���_|����iP I]��:Z�IZR.:04�X@�F5cA!�q��Z�b.0�H�$ 8�?�~V��'"�U�9����a�o�s� �����"��JFa
[HX�$*p~bF �0n�
l�����X�6i���� ۡSm��_����VT��aB[k2��"�$����#^K�������u�OA��H�7�e"�h�uT�T��e2 i�D�
�#)�P��B�A2C� ���G�
��/�`���B��B |f@�aB�I�Ϙ��RP#V5 5�aF3[��f�5�KpM�b<o�Q ��0j�G��f�����)��?}�'��G� ��#�\7�^��
�":v<ESO�b��������ٛ���}~ϾI.v*��b��pQ��ORI}ɱw�%�c�i$��;]�K�}���y[I%��J��r$��_|�\]��RIw6v�Ԓ�{��]�l]�I~�����?����o�b�#˖�^�횔���	v�Vü�ܲZgj�͕:9m�`zt����o}���9m�\�n�o>�}�_�^�$����ԒJ�{����A�&����$�^�m$�s�z�X�:��K�����%ņv��6�mFG"z�K�N�ޤ�-���ꪻ����z�Z�y[I%�{g��-5�E35�5���-�ʠ�s߸f���~��[o�;뛶��� f��o�$���K��E1'&=I%�6v�Ԓ�ߪ���+Ē[9�˽I,[[ ��q������M��X���3���g<�v�m����<�Gb`�V0nzW*ծr�Ԓ�{��]�l]�Ib���I/���}�Is�U���7��F�=I%��������j�um$�l�k�I,W�=I%y1.��mȒ�i�}�Iqv�[I%3gk�_����U�+i$����RH]��L�##�M��R_߿7��s>�$�\�Jf�w�%�c�i$�vK�]���_���?��������s���m��홻m�����[l��
�`�(S G���5�`Ma�a�.��m�����{(�;nW�&� l,& v��\/'Yے��J�������7�gE��a�U�Ю.*tt=:�<�r�d=0v�<�m�j��4����7iV�h�	sb7<r�m�k���ju�7�y���'��A���`;<]s�cW/W[+O� {jí]n�5�g�7a����ԖMѻVzc<s#.kR�d�Cb��[�#��Y�RL�SOl��R�C������g�{Y�f����y��s�iL2@����Q�ȟ�$�����űմ�S6v��}�i-W=l�r�J�Id�1cq�ㆁ��@����8�����h��K��E1'#�&lt�ś-���/l�-�����!#F�4ԙ�����|�v�˖��s@�z������⍠S�`>�`z#�����mX�� ���?�b��{n{Im��M�u��\�s��z-)���ᱵ�W��8]+@W240:�K`L�運6[f�v��L�##�M�����_�?c����P�j���ڰ7w�XO[� �b"&E�$Q��h\�z�e4�-z�n�ņv�a#s6�#�*���+�~�`d�z��v��qց�Y��b�&,�3p�>\��6:`b͖����t�Q+��Ü3ؓT`H(�ӻls;�ш�^�W@�ٜ�nӸ�1�~��Ԛ�7�9"$�9�{��LY��7��_}��޶�/	>L��*x�jy�`v{��TB�	L���X�ݫ���(Jd��f꧋�T��<���r���,��ՍDz9*,J3u������@�x�Qr6�J9�E|����-�3c�,�l	��0�Wp�"&F'0M�������g�ݬ{_��������=	D%{3hUG?�`ӓ��]EnC	r6ͬrH/l�������6K��8��ƍts�\��~�ߊ{��&o ���-�3c�*+e���ڌ�G�}�ڷ��3?$qw�z;}��qs���q9�G2c��|�`ud���lt�ś-�ܽ���mȪ����ÜD�9V��%�}չ'��f��;�>Ұ �P�¤D5�潭�:{��f�-��ʵk��,�l�f�yt7������-zO�l��G�l�k^�����)6��=s��A�������||�Ҽ�Q�
G��Z�-�����9�ڴǉu��c�n- ������2�&r�&�R��q�Q��U\��qڰ;��6y$�^P�~o���ho���^�""dX�E1�w|�e�L��L�'͎����,n`��b�-�>ՠf~P��ޮ��}j��k����!ilj@�T�0����/�֦���R<]g�y�:�9^؊���m�+�)��B�r�����l��3� �[.r\z��7�u�\�jQ%n�,җ<��c�v�Z�k�9:����[���CZ{a�I(�@�Lx�'[!ٹ�Wa�7+K�
NKm���z.����mР�9�q5�4�s�9�z�+Nv�v�N���4����n�����iVtZ��K�;�h�b.�z���8p��ꔲ]kW&YrEպ�Mų�����;�Fw�Wm9t�\��K7\6ɏ#�qȾ�����;w4q����:k�K��DI�9&�����*���7ny03ny0:�K`w/UC�`�<�1����}�@���h.Z��۹�s��jjdm�qFЗ8��ؘY%�;�0���-�O-��/2A�F���R-��^��lt�̽��ܽ���6+J����*��`�N6Q�7%��(�"	��S��n���FcX�y#��$D���n?��o�4e�L��_���[�[ �OX�#��O$Q���h��[��~����C���y�s�s@��;B�F��F)"`w/b`ud���%�<遻sɁ�%�̘�8��C�331q��z;}��s��hq���}*Ȱc�$9����lt�36q�ܽ��Ւ^������z)��&H�ŐM���<Ps3�Q{F�8�
,�蜯W����������~y��Rg -���>��Z˖���9�2���C�hq���@�s��5��`w$t�36q����/_+�9�c�H������;w4�~��셐�/�'>|�:��bt���I��򋻾q���運6[�{�_~��}���@/������#Q���hY���7�ˠ��͎�J�ܾc�/;2�#�����x[�6z�5�Q���/^���:�&S�õbhI:i�mܽ��Ւ[���l�d�|�#�1�q�9����bG;}��uv��q���Ď�O,�9BL��l�,�l��L�'P���3�ƚ�4?�~����s���I������b�0R!�P�-�7��}ݢ��'�%r�v�s���^��;�q���運6^��ah�KcC��5���%�N@��<�0�#n���pgͪNH�,�I$�s,�5kY�B� �I�sc�,�����۞Zny�	�"dbsۓ@����,�l��L�'MR��r���E�3@��k�/j�ٙ�9�zh����gn9H�FG#�.^��;�q�3c�,�l��
�F)2b��r- ����s@��nnIﳾ��@cn���F3�,HbO�-����
�P�*M1-�N�!	!4��`�l����$�" m��	0҅���#1��D�=��8!�%��tz�4$'���u�C^�l݁�LZf�"I�ӝ�ﻺ{﫻ߛ����x.�g7Q5��, �.d	VwTFq(��ry�0��x�Q�#��]�,^��޺�7d��ۮUX?�~>�]wf'�;'��e���Ӈ����L���n������ʱ�e�V����]�%%3M�6�j-�(r�.�J�@P>Y�L��٢uɍGa^��g�r�1EupmPNݨ��*5�&J�[!����u���xy�J��1�V˳��5RN�TMs�3㭢�su���1�������U�'5��9��E�*����uu�W.磧N�9&�0�VV�)�uX��]Mlr%����35��cls�^�0�%_VՂ�gbYY"@�/"m�7M��f�Q���sa�M��UWl\{���`p�����6� ��u�����X%\���:)�w:Rx�I�Ό[���G9+�I��/nڷQ���u�vM	lN�tFL�S���&���I�}q����[�H.UV�N��s�W#�p�8n	덮\�fڋ�W���N����*�8���z;�6��m�Is������ؙY���嶵�l,r�@s��Õ��- @���굕���ם��6���|�>N ~�NS��v�M�r�鵰��w��C�����<xʇm�q:]�-�n�7[�����zIɪ5�;%����ggeE�6����n͸�Cl�k�O��a�-X.;d��Z�Y<2�h� l9j���n�6�;�Z�CbZ��>���VѸ�[l�4���ջ^��vݳ� �X��t�ۛj���Pz� 0d���Ae6tҗX�N�ti���UD�xyw)ҩ�ѵ�n�@��X�烵�#���uvs6�PJ�`�[D�%ݸU�[��tJ�;nV��C��YGr��r#Z�۷=.ä�R[�� ��Hڦ��҆7�lm:{-�m��P�7OJ��%r��V�T9g�jě�y��ۭl� ���P��6�It�Z{<��z�i
S2s�!�sU�g�uW{���}A����Aӊ�
��'@à����*�@N��<u<R��ְ�FkS53YgX���E��^�0�kn,ɧ�;O�e�P�=���h�5��e�M�^W�;c�e9�m�C3�n��[s�givsi�m�^�|Q̽�V����Uȶ��d:;i[u�q��r�f%ܚ��X�n�t�v��ɹ����W��٘nV3¬L��u�:L7(Tj������$�l�7u�E�֏����k�7\kO3�S����|}��a��]>n�Ӹ5>H���9�)�H;)��qi�uٲE����wtV���涡&$�o��4.v���� ����N׭�I�Q��8�h\�{���2nSٰ��,�v�RIy(Q
�{��n728�㍠R=��- ���<�!D���VN=���$�.ʩ�qR'�� ����}�j���Xz%�{��h秂d�y�����/;0͜`L���w$� �շ9k�Ǘ��l#�S��&�ٍn��\���X�ï3��s�/
C5��Q9�n�m�����	��0�`L�遈�"�._8����5sZ���;����<��";��/ܰ=�֬����!%2ww�
@D�1cq�9�s��@������4�ڴW��E��!&$���$�DW����1�`>�9���h�[�<x���Sq����4��0��0&lt�+*KV%J�Y�K�鋵Q��yʱ'^�F@�\��Z���S�t��D�cs$�q��I4�ڴ�����֨Q	/���X��N�\Pq��
E�s�o�f~H����v�hWڴܲ���28�ۓBw��f䓟w���?DG�;�S�	DJxU�_���rIϽ�[�O�%�9'%R�'�RT���B��{�X���0��076:`b4��K��$,�G�hWڴ����.v�|���}�٠^��Dq�I' �cn\�S���n��V�L{�;��9m�ݗO9k���w�Ѹ�8LX�d�E�;}4�s@>�l�>��h�;L 1�bO��sc�����6{���&����[�<x<a��f�}�٠}^9��"&N��Xڰ;�Z�U�UʑGX��C��ff.z_-��=���ܔ��®ﻯkrO��Y|a�Yu�긨'���qՁ�������X7ڴ��1��HF���1����F�Z��ț����r��Y{^m)��Q��<E]�-���� ���e�LY��;�q"xE#Hi���l����RFz�-����O��D�J�%	dj8ܓ@���:�������3����z�hWK�@C�ō�H���՛-���� ���e�L�2� 1�dnG�w����b篹��{6OqՁi$���P�q�'O�Mq��9#��v{=yng�9*�6-��6�&��\�nvg-8�Μn�4��S`�<N�3)����k�{U����N��v��3i�l��$�A��8Bݶ.L�Dp%$r�XM�S�1� �uer9A����v��l]bQ�n	�xn,�Lk���=���h�^1��tR�Gv;i��v	wS�v[m���B0s+�u�)3�~�Hɫ�r�fg	��F�.��K��t��^[�3�����q��3ζ��!�G"xП���g�>��hWڴ
����s@����s�
8ڡs�`v^���[=l	�Θ͜�H�ы��F�J9��@����;��� �������(L�##����76:`6q��{W�R����ڽ����)CNf�^v���&Y���07u.Q��r��ݝƞ��q[�%Ҡu��V��}& ��F�t������pZ�:I���߯���}�w6q���� �l��b�|�"�r�s���+�� ���dF��ʸk�Z���M��V��ʫ��BI�bNI�nlt�;�8�콉�w6q�*8���Sq����4��Z�;f��v�h�W7��hQ��%$�;/b`͜`nlt�;�8�6K���۶�n�
-�v�0��'�u��)8�/��w<���.m�����> �l�sc����WPg�y0=*��24<��!���;������@��ՠr٠�U�DL��&EI�rIϻ�nIﳾ��8hEM��"��,� k�)�T'7.�M����8��J�I��8�rF��{y<�l�6:`͜`uv��@ME1d���@>�l�/;w4�v������T�X$���ؙ��K���q��z3�����U̠�^y����z�(I2BLI�>ݾ����4�ڴ�v��j����jc���0��0&^��;�8����;U���'q��I4�ڴ�v�=�{�ۚ��M�����(�]�L���	�;���#�GԻ�8ӑ,K��  "� ��[�z��Kı=�]��K�p�Mf���ֶ��bX�'�}���X�%�y�}��"X�%���=jn%�bX��w��r%�bX�Ȅ��vC�?^%2�$�1��E���&���?{G�cs;m�q_�w���:5���Y��{���o%�}����ӑ,K��u��7ı,Kϻ�m9ı,Ov�eMı�{������ˁձ�f���~���bX��֦�X�%�y�}��"X�%���l���%�b^}�kiȖ{��7���~���ꑚw��D�,Kϻ�m9ı,Ov�eMı���/���m9ı,O��~�7ı,Ng޾�5��Z���浭�"X�%���l���%�b^}�kiȖ%�b{��Z��bX�%������bX�'O[���)q�eї.�bn%�bX��w��r%�bX�wY�Sq,Kļ���ӑ,K��w�17ı,J���)AU�'�3�?̝��C�]�v��A���9	�����n�ۊM�()�#�T�!�k`C2��N��0\=��$5lv�.����]�v�-���qnm]�m۰��Sv\<	�޷����.q���r���5�<���5�p\�[z��v�^�\թ�U�i9���`��!�g&���ތ��������e{:P6�I�&G��x4W�Ӯ���Z5�e��5.�)�P_�7ϵ�M:�jI��=:�\���v��۫�q��m�D��ۇ���X��f�H�������{��'��婸�%�bs���ND�,K��l��Kı/>ﵴ�KǍ������6�HM�b�����o'>ﹴ�?��DȖ'g�l��Kı/���m9ı,O�������S"X��k����˅ѬՖ�kiȖ%�bv{��Mı,K���[ND�,K��=jn%�bX����ӑ,K=����~q�]j�8[�w��oq?�Dϻ���r%�bX�������%�bs���ND�,��2'g�p�w��oq��������[fi�iȖ%�b}�g�Mı,K�?w߾�}ı,N�~ى��%�b^}�kiȖ%�bD=���oV�Y�5���n�\�9�z9�N��s�=�[ѫ������J�s;9�����v�������?/v��	��t`�! �wI���bX�wY�Sq,K���ߴj�SXfL�3Y��"X�%���bn!	:���P�M�'"X�~��m9ı,N�Y�Sq,Kļ���ӑ,K���foZ�0���˗Z17ı,Kϻ�m9ı,O������%�b^}�kiȖ%�b};혛�bX�'ݞ����S.��)n���"X�%��u��7ı,Kϻ�m9ı,O�}���X�%�y�}��"X�%���d��4k.��f�%֭Mı,K���[ND�,K�{���ND�,K��~�ӑ,K����Z��bX�'�{��˛�� ����g�m`i� (�Y�I)��sn,1=� �IWN�I.�ʵ��~����{�N���Sq,Kļ���ӑ,K����Z��bX�%������bX�%���f��5�ִ[��h���%�b^}�kiȖ%�b}�g�Mı,K���[ND�,K��l����}���??�?���c�����~���bX�������%�b^}�kiȖ4t������>��)��8@*>�j� ^(O�2��MkZC�l�m�n��x���\6پ,a�mNRf �_y��#+��0"/���϶xE�t~�7�`��;¬I4PIJD <G��I�Po~X2�Є�Ay�G��S�<�(ٿ �9"Մ���BݟB$Pa�*�b��O"tND�;LÉ�S5������fSY�0>� ��oi�"���w��t��R�./A�vਾ�O "cJ
����c@q@�/Qz�b�b�PD�'{}���X�%�}�}��"X�%��;�Y&L�h��Y3Y�Z��bY� �@ș�}�[ND�,K���T�Kı/>ﵴ�K���"w��֦�X�%��w���.ŧ�V��߭�7���{���eMı,K�9�}�[O�X�%��k?Z��bX�%������bX�{�n�'�V�;�jM�t�E���00֬jy�m��:a��i��9봼qGT�vx|�іf�T�Kı/>ﵴ�Kı;�g�Mı,K���[��L�bX��l���%�bw���kYsT˫u��Z�ӑ,K��u��7ı,Kϻ�m9ı,O�}���X�%�y�}��"~A?�GX��bO�����Bn{ﷸ��{��?������Kı>�dMı,K���[ND�,K��=jn%�bX��ﮌ�e���j���kiȖ%�b}�fț�bX�%������bX�'{�����%��X1H��!�K`$R�H�P+J$W2 >��D�[��m9ı,����Y�kje�33DMı,K���[ND�,K�����jr%�bX�������bX�'��l���%�g���~��u��.R�im\�-��n���a�Ҽ���n�z�;��K<��F�3Y�fӑ,K����Z��bX�%������bX�'��l���%�bs>�iȖ%�bw�D�I�5�)��L�kV��X�%�y�}��!�U�DȖ'}�6D�Kı/���m9ı,O�������TȖ'����Z�D�Ma���nkZ�r%�bX����q,Kļ���ӑ,K����Z��bX�%������bX�'O{3z։��5�FY�h���%�b^}�kiȖ%�b}�g�Mı,K���[ND�,�� %�O~�ψ��bX�'�O��֭ɩ�V�6�Z�r%�bX�wY�Sq,Kļ���ӑ,K���͑7ı,Kϻ�m9ı,O�G��`�n�!��3�WZ����{J@�������I�Ʊ����q�� z�Vؠ�O# v��:�s�����s�;v,�ۍ�U��In��b����Zz�(q&�Rܼn�^z[Gll�Rs�ե��A2)��=�����3��M�S�W����mp���R��n{F�-ff�'̗b]��٪�6dT�0���e:$��m��u��^����W���{����_�߯����l����K���"]��g]j �eָ#�	:�OD�t�LҴ�j�u�2K�Z��X�%�y�����Kı>��dMı,K���[ND�,K��z��Kı=�I�]�˅Ѭՙ���ӑ,K���͑7�T�DȖ%�����"X�%��k?Z��bX�%������bX����M\�kk-̙��&�X�%�y�}��"X�%���=jn%����"dK�}�[ND�,K��fț�bX�%��� �F�Q-5}��oq������Y�Sq,Kļ���ӑ,K���͑7İ?�fDϻ���r%�b]��{���N�mq�:�w��oq��%������bX�'��l���%�b^}�kiȖ%�bw��Z��bX��~�#��ΒL1@m���wO�"�G[u��&�\ƃ�5��#d؝�p��#v�][sZ�ӑ,K���͑7ı,Kϻ�m9ı,N�Y�Sq,Kļ���ӑ,K���foZ�0����5�7ı,Kϻ�m9��!�p�(�SO�2%��k>�7ı,K�{����bX�'��l���%�b}��.��M][tۭkiȖ%�bw��Z��bX�%������bX�'��l���%�b^}�kiȖ%�bzwY/�M�fK�ф�թ��%�b^}�kiȖ%�b}�fț�bX�%������bX�'��z��Kı=�I�]�˅Ѭՙ���ӑ,K���͑7ı,?1ϻ���}ı,N�Y���Kı/>ﵴ�Kı?�s�_g�IvڰМ�B�6���i.p���X�ï3�cl�����z�]��{�Q,KĿwߵ��Kı>�֦�X�%�y�}��"X�%��}�"o{��7�������~v���Zj��Ȗ%�b}�g�Mı,K���[ND�,K��6D�Kı/>ﵴ�Kı;���tK3SE35�5�թ��%�b^}�kiȖ%�b}�fț�b��G�E�<#Q4��j%��m9ı,N�Y�Sq,K��Ƕ{Z�0ֵ�kWYnkZ�r%�bX�wٲ&�X�%�y�}��"X�%��u��7ı,Kϻ�m9ı,N��f���k.��Z�q,Kļ���ӑ,K��{���S�,KĿwߵ��Kı>�dMı,K�t���˙�1n�)��p�ۛ����:tȈ�V�S���14�yučΨ��[^�}����=�{�O������%�b^}�kiȖ%�b}�fț�bX�%������bX�{�7�q�຃Ssؠ�}����d����ӑ,K���͑7ı,Kϻ�m9ı,O�������S"]���[~K�G���V��~����{�����q,Kļ���ӑ,K����Z��bX�%������bX�%�Ox�[��Z�2L��q,Kļ���ӑ,K����Z��bX�%������bXM�S@TH 2�8 ��!���t���%�c�����A5u_{�[�oq��O������%�a�*W]���m;ı,O~�͑7ı,Kώ�[ND7���w�?��!�0
��j����
vR�Ǫz�!8=��'=\q�Kv]��y�k�:��j�浭Z��bX�%������bX�'��l���%�b^|w��r%�bX��֦�X�%�Ϗl��5�kZ�5���5�m9ı,O���q,Kļ�ﵴ�Kı;��eMı,K���[ND��2%�����Z�&�]f��&�X�%�~����r%�bX��粦�X�2&D�wߵ��Kı;��l���%�b}��.��ѫu��ֵ��Kı;��eMı,K���[ND�,K�{6D�K��#2&}�ߵ��Kı?o�����M�
Ow��oq������ӑ,K���~�9ı,K�O~�ӑ,K��w=�7ı,O*:�(zl���fd���Y�s5�aܼs��kP�=�rl2�#����?ﾍ}���מ��������ʒ��q�e��h��QA5s�MI��8�4�[�W�"�÷]<Ac<5��n����-����as�۶��.v�]��R8nܩs���v��MA��+�#���*:Y�ZA�a&���qd�5��@�u@F�n��+e@�cc�e�ݽV�V+��ww{��������ϲk>�r���)cnjI�,˞�m�cJT��`]�u˸�n��63�ꔃj�Vn�ʵ��~oq��������7ı,Kώ�[ND�,K���P�r&D�,K�}�[ND�,K��~5�0�XkF\��h���%�b^|w��r%�bX��粦�X�%�y�}��"X�%����"n'��2{��?���7��lu��}��oq��%���~ʛ�bX�%������c��)��;��l���%�b_�{����bX�'L/g��l�MS5uu�ֲ��X�%�y�}��"X�%����"n%�bX������bX�'s�쩸�%�bs��=�.��k֮��ֵ��Kı>��dMı,K���=�[O�X�%���~ʛ�bX�%������bX�%����&\�Y�.��g<�b9+��C<��s��pt�f����g�z�3F���ˣ,ִD�Kı/>;�m9ı,N�s�Sq,Kļ�����g�2%�bw���q,K�刺NSY�hշM����"X�%���{*nm 0$*A*�B(V�� H$��(��\lMD�.}�kiȖ%�bw�͑7ı,Kώ�_{�[�oq���~o�����&������%�b^}�kiȖ%�b}�fț�c��"dK�}?kiȖ%�bW_���~�~�~�~�`v�m��9�@��ֶ��bX�'��l���%�b^}��m9ı,N�s�Sq,Kļ�}��"X�%�gӾ5�0�XkF\��h���%�b^}��m9ı,N�s�Sq,Kļ�}��"X�%����"n%�bX��m���	�f�]^�2q:�)-�X惸v�`
N{4m3͈gvƹ����>����^-`���=�{�K���U7ı,K����r%�bX�{ٲ&�X�%����ٴ�K��{����߆�3չ�*����ŉb^w��ӑ,K���͑7ı,Ngݞͧ"X�%�{�kQ7ı,Nt��h��5��5���5�m9ı,O���q,K��}���r%���}�A��AT�&��O���"n%�bX����[ND�,Kǽw�5&�h̓Z�q,K��}���r%�bX���Yq,Kļ�}��"X��"w���q,K�刺NZ��ѫn�.��iȖ%�bw;�dMı,K�����bX�'��l���%�bs>��m9ı.����M:�T��2:��K�kb�/	��c�㶆q���r��Wj�w���ܗL�Z�-�dND�,K��~�ӑ,K���͑7ı,Ngݞͧ"X�%��ﵑ7ı,O{Rw�335p�Z�33Z�r%�bX�{ٲ&�� +��,O����iȖ%�b{=����X�%�y��[ND�,Kϧ|kVa��֌�e��q,K��}���r%�bX��粦�X�Ua�2%�����"X�%��߳dMı,K?b�J���LH$J7$#������T?�(j'���쩸�%�b^�����"X�%����"n%�`Q�@?���v!�y��ֿNfӑ,K�w�����85չ�����{��7��y��[ND�,K�{7q,K��}���r%�bX��粦�X�%?e˗S�BF%2`$�rd���n�G`�oF�ti��ں[�ɷWE�g�,�5�m9ı,O���Mı,K��g�iȖ%�bw;����F�Q,K����m9ı,O����4jL��E�kZ���%�bs>;��r�ș��{?eMı,K��~�ӑ,K������O�eL�bw�ߧ�\��շM����"X�%����dMı,K���[ND�,K�{7q,Kļ�ﵴ�Kı=;�?8+0�np3��oq���w{w;ݟwߵ��Kı;��n&�X�%����iȖ%��2'���ț�bX�{���ߟۑe��U��߭�7���'��n&�X�%��\���kbH$��_�5�I�}�lI�?�DTW��DTW��*+���*+EQ_�EE����*+�
�����
��E�(��0��D�Q�("�0T��PP � �H��0� �D�
,PE?�EE�EE�Q�EEh�*+򈊊��Q��DTW��Q_Ȉ���
"���(���(����b��L��[�*�� � ���fO� �Ͼ                  h    8 z��    (� R�  *� UAU*�
�  "�*���   J   �
�TQ�       ҂��� S�_jry�O��yi�j�ܚ}^� �y��3�omx�rn,��<  +��� h�   $h �  ��@,� >�� �  4� D �@   A@   "(
d�M��2 �1 2 Y� C�tp  @ 	��� :���{���������WR� �Rͻ��{�˛Sֹ����z��l�ҦMJź^�'U\ >�P    
((b �����  �  v`u{ń� }='��qj�-T�ju�<�J� }���t}z�y��p�۵y����U� 7.���R��v���ryN� 7^�sjusr��o�V���Ϡ �  �� xW����W����۶�6ꗞ} �K�;����z��þn��m��G���s��iw��o �^-�V�ݶמ�}����`r�m�p�n�g�����zW��]�6_^���+q۵� x����  (Aɠ���mͺ�q�}��6�S�v�� z7%g��o����ӛ/��]�@4�ʕ�wە���  ���+��ۭ���7zj��l���wo����U� 
g�K��6U͗Z���{��뭯 =H�S�JT� �T��53T�T�@h2d1�z�R���bda0MOb�Q�&�   5O�%O4�*��db40��IJi ��t������������,���W;����**+л�EEEuQO�EEE슊���**+PPT�����_�'�d����0�Є�`U��G-1H�15hFrG�5T�@`�4�T�=asS��T��dG(���y��{��Oѣ� �uⰮR�b��r�0��I��!y�=��Ny��f�"Vq�,H W !L4)�ώ�����r;���s��|~��y��#_f��`���:�'P��%SM�hK7<aV6,p548��	 �&�[�����!P��2�MM[��Ϸi����)��"l(8F�X���,R��0�r�HG^!疴���^>$
�(@������>��s�&W��< �"4qb�3�� ��A���dͲ�U��<9# @�`#%*_P�0�ҜHBb�p#Lt�F50e=��������FNKo�<2���!�Gӄ)�i��4��o�L!�E���ȔLc��$j2���z�Ԁ�!�H�T�)�2F���R����:c�ā�XX���(˼�qӄ8����_B �  ��%O��
g�ρ�+��)�jD�@��*2�pǚs�g�nߦ8���_}B	T#Xc��ֵ����EOG=<ͳ��5,(s���c�}��R�v@�rM��ĞZB�������e5���sd��d�@�
a�8�E���W�|��������W��A�l�MB�Ņ� �p��q���h���
C$�c�`�+�����c
�����b�� kCH0(h����y�b���J�7��i��L�����	<�D�R!�W�� Wd���J�8xP���D�	��H�T�-��hp^���i�N�-�,$����A���@�c�{����ݙ�Q}���r��G���#P�5!22E�I ��T�Q�� P�+�H�F!F41u!�3ōH����y<��B	_Mz	>r��\<���k� @��!�6��FI�>D)�>ߴ�iO�<щU��&�����K�����2��4$���B�1���T�F4���$$ ŖF��> �x8�$�8A�'�CЅ2��W��$�MxM.Px:�,*�*q�^k�
؍I1�$�M��TȰb�vN�~#fhp���:L��,C�x|M̐!L0�oG��.Q,�8���!L2x@���FF���Ǆ5����78�!P��'|���6Č�4���ϼ��)�F).\����y���w�6�$a0c����� ���Ja���o�u���]�8F�JY4���<�"A�o	@�2y��7=��Ct%�|�>�X�5!��0��<Ip�8�T��2{��\���[��[���{xĀW@"���<!sN_�!sF��%(p�`V$p5��CՉ#G�OyrCC�ؑ�� �U�X"'��HՀB!R4f����d"GO��\1��p�i�����I)[��k6�l�a�!��{������0)�s�����q�Ü%͑8����{�F5N>�6@H�㦔�.WN:��w����M\7f���#=<=�5������i��5�Iq�A߻�XT=L�Bx��=!��!���:�y.q��
Dc*Ka�]�_e1��	L�zS��<�$�[
(��A�'��p��S4�:K���,�OBB�x�.�$��⇠ీF� ��`���*®��B�a�E�b���=x�q5����i�xo����-��G�@�rn��y��+�_����8�$
i�'�a
$�0����@�����I9ȱ��f���H����i�|� "�)V @ 	S���$`��+�C�%q5�144ĥ0�(q����K�O%�<��'���fO/3�/�� �%pu9���/ϧ������1NQ��� �A�"���,�������<`�)	H�F�hB���$��J@����� �@�Ō���C���ő�(�	$�L�7*8��(� `j�X�k�Fp�F E��0���qO=�=���
Ip��5�xCR�ݶ��q����FE�ѓ=��y���04>4�� �����a XSNM \7�S�~<:!���?	�x���O�6C,ѐ�ᦋ�A)���<	rC�)!!��L�"D�$k�¡S4��)�)�9<b�H��o9�5�r�����(�b�O��s(D��0����}G���㦜<!���=�q�60���
�hp5�T�M�B�i9���!�"4`F /{vF\.���T�=�P�B\8{��`xMp%����&�p U�#���$
�((��Έ�}�\�"�!!\�D���J��@��=���WԊP��d9��Jc�p�@��= ��'U�@�JƔF Q�ƌD�I1�0��L+p��<@���	B{�z{�'�pXH4N*D�$�n��s�"A���ar+!X�a<s�������H(c���FP!|P�%pcaH��ᑴ�͵�)aj��Ǉ�C%p!w@��q���Ѕ0Ӂʛ���&ݴ���RE �o�^߰Ez�/͟�J���HB�4�0��ʘl.{�6�,��e	�a��-���b��b\�g�p���Ä�4�e�BD�ϼ��x��kB�)/�^ �gǲ��y�F�B�Yy�)���V�}��<�\��8�pN���VK2�a(Ƒ�5aH��m�,�Z&a��4���� @c$K��%4��H̙�ZadC���=���V-C �a5��76F�Q�U��7Za3�䲄�^2��+(D��3&k�xyM��y�rg9�Yο}�;���(�XV!4�`�-4�aaG
�X!��p=:�J&J�)��0dhF'��F�: @hy�'>�ι�%aH,� z�34�r@(��������z����O=��-�xz`4���\>�;p�O�P�$b������N� �A!Y��ԃ�� �
@��ס����,
Ɔ���N��w�P=#Eh���+�`h��$�T��p1���	��R_v��0��@*F��I�c"�jcM"H0�T���avr��C��ˉ��y�`R!"B0�1�4�7�=p��	aI|���Fh�a�^�!�w��a���B�ԂG���2Yd�\�������}!������¨��F/�D�:K��aM������ h  [AJ?`x �  � m��   m�h  ��om� 	 m��`�ڶ�m�`�m�ڶ�s�!m��ql�	��  �`  $��\H sm��  m �Ijڐ8� ���cj� �� ,T��UV�z����$V  � :S[�[�,U�	��ܗJ�`U�SГ.�.įh����|'��5�2�X6�q�
�VU����_�sڪ�)�1��7IV����S-ۀ`�8�]6�� ]�Ia�  m��-���i0   8�  ,�� 5����6�cm&۶ΐ$�uU+�쵵HL�49iV��uN̫.�NP��UP[J��,� �+���c��� �[p٬��;m��` ^�!Ƶ& �T��`���m���A M��m��m� ݶ�e�M% ڶ�gE�\ %�` �q� $��km�� [@l$  ���\�M���kև$|$������Iu\��T���� 6�`�� ������5��   [��htӪI� ,�m�mm�j�Y�P ��X@-�  �6��m�� �aa�H  8���m��ڗ��x �6�$6� p[BFٶp� ���v�X��m&�$p�m��   H p[@-�m�    6��7m�kl� ۤZ$$$-� 	md2�`�n�-�6Z-�� � v��,���e�� ������ݖ�@   �m��4[����8I�m��`�I�m�� �`   �6�ɥ6���o[%ͷm����[@ m��m $��`  n؛\8H^�����H��Z��궕{j������Uwm�G8C���m��   �Jm�m�ض� ׫q p mm�ݳ�Ih�m�imd` Hv�(	��[@t��.���$�8	�`��pAt�Ԭ�4�:��u.�nͻ]x�o�[n���� n�>��ht��I{ �p�.h�[y3&:�s�mu=��R)j�H�m[x� H  �$���   䜶� 8  @ Hl ��������   	M�	� [@j� -6p�!�l���`'AͶ  u�8H n��cZ��a ��mq����$$�8��� ����3/t76[l�v�p��J� p.Jf�6� �J�J�+��4@�9�� [j�m���m�9��/;F��z�t��� �X�s������6�   nܭ Hm� �H�c[rJ�n6ط�:� sm'e�   m�Y$�c��� pm�t|��$��׫m�N �� ���I#mRt�6�e��f�l !�@��`U�].
Q��8-�䄒l�� p $���[̐�)p��$�Q!��Hm����+��ѭžm:<�9�v���H�a�� :BC�-�M� j�$� l��-� �x �IlXa%��e�BA ���@�c� �dڋN��N� lݷ7U`m&nݤ��ko[h�ow�@��$ [@�bගN��ٷs+m�[@ ��mm�` h�X6�&B�`�$[��ݛj5�궪A���p�P�u�z�&�  9'[D��ڭ�Ut�S+-�I�F�d��e�59 ���mU@����U$-�"�n���pH �����H���M�-� �Tm6P�j*�zH�r]�f/K�mbE08sF�5z]�hn��UQ0�&X�^�Z꛺�Q�b�	%��y,�@Uq�z�U�ڕ`��We8�͵�d@��1S*�V��luJ���˲���Ú��U��'�nb�� ��l���e	�v*�۫V�nTz����T�d��-�n�s����I5�
���i��W�L�,�f�(uu� i6�Y��n�	-�����c]�q��C`u��p-���b���BM�5Cm�m�j]b�l��B�.8X[���) ܄�ں�T���Kjj7`��m��8� m����Wg��P�bU����۪�� *���VVh6�� m�ޡ�*� � ��UR�T�Z�m,�"�  ۶��m�q"@nѺ�n�$�d�V�5ꓛl�<����[pj�8  -��sm�   $H 8  H[CE۴���e�U3jV��
�W���v��۷Ӷ�� �F�CZ�`p�$ Nk�[׭�� I�kX��m��� ��U�S�D(���K�d�   �")kV� mH!S�R�f������8lm��)��m�` WR*��c
�c�p7%�^�n���3U	��Ҥ��³���>|�Km\Rdj���2rҒ�UmP@.ݲ�� ^� [A';E � D�kn-��H�@ [J��j�n �ڵ�ۜ���m��A#m��ŵm�����m��p�[(��Ͷ8?'��=��    ��]�  lm�Gn� ��{�IͶ�q��H  8$� im�n  -�8p	$6�h����� mI�q�];b�g-�m!'�s�    %���m����]e�$��֊W�Ӷ�m�$l�R/Zs�Y-кlڳnŽA�e�͵�ڴ��W/��{�:I6�H-���q@W*UuK�<�NPU�O
�UWJ�J�́<6�*���DQ^*�a���V7n�oi�n�mgfkgv���������ma�-5Ӷ�87b�b���nw�{ӧIm�E�mݶ�� �� � $     ����*�
y[���n�8���  q�6�^�� ���Y�PJ�6���B۷lm�s�q������{޶��2�JUU*7UuA�*ʵUTieUj5�Z���e��� ��m&��P�z�W�T�5�ڦ��h�`���n"`-���g2��e�Ҟ�U�W A�q�[.:�
�؃�XеS���ş-\m�p�L�	�݀���  ۲��e�n۱��kn�`p�it�D�e[B�$� ۶[@ 	��6Z� �m	8�� �t�Lٳl sE6� $  -�-�  6��=oP  $    8 հ�	 ͫ[p�kMm�m�r��  l�v  m�@   -�   ��NK( l   n-6;mme���mf�6�m�-� q#�[@ m�� Kh m��m �    s� � �����ڐ� �� [@V�      �`�� 	$ )@�m��8� m�[�6�,ۀ�}�  ��@H$h�h$��  8 @��e�[M�m�$m��  � 6�h $�ce� m&�m�6إ�� p    � �`��I�-� h�:ڶ�llD�յuK�J�uR�U*�9��$�@ ���    B��;����C �	z�k�� ���l�k�[�NHlm����0�\�٦���N��p�v�6�� V� 6ݍ��q�l6ͰN���[Cmm� p �m����a����m�H   �œ��m�q#[��K�� h�`�2l�26٭�`A� [@  $    m��$!��)6���٤��m��-�  ����6�!#� �5P�b�q���6�  ��Kh kt�`[KjB@C�ݝ�-�oP-�h���� �l �am�	6݆�&�m�mm�p��  Fչ��-�n� �N�d�K�p�cZ��G$�6*�Q�^n�T	�J�U��[́�` ٶ�� �#��m� 4턄��V۰6�].  mm  �I���79�ڪ�հ�L�r�M~���Ai&�h� m���$N��� m cZm&˒��� *�����@�V�G*  [گf���@m&�72�N܍*ʴ�O*��l����h�d�z�1��pRT�)q0J8Zm�5ٶ�u�sf��< �N�*���
Z��M!R�uP$�� �i�5K��P74��ۀmt��@q��M��� H��od�� 8t�� 8$�m��ۻ"\�*����ګwk��   �m����  �m�M�"Cm�6ͳ���wwtݶ�e�͓wm���N �� E��"����)��TO���tWU(�R(EC@�|�qO��_P|*OAR���N���E��poS��EP⊞(��|S�=D�4AQ=�@!�����C���@�`�U�z 8�D�|�@B
DV
����@S���Q��`�B�� L��bE"Ez> &���S�@x���-AF�'R"$�b!��T ��*,ASE=t�c �@	��(��D��S� ��<�z�qD:*�YN�D��B"@��>��t:
41@N�|�*�� � dD�U�D^�+�����>Sy@H��Pj P�O=z{Q*4@F����=D:����&��� � Q ꇠ�(���(D ��
�C�S�訨� O�"�@ ?n����}���~<5mR�ث�2qt��n� 59J����m
5T�̀�m����i<I�gR���k�+HZw@��ʢ������v��������:ؖ mɠ�4�O���.^yXHM��7��^1������<ǶUv��i��mլ�9%���6Zښ�:;�����gu�e܃p�H"G*��pJ�!�j�����P h
���l��v��[��Gjjy��)=�-����h|�t*7k0���c<[��=znPg�&ڶ�hr�ю��r�m��YC������[d;���u�pnȚ���Aٛ��z��-;c�Wkp�7�ѭV[0Ѻe;=�i�heh���U��K,
��Gq���i�5���Դ�����v�֦��{=�u��i]�)�N(1�ݓnV��v��7�hĘ�m��h�n�F��xH��)@�G7l�"��;!����C��i�2��k&R5�3�,:p�	�%�W�&(���vq�t�˲����^��{�5��L���v�$O���9�`eՃR�D��rD���yCn���hT�a.S3$u����\�!s�����w$R�p���5͵���;;���)C����z��XCCm;��1bQ(�:�յÁ��p�݊Ì�p7�F�G��V�:�Ct�{p��vn�Y@��K���\:^���_Z�5Ss�-BfƤ1��TKNHH��k�.�	��(�R�P[�����0� & �Z�� ��J�q���%Z�6Uݺe`6�t�@�mR���Ӎ�Wc���) ��m7-b�[�(h�f�@6����]r���˷b5c!s�4u�b-��q�l5�j4��Y�v�-�h
�v
Z�1�p�v�H˘	�s��QmYx��f�V���WAT�]�c9��uҦ�R�l����7!s���lUs���eR��>oo=���u�gқ,���i�S��c�n�z�%U�Lu��2۹�7 "���DN�B@ �B�# �D5' �����zDb��<�Yxu:kX�zv�a3Ӊՙ9��`��"�3����s'���%i�u����M�W2�`�V�B+g3�';�u�۩��.�0����r���x=q�Mձ��;l�ĭ	�gë>�O'. �16{P]W�a�ܱ���mK7q�^G\cjH�`{e��Ϋ�&[L��L�1�A�H�+M���;n۶Yyow{�Ψ��G�<��k0�72�Y �y���rg�99W�ܙݗ��C�r�����Cz���N�?_���3;��*U��rkL	����ƬVƄ�%��מI}��|�Vn�X&��3$���;�Pp�ŕj�^U�0�c��L�L`~��xwQf�8G*r�[p��&0=/�0K�K�l�P�S~%R:�k�� �wn�gu�7v��w sMd�6)~+�I%tXρ��	����vF޲<9��n97�Ͳ�wcv�1v�֚���������wv��w s�� �u�Z�7,�׀O~�w�����B
#  �	�� �A�'ϫ�~Tlz� ���Ҙ��UuQe)mn�� �;���ݸ�׀���?'�-��m��u�V s�c��S ޓ�`v�T��.�����r����������;��, �wn�M�R�8B�5o6g7fuf�.Yͤ�5�5�Z��N㶵����PBJ��E+��;�p� 9�ۀ~��x�m���T:������LzL`z_J`�c���kST�GY-vՀ���?l�60L �
+H!* �l�5V���� ��|�D�vn��;���j�J���]���K�LzL`v�i�oI��#�Z�7-�J��ݸy�ŀ���?l��|�������ky��h<;�7'/V�#u��/{n���v8�;Hi�}��������m������7����LzL`yWP��T��ʻ�Ex������)�oI���� �'^ګ�V��c���n� ޓ�~�0�1���:�G*���W����;��, �wnI��1b<x	��|��}?f��I���Ι.ffi+fQy����� ޓ�%0� ��{�s�����J�b�9e^8Q/B��o[C�ʜ�s���6�&@�X
�w��;���qb��Kl�`w޸훯 9��������w}� �`k'�i�e�r�`z\��7��oF�����]h-
_����m� 9�ۀw��X�������?>v'�Z���q�����S&�L&�X�2[ �I���-��c��TX9V s�� �I{{6� d��=��*N�
��AEĊJXH �L��3�n����C�V�mr��n��6�X�:��θ��ŭ�:��D[��[n�e���#�9�ݚJ��ѻ:w<�Um�vv6�j���et���(���X��{n�uq����4�#�SeF\z)�[�
V��ȯ/RmVN�1&^qÖg�[4�d9'�N�<�5z��,:c�.m�5]%�9�������\��%�}����nI��{��Y��M���E���u:��c\�jőJ�<�Wq�li�W�^6�����["�Z@N�-���� s�� �;��/�;�pۺ��Q#����yLzL`v�i�oI�K�L	�l�$��ꮄ���w s�� ��u�;�p�ֵ5AؤeR�y��oI�K�����I~���� u�lhR�ܶ���׀����� ޓ_�DE��(��ƃ���;h�����vO7V[u�᭼�󲚤�"+��R�$E�[mx�������wv��n���bq�U�mn��7y$��ß�U�E�����T�Z��U����������=�u��~}bٮ�Z�����X������&0;�4����.�Z΋�}��a������`7z���� �wn�wLqTH壩�+��;����UR�o��2n���rK`{cߟ{D Wf���=�����6KqvS�m�ە'k� �󶇉�«p]f�wF�I1��rS �&0����GZ��Kl�`wv�K�9��< �{� �{���4jsmhR�w���`~���I:�J�j��V�$�EI$�UU$�*_��7w�����)~�"�-�� ����������?l������U�ku�1��oF�I1��})�t��1�b�a�H�n����\��)�gս��:Ny�4^w/vģ���{�1��d�ҷi*�0�c��S �&0;z4����ʬt��_��[�~��x�ݸy�ŀ�۞I%�l��8�$rұU�ʼ�>��`v�i�t�����j��ISt��e��������o��&����rK`���IR_o�/�׷ sZַ�
Ԍ�[e� 2I��K������L̍0&/�u��}��C�/�'���][u.Օ�#���˰�=�''g���2\[��%�b{��ڜ�bX�'{��q<�bX�'�����Kı/{��Ȗ%�bt�ܐ�5��n����S�,K��{�'���dK��}���bX�%�{��yı,O{��S�,K��=�\6��۷2I��Ȗ%�b}��
��bX�%�{��yı,O{��S�,K����Ȗ%�b{�Yٗ72n����3H��bX�%����<�bX�'���Ȗ%�bw��Ȗ%�U$��׼*r%�bX�{����r��v�˛�O"X�%��w;jr%�bX��{���%�bX�}{§"X�%�{��x�D�,K�'۝���2ܔ��wJs�n�LvyU��ⷌ-�mY5���d���L�5���Xt�P��1X����xk�ӄ��;t)m���ؚ�K���]��1�m�Ip;�s�Vv���k���`�&*�s3z��x�%o6�ȭ�W�.�1B���-��]n�U��2hmY��u;\a7fPOk�������[�q�,��	RrC���nnk��t��V���3��7"���Edp��dL#��c�&hz�t\������oq������É�Kı>���ND�,K����<�bX�'���Ȗ%�bw�̚��V:�-r��~>L�3�ϗ{��ND�,K����<�bX�'���Ȗ%�bw��ȕ@�bX�v�S���fY�n��*r%�bX���w��Kı=��mND���Dȟ�~����%�bX���§"X�%��v��gwi�ܖ����yı,O{��S�,K��{�'�,K������bX�%�{��yı,N����f��Mۻ��jr%�bX��{���%�bX�}���,KĽ�{�O"X�%��w;jr%�c���Ϧ�9��ugY%�s�M�.a���ֻVW��Gciݖ��c�+���p"�ѷ76͹�L�8�D�,K�xT�Kı/{��Ȗ%�b{�����2%�b~����Ȗ%�b}������)��M7%�*r%�bX���w��8�>WblK��v��Kı=����yı,O���S�,K�����7.�7a�ܹ���%�bX��s��"X�%��{�'�,`$,K�xT�Kı/��w��Kı=����I�sM�f�6��Kı>�{���%�bX�}{§"X�%�~�{�O"X�%��w;jr%�gɟ-�5Q�$�uJ�Y��|��bX�}{§"X�%��P�~��ObX�%����֧"X�%��{�'�,K��
?�r��2�e���eE��Ivj{Xp������O��v�Y�.�\R�:�h�5�q��oq����}����<�bX�'���Ȗ%�b}��Á�D�,K�xT�Kı>�i:\��!���ۛ��O"X�%��w;jr%�bX�w���yı,O���S�,KĿw��'�,K����!�6k��ݹ��jr%�bX�w���yı,O��p�Ȗ5�7�R� �D4?)����Y�ԍ%H2IC�,����M�I0:a���b�Py�
�4JŅcV��|��DX�q@���*J����8=K Х� �B_BOL�}�"�A�$������I�A
+��� ��
����U| \aQ��:+�#���D�P�#���AG�>x��^�?(����b$D �Q!�;��o��@'�2%�b~���S�<P*dK�����m�ͳnd&n�O"X�z(�2'{�<"r%�bX���~�'�OjdK�����S�,�F@�ȝ����Ȗ%�b}������)�n�g�M��"yı,K�߿o�~9"X�~��jr%��ș��~��yı,N��p��c�L�bX�����?a��,)rM�wf[�]qqdv�#*!�u`{C���_n��Q:��Ig�a�ܹ��{�!�2%�����S�,K��H���ޜObX�%����9�Ȑ2&D�����<�bX��(|��C�D�UG\R�[�a�gɉbw���O!�D�DȖ'{�8D�KR"_߿~�'�,K�����O�".�Ȗ'��ә�l����]&�m�8�D�,���?~����bX�*G?~��x�ı,K�۟�ND���"dO߿~��yı,K'~wf�2�ɿ�n�O"X�%�~��x�C�$r&D�>�����Kĳ� ~����ؖ%�P� � ��T �C
Wਞ�����O�y��9�ʙ����t���Hf��ws7��Kı>�����Kİ�G��u<�H'�w4�H$���}��$�y��vnn�\nɒs�Y��w&�fz�\�sŞ�$S+:�s����+ۭ�y^�+A������d�{�'�,K������bX�'{����%�bX��s��"X�%��{{��:m�ͳnd&n�O"X�%����9ı,N����Kı=��mND�,K��|8�D�,K�>��37,�ݺis3H��bX�'{����%�bX��s��"X�%����O"X�%����9ı,N����f�ن�5���O"X�%��w;jr%�bX��{���%�bX�}���,K��{�8�D�,K��'&L˚l�p͹��"X�%����O"X�%����9ı,N����Kı=��mND�,K�N���0�H�o"gq���mx�� ����d\@���^yy��2.�[c�j�]��AD�1�)���f���2rr��t���"Z�TW�|c�H���v���Аn,���e��۷Kcl&1�R�J��M�8����䴌���ї��m�+W.�g,�z��av�[��&�Ѵj�:m��J�9�Bk����"���unɔ��p�/=�߮�J��z�[�;/[[)��1�/N�{N��u������r:�ˋe�«�+�{�{�oq��O�]�*r%�bX������%�bX�}��S�,K����Ȗ%�bY�p�]ٴ�.��w6T�Kı/��w��Kı>�s��"X�%��{�'�,K���{*r%�bX��iz\��!��Kn���<�bX�'�nv��Kı>�{���%�bX���eND�,K���x�D�,Kӻ�C�l�3	�s3v��Kı>�{���%�bX���eND�,K���x�D�,K�;jr%�bX�g���C����6�I3t�yı,O{w��"X�%�~�{�O"X�%��۝�9ı,O���q<�bX�+�kj,�N����Z+@+i%(�7h�I�H��v�ԶC]:��x9�J���	�4�tE�e���"X�%�~�{�O"X�%�~�;�9ı,O���p?�{"X�'߷?Z��bX�'~����7m�u�37x�D�,K��wjr� dE(��blK��~��yı,On~�9ı,K�{��y���>^���#�Q�-,>LK���߼8�D�,K��v��K���/~��O"X�%�{���9ı,O���t�s33l�m�ۺq<�bX�'���Ȗ%�b_���Ȗ%�b_���ND�,K���O"X�%�g���vm3�6ۻjr%�bX������%�bX�ﳻS�,K����Ȗ%�b{��ڜ�ϓ>L�y/��{L�~���@W]��[��G*k�"֢�wNLᵧ����)�v7i���.n�!��Kn����ı,K���jr%�bX�w���yı,O{��S�,KĿw��'�,K�����6뙄ݳ3wjr%�bX������%�bX��s��"X�%�~�{�O"X�%�~�;�9ı,K糷0�M���m̖���yı,O{��S�,KĿw��'�,h�_��=S�Tt�O"_>��ND�,K��{�O"X�%��Xw��)�n�e��S�,KĿw��'�,KĿ}�ڜ�bX�%����<�bX�'���Ȗ%�b}���,ݷ5�����yı,K��ݩȖ%�b_���Ȗ%�b{��ڜ�bX�%����<�bX�'�t��R��2~�fM�e��%��jr�ݸqrCi<���{�]�'�ZɅ�܃��(��v�=߭�7���{���~�'�,K�����9ı,K�{��yı,K��ݩȖ%�b}��5V�rV:�����~>L�3�ϗ7s��"X�%�~�{�O"X�%�~�;�9ı,K�{��yı,K>�^��ne&��nm�Ȗ%�b_���Ȗ%�b_���ND�,K���x�D�,K��v��Kı;��t���!��Kn���<�bX�'�^�Ȗ%�b_���Ȗ%�b{��ڜ�bXj�v&����O"X�%����!�m�3�374�Ȗ%�b_���Ȗ%�b{��ڜ�bX�%����<�bX�'�^�Ȗ%��{�����}�q�2��x�:g�>��qY���p�tW�+���"4�&�㮆bm̖���yı,O{w��"X�%�~�{�O"X�%��׼*r%�bX������%�bX����p�̓�t�-ݕ9ı,K�{��yı,O���S�,KĿw��'�,K���{*r%�bX�z���K7m�u�37x�D�,K�xT�Kı>�{���%�bX���eND�,K���x�D�,K�[��2��.�0��*r%�bX�w���yı,O{w��"X�%�~�{�O"X�%��׼*r%�bX�}����ff�tۛ�t�yı,O{w��"X�%�~�{�O"X�%��׼*r%�bX�w���yı,N�g��wn��f�K�=�{`���챖�g���-u�[��&Ϭ�;]mk9��X���.giKpv�]pJ��c/gr�(�[�ێ_KǷFP�-.�q��û\�j��
>s�iW`v��j-Ѧ��jp�A��k����gz�f϶x��!�+I��5J��Q�D\Ý���W6�	]�iB1#�E]�Ӭg�g�����;)�/$��䢹�2��X��"d��x�D�a��m�ͷ9�Ͳ��;�G^�Z�rm��*{ı,K��߷��Kı>���ND�,K������Ȗ%��뿥ND�,K��d�Oۻ�3r�n��Ȗ%�b}��
����L�bw���O"X�%����9ı,K�{��yı,N���!�m�3	�s74�Ȗ%�b}��É�Kı>���'"X�%�~�{�O"X�%��oxT�Kı/����칻�m̒f���%�bX�}���,KĽ�{�O"X�%��oxT�Kı/{��Ȗ%�bzg��w2L6��K��D�Kı/��w��Kı=��
��bX�'��|8�D�,Kﻜ"r%�bX��y`{��x̣�X�.:�g�G5iڍ]�Q#�ee���{G�cv�ƴ7>,������%�b{��9ı,O���q<�bX�'�w8D�Kı/��w��Kı>�0�3.n����ҧ"X�%��{�'��!�(@�B��(���1�'�,N����,Kľ{�w��Kı=��
��gɟ&|��2j��IX��s���1,Kﻜ"r%�bX������%��a�2'߯�9ı,K�߿oȖ%�bY�:�ݛrfۙ���D�Kı/��w��Kı=��
��bX�'��|8�D�,� �"w������ϓ>L�{����lD,�����O"X�%��oxT�Kı>�{���%�bX�}���,KĿw��'�,K��ӸgM�ad�3v�����;jq�������S�+nyy59.1���4�u��n���*r%�bX�w���yı,O��p�Ȗ%�b_���Ȗ%�b{��9ı,K�c����a\�KV|�&|��g˽����r&D�/~��O"X�%�����ND�,K���O"X�%��[N���)�n�\��'"X�%�~�{�O"X�%��n�T�K~V���"r&��xq<�bX�'�w8D�Kı>��;�l�f���3w��Kı=��
��bX�'��|8�D�,Kﻜ"r%�bX������%�bX�vݘt�37ar���S�,K����Ȗ%�b}�s�ND�,K���x�D�,K���Ȗ%�b{ٶI_�I�$��3pn(��V�=-��FU��ñU����<`�n��u�V1t4W|�~����{������"r%�bX������%�bX���eND�,K���O"X�%�I�:�ݛra�-�4�Ȗ%�b_���Ȗ%�b{۽�9ı,O���q<�bX�'�w8D�Kı;���m�"J�v�s���3�ϓ>\�vT�Kı>�{���%�bX�}���,KĿw��'�,K�읻�:M��a6nf�ʜ�bX�'��;8�D�,Kﻜ"r%�bX������%�`xy� i"����j� �U�Ec E � � P$P��B� īB@�bE�H�w�O�7ؙ�J��bX�%���\��˻��nd�7N'�,K������bX�%����<�bX�'���S�,K����gȖ%�b}�ܼ��
lR,�+�ӕ��7m�� tn�w�R��#�/�N[�F]����[����X�%�~�{�O"X�%��n�T�Kı>�y���(�bdK��g��bX�'~�C�y�͛sLn���'�,K���{*r�9"X����'�,K��g��bX�%�ﻼO"X�%��mهHff�.\0�͕9ı,O>�|8�D�,K���Ȗ?��lM�{����<�bX�'���ND�,K�9�6\�̛v�̻��Ȗ%�b{۽�9ı,K��wx�D�,K��T�K��"{�߽8�D�,K�v~;�i�m�fnʜ�bX�%�ﻼO"X�%��T�{y�T�%�bX����'�,K���{*r%�bX�C�(�P�E �BBAB��> u�c{��,�3Qp������>��~��򟩠'� ��,P0�D��Y�����,�1�!�v�M@��8{��#�EϘJ�� <��8�=ďW��I}c�$K�{'��@�#$s�z���<�4��V ��,"�b$b=:�"�b�<_U�:u�D��ֱ�#
o�5W��f@����b� �����?!�D��/�<�V(D��9��5�0����T'��S�	�z��P������F	ȁb -���oo{�~���Ǖ�kj�*���6���ڮk��(H[5j���5������\��К�Nd�I۷=���QtUe%[�Q��:����7t�%�6���[Tl��R����$ I($m*��Km��H�a;:s�rcZ5ń`{[�1�-n��t�S��Dm/=K�;r���E�۝�R�Α�p�۬��+U���q�Tkm���oU)����D�T�� 5)t��2z��[M�ݗa\�V�>��^ͱiD"�Gj���
 r��h������3�jv�w�j�%�޳�v�6W��z���wYx틶�K.^�%��A���m�`�k!�rI�^���n�u=u���E+PW;��?�ջv� �q�>s�[��Hrnw��3.36[�է{Tu9tÔ�8�^�0�{si��Y�c��u��\�A�vx�l8�y���g��]d�/cu�N�G]�é0lOi�<���[@;Oi���s�(3���]��e��]���R�*�TaB�#V0���mXs��r��È�[Bm��W4�&�2�#=x5�R��J�K��Ol�Gl�Nɢ�Jl�۠�٥m�f�R�Gs��SR��թ��6;eUpv݆��>˘H�˳m�;�����B\��R6k�๷h
��Ǘ6L�`��5vش������_$�א�v�y��:��m��;���v�Ss�6{ �h�� v^�;0��[uV�s[�YfN�z�z�ŵ��ֆ�g!22�$��	�ۃ�6���t�������+۷9v�\b���v���m���^Uぁ�$2 m�F����]��z��6YĔI�v;X�3�۝'6�`��U�̶���V�[���4��m�2��pO0��#�;h0$��h���KKM�*P�6�pS�,��P�k�6�<TBnS<d2@I[!�H)Ie�.�v�}9�Β�]Rg�����/;-�M�n�8t�tm��*�����@���w�@(�8(�A��x�'P�O�Q���<;y�Y��9�Ƹ��W����FX�,�੹ƛqOU��:Yh�+M8EicN�!����$��l��CΫ{�v��oJ�E�Y���9���ꗶܻ6d�8��d�<�[�M�]�K �g�rI��3����ۡ�1�3	k�7	�A��l�������;m[���vy;8�K��A،j�X�mT�pG��k/<n�&���+0�98i]���̻�nI.6ԓ�ݒ綢�]�t�j�K�g6����ѤTe�"J�v�}���gɟ&|�����Ȗ%�by�{���%�bX���eȓșı/����yı,O��w
~&�s0�73seND�,Kϻ�'��G�+�6%���ҧ"X�%�{����<�bX�'�]�ȯG�ɟ.t�8ʻe�r�jϗ�%�b}���S�,Kľ��w��K�dL����*r%�bX����É�Kı=3�iۛ�%�vi�[�*r%�bX����<�bX�'�]�Ȗ%�by��É�Kı=��ʜ�bX�'�ޔ���3l�5�37x�D�,K��T�Kı<����yı,O{w��"X�%�}���Ȗ%�b{;&�l3����7p�v V�rk��1���:�FLP&x�&�m��s��܅˘nfʜ�bX�'�w�O"X�%��n�T�Kı/�}��yı,O���S�,K����gM�33&�.廹�Ȗ%�b{۽�9Q�@J�bX�~����%�bX���ʜ�bX�'�w�O"~ ��,K;O��vm�3e̳7eND�,K����'�,K��뽕9ı,O;��q<�bX�'���S�L�3�ϗ4���(�r��[n|�	bX�'�]�Ȗ%�by��É�Kı=��ʜ�bX�fDΝ���yı,O��w
~&�s0�73seND�,K���O"X�%��n�T�Kı/��wx�D�,K��T�Kı/��wlݙ,��s��ʏ���lk�����piݖ�����vr���d�ĵ�=߭�7���{�}��S�,Kľ�}��yı,O���S�,K����É�Kı=3�iۛ�%�v�[�*r%�bX��ﻼO"X�%���{*r%�bX�g{��yı,O{w��"~ ��,N���?n�&���a����%�bX���ҧ"X�%��}��Ȗ5���b}˽�9ı,K���x�D�,K�K�����\����ND�,K����<�bX�'���S�,KĽ;��Ȗ%��|�קʟ$|���TrI
�v:����Iϯ�6	 ����'bX�%��׼�Ȗ%�b^���'�,K��N�W�8K37i32�Λ��:xr�)���O��E���Vn���We9��Ѳ칖f�Ȗ%�b^��w��Kı>���9ı,K�{��yı,O{w��"X�%��f���wp˹srY���Ȗ%�b}��*r%�bX������%�bX���eND�,K�w��'�,K��N�&�30�73wjr%�bX������%�bX�}���,KĿ�w��Kı=��*r%�bX�{;˒6��˷rR���yı,O��p�Ȗ%�b_�����%�bX����9İ>T?EAC9�����yı,W���@N�u7$��a�gɟ&%��{�O"X�%��oxT�Kı/��w��Kı>���'"X�%>_�k�1D�16���(�1ۡ8�EP�:��v�u�/m�fyL��f�l�fn�<�bX�'���S�,KĿw��'�,K������bX�'�{�'�,K����ä.n�.\�st�Ȗ%�b_����~T9"X�����,K�����'�,K����*r%�bX��ozl���6鹓l���yı,O��p�Ȗ%�b|w���yı,O{{§"X�%�~�{�O"X�%�~�^��l��32ۚD�Kı>;��q<�bX�'���S�,KĿw��'�,K������bX�'��I��wp˷3l�����%�bX����ND�,K���x�D�,Kﻜ"r%�bX��|8�D�,K�jO��F=�y��34��d6�J5�rt;/Y#Nћ��
mLn����bt��0;;��x1�꽗k �PB�ڇ���w��Pk/w��{�M7���[�Zv�Y`0�{ZE&Y:KF�p�Nr#�gc��<C�%�sI\Gb��"<�i�L��Kdy���*r=S����Z��xz-v���6�3���u�+pk�S�RyڇZ���+h`A�0_|��W��w]�vK�U�^շN�Bb�*l&������=��G
��3���W��u�M�&���ҧ�%�b_����O"X�%����Ȝ�bX�'�{�'�,K����*r%�bX�{;˒6��˷r[st�yı,O��p��"!��,N��~��yı,O�_�*r%�bX�w���yı,Os�i�ɹ�f˥���ND�,K��Ȗ%�b{��9ı,O���q<�bX�'�w8D�Kı>�zS��,͹wd1�4�yı,O{{§"X�%��{�'�,K������bX�'�{�'�,K��K7����̙���S�,K����Ȗ%�b}�s�ND�,K��Ȗ%�b{��9ı,O/�}��Yz��g�^�g5���zu��t�-r�����]Ǒ�ۘ��ź�u�WE�뢻��Kı>���'"X�%����É�Kı=��
��bX�'��|8�D�,K����vm-�˹%ݑ9ı,O���O!� �DȖ'ݽ�S�,K���Ȗ%�b}��dND�(eL�b{�m'����2�Sst�yı,N���T�Kı>�{���%�bX�w���,K���{���%�bX���S�.�favnf�9ı,O���q<�bX�'��6D�Kı>;��q<�bX�fD���§"X�%����̰�m��ɷ2[st�yı,O��l�Ȗ%�a��O߿zq=�bX�'_�*r%�bX�w���yı,O��n:]����x6��n�gP���&�ԶCV��	��Ή�S�K�6�p\ݑ9ı,O���O"X�%��oxT�Kı>�{���%�bX���,>L�3�ϗyu����]v����Ȗ%�b}��9���,N���É�Kı;��6D�Kı>;��q<�bX�'~,�:B��2d�nn�9ı,O���q<�bX�'��6D�K���؟�O"X�%��n�T�Kı=����s33m�w&�wN'�,K����Ȝ�bX�%��{�O"X�%��oxT�K���ȝ����Ȗ%�bY;??�ٴ����f�؜�bX�%��{�O"X�%��oxT�Kı>�{���%�bX�w{�'"X�%�ߥ���c��h��km�G*A��5��6�l��j,�,e�O���䉸��'�,K���{*r%�bX�w���yı,O���S�,KĿ�w��Kı;'�p�v]������͕9ı,O���q<�bX�'���Ȗ%�b_�����%�bX�v��ND�,K���e�v]��.�nn�O"X�%��w;jr%�bX����<�bX�'ݽ�S�,K����Ȗ%�b{�[N�nfXn�.��͵9ĳ���2&t����<�bX�'_�*r%�bX�w���yİAx'Q�s�3���'"X�%��}�;��ۛv��f�3w��Kı;��
��bX�'��|8�D�,K�~�br%�bX����<�bX�'�I��R��?M�fe��*u�]N'���m���}�sܺ�9<u�Ʌ���/]���-30��*yı,N���É�Kı;���'"X�%�~;��Ȗ%�bw��9ı,O=��tۗ3&�ٙ6���'�,K��ϻq9ı,K���x�D�,K�^���ϓ>L��wo�$�p��{�J�%�����"�ް'�i��]�wz��ɯ ��h���u�SMYn��ŀ$���L���������"��*��0�cu���I�	��X��[����d����"i�Y�p����mLNƲi-����n>!x�md���[OG2�`�[��:7%v8z��#�f���y�R�v^t�9':��Sv��cV�6���*��r�9��7#����
��A��6�m�Cp<ǔ'mYi,-��8��n�jv»7½c$gf�*��=�ۏ�jg�g�^�[�rx�,����{�w�����q�mMN���9�v�z���Q��r�t7�+��	��"�0�I7]Oj3�y���)�r�cl�0�c���{r5j�����V���|���ذ��� ����;ɭm�m��:.s�`OH� �'Y����5���s�K�9iREm��/�{��`l�� �$�T�sw�`�9�W�ڝ���p�w�}���֘��`%J�5�ˮj��s�rI�2��L��ᔖ��;������j������
_�֕�Kk�r���޸�w�����0��`�<���G]��.��I�{�R��"�;��0'ti�r�1�{���
+��]Y].�Φ��0&di�vE7z���k ��m�Z��X���{�ŀ�N�'�i��n����˻�xm����
�Aw��r�1�6F�$i�;�ŀn�g��yc�(�pjJ뫕��I��R���������G��Y7��m�*�1��As��w����0=24����⤗���� �M,^BrЍG��gF��4�9l���#O��6|_ث�K]R�Uv�۾ŀ]ݸU�j��=����p�Ukh:��A"��9� �@�]58���}�!���-MuG�@8����x���|9<j1��"c5Q��� �GH�ubpU��$�KR�p��#hV?/"@���]A�Q	�`	]x�DC��� � �@��D	�
��4=G� >����E�?!������{ p]߷�
�%��9S����X��0=$i�3#LЍ��b��*i�m�7���}�{ߗ��O�`�L`u!�V�b��]̽=�Ņ!�% �qq^�W6H۪w4y�ۗv2�NF�Tv
8:6�X7w���`�N�J��ɭ0<����/��x��.��oF�)&0&�i��w���6�j�F_�*��ݬ	�`t��ލ0;nR��UU�ef�,��ލ0$��ލ0J7�7n��K�9iH��Հl��ލ0����Ѧ�Z+�}���`�uQŻY��e�n�[r/=u�kg�����)<v���h�������`	1�7�L	$i�x]?O�fUy�X]^&Гz4��F��w�Hѩ�(벦�%�ލ0$��ލ0����Z���Kr�$���~X��ŀ�v���,��� ���b�n�oF�BL`M��I`w�[C�`aL>��C����m��a� =%q;�nL�=���q�:ۙ(����]�cL�A�QخVs \�(�U�.N�����CX.v�[*oM���N����`�Jm�=��R�V4sHj9�h\��\�'`�q<��;+E�ki,mkq[t��7Pc8�5�T�OW�+:�[;,���*��cB�xەLv�4�Ig;��w���wI����*�f�����a��f�j�u�����iT첾�GƔYC�$��~.�pi����Ѧ�4��Ѧy5����]����� �wq`$i�7�L�&07N2�B���t�e�&�4��ѦГzb���6���a,��V��������Ѧ�4�<.���*����� �$�ލ0:H�oLX�����շ���I���ROv�-ϒI��I��j\�����n�vMR�Qx�Z��`M����0&�i�r�n��}�F�,ptmʰ��,��/�A`b �R�U��ɾi�~[7�	�0?/��,ʻYvUy��7�L��{q`��X:A���I[�*���U]	xލ0;���i��o�m�m��`+a-�7��Xww7�LBL`rపO�H���U�Ole���P���Ȣ�e���v�b	g񙑂��U
KB85���o��X� 7Mۀo;���z��\r)jvZ9��7�LBL`M����0=K�ſZ�-%rJ�V��y�ł�T8�� @��*�8�4FbA��@|������{�߸`�F�z�qGK*j+-�7��X� ��Ѧ��U�B"��Օ�U�&� ��Ѧ�wq`�׬���%v9
1�kqW��)��*�˃\��y#�ć\vz�
	�7^Z˰���`N�� ��dk�������#g��cR�eTvՀcl�0:L�wF�l�̣n��P�!-�7�����0�w n�� ���Ih��Q[j�2rK`L�� ���QU$QUI$��}ܝ�ŀ�Tګ$���eY����ѦГdi�%�L�S�('�;~D�ȅ�J9n^���|s�ӻu{3�uhy�(/:��ag0��BL`M���%0'ti��[F�v����5)-�7���ٺ�	�`	1��]t"+��]YXU]�`IrSwF�BL`M���u��SS�X��r�{�ŀ�L`M���%0=���Yt�(Ņfb`	1�6F�\���ѮI0K�
�IJ�@��t�0u�ݲ㳵@A �ֵ����Ջ�Ѐ�zLL�vj6R=lt�nftYy�ݲR���Mu�@�<�X��r�@m����͹۶�-�Lt\�{��Ozʃp�(<���H�Vث��3&κ�X*ON`�c�F��p�X̓��G#���D�2l�ظ��n�#Z2�v��{���:�4-r{��ݝ�nXB7&���)̶�8e�l��=m:u����ќ�3�(oA7h�]�+� �OdJ�ѷKc�R������7[wF�BL`n�aj!]���V���0$��I*Wfɭ0	��X۸��:M��IH�vUl� ��q`BL`M���%06�%)�,0������ �I�	�4���������^�\D�ʚ�����L	9%�	�:�2u���^��{˝�����&l�����=r=�C��A�p��9#<��g�7k�w#� ���>���7�0����Ѧ����)��,���r� �wnw���f���*K�a�I�ލ0$�)��]Q,&]�Y�,X���Гz4��f�������mt�:�)	n7�L	&A�M��&07z�����c�[j�7v�{��O��_��޸� ��7蚱����ð��9���A
9znC[��z�^=�mk&N-2��Y$�u;*�� �wq`tݸ�w��L [����(ܰvBLL�&0&�i�$�0&�i�z�^�\D�ʜ�� �wq`�t���~_��oF��&0=֫�����Օ�U�&� ��Ѧ�I�<�_$��{��9�7Zjy;e��rQ�;�L��di��d/���ĜI��t�uZ�7d3����m=�ڀ.8Ol:�������;|���u�Wy��}����#L� ��Ѧy6�6�l�}(�� �n��|�I�7{�d֘)'X�\w��_;юHEe� ��׀o{�����5{޸��b���mU�JGS��exI+�7�`n�X�4��UN�T�� >�u<����I}��騣��Y	*��ݸ�K�w�������7��X�ɴ'ҁ[,���n�VM��5sn�=ɮ<��{���*p{O�:�q�*qYn��ŀwf��7��^I|�05{޸{�6!yW`�����:�9%���%J���ߚ`���o7q`΍ؚ�����m�^3#LRF���U+��֘y�l�6l�(��T�Ձ����z��~L�֘9%��%T�^ɿ�g6�6�l�}(�� �n��;�u�߻ÒI���y$��)Pn���������S����@W�bj�
�j�}T,X�2���$@�J� �5> P� IQ1��b@:!��D�>#�<!�5WT�^�B@�>��O~U��}�\Q�D�4���(D�^�TO����2qH!<�>�BE:�D�)�PMB$���2��`������~ H ��e+m�q�k�ګv�lW]�m�Y��l�6�{m�خ9x��knG�-��k�0J���`{2�؄�e*���ͫ�����Ie�84�XI��&�N{v�y��\ mYU3=/  \YZ9܁����s���`Ĝ�2�uٝQ5\��'@�+�{U�.�	�KV�]8�j�\�P��.�]h�n�E��l��d �<�)G��olN���GmE�.!�hC<j��ʰ�<ݱpl]!gC�A�n4g�D��`�j�S�K�iĜ�Vm�7g����Z�nݻ5Sv�.+{{ �¬j��N���+T�k!\v�ɜ�X]��V�j�뭌��9�v.��/gA�v�oO[��\��k`�����:��v�ն3��r���k�=����\h����ݰ*ݽ����y��	�-����)�.�#L�p����NGs3�+N�F&����3s��z�9��b5����U�U+�Ϫf�3�>HJ�ES����\�#m���O��ӝ���`����B�T7L5Z��;i���|(��nk.y�:5��;R���u�[(��]J�9��+��3yy��a��:��<4W���%T�֛C��`c��К�;;�m��;r�Zbv�6͜E �.ɻV�Z���U-N��ʏV6���X]���3kI��qZ';� �M���r��ە٪���v�v:�лJ�U*Ú��Ŵ�h�d��Zۃ���c!��8�*��Ywn{.�f�j�Ӱ�ղ��͍*򪼰<Rҡ�xK��HJ77d�Y�%�⍆�61X}�+�-J�m�ΓG6�t]yV�2�n�[n�Mkf�V�4n3�s�y�y���b��{��+�9�����@l�D�����6��դ�$F�v��[7e�nj��<:͂E�QݝOnۥxζܯ#ps�{`�r,�S�U�b��[{hS)���d�f�ܷ4����8!��ujE�1@B��Ꞩ� GU�����͓&���h]���a.�۞
�p��j��#�z�:t<��hP�:��9����9����.:�K�ۗY�/H<a�ܽ�]J�UL��8�g�s��p�+�����*pͱ t��	^gZ�חtb6�r�Efwmpι]ǭ�m�J�z��]��r��Z�����[]���[�������a�P��n�̛�v4u�۞q�y�v}�\q�+f˩�h�a7]1v:�秨�g�W��uϗ�ݹ�\�����w�>;��ӒYj��=�����ݾ_|�K��=�{ s�'���TGS�I{lfN�1I`OH�'$��U/�l��~�E��]� ��{6F�.J`�cV��*VeZ/�}�������RI^�������`2\/��'����w�Sb�lptw�u02rK`2u�UV*J�T�E��|�����~����llli��;2Rɰ�\��n��7l��D�')�\r���U���3%���ۓ6Knf�>A�����o �`�`�`�����|�����~����lll{��?N>A����m��I�nL4�it���|�����������G�C�b�Q�T8�{`�`��������lll}���^>A�����o )� ��A�A�vO�ݖݛ��9������lll��xpA�666=���x �[��o �`�`�`�~?~��|�����v��鐹�is2awt���lll{����A�6667����>A����~��x �[߻�Â�A�A�A�A���g�6���e����A�A�A�A��w��A�6667������ � � � ����|����{��^>A����v�^�2陴�j�sJ[�y���k�o;'8��[x{xi\��C��Y7l5ݐۗrf�ww��A�A�A�A��~�>A����߿xpA�666=���x  AO`��A�A�A�߿o �`�`�`���%'��wn6��nn�A�666?���Â�A�A�A�A�w���� � � � �������lllo��߷��A�A�A�A����M܅�.�s4���lll{����A�6667�{�x �yTa�����Z��Q�Ox��v7�������lll��~����lll}�o0�~.�\�d�.m���ll_�B"�����x �����x ��~���� � � � �������lll{��~�~�Ɇ�M.�3w��A�A�A�A��~�>A����߹�pA�666=���x �����|���|��_{}�j)�s�d��@�P���ˊ1l�VtAܚ�Y���W��<.,�Uc]���9����A�666?�������lll{����A�6667�{�x ��������lll~����L���K������ � � � �������lllo����A�6667������ � � � ���?N>@S�9�����?��33I�K�nn�>A��IU�T��߻����URJ�s{�v{� ;���hQ��U]� 8�gXӰ`frKa�R��z��K�UJ���9��\{���W��
�� �2뒘��5I1��������tl���3�n;e���Y7����S�V�S��8���s���ظ6�ڍ����K��`�c �$�ِ`z�55:�8�+��v�I|�u{޸��� �f��;�֍�UZ��� 8�v�ͺa����� {w� �!��F:�O���ͺ0;�J`N�� �$��T+�`�����x0;�J`N�� �$�I�{���`=H�hUD�p�I0\�a;u������nΜ�Y����.equn��h��d�綴�磵I�Y�h�V��r�t���\e�9��gdባ:��MM��zɜjh݃��ݫi�s��qr��;5�o-i�ɖL��McVr���|v���$@��		�7S��ۃ^Mι*tQ��l`΋��P!�Õ���V���">��x��1��1J�_z���A+*�;[f�M͇���ss�N�rsո{FU]p�c��هa-�rJ�`�VZ���ŀ[�p��<�0ݞ���3~�Tr:�����L�I��I]���0$��$�ş�/�<�4k��2�F�����`wL�9%U:b�RL`n�?r��� ܅%�I���`��, ��ۀn��~ӣv&��X��%0	24�ڪJ�����vwFd������Vs���Z��E�6k�G�h^����紊s�v>���^8�����S �u�=;d�>�J�ʪ�^�{�ذ�/��`�]������y����T�����`RN��������AIki����7}|`�`����2ڥܺ���E��W{ތ6��U��0[������0��߶���e�ڰ�I�ҥU��O�I�с3#L	2��@z�uY��um���=��F��YQ{q�v�:�k�6�3���=���u�=;d�25�����Ż�`sc6D/�ND�ܴ�;ݺg�fɭ0[�����R�K�J��3�F�MO���7$���b�-ݸv�N��_��w���`zg`��.N+W�BR����j���&���\���w�t�7��X9�lj��>tS��zvII�O�l�� �u��αTئ�$�-j���l��5¸9��Ɍ���ƫgP�����_�P�(���K[NHqw���	7�0&di��H�ʿXl�� 9ղz6��ڭ��7�����Wa�n���kL	��{J�UK�\�O��W����W;���ަ>>��	�`N��`Jґ�*�e^}�����W�o��ٽс=#L�m���PO<�'�7�I�e��C�J��N�r�{�L��w��� wǽp�w wzm�Y$b%i����Ux�sPV2Oa��r�9���n����0�MJ�m��%0��, 曷 ��q`ݺ`����Un��KS �$�fF�'`�����UI/�[��lj��>�����ŀnN��RUw��� �7z����gP.s��W�p��{���ٯF��LBF�|�_'��~Xέ�ѷ$���m�zF�������>�����0��*~���d��/72��.Ͱ�Mٍs��>�Y2ŉ���P�c��I�wB�Z1��#�H��e�Ix�+:8-�ҩ�/q��	�m�K�(���z�;���X��բGurY$�O/v����v3s�=���u�f��M+$��tv�Y� ,��X.7��]�٨�ـ�`��u%��E^N� ���l:C��NJ�\�vJ�������u��{�<��G>���^��7.+���]���>8�^z׆v�78.$m��~�q��������\fF�����a���oKD���;}��{}�fF��U*J�������ذ�������&Ú=�Ȗ	ȞU�`}�g�l�0=:�L�4��í��SS���7m� �����'X�4�RJ�dz0&
_B����YU��fb`�1��#L��09�����b����6�T#��/�t�Ӹ'�6U���%�lu*����J��7<�IU��-�mZWP����n�ذ�L ������%���o���W��V'$#�t��~�u2
�O�@7d�=�s��X{��?�͜����rJ�ak�G{��3wz��24Ϫ�%Wrn����`�&w���[J���i��#L�F�}I*_U$�\��~���6��X�+���V�wq`�)��/ I>��F�}Ҿ����w�m!m;W<ex�26[��G��pvh���$g�1�w��Ey̜��	�����\�=�}>�i�wt��F��4��:�V��m��mX��n|��_|�����i��}�L�F��'l�v�w��}��ް?L�0?IfUR�U!�d/>��E	�DOj%����K�D l��y�P0"�6xR��x�%@=�6�ҵ=$qA�DS���j��"�u$�P�S͒.~%�P���Id��Q*$X't ���U �S�N������ )�*z�Q^���3�b����?.�n�ڴ�O�r��_�o�}���>i�wt��F�޵v�RZ�rBBZ�� ��俾T�.n�������������k�Ў�D{Y�5��-�'�ۖ�{�zJ�y��n��KZv�7$��Z�j���p����#Z��W�	��0Ef��U�Yyx��1�zt���0;{!��v��|�<���&��M�n07�i��Ѧ���L`�hZ�a�X��`y/���, ��o$�����B Db�H����S�w<�����]�gK���*�3 ��Ӧ0=$i��Ѧ�_%;p<� �i�Ӕco���Z�z��GWF�ݓi����]z��Y/�:����i��,�٘��W�����0=$i��Ѧ��n�vv�6ե��[�~ݍ=�Wd���z�?L�`~�Z���B��lp����� ;����&�{}p{�ŀ~��C�P��J۷�>�J��I�`ٽ`~�4�ꪻ�=p�ž��W��H��{� ����{w/�&��fd�j�R���`���tv6�nD�ƹ���I �[���9�N�N��,e�\cOc��E�ݸ1�5���e��*��!��=��jӧ�.��[mPzƬ�rM�m���[���D/fZ��hݳN1ᛨGj��L�j��+����6s�C��	�v9Ss�6֜�Ҳ�aϋ���<�d5nX��i�%�i���V�]nM�r[���h�o�m{���"1������JI�=DZNm�g�5×9�kݞ��<�v�����&��B��]��m����ذ��� ��Ӧ0oT�yg�Yj��0ޘ���� ��I��I/�JC�Ǜel���M���n�{���d�>����&M�xD�N�Z�t(��|�M���s��,��׀w��X��-�aV��VIz��$i��RU3�o�Mi�~�:��jI��E$,�en�5T�k���P�Ɋz׋p�+g8�PUܥ��˙�U����Ҙ�`�3��^�߾�,��_����jPv������J��R���UJ��ް&�i��N���L��_�����Z���z��$i�T���g&�I�0%˰:�;dv�%����X�w^������$�o��\ �u�м�a�p���S{�-��o��roX�4�>��NA�RB��lcV5-gm�twON�Sr�8C���]��Ph` 4������{l	�`�:�����*���ݛ�oDz����� � 7��`OH�{�[fF���+��z�6�-�������`ɺ���;�LwL`{z��Ye�努�W}�a��U�wv�&��&d��+��~X;�~�rJ��A���w�����nn������T�vs�_��fqV�v���2Ga���v�8��[x{xP� �@�<6`�=�u����zSN��w�`�w�'�i�=�-�3#L	rբ-�����m��w{�g�=�l�� ����UWa�.�е�
���Y�u079�l	�g�Wfɽ`nn��;ζ�ٴu�p,����w L���0�_RIv��WJ���$EO~OQU9���������,�P@��� ��n�����~ݛ�o{����iT�9�2F)H��@����Q�.��S��A�eb�(�`��7d:������ذ��{���_|�ː����;��UG,ljKV�})�;�LӦ0&���ߪ�]�EU��)YwX�0o^��i���׀�3��~�1�m��`���l�0;o�0'ti�!h��WH��-f^cl�0;nJ`N�� ��w�J��HT��}��3ww$ْx�8���@��:cu��:70ɗ��;m�Z�C<gj �Ԯ`�8x�x�����ep���Q���ʹY�C���B���vGv�w ��{v�`�v.�U�78���%� 9<s��;���U�<ഛk�#[�@������-��Vڸ�f���7:N-�Y+�ŋPy�Uۧ�E�ֽ��q��8	�s��|�{�G������S��<����% ��ڻkT�(۪w4(���0X6��[�j�ŠN����Ѧ��0&��y��[6��ӁdnW�o{����di��rS�D�(����/��`�:����|�UJ�g&�۾ŀ~�Ͱ�һ`'I-������&�S ���L`{z��Ye�努�Wy���})�N�Ӧ07������7`�֑J��nk�.{(�f3��z�nW\=�γq&����]���)Z�̦;�0N���#L�w^ ~����T��i� ���O��%�]�24���'t���դ�F�j��j�7����w^ o{� ���X�tl4	->�+��UJ�+�ٶ�$��鑦�#L�[el�:�N��^ w�ۀ{�>߼�}��03��l�Yo�guއJ1���EFxk�A�2Z��Pvg8燭����+l�H�A!�p��ŀzH���S ��u�\�.���TU�`zH�m����{q`�צUG,lp��y;�	'�}�����Y������
]ǩ��WmR�)$|����4��~���Ε�$�+��^ w�ۀo;��I`M���=ʎ��X]ٖfau���=����Y��yx�7�`�:;�~_Nx��)�l��� �>��smv���'o3��k�qSv��&�Y���t�f&��0&�J`�3���t�����x	->��'%X�w^ w��`Odi��H������2_K5v��]�;�]���$���F��J�ۺ�ݞ��7�6��T���"� �������$���J�i**���Y���w�^���Һ��U�zH�m�L��0'ti�˺��7?}������ƣ��������1�u��+��2�#�R�G,lp���nsv�fN�&dk�I/��֘Y�s��%m�W+���p�w�H�{�[�T�]���GWNs�xfauy������0&ܔ�;�cV���'JY-�`��$�|���`nsv�fN��*����0�6[_���� �M׀�v��������9$��>�5�AL���D��=<��e+�(Lx��N� �Q�����{��ǈ��`j�q`�x��|5�&�!2���Q�����"���6h&��70;������۽�����n�ڥy��)@�q	n;<��3��I�td����"��h����(���Cu�ӝ�X����+Ų��r�svK;�Y�MS�@u, �.�'H%9ۖ��ծ�B�;3���ɍ�:�f\pAŕ���;����,�Ga�f����c��"��� �N�'U*b�j�Fݺ��z�k/��흢ۣ��x:�vBjv�4� t�5:*Y�;�S1b�u
lu�v�w:F��l�y� ��n�Ӽ� �(��m��3��\�m<��؁�.��s��uu@�.���l��u]�n!U-pJgO0�t��)�:"�d���4GD %��rI�1����<�ocx��+8M[F�&�lU[w.�tm���>5��Ai^ݐ/$��͝Ɏq�9��^��F���eWmk�Qn�xmA�tj�@�l��)wp�!]Ym��ų���K���]G�[x+�5�;Η%j�Mf�:��r��v����x�SV��]J�;��� �:ƣ�����CiB{u[(nN)�h�u�Cl�6����r�+qh��8�F�hj��M�a��t1�]�N��@.��+��|��Z��J�XڥyB㭆Xے�X�ΣAɐ��wm�q��\�>wZ��K�sX΄&�����p�p�c�m5�$�<�mv2Q�SQ*ە��5g�ZU��FǑTɢ�8����R��6u�̻e%C0�ųr��ۚ�N��1�  
���3j�t���`8H6B�Lm��	�i;i-��k[8�M&i�ħU���sl�@UZE�E!c����+k���;*������R.���{s��OM*�F�k�V�;IQ�^^FWY٪U� .9Y�<�ͷ���NjW�#��X�CBT������J#�T8�!'mnq�˞Mɺ����+��mYGv[�"A�ų�4���Msg��m`�����{,�S@�9�}�q4J�dvL��7�`
;���C� E@�T�T���j!��@@y��'o���fm�3)�s.	Ҷ��)�l����!V��W[s<Ps7Fn�h��J�b����@�#�l�j�x��V�V�Vp�ԡ��ݝ�݁L�z\��%��ɵ���@vl�2���%��&�Q��%�SA���Q@l��.6tOJZ^���e�;qǦ%-�hW����HM���ᖸ8�n8�VI���hrb NSp���c���E��{��t�YWŴb��FaW�yC��Ⳟ'���<���Y{<�ScO�Wq���ԃ�=2u�3#L�F�$��Xnrm�=�*g���2C����,����7�������_/�l��zz�7J�6;L���`��x��n��� �:i�B�Ɯ%����ʯs�m�I7�	��|�*U~��Ɂ��+�C�P��E]� ;���7��0=$i�6�S��(��ح��*�{sЪۮy��x�5�j7�q����n�盱����|���>*�qX[H忀�v��=$i�6�S ����te����w7wg$�w���H�	@���I/ߕ$ٯ�m�{�z������U%l;�G�Ii�t�9*�=پx�����0=$i����ee���2�)��Ѧ�d�4��_�{w� ��B�AꤥL�Հ~��0=�4�������/�|J������;���]�N䞜��oA-�b�9ۇ0S�?����w���m�
�7�`g���̍|��l�f�T!���Z��w^��q`��L�wqg���������R��.�{l�Z`~��1qU��ERHH��UU:J��$i�'$�_�̔b˪��fb��LN�0=�4����K�\��y0>_r�~{�|s�y����#L��L�0=; ��MOU����Y$� Z�IEj	n^�+��pvh���:0��ڎ?��uV�|;e�䌵Wx��S{�LN�0=�4���Ɯ���
�k�9��,�����$i���K{J�ͼ�7�7���Y���L�`{�i�6�S{�ŀ~�Ͱ������ ���L	�Ҙ�`�\�K>�o�I_:��_�m8KV��� �{���n�����9���j(8�I��-g�����)},p�;���(�����r�4]ph�UݬW�TZʼ��F�� ��I��~a��y��پ���ⴶ�-X���J��=7Z`nsv�̍=U_$�<��=�[�$�;%0o�� ��ͥw$֘'t`�E�h9�O����V��}�n�`��0?�=�~X�l���U�&�VY^��i��*UU�=?��i�=�-����,H,DX�aX�AF*?�w�d�o��&��̷!.�&�a��[-/��&,:z{T�e������mUd�^�iӁ%d:�96�A�ۇiWa�hq��-�c�g{v���s�nݢ������z�������Yn�x�Fy��Q��G2]O���ю:닍�p�z����L��v��)S�f�[�.�8C��АJ���{n\�*e���юcl�:�۝؇{�w���SFGp��1��Z���wQk�@l����][<q���s5������h��خ��g��F�nJ`wti��b��ߝu�P���wq`ɺ���� ���~�]�Sn_�m8KV�rS��L��`zH��a�1wk�Ak*��`l��LXy7^�����V7��9j�=3�`|�����&sv��`n�;?�ǫ���M�7n&��L��+]�g*sm��,�(�úA"�˲��]��߾��m�L�0'ti�n��)��GK!� �MמI~G�$u}i.|��|��F���j��,��UXeyL�0'ti��#L	�%0	��\E�B��f&�0=$i�6�wF��)p��eee�
�u0?I`7;���kL	������i�6�:�؆A�Hk�ю�7[�����췪Y�I�ƕ�)E�o�UJ�����rS��L	�`zMŀ~Ӻc�H��MJ�x{�ş�]�&����������ْ���qZIc��{�ŀ~��XUW���U�I��$��=��Mi���bz륊@�Ud������{��S��L	�`܊D�a���Wx�nJ`wti�;�LI`o~~����Ǐ���q����i���.�N2�A�.��yv�V���?%2�D��h2����4����ے��ְ��+�S�ڰ�wj��)��P=��<��W�/��6s�[6��]v��U�s��ŀo&��;��,{�ŀ~�]"������Ձ����%\�?�����fF�e*U�J�EU��	�)")`,D��D��X��K7.~X�;�;P䊨�^�Ѧ�0=$i�6��U>�u�?��⭖6��0�湳[��q��-���Ak8{$��f��������t���#ޯ���0'�i�=�-�3#L	�lOYKbp��mX�w�M׀2u�鑧��UU�d��h�zW)]e�^&���`�cgF�dk �N��٪�8��+��v�24������*W���`K�Wkl/�U�e
Օy�	�`M��ۚ��n�������"1�6(�g'co�yO���=�PG��W$�<g�^l/`�
g�Ƭ�m��*��Jm�gM����`����l0�\�w/A�+Af�=P��pu��3�Bm
:�3��:�Gb��.�̣eMm��8]��ùr`� m2���ϭ�+�@�n)z����ʽ"�9����#�n�)��tEd9�O\+ �u=�l� ����+>��UAW�&<xW�y��&�k&Juճs��
եa�opGhx2�G�w����hN�����ͷ����0'�%�&ga����~��5��_����	�%� �M׀o{t�7�4��#LC���*��+1R���`d�����_RIR�7�i����[ ���U`�+��-X��L���ے�$i�6媔feں
���{Ό�4��T�nwv�7u��n��ժ��m0v�#w蛎8k��m�ӵv�;R��'Q��8�,���ݰ��;[e��t���m�L�4���n�,��ppf���q��W�wwqs� ���1DƎ-Q�D��0�EF� _uRU��W���٭0'�%��T�6k�M�l�C��(��X�o�$�3j��s�����������;}���.��F*J���L�n�$�`��0�^�7->�KV��S��0'vA��F�Ţ�t�jQ�t��mֵ�ŞS]�N8��ոo9z����]�l)|�N��;P䊩[d�W��֘3�`d���$�<Y�����.���wd$i�6�wwy$�8���֭��r�ݲ��֘ܒ��~�JT�I1/%Tb�#`Or�����(E"A�Nx�0�H�u� �$�xt%B^4b�} X,b�s�xJ��
a�Dآ���{G �MY *X��E`�`�����
0Hݺ1<��c`���)a��bAC�j��"f��HP�IeOrBZɠb��0*���D �D��J����)�aT�aE�X{����D��J��W��(��Q���~Q�>Q<Q�PNw�Ax
_�/ڕV_��t�06#� ��_��/��{�u0'�%�2H�ޝ��I��� �����U���*e��ݍ0=��02H������*����]�PJ�1�YA9lu0�K7A�(=�;,;�<:�6'�.#s����с�F��$���UK���`o��O�H:� �r���� �.J`t���0&�GX��������0=�Il�4�J��f�L	����;�;P䊩XԮW����/��w�`fn���#L-R\�{�K`e���VG,,�Yj�9��X��������@������F�z:V��"�fZ��\s�Q睺�k��\��d�@v��bMs�t�W7W��D�[��V�*�;���rl�I`ñb�o2�]+��w��S����]�wZ`fn���#X������2����,vd$i��rS�i論UYނ��|�a�U�kс7u���-���ŀs��m�u�4;L���ꤕ,����&����`�UG�? DuA��D��1X	��4`��g0��sm�,�wfA6�G#�\��AZ������HV��1�{>9��)��uƝ<pm��U�2K�\�ѶT�[�V���W���	�X�JD����cu�q� 1)�O0m;�\q�é#��[�$����;k�*�����X�%	���j��r�&J�;E�Ւ��=��f�YȒeA��n�gC��;����ϳ��gq�U;������;���)7b�{�Gu��\�� #� �5�G;n�%G�=����pP����x	���`d���;�*�a=��cm�t���rET�jW+����#`ꪫv8{�U]&4:����+ު����~*�r��e��6��74�����q߾RN�������{01���[ҵ,#nZ[%��ͷ�ۈ��|���6�wsm�~��|�X-D�_Ѩ��Q���˺�~m�/���߃�m��������ۈ��o�׶�d��,q_�$�v2''RAh3Ş)�̀l���/���rਸ਼	��c,���������|�柿6���F6��.�����ƶD9�2�a����m���vy�(xB,?I6�wz����ӳo�뻹#`�����l�Tu�4;Oߛown#m�u����%$����o���/ߛog^�7->P���/�_I���~m���+����������ۈ���wO��I"���+����{���o����~m�ݸ�m��]���m�J֦��؂�ڑ"�p��U�p��k��8�ֺ}�-�fq�������{�j7s�#�G����{�~_�6��ևww~�d��������`���ܛf��nL���n��ym��w���A̷3�����������?/߾�UK����/"e���v�m���o����ͷ������_}�|<��{��	�m�g�H3Uv
8�e�[��o�����~m���<~��{�q�m�������Q��Tr�6��74�����������?]���n��뻹#`����UU4۾�9w6�
�;���m�մ'$���=����;\�b|s���HqOlv+~�eU}���ꪪ�d�z��H�:��ݎ�6��\�TnZ|'	*1���7o���}�JH��f6��}�?~m�ݸ�m���t��D�T[���ߛl��Wm�~��{�q�m���To��U��ü�y�u0��UK�}�ၻ�4�=�:�C�O!�D"	Z�G>DV�ͷ� �[եt�m�i]�S �{���������06��U\�,9���U�ϲ�N�C���%w\hⱲ�c�e�ܵ��w��u��O'%-W~�ۻﱁ�#Lِ`wti�հ�(��n��-�7���sn���� 9�ۀk�Z��X����S ��`��F��T��U*�	>�����;�i+��C��7wq`���d� ��r�V+*�0�+��u0zN�6���z~3{�N��$����#H�~�㿶�\�k����\��Ѩ��l�u������8�,��,ť1e�T���&���x'@hgC�z^�۝�zڶVza�n�v�n���W\m[/OlwWkJG�r�UeF4���ŷ0V�9�;Ge�)Mb�(a��f��	LY����������r��Q��P���X�����xuϵA�D6W �`C3v��|�A��}J&_QG�/�O2i��<n�&+#E�PS�l���v͉S{�zu�=�����&CEĺ)E*+��������9ͺ`����ݸ����Udr��G)�{Ӱ�J���i�fn��$�K!�	��딲���, �7n��L�ۦ�DBК��E�[j`��`I;�;�ww�`K�L��GB�-�7v�s���	$i�nɌ��AՕ��Q���8��ul]��.�i�p�=�뇎6x�c-V[	����!UA��n��7wq`9�}����� ��zx�D���hw��$�8��;����`n���5�uA��T�J��ݸ���4��F�ӖL�]]�2�}�v�)+�ף3u��4���%�?.��w�#��9L��ŀn�i��rSI�`N�&~�WXXP������K�G6��u��ʜ�u��� ��bD]���W-+���ww�M���d5z�dŀEօɇ�u�]��&��wvp��#L	$i�&�}��g�v
8:�ex��b�9���'�	 ���& �s{ÒOy7^��k���!U�U�s���24���%���^������o7���31"�wF��%0&���n��?s���`������2�A���V�E(���GZ���nJl�y�ir�YJ.
��� *˼Lے�di��#X��� �úc�IQl����?�]���06Mi��rK]�Qr�}�e�����V��ذ�w��� �n��u=z�q���T��`|���06N�����RI.R�������q`����S�v�m� ���`M���0����>=�Q�!��A�����t��l�ú]yb���<҅��n�'r8��[����F��4�ɑ��/�'t`m孾�E���̼L	�4��Ѧ�`��,{Z�KPAʰ�`L������٭077Z`e��]Lq�J&�	*�7��`��,l�0:ti��:�uw�˲�yx0:ti�6F�:4���V�'<���P�5"�w� 0�����¦���F!<QΠ|D��>g�=q��0Z)<�a`��X��a��u"��!��}|C�H2x�(8.p�I��%HP%�?#����,�SCD�X�  @�F(��!V����要����T M��巽ݺ�V�mR���� �qtϴ�u�a-��Q5W�2Te.N8�~�۽V\���M�׮��^� `���}�lv��v��b6�I�1�l���l)�-E+��@���e�۷q&�N��*m�q�n�5�S���s�����g�U��<Dv��]�ƥ��=f2�Ӄ��6�ز
M:�۰e�K-�'JA��� �KSr�ZMh9�X.�j�) Z'�#O/]�s�C����mT���*��|�7f���&��mв2e8��F��%�Fe	Ҏ|H�Ͷ���n������EV ��1�6��N�Tt�cv����عn�Ӑ�Nŗ8���ƶS�nv�b�sk;S���%Β���"�K\�$� |�Z���z�x;b6Hy����~^>#�C�㦅l:p�mmT����E�v` ��,��p�m�Ü��l��q�Y09���B]:��Mnݣ���s�㝞$�@;��nf�r��v�e! �Wf*�@vW��[q��A��ʪ�7�GE;I�<��M�:;V3�lU��e������M)g��j�	E�Ӵ��p�)T��69���q�hY�
V=�,�r���ں��;A�g$���eb�}r񃍴�0r�qcm���#IN�oTƤr��쎷,�Z�r��n�J�6b�ܼ�ͷ�,�x�"D���:�����J\�v[{rp�/N�&�1HKj��7f	By�s����!�=�x-I�����e٨rޮ����WWT�Q���"���*�hn��Y]��=�]^�K���ౠ9������q���{-˻���L�UVmƮuQ�h��&�V��*l�b%%���Wgʭ��\�v՚�+�"Zk1�yGm�;c�Ӛ��jx�"�вn��3�n���[&��%�z�j�,��uv��v�5O*���'m�qm9&:�7=�1�t٬��'X*�l����w��eyc��셻*�V3��m��v�� ��
"h'��O�����S@�~�>Z�I��;H:ۍ;�g$u:L5��i,�-:H'����r�)���K�\�d����{�v/Y\��W<1�n$���F+�;t1��`K��Ax�M�S��sq��d	RH���]�ְq��j73���~rq�� �G���ы3���R���i	�ܕ�lT�8�s��0W�C��4I�:�Ѥ���e�k����=��,M��! ���/���F?��Kep����y#`�^��g[
���m�( VC.��lu���|�J��ٟ:�$�vGeZ���XN�0'vA�ӣL��R�*�U#��]���02di�)RUWf��f��o7qg�K�l�#�!�}"��-�S3�m�����%IU߳u��kX_4q�Uv
8:����� ��`~�a�Uy��l��o.�V"�X
�]^l�0=:4�ݾ��w��`κ���PW�U-B�t�յvn1ĵn��poq'��6�)��,#���1��x�|�v�S���ۦ���]V9[��h��`�2[�JJ�T����%T�;����L��ş��l�M��G%E�5+����Lލ0:ti��})����Wxw�9�/����L5}T�%\ٿy07��i��})�ӣL	R��U�]"���eef&N�0=/�0:ti��Ѧm������\����'v�Eɶ�z���j^Ԫ�IF�p`r�n݅ݎ����^K��;ަ�̖����=���T�~���ذ�xq�ʻ[^����&Mi�3u��̖���E�w����\���L�F��gj��,�E���f"+��m0��7��xw�� ���׵8���T8�L>�IR�����ɶ����=��_u�BV�(�$r�����?�����N�4�푦qh��~��uJ��]�z�=��>^ɜ���q�n^�z�We�g�I�Q������N�;Q�(ԮW�w}� ���oF��Ҙ�u�?e����YeXy�ş�|�=��,���o;��z�^�\hed���X��̖ϕU]�Mi�2kL��6�H���[V����]��=��,=���\BB�T��ݹ�02�G�W`���e����,�{�����`�w^ ou�j�T?�e$m�ܠ��D]Om����2t#���ӐY;vtWT�4:ʬUAEk�`�w���`z_J`M���uJT�vU���Er���������o&�rkL�F����k�uZ�nҍ�$� ����ƙ�J�]̚�rkL	�D�G/��e�J�)�7�Lލ0=:4�����?.(�o�I*n;]��wq`�`z_J`{fA��`�t��U�5q�xyݍ�V����-��i!���8~w�b���+��5�$�M�;O�\�fG�뫋ۆ�iSuB�8P�A�6��A������\C�NݯK�T�8�8%�@�i������UN�j���%Tv�v̝�rk���-�&���5�/U�����n�n�"��vz���.�r��m�ΣZ۳7kbބvIK������TM�yi�t��s]]�쨻=�c�ڸy��<�;q�n�&����V8���� �]���?>�������̃��Lm�pY0R(�C��V�gu������owذw��?�6u�Ì^U�)"j�[^���`v�i��Ѧ���u�K1e�⬢Օx0;z4������� ��t�?v6��RKF�r�{�LK�Lt�0;z4�շR�m�}�R]3�­:닑ru8�TN��Cֹ���~�,Oe�����ݝ�~��07z4�����#L	����2�i72S6��I=����?���P	~�Ki6l��l�03Ӱ`yr��?V,Ww������Ѧ�F��n�9�ŀu�zk�ƇX�U�f&�F�� ����gF��!uCh�Qڤ�ڰ�n�9�����L�`�W
�ʻ�ԱY�=zrR�.��-�C�c�����pk�x�tr��U����Cv�9�� ��q`��/���_��Ъ�:�ȳ*�06ti��#Lِ`n��_X��N&��U9V����;ͻ90@>`��`�FH�0�K�����%�����i��Ѧ��X�r�mhNU�w�t�7���ou��0=$N�Yw�˲�yx07di���L�`ṽoKv���Sۣf���.zК1��OB:���8��Z�����@��M�~uU$�p-�`�Ƙ�4���0:��J���T�]�˺�L�`ṽvF���,���E"���Հw��0=�3n�f����i�됾X�K틜坰��F*�W���03f����i�䒬*���R��/ߛ��g2��*��Y�U�s{��sw���ޑ���� m���;��͚���ut$�ڶ�䞜ݸ�vŨf�6�n��^��̒�GqD�B�qʿ��ذ�l�4��Ѧ��X�*�0�T���d�4��Ѧ�0=$N�Yw��WJ�/�06tŇ�}ｋ ����?-Dٿ8��Tܣ2�06ti��#Lِ`n�����\�:Udv���ŀw�`���i�鑦_����$U$�T�H�ER"� ��v�w.kHZ0��8딻X�/8s�CE�s���mʇ4�:�&�;N�ȥF3�W��[{F�,ȋk�A+�n�!t[��N�Y�Ż<��mrvtm�Xu�Um���c۰��[��ܥڞŦM�<gva 6��etn�[��^���qkn{"�3n8邁Y�{i�\\��/ 7d��-�x8$�u�ƺ����&6�]u���<z�����fe6��p ?�ܾ[s�ۆ����sOc>¯0F�-n^�+������n9�vy�T$R�
�T-�r�[-^����vF�:4�ݑ���*�S
3�ݬ����4��Ѧ�0?l���hzʚ��[��*�;��&�0=/�07di�*�-\���`������s�|�sw�_$���� 惡�iHWi4䩁�})���w�yx	���4���]�Q8ފ�!
6�Ukv�ȕ�]M��Ҧ�-��1WXh7n���m����v�
�+�wLX�y�ob�^�0;�E�GRJ��7j�;��,߿|%�����!�E[�U�^I/���`I̖�������ͽ�r�4�9U�ڰw�ŀ~��x�F��`z��ɂ�.�.����Sw�Lލ0=�4������I��׀s��X��䷧�^{�`z_J`�uQݪ��9��h<;�]	�L�$���4�n��x����A8��*jʭn+\� �;�������Sw�LWP�Z%���+ ���������Sw�Lލ?���M���=U�vƄ�%X=7גO}��9>�4�y��BzTz�uB��!��X��d%X�cH���=7�B!�\\\Ɨ��J�%�H�!Rs�#.OՅ4A��rsTHY�0Gǅ�U���z���3
7G�B7���Ec��"X��H`! �@�)�~D�c�@8)ĕ^ �3�2��C�� E��
0"E�I(Z�B-���C���A�C�4�hŐ��SU D�2������xhA���Z�r��`�ЈT �E�X1�T}]qj$&:��=''�4����xE�>aeI�`��B,�@�-XB� �w	}�m��>+�E�Iߨzp�TX�� O��p�wD�����Q���� ��O�S��X�/ߵ$���i��Ѧ���b/�Gy��;}��%T��&�L	�Z`~��,����7�j���%M�Հg�4��%IR�n�_���m�=�07�w]c��F�U,�K] �F�L�+��.9�n�����G�Ęu�ͨNe����������Sw�_����0=؅��p�X�Uʰ�;� �;`g�4���{I|�RJ����s�/�n�W�#������~i������k �����`�5eV��U�g�4���`~��l1$�*(���!��_'��ӒO�����e�����S��i��UT�{{6��=� �;��uA�'�v����Q��g�bȥ<��y�]�9@����;O#Ʋ�FeQ��tQw���})��ѦwLX�n��?ouc�$��F�r�����UT��5��u��̖�T�g����RJ�(YV��b�?l�0=/�07z4���.�e]*��Wy��S��i��s%�=�0ڪT���|���q`����5!,r*�LK�Lލ0;�4�ݑ�_��a b�RP�@s�����ɛs<��'/k���F�nz�[-e�k/A=ە����q�q�i:�t��y+u�V;dKK���v�� ���e�u���uo>Ź�p�;t�qAl�����&�z�0���
���P�`��[Xź�WIh���v�^��:�F-�d��/9+(�m�6��]�������dҥ��q�r�jpSn�y�����A���9ù��������3�nYZYrnm&�.vڻA���78۫+W���&x\�������*�YE�L���0;�4�ݑ���׀w��[�ʢ�Ҏ+\� ����%UWff�Lo7m��H���6�ibnX�`�`��,�ۦ��|�{�b�;��,�:��Z�]��J��0;fA�;�L�a��_�}�~X=�X�A	*,�D��{���ݑ�l�07fA��&X_눺�El�ǳn�^��ɮ(��v�(rj����g����ʛqT�r��X7�� 푦l�06ti�Ժ��e]*�&f��wNI>���Ψ�X�'P�	���'��|��9$��q`��,��Z��MHK�eXl�06ti��#L�`�.�Q�+�YAU�0:ti��#L�1`��0l���v�IiG�U�{�4�ڭ�/�fot`OH�=��[���̒�F�J*�Wn.MIV���7�:Ny2��w/p	vC�Ł���7~��O�`ñl�07di����ZZ�]���%X9�Ly�� �7q`��,�I6s������4K�9$����9$���� #���-P�*�I+IR��G��d��2�EuX���/�vF��4�ݙy�� :.��Z�MВ�KV3#LK3^��77z���i��W��\v�v��gm�7�!cgq�WmKځr�ۂ���.�����瘎9s �70=.J`d�wF��4���1j-��*��L �n���ŀo{���7^y6y���ߩr����0$�4��Ѧ��Ll���}b٣�r����{�ŀ~ٺ�I;�{��*��(@��G�!���n���;��6�֝-�	*�?NIl�UU�s������L	�`g���n���Jނ���hӛ<dȜ���d��We�&�*ڍ�!]�9n���^S �&0;�4��Ѧ��L�5F�uG*%	j�;��,{�ŀ~ٺ���,�ɰ�����GBKxs�L�7��v��+��֘Mk �D.���Ԅ����`�n��0324�RJ�y&�r���~�*�r�y�� �[����{��$���I 	"����gr�ƛ��;n�-h�v6��BOF����b�Ue���Ӆ�#�mO=�R3�����e�0֦�<C�ɸ�ev���r����E�U㙸eۛ5�;ӿ��> ��k%ȻHT�8�Z�T�b��֞==�ɞ�ϢA���pWA�*�\�J�S`5vz��vK�f������s/q\r�iB����a��l{{Z�q�l��n��E>AS�}TW�}�M�3M-�4٘smb��X�n�h�9V�D<0B�=���E[E\tpuX�����ʰ�}� ����?l��_$�0�}�X�פ�/���/Wt���L	�4���qg�6w�_���:[Wl�9���3�I$��I�06��0?L��!%U�"�����,����5��0�7^�t,���IQ(KS3#L��I������������z���U�=�g��-=��\�v��|t���N��D{�N���K�Ff͉�+�[���`wti�6к���R��Y�~ٺ�I_��� *!!V��R(Ȑ
R�Dk
���b��x�������Lt�0=]���
/Ď�e� ���,�����$���Oy���8�V)%e$ �L�0=]���%0=�`yWP�F��)�e�`�{� ��u���L�05it����U"��x�uUθ��'S�eD3�����Z痶�f��D���?\ym,i���t�������ۻ���Ѧ�%�=:'Y�,�ŕj�^U�0$��oF����������Y�7Q%RU,� �;��{�����J^��p:
����K���~�x���b����dQ�ɗ�Y��*IlK�L	$i��_�N���v!j�u��%��-� ����	$i��Ѧ�%�t��^e�_����NF�x���&g���y�Ƈ�4����ι��,�����p������\����i��Ѧ�%�=; ��J�V��)%u�;V�wqg��/�_6���9�0n�,�}b���GP�Φ�'X�����U�n�L	&��w��m����D�[���￾��U����	��4�����HT�)	D�`*~�EO����o$�{��.�.�eZ�W�yL�4���� �0�7^��7蚣���aU�v���]��Џk�Ƒ��z�]��-��]��yx��`�c�䯕U%�I/p'�|� �_Z��;��_l�y��&�&0=.J`l��wF������R�$�ۀ~ٺ�n�&wF�t���U���~.�++����iRUW���0$�� ̓�>I���x_���Z���!j�;�ƘUU.I���6���i���UIQ_��QQ_�ATTW�dTTV�����*���Ȫ*+�EEE�E_���E�A�E�@E�PE�P�����QQ_��QQ_�EEE"���U�EE���TTW�QQ\��TTW��QQ_�U�U���d�MfI�?Cf�A@��̟\��� _@      (;�        @ x}  %R��P($
�      � 
 $
  	�A T @  AED,   �  (   ��� S篕��o)��������y��g� Δ��/T��������������J��K�;����RX�
`z�w)bޚ����7��VM)��K'�g�ͧ�9h��-*> w�( ( R� tު}޷y��:��ɮ��� �VYU��ӫ�����}N����z�J���@�Ƅ��uT+ V�w;�DŕOs�Ү�uJ���� =beJ�Ƥ,mU$e�T� �  �   �0 	�*���ܩ)�n� ( �{�   : 
 
 �8 =     �)D�wT�VZ�H�ҡ`:�_[w�>����� ^Zz��Ϋ� =z\f���g����ͧ�� uO����n���k{��Oq���� J �EPIC ��+�]+q�Uv�Ҭ\v�>�w�=�w֗}n�Z����ɥ^ ���n;}y�ﳯ����gOW�5����JY��7ԧ��/��:.�z
xf ����z���{����}� ��(( %A��������y���u����V�ε� �L�t����Y_Z�ҽϠnzz�/�S�g^ �����z�ۀ���\���.�;œ����jW ��>�7��{\����-��]٫�5M�T��!����T��56T���!����S��J��G�4�تT4RP O�$d��  h �!IH� ��'�����	����?�?�����+����G��c����TW�����DTWj(*� �+�DTW�����"����������BI�,8�3�$L ;�{�?���9�۞�lכ��/3�5��6��n5�y��c1��4���#4^sY��ٍ�{`��8�!��	���I�s[3�0f��/0�>4i�K��@c�`IJc�6��߼"��8i�8�ɉ���i�|;$@�<��~~5Ǚ�o;(= k�޷�A�0�%�#$���_>݁XY��|���^LƳ�m�l��I��|Ǒ��{����'�JI�3��|��ag"A�Q�j�W[��ʉ��1�B|+|�=��#p'l��W��ʜ��"���;�);�rpl���cj7�x��s~�5������|����c'dA:XL0#F�4�2�8h��5����5�Y�{�ޑ�z���z2A��=5����zo���;e$�d�pьf$��8��	1t;p��vzxg���M�p�=�ƏB�lu�������	�A���@`�΀���A�����<1X��pѰ8��H`�cz�b�V��v�&:I\%1I%�����!���aC�� �I8��s#��qI�(�=4�����i<��������5�}�q�u�'4���:�kcf�B;I�	��,��0���q���n��A��~󮠒~CAi(�$��E�wU:���ֶF�o4o�H����H�#e����Il���}����+�1��`��.##@���#sF�ڲ��e8h60���,��"ʒb�b�[Rj4��%qM)�ė�fI 4)8����A�xlBV�dŀ�%�$F�� �Hlx�����ËN!&	.*��I��ڐ.) BH$.�Rt��ɏ(�T�CH����!
`�5*D8&�f�L]�58RpӴ��&��sH���x㭛�$�;B2�0�m&C��a�g����<��	 Ã8a�<���ͯh�a����\cG��tU�$h�����$f�a������a�`�t�b���᱌ѽ� �4�83���#)YXӰ�o�M��Hlx$8:v�����C�Ӂ��d�NÉ�
|,8l8��KfaD$�b�B�;X0��,c8�`�$��,b���ma��b6�y���>7$<	+EZ_XĲs�o �>ӯ��,�2`�1#����;''���6ˉ��1Hp̎L2��ӆ�d#�L�'@bH�+��'Q�F�Ѱ�F61:Ꮇ��N&�����a��	,!0'g�g�N!��I���!�1� ah̵���C��i���l�d�5�E�3-le"qd�XhČl��0ƒD�@NiٙI�ܩ�!��T�B�����\9S��rR�P�8 e>q;���.����V�EN԰�cq1cTc+�x|��_x.EE.]��:��N��2I��m"��Y|G8�}��/�K����>V�g��� �8g��g����l/s����l�GYrt�W~��yn%�qRI�.�YJ:�WB��Kn��c��{�;'�R�ޕ�I�c�]qok�+8���C�R�ZpS���6w����i-�u�E��i�ȉJ5�U.�[��ۺ��wZ�%6���~��*x(�$�{��u��w�s�^S�W*T1�1B(�����u7vV�R���_��_}Eȫ�Z�Ⅹ|��֧V��	���Z�_s�k���d<I\T��o�Fky�Y��.Nfp���v6h��Ca�kf�����C�'c�-a�3N�6!�|RLuQ��b�Z�� �|4Ǟ�W��}�E&i� �v	VX��^ b��+���� �1B�FVd� ��l�c��w A�ap	3��QD`h�'"�A�JAbp��a�<R0Ѿ2�&��y8��8N&�pYE�X���Xv��3, ս$�3#N�3Z�Z�1�0	8�#9�[�D��ް��y�5��#�	��Xo�UFK7���tx�pѸ�� �����o3'(�0t���Z�2��Lf��0�Q��vV�@@a�u�p�a��da��I���c��0#q����`A��q��*04�:6��v<I����y�<7���u�����J�0��1лN"Fos���dɣ	���a�07&K�B"b����:���1 ă,��FH&bD� ���H�K8��f��N�d���9A1Q�͞��z�Y{���ٝT�7>fϬ�Zl�sZ3
ѧ2tl-ְ���C�1"4�� �O��"&$����#�'�e�[�Yh�(��QV�1����&���"̴o�$&x�i��jr��c�����N!�2�1H��x�+	�H1���C�$�_W���F�ѳ|�KѰ��Y���6Ύ2��4p�4h�m# ,�����t���p�����rjgA��L8`Fa$��CHJ��)6�0Ɉ��tq6�B"o@o>3#�:x���$�6ּ�H�������I��ȭlHn^Yp�= ����Œ3{���J%�n+Ă 秌kd�<�g|�#A)��sW�����2��a<R1�&ė��FFx���ё�0�Bc������v�� ���	ѹ�0{e��8�7�����:5��i*qК����,4i�6���h#4f��o�bI?q ���|R0ӂI�:��$�a��X�G+����F��0v���"�	sV�Z9�y��f�њ��# ���Pfi�4�$�b` �e�! ��ы@�),$.8�0։��k
��66i�o6f�F��'Dh���1�
SN;wͫ��3�q�Vs���&	!>3� k�bO% �\ !)�`��t���		��F����f�s�<���m'A!�)�x0�h1X0IaC��$�dӴ!�&L	�14�HLEpT��R�0G@�XG�0RFC�p�zt��ך��s\!٭���a�p���A�цBF!P咪)2�ff�ur�
_�R��"�f�ߙ\�##F�X�a���� �[Ϲ�"כ���{�:������ɂ�A��K8�L��t�1I���c��h<q�� �k���A�H#YųX[4q[�`�K8�p!�,�}�>���^�|E͞2c���A��A	lVad�e�&�d0!��`�	!��+J���,������w���_���,���"�����u!�l��}�*��f�8����IΤł�� ���c,I���HK���K8�6@�h�pY�{�����u����~~ �  -�Gm�       H ��|�  }$�N��n|<@;��9�W�6�Ͷ��T�&       H ZӠm� 6�-66��z��m��i��ÒI�I�n݄����=� m���m �� �m  8p�d$^�l�v�` �	   m�  	 ���  H �k� 	  R��@9�-���eicm5[z�*8 ��k�Ft�*�dZ���d�Z��  -���l��WT�wRJbn�m���5t&��<H �  $ �m� ���[4�J Ѷ��ڶ���l-H۶V�	  ��`۶���۰�@m�A�D��[m����R�&����(6� v����]5U�Nֲ�$  � �X­Ul���Y���:m��]J�MT�5�\��.{t��{n�*N�Pu@�-���Y��m�j��V�r�v�YW)UW����"� �U'j�����/���/V�U� �:ۤ�#P�t5s�r�;t3�,ݧ�k�gi�΋��1a[�k���ի5&�D�$��e1��9�pX�8^�[��3��q��*��F���)�\ڎX.G;K]۶�ۓ��mDpqX�ݞ��ۢ��UN��]�����ݶ���(��U�H�d+����UU�vl�;v��ͧ5F�C��,���aKsq	��ĈHL�)��i��b��M�m��$�[]�o�jC�6ؑ ܝ>���  8�$[@p ��@`+�i�cW5*ԫ	� m�h$[@[Am �[@  m:�m�F �	�Ԛ��p9����[R C];h@���R�*�.Ҭ�U@8 m���m���cm�ml�f� �b�m	e dz�[M���.À�p ]�-ϥ��$��mu��h����^W�j��j����=Am]m*�U*��pi�t�{�ݶ�m�%-��  sn�n�ܭm��   6Y��i�[AmKh@-�� }}��#l�L��	��m -6N��@  ��5][WJ�J�+��v�魸� d�����  Hm����$H�e��ޡ!�� m��m�iRbY��ظ�9�`)�!ݲ�owm�d� Htj[f�e���F��� ��}X�.�j`������cm��	ۙ[.�eYP�-�$rC�2sm'm��m����P	e H�����H�$[%6�[4���۳ 8[@ �`[[lm����hp[d  6�m���n��m��� �` [Ri��֝'l��l H	  /N09n�s� �	l �H   ����  6�  � m� -� ��n�8  $�kd��$@p�� m�  H����Ē ��m�8 �m�    �ۀ�m�   ү`�Ͷr�:  ���� m���H�h rM� ���h� 8  �`$6�m�   �� -��r۶�8=�����H     l  6�    @7!e�-�`��� ��� -�l�  8  ��]6�  qm��   �@l      �       �� 8   � �	t̀[@ [[l,��m��� �a��-�$    -�m��@ �N�u�\�&:�(�j�V�.�l ���m&  �[@  z��k��(�#� ���m��᜼��9:4P�u��L��m�`Il�$9��k�lm���$�  �� ��m�#m�I�%m�Y��V��@�ۀ�6�@��E��I� ��6Z��V���X�� �q�٭Y�ۥ�:�� e�@ �#Y�l z�H� t�YaV;`��)j��(�umJK�A�S+g��` �M��m����n�������~M�m'6�-�H�:	�YnC � F� ��Iiu�����nSd���`�l��-�6�� p[@ ��Ӷ�6 �cZ�l�lYA��p����� *ۢ���m�j4��uUK*��Uu7m�h -5�� ��� �].$� �i m�lm& ձs�5�8km�� -��-�m��qm Ӏ	lm[�L�݂@8��9m�I�m� m�M���rmm8��Hk՛l�E�a�ojt� � �;M����i&a(�WOj��Gi��i]���˳<�I����+�-��K���m�����r@�ڃ�֤�g-�;]�/X�f���l�� ,�� �u�mZM��c�-�m& ������(!�ջPl+���m�-�m��v ����C`6�nHI��l ���@4R� o��6�y��	mq�m��Q��k5D� H�`�-ݪl�礞����(����v�vW@)�"n���[] q'�� �\��4r@  ۲B�$�$�"��p�`�����N�[� #j� ����֭����'@ g$  �h8H�n��[E���  �I�l�m H   ������ ���o6�:�(m��I�@l^����M� v�o�$� ��rڷ�-� 	C���-�&�m�j�L@-�m���;e�&�  �f���mm��B@  +k�9�  ��Z�&����w1��[� b�EK��!��6ъ�����1,s�3nya!�K��
T8jI�([v��%�������p88  ��-�� ,5�իE*��]���U�
���� �ւ��d�� -� �g����UUUQ<��� �l�4�@�`4V�p !��m�Y��f[��m  ��Xհ-��M��mD��․�����6�tRY�s[I��ƓIRl��[% I�l�S,�@�����{��@8[x��m �M�o�l6�@�G �6�R�ʵV��2��muV�e ��Ā��mUPl m@p�ְ -�� �gm  ݶ��lAm  ll-�&���%�  �'@�rXn���\ 	    H t�HHΛ]&�c� ]6 kn   	  -�   �  8� `� �ª�
��U�WFU�'� 8�XKɭ�lm-@���[j����n�	/m��z�8��m�#���m�  -�� � �  Vā!m6[m6�  m��m� [V�~8x�m� �M�  �i;GJ`�h [@-3l  9��   H  k�k	Y���ӆ� ��    $�@�  �  ��    p� 	   � �� �H  8  ��m��m���@��j�	��T� *�^R5���   $@�hl[x -�H[G HM�k�l��sY*.�  $ ��M�sn�Y�� �mm�ml[�  y�D� �h�H[B�"@��k�i� �ҭ.�V�� ��UW@<��  �`    �lm�         -��� ��Ͷ-� �� �  p8 ���  jF�<    � i0m�i�ŵ �v� [4�6�` ���[�l 6��6�-��� q��kn-�-��`q�ٛR�� �h
�m�h�"�݀ 	 �  �J   $   h H     ���#��   6�m�m�� �    ��@    �`` m�����+U]*թyۙ�s��[E���u� �@ kt]f�p4�[V�p ���m�� �5l8-��p  -�R�l����+��,�9j���ڀ�+8m�m��u̓�Z��ic��S"��҅���V�bq=���    ZYчA�̫UUR��q��kA�1�N��v[�����Nmnx�<=�$��Wi)�9$X��o-�����yR mm�66KN� >��  ����l	n�N��u��	�V�U���ql0S�][u��oz�o{��"���?�􇾇��?�y������)���������ʎ�]*y�v��MI�0��AO@S�"�uzq8���Q}C@�6�b��z��
�mO6*#�H x��4�A�mN��Q����<:#�x
m5&�Φ�K� u�\}|�u��ꧠ � ��"��^���9��Ee�S��@Q�O�p��- �i4�芎"�}U4�t x\4(���0?��DMPM �(����%�
b&����t	�pA9�x*��E �p�ޢ�zu}j�����%���G����M\t"���H:���P>|_���G` D��T _�__�	<��@� x�� 	�G��P��Pt�P8"��|��!��?hEQ�� Rq��sJ�l���	�� h4�/8�P�W�'��D�נ�"� &������@E}��Lda�o{�ww����?����B��TUt�\��;t�m� H6O�8�P"�ݔU[����ZJ�߶�thI��2��=CxV�ga�L06�9yb�R��b���] #c�݇�i��j��s�*݁y��'�d^�\sP��6����M���zi����ų5����î��Ak9�`9lG<�0uqPW4��UCӖ�	�T�r���x�֪*�<�Y&%��������2A[��=���s�A�=�6�2�t�N���a�Al�Q����e��nC��q��@l��:�I�Q��t��ӁY�K�U�Z��SZ�i%mm@]��Ítd�ڝS�fv���:���ڹ�W�n�H�i)V
�Z�^RU步Z��a��p�vK���v�(A�����x�9:ν�v[
}\�ͮ,��P��c�􀳹�(��bj��t�>zy�->}��k�9��y$C<����P�N�J�{���T�v�+X�f.�,�G-�rj�rg]��My-ڳJS�pm4����{Lݭ�l=q��}� ��:��]����%��mn�l��AWm,e:g<�t�]����jx�ɖ�h��T�ó:]�5�a���*�#Jl�e��B�Ԧ�Z'�E\�I�ѩc����sjm���
V�uUG<'�5�m�t*�ܮ��n�J�t�\����wjޑ���K�^�kJ(��M�7��&�AJX�z�%w*�V�8iP*�'N��6�P��c�XA�<��T�͉ٻ:���
=�V!(mL�qy]�j�r����k�� ̰(J�񀭱�U�٠[t���'��ŉ��	��z�,ױ�Žl`m��$q�[#p9��K�#<�Y� �e#�s��t�4�z�l��!�˵�Z�[d��Kh�G=�������&�C��$3�95���i�N��JH��%X,���&Nm�����y�m���A�ӑ���[DT��*hҎ���CB���x*��/����D>_��^"E�s,O������pg��s��:e���-�ٔ�J�U��3�F���\f۰;�.Ɓ���i��ٞ�v�۔pk���k!;�B��e�[�6��d���M[�ۣ�1[�A�sӓvݴE�o.�����Ѣ]M�Ko).]��ZG����nv��HA86�3�
T�.� p 6+���Jv"k�蠦X{fݠ:#�e�{��ۻ�8�����N��ߖ��E�f��'' �Wrgr���M�÷�d|�wc"��&{��U̚X�J�w;�_�������=��V|{ͫ��$��pj8X�۫�i�kSi6����V��E��������:r���8��76���bǰ@>qR�m�0�6�t��7ww6��K@8��*A���~�_,ݗV��#g�]\�W)��p�߄G qR�Ih����(��T�h�\5���;tnT���m�tp�s�;n��C�x�r��[}��� qR�Ih� N�7n�&"�R"iX�V�m�����N��HbP��G�(u�_DV?Uzgz�=����짘J����IB��3�uXܚY�,�����l�`s�["i�J�n+{��꫱�>T����@>�-�I�j���'I���`wsn��U�Un)���{��������z�R�Q�����#mf�lv.�QD-oQ��;��0n��ӛ7Q��NQ"����`f��X׺�ܚXܚX݉�JT�u!&����Ih���HT��M�2dv��b�j��]JBj��������
�� ��! {���o%�������nՁ�N�Xl��萔�M�D�p�;�4�3��Vu���KWul�)"Q7%
h�}"�������?^�ܗq(����N��-�:uC5,Wm)`�'i��1w{��],a�\�w�H�%�'d�����U`s�["i�J�n+z�U��H�l�`fl�`g^�;Y���QD�ȕD�;�4�;ܚY�U�}M�?yX��+7j#hu H��)��`~�+K�nl��V��5
��i���C`*�x'� �<��煁�z$k�)RA�T���s]�9��T����{*����r6N�Y��mq�x�V�䮣��[�P;��1�҄�W��ą�5?��۫�D:qǀ~��� �����^���}���3*�%7dQ(�,�mՁ�ɥ�Ź�����ʠ��q
H�M�IBr�	�`���1��- ��HyS3i&�)IJ$Br������`o^j�3��V�6���ZKtR�d�:q��v9h�~��}��9��9���]v���Q6!4�r�Q�H.6q Qۗ���7Z��gn#%[��{*Hd�T�rG��4���z�t��)�C\Ơ�����N�k��8���Q"�l>ۥi�����Wj��1Q1�j�I=쫧����x:Q����usۣ�}��ƻ\�����֛y��̕	��9��%أ[.Zv���c��jF�tr ��Q��V�;Z5�z����wu�{ݽ��}��\Nf�1!)Ӹ�ہ�j�����fwGm�v�	�q;	�%ʈ��*H�N,��]X�۫�s_>� ��U���%�:�$RS��p�'8��bv9h�*@ze���I�$N'*����`o^j�3�4�9ܚX�ͦ���ۧp�t��9����T��=���s؜�ʔ�M�
E`gri`s�4�8���u����<�j�JFܕ�hs���;\�h�lkԍa��x�٠�r�ڶ���q
H�M)RP���������9ך��6���:���jR��	2�l�^g������H�f$ `�

���'��@s��7rx�7��V:�R�d��l��@N�-��	�*@z�k�9Y���Q8�I��a��噷��o���bݎZ��(��	��8�,�mՁ��o� �=�3�4�5i��u"R�����m\=t��u���}�,�W%�tF4<g���v�5�� �D���X[��ܚXܚX��V�3i���]�N�1ӎ>����&�A��Ł��j���6��{JBSq:��J';�K76�0Tz"��U� O39����K��Sq
H�m����㊐�� {�@{��d����)N�I9V���K;�K;�u`v�shQ�q� (�c�A�r����=��F+�E-r���c;7*���
�%8�Q9RSR;��K;�K{�K�s]���j�Q�*H��}���I��\X������i4�=�Kht�D���N9ٳŁ�{���������X݉�JT�NT�M+m��Q�]�`omq`}���^�SӋ���#�����xr��$����RՊ�FƤ\}�Ł�=��o��Vu�7	��r�����U�-�5q=`��V��,QR6�g��]��Q6�)	M��J�Q8X�۫#���K@8���7v��۽�QJ��͵|�MD����w6���]c{I5)JQ��NU��{- �� :8� ㊐m�M/k7���ݳsm �� :8�����Vsu���j7����`wsmX�ݷ��7'�,�+K��&�?����s�P��i��,�/\����3�Y;s�WI���I٩"�\���Z(��6pD͸y��駶%�u�[8,!v;�٭UI��$��� س����i�=<�;�;R������\q]��,]��m�[���}�gMz�m��:I����l`��@ݐ��ŴR����U�q7U.;�t6��Px�C6G]P�m���w����j5��>(��Z�<�a�%��$6�Z���)��.i��D�DN�$t�t1��q�`{<ݨznYn���@>�- ��T���vk�)RA9D�':�U��ɥ��ɥ��ɥ��1%����]�u#cRG�;6��>��Vy$�Gf���E��z�Ґ��N������ͺ�3sn���VKVM,��Q�)"Q��*��,��V&�ܮ����w&�UuR�Z����G*JNA>wW0��t8�Z�0k�5��뛆�K�z[�%)J0�NU��{���ɥ��ɧ��� �o��[��
S���"#������/�hm}m���ۭ,�kK:�U��������R9"p�;�9��K@N{�K�FS�H�G)D�`ori`g^�7�4�;�4�9�5Ĕ� �	�U����� =���H��������@�:gD�9ɚ�WN�%WG�{5n̔e�H��v;	d��_��O����������T�}�Z<������d�J�p�9�4�;��Vu���K����)"Q�HR��͵`gӛ~_�O������ey�S��wѼP�q'��G�Wo8�~Vo�h�6n�8����Ec��s��~0�w�G �?*�4�(X3 Fd���1�"៴�,�C��Ut��h0G<~��ѠM/�����M�|
��^ RDe�D?Ҡs~w��ࠧ�_���������#��^�RMJR$ۄNU�)4�Q�[�`}�\sI��@}�\Y�&ۏCi9��|���#�)MIJ�iUrM71Wq�����j ��_v��ɦ�3w�X�����K��*<��.�%`��Ӧ4����kt}8:ӎeH��Z؝6n����|��JIj�mM��po���Ł��j�ϧv<�k��!���`w��P��$l�R�������~����~������r��5�2g�Q����UQ2%i����ߕ��ɥ�K=�Ł����޵�-b��Wv�Ԏ��p��+������V��n���CN�hi�O/ܓM��w��N�ꊢ��A2R �Vw&�W�m����VqM��?{2��8����]�3"�q"�塹�6ա��9:��F�7�XX�A-��� =�l�K@{��@t{{��9I5)H�n9Vu��G��������X]�-�)�J�BD7����M����Ձ�ͺ�3�uX���Q9$R8�qX�۫���%�=����(�ͣw��`s�4�?nOyp��+��u`N�shgq�M��SL�3���gVx�Ñ2C��3��׷Uo.z�]mҫќ���	�q2N6��dya��D�K��b�ʜn��@��ۥCl�	)�c�ض��ք��:^���a�,�p�t�l~�;ݽ��n�!	�X�.�dY�x�N�NY�$t�N-:}���J�@q�hT�(�6k =	&G��HlmU�;n۟���e�N����]�����f��I��v]�u�ԗ��;UY��)��F�oV�|o�1�C!uCl�#o�>���r���{췉m5=u.ں�	ȸq�ɥ�����ν�`�KiHJn6HDAʹG�@{�� �$���_4ޡI�H)PR;�K:�U�μ�`wri`w�+c��R��6�� �$���G�@{�� ���qN�J3��zy霵���fWN�mƛp��sh��.#A���r���u����ݎZ�� '8��U���#Ͼ���.��rH�q��;�4�_z�i6�W)��n��޵`o���9�`fi�6JR6G)D�`osn���V_�Io^j�3�4�9�bZ�Iԑ��^�n���Ih���=��7��S�Իj�'"��,�+K76Ձ�N�XM��*;�DvusIjt]p�p"L�tnT���m�t
\h-�<�Y�M;NAk��hE���$M�@8���=���_��7�)"Q�E*	À{6x�8�5�ܚXܚXܕ��I�JDڑ6�ʼ���r����r�9!=��t��Ug�t��� H� sw�*��p���wj�w=��� qR�ۮ�3wIC�Q9$�4ԅ�����������gt��ZX�I�=��CVavn�MAq�1ٱ�v���kzN��-�X��
��5�c�n!���O� =}& {s� %ǔ�D��#qS�ʰ8���ܚX�`�q�H	�v9Y{��RŁ�F^�x	�߄s� qR��b��)J���TN|Ӆ����X��Vw]��|���������:�Sz�$Ks4����i ㊐��=���u`f��BEA9�"u$!�ݳ=InIӪ��5v���E��j��خ�0��"RG#�`qwu��4�;�۫76��;���R�d��8�ܐ@w8� ㊐��/W볭ŻFiNI#�5!`gsn��۫�s]���K;�3hn!H�nS�ʰ28��bǰA�UW_��}mJ�7�9��s]���K;�K76�����sQȃ���GK�\1����SU�q׻	��(��6]9�B�մs�ǭ�mNqD��9uhz�4E'X�pf�N��Ꮶ2+B�Ƒ�C]���l�k�m���v^��b!^{Nu�R�gǱ���<��^�%�Z�U[���K�<�k�0�t�=��m��L@�,f%�Y�N��-k�U�h{�ݟ���e�-�����!{9�笖W��ww���}��v�ֆ���uX��-��h�����ND�ԝ&6��t`)�=���Wk���� �q�����`gri`f��X[��-�JR�%5$����;�K76�����`f����dѸ�$J7���D�*@z㘀q�����vV�)&�(8��a�}_}_.�o؀�M�@>{�*@��J���6�p��/w=��� qR�s]���U��)I(�G"# �;��j����\�vɴv��Bq���UvhQ�$R6ԅ��ɥ���u`qnk�3ri`guFm�)��qHX��GJ$9ꅌ@�p	�X�m$��DM���ZX�V��6��6�I�r�N�{�K=T����g����OҮ�ۉHn�nx�߄s� '=��9h��m)RSQȣ�"p�9�4�7��@>�-9��.Yu��{�m3<��iKng�-٘��e�5Ym�`�r�ڶ�E'!$B�%�$#����ٷ�G��@N{�� =�jn�]��^�8��B�μ�~����#ٳŁ�l�`ori`�M�q����b�X���ʼ����!z,H��j�<�X�uX�6J�F�8�R�`�q�H�%�{I��hn!H�nS�B�����ν�`ori`wri`V�(���J�2D4��v��rSfz����Ƈ���]/lP#��$mʒ7�F�,��V�&�G�@N{��Q��I,�mE�=�<_�RF{g�ٳŁ�{���w|��HJnIR8��=�Ł�ɥ��W�����`~�OŁ��ܑ
H�sCt���9��K@N{����o�4�Z��P�m��~������I)&�(8�9:�U���m���,�M,��-Q:q�"˦�h��ύ�蒹eȭ�K�&y�mȐ�{W�ۂW��*)NF' �l�`wr��7�<�M���;gދ���MD�rIi���K��W����߽�����ߕ���K�W��FרnRRG�5E���j�ϧv,䓈��������9�F�r�����#�a���]�`omq`}�ZXsi������tȯ�Ww7!UD�UG�7���<�o;o��ooZ�3�݋�H�Z�6���*b�t�� ��}�=HL5��AG��3϶�������6�!�e��$%`� �sې��q����� �$J$!$�V%��\4��0@�z�R�@�F$�&�&:�,�S�F ��!$B �2H�b�����o���7����m$!��U���
��N��9� ��#�#�*�TJ��]����f�ɂ�m�q ,��N�Uڍgb�8mi6��Fq%q<��Z�m�v� �s�]en;'$�\:�(<�<���j�Xm���<5�l
�Yr���vɽ�D�,r�����C�Ʋuv�Lv���N��S��i�`Ⱦ�g��0t�n�^x5���+���M�H���`�=�m�9����j���2@����һ��v�g��2�3����qٱđ1�Yr�����ӞCkl�L����S��m (=��U�r�h���%m@@]���k��[��V��xꈍ��^�[T��ajU��MJ uP UT�Ͱ����N�j�Ri���[�Բ�x�r���Ry ���^1���Y�~���L����T�r�����k�GF{+�gm�t�F#��g�6��A�y�ܽK�m0vW��; xr��Y#�5�R]���^��;u�vҝ�9�Ր�:�R)T�vv��q,��//e�V�x������������n�o�zGζ�t�#�٩�7,-��3���5.ڍ͖�9�c�f�bл=;5J��+���6 !�+�(di�$�vն�]��1]H2�[솠���`;��ۯX�n�̵km�J�t�ܽ)�3�Ā6��;�EḎ�5[W8q����h�ϝ��.��٣-[AU:��@�/����&��U��Pɲ���[Ş{5�S� L�T��1��4�9�U��^l���x
���V���j�49Y`P�U�0��t�:�"�����g�I��;��9�W[@(���A�&!�4^l�m��l ��HㆶF�v�H.���l�ɂ��r�fKR]7=<:Mf5�I����m��l�ݚ��[d��Kh8�S�6�{��J�vʵ�Uԩ�k��[�9�G>����k[�V�b��I`22�a��6)n��v�=�f�h�ͨz�����D�|�������Q~(~�I5��M7+b�
�����&fT�� �GJ��,S�2��f�hjR����m�o1��7���&S7C�+����Kg+ٞ{y����[�2탛l��Y�9�lK�E兢^Lrj�a�`�������h��̐��b�ȅc`j���a��蘤S��oe%�!<.��T���78ڶu͖���]�N��SZ�6�ѷ'��w�}w��I_a�ͫ;|v�ehz��,%isL��)����p������Te���G���`f�ڰ3�ݎi��}�Ł��O�
H�r�$�`f��_�M����;gދ�����r��M7�?�!7)F����,��+{���^m�ﺼXޯ��&6���UQJ�1Ȭ=�Խ�~,�g�{�KURܛ�`j��J�F�H�R�� >��>�z�y>��`�v���v�Uծi!�g7]-�u�%�"T�r]2D�"Gh�b@�?���S��pT�s��x	��R�9h��Xw�~w�zHە$N�9NG*�μ�o�u�J�P���m��Jx�oui`guq`f�ڿ6҈>Q�o"��]�ښ*�����}���G�@8��r�r�R�Rn9��,?�}����o����V�W�_-�ߋ��Oĥ$J9�m�耜���'=���o�ߟ�����3a�٬;s��L�J�Yb��\�5�6莺�i�v�S���+:Y���8��+{�K��O�}U�͞,7S~�MJ��#������gmq`vmq`gӻ�n ���9��	"mHX�,�M,�o�}�W~��1K�`s�4�9�[Cr�m6�8�,=_/fߋ���`oria�Y�H��[$mʒ6Jr�Nz��?v��6	�`��.����R��au�f#24Y`^a~��lt\�8H�l%(�(�Ү��8H'$\ٳŁ�ɥ��ɧ�n=���)%&�R@�����������μ�`ori`s�uHJRD��B��ͺ@z�L@8��@{�wl���S14�MM+�MGӝ�`omq`}�V��&�I$4ۊޞ�Xf��P�R�E ����ɥ��Ϳ}���8���Ǵ�Y��:jD��&����M��n��m��fɵ�J���:ӕ�D�F�$JB��ri`f��X]�vnM,wbkhnRR)�␰3sm_&�i�d��zl�W�ﲴ����#nT�:���r�-�vnl��s~9�\�r��*Ib��A���ǾVw&�nmՇ�]~�;�|שI)7��ۊ������K�����;gދ6sb��i?4�H����f��'r�IN8H���ļ]C���,��U�g��-�%.�!KK$[�<�W�{r�2�u�3�۶	��Ns���Ӳ��[T�C�ORFܽ�v9c��+�n6e�A�ev%b;X7f+k�v�������ۇ^�����Tڰ��K!6�m`�]�+l�Y.��9��je�s�ĩ�$�ݶ��#���w!��tn'����#���^���׼ގ�i.8+=t筑-/ʊ�%�)��OX,jU�^aw6�����|V��$�
�j��}�j�ϧv,�͏�	�{���ޟ�5�?Iی��)ҎU��N�_�i��zw�������͵~m$�՚%��nT��IȬ��+��K=U_R^͞,ǾV-�����*��**j,9�ӏ�o��k�>��a������`wZ���JE#R�"��3smX�M�V�~zw����ZXkm=�T%H��ƣ�cL7]a:R��cEE��pW��q��I�>�=����������ʒ'Q��F�tk��`f��`sriͤ�@ooZ�>����jꦨ�TET�~zw��_�i'tg]q`goZ�3�u_���l����Ԥ���T� m�`o��X���撈ܞ�7�z,̚6JRD�NQ �,?W{�j���ދ7+K6���~�`fϏUT3Rnfmn���Ih	�`���	ܚX����)&�eJ��l#����K=J��q��,�����)�kp���}��ʕ��7 �l�`wri`ori`g^�2���C�(�cq6�,�M/�D�\X������ ͘��K���Tr�������ν�d�������������9��$mʒ'Q��s7D������U_�/��}�.]\�BT�qH��g��� qR�Ih��!,�3v��]iu:���2�ѹS��j�e�oY��m2q&4�mJRJM��Ӆ��ɥ���u`g^�����q��RD�^mm�f�q�H�%�{L�_��W�����$Bn"6�GDr�nZǰ@t{�*@�ܙw�T��q�n+-�ߋ=�Ł��u`�R�m�p��~�>��D�DT�����e��`�q�H�%�����_W��y��J&�R�)%�VHU�6�:9��Nks��Z�ҬG����-�[���JE*9RD�t����;�uXܚX��Vͭ�#nT�:���r�;�}vmq`n�Z�������j!�}�w�Eڹ��)UL�MB��6��^-��k3v�����+Kmh�cv���ѐb٨�&jh�����-��	@��u7ch]�\[e)I�s���)�~�n)JP��F���*f��"*f�����+Km���;�JR����┥'�w�^JR� FM��k>�ڰ֍fZ�f�'X��=FMz�N{n����b:�m,��E%li���k�lpS�<�ՀS��DU�v�&����Z2.p]J����

����rn�s���뱙,�lec5�B���:��x� s����k�ut��^(!;����xg\mI����F��8�R���l��Nك�l`��X��/�3��t_W���گ���𮣝�ܕ19�jV���g�,��t�:��ݭb{`E�#b�_�/��UPD�AS3J���?6��}�ބ�mk~���@��7i>g��ͮ-��kDoLD�*USS3P����}�}��)I�����D��?}���@��������ͩD�DT�UT�LLU��5��蝍�mo�Z[h��nGt'ch]�\[h@��F���QQJ*�ABv6���f���5�Н��mo�Z[h@�ۓ�v6��gڣj�&iT�J�)TD�m�mY�f�v6�%�}�|[e)I����<��>����)JO��������Fz��L�"B�uX��[�t���څ�n��F�$�N����`��A���-�UL�MBx6����W�m�m_nN�إ)�~�n)JR}�w�<��=�_a+f��3UJjjT��m�m_nN��g�蹑��`�*qEw"���<���7�┥'{��`�R��oKmrN!�	��oAUSSTLT'���﻿��)>�;�H��B��oW�mh�t�N��6�}:mUA5L�*�����6���7a;)N���qJR������Jʄ�;-��O��3J�EQ4B&j���}�}��)G�~��~��JS����R��{��%)O2�������Lݦ� %����՛׆,�t�ȷ�+����,��{������4�ԓG��6��������V�)>�;�O�G� 3�JS����\R@׻���L�UR**��mk76ն��gѻ	���nV���5��蝍y6��M5	��3�ު���SQ*��*�i[h@�l{Н��S����R�&��qy������
F��A0�CHt�6���}�|3��#8Y�u��QM{
���JL�"7W��H%�Ą�Gx��o�G�4P<P>^�� ]"�ڝ`����*��U�@��+��S@����v����/}� ���N���%)O���R����F�D]����J�f�j�6�ɦؚ�u���6��������V��5�F�'ch[d��i�*UI;�f�qJR������J� �w���);�~����������-�v������A1�nzei��Wk�5�=In��p�t��L�d�=\���JN����q�1UQ15QTEP�����V��5�F�'chY�ZZ^�I(nF�5��𝍠mf������*fiT����R��{��%)O���qJR���:'chY�����8��'���"f�*����5	�������5��蝍/$ؠmooZ��6�����mk�[�(��������SE���������JS���R�����py)A�@���yۊR���ֵt���Q0MEP���mf�ڶ�6���;�JR�w��┥'��]�����~�??,�&Jl�ҷ�ulk�k�U]0ٸ�SNȺ��pWl���|�}P�LJ�J&f���6�����mk7+KR����k��R���w��)<��?��sQ4��SP����-JR��ݯ%)O��xqJR����'ch[��iE)��RLPD�m)JO��v���>����)JO{�����mf�im�m_FlUQ15QEL�v6���5���[h@�twBv6��������fn�v6���e-��"f����R��V��5��{��JS����R�����k�JU��j�@���J!&�F���fi@<+Jjp���GG��:���q��V� \��H���^֜O��F�螤G�mv��u�]�p�4�4Mq
أF���E;⃐9�j��du�En�R@#2ɠ�z�:ɻז8$.�`��"c'\W;zwNdr�m1m�H�w�X;2�#Դ�وw۲ěL.��4c�v�pPkE�VŦ�gv�FGE$9�lw�n�����O| ����T���]ٺs��]Ĩ4Z�F�=�hں�x;;�T�3J�ED�L"&�=@�����@ғ�ݯ%)O��xqJR���{�ch_B�ڤMTDL�T�I1T[h@�f�7chY�����k��N��6�g6-��ksI�Q3PETL�3z��R���w��)=�w�<�k6sb�@��7i�@�3�Q�DT҉��J�L�+mh�cv����͋mh�ݦ�mk76ն��i�0Gtj�iR����O�����E���fn�v6����j�@���݄�mk�l�*�E*�Q,ڳHj�աZnH�(�O,ѝ����;9����MӒzvc,}�v��m��;ݯ%)O��xqJR���{��JZ͜ض�6���#6�������T�y)J}߻À@	�@��� <y)I��`�R���~�qJR��ͦ�mk~�[3PD�U5U(��m��}�w�������)JRy���v6����v��'��'d��T�)Dԩ��N��	!5��M��3i��ϲ�kF�df�v6���|f�R&�"&f�gvo{�)JRy����R���w�R������<��>��qJR��w��~vt��5��t:�Rsu�sl���X���y��k����BE9u�c"G��R������)<�>�%)O�sb�@��fm7chF}�6���Q5�R���mh���	���l�s�R��}�v���>����)3#fH�Av�j&�Q%T�'�mkzw��R��}�v����D @!�(���$*)�*�%q@�f�J}�w��);�w�66����1f�I1R�Bj	��me'�}ݯ%)O��xqJR�ϳ���m_��V�[h@�F򈪘������my)J}߻ÊR�~Y����>JR�����)JRy����R��J��*H06Q��$�X����#W4�K6���7s�z�lt>y\���*j�*@��m�m_�3a;@�͜ض�6��ٛI�y(�mk�޵m�m}�>�&��QQ1D��Jv6���9�i.Hp6����n��6���Z^hn�5���'chY��R�������"���@��fm7chY��qJ�$����<��;�]��R����&MD�AQ11P�*���К����@���ބ�mk~�ض�	�i�N��7�;�<��R���TmQ4�j%R�1E���~�̈́�)Jw�}�┥'�}ݯ%)N���������N�b�R@�(� �ٯ�L�tcj(<��f���J�ۖ�'<���-���"�\�M*�QU5	�6����[h)<���<��;�����\����ބ�mk�͒M*�b�E"j	��l�)<���y��ԧ�o�┥+:=�N��6��͋ms�mlF򈪘���
B��n��6���[h@ןg{��JS�����)=���y)��N;T�5U TҶ�7�P3��`�R���w�qJR�Ͼ�ג��$7���[h@�򍞒&��QJ&�LMBv6���9�m�m_�6���)�~�)JRy�}�JR�E>����ĕ�ۂ�������������ӕ�β�V{i�\��A���,��i�u�K���sڶV1ԅ���b��<I�1�;:���ο��}�*��a����m��kSH�io����%c��4�c�Ϸ��3J�\��b�ėWmB�S���	k��->��f�!�6om�n&�ll�puiOH��0�B8�El����x�qD��D!�ԪP���(t�YN�y9˩Q���Yh�:h��Q��j�f���\�Ґ!ͻmӍyB�_��v���4�0T~���5���mk76ն��}��	���l�Ŷ��}�i���"�&&**f&�����+KI5擇#h�G�	��׶{�m�mY��ݍrm	��79GUSJ&�U*ST[h@�twBv6���Nl[h@�f�7ch[�V���5����j�iUUMB��y�&��ދmh���mk~���@��i5��H��=�N��6�g���RLT�J&�����)I���ג��}�}��)I�s���mk~�ض�6����N�3��Һz��Yۊ�ʈЭ�)���XjU��:]ſ��}c낐���-�~���y�ͮ-��k��N��6��͋K�M�r6���z������g�EMAQ�����{��)I�s���x����ܧy���R���~�ג��}�}����Ch����"f�*�Q5*bj��J}���qJR��ݯ$?� ������@����������TU3US3T[h�hJ�{��D�~����)=�w�<����/߶���6��؎�D�(��"f�fbi���>����)J?���~���)�����)JO��v���:#��l��]@\��O/3�;ZR��gAQ�9�\9�u��ٺ�w|�V&��p�߯{��������ٵ����fn�v6���fڶ�6��>�6��W5EQ(�����m}�\ZKÁ�nw�%)O���8�)I�s���O�06���&�Ҙ���U8���@���߶���=�����Q�R�A������~��R�����q��k�Ɠ��*�"�&����n��y������@���z���ٵ���5�@��u7ch_F�T�J���E���}��	���ە��)>����R�����)?��+�f8������g+s���5i�8�,���q����%����q?8[���jT�T'�mk;k�mhϷi��=���┥'�ϻ��JS�=�biU35U3T[h@�}�Mؼ�8��;���)JRw�?`�R��6���6����!3J"�������o����}�R�����py!�c%����mh���mh��Q�DT҉��E(��V��&%Yѽ	��J{���qJR��{ݯ%(5���;�؇��Sρ�m�8�)I��v��"�\�U�TUMB��6�ޮ-��_��(}��7����zն��}��	�����{��j`�%QS%T��$�6�ʎn���Ͳ�K��uI�,�q�gf�JiLQ*�U(���@��7i�@��}�R������~���=���m�mY�<UR������UJ�i�R���xpʉ9)I������������)>����O�a�Os�;����Dҩ�14���k:;�;R�}����
)�w��my)M���V��'�(��"f�*�S5*"w��J�!=��~��)I�����)��w��?�D�O�g��<��>����&����*j�j�mh�ݦ�)J{����)JO{��%)O>��qJR�W�$:Fh|`,ll���l\�����h�B zN����a�I�e$��-�RI(�A	��`EY��:!�4�4Q:� �Q�A$.2���;31�ZtJ;�!R%Ċ�|�Xd���Pن�{��y�D�d��>�P�<&=6H��I�|h �$�,��,+`���CI%^��#DC$L�I#$�Hh_|�YT�U%YP�I"��XI!�[����~w���ߠw�I�Z�[j���6M� �fѶ��ƻf�f`1J9��X
�
U���(&��L�4۠X-���;��*�]B��ڨ�iv�=���fkReƃ�V��cV�F3f�J�K�t�U�;KtOc[u�RW�uź����a�)Ghvm/.{n�c��M÷�m������\�j�m��6m��M��kz���n6�4��l��GO���',Ƚ��%IR�,>�Y@C�*6�$l�R�VکZW:�TNм�W �$Z�c��iӮ�+])�[�j�VD"1&��� ���@L�U���KF7�'6���<�-: ���ZJӶ��6ݖ�۪����f�,�6`l6�v����\�ջJ��lPgU�5Q�@9R:�m��A�UUl ���8�W�8 ���oS��+!4t���ާ:�Ѳ���J��*����T��3���=a�C%β�;�x�f��oU;LY��֌f
"y����gTTn���w�s�	��f�VEPn��Cs�)؉��8�v�)0���hLt�p��+hu�q��\[)��{�\����7At�:2�*����c��qZ�Jaz	^c�J��`Ƶ�=h�
��
I����jq���l�踲�ΐhꭳ�k����T�����)m�n���ҩ�֚��0�@N�A��[M��Y����']/Sѫ&0eݣn\�P�UF��H�2i��RP�粋���nJ���1��.��@NZ{iG&7,n\�cD��c��K=v�"743e�R�>uO6TUۍ�*��k�ul�j�Ӗ��(�E���45+lhM��\�=R��sR�0k�
 F݈���EJ� J�UPq��յ!�ԫV�=,A�ӣh�]�ƭ����{g�)��J�Q--UKv��[zڐ5�8{n�XHemS�.mu<��j�qΩv��s��]`�Au���[��f�mx�ꎤ�ҹB/m���w�#�.� �&
����Q��(���S��"x���߿{��n7�)�r{���Gn�Nۤ�e��rp�-%r)�s�]�al��YPql��y��ȅN��#�j0�aWeP�����R�c�@�kB��i�]s�ųЭ:��n��h5��B�;lu{Cjn�\�������-TTǶ�;�8ׯL����S+���6q/*vݰGh�P�+Y$��U3��hXZ�I����G8�C�k���n��!v.fڝ��X��m�su���$c�*T�{^�O�����Gݖ૰�#{��JS�~��)JO{��y)J}�}��~P�%);�߶���/{��n���QT��5SJ�@����N��6�g6-��k3v������V���I���h��Ҋ�SU$��ED�v6��ޞ�[h@�f�7chY�����k�ݤ�mk��A:M)�9�[���5����*#I�����)���ÊR������R�� �{ս��5��T�&����UT��%)O��xqJR����JR�����5��M���=�f�UUt�δ�g���fz��++0����i��y�#;��wv�������	���)?~��%)O����R���~�n��6�sm[h@���'d��T�6k[њ�ǒ������	��	*Y Chi�m��|�����6���3��[h@�ۻI�כhN�B��4��"*&J������6����n��6�sm[h�P5��I�����E���}�n�L҈��D�ELM7chY�����k�ݤ�mk6sb�@�����mh�yTEM(���Jj�����}�����Ir���8�)I�����)�~�)J[����0~�kzy��ڝ��i�g� �J�EF+{.�V4�>���ܵ	�W�Z��R������)JO��v���Y���/4��7#h�w�;@��OA>&�Ҙ�h"�"f��@����n��VC%;���qJR������*��6m����#�&�DMI4��F����?}��8�)I�{ݏ$0�R����)�u�s�R���ݦ�mk�a�EIJ���iDEM+m~mz����I���z{�m�R��ݯ%)O��xqJR�����TLҥQJf�D�'chY����5��M���nm�mh�wi;�o{����py�r��%���v���ƕ�X��/c5��c�A�76�h3�����X*"UMLMT[h@�f�7chY����)I�{ݧ��JS�����)JVi�4�*�4ELM7chY���JR����JR�w_w8�)I���v5��hN���:���Q5SJ&���l┥?�BP��߿�pJ��(O3�(J��J��(L���(J!(J��;�}��x%	BP�$BP�%	Bf`�%'�#BP�	BP�%	��(J��?��q��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	B~�����P�%	BD%	BP�&f	BP�%	�%	BP��Mh@���'AT��"���vog�(J��0J��(H��(J�������(J!(J��?s��y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	������(J��0J��(H��(J���(J��"��(J������(J��J��(L���(J!(J��O8��:�t���3�(J�������(J��(J��"��(J3�(J��J+�
��������9MA�R$�\�%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B~���x%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP����x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B~�����(J��(J��"��(J3�(J��J��(N��g�	BP�%	�%	BP��%	BP�$BP�%	Bf`�$&�4	�z|���J�������WF��R7L��vs r3vP�U�[f��G2�����8��t���v��۽�w�n�~��(J��J��(L���(J!(J��?~����(J��"��(J3�(J��J��(L���(J���ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	������(J��"��(J3�(J��J��(L���(J�~�ǂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�ge�ճvovl��kg�	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP�~����(J��)��!(J!(J��5�%	BP�$BP�%	B~������(J��"��(J3�)=L��"��(JY�P�%	B~���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'����x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B�11�&iR��5R��V��&�2��0J��(H��(J���(J��"��(J�����P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'~����(J��0J��(H��(���(J��"��(J������(J��J��(L���(J!(J��30J��(O�w�	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'��E"�����SSU�&�4	�M�	BP�%	��P�%	BD%	BP�&f	BP�%	߿~��(J��<���(J!(J��30J��(H��(J�������(J��"��(J3�(J��J��(L���(J���ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	������(J��"��(J3�(J��J��(L���(J���UH��*bi�h@��&y�%	BP�$BP�%	Bf`�%	BP�	BP�%	�����P�%	BD%	BP�&f	BP�%	�%	BP��%!�d%	Bw���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'�����<��(J!(J��30J��(H��(J���(J��;���x%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP�"tD��C�b
hQ?o*9L����+�����ټ�݄�q�$�ݱ�m�[N��C�����m�yɢ&�pU��SLq���t�ײC5V�e$��`عN8vѭ�'����n#��5����v����{q�Ůn��[
�c7 ��ƶL�`#f(��RM,d�j���A㶚�S8Ɗ�72��Ķ��ۮ�zJq�"�?���W����8D� �=M�8�)�ZF�8&"�"k×SNɴE[q�il:/Ht��3�v3����;%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	�����(J��0J��(J��(J3�(J��(J��;�}��x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'~����(J?�L��0J��(J��(J3�(J��(J��?~����(J��(J��(L���(J��(J���(J��?���R��
SH&�j�@��&�O3�(J��(J��30J��(J��(J�����P�%	BP��K��%	��(J��(J��(L���(J���pJ��(O3�(J��(J��30J��(J��(J����<��(J��(J���(J��(J��(L���(J����	BP�%	�`�%	BR�	BP�%	��P�%	BP�%	BP���r��[5�Y�[��vk[�<��(J��(J���(J��(J��(L���(J�~�ÂP�%	By�%	BP�%	BP�%	��P�%	BP�%	BP����x%	BP�%	BP�%	��P��"J!�����؃�h;�]��|��Ι��VkV��kb A��%	BP�%	BP�'w���	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	�����(J��0J��(J��(J3�(J��(J��;�}��x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'~����(J��0J��(J��(J3�(J��(J��=�l��f�n��f��ֶy��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP�~�����(J��(J��(J��(L���(J��A�(J�����P�%	BP�%	BP��%	BP�%	BP�%	��P�%	Bw��p��%	BP�f	BP�%	BP�%	Bf`�%	BP�%	BP�'w���	BP�%	BS9	I��o�o�=-�;U��6z������˫�M�N�<��6�B2�e1�p�])�9	Bw���8%	I���ǐ�'�͵i{�&�'"h�{�Չ�Ml/{�iTDTD�������&����N�B(��%)�~�)JR{��c�P6�g6-���~m��[@����(��D�SM���{�j�@���{��)�u�s�R��}��y)KG��mQ4�j*�4��i[h�lJ���;@�ޝ��6����n��6�sm[h@ֆ��T��!R��[�ly)J}�}�┥�{�߶�JR����8�)I�{ݏ%)O��m������b%&v����ۓR�ՎQ�S�ΐ�\��M¶Û��͵5115��5��M���nm�m�����~U/%)N��g�)Y���(��"�f��*&������V�)I�{ݏ%)O����R�����nƼ�M/4�'#k#��A��H�S13J�@����'chY���O���� ��<����k�JS��~��)J۽-kf���ojI���m�Bkz���@�����JR�w���'�Y'�����)��x�D�4MDMT[h@��m7���Ow���)>���ǒ���9�m�mY��N��*�)M"d�Et�Nn�.m��Pu��n��V�^��S���F;Ol�@L҈��MR���n��6�sm[h��~�ǒ�������\�����M����puQ4�j��M)��Vڥ);߻��I��d�k���R���w�ג�����8��G�֔��6<zB�UP��P����mk�=��R����^JR�w��┥'��i;@�72"4�SJb����5�%�d����^JR����8�)I�{ݏ%(=A]��<]�{���h@��M�QRED�QQPD�v6����j�@�懝�I�@�ޝ��6����n��6���C�T�f�*��Do,O"1��Y�,QE�\��Sc�������V(���nI��{���ow���JR�w_w8�)I������JCk{zն��	��;�3J�E)�R��ǒ������)JR}�{��)�~�)JR{��c�?�D� pu-l.�TEUDTD�55Qm�m]��ג�����8�?� @d�~��c�����mh�"7d&iDUR&h���n��y6ؚ������k;������q���Xo#����QT��5SJ��wn�漓�_z>�޵ʾ���ʿ�:/�����q����ݐ<�u'���,�n�fӋMsg��`�\���Wn�����՞�m��46B�n�ݽ��02�{;����YU�ѷ
b�q��h+���T2�a�y&�$��+��K��c�u���U��Y���lsDm'P�h����q*�(�fT��G҆�Ldg��sG!��Ҁ���ѧ�\7J�Y/߸�����?��:�Ӊ����)#[�Z7:��qW]�W�0{<�Dt҄a%I
R�*D� ��j�37mX����K�wu�n�GJiLQAT�f���ݵ~I6ۈ7��X�z�ך��W�$f=�$�Mʐ6�i>�*@t� �- ܊�ף؅)ʄ�6�V�m���b��͵a�&�{{���r&iR�����75 �c����HT��Ͼ�?��v����C�EU���ې����ٚ/X�gn@r�5}�wg���b�(���S�p{}u`f��X��������}O|��[��JII8�iÕ}߻ÜiE�A��WI�
Rw~�;�E���j�����ELҙ��D�&��X��`fɛ6y�����]X��Ձ��Ma%I�R�r�͓6l��Vnm�6��m$�}�v�?{�/�R�7�8F8��۫�oo~_���6Lٰ94�.�'�gV���.zrE�����R��Uѭ��9�b�;�Hj�{�����챆�Z����>���RG���*@{gIڂ)M**��BfiX��~I%��IL��;�`{��^K��������DR��q�5����ͺ��}��y�+h��M*��1�p�qV���!{&�@�h�`eqݭ��l�kT�ma����V	%$��d��V	%��h� �"pQ>x(c��ZP��<�50*JL)�!$��ǁa!#f��QFY��
����d�T� �z(?:�	�J���p ���+�h|��yÕ{��u�:����%pq&H�=_U~����=�����w�XF�́�&l�d���(���&�*biX���y&����>�����`fn�X��jp�p�\���O/3�;]:��g@��찃�9	�wV���ﵤB7)��Jr�Ⓒ�o����ٰ7smy4����j�;:}v�D�HR���7��;w6���ͺ�:�u�ꯪ�n��5*SpN�c���� qR�I�0s�ѲRr
&�IQ9V�殺�}ʰ1{�l�3f�����-��!�����ͫ��1=�Q��$�nU�ջ��s1 ܊�8���>�}�w��uK�S��3�� ���8�T�v�l�j��od��?��w��g?vV�4�?����}���T�q�H�& :�nĤ�D�I�;3v��T���]X��;5����5���II)�)Ɲ+7vՁ�n���DoI�6�u�t2lMʎ'R��8�����T���v���`fnڰ�����;:�.�Ȕ	
n8����?�w��p��g*�;��z��EN� b���o��l�7]���	Z^gX��v��r�D8��ך�Z�ׂ�<��[`:�vqv׷/%'gO63����w��knÑ�b�K��ng�Ң�h8cY�Ӈ<&�4q��-�ؕ��������u�qiN���n���[LF'�H�1�ͤ�m�apR�J;�s��� �G<Q۠�#�6JX�#�� �uϬAܸ;�-���5��wo��w�[�����]��=uz����ܓm:ݒ���ܲ�s����JƥJn$�R�d�@�~�Ձ��u`un��U\A�g��n��' ����6�i 䊐rL@9���nm���͚�~O�B�"����V���6l��g�D'���~{�Հ~�0���($���v�[�{��������Ձչ����i$JH�I����>ݵ`y5����_�����n͛~��G��vRع	�v�FlXn�9X�y��uI@��ЛZ�������q�*��ݺ�:�5����꯾��z������7*8�HD'�`unlݤ�2������ۋ~s����������۫�kM��]�Ȕ�B��>�f���۫?R[��Ձ���`��ѩR���"(����U����V�}u`un��T���;1��NAH�jPӕ`f��X�����7������u`enq���NB+S��H^g��8Ւ��:��Z�u-lFfBd:Q�d�HH!7*����`f�u���_����u`ye?P۔S��Oq �b� �R�I���vb��߅$I��qRd�������۫9����V�5����5���� �iʰ��K}�r�^������a��n�ܫ��#r��ԧ(N)���b�$�r*@9"�߫�ߟ���W~�[�y��Ԧ����}|����tTb�:�E�Uy/$������G#�ž�x��@�=��g��;3v���ݺ�:�u�7hԩM�:R������W䒈7��X�6l���i6�ݯD��R'NU�������v~�K|�y���Ձպ��(�!#dLҰ>�ݛ6Mٰ37mX|�5搐���`��E������8���m�"��i9%����`~�ݽ�~{�Հn�Ձ��x�Rt�U�s+��֝9n:	zl��[�`�\f�5�fzݖA�!�N	�#J&�#�� ���Vnm� �ͮI{����;��	�B�lrHӕ`f��X�l�3Y���۫��$���t�N�N�[& 9��@�mR����I��J�AJR �q��7���ݺ�3sn�?|���v}�'�R��r�vr*@8�\�`� 6���w/�w�9�ڲ�@�m�^m�r\u�òqve�������똵�����K��3ѝ��Bd.����,���й�P�Nv�2vU�6���3��`b�:6li�M�II9�7q��kX�9��h�N�۱H�h��\�u#m�i���O0�F��M�ں|��f��x�u=��.vTΓc����Z��cj1��6Z@<���������}��+�V`��Bq�i��n��4UΙ橳��v�q��en����٠��F���ʐrL@9���nEH\����B2F�ܫ�w]����`fn�X��W�H��4���(�S��D���oM���j���iDooZ�2=�;���z������$v���Ԝ�{�+�޵`}�6l��`nmD���c���X�۫�w]��fk�37n��_R�~N�m����׫e��:�-�	d�;t�rZ���&���wv����ܰ���W~�߇���~vb� '8� J��봩n�)U@A5Q��7���ךJ ��`{7�Vq��ȓ�r�'�S�Ỉr*@F�<�����4r$���ȜQ9V�W�������ݤ�?���m�A�_�r*@;�y6Ȫ��*J����V�;�`y4��i5�=�Ϡo�~��9��V+��k9v+[5�1k%��:^-)9���mU��CKZ�H��4P�(nS��7M���{��q�ȩ �9hpp��sw/"d���Q`f�i|�MD�֬��V�=�`n��n!H69�,��Vl�Ş��|ܐ妔���^M����S�V���X݉-�7)��Jr�76�c����K@8��T�9Zn�%wW"��@�\�O�V�m���Iw�����{֬�͋~�nyLk�6"Rgja�"6�v�洹�C�v�}����n���d�<U���qXzt\�X�ZX����͎m4�@v�����Ȓr
I#RB��ݺ�3g6,�9�`f�i~m����'����#i�*��=�7)�?}_WԖ�g���]Xh�v��:�S��6�7�Ł������j���_RI$���'ʹ�z�"��ø����bbd��ʼ�@8��T�s�u�Z6���o�~QE��p���f.�dm�v�ۉݦ2��
�1�q]����j�����ݵ`f�lX�wc�i���l�`g�^�7)��Jr��U����ޏ�v�ދ7+K~ݵ~i�/��Wur)N�E�?z��+7&��v���y���x���JA85"��E��m$�{o���Ձ�9�a���^ڛ�`o�x�!9#$q�B��"���#�r�=�TTw��H8�����{�Ow���О),m[ �!�	�c�b�)H�
z14�bf������k
]���n��\F��ξ�P47��*AB̤z""�H��"�"!rW��3�b6,�;�����~����U�U���v�8Vj����[�6M�l;i#���h��Y��`*y%��
��h6瓎@Kks`�rp9�EҮӢx���a��>X���6�,6�/
�� Gd{;OGN�����z���e�sf�uJe�[j㗤����#O-�-p�Μ\�0�h뱷`�C��%�kA*4�۪N�զ���V�6.:��,�ۧHEI�r�Hi��Z�%񹺒[c����>�e��B��ƻl$m)��y���9rm1�ݺ��]��cc��4'8۱�k�p]j�۱�|q%jŴ;UA8$T#6ؓD:]&�89f�� h)h�@�/�J�������2��-�f�.��v�b��-T���y�^^jݥZ� 
��D�ʻJ8T��F4�A�UUm��'-�*�W!�d�(lɚt[Un5N^�N.9�쨛��Um�U���$�����]W�e�k�EH���k]%� {Ny����9_6�T����GI��dٮ���S�x^B���X��n��%[����

���Қ���E����InY�3�#']s�\� �.��B���Ӝ�0�҆���垕�X����u+�,�����c��R�$��j�Q�!A�4�H������ �L�,�"�M���5��n�8���7iP�#:i�ہ�ex6�s� �wk����v�7N81��r�A8�t��b��m�A2֝�5�f��[�pd�L�(t���(h�24݉]:fu�d�[��P�G��B6hr�	Ƥg��+ ��l�X:��q��V���5+(�G���ٖY+l����I���H^�m:ȋ��*�r�r����� -��Ԅ���#m�H-��q�t�`��:]���������+�v�MU�s:ڛ]�� mZ�J�6�����AӪP�������Z�n5ɫ`� ڮU�:����η`ygp�q[m���dU��ܥ���':����@D��B�8���lEG�� �*��|%�p��,��7f��.i���"v �e)N{T=$W����!WM�Ƴ�������/n�m��J�cO]���N�c�+�pYk�J�����C�	��%���l�\�s��V�Vr���)B���Cǎ�����.q���u�L�z��ユ��a�<�Ƀ00E��酴n{&�eI���ɺ���/6�]�n1�5{/y�woz8j#���k,ө�� �W9.	��6�h�
Y�y�ٖ�-�"2F�nW@�^j�7)�7&�����6����֬QǼ��R�)MR�35�$��`��EH1�_UUUZ7�|G�q��n����l�`odT�s�u�Z<�036�����Ҷ�D� �-c��W�����v�^�z6ܨ⒢�8�X�K@WҶ}~ϾT��"�����7mX�l�*�@�6���\��Om�9�|���)�T�/��UUe��ur)N�2�v���o���"���UW�~�7^��C�)H'"��Nsv��iCj�6Ձ�N�X�i�4�A���8���"E�`no����V7*i`w7n�,��!I�d�134��wb����K�ݵa�&�no�V�7W��)�R�����ʐ@s�R��K@~�������ޫ#�l��U8�$^��\PםU�΃h��n�vB�:3�����W�U�g�5��Z�77mXd�ǚi/��{����?!��M���X��Vrwb�ߔ�Ł�nڿ6��3�����R⒢���Vk����������\���I)��Z�7wmX�����j�R�HiH��U���?~Vo�u`nfڰ�_ͦ�z��;g�cȚT���ݽ�j�m�EH�T��Zv��
ޭ�dm6�$n
�&:���!{<9���f�]mԫl�NʝaB�������p�)$D�)+�{w�Vq�{OuX�۫��{��B2F�NU���-:�K@s�R7/�����>>�ӌ$�$�#���S����ݺ���%��]X��V-�*HFӑ�i��f�������$��uU��+������`fj�PӌR&�qʰ#qR�IhU�1�EH[u&6g6���Z�NQ���z�.�S5�G Q��+�Z7�������hV��-w�a���@N����T���H<�T���WTE(� ���b��$�n ��`v�Z�>�݋�J ܝ��DҥDMJ*jl��V�͵g6�Q��Vin���4l����H�"r�n*@s�-�� ��~�s�H���!I�d������U���N�O�3{�X�6Ձi&�v��M����~~~~�(��lZ*��ʱ�R%�{9����1�h�[]2������Af��'M�7Lp�k�;�������K�*t����Wv
��v��1 ��f�t��%�eL�"6�p�Fkml.���R6�8��/j���k���yֺy�Խ':����ម;lmϪ$�%�Ǝu�![��'a�d��ܶ`M��kA�+u�ݺ�	�ts+����<�f�77nf��;F^V��l�b�U,<�lr�4�&���8�FI)�n,ig���������72�ksk/6��@s�R��Hy%�=V�]������q�D������@s�-�� 9ȩ �6�3k2)*(�ܕ`w�9K3]��ݺ�3��Vn%Z�%˫�Ju �R.�]�6������֬�͋�I�ۏ��9}�H�I�
:	��ʭ�M�B�^�sHS�*,�������qXgMɛ�ϾT�|�<����b���i9#��DNU��ͺ���U}���U!e}�ve�u���]3߿k�w7n�]��!I�d������Z�q�@s�R��p�bq��ܒ�qX�����n�X�۫��U��wI$M�*9M8�N;����T��Z�q�@%M����-�����jtf�f��[q�Ș��aK{N���b8 �Bb���M��*@s�-�� 9ȩ ��6�7�Q
9*��=�`r������T�q�L���{YY��wU��GoM��nڲ�4������7ʹ����ڰ2;�l�r&5J�UDQ�{�y��T�|��� =W3]���[��F�9Vw6���Z�d���"�t�/כ��[�kP�y����gL�V`bk��n��T*�M�[�'b��)Tn�m�??����$��*@tqRݓ.�^n��������i#se@;��V��=UUT�fa�D�r�9N8Rn;}>T��qR�s����8�"l��G*��_UR�ܫ5�����_w9]D^�
�?)����喙������*��t�nTq:�����@s�- ���@s�R��H}]�}�Q�e8H�M�F�Q����m9��9~�;R�g"Թ��`�lN��}�ѿ�=��iH������`w7n�nm�����V�bo�9R��BR�SqXr*@z8��$���-�~�#�fy
H��)R�����]XǺ��<�`w7n�,j�(FH��r��K@>�r��T���}��Ԁw���dR
F��γu��ۤG �1*�T���nɚm�v���BvM�\�6�d�%s����K�v���+!�.��^�t�/#��k��Xg=��r���2�Gr܎x�T�	'5D*��:�����|<})㗠�X�h�V5��b:9�b���2��Y��%Ҿg��P�sw�GF�j�3��@Vq<��v��pKJ�2K����5#Ʒ=sΌ�xdgs����w^�;�n�اb�WY.��t6��ͪ�'c&�蜶�5ln\�@.Ū�nT�)�"c��o��Vw6��Ź�������ߝ�����r
D�ȓ#�`tqR�s��8��#mʎ:r��7%X�5��n�?RI�L��֬�zՀn�A��v��f�3L�����؀q�H�*@;�;��Ohr�)������ͺ�?������7�ދ>�vl�n�1vj�f%�ul�q�i�ݙ���t˪[:l��^��-���e�TMֆ�߸�<�����T��e�e�TE%T�1J��'v.���m%m$a�$�থ<T�y�r�ޮ�\��ݵ`}����6�@fq<MRTMR���7�;��ug���o����+ ��d���Jr�r(8�=����Ԁ��*@s�- �1�m�̻�"t�MG*����XǺ��3]��ݺ�1i�*St�6㑉�Q�8͛F�br܊[����vG�"�S�!���|�ܨ��7%p��+:��`w7n�nmՀou�����pnE�#�}�r*@z8��$��v?�����)ȕ:�c������nm��m�HX�0� �h�H�/P���0�)�	� ����LRLH1y�aF�e�F#0˅aw5�> Jx�J6��47�kf��ıM&��,* �+�e��u�����5�g*0D<P�|ac�ı2���$1�0O�8��	� |���\7�Ә��`	8��i�=T+�6���=_;�%�:U6z���(|?����=D�V��K�KJ�\�Ł�&���4r$��9s蜫��u`w�3��vY��*���o���B2Ff]���s�s8�����]½~AJ8�LR��$29�v4]*6�.Hk��r;A]Ar�Us�6l�蜥"�G�7�vn�Ձ�ͺ�ߪ��<�~�����H�nT�*G"���rEHG �1 �1 �۹�)"R&�Qʰ9��V-�v{��v�޺�ԑ�y)��r���r��R���q���`nI�6n�	�����X��=?�����T�ܑ��;�`y�%���_��Z�27vl�c�獞�\`��΂�R�=t�L`�諔��<����d�4�.������6�H����& V9h	�4�!Ir'*�V76��W�_�l���6j��X����8���7�����$ci9V�{�����Vz�-��u`w���q�$q�9JE��άr�H����& �7Mc��%I$*H��۫��}�o�\����r��5�s�h<@_��J� �����~~�c{����Q;jhڶ�cr�vRu���!�sB�^��F�f�t���;w�c�U��:���Fon.[TԖ�+'�t�G<�����	�xv�su�#�����ڃ��vӶ�qpZv�tJ�rIc�R6�E:i�gO\�^#F�?�=��M-�r�q*���<vҪ��E�6
�W���M�c%�U[���4����w���}��~i���G]��g)�2�ۛ"Ɛuۢ�VyR�'[�*�v
��AB�6����T�w$���- 䊐�Jkr���r�ܕ`b��`gi��� =T�$O�ҥ���n��f�}h	�*@z8� F�7�Y�ԩND���)'��^�{�`7>T�w$���L@N�/sn�wosv�M73i���& =W�b��Ձ��6G�q�pQ� Jr��v�F$s��j�)��kF�5��'A;�,Q��/kw32�i �I�ՎZ� =��V����i�D�$qH�#��rզ�Ka4�6��胯�Ձ��Z�1n��6B1�J�E"!#�3wmX�6՞m����`nI�6nlZi�$JFڑ)%X{�]���`j����3]���u`su)�m�r:����@;�b�b� =T������.b� ��Ԫ�2AV6����Q��4s��-I�^y%����m���>���ՠnH������۫��u��j������jT�"T�JNBG`f��_�I4�A�oZ�6;�l�Lٿ�A�;�H�$QȤ��r��}u`b��c�I�$�RiV��������:UTUQDҩ�&iXy��l�t��oM���u`ssn�{��ی����*l�Lٰ<�{�ߗ�>��VF�́��ioj�9UN�T��
T�*�j*��gƜ���2}�RM�Bp��B��	lڭ9�*FI� �{�V76��Ż��γ5����LNA8�R%$���j��j ���7$ޛ7vՁ�v"���NGRH�*�Ż��γ5�����{�V}���$��o�+���N"f���M���n���������Z.#3<�����̗�$ 4� �)�����������͛�2"Rr>q$�v]�K�����ޤ��z�i$���|�I*]��B6ۥ�Hz��\,uӷF�NZ�4u-�n�J��hxM�'�
���p}|Tb�X��nߠ��r�Ēǻl��Y�f�q$�v]�Is��
H��G)��K��Iga��Ē��tZI.no+�I%��1��#�FZI,�3_8�Y�.�K�$��M�V{��~���\�����BT��1�>q$�v]�K����K��Iga��Ē�z�4����"RJ-$�77��$�����g��q$�r����"#7j�q���JN� B �)��H�t����<�լ��a'��Ͷ n�E}{�ztǤ�p��h-��X�]5h��d�6=x��z!͛Rt��3N����Y ��6�$�w7F����/���:�&1p��FET��/:dj��m�4��ѣ��<�"�I�bgmۆv��찠X���o1� �G@���+��������d���o���f�7���*��/FY�.n���ΧۺM��GaacM+b5��V����R�3[�s���U����o����3����R)+5$�?��e�����f���%���-$�77��$��o�Wur$�TcrFq$���>s��_}UU$^��]�K?{�+�I,{���Sm-�+�jT�"N�F
8�Ē��tZI.no+�I,{��I%����I-O5HJRE9 �ܢ�Issy\�IcݶZI,}�|�K�}�|�޾Qi$�M5�
H��R�9\�IcݶZI,}�|�If�-$�w7��$�f�|�Mɳ������%>1�Ӫ1�u]q�KG �.��Y�����Κ�c-$�>�q$�v]�K�����}]�Ik����K�u���r�M�ӏ�I,ݗE�:��`���r�Ēǻl��X����͵�?;M19�mH���I%��r�Ēǻl��|�ܞ��K}�tZI%�Ԟ���E!"��ė��ꪧ���-$����8�Y�.�I%���s�%�Pm�%wW"t�D7$gInOys�%��贒]��W8�X�m��K�ޭ49�C\�d]�.
�3l�u�+M7Y
໮��"S���lWtԩND�J�#�t~�������U����/@e�*�E9 �i���d�;ܺ�;�uX͚_�H:i��REqJT'*��޵`gӻ|�i�m&������9��V5���&�#����U��{�`~ͭ,�6Շ�Izw��+:zOL#���q��`s6i`wsn��mՁ�{���vlD��H�Ɣq�RCE��6ts��9���j���9�ٶ��ݮ�ee�N6ԉI��u`w3n���V3f��Ԟ��)�#�9�����U�O����@z8�~�>� ��%wW"u!7%pk��X͚ :8���H	�[������y[[�SU�G��Ł��j��3mX%M~��UߥJ��d����&�R�(�$iB�m��H$T�}�Z̒��������v�:#���YA.��S�]�Uٔ٫��ɣ,��UuDM+7vՁ�N�X����C}޺�5xK��&�#p�P�`g^���O{g���u`s3\#�D���j��͝ذ?nV�y��F�u�q���9��&' �m�
��`w^� 䊐��@9�Z ��y0�r��r��8X��Vu�5���ܫ��0RY�p|XH���֕nԒ}Ҿ�.�WF��S�Ӗ�Nl9{���a���
f%CYP�
H��.(�R���D����: ���Q�e$e�JRX f$a%([I�Ѡ��G����Q�P�W1�A��0�H�`A��� �Dn�s����HeZ�-�}@mp� �j�:�ͭ�7Ke^���٭�m�$ ,��u�1�� �����4#�U 蔖r�{m����q�0�[�Q����8�Wf�V��r�^7
��|�����׀�GE��d �Y��[{CE3�qK�i��Q&�`������:S�FV,�#����eUh6-��W/k%c5T� �������I�U���Ζn�zʛ�n��-�R%g:���<=���� `غ��Ԙv�5�m�+u�n�n��)�v�Q�8���Z1��D�:�%D��k�5���C�H�T��$�`��On���U�h����������6�H��eVȵH+��մ�U@m[f� -*�f�y��@�UUV� �v멩{nxU��v�n��L�	`��6ĺGJ�v��>��r���ǱQ�lO��N�n��u���b�4��К�~��&-������:����,r�M6힞��S��Gk:��n�-�v������%[���M���< �9VNHג���0�ݵ���� -�]E.�̧fv�Y5͑e��66.�FD��i�-'e�2튱��� �m��6�i<SB'#M�����v������z.F�ֈ;HG7ZM��g��K�u'nq�fmr��e.��T*�SV��j��Sp�*]��d�fg��)ƌ��t9�4�<��h�����Nܣ@�Ŧ��w\�BT&T
�Rt��q�ںZ��em�u��M��U)\�1�� f��j��V�nvxJ�w-�.�K]��e���T�q����2Ͷ�\���[)�.��:�F�v6#:��"����.��T���l �nImt���}�����Mתvi5PØ1��j�3�.h��Hv�Im�vi��D1�U\���Tw(��(�s�$ɒ�j�]�:m�[m�y�u�3նT�U<�3�l8,Ȯn978yW���/7E����~w{�߻�܂��)�g�q@��+�D�>
k�J�㊀`�>���?o�䳍���nׂ!pi\�:��7//�ȓt����V`�ӓ<��1�l]+Y�mۅ�H;61��v8�9�� �Xa����v�j�{\f]����5��1�g����r��ٕ�]I�F�l��>6T鵑���kq��s��u�y)�I�ƶJ�=6�JY��������蚗��:b3����H�:�&�Oj۬�:�Z�Z޷��P�p�>�]kE*.eu���o��&���o�N��Ț��b،�T�������KԮ��N�"�k�	������-��H�;�MJ��IԨ�9���U��UU}I�\X�֬�wb�5��m)����?Tr8�$iAH�����3wn��In?yX��+ �=B�(9JJ(rn�>�ذ3gv,<�m��|X�K�cn"7�8����������/� �߄� :��]{ZN�Α�u��ٗ���9W�h,I��U�K9������k��bg����~ds� H� �����ay�\���QU�����͉.�*z�K�&�N����Vl����r��8����r��r��8X��Ձ�y����G�@N��J����6���_���&�I��_����ux�?nm�F�ʰ3��MJ��IԨ�7�������T�}�Z�0��7��u��e�unډ��z�$��]R�Ŭ���fc ؄"1H�r8�$iR�76Ձ�ٶ��sc�6�O���ŀa��!I�%7*��sn���U$n=�;��,nmՁŢY�m�Q�T�U+>�ذ?}����M����_��UU�Q*@w8���&B��t�2��TMTXy��iG��Ł�oZ�>�6Ձ�y��;���N69	���͵`zhmfoZ���E���i`a�?�5�"�v�+��r:�Ӗ�!)�D��'U*�er�����w��r�4#�!#���u`g^j�;�4�9T��,"?֕%����Ff�׀�'�ʹ��,�zՁ�r��7�#5J�)ȓ�Q�n+;�K��ug�}_}Iw�<X�|�]ֶ%�&ȉJ�h��N>��������3�͋M&��}���Y`0ǨRE)IEʰ=���������� =T���;���e���3X�gNti2�ZRp�%�\�f6�JHغ�\�H��n$�ˢ�9h�`��qR���^�S��:r:NE`wri�������g�s޺�3�5_�H��+lNA9*j��*h�>�,�v՞m��7'yX�,n���nS��T����}"��r����	��#����'R�+�n=�?���~8{k�>ݵ`BI�I'�VG�J�&�#nI<팏jϛ��QOI��w41�A���kzu<u�Z�J��	�N�$HV�n^�JY�nF�
�Pl.�'ob^������P�5�- t�6k;�mU������]�n{A�2����� iբ�%D�( ��7l�ZN	Y$�i`��7m��ɦ�k��*�B��:�ƗR�\��M��FgYp5c�n��FÅѮŢ����Ͼ����v�t��u�֔��U<�d�nzt�ky�*��f�A���ð�!TԩND�J�#qp��7&�wv��μ�`b�kbQ��l���p@z=����?�T��>��� xflIIjQ%9;�u`g^�;�4�;�4�8����m�Q���M�}�Z�� :=�����@u�<�)NBP���7��ɥ��ɥ��ɥ��{���3��q���=�"�f .�J� ��\��稜��K�QDdy��br
GN9J����������ν�`gri`wv7�i�JB9RJ���Ϸm_&�iG6�D��]v׋��Kt�����t�"$��#Ͼ�G�G���o�?�T��˷)�R���Ta�������������X׺�f�NF��I�*(���T}�������ߟ�ʥ洬�ؖ����;Jsq*�.jnqM�B�XrN���B��K�v���*@>�-���`���vw�F�۔�NS�7q������`����!�f�ef쨚��3�,ۛjĩ&�i� Z��K�&�֓_%��ȫ���ܜ�37R�' �t㔡,nmՁ�ɥ��y��������mm4ԥ!�&�� H� ��G�@z8� ?���3�����ԯ+��gh��zwG�}��;+�mu�^y%�km[�}�}��1����G��@>{����T���f�R�9r$����������X�۫:�U��٪H�r��:$�h��qR���@t{���RE�HP�,?W�UKs��X]�]������ܯ �T��2�}�}S_j��,�ѭ�m�P�+7w7i ��G�@z=�������ҳ�!Q��N�D�#7V4�tN����m��m;��n�m�F��i�iC�#��\=�Ł�ɥ��ݺ�3�5X�ԕ�9#��ㅁ�ɢ���@t{�]�>ܻ������r��8X��Ձ�y����������ը5�����r��29\qϭ���`�}"��X�e�m9r$���������������ϧ6,P�+p�i�~�+b��T��b���2�-<�q���gQ�+�;����n�q�aduUrq"F��Y�dv�6�"�X�Չ& .*� \Yk�.�Od��M;%�ѹ�M�q�s��[�\<�:
+��(��QH��×g�I���]���^\
\u��#�щʽ'R���C�[�t�FxP�f%�[�Krn{1�Rh�t<7HV�-�����nRx9�bsI���V�KW�0��J���&�*t=p�^�N������d�荪^�Γ�D�ml�) ��I��(�:w'���K:�W��͞,ڼzD��F�f��{�r�����.��"MJP�GrU��y�������������X�K^��BP�8���XnV�ە���nڰ��J7+�X��J؜��ӎTq������}"���� �gC&^�xn�.'���j�����t@����U�MV�ݘ87��|O�ȗ�꡷�m����`�cv�}��<�X����R[��kz�V��ʻ��~�s�B�%1�����!�o�� �EH\��/kjH��!�H��M,�M,��ՁŹ���l��r���r�ns� H� �$�G�@�2fݩ"�T�
���ݺ�3�uXܚXܚXf��)T�����S:�IO��jѠ�l���v^֎�Bz9&1(%Q��(J�9*�ν�`wri`wri`gwn�u��H�!(t�t����� H� �$�G.�ay �t�p�;�4�9�4�6�ң��$�^�`�BQ��)���l�:#р��3tP�wBhµ�43	��(�,�`Zֵ�l�]��؂b��$�HB�@��t�
�����@0e>�!�H����0�*Y�_E!@��l�̈́E��$̔ L2���ZS	��$!IR_RN!"&'�T�A�]�!����p6:\}Nbg��pP����)��G����3���Owѥ�i�JH���N���UW�E���'ր|�G�@H����܎A�*�Àn=�3�4�9�4�9�4�6�����j*dn$݋b��\��x�J����V�ɩrvw0�v���T�"	N!���M,nM,nM?Wn=�=���9M��9E��G =� ���_~��H+=��RE�R'*��x�c��|�G =1�sl�ͫ�h�ܼݤ�r����uKJ��y�`��������u��^#��ԑ�r+7&��w��W �o����V�{�0�%%)%Δ��,�u��ӭ��-D*)�Wm�p�[l��IxfDJi�)8�G8}���3sn���^� ��x�7=^�����ʏv�i��K����}h�o����l�Wuw"���J��|�װ@z8� ㊐��/kkww6�)�E������smX���?���?m��7����8�7a*R����qR� c��q����*��{��������<r�%�h�\p���+Օ��4�����k��+R���؂�mۛ�vX��]���ð��,�l��s�nݗ+�v�1���[�Qv�� 1���l��m1`���<��Y]εΧ�B�Z;Z����cRFє��6݉�`�
�V����ݷ7}W+j��:���R���+dnq��sȽX��U���j�[�l�fl�f���u?���o�y{wZE݌��v�:e��8�׮r%�u�:ӛ(-�W	�#Qm�g/K�����T�}�Zǰ@z8�;��&�(JJDܕ`g^j�}���,�}u`f��X�K^��BP�"Q5Q`f�i`~��V4�Q�֬��+{�)M=b��RT�,nmՀ㊐��@8���%e��^��mnn�� qR�9h������z��d�F������)8O�$�z��:��}L�v�/��^�,�M{$�RL�����HI$���~��ܚX�۫76��7�kJT��r��D7���nuQ�S�@A��I�G�>���UW��-�*@w��H_I��/$r����)D�`w��VnmՁ�y���ɥ�i��D��F�ʊ�� qR�9h����U��y��ܥ	IH�p��|��M,nmՁ�ɥ�着�)׷�H*RM��#L���Wd���غ4��T��&qת��r�h�G�!(N�T���{6x�9T�����#p�U���{�Yy���G '=��9h	�a|���f������ʎE%X͞9W����/�O�������j�r�OoWŁݽj�����j�5#R������������XܚX��=iJ��&��H��M��}��9���'3e`f��w39n}Pvi����$��k�R��=a,exZ�l<�i������m�T�����'=� ��7m)"�jT�'*�����μ�`ori`ssn��J��r�NU����`��qR� =�w2�n�Fa�uy�h����#��Fo�4�|'�W_�y�3�}��yMDI4�p�9��V��}��pǾVnM,V�5%�:l�;m#U8ͅ]Vh�dRQݭWi�+u��dVt�J(4Jhr�#�"D�p������lX�Zs�>�,���?��]�5�n���^��� {s� {u�UT�g�Kȕ*9MJ�$��ߦ� ;��ꪻ�O� :��b�9z�9R���%G�������ͺ�3�5X�4�
�,ؒ�(&�J�)�*@W��}~}7�����}_|kM��!I�\�t'i�#�-�:�lq�p�x�<�G����y�J��Λ�Mй�����ɻ..ݰOlq�1��4̬�yl�(��^��c��WS�㮻(&㭆jZz�������u���zȄ�=97[p�+�2j�͕-^��@b�`��k%u"dIึ����Z���(���:�Cl�Gls7��3!B�����" &�I�U�&�6�Z�< ~UC�3�_k3Fo5�k[�n�:�\��ѺcF�K�sh͕��+-�Wg\���:��n!7)JDQ9]���3ri`sri���\A��]XƗ��)�J�۫��@8�G�@8��r���#���2騉#��Q������͵g�M��7'z,�,�J�T��$�S�"p�3sn���VnM,nM,֑��^����	��������U>���w�~�� �������΂��7#uӣ��[��)O��:I���)5�M]���'=����� ���{*&�)���R���,ە��n�x��)�*���$����,��������4%$PMET��V�����N�Y��vmq`go]Xܕ��&�)B��'*�μ�`8�G qRݗs&�^nE�n�^n�ǰ@z8�9���?���zm6��2:�bR	'�$EF��<���`{uW+<W��i���m�������H�#��Q�����������μ�`ori`gt��9D��r�RU��{�r������vL?����HH��8��+{�K6���PA�&�D��"~EaO �}����z~,��Z�R��Q�6������A�}�O�/7�:NT��n�Q��`gsn��M,-�v�&��׵�	')�t'�]9���Ҝ�H�df��b��� 㮵�;2��}���IIR�J��?o�����19��T����f�y�W�i�TD�`~�͛�M$�Ԅ�Jd���X��76���ZZ�6�d�:�&�q �� <�T���}>T���@{M٘�1PUTJ��b��i��9�����U�}�u���`BdQ��~M8i��	5������yT��SH���ͭ�ݤ�*@zۘ�q�y�V�Ű�JN�J1��1�1,l�z��Q���	�Wn�[�h�L
�i������:��H��ջ�`f����f�UUS_�4����� �� �*U5T�&����@8���~�:O� '��H[s[���!)��	���ͺ�7�4�8�5�ܚX��RE�UAJ��$�������7zlܭ,?W�K���X�Z��NAJJ�)�fl�ͷٿ��ޥ@}�e���
����
���������� 
��� *��� U��@�������� �H� Ĉ�H� Ш0� ��( � �)"���� U�� U�� �+� �+���� �+�tTW�PQ_��
���@E� U�`�������(+$�k=�\@�6�0
 ?��d��-?�
   @ +l              �I)@
"*HUD"�P  �� TJR� ��T( � A@ H �@
@H,    4
  � �2+/yNO.�{�w�]�n�e�{�>�{�_n9�z��n{��Ξ��}���x S:鸵*��� ���Ϸ�\����O.�׳ɯ[�8��xzp ��w��x�֜�\��� �    H$�����rｻO.����ɮ�� ==��s�vۓ��Ϸ���av������s����3O Y�y��\���� Y�Z\Y���i͸���� ����7�5s۞��tﻼ��[� ��   �P� q����K�y�����=z���r��{�O����@  O��P q r{��x8 ��i@�  )k  ��:" 73�M R�P3� w �` "��(�gM4 ;� (   J����h3�:q��� 
M�:Q�� �� d
 ���� t` -�.>�=��&� !�oJ������ �yK;z��>[���;�����8 z}����^���}[D��@0q@   B��,` {�X��wv�k��Ξ���>��� Ξ�9�.�Z��n^���8:��Ӟ�[�����ۼ� 7O��������� �=*��iqo���r������ G���.���C�oy�����>�ת� z�)�*T @����iR�� )��T�mJ@ ��UI1(0� *�Jx�)P  !�*#FA���������Z����3��g{���w�?Ҫ*+��_�*��������*����UEE�U��(*)�G���0���@��A�jB	(0d5���#d0�'�+�?�&���g#��V\����Ь�!�$5���!�̱!"@�B2�G�%���K!	���w���x2��D��	Yk%���F\*��I���޴J��U*����!"A��	>+I�)&X�Ot��� �����y�#�K��3�8���%ɰ�w8g���S4!LД��.1���HT���+ �#�\�>)�� T��^J���4%0<A�6����H?)��E�h�h0H%R
U������ ���
�J�<ZJ0X��74�0a���!�D	<5�
z���$bFF a�ub��uL���� _p�QĂ�0�1�:/ �s���h$P�<ό��=��s�懣/Dk����2|B��$
��!#E� �H�� ����Cjq��RI9B���J1Ia�K�Ł@ԍH8@�[�I]�9��Za�ŉ��	,<<��$痁(`P4� ����º��0�^r�iÄ)��!0��� P�
��BD�;�#2y���xyVR)�0��<>'���H���cRY8^z�JfӋ
F���B�K�xy���^<ˬ�j���wng��J}��%G�O���ҧ��0��ϩ.z���a�2�$���8���s��%�w~ _N_Jޓ��~�O�&�����7�=%�!X�B���!�M����nq�@����9$!xz��*F���I�y�����<�hĩ �Ni8bl+o<|'۬�}�F��!p���F��Q���8Gƞ>+��੥�y���{.�ĳ��2��B����%!"��U}�����օ)ۤ�VM������V��9`�8hAJ-��RA�ѯ�0�p�W �<��Ϥ��x2�rS �T$�Ƹ|}i����kV!��d��\5�b�\H�������'��6$L ����5c\S,j�H�h
���T�D�ą0�x��R�碌�D�))}�H}��xӏ��'�ą	!FP��Ŧ.ʾtn�i���S\�_Z*�N�K�B%a!L���<ć���Ng!t�䥔�.��\���>q�j�]QEH%EeU�Q_Yq�1\.@�T]�:��0��O.d��Ħe߼���`��瞜(F	�Ʀ]��������o0X����3ݶ�LxO6��6}��JX{�G	X�I|��a͙up8Յ%O|`Y_�]�5j@(�P>>�,�����#�"@d�Fg��}�/ "��A/��bF�M�ͯϠE���*T��O�,����Y4�(\�!,�OCOcd����XD���
i�஦��n��J(k�c!Lu���e�$J��:�F�`ă��B6R�	m �B+G?h�"B?0�F㱠�G����3I� ��C�B�pӢ�<a�ʜ<*F�0�i�pS�La������ fp�,.I�l����I)���G�7!CO/u� ��]�d<1��A���B�X�4�_#��1�p����)���s��H:�(N���`B�� E)����0Ӑ�a��i�>����8��N{>�>���.�Y
��q�k���7Ò�E�K��IH����C��n{��'���>1��p�f`C�0��jF�	�5��0�
0��a[��;	,�$4�.i��p'���8���HbNZ�J�XE�C�C}2"A"�O �e�d���v<#^�(��+�E��|`Bᒰy��@����j��c}d�LS��*�k�8��(� �� Hbj�H4%�4"E�Dx���п{��ȋ
x��`8�:�jF��2�Ƙ�
`��Ƙ6�4`�6���>�g�����n�@��+�"t�1�n���X[��g�������V%-X"�(@1W�!j`���
8��V* *�"�.��(��!$�hh�;�!  �qō�A�FA�" ��0�A1B � 1�Id-�
�(i	��>HB�C7Yk����
1�6e����@��B&S��F3�I2��0�D�Kif@�x�A���.BT�!���)ą1����y`D�̤x��0��]�l�00ͥaF,�	�,H���fR�`R���Lǖ�(���6I�
0e���#M!D��XT�%�Ip"�XSG��.FK�OIH��A��W�I�1��I�xy㬹���dfW$�����6�[�[�"h��}  C4o�.<5d��h�2�t�6���u!L�a�r�fa���6d�p�B��OO7�����$
oI�-$�%	!B˄�HԌ�� �I $,H�<t W�]0#|����8n㮼�ˡaR_4�
0 ��ŉ��i�%LXDсrMv	R["҄(I
:���Ah�4C���Rİ�s��#�$�$���(@�+I��@�Jp���!��"�F�����>>���a���K�$(c��,%JJVe���-���a<�04��i41Ni�@#��!�Rp��B0@�<x�� L��WزOx}
?;��԰��p7�夋��<$BH+�Iq�r��8s�q+L<	r@�0aLI���dI��@�C.�̹�9�B5�@�;Oi��kƾ�3J��ƌ��Bn�3pɖ祸k��ː8����r�^0����)�)M�m��$b@�Ė�i3��o���!�f��0�!	t��2iO<��� C&�7��B&�&�=�q�#�K�y�*x�O#rK��.[x@��5kj���8&�Ё_	\e�bA.e�t�A �1�0ĉK]$���W��J���m4�sLR	�&&�d�I��,��^Á���F�ȅ�GCV�0�a@���Y��d#��7,$m��i,�����d��$s$��g�й���
����) Y��w�*Bw��Z]]�\�躈J�8��K��C�	J1@� 0"� ��B�1u� m��b��m2�#A�a�F@����j���, ��D�
���$k���y�����E)2v���C@�C&<�Y	2#�paCBa�$}X�05��%r@2��V����B̌�K"o(fR�m���"�2Aӕ��N!���ym�0u�E�b`o<�2!��y!	��#�y�y<W+�@���K[嬘��Q$����V���dV�����Heu��(*x��'Ǉ�z}2hD�},ٖ_�kl$E�H��H�B>�JdJvS:$�2(z�E�$HH��&jx0(a&ڕ���2�i��7*QІLe�H���]�f52[�͉2V�>����:��}�}~��w~���`?�= �b�  -� @  $   ��    Y����R66݀LK�m��R��C�S-nTh�� �W6�GI������UA�l9Z�{,�uI�p5URM''i�ҭF��Ev�J��� 94XK]	n�l��d���R�J�uSd�(�2m���e*@[N-�۶�^t�$�P6T���T�L�#�%C�QW.ԓ���6���<� �uͤ(e�����`���qo��ZB^���VUldP�� m�h��kh k   �cU@R�E�z�mکU&�V�$��̓ucm�	 �   9��   ��@ .ݛf���[I�Hs�9���Q&���am��� -� l�   H   m�s[�� �.�� �m�`�ni'Ll�p�5m֡ڥ@j��*���mp�?�W��@     l��	 @6�� u	���U�v��Z�V�nC�R�9zU�Ij�R�:#��ݪ4��Gh���i1 �d6�նm������� 6�۶��^�\��S�ݺl�FN�A^���U���v:n�m/K�tnӣd#h[`*��≕�F�[O,ͫ0e���!��T	UN�&�Z�b��� �5��:�U��]e�%�*�lm���p � �m6�� �` ��I��a�T��ԉ;m�D�D��k�.M6�^�s-I㣆�p[5ZJ'���y���a�`]��R�w�k���p 8u��s��  ��m��l���H $��~���K����H�p��[8�\5Qr�]:*W-�kGn�I���m��keV9��
�z�Β�׫!�N2��<���)Vڶ�aZWWK����m�� ���
�v��AU�+��W�����]-�\���l�$N�8[s��h�������G ��l c�N���Ԁ� %݈!�jyX8U��V��ݫ�'\/��
T���e3/}?:��U�=�<�M�vɐ��n mL�Px4ҭl�hI]56�oNh�8Y˶ I=��^�� 4Q' �`6�m�u�m�l��h  [%�n 6��n� $ <  �Zc�6ݒ[AT*հp�UJ�U�9 m�  6�  �`  ����� m���[VK���m�m�hm�M�M�`�  ]6 ��g����h����m� �� ����:�I�[t��-�m�L��h���E�	  H �l��� 	��$i   l 9 �� )m��  m���  Y,� i�}������ۯ ��am�  � �`p��$  �l  6�	 -���-   	 �l ۰�:H�6�  	3���K.m�H������ u�v�$  ݶ I��h  $-�lm��n�a�-6�i� �i[UPU�`JY�\�-L9͖����������ii�]6\��U_U�j��*���ڎ��%���*��6�Zs��  6�&#-��t���>����<�@�I���WN8��E�I|�:gI�u�\�:1�������Z� ���$  	�/���ڶH$  �I��� H   �mSf �[@-�-�m���bj�vl  ��ŴrAn�\H�` ��E��tH $�`-� ��   ��ڭ؛\��	;8����
Z��4���]"D���HGq�a��sq�1.�EϐV��i֥A�!5T�J6,8��ꪀv	�$�jO H$��m{�  Km�Ԇ��q�ӎ�Kpj���vāR
�4�u�Z������� m"���@�M���J sl��hm���  [l09��%\b��E@Uu*�@]@Z��(�V�5�=����$ h-�kn�[y��h�&�DD�Ӳ�r�UH@5UU*� d�$%KٖJqJ$6ٴ� H[Y-%P%-�U�Vw "���]0�j݀���If�R��qP{>z�%��a�j�"6ݢQm�N��[r�2J�e��ɢ�ӥ�5Hl	ںl �[Y-���ɶ�h�Ju���6�2[�m�bK�I��{ﾆI$�mm�� mj�� [��tp �2�v8�m�HN��� �M���ei��7 #�J���`��{kh�h�mp �zr� M���q�o[m� m5������>9�e�r��T�h��-�;a�i2� $ km%�,����.�V�� ԫj�8Hr!5C��16�V�d8C�����h�m l  6� ����]�VT)jɕ�ti�����n�lT-C��
�8�;vU@�����Ii�(K(j�t��7���L5��'Am�t��<�٢������|�D�V�mU��Nx��Mh�ȩ�608�ؘٕ�������>T��C��Z�t��iZP�0 $�eMu,�[�q�V�cR�vCp��mհn�   @�2J�ҳʪ�Q[]��ש�/<^P�X�>��#U]T�Ԯp
Q��M�fL�l��m��;l��� �`ͮI'��4���v�v�Y�UW�ۥZ��v��]�\�q&��)�o1�m���@  v� j�l�=w��}-6��   �-�k5�^��8  $��G�u�m�&�of�l�� A�h   �` �`n�[@ H �:8��]i��l#��i1�l�j��f�j�zVvZBA�  KL�[n  xllm�m�k�}���od풱�b@�cm�d���&��8r�Ӗ� �  �  -��    ��p &� � �mm8$!mv�z��kmm�Ym�m&$h  h�   D����  p6��    $ h �   �p �  8$�j��(�� [@h h  *�d����T�;,��j��24jj�������
V�\�z��gCr�-�m�[v� m���[Im�v�� p�%Q�ؐ6���-�6�X8��rCl���[@m� n�-�	V��ݵ:j�\��u�m  �  $ � ���9� 	޻�֛   n�Ԁp�` m&m�[@�a � �Xg8.�  6�  �� ���`m��6�& �  ��  �   �  �)p $m� [Cl�m����k� ��n���[,��h��A��J,�U x����������C��Y$�5J���YL�Z� ��hh[M����  m�Yp8�D�6�I �#�ͻ`X�������"@H6܃` �kh   �G6� 	I%�� �[$��u�ր�  �;m��: }��  �f��	���[� @ �` �  �  �	 [W�� m�f�p/Z 9mY/U��4����d���_�)`��-,�s �[-�����4�T�U�l�J�Ҷ݂�m�I�    -�ޢA�yn��jK'm -� ��l�`�gvZ���iY㥶�SB�       �m�m �   h6�m��Ė� $   l  �� �      �t�8��6��˯_x� �a� �*[-UU�lim�4�d(巴�E���6��`r��r۴�[d� CIs&����� �  �       ��p �l�m���    p�#�l  m�z�l�&���� ��Z�I��צ�訤��j�j�f�.   -��7{��l� �5��*��R��	��*��Z�%Z�
A�3�.�t �P�-TP
�͖ (-�M�P.e%�l�g��q�}-a��e�5
�4�O��Tz{q��VV�clP���*+�R���(�J�R�+U!��p6�vJ��UP[@�]6vצki�\�R���檪��ԕ�E��Hm��@)��^��\C�v�:����*��z�<�s���E���� �&�����,�&�JO�}���Lݷ �l  rA����/ZH�`  �fٻI���Zm� m����R���iV�͗T����|�u�*�
m�N����5� [%�)��7J����X�Bۣ�$�U�M���K��u[n��!�  f]���T4��Q':����MA�%A	�/P��q`(9j"�
�? ��U���_<8��G�pEG�>�V���_x�OF�D"�)>>`�>+����A�#�"��
�A� ����u^
���<^�z�����T��@���s�@ǣ��|��k��g��� |�p�@@=,T"��!DE�!��W�W�~C�Z��ʇ��A�����x"�G�)��P ET�"�$H1����D�TG����*v���:�"�\"
�"�J`��P
�
�����f���@O�a���P:(���
��X��T>J��|� �t=E��$T}:?�:�|*���:qx'�'�����=@����=H|�����o�
�N�>��ĀDAz@E��tQ:��k@�A@<A|P��G��C�$�P�x(:����Ҟ����)��
|'����  u0����ꪊ�����A� ����;r�U��h
��&焈$�6c��q3ݲ��s����an�]����.t��R%�vI�t��͕j˰�`��8�89�ͦ���Y��,DgCml�p[���\͝���MU,&�Չٔ��POl�^[�ynt���:앵È����Gl���͙��:]��ci���p�Y1m'JZKRm��[X��&�b�9���9�p��k=s��
@���;3��	W��ހ��qٱ�{^��jFf#���<.�]U�:�P�	�خ5�m���jӝq�ղ�»u�S�Ybtӂ�������K�1"��GU+�dZގ��S8����/9�t��}Fu�۵n1^RP��N�e�ƕIf�ud�F���R�˶��j8�����U\]��\��m��.3"d�P�X&1�ѱ
���Wd�� t��^��vz��g�ݺ���i�]��ADA=N�C5-��cC�]���X���[Lj9�M1������ݔ��#Y�د�js�u׷���ǵC��r�ܛA�Lm�l[�Ѻ"y96�^x�GZ�#lG-L���--'d0�M��,ۊ��S��@n��`v�dG�:��TO3"���	��RDsn׭��z�Q��6��yط�Ol�g��"y��[t�V�h��yg����b@A�[v��Pm���'L��T��:�0\�*�m�OF�6�96�^8eV �3���Jў2��A�K]5R�r���Z����)kl��uĦIp*P6Z5=�.��[����p���+ݗ-��K8����]6�:�4�U�<���1����pm���t�ԫV˷;7E U�Ỳ/���mζɎ��UuC���E��l�;h�b���@[�Q��X�]5�#L�V��s����+�Ac�C�����ƴd��X.��>�:4�ڄ����Xj��㧧-��mĳ�-�wk��l7E ��<¦��vA�1[�m��h
�|� ?�S�(��� !E_(����⯣�O@i��`����7b���=I������ƯY�]��ʸn4S��2�PVY�fBw=�ě��g��g��])��2ԩ�zi:t����)zrL�2E�4gAN���,��E�N������ܗd��ǹxd[azwZr6�մع��V�tt�/k���S�$8ŏ��X�b�ݜ��%�X��;�o>�:�sv\�,����ݴ�Ȉ,S�
�*_w<�	�3
L�ɐ�ٖ�e3�0d��O.90���v�,Hn�M�'N�b�عTp�wo]X��0;�s����>���f́����i���)mSL�s1ޥ
!v!B�=�yXZ��`vl����)�Jq�JN9J$�;�2��+�g��,�q$�n5%E`ec�H�l@���""^ݹ@nVӸ. #�qRR+�g��,Ǽ��}����\�NTB�����T��q�i]���zںN �"�mz��QY��tB�I���3;���������X�8�7_!�	�T�HGrXN��v��� `�%\Q �P��w��3�o$�w���gt�>ַ�JH�n��t܅���ܠm� f7h�l@<��.G$C�$L��Vf�/��zXޞ,�r�;�uZ%H4��IDi��3�DG�kt���ܠ5�P���ߓ�yu�\�\���=�����l���Lm\A�M�qն��`��2���lU]�5���ܠ5�P�3���IQ��n7"�
B���ܬ�� ��v�-~���$n=}))	�ӧ*e��3;����vJI&�Dh�b�T+)P�'��b�B����:�Y�`w�d�D�HeIR'��fwK{gV>�`ol���|��'R%!i�`ol���ܠ5� f7h��#���)B�mč�4�Rl�f��73����n^*�&ϧtu�wt#k��G��U��7k���Z�����؀�iuuJNF�H�I#�7���ߒ�Ԁ|�e7t���p���*j�Kh��Ձ��r��^lT(�����G`w��Vg%:�N6IR
O�q�μ,r�X���(�U	z#����'�?�<�y���g$���J�ēq��Rc����P����������OHPM�T��^k��3�3�svݛn��i	�gW��<�I;��s3��cl:����m������� �m���Gސݮ��]>�)�*E��[��͜X��KAٽu`w=C�����D� m��M���n�u/��U5U%4�-�
(Q������Ձ�;��ٳ�����)9i�M�����w-X	Gk����zY'��{y$�S�@�#��ΪQbń��c����ԝ4;.gY����v	��*���w \ubh��N�}Z��k�'^fGlK�]!Ȧ���vJ9�Mt�Mh�Ol��u��Q������:�n-��<LC;��/)]��#�䣳�c<���),n�rn�&�if$��Rd��؏B-V{g6�������k��P�Filt��,���Er����@7��8����Ѻ;4��I��y�wq��ٷM���lsЩ�ɍ��y�ygt�["�i��K�m�"R��J%:�i��%rV���:@=�b2��DDG�6���m�)��	RP�vn�/��7_��o�u`b��`v���M��R!H 3)�@<mB'�ݶ 76�&�	5#�$�VguՁ�;������aDO8�&��
��Զ��m777w�n�v؀̦� ��w{��ߟ��.���X`�]L'O;�ح���Z����N��;X��*%��gu��"q����1�+����ŝ���r�)#i��jp�3r����BpЈDG�TN|���뀧�3����'�����wﷳ�H�iuuJNF���
nE`vw]X����8�3r�75uN�q$�C)�a�
{]ݫs�9Y�`fw]Xw%:�l�(�H4�;vp�ﾯ���7S��;;� cv�3[���S�%���SmH%nPۛ�p\�t�8���ږ��Cc���e�f%X�̭r�xڄ�n�v؀��])� i�Q%"�;;��߿$���=�<X�yXk��)IGD��ڰ����^N�	A	Dr��PAOx��g<��~���V�>�8ʑ)8'%����������w]X��,�.�Ғ&��uWWr�̭r��6� {�ek���>���fjӔjjy����j痙�7�!nr0��]䂓6ivݴ��fi�.�Æ�wZj6�)��fw]X��,Ǽ�Ǽ��]Eө�ID�`cv��V�@fV�@{5�]G�&wLߪ!��$89,��Vc�Vٽu`gt��}R8��qȤ	$�lB��IBIW{y�`w����f>I��"r��U�5��J�\�Vݱt����r�JE`}�� :#����O��Z���ݹ
ڞ�6-Ѫ�3�����N�e�����>����6pkl�Juj�QнU������(ek��Z�θ�M����S%�`}��M�$�(QFk�+s�u`f��>\��JH�I��*�P��(f�ٮ��֬֗WT��i�����Vٽu`���r�����"}��P�\
*$�S��9*�>��`{�l�/��y�`}��T$�
u$BGng�h��aX^3�k��7����@케lsǛ��ѫ����ひv�ϧD�Z�Mڸq����v�g�e�
�ۊ��1�|��6�Og�)sV)����U`��F�Y�NsK�kn�K���gt/�O�0�!O!�V��bd�W������ণm��]j�,ktg^0���]���ln�l1Sau���6�ԂTs�p68vz�oJ6Դ5���%�Ȱ���URT�Z�}O�H�3���85�S�q��Q�gm��s������H:p�p������>�� �7��ws��G#�H�.�P��(f�ٮ���*����H�غSn ��ܨ��X��V�;��DBJg��ٰ9�͛���&��:%H��U�}�����>Ǽ��z����>%BD� ����Z�ѻo��f�� {��:;�I�(1T��6�j���m���\��ێ�W���c�K7�����6x�\4-f�@fV�@{6؀=��D}��}(֗��)9q&�)���l����K�G�D��h�nP��P�\
*.p)�B��}��������T�c�Vf�,����'$�5Whek�ek��m��ݠ��H�JH��85!`f=�`{���^ָ�ou�m��w��7P]V����=��/3O�,��ri;+�3�F�J�m���@Q������wͶ�7h�l#���ek���������CM˗L����R�2oq�`w���͜X�����8'%��~��I=�>���*�a+
��tm� �e!	V�ZZ��-o�=ʃ����J�$bj�H�1���;��̘�`�B&�0׀�H\�#���0��Cy!&��qb��X"�����dlm�xA���UeXѐdIIe���%ZT�YF@�1�������H;��	$�k*6�V�%d��Z�0�!+F����=Y2(�BB��)
"@�b�(B�	�d�0@�,F��-!!�E!U���� � 'E�]��~�8��0��}��pWO@�"��J�pTH�Q��}��߷���{�o<@-������Rn���R�a�Q=�͛{�MID} s��Ϣ!D���[��Ł���Z��n���S�aBHn�~{�K�Q	L�����
!L�q�`w��:�G����������G\X����*��Z���t�;�[Q�îգÔ��]�z�V
�D�L��$�C��;�Qܽ>��ٳa(���=,>�P��vf�T�:UM�I�T�v���
<�$��̭���%3����9�ש(I/��l$�=^�&���nhm�r�a�JD�=��DB���z|��6I)��=,n9֦��TT��j���������%2��>P�or��&c�B�Iv"?�MtT~T{��|�~���A�{k'SR�Cr��M�,�)�w_�dG>Q�zCv�J}/m��D��_�ҽ�J��ga�s�icm�k��'F�!t���#�cNԺ��Ir�th�����l����@{v�O��w�:d��uOqq2F���$�(�π�}�g��w��7ޖ��,<�b^�TC�9qER9(ϔ.���F�2����(�]Eӧ
nT��������,Ǽ������I�M��M]�5��Z��Z�9�փo{��wo�߻��?��s4�V��N%�%hs�YnV/n|C6�%����1��<�ns]��
�ҒIq:���k<'��86��q�d�0�c<;f��fn4h����s��$b*O2���G1��]r>�Yr#9�[-,�&�-����l`��X��\p��[��g]�cl�. Q���WD[n�Vݶt�#��tn2���<Z6ͷt�6��K�i1���:��7�/)Z�T-Uۊ[�n�x޳v���>��ZY��gK-R-��4X/a4R~I�	O���l��Z���wu�/��DD���,�E�I�cC��N+���I��ou��;��v�J6�z.&ID�%H�rU���zX�=���V{�u`otO�H��Dd$��׶�ek��jWEVou��]�R�7#q�HX�yX緯�� 7���������6t��NR(䙃 �Rٲ��N��F6��nۓ�u5a��H�u(�䎤j&�G�ٳ� �7�����Hs��6{���I�����.�͜�O=����' b���zX������Uݙu�M9M��n�RK����������7��z׾�;��`fc��B�m:ں�<m>�Ͷ f�@<�bܹI�CN0i8�͜Xٽ,͜Xc�V�W�������� �nF�Z����t��	'��qְ[^�$�E>�R�)%�J�&䯀3{����Ł�=�`oo]X���~��LtM����@fV�@k֡ {�s]ĥ$n���jB��{���޳�D�@��τ�s��̟s�X��X�.��S�:��ک$V/j؀=��^��ܠ=��E�M�.�T�K�X9��Q�y���ń����؈K�ي��55X��h�f��g�Q�W7=�Sѵq��Vc�$��"��q
:R�REI�'�{_yX�yX�8���X�:�d@�*8F���3r�7�q`����{����.����$�JE`vl��>��`ol���{���:.�I�Q@%H�n�wK{gc�V]�U��>��~���3��-�� 塪&����؀���>^���@?��/ȥ
q�6`�Ҩ^Λ�p�e�:��QW�ڒ6ɳ۴�Ն�l�R��Zn��@fV�@k�b �7h{l@n4���NH�(�?I"�7�q`gt�7�q`f=�`}����ԃ�q%(Q��>��`v=�cK1�+�ga�G�Q�`�H�4�7�q`g+�6s��3��3��1�N(�Vc�Vf�,��c�V[ܸm�rA2��M�2%8ᱛ�X�g��;5�)�v�s٦H�[J΅.�(�帡�˸*������nI�&��m��$ x{���#g���7Z��8�Eʗ=V��=I`���3�ƶ��Q�r�m�P=�u��]v�/Kӭ�i��s�c�.�t��َ.{Nb6�1�Y�bs;��W�p�(�G���<<�ϷƦ��x]q���]���ﯯ�П�<�Hj��Ϩ��!�%n`ۛ��۷S����l��g���up��.�r6���@�� �����Hn��@kw=9*(D��6�`gt�UU${_yX���͜X�֤"��Q)���@<�r�̦� �m�1�@5˸t���$�jB��}����ŀfwK{gcK���䎢�S��ܠ5� f7hz� 3)�@���qR����9�񧓊y�wTt8�w.Ԁ̥׎�]΋��Vu�ؘ@��q��ܠ1� �s.�It�*lRU7`w�����
B�W�U������v�I�og 3;�����J��$T�Q�9VcnP�؎��w��{� =�c��� �mȢN+;g��,��W���g�����
IQB$�I�) f7h{ˏ�]ҀǭB�k��=\���0AqD'wc��6:�k�tn�9�X���5�Nqn\V+a�b5�swh�l@fSr�ǭB �n�Z�)#p��!`f>�~���7�� �����Ӌ�˫�R���Q	�ḿ��Z�s1�IE�|�&��_N,׼����]:�d��%wp�3�� 3)�@c֡ ���(�S�NB�ܖ�N,�ܬ�Xgt��z8�)��r%E���궗 �Hm��&.�l�s�{tF�`&{*�2)*J��%ENH�$,�ܬ�Xgt�7:q`}����ƣ��n��m�1�@n;b2����t�H�(D��6�`�����ŞKu����t�`}�NR�qR�Ȓ�����nP�؁}1}����؈Q��o�vg����T��m�Se��Vd���,�����;�8�>�R��rT�CqG#t�M�{W�^���zqgrX� M���\�,Y{i{,���{ގ!T5T8m���=,��vy�(��(3+ޛ�l��6*l�T�e�s����yEQ����̯zlg^�&���pht�A�`v�x�3t�个���`��;޼M��m9T۩e��'�{�`wq�`�c��D(����,��MS �u.�:���Ƕ�D};������̦�p��z��!�jB���`1>��>�##!!%-�
�#�@���2ʏ�c����j,D��#H�1D��@LT��"���a������	���"O'@����	WR$$HH�F,y�!��tB,�t E�}��$aE,L-P���>��	�PM�� �@t���F�Ƒ��T�,�B`�,��H2�$B=O1�Faa�@t �'�0� �DR,$ �`1"A A�	! �$H�$c	�F$S���:(@"�$=%����� l[@,mKQ�Mr{F3�g$�<��Prq����)�;��CZ���ZM��������^@�lڳ��1�8���d�����h�[H\�5�P�&�S8�,�����G[16��p$�����4��%6хMї��]'�E����;���Ut	��p]�h�f�F:I2�ס�+;��@uӧ�]m���z7X.�.�G,��u�o(��p���9_�����<��s�v�������,��n���J���ōH�  �+�D:���c����@���pmm�!��h
6
�Sv��TxA��U�j��%Q�Au���T �l�e��*�`����F� ����:�2ҍ����3<�[o	
�vM���3�Q�ev�5s��=Wr�a�UBNQ����t�cg]�ks�4*)GM���1��O�M�����q���2��k��d�V݃d�ܙ�n$�瓎�����0��s�\�i#;v��/bu��C8�nF/V��V���5U.z}�bZ���m\��4�v�>mľ<��7�<m�彽tn�ԨN1��OLh������@�دj��A�R���ˉ僁Zq���V�jl�)3�Iˤ4����U���l����x�@�0��l�才%��6�F�R�m�r����cY6d��5FE 
�v�^�s*�QƳɀmu �/be`8g��r���ّT�]�rm��'�F��(���.�`(	���ꪫT�ʼ�V�	�+n��]l��М�Q��!��rʙ㛶�8*{\^���6�oHr�M6k�9Tjay���F�La�s˺Q]�*L���JR��;& k*������Ď��elH�;iu���M�0]�3U@[�Q�Uc!]W���?)�M�n[&l�Rga��@��.�Mٗ74����e���r�z����(3��^�ݝm��������͖��.#��>��R��CN�XB�v$A�Q�Oq��D(�`���U�x�T<DO�!��D����)���.]ۀ�ϱ���ڟ����+ɻ�;� q�a3���QZ��]9ʷnΣ.ڨ#^�]&k4�ż�$j\䝧9f�|�:��u��	P�X�[�NC��h�ω�=I�n�1��n�:Ƈֺ˹��m�C�g�����uvW[d�h�ju�N)6M��mۀ���;��[1z��X'��p� ���÷�\[vfҸ��<�ȯFs,>=����ʐյ=8{Q�j��hq�zӵ�vԝ��Lu�]-�\��=a���v~G˱GQH��I� �����7:q`��b!/�;���3��Zji��S-2�m��</�!(�K�!6��3��X9��b!L�;;�)m�7.[�T:e�w����u�g�/B��3�v矋��ňi����Hԍ�a�=ܽ,��vy��3���d�-RlM�����cv��؈������zX�8�>ݏ��ԡJ�7$��$uy)ð�szҘ-�x�Q��U�鍝��w���B�EQ��>��ŀfwK;�G�{���z�M��r���5�$���ya�� x��v���h�l]}2f�:�j��Cn��݁�ǥ�s���DDL�����`}�J����I� �n��؀3�}�G���}<�JN"
"T���,3�X�8���`o>N�D8�#�JV����5i�uS��Ӎn�-qİ�`mq�oF�)#r(����,3�X�8�s1�!/�;��>��X����ܒ]ݠ5� f7h{l@���5uN�*H�S����fwK�ׅ�)P���Y߷]��ׅ��rQ���J�m��`ol��3;�������y�7vuIR~$��9#.�@ݫ{f�@����{����t��%k.��0\e�i��3FL8�N�o<1�F"�up��Q:���@c�b �n��؀3���t�H�*r��&�,3�Xv�,3�X�8�7:r����22r����ݣ&wn؀3����JH��9*I~�[��VoM,��v�"����|�zX�O���!#tF�r+sg��,�gc�VR��FۅJ���BF����++�EU��7�l�v��[��+;E(��B��%:j8Xgt�>�X��e|�vN,����܍�22UM�ew&�DD(S'{[�`gq�`������%I���G*7����sm�1�@yֹ@{+a�MU�8�j'���� ������������t�8�*r��&�,3� 3u��ܠ1�P��&"";�2��Th�?s�fO�]�0��\ܛZ�냺�?�7�O�nܹ��g"�VN,���,fL�])�]M.�sָ�sΌOOn�M��;�y�v����&]�e����h�b���������k��&scqp��Ӎq7%B���n��"Gɗv;<Bguv����o\���4.˜�gцV�τ�˕70EP9�@����mMq���D����6��k�-{�%��D(P�%���WU-��h�%;78��!3Y��Z듣A��l(���7���b�#t�A�I�3���1�+;z��>�;��`l��Tɦ�l2�̦�t}��Dɼ�B ���/�d�����S�܊��w��3�X�8�3r�>�WQt�B���T�� �����nPw����`g��~M9$���F��7:q`tDDn�t���cv�ͦ�꫐���t^�p^�����Fj��jVD�3l݌K�����]��pRl	mITπݮ�@c֡ f7}��DzA�_�kZ��Iˑ�SNlgrեң�(3=�`ny��9�̛��*���>h�t��je���Հf{���1�f�S=������]X�9J��D��T�����v���Z����\�)Kn���T�:e��+2l%���|�ޖ�N,�6t�5��)%�0��e�&{W-�#VS��-!�nc���XD�Y�)(��H�D���X��V��,ΜXc�V�j�.�HTtBR�������}�L�z�@f�t�1�]Xw%&���i�Q��,���Vd�p�*��v!%+ﻎ�X��;wgT�'�Ԁ���%X��X�֬��v���X�;�j�4軛�n��Z��n���@fV����������1�Z[qk�P[�bR%�nn�lֱ��v��rA��ݸ�fS����������n���@fV�@c֪����T�⊥B�RKs���̭r�ǭB �7k��铧���������p$�������޺���Fo�,�,���STꔺuD�����"=��qXs�vy�	�(Q�DF�3�l��:�T�*X1�MԶ��7h�j�ek�=� ?}G�)���u����=���Q�=7��1��n�U��R�FNE�o��>?�7"]*U������({l� f�Z�=M������Ձ�WrofN�=,��vy�j���*�mO����P�i�ɧ6{_� ����%䢫s޵`fV�l�Y8�-�r���ꪙa�"g7��{� 3+\�1�����'URڒX��V�~��;��;�������+�	s�t0�R��
��|�o��
��c8�y4��e��e��5/��o�$:�R1�g)!�a�qeg��;��3՛X���.��N��I:e��GXĸR��D�vR��v�Y�����>u�=�'�Ҝ97C�"���b:���Ͱ�i5n4[΍���\�)e����ݜ��L�m�Z6���X��ѭ�;��X��F9��9*ꈄ�vBX����*\�TZ��ոwM&�9�gd�\:�[����Δ�<�i�!E�K����S�Mx�͔=� cw���zA�r�K��r�mD܉Sr+;gꪪH3}��~�Cs޵`w��6y��Z�9R��JwSV cv��mB?D}3�O���Ł�rQ��9C� �NK~�UK��ЀݧҀǶ��D�ou�w��n
�L�Z�[V9]ɰ5(K������;��V�fl��8�-�SUs��TB��%n`ۛ���r!���jt��p1��n����������O�o;�̵�P���k6lf�։�HN�77r�l�y���bU�}U���	�w~�uߥ�m���:��������:�n���ڰ>�w&�%�EV{_� �o�����R��R	mL��i�r�Ƕ���h:#�{��@l�i��sT�ʪnlg^�������z�����|5'E"��o\e��W�ӽj��I��޶�d�t�L�){�����j��K�u4π9��`w���r��興�(��{_���˯�7$u)ӌM'%���u`f=�`fu�`s1ߒIyDDU���M�Tɑ�TKj�̭��μ,��gD$�IXF5HB����C-�E��78p��1 CU�!(b��@�^0T"O<D���<�ՂG�7����a�����~ՊQy��+d�XE#����k}�C�������T�_ �� 	�1 F� z(=S������A����D%�"#,���ݵ`gjs�0E��ꪥ���`���7;��Ǽ����Bq�T�7 ���{�}��{�v�J������Ϟ��G$�vJ�%,빹��V͎�:6{]��n{C)�vUmˊ����?#��f�b*�7-���Z�9��M�����	*�Q���O�<R��T���M\ 3+\�7v؀=��͵�>��\��%HHډ���VwO�3�^���޵`fV�l��"�cuA1w]�Ո�ݠ<�P�̭r�ޯ߫��]�`frQ�M�$���i'-�ڄn����� {���6��Nu$4Z[�ܳ�q[�6tgtf4�>IM���f�)�)�M�^W����P�l@���ڄږ�7 )ԩPPN+wg�wK�3�>틠'%ENr	�X��@y�r��̭r���bζ[DӪAT�m�z!O5�́��l��8���X�w���D�9N;�ek�}��<��h:�(
+�*΃?w=�,��nl�2�[�k����:���Q7f&:7�yF�v��-�s!pf��>6��X��ܹ2kg�(�l�s�X�� �OmZ�)���\��T��,�X8�цK�&i���G��m)�J�8u���׶Ș�2���k;���kc��b� H����/#i��`.�^d�^x
pk����RL�WGk�z�Y���u���rn�+<Oi:=���{��~?�f��e���ܙ���y�꬛�N#��M�n͸����9��7����a"nD����z�wK�{���{���事�	RQMG �;��Fs��Ǽ�͜Xڣ:���D�q�'%��>�`f=�`n���>��`n�꒤�9(U�9*���@n� {5�͵�-��XU�œd��wm�ٮ�m�@{���)$�8$�(�)H�2K���4c.qX�����_6��v���kP��+a���
��j��k�@y���r��޺�>童	��
�H����u�(�� ~T`�t�'s?{y$����Xٽ,{�t��Д��&�Xek��ٮ�m�@d�Q�l#�*nEa��z� }����vT�y�����u �`�)B7%X�]�<�P��V�@n�P���uH��j��#�rW'<�3Þ���J�e��!�f˛�v�ޡu�Y��
�`�mB�Z���B �k��f��I�rP�)C����+wz��>��`}��Vc]ԛ�QQ�GN	�`}����$�߻�� �TJj ��BB�J&�U�ݵ`fWvl�b�	�Q2&���U�}���������+wz������'�S�Wh6� =��P�� f�@\}���W6�V�W��׍Xp���i�GWi�}N�c���n�+<T��닪���fֹ@n�P�=��=!�ܡ����G)Ӄ���V�7w����h6�w�3i��;��(�*ꉛ����� {5�͵ek��ˣSe6�ӗ3-�����w~V;Y�`w��V
$(�JQ����o\�74�RT�5%��9*���@n�P�=��͵�t
�'M�R^�r&��4�é�L���N���x�clS Wv���b��o���ϝ��ݠ<�Q�zCv�J9�����Zpm�
IV�wK�����{���޺�>틥	�ڊ�!R)%��w\ 3+\�7v؀=��˖ʒ��Iԧ)�*��{����ŀ}�������Z��T��:pq�Ԋ���ŀ}��>��Vܮ��
"���?��:>��a�un�P�Rg���d;{v�t�{p��'���z�ò��o7GFa�$��cq^%��еj¸μZ��W%ο�z1�&�����m����p�S��4�OGY����b�ݲ�c�ɍcm�B�\����[WA�KQ�������˔-���G\X���.���06'a�M��a��i1Ϙ�9=���"M͞.�D�{3<��?=�q�����zy�y��8�t�(jV�g�)Яknz�s�Q:�ȥd$���.�I��m�wZ͵ek���܎*�jH�9R	9,������Fk�+��� �7����RT�Ғ�MJ�`{+\�7v؀=���B�Kp��EGN�����ŀ}�������5DD�6l�9�M�4ʦ���X�=���B�Z����wϝ~[��{�w��������g����kV�ԙú݅��d7���R���*����ߔ =��P�l@�v�k�p�$�*2R���`}�yZ�_����5
"��ǥ�}��`g3-X��pJ��N2��X�8��zY��������Vk�+���IJ�����]�6��r�{����GSr��r�rXwuՁ��o��6���h�]�~����P��,��ԝ����=[�e᱋�b�C�h�"rӎ;Ztv���d�_{��}������h6� �Wa]��"�7vq`f��>���{����.����H�p��zXfe�)DBIl(#��}�{6s�ݱt�8�D�I*D��*�{����}(ݶ �DL澴OOqR]�a	�6�Xc�V�wu��7�,�����z�q��J`��$&�].��j��jGd����\�<r3�+�o��|>|	R�����SR/������f�>���{���w5�*A�Ģ������_��J���Vr��`w�xX��:����J��I8�������ߪ�����Ž�`}��T�%5���૸A�����@6��5���!���G��w�$�{�gt�ݐn\�n[��������m|7vՁ�=�`n��R���"m��*:�sP�Q��%�'\n��=\v5vw��4^98sS��EN	���7���w]Xc�^�Hfc����h�uE&�[j�ӫ��}��&m>�n�@zs]/�'//xh�GIG%&�X���ݜY�I(���6�n�����)�M��-͇�'3/K��ڰ>��V���U,��V/y��4E)5,Nk��j��(ݶ 3�>���j@���#B!$H�c"�"&g�_�W�L�b�	.SG���r�'��1��_<>8�]P8J�B�,d*�, +>�� ]����+�i=)��V$I�� $@J{
�s�`�|⇑8�R�b��*1�H�HA $I0�U�$�
��2�!$&B�&Q)f( BJ'��A"�*J$�h�!@lE�,�`�`�"�@�H0$��l`H�d $OT�!Ib��|(��x:H�S�Gs�`� *��T�(U�%�뿘��m��[Gm�eF�`ŗ�Ӎ�.�SY�G����N��̶�:���s<�ڌJ�;Al�-m\�����t�g��"�z�v��@����s�t5��c�O�j��nNiݭaQ�X�v�:1`Q�
�9�8�-4�3"�wm�jq�p�,l���8�ڠj�3ً��6l�.[A�\+ζF3�qy뭣���z���j��ҾMt8;g�.u���Q��l����V4�K�䭲)��M�k+ZX���̒�g�^��J� ��q.�#�ǈsv�8�f
�v�z�\�&F��bFZ�,dD�m�Xr�H{*�[+j��U�X�'4YZ�۱OZ�=,m����;8��Z!�6����Y+n�I!��1�+r��^���b�z���Xt�U�+�1����7���I>����;1�"���N��q��1i���}>��-lv䨩y���%�{�#��W��*`����)�l��Ǉ�:Ԁ�ب�)I�+r��P�N�Һ��ӹ��6y��Z�(;�ձ-[�B��`�u)���滶��Y3�.�`; ]9�yW+�����K�![�Kns�[SW]<mZ�;r6�r�ᶓсxۤ�D��:�h
�k���2#箘�yɨZ4��e$)@j��V�R�]+;���N�Yg���5MQ������3�e]��OJFs���{@s#[��t���iVn$�2�)��=6�6l��Ee�-yj�U���$U]UU�m�xj�� �ƛY;"u��q��8��L���;�����)�P����V��ʩ�V���WfU�U�]m�S��On͓nlN�&��k� e*��� &G`��uG[R8��I��ٺR�Hh��k�����: �m�Κ�WJ�}�T�@6j��c����؛qåM���l��<1h]�j�bK���l�X�It�]v�'v��)�X�B��۟em����n�u;4���Sǀ��^"�JqQ����� D}}�����CD1>$�BKt�=�R%]#�Y�N�8���\�n:�]VM�5��$�v^37E�cb�8e܏��['m4�Q�3�F���E�m��6ݰ�r�n7��j��G$�*^q��,Y�&t[y�+���\<�и��ƶ�\��qv��A��
 }�Mg�ۗ��b�����[��8�	����C�IĦ�X�"�N�s��d�I��V����i���L�:�E�-q�M=��b��d�ۭ��ܧ8�uHmJ��;�n������|>��K��%H�q��z����7vq�ߔ$����Ձ��z�M��m���M��Z�����5�͵��G߾��(�=���SBn\�n[�w_��5�͵ek�ږ�j��R6ܲi͆���
y]ͫ�ݵ`}��M�����{�`sqδM:��s-����@f6��r�̦���t�~����/���N�r��K���k���5�9gv�H*(� <�����{�����T���)R�r����`f>�`|�y���V-]�*A�U%5?5"�3{y�*?� }� �N�2���`{��Vܮ�ߡD)���S�ԃ����N+�������Ku������`vr�]NH�q)*D����D};�ބ�>�e7(?G�9[�V�M��L�h�N
mX�w&���v���d�u 3P��sr�~���
�Z��wAQ�x������r�kX@]p�n5G�	
���ܢ��(�"�X��X�n������>�s��	��.�D�F�V�wK���#w޺�7_yX��_�RF{���c���NK~���y�}��5#������k���{����r�$��JS�)�5a�DB�Uܽ������>�q��uՁ�WpJ�r��n~jE`f>�`t澿�ܡ�r�=�4ʋ�*���x�n�G��\;�q1�L�;9�nâ�{ny�2[]Y�����m�����lfw]Xc�Vc�Vg(���nG��rX��W�H�}�`n�yX��;�(Q&�M��L�©8)�`s��69Y�f���������;���ܢ��(�"�X��Xٽ.I��I<�#�bB,H�$�|��^�_�+���������W�9(�49#�qXٽ,���Wrlr�&��DG�֪�c��S�l�&h�3��v,��˵�M�&�n;J�F��V)�BN���M7E&�[i���g�j���3r��zXs]�D�2$ӡ��j���ܛ��%TfW�6qL����o�u`b�����M��H���(ٮ��艜���}(ms|�MF�H�qXٽ,�������W�[���o�G��r���3Whcj��(��(���I����_�
�w��n�̚L�^��D�<�č$^Ӈ[)�ֵ�9�a�Vҳz��F��fŬ��B-Ƥe��'����^�\]��s�[[hgū���ʦ�^�&�#GB,s]I`ݍ�͓]�������4N�]�U浉^2�b.zڶ���#Ǝn���p���w/P+�n;���8L�3�,��ne4%�Ԏ��^��,n#WK��_U�7�<盛��e�6�f��--�enY�rީ�p�[[+X�+���eex�z�6��ImMRhk�7k}6ܮ����~���A���`{+k�K��Snf��������#�C7���� 3+�7�航=�>�M6�N���2ìu��h�j�}3�L�=�ܠ=�lTM4&SM��U~Y��U����`f>�`gt�>滈�$b�����2��`lBK�{��;��s��P�������3�.ɹ37s7w�<6����S���'�����n	�.*=m��V�Svf��wo �`�`�`��������lllo�~��|�����w�� �*�� �`�`������� � � � ���?����76f������ � � � �~��x ��<�����?N>A�������|�����o�ׂ��T "����,�37nfi��n̹��� � � � ����8 �����|�����o�ׂ�A�A�A�A�����A�666?�~��t�2ۺ\�Y����A�A�Q����|�����o�ׂ�A�A�A�A�����A�666?}�~�|����ﷹ�K��!sw.]˻x �~�߯ �`�`�`(�~��x ���?N>A���﷿� �`�`�`�?X�nI�f�\1N��+z�p9�����vw���J�d���t�F��I.:3Y�nm�A�6667��o �`�`�`������� � � � �����ت>� �`�`��w����A�A�A�BQ�˝MM7ClN�N��j��	666?}�~�|���b!�A� � �����A�666?w�� �`�`�`�}������?�Xdr6��s�Fۦ)m9�Se�J>%(�����ׂ�A�A�A�A�����A�6 � ��T��}T�A� �������lll~����� � � � ����I���.�5��x �B�߷���� � � � �~��x ���?N>A���﷿� �`�`�`������M7fnn�n�so �`�`�`�}������lllQ��?N>A���﷿� �`�`�`��������l�n�w������������j���ҡ�1C�S�,�h�+mZK�j��۵��	�sv���͓ve��>A�����ӂ�A�A�A�A������ � � � ����x*��߿o �`�`�`����~7M�-���5��8 �����|��!����o����A�A�A�A�w��x ���?N>@S�@ ����w�iw6BK���v���� � � � �����|������߷��A�A��o_�u�����u	�Dq����aL���q�`s�ܛ��H"!-K�_D$�s�l��s��m�t�nJ�I,͜X�_�gy|k���}�����뤤�jR�I��`ĝav�hI:�N��1[�/q�\���Eh�L���91�+�}��>��ꯐn��`g5��)H�s�r+�ɰ���s����ߢ!DB�$������	R6�R�I8�{��X�xY興S=�f́����̗&*��q�n����T�z�X���t�Ԣy�����K���>��n'"X�%����~7M�-���5��8�D�,K�;jr%�bX~A�R�w�����%�bX����q9ı,O}���O"X�%�PO��W�A�}ݻww�����x��³�q�k��Cӷ�����q]bd�e��^�g=e[d-m;�Jm�r���=hk)�Sjj�B2f^����]�0�nm��%��v��u:���gt�3ƪ��"W[q���X�k��_*���Z�4k�q<4��]��۷k`��ر1v��X��<C�����q�z�b7;k�u��\sõնL� ���w���ů�$v���-�]���4����6�^5�j����j�h0fc]��f۶h(=�7���{�����^'�,Kľ��q9ı,O}����I�L�bX����S�,K���yi.nsr���ۛx�D�,K�{���?�c�2%�������%�bX����S�,K����oȟʹS"X�~�]�3sfL͙�wq9ı,O��?N'�,KĿ}�ڜ�bX�'��{x�D�,K�sB����$/��`�m��aM\ݜO"X�%�~�;�9ı,O=���<�bX�%����Ȗ%��AB�s�.�)!I
H]*wB�e5-�sM���9ı,O=���<�bX�%����Ȗ%�b{����yı,K��ݩȖ%�btϾ�ܸf��^&�Fy���@�ƝҞ�Qs3��={Chz;(�?{�����������w�{�KĿ_߷�,K��߹���%�bX�ﳻC��L�bX����^=�����ow����Ӛ$f�{#Jr%�bX���;8�C �TU

�j/� c�L�b^����"X�%��w����%�bX����%���T¢��v�6�U2�j�83��Kı/{���"X�%����'�,�HdL�~��n'"X�%��r��_��$)!g^Sj[hAUC��wv�"X�%����'�,Kľ��q9ı,O}���O"X��*
7bo����9ı,N�~���\�&��˛��v�<�bX�%����Ȗ%�a�~��~�ObX�%�{���9ı,O=���<�bX�'�O�5�%��O�����Is��.�ш�q�D��,:'$1�q��o%����q1��lff�˻��D�,K������%�bX�ﳻS�,K����oȖ%�b_o{���bX�'���ͳww6f]ɺ\ݜO"X�%�~�;�9��,O~�߯Ȗ%�b_��ہ�'�2%�b}�y�q<�bX�'�/��a�晻m�2f���Kı<�{���%�bX����'"X�x{��B@�
N�0�$���0+`�¸y*`S�0��n��yɦ����ڃ�@�(&:���b�T�x�@�PqԉX���
␃E_��Ǭjʒ�
C�5߽��!a`B��X��/�A����(
���"�����Ǩ�z5�{�J���OE���O;�;8�D�,K��wjr%�bX��{��4ݙ�0ۦ�6�<�bY�"2&}{�q9ı,O��?N'�,Kľ��ڜ�bX�'��{x�D�,K=ߟ��NjX�>��oq��O}���O"X�%���*������Kı>��^'�,Kľ߻����oq��}�}���״���Ί����
�Y���7kAh��h{3[����q��n�͜O"X�%�}�;�9ı,O=�;8�D�,K�~��~DY�L�bX�}�~�O"X�%����ۦn�	0�4��ݩȖ%�by�����Kı/���'"X�%��wÉ�Kı/�gv�"~L��,O�w�����7n���ۻx�D�,K�{�q9ı,O}��O"X�%�}�;�9ı,O=���<�bX�'����m��F�w��7�߾�wn2'�w��Ȗ%�b_����"X�%���gȖ%�'�}`�A� �zg��x�Ȟ�{���Kı;ݽ��7wrm�i�]�8�D�,K��wjr%�bX�{���yı,K��w�,K��߻���%�bX���ϝ>>�E��%a2�vA�r6�[\F�S���'P3�C���iNf~�����&�3��d��Sؖ%�b}����O"X�%���;�9ı,O}��O"X�%�߷;jr%�bX��{��i�7r\ٙ�mͼO"X�%�}���r��DȖ'�w��Ȗ%�bw���ND�,K�w��O"9S"X����ۦnnf�fɤ˛���bX�'�w��Ȗ%�b}��mND��"{���x�D�,K�~�ND�,K����d�����wN'�,K?�X��~�9ı,O~�߯Ȗ%�b_o{���bX�2'�w��Ȗ%�b~��ۦnl��0�.ۛjr%�bX�{���yı,?�c�_߷Ȗ%�b}�xq<�bX�'�nv��Kı9�'O� /oe�9�ݷF
�:Z��^�]m�"��˞Mp�8K��N֚���X����ܻ��l��ָ�9cjx�4�K����yN`5�j��(��l��Pq7Rs��j�qsN8l��$�&s���n�1�Uon2:9 ����K�؍vv����IM��B���V3�pIg��Z��q]�G�XK<�;m�x��<�CmJN�\�k�F�uc�Y'\�O�?	E���2�f�6�f�f�p��S�F�KN�ݲ�`{ph�wb\�mn6Y+��>_�a��IS~������{��?���}܉bX�'���'�,K�������&D�,O~�߯Ȗ%�b}�r�4��f����ww�,K��߻���%�bX�}��S�,K����oȖ%�b_o{�����bX�9��#m�&��ڗM\/�RB���w?�ND�,K�w��O"X�2&D�_߷�,K������yı,Of^�atۦnۙ���S�,K?�D��~�x�D�,K�~�ND�,K�~�Ȗ%�b}��mND�,x���������N����7��b_o{���bX���^�����%�b~�w�T�Kı<�{���%��{������{$��-q�F�^�G�I�&�tvz�r�k=�m��ٶ�NE�f%��7p��2��'"X�%��wÉ�Kı>��eND�,K�w���V{"X�%������bX�'߿^~7M�73v[��sN'�,K��뽕9�Lqg�'��9�������Kı/��ۉȖ%�b{����yı,N�owL��I�a�]��*r%�bX�{���yı,K����Ȗ?�"}�xq<�bX�'ݻ�T�Kı=�ܽ�\�!����ۻx�D�,���3��ۉȖ%�b}�xq<�bX�'�]�Ȗ%��E��ݛ��
HRB�u��ji�O67Mۛ���bX�'���'�,K��Q�ݼ�*yı,O~�߯Ȗ%�b_o��ND�,K;�t��č���f�;=�c�e��Y�-H�L��mHyk�7d�.E���\�a,K��뽕9ı,O=���<�bX�%�����I�L�bX�ﻮ�|B�����N�JZr�73T�mʜ�bX�'��{x�D�,K�~��r%�bX��~��<�bX�'�]�0���*aQ
H]׵Z6S�4������%�bX���ۉȖ%�b_}����%�bX��w��"X�%����'�,K��{y&i76Ệ�	�wq9ĳ�2&}�oȖ%�b}ۿ�ND�,K�w��O"X�Њ!Wg5�+!I
HRB��ަ�j�f���ܗwx�D�,K߮�T�Kİ�G߹���{ı,K�����Kı/����yı,O�#>�����sq����.�*5������WnU�ȥ�k��q������_.fq��ts6T�%�bX�w��Ȗ%�b_o��ND�,K����'�,K��e�0��$)!I�ۜh�t�۪������%�bX���w�,Kľ��w��Kı=��eND�,K�w��O""TȖ'߷/�K��nl.f�ۛ���bX�%����'�,K��뽕9��"{���x�D�,K�~�ND�,K���fٻ��isM�3wx�D�,K��T�Kı<�{���%�bX����'"X�����A���"�x%�
{��p�!I
HRB�Wt�-9i�U=���S�,K�����'�,K���}~�O"X�%�~�����KĒ{/	�d)!I
H^QיU�&�W�1�<e��s�ڡ�x�nG7#x�.�f�.�U��k�35ؠ������{��7��?n'"X�%�}���Ȗ%�b}������M�bX�w���'�,K����O����{#O����oq���~��<�bX�'�]�Ȗ%�by�{�Ȗ%�b_o{����&`�'߿_�a�.f[p����H'{s��H$��>�S�I�K��w�,Kľ��w��Kı=��t���e���s6T�Kı<����Kı/���ND�,K����'�,K`�dޓ
�RB����wQ4�	�����7x�D�,K�{���Kı/����yı,O���S�,K�����'�,K���当�\�se�w\��L.���z��c9[n6�p�ڜ]i�7M���v%�K#����[��G'e�ՎxI��2]�l��j9'��̥��\�9�brm��j孜'X�t�'=�A����<v9��ű���\�$��[c 8n-@�/��D�=m���i�<����ɳ��I��y��۝3�g�m����QӋ����[1�fc��>�������z�������9�6;ٳ�F�P�fϊX�g�����ⅿ{��|�M6���1�m�.���$)!N��<�bX�'�]�Ȗ%�by�����Kı/���ND�,K���d�wl��3M�3wx�D�,K��T�Kı<�{���%�bX����'"X�%�}���ȟ���,O�_ߊ��M6ʦ�:d²���$.u��Ȗ%�b_o{���c���/�w��<�bX�'{w��Ȗ%�b{��gM�4��)�m���'�,K?	Cboo���r%�bX�����O"X�%���{*r%�bX�{���yı,N���ݳwn���L���Ȗ%�b_}����%�bX�}w��"X�%����'�,Kľ��q9ı����?6���L��2�M���� �Sg�v�]%�^�Ԗr�r�)T>����G��ή�g7mܛ����Kı?~��*r%�bX�{���yı,K��w�,Kľ{�w��Kı=��t���[�i�t�͕9ı,O=߻x�G��EO�v&ı/o?n'"X�%�}�����Kı>��eND�,K߷��%�������6�<�bX�%����Ȗ%�b_=����%����;ۿ�ND�,K߷��Ȗ%�b{���K��nl.f�ۻ���bY�O��߻��x�D�,K��ҧ"X�%���oȖ%�ّ3��ND�,K���d�wl��3M��wx�D�,K��T�Kİ�_������}ı,K������bX�%�߻��}oq������ڽ�ыFr���ָn��7;%cy��wZ�J򉹷$֔���3z�b�74�ٙ��͕9ı,O=߻x�D�,K�{���Kı/����yı,O���S�,K����Λfi���f���l�yı,K��w��r&D�/�w��<�bX�'{w��Ȗ%�by�y���%�bX���΄�5v^��������oq����Ȗ%�b}��ʜ�c��|��9�@�����8� z����?w�N'�,KĿ�����Kı=�o:n��Ywe�����Ȗ%�b{��ʜ�bX�'����O"X�%�}�wq9ı,K�wx�D�,����~WS\3t�=�7���%���gȖ%�a�?�w����{ı,K����'�,K��뽕9��{������~�F�6��@1N��+z��3�{)F�:��n�7n�INJ�S����ݻ36q<�bX�%�����Kı/����yı,O~��C��"dK������yı,O�n_Ɨ7M��eݻ�wq9ı,K�wx�C�c�2%��n��9ı,O~�?N'�,Kľ߻����T��,W5��4ۑ�M�r�[w����$v��S�,K��߹���%��ș�{�q9ı,K����O"X�B�B�	��M6ʦ�:d²��K�~�gȖ%�b_o��ND�,K����'�,KR?d.��I�d)!I
HY׵Zɚi�O,�6�͜O"X�%�}�wq9ı,K�wx�D�,K߮�T�Kı<��vq<�bX�'{/y�L˻.چ�W
���PΘ�ϳYz��hPsK�9����z5�<��<%O����o%�߻�O"X�%���{*r%�bX�{�;8�Y�L�bX���ۉȒB����7��ک%�&��[w��bX��w��"X�%��s���Kı/���'"X�%�|���ȟ�����{���k���k�n�ǎD�,K߻�Ӊ�Kı/���'"X�%�|���Ȗ%�b{��ʫ!I
HRB��"i�7M�2��Ȗ%���^��ND�,K��oȖ%�b{��ʜ�bX�̉������%�bX�~ܿ�.n�wi�v�����Kı/����yı,O~��S�,K�������Kı/���'"X�%� �+�p"KBԕ%%#P�T�B� �N�xB����b0)�
�M�a	m$��gۤ>���wQ�ւ&�����@T	B�#V0�@�$
�C4���N�<��߿r p[F�2�\�6�E������sl�=l�c�vj`��]�m��Pt���U�]�.���n]nЕp�e�ϑ�`�T:��nvKN�-���N%]+y���UUAN��2����;���ɹ"�+6ݰ��t�Vn4�k�c��C�����9`;Q,��Sb}st�s:`�rJ󭩜���Z�Xd�Z^�@��F� �ęB���8g�`�헬��l�q�ѮӠ��.�̭��>N+�%�u�w5*�����]�<�Z�!┭u梱��e�� ���[R�N�m�h��� yGb�[^����V�5�Aj��Q��M���=!���t�ڨƋ��=9M��8��T=;�T�g��;:%gH^)�G��D��\�Z�eYV�5X�C�մ�t��5�]�1��*c0�:��a' ��,�)NY�W��s��+M!T�h�]���&�"uxH��{��^��`�n|\F̒���3dL�WSmT��5qJ�izș��gS���w"U��[]-K��	���8ر�y'e��vs�sX�s�l9�GQ�T��XxY���ޫ8]ź�pj���M��Nˋi�Wn�p����櫖
��F.;z�l�@T��죱3��s��cy�q�p@ �=�ֳ��[Y@��j����Uݹۡ��g]US�*yZ���ү*qj�n%]��@��9eܪ�jK�q��"��{!]�)�Z�FzŹh)�YB̤<T��^wl�K�uU�n�۩��^v�;Յ{a�*Q�Y�v����7-���k[u>����!���j����JQ.R+1�ll�̍@Te�K�RY%n��zK� L��^Du� ����v�!��=l�g��n�rd_�D�(�h�Lv�a�c�'y:��Ų�ֵ�b��M�	�����I�L�v�,�p�ŭ�ڞ[\<�ҪWтq�T��b��mۧ��ܐ�q�\3[�w&Svٻwvd�� _D�hz�P�	�� �����w�j/(��Ec�>���(*�?*y罤�=&���,6�8���Dv܆�ɥ�m�s�]�a����A�M�������Y�ΔL�:�u�X����k�s�mź �璶MҚ���͘BY�0�Ln��8�����9]�ټ�ӫ�vXrc0U��u�U�e��m�[g����T�Iζ�g�f��Fy�-����ծJF�NS��c��r��^.Mѝ�1l�������w�u���?Z�a�抦��\gP�#Q���8�R7�b9Ksq�n�\��EI��ٔ��v�]��>�bX�'~��S�,K�������Kı/����DȖ%�}�����Kı;
�&F�4�*���
�RB��������Kı/���'"X�%�|���'�,K��뽕9��L�b?/���na] 1�������o��ۉȖ%�b_=�w��Kı=��eND�,K�w��'�,K�fd�&Zm�9i�5T鹅d)!I�"g�~��O"X�%��n��9ı,O}߻x�D�,�>�~ڜ�bX�'߿[���t�.l�&乻��%�bX��w��"X�%����'�,Kľ��ڜ�bX�%���x�D7���{����r��M2�u�ۑ;���}e���M�s�����[I�e��#�_s���t����l��Kı>��?N'�,Kľ��ڜ�bX�%���x��&D�,O�w��Ȗ%�bw�~%��6���ٙ���Kı/�gv�!�	�1I�����/��<�b^����yı,O{w��Ȗ%����v�_�S
�RB�ժj�sBy��6nn��Kı/�~��O"X�%���{*r%�bX���vq<�bX�%�����Kı<���M7v̦�۷ff�Ȗ%�b{��ʜ�bX�'����O"X�%�}�;�9ı,K���<�bX�'�g{-�ni��35��*r%�bX���vq<�bX�%�����Kı/�����%�b�����aY
HRB��e�ө�Ll���Q���u���f�N��v�5�;54]������a��-��)t�o��{��,K���q9ı,K���<�bX�'�]��)<��,K��Ӊ���oq�߿����<�Og�h�|�bX�%���x�D�,K߮�T�Kı=��vq<�bX�%�����Kı>�g:]3fYp�2i���Ȗ%�b{��ʜ�bX�'����'�,p��x�i�O"_���ND�,K�߻�O"X�%��w���텻t���76T�K�ʄ������yı,K�s���Kı/�����%�`~I�>���S�,K$,�;��t�4�leS.�)!I�}�;�9ı,K���<�bX�'�]�Ȗ%�b{����yı�{���{�ݛR�v�g��x������I|���[��k<\˄1��S��k��U���ݩȖ%�b_=�w��Kı=��eND�,K�~�g��&D�,K�s���Kı=����4��2��]��7x�D�,K߮�T�Kı=�~��yı,K����Ȗ%�b_=�w��Kı>�;�l�sMݙ����*r%�bX���v�<�bX�%�����K���/�~��O"X�%��n��9ı,O>��wd��囹��e����Kı/���'"X�%�|���'�,K��뽕9İ#lO}߻x�D�,K�v��ze����T��oq����};��yı,O~��S�,K�������Kı/���'"X�%�����&��(E4E��e����ەx;:0��̒[ZD���,:��-�M�q<�bX�'�]�Ȗ%�b{�����%�bX���w�,Kľ{��Ȗ%�b}��電��fͻ�f�ʜ�bX�'��ݼO!�TF9"X���ۉȖ%�b_���x�D�,K߮�T�O���2%���~%��6�n��woȖ%�b_�n'"X�%�}���'�,2&D��J��bX�'�o�׉�Kı;'N�8Ӛm�,��B���؄%D*�w_Ȗ%�b}ۿ�ND�,K�w��O"X��2&}{�q9ı,Ol�M�*h���*��_��$)!s���9ı,O}���<�bX�%�����Kı/�����%�bX���'�L��܄�~0�]�B���\lq�{[]��n	2�16\�x���]e�ñ����g�]V��
�Ŵ��ڭ�q������tr����t]=�{V�ҥ ��ܮ�v2��&)��M��v�І�W	��$�X���:��(��눉9\cŶ�%��I��q�Ck��b�@Vѱ�lU3N���G;�q@<�GĘ�=�ux&\������=��*i�띉X`�FKa,�C�;,5��\l�'5�y�2�f�`�Mۻ33Y����,K���{�x�D�,K�~��r%�bX��{����L�bX�v��S�,K����3��sM�3s7f�soȖ%�b_o��ND�,K��{�O"X�%���{*r%�bX���v�<�bX�'~���0ܻ���K�e��ND�,K��{�O"X�%���{*r%��F"}����yı,K�����Kı=��s�]7r[�i�r���yı,O~��S�,K�������Kı/���'"X��I�3߿~�'�,K7�����jw������oq�X���v�<�bX���}{�q<�bX�%��߷��Kı=��eND��7�������߯�.��
�ۚ�j�u������6�g&=�����Ѷ�[����b��.K��v���{ı,K�����Kı/�����%�bX��w���,�&D�,O����O"X�%��O��5m9���K%�P��$)!I
~�c���Q��#"dK���*r%�bX�}��x�D�,K�~��r%�bX�wo{&��f\��mܹ���%�bX��{§"X�%���oȖ?�ș�{�q9ı,K�߿oȖ%�b}2��,�sMݷ3Y��ND�,K�w��'�,Kľ߻���bX�%���x�D�,K߯xT�Kı<�y�ܒ曖f�n͖��'�,Kľ߻���bX���}�����%�bX�v��S�,K����oȖ%�b}���&]3f��v�n����;,;/'���h箬p���sv��v�;�nق�f��v��i���'"X�%�}���'�,K����9ı,O}���<�bX�%�����Kı=��p�t��n�M�sw��Kı=���NC��+�6%������yı,K���q9ı,K���<�bX��o��sS�3h����|��{������oȖ%�b_o��ND��x+P�	�.��"X��s��<�bX�'ݿ�T�Kı<�ܽ���B�f��ݼO"X� @ȟO߼��Kı/�~��O"X�%��׼*r%�bX�����yı,N�ӥ�i�6������r%�bX��{��yı,O���S�,K����oȖ%�b{;�br%�bX�|}y��79)6��i6�$�v{\��1�p�7k�"և�v��#n;%>wy�����Ͳ.T����X�%����*r%�bX�����yı,Og��'"X�%�}���'�,K��e�fM��w-�nnʜ�bX�'��{x�B�J�D�~�S`�	>����)"{��&���!I��U�M:R�ӡ�4��|B�ı>��s�,Kľ���Ȗ%�b}��ʜ�bX�'��{x�D�,K����tܻ�sm�Iwq9ĳ���؛��oȖ%�b~�w�T�Kı=�{���%�`z�� C�r&mȖ%�by�l�It��nl��r\��yı,O���S�,K����oȖ%�b_o{���bX�%���x�D�,K������پv��a�3xP��l�����]��Ћ{<��LGn�k���3u�f�ʞD�,K�����%�bX����'"X�%�}���'�,K��뽕9ı,O;�/t�6�̓rnf]���%�bX����'"X�%�}���'�,K��뽕9ı,O}���<�bX�'I:t��6�-͹���'"X�%�}���'�,K��뽕9ı,O}���<�bX�%����Ȗ%�byݽ�n�3v�ۓ3w��Kı>��eND�,K�w��O"X�%�}���r%�`*(�]��_��$)!v�wF��-����\�S�,K����oȖ%�b_o{���bX�%���x�D�,K��T�Kı*}��ϥ�oH���A�pGc�x�)FD�� GSC��Ͱ��`�zծ��֡;=�Pz�M�x�4�S �z�����.v!6����7#�u�&?�'>m��+6:���ڵf;W;���,7n�}gm��:����k�|]k`rlT�nN�n�:��k�b��2;��'	&�g��\�u�K&yv�6{�84-�ʛh�N���K�Th�3��!��~�ܿ��]{�狟.��s��\���<��#�m��ˮۅ\�ig���wnnM��ߓ�,KĿ���yd��1��^���G(3+ޛ��~&ZnZm������`fo]X��Xٽ,�D�R�bl��NK�ׅ��Vd��IyB����v�������N8�$�ܧ)G1�+ �7��}����6q`}�JI�E!�Aě� ���`yB򄫹�>�����+��ͷ����95t[�1S٢7&�Wf�Z��\P�a�b/3K�\ǚ*��熺��6Mݠcv��m��Z� {5��k�%I��)i�`}�8�����0|��T�R"Ă��"�� �:�g���߯$�35���w�I(�;9;�Rܺs.j��MX�ݧҀ=��&ou�3]���1��"i��-�:3Nl7�]��@�~��m���(�m�7q6�r1SI�`gt�36q`f=�`gt�7C��19MG�BD�$9�i�X��9�Bmӈr�bK�܆-c�3w�w�|M���T�M�F�I���<X�yXٽ,��.ޔ�R�8�%(�`fV�@�v�=��ٶ��DL�ݯJI�E(��8���3{��>��ec��a`@� ����"!ՁF!IbP Q�Qe�W�����ZF�J�d���F��B� �J2
J��0�Jє� ���P��Y;�n@��Ć����ր}�$�C��!��&�]��e�*����h��@(E^�P�D�P0< P^���C�S��*�����@��qT�ꅑ�ྟ>��o��O>��`r4��NJ#Tۂ��Xgt�>͜X��X{�Y��`g�^�)"r%"m9,�gc�V�oK �;���U\�ޒ�JJCqG#t�&�v�;<���t��i�^k!�͹�cSF3wZ�s2��-���l���; ���Tz1����`o��΄�7JD� ���=�� �7h�j��P��&n��NF*i9,��f�,�[���7ޖw%:�*66�8�i9,?DN�\ 7i��cv�D}�菒Y���>]��R�S��p�3�6#ʻ���s�v9ׅ�fw1΄�vh��ə�W��-j�)9�7���%��ˮ���+���2�����>�� {�f��ܠ�8q5v�R���ɦ���w��(��35��3�����_�F���rNF�M�-��e7(�ݠ���5�)8���~jB��n�yXo�,3�X�8�>ލ󤜤�H�dv cv�3�f��؀���>T�5o�U��H(�_��ë�[q�Y(c+wb`9�G�ذ8��y�
�%0�+j�gL��y�8����q�4�/gA�ܺ��QN�J��6Ʈ9��h�}=\�����Ɲt�V]���0q�mn��,`�<Y4m����:��nF�t�=;[T���a����HGm��N�Lnr�:g6%θ)�7)�6$0h�A���n��s��j;o2�q���������f>}B�:��5Z�UnUt�|ɎҔxl�T�:�Ѩ����lW����o����@fm����ݠ=�K�qwCnT�ȓ����Ł�Ӌ �;��fwK��Ҝq�I��C��,Μ cv��&M��@n���ۗqUVQM��JE`gt���`fl���}���Z������6ࠜ��7h��k��O� {���S�ƆGJ5S��������션ex� �f ���4�J���Kr�dc�&f���P��@���5����͗I�����'��ݼ��H�؎��@�h[�@fm����MU)njZd�s`gq���v~(�������}�`wj�ȕ"Q��b���A��g7��]��̭r�<����N�J���R7 ����,Ǽ��ޖ�wK��*q�� �#�ۮ�ۗvo�Q�/b�\����)-�+�9+A���\�)�����:M��7_yX�v�=���G�w�z����XU�2����w�����s��������+�7�&Ɇ�M6�QUL�M7`��9μ,���!P��P�.�-�+ ��sK��p��a�ﾈ�ָ@n��@�� {���`�N�-N�,r��`z!(�wu��������jǛN��~�����>�ؒ����ӥ�՞�<ڕ��Ƨv.ԥ����n^-:�[m������wK3gc�Vv��R�t��UrX��/��~�H�����}�`gt�>�Ju
Tl�G#r	�`fm��Z��d����hK��:u*f��h�5L�ԗ�"f^�l��; ���ê�(�Q"↩%��@�fy��'����6�3%���f�P��@~�������eo+WurQ?�,n9(��� ��K�T�7Wm�#ڮP��.�+tl���_����s͆��J	ɀ������Ł����}����iwrn��9,͌@fV�@�� {��u�����KDӇT�������v~%QToK���V�Ѿt')�R7���n���@fkP�̭r�of�i�K�ꓤ橻 ����؈�Y�ߗ�w��6�w��
�
!.�BG��ߟ�'}����bkݍ1D�4<�)�a��Bs�tK*�Ӥ�TrA]��Vx�&ؗ/8�/�u�Nȧ)b��wό]K�W8�x�j"�;���X.ݵcY-=�����fN���)6}6��.k�In����ԱJn�c0ef��5��i��U�<[�G$@$�N5�X¥��b�ی��H�.�X��n�����p���I2���e����������p�)�ᴳ�Y��Tz�Ln�=�`���Q����ݖ�W)��q�I�����{+��zX��,�wJ�ĩ&MSE)�Ձ���M�(�Jd9���9���77�����Q� �'*:I�`z� {����r�q;-�rQ�6(���>��`fo]XX�������}�`o�^�' &�9.���� 22�� �7h�ݠ?>�~~|�tWgbF�h�,�I�9�9Y�sf��ۘ�;l�aM]R��h�ͮL�m�`qr��`gq���{
!}!��]X���(NSt��"���>��O��D(�䁼�@<�P���nP�%*AF�q5M7%�fwKsz��%3��ݛ ����cN����L�vQ��s~VWkvl�w�fwKoJ�ĨM' :NJ�2����n�cv��֡ ���)�{B��滊'�8�U��:�v�8\�b9-���chv^�����ϟ>.����<}�$����I%��>�$�_],��i,}��$��]�)�q��r;I$�5ݤ�cۥi$�����I%��;�~�ʹ��/x�pM�'�$�s�Ҵ�Y^���yx��b��!3.g{��m�w�}�Ick�����9�9)ZI,�{��<���w����}���<��"��&���������W�v����p��� X����_�_��3K���ZI,�����~�> Y"��Pp�ۖ����ɮ���V��c���Vݻ\�)v���Ʀa%4���I,����%���ZI,����Ic��I}ܕ�)RBT�8�I���%���_����Kkg���$��z;I$�;��U~�m�~�ʑĨM' :NJV�Kkg���$�>��$���|�[��� �����(�<������?��EW^뫙���w_�L������d���Cb��GT�S�~�ym��d��.k��(���I%��>�$�_]+I%���}�I,}��I/����I��H)L��k�);y���Q���nK3HFΌ�[>z�Æ�����4��������򳯏�I%��?��U��m$�}���%��x����'?'%+I%��|}�I,}��I%��>�$�_]+I%��o�$�'I��M�}�I,}��I%��>�z�W����~�V�Kk}~>�$��]�J�R$�%)��v�IfwO�I-��J�Ieg_|�Ktv�K�䮺���J�r�����}t�$�VN���$��Gi$�gw|��~>8H;B
 �D��������,[�=p�$k	��;}�qT��L4�B>s�
�ď�eh���B/St�Pbj�@"<�U"� 0�a���3�P�� ��`Ɉy'��M��`����,L:����rv�p�X��]��V�ʖq4Wl@؅5;�9��J䀁�U�u[c']E���(�n�:DםC��h�&vvj����ѽ�q�Z��X�&�7l�sE+��q]:�x�s�x�TN�
gm��|u��v�;[�09�VآYk��<u�^t��!v�`���:�cY�3�gY^�>β5ǂY�8-̄�/�0��`�f.��8A�n'n�E��$A�z7<�t1Fw8'<.�K.t� ��4uq��GZ�m�A�s��3A���"mκcb��ƣ��UBCB2-r5Z��"�7*�ꃈkv�B%��5ps�Y�]��@�m�I3��Ÿх�Wcm��k>���ҷi�-\�;>��5�W&f�Ru�=*ʵ]�nv�t�����R"����<1�lGv��qU�s�D5,�����Y^�������A���kMv�<�r�����ձk�ll�k��5�1Ѳ���n�;U������]�V�G�
�3����= ��a��ӻp�G�C�q��=D�.6�\�on���c��dŻt��1�h�;H<�!$���6�+���s���Ѿ"��������cs:by[����4�2����Ο@TS��g8 �.z @��ـs�ݘ+F�����Z���� ���,v�ꪬsV�m�m��m@uQ`
ݧ�#HsR�I�l']8�֔4\��Rl� L��g`��)VE�p�R�r��s`��R�7m&Y�i0σ&ɟ$ �����gs7s�&%�-uun��܅ ��WgmH�*��Rd˃�L�Lϋ���u�6�FO��&��0跀��n�-�b�ꫪ�x�+g�m�q��]dVRʯχ���~: m�+��T�!�ki�/��Ā����P696z���l�Ofq��'H:��>|�;���v��Ρt]0tb�ݵy�O*��t�u��RJ�g���r4<�Yo����K�?`���T: z�ϝ�C�7��U����ze�\�3�9f��se��[v�n���;]�g*bӝŦ��B]cGa.1r�Z��2�fCm-�ʻ� W�F���I�����(.��姗�K#>�6G�mV8��n~l�E&����[^"^˷m��)O��;>ݱ��B|A�1\�I;(�cdZyI��K��Hݷ,��(����l�L����d6p��Mf�;�[�6����0���~����W����4�I-6����Z@;5�Cgk�')Ѭ*�ۢp� �{���/�����B�<5�� ��������	,}��I%��>�$�_]+I%��])*3�"������~O����r�}��g1��s33�Ǚ?}�	%
��T��9(��J%▒In���7_r����R[Z��`f�yX�.�N@I���4�3�2��+�}����Wꨅ3���S�5-˥N��p鹰8������ n�Z2��Χe��j�TZ^�s׵nyz+�y���9፸�G��c��c����p�Vw#6��nPcv�̭r���nP�h�i���i��f��9��#TB�ĥ(���iB�BI(K�5׾�V�zl�]ɿ(�9�2֩i�M4鲪f��9�͔FSr��V�@��j��f	U-ԍM76JP����ٰ9�͛ ��������])))4�QD�W(ek������(dSr������X76X-����]�=k��LX9x5�:�As�[=s��K<�l5�Ą���9��>�w&����'R��J>��}�`o4��N@R��4�>ǮW菦L����O� fk�:��&[��6��æ����ܮ��ԢUA���"P�� ����t�3�>���Br��8H7*���P�����37����ܛ+:q`wr�J��
��P���3�ﾍ�K}>cz�@{+\�7����6��!u��e&I��Yֳք%;b��<�e�P�K����{��]V�TNSI9>5�����8�>Ǽ�3�Xwt�#�&:�R�9���8_���&L�}(w����(ml��RRi��T����=�`�������W�_yX[����X��I(�I���z"&{��`s��61�aiD��p�� ~|U��~��ϲ�ߤ��*hiӧSM�r��`yD(]]{�����3�Xv�#P�n(�Fք׎��g��o8��x�[Ӛ�וӶ᥇uQB��D�����XX����=�`�����>����9M��G)Ӓ��V�_������@f��@de7+�$�d���&Zl�Щ4�2��{����(��G�L�mwJ6�J���8R���Iʉ'%��=�`ec�V����fwK �q$�*Jr�"�22���>�ͷ����@{+\��������$'�6�ۙs	�3���f�g�q���Qj�X�p���m�����1��=X��wk�k�4�^2��X��x:hs9��8٪z�5��ݲ\X���WFA�m���:8��{vn�7�l:
�"r���q���������n];e�7��fb�l:�<s�ٸM� 2�5t�u��^��L�����r�n�+qӖ7N#���ϴ~�{�����}w�������	V�K�����/%G�4)R_���.!W��^�a�P	\I��QRN/�3����3�Xc�VV>�`uc]���~��%"���1��}2f��@lmwJ�Z�1(�4��NJ)�*8�NK5������Xc�V��,滥
F��S�Ḿ��̛�Wrl��v������=���J��j')�ӊ���@���Z���ܠ)�.�]բF�W  =c6#��9�JJ[��,�ck�F��oP�.�u㮻6�����Z���ܠ=��Pnf���m����L�7`}��Mߔ%D$�G�B�rb�����Vzl��v��m7Q$�)�����Ǽ���+?�#7ޖk�+�z�RRRi�)T����}D���@�ր�V�@dek�V5�	�G�آPR+ �;����;��6�����o]X��t�	5!R��DC�9r5lh�<�[ãU�z�
�qg)D�rQP�!i�`}�yXY]ɰ>�r֯D(\�;��L��y���)Bs�r+k_yXf�Հ}�����;:6�P�m��e5"�>����y�{�����E@!R$d EN��j�U<�������Vw.�)RI �&�%��<�D�;��v�f���w&��7���JWR�$�")�rXc�(��r��kP�=��]71TM�Ц�m��e�/e�kz�a�r�B�,Җ�9҆�b�o�<�o}��-����1~�66�J٭B �7hek���]�RRi���*I�`}��V�wK�{���Ǽ��k���ѱD�$��k����;�g�i��3_(@y��a3M�7#c��:��μٰ5}��y$�߻Òt� s�+/�!��W����>ֽ҅#n
P�*9��+\�=�� �@{+\�;��x���͢]ф,��b,���F.2��uu�1ۀŷf��b�Nc_�����vL��B��`����9f�>Ǽ��{�����%*G$)R�$�`r��`}�yXX����o]Xܔ��*IQ'*6�v����ՏyYꤳ{�V����gwIR8���9D�XYZ��֡ �5��Z��.�f�!��GM8��z���������]ɰ1^B�BUu=�(%���+�����kt�7�6a��3ds6�=����lK[t��UlVr1��\ɣp��U�:8ڣ+�����v����6����sجm����m�%�%�鈂u��������7'I�{-�씒�lg��84��ݹۆ�/��.�6��K�)�7�^�����\��Woh�5c	)����(�L���Aظv���r�ܳ��+e�Tz����{�yn��/79�n��{Z^[���Ժ��G�N#�(6��qnQri�NJ?F�������v����ՏyXf�Ձ�4����T����WHek��}�D�Ѵ�P�� 溿ș;�;H��9h��鹰5v�f��7��[����+q�k�
F��NT)�����.�;�{���Wv��7vvɖ�m������VOu��f�����٭BccF��[�$s'E3�I��Tz͙�Gk���7�Vi�Ћw0V��D@�*����m}�u`}�*�3]�}��T�m��w.i7v�I����=(0I�(R�q$��Y�s-X�w*���ܛ؊H�~^�����I�)%X��������6� �*[	��>��D�$���;�{���Ǽ��z����]�NJ*JR����+����3_(@9�t�܂��]�m�6`�!I�kg�u]s��c�7jܦ�T�&�n;+�u�ەړ��$���(f�9����(�کw��iʅ4�>���o;�{�`b�w&�DDɻ��L��m����Fڰ6{�Vܮ���V����!Z��e$D�z�,�9��hDJ>��'�Y�bl�"}��Grq�=�D�ٚ:��1HS�BE-#
�A����E�!**'� )"�ǜ ���Ł*���7��X! �!�X	�őBH1�	�A`Ȓ�Y,a �U �H|j'PS��%L=T1� ����P�U�z �Qk�D>Q�'���*�va`}��Vq�p'RH�"r�m�a�>�#�ͷҀ����js] ��*GT�Q�(�+�6q`W�������{����7�E�j�iN(V���qD�e�sθݳ��L������<-D�m�)G(q'$T��`}��V��Hek��}��|�ѵ=�5w���$�`gt�>Ǽ��޺�>�r��P�	U�L���6�܍��M]�5�~�FkP��kP�=��.�IH�$�*B��XY�u`}��W$�{��$��?�h���HF��R
���:>�����O}�ٗ��i���M4�Tڰ>�rՁ�Q<�����VVo]X�y5'*2�r�9w7��b��̇[��6FMǵ�엮��p��0��$��%$I*�>��`}�yXX����o]X�)]IԒA�ܧ3-��WroaD%2qw^�;�j�9�����$�zJ�ĕ9I�$���޾�jf�@{+\�7ki�]U�'d�Rnٽu`������	yD(����,,���i�&R���� fk����ѕ�P�j&7߿S)���M��$ݶ� ls�G{Ma;Gc� r��z�k7V^����U��+�U\.��m=&Sd֫ifnz���\v��1����ct���T�[����.*:b��Su��6<Z ���on8���ӭ]����t��uEr�p�r�g������N�H�6�C�tٳ��N��,��2J�/n��%�@��V�=r3�
I�8=��{������������_ma�eۋI���&�ڠ�:�\�amt��h�M�r�xqV��5ۤ�!$jI����VՏyXf�Հ}����k�����Sr��$VՏ\���"d�|� f������:�u)9iʅ4�>�� �;���~�T�k�+k_yXܺĥH���	%Ո�ݠ=��PZ�ﾈ����`o�)^��H�5��NK�{Ҁ���(f���@������JIi�=u0VԀvkp�����y����8]k-�I�Uj�`9�������\�=�l@���r�ܭ�quW\ͷ7v���I<���稊y>�uV�U���{�y����}����V=�`uc]���T9�`cv��V�@dek��m�K��f��DF��������yX��V�wK�kx����$�ENH���r�菻_z<��h��P�������O��N2���;����^���zq����;S�m�	C�Ս¦n�����3#u���|k��ݠV�@dek�w.�)R*NT��RU�}����{�`qr��`g;���2wM��M&�5Rꚩ����f́���M�(�MB��E(�	DTM�o-X3q���m6�I�JJ$���Ǽ��g�wK�{���z�Tn '�5IH�f���7��m>�FV�@d�~~R���t���T�獙�&�s�����7[!,:-�<No�i�����[�i����n���(��r��m���wrP�		#NK�{���Ǽ��g�wK�RF��x�����YUwr���}(f���@{+Z�;���)#C�9P��Vٳ�$�{��$�{�v�N�4P�����舎j��M��2vɖ�%4�uJht� �7h��D~ֻ��w�@<֡����?>}*XI\͂\�����jk=hqƽt\��N�Ռ%;l���uM�-35w�;i��22���jcv�>��*7L�Ĝ�H��}���޺���`v=�`j�|�7 8Hڤ�Vf�ՀfwK��++r�;M��	�D)ӑ�� ����(���}�DOk�Bg��	��B%!$i�`v=�`V��y|��j�9��`r&"%��Y�4�UMJ�wigk��\�ԪLl�G*�٧l�U��j	O-�BR칕���f�'�jt�v���:�2q�댹��[Yݰ��x����;�:�͎�q�v#V�9�w��]v�ٮ%�s�v�a�a��|���
�ݭ�x��c%�����̅��a�Ĭz��K<B�#�+�}�6u��:6�����ж�-���i�sk���]n�"?�N'���yMݘN��H��/N�O���t����R�����n^�:���qP����ͷ�+zP5�@���}zC��J����JRF�!
�E`}�8���`}�8�2��+��X��#"��N[V�f;9ׅ�	BQ
g���6�z����R��$N�jII��;6p���nP5�@�� ��wUs)�JJ�����X�{{�W���`vl����e����QH��H�F'y*=i�H�c��壋cV_$�e�V�� �rEIH��޺���`vl��B�C���6�u�i�AMԺmrI=���r�� EJ��+�8��Ev"!K�p���`j�ݛ9ܵ`ry�'�HIrX�8�2��+<���u`���>ַ�JH�n��qUv 22���jcv�y��c9�QH�!
�E`vo]Xgt�;6q`ec�Vp����G��\ ���dq�T�ϙ ��[X�:q��V)��"�*A2@�RMIV��,͜XX���ٽu`}�)���M�Q�M$�;6q`ec�Vf�ՀfwK �{���I9�IC��2��+$�w�&	�G�u��}Q	D������~,�X��r�6�ʙ�6s�j�9��`g:��DU-���=�E�Bq�
t�j9*�3�Ͷ 22���j}����	�	UUH�i�u\�F�2g��fB�;o.���T��y�=Y�.n��H4�����M��1�@{�=��m�T�T�J�����fM�(���2osmX{���^r�gTD�!Ԓ&TR+�z��3;��
!)��=,�����8�F�&���S5-���
�3�v�_������� E_���E_�_�b}��������t�r$�rX�8@de7(�� ���Z�*���ʅmæ�������T��*��c��F1T�ua͖�l���������� �3�B�^���k�`nW���D	DIT����޺���`g:�8�Y�~��2n�Z&�!����������6؀�e7(��X��1N��r�M��v��S������(�� �;�ր�R����55J���Se���̛v"#{���'߿f�>���rI�QQ_�QQ_��EE9A��TTWQQ_�UEE�U��U��QO��AX
E `�E b ��,Q@��E `�P(��1E `0E `D���UEE��ª*+�U������*+�ꨨ��������ª*+�*����UEE}UEE�b��L���g"�� � ���fO� �ξ =           �   :4      �B�@(T"TH!T�� �T   ��J�($ H@ $   (  *T !TIU   ԁ@
(�@� @4��/����]��-{��k��i]�}��}����ד^�=�w��>N�m� 4��Js��z��o ��AL{ʹ�>��'����˻x��ܮ��+� ˗{ڗ�ONN���ˀ�  �
	�R��@(� ����׷����Һ���o^� t��w��朚�\ڜ�\�[�ӝ=ngJ��v����\�^x }>�K;w�/qg�L��M� .�M<�N�m=[�o+�w��l�� �@P ��( b� w�����\ZqçqwMn N��st�qwzN8 �  �   �/}v��< Z��N�x�K�� �>��6���n�f��p�{�6�ιn,���S&����Q@� P ,m 4�}R�޷��=�o]�˺�ŕv���y��W���շ;uMź_m�z�� ==�h" z>� 
1 7X ��
z@� z�� � �)�@4`� �vt  p�  P�(
 6 @��ѠD�P"�`:  � � 	 :@6�� �<����\�� �y�{{�s$��P�|S��=<�鸲��w*��@>{圻�z�N�����v�:����*{�P  "������*Pd ѡ��=U*D���CL#��R��UC#�������R� 0��$ �S�N��O��?�������S���G����d���D?���**+� ���AQQ_����'��g�B��		%�iō1eȰ�p������"el$��i��$\v��=j��� �#y����>D��ɜ�{h���$7��a���88n��2�c9&y'�1%�̗$�̦P��f6VH��$���#�3YLMg��Yr�tԄ�L�@���ݫխ�ȝ�A�8�����B�<�<
f�L1i�S	Np�	�n�@�9�Js	I�
��>��<l�d82���M����J�>�������>�� !�MOGjƉ\4��e�8x�4Z�s�nn\�g?��S]=<� ?y���#2�ja�	�
.dfۿq�y�ϐ:y�����b`V�������Jrky zDؖ`nȴ2i��y�<�<`��� �]c���	CM$�ς��u��=nM��b[��咐���X��+�F��X�#�X�!��l��H��e�-2�X�KI��C$��>�	c��4)
Hf�M��M7�jy�GI�%0כ'!rں�%����L������L�W�����(@a�!\F��Dp�B�1�4�Hؤ�=����<3-�r%`�+_�� @��%3J� �h�l M�XP��1X��!T� Wь	�=)�B��bq�ߊȞ�W��	�4!L�ZHz{���
a�@�XC5���p��B}|x�>5>��$�R&�O>�dH�o����4c F��b�X@ �4$��D���\�Y����x�xR���R�A���\�R8�� ��hĊE�!�c*��b@�E,��N]�O<���B�����)⑩��a���H)
b�	�	 j$@�!���
�!�$@��
@�E�8	�D� �P��ꑤV+��h��P���hJF��(��@(�	��+�b�"�qcL4����qВ2���Q�Mx�''!�.�Yt"�]afi d�4er4&-��HY�!���,�F��.l
���8p�����Y�	�
e|�9�0�4a3j6L���762\�5148�:zB���H;�H�SN@����,<`A�Ƹ�MR BQ��@�C  S)@`� �'���!�|Al����C��fo<��!���ܱ�=��Ӓﮇ `X�������B�B	)��z�h,D�� " �Z0b!���"�0��sė4r%��#BR%͐���E*�/	�L�WQ�Ir�\�F4#R53C��H���BR#n����brB<��̭3x��e0p��fj�k90	Y��¤����8HC��'��7����`F1%kX`E�8q�	sxU����t�)Ni�4�a���
�~�-��)(���� ]s25	o�f�ai��5����k�����/�)�>s�1����w���%�*F��c����4��㻖�^g�#HH�
�rF5#4�4liB�!�i�I�-����$�HS\+ ������E�z�<H�˃��N<#���� sÂp�3y�0�!V�s�%<��%� I �!VT2s�B���,݆�4h�!�
��Q�_����,�^B���"}Iw��M5xH�. I9a�X�]�\w|6���5�)	 u�V �=�	߈q��	��>y�ᵟe��F�!�,i
���.jK'�i�9MS:0�dBG��yBI@	7�
>D��LMR�!��$$'23b�) HBHXT �!���U�$�"�&<�j��߯�L<`p'ޘp�́��/���Mk!��7���Ik���rrb5�,��ؒ@�YVRA�׀K#
��M�$4�d���zy��F�J����v@��d����9�K�fI��R*�5��FSB!V(E��~��!LB,�XX+�P��Tr��6GB��CU< Pqux���(�K�U���&bq��	��2\�0		�<(a�$���$�`T���᮹H�c^>BB��'���}7�L\�_Fs5��@�i��[!�g���17���Ĺ	�=���47y�a}���F�������m�li����%%���_c���f!��##&����H�-5�U�1�dB1#I b�`Yn�E���
�K�Yi�F;�2(0��0qYr�$�.��B�
�<cL	X�H����e��k
0*��$�ĀCc3�X�]�$������:�)��|�d˺�����x,.O�0э1�F�ap%�$�L065\XcC	P�HԃD�u�0�ub}HJl5�ݢkN�BO)��+r½up��)�m�p�4!L|�{�L-�>l��]ü��l�=Q�wy��8xw�g�	FF �"f\!����"�6		Y $_��&�Pq*��BWd���y0�C�$������)��I-��CTa\+K#�%�֯�%! ���}�4��˚y�9#�ql$� RE"11W�}H���,!)`L$���F�r&�s�2!D�_<o#	L49�
4�D���z���|w�I �
a�y��'�~�<���뇼>X\��f���s�'/c�!�|��Ξs�0M=_CX%H�F5�I%L��rIqі�d�̙mb�����o���y�V<�c����3x�a�S2FB�XG��d>g7��O0�WС�B_n���
����*p ���ȑyJ�ř�Ǹ����c� �	����Vv�<%���̌�̻J�CK
�$������T�x�/9	��8���c�D���C�ӂE�;�"B�K���|З�IsY�����S2��M2\��I�#s\BR[���5�S����p�)fe�i.0���C.e���,	��RE%�4�2�.�Sq��	���(ĉT*�$(aM�5k�>�HS��Osb�Ip�B\�*�
�zR���,��!BR2�K0B0h�)fB��X�Q�c,0�� �B��hB$�����\�$�&dId`%�4���� ��"�d#P�H�#F$ ���	��c0�`����}Y���%0��Ra�
0i T��
������$ew�� Hfp�� B0�p��.�� G���y$����"�`F�WZ�E�,3H�$��2�!(Kq�>8|HF�Y�� "S|�)�{�@Z0R$v�Wt� `����
�c�$��n��r)$��!P������5	�y�S�xb@�x.`��r�J�8����BY*�0����2`F��ǿ)�D�� ($�'�f�+���X�q�!ώ���
B$�HKRL�`@(J���$Ri�[<!"F���)�*Aׄ�
� z�$J$�SA�t���S-�h0$�g��L����$$hƇ���Gw�dT��D�x;}fDvH�)'~�� H         �*��vA�7;����UK�1U#*�kXW�4��   )��ɟ��?++UUl���1��GU�u�]���� :v��X��F�9��̽@@�2ÚU��ۭ��V�-��$CAJ2�a@eF�d�8���U7Rh���m�#� m�\���8yyP	�Ԃ�U|���jT����[P��+UXpܫ�ZVSynR�4@�ݮ72����kd�em�6����c�����k&�W��m�m -�� m[n�m�f�	6ۀ���V�H�` :�a�"�m���im��%��� ��5�  I Im6ؐ� ��l,�V�"ջ��۶���/.  �� �-��nٶͲ�� ��1�jɕ����  [I�$��L�	M�p H��$�6ٶϯ�}��` H@6�m� � ѵlA����M�m:`��4i�:��  hm�  G�$$8&٭�;U[Ru���E�p�;URq�j�髭��W�(�m��m:��Kh $m�kv����&5�I�fV3�m��$    m$�  � �   ��  $-���u� � mٴ��@p��˦��(�  6�Gb5X��*ա-��>�` $��@6ۧ]���X�j�^ͨ'ɱ�j���Z�Ny�;��T��K9v��櫩V���� ����m�  րڰ��85���%Z��+�6ثj��T�v�e����S�s���m���5���`�ԁ<�e���ιn�� ���/ZL� ��H�:���z�fݺ���;9z������^��W�F늪��ЭmUW�K��U�v 
�m���69m ��m�g:�ܼ�\�  IJ"Zַ����o\pH@8I�^��ݦ�yn��gix�n�[֨�p���wb�]R�Ul����b��p%��'!u1�Im��]�aU��pЙ���֨�:ɳA�,m� v����K��M85UA�ջ<���l	�a m�6�H���n35*�-�� J��nV���{h&U��;J��- ݦ�eč�r���ꪪ� �cSAm�8�/JM�e�%p2H�IĀF��9��&�+z3K���5Um��UWg���#<��U+�O*�⑷i��8d��A�<@�����̼��UP�ʬ��m������P����Ii]��6����2xl�NuAʾ�R����$�v]oT���4T��s"��`�n��v�LH$�� ���6�kҎ�J	 m��V�km���`'��դj�
����_^���d[\�$9�mm������]�-���Tv�¸؛�� ���$�� �I�m�ٷLҮ�y��� B��U� H�k٭�[��)RV�1my^z� G:������`��٤'��<�N̺Ĝ�ȃq�k�L���[���ڧ�U�J'K�f�  � � ���U�l���8 m��;m����� �i9���t$���� ��X��  m�����-��` �i?u�}�m��� ��` ֊����t;]�  	mm"@  �6Ͷ l���/�/[��mH�@�pޠ��׭A�*�u��s� 'N6V��mt������ ��-�m�HIgl����[@H���i/MTM�� ��   M�o`	j�RK֕�(�צ��ht���f�t�Am�@   m� 	�� #�ض���;Ͷ$���p۶5ʣ����kh Hp    K)�:v�,�8m�HI$��Ͷ6�m� -;r��UV�(��T�� p6���� *�V����ܪ���iWE�һH  �m�`H6ؑ $�� m�$�kn�	$ m��Iz����UPqQ�R�,r�lm�m�i6*v�p	$2 ���,0m��V��:�Kgi2WJ��ʷj��p�M��52�970��m-�  ݓ3R��m&ƶ� ��*��$zS�k��!2�5UUH  �m�ڪl�@P@�
�P��.��)kڪ��-� ��:�6�a6�ur��6�$��ٶm��IoY�<$�9p ~�[@ڐf�cEkom�  	��   �ޠ $M��l�\=���v���퐃�:��ݶ  d$t���ƶt��ikh�0�a H���c�[�R� �m� �R�m��� 	6i� o,��vl���%�)h
�n��T�ҠA+@Tpb��RWE��O��$m��-� �ݱn���@@[@ �	m��[@  �v4^$ �  	��4U� �I���$�   >�m    m�l 	-�m� � �$�Ұ  $4Ps��+�(Z�t�^UUi2J��/-+/62lO����V���  6ݶ�     �h [�C�5���E� �6� L�-�nڷ`@/[���Q�[+m�[An� d���m��'m;]��m�  -�h�� !� �m�  H	U6��L�R���C���݀ ����]��ѻ  p��3m�m�m��]x�I�6�lNk��mհ�`���@ [�H  �	m [@  ݶ�@$ H�`ְ     l�am  $ r��[8    �   �  �H6�$ �      ��� 	����N  6�H�޶rmm�yY	I���� ��b��UnճU*�  �   � [@ ��ĀA�6�&�FGY�,�v�� k�e� [K�����>m�V�\�6� M�,�0�H 6�H��tl eS�[� � �` � ��m�  m��I�T!s�l6�@�m�l l���8�-�m6�	�	-F� Ie���m׫ m���s�-�m�ٶH �` mfb��V(��h��R�jIW�}���j� A�m��� ��N��KL�  ж�  �� l � �l   8� F�۶ض� Ѷ� m�۴�h�����p�-�6�v�� �v��m ����  �6�� � ��
��T��lS�A+`         ��6�IU�m�� l��m[`�J��$6�t $� ��damH�n����`�m� kY [F�"0:������h��Q!m 	Y@F�7E�埔���i���f2@� nٶ �%�fu�  �M�   �  �� �	 �mͪ�ke�p ��f�m�l � � H�[dӲF�l �J^,6ڦ��H�    m�!# m��δK(�m�2�&�����:@�@Z`FG.���iT�olm�,&ԤրU��!:-*��b8wf\a�f����-�d�Hf�\��`��IU26݊���;�i0   �k]�[Ĝ޵�dHܽi Hi5nĂIv׷l���n�5rmt��7l[Z�&�d�M�h�-��ڰS[U@Tٳ�@毃m���kj�$w�����^@|s����9�Kչ�RZ�[[��Poc2��x᪜�������l�K�M�ʥmtU*�W����_���mB���+,MR��T����8�9��u���UUe�cd@��pd}'�ָt�hZ,. �a������.z���mF�d��Q��[ebM*D��$�j����Ѫ�>7m�lI ��ẫ���-�F���H�]����F�m��i�۷_6Ijf����	�m�� *����FJ��gf+g s["γ	�$;m��ڕ��$
�
 -�j�[�[Ci�� HIl��n�[d�"�m&-�j�6� ����' Tݤ�d  �6�� �kjUU�]�[aUk�A�TZ����C�bZ����R(*� �@   �Nsk3X���u�Hn@��6�k'�l�o��}��u��nV�vee�= �X�ȵUW�n�� 0ʲt��VүK�=��ZBI��%���m�R��Rdvˆj����gkn;h��@�UU2�L�f�I"�kl�`Hm�\�NHmu��fZ����@ ʶ��ٶ���)Yg�� 
IE� 	.�dҭV�O+�WV(���kB鵭	a����n��஦��W���	�;u J� �:F���Xs2���,�;K��WUS]s�ځ����L�n������s?�DAAR('�X�0F!BE���A��A8��U*�`��"0Q�e� �?�OA=4j'����JQ ���9P���(x��xA��oȠ�M<�U<�O@C�T�����p �#��PO�Tf#�A�@|S���'� �	!$�"$�B"�!"F@�"b� �R&*�4z��~��^�\T����*q }P>~�ڢ ����Tb�A|��T47�,b� H2$FX#�H��ĉ �S����Q�B �tO@�@D���< �EP�� �||�T�B���@O"�|�X�O��`(�E�קy⊧��/\T��ê�R!$SǠ�PN�T���|P~AP>N"�� N �u|^T��?�#���1P�W���-ATz)�z ������_�@���B��+ ��7wwwwv���9ed��O>,v�ryӲ��r��m��ȱ�[�cܯ�XH����5��xe�5���N]���u�MĚͷN����Ok��7&m��֠ssm[hH�e��[�SJYFӷI�Zu�4u�lkm���Br����F�V����vh&���X�k�e��0̽�ӭ���gz-HR�X_HN֩��M�7]�aN�v§ s��&��bH�@3�ڹ�[��Dt��'I�-5�N���#��I'V >U�1�ce1̭�k�)�z������X��:���zӨ9��s:�y�;��Ƕ�B�S-�]Gn��b\�n����u#^�;Yֺ��{YklV0�A�؉�����ۏl���j�����rN�$��s���q�JZ�l���Tm=t�{W`�5lٵ+�+nC�a�m��U�a��M]1�Ї�ތ�HY	p���W��1��{��2sx�cT�7Z�H���n.Vü[�������n�pٵ <;�{�{]����n�d3"��Ӽ��T������V�)� P�4�ݰ-�:4��pY�Ń�Uv���l���0T���؄��k[6��@�W��u�òf�H�,���D����Q'$��Y$7[!����u�%Sa^��:�8�RZ����`��R��a��ԙ6Uݓ�BĎu/h88e�k�q]!u�4���VIvq��[\��tW:إ�ۨşe�欷�m����$�	  bҝ����k����ә��%Xd�}#���emmHp�E܋*5�˘���(��m
��;mp�U�7 !'�r��w	Ն�+�ӝ[�E�r��l�l�n���<�������f�=�����Z�������i9#vF�Z§V�^��6�g��%J�V��4\҇{iM��X�5&6�*��Z���Y�9����"���ڰs8#�7Y�:���]J�S�eTqf���k�3�zv��i�$�Ywv�]�)����1A��BB$�`Y�  �@��qA�,� ��䙆}2c��/F��g<���'��v똖pV�+%��l�����)��� &��)�:���/l-��v0��	�N&OF�a1�<t^��e�����/��l�KLkm�4�μ[mrKO<�p�Ur��Լ��v��+��٥�-B6,r	�.ܻ �v¥�����8��ݺ��'X�m�5n�0�M�d������t��E
pG9���˓-��ɐəd����=�q�P9�)�۷)	�4<HM	��I�!��@�ܨ~̟��J?0ݝ�`f�LgS�M5R������B�a(�1�t�]�h]��㋋`�D���,�C@��1 ��� =&� ܹW��2$��G�r�@��@�l��fb�v����22G��K6�m�@zM��$�x�>�ߛ=��ݪ�ћj��fE�
��:ry
z��H�Vy<����+g88�Xs���w<}�� =rL@6�m�@K3S��UP�JN�iX����BQ)=@�<_��Q����~��v���$�[)�_0�X�LS���#�@��Kf͜�M����<��l��R{.iT�M:�*h�1�l�6{���<��zwJhňE�J,���R=�l��WdɈ�� �t���z��5�-��U:�\nP���p���h]��lSq�76��:��x����tP���1 �� �1�"�d.-����G��Қ.������y�����ByfF�M�v��I>�������98��**�)@�  ���&��EO++�/��@��%���I��'�7w�*@z䘀o��� %��QC�y1��h����)`c�ٰ?nm�����3e9���K�"K�uכm��I:[�+U�7^�~ǻ,v�	4�R�܅&����T�j|oWŀ�G =rL@w;6�e����9aUE��3f�l�oZ�<��lΔ�;��ۋFH�����$�g��v����@>*֏$O�@�F�h����)�r�d��"�U�p��5@���B�B��w�`~ÍN��U�S���o`�v������& >�U����������۵QD�;��d�J.�3��rGv�����.9�9���s��=����}n�)on�_���۹�~V��g�����+�,H� OI��ک�b��@;nbXu����� �LQ9��mzwJf�˺���s@�aزȅ0N,q���UW�}�] ��qR�$�s�b����M����uz�ٙ����}�6fV���PA!�*�0h؀J�X����8�����s=�s�YӺ��<��t��]�z͖Bb����p=WP��s�>�1r�[l;�ǫ�mݢl]�Lq��Y�jv�gr�mz��γ�w�©�h�s�nfְv���`�tXą�β^�v��gL�Y��P�����9�v�*[f-�����q.G[h�tu�{s=�v���4oF����"\��^Ɩ��VKW.=���k�ws7����d�pr�'=h��'v�9�WV��s$��a��pے�˽��dH�l��0�������{�ՠr��_�(Q����́�0���(�1Iӭ��@wd��v��@u�����R��ű9!Ljȴ^��@�^�����;�ՠ~����	DԑʙsMX{�6�͵`g�u�8�	>��@/�X�(�(��$���m�ޝ�`g�5��۳`}	�c��]�3hHJ�tNx���(��Y�ʳv�p�{]L�/�Ծ6�q�f��lKw�l�}��c�H���*@N�uu�4�-ͷaswo$�_~��(x	-�S��>=���y��w�����j����H��D�[rq�m8���b����%�d�H��"��D��=z�h�h�k��ֽ��\OXB?�aD�X���(Q0�Kk{�x~��������$�d8�o���ڑ���y�ۂ[�{�րU���M��Z�θ���"AI�˪����^��e4yڴ
�̰�4� ������I6gOs�<��lͥ��~�m<ʰQD$�H�Wj�?+k����Ǥ
��<8��tV�-���@���T��Y��PN�E�z䘀rmA �2K@N�ut�17#f8�z[2�.���ՠ~Vנ{/CIe�FG1�y4V�%��m*�mZWU�v�#ɠ�&�ݲo�����cɋ[s&6�H6'��/uz��h����e4��!ԉ& L����L���& �P@;nb�&�[���R��I�USN����;��h���=]�@�)qnF܍�ܪ�����	B�U	$����Ł����'����Hl�~'�·o��3�y���Pppx�y�uz��h����e4�$����8㈛/�j�\����uGm�����qn}]q���(%�dX(��<D�=�ڴ����2�.��
���1I��u5E����ܨP��3ii`c�l��S@�aة#��#q��dۘ��"��I�p�j�fmD9���.��[w4yڴQ
f������3i�J�E)T��lS{���$�k���b�~ b�~�WU�S�NK'����t���U��BN��Z�id�\,�Ж]J���L���]s�\E�C�K�%�8z��q����Nɑ�7��n��E��d|�%F��d����nȭ�x�[J61g`E�c-.�97J�'����@d�۱&��Lq�#��Z��������2R`L8|��9o%���6����AwB����KS��p���볺z��O��k�ۤ�-�n�7w,�4����5[���������`���@���8N���\M)UL���uE��=�36����z���;�\[�4�S��Zsj��&�ݒZ�ߪ��ʹ�w1(8౨���z���=�j�;�)��,�U�b������I�@wd��o!_I�
���29��(�4yڴ]U4/Z�[)�_3;D�9,����MvQ�結wf�ܼ.ܧSb�[9��p
=�+��t�PҺ�%��I����@u����6�r����̼�ܹ�Ks.d��'���9<�8*L�E ;��@>�P@>e�y2��@�����G ;��FWꪻs��z�����������}m ��R��b� !*�m��QMҚnf�����X(�NwO�3��X���I>�M���C��*������іB!��s�(�^7]�r���,mrl�9��Ǒ�cnO��yw�=����9����fmŀo�k$֊��nPn���EH�r�ͨ =}& 
r;+J
0��lNf��>�@����`Ō�RH�JIa$	IB�B¤���
����R�I�3�9	*�|04��lHFQф"��~�e ��!��0�|��y�c	��
@�U�D�`FT��I"���#(Ddj�x[��<:�HB*81"�<8�Jp�d�d�I���|}C���H�1B0�X1�H�
������� �Oʠ���t�@=A��!��?� �P(?�����s�,�������쓩�U-ҪSJ�SN��(�{�k��;��P�0��g���I
'v�5R}.iU9�MMrP���?��}	Bli,�����P�̝�`fw\t$�~f��������f�nM�Rxj���j�==��96zT�O/j�mw�#p���]�z&���J6fwZ�?D(K2���3:�]Z��~��9'�}���s��1������;��BQ��\+?D%ߞwM���k�$���JUQ<||��sSTP�M7UN��
��~��Q
2s���jΈI&�'������5!SC\�!]]�~wM�fgu��P�}��_$�
TX���o�~��M����O�*GC�ʩ��?%���~RY��(��3z����t���g�?ͻ-Wc�)�z;]��E�ݕ4�5�1��=�2Lpcu�o�Ѿ7�X�����ͯ �}��;�_���� ?V��INd��#�@������zנ~��������i�rHM�������1�"�v9h��{��ׄ2aD��=�w4y�h�����s�W���l��W�M+ޜ�`{ٷ�/�<�l?(�O���X(�P�G�H�8O�ӥ$���ǩ�q��g�������p^��3Qt=5�3|�������v��0R��E�ȽTA��w
���k��vǍ���X�V�[�I��������5�m��g]��Q!����52���݁z㝰��K�Y�m�Tx���ΗlS�:GD{]�{N��N �1qkD>8��s��c�k���2;���A����f��w~x�;����wo�[b��Ef ��\�p�u������f�O[����9����7lk����ә*YSO���O����<�y$����V�By���|�Ru��������䡳�;���wZ脿0̝�a�C�����OW4R*��eUT�B�l�wZ�3'y�(��37�,?(I?NwM��1��
HS�Cs4��Cfd�;3z�~a��a����=��O��n��4�U4�:f��<�l�ݵ`{Ӛ�~a���r��UL�J����u�r�hٶٞ���T�]������ݩ�p,x�$h�Nh]��@��w��;�_��{e^L���h����'���9��8"�9>�;��������(I�3_'6�&��NX4���v��qg%
D����|�}���;�\[�DbO#�zn/�m�@wH��bܱ��0�#rh���=�w4���z���>�����$�G1);P]��ȼp�Wcs��p
�r��PS�T71[r���a �i�$���}��~]k�=�ۋ�3f��!��r)����`�6�\��@wH� :ۘ��Rѣ�RF���D�Ǡ{������_ ��  ��� � �H�$��,X @>��UP<U��y�I=��s�O;>4�#��J8dM9��r�@�l���[^��n�h�Dbu�R,�'�����舄�������f́���<��k�[O<*�θ�g���rb��	��"�h7g&�d��v�Ϯ���b���� :M�����4�<�Ǡwu���uz�e4���
���\�<aF��@;nb�l�& q~@�KeX9�14�$z�n��[^��n�X~J"%%
�+/?l���SD��73@���@�����uz�n�գ8x�+���I�Q�^���;��6ɮ:1Y�ղ������C�v�=�\Z�������������v��t���k�?S�b�s�ǐ�'?�]���*@z䘀�~@I7�����*�����t���&#������o�@��W[�4��0�f��[^�����v���EH�J�[�{���MUMM��f�X͝ޟ�{;�X��́�'�UUK���5MM
e4v6wq)�li8�L�c���6�K:�,�ze]g\�;hcv�{i�V�u�xK�I�v'��l7����;�η!�����v�y^jK/�\�t��m���b'������n��T��eJ�e�<����3��8�d��,l[r6�li�e��\7`Z�N�w>=<�R�ݵiq����a��wus�����;l6ݪ�R����yQN�K���yMl�Z����v���t���Fwַ)��M^��g���:M�\��� u�յ�EI32"����nڿ�I%���������vw]�g0�k�aS4��6�_�}����%�;�T���ة#S"�%#q�����uv�޷sC�_�|�|\��#����ͼ��2K@zM�ܓ��-��o�痭�v�<���]cl��v=,� f����]:y,ex�x�&ឧ�csm�6rL@6����'��րy���hR�U$�
���Ǜ�~�X�B�₠|?L�s9���{����=�w4x�Ű��6�y�@��u��;�ϢBo3�Ձ�{���W!��<��F�Y�y[^��[j�Ǜ�a�y��Հ{[i�抢�������mX��ﾟ�?|Ձ�mz�p�XV'pJdmIқ���ڭa gr����,��s�Z�^6MV��	��.���f��mz�n�գ�RG��$�q�����ɯﾛw�X�vl�b���"l$�I#�4+k�=�w4_����*���@�|�@����בd ���EHnL@wd�H>�������Mn�C&6�#��r�^��;Vh�ՠ{��h�0;/��O��3�|��B��ʫ�i8�z�%���S��=y�ތ���E&Lbn,������4�ՠ{��h�נr����,s�ni�۵��fgu�_wM��N�V��,]�a?��H!�{��h��@���4�S@�<��FQ:i�Ұ���`fOsVn֖B�J�$�F|��+H
0S�H݃�H�w�$��E[��`~�+S�jF�UMw3qݒ] W�r�� ��rۚ8�Y HG1�xHӑǻQ�`.Y�1�S��$���v�\;c��f��<Zn��Y$�Ś���=�w4]k�3? ���P禦d�@�Q`{۶���'>��7g=�ZX�=NnBA�A2�TҰ1�����g�Q�"��Wgu������N�R�L�R���]�X�\X���K��ﾛ�ϙ'ʄ���j\�V�kK�;�/�k��=��j��D%��XH1�h�� 1"�'���1�``0"�!!:�2���B�Mr��#��)��4�@��� �) ��@�ʮ$���)�SF7H��`��Ł��� @�3 �S��H@�*zЂFSu�`A'پ��H\bAe�S,Sz1�R�����J`D�@��H#(B��LIB�BRI8�D��1Z�h�55Ѡh$!�sl��l -beX�>S�#�1<�I!��_ ������1t��b@�
�$*1R�{D��H�'��b@�qt8DJ���au�>0@ ���	%�cL
`��b@�d�O"�����`�# C�㓕���i	!@�8�d@�RbF��H\�1!.�y�i�� M�L�:�ɤŵ�l�S�eu��z뭮��� ֐{A��6g��iX�V7(n gC�r�e��9�zнEp�6VV�Uڪ����iMkZ��C��\�Ą�W@H9����]3�InYգN�\Nr�-�,յR9�8U�|�NN��8)SN�Y���0��ٺ�;���06���zm��(W&����65�(6Z�,���ч:�G\\)+#��$TY%�Y�4vu�\�ˬ����x��P��+�=�:p�69�]�vֲ��[cp8K���ão�u�<�T��a�=*�1��pf�<��s��Ƣ��WRd�c�]6�ӞIG6��ᓜl�ئ-�Il�J�%Bt�I���z�jnYZvXԡ1e�1�D\O�E&�VS��DSv�)�eڥL�tN�� D�lڻ[v��a���D#eJ;j�H�n��K���k��8C��v����;�k�m�Gɡ�a�&ܽWc�SkbˉN��v\�b��@�&�2jR��pk�`�=:��^Ck�f\s������0myE��Z�ݶ�g]��UuV�l�.�^ɘ�	U�X<���u����Nj��RL�e#m�s��W����Pҷ�h�mml\IJ�i%���|�}~�R��l� @
�z�@0�է����S�Ż���m�� U8��Dm�bN����x4\S�@\�:��ûm��mZ�时@��[��<2e��G�gT�[̝9n�` 6�6}Is�\M�-vxwtM���J����|]r�mT�ˢڥ�qb��쬦�+U��c$���u�6�k�؝��z�Q�f���mj�;;M���l�ۖ�nN��Z��8x��v�m,O3��9���c�+�ו��d���X�D�6�:��DO1����ӨQ��+��Cu�ZNr8�Ի8�"�j�90A�H��D���4[���.B;FO��}.�l���y�p�<��tjۥ�;����9&�[���rb���T�@��Qڃ����0��DQ�vf�<��2fm�&�ۘo\2;�t3X3�3:���b����l�U<��U�;,�b��'�(v����8�z���ʺ[<�j�92�G1���gu�.�3�Cmň��1� YƇ6cn�)��x<��Y��n�ՠ�¦�cn|�Z���GA�=#ׄ�m��`���h����K�{n��vGn�8ml�v��J0ݳ)�W�������U�?_ ����f%�0�H�r<���g�n4�Yz[Xl]���$uvSd.��ZvCb�����߭X�vlzwZ���wW0�o)mI�Ni�3J�Ǜ��Qi%�7g;��ݵ`f��=*��rN���=�j���i�K��4
��=�;&*G"O�$���@����n�˭z��Y�^�'�u��NR�n�����z��Y�z�M��%�+�)#Cȅ!�3��vɌ�z�1�u�y��t����,�zܳ�v`����9u�@���4[)�~�S@��Ű�DLBy�zv}�s@B�A$XF@ H��A����{9$��og$��נU��e�$ۉ�'�4[ ���u~�Wn�L@7�] ;���(L�`�!�~�S@�ֽ��aТ���Ł�1��[D�K���ͤ�& :�H�`��{��?=����lԌ#^�죃=�
���f��:��h�Nc�����qɞmL�j�/73q ��@t���uW�X4�z�vLTRF�ș#JG����?nV�<ݛ�e_BP�l���?��!�H	8h�ύ����;DEB��u�*������f������f�˭z���@������@?{)ql"�26�F��<�� ������T�w$� ��ٗD�pӪ�&'r6힗����].{�Zvr�n�6OV6)��Q#cD��4�`�}"��& :�H�wun����H��޷s@�mz���@��Zp�-Ɩ9�8(�73@�d�\s)��~�s6Z�e��q$�#�q��+����Z����8S�'5��`~���T̵$iH�@�v���M�Z�~͕`~բm7pUU74�5Q5$9�,�kV}X����öx�}m�q�5=�]�8φً8���@z=�ۓ�̧��~���U�v{��4F��E��h��|�BlכҬ��v�����妧p�$ɉ��ӏ@��4Wj�?^��9u�@���uC�"��#��IhG�@;rb�9��Yi�4)K���¦���ݵ`zFKݞI=���rI�s���x�~"�� ����BY�P�9��e��H�]-��.��r���t�t۰I.�t9w9"�N5��g�1����m����-�}Scn����� �;g��@kr<�e����,l��sn,<�Х�V�Ick<pn�v;(N#p��,벥I�l�[@%q�N�m���A9�6���6;v�v�3��s��s����ݑ�Qн�rZ2�^ez�����w{�;�ܘ(	���&0�HL��]�Sn����z3Xr����=�n:�9�IMn����nɪ����-4�>��<�6U��e?�����*>WĎ4�#psS`y�l��	&��,v�<ݝ�;&*)#b��#���h�`���Uv�$��wp�d۶ADH	Hh�Jh�נr�uz���;=Չ��Hb�dR.��r�&���s6�λ5s��"]s�DhN��u��u�9���q�t�rkc1v�1Ƹ�]p�dg���r�&� �E]_�z��I�rƧa�6U5#�E�����%�_�V�{ʐ�& :�/�å���>đ�)��nh�נy^T�=l��Py�B�H��f�ˮ́��u�ݭ,9DD'���X�{�ᩑ��Ǡy^T�;�:�M�n�˭z[��G�o�D�R�a���h��ls�MPM��-l��,mb�oac�$f<��AŠz�M޷s@�ֽ�ū@�DO� ��&����i}	�^�M��y�`{v��?g��5��MŃ�#��9u�@廲��ߚ��%	z"6=[�VX�\X�K�aI�ܙ�@�my�z�M���9u�@���w �$I.���ܤI�@yȩ �Ɉ�����xt0�I$�0R�p�՞�4���6�{[�3��V� qv��]�a{��EHnL@u��H�ՠ\Y�r��s�Hnf�˭k]�|�Rǰ@{�T�w.�\2�(@M��/uy�z�M޷s@�ֽ�;&*G	�	1Hґ��By�|X�֬y�6��J&!D/B��!&�oeX�FTmP�
�T�u��ܘ��e :M��߽�߿���q翼�k�*NxD��q�Bʽj3������LD�C�k����.E�\ɛvͰ�����b�9���6�*�=��)1LbrdN=��y�z�M�n�˭{�E_"�� ���	��J�3���3۶���׽�`r���@?rKaB4(4�)��OR�I���)�l��Ʈ#$J,M��9u�@��j�۵���fڰB�wZ{Κ�4�N6�v�KÌX�f���sUV���Y.2d89��9��c�bՀ�<�%�:+t�u����s�ʏ��wn�9�1�XM�����3��=���w�q�skNx�;���WWT��u��Yy�k��C�$�Z�!0LDJ�u�����b�6�6ϓ<pxv]v�:�c��cH����md�}���8���=�7B�n���{������'AO��ߡ�	�B����6�θ��&ޝo�.��%�j�߁����h��K��6J� &�t��,�=l���u��9u�@�NɊ�Ħ"LRH�Y�z�����m}�{�6�{��74eF�&a##�4{��˭z��Y�z�M��MnH�p�4��hܘ���.�&��"�q	W��Bbi92'��;Vh�S@��mX�vlQ�oZA9�D�T֤����
/&�)�4�yMӍj��]�.�^��9B�&H�8�Y����{��h�נ{�՚��X�
�(��{��EHnL@wd�H�`�����q �Pqbnf�˭z��M��h���b�c��cm����f��!I�@wH� ����옩#�8���h�*@;rb�*K@:�p����͆B.˩������tv9抵�K9y�M*��h�N��Q�A3	1�Hh���.����V���Z�Չ��x(�#��r�^��;Vh�ՠ{��h�K�a$���rdN=�v����{98|#��-l���5|D�<��>��B<f$�`�V�Ry�'���"V��H��} ~������I��5>P�C�!�����a�� ��@R�衇PU@ z"?(�(�N��֬<ݛ��Kbh�Uw[��t��6� �1��/4�$�vT(�N10�-�빠c�ٰ?zwZ�=�ZX�B[��7-�xflN��gD����6��� Z^9���i��7����y���ud1����~�������l�*@:�N���m��6��=�w4[)�{��h�נ~�d�H�S#P#QI����=��VtCz��l��V�[*6�XȦ9�޷s@�ֽ޷sC$�D(͚����dd�uS.���ͤ�& ;�T��"�t�����=���;�ܾ^��ݖu��Z6ۖ�gI8ڑ�m�B��ns�+-Y��*@t�R�EHnL@;�v;� � ���z۹�{��h�נ~�����Y��(�G �M�s��ܘ��H��EHa�f�mU�Tԧ3Já��t���Z�����s@�T�tqƛc�Njl�ݵ`t([�ߗ�37�X�w9$�O�#�*�H#Q�D�Gs�l�s��&�nL3,�ݺ-�����CAU���6�n�kM�ca��Jg&�J�ɖ㓝�չ�vi��Z$u��]K�������:D]�`��#�4A�c���^�k�V1$붶z�:Dq��p=�}}<�1�f1iB� �tJ�=rN, ��g{=3k���Y+��rl�ݱ۶�j�v��:�ͮ�����@���7�X����>�w}���:}��m�L#4�%m�v��qӆ����Yre{Cد;c�����<Zbq��n���0>��s��䘀�K��u���/� 9�3@���h��@��w4��h�W������76�䘀�H� 䊐�,�=�-�r)����n=����:۹�{�w4Vנr��v5�J#v�sv�H����& ;�]��~��������Tų�is�F�K��=�+��z\��s����N;]�M���б�v^m ;�T�w$�t��H�@��غ� Ј���������@�@� ȳɟ��9$����4z���g�qc�6�
'��R� ;�T�w$���j�r&H$�Rf�b��@=.� ��ۚ�"Y��c�s4y�HnL@{���EH�tiS2�}���F+8w*$rlf��K<�ý�WIԹz�ʹf��	qlٶv��[o�}� =�`��"�s��].U�1��8�޲������s@�ֽ�Gc���dD�d��@���$���xr`�E �bA��$`BTJ
QOH� ��<������y�߸rI?g0��F����{�w4]k@{���EHW]V����.�ܽ/3i �ɈvIh�*@w8�~��������[f�aխ�]��g������b�W��n��'��<�#ٮݎy�h�"���s�{�T��"���_W�%Ͼ��&/�"qD��9�����fڰ1������V�6TuQSH{���H� �1�qR� ?{vGn�	�h�TXr�J���=�֬��V���K!Nd֖gUql��#�n=����:۹�{�)�r�� �rk�rDuP���M뉥�u����0f;N�ٗ���ͳöH��b�Q% ���u�s@��S@�m~A�|���X}�bQ6�{���{�& =�%��R��b��!��25�4Vנ~�hm��=��;+��\m���s7� �R��䘀�;&*HI�G��Rf������M����n��YІ(�&	�\l��5�g��s�mVφ3�%����CM�Q�����L��/�nF�,M4�;X�g���xS�fՃ�X��'v2�lݤ�d��]�/aշ�{Vmc��m��X���%�ז�F�b،HY
�v]�;*h�cj&L2T��U�cv�9�6�Ԕ�	�8�'wn�;]�q��Mّ9�k��^� s����J��л�]t�~�{��c}���瞼���&89�V�h��-�و��o��&��2:=�[7���+7/6�	>� �1�{�,�?z�-Q p�ф��9[^����Cg�w����j���,/k�j)�Q8��v�����;V�˭z^Gc��2"A'��[����-��b�9h���J��L�8���;V���^��}V��[��Z�0N�H�I�����On��UX���H'n6�]\�c�vH�p.���h�b�"qŠyzנ{�U�z���?s�h���\m��#`�q����EP�j ������'��{y$��k�=�b��9�'#qh�w4��Z/Z�s�uA?��M����@y䖀w�b�9h�nh��Z�@�&	��E�r��@�Z���y%�=_�\���M\�a�����r=t��\L�,��Ҿ�qcH�"0Jb�m�H�$q��s�T���- �9�	}c��G��� ��@�[��~�j�<�k�=Ϫ����.)�17$q9��v��۳g	BZ���;����`bk���8��8�/Z�s��vՇ%����Y+���́T*jS���<r��*@y䖀w�b~1��Ǳ����[�C��F6�/���xP�S5�ns��=�7i2zK۩E�l��hG <�K@;�1��rȌ��jA4�h�ڴ^��s�h�]��z�#r(�8�qd�m ��<���*@s�-�����1L�F��=Ϫ�/��hO>���MD>� A5U8��G�F�^z/"��R4��@�봀�=�_9�v9h	�h����a�$�])n������Nvl��E�&'r���v�x+n�zv���-]�m�_��� %��c������V���*�t���f��J?�d͟�v��nh�Jh����i1�Ǡ{�K@NqR>��v�߄��؀����Q*���u53N������ͮ,~͛�!$����ӕ3��r�#Nf��t��W�����@�fڰ6#".	 �!4�I�mY�"H�
 H�fBBZ��e�ecBH0 BA��O�ax1��TƄ�9HD�f(m,�@J�a,*ƄjZ�T�!V5`D���D< ��@�V�#FH��
T!i-A�`ċ�8� �!P�(�	#�� '��IBe`�B;�B��@�e�!���	!�V�@�$Ď��b@
0(D�A��������r$$����JH�)
��t�a ������4gx 5��$
��0
�c1 !(0�R�����Y�$r�RR!�AI�4C@�D��Z��}$�$Ǔ@�)R�hf�Ot�;]�ߘ 6����6���![�97W�k���ϸ&�UH�vp5�]Fk=����R/mЙ�O/	T�qJ$�͕m9�R�ڪ۪��g*���Ҙ�O7YHc#AV����8�`X��$�4re�tʱ��m����]���G7f��:C��Йn��Kl���uu�+�W,%n{f�N�˵֙��{iݐ�nh����P�82��b���Ê�k��g�*WX�Q��pi�m<��v�m%�m)[D�`���:���Y�t��6�8�v��nH-n���[m�ѴU�]��j0l����lb�����H��d��c�5t�ԛ(��V�+�K�m-7��
v�]�fft@k�5�d�`��&��k�����w+�Խ's���c�8s��"|v�l�2�R�g�m�ۙ"h	��t�.��U�z�
���	(���鱸�\R��e�f��ĸ�"z(�.g���4�g�۲=�kշJ�8z���.I�a�i���l�]�x�n�5���+O<���W;.�7OL�;P�+F�]�R�K� N���rE�F����v�k��*�UJ�N�����᝱�N�����Zk�P��6��{im\�		�mq�E�N���o�r�4]�`	�r5�rٚv��`gjk������4� V��(!J��C��˥+n�\�0F�]%ĺ�mX�˰2�CT��w�RZ�pxds�3��PSnC�ץZ�������V���,;��jr�>��bz�����P-��[4J�7npnZV��q'jb�p�r�; ��^n���zۗgPl��*�CP�#���r���k����K�˷8����I�Y�&�8�/h��掉bu��zD��Ȫ���*��h͞-�Œ�C�LۙS1�	&x@s�J&�|��1T��R�1-��j�P�V�ء6݋iN9�YrМ#��L�)�Ɲ3p��eĘ�Z.ά��$t������DG�� *"|�: |'���<U@�At����� qV�&Or[9��]��.���۫<��1��J��%�f�ti��齷M�p�z'T�m�wi�[��q9煉�e���8ԃ��۩��ڎLv�ґ�չӳ����ru%�n˭;��:=�0��;]t�Yڲ�cN+Nm[�S�۝�u�ƹ�-�M�E����e�5��ΰ���H�����Ŋ]�u�ѷ�Q�K�g�簠��Vw��Eu7a*�zwa��I���Ѻ�p��<��E�0�P�Lcmm׭�[m���w{����qPT�UQ�s��?{kK}�k���0��@�}�`�I�d�G����@NqR����_UW�%�d���"$��Š}�����M�uz�;V�~g0�b�Pxԙ��D'��Ł�7�����v�!�o~V���O��<����h{��?zw]��͵`{�ZXD(Id��ÙGL�9rݹ�̽����,E�F6z�V���������mj�Ó�~eP׫�!�������耝"�s��X}n}����m����5SN��fھ�P�Ji(�P�$�!(]	B��~�+�x�<�����u��r2��j1��h�Jhfl��߲{����j���쌵NduT2TX|�}9�6d�;}�j�����ߍ�_b�7���ɑ���=�`tGf���ή,~͛6`��۳Uud�b�����쁛2�U�nYMWE{8�l��r��r���V>�~~���+��������!(_�fOs�-��#�n9�I��e7䏗_���=���Nk��;	M=�&K�2�����9�����>����$��I4�(J(��`{z��5zV�ڧ.f�j�Rt�âP��wo���;���������LV)Lc�����%�>��_��@wc��u��X۴��!e�#�cbAǋ�<X�E�N���8��Ӓ��g�L�}�.Y��߯�֖�͛ޜ��%��d�;ٽ#-Sr�R�S"*��5�l�BP�fd�;�{����Z_Д6f��5J���T��������9(�(�3��|h����r��)1��rc����;������1�l�RP���aGD$���v��d9T��.iԓ4��@;nb�$��Ih����}�"����3bt�^M1�W��kG%f�=
í1��tsZ��w���8��1���ֳt�>����v9h	�%�=�`���q7$��L��q��o�3?�3�
���|��&�~���oM��q��Ґq�̑9#�@�}V��YM?�|������@�둕��mH7Zt� %���r��af�I�&F�$��W��޷s@�y������F�	�J��{�I.#Y�Q{rs�\oAg��"�ٛ�kf!-��M�XN�bQ�{��ֻ,N�����{%�덶����[ �:7ܜ��\sL;��n97:w<�۬v��+=��-\�Sֶ�lVڍDְ9E��ʝK
�qۭ؞'q��g\n5�ܽ�SN�m��A��B'p�t=���pn�D��u<��V�a5u@�<�:fn�i�f��?���Tѹ���y����CL�A���3n8tx8�Ke�'�#S�x�&<Rdm�@���_Nk�=�:%��<ޛ_3z��*���.�i���w���\X�zlyڴ�{9�FD�'���z���G�~���'c��󬫫`�a��I���s�?Wj�?/Z�z�h�<�뉹&92d��@�����b�l|� %I)����j�;5ĉQǡ�2/#�d��NWEl�؋��'/��4<R)��c�C@=z���������_�fuq`j�*N���1L��h���ؑ���z�� ��7����x�ɑ�	!�T���%��j�l*֙�$ɋ#�q��Қ��h�Қ/Z�U�E&7�'&	��z9��@;�1��- 8��2�[�3j��i��6zWkgs�SԸ�֎zqbz�;m���u�JY��߯��`�w�bݎZ ��9�Uչe��R)��f��1�l�(�����v~�M������qqq��nHǒc�.nrI���ӒI�~��AA5A*��e����IM�^���&+�LbmƣR׬�?z�h�W�{�ՠ{:�eq�di�d$�@������z�e4�Y�w�PĘ���<��Z��D�@9�5�F�M�{T�A���x3�Q�I�N1"�c����9^�@����u�4z�h�\[��4����=�/�,"d7��X�\X�6o����&�|�]EU'*jf�T��; �ޫ����舄�	F�oM�J<�����~���� � � � �d��Θ�mٙnn�A�666?}��� �`�`�`������� � � � ����x ����s�������lll~�4���m&K�wnf����lll{���8 ����Â�A�A�A�A������ � � � ���~�|�����פ�ɟ�&n�0�3��]��ˉ|<�M���'㫡v^wM���z��3S��x�~�w{����0�`�`��߿xpA�6667���x ����ӂ�A�A�A�A�~�����lll}��8_�wr��n��sN>A�����o �`�`�`��߹�pA�666=����|�����~����
( ��A�A����O�.���6f��A�666=��?� �`�`�`������� ؃�	r9���Â�A�A�A�A���o �`�`�`��������%��nXMݜ|����s�߳��A�A�A�A��߼8 �����>A��C�A��{��?� �`�`�`������lɛ�vᙥ���|�����~���� � � � ߿w��A�666?}��� �`�`�`��������lllz*ƈT;�?�ٞ��	s�kg�s�.�gb;p�Y0����XKv&]�*fWUZ�ō
)��d�cٸ�u�.j�{c��cuVlem�n��Y&���]�XѸ���5������l9E��A)��x��z�QM���0��`4�cv4p�nn�*�8�UtYn �\l8��흙�$���6�'v}cm�==���\[K�R���;YhƲ���l��u��VMy������N�u�jG5)�l��Vs�rZ���my;\nt#�=����]Zc2f��r�?A��������A�666?}��� �`�`�`��������lll~���>A����'�L?2�ܥ�sw��A�A�A�A����8 ��"!�A� � ���g �`�`�`���xpA�6667����|������){?Y2]���۹�8 �����>A����~����lllow��A�666?}��� �`�`�`�ܟ^��6�n�L7rK�78 ����Â�A�A�A�A������ � � � ���~�|����s�g �`�`�`������ۻ�\��۹�vpA�6667���x ����ӂ�A�A�A�A�~�����lll~��?N>A����ߡe?ao��ݹ��=y��{8��5���Ε:�3��F�F��z;�M��ݹf�&�.n�A�664���:���ޛ��������V,ޑ�l�:�EK
�,{�7*!(���A ����[ɜ��m��e4���܍cne�n ;�� 8�;�� �9�U�	�l#��Q8h^�@�����sf��	�u�`Z�tS&*����n�;�� �9��@9�����؃e�۳Q�pF�pޗ�����g��mۤளZ0��Rl�N����u�m�gt�jD7!�
��YM ��4z�h��c�'�<�&(�z�e/���7~���́�q��Ӫ�JJu47N���ڰ=�,ȇ�����BI"FF2BH�H��؂	�")�>?�)h��X2�18��XOR	H�`������V�$'�F�d#"ɼ`p[���>"F0��F	F"~�	����q��a
�A�`Ă�� $�h�OS�N�� ����P��O���)�<�rI�{���xw�d[UN���R��U��<ξ,{�6�n�z�4g��P�R<#A%<͛�J>P����/ g�}V����i�,� 	����lx�j�	�����6��t��(�+݁��7o&���Z��۽��t�������U~��WWȹ���1�1(�� ��P�`�v��t�����밁*Vg���rh�O����������ǋ�ō1H��49DBy���ή,ٻVT-�0�B�@>QOy���rI�{>3�m���,�����@wM� �&�;���$�������������x�%��ιƍ���Ƥ��b����2�k��0:�绻(\?K38�5!����4z�h�j�=�)�~��3+��jL�rh��@s�-�6�����0�����	!�{��@����{���e4����QbnGZ�d95�6y%��M��[n�L�R� �nՁ�������������!(Kp��顶T�Z:��2;Д^�^t���,kn�S��`K���oF����ɭ�jx�<{/Gct��KIb�4m��u���,M�nx7<�6z� r�.Ѵ�[b��۞�7X��3p��Q�JN��Scq�T�`���y�,pc��ov#e@͈ѷ�j컂Nwdy� �f.�[���-b��vS�U�Wm��Y��3������_��݇�+T�l�pVI����z3]�8��k��Ocnŷ�V�l��]�͹Wy��H���$��l95�ǋơ�1H��4s�h�e4�l�=�߳�"������$��qh�ƀ{��|�u�W��@��ĝj8(G�Q��%����y%�=�`��6n3tک�*�X�V��}������W��u�@���13��ɑ��ś�K[r�:F62��g�c5ɵ��n�C]m"�P�I��Z�YM �[4{�4�܄�mbnGZ�{����*� )� �'w���'�gƁ�v��Ge�5��Q�Q� �nՁ�eig%�͞�`{:��
��.ǐi�$��=��=��`~�֖�Bo7��j����M&�fj���,d��ξ? gwU��t����ēxXbrG$�&LюM���Y����/#���}�Ε;��C�5��i9������gW�ݫ����3�_�-�|�6��dyy���j��䖀�H�}����vuZFg�H��a2ɠwY�w;V��"~ʭ,ۻV��dr�%:�Rª��Jݮ�`{;�X�v�{�4N.-�qȣ�܎8�޶Հ{wj�����3'u�ȍꃐ���٪�Ёx|���qg��l�ݱf��=�g�*���{Q��v��+ĕ߰	�����@7�Z�6��j�ܪ%����X�V��	Blݞ�{���l�?v<H�P9��UUd������B����Ve��x��#����qh�e9$����I=���䞯C��z+0�J�Dz_���٭�n^�U*����]Q`�v��B�������޲����9?���(�#Q�`H ��;-�v��:!sF��ewMi��rL�X�V�d�����(I|��� o�}V����
t��:aUE��;����,ۻV����#�DL��bm<X&�j��|h����N4|�Z*��1'�<Q� �&�;�� �Ih>�U|�_��1���2Dܚ�Қs�h�kK �nՁ1
�Inٲ�L%�'6ڵ�����u�.$�c�\�U������0�&N�:��.�=�h��-Џ;�,�]lա�7��{m[��l��'�����m�a���kJ��J�ٹ
�v�V�M�۳��"m�ɶ�r��]�,�f��ݯ�I���L�+��M�'�<v��s�W�����dP��m�KN�2km�	�]��<f��vzkU�����|m���g�4�^x��x�f��mz��i�Y�����}=po����u6�t��O���M@w=�����#���$�@��)��f��t���v��=�%1&���E2�j� �����ϡBP�͝�`{:��<���[5EIT))Q3Ua�(Jۋ� �O���&�:�L/�&8bL	!�{�U�~����v�{+K��&�ˠ��n��*�#�a^��a�V�tok���;c�jKj����:�A9��'#�/�{�����=��-}V�ʣ��$�1'�4�I�Z����U��	1�@{�� P�v<�1�84G��t��k�脓y�\XӼ�ڥ6c�I��sM�U�!'�[������ݜ�`{�S@�y\u����rE�{��.9��@I�ZSu�L���5i��	�5�x���\����]�u�PƖ�6���;a�m�a�H���s���1�@wM��r��`���[�$�q`<J8�z�h_U�{�S@������=A&8bL0�l�����\�.]	z^�(��b��WE�?!������'�����8��ȦG�Iqh���:��@������Z*��)$�(�4���=�)�u}V��YM ��r�rD���d�dq�vx��%�:Z�#��˥�^T�7tE�.�c�\L5F�u{�h�@9�Z�l����9T�E2$�$4���=�)�z�޲�^J⬍�Ԑ�-޲�׬�?Wj�:��@�rSj��9�&b�C@?u��6x��U�~�;6K@us�G�H���'&���V��}V���� �����7�_��x�
d��F���)a6<Խ��]�Pj�/Xg�Ei�$�@�>�@����YM��Ű�Bcx�����9���uϾ�<����@K�vM�J&G��������ڴs��w4���qG��D���B~ξ,��v�fڰ�'���5�E_!�dS"��Hh��h��sd�_����~��I0�*�F�"��)�H� D@C��C,!ARX��)%���E�j� �R>�0 B+�'qM4���4# ��@����o�y{�H}��L�DBp������}0M�X0~�� ��F�������#������ lYd�mn����Dݶ���q����d23�� EȖ�-�*E��F�r��բ^F8 �r�6̈́8"�t�K���񒺸<��I�Y��{Hvi�f���UV��7=vIju�L�oD,�t�/Z���z�6ñ��J��ss�u;nɊ�����d'mqSқػsWm�1q�j��eF�ؖ�˴'��I�䥅����U���Z�
lwVb*㥶r�lnY��i��v�l���S'Cs,v����vbB8S/V6{a�Y3ٷ��=<�]����^ٱ1H��e˪�7mt��N��an�`�#rf,j���lG�&���m�����n�r]]�dzՒ�a�N줬�9x8A�4�U��M�v���.ِ!���,l�qH��Yt4�.��6��m��uX����,;n[h!5�t�1�9Kf�ܝ�[�B!� �(9뭻]��:i�˭�#8G���*Fu��hz������N�z�+;-�Z��l��2�\:#vOon�K��(�z�Y5��i0[aE����"�V�` q���&�l���i��ʮ�PZ��lO3�͹�t�间\�Өy��T� &G��We�X3�sCZ�XI�K���J�N�E�\@ s����4Wb55�Pl<xB�8�e7j�ZBSwi�"�n��&�ng��E�:���^2v6�ܔ�E�,s��S]O-��n��V�BzR���܇IoV�n6 �Kn�^K�fz�qt����.&���XHj�n�e-��E�b)+L0��U�s�\�Njz�ϱ�G�e��c7U�bM�����9�I�9��{����ֻj�rYpK�w��Ͷ�sc�6���P�@A�^L��:SB��N��L�eYF�z��3U�e#Ti��,��ny�sY��!�;,KK���*�H,:89��Ns�jqBN�Gvnq��kn�Ɯ�r���v[b��Ǜ'X�GQd��.�3w����*u^~\�!A9���!� >tT�x�z!���=�˻-vkl�;��l&�=��פ2Ѝ�y�*�ڦ�Z.K:����)��O��z)�9YS��s��O&4���4�p$=��M]m�l��`c1Ůj���/nuvE�Ե��ac��]j����bӰ��^	�p�l0�=rN�m!�퍞Ռfݯf�vn�胂�����=��68�3=7,ln�l�@�Z���sѥ�����׏<��ƙ�	���6��nb�pt�|�1�/&���䓵;�:@qFF�ț�rE@�n��u�@��:_�f��=��NI�n�&I[��H[��@s�-�qR��M��j�:jj���*���ͮ,x�=�*@zܘ��I�������UQa�I'�[���oZ�?<ݛ|�!;,�9;U2ʚT��u5[hs���7��s����Z���Üz�5"�I��`�k�ܜ��y���wk��9���;���w|o�.�]���76�	���s� 9䖀�8� hb�5:�d��$*i���w�DBł1T l���גN���I=�+K�(I6kONa3R�T�eUM;�}��9ȩ���@;����q�$x7$Z�u��=�)�~�V�	BI�k���e'$��7J�$��ͤ7�@{���Z��'�(��?���%񻻷3ra�eݎf�d��7X�i棬9ܓ�'<ɋRtY���;����Ӿd�cp�!�:�?Ɓ��V���)���szՁ��ۡ9US�UE��Z����=�`��UU~�)�-�$d��G"�-�~��;Ϫ�t(�B!ry����'�ϻy$��Ȳ	�I�q��;�ՠ~�Jh��v(��DD)�Ｌ���|�fl�6��7wP�@t�-�qR �[4���I"��%Y#s���ݎU�Ӟx
���u�s�#!��ӻv������۞��P8�)�F�I�w���޷s@?fm|���=�\X��O����d��Ff������t�j�߄�9k��=��Ne��TM"�U9�`��;���Z�6�n7w34���@w=����ls��QU;}V�wH�М���r"����-���=�`��H*.�j�3s�Şn�|�A�����g�ₜ�5��/n�؛����jq���m���� �sP���UzæO�/�uP䪕.]'SUE�~�ڿ��Jg�k��;����/�M�͓�J�R�,ͻ��9�<r��@nU��1d�a4�:T�e�TX|�"~�>�9���A�UW�/��w)|�Ԑo$x7Z�t������^����k��Nk�-BI(�P�HD!
�,+Z/y?Oٓ�i&Y�Y9����ݻ]���:v9����͜�.ٔe��f�/71r�Ş,+q�!���ư�u�����4���S��`���h�s�=b9Sx�i�g��s�N Kkal�2ۮb#`�f�v,�n�rm۱&��4��ۘ-T�ݎ��icv��c2&��yc�n�:�S� �8�Yc��1���w]��k\�xb���!�]u������n빻�v��ۨ)s�.9�<�$���-j<�k:,o0�[��Q8(�d?�R���h�Қ�}W�33�u�u�1}2Lm7��D��x�=�`�<���*��t�nbYU1.@������?{+K>K1#��4u���Ź#��Y�/6��@nj��>��W�gנU��A2G�������h��x�=�`�q�^@�wXk\��ҹ�j:h���^��aqڱ��u�N���B,�Ȉ�Ơ&���t����-�{����s�@K	S+�3qS�5.e�TX�9�����Q2{6�4�}4��M˒�W���
��ʹ�������w�o��_���/d�گ$��E�"����h�@y㖀�=����\�ݬ.�9�SU`~�V�(��mo?�{6����h]���.0N8�A&�x!tn���z�lf"������rG����h���s�^�����������S@�8��$pq�$�$��?z�_Т>P�)��������?d�^���&5��1�$4�����M%L%�";�RQ��l�������ּ�e��cq%�5$��fff.�W��@��)��f��;;,�dm����K@{�� s�P�`��~�ͱ���jj�:��CoEujT����G���յF8ݴ2����i�����^��������T�<��s� 9�@�܉���M�`����u�{>J"&M��͝�`~̥_�Q	���Rvd�I50RI�w�Ɓ�}V����h�h�Z���I���0�(P���N�������V�7j�a(�I�QQ�Њ����O}��w$ps�q�����h�h�V��s]��]��`�+����UM��r�{���#�y�0S�\�茁S�?�{�0�j6A<��C�9� ���{�)�{��@��w4
���v&эĖ����@s�-�R �&��3?�*��!Ʉ��ŊHh_�$�EH����{�w*�f�eɆI��-����{���ҚdD$�k���e'�R��&��UN��rj���K@{�T��WBcg�+<�����WMs������;u̵���P���s�*���u��h5�����^in�z��X��ܦ�Ӷ,4�c8ڑ�;N\V�Ӗ���֎xz��}�}�6�[g�s�s
�q��f�ʥ��D��<� 唐Jr�7&K�uY�Ua�&��W��I�c�h�@��9�'s��Jn�n�X�+��9�^K2ݗvL�Cp��IsL7|CNo8�i�E��ytH�<�c\ u��b%���58���ʕ��̏%&8��0�"I4�>ؖ%�b{�����Kİ}��h�&D�,K����O"X�%����%�a���r�7vD�Kı=�����Kİ}��jr%�bX����yı,O��6D�Kı=����n���)�w7sv�<�bX����ND�,K��{�O"X�a�2'{��"r%�bX�~�߯Ȗ%�b~?�o�Ò�m��^ﷸ��{��}��Ȗ%�b}�y�'"X�%��w��O"X�%��w�S�,K����I��.Cnܛswx�D�,K�͑9ı,?*G�����=�bX�߷���Kı/�w���%�b�~�o��~[�3bt�|�1��z��X7��V����k,n�n��֮6ztf��MK��'"X�%��w��O"X�%��w�S�,KĿ}��Ȗ%�b}�y�'"X�%���/M-�k7]�����%�bX>�{59T$@�R�u��4(+��5@Oq���O�X�����O"X�%��߹�'"X�%��w��O"���2%��٥���nl�m�ݻ�S�,KĿw���yı,O��6D�KȀ�ș���׉�KıFuqP���L��_���s�Ԅ�)��&��Ȗ%���ȝ��6D�Kı>���x�D�,K��f�"X�%�}���'�,K����%�fB��s1��"r%�bX�����yı,{����bX�%���x�D�,K!fm�B�!2!}ڭ�h��UU6Z77��0ɳkDp]v�K���E]�t�Dtl��zߧ��O��͚����~s�g��u�������bX�%���x�D�,Kﻜ"r%�bX���v�<�bX�{��7�"ܷU�w��oq��K����<�bX�'�w�"r%�bX���v�<�bX����ND�TȦB|k6B_��EL�U��Bd&Abw���'"X�%����oȖ1=HA@��pb���1R*2 "��Ѥ$n�H�+@4�=z@��O�"������� 0bRG���S��		Uѐ��S"�x����� �N�x�?(*�U�_QT�*	�b}��S�,KĿw��'�,K��Iӹ6���ws0��"r%�bX���v�<�bX����ND�,K��{�O"X��H[�����	��g���R��&鹛�x�D�,K��f�"X�%�|���'�,K������bX�'�oݼO"X�%����)�~̘~��X�i�-�Y0sڜ��6����4�N�[� �m�
c�(�-��׻��X�%�}�����%�bX�}���,K�������ؙİ~����"X�%���8[���&f�n훻�O"X�%����9ı,O~߻x�D�,K��f�"X�%�~���'�,K����%�a��w�f�9ı,O{�v�<�bX����ND��
$2&D�����yı,N��p�Ȗ%�by��t�rni���价��K��RA��?MND�,K��߷��Kı>���'"X�%�D"HY׼��!2!t����[�e�&m�٩Ȗ%�b_��w��Kİ�D�{�͑<�bX�'߷��Ȗ%�`�����Kı/}� ^ߝnYj�]@枔Kڄ�Z����ƒsN�޳6��pi�-��m���'�,K����dND�,K��ݼO"X�%��w�S�,KĿ{��Ȗ%�bw$�ܛf]�7s0��"r%�bX��~��y�?�P+�6%�������bX�%�����yı,O��6D�Kı;�����˹&鹛�x�D�,K��f�"X�%�~���'�,K����dND�,K��ݼO"X�%��ƙٻ4�ٗd���59ĳ� $������yı,N��p�Ȗ%�b{�����Kİ}�xjr%�bX�����;�d3vf�ݻ���%�bX�}���,K��@#��w��{ı,�~�Ȗ%�b_��w��Kı?'��*uP:�U]��:E�B��< #�0Y�S�	�n��B\��P��&i4ܳ���m�����'X��{W�n{vj�l5m�S;Gn%0���/#�ۙ@lWn�sn0#��Vo������j��[;N�k���92��T�-��-�v�q�e�� ncrv�[@F�܇���ʵ�45��ۥmw,��b���u��i����ɷ	� j�n�6S0�\ԉ�
�_*�/�3j9����ɰ���c�����3�]5+ڭ�ߛ�oq��'������%�bX>��59ı,K����?�	�L�bX���l�Ȗ%�b{���_3tܙ�3l����Kİ}�xjr%�bX����yı,O��6D�Kı=�����C{��7���~W
Kq$�{���ı/��w��Kı>����, ���;�~�O"X�%����U
�L��L���̐��2\�N����Kı>����,K����oȖ%�`�����Kı/�����%�bX��:w$�n훙�]ݑ9ı,O��v�<�bX��R߹�jyı,K����O"X�%����Ȝ�bX�'�{�q�vBfnՔz�h�F�9��9�ut��bì���h��Y�-�]$�M4٦�����%�bX>�{59ı,K�{��yı,O��6D�Kı>�����%�bX?O�)�ٷf�6Hn�٩Ȗ%�b_��w��/���Dqț��g��bX�'﷿�Ȗ%�`�����Kı=�ㅸw6�.컻v��Ȗ%�b}�s�ND�,K��ݼO"X�%��{�S�,KĿ{��Ȗ%�bz}{���[���f�sH��HL�BRBν�p��	���:��9ı,K����<�bX�'�w8D�Kı<�}:_3wdɛ�d����%�bX>�{59ı,K����<�bX�'�w8D�Kı=�����oq����~�q���i��j�r$m�`�krŜ�b�D�(E*")��Q%H�'B�n]��nd��\��]ݚ�D�,K��߷��Kı>���'"X�%��w��'�,K���٩Ȗ%�bw��&^�)��6ݹ��O"X�%����9��DȖ'߷��Ȗ%�`���ND�,K��{�O"
eL�b~�?��.0���ND�,K���׉�Kİ}��jr%��'���ȗ��{�O"X�%��g��bX�'r}zgI4�vM�m�ݼO"X�~ d�s���Kı/w��<�bX�'�w8D�Kı>�����%�bX?O�)�ٹ�0�$7ni�Ȗ%�b_��w��Kİ�F=�����Kı;�{��<�bX�(��d&Bd&B�%�14���P�=Y��4�ll��q<O+༗I�E����G!�M*�3�����4�W�����{��"w���ND�,K��ݼO"X�%��{�S�,KĿ{��Ȗ%�bz}{�����t.�74�Ȗ%�b{�����?�9"X?~��S�,KĽ����yı,O��p�Ȗ%�by��t��t݆�͓woȖ%�`�����Kı/�����%����;���'"X�%�������%�c��~?�o�[���n��oq���D�����<�bX�'{�8D�Kı=�����%�`��@�� 7�o|�jr%�bX���>�3�d&f��nn�Ȗ%�b}�s�ND�,K��ݼO"X�%��w�S�,KĿ{��Ȗ%�`ߺL��;!7v�nH�bۦ;`ȍ���uU 7p��a�9�H�����q���]]�&���oq�X�'߷��Ȗ%�`�����Kı>�{��yı,O��p�Ȗ%�bw'oL솒nɻf�����%�bX>�{59ı,O���8�D�,Kﻜ"r%�bX��~��yı,�Ɣ���n�$���59ı,O���8�D�,Kﻜ"r%��!�2'߷��Ȗ%�`���ND�,K߾�-��d��������'�,K������bX�'�߻x�D�,K����"X�%��w��Ȗ%�bz}{�����t.�74�Ȗ%�b}�����Kİ�	�߼5<�bX�'s�gȖ%�b}�s�ND�,KuD���P?�~����D���5�ͷ���I���L�3����F�-f�ꧬV���Y�KnWt�pf뮎�s]���փ#u�����G�!�=s��+�gv�n8�c�\�\c��L�1!���u�v�L�,���ߜ�}`�l�5"�r�N;B
��u��mBC�ö赎����w^6wήm#�u	�1f�����
�
e]ZG$�]�����}��BIq��[O<"ݱwa�b�K��H�]P���ls���������3]ݛ&�ާ�,K������"X�%������'�,K��g��bX�'�߻x�D�,K��&��B��J���{��7����߻�O!�G"dK���"r%�bX����x�D�,K��f�"X�%��X̐�R6�J��j�n�!2!g��9ı,O��v�<�bX����ND�,K����'�,K��I��m���۷2awvD�Kı>�����%�bX>�{59ı,O��w8�D�,K�͑9ı,N���Βk7dܳnn��yı,{���bX�'�߻�O"X�%����Ȝ�bX�'����<�bX�'{۸�{x�*��u��9ƍ�Ae��ZY��ۧp�N�����q�3N��ujr%�bX�g{��yı,O��6D�Kı>�{���%�bX>��59ı,O>�p�݄��sww.�q<�bX�'�w�"r�^�M�b}���8�D�,K���S�,K��;��Ȗ%�bz}{����4Й���"r%�bX�w���Kİ}�xjr%�bX�g{��yı,Vf�+!2!2�0��T�t�*��\�'�,K?@�?~��Ȗ%�bw>��8�D�,K�͑9ı,O{�|�yı,N�lû�2�4���]�59ı,O��w8�D�,K�͑9ı,O��|�yı,{�U
�L��L�����"j��T̳�.'m[-��4���6��"��;8S�|��ѲMɛ��ۚfٗw8�D�,K�͑9ı,O{�|�yı,{�B�H�{��r	 �^���l��&��ɗwdA$O>��ND�K����Ȗ%�b_��w��KıY�t���L��_���QNB�\�'�,K����Ȗ%�b_��w��Kv
tT/AGD�L���,K����Ȗ%�`�>4�wssw$�$7ni�Ȗ%�b_���Ȗ%�b}�y�'"X�%��~�Ȗ%��Ud�~���Kı>�gp��n��ݻ����%�bX�}�l�Ȗ%�b}��É�Kı=��ND�,K����'�,K�������;�n]l盶띓����`v�s���]��ou��u�.E�P%Ǧl&�Ȝ�bX�'���O"X�%���xbr%�bX��~��<�bX�'�w8D�Kı=�}:_ͷvCw&ə�Ȗ%�b{;�����G"dK��oȖ%�bw���'"X�%��~�Ȗ%�bw;f��ݷ7&i�f昜�bX�%����<�bX�'�w8D�Kı>�{���%�bX����'"X�%��>��d���f�����Ȗ%��D����S�,K������yı,O���Ȗ%��7bw���8�D�,FB}�k�)�UN]1�:��Y	����~�Ȗ%�b}>�ND�,K��{�O"X�%��oxT�KǍ�?{߳~��S@V�u։x���X��Z "jG���mRaѤzΓR�'^utYБ�ۙ�q<�bX�'�����Kı>�����%�bX�����DȔ��[�ߕ��Bd&Bb�9Rk��j���&m�19ı,O���q<����,O�_�*r%�bX�����Ȗ%�b}>�ND�,K߾�-��I772nn���Ȗ%�b{��9ı,O��|8�D��XdL����19ı,N����'�,K����%�ݙ�J��73J��bX�'���O"X�%����19ı,O��w8�D�,K���Ȗ%�by��t��.��d�34�yı,O���Ȗ%�b}�����%�bX����ND�,K���O"X�%�H��d"��'�F"V&�F��	0��e
	�<�&,bB��c ��b0X�V}>�zK!�0'��7��p��!T����1�!�P� hP:C�"��1b_|=WD�0�����YNv�j�XS�{9L�냼{lIuyv$�59�]����n]˴H��S�sգ��M]�:C�$��R��(p5�ۑ�TU+�C��-U���3��������L�#pҤ�V�YSYh�tگQ�d6�v#sIѹ hW2��۶a�{g�Z.��Ԩö�g�`g�l�@I��jM��6���9g�c;a睼њ��⣛�@�q\0D	v3#*܂W�/iG�����(6u5[V�k$�+���`���1��G<u�K]b����m����Z��E��N^����,��.��v�n��L�dw����4��c^�lb���'�����k�Ru��F�t���D�/����;[/oeu�1���d�@s�n�m���)�N}5mum6D���pU�fю�����e���}�N���vN�^cm7.#c&�`4��&���3���?N��������F� J��r݅"p��\�r�j���k�i�Pxݡ/P�J�a���(�ƺ��=�瘰©FMT���m����6 �jڳk�Ma`k'6�쪭PK�-�kjۅxz�n�]����`T8��\�M�������d�nH-h�5�YA��ש������kfkg[�)9��m[8�����2�q�. ru:Xڠ2���̎p-���V�K+J�qB����lu\;{a�Z��9�ErR]uS�Cz�qմ>kd$㵷l 	:��^aۓ��z�'.�����BŌ�rEK�pR: ���J�"�oYF��ݹ�;nz1r��"�;v�jxv�M�+��7�����K�֑��Ҝ+��d��`n��\v��:ޒ���Ftmc�a�.��/��l�!`�����
�fj��C���պ٦29lj4�pFx�{-Fm-ƚ^X�c@D��%��sC�g�����}Z;��SI��t�t�:�Y{v�tm�[��-�tT�P~E��Ј'¡�(����3�J
<~DM���z(�rYvOp�l�㉎�kFzr7Ub��;&x����%��S!CV���]sk·�>�1����0cI�����&G�78o�Kz1�j��m�Ŏ0=�mNہ���xu�7l����5���x�Nۡ��gS̅��jMq��2�cR��=�A*��pE��iػ\�Zܤ<C�����>ﷷ�5�ȺKPW��m��\���6K����[�������<�׳U:�B��]�Zɺ��l��T�<�����mf�L�7����/�|2J#vl��1;ı,O����q<�bX�'���S�,K����Ȗ%�b}>�ND�,K�{e��:��ws��Kı=��
������,O�w��Ȗ%�bvw�ND�,K����'�?�ʙĿ�KK��n�m��,�wJ��bX�'߻�É��2&eL�g�ẜ��_�v�w���'��ș�2'r�ᘜ��S"fT����m��w.K�s4�{�L��S"Y�xn�"fTș�>߾�q=��D̩�>���ș�2��*�/wv+��8RB�p�QĪMuT�M5n2]���r&eL��S����'��ș�2�{���by2�D̩��߽8��S"fTȖ}��ș�2&eON�~�=t��!\��H�=��Lh�u���iܶ�܎��n�����Y�xn���Knq=��D�S"}��ɉș�2&eO{��q=��D̩�2}�l��Lʙ2�}�{�O}��3*dO��d����\ͳs7&'"fTș�=�|��{�? ��� ��	�"g*dL����S�3*dLʙ�����=��D̩�>��d��O�wbfT�gg��nl�k��7g�jdLʙ'sf�"fTș�>�����ڙ2�D�oy��3*dLʟw�vq=��D̩�>��/�:����G�������=��{��ڛ�߿o�jdLʙ�s&'"fTș�>�|��y�L�r�D��y�S�3*dK�;��_�;��ݛ����'��ș�2'�{�19�L��S����'��ș�2&O�͚���S"fTϻ���jdLʙ>ܲ�����'JU��\����Za-�6�y]i�t�Z��e;88����������=��S����'��ȗ*dK>�6jr&eL��S>����@��SbfTț5<�aY
e˅ʖ���P�ҙ�K��8��S"fTȖ}��ș�2&eL���x��S"fTȟf�nbr&eL��S����'��ș�2fS����!���or��{��?�����{�L��S"}����ș��@�z3-�@� q,@�,#*�*C�@HU]F 	��&yS����jdLʙϻ�u92�D̩��Op�ܖn�3v�n��jdL��("�9�<�똜��S"fT������jdLʙϻ�u92�D̩�}���jdLʙ����'N��U��{��;ݙS��O}��3*d:���ẜ��S"fTϾ�w��2&eL��nv�'"fTș�<��m'�Y����4܎������v|�nxH1��9����F:����ww�Z�wΘ[����w�����{��9,���ș�2&eL���x��S"fTȟe���Lʙ2�����O}��ܧ�����<}MqLg�����o�2&eL���x��O�R;v�D�_�3�3*dLʟ~�jdLʙϻ�u92�D̩�=��sI���wx��S"fTȟe���Lʙ2���ݼO}���E�6%���u92�D̩������2&eL������@28�+����)�w�ʞw�v�=��D̩�,��7S�3*dLʙ��wx��S"fP�?(�ȟ��ᘜ��S"fT�i���-�ɒ�wso�jdKĳ��u9ı,?�F9߻�x�ı,K�~�ND�,K��ݼO"X�%��?��\��٫,�`-�Y0�y�mn9��ؤ_:1���c�:�3
�b��Kı/����yı,O����Ȗ%�by�����Kı,�{���bX�'�}8[��乸I��s7x�D�,K�{���Kı<�����%�bX�w��ND�,K����'�?*�TȖ'��ܗ��w6�ͳs719ı,Oo�׉�Kı,�{���c�C"dK����<�bX�����aY	��	����IR�Ҩo.ɹ���Kı,�{���bX�%�ﻼO"X�%�ܽ�br%�bX�w{���%�bX�}ۅ��ݳ6��ۦf��r%�bX����<�bX�ʩ�~�O"X�%������<�bX�%��wS�,K����~���I�!؋�<x��[9q;�u��:Xk#sJ�v&�ANSUs��1�5h�(�]\������&ڷ��^��M���z��0�S�V,�w5Z{nZ�${+BK���q4�+K&sKe�ۋ%��������<��+����=����!GHY�ym�Qu��.����s��O5a�Ww[�U1Ѷ^��b��ͻ5��w��s���;]nR�mH&�@k�����iV��Z�vZ��ZݚK�Bٹ4-ݛw.\��<�bX�'�_����Kı<�����Kİo{���Kı/�}��yı,Os�izm�f�wrd�ss�,K����'��9"X7�f�"X�%�{�߷��Kı;���'"X�%����v͖��%����'�,K�����Ȗ%�b_��w��Kı;���'"X�%��w��O"X�%�هJwwf�7md�����Kı/�w���%�bX���s�,K�����'�,K� ����ND�,K��p����7	��3wx�D�,K�~�br%�bX��{���%�bX7�w59ı,O����<�bX�a�;2�񙻹p���V�VY�΍��0I���Y��ust��s����XpYawd���ND�,K��ݼO"X�%�g~��r%�bX�{���yı,N����Ȗ%�b}��t�&�ۚC7.ɻ���Kı,�{�����X �D�SD�K�����O"X�%�����br%�bX��{���%�bX�}ۅ���3w&�n�swS�,K�������Kı;���'"X�%��w��O"X�%�g~��r%�bX���>�aзK�e�6�<�bY�H����ND�,K�����yı,K;�wS�,K�������Kı>ϥ��ن�t�[����bX�'����<�bX�%����Ȗ%�b}�����%�bX���s�,K����8gI&f�t�ś[����>C]����\��q���8���M�e���.���x�D�,K�{���Kı>�~��yı,O�����A�o�6%�b}���׉�Kİ��n��0�]����Kı>�~��yı,O�����Kı<�y���%�bX7��59ı,O~�p�/t�sq�e��x�D�,K�w19ı,O{�vq<�c�+�AU01<ӑ2��ND�,K��ݼO"X�%���,�X]�73s�,K?*�"}����Ȗ%�`������bX�'�o{x�D�,K�~�br%�bX�}>�/�����e�d����%�bX7�w59ı,O����<�bX�'r����Kı=�y���%�oq�߿�9C��7"��t��p�[`j�mZt���a5�Gr	�%�ɗ�(6��y�wL��t��.njyı,N�~�O"X�%�ܿw19ı,O{�vq<�bX�%����Ȗ%�by��Yp��[sM��͜O"X�%�ܿw19ı,O{�vq<�bX�%����Ȗ%�b}�{���%�bX�}���6Ɇ�t�[����bX�'��;8�D�,K�����K¨C"dN�~�O"X�%��/f'"X�%��OCB�SS*])��.�!3�)!L����r%�bX����O"X�%�ܽ�br%�`~5,O�~���yı,�g�?n湄В���"X�%���wÉ�Kı>��s�,K���gȖ%�bY߻���bX�'}�r��%񹻷6nd�2n��7>6y�sl�e�sQ!�ȣ�b7Ln�:/��{���s6\�����'�,K������,K���gȖ%�bY��u9ı,O���O"X�%�ӷrY�7wl���nf�'"X�%��{��'�,Kĳ�wu9ı,O��|8�D�,K�~�br%�bX�}>�/��͙�n͓7gȖ%�bY��u9ı,O����<�c�@a�2'�}�0���L��Y�|\/�&Bd&B�����U�8�.Z�w��oq���>���<�bX�'r���Ȗ%�b{��É�Kı,�{���bX�'����;6R˹3KeͼO"X�%�ܽ�br%�bX�����yı,K;��"X�%�����'�,K���C�0�ʲ���g=ݖ��i�7Yp;��x��=Gn�t�S-�\1�5�Pݼ<3�����K��V���
�{Q�Y��4�ݰEv��Jvچ)܇��S��clk��/SX��%>^7B�f*-�q�:0sn{*qU�x&ť��!�]��+���o-	s� ��FP��պ���؇��7R74!���Y䭟n<�ո�+C����<��-/����O{������l��~ۢ�c�ض�'df0؝�s�\�ny
x;v�v�o�����=x��[����bX�'�����yı,K;��"X�%������=��,FB�}�0���L��]+S��URT�ۦ��Ӊ�Kı,���NC�(1ș��w����%�bX�������bX�'��|8�D�2�[�,�S�ȅ36��-|�W��=m���f���!6�18�F�NE���Ē��{zl��V��V�I'�]�@�~�G�$�c�#����hB�{�����v=͛W��/��=�����ɔm�����B.m�%[��i�0vD�ێK�f3�.�6��[T~����h|� =mށ���\�[y�8�̑�M�Z��f\31�i[�ll� �n��l�N��؆�L�I'�����=]�@;���ڴ˄�v���Rb�z��hz٠w;V��z����B�) ��SS4�=�VD%�]���zl[w4�c1x+���I���_�ܸ�U��YC{VZ��cf7�M^�wS��k���/�Y����K@;�b����n���!6��䘜#NE�r�^��n�u�4�j߳?�"��1D�"�MPT�M���j�3sj��
D"�"�,b�o�2b�a���BB��J�
�� �Ő��"�lb�@�CQuA��C",bs�2BBB2���'!`��� р~_X�
Jb1!>��! ���`G��!�dD���P#� �0'6MA)�!��> �9 �4(ѩl�꼐��5_D���	!�)JҘ��8�H�)GP~ /$��|p����<!# �\�����H	U@��'�T�.x���S0_E4��?y���uzq�Ź0X�Ĝ�iX|�7��V��=͛����?z����7I�rM��Z�B[=�?��޵`��`f� Ý�E��.4��|�ku�.i.S��������;sI�D��b�)�I8�W��=���76����r{���i���)1N=׮�u�4�h�6o���j|�LuJ�ۥT9�`���d��w$�I �^Y&���ۓ@�v������9 ��@�^nw��7�O��)���f��j�9�`c�ٰ>J3��/�k��3'u�^�ؚ�)H9�n����Ny���On��+Pg��Z�b�t��ö�_e�X�D�na�@��s@�mzs�h��@�8��&�xԃ�1���DD6nOs�5�t���W�QٙϙuUN���4�[���5�t�Vנz���9u�@�|��E���!8�+k�=z�h�ס��"{~��`c��|6�Re:����=�ZX�vlܭ,=ݛ��
" �b�TO�;�f~�fdܳr�1�D�Fq:u9ٛ��Θ�1��n�Vn^t1�7Jv�ҩۧ]��O/)[\t���Z�y1��m�,讌�л������
k�n�OɃ�lanx�����n����%��s��]�rm�mm:-�.�Z�@]]cZ���6���qhf;���}���F{n"�4�lu��S�ڲl�Tv�Vލ�t�dl�F���������w͡#5�Z'>�۬:�:�(�vz�c���/������Ծ:���4��K�������`��bǰ@f�55�T�5)�56nm���Pً���/�|h�k�=�DB,��c�8hW��:����f%W}��/�|hα��4��s�z^��1�vlܭ,>�����`f�rv�!7��Hh���:����[^�ץ4�I	r/��O�j&cm��#�۲�t���'v-�ݙ��lH���i�U���I�H��)�~Vנu�M�uz��'�"ŋ&F!6�~V׾�X�!�(�$�W��׻�`f�k�9p�.�$�L�ӏ@��s@�ֽ��+k�.,��T%�!^Vm��ۓc���b� :�\Yd� �3�=��+k�:���9u�@����L1��Es��#D���c\��BۚE�^11�t���E�0�Cģ��rLn$ۋ@��]��Z��)�{=cbd�J77q ㊐ܘ�q�rLR�Ԧ��Ppx�2'3@��^�׫K$�+��Bj�wM���j���-�H�l��z[)�~Vנu�s@��@�_!<�1$)��[�����*@;�1 �� ���{~[�3ؙ}�S����A,=��ݫ:ʃ�\뛉�nd��L����N�;;m��� �rl�� "ˊ�B��� ��������?+��m��:�v,�L1c�F�wwu 䊐rL@9"� ۚ���Dĕ�1��H�4���^��36�%%� P%�脅}�ج[�#:�ܪ�n�SU6�6Ձ�({�����V绳`~�$M��5U,�]dw6PYm<�w[X &�K�a^^]�N���d�1L��Xۙ��f�޷s@���@�빠~�W�$j6G��u �EH\�T�sW�ٝ:�+�1���1��V�wM��͵g�$�f��X�\X�m<Z�r�l�.���@z8� 6�=��D?OwM��b|��uT�mҩ&iX�5 ܊��� :H����ߪ�Tr Ub���:��Snͻl�7#k4WU��=��P��[�;F&�(���v�9�]��^!�v�(7�-���;r�&��k1ˬgu�k�껷lv��I��m����7F��\��ơ���!\�Wlд�XjW��<���T�z6�2\���CCǀ�6�6N*��S�bį=�{Xi�Fs�b�vo�.7ǻ�㫐�-{Xiw[��3\7-&��d_W����_��d�l�7v\ܻ��f�2�E1�k;ݙl�j�1�Z�&�^m��۪�x�Ƞ������4��z���������~���b_9Iő���z㘀�� ��@>�R���d�74L�SU6�6Հg�j΄�D$��u�Ϸ���0��:&�H�T-��@��� =q�@tqRު��$�y��;��h���^����4��cXX'"j7WM�������5��*շu%G;�k+���;<�M	�ɈY2F��p�?+���w,=�\�#���V=OW4ܴ�arM���'���9���pH	��OA�q��ݾ��:Ձ������jw$�������f�޷s@���@�빠Z���	�C�1�"�h�T���1��H����vmZ�ƚ�Oɚ���^���ݫ=�j��w�sM��j�\�%'��n\�S=g�Gf[Qɳp8��7k��=�.�����ʩ��5S�7ﾵ`�ڰ3ٶ�=͛�0��T��CT�T敀gI��*@u�1���\�[���R��2UVf��sfϢ%�yEj�*�O�����s�xrI=���4���O呑��&h�W�~��V��V(����Xx6��i�w�U��n =$T�w�n*@5z����c��r,R`����nշ9]v{WIζç�qt\��Ob7�۞��|��$����
��=��s@�z���s@�<���d�bk�=��j���"��}�6�zՁ�sf������y�"�4W��?[w4舆��t��֬x�c6�9
l�
�����S�}���Ͼ�l��V�IB��rP�(q�O���ӏ��R��^����HnL@>qR�I�^��=�1ci\�)#�cM��F&�˝���5r6�W0u�[��w;�Ϋ��m�v�f�]J����36Ձ�sf�����Q��?��5�Õ�EIS3*fj���9�I �1 ��K��U]�l���i�n�NPS����j�ǹ�`wu��9{��.,�.+�H1��J�a��S��}6wWŁ�3f�������ɐI��r8���/����$����'/�}�������@����**+��**+AQQ_�EEE�
����
���Ҋ�����@UA������**+������**+� ��������
������TTW��������������)����*��*,�4( ���0���  >� vV�            4   P ��T��@UR"P�RR�AJPB�PP$	��T)E ( )@  @�
�% �  P �� ��o��:R�X(M4,��� :��:Fv��i@AM(��(*�Ϸ��ɮ -{ͧZs�)� �Ku�,�j��V,���7)qo6S��ͥzݭ���  >�   ��6AK�m5;��ڔɧ{<�=n ���q�ҷ}å�n�Ŕ����X��-\ ��R�ip �t�O]+�]�u�����J�� {{O-�zy5ꜝ;��ۥo  ��   P  S �)�ն�gתy5��}�r����kp ���}V󺮧.������޻�z�. =7W�ۗ�  �  @�������=�������v�j�r�7�y��\ k���׹��{v�[���g��|�P       �}���ާ��n�9yu�o6�-pK)[�ﬧ�]7WNN�`Ӿ��=�^�nx  -v�Z��ν��� {ޔ��rj�-�on���׾����U�ԭ�sﻯW���p ��     6�e����w�.{sﲾO\�x�� �=���ז���{��zk��_c�r��Ҁ^�   t��(�3�)K 
f�4����M�S@�P{Jt �:R��A� if �14�� 4�6*@� E?ԛSe)J� hǪ�E F��`=��J{B� �T�BT�J�� ��h�II�▓,�����U�٫�W��P���2r�6NNZ�I �+���`ATW@�(*� �+�� �+� ���AS��1?�BA���� ���HD!1E�D��D�
H���I]#���M$n��B$X4����G���M�5��4��A�����EH@�1�!�0HXY)j�bƐ`�8��"����dK!@���@���5�m8a�(�K
$R�
����)H�W�Q��@B�HӆϾ�T��so!X�aF2S�G|�$5	p�80�����WI����j���6p���H�Hs�tƌ����T�	Ma�Ã
��o
����M��P�XS0��#E��q>X3|>)"h2];�ڐ����
�!���'J0�����@�
�$�h�0�t�t��|��B�ԆMԲh��-&���T5���H0�K��8�)�6Q�B��XI	kv��alс�B���!\&Eq��3�ʖڜ!%�LH�Q��! �ԡt�ђ�XQX�B��cB7N1#���0֎_|:�K��}���oI��A��`�,"&'A�H40�	P!)XfפJ�j�2-f�3q�Hf�96�d���H�!�H��`#P�	Q�!HR$@%KJ���P�K�l-������ԉH�M+
��R%"��0!]D�������X4�H�����AȒ)�X)$�X�c�*B���"F��hH�a
jA�	3NF0<�ApϾ+�6
^��/0��i�ox'�T�~������Z2d��T�Z��	¾�+y�YO��P&�i���.]�����7wu
�w�Z���s������4g��>����̉��Z�%YȢ�\�ö�{��
IzK���㿱�=�H��g���03j)$Q~�|T�ڲ���ɗX+��;w�Ѻ�"���o���k)��3=ۭپw��㵀�"0Ha����o��!L�d�ɰ�%Hpԡ�сMZGsImu5��]B�L��!@�P��*R*�� �D� E S�ZR"b�!��!B �F��5+�ؚ�kR(��,��R��K `� �)�;��(h"E�*A�!P��Y4+�b�W#��H-C�
�ʚ%��!t��5���Cr�cL��]1#�,�5�	�*�B��k$b�8������{)�٦<C�bWS8��H��ɷ��,�.�FO��#R����	�2����ԓс.�MF���"3BE��lbD�϶`JhLqٲK�s�|58m`�m�V'��%���M��71�"L������b1"iH!ts�.��F5��9
kg���.H�����u�,'g̹��l�5L�u���扚�>��K��s��0��F|q!N�e��h�ь(¡

ʗQɘ�Zf^2���f��c�fX��#R��O��Y��
$ZƺL#]��td��e��CB˪�t��.$�0�)�c.�%	R]@!)���Ѡ�P�ŅXSc
�.�#D�]s���lњHV�F�)���J끩�ә��B�SL(F�J��4�D"š�-{��8nJ��a���i!M9�9�aY9r��d��&�����r]f�"D��� Ã)�c��ϵ����|S�
� h��M&]���wS!s���4l`�o-a����s[�8||(�a��g�с.�f;x��A��� �H��DH��AGS �Aa�SI��ϙu�]lwt�e3C0����`�^l%4sF��{��3S풚&�6����@;x�
h�$.�D�HkF0��8�"��P2$v�BSFk�u=4CFgRk7��+�ʰ"*`�ǋ�j���m�ю������ͧ����l�b8R]�p۠�C��ԈA�GA׌.���A�(H`�R�Q��b�O|B�"M�ot�8�9�u�!H�m�8t4]�*0h�¡�dZ�0���SW��ٳ�Ol���ђl&����)��C�!
ka
B��t�l,�l�	7ϊ���2�Iu�Y5���rH|k7��7�p�����g�+h��y���]�}������ȌHU�bJ���,�;>�@�pdM�)�SAu��5�V{W���ąP��"�`�t�SGѦ�];N<h�SF���
�b@�40"@	���A�Rl4$�8��\�ri0^h���&�p#dX]�p�Ms�e֌�i�8ˬڄ.�aMF�ąt8
cA�WC�)F\�]f�:�^��
���C�Bh�(���F�bST��k^�c�ؓD4�.��/�
��&���(Ah�u��B��1��o�}w���>�&h�-�O�k���/Қ%	X�� @6�� �����.�ϳ;�9�ϵ]bCqhB�s��^��aHR$!W�$!X���t!��D)��';��u�8s.����
1��1ܜI�6q�E#�7�2}��,�^k��o�s�����r���ަs����*<`��##��o5u�Ca�2�3Z�SM�MZ	��L5���%Ia�.��Ĉ��~
�"��7��l!M2ɠ�M,b��E� ���44a�G��G�s��%3G�eeesYM��7oLމu�]2�ф(J���c�A���č4���o�81)����aR��
:p�E��7�	�D����uϳ�MCnk3����\�&�k��v2�8Hh��Ň�k!"@`D���tD0b�ns��z���Bf��)/	u�+(K�]�+�)�SD��t�F�##0(F	����4t��ٔ3�i!���k3&���V�����J	5���W0EB�3t�/6�>Ђ�2�%4BA�H�#BB� F�%�(B�	���.s#�:>����P����dHD�"C��h��8d)��4��4����1�}���?��A��
H�G���H帅s���!�2]|jS�7xF�Cy����#H�Y��aRa\�u4�)���љk$�n[�8;����@F$���.�s�r,��kIMc���(ħXSF!+�o�l��5Xh��;���]�U�D5w��[�:24	��i��t�b���@��,
SXl%�wu�cw�Iu����%�}�mֆ܆n����0��N�c
��{�:�Zd�i
T#���"P��cJX�XT"���
1!�c��4!\�$`T#M�7Ii��!!M<X��^�>��)��3P�UXY���>$�k7�00 Ɛ!�0�1w��6�4}�f��@%����	��&��pe42����	�0�T�!M1�C�p��@�!p�B��SH�X�u���%ta��ٶHWN;6la`׉)���{��цv�4�cs|n�zC`MJf�2GL��s�f��6�Û!N:N	T�9͑���n�	�� Q�Xd�K��n7Xva�N��X0����T��9�l���j̫+Y�>G�����QY~0�rp��M��6f����5��<�Q4�����qw��9�6��3��;7�8,�i��q��%=�Ն�h۳a�-�M�)����D��Gcs���n�%5!�i���]1�,��]Q�|�aX�C7i�O˜���|oe.�'C�i�w7�6�))�|4�H:�|��Qؐ����Y��F4$���D��0ټ�q�Ѧ%cd339�.�!s7�a��4�sn�H]a����6l�7驆�Ѹ�s.���(h̹�&�T�)sy���b�HÙ�ؐ���08|}
kp�͚��8a���03�db`Tцݰ*���c�J0��vn@������  �   ��o�      �          �m�     �Y���m6Nh`��rM��t�����v-�k�y��.Mv���O	��Drfk�#�3��nH��Vج���-e4�Z]6Y���E�Sg�/-�
�����"��&��$v� Ft�� E��2� �� UUUm�i��H�    H Ӏ:�7-h ��o0   �m�m6ۇ�����U@uT$mY�5m��������b�<��α�@:` :A�2V�oep�^����UV�U�[����H ˙���� ]�&��\��`�Z�X9V�8{]/Ե!u��h{Z��K��[xd-���`m�/[o˥�}���mְ �UWK� )ҁ\��5+�i2K��&m��NY�J���q#�������:��#�6�  [@Kh����\�����}���mp�l;�n�ݞV�U��vU����PuKuT�R��u�	]�m���/Z�8h m�����@  � �m:m�mm�zV��-�Yzۀ 6��m�v�q�Z�t_U��ks7:� 8 *Vyj�P�i^��� � 2-�[E[R�(�29G�Wiۮ7V�����p$'M�W�w�T�� �PPHN���vF�l�Q��m�-�plv� �4Y��q���DZ�X
��uSh
�.�N���i���e%���lm������h ���m�۾ �@ �Ӳ6��s�{l5��l[V����VʴAKU,��N�[AN@���H ���*�r�mTUUT���@U��k�+����J�*�U�A:�g�#nLcBki�髩V��m �K+�-A��m �V��y٪�R	s�M�g�����#\�6C�����m'��l�6Ͷ���<���F괓��k�@%�S��D�:��_�~�ຩc6��TŪU�HU�WZ�z	U��sH�����	9�[t�8iɬ�-�8�mP
�W!5.�\3���ڰ�{LY$������lm$�� �oE�nͶH,�UTݪ�M����^�nר ,l�g[l��U��*�r�īUr��Z �	fL��f�rK��m�h�(l��T�NdC$+]tdX�'T��4\zZ:@  �ɬ� Y�Ā�l@K� l� ���k7Tn)�m��  2Hm���h�j�lK 8b��dLfU��Mۤ�5� � �ݶ۶-���t� J��;l�J��Z��6݀��6�m�6ِ��'X�&���` 6� ��o���k�$�v�H�X��e\� �UUWU� ~�j�ZHm�`�y���۴�ؐ6���j͛`m'0�]U/!QР5*�][f��Y=j�8ޡm ��ke����m��'��$$ l�A��5�Ƴ\@[] lH<�`�$�mz릸�m�M�/Z@��@u�K���( h��� IQ��ۅV�&3��Smq��� 6�� �!�� �,����[[` T����m�[m�8	l��E$mr%׭��ݖ��ie�@�a���E8���28I�:#a�$i F�^Wi1��-�6��� �$l�g-� r@<6���}�N>���@-�� n�v�uGU�݀I��B@ pK$�� �v�*�Y-�,�.!�X*��'hC�*�V�U�#����jU�%�W�t;�������ѳ����l�q�8��e%@�v���ӀFy^��P����6ݚ�����"�$�	Ibt6�:2�Jl��z���,|���H�� ��JH^�n�i���l�^h��� ��%���6� ֜ ��u4�t�����n�P�� q�b�j�y&���&��h�H~��;g�f���WU_+��� [@m�����z�^�ie� ^�R� ���h�nխ��jP����ism�H��R���U�pI h��Y��`   n�4jʶ�,����зjD�Ulp[wI���l�l,Xh %��t�%�M��m��ll� �  K�$�  �im�F�  ��#� m���%Z����*�l�m���V�H �=;�u�Ue5R�*�m���g  n۳i6  ^�j� ְ 7m�/,���[��@����\k�lҶ-�kDd�!�e�l 6�m�9�8�������EjAT٪��j�-i�TXkym�M�lv���K�Kz�&�\ �M�!!Ė��Z�nm��`m&�%-��Ӷt��6� ��j�m'8'���@8�c^� e�����zT6kj��{=.�-�����1�iI+�:tm�8 ,g[m��j�v�F���Ĝ�  � �� ���H�[Kh�:A�y��^�IKm�,�I7lZ�i]a�
�xq� +U�����`���4�qn�jL�]6-�gK�zP��Ѧ�g��}�_Tn��zPh:��j�J�{����-e���ҭR��<�/P�	��ll�g���n��Anz�5�ڻMνoY"C�ԉ2YXN3�s�n�ɗ���f{g�m����1�8�2��Y��k
���;Wѫ4�������	�ggng66۝�s�m���p� UB�N�Y��T*�!��i6�����mv�ͼ��ې�m� �i2�)�=f�6Z<qٷ\����$� r۞87`�% �/��d� �v���db�$n�O`I&�6  �6���UUR���c�١��!�m���6_���H����h��� oT��rAm �K&ۧͺx ��H]r�Q ����ŲY�  ��M���ض�ZV�ې  m+�FT�V�VV��s78�>Ԁ�ktڛkn @� p�f��;��:�v����\x�I�h�[l4�⸴�ܐ3��;: q	9��d��'@kX� �`[m�CE  �|���Ț����v��l� ඥ���K�u�  q�,m�� ]+I�m�ۤ���qv� 9��巶ʭ�˳]�!���4����5T�%^��Sfۇ;cp��0�U*7j-�n��m p-�d��$�]ؼu�u�����#�ٺ�+g��jU�o^�g@?�ũ��~'��K���6��ֶ�  �����l � ��8,�ས��l� 	���&����md� �6�������$j��`�Y{smk8 کh[m�m�ݦ�:@R�Np��-�`�m�Cam  Bڴٶ��ݤ��� 9%���fZ-�� T����  *�m:���d`�U�6��$�ٹh m�魸[% ۶p�[P,m
�UG�ⅴ�H�H���l6�_Nԇ8-��� H l��$�ki�u�d�$	��    qm�  H[d %�-�m�m&�d� m�m6[!�V�Zl��j��   �����H�$�i���r@�[@�mm�m�-�m���6݋h	9  6��Ė��nm�I-�9tCt�6�K/m�n��m�    9���   $8��\�E�Kh �:tn  6� }�>� � 6�̒f�޹q���Nގܓm� -��  -��    6� 8��� �    ڶ�nݶ�rA�^�Kh��[s��g^6��޶�l pH	�p$�   I
�jr޳k�m�*e����֍!F���I��kY�m   �Z��E����n�޸!�� ¶ÁoP�5�ݶH � [@뮷a 8   $�[\e�\;v�-h�E���]�8�r݃�����`u�m%�����g�m�w�}�� I#�HHBtkd��K&��n��k��δ*A��d˼��se:��^�V� j��;m����ammC^���-�6�
鴚@��6����8 �UHMC���%^40Ni��sT�X�Ā�� �۶��m�&( �-�Ͱ��p�[ �����M�ڍMK�[R�+6]��8�\��v�\H�ۀUjڪګ��4��"���.��ۚ�N`��Pm*��v�$�N�MkA��m�/P�m�t��2bZ�`%YN�1��eh)jt]�`�9#viҾnj��Uڪ��@�[vͶ 	6�m�-�[+ ���L�Y9V�թV���T�eP#����h���ҰZ�@�i:M���İ�ڶ����h���~����+��HV��,@�K��
�/EJ��V�UVV8�H7k����e�99��0;��p岶;�7W{u�Oj�;���{܈�����E�O�m1C������D�W?qC�� !�U� s�&!����yC��|��=�A�_lt�\D;���Lu���G�������B& G����t��(���P��
�v���,��DX�vyA�#����E<��Dw�#�Wa���Q
���<��U��bU���� (���@�(*����\bM��� 'Ѐ�PC�|)_�{h�T
��,���1�� �Dv���@D8� )� 'H�!����@Qy��>|�ĝ$���)�C�
z��w��Pz�(��<-:")��uU{�7�I�2 lހ�(�E�&����Q�Wh�U*l���������Q?�Ex�y�u� Qb�P8�'us�2L�����-�hIm��M�.��5��J��6�.E��l��%bzZD���jm�w(�=:����]c<v[����*����p�qa� ��׶��7������1v9ݙ��n��6��{.�b�j��
���n@s��e()Y�õ/cd�Tq$�9v+���h��/�I�sB�ݻ-n��NYҁ�ڳ��npS�9��M���n���lF�2��N�E͞��{m��v;5�k�w��Ѧru�eL�U�t�۬�L���o.{�g�k��z^����W�x�x^�s��4�Ꝏ��v��#�ݻY4�<��&1v��GnƬ�mf�	�Gn�5�Y�!����[�s��	�F,X׶κygf���[��;�YV(Q�ێېv%�� �;&ɋl]ptd���F�<B���bhv5�gd�3lF �(֬K�ƈ6��ر$4�:tFl��1M[���,#�p9�U-ѐ)�Z0=j 4��Šob����n'r��(���0�.��4=���tN2,�󮍹uэ&��[g��qzH�q :,�q:!b0��r]j<]�\�I�条	
���'Z͝�K��y� =�۪�W���\[*L��;l�It8�����.�6wX6�#��m��T��Ԭ='l�\����Gl0vi;<�uX�X�e͏f6�t�D�l�vE�n�6��nBz�j �t�냖z��kHJ۔5��0�����ҝ��c�]ե �{'��&��'�J)�gJ����vs�Pn�J��R�5�y
��<��p�����V�m��Ѕ�l�ٲn�Y�P:�5��-�*�Z�l^��J��4�+ d0��κ�MN&���J	Yy[��V�[m��XEz�^v�pl�8,�C��<�j��L:�*��GZ��+<v]="�ڞs�2��[Gum+�f֗e�nƎR��̪�	l��\�bk[���kb�]��x|u�������ʇP ��)0���@�8 '���'���| I�|��qcm�C#�*�R7FV�M�c�l�k^q�U#n�>�����\�ܶ�z՞�vz�ݍ�u��3̀{#�v(��+
���8et�]��r�[��(����샆���&�.�rM�k��Wg]t�3���+�pm�k�nz�;��n�ę���BH7bGR�gq�N�ݦ\cY����5����x��G^�h��������&�o
]�]��&}�A㜜o��SP�j!��RdA�@��� ļ4TԤ�L���t� e^���A>��
����MD�,N�߹�w�{��7�����	Bb�]�b�7ı,Nw���? 	H"�uQ,Oz��Sq,K����ND�,K��{*n%�bX��w�kų2e�榲�5�ӑ,K��o�T�Kı>�}ͧ"X�%�~���7ı,Nw���Kı;�}���,�K�,&f7ı,O��siȖ%�b_��eMı,K���m9İ=5��l���%�b_zw���K�Y�j�iȖ%�b_��eMı,K���m9ı,N���q,K��{�m9ı,K���I�fk����HuOF�rh����r&^�����\�=�D�;ڱ��n0�cG���7����ND�,K���D�Kı;���ND�,K��{*n%�bX���:R_��&��6��bX�'{�l����J 2�T*h���jw�,K�}�m9ı,K�k�Sq,K��}�W��ϓ>L�=հ����Kk%r��%�b_��fӑ,KĿ{^ʛ�bX�';�p�r%�bX���ʬ>L�3�ϖ�q�j��[KIc��ˑ,KĿ{^ʛ��:���'����ӑ,K����7ı,K�{�ϗ��ϓ>L�s�i\e��R�mMı,K���m9ı,O�}���X�%�~�}�ND�,K��{��>L�3��u��U R���VG�
�/mS���s͵���<��O]��Y%CV�6XJ�~�p�3�ϓ>]��eMı,K���6��bX�%���T�Kı9�{�ӑ,K���}����Ѣ��Mf7ı,K�{��r%�bX����Sq,K��}�ND�,K��l����U5�?i�n�Z!�Z�mϗ��ϓ>LK�k�T�Kı9�{�ӑ,`*���p�M��^l���%�b^��ͧ"X�%�{�M{55��Ys0�]feMı,K�{�6��bX�'{}���X�%�~��ͧ"X�%�~���7ı,K��:R_��&��6��bX�'{}���X�%�~��ͧ"X�%�~���7ı,N}�p�r%�bX��T;��,�[���齞���f���{������Ox���nW��Tjr&k��k�[�w�{��ı/{�ٴ�Kı/�ײ��X�%�Ͻ�ND�,K���Sq,S>L�n��B��YiT��n|�&|�K��{*n�:���'����ӑ,K���kdMı,K��}�ND7���{���4&�ck���}��%�bs�{�ӑ,K��}��7ı,K���m9ı,K��쩸��3�ϖ�rI��멲�W,�>_���bX�ﵲ&�X�%�~�}�ND�,K���T�K�U�� -���:�@�?0�bg7ΛND�,K��s�k�ۓEԘ\�"n%�bX���ٴ�Kı/��eMı,K���m9ı,Ov�i���3�ϓ>O�f�P���j��H�����9+��j�5۲�Fa�([�.��Z!��9n|�&|��g��g���X�%����6��bX�'�}���X�%�~�}�ND�,K��$�KcLv�2Kk�a�gɟ&|�ww�ӑ,K��o�T�Kı/��iȖ%�b_w^ʛ�bX�%��Δ���f�I�s�"X�%���l���%�b_��fӑ,Kľ7ı,Nw���Kı/}�e���`�?�&|��g����r%�bX��ײ��X�%����6��bX�'�}���X�%��N��*�������~>L�3�ϓ�͵7ı,?1�߿|m>�bX�'�l���%�b_��fӑ,K��U��B"�.�.�`!P�	�E�!P�"�#A!H���$�,#��_|�F����;d����-	�.ѧl�ʕH�$a�q��b۳��V`�v��5g�����N#����ݝ�u����	mR\iSg��5�u��#Iٗn��2g*�eq5{F�к�����˵�cO�-::��å� WY�%9<q�oF/6�{lV&g���FDZ��x�N�`��RS�痚��T'�-��<ۅ���n��o��b���1�[V�kp��7���q�qvNz�m�ay� ���J���˵�T{�{�d�,Nw��ND�,K���Sq,KĿ}�fӑ,KĿ{^ʛ�gɟ&|�{�Mc���,%rʳ���1,K���Sp��r&D�/{�ٴ�Kı/���Sq,K�����"X�%�ӷ��\5��-�D�k0���%�b_��iȖ%�b_��eMı,K�{�6��bX�'{}���X�%�}��K�3!.j�I�336��bX�%���T�Kı9���iȖ%�bw��*n%�bX����s{��7��������@n*�a��}ı,N}�p�r%�bX���ʛ�bX�%���6��bX�%���T�Kı?(����R_��RMe�氯INk,�Q�Z��Ҽ�n���e�eͭ���N�	�3f�B�1��I-���%�b{��ʛ�bX�%���m9ı,K��쩸�%�bs���"X�%�}�H�-�t���\����3�ϓ>O���Ӑ���7�z�ϑ6�,{�,K���T�Kı9���m9ı,N��eMı,K����.d�j�&k3iȖ%�b_w^ʛ�bX�';�p�r%�bX���ʛ�bX�%���m9ı,O���M]73-��L533*n%�g��}�߾6��bX�'�~�ț�bX�%���m9ı,�=���X|��gɟ-�rI��l�e�e�fND�,K���D�Kİ��!w���O�X�%�{_���X�%����6��bX�'u�{VK�1�1]`z�st���n:�<����V��z�j�{��܃��,$�I�,����%�b_��fӑ,Kľ7ı,Nw���Kı=�kdMı,K����$��sW2L����r%�bX��ײ���#���b}�߸m9ı,O����7ı,K�{�߻�����oq��r�����Yj���%�bs���"X�%���["n%�ɨy8�yC�Ñ>�y���ND�,K���T�Kı/����c���[s�"X�%���["n%�bX���ٴ�Kı/��eMı,K���m9ı,K�zFEmE�;k���ɟ&|��|�w6��bX�%�u쩸�%�bs���"X�%���l���%�bs���Z3fy�=��t ��k]�:�b���UA:�
��]����̒��5������'�,KĿ���Sq,K��}�ND�,Kݾ�Sq,KĿw���~>L�3�ϗ;�hI�mm�
�m�7ı,Nw���?�#���b~�����X�%�{�~ͧ"X�%�w�k�a��K��&|���O;m����f�fa��Kı?z��Sq,KĿw�ͧ"X�%�}�{*n%�bX���iȖ%�b{��̓a-�kYm.�
��bY� ����{����bX�%��~ʛ�bX�';�p�r%�`f�*�� !a'>�¥�Oe�
��bX�%�{}!�����fkY��r%�bX��ײ��X�%����6��bX�'�}���X�%����kiȖ%�`�wh�\̧��}v_g2U	V�9�ln�bn8�;�\ێ,fr�ŋٲlZn-5ﷸ�,K���m9ı,Ov�eMı,K�w��ӑ,Kľ7ı,K�{f�B���k$��0�r%�bX���ʛ��#���b^�߳iȖ%�b_��쩸�%�bs�{���oq����~�?�b�Q�n<n%�bX����r%�bX��ײ��X�%�Ͻ�ND�,Kݾ�U�ɟ&|���tnT�v�n۟.D�,K���T�Kı9���iȖ%�b{��*n%�bX����~>L�3�ϗ;�+mm�
�m�帖%�bs�{�ӑ,K��z��S�,KĽ�fӑ,Kľ7ı,N���Tw�Y$��Ɍ����\j���ﯘj�l�:؂���C�t���S��8͑�lrW�g-�[����k�'+Pnnv�6r5bQ����{n�[n�<�vp�Y7*�v/`�#�U��t���68Z�s�M�.�X@^z��
6�mַe�{\s�7�+5ٍ"�v":�\��7���dv�ٹjS�{w6��!7Wl>2Q�!�wln6��~@�@��
\p��m3$ֵf^�Y�-���5��9�ƢN�;2���̅l�s<JIe��*��,�~^>L�3�ϗ��7ı,K���m9ı,K���Sq,K�����"X�%�����iX�$U������ϓ>L�>s�ͧ"X�%�}�{*n%�bX�����Kı=��7ı,K��z�	�5s$˙��ND�,K���T�Kı9���iȖ%�b{��*n%�bX����r%�bX�����R0t��K-��ɟ&|������"X�%���l���%�b_����~>o�7������	�/Õ�w�Tz��ə��6~ �͚�fb�;�m��
�rP�MGTnA���Y���ۺ�`�\�v�j�
皗$
���s��|�e �1 Ms� &�� 㱹S�ڊ;n o;�*����E�D�A�H�ȑP�@1�s���ة��똀�e�̻�����슐dT�7\�� ��rl��J;%�Kj�7���u�@��슐^L�32��9�wW���7\�Q��슐n�{�K��O6���Y]��j��^d���(�/�ݮYN}�3������a*u���%��������?sw��ŀ�v�w�Q�4:[Y]���ȩ{��9�H��A�9�@K.~E�r��ڰ�w s�ۇTP�R	@ D��H�"���$�Č�B+�Hd����מlM6�ɠ�P�`W_�M�D��������P�!	�
$:Aj�� ��	��d�A�a��h�e�DŅJڄR$3P��B�6�X�*U?|��c���N� ��ED�s�"�@B��"�
Fo@���Q��z ��X
���'=�f�=�{��mŲ��Ij-�S�|��@�ݑRW�z��������cv�J�#v� ����=�˝��/�{2t�z�hI�$��>�?�Iw���5]�mtv��^�9�y<:��gYs�g�H'�T����r��7i�U-����ŀ}w8P�y?�z �ޚr:#�fbd�t��-� ���3�6���;���n��|��뾪[Sc��r�`s؀;�b=w��T��3� ���QPTՖ��p<�;��;�b�>���&Vɒ�&I2߾��M f�����-E,����� ��ۦ s�ۀ��@��w�	h:�����ŷU�ݱ!9�:hQm㪜��1�U��^oc\;qQ�̺8^e &�� �su�@~��, ��6��[n�-Cn� 9��@�1ݑRl��rr_8g.�+�U`��O۾���}�X�w s�ۀs�f����$��[�~䊐o �7\��� �s���+�n�ڥ�`�ۦ s�ۀ�ݸ�n��|���͍�ޖ�%���B�Au:�36�t	���U��$��H����֜X�va����b�ުrs�{U��Es�\E�ԩ��� ��wn4�v�ɺ����+u��l��9朝��h$Ͷ\���'8=�'�~���t����a��gc�csq����A;�A2
t*���]M���Vq-�81���Y8!11�<��Ѳ��Ss;\g�c�;��o��z��֯#��r	HV�st[�Q�7/�����شmmsn	�* �K.�� �{[���ȩ�y)�EASVZ�Km�����7q`�ۦ s�ۀΌ6�cC��+�� ;�*@u�� �s[��:�m=U��h��`��X�wn o{� ���X��mŲ��NZ��@�b ��@wdT��"�r�/�?���b��\���P�twj��m�1j�v�mXy׫�+e��Ⳡ�؀�ȩ6EHu�@k��n8�,��Km�;��,IE�_6o7q`7�p{ݹ��f�zO1�U�jbf��@m�Ҡ��hԙ��d�M����7��X�GݪIX�K%�̤�� �� qR�9�E
Yj�� ��n�wq`��, ��ۀy$��HWP��gg�a�h�P.��9nD˵�cn��SˮU��Y`��lac-E$��{�ŀv8� Ms�b�}W�K�������e�̾et	��H71 H� &������[+m��RJ�yݹ$��}�� ��R*=h�]��� ���X;;5�Xݡ%*q٘�$sdT���Hk���d{vY+�GU�ۀo;��}��}��=���� 	�ep����+]�*.�DQ�q������6��6�kW=�+r�m,�4�U�E-��Հn�q`�1 8� &��7��s0� �s9�Ù��#s�bl��9� �9�E
9ae� ;�ۀM�R� ����S�FfXs�fQW|�@M�R� ���\_.[��p~Ӭ"z�J"W*�qR ��@9�	�*@��@�v$��]�F{ ��}m�;t�-��c��0�Nx�&NԠ=0Jv�n���sdT�q�Ho99�Xݡ%*q�n w{� �n��;��X����M�6���e��d�Rۈ	�*@8���s�\���ȥ��Z��w o{� ;�ہ��}�� ��{=�4�I,��̤��sdT�q�H���wq�߿� ��x�����S�����K��`W��q��:C7\,�ɳtfݮK�1�[U�sd�m��6��"=����9����η\��fy�\ϖ�5��Ij�d�zYk���@�j����^mwݦ�1�B'î;iٳ�Nu�]�/R��m�] +�]
La�N����p�	�v57lۭY�4C�NN^�u�VӒ��?=ӽ�X�l�
ӫCn�3�ڍ�r�Vy��c�G:�M�c.th]r����GM���#��� &ȩ ㊐nbll�����V�7-�7����w o{� ;�ۀt�#�����ʐ8� F� �� -��V��P��`7��\ �o���ŀw{��w�l��;BEhBˈ�16EHT�#sh��� �[������plu�BP�<���d��h�/�L����]2�+u��dT�q�H��@9��\�YU��Kkd�`��,��KR���`C���M(� � "��P<
)���x����*@J�[���WWArW,�� ��ۀ����/�������b�:�6h�QT�*Զ� �s\T�q�H��@m�C2��D"��ۀ~��,������� o;� �ת4=���tT�ӻT�e��t�G{p/#Q=h{�!9�ɖ:�%j�=��/�������9�{ o�7!�[�7-D�U����2ffwnl���T�����J�v���Z� 7�ۀ~��*&^e�;����6h�$���y����T��>w���w}� 9����~������)dR�Զ�y�T�7\�5�@wdT�w��_2�'�\�n5<����$��,��V8h�⹆��C/A)-�yb�vdr�h%q�j��=���@wdT�z��|�0�*�!�XKm��ݹ��w�ŀowذ����t�а��;QGm�vEH�*G��۞� �Ob ���Ǫ�߈;V�{���u�}0	�wٹ4��ƒ&�z(�G��w}��X��Ѹ�e�H�IV s�ۀz�糠k�� &��ݢE�+�fr�&1�;�;�;����x��ک�A�A:�����V4�VE����,t7i��B���o�����슐א�����@?L9^�앻��[�~��,�I���� ;��������6{��ΒХ�֭��^N��^M�2\�D��@^wb�5r>͎J��rW	e0<�ɾ�6hכ4�̥Aܙ�^o�P�68�%K���L(����y4.I^wyx͞(޼��$�
!$�î������B�X�X� L�X�F!�%H���P A�(B�D Fc*��P�Dt&ȵ=`6 GDh�B��%!�a�ta0!�0��!Hň��q4��¡�����B�0b�I
�`�L���eH$()�T`@�6+�����g�N��׺��TԮ���@������%�Ye4�	��H�VT ��$)�)@� Q�i,X�t0�h6�#%�%��A#��]R�#�H:���l	I ���#HH����RG�x��CN�c 2CI��a0�!	pĆ�D��ne��m_s���*�HpN�nڊP�}��L0�������mej�pN�#���-.�bVA�0"���&�FB&��6��U�`V�`BN�!��w2L��� ��I o(�q�Yn��frf�vX �V��Tu�ԩm���a\��x��<��9��ndV�s����2L`[F�n��b�/<kc�깚�n`tz���1M��#�IU[i!�������]X2�WQʙ_O2v�&�R���n�fֺ�]�Ҷl��*�u���\v[r�0���������L�T+9�qn�*�Dg����e�6й۶�y�(m�8셺>���m�.�״8u&������n��.Ϫ)�ۧ<e-W \G����񌦨.�k-�v0�ь�d����G<�ۘNvǐ��Q��Y�R�Ϝ�r�
�ԁukv2�0��	��&�ę�����Zv�;�	JD�h\Q���m����F��&q�3���Svݸ�����j����-NS��i����b�w.Ux�6�^$y���¸�j�|��n�q��n)�@ZU��C��򛷓m�t�f��4���p�^�)�c�J�ʽ72q�v��d�*�f�*N�vɝ��mWn���C�]��2����[�/Ln����H�i�s��v���=��I<e�s�Kt�n�%�/��[&N]V�b�q��2C��bl�-��r0�i���h�$�`8��ȑ��%qJ�25]��
��-�#�m�h�
EV�{]�[��-��k�s<��ݸ���BZx��ò���^`T:���[�U^�6jC�홌��VՌˍm ��y�;T��U�̉C۵fCr]Z�!�Iwi�6�iP����2LR��B�v� lŲ��:H��b�b9�:�Bz��g����e%��묿&O��VZ�ͅj����s��T�3JJ-��S#�^`�����CGA�m,Jb8"z���-�윪&g˪8��Q�ն���v�[pm!\��y�m�H1��}r��^�b�͢8�[���m=R�6�T[J�O�ruN; `7d�/ N�v
9�R�3%�-֞*k���[DS�� *�W������}�Nۚ�.�Q��*�9�X�s�� �9��%�Wӻ�Aj뗤U6��Ӡ�ݒ���nɧ���r�yA황u��Y�茗��9�<�:�Xۨ^�ъ����5gr�����EB��aqH3Q9��6񮚆-�Gnۚ��њ�8�7'N&���l�4 
b"��8�5!��Q.�#@v;��p�����ܹ �[vM����v�RQ�4���"㸚��i#��d-�=��M��cn8�q]��4㛯.{mqq;��tɘ����V�r[t��b�?s�
 ��'S7��6hf�8��b'>8^e ;� ��U]�s؀5�b���=�I��lr��F�IV v�f�>�ɣ�7$��ԨΞ({̒X�����K0=�M��s��,�;t����w}0�l�#��c�Xg3� =_k��@v縀;�\��4��N1�аQ8H����{>���t�6����7Aj�ӣVM\���ځ]f]ffW@�3�o\� ����.���IPЇp�S ��veB!�QC}TA� ��I��ٹ'{�l�?s�L�K�����zR��"n+�� �=�슐א@�b �#����Eeev[p��ŀo;��޼�d����f��9>���L���)��u�@�1ݑR�٨���%���%NFHRЁFY��Bw#<#���Xf������ؐZ�y� �svL@wdU꯫��ذ=���BJ�KQc�� �n��"��� �1z�����9W�]����)e�;�b�7��Xj�JA�r��pwu�б�!mj�V��{����5�Aڽ�V7����PЇq�mX�vP��n��ŀw���v>��Dݱ��%���{sJ�x���7`�M�sݸM�\B�jƔ�/�b�Ud�*�m�����7q`��,��ـޛU�eD���ݷ� ȩ��q lski�{[K>(�Xy�� ��v`7�p��ŀ��I6Q�ܖ��*����{�4��J�S/$&L����1c9P����'}�[�fc%U��X� 9�ۀs���� 9�ۀ�P����@Y-"���);x�ո�n8\�ˡ0n�"�3�'VGV�?��#M�[��Z�w����t�sv����\���d�7$-��Հ}�+�&��� �ޚ��µ�ˏg����;#%���޸�wn�m� �ͺ`O��Z���!�]s31 n��ِ@wfA�������²�H�D����0s�Z|��4�^M 2fL�	%�������7sH��(�p��D1�giX' �����sv�H��ӫ�0�l=��� �4dv�N-���h�js�9>{�j�����s�7����mm�����r;}м���lfɸ�#���^X8�+��ا����-�x��vx��S:�!c]8�"'�2;�;*n��h���EbY�����3j�:������H��*&�\�o{�&�$�Mf�ׇ.�̮�2�r� .+��Vۉ��۞��!L����r߄IM���`�2h޼�o�&��v����*�nKQ���v���/��}p�o����������-��VKQc�����ǐG��T�#������7Un�ik��y�۞0�� w��ɾ{}p?{�nU,���^$�/ה�\�s�|}�4��
6��m���]պ��s7��6n��n�����l��H9鴸6V����+v;v��]̮�G�b �sC�]��{���Ū��"E%����܉3kD�:P�����5̙tA����N��MH� v����6釛7����}ps�����"JPs?�kJ �ݚ ��&�y�3��(���F�𫭹-Dn� ;�ۀ�f 6<�느J����¸�3����������&�5�<�Ds��,u���AN�!&YO�iT��Z�,���pon�y���0��z`�蟠�uV�u[d� ���M���,_}���s�|���z�ʥ��+k��`���������a���s< ��rT�"�\h��7��� s��s{t����,��g�UU�D8˙���@ly� �b ����Θ�\[^0>f:���Α%��;\��d�C���*��UU�<]qp�m�1��\T�ɞ큾��O�8�����D"J`��L�l7����٠=�8W�K�Dv�C�KK˻�L��J �� ��&�L��rt�=~�0ݱ���Z���F����sf���Ҁ��8PJK�L��$�%7��0l؞���[��Z���Dvd�N �1���FO�[h��F��秙��T)(��t�=	�k��ūn�`X�p�Mѫ7"�P�o���~���N �1��x��_9���c�2[L��� 9���9��`��L�������Ū�� 8We����@ly{����}3�[������H���R+P�m�9��`��L��� ;����!4�Xϛ���s� �@�bc� �1S�v�m��׭����d�'#8�)��KN�Xwk�8"z�^D��@)�k���;����F۬q��$��43�a8�F����kn���遍�������^�᧓ͽ���Wa:za���B�8̠��7m�0�\���7MW��T��tQ����k��&(k�N�6Hi9whJ������USצ��K��/=
n����(K���5�p��ۣ�Ӛ��%�3g�ӻu�7���oE��'n�IFWb�]9i�Mݎ���b�Ԫ�Z�#w��������1� ȩ ��]�&^W)S��rY����7{t��~a���`~�L��a����n��ǐ@K�q =s��e�ʴ�H��W)�~��0{ݘ�wn�ۦ�Nͩ�[m��X�`�b z� y� =UUW�Y����-�6��ur��آ��n�]�+C8y�X�v��6��N]�Ag@��#� ȩ H� \]6*����m�7{��*�_% �EHl��69���WW%�}w̺�� �EHG1 ls8� n�H�߫��-E� n�n =s8� �EH&r��L̮a���\��f �bG ;A H�}���ߟ�[E,�R��r�q� ����p�d�6�7Y6��@��ÖP.]�Vfs��	T��y �������q��H���v����9�똀q�K�vl99����0�-�����yݸUW�I!D#>V�I����� @���HbA#"$XĈ0��NM�R�ð�5�Ҁ�
$� #RB�D�O:`HU6*%D�#XA4���1�s�����lbB.�f�o��i Č�I&��R�	Mid	�B�(:*��B��$�Z�(�	���`�j���C>M=ڎ!���V(DD4qS�a�Ew����h�J�jf�}��}J����fJ�Q-|���2�33�1 ㊐dT�;�ۀu=]6P��R+P�m�;���dT�s�1��W.�\cm�1��t�;��s0v�Ӻ�	�^��(Gt=�o�_��EZN�3��h	j����ݤ==�c��q�HG�r�g�Q�-C�U������y�ŀ~��0���mR�]��Ie���@MqR=��W�{���1 ���"��-u[d� �wq`��L ��e�ߧ��7���}٪9aT�Em|�̤c� � �bk� 5�Z��B����Ubd��������ͫk���ënk���-�Z�t`�l�fe � �bk� ȩ���Ka~$jI[	l����x�ǐ@9�@J���8^e�s��E��	� �{"� ���ˀ��}��cr����{�{����\ ��n��� 7{"�/�"BZ�\� ;��p$�������߽훒`<`H���1 *�M�J
�ݝ�O[�I5l2�;k���*�Xtf��6U��݋��!�q;�������yՀ�M�'X�M$�kvrz6 8�p���8�
�\�k�s���3�!Y2Z�v��6�2���u�L�7>����ug��z���H��&�d �7;��u��u�������f�iHF#�����v&SkR�z�2�Y��E.�g[���ĝ
��i����{����%���©Kd*q��BX�s�L�q�Ӳ�B�n��^��_y
��`,�m�Z��I,������L��ŀ��;���U�Z��n5�� �w1 =s�%d%��#���r���� ;�{p���{ۦ����Q T0du[(�w1 =s����{}�m/čI+m�]��wn��� ���`w�n���U���6���[%���-������v�n�a�Gk��.p\tf�OOĶ;X+�C����0�ۦ wz��yݸ ���u��ܭ%(��
u���0�!�������9�\yۦ n�M�VHKP� �� �b=w�3�?yRd��mR�d�������7}(�������}�;�b�Ue����s15�dT�6;��69���{OʍF�����M��
�[�_�n�,���d3�W.�X
��;i�Rb:��s��� lw1 ls?Wl<�x@ql�J���p��� �����bk� �� �m�2�˾r뜉wwx�����h��=!���$0�h�~ ��{�lܒ{޾��;�ߵ�nQ��h����0� 9�{p��n .q6��o�X�_0@=qR ��b �s^Al@��]ܰ,�i�(�+ ��sƞ��ld���<#��TcX��r��n��fQy�etc����@My߷����,��s��b����� �������*��l�~��gY\���Um��y�ŀw��X6w��p��\���;+,n�j��̙�3%��T��@e��c2fIs��ݱ�ŀ~�M�A��`��%�@� =��{����ʐdT�~�����a�5��\�u�c����:��v�����jШ��ݾ���v�q�9�ww��g@����dU����\~~^󔶌V+@� ��qV��4A��J�3��h�y5��������b`�#�`�{ s{��7�p�w n��rV�D��/�5&fN���4{�4]�*��O{�~X�<筶+knZYpc����H�*@� B�>U6�5��$�Z4K���2�&\�뮵�	,�z ����#����t���MXlra�GI&]�r�[h�m�a�n<����aV
��h2��q��;۳��y�������;\�g<�1�a�m͗���3��P외���*/�fl����;[�X�獞U����u��9�GL�iw
`��xCgj��Nw��X�6��Ϫu�"�n;�޻����ߨ��՗��+��������u���z�[�T[P���������S��t�7��~��R슐�9�c���W.Y��֦��nI߽��Q?�";z&�3���˼�Z̝�`F�H?(�����@�����@F�Xy�� ��鶴�Ԓ�ۖˁ��;�����J��fR�ԓ��lM�?/��VՊ�m�7��Xy�� 9��p�ݸ�&�B��R�9��g��c\�h؝�-��8�+gp�ѕ{sl��|���X�a%���~{�b�e�M {/'�����Ԩ�lt��M&�5�K�XnI=�����?'ʪ3˷ ���,��Ş��ޞs����-#�� �� ��qa����ŀ��;��"���9d����=�@G�*@�x�69��%�+*���U�w������� w��o{���|���"�AXJ8��b�� ��ֺ!r�cҖ���a��Y�a��b�����P�T4Z��۾w ����7��Xy�� ���6���Jۼ�e�n9�n*@=�R ���~z�\����V�� ��q`��*9&֦I��+f߾+j�h�sb��6�����K7j�;��X��y�<�y�$���* չ/2�萖��U����g�����,��ŀ�S��Ɲk0r�Z�� ڳ2ڞ|M��DF�綝1�X5y^�+�俽��?55�ZG+�_�������;��X�s�a�RTY��l�`��K�vG�*@�׈��\�g��mJW*�;��X�����`��,�Dݵ��YmX�﹚�@[��Pw��*L�)�.��s�{�Λ�r��k����ֲ�r&^h�ّ@~I��v�yx��T��w ?:֫+V�EdE�����t�N�>��u�/N�mXL�Ћ��I�:���6r���q���*@�x���v`���gV��Ib�X9�Ś��73^h=���yJ�3�j̍���Ӑ���*��}.��va��o۾ŀw��X7l�e��krZ�Y��L���/v(��T�yJ��$�~��s}`{�*,�YS��0�w�"�& 6�N �f�_R���,�H#A �B)! 0#�H�$�����H0`B�B!$I#`E$�#�X�T�g�hӤІC��h��-�2Vn.#`E#!�� � ��`$PڐO�AR)���PV@X$�A����	�4�"�Њ@�6�A�<�&i):���^� ��	�"-1`D`A!Si"R�1#$B$C�B(Q�H �C!]� �5�h-Gw��330������ h[m�:r��$z�,��&�QE������e��d��:D�6�&���K�V0I��#+�էU�*�ȴ��z �v�fAp��|9M� õۓ���&�ntɆva�J9�N!�습U�J��Nð��e����u9�]��N�ݤ��;��㙚8rn,�XYMf�jKr^�=���0�	��1n���f�C'f!m��u���u\�.�� 8��Ƌ`�س�Ʋ�c1v^�Zu�HWM�㎰Hr���vy3��Na��덈�� s�<Ψ�_.��D��SVC����1v�>�81b�MC��FNE���V��.6��vݙ�WX��(lVQCE�[W��7#�U*��<�݃8�I�jSn�₵h�;�0�6��e:]������eݕ%2z���.`�;"m9�d��{]�%6��I�ѷ+w;��b,�Z���)0�Ѥ�e�g��Z�V	��40�JȈ5�U�����Rƍ3l��tT��eRs�=q������{r�^�r�K�!nL�qU������j3b��M���Lb��ۉLݝ��Xa����Ej�/�����ϯ\��!���ɎǷCT�T����h;��v��F�zO9�"�z�̥����T��v�y�R��<qS���BJ�^�8a��NqK�bl�&�nKg*v��E�kmm(=��v��8��1���h�f�q�ƶ��4��=l�Ku��\Aהg�V�3����=i,rDӧ6M\]<p��VV${u�/�	v��Þ�M��.���DuU;,�I�Ѣ�)� m��EC��@�FN�n��gE��X5�X���t�FdVZ�ujV�����v�[��̖؋fy'UfW&�B�K�K:Eq��i�e�ӹ�^^W���g�'	�c,\��,�d��7P��nz������d�W������<��d�;'E��*��tXӤ��C �(9�/m�B�[xz�.Vkq�Dx~�ܠ�<(��tC�<Ui��A�6tU�G�t��o�w�G�b�
ZӚ���:��ִpsV�(p��6Yi�`i�0o>�rA/=�֬�I��x���<#!�[���Bǂ:�^:5ە�nG^S^��.r���*\e�lA��{[��،� ������avz1�u�WT�o^�d�qgq�z�0$��"$�Ob�d�`�J���3�n.������g��v#�<�]az���':�O;�)�٭�V�8�H��t�=	�[�V�t;��-o�w����N:ʬmK[��~w�ŀޙ4�ّ�ɗ�y���F���.��������#d����� 9��Y���6k���_�#�I[n�[�;~�\T�ݑR ������e���E�`{���wߖ��ذ.̚L�� ������D��Wy��ݑR ��{'\T��_}�]���WQZjB
/5�h�mlu�&�9ńs@�#:^�75�������o�(��9h;%\ ��?�q�v`��,��ŀsv��RZ��Y������9��)�Tk��M�X��, �wK�s�`o�TY�ʼ��q���*G���1 ��� ���S���R��ʰsw Mp����n*@n��3�^]6�jUl� 7���ٻ��n��wq`����J�%��,�rm����we�uDa�ݵ[u�b�NH�:Yz��ˑI[n�K�u��0�w�wq/�I%���{��<Ed��Eh"��7/U}Wf��T�<�@;nq ~80k�[M��ݫ ����y�L��Y �Rݨ�@6���{� ��q`��-v�5$rЭʨ52fe�������w���2���$�aKk��Hݥ���pzOv���T�&�b�D���3���cnX��%"NT�2��ͭ����6��r�Dt1*"��XԕGl�J���� �R ���1�$�wyfVrw�3)�"�5�nbw��?�_&����n��bjUl� 6�I�-��(�\�;w�P�ԨO�Ŷ��QȤ���\��ـo{������nM���Q�������}�<Ϛq
b%8��"bb���H� 	��v����U}������v��n�"�Ok]av膜�Ν�^�W������&o����w_gw��i�*�2����Hk� �8���X��=�"rЭʰy�.|�7%k��Q�g~��T�v��ɈYmmI��V�.����7��X}�|�� {��p�n�5%E��*��g\T��qR ��b}��9� �{�ʭ+mK[��`��� 7�Y4��"��^R���,ďO���U"���Mv�nȮ�i�p�r�͎9�q�!����׌�l�\\�t���X^��u�)C�/d��*�Y��c�c�����	�i�8;C��D]�k�
lj�r��.��;/7![�[9�	�=���c�r)�kg);<jcm�9�f6W�嵜����J����A�`�on�wK�ּ�Pa}�k�'��YJ�f��C��s9��MGE��-�v95�M�<sƤx����S�UΐJ�#jt�L��F���U���{|�p���=yK�K��7�/��P�y�a��!DH�^I� �^Mrffw6�iP��T�fMrd�;��xiDJqL)�����c��߾�#�0똀><8:�Q	�xRə����* ��^ �b7 	9��Pe_8rd%�%P]���$̟/6~s6��{��ڍ܅R��Ua����u��r�����޲g]��@C�A�@��T�y��f]������*�}_}_��2K�f�4�wL)S3/*c9��n*M�}�՘l�T�$r� _�&�.L�2Qzw�\�0�e�	̤��ʐn^ �b7 �n�7YA���m��}��|߷|� G=��T��qR��y���9$RQ��w ;���=�_$��}�~��b��u���Z��أn�[Y\Vy�f��xl���v�n�c!����ظ���j:����h����,��q`��ΦL��8y�@,N�9���13Aw�H�/�a�=x�#��n*�d˒dɢ�b ~�R���;�J�I������'~�s|U_�(� 5��߷�wq`ݲ2Mu7v�Gd��jd���/6h��T�yJ���3����XI��%uYd� ��q`ə�ۛ��s5�/ד@}�.��&�Lm�>�燔5��-�Y&��9�˖���B�=V�nN�t�Ԏ���~�T�#r� =s=U�}U�I�H����u�m�U�� ��]���s�4@d����J��/)V����2e�z�����1��U�-w =�\[���*@�x��f�r�y���213A��2O���=���.��rh�XlL����!ޖ����t<̧!�U�fR�5�&f}�ן�3w� ��q`�١eCN�Z+����gӞ4�M*�8���6m:�m�0�䍮 U��dD�r� ��]���p��Z�2f_8{wiP�0BْT<<��a��e� �� #qR�EH7k�33.L�d�A��D)�f"%�L���{�\��n^ nb �Ӻ�U�X�V�j���/�I>o��P�k� ]�M3&I�3~T�6cBT� ����L̪ ˼y�5�372L��n�O��ޥ@}����%,�˒K��%��o$��TvR���=r���zx|9n������uѸʮ2sy��=��x�f�t��g�QlNC��)����/B'N�.���Ճ�Lqm%Ύ�l�U�n�`�F��M��l��A�qS�M���3�@��װ��l9����ɞ�i��^Q�Yc9�����yN݆����W$�-���ʂ�vv�.���XY.��54gw�9�^Zl֤5r���"��ne��4	�ד���үv�{b��q:G��߫v�I�2J5]���]�*�̥̒f_8��4�/ש���V�Yn�������6s��, ��&�.�&���'p^����t�|̫9y���{ʐ�@���ŀ��ڂ��v� �wK�w�@e�R��d����*�fsee]���f��1 6� #qR�EX�� 7������a�ZE%�F�u���[p�a�{pO%gg&l�v�����w�NL�H�-�WU��x�_������666?~����A�����L؃� � � � �{߳b �`�`�`�~���T�0�]h�����b �`�`�`���߸lA�GJ�|� �U	�U(b�� �67��}3b �`�`�`�{�~͈<�����{��<����APA�A����I�\���W��b �`�`�`����f�A�������y�������A����߿p؃� � � � ��o�]~�:4K5����L؃� � � � �{߳b �`�`�`�����b �`�`�`���߸lA�ll?�U�����~����A�A�A�A�5=�_노Xf��$�flA�lll{߸lA�lllP�X����?A����{��͈<�������6 �666?�ww�����n����Y��3��ry���=���.�K=�@Ͳ��m���������af�a�� � � � ������A�����L؃� � � � �{߳b �`�`�`�����b �`�`�`�{ں/�$�5&�$��y���3b"*X � � �{߳b �`�`�`�����b �`�`�`���߸lA�lll{���5�W2�˙�5nd͈<�������6 �666?���6 �6 瀂 ~b���O6�]����iܭ�-%�d.��
@�L����$$GB0
�X!�H D�+�J����t��s1y��L�&SJ0�P+!Q�ivB֢"0�@*����+R��SL��A�kpf�Ł�B���Z��D6��H�� � �"�O��*E�UV���Ȫ �?����w��A�������͈<��|��_1|����XI���Ues3b �`�b�*���~��؃� � � � ������A�����L؃� � � � �{߳b �`�`�`�~���jL0�]h�����b �`�`�`���߸lA�lllP�QX"��߿�lA�6667���ٱ�A�A�A�A��~��A�A�A�A�d����ˤy�����T�f�����vҖ�3��Fy���Ů-Аvf������U��A�����L؃� � � � �{߳b �`�`�`�����j�� � � � ����y�����c�	f����ɛy�{�lA�lll{߸lA�lll~����<������~����A�A�A�jw���K�����Y�y���y�~��b �`�`�`�wߦlA�lllo��ٱ� �C�։�~��/3*Ù������H��1 6� ��8�<SB�߽��ܒ{���fP\f��R �!��15�*�̥@s$ɓދS����*B�����<��e۷����qu�ms:�y3nM��m���e��ꪺ�ҷiz����\y�ŀ~��X��.ݛ�Eal����_3\T��R �!��3?��l9������mr�V��ذl�#�U��=�9�H�&rQ��V62;Kj���/�I�w�. {w� �^R��O���-�66^�!ȅ.3$�]���d��~_��J�7���=��	$������;B�Qܲ;q��\Nkۚ�Ӭ2�Q���[s�<Ev����`N��s�u�y���s�����3�-'��&7c�V�)<s�2��[�7��]���T����;FE���ݺ;p��xy�Ie��\��Ӓ,q�6)��ƴ\��Hd�4�����d��Ky��m���|�v�R�;g�GUtc
"UXZ���,i�%_O��`\}qZ�<��7s���pGk����b�n6�V���Ћ��@�����?c��]��[m|�`~���6EHG/?v���� �ղ"O6��-X�w n�^h.�h��*ԙ���͂D�%���ePv�� e�M������b�;�c�UW]��Wew����'��<�6EHG/rm��X[$��+����,�%��_%������ ˼�֋�u)��y�����Y�[��i�ܶ&�N
�:������j!]e����v�y�� $r� F� &���D�L����SW2fa�$����K�'�L�U����}'���nI���l��w�p{�D�&Ԋ���p��h��*5�&d��ݥ@��4&s�6����p?�~����9�m* ̼y��̒I�36hz�B��uuw��fR�EHG/nby�ŀs��6��eqV�"�;<D�[kD	�ȗb�:��&��.}�s%Ъ��۵`�u� �{� �wq{����Þ��`�Y�퍪��H�x�s\T��R ���꯾�|�7�ް���J겹n�� &ȩϪ����p�+���:Ǩ�hY-�Wj�����?w���w5�2�&��&d�o7�@]�f6G{
6ƣ��V n�]���p�w�wq`�;����Ej��VG9�C�ix���Ny�b�q�5�]1�DpV�=}���w��&W�R*��]������"�#��	��8L����U� <L���U��$���ݥ@��4wy5�333�/Z�P�5�:w��̪ۻJ�3/h�ə's36h��X��[�Xܴv� �O��f���ٹ<܎ ��Ax��U�!���tܓ���^��jh˗.d�1/4뼚�2M����f�* �~�7r���mv�DKe�0�sP��Q7X;7nس�i����Y)�yF�͉�^T�13@g�)P^e* ̳'�3&nL̽ f�M b��8L��<2�/3H� 	1 ks��J��W�Hn���E �P{O\ �;(�;� ��n,��vƘDڒ�Yxf ��n*@vH��꪿s�z`��I�P�X��-�7��Xd���'nb}TW��o%���Lnm�Npk��!�D�<�5��mc�M�����p��Hݎ9�u�q��muC�xۛ��BHR��K����C�vpv�-��ۛ��l&ܽp;h�2I�6_i����Sv�n �/&��	 �^ͻ6��Q��͙���'m�s��*���Q˴e��-A��J��n�4�9�q�r(M��м�;K���ً��ӵ�gӧVwT�k����(r�g���e+*�q�Hsvĥ���,����hv��p��ŀk����n�����T��P���wy��$r� 6� &���"��K�������u�m�vWpw}p��*9$��ۻJ�7s^h�̕/$D�DKʘ���L����Gf��}ܩ�$8�skd���_̾e�R�EH�!� ۘ�{"����{ؚ~�P�n�6�S�l'a�<kh{q'@%si����F�yn������j>뉂A�O����1��� �����K ����&p��6��jJ6YI����s��ȨtE_��O���X}�b�8�t��s��P�����b슐�*Gﾻw�x� �l������2���A�̗3&f���*����ɠ�$����{�C]L���۵`{�L�$�\�I(�ޟ��J��3)P����fp�=�K>8�(��*W\�cɚݻ&�w����AIp�!2����-g���{dT��RnHq �$ʒ�Il����[�w������6s��,���0��� ��t#����n]e�7$�����>����:���T��	����2K��$�e~:�&��Υ@s���T�6��imX��{�& zOb슐dT�ڳKs�×n�$w&$� ˼�RI2�2[��\���`{�L����IH�rU[��v��۫�y)C��خ֎�q��
ϰ����KJ�PX����p�w���@y��fd�� �͚ ^Ր�Dk�z/3(fRl��q� ����Y���/�l=�~u2���ݫ ��ؠ�ɣ�ffw�ݥ@m�Ҡ/f͒��]u�h�`��p�w�̥A�&^fdɵ2M1;[�O�n�Il����[�w�����,�{� 7�ۀ~��=TMD�alv�vBէ��8����p�ǧh���ױP֝7ݺd�#������X�wǽـ������7��,�G���Zm����2��������� ȩ6EY��:���R7�RQ��0۾�\��dT��nq ���QyA0�%:&h93'�n����T��"��&����[Ry���D�`dT��nq F� ȩ ��_U#H� ��c	ZR����-$ A�V
A"�# }��������)�k�x]��%7��>,"Cb%V���aeF�	�E���j(�����T,��
%ӾQ8�*V!����T5y�����333 mm��m��6o3�Ӽm����f��\p�t��v$��:ۢ�]&�eR��7Q��E֯9��4,�d���@N(]I���m�n��S1�mm{#��4I{qM�c9�������vEYz�ᰯ��i�������حs��mi8����:ӵ�2>�%��78�i�����vw9�V�\��a_a�YN�kp#c��n�qT�t�Mm�Rk����ܙܣ�7J3�-�1��2�.y�d�Z�ը�&�=(s;���b.3�����q`1��=b�k�v��������E�s�[]��q����GA�7l��I�������[s�sMg,�mm����l)�ݪ��imۋ6M	�A�s����SkX�-����4��uϫ	�ak;�ɮQ���F��NE�@�t�ͥ]��Nvz��{a��v5�w��׉���9��C�[�SlЂQ��4Ơ�s����*�1])*�RN�B������g����Vݘ03�{
�r�G*c�\윺g9G�n�x�'Z9,���p%Ȫ�v�K�v�C�e�\a :�uۍ�;��͇nm�q�ۼ7]=�����j^�̫(�W����!2mld�m�(I�����U;���z�2��w4g��:5����-c���\��g�֞����\q�2�N�IP��clD��͞B3�k�z�4�3Y{vxe�R�n¯m�iG[];[Xӎ{sG"�.DׅwR�tP�Ilh��uʸ�����s*�	�<�Թ�[n�e��@�ۓ���rYT�iuڇ(���e�Ǌ7:�+.���i���V�=HH(�s�W5 ��V55J�ZRZ�V퍵[�*r.\��,n���I�k�(؛A���ʸ�l�+8[�nTUm�P����/Ѳ�&D�%m��9������ۖ�v��0�TU�e�k�ە��r��B�v;c�J&Ct��A Ơ�F�v�����d�.f[ae�%Į�d�3K��͢8�6�AE8E@
��Q�E8�q)���ou!\tݹf�Jbsi%�nM'7��F��5�a���xn"�̦i7:�<�\���:I��煍nu���B20�N��nʈ�#�5��
ɑd��PeJ�R*�\��ܚ�Πg׎ɸ��vn�x;5���e�.�ד[�d�f,[>���y� ���U�j]<K18�x���h�Y��i��[g��\s��[Ϝ�rN�z#��Q~x������c���yW��)�˞#=c`h.v����;���]q�v��`ÅD��U��P��~�����v���.ne���T�ts������fG��� ��@=�Rl��q�/}v{���뤖�+�����ŀo7q`{ݘ���������,���9>��ʀ��ؠ��h%��IF_�ŀ{Q7Щ�Zm���mX�b��΁������!~��vM�l��x�"�UnGH^p�]���l�F^�[�wv�;}��y�����zh�e*뼥̒f���sb����x�u�ʚ�[�w��������ə�U�� e�M }w�\ɒwέ�)<�hv��`��, �wn w�ۀo;��w��J�U�KQ̤5�@��	�*A�������V���r����ѷ-���p��*�̥@�ɠ9&fI>�񿣭��]H)�	�����ܜ���m�<��-�N�צus����+s\�eŁ�{�*�̥@����/��٠5�cr�adr��r��������ɠ2�)W3�v���C�ø��%ə�@{�@w�E4��X̒L�Y�b�;��X�]{BH�ڒ�[44�m*�̥A����4�g���`��49n����?n�, �n� �{� �v�[,r[a�]eƋ��'�Wgv����)P6�g�(p�e6�����Nci��P��{�ŀ�1 6� #qR ���C*̬��p��@d���$����d��ٰ�h�lm�A�m���p��*5�d̝����o6h˜��L�G+���� ����yݸN����7���7$����WY����]g2�/�H� 	�b �s\U�onƪ�u��CDu�U�O�2k�#k���#[tgyul�ୠ�:��	j+����_2���@\� ��@MqR�İ3�M��|FԔj�n ~�v��$�m�Ҡ=���=y5�ə$�jsu�*Ab���-�=��,��qa�̒N��l�^l���D�;�C��&U�&L��ߕ m�� _�&��|������؜�S"��j �X6L@z��'��zO*@vH�U�r��s��n֡ ��:�P�������"`���]t�Ŭ��D�:�^vNxM���d���n0����V\�:�l�**nwY�tnP����N�k�f�6̯�L��' �	@���m׃��ͱћ�]�8g(m���]v�2@�(�*�7n{'<�0Q�p���н��Ę0�x�v]�k���q�ѻz�㇗3��!�ڱ�O�Yb��J8(�*ǙM��ݡ��v�ʶaݻ�\v�]q�\�n���p���*mYam���ۖ�n�����#qR��Hl��q�˻��a��9��s/���T��qR �& ���M�}�W���;K\� ��X6L@���T�ݣ�s*�`]�|�33) M�nb7 ;���3�G��DFӕ�m� ;�� &���"�5�@��y�-z�'d7�9���۟o,�Գgi:d)ά,�%�k�֩#�T:��e`9n���@vH� Msnb ��\�_%�R\�$��7$���n
?mC�D9��}]�L������#�_!��X�v� �n� �;� ��q`��� ��]�Kcn��ݷ ���T��qR �& �˻�u�%���-�7��X��������p�Gn�!Q�Z��m�l;i9�l�'��mMù�-���T#e��v��V�{��y�p���{�ŀs�E�jN����mX6L@\�n*@v8� n�s�e��4�m��0�����ņ(��T�y�����r����,�o����4In�n��?owǽـ�v���N!�Z؀���qRn9��� ȩ4��E��q��s�8kdG�K��8���%��G\W �v���N�����zE��+���9� ��@=�R��H&r�L���ܴ$�� ���Φ�n�@���,��w�6wgv�ܮ�d��Q�p?yR���s��� �/9̲Gdqʭr��;��=�� �;�r|���� �M ���͛�{�E�jN���ݶ��{� 9���;��X�����݌$��b����9�Ky�1�=By����v�h�
��A{<�:h�Kk�6��m��0�����ŀ~��,�{� ���֪,�Z��s1 �EH� 6�@nb�W��s�N�b`�	j�9��X�f ~�v���, ��'4�QX䶎�H��u�@=�R}��W�}�`��7<Eem�k$�� ����:�T��qRm�����XL9Z�B�扦z�s����۶h܂\������1N̸�:�d�C�V��k�N;F�ޕ����ɧ�2�M�dz�ms�E��r��k��\r�P�x\1�呜W5J��^$�x��z�'��;�����ff8$u�A�Ҹ���4f���q��XBiv���K"��5R��\鶇WG����:���ˣ�;F�ֳ$,�Qh��#to�̲�5ur�r��g�(usJ�-g�u�;V�c����<��R�7%�5-,��iGm���b�>��*�w����$�/@��@k����#�8�R�V����>�f s�ۀ~��,w���M�[m���`{�� ��&�L�d�3&J"���{��� 9�u�]����ـ�wr*@wdT��nq*��]e�b&h�2���˙3+��/������ۀsMՑ:��B��N+�5�&�y����uv�dU5 �q�Y�V\\��p������;��>�f s�ۀ~��, �z�qm�rZ�;��^���J�#Tt`�V���J�.sf��ͥ@}����$̓��y��F++m�Y$�`�}p��Ň��%�o��b�:�}0l{�ƥ��D�ʙfh5s2M��T��*�����p�n��#�8�R�V���s�똀�RnK����݃T�zx�Eۧ����Zy�� ����)����5����{��v��*�32��=��� :�T��ȩ s��-q�4ԅb-� 9���?wr���)P{���dɝ�Nf>����O2�L���T�̥D�fL�ٍNB=�w70u�kN�I=��9��$K�5o�M(8�h�P�2h4!�"�)t��D��B��ʐ�+4��` ������!
�
�!u(B��LMcRV�1!a-jjHA������
��,h£��(D�@��ĉ��FkD"����tMk��	�t��kq���P]A��-���	7H�� &�IH�c5� ��ml�P�ԣ����6ehX0����h�!!WѪ��Z-#V@����q*A#"HA!\ ���R��phK��,@��Hh��ś B����`�ac&�UMkN�1�H���*�k��!é���H��^��E] ���8 ������3&e?2�I3���P�y5���<�L`�D�`ｋ ��v`9ܚfL���ߕ ^b��
a�&Q�Rm���� :�T��ȩ�����[�o�P��6J㍦�U%�8�g���7<��&��Ï��w��륤ՙ�"dzzļ�L�1���>��T�̥��&�}� k���������;J��h�\��� 6ۜ@�b޹Y	m��r�\� ���X{�%�2Iܻ͚ٻJ�'sw;1(x�t��kvڰ?%��$�7}0��\�wqP{T�d��Օ��@�M��!<:uK����z�hI�L���/���Ҡ8�ݘ7]B�U��b�ʇ�k�D�<#��l�(�5�'l��5���t�7�ZH��"�eM9-�?ww����>�f s�ۀs�����X�KV�{���&fnL��4A���@��@}y���|��H��Y�KQ�`{�� ��@uȩݑRIf_!�Ùǘ��""&(9&d̝��f��nҠ>�n,��ـu�ݮ6ZWe��Gm�:�T��ȩ��� �sʯ����H	�޵m���HkR�l�ԞrWem�&6�&r.���:�Z7��/���a{7:���C�'�.�j��n6��]�#���Rs�;v���lQ]��.�:_l��́�M�]u�qW!��g=8�mz̕�y;k��\n�+7M9ڶݸص��nmj�2�	��C�m� s��N��Б�]�&���g�GJ[;@d��ݱҏ[�)�ǽ�w�t��9�p7t[@vNeܻ]��Oi�ơ��z���<U�lWNfZUD�J�=���=�E {ד�̙&�Û�b�=�E��V���ݶ����@�b�EH슐캜̳��MHV"�0����wqa���/�|ｋ ����53�z�EQ++&b�EH슐m� �1 C_Z�mL`�D�`��� ���7}? w��~��,�wr��XI$f��Wg.l���2�`G%�̚6JE7kF���jۊ')Y�KQj�8�ݘ�wn������ŀn�+&�Y[v[��� ��&�2I�7�&L�Rj��~��o��X{� �ǻl�We��K��\���#�_U}v�Oq 7=p�vj�Yd�I��*���%��w���_���u�@uȩ#�&f򲋠�˼��@m�8�7\�\����� ���jAS��Emi������q�]gk[�V��f[���N.�/b��wC���jB�����\�wq`�������^�����,�eM93r*^����5�ʐ��똿&��^��1��!Հs��,���6�����nb�EH�\��VUc��Aڰ?��>��L ��������ŀn�*�H���md�^ �1�"�vEH��������?��u����v#DS��+�#u��uӇ3sm�9)�]	�u�]7`�CV�b��y��?~��ݑRm���� :�٪9e�Y$r�\� ���Y��Hk����>��Te�DK�����32�m� �1�����*@k��`9�9��9R���|��䓽�l���TיJ���,$�30
�� $!��#� �Z�k��.��νu�	�U��3r*@uȩ��� ��`�N��cv����+\�0]����n�=�J����mó�
��,��k�l9�(�e ;$T��nq ksr*��HɥeV9-DnՀq��0[���R�EH	%�S�\�̻/�(�x��]��^e*533'f�*�w� ��݄l�Wd��+������"��s�[��v�%]�9���#�Z�X����8�ݘ��n�}훒i_�Q%�~���dݿ���K�*H��n�������C�W4�=r\a�zس��v���J��C�l�˘-N���wV��%=6n���@+��U轍ge�<��lV�j�U�h����<�N�{u��<�-��3�4Y����<��nV"�]���n���f�vw��cc(/O2�qd4ifC�3�g���N6��j�W\�;r��4��c/o���y��\���,�Z��Y��(F��7h�v�)�1��N�-�F�j��*P�&	w��X?vE��y�?���{�o�� ;�4�VF�#�E��[���ٳ�T���*@m�8��vi�)�)*�r��wq`��� ��v`;ݸ�dDژ���fR�EH���1�"��댚FUc��F�X{� 9��@uȩ�"�*��J�Z\�\�fvu��ԩ��>{���@��q�.����w4d���YTV��-E�Y��������?ww����9��a%U�+�̾f :�T�s�����⊐m� s�s��^����,�9U�U�s���s�[���R�s(/2���w��H���1�"�����sZsXVF�#�E�`���R�EH�����a=͊�=9��hv����H��%d�,��l�'L�i�N�Xƪl�ӋF��v�5�6{ʐr*@m�9���� ��dD�����j�?w�P?>s� 7�ۀ~��, ���M�U�KQ�a'׽��$�}�f��j*E�0@1�L��2UW�T��J��ɇ|�Q$�]�3(�_3�u�@uȩݑR/���}���}�(�*��]VY-@uȩݑRm���� #���m>��m�������F1���{n
���ݨ��b�p��A��ʣu�슐m� �1�"��9yS%U����V����s�p��ŀ~��,��&��Ƥ#�-�@�b�EH슐m� %���E���� ���X�n���^��ܟ��HE�,b�1b	E.��~��'���O¤ܱ���7q`}�� �;� ���XV�����&:��T���C���>���{8���H�=m1�r���;"N2���Հq��0����wq`��� ���T�u�-E�Y�\�\���*@m�8�s��W.�evJ��n������ŀq��0�������,�K$�Uk�`����� �& :�T���`�i��e����ـ�ۀ~����=��f�C����X�tO��Jv½���o��|�H�Sqө��-�gKΨ�E�4F0`�Q,�1��YXZ�
H�P�"KH��JA�)*@�����D��J��8#�KF��FtJJ@��R����*y�J�	QdCB��_*�`�d`I�!X1"���bD"��!"�"B	��B�`��-%e
R��0
B���~~$  mm�U:�{���mq9�n��z:k7^t���ҝ��$��EUV]�ے�V*:HA����6�M�����7�J��M�1>�=paŨq�p�A���g�nՎ�v�N���:��q:��٪�'3�ʻp�s�R쫘��ԍ�b��o]`�j"o,{g�ٻu��S���m�p!/�����7a䙤5
k:�Z�l�;d���C�vh͇]u����N�\[=7<��:���8EYc�U�Q�qΫV($B�;�Hl��^r�]�m��a�-ɮ,����5�p[��Z�;Ta+��-a^�Z���:Gr�q���l�O�k8���A�0�켥9Q�ε]���pgjq�kciɩ3��V��N�\5n�[$�u!N�� ��M��kWnRt�ɞuu�qvaK~�ﾝ��ҭ+�`"��.��3����~�R\�X5r��� �<���G���璳�M˃���9 �����n�Ѷ79�0s�]:�z�S�v�i 9��Ֆ�;[7=��Cm���$�ɻ2�EĪ���+�����P:�G�GTp)@k�Kʎz��'(Y:����q�"aV3��c�"�2��Z�:;>�u��ݤ9�e#!؇r��#h3�eď�L��H�÷i6Yq1���;
�#�O��>�:��ѓkD���+/���<"}����ϛ]v^��QU�Bā����tNX,��ŒB�T F�%��Om�}?<|��ݒt��Ѝ��'�M��e�lq��j��Tˍ��cal`��n��,��5D�vl�J�m��nV�@� �cvq���'\���vSs�·!YyceU'����p�s"����E�]ST��$KW knwm!(�@¸ZH�X�1qr���G[��W��!�5��l�gi�BуDͰ[*)��ÙA!�>��u��v�ajܴ�<J�����q�6��m��gnuX6��]�)M��D3��^��󇋧�u!�u��ڹ�f��ѣ3$�� � C���x�@�� �*E@�#���0�E	������?G�T�9�4�ȳ"�:�݇l�.�nr�'�]�lG��,vtujR!e�N�źuz�����Du]��U}��r�X�Ж�Ӷ���Nkdݎ.3��.Z�ga�d��y���G/ljͶ�]�\������3���K�o;O)nx�v噰�M�ҵI�gBM�p��ρ�;-�R��*^�NćH�"�w�iY����7�$�S??ߣ	*n:9`���k�Ŷ�5�k��8�-m��e��@����/���V��[n
B'S�� ���\�wr��� =�c3��e��ʺ/���*@F� �L@K�8���%c�t����0�Dʠ;w�P{��92d���v(f�* ����2V9-D� ��v`|���wq`}�O��~X����R�ܱ9f �\����l��]}<�����ߟ�P��\�rk��u�s���V��nӵ�I$�5�\��T�d���8�bX���3�� ;T��nq �\�����,�K$�Uk�`���<���T���+�I3.I����"���ؠ>��X;�s*��ƘX�*�8�ݘ�s�� ;T��6_C�Ƥ��vف��_=��L��b�?ow����5�;���TX�PY�uȩ���s�z�	)r�����}r=a1U\h�Mkq'n\V�l
��Z]��������+�;��Ӧ;�'c��m� ���UWl6{ʐ�q��U�KQj��v�|����ŀ~��,�l��c~�JW[�!��nI��~��{�ٹ�x
�QBI62Z�L�C2�I��yڥ@�٠:��ln���Z��$�}���{}� ;�ۀu�0z�P�Id�x�2�*��/)Pe̓&e�S���L��ŀk�Ӛ�O�m�[��<�a��^��m��2)��u4�"
�B�VZ��������,v0�+�U�{�\��ـs{����ŀq��	�$���s1 �\��v?O*@o�� 6ۜ@k:wk�Ш�;PY�~��,��iQə3��f��y�@y�2%Cİ<L�2�92d�ۛ�-�6(�y5&���ʉ�w��$�޳Z���V9-D�_f�Cm�|�����l�{�����~��{�m��	Fr�mlm�eӷ]l3�	�3�F����u��j\��EBnm������?���;���m�����~m��܆6���ٰj��I]��Y��m���q���n�_�6�f�Cm�s�?~��羅v��쥒�r�\��m�w���~m���^7��vw}?~m���Wm����%���;
[*������x�o�����m���q�����_�6��k��b����k��|�^G�;��d��7�?;���w������ {������ ?3�����$F�SfYswl���hfR�Ѷ[,��d�FK��[�ݩ��M�z-�)�^�.S��5l�0ɱ�X�������se"�=�v�,n��U1�e�, E��zE��f�݂�j���iK�5���mƊ8:^Eӌ����j�.-B�S�{;FY��r%�<2�M�qEƚ�ͻ[u!�Yv��c�6������^�{�����z���z��O$��%c�u�c��Y�J;m�x��;�$v�2W3͜�������Igz�g=�Wm������m�n�1��';����zG���%�������sw�����JH�{�m�����������m�z�q�X��W�ͷٻ���|���ߛl��+���sw�������TV��bn9a���9ݿ�6���W-���{�9m�W�QL����7m�����0*���ik����gwq\m������ͷٻ���o���ߛl�j�qF��<��g�OM�\�2����:�ۍBoRgD���h�Ka�n��� �����w�wo�.
���u��n��"�Www������:䔶U��m�n�3�/�_|�@?"�f���s�s��=���ݶ�}�~_�6��k�aB}I#,��m�s�;ۻ�ȫ���d�w�wo�.
���	;�rɆ4f��ֳ9�o�Eu}���m�w���~m��܆6�|�v���oH��I~-B%��m�����~m����~m�����������ozkП���'uj-؄�h�m�ʽ��,ilƧU]Z�l+�4(F��ʬrZ�;W�ͷٻ��m������m���g�*֭�~����FR3���+��8�6�{�������U�������dT����×��-v��n s{� ���X|����:f�2e+�7�z� ]�M�̩O1#��ü<J�x����ɓ��~T^�* �;� 9�ۀs�ܖ�-�(�R�R슐똀69�슐�Y�vk��&�c�땝��H�K'�]�s��\�N.��O��{�O���g�T�U�et��@�vEH�*@k4���eM[����?sb�� �1 ����'9y�_3(�����ȩ �EH��W����� ����]eV9-DnՁ����w~Tw�4켚L�2��l̒J(R�!
�Z-J$�"IP��P��
��~�� ?{�g��¹,$� 9���G1ݑR슐�s�u|��VXf�qx�3���k�ݷlZ��&���x��X[�t������Yw���V����?��� ;�*@=�R �s$YW���m��*��p��ŀw������ ��n�����S��(�R�V��Ҡz�h�L��{�4�v�k�1`�AI��`9ݸ�����q`��,YӺ'S���� �� ��@v8�6EH똀>���ԒZ.����W"j�m��QV����J�Cn&I��jFv�GF��e쒸T�t��՚;s���q}b�m\�e�x�R��}�o��� 6�,�!�����v�3��ܖZ0U���:4�j�f�In��/��' ܫ��ş=;Y6:��ϕ�.n��g��U�]=��|vt�9���C����ܜ�|�j���gE�f]%���D53Y���?�ns>�u2o�i�
�Lqphz�v�Tz�;v�g&���»j̧�#��톻rU����ʐdH�����؀%:��2���Հo7s<���l7�����?owgɟ'��2��sY�.�����%�b^��fӑ,Kľ7ı,N{���K�g�{��&|��g˳{!�+��-y�2�3iȖ%��E j&�{_���X�%���~��Kı=�kq7İ?5^�fӑ,K�����Y��s35n��ɚ̩��%�bs�{�ӑ,K��}���Kı/�wٴ�Kı/��eMı,K!�쟟��.��8�Z�c���yBe�;�6ӝ�k�v��-���]�k��y![Sw�I��� �	9ϻ�D$�{"z%�bs�{�ӑ,K�����'�RB+m>X|��gɟ'�wsi�Q6�i�L�b_w^ʛ�bX�';�p�r%�bX�ﵲ&�X�)�-��ѕTX��[�/�ɟ&%�}�{*n%�bX�����Kı=�kdMı,K��}�ND�,K���]K}���3j�eMı,K��m9ı,Ow��q,KĽ��ͧ"X�%�}�{*n%�bX��ǴOMY�j�Y�Թ�ӑ,K��}��7ı,K߻��r%�bX��ײ��X�%��w�6��bX�|�7Dӕ?�$Ʋ*�l��K-��U:�^:QӲ�K��\�<	�����NM\�6[R]kXD�Kı/��ٴ�Kı/�ײ��X�%��w�6��bX�'{�l���%�bw���L�2kY��ֳ6��bX�%���T�Kı9���ӑ,K���=*n%�bX��wٴ�Kı;�kyfk%��պ��2�2��X�%��w�6��bX�'{�l���4
QT4H��BB1��iI�Y��sLJ3��KowF�-W��2�)H4S���O�1!HD� �M�|B�4�0�#z�,�@�n�h!��,�0B�AP�a�$�A�m�� hIj:�΋���]MuB 'F[��7�Q��Ќ��A�,R,d @�:�M�	�ް�.�EJ�D��ևʟ1l# �1!MAFeCHT�l &&�BBQ�m��(XҒGb��/3x��	�H�c7F@�����c�D�
���iDh"9�<�Q@ұC���"��v���D�D�%�y�l?�}Q,K��W���ϓ>L�ww��e��(�#���iȖ%��H��~���bX�%�}�6��bX�%���T�Kı9���ӑ,K��ۚ׳P�$ɢ�e�3��bX�%���m9ı,K��쩸�%�bs���"X�%���["n%�bX��w��\�3Y����I\^�{,�m��la��%&+�Ċ�����BH�I$������=�%�~���7ı,N{���Kı;�kdӑ5ı/��ٴ�K�&|�OBDߙR������ϓ�bs���"X�%���["n%�bX���iȖ%�b_��eM�����j%�zt��~��fj�Y�Թ�ӑ,K���kdMı,K���m9ı,K��쩸�%�bs����>L�3��t���%#���*>Yı,K��ٴ�Kı/�ײ��T�K�����6��bX� �'H*�Z"VDB(�R!R%bЀ(`@������PbYA ��=u�Oܽ��7ı,O����!3&]k2ᙗY�ND�,K���T�Kı9�{�ӑ,K��}��7ı,K��M2�d�'8˵�;�!0�	�0����v��p1�0�x��u�uv�l����NF�Y�H+u����oq������6��bX�'{�l���%�b^��͇�D�KĽ���Sq,K�-���X��7dt�U�/�ɟ&|�N���q,KĿw�ͧ"X�%�~���7ı,N{���Kħ˫�ٶ��1±�Q���ϓ>V%�{��r%�bX��k�Sq,K���ND�,K���D�K�g�aӺڪ���� r��~>L�3�Ŀ{^ʛ�bX�'=�p�r%�bX�ﵲ&�X�%�{��6��bX�|����z!��m,>L�3�bs���"X�%���["n%�bX���ٴ�Kı/�ײ��X�#>X�I|��HK��o�H����x����:����z�:����g�r	�.��oZ;G��9��4�w\�г̝��:"�!5�o��_l{�j�`*��Fzw-�㓎�Y��2[�������2�#u�cc4eL&o\:ۦ�=�[��nK��3��6F��Y���8�3�^`P���0�D:Q�-l�;�`�皽�I���Χ�gYی�`-��ݷ����?=ܚ�ߙ����B	���_��j�)��%���`x�c/+:u�:7PZ8��q�ۧF�k���8��X�%�����q,KĿw�ͧ"X�%�~���7ı,W�������3�ϓ>OwH�IBR;k�5�"n%�bX���iȖ%�b_��eMı,K���m9ı,U�E!��C�����q���%�&^fe�fm9ı,K����7ı,N{���Kı;�kdMı,K���ϗ��ϓ>L�s�r��ݶ��̹�Sq,K��}�ND�,K���D�Kı/��iȖ%�b�6m,>L�3�ϖ��J[mr�Mf��r%�bX�ﵲ&�X�%�~�}�ND�,K��{*n%�bX���iȖ%�b}����XK&��9�����]<�n�;Ć�G]�h���Xg�N�u��E��&��{���{��7��{��r%�bX��k�Sq,K��}�ND�,K���D�KıOzw[��`��
�����gɟ&%���T�6Q�x](?���9���p�r%�bX��~�ț�bX�%���6��bX�'M{R�/���Y�Y�Sq,K�����"X�%���["n%�bX����r%�bX��_��>L�3����&��9-D.a��Kı;�kdMı,K��}�ND�,K���T�Kı9�gʙ|2q���e�3t�!TH<�13�k��bX�%��6��bX�%�u쩸�%�bs���"X�%��و�a�gɟ&|�qn���),���8���g��=�+D��Ǭ��m��8�7�V�6d!��B�ub��߭�7���{����Sq,K�����"X�%���["n%�bX���ٴ�Kı>�������Z��}����ow���p�r%�bX�ﵲ&�X�%�~�}�ND�,K��{*n'��MD��;՛j����:K*ϗ��ϓ>LN���q,KĿw�ͧ"X��Xh?��m44n&�^��쩸�%�b}�߸m9ı,N��絚���l��e��&�X�%�~�}�ND�,K��{*n%�bX���iȖ%�bw��ț�bX�%�g}pљm�˙&����ND�,K��{*n%�bX*��߿|m>�bX�'��["n%�bX���ٴ�Kİ};�����2b}v_n��uoj�x5�\7lF \*qn�p�Ƹ��X�L]�g�f�ݸ�%�bs���"X�%���["n%�bX���ٴ�Kı/�ײ�&|��g��qv!l+,rZv��r%�bX�ﵲ&�X�%�{�}�ND�,K��{*n%�bX��}�i��3�ϓ>OwHȭ�t�[Gd��n%�bX��wٴ�Kı/�ײ��X�%��w�6��bX�'{�l���%�b}�����.��p̗36��bX�%���T�Kı9���ӑ,K��}��7ıs�C��$_ƾ������r%�bX����Ժ�r�jkZ�f\̩��%�bs���"X�%���["n%�bX��wٴ�Kı/�ײ��X�%����ߩK��ǳ�Vҡ��hWn����픢N�6b�&Ʈd� cM�1�K[T3����X�%��~�ț�bX�%���m9ı,K��������%���~��Kı=�o��,մ�K��3��bX�%���m9ı,K��쩸�%�bs�{�ӑ,K��}��0�3�ϓ>Ozw]QZ��ЎKn|r%�bX��k�Sq,K��}�ND��D�O{��D�Kı/}�ٟ/�ɟ&|����=D�X�9mi��%��j'����iȖ%�b{ߵ�&�X�%�~�}�ND�,K��{*n%�bX������Yu�&��6��bX�'{�l���%�b_��fӑ,KĿ{^ʛ�bX�';�p�r%�bX�D"� Oz�59s��ۤ���S4�)Pn��/fKI,��I�l�d���o�����X�S�C���]�F�m�CJ,[��#��.�+�s���w��������b1�g���rX��g���p�cd]�Aƺ��E�m��눖D����8�;��7��$����]����q6��O�+'$��,\�ٖr�D%��u����Meh��M�U���S$7��&je�7ixs� \��u�:�շ���p<'�����y��̋�=Wb��$7ow���bX�����m9ı,K��쩸�%�bs���"X�%���["n%�bX����LɗY�0̙�ͧ"X�%�~���7ı,Nw���Kı;�kdMı,K���6��b]�7��~�Ϥ"�.���w��oq���ND�,K���D�K�B�������r%�bX����*n)�&|����$��kv�-�g���bX�'{�l���%�b^��ͧ"X�%�~���7ı,N{���S>L�3�޷�%aS(ӕ���,ı,K��ٴ�Kı/�ײ��X�%��{�6��bX�'{�l���gɟ&|���U�;lV�#*�9<���$�_L�p�n�q�5����{I��ј��-��s$�ֳ3iȖ%�b_��eMı,K���m9ı,N����!9Q,K����ND�,K��j���Z��Y�Y�Sq,K���NB�16-l�B�A*���Ex�'�,N~���7ı,K�~��ND�,K���T�Kı/O��I|e�\̓R�ND�,K���D�Kı/~�iȖ%�b_��eMı,K�{�6��bS�ϓ��2)jn��`�,>L�8�%���6��bX�%���T�Kı9���iȖ%�bw��ț�bX�'};��fd�fL3%�ͧ"X�%�~���7ı,N}�p�r%�bX�ﵲ&�X�%�~��ͧ"X�{����~�;��ùi2Zt�p�7U�3^��W�b�β�S�'E�Q�i��N��ke�ʜ�bX�'����ӑ,K��}��7ı,K���m9ı,K��쩸�%�b{�޵���,�55�Y�6��bX�'{�l���%�b_��iȖ%�b_��eMı,K�{�6��bX�'{o��e�e�)u���aq,KĿ}�fӑ,KĿ{^ʛ�c�^�QO��v�}��ϸm9ı,O{��D�Kı/�;놌�l�\�5u����Kı/�ײ��X�%�Ͻ�ND�,K���D�Kı/�wٴ�F|��g˪lmm���r�"[_���bX�����Kı;�kdMı,K��}�ND�,K��{*n%>L�3��.�YY ����T돩��2�q���+d6��W\ƶUq��������Y5na��Kı;�kdMı,K��}�ND�,K��{*n%�bX�����Kı=�ۓFf���a5��aq,KĿ}�fӐ�c���b^��쩸�%�b}�߸m9ı,N���q,K��w|S,̚�Ɇd����Kı/�ײ��X�%�Ͻ�ND������kdMı,K��}�ND�,K��n��]�q�J��ɟ&y|����}"X�%��~�ț�bX�%���6��bXO0� �S�#�D�s_���X�%�����k�)�2�sSYu��iȖ%�bw��ț�bX�'�w��r%�bX��k�Sq,K�����"X�%���\�]9e������'��q���0n+O��tX�%�a�qJ5�,�[�v�}���bX�}�siȖ%�b_��eMı,K�{�6�>���%��~�ț�ϓ>L�?i�uEki�KU�K�/��ı,K��쩸~X�&�X�w��ND�,K����7ı,O�ﹴ��3�ϓ>]S`Ͱv��Z�Kk�`�%�bs�{�ӑ,K��}��7ı,O�ﹴ�Kı/�ײ��X�%�z}gJK�c.e�V�ND�,�Q=���Mı,K���m9ı,K��쩸�%�bs�{�ӑL�3�ϓ�[)jn�[Y+�?�%�b}���ND�,K����_�� �'���pI���$�H?� �+�� �+��@U�� �+AQ_�PE�U��U��E��DA�E `�@�E�$B �E b�Q@�P,TE����*���*��� �+�U���Q_�TW�Q_�E�U��ATW��Q_�PE~PE�1AY&SYs�8�O�ـpP��3'� ano� �  �         +@   	 4��I@ �P�D��D 
  
@PU*"� �HP���QR(I�R�  ����   Ò�@    � >�b���x�ɸ����zU�>��RŽisۯ��MO��ۤ��;��|��)M1@  M ��  t0R���@&�J=��
�4�Z��Y� �P��
R� 
/cJ@ �     �@� 4��'` � ZD6ʬM h� s�)�vEQĭ5X���H, p()����� �ŕM��^x�{Җ����u�W{���rgm8 �g^��n^����޷+��ju� <>@     &` 列��N�{��n���{�|^�{�������N�{��������}o��k=�>���M;۾}��;���ܼ��  � �` �������m[�����s�G:z���[j�g���{��^O{==o� ��
 1 
o�}i���^�������^���{]�	z���w��g��=�����nW���wzҼ���;ŝ� �Ͼ�Ε��=*���kͺ�o�/^�&�^�� >�K���{�__]�n�{<�z^ �  ( �� �}5y�������/�u:�Z��� ���]Է=�C�LEz�O�W3_  /]�Ҽ�y=+�� ;ʖm���g_K�t��YK��L�vS��zo����{������� 4`����iR�  �'�UJ�=��C@@��T�iQT�F�"�����R�  �!2��@ N��-���?����s���+u9�ݭ�I&�b���4TWJ
�*��z*+����PTAS��/ļ���&�_��P%WH�w#U4�y���G�k\�̺v?� �y��@o�6v\BS|���Χa�X=c�gw�Yq��!C.���Zz1�&y�0$C�~�)�[ov��gt�Bg4w�t��#��Í�|;Kvć������-��Gk�M|����5�pt�'%.B�]�h&�s7��6�asYL��|����K�Ä����P�xO���99��ފi>�1����M>7�s����A�^��y�G3_f�k\8oA
�c�_��&�wߍd�Ϸ��ٓYIi�4K��4R&kaoI.i�#\57��X[���2T�ӳS��~���Y�bC�
�ka���s���J%$T�)�32�*�u>���Aԫ�s���42><�ư�!	
�|�F��1aVR����������~f��XP�BYՍM�a4abL>P�> ���t, 4�8��X0�&������$uB%Ԑ�i�HR���\Y�E�aZ1#��Se�2�,��Hô� ���~3$ �����HB�J�`��#�;�$��t�|͕ݤ����N�b�o=��i��	RX�0� FB�#Y�zIZx8,�$k�������<�!bB���B1�#,$ɐ3Q̇u�C9�ǜ��	��C-��O�$�8= �1�BE�H���ϙ5�L)ѭᜩ�� 4����B��^kT�h� ��� D	W��
�+�r9tڀjH\X��p�N�1��W@l�>:t!N8M��9.ivC��GP4$1�V�
ګ��W�0#�HSf���Z�$�iHa��"fw��̔ čQ��O����>#R��	BA�!H�XD�햎'I7�
d����a
�(B�@���Ul�.�"q�B�Q�A�h�ˣE6E`V0Ӡ�@"�1��X�v$)�X�meB	aR4B�B��aV8v�P�Fٱ�Hh��Pަ��G��H~G����c��S�#���N����)R��1�v2ɧj�4����U��v!�G8�4$ğm�� W+k��ŉWN̈́/�,�H\��[�~�-���
B���|t%glo��HA�+�R߻t�dr�D
�n]RL<g~���u!X@���cF�0Ѣ��3F�^��&l�i#	.0�Ha�9s�PͤX5��}u�]��a���S3\�8��8i��0�;��:9���#߸^kl�Ip��{�f����[3CL&f���p\�%��p%2B\40c�0�ݟB�C.j��5�,-��`�N�7599��7l�G4X�%ָNM�c�l&����Jf�\Ѱ���uu�	�Ѳ7Z�.h6��}.Jh6cϹ�K�[Is[ɠ�Ѕ�����\�˚����L��˭�.i�5Ú�N�sf$��9�h�|�eޒf��g$)�F�0�$�0�	
`K���a���M��y�o>���_|�h���]��aM�WS+
U�iLH\+-�A᠘h����+Jq��\6|�Cz�i˗�r)�\�ۤ�S��)R- �) ���
jE�anMl8� T���x$J�B�.�۽�}��=���@��HE�0b"�H�� FX��`SJ�,
B�4�����5
A���`�H$��*J�"A�����@p4Ī�
��e�I[B�5��sP�p#r�fX@��JK�&eV����m�$�b��$6�F�2��kx��0��u��5y��	�D��A!*E�#@�Qbѐ�M6(a(�]���ނ��}�i��sm#X�cv�g4:����7�k]%HV\�B��7�[��ַ��ƛ��H�ߓ���ެ01b�3L̎��HL���@0+���ŮM��(Kp��hѯ�y��Cr�A��b�:4l�M��C�۶j�X�1�)W-0�#j�Ņ�+@�V4�0ѽ�ɲA��q�|y���x��f��{g�݌�:v0&����M�'2W�l�h�.�s��(��b���4C�6m];4<��)`V�n	p���\P�[��e�vpϷ�9sZ).R2\9��F�O���CO��~3.��7�f^	)�(�.pː�oBA)��SA�5��f�u��4��\7Ձ;�Yˠ��I
c�+��+&��D�@��}���o[��p�v L9�Jvx�}�$�(Fc
D�?@�`h�>���]l7���}.��8g4|��HĄ!U1�rHSP��#�&�d({ﾺ%8*�k��*�4xa�p���`c�08���8� Q04���#pЛ8`Ƙ�C|� k[�k43�
�@��(��,"�i�pX5"6@`����ώ}]�O�4`h�S�� �#�#A т� W]	
d��e�HB%�5�}�5���,�B�B�r���@H��N>����W<��\�'&��5�	a���I�G,&����f\�����i,��
i�!L4» W	MgC��l�̔%�!R\�I���0����}a�7�5�1�Hf�H�����e`�to}/��J�B�K��L�a,0�`�.0�.�.����a�)
@�+���,���9�b˶�S�| !��8�fZ}�(Fhw����s��7g>��m��ʹΪ��g�8��+U�������L ��1"т�cC1�T0�FH`Q!cL�X�%��P!HS����cLHSxu�H��HW��Q�SF5�%��|� k)���Ʃ*��Z$H�X,V(@*��@
�!(A�B����"1 �!HЉV	% �"�XъF	!  "ĈU D�Ĉ�"	�E���T0�I�ĉFD0bE�A �X�,E�q��b@RHD  �����\։D�P�0�a\LH���_&�Bh6萍0�!�2�C2\!L�F��4o��La �7��k����1 Q�H�X�q�9��ᧉ�`jSLi�d)�R�˔��]m9trrp%%2�p�~�HD�`D�[ �"HJ�(
� u4
0����lv��ЛEڡ�`���a��D� mB\]H!��SjŮ	�� �@��`F�f�ŐJ�����A�b�\��`a��j�)�.�k��\tl�͚$�sF���ݼ$H��NÆݛ#Lѷa��p�CC�xJ�*l6;�L4�ٲ@ă\v����2P��r�:>ϩ]�G�J����GŽ���t}�?����*
?7�E+��$n|n��I�������}�\�0���nsd.:���I.i����c#!YIF4(B�[���J���T�Մd�(�F��JƆ)R,P�F!��������$��Ϲ�r�K��o7/.��ۣ1�
B�6���k)�����l�k�␦�J.��I�J�ƌ
��#m69ϊ���9��2\Ѳ6pH"�)��؈�_���Qj�#���X�K�L/Ĺe��ąaFP�3��9F��c*�h�A�!�$HRSHu
�z�K
`�n.t�B���Z�0h+�"�]!�
i!	�)��"0v��R��|��o������Е�2���r�.�>�D(D�\;{� �`      �   �  �  Y`����l� �� $Ioku��ඃm� Wf���� �l�x 	 ��@��������:@9J�nz�@ p�I��6ݤ���m��n� �i�Ͷ8 �m��k�[Sk��P�jCm��`��6�~0�U�x�@R�Ͷ [@��6�v��x�Ts0U S������&� �ݻ16Ž@K-��:l�q�J�cC�rWm�� �]u��b[b����h	T���m�Ӥـ H�>��� ��m�� \���٭��    :� H ڶ�im    � 	 �m�� -�e��Im�hv��خ���Wj��D� [M�a��      m�  Hp mm �         [@ $�R6�m�mͶ>�m��!#�fض��@  �n�m�p [A�$�������p  m�6�8[@���� m���i2@�i0m� ��h��ԓc�vZ��P�@l��vڡ!� H� m�l�    �  ���vP -��$��l�l [Cl�[m��&�  � [C!���[j 
����[!4�@� $�\��Ã��   $ &�[cm��-Քpm�m��-�Ͷ[;
Yi�jU�F��R�'�G*�]T�ð���  �ͮ�im�v� ݼ^�����H+�ڦ]�\��w�������:I^�e@���@mm�Q;����m#�IӤ�n� ���M�����m��-h�����v��`�n<B�G�$�g�P:XZ���9�]'-�#  4�� h��(�P�zq�f�Y-C.���j-lT���(��` [[l�mt�N�e�t��Z���؄����&�mە������:�-�6�pl]Z����T]mU*8ڱ��H�����^�%�Q %�૭����VZVW�&�A�'���+T�����kj���P ڧnU �� � p�D��m��M��pӤ�t�j6��zt�-	�ؽ[��hi>� �� �m&�@�$�� [@     �  l m��8-���@��   �� �L�x��8-��p���r��h����  6��geʶ��^Z��j�m�Kgt�`m�C����V����eZ l-�Ix �` %�m��cm��� $� m�$ ��  � m� ����   l �  m�-�ݶm� [Vյ����J�kέ�h)�t��wI2�  �-�9j�	m����h�@�k"����a� ���#��m�t9� m�   �`l� |   p p Hඛl-��mm�@    �`  ��� lh  6�l   �ă�hv�Mscm�6����ඖ�E=�¹��c�sU[��f�H� �٧l m �h�6� m �` ��}���`� m� �`  [x     �l ˭��C� � p8�u�Y���c�:���L�Ihrԛl�	 $   p$�6�v��"�����-�hm��-��d����$��\�wE pm�i��� K(�7�o�l-�::MK�)���
ۖ-���m-�$� � ��  -��p ���^�m���M�H���   kn6�C� �h�	���}��'͐���xt1UX�2���o-���:@��c\Z�-�wn��s*�I��pγzidt��-� A�6�ٵВ@j�l��U��`Aԯ)�O9"�M�9��g�m�w-UVҭt���(y�]%�����-P)z�����ne3d�T���̮ǌ��붜r��.�RM����"��F�8q�g-@V�B��?.ŒZ�6�\�q)[a �lcfZ�Ͷ:8y=n����bǍ��;'Uv�������m�*�v��J�e:�� s�2,��[`��6�M�v�6��&U��;v@}lWnʽ��#��h�}�ײַH�Ak�6:�z�[�p�b� �/[б�9%٩�bR���E@�a��*�e�l�l�v;ɡ��Z����_�+��v���I(m����3g��Xg��ASY����2p $�`<-��W-�i �J-�ɁSlH-���H�pk�-��`����:�\�(n'R��Y%sm�$�����!�E��9�֯� � ֻF���f^V�
Y���b���۳����U�ݳ�N��$m�pԩ���j����p�n�.XE�5uf2֣t5���� 	t�� ۶6�m$�$p   Ѷ�,K�^L� @6�mu���:/� L&S���U���і�]z0;�퇒6��{D0[ն��A��r�h i6�[R H �4U�z��@nQ����ϛ|�\�A�Pe�Wm�kA/3P�J�v�y��:#Gj&�iv۞m6���6]�ι%�� � | m�� 	��ᲀ�N�+�@FF�VY��Uڱ��,�{c����ںWL7l�rl�s� p��m:[p���m��i�[�λAn;U�[���X�2av8��� H�kim�s�E+�N��g�a�J�:Yy�]��x��UURc=�!k*s�lڵh�^Vv<6q�m
�6�n4�3����&�s��؝�zV�[m�wN��X�� ��MmK�# ޾h� ��]�$ �@�j��Gkm����g-� ���I�h��.��#E��$/RA�-*�mɸ­U�B@ h�&��zKit��I�	*˶�۶i�v��@������Z<��UuUT�  �k�%��ZR��U%ڕ@�8���m+�D�\�U�[Mڥ �UHqi�����H�� $���%7[r��$tv�� Ӛ֐���uTWPRҲ���k�]m�0  m�ݶ�b� ��m��%$�q]	�֛ g�޵��:��m&*�|�qۍ�`�@*�[mԘ�l趀� x�i%�ۤC�g��Q��g��Y-8�Nm���� ��UR�[M.�a��j�x㞖 �PͬcT *���;�E��,v¥�P*��m���5UP��t>g��@��V�-�z��H 6�	�m��4�m��if�/]n趀�� 8�'^��X2-�k��&�g>i��7�jޠ -����Y˛`[\�-��m6F�G���im���N�i�P�*6+��p��+m��$��m�A@$��9[+d-`�kh �%�,��,��$�Vmm�-��mY��:vrF�ے ;i3i-�'Z���i�vH  �F�Y$����9� ��&� h�p�6̈́�	G ՛`mq6-��mm��h�	����k�rl���[`K( >��  � �"����K[T��R��l;�m�R���6�l*��]@U��\<��gZ
���VR�;`j�ge�*���M�M=4�m�X7l:�,�]� �����ǩ�6�#fK9,��0$㦨9U;<���Km���mp��[I   ��Vͽ��,��N�]��p �*� ]H`$e� �� �� [R��-���m m٤�F 	$� հ.�m��^����q�ÀN��h�!ĉ��  kER��Z �lm$�F타h�n�p  VÄ�  [@����߾�A�kj([m� $�l ��� H6� $8 kX&� h   [��m96�[x 6� l�$��	 l׫��M�{[�kH��  	� 	m�����iz�m�i��  ӧe�p�� H �hh� ְI�m�d�j�mσ��cm�G�$6�d[2��u�6��z�Z�����R����e� 	�RҢU�t^�&�����4]��ԜJj�l��*�f�pl��gZ�&`����n�$�d�L��f��N��nZX�lJ��#-UU_��}ָm  �� 8� ���%�l�m�H!j���P $k��]6��dZ�o � �u\lm@ յ�mwl�(�F�jw<ك���ݠ�j�jV��]R��� iI� ��(�m����6�T3R�)�T���$  	���� 6Z �[KL�+m��`�BUʹ�������H���6�R�@8��m�H  �.�w���w��
B"q6�Th�J��O��8�� |��F T��(�z��\ ",D�ľB���x$<�Q��#�U^���]*�������@ڎ�CK�z��v��� 4��>5�W�!�/����+�ʋ��
�� ت!�� :�p(�(|�"0Z�v <v(p8���u#�h>;���h�PO"�*@`)�u |� ��E��E<�.�W�(%@:p"��	�E��ت�]3J�ʎ����(���H�T0�F�mA^'A�!���X��QT��E #�*��"�|�E�9��yjt"1 ��>Q6"qUB��U` `��C`�D��
D�lA��(-P�V
|�ys�Q� y�]� mGI�hTΠ��E��h �>

|?����
<v�TGͪG����~A<��G���(�SH#�� "��T�v�iy	4!�@�ꪪ����UUPq2�� t��5��O'Z6�b�+�QAZص��7"�%ys���(ϑ7<@3��%6�C����Y-�`�6mw�j�Mi�`e��z�a�N�
��ExƧ��ڰumҽ��K�Ƭ���s���\�ڦm�N��i�{@��Z%�kkS�t@��� �ȉ��]��J[�T�,�ͨ��v����Wal�4�Z�;6�զn؀�VkXэۮ{^�ӳgU��;X�|� T�4�:�t���Xp������Y%Uu�Z�s�%vGB�Y�Sn=
N沲�4C�y$"���b�	�rҝLMl��[A�;	TR���KvNeU���
�L�h�gg�����^0`J%N�ݐe��Uu�*q�	֭&cfP�
N<���+s�-%���e�(VXFG:�6�\�B�fw���o`�.���t���M�6�w�Gkri#����������vV�'�/.�ó����Č>y��	7�V�m���4e6�J��gZ6��1��i���iYU�6��(��{n�&�]�3��W�Ӎ6bke��`�p �uĉlnd�3��Ս�1�z�ul�H'ֳ{q�I�^��Z˴�
����-�ò'a�f�ܴ���u�:Mh.�
��q�,����1�Xd�9��]�ҕEu�vmF˞����S+��C�û�����&^ַh)�.����
ֻ{v��c�㞲���=c�}�����q FU݌�9�n�e4fx�9݄z��X.�i�����WP /�dnrE��k�]��8꨺[Ms�çv�^ݽ8��6�9�1FE���Wv��cNhN�-�i�s��q����a�W]MJ�ڔ]V0΋����u�_ YM�N��{�����%��.��]�7�F̨�5�p�<eHD��6pe����N�ڶXl�ŧG]�3���9�M� Ƽ��U�\Yv���뛱<�c3Z���u��T|���/H�	,�
+����� �0Cȇ�&�V�O(������k��s]�l�ڑ��t��q�q�v֢x݉�J��gf��{f��'�9��nRs���9����U]�lt���#�C�4ju�\<�����s�g<�-����;Z������ݷ����#�n�6�����ݽ;���3�\E���&n�)W�`ka���T��ۓ��,�"�n��d뛶���w�׽ǽ�F6�dw>�;S� ��+��˅|/
�	��m�Ce$��?C�޺�>[���5�«����u`gw����������@z^�]�G�&ξ���guՀ}���! ӃH���1f�@nkP��6��z��֪n�&(D�(D�77�������v�1f�>[܇R5*8��IV�ܡ�z������B ln�.'F nӏWa���ہݘ��n�PD��k��]kG`f�����Y못������@d�@nkP��6� c�S7e�MPQ5SUS`r9ܛ����$ƚK
%��D`r{9͛�w��������v�I���*
H����֡�mB:g'�Rg_R�U7bPmH�)$rU��w]X.�v,�v��Ձ��[i�n'ӎ)*���t���t��֡�mB��]�۷,e+�WU��u�.��f��d�h�;eKn��(���9!��������B�ڄ���ZjIJ�(D�(D�77�������v�1f�~H��y:�)�TQID�V;�j��3�6JI!���4�M<M6�;�6{ܵ`s��5Q�qԩ$�����ś���޺�>�� ��iJq�P �����7����B�ڄ��G�}8o�W�/Z&�O8��a�Yd�6�m:c�J���<1��\L왧4mg��TL�m���P��6��z�����Z���UD��RrG%XguՁ���`b��`no]Xn�����"r8⒬K�H��H舏�^�P��|� {g�����H���>Y����$������J) "� �U1hAOrs_���s����֊a�5r�e�] 75�@{5�@z^�@��[k�e�
)@ER�SJ�UL��I5�"���X�7�3�T:�ywId�ED�t�ɮ�.�����B��� �n�����MȔIJ��R����o; �n��� 3[P�1멛����&���kv��֡�ڄ��;���G��P�NK~�T�{ބ��K�H5�@c֪�왈���NH�7������������krN��lܓ�8�
�A����S 0X�#$Q���"H���z�rG.���φ��h+��c..4+��[Xwk�����s��r�|Ϡ'� �b6C��(��m�v�O��l،;=����B���]sy&�{Vn.|� ��[Αiȷv�v�{"�H��^^��p�Yocԧٵ�@��v�:2�'�Ž�Ț�'k8X"D�]�4pY�xkc�]�����%Nj�f��F�m\�dAkf�<h�3��q1�ܮg
���K�Yl���v�N~|~|��2�Ȳ5�����l��@��sZ�n�ڻ�����$�N; �{����u`f�]X.�vٽmI)S��&�HUݠ75�@f�P���t�=���ky�0��QJ#�`f�]X.�v��Ksz���޴܉�qԫ��@z^�@����B7Z���w{������J�V�mX\*u�ݮ �{QO�.7]�5��uι痴k��p��(�$\��]��׀1�ZsZ�n�Oo;o%B"���"rX��W@g �q@�S�K�of�^�v��K;z�R�d�RrG% 3u�@z^�@����Bj�r��NB�q�%X.�v�{����u`f�]Xڻ�ܦ��$�N���������k|��z���}�~��*��.�{c�d.Q�ó�9���wV\�]E�<ۮ�ڲT���ۛ�H����@nkP��֡�z�������h�)�TD���X��W���I�ϩ�����BwZ���K��jU*��`}ܛ��d؛ƞ&�[�R7�u`f�]Xv�%5R�����n��� 3u�@z^�@b�䔀��P�'���u`f�]X.�v-�vg�;qE�)(�8m�ƫ�7f�o=c7k�bz���ۛ�{��cj@PL�*NH�7����v�1os�77����m9I(����r���z�w����ɲ�� ��kj��T�gy���$�$H�q��ޤ��� =/] 35����&*��&���tD}/_z�� =/^nM �� AD E��H=�v,��J0BR�$�G*���P����+�W��}Ԁ�֡ �u�����s�6C�=˺�<b�m�/'<ӗqV���z'7\X��nL%��l��;�=/] 2u�@nkP��mB Ǯ�H�D�
Q���3{���~�UI��}������fn�K���n˚�@nkP��mB��� �n���ڐ$J��9*��>]��7�X��Vwu�9M��!Nj�����kv��֡�ڄ���_�fr�S�"��CI~pN�K�����9؋6�q�Өm�k<,q]Ck����{=<�x�r�͕ݴ��v����Ҩh�b��F~Q�.�����f�BNJ�h�ʝxk�r�:KGN2��gr�ή�X+,��IvV�=���m#�W9+ǧ`W$c��.l��$�kI�5�Hb�ӱ5r����1g'&2z�6�]g�떸��c��$*�Ee��{��;�{�|��L�:뗺�����|0m�dļ-��L��+t��lC$<�3 ݎ�i�.�殘����B5�K�vf��䢕7De)$�77���� =/] �����Q7A$���wp]\ 3[P���t�3[�滫w��$J���G%X.�v��U��w-^(���FZ��j�{��?�~�̚��M5?=ߛ�oqĳ�����bX��Qc������%�b{�����X�%���}�Noq�����g����Ӌ��dܛlލ������1����V)�0ݲ���%�ݥ�Z][����SWZ֓q,K�����"X�%��_l���%�bs=�f���H�@��TՍ@�@�w7钰J���S]�������ow���Ω�l�#@b!��Aq\GQ,KY��6��bX�%�ﵤ�Kı;�}�iȖ%�c߻���kr3Mǻ���oq����6��bX�%�����Kı;�}�iȖ%�bw��*n%�bY�??~�Pn�e��g��{��7��g}�i7ı,N��p�r%�bX���ʛ�bX�'3��m9ı(�;�5HP�QR(�&������;�}�iȖ%�bw��*n%�bX��wٴ�Kı,ｭ&�X�%���ww����������yE�ͭ�9�k�܌]���nM����J���N%h�����ѫ5�Y���Kı=���Sq,K��{�ͧ"X�%�g}�i7ı,N��p�r%�bX����ֵ,�4j�љ�7ı,Ng���r%�bX�w�֓q,K�����"X�%��_l���%�b}�ﵭf�Yf�**f���m���j�j�U5cP2ı;�}�iȖ5���|��Hb��O)t�G>P��M�{�!#	%� ���iy�,����i�Κ�?�s}�4<E]04I�̲�\I�&�����$e`�##_�+
i�\c\"\�R]��eps�!\!0�����e���T��V\! �%9�\r@X�l�B���c�@�A �R(�! �@H���E�#�YBr`bdJ�"��K�#/��(E� �xU�On4k������0��j��f�R��'7s���D�8�tJ
 :@z��DGbQ&�4��� :8
)�	EF)�Ț��_l���%�b{;�fӑ,K��=���R][��5���ֵ��Kı;�}�iȖ%�bw��*n%�bX��wٴ�Kı,ｭ&�X�%����f]j[��5�K�kY�ND�,K���Sq,K��{�ͧ"X�%�g}�i7ı,N��p�r%�bX�������'d�3ŭ6�+�nfe�t,G6���z���t��h&4�T�-� ��3END�,K���ٴ�Kı,ｭ&�X�%�߻���ı3cmCV5P5Q��و�D"f��+Y5��ND�,K����n��DȖ'���6��bX�'�_�*n%�bX�����Oɕ2%��k�˭�a5����kZMı,K���ND�,K���Sq,K���]�"X�%�g}�i7ı,NgN�tK-ѭe։�Ѵ�Kı;��7ı,N{]��r%�bX�w�֓q,K�P��P)���UC���{�ND�,KӾ&f�F�\�35���bX�'=���9ı,*;�bn	 ���ٱ$D���5��w������]��Jv�+mX�OS��g��W�$P��թ[t��8��Z4�35X�*f�j�-�����;�TՍ@�	bw���ӑ,K�ﯷSq,K���]�"X�%��{=f�VkVk5Mfk5u�i7ı,N��p�r%�bX����n%�bX�����Kı,ｭ&�X�%����f]j[��5�K�kY�ND�,K���Mı,K��}v��bX�%�����Kı;�}�iȖ%�bw�^�sFe�sZ�]\��Mı,K���6��bX�%�����Kı;�}�iȖ%�bw�۩��%�b^w��4L&f��kY��fӑ,Kĳ�����bX�'{�p�r%�bX����n%�bX��wٴ�Kİ~�,"�zzYd~��IݚX�I��\��΍���);s�7a�.��]&�l1c!���0�����~V(�(qs���FQ%�2��MY	�+9��Ɨb�:%��P���u�v�������6c�%�F�-��v3Zw�qz�P�C����5�=/l�S�v��F�5������/kGn1kg��mӤj�G9ص�ڭ�\��gM6��}���]��Ә�X�T�d�V��%��WF���=\���j�o`�dh�P�ێ^Ӹ��{�w���{������ND�,K���Sq,K��{�ͧ"X�%�g}�i7ı,NgN�tK-ѭL։u�iȖ%�bw��*n%�bX��wٴ�Kı,ｭ&�X�%�߻�ND�,K�>��X�륞�k�w��7���{�wٴ�Kı,ｭ&�X�%�߻�ND�,K���Sq,K��>����#]ij������{��7������Kı;�}�iȖ%�bw��*n%�bX��wٴ�Kı>ϯ�5�]1�ٙ}�7���{����w�6��bX�'ݾ�Sq,K���]�"X�%��^�17ı,K�����g$�S�ݐ8dշ^�'L�Գ��d��+���@ҕ���*�kFӑ,K����*n%�bX�����Kı>��f��L�bX��p�r%�bX����4f\�5�e���7ı,N{]��rS訵�MD�5���Mı,K�w�6��bX�'ݾ�Sq?!�2%�~����n�`5:c��{��7�������n%�bX�����K����;��eMı,K���ٴ�Kİ{�{2�D)�Md.��k17ı,N��p�r%�bX�v�eMı,K���6��bX�%�����Kı9�;��-ѭL։u�iȖ%�bw��*n%�bX��wٴ�Kı,�}�&�X�%�߻�ND�,K?M��u��  ݤ�6��7m�6�wf����%��^��*sN�%��Ʉ��7f�T�Kı9��iȖ%�bY�{ZMı,K�w�6��bX�&�����H�H�H�X�zH�E�ֵ�fӑ,Kĳ�����bX�'~�m9ı,O�}���X�%�������#�#�#�c��r
���s5sZ�n%�bX�����Kı>��ʛ�c瀩���E6�O'DN.D�&��}�ND� j��ʦ�j�j��Ϧb�*d�Z��ֵ�Ѵ�Kİ~��i7ı,Ng���r%�bX�w�֓q,K�����"X�%������˖���3F�q,K��{�ͧ"X�%���O{����bX�'���6��bX����&�X�%�{���S�d]i�@E:9�u�5�Ӗc���"Iv^�n&wb�JC8�<����?<r%�bX�w�֓q,K�����"X�%����I��%�bs=�f��{��7�����ꕶ9{N����ı,N��p�r%�bX?{�4��bX�'3��m9ı,K;�kI��%�bs:{�%�2[�Z���Fӑ,K���٤�Kı9��iȖ%�bY��ZMı,K�w�6���oq��~��v��g�U׻��bX�'3��m9ı,K;�kI��%�bw���ӑ,K��x�A��I��%�bw;�kY�5���jk3Zֵ��r%�bX�w�֓q,K�����"X�%����I��%�bs=�fӑ,K��=��1�
h֦��kcg�ƺ��O�=4��OUr�c���.frK�,e��ٗw�{��Y�=�~��Kİ~��i7ı,Ng���r%�bX�w�֓q,K����2�ѫ�)�Z]kZ�h�r%�bX?{�4��bX�'3��m9ı,K;�kI��%�bw���ӑ,K�w��}A�T�nKu������D��{�iȖ%�bw/}���bX�'�{�6��bX����&�X�%�������a�aY������{��"w/}���bX�'�{�6��bX����&�X�%�����ӑ,K����ˣD�a5�������Kı>����Kİ~��i7ı,O�׽v��bX�'r�ى��%�btU�#!���.��Rj�2j��$���;\rq��#\ʷ�b"�8�ҝ,�Rnwf�r�m�{���/ku�dB��b��\:;d�r���vů�DMg��H�j��GX0Iʍj'�b���v��ۜ��8竊��F���	�5F''O>n�ɥ�ӎܝ�pfՍ#B�9�bm��=�����2��J[��ܐ�m��f��'A!�\디�ݽ�I��KVkbk�i���v0.q�`g�&�YX�Tsz_i4D��IP�	+�����]h�v%�bX=��f�q,K���{�iȖ%�bw/}�ӑ2%�c]�����j�j�6n&��
UDMQ�3Z4��bX�'�k޻NC�r&D�=�߳q,K��~��Kİ~��i7ı,O��{WY3Y��f��55�j�9ı,N��q,K���{�ӑ,K���٤�Kı>�^��r%�bX�g��W5�SF�jk3Fk5���bX�'��m9ı,��Mı,K�{~�ND�,K�{���Kı=�{�nh�֭̔.���h�r%�bX?{�4��bX�'~��6��bX�'r�ى��%�b}���ӑ,K��=��jS2]f�s�yX�t]\��������R�-<���p�B+8nU3[���{�oq���X�����r%�bX���f&�X�%����ND�,K�{f�q,K�q��>�qYr�����{�7���{�N��p���B	 �(������Z
�(����Q�ț�bo���"X�%��}�I��%�bw�o�iȖ%�`��z�ѢS0��]]\�bn%�bX�{���Kı>��dMı���ș����iȖ%�b{/�f&�X�%�y��jK�d�F��Z2�Fӑ,K���͑7ı,N��z�9ı,N��q,K�����#���ow�߯��]Xk�j����X�%�ߵ�]�"X�%���W߳�,K���~��Kı>��ʛ?R?R?R?V��Ô�P	�*M���\��Z�����BJ:�^ѬrS��UZ.%�֖�G�w���oq�ߩ��}�2X�%����ND�,K�_l���%�bw�{�iȖ%�b}��]]]]h��S34f�Y���%�b}���Ӑ��ș����eMı,K����iȖ%�bw/}���bX�'�￈7B�8���{�7���{���}��Sq,K�����ӑ,t�ș�{���Kı9���ӑ,K=����~8��f�$+q�����,N��z�9ı,N��q,K�����"X�%����T�K�q�������r�aY������{��'r�ى��%�b}���ӑ,K�ﯶT�Kı;����K�q��~���F�^�MU�LW5�-�c�#���V���ֹJ+��9I�h��a.���R���Y���%�b}���ӑ,K�ﯶT�Kı;����Kı;���Mı,K��ԗD�n�]]h�֍�"X�%��_l���%�bw�{�iȖ%�bw/����bX�'��m9ı,O{ٻ�֥��Z�5�Ff�T�Kı;����Kı;���Mı,K�w�6��bX�'}}���X�%���ޚ�.�5r�Mfjk5���Kı;���Mı,K�w�6��bX�'}}���X��,c�Q�N��Mg�ɴ���oq�߯���t�:��Ծ�,K�����"X�%�����§"X�%������Kı;���Mı,K�v_8f��Ԇd�#9�����ٱ��SdM���v�w=�[t��Jkp�֭̔.���h�r%�bX�z�eMı,K�{~�ND�,K�{���NDȖ%�����iȖ%�bw����d]�ܐ�ǻ���oq�߿�o�iȖ%�bw/}���bX�'��m9ı,O�}���X�%�y�>�pܹXCVJ�=ߛ�oq���~��q,K�����"X�%����T�Kı;����Kİ~�r��)�j�.��k17ı,O��p�r%�bX�z�eMı,K�{~�ND�,K�{���Kı/8��@L�**�ER������e�ʛ�bX��Qc�����%�bX���ى��%�b}���ӑ,KĈ`�����p�:x��!�@��1}{��"���i ׬@���IM�$b|l#fT��1����!����!@v�h6��VlE�0�ޑ4���$
P5�A��b�@2$F���1�D��@#
�DgP~.`G/���x	���A�$$XB0�$~:�2#S�H�UbT��%
�aIZh��UN�.��#	.pBb�`"��l"@���� \AF)Uҩ}ʑ!5�@XD`�HD"E �C�$�$#/�N���Ξ�t�wowĲ��� 8�\�V���?�����
��<!Z;�΍mL�r<�P�]k�v��8���m�C�
k��Dp !�&����e�`��u婵�eY� Z�趋U�Ux�B��%;D�����������=o"��ʪ��cdH[m�9���"�c��Z8Ƶ��j��1�Vw�k�v\��������`�W �<��[��ꑫ:����{k�m�4�nɵ�����;-��k9ٚ��.-ݻNm(��Mh͆�6ULʯ[� i�|v�2&��X�Mqã'ݱ9`� C=�\�Q����Q cp�k&V���=,n�ym��`*��[v������Ҫ��e��m�n�^�cHJ�/ l�Yc"�M���R��%ϛk��: IT�/���q��9��|��u=M�K.v�C+�Ѯ��c�{p�wn��Դ˴����	�8�'.����q�N�d�×r5���w?2n��q�����r�m��%�Y���EƊ��m���n}�L��e� �	Ȥ��(�X!�p|��6���۵+���L`��y�>z5��Jk홢�+��S9]�Mi�{g�Łڷ���>�0].�W��!/nN+��^M�ݱ�W\����<q]��]CV�p����St�t���ãk��p�oc��=�q�Y�he��.�:��z;BJ����l	���m����WC7��ŭ�Th[q������k���i:(ݎ�]� ��8�c7��ϳ�-��4�rmy$�FY�,]&t�� �`K�ɳhU؉]��B{lhf�&m���qL���ʾxpɍ�x���]\�-Rp ��"��g$�L��:�nN-���CJS��.�U�]�uU��_5������*�g��Cˎa�#n`�m���]�j�i��m����dt؄M��Mjݭ�)ʖ���E���n��lF��g�Tdn�f��Wy��N�s�/1[\V�@H�ETq"�:"�#�b�v�D>0P xT?�!�$=M�	���M!�sF]�7��p�rm�T�(�6˭�l]��ѓ,u��N���X��;�8�9�-u�jE�sҧ�U�7$Oۄ�vz�c�Y��{jl�k���rY����46lu�ѧ����n���:�����1���sӢ�at�@+����=��5ùv�)�kѳ����x�Z^�df����[��Л8A�b�nڝ�����b5ױ�9�#~|�|�|��=�m�9� ���-��p݊S��We�ͷ9�^���Dld�.ń��lu�}=�{�K����iȖ%�bw/}���bX�'��m9ı,O�}���X��������q,&���>{�7�����^�17�DȖ'{��"X�%����ʛ�bX�'~׽v��oq������Y���+s2��ou�bX�{���Kı>��ʛ��Hԍgkv-���j�k&3fZ�,K����f\Ӭ�e�ֵu�ND�,K�_l���%�bw�{�iȖ%�bw/}���bX�'��m9=���ow����Ȼ5�����%�bX��^��r%�bX���f&�X�%����ND�,K�_l���7���{���~�w����������u���ؗ��B�%D�MI��8깪��ډ��55l֦k5v��bX�'r�ى��%�b}���ӑ,K����(~Vr&D�,Ow_�]�"X�%��k�ˣE�0��]]\�bn%�bX�{���4
�J�U>AO�tP�"r%��_l���%�b{���ӑ,K��^�17�TȖ'�=���Y2�.��j�Fӑ,K����eMı,K�k޻ND�,K�{���Kı>�}�iȖ%�b{���kZ�e�Թ�35���X�%�ߵ�]�"X�%�ܽ�bn%�bX�{���K��ȝ�p���%�b}�_ߴF2F���>{�7���{���O߮&�X�%����ND�,K�_l���%�bw�{�iȖ%�bzL/�}c�T&�3�e3��AF�n�֊����6�1J�n��g.a[����X�%����ND�,K�_l���%�bw�{�a�@g�2%�b{/�f&�X�%����s2�ui���֮��iȖ%�b}��7ı,N��z�9ı,N��q,K�����"~2�D�;���K�L�	��2�Z�7ı,Ow_�]�"X�%�ܽ�bn%�C�@S���5����"X�%����ʛ�bX�%�o�e�0��L�kS.kiȖ%�ʯ�	P���jƠj�k3��[_@�����*n%�`D?�"w��k��{�n�~�����8��w�n�"s��pI�,~��ʟ�X�%����ͧ"X�%�g{�i7ı.�~���c1CD�i�6�q��]�������&�u��yiĭw{�����&�WZ5u���Kı;���Sq,K���m9ı,O��ف�T���,K���ND�,K����ֵ,�5�sZ4fkEMı,K�ﹴ�? �șĳ���&�X�%�����"X�%��o�T�O�TȔk�Q�TTLTDL�M[_@�@�;���n%�bX�����K�$2&D��7ı,O�{�6��b]�7���~��,\³-^��op{�$�*��u[_@�@�lz�5q,K���m9ı7��
� � �&�:Q[s��MX�@�f��1J
�LB���֍�"X�%��o�T�Kİ����[�6��j�j��5cP5X�����Kı;۫}[�f�.,��l�Æ�f\/n+qVΰ�[�g���v�A1��{����>8��٭��7�̖%�b}���6��bX�%�w��n%�bX������ı;붡������cuLR%TMUMF��ND�,Kϻ�i7��T��j%��߿�m9ı,O~��*n%�bX��wٴ�OʎTȖ}��.�����u�sZ�n%�bX��p�r%�bX�v�eMı����>����ND�,K������bX�'�=�Kud�4h�Zѫ�6��bY�H���T�Kı>����ND�,Kϻ�i7İ?Ȟ�|m9ı�{���~5Yɫu�\{�oq���bs=�fӑ,K��G����kI�Kı?{���"X�%��o�T�Kı:*:�ٻ�{WVf��SY�/c0��ʇU+4q�3��β�[�G����D�D��h�����v��ݝ�#=p��m���mY�iZ�<%��9m,�b��q��B'E8ݷ7����=�t��!�s۝�\(�tZ�m��N+=��Yk5��O]�v�Y�h|�;�[���4�Ɋ��SӢNՁ.Gi�`c'��n�f�Su!]2��� �΁�����{��wr|�M��\8�ђ���qc�77�/n]s���{=�QoK��,e�jQ����X�&)EEL�UMOZѨ���}�MX�ı;�}�iȖ%�b}��?� _�j%�bw?�fӑ,K��?�n�aY��w��7���{�߾��?�9"X������X�%��~���r%�bX�}�kI��%�cߟ~��A���tE]�������d���*n%�bX��wٴ�K�dL�g}�ZMı,K���ND�,C{�ߧߎ+ �kr3Mǻ���o'3��m9ı,K>ﵤ�Kı;���ӑ,K�ȝ��¦�X�j����)�&�QT�UM���@�A�ʦ�j�j��w}�mtjı,O߯�ʛ�bX�'3��m9��{�����}��뜱t��l,��p��9䘬��.���7*�u���@��]��i���Xj�Z�Z֓�,K�����ӑ,K��o�T�Kı9���a�'�2%�bY�ߵ��Kı/|{���[2��\ԙ�ND�,K���Sp�<A� ?W�2%����ٴ�Kı,��kI��%�bw���#^i���KT5Y�M��Q�TD�*Y��Sq,K��fӑ,K��{٤�K���=�~��Kı=��eMı,K�j��Vh�f�[�5USSm|5PjbR'=ݚjƠjX���p�r%�bX���ʛ�bX-$k���m|5P5]�������%f�fkZ�k4��bX�'{�p�r%�bX1���9ı,O���ٴ�Kİo��i7ı,K����k��rLԼ]�1�`.%qý:�nĲ�!�Ѝ��%�N���<�>|A�%z�
�������%�b{��ʛ�bX�'3��m9ı,����NDȖ%��{��7���{����|�٭��7�ı,K��{6������MD�Pg�TՍ@�@����m|5P5;��7�eL�b}�~�e�0��L-��j�Y��Kı,����n%�bX��}�iȖ9�"� �?)��5޿�T�Kı;����r%�bY��~�]Wi�+^��oq����2'���ND�,K޿�T�Kı9���iȖ%����%�{��4�5P5Y�}�EI
`�
��	�V�"X�%���l���%�a�c�n��\���8���V5P5]�}�iȖ%�b_Y�j�a�ճ0�j�ǘ�\9m���ö*���"����;��3RՍ���\{�oq���������r%�bX7�{4��bX�'{�p�~@�DȖ%��_�*n%�c���c��3�f�4�3������Ń~��I�~AE�DȖ'���6��bX�'�l���%�bs=�fӑ?
 eL�bw?g�3F�]\�ֵ��i7ı,O{߸m9ı,N��eMı��,2&D�?~��ND�,K����n%�bX��}�˚.�2�5mֵ�֍�"X�~BD���7ı,O���ٴ�Kİo��i7İ>Ch	�:«9�f�[_@�@�r6�EQQ���T�5�&�X�%�����ND�,K��f�q,K��{�ND�,K���Sq,K��@����ua��ur�D��N��i��ˍWj���Vw��SB�
0U?��ϗ�K�i��������2X����i7ı,N����Kı;�f�����,K����m9=���n����ծx���M���X�%����6���c�2%��~͑7ı,O���ٴ�Kİo��iV5����j��7芒�TTI4Z6��bX�'��6D�Kı9���iȖ?�	��5Po���I��%�������j�j���S5TAPU5T�j�5cP5���k���m|5bX���٤�Kı;���ӑ,K��o�T�Kı9���3Y-�4j٬ֳY��r%�bX7�{4��bX��c�{����%�b{��ʛ�bX�'3��m9ı,N*;$�j�I�L��:�
T�j�%Mv]�w4��xݥ�|d�.��ߕ�|Ō��$�{\�n���[���=<����l��JtwV75Zv�N-�m��Ta�L��`�m!�J[q�䔤-�'��{g��3��v��]��96:�I��B��v�;qM�c-��.�uls�=����H�]���h���ۭ�s��l�q&$�4�&D�����aHNK�����uߟ����Ѯ�JK��k�ҷ��&n�+�7m�/���)�������>_>�&���k5��r%�bX�~���Kı;��7ı,Ng���~Q'�2%�`����Mı,K����˚.��4jֳۚZ6��bX�'{}����T�DȖ'�����r%�bX7��f�q,K��{�ND�,K��l�ՠ{5�)����{��7�����߯��bX����&�X�!�2'���6��bX�'�l���%�bs;��5����5���m9ĳ�@�9�߳I��%�b{���iȖ%�bw��*n%�`��E����f�ߛ�oq���?��v�s�A<]�7ı,N����Kİ� �޿�T�Kı>�߿fӑ,K��̚jƠj�k�>i�iPLAS�R^�Wvغ�P�6�JQ�.�*9��wnb��`���q�V�6�w������oCs�'�DL��� =8�~��H6�B ��F�"$�TrU����s�W�N$4�֚$��}636Ձ�fZ�o�F�����9q���v��j�4ךJg3޵`v=�M��gr	�I�Mm����޺�3;���w;W�}�`g���u*:N�D��9*��֡��WwW����@n�P�����lr�E��b���r�5�NGrT�+����7W'*Ժ]��|��:R�u��L���=�HN7H�j?��zCu�9��R�F��C�)����`n�P��֡�m��wAv\TL���D�\������"�#������	��C��Fl� |�a1��8H$R��o�bD":Q�1�d" �P� ��0>da	 �'FF1GFЁ@ �-K��"�R+�.7�*XLT$�D�R$��;XF�) A�����*b,���[��MrP @�d��@�	(H�1���"H@�T�XB#<��0�@I�1
T��eJ��mD�E�D������;� 
xL₺Du�E�`�GJb��-*/�Gh	�
�����W��5����[�[JStHSVw�� =-�@d�t��֪�>��ܐDD�rJ�J�>]���n��� 3P���ﵾ�U�UT�[h�9�P)uv�vܖ��D;��]��Wp�v�c�����ʚ�m4��m�O��@n�P��mG}�}����<�G ��A�$r;�޺�3;����;w;7��N�GIԨ�rG$ 3P���GDG�}3��Ԁ��E��o]
E)9
jG$�`|�y�8� =�� ���"!}�ߡ���NP��q�#�1gs�>��3����n�
��ɦ��q��JmH�Nz�srl��Gc^5�ٚR��n{Ll�Wf��IJ�*r���n�Ձ��u`|�y����Y�XԤ�I����� =;��8� =�� n��� ���IRIV�w�����`}��Vf�Հ}��ID�AHӎþ����7���@zw] =/yE#N�R�ے9���]X��V���nI������@�1U@�j/u$'��5ML�ԗZ��0l�ƫ��1�f� �L:!8�㳚��+������{\�f�0�vS;��Wh�-�Q��m4��{g���[�\M��#-�#�O(��x�k#�1!�]9�T���ݗ�1ú5Zn���ϓ�mL�/<�n�p�r����ݴ�Y��t�}")�ugV��Q��t��L�N�W]��f�v9[a������#�p߾��wws�����|?9n��Jۗ/fr��ίX8���ܸ�ջC�ӫ��q/b&�[#�O]����0�(@zw] 2q�@{u�@}��B�AJNB���%X-�vN7Hn��� =��WL�PIWWwt�����֡�ڄ�u�5�5��N�����v۽u`f6���t������5S7P]��Յ��1��S}^g{���u`u,��ԏ�M�!��E%�S�e�V�a��^�]\�Jt���-M�61CfYrJ�J�>[��Y���z��_ ����=���Tn���`b���J��0h������f��������v�%(�*�#���Z�cj�D�K}H��n��:�'R�I��a�z�=���K}H�ٰD�u�ϔM�ՓQ5!MH䒬��;w;�޺�3;���5%ʙQ4HӨڂM�?˰�˶nƸwb^�]���l'm�8�*�\?]����l�I:#�9$x.��v۽u`fw]{��߾A�����~�Q�L��r����j��@zw] 2q�]#����)�$c��w޺�>[��6�@���Z*u?"8��;7޺�>��m�""B9*Tr�������7Z������z{����(�7RE#�1gs�=���o�w�Bӭ��Q;�I����ŝ��JK��nu�'"N[���]G�a�A�G�!c�E#N�R�ے9���u`s���������i.Hdg�6w}déQ�u*$���Vgu���~�H���5o�������
RrԕwwN�H�n��}��L�|���j��;�U@�%(�jj����6��mNV{�`f�X�e��J�lHi�,mKm:��ɰ>�k ��&�Q0��ET��rՁ�&�{���Fń�;��Ԍ�PR'"��m�D7O��6u���V�A;�&�.�u�ݱ<4�V�����=Z�)MQ*1���w޺�>[��Y�����޶Ӕ�R������~M���I��ɑ�����V9�j���MD7v�bj���L����@l�u 3u�@f6�����{�)�JT#rG#��~���~�[����wmXGs&�Zi&��ٰ9��L�*:N�D��9*��?��{��5o����W��Ut�V�~k����x�h�3a�n�,�Tf�$��!�X��]a�]��h��\k��֞���5UqYrl�n����PӴ�W;MO���n�n�N��X�l㛑��G]�vvh���:��W3`����.�'F���u�.�R� 2m\��3yΎ���.�-�x�e����ZVm\�N��<s��[;����v�e���dfv��H��V�n����w���߇�k4�陸ܦ]��(�n�n�p�[���{tݥ�������W��]�%#��r�I+�<����ŝ���޺�3;����"H�'QJ�&��jlG3&�i�4�s&n�Ձ���u`|��߿W������)НD�97t���B1�N�H�n�]�$R�E*�I���a�7�����f���fM���I�n�����f&�DHG%J�J�>[��Y����3�����U��/�R�RdmTm(����ٻa�\^��5���QoK�x.�j����ω�#�p��I� ������޺�3���ד\��o�6c=⢨��b�3USU6;ܵ|n�Km��ݤ�˵`b��`|��߿$gw�m����D�]�]�u��[�~����@k|��o]%#�%9
�G�a�K{�����@f�P����ބK���j.n&J�������o�u��{���N��F2SIȇ�
	����p��V����͇��Lt7n=�������&��r�����Vf�Ձ���`|���[�]5(�R��9*��޺�=:� =8� 3u�@{u�*��*j�*��`}̛��d�)4�i�4$&�r��3�V��Z��2�jj(�
�ԑH��w;7z���޺��UR���5o�F�8�Pm����B3Z��[����؁�D��I�ٮ�!���cQfj�srۓ�N��4h]EVn�h����Bӭ�Ӎ�7Z��jq�JT�TR8�����1o����Ձ��u`|��D!:��9*������B3Z��[��g(�cBuT�E#�3w����$�｛��s@De���< u���M�9�s`g�Z��(T�I&�j���w-XM��\�ݟ��wvlwz��7��~ 	ҕ*S��(���#��cخ�8MƠ՘�z�yI�C�DT�a��MqqwwN�HN7H�j?zCu��o��NDJp��7$v�;���5�P��|����~��&M��&j�ꚕܑ����Ձ��ug���T�.����}�`}��6Ԩ�8$�J��I%�o���f��G3&��$�w3�U���]$㨔�"��rIV�{�����7Z�cj���g�@8��S���� �a��'�#�Gf(q�u!!$�!��1 Ē��D�@�B饬M28 �!��c�*�  �� `�1�BDFE�>%b�!FB0KhT:VAbAXD�֝ O!����"���	��G�$���� �`���O@��`֮�p�< ����!��(D�2�M�w�ֵ�UP+���V7!�۴t
�@bljV6:��c:4:��M��˒����%@��]�N�#�DYv˜�����*t��c���9Ӣޖ[u`l�KmUn����m,BJ��:�L5��C�yyƺ��).�:UU�³/����I�]T��gnz�k9��6��F��<�J�`�ܔ�
���u�V�afR�b�n�L�@WJ�����м��ËW[q�{�v�'�lV�8:[iZ^��H��V�H݌9ťPU�u[�j�y��@�T�s��,D�6đ4����!���*���=:ݍ����-�au�tJPU3�[h`X)Ih	Y�N[���3�l�v�t�!��e�V���!m�*e-��E(t���]��Q���I��a;]��mK+���[�i�r�zy���1��#�i,[.s��ۭ�3�u��q�)õc���/�xŀM�������'��K�&λι�������q�ݳ�	n�����ݷl���6�"6zn��qf��ے���cY�n-�;Sd�u�xzò��
��P̥��d
����<��v�K�1��l��Wi��c��%��u�2ოq��n���M�Z��ҡ�@��gg�_7f8������ƣ=`�&���j-qv���@�� leՃ�#��e��3����,shq��+���{�^�l�S���*=y��g<�q�6��lδ�u��I�tX�fv��	[�	Y{]��q˭���Cf�/l��v�{6E�kf�n��6��k����=����0l�9�����X�8��E�DU�gHf�Y9�No@틮uU���Cpl��52�dy�eV(��uU�6҂K�
.�Wq���ˎƘ`OMq�9fz�]�	V7#�DZ��N��$i�U�ûs@m1��0pt�Q�r�(���[[U����FF����D��Jl���u���  Щѿ'B ? ��"�Gi�Q��46�����{�/����Mi/
T��ֺ��u�v:���Ѵ���:�s@�]&"7].5!sf6��ga�{!���n����`�k��5�Q���[`�]�i��Im�w;���TDn�-��6�c<l��Sv6.�9]�<;փ]5��.�-�3�7Xt[�vJӬ���8�"xz�����b��AΞ�q�����R�40(M��n��=��=�����q��H��0u�����<��r֛���ש��Ӂ������_Q�=��g���H�j����#�/����E#�n���vn�Ձ��j��;�6#��~m��S&��)�Tc%X���V�{���;����u`}�ք�ARp�J��a�ߪ"r�u 6w���� ��'w�Ѐp��ѧ"%8Rn��;w;7z���>[����!7Q�dc��p�ۮ�a|u��Җ��W��u�pK�4`�u~���':jTrG#���Ձ��u`|������oC�R���"Jj�j���fZ��K�餒Cj5�Pvo��;�H�j舙�\L��C�TR9$�{��ŝ����Iow���z���or$�Bu���;'�n��� �r�u 7i�s%'BpMӕ���޺�=�w���{��ŝ�����F�h�ҩR4�OFm�غ4����eS,���:]=4NYڥ��S�R�N�������ř���IyrC7}j���&��UT����� =:� 2q�@f�P��mB�H�[��ӑ�)7MI��}�`g{훞J�AJ���E��I9���bn�yj��w�6���"h*T�*&f���l<�o�Nn���������;w;��sjTt�DI;���@f6��O����R7Z�m�����&8T������6���[����Rp��)�NT�t�����S%��7r����x��H�n���~��r�.����J��`b��~��o� 7{� =:�/��&�>.��*�f�*����(@f6�9/��[�;t���(�R��ԕ`g3-X��M���d�	��4�M�)	#`���I�/�=Q����'=�l�4d��Z�a�Y��ηH�n��P��mB�������~VU ����\T]vN7!�3����j.	h�e}q%;7���?�v��EM�� ���Hm�@f6������n":jTrG#�3��������7{� ��@d�t���T�]ETDI9����V�;?�վ�7��Հvk䓓��FTR9$�V�R'�6� 3P���䛲d�)Jhq��1gs�3���wzX��M�M��6��G��*���
�Un=��4f�k�Spr��Tf:Wmƶ'Jb#f�s��QZ�v�v���8�dSsj�6w*�Wm��6����kp����a�Nך�f�Wv6�gL����t���ݹ� �N֚�`gh�ɉ��Ɏ:/O�c&ͥ�FȻmB���.��]2�s�f�0E�D�0k�n1��q4�6h�� �����4 ?k��.Y4d��0��3Y� �[�1�l��Ōq�qU9��1twfl�t��J:r���{�u`���ս����\��{ޛwOM�2)T�&�1T���U�4�A���`r7vlfe��k�F{޺I�i$�7@RK�{���gs�~K{�@��`�4�:LCq3U6>�n��� �v����`b��75*	�����VD}�����HN7H�êQgN+���f�E:z�ۛ{�3�=;Z�ht�:��7�"�Jj��B2D���*�37����d�G3'ɴ��MrC=�Z�fϢ"j�*�EQT�����w2o�����S'#����� �;�~Kɤ�ɱ�� ��DcN9v���vwuՀfoKV�;�{ĎP������þ���{�Ѐ7_Zg[�����4�S�Q5NIV��,UW��sv~��ٰ9���q�㘪�)��^��gb����ڴ��L	y��^4�3�$��b�r(�'*$���uI,[��N7Hm��">���/����
SD*"����9�7�QwvՀw��`v;�7����Nd��x����LR�&j�j���{֬��U��li4�C���� �8�k~��ٹ&��v���9N�D���*�������}h/���n��P�m2T��Ԍ������v����X������3zXn��Tʈn1�Y�=���A��q!���K�벊t�[����١�G#�B��8�q�-�����j�9��y6��#7f��g4��D��DB���jlfe��I���ͫ#7f��9�7����M��wOM�̐�R������}��:� =8� 1������(��5R!I,=_���Ͻ�`r;�632Ն%�Г����	��������k�r��35%��52�*�l���`kM4���/�����[������JJ���#)2`���ͮ����of퉱:��!�n��#��N��M�*
9����Vf�Ձ���������ٰ9�F��QEMAQ7uwp��֡���Ӎ�j�I4��M�2͟UR��ET��$O~�HN7H��L�w(@n�P��}�R
���8�q�~�����K���ܡ��B�G�D�}Ԁͧ�7V��"M3S`s3-X�iy&�y��.����G3&��k�I	!&(Q߈M��	���M\��3F�����v3��1i곣��7)�6.�G��98�'^Mg�s.ˑ���������&��Rd����v�x��ݶiCuXݛ�������zc��m�ŝ���������;tΛ���b7&s�C��]K�θշ�7dz;\�êm=�i����^�ɮ5cq��u��qoq7Xԧ3aj����������{޿�������#CD�G��Τ�u��%��d���7gՕ�`�ӉZ-+�z�Nl�q�=����Ӎ�菾����ʬ�^�۔�JD�ID��[�����r;�6wvՁ�w-_�M8���&��iJq&�)#�1o����3z���os�1grnF�iJ�nH�vn��j�n�tG���Ԁ��=I�R'NI$�3z��Ž���gs�3{����)4�:����3��њPF6K�I-��ӄ��ZH�Sߪ�
[���(�%QH㒾W{����t��mB3Z�m7D���7uW.\�kY�ܓ��{7�B�U�D��HE\
�WS˭����^ڰ;��V#��~M��vs�'*:#�*N���z���޺���U%���1o���9�F�R�j��+��Z�9�6��ɰ�I'�?{��*�����܂$mT�9*������}�����P��֡�z�˵��'�O�]�v��vR�\!չ-�*ǛqL%���{���m���x���Ԁ�mB3Z�Kn�8�rF�h�ܑ�������������]X��������`}�C�$dJ&���X�rՁ��ɳ��!!bD'�����<G����<�`� DXtT9��`���-��A{�a�_a�eL�!��,��bQ1����/�SF��@��%�$V,`�&�
��^�4�m!Ë�ȀV ��'ʮU�,�+S9��
Eă b$>P<�)�uW��@� �U<
��� t >Tx*|�t5��#S~vٽu`��'"
#�TR8�+6�o�)���6c=�;��V9�u`f��')P�M6ӎ)����`y4��{�� ��Z�9�6c�N��g3Û[6u���-�a�ַnu�s$5�[��f�a����p�Y��j�� 2[u�DzC'{���w�R�j�	%X��V˻�����`n�]_��$n����#j��Wp����@zq�@n�P��֡w�X � � �;�%�f�ˬ��ssZ͈<�������߳b �`�`�`��{��<����{��6 �66
8�|DQ����]'�=����y=�~�����4���w{�w��n������6 �666=�p؃� � � � ���~͈<������߳b �`�`�`��"������ۘMkIK'�3!G�.`˴m���,�9��ݺb���w����4[p�}����A�A�A�A��p؃� � � � ���~͈<������߳b �`�`�`��{��<������~֦kVI5��˭f�Z6 �666?g�߳b"`�`�`��w��؃� � � � ����b �`�`�`�����<��� �r9����K�)n��s2�WZ͈<����s��ٱ�A�A�A�A�����A�F�����y���ٱ�A�A�A�A�f��Z��XK������f�A���X�d~����A�A�A�A��p؃� � � � ���~͈<���-���߳b �`�`�`��z~��C�LԚ֍�<����{��6 �666( 1W����͈?A�������؃� � � � ����b �`�`�`����&�*��{o����V�鵗����P�54rC�-t::s��l�!���k�H�7/�$������D�`iknw*�!mֆ��[��vD��C��B�ӧb8�7N�����b3j��xn���rZ�����63آ��>6�5�|;�ֱϐ�Ÿ��$�D1jCO\�&�MЙ6|��/ƪg+�Sy�F�T�K3Re��#�ؠ<�&sR�#�������5a-q�{WQ����,�O^�)<�萇���}�%��}���lll~��f�A������ٱ�A�A�A�A�����A������yg�e��ԙ�����%�k6 �666?g~͈<�������6 �666=�p؃� � � � ����6 ���� �l}�������̳F��kY��lA�lll}����<����{��6 �6 � ��A�~��͈<����s��ٱ�A�A�A�4�3l5M*�SRTDMUMR��	�� ؠ�=�p؃� � � � ����6 �666?g~͈<����}��6 �6667�}�Z��Y$�j�.���h؃� � � � ����6 �666���߳b �`�`�`��{��<����{��6 �66w����������ֺ4\��/:c��ۜ<��ֺ��-�s�ѽOmv*h&p�pVL̷5��k6 �666?g~͈<����}��6 �I��N���X�ݛ�Or�&��DUDI553S`s��W�&��6��j��"� $����lܓ׾����gs�3t�����IVgr���H�""gg{� ��͖��4H��(rU����y���v��j�Ͷ���X��h*�&jfeWt�����ޏ�ܡ�mՁ����&�F���T���u;�|u���0���e�:���n�0�P����"��f�l��j��3-XFfO�m��5o���@�%E)�D��9*����m�'��������}jG �*jG$�`b���Y��T�i�
;���̵`}�̒&�(��*�f��n�};[�H�� 3J�ɦҎ��́��mTMIT����jj����B��>�w���2{��8�X�߫<u����Q�R����B��b�nD6�H�����0���9��wj:��`���������M��TMS�$�������ws�1gs�7w���K�9"CR6�J�`}�7����;ݛ36Ձ�fZ�5��~H��iz��j4�$�v������-Y�n#�ݵ`r7vl���*��m������u`fw]X.�{���b��"�P�|�U~��U������`y��)�D��9p��mB��D}]�^g{���B��{�������6W<g�ƨ�s�vz�v�#(�콌�h:���G���ɥ��(9*���pǽ�9̛��Z�m���w]X����r��m��G`d�t��֡�ڄ��K>����*�Oy��鶩6�p��Ձ����u�Y���9�F�A*&���R1�Kn�8� 舉m�� ��~i�7�%J�>]��Y���j��@(��"5�e�����ڲ��i.��y�׍�^Od^y-�ʛ�=GV-ۯ=Zs�L�t�ɯ#��$���� r���U�=:&�e����3����J��Iu��e��2]��.�����
��>�E`���-� D
�/��N���x3c����nۇ���z���-��Y��M�x����nȽ��m�r]�����W!t��b�j�����ϝ� �G>r'aYQ�w��b�ú����m۩:1%;�����R9�MFۡ9˻���޺�37���w;w6Gm������B3Z���HN7K�>���7�<�D��"I��`n����w;?�~�K�����]X�ϜnD�*jT�U+m��J{^�����zl��j��>���r�JH4��G`d�t��֡�ڄ��H3t	�Ξ�Ӟ��'6���0����A�"Bf8f:z�v.�6�������(��L�Uu�|��ڄ��H�n��.���TJ�c�$�3�����W_�i�	��$���wfE�́���`ww��ݍ�NH��JT�I*��ws@zq�@n�P��֡����V��TL�"j��ʹ��M�k=�7w֬������ŝ͑ěD�(�n�l��j��i7��o3}��;����gs�;yu6�%�4S���ME�o�]���#�GSW;�7�D�%�����)'$rU���u`|���,�v��Հgk䓔�R%MH㒬�����DDɓ�Ԁ��B1�m7I9C�$hq��1gs�3w�����WP�E� �1A��^*��<���>�5�훒b���`�ВA&�"c�7�����@n�(@zu�@d�t���Z����R�$�
�V9�j���O�4�k}��]������#7�B���U`��&P��^��3n`��5׎ܼ�I*����i�&D�IC����;wR7Z����Hn�(@9�S�U�M��M�RG`b�����7��������Y�������^�:�ƣD�(�nF�m�(@f6���������@l�u >·'INS���8�X��V.fM���d�q��Ba		KBMBi'm%�&��Y��`ݝ���@�E5#�J�1gs�1gs�7w�Ձ��u`�G&��A�M�9)5�r;����.x��]mr�C�n��9���2����GJJ�hq�#�[�;wy�X��_�U��A�}�`{�"pI:�&8�wH�t���B'����L��/]DЩH$�G*���]X���,�v��7v7�I#�N
*�UR��i�g��`r;�6{ܛVO���}V�����c�7I9������� 35�@d�t�P{#�}B|N��B����А��Q��C%Pb%b�%Tb�! ���\�$B@��D�8�S���`Ў�lx�R�p�>R�Ҕa���1�����k�ap�䙄#&JhF�R�I��hȰ��DiA�B,5��"C���, 	��ʔ! ��s 1 DG �!U�$ ŁP Q � 5�P�w.�+��T&�06��J�F#a�(1���%>kZp[xҷ8෵�m�Ceɬ�섶��&�V��v�nVz3�SR�&;mm���\l�y�s��ί-	��[N	����]�@j��k�b�A!�v��mn�:a��2�S�^�|��[<������iUU��3c������	GF��6�!;sv	9D�q:a3Lb�^GN�qK�]0g���v�,#��q����.���6U�9#H,z�tg��h��ۖ�p�����^P���^V�(�\�&f2eb�5���UI���-T�J�Rӝ�wh����e�H�<�;-P@����T,Ξ�g���`^u�[n:P�V����[���jX(	Y�N[��͍�Ƌ[���*m��e��Z��m��r���m�m���;);�l�]e���vWM�<�0����&Jt�F����m;�.�T�k;��3�¼d�Nb&,�����󜽭��s�Vzv�'>�H��zm�Ng��&��b��MvVugIkӺ�m)ո�:u�������%�.5�n�b�Ǩ�'C\n�gH��̝!�E����g�Eʳ⋚�e��N*P��HlKv�Bݭ/.���ptq��ճ<=��v����ķ/ce�c�J���]���gn�%Ι���*n�s��F�k>�x�)�3�9�JW[��*.�n�r'dݪ.��z�Y�[�E�����W!�9n�J^!�09��ˌmܖ��=��u��3N[� �u�i*�92m�� 'Z�d�c;�w�8�r<YVkI���m�Yk[Utp��$&���mÉ/,�v�+d��Ү�ݤ���+��9��t+ڽ����fiɱs-ܘlJ���
�)٪������HC[n�R-�e� <��5�q�X�۶�P!��LP��YK���qIӘVv���u���B���,�ٖ!vW��N�Ʈ���m���V�pm��QE ���.��b��љ��Z�<���m��p� qB������A? �S��(��P=��~~T��IN�ɒ�8u��L�	9��շ6�6�v��3Z���y�EC9�ٶ4��m�p<�πv�G�4��۵���pq�u�g��"pLٱxs�Gv�"oH����U�����k��m�@�u�(}qWd��<S����ݵ��Vǝc3�zá�,��w%�V��=�5��#��QG�T�mf�v��{3]N�r�6�bٗ1��&�2�R(�TMI���I�3:�J7&L��ٚ���Ct�ٻblN�qY;6�Xz	�)�4,'V67�O�����w-X�fO��i�C�����Pzi��9I9#�U���u`b��`b��`n�;��A��D7�8�jG$�����@d�t���J��@c�擔:RTm$�Ga�U_�������6�s2Շ�q����M�*&���R&8�q������1gs�1gs�9�]qpt�cT��G�)��S����on8�q\>�����KW��P_:#PMӁ#����Ձ�;���;��ꪯ� ��;���~jI*pR���VI���͞6'x ;D������;�����ꪤ�-��7
S�GS5wH���P��mB'�˷�H�R"B�r7#�7w�Ձ��B'�G�9[�Hް����)'$qʰ37��Y���w;{ܛV�m����h�J�PTUMEq�L�tf�Q�p��.j	���:�:Z�YcmO׽��n�nqԎ9+ ������gs�7w�Ձ��u`g=擔:RR�I�\��Ӎ�w](@fkP����w���$�Iq����>��ٹ�,��h������`j��`en���)�89H?DD};��w���n�t}���X�w��GJ��J��%Xgt�>Y����u`fo]X���R�Ԑ��@j��ۆ��򵬮μ��a;`�3�"E��n�����;����� 35���H�ր���uu7rHR�F�v��U~����Հn����gs�>΁� pr�����*��;���̫5��q��́��6�;_$�
�)�rU��;�����ܓ��f�� pT>D|��Gٛ��Ǽ�r�JJQ�8��,�v�P��mB'�ˍ�s1W�p��f�����-��^�nn��<2<���ϱF�!jBG��"c�7������w;�����'JJ�	������f����g{���Ԁ��wW����;Z�8�P�T�I*����@zq�GG��D�o�Bu�,�̒RDc�GI9����`n�M���Z�֚q�����͉U%D�dM��U� 7u҄G�n��x����ɰ)4���F`�f�15�ږ�f��3�R�M�oN��SNTn��	ll3�sl�]7nnُ8��cm�m��L�
v��ٳK�ŕp^3�kF๸ݱqY��N�<V�M<sٳ�V���v��0�G��a۲���gB\w�����G/n���=���WiΉ���s�������we͍v�!�Tx㹳��۰���[&�z�rՖGr�T���#H6���z�xg�QKn�8U�+�%���K�Z�v[u�v�y��3
�1��qD�]�]\h��8� =8� 7u�� ��ɷ�8Ԏ9*�ŝ����t���J�� 1ֺ����j
1'R;�����wVf�Ձ�;��}�x��*u$Lq��7w�B3Z�N7HN7H���]��A7N�U���u`~��~�?�ž�3w�Ձ�l�R��$����H�a(9��1��e	��wcud�O^O,s�c�$WALrH�r�*J$�`b��`|�������������y��JH��q�ֳrN_����H���LDhټ���o;o'Q8���������=��%���`b�y�o@�:RQ)'$qʰ35�@d�t���t���J=�5U`�&�LUMMR�9ܛ[o������37����oGD
BSL�/:�0Ztv�"�N�����6�:�7H�fk2NP�:�!'�;�����wVf�Ձ����}�x���	"c�7t���J}��}2n�P���Ԁ��t�����*$t�H�X��V_wٹ�`��Q�� ��׾�������z��䎇(r��IV�Gӵϩ��Ԁ��J�� ���Jh��q���,�vn�37��]��͝Q!E�P%5�.�θ�c!��vr�nVb�Rĺ#�Yb�Ŗ˞���]˴�J)(p����{���j/] =8� =����T]\L����*��޺��~�͇���}�`f�?��|�p(�MH㒬��Ԁ��t���J�� 1ֺ��Q*h��"jj���So���zl��ڲO��nO/��3�0QS�orw��35򑒓	"c�7������ 2^�@zq�@~���/�n�_J:�ˬs�n��V�s��f����#s\K���b/*Zg�������4��.ݒ}�B%���n�P�ܭ|�rGMJNT�I*������gs�3w�Ձ��u~�ߒ<���RSQ��n�;�H�t���B%�.�nSp��
Q�܎���wVgrՁ����km8��vlfѳ5!
�R���8�X��V.�v,�vn�>�՚�E�m'U$n�M�7#�9��ʗ;k5q���XM�y�ڵ��up�q[['$�HQ�X��;T��Xu����;%�����ձ��F�|[n�jp�M��ٲI��䳯d�I�q�O c�m�H�72���V������d���K����m����}E�s�)�,�Er��Q1����y��v��[u[�3#f�������
|Q&(�����=������e���^��K�[x�g��v�M�)����8[[�'*X۷���o�fm��4SSUT�#��9̛��M��M4�����c�������nRt�bN9�'�n�P��mB%���(��Iq����u`fw]Y��m/4ڙ���l�������`T��A7N�U���u`b��`b��`f�;�q��#�:jRr���V#;�`y���m,����f�Ձ�fZ�;��JR����:e	���IOVw��	�Wp��dt��/F�٣CE�X�䌳uPM��'�n�P��mB%�v˷����r7#�3w����`��j���:"���oB~[s���ڰ9ݛ��ɿ&�Q3h�q���)I9#�U���]X�y��ߛiDv;�6s6mX3��3T�TMH���%XW�����[�;wy�X��Vs�i�I�pR�qH�Yΐ�-B1�N7H3t&Y10g���F��(�\� ��Aۮ3�'Q�1�ל�괹����,��K�<T9�g�6� 3P���t��������0TJ��p"�������ŝ�����W�ߪ�;_?8��SR��T��V#��`r9�6J>�	��0��L]A����GF�̅�Q�4������gC�(����@��A�:`jRձ�+l��9��B�%RQd�٦P�!B@�ۈ��n�����a�;LqL@AV�IHD�!����c,!
F�(K��.�.�"��՗�i��vM|�z0�9Msꒄ���(J��;��ee�T�%ն[IX��Tq�ll((k3�5��I�AJ��)"0#����������+��@�UC��@"�PO�� S�UP����)�@���٫�7z��>���Ԥ�q�)wt������� 3P�����+{������t8R�F�v�3P���t�����興�}=^�;\��"n�z���J���wZ�K�L����=nܺ��v,d����:�5;�!��ڰ>�fM���d�6�_@fdm� �w�jJ(��SR9$����ŝ�����VguՁ�=曔�jGD��UM���d��c-Y��҈�wmX��v���l�t���8�v߿~n327�`w������a�Sm����x�>Ϯl�Wk�!�&�TU+�̵`j�m��Y�O ��zl����6�x�������<��0�tP�3]v�[��uJ�3�s]yyڒ5�)cc#pr�T�9*��gs�1gs�7uuՁ��u`gu'%	�nF�I���;�����i$�MݏZ�3=�V��ɰ>]��(�N��(�nG`n��3�������,[�;V��������J"j�b�Xy&ӎ�w�`r;�6#��`n��;z�N:���rIV����������� >��>U�H
��箦s&MY�M�]nˀH�#��Ƭ��g��yNF���u����c�-�汮rWu�<��mj��"���9�ê���[���ӛ�\%��Dq�����Gis��#����9���w<V��y�v�c�t�s�,�����s�<��=S��n�۹) ��=h�����2�z�Ӯ5+��Ns��k��2�Y�oo��
��Ut��9r�[��3=�����������o�|��e��	����%�ώƸ��Zi��<Wn��W:cK���n4�48��]�v�37����_�W�1o��9{Ѝ9N��1�����j�� =8� =8� 266�F
�Q5NRU���u`|����ߪ�ž�;�z���n�I%DJ��.�>��r���;�Hݖ���u`gNJcq�����,�v�#�m�z<��N7H�D�7h��v��dج�Nf�4y��ۓ]����ӻ6�h��hi�7a�KOͷ���P��֡�����2w��{���٬.��nkZ˭�}�}�t�D !�kI��K�;{6cwf��{u`goZ�BN�)�rU����`zq�G��"e�<���Bε�����MTTL�SQU6�my$絞�����������>��QF�JRDʺ�����P��֡��������V�tT!�1��m���u �-Κ|xG�/!�:勵��ݰYhĵw�u�ϛN�j�QV7q�7_(@zq�@zq���ސo���[�q9$�R�*J$�`|��ަ�Q#��`fdm���Z�i%�ܰ��?��Dm7n	����������74�A� �(�`1
#E?��Z��u`j�y��y�JA:N��������������gs�7;�(�#�)�I�������{�?�����c-XMr{��F��Ɇ�'x@�f��.e�kM%5���q�`
��5Lm���L�~��Ԁ��t���j�� <�]�ș������}�������;�v�ǭX��Vr{�~M5��U3U)Iq���/]X��Vc�V�;��յ��0TH&���J����iy6�3}�`{'}��ɰ���IA"�H�Z5WPGz4 ���ݦ�i}q�V�Gs&�j����M��w��P�������yB3z����V�HM�1�Fʉ ������L��u����	��cQ	dH��{��]��M�ۀ���1o���]u`fo]X�yX�y�))8"8ۑ��Z�f���P�n����բ:R�����*��;����R^I�3�����Z�9������D��RR9$���+w;;W]XW��w�����5M��48�qX�fM��4��Y�qp�zՁ���Y"&� H��@/�dD{��o���۩J؎݆���0��'�5gF�G����%��U�Z�v+�"�]h#i3�d"�lީ^4������Cx9ώ7T�8*�b�#����@�:��g�nFx�v�G+�2��`��Y2%6
W� z�lsٹ-��&G���Y�cj��p8g�9�U½3u��晛;	$��]snq��[nJ]��߃�|S���Z�7`�k�S;, �{�������+��rsr�p��ڙU��v[iRTR�nn�U�;/R�s�Q���7D��P�e��o���B1���G��zCg{��㧂0TH&���J�3;����Hž�5o���]u`|�y����*\wN7H�n����� ήD�H�q��ܑ������Ձ��u`|����y�))8"������j�n��n�m�~�����D��i9G5t:��z�J,�J2U������3;&ih�t�s)'$�`fo]X-�v�;�����z���w�	Ĩlq���9*��w2o6�iJNNGo&�����Z�����$g��Ґln(�C�)��}�@n��#��;�� 2_u l�S��$���8�v�K��}V�z���w2l5$�r{�6V,�
��U2����@fkP���t���t��5�@jm$�L�UR���AE(&]�,�ɞ�e�e݄�(��m�[��ٺ��~���|�.��*J$��j���>Y���z�+��* vur$�F��7���f́�f�@<֡���t}�ɳϪ�R
S�q�#�;��Ձ��ug~+�@��"��M
��Gq)|��w;s��n2:R����uJ��;�����`}̛&�O�$��{�*���[�P鸊JG�`|��@~�������� 35�@�����kk\���hc��8�&L���|��o#�cu=�D����S�˖$L�S�N7Hݖ���B �7h����IG�n;wW]_�����޵`��XG3&��N ��9�T�"������@n�P�=��Ӎ�wW]X۽$rJ��Dd�I*����ߒ�wj��wvl����=�hI$ "#�=U������Ȓ�n4����gs�7uuՁ��u`gt�3vuD��C�M�M�f��`uñ��n�k"\�=t*����G-8BrG#�G���#�������;���fV���I.Hv3ޛs޸��#�)�I����� �;�����`n���g4�He%#�\ cv���t�����������1H:mĚlrE$�>Y���]u`fo]X��,���GND�Q�M��] 7vZ�f��ݠ=8�nIҩ����M��8�tH!�(�"��!U~C�$2A*�@���(JbF��0"`B��BY�F�dc,X��,�����R�B�$*����
1���>F��1�aXH�XѓF$*��b��ҁQ!Er�I#������"0��F�$ AHB��B"� �D�$�HO	�bA���v�!�/������N����-��m��T����	FQ�ɭ�/l�l�h�"x�y��Ljձ�Z�� �k�һ	�]�9���H�U���k�H�X�ܖ�u�kX˦ie[E�	�u�2�vx�!hKh�C�v+���Fd��v���U�Y\�`��v��v��y+4:$�EZɇ)`���`W)�����>:�#���di͙�<YG#���g��,#�=���2���a�$���q�h6�n;s�:m*z��]�Pp�֡��:ڜ��ۍ�[]QF��U%V�-Tc@T�[�k<Q����d͚�첂5��x���
�ʝ,�]��y]���'�cu�ڐ'm~���N�I��X*��%ge��u�iW�9#�!�M�:)6��`�j�������q;m5+�e�8��6��0A���+Ƹ���T$����5rOA�����|����t��n2���l��H�t���j�9]�[��7��j�>�q��n8(��nB%�x�X�9"��y��'=�kY�L�,�K���	m�"1�8�v�O�<�D��1�<�t&�[�j�H�6^!��l���võ��p��T���F'=X�P��Zta�Օ�|��]�=`��@j܏%�u��<]K8�ٺEv�Du9�U�>	��kn�[��F�/��6d9¢�d�su��k0�Jq�1l�-T��+��`+�৙͇ ���lj�U�U�9�Ca|�r���������=���um�K������:QM'Lk$�3V���i m�:2�ݭA��V���V�C�$6�um�t�UK��c@	8�PڣA�	�u�]d�,�{�Z�<Rc��ȵSP]b+��t�������WZG��M��
�.vFۖb	�ڔ�I�@Mӊ2c!���٧�|m�Y( 7+-P,"��b��,�M[af�6����ٽ77]Xd���R�̂ݸ�^�Z�����v�[�[F�\��R� ���܊��\�~��������
�^�� ���\ �G�T?/�%��./S���}�����v���t�͋�^D"�����Z���2D׎�n��D���Kv$%v�t��u���3u��B^X%T-�+f;V�.����r���jïk=v������uۇ�Tl�<v�cd�m���N˺s��6��?�����<8c�ݜ�$nrū��,.�qŷV�� �@��������.nɺk� q��[�jr�4�@�z:5tH7Xm�{���{�Û�(���v�����unn�Vwc0u���Gh���v9�j*l��������}cIz��"�����P�=��Ӎ�we�@���qӀ茒�%X��,�w;��e���Z�ē�I)��G�R*��#���KW;t޺����ߪ���]Xw�,]��rA��ܑ���t���B �n�~������@=��F�#D�))$qʰ37���߫�N�u����P�{R��7Q5{b��5ͺ�8ٷ���8�g��q�W[�Ɨ��|V���q lQ���9+��zX,�v��37������:M�$�TUU��s2o���I'-��&�����z��ڰ7}���̫�q���j
4�Q�Q��;�����޺���`|���[OyЩH&����V��m79��+ �����9�6m8�͟��s3jjf�M���"���f7hN7H�t���B��]����s�4�ĺC�[�Z�i�q�L�#����n��qR�+���&�`}̛��M���ZԚKͤ�$���`r����R�B7$r;wy�/�DDɺ�Bg{�����ڛ��F��B�G�3z��ŝ�����qx1@+"DFʰv�j�I}\��͛Vs����@T�2���%XUW�}�`b�y������޺�3�s��6D�c�)%��s2l$�o36~_��ڰs2�6���ݏ�Z��zslw%�g7 ��҂�\F�:Gd��ל��s�q3�K:����� ��P��֡ f7hN6������T�t�H�X��W�_D�n�Z'{���� f��������9V��,�w;?��]��u`n���3�8�)����K�ӎOwf��͛V9ܵa�����W��U��I�:X�y�$��R��9t���J��u����ր��t��������卩s��wK�����G:rDʃ��
�鷵��K8�Y�i�b���@fkP�3����P�{��� 6(�JG�`����$b��@=}J��/�}&��j�6��I`b�y������Kw�u`��`w>MAF����`noR�f�3]�=8� 3b��u*R	�p$r�����R����b�ٰ;��ڰ%6�K��(���I�1T�4n�4P��<.�Ѹ�3�Ѹ�ۣR��z��]���GK�p���k<�Ζ˹��8�\�Ȝ\�͛m�Bi�I�ӪM]J;S�b2��&ٜSً��j��<j���⻞���g[QGl��L�ͣsi�g�t�pO1˹e��5Yz�l��������m$p�2;M�x��ۧG��v�f��<��j^�n�r������w���w�~k�搳IX��TB�R8�u�#y�tr�g*�]��J�G�F&��98�NJ#����K����37��3�8�)����U��s2o����3=�Vf�Հs������H���rF�R�B7$r;w޺@fkP�3����jn�躒2P�i�Vf�ՀfwK���ԚI��s��qXݯT��"(��DU��� ������ڄf�6����辉a��j����w�*	��c�uh3S��eڻt��LiR�g�+�9�������cj�� �� }����m�C�7���uj������&�^M����Հw��`}̛6��#��)�9R9Vf�Հs��g�m������� ��2��aD�"��"����i���6�Gwf����Vf�Հfo7��M�I)�$�=8� =��@fkP�35��Q;�}�g6K]v-��6�Y�ɷ=]�m�h8�=:�fޜF۵V���Dl1��fZ�9�� �;�����c=�=��֣q�u(R�VguՀfoKw;�$��K�o�n%���rI_|�Kw��Kw?�WU�UUB��M����h���k�[�%���}�IoI�NS��CM�H������7�}���$o��i$�;���I%��I$�y�����$8�q��IӉi$�;���I%��I%����$�3�n��3�*�9�h�c�4��R`)Nx:s%������ �w��|�i����!>I%�����$��\-$�Ϸ��$��8��K�sq�J�J#$�I_|�Z����K����H��i$�7���I%���r��nIRIi$�}���$��Ks{���׽l��X�yG �R�B7$�?�I#;���������$�;��ݷmx��c!#*2�,�d!!"�$ T�*"xA���j�y��Ir޵����B�'%;I%���}�Is޶ZI/�w?�I.[�N�Iw{������9�Æ�w8�՚\��f�Ζ�8ˢ�yn ����4Ҷ�%�IH㒳KϽl��_<�|�\����������$���')��J�8�e����s���t�$�f����%�z����P?���7i�fY�� �>���I,���K����I|���IfԜ��JD��NS��Y��W�$�=�e����s�䗪�~�������Ǿ�jF�S�Dd�I+�K����I|���Ir޺v�K3{������T�2POD=�gh�ݼ���b��W>�nԕp���n��q��:�NΫ���4N������T�вsM�nכ\�_n.�s�D�58�xb�]<��L�ivn��3���m;��k%,��q������\����y���C�E��ݴ*�v��3�C�j��%�]ɓX���g�K�v��M�E�:c��
���������I�����C��X}f�v�v`k�<+�-qR:wc͍�v,.�F��&�M��#1$��}���%�z��I,���K����Ic���H�*�#���Ir޺w�_�in����I/>���I|���Ij����N%"NJv�K3{����l�����`r��`v��ۀ�����q�V����/o{�2w��s] ﾉ�}�@w>U3WT��)���`|����y���Vf�Հ�_Ws�q�rRd�H0���Ȃλm��u.u�z��l�	,���H����[��ٷV۲���v�]9��27J8�vf�������m��s�j��s�6c�ɰ>[ܚ��T�Q)�Dr��z���v�5f�77���z�r%29WqUwp���t���t��֡ �Z�o(�D�P��$������֡ �Z�����ED��T]3K/�l�0묶|���su�H��yᴩ���r7"��BT�))r;sz���޺�>]��Y���p�q3wWWp�y�B����k��v���������RU����`{�����Փ��N���I2݋��Ȍ��=�=�촔3	~iB}���g����BD�H@�#
)�°�0��U�!	A�� �7� 3UKJX�X�L��W�О	Ca"���HBЀRR���B��}�$4J��A�v@�A�@"Cz��YP!|"E_�|ń��i�Q�+�`A��t����4�Z�i�lIX	����
I�,�	��D!0䂧����xf�@�'����W�	�	�؍TC��<��Т�؊�"bꮁ�)�-�*��&�6�U_�C~�뺰>�� �y���2$�#�56�wr��3����2Ն��q��y���Ȍ�Q"M҃R��Ձ�ڄ��ek�3m��q!wWN���u��2��`N�M���E6e׃��,OTRE$ME�Q)�Dr�������t�̭s���� 7{��]���ʎ9)9%X.�vc�V��Ձ�w]_��~�������H�*�$����P�� =��@z^�@��K�����������>]�f��1�_ĩ$R!) �$F	+(M�Z��-�4�Q-��v�z�6�_E���ڙ���"���%XguՁ���`f=�`no]X�ޯW��
�4@���D���K�P�ܙ��չYl��%���ފfj`��)&���RW�b�y��yX��^�o�u`�~c��FD�$q8���W}�D���or����G���Ȍ�Q"MҁVoz���;���o;1�+�ɢB�u(������mB���2��sZ�gu��H%J��)9%X.�vd�"��;����j���ik4�g�����m�\>�ݘd�ٸX�*@��6˭��P\���p�V�m���Mh������ d���NGKY�)$mûX��j�J�iŷm:�/`8n;s�Зb��!��y;iS��a��5
�696m����|P���mv�:r8�-�0v�e�T�y�Z^Nd�p�m��˸n��w�6����W-Y�gf��qmh�������������C	�-���7��AñۻZ���5�trIkb3�/h�9)���E��%J�nI$~�^�+sZ���K�H�*�K�.��n��P�� =��@z^�@fV�@wl�ۀ�D�IH㒬�����^�G��"gv�J��n�EU��U��F8⒬�o;1�+s����;��7�1�H���D�'����q�cj/] =suSUj����w=��n�e�����։��\K����)6P$�����JD��8����������P�njK��D�Mh���s�{f��C�J��G�����*W�H�n���@f6���DD�����U������7����u`}��V�o&ܦ�*T#rI#�2s] 7P��6���� Ǯf�"4)R�$Q�`nw]XguՁ�����7�����Nӌ�' Pn���mQ��8ٷ��X�s��2i��׎N�:6�����+�I%�JG$����Ձ�����7����u`}����$�i�4�J�2^�@d�@n6��mB �t�I�H���1f�77���߫�TИ�S���﷟Z�;�6�]��0)n�"q���V��u`|�y��y�-�C�
J��(�U��3-Xi����{}<#7�`w��Vm������j7\��x��̧N�x}��
5�9�#=;�]-�����F�����@z^�@d�@nkP��6� go6ܨ�*T#rI#�1f�75�@{P���t��g�L��]D���5w7WH�� =��@z^�@d溰;��4��J��9*��;���;�`r9ܛ
k�!$6&�Ow���`n�[��������`|�y��F־� ���jflL����t��w%�M������Be��h��h앺z�6!��Lܷ&��50�ͷ�5�sZ�����<����jn�T�T����޺�>��1�+o;����M����u!C	Q5%\ 5����M�'5�1���'#DD�Ӓ��U������7����u`}��V���r��T�F�$�@d�@w��������ܠ������c}��(2ia�2�ɞ��sj��lX�S��t��g�Ů���K�:xc[�a�:�-�����Wn֩f�k�:�]t��ձ�ilq&���5r�it3��(o;'n�׍�U���7v�z�U\s�6�d�;gF�\7#�9ͣ���p����R����[f�عm�9!�Og��]Sqd�<�-l��zݻ����[L� �q�֕ZV�w{�����{��Ώ�_��!5"nMc�Zȓ����Y�FGBe���M�:X)�[Om��n����cj�ܠ2s] 77�D��i���9*��;���ܬY��������3����$�i�4�J�7_��Y���+�~Kw޺�3}� �y�')�6�I8�Y����@{P�̦���sSw*L��P��`fw]X߿Vo��|������������iA�#�A�܊��T@��l�vu�K�Ҝ�;�J�炜KV�3�
J��(�U��w]X��X�y~��_ �����z�r5R�ܕ5�hܓ�޻��� �JB�f�y�q�cj=uUWMJ�ܒH�Ǽ���?��,�z������䓩Q�H�F�75�@{P���t���t�ǭUMؔi���9*��;���o;o;sz���{K��H'"pl��9�|���p�6&wd"eܖ�ݎ���.�����{��[�&�NA�RV�����ś���޺�>�� �y�')�6�I95t���t��֡�mB���ٽi�(�I�5J8�������E�������>�wٹ'.�!Ԁ�DԔI*��;���o;o;sz����D��7%Iwp���t���t��֡�mB�����\}㿽p��.���\F�L[�'l��v��ٱ�ͥե�[۫J�lU�ʷX뮴�wwu�6u� 75�@{P���t�3��N�AҐ$Q�`no]_�~�_�L���<��9������	��$))rU��w]X.�v,�v��Ձ��[�&�NA�RU��~�\�͛��ٰ;��	i'��nm"|
g��rI�o�Lљ5r�ْ�j������B�ڄ��~m�����ӣ1�XzT^wC �s���aT�f���qea�y����7Y�fV�qš��.j���B�ڄ��������]�!ԁMJ�)(�U��w]_G�2d��@l��@nkP��mL��M��F�RIV˷���7����u`}��V���r���Tr9#�1f�@nkP��6�}�NW>���fiR�TUU56yܵ`N��|���N�߮������'� EE􀊊�� EEꀊ��TW��Q_� EE򀊊�� ����@H$TB#P,@E b�� D���@U"�
'�Q_� "��� ���@EEj*+��@TW��Q_� EE��`TW��Q_�Q_�����)��#��l�8( ���0�/�  )�����@ �� �� P��U ��ݺ!@�B�H ���%R�T�@�� %*�*��T(��@")A"UP���
!(P��R�"DE*��  &   �@  �  �x�O�]'Uӈu���ط3U�=�f�0 }>�v����3\�  ǓK����� =�����>{=�L�� }�������u�sd�� � � �)K0�;�Ynl.���^ wn-P�@�X���Yu��T���� y�z��� 	�   $  �  �� � "   �   ( D���  �
  U
 �C F( D )   R'@ ����   �`� � M���7� 9����Ҿ���(��H��  d  @ �}p�{���v�C�d�����^� < � �� � ���������:@�A������� y�'�K�. 	�l�3���� ܽn�&����{�q]�T���s���j�nN�\�|(��   ()C; �>��ה��+0}ی� }�M������K��9:S Gp���`  ��vr� ��o@�>�]�}�>lQ�L]��K>��-�`� C�7��J� h ��51J��� D��R�h  !تT4��� EO�	G�JR�  ""I��)�@��G�z	�}���������S�ۓ���^�;��J ��C9�QEu QO�(����QE���*�����?������,)
����i������`Uf�!!,�$��5y{�CUU7tA昫ʜ8"i��5i���Tׯ�(2�Kڡ$B���J�k6�+=����ifb�+=
1j�ڛ����)e&���N$&�"U+&�M^]�V;D�56M�>��j�E�U+[!�^��H*�:�s�^M*�:6^�شA��:^���̸*�(���J��iKj�j�Y~���:!�u��"%T�B�H�����O}Y3~�H�)L���D�W�L��5���\ܴM�E$T�+B�h�pca"Rֆ��I��<%���1(1
�+�R�hP(E+��Ѝ:���tq"SP`%qэrW��ʧ�������a�X�"� ���Z�,��랦��^�Id"n��)��BR�����7��.p8K�p�1#FN�k�$)�
b�!��J��BF^F^{���+LN
T�|�n��R���)��E��7E����0MZҸM��G��~ENN 	�'�y(D��[P�%��P�$�T��BM��v��D��C���$���RL�wH�q��7!i0&��.J�˚�F$)
ę
�	���6�� G�� ���B���x�1��Jc���:{Mt$dؒ��J@�# ��!� ����DZ��D��Y��
B��D�C�P��U�;z��/Ә���g���Y0�!�L����o4��d���!��aaIi��˜�9�2l�J��M!J-�n+B�[����z�{X�����$F�~�[s��y[�j�E��R1�V%�J�VX]�S8�.��K��h\6°��IsaX\ ��R$e\	RCB4 ]:B��<Cd�51��L0Ò#��$���=$jbF�l`i��p�
�YbXI�\�:a���$��|!p6pԍ	0З��W�n��5�x�.)�.o��ӌ���w�F�k��6�3����?>�XRS4�=�Ԙt��o��\����Ǖ;�^S*d:h�*b�*~K�=�^��D��'f�����wҦ�٤eh!z��������9]3~X�e��z|���~�#�5	�ׄ0�zM=�u�A�v���e�0��<�/
�ئjm��[��%��eՉ���Uu�ԩ�)�Pqy(�Xx�s�|�@�\��^d��d������;E�xUs�o��L�_���P`U��{�
��إY%^�5X�4�R+V�(��<no�B�~Y7��"R���V��&L�6���ܢ�'I��{�� ���z鬄/*�)�^����M��X���f�����o�2NM���`��Ue*�4��n��ᦻ�<�~�´� �D�[��j�(��R�*���ɫ����s�B��Jd/���y
�+�B�fq�������9�Abº�RKa
%R�c1�HB���n��0d) �,+��
l�B���`F! ��jᡦR�$FWd"���@�Xz���2D��`Da���r�D�w�,���7�����v	D�R	Xԃ�x��"�0Lt�s�$JHӄsCLH�I!n�&��kfJA�0�M!DńZ,�9��!6�K�)0e1!p��D��1Jջ���7&S�U����ZJ_�|=.y��{�����zP�%3�8ˆ�nhB���9��X)?n��K�1��B�B���V�i�-�JХ�����\?/{hF4�!�翏3��ݍ�IH[XJ0"d
H���f�NG&l�!BY����J�0�.RmI��{���S����I)��.�C��4��Bq�Cy����K��(L��NSԐe�8y�F0��B�F0 BNLL�f�RR�0�,�H��Zb��Ni���ڿ�s��q��_�-��+����Dus0L�%��u��8����7��K�f(S���JځM+DӻI���m��F�j
N�G�J�N��W�9��(X^��e�hnn�UL`M7��y��~�,��HY%eˮf6Z��'�d09��VR�	I��-��i��!M+M"j�p��v�>̔�z�8DM[W�z-�ZB��H���9.:p�pt�1�L8�(F�x���1��Q%1ԅ盟�I��#YJ�HQ���Hэ��H��
$H����
a���p�¦�(g��p�FK�3^��� �T�s��
ư��f�)IYIe�Ѕ��! ũ�B�.��(˦ĩ)��s���Ӟ���0��VR`��$2�����wY���ͅ`@��<�5���  �R�!WH�R)�!@m�ܯd4����Vܭͯ%����1�)Ǆ10H��@#�������H\5�N��
a�4����Su�É ��۪�sUIf5�8�.:;��
�`�)��7}�������w�B�Ja�)�(ƌnx�Ls�g��/.i7f��&p�
�Z�0�J��X��)��!\ՋS��4�e�HW�Ƙ�
a�B�1n8HA��
����\%�/����P�dH�HH�"�$@�bBH����J0b@X��o��e�;����NkE+s���vW���J� ���)��kYJ5_�n$-8"S��!ۼxC<��ssy��K���.y��y�)��9�8�f�.o8���F�	�ׁ�Á.:���.h��.o8q!Lӌiyﾄ��R��1�a��u��y�k�J��w~��Q�w9��*bI��!ղ�p���p)k���Z�����I!
sn����~��$���%��\��09syŗ7�
�
a�
`B���V5ׁ�9��g)rFS�?��!.�y���CYt�C7���\�F��8漍3y��7�.��j)�xB��{��0� ��aK�a��!�zK���m�j�w+�^^��	��[R�(F*'��HF{hʐ+8,�����faZ��$H�s�q̲ٔ��V��l��˄0���o봵��g1�\�k��B@��W%b]�#LM\5��04%�Bwdۜ|B@�n��&�X~a}8�1���ЀW�C��Q�@�8�� ���q��/�o���q�Ajʑ� P���������7��H��QŮ�a$)΁�׊@H��x�$JhrS��Ǆnqݞ�Yx~�Sr�)?d�i)��B&g}�m>��󘻳����j���p\7�%��.C?��ۃ�"S����6���(��&��E\K�Z�өDD���R���*D��buqP����l���R���)�&��CL�P��� H���l��yB*�o�V�U��ᄕq �Q��J��<�3���
��+B�L����3S��4���+^�k���������3�_��QK"�L�G����v:��x.�e\�kb]ISw����Є�!/A���xA�k���<��};��H����n���yM��ǯ|� .!z�}j�ے�.�5cő���ŘkD����@�u�M*�
J囜S8�������XD��vm��xyy�RĄ]! �= BS59�u����d3�3t��ԅck"c����?�Q8��/jz�q^fDJ�%]���� ��48= �%e8x�L��RIG�IP����0�\�~忆4��;���}����1�����k2i���!ŌXR����!O=?�~��?5�S
����+\V²~�9��L���`� Im�,��fb��;Q�mB���\�)��!J�J/3��{�>ԉF��BB BD"
UR��aE!i#p�/�<��{��ZD�@��<��?O�Kq���Ӊ1
c䫲&��\�5��	"s7��rO�ķ,"�RK��y��x��u U�_cI|�<.s�N�s����o�H�@��M��%��ʖFy�9����m�b�ҬB�3F5b �\�)��"r�z����%"PQ"I3�o�̼�
H�H����8�<9đ����a�\!L�9t�?R��K��5��i(K��D�	#.lk��p�%Д�hL����2T��<��l�oA�%.B�\����rid�n�.xi��P�B�� d�H]���n���8э0"4��"�]!UBS	4��3b�噘H
$d�)�my�ɬ�F�D�O#����O
P���7�.��@�%[=�[�Xi����R��H�c"��(q ��C��y4�3���
�ȴ|	R1LP�;i*҄���C�J8j���DH�b�b�k"�H�A����F�:�&�e���k�F1@�:�����haӛ���d#E�q772bf�����:2�<�Gt�B��fMT
�U�M��DO/�;��B`�{A��Ӓg��~0�i��sM��� �FE���Z��")$D�
y�X�T�u���*|���΂o�l����eLբo{�0��1#
 �>"D�3��o�H     l�  m|���c3�;FQY��<�I$�qv�����H3�6��k![��BWq���RM��K��}�|?vS�dN6�;�k�����8m�Lt0n*�v<[�U+���r�R9Y�<�V�m���']�grГl��-$$�"��i	m� *1u�]6�lP�u5,M6�� 8�;�1�l$U���*��UJ�� ��e0�qm X�m�v¥�[��;]�@����D�,�8��n�h��%��l�R���` �[G2[K��Z����ܩ��iö����'���t9�V���W]�&�a"�#�R�A�*�bɰ:�j���Im$�v�Iz��i��j��Wl�T�tFl��GjUxsm(H*�d�H���W6��f�I]W�c��l��dk'(���
dL5Vأ����-�.��[�I�p��u)Q�p�TU� &F ѯ\l�[{|���   ,3k�Pp�A"C��K��t d]-��k@8 [x��i٭� u�ӈ�-�e]��_��+�p��{]��K%�m�-��6-�  �e��|  [@�m-�m�M��V���1[[T����v���  Io[��ŵUev]�j� i�5�n-޶��-�&�`8 v�K.��U�n�%U��-+k���oN�U�N �fV_4F�6��mh ma�8��5��m���iҶr������Ͷ �^�\�"�kW�Y4���� ְ �bmsZ�Ht��-�k��vmSiKnۀ�9��C����+�9���er���HL��R�UF�p��g-�  �����r�˥�1���[C�T]qEJ���ڬ�y�Ű� �m�m�+�=���ۖim4�i � �[UN�6S�!u'b)^]�N��,�� %�4�vQ��l�԰U[,&�cf9�[��vEm`�.]�Z�V��
�����V�b��T�UiL��%!:q+vkv�Aj�H��v^]����atG����΍VSnn�`��y���"�����ut��Y��PqjB��!�UpR<Ll��.��*���l���`-�LS���:�{ *����o������*�j��-m��J��Ԯ��U��fUU@�m���j�꺤gkGs��Y�,
;���5UTm��˻-��n^F�`&�mP��s�*�[UU^��1mJ�]T��m�����hC��Rv��ioN�m�`ְ$6���2��k3-$�@r�R��E���ۦ�k"9�V��h�r�:Gƚ�U�%Ir��)�	����	7���N�Z�j\�mk�P�����*���NV,�u�UCb^` K:Y�[��]�^����;`6z�d�1V���V�
T�}�x	�\q��G�i�����yjxp��)2KmuTk9	v�E�dP�m�I�i0�ܻ4�J��t�8��hU�U�;��]�*�B�eZ����:���l 8 -�-[�-���R��3p���*�e9\�x�����g�m�$�v�vk��n�i�m�^R�8���N�Rrl��-�\L��+j��g���ƪ��U��+nN�v-�){y[v�O\�]*��+��Z�nMJ�sv���b�3tꭔTf^8:ci�� ζ��N�m#��u�6ӳ�L��f=�ɷ��*��7*�U*ʵ�q��lc0Y�K�p�m�n�#�i�+)��+�(j�:���6��m��n���n3���2F�t�v�7W
��mH�0���:֝���
����˒�藬Cl86�@%�t�n��~��~��{ o� -�[B-�*M;!t�2H@j��6ZU�(��������Raw)S�2��`z�سUA�U_.�+� �m�f�}�p�oF.K��s�+�V�X"ʪ��j@z�s���g�D��'��Y.  [z٭���r�t��T�RHn���, �c�2���U�Goe�\�*^��;j�Mz��N�mv�b�S�d���\��UUu���U*�   N.�n���m���-��:���5� YZ���N�&���Uv�y��1U�PUx�벁W�as�ƢA�[v��$.��Hm� � D[7Y��Gn��Lìj�@:n,��/'M��
u�R�� x]V9�{-�n˽�m;�I/��|C�[\��z�vp�M���Kvn�km��J�� [��`p   H�` z�n��f���f� m� N���$�oU�8��0O������	�LIxh6ؽ��x�˖ѹ{u�� �M���I�<.�f�*qV'�[6�R����椝$��m�a{r�I9 �-�,�;h� 8 �   �ٶt�� �Yz#h�����;V":�s��)�v�����&[=l�u��ʲ�PT�Qv�Qo`��
�ʫ�mUu��t�A��%�m���
ku�e�K3˰ײ��U�S}@��m� m�8[@]�ӂN$c�'km�s )I��bFt�e���A�-��l�襴8 H ߍ����ޫd��jT�N�V���yj���`'�c���㚞yj�-ւN���9�vKypӗuY^��ɶ� [x 6�@�i 	 -�g[��%^�hI3�V�����4�U�eYV�mC�ӥ�N�Q��'[B�Lm�@�դ K:N�m�A�/I@^�L�ޠ�w�M��ā�>�A�V]��8��UU�� �`��avT�R��d��Z�$:C�-�4kd� �h@f��n��Y*��Iv@S���
���^���UU�Y^j��0�UR��PV�s�j��d���H�#A��鳇dH�! �i6�����d���m��a,�v��
b�j�j�Wf��M̭͞�&�d�U�S�6�R�������*�n{����\�T;x��9�e�m�bœ�' ν,ުsn�mJ�@8_T��r\����
���]��VΡ$�Q��j�:�@tv�����"&��r*�!4s�	�V�L��MPi�I2�V�#�w��+��� T��ږ㊪���eeP��~�{|���w����M� �i-��l�X$��@�3G�����Sk8�Å��,c���	�����m5d�k������6�"�ٶ
�m�M�ҙ�����ˀו�%�����۱�7eZ�&��W�=nD�zM��m����7 �UW���mh�������!����@Z��Z�Wq�Ä��m� ��e��u[n�i1�8�"F m�-�  �Hij0C�%�OY���mJ��6�6ہ#��Ĝ�&���gIm6ʭK����b��؀���    m<�8 ���]t\�Ai���Ϻ�6�� �$ ���ޒ٩�N��m'�_\�4�-�� [4���H�bKk���H    1��m[F�ܶ��('a�
����l�hv����;'����lx�g   9��J���{u\��-�㏋km��<�e�[nZ����$Im l  p  l��`  h�� �tܛ�m:j��ػ`-�[#^�[@�[N�j��u ���4J�Vڕv��4n����pF�Yi5��`� ӭ��k���[Kh� H�`�/'p
�2v�
�A�@6��lb��(��j�^�a��.��am��;K`ػ2�Qg]Am H�6���\ZI^�F�9P*52�c)�J���A���`+������W �V�.�f'm�����L��� ����al�pM��K&E	 :��f�#H�b[<�8�<S��}�����ه���bKm)jb��+Y9�MW��Fu�յ&�6�y��on<s�v��f�S]�΃7m�/�)$�˲�S�O`%���}��J�m�i�����^ �ڶ�6 dH.� pjӶ��p[R�7mnvm��m�� 8  H �H���eZ��(lJ��@:���  ��  ���m�m� [!� z� $ �`e� ��-�i0���kjA! 86ض�m���پ�W,����p�]. �]4���  ��-����M� �p�� ��jC�	����b���uuͶ6ٶ�l    �Yv[��D6�lh � �[@ ��`   �n�$��oP  � � 6���� $[N��� -�4�l�b2to$�,�5��l�0$��٩IB�UCnݎk�eZ��[%��h(I�[-�m��[@8    6݁��k��ﭧ[HX�����޾�$6틦Ŵ~�����7)d�6�r��(D��]V�@�j�lim�6���۷k��Y���I(	zn���M�Ċ�U�l�ζL<f� ��Fդ�l�I6ٶ$�  VƋm ��.�L$5��  m��m� 8��d�M�UHŽe3d���K(g9����3�)��,�"e^kW�Wl��B��3Ê�����{�ܩ?��	�((���ʀH_��<��QU8�@��; ~
��Qa�b@N5��<GEEqQ W�8����<Q]_ȇ�A|x�?���tQ�PDx�����)�Tt}@↡H@� �P��������_8��������Ӣ/�~S�����_OQ�C�T�`���E�W��x"���+PZ��x��"��C}��5����:���z��(�

Q]=?tT:$(��D<�^()��A}� C�A}A �⪞�DTꪸ��+TP���"����@S�_Q���'48"	�D8 ���U��_ڰ����'�D��C
�hz=@
� C� =P���h�:=D��D���*+�?��D���4H/�DCE��X�d��������r�c���-���-t[����
��k��cL�ommFx�HU���Ѹj��d[�
���/O=�Ɵ%�OOvú�%k�Ƚn�FV%'�t�u�È��(�,�j8�b�iSY�@'s��tQC��{AK�������۫SkM��|v��@u�d0�N
�l�6n [H[:N�s;��+gEAZCs�8v՞knq�A�d���Z�ӔsN���*&�LñyN��'�cmՈ�^φp�c�v#�n)�8Ƨ(����増�rn�9���,׶�kR��@^��c�ƭ�йp���Rsq��3l�iI����;$Ԡ-T�8 �����������]m��{=@6۝�sk��]G�[�{kS�֠n1�`T���N����q/����u4U+vα �h5=�k<�l���������$�G;hx݈m!]i���z6;j�k��c�k��)r�b['-en��Rڲkm�=����4"=&�\]uK�\����u[c6w���w�Z��m��N���һ.{�̼�p<x����n7%p�m,���l�˼9%���-��ѯ��y׋��Y�H�U݅͠�<C�ismi6œ@��1q�����F�vy���۵ۓ{&��x�/s��oOjZ���&ʲ��+���7�@�R�i#y��\�:r=�:�gp�vʶ;s� �W+����=���]��vj���'Y��;5��r�BX�Ț�8M�9�;Mmx�VpG\���j��WiYTț�xw.ŵ�^+��e.�´e�n�ػr��bۥ[m�mwܽk[(W�{-��V�:'<v�n���l�궳�fͭ���h�&�v$
;W�D�O�U�E�m�N�9���8�[c���Yz�a �b*����W)պ�j��A��`G�S�gQ.�\�*����؝<�e�
N�1�!�ZHڳ�b��<�&h�:�2M�i�pȡ�	�GU�}85�<P�O�!����
(�D��Z~��s�p�I&i;)��0�^ݳ�Mv��su�m��g��\��9�>�ٝ���v�Í��#u�̤��.E�HD��to�t�ݍwdݻR�{��9���`��ne�v�p��=��ϳ�k��2�Q퓖1����N1�o1�ث��M.f��)g�[�N��i�[iz�tnP#����D`��Ԭt��w.���ͪ�>-C��<�e=�v�`υ{ w(��W9���=��ܾ���ù��*(�MUҳv��������+��%���h����l@)I$Zz٠Uz�@/[4]�@��ex ��29$�*������j��� �s�x�Tc���Nc����j����n=�h��48��NI4]�@/[4
�����@=�@<�1,S!#�:�9��.���٭�苢&���n(4�"��lY�܋@/[4
�Q��f�k�hQ�R~O$ēX�I��O{�f�E�]��)�����#/�@���@�n��|�AZA�X&5!4��@�ڴ��h�I�u��tɌ�L�M�4]�\�P�{ �fh�@�*Q�P"Fń�I�^�h�I����ՠ}zg�F%2&H�(�9m�]]��ܑ����Z�b���ݳ�d��u��F�DR
I��_�����ՠ���N����N'"�� �,���@%� �#5��LU��!���N94�|����x ?� ����a�?H[�@/���YVb��"bS�h�f�[Ԛ�h�V�����x����$�}�M ��4]�@�s@�vp�d���ۆV+�:.�[� �[��w�t����iI�6$�Q�8�Lq�4�l�-v���� �ڦ��;��'��*�ʫ��+J��	7�������@�8-�1b��ń�I��n怫�Uz8����jۭ�n�q]EB�"�73@�ީ��j�/]��/��US���_��39��4>�>�����N&�=��Z�)����z��縳�1\[�Z�W�k�	�=��2;�����g����v��=��FM,�fj4�+S�����w����z��{]�@�QR��H�%1� �h{�=��Z�)�y��~I�I#�$�@�ީ��j�/;V�w[4+�b_��dY�Wu��z�����րշZ�l��U4�߮��!��L����l�zm��]�������y����Q$bMB ��r;rVH�Plpq�SR�@�s��mq�ܦ�5ٷ��3%���1oP�^;9�]������v�e�9��3���v��nz�N�Z�$��K�%�61Z0�r�"\]�;�w,>p���3C�����/K�Vu�F��"���r��h�P�b"��5����i���,��3k����3Ϡ����ɓ&c�3d�̞-T�'%�9s�R�'n�B\�ۓ�lU���3v�,��6�N��t�kFm�i��y�UG�m��w�@/�T�=�ՠ^v���#��c�"QH)&�_z��{]�@��Z�l�s�lƂ�q8��E4k�h��@;��}ꦀyݎ�#��1�$qh��@;��}ꦁ�v��eTP�Ym�rC@;�� _r��>V�h�#@�D�G{����;�]����5j:6`��S��[qn�"V�Ć	9��Xn�d1��y�7U�f^�'Y�|�*�ZT�bg��O�ߝf%�>̘�	�H���v�|t�T+�A�@�����L	0##"FI!BZ"ʣ�1=9�&f�(�y�h�3@U�*�qT'
^���YDd��eh[u�w)M�z��{]�@�����<n<X������sI=f�듫�>V�h�%�vs��+9�"Q@r^�O@q1���V�hr�h�
-e�Y�-���M�ѪI��uνE��Z٬�r�f*.Lk��r�����T?m������j�=�)�U�T�/d�ɍ��1�$qh��@����W�S�=�j�9QX���#i�r-޲��zm�:�,P�Bu��uoK�U�`�8��'�^�O@���@��Z�e4+]�F̘̘��h�h��@}ꦁU�	<i,#Q�F���=����q�� cT/��o[b�93v��:���A���v���h{�M��Z�8��USb�H����`n������W7W�s��@JҭuB�r�wQW�X"FC@�w�'�{]�@�ڴ�)�Z���t1��nG�=�ՠwWt�7z�`G�Z�R��>��7�V���d�ے8�]�@��~����OY�\�^��@�5��t��3";s�9����YI���v��n���Nm��]�V[��	AI�6�H�`܋@^ڞ��v��j�<��R$<y_���@/�T�/;V�yڴ�S@�߄~.d�d��$S@��Z�j�/YM ��S@���S�J#&
4�Z�j�/YM ��S@��Z��˚(چ<�I$�h�����w����n�֕h3����Y��м��P:V7�z{nz�]�Pxyxň����d���۷9;k�۬rs�`z.dv�ͻk�[c�R��D��w�}��~k���5���d�>�a�8؎{a�c1�A��Ѭ>&���r��M�'bʙ��si���ۗ�����)m��;m���uu���/M�%K��4����֕}�fv��\'c%��׬Ps�z�����l��쾇�. �<���y�Se��.nü�vܻ�nLQ�܎
뭐q�p���eq��:�x����'1D�FC�>W�O@��Z�j�/YM�.C�VLX�q7$����@��Z�)�U�T�;�V�S"y1�m�Z�j�/YM��=�h�Tvb���6�7"�/YM��=�h��@򏪑6�����G��=�����@�e4�t�501`����giZr��G[ vM$i.�4]�^ݢ�\F�1���Y�i��@��z�h�#�1���n/@N����������䓾�{y�J���X�I4�^l�w�ӛ�����`{��sE"Ǔ$�-���*�^�WZ�_U�\��v*�sI�h{k�/;V��}V�z�hq�c�VD'r8��ՠ{_U�^X� ���D��p�����+6�dW2�4����V���T�9Y73���:�K�0d�ȦD�B&��x�ߖ�z�h�٠^v���ómb����2���"�7�V�h��h��Bc��G�r8h{k�/Wt��ח�ړ�b���BOU�Z�JT��z�u��]��9G��mݪ\��|Wà� A�H�P�����4� �f�����U(Z_$��z~f��"hz�JB�t!�%�͜��:�$(�����@� �
��#073���9G���Q"�&Y�!A'7�$���	kam!	#�.y�HA���@`��a	q�L���!Rɂ�� ����XD��-�p���04>�>���4��$!"1`_§����0�l`t8$�b�4��� ծ#����<!$CmU�qDї���+G)/��`^�<�� ��X���Bf��ƙ*\``��Zh܀\!S$%��`�«�c<ˁ��_1)y�
V<��B�IJ�*5$�+jE%J�!#�<PĽ�è�S�u*��AH�	���RA^(�?�Xn'EP?D�/�y��<�h��{��͐KC $I��1�7ZV�h	,F��b#�3�Oנ/C�m�NTVNAyuy��/��h&[z��:��@JҭB�ER���;Y��m��
ۗ��og����M��sƵ�k�]�9��܌�*�̨��/332� ��h
��zRJ�11����߫@�;�y,Nb�d��!�U�W�g䊾��}֝h�#}>��ދ�eǊ��//
����{޽}|�G3I�f�듽ێ�$�4FD��-��/�@�}�NI;}���4���ȣG���G����{�џ?�k�6ȴ�S@��N� ��Z}|`�Ev���Ie��{]���C̼T^�V�#�m���t�l���'5�U��7��e�����9��9ZU�/��?��f��-���b�q`�z�տf$}����x�Wܯ\��ۼ����(�����Zu�$�9��\���u�t��U�eAfffV���޳@u�ހ��Zi�'Z�qB�UfF�]f��^��n� �ӭ%�О��OzK70�n���.�
9�[b��]'Lt����Ӳ�g���GV�㮜����N��Lm:���z�s�H�����pm��6:0�{�~�>{y��0��&m<GGk�v��<�I[��vh���#7]Bǵc��ض�a��m���n:fN&x8IT�lλ&�.X��dRR�ݺpÝb�f�۞۲��tG#TR�8$����q��{w~������~ﯼ�w�q���a��X�t{F�nĦ�y\F��c$�3�tf�����3b�x>���@���@��h{���:�s#��4�$�@���@��h{���V��p��X�c`܋@��h���-v�����j�!9�q��޳@��Z��Z�)�w����D� 8�X��@]iV���؝~���}������.�m��x����
�.UOLs���y�t�����i�/�^l��^�5��A}|�@\���[��[u�(b��t]�HZ*���X�|?B�KU`�u^����@__*�31T8W(uP�!�$`�4�_��yڴ_�+���S@���?�LC�"����ՠ__U�^��]����Adn&�LnH��h���Wuz]k�>��>����#Yr&�,�a�L�J�k;���T��]v�Ք�'��g)1F�'�7"����@�ޯ@��z��Zٟ��𾉓�A�NI<���Uֽ������;�v�x�iX$G�WZ���hu$$� 4U��DcUF(Ʋ�Qe�(����S_9F%Y����l�����Eu5r=�������Y�Uֽ�^˚<�H���E�{l��_z��iV���U�8�]��Ed^�� g2ȶ�m���Ƒ��+��G���yn��H��bd�,�����M�h��h���UG�PLMG�H��j�/���/YM �����+rA�r&�M���/���/YM ����j�;�ҊLJ3�o�h���_z��h\�ٟ�
��/([��K���\�r]إ�9$p��Y�^v�������>�l�,��1�8���Xb٦��gT+\��$����l�Ź��L8��g)�8�X���>�}}V�z�h{��=�.��D�"4�NE�__U�^v��z��hL칤#p@��I"�/;V�W�^�yڴ����ز�!�$a$Z^�z�J���Mcu���Q�Yq�yy��*�@s/�:�V���Y�,�߳<~�,m��&�X��obsg��yY /(�m�:���0�R��n��1�4�<8�+���l��y�E��n��pk��y7��V�q����@�{YLl>.�9�f5x��#W.�Mqn�`ۉOn�)uc�H�>ݦo�����n]3�Cӎɹ��㔳�Ց��ˀݷ�ˮ-^0|����ժ׆{lj���ᇆJsX���������m��Y󣭗�t�9=R�&S�,k��p�?߮�O��ry<�݊��jZ �Ef���@��Z^�z]k�;�U�Q�cx܋@�e4
���Vנ__U�_YSjƛ���R8h{����@���@�e4���1��,(���33�*���}����S@/�f���2W�9��q7#�/���:�M ���+k�7���[�0���uk��8�<�-��66��n��$Wqd�9�Ns5���@�e4��h]�@���@���%t��l�]�L݌�z�(Q�@�(�x�	qDE�c�*���;���ͭ�`ou��9r�?��!��)�@��Z��Z}���}>4�M˝*r(�rFƛqǠ__U�u��}�h��@�]K+�&�����Z[)�|�ﾞW�|�Ϫ�<���JB8�1�)���$O� �l��۴`ͱ����뭁�v�&s�fF`��@�����xV��Ϫ�<�S@�qےC�,����^���N���h�,�;/~��d�1�����U�u��+��	�$�9�;��9�L\r�=�I$�@�e4�l�9[^�y�Z��2�X��6���_m�+k�/>�@�e4ӱ\o�+Lg��zp�[N��2�sh�1c��ũ.s:��g��=����[^�}�M����Y�ys�M�nH��n8����S@/�f�����R��I�18����b4w,��*mހ�ۭ}j�P�#23��K�~�_}��/���O� b��|%���NI=��!�M@���+k�>��ߢ_cu��3@U�+�>��XFE�^۴���^�����m+��uk�&��n����Gs ��nG�U�^�ܱ���~��mހ�����eTf]�^�ܱ�u�ށ�۽Wu{�bGةY�ŉ�%���C@�w�=�mz]���S@=˝���f\efffh9�����w�w,F�ߒ����=���mEnEi�zWʴD����a�~�����Ԓ�	������B+{Lg��!�������x%�c	 Aw���k��'�<��RFR~T�q�I`�cXB�!A!=(V�`Fb/!'"#�#�fb�"A�E2~���Oށ�@ &�?P$!BH"� L (؀O���%��2X�����K�
wh�Sa�G
�xF�FA(V�y����~�$�FC9t!��X�C]�$p�~@�����}���}��ꀫ,�F$v�7�#/=�m�{Cdy�E�v�v3�:]��흹�V N�/Y^ή˶�l㎎-6�.�i�b�Lg�8�}���M͌��1l��6d��@v��	�rM%8ӌ���A����^���G,$^K��%'fS3�����P�*iM�퓘�z�aϴc���~�*��6m8�f�]����+#��mV�ݸ�{����	��O](%ȭ(kG�,v����Gp'O�@�Q�F9݁㌶��/(��{u"�g%�f퉛�zp��d�#��n��1vWq��e�fDy�;]f����Q�nN�a��I���u⍘��ڜ��NH��Z��Z9���\ts�iܯkJI&G]��㛁펽�=��(ڄgt)-�r:�+ڦ�:k�a�a;Q�֭=�\g6��Օn\�Gf:��z�=m95/���+vN�Yej�^%�>2�^�W7fj�]�xŬ,��Җ:侎C��j���r�Q=��-+F�Y3�Y���7nܥ�0�狮���`9���;;�
����ꩀ�n�y�p�.�Ի2�ԬOo<��0+���uriK��9ę
��^Θ��;�6��;5!�G`��'��	sU�GE��7Of�Nz�,����s��X�Q7����zۇ��ۨ��s	���\u�t��@uִ�
��Ƿ1�㋮�⚇����v��MkS�ZU]���!p�pu�}���[<ä�\F��T]�4T:'3i��&����Kmm+H��J�������T�F�>4S6�0h�*m+�U�(4N����]���Ճ�-I�y:�[���)�v玳�mc�$8W;�)˥X8N;v�i{�'!�iMD6��!���۴�n���;W�cˋiܼ���Ķ�T�[��R��Ű�/[��^�܉d�:w/I�R�؆*���*\n[���� �����������gH]�V��L�Z����Z�X�SL
����%��T��UJ��ɮ�]��u^����W�uExqQ��~u_T�)�� � *~	������������ـ�Lɔ�>��R�ջ&a�TK@�/<�s�pK�Y���;��p�{�=����n׉:�st��u��s���Ĝ [�8�L
���\]b]*����6�n��g��t��hx.^5��hLY"�7 �_2#z1�p�n)�.��6�뇄c9��������k��]�6��)	�a�|�ڛg���ɻ���	��G�͇+�e�UF]�V��:��^�\���'V}���S;��h7On�[�����|�W�Y��G�����4.Y�u$��G�M;�X���fF`��@-�7�ى���@tӽ��k����٘��VU�Yw��v�h
�+��雷�g� ���@�X���/#.��+A�;iހ��h\�A�Rx�hL&�k*��32�2�V�hf�O? ���
�W�x�/���?I$#������M��]e�עq�rL�/N������<rc��F�qx���uv����~��������V�(�8���Qf\eff��I�s���5�1�� BP>ݟ_��rI���גJ�W�f${�>��RF�J&ۑŠ|�w�r��G3T�zv�huªW�]�T]�qY�z"���@O4V�h8�vӽ����Y�FY�efV��r���x�~�N�V�h�k4� �mF��$��'.Dx��{.�9��RF�u�W];q�����������'ñhm�#����Z����fg�LD�a������Vՙ�fQw�Y�ZWʵ��EP��h�w�r��\LL�L&�k*��32�2��3@T�^�&"fa�D�Dݼ��@nӭ��{���L�ɻ�n��ȡ�*���?^��~�h	_*��q3޳ ;>ˉ�k�c�8G�@�ܠ����b!,�_�m�4K���:
�����k��+Og�a�kkm�Ľ�f,�b���qq�O%ћ�������|�V�HUf ݧZ%��.V�ff"P7mց�	��0��.�˸�̭%��3335C���	�u�%|�\��L���E�̻�������@t۽��Z9����nۭ7��?E%b��2r�����/C�3鉈�����@��ޭ���I����#��*�"������￳�kDd#ȓr)"�-v��LL�oY�M;�9ZU�~Q����[�,v�sӲ�v��sڞI-�nND����g�0ur:][���{޻�[s��0�l��&����V�8����@ݧZ�^+�<X� �FҐ�z����>�����׽��=�~���k�������.'��5�1�I$�_}��/>��������3@7���գ#+0�ʻ��3/A�LLSX�h	�f�/��31I�u�*�����pU�q��Z%��=33鈈������ޭ���=��r6��lh��M�u�.�Bk<���S(���#�\Y�]���w<�go+�n�N�9���X�7V��wl޵G�[��������k�i6K���U�nyՎ7��y�7;��t�9۰� -�-���N�vv[e��˓	��nN�e�?C�:ϲ���8�u�����a�qk�l\���ź�����b�KOZF(*��ʤ��{�������.;����\m�Y��k�%�&roi��k�#�g�9�گ�����k�����xp/{4V�h��9���@�������o&C�h]�@]|�@� �K5��U��J2��r)"�>����SO�g�ľ]��@����@�e�"��bBr'"�q1M�f�>o4I+�s3Mbk@�^+�<X�Q ���4�l�?�1>���g���;~�%��>��o�������ѵ���L�
�m�pݒtnǲ���؞^��yn����ݏ�����c��33��{4�ʴK�bg� ���>����2)�m�I�y�Z�~ə؉S33.b&wKo�&�@JҼ�_�G2}O���3wn\%��p�ݼ��{<h�,����P�y�5iց��W��dE�f^�LL�ߗ���~�h��h9���m�4��e��&2�9$�:�V�y�Z[)��f�}�ei`����)�{+؝�GI<6���vs��e3�N����������h��&�RE�W~Z[)���L�~�Nۭ1�2������2�2�K�&"f�7�v�h�U�~����qQ\������!�~�}�rI��{y0آoU߅�k�-����n�ƞ;�Ō�I3A��D�X�hZu�.X�zfff����@�������B(�d�E�^|�@q311=g��怫�� _t~@D{$��30�7(=(Wn�!�T9[6�&Z!-���$���-F^&Q�@\� �,�rV�bb"P7iցVw�/��F�oY�g옙����h�u�w,F�}333vv?��kL�i�7$����4_Z���LL�$� �y�wt�����2/*�//34DLL�7�ր��h^�y&�%ê��?*�f�Ͼ�I?||f�rLHND�Z[)���V�h	_*�=330�<�Ȼʬ�3�:l��\ɶ�+��goW�3pvt�7l�?���9�.�ܲn�[�?I'���۠r��@J�S�����	�f�swEYp�*,������Z�"fj��:�x� K�o��7g�~.��w�VUݗ��Z�oՠrX��L�U��@��zsʫrD�	#m�r-4��h��@�I^���V��ap��(%�C�G ��4�3���m����@�D�0D�L��w���g��,�㷴&�nN\u�p����!L<ז��h�6�B��S��S��dѡO����45�c���F3��=�H��v��q.������0�7��"���9����Zy�x8S\�	�s�rgV�Oc��]��u��8��	����N#�lh��� k��p׀Ά-v�Krs�q֤�Fꇸ�ua%�5���GZ�{���}���H�U�g�Qv��5ť���7C=�$�0�˺���m7W��{��GW�I�{Vwc �{٠.�U�rX�133��|�ho�}�(̓!#�9�y�[�~��Bo������� �y�t.�F�rLHND�Z[)�r�^�߳���1T&�h	�u�(�+�\TVee�f]�fb&&&���@o4Wʴ=*?�*����NI'O���)��2l�̽ �hfb"S���	�f�Ժ� ��䑕1	LQȖ�D�m#��գ��3�� �~��.�M�n��$kNZsՒꪊ����W}-Đ��$-�|8^!X�%�ܾ�0?�@�DȖ%�{����w�{��7�������5
��/M�S�,K����g�x��t��8�$�<1O�;bX����br%�bX��}�O"X�%����S�>Ar�D�>�ߤ�\ݷm�l��w6q<�bX�'�{�br%�bX��{��y���lM���]ND�,K���N'�,K����r���n�Y.�br%�bX��{��yı,罺��bX�'��;8�D�,�	�>�߳�,K���'>əw!�l������yı,罺��bX�!���N'�%�b}��f'"X�%��w��O"X�%�������:J8L,t�nX=�(qPm�y6,���l�4���I��?.����}hu����۩�Kı;���q<�bX�'r����Kı=�����~��,K���S�,K������,�vݶn�[�8�D�,K�}�br%�bX��{��yı,罺��bX�'��;8�D�@��M�b_�}�e3�C&�����Kı>�����yı,罺��c � [H��i�Vx���`��~�O��)zR��T����(�#�G��P��T�XA��@=�1c�h%��Wu�sa@�YMU4$$HXFXOɊ`H�4]RD�c"45�BR�6?�V4�#e!T!x����"�`�2[��#<�B�$���$້P.�֤�A�JR#�JZ�
�$	,^J�s%"	s�$rV6�j��`�#�!r"��M�A��N%`��TB��=: >�y����R���T
�~ �P�E>G��&����Ȗ%�b{���,K���vfm�ٛ��.nnq<�bY�$����Ȗ%�bw���yı,N����Ȗ%�b{��s����oq������k��4��E��%�bX�����yı,>?m�ى�Kı;�}�q<�bX�s��ND�,K���雰ݙ������Q������.�zǣ]��c�퇮6-�����8N\3M�I�f����~�bX�%�w���Kı=�����%�bX=�{t?�D�o�ı>�����yı,O�.�f���݌����Ȗ%�b{��s��Kİ{���r%�bX�����yı,K;�wS�>��,O{�s�32�l������yı,��]ND�,K����O"X�
!�SblK?���ND�,K�����'�,K���N��K��e�wnn�ND�,K����O"X�%�g}��r%�bX��{��yİ:
�+vo����bX�'rv�'r��ۖ���wgȖ%�bY�{���bX�������ı,��]ND�,K����O"X�%��vP�;.��R���집�ͽE����#[Jg逸m���<9㗧=��5^ﷸ��%��w��'�,K��{۩Ȗ%�b{����"X�%�w���Kı?{��>��)�2�fe���'�,K��{۩Ȗ%�b{���Kı,��ND�,K��{�O"X�{���~H~f���^�/w��oq����gȖ%�bY�{���bX�'���8�D�,K��n�"X�%����I;�i�e�&m�͜O"X�2&O���r%�bX�Ͼ�8�D�,K��n�"X�%��w��O"X�%�����̰�6�Y�37wS�,K��{��Ȗ%�a��?�����ı,O����<�bX�%����Ȗ%�bq?�}�e'�.�ass7fL�lE]���ݰ�]�:3�t�p졮u���RՌ8wlf�����u�q��]ͷ]�%Ka�ջZr���OWl��77	��v�&��UTԥ��ǰ;��~f�f���c5��c��g��X�<�1N<st�6�ӸD�z���l(u���]���;X4<.˶"�aΘ�c�fҚ���b�3�tCE��$]�[n?=�w���>��������n�=X�yw)�]f�������m�8�۷\j�@]v���C�3h�[;���������%�bX=Ͽ��"X�%��w��O"X�%�g}��r%�bX��{��yı,Og�휚L��e�wnn�ND�,K��{x�D�,K�����Kı;�����%�bX=�{u9ı,N���'r��ٖ�ܓwoȖ%�bY�{���bX�%���<�bX�s��ND�,K����O"X�%��vaK��0�M�����Kı/��w��Kİ{���r%�bX�����yı,Jv��&B��������VZ.��������yı,罺��bX�����N'�%�bY�~�ND�,K���x�D�,K��e�m��n�f�P�13�t]�V���^�h�<>�j��n^�Yu�X$,�iW�������oq�����vq<�bX�%����Ȗ%�b{��s��?DȖ%��w�Ȗ%�b}��XO���e.ɛwsgȖ%�bY�{���� `�� �|�lND�>����yı,�߮�"X�%��{��'�,K��L�v��3n�������Kı=�����%�bX=�{u9��"w���yı,��59ı,O��N�%��滹v�n�Ȗ%������I��oӂH$���q6	 t'�;�}�q<�bX�'{~�9�并ɤ�ۛ�S�,K����gȖ%�`���S�,Kľ���'�,K��{۩Ȗ%�b���!�}ni�f�s;��u옮�i��t��\��!H��k��<�L�a.m�n��n���ı,K���jr%�bX������%�bX=�{t>Q�DȖ%�߾�Ӊ�Kı;	��R��.I2n\���Kı/��w��Kİ{���r%�bX���vq<�bX�}�59�S*dK�~9~�t�nL�̹�����%�bX?g~���bX�'��;8�D��a$!$!!	�@�5U�*p>A,M�g��u9ı,K��x�D�,K��[ٛ�72�l�77n�"X�%��{��'�,Kĳ��u9ı,K�{��yİ>QY�~��u9ı,O���	�i��dͻ����Kı/o��ND�,K�V=߾�8��X�%��w�Ȗ%�b{���Kı ��oc�����u����,��k�(���]:�]S\�nZի^e�<d�����Ȗ%�b{��s��Kİ{���r%�bX�����|�3�L�bX����S�,K���'>%��滹ws7w��Kİ{���r�r&D�;���q<�bX�%�����Kı/��w��Kı=����ܹ�i4��sv�r%�bX�����yı,K�s�S�,~dL�{��oȖ%�`����r%�bX�=��;�K�\�n�[�8�D�,�@��3���S�,KĽ�﷉�Kİ{���r%�`~�	肓b^�;8�D�,K�e=%.v��&Mۛ�S�,Kľ���'�,K��F�߮��,K���s���%�bX���v'"X�%��g���rd�0�il�4��'gl	F=�u�m0�Qt����]���{ܯo��k��TVk����q�����{���Kı?{�vq<�bX�%�݉Ȗ%�b~�{��yı,Ozi��M&�R�w�۩Ȗ%�b~����y�U�+�6%���݉Ȗ%�bw>���'�,K��{۩ȟ��*���,O���a?��L��73sgȖ%�b_￷br%�bX����8�D�,K��n�"X�%�����Kı=���-�2ۦm��7wbr%�g�!"g����yı,��]ND�,K���gȖ%��2&}߷br%�bX������5����w3wx�D�,K��n�"X�%��{߼�q?D�,K�߷br%�bX��{��yı,N��������|S:���i�����+OR���1k8����j�ʝ�]#��t�}�E�c�<��n�pdv�Wy�n���QN���&�<�V/n�^:*Όc�8�5�a�t9q���Z,b�XN���x�a{C�MzR:�)ǝ� 8��[-t�z�n�g;�ݮ5s���tCc�8�H�t����9��[=3���I��uw��]U�<�ɓwl�[�4˹�5�9�<����p�
\u���{�r�ny;q�
-���=\���V�{���o��k�CF��%�b~���Ӊ�Kı/}��ND�,K��{�O"X�%����S�,K���L�a.irY��.��yı,K�{���?���ؖ%�����<�bX��}�u9ı,O{�vq<��TȖ'a��[.}fe�&��݉Ȗ%�b^�����%�bX=�{u9ı,O{�vq<�bX�%�݉Ȗ%�by���m��&d��˙���O"X�|� ����r%�bX���}8�D�,K�����K��C�.��������%�bX�g��i���m������Kı=�y���%�bX���v'"X�%�}�{�O"X�%����S�,K�ﳽ�	�ۍ�Qײnٔ��չ��ճr�+ΞoN�Mq��RsY�k���F��$l��i�~�bX�%��n��Kı/�����%�bX=�{t?����lK����N'�,K������m�6R�7wbr%�bX��{��y�*�(���L�`�<���Kı<����yı,K�{��,K���e��������w3wx�D�,K��n�"X�%���gȖ?���/��v'"X�%�}�﷉�Kı=�۷�m��.�wnn�ND�,���;߼�q<�bX�%�����Kı/�����%�`|L����Ȗ%�b|ggL�2K�f�7s%ݜO"X�%�{�wjr%�bX��{��yı,罺��bX�'����O"X�%��{/L9rf�f�Ke���˘�9.�]S��pv=����v�z��tf���@�Ρ��}����oq��{�O"X�%����S�,K�����Kı/}��ND�,K�{�߀���������{��7{��v�r%�bX���vq<�bX�%����Ȗ%�b_��w��Kı=�v�4ۙ��7�۩Ȗ%�b{�y���%�bX�w��"X�z�P~X!��E8X�D�o﷉�Kİ~�~���bX�'L�v�t�6e�m͹����Kı,��ND�,K��{�O"X�%����S�,K�����Kı=���-��e��!p�wu9ı,K����<�bX�s��ND�,K�w��O"X�%�g}��r%�bX����Ky��1ɹ�B<��br՞��9RnpG��	�n����ڜur�ön�+KW����X�%����S�,K����oȖ%�bY�{�3șı/�}��<�bX�'{e��70�Mݹ�u9ı,O}���<�bX�%����Ȗ%�b_��w��Kİ{���r'�S"X���>̖���f�d����%�bX�}߷S�,K����s��Kİ{���r%�bX�����y��{���n�6?"rlꚯw��D�,K����<�bX�s��ND�,K�{��'�,K�?(�W��0\@ �x�qCr&N���r%�bX�����i�ne����'�,K��{۩Ȗ%�a���?��ؖ%�bY����r%�bX��{��yı,K?t�ܻ!�$pU3)��{9���\v��D-⹌&A��S�E�U��˶걤b��Ou�,K�w��O"X�%�g}��r%�bX��{��|��2%�`����r%�bX����|e�&m͹woȖ%�bY�{����șľ�����%�bX?g~���bX�'��{x�D�\��,N����d�s.�\-��ND�,K���oȖ%�`�=���K�F"w�s���%�bX�}߷S�,K���e���,�������'�,K?����S�,K��~�Ӊ�Kı,��ND�,�T�=�﷉�Kı;�7�6�M&��ݺ��bX�'����O"X�%�w��Ȗ%�b~�����%�bX>罺��bX�%�V�YA�IC:Ed<R
��Z�HFU�4!c�A�H�#�V�!^�ܴ�����X[����
�� @ "!@�������,'��z������� $IC�"B*B�0)�� �R�ea	&l6%�BHE���"�!	��@�@d�D� ��Ĉ�	$�@���`� �1!,�
� ��s������2��&�zF#؉��Q:nM�m�n��;pc<�ݎ���h�/VջAmJ�8(�څ��7X��e^����an������D��q]�t�56�PEC����2�M��6�C��%�q=F�l��J\����:ӎ�B�f-�&p]�;�IZ���Ʀ�d���P�x7Z�*LH��W�T�l�	��;ve�x:�g��ۭm�d�"Q*�=<�@p�0��N�� ��5�3�i��p���8j�oku��1:p�O[��4��Vٯ;.���6�j厔�O'8�I�9�v�����E��3ȰfW78t�;ql2�P#��T���l=��B�q�&�ڊr;�s��u`���8g]$���4�euĬ!wX�g4t�m��s��Or�؈�;.��U{����ݷLvz�:�FѰ��:.v&��:���l�%<LZ=vY�/C�L�U�x��']�۰b9j(�yy�Yq���� m�u��n�5ιm���ۓk�Tpl�̔���3b�'&���2'Ji�If��<u[y�p�5+�Ѻ�]x��n��Q\v��$�Y�Iv�Ħ�O%YO8:�ؒ8�]�%��Sm�\*.��I�D�]�>�.5;�t�ۆy��v�%��Z�@�ێn^�q�Erntn��3���"a�m�n�]��]�����W�V��ƕl悎�'�sD�⋞]���v���O5������b�ݮ�=[ꬔ�ܺ�ظ�T�&q�y�6�"՝ˢ�.D�V�VҼ�J^vT�{qsv�=np�%�c�-Ճ�hu���ms�]�\r�ͮ�w;vhNI�M���]zGi�:��Mm�Y{rt�T��"�!��	�zv�r�74�$�&�.�R�����1�4٨��ʭ���G�7n:C�gV�(���vd�:􀍯]��-�נ��;����m�S[;�@�W'[� �6GSE6����bɌ�]�V%��mT�N�U3{T�l��K�6�s�kK��ET�D=�������j
� E�54<E����!��ts�����=m�����[��;O]�2V�<l܋aέ����C��ݪ2�C�[�!�S�c����9�:\'i��N�a3�2[�6ur[&=m�2Eղ����U�s�1q5�P��n�[�f�� �wmŒ.��=�,N�]���;��HVx�㣯Y�c%ø8��-v̰U�6�j-�d�\��5!�E<~������xw��r�����d��Z�qu���W�Y���b`6�R�yn��>P�0�Ne�晶�������%�bX�w�n�"X�%��;��Ȗ%�`����|<��,K���N'��{��7��;�m�m96uUW���ı,O���8�D�,K���S�,K�����Kı,���"*+�����������77.�˙���O"X�%�߷�jr%�bX���vq<�bX�%����r%�bX��{��yı,OI���dۙ��7$�ݚ��bY������Ȗ%�bY�~�ND�,K�w��'�,K�I�{�}59ı,O���d�˴�%�ͻ���Kı,���"X�%��~��^'�%�`�����Kı=�{���%�bX��ٝ�ٺ�V1�'��$)�;Fb&hХ�<�:rZ6n=������u}�K�q�Ѹ���D�,K߷�Ȗ%�`���jr%�bX�����3�L�bX�{�۩Ȗ%�b{��ߋm̒��&fۻ���Kİ}�{59�0
�OTO�LybX������%�bX�w�S�,K�����Kı;'�޻%�0���wvjr%�bX�����yı,K?w��Ȗ?ș߾�Ӊ�Kİ{��jr%�bX�0��;�-�2m7w&��'�,Kĳ�{���bX�'����O"X�%��٩Ȗ%��2'{��N'�,K��N�v{Z6uUW���7���{�w���yı,}��ND�,K�{��'�,Kĳ�{���bX�%��w��݀5��3��8X4����!�N9i��^�l�q,�%�]Ya�:,�7gȖ%�`���jr%�bX���vq<�bX�%��������lK����?�Ȗ%�b|L>��dۙ��7$�ݚ��bX�'����O!��"dK�~�u9ı,O~��N'�,K������Kı;�z[gL�Hf�\��͜O"X�%�{�sS�,K�����K8���2}��ND�,K����O"X�%��L�m�e��k�d���ND�,K�{��'�,K������Kı=����yı,K=���Ȗ%�b~�����n7a�3m����%�bX=�{59ı,?����Ӊ�%�bX�}߷S�,K�����Kı=�(�m�r�E��e���l]����)pD�5������kFm�y���ڢ��Ȗ%�b{�y���%�bX�w��"X�%����gȖ%�`�����Kı:a�wrK�݆�仳��Kı,��NC��L�b{���q<�bX��ߦ�"X�%���gȟ�S"X��w$�|fm�$3wwwu9ı,O~��N'�,K���{19��!�2'{�>�O"X�%�g��u9ı,O:t�fe�4�n�ɷvq<�bY�@�?w�MND�,K���N'�,Kĳ��u9ı?$��
*đ�A� ���HA�H�#,c"F �_>"���!$� Ȳ��ĉ$d� DaA�!E��BI!8_�?(�'��Ns�?�Ȗ%�b{����C��&�g����oq����y���%�bX�w��"X�%����gȖ%�`�����Kı;��?~�c�q�m�魅�5�:�4I��<��$�	x�#v�{���o�;;[��n���Kı,��n�"X�%����gȖ%�`�����Kı7y��x�$)!I�E=D͔��rd���ND�,K�{��'���J�M�`�}��S�,��>���Ȗ%�bY�~�ND�,K��ys��s$ͻ\�n��'�,K��٩Ȗ%�b{�����%��C"dK>�۩Ȗ%�b~��}8�D�,K�=.u��l�����٩Ȗ%�b{�����%�bX�w��"X�%��{��'�,K�����Ȗ%�b|wN��,�5���ͻ���%�bX�w��"X�%��}��N'�%�`���jr%�bX����8�D�,KN���{����6^y�
�3��WP]�ϰ U���W=�����v�!`�m�Uv�-g�X�;N��9����JѬ�'��:��N��;F�K������TV�"��m�v��פ�yw��lc��-�:�� n�uK�vUN��e㮮�ݹF�孳ی��:�l��%��ƷW��V����+<��n�38wF�]t����51��\\�S03g�����w����~�߮�IB'V{{6�집�!�[&�m��.$
vȅu�٣�nݻyfE�v �~�bX�'}��q<�bX�}��ND�,K������/�6%�bY��ɍ&(��b�����2�ʬ*̬�'�,K��٩Ȗ%�b{�{���%�bX�w��"X�%�����'�?���M�b}�f��3f�̓v��wvjr%�bX�w��É�Kı,��ND��ű?w��r	 ��;5�
B��6hD�����1B�G�2}߷S�,K���~��Kİ{��jr%�bX����O"X�%�����R���Z�w��oq��'���q<�bX�0>�>��D�,K���O"X�%�g}��r%�bX��{��Za��i�f����s
n�gK�v���ݸ���v����|�KY����ɶ�oȖ%�`�����Kı=���q<�bX�%�ݡ��"dK����y��%�bX7�I��Ie�ۻ�S�,K���{��� �q�D�,K�s�S�,K������yı,������"�����>���IsZd�ܙ�q<�bX�%��?��"X�%��{��'�,K��٩Ȗ%�b{���yı,Or��cۗnܐ���ݩȖ%�+"~��>�O"X�%��w�Ȗ%�b{���yı,K�s�S�,K���Iù�se�3mɷvq<�bX�}��ND�,K�#��^'�%�b_��mND�,K����O"X�<ow���׎,s�mٯr:�R6;&v-�l��wm��V]uj���H=�7wf�"X�%���oȖ%�b^��ڜ�bX�'��;8#?DȖ%����19ı,O��-��7)rM����6�<�bX�%�ݩ�ș�����q<�bX�'ӻ���Kı=�}��y���M�bvL���.fn]�ْ����Kı=�����yı,N�w��,t��"A$@��H$"  #$`�@$�"��h	�D)� *:!�P��,L�~��<�bX�%�����Kı<���&�6�r�8�D�,�H���Ȗ%�bw;����%�bX���v�"X�%����gȖ%�`���u�nͤ����٩Ȗ%�b{�����%�bX|ϻ�mO"X�%�߻ϧȖ%�`�����Kĳ������NؽYgO;�V��u옮���)�Ӟ����<
F��\��ˈ�cvuN��q<�bX�%�ݩȖ%�b{�y���%�bX���f��&D�,N���8�D�,K�N�c��˹�����9ı,O{�;8�D�,K�����Kı=����yı,K�s�S�>ʙ��ߤ��2�6͙��ۻ8�D�,K���br%�bX��}�q<�bX�%�ݩȖ%�b�9��x�$)!Izʞ*�n��.�k6n���KϘ��~�'�,KĿw>ڜ�bX�'����O"X��� �FB0@�T�X�D�$@�`��j�H����ND�,K��岝��\6��ܛ��O"X�%�{�wbr%�bX}��ϧ�Kı>�ߦ'"X�%��=����%�bX���{w!��9S�ι����b��!��M��Ѻ�Z�$Jv��/lCT��-<�n��k{���{��'����O"X�%����br%�bX�������L�bX�����,K��ޜ����4�e۹�8�D�,K�����Kı?~��O"X�%�{�wbr%�bX�~�;8�D�L��,��>6Iw6�˻7wf'"X�%���É�Kı/}��ND�,K���gȖ%�bv{����bX�'rv�N�&��&M���Ӊ�Kı/}��ND�,K�}�gȖ%�bv{����bX"w߾�q<��{��7��;����)�4�ow�,K���y���%�bX|�w�LO"X�%��~�É�Kı/��v'"X�%��(~��O� �)��~����ɹ�aM�f�q����ɱ�Ƣ�r�E��L��iYA)�Cv��]� �Y�/'����l�@`٭E�Z�i�VmE��e����E�j�l!�1�5��עt�۴����ǚ㉻[6�������Ĝ�#� d�,�����;t�s��K��6N�獏]���c�K!�mS��s1H���yX9|�པ?��������w��ݿO�sݡh�v���wKv�Yi5���:�:�\��dr�F5��3tT�gXv����%�bX��ߦ'"X�%����É�Kı/��v��&D�,O~�>�O"X�%���2�fm̗,�˙�wf'"X�%����o�*�"dK��۱9ı,O~�>�O"X�%���{19ı,N���d�nRᶖ�乹��%�bX��{��,K���y���%�bX��w��,K��?w���%�bX���2�2��d�.M�݉Ȗ%�b~���yı,Og�ىȖ%�b{����yİ?�D�~�v'"X�%�����������m����%�bX��w��,K��?w���%�bX��{��,K���y���%�bX�����.駧uL�t�6Dvc�'1��q���x�B��py�;&��dW$�e�e�{���ı=���q<�bX�%�����Kı?w�vq<�bX�'�����Kı:g�ӻM���n�n��Ȗ%�b^��؜��/D\>�bdK�}�Ӊ�Kı>�ߦ'"X��������y��L����L�k���h�3@_v#OU*��@>i�}p�<\Q2	�Hh�Jh�������_y��:C��ݕa�uvefa�u}��L�LW�<���}؍�Kf6T��QTfeFFUT����]k��f�<+ΞoJ\*\y�9��u�K�8O�I'�~�w���@��)�w�)�z���=�\mFH���I49b5��3@䱚�r��:1E؋��Q77Wcso�n�L،\�HFy�1�
4�saʆ�d��E�P��c$������y�M����I�	MRYBqn&EVU�E%P�Z�c<�`�$� KP�B@�R�R1X�!U"~0�"u�00�I�_�I����!�Fa!D.Q
6�ŉ����<� DNe0B&��97.���[a��1�3��Ƒ��$��Ѕ�j��ca�(�/�(�_�8���,Ex'PDhz������z��^�)�Tx*��]�y��o$���F���+�eU�xff������hy�4�b4�� ����n�$�nf�yz��e4��;��hmǣsh��!�,�A~�u�i-g�lg�՜٭������g�y,�Fm��癘�E��M������;��h�w?�@}���(�4}��&E!�_o�o�f�Ic4�y�~K�/����#�F�"r-�uz}�4-��/���/��¸A?�$�dq�z��y�|�3@__*Й陂>�fb��>�4l���'���L˸E�A���h[)�^}V�˺� ��4����d�h��x������.dl������I^�Y/G^��;!��ꎒL�YD���}]�h���-�@��M ���L�p�#�h]���A�o4��h�ʷ�35A�R��D�r$�)�{��M�e4�J�~ZV��Wg<7f"�y�y��蘊��f���ZWr�U>���(���aqHh�U�l��0��`{��`5�!(�Q0� ���3��@�	$R`�#����ٷf�bl
^pfɌ]6���*\c�Uջ"���y�Yր�C	W���<'��G���nt�4��$�{v'bI\	[<Fy��Gu"ѹ��X�n�h���cns�����ý�Z;i�5�E�ՀY�ձ;�^����y�v��9gcL���Ui���ۗ�h�eqg���'ˇD�Âq�"�jwn.���t�^��Krw�{����3����u^�´kQ͠<ruY@:��;fƸH\������{���FH��D�\��z}�h[)�^}V�}�\����q8��l�?%��_*�;��o�'�v%�u�E��I�w���4Ϫ���ύ ���h��."~��•RCC�Mbu�$�ƀ/���X� ���aU�QY�^eh�-��������;����Z}h��TF�^drB�:�b�C<]lۃg+��;6X����K�tg �L�D�r!�Fۙ��f����9'�%����x #?A �`�`����8 ����&s�LҖf�f��A�666>�߼8 ��o�i�z�)�P� ���{x ����g �`�`�`�~�ﷂ�A�A�A�A��'e̖�L��v�m�8 �����A�666=�~�8 �F�����o �`�`�`����Â�A�A�A�A��˟n��6�fdۛ���A�A��X�d~����|���������A�666?���|���`��w�^>A����M����LvK��ss��A�A�A�A�{���� � � ء�	}����pA������ � � � �;߳��A�A�A�A��ι��ve!nc�nᙑ̘�G���N׵Wz��t�z�ۡ�9��7�Ν�f\&�� �`�`�`�������lll~����� � � � �;߳���lllo����A�666=�>&�nM6�m��pA�666?w{����lll{����� � � � ߽�����lll}��|��`�`�`�{��4���Ywf�����lll{����� � � � ߽���� ؃A�B��r9��xpA�666?{���A�6667�gO��͹�fL�ͻ��� � ؊� ��w����lll~��8 �����A�66
� ���}��|����s��2��n�Y��3w��A�A�A�A�߾����lllP�V*��}�x ������}���|������~�>A����?���۶�d8�/�u�/k�,լ�\�^ʓv�����g]����ԗ����|����ݹ��A�A�A�A�������@lPll~���pA�6667���x ����|����}�v��nٗn�fM��x ���}�|��`�`�`�{���� � � � �߾����lll}�{����?�`�r6>��$�a�M��v������lllo����>A����~�Â�A�U�A�A���ׂ�A�A�A�A�;߳��A�A�A�A��{�K7&M�p���>A����}���O}��y$���s�z����a�"x!Qr(l f���_w�sy$�N���a�iXVw��}���.�w�����lh���m[Ƞ��#&�(�*�T4�d�nr[Z�"��Z�ጜW�Z3}����HG"���= �������� ���h�\�"8܈c��#�oX���i��]�����{�:yJ�J��i���ۚ.� ������P|۱$��HD�h�j�9wW�޳@�۹�_G��n$�Q�Ȝ�@��� �������}��&(&N���̺nXY&�fm��&Q=T��h�7�b]��%ݷ=t��GcZB�Ö�y��&�q�Y�nL�t�@��l�B0cgmX8��q�;X
��{A�7M���$�J.��i�f8�E�WsX�(�u��'��l)�������n�p��y�(	��
�In�tpw\��Q ��P&�$�;l�r��a��gQ��v�j96�$������cq:es�0;�c�M�kj���%,V�	��=�tn2^0Hݬ��{/\��a��� 3������r���ӻ���O�����4�'&��s@�_U�r�@<�f�ݝ�FFOȑ�'V���,�ަ�޶gsLؤXNe�eVa��Z�v�� �������}V����)�LR8��{�����i��[�����`}������|:zc�;d^�N;p�a��l�z�u&K��!�Â�κ��y���nO ���s@�_U�U�^�yz��>m�	��Is4��[�3���I(J�@=Θ�z��|0;�ڣq(�4��@��� ���}��ES��Zu�~��'Z,����ʺ��`zs���|03+zXlDOWs��γbY�4��@��M�_U�U�^�y�@��I'�~n)��z��MLy�G/I��s����Y6[�v��i�QqB�2a��b$j	�h�������m���h��̙&!HG"�*�@=�٠_l���ՠv.]�!9��ؤqH��m���l��>\(� ��Ax s;��h+~z��������9��<�S@�]�@��^�{z�����M(�2B'3@�]�@��^�^�4-���߃�ĢX�Nx�7��(�]���s�nUc�e6-����˫E`��,'�D�nE�r�@/�f��s@���@�����X�@N28���5�LL�7��Zu�urW�""��+���i,�di6(��>�O����������;��\" ��;�5v07+zX;�Lݽl*��	��"EL��/Po���I;��_�
6LB��E�Uֽ ������;��h����Y$�[�H��u�X.h�����4\�����5�m<�	�c�
G�@<�٠Z���_U�Umz����򡀇"����x�~�ӭRJ���f�n���#��!$Z���@����m�Vנ^g,���9���Z���@>��@T��ﯕh{��Lb��q�Ǡ�l�*���̮�`t�u0-4�a�)JH�*D+$}B�@"# z�708B�H@$da$HE�#[`��!	!�HAT,\��;a�8JB�xe^�Z�<�aBHA� �H�3	���Y��ZK��fi�
�-`�Oߺb'�U?$Jd��+,�i �q�		��C���aB0�W��0�!	��8R$� �O)�����$HD�@�ŌF2H�F2�0"B0gc$�bB�X����rC�����ԫ�mn�u�t��#��<r����� �cy��IQ��ƨ؏Yv^gn�aM�u�[�v-T�p�`�B��3�[�i�����j!ޠ뫭����W��T�����f�A�:����
٭ڪ��1��7Zn�OJf5�i]õ������ng:ë��=�0�Kb�J��Ha���S�����[�2�Z��Fz�������ԫ�Vˠ|��X8�AT�ɷi��b<s�-�����اp3�/)v�����-����g���[]�Y$��t��X�/3`�/.��oG6��|�#H�3�c��9�<a�C�;(�ܽ�!�j�UV��� �5x��Lc�4Q�f�s��8g��8U��l�e��]�:��-n�A�X�&���wO#�M�*�\V;Gm�-���iey��1�v:.was��a����e#i*;[nx9&8��9�v����ԣ�2CrZ�m��%fm�UT��v�����v�r].�($ơ�S����)���T��9�Z��<��5��q�͜�ST��:q38ϡlv�Nt�pmi:�5���8�H]�f�-�\�oXs�\�u�)AŸ-ˍ�F{*a�p[n�E^)l�v��C�1�s���d�7cv�ڷ���+���dm��:)�S��8x;*,2�:<m�5^V�VVG\���]5����z��v��V�M[d5�6��I�-!>����m��*�Xݝud1�Q�U��3�e^� ����eSa.�r�"�����%d��ܺd��$ΚX��F��a!�c���㫃���wA�v͜��ƀ�u��یg*l��R��2���E�랍�pd�k/M�x$�#�v�,��1qnSB�lR�Lj{�T�C�����ήy�p��s�p��mć���*��	Z㶪���B�h��;S`��s�2�.p�-Խt�{�q�μ��PD9\��_�b�m�:f�S:�!�]eθb�ٹ�t�	���^�:���0Bx��!�AB�U^���z��z�D�v���d��0ٻ�r�g@)��u�s��I�ܐֹ�ev�WlŽ�����I�c��qm-�q�֭�n�57%�ۖ9I�vV���J��r���N���]���.+se䱛�1����qT���8��ݝ�R�b�N��:=��4��C�l)��;#݅2g�&M�B���Sq�KnR8�r�!�Ol\ڄ�I�A5ZfY+�gn�{��;��]a>��21֮�Fݻ4�n�;מƍ<�b�h�z�z�^k6��9�9e�d�<]����ZVנ�l�=�p�&)��y�@��j�*�@=�٠U�@�܂�"Dl��!�@��z�������Z��]��c���)R= ��f�WZ�}v��Wֽ���كyQ�9rhu�@���hwW�{l�<���ߛ�S�r�-;O-���˃\^-�v��>Nbl�G�Ήt7jKrH�BM#;@8�}}V�Wuz��4
����q�VUJ�UU�w,�ާ�
az!%s�`zs����,j� �����#�@<�f�yڴ��Z]k�<�w[IA��	�94�S@���@��z��4sޕ��1�~�ǃ��;��hu�@<�f�z�huS��Xّ̑�<{N�#�x<�{u�lL�7dlhL��㞭����&!HG"�*�^�yz�����g�/;��=����
D�����#�/Y�^��z������ˍ���r&��/YM�}V�2��X�US-����$����I=�[����,2�,�����s13݉ր�7z���h���pl�cnE�Uֽ ��f�WZ�}}V��?��ۮ�',�B8����tk��Q����8L����]����Kt�݆$ϭ�tǠ{l�*�^�ﯪ�*�^��.�ڬiD� &D��*�^���f~H�w�|��= ��f��/z�Q��f(�xԏ@���hu�O�=ﾚ����<���@��Bp�E�Uֽ �w[�{��ĥ0��	N�b�r�)"ƈ�R= ��f�WZ��z�����Y��'�)������΍�m��˻q!֦�ۣ�1̘#;��g��X(ɍ���	�''�|��=��@��Z��4�.M�&0�c$����u|��&�jۭ �h
�+߳�GZO�'��9���@���Z}�4
�נU�W�y��`�I����q8���hu�@��W����]���wg��ڌiD� ,�I�r�^��ޯ@��V�yz��(��I�;�8�A{tVؖvN̛IqN����r���ly�+iɳ����l� ����3��2�݅��-�3I������]��!zŚ��&��N��n��+��,���A����=�sq���`S�Nz���vݠ'�c�H/:5,[y��^z��l�`��Ǟv�s t��:}gN���:����]���tw��]U���Z�A=�I���c].M�n��k`�i��K�3�h��]v��ܘ��Νũ�S�H	�q�R? ���@��M ���s�h�+�"M������yz��)�r����qUs蒑�DH�!��~��S@��W�[e4����N$��q���-��/z��)�^�@�Qؖ;0Y#�I!�r���-����4l���~����C���H�c�ɍI1���a�'N�3�U�4���7����7^���,s#r)�}���@=�f�m��9{k�<�_�u7��0N8�4��y��:��I/s���yw���V���i��(�p�cRM�j�9{k�*�� ��f��z�(�df(�y#�@�{��[^�y�@�ڴ��W6(�D'$zVנ{l�-v���W�yyLx��&O�*`f�E�)��{k��ڞ9���%��yn�۴]@Rvz51O�m��٠Z�Z�ޯ@�������&&$�i�4]�@;޳@�����h�;�b��$��hf��:{��jn"�P�DA
�v��<��hۓ�^D�9���@�����h�V��ޯ@��TuA�4�#�@<�f�m��9{��[^����ΡH5�$�5p��#d�"����d�����l��^n:����t�n,�I�[e4^�zVנ^�@�=�V�m�Oѧ&H��9{��bEV���4]��~;�"@BpRG�uv� ����ՠ�Y�y��e�)DH�!�^�@���no[�IDMN����\�B"	4ܚ��h����)�^�@<��d?92AdD����\\���m�:ճ���o�&����c�쎮k+����r!)2B) ���@��M ��~���f��v:�*/#.��̽��4��h[w4^�z^�@�Zx�ӊ7 ��f��s@�{���)�{�;[y�`�c�F���NwS6���go[֪ҍ�)�Ȇ�h�������hu����2��u�&A�8�9���g/���]����b���<s�3B� -�+��6�:��d��v�5��	�q�A��2�l��<���;M��Vpg����P�b��l�'k9������k4i�<��J�['9�5ێ�yk?ȵ��s���3�lb�[����c;���;h���;c3��;�>/G6تn
��Pꎱ�w�h�F���3��\�BS�v����{���ݺ�cl�l;&�+Z�b$�V�˺��[,Y؋���Tt�؋��*^ܒ�VM���]����`{{���(Q�*�zت��IL�	I�H���hu��/mz����q�&�i94:����W�{Ϫ�/Y�\W��yf%"�Is4^�z��Z��4����a��I�HF��@���@<�f��۹��Y�r2�GŎad�ɒc�u�9�A�!F{(c�r�=mw��fV�fq��Ø~��Ӌ@<�f��۹�r���=���=��c���m("�h�"i�J8�)������I;�ڴ��oߒ;�}��o��8�7�{�`gV��v��7;�`ftM�X���=�����s@�m��9{�����bjFL�H�����06sz�=�L�i��np']6�Oۉ�֫���h�\���i���wN���˥�n���]���06sz�=�Lv�LS�0yQ�$i��9{�����^��{n��0�v&�HF��@���`{��e)P��Q�
�L(��B0��HB�@�P$$d/r��t�%�Hd_� ��e$��H+�I0cB!		B҅B��"�0"E���t�~���p�B	䟂��d�+F�#�%�`!0#�����fL�D�*`��e�� �!	YHU�(6��HJ��`H�đ�)A��1H����Q�ASPo���8�x�G9Ǟ���1UG�t�DA⪥���4�7������UWMR��&j쪺`{��`nw4����`gV��3)*y#Q�M��I�{n��ޭ��[���w4��!}���E*�Jθ��l��5�yܕ�������Q�[!����Eӂ�2ao��8�73�9u��׽,����0;:'�e�қ&TՓwt�έ�`fw4���i������]����"�)�h{n��۹�z���k���G�C#�%�ݦ(P�����g{�`gV���I��T )*H�HX"�R*�D0����$��1��Yd$i��9{��w��� ����;�w4��vdi��,A����Zֈ����2��٫��燎sv7�R%h�(��D��"n5#�=���/Y�w��h�����cu7���'%��h��5�L�P���W'z˱�bGw��<���q��)&�{�4��^�"f"���h�<�E�(	Ħd�<M��9{��ޔ�/Y�w��h�+�#O#ı8��h�|0=��07;�`����B�$'��������r�s,$͛h�[�g�M�r�o$m��p�)�66�'n���v�$������3�1Ւ&��9�p��]���ͱť7�u�m�� �6�V�"�[���"�n��=?�:죾��g�N�W ׵�oVL�.�D^ش�ن5����[/�󺼆-�D.Cu�M��\n�vm�[��ͭv�s���<��.�Rv�vR�u�L�iBJ�f�{����ݤ�yr��t����t^�m����<RF���B�t뛢1��)��Kvx߾i���� �޶v�ނ��y$Y ���w��h{�h��h^���^�<U�C$j�06sz�=�Lv�L��ۑB�ʹ��3.�.�/C�135�ӽ��4���i������\�Q�Jj�%9��<�w4�����^��^�������Gc�4cV8ً���۝�I��:dXX]<=]/5�T�U��/*Y�WUv���i�fo['����7�@����bS1�&�h�����
�
�ޖ���sLi�Nf%1ǍbpRG�{_U�y�]���s@�{����b#��9�h8����?Ѡ.oc@�]����%q��dxd����s@�wW�{_U�wY�{��VnF�H�"%<V�+T�5�Z���Jy|봖��-`m�Q��B�Dj4�hwJh��h��}��}��}�#>r'�	26ܕ�h+�Z�"&&�>I怹���vvs�Em�����nS3knn�ͼ�L�����3���H H����A1G�B0!$�H��`�� �`)1P��B5%���論�=�,�(��DNM�f+�}�hl��=���<�w4���Dd�0jB��7o�moKۼ����������u���)��{7��br��[��f���L�:7�8z�z�p�����f���]��=��07;�`{v�`f�&��.��U�Wuwr���4���"&E��h%��>Wʵ��L�P�]	�H G3@�����t��~��+~z����Z��M��A���۷�'w��{w���" J�(�Գ��ѫw4�Der'�	26܊C@�wW�wY�y��hwJh�v�Gq�;	q0v���\=�۪�x�؁M�-S#l�c�'sI-Ӹ�nX^x�?lwY�y��hwJh���1^I�E6�h�I�y��hwJh�����4̷ �ǋ#2B9���F��w+���L�Q�O4�{\*�cf'k������뱠~�4��L��k4vP��y��AWuwr���4������/�������g$����a	�����M�Á�l�
V�g�kf��X�v�s��t��vVۿ��^��\�'e�=�l��z܍�0��,��]eq�\��-Ne�ֶ/:��BCd��r�at�N:[����;k��"A�^�ݱX���Wbm*3z+�苴�9�8u)��/.�8�	�W�����|�r�.�O&x��6���q�}�lxy1��]�7k�0˻uڥDg9}\������rW��]��n�0ƱLvFً�v�:�:v..H��4l�Yk%"#Ƈ&G�H̠}�����O�k?�,c�����$�4���\>b#Y��y�)�~ďzύ�~��<�����"����I���Rf�۽lf�Ln�S�eu7���N8䆀y�f��w4;�4=�M�W�t"�mA�%����i���`{6�`��`fr��7/��y�Tm�&(�<�Y��O�	z�';@.;r��CK��Iv���t�}!��`{v�`��`{w�`r�w1J�n�����X�ާ��P�U^��37�`{kz_�D)�>�N_Z�����9�h��4;���>�@�wW�Z�\X���(�)&��u��?u��w+�s333_$�F��j�ľb#Y��yϪ�<]��wV���D(�;��>��!W5R]^�:�^^{�us�^���N.-��3�K��]^�
dm�#��=V��;���u������{����D�O ӎ)%0=�j�y���[�����0<�:GLq4�4��hw]��}V���
��B����遝�����L�b?BF�&hs�uz��cA����?Ѡ7'�e�Y�^y�����0>�Q	Nw�_���`f���-���+�qLc2F`�$9����N�3�<<�nz\���3kupf����H�ζh{�s@�wW�y�Jh���7��E�4ܚ����9w+�?}؍ ���s3T8V���*���##s4
���{Қ�h{�s@��Y\$��q���(�=����o4��	E��IRM%�m�����gѤ�y�q� ��[ټ�gw�������S�J���/fk��8+����n.�eMS�*�C0`�18��#�cDnM�z�h]���v!���D��>m�ݷ,�"~��
L�9wW�bG�ύ �ﾚ��s@��[�1I��H'#�<��-�@��h���/��b���	I��-�@��hwY�y�)�Z�V?�c�",���=��0��`{v�`��`z%B{� F(�Q��$�! Đ��	<�Qh:�!!��F ���b�B�a?o�w����_I��4<�M�Si�b
�R�6�6BR�(  ~6�AO�*B�T�� ��E
��P!  �H��`���k�����p�b�$�J�
F�����"K+�/�H��S+�G	��]dY]!ʒ���$��@�]�3��18!�+�%�x@b,I"�c2� ��c����7��^��NwW\�t����з�9�/�SQ`�<R���W<�U�����v]�ҭu�\^�.kD�Hݷ���l��E�'o7��B�U[nE+$�R�h8����F�5�|�c��"��/�(�*BӥxA�i��A��4e�W%�x��ʦ�D��&�z5ԭ�n�%H�G9JV�
�m�$���չ�n���q2�;�mG�am&����brRl�ȁ�ϑ��2;�:��i6^I+�j�v�^T#�H��k48��Y�6�vKLlζ��؎��:�+�uLv�'.�!�gk'Goi	��)yŁcR�{�o�N�MT�V�TɹȲAZ܎�h�n��ݜS��{{h�����E6 N�9��6:wj�:z�a���7k�g��{r��V�\��l����<Yӡ�)$���޺9i��ϳٌ�kL�xyvp8��g4�U�]WG��c�7��vv892�� m<YCe�[����(�d;a;��5]�cZz���x2=]A����p�[#�3����Fs�#��gF�����&9��մ��scsF����3r�p�M��sm˅�#e��d4�fwC�F�V$�C�IciFK��F��c.M��ڸ�.ml)���e9�m֡�u���͝�*�ф� �cYq����	��n�ɲNz��ұ�Ƭq.\��=U���ώ�J�3es�&��@�<�ij�줹�헡h���)�U�4'n1-� ��t��*��7:�'�<�1r���#I�L� @��k��zv"qj�4�n�,Q�*�u�0F��.3�k"gm�U�:6.kȄ�����2E<�rk�*�]�	���6L�s�nX���ˮ�7Z�75����Vd��V�J�	:Lv��;8J�/�ck	�tcY�u*9��ѻ^�6�m�t�ԋh�,Y;>K�]�i< ��@��pJ8@��pܵ�*lR��T�<�}��|�E�����h�u�w7/;��],�'��CD��Tj�~8𢈱uL��� ��aD'��M��Z���VLͩ�,� ��w5�Wg�{pW1����i�k�����뭝���j�㞩�,���;���!�u�F�;���6�h��-�ԧdS�S��,�.�F���-�� \���o9vj�[M�dk&5aOmr>�v�����>�����w\�MU壠��rf��Lh����?x�{���d6�f5�ⱝSm#u�%�dn�������۱{�u��8�#̩����ʦ�g�~��v�zނ"���2LyCI��#"s8�~��Қ�hu��/R�yT#��drG�{�)�[f��[��r��/1b�щ��q�$4��h�-���*Iށ�c4����X�4,���@���9wW�{�)�^�@��Ė%1���D��06sz��|0v��=��0����ʡ;S���7bBn��F�^�{fN�Fc-��1һb,':s/7Xu������� �o[3���oSV��/e.n�-��svrI<��u ��PP�DBUa7|�g7������B�}��>c��8�"�rM��4^�z��M ����|��U�L�%5i��������{���В�S���f�Z,��@�L��G$z��M ����۹�r���*2�H��M��j�i�*�ts���T�y�a!gm{nom�[�dIb��o����/Y�{;�`���IB���_������4,���@��w7�ٙ�"��=�ύ ���W��B����$H�i���������D)�BS
"R��(Jɿ}�`n}�L.��V*���욻�f�ݽlgsLsz�;�a$OR4�4��h��ù���l;�]BథgC������wWb���۶[Y��N�k<u��cJ�$��#!c�b�Hےh{n�W�^��)�^�@������4A��9�/z��#�ύ ����<��� �s���$m�I&��)�޳@��w4��h�ĳ���7�.��0�sO���oc@U�+�Ʌ��kၘ-�E�U�R�J.��{n�Wuz����_m��?=���q�v捐��j̱c��x��Q`Q�b:y5�H�uv+ b�t���탷z��|0��`{;�`f����Uȩs5wl;СL���[;�4��h;�R��oR4�4�������U���c4lbX�ȱC$i�4=�s@;޳@��S@�^�@�p�u���22'3@;޳@��S@�^�@���/{�����/~4�6��xqv�B��i�4v+���J�Gn%�S��:zW
��ce�<l��Z�F�ʐ���1�ʯ�,Y�g��ۭ�܁¹��@���:�y�6��ʙN�`��8Ɏ�t<�VE^1(���vg*�i��n"v���/<n+�v��y����R�s��a:��C%�q�D��:'/#k�V�N��=qVb48$������{���mg��Eݸ��z����Dta{����u��÷q^�5�R�d��+��Ԯ*������v�^�huWs@/[4oK,hm '$nm��?g�H��������b5���LU"0̊�̒Ș�nM���s@-�hzS@-�hwQ$�?,���D�h���b4rY��"fbb�N����8�1�?<$I�4�)����U���� ���V
4�F����"���t��}�Kkcql����k�H���UsG���x�oR4�4��@�ڮ�^�h��-w��X��7����N�
&C����|0��`e擱���22$�h�f���M���EP�y�}Ξƀ�URWW�@�F��M���m�@�ڮ�[l�=�D�$m0y9p�:ձ�9�c��o4�b4�����\�F�]lፄ8�)r�M7C�)�e������qͻ �8Xu������I��[�,�;��ocL�P�ϱ4
b	�(%�f�_��h����`fq�02s��)�B��]�Wt����ow[2�H�P�
�	B�P���*s�i�oo[лH�1%#NC@;�����h�٠w�S@�����"A	%�3�i�gw[s����lY������n[��N8.-��w�V�/!��.��6����-`m�ԣO<�Θ3@=�� ��hu�@�iw4=�`�(�ƣjG&�u�4�٠w����h�}�RF�ƈ	̑ɠ������m�@:���cꢘ7"��5��4>��{��3@9��˖htD���b.b&f�I��?��7�}��}��r��,�]��Nf�u�h���[f��]�����H�4�F6I0X6�\�;�c�s
�2�
Z@x�ާsh�깞�w\'^0�'$�9{k����j���٠{���豩1�)r= �l�?|�lh$�@��+�31T*U(�k��I�{�)�m���4��h�&��6A��) �h|�h���s13���h�L_A����mH���٠u�s@��Z�٠{���<Z&�x J�j�7P�l�\�xP ������I�M�(hvvѫL��p5vRC��n�I����lu��>e�sзj���;[n<Ě��ض]��4r���.AP� ��?_gj�U���m��۷m�7B����x:���P=j�-��چ���[qˋq��4c��bl:^�ɉ#�aw�X:{b槵�iȽ�S
��7f���b�n6uӔ��Hd.z�Z�h��Y�Gh�,�[�t�Ơ��A��U��U�y�����>�e*�Ig�?P��h��H��#�i�&h�b�@:�4^����h��ؔ��)%�E�u�h���u�y�I����Kۓ�_�O�	rO<I*�V�$��l�Ē=uW5$��l�Ē�u6bƤ�4�q�֤�]m�x�G��椒]m�x�U��jI'��x뎿�7�/�=.3�j�Z���K�J8熶VK��44mrYn��h.[<�mj�l�I!}�q$�����$�$���3�H���4��NF���Iu�y��tb%U�9���ݼ����[Q몹�$����Bƣb�I�$�K���o��$z�jI%���$�{�������-I%��3�H��\ԒK���I^�-I%�:�'$��cNO<I#�UsRIe�}��Ԓ���Z�Iu�y�Iܯ,�0b���`{O5\M�/;��t���v P$6�2桎\F���&� �?����IWҵ�$�[gٞ��G?��jI.�.i��B~X8'#�Ē��kRI.��<I#�UsRIs��<I.�Qsf&)2)r5�!.��<I%�ɩy�Qm�°'�\6� ��̮˔%�$<�ܔ��P�L��:X�Oƒ"�KJ�./!$���Za?~���XF��p=�9�!���$!a��~?z�Ĕ����̚C,�/ �0`�u�K1�F��	$	DX�c��i,b��	Ȥ�b�)�E�u����sGyLc ��� �~� B@�� 4.OR���z���)����5��<b�'�$ehR1�3"��6��{�0�*�Oʶ!T�%��M�z�p��A��xNO߉e��]9��x������!����0BM����as32�%�)i*�dV��L�1�D=ˁ*@�������P<? �Q��P� z"��u�F��A�A4|@���bJwt�Ē�t�Ԓ\�K���)�$c�y�K��}�RI+��O<I*���[~�������K��f}t�2h��95$��l�Ē-���Iu�y�I/]�MI$�=ŝ�h�0� -�����j�j�G'I���h�{r���\ѫ[6G�d	�F�$��H�RjI%���$�v�>��}��Ēg�`��bP���K��g�$����Ԓ\��H�Roʹ��K򑉹a��93�Is�}&���-^x�E�I�$���y�I^w^,H��"E�dqI5L��wKݷ�{��Q�"!o�Q1L���Y��g��'~>w�p���q'$�-�M�����f�u�h~����*�x���4�&���a��인��,�m����Ϧ�=:�Cs9��mbd���d�H�<��ۚ��f�rK��G��3@T*��*�(�̼����?RV�\L��EP&�h�f�u�h[��v6��22F��9[^�oJh[f��٠�*�x�0��l�H�zS@:�4�������`�ŎbP��If������,��F�31' �����`z�c,����<&���;o.�[r�ܮ���]�`V��A5�1�O1ЖL���%y�x��묣�K�n��5��M����u� ���.��p�6�2�m�qλ$�4�v;Ξ���5��^\W.Rŗr�Q흥���n��������	��Nj�q��9w=��+�N`�Wp7j%3)�]�Mp�1���i�vz�����(߯�s:�\�5N�qdNl�'���یl�# 7nV�!a�Y�7S��C�r5���~����`�l�-�M �l�;�u�)�"!�qɠm��)�m���f�bG}p>�3Q��Q'$�>�ύ �l�<V�4��@�-E͘���9#�����m�@�mz�S@�r]��19��9��<V�4Vנ[e4��@3���vrA��wri��������b��}�ݧq��q���9�ۦ��mF���I/�}4zS@:�4����b�;�K&�w3sss�N���砪~���X�;�@�Z��9[^�g�K-�6�q
��٠x�vh��@��48��H�dF4��<V�4Vנ[Қ�l�<�ia$�ɠ{]�@��4�٠x�vhٙ�>��#0�j2�#n�t�N��k�}�y	�;L\dN7ظ����B3Q��PnE�}gƀw[4����Z�j.l�Ԑd����w[4����Z�)�����iv+�s�ds�h+]�OwS9��J<�$��J�k��`oo5�nv��� ���@�[^�oJh��h+]���
�$���yyyz]���DRm��>������.���̂X�ɓ�Fd�e8���6�/.w&¼ΌN����gA+����1�)�Hh[f��٠m��)�y�ꤒE1L�,�I�x�vh��@��4��@��bXV��N(ܚ+k�-�M �l�<V�4o~.��f<����`ow4���u���")H	X���0!+!$�������ꚫmށ�·�FfFD�rG!�u�s@�[d�9[^�m��?�9��}�@Y�<�&/�)�w�k==�c���Ê;��ֻr��FN.���<]�k���������:�W�$�&b|A~��� Ͼ˃�ϒL�#$rM �l�-v������&���33=�p��ndM�n8��>����:۱�������*mށ��EE#���Jcr- �l�<V�4VנZ�Z�>�I$Sb#�#�h+]�Wj�-}V�u�h;3?a���R�jq����
��⓱�A�Y�g���s$v���!5��ǜ�;=�덃�&m��[1we��gvm�bp8�Hi�N����7v�b�d�<.�i�@����;7��W��c�vs�]fMLk=����*X��=�{[�:��=S������܂v�Y3�k{;l����m�1<Cri�;N��[��<USz-���|U�Lr�Sr�J��F.�r��Y����nf&�ģ���;��q������I��\�*'V�1,#Dd�'nO ���-��h[f��٠{{�t�Y	�x(7"�-�M �l�<V�4Vנ{��sb2I<��h[f��٠r��ޔ�;9��$1�9��<V�4��@��4��@2��6T� �jF��m��)�[n��٠y�p.�ŉ��\kb���Q�jѐ<Ҳ��K�8p;�Nŀ�T�I��7 ��M��@��4R��?RV�������
fUe�e�n����N����qQ�O�����M ���@��4(��$��Fb�,nI�x�vh���Jh����İ�`O�$�Q�4�f�ץ4�f�����=�tɌ��<M�4zS@-�h+l�m�@���:~���ď�k�iL�ԾM��9���z�Ì4��x�����Vz�=F颃��$�����x��h���j�.s��^�<p�B94�M�k�-v� �٠nv*I�q5#�h[^�k�h��߿~ΟDD�z���S癠}�p�E�eQu�6��@��Z��h.�� �٠z��*D�k"bS�h���֩^�.K4��h�����S?]�^s��mے���y�]��zB�ݍM���['<ѷbd ��\��߉���zz٠Z�������IaX����7Q��f�oJh�f�}uW�u�˦Ld" �rMޔ�����@/[4r�nQ����y�y�������t�I�{��D[h"�@h	A��B  ����B@%U,Em%IJƧ�M�I1��f���S�paq��^Aw3@����*�^�oJh���=������V����nZ�%��g����f7���9U���n;0ܖZ��tu�ɠ9�����h	v#@;��LL~�}n��Z>c�$5"i�$��)�~H-��|��@/[4{D�����LrC@/[4
�����@��hQ�Rd$&��L�I�UmǠ���S@�n��|�XV<#"򠫺���rY�S�����|_i�Oo����'���D�*+��

���D����������

�����T@W�� �E b�P*�A�P(E�EA �Q@!P�=QE�

���(*+�*+AAQ_ PTW��AQ_�E���PTW�AAQ_�

��E�1AY&SY�!��,TـpP��3'� av�  (��Q ����   �(�@e� 
4  �
$ \x �UH�� ��@�@("�����$R"�R�P��R��R  �T$*�B��QA   �     � � kO{�\��׷�wf��|��c���G����>_K޷��f����������p{��^��  Gy���w��1�����X��[����<�{�����w>G�܏���� � >�%  
�h �>�vp��m*�,>�>�{�J����C��E����w2��ܪ7w>��}��� ��Q.YT���>��������U粞��x�� }�o���\���\���>�  |  >�   ���R�T����+�.���>���K� }+ϟ-�u��wu���ұ��>����)�=�J�۩@Bݺ�J�jU)�u*�r�U)�R�VZ�@� h P     
 
 
 v��Jsj
W��Vf�J   0�      b���C��U3����Z�MR�� ���:�;�(b�1iUL XuB�R��  m]��.���O�x|����9e�.`�7� p7��{�����zr���o  >�� ( 1� ��C&�������� u�zWG]���ǈn���=�Ӄ_qz��� �<��/�Ͼ���g�	{����L��k����x`Z}�6o{��{�y�}�w���IR�	� "~�
JR   ���R�'�( �'�T�i$�
����ڕ%T�F��!�)"#@�>�O�����X���������{p��{=����'���`QTW��$�� ����PT�pQTW����������*
���8?��H0ѳ?���f���}����f�1ѳ���?Nh����Bp4o8xz�f�������N���>W�zپy���H1�m�����$�kxx���06�<�p��#Ѱ�FH1��N��3��o����,���f���O���i�p��ÞC&2b�8�w�<��Ϗ}8�a�2+y��bF�`Y�4ٯ�4F��Ē���C���6�r�0ٲ1�;vFH3V��oA�L�$F���3D`i�0���ʳAc�F�f�d�	�(�P�"qQ�Ó�A)˲	l�3F�f����f-��מ�����,4G����h4XdD%�q���1j9lك㱐�I'dăLa�(�l�4X�b�l�h��|�#5��c��&,��i,р�&�v�k{LM4y��f��p�������hۧ���Z�\��39�B{��*T8J��p���@�m�+�J�E@\��@�B��d(,pz��a���8xg�j���i��^�.eД4���QP*�Jb*�)l��'���\�]����FYH<D�����-����KA�`C2A8C2\4F1�d0�Ju��RHH`h8�`P�qf#8�vsC(c�4��>�no�q��h��f�4p2�M�Ȉ"6�Z1�`���1�h��5f�ϼr��M�kWhp�h� ���,�!aJ�HFi7�Z>-�,c�Š)�Ř�0ZH��5�h0����F!9����\�y2A�'<�W^�uC�U����߻��~X  b�V9cĔ��m����RbP���ՎУI�l>U��n��|-]v��!-��jӕB�!��F��F��� �@�`��}W�A���m�_�)����c���H-o��t���.�@��K谈A8 �|-]Wh�F��ڢ�p
��`��[2�ØW��Ē9�l=R1�9��ס��0��o����9�c�Bt
T�8M�ڀ�����We�V
b����. m��Qパ�,�-�l}}gF��>$F�s��r��h�Tn�a_AN����
�]�m���)���ŮxdYk[�,4p��q�l��I�r3[�\=l�~s��X'-�WE\vXVi2ti1��Fi�cXm�վk�s��9���Z1����7=p��3F||�0淖g����g9��)뿬��:��NA�"�vC��c�h$��>#4�|/^$eMV�֎�"���y�
y�P��'9f��������X�G�xkf��X3F��f��ᤃ0�40a�p`�N�L����oa���c[�1,��c0�F��0�F	�La��'�xp�&hMC�)"b� �dŃA���L+�('	&��`�L�6D�m4�$�0e�F�>$����&(�`�0`iG� $�� �% %	RJ�RD��	!8� �	&Xp�d��PC�.�ۢ�� !~#F�	04��A����8D��4l�ɳA8i�K��1�*BI�o`�ѷ�N�HI��5��q��4F��A��u�|
��(�Xjs[�4h#5�4o|0`jb��5�Pa��͜J ��F�0Ө1Ѩ��p`��5�mf4i,Ѡ�+8oq�ca��F8N�h#Fͱ�K&&�l�9�c6[�h�q�e�h,�[��c8��HF�A:��FRE�oތ��q�֩�m�X���mщ�0֖�DQ��u���u���)�PL\��E�$Vh��(Z6h�s��VK
Mk��a�;�x���9y����R� ��xm&=	*'5�qڱ����<<8A���7����3[8�xl=I�X�������{�x���l�F��=�֋`�O�Fv�y�l�����C'E1�  �v��!�AD!p�gJ4�͜3{L�pM�6ca���0u�'�&�1�lpM hd�40ZϏ��'��>�6@���[�<r2��[9Jy��e��m8��L!��04Pm�C)'5���$�� �`U��wur���^1�<���7���G�#��z�Ǆ�"n3����O�M���Q��i,*����I����	����$+l4<K;Ki,���rLe��xFiѲp<��/����|�4������
l�N�[�B�1��z3*�[���?I�v4� �L��@q�	���8��v�\�����2�Nz٨��i��4�m���#c8Xh�!06�h�!8'4Xh��pѶ�Ę�c�a��y�ki����٫4�h�Da�,58�Z�M������3 עD�0z!"2��;��JsKK�DVkk��8f��yz�a��l��f�Č6�ko�������}��<9��
c3Z�N��2�,�f��F��0�j�fjѦq�٬զ��ՅF�A?�!�C@NbAg�Zti1�)���?,�F`A�G���Y��v
�:&[`��
� v� �@9w�	�,p;�v��$6��Y�&��$�e�p��������@��*���z�U]�G���k�ـJI	1��<�,w�p��&�����bFb��S G,>��T�� ��|�Tt�T����Pjv$��c�.�P�|]  BT��I�@��)�
v�M ��D�]UA�Hy�	��a�L4�k1,t;u羚#-F��|3|疈���!��#��QﮞzAY�6q�[���Xj�f���fr<|�6�@Y�VjČ�Rp��x\5�k��\4G��٫=���C�<�#F�M�vFx�M/Q�Y�1�ߍ���$�	���Ab�&Г�A�^h��p-s0���!6k~^h���5 70�
	xU�?&� i�����xMa`Xi1���=S��Y���o�����D�ϼ��}���Č^�p!#gǠN6o	�Zu69�k{���f�T�d%!�tF1H�p!�qc ��[4f����`n��R�4X*7%QS��T8+�QB`��g&|k��Np��\�f����|���<�� �1t�N`$�I,�Xh�F�,�ff��e������sI3M��f��a�K�qx�����1xI���}V�Pcn2�
(AQ;}�zl[6o��P}!1F��9V�`�����`'�
���� �0
��Ф;lb��� ;�p:"x���y:pe ����
��q�Y�E����	 �5�FxY��,�~������M�;���4����4F�Y��03[l
ٱ�M�];fpѱ���bf��N2���t�$�8d[8�_{����f*�TT���[^�����*� jXf������y�|���z��o�{�fY���sGƘn1���������+�N
"��3c����F���Z�\,4i�ּ����qtp�����06h�3Z�s�|���������[׉���3�S���L,�Ef�����i�祆���繜��y���y��&:�sßY��b`Ŝ�N�0��� �#i�$0I����.��R���C�q]#!(x�4:vs�zz�70�Đ$<HORAƉ)pI`p)�H@��� bLt;^X����A��u$,�b���	�#& �`���8�4J��@C8����jc6Xm8HrW3I��WF��c8A�y�'�o��p�8�I�hs�|w��D�'S����f���g�h���,<,�S���t�:QKM�@ �� ���%�ՠ��hr�����'(jH����� C�DS�i�W�Ȼ����p��O��<����:��Xˬ%��7�y���.�cg�q���'Q�ꆪ}q��/ɕu��D�q	OT����Q7$)�Y�L\W�k­���Z�K�#v���j�߮����H��U��@�S8%������$ �|US;�\b�����Bw*�9���dE����XD�v[2^R�r��t����`�q�5C*¦��Y	X%�S��9}�����컺m���8.��@�Dc��R�;R>O���EWfd'w.�)����� �#�mD*&e5u�NVz�"t8��E��jTE�^���xҬ*�/"Ⱥ�"��J��Zw9��SXLA���VF�"��B�PW9,�����cSg����U�=1P*��w����"n�n�us�lRԨ��j.	P]��F9��mx����)]�!���ʉ��sJ��uz��V�	ʯ
��Zsn`��W��-7wSؾ��J���k�S�W��j&g�L&�w�M�
��+f�wM����)wɰ��s��"-p��B����I$��`  Hp        � [��g7i{Y����T�]w;��T1���{D�F��s�w(��J�!������yl���+�5n�š.�����7&�]@�DT�]�]n���r�p����cg-�-�W�N�늗�p�8I���[m�	�܇[ѬZE݆�g��ki�bpvc
v{$Y�n���Q�@c
��(>I.���GYk��x;b��nzι-���>:J�B�@od����]��-Ԗ��"���/m�`��ɝ�n�˞[�mEQ̼v�=��&v�vB�{MdI��\8 ֧N���k{GN�Zew4���\u�lY+��gQ�Ӎ&�-�n����+$�<����{g&ѷbs��*mf0�r;i֎Ӳ��y�;��N��V������m��6�si1��l��Y���T����P��r�<�%�P+f��[@���V��<�����͇.7lC��(�Tl�3�W@�j^z�-utQ�MT�W@f��X*��^���o;c���׮5�;[R\a �(�e��� �nWf	��ZtU�p����u�l�6�@o���ψ�� +�R��R��sF��m��	z+gevZRkA�q�Wm�G\3ҽ/jt����;v��\��A9v�۶Ѻ5-��6L�.ʻ5\9A�����n�u�����se����+�ͯ`/��K������0����7��.��m���E]P��#�^Whn�K�YoX��Ӱuu��ݞ>U]��ZN��ث��)v����i�6}��Z8��{lSYUm�m  mm��ZKd��〓Z� 7^r�]9f�p.��S����f;{jj��X�D��۵�Hm-��z�v�q:i6�I�Vwjv۵�z.�iY���Y\t�ј�j'�Vۛm��0"@�u�o\m�� [@k��n�ERz�dj�3����v���!*\�La�EP2�R��q�R�T�khi��l�z۫Ul�H ���m��M>�>�  Hm���h�$	m�� �5�ʾ�[p�t��@hd� ڶp���e�1b�m�l�����m-��,���3�VvѶ���D��a�7d���Ӏhm��m�[@ ��}��|�`$�B��` ���?�A#E�8ݵu�ŲS�m��m��I!�r�n���#��Ͷ@�����@[y�� 6�n  
���ݪX(�
���,۱�]dV�Pٗ�v��̀[v��m g[{b{i]�ô�U����(����"�nv��:K��[gm,
�s�̥紛�H�g$����	Ӛ�hM��	m�    ��6-�@�  �hH �H 8  �8lְ m  ��� A���  @��Է��A�қU@�d:_i��"Lpڗ�s� m�k�  k�V���^)��BR���  $$m��l     86UX�U����������0^���R��@�n Im,�����6�\����C��2ѻN�������;��g�T Y
��P�q�*�� �l��� 	 �  �����l�a��m$6��  m� m�    l   m� [@(  �f�h  ���6͚���[,�UM��� �[���8���o�|�6� [%�-��ke� h��  ��h��l ���i8I�*d�,��ZE�2���N���m���Rۺ��kdְ�2�R���l�U��jBz�)����`�`	 b��mmm ݵ�  9  �g�Tͽ���T�^Wl���+�6ٶ�  mJ ����@	t�b����-�p�3���@T̩� ���uPT�7J��T�
��col{j�P������2$7m�	�R�T��P Ә_m5K3�+mҭ]�*T��HJ���G[T��յؑ�[!A:�iM��ڕW��iV��6;gc��)2�v�#<l�t�k4p���s�;IZ0�K<�ۤ�]X����Xr��k�-*T����UV�4�� ���-��	UTl�8�F�Uy8��#(�ݕk�H�F��	��^ˀ��r]ӖKx �jF�[Bz���*8�h���m�� k� �#k�&�i�7i�	Ѡ��Ip6�ږ�$[B]�n�^�  ��#[��U�P�/�v��.��/MI��i:�M:���m[Vж��gnM��Fđ���SUJ�@��e�I�V��l��u��$�M� m��Ѻm�D�ɭ��8 L뮃�m��n��i(;9������4�Y��9%�mm�۶δ�պX�ɸ�H8sU�d�*�,J�*�{aj����Z��J�-B�u�A��*�C�����dmgM̀ m��w}��gC;m�sm�V� 'K�Il�[l��ҰH��V�J�X+�;&��%�n� �v���ۗ�=����ź��M�e��ր6��5��e��l���:r۷kF�@�aY,�u*�T I 6��'��M	$Y��T�\�M��J��.{LQs�l�UX²�̪SZ�MjJ� �+k���*��e�b*�j]cj�Ŵ�It̓e�v� m[� ���T�Y�` 	6ٶ�lk:uڪM�:�Ā�[-Mv���q+,��T	ɞv�SU�o7:6�Z  ����bG�Ջ�d��ܕ@P�l�Ҡ7��\m�����̘xZ����8*��/.w�`}m������z^�@ �hض����t�Rm֛��7@UU[6���Rj��]�b^*��	�M#��V�����#�͔@e�n��lۉ�}o��n���l�m�  ���cm'6���Z��.'m��U��8����m&���`-����j�e^�k��r�4�h���z��� 8I��U��,1o#AUl�̕��@C����M�h඀[��4�MVֵ�   �4!�\2g� ؕj�����I�rl��rI4*["㮫p�Y��!�Z;@5R���3sE+�4�u����8*��2�b&�U�V�
徾Ի}UQ)@A��w[z�y�4X`�k��mtӭ��������5�d��*�7j鳒���,5�y�#���F�����նk�j�������Jmm��  K�n��]�$���Ͷݫ\$pӧ@�hm�m[����Im� ��9� �j��&�I=@��s��m&���v&ն$lE�!mm�m� q�z���8���	e �F�se�o Hsm�8��mU� p8p$:^�#�@��    6ٶ�� �0 �����B@q 8m[
Ix�%� 7�a�ݱ��ۮyz�@ �i��9� �J���URv�t���j&3�t6JA!��WR���y��U���*s�h,��Cݻv$��l�*�R�h�I@���T���TYC�(���Ā��WR�5��UV����n�@ݡ�-J�0Eݷ0�m�gMj޺J��I˺V̀J�I)yj��ji���*Ut+��U[U��<��`�ۗ4��l��m��GinlUGd��UM�}����+�N��!�Yl�t�o`[%l m��fNm��޳$�uM{ �i]  �u�m�`����j�W(ܼ�λP
�J�ԫ��N� i��u[1�N�:D�-�H&�-��� ������ �mmmK:�ݶ�$�$���Uy�AH[*��jgIy�,�� ��{6#V0�Jg�Zl�=� [��mmӖ�-��N�I������vc�[A��
UR�6CK��8�$�)�X.���
�v�ض��
��F�����[%| j�ۀ�JE�� �s��;H< h�$7 mO,�ݞb9�%mp@T� z�I��Ȑm�����*�ڤ&���j�t����^�[�d�b�S�m��;C��0u�m�Ԍ6��[@��9�Ӛ�m-�4�徸@�U��6S���9r�T�U*ʽ:v��W�4%�m&97N�m� �aŮl �ɵm�i4�$���g�8�dt���t�  �g$����ں���<� �܁UP2�A��2�m�� m&p!m���G��6�� %P%Z���b� ګm�`�$N�m�6�Ӥ�6Zm%́�Z����]�r�C3�*�
����k�n��k@�������h[P�v�S!�V����]mJ��lhpK(H U.�G+eN "]���4P��݄:Ce�zֵ��l��n�9�d���J��}��u�~���8&P��֑��j�[��%�K�M�M�n�H[lk@�É���n�8 qx�    �I$��ͺMشS`r@۶�[�[��U��.^�޹/=	="҆vݛ%�J���ά��Fw�7_Rq<(D2hBs�g`n��OCٜm�IӣZ��� �*@)��>� ��4���l�L_M�<����|1q��#��!�q�������x.�(�#�A ��,����W�3瀧�" iqN"�a�P<PS�O�RU�
T�9��E�Q'UP�P�k��(����Mz
q�?pN{�*mW������Q@ү��'����<E⦼C�Qמ(U�	$4���z�� �=x(��:"�����x��<P��C����P�@t
ʇ�+�.� �H!�Qu�� s����iD8'��m^�@M�N����:uت�tM�/C�/>t���0C��==�Aₚ�O�A�O�T�X�(U�������tD�@�X�a�b��)�DN���4D@1
�,Bğz�����v�z���
{��up�d � >��*t����	LV���fb�NC�RXY�> ��gC�A6<	Z~}6����.�Q���D�!��ꦀ�ࢨ���&�$@� (� �����$ےI!l��)7.6�d֞�%'<<��Ξx9��=�z���.�6��HEB��q�M�KQ=�US�2Dɫ�S��Gw<�U�m�`��;n��;#�ae��2���k1�M7q6C���r���ۣs�&�7+�˥-h�l8ݚ���㮹�۔��q^/t�N��C<��uo4�֤q��kQ;ku��4�9����FL�%���:�&�/c��Yj1�Ct;>\��[t���\N6���r�\�6����Nqù�ҩ��]�']��@\1���$�	X�B�UmJ���0iۘ�\(��[dY�� �U#�S76��O;��B�'=�WA��Ni�CB�&��ڶ�^��s�M�Z��\��f��lr4�@�bq���i��6筑��'���(�\:�Ě�7J�ۤ5�[u�ZG�5݁0
�E\`i3�]n�C����g�5G1q�fLDq^�g��=��YI�����Y�R�K���������-�g���h%u�_/\bt�s�v9K�s#�=�@6z�S:u�\��V�-����7b�]T[����ۈ*��ݱr(a\/Ny7vh�r���qu�J2m�ݢ�g+h����l��'F$q�v����@��í�{p�ڤUi���CPZ�.� [D:�c>�m��b� P ��gxW�u����]� !�\1�Z����v�i3��gv��\��4��μ���tBm<�:��:�m�W(�zv�,g�{/��v[j�܋ѭ��;��%�)��R��2:�6�����8J�[�v�l^j�Ʀ�x�r� c˺�x"�ѡh
3��(b�g���N�m�N� ��t�Iz��I�����/(�A���r�p�g�[��K�X@�Q<c­�[qֱG��]hy8�I�m��W�=r�[�2�P\����nE���9H������<lt�E�Q�Csqa'���ܸ�'c]��s5������>;T�� AU�� x�����>�>TP�
����{{���~�ԭ ˱���ex�mB�Ӷ�ѐ��n�7[�
�1��T�<.��͸ʻoP��+.u�K�P�*�<r��u��l�(����P�nޫ�ȲoO=�.;m�M�v�g�0cl����-
��u��l�\����x�������3��شg��a�H܅qr�G9����Mu\���n!.�8u'np�Ƙѐ
qS�_C|�����ɕE&NG<�{n=�3�;����QWa1���!68�.eD�gt��T�v�W��
��O�n�$�Ku�D�#2���k�s[��U�y�ݶ`.��$��$PMI#�;׵`�� >� �mx�W/cM�I8�V׀|�k����nˋ ��cQ�["7D9#�Os���n�`��`�� ��p���Q���A2̜	)v�.�����6;c�@�D�h�Z�Y���e�vÒ6�M8�I;��K$��j�5[^�� ���i7"&���k{��W����=p0�<GH��" ֡�S  5w��B	�W�D�-�<�
�׀m�v��ț|RA)܋ �mx˶� �l�;׵`��[r$#������x���� H��z`��`k�`����p��|)�@b��@f=�@^��@Z��D� W|t-��%�!��I�j�s9܆^��mjQ��i�-����N͎X�<��A5$��7]��>�j�>]��[��qP��lrH�������:��xV�xz����662fe�̪�w:�:2=>ۃެ R�@s���}ט����,G�������r|�|���X��X�v��>��T�&�D�Fܑ��yP��P�t��y�Gl%����-W:;l-����2[	����+m]iu�RI9n�x�
���V׀vـj���{Vzͣ��#������O;�/ꠑŻ��7]��5[^z�k��9$$I0V׀uwk�5[^ }�f r�dI��H���G�uwk�5[^�{�����LA���jQ<T���m�E����u��=�_=m��#\�ǀ}�ՀZ��@b��@b��@Z�@ rLNZ�v.ܳ9��l�n�����Y��� �g�]����I#�bG.uS�٣����~4-�t,�t��T�����M�I|M8�U�xWv��v���^.$}����Q)��#�;׵`k�`.������n�12�1Ir+'�T�M�d��n�$�n׀w�j�/y��K��NAIk;��DF����@Z��@{��� �8t�v��F�ֶh�އ�]�[��NBI�G+sJ�-��q���K�#��"6�TK&�8=v�n�*x�s��;�P����.�ɪ [��&�v�ɒ��c�y�z�y���<��뫋g�<��ۍڙcE�ۋ��{��Z�ݵYV��<%�v��Ž�dϫF\�v�k�v�n��Ɯ2N�r랊ܰdm��΅�$�vp��@�,�P�D�o�mD�ƫh
� ��{���z�}$�;���j8���p](�L�qx��iu�6�DstV��\���H�$�<��<�{V��^ }�f nԫ"S��E�$� �=�_�	�� f����yդsb�P�J4䑠#� �m� >� �ݯ �^Հ[��H�k�H��� ^wM�w����k{�y�W���j)$O��'�j�� �^Հx���y��d��!��聓#n�fĎ]ո!�:�1�,��ޫץ��0�ݜ���H����"Q�$����^ }�g��V��_�߈��$�)%���ʼϻ�s� �\�P=:�� <D4�����o�{���r���X�6�Jq�����ݶh[��Ǽ�[��ƹt8jT�H�$���s�]�x�X�mx�m��ڋ��$�	�$xc�T����|�Y�}6����<����k�!ӓ]�]�;@��Lii*M�\㧄���q��k�+T�i�k{� ^wM�w�����C�e���0�R;$�w2^С@$|���7]��>[k�>�Y�>���re8M9v������0�0#� ����	��s~k�{����^}j��bc�$��� �^Հ|�׀|�k�:�k�;��F��$�) ܕ@Z��@��@b��@f=�@���օ6�v�V�l�̧�x��cpX���V
.[)�&+k�bErQ��^wM�w����k{��t!0�$�BJ�Y'���P�T>��XU�� }�f{��m�{�7 IRH��|��ڰ��0���e�,	Fܒ4I�+'@�콼�W�~��U�}�u��t�o�~Ec�@�T%��+$�c2$�M�$�.E�vـ{�9�v���x�>�i���������8%([0��K�?������ّѫ&�h�b��ԝ\���J����rt
���n���V }m��2�F.6�#M�$x��g���$g?�T�}���y����}�#�I��>�j��� �ݯ ��L�=�M��E9�X��`[���)�}�Հj������$$I0���~��[s��v�~�Uy��|�������5�������؇Oi�MNŷp��s���t0��5�l�\qt�#���m�8�[�s��۱�.�*�%;$�(Sg�碵%ۄ��&�����+u�s�.-�u�4�[n4nׯ\s����p��srm>_
��=�-C��mpD	���U���S��dAzo:+��^���[��y{-�:�4�A�ӴݝaÌ<R;N��R�S��:z*7�WB����[�fY�vh�� ۠,I�Cck�<��2v�,gITν�)��;���Zڢ�U?�o�����V }m�V�x�5;�8ےF�����V }m�V�x�ڰ�-�4�L�G��Ȱ�l�:�k�7vS �]� ��M??�x���r|�|�ݔ�>�j���Vـ}�-ci��D�rG�n�������/�;�z`[��ծq��l�>���ۧ�َ[���Xp�E�í!Wl�-��[]&z�2����P�t��y��Z5��\h��&(!�Ed�]��`b��� P�)�쓙�Y'�y��<�KJ
%�HI�I0���݊��v� ����Ӝ$�	�$x��V��V }v��v���H��mF��5�)��V�^��d��{�{ֳ�tPѓF�l��n�3�&b3�m��,�j�k�7l�F���X�n7�DuS�f���?����y��w:��*3��.���g����V���7Z����U�����/���sC��X1țnM�}����r�>�{��4�D�̈���@�f�D�F�Y$���0֩B4�	�m�e���D�m���(S��،a�#4Y�3Y�m4G�(a�4k�*�A�d�Ŗx�,*fc�Ha%��F/�i-0� ����f�ֱњ5���Y��kLf�46�����05���y��I����Xa��a.��V�Zӆ`9�h��bH�f��و��h���xq���|[�����͑�oq�:0Č[#�17x�d�Ϫ���)�٢O3)?a���!�p9�z��
�~=� P�G�� ��~� Gb�� ��D�w���*���OٓQi�����$-�	���^����'�͖I����?| �Z��d�|��c�d�1Ȭ�{�d�N�C���v�_|��ܨ���>N�zdb��� �H����j�Q���^d��[�5g���$%|*�V�6J�0X�RN�q}��@f5���ܾ���7{����p�5$��=�Y���G��U�O��,�{�d�� ����|��ܑ��)��� ;ݳ~H�}0ֽ�o�ͥ��lD�>((���n�U��w|��u��Xh��&Ab(
�P�TU����|���σ_���فM���m��7������� ^k�7��nd������pu^3~_>ﵚ�=N���e��7���A�w:�6���M�$���x��X��V�x�i��P��$N<�v� �v��v��j׀^��qĉ$"��r,���v�|�|���^��V�iR��p\�pRL�:1��@^��@b��@��d\�q15$� �Z������f�$�{����P �w�HBlJM=�{9�5nx��`��W�F^k��3�v��;sk�8�MŴ�+6�>&�8k��Z�gP�ڇU��S4m��k����oB���� �]B�mz����-�t8�I58�5��R-v�{r��ڜ���^���ut�<��︱�nܚ��cVjȉΤ.�p�%U���c�z٥�Y���	���v�mD�hP@��\-		q �Enƀ�)ڗ�ڷJ��9����Q%G��nՓnMq)r����H�׾X��V�xzկ �˛R�M��$|PQŀ�ـun׀w�Z��ڰ����.M�b8�mI8I���${�{� �~���ـ}��\PM��D�rG�}֭x{�]��X��L�v�z�j�J)RA���>�j�>��n�����t�]΀��
��ta䛷57L#u8�3�9���z�UuN�
YKnU�vj�K��W#�!��4-�t�]������|�Y�J�0X�	)�d��{����կ �]� ;�fu����9LQǀ}֭x��Xy��f�0W|�ָ��9�RF��x��� fwM�w�x�s�7�c��iH��, �m�V�x�jׄ�y�+$�P {!(-�I��#	�dS1�k��X&Ĺ:���v�<����%qKf���;�"B�a�$�'���<�Y���]� ;�f���9�J��M"9m��wZ����V w���v�z�j�J)RA���>�j��2Y�P��PU(
������'�k���YyI�!9�7 w���v��k�>[k�5m|�L��䐐��:�k�=����{��:���	�s%�v��� ��k<�%�Q �V��k��-���z.-�+X]�.�M�w73���`s8HEË�D���k�x�mx��0���ъ�$R&5#mp�G�|�׀� �ݯ ��Z��7��?4�I#DQ����`[��u�^��^{y����3�7	�fl]�:��@Z��@dG����&���ԉ(���� ��t��t��4��t��BϺ1�����!��
�H�3Ū�HNw]&.;/Z��H+G:"S��ND��5�g�:��< �m�����կ ����!9�' w��V�x˪ـ|��>��V��"�A9#$90[��.�fK�����z`�lK���D��x˪ـ|�� ;�f�s��v���o�I$cR6�"RL�mx��0[��/s��*�	�D� i �)ZT�BC$f&H ��l�~�6���9�1Ʈ��q�R�m]�Yj38��E���)O+�1f{*`�sM����m�1�.�w@�mRmȐ����1�g��;������4fƬ]zvCf�/^�Roh�iӷ��"[�D
�+�(���;lM4�Vyҍkn��n�K=�X�w%��Zi �f�pL �[f+O7u�N�������^��N��`��%I�Lv��T�ƸE�[knge0ȧG��K!��Z[��q]b�f�]]aΪM����?7� ջ^��`+k�/oy�q�8���*�� ��Z����{l��F�,�ԈPDr&ے<�׼����{l�5n׀}��N�q��m8����{l�5{��]�[��>[���pA��t��4��t�]΀��΀Ղ?��"�1#���%1e���ˮ˨r�u������_����G%�>U�x�j׀}������=�i�QA	"eD[��<�Y��PBu�)�(; ٰ7m@# qة�C�p=<�<ם�U{���*�>���G�9��)�jF��� �~���ه���[�wZ��o,/��D�$h��%��LU�x�j�-os�;:g��s�R)n�����>�V�嶼 �m����h������p��\n�����κ��.:N�5v[t�/�bm��9�ݩ֦�]���ҿ~v.��@��@b��@^����$�' �q�k�g�s�m��0W|��կ?�5z�A�"9�"�ӊ�'�ݖI����B��]U�\�*��]�s�ڬ�Չf"�$�H'$�:�k�>�V��v� �m�洊���$M(ǀ}֭x�l������:�k�>���P�Q�OV|����upn{HY�V�Ol�-\㧱k�6ȳ!emG��R8�jF�)	=Ǻ���`]����^��7ǽ�R8�L�F�r, �m��[|��^��O:��G}���fJ���ʒp��7�d�u��g��7�|��s>�Y'����I1țm�읡K��u�'�{�9U���gUG��_ 0�?���~���;��
�����vI�^b�O�_
3�I8�~vI�Z�vI#�̉���-������n�#nI����T��Ct0b������9���]���ln����y��w?�=h1}�:W�n�b�$�HS�Y'˾�zRG�ku�'�s]�O{�/@��ѭ#�B)$M(Jq�'�۩��%չ���@���L�|�
�����'���E"x�����|�w~�Y'���d�_P�L��쓿���F�rH�.8�}��@}�DDs����-ws�o�. ��d���`b׆����hR��B�T�%�(bK�����ll̰��1����1�#1��1���,����1�&,' ���q0"��,��,�JA �����K$2�,L�XK ��8��А�.�eІ
Y��"f!�'^l��Y1xM>$��Zf�-!�Jv0�����!���[&��6����J'���f(l%4K����c1��	���'1D�|}���	�B`��I�4�nI$�G-�yn�w\�öooBu��ݧ���y4�5d�8»����\;۱�/��[��i��.;f�v(����tm�[�:���v�'����m�����q�ptT������O/���[y][v8ˊ���6�볞�vo[�q��]�g7�W�m���u���&�v:�ɱ��$�{1E�@��н h�	=mq�`�5 !�Z�HL4V���dku���}�����ˣt��̆(W:�t���x��;<F���n
�WP�	��<���m���h܁�@�m�^�����c��Z^UZ���t�eW}Ol�%�)i
�MZ��J��sͮ�㓔7��x�8ڴ�"A�75��j�p���m�[V�&��ιnmb�l��m������Zn9�zl�)6�#h�MRf�L�N�q)�ܜ�j_`��a��k����
�{�б��q�Y�T�Z����h�&�M�=���y�XZ�.�=ΗF㫥[k����A� �Mz��f۴�ΏF��P/a�.�=<^��;÷����e�\5��r%Y��q� N{c�b:���x疄{l�x��v���e;%��y��Q��gY�-��/�/`�(�nS�@%��}-�m�@�����i737�.�nrlQ;v��tƦ]�S����m��6�qL��[l�5���v��F瞷[N���e;-�����?css�g�;,���g���$�X%mrt�q�v9r��v��A���՞��	��7<s���sx
V6��ɫc%���ݣd�uu՗��i���`�:��@B�-Çk�#�!s��<���\ƻ7�wJ4��p;\�n��t]u�D�Ĝ㤋�v�<���ۖ6�	6�/<vjDvK�+�f��<��e�WIy۝b���6WyAn��h�C%Cc�W3ٜU�C�{kn�=���n�`�L-3#�p�v��]������T��\���.֒t�:[R�g74��	�͹gNil7F5o]z^������"�}~W�<D؞ 	�G p��t*?�ΞjՆ2s�S��Q��G Qm�[�񟟭�,�Y#�3m�wGh���t���s9�i�X��0���a4hr��X�q��KҚ�z�=�kS��⌖d��I��N�s�������wXyճ�4U��w�ַ�kȵ��z7e�uv�trD�/m�lmZ��c���e^���6m��k�1	��tg����횜����<��� �����;��st]����JjƧ[]9�����y>���S��֐��(�o\Z�XC^�w{���}�,Cn%	�$�I��~������ř��UU�I�ݖI�#FB�4ێ;$�w1;�� ����'3vY'���z �=͌� ܎(����:��< ݶa�����Uo��۩�'���H�J)�d�V�� ��<��l���s�����^K���9$$�rLV�x�s���{��:�����`m�(N&�|r(R-��h�m�rD�&�<�:9�Wܽx�n9��+p����ŐbA$M.F���^��>[k�������|�+�6䐐RF�1)%�x���U "�Pb�����o۲�=Y���ՙ/��|?|>�rG�F�q�d�Y���>^�;:��ݖI���d������.n%-�]�˻�@Z��4��t�x~y3}����ي2����Y'��ـ|�׀� 7�f ��g��������݃����ǭ1�+]6�]B��x�{����������~�ߵ���'�̖I>�}B� q��,��ʿ)����S�x��3� ��Y'��vY'�َ��*�����_|bEB`�!NId���K$�ufK>
�{�����< ��0
�IU`��!�ܖO�B�R��ݖI���d���K'�/{ �5P���
H�iD���u@�٠��-bޚ㙱�R���Q�Y3֣n:z�!��{bz��mCK՚��ۍ�t婖�6J~�o����h7zhX�����΀펎����Y�b�|��`.�� �n׀vـwlu�F�rF�qɀ|����^ }�f�ݯ �ظ:nGNA5$�>[��ݶ`۶r��A�"� ,�����?<Q�k�nrr)�r< ��(�w���|�t��tgG(qP��[$u�u�l�*H!��9,<�Đ͊�5Ӷ��s�����q�h�I?�ݯ �v:����������e"d1�#q�'��x�@� $z�u�^��ջ^�sU�y$$���� �m� �[^.����c� ��9 �F�$�q���v�����>V׀m��g�А��(�A�	8�5�'�*�{-j�'�w]k���4\҉���10LpCwf��b�w�[�kdt��ݰ\�����jܸ	��j�� �I���#7$���X,Kv�mPc, i���a*��-q�kV������t��<�s�ݸNy��T�{��8��r�6��A����ˮ�Rݞn��un�a�w5�M�<�:ۮ�n.����גνvY7c�:tk=��@U�f�Jv9�����g]���3��^�}����}}��t_S�es]�u��GC��,BuFoI:�V/5"�?�o����|�� �[_���s�*�� ���S�E�)VI���{A#վ��*�� ��U`+�������I������k�>ݎ��mx�R�D�''$�%x�����V��v���[Vh��\�ǀwv:����+����ߟ���\����:-�x�Enı�î���6�ķ$���i��F��H�cqŀ|�� �]� ջ^����-���"��I�<�v���*�������'ّ�Of;��#�7K_rb��q�w�wv:����+�����pn)�I������ �����`{��v���.� ��F�d�ŀ|�� >�f�v���Հ^u�ò"�.������̭{|ryY��/�5����� �5:�5�U�:��n7�]� ջ^����>V׀}�mm"rrNG"Qɀjݯ ��u`+k��ـ^V���iD7���P���^�����;�hWk�>G6���AN)#i�� �[^ }v�V�x��~V�^X���$�i�9$k�8��l�5n׀ovW*�w:�b�c����LH�Cu�%#�¸�v3�Ѯ6t�S��"m4�5����H���*�� �ت�>V׀]� �o.�m�$�F�@n�\�]���zh[���z"-�\=8A9�8�qG�u{�x��x�����^����9#�|�Ĝ� >�f�v���ׁ����C�� ��c�O��aq��H#�(��5n׀w^������l�N�Y�ָ̑��D��
��Ӷ��zx{(�ل�<ͣ�r]1��ݮ�ɀ�.�x�#J!��k�� �[^ }v�V�x����y ���&9x˻� _oM�w��������~>�$P4�pI8�}��,���c��{=vI���d�`��pC7�����?�������<�mx��0�ʒ�����(�q��Ux�W^�Ow6Y'���d��B������I��w:�b��[�Bn�-:�bU��[����V�O$�ü3��2m�ʺ-���ӣ�[�a%)��:E�gL.��6�qj�ɚ�U�b4<���4�V�S��b�O��&�e�qg��{4�v!����֣nL��&f�F�.�=]\��^x�;�W���!�^yvغ���uF�u�C��V��K3�]pɳ���R�g�uNG�߷�\g����x	�b���6�z千�V�TpKpU�b��&S�����;}r.'"��N(������l�5o��>Ǐ]�z��hn($p1#�9�O3�/E$qfk�T;�W��=[�����7�����G&�v�������	un�I���$��H�$$H�ǁ�s��W�u{�x��Y?UP�_
 Sٻ�N#���fB�RF�e��Of;$� (�ݜ$���d�y��O�����!�nB�o��sN%�����;0!"S]�ӷLu��LF�\�I#li6�$�q��u{�x����?<P��8����d�њ?G��26jG�N,�w��!@U*-h��PΈ*�����5�W����$�fc��*�#�=a����8�n8쓋3K�Of;?����U
o�|�/{���X$�q8ӎ9 �]��]��[��>��G�>�@b��HP�BĎ$�vI���d��UU]�U�����q��ċ.�A�kKBt)s��]�Ye��9:�tstV�d����{��}>F�G71:������d�/{�O{¨��
��q}�����bܑ4HH�� ջG�Z��@b��@j��_z=�z! �K�������i� ��_<���||O� �U�%C�! �1�B��D��p�/��A�%1���a�ADELL2I%1EAQ0�0L�+e��$�wJ�D���	$��Y�XChL�(�pTغB7�6$���F @蘂�Bj!�]p�B�9�P�6�$Q-(��!��*�6�:���"p�c�DIQ��4Z��b"a�)(�	ih(X�I v�j�5��3���rimk4樾OQ<WҠ�s����|��@�E�EO� �Dت�|O�T: ����*���-�]�|��]�s�"Q��rH�rGd�
�w]�q{5�'��x��Ş�$sFh�,;QH�A�	:�~vI�U@P w2ޮz�5��=��d��n�����AIE(		�vɔ�q�d�e,��4���M��0���v������{��O�
)'#�F��?����|W�� v�M��*�Pd����'p}
O�IN&�rI$�^ v�0]����*��P�H��-��B�0H�R;$�n�O�}���P�T)�׿d�/��d�.��1�!���$�tAc��v��������0
����4HH�� �v:�~�ο_?�OwvY'˾�d��v�m�D��@ƤO;CvV�pV��Zūh�q��X�똖�em�m�| j�L�#a��.�|�ߝ�[f��_�A�c��=�x��Qm�#\rG�|�� ջ^��u`/f;Ԏh���DŖ�l ԏ��[�<������u_y�}�L�t���j%R;'�
?n�����|�}m�V�x�X�q5��8������{��5m��7^�`����@�g�8���Y�	ڿM�O��@;tU�8Ms�Y�g�<�9�IZ t���ә���r��p�Z�F\Uk��`X����X��)�=u��{9� �:͵pO;mƈm���<;�k��u8y��v�����Ȟ6�2&Ҙ�{�`m{p�l=1h�ݺ�B�y�����Y6�l�Lfn��0U�dm��M6&���<9��l��`��%�6�����ww��C��T�s��Hx���������3���
4����Yrt�������k���F�����ݯ �{E�|�׀ov*�k��4E �$�5wk�~H�� �����f{�G�z��8�$$H�ǀv�������?$w���*���V��i�$��i���>V׀[f�v�s������'�H�nI�< ��0s�+���3Z�k��x69���	���m���`�}�|o�3e�4&.��ޢQU;�tFA�;���ԍ�ʒt��w�d�u�c�>V����s�wޘ������7��kz޹W����s��� �0�5F�� U@���o�;$�}�K$�{����������>[k�����Z��t�3k|�p�r$d���j��넟,�vI<�@.?f;$�-Q4#20���I0����ڦ��^ wm�������le�HT�����Iֶ��=����l;��
���Zcj�[��;��t�}��ʚ$$H���}����^ wm�� �D�fk�I�X5
mI#��4��ty�4-�t�[�_{ޏ
H�"i�Ɠi�#A��O}�,������@2��&`iQN�
(��bv!�~ �AO(�e�|�5�'�}�\�&,�%�LS3`j����oMk{��z"�%�n�$瞵��r0�J7vI9��h��z1��; ���1n�*U$�ņP�
iHS1cq����N��Z�{N<6�v�:�:-t�k��X���ț�O��^ wm�V��� ��I�ߔ�Nc}"-���##%��{��z �)#噮�'��S�\A�}�{lG����$�V�;$��T��������O�f�$�'�Z����d���vN�%�f�d�s��k�{�}�r�R����=���z��d��RH���L�mxވ�{���v.�����GT�Ѷ���F�md���@f]	�t��8'�j����V�μ����{���n��U�Hje���t-�t,[��=�}�O���_�K!�4��'�3]��($|��e�z�u�'�����*�6w�&��6�D�q�d�X��d�/f<�ݯ �ݯ ������B��Y;B� ��u�'�ٮ�=^�;'着�Sɋ~�I�`��Q��rDdd�k7��#��k���o|����Ί�� �*N�ؠay����lX�[J�sXL��T;3��`ۀ:��I���iñ�g�V�G%�k!��+mtc%,�2t�%mU�N��B�4tЫv;�Vd����g�[5��GmG.��YS�qy�����.퇶�kO����]���������x8��ܣs��6�>:��S�N֎ݥ�2n^0����4��kQ�=� ����m�����4��q�{��u9�z��7�gn�ˢ�;'"�g����;J�4Rr�T�l4�λ��p 	�j#
R0���xI�g�;$�wj��mxV�xA��x�C$m&�OWW�_ꪯ�P��/���'�>��$���z*��"skI��jIM(�� �����v� ��0����>�(qD�M�#h8�t
�_�]�Nfl�OW�Y?P���
�>��d����~�n�jF�H�I9���<][f�^�� ��U�Q�s�q��YO4כ�}����C���ݺ�ӯ:7��$)ar[���U)fݣ"�
q(�rt��~�I��΀����{�h��h��A�JCfC����I��c� \��PT(Gz"=���@��@^5���H�|9��0R< ��� 7�f�Z��������%#ℂ$�߹Į�L����>Wk��?q.�0 �b��HII�0��׀Z��@��@��@o��=0����s�-�!.7=�n�%��'�F��꙳/����ձ���|·iJ��O�W�� }�f ov��Jqq\1����9#��l�~��]���5��Ş�{A#�/4}nݦT���7��U����ʽ�~�b��%(J¤B�������7�k���'�ݖI�Fa�bA"N%�K'�/=�xW�� }�f�?%v�`y��Hl��q��x��x��.�>��xWv����$�jF7���h��X��<�8��k�4Ik��W��qK�ܜ�O��"F��wޘWv���^�� ��¤��|P�)$�1f��m���t���@��@r�^&�	#bn<��^�^�6}�},��7�d��%���ҒFQ�읥׹��'�ݖI���0U)jP4J��z����fo��w�Ae�m�#h9#�I�s%�~�T ��7��N,ߝ�x�1�'�{+�N��q�W\�\qmX;7Y�F�n8��L�A�(�K�A߯�����J?O��߷΀ś΀����{ր���3O�Ȩ�I)ģq�d���� )#ջ��'�ݖI����ꪤ�xl'`��nGd���vI<�d��,Y�����d������PrDdd��� ���d�Y����c�~��^�$�Nâ��''�
I0[��]�����U���W��D�"�-QD12A�0A%0D,���1C0��	10D�R�L012�LK�UQ�10LQQP��Ħ)`�`��h�`	d�H���! RRXYd �$!����`�$�jT����&A~�8�!��}��e�9'li�Y�D��,<vxS��3!2DCE1��@�P�1S0L�H�$�HB�� JȔ���(Q)I!J�,�C(D�S3Q$Q4S17(���0�9�n�m��-��̲2ö���Z���Ƕ���o��U��/R�خy��7K��0\�b�+�ng9�wn��
Vݛ��k��"�Bc��7(�]\����8�Ar��^v�ht�a/q秷8����z���˶=�;�D��9/nM���c�(6ts�<ݶA��g0m��l��p��������m�q�ۇ5�m��q�os�붇��U�6����;&58����oR��K<���nw��CɌ�4�Nր�l@e|�X2�څ�օ^z87:�.If�Rݩ��r�c t�&��lU�݀5�8n�T<;�y9��ma�0s3i�r���ͥy�vU�UQ��@p�v�k_5�u�s:��l
� �n��s��v�sm��Xp.��O[,FH0���mp:E��۶�w��VԻk��� �K�mk��f�n�����nU֭�$	�ŷ�rO+w.�̠bz�O-����٘N
���p�i�H�xv筜�[�kmVE�k��7���I�ۭ�¹B�dԔphݎYy]�u ��*:6�;g�8v$b�[b��^)B��xN��۷K�e�m�^�s��ovA�L�����KL�P��qc����`v����Υ��a��*�%Yp�[�F�M�Q�۴��K3��-���m�����{��Vp�MY˄�,4Uס�t�kۄ�:ت�����s;C���E	���H�����bvͷ=7��[oN�� �;�X�\�&�(]s&畣.�ku��i�g�`���&0�z��u�i���5F:��koT��{s�m�k��]qڧ@�d�j��f�],�e�u�c�<A�#m�O��kӲ�sѰ�:�S�����i���]�ӻk�����n�Ӭg7Lb�b㱌ܫp�.f�KFu�qɸk%/.��	�S�N6�5�dn�9�{���2.%��=(d�&��8�vIm�n���&v��s�����(�Շ�[2���:��D<��˼�;���:�ٹ�۞��ٮP�P(Tq�0�d�A
@��:C�"}� ��UV<@<L��:'����k��_~��u�s��!}��Z�F9���`�|Zu�u���3C�0v�z���ئ�[e�m��'��Z�±��:��7m� મ!�@�kw��^�]t�����3�v����P�;E�v��qGg��s���m��|`�;��)�m֋.b��Sd�5J q���m94Ҙ�������[N�pVz8͖Xh��]$����[�W����뻽����Yi�Ւ{E�nn����K��i<��*����:ɱ���{�G��!�mR�g����n�$�g��$��C��Y�;$�>_��q�RH���G�|�׀vل�.��O{��
�����Hρ��$��8����� ջ^ w�f���d���s��v�QH�	�$�?T Z�~vI>�l�Of;'@ PK�ݖI��/39$�	ģqǀ�ـ|�� >� ջ^ oo*9 �NGv,�S	�p5z�7f�����DlCGi��tD�i���M�aM�4ܓ����v}�4��t��4���>9ݳ{�f��Uy߻�z!�!������*�����m�ܮ�N@�P�$�N,�vI=�Y�;�� ;���>EU�(�	#bn< �v� �ـvف�s�����5x�q�8�q�%�Nfd�N�]���^�� w�f����i��G��-c,��Bۍx�h���,+7nvk�lWM"�'�&�#k�8���0[��I�}���'��vIϏ��o�U�a2��$���������e�z�u�$����ԫ�E��q(�q�{�|�ϵ��,6��`b��W�����V�<�=Ћ���8�MI0>�5g����L�v� �v�����
�12Ɯ� ���x����X��#cq�P��շ*��A�X9��Q�]Ȇ�4�)L�vL�%��"q��H�I98�PRI�un׀�ـ}�ՀvـTj��D�8Iq�{�g�;_����L�v����՚���l($q�aNK$�f�C��0�9�6_{�`���ҐM�HMF���ݶ`wl��l���)�����IL�@��4�a8`>��ں1H�d�D�D*wת
i��?�����?�a1%�G���� 37����΀/;���z}�ɡLJPZ�bV{i0n��q�u����J�����5{-�h��Փ��u�k��!��m���������^ }�f wv�{�
���������Y'�َ��W�ϖ}�ڪ	����o�޾/'�q�NHƜX��t��4,�t��T��p�Q���AI& wv���^��V�^�� �+��N�����1f�?gO�+ ���1n�+��@��#�^;���Y���wn�Y���t�mu�ي��-�KJ��g6ډq��p���1��l9ۚN���H�*��c[K�R��l�= t.x�d����j�<g#nr����HY;�r2\8^;h9�B�NݜV5� �`Ԛ����8�x�r��<u�Z�ӭ]�U9-#�M�go-����h�I*:6��/b=1��km�k#n��X-���.�sm�:v��r;b�z����e�/��N܋��Q�0����GC*�H��D��׵`ݶ`[��]���
�ĒO�F���ݹ/h��f�$�{5�'�َ�UP���9��/��Y���#�&T���_}��'���G{�b�Ry�4椥��������X�y��� ^wM�w�����F@�mH��<�d��Aw}�����:���6�yI�8�B�8����P�v���zs�F{q�i����\�K�����>9	�Ӌ >� �ݮ�=]�?�@u��|���7�j(�rBr�S34-�u���\y���ts�+$�w2^�GQůB��L�H�� շ� �]� >� ;�fW����0I#��vN�UK�7]�uo����`]���,J���F�jGd�.�;?%�P ,��p��7�@Z��@^@��0�0���s0�H���I"��}�d�v�ƫ�4i���[����h�,���	��G�Ƥ} ����:���-��
\D�{u�'�����-#q��s4,�u�=�H��|�[�΀Żζ�U� 6}��O�B�)q�#�������^g��u@?�Za%@B H!IBI@S� �;��u�-�xz�P^N�"F4��� %�n�$�fk�OW}���R�M�d��zޖ��� N [��=^�;$�({���v���P�t��5�L!̐�3д�Ȼ9�$����o<�׷gJiQ���!v:ۮ�YBڵi����~���؜��VI<�d� P�'Vf�$��L�q��H�"'�s�1_�V�l�d�d�Y����c���@Ώ��/���$mB8�o���*ݯ ��׀^��d���f�,��#8��?P�|�~vI9��d���VM
��{���%/ i��� ov����P����t����쓋��d��2�,�d
��9��ϭjwFG6l���N�N�7f��m=�r�U�����~o�-v�9n��=�@v��@n��"`s�D�p�>Wk�*ݯ 7�f�ra�� W�B�g���\j"��8�8���< ����>Wk�6��x�P$$#��=�߹�+�� ��O{��off�$��V��F	$aS��<^�vI�B�� ��~׵w?~��*����@+��N ��۽����A���8+�r�ljm�r���+;����d����>-�F�l^Ly�ʚ��9�0E��kgT��ŭƘ㠕ySj�m��sa�[�P�-��;.����;m����k=��&����vba2Nݹ��/��-�s	�c��k�uN�b^z��o[��-������7;&�-���LZ�i�8ι���%��d��@�I¢!����W�U�q�dD�pM����&�aN�U˱Z.�ۍ�Ni��f����Ą$>I\jG�uv���{�O��
���=�d�i�c��Y�7rFq��O�f��(
���f�$��O{�  =�G��P��� ]����X��xV�x���qq����ԓ �]� �_c�OW����Y��d�y��Q�����iŀ|�׀un׀ݳ �]� ��r�8�H�98�("≡V���)��]��x�*]Rr��8��M�ן�w����o��Q	�����V���l�>�j��ـ^-�� HHFq��������!�?�M�w���9D�ٲ�=^�;�>���44��ٽ�7e�5��%)O{�߳�R��]��H ���g{�\R������Vj�5C�F,n�$X�6�r+��I��{��)�}�u�)J}��JP�ȸ�~���qJR����Z�����0�R1\5@��噮�4��0}�l|��=�~�)JRx{��Y�� P�F�#jD�0��m���w��ڢ�2OF�&��z1>��V�Q�`[�������	M�biFԏ��F�+�JR���߳�R��^��O�y4	�^�wT	����Dq2�I���Y��y)Jy���������~���)�}�����w�ǒ�T3�D�ԀȋN+��Es�ݏ%)Osﻮ)H)���!$��S,�C���З�X�E4\ �<(����XJ�Hy	�k��l����"Ya�&��i�b!d���!�Z�#�Og#�;y�X"$�c�Y��VfN�PZ7�옍�a�dc��ff�3���	�%Jd� %	�"E�b�`�TM��� I��@:(h�G�E8����/z���S�֐<����JR�wY��5@��ǐ8܍) N"܂��_� ?���~���({���JR�}��8�)I��ǒ��L���Z�ٽ�ݽU�o\R������y)@ �&?~���qJR���ly)J:��wT	��Ã�D���3n�������V��M��:�.e�s�d���]��J#�B���*�P&�s�1]P2��{��y)J{�}�p?$�)I��kf�T7kV��H�$m�WTR��{��yĆJ}���qJR������R���w��?��R���{QrH�8*�P&�yfk��MP%=���JR�}��8�)I��ǒ�j�=��BTj�Q�㺠MV�Q������R�����8�)I��ǒ� �K�~A[{��⑪����8�r$�n6�b��j�>�{�R�����c�JS����S@�=�1Vj�5C� ��4��M�.N�qv�^[��&`��Q=�M�k��W��A| �m�R"-8�T	��w��c�JS����R�����*�MP�b��MP&�<��8�jH�Z��<��=Ͼ���JO���C�JS����┥'���JR��x��Hd1�[��5@�=�0�R���w��)���{���JF�yfk��MP&�ymq(�H�;�oC�J�PO{�߳�R�����ǒ�������?��O���C�J�����$X�6�r+��hs��JR���w\R������y)Jy���┥'� �?��B�;ߏ�e>�r�$��3f8v�w:�۷V��#�񵃃k\u��v���3�+.���Ǒx��,G�'��)��R;��">��➉N��J��4�>�gc��i�����u͂ݍv�pc�=t͒-fR�F�e�]�ثq����:�;z|�g�v�Mۑ7:B'IR	)$��Wn����/n���j��e�Sۇ���{��a��k���Ѻc�	�,Z�>K������Q��)r�b�����`���m�#ச�MPŻ󺢔�����y)Jy����	.JF�}�Y��樞�m8biF�┥'��wC�JSϵ���)<����R��>��⟅�ZR��?3�j4\�����5@���|�������c�J_���w���)J����*�P&�w��G��r"-8��/�I�߿ly)J}���qJR��߻��)���s�R��}��d���R@�E�Y���{�j�?�?�{w����JS�����)JC�̂��j�{�M�I�EĺݝԵO1u��:ь�dn�uE�1��Ѯ�l�P��C!���wT	���ﱊ�JSϵ���)<��� ��JT<�5�P&�Cqm��H·�އ����k���-�#�TT�v?�$�)I�}���)�w���)JOo~��{Xf8!"đ��]P&�C�̂�R��>����  2O���C�H���WT	���`��B�rH�z��R��>��┥'��wC�JSϵ���?Y'���c�JS������m7M(�q�P&�CǾ�*�Q@ ��w��qJR������)�}�u�)J{�܍�-�3U�6oq�4�r�i^|uF8���jDؖ���N�a8�R6�j&����j�<��j�'���JR���w\�B\���ٰU��MP��6
bI��WT)JO=�v<��=Ͼ)C�wc�JSϵ������'������5��̐'nAVj�5C�3]�j�"��wc���0ԧ��{�R����Y���x��Hd1�[��+�X2���%)O{���)JRy�{���(K���┥'���Mh�"đB�nH*�P&�s�خ���}��폒�������(���Y���쀣�6c0�&�к��u�b�Rz�Ve����J�[�����p��rF�(�$m�\��hw۰U�)O3ﻮ)JP�����R���}ܺ�MP&�{&�%�F1�Vj�)�}�u�?$��w�ǒ����g�)<����O�V��[�~5m��iF��5@�^�lf�Ty���qJ���=���%)Os���Uj�49�md�4ԍ��� �5B���(O�s����(J��J��(L���(J!(J��30J��(O~����(J��0J��(H��(J���(J��"�r��(N����y��%	BP�	BP�%	��P�%	BD%	BP"z�pI���#��<C҄�0J��(K_����(J��0J��(J��(J3�(J��(J�(nB0}	�1$�H�N.pP$P$%	BP�%	BP��%	BP�%	BP�%	��P�%	B{�����%	BP�f	BP�%	BP�%	Bf`�%	BP�% P�%	������(J��(J��(L���(J��(J���(J��/����J��(O3�(J��(J��30J��(J��(J������(J��(J��(L���(J��(J���(J��?�_~?�����uwm��͖4e�8�Λ�v}�j��ں(�]�B��MWe��%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	�~���<��(J��(J���(J��(J��(L���(J�����(J��0J��(J��(J3�(J��(J��=��~�<��(� w����(J��`�%	BP�%	BP�&f	BP�%	����(J��<���(J��(J���(J��(J���l_�4Dd���D�(J��(J���(J��(J��(L���(J�����(J��0J��(J��(J3�(J��(J��=���<�J��(J��(J3�(J��(J��30J��(O~�����(J��(J��(J��(L���(J��(J��]��y��%	BP�%	BP�"J�4 �tj�KE��M&�*�]ǚ�44 ��{��~��30J��(J��(J�w���P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B_}����%	BP�f	BP�%	BP�%	Bf`�%	BP�%$P$P$Pݭ��(�)�$m�\�J��(J��(J3�(J��(J��30J��(O~�����(J��(J��(J��(L���(J��(J��]��y��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP��w��%	BP�'��P�%	BP�%	BP��%	BP	BP�%	B{���y��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BDP��)�l£RH�9b�"�"�"P�f	BP�%	BP�%	Bf`�%	BP�%	BP�&{��ߞ	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	}�o�P�%	By�%	BP�%	BP�%	��P�%	BP�%	BP��}��x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'������(J��(J��(J��(L���(J��(J��y�ޟ��.(�6*,��s���;Eӵ.�<;�Vgn978�W�� mA��{g��b��6u�Fl
i�5�)�8�0�3��LgͰMԑS����r\l�+�i�m'�Jv�׶ܑpn��"����j�7=u�:�f�L�l-�`e{��ł�9�/1�շ/ksX��E�;{k	\6��UJ�H�cn��gOH޸�9ÞA��gt"�.a���e1X�:�әM���j�x��n�=r�3�8|-��Q�z�u?���?s*,���?]�۽�w�n�m��%	BP��%	BP�$BP�%	Bf`�%	BP������P�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�w���P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'�����(J��0J��(H��(J���(J��"��(J�w���P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'�~޵��Eț����				y�%	BP�$BP�%	Bf`�%	BP�	BP�%	�w���P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'�~�ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�����P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�%�����P�%	By�%	BP�#�%	BP��%	BP�$BP�%	B}��C"LI R"ԋ�				D%	BP�&f	BP�%	�%	BP��%	BP�'�~�ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�����(J��"��(J3�)?�VL��"��(JY�P�%	B]�����(J��(J��"��(J3�(J��J��(O�o��y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%
�Z�!.	�Cr			��0J��(H��(J����Q$��(J!(J��>������(J��"��(J3�(J��J��(L���(J�l��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	B{����x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B{���8%	BP�'��P�%	BD%	BP�&f	BP�%	�%$P$PׅizDA!��q�!(J��J��(L���(J!(J��31
R��(K��g�(J��0J��(H��(J���(J��"��(J������(J��"��(J3�(J��J��(L���(J߿~��(J��<���(J!(J��30J��(H��(J��]��y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP��� ��Y� K�R8�f8IY���`[6����g�s���v犹�Tطh�oǻ�"�vɈ�$�'�				=���(J!(J��30J��(H��(J��������(J��J��(L���(J!(J��30J��(O~����(J��0J��(H��(J���(J��"��(J�w���P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�%�����P�%	By�%H ����l.4h�@��)I�߿lyѴP>+�<��~����)C�����)�}��R����)��F���"pU��MP���\R���߻���d���ߵ�)H����Vj�5C����a�Q��s\R�����ly)J}�����)JO;�v<�������┥'�����EH����
�T	�^�wIJQ�#�#��߿�>�R��߿��)J���JR����ճy�����j|�iTQ(�"�u��x9Y�!m�U��v�2 b��0㺠MP&�;���������(}���y)Jy��wT	����k$��Lp'�*�)Osﻮ�rR������R�����8�)I��ǒ��s�;�4e�{��z-kz┥'��wC�JSϵ���H�T�C�ӥ�-)����� `������R�[�;��ht�"�`""Ē0��{��R��!?}���)JR}���JR�Ͼ)I��{��)ކ��M�$mB�7T	���s �5B�������߿��)JN�����R�;:x�zހ�^�C��C�L�X�0���$�ezЅr�v�2͈��լ�Њ%$�"c���j�/{�j�Oo{�%)N����~e�JO���
�T	����%ț�F��*R{{��y�)����qJR��~��R��}�u�?(�b�����Y���� J�jF*�P&�o�i��MP%=����C�X�O�����)>���C�JS�u4tݚ7�l���Z��)JO}�v<��;�}�qJR����C�J�0�2A0�uT������l`�Ff)���i�JI$�H�P?ms�����)I�斎��82��U��MP��c��JR{{�t<��;�wۊR��{��Vj�5C���b!��1$�r����b��v7c��nrvζE���4��\�W6_]&[5�{�u�o\R������y)Jy���qJR��{ݧ�B�R��;���P&�+�;���H�hG#f�P��^�}��R����߶<��<Ͼ)I�����O��%?~ua��)6F�n+��hws`�5@�<Ͼ)I�����R���}���hg�nF��)#a�f��	���┥'o��C�JSϵ���?��=���JR�����V�L�����j�4<{�b��j��k��)JRy߻��)�}�u�)JH���(�ʹ��	&c4,`j����6f��-�卜,q4X$��$l��l7�v����f�`M��f�4���LH ���ј�HhY������Ї4�M��1����f9�Fa�XXDba�a`X�E�1�a��Xض��caa`IFŁ����fa��@L�(H##���@�=O@OA=0g���M���0 �O�Y�y�5����л1���Æ�AbiCS,g =������D�r!��5Vh,�Fm�HZ#[cs�f�4N�bX٣0��!+�P�0>7l��xak\(\�ɋ5�$X�93��f��V�f9�4�&of�bi��	�3�5�2C�`�6Y8�Y�D�Da8���� �"��XX�@PD��nu��l��y����  ��&��6ke��63xh������[��DP>�a�.e��9���{��UYF����Q�8�,�v\q�zzq�5�:=X�mۅ�'k����2>0hc��ᛢ-M�X�'n�Ѻh�&[ם��F�sқ.��cnݽ��<^�u��,g��68:�bx�����îx��K�����v�ݽ��9�Od�h)����-]s>lu��"m�t�xy��.w-8�Խ��$��*h��7n8,������1�C�lS�gWFPr^�-϶�*n����H�:9,����U4��v�h��Ω:į���(�(�M�9a��V�^�nɍ\cV@f��s`E6-���^i�ٔ�Z�v�eJ�OCJ[+W=EHJ[�7Y�ʶLI�^$KRh���!Z�`��]U[W@\��FO<nHm���j�-�R�ݔ�֦�p觞6=�S���Ȃ���J����iR�<���9	S$W;�q�/G>��8�K8�T3�4G]:����w��^�3�k#<6�xc�fse��:@�:B{n7h8��b��s� m��/.:9n.�q�e͆�m�;9[�sHO!�Jr;�'�z�����2FŎN��:.�^������/Gm\3������I��V4s�����2uk.��lE�5�.�^��ئS�E!��6m��-V=�WL	���.ʉ��j.�ll1F��ڰ���n|t���F�۪��+�L�)eUs�um`�ڹ�D���6^g]<����qΐ+�l��l6�^e�ڤGU�ouȹ΅�ܝ+��b�=J]�g9�&�ڝ����s&""D���s�Y@(A1�pQ��%�L�qٶwm��֙r����˅xvBV����\�]�2���I-1�V64ke�:�d��ѳۓGY�����-�R�T3nX.hv;ٞ�v���n��S�j�m���:���g�@��v�v�JY&亗�,v%�n��zW����ѰX�Vwdh� ۓ0�
�����������@9�n�ӥ����\��s\P&䜥�|[goߨ��:f;����S�0~A�@~ء�E5 ���8�爏ފ��_=����-oz��a7��:��3��Eϙ�8C�ѷ�5];\��t	K۱���Wf��\m���������@$��b h㓮z�:�0�ܺ�3���H�뫷��d�÷nw&��1�qۚ��v����ϰ��CO:��;b���'V�_V�ӱ�A���kn�N��'NՓs�n�F3�-WbH/<��a�9)� v��j�/{�����90fw�}p���Fa!v�O:���l� � �Z�眬f&�36k7�f���R����s�R�>w��y)J{�}�p?��DCR�����b��j����c�BbG��WT	R���ݏ%)Osﻮ)JR}{�t<��<�]�qOȋ��'o����Z�o[3v��oc�JS��k�R��^��%)O��)C�~�ǒ�T8����08d*�wT	���}�JR�}��8�)C�~�ǒ���b������)I���k�o34o{ތ�f���)���s�R�A�����)J}���qJR��~�ǒ������:�BGc�V��C
�U\���81��Y'4��	[�֤��O����G�u��ʙ��z����)JR{~��%)Osﻮ)JP����+y)J{�~��R�Csu5�bm\���r
��g{�\� JP�����)�u�s�R�>w��y'����~?e�ۄ&H[�F��5@�Y��U��MP��w��)J��v<��=Ͼ(&�32G�� J�q�*�P&�yw���(|����R��;��P��
�(��f�Vj�5C�kJLm$pFoY��\R�����c�J'�w���(}���y)J}��u�)JO�{������ݝ6�.ٓ2���^=t��kM/En�Z���v�����{���o�J�
DInA]5@����wT	���ݏ%)O����	.JP��߶<5@�����D��%(�%�j�!�ﻱ�)�w���(~����R5@�3%�����43�[�I1$�3y�oc�JS����qJR����C����LL<)�E6rR�;��JR����JR��k�k#Zћ���-oy�)��;}�������{�|R����wc�J�/߹���R��4>��*O��q+���R1\5@������)JP�߻��)���s�S@�=�b��j�x�m����&�cݝ$k�;�nٚșqlO��U��hi�{r�������T	���s �5B���w��)J}�v<��/~���j�43��9MP5RAVj�*}��u�)J}�v<��/���R�>���y)Jy��Z:�kzٛ�����)JP��{��)�w���� 2���%)O{�߳�R��Y���$��"$� �5@����c�����߻��)���s�P�� pE��!�7ݏ%)N�_i�[-��7�����R�>��v<��<�]�qJR����C�JS����R��~�����Q8��g9š:��E�y�F,ce�з75nz卧c�7 =[ތ�f���)���s�R�����JR���w\R�����c�JS�@���(�$h"��MP&�Os�'�I��;��┥�~���(�,]P�(��474�O�&D�F̵�އ�JS������)C��ǒ�d������)>���C�JS�LXݺ����6��5@�]�df��<����)J=�v<���*�^y��T	��ѪF�jFJ����c�JSϻ�R����~���R��;��┥��ݏ%(D�wdw�Vq���9shr#!���ݯoj���;Yz����m�0ft< �#��ؗ�w&6��\u)����Pe��\�KƭZI�ݼ���k�۞3q�.�	-�@�0��#��vL.��S�đa|q������d�ñ��O�}�dyZ/%�$;�y�'E�sV��c	�Vq9���u�Ӟ��t��XeΨ,�s�Eh����c�nR�ז#RJ;�H�%��7m���2�ih�J�3��3�a��ٽlַ��)J�����){����(}���y)Jy�{ÊR����,�F8���b��j�����)I��{��)���)JF�z��4?Q�P�z�Q��\�%���R��_~���)�{��R�����py)J}��u�)JO�˺��8�18�Y��{2��j�O}����������)=��t<��:t5��k{����l┥'��{��JS����R�����JR�w���)JO�*{�w���ڦ�Wh���Xxok`�)Q]ӥ�s#)kT�J�
��a����u�����ԧ������)=��t<��>�wۊR�����%)O{}����֌޷�ֵ�o\R�������E?��h]HnS��o��)JN���%)�噎�5@��P'$�(����%)O���┥'�������\R�������R���Gr���[5�z޵��┥'�������\R�������R����n)J	�$1���"e8�Y��.��┥'�������qJP=gs�Q�@{ѻ�R�b� �,��3���K��r��F�܄]9�Lss:SN�*d� 1"�@Kq�P&�C���U�)O>�xqJR����C�JS���h{��l��������*ʔ��w�8�)I��{��)�}�u�)JOo{�%)N��w��kY����z�޶qJR����C�JR�﻾)L��D�_ �	�	��Ɓ�<�Wy�C�JS�����j�4;��>�LB���A��JR�w���)JOo~���w}��)I��{��)�o���-�z�ky��JR��߻��)���n)JRy{��y)J{�{�)JR���ŷP\�m���[*��7<����B���4M���jE��u:b��e�璔��w}��)I��{��)���8�)I�����R���]�4u���l޷��{��)I�����  O~�v�����/������)I�]��v�H8�R(��
�T	��ۺ�MP&�o����w}��)I�����PMP�?2p�FH�P�%�j�"�ﻱ�)�w��)>�;�JPH��|���"���������j�43��OBA1#�(��U��e<���┥'׽�������(}����R���]���-�h޶v��e藇BV]�3�=k��6n�d�)e�0�m��j������{ݷ����t<��=�~)C�~���/%��v��j�43u
~�LB����Y��|��>�����)C��wc�JSϻ�R�������O��%=������wT	���f�Vj�)���)JRy}��y)J{�}�q�MP&����␧q8�f�O>�xqJR����C�JS����	4�+ٛY����)1����k{8�)I�����R��>��┥�}ݏ%)O>�xqJR�>�����]u�Nu�¤b��a��gG<��s�W��4�s�:3\vu�H��خ���ܩ�M6�V�]�vʥ�qh�h�U�u��Eۥ^7�Λ<����ۇ�ܗi��c럽�x�g.:9�[�a�燣��L��&)�x�KE��[	���GS�����p�Y1[�g[X7+�3�N���F:5s�muR��z�,O7L��	�<�%�2����xo��Ӹ�x����z]gnL��Ӻ��עD���vL�,
퀎�r�9��"h�~���)����\R���ﻱ�)���)JR}{��y)Jw�飵��[��y�+Z޸�)C�~�ǒ���w�8�)I��{��)�����)JO�˶�/A1#�(��U��MP�fX��M%'׽��a�Oߵ��8�)Y��Y��`$d�m&\�4{8�)I��{��)�����)J{�v<��<�{ÊR��v���Y��p���k7����{���)JQ��`w�����JS����R�����Ы5@��y�q��)�!lH`JBQ-Wu({;krb�������5�-��-�hN��������wT	���{ �5@������)JO�{�%)O�ﻮ)JU�<�)
�B�-��U��MP�fY�=C@x�̪~|E��H}~�������C�2S�����)JP���Y��(H�xd	=$��rn┥'o�~��R��w����+�����<��?~����)<���6R8�D�b��v�������qJR��߿�<��;������X˖���NIJ4�X۶`�LWmx�Հ}��'�q�Rv��복k2inĴ�]s>�kn�sm�El�Z�1��.�1���H�q�'	;�4��k�-v� ��0�
\�B��$��`�ـZ�X۶`fe��)#�to�)F�iI8I��������w|���@(�$h{��T�0I0I̓2�$���� �	" *%�`���!�U8H�30@I#���D�敋�C㏙c1Ė<<;�ce�E�RXX��F��,�cŃf�Z,PAq/��y�X�cfi.�7����6�����z�����`)��i�$C!K12L�M�!¡�#ׄ@�3�s[� �ͳ,^|o�Ĝ�&"��X������T_Q@ͨ>��hE� z�_	�G�1 ���T�O?�+۽��U}������^���8�8((�NH�����-��}��d� ��7U�w�ؒ�)p��L�)��fk�`nف?
�=��(`��"M�P��1��k���F4�e��.��`Vm�uI(F:ܝ�l�eА5�z�u�'1�+$���7� ��~���O�;��8�%$vI�v����m����� �m� �r�D&	�H����OW���9�0��
�K�7]�w^꿨$|�Ť��L�0��Gd�UR���Y'�7]�}��VKM
��P�Z ��ߝ�y�#�P�˒F��$�{1�'�>��o~]$����'�ns �A��ls�h�>'?>?̒(/.��}<|�xJ�ք+�gO1CTM2�����j�������������d��{��ݽ<$�_y��-�G�A&Ԓ8����G�T�����>[���'��K�
	�¶"5��7�<���|�ׇ��~�?$[}0V������$'�nN`qu�y��0��������^4�q8���{l�:����^����^g��WȧD�������;gt�+�=fݙ0Ou�m�<ñV'W��]cv��!�����{p�e	zf�eQ�x̪�e�&A%���2 ; v�=�Ji�)�ݖ�pv�I���d��^շ6ہ;�<�$ؔ9$�:��m�C�F�7�%��Vv�x7<�T�z�7��k����z\�ݖ�H�9��K�$��)�0ݵN�ѱ�P��i4�+:n�@$wg&���8�e��m{/sv��:���9�䞄څ���|�'���(�$�
�����嶿�|�V�� �Q{�LM�9RH���� m�`]���� �Zس���$�p�s 6�0'���Υ�w]�}��I�3�(�,I	�$�?���}�N-�vI�s3��ـ}�6��ࠓj6�x�k�;�s��ـuv׀}Z�6��U���J�h�H1mrIQ5d	e����CJ��K��Cs��Ke�g�������������^��o=Z�EC!��ܐ�'�3���@^ǣ��Kw��;�}��j�K�2r)#�<V�x�k����%�٦�'7vY'�fd��&"�0T������w]�{�4�$�3%�|��vI���Ȑ&(�|MI#�>�S 6�0[���� ��[���8�' �,v94D`��
��eoH�hx�����n�u�[4�~��r�I$h�C �mx��vI��ǵC����6I��w�)F�.H�Iř��*�G�$�۶,V׀}�6���mFӏ ��΀�z=��G�|�s�1gs�=���A���-����UT���!W��uv׀j��w�7[�
�N7'0�ڰ��������$� ;�V�����$DC�T�fWp�y��x-����K�:����Eٱr��I�Er/�7}�un׀w��0�ڰ
�m�����"�0RL�v���9�}�Հ� �6�I((�|MI#�;�s���X{��$n�� 6�L��
I��I����K�7U�|���{�d�H�X �@
B�P��X�Nf�58HJ��G��ȾV�� ;�f�ۜ�>�i������?8n��{�1����>�|�s�;����ș�k�lє�B��m����i�Z���o��ۜ�>�j�:�k�>�x�g"Q���q8��;�s��k�:�k���w�7c��N7'0V׀uvׇ�?$_{� �<`.Ex�\jN�8��5n׀m���`�� �r�?	���`��O�2Y'@(wv��w]��}�uʿ ��$J%4#��*JJ\ß��ͻ����u�a�	U���q�nnxck�st��7�	����3Gm�O'e^=����t�wC�4.]��9�p���ۖ�OD�%�PP���X���l�5�K/0#�6���z#����z�6�$���qU�mҷYK\��P�od�q��Q�ݽ;��̝���Ңܺc��Pm=nnl��a�LŭT\܂�،��毾��6bV<V�*2�vn71�|]tl�5�Bܕ�Ty����N�lN��U<B��mϾ�$�*��up��3]�O}�I����I�&I$h�C �]�=��[�o������+����H��9�Uo� wv���`k�`ӛ\@4�M(�q�wl�;v�0�ڰ{l�>�x�g"Q�'q8��;v�0�ڰ{l��نߟ��to���i�g���Y�z�0���I�i��lb*�,��gY�ZHV�S����v� ��0��`�s���\t&!��$��.] nwM\\{��$�� �ۜ�5[^W-��� 7q��`�f۷9�j�� ��0E�(��$��&��;v�0m� 7�� �l�/;��:	ĜRF�"s��k�� 6�0�Œ~(
�͢ƦT0���b�u;�.�DɵN$er�坄+�00ک�6�Ʀp��7��Ⱥ���0��`�ꋋA��H�t���4�i�)�3@b�R��E��� fwMz�,�J6D�&��;�s���Xw��ba�ޑx�2���W����*�뱻�9S�N''0���{l�=^�;'�@
ۛ�d���^��E�8BAI om����������^n��Q1p$j5!Ƃ�ѶR��Dv�p]�����H�73
��꽤��q��`[���S �m� .�kV�)�"�$�������/_r���1n��H�}���E ���9��� 7v��v��e0i�s�L$��pr/�ջ��=^�;$�d�d�T.�
 к9U�BU rz�Y'��b-�M&�m)q�[���L�v��k��~~o�Bz�-۫���l\�xOq���gqVS�bh�r3Q��+���]L�m��>�j�*���v���X�IȢ�j7$0�ڳ߹Ă��j�� ��L�ͣ�؆��	�X�������)�}�Հ|�l��|� �ݯ ��LU���[�u_zqFH�	$|Dn<�e0V׀jݯ �mx����2�%0�@�æl ǁa�Gv|��E1D�AD��LD����$DP̎�<F	e��X	 ��d"��efY���d1 '��' �I�$�OA="&BY�XH �`4m�-�LZ{���� Nxz'0���g�{�����`I�!&cd�P�3d�5$��yp{�j�w]G;�Ȅ8A�����"A�� �j�v;�*s�sΟ�CI
*s�h �&A���|�g��ͅ�Ȗ�#3��swqF��n�
�U�]zU�+wW�k��.�C��]w;�+@֗<d����=�]�6D��]�Z�����������q<�L�]��m����n�N�������;p8-�ϭm���9�uu�[l/=�>5Z�L��ۮ2�Û���Z��v<lz���n)���s��9.��]��mh˜<�\��g�vC<ݰ�<l�1�l#j&Ǝ�ṰՋ$����Vʉ���2�e6v�F@�.Xq�6m����t��B�b-�5��.!{]��=�����v]l�z�I#�X�@;JhH�M%��Hֳ@�[&�]�/D������	U��G1ZZr�p��n$�]�%�vq�8���������]U]]*Խ�l�T�<��kd"Ӳ�m�T�x��5=;v��řx�r��U�ų�1WM��D��,�����~��ֺNz�h���F���wN��W��wX;zU�E��ȼ���=�vs�c��8�C�ez��ɠ�Vz�'ř�U]��em۶�-\2&�M>�'\q�{:�f�9N���!�]����j0R�p\�Cb놵u2�$u�O螧��=u�ͩ���|�l���L��w�b�,v�#�U��:�b�<g'��q�w8�f9�ƨ�j�rE��6K�.'vo	�e�.Ћ<Y��-�uq�;J�Zǆn���QK!5������-�r��Zؔ�;�6���{D@#v�).8W�b�L�ڞ����I��쥏]b�k0���,t	��m�J���HZ�5=��v�K�Y'��"[��nA���z@\�K�����m��Nʓ�I��L�<�kinA�u�B��v�����cn\ka�=t�C��`�βуe��S��
��h%�{Dvv�j�83acss���qlZy2m$�����s��rL��y��^4Y�s��h��<�줚9����8��]�[��b�n3>�.��T�0G)'��
"F��y�t2��KǍνǿ�!����
zz��ʋ��*�*:^�+������H�?e�}�4Z�kv�o*�������6�9�TI�-�yպ�n_��|}@mЖC�F�;�v*��=��M�ാͻ��9)�͹�0F]���E	<�a��>I�9��C���`*^�\9.���mŌ�;;�+W���֋Jvx)z丱ceMuӱ-�����s͛ڳ��q�bݛnG�m+�s���ۜ�����f�^ݸy
Nզ�'����׻�����1Yb���9!	qՋ��G.�l�h-OTWT���A���3rR���`���jݯ �mx��`��y��$��H��|�V׀}ra�O�f;�
��ӑ���I��m8쓋w]�y�0�� �n�N,�xn���%'M�� ��LU���k�5[^ݪ7cQ'!�Q�!�j����+���*���������L���O�QA��L�n��0CŻ��X
����	�tQ�]���\�ʓ�#NG�jݯ �mx��`�� �ik��D�>
G�m�@��]�@W�*�d��d�^�vI�������i��$�>(�� ��LU���ـm���9gq9��m�9s�8�g����ݳ ��Lio?����cD��.E!�[��f�����`n�>.H'�+�R�	��x94vL�sV���b+�Y&����y-Ƴ�vr�J3��?��� ��L�e?��� ��<��'�"(����NI,��Ɇ�
�����d����ݳ ��rHB)ƣrK�y��*�>�����(~�B�`àB�� �D$}����}s@^�?�[|�*d��M�d� X�5�'f�?%�٦�=����WȈ�|� ջ]�v� :���Owf�$�{����}�=l��m��ݮ�a�޳�����	õ�Ism�D�1�ݝ���,���\��F���{9�}l���^�v�;Y$ԎB܍�"pY'���UI[�<�|�ݹ�ie�E&D��.E!�o��[����[����zx�>GJ4X\iFӏ����;$�slY'���j�@��  F�����QP�q9�L�ns ��LWmx��`>ݰlQ�4�8딇��<�1�6�Z����vQb�%�*�0�S��r\5�m�_����m��� ��0ݹ����dR	�l����{UT(PH���d�{v��}l�V���4@�F��x��`��=�����O��� R��V|rH��nL��9�}l���^ n���V�r!�k�9�.��� �����*�� �ۜ�;���;��q�A���"n�G'C���z��aGl\���Ca�;۩��Upk��ӡ�6�<c+צ4� �1�Ӝ ��6)�vͱ��?����L�����;��]�fجm��k����۵V����q�h��D��n�N�ۘ�p�t�#��u���˖h$�i�˞�Mp&-��
�k��:\,n��e���N�r!�'D��l��QI"e/P�G�+����լ�.��xj�ݤ��u�~��&r:J��&�t�
ZF:"����MR��[��������[�������ќ��"P\#iFӏ ջ^�����`��6I��c���ƨ�p��r7$x��9�}l����V�xv�Ҳ.��Ƨ����`�k�>^�;'h
�ۛ�d�/������&�j� ջ^۷9�}l��o�����k����C6�2�*uv7U�cm���U��BЛP�٬
Q7�k��rA7�v��ns ��LWmxKD�x�|rH���xn��g?��*�c�}�4�'V�$�{���#X�n���\��`[)�j� ջ^۷9�m����h�7�Ȥ>����v���9�}l��6�0}�IKiˠ5n�?����}�� �� �f�����P���VMh
Rѥ1���7	Վ��Euf�4.�RqA>E��'#rG�w��0���=]�{�N,�w�T��ؙ["8Z������zx�:�k�5n׀w��0���5��#8�� w��V�u˞(z"4�x!����;�� ����X�N禛$��/`&#8FF�7&�v���9�}l� w�� ��>;��d��"7�ۜ�>�S ;�f�v�c�TqÎǌ[r� ^;fd���1㙌%=-�i<ڀ�f�����6��S�������S �� ջ^�ۜ�6���O3�D��.E!���x����������U���CLJ6�x���������Wmxݰn�RF\NF���*���n�Y'��M�{����u@y�"X"I��?
F�(~�� (�'�vI��&VH��N58ܜ�>�S �� ջ^��X�O�P��e!�6�)�Ȓ�IM7[$*�\��1m�;����ѥ��:2[��p��H3��|����v���9�}l� n�o"B�'jH&��5n׀w��0���:�k�
Z�㼍6I≹0������Wmx��`S����P�RD���� �m���`��h��F�8q4I��?�7}��f���9W��{�UӢ	���=�n�%q�y,�m�zȷ=R%���n�){[����u�Ý�r˶0�`qm����E��7���6[��vxNIs�C��Y�Q��Ywz����]3ЕZ1�yNv�gK셮]�#N�-�$��F3L�;��b���љ������Vװ7`r�^n��c=���4��7=V����Zn���F����{6��k��@�k*��U�`���8�3$�,��u��>��;��E�MŬ3�]�FR�ENk`�8AD�IDӓ@-���;�s��m�~���L�~�Ȕ��'"rI�w��0�����`wl�6��y"��Ƨ���mx��0��`����t��F4�vN����d���,���X�tUP�� -^^Q!N�2H�r`�� �5ws�1gs�n��t�G
+6�c��ĝ�v܄<@]q�j���i�Ly���狲b���x���m����@Ż��Ś�[���B\>a$���Y�޶r�����(mBT���o��3Y��w΀�/x]�iϿa$o�?�վ��5[^۷9�j����x>;�D�D�m8�V׀v��`k�`�k�7�*HH�����nH�ݹ�U���k�5[^w��p8���B��q�'f����>^� �,b.�)qr��עjdnD)S�N''0���� ջ^۷9�uS]"c|j@�~M� ��^D�[��m�`[)� �
p���A7& ov��ns��zl��Va �0�M$LFF1%��.��,I�PDLDDD�PQ$0E0@�4D���#�$��!	a��Ye����Id��d��OH%꘾1�P@K�FIG�'�d8ȐX��:��	ٽ<�C�|�|��[�;��򙀍c�EXf!!M�=����k�!>�!�� b20��th"�*ՌL�Q��!�-B�X� ���i=zE���>�96�9��NHl��3Ek5ѷ��;�2��T2
'����T<TG�W�E���; �!�_���@1]!�O���1^��P�_���D�}���'N�l��đ��nK'@����I���d������ �6z�6���>�Հ�f n�n�����7���֤&��Y��ڍ�*�.ۊR�Vt�Ɣ�d�w
�%�WgޖiХL����@��@goT~�{��>��uj��qH�Im4��ݳ �ۜ�>�S 7���?s��7}�	�F�NI0��s ��LWmx��`�Y8܈R'��rs ��.�HY����K������ޏ_�y�K���FD�� Q=@UW���}��$��:���A���>M�v�B��4�K^�;��սP�$��Wi%���,NA�%��}���cd���]1W>n�;f�8Ѫ�vv��V���9#��bI-{���Ijۜx�K�r�|�B�bI%KSc�bq3)���ݤ���I$����I!gW1$�����$��$���M���:I%}���I;��I-{���KV�i$��8���h�@��}�I���$�����$�oT:I%����Ic�x�24�I#m�㘒K]���Ijܰ�$��f.q��d��I��U���T@P2��ҤH$�a(�`���v.�zx��99��Z�m���5�ꎳ;.&�eh��i�����γ��x�6&�'��R%�*қk�/=c�.�f�ɺ�p�E�bc�^���sF�D�{n�9J& Y燴Z���`t"���ݷlPnzn7''E�M���=s������K���eb㚹�R���+L\/Y��M�TN�)�A-�$�,����(!�UB���'���i("CA�U������<llZ1�,n'p�zQ�^\��vsk�£D�nF䏾I/���Il�}�I���$��_�$��Y8�����jq�8�$��j��msIk���I/y�i$���1���R�8�Iv�1$��k���w8�$��j����lS��s�M�1$��k���w8�$��j��K�ɉ$�{Sc��'�H���|�[��$��Z��$��d��IffNq$�2@�t܁��� 4�]a���5�K�0����r�[C8p.p��<4)���������~��dĒJ�g�!-�q�K������H؆8�Ԓ+ۮ_@ PT0U`P	@��e+�l�K2m�i$�&b�$��LZ<��1��M9'I-�z}�In��X$�����I.�&$�݆���B&܉�'�!-�q�J�j��m�I+m�|�����<���q�nDx�Kvn�q$��c�RIffNq$����ڪ�34�"e�=�wVG��9 ��{[֏m�.�39���b�d�Z1!	�r.���얒I[l���w8�$�����%k�UȸN�1�LI$��`�ՀZ�X˶����|�M�i��((���^�������{������˴8�A�N"���C������*������(��M�9h��-v���^ [l�;׵`K����"�6RE�OW�]�UUP���8I��j��V�;�(����"q�����WMn�zK�mי��k�a�i�yi�3�&m�GO�� [l�;׵`�V�� �f����nF� �^Հ}l��� ջ^ݲ��$k��")��X��`.��[���yP�6t��53��ܔ��uʾϾ�W����+�`���W�&�
y����ʽ��w����b��7.�Ż΀�{ʀ��΀����?U�ޑ)�K�"F'0'�,�;$�ɮ�@��c���s]��J#sMutM>>I��7]��>[k�>]��wl����Cm	ț@G��^�� ;�f޽� �����p1�I#�� w}�ݳ �^Հ|�׀}�Y���o�8�|m907�k�0��X�mx�m�����j7M��L�{V��^ }�{�U{���*��X�N��ެ���=kE�˞d�g��M���۞�:vwv�B�s��q�q�6�I�b��8lGh��KV͠s�D�I��X
����0���Q3�^lN�M���68[/�0m�MS�n��/F�<�Ѱ՛9��ⷋK]��2���40�,�����-r�i3���[�Ӷ�+65��$8 b"$*�I0��n-�kR�3�Ny�Z������
���
�@矱2�%�g$o:�k���V�uπڛ�3F��Xꔴ�"��蒲���9b�i�o���l��ٜ�{V�o�/=.7'O�q�wޘ��0��X�mx�8�ȸN�~� ;�f޽� �m� �v׀UK�g���ADܘz��嶼��^ wv� �J�n�r&�ŀm�˶� �l�:���s��w�<�g��O�s�Wci�ퟯ�,��if��g���ܝF��5�ʩ,;���g�Z��I:����vـuwk�~�>@o��=��n5��m0�q�'�َ��x)�d*%���(2!�N~�!��< ��� �v׀]fԤ�D�n6܏ ��׀�� ���V���aLrr")��x�l��l�5m� ��׀m|�>X!q�)Ɯ� >� �mxz��}���?
�����2��('����t�������$5p�b4�j��xnm�p�$#�)'�U�y��ڰm� >� )tu�'��"�jI޽�>H6ܘ�m��k�>Z�x��cmI@G m�`ݶa9+�@�<X2�o��r�{��`�g�fD�$��������w����k{�{������9r�p�s4-�t,�t��t}̖I�혴&�p'��!��.MV�7T�6�m�j��Y�����<�E��q�$����V }�fջ^�`�"i�NDH��X��Y�z ������@f=�@r���KK��NB9�� �ݯ���`k�`Q�Ӄ"	��#�����|���*��*�DDA~��(~EP� }�{��W�Z��y���E�L�{V��V�� ;�f۷�2rrr$�$��Oʹ@�y,���g^;x�P%W-���j��'���*�e��T��T��t��?�""�>��VI�{���l��n0�.E�L[�ο{ބ�{��u�ʀ�}ʀ��P�q>8�i�4���ـw�j�>�j�>]��kV�$I)��ӒL�{V��V�� �ݯ ݰ��&�RB���"�O�f;$�  =�߿kڻ��f���{�r��QTW��QTW��DU��U�TW��EQ_�E�QE�QTQ��%�PE d !�PB �PTBFP	Do���*���
*���(�+�
*�∪+�*���(�+�@��������
*���(�+��"���"����(+$�k%��@]�k0
 ?��d��,��@    � 4 �            ϨU @
��T�  )%!D��R� J�@��*�Q*@� R@Q  �R($�       T�dh���RŜ������\ t��z���}�ӓN���p �7=/���{rk�  l��+ӗJX@9ҙ5��{:��o'Jdһ� ����m��z��Y_[�=7� <     }
�@� ��n-糧�q���J��r��#�;�5͗3���p ӫ�k�9��דI�,�{����b�Z\�v�6W..R� >����ͩӓ�[�v�� }�  P �*�l =�����q9:��y��� >��Uf2�Z�Ȳ� �{r}�&���r���=:� �9�N������|�2����} <���w� }�  2  �j�m���( PU  � ���s�=��Ҝ�N�&Ϫ^���./�{����J����W�r�x#� �
2(�0h 
% �h� ��c �@� ��Pbi@�� � 4  ;�  U  �Y �D�� M 
1 2 �0 hh�@� �  H�`�}�f��;7=�W���zۋ��m�[+l��0 �wRVO�=�������'�� =!SoJ�* �T��5M�UJ�� D��J�Rh�F�D�*�&�J�  ?�%OmT�$1 ���&Ҕ� �➢����?�������L���v�;ޏ{����AQ^����(*+���*�(*+�dPTW�AQX�(�����I%_������?�����0q]|c$�ĄR2H�E x�R X�1SV�qH�ׄ��I�54+
x@�3	�)� �R�f�%R$t�@���).n�^��l����T���?=���D�zYa'�s�$q�$6C�Sf��H"�CAW��M}��S@	 ��vB�y�|<!$$��52�]pI8J@��0�JI%���99��
�<�3̓�a��2�.f�����?O���?���OJ���\ǃ�!�����e�e���o<�!syM��y�5��_3^M��3��	"G������n␦o�O��a��K2�p��������$ ĲKRP!?o����NZ�$jd��$&q�BS4���F4�Q�45A��JzT�H���8V����Ar3-�Oxt��%=��ą�H�!p�7<9��[�y�ʗ^B��z�Ɔ֩�荤�����涘ÞDŐ�E:$B�+ ! �  �b
H ��"*BE*���  I,���(@���X9E��H	� �"*�����@�H�,jL�Rd�����Z�`�X��T!��#
H�	D�c���P2�S�k�J
I��;
����9rH�&]���#�K$k!R0��Č�HT��$<�B�X�#�����Sl�0ɕ�сC#�:H�Bᧉri�	�9!	Õ��H�䐸:D(f�����X��2ۍ�L�b� A-x�Hp�FK��H�0!\	r��bY�I	72	d�R)��.q|���o$$d!WNJBf�X�p�FJ�:���LuHC�P����#�!�*L�x�,خ�
����!��FB#A�S���������}�!O�F�
������#S-�\p �HT����P���``��©�A���0�"��4�p!"7!G$-Q�P!X�0��))���A�B�8$+Ё�e��mXA�5��5�a���N0a
�FB��9J�jK�.hK���/%a�З^Go
������b�4!�R%pӔ�1�L0��%	t,F	
WB)\4�5�B�HD�I!D �%|=���Ng��|�ᄧ�.{����f͟{�&��|�|�]���^��/fI��B��ⰷ7�S9�ā
g0�]�)���J��`B��_#6�����(�����[��w�L���Ņ�-8�Аe1�H�#�1�>�i�bjj���zO8��ۻa!��ß��R6F3YL	F!b@�eIRW �P����ksx��w63�:g$ns@4�$��A��H�!$��"!�ࣷ{�#F�	dI��c��S��u��Cة����U�m�Ѱ�fv��O���XӉ��d�CNB�d��K�L愈?��S�)���G�XB�iU���vp��~0�O$aH�9�"g�.H�	/��c"y�a$����8Ă�A͉���d�1}C�JBQrL�$#HS������Hd0��!��!��� b@�ږ@��;Y�\@�H�	�S0����n�~��@ؙG��Z��7h_�۠ �Vd�y/$4&ߩ������e�^�&$a���s��8���8 i�?7��jf��y�Hܷ�=�z?�{)�H)�)3e������s�9�����9?p�)�Y?�?�����H����G||��<忆��9��t����@������I)���! a�1!]᧾��Cy|'��$�KI�-�Y0������ �I�F������` �� �����L"(H 0�������$)�H$
�a!@0�# �2G�S!�D$��:Lń0<�"X�XF���$�
c�E9��$�!F`ڒ1���,l�!0$a� �%� GI��$Yk�F���0+�ZR�A����M��$nU�a
�hN��:q�9k-(I��8�F�$$���3��"��&�0�#`]98Y�,-
0�d40�V@Đu�9���0��u	�YkF8�a �J��hcŌ!Vq#\�Ip���)�� �� ����N�o �$729I%
y&p�($�
CxxxF���,)�ā6	t�$�k �$�D�L5�\�2@��$-I	L9��$�4�I��>bJBŦ���� �$FA!L] P�cY%�ĒHf�|�CN �i�%!���I�%3��Jpe���\�В21��j���Is��-��:鄏H[�2���w`q9�Y��3C0��*H@���CHB�<m�3&��\7�H;�@�lS8p�e�B,y�\�)�2��qӄ��I�D��;�ʖcP�ty.;�:K��X�i��rH\�_#S�x��¡\$H40�I-0ԁ	�q���s)3x��#C�M����}�s�ɔ59�|��.��z��F $-��D�X�����ٙ����B[F���f���i�p�BLxpX��~s7��B�//���i�xxz���O?0�o//���ya8�j��%<�2�	�7�����7����?��čq��y�>d(d!�u#���S���^d	LH��||!
�p,+&o	�F䆠B��'��
F���H`e0H�G�C��$Jf������ĈB�̥r&�By9��%	C�\�ߠI��|�}��㯀r�eb�'�I*mI3��u�+��<$�Ð')��I����?	
o�$?B�.:p���+����"D�0ׇ��@��;!����<?BK!�
HHD�ke0��\u�x~��
a�'�~XI48@���*I�&@sm/���y�D�-��5 d�|?"��(b�J��(ἑ�S�D�@X�!	# dZ.0 �	!� �������tg�Iz�'I��J��# �CÐ�����?�燛K繘P�u�������1łE�@���믒�����%`4�L͐��V$�#S�y*��.I�	��i
@.a�a��1Vؐ�H���ra�rH�� R$Lb]��sE�ȵ`�% �5��Ŕ�$�D"F,������H���-���@��*F$(�I
0(b$H��~' B�%�p�##^!Z&�1P�`�$��惥�B`��oe��m5�)� �B�?O1!g$����܉!H�0թ�F%X�V�`��;�
1�ӍT�H�Jbi�hK3]x�F�F-�,���9$��	!p��X@��!lK��攄B5HQ�jf�V�A��
�4ז�ĦB㼤JJ`0��HGHRa�pe!���^H�L1��0��iȑ!)�0!�!X���!
c3 �$�C�7�a#
��C� �ӟ�~��nÏ��`T͜��?8:���8¹�)]���	��B��B>)ǒ�9��2��������"D�@? E��	+��ѣ���¢`X�@�<<�	�q߾s��'��̛�{oߘ����$�I   6�    l]��n'^��S��ӡ,���F�(�h$�jmp)"�4��7H���b@;��=N���q&E�ݦ`W�{u&������thv�����ouW]�s��:-�[�gmm�P`�)qr�O/2�5��ˢى�&��[����uA�h�,V�����R&���%�8�ԫI���ltR��Z�r�/�����ةݕ�8��Y]�۰qڞ	M۾�?���u[\k-� ��u��m��i.�yڕ��������A�Z-.�
��`B�j�{:�6Z�	o$��.�   ��I����s�݀rAi�N�n�km� m��ۜ	��lH�n�6� �   n��D䴶��Ü}��	$�g ��@��:0 l� �@ $�b��ݶ�` �m� 9�аÍ�Ji����	�/]3��5l�P�@U�+<�ZM�N�m���J�N�h�	   pK$�9f���`[Ad���t[�pHI�f곐�#�I� ���u�Z��*�q�� Zl �`۬֝%���|m��nM�$f�l��л� .�IͶ���\��6� p6� ��������Mˈm$�ǆ� �o]-��b�_ ���N�j8�Kv�` ���2�P��!�*�����˴ʴ�P�2	$mmͺۛl�\���`�А��`6Z�@�F�'*�yY^U���Z�i�m�܋S��u����  ��-�6��Im ���n�qă�$ƻ~]��  Hm�V2Y�dv[���!�ͣN�Hm��6�Xcm�  [%�k:@ �sGY�6�OP PA\�TU�� 8��i�h6*G5�[M�7�?�m�Y�%��$�k'Kz��d:�x��!l�,ւ@l�m,0�k�L`%[��/��UU.bquY��m�v�P     I�]��յ�� A�i �mr�%�Ӡ��:]mÜ����I��P �J�S����n� ��+Vܤ���̫�S�Y��8۴�$�m��,H�nm��I� ]�/m!��'@ i,��j��YM�V��YD8�^j�@U[UAڦm[m��9'i�Hmt�\��Sm�Ӎ�m�k�Em�� -�t���C������ջ[ך�f�     ���� 9m�  �� �jg���m      n���q��I	&�|����8�jC��h�m��l�  M�F�/Yim�  @ 8[M�I��dKd$4P� �3�  	��m�m�o^)Km(-�0� �a v� $�Xkh ��se��6p�ɹ8�[d-5�\%�p��u,�^vk���(8��;�/'<�b���K�4��-J�U&m�;�����W��v�#�VcAhW�Ci�V� 8�@ Pq��Y�F ��1�"	�=]������� YWk1� ҭ�h����X��a�T��L��m�m���d� �]�n�#�j�B~���U�j[���j�eC����V�����U�k<�Y^b*UT�me�6  7m��m��z��-6�1���L�P)�)YJy�m�&�q�)�*A��BIu�dr��ֱ,�PT
�@K��p%��J����� 6ؚ�����hp�I��;md��ؼ��gt��a}h�	#�p�ݷb�֭U�,��YGjRZ�� ��q�ŵm[%�mXl���h $�k ��   ��j��`���F��)f�Tpj��d9��M���l��#^�gWUԻs�Y$��ţavi>>[#Ͷ[��R��J��D��m2��J٭�azmX-� m��v�kh�D� @  [
�K(Hƶ�۹X�.J^�/N�X�'@���K��f��$�l�[um�      6�f��J��p*��,b�I@�@��� -��,�]l��p�X�B�ۜ�]��d`m4�Kn��-0�J�g-F��5+(Ȃ�
ݰ 8@� � m� m�H�UR�6/��~Z|�X@��k�4W�Xd����	��UR��P��7mK��,��v¦jw�%��R-���"�ʴ�L�J�*� ��Դ��L�T�j7mm�F��n�;,d��[GnL��eL����� Il�͕��[S[u�   �  @6�$ gY%:�@�` �`�jBI-�km�u� ��m�����j�$��m�Z��0�	�@�^.x@6B�h�J�u�_���:�`U]�dsʲ�U@6��5���-��� H�^�$�e[x8���jP+�.������M�b�k�˒�z�g�t��k4�-������|R���� 6�٬�:ڤx�l��E�9YN��(�[t��4��kgS�u��V���u5UO$�pb�[;�(�Ԯ���Z�[�wD�і��.��#���:+K����5UL�@m���<@���4KJ7W]t�R���P (�[\��vƊ�㜰lIW�	���8n���9��(M<�6���I:�m�v�.���Y@ �y��R��e�+�d�[W@yYҭ`�d!����T��t�,������$�荚�P%L���Yy�� �m�oU�]��\t��( �$��d�ܛ0�Ce��(moW��}Wo�[`�l��q�mKnӥF����,l�mT\��U�v7D��Uj�n��������` �!�km��� R���['GA�F�m��XK+l�5J�ur�5/[b��f^ۓnZΒ�ہ�:MVVP���@@�j�ڤ�$��j��X#[ۭ���fͤ�6�-[�pӀ���4��	�\��]	�p	8X6���Q��mf���ɱQgZ63)\�v�  � ��g 	0i��5�d[h[@�f���u�m%����6� ���@ 6��m��� ��@�kn��ڵt���� 	���I�մ VƸ���S�m���v�p��m& �ږW6Ψ�S(sUtu 	�j�a���[0��#Tjv���e%y�^�h6�j�� �ĊMeդ��a��v�l[UU��ʳ��@8
v�[�eɰm�b` ��VULe%��@ s9S����WF�����m[Cz�`�n�ڶ  �` hZ6 = m��� ���    �f�  5�0ٶ�cm� ��� �p�V���m�����[%J�o+n�ŋ6-�Amp��-�mEUU)r�J�*�F��vKm��g��یSU����qִ8  �[}��ky�M� �h   �m�D�I���gR��mA�0qJ� M�T��'�8��v��N�P�ľ.-����8\ʖN!�U��%�J��Z�m������GFoD��3<ҚJ��P\��m�;m�А�[��0� 	   m�  j�  �l   �6� � p  ���`    $H6�@  �� @� � l   ��l �[N    �۰ ]U*�UU*�U]0 6���	t� hlM�N�Pevey[�*(�P�I��ib�(��ZUk��
ڝm;I��t5U�����g�Kl0  m m�  �  �   H�   �Z � f��߁�ڶ�8�cZ��jU�J*ڥ�VB��Hn��.ŴHȶK�u�8�5�1m 5�$�n�$����\��-����5��Wf��UUtt�`ت�UV�p��ͫl  6�  m�	�-�H  -���  �` �   �`m�  8 I!z�P��LF� $�m����+m�H�H�t�%T�%��[J�n]5$� �`k�q�sm�@ �  qm�b���d  jj  $$ ڶ  -�UJ�쵷VʍJ�Q�aTv܁J�!J���U*�2���{YehYVUi�9xq�����j�]�8�U�S+����  p �����m�,Z{f�֬��P �ٹ�b-b�� �`�m�l�h 5�E�[@A&����2�D;+Q���V������\��[ �lu���&x�N)j� ���I�[[i4�B�Z��V8�ِ�-��@s
�R�t�R��$J�{���r�WT��a����,!�S�����z����E��I�Ri�iWg������Kcp�"ruH̺�a��ںM�f�kh��-��;-K��Xlͧk(ԫu �`��uc'A��{f۾ -�e�k[�V�(t�1
AR���xAS�@x��b(UW�b(y� b�� ��@��*(p^)��
 > � ����H
��D����pT��@E���O�bj�E@��E��D�X��_E*����!���x�t D5C���t|q� �P������Tx��T4�� ȉ�����`���1F,B��:�� �� �@5h�q8�`�� ��~E<@ML@�_@��{� � ��@�"1b `���A@:*���� W����US��g��� N*�ꊢAz��
U�C���EEx��⾊R'�PH�V� ;�n�f5D���`���2��t�	2�u��dr�K���5��*`�I��-�`�8�>����e�g@�k���v�s�V���ܒ�Y����l��l^K�D��*�.��v�5<���v�1�F燞�lf��rt�����IpPR�';9�9ŭ�6�)��j��p�i��A���Q�llĘ����q�*j�C���r�N�mت����ܽg����ܣ�YV��J�W�Z����"�5v�F5�bwo��s2�Wk5�Z%%tqa�k��σq,M�^Uj�7`����\�.W�a(6A�ZְVQ�q(Au�����g+�.8��O���m�M��`�mvu���p���÷oWHU��X�749��:c\���d�7@�UV���G/X^�U����<�����&8�����m*��#UT�H�*����鼗��`��&b���.\��;&���l:�cma�S&e���j����4j�����]��4�uǣ���Ӭ��䴬�箂^s�M<��t�+e޸�GC3�H77�[��!�;�1g����[bF�4su6+� ��`��x�8V�;l�\�V��T��^Q�W#(cT�:���������V&���cLr�;�����<��j+v ګn�|��ʰ���Ch.'�i�]��I�P�����Y=9�!����j�*�*��J�<�Z�:xt�<%�p	�(c)8M�(�jBjݪ� C��qWcY��2��l[7it��ル�� �mY��� 7A���l�$�6��kI�V��9�j۴��Վ�l���6� ㄍ�ヶ7<n2Ĝ]X�k;��xȗ���#�VVIki�m������I(pݳBn��2�j�Z�ؖU�mJ���0��۪hݰ �! t쬽P��q.��V��C��D��.��ٙ<tO�`�2��h^�bs֜�Kl�͵r�:�{�����D?9�G�q@1EMQ��HN��Ɨw33f�4N{]��(��%���s��65iν]�����Vnѕ�I��6��=n�j�$���\GG9�2{K/gu�l��p�u�����t ;�n����uθk��Zݻ��P��2�ތ����p2-C���H�;�� n�ܚ��3�g"���29��XY�N�6��sBu�wx0q��$����?}�<qϑ�M�r�nr���l9wn82��m�d������bC���Y���9{� ���r��@�RW��5�������#����)RJ�	���9���׬�:���n8E1�8�����.@yv �s�����k& ŏ&(9&�W�z�[4Ϫ�z٠\�`��Ȗ�Ǡ������� oː�3pڸ�\g��Ζ��tcvB�����K�K���]�;��x�uҵ�����p�]�7�r y�`�_�z8�I��@;�Ϳ3�����@=z��ڴ��
�kp����\�y�������Q~ �"�D�A'�z��]��z٠U�^�u��_�ci���v �.@���\�W`����v���-f��CY;FH�Gӱ�W�ĭ�S���@^�f-F�\�QY���܀˰�r y]�=��ޡ�;1,KL�rM�Z��٠�� �h=�(%B�Iyz��� ��4˪EU*�"�T�*�R�WJ��>���G=/@��CX˒60r�ɠ���hu�@=���A|�G	0MH��I�~���I�~���R��?�߯?�#�Z�g�m}���7�{��[�2x؎)Z��-��oFx�cV���W����@=�� ��h�٠U��`��A)�{��{��u�@��^�u��pm<�"�I }�pܻ o���]�rge�$B���(��u�@��^�?{��$�A��r~���I=��s�)�ǉ���$�*�W��f�}�s@=���\�JA(���j[��S��1�ag���`�5ɜ�i�����LO��8,1"F)z�h�w4�&U*����9�����>e���kwsv �spܻ o�� �.�-�4��q��@=������l�/�U�}�\Pĩǋ#�o349'��נ�٠O�C@>��heG|CW!��L�N= �������zf��/@��P�!%S��6߈��/Y��GoOc���㝺��ڝj�ra�΃N7Pl��c<�yywT�3���Yˉ=F� �8ݲ0�(%��gXy׵�H5�vĜj^�n�gA�N�]�C�	tby�n�z�ݸnB��%���t���6�m��ݭ�wl�p������j��w�}�l�? 1�l2�v��X�6�-��JbSp����Z8�n�l�O�wLm�6f��&�h��]мBu�7�u۝�j�m-Ht;NŒx�pBd�rO������@��� ����4vU#"&5 3j {��}�@�v �e@;�<�X@&ɒɠU�^�}�f�}�s@=�f�s݂�T ��F)�� >W`�� ;��~� �YC��X���@�}V�wu�z^�~���'��;O��]�'oCՒ�P��u)�v�7y݀���{dtc��R�˱_�|�,N<��Cq} �M�uz�����x���,><X����'o�{���(�*�����I��k�wY�U��\�b�1�H��]�7����`�9 9.����Ɖ��I�U�^�{������[4�4vT〦
L29 �s����r� |� {:���L��vM�ݡVs�4��BKBv�F1��,Pv�.�V҈���[��g�������r� |� =����<����1c���ޓ7�U$�w�������f��;�T�hŎE�����3@>��i*�uT��L��٠[�͑bq�LjI��v <� >�� ���SW�]��<Hh�nM �l��l��� �u�sn5�9���6�s$� �u����m�b3\��5��Հv#e`��`�s�qta"S"I�����Uֽ �u�]��Q.��(��8҄rM ��`w; o�� �]�rVY�nm�LJLNM ��4^���hk�{��XF���nM��/@?I3@�/��z�*�K�T���&h��A_�!�@S	z��4�~���m�4^��
�U6���-Lbvᬼ���j�<�g�$.��]�.p;A౨���ɒ)&����@;����� �m���_6E�G�@i���{�7�I&��:�����}V����$˘�76��9{���g�l�9����:�i�˱�0�)�JG�m�@�_U��f���^�u�X1�یn6���� ��`~� ����~�_��������Hm{;��������1��5�p�<P�wr1\���f�pqm�l��莎T�lm��=`uŹ�և�y2��ڭժ۷KW�u�n��\�G/H v��0��M�/2�qZ����i�N덭Ƶ��/���6�o[s3�n[�:9�ȶ�P�bYms�t�A�pp�3�14n�����}�>���2��7�~EZ*�y�ᴙ��ԜA<%W:��f���6���X�rs������nq1�3X�m�??�� ��9 >W`9��=�2�J��HHG&���^�}���}V�wu�{�Y.�$�Na#�@>�s@�/���J�&�;�@�ӯ@���j*���ɒ)&����@;��/uz��h֡|�)$����I�U$��u� �N���G�I�?\�����vt�u�9{TWv�qÎ�9��4�"�I-�-�����l�T&���r y�`<����{��`R��Y�#Y52	8�׬ۙ���Қ޶h���Q*�q��5znf��P�� ��9 <��4v'a��&��� �[4���<��P�FWa�i�x�a�����4UT��~����v� �u�W�j�Q��"m8bGV�҅ҺGڹ�a����LD�g��5��H�LlsnM �m���s@;����4�v"���'�ɠ}����Sa=ݚ=;4���F:�(�S&<JL���@;�f��3{H�
V �$H22 F
@��B@X(��B(� @"�F
H �H����B	H!�B! BHH$B DbdF+ ��`$P� �#`āA�0!"�2$ @�$�b2`I��!�F%��#�#5!b0�B�q =�����1%��2(�
Ŋ$@��1�`��B�R "�Q��$D�$@��#d	�B0�B"H�� BH$�$H�@�HH`HF"�bI$�"�b�$H,F0`�+"�0 BHH� H�I BB��H��B �� �� 2
�4����5C�$ � ���  
��ߓʪID��/��~�4�&��"ˡ��!Ʊ�&�w�� �[4��4�l�.+���D�L�'&�y]�y�T �]����W�w���y=Trp�H�k#<ԡri���t�.�c�k]�A��$�:�p��U����� ;�`yv y]�rSE��1Li9bp��@;�� �m��Jh�;���Bn� �s����9�ܻ �v%�H�1��rh��@�_U�'�������)ꊫ�!���٠_��E\S�$NM��Z�mz/Z��� {�s�h�ЌRWa�h̾3i:��:�p;1��i��l�d	�H_�
G	��@;�d�.@�����;�W�٢X�Ȝ�^���Y�^}V�w��K��5a�P�5#�^� {9��]�7�r r]�ѷ��8҉�&�|�� �h{��[f��Ǝ�dYH�&D����s��v�ڐ~������;~e�WF[�-�B@�l�oa�K�K���6�=A�@��om����YY�&��6� zIꢗ�d�hwE�mE�g��Мp:�5b�1@m����eس�J8��48�'];9�d��tXn�-j�r�v7��b7fk�q�7F#q�4���\��#��Cm6s�|�0HlJ�2�[\������&>�$+�Î] ����;��[��=<�uٛ����\���!�e�F3�S���%�J�Lhu��Zjy��.c���2B9>�W_�@>�f�����wu�{�Y/�E�cC��q���� w; ��9 �E�ݑLyI�@�z�hwY�r�W�m�@�p/��H�ɓ%&hw; ��9 >W`�� �^�88ر�#rh{���٠}�w4���9{��`�c�1�QƖ7�����ۮ�;<�{k�`�b4'F۲�/6�\�{$�2<$ ӏ@>�f�}n�wu�]��Q.w�$1ƒ�I&���P��w; o�� �]�rVYج�#��19���hwW��$�6}�٠w��h|�^Wqf&���L���}�@��� ;����de�AA�sn= �m������hwW�Z��1Db����ľ�s�BZ��6�N����\��X���*�QӜ,4�&8<��&�}n�wu�]���l�>�!|������3j ws����+��*�.(apq�0�ԓ@��� �m�
 t���A@˟���O;��
\]�c��<# ӏ@>�f��e@�v �.@K�Ʈ�v�����<���'�ՠr���rN��s��=��z������&�)�r
H�X�dL�l&g\YDOM��e�	- ��p�M�3�$X��"���_�@�����z����;�"�R7$�� ~\�>YP�; {����"���i��^����h�Y�U�^��;�YdRa�@|����}�@:�r�uݙ.��1�9��l�*�@�ֽ��� �A^$�Is��~���|�Z<�+)�;wW;�HU�b�8ɞ#��p&6���o�r�^�}n�z�4�|�C#�B8��� �T �]�7�� �]�A�'n
8��w4�hwW�r�@�1.�dX�3$i9P�v �s��� �� z����H�d��)$�*�W�r�@�zj���4	J���`�Ge���k4��Z۷�nxcq���ڂa�v��<jҗ[]�ȭ�z��V�95X�+.��ѣ:�f׃y�@O������+�o'&k� I�糱1I�c��z#3ն���g�q�auڸ66�۶��z���O*�g��J����k�*��GW;ƭ`YE@��6D�9ٸ��ŷ�#�i#s;Uz�n�X{[����WbQ��.nU<�	m�����k����p���@+9�==�']b95�w���:�	��� �$��J��]=Ը,��R#��G#�/��h�l�*�W�r�@�p��8��<jL��٠r�W�r�^�����=�C��)0DĜ�/uz���>y� >W`[��ҷ(�ݼ�܀˰�e@+��Z��� $����2(8ծ6�-6m��՞�N4𽪍m��	a��qGiƜ�@�빠����� �hF%ج �3	�&h��r�RC�IU�ޗ��&h���{���pX�1��h���u��̨�v��/CJ�C+6�����&h����&hr��I9v�z�pY?1�!�c���>�w4�����ܻ 鼫t�1n���}TM��>1�"�yȞ�Њ��$���[x1�$B|N)�cds4�٠U�^�w[4�w4x�P��Aɑ[���h�������N��;ݜh��@)qw��$Px�H�q�u��O�CE�R��T��4��z�%l�A@qF8Ӓh�S@=m�]��u�@�1.�a�@Œ��@+����u��� �����74��Y���uLnlb�ƺݕT[�i1���;3�����<a�u�s`�f�ww`�9 ����R y]�^�e����i��]k�/���z�4
���>��,��p�<�����R y�`}�@:�� �p��q�Q�ǒHh��@��_$��{�䟑0"��R���u��qr?����)�rhw9 ����R y]�wV]�e�_�}ž�a��u��#�m�m�Vm�qcX�qXX0�ֹ@�Im�u���ֲk���o���� �H�v �s����kr��D(7#�/��h�Y�U�@��^��b]��"��d�5&h�L�#����IU%M����;�ڴ	�/;������M���^����h�Y�^�t2Sƛ� ����ʀy�}�@2��*���$I�$ @�$H$@1 I�4(�D��dH@�		1�B�XTp\%9�41�\HX�p �%0!HT�	X�D��	B�Ip�?�
OC�B0���"y>iB�1 %H>FB@� p5*�%1�y�Da$<=̄PX@ A���X�R@��DHH�d@�qR�
@�
x�
��8�d$)�,����Hʑ)$�
bń0L
`̐2�J�F�J����-X��P���$�i1p5�#��a"� � �%aFc�X$a �	$�!~��J�S���s�&��m�5���iܶL�lg�j{6ZYF!|)�����5�m템h�c�2=-ki����Q�K�����}���4d�l�kaRd�����E�6��g8	�w&�R�qx�gXE:3Ű��q��[�l���٧�pm�˔ޤss�J��d�U�!��H�nk�lKH�tc"]�s�j��Z��|��Q�4��1;�ص�[Vnv�US��6ޡ��:�F�;��e���r\픞�SHvL��Jz��3��97$��V.�lg��ee[W>iї�[j3%�q�Q�:ō"+��y�.��rN�c�^23n��.T�V���氵��U�<OB�m�2�a�8�*+R�p�R�����aW��l�f��e�٬m�/V��;0���q�"�U�Z;$�#��nҽ����ʽT��6�ݱ��p�UVm ����Y�nGsc�e������E��Ϩ�%���[��s��5���%rTpp��ٷ.��x�1��K5�٦��Y�a1��e�0��F�Z$���Bݗrmu��h��6H��Mȱ[1kM��ڈ!入;tʤ-Q� ��]Z8˘f[����ey9R�!�wkD��j�U֗f�Cۘ"⛲�񱪽���5�u�M���*�l[�.�G[p,�Qq�m�۳ЯH!�nQ-�rt���i�M�5�����1�e���Ժ�:j��a:^٥�U�b���T�KX�f�e{;�gVRB�f�U�A���L�l���.�:;4��<׳��E��h�UUJ�Ҭ�� ڶ6�|v�v�kg�N�6H x��탎W�;��눛�Z���ZGsT��ό�P赸h�:r�#<�u��Nd$u�޲e<�gn#�y�^Ec��T���~��
\��{qrs�]�m*��P*�U�u��ڤ�7*�^�[���1��`tv1[؇�ㅎxn}�u�Gv�N��ᙻe�͆�t�R����TT|�&C�ff�Y��=7gl\e�:�k����GP�v"iT����g�<!m�v�6a�N�FNY�S���u��֣���um����ɰ6Y�%��ku�]��9�@Mt=�s7#����`5���m�	ʜ@����y;d�V��s�퐕+��a�m�q�ק;$Z�j�"����nZ8��Բ	�ܜ�5�\,��.�WD"�������=�zjt��	�Z`+`�c�\�� ]�Bw[ �v8ȵ�' �u�{�s�q��[?���� �����@:�r��ل��V����/��^�R���N�����/���=�dQ#r,̽?z^�����R���ڴ>�zK���B<O&F�q��k�/���<�W�U�^�u�0�Lq-��3w �T�����u�s���x���9�[�F����krM;�����F�B�^���koO X�q[���y�^�������u�r �fh�<�N�Ħ1�ɠU�^ϘPB1XFD�  0��,0"��H
H 0�J���^�=�@>���T��!�c����)�7�W~���w4׬�*�@�r���ŏ&6��/�� <����u�r�����ˉdL��� ��4
���9zנ_[��w_��,�LxIn)1��9��}$������mb��i!�n�l.�Ż1��@���v �s��.@�P�Y��]�˒F�A�8�^��zj���h�K�IRI��7-rx5��.��w�z{�V�}=3O�*�_UR��Y������z�c~N`��X�㙠�f�Wuz/Z�=��܀_`�;�)�d��ɠr�(���w��h��@�P�M\J+1bJ���W"�qt��#V�=��}�ю�� �AȦH	�90��1���9u�@|����}�@>�6�lҶ�C37 �T � o��_Z��	���P�f�z�4
���9u�@��s@���QF�0O��*�@�ֽ���٘������4�NQg,Ǌ٘Y����\�>YP���� yj�/�w��N��`�`���t�$gJ������s�����뎎��H>�|����}�@;�nɅ�R�ȦD�9��f�z�4
���;��@��s@�A�bw17�51)&��s��[�>YP����[va�'�cMǠ{��@��s@=������v%r<�I��h�T ��`�9 �b�����~��p� 0�LXL%&�I�c'���NFѮy�D���ƫ�͎0�2q'a�O�7]����_��j	���ۡ�,�.F{֤��;U��e8ys��E�\kZYz�3�koEe�ƅ������
v�
�s�l�(½mõ��s;@����9�JG/h���vɋn�*�buE,4�����r�ѫ��������)��2�ڹ����ww���ٺnet#�+���{\�Մ�n���u���-�v�,�`$'92d��RL���M�� ����T�^�f8V�n�e�����{�n��٠\]�QI�H�"���j�,���`�9 9���j��r$�܏@�m��u�@��^��ֽ�Ļ�&A�1&�h�� ��r���� 9��3sxȓ�yu��Wwn��d�k�\�ˮD�G�m�B<)����1�&�Wuz�� +* {�`�E��c[EY{F��f� �.�,��]�7�^����A��LfG���/���u�@��� �[4��R�rd�71&����f�Wuz�hgʤ��ߖ���
��e�vۼ�?z^��U^�����ՠzL�'��?6~ۉ��E�V���8��4���L���h�[��/d�=x�q{7��C?`�b��ʀ��}�@n�.D�c�1Ĝ�@��s@=�f�Wuz�v��Ļ��"M�#s4���?z^���%M�^G�O�ՠ}�yخF)�	�#�*�@�;V�}n���^�{�Yw& ���f���n �e@>�\�7��ۗb$I����n)��	6�{gVwc٭�v��a�<�g���rζ�L]^n��ʀ}|� o�����*�&1��5$�˭z]���j�/���=��4��) ,��}�@=ط |���\������x��X�y���*UO�;����ՠ|�%��JRH�/@=Uar%�ő�$�Z����Z�
���=�ՠ�a`D��`��$�Zegln���������֢��2m�=���<N|H1���f���^�Wuz�v�������`҃�$n%�����}ط |���� v"n� #$r=�;V�z��:�I7�'^��w^���!�v��V^�y�p�T��r �.@>����*�&1��5$���^�_���_��'�ՠZ[J�R��Ov���tF�"k�9�8���V��-���F��!V�[�;W#���j������o�����v��o<E�������N�ݨ���p�N�[��=uz�R�h��΃\κ�Yf�����2ڥ9��m��:�� ���2����!Z|�Y�cR��N�5�1��
�/�ݲ���7i�ikb8Z.R
䞎EZ�xڼ������
X{�$�g�[��_}��Ǝ��.�{kkv���:�lr�l�6.�g�:8L��6�N>�~��s���hWZ��|j��c�	�R=݋p�T�ː�r swm�r%�#Iȴ��h]k��%�[��_��@�1.�a��rD&�hu'듯@�'^���#��{���>������	���Wuz��������ՠ|��z��UT��F^7��S�!r`��6��a^������M9̠���ݎ��۷M"��6������	$ՠ|���~aϻ�@�"�2��o,Ww�@��V��U]TYN�����G�I�H9�w����o3��'^���?�������������=��d�&H�CR=����r=zMZ�ru���|���m���Ÿ�*��r �5�=��"A$X8����QAƨ����=��Vn�p�5��kh�<	~�F��u�z�����ݫ@�z^��/�RK������@����?�<Yj��n����@�r �� |���U]�C+�/�
H��@����zSE��T���F	T�
'��,`���H����$@ "�0�!�a @����"Ȥ~X�
@`��aH�����E��@�C�`��D�:!��Q?��	����@?�Z<E3򊮭���ՠ|��z���[�� �2���/C�>��4�v�9�z~��q�(:ڃı9�'����ϧ_�'_s�$�C@=��9�"��!U�/���m�g�7�E��t]��$���m�����3�n��e�1[���}�z���	&C���W�����@��'��fb̑�6�N=��h�M���rK�UI6
.�o��y��o���ݜ{�$էRo�w^�:����*�d��B�����Vנuv�-���bW�E2<qē{P��8� WR�ʀz���W5��\�v{Vۨ�9D7VЇg��]��G���n��י���]�q՚r�-�Ԁr�����D'q��HܒE�[e4�w4
��@��������<I�bi� ^e@W ��]H�u&�'��"rf�U��_U�[e4z�h�b�#�Ƥ� '/@����Iwv����ZrK�-�_E{Od��d��2ܚ�q��'��=�֎5�n�sA�L���ی�K����q����[��X3�m�c���/l�`�v۷-�6�i�'8(�$�-���ۜ�u��V�S�!��YBc�A�
�ݪӥ��<����kv����ul���;h�kd�޸Y��q%�ͻ�v����6�6(ƚ�tP@M=����k�����ZT�\�:ø�c�4R�'kNק�}ן�W,���ʆٻ-�[n!�I�f��7b�;۷=>Kj)��6�������-�s@���]�@��1O�1I�@����k�-v��k�=���2)�L$�fm@W �p�������8�y#QF��-v��k�:۹�Umz��dƝɆ(��swn ڹ �e@W ���������@V���ex���q(6�P.;��l;���q�{e,�2ݗ�� U� m\�.-�W �
��r#�L�I�V׫;�f|T��*T��X__s�9�u��nh�b�s�$�$��:�V�m\�r��������ѷ��{�����Uڠm��9w(��- ���YrS�)$��m��*W ���r�]V�ں�skC*@�3>�zQ�{U������h��e{:�Ęcd��!�)��N$���k�9Ÿj��e@>��j�6�3ks37 �7 m\�r����݂���<>)#rI�U��lբ�IUSq�/@��G�~��<.]��.�ͬ�����j�qnU����SRn��I3@�ېŸj�VT��`iy[j�g�������̉����4Lr�0�� j��@�����71%#�-v��[�*ʀ7ː�{�9F�晸m�� {�
�����ՠT\YrS�)�h۹ o�����-�=�m^5[x��w�����IS�נw_s�'�G��UI~J���'�}���c�^�n^n@�:�YP���m�~�L�v%f,H��r��ԯ����<Xb��pJPջ�Hg��+w]�n�m�:�YP���.-�=�`�`�F�71�Š[n�Wuz�ՠ_;V��\56�>9�%�� o�����-�e@/��I��Ĉ�z�ՠ^v����]��\�����LS/36��n �ʀ7���[�M�T�sB�`�V�n���̻�:tv�ƫ�k�I��3�Xm)��D$%���v���shۣ��z��]`v��I��V�ǭ��=�u�j��1�Q����-�m��8�E䬹mQt֌I�H���nrZ�
x6�Hhp�\�q���٘�r�N��a.6�rR�!E�,�тCh%�m:��g���4=ͻ`M.]��vn�	�f�#t�r˺���3e��G�u�\��F6����n#m\��/^�n	��:�8�HQQ��~���Ҡ�9 {��n�0�k>I�n	��]k�/;V�yڴ��h|.+	X�Q7�y��Ÿ�* �.@=�E��c��N7�yڴ��hwW�^v��v
4�hBs�Z�%����#�?�*O��]vzi�B7���N:{mvx ��O����-�ǷfK�nàZ7W]vj��ֿ� {��n �* �j������e�\�u-UUT�]�b��YP�r SO~�(�k4ڽ����ط ������\�b�ڑI��s@���˭z�hF%q�c$q��s4
���9wW�_;V��۹���18�1��&�&Li�H+��ۖ�[<��A�g�uW>�����<�k�T;v�ͼ��_s�ط �YP���wv&7aFL��8��j�>VT�\�u���:�ѭ�ݲ�nd$�@��s@��ק��Ĺ;^�yڴ�`��7	��0�L�..��?Iz���9URI���-�rj~Bq0hp�E#�9u�@��Z�]���^���
�����i%��4�>8�Xnb�nO�ϖy�]bvפq˳ׇ�7��D8LSN=�h�w4��z/Z���ŗ �2�"�-�2�_.@:�� {��]�X|�x��Nf�qu�@��^�yڴ^���ʋ"`ڎ(�&��<���	��OMZ�j%J��SX�נ}�`�cv0D���@��p<ʀ5|� ���T��鱎���*Vܱt����;tuat�F���D�Fd� ��dȜ���2
E�z�* ����ː�n��z�]�[W��^b�"~���6G���:_��@�빠}�qd�N&���R=�ː�n�P�� 4�`�&5�'�yڴ^���ֽ��z�r�ːby>FF���P�� ~\�=�p��?H~��$ "D�HE�0��	�$b@������d$�5k��A�� �B$P�+Њp��$��B�C�O9"�"�0%��2FBbF0�e�)RH� ���i$ T!d!#(��21 �H� H��B ��D����H,��I	!"D�)�P<? ��X���*�$R)H������21H��=�;���Ѧgz���wM��	�qȜ��նwn�v���T�Л���w�j�9��=:��T��A��̉eѥ-��ե6���ܡ���:��gd��}Gdc��Mڎ��n��5\B��4[�!٠yݛY���\���,��J칕���1�������������i�Kn��:j$�֛������pv���v�UXړ���{c[����y�"������ƷV�=a��$qfB�x^�UT�n{d5*ʷRE�s��N���PSi���cUp!b(a�G-'3Jh1\ ���q�@�9�����`�y���8�
�mŮ��<ۜ9��SR�`R��L��wOdCdn;����I��W'���iH��X:o�siѣ�����M�*�ܯU-�vf�t9��Vj��b\(�m�j���DU�L�fVu:��^]�/E��j} �m�ΎŃ�@N�e��l*�K3�#e�e�l�n�p�
�qٚ��wN��<`��4,�/6Ժ�˧��f�r��#ny-���8��cP:�n2��ي6�9B^k!�u�]ʹ8�����,y" rLn����!�`1Z	�,y��Q��m�aۻJ�v���Cœ��W�0�7:+9�mEam���r0�J�̼=�E۲gf;b{a&���g�Y�͊��K���r,�.�@�ī�)c�|;r��=tr�eY�����$,6δi4��P��om�kMPT���ll;8M��g�GuT�UTt�*� �ݶ٦�ЖuJ��m�w@���e3�a�uDp�j�U��ZA��V��ە[�m�9ۧ��ۛ���e$��t���z�$$`׬��흷�z�ϗ]H���Ri. ��X�)+��om�m��x�怹�˅�`�mU�"E���������ۇ �p�x���ln4���RstfN7n��&鹻��4 zP���� 
�����3HC�M����l�yyk��Q(�.�Ө�lᣌ\������٤�8�=��vwkRm9�BH"+G7�.�R�;L=�6�GI�New)fi�vy� ��-S;H��WH:8�uEϞ�r��X{�f��鍌��֛'T��^;�ѝ�Y�,�c�f]�6�p��L��ʬ����OU�4�ny�R��:x8w:G�;d�S�����훴�#X���	���ܸq�� �(W.���L�:��g�ޞg�84�p��z/uz�j�>޻��ʋ"`�����@��@{�<ʀ5|� �u[Y��iE������@��s@��נr�^����B���a�̄�h�w4��z/Z��ՠwp)P�r,r)�#�4��z/Z��ՠ}=5h�U*I��Ӵ�#�am��ź[�����c�v�n-ۻm@Ul�f�-�;n+v9Œ!8��q�R?�_��^v��]���^�ge����df4���[�U��ج� j�r ߗ'�6�rk�X�2��y�@�ݫ@�wW�Uֽ�ڴ���A�'N4����@����ڴ�ˊȠbp�����
�k�b��e@�\�u�ѻ��s�n�t��0�ه�����յeq�q�,{u;-φ)�ɉ�k)���yڴ�� j�r ߗ q�^�f������� j���7ː�j�=܅*�KG&huz���=J��I
��Ud��z����Q5��xZ2�[�7�zT��'.w^�޾�}$ՠD��z ������<KN=�ڴ[w4����Z��G���`�'&&AG�T�r�76����2!�N�]�t'X쥍�x�L'�ܑ���h��]k�*�^��ZJ��Bq��ۙ�5o9 ���o9 �pe6YN�1��˭zW���ϟ������h��w���CX��x"�X�e��K�'�ՠD��bWJ���DP|x���_�o�g$�}>%��[���ȣ�@�n�q^�@��zs���T��j;O��]��cM⻻��V[N�/l��k�m�q��㳟my݃���{�1��m�c�" ��������*�^�U����hnv,���ơ�Iz~�����W�%v?�������h9��v^���AA�i8�
�W�OI�N�M�}:�s���g�����F8ے=����z����r�}}:���}e�<c��w�wx��� �����<�������g�O>.c*�֔.�nף��:)9Ã��4�l�g/;��p����`�ѭ�B�mƓ�E�����d�v�&�utۨyq��B�ƨ��S�*zP
ϗJ�ڵ�pMآ	��8�6��T���75ǎy3�����	T��E�:;h�џk��B��')��܋9Sa���ԂX䆶��p�J\�fNjpu۝��Vz_^:�~��|�c���ܽ��֨\�q�D�Nl^�mݝ��L�Ѣޗf�듐��I�519����zW��/�����J���O���@��CX���V���-�^������M���Z'ӯ@�ޗ�K�*��q�x[xbfb����?����q^�O|��]T���|�n�V�����ʒN+���y���*�^��۹�_a���XG1�bS/@�����*������V����Uȷ�?Û�&��Db AF�V6���aϩ�&`�qщN��{�n:|���c����>�z�&�'=/�T�/�R_Xs��� ���Maww�ۼ��̽��Vڤ�dNz^������K�I$�"撬����m����/���<���*�^�����>�<���O��&�;̽��T�ru��u��&�':���,�Ӹ���)�)�U���T�ӻ��'ӯ@������g��B7@ݎц�S�ۇ������ݻk�P�!��.�g��5�ܝ]3?m�I5h9�z��/���0�ӯ@�D/�f��"1�3@��W�r�@�z^��I��*K��+��!g����/x�y��s���9�zS��:����h�N� QOU�E��o�o2�?�I����>�ڴ���?�/@8��X672$�NG�}�w4�Ir���G�נG$��bj�k��I'�㦎q�OD#ա中@��<ܶu��/)����Y��~q��/@������%���;V��\�f5���e�Ww��y��{��*M�����v�'$��T��*Uvt�5���m6�Ȕ�@�_���@�z�h�����x�D&2L�8�?|��?���h�w^�����=J��J��RR���IV��/@��!m�^1e��b�"rK�9$���u��w^��z�ho\f���)$nLr@��6җfD���T�6g������-��c�3�G0qbN=����k�>޻���|���'�נ�u_Z-e�1�����#�^���5h9%�?�/�K�$��a��G� ��m�BLI����ۚ�mz����k�;+Is.@Y�wx]�-�UI>W�נG'^���?�J����h@���c�v̳+���<��z*K�UUW�_�{���V��^���U@��Z�]�;�wy�e��ɌZk������mU�9���68����p�^�c�v�i6k@��7Eڝ�j��C�uűk	v��ݳ� �	Mڹ��:�lE��w��rͣ����	ӷz�D[�}�	�vLx�nCv��`�XǶ�7lhd�ˮ�j�X0sׂ���Ȉ�mۋi��$f͸v��,�Mp����ktX�l�'m� ��e�7bV���Y;uf�V�9�u�O^���&f��۰W�y.�:���c��FU�
�o������MZNI�T���9:���#5�dqǠ}��h����zrK�UT�=��<��X�3���u�~��9%������%b��9��q����*�^�>�V�U'����Eү���zYw����� j��}���gQ���XЛ��E�9�o<�;�m[�i��9D�K�&�[]z�c���ɾ��Xz�<kr?�{��ۚ�mz.��
��@�%̸E8�pnC@���r������P�>C�u�����M[��M�@���bɍ������V�zWj�>�w4
��h݂ɂw�I$��)��Iz�2qɚ�$��נ}т���Ƀ"n8������4]��[^�w�֠�R���Q`��<3z�|�{m�O;S�+����=]�)�9	���q�@����uzVנ}�S@��%q��9���h~���I��w^��vq�FI&�e��y&<x��ґ�[^�����OWı�8@1�.�Ȅ��+(��pJ�AT4�
��XAU"DE�H"A� �H@"�CDx54T@<_S��$]D_^!�l���9u�@8�����8����Τ�]�7���r��öƱ;ye�w�h�L�9*J����}�z�2�T��/-�8\%ڥ-���g����-�莝�[Ll�B��&ǊH�Lx���ܚ.��
��˩ lW`�E���n]��ї����˩ lW`}��>� PV5 BpL�=�v��]�u�9 m\�w�-��m��ѵ�V^���_s������b(/�w���'����.�Ƞ	ɠr�@����j�+'�hJ�%�4>�S��cǘ�+�9�{h`n�-����0�P*�ڸ�Pz�<sy�H��CJG������ڴ
��h���*;����x���8� ly�_s��r��wȸE���prE�T^�@�ֽ������>�<���'ŏ$	$��UI9~��N��~�@����w��qdK�)�k�ٕ^�ߗ�9���^�)u�Dp��6�l�X,�GSgn��sF\t�]e�X;\���+�U�e�p[�\���){;\�õ���۬c1ǘ:��V�[�]��<�l&]�3���T��U��om��G`���g�a�y�ΉX��n�Q��ݻ����n�&�1�����r��J��49E���Pj�n*aF�J-\����!gGI'���:qzE�	ԄWc5��]��Ӻ�0����;G.v;P��{U�����6,R[cD�}���4
��4
�k�9^�@��W����G����\�u���R �:�ݬ�o`���]k�9^�@�e4
��4;/|u䍤�N=����Hm�����߮���p�'�9�}e4
��4
���9^�@/��"NdƤ"��&F(dńI�I$r����4�"̧K!s#d4q`Mv�LdD�9������W�����g�-r}��;i��f[��?}�s���Q�@���s�N���rIU]f�{�Y1\�F�"@IǠr��� ly�}�@=�az[���ȡ$z���*/Y�U�^�U����fȤHdp�*o��7���� �T �vU�[�B�B*[������q@A�������z���ܓ��Y���L��+#�*�m�m� ��@,�c��
�{�9�6�phiH�
�W�_[��T^�@��� ⣱��QĔĜ�@|����>�߿U�}�@W U�r.dc"i��E�hw[�#�^��R���ߖ��\�f5�E��fy�~�������{�V�UV����)����$�uL�ڻm�`��#����;��sv��n�ekq���И�dɑH�Vנ_u��*�٠U�@�y�����z���8��?�/@�^�UR�����1�6��/1h��f�ޗ�r�����|�J�Ǒ)�'y�z^��$�}�C�YUU*�-�T���&h��2��we��p�r ��P�]�7�r��������1Ü���Gh�=vіeh
���v��#2��b.����L�n`^�r4�6;ӵh�&h��|�U/�#���&~bW�Q"c�d�'3@��f�W������w7�|H�,�X�4<LM�*�W�r�P����9Ul�/��+�$F<S&E#�9[^�}�s@��f�W����
*���R���; m��~� j�� ���HN���f�̳6G3\����`5��*뭸��<YŌ�:�z�:�U�h7$��w^2b�Y��Y���p�r�H��N�=�ո�j�:L[�3�8;lӐ\�t��y�!N�-�N��Y-�@X�,%�z�x9����<Ǜ\:q'J:G$Q���.�!cc ns�^g^����+�G���@U���ѱ�t�,�E�{ǉ^v%��z�-*V�M��c���=��#1��v.��Gݗ'<]��և��	#@��ӓ�UV��uz+k��@��%���w����@:�� ���6�� ��~5BD4�I��z+k��N�T�&�������@!)�(���]�e��7�vh��f�ޗ�r����.EȑX�I#rh6� o���\������v�y�5�kGF뵚�J1���k���۲�%��*��N.�~������1uɞn	��s���<䗠�L�#�LөR�A�A�A�ޒ�>ɳf�]ɥ���� � � � �>�����F"�t��A �`�~��o �`�`�`��}~�x �����|�����d��f�i	0�ݙ��|��������|�����������lA��9��w�����lll~�������lll{ޒ�C͛�ۛ-������ll_� �d���o �`�`�`�����8 ���}�|��������|��������n��fl��ۛ�|������~�>A����*�����A����w��x ������� � � � �'^�2��7xCy���q�/:ݴJ�ݽ�'f�Ǯ�����6i*Ö:���ۛ�웥ɛ��[��?��`�`�`��g �`�`�`�~�ﷂ�A�A�A�A�>�}�|��������|�����}g����&��L���|�����߾�>A�A�A�A�>�}�|��������|����s��>A�����-�n�e͓w77w��A�A�A�A�'�}�|��������|��>*��C���,���`Eb�0�(�����A�>g���pA�6667����>A����dߤ���.d�����>A�����~�>A�����ﳂ�A�A�A�A�{���� � � � ����>A��������m6i�ܚ[��|�������g �`�`�b��#?����A����'����A�666?g{�pA�666?g�^���n�i����klqd��\��Kv1�1���O*:\ml <[u�a��f�4�ݗw8 ���}�|�����>�����lll~����*y���>A�����/�<ٳv\ٙ������lll~���o �`�`�`��w�g �`�`�`��}���� � � � ߽�����?�A �`�����v��77-�&n� �`�`�`���}��|������~�>A�Q�A�A�{���� � � � ����>A����>��d˛��[��|�������g �`�`�`�~�ﷂ�A�A��>��䞂����~�;��gU��`�X��e��L�"-�@����k�=�쎩��A]R�.:h���F��]��oD����3������%�	DL�F�rM��4��z��|�%��������2d�A�4
���=]�@/����3yR�l��'}Xb���M�d�������_Z��� =`�[��y$q8��٠r�l�#���u%I?L�z����x�^��:��`�9 �b� |��'=Ut���@���J1�����
�u|�x��b�@a��X��HH�	�H	�'�@��B1��y<�����n��m��87fݜڣ�wN�F8�Lyr�enx�[crez�FlN4�\��3۰t;�睸.j�%$��qJ��ܚӴ�G)ڹ���V�4R�ƞŵ^:�*��'*�$��p��`:�܎���e�N�J�f[�[Q,����6�:�����*�+>^Z���e��h	�:[��R�aC7�jT���ƹ�l	�V��]���UQ�A��w��6���һ�l�R�W:.Xt�v9��sgv(�NF_kt�������)-��Y6A����H)�3
�4e��Q��.'ذtem4���CN�P
���˘�gD�v�YԲ�l�ӷ�%k <��Sl�e�`����sg#�l���[)T��[� gv�痩V����VU��kZS�	�a�]��l�#�.�r�M��,�v�vf�oe�` 2fyYeu�y��%���h�i�Y����]W8�������hG�.8��!��<�iJ�5U\Q]��Ѵ��ݨ6�Iq���ɀ#�v�g�v9b�͞rpev������V��X@Z�px8Q��fn%]�Ѯan�Kr���%s�E�wc����y`h��N�r`���n:��F�7�
����++u6f���/lb�FNZ!�r�+�cqrQ��۫V��W�;D��U�#�R�q)fH^h,�t;uIŘ���3�b�&�\gTcvRZ�P��^e^Q�T���Gkh�t�n�S�^�����e�Ʀ�����]P�<�s5;:��؍'l�����GW	  ��m�[A��-$�
�j�8�GM��ۨvY�gU�]�nr�S`�Ҳ�T�NSj���e�I��S'��8�9����m��lH-�`��2��<�ϰ-�P�SJ���j�Z��ܬ.Φ3� ���zl��ö�୶��Hf{u&%��9�IX�ã[�p��j�h�u�Vt�ݛ��qtgh�5l&�컴��g�)�(8�DW��� p'}P^����ٷ�w<��k�]�gks�]�-q����y��k0����y�;`�H.]���}���c,��as�����p2q�ڪ3���0�ki�v:�]�F�Ni�S���-�[\��Wm{���M�{b!�Si���>9䵍��t�݌&!�kQv���ً-)�kz�52��%�$0#@L@�Q�<E��kt�(tl��S�'���Z-��pKQ�T4e��X:1t��rDnf�95d�2K���Y�4=��<`�����Umz�ڴ��u*��0�>��u�3n�ۻjG�{��@/���.�@��^����6�]�V�ʻ�f^c����9r�4
���yڴ�Ĺ�e��f��R���;4~�z�\�C�R����٠}��1bŌ/-���� o9 s���`����؅��Xe��"�:s�V;U��WAC<cN����V�?{�����u�QֺDdĜ@�������*�������������P���BA8����t����B#
"A�X� �ȤV!"(Ҥ�-I#q�٠G���s����*T�$C�-�1�3x���>s�@o��[�@˰�CEM���M(�D��*�@�z� ��h~�T�}|�f�(�Q�e���o2�9�z>�4���?z^��J�����߼�m��&�\�n3�z�禱v:
��ðb	��$�f�]e�P^l�q�8L�\���#�����Uu�]���W�u��a�J#&8�hU�h���9�z>���Rl��_,̘�!#RM�����W��f�U]f�{�dM\�"x�N=��� �zf�rf�*�O�ӯ@��� ��IǠ�f�Qm�^��
��@-�)2"8��F�rЗ38�\��8%�pr�b��9y4��c����R.���x"���g�9�ݚ�s��� ���w�!��X���� o���r >�`�3z�M����/.�,�^�/@��נ�L��R�M�;�4~�z��Syph��1��z}�h٠U���b��R�U�;���-�>�ZL����m�PU�@���@/�� ��lܓ#Ĝ�lP�7)�\v�	�˳��G]��v͘cg�:�XM���];����rh{��*�� ��4�f�{�dN�0�&�N=�k�	���I�~����T�g�0xs��1�^aw�����	$�:�Ro��z>��x��ř�y��ʪ��&���@�'^���}$�;���$ɂD�	$�*�@�_w_��vh�f��J�-UBIR_�?����aff �MbgY�Ǳ���n�n#��KD��k.A�#P�5Φ�d;e�$勬b�rv�{su��3�8�ʉ���rz&���k��ݳ�A&����f����7�����9��)�,�9<��ܔ�Ń��u�-��mc>�:;�k����NpsgM\�Z]�cj[��6;I�Ü.m��$�]C�����偭�E�[��������y#�lu�c��6�v;�lf�]B �N�E櫵�qS%���e��q����l]�����r >]�
� o����Ve��)��m9�_[4�f�WuzVנu��a�� H�h�����6�@˰�1kv)��Q�&�WuzVנ�� �٠^�F���!4��*�^��J��wg����#�����~xh��j9�Q��ז��3O1[�랸��<"�� �^��&�TY7(�7����� /; o��o9 �p[C�2'�8�rh�f�33s*�^�W�� ��h��I$��X�A�� o��j� |� 9]��{�L�)1)�����٠m�]��*/���8�mf�@�� �v �s��r {���v�������C��`�.۩V8���z7AX�vZ��!rm�x��c�ڭ�܀���r�-�������Xۼ����#���R�T�:�����נ�f�=�5�r���1ۼ���zIzj�K�J�Ņ����9z�z��JNG��D�P�� 9]�7���[�w�.��E�8$��������ՠU�^�w�	��&�D�G0��~���d�)�ہ�;n���IR�v��+zE�ޗ��ɓ� E$��o�uv��Z���@3��µ1��)��ڶ�A�\ �l�{�����1 �E��V!Dd�i���~�4��@�������yج����q��UI��٠s��@�^�UIJTD�������I?vL�grnܥ�m���� o��j� |� 9[�������n+%�wP�.\�u�ڊ��	���!�M��00��gj�qv:Ϸi�	��*������ �l�*�^�������� �zz٠I�~��䗿�I�H��pX[ME�z����@��zVנUֽ�p�lNL�$Ʉ�hu�@�Iz~��9$�wvh��s�-F�� ��@���
�נm�~���J���'��x[y�O0lƢ��s�vU�\Du�N$�s��y�0�Kn�㤍q�����h�9Y��Y㝜M�B��Y�֮���:,/`��a����|9�l ����m�l�q���/6Wqo��q1��S �e�:|�������Q9�e�RI�v��[v�Z�S�9�&�Y�mv㧻%O���x��2�I	%ٺd�&Wm�7Q�UD����M�8b��ٵ��Y�n�;,t��v�إ�u���$��ƌ�z{����^��w^�zI�~������u�=p�>�X�yE�e�^�zI�}k�*�����h<��D�$�/^f���9%��$�W�IU�����@?�����{�Y��1FF(�zj��[�
� o� =au�w�1�^'���O\�@�K�R������x������� �g!�Lq<���7b��&7 :4I�ݟO�8ݶC�X3��<!��� I�[l�*�\ U�ط |��6�v��[Y[sw�N�{���@Db���m�wvh��I3�US`��]v��X�,n����4	���IRM��٠s�נ6�]�xݻ��y�����}3��wvh�K��I��I��$̥�&Re&R�Naan�swn��'�,Kĳ���r%�bX��{��yı,K;�wS�,K����'�,K���電fn�:��c��hY�n&6^PK��K[9bև�<
�څ77!����~�Bl�i����bX�'�߾�'�,K�����Ȗ%�bw��oȖ%�bY�{���bX�'}���Ι$�ܛ����'�,K�����Ȗ%�bw��oȖ%�bY�{���bX�'s��8�D�A2�D�=��S~��f��.i7w59ı,O��}x�D�,K�����K�c"�z��S��!%�BIJP"B�)
�²�HJJʅfD=�'���$R��j�P��@6� $S&�!��` hLAEQH�rI���5P8��p(IRx�<a�q��@��pD !��GP8 �ED����3<���yı,�{���bX�'��%�3��n�l�l��x�D�,K�}��r%�bX��{��yı,��ND�,�J�)t�紿�I���N,w�(�4�nn�r%�bX��{��yı,���"X�%��w��O"X�%�g�{���bX�'����e!�n���E[��;m�^K�nx����u���V�*X���;Xa��a����t�nnx��X�%�{߳S�,K����'�,Kĳ�{���<��,K���gȖ!���~������.��M��{��ı;�����Kı,��wS�,K��{�s��Kİo��jr%�bX��I���̄�6�7n��'�,Kĳ��u9ı,N��8�D��a�2��f�"X�%����׉�Kı?I0�:]��Zf�vnn�r%�bX��}�q<�bX����"X�%�����'�,K�������)iI��I���CZ,w�f���yı,��ND�,K�#������ı,K=����K��J_�/i~)2�)2����d�ym��@�k��l�{ �= �8k��Y];�,�`�c��!���oq��%�����'�,Kĳ�{���bX�'s�{�O"X�%�}���Ȗ%�b{��/I�͆��ɦI����Kı,���!�����]��,O�����yı,K>��u9ı,T�������L��^�,w�(�Ya�7u9ı,N��8�D�,K�}��r%�bX����q<�bX�%�����Kı)��^���7ffKws��Kτ��2w�n�"X�%��{����%�bX�~�wS�,K��{�s��Kı,�/\�wi�2i�n��"X�%�����Ȗ%�bY���ND�,K���'�,Kĳ�{���bX�%v�2~���1���Ф���A	�R�M\4�gw8ƛ�Kvh9K��`�x�'�9n���p��{kHz����;{u81��g�a4��ɼr�q��]�WV[ M.4F�!�,�i8��:�띴� ����a�m�&�{x66�viU32�i�k�� F����۷��"D��~ �����$%��7	�����\qFb�q�c�[��3eɷ�D=�.�4�w7d�U�/b;�Og�(�W2�]z�f�k�#vT9ۀ��\V璶�SO�����{��"Y��S�,K��{�s��Kı,��wC��L�bX�g�}�O"�oq�߻g�?�Ҁ3��W���,K���'�,Kĳ���ND�,K����'�,Kĳ���ND�,K��Js3�Bl3vnM����%�bX�~���Ȗ%�bw?w���%����,��n�"X�%��w�gȖ%�`�����\&���&f�"X�%�����'�,Kĳ���ND�,K���'�,Kĳ�{���bX�'������d6�nBf��yı,K?w��Ȗ%�a� G��~�'�%�bY�����bX�'o{x�D�,K�N�r�nn��fjqjT6�i$v<-���\�mL��u��l.p���E�^ﷸ��{���}����%�bX�{�wS�,K����oȖ%�bY���ND�,K����a��]ɹ2[��O"X�%�g���r"���ȥv&ı>����yı,K;�۩Ȗ%�bw=����%�bX�N��w�̹&��wwu9ı,N����<�bX�%����Ȗ?�C"dO���8�D�,K��̥�&Re&R��&	���2���yĳ�D��2}�۩Ȗ%�b}�����%�bX�w��ND�,K����O"X�%��I�s���,��w73wu9ı,N��8�D�,K����Ȗ%�bw�����Kı,�{���bX�'��w:iw3z��,e�l\��[/uƞ���ҁj��8X��mn�Rx��w� :_��ƌݡ�����%�bY��n�"X�%�����'�,Kĳ���r%�bX��}�q<�bX��IM���6]�\�77u9ı,N���8�D�,K����Ȗ%�bw=����%�bX�w��ND�\��,N��)���eۻ2�ws��Kı,��S�,K��{�s��K@WU(�A��ؖw��ND�,K����'�,K����fK�5���m��ND�,K���'�,Kĳ���r%�bX����8�D�,K����Ȗ%�bSӽ{��ɻ�s%����%�bX�w��ND�,K�#��߳��%�bX�}�۩Ȗ%�bw?{��yı,K���6�L i�v�qǜ<�W�k4ch2�Њ���:�؜qy,�*���9ı,N��{�O"X�%�g{���Kı;���q<�bX�%��wS�,K���M=/w)7srL�����yı,K;��!��"dK���gȖ%�bY��n�"X�%����s��Kı?I3�:f�S3n����ND�,K����Ȗ%�bY��u9ı,N��{�O"X�%�I&e-)2�)2�������xs78�D�,�QC�(lM���۩Ȗ%�bg����Kı,�{���bX�� �t
 �bf�{�O"X�%���S{�L�nf����bX�'s��8�D�,K����n��,K��;߳��Kı=3)iI��I�������<y��ԣt�	rv��;V�'0V��^���I�؁x��ɮ����\��7'%?{���oq���g}��r%�bX��}�q<�bX�%����Ȗ%�bw?w���%�bX=�m�%��f�swS�,K��{�s��Kı,��ND�,K����'�,Kĳ��u9ı,Jzw׹�᥺]2[��O"X�%�g}��r%�bX����q<�c����,��n�"X�%��wﳉ�K�7���ߞ.g�K��w��o�w92's{��yı,K;�wS�,K��{�s��Kı,��ND�,K��4���ۻ�nn���'�,Kĳ��u9ı,N��8�D�,K�����Kı;�{���%�bX��!���l7wrI��-������W7\�T��6�8�;��.�v���]q=���;�cN �W[͍�nc�#�g7Vî�.��݁L�MY�D+q�V���ة�(K���XvŎxp�Sm�@�Rۄ-Z�b�s��[���;+�.�̅4�����:����/P��v\�vI�l��q6�Ŵg�e'�rv��J�yw��j�;�����{���$���乡�n��$�O^���R�G.
)7rŨ�Nn��&����Kı>����yı,K;�wS�,K����oȖ%�bRzfRғ)2�)O�mǍe���s78�D�,K�����Kı;�{���%�bX�w��"X�%�����Ȗ%�`�����\�M�&nۻ��Ȗ%�bw�����Kı,��ND�,K���'�,Kĳ��u9ı,O{%:\�a���2�7oȖ%�bY�{���bX�'s�{�O"X�%�g}��r%�`�"w���/�&Re&*���c�2�Ŋ�<���Kı;����yı,K;�wS�,K����oȖ%�bY�L�ZRe&Re)�48�,w�m��A�jGc�7a���<��͑��[����y��v��v훓e����%�bX�w��"X�%�����'�,Kĳ��t>�DȖ%��w�gȖ%�bY>��0�6��]3-����Kı;�{���QB�"X=����Kı;���q<�bX�%����Ȗ#)2���ɍ�2��32�1�/�&QbX=����Kı;����y��dL�g��u9ı,O�߾�O"X�Re/2��B��yyt���N%�����Ȗ%�bY��u9ı,N���8�D�,K���'"X�%����Nͦ-�4����yı,K;�wS�,K��~�s��Kı;=�19ı,N��8�D�,x������1l�=rEuk\u�\���n�� .曘�GJ�6yK���U����f�����Kı;�{���%�bX���19ı,N��8!�@�It�T�R���w�,wj�Ɲ��	 �'��jlNı,N��8�D�,K�����Kı;�{���)��I����Ǹbŋ�˥�&%�bw=����%�bX�w��"X��0��!Ȝ��O"X�%�{}��r%�bX���nM͆�[��ws��Kı,��ND�,K����O"X�%�{}��r%�`��"}�����%�bX�O��ϴ���˦e�����bX�'o{x�D�,K�����Kı;����yı,�{���bX�%�����N��Z6����� 'Rչ�3����6����\�l�v�3�RM@���%�bX����'"X�%�����Ȗ%�`�����Kı;�{״��I��K�\-�XZ0��e�3q9ı,N��8�D�,K���"X�%�����'�,KĽ��q9�2�D�>��S�fܛ[��377s��Kİo��59ı,N����yı,K��w�,K��{��Ȗ%�`������ɴ�4�n��"X�@ȟw�}x�D�,K�~�q9ı,N��q<�bX���
v�߳S�,K�󽒟�6�t�����%�bX����'"X�%�����'�,K�����Ȗ%�bw��oȖ%�bY�=�?��-d5T�LQ4s���:���Gq��l�b�Q��i��)6��]��w��bX�'s��8�D�,K���"X�%�����'�,KĽ��q9ı,Jzw״��s.fi����yı,�{���bX�'s��8�D�,K�����Kı;�����%�bX4�{�f�M�2\��ND�,K��{�O"X�%�{}��r%�bX��{��yı,�{���bX�'��i��v��������yı,K��w�,K��{��Ȗ%�`�����Kı;�����K�L�������o0w�t���N%�����'�,K���sS�,K����'�,KĽ��q9ı,J��z���@a�$������͡(�� , ��1��,��dB+��HR! ������ D�0c<ex`�B
NJ��@/�k1m�#ļ )|E����N��$$c$"�H�,Y�᠐��ȑ#n��)���Ԡ�X(@��@X�P�B D�Ă1��!1��A�$"Ċ����+���`ł"�H�"��9$�F)`�`�0��! 0q#$ A�U�DF!��T�ՉȲ"A"D!%@�@)i�D��	!H��O�N��������:�6#�d��Xm��
t�sQ#r�=����f�o���}
���n�㞙�nټ8���l�v2�V꘣�<
H=msn)V�w<-s�m��z��&�ir��Jܬ7��1����yˇ��쩺s�U1�ͣ�9akD��ۛH�%=U�N�;6@��܎�{r��*c]09�ӗ`&��qmg��n�����[Pnvu��y�=���z&*��u�)v� ��:��lv�d9ѻ[:�Q��}E�O�p;W�=X]�Ү�B�j �'+*˄{��v	�����'m��Vg��h�9T%V�N۲K];�}��=��������e�qv�{ܕ3�X*0�3������+W�˴�[|�����#5����p������jRn�TH���f��n��8�O������-�,qmO6F���$�Þ.r +!0bU���a�tp	�4��lt��.ª�p#�A��2U��.2�*��e��̻\�U��iι�5[��N�j���\jlNݢL�Ѧ4�U8�P6�]<��ķ=g�`�6$�4Aۡv��c{�a��Β�ò�h1V&D��Y��G(�j6���݋��k�����,�x�&ێ�`g���nPR,a{'P�1�E��!�̡�h.����RX�]������l9ְs�g.�*�W���s������u4� 4ԙ�J�-�9xd�l��jԦJ�q�f�|�|���7n��9�ٕe_mC���b��N��ūb�}�A��,�UTU�]�mv1n��,��K�Zl��6ܒ�'"/U�� �6��k	  h�8��*�[T	�*�M��[h�V����-��D��ې` �ao��a��E>��-v�u��ֱؤ�"�R�f������8ڠ6���� ��j�V�]����@�� j�YkQ�CX敭������I�$5�}F��ϔ0�:��nBgC�m��4&x�^s���'a)����x�v�	k���󻻻���#� �u8E]Q?QT>QTO������&�I���Qgg�����7`�1a���ܥ�ʑ(��⩒n�|�sr��-��5Ԣ�x؂ц��4s�E���5s�ۮ�[�;��-��4vw+�tc�{�*@���&.��h�gO]�$#�ǅ2�F�>y�Ʈ+�<AW9ٳIJ�wF��S�|�A<���UT�1`WWcG
��� �[v)�J���fa�ffB��M��nٿ"=�s�$��\�a�����n5m�H��PN�݀�7n��Vҩñ��#��i�x�Kİo��ND�,K��{x�D�,K�����Kı;�����%�bX?�%7�n˰��.����Ȗ%�bw=�s��Kı/o��ND�,K��{�O"X�%�{�sS�,K���d�L�6w�R���yı,K��w�,K��{��Ȗ%�`�����Kı;�����)��I�� �fن y��2�.���K��{��Ȗ%�`�����Kı;�����%�`�̉���ND�,K���>ͦ�\��%����%�bX7��59ı,N��q<�bX�%����Ȗ%�bw=�s��x��{�������M�8uJ��u��ն�+)*:�g;�޷�+Rw�Z�L��m��i2\��ND�,K��{�O"X�%�{}��r%�bX��{��yı,�{���bX�'��i���wd�������%�bX����'!�|�@�D5�'�,Ng?����Kİo��٩Ȗ%�bw=�s��Kı?��ntل�nK�.n�r%�bX��{��yı,�{���bX�'s��8�D�,K�����Kı;��)��ܻ[wr\���'�,K?���s�����bX�'�߾�'�,KĽ��q9ı,N��q<�bX����^�n噲f����Ȗ%�bw=�s��Kı/o��ND�,K��{�O"X�%�{�sS�,K7���?�S���sA�	�����x��Nκg$��q��V:�C�s&�<��n���x�D�,K�����Kı;�����%�bX7��4?��2%�e.��{K�I��I���6Y�a�.�nK���Ȗ%�bw=�s��?��2%�~����Kı>���q<�bX�%��w�,Kľ���������f]��yı,��59ı,N����y�
�� ��Q���(V$"N�$1@Hc0\dI�*�R@$#XD$,q 4�,K���ND�,K��{�O"X�%�Iӭ��ݰ�4�.f�"X�|(��y�׉�Kı/���,K��{��Ȗ%�`�%�-)2�)2���v�f^f]���ݼO"X�%�{{���Kİ�Uc��ﳉ�%�bX7��ND�,K��{�O"X�%��;�7v��3Y�`�k��9f�Y��su�uu��u'Xw���M��v,�v���T����{����{��Ȗ%�`�����Kı;�����Kı,��ND�,K��t���ݙp�f�nq<�bX���ND�,K����O"X�%�g}��r%�bX��}�q<�bX��IM�뻅͒鹻���bX�'o{x�D�,K�}��r%�bX��}�q<�bX���sS�,K����S�y�ݗf])sv�<�bY�,�������bX�'����O"X�%�w��Ȗ%�� �V�N����Re&Rb� ٸ���Yw�3/7u9ı,N��8�D�,K���f��,K�������%�bX�{�wS�,Kľ��ٖ0�n��f����;n�pul����^9��rk�aZ&ى�kv:}�.�ܛ2��Ȗ%�`���jr%�bX�����yı,K=���Ȗ%�bw=����%�bX4�:����eɥ�nnjr%�bX�����y�DȖ%��۩Ȗ%�b}�����%�bX7�{���bX�'��i�s���̙�w7gȖ%�bY�{���bX�'s�{�O"X�%�}�sS�,K�����Kı:C,����j����e-)2�)2��z_Ȗ%�`�{���Kı;�{���%�bX�{��"X�%���:rt�ݛrM3s78�D�,K���"X�%����ϧ�Kı,��n�"X�%�����Ȗ%�bb��� d ��{����r��n���M��z6��p��ԝ��|s k�z�sd:v�>ݬ���.1��{���7g���}ur <�{:��q.krn���Grt���^P�m;�������м�Btmh�v;[h��˯;�����n��,F��W(u ٸە��Һ �Ӵ���A!�,q�5�B[F����N���K271K��ڜOn�b|���a���;��у���D�lS�v:�a�]��{l7W<�M�ݚ���rkn�����njv%�bX�w~��yı,K=���Ȗ%�bw=����%�bX7��59ı,O{%:fy�e�&L����%�bX�w��!�r&D�>����yı,�~�ND�,FR�I�m/�&Re&*�f��e��ٙ��Ȗ%�bw=����%�bX7��59ı,N��|8�D�,K�����Kı/�}m3�]��n\����%�bX7��59ı,N��|8�D�,K��n�"X��ȟo{�q<�bX�>/��s3fL�K��njr%�bX����q<�bX�}��ND�,K���'�,K�����Ȗ%�b~�zs;t�w7d�s=R�F'�Ֆ��v�ɖ�E�bLv^S�!m��K���ķ}��oq����罺��bX�'s�{�O"X�%�{�sS�,K����É�Kı=!�v���.ɻ�S�,K��{�s��(���D�A�M�`߻�jr%�bX�w�}8�D�,K_��ZRe&Re/�ZL2�kff�Ȗ%�`���jr%�bX����q<�bX���n�"X�%�����Ȗ%�`�����7ݷrn��"X�|�"}��~8�D�,K�߮�"X�%�����Ȗ%�`���jr%�bX���Jw<ɺ\��i.��'�,K��=���Kı;����yı,���ND�,K)O��i~)2�)2����[1�^eݖ5v3*�'tc�j�u�rp��xٙ�6]��8:�B�gf�j�����oq���}�q<�bX���sS�,K����Á�(��"X��߮�"X�%�z}�ܟ9�s7f����yı,���"X�%����Ȗ%�`��{u9ı,N��8�D�,K�/Y۹���l�759ı,N��|8�D�,K�w�S�,j��S�a�6's��q<�bX���sS�&Re&R������.�m/"X�|�! ����r%�bX�g{�q<�bX���ND�,K���'�,K��Y�3��%3v]�wn�"X�%�����Ȗ%�`�����Kı;����yı,罺��bX�'�ӷ	:i.�.��,i�`�
�y_d�[�\�v=�.#�`*�=S�?{��&�9&n��I�����'�%�`���jr%�bX����q<�bX����ND�,K���'�,K���)�v����M����Kı;���q<�bX����ND�,K����Ȗ%�`�{���Kı=���yr�̦�i-�8�D�,K���"X�%����s��K�THdL�{�٩Ȗ%�b}�~��yı,��[n]�!pۦ����Kı;���q<�bX����ND�,K����'�,K	x��*+-E�����Ȗ%�b_O}�u�s%͙����%�bX7��jr%�bX���|8�D�,K���ND�,K����Ȗ%�c��������m��M��s�v՜������ٙ84���\ɛ2�!75�n�_�Cvax�nfl2�i���j~�bX�'�~���yı,��59ı,N��{�O"X�%�{��"X�%��d�zfw!w6�weۻ8�D�,K���ND�,K����Ȗ%�`����Ȗ%�bw����yı,O�&�:nRn�vm��ND�,K����Ȗ%�`����Ȗ? ��"dO���'�,K��}�jr%�bX�~��'d��6W7378�D�,K���ND�,K���'�,K�����Ȗ%�bw=����%�bX>�Jm�M��l۶m��ND�,K����'�,K�����Ȗ%�bw=����%�bX7��59ı,J� A
�A")��$�nO�06ϲ!��=p<C�kn޳�g��! �xN��P���;<{hFOr-nw=huN�wi�v�mۮ�D��Œ�q�d���!�.[�pp�d� �� �P.�JM����Fخu\�s�q7n��,p�wT�nv�3Ƶ�i:L��zw�����n���ͤ�h�2�5V�-���:ً���8�5��׳�ݣI�s���R����-_�yy�&nM.ݻ�نٙ��$�\�\��̈́+�޲O\����f��d�ۘ�볱˦l��&l����;ı,߿�S�,K����'�,K�����Ȗ%�bw�y���%�bX?��l9�w,�馛ssS�,K����'�� c�2%�~����Kı>��}8�D�,K���ND�*dK�Ҭ�]L�woy�K�I��I��w^�"X�%����gȖ%�`����Ȗ%�bw�{�Ȗ%�bY:^���6M4�sw59ĳ�@X�y߯Ȗ%�`߾�59ı,N���q<�bX(,�9��f�"X�%�ߤ�w&|ۻ�K�]����%�bX7��jr%�bX"�~��~�~�bX���S�,K����oȖ{��Y������IA��ģ�9�;[r<��'=l,�z�D�P�:;Xٳ,���vm��A$N��u9�I��"�{�"v%�`�����Kı<�'NNͻ��0�m��yı,�{����+�9��Ȗ'|��x�D�,K��sS�,K��{�s��O�*dKޒ�a�;��[�m��ND�,K�w�Ȗ%�`����Ȗ%�bw=����%�bX.IyKJL��L��yK��+�fn�'�,K�����Ȗ%�bw=����%�bX7��jr%�bX�����yı,{�l9��aݓM���Ȗ%�bw=����%�bX|*�~�O"X�%����׉�Kİo��59ı,N��%�/��s`�D��jyz��f6w��.�m���Y �N�ql�a�=^���;X������{��7~�� �H~� �9 ���MǍdɐIǠ_;V�Wuz]������*���\-�Sy���+��4~�z~��=��%K�T�Q���T��� ~$RH�����CGuX�}�@a��Y!�X� _��"@�! ��<�B2�4��Q���
�D�V�шꧡ���=E@�'�D�?"�"D���W���@<Pyo����y�����\w$Y��G#�*�@�ֽ��hwW�}�\�"�CǑe�����z*�T�{;��9�u�wW�u뚢�H��I6�p$��v!v�"������m6EBt�7Wm1�=]�M���F��#�@�v����
���*�W�wv.5�� nE�UG�K�#���	������_ʪ�RWg���s[F;��o2����z~���j�*��@3���dDY� ��@����ڴ
�kп38�?�$jT��B,�J�-����9���w�6�b����'�#�?��UUW\��s�נG�/@=�eq$@ԑ'#�����V�=Q�닺n�v��UI���ˑ���ͬ�ݸ|� o� ���[�vPyq�qdxGY�@��{�3�UI&�ru�;8�#����X\D��_L���
������W�z]k�/v"1ߋ&H�=���%��K��UT�>�:�	�����##���W�z]k�'o��rI�s���U���X"0JHI*����`�V�yx�;_\-f8����m6�vGUQ�BqͲ�S�P\x��K$x��d�3�V��|<���ok1�k��*uy-�ґ!t�lF�ZI��{�pݓ����b��h�y�s���g.�Î�m�}�ۧj�v]���'��s�r�v2�t��uR�ĳ�8��m0���=YPv��T�l�q�������w�����x~�]8����V��_�9�lW\��۴`�֬9�CF��^)�l�"��	�8����@��^�yڴ
���v^�\S"�b��y�zz^����U*l�}�@��נEֽ �E�^ǉcɐJG�^v�~� �����-�x�^��71�"�*�^�WZ�
���~��IS��@��j'��/+Y��<̀7ː�r �-���[��f�\�u=���,�[Z�%���v_ZN- B�So^�H&v:�D�9ѥ�����=���s��� k�E��ݶB�Lۻ��w�w��<>R��a��^���u��K�=���W�B2c�0mŠUz��Z�
����U�[�͑A�cN=�W ������� ���x�`��x�f^�ޗ�rT�t��~���U�^��W�Y��4qbd��8nۜ�7���ة#u�1�M0Ճ�ifl��3�>��G�Ǔ �������U�@�ֽ�uz\�cQLsNf�W���$���jI*�����K��7�3�|�C�{]���4R�OC?�� ?l��r����RKUw\��5�ܙ��}I/v#N�����ےjI*��Ԓ^�ԒUޯ�ԒK�dԒW=�,�6/���_�Ͷ���5��*U]��~~�I%����J�k��$�R��� ��m ؟'���z� ��l�u��9�vS�]��Wsg��3�ss��*� ���ԒK�dԒU�_ߩ$��a�$�Z��E��&�~��^�&�����6��M�[m˒_��UUwl\�S}��s����������>������I%�jI%J����a2	8��I%RI^���RH^�椞*(`�f����[oi�zgt��I4�.�i�������[o��*��w��Ͷ�����~m���m���9�a��#:��5�J}���njv�oG�����ø�]�kk�-��5�e�����\ԒU�W��I��RIW��Ԓ���n�,_Ǔ#n9�$��W��IL�km�I�6���y�T�]�|�B�O�0��S����I�~&����?�+��y����u���rD5��
O�a29!5$�}k��$��\ԒU���~m�URJ������}Ӂ��ǅ��<c�̿ߛl~����ԩvN����=��km�~��~m�IU%^�lB-���6훩�����E��N�p0.�p�'O;0�,:�Qc�&ڸ3�Լ���JU�:p<�N�AOK	v��v7hݵ�[ �^:涄�9ك�z�v�p��򰙹s��;=m��M�7�9�ډ0��b����>��w�wX��ģ���e48`���m����)��;�Y��s���]/l�m���\>��e����"�r����<rΟ�O�/gd�w;v�{]k\n^\]�GO�=A��D�+�6웶�O��1�ڂn9�_������G�ܚ�J�I�R��T���c��5���)����L&A'ߩ$z�ɩ$��_ߩ$.�y����K����V���n'|�A��N�34s���zf�ʩ�s���:h@yq\rA��&G#���hu�@>�Y�U�^�݃�v1+F,wy�Iz�RO�ݟ��;�@=�f�ʡ*���m��Ȥ�|�7e���s�s�F�2�u�@�$��[����������#�@>�Y�Uֽ ��f�WZ���d�q�18�&�WZ�߿UU�{��|� >���_麠�@�&�z��4
�ק��ď_ߦ��_ߞ��#�+1�ڂnM�\�r��\��v �6w�EI��$���l�*�^�{������Q=��$&1�y$O%��'V^�G+���C���6%u��e��O����-��0y$"Q�>��[�����*��@>��@�ˊ�9�H�ə� =˰�� =˰�r���7rA`,y1A�4
�נ�f�?�0
'PC�<���g ?[�h;�YB$#�@=�3@��^�}�3C��UR}s��	腓?3��	$�@��Z�hu�@=�� �rdmD��W�H:ݴ�U�E��E�ν�L����ã�d���I8�B!&��u�@�ֽ ��h�U�w��W�n,Nn��� � {9�ܻ n�_�,�& ��@=m���i�*J�$�'vh��z�m���b-��y����T�}:�I٠y�%�1W�g��o$��I���29�qAG�wu�^���l�/>�@��l��Ғ4�&8(�5v�C���oi5�!���k�s���n8���ܰHy1A�4
�k����/>�@;�f�s݂Ȍ�X�&5#�@>޻ {9��]�7��{��ڶ�n|X��D��/>�@;���Z�׬�-�͑Aŋ$��@;�f��^�~����I>�9��}���n�N�3@��/@�UU~������$���$��(*+��(*+�Ȋ
���
��PTW��AQ_�EE�EE�P��A�A�$B @�� !P(�PA
�P����AQ_��AQ_�EE~EEj(*+��
���(*+�H����"����
���(*+�Ƞ���PTW���e5���} )���� �s2}p��                        �T��"REP��D��	��*�U*B$�%)P JQ @B(�(�TAHDQJTB�B����   h  $
   ٠�Q;4��H����tH)JR'@;4Ѡ� z3�@ `R���l�t   ��V��3� ��A���O&�i�k�'J`"��Jr}�&���iu�������  P

  � 7����皜�s\{�L�W� >�y���uɯ��>�^g��ǠO����� �<�S&��A'�����q��qaӓ�w�:z������>�=:�Yv� �� ��@ 2 w��oZ\c�d��9W� S��fҕ�;e�%Ӌ�V�}=9o�K��ڹ���˾f�c蠮t�O]_x�*��{��� ��95+�x�ŕ�s�   0   
 @� ���x���o=}>Na� ����4�����y���{�p}���[Ͼy󯓯 ���^�}ξ�� �m���zk����`�ϓ��o�ӃՋ�G�w+�����    @  @#@4w����m��xڹ5:ܞ�� ��95�n;�]���_[�7*���>�w������  D  R�C� �DA�)E) �� @�%�D
��@��   "~��yRU	�#@
��'�?j�U4�# �=U*T�T� � "{RM��Pd21����j��@ 4 DHS�JI	���W)�\����_ι��?��ʰ
n�:�Ǎ�>r�TW�
 ��@AS�� ���TAQ_�Eb �
��C���K����S��Se�.�s�ę��6�0)���cB����!Lй���H�F���p��e8��
�3N˚J�57YM)�k`�A���h�h�3��ݝ�qe���nl�������(���ܝ!po�q��6&�!%����	M�0з]����s��Z�U�C1�7�����X�@�`L��ba��1�!XP�\��f���~I�~�5��,���q���o)�߹$�kx��.~�:��#D��04�!K-�N1�?�1a$ �#�WY��7�Ȕ~*"v?p?$ۗ2$JK+)� ��\$Y\�"H!����!���#"$�`��7A���	s�g4s�[���@��띦�Xp��?8턏�\�!�ʒ��I ���DֈIv�����! ����u�� 3o3�=B�Ƙ��$���ܳF�t$(am�ݧ��?�H��0�������&�E��KN�� =�e-٩�F�~����������p�8c���(D�� Eb�F&�`E�5	|rF8��p�a�p�H�.�dd$�����%��M�W5�;��%���u������7W ?BBB�xNX�l�h٥�C���'��Ďx�n�4ey����g�иKK(h7����FF��,��� ��0.@��D���L��,s4\� �	���A��C��i�`r4"�@�,IB���F;YLa�{��a�6�	.8��y�l���A	pӲ�[ �IBB��g8p�WHlK�Bѹ1�)�D�#]!��2���l5���+�$�4INZ� �ld(C	 ��,#�������HF� B$�+Xf��  P�I�SA�!  =�6sAHt�!��7��a���ќ�_\;5��N�0��JB~�=�������21b�f��Yn�#��S~��^�!$'u���HI E���s���|M����&%�$՘y�5�.	b����6��mHW@Eۢ������Ѳ:�D��@�!$�f��8o�d*c�'�	)�CCn�4�Ef��ɨoo�ɨk�B�"�ȒV4 ]�6X��.km��b��s_���$2�6l��L#�¬���?�� ���9�r6BgM��1h��KLѼc��	.vW�e� ?�Mnl8�.�/�r٣v%+,�f�!P0��jr��5wc�� �j�6Fg�u�q��-����
�6SZ6L���j�[@�2 �$���p
D�� 2F[�o�q�l#M]Vd�*�`�)_�04o�R������֎A��7�r�߿csp����"��\�35u���~޵�I F&�]����1�)Cyλ?���`���s���i=�h�/L�Eï��=��/��֫D��'�)�x�gn��u�a��ъi��C���bKi`P�����bU�!I	H��+J5�h�7# �V�:7�m���a"�89��4���� Fti��.S���iG[IB�n�F�,�0!�j-r)	�d�C�SD4Ź5�`d2ՎR$��p�l�)74BE����{��ԂF��tna�#��~���'����jr0�B6d��	�W�ra���r2d#�5�!BVE��	&.�B��Rɦ�6Ű$`8@�(B,2w���:��)\�!X�0��Nэ1��0[�+!����*����q��tH,{���L4s��%�a���X�k�ط4MHo2������kIH�I'7��0LWC6T�]����W,�A䄜p��W�aq��Ͱ�ՆL�MP
Ԅ�۰�81H$RIH��P�Ń/;Ip�`�Mhf��BBG�9�~�nh��Q�Rr�R�`���9�aL�[��m�5�٪��}9B��'�� ����~ ��!�pM�u�,w!$)0ԃ@� ������n�$�,@��$4�(u��\;)�}��\�n�ơ�!�xHr�<��\[��d�g3s������$#�FjM�*HkxXll"Y&Q5#�+�X��e.L�P��š�����_�$���HV*�t�B�ٷ�\Cp��Rpi�&,m��@���0�ȑ!	G7��8HB?�)HH�@1!�N�;BZ��CrA#[	 �hjU�a��~���H�JB��!F�HF����8�!K!��S|���[;ý�~l!����1�F[j��L�2��7�D�C3g!�B�6�&�L,"[��ˁ	��	!�	[be5��Q�
FҰ!���SZ���hB��w���~���y?^.�-�� ��R�,٣A�{�p���`���p܄��4�����&nh�rW���u�c���s��^�~�����z�vn��6[���%���$��F@�gy���%p���v���$.	�G�����)S
I5!
W,X�\�1ƬR�LlrTM�t�0M��Ə�)�,ˠ�"2!��a��q$$b8�M��A�,�`�۠���.R艧 �F\6���p�)%�D	!a@����$"�F�.݅IK��Z�j��96f`�8�̒l�7.��;i���kG�HE�nfjL\dX����I	�5IT�(fMu��!�IRI��ِ�2�+-Ʀ���Ԋ�_���yj:#\P�3\�D��2�H��Ă����&�-XA(�)B D`E"��L�`,$$b�@	 �	=�1��B7i$b�X��`@��X��HIY�(b�[$d�$B:"F�0
[$�e�!����5K%���41ݶB�o%�n� \��BĄ���"Rf�6HJi�1aq$� �d�m�bJ6Cn�5�
�ㆤ����aa ),��4��i5�&�n����#���HI��t4HB+�,)�������@� �Ā�CB��
� H�(�8�����(�J��� )�Yva�E�Hl�:�6�)��6ZjM�ha�46�� �Lٱ�k-���h`h�WI-��S �G-�d0��˽��m5�Y�?�6 t:������H�.��0�@��IYi$4h�3����I��HX2D�Bk��P0&�c�Y�����5�_�P����0��,����H��$cRBIL��� SH�Ѳ�MI��뻑�r��GӢ;+D���t�9�iăSN��-s[��vv���	�Is�������v����s��= �*��x�X$�����!��f5J�R�1ذNl �F�~4�3G�!2����iMЁaJ@#1��@4��+�Z~ z
_W_�dp�!�ѕ��P�I���$ ~ ~"E6�H�@1d9G!��1�j2�~��L;)�,B H���� ���5�B�`c�
�f�Y%IL�OԨ�i�ݖ�a���Ɔ:vYC��
�4Jh ����M�uՁ��B����!�O�::;6����HF���I�p�#l!���
H�q#԰b\K	e������8ɢR�>Q��<�L4���$�&�g� F��Q�n�m I.�9����<:~P$o�A�LcT�(�.�v~+!$�&���
F���D� �!D�á��a�;HB��0tm!$	W$ѻ7���$��I��t�Ύ�v��[����w���z~����( ��      ��}�sm�  $�L/*�[�i�a��
��I'6���ki���X�1�W�j��V��Z�BG%�2֑6����Se 8ZM�� l�Z�X
%��IKS��M�Z��A�$m[�Y�N��/Y*�Mn8Uj�bͫ	8�h�UN�yUkj�*C�[������˭v����[[�ĥ�^)��h��g�I��I��8hW*1UJ�-T�;q�����R��� ��N�` [[mm$6�z�vs���ۛV�$kխ��UJ��!�KW++tp�Tˑ��I� ї+�8*���u������NڶZ���v��r� ��M��ݶ��m��J��Ĥ�i�t� �ڋ@$-�z���h���N��  mp
B��Uj��X *���+S�*�Ut�W�y�e�^�b�[$�o ��m�LH	Em���'6ͻm��x�m�7(*�t�NʵT� aM��n�6��Ui4��Sn�
�i6P��Qlm��I$�)��}o�����am��l !��[@  .۱6�� m���I֬���m�hf���esj�tޚSa���p6̴u�[
 �-��e��  ��r�������9���m�8�L^��1��\�K@K�����Ad��G[m$��u�A���mm�����-�m� i�MkTn�j55w��Z��2�.(4�TpJ�U*ލv����@�Cd̐���X4�<��*��6�R-�6Ͱ  Ye���.�A7a¯]uS��uz'$p���m�H�+[m�Dت��-g��t�fvs%aע%�V��Z�!'���U]Q��e5�����-e�wH��Itͱ��	5�2r�J59F^؎���g �shʺ��v�U*�*�P�p��N�p �l�l�0�Z����I��'/*�
[V�-�!�܍����4ڪ�sX+e�T�����5��ҙ6���O�[ls6E����b�+��6��@�i�Q͂�1�g5������<H�;V�B��T��,��UeQ�UT��r�:*;k����$l5��h  ��җ[yi�U��N۱��m��خ�y��5]�ʀ�����tV�BH��U���� �[@�Żf�AqB��i�
iVU��m��aSf�qN��j��Vv��v�5݂��m�m1�n��@6Zmm��8l�#m��V�r��l&�u��*�\�uv�Zv�k��R��[m�r�ڶ��ȠY��΅�6����t��Y' �ku���w�sZ���[Kz�_ë���� 4�j���S*��xrRI��Wa�Wmź��-� ��\�AKWUJ�<���`   n�L�X��
�>Wkez�  &�j��6�(-�l�	��U�BN�j�Iĭ"��[��cf�����:ݭۅ�	L�4�U�/*�UuR�@8�ۭŴ�I7<y��k]*�R�U��B�,���Z��҃��JH�lۗ'$�&�Iyv^R@z�3��YZ��8����-�˅*�܁��� ꪥ:�eN���@UR�R���^�6�<�	i���nԴ���>�6!��[�pN�ɻV���ui`�� �Mp  ��[m](X Z�25n�=���\v[<:*�	��ё��uJ�0ؔ����@[\׫h$�m�[%��A�M�m�S�P��q��iyٺ��;)�M7��J�� ��X۶��^[�3	���I�I�@�N�6�s�������U�����X�"$ �6ק.m�o�ڐ�  	 p�붽����S�jNJ$�� ��$HMuT�]�[H�J�y�9�U6:We�Ѹ
�	��m�}/�}���$l��7&EV�wl��4�DP [b[��+[��O+U;J�ky����ھ���J�,������-��6A�\��"��kjU��;  	m�8UJ��hk�*��6�[c��c��Mv&��ݗ�  �t�t�kN��6 kn�m�۳l�khm���h 	�|��M�j��@���L��i�   ��p�68��bs�in����{��sVl m�6̽5EH�R��r�+Z�m�m�kdF����l�GlHl ���B�4����&��ҝ.I��Ͷm�`HzKv� sUn 8-��m��V[@�l-�^X�8�m���K9jڥ|��{���~I�Ҫ�l�5R��63+�\�UU*�.�v�*�t�W���cjr�c�� l��t��ͮ�P�����m��R8�`�j�S�Y��,��%鶻��[^[�H����r^ޓ�뮬S��j�_���UJKT���Y-�^�H��tLrU�mvۤ�m��  �l��ɶl 
������Vy�����jk��ؐ��2��[F��-�:.�eYn�;k��m���P�H��m��U��v^6�m-� �:UcE,0m�V���J�f�}nJ ���M�>��rtj���&0 ^N�	4Qi�G X�i��m���Ckh��` -�� �j@Gm&�Uce�m� �Pl7m��m �mI�M� p�Tۀ2H H 4R�'n۳����U<�C�M�V����5�M�`�k�YZ����8��.ۑY   p r�v�`     �HqE�L�!��6�6Zm� m��RCm�  �n�'om�[D��N�P [�v m��v�h�̎�JQ�U���y�LB��1UW�I��jyek�|�����e����;�	�*�֪�[LU�������b�   ,m  l��� -٢� �`�Uj���VX�U���D��H��26���vp٪ٵ��cm�  �U$�� [sr�U*���UJD��%�$��6�5�t� .�I��kl M���m��U�.� )[���[[lm�  ��E�[���s�݁���69� � ��%����UK��U�xpn@�p#m����J ���!%��d�p]*�Y��-zD���n��m)m��lM���b@ 	d�SeW\J�De�m���[zM.����j� �` � m�� f�jV��� ��:���$
�`mp�`pp	z[LGm�,�\[@   ��J�֔ȫUU*�T�%vjuKV�R�mpq#v�I$m�v�yj	2�T�P��VR$=Ju`;5PZn�Nk�Ʒkc{Cm�nծP A��� ���-���  ��-��$86ٶ��c  m�    6� �h%��lY�]+]J�YU�!L��2�V6�v�rJ	'5�`�    %�6݀�Öݦ�Ma����iYW�L��m�Y��j�6��
~>���ێ8�\��WN�l���7&uI6�k  ��$S�p�� 	�6�m�    6�+@��e������k~���ūaB��N�Va�n�-�ֵ����  ;v�   
���20Hl,Q`#::�϶�lk6X�v���S�&gg��ڹ25T�Kt���/6�*[������t��Ӳ(8 l   �psiz���e�7Ym�Jz�PM�*�E��ī`����M�p*�+#�۷*�hI��Vv�V��-Zi-���w�&�ߙ�1��%z�WPU��yBځ����%EH�Z�e&��8*���A��Nm$�Y�m���6�Z҃������9۶1r�PA5t�;���C�� m�6��n`lNiVV���)�r�� %�J�WV��53j��V��mDc\UJ�ܡ4�;KV�A�m�� #m�Cm�   �B�6�׀8!
�n�~������ $	ko^� lշm�  �ʩY��A5UU/-li'�0�$ :ٮ`�ԷdZW�A����a6�X�j�k�
� 8ְ�MU��40�    ����-���@:B۴�
�	�:�M�=T �m��X����Pp�U[GR���R]64"�\ձ��[`��m�m�G�q%Ӵ�]�a8�
5U:BV���`��v��Z/U��%*N�kX�m� DmN6�k�l�$�[(� �v�n$���&�� 8����e������h���o� 5Ɔ!r8��m��J��3#��m�t�m �3e����ض��`SPvݰ��� ��4�P9J�����d�5lH-� H3��hZ���U��t&�WUR�3\rD�R���fڸ��RZ�]+I� X�cm� � WfVU����P���61���Q�#*�Am@GY���m�p�D��7`��6ph���lG2�v$�*�ֵ�kZֿ� AS� qP�IBQS�	�J�'?����)�(�8� u6��J���E�)�H�V$E�"- . A
)+!��v��@�B!	$�HA�$	 �H�	!$Xŉ @�c##!"�`�� 0c		�2E�
��X�bH,$T�� D",a B��! Y �E�`�*
�@N��U"�D��
��@�>UW�lN���T4.�hl|�@GȽ��@:tA���`�y^pXȅ��4�u�?���"H)�:)�b� k� �z"�Q<)���
���M"�A�$]���Qê?��b 4y�CB��"!$Tv� 8���0��/����� Sj'�@8�bhTҀz:���C@A�6(��'Q���tP?"@
5M��� ���E��bgD�~6!��DH�_O�A�� ��ACJ �=�@
Q?
'� ��QEv�o��|	��G{w{{��r������GS�+(7%��Ћʡ�wj9۔か���5���������US1��O5
���\�Ϥ8y�a���˞bk��:�v��l��M͆NrH�i�n�8�Y�-�^5m���8t����X͚�ƕN������]x�m�eB��y���`�]sc��QG0#ͮwc�ր���Z�.��h�^ۭ=7�p �OR��0ᮂ�h�Fk��ú.�*]ִ�	��s��8Φ�z-!geݕ{�m���Ѹ�+ $X���M����vFí�1Ph�"M�-�md�:� �6N�|��O�5�l�r�S��k�Ni^I�N��9'�p�c�96˻p�u��k�{F�an���痳�����z�Ehfy�⍗OU���{@8�v�C�/t��cYb���\np�n��)��@l�1彭��ka����t��t��3id3��74��Em����%� s��uK;nj*�D�0uA�j�ݺ�qmbW���n�r�.�Ym���#N����
{j��t�pa4�#ΡضkD���J�m��Ek�EIpI�/K�f�v��]a����ˬA�;)�V^@�km�����<:1\�^X�n3ۇ�ŗ��3Uf��(�U�
@Mp�����Nb��٩��;'�#���\֚�k��Pg��Q����n`Ս�ێ�0��ܢ��5�&m�َ4;���Ԯ��mn9��O�z����5UJ�����J�[Q��&�eC���-�u�ij^x9@�ٵK��UW]&G&V4��o�m�'����<l�`��ҫ��=�=\:+F�v{<\j��`�f��ظ�m�sĻ&��:|��i�.p���*�f����*�e3�%db�v"�:ݷm���73U�N����c���&S��ژ��W�Cm���-�v�t���ʻ;)�r4��tc3S���B	�Em�j�,���v4��]9�;^���l��^��O�O���; 6 �� (u �݆��kSW �NH��ilOn��;eel�Bq+��v]��M⣆� v�X�Y:4j�d4�h�&�M��)YN38�;v([DW/5M(X�{N4���Zsڳ��h�y�펊6�4$�A���V7m��7k��
u���v�U+َ��Cg��[s��k[vb��fkD=X�Js�kg��p�׮�.r�<6��}�݇q�:s�㇜!�&�^Npc0?���cB�ٙl�̴��?G3X����{�bH$�����A'�w��z%�bX��{��{��7����~��}�tmRQ��Kİ}���n� <�5�MD�.}ﵴ�Kı>�ٸ��bX�'}���9ı,N��sF��R��Ֆa3Zț�bX�%��m9ı,Owٸ��bX�'}�z�9ı,Og}����%�bw?wڶ�]kV��k5sY�kiȖ%�b{����Kı;�{�iȖ%�b{;�dMı,�2&g��m9ı,K�{Z��j]h�ѫsY����%�bw���"X�%��ﵑ7ı,K�{��r%�bX��q7ı,Og��L�I[�̊\p\qp�2��6��z]�������ڙ6;3]WGf0�D�|�~oq��%��ﵑ7ı,K�{��r%�bX��q7ı,N����K�q��]�~�uul+2��|��{�K��������+���b{;�dMı,K߽�ND�,K��k"n%�bX����iə5ur��2fk[ND�,K��l���%�bw���"X�%��ﵑ7ı,K�{��r%�bX��}��ֵ�e33.��&�X�%��{�6��bX�'���D�Kı/}�kiȖ%�b{�͛��{��7����r�z���m9ı,Og}����%�a�#������bX�'���D�Kı;�{�ӑ,K��d��u�][sWN�v��{&+ۘ{2[b�V8�A�v7F^���.��Yp�VH�Y�cOw��g��u�/}�kiȖ%�b{�ޤMı,K���m9ı,Og}����%�c߯����Z���{�7���{�����"n%�bX����iȖ%�b{;�dMı,K�������ʎ��~��kS��qr����ou�b{���iȖ%�b{;�dMı�n
E@�QG��x�Ț�u�{[ND�,K���"n%�b]��}��z��Ka��n�����{��"{;�dMı,K������bX�'���D�Kı;�{�ӑ,K�w�}��Ԁ,��;��{��7�Ľ����"X�%���z�7ı,N����Kİ}���n%�bX�
�=n._�n���R�j[��i�� �Go�rd�#���<�Ce]�S����.��3$֦\�fL�k��%�bX�{��D�Kı;�{�ӑ,K��w�I��%�b^���ӑ,K��;��H浬�)��u��7ı,N����Kİ}���n%�bX������Kı=�oR&�X�%�xw�2�֮[�E5�fkFӑ,K��w�I��%�b^���ӑ,x�0ș���"n%�bX���p�r%�bX�����6ӣ" �������oq����bX�'���D�Kı?{���K���+��Щ`����Kı=���VܷZպ���\ֵ�m9ı,Ow�ԉ��%�b~���iȖ%�`�;��Kı/{�kiȖ%�b|N����d�WW�!�:�,�-�ȸ]���kv�b2�[��O�6�n�������Rv�4Y����%�bX����6��bX����Mı,K����*���L�bX�sp9Zr��G)�2K�̬Uk�˽]fh�r%�bX>���7ı,K����r%�bX�﷩q,K���{�ӑ,Kľ=}�P�ֳ-��XLֵt��bX�%�{�m9ı,Ow�ԉ��%�bs���"X�%��ﮓq,K��6{NL�4]2̗Z�ӑ,K8 �Ȟ﹩q,K������Kİ}���n%�bX��ﵴ�Kı?N�y�9�k0˓2�f�Mı,K���m9ı,>@�����r%�bX�����r%�bX�﷩q,K��o�/��.�p8�_t��=%Pm���δ�"a:M�bm��g�K<6#�\���J糗�Z�p�,�w�&��>
Yݎڛm����ݱ�ے㱫��掽	BI�l��y�ל��t�u�C�����9�d���C�km˪"�Un]Ņ��-�1��������v�iDK��3Y�6s��n\���ۧ��9�ve�2��z��� L�n�\�G����5���t����.���{6\��j�̗Eֵ��OD�,K���I��%�b^���ӑ,K��}�H���,K���ND�,K޾�������b�|��{��7��������bX�'���D�Kı9�{�ӑ,K��w�I��%�bw?{�U�Za��{�7���{������"n%�bX����iȖ%�`�;��Kı/{�kiȖ%�bw�ɽ�f��Sm������ow�߿;iȖ%�`�;��Kı/{�kiȖ%�����5"n%�bX���߯U��B���������n����I��%�b^���ӑ,K��}�H��bX�'=�p�r%�bX��_�l^��L�M9��"��n��Ľ�����ꓞNS�aK�-�����Oa	�֮��,Kľ���ӑ,K��}�H��bX�'=�p�|��L�bR�-Ŝ�9H�#��W�j&r˳��0�u�m9ı,Ow�ԉ�|=:���n%��}�ND�,K���I��%�b^���ӑ89S"X�����9�k0˓2�f�Mı,K��o�iȖ%�`�;��Kı/{�kiȖ%�b{�ޤMı,K�;�|kW2�њ�����r%�bX>���7ı,K����r%�bX�﷩q,K�罿M�"X�%��_na��շF�0�%֮�q,KĽ�}��"X�%�#�{��9ı,O߽�M�"X�%���zbn%�bX���M�h�����t��ۦ	��s�l�&�}�֕�1Q&ˋ6-��*#.1���ı,N��ԉ��%�bs���ӑ,K����17ı,K����s{��7������|�[�iŵM���Kı9�{�i�|���,OO����Kı/�ﵴ�Kı;�m'����g��w��������-�ND�,K�����Kı/{�kiȖ?#q@0ț���ޤMı,K����iȖ%�c�߸~�s]=�'٬��oq�����{�m9ı,N��ԉ��%�bs���ӑ,K����17ı,N{�g��̓Eђa��Z�r%�bX����q,K���]�"X�%���zbn%�bX��ﵴ�Kı��'�co��{][M�^X�Q��U&n��R��v��q�^�������>&�j^i��u��9ı,Oߵ�]�"X�%���zbn%�bX��ﵴ�Kı;�oR&�X�%�=��5��rk$ֵ�5v��bX�'g�鉸�%�b^���ӑ,K�ｽH��bX�'=�z�9쩑,{R�]f���Ֆa������%�b_{�kiȖ%�bw�ޤMı,K�׽v��bX���M&�X�%����jۖ�F��fkY��ֶ��bY��Q���}��H��bX�'k�ӑ,K�����K��X�"����?�|�n�ٿ���#�#�#�[Y�Rے"L�ֵ�&�X�%��k޻ND�,K�צ�q,KĽ�}��"X�%��{6D�Kı=�I���&a�A2f*�:���=�)]����[�	�����V�p��ө�~�~'��u��;߯k�I��%�b^���ӑ,K����"n%�bX�����Kı/~����l�\�������oq����r	�A�&�X�}�l���%�bw����9ı,O{^Չ��%�bsޛ=�&d�.���Z�ӑ,K����"n%�bX�����Kı;�{V&�X�%�{��[ND�,K���RC5�fL�˭h���%�bs���ӑ,K���X��bX�%�{�m9İ8ȝ���Mı,K�����\��Fֲ�ӑ,K���X��bX�%�{�m9ı,N�ٲ&�X�%��k޻ND�,K��|��s�Y�-�#��Wd��mٻ:P��L���O&�S��+�W���������Z���ujK+f`�V��PW/1�B���xk@���kK�(�q�i��V��,���E场un,��,^Z�9��es�ݦj��k��E�H̵�+[r�'/ �݀8��hx2�{n��-���j��מ�;3�\R@�zy��������`�Hq%�عq���{��Vɻe�=�Z·`]\�M�i�ù۸Ё�<Ƅ��p ��c�m�պ�f�Z�;ı,K����m9ı,N�ٲ&�X�%��k޻ND�,K�׵bn%�bX������n�j��f����kiȖ%�bw�͑7ı,N{^��r%�bX����q,KĽ�}��"q\��,O��l�c�ki�Uv�|��{��7������ND�,K�׵bn%��
ș���[ND�,K�}�"n%�b���~�z��V�G�w���ou��kڱ7ı,K������bX�'}��q,K���]�"X�!����>��jNk�F�|��{��/w��r%�bX|$}���'"X�%���{��Kı;�{V&�X���~}����s���a�8�+�4��)�X㛈�"jN^���ԉ��w���w!��&d�.���Z�ӑ,K�｛"n%�bX�����Kı;�{V&�X�%�{��[ND�,K޾ݤ�kWXfs&��&�X�%��k޻NE8���D�K�׵bn%�bX��ﵴ�Kı;�fț�bX�%�t�fx֮eɣkYsWiȖ%�bw���Mı,K������c�a�2'}��q,K������r<oq���}�~��AEͣ�F�|�,KĽ�}��"X�%��{6D�Kı9�{�iȖ%�bw���MǍ�7��������Դ���w��bX�'}��q,K��?���]��%�b{�}�q,KĽ�}��"X�%��}��O��K��^��9ڳ�̖砵�q=tbJSClWcVxq͇<�³�Lr5���{�7���{����o��Kı;�{V&�X�%�{��[�,�L�bX���dMı�{�����~�WcVF�G�w��ŉbw���M��c�2%��}�ٴ�Kı=�ٲ&�X�7�׽w$���Fd��nO�H�
��@�n杂4����8���j+*�DŐK,(B���*B
�0d2#"0b2@��X�HA �� @�V0#�6:����6Ej��A ��`Ā1``b��&#��eC�t	�C\��D��/$a$��$ �b� �$�F`8�#�dc"@�@�Ȑ� ��A Đw�F`@�$��H�HE���bA+ �D(2	1aF,��D�@�	!AHF!#!�$H���$I$Hb��)H	 $ �`	D��`1�"�$R0	���X$�HŊFD�$I$)�$0I$ �  0! #biM��	&hA)�1&V�� $ b6
�`�҄�h1��G	@��db@b�0YL� A�0���f� B(��Q�*��'�@ؠxP��
p@:��=�m:~pO!������EY>���o� [?}�[�U�vVU��j��<�Ur�u��hM}>�O��_M� ��g�f�ɩ!y�wV��ʪ�+�׀I2F���k��D����f������˷������p��vү3��k狾*��Mm����hh���O7�;+���J�C�.՗w����$?�g�@�\���ͭ%q)&CC��R���V%���X�Z�xhI/eUr�:�����URRL����w������w&�����q]�KH��+�\�.�<�ʪ�W$� �̆��
����rO��ۦ����Yp�* n��x�!���W8��ʮW9.I��@��A�H���U?�<�������?���������h�Vjj	�@�\��͇�:�W%ȥr�� �skC���������q�<b��S�k��M:���:�t�{[\�[U�r�%�n	�+3Aj���5�II/@��u��x�"�Ur��̆�옉�e]���$��@�f���w��f�£o�g�]�2��r��I/Cʪ�U&��Ty�.��Ֆ�2�	.E���W)#�r-���f��9$������?=wr�FY�,̵x�9�s�^̑xRK�r�\�M���%ȧ9\��{$�U��,���,š�r�\R䗠6�Q9d����8�����rO�!�"@�!	����K�.p�fh�2��K��Yz�w�xv�CYqmm��qa���]�qvc��x7^�cvx�������m����D���'QAȇ��e특��u��Q,�b�<��{1Ѣ�6�kk)ǐQ
,4Dl1=p�  �mf�������Eݫ�#����t�yv{l4�8�7�m��H`�p�����99]a�m���۹v�$3Xe�i�hִ[5�@�$�/}~�r��,n��ǜt��=��݌���V���9;6�1��E6$�q]�KJꯡ����/���4	.E9U\�x��n'�Ux�k��U)y%�nb�9k2Ю�̼6UW+�\�@�[�UW+� �Izf~���]��:���	�rF��-���RG��ZRK�\�^CC�W)I�-"'+3�V��31l�W)")%��!+�^ ��Z�r��r�ٮ-��S*ʻFU��j��'*���h\�r�A����n,.)#��b`q����RSv�F7`�N��'��B�k�����7LO/+�6��ڥ����@�[�H�RK�^C@<�k���Z�&kD�kYsWrN{;��j+b�T��@���b1@H]�I/@�!�7m�ʮRC��bY��-e"Я�׭ށ�{��W���@��~Z/k�&)0�F�c�=�z����� +��Hw$?5#Ba$��-v�����k�;ޔ�9[[x�r?Čn1b�iܽ�Q����{l^k.�6˪`������{��Q��<�(��@�@�����4]�@���fI	�nL$�r � �^�ur���,�2�S,M8���4]�f� hȧ�v%҈)��g�-�mzp�Y���x�6�����9�9��]�@W`�Ԁ�����nF%$iŠy_U�}��~������/Y�Z�Z���W#ly7nq:1٦yv+ۤ{3=��v�a
��7`��!�.�MV:
�R�&���}�����zS@��hW�h�U$ų�&�h�=��M�����Ċ즁�}V�U���SH��H��H�[��]�@W`�Ԁ}v���x'1�F'$Z��ZVנw�w6O�T*�}����}~��L�����[p$�h[^�33?fw����hW�h�眓bj������ cXɅ�4A.֎m�ѻz���#��<݀+]�z+��D�?%�������k�hW�h[^��;�b197�1�&h���k������}˻�;�nHƤ�8�+�
��I��~�ؗ{�s@��V�ݎ���&�!�� � �Vr �� ������-��Q�F�$z{�s@�ڴ+�
��@���:�n)21Mq�
�^*��Ո�Zf��O�����K+s<L�귡p;��9B��z�:�6���^)y]��\H�s1�vzR�V��Mqj�����j��w�/(�"�Vt��ڝ�֛a��Sn��W=���󊽖q�9l�i���Xm�W�{�t�hm]Q�:^��:G,�X����;DtN��6�7s�p\�c�l����}�{��;�~r)��'�3�܍���q;�YbTIk�ʷM<t1�p�EgqP�332���Z��ր�n��W9��r�g�����}u|H�Nc�$m'$Z�� +��g ��ʌ�!1cM�IzVנ^�s@�ڴ
�נx�UfC"Q�&��Vr �� ����<�<�;�����F)Ƙԓ4]�@�@������g���$d@�"�����ng��j:���ո�r3��"�N��1��ۙ"NG1�#N-β�Vנ{�w4]�@��^XGS�j�䞾��tE9�'|>��3ɵ�y.E�y׌���*��e��$"iG�{�w4]�@󬦁U��{��)b�&�RI3@n�Z�x����NUs��]nyZWWď#Ȥ��rE�y�S@���{��k�h���x�V(�GW;]�)��m\KѠ���q�ێ��˺� ��o���?~&�4fF�,m7 �W���빠Z�Z�e4ʬ��DV�*V�/@��{[*�$����k�<�ܳ�Ġ�5��L�-v��9�k�r ���������~�}�r��sn�8�I�"qhO߳�f/:� |� ��r �� ���ǧw���k�Uz����k�:�h����Y���X�I2,z(�m<o\��u��I�{+;�n-V�-1r6Gnh$�H�=�빠Z��β�W��<���SXGM)#��k근�s���� }]�}k9 ����w�#q�'$Z�e4
�W�{�w4_U�UR�c#p6��Gƻ �ޤv�|�����3�9���� ������{�}>ө��f���7;݀}oRy�����@z��V�@��Q'��I�LX�cf��ۍ����vM�	�����jC��^��Y̵Ƙ�p�-�Mβ�W��=��s�����HE$m�@���W)"(��o!�7�f��ջ���∘dNW��=���߿~�s9\��o!�z�C@��V^�*��J���v��Hޤ�� 5���3Y1�F&���@��4:Ā8�`[Ԁw���9�xxxxpx�Ӧ�
_� �+(J�1�ۘ������!# ��$����"�8�'��NSW���OI	
)���{Cຯ�>/�8���Q ��X�X��O��@�$F'kO����) ɤe1#�K�$�� �ġ
bH�ڑ	Z7FBB֢� �
m:�c�:A�� �c��5��Sa���4CB� D�M/��H�C@��C�ޝ�:O_w��?ne��J�I�լ년�S���m�n��ΠUM��.�Ѱ�z]���I�n�>�wC]�;�Ǿ� ���c����^�q*1�`H�m��T�f:�n,�bخ��d��[N���#؝�L�\MSi˻lV�Q�����n��	�:6���J��=l��(-����!��nUV1m����,.�1�8U��*�,]���d�z��<�òۏ1����i4;��I4��L�uX��)��e�v�=qۊ�6ҩvUZ�C4v`��b�����/Z��jz�ULq-*➛�FŌ�-�խ��BI��x��j۷e{n��:1R�ș�s������;_>x�3ZF�NIf��� o����u���<�Ҝ	�;<��p�z�x���:�p<S.km��C��cE���b@�y����6!i��3���j�����!��:���L�d�.щ�� �[�ڭ�D��QL�:�b^t�wZ^q�C[�d:�Y�N�ݵ<��C���cs�l���J���>N�/)�"E �J�7��YMz^�;f�3"�Ԛb�@�]T�F�[�AA�����;Tqc�4��mC�O>��#�NCb6���܎���+�]�8۾+��cn�W�LqT�k(�������P4m�t;n��K�-��؄��v�lk]�<=3���T��ح�ٱ�,gf���5&��\�*���v͹K�VVRZ�vf��Uj���*�e�àوԒ��y�W%�%�ݖ�/�l�Um�[;*��H"5n5,&��ه��s|܏m��&Wg��غm�-��;��j2n0�<�A#;�W�/v��R�O*��8�Ht;	7U�mnn$��h��t-�&۫,�%�:�˝�p=��Ul���Z
��[.RiU�X٭71C�cK�(-��H�)Ũ���n�Z��b�G8Z7j����t��<�R����ֲt���t���X"w������y�{��EP6���B�t��P?���O�@9�I�kZ&L��ct�����QK����x��+�[];<�`o=UB���;��[���n���E\l�'��m���3�[ۇV�k���kj�s�9�mk��Nm����y4Me&N;t'9�h�����d:��]���D��$&b�	vf�� ���6bv�ɓ	Z��l����ϖ�P�ҷ ��M�8z�^��v�d��{N����l^>Y��V�Ȏ��l�h{2�m��z���:\�#���6v�vi�Cs )$T��>4
��@��S@��hT������&p�*�������{�4��<�)�yYS�A��e��+W��{��4�3OܪK�2��z�af##�<ocQ�@�Ԁz�H����@y�.)$�RF�4-��;�f~�ի^���s@��h{�1�0n���%��r�Bh����FÝ�]�Hv�	��ne [�]G�RG1L�	�@�����-����h{kI��I�a��;���x�� ����B	 �0
�A~ ϔ��W���"�'{��m��W=n�e#��E�˼4	.E�x�3N�9_������=�ʒ<#���Y��@�f��n����	T����W�$�!���'�k�;�S@��h[)�yr�JF�V`+�zce�&�����Y�������'��v0F&Ɯ2āO�biǠwt��m��<�S�3�~�Nנy�b22G��Lj8h�Mβ�Vנ{�)�f~�W�͇eϛ�"�E0�H�7$������z���Ο�)��J W>毳���>����<�k��2��2��+�BUR�$Z[�h�kC�*���� /}��&,�`�ȜZ��0j���M=g�{&C@n�Z{E:;}�o�X"8+g��q7a���V�� ��II��]�L���'uk�b�)m W� ��H���z���I&�(�r�e4
��@��S@�ڴ
�����X�ܘB � �ޤ/9�9�c�� ��H��:d�f%����t��k\�{^���s��9�/� �����<M��G�)�y�S@���{�4�ČW64��,��xt?�>zw�b�I��#���sP�xۋ�{s���\���rFI��{~�Vנ{�)߳?fx��)�yݒ��6���d[� � �ޤur�z��kI��I��=��-v���h[^�wZdd���r'� �� �z���� ��T��na"�A9"�<�S@��߫Wٹ'{�lܓ��z�IC���D?�������L��vX32犧�v��G��]��݈���Nx(�ļ�%��d�{g����|��n���U�Wr;�C'X�P�Vu����c���ƺڱ��s`]��g`x���k��d-�6T��7G.�+h� �Ǧ��Q}������Z���vt�[��	ml��6�p� �@��e���cd�nC`d�̞��t����Pu�Z��"='w{���[�F�RD����j���3hu��y�qK=������8[���-v�߻o����:{�f�ݶ��+�ɐ�=�Ep���KN=��4]�@��M�k�<�1Q�lLJ8h���ԅ�s1�]�[z��}�۹"�HȤ�8�-��*����4]�@�{%�5$M)��a4��� ]\�z�H ��C�Qv2j�qJh�t��P�fv�GctQ�s��L�k�#њzXf��1��0oR �\�z�K�9�=�sk���d��dR�Nf�k��G��h[^��қ�$uu|H�70�G �qh����*�^�˺���h+Τ2I7�I�)������-}V�岚�,���N%J���]�s��9�\��8��'ƁU��^��$�p$yō����K�?�M�]�3nݭ�Q�mV�L��m\n�(�&!H���-�e4
��@��^�y��ڹ"�$�$����x��"(��7/@n�ց�{Or��"iL���Uz��uzo߳�M"
k�Ͼ��w���nI9�zېr �$�a$z.��]�@��M	\�.Iz�p��8��E^^^^��� �z���]�WQ��i��k��N[�i�uq�v뎎t'+VQ`�)N�u��n�t7K�#\� �z���]�.�@�Z3#s6�&&�4
��g�Ď]���j�<�S@�㣤18,��-���.Z�ur�� +�z�yH��2�]��%�z�\�R�$Z�d4�w�9\�U{Er��sk_��z�>M��F�G�Iqh[)�w�Z�]���V�xh��q��ݹ��q��䉎�G�7�۞���$��[��)�"�(����ԑ6�G��Umz.��]�@��M �mic�"	"K&G�r�@�ڴ-��*���}D5? n!�=�j�<��i9\J)%�M��:�Lyte⼑�H�ЋλM�mz����j�-u���q81�h[o@�w���y׌�7��n$�}�;?�.]�ɵ�[�KlRp"C��ӹ��jM���,����oK����>�a���C�L��Y�,�&ȯ����krm��[��m��Fsv��e���cۢ���q�2B�WNAvѮ�V��^q� w��S-˓�1�i�HKp��GZ��,6�g�A[�mM��Wgvсz�^΀���هIۉ�%:�5�ȣ�:zr��nfML����:���L\ڱ.��;��=t;h���mnzxv�O"�!��a�bi������k�h[)�Umz�af##$x�Hi)�k�l�H��M�mz.���NM��F�G�Iqh[)�Umz.��]�@�{.�MI w�C7� q]�\�� ]\����vĠ9IY0�=��^�ݶ��ךM��>�s���J-,�GN+ngG��CP��u�f]��֮�J���aPڐs.��A�������~���O� ���Vנr���9z�cĜ��2�Z�4�כ��r�9ʪ�"�^�����-v���Q��q8I$�Vנr���-v� ����,�bpX)��M8�^�z�ՠy_U�Umz�af##$x�I�3�����k��ϫ���߸�=�]���s-<��b��lۚ����p��� �v"K�/ˑK�^�UV��㾵�4۽�޻����"�/\�f&��)��8�
��@��W�Z�Z��Zz�@r ��Ʉ�����]�G����f~��g��#!0&�81V��aD9���mM�DX�k���i��� ��"�F���F @",� , ��B@ZJ!�D�hE�"E!`d#X� �@!!�
� �XB#21�K��H"F)`�����A����T�
���hmX@%Q<����)D ��A��S�����
����v]k�;�T������c�8�ur�������ϱs���2<��	���}V�U�����]�@=�%��`�QE��~s��������V]��-�9ضp��-0�ݴ�wK��N��U�����]�@�@�㥙N?M8�_W`��]�@W`T�=���	���#�-v�����k�9{�����W$��$�4��<�\�8��.}]�y�9�5ޮ@�؆IR���*����^�k�hW�h��bVF�?�Bq����9�x�Y��;�'��H�i�t���g���""�#&G�r���-v�����k�;�T������C�8����� +��W`>���	"y$Q�qŠy_U�Umz/z��j�-3#qcX�Q7$Z��������k�^j=�x*2�,V�/@����	\�$^���n�y��+-.w���5X�v�n�h�ʔq����[]�щ�qmW.9�c�|��ǃ厶Nζ�*8ZpqƼb�hư�Fx�8ܝ��wf�ն��U����w-�bP�bK׳��� �����'A���d��;'^`��r����N��v)��öŸ��g��X]�zݏ3�w[��K�E�lx
c���Mn.jYSXc�G.D���D��f������d߯{�۽��H���e��ꛈ�pؼq͡�^1�k6z�g`9z�|v�Fm�ָ݈q\��Ƞ�X�R:W�Z��ZVנr���<^�I����G��qh;\�8��.}]�.�@/׌�InchhN-�k�9{���V��}V�޻bP���?L$�@��v �� ����vn��s�F4�14��-v��_U�Umz���ۘ���kHdC�5�s=�CسXxI۱��gs��ذ����q���R(��@���h[^�y�@�ڴ�s���q7rE�[�{7��T$@ F �D*0� g��I{��ܓ��]�{��.:Y�	�
~�q��� ������v צ��p��#���ɡ�+e ����r��t�)ɵrH�H�9"N-�_\�8��~^�W W���L�x;V9H�d�/hML�t��ʯrB����lu��m̦�{k��*���1�m����r���-v�����vĠ98O�	#�9{���V��}V�U����,jf,n!�=��h;�Z_6r������*�b�o@�v^���j�"$q���@�@���^�z�ՠ��fF������{��ϫ����k�7��?�v��ڳ��ӮV̐��d��:X�q�V�fS����<n�.�X`�x�77� =�{ ]�@>�k��ZGfL1�G����#�-v�����������NM��(�ɑ9"�<���*�^��ޯ@��ZwI��&ۘ�0N-�fb��~z�d��mh{�r�K�\�����w��"$j3&G�{l�-v��_U�Umz��İ��	�M�Sp�vk�X�T�<m�FL[[vqYm�X��K��9F8�@�ڴ+�
��@��W�r�Z���F܁��� |� +������ ��V2'q�p#��*����@�ڴ}���,��B�Ǽ����>ϗ`���z���H�Ɇ6H�6��#�-v��^3@i�z�o4���s���$���ͮ�����e�[XI���A.�v����t�7[�5���W3EY�-$u�[[
���r8;5���E�����[6�*D��7%k4u^Y��^�7ER��e�r�"8��z|�����ax 0u�F�N�*�J`��q�]������rnν1�L����y;	˄��#���zzzv�#��窒��)�L[�����w[uƝ�Kΐ�gc���ű���i5�p��D �hM��nvW7u:&��x�Ȝ�qP=�O�@����l�-v���q5$L�!�H��@i�{�$�3@��Z{׵�w�lJ�4�鄑��٠Z�Zw]��k�=��X�G�b1��{ ]\�[Y��� �^�>�U�<��HېNH�Vנ6�@n�Z�s��R�hU*�Z��\�5��b�{S.�6�5�[&�s��g�j[`���	@$�#�p�� �}��@=W������z�Q�3{�]9�f\�nI9�{[�W�~�Pvo��Z���U���#� �<��3�����g +����=96�Iy�N-�n�U�����-v�����'2H�A$��k�9wW�Z�Z�����TV$6%$q�$�Ҏ�˛�t��IuF�K ���Bf���\�a�[5��郑����-v��n�U����5���q��k�h[w4
��@��^��>V(�G�I�NH�-��Vק����ҽ�j�N�c$qc�`�s4
�w�uw���9U�/d�V��)���HS�oN= ��f�k�h�n�U����	'�ƢDpY#�[��ľs*#:������v۱�#<�W�m��:k��4�xa�����h[^�{�@<��ڹ"�� �bqh|��������Q��I"jH�&L�*�� ��f�k�h�n�޾�(�"&FL�9�{�y�7m��[���r�H*����\�f�~��Gm٠{_T����8�CM9 ���Y� ���]�{^��n0VwD��-$����i\l���VXɭ�씮ۑљ9�d�z�*&�U�U��
��\���� Rر�8��&F�� �٠r�@�ڴ-����Y�	ą?&�i��.Z�ur곐W�
Ӷ��+Wab̽��)2E�{$��m�.���NM�"�� �0��@=Vr *�r�`���D �d tC��*yVo�$��	,P�71d�wo �"g奅?�M����E8���� �#"HM)��"@�l`Lce�[J� %�e�VB	*2IBB5:�D��R3`B���R���r�HL�S��N HЂ�lf��p�$eJP�dd�*B� D� �BFHF,�a�$H��`AL�$ !�����B�f�ȤE4�
D��VP&
b&`�@i�r̿������]��Kf���ήݛFx��g@�[Yݓ�Л�cv�S�Y���N��e��1��yA��6S����wf�mچ����j�'\9�Uc<����2���q�9���^���¥��$�U]m�D��:����mԀ������2l�:4cv�D���Nu.j]��_�<ki��ܯnm�;p3;��pv�pJ�q�k��s�y���M����v���\��F��Y�c�۷�����Wkm�ְ��pQ��vܠ��a�V�yk�[�q�RpsG���dp�n��ԁ�����m[pn�cݦ�Eˎ�X���L���n$��9K�.�P!j��(�x6(����j\��B�n�Le��9���3s��Ѵg�y�G���ک�����@�e��Lh�r��b�v@�N���cf���F�y^��*�:��J1�g�5��f���� ĕ8^�tv�y�zP�m��T�
�n�q�
m��D�� γ��Ĵ�灱�\�k`{�u�ى�\��AkR�;!�Yӝd��1�be�m��+:-�2U�[4@@-��=0��[F�j۫���ݍZp��*�5m�v�\�r��T9�,��+˶	u�6�A�iwg�`����aXu�s�in8�\�P�7j)ؚur=m����
�L"g�@G��ҽ���L�6�(��՜�-��MR�e1˧p������0NI-�m��u�Țɔ�
Z��2�WT�q�Glm^i]��qN#�(l6����8
�d�Uum��sE�5Ķkt��'q�b�[ks�\�)���X�e�8�v|<cX��qó��L�\����a6lc��b���pt򹍸/X��k���Mth�v۰��4U�T��Ps=���pX�U��!��x�tl�]�f�뗒�l��n�ޜ��р�.���;*:��QG��'q`�]��ȨEȦ�Mn�rZ[��-ѮT2ҹ&��ӆ�0P�r�Y3V�����O÷��w��� �D�wR�K�32���X#Cc���Z�m�e�Ż��.9t���МY�8y�:2n}��f�����f��7o:/9�[^�rk����]����۟U�\����^��,���`XT�V�[���N�ݱr����.i!㧣 � Xm������ƕ�͛;ce_Mۡ�"�����m�^v�ϲ�����;x^ٍ�g��}tW&J{�ε�A$J�:�1ѝ��#�/F����ng[�tQ��/,�"٣:�*�������� ]\�z���zƢ��29&�˺��j�<��h���}RƢ?5X8�.�@=Vr *�r�`]��H�I�
I��s@-�h���-v� ��2GJLr'9 { �k�����@?s�s����f���WX�3�4`�͘�k%��ǃ1ms&^T��k�hE�۬0Nv����_� ]\�z�� U��D��dQ4�R=�j������*<І�y'���nI>����9wW�{�4��)2djD'��r *�r�`��h��{�ә$���4]���V��s@�zUc��!��@���ur곐W����[u����.z�P��uք���X!$��D�h1S���5�����}���h[w4�g� �ߞ����Qd�d�I ��h[w4�f�˺��j�N�c�x��!"s4��@��]��W++�p	U�W=��.uh�6��<��%�awE��М�r���z���<m�h}y�w�Yo2 �EM��@��Z��� ���9wW�y���[D��ȤK#5�R�<Ɏa�m�jy�3�uq�i�]w2�S�^IRd�〜Z��� ���9wW�Z������'$��a$� Z�r�`����O����Z�p�"�,`��V��_U�����I��9�}����"�W�"�///@n�ց�x� o�42��U.Us��?g����v��@�u?�Y$�$�H)$��Ԁ^�.Z�v� ��s>۷���n�Gֺ�5�L�4�O�mA�L��v�AۮM�a����|�䬙�D�C��￦�˺���h[)�ylE�����6��.�����~l����w��@o4��o+ WX�Z�e��k@�f��II�V���y&��D�L�H���<�3@����w�*�����&�,�7$m�a4�f�˺��mܓ���7$����A�z��K�R̸{n�C�n�:���N�A�m�d���[:�Y��+-�-Gn��8gr��{Gkun�roi�L)z��^\r6�Y���w#pϪ6՛/Kd��!XcY��y��5��"0l5���<��ۭ��VU�wf�u[�V�(�ۨ����!ꔺ�b���'`�1aA��fC�ٸ�۩�l����\cgh�Tr��8AT��O�3��as&^a��:.��U�(�m<o����s����l��FV� �'6�ň��fc.ϯ@n�Z��>����X����@����Ƣ1�����]���H�L��I&h]����RC�ɬ�L�)$	����O� �٧��%˪�[e4��b�!����	��q&����^���h7��<�"��N	LClM94]��~�\��l<�2 �y�x��@�<�v�xz���WC��kqh�ѫ�|q����F�3�G��ǐȆ��b���M�q� �y�}�r�^�E'נq+K�ō�)�4-���?g��f�˺��)�g��ċi��2Hܑ7�a���I&h]����<o�wޖ��D)&�߿g�ث��}���@��M �٠w��LQ�ۏ2��yyzm�h�\�{&��	$��uz�i�W�ȱ<xHdFD�i�r�\]v({CH�8�b:���9�ŷF�S�94�/K�q��!�yl��[l�9wW���U�I2 ᅖ�.լY�x� m��:��zo�x�3~�*��UW9vw�g,W��.բ�^f��^�{�צ��8*�@��}���nI>��:��VL1<�&���G����fb�l4d�hm��޻�=�V��Yv^�b��<o�J��)$� �ߞ�k�hzvLHƝocp�s�0qD�t��ʩ�rB8`뭶�ɥ�<�� ȆI�&��#��[l�9wW�7m�\�x��2�Ʌ�^��ia`�3@��]���RD�"�=�!��7�������4�����=���-�e4�f�˺���M�Wyf]�ᗙ�Bs��� �L�:��f���b "���*���r�d�ՠ�Yj�Z�Ř�0�����)�r�K�h7��<���ݨKk!Y�Wc6H�fHuqS�͂�;\��pt���z��eڼ�.S<ڼ���w�7m����I���,�cy�'��@�ڴ�hm��޻߹�r��U]�NZ���F�dq�N-�����4]���V��r�Ld�H��8h}\���4���7m����a�>��8E2H�)&�˺��������w��@o4�U\⢹\�We��Ots��-��{$&Fvn��Vx�<x���Wn�$уj�����a��m��k�l��2���t�ݖ�8��
�v��i-�j��˺�v��9��ֺK"gD�EշLE�ӧl��e���t��m�;��!Gcsm���ds����A��D����Wg�A%��J:�ؓb�ǃf�c�$Z���:k��8�����%���ͣؠ�Eh2Y�P�g�m�r4�u�iX�m�B��}���yl��[�g�Uo�@�ؾ��QȒp�I$Z�Ԁ
��\������s0?~/�kpm����}��h���*�^�岚��Y��LQ�񡥙�Wz�@n�ց�x�	��R9���,�cy�R=��h[)���.��8��C7%�z�w�|�]���i5��h�c;i�뀱��{9�س?�g�Zil�8I�7�~��������@��]��+�����6ɦU����j�2�Y��$���o`iJ��`�D�"/9=u��rN߽�nI�{^����~؜�D�)&�U�=�Z��K�2$��u{�jŕv�^f,crG�Z�Z�e4�f���ٙ���￞��k��7�9�&E#qh[��>�)$� i�zv��:�vY���8�v{F�n�ë������ҷh�iz��X��wo����'%
�Xf��I�Wz�@n�Z�x���Ӓ�F�30�乭nI�����(+l��h������]�w�R�Ŋ��.���{��]�9�k�s���$0�@"��'��b�B�L� ����b:;��>M�q	 "AR- ��*Q �  ��ĉ$	@�4�����9�*��FA��b�BT`^��� hCb�?�
i�|�t����������/-�h+��/W&ՑL�w��+š��͆�I&h��ހ�ڴ{��c$�)��#��[�hUUq�r�Kqh7��;Bby��vf��mBIq�����3�K�����n�2u�	͛$�"�J>�~Wz�@n�Z��>�9�]rՊcdd �����@��M �٠r�~��"�����'R6E#q@>���� ���]�.�@*F��i�1�$��ؗ�_��U�=$�����(��H#�� D�QU�߹��'~��NE&F������9wW�Z�Z��hm�+��R�i�J�1,K�W];���>w�F拴�6�m,�'��&T��N������u�dDƞR>����-�e4�f�˺���4Ҳ)&I�7����x͕�H$�4���4�z���1�FI��#��[l�:��zJ�QI/@�L���z��^yX�`�ff���s���/@��z��4?�����*��LS���1I#��w�}U� #�4��ށ+��x����m��� � u�]ZՐ��[������k=`8��=��U��ȼ�.A���{jN���+��,���1%����_cȕ�8������v�/S�c]mX��t ��������N�Ɨx�whڽn��9�[n2I$�izV�s�L�ݠ�ۀ��a��-��a:�n6�Ǝ��]��ib9�,��ۆ�Ȃ�ӧ�]�޹砶X����^rk���%'�μL.WI	�q��k̫$���gv�%v�y�MR�$�2A��߾�z٠r�����⪤Xԉ4�r8h�f��۽��z[�l��������
L��ǉ�ɠ|�����WZ��S@/[4GΨ`6E�7�أ����h�y�u6�@<��ZVD�Rd�LmŠu��ؾ�}<������@��;����b�Os���7%���'�L�p]�z.%�ێR��.�p�$n8�7�p��������@�e4}�8EJ,JI�'o���qE8 |�����n�w�|h�f��ޭ1Lcx9�B�G�>�k@�x�'9Ĉ���%����M�Q�R&H9���h�f�ɷz�T��/@#"�1U��v�/*�ސ���v �]�U�@>�y��{�ո�-y��e����K��.�᎞Q����7Z�\t"Y��q].Q���4���u��:�2W+�rf��ï��dD��!��
�נu��z٠r���;��4��(7�917�~�|h�f����
�נy�+��I�1��4>K���@jIz]n�>�+�ɰ�;ד��.EX�JI�r�����l��>���Ty
�X��
�H�B̢����]�W
�YΙ�;i��ۥ�bC7]BE�2ҘǊBQH��~��l��^�h��@=�j��A���A�#�9�f��G&hI/@k����W9Ig���B6�s��@>�}4VנUֽ��h��O�RF�M�37��}��ʻ ��@��'<���瀬PWB)�L�}�nI�e�z�$l���7�WZ��)������qzp�Dв'd��.�95Ρ��Z�Cs�j|��v�s4l9p(�Af�&�7��e4��@�[_߳?x��~���_i1�F�m<��@/[4U��u�@���͝~�<Lm�`�M�9}��@��(���@;��h{�X��1��1�)�WZ���4��М]�%�[�1]�L�qH��)������
�נo�����%�6��D�A
Y��mvad&��晵ϵ�hlclD�p�.k>�鲭y�WvnK��غµ2�k;r��g+���
��wmq�n'�f���u�23�\�.� �D�,���M��m�#i���k�q���͓�|l�Zva�xo��.8U(�<��[�H��p���ɧkm��3�<;
��nƇ7�N�p�t�ғ%I�~����|���̫˛ӫ��b).kKbz{v���h�6]t<a�v��������Q�B�J�Ҁ[��`b� r��-z��O�RA��Ęܚ���
�נwYM �l߿~ď�U����1�t���'%���i�r�(���uG��=^�I�dJ$ӎLMǡ��?f+�l4���z�]�u��=���fdnL�M�]k�=W��*�^���M��щ7[�#��1)�I��Bje�O���گd�i��˝gr��g����f��	țxA)�w��������*�^�g����1��E�bs4����s��r��9��&�ŠD���s@�w%bo �!�@�����z}Ĝ�k@��z �����W�wx���+��_�>��	��k@k�zW�h��W�) ؛Ʊ���׵�}ʯ�U�O��@�\�hu���ϼ��+�O*3�z��:�e��Xq͂.l��������&�=��Ddx����*��\�9W`����ԚRD��qț�@����?bDNK�sk@k�ށ�OL�32�2���4��*�^�׮�ٟ���s?��@$A3 �3ziU�!�T��B �A(AJ����_����w�?��䟿w���I�$�&��R=�]����_U�Uֽ �{�YCk$���hsw�}�}S�/@�O����k@�8/�~XxIݮ'0ɔ���ӡ�����WL�y���@�r%��[Y�~m�~�Z��w�u��J�NK��-a��m�ۉŠUֽ�]����_U���31#�e_/�RA�f%��/@qͭ��z}T����"r^�kV��a �Mɚ]k�:��ܟ6?g��6 �66
P?�F .� 1Y����؃� � � � ��_g��n��M\�ֵ���؃� � � � ��{��A�A�A�A�=�ٱ�A�A�A�A�����A������f�A����w����s��2t#q�ӳ�Y�j��\c;����!�I;X.�׬�s�i�æ��2��A������f�A����{�y��}�Qy}�}v �666=��jL�ֵ�s	�n��y}�lA�lll~�}�lA�lll}���؃� � � � ����؃�
� � � Ӿ�ڦ��fj�d�ѱ�A�A�A�A�=�ٱ�A�A�A�A����b �`�`�`��{�b �`�`�`����<������e�]:�jL�SE�ֳb �`�b�1D� ������A����>��͈<�������6 �66(%���͈<��������jkXk2ff��W5v �666?g��6 �666>��p؃� � � � ����؃� � � � ��{��A�A�A�A����dC����=����.� x�����ǡ �P����!	T%$�K:H1ь �	Ƅ�1\���#�"�H��$�P�BFE�,������� *�yj�^�l݅6.%�rFgF�F볍�zm@p���;��Ԇ�۝h���`����`�+��G +�mYT�.&'\膩��(�zc������
j��gi�h��[��*��Zڪ��(��ۓ\p���c�S���S�e�R�� v�5&�<P;��v�;	s�2�ZJ�����Xs��y�n��vS��w��,�W�Y�5�]�c��%�.��;[Ÿ��d�7�ѺG[�8��v�gT�h�����:��Rt�t�}d��]*���u��l[B�#Jˎ�T���!cN�jv`ݖ���^S��1,ʢ�v�bv�q�;[�lK`ܹ��KLh;4��!�kNLח��k�`�F[�x��7gs�H���z��K��|e�w.\p�f.���d�:��0�+iN3�˥�R���J��c��K�����[/l���VԌ�(�Z������X5� ⪢�ID��x���q=��M	ڥ�W��SVŸ-J)�8;�vH*�ǧ��7<��� �cU�3�Ù��uUͩz����b�s��+٬nss�i�UTs�:]��x�A;u@,�en�Ȳ�#8����,��R��ͨ
���û2�_3lڹY�=��!��Kgk�p��5���f	K���a��]�#�U�T�����7�*�L�{gj���zQh7ls*����A��v�Z����D�ՃY��l2k�"t�Z��Z^�䀕R��X���H�ej���L�UmK�E�q �%vb(��l��v%H�gS��&��bC�͉kMZr�]�uL̰�t�kqv�hquĔS��P6�{L��=T]'Ƚy
��f8H�8�]�s<J�UݏN��c��;`�h�v�q@��U�r�ꬷ=5��C���j6Ύf��m*�Rc�͉V�^��Gvݲ����X)����99��8BU]v*��c.�Fǩ�`ی��օ�:v��]b�k-֍L)�In��5DO¨qU�q��mh�"*��ׅ�"��@���a�:"3`"mPنzK'd��K�(ݳ=t��V�h��l�N�W��Hv�ƶ���ek���7f'0���%E�z���G�;���b��!أc<V�<�JK��
wŉ�&3�Tk����ͬ�Ů&��ɽc�n�غ,���v�4v栻^���j�^�<:%�K�i	���&,spғ���u��a�1,�7�msudá�km��Z9���;<m��Dڙ8o�f�ɩ�u���ZԓO\\�-�!����t�M��q��k���t�d�֦e���fk��Q?A����{�y��}�y}�}v�������͈<���������d�5ud�-�֍�<������͈<�����׾�y��}�y}�lA�UK��?�B�t+U�~w������7{���}�}v �666?g��6 �666>��p؃� � � � ����؃� � � � ��ܚ2kZ����3����A�A�A�A�=�ٱ�A�A�A�A�����A������f�A��P�A����b �`�`�`����j��K����j[�f�A����{�y���6 �666>�^��A�lll~���lA�lll|w�e�擄�&��4a��ڻ�=��,�lҖ1[؃,vmd�r���f��ꚺ�ִ�5a�3F�A������͈<�����׾�y��}� ?�����A�A�A����y���_�t�kRfj.�k6 �666{�{��� X�'�l"1 �X�BRT�1��b�	"�����D�ĀH���!" �x∞W9U[��>��d{Z]���� �2���MH�N-��|��w4
���:��@���W�)#CMcM�����9k�
�r�s�����|����0	&�nL�*�^���Z ��h��4���*��%�ĻTn8��7�#|2�m&��=�և�`;n�V��s��?�p2|0U��j�����������׭���4
�נ{�]&2H'��ƜZz٠_zS@��z��[�$w_����4�D�$�>�|h��I���n�޳@3��VGR,�#���h]�@/[4?s��<� ���e�P�
�Ff-��@�`���� *��o��FR�XѮ(�C���{N�A����AE�w\+WHӤ!�!�]�r�$�^�+Y�ur]�@�]s�q�McLnM�]��h_U���UUS0	 LI�3@}�ց�}kI��Drf��Z����d�Ym��@��� �l�;�����0��绞�ܓ����5�9!Oqh�f�׮�yڴ���-K*���dM�cr
 ���ufn{m7d�rq۷L\�K�Dn�ft�Q�7�Ē�hm��/YM��h�j���Ց�I��73@}okbC���ԋ@�����r�I���qe�.��fa�9n- }M�%$�Zrmh����ay����f,W�Bs�UIF�Z�mh��u}V�^9���H��@�iŠu뵠J�r�� r�Z ��Z�U�����E��F)��HN$��!�.��u�h���A.�[��b�<YA�s�&�������Nؑ��r��3K��j�NE�뗐����=�<kT�	bnJ�h�ƦL��\���;�pm��rjKpV�m�����]N��Յ��zgڢ��[`q�8��rO-�N{;d��*{�SbG��;VrCf�f];=�H�{Ӟ
`�N����w����&��i����m(+s3��8�q�[�����<�qX����]�.հ -w�����
�r 7 �����p�H�I�ۍ�@��� ��Z^���)�yܮ�$�D�ƜZ �\�V���Hv� ���(�r�BIH��w4�S@��� ��Z��X�)�q���h��}UUUT�8� �H�����~~���W/I��v��x�q͚�W5��>���i�V)��<��.�݋��a�� �� qrZ�@� �:�H�H�qhqj߳*���r��ʬ���ց�hwִ�ί�RF��,i�Šu빠^��W�hqj�*��ـ�H	5���� ש �� QrZ�@=�����"M��p�:��@��V�׮�z�h�%Ռ�Lx)���E*��qwkY�"wm87OgT�'n`vj��E&<d�7$i�4��*�ՠu빠^��W�h޺〣S���H�Z_^��r�I̆�帴
��h{�b��)jc�����'}���٠O�@蠜C�"�E�Iٵ����V
�+�oz@+���\�V���H�ή(I#��)"�ŠUū@��s@�n���Z��&̩�F�C\k�ȳ�pى{N������5�c<,qv����`��W�)I��lqx����^�s@����-ZV�[0	�i7&h���Ċ��\Z���O����${yE[$K4ӎL�>��� r��
�r ՜�{o^��7r�3,��J�h}\R�"�sk@}oM��I?@�&�}�z�I����N�G&qhz�h���9�Z����>�N� P���*E�]Ɛg����:���u��A�=�ݸd���eŞ*�w�|sbȤi��3��@���W�hqj�:���xu)�M�7��n��
�r � ���R~�<�$�U��32���fb�x��"�+Y�^��\�.����p��9��orZ�@�`���yJ[$ZRZ�e�f	%h�̭ j�]�@�����}�<��9϶�w}>�k�n-͹(]Ŏ�xK����9wb���v�-&��v{I�$�.����ά;����dnf��nݲP�q���)l��Ր��C�wN�p۷o	S�i���P��z�˥�q�(����}�^��XYm��/�@s����;��u�[� S�1�69"�v��m��X4�*kp�ɩ+�v�k9�F�^70��X+�c�Ѫe��T~P�vټX��]-,o+�s�}�9��ֵ���g�n�n�"eΨ,r�3_ͷ�����6�N����k�ɚ���t��WxI�6��@��V�׮�^�h_U�{z��(�slxcq�z�h>���*������@�W���{ה�)�6�1	��*�^�˺���^�}�s@/�:��Ʋ<"��w���\�����}~�ߧ�ZO��߿����r\�u�ٷ7fS)"�n��9ztGWmmX�G��蘜�rԃm�Ԓ�v ���g 5��]�gs��u��2�L�]k7$�훪�`X��Q��n}~�ٹ'��}��yS����U$E�젻ĕ�һ�4���u{�zNr��U���ցު:��"DM��zي��=�_���빠Uz���<D�G���o{�8�`���8�`>��s]�6�S��##��2&&����H�n��E�yʚ9���wf�\�I:��Kn? ����U��^�zYz� �z�Y�H��1���*�^���]�S��׵���H'Yqe���,"��u��e���}�	BI�)*@���ʄ�Ɖ(��!����ĈR�%#��-+hƁ
JJ�RW��@�`��s��F�Mʙ�E�i9�!���s����b�, �ia�HV@`Q[p���`T`���PК�5$h��E���P5Q3Tj��,P�L��B� dB0`H`ԉ�tP����>E<pA���^/O(�D�#�+�D�������r������i����݀9ƻ ���ƻ�9�y�����_���dy$�@����U��^�zK�����7�Q�.�W��^���].2�m���덃����.�."���Iwl=�xVߛo������޻�>���\���4�]�c$�6�dq�������<�)�Uz�ηcx�"R'"MG�}w�x���Uq(���5�/@���1�Q� �M �C�?f/~��|��ٹ'o��7'��T8)����}�7$��}1AI��3�4
�W�~�����#��x���<��8'W���w2-k�e�z�mv��/I�M�Z�F�i�H,i7fD`�")��ޯ@)z��ҚW��/.<#��/0��=n���U}U�]��gƁ����r�����cq�O#�!���@��ϫ�>]�9��lO	m1���~�_;~z]~zOmz��4�Z1�$1di]ٗ��u{�z���~�y��ٹ'�ƚ5�g�-.d���Z���6��-W�i�Ù۰ī�wk`;I	��.��^�8nܢ�]��x����$��9{Dl��풣dk%G��r˭N����df�]f���|��>l/̛��r�@y��v�z�`�cc�,Ja�]�1[n�<P�A��n����ԣ�g��vJ�'����4.��=�-۴Y8���]k�6V��;nr#�ݹ�휼-����޻��׽�_1��e6#��s�\(�KWI��	��[�6����F�o:ixԉH�hr= �/���<�)�U�_����
�����dǑF���Cs`�� q��.}]�	�� �[1AI��3�4
���9{���q"��=�!�u>���0T�(U��w� ��v #]�zޤƻ �t�xI�����
^�@��s��r��z�@<m�ݖea����j���5�ˡ�&/uv�����K���(��;�H��qac�1Oͷ������vs�� F� q�;�s7��m1��Uz�_��y�?6r}^�R�z��4k��3$�F�l�^���]�]���{C@�9z��cx�"X���'#�
^�@����U��^�z�&<�5$J65����=k9 q��.}]�9ƻ �/b. Ց~$kI�&L�.�����M�&k<�wb0��v���n,TX���I3@��z/z���_� ����W��2�(��G�r���*���^��W��/.EF��Rq�e���SO3����fa��D~R"0T��b�T���O�z����*�u1�LPm�y�;��H�.���9k�ex���	��G�mz]k���ހ�����eb���n,����*�MlJۃ�5�]��wf��D� D�4̒%�i6�#������*����S@��^��cb$�aND��@�;��/YM�mz]k�-�cȣJL#CK�@�e4
���u�@�;��;޻�
H��x�1]�W)K엠D���]�t@40ȇ�J���~��v���j38İ�#�@��zY�^�z�h{k����ԑ~j&�)	�,u,ʹ]$�t���::F�ː�-�Te�� �Y�������
������*�נUֽ��S�DM��#� ש s���v �-v �t��56��U�@��z}��q(��zs!�z�t��b�[�g{�*��Z�ֳ�>]�y�v<iI�H9r=��@���hz��^�ށ|�Nr�+:�������=Cq�Hm�D6���n�<�@�7�K��\�=��RF�����y�a�m��m�6��س��]a0h�v�,v6tty��u�4K2;�v:�I`��l\�e��]-�Au۱�9�c�3����ֻq�:���;�����.(�(�ն�7#����by#K�%��m�e	cQ�uP&��q9;;2�r��v�:k�&���qMn[nK��&L��1r�v%��b����3�,W`�-����vݬ񮖤�cȣm�A�K�����ۚ^��^�zW���븠����ǒ)&h��@��W�U���[w4W���F���=�uzY�^��s@��^�}:R(dN&�����������@k��נU�u1�"M�Y�#�<��h5��]�9ƻ /�r�o�N�W<-�w�5|4���K��q��i;vzl�\.�%�!�#N�{p�[*��ߛo������� s�� �Y�غ=�9���W%�&�Zܓ���o��o�ost��z���y�f��vLiI�H�7����]�z��ϗ`-v���EmL�Ɩ7��빠U�@��W�U����{�
H�r)&h{k�9{��guz����ϥ�
�ؽ�5����[��i\n�X�ʮ��q�l4g�Z�<�'S��%"�����
����җ<@{k�^:P�"�6��7�g��o{8�*�נr���� �+�R"	����z�Y�U�O.fy���|�yʮUsı�zT۽��*�WM@M16�Uֽ��^�VwW��W9����ƀ��Y�++3�V+�e�>����[Ԁ9W`�]ߠD��7F�gE�Y��BJJT;w>�槷=�] k%����6[�� ���� +��W`zɋ"���A�$z��7䏗�|�
����נ_m{��H��NIw��vs�� Ev�z������IM��$z~�__��|I/@���h*��}�r�QW1d����@�4�������<�w4
�W�r���=��%���J��rF�4Ys�ѷAz���i�s�����
ô�	�M�X����<�w4
��@������EQ��$�dʰ�eһ�7w��ƻ ��v ���g4�X��D�&&ؤz/z��mޓ�I{��"�^���ebY�,i̍��zYmz���U�����z��(�r6�H�/Y�������W`���<�8s�P:@�.
�h�!	[KR,�b�Ry�	�(��X4�IT$ D#XP�Q���dB!A�bE8���l$X����?H�ň�"@��V@�bbȕ Y"QaH���6#$ HB)%���Q����,��!O�?!ʚ(��1c)��a&`B4��bDIp��@�qw�T�"a A��1p �U!"D*��"�h4�
I��GR1X\F%�)�q�h�P��!�a��Fha �d`�p���D��0	 H"�$�$H$@�! "�R*�`���RX��H��b� �6 �"\����afB�`JbD��G�Pŉ\��G4b�0j���n;��r����w���j�S��x,
AHm:7�x�T�%[6�gB�H���Q)Ըj��m/j��l�VE �vs�FDm��l��v�nD���@[M���kr��Uȴ�TY��Z{L���i�8%wj�q�B�� ��k���K{pm*��=g,�W[���
��U�<͘ 1n��s�S0*�pgp'=�ؒ2I�F{X gZ���ܩdVۣb��z�[�q83�v������,�A^�gv�ӷ']H5<�]�5[���o�ʹ�ze���;mY�vN�Y���M�5�Ҋ���Z뵴��e��MF.�$�Fb�w[/g�y�e�:CSv�m]@%�l\�����r�gQm�V�V27=��%�.d5��s�y*���80e���v'�����]��Yٻq�r��"Nx{y�����j
���׭��[�xl7�s�Tkin�P��`Z��؉ٻD@[2DF�qQVV��G3*�m�F�v�V�{D!kg��:z�Dv�t���s��s�@�_;�?7d/gh)�^Uc�7\�Y�@o.��#weaⶓ�� ��]6uȣ��j�NpM�F��u�	e��n����u�d�U�@Um�!*��M�SR��y�lݰv� �`8$8kj�d�8ꕀ�r��p�p㫜��UNl6%�����U�뎲;������=�Գ�@�:`�1�[mt+]c�ٗiUs��-�� ^��ո�Vɸ�)�uPz�{k�����%����J�UmK�Zks����Iٌ�:6]<ʒ�mg}���֢Si�ph��t�;jfղ��dj�;��W⹱)�c��Uvk]kpcc�[�J'I�<n�|9^�0�x	5��b�خٯGr���q�6	�YtJ����qd�� Q.��\ܮ�Hn�Vݖ��\ �Z�S����Q�[�-�]�Wmn
����h�L��puV^v�:L#�H���.t`�>i���N�P�{`B嫍a$]c�z�nn�'\q55<'��Qb�͠��"�� A�BP���w|�Ɂ̧�]�m�dU�`���`���@�d��qp];�.^յ��=:�έ4���/��2��m�f�3YŮwq��AƟ�Ϝ�;�Ս>�L.�[GF��wrR�ok7�܏`un�`tR��F6�ֹ�;[iZ�U��d6�.ig�Ni�-�m�鹹!ۣ���M��G�X��凂6ѧ��r��]���\�I]h�a������'$%�4�����:z;t�g����A�p��ݞ�2Q�ʍ�+����?8qQ���Ϳ6�������W`r��=oR�*i��YYYkw�zW�w���\H����{C@i�{�U$v<�*��ĭZJ򋼽*�^���3O�(���5�/@����(L�o"��7���M���^�އԥԒ�	-�2��WY�J�Yww��{޼�>�)�\� �S��/Jh�9+h�<�	�Hk�y��H��Jݲ�sƳ��0�M�l:�ղ�C��,CxG&�˺� ��e4
�נ{��D��ƦH�RG��w����UT�uϫ�	�g�����^��ޯ��G�Y���(�nd1G�{��� q]�\�� ����9�g{�yyy�yxhNW9UϪ�Ͼ������נ_l��궵�L	�&F�{݀9k�*���@����7��.����-����b�I�mm۞.�r�^���.9��u���� 7b���n��{Z]n�"n^��_�b��%���@�۹�Uֽ�Z��k�/�vX���G���35�rO^�ٹ'o}����B8�6!��0
�j����LimV	�x��k���?{�ٹ'+v<��f%YwJ�řzs��}s'�^�=�n�WZ�}�\Ȕ�X��.����u��>�vI�xNK�:�נy���$ڣ��ᑊ`�9&D��h��O�(�ۅPa��W.]j;�K<����I7�c��}�ۚ]k�9u�@)ֽ�W����
G��3@�����r^�A�z��� ~�����2dq�8��9u�@)�^�ىt�k@��^���0�2��K0e�}��)(7/@�k@k��As���+�*�*�k�o7$��N�5��PV�U�2�n��_d� i�zN��n<�݊c�26ڊ7xI�sŮ�q�ԍ���S6g�EOny���q	���񶘚N=�mz.�����+k�=V���I��H�]]�	k�q]�9����ao��{��s#iI�|[��<VנU�@��^�oK&,�$���1��q]�9�������VpLrH�H�G�U�@�+���	�����9}�f�B ��b��Eb?z�Lɗ>��WS$շZ�%�떋�!Wk�v��/ZKi��ð�v��p���	��@��7���]˷0\k���	�9�J����ۣr�]��u�fû1�8�<:Ǘ��LC�g���p�ԉ��c�F#�Ɗ#����۶�F`��ϵ[�uƦ@�&��ɰʵٰ�&���G��pö���`��dw��o�S�n��ۃ�=��c�������{�Ѷ�xa6cu�Ҏ����i��*�M�F��GT�i�lfW9,�F��q��￞�S���mz^��oJ�2A����@)�^�������z.����P�1&�s��݀{��ʻ �k�*���~bp�i����*�^��޻�u���_r�����^����}�|���H�]��:נx��@��z��HK�&	F��0N��=C6�#���֜�gv��^�s���T,��9�S�z���
�נr�@���E8�O�#�<M�ݮU}\��W��+��>S�/@�}�נ�^��w�$��9 �z]n�.Z� J� �� �h�|;���X����	\���z%�'k�*�^���H�I�7�z �v�+�*������ǕN�ژv�s��=ug�0��akk���z;6^5u�yx�:8�6���̚���'�z]n�����s��K�;�Q����6�I�ǠUֽ�uzN��+k�<V���I��+�e�^�z ηz{�>+���\�y<_}��=^���=�lM���"s$��yzUr����uG/@k�ށ���@���EnA��#�9^�@r��.5� �vx�f<Йͽ"6Xʄ��L��5��bX1��IKxY��NYV�?}�u���"����~����.5� �vq���G;�17�=�������W�U�@����	�	țqG��]�O����URQvK��^��S��P��$�@�z��kܓ���nN p$��Q.�[��/>E���#ƚm18�
��@�}w�mށ���@��Q�P���}8�۱��w�����]�(v�\�8�K�ňm�
�)����{����~/���qW�>_��z ���O���w�{^�6�F,�s#q)�R��W��*�����zY1dQ)$x�1��zS����9�s�5� ����wi�$�,��9�U��O������UI�r�FYp��)�@�z��k�9^�@���nI��PH�R���ˬc�ǆ�::pKW/;f��3'`�jGt���sv̵���1�w@���6mh�q;׌�ݵ��� ���j�+nu��͖��U�_��Z��ꆗ��:�GAj�,1�>9�g!��n
g&\ِܨ���'w:�v5�m.��|�î$���4����\�;uxm��m�.�lA���6�GA�Z�c\hr{YM�mvmOYff���*9��<7�I���jU��mr��á�uq���4ME�e0�a�mzn�OF��t��v������6.5����]�<ĩΙ��в��^]��O���W*�"�^��r��w�s��$vY&r�y�Wv�ڱ^^����[������z���w|�ī.�]س/C��Rw�)%�O��')K�^���2��e���*��e��6�@���Wn9~���zހ��TW�	9��1�X6���n����&�<n6�Lkݮgm�z:<F�:���I���r��r���w=�]Ěr22)$���[^���~*�ę;u�f䜾��rO���o�B�>���L�s"q�N8�
�U�����[^���IDc�##q���v�5����˰:��" cq!���=W��>�߳���vK�mހw���ub��jp�O[�8m�ʊ���ob�Yr�ݘ���^hmc��+k��\���6��������%�bX��wٴ�Kı=���&�X�%���}�ND�,K��3َ�V��\�.��7ı,N���r%�bX��{Yq,K��{�ͧ"X�%�����7�DL��,N��o3>5��Y��j�k6��bX�'���ț�bX�'s��m9Ɓ���9i��PĤ)N!�8���#�:��"�{���V���S��<������N닰<��� F!�	"E$!�"�q�  H��)����"�|������1�݊��ͅ :M��ز��Wg")�D��Q��� .(��`  ɡ�����MD�~�&�X�%���}�ND�,K޾�֋��u�k2fK5�dMı,K���6��bX�'���D�Kı;��iȖ%�b{=�dMı,K��[�5�Z˪f��LֳiȖ%�b{=�dMı,K�T#�}�i�%�bX�g�k"n%�bX��wٴ�Kİ{1��SFt��ܗK�nmC��չ�,ђ�x�[<�Ah��Tu�Xs��-�e����bX�'s��m9ı,Og}����%�bw=�fӑ,K��w�ț�bX�'�w~��Nh�5���Z�m9ı,Og}����%�bw=�fӑ,K��w�ț�bX�'s���ND��D@�&�X��L���֋5��asW5�7ı,Og��ٴ�Kı=���&�X�%����fӑ,K��w�ț�bX�'}���rfkT��s.K�ͧ"X�%��ﵑ7ı,N��{6��bX�'���D�K��xF0�"X5�����U�e>?
&�D������Kİo�d��][�L̹.��7ı,N��{6��bX�ʠ$~׾�D�Kı;�{��r%�bX���Yq,��ow��W}4�Ku�\���v�]C� J�۬� ��`��r���a�&U�e$��5�.k[ND�,K��k"n%�bX����m9ı,Og}����%�bw=�fӑ,K����5����kZ̙��ֲ&�X�%���}�NC��R����'�}�����%�b^�}���"X�%���{*n%�bY������5B�UY���{��7���ﵑ7ı,K������bX�'��쩸�%�b{?wٴ�Kĳ����gS�[�$Z�������d���kiȖ%�b{;�ʛ�bX�'��}�ND�,��@���������{��7��������y��[���Ȗ%�b{;�ʛ�bX�'��}�ND�,K��k"n%�bX��ﵴ�Kı?�t�#05�I㿫�gx�^}��vb��k����N�3��W��7]���k=�Hgu��ŷ���6՞�нvK�Vp�x�v[�ӌ�݉e�	�,i��-���b9��&u�uƬ��8�>�'a�[�{n��]*�d+nN�s�e�+g$�0s��:C�9��zuA��g�҄�=V�q�N�3�X:-��f�6�n�f¶Ws������~��{���ϝl����N�Ӟ����m\K���=T;gME�=�ec\haݬ��Q��ə��|��{��7������r%�bX���Yq,K��{�ͧ"X�%���{*n%�bX��o���'�r��w���oq��^�Yp� �L�b{>�ٴ�Kı>�g�Sq,K��{�ͧ"X�%�}�zuu�32��D�Kı;��iȖ%�b{;�ʛ�bX�'s��m9ı,Og}����%�b~?zo3<k+l։sV�Y��Kı=��eMı,K���6��bX�'���D�K��P����f����{��7�������X�\e���X�%���}�ND�,K��k"n%�bX��wٴ�Kı=��eMı,Kߵ�zB[�j�d�2i�v��ۦ	��w<�<��t����U��t=V�,aZ��U6i�����{��7����w��Kı;��iȖ%�b{;�ʛ�bX�'s��m9ı,K�{SSZ�k4ff��3Z�D�Kı;��i�x����w"X��g�Sq,K��;�iȖ%�b{;�dM?b?b?b?g����&"Lh�qG���,K��w�ț�bX�'s��m9ı,Og}����%�bw=�f��{��7������n+�Nd̳�n%�bX��wٴ�Kı=���&�X�%���}�ND�,K��k#�7���{���}���y�G*9g�D�,K��k"n%�bX|�}���m?D�,K���ț�bX�'s��m9ı,N�{Km�I5����V�d.�tcH��G,�0v<�t�ŵał�y������*8�{�oq�������ͧ"X�%��ﵑ7ı,N���r%�bX���Yq,K��������6⠧��{��7���}����%�bw=�fӑ,K��w�ț�bX�'s��m9�2�Oq���������R�q�w����d�=�{��r%�bX���Yq,x�;�	?����
ḛ���fӑ,K��>�Yq,K������aZ��R٧��{��7����k"n%�bX��wٴ�Kı=���&�X�%���}�ND�,K�>����7Er�S��7���{����wٴ�Kİ�AR?kﵑ9ı,Og��6��bX�'���D�K��{�ݻo���*=z�M�Nz������f��m�e�j]0���:��{pZz5f�3VkZͧ"X�%�����7ı,N���r%�bX��{Yq,K��{�ͧ"X�%��=3�P�h��L�Y������%�bw=�fӑ,K��{�ț�bX�'s��m9ı,Og�����*��2%�ߵ>>ӓ3Z�nd̹35�ND�,K���dMı,K���6��bX�'���D�Kı;��iȖ%�`�w$��]]aL̹.��7ı,N���r%�bX��{Yq,K��{�ͧ"X�Q0x(�����7ı,N��y�|kVL։���u��r%�bX��{Yq,K�� �P�����6��bX�'�k"n%�bX��wٴ�Kİgf3�cKv�݅�r�Y4RM����nܪa�	�˘�s	�7�����QS��7���{�N���r%�bX��{Yq,K��{�ͧ"X�%�����7ı������aZ��TVi�����{��=���&�X�%���}�ND�,K��]&�X�%���}�ND�?�������kS�n�Z����X�%��}��ND�,K��]&�X�%���}�ND�,K��k"n!���������UљE�Ʃ�����İ}���n%�bX��wٴ�Kı=���&�X�� �2'���fӑ,K��'�>����5r��-�kWI��%�bw=�fӑ,K�� ?kﵑ9ı,Og��6��bX��޺Mı,KB���~���=K�p�gb�wqH��&@MOnw-�:�!nn+�3�ܖ\�Pi�S���Y�xS�nKi���u\nWk�ey��S�`��b�Y�ی�J���Wϫh�geHΤ-o9ڻ�r��t��Ue�q�.b(M�Z�뭠2���`Ν��r�;��I?�>c�ύ۰gC���l����ƺ�ۓ�M�7���I�Giq���I2��u.e.�!���3G�4ga��'<Z�q�Ҳ2K�oc�q`⤱n]���\g��]�aTr����,K�ߵ�7ı,N���r%�bX>�z�?� Rr&D�,Og��6��bX�s��>�]k0�f\�Zț�bX�'s��m9ı,g�t��bX�'s��m9ı,Og������(9S"X���y�~5�&f���e��fӑ3*dL�?kﮓ���3*dK��[ND̯�D֪}���D�*dLʙ�k�fm92�D̩�_rf�3�	�����{��S��p�����3*dLʞ׽���Tș�2'���3iș�2&ek޺Nr�D̩������j��e�M�����{��Z�׽���Tș�2� ����fm?D̩�3(����Nr�D̩�.{��m92�Ḍ�I
y�Ը\՚��@#�1�ڠ�C�[�I�|�U#��.ٹXj֧t�U�Z����=��)�w��~�3iș�2&ek޺Nr�D̩�.{��l?���L��S�}��'9S"f�{�����Uѳ8k1�_����S�Ḍ�{�I�S��5�jhv�.�dK�߳[ND̩�3*{^��'9S"fTȞֻ�ͧ"fTș�=��~�uZ��5����;ܧ��.{��m92�D̩�{�Ȝ�L��*0֪j'�׾��r&eL��G�{맿?s��{�����|﷜�#
��u��Lʙ2���k"s�2&eL��k���r&eL��G�ﮓ���3*dK����ӑ3*dL�=��$�5u��d�̗ZȜ�L��S"wZ�6���S"fQ����*dLʙ���ӑ3*dLʞ�}���Tș�2'�oͰ��؄��Wp��PLZx����X#�ɞ�v��C���o}�����*|�l�Ak3��&eL��G�{��*dLʙ���ӑ3*dLʞ�}���Tș�2'���3iș�2&eN���F��R��L�e�]'9S"fTȗ=�f����S"fT���dNr�D̩�=�wٛND̩�3(�]��s�2&eL�{�r��Z��M�����{��S�����'9S"fTȝֻ�ͧ"fV��!А �� �"��H�#�B1� @�R
�X&)bH�$@�!0�B$�Ĉ�l� ��C"o�����s�2&eL�_����=ߛܧ���=��߶�;��n��ֵ�9ʙ2�D���fm92�Ḍ�w�I�Tș�2%�w٭�"fT��
Z�����'9S"fTș���������*���{��;ܧ>�}t��L��S"\�}��r&eL��S�ﵑ9ʙ2�D���fm92��r��}���*�kmV㢜`�Mssi�W�]#��v�B��vWC�:8�����%�[��c�9�����{��;�?�߳[ND̩�3*{]��'9S"fTȝֻ�ͧ"fTș�}���9ʙ2����M�?1��i�N9����6�c��S�ﵑ9��Mj�D���6���S"fQ�^��9ʙ2�D����o����{��S������tR�r�)��Tș�2'u��3iș�2&ek��Mı�D�Dȗ���[ND�,K���ț�bX�'��{3/�j�fDֵ�Z�ND�,�Q d�ﮓq,Kľ��kiȖ%�b{;�dMı,
�(�"'�5���{����oq���ߙ���b�|�bX�%��m9ı,Owٸ��bX�'}���9ı,g}t��oq��������9�gv��&�x䛝����jd��G;v5��\�LܯEj�0
Ti��_=ߛ�oq���}�����ŉbX�����Kİ}���(��2%�b_wﵴ�Kı/��Z����F�F��fj&�X�%����ӑ,K��w�I��%�b^�����Kı=�f�n%�bX����jkF�պ34]]k5v��bX����Mı,K������bX�'���Mı,K��}v��bX�'�z禡�ѫm˫�浫��Kρ=���ӑ,K���f�n%�bX�����K��Qd�ﮓq,K���M�iə5us0�2fk[ND�,K��n&�X�%��+��ĐI�}��$�O���lI�?�TW��TW��D�ʈ*+TAQ_�QE�D��D�� � �B!P	 D�B(A��B"��QH����
���D��TW�TV����DAQ_�E�E�D��TW�DAQ_�QE(��������)���3,�8( ���0�G�          `�:  �:  (  ��   	%$�*�%J
"�JJ*�UP�$@R$@  P � P) 	 $(R�*�   H  	�c`�4��Y������s����=ܵ}� .�^����-���:�������@W�zn{�^�>]�   =}`  ^�� �1JP-`PQ�AJJ  ���S����3J �(( T  EA) 1P��F 
Sn��s@� Q� �   ��4�AD �: �h n`  }�n�;� ��3�]��ϟc�ұ4;�J�������:wg/}�}�T� w�
  �Q��P� �D�{����{�}����G�x '�f{����}/n{9W� ������m��u���n����;�ۀ \�m�y���;v�q���y�����Ҭ��W��篶_|��mť<�R� 
 � 0�lp���  7�    gy��� �8���9����oz�A� }�'�Ϡ�0��s�{;��F�����>���}��ݻ}����������V�=�]��;3��{_m���L���H ��(��!�6��Yo�{��;*��z��w�|�8 ��Cz���G��� �g#��>�>�}J޷��6� /�ǝ;9u� ��=�'��=���ۗ�\�{]�x��z
>�ﾓx�v���ܗ�{=y�o��� iꌙ�)S@  "��d����@���R����   "{RM�EPd21��*{JT @DI6��A  �LJ��%�~~�����ڻ�k�M�����AQ^�����*+���*�D���*+�eTV*� ��'��	��0���-��I�2_^��3'����2�'��
�!�ňQÇ
cV��R�:��-�i���d�O|�/��B�/�?���q��@��d��%���Cԋb0�BQ�������M�+Je��x����$�>b~�!�9
��af)��0�U�<��!�s�ꧏ<?H0)�	�|���1�k"R$}D�0�����������	%2B\���� �(�0!�h:<!_�_48p�.v~4^r���u5�D��xÇ��?�%e
�mIC��x0�Bi��;�<���Oi湗N����R5Z�&��K��˦�$S"D��Yp��d�˾q��d¦@�q�rJ��P�6�,���<��O���K|�Ņ%�d��xR�xd'�h�X4��ՖL��`����8��4�I`@���?"q�>����i��|���\#ia9ÒR�:Ns9�8�L�a��
�p<I%0ׁ)��H�#��MOHI!���OP% HaB��y'ԉ�C�p�"P��3X���c	��R�ajY�l$4����<��
Db�'���iB~��$���8A)	
{LO9dΐQx�Z_ߩ��ǐS��#�l����0<�T\��ȍL?@�	̚ O}�bbB$���q�A8�w����!P�e��	S���CM�r��s��#L$��N0#,I�?T`�q}#�A�J-A�ǉ��ѐ�!�
$0��)�"Q1ׁF	ii`��aT
����C8RB��!���P a��$H�hXbD�҆���F�rGr2��<?�����̔2x�S��.I��&�	0�/3��a48c	F�G�,$@��e	�bH:qH�3g9������!����H��4��#]	S�ntC��!H~�D�5S�:E�@�-�а��\S�$JW�����rԕ$a�1$c ׂD����H4(`$�)�Re4x��H�E�I��bF$aB5��p!�&�F����9a�7f.b\9��#ʶa�S^ ��rF0$�(:� Bsy%� �	�k��i�@�--�)�t�q���XԂH�����ф��禅��=Gōxr�8��"$�2G�#I�dh�HBD���BJ�$���@ ���3���sI��osBHg�{L6@ڐ�~$�	�ji�0FDm�����]?W�_7���8�F�<9)��a$�N�&Q/����_m&o\巛���%p��?~�`a�9��%�ľ���|��#}t��B�$<<SИ����) x�)p�dC�(lK@*N,F$X1�rr��V�HH�@��!�Y0ћduy�"F�C`��2��H�3��dHP44y��7"l6�$$�&�E�JX�F���i,�k#$Y%��)0���ld������F-���O	m�&�Ҳ�mѲH�k�$V�(B�F��F&��$�0��$��ܰ����m��=d��?^�����!aoh�[�z�(���Q�]"�u��5ӗ��/���}c=>Mʕ�F�fx�t_�
~����y�z�=�x�iWXk�W^fr�ض�/�|��p�ܥj��׌�CTVc�U��}X����崈e���y��|i���"��a�� wZ�v�<*�+��T"���b���藲�xƭk����u����δ���vV�+ļ{Ζ����8|l����w4-�����^e��6��}UV��Z�+���/ޯɴE�_�,�M���5E�WBT��꬧�*ͫ�}�w��N{��~��g�$pT�N,�C!d�����XT%�� B�"5��$lj_��üFO�}�H�W9�G|��Q�	!K�hB�c�&�X�c
!"t�\&ְ��ڱ"8�h0�@�F�A*a̅��"A����1��KP�-L�,-���k���r�@� �u��H�HB{���Ǵ2kx�x�$8�II͵�����<L?SI$�����q<V�^$.[u�����~@�0hF
DH�P� F�
�h�"E�� �b$$c#��b� ��0)�"�*�2C @���BM+�"����8E�h��䎐*:�"E��ŀ�R�U ��H�T*
@�bXRX�"?�������A�d�1k�Sf��8����i���p������H�0�g0��<�;q�{؟j�������a�p���eaHV%0��T��(�@�J�� �"h�B�@��H�D��P��A�E� "�R-tB\��y����CHA�����n�����~��,��*��Z��ۛ���V����%%Jy?r�D8�BK��Ё �R5p�@��$H4��\B�iLH�C�G�o�_5��X�H��-q  �D"��1�q�Ub�%$F15V5��@"Ձ@"С��B�?sӞ_�#,���H4B\B�Z� �P A�V@�X�T�C���y�?�� ���g���^~�9����!�ǁ��e��y�(�i�0���i"��q��I	s����R�.����8J�i�`�S4�	`�&�I\H�0`�8��
�$B�hh��#@�уG�P��BN#��G*E׏�\���%�8N[�-����Ό����(ǛF$�Oj�G���n��sܾ�0��f����!������K���a�Ȱ�r#fjJlu�jJd���Ćl	7	L6D���WB5#qeP�7�CH���\ro��ݓ��+�+�jB�@i���hI��r�9����ӄ�Ӑ)�2�k�cF`P�`�XA�� �-�A��B�!�A ��B��bBAK`��R�bp`�00#b�N\	��R�:�8F�h"A8�(`h���*F:�����q���ӏ�@��fP�����t�Ǉ�@�l�xSGS�4G��pt�P15��
��@�@�cd�+M�h`:�a#D(bh ��,�,�`Z`i��i���F�l!!8o�.i�#CD8�(�
a�'�@(b�H�)/,�LM9��/��N&�A��{��}#��       � m�  ��        u��:��,�
�$���;>��˳��,b���UmQ-!O*�P/ET-6���z��k�P*�͆8t*�Q�P@    6���`  �E�v�!��Z8l�m�n�F�m%��  �     ���m�0�m�֤z�k2�� -��` m�Ŵ6ض�m���   �a#Z�   p    � 9�� %�m���m�������]v�ç=�h�%��`�  �k��   �ll  aw[vmqu�� 8H� m�   m��� H	 �����  �l.�8   햆��\�9�	 ��m�      �)����,�i:�H   �`l ���h�m  .�ۀm�h  �K�l-�=&a֕��j�'`-��T6�_5Ut�uA�	��H��}����H騛k��K-�V׍�hzN�n��Rq�;v@�7`�7P��R��1��[���M�p�[Vr�ˢ;%�Ⱦ��8t�<����AU����@S,�sڧ�Y\1�nRZ��)i1$Z��	3(@�F8'ʽ<�$�/dz{%���#�� Z�84V�:E�AZ۰�朠)4�n��ԺH��m6�;mo]!m  �RA%Y� a�	f�+*�
�<��<�h��%�G,�N�V�F�G		�k�@#�r�:�` ��m6톊�P�1�!� [Rp����9�v��a ��m�*���WJ���خ���`5PP*�E������@ l�`��+m�'N�)U\�K��4 VҖ�+�\9j������-�-$m&n�[   ��r�  m�m& 8�m� -�$d��l΀6�շmSf�l�d�A�1��d�ﾶ��m���m &���R!��Z�jW4��)%����r  [r�6�M`�@�d�Phh��$ K��i��l�'Iѹ6� �K���f�-�k ��avX�s���*�n�m�[� i!� �8 �[m��mねc����� �UJ�UO�B�.]�	TZ
Z��j��m�l�dY;K#UAí���)�UP I��9t��� �(�[A��� *Լ��+�=�l���m�ڶ<�VK� �� ��h$Jm��M��$����   �B@H�����u��YeA��W���Y]�� �m�`r)� sm�-ĩ2��i�N � ��V���Uʀ��e�jT�V�vW��eX *�U��!]fzB�OT ��� ��knd>R���U��yJ^vUm��-��RK�`�I� ��B`�2:�U���ϟـ r�(�� mpl[F�l��UԨf���(��5U*hِ�n���`�.p08p  m�
���UVT��SMr�˲��&P6j2-&D
8n�kȡÀ ��-��]��:iX���omXçF̪�L۷5l k�` Y`�(�z�m�kd�    [o3 ��]�:�8�M4UtZ ��		7ju�m�+bzXڐ�l`�6���Ni��J�%  m��sm�[d�� � [`��( �`�m���p�,����v�T�*��U��2�f���`#��X��ZU��gE*�*שVSi�n��mV��!v��M����4�Zhj�#a���,���o��(��
��M>�Vk0F�z,�d�-�� ��L��f_(
�U@&"���)^�V��lM�R%�U�v���XIC�U��-K��WC�S^�����9��Z�.-%H@!�pHk;P%�u�F$��7f���B��Iݭ�/f՛q �A�sPSr�*F@؀�Z��@UU++J�+P�RY����� �ؖQ"Aa��fX�C���B� �ڪ���y�Un�mT���_���
�9ʜ�?:�U�!|_��M�	 6�ˎ6�   �7[t�ѵI� mm��    -� �[��m���`	6�&m�   l �Y. ��j�<�9��檺�WjT����� [F���Z �mp �K&��GLݣ)6S�KT������4s�˲�K��N�&NW����U���3�m�
�@l[Kl�D�����$ m*�[[m��:�;
�;vrN�v"�w=!+��K�v�+q�WWf�;&Ԣ��v�T�A��j����5�m�8 ������ Iq����l� �oml�6�v��-�m�� $��     2 �` @��Hl6�	mm���[#�6��ѫM�n�xݶh �-��  �Rh���5�Ujc6ؐ�  ���-�����`86�� ö�6�  �`    �	�8[yËiW��/]�Z�-pQ�Sn�n��`H$� #l���� H��cm���e�v���-�BKhm� � 8kYa�lp�nh8$^��S5��m��G���Y�  ���  �$$H�w\2k#m����J�UP�v.z��Çmm��m�m�8��e�K��ޡ�5���r%���n�t�N� �D�ʨ!@ �5�v��&�m�#m ��6Ͱ��l8?V��� � �Am@  � ��m�   ��    �       6ؐ�$ �$h    ��m-� � 	    �� H$    [@ � p       @� p      ms��imt���*QJ�n � -����*����Tʷ!=	 ��bC��	-��i$���H m�@ k�o���	�m��[@�/ZHkm& -��ZlH ��v 6� $ :k�ZXa��[M�� ��� �� � [x9m$m��`� $ ���l ���H/[��Ŋ�UYz0�]l��@�[v���۶ �	��( x� ��6�  �� �� m�m�ObG  �͖)mm����� $�p $     �a�     H� *j�m6��t�m]m5��
Kyr����Kh $p    �l  8  ���|       l    $   -��u� ��'��)�+��x�f�� � [@m�    �l*����/�I�
��[VQ6�keZT7��6����Z�"V�
�j-�   �� ��6����6� �N� >��6� �      �     [wZ��    Hh     �          �`  	         l 6��   m h 8-� � h �� m���s�m��t���T������Ar��'g4Y��Q��R��u��dm�m����h^���n��[4P �H   m�� ��A�@[V��� H�m�p  �-��I���۳m$6Z�6Ă�[@ ����h�   �[@�p[A���b��8UU���h
���eZ�K�t�P  � � ͷ`   H   �����H    ��Me�ͩ�lH[�
���5�` m$��]�bސض�6xI�����S`v�Hn��^Hkm�6������D�*�WWG��������k�a��kY&�n�M�[F�m��6��b�XUz�
����Qf�l  e�������5��8l�� B]pm� �oN�BE�5���f� �k֜q�m�	   �Zj�H  I�Ѷ�v�� �:Xe���s-�k� �U#[�$�-��z5�q&�c`6�:o�� �h$iMn �ݖ��ԗR�m�k5����'_^�m,需�L�3�VP�����v�k�7QH֧4��2�y�ۥ����0��h63�:I��ރdTշ�R��Uʴjo  q h�gN�n���/YH���� /:*���6���VI�5u;6��p6
zꯉq?+��\�4 [/mJT3�l���� (���0T�C�ȯ����p�
!��#���^���_��j(h��0@=�8���_�
%�<X, ǟ���� ! �R��}���A��D�c�"2� BA�^�UC� � @H�|���] 0C��TD�QUT4AY��@:��tO8�A<!��`��T.( ���"�bz�rztOA��(��B"�Ј! ���=�
�Q�#��j��' ?*
�(R�}j��T? V�����?��<|C����x���⯨���Ԓ+�Ob�P=U�ꆏEG�b�8�������E���ECJ)
 ?��?z�'���/���
�����t�*T <���t��P�4PL�j�ǂ��T

'�P��?�AS� ��"u�S��������DA�� d�� @��o�z[@��Z  �,�;��ǳ�la�\�CUTQk�M.�� ���ӑ�k����t ��(m�O[�kp���h����P ��k�@ gUt��஬����8�x�:6�n������ey�b��c�Շ.eARr�6�U���G�x��4�)r���r��nۣ��lF�ʜ�հ�
��a�\�5<CA�C�H�S�[�W�����B�z�ڴ��ɐ���U������\Z^Ɯ�H6�Gf�l"���+u@٘J��3E �zJd�[r$��&�MC�+pU�j�ٶy��/��c��A�n�x_c�,;�Mzh��ݧN�5�q�H5�����5�j���:���=�A��L)c�m�l���Ȝ���@R�8�z�UV�mY����j�i,9�m���v�vyK#�ŝ��@�V�\j�U��M�T�z��n�V�S�(�V[U+e$��]J05�S	���h��8x$[���h�wlݛnn[�j�]U�������v<۲��{#<IK���E��]���mh]�͛��郪�I,g�m�lM��-�yݹQ.�T��	�+��ܶ�)�:�H2��Z᰽z��5�Z����C�8m��X*�B�n�Q�	�e�pm2�R���2ݱ�*j�%vf��-������+�`-bx�u]��RN=nCn�4��5U@UG;p`��K��*�h]6�$$-�i�ݧM���m�m�'��l�%�m�F���I�8�a� ����	 ��i*ԪT���uU@K����ՠ9��VŰ-��
vTp<�8Y����:�|�n� ��eT١�i�h�K&��t�t�ц��v��un�Bخ�g��ӡ[E]v����kn�8�l��8��t��N�+�[8� �\��U����țh����;��.㳶a���չ�����O@��C���05 ���+��*tQ�_?o��6]�n[.Y2뛅�t�^�^V�4��{���k��Wn��]���7a���a'8��b�vu��i-��/�m�s�]t���OJtf��ļ���<v�`��H�Z�WO[��y�Z�gh��EF�*Yhƌ�1�jW��v�\Fpu�gZ3Ӣ��@���U$�f�@���G�m��l��ڄ�n�p���7M.]��A�7���d�S2�����>�N@{+�Ƞ�{*y���y9x9���TW��.��[�.�I$��wi$~~�-$����_�$����-��G�M�%�I{3�|��$~`��6���]��}��?$��e�i$�S1m%I��i�Ԋ~��G�j��K���_�$��e�i$��5_���ۏ�:t1L��_ ����<����xN[m���s|����(����� ��~������Ew��������Y��~��F=�-$�����~I,C�]���猊��r+��9���R�76�d��4�؝ �պ�9W�&�%IMi�+I$�ٮ~��F=�-$�����~I,׷J�I~�6���	G$��~��Fg{w�(&���EQ�����y�I{^�+I$�3\��$��Bv��I�7I8�����W��%���ZI%�����$c�R�H�X�kI�Iqē�`c�el%�7��wy@]�J��~Ŵ�#rA&��`��,��覆�K�7d��=�2�	+��$�^n\i��y�5�	���3��y��ۖ�#�&�El5\�\k�c�iJ/�o����|vL��&V ot���\6�m�i��� ݓ+ �ɕ��-���W�}�����G�m.�(')� �iM9$���p�~�����	��*�X+�
*a 4QR��w��'���۔��F��H���ٚ�����vL�vL��Ĥ]���n������vL�vL� �����|���)ϥ�0��І��ۼ��5ֻce�萺�Ϋ�b�@o5���nm�����N&�RD��N/�fw]X�mՀwtO ��/ ۮ�+��M6�n�oL� ���]/ ݓ+ +j}�)*���]�f wtO �R^	"��3v��gJˆ.&��!&�V�i��K�7d��7���Q�q]���b/�~�,p��H�E"���q�`{۷X�p�މ��K�7��%����n;���n��w5\��n����G���a��v!6����|z>M��3Y�+�x����@^u�jJ#�Ǵ�ݥ95�E$��%X{5���K�7ze`ޙY]��",�av�CmӶ��=����e`ޙX�����P���$�I��V_}_U*P�3wʀ�{J�2��h_q�,y��dRGr6���n������y@]�@d.(�I
"��>�RJ٧G^���id�u�m�����;'�����=�d��gD�hk�tYk����.�����>�l��.����d��ΐͲ<��]�6��2�������F�V+3��f����,�Ai(�]��B�[��P�\v�h���z��e������'�+ �Ʒ2�;mmT�G������%cֲV���@[-�U�Kڸݻ{��ǣ{hx𒻫���,]��Id�YH�s��Ӌ�(�ن|����_�Jm� �Dp�����{��ݓ+*��z8`�:�K��&�Lm��o)/ ݓ+ ގ��< ��v�nӶ�I�Ӽw�V�0��x��V܉�I�i�4���=�2���x�H�
���{6��̠z�5�E$�F� ��٠=}���*׎��%
9����%ٺ��;;6��n^���(M.m��Wc�+۵^r%F��^�6�Ye��8���~�w�V�镀��=["��$�I#i8�{6���QUU]U
��(HQAǾ�@�{4�w�/���w>hl�H�Fܕ`n�Ҡ�}����w�� ,Wƺ�i6˵j۬ ���$X�L��L���Y	e	4ؒbm<����	(B��|��iP�>M����RH�Ё*H�)ҍ�u(�[2�<����ᡒ�����[+n��}IҤ�����i�vL�zL� ��o �����(�ݦ��bi]�X��V n��]/ ݓ+ ݠ]rյn(��ě��{٤�=�uY�U�|��D�!��(����͝u`f�����k,m�rIC�����2���n�2��-e�cm�m�v���e`�� ��e`�K�6κ�U.��bCi.Ξ�����%j�\k6uZs�J�u�kiU����[W�v��m4�i&� ����7zX�t�vL� ڗ�JU�M��%m�����=����e`ޙW��}�ԑ�A�p�&�m�i��b�� ݓ+ ����7zX�j�L���������>J*�����$��߸rI����9&�=�Tu:+F����x�4���4ؚWm���@jQ�����{��T�����!pkM��8u��t����nF��S�c�����ٮ�s�)	%T��|�n�2�^�X�X��V��+��t�3vf��ݚrI�����	TD���VoN,{4��=����jD۴�J�;�7d��7�� n���� �EDWv�i��u�oG
 ��&���|����w�� Z|+6�7$h��f����6ws�fnҠ/���Q	LBI�t�ۂ֎���-�һ;�����r�\Zs"��E�ܲ>օ3�ָ�u4������94�Ʒ�x���+��nޅb�u���K���&ܒ6Y�v\6M�ŭ�	�:݂D��2��v�]���Z��k=���:l�]Ƣ���]��Q��k�y	���[%���lEnm�4c�H�{\���N�I�^ղ`��x��#������r(3��׳.�%�ڸ��D�sK���7��G�^��g0�i�%M���;���x�X�p�ރ����SN�V۶�i�x�t��,��d��o�$�!$i�4��v&�J��6G ��K?Ͼ��KV�;3�����#Z��jKv�h-� =�-�}"�7ze`J��2�w]���bmЛ���@j����������&��`~���W��������x��vk	��d�s7�H�u�]������i�4j*m�I�vL�vL� ��o =$x�Ȩ����M6�n��YU�=�%@"!��3$���w�I�#�7d���eHĬi6˵j۪ ��M|��BP�BAv�*�X�ÈK(I��hm�<odX�X�X��x�*]�-[�G"rG`{۷VW��gw����K�ۮ����+m��S�B4����:�sm�ˆ�5�n:pOl��䶤��6JN'�q����fw]Xfk���0�DDPmҠ3 2G�{ɞO&fz�� ;�'��<vL��B>�����yı,O���y2�37r��3v�ND�,K���x�D�,K�{�S�,h
�2 ��Lp"a4��b�� ����Ec�13SV����)�D���I���p�F$a�����
(XB��G}IA0`��CT @� $P��!��l�lhZT ���r\��	$�AbȤX� �#$Y"A�� [HBBE�1�StтX,BH`1�#�*�)#�B��"F@�`"�a �1���,@�F$�d @�2B$ �/�ؙ��&2�2�Bd�𢘥 ���H�	�	�
!J%#B	���K�UB���V'�JJ�T}<3$�+�y�f[0���$ F FEB�z����*`�UG��)�(�@��~�������O�=T���TI��%P��>���}��� �?DȖ%�{߶�ND�s����~�(���*�Z�{�7��g�X߾���Kı;�����UC�L�bX�����9�F@��QB*܉�����yı,�>��L�������(n�8jyı,N��xq<��$r&D��9߾۵<�c���/��x�D�,K߾��|��,K�T������lkzx��Lm��թ��:�GN� �nmZ\�]r7e�,���X>o�;KV2[�~Oc�@�DȖ%���sjr%�bXx�G?}����ı,{������"}���O"X�?�a�:l��?����ݹrl��ڜ�bX�%���o�?�5؛����59��D�Dȟ}���Ȗ%�b_�����Tc�H(�12%���3섹wv�n��n�<�bY�DFA��xjr%�bXx�G��ߎ'�?�"_�����K<TP dL��{����%�bX7���nݳ77fn|*"ng8jyĳ���=��O!�A�DȖ%��6�"X�%� ����}��?D�,
�����Q�(��^|�����S�<TPʙ���O���r��]��۹���%�bX���~�ڞD�,K
�����jqT�I��i�H�Yb{����A?R��$Ͱ��϶��aDq7��::m����jm˨���p��l�O31�����ș��wﳉ�Kİ�,{����,K�����?Dɉ"dK�~�ڜ�bX�'���3�f��ۛ�~B]�g��%�bX>�����ȕL��=���yı,K�~��(șı;����yı���wy����sSLҵ׻���o.	|?����䒄GH]!p�Ϸ���D��/��2b ���ﳉ�%�bX>������L�b_{'g�nI���.e����%�bX�Fg��sjyı,N�~�8�D��@dL��~�Ȗ%��Ȟ��߸~����oq�߼����;,�GY�=�7�ĳ��߾�'�,K���p��<��,K߾��'�,K�2&{��v�"X�%��{�_���p�fْe���+��˭� H]���K���k�GB�2i۵�9x��l4��S�[��c8֫��+r��ҫ�����ٺ�ۍ��h��xݒն�f���t�����lt-�v؜��j����<��;:Զ�j�tVQ�.����s�ힹ��Y�v�9�k���~��_�׫l��^V���FW	�p���3��%nӳ�xAۗ1��߽?6;����y67X�ѡ��(je��l�[�mV402¹�A���%�w7nn�z�D�,�2���ND�,K��}���?TȖ%�}��C��D�,	�=�{�q<�bX�%��?��̼׻���oq�ߟ��É�Kı/��n��ʙı=�{�q<�bX�����"X�%���x�_�IRS(7|�~ov�{��2_~�n��Kı=�{�q>S�L�bX>����bX(̉�߾�q<�oq���w���sӕb)�b=�7�T!�2%��{߳��Kİ}��5>�D�,K�߾�'�,K��-����ݩȖ%�b~���g�7.���ܓ3s��KϖA��xjr%�bX���}�O��S"X�%��br%�bX���8�D�,K�{{�Y��b��Jc���g�IO�R�h�:3\����:z�Ӕ�e�m�M3J�^�,Kľ~�w��Kı/��v'"X�%��?{��yı,}�ND�,K��{۞\�f]ݗ0���'�,KĿ��؜��E�*�B ��k�*�ș��w����%�bX=����bX�%���x�D�L���~����Y^�������bX���xq<�bX��{�S�,x�2&D����Ȗ%�b_}��ND�,K�?JvL�n]ݷwnn��<�bX�����"X�%�w��'�,KĿ���ND�,K��{�O"�oq����}
љ��׻��X�%�w��'�,Kľ���9ı,O}�|8�D�,K����"X�%���oK�͕�a�fS&�i�$Z�A�H�%���lQ�dm�n�	�������<n�	*Jf��{�7���{��?~����Kı/���x�D�,K����"X�%�|���Ȗ%�b|����T��j)�սߛ�oq��������Kİ}�xjr%�bX�����<�bX�%�{��,K���oK�<ٹwv���37x�D�,K��ND�,K����'�,j��������2%�����Kı/��w��Kı,��p�����������S�,K"�,K���x�D�,K��݉Ȗ%�b_߽��<�bX�{���bX�'�d�nywd��ݗ0���'�,KĽ�wbr%�bX|��}����ı,����"X�%�|���Ȗ%�bt��2L̚I��E�a73e�97JY�b#g���e���
�4ܬtm���Y^�V�|��{��2_߽��<�bX�{���bX�%��{�O"X�%�{����Kı/7���ܻ�n�����yı,��59�Fı,K����<�bX�%�����Kı/�����%�g����������̡]{�oq��K��{�O"X�%�{�ڜ�bX�%���x�D�,K���Ȗ%���ݱ���IDU05������,K�����Kı/�����%�bX?��ND�,��H �ʪȜ߾�x�D�,K����4�����w��S�,Kľ���Ȗ%�a��ND�,K��{�O"X�%�{�ڜ�bX�'������pd饷x�X��:s���D�:�Ϋ�b�&o-�%�sG���XJ�����O"X�%������Kı/����yı,N�{��,K�������~oq����o��q�n�)�V�S�,Kľ~�w��Kı;���ND�,K�~����%�bX=�xjr$�,K��{���&e��nm���'�,K��w��9ı,Os��8�D��	��{�S�,KĿ���Ȗ%�bw݄�;m&f����ww"r%�bX���q<�bX�{���bX�%���x�D�,K���D�Kı<��m�g\�wv������yı,��59ı,K����<�bX�'s�܉Ȗ%�b{�����%�bX���6\�f��.�q"K�Y�f�q����I�vݠ��I/B۷,�9�9��[u���{(������&̆��6lh�9�p�P6c*�Xx�ݓe�ڎ8�`����έ�%-]�`�{na�-������b�ڬl8l�jM����H�N���ߟ6d~`�9"����S�8$(6�e�L��cpnu�Z�U66]age�3o����w��>A��[tm>vy�g$m�]�Ÿ��vH飂�F{ss�����x,f�vnn���wMND�,K���oȖ%�bw;�Ȝ�bX�'��{��j ��,K���jr%�bX����%�ik��{��7���߻�9ı,O����Ȗ%�`���Ȗ%�b_?w���%�bX�;�G�p��S�h�|��{��7����~�Ȗ%�`��xjr%�bX�����<�bX�'s�܉Ȗ%�bx~�Ify�r�����378�D�,�BA��59ı,K��}�O"X�%���w"r%�`EA�'��{�O"X�{��7��<}۪�f����7���%�w��'�,K��w��9ı,Os��8�D�,K��ND�,��~~�߽��9x9�:n4�1�{v��M��dy�)�$�:8�5����!�j%��37x�D�,K���D�Kı/����yı,��59ı,K���x�D�,K�N�nv�L��ٙ���D�Kı=�}�q<�ʩ�DB(Qy�,��59ı,Os߾�'�,KĽ�wbr$E��ow����c���f~{�7�İ{����Kı/����<�c�2&D�}��ND�,K��ﳞ���7���w�����3Y�+��Kı/����<�bX�%�{��,K������yİ>����>�>�}H���y��t �d�773w��Kı/{�؜�bX�'����Ȗ%�`���Ȗ%�b_߻��yı,K���rH]6�.��"�A�[�[��:�&����6K��zt���!��{��ݸ��mvX�{���=�x�>������ı,O��p��Kı/����<�bX�%�{��,K���zB��s.�����nnq<�bX�{����G"dK�{����%�bX��݉Ȗ%�b~���8�G��7���~���ݺ��iZ���x�,K����'�,KĽ�wbr%�T��E�"lN�|�8�D�,K���Ȗ%�b~�N��t��we�ə���%�e%�{��,K�����q<�bX�{���bX�'����'�,KĿ��.v�L��ٙ�7wbr%�bX�����'�,K��{�S�,KĿ���Ȗ%�b^���9ı,O;;��mݣ���t&m�9���gX:˲u1Ѻ��Z�:$�N^i�2��F�}��O%�bvw�19ı,K����<�bX�%�{��,K��=�s��x��{��>�������̡]{�o%�b_��w��*�dKĽ�wbr%�bX���q<�bX�{�������oq���>���W+K\O"X�%�{����Kı?g�{�O"X�%������Kı/����<�bX�'N����-��7wM���,K������yı,��59ı,K��{�O"X���+v&��n��Kı?{߈g����ۛ�r[��O"X�%�����"X�%��%g����?D�,K��۱9ı,O����'�,KŽ��-s�+y4��i�d�u��J9��-��j�CWM �@�<[uQLҵ׻��ŉb_߻��yı,K��v'"X�%��?w���I�&D�,����"X�%��d���&�3.�˙s7N'�,KĽ�wbr 1ș��=���yı,����"X�%���{��w���oq�����/��k+j���bX�'����Ȗ%�`���Ȗ?�i"dO����Ȗ%�b_��v'"X�%���!�nu�&�ۻ����O"X�%�����"X�%����É�Kı/{�؜�bX�%����=ߛ�oq���L}�]9�ԩF�"X�%����É�Kİ��}�۱<�bX�%����O"X�%�����"X�%����S0�}�C��0����5a�,#!a��p0J4!�,�� �	�0 P�0��l�4J� ��R$U3P�烋�9�)�`H��H"B�E	�D�$X2�H�"���<3���R�b�# �� ��Bs>�aM�����`1X��� Bs�
``F@$"A�L`+a�,X(�=�g۶��7vivUZ��:�3�ݍ䞬h��;J)qae�[}h�E[RqON�H��D�8�CBۯ�k���qջY�^V�EQ$-��U��������n�5]*�0HF���8l� ���-�۝��+�Q�pV@}����+:���H�X�T�ug��nG��'��σ�So�:b+��z� k�.��mp�'��\ۦ݂�r�.z-DیJ���l���N7lv}SR��L�B�]�Z�8 4`3�˳ �`���a�9�I���:v��.vWhPF��*¬� �vTA��o]��J��F0PN�(��8�>u�(ݤ�lU�ε�i
^-�ݒۤ�5v���Қ����g86�'F��K,����U�=6M��73Q�5u�"�����0M��zmR�5 %:R��8,h�}�;Xv9�ɇ�m��;�::�y�.܌gd:��;�h�n�8��;�6�z�'�Pٓ��M�n�m�Hm0�!;LN�\�i�d�C�5�<nM�Vz��0I���Q��i�L�V�f��[VѾ���ä[%�F�w��yZ���HY)t�*��D�P�"AvүΛ���e�n�#cؽR�u�1[�cAg2� >nd*U(�z.1��uk��Y ������ u�68���F�Cm��#m��&�U���(��7@T"\��ݺ�sv��k[�K�gk�q* 3���t+m]F�j	�P�p��b���=���ETs���6�زc
� �j@HH6�6���Ƒ��j�9��kW=t���&N`:����V�:�n�@$ Hm���c����Z*��a������H�։]�Vj�:���m5{i�='l�lƹ�C�ݶ�3�j�K-R�OjuRn�(T�&-���ʔg������u]�yG\��Tpnz��к�(��Tv�σ�G�ە,�����U�:ۍ!�pr��I���^M�b;�1�b�]46Sp�\TL<@P���b����8~@�A�W�|�Q?
�6_�Iin��I�M�m��#v:�	\m�\��qʜ�Y6�;�Q��1�v{W1u���l�E.���m�O]zE�7���zctH�f�1�<�mѰ��zc��c���0�3�R�{s�h�@��6�]������9�(6���~n��4�^:���AA�j,��M�,��e	��qk��-umׯ�p�����A��h�l�׺7U��//��GDYD�{B%��8u����ftVˬ%a���3x�<v{���:�sR�7~����D�,K����,KĿ�{��yı,��4?�șı/�~�x�D7���{���? TFuS������%�b_߽��<��L+"dK��Ȗ%�b~��8�D�,K��݉Ȗ%�bx~�Hg����ۛ�d���yı,��59ı,K����<�bX�%�{��,Kľ������{��7�ߧ��:��iZ��"X�%�w��'�,KĽ�wbr%�bX��{��yı,��5,���#�GԽ���$��$bRK���bX�%�{��,K¤g�����%�bX=�xjr%�bX��{��yı,N��ܜٻwim�n���&��s����+���.N���J��^���2�e��ګ{�oq����~���|O"X�%�����"X�%�w�����"X�%��br%�bX���,��.Mݷwnn��<�bX�{���ʚ�-�QJ"|�q"X�%�>�x�D�,K��۱9ı,K���<��2%�~��.i�f����˺jr%�bX�߾�x�D�,K��݉Ȗ4��b_}�w��Kİ{����Kı?~���?]j��Y�����{��7������Kı/�����%�bX=�xjr%�`|�2&{��oȖ%�w������Ej)����7���{���{��yı,��59ı,K����<�bX�%�{��,Kϫى�z1!1T�*�BJT""c�gGM&�p6A��'J�'6�j���e����nn�<�bX�{���bX�%���x�D�,K��݉Ȗ%�b_}�w��Kı)=����&����Ͷ暜�bX�%���x�D�,K��݉Ȗ%�b_}�w��Kİ{����Kı?�owpݙs76[����yı,K��v'"X�%�}���'�,j)EtHdM���p��Kı/�}��yı,O���7Cq�6��ϩR>�}K3vZyı,��59ı,K���x�D�,��;���BE<���r���wm��www�H$���lE����w�ؖ%�bw��D�Kı/���x�D�,K�l��nR]��0����M R�Q�f�Z�e��m�5=�7�$2����3Z�+�w��7���{�?w���%�bX��s�9ı,K����'�,K��{�S�,K��!�r�rn����a�w7x�D�,K��r'"X�%���{���%�bX���ND�,K����'�,K���[.�i�$RF���gԏ�R>�{7���%�bX���ND�,K����'�,K��{��Ȗ%�bwޔe�ۛ��Y��Ȗ%��ȟO����Kı/�~�x�D�,K��r'"X��z�?�"w��Ӊ�Kı,��.�wnnnl�4��Kı/����yı,>�}�۱<�bX�'���'�,K���xbr%�bX����e�ٹB5�SM͓+�{ ܾ13�$t�gJ�$἗Y�z�?ݹ��=Y���-ə��'�%�b_��v'"X�%������yı,N���	"X�%�|���Ȗ%�b_�s;.annn��ٻ��,K�����q<�bX�'g{��,Kľ~�w��Kı/{�؜��2%��>�e.|˓wm�����Ȗ%�b}>��'"X�%�|���Ȗ?ș��۱9ı,O}��O"X�%�{��\�l��ݻ��t��Kı/����yı,K��v'"X�%������yİ>&D�}��'"X�%��!��_�:��ik��{��7����߶��Kİ�}_}��O�,K��}�ND�,K����'�,K���H�E�PA���D��;�o]��^�g#��
���Dma�zH q%���;Vi��nyvcj3�hx�u>�&�1��&�C`x��V�w���6���T�4V��v��X}�t�TX�a��{]�c����ҫ%��=��$��^�n��-�:���hL�nN�m:���-�T��c�Y*Ոi,�-
X�Zx�ˎ{\��7
;\Ы˔��Î6�q{�����1��H/���M�o[K���x�R:m����jx���_�q�>r"�г����o%����8�D�,K���Ȗ%�b_?w����	����K�����Ȝ�bX�'���?�ͳ.�������8�D�,K���� ���,K�߾�'�,K��>�r'"X�%������y�2�D�,�:fO�ۻ�7.�4��Kı/�~�x�D�,K���D�K�i"dO}��O"X�%������bX�'�����r\��-ə��O"X�|!"}�}��,K�������%�bX���ND�,�fD�~���yı,K��ϴ�e���30��Ȝ�bX�'���O"X�%��� ����ߌO�,KĽ����'�,K��w��9�q���~���o��f�Qr�V��Y���Z�m�\��l7��h`j��������-㙓wm�������%�bX�O��Ȗ%�b_��w��Kı;����_"dK��~�É�K�7x�����\�jD�}�7���{�K����<���]��,O��"r%�bX�}߼8�D�,K���ȟ����lK�6Ys��wt�ݹ�]���%�bX���jr%�bX����q<�c��2&D�}�ND�,K��}���%�bX�;7;732�f���ݹ��9ĳ����;߿�8�D�,K�p��Kı<���q<�bXș���S�,K������r�����,�Ӊ�Kı?N��'"X�%��`�{��8��X�%�{��jr%�bX��{�'�,K��w�m�~!˶�nQP�;��7<���"�vY�����oS���G��{�X�P�ݶ昞D�,K��}���%�bX���r'"X�%������|��"X�'��br%�bX�ӷ��rܻ�.[wN'�,K��w��9���ؖ'{���Ȗ%�bO����bX�'����O"|9S"X�gK/�Z]��ٙ�fi�,K��~�É�Kı;;���c���1��C	ȝ������%�bX����9ı,O?om3/\̛�l��ۚq<�bY�2'��19ı,O~��N'�,K��{�"r%�`�b}����Ȗ%�`��m?�3K�nn�ܗ3t��Kı?w���yı,>�{�xD�%�bX�����yı,Oӽ�Ȗ%�b~�N����xy㲆�	ޑ���N�k%���z(�[,�fM�c�t��*�v+|�~d�,K�{�"r%�bX��{��yı,Oӽ���"dK��﯋��R>�}H���\;m�7$R8��D�Kı/������b�DȖ'��br%�bX���>�O"X�%���9� ��,O����n�3wn��a-��'�,K��}�ND�,K�{��'�,~�Dȝ���'"X�%�{߾�'�,K��};�.��4�Pϻ���o��� ����8�D�,K￳�ND�,K���w��K��@N���*�?D�y��,KĽ?�ng�r��͙��Ӊ�Kı/��v'"X�%�3��{�O"X�%��w�19ı,O?w�O"X�������L��d��N���t��	c���mg���e�&�v��bW�����w;�/�w77ff���<�bX�%����O"X�%��w�19ı,O?w��	�&D�,K����,K�������\��l�7wwx�D�,K��xbr	��,O����Ȗ%�b^��؜�bX�%����ȟTȖ�����s5���>��oq����߾��yı,K�݉Ȗ?�4؛��oȖ%�bvp��Kı;��ne��m��wv噚q<�bY�"g{��ND�,K��~�'�,K��;���bX�'���'��7������������=�����X�%�~����%�bX|�����D�,K��}���%�bX��{��,K��4"@?~����v�ɗ�M���i�͑����#�gXb��0�(�n��s��:�;g,:�ö���p�W�c��HO'l[g�S��b��\74�n���},�dz��&s֐�o٠�.�4.��ق��Y��d��um"����Ƚ(�]��܊�::�hK 1֮�-�q�8;j���Ph�+��7[*	�y�����I��q�w�������ͮ��f0��՛�!���ێXh���k/*����Nh�������n�3wn��afn�'�Kı=���Ȗ%�by����yı,K�݁�șı/����yı,K>��񛙻��wm��'"X�%����g�|+��,K����!�L�bX�￿���Kı=�}��,���#�^�4z������~>�%�b_}��ND�,K�{�'�,�XdL������bX�'�}ϧȖ%�b_�essvfa����,K>BD�~����%�bX�Ͼ�Ȗ%�b~�y���%�`|��ș����,K��>��Ϝ�7v�rffi��%�bX��{��,K��#��}��~�bX�%�~݉Ȗ%�b{�{���%�bX=�'eû��<��N幃�i�l[��^�x(dg�71YY;	[9C�n�3Z�-s��Kı?w���yı,K�݉Ȗ%�b_}�w���L�bX�w]?�ϩR>�}^����NJ�D�-�8�D�,K��wbr�`�dL�b_}����%�bX�Ͼ�Ȗ%�by����yı,N��g33��n�wv'"X�%�~����%�bX��{��,Kľ~�w��Kı/��v'"X�%��}�<ݶf�����nn�<�bX�'�����Kı/����yı,K�݉Ȗ%�b_߽��<�bX�%��L3�m�ۛ�vۚbr%�bX�g��8�D�,K��wbr%�bX���{�O"X�%��w�19ı,N��g��6�&�.�zk-�7���$�׷\�6�:�$���)��ӯ|�e^�)6֏׻���ı/��v'"X�%�}���'�,K��=�ND�,K��{�O"X�%���Z]��ٗ&���ND�,K����'�,K��=�ND�,K��{�O"X�%�}���9�ʙ��>��ϛrn�-ɹ����%�bX�Ͼ�Ȗ%�b_��w��K(�$�J�H�����!		#5G ذ�"�Db�� �$A��DaF$H�IH�	!�,XH� 1�B,	F� �AH,a i�����Lɘ�)��$�"���T �U��A��la+��Pa`$Ï�D�Ez O {�x!�!�0�����h"�_JC�~yD<���z>�
�'"_��v'"X�%�w��'�,K��ݴ�\�i���w%��19ı,K����<�al���p�G�nɕ�z�b�)Wv���ID���n� �ݖ��ug|���,0�p9I��'�B�N�F�*�7Gbu�Z��+Bm�{v�î�k�ێS<ʼ,E=�fh1��.ۥ@��R�	{�foK�y��9"�FĜ���u`� n��w��
��J���m8ԉ'*�?{vX��,ﾪ����`fw]X�4C�4�m�nK ���.��w��$��=m� +P����lV��o 7z<w�V {dx��*YM�*����\iycfLU]<�q�Sf��#vC�vִN�'KO����wWhi��ޙX���G���ÿ��M���i7X���G����+ �j�
S�M�m��k �ɕ�m�E�n���={"�%o]�Yi*I6���X��X�L� �#�l� �H�Ě۶�J��X�L� �#�l� ;�x}]�QxXIҢ����u�s֦'U��;�i���/'\�-ӄ���6�n՘��Fܙ���<M���ӺM�7�)��z[r,PH\b� ݲx�q�u��k0�Z�]uX�·\Z�=�q=�mӡړ���|o��^��q6,����-���&-j)^��8L��v�!v.�,lj��8m�Nn.I��3m�u�n:WR{3
���o;D.��U9�sd�.鴻3\ɛd�5��M�J9�7d�t����ᣎ*�l]/"㛘܍ƤI9^���~��{6X�2�k�b�m�*�m��G�:<w�V�&V W�!wV�M���M�Ώ �镀vɕ���.��ʻCn������+ �+ =�< ��������M����M��&V {dx���=�۫s�͍����9$s��n�=#l5:�h�r�ۆ�lM��yV�ݞٺ-7I��N��#����+ �镀zW)e��$؛t�����}Q���/*^
Ǵ���X���Ux��M�i[��7ze`�2��#�t� +��]F'i�M[wv�`J��)�n��{�������Z��+N�I&� 6ۚ �74�t��t�Q��}껶ʴi:r�*j9����	�1t�.7]�	sڭ�뗣N�����efk�����.�Ҡ/1Ҡ���0��U�wWhm&��2��2�vG�:<�ú��C��bj�&�{����$����O���

��BD��d$�$���j�"�]������S=���ؓ� ݑ��G�nɕ�ot��=+��F%t�lM�o =�<vL��8`� x����i
�k�`�����aV9��3�-뮞�3rv&��f�4�m%CV�&ݶ�@�~�L��8`� 6txSnU�bn�M2�:�;d��� l��}��3;��k�D��M8�iG ��^ l���2��X�ڲ�.��i�Zm���#�7d��7�e`O�}_}�:���`yi�ͅ
)"��#q��e`�2�vG�����=�طK�c��^�t8M�D��1u#m���cpÌM��0�bMţ�+����)��7�e`�e`�G�nɕ�mY�te��M���I��Y�着��;zX��V{v�����;Q�m�&ڱ�X���7d��;d��7d��=�)V4Э�i��&��&V�&V�&V l��mԫ��	��V�I7�vɕ�nɕ�:< ����I����C~�̟f�mn"q������
���s���N�0n!c�y��n������v�V�g��G]�:A�^:��}w˗�<[�7^��P�����n�m���]�o]i�q2�f�0�ܜ��n��.��y�l��9*�e�U���m����[ю1u�q����W���3T&�wV�i�$=o��}�i.�i��]p��0�]��BB�i�������Ŀ1�ƽ�[/U��g�[��v�h��N�v�F'Νhn��#����'C)�9Vw�]X�6X��,fnV Cj��մ�bI+N��#��B��3vhoiPmҠ=�#�ȋvۺ�Ci7��<{�V�&V {�x��t&�WV�x�L�vL���, ݑ��m;��I��%v�`�e`��`���f�XU�Ew>�&(��4�n�{c�-� �9��D�GGM�4]���O�(��ICr���I+�[���ݖ�ݝ_~A��u`fo*.F�RD����I'���������A�$����w�ntX6�\whM��i��fh-��.ۥF\�s^��37g :�
[�V��$��x�L�ntX���l� �[V\��[M6$�Zu�m΋ 7z<o�,�&U�U}���X�)��a&��V�ݪn�D8��q�n�%�K����qzUWhM&�w��� �ɕ�z�E�zp�*㫺M6&��&����=�e`�"�ޏ 6�BAݦ��RM&�l�X��X]�f�G�m�E�J��t�iU�� �����n�,�vK�����TNQ��v������7ze`}�`�2�_H��J>X�LE[M�4ݢ��{L���R��
��d�
�#�<h���F^�Ԍ�D�M��v�`}�`�2�_H�ޙXоV���vؕ���=�]X�n��ͺ�<�5�RG*�IwR�9�iʰ<�����u`yfk�=�2�]q]T'm���&�X�*���@]�@ҡ%P��(U�������rI��v�^�i���7.�i�����+ �� �ɕ�w����ƻ	�s�����O��[�P�iٗ���E`�.��Ru����:h��d�k ����=}"�=�2�����K,�'I��[n�_H�oL��3]��f�_Wԑ�ʉ�0�G$iP&����V����+ =�; �-�\��㑷%�U}T����7����, ��xоV���vؕ���=�2�_H�������9$�i�k4x�� H�0���d$�a[6�_!��c�+ ��50�c#�f���
�+h�yP�KP��
�� ���$,	J��c���� ���n�`H������\��^�}��y0�/0i��[Je0�!��$�BE @�A�V �#���#` D��TP�(��X�>� �D �Dx2	�VE^���@�?_�[@���  �t�v��ݐ,��s��Y�UTQP�Cd8���Q��P�f�ͤ��p�m"�t�0=��^6
6<�0U�Q@�2��r��y�`*�Al��J��]մ8�	9�ݘ�Wa:Sp<KU���Ov�#,Q;�\f#�����;ۓ`Y�QcMt�,�2)k��:����+b�0<�݉�%�T�%qے	F(m��^@e为�p.p;Gi=[5Q�C� �x���l�e�W6��౜G;�	��tn��k`{;.ȭ�їa���Az����ts<�]r�p�ʛl
�ܷmq�l����*��k��J��8k6켽�P�b׊�݁�S��;�x{M�>�Uu��k�8���h�4;�p+[/B�'�����nZ��4ge���m�[R.1��S\O#����KcH�	�Qvk�#\#�ƴ��nW,1N�'Q�[o$+A�2۵T�[�R�j`#�	V�����Z;Q���+RV�;�5�uX�g<��ބ�u�s�`nR���eWWY�t�06��L�ǭq�nNId+�2�X�`6ݯY�u�r$�^8tNn����F�a��m�=��籠�9��R'R����V�,���pP�x K6Ic�08��j�ƀ���m'6��m�:�M�v�j땶��j[�#���vm�k)�q]��zV�4��l�g7Y�he�8�K�-R�챏b���3�@h/�v��j�֑m�`�]7`�Hm�m[U�����������ŶZڸ�:ڥێm�[@$6�h$�!���%�l[du]R�*�m��r��&j��0ͬ�j�Eճ��t��b�<nـ;b�|z�iV���M*Ի�uR,�)����WM/;�-�.�P�%.�/k]��nIz�`�Ӭ]�P*�'�V�Ŭ��v�,�۱�A�m��8��ٶ�mγ���ü7HЉ��4g�l�&��,2m�%�ݪz"#��C���Q�C����"~��TƂ'��ݖ뙙6۰�rAJ�L��ŵ�rvݛ�����4l2�;=\y�O\P���ǪMA����3�N����G�A��K��2*Bw;s���������Ig�������r�r��s�y���a��ݺsg�UӢ���[U���+�2n�0��p�-\pv<��J�Z��`Ipݠ�d�礉 i-��mХ]7Vx���q�g�mʗ=�{[m;qv;v���V닖��v��Zt�e�jt�-&�Y���V�`� =����镀MU
��Bvۺ�V�k =��ٮ���۫�ٮ���H�>HGJ�M[m�}���=�2�������%�M�j�i5�{ze`{�`��^Ȱ��BYe�JrF�I*���k�;�7��<�����u`��I�#�B&�JT�m�ճv��,4I��쵪Nš$��L�CJv�J[i��ݦ�^�X�dX��V�� vܫ�մ�m5m�&�vGτQ`mEJ&)�'T�=���;��k����ʹ���r�V�x����m� ��E��< �u܂���lV�V�`{"�={�`� ����=|B�mU�wWi���={�`�G�{ze`�l�?f�Z��R!�"�I��K�5ط�6�	<4��:g:�Ჶ�˫eP�6�f�շm��ޏ ����oG�ﾪ���o;����I*I��q�����ޏ ��E�z���:�AZ�b-:M���u�ޏ ��E��ﾯ�����f�Kٽu`~��E�ڑ���NK���o; ���f�X�u�mԫ��&�i�������镀�<׽'E���%wV�qԔAqq�ʘve��l�6�:�$����~|�t�iFڄU�A������ ޑ���zG���WV�M�*�i� oH�^�X�#�=�2��ꯪ�1Vr��:JEI9#���ǽ�=���6\�c�Tx�hfH
㢭;lM[v�X�z,w�V {���I����b�W�9�ދ ���wm�M��&�X�L� ��x�dX�z, ��p�	�M*Ğ�;��vrFKz]Bt���V�خq��-tIDv8�7l�5)��m�����^Ȱ^�X�L�t��CJH܍�'%��{u�W��G�o;?U|�f�Ձ���7�h[�9#�8�q�� �镀m� �� 6]�IA�;N�Wm�w�V��,ײ, ޑ����մ�b�%i�|��@o3wg��f��n�1E�U;�˙6[$�!��M�3�\Ş��h�I��v���(S[t�p�<b;�It��燁��cmh].ê�h�d�v�
�r!t.��$vg��[�1�LOk`{	��-,�,D[)�.v�9svA�%gn�nƞ�b�%���78nG��[Qz�:�I9�U� �mnq���&؀�n%�nX��`3��l�ʌ��#$ݧ@��s��\����w{�=�x5�����i�u��-�i��V��)�zY�Vٸnr\F��6�t�T�1�uv�i� ���� �+ 7�x��������-+bI� ޑ��e`� 6H��Q��t�i'v��;������gH����.���$�IS �o< ޑ����2�	Ү�m[��m��-7��<׽�&V {z_6ߟ�~�;'�C�7�:�ͷ���D�l��2�<U�7S�LZnT�536�u�z���7���oG�oI�����A�;N���X��X}�P��`{6i`~^�w���|�v�%�5J8��I:������ ��E�oI��z�H�6�[wWi���7���ދ ޓ+ =�躂�:*Ӷ�մ�3 ����oI��ޏ �٥���ң6��(QJS��(&�T���=Lb��e��m�V6&��V�y0�Z�6դ4� ޓ+ =��0^�XI(�R�cn�m6���oG�^9e��>P�ҭ�Q��qN�zE$�H�rX����k�����UP0G���7���9$�����$��i$�m4�i&� ����{ze`���=�2�eKB��v��$��� �镀ޏ �ɕ�{WK�;ۢ��Wv�V&(Jc�7M�$h�Nܚ��W7:la�Hҷ��Gk�k�ӱ��8���I:����l�X�t�w�V���t�wWi���l�Y>��7Mw���^>��
8[�@��i�bj�m:����ޙX�z,��+ �^����t�j�v��=��P�����J�a/A	w��(�E}_T��q�E:N�JrFԒ���`ޙX�#�=�2����Q�x�<�,;k1���α�3GWnzw<6����ĳ���^3E[���I�镀�<��+ �� vԥ��m��m$�`� ����6�G`~�m��}�}T�gW7O��'�m��`{7���ٮΪ�/f�Ձ���+��qKWV�M�դ�`��omՁ�{5�r�o~�˻��$���M��oL�׽�镀ޏ$�(���J
U}�^̗�W��{a��a���6m��7&��d�v;!�^[v��-j㋵;�V0gۑN�dWu�1\��Jn;un�z�I�[�S��)���tLY�V'���i��n�K=K� S[�$�z����
�璌h�ێ���j���//��R�C4m��v�ک`�m5+<�:6�c-n��lr�z�NR썮7mu��.��E:��˹��p�݆��3k= �Ţ]U��Um��f\b�m�'�ݷUۄ�v��M�뀗���=�2����ޙX���"wbn�mZT�5�{�e`���=}�`�����St�v��X���oL���+ �镀{z�cM�m�m5i��z���t��t�?�/� n-�e��m��m	5�{ze`�2���,�7]��B��Z�*4�$jQ"���%�1���qzl�]RN��#vn�ʿޟ�-,Ӵ�$�n�I�+ =������}�W��� ����r<��rI<��w����2�׿}��{��V�6����5:RTp�*Iʑ�@{��h^:TlB�s�Tx�h_PY�i��5n����镀otʰ�͖�UR[����Z�C������9�T6�PD.^=� =ݚ��+ ��*�_$��J�o�ت��I1�g9�ɟNtqF�����n��2'�{���ö�VR-:m�n��?< �#�=�2��e`ީYm��m��6�s_G�!(]�~�@o�}J�=x�&�A��i��i��m�ޙXI2�=_I �
Z�'"g(��L!�s�ď��
 R%���$Ձfꏏ� jB��E��1pȑ�)IB\�x�(}�7�y�~a�����E��Ċ�z �*�>!�K���@�SUP�4 Q]A�5UC�D?�@��!�������?	��?����� N"T�lIw��T(Q��wʀ/� cnh_L� ��W}um4ح+I� {z<RP������iPۥ@[B���N3;��b��k.d�j�X��Pr�v٫���3�2i�e�Nd��1������t�m��J� �{4��wȤ�N�V�I7�{ze`$���͖��/��H�U��$9)��E�X���V {z< �#�=�2���m�wLNT�(�%XuW�{7��=ݚ׎�(ID�(�!A
"3c��W@83�y�I>���-�;M�ݴզ� t��ޙXI2����]��j�LE[O�-Yn0�����5�ٛ��$�j
ъ�:�p2����0�m�M��I�v����V�L� ��x�G��hPwCM6$�NU��U�s�x�h����t���_RA��-�� ӑ�*�=���1�4}���T��T���*{#n��:m7�$x��V�L��|��zX[BU��NG�JrX�*t�׎hs@}
!*��w�������}w�E��ֻErWju����j9V�v0�.8��8�����=�<=c����	���`�X"ydƳ=:�v���Y�:����P1[�6۠�n�X|ۘz��k48-w`ʆM@e�6J�9�p��n�瞐ur�s�<	\��ga���nu��A;%m�-U�^U���C��Q���n#7l.ˍ,3=��4p��'��護�����;�7�a~=�^WƷB^r(&��OY(G�����Q�PT!skn.9?�w?9;�|`�sR�w��}�Ԩ׎hs@z�Ҡ3G:��e�M�n��X���I�0	$����"~�����6�m&Zo���}4�Q�9ķw|�q���?a�'$m�q�%$�����{�X��+ ��E�H��D����l]����@6�*�}ǽ�����wV�+[[M
*t�7���,��p<@2�gZ��9�NE��٥jNs�U�Y��$� ��E�H�oL�I2�đ!7M1�uv�i� �G�G���Ӹ����J��/hq���!	��պM�ޙX�ea��ꤏf����`~^Ȑ�$it9�T(�����@�f�nh>�U/f��7{�L�7)I�$� �� I#�7��$�Xղ�-��V�r� ��su�Xh��vvZ�š�z`\��C�S��U/@��m��nh�,�n��BI{�cݚ ��~��I6�M*o ގ�e`�vX������� ù��EJ8�;��92P���񹢢IG!pm��3sn�յ�k~q� ӊI*þ�(P��{�@��@^9e �t�͒�&�6�&�o $���UW�V=�<��* �nhIE���s����[�l3�8W�.1ng���V8�4�q��r�[vrDo��ww�c��35�.ʷ�t����I&V {z< �G�{U�K\@�$i0NU���u}��U$��`�����۫ٻB`��9Q��\��@�s@�4lB�r��*we`*}1�i:m��ݦ� I#��~��9$���I���A(�Z#s�����-���m��T6���@jIn��x���m� ��t���e�ۧ�����g��eħ匬n���Ɔ���.�[�d�R�6F����uՀ{z< �#�=�2�jWRD�4�b��m� {z< �#�=�2��eg}��Vʊ��I+���L�� ���vV {dx����"��biJrX��u`fn�X�f�䳻����\�prS�4�'*��ݺ�oG�$x��V���4����k&NU��i��r��b�Y��棘�R�4�����^#�sBzw-o\,*1�Y�!�d5�1%^��{.��=)�!Ⱥ`�KwU�!��rl*9z���e���Nb27<ce��`um"���Q@%F6s<��ck�:��t�c��Ğ��Kfw8A���U���h�82�Glҝ�юqS��ů��C/�Ȯ<� O�_99��2�3v�7I��iI}8�ɞ�Iu��Z윂lS�k�m7�z�k������F��m�M�nۭ  l��ޙXt�X�A1�i:m��ݦ� [nh^:Tct�׎kT.p����6��m��T6��?e`�e`����< �.���M��`~}���֨�4m��=x�P�GRD�4�v�$�� ��x�G�z�Ҡ3�@}�vy�(��x�#��wݺ3�.�����ѹK����V$�f�ٶ���N����O����p��$�������2��2�zG�{Uݕі&�q�nKٻuh�����h���`��`yz��	�n���t�X�#��< ޑ�!.�:������IV_UU%��,;������:L��T�l�N���Ps�4���	G�����7~���f��E,H�M8آ�ڸ�M`l�{K�J�q�S8������u�jܼ��V�m��6� oH��2�zG�m� l����[M6$��o �n�jP�.p1�������s@K���S��M��I:���$\��?�H��(�b"(�"3�Q	W{�]*w�P��+���wWi���6� ޓ+ �+ 7�x�]�]bi�m6+I�y�(�DD%򈄖��Z��}4���(Ʃm�#Jl"��R�wMٙ��m7f�ٷA���2�pcpۃ2b�a�զ�zL� ޑ�}"���^��o]X�r��jJ�FԒ���e|��3�w���T�t���S��	'M������`ޙX��X���u*�v�m��m`�t���P��lB[��<�RT�s��-؛�r�$r�f�Հ{z<o�X��V.IG�u���켣[���r��nm��֖�{vZ�к{N��ݗ[5��י����Ͷ�~���`���镀oI��K���[t���q�%��U�=���w]X�۫ ��x�1]Ҍ�4ڶ���x��V�&V {z< ޑ��Z��RSp��9V�UR���V�ޖ��X��V��K)	�I���X�����`ޙX��Xү��� ���Dg�\�1�q�j)�xA"TB�0�DI`�MG�<P i �A��8S �T&մ��a@��4�$ہ��B,D����+A���pD*� ���#�01O{��m���I� f���VI�vU��{$]�4Q��m8ö��[jWh%���.$HD��V�ݹ���l����Z5=R�*2��;;[�GJP �ɓsm��I,��/j:ͳ��yy�s�m�on�����&����,{Wtݢq���K�.�����ƕ��ؖ�T�B��ΐ:�l�������1�՞�jq�Ĩ-�)D���S�u�\�S���.4��kj�ڧ��t�k�6��,=<��j�0�R`q���n�k��]A�a����m*�:��\�[�`�F���)ey.�	i
�/.�cl��m;P�`6�V��m���F
�8ŕ�����{�kj%(�pF3��Q�l�19�I;Ye�aw[I��N��9*:�`gB�[��L�ζ����h��;rbض�v�{�ت�n�w^��آr&�fy�Si��b(h����,�Prc=Ėz�\�����4��g6�I�u����	vlѹ@�v2P�1P&��:`l���c���=�ӋO+�-ٙ�R�/2��փ�XRR/�N��YV��v;gk�v�F�lN���.�&f��2�[�-�6m�sQ�y��6xKiq�E%�l�UM6t��F�\�mڷ`z� ^],��H���,h	]UU+�*�Ү�4��2$�v�mc[K+�k\��u�[mS�q�+�w6{U̬�Of�*�����g���`�.r����%צ�,�M����.��-����Y���*c$j��\κ��L�lq�-���Ͷ��K(@	����l[dR� ���^5���.�(n7=��u��,���l��ayj����rD����6�s��ƥe�h
�В��ny�,�l��L��H@ѹ�9:����*y늶��tc�,b0�k����7Ν7>ڹ�N�)�6�/[c[;k��1{G�����oY�x�ٺ됐��۔�^��� '��qAz>b�C�T"@8��"b!� qD���Pb�X*�����x�����.��{q���s��C����9ݺ�O�=�n���;���L��b���<��C��f�.K8o=��*�9:X��g��ncvmc�v��L�F�qm��p�.�Vs]�1��)��]N ]v�u@�n��Ûc�v�%���Lj�;E���/N��!(]nr7i���*Vأj��m�N�N��I
��Dmf��M]�2n�4��7s!��͇<�M�j<v^�.v��1�z��/^-q�-�fx(�59(���GV�톾m���� ����6I��ޏ �m)bI&�i���x��V:L� ��x:G���V�M�&�N�	�e`���	�<z8`��S��N2IVIf�K ���f�X:��t��_�n�cn��6�x:G�{ze`���oG�t]w.�<pO�^}���d�q���ZMm�+�hs�q����X���3�9�I�V�m�?߮� �T��:�G��٠��w�>�.陳d�\ӒO��~�Â���(�	B �V"��H��C�* �^"667����|��������x ����>A�����~��'��4�����pA�6667���x ��~�x �{�>�|�������>A��������m�34��̒�� �`�`�`�~��o �`�`�`������� � � � ���xpA�6667���x ��'��f��n���3ww��A�A�A�A��~����lll~��xpA�6667�{��A�6667����A�666{��{�;�:�$��Sޝ��j�DlM�nYצ����\�]dn�n�S����L�P\ӂ�A�A�A�A��}��� � � � �������lllo������lll{߼8 ���L�󛛛�.M��� �`�`�`�{߷��A�A�A�A�}���� � � � ���xpA�666?}��|�������ۅ�76n�-����>A������o �`�`�`��߾����lA�@q�@5A�A� ���xpA�6667���x ����̟lɛ��w7rL��>A���"��A���ߎ>A�������Â�A�A�A�A��߷��A�A�P���s����x ���[�g��wL͛%��|�����}�� �`�`�`�{߷��A�A�A�A�}���� � � � ���xpA�666?�����*�����ص[t���L�%r�ӹ�m4=a��O�6��Y������8 ���x ���}�|�����~�Â�A�A�A�A������lll~�i>��ff���������lllo�}��A�#��D29{����� � � � �xpA�6667�{��A�666?�}~3��������f�� �`�`�`��߾����lll~��8 �����|�������>A����>���s0����wm�� �`�`�`���}��� � � � �������lllo�}��A�66
����� �s~��!�����ݙsi�2�1��m��n� �t��y����\nxy����&��� �\%d�]Pv䣶	a�c;Mk�̂�����	$x�L���X����W�"1	�մ�7�{d��磌�7���3zXn�ى4=�RS����ʠ1�J�.���8=ݚ��u`n��6]	9Qȉ$� ��< �#�=�e`�e`8�#ē��H�M���+ �&V {ٲ�_UW�K��7��&ƾQ&3(dHx��( Z�Ӊ�%hWg�pAB���z�Pg�g�2f�6n��a֊�;vDvO����Ǔ��]V�d�j�u=�Hݻٍ����M֊l�i����B�6�=NR{=��o��u\5̓����m���v�Ɏ���+u@.�B=�h�2�	��ՠqjG��9�$��]�Iv��m�:�������Y|���9.=���[�;t�Vm����.��fn{,�͖ъ�:�l6�书��e�{���L� ����"�
Ӭ脪�i�m��u�wI����$X�L�����҉M��M6+M��`t���"�=�e`���
��:��6��M7�K��+ �&V n�x��-�m��Ҟ�{@zۥ@jZ�|���h�o���}�l/״y\x�6km�#2c�=d�NĽpQ�V����	*p� W�,-:�'I���/�X�L�wUm:h�r��H� ��e�U)�C1qKg׿}��{��rI�d��6qDF�'M��v��%� �ɕ�N�+ 7z<�D���m&�M*��=�e`$��ޏ �� o]�DZ-��v�I7X�2�w��%� �ɕ�K뫨�ϓ*�s�زح�:�\�2a��/-��v�1��t5��ґQ�)Ƥ�N7$� ��e���,�&V�&V z��j�+m�]��o ���+ �&V n�x��v��Bm�����X�L��~�{Ò�)��WAD8�1d��~vݽ,��t�ē����`l�+ 7z<��X�L�d�U�W�bt�v�n�w��:�E�{d��6I��tJ�T:m;LN��!$�c��w�ڌ���nb�L�է�y��'#�Ŷ$�6�E�o ���8`$����+��M��T��l��'GL�G�������h��m�n�`�2��G��x��mJ�h�I�m�l��`~���ovh^��ܲ��%B��(��� 뻽�$��?{ۖas.����i� �#�6Gt�X�#�?o��ݿ��ۄ�[�I��p\��L��\�-��M�����em���q�	��Za��$߀�ߟ� �&V wH�t� ��$�{NRp�Br��ՀgH�t� �0�%V�^U��6ݶ�� ����8`���7�땎�ē��H�M���8`�����K���m&�M/���6Gt�X�#�	�<���{����V�c ��d�&�9�b�ԍ�����V��K��v�:��Ŵ���8nܣ��X�ܵS�\�y6�q�K���n0%ɻD�՝�;�jǐ�+�]�n&���f��J��0��m¤�W�Z����rs�Ƹ�9�u]:-���G[U��+�TY*,i,
 x6��&8UB���p��a�;m���̹��o�_�������VpX�Bco{���|�S�὚�m�<gv���Zg�-�V7L�FcB�/����� �9x�������>߾�@�� <nI(�7�WV�g8ԐI�$�`���$��#�$�X�oP�J�we��o $��#�$�X�#�']�nЛnӴ�o �0	$��� I#�=²�;�N�� ㅁ��u`w�R�;����٥�f-�1�IQER4�/^E/��Yyf��d\���5q�wM㞦*�e{�Yi�m�m��� I#�=�e`I��{g�)e�$�6�E�o $��pS�	���Q� p���=$��ޏ ;Iqm��M��m��&V$�X����< ӯ�!"�i�m��u�I&V n�x$� �ɕ�mJ�h�I�m�i�m� n�x$� �ɕ�I6����Rw"�2��T��U!JD��ڂ����n�/C5Z]���s�mm��'�Bg��jěm�\�`�2�	$��ޏ 7�K���M�i�j�M`�2�	$��ޏ �$X���}ݻv�eՖ�`I���[�U���	$P� �c�D��j��ժD��� hH,H1���_W�����,d��;� HC�� �0@�E< ��CO�g<�1e���!"A���RU�c@ XP�	� j�(D`1#� "0@?�����8��}R�z$A*x��>(?�F���!��P�=ID]�߻@e�Z��5�8�ʎs����V�`t��	rE�{d��$�+ �ʂ��X�t�ii�\�`��P�J�.���	B��szs���ZZ[E�--�Lg�J�$A�2�{U�T#R�u��N�5vP���$���+ �� ���\�`iܮX�m[m�wv�`����,�&V mJ�H�I�m�i+l�ޏ ���+ ���Wf�E����r47$�X~����y�s�=��TfK(8�D�r!x�o�ɔ�M�i��6��=�e`����,�u�"0v�lb�n�����32V���6�-�lW�.�hq���8�MD�Br�̚X��,�H�l�XΗWh��Zt�iX�0������y�J���e�ur�eX�t�ii��$X�Xw8`� ���Cm6�m m��&V������"�+��Cm9mH�r�̚X��,q���T�$��%�����B��I&�xK<&#��ɴ̒M�ێ�����^˞JCv�Kg�����n2�r�Y�%	��`�ړ���I^t`�{x�\jzO͘��x��sTF.�M$�%��X܋�-�q��eYc��C����)e�3��Z��yǮ7g�ڠ&�uJ[�vn[l�6�)5A\�a����,<����:0/?MVH�%��3I�wb�|?y�	��'	̧�ɞR�-I�K�͹��t�J��`��K��Λ:W�7I:j8ԐI��0�������&W������0	ʉ��ZM6*I���=rE�nɕ�ws� n���m&�I���X�Xw8`� ���\���S��.�Ӭ��0vG�z� ݓ+ �����+N�n��L����
��������Ҡ=Ƹ������:��8�oblq\e;^h��$�m%�/3kQ!��\�n�\|�}?dX�X�8`� ;���7������&��$��w�9�p@(!��#�`I����`�u(+M�J�.Ӭ{�0vG�z�E�nͺ�5e,cZ�A�����K3�`s��nɕ�N�+ �Tu�V��i�V�M��K��&V���#�&�8���]:��Z)�ݵ�eG�%�ZX����4;�b�h���\�����ωjI��jƩ�׀���+ �� ݑ��}��w;���&�2:��I9V�K+y��ݚ��{@]�J��QޟO�ʄ�ϒN�m*���<��,��D=�*h�3߾��'~�{9$�����F�I#bNK^{����{�0vG���);m��M�Й��mҠ>�M�����@{��`W�}Uϗ��W$�n6�J6�Ξ^� �t��&�淧F`sIr7��%�-��.�*�v��˴��I� 7dx�H��2�jr���M�Вl���|��L��}����@fd���̕j�&�UiSM��z� ݓ+���Kwg��,U���H�q��O{=��B�f� ۝(���@=( A��o9�����,�3����I9VfM,�Y���]���2���R�IZ-P��-]'I;nN�����Y�\g�V��Q�i�.ra�l#"��������Z�����BI� �����"�7d��;�� ��D�e�4�6ڡ&�\�`�e`���< �u�1��m6���7d��;����]�������`=��Dm�mH$�X���<ײ,vL� ڜ���8�i�9 ��e��_y�s�f�*�%��K�" �P��@�	�F���%�m۴���C��E����z�����;VG��.��ey4gd���?�l:��Y�&mz�c8�k��c���� �����9�=�w"<,t�-�Zғ4�̮�.��6	�@��rP�m9Ƭ/%a�s�]�P&���2��:L�u�Yu��mu1�kj��8m����N�NmIv=BM[�y�Rf���s�r�OXn�2�Ywa��,��n譈����t��%�:�8[%��N�%��1�����#��G$����`Wՙ�����������`v:�l����q�8����n�~B\��J �ݚܶ�Q o.
��lj���uv�`���<ײ,vL�g\BBYM�um��L�����&Vﾾ�X��u7ldnT�:�������2��p���.%����sֹ�l�O�k��Xn�%�쳊R`�1^gYn��,�Mm4�M�����2�{&��nί� ���`f���$i� ��`{�4�W�:�;���� ݓ+ ڹ�+�I�m��]�� �nhr��.s3v���J�5���n��K流�w;3����� ݑ�s�����m4���M`�e`���<��,d�}��ӣ.��ŭ���=rQ����G;E`�a�[;�_��װ�j�3T<�׀���<ײ)^���6���IJH�n�1�-{1���Ձ�ɥ�$fhpUԔ��䎎�f��=��mҢ,Q��%	�$���'����˒��n�m&�@�X�X�8`� �� +wZ�ے4��JJ�=�4�?�Y���[��{v����X�5�NH�7M�]1F�Z�c8,I�Ŋ�n���:C�+�����ګ�ն˴ZM��#�=}"�7d��7�� �����Zi�V�4���c}���3v��Δv��Д/�#�usur9n5�;3����� ݑ���`˨-%.�rH�5%X,ݾ,3�X�n���"�_���ޜ�}߯�&d��cm��L�����&V�ɥ�m{5�:���9LB'm�Q�Ǟ^������C�TY���O#��WgI��I�ײ,vL�w�?��X����z�PIr7$l$����mW�9�1Δ��4�m��,���ӒD�q%%X�M,�ݖUW�ygs�3;��#q�*q� �����n��^Ȱ�2��p�=a���4ڴ��m���`�e`�,�����ʈraz�a���"1��x�	�Ȥ��* ���y���`~�HWď� 
D#B(�IV~I0@qH)�X(�i��J�iX���IIaでl�c'w�ٻ���d���6�����M���[�@r�pvv�T���Hc��������F ��B�  xH��"�G�`E�������ݶۖ� ���fg����Gd�g���U*԰1�:  ��X�ZΫ۴���h� l��,'%έ�7F�5��`�I怊:��`�U�����vt! �U�3�n�Uʅ�ݴ��lCd�oI�盬;f��qH��X۵׹���\��nsӶ���Q�Z4�i��F�9:Qxx�䌛��+3�DЀK��m�B�q��$JL�)����!�J���+<ڳ܁��j�I�&�f��b�����%�4�-�tɸ��qk%�kH k�̕�3i��`����)�s��u�f�*F�B���:T�R�r�'n����ò�K�RhU�ź���,�Į�T�⭜����	�J SmuW�X��5����<b;j�p��R'i�{F)c,�Pr��cn���ץv�� V�f� �gD���̓Y�2����m���.H��]�'5i�yPҶ�:��F�{��m�[�ÂZns�Լl��Ι4�˩�n���ëy6����s�������[���H�f%l�j�6Z۲�'=�Bv�j�]��K�U*�m���k���srU��Y�A�Ol��:���V먷([q�s���F��qq�����Jy�pV�m�v m۰ ��Y		�N�$	f�q �UT�kƭ�"S���-�CgP+�S-Ԋ�6ڦ��= �0�nA�%@�U��j:Zz���΁��K�"˳�UR�T;l��q-�5T���BCm��;fݲlܑ�ڥ�K��O��sk�Y��K��k��6ݜ��a����J�%Z�q�-�UԪ $l����=:1Cqd�vv�
vUI[��nm��: ����0ZZ4�.�@TX��&d�fZ�#+��7:�v�v�<��)1c�l$d���[nĻM7m=�eZK���H! ֻF�\�̀� pJ���8������nC"rX
�'	��w6�v��Bzw�6�k�|%U0"�jǊ�^�~E/� �q���	����`��O�
L=.fn��.M�:ۢ��H斷j�jzvy`�:CmuW/�����nME�5a��a�`�\|7ϛp�|�OA���ձ���\�]�kI"��m�g�7'[�.&�	s�'&�vH��(g���X��"�\һsm`�x��܎ح����hd�N�np*�'�A��F�q��i�
n\�٧:��՞��]P�g����������|����;�	�<�6��[��tpr�5f8�=7]�:��m����:O�������f�i�նƚ�we`���;���`b��`�AS�G�)*��d��D(�3vh���v�*�(P�Fn�`���#�)$M��3;����E�nɕ�os��:�v��V�CmГx��X�X�8`~����K3�Xi��#�9�6G`{۴��cu��37f��1��y+�;ӱ���n�a��Qi8����-�F[��7U@��Yf���|��\�̃0ߛn��0vG���&V�ND�)��we�.f��~���?��N�R������P�����@7�Ԩ̖_�U$y�'�6���=���ݓ+ �� ݑ�T�i�&Ӟ�{=���fh5/�(����֨�?�۲�����K �ܴ� ��#��N��p�l� =�<w�V u}��ݭ���K�:��@���)<ʹ��V6�q��9�Y�^ۜ<�%�i*��P���cs@]��B��f9� �%�FU�I���Zo =�<w�V�����\����v�}�34�:T�K(�(���":� {dx[�
��j�4��A��B�{� ���@�总�J��'"[.�V�.�v�0�#������ޙX�8`!w1�[(��v����c��A���ĉ˘#i�8�4�zs����������|�x�V�_�c{��n���7�� =�<U쨓�rH�i�$�=�۫���#7g����t� =��#lT�lM&$��/2Y@�揢"9�����iP�D���M����&`�G������{Ò(""�q��|��U]��e�� �2�D�d�SNK �74�Fc�/�Δ�nh��a��r�T�O���k��%c�h�e;U�UbF�^���dM���ށ�n���7�� =�< �H�v!@�n�j�M$��{�0�#�ٻ,{6��#��(:q� �r����t� �镀os� v��K���j�Lm� �H�ޙX�8`�G�M�12Ěm�������+ �� ����#�3��~w�~��&vKY�GR�3ON��ʺ��r���ZW[l�s�n5��ܳ&R��9�M�=��Z���PkGd�^���������*�C�����;kMTİ-��$���e�ˁɎ��®L���Ν*��D�Q,5�۪�tv��ltf&�yv�y�Tx{-���l����h/h��5t�j��d͒x�hv:S�c�v[2�s?�P,�$��/lqjZ`�)��ЏBݙ���vh�͸�/��L��JՎf�K+wͷ����� {�x�L�{��b��V�J�L���� {�x�L�ٓK�+�H�j9	��q�ICr`�ߞ�&V����ı�Vݦ�6��m�w�V�����G��
�v�V�i$�`��� {�x�L�t���(���\
Z���kxw�u#��M�K��.{W]��=jr�<�3Y-o��٠cs@]�@^d��<��;fannn���ۻ��O=�w��(4K":s7iP��@m� ��u�V$�m�ժI��nɕ�os�����gt�ot�?/
����r9N��p�l� ;z<w�V��h�^Rn���i3 =�< ���ޙX�8`�EԖ��t��N��ܾ�9�ب��U����K:���3kT��E�N�$���BM��G�nɕ`~��,��e�U|��r ��ND�i}v��;���0vG�� n�v���I��=�� <���% L< T:x���Ovy��2�r���IU��b�j�0�#�ޏ �镀{c� z�:X�]��V�cm��G�n���=�� =�<m)v�;Mة"��A+r����3k��p�X{�9�V.��T�I��I��BM��2�lp�l� 7z<�T��Fˤ�bi����0�#�ޏ �镀{zZ-]�'i���I����G�n���=�� �����*�I��t%3@x总n�v�$�%*'�=A�<�>�y$������ݦ�6���n���7c� {dx�#�:K�����v�m�n�b�[�l	԰��k]�,�Xl�\��u�����:n�V�����=��� wtx�L��uEJ�*�i�Z��x��wG�n���=����6�4�n�q��nI`�����n�E%��G�N:c�ڶ�m&�*k �镀n� ���?_s��������N9��V��K���π���(�t�T�,�,�z�Fw^\φD:z.�Gn6Ӷ67��rZ'��MvCu��n+�E�hV��wK�.u�X�Y!cŴ�X7,���*�:���2�=Y�w*ʹ��]Y�NF��Wa{'0�kcu٬��d�	ڬ8l�mm�v��m���O6N�n�v�.#n3t�2clq3�Yq:3�v�CV�V��t��ة����]|�s�a��d� X\0��̔�LA����zC�֛����1u�;T��7Mऋ@�RdD�)$I�x,ޒ����=�ۯ謹 ��Ł��p����q�ƛx��ޙX�p�:����$g�D�8��JE`fo]X�� �ލ��K�6U�Bv�����7c�׽�7T��n��X�f�7��r4G��ٲX˥��2�E%�]]L�:ˏPnF����]`y�zse�l��z���N�ΰ�cMʵ�ֺx�WEW�����0=��ܸ`m�y���e7�J����n[���O߽�x��`# ��UU_cC����D����ӒBW�M6&�I:�=K�މ�����2�l,�w�bm�m�m7x��<�t�w�V褼݂ԕ;�����q�1��7�W�=ϹX{5���O�i6��>�ͳ�K\oa���a���u�gU����kY-�#d4��M��M����7ze`�� 3ٮ~A����a�]*'�H�ݷX�p�މ��K�7zeg�}I��I>�6�i��,sy�	��w����q�u�_8	�â�$kB��T�X��#'	���	�S�N.�H�9\p�$d�w�o�(G��d�0�̐!3%̳-�)BC+��s���8A$�'�Z�0���?Q�@���D��A�BĊ/�B�0��&]%}$`�a##1�D�!`��	���D+�A�/ h��/�‿
��hz"<�� �*���o�� ��ŀW��G:I�#M����j�J3'w�c�TۖPj���7��7v>R}RI#q�M�`z�Ҡ>P�f֞ x��@]��P���>��p�����]q�CǞ�͸+���Ǝ�8)趍��r�v6P\9e�f�4�X�p�މ��K�7ze`�V\��N�m�m��f v�O �R^�f�X��/���#۩pRwBm�6�4�xr���ޙX�p�މ��%tJn�v�i]�w�n���=nY@x�4DB\����߻@�����$�GRU��l����幼��3r�=�۫�zR�B]P����:6�֩��k2m4,�<7�[���U�������Lr5J8�m����X��V��u�_�ft��+�f��#MӉH�����_Wԑ��u`ft��;z'�v��4�m�ڡ$���+ ݎ��<odX�tU�j�M���N�����6���}��D(���Z�3~�t�y�]�ve&ݫ�����6�E�n���7d����ٵ��L�IBCi52�Vճ��t1V�k��:w	��0����s����zi;l�����0Tmp�Z�d4��r��
�]�Ӏ�{k���m��j.�����	m1#.��8�tu���H�r�k���l�s�5̓��H��۵�+*��]P�r�n���2m&�!�L !4���f-��v6�)p��c�( 6ѓrL��$rMwm�r��?�~PD����xhj�II�P���*�1��v,.h�a�;F�U�E�7[�̈́�7`Y�%F�����f�X��,=��xըbڑ9�1���f�_U}�}I�8���,/n� ����m�rH�q%%X��,=���}�X�����Vz��FƩ��M�!`x�4���w��В��f֔�WO�T$�jҤ��O ����+ �R^ v�O �\]*�)��,��X��z{q<M3-#n*͛�Gk���m��SۦӫM��mP�k �镀z)/ ;z'�u�E�n�e�m[t�n�����9$���)�>z�U7`���.O� ݓ+ �IH�w����6�
ۼ �����&V��U��0[HN�I��$��r��y���n����@��4ˉ�:sT�Ȝ���~3��������t�_�7w��1fk�=��$��iP�*8lC����J��;F��FK�#\Ω�V���}���C�E#��%~����ff�`e�E�nɕ�um(Q�M4حXӺ ��٠3;���t�>��iG�/���+�~�CrH�t����{��~�����"
H!�(�Y	$*럧��=�f���7�\'���i6�&���e`�� ����K�7y�ډ��M6&�I:�7\��؈}of|gwy@]�J�/gݯa�H��x�u`٤��n�I��iOY�����ũ�=�<��0�5-�lu�F��%��e`�� �qr���]�Лl���7T��nɕ�n���ř�_}Iv�!��D�NH��xw��X�p��)��"�6��-�v&۶�I&� �� ݒ��6�AJe(!H���B�{mP[N�9�N8�m� ��jX�Q
�d��ݰ��TfK(p6�N����20�麃��::�E����k�%�a+��u�=����T���ͷ�}�.ۥ@fd��p��4�t��$��m4�&�X�X�8`��_H���tuh_�M�i�4�I��?� n�O �� ݓ+ �Ҙ�`�rS�6��a��guK1�*�T	(�^mi@[g5p�i�{,rJ�,y���3��~�Ӌ ݒ�����F��.ĒJ��j��gB���G�Q/9t�!�v�v�v��A��U��x�h� �B�\��n[�on7j8ά�[m�\�.��n��^���P�j.^��2��T�ALE�m���b3�H:�ktڑm�j�]ҋ�v'm:����@�I��j���P�v:�9���xvە���/`�3K��ss33-����N]�d��g�� �A�w����;�;���%��4��V���]]���٠�^S�:����u�]�k�W#'�3=�9��(��*��vڟ����Ǽ�U��Bj)#�9rU���%<oz,vL����%J_�T��A�ڐ�����U��UW�Ifw]XΜX��F-�CrH�I��x��x�L��0vJx�t�e4��m4ݦ���e`E�֞ ��S@]�(��pp�Z&�[��]x�00�v�Xg���9�e�x�ӧ6z.lW3Y�+�m�?�o��vJx��x�XΫ���;OL���˻��I��7��q`���BĔDDZ��IE���@<ݥ@z�� �qe���&�ۧm��n���{۷Vu|����ޒ�7+P�5���J�ӼvL��0�����^�[�]��m4�i&� ؛���s4g[�v�*�����C�=su��7c�:����8L-t�	u��K���F��c���z���/U�4� }�ߝ�3��n�o��2�*��]	6�I&�v��%��e`���-����44�i�s3��T���?"<D2"9�⏔(]Q	B���~��s��h��w�z���i�4�۬b����x_H�?����Y�ߪ���\�i�9)��H� �� n�x�X�8`���������qf�]g�;3��l-<#7b�����K0�'m
�_�{��F�n����mӶ��	?<vL��0��x:��%lm�m���7�nɕ�ДDG8^l�@����9�/��9Whv�M4�I��=�� ;�'�_꯫�6c�R�Ifw~�ߒIVS��t��A�ڒ�Iw��UU}$���?~I#_)�m��w�ym���k����(Q�z$Q�s�%���������nn�I6���]ݜ���ww�'�޻��.�I,��?~I-ͻi8J���C(� �ƇG��*�f��l�
ҏZ�h`f�rP�\���2�1| ?��;����}��^��;���y��}�ZI-���I��k!ߟ��[�> ����~~vr��]�{�z�뻾���Ct���7��Kٚ���$���i$������I{6�-$���~t�@j8�$�H��,�
�_w�]��}��<����xN[��n�$���&���E$��N)i$������I]vo~�I$�yݤ����m��TW��TW��D��D� ���(����QE�E�A��D����"
���
���D�D� ����*+�eTW���"
���D���*+�
 ���AQ_TAQ_��PVI��c�S���` �����Z�                        �@( @*R

D�J��� (J��
T�TIAI  P@D  Q   M   P  QL@>��9o=ί�-\Z�[�U.����)b����;��rt���=n}O>�f}t��� �Ν��yK� |>�yr����+�ç'J� ۴���}3T�,�'.���  �� U  P �d �������{w�'���Ïx>���'%2:���n�`�{�X�z��y���{� �,`�P� 6� R� 9�( "�0 � m` 1 :M s �p @
� PP1 � @�@�n� ,΀ ��
2( ]` ���QZ� �` ��  {}k�ye��� �{Z�=u.[��ז��r�/\@�y�NN�m���5���n.�^ >� 
  ����}4�=�x��^=�x   �P  ��޷��'K�����m�
�}��{���� m^m!}�ԯp ���={Y�o���..{y��C|�\_v��;��<��NA� x  @ TS�
��6����g��Z��+ݥ��N���Ի�8�WW,�7 �����w{���7��/sＯo�����S�t������.���{��ޥ2��Oy[������� ��iSإ*��db41S�#S5)U4��D��IS�hi� تT4R�  U?�	S�T�T� ��&Ҕ�� )�'����g�������rv�����w���g/��(��������(����QQ_�EEb�

���葯���,�
����W4��I��NM�-�r2Jp!L
m�BB��[�4��J!$�� F����.n�+���֬����,(d��[�|���ǐ��������.�o�梨V�8F	� �	"I$�$Z�	Sxg�#HF�����%�S<f@�0�#$�X�� D��
0�zт�R��p�� S%M��0$GҒ�"1	�%�CST?$
�)āS �q���� �!ȗ V�"D%C$&��b�%��F@č �uabV��`�@Ph�c�^=ap�� E�q}�H	`�� $ā,��@��D��M�F��S�v �`s7t�H���"��B��0��]���d��c��C7�Y��	 �*x�~=Gq?1���� �p��g�KX�EjB�@!���j��E�0�ЉJ������)�ā$��F��@�@�	�� F0��xC�itabQ9���h�)����!H�"BbD�E���	dy$$.�`��F�B�H0�H$)�fi�XV��	,jB�� ���
k�@H'凢�A0�,������"�(lHB�B1���Lp�!aL\!j*ę�r%�9��H��D��B��0���!#���"��14/9��9�$.d��\�0���2�~4��$ ��é�;���s��qax������V��Y�IXTt��~4揿��6�����㿿P���.�5���n$�&���\�p!sB\��]�`P"j��)���E4u"�=Ŋ�8���qz�
���8e8�R5���7x�F�^<4���Qi��p9$k�nP�ዦ�HS�s�\�<��efKm00549�i�7��dm�$�4�
�k�F!��c Ґ���q��@�Ӈ��$���c`�&Z�Je)��2�0�#�5�^�sm�D�e}8�t_CQHz%x@�X��`N��#$���H�|���T��?+����L2�0�e%C�Pawa��Yr$���8j�@�F���x�n��x	�=�5��eמ�?��_	L���ee���lК�I\��7�*�#��B� xk��B����l�;�*�
Յ��MaL�j��!kI�2nq%�7�~�ҘI�p$��)1���͹9l���3��@��)!��wI�3<����1`I?r��%}j��w�I7�$4��|D|7�f�Z�f��<t�|OHT�S7�B��3s|�B\<9�<d��0%3ד�ZKsBfy�,I���_3���
�b�`K��
�*D&�U]8&F�i�8���}$��y!�q%S� T�D�P���L
me�0W"�XP"�	N~)���C�Vu�LT�!]��؄gX�R6a��
�#�����HnjD����	L�B^08�B����f�~����ݰۛs�|G�@�L��Fxa6�wf۾=�<8�p������9d�bxQ�s�7�Ǡ���)��燧�M8>�R�L��r~��aY}b@�64�) �b�q�@�2_o��,e�y1ӞO���<�	- N��!X���������DԂU�HX���!�AbD��w�Y�~ل�C `Cx2���'�.l�y��Bg�<���ƙ
2\�"���$9˻����Ĥ#��^�#L7��K�iL0�g���X\60i��4�%ូ`�³3�Bȥ�)+C^2K�ʤ,�����Yn�O>�J��xy�H��4��$��dHBxg�0t0�B!6%34e3\Xԉ1�����;�7FE8aA�YRW���P�����|�	~&�6Zy&$�m��1��x�A��xNGskT���P��T�KXSg$<HP�fpy/9�x�F��qcp���ՙ��O�����F�+�o9?|�����-�t�����.���e=!���j�)���O��8h#��X�Þ{��:�r�2�B$H1!���+��3s$͡��{��,^�$k�ɥ�8��2� \�B�1!V	L4��V4H����uO��~?jbB�/���S�3���8~#$%�g7�ɼO@?����U֚� �� �/�R,#X�DB�R�x��q4ND`�"��Ոҥ`0�F$$!# �$X� �P*��R��$Z��8�
0����S9����j���q	d�ל����Ӈ�i�5w|����cI"Ü<xr@��	\t�D8��$��B㤻�4��8�����)��FR�f��A)��4#XHK�7�4��C��!J`o���.f��]��cr��~��j� �`S��ᥗ(Z/�~D�R�s�<9��s9���p����矿~��֑���E�!L�?o������)
B��	BROߥۻ��Bd[�D�8@�~WvS.g�<�̳̗%	9�&���)� �F��M�O'�BSS]#G#I6#%P�p��$�|�3?��c����X-�$y�;.obH���J��k���@+��J��Ȱ��aF[����x~V�iT@������q4:=���B3��:i'����HWăW�n�x��yIXVR|���g�,�����!��Ō�B�,�
B���PŁL=p�pԉP�S>0���!HPă\#Lc	L T V	F%H�LL1�!L��qcXЈD#M80(1i�~��n�x���B�F�HD��H��+"X¸$.B�� ����H�H�0��߬��Zx�B�k`JB�C!/��g��)�4%e	M�<��&Ò~�?��9�?_*VR�3)gvq��&�JJ�bĩ � *a�Ń�)����x�HS�+��� c6j@+.FL0)��8K�cF#p� \�q!LbW�B��`�bP� �e̮$�O�&�K��:����Ka�Ć�b,%p�B��k��H�P�\�$���V�9�.s�)!�j�k(�(F�!4�L�%bBT���8�8�X\l���2B$�B�! D�&���cK�`�� �X	P�T0��F1B�T""�"BFB#\s������DZ" ��2 �# ��YH��C���&:c�a�!l�D���ӻ��~� ��  ����|�p     m�     ��� -����-�$�L�l�`��Hs��  .� �L $ [A       @   m �`6� 6Z�x m ְ -�m�I�8       ��-���)�M���H@   � m�m�����Km�P��
�m�m���[d�-��lt]���h �d��n7i6�6EH[@-�m�ԋh�U*�@�Z��ө��1^��T����,�[C��ZlH���d��lUYF�V��f��%vd�� :�3l��EP��*���T��eB^�8 8��`-�À$�CK��@�n�kQ��p@h�  � p(�h�H���|�]h��ok{[��?>�O��� Ԁ m�В� 8[m���l 	�݈���PN&�vj��\N- ��m�V�     ŵ� ��(�^.�{pܖ�btK.�Wl�x��@m&�lrޫhk�  ��H-�	��p��3-�h��l�ۉ �D��D���u�I��96�9��7m�5���m�Am$  �   [@�n�k��m��� 6�N�in�uQ�i-�yvk���}��U���m�۸ -��	 q �$[d-�Z�j����H6��m��Xi ��А�%��BE�m:	 ��)��S-6�[R[[m H m�  mtk�'I(k������H ͇k�۝m7/�y��JY�#���ճ�1�P�l�n�`	ie�LH���Cm�  ��	���m  -� I���d� $[v݀ nԷ׭6�6�v��f�\[@   $��ۤ�l�R඀�ժ��ںb�궩��s��r���-��]6 lv�v�*���\Ql�#�i���\	��;u�ʮ�d�[�յ�Ŵ�-�+I9�V��a.P8�0>&�ڲ�\ �+/3��Q$�ѶrZl�l�X�� �aiJir�͢P�r�H��`-�F�"�r��.�4P�-�    -�"F�m�m�  %,��Ԩ�b�j��� �m$�`�Sl���Mm�� -�9m�d�J]:��|6�[@kX���I�  �r�s��4�,������f���Zl �j�[@ -� �� p�`  u�t�g�ܻ-J�kb�` �
�gl  �6݀,��L6�P H��rݦ٭��h6�p  ��v�tp @m�l�lr�t��m�Ŵ �m�e��c�ek(�WU�+i�[���Ԓ�m�  �ͳD$�  ��p ��3m 8$$��d�HH�m� ���9����U@!��$G.�x $-�km�	���m�� ����� ��9���b���h	6�\$��X-i"N���	��%^������jӖ;@�FP-�٦���Km��i�Q��i.䀰�ۖ����t�HӶ��n l�vY����� �-�Գ�5� �릚I@:t �$����̒��.A�msk�	UVΞ6%h +69Bp�����j��ݨ8����@m��u��]7����/I,���p[I+ccm&�P6G6ݣ�ڠ�)��͵+��j�!���+�5�Kۚ�%�C�� �K#�Б:�����@��^iv�I�!�m�����XXm�cm��� |    ݻ0s��zQ��#��v�CP�uӢr��E�i�NRP���Mnݴ���p�[�m �hV��ƎQ�Gvp����d�\!�m ���TqG;j�p6N�')ʩ�eA#�2��꧕����k �2�!�;`���m���]�j�κ�W.��&�I�pT��[*�a�M��A&�$�/S��6:yʻ~���-�dX`mZ��`�>���iT8U�����*��;m�ac��n�@N����H��� �^6�(  �4��"tm[ HHM9u�5�r@� &�Ri3��m�ì����  �mm�AZ۷�������ۖ��86� [4�������f�e�H    ��tݠ�I��m�V� �[@Eq��Kh s�+��bc#@+�ꪨp��i����sa�ۤ�  [@&��:��q��u	�.�n�kn�Nm���֎��J[�6�Û��� �+�c!��afd�q�j�X9U	����[SP�v�X`��UG=�B�t�3�-6yY����YC�1�V����g`eez�lk��]��Wf�T���-e` �� ڶ�m����6�W��:m�i2�6v� �e4��4�m%�9��n� 8��6Z٦�   �{��庭�Un�Y6ZM�s` ���@��r�e�      8pm�۰ ᴖ݅�hְ���x6��*�!5J��\� p 6�����I�V�G:۶���Iӵ�m	�  l���[p�    �&B����%����T� 7l�I��c- l� �d�ᑲ���G�W!/C�k2]�Wj�;ev]�<�,�U	Ք���퐃j�e���X�V���.U��&Mhl:�+��m�riy����ؽ
^H��
�J����S�.ܵU rD��m��d���^'kj�vTc�C`F&��X�e� �-����y���
��� ���/K�K(l-�����z���I6  �n���m����$�9���pH�n�[@ 8OUҫ��+jpo^rA�[rڐH'CF� �j�����s�4�Ul�-�  �o0�[��u[�  �J��UUUS�xi&��  �   m$�29ۢ�@�f�@  �m��E7���ͤ�m�q�`�`�V�-��	'%�ev����� m�   ��hV���h���@����Ytk�<  $ֹ��v�[�5�K�U+���)V.�2�SZ�-������Sl��=]p is��\�5;s��%�r�EU����˦ć[]��KXE͝����|]jiZ�Bv��F��ʹ��ޥ��˰��v��P 	���ZU��������$��[B!�5�7n�����d#h䎴��j@8I�m�CnBu����޷E p   [Kkl�Omյ��-)B=���U]ɆjBCns4�@�U^86�z�h ��[��(���  g��7�Um����$�֛l��  X��l���� F�m�l�[�� $I�m,�V��.ݘ+7[vؼ�$�Z��N��t��Իl+1jN 4�� �s`��   m�[=��j��<2D*�UŶSvia	m�����Em��MVa�%�$ m�m�` ����E�D��5�ؖ��.�[��-� H    $�b�nt�#m�i%�iB� k��[.��޷�9� ������ ݧf[�m��m �-�p   �mZY%��[m��m    GJ�v 	H��m���/�5��Im8A $	�m  �  ��z�m�"H [dp�]n$����  *Լ�VյJ�I�p;v��А6�X���ȓr�"ն�  ��    �m� n� 8 �      �  $p -� 6� � �c�@ 8 8  ` ڐ m� A�[E���oJn-� [d�``*�k��iV�Y�hq��   ��m��$  p ����� 6ZH�D�Rf���     ��`6��A�oN]h��ލ�A��}�}� =�zJB�I��%�����d�W��K-,l[*�UP#-R�[��8�-�]�Am�i1��@%��-�Z��#^�m�E$� �M��V��ŲP ���   mi��o\�   �km�ۀo9��� >7�O�W,��  ����Im�e�amh  m � �`�   @ [d� $j�kViE$p m�i�g i��8pl @ m�� �  j�m�Uz�$�����l  � m�^�@ vٶ 	gIK���S��r��R���䖅�q��u�m[@  �h�l �ą�sl�o�ݻxZ[��U+¥��QJ�UU�l�� �2����5�}]��ʫT�@7e��-��]8����ww�ܩ�"��D��#���h?�"���O�x�����$D�?*5�����B����TJ��g�q��"j uT5 �/pG��H�A��> �@P(��]G���W��A��qX�D��9�U|7�@ �����ģ�@D�TS�?�� ~��ő�E'�Π!�A}���� � *)�+����	�*��^���(�8��G�>���=@������01�"X��� ��A0D}�)��A��^��0T �����@��z#�� �"��}DE�U}3����:�AC��T�Tc?'��>#��A:"	�SP#��A?!�pOھ���DC�	ި�b#�QD�	��]x~C�<�DOʑ ��\�/�C��A���!�� ��?�EEtG�?�!:{ޝ���o�|6���m�����o6�- �����^]���v�����zI%�]�td��Gn؜���N�6�n"4����u�T�sv�8{���`ۙ����;�`�t��˳6.0����V�d�ܶ�#B0��ٴ3v�2]��"�J�bL5]-�sѧ�ݎ�yR���!�-ce���8��SrNe�:�xT�x60�����Ry� #2�Ns��=������v[n6�v-�
l.%�t�l�� �UW6
�x⇴����q8'f�ƙ�:"ZYY٘ڮF�9	#��=[���J*/!���Q��r��.jTqF�&LՔ�jk�]	v���� �8y�� ^J�v9�АsY��ç�&��\�Mr�Zq�ݗ.8�U ��l�ƷQ�km�Gӓv���r��[��teZ3*�#�24:N�����s�杵ӂl���OYC���-Z�=RE.3.��g����#�f<m�qՙ�iŢ��O�y!��
]{C�b;m��V���vYUzmPS<��w]1s����p��M��rtRk����l*�-�7+.��U"�/;p�2hC���nɻMU�,Z�.笜��!y��#H��غr�qۜ>�x�n-՞Y���<�R��TU�e5u���=Y5l���wkV3�*u�z�Z�&F����h ��62�z�mƦ���0��܈l-��8��G$�D�nZN�,$s�;	\�Ƭ+�V���]@�rd��y64VkhM�v&����X���K8��P��#M]*��Ŧn���v���djO����ݴ���܋���UUmۣl�� [:�V��<��R�J��͌Tp@C�;N�����,��z,���H�n��l�a�`%6浅���5p�1m�I��
I��T���ś�h
^en�0*�%\��e�IWI���,��۲��V̧>�:����^�72n�7�&�^[���]%�]�@S��=P�FAE��,UH"���NQ�����^*t}�$��|��ݣ��Q�af���p(l�9I�<[�v�&��N�"���xg�f�$�S-�W���:��m�o�&��L�<�:[:�n5���/	+:j4\=�n�.���'���&�s���pta�p��O9ۧ\v��e[������'��/]�l�����֣�����77%ȊqEZ�����lg��4l�5S&Y��K3&�7Kw7j��^i����>�/c'����^��wm��'*�)�&���òbm6����C�Қ���wO�D$�~���7Pj��ܹtQT�I�X�=/�%�d;7����7�)�v*����$�di8h�Y�w*D���f��!�\�-pSQI�~�h�)�{�)����Y��J%�`�$qh�S@��S@/���;V��ҷ��H<M�X�z��k��r�`99#�mϫ�=�D1�:�#�i8�Ȱ�1b��@��S@&l�r�L	�p`b�T��⢓si36rI;���0�D�����f$�T ��AB"$����J�Q2<�ٰ7���=�zX��.�'0�8�@���;V�{�4�.�>4���.�IZ)25$�]U�ծ�$���4�Y��ޤ���$��KW��%݀�J(�k��ԒY��ޤ���$�r�]�IE�
`��������������.�& ܨFx��:��K<]�N�}Q��!a:�:;3���T]%Vf$��󱤒�\��I(���$���OߒK��h�I�`�4��4�]ˑw�%�)�����$�ۖ�$�v���Q,S8H���$��L��߽�g�\QH@��X"����y�;����oߒKϮ��,&LX��pz�Kٮ�I)���Iw.Eޤ�[p��Ix�tq�����,���$�]����\��I(��M$�dp�RK�}�%OWx��:��f��\�)'k�s�k��峻�= �٫�]m��#�= S���o�$�o�]�IE�
i$�#�z�Jlv4�]蒵)2E$�F܎/ߒJ��z�K28w�$��cI%�;Ԓ��W�qG�����$��v��$��v�ٟ;�������$��Vr��0hqA8~��J��jI/zZ�~I+�v^[j�|��$(�*,@�R!E4)��
g-����$�ΣF�L�1�܋RI{.Eޤ�ڸ&�K28w�$�ܴ�I{������w��]!�,\�^-�<�>g\���W�>�����^K�ϳu�2�й��-���n���U�I%���I)�-~���[I{��/ߒK��Z�y&,RF������$���i$��"�RJm\I$�z��o&&,#����I+�a�$��"�RJm\I%���IF#k���8�)!�$�zZ�~I+�QjI/{���$��v�K�V�&H�������ޤ�[p��K�svw�@�O>9'����I?�b����j��(!B����ɦ�QUOl<�j���#��A��'�{�[�� �WcXl�|�Ƌ��N��z9��).t�ťۈ��.R4������s�i�`]�V֕m��9f]�$�K�Nt�����u��un�ݬ���bO+<w��Aꨴ��vҲ�������:w&�p#/��8ڲaB�t��R�A�*2rn�z���x��w;1cgd�,�y��{�X�:a{y��Ɣ֗W\�ҍ�P�h�w0p�.�
���V��[12�l�WZ�~6���T���$��U����''ץ4�v���Z�Қ��(�I�`�4�*�`fK�r�L�p`dۃ+[Tx�K��Hh�j�=�)�z����YM��A��	�)!Ut�̗M���p`j�)����������Qy��v���j��̅/ƶl]�.Rz��m	�n�ӻOIz��j�p���o�����ՒS2�Lx����"i˙	mX��.�#𖇦"h�\QB�[��rI���o$=z�h�kRd�I����4�03%���c��.��qHj(�C�IŠ{�)�z���?z�h�j�;Y�`�Hpbp�=smX	(�������6��K|n�/F���l���CE���S�u�.'[���n5p7N�Yz�;!l`w%���R&elL�H�S��X�4����v���?�3;jy07�ό�0;6:VUp��_��M9�=�͛ۛj̈́�KQ�9)�w��@<z�"k&(,#��02l|`w*D�ܩ2�&�=����18�)3@��j�;�ՠ{�)�z���;���<�x�'
S��yXS��hV:.���*=k�s��^'X��S�I�"�b#rG��v���M׮���ՠ{���E!HpiS��ǥ�P�L��֬ewM����߳./�/�X�,pbp�;�����ՠ�f��t�����7�dXKU2�ՇBIDO��M�nw;����=U�"
~������N���ʜ$pp�C@;����M׮���S@�}\���ӑ��1��M\5��u��t�Tl�uvD��6�@�Hֻ-3��dŊL�ɠ{�)�z���?yڴ�l���5�Ńp�=����%2{+�ls���=,{�]TNa��Q Rf���ՠ�f��t����s@�<Jؤ�$��ܑ�`�[3n�ʑ03+p�B6��94{�4^��?z�f�3ۮ�"D(Q���j�ș%��W7Q�t��綺�8�v(�K���k)'T;�r�&Yxzړh���;�⫮z�G&��mp��q`�����fp���[�؏NQ!��X�N��onr�q�;\��kZ�7��Ս�[���gD$X�ɰ��O3sQi-�ܪX��'[�q�6���c����E�8
�c7+�q�$lB׭���[i��X�������9%ݶe�v�ٗ<�ٛi�t�Q��:E��)���JsѮ��(?���H�M�����_Y�~�hz٠{�)�~����
cJ�*��ܩ ̒��p`fK��[Ty$Pp�Š��@��S@������ՠ~���
dŊ�Uv��ۃ2\ʑ0�-�x�U�K&(,#��{�S@��0�-����M�Z���3C;�q����;t�.M�{u�ym���d�r�ݰ7XǊ!8�sC�$$�~�h�l�=��=zS@�<Jؤ���n��{uݥ��BIE�g���t����ՠ{���E!Hy��f�6���T��nIl⋄�cI�818h�)�~�hz٠{�)�~����
cJ!�ʑ0?s�qM���n���ɷ��{�������9e鷃�N%%��3��gy5�����q]u����鄳��2U�uk�}�`fm���n�H��u�ƅ2`��#rh�Jo�ى���m{ɀnIl�U�._������6Ձ�ջ6yT%�"AH�I(�A�&�!�虤I�(H4B �m �8:P]cP��.B�h�I�$Mz�a K�� �hĊ��.�R���<��b_��)��L1"@�ddj"�1$D�#��2� ��
����
�k����
�����Iy���� 2!�""�߰01@G��@��QF���Bb�?�C�#�@AP�EP��
�X9'?~����Қ��TG0�8�@������nIl͸02m���\JKWvAɁ�8��l�=��=zS@��ݛ��s����̶�*N	+7�ܼ�e����gø�)�c6�ӝงgm��(F�A�'�;���=zS@��)��f�ت�YbLi1�����r\���ۃ�Fz��\�����n������@��S@��M ��^<�&"!�	Z��v��KۏK
Y
1@�	���:"����{�גN���ܹv�4�|���f��K��R&��{o����(��!V����Krr�e�.h�u�I=a3�%��bz�ɤ���,v��ª�vG�r�LrK`fm�@3�B���H��~�hz٠{�)�z���;��#�&�]�Z`�[3n�ʑh�0V�#�0A�&��t����s@���@;��⫁e��i6���V02l|`fT��nIl�rrI��"�ߗ�l�3<�ɻ����?|۷���=�C�y��A�ƞ��,���c�.���t�+c3l;�a����$�.�ӓ�'^w0g�٘+�[�Y��-)�0qN���/T��[u�vMַc]��<qXfk:$q�.�5���.
�h;��v��.GJ]HZ��Ǟ�'��a�l�n���S����k�2��6�n7#��1���9��-/��}��w�����B��quۉE���s�]rI��z5��M�������i>�v�:�de���%��rU3��?|��� ��|�Hfs����o~V��]J�iĦ�i�t��d7;���ϋۏKJ'1�M��κ��,h�6�Sw�2fs����Ɓ�;V�w���ܬ�Y1Aa\*�`dۃ2�LrK`fK� �GVG0�n(�'�v� �[4zˆ��Қ]]s���bN�=�H�nN�z�V�cB�����V,@v藌lV�gHR29��6܎- �[4zˆ��ǧ�_�3+�l����7N]*�I�i��ר�%P�%��zX�[���f�qU����4�C��h�zX�n͜���ɹ���|��wM�)�(��{�ՠ�f��Yp�=zS@-�׏$Ɉ&4�QŠ�f��Yp�=zS@���@�,����Dl�$q
n8ȸ���)���;���b�l���H�R�	"�L�ɠ{�\4^��=�j���@=�ŐK&( �,#�h�)�fT��nIl�s� �p�l���}T�̄�,z�f�3ۮ���@�^�����	B�D?��^���ץ���'�#��ɀ�r8��l�=�.�Jh�h��
�jF�A���k�X�Y�|~2���3ۮ��3�ۿBc����@psȅk��q�Q��ln�΋�Aw����Z�똶:��EYB���7�όʑ0�-��%�@�����2 S����;V�w���e�@��M ��[	2b	������@���h�)�{�S@���	0ń��@����=���=�ݛ�
���v�N�,���8��a�z����YM �[4zˆ��}��ĠI�$��mb�Ks�V{֡p��(����Q�7nMpk�]���$#�7H��;��- �[4zˆ��Қy�uq9���ۗV���̗802m���R&x+pq�%�!�@���h�)�{�ՠ�f�qU��co����B���ɷeH���̗80*���2L��(��{�ՠ��`{������B�!(�Сx����w]�o��C��T�]5X����j�٣FM��ck��lc���+��n�S��fɡ��d�j�>�񛳷���7/->ô�+v��V;X��g\��m���+D^p%'>ݮ���I��>��o(%�B����&ܜ�[��˙�3mGc�M�n4nxƛ����6�.3�Omm��U��;�-���o��H��m�GL���꿷���kw�ׂ��vh�7;�h�l�˗��~7�"�fh�6ϳt1;8J��v�Zf?6���l�s�&��"`E�����m
P�uM���E�$�L�|X�w���.�Y1CG�M�03*D�7$�d���s��u�9��qD�8h�hz٠{�\4^��;��"s�91�%Z`�[2\��ɷeH����d��:L���S�Ħ�H�ㄔl>Nh����e�<��f��M%:f��{r.[2\��ɷeH����Rp�:�*J��Q4�`{q�j!+HP��&�)�0F(d��R�z�����s�:/ju0��`fK�DlWwi�L�	L�=�ݛ �n�:"!)���h��mT�#y1��nl75���E���KJ�>�:w�����hR�Ӛn����,������6���ڜ�ܸ��i�F�p���N�sg�D.�����ip��M68��x�1���1dqa�@�Қ�e4�Y�{�\48�s�Na��Q �e��k��%2�����Ȱ3q�w�%�D��cn) ��h��E���B��u�`~��,x('tJF�A�&��Yp�:����YM ��h\,V6���819���n�p`6[2\���sn^�M<�$a�ݠ�S8�:�
3�f�s`�:�1lf�n��=UaF�Ӗ��p`6[2\��ٷ$Yc�9�I�#R׬�=�.^��=�)�U����,2L�ݰ3%��p`fK� ٲ�bẅ�1AǄs�Jh���$���y&�r ��J��R���
U�� *T�fwΓ�I����G0�n(�'޲���~����}��ץ4���"O$��3jP݆y#�O0�my�Ղ\u��-��X���H�)$n)'�m8�4�Y�{�\6�����`n����t$� ۓ@���hzS@����u�4��+��Ӄ�hzS@���gDL������Ȱ7*p֛�%�q%���@����u�4zˆ��ӽ�ŀwt�t��ؚ��n���3s]��Q�|��ok�����`J��<"b�G�����H���ԒB13F0"��$�@8 8n��TM��1"$Y�&��)
�	.$`@�q�d$�V6B1���&,@"Eb1 ��,����LH�08@�H��B	#��F$H�����cG"���GXVHH&���$�B@�D}_!9���T8��F0Z��@�*1(D�)
J(F����<��1�����'��p�x�� �
HH���	OI!%�����HLx����M�	��$`G�4|B0���HC���%����o�xЗ %1%0�!,�4t�2I	�B$%�T�5H��D�]Ѕ+�x$!�N�=R����i��"q�$���Q!1�<�0$&�ܞ��dB�
���DX�dXDЁ!1�L X@�HP�H���s%��$�RRT�b�bDHH�#0P�c"!X�%HUcB-$�d�1���(�"R�(�����������}�~�&�n��m$x[��v6��
 Uvg*T���M@c�3�n�t۞��p��{e�{��j��ܩl��ݼ�g��m�ٲ�(�����a����Ot2@+g8	��{p�y_N�V�I@���]R�/:8�)��tGh�h)�����i��^��y�������`N�qtcJ��;�ݐ�:���c4˘�j�������%�&;:V.�����1��6�{v�8ݡ�n�y:ժ�͉�����mY�tnҞ�e�ƙܩ\h��L�#5�krd��,u��rG`�#I���3I���\'j� �����3Z�Gl�$n{�D�(p�r��^W��:����j�+tpŞ���n��;t�8:��h�,��ohQܹ@�2.20���� _U[��е�x�W�#@�9.��vm�p9�����r�&@��3����ҧ�!����e�;v�h�5v��3�n��gt�/E;4�����ܜu[�8p�UX����=vd@ܱ/l��C�~�,�m�]�,�N�t�2�-��`m���Vne��5M���j�V�C����K3i����x*�N�\��w�>���O�q;&�wBBqƴ:x.��[[g�K=Bɶ��5�y|9w�Vѳ[a�L�������V������clU��a���N��U^�  '9W�7C��2!�b{;hN	�[nh4RM�i�6�Lt�6�V%)��]�'�eʱ��x�y�6��t�^/=�m�R�N���J�3;a�Iĭ�:��L���h��z��0�U���p��JŞֵif thL���ζv�ȣ�UU^�q�T���
:e�
�Fv�V�٣����RID;�N7CG�-���I@��!�cjI;�����&��7^�� 9%ڨ�,����c���{b�[m*�e\�Ԡ�uP;�Km�E8I�i̎�u��O7f����."R��K�N�Uy�UK�������{�߿= �S�T�@���T7�?�⠞z-�I�{�v�d�s.�˒�U�F���Dl��p h�e�N�ٶ�\;��@�Pi.�D�������lU��lP�����n���p��v�u��g�۷'V뉝�>�\��s�qp�N^"�6핳\�$��}���ۖ�x�:����`;r;�wg�4G^ݫ��t�V��7	�ӹ]Z]��gQe�g���%)q�-�烛�7j�n)�t���W �M���㣆�݂^�'$Л��Г�v�Ȼ����k�Ysŵv6��ց���͸03%��l�l1iTj�ԱK)�4X����'Tfs��7�]��k�X��5��DU9��U��p`6[=�����zO���+dn)'�m8�4�Y�{�\4�)�{�S@����$QF4�A�&��Yp�?gU)�{�S@:���AJ���#q���Hq�=d6�Tu8�G2��ha99#0�r��m�8��c��@�Қ�e4�Y��~A����:��#dm�%��@�����/� �������o;w"��ǥ��d;�xt�RpȚd�8��~��e�O�u���e4�:��@��I�94z�E���K�ץ�(P�w���fN��bɊ8��a�u�M޲�׬�=�.����x�br(���I룭t�I���׎���^��G�cv��ns���'H���YM ��h�����Kޠ�o�g=�UN%�U4���6l�d����n�p~���H��Em!�rh�O��3q�f-Q�C{�����S���n�&���D�E�BQ��Ł�ύ ��h~��.�gW1�Fډ,�n�� ��4�ˆ�ץ47����Ø��zw��`΄�gl��9��$�3 ��9X}1OW6���]�f�`fK�6��̗�lx�I�L�ɠ{�\4�)�{�S@:���ܛ�Y1B��_͸03%���|��;`fK�hq��2'0�N(�'޲����{^�(���"�%!:�{�`l�'���Ķ⪦��0�-��.p`l����.�_��]�F�e9�۝1��^J��b�nM3�|͔V͸�tgx.!��[�(g��|d�����&eH���dv��Up�co�61���4��߳�?�;��- �_���Yp�/5�\��j$�18�yڴ�Y�{�\4���j���LI�$qh^�@���,�͛��>�;y�U��h�Ni��ר�>I/�}}�������`dD,�5WT�L�(d�'n��ܐO�w��ҥ��Ց{;���x(:ȇ�;v]����X�q[���ųlh�"���b�������yvP�`����V���^gs��i`:������8�ݠ�J���q�z4��u�U۵�;��gg\�A�֥̽.�\H�Ջtn]f���W��Ӥ�ڲ��88�L��T�{y�v����K�7s �)��@G�˙�7.�7e�e�7wB��.�3t�ɛ[-�D�]�`B�ƙ֩5B;Xj9�d����9������yڴ75�~���Ȱ�-�MT�̅U�eH���OO[w����09{km����i�#�@:���e�@����v��
Є�m!�rh����h�h[f�qU�����lc��h]�@���@:�4zˆ��u؛Ș�S'n'+T�:��D�=F�m�̫{_�����=1\\L�,��m��K#���u�h����h꬙&8E��6�9���~P�BP��(r?k�X�[�`{ջ7�$�)���uQJX6�(�"rh�O��:�V��;V�u�h�r�bY1B490�a�uv�ޭٰ��aДNg_"�4żӖ��Q�r-�v� �l�=�.Wj�*���2c��?�"��� �5ck���V�.l]V�7���c��Ga�o?�i�����޲�uv��v�����Q��A�&��Yp�:�V��;V�u�h\,m�*��V!U�`l�2�L,�⍗f����U�9ٍ"6�Idb�h�ǹf��ר���]��������mS��j�n��n�9(�ξG�7��lz�f���S��M��^�S����t�2�`99�*/;GQ�!�%��dG(a�	2'&��Yp�:����n�BQ���`f�SS)�M��4X��7�Q&ewM�ow;�ר��	DL����r�))Ժ��s`fWt�nk��"!L�s�Xս6O�w]U8�nUUM7Nl>J>J*�����?�`f�l�$�Q	-I*��.���~�;��w���uS%&USl�s�elLʑ0�-���s�������\�p�;&l�V8 �	���)��MO]w7���4Z���w{�>��|(��$�G�﫾�ޭٰ��пHw}>�@�U����j$��n-�{�}2�����Ȱ3k6o�C���M�c���Smӛ ��v��Qg�(��J���@�|��:��@�XI�94zˆ���Z��Z׬����1,��G�Ƀs���s��������,�JJ�������Z�gvZ��5{4Ցk2@���������V�+��v��`��6\����7V��sq��@'n�k��u��]�a֭j���̻	7S�������)��z4h���u�df���F;�<����u�v���{\��v9� �0�C�U�v붝qs�k����Zg��c��G�Ё��Q�fe6Ͷ]�.���~3|���74j�3lv�.K��ۆ��T�Xĳ�2m��Z�F��bū���2K���o��z&�e��9l��05`).����r8��Y��nM��y�Zw`ԎF���4�'-���&elLf�`N(�X��M��Lnd��+��-�ߖ�u�4?ᙉ{��&��*&�IaUi��[ ٲ�rN[elLﻻ��������x)��K�Db��qh�¤ά?���ؚ�m��n��'g)WW6�53T�t���|���S�3k6ly�Z�x�$�dNM�����h(@�Iy���'����@:����; �LX�Ƥ�Zؘ��3�'�������i/��C�F���y�Z׬�?zˆ���ZY�V���Jm�#�@6l��|�àOT�`fV��ͥ��BY^�%y�Wz�`:57=�t���m���^�-Σ����z��{���kc�%4㞲���s�X��6�Y���>����򟧂WΪ�j�42f�,�͛2�&�e�;�����Qr*�(���(���;��h]k��0���}X0�X�0�JRE�$) 1d��hJ�����H�HF��M�T�*��N1��z8�T��h0"DH@�<��4H!��/�����
�H`�X����'�`u�3\�IiD�h4q�D�A��V��P��9L�HB1�`���"z���	�wMN
)@E"��QD��T S@��q_A�z�"�?*1q�dD.P�W~�Ȱ7k�l3gi��c�䚖ۧ6�����"HRBß���Kı?{���yı,O}��Ȗ%�bw��;�a6M�-&훛�O"X�%��wzLND�,K�����^'�%�bw�~�9ı,O��{�O"X�%���~�����sw.�Wk�0n�yg�"����[,x/MԺ̴N�W�v����~~�q��V�v}߽�7������x�D�,K�n�T�Kı?g��p?��ı=�o���Kı/��i�vB�ܻ�&f�'�,K��۽�9ı,O��{�O"X�%��wzLND�,K����'�,K���;����6feͻ��"X�%��=�s��KİwzMND��XdL��w�Ȗ%�bw�x�VB������a:ʖ�%Rn^�q<�bX���I�Ȗ%�b~�{���%�bX��w��"X������Ȗ%�b~3��Sw3��m����Kı?{���yı,O}��S�,K�������%�bQG��+!I
HRB��C�xm�����<����[۳v�#8I�Z��^��3d1`�sp7N݃������r������{��7���ҧ"X�%��=�s��KİwzMND�,K����'�,K����ɛ3f��L˻�vT�Kı?g��q<�bX���I�Ȗ%�b~�{���%�bX��w��"X�%���[J�	�7#�W�
HRB�G��I�Ȗ%�b~�{���%�bX��w��"X�%��=�s��Kı)?{��-4��	wI����KϒD������%�bX��ߥND�,K�{��Ȗ%�`������bX�!O�Y�9l$M�ꂩ���B��X��w��"X�%��w�}�O�,K�������bX�'�w��O"X�%��� *�E�	���L��B@"�$��L���:��
j׆�*Q���q۪4���ۥu�h4wE�X�n���81�Q��8KmY��ҽ�0�+�ď����yv�8y:vNY�����\�\:�c���k۳t�]�m֮<,p�k]=�i<�����8�+t #9�q��W=GQe�$����%��{T�m�id��A���޳b�is�$�ԑ���ܲ曹�}�S��%��.lۖ��UWMm�[)�@�����ub��9:r;HY!��GF�K�k*1X�~����{�Os���O"X�%����jr%�bX�����<�bX�'���Ȗ%�b{ﳔ���w7rSۻ���%�bX?��&�"X�%����oȖ%�b{��ʜ�bX�'����'�,K�靧Jn�cs!rm�4���bX�'�w��O"X�%��{*r%�bX����8�D�,K�w���Kı=����ܓne�rMɛ���Kı=��eND�,K���x�D�,K�w���K��&D������%�oq�ߟ���h�p���w��oqľ���'�,K���ω��Kı;����yı,O}��S�,��ow��ːx�U�<���-�v{y�Iz��:u�m�{s���\E�,��v�-&�wx�D�,K�w���Kı=�����Kı=��e��2%�b^�����%�bX�����2�\ۄ����jr%�bX��{����| �!l@�T`���"~�b{w�S�,KĿ������KİwzMND�,K��{�6饆�M̓sx�D�,K�n�T�Kı/��w��K� ���MND�,K�}��O"X�%��=�3��[v�nmݕ9Ĳ���� ����j(A٘�X�]�f��VB�������'�i���2�7x�D�,K�w���Kı=�{�Ȗ%�b{��ʜ�bX�%����<�bX�'}���m�t��v�䇱��U��'e�]�5�=�IYN�7*gF'Q��݋��y7.72&�sI��Kı;��y��%�bX��w��"X�%�}�{��~��,K߷�jr%�bX�giۓ�ne�rMɹ�O"X�%��{*r%�bX������%�bX?��&�"X�%��{�8�D����w�?��uuh�r��w��oq��%��}�O"X�%����jr%��F"�U���H0���*��|,M��o�^'�,K���J��bX�'w��3��KI�m��'�,K����59ı,O{���<�bX�'���Ȗ%��ș߻��<�bX�%'��t܆�v�3t��MND�,K�ｼO"X�%��${�ϥO"X�%�{�~�'�,K����59ı,K��=�ͳ�[�]�1u�tc��\Et�Oל��#�61�v��n^]r���.�{�[�o%��{*r%�bX�����yı,�ޓC�� o�ı>�߿�=߭�7���{��L��ا��'"X�%�}��'��@#�2%����59ı,N����<�bX�'���Ȗ%�b{Ｔ�����nZa�37x�D�,K�w���Kı=�����%��,2&D�n�*r%�bX��w��yı,N��t��f72&�sI�Ȗ%��������^'�,K���ҧ"X�%�}��'�,KS�@T�����y�jr%�bX�����zM��f䛓3oȖ%�b{��ʜ�bX�����x��X�%����59ı,O{���<�bX�'�{�ۓ!����9����9�-�{su�J��vխ�ـu���R�����}�����G���SȖ%�b^�߷��Kı?N�I�Ȗ%�b{�����Kı=��eND�,K����3��KI�m��'�,K��;�&'!��/�"�؛���~��O"X�%����ND�,K��{�O"|�.TȖ%&o6�	�ni�U4T+!I
HRB���x�D�,K�n�T�Kı/�����%�bX��w���Kı/���vm�Kܛ�&f�'�,K>VD�o>�9ı,K߻��<�bX�'���19İ>@dN���x�D�,K�'LϷ4�.��sn�Ȗ%�b_{�w��Kİ�H�>����%�bX��{��yı,O}��S�,K���?s�vssvj&II˴��ht�����Q������=iƩ���1��pD�J�+mn��Ey��]�XκY�-��nM�˞.9���S`$��5v,���n�`$&��V�z�1u�l�p��õƣ��mY�f�m�z�p�u.+�[n�vw�63�-�ֵ�]�9�d���M1b�,��T���1E� B�5�mp]e��H�=��w��|���j�$,��,G���0i�[�L�s����^,I�7;����w����p_!S!�-~{�{�oq���}����Kı=�����%�bX��w��"X�%�}��'�,K�靧l����2\�-�&'"X�%��w��'���J�M�b}���S�,KĿ}��O"X�%��wzLND�P2�D�>�ӷ%������7&f�'�,K��n�*r%�bX�����yı,Oӻ�br%�bX��}��yı,{w;7Mٴ����˻*r%�gʰ2&w���O"X�%���~&'"X�%��w��'�,K��K�>���*r%�bX��s?��6�M-&�wx�D�,K������bX�'��{x�D�,K�n�T�Kı/�����%�bX���o�&Iʓ��%n�ɞ]]l�8��v�X5���5�����v��F��]�6L�&'�,K���߯Ȗ%�b{��ʜ�bX�%���x!?DȖ%���~&'"X�%�{=;�M�kfn]̓3oȖ%�b{��ʜ�'��1qؖ%�w}��<�bX�'���19ı,O{���<���L�b}�����%�7&\ۻ*r%�bX��w��yı,Oӻ�br%�bX��}��yı,O}��S�,K���m-�r����L�e���yı,Oӻ�br%�bX��}��yı,O}��S�,K�3�w��yı,O���Rn��2d�6[�LND�,K�ｼO"X�%��{*r%�bX�����yı,Oӻ�br!�������??P���օ�s9���'k�vM�ɩ����[s%��V����F����|����d�rMə���ı,N��ҧ"X�%�}��'�,K��;�&'"X�%��w��'�,K���s�tݛK�.]ܻ��"X�%�}��'�,K��;�&'"X�%��w��'�,K��۽�9ı,N��e;�m&ZM�n��<�bX�'���19ı,O{���<�c�#! �b�G�,M����Ȗ%�b_;�w��Kı)?{���MKt�SaT�P��$)8J�[׽<O"X�%����T�Kı/�����%�` ̉����,KĽ��Ϧ�5�773$����Kı=��eND�,K��{�O"X�%��wzLND�,K�ｼO"X�%���ɼN�tW�&ݒ�۞��m�^b�V��hx�5����QXv�u�g���N��weO"X�%�{�~�'�,K��;�&'"X�%��w��'�,K��%�0��$)!I��S-��d����O"X�%��wzLNC�9"X��{��yı,N��ҧ"X�%�}��'�,K�靧i7ncp�rl�4���bX�'��{x�D�,K�n�T�Kı/�����%�bX��w���Kı;����zM��v囓3oȖ%��"w��J��bX�%���x�D�,K������bX�� �@�MS��s���<�bX������m.�wr�ʜ�bX�%���x�D�,K�U��y�1?D�,K�����<�bX�'���Ȗ%�b~����2\=:T7	�ڎ�u�hDݷV�:9�kG\�E�-�[�v�˞��\����߭�ı,OӻىȖ%�b{�����Kı=��e�y"X�%���x�D�,K����7!���ݓ3f'"X�%��w��'��?���ؖ'�]��9ı,K������%�bX��w��?�*dK�zw>�t��773$����Kı;ۿJ��bX�%���x�D���DȞϷ�Ȗ%�bw��׉�Kı;�ze��%��.\ۻ*r%�g�*@ș߻��<�bX�'���br%�bX��}��yİ?�FdN���S�,K����T�m�H�5M�/�)!I
H_�w��,K����oȖ%�b{��ʜ�bX�%���x�D�,K�D�ԕ�4�Uc3�#cd������B$d�!��=@�EW������`5R.&�P�t�HM N��� D�@x-�
`h�������J$b@/�a��$W�OOH�~DD8�`H� �F{<``�n�(�"���swI6퀛\[vZp[a'9�cj�`��u��)�*�J�F؉]��6�Y�������sZ��(8�u�.\n�B��6�*6��^,�r<�P���m��7�Q�Nh�/dM��v��
ו�q�ے��G��6��"�i3V�Ԩmo]�٩c�B�Y�2t�oj�<g$ƹ�%�{��n��Ky7`W�n��D�.	�*Ν�$ɳ�C]Z�$m�\��ik�k���p*�F���6�y�H�!i�vJ�qu��
��B#g�i"[3�lź����;wQ͞V��
e�//���+gcbj��oe�<�k��:Q���É)�����q��C���:f����qd��׬ձ���_#c��J�x�y�w\�Ⱥ�q�j�nʹd�ll�����
j�����e܆�j�s]�:�-�]�Y���F�n)ٰS1/�s��gj�8���l��T:�uc�.��8�Vӧg����v"��Ų�vm����Ul� f˔{{m��n�n�'u�E2v�֚u���8d�ڢ���͞i;U��a���t�՛EU��.k΋q{+U'�oR��z#	���
��j#�K�ю��m�ۥ-��Y8]���G�!@�Uv�ltOYu���'��es�+ļ5��М�c��z,lQ��ء�^�;-R�������nm *��^k���v�� �x�.K�ڈ�Q��[��M���� B��ɞ{<O��JN�`��v6�^5�t�hv�s-�6$^�R�Af���!ֶ����q+�����[8��8�i�.���Y�kR��"����U�UlYx�;2�]cY��RJY]�v`r�L쪵u��Y]�8:� r��R�� ۉ	کVB@6�C�v�,I�`)�ح���'d�k%�%]�1���%ԫSn]��k�52� ԠGTڃ����Զ�`���e�N���;3,<�ݺ�Q��i����L�M�sws6�@S�( V��+�{�=T �z�4�*��u��x�Q���3=�ɻ���C34���v���*��4���]Ͷ�m[�dx�qV��.��ؽu�Nm���ŶDFp�7,i���k��z�A�VU��,�N�y'��c���Y���2eO7s�v�x�T�d��C��Q��v� ����`AvM��"�V�nVn��קq9\z��#��xV�FN�h-ӌ��H[zS��i��gV��Ӻ5��r�j؊�]����7��vL�v�v,n���rf.�G=��5;Vλ��7M�i;��ww��;�оq�m��SȖ%�b}�����%�bX��w��"X�%�}��¨O�2%�`���59ı,O���d�s2].Y�36�<�bX�'���Ȗ%�b_{�w��Kİw{59ı,O{���<���L�`���n�K�3.���S�,KĽ��oȖ%�`���jr%�bX��}��yı,O}��S�,K���[;��0�Y7M����%�g�02�s�Ȗ%�bw��׉�Kı=��eND�,��;�~�'�,KĤ��f��ivn7I��S�,K����oȖ%�b{��ʜ�bX�%���x�D�,K�w�S�,K������O��:m��kf��]H�N�n�\uKŌK])%��7t<pF:R������w�]\L����\��=�bX�'�]��9ı,K�}��<�bX���f�"X�%��w��'�,K��OK���d�fܹsn�Ȗ%�b_{�w��?U�x
�U�q�L�`���jr%�bX����x�D�,K�n�T�K����	ݩt�UDԌ������K�w�S�,K����oȖ?$2&D�n�*r%�bX��w��yı,N��v�6�n.M���ND�,�D���׉�Kı;ۿJ��bX�%���x�D�,�}��MND�,K��;�/��̗s)w&f�'�,K��۽�9ı,>#���o�Kİ}�~���bX�'��{x�D�,K��w9���3۹�]�൲���V�WQ"��ɱR�t�[l�cU�n�<���*+ﷸ��{��?���ˉ�Kİw{59ı,O{���?�T���ؖ%����ND�,JB���%}I�Rh�m9m�/�)!I
`���jr%�bX��}��yı,O}��S�,Kľ���Ȗ%�bR~���r]ۄ��fl��Kı=�����%�bX��w��"X��� jX$��:�,L�{�{�O"X�%��٩ȖB���,ֆ�TP麠�sp��K?�?�ﯟҧ"X�%�~���x�D�,K�w�S�,K����oȖ%�bw'����2K3n\��vT�Kı/�����%�bX}߹���%�bX��{��yı,O}��S�,K����zKv��e�m�w\������X���Þ�g�k�uRɻH�s8i�6�i*�ۻ���.f�Ȗ%�`���jr%�bX��}��yı,O}��C��L�bX��w��yı,O���Rfܭ�%ɶ�٩Ȗ%�b{�����Kı=��eND�,K��{�O"X�%���٩ȟ�TȖ'��w2_���.��w&f�'�,K��n�*r%�bX�����y���)�6��jr%�bX�o�׉�Kİ}�ܽ�.�.�̻�weND�,K��{�O"X�%���٩Ȗ%�b{�����K����"�x'�'���"}����Ȗ%�bw�/��i��n�ww��Kİw{59ı,O{���<�bX�'���r%�bX�����yı,O�>�}�9Zs�C��f���4g��aj�gU j$�h��C��zhN����e٩�%�bX�o�׉�Kı?L���,Kľ���Ȗ%�`��z8VB����8yeh6����PU;��%�bX��{ۉ�
�-v&ı/��oȖ%�`������bX�'��{x�D�,K�=.N�i�Y�r�ٛ��,Kľ���Ȗ%�`��{59��Dȝ�{��yı,Ofw�Ȗ%�b~�m����������n�<�bX��w�S�,K����oȖ%�b~��n'"X��L����oȖ%�btϩ�&m��2\�m͚��bX�'��{x�D�,K��{q9ı,K�}��<�bX��w�S�,KĂ�S���w{w����	e��U*�MV'�T^�g�g�ހM�����c�Ʈӳ��kN�ɺ�8�]�/b�];�%ӫ8��8����˅D��E�|�\)q<�ϛng���1[#��ù=Tv�h�7�%�˅��zd-GX
��$��{nE���2�6�ۇ�!t��9V�YN��,��׎��E��{ETQLnG����{�~�{����$��k]7M4�GH�Y�:c^F�N-(�5؛��k��@7.�O%ٗ7(NX�'�,K�������bX�%���x�D�,K��١��ʷ�M�bX����~!I
HR(�_S�M�uU4���Ȗ%�b_{�w��?�@�DȖ�ߦ�"X�%�߷�^'�,K��=�19�ʙ���s%�a�M4�7M����%�bX>�~���bX�'����O"X�b؟����I�����I�}̖�S)s	s`�|"0>�߻�Ӊ�Kı=�����bX�%���x�D�,K��٪����$)��+A��T�T�i��,K��=�19ı,> 9߻��?D�,K���S�,K�����Kı;��!��rfY��ݒ��+h�v���R�o�ؓ�#�m:��]tk����KL�r���ND�,K��{�O"X�%������Kı=����"�_blK�������c��������S�I�k�w�{��%������"�DF�%�b{�y���%�bX��{ۉȖ%�b_{�w��O�2�D�:g���6�0˙�6ۛ59ı,N����<�bX�'���r%�bX�����yı,��f�"X�%��v�ᗤ�̙�2]ə���KτP dOf��Ȗ%�b^�߷��Kİ{����bX�'��{x�D�,K�˽��7i���7&n�ND�,K��{�O"X�%��(����jyı,N����<�bX�'���r%�bX�����ʡOU�=M���L��Ξi��ר�e��ܖd`�2\rˋ=]��q�ѻ�O"X�%������Kı=�����%�bX��{ہ��șı/~����%�bX����nܦ��ist��59ı,O{���<��G"dKٝ��r%�bX��w��yı,��f�"|���+��ĿN�g�ۦ�)���&f�'�,K��Ͽ�'"X�%�}��'�,}E?��OG��|�`���jr%�bX��o~�O"X�%�ܞ�&w4��&�˳7n'"X������oȖ%�`���jr%�bX��}��yİ?�D�o~���bX�'������SM��n�~!I
HR(�=r%�bX"����׉�%�bX�����,Kľ���Ȗ%�b?��c�38�����0��y�vzu�C8��sp�:dd4�;f�od���#ȫ[.l��Kı=�����%�bX��{ۉȖ%�b_{�w��O�2%�`���jr%�bX�wi�2�L�ɚf[�36�<�bX�'���r�G"dK����O"X�%��w�Ȗ%�b{�����O��wg�������h�QӚw��oq��%�����yı,��f�"X�%��w��'�,K��3��ND�,K���/f��HStۻ�O"X�|��2���S�,K���߯Ȗ%�b~��n'"X�DP0 ["gw��Ȗ%�bR~�sv�7fl��nl��Kı=�����%�bX|�1�o~��D�,K����O"X�%������Kı/����6��n�bol\ӬvX�<&눮���݋�����[��|��]	�˲������oq��{q9ı,K�}��<�bX��w�C�P'�2%�bw��׉�K�����9���=Hh}�oq�ı/�����%�bX?���ND�,K�ｼO"X�%��g�����"?��n&ı;ݶ�e�ͳ76L˛����yı,���S�,K����oȖ%�b~��n'"X�%�}��'�,K���Ӵ��)�\�Ͷ\٩Ȗ%�*	"w�w���%�bX�����,Kľ���Ȗ%���2���S�,K���N�K�.�Lܙ.�����%�bX��{ۉȖ%�a�)���w�￷��Kİ{��MND�,K�ｼO"X�%��� ���	�I�y�:g�"��c8D�Z��m"�:�}��s��*�a������v�\b�v�͸��-=�!�N�s�v&��;=n�c(r\���uF������{0��Y��;c���u�잛T�I�I���u�L���]�"�m��ccm����:�F�7bԫ�q��s',�Q���D�ԽIgGv՛����u�0ti�qOS
���Q9�mɺ]�w0�Mܔ�ɍsnNu�rgh��U�eD�f��tK�.�)���]̹7&n�O"X�%�~�߷��Kİ{����bX�'��{x�+?DȖ%����q9ı,O��2߮��KI�m��'�,K����jrʃ��,N����<�bX�'�;���Kı/�����'�(�U��(��njhj��ht�
�RAbX��{��yı,O�=���Kı/�����%�bX?���ND�,K�{=3;6�7�ܓ3oȖ%�b~��n'"X�%�}��'�,K����jr%�`|
L�߹߯Ȗ%�b}�����$���n�ݸ��bX�%���x�D�,K��٩Ȗ%�b{�����Kı?L����7�����~~-&�̚x9��[�#��P�z�&���#9 ��A�s�.!���w�|i.������x�$)!H�5��r%�bX��}��yı,O�=���Kı/�����%�bX���v�v\�e���e͚��bX�'��{x�B�P�(�@�0�P�P�B6&ı=�߮'"X�%�}߷��Kİ{�������S"X�gi���K��7&K�36�<�bX�'�;���Kı/�����%��$2&A�����Kı;�����%�bX>�w/7ͥ�˓rf���Kı/�����%�bX?���ND�,K�ｼO"X����v'g>����bX�'�������HStۻ�O"X�%������Kİ��~�~�O�,K��g~���bX�%���x�D�,K����²[ؓ!�6�nv��U�N��
v�E��j�YM��w��|Ў��5]�f��,K���߯Ȗ%�b~��n'"X�%�}��'�,K����p��$)!IՆ*��i�:UM�U;��%�bX��{ۉ�|�"dK����O"X�%��w�Ȗ%�b{�����Kı;��L��$���n�ݸ��bX�%���x�D�,K��٩Ȗ>�A<U�� 1"1"��&�`G q`B0 2�$�c)44(]#�}:�!~Sا�=0F0�#=�=���S�a�x�GO���4�pB0V$uU=�B�Oԩz���F<^ ��]��B\�:)�(��$`����a������E#�({���#�}DzQC����M��~�O"X�%���{q9ı,Oߦ�ܽ�.��iw6f��Ȗ%����߼����bX�'�����yı,O�=���Kı/�����%�bX��i�M�ssv]�6d��S�,K����oȖ%�a�
��^�}�q?D�,K�����<�bX�{����$O����*NhleK���:�ÄM�i�`*N��nr����ٶ���j�k���F�Lls�Cq~�ߖ�u�,�=>��ս6oSn���K��.��Lf�`nm����&elO�)���L�Ҧ52�Ӗ݁���+���Z׬��Z�M�c���:e�D�=�=ս6���?BM,����h�$�}��I?_��o,&D���`�Z��� ��h�zX��6�Q��N%Ӓ�1M�u�7m��c��z��ڱ��`�s^{<%<�����VR�趂f)�2�n|�w���c����Z����+U�N(5�89$�;�)�bE�ߖ���h^�����2d���s&�72�i�M2�ީ��쭉��'���6_�Z��\S���Z��tU9��!D(�sޛ ��vf=,>�;�zl�:��'IʗU4:)����`}�Q����7�zl۝���U}���B]ϳ�t�&˦�nt�n�m��ql,l]�L�4�7D];�{H	D�u��Ф��9�4A�����OgV�q�l���vY�3�ۮ�C�1���\�R��g��ќ���˺��b.#m��/F���ؤ�\�v|jا�e%8����V�N�b8�����e�C�����'�X��ZEwsy�5�j��&#�)��q�{����W8k����g�]q��-�O'ltsd֎/]�+e�F���hg�����͵��������elLʑ0�-�srJdmAd�"p�:��@�]�@;s]���K�}
���R��9�J��
�L�_�&�e�7v���[��%m�MT:*YM͇B����`n��u}V���V�{�U��)I`��vf=,J�ޟ�{��l�Y�[��c��q�xԉ����n�=6��#��V�4k�3�hX��T=1�ڷRAc���u}V���V�u�?�����|h*����#lQ#�I<�w��QB��D �?��>�~��>4���-�ő�X�m㢛� ��v{�t(�S;ս6�ߖ�zƫO"&$dNM��4�͛����rQ;���7'��.A�L��4�6�f��G��O���4��<��')?�(�Ԏi�^�����W�h�xmy;���JYy,��)�8�7���V�u�4��B�K��oM���2r�h*�,���7$���+b`vT���}�bAܒ�?��"�,#�rM�>4'�罼�����""�~�w��I��������b�r�%RtM2Ò���9�M������!D)��������/�Q��cQŠ~�ՠ�f���K�Y�`rK�]ߜL�ES�E`��#����$TH�����Z��\�`ۛ��n����B*�*ܧIʗUT������4��=_U�~�ՠ^����	#R�6�Svf=/�DD)�:����Wt�{u������iːj��MӚe��[�`~�ݛ>��	L�����gƁˎc�O"j�����ڬ=���zXz"�D$�HP��	 ��(�@^
}���I��l��h*�2�����{u�DD%����;�~Z��Z�}A8&��E'�ywv���=��$��V�kdz�W-�r�=v�0��1pnI�wt����Z�ퟢB_BI/P�|���t��)�.�,yN����Z޶h�_�9D%Tt���R���!Jj��������Ɓ�v���ő�X�i�E����Қ��h}�	O��M��Χ�i�r5*Si�7`g����R&elLvK`>}�}�p�"@�	F���t6�T�sM�幔*�]uVT�{k\]�ӵ��l��sme����s]����Lk� �����ٌJ��`e=��"��]t���	m��	p64d�u�&���zgGttbK�$#A�m�6J^b2B��y�&T�bCL�v�q4�۞���s�T�������7L�s��[g��v�d�V�KM��J��n0k<=������a�T��ھ��&r֯�ʑ��n����5T	���EsS���������M�z��a�������LvK`n����M����MA�9���V�w[4��=]�~H�hG���$�1(��Z����zY�(�9��6����?y%S�bqF ��4>����mߍ}^�`vT��n�lQsW	gZ�bǑ��@�v��v� �h�)�_+��GILbdY��6ձZ�z�*p�g�z�4�^��[�էo��^>��1�D9�=�������4Wj�-�cز<�M2Aȴ��(���Q0��RX��=��6�@������"bA&F��;�S@�R&~�,�{ɀI�[ ܕ/���	MӚe�(J�>�=��6��4��9q�t#����l�@� ݒ��p`d�4��9b�e�T��ۖ�$�Q��Mv���V7#>9��J�X�Ӟ��f�ۂ,����%�7v���R&eH�q$J�jiˢA�*�vf=/�IL���6�|��٠yU�����bǑ�6rI����I<�w���/�@��(�A��(b0F)Q�C�$����x�/�`{�Ł����N�]QMQR����>��6����zX�ՠ[jǱdpA� �Zٺ�J�Gw~���}����f������䫪���І�>N�t�ɱuW�	�f�@1����RG��\q�����ۃ%H��"����	=�`�L�����N��o�#�?�� ��vf=/�$�)�gM��'I�Y���h�����f���J�>4����=�P��&�$���hf�31�`{kvl!%J�����R�DGB��>�ٙ:�Z�婙2����p`d���LvK`f��?A���jv6�������z��ۇ2�a���!�s�b��'Gj�17�᱁��Lʑ0�/��_��啼_`(܃�r-�v� ���zX�ݛ�P�d��m��$#I��E����;�S@�v��v��VX�G�	27&����~,������|�%;���7:���,���n��h��hw{��{���'���\a!���P��0<B"� ���U ЌbȺ|WC�h����@� A!������+x{�D��sԁ$<�Z�`��N:a�&h%R/8Oy��@�$nK�r'��=@
���.:%�F��$	D������a��*A8�)�F����␀�,dB2!@Dyp��� ��۴ض�Am�sSM�$e5��z�@j�L���6����֭�-�g�� �d�u����p%��,�#I��L�.��:ē�e��F'���F�9EN��\���̝�g�n:,9"U�@�ke�Z��k�q��4O[�gj��݆:����������byx0�=2�L9Ի�v۳G4�Ʒ!�Fr��L��6���ِ�g��Ҫ�28�Gg�<ܰ�s�̠��a�#�i˹�3UC�3ӷq!\V��k[��[.{���\
t��(Y�93�A��Nu������6�2�͆�Dٳ' ]
WWCp-9�H��OQ:��cnvsgJm�m��\����y5�V��Wp AM����2n��v�w��M�n��!�2�HA;���bT�%��j	�b¬�7	ӻez�N��� u�`��r�OK�8�;����x���e�z�Þ�Ӎ0�+���p6��#`m��ɒW��n�/#�cnݪ�q�:�1�n�t�r$f�5�B�=�1�����W)�oV���[�9��2�_f�q5ڹye�^V3M�B�ל�&��;�2%	j�ˉ���s�ێ�<�7��+�nۨ�+to4Xr���Mm/.4:9���v�m�mpm�`�m�q	͌u�L�9�-S���%l[��֤�S��f���j��vNhu�ܛ������^��=;8���k����K�N#��:�Z��ک֭
/�6B�
�e^�{K%�i�3H��y�ֳK�3��N0Y�W�5v�	�y�R��&X�RܭL�pS�=����K l��wџ6U�ʪ�*���D�A���C�L�HI�f�j�
�86��kh���$������ �vݺ�t��^��@��ݩ竭��L���r+cgdJ�@��ۇU[b�Fg@+<�Sj�M�<x-\�V�ڶ4���1&F���/Zn�G
6�)g�`3un��ܹ�ww������@�(�v�� 4D�������	�	<��}�ٙ�eɛ�Z�`!���\�͢K�3wM9��X݂-KX�6�D�Сiꢔ�<R�e�g�H�I7��$��݃��Xtܻv����� �*�@�rP�c=vi��ӷi��iAq·Gh��]�ָKFg�w�;6ܗzz��&y�s�yͺ�VGPzvݪk��U%;��m����Ai`rd�PG3�7Uv��w{�w%���
�Ksg5���Mt�;���O]p�q#٭��V{�Nz��N�\Ss`~�ݛ ��vf=>Q�(I/P_����kB�!��	����@;����*D���9�}�5jI?�D�b�M�>4Wj�?Wj��f��W	�Q�L#��Д)�}�`{��l3u�}	$���|�Y[����1��"�?Wj��f��Қ��h����$�G�]��K&l�����]-�n��YT+�~�{��}�׾'2Y��1 {���ۃ%H��"`E��sJXԴH6�Svf=/(����(Jͺ��`g�6l3u�(P��nutȞ,���n|��h��hu�@��M�Ǘ#�ڃr0r+����f�31�aВS�����x��L16�2(9�w[4=��6�ٰ>J""3��K��\��@�wG
�r�/V��>�gZkZ��[s�.!����v��?���5�����%H��"`�[Z$K1����F'�ڴ�ڴ��`fc��!%2t���S�%�6QR䧷�O�g�^I'����
��X�������hڳ\��#M�E76����zX�ݛ�}	Eg���`};�9�,jZ�Ci�7`fc�@��Z��Z�٠_4��q����uSU������<�a�/K��˝��SN:.��h�7}���~�:�ݎd�~�ߟ��L�ؘ�/�>�PM�ၪ�dy����h����@�t���ڷ����y�_1�0���Ƞ� ��v{�|�!%3�]�`{�zt/$�]Q9�`�jI�w�S@����I<�{��;QJ(�f}Ͼ��666>�ײٟ9�wv\�r���� � � � ������ � � � ��{����lllo~�����lll{�y����lll=����������gv���F�M�=���bJv��b:�����v��P%٫��Lt�^Td˶f��A������ � � � ������ � � � ������ � � � ������ � � � �߾�L�we&�f�7o �`�`�`�{��o"?� �C ��A�A���8 ������A�666?�߾�|���*�A��;���nf�l�͛sw��A�A�A�A���8 ���}x ���9�����x ������A�6667���i�
i�	Lܻ�8 ���&A��^>A��������A�6667�}��A�66
� �߼��|�����w���72�ɛ�&n�>A�����߯ �`�`�b��!s�������666?w�N>A����o�^>A���UO"����~�����֗`��=L]Qpu�O)��bP���ҩ�dVlލ9�tb-i�\�aI�5��c]���ۂ���іq������F]�i��c.+��<�ɽNptWn�yz㰝�Ɏ��mڷ.�ᶎ��t�pc4�k�K����ʠE�l�h�bg���R�N@��y�;�XLk�ʭ���.��Ϫ>#=�jŀ�6�sűr�um���I���{��f���<OX#R�7m�ѯ:��╷8���Y�����N����v�:,������w��nA�A�A��~�7��A�A�A�A��ӂ�A�A�A�A���ׂ/�A�A�A�A������ � � � ���l�>�f�l��˗wx ���}8 ���}x ��o~�|������}�|�������g�˷se�7-͜|����~߾�|����﷿^>A�F�����>A������N>A�����;�_�vn�ɗl���� � � � ��{����lllo~�����lll{�y����lll{������lll~��_&k���r�fn�>A������>A������N>A����o�^>A�����߯ �`�`�`������~�,ͦ���=u� n�<�5��͓]���<�Lb�^����<Z�\p��w�������?� �`�`�`�߷� �`�`�`����׈��lllo~�����lllo}�>ݗ4̈́�n]͜|����~߾�|���AuWPQ~߼�|��Ͻ��^��@8�<W"��x��C�h��0�[=ϸ��~��&�q*�f�ddQ��u�h��:�V�~�f���+�"G!�Ԗ��ۃ����ˠ��`$���Ϡ��1���̂nֻ�.���ӎ�E�-휸�^H�I���,�rŃV&ô�V06T��vl��K`nm��'%eR��t�sEK��� ����_B�������,�ݛ��MCl�:��ꦛ���`g��e�(J)$B�r" 4@\Sf{��o$����y!W�,O&"b��ɡ�f+�~4�����@:�4�]`�	� ,q��uv� �m��٠wt��o��?9��C]l[q�]��[���N��1����.�����0=��g�`�e�܈r/��呂[l�;�S@�ڴ/	V;0��#"QI4�f�}Tn��� ��O䒈S'��3;:�d�ChrM�l��-v� �m�m�@�䕂qI�18h|�/�*�����n�P�b�H��^�EIQ�E���.Y���<�&5�Z��4�f���M�j�/���)N;O<Y�5�nz2��6n�c���M+��ĵo<u���r�d�6�C��N�[~ ��v��T��vl�Y(�����L1����;�)�Z�Z���n�J�ήl��j�	T�]2��y0͖�$���p`ͮJ��'19�Z���m�@��MP�)�}�`d�3<�����s.[�$���ۃJ�0�-�NC�_�uKq�s�<v��Z�+)Ů%ۇB��&ܹ��r���iw$�$��gt&t0&�V�*Q�q&Ŕ�;n2�n��=�*Y�Wh� �4��ε�d�e�-��<n��<�SAoWc5ƹ쮼�g��7&܀r]�8㮶dVnxݷ#xâ��h�/q�(���|z6��''�]Ӧ�N3i8���ާy�{��|������dݒ���S�zo�|�K72ip�ow'�M�g�8��x:���U�e#���OX�I(�q�9�`������Z�f�?n��J?�J=@}��;&~bj8����@�ڴ��h����4\����y$Lj!ȴ�� ��v|�(K�I%U���������������yRM �٠wt��k�h�l�*�udxB,��r:n��ǥ��(K��O�ws�m���q�'�jO��4��)�5l�����	%��`!�^��e�C�MX]�yc�7�j��٠��w]� ����Y���r- �m�q _����W�)��8��
"�����|X��7�JDɓ����ԩ*�T��-� ��vf=,�J"�ޮ�ws�=>����N�m�(���݇�(P�wo�z���?n�����K��D�q��#����L�K`$����ki�J��&9�cnk�*27ejp���V[���u�]�v����݈������] �{��6Ilݸ06T��������yRM �l�;�)`f�����wВ��N���N���4M1�7`nk��ͭٱ�����!@8E���I�O=�
�$Ir�&b��)�
H�$"⁌�-*t� <	|T P
C"�VB��%$%HQ�%B% ��VPH�B �B$���R_O߿sÇ �i���0��C�`J1������Wh$ H���7y�J���RՊT�A� Q�B%	m�*J���`0"X0��H�#P�O'�P6)�*@�
���*z�")
F�������C�Az舄@R�/���i�@��A '����T�������{�{����m@X�Q�@��Z��v���9(�Jw6��3k�u)��М�r- �z� �l�;�)�u�ٰ>J"����L�RQ-Ӗ�c2�F�����f{7;��ۚ=��	s�LqCF9,	1����RO�ﾚ{�4�vy}���w���ٙ���N�m�"m5$�;�)�uv� �z� �l�/4�J�mĤI�bp�:�V�~��g%&�s�7w�X9+*��eRuSEK��������w; ��vfm�S�D�7��lv�jd���'U-� ��v}	DB]���������٠r�x�53$�$�񫢥$�iڧ�^u�n����^��YVn�3��I�L18D��;��h]�@?[f�u�hz��6�1��c�93@�[�$�P�(UA�}����j�;˝$k&7$�c�h�l��]�(I)���V�wM���3;�j��N�\˖݇�DB�3�����V��Z��4/$��9$bi�&���j��"3�t� �w; ��v�q@"�A�#�f����׶����%*�KV�ـ�]
ͷS���c`ۄ�W��X�8�Ր8�gѢ2՝\٭�[*�5۸� e�z�tv{vk��Fv1����t�4���q����.|mu���c���ź�v\��G:��O;�fz��32l�jjnr���a<dY��2�њ�Ϸ�y�j�N�+�U��s��w;��+���=h��o���b�h���wq�{Hƛ�ܓ��cn2���8�rz�hcn&��%�N5�v��;8ҰP;N+��o�����?n�������7w�X<����	�m1��"��٠����4Wj�?^�ڟ�pXF��ڍ�f�33mY�!(IL�Wt����;���!7i����J��w��{ɀvIlvK`��_P5I���tڰ=��6�(������~�h�w4˪��!�3�)?�,�$,�&]���w)�	����n$Zg��K�,H�LMA��@�ֽ �h�S��|��h�I}�S1�2,NG�$���y�	�QP?�l�{�NI?|��h{��<��V��I�M��͸02T�����yl�0	=�`o�i�736��rm�sg$�?�L����0?J���7d�͸0"��U�9��bQE�U�@;���Jh�ՠ{���1"6��Y1��n�5e�����V
��&��YT:���w����'���7$��-��~��=^�����vOmu'HT�0&�꛰?f=/�$�L���6��v����IL��k����52Sn��uwM�~��e�K�P��fo�`f���=��IɉǍ8��Z��� �h��4Wj�<�%]�c�1�D������>�l~:����;�-��������M���:�:��G/7rpN�˰%�I�0s���Dm�ŷ;�5���K��pҫ����/�%H�se��-�kK*,Q)dLN��o�?�u�h�}4��M����r�b�U�`͖�7d�sn�6lۻ5�(u3C�m��!(_*��vo?��[�a	B�!$��BR�(J��v����N�C�0&�ꝰ;�p`d� �l��%�&�_���]���X�\އ\L2&^�����[r�]E�F�G&�*frݕ�i���V�"`͖�7d�sn1k��d��`�#�h�u��l�?{�4Wj�9xJ�Y0cdI��fn���mY�
>�߫��3{�`yy$�#b�!��N94�빠z�V�~�Y���֖TX6�R%E��*D��ϖl��Oz��{ÒMPO�@%R�,D�B��r [���Sc(��T�U7MU���P�Gl�=�.B�D���^b��l�ۈ��V{rܰ����&�۹J�ŝy۞��6�X�r�B��Z�չ��\ݣ���Ɔ���9q��m��[b-�����ԗ@�9K�7�l���*i;���n����:K&@�3ls��k�Q��;�)�[R�rZv���Fגr`h�����ܭ�ｋ塀��v�9�p8�le�4��%eۂ�7'_�~�qv����#�鎗���N0Fh��}���3u���k��uwM���O�8,#KjI4�٠~�]��ڴ����μ�E���rh͏��"`͖�7d�ٵ�l&<���RL�=]�@?{���f���)���Iɉŏ�9�w6[ ݒ�͸02T��f������1�g��ٖ����תF��͝��yF.v���pɳ.�)�����vK`w6���R&��lX�R�]ܳ2�˛���y����O��2w_�- �_��w[4ZYQ`ڂ��-P��J�0��`�[���@��o�6�J!ȴ��� ݒ�͏��"`vI�U�Ջ��\��wv�7d�sc�%lL���'ʂ{�������3w.L��7a5�c�+�N�����h/0�Ț1p�����Ό�8F������z��@?{������ ~��bx�cɉE$��ܬ�6��-��ۃ �[P�9|�Ji˪s`���=��!(SBP��H���	v��{9$��o r������q�'$�޶h��K�Y�a�%
gټ�NL���)i���@���=_U���hz٠_uؓ�(�1d���.m���=M��\���t,�z�j˛�n�9���:Ⱘ)�LN����� �[4��M����r�M4�cqh�����ۃ%lL�>j���aX�Qɠ�f��t����� ��f�U���E�$rh�^�~�{��$��{����T�VAB0r�)��﷒I���ےᆏ&�I������޶h�Jh��)��''��Ja���ݛ���md�q��3��є[F8��x�mI�	�7�~��@��z��4_U�ya���s�8ȓ�M�����-}V�~�f��y$�$�Q��x܏@�t��k���3=~�h/��@�����5 ډ�&hV��;�[)����sj��A�����Z���W��=�rI�罼�~*~O����CODHF!jBp�� hKKR$�\
�	%��0�*1b1 JB���Ќbf�����j���?(��a/�!��0���� ��E)B$��0� ��i
x��J~
��;^)���!�X���$�C`<X��>� �O<�"��H�H1	��Ξ��ɹ�t�� `H-���Z����vZyU2t�R��ɏ�{�6s۴M�ڦ�s�q<��Q��8�]]��F�qט+����gVZ�v�E��o�{����u[;u��=�%;1ǰnUhq��� s�-ʵ�e	�m��vɐxq	
K�A�mm�ɑ�)nK�����pAq�9s	3N֦�v�nω;��'��l��.Zڶ�W���Ga��ʹ^��n1�&�UY3��D7fҤj��=E��d�7�b"*{�rN��6}+��F>�]��db��v�l@�%�M�;�U+/������i��Ge7C�d�Y�xK�˫I��u�)�e���8K��ۧ�p��OQ�΄@ݳy�r�D��y/V��m�9z/=nխ9��g�8l� ��՞w8���"�k�S��2���� k�af�E��9��e9��=>8�Wn�6���4�å	��{`��T�tV�ns��g^���	����m���/v�{^��Vw�l�u��Vn���B�)N�P��M�9�jٚ�YP�Y	���Z�����%UJf��l�`ە(7V�=�2Չ���9��sZ�]��n�.|tkՎ.��=�l	��Y���(S�L�j�j+b�(�a=Et�fhҹ�D��*�0�Ny��u%2�r��筴]�����Xĺ���������H c��]��.���,�	' ���.µH�zu
Z�i3���:m�l�[EY�U+�>��;FʛV ����aLۻ\�q��N�T��;k+�i�h3�ʝ��L�ee��d���Neё�A�� $�:Z�(�h ��8��Lk[��!m�z���v�(�i����<\� $ݷk�Ybq���.z���x��h�Z�v�\+�<���}/��,ն!s�*�/R����g�zIlY�$p��K�u7Pu���:zn� �'h��^�6�svx���@�D�����p@j�~OAU�'��Q�Q?8"'� �G�琗�{��`L�)]s����::�m�c��;;��mZ�,�;eP稗�:B��3`8�9!���{i��C��e�=�c��k��qXd��y�G4���m�l٨�v㸵�<+���m�m&�xG�3'c7��œukr��d�m�y�x�s��ta�W%��{�|���m�j�贷f�́��&M���X�<��j��p�������6�M�e�q�)�mi1Y��ϧ�J��NG��e/7t���{���ap�WJ���j���036>0$���~��@��^G�"ȁ51I��u�`n�l��n�gsj���$��~���4�5I�SM�6����l��]�DBS==�Vf�� �NR��SSC�&�]U�ܒ�M�������9Ͼ^��-��H��#N2$�@��z�����{�<�rK`f��.�-qx���=i}a�e����v�V8��ۚ��A:�&�� 
�tĈ/-?m�����JؘrK`E6S�ZT
X�pݗnܗt䓽�{y�?�ڠ�DG���������=��W�2j�+y�27�LL#�@=�}4
�Z`fl|`I[�O����\.�*��7a�%	D�v�X���7k6l����]y�"9����Jh��@?z٠Uz���sۍI<�N��Ԯ�K��u!�:[����j��"�h<r7#ǓLX���h��@?{u�;�]
""?Hfk��;'k��T��МQ������H�}~zu����9���@���8��*��I?~�{9=шU�+���� z���1Ԃ�o��@;��h��J�I���Ho7V�|�J"�{�Ł���M�~��`Uz���<V	ǒ%��4_l�BJ!O�y������c�����EՊ�� f�p�����K����f��;]pa�v�{��؎���u=#����M�����-}V������G�f'�M�����#�ύ��h�[4
�u�x8�(�T�MՁ�c��ݬٳ�
���vOoU�{r��TRj�R����X}	(��6��v��Յ��ĢaD(��)��s��d���91��~��@�(����f�,�͛�	�'Dp�P��U�.n�z{Yrgƻ���k<��8A��&�5�ց��m�~?)�����0��`ubIH]�.�����U7V�c����d��f�4
�W���H���q�$�LNz�� �l�~��K����͗ၫ�r�Y�<�cxF7�~��@��z�Қ���?[��#��3�]]�"�)���n��{�<�rK`RP�/��Ϊ�6ꩡ�m�M��t$p�[f�[	)�K�L���W]!��6֫ ];Փ[��J�%��X�^�m�#��th���:^�>��w�^-��`�ݑ�4����t�cl��nG���3���ӛr��R8��9����{m��nmv���q����r�"��Imf�\tn�'�V]4��n���6�����1�1��O5������S���va����)-�%Iݝn��0HU��fÛ�����u����]�ݮ��_�%lL�%�"�)�e�cLy1br&�Z����f$ﾚ����=��
{�k&&G�ɍ�����W��=��-}V���:ȤQ9��M����=,�͛脔G�"�7��3?|928�m�r=��M��h�[4
�W�r��9��b&H�ǈ1/<6ݱ�Vy �wm�ٮ��� �ܞ�Ob�����0R(&D��Z�� ��f�U��{�4\��5�y#�1���滤�!B��	+��v�,W�h���fI�5�ģ�@;ֻ�ǥ�DL�V�����;���"�ʖ�hr�7a�Js6��3�zl���޶h�u���Ǔ'"nJؘrK`�[3n�RZn4���ڮ�P�eԗe�&Z�l�Cӹ����xٴ�\�Ks��ٓ�<5���rK`�[3n�>��O&F��"�1D�"N94�l�=��=_U��l�?/$���#��i6�m��=,mf͓
Q䄈K(�>\(�̽�`������z�m�̍�M2â"s����y�{u��ҚUg,j�H�F7�cqhse��-��ۃ%lL¤�Ux{Hk���z �8��v;^cx24ZѶ��'f����]��{����˺�t!���M����ۃ%lL���IU�x8�)�2)��t����� ��@;�� ����o&<��9p`d���w6[=�s�$M����/� ��tq������ۋ@?{����`~�=,<�$�~P�B_���ٰ6MGY��n"$ܓ@;����S@��l��f��P���]8�B����A�z�8��]�`ջ!G8^��Ԝ�j<��v�!$]�̻i�t��j��7�3y�X�����4�l�:�X)pRHD�i�@�}V�~�f�w��{��:zt�U��&榕:*���z����|�I~�L�8ʣ� ��MFܓ@;���Қ����4
�j���X�&�)�{����w]�g�]��bP�~������~|�Ê�*ӊj��Űݼ���[.�x�4q�4�4����Pj�1�]�=.k&� ��v�Xv�>����/[rt*W�����r\�ݲ���[�8��s������O}�b�6�6��T��'�H��ؗ��L��7U�q�+�NۀR��<���-�=����;R���1���;�:�v�7p�8lk���R'J����;������~�>�g�Ɗu��<vI8�mӛ���p[;:.��4E��U����Y^��KoͶ~���%��-����mB��5T��M��e�~��С)���v�|h�)���䏗$��)�D���M�����M�0�-�������N��U3U4����
wv��3��`�u�t%
gs���
T�	�Ls#b��X�zX)�w?��}4��wu�Ǒc�"�8��$�m��Ӥ�b�iYv�/V��~��������,n3#��m(����� =��h����8�?{���8,��m�4rKw��q}�wv���.����/�k�<K��8ܚ���Jh��4�l���M4ɏ&,NEUcn�we�	�[������Y1�PNF' �����_ws�n�,�zX�6�K�$�N�0�t\\f^�>���e���H���M�t�I]64�9)$R�"M�4�٠{�S@�Қ������I296�iʻ`f���7n�%�	�[�9�G`.R�%��):��X������'�"�$C�5*EN�! #$�؄HD� �b� bFă<	@�Hl
i� �ljA��"F�b�b&��HJ0�(�$J�HF�K�HĄ�G��$�D�)��v]R �F��"ŉB2�����?)!^?�Vf)B�$	~^<���
�B����7�X��:������D�hJ��)�B!�O��xzR,����1qX�XE����#"� Cc�$N���QJR	���ɠx�pD�,H�W�̓�</�&"��x�����P`(zB��N����DD(��(�/;�������T�Щ���L�SL����n���`~�zXrQ۷Ł��Ss*�d�iUK���L���Ϲ�?�_�ݒ�����(�C�+�6����n���lrsd�h��^�2Hq�u�ZZ�T��`���T݁�ǥ���K ����_���`_��4�&<��9p�/t��~��`��`{1�}	DG��6{�m�1�PNF' ������Қ��;��"s1�D�rh�u��zX�n͆��D!!$D �ċ�D
,051*�h���ʸJ�"y���!FSD��~�&�˒K�&G#�6ӎM�Қ�������v�n������R�։5s��2[�6�������`�;�v��A͡;ev�N�I)�%��ܟ�5o�L�%��-���Qh��c"�$�n= ����$�}4�|hW���G���Z�9 �OQ:��7޶n���`�-��R<K��8ܚ��4+����v(Q3��������������UX��6S ��lrK`fm��8���*D+�A!(D(U���cPL��eM*t��E�h�*a���f��P�������x��j���		�;]��G�u�5XwLWN��[q�RR�u���\��l�㋟�6�qǾ�ͮz�6�oG�4[���!�^nBxt��	jj�n�70�->��cr0����A�y�l͵ہ�.��� ]��Z���:��Nn�[q�+�Hm���l#Y��kQ���w�_����^n�������K�fB��ƲAv�kp���t���:����łJ�X��?��~��%�36���6S2����(T�.�������2fk�������[4��%i$��x��qݰ36���6S �IlrK`L���D�'�	�@�^�~��@7$����������QIU*E�*�`�-�nIl͸01d��~~�~~}x)
m\�L�']nɡ�HN��z�|t"��˳ڷ��\ӵ��9����UW} ������,��rK`Uլ��X�q���=������(�IB��D/�s��V�����v�z���2b��m�@���@?z٠��@��S@<z�YX����%WL�%��-���eH��ĺȜ���H�nM �����ٷ��3+�l��v�D-��!�Rj�y��A���baM��k�g����b6N���}�Dk ��� V���2�5��?�����̩ ̒�rK`n'�Ut���E�U�ʑ0�-�fIl�)�v*�X�cM��ӑh�l�$����H*0���%BO߻�4��h�\Z�9 �'�(�rhd��̗,��d���%.K�:�KE�]7`{���:IFVwW�ﾚ�[4w]s�B�g�s��+�Є�י�p:S`[7q�Sur�s��x-��Z8��2b��m�@���@=�f�{��޲��ܞ;,PPNLJ]0͖�̗r\�e03+�u�9�1�����޲��e4/uz����䒴�dr<CnE,`w%���6Sl���|������-�
��X�X��M:��UI�01f�`{�}����3}~�p`o�~w��mV�.y1٧����%P\�@���SrݧN�Ӌ��<I��X��DS]U]�l�d�0;���̩��R�$$��z�e4z�h�h^��z��<#F)��X��,z�f΅99�Vg>4˺��4DL��Ip�=��h�J`w%����n��`l�+ָ��\�W\�`b͔�̗r\��o$��*9�;.fw0���,w�$���X��n,܋�	�:L놛�m�+�mm�٠n�c�[����NV���� �.hs��v{)����1��Qg�6n�'\�2�o��ό<�gQv䮕�6���Q�q��������j��`�����3�.մ.�l�+�IӒ]�=yVS[��fb,�˵h�@�܃ǟ73�{%l��NN�ƚ�w��󻿝�u��}��o�V�.���N׳\Cacm ˓g���Y��5������78�x��Ϋ-]
�遳|���K���/���u.�=ʤ��L�G�m�9��[���&,������U$1��N��� ���>����_�4�|h��*��3i�F���vIl͏�ݸ0;+b`vlF��X�ƔM94�]��Қ�Қ���������<�6�[�ƛaӳ��wNq���qt�2f3k�����J9�{�4ץ4��Q	~��޵`z{��ҥ,jT����I<����U �|`� 4��a�vh���;�S@?�7bŉ�"q��4��hwJh�Jh�ĺȜ��8�m5$�;�w4��?^���٠~\�V�L�G�m�9�wJh�Jh�l�;�w4/.�I��L�G�o�O�+.8.��Ꝺz*�3�n��Nw��g{]�b�L�q$�4ץ4��4�]��Қ�rʰu�ƚm���[`nl|`nm��ٷf�1QWjT�U2榛�3ٶ��=,بJ�(Q�	(q$�zX��v��
����M�*����͸0;6��;6[}��w7�+����)`�R��U2���)���@�u��;�S@�Ү�1+պ�N��9��l��u�<M��m��vvӍ��S�-����8q�c�����l͏�͸0;6��Ղ[.�4Dӗ5SR۰3ٶ��(J&M�|X�ύ �m���%i$��x��#j��ǥ��q�gDD���v���}!�6�F��s$�,:"����'��y$�����5Dx ,"�������\^Y�cI4�N�%�76>076���ۃ�RR��;�]v�Q��n��]D�z7$�&��ˎ���zk�Mqv�Lk/6���B5��sc�sn͸{�}�zz�^�
��˙R¥��V{�Д���ŀ{����͵|�L���TR�5*]�*�����L���v��?p��&,#�����Қ�Jh�Jh��]dNa�q�!-�=�K�(������0����'�
*+��
*+�ʨ�������TW��Q_�EE�EE�P_���(!  c D�EA#P	 D�U@"���� QQ_��QQ_�EE~EEh
*+⨊���
*+�@(��� ��������
*+��Q_ʈ����(+$�k'�m� g��0
 ?��d��-�  >�   		     �    ( A@���P � E@P�� )B�(  � "�(*%$�D�
 R��� P�
*����  �   
 �� �Ëz���ﳧ�n�{r�^O��'��}i���\� ���o{ϡ��8� ����^��0� ��}]r9�+j� v๷�����ڜCy��cx  }�	   (�r ��S��}g��ڥ�A�[�8 ���{^m+�8�-+�w��v�� �AfҖ��� Y{ے�l>���}��Vg��=���|�W[��j�>�9׶���ͺU�w����=Ϋ� ��  �  �1�=�W�[�9n�n��[������@�Jn�=[sj�Ӿܾ��ݵW ���6�ι�ݼ Z�}�^�SͩT� ��Yj�A�U��9�==)�Y�{i�� ��
{�zV�!�Cs5�B�� /x 
   (@ v��*�]4�]73]4��ΕTp �znn�     @  @ �  � 4   /w:)V 5J�s��@q=P �#�Wn�� ����}|v�s�qgZ��;�}��{�s�J���u}�����n��{��   U �` ^�[n;��q�on��wե�;�� {���l�ݫ\�ϡ�2���B� f�ۙ݇3^  ^�Yy��=�-���/��\��Y<��=�\]\�r�o�H��h��9wi�w���x��*oi*R�@ ���������  �'�UJ�'��@ё���R��E   ��J�iRT� 4)	6��4� h�OQ?��������;Y���.@��������;=�?��bj��DTWj (*�
*+�dTW�QQXO�� ����FT�C��@����E&2�Î��4�2@A,��`���,
�0Ōk�0�,޵�,�0#���c6�1�dh$���r��f?łR��bF>�I(��/����� � ��6(�IH?1ѳ�ް���0��ѣ{�r0Č��pޱ�ű�c�tk|��,׏3If�m��F,1����ı-�g8��f�;w�$���ѧ1�N�o��g�o���3Zپ%B`:R�3\4aY�x��La�0ѳ��f�l��TsG�8:w��h��\�N�q�Y�7�',�ލ���5�><I�[8�o�9�Ɏ���"�;A�p<�oμd�^�8oo��x�D����$:oVw�,�U	��5�-�,�k\O��1�����x�FSfK���fq�o����#5��4b�P����ɉ�Ԧ2��C���N�6s��A��ѳaÄ!���ǔD0��(N��/�Xo��a��C�� 4���$�xZx�H-���� �B�q`e���y���6:=�A������Xe�$�s\<*Ѿ#6���n!`bhXq`�:BC Ь��I��n�	�N&�$�L!F��!���8I8�0��!���4��N,fka���s�81���|H�[n\t[��ͅ��5��O�y�Pf������o�ji{���x�A�g?9��9�|K���1c4����s���$�B�߽�4`h݆�-������OZL;88�v�Vt	R!�'+@�����M�C�iBA�h�9�iE�'����C�A���xsg�a�i��'���g A����É8��7�͡�N&��ORr�1Ӿ�Ï��F�s�s����5��������c�o9���-��~I�%`�ma���?1ӳ��F:��ēA����l�]l�A�6����`���ѱⳚ6���[��8N�Č4�e�9y��8~�,�p��m����s;�E���Uߖqo9����~FO�'*�_��M�c��E08:�a�L,u8FL�$�z�kop4m��k|��LFM,h!�P�4i��Xj�Xa��Mh���L������}���Ĳ ����~���Y���߿e>����������FRX~� 5)�$N	������8�3S5a��),��`��`��C�D���Vc5�8��3LX�e�ae��T�}M),'㿺�����%�K4����?�Ф���I�&�J�,�i�4$aHa��6Bפ�|�
F�v�Fkn��	a�ӭ���ڍ��$`Bɧl涄���٫<�X �# �ˆ��$�����jPӘF��,��b>YoM�с�Y,A�c� 0�hqBX!!#�,�8�YZᰌM�j�@�5��s[4I,�
̱.�$���{�i<�"@�v�f�?1/��+Ph'v���h��mx�>C�i	���VlL'��h7�(q��"8��i�¢�l6:H1�A���8��CD��`-��i�(XY������a�Ԍ4'5�5�<6`xse�,�)�h)��ń�B �g�L%Y&.���Dijf0������(l�7�sN����2��<I� �p�f�1$�(�۽�B0�jLގ2ٳ٠ؒ�&4�kD�p9�؜,��xnNN6)��6�#�2N�`ʐ`�Nb��N�62��6�C$Q��P``$�RS��a``M�����c_������$�KC$�L�T@�̀XA�1�qH�Ò������kAdo�6:Ф�O�pq@��ȑy�C�<�a�0�&��C:'��9Y��%��e����V�	���\��' �&�<Շ�4��9N��ȕ��F$bo�6S�hw�� �h�F������d37��!�hq��zc�|0��0Ń0Ӱ�Ś��Rj0� �0�o�p��A���h#�d�
�0���0,#��l#��a�b2f$�~��@~�!I���Rf���N&�y�,�k��rZ6Q��ܻ���@P[�� ͐l}؟�^0��M��5�sy�o{��P�֧�h,����4�X�Xj0�-!�3~�<=��Lȣ�~M�c�a�٠��'�q0�g,��sC��ׯ<�q�9����p�F84ld��f��I�q�Ӑe���+[8ߕ.k���=5�G���0l��%&I	���\004(�t�d$"\�)LC$HRH$�L@�3Š�q04l�n1*5���`k��1%��q����4o��Jh��m����-��.�L).��fb	`�4�BXR��|�s<�| �\]��H�ґ��������MQͥ�]᭬da�#				��1ѳ�&��p�KX:1I2+0�!�3,"����nh�Nl�Ef���s�6f1��o��q����ZsXo��04�`k��S��5��.уk�g%�@�N�:�a���� ����M�r#L�A��9��ϗ�A|��}�����\���G�����i۴,�0�اn�1#8x���t�,4l�S<	 tq<�T�-	0�u
����9&;#��HC;��l ��F�s�do<:�bi�'�"X�Isz��Q���,��X�$��yj������5�TƠ�8ki�-:�T��J�DF�L�#!���#��I��;�Ǐ�,7���6�NFi���ai#L8lA�}3��.:�t�l6��<"�&ތ`��bp�5�\.��"�N�a7{#F�1|`6txc4m���� �@�(�K��4��Id�J*��Ey�2�ъ�'0\H8�Y�(�0J�;4�;�0a���mM�#�8KG��ڼ-��b��Y�e�H�'F�q�v'�N:?x����g3w4�h���q,��E���lИ.3���)UHNZ�HI�V�Br�&#o��o�8�э���F��b�%0���8k`�$8�8ˊ@��;0t�+��1� A!8��8����a���XkoH�!��[80��,<I�I`U8`�`���v���c��| �=$�`m5��5�\��cf� �\?!8��<n[Sl��1�q�X[�*Hp7,���B��A��N��pf��C�H�(+ۧ���   �  �p�� ���     ��  H         :E���N^�6� ��eZ
v�t�qT��Wel6�wFԦ���l �`ݶ6ٲ�:K�ڶ���  ( n�I�e��:�@�U�*�eZ    m�kKX��o��-� �B� 6�[@  �@	l 	�I� �i  �m�6�H[@� �bE���[oZ�z���ā�G�@uR�����J�m�`6�@ +~���2��j�4�uUĪ��Ҁ���:�v�:�6Kcc�u���Y�3A�`[dE��vm��:�l� H�۰sme�7!z�%
R]�*yUZ���e�k���8m�HIm �� m� ���MZ�$�m	 H��Kh m&��rY@l�km�ڒ�^�8��a � m�4]���R�[/k�� %;6v��ko`  [Ce��^�C��`  m��Չ 9m����� ��6����"�  ˚ Y	v��W��r��tu���Y[TD�kU��}۶�p  �����}� pZ���  �\�	:E��$Ŵ�  ��dN�m��   � V�؀ �  ���q&�v�6Z6ٶ��Z     ��` �  ^��� �m�6��`h�.�Ú&I���Z�̜uv��z�N�[@  �e�\�հ   Ԝ�8 j� �����ݨ࢐D�L�T�j�Y痕jU���V�%[���m���(Y�� ���I�X�{	�]��.�����8��Jq�GmUX�]�����e~X���UW���8�v6�����/;5z����B��]h� �@H� �$�� HH �9�V�wK*ީ6�%v�H�h�`m���� �v�m�A ��� p�    *ݸ�	k`!�8�Jk)���m�6�8�$ �l�$�$H   m��  8  [K�`U��WUV���+�2�0	o  $  ���  ��U���P*��f���ܦ�.�[i��m��q�� 8�s����nSk8�3l�t�-��u��[4d��Bir`�q,�1 $[�:��bA%(��n���6�׭I�I����zn�����-�� ���I� p��[rAmm/Cimz�8��+��U���U]��v'`^z�T�<�m�Z��u� qSi0 H��&��d�i  6ڤYjN`��҃�ݬ3��m�� ���UV
@�nj���9�  �	��@ &ص"� �f���U�.����U�  �`�U����J��Wԑ�+J��5UT�t�����J� �&�mhm��.��J�B�l����-�q�f�i��	 H',t���'Yv�l�ۄ��i$ 6���p9���&^��  ��8  lm [H1 ���΋���[,3m��`6ɺ��m�*@ @ ���m�����0�ة"j���j�q��6��m�6� -�}��:����Ac,�M�bY��  �m���m z�,ML��ܴI��ƷZ$ r@ ��m���6t-�\�j�f�yl�õ/l�e<��m�[��� 6���\Ia�%�h�l��m�n]�� 	օ(��` ��m�`Z�����
,��J��^��lu�Mk�-��b@mY��շIJE�H�^��H-�`m�	��9r]�6� tZ �mF�n��m�tq791MUR�mPR�;ih�5���Β^-��$6��G>���jI�����N)j�҉UUm   mm��5� �;l�m���6� ��m������i6��յJA&$e�  ^��`�$5V���8���m�$��m!�m�6��`  l� mm:[I l���y�I�H
R�h �   �`pm�6�� �mp 8�[A��3m��I���Jᆽm6l�zԁ�ֶ�u�� �F�  ��� �  H�|���pz�  �ۇ�h�� �Ĳ���K�n��m�T}o�}t�� �-�l  .�l��@  [@��V�րl& 8���ml����i3�l�6�m�nZ��Ǿ�km��4`n� �` l l�Cm��[@�o�u*A�ѻm��c�sB�N��� �`q,�9d[E��m�` �����t�h�`	 ���@s��vÛl6�۶��� mm�2M�mJK���mR�Ի-U;+Z��ࢥ[Ҫ�J�ݶ����n��Z�C�����N�a&�o����n�Zڶ�U6UyZ���ZL-�E�n�t��.�8 �`H�
l�e��l�a+. �R7E�i1�NT�鄅�m�h��m��NU�ش�I�   � m���yZ�6^/+@M���%�aɵ#���-���	�-�4ۭ��Mr�G  $��6&��̀�N���K���� ���d��8
��UZ��۬vL+��*@�%���� m���f�4�x�7UX�1�[*1K�J�r���q�UTpnҭ��5R� շV���V�h��`6�Y�`s�-;kw'u�Np5\�@U�@B�ۧ�� ���.�-�vh��0��T���A�a�����+�s/a�r�rk�{+^[��Q��Vۥ�mI�&�x��f�6$ �WL�m�3❶��X*�˴��2�H0m6Ҭ�U^iV v�I9&nNIR=�mrCn�N��m�m� 6��m�m�� �m�U*�Ҡ5U �V�86���  ﾅ���ͥ��:��l �5����h/S`IG�8�U�bϗ�[��7R�]a���U)8�p� �`��Hp9�ж�� 8&����8   �m����-�n��F$m�i�[`����igjl�w[� �&�_+m�i4�sm� É  Ӌi!�-�H	�n�ɶ� �ۇ$H� 9d�$����{�$  �Z�]��P�7UT�O	&��X�I��O)mxm�kHqM��Ѷ��$�MW��z��J l	[%[v�ڻ`Kh���K.� �`	8H7m�-��l �j&��-�� -���%�m
��l����5�$��-��.�q����@�em��v�-������;kV�l�a'h	8�& $  �m+6 6����
� h[VյΝ-���I(u��Z��M���UT8٪���c�@�E��I��k��IÀ9�5���G/]nN��C
�*��U��Z:ɪfm�m�� �� $m�Ȑ�` [@�I� ���u�]���m y(�b@h �m]6��  m��ŲƲu�kWXu��[BD�l$�m���ӶH  �i�M��ci+`!� ��\�� ��Am���[���V@�j����� ��ͭ�@���s�  �T��m�	&�۪�'����  �s�g����ߋh [v�6�p �J�V�6�e��� H� C� �`��� CF٫a#�mj�  m      phm&���5&�  ���	 ���3H�ōsi�eNeP+` 2KD�� �`   �v�m׬����\$       $l[~�}'O�7 ���l��{ ��m�ӧ��Hp  )y�ޓi6���z�[% 8 l-��Zж�5���i*�I�@t��sUUUt-���$ 8[]��l6Ì-�NP�I�muh�h�Lݤ�t�iv�V���K(8Iaz�Mμ�nĵK�D;NL��dÒi���HNNd�r��Wh���y!�,���2�6݊�J�����\D�t�Y��$m��
'j  I!�m�m��&@i�j�`[Z�/e�z���ۮ���[[vn�@  k ��E��πl� �l	nڪᶪ��YZ�v��| 4jΠp *��ivZ�Z��ʨ ����m -�H�M���'I6    6�AؒJj� �$  ��i$��m�H�8���	�j���J˲��v�$�n� m���n@5���KK0��G.l�G���ګj�-�ٶ�ͫkhm�'�o���u�&�b�v��e^�T�mT�,ZԬ��eY ^Km��� �^n�m�)�guK�ٶX'�=��w{��SO������:Q��؀�����O��@QGo���(z�� ��G�Eػ@�Ae�鰈E|6��A꿑T1 �l������~6�+�~<�w���z���j�p@i`���Pet��PB*�
���!�}舞 ����h �"��uC�G��W�"��lA�hQ_|�}E} �*&�OIH%Ba`�VH&I%e�A�XT� `�!�FiB%��&d!ڂ��A��1U��8�#��҈mȧ��!8��< &!D���O������P��zu@����PW��� �Q����B��$� !��:t=�`~@Q�U_O vz������@�?/�QG��dAj:������a@�j���(����#A@��}���f�����*�k���*[P�5����ؓs�8vɇdv��WU#�p��r�(▱��������g���9�S[�8�M�p�.$�s�Gݨꭓj�Wn��
�:���v�iJ6
��J��퀞�[\��v'���.v�m�:R���i&FEn�A�Q�}I��b��*��0��FmWE��g�t@�m/nv��X����D��کV�#���6�@�,
�muAˁu��mU
��ԷԄ�u��[vΉyَ�b�Rƶ���=��Pۇt��u����6�QB����v@���s�$���q�r�5��N8�kpS��n��P���땨.��)�2�K�ew>fU�jn9�th^�7.�RSu��j����N��b���"t󽡐��Sl���	�ۍiA�]sp-�*�,y\pU�) |�6qȂs�4h�ed�$�V��m0nr�	-��C1�N�3Pm[���]�䖭��;B��{�	�[�ظA��W�m�Ka�Ŷ�l�v������^�gg��t5w@�!t��WMˆ�	��\du3m�uma8�vg�r��Ghۜլ��uY�g�d3�ヴ�'MAz�@���Y��#�ۦᕻm�aj�Mpc�ê�N���CjUΝ��	lܭ�ݧ�)rT�A��2�P;����U�gXh����x��������c���i$�&�E��y��4�i*)ص��=N��}luÐn�m�h��*�zX,,r�ya��vv�[T�.`5�p�ہ��]��՞�N��j�U�#ڶݸ��ZAxw
ۚtZu;d�G2�6Rں���3]��n��l���@F*�xsU]C�1���f$�p[r�؞f&�5sԎ�;{uv�6�\z���Hf�a�p�݌�P.繳as��P� B�u����l4�v��\{[L�����6����p��%�z@����h\�0��]3uN�2�^tQ����x;
@0 C23,, � L$#1�0��)$��� C���v?
����;�.���T��4�:�u�ڲ5��=`�nN��5�\�G\�uXe.ƛl��&�kL)<�6���G�8��r�����`��v��2�<m��Ӻ/	��u�q��]�u�1��`��@M�&�i6v	�O �:��[�;;0\�Ǉ�m��n^s��6]����lⱽ�;�U[�n}�<.�Y�i⫙�9ɦ-�{ݯ{��<N�� q�7
/`|;�; ���t�������DD���r�Oﻸ�۶��۷����@�� ��Z���u��V�v��9�Ϥ���p��� >ޓjr�5#��!�zZ������Q���W	$�f���ܓ ������֪0KSH��r��Z�qa���0=*�׭��j`Z��o�z�;��u��cQ��8 K���]$��]md�-�Tl���vzF�d�`z���=-LKSӭ���HT^Z��˗��r$���K�4@82�k@��5Y��*����׀oӻdU7Xʠ�Q�n n��M�S?uwN 7�x�zmW�T^2:�$� �f��?l�x%��I*`N�p�pov�;W-`}z�`Z����[��M����j[����ip�rϴ�p�Z�T�x�%�㛕�/]p�K�-qZ�ȅ�c�	-LISץ�׭��ڳ�ԅ����ܓ �T���u���u�OZ�$]{�����K�_��{�����X�� �(Q�P&$$$h/U��&�e�i8�//|�w�5�v`��VUc������[�z���-��K�	%�ܴp�Dj��M=������-��K��n����>S���;�Ue��#e�����۵��1&.�\eX�����ui�TT�0�T:�	���^�� �gu�l�x߷n��M��P+9QIl`z�����u�OZ�e��$�j�����»k�>ٺ��n�=�qq7�}�w��x��ͩ�j9n�U\��w�l�u�|���
9DB�SBH �@<9�$��$��I=�k���X�����ܓl���Q���� ����3z��NV�WQ%v�6�AΙ�4E�.�ڝ���[��5ȣʲݎI���*����`:npu����0w�2�ʈ�r��L훯 $�0&�y��Uҏ�h,B�F��4�߀-��L	��`z�F�n�~��"����Fʤ��������u���� ����l*���J:��ـ}�u���]����6��������u�{�<���D܉�PĘ�����9�s6Fj�VZ�q�q��ԑ�,p�[9�O�r��hv*���7d{]�ݲ�u�����7\v��/�V�qp�a���ŧ��!�R���PMs�����)c��@5\����B�n�9;v�;���#vam\�t����=n 4�neQQ��ved�-j��4���Kv���q[p�����ε>�-��#Hy:Ց%i�Nn��������p�9H덣�G6�'W^Y4���^�K�&i�9㶰��+����mn��ލ����������1��gwg�Ͷl�wm��vmV����I+��������H�����Ͷzo���m��6�d٤�U��mNK^6�������͝�q���w_�Ͷ��k��}]�M����P�r�ߛl��+���ۺ�~m���^6���v~��{ݦYYTe�Z�9����U��ۻ�b�^��Β��n�\Wm���-���"��2�Y)L7f�rhC��k�3GK��I-�2��M���[����Gg�\����{����}���ߛl�w����ߛl��j	P��j���rffv�]~�ԭ�d%
�I$�>\���.*6{���o{{���m���x�o�ޛU�
�uE$����;��q������m���g{����{�6��n��»k�7两���?ߛl﯋���;ݟ�6���ٍ��ڻ6�@RF^I+�����v�m���ĸ�w}~��͛�q�������m���5I$�i]x��kp�۵��$De���8X;a�vVή�el�Ƭ���4| ����~���'K�����[�}���*�����Y*��
�m���͝�s�%�#m���Ͷ����m��wo�ͷ��e��FX堣��m�ۺ�~m���^7�u.���@�<�o�o�33/����337���J��T�+��3.?�m��ow�U�ۻ�������[�}��N�rX��#eR[k��o���ߛl��.6���u���o{v�m��w	���U�X�b�xh8)���q�]r]���u���H�#��B7���n��]ٹ���~~��| }+��n�튭{���������K;m�NGY���?vn���I&Ͻ�� ww� ;���$�}�g���A$e��Z����T�=�S���I�Ih2��ԱG)��s����w����ʼ�]�r��4�'���+Ē|�v�|`��6J���J"�$��j`}:�`{�Q�zJ����²����;$�4A���]��m���r�"nL��۞{]��4]�mN��Zۑ��^���ު��T�=�S�q�SQJ�Eu�2f����3���w� ��Ɂ���zU�`j�Vwn�9$��*`�������Um�X�%�/�j�{y&�J�J����Q��~���0-�����vgr��0>�Q���� ��0z[�b\�Ot�����,!bV7.�Ƌt�63���֕tv�����E���ݵ���5ë�v�NX|���R�7HXݣ���Oc�;q��M��e(;7n̈́�z��0O[��!�3���4��+:͹Nk���/��ہ���NOn��=���P�q�ϔkS��97"qً n���ݚ9q�(�h��4�v�|c�m�r���j�a�r�~�w{�{���w���~�v����a��qF�jɒ�x��t���MJ�UV[��,sН&��~��@>�IS ��0>�S ��f�h)h݊X�)�w�pzT��UF�*=�&IZ�Xn-\��mT�� o�� �ݳ%�~�|`��0'���i���5,�I0>�Q�����T�'�L%z�_�:ɕ77>̬��s�0N������?wn�t6�u�D��w�7QxWD�ӄ�m���D�h��]�G[�����{��c��Yݺ,�I�T�'�L�T`}b��!f�4;Vڒa^��w�(=��H:��7ەy�U���dU,�� 3�yi��&�T`}b�7t��0	�S ���b�#��_�y�T`��=*`zUF�^��$�wvjXw!�}���	K���}|`��0�I驞�`T۲�Ya
V��gk�7���s���]����4��׵����;�v��K�?��Ҫ0=b� ��0'���g-��7{�`}�^0=b� �Ҧ=j`_J�r�;9��V�s/�7����x~X����*BRUEi<Q�I34a���|I��`I�5@��@�IH1#A1?a�h4��1�����=ݤ�y�����4�$���{{&XCA3��G�#���Bc��<Q��V6:AA�DC�S�𢚄$��/������ŀ��uV�Vwn�;�C �Ҧ=j`}�^0>��0{�j��2��8��7x���>{l���x�Et������,���zz݋uf��݆���o7	=i��xն�0U~����b�>{l���}��׀��Z\$`wv��c�*0zT�'���۸���f���v���$N�ILD�}��?%�����ŇL����:��e�U�j����e��{�������U���땇�G�>(��������{�u�Q�JT�� �ּ`L���j`���왭X��[�uk�}��ŗc�����ӥi�]`�&ۖM��S}Ygn:ު���ϻ�/��=�S ��0=�^0e�܀�j�w$��Z�����Z�����b�,�~��Xiܓ ��0=�^0>�Q�{֦�T��D�������X��=�S �T�=ruY�0;�V�\�����޵0	-Lz׌����]K�h��s�+����䑖��C�mA���/I����2/h�l�td�ٶۮ:���Es,ݩ��Z\����k"p�v�,��:Y�룵�a�Q���j�͍���bt��ɲ��WD�Z	�J�Uɦ���Q��͈�;&Wg]�V��������ݠ��[���PO7h�ۍ6w.��=�e��72�KҌ�3ٹ�<��[(M�ms72ƴE����ߝ��_��V����]�5d�Ƚp�R&ۋ�"��o\�J��m����R�Jt~�� ����Ҽ`z�F�ֵ˃qjIg��I�Ij`}�^0=j� �Ҧ�Ww����,Y��$�zW��T`zT�'�L�^�Zgg �Է����=�W��>���OJ�zW��yw 5��E��!�}�S ��0>��X����fʷ��,-��!�t��,����<v��Vݑ�k�p���"����S/���ۀ��p�k��*0z���.�����9Xܖ�}��/�\K�H}�0o�LzT�>�:�\$~;�E�\���� >��ÔB�2=}x��X��W䅆nrùz��'�LY^0=b�g�k��\��r�ԓ ��0=ex�����j`~��2���ݚ��i��[#g���vv��9�r;�F�ڵkhm<qFJ�`n�P�݀����`z�F��0	�S������۵�����o� �{��OZ��Q�[o.��Wh�Uݘ�n�~n�p�Bq
"!*Y�J2""���f��f�wGj����ڰ�ԓ ��0$���T`���u\$�����I�%T`}b� ��0	�S����oZ����bA��k�m��u�1`v6��ں.�%�M��xӪKU��	*���?on����'�L	*��u�9b��Xf�y,`��=*`IUY^0.IZ���˹w�����%T`z��zژ�]�Xv%��W���0$��Y^0[S�ظ�o�n�{���
)A�+������� ��0	�SJ���=���hMٺ!�c����٫�m���25��#Q��Mv�C�hv�f[lX��\�w�Z����eT`z����U�� ��Ն��`֦�Q��+�e��d]W	a��ˍ�I0,��X��,�0	�S ���b�b3��Zq���T`Z�����\���<`�{����N9�,�0	�Sʨ����?b�q#�K���s��UN������Ճ.�֍5�Ϋ5����]&��fM56�u��l�ʈ=]�m�n��j-[{nv^��N���nUݝbɧ�OVw.����ܧl�Zrm��:���4u��%�[�K9��q�O�v��vݝ]:{f}�2��3sZP���FDt��Ƅ)�M0������m������N|���';����D��u�LJkW/9L�]O���{������	�^�\�࢑�#ki��EHD^��A���Z't�U���S;�yU]� s}x�l�>{l�$�H�� ���r�+\��Fܖ���X�*0-LzT������4�\����=�W��,�0	�S�^0e�܀]���E��!�Yj`Ҧ��`}b�퐫�@/۝�9$�'�L*������!�%D��J��5T�USX:�ѷ=)ƭ/<��;Y��OGH��K�Bӳ�������I�eT`}b� ���'����ͪª(��1�`��L��L$P�� z�.$��
	(��+�;�����f�j� ą�nr��C ���=�V�J"g�_��� ��˫��WE����I0zT���0>�Ta���}���;ݧ����%��-��n�}��~ ��x��� ߶n�"�ɫ�\��m���s��n3�Ļ]���p�C.�5tg`�-n�QZ�9a��.�������J��Q�[/.��.�(�Wwf n�y�2�� ��� ���0�zmUJ�*dn�ۀzT����?{3��}�Q�Ij`[m�+�NV7e�۷L��t�	-Lޕ0\�ya���v�ۼ�ު�KS ��LZ��.{n?����.�P�v��7]�Z����L��u�X����Ͳ�s��=�ӛ�V�p녷�	-LzT�=mL�T`L��˃s���GrI�OJ�������KSz"� X��Z�����׌�T`Z����=(�PUZ�NXfL����� w�� ;���#�bb�HB�H# @���As��xr��}�z��uSD������� 򗯯��ذ�ۦ�.�]�7q��[jŹں2n�\s)sy���m ���#��Dog��s ,ӷVrI�OJ������ٟ����=�g���T�9Xܖ�z�g)��w� >}x�k� �VӫÖ#7C����0>�Q�K*`Ҧ��`}�q�HXf�{��%�0	�SY^0>�Q�r��mCV����� ��ۀyqs��o�/�~����W����\6��H z�Ic43����`'CW�`�H�T�i]kz3F�C�RŜI!�Ha�l�01���i�bi%X�.:M�)5KpQ��,�,�*0��˚(=�&��� Ě��, q�e%�<]2ca.e��,0cAi���)$����6
A��Te�0X��᠛	�F��������FAPX��Lcea��folE��7�֦{(�I[�a�"04���Ve0�,�D i�l���z��"b4���F��b��j[�h��:`��F��.mv��H�h,َ���6/��^����`p͉������6#��F~M���y�E�K�'������?�_��]���	��Ž�( �f�z0���#��L10M�4(�U��$ K�G,#U�;���Zѭ/ !� `�8�̬< �Ş�p�,4,a�b֣!$Ι�e��p�2����i�iF$�L] �CaX��h�
	�����6g�5�i��BW��H��8���S��p�p��}���m��Ӄ��im�����wo#���8��R��mɲ"��@t(O;=�<�2G��N8�����3qc@�uD�j���c�4uZ:��cc�L��d	ٻc�Gfe�+ݗ8ZZ7\��p&6jǴ�RU�Z����Ύ�E�1)mM-ɷ\����b,��y&�	�_6j��+�wD;R|p��L��a��n���M��#U�J�R��7%6
_(�U�lx�!�����W�@���Ё!4�sh86�9����z23H;U�_\"4s"�>ݖ�s��N݄.��T�b����5����Ƅ�ר����8j��i�n��ݻ���-�kF��@�z�flT����WR�B���.#�yo<��
#�ظ;c���4�i)I����ggJ�����d�k��\�x�c�\��8P���tx6���5��(rֳ�;��eg�JF%��P�U: ��0��T��V�8
�]�98��UX8�S +��raQ�Ց�q�7�E���5���ѷ�qc8Fv���n�2��7& v��\���y�1cS6�l��P=3R�Z-�٭۳S�4uI��r+n�t�[t �ݸ� �å튣�&+�r:�(�y1p6���m<a��&IDge��UÓXYc���һ���Fs@-Ԧ��c�'Oh{7$��*X����'DܐL�N�hu�aK�,(u��n�ʛ��ҽ���Ͷ�N^�Ɍ�.Y"@�by���˷i�Ͷ�n��hO<6�un%���<���/�Hs��������?{}��.�1fb�ɳ�$P��v:^�&��yW�r�J��׍Pl��m5�U	�eR�֞�D�4�[qa�t�۷]H�5�q�g=\�g��q0�(U�*t�����$��RgӑY�����)����Е���P��Vz����R[t��^VڤV٥y�B9�c��ƌY�6����Kf��f��a�ۆ6��C�{�iC��S�P��������T=��j˛�e�ӭ�km������*�����-�d�9��M[ ����� NLpOk�ݼ���}����ig<͎6Έ�z�x1;q���C��7Yu����g�y.�q�V�Oa�Q7'R=	� ���<e:�����㠓+k���K=0d<�'HA�	 I�V����8�@-,ó����bw�Z8�G����Ւ���5'q�R��5�c��*V;;��ӎl�]���<�6�)<\�����b�kEۆ��]DЊ/%�x����YS ��0/�1�
�Si�Ws�;�3�..6�׀{� ׯ 7��n�]+EM"��ݘ�]������W{�� ~�b�>O�j��T��D�ہ������>ŀ}�x�9DL�}xs��T��Rr��m�;��X�;�{����\ ��ۀ�f���"ڥlvᇎ1F��FԬ��x�YZn�[r�RY=�n!c��r�f�p�ur��k�,��{���?0�o�`�zz9P���RZr�����S�*>*#�9^��w�?ww�۸�ˉ6y{��CV��7���`&��`{ּ`ʘ�E�@�-]�����I�,��x�^���P�L��^��ɻj֛����ڛπ���� �T�=�S��ŀwW^�#�����"n��bOi�7[p�b6�D�ק��L�#c�o)3�OH��Z������ ~���5����ý�b�:�t��V�S#u;n ~���5�ŀ}��X�]�B��Jd���TV:�"r��m�7��X�wqa�RP�,�H��������m:�U�+TZ����Т'u���^ ~����������f�*�>8U%� '� �,���.i);g�oS�0
s�`�޳E�!��C��"����׵����]���#a���_�0%��ޕ� �T���.��j��ݽ�ܓ�^0=%x�-�0���=(����ӷV�Sy���YS �Z���K/-H1vj�;�˖0	eL�j`K+�	4�9�	`�����:�t�T�����8� �Z����+�l��<~���c��7.���5l��O]5ۇe놔��շ2�Avr�s�\�3q��Lex���� �T�>����͕�&��M�V�{����I%2�׀>��׋ ���\աRY�����c �T�>����`zJ�r��j�q#��o#�$�>����`zJ�[j`OEwybZ])�*��� m�XB�I�~����^ ~�� _�A
#M8��
��dSq�t��,M���W�^�mK��8���nI�;.�k��n�^�NŎ�N��sȫ��[��e����ɣ�\��ƶ��ݰ�`P7s���m���3ǉ�<����sa���b�b�7Bm�2G*ץ�ñ������=8�.3�^����e�ݖ�nh��=�vN�h���'�`
D:��BW�Bs0�0�RR������>.$�qs��&���Q��U#�R��gqvq<r��N�ݸi�]���5�{�?����W��������� 7wn ~����/�=�{ w��sv
�]L�E���X �w�I)��{� ��ŀ}��Y���}�֩[eヨ������ �x���}� ;�� ׶��+��A�r�W$����J�[j`{v�ڻ6TJ��j6�X�wq`����Lmx��̆��N+)�Z๢a�E��`���1�vm�w �\��7f�E���T)j|p�KV n�� �֦��`{Ҽ`\��ڰ�K��9I-��۷'9�$���� ���, ������M���7(Ejv)a$�&���x���x�-�0�j`OK�ʅ��5W�;����`�v�DBI)�}�`�꺻t������X ��xB���������X�z��B�J��v��!�ݛq��g��ݴ������l�oc�y��j�����VrI�}�S�W�zW��T��-�;���.5rI�}k��+�d��}�S ��ז�*U�n�`k�`z��IF~���f�~����`i4ڥB���
���Q3���_u��Ł��IS�~�y{�˩�J���TՕWw�kw�rJ;�~_���� 7����:���(�a�����G�6Dv�#�nIӵ]l�SO<јg"���i��E��ߟ��� �]� 5�P�_�}׀v��r�EknU���/�w}|g���8�o�^ k�^�Y��СBUA����
�]UR��T՘��� >���IBo}�b�;��0����+M���GWx^Q
S�z���� �]���ʢ�h~l��}�U��}�F���v���W$����U���wn�������bV�+�uKqe��^�
���[<�g#�����N�����������d��Q4�*nʾ}�� ��� �[�IG��ذ⻮��+�SE��� 5�y�D�k��v,�v��I����X�l�:(���w޸��a舅QT��� ;����m�B+S�J��Kp<�����﯌ ���=-L%{�����7���_�����/������5�� Q%�}�Omv7l��aVkFo��'��:.圙R�R�H��OA�=�n�h6�gZ˥���F6is��q�l ν�n�����1���v���}ǚ��5���q�M��]v��<0&ey��9�ݵ�
: �x��� �3Qu�S�Ҿ)�t��E�ݜpA�p�ɜ ��ƵSa:֍m����v2g^���IJW6_��GvGV=��w���?Vڐ��S1�s�wԶϷk#��wN�h1�Hv���;p3-ۧ�^5�o"�{���j`Kk��T`y?�m���x��$r� ��� ���`zUF-����bĵv�����&��`zUF-��zZ��'^Xr�f��7W,`zUF-��zZ����u�;��f��j�0	mL����׌J�����$�C���p��7hݶ�MPmj�a��Y�=��$�nJ�)WaW���Z���or_ K������U�������e��$r[�wwqcOOJ��%�0KS�^�Zvr��;ug��7�/�����j`K�� ;��ʯ,r �G)��ۀ����`zUF�}
�-�զo���I�zZ����Uwv�}�)*-+��YK*�R<�\y������c'֜��Ii�m�ڜ�wjӗ$����U���}�w}�j��Q/(�P��*�>�����j`Kk��֬�Xb�>8T� wwn }�ۅB��J�XH" ��$ �� BQ! z��P�h�C�P�CI�zD6�)�;�L~#��b8)8�H$�C��&��*&	��$e3��2(<4�h�E�r1R/�q x�`Fxb��u�Hl� �/�`�����j��a,\#	&J��P�%$���5��������<�AӰ	 3�=A�pC�	��P�Th�@T3^w��0�n����M�ҊIG%��j`Kk��T`ژEwybY���wv�$��׌J��%�`�ݸ���XW���ժ��F��ǆМs�����u�q����V�db�딲8F����/�w}|`wv��ݬ	mx�%��$-Gw,]��-��Ij`Kk��T`{7Щui����$r� �wn��Ň�\�M�޾0}�\�ν��]�$��^I0%��Ҫ0	mL7?g������]�*�j7eX۷L �j`M���^0
\�pK�s���HQ��)m�`��8\>zey����3v#'P�V�	-RT+*|p��L �ݸ_wy�m��Q�l�n���V%�����e���׌Z��-�0$���ė%����˘���U���o0$��r���ݼv��T�b�Q/����xηXm����eU0�� ��)��� �O���݋ ��fIBi$!	D��I�DBC��RI���!##T��	J#!II����e�T�L�MV_邎� &Xۣ������ݹ��)���s	϶.wr����]�a&�۴��F�{nl�=ݜ�v+�.�P5\�紪��j��id�9ӝ�x]m��ll����sFN0@U���T3u�k�a)ʝ�����kt�@a�J�\gM�ě���!s��f�a�	�uc��m���v��n���p�"r��ox��(e�2'a`�]����,竛���2g�{s�:����`[��Kl�7X�D$� ���`���Z��-�0>�6�X���;N\�s�^0>�Q�[j`M�� ��vʇyF��M�V�v��� �-���`zj�H1r���f�C ����-���`z�F���Q�굩%$��}ݘ��,֪0mL'mŠ,Y�klF�������9�9w!d�.zɉ�\�s���5roN�p�r�V�j*�I,���b�>ݺ`���:��0���J�R�"����p�~�\������'9_}Ϸ�:��Lww w��*���8V8�m��6K�mx���F�}�m��������u7��n���>�$������ۨ3�� �K����U���o0��߷󶺭ڮ`�a�
66���ms��qi�utO"���tpX�kɺ���������Sl�����u��bĖo��f�C ����-���X۷L~��n��uZԒ�Kr�s��\�����+� !�FA!�de� +�����w޸{ۮʜV�hUf��� {��v� 7x
]>��7w���l�A��ˋ��������r�� m�X�<������./<F�TκA��^ͳ��K/#Ӯ;=\��^��E/$v�eU5]����r���p�n��������� Ծ=wVJv	��%�_wf{�6{��,����� ���*���A�UR�0�ŀ|�áDL��׀9}Հ�ݲ��V!B����I���x�}��W��{�R	#$����{�Q�I��!UB��x^����I���6��v� g�MN�	W�.o5Уۛ%���]vyt���b^!�:��*~�Iܱ�N�W��g�5￹�$��Q���y�$WW,�λ��.ɩ���7u��B�	y(������ ���XηY�IL��d��4��iIk�����ޜ�m����������eU0��ƪ�J�?��q%;]�X��X�x�9%	)޾��5>��ev	��$r���� �[ŀ|ݳ �[u�$�	5%�� ��k�g��}6$�l/�8:׆i��n�����l�nڹ��g�1ѽ�륋�ɰ��n#V7i5m�ɹۜ�9q��2d�ֆ��e�lT�*ٷJ���Qm׶:ᨳ�H�rE�nXY���'U��k��|��4m��v9��7Q�v�=�ܦ�0J�H�úр��Y�!��۷T�8�Ս{z����kY��V[�3�������5��in�.���c=[6���k�� ^g3�p��9��S��w���|�t���*�Kg@���ŀ}�t�?=ݘ_wf ~�ٲ�D�B�N�V���?�DDG�$�Q��z���� �׋9BM��{ΫBVP"�S ��ޘv[�	%x�����Z�Y�٫8EM\�U�(R��V ��X��09$��������\N�c-rY�w�x���`��XηX�7�R��(h��9��s�k`�<;6�g:�\�6Ř�S�f��ӿx������wH������d=�W��N�[u�l�u�H6� wwU�T�]a��+�?=ݙ���^`I+��[��7K�i��#sW�ڰ��\��o�0$����������ŋ�V���f���$��n�>�o0&�y�}2��vb�3����0=z�`}��`���q`}]&�K
��H�n�[%t76,����<2m��Ol$uv�u��=��][1�;;�or��m��j`I+��u���YT�N�R9[�� �wnt���Xu�8�m�����\қ�c��7-�;��,���Iq4�9��>~�� o}�o{��ڣ��������p�۬ ��xJ"[~������T�YH�U�S ��v`ӽ��m�,u�0�Z��UTr��&d��WWv�N�ۛ��`���^��������%��W0�ev	��$r����p	%x���0>�o0>�6�	n���囼�&��`IU���=�� ?ul�Tq'Q��*�;ݺ`����&�u��ŀj��j�.����f�!�}mL����W�7�c� ��o��U�z��������YT�RUHIK%�������I{�w�_����w�|�)�����^��לsy�d��b��J]��[�"ڹh
EX��������~�}��x���0���zژJ�$ob�G_�1d���_�I&��{� ;�z�=�$�w�����+,h��� w^ |ۼ?�Je�݋ o������4�����p?���}���]ذ�l��
g{�����е��*nYnޭ�X{�L
��{�U~�{�U��WH&�/=R$BaLPYH��E|U��a�g� �M���:����� �d� `	I@��!��$��"!�e$!!�H  `�	�C��$D��0�a�A�<,T; �����&
Y�^���)0��$\��fI����b� Rq� (��$4;v�&%�G��A�eIl�s	��@����v*qX� ���[D��������mL5h2��;`ԅmc�`R��l�Z�[-lIW�ny�����K�]�m����X�mv�d:�\��h#u����ε����7 X0X7U��s����tl��倔R��x���ٺ���@S�*������m��
H3U&�j�xR��_��LH4���k ��g��۪��ǲq�;=c��2��n�jk��#�]Χ�m�tϴU �#�$ssU\jUv7�:aکv^�7N�HN�{���e�M %�MvPk�ܶ���N���V^�TS��Oq3�[�fY�TJ�EƷgM�V]���
�/Ar��Z�۶͸L�K�nɞkd�ǉ��Y�)a�zM��q��s�5JD�=�n�v͌`@ᢎB���:�ۖ��\n�Í"��)Z.�v�&L�`�$�j�s��  1d2f@���n�%��`���]����\哂��5�;lsh�eޤ��e��E�ת4�[�T�nH�U��Y.�U��zK!�[����l�tt�]Ts�n#=�tr�xr6.�v�����Z��n���]�P��x�dx�dܲ�Ֆ�#�Z궥,��]�����@c�tZ��1n���Ñ�W�����*ݞP�:謽DgWn�Yյu�öw���(�����qS���u�d���qØ^�,F�p�Z%���&�	v�<枺��:y�)�������WmV�JVܙ#<���m�m�i�h�=99�I'8��ۭ1�^-p[u�H�\m0sY�+�ݶËkql���[m�"�Fs۲�Ƹ[��8��!��J�,q���T	�v���sp�4Im,���9͗��ǭOUt�L�KYw;�:��*��<;C�=��n�0��&T�N��bwZ�����2�i�*�u�xI�s�[:ιb��&��)2��q�M�m�W%��N��
Nܴ�f�ʵZ�f��u�7��D��^
"ʪ����� z��@0�~P�(ʾ��nu��F���v���6��8�]���jq��>+:�]9ung��6�u��olbY��E��T����:��.��Θ9Xsa3�-�c!��n[�k��7���tMMx-�c��Z;0�e�����C���z|X<n��m[q ��n�\�(r�	��ujuuj������8aon4��c��$K��M�v�ű�"�6��ٔ���q[~��?`~�������5�=:2��[v�aVs�' 9�ki���s$�o_�{��}��7C�]��-UZ�;]�6� >m�DD/���,S�~V���ISr���f |ۼ��ŀn�ft$��9�˛U���n7m��{� ߖ�,�ۦ��� �{uګ��kr�G-��BI)滿,��0:�`r������p����mND���_������-��j`Y��`}3�P	v��F�����ԶϮ��D��{��V;c9����m�Y-��{��o����	�vҶ�lm����j`YJ�%T`{7Ъ�'P��`ۻs��8����K��/�{���9m���˻E�؆�Sr�p �v釗���0��� ~��eUĝDj�a*�7]� r۬ ��x<�w�4�_��k�RTܦ��� �}���^�,�ۦ�g�Ѧ�Q5\/�r�;QŤ�K��#@t�ɹ�c��_S��*�m�����n�0�ݸ�n��7]��!BK�Pz{ެ���v�iM�Zr ��e�u���-�����f���h���+�%O1~�k��9Ws��\��`��TN @ O��/�]L\����|���Wn�����B�����X ��^ �7� �f��:��6�Q������ �[�������t�u��?}Cus �]���I��,�z�v��Ԋ��(kb�$�V�T�XJ{ROc�p3_m�57� ݦ� s��/��u�ܧ���$ꍪ�RU�w�u�<�ޘ���,����YwH%UZ������ >z��Q�U���X:���7{�]RE-8�n�0������U��w���G�N��������0�ۮR����(v�{�ŀo����� >z� �J�c���vz�j�9����=�4n���8��g03�cN�1�� �+��I��e������k ���=eL	)^0>��%U5[v�9^ wwnqs�$�����xr��`�78��Gv��v	��H���nޭ�Xy���� w���?ok�luD5*�[nٖ�`Ou��=mL�T�>���H��Yۨ9gr��[����=e�u7� ȍ��1,��*�SD�ھ�6۫,	m	�^�HcN.I�y-)����i)�F�f�)Q�^�B�0����s�k��a�]��-��\v�;99ƚZ�-*m�qlu�Z5S�vD��bi��iA�\��8(�� ����=h�kA&^9���la��mc��z�N�8-�Ԝ���n����z�۞�"/�Sn���c+ �U�	�����{�����������t�r��$(�s�B�ku�\�t�N�ә�UwoRNY{+���Wp�%Tښ�� �{� >z� �M��� �=�{w�]Q6�k�p�[�ov��26��`k�p����۾��b-�9@#����ŀw���q����}�ۀw�U��F>O�j��K�� �w^ |����ŀ~m�J�tm�	XX�x�����}������X~�� �����ȝU�̓�����94�\��w�ص��C��+{<�"�N�8:�� >���;�7�Ss��D(�(����� �uϮ�wSj!�Tr�p��n~I~�l�x�n� �wn{��8�}���[�Td��{��X���j`IJ��^�A[_���^���7��� O�������N�X��,�;�IlL�uWx�n�P�6��/�7]Ӏn���O�U`EW�y�Vԥmn'<6�.�\Q�b��c�8���𖝝d�p�ݧ�U�� ����6��`���ͻ�(\����{w�E*���W��<���p���ͻ�7Sx��%У�C���J�u�^9`Z�x���� �w��/ �8��7�};��*��[� �w]��T����p<�}���]ذ�np����ܻ�]���G,� �V�,�%�}����� }�� 9�f�duZ"J�`��:�3rA&�hܗc���&�N�ٯ���c�Udg,#t%RU�w�u�ۻp���B_�Rwx�,��O��+��%Tښ�� ���(P�L��u��ذٺ��.qq.H����ʤ�,����k ����0$�x����-��$Uʋl���������� ݞ��m����""���^ �fR�V�u�ګ�l3�7g���q.=�� w���;�7��r��NN�&]q�6�#�myҍ�b��:���ct F��i�ʪu�^I`X�x�ݸ���u�D(K�u�8���W�X)�V��0[SJW�	:�`ݹ��8������_���;�*�Yn��ذ�np�Q2>� ����׵Y�:���`s�s�{��x ������zID��~XR��m|��%x�ݸ�K�%�s�}�_�wx�,v����BI
!��r�߫<h|��u�I�]�9(�iݺ1�t���[��DLW!�w$����R���+�uw5C��7p��m��p���#s�a�7���T�c:{n������N�.�r(�6�"-��Ŏ�2��69�N�����=��&��h���-�G���UNn�k�����Qq,��Ƹtx�ƹC��5��e�]V��f�S�����{��uk��ߩ�N1sy2�Nh��b6����pp̝��t�	���LA�=�-m�U$��U��[���� ݦ��!D/����w�V��]թ� ���u�Ş��S#u�8 ����ݹ��s�����ȥU:�S����'�;�ޜ ���ͻ�7�<X��}�[�/˗p���,��zژ�,$���pS���-J�SF�;�$�=mL	�W�	:�`͸��7k*r
�aeU�Z'�ճm�{L�@��ϛvy�ls	�dI?�������Iq��,[˒�2�<`I�� �ʿ��}�\�Q�Ulg,uIT�`��s�P<PV�r��o�\�^�-x��	L�[�UhWw0J*હ��������
e�� �wN _Z�,���VbӅ�&�j`Of�X�M��B�D*���xx����\E�W(+%�z����s�}���{� >���7��@��y	hY��ջ]��@�
��ے���=Tѐ�Q/���{��[��UN���,YqtO����ݸ�j`I��`z�Ϲ���˸KyN ~m���U��xw�b�7i��>�wm��5A8:��� �wn�ռ9B�H8�%)K���	$���@�4 �$�E,���D�H�B0K�tm�����Y��<ـtF��  `X� �%�� ��	!3@� �D��!����M��I�4�		L� K4,��B�bF $"�l9���_C��RJ�.�Q?!��T��@E��qqw6\x�n�������9��uWWxJ"#�Uw��xu{Ӏ�n }�� ���ګ��F��8� ݦ� �
#�%]�z� ~�� 5�� Iw���l*��U-V�]��c	m��'��i�d��:��tv�-^s�5vtፅ����┥��v<��/��w�)J}�ݧ��JR���8�*�{޶U$�u"�Y-\ÜA�#���R�>�ۻJR����8�)J5�j0�ВB�"㺊����W5do5��JR����c�JS�����(}�{��)~�{�)JRw�{oJUS�ȁ����*��A��฽=��8�)C߾�c�JR���|R�ꁤ"J����9�.�y(��wfIB�2��!K,�q8�s��v<��/���┥���ǒ�������)?��|f}��Y�E�[⸭mM�Ya|�!�]	k�Q���p�s�q]�1�3?�ąnew�5A�u9�s�A�#��o�R�>�ۻJR����\R��wv�a� ���6�KSnJ��{��(}��v<����{��┥~��%)K�}���򀙊R�5�U��`�T����9����zqJR����H1���w��JR7|z�a� �_�z�B���9g��`�{��ly)J^�߷�)J}�ݏ%(?�{�~�\R����z�T�!Ԋ�d�sq8���s�D��{����JS���k�R�>����R��W��� �-���s�'�D�w=u{cGF�����l=f�KѴ�@�t$՛�j�Ǖ��3�2��;h*$wm��S`O����Ѻ��+�,&������ɠ�Sd�М�q�&�e��l{N���ktt�ma,:M^w1�v��vk	��*s�M����v)��=�4��с���ga�(��V�zj�Ոي������wj�v��mcFs��a���ik��^�m:���d���x����1y���D��Y����S�����/e+��*�M]�B�
;�z�a� �=�u�)J{��y)J_���S�[��qZEc�u��e\�s�9ý��g�(}�{��)~�{�)L Q��j0����E	�ެ��])���W!u5s�"(�{֣���x�?�~��c�JS���g�+��w�]�aA�u9�sq�8.'��}�)JP�<��=�]�qJT��ڹ�8��[�l�,M�*�]o|R����;����{���)JP����R��w���)<��3����y���s:���݋���%���K��P�C:[Ӯ�tA��nT���)��s�R�>����R��w���(}�N�y)J{���5�7��Z�k[�)JP���cȐMx����VPC�!���}���)C��ly)J{��┥��$C�B�j��qov�8R�>��v<�������┨7��\ÜA�.�	E]��AWw�)JP�ޝ��R�����┥��v<���%�~��┥'���V; �W��VU��8��[��<�R��w���)J^�߷�)@\��ڹ�8��]kw@*�NR�m����čC���O`˫=�Nz\m�s���r[K%E��J��+�q8�s��W0R��w��R�>��v���7����t�B������XIDښ���<��/���┥��ݏ%)Ok��)JP���c�>EV���g�D��%Q�m�q8�s}��JR���{�R�^"! @��jw��y)J^����)?^���Y��6�7��f�����D!;���8�)C߻�ǒ�����|R��Q�N���%)N�ύl��x�V����R�>���y)J_��w�)JO{�ݯ%)Os�{�)JRzW�Nّ=�W^.�ta9-ֻۭIZ�+5��Z�nzy���m�w����σ�ۥru�5��|��/~��┥'���ג�������(}�{��)�n�V�sF�����F�{��)=ｶ���$2S���k�R�=��<��/��y�
"&bB�|]+����Љ��S�\_%)O����┥��v<��P�����o�R����[^JR�n��V(�!+ErY��q�wv�������|R�������R�� %@�@���D ���s\���q�}���"��Nk7��%)O���┥�=��[_%)N�}�)JP���c�JS��ߟ���]���Q58s\Ȓv�]gf��mUu��*0h���U���ܲ�{�)I�}��)�~�u�)J{��?�Q?��Ҕ�����)ǽvs1775%�qD �[?7YR�>����R���{�)JR{�{my$/������5���f�
��҈��m���-z��a�!l��dBq���j�D:�i��j��'���qJR���wk�JS����R��D(|��a�!>;��YJ����Y��R���ӻ^JR���{�R�����c�JS�}�8�)I�h�s��=�ҦDpp���:�]��n)��P����.�5碭k�h�az���x��f��%��L�\�N�j"㚛:�8�s��a;;�%x�p�8�α��e·��lH����n�y���c+�Uv���=v99{nq�got���D��(�̙�����e2.n}�.�u.�]���}�X3S���`�v��]�8[M�btO�kvh:��w|��|n�^M]'<�v3���rМ��ԙ�I���n��o\��m�����.�ͩ-]J&��M,ȆD �[��NBR�>���y)J_��w�)JO{���a� ��ݙ-E�G�Yd��8�J{��y)J_���R���ۻ^JR����8��f)I����6���f�6f���ǒ����}�)JR{�n�y!� ������8�)C߾��a� ��{j#��ƥQ�-�q��$�~���R��u���)J{��y)J_���R��^��w�o0�n���o-my)J{��┥��v<��/��w�)JO}�ݯ%#�B��j%�֣��+��¨�t[��s��=uN"I։���YtGA�]�8_[&����R�>����R��w���)=�N�y)J{��┥'�Iꭧe��s�9�}�ۉ/��@�ӹJL�O6���=���8�"(�ݨ�!B�7ER�UuvM��Z���)JO{ӻ^JR���{�R�����ǒ�������)I���7�W6��n�G�M,ȏ�BBJ?�B����8�)C����ǒ�������)I�շ�ÜA�/�vd�����,r�)JP���c�J��w����JR�����k�JS���s�R���r��͉���I�w+��ȗ�v�5v��G93���]�0vu�B^ҵ���F���}��������)I�zwk�JS�u���(}�{��)�~��쵛0ۆ�k5����)I�zwk����O{���)JP����R��{��R����6���/,�2�y�9����u������ǒ?� I�>�*`�z��ԥ�����*y�\F"Ӧ�V�Ws!WU�)JP���c�JR��{�)JR{ޝ��R���wۊR�������k5�3[23V���y)J_��w�)J?�������JS�o�┥��v<�8��O�U`EPK\�*�h�������w����F�������:�d�v����ѭk{┥'��ݯ%)O��}��)C�{ݧ��){߾��)>��v�]L�4X��3��s�9����/�	�J���JR�����JR���qB興I�wVU�&�.�$�oY��R����}��)~����� 2N���ג����\R���w�*�
��u9�sq8���qJR����ג���{��R��,,�|kp�����R��;���l�ц�k5����)I�zwk�JS���n)JP���c�JR��{�)\��u����h�*���q���U�t�7&n!�n�ӵhu�p��lE͖�t��Z�f����?{��┥��v<��/����|K������%)Os�~5�5���f�qJR����JR��{��JR��{wk�JS���s���M�8�{ޒ��Lv�N��W0R����o�R���ۻ^JR���{9�!�mڌ"D-ctU,�7Ws�޲�k{┿�A�w�_my)J{�}�qJR����JP.{߾�q��v�]V:�?����?�'���g�(}�{��)~����)=�N�y)B)�}Y	���b	͢���	�Wa��s@��7� ,�D��d~ ��j�� ��hd�E�I��������4a��H̶4A�T�Ha%�"�Y�7�nNK�3E$��6�,C$�A	0m]��)����0@�~O��:�xb���,�0��8&=p_�ohK�`&9�RHAb�8fZS@@�(h�1^��s�IG ���	 ��qK�	#��L�3>�mڬ�%��8t�h���
���{L��.^�m\ ������iib�[k �o*�;�㊻VM����'k�ل{A��գvsq.͉�r��l�=��@�`�%u�f��AWS����T��+q�k�5���16��'sa�=p�hV���k���ZlqSv��2^��@Y�u�����Iq�v���l@�R�&T�K;�.m����kz�h�b���vq�.�����m���T�UƤ��k`�]������\�rlʡ�d��x���붮�X�*����#l#vQ��-ʲ1�pl�(q�n�:utԊtkt[;K,�C������FZi5��#R��=N�hF�k�s�v�WP�:v{Y��,�nZ���m��6�u�Y�z	�`�v�5�6��z�/���f����cc]��5�gZ�]Kv���R�/4�=*�Um���������3ʄ�\v��He���iIj�)7"��\��W�@�	Vy"g�w%U5#�/VX������
b����řR�dMe[c8�+����hHj�v��i[	����V�sǳX:݌��v�
E�v\i��6;V��"n.�g��Ӗv"	�#�i[�G]XA�rN�%(��겒i�G������N��l�2Hl��p�x
�,L%��=���`C�������a	f����a!�Z�	P�x7f�r��|x�Bx֢Ɗ���U� nTd��l��v�2�8nf��v-u]{O�t��@sl��us��'v�WAx�m8vڸ+T �e�8��-�r7�/m�į��+M�U�ݳ]mU@�p�Ö���5�vek��;UOmN�D���D$\�3��7�s��R�.(s[��������Z�=�z��d�s';hp�]�S���*�y��F��V���4Լ����x8��ރ�b� �4���+Y2�\�N��w%����߅�?��(@P�E_X����|UU�Oʂs�������5�mu;v����ڞ,���-�֔�����Ƕ�×oNu�hم���ۗR���;.���u�n��&�@4�ip��9�L�Hvv9�N�f�q�7r1��v��\G#˻aP�<u�:���y�X}�W\��ɬ�l�8�
�D�@#c�q\s��g�,/\��������Z}o�i��yH��뮧���w��}ޮ{�xv��炶��a�m:Iݛe�}We
W��sV˳l��u�K-C�*����W�8��@���ڹ������|R����;����ҁ�W�9�!&wz��R�\�R�S�f���)~����)=�N�y)J~�]�qJR����I�C��>�zЅN�*��ns�9�[�/T�R����┥��v<��/����s�8�6iS+U�k�©W2R��D�����┥~��%)K�����	�(I߾>��R���R��4Լ$�9�����\�JR��{�)JR{�n�y)J~����q暺BMdv9%�NB�uA��f.<kT����WX����"�DEOˉs�&d��"c�bt�Z���s����9��I�{��)����(w����s��n�v�v؜�r[��q{���y�?*ud����%<��qJR����ǒ�����|S��8��8����;j��qWiڹ�8R����qJR��{ݏ%)K�������Sv��[u�v���j�L�[�kw�(w���R��{��R���w�JP|��/���\R9�Zn�X4�U��S��W0�q/���┥'���ǒ���{��R�����c�JS�G�_e���f����7E=����;��rZA���m)�kk�^z��dI?�{��������u��芿�{�JO�?��<��?{��┥���JR��{��JR����l�Xo37�޳[3[JR���{�R�����c�JR��{�)JR{���y'���䧹ۿ�j�n0�[sZ�qJR�߾�c�JR��{�)N�T�H� q4��ywc�JS���s�W8�s�w]���r��W0�s����|R�������R�����'�$�	$���z�a�!w�{.n�љ��Fkv�Z���)Iｻ��)��w��)J{��y)J_��w�)@�ߺm$V�ru��;B����؞yv�k���ڷ�-fWiʥ����WEƧ�3-�|��=��8�)C�}�ǒ�����|R����n�y)J{���j�U#N��+�q8�s�ݫ��!������JR���}��*�]�"�P�bBѾ��T�W%f���ǒ���~�|R����{�H(�d���\R�����c�Jx�?�mUB�S	*��ns�9�]��ly)J~����)J{�v<���`�~? � x�wϿo�R����<T���k��㫘s�9��v��%(}���R��{��R������0�s�9�D��J�qʬv<�v�<@����^ŰX��=	�]f��IdT��Y���Nѷ3[��)C�}�ǒ�����|R�����6<��?{��┤.~7���ӗ�t�Z��8��G�ݼ�	�JN��c�JS��ﳊR�>���y'Ȥ9)߯���{7��')��8��AŻ�:��8��_vw��)���{�~��R����o�S�[�u�UuX���뫘s�9��u���(}���R��{��P�.$3�w�usq8����j�AUcOyoZ��R�>���y)@|,����JR������R����┥$�b��� G���̌�_MQ���{>�<M�_�-�J���ԝAv��웆�m�7h�N��nn�'{��kHKMm��͇<�8�؜�и\8\�����Wgof�1�6[1�sX�Y�*�l��E;a��&;b۷7�h�×�"��vǾS�ۗ}�a�M�&U�;��h��<9#rm�Ц��gE�(Q�m�3�չ�Ɍ��֠mٸ[����7v�����^k<�ٱ�uE�;N�'�Q����];v1�2��8��n�\��?�)K�����)I��ly)J~�]�qJR���ݏ%)O3�N�٫f�ek[7����)JR{�{�JR���{�R�����c�JR��{�)Oq~;�iS#���+��a� ����)JP��{��)~�������usq8����B�ƤW�K�R�����c�JR��{�)JRn�6����"D Q�z��ɩ�5�,ݽ�{JR��)I��ly)J~�wۊR�>���y)J�L�ձ�Ud/-eV�^T6�r��%]�������� �-�<�q<NF�Et��Xֵ�qJR��{wc�JS�{��R��mڌ"D-�n�!BO�swe���k�Yf��JR��������uCn�(w�{���̄�(Mf	BP�%	�%	BP��߾מ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP����ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	��}�5���j6n՛�z�n��(J��"��(J3�(J��J��(L���(J���g�(J��0J��(H��(J���(J��"��(J���k��(J��J��(L���(J!(J��30J��(N�����(J��(J��"��(J3�(J��J��(O~��^x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B{���ެݣ7��e�5���pJ��(O3�(J��J��(L���(J!(J��;�����J��(H��(J���(J��"��(J3�(J��~���(J��<���(J!(J��30J��(H��(J�����P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�%߾�g�(J��0J��(H��(J���(J��"��(J����f�[7�-f�l���y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	��}ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	��s���(J��J��(L���(J!(J��30J��(K�}��	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'u߾מ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP�����ދ4k[��pӛ�$�c^��L]%�;��4;%��.�uQd�эO�q���m���	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	������(J��"��(J3�(J��J��(L���(J��}��P�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�w��P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'{��	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�&{�]�٭[ޜ5�nf�y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	w���(J��<���(J!(J��30J��(H��(J������(J��"��(J3�(J��J��(L���(J�}�	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'�o���(J��J��(L���(J!(J��30J��(�:{|뭄Q�BR�j���$�<���(J!(J��30J��(H��(J������(J��"��(J3�(J��J��(L���(J�}�	BP�%	�`�%	BP�	BRJ��'@�����y	B~���(J��(J��{���<��(J��(J���(J��(J��(L���(J������%	BP�f	BP�%	BP�%	Bf`�%	BP�%	BP�'~�����ۮ��I,��q���	BP�%	��P�%	BP�%	BP��%	BP�'~��pJ��(O3�(J��(J��30J��(J��(J߷���P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B]���(J��<���(J��(J���(J��(J��(L�~�~x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'�����[�Y�F�����%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	������(J��(J��(L���(J��(J���(J��.�����%	BP�f	BP�%	BP�%	Bf`�%	BP�%	BP�&w�}�<��(J��(J���(J��(J��(L���(J�}�8%	BP�'��P�%	BP�%	BP��%	BP�%	BR����M�V	�T�mq�hͽ�ZԩnN�����;6��E�rݍ�{[#3]�f��o-�Z�y��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP�~���J��(O3�(J��(J��30J��(J��(J;߾ߞ	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	߾����(J��(J��(J��(L���(J��(J�����y��%	BP�%	BP�&f	BP�%	BP�%	Bck�. \@���},"u���5����(J��<���(J��(J���(J��(J��(L�~�~x%	BP�%	L�!� Ѓ߾�b A�A��}�q)DhA����@��C�	BP�%	��(J��(J���g���%U��Uim��. \@���(J��(L���(J��(J���(J��>�����(J��0J��(J��(J3�(J��(J��=�}�x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�%߾�|��(J��(J��(J��(L���(J��(J�����P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B~���c-��� �.. \@��q���J��(J��(J3�T���(J��(J���?����(J��(J��30J��(J��(J3�(J�������(J��0J��(J��(J3�(J��(J��3������%	BP�%	BP�&f	BP�%	BP�%)�F@�e~Pҁ�D$���`�%	BP��>��(J��<���(J!(J��30J��(H��(J��~˿3F���Y�5��	BP�%	�%	BP��%	BP�$BP�%	Bfa'~�폒�������)I�{ݏ%)O��{�R���Lz�v")!x����\t$Ds7՚��שЛ�)�؂:��Y����3����[��)J]��o�R������R���w��)J{��y)J{۽��uX�d�trKs�A� �����9�O��{�R�����ǒ��������)I���7��ͺ��u����R���}�qJR����JR������wv�a� ���yj��T�Eeֵ�┥��v<��/}�w�)JO{��y)A�/�oﳊR��۾��:6�*r9j��q���%)I�{ݏ%)O��{�R����ڹ�8��]_mÑ�������!�I<㋷�.�����絬q��'Y�h9�l�˹!͹qn�{����;u�k��Y�K�ڰ��d���k���r�;��.�v�&NK��5�
�
ѝ�:�m�kN]�[n�C�8�־�v�UY&��֍�"�L�g��#��'{^�2%�ͨ��8��GDHXz휓�l��ӻ,b�<��*�۩��������V��<k��b-;V.+�����9��(�0Wm��V��:򣫯7F�K�5��R��~��%)O��{�R�������O�@3��)}�����)J���V:�PvYYW0�s�훯�(}�{��){�{�)JR{�ڹ�8��GڟuT�pq���y� R����JR������ )� �>�����R�������R�?��]u�����Z��8��G{�s�D�'��v<��?w]�qJR����9�8��]�w+�X�NI`����s�'��v<��>F}�}�R��wZ�"D#u�Ȅ!=6��)\�n��n;;�6�S�jL�]�胛6Mм 'k��vI1G+��7Zw���IO��{�R�����ǒ�����|P"B�ݨ�!B��N]���Z�Z���ky�)J{��y;��(B&Y�LP�Gb��|���.���R���߶<����s�В��AF��T��7$ԙ�5���<��/{��┥'��v<��2S��ﳊR�=��<��<��wf�l�FkY�{�o{┿� ��w���R�����┥��v<��/���┥'��u����՛���-�c�JS���n)JP���c�JR��{�)JR{��c�JR=;���ژ�G�x`�+Lmv�tf0d�3���ݶ�u�t�f�;��{�q��qu>�u�n�JR��}�ǒ�����|R�����ǒ���{��R�����L�a(RG)l�sq8���s�A� O{��y)J~����)J{��y'ˋ��\g8�ǽ�ڬC��9%��*R��}�ǒ���{��R����`��,�o3�JE1b�҅�8*�����Aa�
	��#3�o-�����,��F�kx�(�y�3�� o(%.���k6� ���$�$lD
�򨯈�z���Ȏ �G��'��
�6:@Q��Ы�������)~���);���{�fZټ�޿�Z��JS����)JP��{��)~����?�E�N�߶���qo����]�Z+,r�� �.w��c�JR��{�)JR{��k�JS���n)JR�"����o5�����&�Ɨ[0�Z�v+�.8���r��q{q�֞K�Vgb3�������m�v��}���)I�{ݯ%)O��}�����������c�JS����ٷ[7���l������)I�{ݯ%)O��}���
5�q�kw�}:7vs6Q7WTI7k �]� 5�xt(JL������`�O��u[8�䒘�IB�|��_u������!(j���0O�������9Ke��wnބ������޿���5N�Q�=w�_fu���Y#
x��^\\��u�-���YPt���Et�0�����m���<`YU���o0/�֒5d�j䛮.��9��I% ���=����ŀ}����[��U�:� 5�x�n����_wb�9��|�ݖ�:ۂu9���.qq�o���ذ�ـۼ�����r)��WW7u�ko���? >����\�@!�DL �F������\u�x�ۨ鍵��x�a6)j���BtHs����gRg�z���jI�u�R����d7(d�M[�]t�1�����_�������[�M*m����;��\&Bom�0�-qv���j���v�;jܧ����ҧ<
[n�Z��\�[2D;q�ي��li����c�ܷf��sac"����y�ӱ�9/P,���]Ow{���r��3s[��F�aӻ��aw7e,�b�=�u�Y��b;7#���r��$�����-�,�@���� 5�x��(Q����Xܥ�)�v��w!�Kj`]��[^07f��ƽz�l����[-�5�u�ko�(���� }�x�ۮ�bm9-�&��q��� ����[S�Ҿ�{4�M��5Vb�uwN��"_w_�:{��oq`jչh�ph�"n���RN��Zr��y�I�&�GZ�ymdɣ#"�J��-o!�Kj`]��[^0-�L���:4�!�#���v`	ąz��P\����ʿ}��`wv���گ%U��겻f��Xnه�w^��Հ~�;��WD�]]�UZ�脗�(P������� r۬[x���ժ�.���_��YS���mT�5t���\u�%Q�R(��A���ݝ[��.� ����DEO�Is���v8�i#����?{� ��q`�t����}p[���D6Kd�7,�;��Y�
d��� >��n�Т"d��*��iIV�I��.��=�_� �������ٟ��~�����K{ZX�V!o�uwr�,��v��	ex��7^��vX;�@����ݬ�B��ߗ�;��p[w�DtW)�#<��ήj4���;��u0	=�v7X:�ݣt�]�:�y$�j��єK�)���Xt���� r۬���k)���\$� ݛ�?����}�\����;���uvj�ZY���#�[S���o[��v=R�ʬr��p?�Ĺ�.I�{��{޼���J�D%j"�%��v�_v붑)Ydv� ��L�[�[S �T��VwbF�T�b���uqv&�y��%юͷJn��C$[߫�{���%�fr�_����I�}�?�	mLIS �����ZX�W��Wo-`ژ��-���f��>}�� :�P*r9n w�� 5�x���V������x�z;K�,Zwoj�GrL[S��� ���$�0>�w�ӎGjԐ�-I0?:npDy(��� ww� 5�x��_�2@`(����������t���]��ڳm�x��e擋c@�i�����HW�mw($i9�l�;A��,�q�v�P�<N�m���n��}��z��շ�d���a�7��lTq�����n�[g��F۱��B�g�oX2�v�an�4��Mɶ�)ݮ����6��]u\�,�Ic��	&8�׭��#���]4�k�
�i'/dɒ=Y���9�	M�fi�����8���Է�t�<���=ay%�=��zOa8
l��� .�9��$������o-�O��0	%L[o�_�}��< ���򔑎Uc��[��w�ЦA�u�uwN kn�R"���ob1wjI�Kj`}z�`ژ���}+䑽�r�a��o$��z����	mL�T�%�0/�֖-\bոM]���Kj`��-����u������X�Rζ�'���O�GgTQ��d�[q��֚���y�XY�"����{� ;�� �u��%�0>�
�~�N�9g%�w�ۼ��D%��{M� ~�������˽V�r;MIwo�J��%�0IS[^0.�ӒĐ�(�*�UY��
e�u��׀ko��u�|[�s��o.�rL�[�5�� ������ �I-U��Wa;]*\G\W�����^:I�`�Z�0`�멡.�vj�zr��uq��7O%_����X�M� kn�� 6��kʛ�;4��������]�P���I?�[^0$���1j����Z���{�U{��/Ey(� �>m�\%۸��;� ���,,�vGȪr���w]��ŀ~t��z!$�L�{� ��OUy*��	T�����X(��� >� �u�����hY�I��j��nY��]�Ү�ŵۄ{m[�Q���L�[4�g6MM������~k �T�=%L	ex���NK,]�����o-`ʘ���,�N�XŽ�9�ڳ���&�*`K+�ӭ�,��2D^BY��\��0%��ӭ�,����^, �J�x`
�߽����}܎�D�B�g������� w{� $�0%�����ڷĿ	.޽-�d��X�t�3zN�ٶv�@�1�8[b�B���]���K*`Z�{t�>ٺ��{��؛�8"�#�0	-L	b�׭�,����U��,Y�vrĄ�`K�n�	eLKS ��R÷��-K;���[�YS ����*0&�NK,]��w/ۼ��K*`Z���ܫ�u��*��V½X��JL��F�]��&���X�	�ibw@�И0�R���$!c@E��LD���4�$$�һb Jm��1X�Q�oZVb"X "S���� �=��������m����6�� 
�������5���&y5�S	�dv��WTg0O$�+B�O5�^�g8����+���@�J����A�r�`]�խ����ӱ;���������4�5�Ys]+=��2O+6S���v���QEKx,-���\ZT��V�=e�J�m�v�A&$Wm�"�#hܝ]˴�m�4�c,��"X�ۗ����ݯ.�t�I���b�]����ܑf����F*��q��	��,�����S@`�55^G2�c[r���t�Fzw6�CbH�w;Ld�Q��Z)坴q�7^�M����<N�gN��;�ﯠ��n��8�`�1�4���C�&��m�UI���[�gC.ӭ8�:�[vl�n;h�͎;f����u��mq�͝���-��ܮ'���Uv�T�y�4�z+�[=M)jn�mg�A[[F3��ix�s�ʽ�H\���QV�*ӎ�K�e�s��P�$��z^&%XغS%z�����3J�nڧh8��Ma8*���.	y��^�U���]lcc��W��P�T�c8VM���إ�ɚ�=n����e�H�B1cͻ-��m�u�um+�۔n
A�3�Ln���9�e��:���c����c
�u�cZ���%�s��VA��u�uYQ�Ik��h�b]M`�ݣ��9xŊ�R�①��v�(�kb4l�0��^^��ۄr�����NƯ��}�|��ژ�ض�`��Zn�z��Ms�f�n3X�]��z��D����7m��5�\h�"ܦ����O}�o\e�GR�n�����;Q�ǝ׋q=�c��6���+�z��u��i����c���ѫ�"�@�Μںڪ���Q*S�;/�6���Wf�N��T��q%�k8�qu���G̋�W�v���[�q��ͳ��e^������L�g������=fD�l���m�yv��|���8vY]�q���m��h8���[
�d#@�qu�\ sm�9g),6�S������"i��_˂�x��D��~t��P����w�Ӄ���	bUT��.�Tpb��ɸ��-��Kt'tQ�Gs��A�˾�0w���v�q��6��sϵ�U�g�sK���n�x;.�nmDN�`،�����ې	����]T�"nX^�=�pl-���t�p�����jv�s�ͧ���k�;(�Yx��{��u�hB�ņ���N�֒r�:��m�V l�n6q����~�]c��lmF9]x�ь�p]�Q�L����Z⺞ �P֩{V_��2<R�HU
�$�����\�ۣ׭�=j`L�,K7P�[�+���>{l��M�0�u��w�IrC�������US��,������� ߛ�?�L��^�O� ��9J�1i�f��C ��0	-LX���ĸ��g�����vGT�� �n�(�y��7������?}[����M�B	�����ky7:�H	��K�R�m�3���Kʎ���q���RLX�����z��$�0	7v�W�]�HKL�ۦs�\^\\B�����Q
�=}���z�u��}�%�ʬQ�K�%0�ݸ%��,T`z�F�om�Fwp�r.ʫ����$�*��z��_���=j`L�,K7P�[�b�I���Q�OZ����ue����u�gy����x�iM�9d���m�gɮn8�U%vxMu���_o������ 7�� 7[�(�
?Ho;� m��ą�7q`,���`֦%�����}�t�?};�Q؛�8"�%�� n�x�m�|�$�J>��S
!�eEԦ
&0��f��\��ۀ~{�j��^9���p=�qqq���	�����'�LKS �uH8����$%���׀�\�8������\��� �f�D���"�J<0�b��Ŵd:uv2L�tݱ$�t�yv�2���rU��*�&5%�r���z�e����n��z����_�,,��� �n��(�7��oWt��j`L�]Kf��q,[�0=b��M��
����_u��ʛ�D�uY\�Yn�����< ��� >����%}�
$����9�We�dʴ��j� 7�� �P�N����0��L����G��;�m��<qY!c���+s�"V����&�׳GX�ۥ��8��v����0KS�W�N�X�����U��,_��5bKRLYq`k�`������D)�z뮂Xʣ��`�_߷n }�ۀ}��X���j�[���L ��0KS�׌N�X-��\�^[S��� ��� �;�{��v{� 7[�Q�)(�Z��.ˋ���\nQ5`��4k��R%´�[R��BO��rX�	��q�������Y�c��is��{s-�O6܉"��5`�ے{;�%x��uy��Q"�5�F-�V�nM��f�p���EG����� �1��ݱ��5�Ƒ�#[#��t���8��jy��N'y�5ml\A����%g<=D�;�i�@�7s�쌛Ep�����\N���K�0���"����k���N��HN��z��B�d5��	���S@]��WO��q,%����<`zu��$�0wv��׎�T�u;I�31~�=��d� ��xͼX�s��ˢ��X5v��%��Ij`z����׀}�;����N:��ۀ��5�� ��s��(I%2�������@���Y�rI�,��n�	eLKS �.��9gr�o,KV�r��3lD-��qVi�cn�^
���v9}�rR�ӎ.�go��n�	eLK� ��q`O��Z�V��%�r� ׮�%��u��5�� ��s���/�ؿ$�Qܒ`Z���Q;��8 ����m�ڵJn�E��-������ �T�$���t�j*q:���[������ }eLKSz*0$˕�nov�o Wl]��]�!#�dZ��!��+!v���k�����9dV�Q���W���pu��7�{��_t>��n����ڳ{�$�$�0'��֪0�����U�� Y�v,�9$��W�w����RJ	�
2� ���H��`Z��:�.Iwoor��T`[S ����W�	�.^K9!w����!�}mLKSI^0=j� ����uӅ����ˤNk.�a �h r� ,E��D�PR��Ec���H�-��Kn w�� �����T`YSH���Yػ�#q,�����U��%���wLr�N+i?������� ��S ����W�	%}ؑ� Ŝ��Ww!�OZ�����fffv��s��n��ݖ�����S��pu���ŀ|ݳ ���+����:��N0�N盢H��d�Ӷ�ۋc�qr��U��=tn^�sW�����n�eLKS ��K�E��q%�or��[��S �v���X_ul�KK ��
I^ [*`Z������ ���	g��勳�$�$�0-��׭�l��$]{V,�]�����`[+��[��S ����_ؿfp�I!q�3c�S�Һ��W�D,�����m�%�ƆW�ӻF[fܲ�a��6tf��)�7]�ݺ�&"��ݸar�5!c<j��5�jŤ�&��Ǖ������c�ۛ�S.��\l��veiݶz�����k]�!c�)�F��!+�l�!nr�<7.��1w+���ǮRGl�{�U�.����F�F�
���Q��J����
�3��{����{������lg��^p�[[C��{<.�]���l(V�P�&��>�e]�ݮ�HV?e}�x�����eLKS�^0$�_bB�,�ݺ�yk �T�$�07{���n������FW
����$�0-��׭���0>���*���	m��q%�.=���w��8�m�DDDDL��x�뮂���椴�\������� ����wq`}��TD��J��u;]Dͣ�|$���{��xۢ�)�\ܐ)Ӯ�n��!vq�ڿwr߀-��=�H���5�Yv�qرr��Is ���I(�P�Q��,�M���� ��6:���%�� �wq`l�x���KSz��X,��v�o��o>w���=��`Z���`I.�ą���]�����y�Ij`zt����u��m	P-��X�j�ce���"���o���Pm��ۃi9��wl]�ڥ���\|*v�f w�� �����n� ��ۀ~{�j����"�B$��.�=z�`KS �������w��eV;k�X}=�wv��j�]��o�0	Ŝg��'b0&`��l!������P��@a7X�I�ڻ�`Fd%  H�$"	�b��A�	���dR	�)I���o�f�~��L�I0�$D�C]�c�� : ��X8�D�`�
a -��C1�I��Y�4�<��z�7�7�k�p<s1$�\? %�~��\l�s��@♶_�:h��<]�lC!]�<l�#8�*��
".��DD�f�#��1,VgG4��P�l�<U6l��*�����~Q�A(8(���_@ �r��k�?\��q`}ղ�%V(9䒼���^ 7�x��,ID�_t��?BЄW�Ub�ۀ���?�;�����{� >���>O_V�8�U�:�-�齐���K.V:�3���E:y�Z�;��e�Њ�mL�G-�>��,훯 >�����u�{�f�)�&�W�U�/�oWt�����w�}���(��/�8�����ZXTVJ�,r� ��ɀIj`zUF�[��ļ��{��K�`Z��Q����z�x�xoH-�U��g�s����j����H�����ۦ��Q�}������� �R��5(�U	Y��җTmvz7!8Jè�<��3�oW)�Rf�롩��\�k+~�߿����KS ������	��䳹+�S5UqUW8���"&A���7��`l�x���Z
EymV)m�%���U�n�	-L	"�ڐv#�#N�����`z���$��y.q��z�ｍ�Pr���s�7��pu���� ��� ��?��F  ��HT���&Ţ�#��RX ����{���;m���}��F�8��QGb�]Xr$>v�pլ�;���1;ݸ�7-��]r0��ۛN�l����̥���˗X��.0����
�FW#pH�� ����36��;���۷�-{X˰̓��E�-�jه=���Цۛ�Xɱ�
i��gQ!��v0e������C��x�*�abrTܿˋ^c���E��=^��;v� 6�^3m;�C���yMD��eGX;]���QY+�������pKS�׌^�X{�y!oi�{PZ*���u��脦M��X�wN Ij`}�b�رi��w�`z������^ 7�x����KA�w$o��n�	-LKS�.q>��� ;�'�����I+�	-LKS֪0=z�`[�l�̈́,���]�끽a�kZ6y!�<󣣢�r:8��8���s��	:�YÛ�} Ij`z�F�[�KSH���ȩ,�$Q�p�n����$��S�BQ]����~� o��u����͡*����}=�����Sץ����嚱[�.�Z�'�LKSץ��[�{�e��q����p������;�����x߷n��n��qWev�DP�]v�W=�<�[%�68�3�.���=cB^T���*����	-�>��x훯 '�LIS �T�h�۽ܑ�Ik��� �Z����K��3���{Iꬪ�$w�J���� w���~A6>+�b��{�{�����s���A�-�Ib��`J��.�>�n����$]yrӱ��������������%��� o{׀�v�t�Ǌ������d�����Y��\<c���Nm��rk�q��<��/]�n
�DTrT�L����� ?wv�{ݸ�K�	%g,��b[�.�C �Z����K��T�ٺI���v��a�rL����.�>����p�zmW�TT�UHIn�ֹ�?:np��x����IL	���v���mZI+-� ���?���z� ��^�ֹ�=�����jJݗ�hya��⍎�N۫W`ˌ�˺�J��3d��#�	�g7kf�⪮ |�� 7u��ֹ��!�u�������"�ۀ�v�vw^�f���ݹ��7v�KkqRX���Swx�}8�M���d��^ n�߷q�B"*9*?�&c�ޞ��������(�:����2�,��b×v����>��$����׀~ݺ`%����q��jlv6vݗgg<[b냒�8�s�ҽ�c��\�rMZ@�V.Ųn@`��u�����< ���BUƝ�n&��3������m�]�h0���v䶕cpdɮ'M���p[^^c�s�Zvn�auJd�=�����_�_�*2۶�\!����4��m��.;l����ݖ+��ځu%E�{�Ȝz�:ά��Jkvc�`�>ng��{�椖s��LN�"��ݕƈ��Ћ1�t�T5Ĥ.cF.�\V��<�os5��uƙQ-���w� ����۷O����޸��z�Ȫ*NHIn�Z��'�LIS�����H!hE$*p���z����p��\l��\�����ڬ��$w��0	�S �T���u�����xH1%���wg$� �T���u���u�OZ�&i..0�Y�7[x�Җ��������-S���:�����Na��{[=�f�h⤰)����o��v��w�B� 6���왻
E+�����\����yR]���K�I*��~�0ISץ����9f�ܰ9wIu5s�����w���O� ���X�K܀]�����7�����T`}z�`KS��ł��w�0=%x�����>��$��_�~�#V��6��,4��6���g��Ե��^�\N��Վ_!)JSVέ��Vo�^�X���$�0=%x�?oI�YU����$����� �eLI^0>�n�=���A�-�$�U�]���>�x���(T�%tM�W����\��%����R5� �u��?:np��x�	L�����nЈ��%�y��������� �{� �����^^�hԑ:ݒ��kb�v�7=�eڸ�\y+���^"�M�4dd��qإN�T����w޸��n�k�֪0>�K܃ui��3Vo]�� n��IBS&��X��� }�� ����yEI�Td��wn���tDDɯ���׀v��T]�IUvMv`rI%��}��0��x��|�
��V�7�w�ܪ�V.X���������=-LIS��׀~ٺ�MO[$�B·%�����qr��N�
 i����!ZT��2DX�U(��j�	$�i�b��I�I*`zUL�v�(�I{���xw]z��WUX�Ԗ����?�l�޾0��\ �{� �۸ݡ�Z��yp�������I*`zUF���9f�Ҡ��쒘���� 7w� ��t�?n�0����ePN�-����+�Q���֬�۷�BTW��TW�����TW��QQ_�AEE�AEE�P@���T�����������
*+�
*+�(���
*+�(��� ���������
*+�H(���EE��������)���y�����8( ���0��� � @
 
   
�    
      9�PJ�AA *)TR���
 H*� )T�(J�$
  (H��	� !D�J�"P�*�   @    4
� >�o�����������͕���^��9�^�w���o���9 ��4p��\ ���^�\���zS'�ww�ݼ�*�s�{�@��f|���U�'m;�^   <�  P
� 2 ��iqx�{o;t���X�Mox ���ɪ���,Y]\λm�Ӟ�b�X�� �n}i�ӫ��G�K>���O�^{���+����3�U^�I���z\Y���Y^����  |    (�%@1 �}[k��W��nx�=���,�ox@;��\Z�������{w[� ��'�U��\��6�t� �+���t��{��=�S����yS��{��:����.�N�^ �  Q@ PT� ��R���۵y�uN\��;t���)�R����׭94���   R   �W�wO| ���� 9  �  P"        >� Q�� @(  �  �@@�p 	  � lh D  (� � � D E � D X   f z��ϧ����}���iɯ��������>�==�֜�t���9:^��>�W�OPL)R h?�Lѕ)TC��Ǫ�T�  =��CH��� �S�	)J� h ��II �)�2�;��~S�������5�7u6��~i�2fd�B���E�P?�E��E��TV"���������␡?�bCe�6����%0H�!T�pF+D�Ī2$k�e'�C�y�&�*!
�7�Cۆk�
��Lȴ�D��M$9�by᧗�`B����	�`� ��-Ii�
aR.���yY#\&y'��H��&�F�?�q��'�$hB��ļ�{&b�!���Ɯ��B���J��!X����!��O����£��q< P0N�
a����)�Oe����Ϛ�L�M���̆x��|�a-�|�a3Y�$�5!J�*�!
aw�}�\���(@��+���ÈF�L���"B)(9��v�����LB�=e͢W�1i��rB�H¨T���$�X48����y���h�q���hJ2�JJ�� ��b��F`Lu8��k8R�&�*b��RH0�Rd���n�±�F$jR!�0�b[rN]7���D FT�H0 P�m"H	 2(�(O7�0�4�8�X��
�F�델o�	w�B��@��hSS�B�Ho%$�LM#L5bT�B%3hH��%<э
DXF����hi��`P�x<CL*JT01�3�y�	���`L1)5�5!\4��X�����Uu�[!
)M&&�%�dSJ�H���=R!F!SЃ)��	r��j`�^�@��/�$a���e@�x����]������.�)�B��Z� �H�bЂY]���
`���|�`�g�ė1�0�f����=�e0%�\�0w<��	��<p�����p49y�a��/���I_XC\4!sL�=>%�B,�i�0�@�o\��hviV��/4��׽uo�f!�$"p�q�)F25�S�� 5HSy�\�(W��\n|>�k=%�!�V��eącFYL�0�0�4#x\�(B�
a��(J�x˚p<X� ��E�sM�7B%e��0�an�.RJ���sY|��spHVB1> �X��@*�V���6B�>��h�o<)�$J�M8�xB�:|+�R�Ӌ�B:�% ���>B�j������3 hK����Ҙ�=}/4!|�$��{�\} t�퇅�<2l�f*
�J��3�t)�ʎ��i�F�:��-��"SB��.����Yp˲�J�_Zpcx>�B��(x�
a]8x�i
`;�rd<��	��e�y��b���&�=a[ωp��
����\�0����s�paXP�7�x��$ጸp�_��i��O\e�y��p�p�#p%1&�y�L���n���.��O�B%�`11=���_�]41������+�ǫ⸼��׎8���Ӊ��Ec��!^�Ԭ|��u�8�X��F\�35��|a�݄<�Ja��nl+)<�|����̸�0�3|�~�8�(D���
�`l.B��Jf�t�p`ԅ���\8��gĹy�.m�%����f�(�����s��ˤ7f��7n�HM�]6�p��0!R�"R\�p�t�!#L7@�L�s�y�D�^��IL�0!BP���BP��%�x�ȱ)�o'�p��	r]��i��r_%�BS%�!L��$9�K��<��7aL�HSLcC^���)g��s%�h9���
iC��y�����Jy~��<�g��F�bhhB��	ŗ~��ģ��M�Ja��F$'ia�n��¤�c5xq��R3��Q����5��'�<�K�n�
B#"�$!%2��a
�)���|B��0���x� @'IBDzU���XT�%*^x���hi�<%0Ӟy��379�{3�3�ہ0��<��}���Lf�AH�X�Q4ޔ8z�@&�a��W�	Ni�%2��|\��|���X�5��}��h�hz���Q�8�
`o�C�&���H\�Bp���0�(�]DЂ"W8�B�Y�n(�#se%B@�7�X�q����4S5$�3]� P��<)Â�>�l`�ŉWB�4x�3&Ȕ�4cC	G��i��� HT H�H6"�"��P�q6��}�hn���o���шW@�\M[H`i�B�?��z�bA @bBe2di���F��hH�)�j�
V$!4�W�,F��t=+-0�M�8�#
D�]�����$��[������	���0(��j��)y�&rp�%!5�pҍ�K [M�D�4�U���kĆ�B�$Ӛ�"F��IsRV�*�L0���d�0�§�xP'!#� h�
F��M��s�<� �, ���Up�##��`�@���`��8���@ ��	�@j��H��T`�P"505H, � X�L�Ih�:�BH��bP� �#\xJb�' �P�u�� 2l��|*f�$�S �"�Lt�BIp7IH��cVXC�
Lk8$J�|3�8y0�p-�\f$hIC$�.M��s���
㧞1µ&&�=��J8��}=e)������e��h��HVc\HP�Hdhq<Hb]0̴Ċ�H� �X�:��\�� %����B���<����;%�5�5�GC�H��t�3���L!��V
'�d����vZ^��*y�#�+ǁ�Į�5;I+5�G�s���&_�f�|���Ja�>���97��ӛC)�>q�cLM8z�����眞���wg1�FD!��� "$�����"B�`�I����3ͬl�����$4��O���<�l!)��.o���ǧB}���2��o�ǩe�k#hS� A�X@ �!�B$B�0 [�Ĺ��B(B��80a���<%��x2���NB�J���/�Oʱ�Ha����,��LÇ7�7rg98a|�8����%�%bŭ8���
�*�B"Dhx��B���
0
Ħf�� �n����L�4��0g1�$�$�L3RA�b3f���J[��ICI��VS����Bz�,!)�Ѯ0B.��K������ŐBDK> }ᳵ�i�!�>6���SU���T0
�Ȝ�s%�$ a�B�/-$��ɛ#䡁�)�����0bFl��Na'I�S�
�P� S�	Q1׏�z��
��o=g���L5���N{X����Hp��4��Pb���jX�@��qB�;L��
����i��Je
�y���Z��I��l�=�g�0�l燫��p9���]��5��hf��t�B�	 �`c������ �.䋄a����Zhy��D����(B���7�ۛ�w�	%3���Sr<��C&2ɇdhW���`x�R�c��D#`s)bX�#d��m&�! B�� ���Y��fa�4�I%e�˒�-�k$�
�I�!2Y�h\3�X�g$�<}}�5`ǈ�b��< ��HWx�`KdK���3������IL�RH��鱹�4�s���Kf0&�jh
 D�h��ufn�N:���$+��h��(�qP�cKf�a�+%޻�4�u�� ��V��Z�#y�Ej�*ĀF��`i+
��K!\_i5�F�j$J, #��a,����I
FŒD�2��VԤ�d(�HČF�#)�$a��
0)������į���,地��6$Ha�g�!sS��FL�q�<� ����9�      ��  �iv������Y �bVb�3l�i6��t�E d�m6��8m&,6��}����� ��uU��qR�� �Ͷt��ٹRI&�����@�V��F����类����6���)�� W��j7]J�^`�N�]R�L�n��UWl�
�����ب����; �TcUUWi�K�^f�;g\)ٰ��m*�d�(�7g\� �d���ٰZ:�������mm�B�$ 8I/ZE��nٲ��� $�h�R�P��h���ҕ+,�WV1u��g��ǫ��l�%���n��R���K*@�4�dܼ��UW2� �5�@�˥��l�Vm��j�� ��$�[i$���:x m%=I)�6݄��gK$�H.h�U��H8�uT�6]�H�j��d�6��Y-��������Ո� OJ�U[��V��UUUګ����@@Pt9W�$� �_,UmJ�Q�R�!�+-l��L-WM[������d��2F�K�=P'�*��vͧW�&��;n�VR{9�����xP�Ap;V��^��]v���[i�H���&��ޚ�PAe�r�m���5�mH���ݰ�@H [@[fD�nD��p   ���5�[Kkm�n�8 $��vU�`�]�[E���h��l�[�(m��!m���*��M�H6�t-� 6Z ��U�-�j�m�^Ӳm��ٕ�K�T����v� ��۪�с��H ��y����EK��2��]��zw[���k�۷`s����6��Jqs²���Nku�`88+�n��9�� �V�Tɼ�uu�ѭ���ZA����ԴK{+�-������t(5��\;�s���G;iW[B��}�M�yZ�l��`{!\��WR��(���ˬp��z츧��٪�WdN�T�H��ٺ�W2pn�W(��yUC8j��k��V�xGM]:+�j�ʱ;����8�nM���@Fٯ7ekJ:���UJ�,q.ݲ���:L����e�&� Z9kՔN�S�r��=c�D��]eW��v�rִ �&�Ě���P[m*�UZ;���Z�^t�k�&�������6�	gP��6Z�	n� E6�l��� ���k��&ڜ�P6�&�6$%yj�x�l(3�:� �m����$ I�À'��X����  ic8$qm( � :�kikI��.m"�H�a  pUUTH�ݲ���T -��~P� kd�l H"�[A�ѥ�:�����W5lj@ �m�d�mz����6Y�5C��ś ��"��m���lH���.�(q|]��.�S�4[M��� 9��$��v�j�ׯ�"Ѕ��K���ѪV�V+�bth�m���h��e�]� $ �	��[%,kBKz�ڶJ�H�#N�t�q	�Jm�O���$� ��5 6�,�����i����m�I8p�H�� m ���� X�k��m������F��\ĉ  UU��U��%���'�/-K�r��UUR�� [@��$mڶ��-��3�� �\��V�r@5� � [m��8�`�6�xl�m��E�X�z�
��]��ʖqm A&�[T��nE�*�(��U*hXwBg����m   �����-�nvր,��n������ �	e�����a�ݷ`�v�-��m����͑"�탂ްTֺ��-� h	-���}�� n� ��n�
�UV��ل�Z����vt ��� � -��Г��b@�HU��&� |7��bB@ ڶm����hm����m  kY�] Ŵ���6�v��À�M��i��#Gkp���"T� �m׭ �i �մ�;`�I5��6�p��#m�!m8��9)�-6�##�����)m�,$>
jޮ[%5�&I��kt�E�m�y$�Z HJ�;gDWUW] �l�h�,0 ���ɏ�5���
�#��T �k*�flK+k�@[N�p�� ].mYֲ�R�󱝶{��F���8�� �[p-���6�  5� [yKU#��g�t�8�F�z	���:�Z��
P8 �K��vӢ۸��(���#Kje:e"��ݹC�Y`p�n�pK/� pk���D�{`��٫[r���O�[M.m%���NIJ�v���T�*�4ڶÆ�cښ]�fr��m�h[[;Tۡ�8���؋��� U�I �-�I�m�ɶ��n�`�x�̗)3��vsȨMT�횪�Y�%R;vf�� l  ��3E9�4� H/CZ��9���۶H�ʪ�@Us���[�wPW!�l0"G[�٠ �6�@ I,�m�gD�:�m�  m��7U�Ӝ�����$8 �l ��:Qem[H m� m��� ��5��^�6Uz� W+��[��m[B޼^������ n݇	 5���/�-��@�np A�	-�[m�� [Cm�@T��J����<������uݵ�����   6�#�%HI � m-���D�;[��N��@ �  8 �� �v #�J�&� -��"Nm�!:H��n���@   �R�6�ܖѷH� ��\�v�5�`$ ���6�Ÿ �n8�v  � �p�        ��� ͳl	 I�  �$Hm�&3  8��HH   �M��ҷ �́ �u ' �ͫpS!�\]�sWe���`*�;5U���   �y�tƉR�r�m�   �   q�&�\�dȓt鵽vm�okp�7K������l�[o`$��	�K!!ͶH  [@  ��ݳHC8t� Zl8   ���D�U�c�l�+�6�6t��(6�  �]w/�[@I'��*���n.$��l�n����8۪Ci�v��<rQ�Lb�eZ�k���`��/f�[Al�m5��6���~��Hc���gJ�Um m��"T���: �!im�fک@Wl   [Sm�
�t�lU;+[:b�T��J�\�v�m�8�`��"�U���d78$&��L� ��}j��b�:��`Hi���p �xu�*D��[N;m��m�m�@ 6��m�h|l� ��r����iV���9ٻ.����j�Z -���E�� m8s�'I)��I�v� H��$lۖ�  ���@ I ն� � �Hf�� �j��	W(�հT�lA    ��N$e@���yj����]n�Hm��� �I�^:�ݶ׭� �   $�	 ��  < 9 6�z� p m��e� � -� m H�����j� �#j�  m�  �5��m� Z���UW�jU#u�&�v��h-�UJ�Y2J�Q�d&���Z��K�U�l���Uiҁ�� ��v�m�   >� [R���9��m�Jm��!���` 6� h     $�m�6�6�MT  6� qn�q��/V�c�Xb�J�s]K�@+�r�`�ئ�)*�Z�vm@�d ]Ut�K�!�d��a`Q�3\��UU�Qh �    5�N��m�%��6�8$�j��I�$�  �&� ��# �V�5;WN���/6�`V nݳ#��$��M�i8:�jk��m }�>&�bݝ��[ZrK���Z�{db���!�K��8ڮ�;,�6�L��%�a�}�IS��.���«��o�:��?�0 vv�I��e�	/��g;�Z��n�+eٞ�n�-�pg�ԫ� ͫT�s ��6�]\o�ﾮ�R�k`*���W]J���� ����M�a��.R+��ږ�85YD
�4[&�ˉtEې���$�u��T8�u@E����uAKKt�(Xv��9��"G+U)-J[d6����F�6�$�$5�l��.�r@��|,�m�B�$  КL֨�P#�5WUl@튶��z�o��}�IJ��hܽm�UP p  	R�]k�Y��X�`6�[% 
�)j���-��&QAp[@m�(���h]4�l8��IMo3�m�Dڀm�� `� �Zm�m$�C�ՂDCvdZ�
醵� �  ��]	���aͧ�N�]@}UUT�J�s�툖�^m�� HKh:J�:[�[h�s�ڪTai�8�Qy���Z�� ���햻Q��
�7g��B�j��R4v��m>�m��UT���]Kka�?�w{������VE�(H'�EpO�U:*�LB" S�����jx���	��8�G�tR T:(��U�	��T�1 ��=T�"�A 'P����R����b�^�$BH��2B�	"0$��P>@�h����$u�PO���G�� G���U��� �`>��A>��E�=Q�����,P��t\�$X$ �R DH*�$`� 0dE^�5 0��A ��*��x�(z�� p�.��pZ�u�US��AW�/���=lA�W�D:	���"|��TP�LDB ��AP��P���Uj1S: � ��MDT ~E47�A~T�j�u��C�� �Ԋ#�����x���T�w���E�G�����@+ ���337wwd�a�̲[t��Lh��ͻ3��l򽧀�yd�=]��yr�N��@+���b�먧q��LUm�7[�NW�X�3��V�m�hvh���ɳ�/gk�ܽlʕv��s�mڣj^{B���-�S�#���\�luq�*��s�pm�i]0�U��/M�|m�0�`�ul��85���9z;� -�q*XU�M�N͍N��DZ:.��C�Nd6�^S�;u�#v��=��=#��=��T۪V�h*�ccP��u�%����s�]���U�ʪ�E��L����k���X��
�V-���6v�lB��Z�3��LHrm�mlD�,"�pYtR�*�+��]ݞ^�G��i�n�v,�T�ga;sċ�qЯJ���q,�LޱÃ�d�7V�!�&9��=�\
I�l�nwc�U�7Kų������ˎ|�u(��-�-�w7i�Rg�s�f�J`,�]̖Ӗ�������^q��`Li�5:@\{ �6�î��Ţ�,H����l󦕦���[�^�ʨNZY��<c��U畯�;nu���g\լ��
�Q��]���#�^z�[2���L�KU��e�:n�d� $檪����`U�Td����Y-n4���:
��i-moZ��H��m��M�{q���j�<�{<�W��і������í�:�l�������ۄ�-�4[I�g\��$,�F���ɺ�\�OAf�JD������P{%.E,��֠�rˉ��.�Y���j1������g�,�f��ZJn��!��m�F�.ң�H-���z�H�����@�i���Z�%j��W�ڮ��sjL���	�ݶ]Xy�]>ɵ-���N �r�[\{�ڸ��.09�nZ�d9!#a�f��x�a�����<,qe��;v�%��gn:l<�ت�]�EY��M��+�n�A�N���� H��5�t᪔i�ٛ7p˻������B F"��"EHA��BA?�� �����^| x!�	��ww�~w�߻vY�6{*3ù��eaz�4֦l��뮂�dAy�J�s�^}R��{<ԝ���wJEU��w.�{s�G7 �֫��8Ν��7klGnƶ��u��;�	@vzq�@��s�=G+��7]$@��D��pݎ������ٸ�Eɘ���v۫6$)YېB�ͬ�uOU�^ʙmF�U��=
'�3=Ҏ���.�{OG/g�TUT^Ó8�xLgs��x�L�݇Ha@�Rt�T&�u�H��l�fD�^���$��v�M i��Dr�p��t�����O>�w��Qz�d�����3w��9��`n:[���:p�I��by�H���7���L@�Ǵӏ�RQ�$�`��`�l�f����]ǷV#3`�"��{.���� �1 k��*@ܾ�~~��k��/^�Nf��u�)������/;^ܡON����{6��n�}�K9X6���aw��5Ɉ�@���� 3���9#(��&����rie}U�(F ���%@*�!Bd$��&^I5x=����l��vX�r�q�����`��`�l���zX͞,�M��d���~33�5���@�� �M��Q�q�CnI`��`:�����@�bJ�=W�z�D4�/�m,�h��:�	�
t7(�U�ẗ0��
9)Pt�R�$�9ܚX�1 o9�\��6��W�����G��~2�@���� rby�-����̓c����J'%�w�wy$�}��&*!�bFEJ� R�H�`�JDd�$�/32L�^�t�fl�j26�'�Q�f�9ܚXs6X;�,�={NH�*8*I��7�A ss�5Ɉ�~���J�Q�"�#�*O�j1܎7)ӗ^��mۖU���wl��1�{v4��3�ݭ��gl�~�8}�� �1 k�� ��]FA&ӓ�I,�͖�ݖ;�K �f� �U����:N8���b �� 7�A��~���b �s,�Ku��N)0RK�ɥ�}���I'�����Ah��1��Uz����sy$��gL����(Q#��gse�s���9����ri`���	����7 :Pκ�pާ F^����V��'vēe�\"����ƾ�͵
�	��rp�͖�͖;�OUW��`{)��p@I�TA�b �� 7�A >s�}O^Ӓ2��
���9ܚXw6X;�,��,��I�褝(�� ����>ss��69��s��6����$�r|I%�s����.�t���z �͚S$$&L�2��X�Z'Vf݋1u���9�qˣ�x{]R!V��6�^z)�j�k���ܒӊ������HZ#H���/��.���ձZ����ѵd���1��;[\��\��f�Y���Õ�QR":L��0d���;Kf�ݴ��T��Hsm�΀9+�eN�s�d��c����C��9� d�n֍v��Ӳ��lv��ZNMm��;�J�f�l`���z�a���6t�6�RV�sjH�W)�t�q�nI��ޖ:�U�ff���@u��q��deAӅJL��ny 6� �1 k��w�ӏ�RRP)�w3e�s���9����^j�1̓mB��Dm(���� �1�ny�~�����x��j$�ED��9��`w�5P�6h׻4�2X٥tC�R�"n�	����]xiƶ��Y��%nnK�u��d��*mJQ�rFQQ�J���f=��1 oI�y�@8�,�]�zɲffm�y���jH���jelܒL��l���:h��z�d�sL�n�� �i��$���� �se�޼�`�l��m��Q�q�E߯1 o9��@�b ޓ���#*4:�Jt���ri`z���i�����^l���2𝬓�sx��N1sZ�� .��[��G��:�1�R�r�q�*JC�`�l��1 oI��@o�s���)"6�NK �we������K1w�����Ǵ�Q**O����9���I=�>����SG�6f���wvX�z����TqR��$�;א@���& rb�ez�0��qXs6X;�,��,�&�\��F�#rH�Q�7%4 �(��m�lWn2�u�m��n'Q��𝯌9z�PI����N w=�`��`w�5X36XqV6�ӥ�nK�3vs��ꯪ�ic�Gi$�n�s�$w&��UM������ʍ�)���I%�}��]���$�ܚKI$����I!W�gL���[�d�ws��Ȫ�3�����߻����m���|��P���  �D
���s�ym��}ݙ�vJH����I%ܛ��\���$�ܚKI$����I-�6+�)H���ia^�k�ʀh�Ǜkd�x��v�����a���ࢤ�ғNH�I%�͜�I.��,I%�͜�I.�ح$�v���$`�J���I#��R����Iw7ӜI%�=��\���$�n��I�����%KI$����I%ܛ��\���$��۩i$��h�rA&ӓ�I9Ē]ɱZI%�͜�Iͺ��Is3g8�K5hڸ:PR8���V�Is���I#���m��~����~����A@�,Pߡ�eϴ�Ҕݶ�	���f�	r��G��h�Z,���:r�9-�"�Y�HX�՜�������==v2���q˳�S8�K����m�F�u�vm9�B�Eڵ�r� r�U��4M��X��v0X"�X�S]6p�x�'j�&����r�m�B�c�\;gX�y����)�؎���s�a�;\����}sHKw-�]�.��ff�ʂ�D�;�<}�VGD]
�f��-���3�p�el�E�[�#��)۫q6ȝR����tG&�$���i$�;�9Ē]ɱZI%�ݜ�I%Y�i�9J1�0�T��K36s�$��b��K��9Ē;�Ii$��̓c�����''8�K�6+I$����_�m���ZI%����I���%*i���\���$�ך���Y���I%ܛ����״��#��&)'8�G^j��K��wӽI%�=��\���$��єO�����Z�0k���uv���V'Q �uίC���qp��0�ܧCMJT�p��Igsg8�K2lV�Iswg8�Gwn����7i����ӓ�I9ĒY�b�����UG]���$��4��Iw3g8�]٣j��AH�*tۑZI%�ݜ�Iͺ��Iw3g8�K�4�7f��*:N���m�`�b �� 7�A k���ʿ8�r�#D�Xs6X�������,�͖���a�/' �NTi�p�^zY��K�{�N��MggpG�\$'`ݫ���lqTqM'' �l�`��`����Ws`�ࢤ�@Oט �b�����؀#��@w8��OӒS��
���wvXw{��>������\���F*j���%1#!$��B- VҊx�pH(��{V��*E��3D�`š+�H�+���.)� �
`e��F0\�� đ�.B	##3&9p���E"H�-)J�XT$!%!+�`%�HR1�0�Y
P��,�HF��D ��E6j)+"F��T-e%��`��X�@�Q}�x!������XsS�*�x ��X%�*|����\)p�����G�$����x)i��=)75)Sm�aʪ�,�zX�Թ7������^wM�o
��R�C����UUO��ޥ\̙�3;��$�ܼޚ ��I7�>e����^"b�[�0�:y����9�W-�p�u��9v��t�ug�{u��~�������I��z|��4s2w�ޥA罚�F�*:N�Q�M�`�����9��V�����ԑ�[��ێ���!��y����@kqR �s�1 r�6�*�"	��$�9��V�{��y���I��S@�8�!�~�����O�IH	��X;�,��k�w6X�J�g+���qT���u��.��RYɶtv�m=���vT��V?��7)�pT&'%�s���7��� �1Νd���X��������� 5�� o9�\�`f���\��ӓ��s6��9�b �& �1�˻��ר=�V~���5Ɉy�@syq�lnB���II,��,�͚3'J ��������3xL�Ao���Mm��%��i�eyvܖ�6���`����"����w>�2���2m�Z:֊��h��U�e�-���:;L&�����9R&��GI�g����Oi�!:	�'�����,��:6��g�fe퉛:�O/�܁����k��0�0[������Ƃ�ў5K͌��k��ʇqX,j�S���a�7m;��e��{��ܟXw�h,ڬz�M�r�[��
�,�V��.�LKl=�;tN��&�l��Br`��,̚X3vX7vXk���$UED�C���A k��1 ssSǴ�"��D�,��,��,��,̚X�x����TpT&<�@$���@6�\���YSe&���Ԓ�;����ɥ�s7e�s7e�����Su�H���C��⡹ny@�v5�nAË�ZV�ű�I�&7RA&ӓ��s6��9���9�����`w��n���7EO�L� �n�s$�C2fL�/{��3w���f�X�[��
��Q��=��@��G33$��7z� ^�M�Y�Sn6J��hNK �f�36��9���9���;]Ǵ�"��*&�/3�� ks�1 ks���~~l��y�s5��I�V�v��<;��*�8����aj(n�rg�u7.`�ڷc=w��5��d��5���T���Ǵ䌢�"��ܖ�ݖ�͖s6��9����VT�I�覤iTD�� e����ҌI$����0",FIdH�AI _T�������}�@37e��3F���m9>��`s2A ls�1 >s��X]d'"��"J ���ə�'�ޟ no���ɥ�ݧ��!N��7N uc��<C�@!�=�z��D������U�*B���dE6�fl��l�9��V�͖��z�q�Q)�&�$��b[���1 ks���*�"�h��,fmՀsse�s3e�gse�ew6�$ED�
&� �b �� �b��Uz��@oi��q�QJRL�K �f� ���� �1�Ό%]g��e��������#A�u�=�ٕ��J���I����4��!e*���tSQDSrI���X�۫ �se�s3e��n����I6���/1��Hy�@���� 7����8:�*)�*�9��`��`s�4�;��Vq��jB�����]�b �� 7�A��Hy�@j�ש� G��7%������fҠ^l��vh$ɄɘfI�n�?�m�N�yYy���8�x-A�h��Ć�������&v�di�rB;Q=������Ք9� aj�u�)؝��F�џ9��h���t��a�(�ǳ�v�ݴ&N���nm�����;J�F��q��-�4��\�u)��ή�b�e��L����n14nT^ۍn�S���BkYs��CC�[�]�P=��W�z�]��Dv��ş���{��gk������u�voS��V1�у�:��Ӷɧ�ڮzR�r�$UED�9%t����9��`��`s�4��̓mAQ+�뼤�� �by������[�R0�&'%�swe��qR� �1Νd��߰*���w��@o<�� �1 l�,�tn�:I������u`�b �& 7�T�4{�aX]�]3
M�{p���Q��ݝ"�vz9�6F��ƁBBH۩	t@�� �se�swe������ͺ�;��cRFl�]��y��y�Q�O�Z	Lb1LD
D$4W��W��gK{�u`�l�5Vk�ێ�Dq�n�rX�M,�۫?W���$ww��;�zX+���H�(���q� ۊ��1 l�}���"�@�}�"�B�r���,��,fmՁ��u`g��jj���0u��ܮ��A��c\b:z�E&����u�1֔ӃR2�p��crX3vX�۫��u`��`w+*l��`:R+�f 5��}^�$�R �>��L@wMѺ�8�&Ӓ�rU��ͺ�fl�~���l�6X�۫{������
�̤��@��� ;3n��[��
��(�*q�`�؀��7 nbz?W�W�WK��՘�uъҺ��Q���f�x�]f3� 3���m�K
ϛ�^^��~���Ϲ��H[��5Ɉk�ʻ3=X�*&��*��f�X36X3vX�۫ ���68��(��`̘�5Ɉn*@sqRu_�/ٖu�W�e�b �& 5����H5��� ڠ�t ^���r���T�I�()��K��u`sqR �� �b �N�]\��[M��+g�f�y�սq���<�U[;D 뙨����)lpn�t�i�#������5��d���|'ʐ��]�,3,�$ ��@�ٮI����h��Vs6���u�ڐ���$(�rb[���U~�_��'ʐI� ��ۏ� �hi'%��ͺ�;��V�͖�ݖ��=��EQ4/7 nb �& 5��+����i��h����&B�L\ԅ�����%S�!a�p#9�i31�������J@��"����2bA��V%HՂ�4���!@ F@��%0��"HBB&�8Ӌ ��HgaHUS%�U�BHq��c���\"f$Q���`FI��`���XX���`ŜU�s��!p�01�E��1��$0��)XFfBJū!-[3�Bn��K�*�q5"��40!FI�R��Z�� �	
hF�$Y$�Fuq T(bFk�	V A���!\`č�Sذ��ͦ��I�K�	�[#6���$E��F4��\ I��P�+�\"�"A�<`�HA�B�Q�b�"'X��*E$!DX���Hzj@�b����B.k
K�"K
ܙ���c�"ԉ	B3a�c��sn7c�v��꿒�U��=�ngHl�5��y�o]<�7��ݸ-sːɤ�X��l�m�n�4���ht���s��Ѭ�^4q�\k3�^�Fƭ�:ۗ�zS=Uv����nv���Ť�$͹�uc�;1��)ٮy:&l�\�l��lZ�*�����1%��۹����N�Eu:v̋Φ[�;l�βh8;V�nέ6��Wo>�!��v���[�����c�v4��!��l�b׏��}׻g=cF�c�۔�Q���*.�3AQ6�k0
]�ݺ�WM�h�$36���l��+*�d1����a	��6v`*�tg���$и��dN�p[rWl. ��w�֟�&���0����x�k ���)��T��g�Ҷ�]q�iY��e�'l^����UqGnqvuk J�]�B�g\� 'g�	�ͳ��;gm� (\�Ùq�6�]�]��e�q�,9���÷���Q�TD�i ��STK�];W:��O/l ���gg765�8��h욌���Pm���r��A��aVpWe�j�l�km�3�p��0Z��B�˵7;Τ샪3ԡ�[pjx��P��[R#9*���ڶ����e\�V��u�Ԣ7a�mG6鶶Kn�0 hq��^��յZZ��W�_ �N��o^���[mۥ{�n�b���
���ݚ��:9�٪�W��qu�=q��^2q��}�{z�Zj6�s�A;u��1�;jA�vg{�kg8*\���̬�IO[S��B�mThS��RJ��ۮ�K���ų��Cmح�H�:�%�Mi����`G�US����;��Ö�,Qn�՚%ڢh�2��3��C&�9g8�U�
%���m���fT[���4I�r�=���l;�8�;��2�\�c���Sye���[�&��Y��\A)�D9's�h���!��=��1�˺�j��4��8\�OYSU��n�KtR����$�Tsv���l.vR��p�R�B���.���&f�L?!�<��@�
�(?)⠞"8���x�����嬙����YeJ�g4v�]���������q�y=��3���E�'kWm=u)�B�;��n�֝��'^	d��-&�t ֱ÷]�sh���
q�t9�:B`�ه\�H�l�#�����޳�Į�'G������Vڸ.ݐ^��l�8�rF��ݱ��z���1�p�ޤp#d�[�Oa��T���p/]��+=]�/>�X�M�e�eM,"k���N]���z���\f�ҽ\i��NH6H�"%@DnW�37��5Ɉo ����H_�,�N�DL��vk�3�{����J�9����VT�I��pq���X̐@6���@$�А����I6��9*��ͺ�fl�n�9�4�9����H�"�������1������������%%�,�8�&ŷ<ۗF�ʖM��:�b��[Rs)[�C�'b������1��n*@�bz��.�/�n˷�����~�j�q�`�aa �D��`�� "@�Z��e�}�xrI<�6X7v_�� �n�Sd�
2$�,̤��Hy�@$��Vf���"Tr��͖�ݖ�6�$�L�w{ʀ�Q��3 ��Q�=y�d���qR� ��`mv��T��T�������:�.6��q���gIS��X���ʸڎ9��m�0'���ד���J�=y�ə3. ;�zX���1�q�M�$������� �by�߿U~�����6��# L��nJ���X7vY��U}U\�ɥ��ͺ�3n��#m�D��y���d����h͞(��VIw5�5V-ѷ�D�t�$�7��w5HzL@$�w�A3 �\B[���.T�v��mE�ح&wO"5^N0W'39(��M�����6I��@M�.��"Tr��͖�ݖ;�K36����׬��S�*I���by�H�T�7��:u�*��E88�MI,w6���ͺ�w6Xg�*�����wf� �թ1�q�M��3/2��� �s�1�⯶߿�?��Kj�{[n�C=-��ۥ�#�)�B\gmun�t��Ky�!W�S��g���� o9�d���qR�X��[RiS�T)%�swe��I2w/7�P�Ԩٛ4���Q/�"Q��I�`s3n��۫ �f� ��� �w��
�"&���?�I�� �>��LA����� �O���ATr���,�_U~��g�}6w}J��ͥ@ZT�I��fkPJ�K����L�#�nd�%ٛ�M�n��vݠ�\Ĵ^�i��;�ϛ�\6$Ƴ:y��u!����6lH �;�өxl�@2�$k���i����TMu��\��j΂|�s�\۶����sX4�[v����m�-z2	ڻ�]�G|]�u�{d-׶K�[e�5���W�N�9���������ZT#���j X�9��HYM��͖�f�����@P�w���~�9��Z3-�`ӱsjx�h�&���!�\d`�)��9���v�nqJD�&������X�۫36��_W���3kjzP�@�I�%�����x�|� t�b �& ��ɎT���$rIVfmՀs3e�swe��ͺ�9����H�"��p�nb �& 5�� �� ��ڐ��J��9,��,fmՁ��u`��`n��n%rD���a�R�^�0.�L4��S6��H�F���5tW5�D�ct����f�X��V�͖�ݖ��=c��*6����T����UW�-���������_U$[��mA	PMʰ���1��H�T��W.z���)B*I�`��`s��VfmՇ�$�w�ޚ5j��D4��xy��7�T�m�Hy�@$��2�hi��=�8��uP�)1C�'n�-0Pa�\�ҳ�h��YH�Oc����� �1 l��*@l����# L��nJ�w6X76X�mՁ�ͺ�3f�� �I�5B�X�1��~�^���Hy�@OV,�h�9Q��'%����X��V���R]��,�����6��̤n*@�b �& 7�T�?}��������SIH�w=:��X�3��d\��ι��&� ���ʖ6��؆��6I�� qRu=z�q�R�*I��n�9�۫36��9��`w+*l����5M�1��n*@���L@'�&9R0i�}Kw}ʰ��X�vh5�ٙ&kI�'}�x�/wb!T$`	�QM�V�͖�ݖ3&�fm*��g4�:��O11��f�y��8ʼ��<��0�t]�J'm\��k�m�A���7Drp�����ͺ�32i`��`j�Y��P���I9�o �m�H[��6I�k��8�p��:t�����K �f�=�2L���t��<P�͒ �J�%`^z���@$���@6����N8�)T�	��n�9���̝(ٛ4��*fk��u��;7��Qn"ΣihS�%ѫE�(��y,���4�e4&��s�v�OX��ݪ-��烞�RZ����v�h���0��`�;��5���&��t�L�՝���ܥm��au� &�tq�]��3����,\@������.ٳg�v�.y���k����j�6s�0e�m5J����1ҏ�.�T�N']��>�w|CCi�!r�������zd݄��q���}�y�!�ꭹ��y�z������g0v0݁g)ӧ%4�8�e6���޺�32i`��`��`�Z��	�/�y��m��1 l��T���˄����m��9���9����d���ɥ���ԄI8+�33�1�����߿U{ݻ�`yV��4T$��m�NK��K��@���L@}��U{�}���棆�uڰ9����X1`Հ��9k���s�k9��[���9�tF�犻����>�1 l��A u70�!R��8���s3e�UtA�ۖ3&�fM,�=z�q�R�
I�@$��� y�� 9ө��pFFSjI`s�4�32i`�l�n��Z��	�4ۂ��@�b �& 7�A mc���f��z� �X\�c��i�,�[��[n�a�vz���6�z;r��5��d���⯫|L�@OC�mI6&�J�X7vX�mՁ��u`��`j�݉��$n���ٛJ��ͥC��I�C)gv�b��Yh�`���&!
����~�L�4��Ë�
�`�Y!��[A5�5cX�B$"0�e�I+���!b&$Z�"�,��NbB	 B
BI	zJ2���Ґ!)
�$� I"��LE#��C �!��)$�����P�Q��`�X�!!�
�Bg�&7P�#�tLC��P;�:1Up�4T| N�_A�U�tE���x"���3�}��N��w�Wq��B@M:T��`ff�X:� �by�H���مf��g���6I�� qR6�{���}�-��q�.��]q���ӌ�۱s�fm]�2��Z[ץ�z�G1pӧ^'O_�y�d���qR� �1�ʛ!�22�RK�ͺ�33n��͖�ݖ��Rc�#1�x��@ffҠ�٣�&L�_wMy�]X���]G�*Tܕ`�l��bzEH
�U��� ����"���I@rK ����ݺ�33n��͖�Ċ�r0Rq�I*8�1��u��ѧ�5�U/:�ڍ:W��Q��]4,�IFۤ��;�u`ff�Xs6X7vX+���R	M6�'%X�� ss�1�EH���eBT(�Dܫ �se�swe����X��V�=z�q�B�
I�a�$�}�4�u*36� ]��y�6B9 "�)��%����X��r���4�ݚR��d2&��F�  ��T���}EWո
�e�P�#�QAK#�ь뗩N�pDwgk���)��*�����{f�/O��`�b�b"3e�L;-�n���ۍ�;F�L^w3Y�nە�ja۷�4�襘�i������)�[n�h����o�&�g.j��<V�$�v�kPJ� ሶ��sڪ�v��\�����V��+�ݬ�۶�WW8ӹY���@�rKn?�d9s�f�S,߅p)��~�h�Z:�d]սq��ݧ�K�Ol*�;Qb���7���|�n�l9���0|��� w9�d��ޑRt�����*CpT�� �se�swe����X�4�1t�r9%6�q$��,d��ޑR��@�bz����T�m�I�`s��VfM,�͖�ݖ��zƩE)��I�Vo �;���L@oH�?7����]=S�qr�,"k���ϝ۬/��=���S	i,�)oa6���rJ��I�1 l��*@6����^n�	M�[���$�����?�h@�	�C�3&�7�J���Ҁ.�f���1�G RSRK�ݺ�32i`��`��`�tL����8ӒU�����X ��7x���@|�����u(����`��`��`s7n�̚XU�Ѓ��*6���ű����0���99�cFw#x�f���w������rJtӍ
�p�����ݺ�;�4��}�f�X�}�>n��^�� 7�T�����@����ߪ������G*&Ҥ�7g�	=���'P��`#V*DX�� @�)��5�d�����7z� Z��"���a�/0@�b �& 7�T�ꯪ�nߋ�Oމ�*������L@}U��s��ɟ��@?�_�G��Vκ�`�k7m�t�u�zu��:��.-Z^��jZ&�n��r���ݥ@^d�@y���2k�3��hߏ߄�	Ӎ9%X�4�W��;�f���t���T���*S2��(P�"J �͚ ���̙;�wUX�<X�n���4�I@rK̓%�3%�}���}J��ͥA�����"$��������I�;�v�K�̃�DBw��׻J��L�����f�X7vX܍���MB�dy��ȗ��ݓ9M�F��g�H=���]��{�����eINRM�I�\w}u`�1 l��*@M�.�٘~2�^"U ]��s$ɝ���h��T�m������=��蜑�B�&ے�:}� 7�T����� ::˙鉑
^T�"fh9�3'���7w�P�l�s33$�}�4�w�3 7N4�`ff�X�噾� ��`s��V�q��'�)�IT:@�����O3�ft��I$d�e�5IIz���[�-p�"!pW�P�l��6�nՀz_]c��e�(�p% �2:XƝsG�Л�:������q���Ga�p�D��Z7m;3����ͷ6#m�v��g� ];�ۻ�p{v��� �g���^U��8Ac&��.qX�d�v^D]��7n���^�M��w��&Z�;;7J�,��Q�yHr���1�:/2����ݻm��~=����˷}ï@�����������L@oH� ۊ��j����%�,��/�_}�_&I��3~����R��ٮI�I����n?���m�NK��]X��V��� ��� �f=cn�*A(ӧ��AɒI>��� foM {wf��3$���T�w��fF%@�$D� �s�1�"�n*@Wҥߢ��a��li+�̄;�/c�u�;d`��P��i����wv����j{v:��6�}����TfN��/8��`f�G褄
j)HmI,wv���2kd�Ғmfk���ϊ �͚ �������|{�d�R��q�$�wg� �s�1�"�:O]�VfW��A:m���T�n�X}�K��ua�[�~,XyzE$�Cq!@nK �& ?���I��L@Il�����P��Wd"�g����V-���Ȧ�J�3��/�����]��H�j�.^�[��n*@�b �& ��XܟJ�J4�9*��ͺ�|�f{��;�zX��Հv�6�IP�2��r�I=���I'��w�E`)�"&&mX̦f'iP������30�H	6�K��K3޺�3��V�����������)��!��;�T�|��& �bJy3��M��uƸ��=:),<'ur<�5�.26���'Tyk��ëE�/25w�8� wI�c���R �Oz�RJT*N'%X{�/ߛ������������X�j���������R��H�L@OSr4��H
6�(�����Vf���=���I�h!SA��*z��VM�%�v���>��(Ҥ���J���3'�� ^wMw�J�<���Z�zY
i)N�=:��X��v�&m��s��Sm��se�z欻���;��r �����W���*@}*��NE H	F��������Ձ�����v_着�3v��RB5#����3;�Py���&w3;��/=�`f��e�)@�8�7%X~���foyP�t��vh>fL���T����GQ�I�V��� �we���xrI�w�$�."�z)"�á�:��ߑp�>�'� 0#D#� ���X�Q��B F!8���Ā����1���T~�"xD(v	R(Z�Ґ���G�g�0
�����U�b��,`�$F+�C����� ��( @I!� E,X�! ŅH"X�"����-+P�`d�#B�F���!I�%`"1$�YL��L��T �JHI!� ��2�� JQ�!$�a�y¦H�� �HB�0����6�d!$�%$aHBHbBC� �Z,0P��>}Xg��}������-�[�n�J�u�:Q�I�!����3���.�Kͱ8�U�Htq�{S��TN�mOl�5v)�ȓF
���Ld�[L��lc�vz����aL���B�	�#���4��Π���q� ���ѣ]�H��\cte�d��Y͛�ts���՝=O乫e�6��<��C�+�����g�k5�9�k;�Ss����H�M��{�]�A���sl*�񵝹�K�.qr�ɶ�<���#�찣Ɖ�et�V��I��"�����8�(Lp����B���Q��I�7tqi
��p�+�6t��L�ȝ���d�ճй6�u��t�cWRjb���\q�%����*�IJ�ut���uq��7=h)��x����r��m�]W�\c�X5M)p@�*k籮������N����]�u=e'LP�m��]r.z�5�M��'=�r�5���g������OmsiX���<��x�:x;i�y��i
�f�n�,�8<��5�rn@�-��\ݷ���@3�p�� .��	��� jwm$l��m��燶�E�&��Ó���k%���Y�F2�]I\����nc���v�!V�$M���7nu۬�I%� �uPA����q0bh㸼!��K����r�Um,:{��v��i�V�eH֯Z(ݓ��ć2d� l:�C�l*�:x��bxU2��k<us۱��܈O�����eL�.[�\b��)�{kŷ\m���@>ƛ�:t�������^ɛl���Pvp���!���=��R�W���n۬Ke+d:�!�76�&JZ�n��vev�{ض�x!��"��Γ`M,�nե�$x��Wfű���6lgn4\�n�������nw0�=�x�+���j�̸��E�.JaF�oV��Ԯ�#�S��(�M=�s�p9�Gd;;���0��<l����`��l���)V��]2�N�4�i.��ܛa�f\ͷ3JL�$&���"�$DC�#����N(
"�QC��"	�!�x��)��gw7bx�Kv1]�l�����4��� ;f�!&�
��MD0���Z�:6�f���.���N	o�L�g��IO"�ɹ)�h��`n҂�ۯqs� I�8ۤ�>�&�ck��J������Uo[��(lA��n�u�7M�P=,��ٵB�'cm�N�5A�On=��'`��5�3���K��mn�c�v��u�?]������P��Y�f��E��Dj�n�܎!㚨밓+��wB�������QR�2�L""g@/7���ͥ@]��ﾪ����{�����5P���J9�� ;�T�7���&/�~���� ��~cr}(Q�JIVs}u`였7��s���9���2��,�u1�9�I���t����y��;磌���r�e??'�@�@J7$��1��������_�U~��}k��
#�.���ۍ9�Ѻe^@㫱��nMR��Ӗ�-T�����Q&R4����=��˫�ͺ�wvX;�,�4L�E(�&��ͺ�L��3+X��3{�3�4��4�m* ����J����8$� �we�r�f�I'|��T��*v46!�eB/�.����� ;�T��qR�~�����5V��6T$���ҎK�ȩ�W9�րs��@�b ��{ұ�Mfj�9ж�^�ڹ	#pu�ݺ`�[e��Ƹƕ��+���"צ6$8���~�n*@�b �s?ª�~���ʐS��5�� ���7*�9��`�l�;�۫�ͺ�ԑ�����8$�9����.�iP�3z�!(34$�%�2PɓQ9�J�=��@^☍y��f�DD����7ѻ�Z�3{�T��� �se��f��	)�t����@o8� oI�y�@w8� :?�;�[T@�f�烴���&����m
v�]���G,Ly�x�.�iާ[�@�b �s�*�|�ʐ}�Q���(���w6X�mՁ���X;�/��$j���l���t�)���z��ͥG37�o}4��M r�64ܟG(ҥ$��ͺ�{�w�I�wy&���C=J�<�^Հz��F���MTnU�o9�y�@o8����W��U??���%rh�p;�Wgl̢n�S��w/�YB�b�KX���'lsv�Z�a3�àe��9� 7�T��qR �seީ@��rX�m��ꪯ��͙��u`��,�͖i�&]I)t��י���qR �s���ޑR d��*J��'%X{�,��4�v�'���;�j臘�et^f �1�"�s��s��'���;{p���!M7L˷r7zxY�Q�+k�d8�Ԏ��4��*v�7{Jw��wi�OsnR���ٶ�]6ôŉ/:�����aMp�8�2�n
�v���<g^-�hpv;m��Q��լc��] ��H7g��2�-�d���ܵ�����Q�V��<.�ε�"��c��g@�P)�-g���k�;S�ط$�]����5�$;����D7\�;���k�c,��J�x�F���-/��!	�nf���]M˺��^&�{g'ʐ�*@�gվ��b ��>ƜGF�'%X��/�UU}If�Pgt���U�$��za�Ԓ�	��B�37��;��f��]͕ �vi`b�i��& �n������`w=��٥�w����eF�H�*��<C���ݥ@s&K3�� foM w���+�����!#�#���ĐȺ5�zド�R�Q^�e��/2�_��:��x�O2�gOw�4{�?�ə/�L��3~�� w����.��ă�I@y�Vɓy&Q�4�m*/gJ����${�Cͩ%:%����D��A w9�	��r�ʼ�ʙxQ	�fh9�&Oy��@nt�@y��;��`���ӏ�"���gJ�32|���gt�{��_��?���7(Zˊ�R7Ck�	���g�.�x��Gi�Y�Ugm�����m�i�$���.�f�.�f��ݥ̙&�gO���c(�Ȑ�I`����gu*3�� �ݚ�L�I�h�;���E%bcm�`n��u`w�4��4j��r{���I<���I>[�D�e8<0�&ePs$̟3�� �� �ݚ��;��8�	S��<H<Ĕy�4�&L����/{��wf�Uwt*9$d�D��j9�]`役z9���fu�s;��Z_e�[����+JPt���;��`s7n��f���������<�7�l��"t�)4�v�|��2w/:x�������E?�\����ܹ�d��.��� ��� sss���"�����HPF4��,=��UIf鹿foM�ݥA�d�{�y�%S�|Pj;��"��H�3@{�@|�$�}�W ���`��`g�O(c{"�8�'L#���b7U�у��uΜ�n�5�.��X�T�Sn)��&6�sv���vt����e�3�h]�D�e8Ӣ:NIV{�K ��� �we��w�9���ʋ�'����\�ne�3I�x 	��� �1 �EH�@OWwRnIN�%(:JIa����K=���u*/gJ��3;�oM��zH��sLˆawwy$����$��G�������@{�@|�$ڙ�&C1UU�+H^���p���aD(�nڞ�']:��Np�u�g��1Qa��C�H��n�q�Rz#�`ll6ᩦ��ڻvD�c����b^�^K��λF�whKwPeݳET�i��۝��q �m&�Z��nr�uK�S�e�1�qڝ�B�k2���vݡ�n-�n�۲;Mkp]�Ļ؃�&�0d���"��ڴ8��,��hR���_����w����Þ_Ծ-u��-��������{%��E��2Y�����:R�J�F�t�(Ҥ���Łoy�@���&I���ԨVlt�3 )�ɉ����د�����3�h��T�Ε�2fgs�F���
]�~�^Z o���H�@o�����F�H�9�ܒ��n�X�Δ�f�&I'|��1wqR��v:#�ܕ`w�4�8�5�{�,fmՁ���J7#%9*'Q�P$�93[���_iq�n��E��Հ�rCFJ����a�GD��� ����l�9��_����s�Ł�[�$ܒ�DFҒ;�O{�w�*�Ą �&ft��2_2O&w]*�g�ϙ����H�Y��g�8�:n��X����gJ>fN�����4 ��6a�B��iRrU��٥�ՙ��;��A�&I�I�g}�� �A��ɂ=�/0@w�����?�٠t��H�!��������2�6����v.h�����qh%ct.��9+�Ƚ�������ﯬ���/�q�=��3v���f�X]�v�ToTR�r�brI`s��U�ɒ�7��T�w�@�٠-n�R��x!	�&Uw�J���lQ���5T:$���8��,ȨQ"`�R$�ȡ����C��^�E�E����b��a��)�2ni�*��ra���A��E B�EF�B$H�B!"��F0(`�b1E��SU^�  �`�D�� ���pP1tQ?*���
�3�y�MO��Pf�d̼3S@^�Ҡi��	S��I���T�I/�Q���Po�M�ͺ�;�۫ 雱�$�Cq(�RG`�٠>fd�|�gw֬������������Pv�q��A�)�a��<t�ς4**��d5�ͽz6�]�]{U�{31��H� 7���������
�f�4�)Ȅ�j����6�����`��9��W�H2�_���)EF4�NU�ջ�`�l�9��V;�u`oi����u��q�z�.����Ԩ��T��$[2�ə�ɒP��3Yw{י�ALD�Q��@k�R��H�r������U�W��~��Dr�b�2"�$�q�W\ڶ�T;p��x�ֳ��7$VS�q�uw�ۖ˾�1�'$�����VVf� �we��ݺ�i�&J��$ȥ'%XY�^wM{�J��ͥ@3cb^fTP�H4���9��`s7n��%����1n����`�T�&��t����}�̞��ʀ�ޥ@[�lP|�y�4 �n�4�)Ȅ�j����6�����_V=ޏ ^wM�ݥ@s2L�N���3&��c$uݓ�������kV�r���²�nmZVE����G�댠f�F��`��]uNFG���tVm��+S�#�5Ӳ1��Xŋ�{���n���[��;F����rX�l`��ֻ�f��m;/*����r��c|��nx�ݥ�Sq�:�k<,ۗEOY�n�ư]����.� �:�4r��ی������{��q�$kt��2�T��2�V�v����݌���tr2�r�)��o����2��F4�����}��;�,wv���sn��y�l�@�A ��hy�@oH���{���U�Uvo�To򑒂7)1�$�3~��9�۫?RX�|����V�ke�p��D���e ���9���}���1�EV�7D�Q��Ԁ��3]��=�����T�6��hs_f^!ӑ72���lu�qPg9w�LӇ����:&�pq�����H��͖r*@o8��rZ����Y��~0�]��I=����Q_R()���JL���"���T{�4�ݚ W]Ǭj��(�NJ�;�۫ �n�933�y�4ou* �y:�y�Q*��U ^n� z�f��ݥAɓ3�o�V������$RK �wf���6ow���ޥ@��@Z�i}V�����}/'?&kc���x�l�����6���&L��`9lr�N�m]q������J��ͥ@���d��p/;���ޯ'WMi�rJ�;�۫ �n� ���y�J�32N�|w��H�D�L� �� ����$��&M�v���ݺ��\RJ`�I6�rPrL̝�;����@]�Ҡ�3$��o�,5j�%T�6��t����f�X�*@���& ���W�u�s˵\�q{3�[%����iҎ27�n4c[��v+7,?�Vs�̙v�an�f�I>s�H\��7��7 �w,��/0:�hu1�ٻ5�&fw��3w�Py���d�;��7���R;��34y�4�m*>dɒw�ޥ@�zXܨީ@T�6�s6�w�J�=��A�Й��䛱33(��2�I��:nh��s"H!�2���Tɓ3=�t��h��V�v�F8�rr��T��C�Z� b�J�+l�d�iܬN���z�a�Oh��q*�=��@�٠/3i|�L��ff���u`{���SN�&��^�������T�͚�nd��yy�6ҡRm�;����P�ܖ��e�W+1�9�ڧ$����� �1���{��i 7/�4ȣ9�U�`�l�wvX�m*�6�,�$$�#5�lDA3*"j�R�Z7�����Y!y{g��q	��;d�����C�xw(�gV�;��Mf��l=�6t�1��1�"�X�;]�,����;=v�󷱧;��1���q����hcs�����2qN���m��^���������Yz�h���[���8��Y6sśe)�� QD���XxW(��͠��z{c�y�{�L6�x��||�˵�l.�Vѳ2����`��>�aOC�%�r���$�l�^8������כּ��{x0���>��*@w8� o=���=R2|T�)PےX�mՁw�J�=y�@�ٮL��V��
`�0����L�3z� z�f��I�'r�ޖs}u`�tL�D�9��aə����h7呂�fҠ.�iPU���$�4�)4I%�s����f�X�mՀs3e��h�����*:�����.�J�h�R물͖����Q��'Lu�,�U�V��I#T�:RI�;���ͺ�w6X;�,�����P������9$�߻ÕE""��3����t���Tj�6��<�D�z��) o9�zLG�{��ʐϕ �f�2�Sp���a����Sy��� ��ʐ�*@�bu_�//,D�yP34�6���n�֬7����� ��V:)��GiBH(���F���8�v:Nj]n(�v�"-e��p�~����Q��������w6X;�,w6��9��*0�*r!9*�7�����{����|���z��q�4�J$��9��`s2ic�W�B0 ��C�Oʨ��y�� �~���3B}"�EN��$�:�� �1 o9�i��z�Zf\O0�bJכJ��&e�(���3}�X̚XY�ll��R�#p�����.�\��V��'�V�(�Z���*9�1�
R�s�ܫ �se�s����ri� �o���[�l(��	.���y�󘿿W��$nS[��D��:rK��Ł���Y��;��`����i���J'wF_����1 o9�'��N��fI t�&����(��	R�$�H$� �f� �se��ɥ����XUݭ�9$� �*Aӌ�p�]c�^l�M8N2��NgR�γp���h���X&�NQ$������K�ͺ�q��K �#|�I#L�X�@o8� o9�y�_W�x:���NO��Q6������w6X;�,w&���=cn��)A9V$���zh�zh^N�&Oy��@��8�aE9>H ܖ����ͥ@z�iP�6hJ� d�L��2,D� 1q`=<�`� H��Y�$�b��
w��{O��� # B5pH�Y��T�b�^���bMU��V\H�Fe�5�0\!q%��0�Wn�o���$)��2��Ħ$�������5�t! � �Z�hȫ�b��dHA��c@ H0!k����0�b`�0��VMF"��H� �]U����A � E���)��+�J���|�n�x杸�
����ɹ-�^�
{*3�\[l��z֭݉��2����m� e�nM�e����ϵ6�vy4b]��! ��w;!�gv�=0�vi���6�;��1�Z�C�� 园B�lD�s�]]�ɖ���=f�E^{j�Ld�C�6C<0M�ꆀΖ�� ��\�lj�Dgd��7i#Q�q���gs��dM�9y����.=�g�{<T���ʵ��n��m;��m[vsۍ+ӏn�4�M�@1�A[AL��V�\�ƶ���7m��۠�ݪYYTj��ץM�M��D��X`U�cis]��.���n��m���ܥc���B�m\qɆwnG�C���p�C
��]�"�[�n���h&���[�*�	�ۖhv{In.�jd^3Mʵ��caX��V� �"ZYٴ^�����8��BcUͤ�;l�b7(35���K��ONQM�I����ީ�s�rĉ��l� �Xx8n+q��ڀ����%��Mv�Y�G�;\
�Kq�4*�>T>4�'��*[��
�9ǎGq��1��μ�I��'M���p�ݡ�<LF3�ؙ��h�e�F.I҆�����Irʷ15�I5�f kV����͂ivͷ�ΝT2�j��q5m,uJ�-�iݞ���U����8*��auYv�r@���]�*zcۦ�{!vT��hn{o)��VSm�5�u�9nE�;t���u���1;�e{]�ݘ*�K՝tH�%@.϶n�#a�ݴv�v�t��ay絁V�\�v���m���*������6 ��N�;3���^@���ɰ���uh�IoW[@#]쭞��-��M����YN�P�q���M]�b�l��d�;9�]�t�3=��Sgd����9w:�={Y�B����L�2���`�װs��'k�Wn-�@#�g)����jF�!�)(�x4����F�e:��۲�c��inxH���K��3� �G���!��� �x)��0E��¡��t�T�����nf�f��4�M�4����s]u��/1˗)��������ڸ�\�ĠZP��t��g���u�a�m>�v���n:�Sڹ�����Umk���^�K�7v������:s�#�5��/cS�G���WQY�B�nX^ٌ���ӈ��с��.L5q<1L����K��)d��=f�u�z���!��k��5��\���n�NY�&rN&�wws��x��$�"κ�Lv��Vsm�l��t���q�r�n3̷N�;Rfi�����&g@�ͥ@z�iP�6~L�L� ���`�~?'�(�anJ�9�۫ ��� z�f���Үd��/���J�"J��NJ���X;�,w6���sn���z�ni�t�Ia��fL�y�4��*כJ��L�����y��I"`ؤ���sn�w6��9��`�l��&ж(�)�r�ѫ%�J�벩��aٵ�9���͹8��}�UU�KwM5
�!Fۥ$���]X�7����s�*@������2C4�v\ӒI�wy����z��d��7���ͥ_$�'p�[�/E]�^�aw��9ϱ���;�,�5�8�(����jI`s���^m* ���3$�;�oM j�<�(��rU����X;�,��4�6��3$�po.�R�DJy&yzr�Q5�-���^\�#��b.7���9�	g��W�W��iT@DBA�%t7ߥ�o9�� 7�T��Sw/2��z��_���@�by�H� �l�UUW�$�o�T ㍃t����ޥ@z�iP�%�L���d�)�2�l�͖��{M5
�"6ӥ$�כJ�=y�@�٠���I$�7��@[�����aJS�`�l�w6X�mՁ���X��&�1��)*)qX5�5/S��g��[�I���su��t�{=l�{�}UU�W�QNO�7' ;���7�T��qR �s���y~��e{*���f 7�T��qR �s��~�� �������lAnJ�37�T�͚>I&N��t��Ԩ�n��T@DB@nJ�wvX;�,�6��P�dړ$�T�ϕo�F��D�i�&�nK �we����X�mՀs���ͧ��8��7"Q�
�T��\�u��ʷ�j��MZ��·W�iF5v��e粋��fby�H� �1 s���;Y�i��D(�t�`w��U��&d���h�h��U�2gp��~cL�R��Q9V��K �we�K����37�V��[�NO�	"&h9&L���h��T�m*����.��X�k|8� p���$�7�T���7>��s�@�b�P��ga�gM��\���fnc��]�雱�ۆ�+m����V���ۗj���NM�/T��HgN;6�=7���+l��S7Q��[L\�S��79
�96^-��?Ӿ����-�9�u���̒�k�WH���cK�vحĻ�SuA���i�n�ݵ��:�ۃ]�uS�rN���j3�pRro�^3��KN�.�M�2���������I��M����R`\�d;1�ݐC'j�[�s�	v���qͭ���K��Z���s�Hy�@�by�Ha'�9Q	�*�9���9����f�X�۫�{$n�M4F�)$��b[���T�5���zJ%H�%&�9%��ͺ�3��V�͖�͖��lq�$Dm�J8X�T���I�h}>���@�Ia֝x(Ɩ�3ι�zc����-c���u�u͸^a�WK�p���g+�x��:��o9�c���y� 	��2fa$3�ɲ��$����抿��A%ə2��;����@�٠6�djq�A�����d�����X36X76Xkv�84���#m�X�T�5��[����`�9Q	��`��`��`s2i`s3n���ݩ�&Ԕ�h�i�:�B�Q���A'`q�MiH����74�)4I%�s3e��ɥ��ͺ�fl�ůiJ�j8�4�rK[�/��W�t�*@�� nb ��lq�$Q�IҎ36��9�6\� MB�����K��`o�4����4�q���7*�7�1 ks�A��Hu?ltP�) cd��͖3&�36��9�6X��AhR��*?[�}�s�i��S�93�8�ݎ��og��g���.��عn'�J�:n98wg���u`�,��,��Z�u���n*R����nb�ٟߪ�y4�Hr�"9*�;�zX36X̚X�۫��o\6C�$���~"3��3�~(fm*ŀ3�~�3{<�I'�^�K��˹7L�&n�$��{�~�|�������>A��������� � � � �{���� � � � �v���74���๓^�ѪR'#Q�a�1��W��;N#dnܔ�8s�ٗ7ݻ���w6pA�666>���8 ���o �`�`�`�}�o �`�`�`������� � � � ޟw?d˓6�5˳3N>A�����g����lllo������lll}�y�pA�666>���8 � [�����$�a��نn�A�6667����A�666>��~�|�������>A��������� � � � ���ٗn�m�rI����� � � � ��y�pA�666>���8 ���o �`�`"X �{���� � � � ޟ��lˆ�Ʉܹ����A�A�A�A������ � � � �~;�x ��{�x �~�?N>A�������g�j�nu��)������U�j�ɍq�XC8��\���]�u�"{S�{68�E ]7@��n_EjᖇJtB�pIX�oE����G^li�C�zy���;�?&��:9��h�'F�u���D�y�Ke۟�Kn��\�@��-�7���s��l�a�m�mvت�h^�r�m[��u����ۑ�u���#�l��s���7n��m�n�a�����p��p�ۻ�ef5u��eU����ckтL<�rV�V��l���)�m�m�7f\�=|�����������lllo������lll}���8��A�A�A�A������ � � � ��;��v�fd�\�����lllo������lll}���8 �{��|���������� � � � �����&k��M�3	���� � � � �������lll}�xpA�6 ��� � �o�?o �`�`�`�~���x ����ٗ7ݷn����� � � � �������lllo���|��������|�����w�� �`�`�`�z}���.L��K�]��pA�6667ߎ��>A���肦}����A�666?w�?� �`�`�`��{�Â�A�A�A��w�=������8.�\�F���Mv�;�緧6�X4u������y���]���/X�a��|��������|�����w�� �`�`�`��{�Â�A�A�A�A��w��A�666=��3�f��n�d����|�����w��"<�P����q�*���b"_T~����l~���>A����������lllo�������e����\ٗ4Q"a�"J;��@��4rd�$�ww���l�`�4T�D%	�����������@'؀��n*�:�X�4��F4����͖��@kqR �d��������\���c;i*���y0W����S{4�-&��㎐Q����]��>�n:lt9' ������� ksW9�����(�7J8X�۫ �sT�fl�;�4�}��_RA��|ę"t�>j��y�=��Bes,�Ǉfbd�#� "�G�@�04+s � �A.�	l:�\��LR��d(�K���YYr\�e��I&�y1Kew�J0����,#m�RP�����c�1L!V"�![�FA�L�e�U8"z�A��H#�0�B�>��A}C@j �U�W������uQ��-I+fI$ٹq�(��T����(�*U��͖s&��6�32L��7�hů�S Kʘ(���@sy� �=�c�`~���V�RУ�F�dEI"��uu��ܶ8�5�C�jg��D[����S�����F)��&�:�߮���R�9���UU��qn���S�D�9���=y�4�͚�'Ij8��N2�߻���%�bX�ge�n��f�s-���jr%�bX�����yı,��ND���,2&D������%�bX���۵9ı,O��~�[�˙vfL&n�Ȗ%��� ���59ı,N���O"X�%�}��v�"X���3�9���x�D�,K���̹���ܸ\.�bX�'���'�,K��@B9�M؞D�,K������Kİ~��59ı,N�N�vfM+sM˹�˛nd�@)z+�s�����\v��U�-gn�)9�����L�)��q<�bX�%���ڜ�bX�%�wx�D�,K��S�,K��߻���%�bX�z}{�3$�f)M��v�"X�%�|���'��_�E
�M�`����S�,K�����O"X�%�}��v�"X�%��O�o��a7rn����yı,���ND�,K�~�Ȗ?�,2&D�w�ݩȖ%�b_w��<�bX�'�zfg.\�fL&�s3f�"X�( �Ȟ���8�D�,K���v�"X�%�|���Ȗ%�`���jr%�bX��ϻ.M7$�i����8�D�,K���؜�bX��s����=�bX����S�,K������%�bX��@Dy=�ߝ����]�=pinX �̼�&D}.8鋜�uغK���<G.v:��t���ٞ4d�;4l��q9�����o�:�^S@ug0��5���]��t=]���y4p�]���Iý��Ev��@Z��HM5O8��<�"'�<C��S�����r�������ɜ����8�0ږ� Cb#��Ő�$�۵h��䒧���KffCnf쎘R]��E���\�k�:5s.��psp�$�8˩�	�]�.z��N����=&Re�v%�bX��wx�D�,K߷�S�,K������Qg�2%�b_�~݉Ȗ%�b~����.�ݷfY����<�bX��of�"X�%���wÉ�Kı/�݉Ȗ%�b_>����%�bX6}�ve��wmۙ�M͚��bX�'�}�'�,Kľ�wv'"X�U�Dȗ����<�bX����S�,KĿ��ɗ&�e��2��Ӊ�K����3br%�bX�����<�bX��of�"X�%���wÉ�Kı,���ffI$��R�0�؜�bX�%�ﻼO"X�%��>��O"X�%��{�É�Kı/�wn��K�q�����}��0�3�uղc��b�����kע�<%�N.'0���7BSs�.��f��Ȗ%�`���jr%�bX�}�|8�D�,K��v�ND�,K����'�,K���L��˺d��n36jr%�bX�}�|8�C����~S_"yĻ��ͩȖ%�b_~���yı,���ND�,K���eɦ�6[�w2����%�bX�߻�jr%�bX�Ͼ��<�c���{��59ı,O{��O"X�<ow����H�쮝�7G���7�ߕ�Q��7�߿���Kİ~��Ȗ%�by����yı,K�s���Kı;�K�r�Gn]�����<�bX��of�"X�%���wÉ�Kı/�ΛS�,Kľ}�w��Kı/l�fv�ʹ��i�a+�5l�#F=vޣN��yD�ԌKa������������﬌��USM�w�{��7���{��O"X�%�}�tڜ�bX�%�ﻼ��L�bX�w��S�,KĽ>�~ə�6e���v\Ӊ�Kı/�wn��?$r&D�/����yı,K;�۩Ȗ%�by����y�2�D�,����3!	���6fmڜ�bX�%����O"X�%�g�wu9��8/L9�>�xq<�bX�%���ڜ�bX�'ޟ^�74�mݘS3ww��Kı,���"X�%���wÉ�Kı/�wn��Kı/�}��yı,ON���\��L�M��n�r%�bX�}�|8�D�,K��s��۵<�bX�%����O"X�%�g�wu9ı,O�_z�{��\�̱\=:���x�[��n��5ҭA��ۄe�+Z��X�wt�=�bX�%���n'"X�%�|���Ȗ%�bY���ND�,KϾ�Ȗ%�b}�/sw.���̶ff���Kı/�}��y�c�2%�g{�u9ı,O{��O"X�%�}�tڜ�bX�'s�~�]���ve�n��Ȗ%�bY���ND�,K�~�Ȗ%�b_{�6�"X�%�|���Ȗ%�`���ٗ7ݷs.d�wu9ĳ�Q�(lO�����Kı/��ڜ�bX�%�߻�O"X�^�O`�5Qg"rw{���bX�%���ܙ��fXn�.��8�D�,K��v�ND�,K����'�,Kĳ��u9ı,O}��O"X�%���M�Kwse.�	3qX5ɮfY6�e��ۉ�I��y�F�vkg�����l��fl)M��v��,Kľ����<�bX�%�w��Ȗ%�b{����yı,K��۵9ı,N�}{|��	��p�fn�Ȗ%�bY�{���bX�'���'�,KĿ}ٻ�,Kľ{��Ȗ%�bzw�fr���\�7���Ȗ%�b{����yı,K�ݛ�9�����ؗ��oȖ%�bY����r%�bX�vw���ܛ-�372����%�bX�߻7br%�bX��{��yı,K>���Ȗ%�b{����~����{���~]��O
�m[�"X�%�|���'�,K��@�N���yı,O���'�,Kľ�ٻ�,K��O��$�XH�g�㴟�a�4�&�ݶ�sւW�v��\6�Yz{V��9��n��u���F\>u��6v!�rU�<�vk�����V0�S�2uۧj���w���'����\\�������Yc0�N��r��*u��cq�+��ԶhK��]n��z1	�̙��6�l-��/����Uv�ǃ[lI�yx0��.���Ս�嬯<ݻ�3X�d�����{xz~:u�
,�>�!�.1u�[��`:�V�C�V�9%��e�if�$�BI�e���O"X�%�g߿�S�,K��߻���%�bX�߻7br%�bX��{��yı,=�:e��wm�˙-��ND�,K�~�Ȗ%�b_~�݉Ȗ%�b_=�w��Kı,���"X�%�}=�;�36��Jm�8�D�,K��f�ND�,K��{�O"X�%�g�wu9ı,O}��O"X�%�g�׻32B�
Sfd݉Ȗ%�b_=�w��Kı,���"X�%��wÉ�Kı/�vn��Kı;�>��sL&�م33wx�D�,KϾ��r%�bX���|8�D�,K��f�ND�,K��{�O"X�%�ߎ�u�fő���<F�e��q�M��<v�.��c&e	��7v^�r�6J�
i�j�}���,O}��O"X�%�}��v'"X�%�|���'�,Kĳﻺ��bX�%󳽗&��e�Lͳ3N'�,Kľ�ٻ��qQ
�L�by߻�Ȗ%�bY��u9ı,O���O"X�%��t�f��7���l�ݻS�,K��w�'�,Kĳﻺ��bX�'���'�,Kľ�ٻ�,K��>���܎ܻ�.��<�bX�%�}���Kı>���q<�bX�%���؜�bX�'���}��oq����o����g���ND�,K�~�Ȗ%�b_~�݉Ȗ%�by߻�Ȗ%�`���jr%�bX�ȉ�:~��͓rk.�lVɞu�+�V�K�M����N����CqFU�s3��N�Y�Cw�����{��7����v'"X�%��~�O"X�%������lD�߻��$�I��ݙ�!ͅ)�2n�$D����ȝ�bX?}����bX�'���'�,Kľ�ٻ�,K��oO7t�m�p����yı,���ND�,K�~�Ȗ?�|�x@P�O^��%�M؜�bX�%�߿oȖ%�bz}ٙ��wL�2���f�ND�,K�~�Ȗ%�b_~�ݩȖ%�b_;�w��K��TP����Y�#�Gԏ��7�5ʌ�L��4�yı,K��;���bX�%�wx�D�,K߷�S�,K��߻���%�bX�G,��7nɹ�仦%�44�v����dRv�g�T�m>ɭ/+P���u>ﷸ��{��?_����yı,~��ND�,K�~�Ȗ%�b_~3�S�,K��>���܎ܴ��7w��Kİ}�{59ı,O���O"X�%�}���ND�,K�߻�O"X�%�g�gL����s,�٩Ȗ%�b}����yı,K��wjr%�bX�����yı,~��ND�,K�{�w&\�nHf�)�4�yı,K��wjr%�bX�����yı,~��ND�,��U���AH�؞���8�D�,K�N��32B�
Sf�S�,Kľ}�w��Kİ}�{59ı,O>��O"X�%�}���ND�,K�ߧ:��u��۲j��F�������:`�`R��S�W3�ힺ�ˋ��{Eg�Z��ߨ�%�`���jr%�bX�}�|8�D�,K��ڜ�bX�%�ﻼO"X�%��gl��4�s,�.fl��Kı>���q<�bX�%��;�9ı,K�~��<�bX��of�"X�%��g{f_ɲܙsn]�8�D�,K��N�'"X�%�|���'�,K������Kı>���q<��{��7���w��=<.g9]O��,Kľw��Ȗ%�`���jr%�bX�{�|8�D�,K��N�'"X�%��}/�˹�vap���Ȗ%�`���jr%�bX�{�|8�D�,K��N�'"X�%�|���'�,KĨTxVW�qI-F_��c ��&�K(4�� �LV0��Hi+���<!-E�����1�>��*ł��c	.M҂�(�R0�@x���$A!�"�O"P���`�v0�� �|t��)J�
q�% �'���3}���wwM��v����gLbx������(�[s�۞�ֶ�Y/ <d}�Obڴ���A��	%A&.880R��'a͒G1=l��]�Q�ĕM����f�Y��커�[��>������5���1�EW@�4M�X5��n��»2ڥ�v��n�y�Q�U,��o��v8m�����`�%�ݹy���jvg!�F8':�M�t�7�Z�ӛ�[�l�'����.ԛl�mm�mݞW�ss�v� ӥ��Y�"e�ۃ"6��`�	�ō-��%A����2�Z�@96�ȸ�k���>-J�<9����n�K\ ���:(7<�C�j�	UU�pR���V�f@^2U�RqO8n^� �[O+r��Ys���7=m�6��nlյ� �d����6�u�4m�D��m�7V�&�J uZ�CjV�N׉�Û#q[>Ԅ��
�t�p��z�Jt���ƕ�ܴ���❞u�q�ܝ�:��kL� 0��y�rl���.����fK3�*����a7�%w���q�jUcʜw5O�U]۬�9�m�b�Cf�g���e"�W����!�`�Ҡt�m�c�X�rtN��y��"�p�]���L X�i6�p�)b�F��ݭ�+�J�e�3��WK�a��xםy���:M�nY$�͎9{;/�K���T�B�;;=תU'j��k�!2��smE�w���Y�@G�^U8���=�����Z]Ol��R��=Ix�X��
�96vz+�kI�X�J`�ݖ���DQUP���.8l5�u֮P*��Õ\v]��8[��|��N�4m"t��;`h��v�]'+Wm.��1u��� �͵��E�1!�r:�3�ݭ��q��8��4� O@��x8畈`�^��-m68�g�5۠+� n���ۘ������kg��l��	�ǲ����r�B�C�Er��v����F٩�Ar�	��f�q�\t؆�O�|��,ɗ<�:���=�D�D��Ds�"'��uOD1@>UC��@<�NO�/k{;[���]�ͭ��Q�Z;=���'*��'��=s���8��We�a� �#����9�R�I�>m�Pܗm�@�� ��c�۔�Ƣ�� ��(68܋��.<��T�K������cl[t�
�t�kɭ[E.%OG97�M�wmØ.�94��S�8cN���t5Wzc9D5<�n.��ʐ�'R���>���t.S��T�GD	N4&�Һ8iK7a,קҦ��u>�n��y.Co�|o�~�gն�e�f��O�%�b}���'�,Kľ����Ȗ%�b_;�w��Kİ}�{59ı,K���ܙL۹!���.i��%�bX�߲wq9�H�L�b_{����%�bX?wMND�,KϾ�ȟ�C�Gq6%�gO��ff�3aJl͛���bX�%�����yı,~��ND��dL�߻�É�Kı/���q9ı,N�os�n�ۻ0�f��Ȗ%�`���jr%�bX�{�|8�D�,K��N�'"X��̉�����yı,N�����4�s,�r��ND�,K�~�Ȗ%�a�!��?n'�,Kľ����yı,~��ND�,K�O~��ṷw,ݛ�����R*�K`�N#�-�s��ݪI�&{,�.��e�2�ܻ�q<�bX�%�㻱9ı,K�~��<�bX��of�"X�%���wÉ�Kı>���ۆ�p��ɘn�ND�,K����'�����A?"��|��K���59ı,N�~��yı,K��wbr'�TȖ'����r;r���&��Ȗ%�`���59ı,O=��O"X�%�}���ND�,K����'�,K��ﳦ\�wf�̹l�٩Ȗ%���Q(lO�����Kı/۱9ı,K�wx�D�,K߷�S�,Kľ���ɔݻd7r�ۚq<�bX�%�㻱9ı,K���<�bX��of�"X�%��wÉ�Kı:�ܼ۷ W.qV�fu�L�7.��v��ۮ�Rqz\\�zC�qtVW�l�㎳�ow�,Kľ{��Ȗ%�`���jr%�bX���|8�Ug�2%�b_�~݉Ȗ%�b~������0�t�!�����%�bX>�����bX�'���'�,Kľ�wv'"X�%�|���'�,K�����r[�d�%�����,K��߻���%�bX��݉Ȗ4ϖ�P�D�E����< ,"�` @B���@1T�,K����<�bX�'���br%�bX�v}�����[�36e�Ӊ�K�ʯ�*���ߏ�؜�bX�%������%�bX��w�'"X�%��wÉ�Kı=�N�n��p�wrJf��,Kľ{�w��Kİ�D?�xbyı,O���'�,KĽ���ND�,K�t�v]�ݸnM6�ݻ�I�g�"����ҩ�-���1�V�k+�EZ��{�ܡ���w#�)vL$���=�bX�'���19ı,O}��O"X�%�{��؜�bX�%���x�D�,Cw���?����%J�����oq�~��r&D�/br%�bX�߿~�'�,K��׼*r%�bX��߳�2��J�̔ۚq<�bX�%��wbr%�bX��{��y��B"~��§"X�%�������%�bX�t��ffI$��R�0�؜�bY��������<�bX�'���*r%�bX���|8�D�,��Esbf|wv'"X�%���:f�&�7$����O"X�%�߯xT�Kİ�@B?}�ޜObX�%�t���,Kľ{��Ȗ%��{����n��f.��\��3rF�����5�S�)�y�:�S�u `nvw7wt�Ȗ%�b{����yı,Kߎ���Kı/�����%�bX����ND�,K�Ϻ\�l���37��q<�bX�%��wbr�r&D�/�~��O"X�%����
��bX�'���'�?�*dK���3sn�˷IL�wbr%�bX�߿~�'�,K��׼*r%����>���8�D�,K���v'"X�%��}/�˹�wp�ww��Kı;��
��bX�'���'�,KĽ���ND�,K��{�O"X�%�g�gL���w2�ɛ�ND�,K�~�Ȗ%�a�G?t��Ȗ%�b_~��x�D�,K���br%�bX�EE���ZN��7v�u�ss����G���//l˭v�:�َ��us�;Ga熃GT<e��շdrvo[�[�}��ؽj컦E��
ǇF0����� n�{n�;J[n��a.)�Oy��,�㝭k��[�����z�s�9ey�&�=��&��.�ݗ�T[u������T�L1�{)��N�4i�����Fs�n.�LB�f[wr�n�M�Qq
d�5�F�7Hו�vjgtU��y��o-�77k>h��������KZ��Ht7}��%�b^����,Kľ{��Ȗ%�b{>��ND�,K�~�Ȗ%�bY���̸I%ɲ�نn��Kı/���������blK���LND�,K������%�bX�ߎ���Kı;�Ι��I�f�37w��Kı=�of'"X�%��wÉ�Kı>ϯwbr%�bX��~��<�bX�'��9���Ir[�.l��Kı<���q<�bX�'����ND�,K����'�,K�A?�B����jr%�bX�O������-37p���Ȗ%�b}�^���Kı/����yı,~��ND�,K�~�Ȗ%�b{��~x꧖�]Z���!�s��{On`�]5�#��Sƹ�a�n�Oa�:Y���gl���,Kľ{�w��Kİ}�{59ı,O=��O"X�%��}{��,K��}/�˹�wp�ww��Kİ}�{59
���A�T>�Mr'"X����'�,K������ND�,K����'�,K��ﳦ\�wfݳ32nl��Kı<���q<�bX�'����ND�,K����'�,K������Kı/��gL�n�+��.i��%�g�U��;���br%�bX�����<�bX��of�"X�%���wÉ�Kı,���f\$����nn��Kı/�}��yı,Nϻ��,K������%�bX��owbr%�bX�{��3wnn�ܹ�M����k:�6�]��Ox�q�^�d�Sn#r�;�d��nI33wx�D�,K�����Kı=���q<�bX�%��w`~Ay"X�%��߷��Kı;���9���Irۻ��br%�bX�{�|8�D�,K�㻱9ı,K�wx�D�,K�����Kı<�������-37p��Ӊ�Kı/~;��,Kľ{��Ȗ5OAc�N�p�O"l�19ı,O��|8�D�,K��;�����ssL30�؜�bY�=����yı,Oӿ�br%�bX���|8�D�,K�㻱9ı,O���ܻ�ۗf	77x�D�,K�����Kı=���q<�bX�%��wbr%�bX�����yı,K���I�i����)��u�P{zՓ6�D��Q4�d��.�������܌��h˙�wLO"X�%�߻�É�Kı/~;��,Kľw��Ȗ%�bv}���bX�%����6lқ&��Ӊ�Kı/~;��,Kľw��Ȗ%�bv}���bX�'���'�,Kĳ�׻2�!.M��L3v'"X�%�|���'�,K����19��"0ș�w��Ȗ%�b_�?n��Kı;�Ι��I�f�3ww��Kı;>�ND�,K�~�Ȗ%�b^�wv'"X���V���D�w��Ȗ%�b{��s�[�d�eۙ��S�,K��߻���%�bX�ߎ���Kı/�����%�bX>�����bX�'��oߏ�&l�3ss&��d����x�N�(��q��h8�P�r�$����l�3l���3w��=O�X�%�{��݉Ȗ%�b_;�w��Kİ}�{59ı,O���O"X�<oq��;�^���z���{��2X�����yı,~��ND�,K�~�Ȗ%�b_~;��?�ʙ��t���r;p���&n�Ȗ%�`���59ı,O���O"X� ���/�?n��Kı/���y��oq����o����f�V�U+��Kı>���q<�bX�%��wbr%�bX�����yı,~��ND�,K�{�t̛6iM�r�ni��%�bX�ߎ���Kı/�����%�bX>����bX�'���'�,KĨt�(�e��s6mծ��W��2��⮥[�1�l�8ʛ�C����jȸ��G@����N����hnGBh�����z��;��M@<�8լc��f��\w+Z������*v�gnm;u�����&*��g<Ŗ�:9�@�C�C�8�W3OY٭��C�x�G&���lS��x;NN[;	��\��
�z���l�3�ïn�wN����˲O<�nܚ��n]�Ȥ]s�q:�6�NlG�x�t��c��ey당�7ve�I��)�݉ؖ%�b_�~��'�,K����S�,K������%�bX�ߎ���Kı;�Ι��I�f�3sw��Kİ}����?�A#�2%�����Ȗ%�b_�~݉Ȗ%�b_;��ȟʮTȖ'��annBY�ne���Kı>�xq<�bX�%�㻱9ı,K����<�bX��w���bX�'���y�w	L��s7w��K�� >��v'"X�%�}����<�bX��w���bX�D�;���'�,KĽ�Oٻ��n�74�3݉Ȗ%�b_;��Ȗ%�a�!���SȖ%�b^�����Kı/�݉Ȗ%�bD>�v��d��]T�i۞@�qZ����1]�q��Su���ܺù�-\2N�<Y��k���ݷ{߻��I�����$BA����ؖ%�|�{�O"X�%����.nl&��˖����Kı/�}��y ��AS��'"X��݉Ȗ%�b_;�w��Kİ}��59�S"X��{��ͻ)�s�sw��Kı/�?n��Kı/��w��Kİ}��59ı,K��wx�D�,K�O�ve�7ZSf��,Kľw��'�,K������Kı/�}��yı,K��wbr%�bX����L��$ݳrI�����%�bX>����bX���w���ObX�%�~��v'"X�%�|�{�O"X���~~w��s�n:u�;^���l�ÜH���Iĝ^^�t�ۘH�ݸh�j{X�gv�,�˺jr%�bX����<�bX�%�㻱9ı,K�{��yı,~�ND�,K����<ٻ��3w\���yı,K��wbr%�bX������%�bX>����bX�%�ﻼO"~L��,K��������ssL30�؜�bX�%������%�bX>����c��H��=�	$ �� ��D�B�|	露�Z$F��i�苄A"Ƹ)��(,B�F n�LP�G�b,@ ԉH2TzʱBK�b�H�`�b��M��K�*��y�Èqb�V��:�H�"�#B����!äc FHB���e��$�ЄHx��Z$�qI	jp�b���HHbE!	GLX�a��YR0�%�!��
$��ŀ���@ۂ�")0"x�h>%DX�'���� ���V��o���> �POaȞD����Ȗ%�b_~;��,K���/�˹�]�\���Ȗ%��2���Ȗ%�b^�����Kı/�݉Ȗ%�b_;��Ȗ%�`����.nMٷne��jr%�bX����<�bX��G>��v'�,Kľ���x�D�,K߻�S�,D}H��Wku��E
R�r L*�y/U��1�.1ȷ����bq\�r)�3rź�ٹ�ɹ���%�bX�ߎ���Kı/��w��Kİ}��4?�y"X�%�{�x�D�,Kώ��2�	��!�݉Ȗ%�b_;��Ȗ%�`��xjr%�bX����<�bX�%�㻱9� ���&ı?�o���$ۦ�3sw��Kİ{����"X�%�~���Ȗ%�b_~;��,Kľw��'�,K�����0�7!,�6ff�Ȗ%�b}��T��'p�[S@�٠�f�a$0ހAJ҈A�I*��P&ɆL�S*}�R�6���I�C���O2�ֳf��$����/7�P�۫��}^�`/y���"i	�Q�i�y�+��{3[p���2+����S�v�׶4n����RN ww���sn�fmՀs��,�K5�Ϣu�0RKy�K���t�*@�}�[��6����u(���$���u`�f� �f��ͺ�1Ǵ�"�QДdʠZ͚ �f��ͥA�%�(�ﮬ�ח�4����Lt�fl�=y��fm* ��٠&M�$2a2X�/�������0�	t��2�[U�Ƨl��3��62�q�����TL��mZس���;��~�mB��V�gٷa��]v���\m��$"�u��ss�N˹����lleOG$7m[l�l޸q�Y�
�`�s�i�LkY0ѐ!����\p�>��v:%���V�B�n�]W�s�6��Q�;
�]�.t��GSqҍ���I��wb�B3���ﾏ����g:��5���X�=P�:&���=<c�����1�M�]v.&拶�ɲ�vߟ������T�7��@���������D�2�fm*���^-���9�۫�n�up�Иܔ9%X:����G����ϕ :O� ~�sn�C�0m�,��,w6���f�X~����`{]-�Q�D�&	��X�*@kqR �s�1 l��٬��5̘K�Z�fą�<�k�g\W���۵��p�v�u7#>��NU���Hy�@����9�A2�T�&""G�T�͚�d�cf�$̒����{��/7�P��T��[� 7PT��`��`s��V36��9��`gi��r)A�I;��@o8���Hy�@����t�S⛢�*��f�X��s}8��K�ͺ�
�uZ9�G	:&���*�F�z�m�zp���m��q��Uu��h{��BGBcrP�`�l�fl�9�۫��u`�X�8�II�)ӻ����@o8���Hy�_~��k��j3��0rK����fn�x��� ���yɞ������ �bͦ�J����$� �f� �s�1����avfz�Hi�%�f�=y�@|���=�t�͞,��,����pi(�)��"6fQ5�L���km�c�\m�t�6�2=E��m��*�rX3vX�M,��,�͖v���"�H�&����y��@�b �& ���ڟt��p��l�w6X3vX�M,�M��GBcr|9%�z�f�=��@z�t����I:�KS�y,:�OiԔ�r�6��و����� �}��y�@o��^��[4mtX&��C�<�eٸ^y��G6�cn+l�ق�#�Iއ��vZ�m�����7���վ��b ꞟSn?�IDbh��͖��� �we�����$u��d��$�Nb �>��&#��ꪯ{�τ ���x���(n�S��9��`s�4�w6Xz��o���O���R�))�6ܖ;�K���N w7��9���I�' Q�zXB�w7r�M��L�/Z6�������}�]yĴ^��u��������=��p��d�&
Ny�s��SV�$`i��Uvy�G#�aZ�t)1�N�t�;�tF��f۶
�u��g���������չ�ʘg8�Hi�+��$W^Ӷ��
������gZ��uix�m�5��Զ^�����u���;v���.x�u�g�\�̗�w!]���l��v� ����{�����-�=���J��F��ݷ��D:uK����<��~�����
^�x�w���I�؀7�����վs�V|o����*i������ �f��ɥ�s3e�4���:�'�DD�������(��2gr�zh���륺�ϢtA�a$�;�t�5��y�@�����]�_�(R�Dp��l�?.��p��K�ͺ�7L���/��r|ۂt�78[�b2v{�5v�]7����o\$�v���Yutt%�rX;�,��,w6���_}�n�X�O_����
���=��T̡2C2V�S2�.�t�nl�;�,����"�8:I��9א@��{�9� �}� E��j|�:PN�͖��� �n��ɥ��3i���*��I,�s�1������T�=웖�N���8չ��a=�.E�us\k�;]:��SXz�����0]����� 7�A ks󘀒��Y�}��	$�9ܚX36X;�,��,��6�q�*J#Dp�fl��6h�[�lfM���K�l¾�M�ߧ���l$U �%�rX9�@���� ���{���W/�6������fl�9�۫ �f� �se����CU	�I ��A���YՐ�.ݳ�]ZG��g��[q�ܬ��=�=��9#(����rN��]X36X;�,�͖n�ܤ�`$�@mIT�͚�2fL���zh�zh^m*�n�uu$T&ӓ��,�͖���=�]��Հww��0�oi�t�o(�����d�|�Dgw�@f�Ԩٛ�����S�~��o$����M��l��&I`s��V�͖��� �f� ��MjqD��%E���M�)�sz������n�p�J�p�m6�s���m�Β���$� �f� �se�s3g�����UU���u`y��lqHJIF(�b �s�W������ʐ�1���Xۊ�IPT�ܖ�ݖ;�u`��`�l�3���9#(���xy�����oyPn���6h>w������z�&㢒t�6�� �f���34^oM�gtH��T�2fL̕��E�������"���TW��QQ_�AEE�"���Р��� �`�`�@�"E��EE�"A �PH �DU@��TW��TW��QQ_�(��EE|QQ_�AEE����*+�((��� ���삊�������b��L��t�ǢHv� � ���fO� �� @                       <" P
�E���R���R ���@J�*���T��*HUP

��H
J���   
      � � )A�`
	� �����=��h1  �@
D
R���� R��P  
"����;��Pɪ}�7=�k�et��]�ӻ�W�o�};Ů�rj{nm� ��  R@   1 �Ԗ�{槖�h�̺�wS���{�g�W��{��x��� G=/q�)eݼ ��Κ���_|}S�n��N�ܽ����r� 4L���erqK}�K��{��� �     >�B���}o��O���{{����=}w��X }��s����ܰ��Z�`юS-ֽ<lx ^�&��o>��W��X���^/v�qq׭�W�x �-ź�\ws�+ͪvr�k/ >�P �   ���O��[nO�ʮm;i��zܞ�`�ަ㳲rӬ��K��&�� :��v     D(�*� �Jɩ{�uM��sn����� ���>���w����_[�)}� >�(
  �
 @4�>�z������ޝy���ϓ�,��@w�,���9|���<�{�x�:ox _=�|o������ ��ӯ�Y�4�  �E)HJP);@(� 	� �����i�E(( =AS{IR��D �U?�M5S�T�T   D��RS�6�&F@=��&Ғ��� �U?�	S{R�J� h ���IH� )�Bq���������_�o��u33*S�mF<x���TWA��DTW@PT��
*+��
*+�(��QAS�?������������&&�o���Ç���4��d4o��5"���T�;�}���p��#*�B��$���H�$B4� Q��Х�h"E�H���$��-0��I� ������d��a59��q��ǰ�dXE$R,�!GC"@�!�SAsW{������=��v�v9�=�}��ݳU���,4����7nNcP�9�o8BVm����5���|7�߈baHV4�T�w*J|B�61"�v;��(D��!n!��K��!����s[w��T��L6 �2�3C	�q(7�a��41�$��c �4tB���.%0�HY��h�� �4l�
��m�f�K	
Q$�"BIG$�C��CF	�ެ�K�[�ɟ��z˝�}ǜ�7���7A����nl��L���YLCBG��B���5�4��:`A�E�9�,��ﭴ��K�����ެcZ�`@�&0�)"Ml�HX\H@t2�xn$��JJx�0�+��tjn\���X�1�Lp�f��ɫl�w!�s휓,��d���"�Ģ@��vqYC5�`E�%�t�6�l�of��i�|��K�لi��|c.G{�aL`�%��rt�,�fI;��!XX�ȱ�¶R�Ys.��O9�3g���p������O�Iۨə9�������&jCDJc�٬�ֵ�}���!�`A�H��a�Gɣa䐁!4*1�ƌ}�~�o���`>�!����5ô��%-�y��:a������Mɠ�*Bh��|o l�K���bK]BnG���~�ጴ�p
$j��Za��>H��D��HƤ#�x�d�voF�d�dv�J!p�B᪒�, ���3U��p��m�Gc$.i��ݜ���bp4m�%���B#X� AT�60d`M8`B�`əY�NƀȐ�T�K��!XY��Q�	���"JB��)"J�����h��0"�4�M,�	7��n�w�h!p�#H�h��B���$F�W�.va �R�:�4�a
B�J�na[s_�0CD8Ů.�4q��s���G
A�
�IP1��"j!M$vT`�Fȑa���i��|+��m�Xӈ�<H1(D���lӎ�
h5,3���ZVV@�8H^�K�;�3T�)l)�C[����W��nl����C�B��h�c7~@�:l�B5�|<�X)�4�JA�M&%i�
��$h���d��N�D~�CP������P��LHЕ�
koi�0 Ӥ���C�:v�+�����e%�s�5��\�K�����4�r?e����/�e��������A
a�7��L������>����&�]�.Ƒɮv�$g.a\�1>M0���	s��4s�oL��7�oR̈́�)
�t�%l`0�� �od�!��t�aH�F�6Jon,٦�{�30��)/��0�F$�L#�p�q�i��1�7�-2a4K2k-q4h�2��o%e%�r�!
&n]�;5�gt�.�H�}��jl�o��t�˾N�9�c/�;9i���Mo]� �Z��D�P2�(S4$�) ��i�Ȅ V	q ibQ�EH,$��\���Q�6�����4����\��kl.3
�! �H\SS7�$vk�l��4�#w�r杼�&�s{�5�I�	-�g/[fs7�fl�ޤ����z��N����X���!�*A(j�)�n�Lt�7\tl4˚�� ��:ĀH��W�K�Cx'^k�R����9���5%�$���\�>���7��5�H}Î�5�3[��(Fp ����������of�	�a��[� �7�\u�) f����7���ϰӾ}��&>���aB$`@��8��H,hvs����D�F8Ῑp;L9��@�ѳ�c���.���ٯ�.w�}��&3'^��!�����Ip��i��.<���K���}��JJ���6r�95�f�v�`E!�P�.J$
���P
�j4#]B�
�

+Jh!F�F�/\>H�!.�J1��$��L�:jWS�h���.�HSWBWH��4�� � W!���9��Xas;H��
B�2�v@i�%��
B܆a)��S3[%�*dB�,�Ja�	5�Z��aL4�R\�C6f��R�f`\��.��ȗm#27�0#��0��F��p�K5���%�|6�f�N^�M�!u8M�l�%���.��$~�!q�aR0���o�'��0��Á�`m Cd�/ҙ2�q�5��qH��q��F�xi��sP�(�ʒ��Z��4i�T�@����!	Hj����t��
��,�9�rk��G��n��#
a1����)��ϴO���H�c�Ç���!)���$�6Ȥ��YCHH���4mC��5B�������� �I�(@ �rI*8
Fɠ#D�M���6�xD �"iXHȒ-$#P���B$�hg7"a�oa ��:f�f�@��1Ԛ�I6�a\ky&�F,�.�8�� �D�a"1�$�v�mB(���L*f�D���l�7�5XB�(k��SR��
8���\��7�ji���c8&b����ċ �� Da��H�����2B�.���1ѽ�Nԡ&&�n�"c�6p�Ѱ�ą�3��*�2`�a P%4laRH���!)f��b����	�C�0��Ry�>;(H&��B4q4n2�P���1�&D/�MKf�wK��q�CP!�,��\8n��zũ�� p:�i�]f�5d)�����X41M1B��40��DsF
FS�7EdHP5��!RT�4A����:�`�$3I�2F�)�H�͐�#0#�B�t]l'ЄFZ$J��`��
.�.0�
��b�x�>�@"hb`h!u�`7�77�[��Y�r0�F?4���~�Ĕ���˒���)�)�Ģa�o�6���ț�n����p#�4%v�B#@�6°�P��.,nkz���C7��B�Ա$0�\����(�ѣ���9NsiVR�7�]h�3#�@�YB[���i�a�=Q߷�hѯ��'�^w�f�;�gx�Z�@�5~8�xT�M����H�����!Hp�KhA����Љ�a��Mq�h���a��^ �P*`ԂĄd�YD��$ђm&�F�,5��ӄ4^�"�+�lP��x.�'�B!l$�C�$�j��ۆ�������	y$���$��,����dH�B4B%R�	��['Ӡl�~�8��@#�k)�_�7����a����#!
&܉a! U���!Wf�d F0����m� D�n� ��`:0	�M�)��I`�A4�t�`P1�V��#"�%I!5i4h6q��I�.ݬ������|����S$�����!�I�
B�JL0#�6M�80ֶp� @��%�$Ӷd�BW�x��5e-�$�3v�P� ���$�.��#D��F���5���-q�L�s[#hA0�hL7�f)�J�����FЍ1Ðj��$!���V�Mh֜��P�������&��L5l܈B���];X�	�I���p���BPe�H� T�$XP�v|��(k�f�Y&��d!����!��r��L!��%˧\�y��gRI��e�%��覉�xCQ��Ebh;��6; \$ѹ-��O��������  �     �    � 6�  �    �۰� 5�$�v���$H�Y\��)TUT�p����  $�[l�ݶ�KRqn���6�݁l��r$�5 ����msI���NZ�vYB�;�UVQ��n5̫Q����,�cq�j��	 �M�x���Vs�t�rm�M#� � l�[@��"�խsm�  ��-H 9ն@�݀�p	kn��� ��[R����$��k��2wbm�m���� �m�v�����Y�� 6� �T�jB�g�
ʽV�m'�I��[�IM�/Im�dKt�֭��  �[vسNѶ�  $Xa��@ �-��  m    ְ  � ��  � k�6N�� �`m��jنLP説�7mҨ�s:�F��a��m�x�����J�@�	�=]>j�ݰj��*�r��KmUn��][[.�]"a���4�:I��`�ŷm#U�.)u�	V�V����Zڪ�:�:�N$1Ͷ:4���� XZ�)N��-�n�@4l�[+$ p#��Y( ��-pm�A[#e���N������#�[M�az��U��Ŵ:@m�ŽV܀H	m�&�&�nm��9��@ H�-��H�n�-�UM�Ĕ�K��;A��v�Ij���^wiR��Ԁ-����%	׆�8�u�۵���P!m����ۍ�i$I� ����-�mK�ʪ�z�)I@��l9t��%^��(  ��HK(-�9�lm�6� [d$/X]�.��sm��0�Aa�'8 6�e�m�� ����(�6�cnZ���l��9$K 5�C���� �HE�ZN�8ְ6���h�7Eogen�hk�6X-�-�f�O�}zԞ���6��I<�bF�C� ���gZҥL�� ��5�0�ƶC��d� �`%�U@��C5g�
४��ؗg���U��݀[Fݰ�������`.���J��r��Um�UU����Z�ɱ@*�@'�prD��#m�������<�UY��]�^����WR��A=H�ڝ���9�p9$��I��S�I�UJv��Y�d����2;-�����[b�RZU�Vye!�\�yԥ��XIm����P'f��
��|���]*џ�4 u���!W]����/@x��weBk����]l�f���[�������b��^e5�vY-$7[%G��N�
��m-��we��Z�R�.i�i;2� ���oT�L�޽;��r��j��J:I$ڶ�Ͱ�ZF��"F�AГU��bR��\%kvxk��� v �����sF���Z+f���52���uY.	����H��Հ$� �m�2-�� IZ���v\ 6�[oN0�z�Y�$m�[C���!ʕ�L��0  s���   �]�����eY���PA�   [M�	���%�4�k�HH� �p-��]��}>����X �� p7n�����  �8�[&y�r�V��浒j�mHڶ��HY�1��Âv�[@    sM�����r��    d��[Զ����T 9oiV�YvWe�k�l��`[R rN���� ��L-`  �n�m�&�%��m�6ۆ� ��X'I'N6�i6M4���|�h�Ѷ�W^@ͻUWmY�8��km��Mҷ. �� �I&׮�F�8 p�n��w[�6� gf��PP���Z��Q��!:�.��[�m3�-h� �1��\&���q�t
�a2+�]�$�c�+A�Բ��j��g��nj�Y}�vP��ꀸ�`��m�m.��c�^����	�Nɭ� /F��޸M�6�66���m�a���`:�:CZI�8��Л\b��[f1��[� �"mr�$��l 	M�b��ֳZtݶ ��-�n��d��-�  ��  � h�\��V��� &��VW�ɳ����h�F�h�m T�R���U�
��Um)(lUT�9�e��:YR8ݲM��&� �� $�  � j�ۖ��:�����@�֥�ZBj�)��N�j�YZU��u�V�U:A�v@�v%Rؖغ�]���R�����-�$  ��ͱ�m"۶��c�� Ŵ\9i	�bvBj�Z�%�J��UT�,J�Y�j�)V�HJ��M�� �v�9�$ ��Xb�e�[m��,��J�H�2 6�BK�lA�h�a�.����Y��*�g�R���[!�u@R���6�E.���j宪�ݭvS��azED������-�MF`ݍ��S�k���d�t�,��+��M 9m<.��(ruYX�@mQ�� Hsm�N���i���p9rTݮ��`8X����U���8%��}e�}/Km�o  j��(
��V�[7]8 ����[ﭡm[J�RU@�u�(v���.ķ 	�i5�w[��7m��)m&�YKG ��z�oPVĜ��ݯV  �KZh�M���ݰLݭ̀A/Yl�Crޕ��� �g5��!�N�V��
���J&I���tm@�UVʁ��3m��:�ԦJ�T���LӉz�|��uג�p�,mUUUJP�!K���!͵�I0�ݰUN��GUpS��9m��Cm�Ӧ��C�k�#/Z�j����l�!��_�ͷ�m�lm&m�6�  [Cnɑ���{���k��T�2�R���U�X�f�[x�7B�nrA!��Mn[͑&�m9@�I&r�YF {	�V����e`*n�y	����� m�mp;';]1zo]�� [�cj�dw6��J��� $��]k�K(�����8���m�� �i06�8�D���l������&؎sH/L�0k��v�i���e帤/ ʽ,U�Rh)j�~n��]� -�ඊ�zڭ��!�T�����ia��UT�G[[l�#�� �n�� 	I$�u[n9��`Mi\��햱Ĉ0I�$���6['�N����M�� 9��ۃ�Z�]^���i���h&�q��H �6�-�q��@z�����)U���^�`�r��[����@�Wh��Z�mP J�Uj��X��P *ղ�7R����Um[z��6݀	��[%��r�[PT�v����L�e����P sm6괃 �sm���@���Zڕs�?.�*<�, 'cb]���*�W��[%��d�.�'$�H -�l�a 6�M�U`-� ����z� ��ڤ�p �`
�K�+�R���U[P$��m��%�p
�V�r�UT���.�t���v[m��KS4!rڪSf��V  $�m[C� u\Cm#v�   Hݰ $���X kXlY˶ 6�$   [m���5n�hěp9��%H"�9�i���8   �VVN
��$�V���`  �lA!"Aԣ�J͐p d�@R�Ĝ���нm@ ��κ�M� H [Sj�H��l[Gj��S�
^Z����Im�ku��4P   ��� i��k���킔H $]��J���(.�֦��m�-�:uN���ѻUW6U�VX&�m����@�b�a�zϾ�Ko4� �f�uq�]؝�Ku�R�l��� d��#&�Ͳ���/-TR�` �Զ�t]t� �  �
��UUV�@|��]@D�hHm�T��խI�i$� IH /[7[��R�Rҭ`��@����z�t[��VU����@p��  �l��nG8�X���|���n�L8����(��e�P�y��H�|��f  m���7iҶ [��v��үU]++UUJ���M��m@U�[ uT�@����6��ۇ6�F�C���r�-���`��[RR�Km�l �i��kx��Àh���[@ �%�ml��ホl,�$ 6��p M,���[�Ò@�UKN[g��~H�j-��M�@(m�� msm��"�[��M"M�&���V�p�e� 6���]!�H�����   ��l��6�m[A��8��s@U*��KU!5=j˱ҠQa�U�L�UT��kX�[��{t��vvj��-]�-�М3m��l[�l��܉� �kz�,L�  䀐�@ Hݻctj�5�z���j������ӥٶamm� kX��2R��&�}��ְ��;i�pm���X8��f���u�i3r�im��lE vZ��U��4+U@�l$�    6� 	 �5.��  ��i�#L�5��kZ՚2��������B"���D�\W�?�L��TB��D6�%�T0CB)�S� c�t
'1@:2?*�P�8�E��;Q�(�-��w�M(�X���W�PF�.�"����	��@�P��*'DW� v����A�����U�"���U�W�#���t�7�A��z�tT�/`/F
1#���^��@"l8"P�pE1���Q �
�{��S���� _��J!��D	$P�F��`�0b*H��  F1`@#�W�� ���H�DCS��>p@�'�/@��z�lM��V��+��� ��X�tz*)�G߀��ttP(�RO�b ��<AM|#��)�t�U>(�=@~S �~оA_�N�Q=�j&�P�4	��U<.iv�!D��4����~A>A򈟕G� |u� *��x��((���
����� sl�H��+�V՜e�їn/$���bs����	\�J�pQ���uʝ��.���V�tfh�Mk�\f�c:-Ce���e�[��X�'��U�f�4���؂6%cb�E2���C��1q�;Fq��ba&��@�n6��l��=j\di'�D�[f�8-�S[����֡v�7o ��V��^׮���U곶&&6���ygn[�ywetJ�,"Z�!=1l�Wc��ּl6q�t��t�uA��O<Gmq��8Yõ�˷k�Q�z�ѵ%�ܱ����pxJ��P��d�s��Aۉ��cv�өv� W;lA֪������=���­��n�b�IcR�G��(l.v�6ȭt�Lv�,����:�8f[�v媢gdf����
 Wv�{)5��˨{[Ӆ Bӭv�]��9y0u�`�q���+��f\��6�muuť$�o=n���\�b*����y�D�+"�F=d݇nf0�<��G u��Jrj�;V���N��GqF����`���hu���l�5ٮ��;gv�� �0�ƹ��MG[k^���hv&9И�6X�^�݋!�tݱ!�v�vİ�6�`�]V�4q�2�\`�Z]���5F��l=lL���H��ԙ:݈>�B8���W,��ےs��v��\bjœ��U�u��k`=A��M��x����e#�V뱮P9�7!t�D;:���S��xt�Gs��v��B��ͧ�c���[V����2��֪��L#Gf闫�k�`�j�'�V�����[t�=��s�f��P<l:�N2���[�8�u���� ��Р<�S�y�⮪�H�����]�-{y1�]÷�	&B�����j{e�I���[J�PVȧn�v�˺�vZ���є��u
�5��M�V�Z��м�!/��۴���fӇ��y���sɲ{4v̦�.�(�a��I�հ؈j�{��n�n��#�W�.PC���� x�qDN�P��~;�ٸ���V�;t� ��x�<��wLb[vJ�n�����\��ɧ���n�u�h�;v.u�Ipc�#��9G��b�8mw3��j����������N6��x^n�u.��Y2�:��C�낃R��GwB��[3�F�Ki��ҜLXd�f{m�#��6�my��sN�XQ���B�u�:�:ϰM���m]rG]{۟wwe���l>Wgv^݃prr� <�����ɐ���.��e����k��� �{4�$D��wI�$�r��A����L�bX�����r%�bX?��˛�\ְ���fi���%�bw���!� �W"X�s���Kı=�߹��Kı;�f؛�bX�'��s-3ZԺ5u�Y�-�ND�,K����q,K���m9ı,N�ٶ&�X�%��w�6��bX�=�����3��CE������o�}ͧ"X�%���6��Kı;���ӑ,K���=��Kı9�����Ff�����%�m9ı,N�ٶ&�X�%��w�6��bX���]&�X�%��w��r%�bY��o���W��]-��[�m�ի�.�r��O'Vb��n���#W#=5��ֵ�bn%�bX��}�iȖ%�`����n%�bX��}ͧ"X�%���6��Kı)��e�CW5Lˬ�eִm9ı,�޺M�a�b����Ar�@���"�dMı;�����Kı=�f؛�bX�'}�p�r%�bX�e��W�hZ8h��7���{���~��~'"X�%���6��K�2&D��~��Kİ{��]&�X�%��������2�~{�7���{������蛉bX�'}�p�r%�bX=�z�7ı,N���r%�bX>���]K,�h���&�X�%��w�6��bX�T���]&�X�%���}�ND�,K��m���%�b{=��Ƈ��y�1�40�D��{� m�@�6��QD67Jm&�q5��:�=��2����%�bX>�߮�q,K��{�ͧ"X�%��{6��Kı;���ӑ,K��Ok�nMY��I��Z��]&�X�%���}�ND�,K��m���%�bw���"X�%�����q*K����.35�]Md��iȖ%�bw�ͱ7ı,N����K l�M�I��{�I��%�b}�wٴ�K��{�߯#��MU7�����bX��}�iȖ%�bvg�q7ı,N���r%�bX���lMı,K��_i�f��u���֍�"X�%�ٞ���Kı;��iȖ%�bw�ͱ7ı,N����K�q����ww}����~Y�.Xš����lvwi�/`H��U�$��}oGe[��Ʉ���;4�J�Մ��~oq���������9ı,N�ٶ&�X�%��w�6��bX�'r�ى��%�bw>��\!�j�3Y.f�iȖ%�bw�ޡq,K���ND�,K�}���Kı;��iȖ%�`��2��5u,��Fj�P���%�bw���"X�%�ܾ�bn%�@!bX��wٴ�Kı;�oP���%�b{��2�֥�WY5�2�Ѵ�Kı;���Mı,K���6��bX�'}��7İ?�*���*�E����@v'��~6��bX�'�~ײܚ�Y��E֋�k17ı,N���r%�bX����D�Kı;���ӑ,K��_{17ı,NwGOkV]fkdѣ:��\	�FpA�z���]ś8��6��vK��޾_>(��P���g������ŉ�{z�Mı,K��m9ı,N����*��2%�b{?{�m9����oq������T��ݽۉbX�'}�p�r%�bX���f&�X�%���}�ND�,K�����bX�%;�}�W5L˫�fk4m9ı,N���q,K��{�ͧ"X�%��{z�Mı,K��m���7���{�S���J�Մ��%�X's��m9ı,N���"n%�bX��}�iȖ%�bw/����bX�'s����֭˙��5�ND�,K�����bX��>���O�X�%�쿿f&�X�%���}�ND�,K�08�D���P1��2������G01�[j�&�9��٩�ېؖ1Ί]�v�v�\�K5sӍ�?��o�ó�#vl��ձ��.�ݮ�]k	<����aJ�*V��h�v���֘��b�(s&��\s�v^�����u{��]��[\��4�z��i�Ms�r^Y�HK!1v��z F����d�,t�|�z$�S$X�d،9�q�vp&�C�ݸ�9��f!q��.����lAŮ4�f��jN:�jC�5�t-�˞ٻo��wa٪yXxb���ݽ߻�oq���~�߸m9ı,N���q,K��{�͇d�bX�'}��7ı,Ow��\�ZԸj�&�F[�6��bX�'r�ى�1ș��~���r%�bX���z�Mı,K��m9�q�����}AѦv��*_w��"X�'s��m9ı,N���"n%�bX��}�iȖ%�bw/����oq���~�ߪ=qT�sv�����ı;�oP���%�bw���"X�%�ܾ�bn%�`PI"w=�g�w���oq���ב���
���"n%�bX��}�iȖ%�bw/����bX�'s��m9ı,N��ЈXB�����3XUu�R*��EgGX.�Y�{*�Ğ�r:М{�i�<��y+��)�w������ow����Mı,K���6��bX�'}��7ı,N����Kı;����:V��%/����oq�߯��fӐ�2	����C�D�?w{�"n%�bX����6��bX�'r�ى��%�bw>��\!�j�Y�&�Y��Kı;�oP���%�bw���"X�%�ܾ�bn%�bX��wٴ�Kİ}�����M�L�ګ����$)8J�O�|��,K��_߳q,K��{�ͧ"X�%��{z�Mı,K�wܚ�5��]f�h�捧"X�%�ܾ�bn%�bX~U����{�m9ı,O~��B&�X�%��w�6��b]�7{���?vuR�ix�
ጦ��DՎ�����7n[3��6�*�!ʹ�&��Z�bn%�bX��wٴ�Kı=�d����%�bw���"X�%���bn%�bX����[���kY�Y�E���r%�bX��zT�?*�r&D�=�߸m9ı,O�}�17ı,N���r%�bX���.{f�\�ˬ�\ɩSq,K���ND�,K�{���Kȇ�+��� 8	�Q,Mg�s6��bX�'�k'�Sq,Kħ}�/�˭ar��Y��ND�,K�{���Kı;��iȖ%�b{���Sq,K���ND�,K�|f{Y�k35���.����bX�'s��m9ı,OwY=*n%�bX��}�iȖ%�b{/}���bX�'=5�뫬�ֲd��ܾ��0\:ï5�l�u�W31�t$ogۭq~{��/˟�;E<�ݖ=ߛ�ou�b{���Sq,K���ND�,K�{���Kı;��iȖ<oq��~�Xƛ����d�,N����? 	��,O�}�17ı,Og�~ͧ"X�%���_J���@ʙ���~���Y�sR���nh�r%�bX����bn%�bX��wٴ�Kı=���Sq,K���ND�,K�w^�LԚ�d�.�]kY���%��U�'��߳iȖ%�b~���bn%�bX��}�iȖ%��ĊFQ ���@�"ow��Mı,K=߿~��p��R�K������7���'���bn%�bX��}�iȖ%�b{/}���bX�'s��m9ı.����wi6z�g:�����Q�m�zvѶ����mO�jd��S�OEp�9��.�&�X�%��w�6��bX�'��ى��%�bw=�fӑ,K��^�LMı,K�����.��˫�fk4m9ı,Oe�p�*�"�2%����ٴ�Kı?e��17ı,N����Kı=��?az��%/����oq�߯�߮ӑ,K��^�LMı,K��m9ı,Oe�q,K��}��à������w���oq��S��17ı,N����Kı=���Mı,
 �D�{�ͧ"X�%�￿y_�+'��%�w��7�����m9ı,Oe�q,K��{�ͧ"X�%�콾���bX�&*��C]��fJB��E�fY�2k+�l��f�얄��l�MָV�'k<
���p��r�v`���&,v..�<&����s:T��x��,�s��+a�m[n���1ڹ����N�]�!*�����m����kk]!p�uur�ɛge/5�`���ջls\�gu�Cdi2&6��l��8��-6Jf�7eE����H焳�2̹3'������z�w�ǻ����/��Ѻ.&fmvM\a�E�q��4l�96�'��h�ܐ3izM\5s5sE�4m=ı,O쿿�q,K��{�ͧ"X�%�콾���bX�'}�p�r%�bX����Zf��k$�u��Z�Mı,K���6��bX�'���bn%�bX��}�iȖ%�b{/}���DF%�bs���p��ZIK������7���{��o�&�X�%��w�6��c�"�ș�_~�Mı,K��߳iȖ%��{�߯#��l*��}�7���%��w�6��bX�'��ى��%�bw=�fӑ,K��^�LMı,K�����.k	�WZ��h�r%�bX���f&�X�%��R>��~ͧ�,K�������Kı;���ӛ�oq����۾�څ���qXz�q�g�佛��y:�s�Q�]j��G�)�ww:yhXCV���{��7�����}�ND�,K�{}17ı,N����Kı=���Mı,K��L�j�չ�L�35�ND�,K�{}17���,F"��M��uQ,N��p�r%�bX���f&�X�%���}�ND�,K;�~�VN1-�%�w��7���'}�p�r%�bX���f&�X�F%���}�ND�,K�{}5��E=��)��}������=�7|����3*dK���i72�D̩�{�ͧ�Tș�2%���&�fTș�Z����L*!UL*!0y�2����-]h�ֵ�&�fTș�;�wٴ��2�C�u���WIș�2&eO~��Tș�2&eﵭ&�fTș�������۾�n��n]��F��\j�3�rdn)bۊ�{P�՗��l><�ݬ�7#�i5�t[��'{S"fTș�����q3*dLʝ�}���2�D̽�����72�D̩�{�ͧ�Tș�2<}�G���U�(��7�Os�ٕ;���i���GQ5��2�����Lʙ2���߳i��2&eL��{}���or��{��=���?[��d�Y��}�L��S"f^�Z�n&eL��S��}�O����N�]�!#� B2B!��(,X�WjԌN�"k��V�8��x�!4X�,��	�)���,.1�`�����1���\&)�)�\c��1��������B$`��P�K�\HD`5aV�qFY0��' ޘYII�f�HB�Ȱ�2	�I��LP���AH@��bňA�	$HHH��b�8j���p�D>XYH��"�01M0����B!,����$� ��i����1H���`�D�FF`I$E� �E�$B���!��h��U��b���k]��mf((��8��J"���ʊiV
�H��D̿_�t���5��2��{����tD�Mj���S���P�	U{�or��E kU=����O���3*dL���WI�T�Mj�D̩������:Z�j&e��kI���2&eOk�3��.M[��Jf�K�o8��L��S"f__ںM��j��fT��~��}�L�Pa�T�L���֓q3*dLʞ��~͟��{SQ3*dO�Q?�]\��q��[:�/�>u �|4%[�Qۖ�X�Gg���]�f��˖�n�(����MD̩���O���3*d:	j�����Lʙ2���߳i��2~��T�L���WI���2<����r�=B�p�=����w�ʙ2�����?GZ����=����O����j��f__ںM�̩�3*{��|l����!@�k*dO�?w����Xv���m}�~��qZ��߿�i��2&eL�@:������Lʙ2��{����d��05����}�Z�n&eL��S����\4k5��]f]~P	������3*dL���WI�~c�T�Lʞ���O���3*d�(@֯�kZND̩�*�����W�(b�]����f���kU2%���h��L���f�\ֵ��Lʙ2� 	����i��ș�2B9=�1?!�ı=���6��bXL����MD�,o�/���ݛUl�HQem�x^r��孶��p7Z;d�T�擣�����vg���U69��K�jI.w���$��dԒ]{��~~ ߼�a`s	@�_ ��W��I%zɩ$�����$�W���K�ݎ�&�б�#���K�dԒ]z��ߐ��u�RIs�_��%_\m��☐��ӒjI.�g��$�u�RIs�_��$��ɩ$����"yq9�'3��K�ɩ$�ޯ� >�zh~�W��7$�{�����_�)u��p֣���b��l6���g��m���86���kV��<t�)�nk-`ֲ���l�s��>�lD��:��gI�����ڕ�6N�9�/N�t��X�Ia����S���#��I��q^�s׵n��g�`w<\�=R7eC:vx�0h.z�5�t�2]Y�΃��$��8�]�/�������;%�Sӻ<0�lnvy��ֶ�n� M��w}����������>��<=i�=U�l�&^p���`��q]�u:�[\A�.8�4�T�6�I�K�Wwl?�S�[�Հ�=|���ذ?g�%��hw���ɑ�H�jbN=�2�=x�عB��@���?(�S_������?<Q���n&ړ}������, ���$�� �V�3���@2�����X��F㙾��䃭��*����Vhz�h�q�q&8�qI4W���Vhz�h��hnGH�L�"?���	3=�Bv;|�W��<&n��.K[���BƏ3�sV�ƒ�8� {�zhz�h׬��ߐU��U�~7"Ć⍵&��^,���B��P�.�y����� �f�1#�}�n<��q9�'3@;ϯ �z�J&N�=x�ذ��L�D�E1�&���zo+4�w4��h��q��#��F�Ĝzl��	ex�=e��*`~�&~N�cV�l�8�o,�ŝ��&�r�V�y-uv�4�]B5r3�\*���	ex�=e��*`ͼ�2[�X�n$ԍ�3@>�f���zo+4�w4�q��Q5"MIx��X �˼5%��/�%��P�S@��@99�ٹ$����$���{Z�i"@�= ���^����4W��9}�ӣ��X�n9Rh���9(��}�sϫ �w�?�����2c�<&x0�(2ym����[�&�u\�+)�ms����t,����z��	�T�-�y�,�ۭ�p���(�8��9}k�yY�}z�h׬�?}ey29	k{5.Lٷ���`��o�Z�X����N5MI�}z�h�]�?7XDB�P�Oi� /�T�f'jF㙠^�@���@��@��������Q9��ȜGV'X�����\ ۥ	��۞(�:Ν�R��2A�b���I�r�נUy٠}z�h׬�9}�݉<#Q��0R&���������So�4��%#���4�]� ���/�zW���tmǉE���n���/0&����b������kmc�%#DQG�/�zW��� |��p�J"~ID}S�A��b����1�\�m�V�z/u�.D�v��vފ�
b&2�_+���-�9��2;�/m,w;1���X=�� ����)u�Aɉ�p�;-�&�9�'z�����K�w\�x��\;0L֝���\�$�u�r�:���h��M���x[AL��ևZ�w-��[7�mk�$�����$�\9���#�A��kp��Rd˗Y��EC|6g5%�f��M3�\Davm�\��lvz�{�qػ�6�6Q�hW�vt�pm��$�����t����>�q`�]�!B_��u`먚�.��$.\�Iw0=ex�=e��Z�^vh}n:�18`�RG� ����Z�lW���`��.[��K�o.L	��0&ȯ0=ex�������nĞ��D��z/��������T���S{/-�s��鹤sYQ�v�e��N'n��LR�{v˻Bս���\�������m�������T���So����Vr\-��Z��f�nhܓ���7�
qC���P(@ 8�H/�A�4_�O����3rO_w=��>�}�`r���9R4EG#�9}k�9nӼ9(�����XӽՀ~����V�I#jbn=����>�w4��Cٟ�������/������q���`K+�����6ʘ}������r�+Q�v�iO`pl>�p�)k�
;iqk���S��3���aJ����}*`M���Ey�,���d8�F�q5z+��3�?�"�W���_�0?zW�E%{ua�x(�	�� ߶]�=x�H�
!)�n�h���/�5c�X��Q��`z���Ҽ`M��=6��VF�<��Ȥē��~�����z�r�@��s@�e��"I29N��#�0�Er-X����nN!�r��;O=u�A7k�G"�s4W�����^����h�v��LRH�S7W&=6�Y^0?zW�	�T���t���8�M�&�׮���^0&�S �m���W�nj�K{�r�`~��l��I6���̘�G�����T8��o{6�q��x�Ym�	&h�W�TYy�,����*�E��]٨nAn^�6�˝�d�oi�9�%VoO�����\�ƣ��I���@�= ���:��l�l��7��A��f�Q7&�׮��#޾��*���z��K���ȤL��I9��w4W����l^�����˭m�r%$v������eL�y�,����?|�M����26�$���٠k׋ �׋ �z� ��jP$B>�#�X@�"H�$``B�?
ͤD��.�*Av��&��``�!�<��`�M��0��@d$-*�Pd#��`S �:�`�Z�(�V�C�$a�$f���c�0��'`m@�#
��1�H@�`,Z��ma��<�
�V
�?QC��GC�X�	\F<:R`YX1�# �!4��#D`�+0��%mIJ�}��8�UKNy����4��ФT�� ~��{��v�����]��VWj����tp3�<n����jIΒ3�m��^��\$m��6�oH|Z�(�d��˘�M�@vá'^G&ӥ�j]fZVjicQ�p�د�6��H�cq��!�y��#u�/p����lEYN-���xA�8�s���J���]�#��;�M�̤����,����pkR4��I�@N��%������*#�B�J�6���2V��i��n�;��p���e�7))���v8�L�eݭ�L5NwC��X��v�5����{U;+����H��]<���M�ʹ`��&�m���/J��ͻb."�sÀ���<
�6�`@
�`��Q�ԤFV�ۍS+dp��"�4���R�|�4�����v�[�cL�ɚ�
��s�U��-(�#jrX݋i]�H�������{gG�v��;v�q�̨���vԡǭ���m��0�#�wU�RA'���"m��6n����/Hլ��-ޤ��
|��Ϝ�C��mn��{gd.L�!���Xj��jE�#�9�^;DN�]o!�ˠ<H�����	G �b�d\��v%S�ȸn�j ��&�s1�n�� ��l���h��؊����@�2C�E���2�]��ѺƄc�b2����h�-)�֌s8��/\�;�팆�Hl�k�:�h���f���$�FK	w0h���h%z�t��ێ\t� ��M���t�b��k�81���`]gK��Ws����̻l��H7`#D�u�{j\�S*����єXڼ�Kl��p�;5u:�[MOix�M��A�T�8x#19�r�g����G��'�p�e�2�KPRp+ŵ�p-52QJ=�m���s99ɧ���P�
[)�`�h�RB�����)��Z�e2e�Fݩܷk�w��*�7&�]�+�x�&��]�pdj�z�.s�JA��H<�q�5<���V���m�-]@{I��ʭZ���s�Ij�2�&�f\�˚֍(�:!�? �M~T�&"lxAM�? 
|����ɐ�Y$�MXb�^`9��apQjݷ-J&������;�K�6���{�]�(�9Ee��E{q��$��n��{bi���ۖ�KK:��Q8�yJNXx^	Zu�����I��%�\@�d�݇�:�.K�hҏBY�\5�yw6���-�����t�n˶�M�n�ӻ�ܒ�@B�1qZ����HH�֔�úxK�tTGe;uX�ƻ���>;w�qm�N�t�gV�&{�SX�GnN��m�=lu,]g�p��ʤ��K���J�7֦���>���N&ԑ�3@�빻��I�T�=�y�,���ś�s�m�	&h�W���O�W�ۚ�ۚ���v$�MB,�#�@?u�@�W�I^0&�So�-����f��v�sY^0'����m�0�٠~��TcyY1G�5���ܻ /Q7�Cv������ݔL�4�Wa�gM�H���s4+���l�:���>V���"JF��M9�/wٽ8��$����{��s�܆�X�Y�
���t�R�7wsE�]Uu�wu�=x��P�gu��6_W�^u��H��j9ܚ^���X��X�D%3�w^ 3�Mu��łmIs4+���l�:���?}��G#�!��q
��眣8rNด烛<EL�{]���V%g��m�	&h�W���@��(Q�G��b�5ӥ5�SW3Se�w.L�����$�l���33�*�z0nE�IȠ����X�X5�D%
RID*ݺ��٠^�[s�82'1$�h{3�?��߳@���@?[f�b�w +մ�Ȓ��(�Nf���P�����wM�^0$�� ���������{j����+,�Ϧ�;ZL՗��\絥���aY1I"b�!'�~���]������z�Xۣ�	���@�W�	%x��eL���-�W�K���˗cI^0&�S.bG�٠u빠���x��n(K��l�u��w�k׋�$���Y�?���Kl�4μNƜI�$	90��`K+���`M���d���;WlN�[Z�M�� ��uWPN���\Zp�նY��ݖy)ة�E��� ��,w^,e릡G��n��.6�$pdNbI��;��o�3�DL�y�`��x�x��몙Ue�F��M9�+���l�:���;��h�}Sl��D��JG�����W�	%x��T������%��ʪ������ ��ŀy(M$�����t�z��n�Q*!G�"��S�?��n^StgiSkWV6�dH�,��{r�dke�%����/&��k���\u�ҩ�rnv��ک0˞���:܋f�֞:��]���@6��^�A<�e��˞::G��v�{Zs����:�\#'*�P�t�N���z�u�����y�c������B�����ۇ�[a��]�;n��v;K<�m�dp�z]�:��]:3Z���� ]*��2�ڛf�B�8\'(Ώ-��=�3��8�YV9_{	zu�O+<��aJ�������ŀl��`���%�7�b��T�dl�"m�	&h��￿����M}~x��W�	jUr���]u��w�|���TDD��X�����ƬǊE$�PNM��s@��o�L���ι�v;������W�	��0��`z�������nϾݮ�]�Ju�$���E�K��۷Cu�g�a݋yj;L�ͣW&��V���Z��o0=ey?�����w4�>�6�I	#���8���kJ#����x�`[ŀl�u��D)���~pm��nM��s@�빠r�^�~�� �q�^<N,d��Z�7u��6^��ͻ��I(�Ͽf�[�kё���$��r�^��BJ~����ذ�x�mM�����9��F�]Wc��N��>�mc��L�N�K[lu��ޫ����u��6�����0%��I^0&�So�-��7�� �ݨ����W�	%x��eL��h�\i�O$��$�h��`/]a�D%��J$���׀=׹�}]���cDQ&������n�z�`z"����>�|E�p�E�R= �m�^��w]������ɉDB(����&9�}���X;�5�PѺZV��E/"��q.�i�Lv$��ݢ]�	ex��W�	�T�?[f�u�ݏ9&�$q��;��`M�����	ex�$���9#��$��r�^�~���]�����>x��Q2�"8�=���g����X�XBJ1B�/��g����r���1�<`���ɠu��I^0&�S �m�ٟ�N3t���q�Zu�k�^��'�m�`��@�Ÿ��gM��N�:2-��+3cKv��-�<`M�����	ex���Rk"$ƈ�M9�+���l�:���;��h�}Rc��R8��%#�ͻ�5�Ň(S-�ŀ9�Հ=U	*.�Ē\��K��,�J���z��4���y&8cm�G˱�$�l��~��Y^07%ު���]�J�������-@6.:�1OZUa�v���7mpɣ�u�����;�l:[l/���������W�ܞ�G=j޺qr˖��؅@��1�:�1�	˱��r�V�C]�n�cf��i䧋',E��+�2t���o��V؋�i�̓5�ʸ�%��>k��gj����D ,PcmͷF����j���5�Ѭ˚-�"�O k�9�jd�).KC��*D�粫��ҎY���q�.�a뵔�)�K��X�]�m�?�~L�����$�
,Ԫn.ӎ�wr`����W�	%x��z��ݍY����LNM�W�	%x��eL���N���Ջ�r]���`I+��*`������د��f����mc�%&4Ei��6^��ͻ�5�ŀn�ŀr���۾��v!�գ\�q�vn�\�`����Y�s��l�ĥ�hNc��hܐ��ݻ������`K+���`M���Xۣ�cm8�Crhz�l���?���%+�����[�*���Gw.]�	%x��eL��hz�hu�\d��"m�	&hl��~��Y^0$��AE��B���b]�w&���	ex��W�+���|XҌ�?�����z�T��n4�V���b�AM';�t�yn.yj^J���r6''�/��4+ν	$���w^��*��4���&�еv0$��m�0��`K+����X�&4Ei��9^�@?[�nS�0X���=�`��@��K\RMU�5!�� �]D�7��BS���0i�e!A;t�B6���C�U�Z!eB![D ��a	�� *d�0b�B���	@�  G�ƪF tN9Z�20��F!��dZ!�p"C"�O���(�A���ӈ ��1��B(�'��� �Ev���)�U��Z��_��(P�?�`u��?}Z�TƢq�$�)�~���]������z�XۣrcM8�Crh��$�l��~�� ��j��AR��z5�6��/ ��h:˹^�qsأ��=v��B�g��lەuL��m���^0&�S �m���`\Ur;��DۊL�9^�@?[f�׮���s@�<M�8��6�(��ջ�׋��IL���ϫ ��SVc��x��Iɠ[�s@��s@��z3��f6��h��Ɯ��7�b�]�%x��eL��`[.�����G�	p$ȁ*��0u�s,ط'[Y��0��k�����*smucPQ����yz���٠[�s@��s@��7�cQ8�D��@/���^0,���0?Y�	.wf�.\j]�ex��W��T�/�� kj�͕eت�����X�����<�|��l�-빠|��댓�M��4
�W��f�o]��=��f�_��Pb�HTM}�91Ԗ)��3��a�l#P�.7d�����s�G9$�棻]���������Ёv;-�$w]vs�����u�q�ۺ=����V�jn�6�ƜWUC�f�:-�W��Hx�X�M���Ѽ��:N�:�ͶY���i/7k1��'�/cF�ݠ0�]GM����p��/;[c!x�)�ͱ�Z��Gv�;-����������=�w��F���\��ڤ$͒yEצ6ӝ�
���u����ta@���c�Cjb�? {�f�o]�޻�W��9}�՘�9 q�j]�ex��W��T�-���\m�F�Ɠ��[�s@�ʘ���^0$V�[�����m9�W��z�޻��{�߳@�����1��q�"JG����s���ϱ`^��>M�-`]HR�X�]n�<�%p��ݮI��i�m�;E�/[�9ۃ�bm����@���l�l��[/0	n$^���32�]k4nI�w�7�� m �p��P�_%wB�/���Հ�u����9Uq�&1Ȓ��3@��x ޻Ô�s�Xs�XҶ��:*,q4�q�}�o��{�ۚwL�Uw��9w��Lx�P@ԌMɠ[+���`]��l���2u�B��GJUPE��NM�7-m�����{\<uA<O13�ړrG�Wϟ9[�ڥ�܃w�ϱ`^����(�!�� �w�kɒcPQ�������f�o]�޻����ď��ɼs��䒦f������ŅB�(�""��(��G��>�����rO�����?^���9&&ڎ	I4z�h�ŀ9z���3����*��n�ب�WsWV����9(��}_�;���o]������RRA7$h�x9¥���N�s�F3�W�K����.�-Cʑ����"�f�U��޳@�^/G�%P{��X���5^��U\��jn���w��Q2w>ŀw>ŀ9}^���Ƭǉ�4��nM޻�z�a�B���}X����mUU��wuD�Z�����
"{�~XO>�	=��[���c ����d�f��;Sk		��F�s4
�Z�:(S����� ޼X�^����ɰ�Gggipp�R�C��Qv��(����[�����w���|��fZ��\� }�����l�l����*�ʫ�Uud�]��ŝ��9�ŀt����w�	DD�>�Tu̙!���)���s@��z~�h���>U\j�G�r&���4=��!)��Հ�׀7�(J"y���.���E�67G�_���w>����,��X$�BoGUD��3	���k��Ų�J-t6à�������;Fۑ��1v�������[P\�6ˤ=�}�d�V�Wpb���[vV�4�m�I���v#@�/�"<�� #A��	��Nݧu�ݖv�p�n`ŭ��qy4�6f#�7���=�]�nl㷍!��Қlr����<��{sю�7Cqn�L椀a?�H�э2�����q���v%!c��r��6�|��7=u��kls6�甭�Ѣ��w��5�'Ғ9(���ۚW����@����<$��9�*��=׋?�%
=	%
����X��^ ޼Y�DL��j�U���Sd�UMv0>߯ɀ_[�ex��W��V���q�"JG�����Ľ��{ϱ`�Ł�(���Հ}��������ˍ����W�ex��eL�w�y(��\��&�UwSW%+�����5�p�:tu���c�ܙ���)^})�i�K�`�����|��ؤ�m<�H�|�����U���w����ذ=<�z�5urM��uk r��jJ��DDE��P`?ٗ�6�,�x���ӭ\�U]QUa��0��s�^0-���0"���1�p�RA�&�����}�4z�s@��zK޾�{���<$���ؖ����`]��l���W�^�4e�LN��R2b��P�:y{Z��o�KuD��.a݋x�����!͵ՍAF�s?������w4z�h�v���$qI"JG����L�ϱ`ϱ`^��S'��*j��U�*�n������,�x���Ȅ���(HI$	/��9�������Rc�1��8�h{?��}�4/>� o]�z%=Ͽ,�O*��&jl�&�컳 r�������ذzS@��D�rcSfH�c$$��u�0�V:�J����:��i��II����}%�UuD��7W_ {���׋ om�W��9}�՘�A) ۓ@��,�Q2w;� ��Հ���M�ZFĤ�ә�[ҚW�����_M޾��;�T��0�&EjCC�z��`s��׋ �I)J҄#bhE0 8��7�޻�&��y�R�WuswsWw37u��Т!/{���{�~0/]`���w$�]֜����^��(wTk�ύx�ۉ�E/9��W*Lqƛ��ڎ	I4z�h� r��G�����UEtݪ�Q5se]Z��fyD��ϫ ;�^ ޼Y�""ds�ʧ����W35WEݘO>� o]��{�b�;��9�QT�l�WtUXM���DL�>���,��`y(��}X�j��R��d�3}�K��l�Σ�0e�IŨl$"F0�@��bE B"� $ H���@�HT$X� ��� �$XH�)��"��A��@+ ���@���S"��!	��T�H1f�6��8�+�)ɂx#%�+��H��%Sf�
�#�T�	�BGJ�,H0!����$A�BD��XJ%+H�<�܌�I�!�3z��pX�4FH2$!�b; EO��ĄB����F1H*�o���<�����	# � �����a��� ��QF5+YA�0|0d$��v��m��������V�\��J�UT��R�����2j�K�my����]u/]N�Ka��tU8��m���랂���P����ŕ5�B�2�U5idkj�����V�OhNyu����
��Wu���y�S��Y9�Hq�V��1��l��������!^�7B���9��m(lN�8k�ư�m؍n�s��`9�����m�ǥ택h˟f��ۋk��g�y�:��Wu.Sd�Wn΀�I��Ʋ�Ъq�e�Ց����Md�b������U:89���{c�5]�;Ɖ�oC��w����4�ƹ��7M{Y�#�����v�ƨ|�`k0�9�M�!�^�ݐ�|U�ۊ{3��ˇE�f�\�`N���K*��R�q��3�U�\q��N�ۢ0��n���kY�1
P2���]�qnN�v�v�G%��X8�[ngJ����B˸ݶ���Ƒ��2g�i���iհR7]�v�R{2�N�sE���j�_C��Y���H�[u����<��Ů��M��h�9#����@��d�H�ܫsv�.���FOj��v�7�/O.Yぞ�pU*;g�.d��n�I�܈�vr��n.F��}g���O�Ԯ��@��z�oA=���Ƴe�m�Lq�L�����:�v���c��\�Y��wkT9�����u�ۃ���X�������6E�!#�6��L�:�X$i`�F���I���\@�O�#�$-#�Z��#Z�N�I*w0��9X�v�	�V%�����l�*�iUV5nOj6=��}�u�wf��$��Fb�8�+ŭ����)�M���s��1���2\�^�5uj�e�:�*����N66Fj�<���]�ID�*���gi5N��ػ,�wBm<�8�w`��+�6��ȁ��jZ�FZ�;�lқM��9��9�ャ�m�����d��Qp��M�0��N��-K�[�ئ��t��^Rgge4�H�wC���QY펻)�V��!9�(������"C�Sʠq ث�v�.y�)�S��lP؈��'�>�aջ��1�����ܑ��-�:���4�5�^t��2�x��\�y��un:�lXS��:�q�g�����y���<��$��8�\�� s��\�����r������c\]��%E�Ւ�[��	����|m�:�yMt����3�\lJm���g��[��g�m��J]s���|�.{>9gD����8�u���狊���������s�zR�b��\Q�VY��n�s����k��N�$"�������6%&6��[<h]u�뾄��!�� 循�Uh�s"���!�Uz� ���-빠_�������w��_��y���j���_��l�Σ�0?YZԪʫ�UT�Y3wx�(��}�`����u�ВIL�>� }ʨ���V*�9��)�Uz� ���-빠����#���xF���L�*vp�Nl
/0�,���x:)�y��l�������>\��Ȓn2H~���@-�4z�h���Wݍ:"��(����[�������(�Y���� ��|`^��6~�R�R����SwE�]��ŀ7��:"!L������}m���F���ә��^�|h<�����yBS����5�驕V�$Ƞ�mHh^�@��b�{�����{�4��c��&dɋre�q�����=��jx�śd8��J���'�d�)"rD��@/��޻��yDB���}A��z��{*j�ʪ������������`M��l�}������I���93@���'o}��И.$���-Q��v����ŀl�j�ک��W35WEݘ�G���ެ ��׀|�ŀ;Қ+�Ӡ�'7&	��ޱ��k�����-L�M�.�^��v��s*�غ]����S*1)���T�m>��`V��y�@�YZ��~�|�7��g[�/�ou���75jiF�I�nf�{�7ؑU���{��}m�������]�i2d�&D�jA�v��`���׌'Q���Tx�H�&����٠}m��=���rm��*b�l��{����؛pi�6�pJI�}m���f��� 7����Z	��S��l�d�g�=܋�T�b��G7=�;it��Ov�@i<l�I��q���z�.���f���s@�UƬbr8Q5WEݘηY���w>�{�oJh�cN��AǍɂn= �]��Ň�{��t���6~�R�S$����4z�h���U��=�{��@�zyF�'���Rbi���f �� o]��ŀTF�y{�����v:qp]�^�6�+۬�j��Ϲ����s�y����e�F��u�^{Dh�e�=���t8�b5�ۃYP����������&Z��-�鴪F��p��/(����ڹ	4��N��vt��h��\�lL�W[<I tn� ���C��ʚ�ҔS��v������dv5�4��U���i���v�EFEN�*���������w��x}�!ن�Z遍]�Lr%��=ۭ����8lzsك�F�ȳ@�k��T6�������������9�� ݮ��RD�q��ٿ����z�s@��ƁU����ى�=�pM�rh���{�4���*�P�o0I�K��Vp}���dt`Uo��_���w4�W��I&Bj���0/]`�����s�X��?p�s��jcpQ�5:�93��v�z��	\i��v�U4��75v�����w�7� �m��
=
!}A��z��ʧ֪�mYE���SWxz�g�E���{���n��w�	D)�{���M"�nd��55k �w���eL�y�l���Գ�*�\�7ww5f(Q
z��`s��빠[Қ�;cx�5!$M�%#��w�rJ!w>�������7���1��m<s��FR���%�s��s8�]ۛI��et<a���z6����iI����׋ {����\�D/�o�4�����i8�㙠^�M�L�<��������Q
#�DB��|��t*��T]U�wf��z�����ب�h�׻훒{�צ䞟�US��e]*��MU�BP�]s��;�b�5��OW>�εS֪��l�\����� ޼X�(I��?���@�z��gJ���D�rH'Y��v�`��E�lTՌ���	�y���M�e���(���ә�u�M������""�ϱ`ϲ�Z�Wj扺���0����S#�}X�ذ{l�Q�"�n��t��we��U�3wXO�Հk׋ ׶�e���܍�ܓ�G0R=fg�����f�}g�䞾�rpE4
��\�_���덖)2CN88�hz3 �J!us���}Xz�`}M�g�՜5�h�G$AR�Ө^�s�\�W�ԜcF�-C��꣝,� ��e��x�(J?H>w���~C�<nO�8�W��;���5� ���B�Q�	(�:_*�Z��PfD�q���ۚ^��?Wj�9^�@�ʣs����s49B��_<� ���p���=	%-���z�bo$&DҎ8�4�ڴ��/%
u��_��ŀk�f���۽����w�%' �]n�@��#n
,�w:z3�ض��9l�Ƨ��V^�v�x�02gm]�p<�y��>Gnܘ7IIm��xM�u�ָ��w�c)�I���U�3�&P���G&n9�9����]��!3�f,��%�� r�l�6ۣu�ܛ�8=��M�nۢt�Ÿ���G<��v#�ɘعpg#�Vy���Y̐�3Y�˙\ѭh��#�u�p��n�x�P�n�{<��˳�� ��q�'fQ���Y���t�by�U��c@s�� �׋ ׶�DB�_�>�����*���u7V���w^,�B�#�|`uwN���zBQ2�Ur��!�'s4�<h��h�W�wu��*��3��#q�C@���6^��7u���K�`��o�xAǒI�Ӌ@�z����ץ4�ڴ��KM%��Q���[E��>|�q��#�umӀup�+/Z]�m�g�7\����{�ٍ��D�q����息m��M��/�y�`�}75h�U�[.�\��rN����ñ`*mE�Q�	G���ϧ ����7u��DDB�;��y ӄQ(��@���Z+ΰ�D)��b�;� ��nn�Z����Ի�R�`M����`K:�?����^J+}����~�j�j����]Z&��x�BI��?�Wt��]���?v.�t�����qm�U�8�^nNݧ{���)^��k�&�X?�{�ϟ9_�6m�3fl�����V� ���J��n�R�7wJ���.��?:ns�
�%T}��;�ذ��0?j��%"ʺWwqSW8 ��x�XlG�""�"P2�� ��J%�� A�jڶ�FYZ��$�$#
U�"1c�#�Qba�D�`<�bA��B��5��!57���h���H!,E`�@�u4�B�k�T!S��F!����	��� @MnI|y�)�#!2!�E��tSb8��U>P�C�(�'�(���:A^�'�*	~�{[��}�����w�]Z���(���*n��B������� �_O�~�ՠ�@�ʢs��L�V����?�ـz���g�? y��4��ƌ�	����ډ*$��W�.Ἤv�-�C�:w�Ծ�K���4��Gn��Z~�4�����=�x�;��Ƥq�ܑ7s��w�n�ŀ?�ـ~t��(��G޳�M��mH��h�nh��`~��`�� ����r�7R���`rQ	Ok�0��� ���� �
��(DLDl%��w� s��K���*.�����u�_K�	%x���F���{������b�ݧtQ�ի��dÏo�\�j���5/d��Śp�5D�~�����}�o��G�I�7 ����-빠_�S@��z��4���HƤ��w3�!L����:y�`�]�7nnj��qD��9���4
�W���1#�}4z�s@��u��"Bcq(�ف���S�ϫ ;_^ ޼XIOk�s�Qc�Ԏ8�s�����=��}�~�������9�.;q�	����	�\�m�]�qd��9�"1g��[�WZ*z�vБ�rm;b�n�p�Z�/��}۞ڶА���؎�;uG<@(��c���!����:��v v�:�:)9hy��v�[sDݩ�"^M��Vk�m����<�u�� ���r|�g=V7ù�n�3c*�vړ��mN�=�m�kka[�3�����<���S�%���)X �����RtV�7tZE�LF�u���O��&�L�6�JI>����s@�t��U����h[��G��N89V���0/]`�]����/B�6}>U>���*���.��:}ެ k�<�e��Xk�0��US��ʫ�$��q��/u��/��4�Jh�W�Z��N�@9ԓ@���л^q��}X ��x����%6���Voa���3q�.f�k��c�\ږf��=\�t���b�٤�n���m���}��T�/����`~���gh�4fj�f�Y���v����R#��+��}xk�X�m��SwR�a$Q�ۘ��@�z��]�=����_Y�@���@�zV&�RL���Ĥ�^�X��`/]`t(Q.��`����<��qȣ��u�M������~�>�^�X �|N�)M�g�']�v]ʏ�Wa!eIe��8��Y���=<�%s��akU�m�O��_�6^��5����;� s�T�!g,\����Ɂ6ʘ��,�h�W������H���6�x�RD���ϱ`�ك�����IU9�u�r���eQ9����G1��h{%	K�`y�`/]`y%/�~Zz�bo&L����7���	�T��W�	gQ��,��a���ݚ��u�sÒ3���K�f�x�x�śd�1�cd��{��w|�_$u�L��%?�~�&��`K:�	�T��ekuU�wj����wX�x��D(Jd|��>�e���A�*��)]X�f����� ����XyB�2�=޾��*��N�ԍ㉹	!�9z� �z� o^,�&"!B^K�P���
h�+������'���M4R�Uueݫ���e��D$���g�/��Uz���X8d�i�3qq��8P1t8;^�v*�[��ƻ�~�t��%���Lm���4�#��}��u�M����B���DG�>�V���nj�H��9�^��*�נr�^��^,�#�(UG>�eUD�L�MU+�}�`{d�{���w��R��]��Gnb�=����w4�)���������>�����9m)1)�d�Σ�L	�T����y���?y�y���]kjB���1i�mW.������e]�9�ݭ���p���mA�NQ�۱�U����:v�s��V5{k��͍y�i\�6���m�6�v2���9��ݷ`���nu�q6����h]��ۅ��sd2��1˒������+l�iJ�cM���];�z�-i�]�o}H�m��2l�tWu���֫���F{	��ś̞��ǣs���k�c9^�w�i�z]6�m����ww���Z<��q��3��<h}k�9^�@��s@���:cR7�&�;�`]���6ʘJ�,�?�3�#ˮ4�ģ�#�IǠU��^׋DB�Je�0���֪�ꊻW3S7w3Uu�Т#�B�w{�w��h}k�9^�@�h��F�#�-]�	gQ�w֦�*`z���������&�Z� �mq��dg��):�ѭڍӍ�`Gg�,.��w���o��^�sg��.\���>�0&�S�W�	d������&)"�$��z+��U
">P�(If3�`��l���?^��n(�1�1)��빠K:�	��0&�S ����.�j��n�`z!G�D*�w�K�� �}^��빠n4�X��RE	!�l��`J!G��Q���|�{�o����￷}ԑ:�r���itƕ���w��Na��ۖ��{quȤ�3�y���n�L	�T����Y�`M��@����lrdI�$I���]��DD%2>w� �V����l��U!Wu"��S3V�{l�6^��""�S0�t�����>X�	Dz!(J�t����;��X�yST��iGn�U���z��z�hzS@��li��FD�Ƥz��XD%	y(����|{������3�����l����F4��r#�Z������֬l����.ru���r�]MTݩ���5�ŀk�f���$�B���_= ��6ׇbqF���u�f�������^,�%�A�&����xE$P�^�z+���ġB�|� ���ڪi���Uweݫ���e�^�X��`}	B��PGJ#�P�~��ܓ����35�rdI�Cq�z�hzS@�z����ݝ*�b�&A���o$�ڃ� ^���u��}T�	t�qڜ�j�Y+#FD�$���Jh�W�r��$�~�|���.j���VU���.K��*`M����`K:������H�~�k�I�71��W���,�Σm�0?YZ�K����l��S7u��{�~X�|`^���DD)uϫ r��⬫W6Uզ����eL	�T��W����ػt@�Z��"+�ϒ,&@,Y1�A�H�1�+�]�t�*B���d~�����_�1Yq�A>X\�T�UA��M%�i%���+I�U���ڸ%�����F3� /6J��@��-M d ����B#$��*��0)!0��#�Ȋ�{���~?`�8m  �ڕ��w,	v�Ӕ�e��ũ8@����Uη]�W�e ;f�`��c�V�����J�T$A��n��z��% H	�����퓭��Ih�l��� :�+�n9z����H��d�eݡe�ظ�%�鑞�L�ħt�n���K8��]��1�1-�6���Umջ���Ƈ����y��.�]�ɵ�L
s��]\ٲ�l:�:��z�g���WN���-�]Om9;wYKbΌt=�ݸi��%kO%bq���cل��F�91s�,잰�94^k�z�u˻<��ƄB&�*��9�a#h�UʻUHt�뱞є�5!l�\��᱓v��)�B�w\UO;<�kEA�l�f�`Ǖ��=ne�$���+��N	W�]/c.k[�H���L�c5�#.uɑ*x4b��.��+���H�v��X�um.dX�H ���[Q���KjC�����б��᫦��٠;a�mq��n�-�kMu&�V�ٗof����δ����̼���ۣ�� ɍۚ]玦)�G:�AQ6IW��r��x�����#�5]�un'��u����1���Eʮt��K�{ֱ�*�&#�m��+mIk��q�K�Wb^�{�@bŸ۷%۲��³����k��9:fԎ#C���i�*c+h���9&e��Y�]ւ��ΰ���v�Y�]nh5����9�u�Q�o#�.��RM�9����-�Vs�Yk��s�sO5�[/c�Y��h:{Q���7#�I��ӝ�X�1:8d�[jɔr�b�;:v�B�ᶋ�]:�ژol��y�,jn��c��Y΋��ѧd��9�$��y5q����Rj��b�QCH��g;aq����f�4���x��3e��S���d��M���4��TL�i���ҫGD���7��;7N�ڌ�8�\��b��j�ϱP/��6�qL��{�����{ߛߞTC_�؉�h �O �
�����3�x���Ic u��N�\��yy�M�Ş�8����{���=�q��ɶD�!��b.óq^&��ll���v��j��ݗ��]�q�{S[��k#˛'�R�uf����෱��],�i!��us�mɥ�is��C$���㱡u�\��g<t�*�t��8I9��]@Q��z��*�ر]Db�:N%9۳h��K���["������w��w����:��;gk!��+�u� �ע8��v.s��츆�g,K�6��)5#17I$��W�^���xz�z!z"!G����"��rAH�n=���z�hzS@��{�����H���5#&D�Q�7�~x��ul��6ʘ��[1��K"sNf���_]�U��l�u��
"%��� �}�5J��*�w�.K��*`M����`K+��tɉ�xH��80��"w89�ֵN��\v%3*��bnw>��=_��{��7�y��F�C�܏�z��z�hz���3? ���@����n)$�A�0R=�;��f���`�E�A ~�! �����(����E��X��� �z�=��>W���x����G3@����9^�@�z��]� �q�����H����l�u�l�u�k׋�$�K��٠U�~C��$$�q��W�|���5�ŀl��`ID=k+�fX�0�?�� E�5��K��Y9�Ӏb��+/X4(��m��?�w���|�y����uu�w���`���6~n����}q���5�9�'3@��s@�z�e�^�Y�DBS'7�ST��J���j�j� �V����*�J"'Ũ�" �ֽ�lܓ��nI�Ϭo�IQcr=����u`����Q	/BIEu�z��{*f�ԒH�Q��@����:���9}k�:��@�#��	̉�8�q�a��\n\���W���מ��ol���3�z��`��{�|���+8���⃎g�/��4
���_U�^빠n5c17I$��w֦�]`Y+��������>�Pߑ ��	&D�z�Z�?�?���Ɓ����-}q�92$�}ܒ�`Y+���`]������_و|"����ߵ�.����o4a��u�֮�uv0%�F�Z��u�d�4zю���@Dm(�ƛj,k3��NN[��n��R0���8�y}��jE�lH9R_Z����/u��g��x�;���0�F�C��@����$�D���,�0?7YТ��>Ɠr9#�9�H�[���Ji�����K˽�_;�~_[���Ƣbw6UլJ_<� ����5ֹ��
?�������c^���xE$P�_7X$�[��7ذ{l�&BQ����w�~���7�ʜ����.4�l���V�����9Ϝ;�R��m��OfN\=p���%m�$ͻ[s۷���:|�k>^���k˻*�۰�]0.T��n\��h���]ك�=�Ӡ'�qw)m��<�޸�	c�t��8��m��anS���x�С�-��왰��4�`�k&�����;��G���:�b��鸮r[+sΟ���ݾl��	C��u���v�.����Y�F�4t�^��hr�<]�W/\�ƌ�n�Ξ*�\�f�5i������8�^,^�?�H9���;��T�vv�rI.���Σo�L���:�ǲH�Y��s4�����SU.�=ex�������'M�����^���Z׮�ץ4�}cx�E$�D9�H�u�p�
7�~_�|�g�� ��߽��K=�uD7yͲ;t�:�\h����wG6���i	��]�0��R#����`z��,�0&����K���j��U��W7Suk ׶̘Q�%p�%��(Y��߫ }Z� ��ŀn5c19(���@���@����Σo�$���Gwj\�w�0%R��W�	gQ�7֦��5&<rdI��m���]��Jh���_U�U�*������n�y1���,zn�ۯV:Ӣ��M������2��q�r'�$Q�'1%&hzS@����*�X��`z��R�]���HN)$4_Z�ؑ|޾��:�������9�I#QH����>z�a*�)����	A�J#-��W�z��ԛrH�Lq�JE�}z�0%�F�Z��u��}n%ܱwr�7�-����W�	��0%R�׮�g�	�	�F���Q^]¦���ˎK+��������W8i�����wco�L	T�����^��/�u	�F�Q)���[�d��X���>�پ�I%27Z�M�x㘆�����:�nhz�h���_U�u덽MH�5�H$���
_>��;�X��8�Z�D">����lܓ�w���5�.jo-�ܻWco�L	T�����^���y���E&H52)�q�4�*��B�ͷ8�l�B&�l�����|���$�D9�H�|�빠u빠r�נ_�]I�$�4�ĤZ׫���`M���*�_ٙ�{g�b]9#M7�9������^���Z׮�u�ӭbr<QG$��l��`�\�=x�:!D�}�`u�o�pL�6�H����>�w4z�`?7X�DG�sUR�K&Ԓ�V��H�J������Cg/[�B�om����n]�-���j�.���ln��غ����t:;��6��˷!�Sf���/n�z���I�CXv�.qnH{l�l�[����h�%H��������Nt�zΦ����-��;�32����s���Yیs���>���wm��YJ�GNx6ԃx7��W����W�؝L7�޻�����|��#V���t2�񋱮�b�6}t�Q�R���7o�|�#*��#g��!��m��w�ۚ^��/����3? �w�@��ƞ��#Q)����W�	��0%R��W�Y_&�H'�G3@���@���?��IG�$���ذ�{���̪�sw|���w&�]`z��,�~���R��$�4�ĤZ׮��z(�w�_����5ֹ���?~���=FF�G����79ܺ_Z�0��X��i�[�W[w]z��Vy�f�������7֦�]`z��Kqj�&��M��͗v�����	\@(�+T���(:~T?*��W~�y�,^�]���(B�%�w��n�w���ܯ�fê`��{��A�A�A�A�����b �`�`�`�����b �b��D�A����y����؃� � � �!�����#g��̵+;��������!`�����b �`�`�`�����b �`�`�`����ٱ�A�A�A�A��{�؃� � � � ����˅֩���Z�n�lA�lll}�߸lA�lll}���6 �666>��~�y���yw{�������
�Y�02�q��Ӂ�.��RwO��\�\�tvu�s!x�w��/��V]e��Mf�lA�lllg�~͈<�����k߮�A���߽���A���߽���A������ڴ��ֵ�VkS3Z͈<�����k߮�A���߽���A���߽���A�����߳b "X � � ���[��ֵ�.L�h�Z�y~��y~��yvy�0�b��0ʝ��0h l`�Hݸ��h��pX�����"��gG��� �E�tF隴�D̢aL��],3 q"���:2�!XX0F�K��Y��B�
a�l�@�X���ք�A���Y���4R%IF4���>��@8�/�	YFT!R�X!HV��E�).2.+0a��2*$��{�8��)KQ���<# �ph���!���(�U�;��_��P�p�����A�Sä���� ���~͈<�����k߮�A�������fk�jfe�f�u�6 �666>���6 �666>����y~׿]�<���)`�����b �`�`�`�}��?L�3XM]f����b �`�`�`����ٱ�A�A�A�A��{�؃� � � � ���p؃� � � � ���p؃� � � � �t������d��n�CЙ(t�����C�9�jzu`學������i����?A������]�<����{��<�����{���>�A���{��6 �666?����r6y���J���������͂�{��<�����{��<�������f�A���ߵ��b �`�`�`����fg.Z����je�ѱ�A�A�A�A��o�؃� � � � �;��lA�l~׿]�<����{��<����w���~B�t6&e���w�7{�����&A�����y����v �666=���6 �66
O���>��~�y���5)�&��f]Y�Lֵ�y~׿]�<���������?A�~���*�y��L�M6d��C��Pܓ�܈��2m�0���gf�:y�+ۭ���٧+Ii�9�H��]��Jh�W�u}V��wQ�8��n8�s4�l�y(�Tt��Xz�Ӏk׋ 5�ӣ��H�$4W��:��O�fg�W�ۚ��4_v6�$Q�5WWX�P������X��`/��-}q��9�j9n-�]��>y�����5ֹ����AD��H�$���d�"������w��y��k�ٍt���h����
N��2�gtf8�]ƆGm���
/e�#��3�(�q��s;�O��Z�j��;/��Q �N󮪋�8�k@�3�ɒ�j^�.ڐ�izP�N^�2vu8��:������iN �qK=�\���xSb�$�mƑ3����,/�h��m�6��ᧈ.Rk��4�;�ݎ7�Q.
�?}ݻ��|�Fq=u�v��{t=l� K�Kn9���͎��Q�ϖ��V(��V�������l�u�k�s��#��ذo����	ģd�$p�9^�@����]��Jh}n�c��8ҐnG�k�s�k׋J&_;� sϫ r���m&8�%"���������h�x�9^�@�����n<jD�n��n�`�ـyBuϫ������h�r�s�6䍲Db�<�Y�S�ۑ�3�[l���g.���h��g����MI#$����zW�hz����<hu�ߐ��"�D�q�_Y�IBU�(J<��gb�;� �{^�k�8<rAG#mŠu빠}����!%.y�`�p��U�4����s7eLݬ�Q�}�|��w�@���@��s@�ұ��bpQ�9�����eLEn�%���׌������p��Y�B�qx's�ٵ�nŃ�k�Ħ`Xy�s���b����|�X�������%_}�	ex��������*���/��Cn7I�9�H��w3�BS&��X�}X�M�yL�K|U8���qƣ��u��4W��?���-P�D%�P�L(Kn]�d��b��u�NG��$"�4W��>�j�:���>�w4_v7bN	�(�Mr���V�Y^0=-x��eL�7S�⦉%U�quv7�K#$���-2��aC��N*���Еe��%�8�����d��������`M����X^����I2% ғ4�����0=���W�Yׄ��f���.������eLEn�%���ט����Uj���jK�UwXP�(�w�8�ذ��X	F�(�	(�Y�?�3�f�נ_�J��n6�s�X���k��*`z+u��'�#t5�U���ۜ�؜��u�,�Rq=40��v�CjŃ��3��U�&�zZ�6ʘ��`K+�-Ů�Ӎ���I�+��s�hz�hu��/��N	�F�Q����s�k׋IDξ�X�}X�px�ȓ��qhz�hz�h�W�u}V���obx������k׋ �:�����pz�ܓ�/�,UbE����.L��8��m��G0��*y�gbYGjݭ����۶�ƺ3ɹ�����//:�΍�4�,S���vA���	�n��R�˘����F���|bI�b��5)`i��s��%�i-��X/8d[+udc����';��ݹ7>ٸ7F��r�v��n����G$`!�^(��݋�c��eˌW]��O
��;m�c�������;�w˵��n����Y9#��|��9m�֦�.��:���Me阜b�H���}�zW�hz�hz�hg�X�ɑ�h���T���W�	ex��eL�tIF�i1�1)�׮�׮���zW�h�uq���G3@�+��*`J����`�Z��8�"I#��r�^���Z^��^��e�������"�,d꿳A��>Q��zĭS��R�X�Ns7hޢanF��#rG��|��w4�w4W��-}q��H1�$i����c^P�(J.��ذ=ΰu�p��{�$x�)���u빠r���*�X��`{�!,����H�����`M���*�X��`K+����$ɑ�h���_U�}u��5�ŀl�u�t%�v��&ꧮ�RKv��u���t�\k�R�ػ��0��.d+��ٳ��Ye3pQ�������0%��m�L��v]�?l�Z�f��$�.[˱�=;8l�LT����s@:�n������9�+��I�g}w4��F"0�U��
?BJ�{��z�`?j�w3VUڻ��wr`J����`K+�fb���@���4��I5#�n-Y^0%��o�L	T����bڴ6�xz������$��BN$�T��%WܻL��\��g���,������W�	��0%R��W�'T%�dN	��m�3@���@�����s@��s@�>�ę28�Mc�=U.�=ex��W�	��0/�+�8�m&9�bR-��s@��s@���nO��B
�E�A׿s���u�ӏpm�j9�^���Z��u��+�	0J�����K�K��������E&-)�Gy(�s�4bq�NNG��j9�/�zU.�=ex��W�	���v��{�ܹr�L	T�����Y^0&�����cN�#��D�Z׮��W�	��0%R�Yq$�f�o���wWcY^0&����K�Y^h�V7�dN	��m�3@���@�Z� ��ŀk׋ Չ\
!"	0�"�d�$�D��1�@��,	�_*d��"� FxIiV�Jf����"��[�R��	B�� � ����L3v�#`�HH�$P ��� �@�0X � ��*� "e�B+�A 
D#��$X@��#��L�$IXF0j�R�Cpٰ��_�I�D�(�©*�&@IV�;R	�$$X���$P"RSi�$T��@#!��Ds����Zֵ֤�m  n�U�,Ų��!��`�ԛ���D�+Oa����i�	I����-:�L�]�����+k$V��n��cP5䣀�-��r]&嗵�.H��f��\��B\aJm���6�Ϋ����8�Cϣm9	��/F�N�P@]�-嬢�m�����t�f�̩���ۣT�:LFB%�9&�\'enf��nYMlf�7��E��d�V��FR�Ƥ�r�ZB����y�:����Z�w�쵞�=�=�܈^L���a���;m���e�y(��n� b����c\�0=b9qZN;8�5�I��̂�����Y �N@k[���_�>��\�5m��cw�l]b�5̪�7]UJI���:�D6S�ۛ�23�)�qa暗��˛���y�	Ta����2���q����um���q�[�@<���bZ`R]R���WYnbQ�ۧD ]S�-�����\2h�/ZZ ��m��Z1�Rjݺ�I*��Ѽ[��S�ڵ��܍����vT5�ƃ׮g@f�'c!��vS��zZ��i���_[�vS�^������ڶ��Z��.�6�5L�ƹ�mS���g
N݋K��tn��J��ł��z�u�`tdޫ�79�^�s�y�k�qϜb�e� 3c@�����Q�q:����	;l��
F��;N���^�==OF�a,��z��RU��:�KI��{揝+����[�!�k*!ms垸��cl�%�S��Y�l�8�[V�]�B�,�K���]��8�3�^ۤ���v��fˀe3���1��(�6w6P\�|������z���r%mlpY�r4p� ��O#U*�*��b����kb�r�m�G��lv4T��f���2��ѭ����kA��r��F9fQ�:f�&�WQ���Rl*+�[oզ���V����jZ^u͐%�1�OG&F`���V�:�U��ya���3��kR�j�TuvFu�?@4��"z�v*�T�T��=t?�)����E^�.�7ٯ.;q�f�m��G#x9����2����v9uB:\�q���]h�-�䋊����gu��T��;&�|���	�u��n#��j�Z����V�����-���Y�^nΰf�Y���?�|l�Ʊ��A6�u� ���b��gY���w6��m�9�Gnw[j{:K�/�oh�s�M������;Oc����<ӹP�1[�JK�s:��{��߼ߝ�˱��6K��cF1 �*�2 ^ln�ė�b�E���|o�:�W5?�o����0z��,�}j`_NW\�!k�1)��빿�/��4
��zW�o�3��������4��m��f���b�6~n��)���p�ذ[Ɲ1��Ԏ5��ֽ���]������V�zQ7 �qU]�����o>�� ��,g���������͵k�]A-ϡ�v9�/:��/��:���+�"����{��r�Y=6��\���>�<`K+��Z��V�׮6�<R(2% ғ4�w5g���@ꢟ��O����?g���]������"pM7#s4_Z��u��+���`{=z��;������U����"W{;Ӏ?w�`��7֦��q%�r�{f�v�=ex��W�	��0%R� �o�߻���P��x���s�x^�܃ mv�v����pDz���\�-��&ʬ�6�z�`?7X��<�BQ�Cy�- ��4�c�5��j9�/�zU.�=ex��W�	�o�Ի�������5ֹ�>z�a�"-DB^PB��F@?���Z� D!D/ݗذ�����T�)M��E]]]�W8����`��,g�� �z��\m�x�Pd#�%&h���<�(P�{��y�`=x�����
�qk��(��F����C6��:��m=�ҁn�����'����x��n9w*[˰Z�?��Xl���+���hg�X�$�$��h�W���5�ŀ>}� �����j���詢n�S7u�}��`���СBI}_��
�|���F�x��m��R�`yBR���|�p���*!(K�4LAE����rI��2�c�3�Is4��Z��3?����[���]��v;�E$�LKqj�B���'qո��9ި#1F�k\m�f�T���	#��-����빠u빠~�ڴ]�N����%M]`}�zd|���t�/]g�g�G�}��O�Ȥ����s@�����eLz׌Yׄ��Y�.�ٻ�������6ʘ��˹�v}e�2dn@h����W�r����~��X��u�Z���/(�(��]�6Ih�4�X���*�8J���Ĺܶ�t:;I��:^��8���d��ocU�_N�p�:=�;/l=��U m�wn��>x� �9��t��i�v���*񓝺��hӔ��CA:��BwMk�J�+I#���K��G�0*N�a��;E���:���8m�/a�Q����;�Ǟ{!q"ć�]>2�Й�vS'gg�6&��=�MW@�����������q�ܻ�*f�MvI�nLd�n�=���k;5c��YSA+`���NI6�dĤ����h��7֦�*`~�J-\�yp�n8�s4�w7�g�E]�=�_=��s@:�i���ډ�䙠r�נM������6Am�[ڔ�H��G�r�^����hz�h������Ͻ�Uh���I2G�8�z׌	ex������eL��^�������k[] P�/jp�����C#��&�8�ě7k�u*i �s�������6ʘ����L�Z&��fj�nhܓ����ډ��$��篫 m�,^�X�;u3D�܀�I�H�W��>����]����@�r�i�#Ҍ���C��}��`_���Z�l���}n-\�yp�K�.K��,��Z�l�@��w4�;��<���2F���u��G9n�I�^�x�n�B�7<���lj�#���N7$����@�z�����;��X���75WsUe�U�0&�S޵�Y^0=��0&�&�x��Ԏ6�z�[��u빧���Ȑ� �
�ܾ��`r���\i��H���Nf�����g�&�*`z���:�I�(�sNf���^���z׮�׮��[�<���<�H�pr,ql<79���i��&�uv�*$�7I���na�z��_L��)1I�*���>�w4�w4_Z��)F�r0m(ɉH���`K+��Z�l���}n4��m��f�׮���^��J�_=�}���i���i����6~n������X%"@�	 B2Ba$I�
F�;[���?.����7����:�>z�`���6~n�(�	�,�����z+km_�����;��L�#��ɑ��.�[�B.���������S�Fa����x��W�	��0&�SYq'��"�HD���]��ֽ����]��$w����INbJ�`w��������}� |��ŕ�ɑ�����W�}z�hz�h����R�8�`�Q��&����7֦�*`\�PE�B^�����]D��Du�]8�MZi�O��<K�7Ri��`˩�7�����ڌ�CG	�ă������i{��j<���Ս8�Ć�lkai���>2��=n�J-ãn,;j�m��u����tӛ<�Z��n���m����<�ӝXҚy<��s�� �-���6ȴI�{p. ��=�ӓOg�Ê�1�^�gga�}T�"mD��[te��֮jV	y�ꓓ[���t8۵�jN'I���X�l�V�*�$Ɯx��m8�Q��/���9}j`M�����Z����	r�#�f���^��H���@�_nhz�o�ă�����p���W������Y^0&���� ���{�b���U]`z!B��ߖ ��,g�������>���SXR���EsvL�Z�5�ŀy:����}X�^,ӽ�4:"S&1(�
'��O��\*t�g1ۦ�1FgJ��F&�E�2�n����W힉��N�����:V���<�a$z+��߳�#�׌	ex���S�t�^_j�˹[�������_�0%��o�LW��?/�ƤxG�qȣ��u����Sm�0=ex�$���˻���������l��`��}_��}�@��s@��R9��D�X�ӻ�?)v9;��=�/N]L�l�G����Ms�qV��[$Mț�M��W����빠u빠r�נr���S�$xƜq4��>��`���6~n����ВS#�ʓ��qAI���__nh���`p(=b���$&��E,$��
@[m6�j@�!�:��B�s���H�T�a��R9�1�kF��:�lH��`��61��Ni#�0�Q V!RP�D�ІPd�b��V��
K�N*@R&�	Ԍ�4�(Ƭ��d�Ą$"�"�R��������-�l�!��H�0��*����C�y��%FB	�z��F��V��BX��Pp�Tz&�QAp�M� ����4��|�Dz
�_�
 �_���{��rO{�ٹ'��X�HD�H�sNf����U���
�~LY^0%���/U���K�mY7wX��X�������ذ?�~�6ߟ�~��1,������}���u`���[�qf�-r	��L���jh�����`=x�z�`?7^Q�
�|��{�ԏ��N9s4��`?7X��X�^,�Q�
J�;�T���UuUw7v���V�eLY^0%��l�����.�Wj������RB��X�XB��bw���"X��!����P#E#`�T����}>�����bX�'���/��ֵ�d�kW35�ND�,K��l���%�a�
�}�߾6�D�,K�~�Mı,K���6��bX�=�_p����vzK3��q�n��Iĩ��J�6x�j�/f��l�ō��j�sDND�,K߽��ӑ,K��_{17ı,N���r%�b����"��$)!=�tJ�����段-��iȖ%�bw/������r&D�=���6��bX�'�~͑7ı,N����Kı>���[�F�5�0��u�f&�X�%���}�ND�,K��֢n%�bX��}�iȖ%�bw/����bX�'>׽�sU4X�pS�������oq���ov�X�%��w�6��bX�'r�ى��%����u���fӑ,K�w����)�6Tf&�������d��ND�,K�}���Kı;��iȖ%�b^���Mı,K��!�~��2?�e�ѣ%ќ޻FMe-�(�wa����]��!�����D�E����X[�8+l��~��yݸ��8�ڳ��q��&���r�#E7=s11�<(�amو(e���n�ѹ��s���l�6��겶=;q�R��m�Z�P��^�c���ݻ;67�!�� �1������zzX�),��l�ɓt��cD��i�/k�����}��x�ߟ;/��ђ������v<"c�k�Su=��{��4�Q���d9p�J�S�em]kG��,K����ى��%�bw=�fӑ,KĽ�����bX�'}�p�r%�bX�����I�W3Z�����bn%�bX��wٴ�?�H�L�b_~��D�Kı=�߸m9ı,N���q,K��}�/��ֵ�d�kW35�ND�,K��֢n%�bX��}�iȖ%�bw/����bX�'s��m9ı,w�\��浅������ԉ��%�bw���"X�%�ܾ�bn%�bX��wٴ�K����2&{��ԉ��%�b~���㚂�n���{��7������q,K��{�ͧ"X�%�{�f�Mı,K��m9ı,�~���j��\�/Mr��aOt�X/7l�7g=���<�J��:4��4mkY���%�bw=�fӑ,KĽ�R&�X�%��w�6��bX�'�����oq��������Q�MN���m9ı,K��5"n ? �8��D��dK߾��ӑ,K��_߳q,K��{�ͧ"Y�7������䧴�Q+T�{�oqı;���ӑ,K��/����bX�'s��m9ı,K��5"n!����~�����TnRY*����,K��bn%�bX��wٴ�Kı/{�ԉ��%�bw���#���ow��r}�HZ�Z_w��ı,N���r%�bX~D9�~�H��bX�'�{��"X�%��~�����oq�ߟu���1d�A[�L]�� ���}����������������;j�h^Jzh��B����oq����}���&�X�%��w�6��bX�'�}���Kı;��iȖ%�`��0~g�,n�$[ow��7���{�~����Kı>��f&�X�%���}�ND�,K���H���"�S"������Ջ�a�����7��,N���17ı,N���r%���X�?�0��������7ı,O�{��"X�%��=�e�5usVM�Y�k17ı,N���r%�bX���jD�Kı;���ӑ,K��/����bX�'>׽r�d�u���w���oq������ݸ�%�a�A�B���t�v%�bX�������bX�'s��m9ĳ�oq��~�ݧ�z�g���@s�����@Ѷ��j�T��A:^t�y�l��2m�]kZֵ��bX�'}�p�r%�bX�e��q,K��{�ͧ"X�%���z�Mı,K���s��f�����j�Z6��bX�'�}���Kı;��iȖ%�bw�ޡq,K���ND�S"X��d��R$-hZ_w��7���{������̖%�bw�ޡq,K���ND�,K��bn%�bX�Ϻe���kZ0�ֲ�f�iȖ%�bw�ޡq,K���ND�,K��bn%�`b®�@8)�o"w�o��r%�bX?w�\�YsZ��Z�[.���bX�'}�p�r%�bX 
�����b}ı,O����6��bX�'{��7ı,Nt�t*��ݪ`��q��r�͒�R�lWOg��&�i3%yajq�X�'M�7|�Ȗ%�b}���Mı,K���6��bX�'{��7ı,N���w���oq�߻}����;\�T���%�bw=�fӑ,K��}�B&�X�%��w�6��bX�'�}���O�!�2%��u��eɬֳYuu�t[�ͧ"X�%��~ޡq,K���ND��!�2'r�����bX�'���fӑ,KĽ�s�]f�f\.��kZ�Mı,K��m9ı,O��ى��%�bw=�fӑ,K�Ȟ��j7ı,K���S��V����{��7����}�bn%�bX(�}����O�X�%��߷�D�Kı;���ӑ,K7��{��O�8㾗=�+l�z3���.0ٮ�\�-�u�n�\����iG�b���,���M�L7�̎!5�������E������wkB���Wf�֞.�M���0�9yI����1�B%�%��+�s�KTn^�&�/lW��;.��Gӭ�p��ݯZm� �1�St5l>6���q�F;Z_`جےoE&������!�YZ�FZ�z�n�{�w�{��>~w�^����[�!����1��;1����\u�VG��vݺ��*�39�Zд��ؖ%�b~Ͽ{6��bX�'}��7ı,N����'�2%�b�OuT,!I
HRBu�T�қ���������r%�bX����D�Kı;���ӑ,K��_{17ı,N���r'��TȖ�~2��5�XkY�m֡q,K���~��Kı;���Mı�XdL����ٴ�Kı=�����bX�'��s-3ZԺ5u�Y�-�ND�,K�}���Kı;��iȖ%�bw�ޡq,K���ND�,K�=�e�5f�Y&��[�k17ı,N���r%�bX,}���"r%�bX����6��bX�'�}���Kı/�C�w\g�.�r���\jC��ɒ��[c��8�����[�k<T#��"R�g�r%�bX�﷨D�Kı;���ӑ,K��/���$�L�bX�\������$)}J���]YUSJoZ�kP���%�bw���!�M�!Y	���@4
6Ȗ%���bn%�bX��{ٴ�Kı;�oP���%�b^��L�5���[��eִm9ı,N���q,K��{�ͧ"X�!��=���"n%�bX����6��bX�'�{��sҴ-�i}�7���{���~��6��bX�'{��7ı,N����Kı>��f&�X�%����_k�]L�sZ�3Y��Kı;�oP���%�bw���"X�%��_{17ı,N���r%�bX�t>�#8:oh���[N�Ít��:'.J�H�Gj�\ݪy����_.G�xi�t֒�P�Ȗ%�b{��p�r%�bX�e��q,K��{�ͧ"X�%��yb!a
HRB���D���m\�\�nh�r%�bX�e��q,K��{�ͧ"X�%���z�Mı,K��m9ı,N��{-3Rk5�h�պֳq,K��{�ͧ"X�%���z�Mı��p���%�z�����ȟD�����r%�b]��O��}�7���{����_~��f��-�fӑ,K��}�B&�X�%��w�6��bX�'�}���K��QdOk��fӑ,Kľ��f~�5��2au�kZ�"n%�bX��}�iȖ%�b}���Mı,K���6��bX�'{��7ı,O��.M���mҖ������0 �ݜ��"nmq�x�cW?�Ϗ̏����%�����X�%�ܿ�f&�X�%���}�ND�,K�����bX�'}�p�s{��7����~����Z�Z_wȖ%�bw=�fӐ�U�L�b{߷�D�Kı=�߸m9ı,O����|��{��7���~�}�j%�Y��m9ı,N���"n%�bX��}�iȖ?�@!�2'r�����bX�'���fӑ,K��|e��.kX�Suh*�D,!I
NIzR�{��!r%�bX�������bX�'s��m9İ*"?�?�P2'��������ow�߿߈sV.��r��,K��/����bX�'}�siȖ%�bw�ޡq,K���ND�,K����D�sP�j[�]kSYgs���]����D).)R71�Ŧ�ڤ�5f�Y&��[�k17ı,N���ӑ,K��}�B&�X�%��w�6� �Kؚ�bX�������bX��~����GK6-:�7�w���oq���������,O~��ND�,K�~�Mı,K�ﹴ�K7�������x��ɪjݽ�7��bX��}�iȖ%�b}���Mı,K�ﹴ�Kı;�oP���%�bS��˞���L�Y�˭h�r%�g�"wW����Kı=�߹��Kı;�oP���%���"{��|m���7���{�S�/��Jж���%�bw��6��bX�Ƞ����B	 �'�{��pI��n��I�AEE�AEE�QQ_��QQZ�����
*+�((���H(���*�"��
"A��@X � ��"E��@ �!B"!U������TW�
*+PQQ^(��� �����TW�QQ_�AEE��h(��PQQ_��PVI��i]&]�Z��` �����[�� ��           
         �@B��J�� B"�JQ � �H�UH��T�T�"B��D�*�J�P( (ER��P�*�   � 
   P
��O�'�b=���&^�V����D���ס��������ֻϥw��=�� �y���`  Kb)DJ��"  �  	�
BP ���@     r  � 0 6h D����� r   :� R�D tgf��� ��� �JPD� Q�@v}�w�T\�S'�js=y켲���Q�z@ޔ���zڹL�w���=� �  @
   b �T����=�G��\��6�m� p��}z�{t�c�����z
>�y�}�zz8�� -��7��8 ��/m��w۫�L_g}oR�� g*b���k�qt�qڕ���� (    ��;��g�*�׶n7K�x����*Y=t��[�Zr����� ���r|���}| >�d9�     @s�fiv��=/y��x���o���_[�ip ��      �{�Ov��������b]�l�{�i�g��m�g��y����M� 
�=}.,�� 7v��g��4�������r}�W�Ͻ���i�_{�U�Ӻ��n�tx��zy5�ܡ�Q�M�%J�2�C�SeJT   D��R�L �D�*�&�*��db41O�BSmT�J�40��IJi ��"w������������;��w���
��,���AD?���(*+����TAS���_�HJ��jj?�FBBD�L!p�)���n��� Q�!p�GD��LR��&��#!t�x
b1�̐�c)�& ��F�D�
2��)���e=!qC!q���)�M�NjɎUː$�(K�.0�����c 4@�S!\YB�Bncy0!F�'�q�aJ�L-�NS��t8�`�&�C7<��6Bi挡�|BM���_x�B�����Li�3Єa���xI$�&����.r���
o&p�0!!��ӐY˦��=$&7�#X0�(X�B40HS3�������x�搹� ��{7�{n�����;���?n�5�&���1�1���IYVP�ژJd.;�$cLӕ��a	�l�)-��+4e����VV����%���f���<X ��H���U�noᒰӌ������#L&i˦�����sx��Rn@�١���%�P#��L���g',,#�/8|��9�I�����&i.l��<�&o)|y����e�G>?�s7��oW����|�~7O�bqm����%<�eÜ8@�'Շy����5t��Y7�������fi�T�X1!B���X�%X%J�� A�!B�+�sr�(�Z�`i��H@ 1H�`
%04cS�\x� �CNjBh@�,H�|aI��8�((˛�E$��r�St7�8�1t���:��s5��f�,�Cх2��t��t%� I���$$�x��H\�Zn]�7�=w͐А8i��H�,�x} O��B�)����|�}�ln�!�2!��j]v��Ò�lI���hH�q�d��nMͰ�G�!H]9c�+�
Aj�X�������tX`B�q��|OC���	�	�p���$!\�C��no����!$s���Lwy-�I,�>S�#�bS4��e�����=	sS��	sL!n�^o\Ԕ�Iq���8x!!p���O=���9B1��f�$��ys8ɘ�uxxKn�2bc$�A��Yk
���2��������5rFP)��77�A)CHY��3e�T��ϼ)���Q�X4a$%10 `x0��`C�WÑ�0()!��)��	@�]���h�y3�zz�I���10�$X���,�(��:�H��8<����d�p�88�|	����0+�hE*���M9��ݗt��K���L8���|��COT��D���8l�I��8y̴=�$)M�jJc<!��
V�(V�2��yn�S[�dy�=f�GYq4�<x�.2��aa9�$*D��N���	�Ѕ2�&�3vp�!M+-�IF@��ej�	"��OL���5�{�=�5dJAai�@����)B-�C�d���4a_4��P����3]9��f����sy��4�F�U��q�1xa32� B����Hѩ
S_�0ґ�`����ׄu�e�L�a��XV��B�p&0�5��s��Hl�vH�y���4��t���V�>�� ����d!P�G�I����B�H0�(�p�\6��|c��)|䑃�B�o-�y&��I9L9"��� ԁ�a]0�p��=�K3Nn�(`8[��k43�u��8i�+H���P��	$y���<��/9����\�|�O>HWĮ�N$J�
z����lV�(bh	��!x��āS4� �X�蜌�V�`RMN, @�*�A*�jby���� WP��O�!t5H�6��фC˗�>|��Iw�o��LFW�S���
����:�<�7n�s���7��w�|�$����%v��&�0#0`TRf� ���{������q˒�$���B�&*b0�.L�y�%�x�y��� HK�������5燧��1��B�D�k
�L���<��ND)��,*J�{����o���0�S ��%0��B��!C� �v�eˢ4�#D��"���yŜ�|�L �9u#F!0��(�q����/�����8FB�(fg	���<��%���d�g��$�nrq�燓<���!��0�p�	s�
F	����ab\-!i\sww�%�8ʑ)�3�aB\ӗ�<�ϟ"T�4�<)C�7Ԕ���,��0��78�q"�8��B�.B��&&bK�q|u!��9�	w��|/y�g4�D�|���L�2�q���I+����\���3|e���JI�.$�xp�<�Kn�<����<N$x0�ڌ
8j���Jc��]��' �\|%b�!B30���F�k��D�q"Ӟ�͛��F!�2S���*���	�`.�'ܶ`r�$�9��"�������g����O����`<>���G�)�aVX�ă	L4e0ЍF2*�S������!%��Hn:kL��������8���41`WD��̬�ɆF�k�����Ja�.L��^!,��	ro=Ix��K�ȅ�Sd��r�SX���B���\R\%���n�%�����xi�
�����B��B���}�ۼ|a����H�0)���g���t��<�x�+r�� ��a�bF�M��\�'�=��!�1e"L%\��v�T`#�)��y|��,)(1�a,c��$JB��a��J������� �rSA�p�ō,�\4��F�k��b`�]�&��А�T�\���#cpH$�0�B5�+Pb�xE!�� �d8�p�>��D�`H��V'���@$d�Ȇ�)�E4H�c�j�n`F�Bʰٴ�L	"��P���NX�}�y���ĭH�#!��Xz�2h��C�Y�cG�-lk�����5�p�$�[J��nq��$�3��A`Q`V�n�_���m�3t��jq�g����<����bT3p��$�\f��(�F���\M!iK�Ó���y0Ӌڛ����&I��`e�;p�K����O8q���J�����������"W4*�|j@�Ja�<9����#���y�a�2L����0�8A��D�@!�%8�g���k��R+P)�A�P��AH,8�o�!*��fBe������-����>O�Bq�-
�4O��!�20�ę"i�HȱNIt�imrR����v@|�;�Ú����).f>I���1������|�y!,���B��|8��I�|�=O�$
�o9��0`Za���"����{B����c�%I��Ri�8Y�V崖�Ym��F�P�����#��%3YÒ.�dn!��f��ͬ����#H�@��cL�ɶ��S4!S �"���
��@�aJ�	#*�f��ZD��3"���b�(hA`�)���e%�:��!
}+�K��Ip�X�F��@bH@bT��2# �"P�X�!�S�+�-�vRP�!,��i��r_27�\q#p2S�����b����o�,�iő�OfL�$@��u�0�k�i�1"��5��'�,���<D��K&.���\I' �	�x?K&+�*¥�HQ� �{paL#6�d	\r�� � 2��4"�>C�S���A"�7HxR�)[y�(\H��s5�`�-7ÀE�
D�`hi�:$H.�D�B���_�W	FQ��.��d��}�ഘ��d	�
lX$�e2f�3ި}�(G���`4��V5H�ĀU"�SB���n!�F��!���������ww@l�Ŷ�YCp9�m� 8��r����}�͒�݊U2-[]T�$   -�ܐ �I6 � �  8�5 	 [@�h m��M�� -��#E ����6 �n   N�i�YYbnܹjU��vS�$Ur�1@j^&��T�U[+�%ZT��2D�]T�\�s}��*۵+��r�e�h   zY[t�e6�v��{����>����, s���&�.��p��$�kzk�cuV8�h� N���[p.��<  Ʀ��� M�K(��I�lA�r-�m��o���8I��۵��0H �6�����[���6�k��c[�Ypm�]6U�
�v���ڎ8�t[R��O5)-J�rs��l�` H8H �I�F� �WR����T�K�꨽im �`����s�8HC�vն[@k3����`-� m:l����߂C鵵�yv-��ڥ�7V�Juʼ�6��:�� �9�m&�$p ��y{eZ��C���^���CN�zJ [d�-׬�m�k�nH<�c�6�M�l�E�@k�����hioYhu�@ֱān���m����  )�@^����-�����[W7` q-���m��H-� �����;�oS@TUT� m�\ 8-��H9�N�m��mB�  H �����$�鵴  }o�wͶ��  -�m���|���l� l 9��kz�� $   "� p#����рpH-���UT��m���7m"��\a��)t�҃mڦ��tV݊��vN0&��ͻ�*�����􌁞��tM�I��8�bC����Ү���ibc�=v�]��$�t�Ԇ�&�vμ5]R� Քe�i�<�f���t�#�n 2�.��1�T����R�l�I�JM�:�f��)UP65�혥�UUUAŨ]���5wl�h�s�ʹ��[v��   p�q�lը7�z�E.��6wC�m��Ua�5Q�����偶� n݉ �v�a�׎� �&k:��ir�s���*UBc+���z(�F�o0 ڴ�tӣM��f��m�	͢��W� V;Q.Ƚ6ݰk[�� �3H =�u2Ei�Sc���6؝���V�T��j��`�#Z$��y� :��+(Ԅ�;wYƻM��nۖk�� �6�&m�-���k�P$�ݭ�ioK[�`8 �T��  8���i6�f�ڹy�W�m��/(�ۚm��[[l�@h	�	 :�jݤ�J]��H\.s��mm������!m���	  �� 8�I�����Am�v�  �]!����� �ܶ� m� [m��P�I$�� p 8$m��`���sN�j�D��m��kGG��m� �h-����4�@���� t�gGgL d�$ ����� z�� ��I� m�E�����XVݍ�d����� m����@�oD��*�ԃ<�]J�8�۵��m���K��E��Y2�],+�`�u"�-R���R�mUVy�3J��C���΀�]X�^��yk��qŷ�m����[v4�B�m8��M/��}�}uc�j|�a�t���8���1�N�]��h�[b�Mb��5�i�[h 8p�Y�pOni+��[R  [%$��3�.�%v����A!5���i$�m� 6�K����!�l$M����BD�4�Sd���[@ p����P��!+��!��[ZE�ʲ�X�f��d Hlp���on�I7m&p8ΛV�e   H8�E$[\HM|�+�̬k8������� -��m�f�$^�T�i%Ŵ�x^� *RU�j�I~~� �I@���-ۜ �u��:�����Ps�Uk�X��Mz�rss��\�9'BHm�]R�[V��=�l1uJ�,�Kr�����.��D7eM��ݶj�׬6�at�nn��kz�^lh�ۙh �5F;cT��Mr�u*�+F��5]6۩q�ku�)W��-��_o��U�������+Utn5*ԥ[Q\l���s�R�I������(!�%-��:������D �f�Z ���YM*���l�$�mpp�dn�wl�c�][
���1 婗f��]���-�[`�GY ,�M��vA�n����a�m������.Q9K�"��i����z�}�Vq �S��^T�����Ғ�	�K���V�  	<��`Yդ�k�&�cn�mp9�*�yU檗�k:����f�,�Cm�U��.�6�K}rI�  [E�H���m�U�U�����uN8���@okլ0�Ѫ�n�ض�Gn=Z�
W�0qx�D�F�v����6ۆ��&-�-�o�/N�VE���z�;�-/*�V8������ծ� �����ަJ/c����hj���Rd,�4��@_+��T��B�kmʶ��kM������rN����$�F9���e�7lV�'m��J��r��ʽngqSv�*��΁��:�m-�)!Ëh  ۶8�5��v춭�  -�h   ��@:��d�&ҟ�ԧܳ�����yS#=��l٦ÁMm�n��rI6Ͱ��6��I� �[@ G$6��M�nE�.��A��ؕn����[8�EPgmĭT	�Un;=��`�H�hqm��� �H�6m��|�|��+���X�+��j��ҫ���*��g'�M@U�P&���f"�۵�]0�f�{/�ͺ���V�Lq���j(���Ś��r����*1PX�hS��vZ�[@9t�m���m[ N�I#k�$��q�kn����ٸį5U��mm�A�q<�R�����[R�UI��+��ݍ�Pe�v��1�	�B�s�!u�j6�����vUY-�M`Hqd�A��fum-הνd�6� 6� �z�m�߃}�Ҽʪ�U�UUR�8�sE��-�,�jC���jys����`. ���蠽Zp�ն���mk��8N�m[Kn�۸$A����r�m#l �kkmؐ��Z���G	8 "Ŷ�-6 .J8���6��m��  hYG$�`���z����6���-�&ʳ�#mm�ݶ$$�	 nݛv�j�a��pӀ��]6$$�-��6��m[ִ�I��K�^�5]tq�]NĨKT�me�u�u�[d$�[N$m  *��{s��`N��-��H��i����f�%��\@R��s��@T.� �+��ɱm��}�G�V�]��R�m�2H�x=1���d����h:����mm   K���g��6���m�  U*�KČU*�U-m�`-��V�k�� m�N�[G��d�M��ր�`    m����[\�����@ ���m3 6݋h -1\�s���j��/ KP	�$� n�.��>  �K�� v���� �J��� 8m�Kh���m�   &�6�  'm��'D5��CI�� mp�A"E� h   
��&Em�u3�-Oh��s���mv�p �lm��f[�T�@ $��6�Um���B�ʪ�p��n���B��U�� -��[E����&�8  �[�mm6ͱl��09 n��u(�4��ٶ�`X�U� 5,i�Pz��m&6��h���9Ͷ�m��� ֲC}�πM��״� {�`�c���I���m �agHAۤm��gm�>���   �J�9��mUR�2#��FtC��[�,�Z�g[�� [A�lmf�m��I������cj�l�h�f�k��,�3l*�B`���WE�*�Z���a��UU���+�UT�A�p��7]&m[-�b� a�jڥ�ld m��[��m	oV6ۀ9my��W�`�V��z���ೄ%%�2��T���B�lj6��f��5출6�p
��P.��v(5�Y  ����am[%�%jR�j�P�l�0k�n�  kNw��V���gkm� ��V���@ �F��_+�i@Z�j�&����5� �&��/ƥh3��h zmkX�Nv4b��b���P�ñ[k��[]7#7GP�@���Bu����"ڥ���[R m�E�l ������m� U���#;,��`XL�c)T�v�**]U]O ����xj�I ����Y���*�ThHb��mn���]Wj�X�!�RI��-ɳ� 3I=�����v�J rm[`H e:�t�m�*�i'�.�F�5A��-�� 	$%�GR��FYe]�n �T
��@$6�m-� �-��mm [S�M6�)�7w?�TAR��6�B�A4T���`5�"� �
��� �_>G��A�> ��j �x�p �U48��<@S�p�D@=�TV�	�H.��� !�*x����<L_�> A�N�EQ2 <T�V�w��ު��(j#��P8�(��~q@`#"�x"|*@8��|��"� "x��j���U`EC�J"�TO�pL _EA��j���t��`|x�A�E~u@}6 ā,�"E�A�#��$B0 10�R"�" F	H$��,���$`D�!!����MQ_U����=D(��'�)�=&��*�Dz8"3�pD|=UN
��� �(���|*�¯���@�@��S�8? �(x�A�C�@>A���T�F�x��*�Ea�
D~P�:��`��EN�+�<ת�wTU���D _�@S�Ax
�W���Q�z� z�%F'QS�Q=�
����/���̷��%�2陹�7fZ��֧Yy:q:�FYf�%�k�'Z�F�Rј����6gN�I�n�VG@�v��6ܹW��s���]U�Y8[iە�P�q�u����O� ��F؅:%��x�v���k�s`��&}nз:�I����8Vm��k�M*�g�O&��np�"mۖA��̤����u��˹���zm�]���d!�gh�\�vf���$�8*w��鱗ے3��� .`��r��L�y+�xfq.C���If�^��dӻ[���Kv���q��8��i�ڤxF�ru�uV�6����j��iݵ��Ve3vcrmV�`�[^%���*��q�k�v5�`X�0a5�8������e�T;\�9��.�c`;]�XP��-j%^�Ƶ�tVK�}C��:Yd���Cf���/6�k���q���M��	���1�}Դ���6��6���k���x���ʬ��[�ݷ�y�P��e��B������ê�����p�Yb�A�F������S��&�Y9� qeLi�����.��آs����0qk�R�cp��7��0��ȯO�7Gn)h�@u�<{ʡ��dR�n�P�f�T�<ѳ��	����b���Ȯ;f7K�۷%�.�g��z�ʐ\U�+��\D-�Z�uf��lp]s�KV�L��Ӄ�EU8�Z��j�sE����[�Zv1��g�]�Gi΃q���m�ҽ����`�� n,,QT�Ε���Gjmn ���%�*��ٹ^R.T��[T����sIOes%]rr`0ܪ�$x�d�nk{D�ʭ���`�N˹�G*���iQ��t���Z�H��8�j��:Q��K-��s�Q�̇�ݝ����!����պ[d׵�=d���[ȓWT��$� Kqv�cRFMr�_/)��v_O[E0Fݽ�\j�Ŭ���lN �Uk�ڮ`x�۞���ؚ8�m��'�����@� X �<5�T�*�qE:!�. /�*uqF�'����S�/���7�[uB�-!��;\X��ѕz������uc�gt�W7�{zB#n��jI���z7���Q�x���=y�
���Oe�vv�`8����hgn]e�S)�s{ny��=L�γ�V2�����д��Kj�62����
�ά��w��q�����&�v�-����c��]�:쾸�6yNa�=�]n�{���w��:��.M�/l�Ƀ��d��a0���#�;�9�I�Z��C�Z��� ��8��?����Ɓ�
���dx�mE$N= ����""c虋�y.0�� ����;܌����Brh�)�wt���ֽ ��4�)d�)y$�;���@>l�@�b]]sgr�IbI�qĢq��4^���٠z����Қ^U�4f�ND�dy����ڴ���βo7�������79��{l*�919RH��q�����@��M��4^��]����6���f��I�~��P<0@�z��E@ |q� ������[^���^�k�V�E �"�7޲�/Z�/Z�^������s$m�ƛp�9zנyzנz����YM݇#%ɑ����Ǡyzנ}��ުS@�����ֿ�߿������-�Y
�q�5ٮ�R���9�"nL�����s�ݎ;VƖ5嶺�24�߬�h���9zנyzנwQK$qE#m�r�@�����ֽ ��4^�׉u%�'1��4�ګH�6���͵����Hjb��X%X�`w^���UWڪC�dfA ��JE�8�N= ��4^��;�S@��^���NH�mLM�& 6<���@>l�@�b뫾������ 6�
f
".�;M�Y��;eף�BR���lu�ծ9Mq)��+�I�7���Ɓ�ֽ ��4^���ʕ���"m�lm�@��^�}m��Jh�)�{��d�26A�I"���٠z�����M�Z����Й#"R7I4^��O��{9$����$�O���EH����?
蠾����I=����w\R86��	!�wt���ֽ ��4^��/�G���F9 �(DBsd��m^9Ԗ�b��ik]a+oZ5��U��=�o��sdNH�NC�9u�@>��ץ:&f?P6�ָ��P�!Z���^u zI�� �m��'PvX�p�D�jbm�&��ҚwJh�k���@��+s"�C�l]�;u�ڂ����& 6<� �\�\�L�&�cM�h�k�?DE}����q�n�f��DE�DI$0�1�X� ���73�.�ɛ�W�@��#��ݷhM`4������q$l�Y���"L1�>Ӽ<��w�ጰg�����Ogl0q�6�v�ɬ�ٞ���˵�w75�5t��lx���Y�
݅�7+��8�h��v�v��5��{A�����q�κ�+��K�[o7=���X��9-��e�����S�K��y;gw/	��: 49y]{dvxx��?����t�n2N5��Ts�%��q=nM\�k����s����YP�G�����=zS@��O|��]zx���L��)�RMץ4��9zנ[f��E+���o��wJh�k���@��M$�52'"�7!�r��@>��ץ4��;�)"�I�iǠ[f��ҚwJh�k�m�������~�RC�#c�[t��+�gU�/\��v��`����Z!�
�,�j�&�&<i����Ɓ�YM��z��z��V�E �&$�&�{���b����$	0D�@Oʇ뺪�3�x��&�1��l��J�1��p�9zנ[f��ҚwJh�;.LJ(&�$R=�U�w,y�0�L�6�n���V�!X��U�)%�|�3 鉉��q�
���[f��ꣳ"p�7 ��^�lq�گb�$�Y�����H5��]�;�l�r8��6��	!�wt���ֽ ��4^��>�KNcS"rF�q���t�DD��ܰ��7u3@�t�ND�q4��}m����r~jz�!�'�? ��]��rIW~�����p�D�j!���Jh�)�r��@>���ثS$�`�Ĕ��4��9zנ[f��Қ^�I�0#	�,�� &�ܴc�:���򱶘��3�z󫴼֑�<<��,�M�lm�@��^�}m��Jh�)�{��%ɉE�9���՝131F�\`����w�T=��P�������7�� �����z��h�R�����I���1
���>w��k���T�kQ(�y���ı% 9��dr/Z���4^��>��;������J�c��fL\��lއ�<�x��)Y'g�̎����n�$�Cp�r(��4��}�f��Қ�Қ/Z�s�U#�'wB�������艕7gͮ0O����h��Z�$�&	Lm�@�y����� 6<� ��9�Q�#�'��h�k����=zSA�b��i�}�v"\��PlNF�� �sA��͓��������?v�a��c;-4��闛���ݡ�����-�Ź����D*O.����Y�w˧mV�q8az��ݵ��=q;��bh{<⓺�98ώ�w�8��Y9��NGi䜶�L�j�v#c�\by��'Pe�h���+|\��֭�z��k������9�����ڷM����mۺw�M�H�Y�Ɨ�`y��n�n.p�ᴐ�$�r���)�@9�*�L���Y��r��[��;g��u��Ԓ�x�F�+]�K��p��zy1���-���1�2��3�7�@>l�@nb�)\RH�x��Hh�)�r��@>��ץ5�fbG�IbJ@s#r)j�# ��� ?6��3U���~4+S�D�E$���8��l�=zS@��M��zWZ�(G%U�Ң�%�|�3 �m��u�נ[f��P�c�I��E2B�Ce�C�2u������v�z���vm8�;���Ք�$X90JcnwJh�k���@��M �\�\�)iI����'V�ת��U�^`l��k� ;�S@�vw�,��br7#�����ۺ�q��@>9:�z;ɔfHȣ��RMץ4��9zנ[f��E+�A�o�I�S0��w�����X�S0��|~���J-0l���tmr�]�t��<ok�q���̎�5X��^q�Kf�n���2�x	���@�bc�r��py���!̐�D�Ɯz��o��g�@��Ɓ�ֽ���#�&ڈm9&��ҚwJi��g�0���Ǝ�z�� �p���,�|F/�|ROa�J0`��h�F��ZZ�6#)T��Oڎx�JƝ %�Fa
.!�1aLaq��\� C0$�q*��q��
1���3S�?(ꑄHBI���KE*T�I"�c�H��U��c �5�u DIIP�U�H!��H���$��kFH�#R֍XX�`D�5�`A! ��PX1 ��I�B�	�S�j�$Q_>X j���W�Q�QU� ~Q?���b��P��wo�Q3��,�11Tw[��	%PZQUJ*��""�y� �{��g��w,?E}37�k� ��ꮅt��uv���Ia�[�y�Twr���o5� �_�����g����0�7.]�4�y�Wj�%s�v�{c�ܔs��䣄�������׳ ��EYI+����A������z"P:����{R��T����c� y����&~{��UB���R�T�$����.с��wg��D;����w,:b"�y�0��URPZ�v�����Ř~��^t�EP}��y$�P>��~�I������*E�����_x�L��Q޶_ �		%WWV� �_wr�Ѽ��7u3 ��ڶ��������l8:������A��K�v+u��]�6���݀�;�̘=��S7Zh�4̹��O"X�%����br%�bX�}�;8�D�,K���"X�%�|�{�O"X�%����d�sv3e�K���,K������%�bX7��59ı,K�{��yı,O��ىȖ%�bSޝ��ۛ�r�ip�͜O"X�%�}�sS�,Kľw��'�,K��}����bX�'�}��'�?eL�bt�v�ɹ�e�s-��ND�,Kę��߷��Kı;;��'"X�U!�2'{�~�O"X�%�~��4� Gșı;����ɚf�۹�6˻�O"X�z#"w���ND�,K��?N'��ș�2��3S�3*dLʙ�{��{�L������w{���}s��:C�;�t��!��銵E?��y��C�&�KJe����l����og6;���n�&f��(q[Sd�mtm�8x��'�rNzѮz9v��.�36�z��N�M�
=f��-/F#�X�h�����u�%�K.��be�t��
�<���v��}i�6��E������gI$�t�r;=y�̙�,�ݖi̹���A9��^M�OY`]Ym�;�20�yॵEn[0/Vn	�w:�a�I]Xf�������&eL��S���Ӊ�2&eL�~���Lʙ2�y��x��S"fTȟm����Lʙ2���w=�n왦�n������ڙ2�A�w�jr&eL��S<�{�O}��3*dO��r�r&eL��S���2&eL��ܙ�	uf�F��}��{��S��???7��2&eL����\ND̩�3*}��vq=��D̩�o�᚜��S"b{���~&:�@��Q��w���{��D�n�.'"fTș�>��;8��S"fT�7���ND̩�3*g��w�粒��=��~7~.�kv[��G�"fTș�>��;8��S"fT�7���ND̩�3*g��w��2&eL����\ND̩�3*w���&�3$��nŋ�ێ\�+���e�vԷM�����Kۗ�ùti��m����s��x�7���ND̩�3*g��w��2&eL����\ND̩�3*}��vq=���r��{�����ҖT����&eL��S<�{�O}�����H)�"��by�L�ݻ�.'"fTș�>����'��ș�2��3S�?*n�lLʝ�t���e�n���.��=��D̩�;�e��Lʙ2��}�g�jd 7jl��3S�3*dLʙ��߷��2&eL�Ӷ�V��������=��)���~��2&eL�~���Lʙ2�y��x��S"fTȟm����Lʙ2���w=�n왦�n������ڙ2�A�w�jr&eL��S<�{�O}��3*dO��r�r&eL��S���2&eL��'���q���m�&fez��qtܜi��YӎΤ�Dr��F�ץ��6��Z�P�#s{��ܧ���=�����|��S"fTș3����Lʙ2��}�g�jdLʙ��3S�3*dL����}����M�e�����w�O&w�����S"fT����{�L��S ���jr&eL��S<�{�O}�;ܧ�������Mn�pt-M��&eL��S���2&eL�{��ș��$IEW��
!�&h���,O}��}���jdLʙ&}��ND̩�3*a�N��m�ٹs4�ff�'��ș�2�xf�"fTș�3�����ڙ2�Dɝ��"fTș�>��;8��S"fTȘC��~[JYzh+����)�w�Os�{��{�L��S!���ٚ�D̩�3*w����{�L��S ���jr"��{��>��<�7�QWS���v�kha{CՍ�l��囓5�,���p���r�t˦�͙�]��{�L��,��jr%�bX�}�;8�D�,K��ND�,K���x�D�,K��/y�wfnm�������Kı>��vq<�bX�{���bX�%���<�bX��{���bX�'��w<�n�f����w7gȖ%�`���Ȗ%�b_;��Ȗ%�`����Ȗ%�b}����yı,K�rwM�rn���ˆ\�S�,Kľw��'�,K���sS�,K������%�`p_�{��jr%�bX����3����s2홗7w��Kİo{���Kı>��vq<�bX�{���bX�%���<�bX�%��;vۂ���n�ls�ؽ<�k(]�
�>[��f���s��Yu�[��U��%�bX�}�;8�D�,K��ND�,K���x�D�,K����Ȗ%�bSޝ��ۛ�r�ip�͜O"X�%�����"X�%�|�{�O"X�%�g{���Kı>��vq<�bX�%!��wd�˲��ݷt��Kı/��w��Kı,�{���bX�'�}��'�,K��{�S�,K����̽�L�m�ٛe��'�,Kĳ���r%�bX�}�;8�D�,K��ND�,�2&{����y����ow�~������&*��D�,K��gȖ%�`���Ȗ%�b_;��Ȗ%�bY��u9ı,O � Q��s	�i7i;6s��^ջc%rb�����/ݜ�n�	ӓp�2�*�bv�ZQۗ�ˮݵx/h�,���T;<MC먝�7`�7O��;z�L$�������'K�^�#�p�h��=�J�ិ-�I#�N0��#�p!���ɻn�m๪I��l�6a�1[*[��u����箱�mm�@._[�h9r5S���oG�gd��(��������{�<�/S��pE�F���%b|��W�������ט��쫹�ykl�nn�����}ı,߻�S�,Kľw��'�,Kĳ��� <��,K��?N'�,KĿ~��M�黻��nsMND�,K���x�D�,K����Ȗ%�b}����yı,��59ı,O���3����s2홗7w��Kı,�{���bX�'�}��'�,K��{�S�,Kľw��'�,K���ٙ4�ݤ��-ۙ����bY�D�{����%�bX?�~�Ȗ%�b^���Ȗ%�%�g{���Kı)��e���ܹ�fsgȖ%�`���Ȗ%�b^���Ȗ%�bY��u9ı,N��;8�D�,K�ӹ�\>VW�tsum����lhqt)h*�u�5�3g�N������k8��.�Zs��Kı/}�w��Kı,�{���bX�'~���O"X�%�����"X�%����;&�tۻ�m�wx�D�,K�����x��D
z'*& ��X�^���"��M�bg~瓉�Kİ}�xjr%�bX������$KRĳ����Ϙ�M��1U��{��7��߾�gȖ%�`���Ȗ?�R"_�~��O"X�%�g�߷S�,K��ޝ�6[�&i���wsvq<�bX�{���bX�%���<�bX�%��wS�,K�"~�|�8�G��7������ۣU4C��{��,KĽ���'�,K����~�O"X�%�������%�bX=�xjs{��7��������:A�a6���GV��O��7��ф+mh��r��ޭ7g��������i�V�V�������oq�;���Kı;����yı,��59ı,K�{��yı,���ƪ;,���}����ow����g�~�L�`�����"X�%�}���<�bX�%��wS�,Kħ���,�ٹs6�2��'�,K��{�S�,KĽ���'�,|>PO���"r%��n�"X�%���s���Kı)�û&�]�����"X�P�{�{�O"X�%�g{���Kı;����yı,��59ı,O���t�.�wtͶ��Ȗ%�bY��u9ı,N��;8�D�,K��ND�,K���x�D�,K�e��sf��އu���گb��	�m�5���H4�ֻ�6�^a�)��K�mew��g��u����;8�D�,K��ND�,K���x�D�,K����Ȗ%�byӽ�m��n����6f��yı,��59
#ı/}�w��Kı,�{���bX�'~���O"X�!�����ˣ������}����b^���Ȗ%�bY��u9ı,N��;8�D�,K��ND�,K��������-*�eZ��7���{�K;��"X�%�߾�gȖ%�`���Ȗ%��QP��U@��*=9�Ns��x�D�,K��ffٛ�d��l����ND�,K�}��'�,K��{�S�,KĽ���'�,Kĳ���r%�bX�����o�#��JI�J�뎷NݜB�����W^L���i��6���V�E��6����bX�{�:��bX�%���<�bX�%��wS�,K���s���Kı)�û&�]�����"X�%�{�{�O!�Q#�2%�g�߷S�,K������yı,��u9ı,O���L:i��nn�����yı,K;��"X�%�߾�gȖ?��`�q��Kı/���c�1D�Llm��%j�	\]Ի��Ȗ%���{����%�bX?�~�Ȗ%�b^���Ȗ%���v&������Kı>�?���n�ۦ���͙�8�D�,K��ND�,K�������%�bX�~��u9ı,N��;8�D�,K!깴��A�Lep!�F�)��+�/tdR�#&a�1"�n�h��	K����p��
�[P+ ��Q���7�i�T�@+�XƮH�A���ʠB��
J�ԀHE�����XJ@�(A� ,e]�tS~T���!"V%�Z
Vi
����V���R$�0i��@| �#Q�H $d�!"B����$�J2��HC`�ʀ`��Q�	"�bD�� �jBE�R)X��/΃,i�T0&8Q�1\IXP�L`5���!Wp�C�c�1�ĉI�K��c2����f�8Ǝ1d`EdH��,8�`(OO/���L��L˹�rf�5��m �m���9�����0���ԁ5�mQ�����n��`��/��h;<q���m��n���f�#�^n�V)�HJ����UU�C�m�h��*��VU�=��x捒�9�\=KOic�+�e�۵�ntoj�;G25��u��+�0�#��UUr�8����\k�vɎ�^u�[<c����u�7c�:e��׫m�۱����VC4K��[c]lq���'WX���l���7;-[�G��X�zv)� ll���J3٘6�K�lj��]�X��;=Wt���CP9��9��F��76���[Y��ܰt����r���i�Y��Ck�H�nk����]�����F����xй��/����������.{7���tn�;����٥e5���[[�&It�9e��/,�ag�	9���<���x���j�������a�²�T��'m��'���ۡ�Z��(�p8�;
!=�v�����g��7k��n���a���i������v
������J�uBҁ�۳]#�,F��6qЗ�7m�F�8������3�1��AAң6���۔Kj� ����v�vW��~�p�Eћ��f;N6�J��-S�wfpøhlѝ�Om����\�����N-�7T��<�6�fզ��FzÎ�g�V;�V�Wu����#9���d��!�H��)�=*�d�zYŒW=15M+[@Z��Z5��N�y�Bm� �[�Z���ӥ�T���f�۔��ա�V��������%U:݊�iY�vpy��e�5ɵ�g7JEQ<����]�P����2�x]�H'������ʮ�Qg�v՗]:T�۝����X�у4��4�@O/��b���^��7&�e�X���Y��v�y�g9:1�����9�"�ۀB����mC��[�T<�s�TJ-�ní��NSi��m�L�5e�0�)&��P�S�)��j���� >�Ojj�}@ ��7�7nf�sf�0ˆ�f�%�Gɺ��ƞ��㜜�=�KI�Zt�\�d�m!����^͠ι���R�88����u��3ge�'r��� ��\ź�E�vc&��3��,��u�Z;=�2��v��۞I;l{A���1�M�8�Z�5�ά� r�'
/Y95Z�y� �&3����=t�����gn�,=����rs��k�W:�]��7nW Fs�{���_<�8�SmXy5����vr;�p������In0����w��>%�8®�s�w�,KĿ~��'�,Kĳ���r%�bX���vp?3ؙİ~��}�oq������~���a�Q��WȖ%�bY��u9�A��bX�߿s�q<�bX����ND�,K���x�D�&TȖi�3l���3$�ffn�"X�%�������%�bX=�x�r%��Dȗ�߿oȖ%�bY�����Kı)��e����̹�fsgȖ%�����:��bX�%������%�bX�w��ND�,�2'���Ӊ�Kı)߬?l˦m�77m�u9ı,K�{��yı,?r~��u<�bX�'����Ȗ%�`���Ȗ%�b|{���õ�#�i�.9�Y�W#gh{f�E+������ӓlk��^;�y>雵���bX�%�g�߷S�,K���s���Kİ{����Kı/}�w����{��7�����5����*�܉bX�'~���O!��W����j�yȖ���ND�,K�����<�bX�%��wS�?�r��q����~�� +E�T�������x�,߿q��Kı/}�w��Kı,�{���bX�'~���O"X�������u5�7�w��ou��2&~����yı,K?~����bX�'~���O"X�����`�z�ﷸ��{����o����*�
��O"X�%�g{���Kı;����yı,��u9ı,K�{������{��7��?��BP���h�ւ(=z�"g[�v�U��N;7�7.������ILa1D�L=�s��Kİ{����Kı/}�w��
3ؙı,����r%�bX����l.��˙�a�6q<�bX�{�:��bX�%���<�bX�%��wS�,K���s���O��S"X�����e�6����bX�%������%�bX�w��ND��x�� 0ț�y��'�,K����Ȗ%�b}���xf�ݳl��'�,K?"�2&O߿n�"X�%�������%�bX=�x�r%�`D%��{�ND$S�|\�nn��ٙ�2K��$�H�{�ڜ�H��}��bX�%��{�8�D�,K����Ȗ%�b^��;0۷v���r[�%l�˵v���|��V�]�Hv	�ޚ6Sq�K��ݛt��ݹ�7gȖ%�`���Ȗ%�bw���'�,Kĳ���r%�bX���vq<�bX�%��;�-��wwwr�nk�Ȗ%�by���'�,Kĳ���r%�bX�}�;8�D�,K��ND�,K��p���sv�wm�w7��Kı,�{���bX�'�}��'�,K��{�S�,K���O"X�%��w�3l���3$�ffn�"X�%���s���Kİ{����Kı<�{�Ȗ%���@ =+�����u9ı,J{����]ݹ�3l�.l�yı,��u9ı,K�{��yı,K;��"X�%���s���K�q����Ϛ� [P���<\�9v�
T��c1�Tɭ��\8��Nس�O;���\�p�ݷu��Kı/��w��Kı,�{���bX�'�}��'�,K��{�S�,K��߬)����͓d����%�bX�w��NC�ș�������%�bX?�~�Ȗ%�b_;��Ȗ%�b|O���3vmɹ�2K����bX�'�}��'�,K��{�S�,Kľw��Ȗ%�bY��u9ı,O���mݛt����ۛ���Kİ{����Kı/�����%�bX�w��ND�,K�~�gȖ%�b_{���ۻ7wwn�2溜�bX�%���<�bX��?�����u=�bX�'�߹�8�D�,K��ND�,K�<*�P{ٗ�ݗsn�n�,�b�<ݮ9��圸r��K:�y����M�:'�5�{=�����n�A�^���k�s�K٦qve��GU�W	��n�ݎ�.u�1��K�vSl�\[�=��n�r%��:�����������j�:^pf8�#�G]q�$n��r�y:���]��j�Z�ca�v9�o7e�\�ld#��.���/�6-�c���|y������ww�W�)�w2�/M36�p�$�9c0�,nц�]�{v� r�{��� {����g����R�F�����{��7�����W��,K������%�bX=�x����&ı,K������%�bX?���.���{\*�{���{��7������O!�*G"dK���u9ı,K�~�'�,Kĳ���r'�Q��{���߸��,&F�{���o%����:��bX�%�wx�D��2&D���۩Ȗ%�bw����yı,JC���]6f���bY�D�w��<�bX�%��~�ND�,KϾ�gȖ%�`���Ȗ%�bw߬)����͓d����%�bX�w��ND�,KϾ�gȖ%�bw��'"X�%�|�����7���{�?5��r�t�\��bz3j�L=�{T�ϕ�a��n�a9ԑ����n��nm̳$���Ȗ%�by����yı,N��6D�Kı/����yı,K;��"X�%�ߧ{��wf�7wws&���yı,N��6D�=�:؛Ŀ}�w��Kı,�{���bX�'����O" �S7�������`+������oq��%�{�oȖ%�bY��u9ı,O;�;8�D�,K���9Ǎ�7����{�*�eV��7��bX�w��ND�,K����'�,K��{�dND�,�L���������7���w�?oܺ�e�p�[�Ȗ%�bw�����Kİ�������ȞD�,K������Kı,�{���bX�'�w��0ܹ�&�+�S�6]�ЮЯ[��;`�t�l���^�kg�w6�u��QV>�7���{�N��6D�Kı/����yı,K;��"X�%��w��'�,KĤ;�ΚL�e�wI�l�Ȗ%�b_�����%�bX�w��ND�,K��ݼO"X�%����Ȝ�bX�'}�0����6[��O"X�%�g{���Kı<�����%�?"M��;��'"X�%�~���Ȗ%�b|O��f��nf��2K����bX�'�߻x�D�,K���9ı,K��wx�D�,Ȓɋ;�)�&(��b��gw�UI
�$��d�ݼO"X�%����Ȝ�bX�%�߻�O"X�%�g{���Kı<�����%�bX>�woL�ݲ����n\c����7u��Ϣć�h�k�s���#̈%��5��$�}=�{��Y�{�w��Kı,�{���bX�'�߻x�D�,K���9ı,{���{�-*���_{���oq��K;��"X�%��w��'�,K��{�dND�,K����'�?9S#��~~����e�p�U��{��7����׉�Kı;����,KĿ{�w��Kı,�{���bX�%>���6]ݹ�3s.ff�'�,K?2'�߼6D�Kı/~���yı,K;��"X�U�AS���ȝ��?^'�,KĤ?~��]6f�L�dND�,K����'�,Kĳ���r%�bX�w~��yı,N��6D�Kı?/������rYJũ��h���%��8��<;���ڰNu�αr,��ݫ�%���ؖ%�bY�����Kı<�����%�bX��xl�Ȗ%�b_�����%�bX�����f�sfe�%��ND�,K��ݼO"X�%����Ȝ�bX�%�wx�D�,K����ȟ�*dK�g��m�t��3773n��'�,K�����9ı,K�~��<�c�!�2%��~�ND�,K���׉�Kı/����m�ۻ����f�"r%�bX������%�bX�w��ND�,K�oݼO"X�%����Ȝ�bX�'���ٳsn�\͓33wx�D�,K����Ȗ%�bw�����Kı;����,KĽ���'�,K��E ����~lZ�K�u�"��֦�.�X�;Z�vQ�㫓m���utgSp۶�c�v#��v.ݶ��Y�Lo������Ao]���E�gݜ��q{T)Ƭ8����3�M�h�=���������Χ'�=8.��O�3�]lQWu�u�;��"�k�g6�;�lY��cu�p4f�ޓ�Wm��v�I�!]�o�}c}�i�ͳ7&k����y�w,�]�٨�ٷk=�z{N����.�ӥ�L�i�9w:�9��A��.�v^�
�^���7��������%�bX��xl�Ȗ%�b^���Ȗ%�bY��u9ı,J}�izl��s.f�[��x�D�,K���9ı,K�{��yı,K;��"X�%�߷��'�,KĤ;��e�fa��f"r%�bX������%�bX�w��ND�,K�oݼO"X�%����Ȝ�bX�'��I'L2�nf�-��'�,Kĳ���r%�bX���vq<�bX�'{�"r%�`,ș��߷��Kı:N��3Lݛsfe�%��ND�,K��gȖ%�bw��'"X�%�|�{�O"X�%�g{���Kı?*~���3���nf���3���v�3tǖ�H�j��4C�����Z7��>��X+�YfXk=����oq�߿��l�Ȗ%�b_;��Ȗ%�bY��u9ı,O����O"X�%���~V	���3u����7���{���w��9�5؛ĳ���r%�bX�����yı,N��6D�K�q�����?�ġ@�W�����bX�w��ND�,K��gȖ%�bw��'"X�%�|�{�O"X���#�[����
�^ﷸ�,K��gȖ%�bw��'"X�%�|�{�O"X�%�g{���Kı)߻K�nnL�����͜O"X�%����Ȝ�bX�%���<�bX�%��wS�,K������%��{��?����9|ԇ&��o�]������]�kE#mz�`�{4���m�:��u�3͓0��,Kľw��'�,Kĳ���r%�bX�}�;8�{"X�'�߸l�Ȗ%�bt�d��/��nٲ\��yı,K;��"X�%���s���Kı;����,Kľw��'�,K���娴�V��,)$�0��b��&7w��%�bX��xl�Ȗ<;�S�A�1!��!'��y��
�8�!,=
�|�He���`��s��PhLT�`�(��u ARP �`�BX�ƪZ��C��H�9>Z���R0`��@`�Q�� 5�8���� x��x�T4Tנ��Ӏ A@��� �E�P���DpE��ʣUD�u<O_�T�b{��~�'�,Kĳﻺ��bX�'��vۺLݗ77snn�'�,K��{�dND�,K���x�D�,K����Ȗ%�b}��2c�1D�LW�ƑT�V�ZWwFi�'"X�%�|�{�O"X�%�g{���Kı>��vq<�bX�'{�"r%�bX����M�pۛr�sDpk����O�fcrmHl��24���g]N2JDZiVl(��������d����r%�bX�}�;8�D�,K���9ı,K�{��yı.�/�K���k��W���7���'�}��'�,K��{�dND�,K���x�D�,K����Ȗ%�bS�v���nK33w-˛8�D�,K���9ı,K�{��y�� �"dK?~����bX�'{�~�O"X�%�Hw�4˦���٘l�Ȗ%�b_;��Ȗ%�bY��u9ı,O����O"X�T�U���Ȝ�bX�'ǿr�ݗM�ݳd����%�bX�w��ND�,K��gȖ%�bw��'"X�%�|�{�O"X�%��2���3.ݛ����v�Rv������A��Y�N�Ln���rq���˓k4�=�Ou��=�x�����%�bX��xl�Ȗ%�b_;��Ȗ%�bY��u9ı,O>;��vLݗw7snn�'�,K��{�dND�,K���x�D�-�����4JIq��C� �����m��� ��*B����*����DLU}�� m�4�M ��4��Ss$��a0m�&��ҚwL��}m���l�_�dY<��'ٽ�4��Ď&�g���pORhװ��պl��p��n�k5(=n�s���x�:y��*�]Ub�N��/V��۫�Q�x�k�^�!��gZ�·�-{�&�;Zݜ-�����b�;it&C9��7"ݷ���;t���������G�����Y񇶈�}�g	���Gn�g��C���l���r����x �a�|�hmg���Ϝ�s����^o��.���v����U��K7�gghp�nY-3s֎L�y�����ʜ^�F�ۑ�Ӈ��3�[f�}m�wJh\�rcS �)�C@=$��& yo*Z�"�"S$�"rh�٠wt����)�[f����u�ndN��� yo*�L@�bΦX��jA�$qI��S@>�� ��4��-t��#$N6���θ`����h�ƶ���÷��J\b۶���H%$�H�m�̆�}m���h�)�wt�h]j���6H�s7w�I�{���x@ §ʕE���;��� ~�0���?m�N�$���(.��X�L�7uC0ꣷ�`�~�4;�����6�i4�طT1 ?�X�v�u=�f C��#�`�A<R!���_[4�l�/t����)�vy�d�Mly'�d��l���Wi��!3vk7E�x��˺�m'�w�mVBUJIE*��� �{� {���gO���`5�vZ��
������7�@6�&Ɉ�L_]���URE�E���I# m�� ͮJ��P��	" �.�&���$@�_��{?o���'�ݟ�@>�Yܑ7��9���f�~m��`t��6�8�_¤$�U�+���I`���:&'��?m����f�_uC#hP#k�hqe�ײK�6�8�Z\�Im�]j��H��$�	�m�4�)�wt�h���1?���`7�Ғ�awi]Uգ ��Ή�����X�w,�Jh\�r`�A<R!���_Z��ma�3Uͮ0ڎ0��S���$��V��&=w��������}��vrOE4*D`N
꣊s���y$���f��m͙��d�K {��LLKo#���� ?6��������$Hr��F�(�V��L;<�i�OFD.��&�չ�FWq�}�������S#���m����f�}m�����A7$M�#md4��Έ�����`�� ���zf&".����	\$�Uڸ���I`��Z��;�e4�٠}�*��$�`���I`t��DW7�`�`����31U�w, ����R������рn�`������X�NrI�%"��S�߿{I����3s6I��hb��hYۧ�4t�7�8�T��6����Mԗ�vji]�yd�6�ԣ��q��XG��N^I�y�]���#. ۞����}k��ݶ'Kp�d�t�0lA������s2k�gn�b�`k���$nJ���r��s�
Ϋu)^��㵠7֣γ%ʹs���gq���tki�p��E3��1�<lBy�����r����F�<Dӌ�NrMy؏kS�N���r�Ц�eلێ��қ�LP������p�, ��X�L�;�e4�vW$Jdn)�JI�V�L�D�bfb.�w/w(���tLLMP��vZ��
�UںAV�ͮ4�M ��h�٠}r�RX�$���������G�ܰ�m`tD�Esy���v���j�,�X 	�b ������$�Q_�w�l�e�vf�\%�3C3btܬn��n÷F��K��y��K7,���޾d��J��T]�]$� �{� {���gLO���`>U�v�$�.�Awv����{wUu�i�+� ��@[f��ă-��~�D�BND�N�+� M������J��8PZ�U´p������wr�/>�C�b��~4�r$~�ҙ�B*�, ��X����ڎ0���-jX۟�$���C�`�Ȇ՞�{h������9h:�tq�h"�_�w��}�p�22r|���wt�h��@>���X��q��$qI���)��� ��4Ϫ�ؑ����M����T�# >���kL~�&b	��&b��&e��m.0�P�]�ؕŤ���E��i,U}�� m�0�P�L�EW�ܰ�*�P�V�`�rM��4�M ��4�l�=m̓���)���m��n�S���8;\�9MY�^ؘ|5��a��!���ֆP��$ӆ���)�[f�}m�wJh\�r`�A<�y �ֳ�v�y`ܼ`�����*�L�E2rh�٠wt����)����إs�N&�P�@���� 	�bvuu�un��:�T�#>��o$�t�{��7vݵi*Ui�f陘��������@�Қ�(��Q�܉F�bN �r�L7����YmřѮ�5˺ѵ�ݔy��`d�9�H�Rd4�٠[f�{�4�M��U�����jI��k:bf#�g�����x��k=115Gϗ]](I+���T]դ�mq�n�a�;{� }�� #u�S���**�*���`z&&�y`or�͵���� ���#�AjW
�]�l��=$�o �m�A-��C�XyQ1��ybD"H��Dg�l1�!�,"Ő@�(�� ��0J0%&�z��<0��X�`��z-�є	RST�@�(��(�F�׈��xƎ��C��dTI�N��@��%%IkT�4\bL�15cQ��A�1_!<Ex��>�:e$�\c���!c��F8+Ub!؍ �Vb$�",�,H$�a(���"Om�F$�J��%�d�0 PJ�P!D��hA�Bcz�A�D�#$$�W�6$e�#�1����`�� �° 	  #C$!0`� ���!!$$	 ��T�0�Qecڥ@p`�ۋ�`�@��5��	�cBN���k��۲�:���U;���msa͂�/n��A�%`v�ƛ`A�bA�7.��1J��;�IW�3�uk�M�򫄇���r�X;�/Ikw�=�m��+��SU(��uʵ�U!��J�+�m����H�:�b�V�\v�Ӭs�拶e���a!���l���ܢ��jigu�`c��'5�pˆ�;$${��=�k�#��u��Ln/;c-C.���Aw�d��9E3&��˵J���њ�� psi�'�WK���q���T:�`8�-�7jMD�r˫lxEXpqsI����&���ܑ�ַ]z�c�F�ٺ��ls���s��c=���B�L�M#xl�tM pu�)��a4���r�[������m�&Hn�����ãh�����`�ٞeq�g��Z�^7��y�û'l�rBewїX5����1v��#�zM����5�;LeLI�v\g�Ke��3�i�>��$�˝�2�x�`6�HN��@`�n.Y��׋E��':ul��cN��͹^�Ҽ�g�u\n0On	�Lۯ6�=��X�S�[�c�$�4�`���ۣn��j�����㒪��M����-�;�v�	�p�ݫ�ʵá���ۃs��lq�Q��Z�ݵe!\��d}dv�Z-�:��ӊw��nq&k�)���.C���uNXm�s��'��b���]��*�U��胳���M�����S�)��+<�U���ێ�fA)k�@�%p`�3[ 4v�#�F�n���lɳ�ݝq���p�JZv��oKt�j�w,��
�Z�;j�dz|�ScH�����-Ʒ<֘� dٴr<�r��lt�ZMc�ʼ�g��^w]�ɺ� 9X�[Npo@�$�K��}���,��{d���iN&�o�,���]�cF�uO+/,�10����i֋��.�}t��@ ��<OU^���W� |�PN �G��v��lݷ6Zd3I����ɩ'�Ű���NK��q��)ÝpԦ�sv�8��#{i1��0��q�}{q��N���n;z��ls6�nx�۶P�v����+���k.z�v�,�ݎ{A's���WXAN`ʼ �v&=������s٣�4��c�^9��f�n��gn+tr�ۇZ��]��`-�m˽]��]��j\�ۊ5�ncd�p�C�p�=;������m�@Q4]us�����'�A�<��|38[�6k[pV��{���w�At�u�����=��wT3�"c��ܰ���98ۍ@NM�Jh�1� �m`��Ή���>��ʪ�$���D��4l�ƀ_[4�l�.�f�X�V��jĕ%IB0:f"&*���wr�7u3�"bb�y`�������cm�&�}m���;�e4�٠ݖ4 S#��5��9����)!��1(�Q��-���q������%�J1�j�m��>�� 	�b ��79\���۳n��r��I>��;9X�����DDOOd�"bv�{>X ��X�L��ʑra!�8�4�٠V�1Uͮ0ڎ0��W�R�Є�V��j���sk�wT3�U�ܰ�)u���Z��t��,�`-��? v�, ��X����ȴ+R��unӹ=sq[ʒ6�2�i��E�ݕ]΄�k��N���Zɉ��f ?�X���3�=ܼ`�=���j�+T�%��k=A�w,�\`����\u򪲒WWj���X�w,�a�1!�&&�B"����O��4�9$�{����i�](I+����ZK�bf"��� m�� ͬ ��X��p�+Wb��Uwh�7uC0Ev�/�w~���*���do�F�,�cS.7�6Z�s$��b���^h���t����d�yd�B	�p�h��@>���Jh�2�x�Ȣ!&A�&�zI��A �ʂ �&/˻��	���98ۍ@NM���wt�a�3>����X�����MUR��RI!Z)#���� ;{� ~m�A�U( <�<�}�g$��r!�Q�E"�!����m��`���LD�6WWb�\̀]��t��:"7kjd�ٶLf�]�֎��s&�iT�
�W�m�����^�M��S@/���ei��H��Ae�W�=��虘��j8�����>Vנ�R.D䉑9�p@6�&ɈrI�o �+fT��	'��o!��� ��4����m�q�=+��T��!(Gy���& #yo*l������ק�d�d�����f�4�wq�S���7���Y3������+w,m����s�u��;�t�hݳ�k���t��G��]���t��J;�`��-�K�=���b�s���n��gC�����]���+m��s��e�ay�O+&�.1�V��!N�9�<q�h�
�.�n�1��^%э�q�N)���q�Ƭ��pװۖI%�ݛ\ɒL�a�}���])�Y�wi�6������xL�q��g"�Փ��μ���uO�0��a��n�`��� �mt��������*�Qv��I
�I�g�""�;{��wu�u3=15Gώ�TZ�J��*J�F v�,�6�3U�l@n즁��&�M$���ٟ��mz�g�@��M ��h[
��#��v ��+�޺�:&"y����|��@>����'1�)"��ɴ�Te�zb8׭V�'^��ʋ�g��]
�UiWV� ��� 6��ۿL�O�&'�u�� !�=Tz�p���1���U|��:���@6��315C�¸��J*Ҩ������~z��h�)����إs�RWv��j�:&&f��Հ6�}l�>Vנ}r�S���%#�,wS0������_�����������:ᒆW�s���qӗ��v^Gnm�IP\;zyh�v�N��R�2�ART�0���?Sn����f"bP[g�@��/ߣLRF�����h+]�o]`�����z&bb=131f���ZBV���]�x��Հn����(�� DN(�}>O}���f�����wQeȔqNA&�X����m��ܰ�m`z"��Հtu�ЂԪHH*р��舘����~�\`���l}n�SW������QN�������[�2e����p�X3�.��M�k]FZ�m�������L�7u3�3���=qJ��H�J�+�%x�L�鉊������`��y�����7��ʪ�]���UI]$`ܼ`���?Sn��L�?kB��T�X���$`tD�MW�ܰ��� �u3�LLʙ��I1! �S������~����e��̵WwwI,�6� ��L�4�� �\`��@/����(6I�`���8��z��I�&�m��斛�sr�إ՚� �m6@m9&�{�4���g虈��@}�� 5�Tt*�j�U�TU�p@6�l��=$�o �.��c�1v��=-J�	 �F y�� �M���f����lR�p�EZU
��K�bf"���y�0�L�����=�X��΄���һPRW�|�3 舘���DDww� s����w�}阘�&$�"&��_i6��"躧8�;&�{4G:z�Zv}rm���ѷ]�-��)��tQ����1��̮�*��T�������OW�1��Ps�'�[crΗ!=��˲�s�T�}�X3�X�!�^�Y���]M���F�8[��ɢ��m�rWCH��LZ��v]K�д�vM�1�'�;p���� pܡ��A�/kn�l�K�:�� 7��y�&��ٹr�al�nmm�V��1vyئ���ә�"�e���;8��	��RI��=z~4�h+k�D�D~�m�0����HV��Uj�F ~m��L�EQ�wu�����������ߟ���r2�*����?{�����`���?6�V���������4���١�3_wr��T��R�H���� �� 91 zI�o ��N��8y�q�����8WU�K��pj�]t���a�n����S�{���]�o�ٽ�ՅZ? |�� ~m����DLO��� �P��%iT(J����mf�>��%Dj4G���'}������ ~��zfbb�m��΄���һAI,[\`����""���, ��ߦ��v]�%1�)$�qHh������k�1鉈�������
��J�V��T�0~m`������7�� ����a�닪��wB�c�a��@t\�n����n9+;�8���8�����Z;��������Bp��m�����=zS@��M �[4��S������P]դ���g�"&}vwr����k >�UR�@��*;��o �Ɉ۵v��������<��"�(H� ]5�Q")F1�D D��H��H1"�"���p �Y��1�#�0
�$V1!�H�$H�m�rZy��Hć�A��Ą�� 
�=�1!1$�0BF0N��@{� A��� ����F���*t1@z)�A�
qG�>(��n������k��s �+eNp��jU$$h��L�D�""�}�Mץ4��/��ErH�"a%]ZX���DD�&f������� ;�����������2(��dͷT�֬sٻn˛Ӻ�GkfyI�uW:����)��ҚwJhz���f#���׀}���*�+UJ�IX�# m��1�I:���껪���ۑ	�'#�'��߿M�mz�Jh�)�Z�Z�ĜlQ��%��1__w^���`LD�@ ��#TW�Q�/���I�~�S����n,k���)�wt��oͬ�6� ��LF�����t]�%E��s#��2��{Y9���w6�v��/l\��Vnv������p�t�.��i�3g�O߿O��f��ץ4=r�r�Ii
­�6��&*���� �k�wt��|v �$hp�&���m����:bj�k� {ܰ��Uc����һPRW�陉���`�� oͬD���׀}���*�(����(T��n�f艊{ܿ�wu�=L�:fcd����qxu$UZ�v�A��4K;G0�Ј� ڱN^<pݻf��O[O9��]�B�
�{X���'ASfں� ��i��x�7	nݵ��\�Y��}�/Bq��ϗ�[ld}�R;)g�/[0!5]۞��g%�pf;v��
y��!n� n���m���͋f4�%-�m��΄9,���<��/5�t�����̹�RMɦې��|��\5L�q1��Cc��g��u�����ِ�qu�m���m�s��կ��)�U$� }�X�m���f�����,I��Ҍc�h+k�=�)�n�f ~��z#�voyW�%IZ���UQv���x�7u3EQ��X����yZ�\�FL"p"i�h��| �}�rI���@��9+թ�HH*р���tD}}����wJh�+0��Dҟ�dɑq�k٭���8��^ٸ������+aVs��ԡȱ�nM�mz��4���٠wg(�QĔ����H�wN�x
0V+����������4�M�mzݖ;�L���%
�0�L���âbj���[_���$�H��8�RC@>�f���w�}����33M�� �UZ*�ꕔZK �M��=1:�q���h�l���%1��"12D��l���)�;I=#��C��/:]Ω���J�9	lmőcr=�ҚwJh�mzf"c���׀mwt*�b�RXD�p�;�S@>�f���ҙ�35A��]��7I*TU� >}؀�$�AuUuYUuVs[� <�A �6(���Qp�i`tDDM}}�x���7u3�5_>�7�r��JG$j`�z��4���٠|��@��,v	E���o	���J��q[�I�؈�Sj���]wHO����w������H�drm�� ������wJhu.�'��E#�E$4����bbj���� m�0�L�D����+��B��tZ��I`Ww^���z&"&������`�V�%I8����zwJh�)�[f������? /U��2���x�ڳ��P]ZEݣ ����13�w/�}]�x�`���%�4gn�0=nF���$�,�jir�<',7Lv,�����HV�M����m`��x�zf"'�1Xwr�~��A?� �E�!�4������n�f ~m��g�ff�l����&�C�5 ��Ɓ�> �t�>]ߞ��e��9��)�'!�wt��~m��6��&"�y���p�J)R)!�[f����4����I4� !;Ӗ}�sK�F��u�4kf	�P�g� �K���첤Ln��|�m8\�c��q�hqή8�؝q��[Wh+Pv�m���ڣ����<���������n��s�]��p�4i�0�a��=�"�[b�}���\��vh<��L-m��"%뵱��ҺWv��Od��k�Lv'nЮι�����V�����6'1^aW�]����i/'\D=Wf�ݝ�c	���iU��cH���{���t%ɡ�!�8/���;�S@��M ��4���"����X�7#�;�S ��� ��X�m�t�EQ�}Vt"���@���`�� ~m�=311��y~�������ʕ��!��U��bb=3w�����z��L�;�S@��%��(<�ɠ|��@��M��4�l�;<�1�uX�G���#�3sگ��n�'��i����g^z�:���|��}�g]��o�g�@��M ��4���vX�4��ssw6������qT�#�a �ܰ��wS0�ǈ���P���"���h+k�;�S@���]�7J�UҊ�-YE��=>����z��^0�L�͵�o�X�Uj�]�j��.ҼwS0D�z&c��x�}�,�6� ?nՍ%�����ti��u�b8�n�9���8�]k�ˎ�j7e���d�(���!���4�l�>Vנwt��e�r1HA8Z
�`��Έ��>�����7zS@���\�O$x�D7&��$�ﷳ�5U1?�)��VS�*Ev /ȇAT�U>��^0��X�m*j��)*��PU���ַ�`�� ~����w�~�j�hUV�+�`���t��z"b"����^�� �u3 5ӶX�`��/l�y�Z�zRݹ���8�%Չ���M��s�
Ej�71LQV�m���ư�ۼ��Έ���@�\`���dMLMcI�4�����;�3 ?kk=33T=�g$��Uuuj��.Ҽ[\`����&b*��r�>�߿=��ˑ)"DRaM�@��NI'�w��'���rO�@�S�����#���������C�O����͗ �' ������wJh�)���?+˓]�������,��Z�Z]Fn+�e��u�N�&}��c�7V��J����wu�n�`��興�����@��?Ď!8���'���LwS0����ۼ陈�����x�#i�##��-��u�@�[^���M��$��9q8������U|���wu�n�`zbbf�yƁ������0i���@�[^��yo �<��)[*���Ue�H�� �[a�j��ԉ�� FB��$!��R,���р��B��+
R��pOEJ�H� �0#�iG� � u0% @Hߥ���<T���ph�����.h���(Fc(�2�F�)��.m0a4er\� &�� v�)4�HQ�X�Hb|,B	��X���|c�a�bPG� Tw=��[���n�[�f�Vv�� +V���.�����8.&�i�5Y�L����mCs^�K�@�k&�	�^��@����h��.z�����L�m�%IyU�e��������&D��s.�>��ny�vB���f�֪;]��=e���-�R%��}��Z {um�V��ä���6ۡ�a�q�8�.��Ц�NI#]s�T������C-�2�ZӞJ��{XɎW�)`zZ��l܉V�Gu�`�B�;6烀�n�cB��e4 �ۮ��lٳ�k�%\v��L�]m��P� ����N1���pm���z�՝��'5�I,7Լ�g�쫵V�9G$bW��gG��ۨ�kmټ�]��K���L�Xz����]ml/l�9���8�DԊz�[��m[��I����˵��ɩ��Bu��t׊���A���:;n��L֮3D��ȶ�zݺ;5e�\����X�]�2(�[��v�v#v�ħ<͸�i!<���hX*�qQ��u9;(�\vݣ&�S����i�$R���F�-ӡ.Rx.Uݻ\H\���j����{[\���-q%�^V��m��.ي�Z&��rf��Ӱ�N&������Q�O9�i�G)مv�8n���{p�Ͷ�7�&ynx���*���b���'-â	�g�+b@˴���Y,��̌�[A��׶F���A��8걧�ا�)T�g%��]���\-F�'�z��z��=^������B�U�I���������l+T8L���I;&���sU�Z1;���\��N7aq���g��4v�1�]m��p�-r쀾�EF��a2�õV��#���&�$ug�
�Z��<�{n�����x�i��m�7�Nݒ�i[�$�8�c��x.A�5G=�'�DI���Nmܑԯs:{8��)���ێ�X�l��s��x���[$���9����L��؀��su��&�X�MBv�ZҖG[�9����w��{U>D檜���~@(q�p8#����z@W��� �����7M�sr䙳&\�zvQvW<�W!!:Y�:R�j0�q/J��X����FDự�T�=;�c�n�kF��y�z��酂<f3��*��r)b������b@�Mj^_<d�ŗ-�F�;m��΁{]XMZ{1Ɠe�<hd�y��f��ɷ>xc&���ơ��Ŝ�\�σq�rn��S��0�v�t���DL�d)��,�d�)�fi��Pu��ɺ]<��Z�;�rX�{@�]�c�4���W���:t	K��P��'w���7^A �� 93�.���z^�� ~�U��RJ�����0�� 91�I:���껪���s�_�1HA88	�@=~����wJh�)�_��\�O$x�D7&�bf���[\`���陈���_ߦ�m�Bq)0N=�ҚwJh�l�>VנU��E5�J
��=���oj���٬���3�#ͅ�Y�K��g���{�~ﯠ\�H�:k6k� ����6��1��[\`>;UvZ�T��J�F ~��DL��@L�$� �`�b0AP��H�"x�&����x��`��������;�:��U�,mEI�4/߿=�ҚwJh�l�;�2��&�q�X܏@�t�����[X3__w^�}V~Ȕ�(��46�wt��}m��m���f鈙�}��Ҳʸ�JҌu�؝��^Ҋj��{g�.Wb�/1�.N���c�2#+*�]$YV�AV��7��~�������@�\`G5�Cd�H���>Vנwt���Қ����3T6�Wʕ�)*��PU��$���m�Z��*ꋪ��]U�f&z[4/Z��,�6726���U�`����k �M���L�zb"b/��x�7�{Uqv��%j�����bܒu �� y�;F~��2����m�p���o[�%gv=u�"�wF������}��<�Ɲq5~����7u3 ���~�>��=�g� ㉶�x�7#�;�S@��M ��X�m�z&b"�޾�:RJ�U%UWv����͵��f""�����-���R���j!8h�L@{�N�y���U]U:���WJȡ�g<�9$�����M�p���33䓨�A �� I1 �a��[�W�&�vf2f۪PZn�����voFq��5�ڹM�&��Q3�į ���wS0�mt������ ��.Uv]�WujҵV��n�fz"ffj���X��׀n�ft���f.���U\]��IZ��$`��X�m�����m�0�� �p�-�
��Z������w�n�f���艻�{� ��g�"ժ���qui^����y����`��x�DD��0 Aj~���]�.n�]�I���N��إ��Ψz��l�{.N��]([g�X7:�N�f��q�GR���`g.����Нvݎ�3ٹ�E���=�my�[NN�˂v�+s�:�sWe-ʃ \]��;�'ce��fK�Z{y�rk��C�ܶ8�I_3�
j��Q]g��vc|�C��K�X�ط'�:Rv�8�cr��0��n��'v0k'�n�	���s#��H����tv�GF�:�l��'H��ݸu��:�u�9�F�2��x�͵�~���L��m�0�W�d�b�(��[f����4��;�,�$�<�i`��x�a�M�� }�� ��G��!8���)��Қw&`���������r�WeڅwV�V�$`���DD���ܿ�wu��)�_r���i"9�#�Ȇ���Tg������y�Rĥ�tm�^�a^isX78�qH���}m������|��?�����MLQIi�4���Q�����;ɝ����{߷�[f�ޱ��8�m�5����L�7u3Uwr�>���n�y��F������4�l�>Vנwt��S�J��c�����bܒu �� y�d�n�h�@��ݠ�s�j�Ɔv$�h�HI�̕�^��3�ֻLeVs㛫.�=FZ�cܒu �� y�& g3��&��2`�zwJo�-������>Vנ}�e��̑���$6I��og$�����MD�T?*�?}�����?�K�I�s	q8�0@�bܒu �� y�+�qF9�&�$�>Vנwt���Қ��hwcTX�M��n1u�]��R9���'�+�Ѷ�]�����e3&Ը�$N8�iǍcr=�ҚwJh�l�>Vנz���(����nwJo� �W �[^����f$�R��(F��N���ҚwJh�b�rA�R���,������� ���rO���h�� $OQS�f�4��,��Hɂ����;�S@>�f����l�j&P�b��w��z��Ĳ�QC=�\���&�ܼ�d���bl��rH�$>�?�6��ۿ~��k���b*�*�H�qI �[4����)�wjfz���E+-E��Uuv��>��ץ4����@�X��q6ӏ��z�Jh�)��f�虯��� �}V_E*�P�����0�A =�䓨� �wuw|o~;P0p�zvz�;	��UdU���ܹ���x��m��۴α�u��6�M��E
9�؃�3;c���1r���g�ܙf�<��5�c%�1�\�|;iˈ�����q��e�"�c`��nu��m�q�9���m�ˮrm�<�B6lֳ[���F�s�,�Gc���4���Y* H�\��7��S��u��t���9��e���w�mV�}�N����rюZ��3ɻ,+��q'c�m�qo�JdR8��18|{��|�w�|�3��k��sP�.ě	NM�mz�Jh�)��f���F�(��50R=ץ4�L��""f=337g?y`^�� �ὃd� �����;�S@;���mz�Jhu.�'��$����6�L��f"u{޿�~�� ��M ��ꍴ�NA��ӌ�dN#3�"�j��Pn0�H\�U�X�;I�X����Oq�+k�>�)�wt����^�ޱ��8�i�&4�"�>�)���M��Q"�"X� )��A�?��g��ӒN߿~z�o��?��#��c��S&D����� ��պ��������>|��6�S�IZ�ҥeZ0=1��^�}Հ~֙�=���l�'	dPy$qǠ_;V��YM�Jh]�����o���&%��己$d�odI��P�tݻ6������ww_F�>�6��2!H����h�S@��@�v�ܷ`�1�$�q��4
�A�nu7�q�2뫮p߾>PI�s	q8������@�v�&Q^,�# @�#B��9�n���"B�,F@�A�*bq�r!N0� @�b8��U̡�ԅ��IHYB����G�;B��S	�D��+xDȸ̊S0��%h�X��S,A�ID�5�%0r1=0#!Lec1�Z��DX�@)�(P��P���=eLR`@5i<��JBJ�B���%��˄
�d�J�7*�(F��e�%LȊ̴��&���H�' LEMN�����b�>�ȪqP><=�tEt�"��ȩs�6N�M�Қ�̯$mLq76��/��@�YM�Jh~�������ߣ?9M4�Ɛ�Zz�hu3 ������`�����u\��Z�l4�K��ҍ\u[�;+,s�e8����Ńp���]A]��ͷ�k���w�?����DO��.0?%��"#QF' �[4�j�=zS@�Қ�;K��A䉦� ��� {��t�L�W6����o�B������V*)*��L��7�`�� ͬ�c��L�DB5wV�G.Uv(IUU��v�# {��z&U�����g����w���A�666?~�?N>A����7{���������\��3���ez7/87I�.�h']1�L�6�(�2�mV��m�ͻ�wg �`�`�`�{����� � � � ��~�|����߻�ӂ�A�A�A�A�������lll}����7f�fi�nn\�����lll}��^>D��&A �`������|���������|�����߿o �`�`�`�߿p�ٹ3sn\��e�ws��A�A�A�A�������lllw��8 ����A� ���o �`�`�`������>A�������g��7-�&Y��8 �E�A�������lllo�~�>A����}��pA�666?��~�|����;����6\ݒ�۹.l���lllo�~�>A���������>�������N>A����{�ӂ�A�A�A�A�j���������,�6n��K��d/�cX�ٺb�N�./�e�c�⋴�k��7Z'3/����{s�%������jw]]s�u�����`�נ�3�\��۱��롰�c/"��v-I%h�4�i�Y-�e�w�Fl�ƿ������/�ZxӘ:ʸz���B���cs���<u�nw˟F)�:��l�$�t�{G7�<�]n��w{ݾo���z�+���Ц{}dR���2F�3r�^�ר��k���n�f��ԻP�~r`�`�`�`��g����|�������� �`�`�`������>A����������lll{�l�Y�d�ɷwrm�78 ���?N>A��������� � � � ��~��|�����������lll}�~��Mݶ�������� � � � ��y�pA�6667�߿o �b�6?��߳��A�A�A�A�������lll}��~�e�\�n���m���� � ؿ��Q29�������lll������ � � � ��y�pA�666?��~�|���������s34͹�����|�����������lll�{�ӂ�A�A�A�A�������lllo�~�>A����w�����7K����wZ9,v^��]\Z�7� �U���}�eé�g3��[�78 ���?N>A��������� � � � ��~��|����������A�A�A�A��e���M�wI�ff�>A��������Ȏ�DT�(��|�����x �s���|����߻�ӂ�A�A�A�A�~����ۻ�]�w%͜|�"b&����{ܰ�}xzf&b�y�0ָ�llp�W	]�Uui`tLO�bf���x�/�L����oڈ<�dRFD��@��M�Jhz٠U�^�q�^$P�dM/=p��tð��n��uԄ�G>��K��j����#͛#�q�7�C�?[?�6�_7~��A����b*�*�
��IRH����GV�^���L�DLMQ�r��HUwj��wv��:�����`dD�����L��f�޳q�8�iɍ&�z��߮�sk� ߛX����wE��P��(.��р=���1O{��:�����`��o�?Yh���Jժ����>y{J9�	���;]QVka����f{/�7s)#�QF����~�^��^��/�S@����y#a"i��:�]�fj���;Z� 7���r �����%#�=zS@��M �[4
����Y��$��V�D��G�&���� ��,���$�N�X�`)"��P4��������|���>�.�'��RH�r9 �L@Nk�@lyא@=s���dmY�U��-�.wX⍷[Ok�Vq���^s��6�l��7�|�hV�U����9�PA5��1�2�;㉦���jG�z���}Қ޶h{��=�V���NM7����6���MWV��y�0;���D�Q���f�W��ץ4��.vpB䂙#a"ui`��xD�o<���q��k$�?�ъ$U$X������V�xȹ����v7u:�8v�k�/����.�j%J�E:,�N��;�v�Wd��3�"�n���fݩ�͍t�8���:y��y�3�v�a�؍��q�2L;z��B����d������+�z+Z�p[F�:^[n5�ݭΐ��V�ݪ�73��Q��'.��sEQ乤[�;�[՗����m��7Q�Mp��v}q�)r�˳,�'㊦�������d���B.t�3��&�ۛGE�N��x�r���[c�m���.���S�m�����}Қ޶h{��;��9	$I�8�p�/�S@;���uz�JhZ]�O�I#���4�l�*�W�z���}Қ�̯Ȇ�F���$�*�W�z���}Қ޶h���q��NLi5#�=zS@��M �[4
����sTI�(�T\l�&�����v���Kp���n
�n�lt�L��+�"�������u�@��^���M ��r8�F�Cp��ٿf��f6U:��Қ�Jh;8!rB2F�� '5Π5��k� 91��bˤȞE$Ǆ����/�S@>�f�W�����!#�n5�^A yɈ	�s�o ������?��<��㉖M�K�NƱQ���<�t^�Z�XGF�k��v�9����i�G!����@��^���Nϐ^� ��,	�̍)�$��8���@�t��}���⮶��NLk�s1��^A�����.�ʺ�ȉ�����b��k ��;��"�4��������M �����4:&&"+[�09�UЪ�����v��& G1��^A'Y<��'�1y��G�^Jv4y��&�E`�Ҝ��c\��s�N���^�寶���@kyo �<���¹ɑ�)&8�$�=�)�wt��}�� ��4�W��!��"p�9�� ������8E�9�NdNI#�Hh�l���@�t�$��$T @b�J���[��@��3��c��)NI�^l�@kyo �<�� ���r�GH-�.�Ͷ���qn��s=�2Wn��c�b����Hhݪ�-gЍr	O���/t��}���Z�V�C��c���M�@�Қ�[4
�k�=�)��T�D�9�F�M8h�����:����A)�3�rB2F�(���*��@��M�Jh�٠w���5L��RLpJG�6��A M��'P�z��,Y$���@`F1��Km�"B�"F,�bB+�#"�@���B��c�#��ZÂH �XՌ� JB#-�e�4�'�:��H�`��%F,�H�R�$�R��'���$,FÇ#"�D��@`�H�S�,�*0�<��H1M�t �D�#	@�D�-RXИ��R@ьF+�"2H��`"B!����_�, ���)���#!�0bb$%��`R�L(AMBX5 ��@�\C�$�@ ���E�
�j��B$*�jCĄ��&��䐄���	b�B��w���σ����WD��b��i���lXy+v8:(�KHT�R�-��\�zթ��r��i��:v%�wTm��zX熍@�^}�P8�q[s�J�fӷ����E������%>LB�nsu�*uĻ�gq��sӭ��n�B�H�p별�m�DڧcA��
��
`kd]r-m=҈㨛	$:�A�n�S�Ӣv��әW���1�.���[��l�\pD�� fiN9�ˢz������������+�:⼆أ�;{�͍V�!.��]����͝��ݞz�}����*9�lJn3;.���D�.z�B�=v�.��F΄sUkrH��tZKe�AԩA�:�N���MSje�F�a:��O4��\�Jv�����H�]�A8�\���V�8:�&X�X��=���Z���,��Wq��Ԛ�[l=��eq�+=����A�7�{.Pk	�WpD�6ݽ���]�=v��<��In/�[�B��H]h�g�U�rͶ��勨ۤ��Omxq d�ll���du����۳60&��m�A�
8C�Sv�T�L\P�^WJȯ5��+վ���۝����WnKv��J��hYv�ގ�8�U�TN��i��6�hΠv7<<�v�ҷ	��l\�H؛����{{F;Yx���9���]C�cb�o`M�A�z�C�N�[a��'C���$984�[Ml���&�3��3�*q���u�pֳ����E�P�!w����`�Zk���8��|5R\$<\c�L͕@�8�ej�PJ��hPj�m@�[���%WnmN�\; +0z�j���L)��UQ���wn.v�4��-��Gm�4��ڃY�/<�/����^%�-P#����������况��^��9�)��Tq�n�ی�e��V�x�sj��)ё��W��ؗvm�n��*Kv�p��˦#�	���ɖ[Wm�Q�!os�-rQC[�t]��
�����SWL6��.�̘H���� �A�Q^��C��D]=��0è�| 3�����h{�����￺(�q4����RZ�l�N���㲳��������ݻfҝv�!�����t'.��<km�ָ�.1�@8�Ev3!�p��*T�b�ga���7+����m��5YC�[����>~�[���O]���=�on�� ���:zz��s�vH�Zv�4쳇h(����q��`��u�Y��<�W;sI6p+ѩ�����$�7-���|��M��2jTX���<���v�%�4�[ �Wں��;<�vn^WI�3Z��2��������f�W�z��>���&�U���I# ͬ��MQս׀sk��gDLDEٽ��HZB�V���X��׀=��=3\�� ;{��բ�q�̉�&4����S@{�� �m`z&+�{� �}v�J-]ݪ.��F �S0LL�or�V���Jh��Y#�# �1
d�q:ܮ��7]��9u�+]u����]���V���.�Ls#�F�p��f�W�z��/�S@���,� �B5i94�~�s�0|��O�� g�;���� ?�X�4̥
�$�Ĕ�@�Қ�Jh��@/��~qIڴ�V��WIUZ0=1����>�� <���k {���ǈI�s#rI�C@/��}�h�S@��M ��m$Ȝc#mHEQq�ٽj�Fv�%�`��9�cv�6��y Lr�#M�4���/t��~�Θ����or�7�����B����mI4�)�_t��_[4���9r*w�HF�q�h�)���y;�F��B)���� �D<���y$��ӒH}��*VZ�t�Uh����LDEߟ��ϼ����?�3 ���T8H�V�EU���k ��DDsy��;Z�@/���λ"m��
!"L���+u\582�C,��]���ls<���{���?�橑<�I�$������/�S@/��}�h��B717�+F ����LD�or��� {��֗`���F�9��}m�~ְ����U6�k\`��w	�!*����X����� m�0��9&���  u��y����N��6�ʴ���]]�K ����3=�8��w, kX�j������NY�r�{0YJ�в��s-v��8��y�D�i9�����p�/�S@>�� ��4�Jh{��r(�24�Uh��Z�DUk�=k����陉�61Tt$R�+�Jʴ��|��S0�Sָ����>��e�\ȞE$���{�4�Jh׬��Y�_\WdR���Ԃp�;�L�=_s���|��S0)��y��>�I�nۻm2l�,�m��ѪK�Kc���F��vs��!�pvӭ��gt�d�v�b�]n��������h4�D؍����vW�ذ�	�__�}v����rp�ng�Ľ��C�H�<�1d�&��a�mG3��B�����L�6�V{s;ѷt]��/�.�{X��]8�3�<F�<%D�e�.ɸ�Q��m�q2Cl7nܷsl�=UuA7�s93`4�˳�mї\:�{N���ǭ���@��ɍ�j�aɮ�ժ��°61?,�O���=�א@=y�eN�`+�J�%��������\`l�h׬�=Z+w����Ci�^A �����=�����Q5Л����M �����X�11鉋�߼`?G��
���5Hn��4��h��;�)�|�Y?�<y	�L���kID��Y��:b�d�0�<:Kc�z%Y��ݧNI��\���NO�=���{�4�Jh׬�=㿫�S"y�B�h�՘���F=�y��o��{���4��h���nbnA�h^A z9���@=y�"ª�%J�$��i5]�� }ϖ �Қ{�4�fW��
F�i�" �s�8�<s>�16Ngo�>�#=����½
^�N��g��e��u=��;���c��\!���H�F����� �=��� '	�rĢj!�7�Қ}�h׬�/�S@3�*W"���E�$�����y߻���@W���U�WW�\�o ��t²Va��
�h*���W��`Z� ߵ3 ?>�@��^�dS"�c�RM�Қא@�b �s�
��a�k�ZZN��=�n�v4NgBvn%X�t�#��Ȥ��)����p�;�)�^�@>�f���M$�H��H܎C@>�f�}z��Қ{�4�fW�$�8�rM ���{�4�Jh׬�=Z+w�wt���I`z&��� z���X�D�a�����}����.En�������4z�h�`W���jf�3/�����Þ�`-�û<�x�]�+�I��:ykb��6�쮓Y�WAtN�$A��Ͷ�?g؀�l�@=y�� 6�0���'��$�7&���^���M޲�/Z�w%�f)�L�I�F�z�&`|�0�U:���6���n)�ID)��p�=�)�r��@>��ץ4u%�'�E�F�rsd�y�u��� ��r��� B��Y���t�7w&H�ɲ��+����dS�r�v�N2��j�?���#�ޜ�;#��ll{W��t��L�Y.y�il��	�F3���H�ۜݷ��ڝ<��q�q����j�dumԓ"�zZ�t���@u%�a�s��;\����W;2#�#ێ̦.#Cme�zۣm�����[��n�ɼ<�;z&�42��h�S�	�"�m�'����w�r�ɾs��˛7f0�au�f�E�I�8����%'^#s�i9�5���2,�SU��� ���x����S0����En�#�M��r=ץ4^��9zנr��bE\���HA&���4�g�@��^��ֽף0�T�U(HWJ�Uգ�&&f)��^ �{� ��fLDL�o<� �p�BE\!\+J�+�6�n�F��>�Y��9zנL�-x�rɸ��(ٍ�7-ru+��^��ӻ`Nz/\�X{m\��P�ȦE$�#N?��f@>�N4.� ���������O#����O}��s�1Ts'o��rI�����)��#�I�$�IrI��h�ﺀ�l�@ly�� ��"#�r4�IǠyzנz����YM��z�En�#�M�19$���S/�8�����������S0U����Mv�[�w��7	[/�pu�[=x���[�t�F�ِ@>l�@o6N�6<� �*�r
d�q���4^��^���)�{�SbGe�?d�y��J��[�x�S0y����A$�$; ��� �VH�O�`H@�@�U�!Q� �H! ��į�Td@}$��H��
�8�
J�����:�0�B#0uMZA����ԉ,��"Ā��R4&��HQ�eVD�Rx�Bb����hH1���1	H!
�� Z��`�#���k�L��`�OX�8�#0�*�3 �.�����B�#�Z�A�F_�G� �Ĥ�	D�!m����� 	��D���"��"��#�#J�zF ��G�u >(���}���z��^)�2)&9q������� ����|�:��l�@7<J�
H��ZE�0�i��!��_�r�ߞ��Қz��#��t���l�q�1#r�}4��.��[z�z�qK��Lr���h�k�<�k�>z��������V�B��J���;�@�bc� ���d����"=11v?\u�UūVU�Ҋ��I`�?Ɓ��M��z��4_"�0�#lp��h��9zנ^�d�C��H@��(@��
R�EX������rI�>��"�]�WWUv��u�z&f+�|�����jf��΄*�PR�QhG-�K�����Q�t���x�Jpj�e�(�+e3c��H'��8�_ {��4��h��=Ϫ�=�,��2FD��V��Zfzb&&�z��}X���»#��NA�h�)�{�U�[f��YM��$�9	i+�I# �o]`���?kL���DǢ&b"�����{!Z+��J��Wy��& <�A �� 5�� 2���X���\�m��˷L�r4[F�������Bf��w�y�l;�:yH��:,�$�^��A��lwBn��]U����7��_}';c�d'n��[����N�r&����][�^Oe�W۶�ֲu&��`��=w��;$�-u���!�GB �)�v]�C%�k����N�0u��Xڎ� ^ΰ�Pr�.��6j2ZpA�l�y��lqyߞ���}�鿏���C�V�s6�Z�'�z���*%v���ѱ`{T��It��3�jbm�'�=z���4s��l�;�En`�F�&��4��������5�����`��`|��B&܂xۆ��}V�}m���^|��5���lhBp�WV��U�@rb�d�A���]�̟q��d_�d��Ɏ!94��h��=Ϫ��٠}�jd�F�""ҡ[��Sy��^�6�Ζ�s2���5��k�[���`�rH�����#����M��� ����e4��`��9䍓wg$���v�"| > ��"�`>ϖ�ˌ���~א�*�V��m��@>�f��YM�Қ��Z�9؞7#i��&ےhu��=�)�{�U�u�@�u���,�(��F��f�3�{�����z���W��Œ?�B2��GI�v^ێ���e���fz���Wiy�y�<<�2H�NA67��z�[4^��=�)�{��%��(�$� yɈ� ���͓�뻪���H��UiE�*��7�� �w{94:H�0U��	c311��� ߵ�u��դpi�r�@��M��z��h�)�}Ի��H��7��9z׀z"ff=����?r�n�f�������Vt�n4�籵և�.��y9��]!p�����7.��Y�+t�EAH�ӏ@>��ץ4��9zנuy���M�16ܓ@��M��0��� ��Y�3Gu�:�Aqi���n�~4^���٠z���g�T�B'��lm�@��:�=$�ǐ@��n�����������_��z���rA�8I���k ��DDG�bf_������� ����?��~�BJ@���b1Lk!�u�)�w�iw2�gl�v�m�d�A�k��iE�*���\`���m|������X|WbV�$���ZB�`���m|�����>z������>|v"��%j��Wj�F �{� ?6����K�Y��-��w��7"q9#n5V� ?6����wS0:bb&i���_�+���m����rMץ4DDĶ��:���͵�G�1��՟����.�kNǴ�s��9�tI��˷ms�qVSo/0>q�m�V��óf�X�q�s�;f�!����&:v��P��[<��g���.nr��~0n��l��s�����r'Z��6���O2��&�ϕ�����λ$6�㈻f�tv66�m�A��u�t�N�.��ܛNë��ڮ���v�͕���A��HtQ���<dZg�.̹�d�fb����.[�n�Y�R����%�n���EB"�Nr���+���lȬ�#����m�`<M�@����6�n��mDL�G���ގ�肎!� �6�r��@>��ף0�L�蘙��5��Бqj�����^ }�� ��f����� u�׀w�t&8Ȝ���@��M��4^���٠wQK"��D�Ē� ����3��� }�� ��M ꫣȇ#�q x�0��9z���Y�縀u�Б�ɸ�A�:r�4ڬԫ�I]�I��� ~m�穞�����~4���r'�r4�iǠO;��)�bʭXa뻪�wW�lYא@>l�@9�屬nF�mLM�$�=zS@��M?�3N�����Xw�;�H��,��h�)�r��@>��ץ4=r�r�6��xۆ��ֽ ��4^��;�S@�^�,l2di#����� A���J�.�]!��䠋�T�<�p�۩����{����u�Vy�i���m����� 6<���@>l�@=|0���Brh�)�wt���ֽ ��4�)dR86�I�wv�rI����H>�dIH��P$B2@$B#$���?". �*�}?��������hu%�'1�rF�/Z��m`=L��LL�So8��ȻQ8��Ӎ��}m��Jh�)�r��@���p�#,J(��E�R��V�q�:;�/V�y�>g�8��������N'���m����߬�h�)�r��@>���ȭ�$���x�F���陘����^ }�� ��f g�T�F��i���n/Z��ma�15[�q�6���	�EŪWJ�Uj�:f&}311w��� ������
f"f=7�9��2�� �]�c��I�!I4^��;�S@��^�}m�Ǫ��H�ě�"d�}k:��g2�[`�3!dy��:�e�)��BG�I!4��9zנ�k�"bc����/���UV�ժ�V�U�`_7y鉪��`�q�wt���ċ���r'�7�iǠwr�>z��n�f�����V��i+���wv����M>y� �\`O]�zbfb���X;tuڅIZQUWv�wS0�10��_��h�Ͻߧ$��(*+��(*+�Ȋ
���
��PTW��AQ_�E�EE�D��A"B��EA" � *@ �AA@� ��EE�Es�QAQ_Ƞ��"���(����
����
���(*+�"����
��������d�Mg���H�f�A@��̟\�ʾ            �       X  ��H	T J�*�%B��A@*�T�JU��*�� *� ��
�*BP�0   `H    �@ _|���4�5�^���|��M+� =�}������zw�z^�>��� (�/N[�^�}��� �y��w���U� �����3�׶����y���� 6� ����������:��=   �P  
  5Gu�9|���S���ɮ[� �T����k��Z�����[��p ���ŝ� Y�-ug;w���    l� &� 0  �G;  �  �   j��
 ( b( �� "  �  $P �  ���@�� @ D ]`  l �޻���ˎ�G����W�\���m^�\ w5n-Ү;��/�nl:� }P 
    1 
{�k.9粮-����o��«� =}*f���^N�yy�=��ov�� �{mn;�=��/ �_}�������k� {�[n�:� <�    ��[{���-�NN�zy=]��3R�  �(   �P�<��n;9[�癫�S��o��o�������rk֜������{���m�}������ 6�[ռ�ǹ]�� 4��}���}i���{wo}{ޕ\�v�� n��.��m���y{�7�ڼ 4�Om)R��  EO�FS5JT���COǪ�EOҟ�4� D�*�&�) S�BS=J��   ��&Ҕ��2�⚔&�#�}�U�J?�]�g��[�I7N��J"�����**+��(*�**+�PTTW��QQX����������!�!I1Ms�Lrk���������D��	 ��8.ҐQpF����P�ܼ$��7ǒ�m�&����B����x�\�r�6@����Oǋ�_P�E�RH��`�5����`��y�����S���T�U�V+sr��"`D�)a���C3�zŮ�6b�<�Bh^A�@�a7$�Ò̜��L)�J�I��;�^I6��!8JC#Y6q���#�*8i���JF���B�S6/"XH�!���r�^c<9	rD jCdr�J�Za�)D��a\Ůx{Nk�0�!S��U��bȐ+��E����tR|�H��H�8�XEb���B(C�,xC�x�.���3���q4"�=�F��� ��+���'�k����W6�@�� &�T�Z�J�@��J, �h�(�F)�
c��"�JT%���!RW������4瑐�����y<��Y!Xq�^i)�aB\��&Q�I*JWy��,:*������b�XR4�'<�����3:x�,1��
F]�I!^jk ��*B�w�p��3�W�(HH�`a,��BNp��!p�BT�$H�0��Q�hP�璓B���
��ٙm!@�*
�H�$ �B)Bk-6�u"@�9��Äd���4!q�+�r��8����8x1��$���勄 P����!L7�ak�S�)-8�HI+�2Ȑ��jQ	l����p�VX)4���#L"�!��P�1"�\0M�0�\\!HXW,��i�;��L2�`[Z#,BWH�0!V=4�F����EH�����(nM�=���y����B����!��C4�@l�)� �#$�$�Kb�@沚���n�(B���!��Sy<��0�Ð��Lfg�sHms(�%7�%3o!�h������XȒ���J
t]5bK����CO�5ĉ X   ҹ!K��$Ha��$�cYJ��8�y/	��(R�xs�.p��d+��n4�Y�a�0�!	q!B0��˧x�ì�N�'Cۜ$x��]�K����X��� B!fJ��HB0Np���\d%�K��CC�="P��L�� ��4�����*1)�k��(�Ð���� ��З����=��d	�TɄ�q%%�yc$$f�� D���'�3YF�q%	H���B�bhh���J���'$xnÅ%�, os0�|�XV�e�@�Va�����7-柏|8Nf8lNR�,b�"� ����)$B�%),Z�����Pa1�xJ���hA�w��� ��.meX�p�1��I �e�VV�)BV��ad
BЈҘ�G)HZ�C*H����p,+`E�5�ĥ$d!Z4���kF~i��H��_d��K�8y��(ċ@�8B�aR-��)�X�!Z���	i�=&�2]4�27p"´���\NOE! �@�J���i�hi������	�$xo�sN2JU�aZ,�nV��i������p9����O9�9��z�������<c\J'�p�i����4�*�����a�`^��J�(@��(
���j�/��
�@5 41�0ᰨ@�뿒\4�B����]9T��JbL!�YD�^>p��{�	x��y�.$9������B$I����as8'���B��(���5�<�8_�	G4��4�_A�E��Ӊ���T��8K���&s<�q��\�+)� D� a*�F�xl(H��?'���o����o<��a�$��B3sg7�\��y�!3ß�'���qz�5�R�~H&��DjB�fhK���%8a���?p��z�P�`�E��U�VH!G�杆��9�-�2�~��!y���H�f���No�~e���e�i�~�Q�L9И���>8��"@�����9��yľĆ%�� �@�e�˜u���a���!<��$�e�\�/�>����`B�c"�ᔸ�H\u����9��p:#���FP�.�����	�P��ӓ�s����w��Lta��yq!H�٬��l��#sy�6 yw�n,hƇ8�0i��I
���0�����ty�q)����$x�0���D�|=#�������J���:�������T04�8xs�H\���0-��s�YC���K���Ș�bH�$�A	xBJɜIe��w4�%e��y7<�����F-H��B"�,�c��c��F�Jd�
��H�}I�hB�4%�s�%�$
a)���_��nHi��j���˄(��t���B,B4�)DĀP�%���U0�0`��	|�I"�S���a|�!caL!L!M9��G"L��M���`R�%8p��
�s�_С���K��d�\ӄ���B�@���,�@i�����~��Yᡔ�s�ҟ�_�� Q������ۋ�B�WC��ٙ�Π@uqX���sv�.s2�s����!�K�!~`�t|�w��-\"�"�X�<�}��~�B�.ax��О�S d`�i��,�(AbbR+��&�I��:�$
���R��(`@�0�����,Z��e$��S ##\��SXS#]H�	L4b���L`�Lܗ)���&�q�ZJ~=�0�.!�>����5R�No=��$�`X��#���o��@�������p�8sf�!��1��� ��
�C�X	��pg{�\qe0�!��P�csr��9�8y<0�0�ǆ��1�#!pW��0H�@�������{)!`G$��$$?^$��SR Q�bP0��=<8x���3"K��HH%=a@"��0�%���J���f�Ȳ�!a\�x�.��&�V�h����35��!���f��S�	C����HSX%i�Lº��p�S6C�_9!�)�9�ְ(R��3u�֌iK�ņ�Fp�^r7��0�q�LaL�����j(i&�7�J`��y�G�5�`Lq�C܆L�d�u#S�h'-)SJ��A+!�n�9��z���y�+���g:��~����=�Lm��_��ZuCt�,���e6��3��
"�Y~.�����aH�X����م�y�J�����}^�7k�Vz�j�R·+��i{4��]W�)Ї��f]5�:����[v��?mU�cX�ݺT��u��j���{���7���7�~�!	��~�B]�t�$O� xS���ZG"�������@�43r�)�<B4�6Nx1@
���5p��y��y��F��!����2�y	� ���c��G��j`hpH�y8�xHH��x�.�<��I����"�a�r�9��˼���f��a�.�_�s��r8�T�� ����x �"A)�F,)&'�!8k���F�º��FɁ�%6XH`Wa!p�% �"��׍F4������y���n>�g�#"��Jl�&�9��*8������h�FJ㩁 �(``i�`B�.�F�`l�j�@(
�c!!&K��
s�o��pb�G�%��HsY ��iMD�2��_H�Ld�x�J���a�Mh��!���)�����^$��4����Jf��SSȍ1t��Y�n��O�),�;ߎ���3�}g�ӯ�_�         m� �8 �`  $ m �����"m�H���Z���N둩Y���
�)YJ��  ɵ��="�v0T�u]R���)����   )����P$O@c�l��ȵ�n����B��UUI��g�b�Vރ��)��m��L���RܭU*�e����U�^2Uꫪ�k� ݈sm� $m:l��ΰλ�g:v�`mUU@eI	�>�Ux��yYV���, M��]��js���p8 m������   ��-�� g�KHu��e���l����I�^bu��ۣ���θmz����<�ô�����-��#Wqc�����]p�\r��2���[H<��^!d�D����3��@��l����`97]���m%�-�0�am$Q�ѷ�ne�q5uUv1c
�V�<��UUN���)@^�q+sf��jٴ���Y���s�ݺۅ�]�OM� �5S���HI۶�)6`����� �d%V����֜�l�$m� �»v6�n�"G����:3��ݗ�Ҷ� a�ZYe��n������M��@ �m!mH��[p蒀� 8-��K���P	  �   Hp什��	a�6ۀ�`�(�` p �[��v۩v���n�G �mmne��R�ڵ�`   ���l 	   	� 	��  #�7��<�gQmI ��[t�L�i� � H  m�8�+�  ���Ӝ.�m 6�]��������#m� p[@8H�g ����i��k��*�Yc�P�
kUUP� �6ٶ���Z��V���rgg/������l+�[05�Q�,��+S]O]�BsUP!̖FV�B�Z�ZuM���@W����lWp�cF��+u:It�6�tI���ܶ�c��%���t�@�Km2I������UW��*��奶�m  � 9����+�I�p�`$�,2e�[M�`� 8Z���l/Z��m�  ��v����mZ-� [d$�p    6���ؽm� .ى�W��Z�ؔ
�]���p�F;UP Lœ��BO�3p�-;�kl-ʵ�nQ��vN7�U�+�����]MUVX���y������ƺ�rڃ v� �P[M�\��D���Q�H�]*����UR�t�D�KN��[C��A�4[Sk�	�ue�:�e�w 4�����m���-�  :)��n�/Zu�զƪ�R�@[M���� �ېv��j���B�*��]���-�U)�EZ��@�<��*:�j�{oo-�����f�ƀ �mJҫ��2�:����[�U]ٷM�����m�
� /]1�I�Ή $�/M��_�
��fWI�+r�,��
�J��u��� �|�4�� ^�-�m�%��jC��:m�,1�פ�M�km4�K+�m�k�j� �[s�BJP[@ n�r��4�$,j�m� �,��l r��*�{<�l�O+\��` �a�P   .鵶Mz�Ŵ�     	-�p���m���gR�Ī���UR��U�m  �Z-�]�s6��-�5� -��A��=�@IeZ��^��6��m-�z�l�n˯Y9of�F�҅,<�������۵,���;vUhvQX�����N�����e�χ�!f��N���@oƙ���t�*��
�ꪡ�V짥�[j�m��� Ā�d��km��$ �Y� $ ���m���V�  m� �:�;\�`s�RE��y[�j��Q���n�ą�@B��h88�F�'Ki�m�-����H�m�ַmHm��$�P[v���֤��؀H�a'��Hӡ -�n�p &�Y�]�D�@������m����V�]ٕ]���
�^k\ۭ���IY�`��m7@UU@]T�*ʠmp9�r����M�	�! R��!7Us�-P��ܬ���  ��amm� -��n�vv[!4延-�Z(F�  �[Kkm�K@;Nif��[�-����vͤ���muT��6�Pq��e�ݕ٪��
�����շm��z�@�r� /[a��E�[�lr��TJ�Ri��]�2��Dm"J"Kh��PR�U++�Gf�d���Y[��Ӻ�VX��geӵ��P�6�`jB��l˖�� �ꪀ�U�q�����R  Ε��D�g:� ݻn8�j�vͶ[D�	�=<��� [N6�^^����� �`I8ᴙ�ai�&Y5���  �j���` �����a�8G6��3�m�	�m�9�e�A��(�n%�ڪ�j���m�m����H$-� �i�-��Z�� �h�D 5] �UU@AN0� m�g�ڴ逶��F۸mm�N��>����j(�V�ą �mm��gK�lJ,%�kc#+uXňV���m�C��P�m>�m����m�[�ض.q�ɵm���rWnM������@�8���g]�����ڴ���m�yٶ��[US�J����a��! �m��9h��
\;@UUVҭU ���m��lNXt�tq�T���˵Ul���Y�Il�_{�XbA����+�v[��+m�v�@q�ڠ �G1�Vİ@ [=��O[UP��/GK�s�V��Mu.�_��Oya�@��ҢL�k5  m�-���-����=:��V�u�\��ޅ� ��ȷ�Ԥ�vK-Um���l�{u�V�+�UUp�U*��SXv�lb�j�Z����o�|���tn�(l�f�& �����6ݘ�9�$kJ���fm�C�����H���rMm����K24�4�p�� �+����z7��Ӫe�`&�I��8�I�V�M�6u���U0nE��2�k8�mM�v#m��8r=kvv�yL܂pn�AvX�L��$�($	-�nH�`�l�G���� �KR�qJ�UUA�u뀏�����),�@T��2�v��$m�Í���sv�`Lي�m�ζ��i�M! ��hm�m�� �|�m8  4}%m��m�d[[2�0  �m�	9�9zL���@:tUT�W�j����m�� $��������e��Q,`�p8`�e9{)UGԫ-e-�` m���X6�  ��knn�ie� m� "F�6ܛ���X�����$rB��U+�T�m#�@�[@6���í��h     88t��۴� $���Hz�+m�p��$��SkA����R�H�հ���m�l m�l���d��n l�	 8m��skV���]K� �� ��m�kj�:kM�[@m����j�pmN.۰ [��slS�Bi�������m����D� m�%�Ү�&�[ U*�,�^-����;K�$��mJ�R�mv�*j�傕v�ָ@���v@���D���   �f�l �l����cl�6�   � -�6�L� :@[Am  �  ںlM�pm� �m�Y�� ��    �hm���h  h� 	 �H �8,�]� �vh���j�  �G̟-\���eZ66*�3��T��>d�V�F*cm[ Y-5�y-�`i���������	3�>-�m��� :��m�p��6��u��� ����Zl6���� �h ��um��2
���lQZW2.�;da��X�l�[G p � p��� -�v��T]�mVj�N0��/����kI&׭�n ��� H8  �   ��2.˳m��i�M���e� I%�.���Si�8���A�V�������W ��Ͷc�-���Z��hZ�g]	���z�Sr�Rٴʽ�UͶp �`Zi�-���5Iv��h8۷A�EU�8|Ү�U]R���*�mTު�R�xV��*����Uq�  qm�(mT�UU/.Ӥ hWq�N���c���e�2A�]�t��ήks�m`�j��V�ʩ�w��F�Of�VV��n*��	xt��q+*�mZ�3]��pX�
�U������4�v�H  Imm6p�f�d��!�UDJշK奸;atێC[m�`�,�� 	���j�&  I���P�9�ڤ�.m� -���X��v�tW]V�,�4�[���T͡j�������Jm�[\�e��Զ@2b�vm���@�ky��z����[xt�� � mz+]��ڶ{�����m��m�Б �ֱ��}���w�w|���UY ����v*��8�`�q_��K~��>����u�T|@=�9� ��j�}P|S�1F��C�*����Q{�U������@\E
,���W�hPSA�����@~}G�x*�(� G�OC�@z�t��?�@�E�A鿕PCN���(`���b����� z!�H�N���Tx�D���MD��@�a��U�*8��P
��E�f ����P? �8�Ah����z>�8
�5&$��H@�"�F�"DI��	0�A��B�1bD�!2C�`��<^�= 1 ?t�U4j	�(?���O à=S��Z � z�W c@���D'��� S��翇�{�/��U�C���'�E�S��A�ꯂ�tW����z(�
�z�.���A�D?��U�u3���?T�,i
D|Q� +� �:Ǡ ~ pA4Q}C�V��EQ�z�P�
<uQ>8 �QN=Qx
�W�j��������`�P�
�P�}���.ض���$�m^�E�\�JXamM��@t�s�zM������0�v�iݭʢ�g�t��{-��]T��eg��(]66㇞�v�t;��Ͷ�.�k�/#U����Θ�=�L/�@���ܖ��*-��[w:I� �I��[9T���fڶcK zW�k��k��V�/F�;@�X��S�[�f9Z)�����h��Wx�9��;i���g�<�l��U\�۰�C�.ʜ�Ԕ �Ua��.w<[��J�P�.eݞ�[p��%�o+��b �\�ǫHQW��)
l��FzK���-�0��M�a띍��n���:�:�C�:	`%�Gj��6S�SS�c<�WX*���=s�*�XE�۝�ƷL�r�r��l�pb�N��&<츧�\��V�՛N��$YwFj��5�@�[&Y�s]l�9��lu�����!��<'hz^���
�-m�\cN.RݷZ�w��Ɇ���ʍ�ZA�e7>z,ϯGqٞ6�"�N6�^y[��mru=n��i����3���`g��o��,չuJ�eu��sY�9�z�˼Rnv�nΫWQqW�*a.˩�{gշ;���J�Uy�:�f�3�;���6�n���Y�/�m�%K��:2�Y)Ka����lRq�le�%�z�byҫ��<�kǘ�r�N��M+�SNɉ���K��*���zd(���9�:rt���Mx�nn�h��fM�1�Вi،�7�/*�Xd��y%[k���<��v��1=���3�Z���hSeSV���l[D����:���\�"JpdS��nZj�.k�\,ꔚܫH\	)��)ݻ[*�B��6�>��.�8�.�T��/;Sj7c;v8;n�:U抄u�vm\� �Y*��^��7R���;m�i��\��X,{�i�B�#U�FtU�i�M���g�Z_<��T{T�i��8���ps�*�.���6M̙�f�d�i ���*�@�$$I �#!*0a ���<*:z+�1D�N�x(`��qO�
Q�1���}��r������l]���ƨ���,r�ܑn�SȜ:*9vm��5�mDvǛ��L!����6�Dv�1�ɮ^]�k��lX�r=�7;]��ms��ָ
��ۯn�a�\�Eu��s����u�g� wͰ�K\0�sv�ڝ.-��7I7���4�j,���6Ռ�Yŷfۮ���q�c11xD7WX^-�{�:���l�9�̙�\�ə��J{dȞ�<��v ��o�m6�1��j���qvנ}�`z{k��!~�;_^�EqԮ�swEUYUu�~��3�BI/D%C�}X��M�{^���X���ěqf!�׽1�n�L\�lP`mލ:�MbRcP�)�s��@�^נ}�)��g�]o��v���Eq�k`z�L`{b��zc ������B~�ݹ`�ćBS�3��5�mul��m��v�ͳ(	i䭳��a����P`u�L`�&�uzoE�E0X��I�4�v��_ꑐ!jP"�Y*(����^��s$�������P`WJHJ̤��2Ջ0��:cv(0:��h]��FEb�8��>W��;�_	}>��"`{h�L���V���Ōؠ���쾘�7dL]�z���$�i��8�NH7k�Fku;;mn��l��WG5��vӭv��<⑉���U���@�^נs�S@�u��%&5���9b`z�L`wtt��ޘ��$F��QF܄q���8��@�{w4�ٓ�`DY�X*H A���$P|Q?(��<�ۜ�p��h\W��E##�'����׽1�zH�����S�$�D���us���٠|�k�7u��9DB�����T���権�"-%v���=w1-ۇ����rl���N4�:>�3��HH��<M���������@�{w4�v���EPQ�#d�)Wx�z�:���_��}X�� ��**H�qH�r)����h\�zD���@ⶽ��Ǐn7UU7v��k� �ۼ��u�DD(��|R �jW_qW������o��v��˝�l2�VZ�K����1�����t�GH�黱�zؔJ2O��k�,[;ru��t�������>���֖��[�D�!m9>���@�,��������3>@w���*��5�<�)�8�ؠ��ޘ�7dL\�݄��Q�0X��I�4
�k�r٠|�k�9�)��nI�<M������:cv(0:��0:�Y�(�68�M�{^��߿w�� �_V ~�w�j���I)(@����w�m���ɺ��v#N1�g��[I[�۞�m�.��уM&��%��6�co] Gߊ�� z��v1]��+��uy���Dy��#uq�cu��L�M(�a�ꉊ[�Q����H|�r%ܻ�]6�3rk��
9{;q�^]��%���˚��v�[\�v)�O:K���6��q���-�v�c=;�6 �L[�HA=u�w�e7K$�]}T(�ۼ�7.r�-�N"ipQu�wƮ:zԓd�*p]�)b��ָ��k���N�43��~�|0:��0l���1��2��r6�Q�h\�{��{�M���@�,���z4�K�S�QH�vD��Θ�݊��H�3.	Er�ӓ@�^נs�S@��k�r٠uq\j��5##�'���D�7dL���~�����t4/<]���K���[��*�'ֈ�̻��T���%�tr�*K��bjO o}�`�&����P`WCwi��\˦���~���1P���0	�����G�D6ϯ�נs��4�[4��X�G�86)�$��ޘ�݊�"`�&΋���$���N=fb�����L�D��ޘ���GE�VV,J�����`�7x(��O������ �{w4
�i���'�ƣQ�!9�u�b�p��i��3�k΍�\s�ڕ����FC�.�*�BBĘ�����1�������@����j6���&���u��Dɻ�� �_V {�� ~֩\��F��$R=�����i���O�S�sy��}~���$��Օ�`���5!�Z�V�s�����r�h�ےE�H�6�#��7dL	{��A�/zcw���eD���]��Y�S��5��un.p���e�Y�6�k�w7��O��q32��L`n���vD�'�R(GIȜz9e7��3�bG��� ��ϵ�rQ'��:�T�ܑ��n�o��s���v�����ӭ,M(�7(����ٙ�3��xO>��v�
I-�
�"U"�B!_��h&;��n���1��l�9�iɠU{^��YM�ڴ��h��2&�s$�ɛ���/:Xl���[�����P^:zܚ�yY�W>v�dsAM�'���~��-}�@9�f�U�z�ueq@X����4_j�g썇{�M�ޯ@�{w4���"ɏx6�jE�[\�ؠ��:[���eZ�Q��Grh^נs�S@����?~K��h訩$���n=�v����O�����u����N�O���m�Snٓ%�3M�]d�&˺�.�N�Am�Z;�vQr� s�����I">cF�v��O+�=o�W�F��zq��G3��un�r۷W[�q�ZGr����1�ͦ��9�<Y;:K �f��B���%�:��X�`��r�D��#��9�ܘ�c`n��i���76+����l��L�Fm�a'O���d��lɄ�ͬݒ�Y�(<QZ���{���L��3ez*m:�v�,'C�E��c�������b�c�Ӣ�]�G�����n����r٠U{^��YM��tk�s�Z�[4/]`��`ֹʈIL��2��&i]M]�WU5w�9m���(�Q*��= ��ur�yLy#QL�H��wGL���D��Θ�:Y\PI�RW;^�s���{^��YM��L#x�1D�<b�U�s+]�:��c3Ӳ4BE�58\� ���ݙ�'�d�dǎ<QǠ�@�N��݊����dYV��%��n���$�^��� ~���Aٹ݃��c ݑ0ip�+A�RYw�f,`n��1��_����������ǒ) �Q�hܶh쉁��1��s���]]ͫ�WeU� {��В[Z����Ɓ��נ{�~�>��d��I�̌���*qI4λ���sM9m�ٲmF�u�5�9�O ܂����y�-���ϵ�D(Y {���|��qj���-U$,V�݊��vD��Ζ�;N��)���85!�us��9{���5 ĄF!�a'�`�� I61`�
H��(X%X��!	E�!!�� 16����y}��3�0��
���A#0�,0�8.�D�jB+me"^%�v��D��8D�*U@B,x~`A��	�iU��j���
c3��
���Jh���E����c��������Ip��~�������''Fs�����`�V��� � a1hX���HAH4�XU �2%F$IF`��HP�@� �� s���O�:~8>�b�:?�(A0U�
t z����4W�B[�7?�������B���]��ǎ<S"�h}���{�M�w�߳��|a�H�J�ݾ��]'])�Swt�nz2����ӝ2LB����u�`���B�ݷ�5VLUU�EQjEoW//<vsF^w)א�����bQ�c�t�N�忽ﾲ��(L���n>o��4�v� ����|�A��}X����M*�˻&��b�D�7dL�ﯧ����|?����wk~߲?ܝ�E�ui�����^�F־��n��D$�\���=�Q�@I��R{��߲)6|�����}��9$�D�{߳�4 �� <�ʧ��"&��������	l���k��+WVZ������Ku���I'O��D~�=�ׁ�BQ>����6n���9�xP"'E�-��ؽ�D�O7(�F1b��g2�@��c��l��p�)�g�V�"!O��� ���9BS>�ۚn{�$Y1����kf��=�|��A�;�������,�YV���V�Ę�A�;��J�U���zyl��**H�o$����;����l����(����A6ܓ4+���٠w�ـ=׋ %�!(I�䪪d�؎�����t2�0��0���3�7E!փq��]�n+�c�0<�;�v佁5<��x�|=�w�Ph�q��ft�gVٮ|-�S��%�
��sDM�m\�rh��H���ػi�nuSJM�m�#ū����m��:����gGFF�g,lu�6��7���%�n�i��=$g��!-�R^��']WT��d�U����y�2�m�srK�i��������ڢd�oUEʍ͋�t�����n����0�c�"�G�_zh�h����g��ى>��@-G�������΅'7|`�b����x�Ao����I��K�Θiwn��v��|�d�� v�_$�~�;{��(Jy�� ;�+���*f��n�j�gB�S!��x��|�B�!���$���, ���$�&<q�L��@/-��d�:`dL���ZF$x��^���;ny��c��6�j�
���9|���D���񨤎M����n�^[?ϐ�4���#���&�Sg$����� )�!,Q�
!M<����x��3�B_�%Ts����<p��&ےf�W/��^[xt%���_�� �ɳL�AV�`���6D��	�05^נ�(ՂA�#�@�,� �^,��� ?7xDB�.zKi��nu��*N�4nk�kk��I��f|Y��e��(�v��8s�U'�o�`������7�ـtD�g�S�I"�&�|W���^[4ؠ���� �)%t�+V^
ŗX ����l��P����J=�(��DDb����� �x�Ѳ;�7F%���%�0'r�wGL�����BYBJ�Yw�1	��`�{{��ou�vـnѵ.eDV^�jF�f�і62�{a��6�����v�莎�E�#Dtf�� �m�zO�J�X�$���}�IT�SԒW��g�$�cΧF�$q<$r-I$�-�|�U>��$��o���%�n�RI.�j�4A�#��K�ڞ�����>�$���jI%yl���w/�&I21�#��I+�߳�K��f��W�ϾJ�ɨ�;��[m�v{K�4��7w7Rng�$�]��I$�-�|�]N��$��o���$[[׋$�����"cɖ8�
�v�jշ`f�l�\����\l]]\�Q�5�IG�$���K�ڞ�����>�$���jI.>~�,x�G��$r}�Iu;SԒW��g�$�]��I$�-�|�]]%#�L�#R'�$�{~ϾI.�u��I^[>�$����I/�L+�<r,�	����%�n�RI+�g�$�S�=I{�~o�����%�ҩ�M�
G�3RI+�g�$�S�=���}[o���'-��*���^��ߟ�|<~F쮘��v.�X7��pN�$�];v��y���}��yS��s�nј-Şz���98�*�qv�;m�=�u�X�䍓7l=��ڰ77���f+��nA��t���9D9��v�J����� ���]$q�F�C�Gm�
��n;yuţ��ٵˡ�<W\X�4i��6��k�R�v��nd(�)O� v�!h;\�cg�:�gl�7K4��-�a6{�@Q��m�~#3�=�=�"ͫ��K�2�s�%�Dj�^K:��96���Ζ�K�u��NY9�����I+�߳�K��g���g��6�^�>�$�~��~��2L����z�J������Y�$�����%��ORI.ӫ�0X'#r$�ϾI.�u��I}m�|�]N��$�{��}�I%ܷ$�&<j8��3R^m����䒩���I.������Y�$������X97rI��%��ORIw��g�$�]��I$����K����4��x��j8�F�����x͋=�����e,Q��x]j��xD�L��H����;~ϾI%�v�I}{g�$�S�=I%����"� �37t��m�����A ���	脀C"Q�2����� z �> +�6���'�$�S�=I%�v��|�U�u��a���Ɯ���l�8����ff~įo�4[�� �QF�D�A�#jK�?N�}��u���J&}ϯ �w=�c��2"G#�@�;w4g-���=}4�{^�p�ւ	Ɠ�i��e��F��Ws�Ẵ�2ݙ9N�[�2,�1�!0X'1G"Q��=�}�|�����7u��6u6��U�U6T�ʙ�X��y�'�_V ��X�k���H���G�`�x�Q�&����n�Ň�$��DBS>�x��n�\:),�^RT�J��wGLoG���h.v�����"�"I�,T���t����^o������߿���D�&rC�"�q�]	���$}�=��;=�֐{E 
��v),��J�����ޘ�������[XƮD�A��M��נw�0=�0I�f�J���VR�*V%�b�wGLoGL���f��Ɂ���@;��abNb�D�������o�9$���������$�h�@!$W��TT���<�������n�&<j8�)3@>��ٜ}�m���;w4�E*�1��?�����T=���Ib�-���F�S�r9��B��;��{��|e]]bJ��X�����0;�:`{u��|����׀l�w�ҹ���v�����w^,�BP��F�}� 7ﾼ��k�g�txW�9$i�3@彋 ?6��>IUl�}Xw}� s�:�I��H�i)&h{31.{ޚW��n�Ł����`wQEO+��eU�73uw�z[u�tD&�~_�o� y��y$� O��<BBCT����^2	@ �e<_�����X�I$��@�AJ9�k�ˌ��c�4���҅d��hh�Bȋ��d!)�T�8A�bD���	p�4�B��cU��5�H!�F,م�)*F���#���dh�n�pvf�Y����v��W���a��bb@H�"�Hā\��$f\�%�ь��R�9�5HU��C�X\�%�s��}��	������D��J�����~�I�SRXT`BIaca���ƞ�$X�[�2CX����%BR��VR7� �KD��B1#�*�$%T9�P�Y������o��$`��5�!L��wpaYXP��e���B)��1H��`�F-�hJ˘iA�z�F)8�(£�(�	+
����>L>C�,D�� _w���������UT�i
^n��	��#9nT`)s�l�5��`�b�u`�y�e8 �fh훊.kc���jqF�>���3p�����ѭ�Żmmk<c�-:-�tN��{n�]�fs`�ۈrf�2u� �N�ܲj��a2�@sgkUF��>�c��-�	�`ٍL��!5T�p�I�tH��z�:md�N�F��v��#�frX���j|��K��M����5e[�pi�r�m `�@;s��VFщ���8[Gm�n�Cq�fr�mk���ܫo"#�s�h`��&j��g/.���qq�9�]Yv�c��+���-����ڋ��ɴ��X�Upbܤ���K^��*���=�
��1rm�|�|}�!m!J���MÕ;[8��p��8n��g�V8Ӥ�K8uri7kx���N��[�����&��]*��lZ��:1�.��:�dٸ�g���C5>��;Wsm�"�<�J� 
�A���;3��y	RJ*{[���e�-�Q��87F杙�H\��2<�kJY���U��[E��<�ѡ�U�t\1����m��u�;X�P�Q����rN��6A��3ֶ��f&`m;V96�s�(ɬJܽp�C�}Y8w+v�p�f���Γ*��(��`N8��Ӊ��:�bn�H���)�̇:�����F�L˚��Ϯ3����l��1屯V׷v׳���QM�{U��R �t,��/=�mRÙ��e�mɹ���(�*��a	;hn�xt{l�=�*ݰqjT�b9e��ǭs�v[���u��=�W P���v�{ˢH�{g][U��t�Us�\�>W�U��4�j�c�j�.[���Y��B�w:�W�6�<P/3��ٶڮ.�C��۩4#<�6�'�����mn��ڊH��m�@2�h^�A�p4H��-c��㶹�sa��<e����ی�������.O��(��e�52v��������f3���uڷXF�[�0�tz������w���C�N �	�y���D� 8Q�p�� �D>�tW�������nJ�EcU�d����]�y�g���s�۝��+����}AP �v[lrRe������_}�M�vpuU�.w:8V��`��k�����-��֍k���qs��E�vlg�e�r�.:�^^��a�^�kd��Idxy-v8q`�Ƿ6�v�(Z-�୞����-a�L"�ۡi�]�\��>��Q�9�y�p���{V^�$:9�A;��w�w��˭g.��n����K�z [���͝N�Zg ���v)���{��\��\��tfi������}� ��� ?6�!��� ��٤����ݷsNI?{�������d7ﾼ�}�`��gBIL�Z|]ܫO�N$�����4.����߳��s@���4.~�,x�c�cqG�
"v�u`�ŀ{[ŁТg��xΏ��r�\Ֆ�K���w^,�F�{��������^�s���Hm"BS�f����(]�S����������[��6�̓9��ٸ)��r)m4�����}m�m~��ۚ����&�7.�wNI'��w��ɀ,=

�� 1@PO�������'�}�@�m��������zm�O ܂�G���wGL�Wr(�zH�r��I*Xb�V�0;�:`wH�~m�%	D�wu`ӑ�XJ��V�+����:`�&ܓ�h�*�H��b#��ې�7'5�%�\/5��Nlֹ�J��B՚�Q�<�T���լ �ۼ�۬w^.IDGB�Pw_b�6v�t�J��UW7WWx��X�X�x��n�%'WK�<�&D�2"H��-���;�ua�(�^Q
.�y���7X��lo�EM8�h{3?~V��f�s���8�k��{w �u��a������{����{���#��o����VDL��v\��]\��v��H]n��9��mF�n.���9���Z֮�$���1����zGL�D��r��YJ�T�Ŕ�,`wtt�ޑ� �"`m���&������+Yv�SzGLl����U��I�	�74���H�cƠӉ(�h�@��u�=׋R����
�(6[��>\΢����H��8�k�/{w4v�� ��h"ښn�ndi�q�M]<�����t�#[O��4NtA���[c˒#ȠE&L��H������s@/-�����%�^����mc�H�T��լ��,�J!L�ou�/�����֎�Rl0�7JI�yb`m������zGL	"0��Ww���Uj�bL���:`oH�^[4����1��&F8�G�{׋ �.IB�;����?��ӭ��"j���);�������K�̺�sW5���R�Kɹ;7d{kW=��6g��!ˋi,r^�tl�QiNA�9jy�Wm�U����}������f�e��dSX��XC(�L���u8^I[�.�.n�r���֛Fy���0pCi����ܓ��*�0����g��j�+�盈��������.^�8�ۮ,�zq�n�;4�ӷP�vܗL���Ӥ9\>�xtN(��/2l����ͦ@�C�-��ؽ���K��^�x3P.-�s-e�}���$�(�J9��{����^[4N�_�I_��w}� 󮟦n�U�U6TՅլ ~n�舉�e�V��,��s�bGWr��Px��18��M��� {���BUO��`ou���y�ɑ)����٠v�ۚyl�8�k�>��]��r)m5WV�kx�S����}Հ=׋~���?��0�;�{Q�(ֆ���n���s�Ԃ���d�b��V鿼?_�v�3�	�����^��� {���Hk�s@�����'�m�Q(��8�k�I%iU��`��`�w��
!L�{<�d�$�Q��[����� ��06�L`��'�WWx��H��X��X��x�[�J�-�}�V�)ɏ�N$���[f��Q��>��o�`��`������՝͸h661v㵮+v$�8%�W:�Eu;6�NpY��<�WL����1����zGL�D��Ӵ�"�$�21�#�;����Go�����4.����T�9�6�r�`��`���(��舄�(���䬯@���h�vɃa�I��ĕ0Io��wGL>��>�z����߱$���(ܚU�z�::`dL���]�X��ɷ��S�X��c�s\Z5�)8�rb� yx���ĤC�ɐHI�BG�{۹�t��M�0:�L`IFOʮ��U�J�b�N����t�����EV�)ɏ�N"'3@=߾L���:`t�遷��qZ1R��SW7wWx
%�>���X�|9 /EP�@J���wy$��{ٹJ�$�*Xb���;��N���f��{^�����$�i���0Vյ�uۅ�햞�ݢ2s�]�탪\�q����%1ȡ#I�π�����f��:cwGL	2ΉQ��*1�T���e��X�x��)����߱$���(ܚ^�z�n朢"�|� v�^ ���Յ+���YK1cwGL�0	�&\�zx\�1bNb�D���v��h�w�l�u�=׋ �P�(P����?8~��M�nn4�6A�"�ڡf�&5�/#�w]�lg�3���.uk��d�=�>.̠!��cc;<<�kV�`:�����\�B�LQ��Y8:���%��-���W�s�����z�Y����k���z���?���g>����+5�q���ڰ����4�jƐ9n��j�V���p�OY�F��U����E�/]��E�^�J����V��]��UUM�8���g��/7mΦ3�ئ�v77��WrrC�g���I	�5�5�DNf�}�Y�u^������GL����ѕ��*�V��� �z�&d{����ذ��x_+�X�%X��+K�0:tt�=$L���*.]�ĭ	5Uuk ׯ ~m����(�-����h���s$����e�u�X�x��IF��r���������qŘ:}����Z��5�a�5ŷZZ�9X�z��A5�m�~� �o�^, �n�>N��Z��uSt��� �oRL_B�;b�{ޚU�z�����sr%iS�GLd���:c�GL���dǎ<i�D�h-�@��@��gGL^�U�h��ĕZV�bL���:`l��l�07f���Ñ���dR�z:�;�m��֩\�Z�N^v�R�;���-P��Uͧ2Ō�06tt�6H���XK���&�LrG�6ԙ�r��h-�@��@�{w7ؑ��}&�8�e]ݬ �w^���KHJ�N2)�
�0��	���Wn ��H�,`�0��I0�c�
K@������ ���@�'��<MX�"� �WA�X���1���^P�@ �,�F�	JV�r�X�Gp�CD�H�H�Suj?���`d�b�:���?���=����`bF��S�qz'���8h�(tC�U���� _�
&*T:������ j���X"��TS�x�	yD(�-P�B��{� ��n�u�A71D��@��@�{w4^�h�٠v��e�1��$p�����遳����]�����g���(�/X��¦n�r��\��q�7�j�/<1f:�B��/-��h&��P`dL���:`m�&H�Lx�ƜDRyl�:�k�/tt�������ѕ��U�Z��`>n��x�䒅3�� �w^�ċ0X�%X��+K�0:rf ~m��B��DT��X�Z%��p�H4ێf���M ��4�����s@;ӭ�br"�#xIEYѵ��y��t���3�x�z�g��ӞE륃Mp�V,T,ı�D��1�����e4��m�by��#�@꽵�=׋�B���L,!I
HRB���x�D�,K��LɦɆ����ٹ��9ı,N��|8�D�,K���Ȗ%�b^��w��Kı=��r'"X�%�z~��L-�.��q<�bY��߯>�9ı,K��}�O"X�%��w��9ı,N��|8�D�,K���Mܦ�f�6ͻ��"X�%�{���'�,K��;�Ȝ�bX�'}��O"X�%��n�T�Kı4 p��F�!"�R#� ���P�XN���#fr���ӥ��i��x���6��W�·�ku�t1�GA{p�>�ܦ����wm4i� l��8!����Ѹ�a�����7i07�&EJN6-ú�T�:�i�-�-���2��[j�$���a=P�3���g����d6����`^Ŋ*ŋc3$;��n��E�ph������`��z�Z����]d�o�;��~�_+��]����r�Q��$�b���[tF�#!��+�MƊ�'i��:�7n�ۻ����ı,N�nD�Kı;���yı,O{w��"X�%�{���'�,K��,�w2nl��f�ɛwr'"X�%��}�Ȗ%�b{۽�9ı,K����<�bX�'���D�Kı;���^ۦlͻ�nfni��%�bX���eND�,K��{�O"X�%��w��9ı,N��|8�D�,K��3;�̐��&�n�ʜ�bX�%��{�O"X�%��w��9ı,N���O"X�%��n�T�Kı=�gfft���m��fn�<�bX�'���D�Kı;���yı,O{w��"X�%�{���'�,KĿ���\�sLл<�S8��Mf5��3�5�rp�	;OZؤ�Me���]5�����oq���bw�{���%�bX���eND�,K��{�O"X�%��w��9ı,K��Lκas4����i��%�bX���eNB��S����"��ʿ�\��%�|���x�D�,K���܉Ȗ%�bw�{���%�bX�罚m�f�6͹�9ı,K����<�bX�'���D�K�dL��{��Ȗ%�bw��*r%�bX����{�fnws7x�D�,�}C"w�v	 �w�p��	"~��`�Y�L���oȖ%�bw,��̛�&]�Kfm�Ȝ�bX�'���'�,K�����Ȗ%�b_;��Ȗ%�b{���ND�,K��{��������Fj���qq�C���O<�y�u���Gٰ���f�v>�1Z���{ı,O���*r%�bX������%�bX��{��g�2%�bw��É�Kı>�l��K�!��M��ݩȖ%�b_;��Ȗ%�b{���ND�,K�}�Ȗ%�b{��T�O�2�D�;ݟL�����m��.n�<�bX�'s�"r%�bX���|8�D��	A� ,x+đ"�`0��"tW����br&�]��9ı,K������%�bX��z\4�a�������܉Ȗ%�b{���yı,O{w��"X�%�{���'�,K�BdN��nD�Kı/ǿ�&3I��n�O"X�%��n�T�Kİ� �}��o�Kı;�}��,K���É�Kı ~�����ݓ�{]�lFF��"V�G%�M��=�N�M9�^��Vhh:��y8��Z�"X�%�{���'�,K��;�Ȝ�bX�'}���	�&D�,N�w�S�,K��=:_�����7n�f�Ȗ%�b{���NC�9"X�w�xq<�bX�'~���Ȗ%�b^��w��Kı=�;�̛�$��Kf��Ȝ�bX�'}��O"X�%��n�T�K�XdL�~�﷉�Kı;�}��,K���g	{n��6�ɹ�sN'�,K?�������Ȗ%�b_��oȖ%�b{���ND�,��b1R1�"��MD����Ӊ�Kı;٦wt��������S�,KĽ���Ȗ%�a>J�~�r'�,K����É�Kı=��ʜ�bX�{�o���H*�+\��sMC��:n�:��F�����d��N�9	��}��������w%��7l���?D�,K��ۑ9ı,N��|8�D�,K�����șı/����<�bX�'~ߋ��77ffnnf�ND�,K���'��U�L�bw�J��bX�%�߾�'�,K��;�Ȝ��S"X��ߌϝ0˻.��q<�bX�'~���Ȗ%�b_;��Ȗ%�b{���ND�,K�}�Ȗ%�b{3��Mܻ&K����Ȗ%�
�"g��x�D�,K��ۑ9ı,O}��O"X��*̉߯>�9ı,Osӥ�n�0��3v����yı,Os�܉Ȗ%�a��{���%�bX���ҧ"X�%�|�{�O"X�%��{��Oe��?��C���y&�[�c5�v�zy�z�&щ�Pe2���^yJ�T��&]�s�����uv�-�,f,	Zy�X�T]�.X+��\1�n����zP�� �6�qZ�r�4�����z�c�[-�]O^�t��Fڒ�Y�m�����b�[�1��͋k�"��鴇Y[
u��N��ۚ̓�X��T���}��w�s���&<��.ۤ���{9tgs�}s��݇�Ju�N�)i�7�����u��nή�3�w�{��7���~���yı,O{w��"X�%�|�{�O"X�%��w��9ı,O{8[�t͙�vM̻�q<�bX�'���S��P�B�bX������yı,O���r��&D�,N��xq<��"TȖ'���?�I�!��m��͕9ı,K���'�,K��;�Ȝ�bX�'���'�,K���{*r%�bX����3;ap�s6�ۗ7x�D�,� dN��nD�Kı;�����%�bX���ʜ�bX�"g��x�D�,K��ᦓ77ffnnf�ND�,K�}�Ȗ%�bw�{*r%�bX������%�bX���r'"X�%��	���~c���VX�ո�@�Cl�g��x:�s�8z�T�E�a�Mv/�{����/޹䍻���i�=�bX�'����S�,Kľw��'�,K��w��>�DȖ%����'�,K���߭7r�e.����S�,Kľw��'�������"X�'ٿnD�Kı;�~��yı,N��eND�P2�D�=�N��p�wt�۷sw��Kı>Ͼ܉Ȗ%�b{���y���Dȟ}w�S�,KĿ����yı,N�'{����ilݻ��,K?� dN��~8�D�,K��*r%�bX������%�`|,Ȯ����$)!=O<M���n��.�O"X�%����Ȗ%�a����o�Kı>Ͼ܉Ȗ%�b{���yı,N�3��̓2e�p:�n�N�im�.�p/Fϳ.5$�GY���9�{�}o����ݦ�ǻ����,K��}�O"X�%���w"r%�bX����q<�bX�'{w��"X�%��;33��3nݓ3w��Kı;���NC�DȖ'���O"X�%���~�9ı,K����<��eL�b}��\4�a�������܉Ȗ%�b}�����%�bX���ʜ�c�W����,(�B��)�6%���x�D�,K���Ȝ�bX�%���g]0�ɷw6��8�D�,� dO���T�Kı/����<�bX�'s�܉Ȗ%����"}����yı,N��Swi�%�ݙ�*r%�bX������%�bX�~�r'�,K��{��Ȗ%�bw�{*r%�bX�þ��ni���͌�c���`k��]���kX��
�X"M4��wW��}�pv*����1,K��>�r'"X�%���É�Kı;۽�9ı,K�{��yı,N�'{���,�t�f�܉Ȗ%�b{���y���bX����ND�,K�����O"X�%�����9ı,O����웙w4�yı,N�w��"X�%�|�{�O"X���>����,K��{��Ȗ%�bwٹ;�&�ni�7s6T�Kı/��w��Kı;��r'"X�%���É�K����*4�S�+��'v��S�,K��흙���˙�n̹���%�bX��{��,K��T������ı,O�w�S�,Kľw��'�,K�읻{n͹�̲������b��F:7/F���q	�b0���g��vup4�]vz鬬�;����d�=���q<�bX�'}��S�,Kľw����"X�'�߷"r%�bX���dϝ4�ɷw6��8�D�,K����"�r&D�/��x�D�,K��ۑ9ı,O}��O"|"�L�b{3�}Mݦ�L�svf�Ȗ%�b_�}��<�bX�'s��D�Kı=���q<�bX�'}��S�,K����Kٻp���7.���'�,K>��>����,K��{��Ȗ%�b~��ʜ�bX�ș���'�,K��R}��L�.�t�3w7"r%�bX���|8�D�,K���Ȗ%�b_;��Ȗ%�bw=��ND�,K��H�,H��"C�%�	� ���%�$�pŁ$є�B@ H@!#F`�(b�8���U��G��F1��Ј@���)!�d)R$� B$HT�X$R1S�B@Y[Af�Ѐ�A�1!0 �O � �P�%BA!HaYFhY
�),J�� B�0�E�#J$$���#�� b��X�0��eiIIB4��0�H�j����� H	 M`�.���S����1R B,�`� �C�$Cހ�"HM �1�X1�p7X$�b�H�H��2FH�D�D#a�ă,�!���fg�UUP�m+;�����ʹ�nI�M�m�"t�:J�iύٴ)��Y%*��+\��4��i:�ņ9J��Yf��i.Mђ���غ��7;�Yꇬ�'f��@��\kv:#;�"nY�J�&Onz���v{b��n����Y`:��H�@��;r�cUԫ+h�8�R�xU��ٶ�����Z�=����A<�\��z �ջ+��\�!Zl�����̮��.�۩kc�4�6(p!ƺ�+��U�5e-�]�D���M����p���f��/q��vܴD�,���&�kJ[NF�k���y�cZs��i�ތ�=�9Ԗ�pMgK���cH��Y�xC����=baz�u�������&�[S��q��5���-i��c�02�1�HY-�E�V])"w.��c����jv�ژW[J�D7��w^-�L���m�ƺ�REZyT6�UU��p1<��k��%䙙gf0:�C[6�� Kd�crD�mV[th�\�;	-���S�QWUn�M@�s�Z�,��;�������%��ݕp�x}Z�m��kk���<
����!I�y�܄�+a�H�A�p�9.�v��cg1�{M�<R*�c��Biܘ8㵒�[�I�\�Fh�S��$�/92�KOv�L�mf�9�Kvt�`Y�m�M&��Uw�.(+pm�6��J����rJ�x��㞀��4l����ҮS�����ݨ��r�0������]�d��^Pm��y��#�u�[O��-�lㆢ���]g]R�x����ګҼ��[]*4�j���vӍ=��*���%W+��tf66ᗳ�Zr9x��8���^�ݵm TY1`��.ʡg��p$�y��\j��ۜ���kV�ԁ�6ݕ���X���Vm�-4��c�0��ѱ��W,s�
��ƫ7Q�&�v.��Ʈ�h-U�ȝ�N8�Z��Fy��&�q�B��$�`	&��Jt�T�6�ŭHu��s�� ���̼J(�=���~E?*�D?"x �E�ދ�^'�(x �g�yo-�ҹ����KKr�!g���.���N��K�u ns`�ۜ�7P<4�7j܆"�'�<¸����9c&�'�z�<)նk=�<Z����r�����9��Бy3C����Y��5�%ԛnZ�Lm��:oI���CӷKrR�[4��ȼ]�"�M�:4��#V�3�,eT�l�S��Gu���feWr��T�[�p��j�!u�Y�{���o��@�������L]�n�/H�:�n����3��i�������{�b�77wl�˹�S�Kı=��ҧ"X�%�|�{�O"X�%�����?��[�&ı,O���É�Kı?����6M����]�͕9ı,K�{��yı,N�܉Ȗ%�b{���yı,N�w��"|(�S"X����Ϭ..fݻ2��Ȗ%�b}��r'"X�%���É�Kı;��ʜ�bX�%���<�bX�'��za�nn���6��ND�,� dN��~8�D�,K���T�Kı/��w��K��&D�{��ND�,K���3�L3rm�ͷsN'�,K��{*r%�bX������%�bX��{��,K���{���%�bX�ßL��0���w)we�Q�V��lI�얚�����;����;W=l����Yy�9Mݦ�e.����S�Kı/������%�bX��{��,K���{���%�bX���eND�,K�~=/f����ܻw7x�D�,K���D��lh����z~ S�?��6%���?�8�D�,K���ND�,K���x�D�ʙ��)>�s&d�K�L��w"r%�bX��~��yı,N��eND���Dȟg�}�O"X�%��}��ND�,K��xK�t�swv˹74�yĳ���>���S�,K��=���yı,N�{��,K��>�~�q<�w���{���;��N��Ĕ�=�oqı;����yı,> ���ۑ<�bX�'���O"X�%����Ȗ%�b~?{o3�sn�&f�r��`���[�:�k����oa!v���k�Map�s6��fnq<�bX�'s�܉Ȗ%�bw�{���%�bX����ʠ_�6%�bg����Kı������m�]5��g{���{��2w�{����ș���J��bX�'���gȖ%�bw;�Ȝ���2%�~=����ܛt��w4�yı,O����Ȗ%�bw?w���%��_�V�q�"w9�Ȝ�bX�'��|8�D�,Kٞ��n�4�d���7eND�,�QDϽ���yı,O��"r%�bX����q<�bX�'{w��"X�%��?��v���n]���'�,K��w��9ı,?������~�bX�'�]�T�Kı/w���{��7��������")�aK���3��e�:�+�x����v�X�'sv�]�]�%��&m�Ȝ�bX�'}��O"X�%����Ȗ%�b^��w��Kı;���ND�,K��xK�t�swv˹74�yı,N��eND�,K��{�O"X�%���w"r%�bX����q<����2%���r}�&�niw.�fʜ�bX�%�߾�'�,K��w��9����b}���Ȗ%�b]��9ı,O};/2u�6��ܻ%��'�,K��w��9ı,N��|8�D�,K���S�,K��*��EC�ؗ����<�bX�'s��͐�M�ٙ���nD�Kı;���yı,N��eND�,K��{�O"X�%���w"r%�bX���?����*їb�k�4p
��pTf�����h�vnQ�fl����w�����y�N۹���%�bX����ND�,K��{�O"X�%���w"r%�bX����q<�bX�'�=����i��wwnnʜ�bX�%���x�C�U�L�b}�}��,|dL��{��Ȗ%�b}�ߥND�,~�D�}:_�����ܻ���O"X�%��}��ND�,K���'�,K��n�T�Kı/w���%�bX��N�s&a.��&Lۻ�9ı,N��|8�D�,K���S�,KĽ���Ȗ%�bw;�Ȝ�bX�'��7$��ݶ�M�8�D�,K���S�,KĽ���Ȗ%�bw;�Ȝ�bX�'}��O"X�%��>D���r�s.��\n�7$�$����Z�=(�ʩ�����[ۛvۤ��+��=[����G N��k4X{q��vzgY��k�w=;e��˵�;i^.t��f�v�SOQs#�w]c�㵁�����������΍n��+q�-�[b:�]���vz��C��%G����r�;v�݅�i�֩�}��.b6Hɺ��p7���-���M���r��D�����Msq��]/S�
F�'s�OUҹ�B��轞�kN;��Ŧ�v�n$����7�ı>����Kı;���ND�,K�����؛ı?���J��bX�'���'�m���t����%�bX���wjrȉ��,O�߼8�D�,K߮�*r%�bX������'��L�bw:_��4��˙�nf���Kı>�~��yı,Oݻ�S�,j�lN��u9���wj�	"zy�}p�f\�nf� �|,�{��ҧ"X�%���}�Ȗ%�bw;�ݩȖ%�bw�{���%�bX���;Mݦ�L�wv��Ȗ%�bw�{�Ȗ%�a��~߾�ڞD�,K���'�,K��۽�9ı,O;����\�6f�M�ҳ�&�gX��܉����!s��5sZScY$�b�&�\̙���%�bX���wjr%�bX����q<�bX�'�������7�M�bX������Kı?����I��sG���7���{�?~�É�6�.2%�b~��ʜ�bX�%���<�bX�'s���ND� 2�D�>���$ܓwsv[�7t�yı,O{w�S�,KĽ���Ȗ%�bw=����Kı;���yı,O�����7$2�r��l�Ȗ%�"���{����%�bX�g~�ڜ�bX�'}��O"X�%��۽�9ı,O};/2u�6��ܻ%��'�,K��{�ݩȖ%�a�������ı,O{w�S�,KĽ���Ȗ%�b_���ɗ <W<;74����Glƺ�2��k�50�)�mn���oWd���]�\/��%�bw�{���%�bX����S�,KĽ����'�ı>����9ı,K���gΘf�ۦ�۹�Ȗ%�b~��eNC�9"X��~�x�D�,K��ۻS�,K���É�O��Wq6%����۴�	�3w6f�Ȗ%�b_��oȖ%�bw=����K@�D���{�É�Kı=��eND�,K�~���r����]���'�,K>��ۻS�,K����É�Kı?{w��"X��L��{����%�bX�e'�]˘Mɛ�ɛ���9ı,N��|8�D�,K�Q����T�%�bX��~�x�D�,K��wv�"X�%�v�.g�e��m��h��mnXq��'Թ�뇡�ktu���;=..9�]�j��������bX�'�n�T�Kı/w���%�bX��{��>I�L�bX�7ߖB�B������:�.�U��uW��*r%�bX�����y��DȖ'�߷v�"X�%�~�~�'�,K����ʜ��?�!������_���`ZKa��߭�7���{����UND�,K��{�O"X�%��۽�9ı,K����<�bX�'{�.�f���3wnn�ND�,� dL���x�D�,K���T�Kı/w���%�`h!�*@OD��H���ۻS�,KĽ��3��e�n��̙��O"X�%��۽�9ı,?��������{ı,O���wjr%�bX�����yı,N��Ojy�Dr=��XIn+X�l</,e��GpRl���vԽ*dꎹ��fnʜ�bX�%���x�D�,K����ND�,K��{��~��,K߮�*r%�bX�署���.�r��n�<�bX�'s��ڜ�bX�%��x�D�,K�n�T�Kı/w���'�������K�����E�:��Q��{��7��/��oȖ%�b~��ʜ�bX�%���x�D�,K����ND�,K����vK�n�n�re��'�,K> H߯>�9ı,K��}�O"X�%���wv�"X��2&}����~����{����4��m;s1�����bX�%���x�D�,K�G�Tk����ݩ�%�bX��￷��Kı?v�eND�,K�����}������8�?�܍��r�յg5���\�ͣ����l[�V�gۖG��V�T\mz�GCm7=	-H�;�G>�kG�U��9���[i���uF���0]Eb����x�Hu]X��{�ڸ�����Si0�gOMrJDg���sk^�%��V�X�7��-�jm�[<�P�V��Y�XM�=g��vwL{t�	.��٤�u�à�s�<�6�*Zu��n��<>�M�'F�T�B���\r�NڍW)��^p����[~����,K���ݩȖ%�b^��w��Kı?v�e�U�DȖ%�~�﷉�Kı;��f��f����w37v�"X�%�{��'��H�L�b{�ߥND�,K���oȖ%�bw;�ݩȟʉ�2%�~��3�L2�M͹3wx�D�,K߮�*r%�bX�����yı,N�{��9ı,K�}��<�bX���i��i�ə��3vT�Kı/w���%�bX���wjr%�bX�����yİ>	�=���S�,K��=��ܸawt��w3w��Kı;�����Kı/}����%�bX��w��"X�%�{���'�,K���?a�Ǌ�N.ۤ��K�=��^S�}8��'�e�p9��#�����?��ws}�����f��ڞD�,K����O"X�%���{*r%�bX�����*�"X�'��ۻS�,K��{��n�vL���nL����%�bX��w��! $ ,@*�"�ʦ9bX����x�D�,K���ݩȖ%�b_߽��<��(�S"X��7'ٲnHf�ݹ���*r%�bX���}�O"X�%���wv�"X�"C"dK��x�D�,K߮�*r%�bX��Ӳ���Lٙ��vK��O"X�%���wv�"X�%�~����%�bX��w��"X�� ���bo����=���{��7������ݳ���R�T�Kı/���x�D�,K����ҧ�,KĿ����yı,N�{��9ı,O�~��2�n��ے��p�k��7e�V݋�x:Ķ�Bu�ϖs����*��O���|�y�t�0�_�����X�'��J��bX�%��{�O"X�%���wv�"X�%�~����%�bX6z{N��L2����weND�,K����'��@��M�bg�����Kı/{���<�bX�'���Ȗ%�b{����ܸawt��w3w��Kı;�����Kı/���x����G�S��T���*��R- ���`�X�A��U:�`�	`�+Hj�'�	$S �"fQ�"S@��AH�+�0X)�Uc-#Ω���3[LL�����$�h�,Y,H�"�#���nI33��l���9@
�"��E"� #�?$U��>b�@�b"�@�?���UB��� �D���ȟ�y��ҧ"X�%�}��w��Kı;���ܸa��4ܙ�wv�"X�|*��-�������%�bX����*r%�bX�����<�bX�'s��ڜ�bX�'���gv˲f��[rM��'�,K������bX�� *�}����=�bX�'������Kı/���x�D�,K��.G���P>պ\mHpr$4�m-�jY��x�ʿ���ndd��$i:b-c�D�,K��﷉�Kı=�{��9ı,K������"X�'{�p�Ȗ%�b{���\�n�͙���d����%�bX���ڜ�bX�%����Ȗ%�b{�s�ND�,K����'�>ʙ����n�0�3ss.�fn�ND�,K��~�'�,K������bX�%��{�O"X�%��{�ݩȖ%�b^��3�L�svf�f��Ȗ%� �ȝ����,KĿ����yı,Os���ND�,ABx"���" � &%O̉}�߷��Kİl�}N��L2���6�9ı,K���x�D�,K����S�,KĿ�{��yı,O}�p�Ȗ%�b|��ﳿf�晻-7fC6Y��1����n��c���t���H�[/������ޯ��ܸa��f������ı,K���wjr%�bX���{�O"X�%���9ı,K���x�D�,Kܤ��r�n��lͻ��9ı,K����'��c�2%���~�9ı,K�߾�'�,K��w��S�,K�������vL�ݶܓsw��Kı?v�eND�,K����'�,~�Dȟg�n�ND�,K��~�'�,K=����w�m;vkAH��}���舄�����y�C��.���x粚-˭��c�nF�'&�U� �J"w__�=����n�P�G�I�fR2��̻�Л��6��o�)����oh{V!�)�Z���Y9J��V�:�������ۙ���B��o�f��C]�N�7X��[v�ΰ
g�c\v�S�n]u��ӯ�!���g����=v^�L�u��=��w\ה��4[����oQ�6�6��R)��k�q��+�nFnl���9��7c�ݮ�iͽ���{�� ��
K�j�]u͔��Ѷ�8�@=�\���搀.�H���L1�㍩rO�;��}vـ���_�:y�� w'U�J�V�1fbI0=9A�{dL	s�L}���EP��ҫ��U*�� 5���^��>���}��;� ���܉������4?�������h^�hܶhwTi��#S"R����x�>���|x_�^ ��ͷ��~[�,9V]�M=:��al�<�fcR��<�>�X��p��>�4b�j �X�Ӕ�D��:$�7z&�}+�c�('p��l��������D-C,!#50�/�-��z�h^�h帵�ڌpm��D��*��h9�4�f~K��ƀs���;_q��x�8�jFܓ =�w�~{l��n�9DD�s� �N���"캻*��� ��ـ}��}��_���D�<oEYE%��9���g�ؑ�����d*F�G��K�^w'$=l�+*;^��nׂ���~??����wx�k��Q�C���]WǑɎ5#rh^�4��ױ����tB�Jd�h�J��m\�sww��� ��ن�	B""����W�M���d�"I0�MI(�>�`���/]��DB�ݾ�<:y��1�'p��l�%Ή0މ����v�,�%�;������(�K�=�=��KF��u�.yׁ {hh��K��ww��\|����'C_����}�� �����=�&L�̧hT��]�U]�U����3�"S'������w��Q�C�:��T��r5�C@��r٧�g�߳����{g� �s��Lx�I"q) ��� r�����0F(������	� �TP�/����>\�Ȟ<�Lq��@��ɠy$�-ל~�� ��� ���]��TNDᕘ��/)ʹ͌�Ү�����뜧&H����0�Ab��9��)$�9��h��0����B��J"���}w�nW��@Pi��I�nײ��-���� ��َ#�B�Tj�u*�S9X^� �������@{ڸ`{�P�9�qki�Q��k"rh^�4{m����
Ϸ����R�Ef*Ėf%��&�(0=9A�{dX��� �
!+I/k�����S�3��lWC�'�V�z��֊QLnM<9��Ǒ�7V�k�`�k���ڵ[@��c����g�7]`8G��퐄�I�p�#Ŷl��}n��vyU� �]C����t��E[�غ�����������Iѳv�=����k�ю}ղ�ۑ���:��pe&^� �l�j��<m���l�9��\��\�֔��\�.y��>����4�\����8��	�'f�k!ɮ�v��9x�$�t���o��/޹�u8ڍ�!�/��r٠U{d�9�P`��YJ���$��C �Ș^����f��:S#����)��7SwUw�t����fB���%�Y�@9�zhwE���F;���J��QM��~����n�
�l��ǝv!1�#I'��h^P`�\�w��UY�/�Nn9�c���s1b�8zS������ٝ�r^�g�S�ζ���V����+H�Q�?��\�w�����ꖶ�Q4܍dNM��&�����ޔ�P�&�0s�0�������Y�<s��ҒM�즁�즀}�f�U�@����<&H�j8���S�y� {{� r���l�ճ 9���a�5�H�JC@>�@�(�(����}���ٺwvZ��n�"�T��0�:�t\]>+j*��4Q��i������x��)k����&�(0=9A�{dL	}D��1cs���h�e7��9�<h;�M��&��q�]�Li��I�n�� ����$�Z�#�%GЅ<�P|�����@�D�H���"�7��{���?2����S!pnؗ;�M���h�e4�e4v�[M���jA�'&�U��9DGТ��~����n���������974�ɔ�4�d�U��0nP� �i�T���m//Wny�hW	$����(0l��߫�_��G�߿LxL��8��>������^����f}	$�CZr��V�5�H�JC@9�zh^�4���w�x�9�<h�+�<x����I4/]��m� ��ـ��JP�������
���xKGq6��Uj��i$����(0l��.tI��>�\h`ۍ�p2G#�l�L8��7P[�q�S�\�{Z���������F�!w����� �Ș}"_UW�;��s���<1�Ӄp�?�;�O�����9�M��M����=���CQ5 ��@����9�M��M ������x�'"m�I4>J�� �;� ?y���"z����G����$q4�}{)�r���wx���!%��!D)��H@� YX$)Z�D��$�E �)1H�7�#B ��&T��RIeF��B��X� �:'� B���X��DbA"�V0��	$a ���|Ņ��GR9�t��zh�"�o��!H�H\єb� �4�&l)�� �b��B��Xʹ(~���HDՂ�Q��+3.�Be�� I�jb��1�{��,)IIa�K����{�wo{��{�G�_�UUPQ-���v��W.��qK$�{f��Ni�]�9�0�;Ha
k�oR��ܸ�^�I��01Z;WI�}�4����2<�W��k�)���;Og��w�[�9Z�Ƕ'�4vז�����*���vg��-����շ,RJ�Gd�v��z�u�RA�M�ҭT�Qv^�ລy�5g��e�+a݊9�Km��Û�k�d��Ή�'�W�NkG%�cR�5�R�����3vڕ���0R�K�p�З���qZz���H����ؔ�a$�A^.L�q������\�;��Mmմ����l��; �hz6$v�n6,5�48�Uv:�����4Y��ű���t�T�^��C,mWL[,;��A!;�쯝V�n�K���v�GZ3�n9��f�@Q�EA�=��ۂ�f�5�dj�m�0[.��e�Б��ky�Qa�P�l.�a�rRA���iN�
I7+A@X0P�]Y��vعt(��k5�Ӆٝv�v�E��G(q�a�@n1�z�Q�s)��m�&�b�s�\�����j<3���3�a�{ ����ݮ��{5ā"gD�z��rmd�<o:o�6*���d��k��kp��GvŮ����-�3͞A��ŭȅ�uF�L��,�v�Vx^���nG�4[.�}��҈"]v�\���=�,Wjٻ9=v=�.㩳�t�e]�
܅k��p��絻V��iÊ7Gl���j�S��.5�yn�Ӕy��Zigvy���n�xJ�t�m�cK��Uڝ�Ùۆq����ˋ�Utm�*�v�Y��ݶ����"í�p�n=CF �V�V����-��u@T8�tj�4�%WC�^S�P��JK;1tu���k�.��+̗9��I�lP`���Fڹ�������2J��i���`6,՝�KX7l8��lY*mֆ�k
���\�YYQ��&�mڙ�,�D��n�S<mn��[�=��͐
^�Al�V�E�펕ggt�]jv�\�������x��5wT��U@�E�'��C�aOu(�?��� ��^O�6gm2a[��%�P�;�]�j�jyR��`��m���i�w[�0Jp�7#m��5ݎst]q�qvC���&�E7&^ӯn��5�Y�e��aTmદ�a1z�ޓ��������^���-�.!�Vq�)^95��:{x�xJ��hѭq�4��=��l�\rf����E�.�v{c�<��PjV��q�q7v�qT�|�nfy�M�ٮ�ܗ	wi��b�3��x9mf��Y٦2�↶Ԭ%Lr1�Y$�Ĥ(}�4
�l���Ϣ_%���� ���)}WsJ��T,J�L	s�L�P`zr� ��7߳3�G���Q��nc��M��Ӕ�D��:$��nWdVM5wS34����"��q�����wxD$�w^q�{�O��i
��Yx��0l��.tI���NS}��??k�<�Zc��<\S�9��r�.�P�έcWg^[O/jt�Nn�9���w��||��5�'�����4s��ײ����;�M���y��19lRI�O߽��x��#F���� �5�H����G�}z`��^ ���P�B�9I��{�Ǆ�DM8h��4�[4
�l�9�M �:��dǍd�'���n�>n� ��ف�
��y��?�9ǉɄr)&�W-�@�;l�?n�0��������U�]\�wޞ5mn�nr���wk��cOv˭ۂ�$�Uj:<����{�}�k�E�nn��W���_��vـ����(�!ӽ�x�^W�Ɯ�$�F�}��hܶh|���m�>�Q�O2�갚B*컚��� ��^ �����G�BILL)�$%b��.���|`���<��I�?&E�RM�[&��vS@��l��(_%	B���׀o}t���V*�J�0X�`n����"`U�d�9zF�JA�����PF]ѝ�WѺ�6ݴi�۞5j�u�q���_�{����o<xL��H��[<hܶhr�4s��˝X�2cƲI�H0l���D�����r���UW�H���眉��r)&���zM��f%
ϛ�0��x�Csu5���,1,I07yA����rJ��EGD@��C>�盼����A�#I'��hw���-�W�M�즁�W�V��O���D⣇����"CM�>�&0���Xr�y�����〞Gm��> �}�U���{m�B��Hy�� �}�3U7E��w$�� ���™ɺ��� ���9%B�To}t���*�5w5TM�� �_��������}�4
��n�x�#�q�!���w� ��^ ����r�	/�T�~����X���5�H�JC@>�@����u��7]�~ݶ`
r��%jH � �*��ygd�>vٹ�m��A��rd�qV$'���n���A����޻*cՓ�J69P��tS�1������h���VҘ�v+;HF��u��Nas�wmga1ju/n8z��[��S-��z�F�fѡy�	i�$4�f��6R7,vi��7^�^�;Y!����]IM�-r��tJm\6�tu�l���9Α�{|��=�� 3Փ�;�u��nF�c�qX�f�@�G�)6i^p��Y9A��zhy�z+J�P��$�����?�z����y\=�h��F9�@�;)�{�A�{dL	{"LV�Z2�,���Y�`{�A�{dL	{"Lޔ�>���L1����� ����H�w��P`l�0��Uf\Q1H�$�*�h�f~������x��l�9B���m�Q�<iF�����f�ɹ{^ћi����r�F���:pu��ZH�+ZJ�0X�`n����[4
�l�Eηq��HG#�l��}��h�r
��(�����<���=�`��T�V�U�I^+���0%�07yA���S@��y\���r)&�W-����w(0l��/���^Xf,.�,I07yA����0*�h�R�F�4�<Q�I�����8N�����K��\<���(�N�m�t=V�4�i$�7��S@>�@��ɠs���>���L1����h�n��IL�w�� �w� ޼X�ۡ6�!�A�D)&��m�@�;)�� ��"�Au�}߸rI9o��m��9�H�drM��N���D�ے$��N3"�*�R�bX�!�'GL�"`m�`s����[1�rF�9���OOnؑ��,�p�+B��k��D��GJ��pL:��*�ˤ���X��{dL�"L�P�-���U�Ȟ<�	9�@ے$����N����}���]�{�jQ4�H$�rMݳƁon�}�f��m�@�9ٖ@Pj4�S%U�
B������}x��w��?���A��@C��~4Q�a�8�m�&hܶhrD�������t�YbV������|aH�8�.!=��M]5����^�v�6,d#s����ژ��jD'' ����� ��ـ7��������R����%y�,I07yA�'GL�"�8��o��#�o�0x���$�Hh}>t�=�nH�w����a�5	"�G3@�rנq[d�9��h{3�}�h��<�OH�&�%��"L�P`v�ײc
�*v[$=�gvS-���.�nW5�KY� ��#Oj��gY�v�lb�vb����Z��+tL�e;b3��OFCƪ�1n�c��q�N����<����v�gѥ��t3�u��s��ۮn���r2��kH�Sn5�8C��m�״��v��@�Cqu=�0��f���.�!���w42��lWS��A�i��!�������[Ml��Tͺ>����������2�d�2�9��;�ԭ<V�rgA;��DN�����A	�ά7w��� �m� �>n���?H9����3��NF�O#p�;��h^Ɍ��&�(0=�WLAx���Uf�|�`>n��(P�����}?�����9{+jbi)jLI�`u�07yA���^Ɍ�q�v ��ND�#�h�e4���߿DDs��e��`>n� ?l�v�ʻQ�T���4�닎n
ԍ̈́��)�)ء�P��SƬ�]��F�m���A���1�ײ$������"+L2��۳n������qA0 0�B���<V($ �	��"`����
�~�r���~����ߺ�0���J�wO"�M�QJ��U��`w�� ��ه(��/]�z{�=��Z�O921�������$��������{"LV� G�9By���vS@�rנur�4s��ܨTm��bɎ3$M6�l;gJ;��.�L�a�k�W���ԣ�=��a	�\�q%���8��=��$���o(0:r�^e�����-*�K{"L�P`v���f�33����o�x�'"nD��@���9$����Ʌ:���)$*�=��+�t�RFp���S%F�"�XQM<�J�����0�
J��"J���X(E �*�7�<�0��<�P�eIRr$�1�XR A %�B�9�d"�Ȏ�%@9����W�
�O,�8�%"ĄH�S�$�ĒG���=� ������<�UX '@C� j�����!΀'���Q�r +�}��m�=�I?_}�� ��ѻ��B8���w���>�n��7w��	$�[�0y9U�Xee�%hV��������`or���f�ID'�r��P]J�����Q�s��:iԊYI�����SS����H-�O�H��G��I'�U�zM����m��СB^�9���<�����5��a�bI������;dL�[&��r̲x7$HO�w�l��w�%�L���y��v�	�#�6��4?�ff%{�M�����%��� �}�72�rۻ������������T�ￎ���h�@���0mbX�3�ni.�s]s�n�R=�c���R)��'U6��A<nL1��8��'$�/{)�v� ��`�j��d�FU�]��*�� �m�>�B����}x�w�@���g�ԫ="��I"���׀��âS=����� 9�pyT��$x��I4?�3?~��=}4�/�o(0	�����^U�b�224��?�n���n������y��I:��"�?��/;�����r��]�msl����qHݰVZ�g(k���ú�s���Нg�v���@v�t���m��]��%q��\�X�Nn+v.-�$���s��G'X�v9����v�x{���N�|Ǝz�n�;cV0�p��6Kn:�6=k��q�=��#V
�b�\���m�J-E�xۦC�	���ݛ���y��n�؁�d��5�/�w{�z�o�����,
b�:Z�LX�C�rp�m��m���hqֱӇW�pg�̒x4������e4�]���ġ$���|`e'�a4,Uw��bމ�{�&�P`}��h;n��Q4��5"Iɠn���هBQ=�ذ����w�y9�ܚ�ff/v��/�7�`�d�2R�*���UUf�vـ|�"����������/*��)�q���bO�G4����ѝ�c5Jٹ�$��Ʊfm]$5q���<k$�8����^��@9o�����y�M �W*���q9&�|��ZJ��%iB��Q&�_�|`;�4��jQ<X��2c��4=��`���s��� � � � ������ ؃��A� �o~��x ������� � � � �;��d�&]ݹ.l����A�A��"����ӂ�A�A�A�A������ � � � ��w����lll{�>�|������;�l�$ɹ��fnl���lllo������lllo����A�666?���N>A������� �`�`�`�����fL��En�3��R���E�]��0[\Ṩ�u��鲝����wwn����u��R�< ��~�x ���ϧ �`�`�`��~�Â�A�A�A�A�=���� � � � �=�����d����fn�A�666?���N>D�"������|����s�g �`�`�`�~��o"(� � � ���fgƓ�n�sg �`�`�`��~�Â�A�A�A�A�=���� ؃���B�]A�A�o�}�x �{�>�|��������v�e7ws-�� �`�b�� ������� � � � �￿���A�A�A�A�߹����lll~��xpA�6667��Y��̘n�nM�����lllo������lllU_}��N>A������� �`�`�`��{���� � � � � }�����鉁ͷ��vs���˻k�X{y�nب�A�3n�+5�b9nn�#_��lll{��N>D������� �`�`�`��{���� � � � ߻���� � � � �=��۲]�77s&dۛ8 ����|��`�`�`��{���� � � � ߻���� � � � ����pA�666?�4�ٲ\�&��7N>A�����ﳂ�A�A�A�A�wﷂ�A��"A ���s�pA�666?�xpA�666>����2�]�mݙ7$�����ll_���A?����>A����������lll~��xpA�66
�dȪ�N�.���>A������A�A�A�A��o�g�C���fə��� � � � ����pA�666(E_￿�A����������lllo������O{ٹ�����N�Y:�Wm\c�3�����^8�s^�yu��G���}��<7T�x��:`m��'H��A�N9e�@x�I#a$4.Z���4r�h�e4�q���$x�$����x��|�9|����9}X�Ԣh��FF��9e4w�{&0t���تb��bĳ	�sV`ݶ`DB������x����P@��*$`H�z�om��������s=�>oUu]���š(�f�)�[�=�ѹ�(�؃\�vhḶ5�5n�|sn���ev^��Q�����`[��6���ۃ<V��#Պ��n�L]µL71��v:�;X��m�L�=�`�G/)-�̇X��{HW��=ŭ��xv�:�Rg�,Z�\v���l��[�n�N����}�odyΈ�f30#�
M�2e�;�˪�����(��n�B��%����.df�vZ�[�.�v"?�����c\Ͱ��+����c �H��A����n��Q4���Ĕ�@;�f��e����/���qr׼HY���y93��07b�g(06�L`�&q�w&�$I��4^�h��l����q�Q+A��I%�	!�ײc �06r�g(}��~��ǆk+����Ч���n�k��`(���f�B�"I�헑�2E�j����"`l��P�����=�h��FA�4^�o3�""�%
��|`w��|���ՙ���4^�h\����{�M��Ɓ�v�	��bQ8h}.��`���5� ��f�����M% � ��@;�f���M���W-z�ffg���R7 ��,=���f�@�덧��� �esV���1����12L1��N&���Y�@�즁��]ϐ��;���0x�đx�`v��wc �06r��$;s�(�I I���@���w�#R�8&�=E�g{�4�z�XȤC�$�$z�n��`{l��B������V ��5�nc���/;)�r�S@���@;�f��T���0q�F����w8�ŭZ�e��3�)b+\�[v]<�"�㑶�F�r�S@���@;�f�y�M�<�pG1&�X���밝�Ɂ�E������SLPi))�z�[4��06r�^���Zʼ"���^%4M�� ����m���X(��@� H�
��=���Q�}6h�z��&�#Ɯ4^�h��0�o(0�(X�W��:��^��
7��͂��ma�u�բN��S�'!""�‱����*�k��٠^vS����4���E"%�w��bL�D������/{f��p�(��s$��7&�ye9A�N�l����*V�,If^R�Cg(0	� �0',���v�	�#��C�{�l��6(06r�S��TU�J�j�l$�J��*á�9�X��%�ag��Ԙ�V RD��31ъ��l�(A!��}@(1&$�0��� DZt�hh'C��F0c� �6ѫ��tX�aR$T E�đ�`��#Q R\�@��1c � l
P���"�HD)���@c#ŀD�Pq��CLz~d'��B����)f��о��{k��=�[}!7�jAX��Q�#)A���
�#��H�Ç��P�ŉ �#�����wv��B��������Y0�c^��r��մt�����o�{R�9 ;v��lEj8�2:�m�L+(��y۶	���oY�<������ss�r8{l��3UCru���pU���ӳ�8��h��+�/��N�P3v���Sz�����@l�c�f�jV���G����I�;f��{l=��	��90���ܣ�%ɇX�=�5�Hsv�l6���n�u��v�����^���t�^�����,����O/2uu���x�f�������M���uɛn;���y�N1l͎���3�nݹ35��R��[�-U�=���y]��F�ݚ��*ѱWJ�\�������>E`���m��M�I�5�{$؉�ζ
�öK�+�!�<V��[P�@(Ѹâ��W<��܄�-�nruG n�kb*�V��I�ڥNdv��&Г!K�	��e��ZD ���x;��v\���tm�q�F�m��IƲ"�m��}��@�����vˊ{���B�6�م3\T6ヴC���}�A�5��e�\��6��.����I��^mbA+D���';_nul|��{��y�����n�B��;I�c��h��&�;d�q�n�O;.T�#��atZN�ŋ�}�	���h㗮���m��[�ɮ�^�ʮa�;W;]g�<����LLpW�\c]�q`�e��1���L[Kݬ���Ui٧����M��qШUX'��#v��=/\���cawj���T���LY�]�(vhaƶc��<�iK>��I��[`���a��HQ��U�"��(u������K�z�I��݈dIy���.�ͳ�ڞ��@e~X�9;�L1m�g$;\��$m��[OW:�i)Eq�ɍ%lCf;u�؝�m����/�dG��.�kDY[gf�B���q�:m���'+���h�秶ڑ�ۚƋ-<�.%u`x�k"q���h��"�p�� �� �&���Q�.�j� �
�q�+���*�
�D���e˞��a�z��Y�]���컬���o����yEz�n��ʑ�Aʃ�`�bwk���"[D�%�����n�Z�p1l���z��,kd���h�h�;�qĩ���g,m�|�d�WY��*-��w��~�2(׮ݶ�5dra��F�*�m�{�\']K�I�m�C\7$sR�]��ãՅ�V�V�du�^�GZu�-,��6��_T@��9�3��ݻ�l��9�i|`B�u�bw��U]W�|X����a�bۭ-��?|4���b�(�� ���h�S@�즀^���q2�1��N&����3��)�y�����n󒈉�T�ʮV�UV��U5f�� �]��2y�^��� =6S�����$���;�`�lPa�����@)�dR!�j5$����(���������� ~u�̨�]�.`z(�dv��l�7m;j��a�Ol5they�9y�PF{-�	#L	�A���\��"`{C8v�U������uV`��3�!Z!R�J"�"">J*G?gՀ����g�'����LĚ$p�8�|��[4�9�M��m8�JA�@����
#������>����fx�V�ޏ����y9�nM������-�{dLL����W&n
�p��H���p7@<ݍt��/sH�pǇ��l��l��y.�#o���ـ?V���n�BI/����eY��H��Š^>ՠw�h���;�ڴ�ʪ�D<��mf�I'����'��{9:z�D0� �.P(�#�0�
#KDDEVw]�y�9�6u�ܔ��.�jn���9D}�Q[�~��9��`��Z���K2G�RIdn�m��"5��������l��EM�LlY1��JI#��;g�w)�լFq��76�5c��*;1������5�Ͳ`��$Ӎ��<�|���4��hw���j�ӊ&,RS	#�ۮ��L������ s�u�k+q1���r'ܚ�e4�d%
g�_V {�^�G�SV��ws4����Kל`:�����
Q�aQw�������y9$�}=�q@Xԑ�1��v��3������=�<h�e4G�#�8d�FԘm�*���[�6�a�R�ٴ8����r��b�<�(�C�&�#�@>�@��w���0:��.ՙF*I+V��� ~�f|�&M�|`:����������?�&<��F�F�w�x�%�L`�o(0=�WLAx,Uw��1	{��D�����hs�6�Q4�RS	#��l�9.ל~u��k��%
)��{;m��,ϡM�L�5��v�a�Tcq�u��i�����u�8�u��-��Z�3���]m֏<kȡ���>�p�{S\��d��kl���f������7��o�ב&kvD(ں^]Ŗa=ћ?~�zzu�U�]׵&����:5�W�-#؋)ndʭ����6�:����l��֮*kˁ�f1�N��aۀz��vi��sl��6CrGL�ꫡ��w9��@4�p��:��3[8���#��sy;�!��kQ77����۞��_�?��|07yA�/zc �Șf�̹��I"s"p�9��o��]�z���@�즀Zueq@XԊI2)���"`zr�w�%v�)�G��H���l�>���=�`""!/���Հt�>�f�U��B���0=9A������"�m����Vϕ�狴s�Z�g��T9|�%۱��=��سl��r���mq�.ի��b��Fb����ޘ�=�&�(0>���LĚq�h\�{����>P�!}�������?{m��9�i��K Ҙ��@>�l�>���>�e4�v���1���r&D�a����0;��`u�L`������I#r�@�;)�~��|� �}�}{)�^tQ�E2'L��f����v�N׊�����Vш.([nI�4,�#���$���:����[4�e4s���ǲ��H��<O,K0�LNP`n��zc��UC2I�nM��M���rTS�T���p�SW89��j���sޚ�K2)��H�1^b_t	}>��0=9C@����0dsi���:����[4��Z8�V��W����DRg]��=��Ε{=��n���s�tGg�t��^Ia=�`���k ҐjG�;�Mے[w:[ozc��W�T����+�e�LnIl��l���,�:�\n���$�ț�@�;)�z}�����x��� 5�����P�85!���31u���;�M�;W$�? ?|�U_�s�w��$�~>��D<��m8��[4��Z8�V���נ{?u����␟�����X�c����g�u`�!�[m�n�u	M�|-��?}��Q&I#"��8k��Z8�V���נr٠}�t�"�8�m'�l��l���"`{rK`{G��`��I��@��k��l�߿%οyh�Zy`ӭ��
@j!ZX�=�&�$��t����h���/��8���>�h����u����~���D!A @��H�c���9��g=!�e��P�N�A�oF���3��z�)z��{91����1�K���⣎�fVƞ���ӻZ���6K1�<�]l/<������5�u�����]��u�ls�]��dѳ\��u;۬�8֚��ql&�q��w/�]�������j�\n���4�7\f��)yb� ���N�kx��<��p����x�a�O�81L3;���� ���˹�����&���t�8lM���:11�'ױ��Y��1���I�̘<RH����<���qs��l����[ �]u1Z�Ib*�� ������{{� ݮ��=��9��-�"�$x�D�= �}�|�L`n�K`u�L`u�]�ˣ$�suUw��IDD���`��p�k�ID(�����Z��U�]T�Y5u�{�ـ}	'Z�� n�^�^��/�?z?o�ebl�P�TV�q�q��S���k���f.��ѿ~z_{�����K�іݖ��>��w&�z��.�����hRRH���o��03�P%	*�P�!*���u�o�� ����߿f$_�����r'NM�������׽1�zH�f�̈�HI+Ĳ�c���^���"`|�k�s�+���$q&�h\��O�����Հn�ŀ~��%Jn^H�lUa8�܏6�)�����nur�m���v��\Ί3��~�o�䉁�1�����zcoh�v�.�����I��1�����zc ��7߳�G;���@q��n	Ǡ6���u���$������%����bB� SRH̥X�jB��*N�v	B2B ~�"��!� 5������E��B XtNR�H�����1b0X�b��cXX(E�L�A1RB!Y��x���U�a J.!�) �"�ĉ��MG�A�4�.\e�U&g1� FA��"B2Hy����J����x+��UBE�1"��@�(H2�ZD	YB�3�s-��t@0N���C�H�@S�xuh*E4���B���(��CQOE^
�R"��n���&�W{^����	�#�&ےf����u�� =�׀~���y�0y�ӭ��
@jB)�s����g�?_?��}<h\�z�J��)���<�LTn}]s3g�|�x��N�����R�����N��`�Ӂ�'"q$��+��r�0�k��� n�^ ��U]`R�K/�Ōؠ��ޘ�7dL[�Y�BIU|t����QWwwVT�\��쉁�1���ے!�q�z�[4��z���g$� !B!�)��)HF�-�V��T?/;���+���I��$dQ7&��@���%�������y��>���u4��Y	�e��E�y�M;�\qkS,��ܙ�}��DN��n]v\Z-��F[o���|0:��0��:cչR$���M�7�����g䃽������s�S@�Ɲm1����G��&�t��P`u�L`t3�i���q���>W����;>�X(J�"U7�׀}?u*��
�ВYyy�,`n�^���"`z���$�" �Eb!b0V��;�^��""1��%!�˰����g�x��o[usC\�ܔ�ר\��P�i��Kj�p[�8���r6wH��Tƨl[������ݻ���E��uDH��k��&є:n��l�xՂsòR9����q�[��oi"�ۚ"�y)�{OV\i`WC�gtʷ4�恘���c.zv��[�]��<�����l�黥����'TC�<�y0�ܩy��L���vw�,M�H݇X
䓔�0�QgF1V�K�&��I?���?��nȘ��ؠ�$�������MU���� {��?�"!D���Հ{��4�v���Q��$��NF�t��(3�~�����`����������zܲ�W;^�{���J!D���`җuXMJ�3�!�׽1�n�L\�ة�UkM���"9�-i)�I��eع�>��Y�ּh��<=�{0u���G;F	
�� w}�`z�L`n�^�zh���p�8GNM�{^�z
����� /��D��矷ɠUo��s���׍ن<��F��Icv(0:��0��:c ��YTPI#�RW;^�s���{^��YM �;a�y#��s7WX�7xB�P�\�������נs�Q�$m&��Sq�ͤ����s[��5�L,�3tid������{\�+2��$��Θ�݊��vY�}�"�䑦��@�,����u�������(�QTm��U�`��M�7��= ����ߏ��
��H"����@�B���)#6~� �}��US��0-*0HV�0l���1����v����C0N�'&���u�}�">Q
!����:_}X����o����uђ�]93t��F�1]]�g[2-u����sHĠ^:}g�i�Y���nzuK//1%��P`u�L`��:= ��eQL'$������@?y��?K�X����	(���˛�H�7QǠ.����^�z9�M���@��T�,rE�j6��>O]`�k�g���@�Q"�1	b��럷{f���RG��F6��z�Z� ���B�}�x_�^�_k�?���yM�H��$M���&�/l�x\�5k�{�V��������ѳ�y�a�$�m�8���= ����{_�~ϐw��h]�6��c&��G���:cw:[�zc��UUWd�������ɠqz����Z|�D%2�_V {{� n��T�
��i,��X��;�{���U~������{�,�`�9$�$�4ϵ��J"{{���}Xݶ`��VP�ld2S;��nY�7\�5��y']��g��z�v�q��,�k��X��v],�q�]!�WuK�����7lq ��=ڮ;/1<j�9��<�`�c�C�:���tq��b�i���F����`�G���}�S�Mx���"�iAϔkT㎍Pp<��шH�nL�k�h�i���긋��6��:ة��5�:P��\�ҘL��&fip���D�������������5����%N��&5�y!#�*�NP,�R�֦��xZ�n����� �/]`u��(�Q�A�o���ڏ(�H��܍ɠ|�k��ŀl�]`�w�(Q'���q�⑍�7��}��us�����4/_=�;\��D6ڒf�׽1�M�0=s�0'tt���YyL`���H��٠fg��?_?�����:����]��#A��u�V�nܱ��wC)��IZCI��5�^mLm8�$��nM�{^�{۹�l�]}
/�ou���*��*WE���������w��J!�"�,��!-�P��)�9�X����u��,�)���85!�us��9]��(��O>�w�� mkWw6��2Ջ0��:cv(0:���]��)"`��Qɠ|�k�=�l�6}��>S;�׀~[���ʊZN]q�M]<����dS��u�[q��oI��9GOlxo��������{1NV�?���/�׽1�nȘ���*L@�2H������נ�@�^נw���.4�I��2B)�~m��^��B�	BB@%"�0i�O��t(��7��U��}lN�"�9�iɠ~���y�0�k��%�w{� �u�k�yRB6�@�,����נ�@�^נs�Ģj�A8���<;6&u:���,3<��=����qim�h?����z�j�`�9$�H|]���"`z�L`wtt�$������MTܗWX��y�B�S'��V��Ɓ��נuv��E�5dn(��?K�X��r��eξ� ����Lt��swEUYUu��
#�	B����t����n�-(K�(����
IDJK߽�Հy����h(�������ޘ�7dL\�ؠ�����⢆�λ	�{Q�0��g�fl^oL�t �\\˦�#x��q9;�բ��y��?K�X��%�Iz���������Er	�����|�"d���9�Հ���u�J��2�+I3,`{yA�׽1�{z��{^�[Բ���H�JCC��K�}X�}x�z��%>לh���!"H�6�#�@>�l�3�(�Ix���5�����X�(�Q+��**+�Ȋ����
���TTW�QQQ_�EE�EE�T ���� �UH� �  �E�� �P�"E �!"� ED�QQ_��QQ_�EE�QQZ
���AQQ_�EE��pTTW�QQ_�EE�������b��L���I���ͳ � ���fO� ��            @  Z�  �� �  �EP$)$�P��

$% R� �AER�   ��
P J�
 
 	0   e   @ @ ������N�:�N�3����� w)b�^LGݝ}�s�ץp��}�}���7v� u�c'=�}N�*��O�c����weo� }=�8]K������  ��(    �@w�>���˼]q�'��� �sϫnY]�}���XRe�l����}9ۊq:� 	�Ž��7��� 
gRe��;͝㻷���n���n �}���n���7�>n�������Ҽ ��( �T 
e����N]���yj{zy7��{�}� z����r�U�n�v^X���{]G�� ��_jry揽μ �>��}o�ܼ��� `� 1�� @0 4� 5� M�΀P 9�      �1 Ѣt 14FF��;���;� �� � X � �L (�
&� d   ��  D�(;�[k���Ź�ݾ��z_n�@      ��,�k��+Ϸ���| s�P(    Q���f��l�w]��x�]�w��^x ����ŝ��ɧ��GG� {��/���b;� {�ۖ����{�Ps����t��'�'����U|�P�{��]���üY��N���y�x ��̕)   E?�5R�(2 h��O��)�T�@ تT�I�Pa2 T�Д{T�* �"$5%)��� zj|	��o�����W?��������w�ý��*��9��PTW@TPT�pTW��"��������""�
���B���Ќ6�M�A�CMM���qԎ�jRF�XHjj.0֛ ��Xi�25�Q�E�M��iiB��Ò�q�4t!4�HD�X[�Mڒ�6�g�2��O��=E�`D��?��LC�cW���9�F@'�\��$!�������b���i�$�	kHa�4��@�����0�t��.��q!Sy�a�nf��	s�R�"��H��kB�h��d�������
�:�1��jB�����a�0���u{���:�E��@$@*b����Y�R6���t.���p��Ʈ2CB�9�$d.��1���$+Lt8�i/�T�
@��dB-1)R���k�)��g�+�I1�H�jq`�� �Đ�1%��9� �H@�Y�Q��$	@���^y�t ��)�!8z2�i�r�B+R��,#	/�RY ���t�8˳�3a�.	$!�%XVÜ��Á!�p���NM�%"D�Bĺ�d�p!p��\�� Rj˓bIa�J��H��KJdI�8��2�+P�	�͉6HcVnc.cR\�	fi���y0�s�aaHU"#HQ�c��DCрX� Ԓ�5禖�9���E�-�_��݌�З9�a��E�
:;��狤V����D�E$X�WP�"R�|�X��
�j|)�1+�7�x�&$4�WĔH�x�i�k�X�65ģ�Ƹ���X!4�E�x@�j�k�K��
6G�>B$ I������k�=�%��(	)�����<��a�FO!#0�%OO=¦����2�wr0�R�"��XO8o���%9��8���H�	|�ăY�s�e0ؕ�aR�f��0�� �!Xԅ0L|%�Ç�WS������tc��<X0!s$cLeF��ĸ���9��h�8_��g�Ȕ�x�X���j���oCL����j|ơ�(G�� |(|�i��Jxp��	����$� /:H���<�|�)q�����3�;��Ѐ��y�8��o7�_p�|�>��'� �
o=�H\�M瞐�`���ac4�H
��i���)������F��4�aL�N�)�%�]%1��"Y�E��7�\%Ny�.��x��&�J;�<%���B�)���	�
&I!��&xs��S�%��H\M8N���I������)`���N�E��OpMT�K��g��HuB)5�H\���ϼ"��Nxy�c
�F�.�`@)�����a ������|,�g2�8��Di���P��H�7\Ֆ���9�\Ճ9����Y���*c�	\4ƅp8I\5,XS\ R0�(K�)BH�Ta�3@߫I���#G��" ��D���Ǐ��!LM?����2S ��4�0����(��RIrIF!���,����bIŋ	B1#��C$��"K�e̚0�0�$���(B��#�-�JZʰ'��D��%�p�xaM�(�Xġ��	���(�4�j�1)P�@#��]OS�$$�B���
�AB�#b5��0�b!Z$+`[ Ky��y����h`Ƙ�sJ��p��ȰvS�s��&d�ʙ���9|�%�%�!4�����BP)�a��8����ˁ/g����|���S��j1�#������o<���_|�g���K�s4��3�.R\X\5�<8{��\<+��>�L��&�#%!u���(B`{���z@�y�0�/�7�+<�xK��3̳���#O|B�������]UԾ>D�&h�\Bs��NU �I�0#B5 R4Rx����S0�f�n�蚰���v��J,XLb@�)sXE�=Hz�ͧ'�}�=p1&�����y����&�}�2��D��P�=$�<`�0+��5~RS"T�0%���L!d0Ӊ��e����Ĝ�x�&��_7� x�1��eq�c�c��.{��y��fe�=�'У�I\^��^��o�s>e�I1:ƱZf�I4���ᱣ�F0����<%3^'���p<H��"���H�8�=�%�%�k	J�hB�s�����B.i��$����f�<���%qap���ˁ�8���w����1� 4@�pHǧp5�,�:��ޓ���q�HД	sxx0� c�|��y�¸��� �S|��Z��K�/��
o���_��>�H���Ҟ&'�=!pЄ�7)���ee�a��.3wn�p�\��0��taLB!!p�cIL!L��zgԅ)q WSR��5�T�r�H�N�ﾹB�,��xO	Ip�9�f���FH#й�B�Z�q!X�!X� g�����]t���N��i0�}T�ϟ>�r��u\�v��\�o��j��������*��)Y�K&��>q�47J���9�Nj����o�����_a���ۇ�~�q�	R	B]"B�$l0!�xj����¡�
�Ib0�d���$	�h��jd
`a�}�$H$�o6L�J��aJf�e3S�3)2�Od��.hpiw<5�"@�L)d1�CW����4�����$��i��f�
s\H����%1!L
�ad0�U�#dHWxHi�&��ff�$X2z���FF�(F���F���]#v\�6�9���q0(�|!�l.�BHM0��`�B���q�1�Ĕ�_<ӚzȞ���߬фX�_�%͜�sO>>:w��qu��x�)
����Rn��^2���":B�!��n�p�$��s%�r�\�RR%"BO���υ&�7Iq�)!�0��!a]�|V0�L�y��������}.i�sI�%eI\�XR���I�.K��e����[ޥ�n����T_)_���T�+��_Č�����\��Wwh��nKo���ٸ�n�}UH\��КJМ���%��H��0�0&F��\�=%ºH��$���©�M=R��z+�N!�BS���W^�.p*xI�!M8JF����1,�8Sx����B��$R�a�k�3nn����4#J��Bjh
��tcS�f�e�/LH��
h�@��Ja�!�<��7����r��\�y�>����f��a�~����^P�������c,0�.k��C)����M�� �r�C6$>�F����&��9 �j@��ﹼ���=��\	R0ee�!�X��߹}k�UN�WR�r_o3�><瞧��Z��{��s���K<����A7p��󤅥i
�K�+�8g�����a��RH
d�BR
A� �(星�F�:&Z᎜`��.��s�*�8x0��A�20��x��jD�<)\�(��8ˎ��oNo9�O���$��)�Hp3��<<�)��M�٘i�4ap�
��o5�^1�s�)�
2�q!^���t|B4Jze�����ԅ�93��p�N2愹�����׆���P�L����=B��Ӑ���i)��3q�	~�������H�:�d���.Jk�w6%0��$���'< B\�ad>%)�m%Rf�p�<&k7%�b!�āA��A4����o=JF<@�_�5���:�Fm���L%�N{�!�%2�|�a���Q$c7�{�=��C�sɶt@���Ќ<] �{��� �   6ضJ          h    p        �    �Y[m�H�N�lUQ��yn�b�@D�U�[F�5]� ����[����6��p�		V ����])�৕P&�h-$؛\pl���          m�[��N�]�mOTR���[@  � ��oR���n�l68�ƺ��D� $ m�t9�2�uTm�"&�
��+VtW.��UUw�����n+�����]D��k�&�1m8T�ԵU�ջT9T���Y��smӈm�"� �$I��6��D�@��8-����x�gZt�I��)��Y]�f�)� $6�.�۰������D.V��U��p�:��cW[6ǐ�V����L�,0��� I �N�T��u������\l�-��8��5l�$�����ngIt�Mwt��M��ޞq.��������#7m
�v�    ��I,��� m���P��a�Ld���   m�t��E��:�[%t0Һv���`    m�> m�  :D�A,�am$*�Z����君f얚䭴��h@ ���or�`ڶ��6��
�"�tUNq�t�+���mE�$�I�-���ʠm���I[Y�LmK<��	"�*�T�*�UuP&���m�U�%�p m��d������w�]6p86���l�'i-�.�Y����uc'd��]x���3�|�]�wP�@8�͹��6� #u��h������9�`��m*�݁���D��œM���g�Nl8�hI�@m�$ �d������I! ���XI��<�ҶL�UQ�uP.�h�X� [V� =,�e�^�6��"S�l�&�  n�Nċz�8x�����+h��q��j��%� � ��������D���!�YYpPu�����azm�sMn��@k�G[�j�`���*�:�'8l]Ͳ@��z�l9� p�Ol�ߦ}:I~��I֛ D���
��O �UWUZ��.˵P��ꭹV�v� $�m�g^ -�v�7m��� ��n�m�]r�MG6� 8$ ���tK�Wj��ge��n��g�ѪvV��iy,� �il   �:�`۳v�:Bړ���M��$s����m�m�	�m�� �n��X ���l���&հ�YL��Զ�8��Vӝ 8  rA����Y�\	 6ٯV^��m�Π-�۶6�`�l9l��p�5UT�Q�j�Zt�̶�8m������-�&�ۂ� m�����:���z�A�_Uz57]텥%����ձ�pTpmUT���T�-�t8 Tմ�[I�k��]�78m� -��wI�m�� ���[n�	6�k�e�m���;,�[R���*Vw�j��t�)��umGdzT�Kh�[���٪���mmAmN�^�+���m��T	� i�#�ka�q+WP'5S�sT��6��	A0]��eΙ$�� � 9�m �6̀�8� � ��J�G�ImmmZJؐm&[d�A�6�d�`�6��fa�8�`���N[:Pi#��   JNK��"t*�J   6�e�gAΐ-�)V5�[%[@	;E�𶺔���$�!$&�:m������0p�K�k9�z@�E����m�n[A�^��Z�\�-)-��. ��n���ݶ�Cy:��t�MfZ�l�n!#��H��� �I���c���� n� 2$IImi6^�89��x�۶�Ԛ�� �d5� q�������/�X�m��m�M��$�	 ��J� $��\�֭�[bi����e��bI�t��l���[x�[m[&�sb@@U�jW�dhH`*�\۸��  $pd�l�8 8h�[� �f� �kd�$��f�!����H��]ٷl6�kht����/Z���n��vI�!�8%]@� m��� �^�&��H 8�f�Llr�/Zmֱ���l ���m�`�ե��	۵Ѷ� 	 �ZR�W�N:�V���61@ܫPUA�p��\�TEb��+* �r��Hft� q�� ��U���5KU�ZYk`Kr�[J�s�-hӡm���I ��ۮUVq¡��\���9ƫr�$��gm���l -�Y��m�z�l����J��V�m&Ͷ����[h-��ݶl���NH�\m"�tB��]�onyS<�U\�UU�T�E�`%���R�vz�%�T�R�$  �;�zN�eU�T�9�ꬼJ�6����r�s�{vaӢwj�
����'xy�S�k��7i+"�m�eZ�����-�1�Z���#-��j� m��[vݤn���.,Y�ڀ�*��\���"��`)^�ȼ�,}�_Uҭ]J�@���!! 	�nu� �^�J�[	���)�P�����-��H  dK4��ۻv,H�n�P 	e �ku�vHm��M��	mUJ�mm*Ԯ2��$�X�l�M p�$�+Em�l�流 �nې�Xm�4Pl�!m��  � �  �I�  m� ����fו�lAk+j��a��l�[��qwE�  pym�i2@���� ���}��   ���:u�I���� �6ؐ[m�l�$qm � �[_rG Hw��`-���[vض�p ��[�\Z���%��/}�I6�:q$a�֖^��A��l��H�&웚׀ �m$�Z/m��t � �E�����kM�n�    	�+m���-�BtZ6�@$�m� �al�b��V�W�^�Ha�=�ņ�ܐ�౵�'T�lq�UYFǷBS�p*�n��#�4]%���aƸR�`6%���l7�q"�R��rA���t�8  m��m��pа��-�V�����j�a�<�!��ہ-�J�� A�mR�j���[h��[@6�&����Nm�[�ZR�  ۴�g��K�ؽm ��	-���`�O^��nm��T�a"Cm�u�[KjB�m��շnKd��6�D�M
ݥZ��UUҭ�%Q�Y��� .��o��n��[��[u�� �p*U��Wf�R��,��-�^� �`    ,��In��	 m�[�m��u�m�7] �  -��6�&���l�\
P  $[@m��d��ԭUu�m*Y`5ȴ�*���*���UWJH
�a�@�l ��UUR�ʰl@��(��������j���Xi�W+�s��j�����Qr��J���(!6ܘR��mI� �� >qh��T��86ͺ�#8 u�Z`�d��R�,W;]�,@��$H8���� �  $ �t��6��8 -�l6�q�  �[%�h��!m i�[Vշ��H�C���M��ԻsW)  ���+���[�`)�V܃�JܼҮ�U��:�Z��'X��.�:v� v��h;�7 ��dm�f�8j��*���&����-�K( %��I&n�3�u�H!i��pk��XkM�� �a� Ӕ���E�Kh�rۑ�&�Ͷ^`���.1U/<������*�!���5r�� 1Xz�F��Z��(�T�շ=GQAR�g�������S@[Tl;cJ��FT6�T�Y��� %�v	��[���� '�UUUK��5�+�-&Fڪ�h-�Amq��Ͳ�)\6��٭c�,0   �ä�LY��[$��q%�� 6��n��� [xsm���h� ��E-�ծ�F �����n!T�W�,�k ��-�HH �Ya���l6��[@ 6Z�[x�6��hr�J�Q����ey�Vݶ�-� ݤ݀ 	l�-�����[@ ZWl�jm&l	h�m�#�$��+\� �ԁ��m�-� m�� $-����2�:�^�l8�@�$6����a���/gV�p�{mv�� H�o��- 8;Z�f�ZI��/ie�L[X5�`e���$���4�ձ��Vݴ=uT���ҭ 89m    -[�� �� p�I��Gp�߾�n� -�������d���m�Hi� i�M��H�1`���$����:A�� j��� GM�a��۷+km	�MZ`H�#�h������2hiX��5��L�e�6�k�t6ʬ4�KIUVyLˍҫWUUT�α�@��ѱ9�Jf������Su� �N�   7wwM���E ��T?� �8���Q�0_�N @N����� /�_	���!���G���D= &��P�(P�D;����ʽ�T�@����� ��1A<S�<O��AS�z��{��Q>�t�= O�U"
u� ��@�
���   ��U��) �@#@��P@��
!�����	�EO�@�U�`�ȈqtA<� O�Q=C�
 @�@O�G@�"� ��� *"t@1S ��S����}�:��0�Db $F���q�E�+�AS�0�Q4Jz�> SՁ�P|�"��('@�G" �P���s�P�ނCN��'UtO�Z�\%�T��S� �*A>@�Q��W������4
"'�b�$,"		�OV0$�����tG���|t�z�!�ASU�#[QH^ :��:D~ES���Sx��QP����A��C�D(�� ����꣠�~E|:"Ꞁ-UtQ�� "�T?�Ex#��/�Pi 
{���  �h�  �-��X�;k#If���{Ur]5�F[@Ӌ�C�Zu��u��m��B�l��bV��v�nxKvZ����5v�]���k\��^��ηvW���9��Kd���\UC����EL6J�����v��E�!HT��� �'n�Oe�n��C&�i0�l;��9��z��G�F�j�BO(�8v����=�[��T�&m�u)����Ų�kN%Ȁ���s�\1�׃=����4Y�=9¶w`[�����iq�rƎg8n��4��WE�1�s[Ϩ6
TWi�(�'�pD������Z�tvx�8\�J�pT��x6q�jy����D�tڠs @��m���ݮ-��ЇWUV�v�6esP��Jݷfɥa�����+h�pms6����=fɢ�Q��iZ��hH��l$��q�ܲj�3����t�h%�`�s�8M��,�nv8TP;��A�m�e�������2�b�ܹ��cX��t�����٨{ C죖�[Qj�1�䛔��n�<�D���m�R r�9.��-ٶ�
�X���q�q��Z�j2]Td���<�KI��$B�}t�N�KoC(\T�/�z���x�bd��)�8t��8�rR'�q-gw���'��R�D���ڹ^V����f�\�Ct�\��v^]�<�/Z��be�FhsƛS�c9斷d��ͪ��;Yq-ҧ!�����l�v ��5���=�M�n�#�Xr^�5�t�������K�<ؕv�tl�7�Б'5kq@�:�5���n���#��u�p��ѬO�㍁/0n��]�X6w.v.6(��UI]v����p��a�Tn�Х�!3e���+�8�rF�][�%�	���`���m��K�O0]`�:�0lsQq{A�E�p�GK��/;-d�'�]:��c �H	CNmc��Ѡ�l<u0�R�g��ńs ���h3�ww(���	������EH#O���/��b����S�:=Q<ES�*��)�0��jY��b�#OXۘ����t��p�q* ��<�[�c�t�g�	����Kif�u�|V�y�Ml���{·��Ţ%1u	�� q�N�m�˷N�v|��t�y�Ul�%��1Nu���s�f�w*�cn9ԝ��Oi��C(�֪|���1gn:�0vl"mv�v`º6'Uså��"'+%�7Ks�g=�w}���=�����+���>ʯ���6��"��c�����6�Cx14��{Ϫ�=�� �����K�̭,f���L���U�Ӱ;��w��!&�=ݛ���������X��Ѩ�2d$N-�d�d� �- �Ih��*g�615��q��)�w>�@�v��mz��ړ����O$�w>�@�v��mz��h �-�<XĒ���k�`��5�D�x^#��gj��W8�ƞ�1��Ĳ~Pyqh�ՠx��@��M��Ze,2��$&M��w6�I��{��| )!� �`b�	�� ��s�e\�|�|���UUWQ�kc��o���uD�Q$�z��hϪ��w�z���z�V�R5&&!M㖀o�.I�I�@qԢx��F�i8��j�<Vנ{l�������5qL#��ӹLV-M�u= ;v�WklN$�h�IRv=/���ky�b�rcQ�d�H�Z���m��;�U�w;V��5�W�������d� �- �Ih\���Շa����~�<X���k�-�ڴH8�� ���1"A#N±@�u8 �9��;��岚#.V�Y�d���(��;��@�[^��s�p,2�i��F��@�[^��s��j�>��3;:�͸!����x�cKp�z3�����kf�"���p=[Ν��5�	p�k�C����I)�w�O���Zs�h+k�<G�թ�	�4��@7�Z�$�d� 8��-���72~i8�U������߳3#w���ߖ��g,Tof5&O�����$��� �-���{��A`US���B��U~W�� ����\��rI��;�qG1E��q���;�U�z�W�x��@�-�(������!�!�i�.�����N�J{q�l�b��L����Bʲ~q<X�������z��m~��0��i`c����mT:%S��`v㘀��1 �6��@IA+I�� 2)�z�����hϪ�=W����C���8$�zUnG�x@N���;q�@r䘀��V�#N��Rs����_��Oo�߳�O���rIT����G�{ߛ���u��ɸ�ܗ�����5��v���2N�m5�Û����Nۜ��e���1��\qZ��k��LZ�q����/We�ɶ�3�R�<sf�^j��ԧ^�^�.ÐT9:v��N!{b�K�<Q۩���z읲C�E.ݎfS�m�i�;�#q:\#<����'Ƹ�(�s��$;�%�U=F�gcwN9�����_��{��y��ܻ.��8��[]	�7gi��T��t엝�'q �h�EkKu���}�@r䘀}�x�:��\3ƦI2~M'�ⶽ��������U��y�2��G1E��q��`�o�n9�\��C�cY?B<xӆ�����z��mz{e4F\�b���A�QŠz�����1 �6��@z�����͌���; hܖf��	��z�a��Ql����q^V�t���r,�ūC?��o�� f� �9h�s��fn�nK3e�w9$���g"�|X���Nŉ1��''�)�@>��sV���������
֤i��1
C@�}V��^�ⶽ���������72~i8�U������;�U�{��ٍL�*�-�M���ɰ5%	,�ޟ�9���^�@�υrG�0�$k9�3��9kC�u���@VU���<j�,�(�t�b��6��;�)�w>�@�^�@�[^�� �9�Ǔ�i�Ĝ4��o�l��ٰ8�vl�+�X�ZyI�P�N���ǝɰ>y�6jQJ��E�ܺ���Nk�3dV)s5 ��N=�mz{e4��h����Ρ��bR=���s�U�����n9�����������g�����\캍a�0˷7-���CJX)��D�)��Z��z�����hvR�{ܠR�Ӱ8�7�"I��wf���i`w>�~�ؑ�*����jd�'��q��{؀}�x�;q�@v��Ԕ�Қjb����؈QQ9��K99��Oo~�rN���J� !H�����DB�'W��7^�� �9�Ǔ�i�Ĝ4��h/�燎z���^�M����x<�&���B��/u�;��9�Lp�Olzu���������ɍ�RbY?(<�8� ���h+k�/t�������\i�b�SR檬�fM�E%2nei`g'5��٠g:�"q�pB�h�� �9hvM@rd��vK���q�F�)��Z}�hWj����W�i�{�J�lM�s'擉 NɨL�����r�UU�yů��H1<I��	S (����r'�1����ڸG����G3
3��fպT�	r򽵫��U,W-�Twc�� �˙7���۷}�ҧ5cv��x�s�����n�{.���k�)��Z�d�/sx�U�g�77iӶϋ\tgN,@��&�ͫ����Kann��S��u=������s�O^6��k@mK0c�����6�f�����S�Q���>s��!�5ּ��%铦nFva��ƛ �c�r��w\�s�� �k���u]xح@?g��#{x�	�5�wK+�cSX�A7�{�4��h�٠y]�_����؂�]y?!�y.h�;��; �fU���o�;�����@�e�1Y�d���(���@�V�{�4��h�_��Ls8ӒhWj�>����������@������,�9?(�bB����-;�M��p%�b�.�M�l�x���{�ޒMc:��c��@�Қs��l���{���T|�W�n@��
C@�����^�@� (��}[�U�od�&Ih���P�Cbo`ې1����@�V��gﾫ��� ��Z��D3�^����e��92K@6���@�j��x�d�?�MŠwt���fffVk�{�V�9��؅��2��D��v�&�׋�#��q��[�.�khc4pc]vA�sM�`�y3x�� �߭ NɨL������XF�eF`�RmT:%S��`�ʽl���72|hϪ�-���ƛ� �Ɯ�By��o$������;V���qȑ)T�DZJ�l)��1��T>��	B U tdc ��*B��(�� ��n�E���B+!���ĄH��$$P�D��OVTXaC�q%u,0Ĺ�/�P Bh�
!	$��bE;�V(J|�ˁrI����߂53>�����q�G�O�挅�J�ł�H0"D�"E�=�D���Ia$%n-z�
d����T�W�/��
��z+
x�2��5�
a?b\���b���Q�p���� G�W�����=8xQ�(uDz��0 8!��(���sڴ�f�pr9�O��pB�h���r�욁�U��}���ʰ�\���$lB��;�U��A���`sgu��k���F-�|��ML��x�m��;�&�f�p�7������Px�I�Ů�%��7 Ӑ1$�����4+�hޔ�?x��~ZZ,>i�ȦI2~DnM��[���Y�Z��@;�kc�$�$�T���zS�M2D�GSNÉD<�ߋ�Q2�_��ڳa%�gu��b7jJ�I:��"������w��D&�;�VСDsku��B?���B��F��V)<Q|�WA@����9���Ϭ?��#�M���T�i�$�'�ݯ�Ģ�֚�B_0��ia�Q�=�@c޿�4������ �^ǲ�3j�'<�p��2���ݾ�1��p�kvϫ���y����;��;�K����fNk�[3��`*+��$d�Z��4��h{l�<�ՠr9aι���e�� �- >ɨu_}��fl�c��<�CCo`ә?$�ZoY�y]�@��4��h�
�ّL�d��94+�h������ ����x�:�@!{y{�ٙ��\�L���-\��	���z9������"^t�έ!'5�2B$�.�
1��z����l=��[����/�����S,q�{L��R���̗�V2#�$=t=7�=����c��chD�d��v^����Cv��a�ms�΄Iv�3� r���X��V0��l��'s1ˡ��N�t;��vg�	5���Ƈ�uFa�κI�@�~�n[�Mnm�I�7	qkLn7N��N��qpu�/Cў��ʾ'���h0�'C1~b�*�t��;�U��+�B_3ϻW���a�ݥ5*�s)�sEꈆ���v��[
��6w]��B{�zXźH��mT:%S��{�a��V6w^�K��ZX}
ef�u�j���J��UUz�͝�`n���;�U�?f%oY�#����D�m�;3�����fVk�w6�+�h=�ZsG#���x�d󎐘7R�]�l�g�on�7�=Y�v���c��Rs��Y�y]�@�Қ���M����sI8��Y���P�|ݟ~��^I?{��4��oٚ��*��M��&Oȉɠwg���k6BI���v��V霐W��_���@��4��h�f��v��0X[1Ǔ1��^h�o�#����-#� ?F���~:yp�]�L��x
�C���Gki`Yd�CY��,�&�r�q\x��G�[�hWj�-�M��Z����q8ԒhWj�-�M��ZoY��w7#dD�S�3;XX�����b�������,�}�y$���o$�YՇ:�RBc��Rs��l�<�ՠ^�M��U�bm�4��SN�3��`lB\��������q��(1���T��R�M�(�/	OXP�&�� ԁN����nX�:��E�]$���x�?�Z��;�U��f�zg$�j��/�QŠ^�M��Z}�hWj�-�*tQ��m�ӆ���� ��4+�h�S@�e�1Y�d���(���@��-� �UUUuUV���@I@��n ��rM��Z��;�U��f��wd�A% ���!���glv�C�����M��S�0�w:wC<�tf�k�Ǎ���%"�/t����� ��^��sgu��h�٪uTR����r׾�?{P�{ր��u�bm�4�ŉ'�_m��ڴ�)�w>�@���*6�Y2I���P�%�{x�I5 t��T�1~b�-��4��h̬,�s�D(�!BB����39Sɇ��J��ƽvu��]I�x(q<]Ʈ��ct�uNC]g�$]˹R��Mn�'�pSlT
c6{���N6�4�t�Ż6�K���nv�lۮ:`1���l�sݻuփ����S?{/�Sv�z�����iiج��*y:nLHf��玕Z�/5��e�2�[l�:�ֆ:�J�E��n�� ��
�aSr�Q�2~����w]�s.�nkN�9;mFC2�q�rK��iOn3͓�:E��)�� Y��&co�(z���e,�s�(_0�����-�H��j�ƈ��@��M��Z��;�U�[�K��F� ����v��JhϪ�/�S@8�wpqF�D��C����Z��@��M��Z"�9�⑓lB��;�U�_l���v��Jh�&W1c��8��u�^m83n��lݝ��y4R7A����h�7�4� `؛sNbē�@��M��Z��;�U�{��z52HkK���O;��爾 ��USU L���%�UtA�`$�#�	�5B��Et(��
y.��rI��{y$�S@=3�
���1G�I^���o2rӶ�B����v����{;�6�J܀��EL��8y�IZ��ԛ}��|�o'2��{9���|�z�:)�mT:�S����s���6ީ�ݏĒW�x�V���$��:��@8A�g��U�3�Η��z ���L���p���ܮ���^l�"j߯���~O�Iu�$���-I%�ݧ�$��dwdqƞ�=I%��}�������$����IWlz�K��u��dSS#Q�ͷ�9i�m��/�)P�!~�$M����{i�%��or$�,I9�RIw�i�$��=I%��$���-I%�g,U��"�$��F�<�$�vǩ$����Ē��ũ$�۷~�@�~���}mu=��㛇l�4���.�l6U���<j�X�P)���\�t�(�z�K��O<I+]�Z�K��O<I%]��I/{ ,��Qd�m���J�w����O<I%]��I+�y�ITc�1Y�d��DQ�Z�J�m<�$�vǩ$����%k��RIyp/���qdi�D�<�$�vǩ$����ĭ�s�/-��"$��1*u<?f~���o���K(#�dqƞ�Km���������ߙ�m�̽>��̜�5$��q�o)���P�0l71�d�jٮ2�Np� ÷V[�a�uk`�3SBd��I�$���5$���y�Iڦ����W�$��Plm�ȓ��$�5$���y�Iڦ��}��<I+]�Z�K���"�$��F�<�$�vǩ$����%k��RI^�$��9 ��܌�?�Q��%�v���Ē����ԒW�i�$��=I%�C�<����eI5O�o2rӶ�{��i�7m���nr�o}���$��b����0'C�#X܉Hb��"\��"#)�H0��
&0�1$#@�
B���@���D�H�!B!CHE�$)�0���F0Y���)��!HLm"C*'�c	�B\dbK��=�D��OY}�fi�wwmwMt���O�&� x�a>y�7@�W�0�T��|�¡���t��B,B0aR*5J��搻�HD�c����_��HHI%O�R�`BB����z� ���D�H1���b�8Y��AW����R��aV �	X 4!��p�|�21 T|����#�����!	���=�}�x�H�BHH�@�4�n�{�����+��_� G �]W����]fu�c���)�R���UU�[lcG:�K�y/���"��R���D�@(���/U.Q��J.[O^�#Yq]��)� :1���3ZXZ�x�E+qZ�&�^i��S[��Z,d��,�gNN�f�v� K�ˀ��]9�͹�J����kl��g���*� \�e	�4���{uS���ƥ8�%ݕ�b��E۩�|�vѝ�^3�����<�Ϩ���'9�V�|vtv�5GGn�8̶���[�8�V�ۜ���k���r`Y�kn�#�6�'����{ݙ�<iݪ-��1�l<� '
1L�J�0H9�����i��K��t�7D	zzv�VM��HҭEl���nغ�`h��v{fKV�.��n.�gK5��W�x�ˍp�"��Ku�R���r-�k[�i��ܑ5\&3@�p/#d�rXՂ$�ʧd�Β��;�3���a�OD����&#c(�eGt<ݧ#cr2K����4���2��f���v \�V�u��^��vσ�K�����CXM�Ĵ�q�on�q�؎v8G��u�YP皍Ŋ�q�f�M���l��]Um�>1��Y��S�(2�V�[��7���Tcpp��8�ūCiPN0KV�m����챱�tu`��.�nz�b��<8�I�r�lO;�-���lj�m�g)&չ69]�Bkm; Yٰv-�ݳ�wM*�CjZ����qؕ�
\��A�*�* gY����Ӥ-�x��s�5���*��K�#�+���U:5lջC�*Ah�u�{tN�:�q��fv�V��c�̚3��x�S=m�we�[� �kUm��t�#l>#m3%�xc��MPC�m#�X����3'e��ݢ�>��Y*s�������ž��s��J��ضؑS������3��ʠ5�6By�a{m���z��w�Y��mӂݻ��sT]F��l˔k3wf�v�˖d�.��U@(�
�_T�.��S��D�8��x���� �O9�ۻ��牖]zvY�eh��%q�{l	pӋ�H��ך�����j�Nͫ=����Ճ&۞z�:�cNֲ^H���雱�9'��P��3�3��ظ��f���.�9���$Y$�N�����z�)�#�qIĈh�[�N#�xis{J=i��;mX�ۻC}��]u��1����0p�I�˵��]f�&{L[ewm�
�c�z����^�z/�RS��38��jˎ�/u�X�3�l�����IJ��4p�E�V�%9C�]	�f%��G2�~�z٠_]Ǫ�77mX�d˚K�UL��̫�Q�	)���y��zՁ�������b���[���(*��l�;�j�zgwkŀ{}���vrj�d&H�E�������[gƀ^�hWj�<��X66�ȓ��$�hݰ@ɨL��ȩ�p6V�n�K����]�;6��3�k���[2�s��;�7p�8�x�բ�4ޑL�d��N }~�P�%�#�W�����a$��]fI-T���MU��Nc�J%B�>EC�G_�y;�w�$�����$�s*�(����k\�t�$�b]S�7>�s@��M9"�f��v�ѕc�Y?8�B9�{Қ��z��Z
!<�o��� ����L�eS�����1ɎZ��Hװ@q���,��J�6�R��/apt�+q�a����:�e���U�^�d�p��������\T�}{}U_WҾ���;���ʰ��$r�$�@�z�h�`���1ɎZ��U}v{Մ�3��)���niXܭ,�w&Χ
i$��k�;�`s����2\�S�UJ��3E���|��v6s]��w-X|��߈�E�|�Y���nE�yύ}_UJv�+�?M����-޻���v|7]�ɶ5�	�Z�nr�6pRܩ&���S����7 ���v>ݎ��#�|~�G<� ��Lr�_rþ��@Ha�H���)*T�SJ��{X^����v6w]��w-^�9�66�LМ�uNj��9���'1��P�%9Y��l��=�Dw�$��)�߱>mn�;�j��{XX\BI@��P�/BAW
�I.J���yu�����HF�$�@�z�h~�ϭߏ ��~Z�ڴ3��8�<�9Ytv�t�������r�k�޷';��4k3�Z�k��fby��{���$�x�ύ̞�>��{	.D%���V�L͒�UR�u.h�>yܛ�BP��L�������Z�;���!����l̵j�TLT����;���;��Ԓo3+K�sf��dC��ɖ�$��Ꝇ�I�s~VfV��;�a�D'ͭ�`fcR=�5JJ�4TҰ;���BK�	,�z�w��;��Z�9�C�w��,�&Y��!7:fgP��u��V3�fn��n����5U��ZsHdK�n޳Z�9+OP.�&�7k�����8CWX�'�b�.�J��ё��au�Jh�j�݊��;��f�/U����v�6�3n.aݲ��Vqѹ�/=���iP��������qv���0]p���k[��{-���iɏI���lI1��b�ݒ�|�p�I	��rM��kp��U�{	�[E��<p�ў{Wn?�7=��b8l(��mEXɚ�,���0��6�9���;��HIyB\����`f��?�O��cIǠy]��~H�~��-��@�^��?bAB�����HF���@G<� ��#�����w�,@w�n3������$�h|������{�%�\T��D31�UR�u.h�>yܛй���;�j���Mלخ9��H��<���V0�������ruʯNx���M&;�-l�Վ�"d���r=��Z{�s@��O���ۛ�"�V̵Q$�7T��j�"2c�5ٻu�`u�l�d�;�-V1}�c#��h��|�6y�l�;�j���2+&hL����ˎb�$�느~���n�hB�5�4䌑Li8�+� =U�+�I7���k�f^m]Z�竀Ӟg�t�������l���a�펮%fݚ�_���>�a�F�ARO��m���a`|�:��9����&4L˙z����niX�k�M�{�66w]��w-^�l�ѣI��.�U*�R��9���'1�P��Е%��lG)�H&�@s��!���ҴϷ3*����;�6w6Ձ�����(^Q=��"�+�-TI3����Z�>��mߏ ��~Z�����*��4Ɗ���H��5v�]�v�e`YN�M���B�����1H��8G3@��K��>y�:�_0��ڰ9�6+T�4**B�f��>��;؈��=ݛ;�j��{X_�	%2f����5S%S�-�M���zl�j̈́�I�̭,/��@89�9�BDH�?�fg�N�������`|�6B�
�����
�Dl(��r�~���։���U4�,I9�wJh+��+k�;޻��q�O�&ML1Iq��KW��x�l�����،�]xwk����wv�����Ʀ92c#n�����x��@�z��	$�a����άi�!6ʡQ1R�w�&/U}_}vG<�$�\roT$�g^!��=�j���T���V{���%	%�L��}6_��;ќ���,��x����1[w�@�}=�\��*@q�O�V�u��n�n�\s�{���o`�* MT-((AH�]������K5��[�;��]����C-�GwX��_�흾�]��K�Mu��]qjCc�#D���H9�#���\�,ܢ�e�'c6�vI��$��{sN���;3��YV�t�7��n��.�8wU�q����%��^��l���Z$$0rj�'��73���_,t��0덧v.7M=�ׁ7N:Lv�%�M١;=q�6�"'V陹e�77s%�Y�S�'Ny��[1Yu�֌.͸^��t�k����Ł֧ɇ�����G6����V������.p���{؀}qR���rþ��@"+��$$��"���]���E�|h���@�[^�n>Km�\�9���@6�Lr��߽�@G<� �K
7���Ɍ��h}��K��=[�6yܵa��<̽,u`Ѥ��N�A����ⶽ�/_�� �ύ����3�}�/Oщ�ㄐ�ȧ=��2�Τ�}��Ƙ�}�<�8�!8	�k��@��.��7>/w8sʐ�����\A��i�c�4�d��s4��qpQ	�E�[
���5��vl�j�Cg1�j��5EHUL�6s]���ɳм�w7֬{޵`s��F���"����*���빠[�j�b6�]�t:͝�n]T�L�:��;��V���/���k�1�d���v���p��E�raWDh0��j�+v#RO,-����ۦ���wu�=�
���M6��n�ڰ>��;fO�����Ձ��h�3u#�U*TMUR�>��Z\��*@I"�������Sn�5D�L�S�5����e�%R]�H,HE��0�H�X�0~0F�*�),²����!J�>Z�HL%����0���6�@�@�# ��$X���a /�&1	%P8�	����FD+h"i��������yH�JE��#��U�M 9I�Ң�dP�b1$H��4 ��3��s�1D����CRCA�8��*<D5Uu+J*h
@��<<@b�h���&� ��z*� ���C
����*+�@~A>Q^	�J6G/��Z�7�����NSɖ�(���M���O;��7wmXyܛ�k�;�|1X�d���h۪�؈������n��;��Vd�&fM�Y�;;[u��닏6��Ԅ,�k���<�Ɍ�3���=��w]o���S;��,���͛2s��fZ�/B��䇽����w��#_�9#D�cIǠZ�Z슐H�ێb�}_U]�g��#��J�M�����Vfe�<�P��!L���lz}�`f)]m�̹X����s4�6'���:�6l��vB�IZ����>�mL�H�J�UT�<�M���n����ڰ33-Y'�~�k8ܒ8t9�gT���j��u�c.+�6U���<j�X����wϐ�?gԹ���ݝ�`w�����Z��:�6lWa^'���OЏ�R-��s@����z��jߒ-1ы鉼��jhsJ��ݵ`q�rl��g5���VWL��榙3M���a�	'��ٰ=잴느8���˔f��$SN=��h�]�޻����䒀�P@"ŀ�]M�{q~�nvP�{�/
�,����G/;�OG+!�2�Ќ�C�.tC�]Oi{N�]������/8Rr�.˜%�ڒz�z�`8�|<�� �\�n:�C�u�©p��,m��cyx.^L�a���*��EO����\��������jK��F.q���1�vs�Qk�Z7+�2��Z�Lk�۲.�n�	m��e�rf�[����Aq͎[n��5͛� 0��p��
[f�bўǧ�b�3�Z�.�k��2J��ų�K�G6SC�45�bd��D������s@����^�k�q���i��'��wy����H\sc��}�V��~�a���(�2~�G3@����c��}�RG ;ߝ�3[��Zgۗ�����느8�ˎf���*�Ɍ��ӏ@�z�h}����W��Uz��m�RLA�)E�՗�������ǉ������z����{�3�Ќ�b�y1��s<�ۚ�9�	q�@>�� ��c���������$�^���C�<*�Q� 1�� Q�BS�k�`n�mX�������#h�Li8�
��@�z�h۹�x�W���S$d�$��B�w �)��8����mz��ͷ��sNf��Қ.9�\�n*@r�6�nf���'��sW`�ͻVX�`���K2�s�HwNo�fI<_fa��ocD�?H7 �[� 9rL@q���}�	&�@?�,�fe�ͭ3����@r䘀�qR��@|�ܛ�	�1KZԩٖ�IDĹ��9����'�}�����j "�8��E�B �)���P�z�Þe���9!U��@�1��f&�ci����;�A�nb�$�����R}�V{*�L:��#�,�{�`lDrwv~����w�)�\���ɋ�ci�iH�܏Ts�#�fYS�����q���'M�d�K�y&��8��i8���;����G�G$:�}6��\��䪒��m����K�_U��ܞ�.9�G��X�w �Ƅә�wt����rl�J��ٰ9����[Bɛ�2�TUK�,6"!�s6l=͛��-\��"!E��h��=��E�i�{�DkB2�i��\s���'�\9��� \Q��\�땻�����Æ���#\���j	��t�܃s���������s�ϲ�s�vO*@>�����.9��Vbo&!�#s4��7��f/$�)��w�`u�}6��Z�Q��#����������4U�=�z��빠w�)�{@�48��G1��l5(����ٰ9���󵅆�IB^�~zB��ɉ�2EIǠy�U ?UTqx��=�\sU4}�����UWny#��m�h�ј��{Cj\��q����"�SZI���u-�n�s�U�O)&%�݃��u��Y�tS+�=�>-��ȑ���Z�[AA���t�x��a�f A�S�Z½&�y�)�V�n�.'��v�zuu��pV�l��N�fĳi�V/��Oi	$l�b%Q�M���n���`$�tdZD�ص]n�,�mDc�����v���?�<<�9nm7:��5m�ato\v��nJ�b�q&we(=g�3�Z�k��w{����8��?u���7x~���nb����;�0���i�J�34X>�&�P�򈄒�:������`w��/T(J9���YD�ӑ����@��h�Jh.��{ʱ����ӎ�bJ37�`gr��>}�M���(���׷�`n�vZ~��U'.X:�Vx�_\�.9�u�H�O
<J�;O�H���nk��y�:���/1`GF��j�o��{o��x�v{���w��W?4��*P��c�~M�����w�k��"#��^4��?�C�<$sN=�z�����)����(K�3y��;������7���� �UO���"�$��=����� 9m�@r㘀vt���e�T9�,r敆���zXy�6�;�a�|�ߕ����I���AT�*��[s�� 8�T�}{�Wg��D��s���]�N�vӬʚ�=�Y�}9�������Ge罾�q�ܟ��Gw8o�� 8�T�m��� :�(ت�A�jG�y�w7�H�ύ�o�@�[^��"�k�4�c#	��rI��NI<�}����,����b�"� D �`{�D'r�nl�vՁ�ȜS�N���e�����+5�{�6��Z��Q�2�4�����9�'��^�����p��@rۘ��u��ͫ���W���-�N�gA�Nc��z9[��[��/��9�hҘ��q12FH�I8�;��������@�@�z,U��riK��`w��/ɳ�3f���k�<^K
=��"L�ۆ����-���� 9�U���yD�ӑ�/~��{oۚ{ҚH)��(C� |'� UD_7y��I<��N��{v�͸�ͼ��H�_}����v�� 91�@~~��㧇�j����Bz��ض�6}dX&Z�mt�g���>w
qB=s�mfm ^��nb�������;"��)#iHh.���#ߝ�h��Vy���	D(l�d%�J#�i8�~w�y�w4�J���ߞ�pr��ƙ$Q!8�?�3?/mߕ��������6|��v3�Od����4&����M��^��}W$�}�xrI��A�$`E`��(,`E �FH�H$3�1F C�H@$$I!#|��  �����ꁢT(��_~���ԃ��7���S�L�O}��"�p����1BC��`������a=A:8P-��iBU��;�'�_6�0"�� ���*?
����<x�[�1 �}dS�	Qv*I�>���	�<[��H��0�����x��q1!b�X�X�
#�={�6�� i6�	oP N���6MVu����(�`#�)�"R��h� �tk�#��}�N"��"�H�Vd6��q=t܋��OV�v�޶��=\�l[gi�k�[T��Z2���<Iv�@)�����K* �X(6A�V��v-���-��]���5���ċ"�j`O#��E	�%�A-�@��!9��E� 4v��'2.��"a6,�s�n3���sC�<s�qr`�뚇+4��� �B���6W�p�����=�N�\�R9B:mʐ'^h�6��Kf[�R�O.�F;kgm�MX���9웭	�;I��4P����*�dv���nz��Z�D�Q��Z-Y{`�@��,D-���gNW�[��
8����*ݸ8œ��q��[g�n�h���ۊF�
)��km�+BE�jz�t�C+A�l&+0��c:��f�M����2Wd��牔��v��<�@�r���u�yN�շ �c&4s68xg��;�Ӝ��=�7J�;��nϨ�j�.қ*ۣ�gw:8J����6�����GFn�6��[&Û���m�Εv��N��`�Y糂�UU��]���c��yڤtf�8-�����Ԫ�Z�t�i���Ӈ����@������9�gk�T݌v�;�xЛJl-�=(��S؋(��sO�zh�׷CI6Ɖ'��eD^�ʤ��p�z<!oT.�Z�[��wY<��U��n3�8��8��Cul�lϭ%�<���O3�m�qmB�� ck�ݪ 8�ە�nJ&U�c�t3��y.���Ѷ��M�%�.�݉�4����$�Y��68��ݪw�0�
��BS�w\��@p<q��i�ى�#��[J��9�i92Ύ:��Dqg�F�3%��������9�Er�猠���V۰Ygv�l�r���vJ��FF�m��ٵ��^^��rb��q��H�V��zNb����˛@m2�aiʝYj����߾�y�{�?�(A� }�"�D=O�G�^���"S�����{���c��/�5fB&���*ƸkYr���k&�%:$���K��vL�']�3[KF��n�����3��[�i���8�ǒ����Z����N��\�Й����]�1�<��n@wh�Z�Ny�h��7N�cga�Ѽp�v��hD�2�L����b#��X+��jݪ�ٰ��M[ꭳ��M���v��i��0�<��;��}�z۾�a���)��(���*r�1��΍��[��L3��85ٷ2���� ��~�1����Ѡq���d���{��!B��gr��=�X}��DA��9��}V����� 9m�_���UUVa=Yt~3?iEf�|fm���R����hW�h�>k���Mnf�ߡ(O;���Ǚ�`}��v�Q���/�;��E����!�x���<W��<{Қ���GDGd��\����p@랞�qB��϶y��F��hNm�����d�nk�4��G �q�����<n*@>����� �ۼ��en�v�ss�O>��9��������MB^�P��޺��1�zl�w&��8,U�	$JLHM9�{Қ���>P�o�wf��fڰ;��0���%*�U��f�<r��& 8�T��UrK���cZz�ة����sU6�3&��3=��3�-��@�wW�\���d�Y�+�rN펣!J�v4�����Gq��L�%���O�R=�빠w��,�{��J^K�~����S��D�ɉ�F�h�)�x���<Y�6��Z��ّ��N�5R��T�uE�Ǚ�`|�2l�|��� H��R��"N<!�*'�{�s@�ޔ�/`tCJI�r,�A꯿}�~���~T�m��� \�Lo$d�$��@��he�~<�o�@�[^��;+��<qE�a�
�M*�������K:�]�>n�a�'pȠ!b�(I"RbBi��;�S@�U�x���{oۚ���z�o$6�����ǎZ�$������	���i�sb�R�b�f��{�6��Z�T%�3��������ꖌW���ԏ@��h�)�yϪ�*�U|�F�ZBBDOEO�������ߌ�R�SO&'A��wt���>�@�[]��{��DD%���3S(R�T��I�Vݭ,/\\y�Vԫ����G�u���:͢:2��$�9�~pz8�<�i)@���@�[^��u��;�S@��б&����'����1~��ﾻ;'� $��ǎ^�pr9���FH�IH�;���Қ%�w�z���r=*�y$"�Nf��Қ����mz/m���/�%���y2L�ۆ��>�@��1��o`����U�?���}�H$���ffg�ݰ�&;�,�3�m�\a�"��t�iMtPV��ޮ���9��%yMb��x���_��Ӏ���1 '�Y��VyȈ���*���<�ŭܱx-�<F9��v7��v�=�xo[��<$���Nf��q�Y�s�.'s�yl�Ć�*�;5�pVy�gFq���WiU{tu%��ƵR%�#e�ۊ;�]̈́v����h��������Ƿ>���Cָכ��������J�+i^�s΍�V�X�g)����z5�}+G�~�M��{��󵇗��vw���R��dr���s�;��-_�$��;���Ǚ�`}��w�"�%2f��l�KO&'A��}~�Ɓ��O?~J������VW$}%�p9m�*�a(Ks�=h7 '^��mܷUH��R�����;aDB�f����@�wW�{�r��$���m�ج3�X�Zب��\SK�vy�:I��=+��M8��H� ���<{Қ��'�(Iy(Q��|�V4zW�UU�c�4���(��������d���{��ބ�!L��m�n�eR�[Znfh�~�~�&9h7 ^�����<N�)������v�$�6�ր�T�}{9h�ˢ���ji�4��ܵ`lD(P��z|1ߖ��}V�媴�L�i���R���v���vŬuCq�׮����N��@�҆j1��0����|hs�+�~JP�a�͵`b�ʗ�5*���w{���&9h7 ^��м�Q	L��6�Sr�U"�iH杁����y$�߻ÓO���ED*-F�PH�!�Nf���9$�Z���[�"�	š��331>w7�`gr��>����6�]�b�F��EU�c�4�󵅁�
,�/ ��~Z��s@�:ĮH�`R�Ům[�e��5*x�ф�+�p��՜��2'�$Kn(�ɒd�F�49�Z�=�`}�孄����V�25���AJ�35N��'������͵`gr��>���Q�J"d�R��d�~�S���h�~T�}{9hLr���H�y$��TԅLҰ؈Q;���̜�`}��vB�	4�D*�Ԕ5D�|���s��$��_ۗ����nm��Q`}��;�Dsk5�36Ձ�vS@��J�&/�6�di8�H�F�T0��am��k��z�F{l�뙶y7[f�6��f��h��@s�*@>���ﾬ��yߖ�P�����"�Iɠs�*@>����- r9���UUU��J!L��h��T��*���TҰ76� 9�r�#���\T�pwWW)nf��**fh��	C�k5�76��ܵa脔<�^�25���AJ�35N�>��X�!B�P�%��qpͯNI<�>��� z�Eb5!R��o�����Ujok q��:�i�ˣ���%���N��^�T�*tk�F�[S�c/Vc��@��=�7t���٨t��,�F�SE��98��-&�;;��]��R���Xap枬�j����yu�(��땶�wR�=����]�u��,w`m�v.��A��5:q����C.Ks�y��e*6��7���7e6i�au����n<�$�k[]��Z�偶���⍭v�,���r����ʯ^y��5�������`w��,�=��(K�76���1|�LR8�G3@�zS�ffbG��]��������W����[R�f�V�w�yw{��'���u�Hޔ�:�б&��nc�@����θ� ��=U_W�}{=h�g͉�2E���w4��4=}V���M��*N,�L��	��9z�{Muյa��sg�NF��qf{n�6x�w{���|a�6I"Q���g�^��@���h^����~��/�X�}�[D�2d#���'��ݼ�P4P 1�DE��-C�\�U<�y���rI������;X_�$�6gu��W5�*&*fj���������VzI��V�;9�����(�ڿ�8��8h{�s@�zR����vJP��D����5N�d�H��U5 �iX�kСs��������;�����^�SK*��u3S��M�<zr�M
��9s�����ۭ�X=���{�c��Z�y'�8�JC��?��h^��<������|h}�a�I�����4�����K�	L����skŁ�U�r���[9"��@�޻�$�߷���x@@c �B$D#�(�`9�H'ϢH� 	 ��+���<�z��U��(�|�"�"��=8�Eb��A�1 ā!�4\|��[�����d�LS�I>$�#Ib��=�`E�D�! H�A�g�wρ,<r�0�Or��8DH�2{�>M���x4H!AH�$	
�(�{ǀ�!�|<�����BBz�OE<P�'��U� <D�Q �_�Q��U���3��I/t��vz��,�D�s����_}�����?3߭��u�H���72�UJ��\�`}��;�K����w7֬󵅁̕�R�:
&�9�8v+���Wk�e:\�m�jK]��-��v=`T�[�����&�l_������ 9� ^��W,:�z�V]332��V�]�u�Hװ@s��<�)�~���i1|�4	����9hG�@s�*@:�=˙���52۪,6|�f������;��'����`/�#�<t*��;�v�uQ��.jS��$sMɎZ�qR���9h}�W�������n�K�V�米�6;j�+S�c�q�vZ���\f디��{ޭ�����6���y����Hװ@s��91Š��,�D�s���M�����k�9����ܵ~��I�ucM=Ss,�T�*��;9���'����{������LYQ��L�����?�/������Kı>����,K��߹���%�`	2'���p���L��]�ML�΂�%L9��O"X�%����19ı,?�=��~�ObX�%��w?Z��bX�'�߻x�D�,K��*i���۝�?���(�/#v�/%�V����;n�1���q�rU��a5���ð�T�3�d�ꒈÛ-� fṂ�i�Cln�v��x����^��1�gW/.��\������ݨt����;"��k/��D�p�ڷW�����g����Ƨ/\m�j��������[9�n�H#�8��'c�1��<izvۜbI�Ab�gn�?���w\��O	�Vul�㐞��3�;�8ۭ���e�sA�b���q���G2>ۛ�&��{�ı,O�w�Ӊ�Kı=�s��"X�%��w��'�,K����9ı,O��s/s7�\��n��yı,O~��Ȗ%�by�����Kı=���ND�,K�~�g���L*!2�G��\ԧSTH�ND�,K����x�D�,K߯xT�K�Dȝ���8�D�,K��~�9ı,K�����d�n�w6�soȖ%����o�
��bX�'~�?N'�,K����ڜ�bX�'�߻x�D�,K�}I{7wwm��-�niS�,K��߹���%�bX~?w����%�bX�����O"X�%��׼*r%�bX�{�\Ζ�8gQ�E��qgG,�nҎ�X�h�+u7!��'=vṁ\�qs)���H��w�{��%��۝�9ı,O;�v�<�bX����Y�L�bX����8�D�,K�����.�l�s3v��Kı<������ 0W�����L�`�����bX�'������%�bX�ws��"X�%����;s33�d�nf�'�,K����Ȗ%�b}����y����;�s��Ȗ%�b{�{��<�bX��}���&�nYr暜�bY�"w���q<�bX�'n~�9ı,O;�;8�D�,�P���xjr%�bX�?���.�˛�mݜO"X�%��w;jr%�bX(���|�8�ı,K��p��Kı>�o��	��	������eU9eD�E�{d���$K�S�}J�� <^눍h�HͰ����f\�.���smND�,K����'�,K����Ȗ%�b}����*�&D�,N���jr%�bX��b�ّ��N�i�f���	��	����Ȗ%�b}����yı,O���S�,K��s���O� eL�b^���������ۚjr%�bX����8�D�,K��v��K_bS� L9�=���yı,����bX�'z}J^��e�n���͜O"X�~BD��g�S�,K������yı,����bXʋ2'~Ȗ%�`�vS��݅�M��fnڜ�bX�'�߻x�D�,K����"X�%���s���Kı>��mND�,K�����R�n��3���J˅�E���6�ŕ���h�Q.��Nj��^IBJڔչ���Xd�nf�ؖ%�`�����bX�'����'�,K�����9ı,O;�v�<�bX�'�}���%��,�sMND�,K�~�g�~A9"X������Kı=���x�D�,K����"(�eL�bt��r��6���7rۻ8�D�,K��?Z��bX�'�߻x�D��Q"v~���,K�������%�bX��O��s&\�.�mə��"X�%��w��'�,K����Ȗ%�b}����yİ �Q|�!���ʈ��G�9����K�L����̍MRsSR�4��&AbX?w���Kİ�=��~�ObX�%��۟�ND�,K��ݼO"X�%��?vrM?f�swl���84�]���Z��N�4��v�yn���`����˹�[���D�,K�w��Ȗ%�b}��ڜ�bX�'�����)��&ı,�����Kı?��ԥ�3��4�5�˛8�D�,K��v��Kı<����yı,��59ı,O����O"A��GuBhי*IR���HT(@�w�^8$�H>��&�$O�{�;8�D�,K��v��Kı=�ҝ����d�m͜O"X�%����"X�%���s���Kı=��mND�,�Ȟ��^'�,K���L���e�2˙��Ȗ%�b}����yı,O{��S�,K���oȖ%�`��y�Ȗ%�bp ����۸��,9e[یPq��Z�k�����v1ʷh�3;�uV��N �s��`���{JD$mpFd9R���Q@��lOl6�u��S2��c��%���Xm�5v���ls9�fB�Wt��sѷV�nn���D4n�Ş��v���l���[��ܽ��E<f�î;Q��H�M ��γЯ8����k7��C�4�!��0��%���
\mն���p;gf�˳��0�g�p<]��]k��]\��{��s!�f�p���[wg��Kı;��֧"X�%��w��'�,K������Kı>��vq<�bX�'Г��ɗ7�vd��S�,K���oȖ%�`��xjr%�bX�{�;8�D�,K��v��O�S"X��b�ّ�T�jjX�����L�����jr%�bX�{�;8�D��@XdL��~��S�,K������yı,K��%�ۻ��s4����"X�~D�������N'�,K��g�T�Kı<�����%�bX?}���bX�'z}J^��f廦��sgȖ%�b{���ND�,K��ݼO"X�%����Ȗ%�b}����yı,N��7��7I��.�rte�8�n0�;�'�5F�m+�Q�F�k4����	ɒ���lܚl�r��T�%�bX�����O"X�%������Kı>��vq<�bX�'s�ܩȖ%�b{񥓹nwHa�q��x�D�,K����z�A?	��<�b~��=�O"X�%��~��S�,K���oȖ%�b|g�i��ݒ͙as4��Kı>��vq<�bX�'s�ܩȖ%�by�����Kı;;���bX�'�~�.vf�I��-����K��O�(lO�g�T�Kı>���׉�Kı;;���bX�'����'�,K��t�72e���ݙ36��Kı<�����%�d&/B��P�x���L��L������%�bX���mND�,K߶Ϳ?3q��psvx%ج'��t�y%x�ET��)ΐ��sԸu�d�.��1�yı,N���'"X�%���s���Kı;��ڜ�bX�'�߻x�D�,K�}I{6�����-�ni�Ȗ%�b}����yȱș���s��Ȗ%�b{�{��<�bX�'g{��,K��O�K�<�ܷt�f�f�'�,K��w;jr%�bX�w~��y��Qz���X��.�<O�*pȟD���ND�,K����q<�bX�'ӳ��9��˦�w37mND�,K��ݼO"X�%������Kı>��vq<�bX�'{��S�,K���^�3�B�7����Kı;;���bX�ʟ���{�8�D�,K��s���Kı<�����%�oq�������^�Emd[�tgn9���ۃ7J�#n<���U�g'\kBn�9,�م�3LND�,K�~�gȖ%�bw���9ı,O;�v�?=��!2�����	��#pV�I�[���6����%�bX���r�!� ș������yı,O�����bX�'����'�? ��2%��Ѵ�.jS�TI3M²!2!{�{��<�bX�'g{��,�dL�߻�Ӊ�Kı?~��jr%�bX��>���d��L�Ͷ\���%�bX���ND�,K�~�gȖ%�bw���9İ9�!i�� z�C�Oɾ���{��<�bX�%��IM���73Kd��br%�bX�{�;8�D�,K���Ȗ%�by�����Kı;;���bX�'�����v/#�dŜhuv��'[rQŪ^Oz�0��.��Y��j0�n��L�u�˛8�D�,K���Ȗ%�by�����Kı;;���L�bY;������L��Xh�:�EH�QNff�Ȗ%�by�����Kı;;���bX�'����'�,K��w;jr'�r�D�>��n~�R�7����Kı?O߸br%�bX�{�;8�D�,K���Ȗ%�by�����Kı>3���7-ɳ.f���bY�#"w���q<�bX�'�۟�ND�,K��ݼO"X�KР���)�d&Bd&B�����p�3&ۻ8�D�,K���Ȗ%�by�����Kı;;���bX�'����'�,KĀA��P�!b0F	�5� c��$!! IB4 %��qCWCHȐ�:��8Q��)�-@�MV+\TX��2
|j��R	HD5O����'��1 �0�L�\&��j�!V��
aB݁% Ќ&���D�'���@�Q�=#����9��̠�L 8Or�&o2�����!'}G�4��2����Ov�__}��~���	 ��  �kν9�%Ѯ���6�v���`*U���dt3�a�q����ma���L���:S�Yƹ����r6��#u��m��vB�Y^6
���+[���p5kdY-���ib���TPV]��V�,6x3gI�ݒ�����_:)��^����^�Z0b��u�q��j06wa�`nخ��T'\�x}WUK�;f�$ɇ�r�J�۬��/3+�S����X�>ܐ9;c�5b"A�q�]���ُ�*+�7X���d�g���Z�ъ�{]V���r�.�`�:�������x�-����]{����&�!�:�5�d�m[��z�z�eZmm�L�ۊͱ�:�`M����'�ZK��a�{,2��ԧ%ny�ϴ8Kƥ�Pu���ݗ���2ۣd��۶�W2��^�P�Փ�z���Bom��h�L�B�9�ݲQ�<�Jh�v�h��"eV�%���p	�ݬY�v@��V_!s�wɃH������8��]��˝=�Dn�6z�:��K���nqn-����m�v�>�& ����&���xTwm��mS�l�=`�{
�uS����
�J�[u\�xd�^���ƛiZ�uO��b�K���dl��8��R����Ռ��z�8M��ۊxC�rY��Z�[���)�t��mq�e�omaݍ��nke�`��6�6t:ܖ@7B9���ʫUR9��d^*z x�CC5�1�&!MHcQj����-�&�Ut���i,�;6G�k�F�Mї��Z=<4=���d��l�S�5[n�PI�q�u�Q��b�y�͸��mB���vn����&�݁�ۊ�l�N��u�jKZ=,�s����=�p6rbֲC�9W붖�9��h˩z�Z�v��"�N����-�S�:�8���v�C�ރ��6!�h�4���g�vN�[V�h�^�J�x����[j�5<q@��!�ͷ.\�d���swwo�"z���|���������R���p�U`�:�� ��x+�>��6�.�d����-2��6�/ej_I����2���w�:�mYk����[l�[�i!�e۴�a�ќ��m�8v��.;p�P���X��e��;p�aӝm�q+�`S��^-A�,�,�JȖE#�u�oE]���y)#r�b%(�줁qESƽ2��;��(� gt�\O<{���HyH�۶��� E����naf�z	k���ND�v��Va�N�낌���:����vͨ23�0���oq�ı>�����%�bX���ND�,K�~�g���Dؖ%������Y	��	����g�#�t��i���'�,K���xbr%�bX�{�;8�D�,K���Ȗ%�by�����O��L�b^������ݛ���M�19ı,N��~�O"X�%���v��Kı<�����%�bX���ND�,K�>����ٹn��\���%�g�@ȟ�s?Z��bX�'����Ȗ%�bvw�19İ?�&D�����yı,N�Є��ݹn�5��ݵ9ı,O;�v�<�bX�'g{��,K��߹���%�bX���mND�,K�~�e�+��[��6�%�*a��+����K��X��y�v�MD���}����qk>���%�bX����19ı,O����O"X�%���v��y"X�'��5�/�L��L��r[R��K���$�i�Ȗ%�b}����y����C� B���%����mND�,K������%�bX���ND�Ur�D�;��ٓ3��fə�mݜO"X�%��?g�Ȗ%�by�����Kı;;���bX�'����'�,K��wgvٗ7��rfm�Ȗ%�by�����Kı;;���bX�'����'�,K�2'��:�+!2!2��d���)��asoȖ%�bvw�19ı,O����O"X�%���v��Kı<�����%�bX�ȣ��ǜ��ɻ�G�]�n^����+�z���ղr5�c�3�:9�_�G�r��sssrnf��74��%�bX����Ӊ�Kı;���ND�,K��ݼ�	�L�bX����18Bd&Bd-���r:�QU.h�_D�,K���T�Kı<�����%�bX���ND�,K�~�gȟ�TȖ'g�B]�nܷM��\�ʜ�bX�'����Ȗ%�bvw�19ǀ��$G�	h9�;�s���%�bX��s�S�,K���^�{��]�1�6�<�b3�JHZn����	��;������X�'s�ܩȖ%������?[��	��	��N�j_�D�(�RMM,ND�,K�~�gȖ%�bw;�ʜ�bX�'�߻x�D�,K���Ȗ%�b{���ޗp�L3n���ué:sբ��h���et���]�=��Xr����v�U-Lۖ��fJn��L��L��S��"X�%��w��'�,K���xbr%�bX�{�;8�D�,K�Iݝ�f\�.\�L͵9ı,O;�v�<��G"dK����'"X�%�߻�Ӊ�Kı;��ڜ���2%�pY;2:�I��69�p�!2!2�߸br%�bX�{�;8�D��"~�����Kı=���x�D�,K�}I{7wsl��-�ni�Ȗ%�b}����yı,N�{�'"X�%��w��'�,K x*'DA���&��'"X�%��{l�w<��%�5�˛8�D�,K���Ȗ%�by�����Kı;;���bX�'����'�,K���;�WWF��c�p�M�� �4����_RnlԺ�5��-��$�#v�5��Z��"X�%��w��'�,K����Ȗ%�b}����yı,O����,K���^�{�
]�1�6�<�bX���NC�r&D�;�y�q<�bX�'o�9ı,O;�v�<��r�D�:gr�/�6eɳ4���59ı,N��~�O"X�%��w�br%��!�2'����Ȗ%�`�����bX�'����͓ٔ3&ۻ8�D�,K��v��Kı<�����%�bX?w�59İ?�2'~Ȗ%�b}	;���2��r��f�Ȗ%�by�����Kİ�)��xjyı,N��~�O"X�%��w�br%�bX�}���ۿ r�Yu�:I!9e�'@��28�;T+���sȉ�J�7���F�*�1�A�p]BC97a��F�F	�G>^�sn�i�+�zݳ�Թ3���9�Lo�3��'L�­��8����l�u͎�]7Oin7OW��v:�h�FMv��U*�v���ݍٶ�2e�֐su9ѪМַ+�s��ٲ�aR��Mq��1��z����禑�p�Oޏ'���X뤮��kau����n�z"9�IK��i�����.�m���Sؖ%�`�����bX�'����'�,K���ݱ9ı,O;�v�<�bX�%�������ٹ�[���"X�%���s���Kı>��lND�,K��ݼO"X�%��{�S�,K��~�K;�]ے�l�����%�bX�w{�'"X�%��~�gȖ%�`�����Kı>��vq<�bX�'ga	w���ܻ5��ͱ9ı,O;�;8�D�,K����"X�%���s���Kı>��lND�,Kߍ;1�݅)�q�6�<�bX���ND�,K�H����q=�bX�'o�9ı,O;�v�<�bX�'�?�~|�rY�i�/z��d��]<q�i�>s!�e��f�i�]�C�5��n]��SȖ%�bw����yı,O����,K���oȖ%�`�����Kı>�w��̹6�̛n��yı,O������d�� }@8ȞD�3��oȖ%�`�����Kı>��vq<�bX�'���v\��\�t��br%�bX�w~��yı,����bX�'����'�,K���ݱ9ı,K�����d��K��l����Kİ~�xjr%�bX�{�;8�D�,K��v��Kı<�����%�bX��!{���f�il6暜�bX�'����'�,K���ݱ9ı,O;�v�<�bX���ND�,����7~}������[�Eqp�eMGCt�ܱ��r�e*�a��[.��iN�v4�����sgȖ%�b}��؜�bX�'�߻x�D�,K����"X�%���s���Kı;;K;ͥ�˳\����,K���o�~�DȖ~�Ȗ%�bw����yı,O����,K���N�gwaJn�eͼO"X�%��{�S�,K��߹���%�����E`tb����U��'�3����,K�������%�bX���\�2�74���jr%�bX�}�|�yı,O����,K�������Kİ~�xjr%�bX�d;�R�L�6̸M��O"X�%��w�br%�bX�}�v�<�bX���ND�,KϾ�O"X�%��3�ۛ��5��d�;s�\�ivt��1�D���ܖ��Z�Ξ��V��3�%٣{���ı<�~��yı,����bX�'�}�8�D�,K��v��Kı/d�gs-��.�m���'�,K�����@#`�'�}�NA$��v�$RD���ȟ��S"X��������ɹ�[���"X�%��{��'�,K���ݱ9ı,O>߻x�D�,K����"X�%�ޟR���6n[�i�n�Ȗ%����;�����Kı=����yı,����bX�| b��"oy瓉�Kİ~�il�6�w.�s33lND�,KϷ��'�,K����Ȗ%�by����yı,O����,K��Ͼ�ͻ��7we�K�����0-t'�����Ξ���ͣ�d�1�k���9L91�݅)�q�6��ı,K��p��Kı<��vq<�bX�'���Ȗ%�by�����%�bX���\:lː����i�Ȗ%�by����yı,O����,K�������Kİ~�xjr'�L��,N�?w)i��ٗ	�vq<�bX�'o�9ı,O>߻x�D�,K����"X�%���s���Kı=��l;����2e�f�Ȗ%�by�����%�bX?w�59ı,O>���O"X��I�;�����K��	��ve����f�Ӹ_�	İ~�xjr%�bX�}�;8�D�,K��v��Kı<�~��yĳ�ow���|����]flVit��Z�&��9�]���k�Nϙ9�z�ά���7dv�ƿ�O���w��L�]Zɷa�A���t����rW+�4Z\c&=[[�դd$)�f6�)�[�OC��^
�lC�t��6�Zv�W`��m�S��d��Ϝ�F^ �6]���V\g�\Bx(v�ۙխ6�8]Ԗ!�q̎���Y].홷)�͘Sf�5C� 9ko���������鲺-�uͅ�pr�qk]�^[����v�gKpn�i��Kı>���8�D�,K��v��Kı<�~�����*�L���Z�VBd&Bd/ykM���n�]�]�sgȖ%�b}��؜�bX�'�oݼO"X�%��{�S�,K������%�bX�G��w�K��f����'"X�%����oȖ%�`�����K�?�R�bwv�\/�L��L���S!Y	��	���f9��0���\���%�bX?w�59ı,O>���O"X�%��w�br%�bX�}�v�<�bX�'�'�)p�Xn�ss4��Kı<��vq<�bX�ȟ� W����b{ı,O�o����%�bX?w�59ı,N��v��&Lݹt��&�cvx<<���/%�L�g��z�gk<��urct���f\&����%�bX�w{�'"X�%����oȖ%�`���Ȗ%�d/����|Bd&Bd.2�)�sR̙t��br%�bX�}�v�<�`�B}P;Q1�\@48���U���;�߿p��Kı;���8�D�,K���ȟȩ�2Bd'�b�ٖ榔��69�p�!2����ND�,KϾ�gȖ?�@�Dȟ�o�9ı,O{��x�D�,K���;����73Ka74��K��P��=�|�8�D�,K����'"X�%����oȖ%�`���Ȗ%�bw�Է�<�w2��ۛ8�D�,K���Ȗ%�by�����%�bX=�xjr%�bX�}�;8�D�,K㴛�n��ٗK�:��mX�T�Oe���r�J�*��x�7�� ����y�%%�f᛹vi�2�؞D�,K��^'�,K��{�S�,K������%�bX���lND�,KޚY�gwp�soȖ%�`���Ȗ%�by����yı,N�{�'"X�%����oȟ�*dK�'fS2~6K�.]�59ı,Ow��Ȗ%�bw�ݱ9��L�b�C��AS�$ ���F2�(�P+D�U�HVYU!e	H�Ԅa	RQ`A8n��r�P����Cv��3!a2BYIi���XYX��e��3�I}���e˺M2h�5極�OBB�s|�,T_#R!IOSP��%!D`��	��/��q_ �E��X��H�s1)���M�g�q ��q�� ��R#d	V	B4eeeHQ�QaIVYuB�\�@��)�� �� T#H^%�S/���*t<A � �U�( &(/��ȋ���ȩ��"Az�+"�� �ER���=�y���%�bX=��59ı,N�;�R�L�4�.n��yı,N�{�'"X�%����oȖ%�`���Ȗ%��@&D��|�8�E2!2DF�9&��K�MS!Y�bX�{�v�<�bX�{���bX�'����O"X�%���v��Kı?�P���?��R�ͶKvi� ����j��@�2<B۳�SNJ�:�n6�G�L]ܶ�晹�Kso��Kİ~��S�,K��s���Kı;����)<��,K�o^'�,KĽ;J~����ۙ����jr%�bX�w�vq<��r&D�?~��br%�bX��{��<�bX�{���bX�'�>������t�n����%�bX���lND�,K�w��'�,�F �����bX�'���Ӊ�Kı>�e%�&m�ܻ����'"X�
��߹�׉�Kİ{��ND�,K����'�,K��<^��ȗ�����Kı;����;��&��7oȖ%�bY�{���bX���D
�������%�bX����lND�,K�w��'�,K�w���.>�״ÖL�5��Н��wn^�D�&�VI0p��5��}��~�H.�2r�kK����D�,K������%�bX�w{�'"X�%����oȖ%�b_o����Kı;���K�.a�L�M����Kı>��lNC��D��ؖ'������%�bX����n�"X�%��~�gȖ%�b{	>�ݥɛ�dˤ���,K�������Kı/����r%��$2&D��y�q<�bX�'o�9ı,K�>��{e��3s6���'�,K?���3��ٺ��bX�'���Ӊ�Kİ~��jr%�bX�{�v�<�bX�����w�H�M���׻��7��by߹���%�bX;�����,K����׉�Kı=�w8jr%�bX�E4?^�����f��M��&��l��5�k������g�����n��/g�Ay&؝����9�Ոl�/.V�v�li.�6�Г�\�j�9�![�����{m�>���V��w����q�O=oky8ȷ\-\�������ؠ��i�r�G�Gt�i�����m]x�H��Y� �v��m �vz:#��l���ێ7/�n��i��*��s�{��������-݊uDt9�]�v��v�`�Pݑ�N�˓����]�qkc]�S��TK�4h�kK���>�rm~B���{��}���'R#�C@}�-��*@r=��l��¦G#!2$�Z��{���4��D$��Nk�3�����֦LT7Tnf��ﾾ�/2z���;��Q�����Ɉi�������W�UQ�����T��{)���x�="��tm�G�\���ч92��k�����F�g��6c��3�������z�*@r=��X9�ր<�ǬsUD��4�Ӱ9��ڱ$�$����!(�B���7��`s'5����vr�G\NH�������Қ���?�bW��h�繠u�X�O^Hɪ�R����Nm�;�`{�W��yzS@��
�H�����@>㖀�\�HG�@u㖀��~�|ݮr��]k
an�
湴:j۱��Wj�˹�����L;��7��j���[w�����HG�@u����X^w�T��E�~ra�73@��a{	DCgvs]����`s�ɵ{	/(Q'���ӟeR�\��Q`g�|�'��ݼ�����0� F����.s�ۛV7���� �a-MK&[�/v�z�����@7=��o`����P�.U&�C�Ą��=����<�!s2������q�Q�v�g' ^ܘ��'V�t��׹�lY,��N9Zޱ��J�sg�����T�&2�~�;&�@u㖀��-޹��2躞���H�N����33�?f6wӾvf�mXw���%�գCغ�����qh�~Z��{��Қ����lf�$�d&A9�����Q�Js7��`wv�X����	Bp����`�b'��L?~�k�h�Ӗ7TX��&�s47�@u㖀��-޹��U_p���� � � ��}?_��,���f�Us[�^&�z9s�eJyI'=���P{u�'C��r�&�i�nn��A�666=���� �`�`�`��w�� �`�`�`�����|��������|������;ɓ��f噖�.����lll}������lll~���Â�A�A�A�A���ׂ�A�A�A�A���ׂ�A�A�A�A�t������73m�6�A�666?}����� � � � ������ ؃�� ��A����x ��������llloN����6���f�e��� �`�`�`�߷�� �`�`�`��w�� �`�`�`������� � �("�{��=8 ���Ғ�fy��M�������A�A�A�A���ׂ�A�A�A�C�b�����x ����xpA�666=�{��A�666?ȇB*@�Pm �#�E�V$yO�fg��ͳ{w�7�q��C�;O5������ �u��a�u����୎��ֹ�x�6{=	��Q�lugi�<��f�H��]�ڝ��Wl��^s����;&��5و�qs�ۮ3�r<f��θݻi��Ƌus���)��lgH�@��ϵ�7;Wm.�Cqc^u�[^�iK�狧[Z�A�x�pv��t�uTѶ������Ѷ/1�����t�}��su�[�䥱]�K��[���0�j�Ll1�Zz�q�	�P���z�.��3.m�A�lll����A�666?}����� � � � ������!�r66=���� �`�`�`����Bf��ٹ6i������lll~���Â�A�A�A�A���ׂ�A�A�A�A���ׂ�A�A�A�A�������lll{�vv����Xn�L��8 ����x ����x �o^>A�����<8 ��?w+r~��&�6�m���lll~������lll}���x ��������lll{������lll}�I��~���fe�K�x �o^>A�����<8 ����x ����x �����sJ\%�4݃y<�� �Ŭt�V֫��,v��V�ո���!.m�۶��ɛ��˛x ��������lll{������lll~������lll}���x ���/音nn��i�Y��pA�666=�{��A�#��P�>���A�6?������A�A�A�A��{�x ��������?���A� � �~���<�70�ݐ���x ����ׂ�A�A�A�A�������!(dD&��ٵ`gg5��C��iȌm���}V��^������g��_���c�����Z���Hװ@u㖀��-��瀞�_��t�%31n1kg�nW�c�l��9ҝ��惀�	r+l��g'����9��������-Ɏ_+�r�������K'��)�|@7���/W��w�)�yp9E�Kha0Oo$�w>���~�p��c�xpZW�Q�&�@q㖀�ܻ���73n�ʹz�*@>�������?b��~ZEX�k��F�4!�3@}{���6z�}�ր�\�Ht�Δ���엘���5�cKΓ�V�M�!m�������6t�\�������x�91�@w�b��� =�E����8�F6ۋ@�@�ޯs@�zS@��U�bGu���pq��miy�h�R��x�91��9�Y�`��bƓ��޾�@�����O;�v�O��0P`�������Aw�����\�p��C�U7TX����}V��Jh�Jh��'4I	�v����q���y.��f�l�WM&��u��xN�(	�EA,q�M�"�<���=��M��O���/;��
�W�'��	Š{�R�{Қz�������j���71�	Hh�l��91�@w��	t\�r&�9i�@�_U�y_U�{�R�{Қ\�`�!�$r#mŠrc���e��`�}�-+�W�B H	�|�E��aƨJx��5��	F0 ȔX�R N��0��,�ĪFd��:��T��`���/ E�	#�jf[R�$�3jHM�0!�Յ-<�7
Ҡb,R z��C��)�H�e����O(;2aCX 20��0�a�ٯ'��P0P6%��bZ��ȟ}�{��{��������  �[� �Xh��jӞx�L�(��6��0*�.����Ӣ�a@��m��s�z9
Hֹ�F� Y����j���G�+e��������ӝͱ�Q� �u�d��u�T�lB�cj��Z��NdW�5T:��&���-�i��M�����*gm�OJ���	�i��&�ʚ�6�i�#�eݿ��F��T �h\�����ڪ�:N�+I�\��c-�\Wkun5rgVێ�7|}����z͓�4��,.��ݺ�dP���8�m�ya�gt��B�0�6�m� X�;Dg��r���U<�Q"���1�:���H��������&��7-��7n��-�C�+�	=U��7*�E�:���k�=b���Y�8Z��B�N�aXa[�Ob�N��Z��&�y�e���vsn�jUs�����%��٬�%�g�J6�Bm��x��-�^s�RZ�S�:�ݡ�pl���VJ��eڴZʑ�����pvZ�%c�n!g1��ף�)M���r��]���Vbs��G�6x䲩�!�6�u�.R�mX��q����}�p�l��!��=���Gɺ�(��J����J�۩n��l��ؓ���z"I��jxZ�*�vl���m�r��!KR��:�F��ɸ��8j���u�3ig(��˄,az��Ӝ�ՏYzI8F���^�����܅	�'mbwa���e�9mŒŇ���5K�pdgm�&�+<�dƌ�e�j��
�Z8��m�abָ۫���;l��^з�n�f�h�9�	����X�3��ԯ5ձ�vv등�Mb�=V��sk�6� ����9��W��z�=�������ێǎ��ʼP��ڲ9��z.�U9��s�N��+e�*�*PX�v��9]�*R���u͞��9{;Ne6'���Pe�:���h1���6˭�Ok@v���pZ;k�����	�n�kH����c �H	C\�����۝�u�i�ӹp�,q�*ݛC��r�_�{Ϻ�8�WU8��~�A>5@>�Q�E?	@pT=Qt�B�?	�w�?{~��i-�-BnH����h�wd��M�����e�.3F��4:�n�$��ÛE2��7��7����힌	���+��<G�����[H˺i6'%g�x9ņ��cm�Էmmf�)��{OjLteu����]�y5�����Z�4M筛m��77+�H(u�0O��O��Ba�e�O3��pE������ŧ��������?|~����]��M���,a��3�ț/X���<<�wP8�5�M)��5��L�r/ �R�{Қz������q���&,˼� ���r���;�{��"!��%ÝU�T�Q`gg5�d����u֖w+K��F�l�)��}V��Jh�Jh��X��I8�8�HN-�m������� �'�ɎZ�,7���f�8c�����<u��{N�t69�m��9����[LT�tcװ@>㖀��-��� $cM�ۚs*���sE��OqިP(IG�P�]]J�����~�M����X�JhrŊ�z����qh+ՠ;�{�� q�@w�p�f���5J�����D%�Q9�x�7'|��{���$�;�60�{J���,i8h����Z��z��)�^v�"��s��$�!�"C�7[/e�r'�Mu$�n�;X��3��ɍӝãu�L�����9h\s콇�����vC^o��� �6��72RS�>q�_��o׾�� q�@;�umT����$��=��M��^��~����b'(��(�?�bE"�������@�}�=������72!	H ���W�1�b<��.9��^�o�S���@�q����P�%�����]i`u�6�*�Nz�U��,�v�p+��qqu{UԮ9G�n���p�<��{��t�~u4nUc����{콂����:��&2Țqd��z��)�߳/Y�^w�x�W�r9b�"�$ō'�������}W}�Ob�^�@u�:H���Q4J��BI�k5�Oo���I=��{9'�<qR x�T�j�IC���`oPu:z6��72R/v��� ?W��~��G7����*��C�1��bQ�)�8�˪��:v�<]��u�׈�p��<D3q$�z��)�w�)�w���<W��9�*��I#s�������(�	�;9����ٰ9�u��(l����z�M�r(ӆ�yߖ��^��w|�Ɓzύ��X����܈��ʹ.9��^� ���r�mV�"i���܏@�ڥ4��6I���o$�^������(!B	�,������3e��훛�[��nJP�y�ֳ�V�Ƒ
�+uq�@��p��>n۳��Ƒo8(���o	�q)�Ӥ;<)������r�c��Z��]08�N�tj�8)lsYLv{���]qЧK���y�#��7g�{M���:�:7�9c`b�y��̌X�Z���0�5��un��M�ԕ�j�Mg����uFa�A��o���{��_���zY1K�ƺ�:��w
f�j�۞�M�i��J��7͜�ΐ]ld�;��' �����;��h+���T�����12�'��)�}V���13�sf��u֖y���;�5T�%�&ژ��@�}~z��)�w�)�r���9a�\�I�1��I8�}�`�}{���=UU����� %��/��)$��hBR{Қ/z��z��j��<��+�,y ��Y˷\�]��}b�<iޙrF�2k]X�qH�E b�8h�����}�S@�zS@���,�f�G"253S`|�7P��U	��Jg{���;�Zh���y�*x�'O�nG�{�u���v��Т"x��6�́�+0ȏ�LX�p�;ޔ�9{��+���T�����1:�����W� ��@{����������g�����a�m����On&Ryɗ�Tָ�������u�����i���\s��װ@;nb��ʉ8�8�I'���)�w�)�Z�Z��z��b\��I#qK�Q`w��,��v8QBI��1�pXY��[w{��)M�%^��R(ӆ�&Ih\s��װ@9󺻈f�G	�H�Z��z��M��M�j�;����s�n~qG��u�I��1���ك��=�㫵bϕ��|�[	���y�(�Y?A���S@�zS@�ڴ��z'C"?91cI�@Lr��� 9%�ʌ��,�ȞD�4_U�x�W�yj��;ޔ�.qr��46��I����l��u���v���"&����'jV�F�������I>��
��#��q$�z��M��M�j�<W��>����~IŐ�E� ����]jm9/In�98����[�8���GVx-%QI$ncB���|h�V��^��S@���T��I5 b�8h�V��^��S@�zS~J!6f�4޹j詚)IT杁ǹ�`{j��;ޔ�-v��j�OqD�����mR�{Қ�ա���~z�8>I��ȁ��w�(��$�.9��{����u_U���_�۴�4u8�ʷjb��u�=j��e̤"�:6�)�\$�c[v��8��p(p���ݳ�t��n#hݬ��.�jݏU�����Z�
mh�vw��v�g���P�)�e�8�V�ۤ��<�am]F�q�\l�\�j�t�jy6���=Wl�U;�"Q�ZJ��-���z7�n���0�a� ���عމ��ۆa�n�L��䪃뀫͓f^��븳lܣ�:sւE���.X����������!�G��s�p�u·����?��Z��d�����+I���CiIqh+��ڥ4��4]�@�!r���I'�연@>��L���� 9a���:uUU3JX��BJ!<�^����ɰ�P��uޖ�7�ni6ڙ?(ӆ�k�h������>4��4�=������Ͷ�7�������c���Vх3;4��bڇ�ۏ\m!�''P�p��������r�hz��w>�{�a�v4�����mR�����U�w�Wy�%��%�9q�@x�Щ:�ȁ��w�)�Z�Z��4mR�#/��K&2'�)�j�/Y�{luh�Jh8�*��"Ғ(��/Y�}����_��/Y�Z�Z��Jۂ�������ntgv-ۮ�����ٷa9���n�[��.R�v�pUq,`k����?��w�)�Z�Z��4z��rIƄ(��;ޔ�-v� �����V��1#僧/��0Q�i�@ݝ�`gr��Ϝ	�B@!"�R#āā�>�����deR�YH�%�Dad#k#�� ��=�Ŋ �#0�`��歌�� 5�<	�����@g���4��uk"��� �C�>����&0:�����t:a��0�X]�}�����(��y?\�Px�~�Nu��!�"�@�1cH�`A�����E�@���>3�Il,�>`W��1 �"F+�P�D Ł#[n3)�	�dO��@��CH?A��|ji�I<C��f��σ�qB�!���D :���A�E�H�U���:����*x��1T���Ͻ�s��N����'�>��r��RM��uN��	7�ͫ�v��;��	<��vrZ֥UR暘ܼ��jM���}^8��Z �vhܪ5&0i��� �7�Yk�rO�W	�����t�����t
�7^�Y�Ѽ�aYy���䖀9��}�,}���*3�c�%�Ȕ����V�w*��̬,��P�%�S&�Tz�SE"e��uT���U��̪h�JhϪ�9`v.W�LQ�e�n�9Rl�`�o��_U��R�1�2� $�FJ�D�����*A)R$XA�Jȋ� ,
�������vɀ�k����iL���;���Fef��9��`|�+�	.tй'T��!zB����ѣ�.�b��i�FQ--�k��@�iΔ���v%��Q��m���Z �P�6���N��^b�*I��N��ٙW�
g�i`[gƁ����k*ǅ�1ŏ�i��T�o`�o��&�;V�!�ɘ�A�8h�)�w>�@>�ʰ؅	>-����-ZH�F�&D�(��;�U�[f��[)�w>��@P?�O�N~���Mvɛ��'NeM����ö���ְ��n�ZA�ۇ�iڷ��%:'�|ld�vնʇc�������dz틟S��gFy����ݽ��@�l��Mm�Fn�slqõӑ��{i�䄲\��Vxx�f����EŞ���)���tX��$��	n��4t$�W�q;F��Z[ �z遶�����7sΪ�ñ9��la�֬Z�^/jw绻���{���~�����2ÓT2ܛ��6.5���mX��1�k����n'Og�u$]�JH�����42�M��Zs�X��4G&�����l��$�M������v�fU���Iq�cb�HhϪ�;�U�[f��[)�ym$ީ18܁�'�r�$���I�A磌�g��*��M��1�d$R-�mz�l�������Z�|+�&<�����n;:,a�dwNo & ����quc!��SA,�E����rhe��s���h�٠{�=*e�d�q�e͜�}�}��_�*4�P����~Z��}42�M��(��LDO"�-��Z�he��s��\������Iqh�٠v�� �- �Iht���7$�7JG�{��hg�̶_��Z��h+k�?������o��A��=6Ň5�ǆ�a�y��aۮ��i��9��2B6�j<lX) �ߖ�����mz�l���X�fɍ��i=�x�9rL@r�� �-~���#�U��̈́c��H�Z����<;����ȁ��@$B1!A^���?~�<��w���䇼�U�*RAE����e��z����@�^�@�A�&X�L�
\�`w��v�IB�(YY�O ���ts�)�^��#��q9�Hc��D�����[;l�P�Og�]z����$��ɍ�9�1,���EZ��^�ⶽ�K)�w>�@�K��p�cQ)�z��zM���o�b�U�.�R�`�90�Ē�����@�}V�����<Vנr9`�֢��5@����@v�� 9rLA�>���Q��TV�P ��FG��'�率��=�	6l��9N-��W�$�^K��zxa��`w��v�Ub���P<ޡ	��ٷ���'[nfƖҮ9È����d��<[���Nmu���ۗ$�zM��r�}��r�۞��y�ǟ%$X�A��凜�;�S@��rl�fM�S&�kS�mRSR�h�7v�X|�M�I�=ݛ�6��9r�VbY1<�Hh�z�癓`s�V	(y���Zj�h���JA��ⶽ�3�woǀ[9����rl�Pt������CfI�a6��k	�1"e�4�r)�d���$k�%���L�&�d���L��M4�^ �D|�u��\"�qnܵ���j�Y���n�;���5;l:V�|����'��μ�Ji��4��@ޛ��t�v�����9���6@�q��v���#%λ-dͮz�{zy��m��k��'	���oŒ��0�����ɢ��pRl�pۦ�s7K2f�1���l�=`��u���.�S��Ͷ�=K�]n�LG&��R?@���w>�@��r"%�=ݛ6�n˧U4ƣH�������W�x��@��+����9���̓u-�5@���`;s؀��1ޓ`�o�e;���̈́c��1�����YM��Z�ޯ@��ʱ��Mc��z{/`�o����\�əWg�k�Ɏƽrt'-pw+��\v%�K,��e�����~�H.�c'M�^a6���=hm�@r��}���,#��b��i6�2��u4���&�C�!�Z�b���|���3�O>��M��Z�,2�Ĥ��R8����e4��ߖ��ߞ��G;��b�Ē���e4��h������K����)x�;m�@r䘀}&��r}��z��-�p�g�4�CMɮ<ܧGK�t��t�:��k��\Y���� 92K@>�`�o�e;�ZoH�$ɐbq�Wj�;��hϪ�=]���XQ��Mc��;�2��;��;J�P�b�t�6ll���N�e!TU9M1�{�Z���&Ih?UU}q�^��|1}1,���EZ�����ZzYM��ZٙY���Dx�D�&�m�!W�ȈG6���ļ�*��݊5�g�x6y�p���H4��~|����s�Wuz,9�H�#Q��;�2��������͛�v���bV�R`�b!�w>����rl�
|��vt�������37C�j�KsN�aBI�s6ll�I>�w{9%@�ċ"F!��!�	��oo$�t���s96�M�?F��@�V�ޖS@�}V�yڴ�-in9�����Q�L�E��l,q�P&�u�/i�8�ᧇ�=l&3�}4�+>�37�� �-I~����ݐ���6S�~n�TU9M1�{=�~������v�́��XXb�F+1,���EZ�ՠx��@��)�w>�@���,Q�JH��˒b�l㖀o$����#�mD����)�/�3���o;��$�s��'/�}���"���@"�����+�pTW�pU��ATV�
���*��� ���+� EQ_������E ���U�TE�U��TW�@EQ_� ����*���ATW�ATW���e5�~��@8o��?�������;���`+�U ��h��u��h J���4j}ž0    P

I@PP�� �
�  � .� �|   s�����V�����V}c�OF]X[t4ӻhn.x��נ�Pz=�lr�q�#��>����*���W�ӡ�l:tǦ����t�'P)��g�1���w�5�G��|��o`h{��i�n���� �8�>te��;�={�-XP4��:ܓ\�����m�ס��85�ɦ����ݎ��w��>6R���|� ��5���º:iѬ��+�G�P�ACo���{`(i��`���  �h�� ��^��ɷ���cT  �Ǧ@�$�ʣ�S���aF
�w���C^�������ѣ]r�t��P�@���B��He$�)�02   S��R��� � ��d��"{J�����  4    �Ѫ�2�(�4      !	��M
zjz@ ���5H��M
~��$y�?T����4��>�?���������?�/��QC\�����;�f6o��N���:�6��؟�������h�"& (�;�m!k�����I�V�f��T��d?��W�����[s333333333333330ffffffffffa9��������������������������Nfffffffffffffffcm�ffffffff���������������������������I3333333333333333333333333$�ffw��{����ª������������W��ק3�����u��M�0��F����ޜ�%��z����i�-��b��R�@X�� *����a����E�p��.D��iu�<�;�_<�2��HK֯UG�F�^��
|HS!�U2r�I�*�!A~�(�L����A��ep�dX��0ӢYv�^�#1x�
HѢA�$�W<�$�V���6�[e[(�Zi
"�"�S�-s��*�\$v�x�u_B\0r�fBO�K��v�l�1��:zy��-�8�OMSP���]�?��C���93���{��1(r8va~�+�3�\�v
�)ќ$�;�`��E9Kze�� �X����Xw����xPB[�`�h,0H4��`1J���F�-�!41����2�����[U�i�F����@B�HH��1�4Pr�R�����h�	��LB�U���aR�!3I��!�������u� D�l����@���j�B�VIέ�#���!l��i��u�Lx�x5����
-�46� ��f�H�����m$�]�qh�.n7Gz9�R�̥�6]$J ���Ӳ�Mʹq�%�YM�%Y�R�0!K
�T�HkICqU������`�N�,�)�F[UF$2��PBF�VY�m��+���E�إ��D���eQ9ta�0�ر|�|��F���Ai��\��s�¼�0�l���u���u<P�"�f<�&�`R��z�+Z�T
�Um�Y*�e\su�UH�)#ز"�g���-�[��xU��pe[���B���m��[�r�Q�c�j-���s��Ӌp6����M�a�SB����@%��
�v
`�Ȥ����*SXNa
!XB��Q)C�M�Ja � K��樅ͦ��H�	�m8����)��	E��E�ܫ0�A��nQ<�[�/A
��i�Qp*B�4]4�"O<�$e�1n75����#��N�ʤ�NÃ8�2Q(�HQ��iɰ�o5�9)���Dh�Qd(bnQz�u�L�':N��u�t$�!��nYi
mՐ$�"BT+�48�:�AH������B��7��0�!L�Z��e�x[W&\��@�4ib�cE��M��F!M���RG@f�v�
ma!"K������m��W��d.�$h���S`F���'Y��m�HA���R�q�B�C	W�!� �VV1��bj���`7�Qa0��.�*�5��~kA�x��^}~:ۺn�i�1�JBsG0�Vʽ΢k�0ᡅ�8�'m8�s�+��q�9�s7B0��R��%Y���H��0\��H�g`$�%0S�)� Z��M�zO �TE��FC
����|M�Đ�E��X��h�#�X�pζ<�w���R��p1ȔjbE��i4
LM&�%6��!���Q���JT"��H�I����4i�g�
l1	� E�"Qnkg8�8@�.ԅ^_��\�lx�pM��4��4o|NJӳ�� RXa��`b�^��h7��X�@(2�k5.�#�RDH��\|�),� ��0Xi R���G^!��0h|B) #Kc ����b[pL�FF��;ӝ-�Nn��ۤ��stv���N,�Y��A  ��hH�a���tݛw��p�n���8h,B��Y��`�X�L"�ZdJH��t]�1����Z�E��c�	Af:6��,�[	Vf�l�HSl
,�6c����0t��6�7��M�k{�^^�1�-aC
1۰ R[�����U�o%]\!�U�B  ��  �p�S�xtC���]Ή~+��,�G�Ĩ�����[d1�&ή#��0¹Q:avp�hp�Ē�ᓜ�c���c��F�M@S�����q!��R�"��P�R`�]%��L�JHq/t����˚+si
��:�<�������	߇�'v(� ���6x�Uy]�	Mr�]�^�?z�U�'E<<Q@�!�Ű��n[�{l	i���rR�	k���]*��\���.�2.�WR����C��1�!�B}v�8A��:$���$�h�ɾ\�N>_�	
�yw�!q
֥�^4�X ��ƚ �>H��@�ųr���NM����3%�%B�D��s!�RBC��UՕup�#t��ۊ�>[v�!9�j�ֆ3ٺX��:�TM.c̶D"i[ƍ��H����V��l�q��!��n���ډ�r�(�I᧞T��s�w�A�����R�C���h1�?p��y�I;�|���g��;�����#�m� �    �  m�    UQ��n��˗>.W�tt�����̽p!�=ujW�A4�JF����*|���N�Yv���g	�!1��^Xv�9�m��l��<�E*�-���&�1�+u�X�V���]�s;l�������;�E�lβ[(��4��U�!xJ�[mt+�m-�`ln�9 �JO5��ㅍ�*���fyH�8Y�G�� �)�mf������.��F�N��=�/'W��N���v'dڻs��H�mu�@ M���� ���� hC��+eb��b���gq�a�9N�ݵ�;, �,�1���h;�B�P�xjWF�,�U��3��mm:�FJ�n���՛��͹���	 t�d�i��6H�m�	>��ﾜ$��i�mmۑ  �z@-�۶�   �`$m�k�:M$�   �  $��mm��L[[-	� .�	m  m   �l[�^�m ��     8    �  m� ��   �� �`  m� �� [N-� ��m� �� ��[A��fٶ�h ��Ll�m����`m��   F� �F�BA���   m  $���m�6� �n�� :@   <�/[hp� 	l�6�#m���3m��%(  �m��-��۶�%f�۩j���;n�pF
�����fm�hH8$�H!&���u���-��6�� Ho��H���m2Ga#6�[��tۆ��[m��I�#m��ɰ�^r��ɰh�n�� ��m� ��6cn�V^h���]��@m���,鬦 �|���tn3�Hm���9"@ �9�\I'-�m���œmm� ��cuͲޠ�%(�][@UC���.�t�  �  ݶ&�l��f:�Wj��b��v�;qb x��uJ���p;kn�iΠ&%�}�G�eq���"MJn�	u���(ۻue����5$׷A�ݵ�  ���m�۰2 ��M& /Y)m���V�$ف���5�N�"�z���op -�  n��E��xq�$�Hh 6�I�	�k%�$mհ�T�mmZ���eW�+[p�[B@[� �@ku�8�D�v�Y�̀]g�i�L� I��Lۆ� k����(�P ���nVj��S[����~�An�R�܁���n�tkl��ll ���lm�  ��%�[�ےgM�UlUn�ʵVʼ&��:%��n�[M,ր� q�0{o��}[WM��  �m-��@n�m�����a���� ��Ӡ �gS*��ܒ�/�v�t�.#l N�lm��Kn� 6�p m8m�� .� �$ XI� �e�8����讠*��T�T�;,ʮ�4n��Εi	�m   H ���Jݶ	  ��$l�fͰ Ͷ l�m����K�ᵛ� Ͷ�am[Mړ��7�<���v�oUSEp [@ ��l[@$6�-�N�[�M�ݶ�9#�� ��6���V�Y0[%8�i�&؛f�     h�8 ���a����IC�^�E�� �tؽh�ʪ���t��I���s���-6�H ���jU��.F���~��v��v�t�y�V�n�(x�g��l��G[M��6�tq��d��$4P9]V�e�=�  ����l��x  p6��6�pǍ5��Y2m N��!۷lp���;t��v�;m{�U� 6�  $�ƶ2k  8  	m��նI�*�t�  ��m� 	H-�� m��[Ii��m��m����%i0�m��6g� ��� ��m�  @�:v�[I pp-�#��\�l�i��  �$  [oZH I��mp�[dm&$�������Ѩ�'+N{dֵ$��n5��g���<݉�q �uT�   �`�h���-��lKУy�t��hm�  ��Ӌhm�m���$ ˒��� ��h m���Hqmp[@��m��B�oRKd�  ۶l���B��-���m�m�*ծoRA ߅�n�� l�d�	@�w�f��� �@�$o5l�����U�5}d3=Ck;v�j�.�X��� �`lt�� �UV�P倪��vU�@ 6���ׯSm��m�h �� 6�۰[@ �з�ⶑh  �v�Wj�kZ��vp�ؗ��l�$R�-��l8H�v��C�����PZ���U6�T��[ �G6ؖVݵ��[{={=��    m�m�m�D-�ր��&� $-�  �m   �`	 m�۰��  ��-��  8h����9i�۶6� [Kl���% ��d��i{u�v�Cy���e������b�]m	�j�Qf��_�I�OS�='I��ݠ*���� *�a q��n��%RVQJ�(�*=�r9̸r�[�[��$��q��Hq4���pq��:::4FD4p�����UT��UU*��UJ��UR��UT��UU*��UJ����c*�[eU+5U*��UJ�����l���_H���g�g��HG���*�x(!
ڒ�����M�<p�
��/L8�ī-BX/Uv�!�Z8"��������P�CO���K�&�q�,V ��L�t)�{�A� �  h8S�n�݊��=�uvx�<A�ǌU ^�%��B���RH��H���x�l@��ҝ P4(�E� ,Yj�P<=CJ��Ǌq�F�D�y�#��+@(�|3�;@ҡ�x� ��J���jDҖ�j��ݔ�)�E�c�@OԿ@x��P��Ph#�So�h�p<ZM
���!��N� �T7�`D�0J�4�<z6!`��'�N����Dꦈ"���!�@�i::R*���-�y�M'N"`dBBkc��#�[)4��m�<�  �|��lg�`��XXX� 7;].�˻���yW�yW�yW�yW�yW�yW�yW�yW�yW�yW���i��m� @�i��5طwe��wv]ݟ������:���l��)"S�I$�@~ v���ou����R@��]B��A& ���F~�k�f�;�S���)~ $y����,庬�7`��L)�+35Z���6�Gn'�[��u^�:��+�m�U�{qudD�D�CG1�iK�q��L)bkpX�Y�K�A�2k\AJ'8��m�`�����h���[x$#�uf,�3��/Zٺ��0��5vl�)A��T��S»G1m)�-�N��� �Ν��2E���rݗ&�6r�=k�Ye��*ǅb�i1�i�@b��.]�^��U6-�p�� $]il�3hʝ9t�U{7&k�q�K�K�uy:Ո1���AVl\8̉#����������mAp�b�m��=��ݜl�4���3�U��n�^�9ds�e"R��kc'�w�O9}�t�R2���nOe+�h�cvM��e8	T��k��D*tG:���԰u6��5�p�����ۧ59G�����MT�-�x� q��G���[ t�o&�j�;��)<�����-� [Q�����\���J:�5�{rv���]J�n�lEnh6���D5U�$"\�힍[a��ݘ2UV�e�P��V�v��t�v�	��F;MJ���ϩ1>��iH
��E ��AD#�C��
<.�~���
�Ta�����u�fVVnT-G/c��U�5h��=	���=�ݲ�R�K�i��Ý�L�����"�V՝nY���⬛e�
�k������'Uݞ8�ؼ�e����5,Y��0�̻��uW��b�A5UJ�:;m6�h��&�TRi��ơd԰�K,��o�f�'���vL��� ���|�����q	$tsڪ�{�vqk��c��z!R=�v���xjz��Ic;���c� ;�u���n���UW�M>cx��ë�s�p�5���jYU(4�$�QQ�"�I8�M�|@�:��1��l��'/2�WY���:��t����hH�Q��@š���Yf5��i�b��q�ِ}P�_D����U��גWٙ�C�N���y�<5��.�&��\�x|zi���W��Y"8��ƻ���'\�1>�Icm$�����L2��.�u�\-�=�h"��i"5��v���X��Jz��R{r���c�0����#m�w_I�G��g������n^Y�v���*���r��z�^:��9����#	�k3���]L�0��^g}eF��������HJX�Z1���
��r�/������o��/=�Y驝b�	�L�ېp�1���w�g1��1d�H�X��]�_� U w���X�8��T�3*3�{�5�s���0�i�
��E-E�<C��f�5�xt�d1�e��:��	�3��Y�)J<����yi��38ܙ�,4QD	�  �n���O���3��^!��4��0��{�g9��1��d��M�Y��o��c;Ë��������U�1��ޖ.���mI\�c��#��3������F�j�l6�#���@�m��Y�q�D�WS�,�4��YȆja�nֹ�V��l�x��?���l��2��]��M��b6�ᜍq�Ռ�ZAt�):l�77�3��øp]c��.(�-9����$�u�$�|򩛁�H[06a��M�5�3�텰e�8�������S1�s���Hd��f?����'7`��Rb�d���wN��<(���W�+<26�s:�Ofu��u~�ļ�A7,a���c9��1��W���� �e�m�JW�f�1���Ζh9t.t�sX펺�ݚOPsN��ydG'G���<7��D1�K���&��
U������i;�3RWwX�#��s%_9�d"I�7q�����k��vC��?T�C �cUU^�u��D�+Wba$$-!($SE��͙�&�.6��U�.��A%��:���@g1׏+:26؀�1=�}CH7�m�xu'�M�<�7��xZ� �5����'G�Fp�}�,w���b����������W�v=5��%����2F�y�Jf����"�`�U��tkU'��2��z�A��\�q'�@�>?
�(=�>�1g��A�|�T�H�nn��u�/C��˘I2Ė3<���0١XEJ؂QOA�(u\w�݇g�9$���s�����u�ޗSx�[�
Q�m��6&��6`�T��	��B�idaܱ�ƻα��W���	`���nF{�z�̐���'>nz�I������/��T��K�r��s��uVs���ĞT� \�w���9ᇼ��w�X�<�EV��ȬQ����+�+7d����Gab�71����ICLj�z����x�h��㱷&����P5pY�C�Z-�5�p�1�'9yh3"<qr�m�[\myMˋ��Fv���[�6\Z�h�$�=Β�gwwFy�J_~ۥ�-@m�ۑG^.5���%<׆[��1�>w��]su��1s	C ��{_|��Vs$F���]�u}U�c�u�s��(�	���Uw�c9��1��%��#	H��b����c<�y���&�7�]u0q�+1.#)����Cm�p�����W�:�_��/�KТb8����� =U�k��_�I��]s�ԞԒ2e�qWy��s��c�[��d�*����vW3��<����K����\�Y�cj����[M.�4�p��{L*(��l���������J���gq�qp.�Fi�,t��s����{�^p�\�'"5��y�;����%i&�I9�wwww�<�j�F�S- `���U�a.�hF��}��a<���ӛn��tW����VEUh�-ZP!�$�5� �cs-�ziΒ�[�F��{�n��:�ΉTKI5��:�֝c�,�ek��&Nu�)PJ�e��$*�����[tL|<q�V�f��[bml�"؉���Z�<��D5���c��ɿ��Gl�b��T��<
@/���T 	�M�8(?� >$oď�'��h#����P~�ۖrnVf���;�����W���N{�6G��{�_4��4Ğ�n�H��;UC��@��w]Ni��#�	+�s`�
ʑs�Y�����oWu$�����:��_��A��ߖ�Hc�l�y�>Gþu��,ޯ�)�V|I��$����^�#٨8�W������&OP�A(�u���[�a�P����5HD"�>����㭟~m�I��D��u��:��'3�8TSi���M��c��Z��e����h�r0��J;�ǻ�W��p�N��Nz����\�b�Mfu�xK�bH���b�I���s�ĞT�,t�U�u��uy�s�o.C��1��cp���3������(�1tĽY�ΗԬ�D�;v*xy�;��� e��lW`�QQtWP.{��n܍ӝY�e8� ']&lv�ns��pY�j�ힶtl�d��3��`�	M�r=ME��k]��un�x *�\F_
I
`�`)2�B	!x��1P�g����Bdz?���J�3��:e�vFZ<	���O7���â�n�=���bI���{ܨ7|� ��ޒ��>#w]�{����U��>?9�Ҏp`��~��P���_}�T���G$ȉv�L�m�[t�s�j1�d�	��+��t�C�w�#������9c�u{����X>��ϣ�^�y����؞T�/���/{�`����eA�Ks���&C ��>�Ӵ^1gH�P;ݸ��G�24ߨ;�şQ�cwϠ��p��bq�˂��X�D��5m�RER�E�	!���_G}����u{���C�x�9Q�������1�v<?��y���k8}�����~�����4��꾠�]�i�߄��7�lHԕ`sA��H����c���M�H�rǎ��=����ovot쯨U��NU�IAb!on0=T�#6����.����H`p�~�X�:����A�g�w��I��"V75� ��1à��8Fq���n�n��y@��;;�~�{�F�A�v7> �y��
�K���D?G�G���g�ܺ��̶��|+���X�} �aqi�D�[O����+e��>y��� �Ii�,�p2Ls�V��U�"���ߘ�@�p� �[�b�4l�6"�H=T7_	>J�U[��y��o����
M�F_F�W��7��E��{��B�08A;��(��u{���:�5�|��&C#2�S�>W\�s+���/��!��?Q<�=�V��UZjd�0RXZV1#��)�V�Z
���mH�j
d��e�L�ER[��9��V�ɷ=Qf�f<\�Ia*��5㭝(�O�L�ܝ�G5�`�E�L`��]+a�q]�*�WU�/�{�}I�Kk9�q���3����B�-F0m���֟����>��~�Gy�nD���x�� ��z�c�{�oI`����� �wүw�Pp�������"#js�~ߝ^c�x~5��8 �i:�2��IsF�����|��_�_;��&L@�-���K`�R`P�҆�M��E%9c�H> �y���@�c��ߦK̘^G�{�lZ�b6��QFĤB�Z��h P��U7����yn�=�8p��.�$�d���͕�͟
��Q}�+Okမo(;ߘ��P��{��xF�!2e
W875�u���ovx���,���[rI $�J���xnyշ)�M����S��>�=�:��Y�NǇ�[<�JE���~wu&:xQ�b'{
�IW�b�H?���k�|�ߪ)�:t�{�3��f1�q����y�W�燳�y���st֥�
X-Z�e�ԋ���U�n@Qp�?z���f�8��ޙ�h��$���Ş���9���/0��v:p�;�3��M�%��}�5��w�u=���y��J�}�q�G�OԼ��*�8>�u�y�p�I�uU-n�(��y��^x0:;qӮ���aE�$l! �J��,��gX�c�|��T�/� �w�g1���]{�n\�^c�]9��0�!��,{����,���V��Ԉc��n�u��
���G�g�s�����=m��m$�uU|�Zֵ�kS�~CA�s��`��F���)�wW〱 �,�	���2r�4q��%,�#�����0��c�R K�� Fɂ[�~Z�	�{�~J��h$�Fa�������9x�'�&�ݻ5�	ֺ^N��ZXNi8�Kb��Kr����F�k)
#bƎ��^��f:#�6�p����c��j���j��ï�������b]ZGh�M=����#J������J*�. �H������^�-���,F8��[%T�	ŘU	��X��@�u6x��g�������s��U�h^D��Y�R����Ձ`l��VR�F�\Ek��T\�M��\C@ؙ;P�B�Yr\�h|����#�NӸܗl8 �Z	S�q�v�.�n��,��Di�xcr�b�C�TV���pq3�!l�m�m�M�.Zy,
''M�L\�8k�gջ�9�3�v����U�!n�:���i8��
,�Bg�L[��
��Aʹ�ɷi0�qp0�,iXH��r���:e:�z�C�y�ʱ���݋K�s+�$O@�� ��
5Ί�25���Pv����X�.��,���Ur�[���8F0eU���_}��d�gœ5*��V��B�6��[M��V���M����s[,�f�Z��#l�����Ul���»URM�sk�R�$8z�uxd�����L�����E?��)�lP��1��
H�G^��X�q�ho� !O� =R�{.����VU�3=5e����\����X��n��!�i���@��Jd1�. �&ft�cm\n\K�q��sw�������箸��<p��a��ݎ��i��s��V9X,٠��7��~�=�k��۞rq`·c�63 �վwsp��r��?k���Oz�'�6mP�wd$��&�D$p�$�&���w�{�!'�Ix*�7ѳ�s,��\$��HI�zC���,�wɒxsI��0Db�U������ۄ�.�I;���{�	>簾��p8�I��d��k�w�!&�d$�;�i[n� N�u��'�Y�x �hr㺁�S�I�L��vv�<ݟ� ��|�Y'�k�A���VI��u���$>S���|������d�.��zQ�<F6ݒ{�!>]l���],���	&�p�0Dr&l�Մ�OWK$�2v��Ч��BO�����D�d�XY'�w�d�n;�Re�e�u���j�x칷H�Y�4�-m�Y L��g�	\������fHI���(UP�Œy��2�PF�o���	>],�{��9̓h͞�����.S��8�,�{���@|*�\�@h��9!'�}!'�kk�B�QY?��V�o�ɒs2LH��'�h�Q'�k�A���VI�l��B��N�j���L����O�@Ț�v�5��ϙL�ե�\��w(� ,�o@{ݐ��Y$�V�TD� ow��O���ڎF�y��RD��4H�l��nɀ$y�06���i"wS$����PK��z����T/�O�������*��7���Ͼ̒r�.U~�� �Hf�������9��ψ4$jK$���	;]xa$��'{�y#��'$2Gb(�J�h�
Y+9s�~}_|/ޑ���'�$��2N�f��v��	;��!a�z�Ku?�@p6sٗd�ﾸI��yA#�5��2E��;�!Թ�!�K˥�N�2I�Q��L��d��ۄ��,�M�T'Է�p�O4�he@�n�=ZY'�T��+����$���ۣ��O?'�V��(9�ˋ�Pl6]�f�`S��B�A�H.���Cͱ����
v�6NŸ62g�]��N4]���oZZv�6���,��$�lFuٲ�e�H,q���:)��X�m��36�]�I��N�'w��{i>lE����&�r҆R�hCgCmn���\Cod��'�(I�=!�\�ͫD�t�M�l�A̲R.~Ϥ$߽!'�K$����I:���H���	=^,��Oɒs�!&��-�I q�'�$��&I�U�۳����s�yR����'q2O�}Y��	=��	�u��<����H��������on�����$�:�����|��������N��I^넓�HnL�I,���S���8!�~�K�e�'ݢ�o��� ��#�#�#�F쓫��Oz��_w�	<ݐ�� sQ0�p8w��U��ɒs�d$��HN����|KD������d4�q��?HI���=ZY$��2O�}}��.rk��R�u�hFh�&f�\>x���lV����7�x�Y$�V���섞u�Z!�@�OV�I��&��}�۽#�k�,r�8lN�d�󳶿�A_�8+�4W���HI��d���:�(�VO�.�Ϲd���I��dषɒM�C|I.6˲O7d$�qᄓ�L����'���\��2�%�Y���m�#Vݵ5�9G�.ހ�}�����|����'�}!'�a0���$���P6X������	<Z_�4U <��&f٤�\'�\$�2C�(���I�&I���6�E%�ꪡT��p�^��I'�����<S���:�P�O��	;��[RH�1�'��d��G��s�!&�$$�B��'�t��01x<�ɯ���-���K��TPˣ8zRG�$������� h�.ꄝ���p(�VI��6�
H�2BOV�I;���@		�P�	%�۲O��BO�:*�6~��?{�	7H���=Q��n���d�~L���:��섞s��S�!G�Nbd�<�ԓ~��=��]U�?�
�x���P����7̻U։��t�i�6�Y5h$څū=D�l�7dp�)����┴��ջ3@e�u�
\�U�%�x�B���u(s�a�QV;j(%�z�@��]L��ܖ�.ik��@T��0%B�h+�i�1��i2�:+���!��6�.�����B���吓�����BM��O�W�'|�'��u�h�"����m��/�~��?s�<��_�}RH���x|Y$��?%��	<ݐ���ͣ	Ĭ�7��'��	����~��'Ŕ�w���f+$�
�>�$�2BO�I;�ɋ�T=N����Ӛ;]������2�e�Qcm���<�.�%���'۰BO�$��_EiovBI�-��w���We�ɰtD\?ۂ��T�{VI���BM��MH���J��V�9��{}���7d'W�,�86'��������O=�	���'�[�&���*�HܲO7d$�^I;��;͐����x�74a�n �L�-��m�Xh�.�����U��@}�ˉ'�L���j���	=���1��J�'q2Oo�BM�	����_P }Bv�~31������BO9�]��o��6Km��d�~�����|�t
 ��S�{��a˿X�>+ĉ4D8���Lj:1��eF1Y��Zm�R�9�s[E�����nh�M�A.[qj�g\���e��b�b��h1� �ţk��>���֒�A��zs,�")�ѝ⁰E=Q8!�*������ON����M�����O��P;��N�L�)�>�$��vO�K�~W	=XY$���}Ao��������r7d�.�I�AyBO4섛݈�^;�dU�2���̄ĥL�r�'v>���F.�<$���=�d$�����q���d������qm�Ӌ���ߤ'����O��I=�
�F���j�N
����	=XY�*�����2O~�BO�|<`�S���KŒO��&�`��P���7ﯰ���6�p'�I�O�#�O]������`G�o�Ÿ�`а�_R�����ȻU�=v�Fb�Os$$߽!'���;��&�!�$�l�$�tHI��d��)�o�!$��C���'�$��2Ҽ�	��˄��#X�7�� +���2O��BM���H��d����8�dH�\$�vd��?{��$�~K�O�W$�&���Ot��۽�&ڲ�nM����-�T�ѹ��c�F��i6n��2^����hN�q�IN�]q����o;I�$�Ŝ�ۛ�
�����e����i�[�(XM�Hr���g8j�L�m��!��͠9\7�7-����䗟l۱��1�P����Q�$��HI��d��L�y�x�,1�NK$�`/��+��o2BM�HI�zfQ�6I9��o���y�z��H�	}q@�VI�d�������,�s��L>C:I.&ݒy�!'�ŒNu2O����$�W���M�H�F���{c�nɛ+�<l0�YhJ�F���BO��$s�!&�$$�<�y�
qY$�&��V��Tj!@v����ݐ�zBI�ɒg>����!�	=ݐ�~����G�L�oɒf����$�x=�w��wS$�q2z��$�u,c���I���'�L�y�o2BOᢅ1��&@�I$�'M]�ںI��ِx��X�F8p�wS$�{!&�D�Ì���O8_F��r$����	7�IԊXY$�S�U*�d��7Ē�m�'۲z�u|r�;�2gx83�e�#M�[JU)HV��|͸v�ª��D�7���š�F��^ZY$ΦI��	�T���N��,q�P�$�&Iڪ�z��ܻ'��K$���?=6�[I@e˹Ƶ3V������g0&}��	�o�?>}a�_�!&֟ߪ���!%f8I��G��n)d���6���D�&H�*��KZ��c�9+َ��6�����;�32U�h�=����3�l�4��� �1O|M}Wg7+��e�ȩ~�ϐ r��]nk��i���E��O�lfE0��h��.I�I�Ř��Ip&�;���꩘�x�hv��]���("	G{N��������������H�fK��S�bn���
pd�w��F��>A���o�-��Y� 	�9�F��1Ic����:Ϊ��V�g��h5�j�uP%"p�$&�sa�6eC\�������l�m�^�
Nn"�^R�T�MD7k�l����@�G�c��""�.�̣�c=3��s��v�-����;g$��H��9c�s�S[\�S>w��x�ش����V�I$�cŞɆ���P ]�J�1��������/8��̣$)�u����U@!��9�ξ����ޕ�`�d-EK��9�8xV�J�U�p��8|� ;�!'َ�ˇ�T��$sO�#G#u��Ǐ��&n�{�t�o����DT��q�l�
���jq��$�Z�#���! \�sP� _���>� $��A����m��` ����\��@\���I���%���(y���6��I��{�o�"�\&��-� rY5Tw5�=�W����7n�'��ݢ�I�88wPf��	�٦���6�p��[F2с�q`��l�,dSܗT��Ɍ��*���s�p�{��Ba�(I�!� �|�#�� G�$���&���A�n�w�z���{���6ia`����
��b�zl��_N����Y.9c��̿19��U��1��?��mD����_��$��#x� ����8Zp��
����ք��j�H �$�b�������z�<ݐ���#�9,�n������	7��{ޟ��"D��ú����ewu�p��32���xMs�2s�o'��S�J�U`�!��'t���C����!��B��5X��A��?�|���C7v��"C�ݳ@{:����RL�"G#vI�섓�-#�y��y�Լ#u}B"}�p��$��ڠ����M���o��_��H�O~�A�<��C^f���s$��USsu�qj[R9 �x���^�����}�2����d��-�Kwۻ�kZ��tĀE��%E�h��FG�g;�d���-�&�&,��&"�R�M��ZXD��T�T>"���*uE0�E�%qCDRA$�D1��(���6EI�bs���B섒�H�Ƭ����^�l�	�=��!J:�8��/���o`�߿�g�>��*��uY�q�9�i�!.�җ-��V��P8�l��[�����!�ծ��A�WV�d�g;�+=U�(�m�^�5s��-z�]P�[nSf�Sg5��ƛ\[�u��m��M�-%�^��jA&<-�Ңb����UX���� ��K�D�d]�P���댚�7`"Wf'��\���a�ecZv��c�0nT�D�jD��I%�]U�p�N���^�]cղz���/S��� ����wk��;ր��[Rl봼��e���"u0ց�V��� 5��\�F�S���-r�v��u�kp�Z�^i�t��o��#�w(�v�u�o(N��7iJvd�At��m��!�9�6}��\�A+�i�t�a�V�s��U�k=�E�����iM�N�zk�m�����+{a�:���2EX�$Sҫ�Ċ�3�=�kZ�#x��zH��m#�n�8����i`�"��ԕ�[a�4���lHV����1�gt�!��x��]ov�P��mlZ�� �����j���t�2�s�<�Z�d�'&�v��mځ�̍�ݎ�NcmR�?{>��e��.�9�:u��un��p�Np�����vv�������H��D����Pb(�08����t��+��À�+;��{�|�?7�5�țfR�e!f��*1܁�] ��6Z��\3@��6V-�����eq�n�[]pV�y���v
�=�`��Ӟ'3�h�5j:�����/Dܚ`��*O��n����ǵŴ�cw���y�<��4a�o`��ֱ�Ԋ�Z��g?�T��E;IS��������T��9»��e�������@y���_�QB�7��t�,˻ѳϾ�#���ɐw�7�o�(9n̈́ �w}��<�2-�A�(P�6MH－�q�
s�������۲y��޸e�~�ߘpl��Y�m���@�e�2�զ�*��wwB��7#�F���������HI;��$���C^f.�z����3?f�?c@���kU/켒~o\$�߱�G��K�#�9,y���d������s�;�[��8I;����%��  �u�y����l�`���d*��HA����w"w��1��a��j]Lm���H#!aB���i�	��߲@N�|*� ����p��#�P�Hس��p�y2A;���#�����Ed �9�A�T��87ު�T|W܂{d&�>��2�N.A���HI���L�gF���1I�p�u� ����&���=�	篿|ɛ��0��Fk�,�1d���y��V�3%���	>�dn��yӻE8Hr��Ly�8ou�{� �
�c23�}���C�}�>�7gP���o�>�ﾸI�k�{ɓ�0P�T*"�GIJ���Ǫ����sH��#��`��u�*��&믴_��߲��3�Dx�S�oY�6e�P��΁n�.x����������u��0P��O�8g���n�������Y��ξ�D\?��j������W�ĵ�8rVf>�z�y�}{��ޝ�)�C�[���bf:�c��� �U���+ت+m8�I�SiIaK*]���#m�GdV��v���\ܡ�%�]rbf2,Ի6G/\�����"�����p2�iz��-krh��h@H����\�*��^��ۊ���a�ұ�ō��㻻�t�w9�����G��bYq�ų:١h*%��?_�^���~��U��7��n������o�^k��i���n��w�:����N�0���E86��U_:��u�͂�1�G�Q��7X�U�һ����U���Y����s��4-6ЬpkD-H{I,;MB���c��gV� F�_ծ!��[�ôW*���U������U �}���-�K���>���γ<��\�LiIChUUn�}�n���:�>X|�D��󭪪��V�U�z�I�ԅ TD�m��zV쌈%�pT�֋-w1�z�O34
 9�u�U�+IE�!'.��s�b�]su௅P�W���M�W������-������ZE`�  ��P�U=��չ�u����j�?� Wl��������c�� ܐ��su����U��&��u�`փ�R�X�G�7�q���7�[��.��X�Z{�s�f�c2b��Ϊ��Y�m!vqi�8������Y��0�'�ΘP��4�u�|�y�~��ڪxW�S�zJ/!	9u�U���U7X��*D��w�E�%��j�Q�X�!!��"�Q8�sX�Un�*Q�Na/��`�K��x�1VL� +�]'� ܁�_}��z���`�Uw�̢�@��i�U���x��;Ҷc23o��(O;���[������E�u�������]M�n����ଘ�"�e��f5/ Fs�i\����i��Ƴt8�+`����҂�c�1���{j�����'3�p=+f�����6��su��]1]]�˺�V.��F߄[����e]�ٞn7]0���L!)��5#4�f C�>��κ�_���ؑ1����hTG|Usu�����߉E���Y���cuU�1<1�)�D�f�ު��>T�\��K^-C�7U_zǱy�^bd�C"��I�Q)2B+N-��k"�O�������{t�ޠ/w�B�\��-�C��?G�㳊T+��Z��>������s���Lf(5��������1� �z� ���Wα��
 �߾u�#�eW~�1�=�n�7UxUe�_�����B��Ѳ��X�
�2�5$�}T,XE�!';_|��u��Uy�O�E=Q9{u�(ߕs�QԆ;��*���;�
�9�P�����[%�JH��wwww���?$is�h�]�U--��v�7�ǃ���ؘ4��@�Ê�����I�fs+[dn��ַ{���xt��t�����6�4�!"��)Z����H*�a2H}��v�[,6��t��47u�G'ǻ�	,>��}�ir����}\s��y��<���$�Жi4��K4��,��,��,�����AJ��qmm)6ֈ�k2ƖڐP�T?�(������b����C�C@iy� �M�OQ�DN��ft��}�j��\(���?�(�`���Y��8�c�\��E�]f*��(�,}���>���#P&,#3v��Ee��c��c)f6b��<=�L������C0�f*�u�s+̕~#;&2�w��M^c��g�/�������u��?l���pN������~e������H���~c�U{�f ?Vo:}IB=p�<�&�]ע�=tT1�&I�	�VR����_��|��� �s	8��1��W��b�
��-�C�Zt��o5�3啝 �#�UUG۬w�u��6��b�ʒfU^���[坝��������;�'��x��X��E�%����;���8HB�N6�X�b��l�-t�+�#Cm�q�!������9nn�8��z�v�a�k۱*=7K�����y��2mr(�=�n�.J��-P�C7K�����wO����D/����fA%������!�E�$IDI&6�_~c�@^��b�Y��O�������u��W������S��{u����}Ϡ�@p^�.��@d�=k�ߘ� /1�-�BLG%w1�����n���.�S)�L@X!�c5��m�)�=�w�Eȓ&X�@X�X�[@P#�5��+��Q�Y����8��^�%�RP����^��>]�Z��2$�wu�;�� �@svi_�H��}��{�n�����2X�@mB��A���Xg���}Ãe���>g͘W���l].�!�6/�r>r��O���z������@r�kHT�K�@*��cm{��#��I�%{u�u?�EؤAEϾ��i�MOx�̕����3���C�>��w�n�T�5��;�\�cu��o���iW�U�!�8�,��몪�eZ�I��7U_:�������8<s�$ciW��EU }�C��n���P#xz>�B"������T~�W7X�5�G�)#5�c��n�`	��+*� 	e
x*�QQ�'T��5��̢r�2X�U�(NyzƝ5����CCMMtl5�x)].c@BHq�B�(��I���1��[�ߠ,}�����H9c���X�Uy��Ap�
i�k۬p��c�Ƥ�^]D�-X���u�8F�*���\w�$R����OM^`c1U� U�XΓ���jpG5v����L�u�f�ln5� �6��a��a��섺��&IL�I�s���hp<��tH�VS.�Z] ��W�*��X��F� �"�r�h�W�U�n*�mm�����1���׾_��#�J��p���(��c)1r��%F3�I����c�c>Uy���A=RH�\=�n��@\>�Q=���b��_�Gu��,Z;���rB�۬z������\��.D��7Pα��\̚~�������p,�Bͷ^Ɋ�5���k�h*й!X�d����uou���WWQ&D�����2�P�� ����XÝ1#J���z�i
\�cuVY����"),n /�c1U�10`���$�{u��U�u]矟.L]G%��s����hV:�U���)�'��������W�ŋG1���J�c�=>5̶3 &��޲�*���;9s��m��ޯ�  ���M�.��*�F�����3�H1c�$ȓ�����A���ߏӏ�?����b2R-�Mm�V�J�Y��J�o{��Og�W����U�=~�E%��6�
��|��su�U y�����V�g�1ު��Lf >X=��3_z�b��*
!]�
-W{gT�nVe�<�l�(5�>3����^��e�k@M��Ȳ�	uևH���<ڽ��7��� /��f.W��8�t��G�?���W�����i�����"N�b��XÆ�1����1(�C� �u�#����^�����")�>4��3^`c����"�ߟ���h]������!��0'���J�[d�% t�B�Q#s�O�q��yq��i�����B���, �J,�l"%��`���I	V2�H����w����x�9�����$�S
�F$ �6�cW�)!L!F��j����bR�%�(��]�U��"�`�bE`DS �,�
B8eD�j!��YD|J*�ja�J�����)�	��,>�m�V+US��K=�������d�ρ�s;@LD[�O�:ϵ�R����+I�����C��
����a��*e��ǫ����R�'iےZ����KV�fO*]:d���]2B���A��YN	6�c�ֵ�m�;l�H�#i6 �`�9[D�8[r#``��8R�%���;M,��\\JO���r�ogl�@�:Ylv��P#�e��\�Z�oUl"�qF����Xѱ��i��y�N�q�[G\�ez�����AJ ��gf�@�m�ыWA��2]�h��"�AN��@������u*�����f�HV̛.�J�`�k�IEB˭�EX�� ��	�M��]�A�=�[��[$�����Ҳ�
Q;�lk+��&x����7X�e�0��{i҂;�jۗ��c��w� W���Kvú�թ��[Uܠ�U\4.��y�,Ǵ%��gqh\�*����lp�"���s$�;@�b���FG��D�x��'i$:'*j���۶VѪ���l���0�J�:{�x�+;im]N!G�˸*�yv3WiU
Gm@�s+�ɮV�U8]j�?�ZW�����AKR�CBkjQ���6�UJS��>�A��-�;/�n��&]T��w&cDL���E���z�F��`�c��4��v�v.���{]�]��$�'/&��9=-��>zs<mҬ�����sn�k���T�m��`�jc�).4a+�b�pm�5sE��ӺI	̟�Cy����R�@e��-���f\�ZY���Y��J���;�Ϛw��w������y�|9R,}��XÆ�1� x8��!'���M^���5;�fd��Gʟ*��<�}O������w�oH&B$���9�8y��Z�<���X�vXWSZEκǙ����^��ޒV6� 9�=O�m_:������bQ�����U�R PS�@=�gu}@3���oЄ[��j��7U^c��$���@�u��U���M:�x���HT|�uU���U^c�p��C�&Im�N&bLLgUC2�����t�>������]���7Ur�wh�
]n��u��W��8�i�1W�X�P���(PC����nj��eOy$����P����V�C�Ty�u�#|LJ6���U^c����H�e��0@�.���R��.�����H,]6�&NVj��X�Uy�L���E"�nl�(�!����u~� �/�>��guW']n*��.��d$�rWs-�9n��w� �>�=�r{�I!H�.�P�X�Uy���9ؒ0`��XF,�8���Il4���h��n&빌N���0�0��$�v3�Ts�cN�_s�U��BbP��{�����3z��SO�܊�ڴ���C�*�<��0\Й�#����;��9���r�W(Y�`�ۚ����������p�u��s���Y�7�(���C�9�5�;�؝g/=�&Ձh�����	��e:�d�j��g�{E�D�v�t0�jA�4c����c�1�EmE�]OP����#�:��y'���d��tf՚Pm.�#s�|�1=�,�s<���I����ڣҍ^c��9|;��!L��i�Wα���8VaA�װu�uy�~դ�v5-�$ȓ������f�1�z�]h�X��:膄Q�����IDHI�&�{u�����Pgi���e_��Vf���@�`����*����䞧$5��;�:y��8iߊ���Hі;���8j��GRN%w1���9��{��\\6����M��>b�ڃ �#�A�2�IHP��OM_:�b��b��
�9��1ή���!�RK9$��W���[��� !����S�u|#:I�&�#��C�W��b�8(p�D��FE,`8h�9}f*��=wջ���Ԗ��,d1�%p:r�%Il�rK��U�|��P��YЩߊ���Hd���ޗY��� n�մ�P9+��A��*���b��q�F���;�3{9�}�a�4W�P#�ߣ�Y�
�6b���:�f:�U��^�l�j�&n����Q���.��s+J(�>^}N��m��W�o�1@�U���U<�3;�"J}���1U�f*��'�3���H�>�w��u� ��
���H\�9��:�1Q��< 4pw��Ӝ��E��+y�m]���)��x'�U����]�kD%�G6��q!��������M֔Vf����;�q�\؞�:�������ю9�o:�]-c\l��t�丼��eL�'w�:t���̙�&��-�&x�WE���s�L���H�f+��rW7]w��w�UP��uW9ïB2�[���c1U�1vW���������u�5��+�(�&D�� k��b��b O�Βb�������W��b���rH�-����!�T{����S\�)�]��\��<��j���.����!��n��ڞ)O�UB�v����+�o�Z��0�%��0��y��@�W7\�GV�N9�Ͼu�*��뫻��@b�.�_OX�U3z��&#A�	�X۷iF2�1	�9��/��	*	�W�_	�<�,Bq �>Y�Iq7c1|��R� �>#<I�&�w��� 
��m��%$J|�I"f�AkZD�T��m�o;ǆ�C=
GlX@tZ�W`��D:hHБ�}4E�5�Nԃ@�"Z	L"1�(�j�Q�����6ޞz�D�	 �����&؝1���C(�����C����n��"�>� ����'�`iB�)_�%���R�"]fY�)�y�DWa9c1U��f!���^�-5�C�{�X�B��c؂?B_3[��#.	����.��[\'mHK*3P�!��U}���3`���q�]�c�^#�ݜ��(��V'�܁�Ҫ��4-�]�b�.�%�$0}T}��wʽ���X��;u8A�ޒK����P���|�7�γ�>��i6�f��uC�=�ve�P�-�P�0��>�c�U|�3��"�� �,s��
uT�s��W��O����aG+��w�}UU@�u��N��g�(\jX����:���D��bţ��M��w�o�뽾N����|
VQ�#�^��r��V�T�Ȯ;up�	n�!bA�Ȳ��jtX�;	��5A���Ux��q���s���kfl�ՙ�&u��[�(�0r��q�u�FH���qv�i#=\qű!�l�d-�x�j�7A�FU��zI�'��;���6Y�E��X�uV�]D�	<�����x���Q���9j?v��U"����G{���%�fd�]{큂��w�����O+��Kʻҏ{@��,_@T�����l]���ɒ��C�Q�q<��Q���.����^�.o�ԩ����(��D�
 �=�T+uU{��
�����$Qۮ9J��͢u����#sW&U�����{j<� \S]�P�����5˜��0��Q�ht���� �%�u�����-GF�{�®���y�ڎ�@��mG��[֫�ܗ/1���|�|!H_����~��u�֣�Uw�K�3&��u�ڏ{@������%���a��7S&��u�́p��g���Y�$���ڏ��.��S��i"Sy�א�!2e]P/;��Q�A	���mG�iO���U^VQ.�J>�@��,_�!$��h�*��9���#
8(U j��nڏ�P.�׸���A�f�_%Q�L����r�|�뽱�D�J�_�#�e{w7i�E�Z�6�@��9�.%V�I����P.���{�֍v��2fa������CQM��r	����S� 9ʯ{$��3&��mG|�|E���mG�h0��xB^Uބ<�{�}��������7n��!k^�`��;�L�w*�y�ڏ9@��m]@{ړ��_>~78� ����tG�Uq��MΊS���{���86��P.��Q�w`��m����^[2����P��,��c�D�R�"D�7�W�2L̽(��~R��P.���tj���*�/,��j;�뽴OB��.��j�ɓ3�ҏ���$y�,q��߾ډ���(�F,F �=��y�{��y�?z����`K�m�`�ɑ�ZD�j�R�q�K��AC����ky`-X�n�C��2�%�E��i�O=1f��� z�aF������j��7��ѹr��dyzѮ;��YA�5]v�̬�K�?$��o=[F��bX3:�<h�ٖ݋N�%5�b�d����I;���,��Ͼ���M{@��;\=%�fLҏ��.��Q�h]�C^C�	�S/.�.!���s����{��L�fT�VQ.�J=�뜵��u�ڎw�]r�,�x@Nw���P.��Q��|��W��]l&�uk��A]��;[@�Q���1_;�|�v	�<��뽵j�z\�̻�㨧;�N �s�PhB�H)�:��P�EW�{�M�1�@W5cx���7͵2�L�S)��e2�L�{����)��e2�L�S)��e2�L�S)��e2�L�S==����e2�L�S)��e2�L�S)��d�H$�H$�H'9u�d��fLЩ��e2�L�S)��e2�L�S)�s��S)��e3��۾�L�S)��e2�L�S)��e2�L�S)��e2����L�S)��e2�L�S)��e2�L�S)��e2�L����l�S)��e2�L�S)��e2�L�P�iɔ�e2�L���S)��e2�L�S)��e3�q��e2�L�S)��g�+۞�u�n�����e2�L�S)��e2�L�S)��e2�L�S)���t�e2�L�S)��e2�L�S)��e2�L�S)��>����e2�L�S)��e2�L�S)��e2�L�S)�χ�]2�L�S)��e2�L�S)��e2�L�S)��e3Ϸ�}��L�S)��e2�L�S)��e2�L�S)��e3�m�������t�1%���r���u�mJvZ�)m�z�t	ҙL�S)��e2�L�S)��e2�L�S)��3����S)��e2�L�S)��e2�L�S)��e2�L�x��S)��e2�L�S)��e2�L�S)��e2�L�y���S)��bf��"�w��+��%�hE_}�W�oy��e2�L�S)��e2�L�S)������S)��e2�L�^�g&S)��e2�L�S)��e2����L�S)��Nq��e2�L�S)��e2�L�S)��e3�����e2�L�S/N3�)��e2�L�S)��	 �	 �	 ���Uyw�L�4*e2�L�S)��e2�L�S)��e2�L�S)��_on�e2�L�S)��e2�L�S)��e2�L�^x�L�S=}z��e2�L�S)��e2������zg��2�L�S)��2�L�S=�;�S)��d�L�S)��e2�L�)��e2�L�S)�}=]�e2�L�S)��e2L�S)��e2�L�I��bA$\�Wj�v����� �	 �d�L�S)��e2�L�)��e2�L�S)�޽:e2�L�S)��e2L�S)��e2�L�I��e2�����l�S)��2�L�S)��e2�&S)��e2�L�S=��t�e2�L�S)��d�L�S)��e2��ʹ��2�L�S==����e2�L�)��e2�L�S)�e2�L�S)��e2�^�N��u��xe2�L�S)��e2L�S)��e2�L�^.2�L�S=}����e2�&S)��e2�L�S$�e2�L�V=�re2��קL�S)��e2�L�I��e2�L�S)��2�L�S==����e2�&S)���* Y��|�MCp��J�J\�Ҹ��s݆ݲ�kN�Q���9j=�`��]��^��Z��H��mG��\�y[:K˹zQ�h[������u�;�L�˺�^w���R.���H�
ҁ)bt:]��@�f�Ԯ�Q.�4���r�{����Q��?�.�r8��;�u�u�qSJgCX�1i�vt2�;�������]w����O}�\��z]�\�u��Q���o�-G�h^�j\ �=���̲��u�ئ�NP.���;�ֵھ�ɗ�f�{���j=�"�{j:�WN��̙X�;c������P�b&�T�|��i�%>I$��uSQUg�������K��ƣ.�!�"B��q�a(,F� Z��V�$E�� �+A����X�e$^��X��e�Z���eF�3��O�$6i��ܫ�6E��QE�BBZl|&��YrLo�v�������D^}��Cm�����(H��D���k�|\�t&�ך�a�%3IW,�R��8�����s�8�VА��WTv)�����R�L�kf��X&#0l�\�XUZ4�� F�WĶ�2@�N[\[B�������������v٤�	$g�� Yzֶ��6���8Gu%��^	��ӌ$n��m�݈eM���B��Rڤ�9w[R:l�\P�f�Wiaʲ�.eQ�Gl9c���I+�A��a��-�Ue�t.�?E��c��m�*'��WlyCˤ�ۅ܂b�4�[e[l�lݱ�v�v�;n3r�@7V�t����)�iIn���ɃR�l�a��\�#2��0�P�_!^y�ĂBcwh�-[���E`U:��n��m��ɐ��w0la(�����6����+�ko��a��-�v�9�"�h�y9��U,[^VV�6,�������S�/l��1Tn�{r�ʆt:H3b�G��I�mupj�r
�J릭�/n���G���m<컗�6�J6���Ui�M	p��zwV�u�T�UgS��^UP�65���Y웠umѣjU䙖��@0���=P-| ]l@�D b��*�_�84� |A�#�x�w����LGU�a6���;[�K'70�ܷKc-�/Y�P��>
ض��g�>6M�9C�5�ͮw�����7UǔB���xn���(�6Cl�-z�6��0nV�Cp��u���7���Ys��I>BW��m�fॖ�J���/
GB�Q��0/(��G�h7�@���P/y��Ü�ɕu@��mG����Z�{J~���|���v��.�J;��]�T+uU3P��Z���!!�
��t�r��^�h��O`.l���u��/3J>�H?���}�(����mN���ݓ7A�h;0��b�ɴ/,lju�qY�.��;�|���s�������o����J=��mT]a�9Z���s��=H��t���fe@_{�� ����{; �	�<��%�a����s|�'b'�_y��r�2�d�]���r�}���{�n]�2�噙(��k���l)p�P!V�Ԭ�(�y���^o�j ����7ﶣ�����Y32���Q�(=��{;͞�uW^\3Y�mG���<��A��"!@:KG'����rO}.r�-��]���r�}���u���\���ҏg`=6��^Z���.{��5��n���г\SXJǮ7Z86��]�Z�ZI����P.w�����<��%�a����s|���^��!�Bdʺ�]��������2	��.y��U��%�hC�!����-G�hr(�>p�.��Q����/��Y�LȁQN�����U{��W�*�ߎ8QR2���	11�3�.&�k�՘��G���X�\�(����v!'`/w�Q�wr��^]�X.��� ��r�U��@m����j�K;�=;��F�v���$���k��^c��܂Kp��XÆ����+�N���x��\��mZ�;h� Vޙ�[�3u�i,�V�#ge��c=mA�Y��1��h����6���J�񗛀Hm�f�nb8y5VG=���4(���)����/��q2�xg�0[tn��g^�����?((�v;HԼ���&a�B��X͸ģiU������f*~��u��-�p����y@�Uy�ne����ߘ�UO�c.��i��1����w�a�> P�;�c�Gv�q�su���e�����>{�U����K"�f�qsք�@X��mz�N�5�u��uy�]����$��`}�T4`X ^qV�	:j�˃ApH$���s�h
(��[�(��LQ��u��5��3?X���`�/	8h��}cuT�b^�X.D�(���m�Af��iO3�����$���4�Ϊ{���t��M6�Q�cuT�XÆ����9���n:|̂�v�\6��)�a�k�=�9�v��d��Kt�9�3L�.����!2DGN,�9�W�����LF0Zj"L	^4$����Q�.<�nB��A"�����0�s_�Βb�����t��c����+��O�r��F������Aw�&|�ݐ��}UG���yW�紐*�����\�N��yQ9cuT�XÆ��ŏc�8�rBKl	��Xˉ��e��S�r7s1���c���$�9c�:�b����z�F��2EnjbuUᩖ�0�K��:XÄm w��F���%�k.�Ɍf*�S��}$��~�QHn��Qw8.�ܷA�6�5Ԧ���]m�����Q�V���ݱ=s�.zƱ9�i'��r�����/]ѷ
G+�J2��#���B,3�W=�L����g�y��;n0�ؙ�+0"�,Sp�2��a�<�v������Y�%��WI a�:>?�:��/��7X��/��Y
8�}���T�XÆ������1���1��fu��}���m�>��y�ǏMn��P�u9�I�G r���\�X�T��Vx��)d�`)0CHFӸ��:�%�&�suحPk3�U<�Tp�79Ѡ�ā���ЖYI��M$�H� w�y]��u��	�7���iN wX���z�b�X���a�,a�]�nt�*��Na/��v����;�Ou�8k�&�Z~i$��D��$%�'8��]p쓱���eNoCpn�"{�C�Ά.��dF��W��zQ�w����1'ڎ@�5���[��kB�{UW�~�u�q%�,�e�h�$���T���!�J�@�J()	����_ɫ>�.Q���J�]���z��Z�C�JA򍜤`������"`Kӻp�fy�5�7�Ǯ�"Y�h���Q7��"����#�W�}��< 6.�2@����[>��8�↕E����N��B�o~UL�.���T�H��S[�Ǉ�=��V-5/t���9cuS�X�p�gX��b�eN��89�T���	�Ιm�r(��A���=5�ݪ�7U^pj�p��rƝ(���f!ff?��<�-/�j��k~���UO�c��w�m��nX��N{�;��S�h���O�b�T4� +~����sC1�Ò��c�@fu��Z4�׋����*l�5 *�tp��NTr��@s��7V�%��ޔƂ��C �Ǵ��M�LqsI.	��u;�	�gX�3���iU�?y��g1W��b~p�ۖ=���z�b���� t����\?�	`"��U��I�3��muSֶ�g�2.S�[�"BP#2n�����p'��+�)��͸����Ǩ[M��Fb��ic6V:�����Ѣ�ϫ=�=����=�HPI^���M��$�x+� ;]�R�q�Ԑ�X?�-�'[vݸe9.|�d�%p���������UO�� �8�g��3>��fu�v�`f7�����}���N�yRH������Uỹ�+�PC$F�=�{�u���8k��~�\7:Lc��uM��yq�e\�U1f|�>^޽��v=�mא�	��˪k7��@"~��΁~8ke��O,j}p�ۖ0��f*��L�Z_z�n�nk�u{�a�Nǆ6��G%��Us�a�Y|�>���드d�m����䧧��98.��×L�������q��,�*�syR	�<p�y�3L� $jJ��Vd��Q|���+�� P4�+����z:Qv����	c��W�1������Q΂�*�c(  ���u��[w��Ȓ%Ȓ&�]���2�*�E �*�i��rǎ�:�b����%����Bݴ���;�Su�4�`�������w�>:k{�]��ȎBܕ���ң����l��z)�����Uzd���4�k�(w�n���z�z��bF�p�	ȸ�{\g�՝(�A�aL@T�H�nk�=U7v��t��.��"2X�U;�0��=s�A��]�c��x >�|��*{c���B7,g��^�n���L�Y_�v���n�޺��p�B�����Tv�4̍�P&�fK ���1�Nί������v�A�]vE��.�k>��g. ��x0l�]f��̲����i\ܒ�u�����e�P��dκ���t�ܦ��%Li�[n��.�fT1�y�t�3���=SҔ���K	n��\4���:�5��]�=(��߁��ޱ��5��d�9���lIW��R�α��x��rI*#c�w�<���+�2Dk��;�S1�8jz� �Ic1a�1���x�6�e���i%�u���5it�j�Dh8!���~>>��?U/UL��עD��{�N�P �*���>���O�%�O�h&��c�U7XÅy	��2��B䱘�s�x�αw���&�J��A΅�*�c���7{�T����t�c�\ڸ.ք�` -EQ�ȒI*.�{�7V� 7X�
Ѡ�	��7��/��1��=k�2ي�b�Μ���V��)�����C�F$��c�&��p�*�����!2��y�0b��X��6�E��pq�������꧰�D���g�r��f�ߘ��{����NE%��W:�@,�%�8$I�u���:�d�Y����IVL����|���`٢IH���@C��pw�| *C$@��1k��y�t��<gE��)
L����^ջ.����Z��f*��p��(!��Xy[�A�6���� >>5��n�ycSo��$y�N�:�g^c�%�^�l �#H9�v�؈��bug���A�;�:�fv�����ۮ_�~?�R��Ԫ�Xl�7��l���_�·1�}ۛ0�	��ȿ�5[���
 ��Q�v��Ì��L�-��\��ҧ�THE@�
fwq�Ǣq�f6F���7�j���	�"����`�&ʹXg���6n�K6ص��屳)�@��Α�ڳd���k0�"�GP@AB����D��AB�(��(���G���N���-��1�b��<����7�5��_�Q��-��"�@����Q�O� R*���C��y���
_���1�`
urg��Q�����������SgL���(�ЧG��Q���̓�����Q�M����c`��'��-����s5�������O������e�g3�x���p1����]�o{�l}��i�
��6|����q�_z'�ǜq��}��~g�ul��<������y��c�s���
����'�l��ݗ!�������<�j RADFEAQ�]��ق#B��l�X�Zmb�d�kQ4��em2k6���65��bd6-�dɶ���f�A�[hY�L�Vڛjb�| �f��m���B�����l���0�������?�����UQ���/�<>-��_��o��3M��|^���>��v~��x��/�}��~���1���y�gy��x��S�����>[��q�x�}/����;�����o��W�~���>��?_f>^�lG�W�?�?����O�����w�b��H�֨G�����~��f�R�e�+�p|�����}��h���?�?)Q@�?���K�|���{�����F�ޅ�
���!P(�` ����C��bp�������!�xl���|����1������ߣ�|p3����ާ���󿃟Fu���GO������?[�,?�so������?6��������6}.�6>^�};�G������>?�6|��>	٣��q�[�u{}�����ӡ��'I�y�`��G?����ӟ�G�~rW���GN~��N@�'�|(0t��h��_�~߇��
 �������<��AC�k�{�>�ѻ8��>��oy��<zGm��=�Z?�!;~����w$S�	�,��