BZh91AY&SYV�n��v߀pp��b� ����ay�
(  �P"$ +�JU 
)J $�EH"P(�@HP�� 
� 
QI �*� P��E*EB����H($��%B	(   J�R* U*J���T�PH8    m P     � S��}{�c\m:Ӎ����d� ۥ-ۯ'�f}9\�R���X�:���!T
���
�5B� h�P�mJU1iAJ�����U)� l*�e�R��hU7YХ1 TRX      : � �V[���W�W��yۭ^wx�^� eUb���u�z���yޮ���g�(ž1��1�4	%M�yi{��z�o� x�ng�ʹ��C�e�9�\�ǀ �yT�S!�&.�x��= ��@  @
��
��ݹ���ӓ+�rt, 3�91��Mw������U�>�K�i�'��=��� o^3K��^�yϠ��S-��ݷ�׬��n-%�� �y�V.�{۫�L\��_o  � �       �
G�	������5& � ���y}�}�i��Ǣ�o��'��W�/  m94rrq��8=2��g&��u�����Op �:��޽m^,�e�ӧ.B��@ ��   �@ s��=�7N�����y4����>��w�%95K��y��=����\ `w}o�!��T ��.���p�7H�g�׽�=}7�;vyo�X nR���;�z�y����ם}��(      :����J�(�zM�d0��iM��zL��P �#  '�UR��C �	��bL"{J���A� @ ����M�T�Q� d�h B��*Q�Bz&�=5�4<�=S�O���������w_������G^����UW����EUv*����UU��*��/�iU���AU]_����*����H ����9M/����������$�0d3��qw躉���nMzk�Ts	���#}��J��x�	�4�0�GI��тw��8�\�q[���ڴZ�LX�$��M$�ʅ�٥�u.�uL��|�k�=ϯ~_&F��g��Tp	�0�έg��)��^�����TD[�]v�)�wQ��?�x�*�3̖�k�|$�*�6.$�Ċ&��U����g����p/>ߗQ�s�y��#;7A�;��o���~y��8�i��|���vK�%���D��9����5�&4�PX҉57��Q�P��	�t�U\�������A�;��ܞy�!=j+��L]1��{���&����/Z�������OZ��~�|��!Q:��Z,L\�ɝZ&�i,g_=d/������.'ϕ-�>j/�֜�P�h�h�E�.��1��Q'�6���qD�`�'��5�|��K���q��P�%V�xi##�bfvv��z�Ja�ۉ��ME78\I�q����z��x�	��������oT\[=�y&K��y<�f�ű��T�ո�%H��
�����n�uI*9����G_~��g>�Վ�NE�4�B�0@��Ϊ)cg~}�"��׊��(�q&�i3hM�b�@����Ý�������4�0��q÷�s��'S��uu���VC�u��T�T>��=�g���_(/*�����/n��'�Z�u�[ą�Y���ߓ}���.�C�ITST�y�s��ŌX����uǹe�"}�>λ�z��۱܆S^�0FXK��(%R��B$lu&��d�bx`���<w�(,A�V����#ƅ�����i*��Z�~��7���t�}˓9~����ۺ���^}Dr���,�X���B����DM�5�7����|�Gj�����?���ϻUj���`#����I�0rl��p�٘z�c�#r�6̜5�v`�u<$�a��s��WW�i-��)��^nt\�j�An�,��hɑ���\�`����φ$�a���E���D"U-w=��]�b�l�wN�BE�xxGd�I�0bԘ�`f"jBt�0��,�xf���#R��c����>�c���yh�/;���&0��)�.����:�_r��bW��1��K�����ϖp�f1b�̂쒬n�G�_%9s��dE��Q�K��䲓H�1.�D�r50cL�y�Km#I��Z�C���*�[����>��u+��5�g0u4��㒶��w��`��Dҙ`�Ȉؐ�)e\"�qwG>M'[�e��qwd��j������^m�Nb;�1���w�UO���y�8F�.���2�v��Ep�Ȍ_F�T�Ljb��s9��'[���{\���onD����<�1���1Ņ�i�<{c�`�RF@kFlpѪ�P��	d���4R�:3,1�l݆��i%31�l�R��Z�/"��m�r���JArq�om�5Q7�ɓ>$h�$�g����Xc����]�B]1TQ&�N
�Pñ]�����P�r���&�V��w��>����#��C���L2ṉjTj*��B�5;���^�����w�04c���	OTs#��|��1�ug8�Xg��J��H�����$�g�OMZ��b�+�S��1!�4��I�c��U���ɿ��&�G�QA|�LX�%>��%��^��T�ٸ�#1��A��^�ٽ\�4j�����~_G�]��1M��Y�2	&�����d���p(�~|'}=��|�4x��#�kcԨ�4w�p��JJ��57,�0����4�Md����A��淎e˔ΡL�Ġ�i�`Nٸ<�s�����(p�Ǖ)�H\��ժi�b�SlQ_gE��3uǀ�g)�����X���;�V��7eՔ�Oǉ�d�}>Xj]��X6�XbpN*P�B��{��nV��z����s�Y��V����w��s�D�0b�4�Ĥ�
bj�5ߗ5k�q�B�b@�h2}�Rs�V*��pH|#�b�'�4]�9$�F��p�����MDƞcS���=�>^���1.�PO&((��	.��\T�̨bxbbL���%�W+|IC����s}�z��z��0u	c���&0Ǵ�nL1!3~L����x���R0�x �!��D�o�:�QT��#C�	�Th���ԙ�5ì[yBT�&,�ȥ[���j^|�T��]/8����%�C�°��y�5U����Q��[�Bg0x�8̘%M1Wv}�|��#��j�>���'W>]K�q�S�}�ԎԘ��s��6��A��6�h0d�"���c[�!5T!&1AA S��4��'>�'9�<�E�r��'g�*%1XҘ�N+�ǣ��g�Nx���y�y��%|o�8��ƶ��ظ�H�͊4�%~$\\��B��j:�7œ��>�|V�D<�#Z�I�1�u[�.�����6�*sGP���GF��S��b0̡�NG��<s�,���3D���I�<[��������/.��>��To���,�E�\ظ���{ ���Y���Q���d�ݳD5���6�#��Ml��Y4�I�wc��{�غ�٢z���ݻ�y���+�5Ns~.�$=���U9bn�R4�g���9Sz��z���ĉ���I��P�Џ4D����Q�ו2����7Nn��y��q���o3����q�Ԛ^���P��rb�D����-2n�%��։�|�m׼�A��q�ƺ/�$1}�'$��O0�&e��7�f1b^�ָ�}wW���_�7�����s˹�q�%�.
(+�1'���b��k��S�+�59�y��x�+� (v/���qv�����U9�0�����R���D�-�[�1<������'�U����P֦�@����3��7y�d%�7��VA�t=\�-���k�����~Ŧ%�>G�u�a��i&d˛Nh����e]q
XȪ��IDD���^�!�ֽ����o6�G+P��h�RD�W�|��#9R��9���mr*%ŕ�f�^=�r�'m�V��uc<������9�r�N�}8��:�2o��&���z�L�.�4kx�u`삈����c�bs04og|�q ���!�W�]F������w�����//���y)�EN�3����Z�ظy=�[��]��p����v	�����w>���z��k��Ŝ��ɟ.�<�W[P�Q#����q`ꪏ�j
���:5kw���:�I+��u>I��dDٙFg�-w����\�K����:��'!��Θ�z��1&&�X�H/��M��R<ɍ���I�֢c����w��o':����9^�,qh
���N6�����F;��.!�}`�Qm*�\]��FU)x�gSj�����PL�����|��t8��s�.�����hg��᳸��ER�M$�ǎ�ϱr���R%GU%�P� ]�A��Gٮ�%J����9��a��p���8k�P�M�u	ܻ5�k��))�Ȍ���En1���W���oMέ;ًw�QcI���>����4�ʝ��S	�a�]߰�ĉ���� Q�����12fc�MBu�����a�9�
4�&l�I��۠�-dDF�^cô��l�Z��e�e��i���`�Ԫ��j*+�.CS������C��Ԅ`�㘆�3:cA�^#F%�=ؾ{��p�D��57��HV�������q�x�m>I�Ύ	1!��T>�����/�u��#����t[�%W�h/��0�i��QjHÒ"���^|��ɪe��LjT���k��~��w�\Z�W����\ݰFU��N����q���K��)rC5������a͒j�I9�����x/����ө	Z������`��QD��3ړ���|҅�O���]y��Y�<4�L� d� GܪdG��8���O��R��4�%t~�׿%�$ӏ%��=�V��p�q�\i��w 5i��FV�!(�A0O8�������o<�9��%ko��+P�j�00���/ �bK�L�����5}�_z��ut\��bb��8&A"6����_#4A�hƐ���DPX��}�߽��-�x"Y�D����X�lRb8LH�U��
�h�m2����ta���_��{ۓV5Bv��~I3.m�f<F=&�6�K,z�b��#d1�h�^πP��l�����.MW�WԛY1T'���w��^M|��l�۲4.f�y;�غ�{�x���+ߗ��L�2$�F51@MBu�%$c�gX&f�����p��1��J�	"2%MInb_'ڗRi��1C���~\�1���������#�r��M[;ƭ�hڔs�V���|��S
�������t���o}�.���"1��:�w*CD��ĵ�����Μ�H���"BiF��}{��w���u*��LB�J�h4WK�k�͘a��a��lP�'�����	�)h�݈1vr��T'��S�C�M0W�s���R1���}�i���D%�ɂP�4�C�w˦>[��V��^'}�'oZ��w��nQTruν�]���N��ߠ�|=��p����<�|5�]���1j�. �/��븋��kS�v��d��~N>sZ�6��!ʍW�>[V�>ϊ��}�����7��K�ky�(0��}���E�#$�}��1V��+k�B�d:�\1��Q��b�*�S�@�d�����x����9���������W�q.]�W3���Tm��Mּ��r>�#>s� {�|�9���v�c�H-��qUZ6��9{y�^��N9z��I>CE�Emt��d����p�a��r��57�?���4�|��>�c�t�S�R3��;w�_f-�I��#N�Ԇd��E�Z�9��oT籩�V�ق|ukcr&T��WE�K��aI4����_��ߣ�B{���X�j$))Ǡ�	k �KvWG�α�lO�P�~Cݔ��Nnj|�O�[�g��)h�s0ǘ�J������9�z���ǋR�n��&`�=�T�qUV�[�1�w�A�n50pķ�Y�d!��>E�s�������N��� ��j�(-�~�ߛ�3�}��R���<J�.�3��z�.Ƅ�%	�x%,@�C1�S��co~>�d�%�e_q5Ϲ�d�>�/	�V���-x��g�w�ًEs��
(�\"B�s�/�^s��ǒ"͆9*L����9ϥcFϜgu�M(@<vo~>{���r1-�3]��̝�w`DN�Q�kT��{��/(4�/4M�}��[�b�(�t���
�w��m�5����߾յoc_j�Ɛ\�s���!������X�	���8�y:vF�4�h�K�ᨷ1=�7L����h��˜>�19�u�������.4��U�����[��B�4X�bJ���*�W�
��_.�Ց��]��w�+�Ι�ߝ��)߶,{�>��������/�"���[5A��Q����*��Z�?������v��}�������\�Q5�6�fͰVkc�N�4��#Xϖ��λ>D��n沢�_�f�r_�}�����b{E��wxq���r�F����������]����A���m ?�> M&    $   :Ym� HA��m�  �l[@ �o�_� R�  ]e� 7l�     ���t� l� 8�l@-�h          � �> �e*@   5ڬV5#,�������kH�iʱUG�����.�4qY���e>.eM���W��@�����V�i@�\LKUʴ�z�5�*�I����� kZt�7HMc
�ʭUT�+̫N�I��US�u�7G�lr6��ݺ����c���KR�ʎ|f��T8�k�'�ZV�vx@�jꪥZU�qA�Y%�5I@���R[x�U�5J��*��H0&a�i��-=�h$;m�K$�m�m[���@ m��k��4����A��UW�����[v�  8     kͤ9��	Yvyظ�*�v^�-U� Ҏ����(�@��x86j��8 �Y)�Ce��5�����c`⪩���m��N����P�羶Y���PlU;r��'d� �ZERP��;ڮ�cs�/��*�Q��ݬ���������ky�I�%<�,��ܐ��;۶���N�x�W�T������D)�`�Td�cN��2]Z�CnA���@m[ ��d�n�&p��#Z�A�Ŵ!l���榪j���;�vz�-�6��^ݹv$� �j�Z�VrӺ�U���4�T��MٜP Җ� Ҡl���n�;h�UZ�@W�(�sM���UWf�'KxmJ.�U	�P����v�m���ۯd� M��;u��J�'+	�m�#u�U[up:�6�m�k�0���$�m��Ē �]�Λt�d5+iN���Ol���xjgKݍȚ�B�t����<���p2�4�]o,�g�Y�7X�<^��67g�v�n4�m�wõ�HI�0jv�p�UY$��˷u��k�v��k�{V3"�c7f��.��`g��\�c`a�.�����=l�O��|m�E.�qx�:r`��Yơ���F4�:����4��r޹	�'TQ���m�Ӫ�sޡ�냶��Uj�l�5J�\��K�gv�F��U֬�,A�Z���uJ� �tZ	6촵�Ra��⪀�DC��q;J�Nܚnףm� *�1q�@US����UGZ	�-��U�`��t�p���l96��p�6�$��en2����M��

y�UWf�V�d�6��7N�F   m�Ӛ(ڪU��H��\�ͥ���[j@V�
J�R�q/�}��U;�*�H6�C�-��@�x
�YwEe68���J�j���`U54s�C}�ϛ��  �+m��n��J�@m�店��qm8[��-l�I��I�"۶�nA��n�	��HJ�UK|}�I��~���ZL]u��i�ڦ� �>�Z����@�m�\�� 6m�5��JiW���ګ��U+l���JQ͖�zM.�8ץ06��7jQŴ   v�C�-4�ź��` ��M�8cH Y^�@��m���m ���v�mX֎/.�`�FV�R��� ����M`N`�m��-�e�ɰ� H 
�.6e��bN�y�c�۝�(
T�;(�EĀ���M-�hH�I6$)[l m�@  ��8A��u���������z��iضP*���J��k���n8	�Y[kn ����Pq��]�
��m�Nw.y�lm�8]s�:p���jeZx��+�uAm�%V�5H��Ʉ��!{R���/-�H4IGkgmt��� k6fCpt��G�P�[����gA\���v-
:v裓L�6�np]5u]mt�6�&h�*�$�H�[T�S���2��IR�KƇ�����7J���ڝR\.6 �Jj,��A.��pZ�Ӱ�:�U�aV�8U|�
����>�( ��ov$x[E�%8��BVWe��mF���0�Ҝ[;mGQe�H��ڄ�9�QnG �нF�.:yR�3MYF����8��k̩��N	2	�DbD��K��@.���q��yVӻ9j����q�#SU�q6��C0�6wkoi@[D�-�rś#�!��n�p��I�c�e1����Q�P��A�6���k��e��H�`v�*<�"��JW]�f:^SV�ppG���kR�l�]Cr�`�p�A��uUJm�cmĳ٥7a��P�[S,^rq ��'G-�$��D�q�>�'ŷ�kj5�`��M`*����\T�9�I='L�56� m�5���#m�Y!��E9v]@\�}8^�FەŦ��K-	�-�Z'Ѯ���2�m� qk�h�U���pW@UUUT���1l/1��,[j�� k5��9'�!�@��]��ɕ��[d�gd^�@cE@�%M�sd['GN�[ˢ�۬�v��/n�m�hi�m�e�KJ��m,9�U�n��h
�ص5kl �b��Vr��ln�*�ڂBڥUؖ��@�����^Z�m�KG*�
�<���-�H^( �n��k=+B�G���u���t��&U��29
[c!�n��v��;�3�$9�h�'mp�$+���y�k	&�u���=>#�:%��\�J����J�U-���n[U+@�gY3��v�T=��.)B�\vݺ��2�[*�U�8�:4g�.��,�5O1�L�حږ�zDu�٭�5*�T&��бmr9G�Α|!�f]�uܓ�Lm�w�)�{�i� w��&:1��&�]s�C�:ٱ���vy��'!�p��{n�L|�5UUJ�0��k�U�������[yp�*���V�Y��[���$�nc:
�����\��Ɵ[��m�����O�Q�+kT�����'I��vR��I�9-�WH5���t-�k6l۰Ѷ�� 6�Y��m��J���COi�͞lY�%j����l��.K�s&c������`jꪕq�T&˰|T�;�^��t*.��4uX�-T�v�6�n�N4aU
L�:�Xy���]Mv�O*R�Vv�ccs���"v/;`�풇C�`brkq����A�dDvI�n���ts�q�H���Y"��B�ZW����INY���v�y8v�YĄ�V.Ênl�L\�[x{R�tζ���蓣D�a#�v�ΪGV�MkGROg�\"��.�k�ڴJ 	��.��u���P�����[\���.�:���t�V�Y-�l�ۃBml�U)l�B����N�P�aE��W�`�k^��F���0����%V��([On[e��jaz�pݡ�[�EP�{VB9��r� �R��3���8uPP;I�΍rd����T��rMJ�`lĝX�. ��uBD�UGS��J�#۰۰33�)�[@�뭭�l@�A���T�Uj�
���[UN�m�qt������vk����V�Q�n�g8ۋvʂ q�ݭ��l�l(u-�5m�n�TO 3��o5�3p<6���]�6�� ���]oP����mjg�n���ڤ�T�
�<������9Ij^������(�*�֎{��Pe1�@�Skkm�C�Y�)�v�4Ԇ0�\��sƵ��dٖXV'�e���=�kq��aݶƙWd:��D�	onВ�\�5,����g�n�cxn��R�>n�[6�n��ƍ�-W#��U�^�Ex��ҋ�tP�ӥ��B��U���WV�m���/$i�`t�-�2�E���H�N6m�F�'Ya�zАU�*Ү�UA�R�Zl-�Ƴ]�֍�y5��U;�����^�]�ؙ&��-(/k�:tuvml!��Rt���͜\����j��YB��f� t5��Rݭ�ni�@V�J���H��lu�����5�{���':�e��v�3��0����+h�����Q��خ����c� uV��0�t � l6� ݶ�m���;"�Zm��$�U�b�ۑ�Ãm����*�yi&s7f�]#��eC /s��}1�JKU@M�q��ћs�LUۡokzM�kn'Zaa�'G��UYP=U���Z��4Pۮ�	�	��۶���iK:T�d9:o+�/[  H$�#$l��b@:s���lgMUK��ɶ�v�Z���Cc��:�����%J�`��.��t��3�a3L* ;U�UUI�mn�  p�@�U���6�T���I�B]����w�|�p/Z���Ce�5��e�V��Sqv���d})y灴�+��v��, �@Ucc[u��5J����8m���%�:��-��-�&�,h8�7/v� t�ճ�l��V�:�'D�u���+j2.S�Z=�Z�*U���e��$!$�vu�oU�[�L$,�27l�:E:�RV1U��Ի8��	2f�)�-��`�ĦX-Y�����꧕4���`���m[�A� � X<�[R�V�W:L=0�n)�*ۤ�Ғ�YM����( v��4Ʊ��c@�;,м��G���U�y4Iז�h����6��-�ci�Z��L��f��������*{N�:f�T
��;��`*��*�tU� �ʋ@;s���]�G 5��@y��!�n��.j�Z�)	U�tٕ� N�Ts�F�eT�ev����pU]P<���K�ɹ-iC�K�6�	 In�,�	 *��TbW��=�uUUUz�Ф��qeiUWn�6��)Y"nF�cL�	��d7���Y�\���|�'��f���  �̦�[@   :����e�6�Mv�oq�DU�_��AU�9�?��������������ڋ�(���
8���)#�e)=M����"��ؿ�@)����������@�s;8B� �D{O��D�G�N����-�D�� >�* ]P�.�}G�D�ۉ��t ��:d $�v���8��(w�z�9�@�	$�v"���pTC�^���xu牱�B�"�*��]({� ���_W�㇠���� hyЫ��;�OECH)��G���N �(�	����ŀ�$!���B�2��zGBx^*�� �����@<LH�v"�(���N�A�A;T<�@|�U=@�$�S	�դz D@q;Q��D�<��pE:��hi���P�t���@���$�44��'��xh�,I"d��"��$�b�,Xě#&� �(�����2T)�u�"iP҂���!���6� b` �t"' {	D��AU_�������>���o_�G��BB�.B�L!�!��B�$T �D�T�#D.����& � cJ�d�4) 1@3�� b��� J�`��B!�J���V���W�� #�!�UU@��fٴ�Ih� �Zٖ��J��5���&�V�Au�M�^j8#A*�^K8G��%gcv��b#G\ӂ�ݺE�'\��x�<֔��ŭ�U�I�U��W����g@;$�ѱ��yS:����4�#�S��j7UY!�!'J�cdg�a�T��/[�ˎ�ݺl6XN�h�v��yKH������Q5��-eH��u�M�kmtq���:�`ur����U�e�R�>;Y�66SJ�xx���h�+D�jH��`(��؎��Mgj�LwK�&��k6ݩ�n�8�WC�=���[��x'��C%%��%��*�t�ҩ٧n�7�����xӂ"�wj��LXzx9M�7 �q�jI�m�����Rjɴ�g]gd#8�w&��Վ&ݑ"ی��;7� #��CM��<٠�{��<"ԭ"�]�9b]�v�h;p힞���'=ּC��q�\s�#���j��L�<\��K���e�[A�.�tC�4p<<[s�-���23�ø�Q��tgX����>n�Rr�t��۔"�y��:���gvFz|ӹ�����cob{[�<Wn���]!�����Q��m����"�璕@℮I; 0�롡�"gq��[��x�e�k����q��x���U͛�[�W�v��nR�Ҿ�g��%{>�p<�mE& �jb�����ΩxL��r=v�9���P��;F���F�J�]X�7!��ƢvJ��+���,P)�ϧ�;[8��=V��@{-Jk�9�M��+�L��m�lt���{m��e��l8T4\i*z�u=�#"gv^.��E��ĺ8ӎ%�njp�����nZ�q�f�vYyun&%w-ۡ��0<�q�Y�NOi�{`Dݹ��5�h0�یi7h��=s��1�l�fv�Q�Vv�:����m���b�*s��=x�G��9`AM:�Ƞ���96�,m`����u���T2m����4��h���z��*��Go-�5����oZÚ�zDD�T�����v�����	���x�z�z ��vhA8���pT0��k?y���Ef�9�5絴�n9�������9��.y���`��;p�8�2s�C�ݥ��M�h���lsqF�t� �=�k�6co]v��Ō�qx�5�n랜7\&��C��w9�՗���������ˋ�Hl&tOm��x�3�v�!ƺ��}<���J{v78�k��3�Mȅ[��jތ�Î�����{;����:��]��PP⩥l���j�
�9��2��P��|'� ;���._s�8�
�w<��5�;���{Θ�{+ ��� Wz�].�Z��V�����+ ���{�������q������@�B�7-Z{�V�����׀{����p&!����� �s� �^��=�{V�߻�Z�E�D�M�	P���.3��ٙJ����T�'
��j=����R{h���VU�
6�]�u�]oS��-]�8��7�sr^]h�e坲Mh$��=��+ �s� ��r�;�o�e1�걶YV�߻�[s>��/p�1��!�=e�}oەy�����+ ��^+�էM����Ӭܻ� ��r�=��X��e`{���2�)Ҧ4� ��r�=���{�h�.�jx�A�m��4w�+ ���ܽ׀m��`}}ԩ��aj��T�p*�VD�z� ��sCr��bN)���gt���.�@�������h~女��Z��p&1~t�v�շX_��m��`��ՠw��V���l�b��s��nc�Ev٠|�{��=�}�O&��Y�y���̑#KTRLL2�H�$�>��V���}4�$1ȣ&��ݕ�o��X_�� ���h�ѿlC0d���ʴw�ՠy������@���� \y�wȮ+�]����amN4�c2/C���t���(<�%�g���N�N��U	�����?���߽� ﻲ��ݕ�{�w}|�&�L������o�Y�������������ޣ�J���ݶ�m�k �)P����\J!�c��{hQ�w�-R)rX��@����Ͻ��:���\��EfǠT:^#׼�ڴ�x%�U�v��Ͻ��8�女��Z>�h�c��q�5�$�=�r�����l�C�{\qӳp�x�E$ȏ|�W�qÄz1�|7������`�vV���R�m�����i+p"�	,�=���@�{�Z�{�q�ޚ:to�xI\M�U�w�����m�r�;����{���M���wwi��߫��}/ �� ������h�6��j%e��bq;�6��`����;�e`���~�6�;�a��������sU�&綍&2F����5��u�<Ȅk�v����	uT����7ovkg��Y�b�����x��
��Զ��q�qK�����1vnd˹�-��w�'3�����z۞/�7\pIӴ��jfn��6y��\��z��BۘS�M���7U;k^�ev��H���Ӵm��r�&�+����߯{�w��~��^���	JY��|oWĊ�uYz�n��knob�g�t�8��eKz9zk�A�U<7m�zL���e`{����X��;쮑������ڴ�����`�vV o��5l�`�m+��� �{����`�vV�{��5���/6��9S��h'��M�d��7�vV��� �׺�wB��m� ﻞ�{����^���h�,��:��7TrD�r�Y+o��U{A�7j�������4r�%�g�9�g,x�$�'#����ڴvw�@���S�ꪪ�zG�J�P��I�m4+�h�~ΐx�1		1<�
H"�"�i\3K��2#3ʰ0��UQbY6a��-a����I6"��%Ĝw������@�����F�<䭵,,lh�����h{��{����^ }�<�Ŧ2շLm���UqzE�}�Xy{� ��ޚ��;�"��X
9n�ϻ�Z�;�q�����s��$qɕuϝ���pg��Z���Qs�c���<H�ֱ�OiA�,Q�:�r�tW}���/��0��< ﻞ�ݕ�m�z��,*ӫi7x��� ;��o���vw�@�]�/��X+e�_��s���;qfn�ʂ�w�@>���:to���W��4}�j�;�� �{��^��>�*�N�m�M�wWm��^���s�=��xw�+@�;��T��Q�R6��v�6�3���mt�v��6%��X�� �^m���]]	;��s�=��xw�+ �/u�uT��1���cJ�x�{�@�:T>� ��M>r j�7��Wt�Z�� ��V�^���s�=��x���V˧m��ڰm��N����]���Щ,YİĒ��ى+�H��s�ՠ|�ǜ�L$n�i���s�%U~��K�'I��wӾzz�="�7dD�5U�
9�C��\+g��.ׁ�kqr\�;m�s���t®�*h���r�^����=��z_��s�F����첽�ݕ�{���_w,ܽ׀m|���Nݻ�ƨ�� �/u��w,ܽ�}�{V����)�*����$�@���`������=��xޣʸiݱ+LcM`�>0wvV���:��Mqg��cX$�����T��t�b�^����
��v�=a2L�R�nuY��֪;5&��zx	mu��w��<4�kӴe�vی�N�f�Vxeó�������w�)�Z��g{s�.z��C�C�#u�9Bg��%�1��#�,���ks�k��=-��ۆ�3��h�)��Q���*j4�,�$nraI���[%簏$fq f��'k#͉-�Dݩ7l�����K���j7'6�<�q��z;jy���n����n��x.^�=��s��l�U�"��QI$�@�߿j�>����� �˺����!�ai6�u�}��x����u��{V�ƾ<����BGS�Z��{�@���z}�j�>��]=���M6��u����^��=}ܰ����X��Ulm���ՠ|��M����:��M��<?<��ܶ�������y��:�$zzVc������C��u�]+��էb���������=��%�r�<ۥ@{�~��U�b��h}����1f$��s32+}�j���K�����ؼY[�!Q$�>������T��wںwޙ�y�^��"��QH亾��R�}�j�����}ݟ��ȵV���Ӷ&�������s���j�ꗾ�z0s�0s-��[�vڥbW��N���{��IT�:.�pv蝮ڹ����5#rP��s���o���w��K�w���=�<ӐQ���9m���������{����ʢ�ǋ� V]�E�������J������84����/�!J޻Y�ظ�u]��}��aof���l��:(
B-%P҅[M6�q`/!�DZ֮-*[n�b\��������j��$8�Y˨ƛj������NlI7��M��mx�oy6Ό�LǨ�[�D��f��C�.�|������?s�>��&�|KG��ĉ�m FA!���YL���K�o��$��O-R�� 3x�H�.�4f�a�=ݻ�°�@����9�|{�t��</V�:��4Fk�̰%`�&���o���m�a���/$0F��T*5�!&�N<�0�	"2�懢�C�M4lϐ}R���$�ًMZ���$�/Iq�f��pa��Q��s[ƍ�l?@�xz�t�}���i�ǰ��$" �&E�d�iF	(N���C ��0��T1F��%/:���JR�����R��g���ܲB�Gi`;V� �A����,�)}��o�R��{��pz�����3����� �@����I�r�X�@ֳ��R����}�)JRy�����R�����)JO=�^��ԥ)��}� |γv����L�0vSN���:�ls�m�vz���A��ۓ��V��:��JR��~��R���}�)JRy����O�)=�R�����┥'�ߙ���b�kj��%՜3f/߿~ո�R��~��/R�����k�R��{��ڳ�,�~���d�m��K+Nڷ1R�����qz��>Ͼ�\R����>��ԥ)��}ÊR��zy�f}��,�k[�����JP?}���)JRy�}��R��߾��(I݃��3�'�ͨ���_�����3�]?����Q����.� R��|��R���{��Q�߽����\ś�=pn���Tu�J=hn��pm�k�9�T�8�[[ϖ�)һt�~�>~\f�YoV����JSϾ���);��~��)J{��s�Ҕ�{��pz������7,��kv���[��1/���qz���d��~��)JR{���pz�b��ߵnb�;���?Gj�؃f���R�����)<�Ͼ��)J{��p┥'~���^�)Kϋ�h��̲�Z͕���)<�Ͼ��)J{��p┥'~���^�)O~��qH�A�ߏ�y����U�]Y�1'���)JQ��߾���R�����┥'�����)N�|�~�o�'�ꫦ��s�ۋ)4+��@���n�9'��6]���-=k3۶7b���+Ƽ�	���{)r�e�.R�Խnf���|�>9���)Og0��W��uwV�ŉ��7F;�8�y���{Gon���q�춇�ɂeH\r�v_	q۝u�5���eimρ����^8�g]j�
�X\l��g�7o9��]�\�,rۮ@-���1b_�Ķk߻r��k������e9�^�N"�-Vꇳ�e9���CY.fbY才�7��)JN����/R���}��)JRy��}��R��߾��)JN�<�1���Lq�AYn�p�A�����nbJO>��=JR����8�)I�{�ᘃ1}�/�����r�nbJO>��=JR����8�)I�{��JSϾ���):;�/�������ѽk7���=JR����8�)I�{��JS�~���)<�߾��)Jvv~�+��VZZ�j���1}�����)@���~��)I�}��ԥ)�}ÊR����j����o0ѳ ari���9��p���n;Np#�}v�seͻ�U��oI�Z�,n�89w3�b��}��)JRy߾���R��߾��)@������ᘃ1� ~�1�8�#��)JRy߾���;T0��B����ÊR��y��qz��=���nb��X�b_������2����tz��>���)JRu�����R�����)JO;�߸=JR��}�f��ڶ�[%�;V� �A����ۙ�1b��o�R��w�pz��=��qJT��w�o�a`�$���g���}��)JRy߾���R�����)JN��߸�JR�����<��Ʒ���Z�����D��kSV;pu�;,�;l�4n�C��I��H�6�{ݷ��O|����)O~��R���Ͻ��՘�1{����b���������Eu�ݽo�ԥ)��}ÊR��y��qz��=�_}�R���}���)����D�:�c�nb��������=�_}�R��22�M!�qRFI�� 1,�&"3a`�d$��$0T,$%�$"r0�1#���!I�w��@�^��ڷ1b��[���
X�Bf�[��)@����8�)I�{��JS߾���)<��~��)J^�{���SӖ���A��~��ڳ�b }��qJR�ϼ��/R���}��(�1%��}����E�C�X�#�͊\vGM��<�ŭn���[@�n�;�Ľ�t�_��U�D�-�B��V|f �_����j��'�y��^�)O~�\������Vp�A�����8����-���T�)=�Ͼ���2S�߷�┥'߾���JS߾��)JN�~��s+>23ZֶZ޷�/R���}��)JR}�����PiO~��R����>��ԥ)}����F����[�� �}�����R�����)JO��︽JPz�݋���,�JC�� "�]o}}qJR�����~q6���.�ᘃ1{��ڵJR����/R���}��)JR}�����R����Ϭ>�oF��Z5�[+��G�O<�ۉ�M�OI"��.�k��f��<9�w΋u;$N���;V� �A�߻�ۙ�JS߾���)=��~�JR����[��1����?�ʜ,�h��gR���kﳀ~��JO�{��R���~�ÊR�����qz�)Kϋ�5�uB�I$�nb������8f ��߾��)��9'�~���JS����nb��~��7�-q�c�m�n��R����)JR{�����R��=��qJ��I��~���R����?kV:9j���Z�1b\��~��� �+���\R���Ͼ���R��߾��)JN�7�>ݕ�ݭ�y]2F�y�x�_=)�.��k����D����dY���/�ks�\���^�3l�]���]^ng�vʖ+�ݟ`a�Wn6]�?��z��!�f��0G�[��(˹��'����e2�̆׸gs�8�xti=��έ��nlm�!��ׁ���W�W��h�ųg]^��v��%�<�:`"7m��q�y�w>3;7W2� �w���w?'�t?����l:�|�qC/b���y�����JF�*씧b�}��(T��=R81�۹�3f/����qJR�����R��~{��'^}��^�)K����_�Z5���ky�)JO=�߸=B4�~{�)JRu�����R���{�pZR���3쟜M��q�۫8f �_wߵnbJN��߸�Jҝ��~�)JRy߾��8f �_�b��;m��ڴ��*���!.I߿����R���}�8�)I�~���J�N���)JP���k?KX�� :9w3�b��g�=�@�'�����)O|��R���Ͻ���3f.�Oɹ�����܎*�9v�H�)r�]Վ.Nb1\n[2�V1������ʡI\���1b]����8f*S�=���):��~�JR���~�f �A�߿?�u�m��mGn�ᘩO|����i���4t�b���т�681�4�ۀ�L�6@�F��$B�h;S��R�\미�JR�}�~�*�������1������Kw��o[��)JN��߸�JR���~�)O���>���JS�~�ÊR����A���(�uB�w3�b�����T�)<��~��)J{�p┥']��ۙ�1b</~����@�W���'�����)|��R���Ͼ��ԥ)����┥'G��>�(��/6S��z�Iw�Rҕ��7M[�d��\8��s��~�h~��}�R���{�)JRu��}��R���{�qB����}��ԥ)�揾3{ַY������qJR��>��/Q�G%<���g�)=��pz��=�߸p�@���<�Z���Jt��g����~�)JRw����C@��MG����,0J0 j����� �!$d��ԧ^����):���qz��/�+�d�h�4��k���/��~՜3)��ÊR��y��qz���������1}�ͯ��2�c��l�������~��)J��︽JR�{���)I�{��JS�>�k�+>ˎ��qk qw���Cn�U���a��X��4��c)�9����w|_=��b�Ή�qJR�����/R������)JRy���Uz��=�߸qJR�����8�#m�e���3��~��,J����=��ԥ)��ÊR��w��qz����~(��բ�ȷ��R��y��pz��=�߸qJ �I矿~��)J^~����)I�w����F�W$��Vp�A�1/��ڷ��￾��ԥ)w�o�P����10!>^�✓�u���)��z/ߕ�0�#��*���1}����)@~�=����)I��}��ԥ)ߞ�ÊR���^{������%���(���gq���6�h����;�(���)��������Z[nÊ��R��ߞ��)JRy����R���~��JR�߼��/R����{��{ݫU���o{���)I�����A)N���R����>��ԥ)w�o������ѯ¬E���W]���b%;�߸qJR�߼��/R(�ߞ��)JR{�����R�����E�3{�o{�f����)K� ��>����^�)K�~��)JRy�����R��� {��)JRv}~p�~�f�k,͙�޷��R���߷�)J?��������JS�~�ÊR�����qz��1᧋���4�a���j�B$�z-�k@h�ք֨���
��ǀ���g9��C��&fq#�s�
jH��ں�Μ�ș��/��k� 6�!�0ia�A?�7sJ���H���f7I)�X��po��8��Z�bOS���	�����5��ѝ�8zW��b�4`��1�id�u\���1Ć��>BQS�<M-���0DM��ы��i"��9�s���N�2��`qx5DDC�ٖ�O�k�Akn��ɛ J��r��u@UPqJ�i]#��}UuT�-y� �V�tT�����ڣ��ۑW٭��cA��]���U������k���۞NlPu�6�I5�k.�iIboc�]�KFe���7�&�m�Hu�nZ��&x�m����C��EK�T�9�穭Q�&C�3x�=��c�SOj�r5���d���;M�k�H�s��xE���w/��Nr��suۍ�mVzvۓ�k�v�qe�vq�qV�f�\�H��ղ�2�OWN:����B�K�9�69�A�a�]���[OVNΗ�v�{�}U|��mU��cE�ƹfh
�Tp� ��	����5\h[`��q������dP�D�r�h�N�q�\OrY��]�^`v۶�[&��Ba���.$��:�+�8m�P�{v�O�?gvݍ�j۴8P��8;v�.%���Sb��nM�W#�k�M�vz6�S��9y����rhs�qO`�v�=��3n��`{3�C�y��6��D�D���cs�3z�h�؟B�=�ζYk�ʵcs8�]���]�3o#�g�&9�2��.�:����t�z���ɨ���<�:|	�ݸ�z��5��^�I��	�*9Km�����$�҆�kg��v.���%����mH�V3n��k��෴8iU�)�n�c�m�v���d����:󶛫k��ۖh.�]�	��Ǯ�6����6���-��N<��v�Ո��s�s*# Zn<��.�l�[��91��u��r���G39)�UŶv�g]�lnƦ%�jS���Ӝ�&�ZN�V��8J{g�ۭ�v#��Ӎ���6�b&�A�a�x�,j�p7��u�s�@q����0�c&�7Z����4���,#���vm��f��Qsk�`m�`�v�
�\�n�4]�p�5(�a�@F��%�zy(k���}�����v��u�*wh��rp�1��&'���e�k���3ʾ�0����y�r�6����n�^y�r�Z��mWb�L�N�F�ޠ��'T%�,ݭ�y���>O�����1:�� �W��@q��ꢉ��Tz�fv��ڷ������˭���2�3wcZ|Mn�����9f"���i��X���^��[�����=�jm������=���7&����펮���LǦT<�=�����d0,f��!��Kv�71ΐ��q�G�Gl����==]v)GWB��\OF�WOY���#�[��ۘ� ޖ�=n{����+��:��Z�MX�u�k���࢑��3Yh��T
�Z��Fu��Y[��RƎ]��g���g���g�D<1�;Z��r6[���`�@��KaTE��bJO�~���JS�=���)=���ԥ)ߞ��R��w��}��34f��Y��o�ԥ)ߞ�À����y���/R�������)<��~�� ҟh��z޲��٬��3{8�)I�}��JS�=���JO>�߸=JR����8�)Cמ�����N�������R�;���qJR�Ͻ��R��~{�)B�{��}��R������#�&Ul����1{���VpĠC�=���)=�Ͼ��)Jw���1b\���_���%2�$���M��^�[VQ�b;`��h�_n��ny�����_'|Q�Z7KU�۫8f �_wߵnb߼��/R��~k߳��Q%2����۠%�*�Lm���7X�鵺x'���<H�2L�,�002F(	 Lb��!&PP8���q@?6�����V�.�J�=B��#��%����������8bă�t��;��Z��PR��);t�&b��po��c�@7�ڰ8�_yt�}��Q:�]�����{�}�X��7�Ұ>�q� �7v���8�Z �G;�[]�U����<�8u�����R��F��:ٻm�_w�����d�k�㨈��nՁ���(��q	q%���������V��[yZ��8����y�݁��Ҡ�v��� ��u���Z�:m6`�M�>�N�>��J�' Ng9��U���{�~���-
[I\��f,����^Ƕ�n�i`}�P4s�\��$��wD���Lm	�7Xw>(s��W��
3��c�@7��0=vL���w)�\�][rm�:P>ʗ9x@�k6�*bpV��ܪqbĖnH��ID�;=�,���3��c�\�J�P�d4	��AE7m�L�f;��\\�}�t��t��d���%��w=�U �������}�V��n�b\�8{%���v�өGI!rX5knU���$��1?��o��;���_{�u�~7~� �\%q�~�T��~�Ô{���e�#�Qv�����$��ĸ����Ǵ��nՁ�c�~ܢ����1�@\*�#:�ɬ�%�#�v�vd)���n������k����^J���@<�w`}�t��n����� �t��@�lV���v��{�*�9�q �mڰ>�K(�����8���%V��N�4[bn�	��k@��,�Iqq{1݁��Ҡ<��D�$Q:��\,X����hw����qҠ�I$_��,�j�]3!$�d�>�c�R\8����mPc�Ӏ}�_Ɓ%y���o��dV��ꗞ����XW�C�����k����oIv�����i�+nY�Y����e.�Ҁ�����t�%^�6WW�a�9�{'m���}�E5�ț��W�z��o���v��mg�UzݵÀ����W)��Y��;��s!�j�7 ��z��ǅ�G��Ѱ�g�e�E�YtX�CՅ�h��T������ӚWq����ආ��M�-]��w{��ｱ���x�$v����������X�8�[m�yk5JD��;���y,F��%QF�
:�9w�~���Z~�L�>�K).$������R�GI�&I�3*������D�:P����>�j�ı�}�m���K��5E��d����;��s�>�t�|�~8����Y$�8�V�M�>��v��J����_{%�1��_�;H��d��wߵhً,\�=�>��J�<w`}B�t'��M\�N�ڒv���n��g�VF����l��o���}��>{<+�+��2���,�>�c���`{��P^;�1��h�FT㳚p���5��.$�q..��q݁�c�@_��/W8�s�� ���#WAL��I3�(���{*�E�t��9e �����tb`Dvn�a.s1�����>�p����}���)�Z�v7m*N�:�7�2ގ�}�X���m�ۥ�@epqE	ev���pz&��Fۨx�w:��J`���=}�{ʵo��6�tU�y����� �{��{�VU~��I���ԑiRB4�(��݉s���Y@[�v������ �t��Am�ګN��{�}�p�7�=����)" ����«�i���wM�w\T*-$�j��I�����o��X{%�}�wa��Ėw߷��:��ߠ?�D���l���}�P8����:�>�K(��ڰ?�w��<����Yh�U,#�w#l����XkY�>9�G=;��NطWX�L��;u12L�K}�n���,�/��K�����O���j՗B
V�����es��@_�������n�Ws��P6��lt��0L�OWI��@{��Ձ��qA�s�=�����}��bk���#�W ĳ;����9��~� �߷�ʕ�C�b�l���tuQ�*DE�J��Wi;�7�I��8`}�Z�Ix����I�e�J�z�'aۍ5ؕt�uk��mn���b{:�"�l*ڗ�ŉn���7DTQ��~Δ�{����\���;����N&�r�ƝTr�>�qp�K0=�n(�����9eoI$$����@�j�*-�V����t_�׀o���\\��{���{� cv85�]��+�13\K�����,�/�ǵ�{���O���ؑ`��S�$�@�9e .$����Ұ=�n(���w�����y�=�`�5t1+]z�D97<�k��zWV/\�>�f�X�c��wVН������1�x���,��MF�v�׈7aG3\7m���X�n�']��y�n�m���{XA��2A�/e�\tv�r.�O�`[����rluu��@�KųF��/b��݀��-�m���Jcu�ԩm:8�4��x4�8n@�Xj��9]k1(���e�u��WI���o3�DH:�{�b�ȴ�4�����)k���JX��O<vW;U����F�j�	1��Q�}O_�����5Yhn�ն��C��g��ց�Q�<w�Ē�=�Y@<s�1����+���3J��u��qq$������t�3��K��qDh&���'bN���G{1@{^���,��\\3���Ix��[�[ӺI��+�~�^�,�3��������s�J=�v��������v`�vI#�P�t��$��n(�7v��(x�9���>:���V�{d�Wdw]M�Y�V{i�i����{q�;���N�5+������߭�g[�����9es�\>�L��/Ĥc�I�n��t���*�Uma�!���2�tlLN��Փ���iM�!����5PaMU����Ћ��ڝ(�mi`{:�R������]�@w����37`{��ϱ�,�$��$�������3���{
Tu��C�����=�K�>����fg}��4����LR�Ɏn����9�Ľ��X�,�>�t�����j?�(Ki��A��,s��Q�u6n�����1����u뮱�G�]�{���[z���Gc��e�f(n�݁�r�31.s�\�=�n(&c(�2�OI;37`{����L�=�n(�n��bŘ������N �V1JQ�h�����u��UJ�=�RGe.Z�O;!ݹ�p�c��ޜ�����aQNӆ��vf¹�wۅ��O�<�q�83���ڧl�U,O�0tz-�PĔU��Wt��F�A�����ٖ�h�)�($_;4h�3�4APR�ff�e�՚��C~`a�����$�@�cF�Yd#N�X�
�&ԙL��J�F�=�����s��[�-�ʖ7.��ϋ�1�Ğqs1"%G �1�y����A�s��vAG���)0PFt�[i�5��1�LsQpw��z0hl��)L!�;�{l0m���Y�8=S���à��6͛������&�<�N��Ļ�Y&ȀlT��ᩉ%4�s��3G$֍�wU!+a6XV.�j-6&�
�i�E AcMcbm4��m�\]�.�sZ�"Hq�x���_w���3EK���5Q>bRIԌ�z�j&8�`�0%�r�R	���>�&�|<E`ݣ�z�>����{P:P#�<^K��$�����z����e�'�i��*uckp�+�~���R^��n��wL��IZ_�HM�Q31@|�w`qs�K��f:e��R^��ur���"�L�e5g>�Δ]��(7v�n��1�m0c�z���]��p�����~�T�Zo4tp�;�L����q�K�W�Ġ=���ڞ�$�0u۵HvـwӲr��Ot��8eW�=ӰNeYI�jʴ5�h�n(?c�7�H�9�3vt��֖y�~m��*�J�Xw�}��Ͼ��*�����T		�$0�,K����@�����7ce�R:G/,7,�$�|�Y`fu��<���7��~~c��Is���Ѝ�̬[�Ǧ�&�u	���{`�ꞵ��^^�w?'�ܻd`�v{vd��֖g[����.%�zG�|(�Ej�S�;{�������;�<ܲ�ϞS,�I ��~��R)1շm��{��bH�߽���Oߞ����?J�L&5�i��*�{���N�h�%���wSP�1;�M���`�솁��g[��1݁�r�R�����$鴸� +h��W!�nr�q��"]tF�k�����1c����۞^�V㺻GB�v��z���ۖBy��R��6��ā�,�r���%���ǣ�.��\l�����u�{;�N[:�lv#�#ٰ���nZ��l����{ztAT|�l�E�q�i���ۍ�:�Qݞ��s��G[=��S�/jٞ��e����]�ֺ�ր�����av��͜A�H1\NFqۍ�+�Ng�]Ih^�=�3q�g��[]I������-�n��������ttp�;�2�W�"�Ŀ;wi'x��t�@{�xt� �H���C�B�Wt�$��� �74ct�?=٠3wv�$BB��ĝ�i��L��{�<�I�}�� ��]D�vQi����@=� W��4�8`�d8��E��5�H�#R[)h����0xy��+G<�ٸTu�^�&���s��&�o ��n��G�L��{�<��-���O��{�}��`�>1C�ZX��td`$��>����,��4�n��)뎌n�&�"�m�t� �tx��t�8`�V)�f~�x�E]����%���n���Hs�=�����(!���v%�۲�o ��7@�G
1�2�=������݉���p�l;xeWn�i
\tFN;(���=q�3����ňZJ݀�ժ:K.��_�@�yL�csK���݀�cj �'e]��e�`ӲW~��:n��U���.�Q;�-"�:C�����߾�*�����*�E��z+���V���&C@'EJ���$졦�	Ӧ�{�0	ӲW����w�ԣe����t�Ֆ��{�0�~�9�@���N�7@�G,����L��G��}��i�Խ��Tg��u��#jK��룖i��ɍ��x�`}�P;IX{%�͵�e^~��XZ�4����:t��s�:vC@�R^%WL�/�;�bfJ盻ْ�Đ��`}��4��߃�uF*ժ;��b�Y@?�S,��(\� �c� �Wi�Wn�T4�};!�~�U_t�X�t����I-�j��V*R�^��Ȏ3�@g�ec�s[���:'�	{v�.�qJ�1bF�W��D��GwN�7J�y�w`{2Y�\�.}����G3�
d����������Ř�X���J}���>��V��8��y�kt�����{�t���'�d4�L�w��ޔԻ�N�i��l�%���ڰ>��P<��糸��$���g�^%M]�yZ�&V��qkǿ|=�(��j��9ġ.	p�#U22 �%)R�(�ҘJJ�%�10HB� �W�і����N.`��"2F�s��v�Ѻ�T`����j݉!h���=fbt����V�N�kf�;��c[7s��$�v�NJ�;{q��C���o<�c'{�=��W���!��V�;n�\�[Gm�;Wc&9�܏0d��rZf��ɩ�3����;��^�Wgv��qK��훰X��ݸN�@���-me���"�1����\|�֨v�
c�����w{�`���H�;L6u�k�ۢ�grm.ѹ��7+��'&����2��j�3X8+�YeZ=�����`{�@}�b0}�j�[�+Ottp���t��=�e`�M��_]tBJ��-����<�X��Pw`{������Ƭ-P�:b��h��&V:Gv��(?9�Ď(׻ZX����5�$��&�`���w�e`��hN�X���Vƚm?Ŧ�*�.��-�2��s�l;u����<U��&�㋜���t�4��ue��{�V:L���n���Z�׻�`c�=؃���I*"	�ʠ7L�\��q%�8��<�Ҡ7�&��2��ڒVG�g�X��.�=�VͺT��٫�\�m�*^��ց8��*�uh�o�v�`���{1Ҡ6�Xl{^ڠ=�hf��J�M[-��{�V:I��}$��'I7@�ҊV
��V���-ں�wɨڛl��۹׎�7kn��s�=�n���u8R�WV�M�m�:I��}�e`���{�e`J+�\,j�+T��m�ht�X�&��X��k@!��EJB��VZn���twL�2���%)����J� �?o��V������OzR��bi���Ֆ���t�c�j���T��1��X�N��:���u�{�M����:n��I��u��.�J�?ɕwm8y��V���[*��q�>:v8s.�8�\vC���̬���������=��wN��}�e`��ց<pҲXZ�O�s2P��ct�7�Ձ�d��D�P�	�I�=�"{7`{7iP;VlFc�({�v@�ӳ3=]��݉:�'I6�{�0	$��������A��F
b��G�"+���Z�_�7����H�*u�x�}��x�����ݥ@cmڰ=��r�-�=n�l�k+�-Ձ��X<ra�����[l\�Z;a�b�]c(���ܮ���@cm݁�7J��۵`{�,��Ԣm�b�ue��ޓ+ ��mX�K(��ޥ��D��Pw��(P�J���U����{%�cn���*�t:T�����x)��V����I�ޓ+ ��mh�4�T��ڲ����f�$��t��=$�Z~{��T��J"%(�H���I�	%`�ƋF�3EL�6�ց�M@�dT��g�h�fd��Y���
1�`i���~.��(fNàR��bHX�� ����s�U:H��&��*-a����"[��	Hb!!l^�9�n.;��6��nc�0�C���	(�aB�).=Au�6�9�,�t�#�V��@��ę*&�!�D��V���hi��aH!��B�<�Z����+i a���+Ƞ�Jdf�#mo��CfF��XRY��h����Č#�b(�"7���Pt郣�Q��
p̣s�3�A�I@DA��I��;.$�b1H������ڞ���[v۵/!�*���mJ�U$�m��9�m� .��4�m��s���;q�N5czMLP7-a�-�#cF���:�YK7;;h�)�{@���Pe����ڐ��;�/UU���Kr� !���s����Q��i�6�nU
oc�]չ4�F6ٌ�U���(�"��_] ��8-���gu��v�*��i]���m�/m��g�1v��*���×u��ۧ��g�r�s���[���kw��I�N����VVz`M*�[Q�ѓ����e�j�D�ǌ	/p��݉-�{Nݛ;)�	s@l֗&��2IO����Qp%V�L�0n�PU���ܷl1�c.�n3�r�'Z��ܚc��z')�0n;)�@uph2Dh��s��Q�ZZc�Q���I����%����뮥۝8�.�q�cڱ;'&�����@>���]�MI�'��N�n�v�;�9�=���Wj�#mvvhM�X�sc	4���Yw��5n���^aîG=��NLq��a[�)��뭶g6�:�PO�#�&v���X���c�u�ϗ�����㷶˳ݏa6���o'm�u�qQ�j眦Ȏm"��˱�l��g��u�)�c�3��m�.0��t	x�K=�n��3<�.��Z�������7[W^sk����+�	u�tF�^�A�%U�d�.���uh#��`��n�Ov�m�ţ�g�uL.��-n��݃��W�g��]��$h�;L��m#���m��pIjD�<�W<ᮼ)"p/��*��N�ѳ'�3��n���u�Y�N�*�2��m�ƗFaa�
�Ӧ���m�F+�ݶ�=v�YG(�7��������������4��[��@�vl08�N���^1�ј;
u������s�n4vNj�Dif�u����m,9ĺnM��]�
��m`�s��j^�gFu�<��s���;.��0x�{d���͉ݚ��!�z�/L`4�
�1Z�K6�����Xݮ ��ř�,X,K3"B��=l� )����x����'����C�?�{��}3�Y�p]ؚFu*L���v�����z�p�\d�u���w=^�ƺ�s���]`����=�Hi�mؗVx��W[�J���m�'8P�q�x��dt�ː��h�C�e����
1�gdwA��/f;����Ӄ��{'$৷6S��&��sb���i��pJ�W!����Ν9z��қ�U���z�k<<G�i�V�5�z=�@%۫��n�?�{�ǽ����~���U㞹�*�/n��٫�T���죦--C������1p�qX,Z�$&g~|����v�����.s���۠K*O�-	��&Zn�n����`}�P��{*�s�K�j4�݀��;Q(&{6�c�(�;�>�L�t鵠�wb%���N�CI���t��+ �:mh{�0w����ěi�-��Ot��+ �$��>�8`����!�EBm�����q�V�N7/;q �Q<]�$�mU�Sz6��/$��.�b�������u�N�mh{%���������lmlU*�:D�I�Obf����YP���$�Q'[�z�镀OI6�	�4�T��b���l�'t��}�X��k@���oW���N���c��@��2�	�&ց��� ��7@�+�YhI�hwm���}$��>�8`���{�4����ߜ��#er��cBt�/D�j��]��IҤ-�+�|P�)�["a�TJ�fՁ��Y@~�kǿ|�wc�s���7��Հn�"�;]��c���P=��R�8�f9Ҁ�u��9e��r�I�m]�-'���+ �~�A|IT��'��o\���M�%w�
W�M]�wi��:j�>�P�c��Ƕ�f���"�V[�S�,m�hz8`�t��镀wӦց*)WwJRB�t�]պ)=��z2����ڣx	8r\�����㮷b���K*�][����f���?�@��e`�鵠}9� ޯJ�������V���:Ty�`|�Y@y����%d	��B�{'f ��Dʠk�VϜ0(��7@��+ �Q눀[W]�=�ڰԗ!�(׻v<t�:�E1Q���M�e��t�1nS,��(� �Ȣ�� � �R	�,!����A;�;���:����$U�P�ح�0	:M�:t��$�6��p�:�A�߮�! �v�4n���L�<��Q1���iGn�ۭݬf4�ڷAj�ݫ�E�{�zt��'�M��0	��t	]H*"1�h�{3�ʠͻW�͝(m��x�z[�2�ݫ�uM�%m�h��N�M�=:e`��k@�{�b�B�b�[��l�'{���2�	�鵠t�z�������n�[{�t�J�ջ�~_ �gJ�c�9�K���ݻ����~��\l?�F�Mz�<����l(���]i�	��I�;]CjwݷO77l���s�a����*�W����\��ug�g�1��Y���v��s�N�WM��0���c���٫�Z�p�q��;'R�s��X�ٝ\+U���������T,n\�d9՚YU<p�Y�t�<�m���A��u�;l'0�"E8����������I#�����v�|��ݗ�<ӷ/�4(^����ōc���C�^�"r[�7#�m��wm��l�M�{�0	=�h�2���r�B`�Ҷ�{Z�K(����t�����9�D�dGa�&d�t���=���T^c�{����~��H�C�h�2���ڰd��o�݀�]�t���R�JҶ�`�M�w8`�M�'���=RQw(��T��ڱӎ3��u���� �������@=�*�n�M9�������wn�0���N����zL��$��:�(uh�
��s2P���"���r��t�|�ڰd��qs��6(�d$�ʙ���n��ݥ@7��X2Y@7�����X�HN�v�n��$��Z�p�$OI��zW]��]����i�h�� ���zL�I&ֆ���M�~G�m���jT�6c�ü<��6��V�xv�,vz�����6e9s�wgU�E��I&��e`I6�	��{��D�&4Z��{�OI��߮��ݵ`n9Ҁm�w� z�D�;�L�Wy+�Lʠ7wvՀ���#�Z��Pba@UPA0Ce`da	S:�b#�h��B���2�($"$C K�D22R��$CC2qL����	��!\W3��� o�z�~��κ�^m*>y��*�EDO$$:vf���%�m����@6۵`}��(]�	��M��M�;�2�	$���K(LBqv:�HJy
&���W��qE֫43r���& p�p��̈�`6�؛��ot�L�I&ց��I�t	et�"����ۻmP;V�%�ǎ��:T��u�}()X�+�?����>��I�7@�t��$�Z޺�/�s�v'}��~n���*��j��ώ.)(�	��)Jf	?W�.��t�Wq�%i�vZ��{�}�Ҡ68�[�_�Δ~�vb� _�tEbm0�+��%��5V�v�ַud�M�8�d���U�ny�8�ܵ�e�J�L̪�c�`{2Y@7�w�Xc�Xt�QW�o�؄�V���
�c��n� ߱ڱs��&u�lB���`{��t�X�鵠{�� �W���cN�ۦ�ot���*�nՁ��e�J7^����'��HM�����u�I�mh��3%�x��6�P�9���䈅1 %�BJ�5J�@A5DL%!P�K	'�hϳZ����[��F͕u;�5f�[H��s�q����u�d�X��=;.�%9��pcg�ek��6����%�&�G	���[����]m�����7���̘��v�K�v�c����X�gc�W�­�EVHuX�4�q���p�Cѭ��N(t��Wrhݔ���rv�t�Y�pG�$�+�ttN�3�u���&ۛ�����ֹ�QH�R'�$�%b�f(���$%N2r���q��h�۴�<)ɝ��3���Ou����'�uL��(�2�A˕���z{�������J���nՀ<���C�V�4+v���M�>�e`�M�ޞ����RO�	��8��� �I��OI6����	�&��)�+�H-Qc��� ��mh˥�1��9�|ۥ@g����TErPJ�m��ܺ^;���+ ��mh���=�����[���Q�]�qq�n˺�^,�^3���9yN@��z���{�=��l��YV�Zn�	�&�I2�	�&ցܺ^�^껺%�;�n�����&W<G�@�XI �Dؽ��*�vI��}��Ot��u���J�Wam��� ��6����?�&�I2��T�
V:J�O���;�K�'�M�>�e`�&րN��X��̝��=��~���ԗ��V��j��2Y@o>�ƅ���vg�����ێ�)��Y��#k��n�r��,��Ѯ3�kZ9�)��MA%���7n�~�ՠ?cv��%���n=۰3V��c��ބuJ&{*�~��_��.r7:P�v��*>o���(]������f���d��~mݞI{���1υ(J5�߲��i۳�@����u�73�3�� ��T��z�3y���a�����N,�F,Daac`Yu�)�p9�
bR$ �Z�����@�tkX�b���F�F�!�]�`h֦l�sR�,j#zxs{�Ϛlk<�K���.J��F�ū�'A�]XX7F��tt u��E�\���u�+6�]t����ml�
s�4.�ƣ4D�`�θai:81���!�o��	���Y��5����5��a�2'k��qÅ�;�b�B��]�s	*5�fr#�2�p�a�I��<��XC�"Fe-�2��ޜ%4e����7����-t�kc�lT;�AhM"��5Ш��@v����`���� 	��+���~��{Õu�}��^|Z����=;؞�O{2P~q#��׻v��,N�k@���o����v��[�����{* �mҰ>�K(�w��~/⟝�;<\�R�3m�>�܏\θ�-��u�Mam��%b�h�t�w�D�ut�i�� �I��}�p�$�m~��t��>�]�F*uj�O�i�h{%��q(�wwn��=�@6۵b�u�K�ܰ��hv��I7@��2�	$�Z�]/ �q�@�իe�- ������P��X{���>#��4�PR5Q/]*��~����^���b��5Qd�@y�ڰ>�q� �7v��J���gp?7�ůV�k�z;3���v�˜]1�ֵ�N�@��'^7l��z���>O�矃�^�7{4��ױ@7�݁��Ҡ�v�JWȤK���J��m�;��*��c�@?6�X{��s��A�M���Ro�v�{�{��V=$��>��x�t��"����v$�i7X�Ձ���(���l{ڠ=����B0�v'�M�hyt�{���t��_y��tuW� f�*�ha��J����,"�!���n���<h��-d��]���<�L�7J�k'#E&I�r#\�$CkkK!��$8��v���4�h㞮/&b�'����J�d��6{+��g:9�:}\���!,�sw.�@u�ݭs;�W!.C��m�� w7�.�@yΉ���ON�-��D�z�˂���ґu��}��x).�M��V����m��,��w��9��s��fܼ�&�碷��~{����w>����;-l��m����VW/Vjn�:i*�6psob���q #�#��+���T������7v��J�~��o9���O��=Љ]�v���P���>�L�{���>��x�I�J�%���vR��eP1�V��8�b77�@�O���\W��e�S�+i�X{��~������P1�V̄ҫ	�Ut�n�	�&�{�V;���>�tX��J�T�WJ���<a�ڷm�k����Xv8W;�Sٺ���81�v��wT�:j������t��6wKV��}�q.q+�~on�p,��]��6[,�h��~���$�y<o�����30Gh��n(�-glX��7@��2��N�L��ZUj�ok@����;��t��V�N�\ ��I��`Gm�����K�|����*�x�XG�����}�����B��@�G~�6�_I4��~� 3�����Z�S,r�Gn���s�ُ\,m�]�]�)��� �;��L��V�i'X�:mh�"�=��n��&V�H�+��]�:��sJ��6�@{�c�1�T��ڰ>κ��	�T����=��n��&W.*ҋ�ʆ��7��U�y���:��.�ER����14�@�+ ߞ;V�����=������= �ff;2���`j�8�ww{`g��n��&V:U��.�+wv�6!^��+�{W9�����b���c)kM�p��J{*p�4ˤ�%B�E�{Z�H�}wI��oӦր}�Wp�倮�����'{���e`��k@�� ߫�uv��6]��I��+ �N�Z��X�t�W�,V��:J�w����j��6�@<�wa�\h" }�s-h�h�2E5�+Mf �E!�ЦB�fR0D�ES�1�7�U�NW���)�;.�yZ�H�g��1�Ty�Ձ�K�Z�t�Ʃ��맃�k���5�7���&�d�����=pW9��SS9;�r{uӖ����m�������3�@?<v�>�/y	�N]X'hbI��&V��6�E%��n��/�w���!GWzA���ީ5��`{;����˰7�@|�6�$P���
����{���I7@�I��{Ӧց��uv��uj��i��m݁�n��<v�c�PĒB���X���G�?;r���*�Y$��k7�N]vv槀���5��5��t�d-�h�;:Z�!�u^8T�ra\���[u� ����:w/��ܶ�Y�/�[�'��֌���u��&�Yc�i4������ʵ�듞xv{]�Lq�PZ�p���;l񅵆��Zݝ����  ��{�����ˍ�,N{6�ٙgU%>4rZ��$��x2�L�݇.���$�b���!Z������Gb��n�<N��rU��r=�㮶��5�QZWlt:T$���L�Ӻmh��w�M�%B[��А�V��N�y�`{���ͻ�=�ҭID�Yظ��JQ1ٚV=�(|���&V�N�Z�*5��J����)��(5.%�����ǻJ���;V�8`��u�ASo�C�1$�@�I����;V��(|ۻ<�Ȉ!���c�l�m��^��ܼ뜜�z��<��j��¨�-�x]�����]����?��c�P��v��T�f'"����T7/ �_��ssŊ��ߦ��e`�鵠u��E��T��d�=�n�f:Tj��׶�=��@����ը�Q��$���l���ڴ�{j�����ͻ�c�J;;�����X�:mhtp�=��tf:T��i�":#d���DLw�$"\9zN�{M�^:��3B��C��"�p񵵻���R�������=�(|ۻ��+ ��M��*5@JT��)*�ܔ�m݁玕�<v��P��뺊���i�$���2�zt����O�a�*�(��T�as��ݛ(�ͻ M��:v"TJ���۬ޝ6���{�&�:e`J��U�wv�M]�ցӜ0�I�N�X�k@���N�Wj��<;��rˎ6�8p>�]���.k'&�m[F�;�t؋�CJ��Ҥ�4��OI7@���k@�G�ߺS��bT#����%��.$�ovՁ糥 ����8��5i�6Tv:w�IQ�S%�7mXc�P��̖P�Ү+���N��i$��8`_y��u�^{���Zv�iH*e����n��>��~���]���%*Bn�ҧi� �N��{�� ��Z�0�/�E�)vݧH���l��^��4M�fJ�{z��91�ds8wl�s`�WN�i����otw8`��k@�G}:n��WIb����:v��N�M��0	��t�X�J�Q��i�&�V�ց�0	��؆�iP�vՁ��:�
���0	��t��N��Z�X������;�����RE!X�%� ����y��XnY@?<w`~�Z|���̬� �A�4%'3Z�mO3Gٰ��7Ŏ����4JVp���!�0��Hi ��l�`��$A����6��g�� �"�u��o��y�7���:#;���+��aKAA��Ʉ�y s�4�}�:ۣ($�	�Y�2�&&	
�j ���"(h*"ᆍ%5��M����u�bDΠp$,��\ڥ]ZP)"�ff��!5	��Ό��&�`��,��\�PAK���ޒC1�D�%��	+�4�Ƭb�,,ӑ�F����p��)�Y��1g�y�����{y��;��HuPBI���֮ 좼��qG~cq���:\�#C�@E�Na��c�� u
;�a�K��K�H��wk,�!0�қ��z�0�'�1MųP䮡y�n)w�����`PE�rM���7�oLeaȁ�لM�9Pc�Y`T�aܺ�7��h#P�`��4Rf.��nc�����ָ��Y�l-V�(t0e��X�c\y.XE���ea����kv�ڮ���3K++[T�UHt��˳�rUUUR�T3y�'ظ#CnҖ��A�u]]\�<^�k�Z9H8P.sO�M�x�m��d6!�{+��RkuT�z�:�K�XV���/S:uٛ=gTa�Fۦې nSM����z�+�Gm'��˘x�����,�qd؈	<&Yt���;-r�Pq̅��ӻF-�;�N�=,=����N�<�������,񞎀x���6��v�Y�#nTL�ע���-�9�m
9&Γ���懶�M��M��;��n��n�<m��S��q�j�8m��v���;Z���.���d��.�ݺ��B��U���]�tu'
�����Z�w[;/.���\���3ɽ�t��L�CeJzť$��6�Ð�u����V*�:�3�sAݶm��2���C���s�S����r�w�9ꋶ�v�v�ۭA� ۞���r�7�]�W��m�/2.p�G�y��
�9�b�$�FѰ�qļ7��;���.� D�̶��Y�Xqm�A ��:7�l���7M;�m����j�9�x׷==�������A�B�g���`���zڦ��g���O;��#��9�͹]ǘ!uC1�[s�z{O��&��<c�����C�0m׳���!�ls��p���;<�"�MM�Zn���`Mv�G���́���3ۧ���zuc����s�˺;�6�ʡfl˚�WQ��^��n˭G�D�ή�pI�Q�N{l$J���ı�a�S�l�s��ͫ�u�q����Ǭs���ֹ
�-�[GgaWJ�6ˬT�AYv:T�r����Ht2\���n�	�b���P�i]�M�ev�mt���Y.݃m�t��$��ᗀ����tOgqgqٶ�W\�P��7\�l�� s�Qѱ�9�)�9�`��m�����м	���t4v�8lے#c�r�98��u�l�Cb�lV�0�ч0<�6�.9y��7]wvs&��j�F�M���ujy��Y����{�B)�G�@�o�=炡���*�*#����x"/h(�<T�u��kGT[��9�a���w;G��`�ͨ2�+v)�=��f8nx��Cl��q3Ѷ��V��:�+͵\�e�f�1��>�r9�n������]â�M�8Tr=$�����l��A�T�n���Bc�u�{M�Զ8��wc�;s�z��c]V��sJ�n8��&�u�S���q>���D2�n1n=�2ۍ��e����P�'JV�m�K8�Ÿ��fث�������i�� �n�m�u�*]؜v�ݶ��K=f7<��C�!w7g����������(��>�ogJ�Di�ve:we����=#�=:n��0	ޓk@��uqYDB�M���M���tp�'{�ց�0	��:�Ke���Cottp�'{�ց�s�������V�t�e�rL�@<�;V�.$��i`o����,�5%Ǎ製J�B�fT̩�PvM��}v��r�qs����)m��n��3��\���;��I�wV��|O��`���8`�ݐ�%���ĕ��T���Kw*뿽����FU�o��{�mh��oߺ����+I]ۡ$�@�9e�;V��(|�݀�d��V��Rt bl�==�k@�G��7@�G�:Uܻܼcv]��Ұ=�Y@j��w�ǳ��<v�y�6P�%Cv��D�u����nqg����l+�n��۔7C�h��XT��O!O{2P��v��(y㵩$��ǳ��1�TH�L����݁�r��x�X�,�=�n����	%c��.�cl�=�&ց�\?g��s�\Ir�2ۻ�r��k:�eGʎ��$(��V��\�ݭ(�ݻ1�(7�Ff����4;�������մ�ޒn��0N�k@���E\t�;�Rl�m�4�:��q��l\u�vnη|,���On�\��s���^Dn�դ���� �I6�H�w�M�%Nup��ںN�C�ـ}$�[�.r ��Ҁm�݁��'�Z��1�]����$R^;��?����Δ潵`|��P�"N�:L!٘�y��r���a�#�/s���v�� ��u��*���i��8`ޓk@�,��7@��%)S�=�sW�]u��\��vZ�_�<Ζ�3�k��e&ȏ.c�^�����`�I��u� �zM�=#��uE�E۫I6Yi=���X��n��0����:�@J�$�Z�T��X��n��0��C@���w뮌�*V�]ۢ�{�zG��L�1���ԣۛ�X�ʅ�ٙ�$�T;M�{�!�H����7@�8`�����	��[.�i��-Ҡ���v�h{c���:��2F��8њ9�R&i�Ǟ!�x�$V{g͚���ܚ�`�H�J�r�v��{<G����5۷n��n��ý]��4�[٨�ص���8㫖�Z�]�㢻x$�t=���;q�K`j}�I��k��p�]y6dp�ۯ'c�z;�����'/ci���ۙr�XNKuOf�����������݊��������Y��7Fp��gV;+�]\����V.Ć��q����������|��W��w��@|����e�x�X>�U�e��V�-7x���H�g�;V}n+�D���&bz�I�1ٻwgJٍڰr��m݁�.�I!�e�i�m�����'G�n�:8`�TQ(T�+m�v���:)/ ����t������3,����C��$dTb�;b�c�j��S���Ru�����f�F��o,ut�vPiZ-U�]�I���n�$p�=ޓk@$����r�Ē�j�ݺ-'��}��\��de  �I�XV��oEC������� ��x�:n���up��ںN��f���Z$� ��M�$��Үn��/�'���xޝ7@�0}�mhr�Q �v��)4��>��ttp�=�k@:H�Ot���E��-[N�U���@����.����c�|�Rɓ�e�$�:^��"�E靌�4;���#��t�Z��zI����I!�e�i�m���mh��`zI��8`���V��iZi'��{���}�&�������5
J�.`�q.*K���!Go�:P��Ձ��W��j�E�I�ޒn��0��mh�� �߮P�We�Wv�I��;����M��Ix��7@�������C�6v*��΄�[��t's:u/`�k�0�<��6,�nN�q3e�������6�t� ��M�'GW�RK��/�h���tY�v{��������7�ʺ��uj�Rm��I7@��� ���k@��"�7�%K���e�cI��s������}���8s��Ns�j�_�����N�.����wM��� �t��{��w�W��V�(:T�]�]�
N�������o��[��Z8"ث�^ݚ+6�۫B��V�-�@��� ��;�=�o8�p�kK�Tv��Ei;V�۬�7@��� �zd4�&V�'�AZ.�I��s����>��X�$���4��Z���f���>��X�$���Wq"��W��YN���a�}��Pcn�{%��2������ x��C�y�q6�Fv��9 ׳��uƱ#�뮂X��mۋ)����);���i#���'L�i�h}��H��BE��l�c�����9������/Pl+��(x+*���l`y�xς!e��cr�J,p���E�;q�mθ�Y�M�����f!Ǝ�CE,:v�{
�n���vS)���Ӑ��@F۶�8.ݭۓ�C�˭���ߝ�{��v_��6H�3���j��1��o�;:,��[�6ᰄ��٪;9��bN��ٓ�?~~~]��d���c�~�.s�?M�����r���$�����P�:e��y��c�w��FB�zGIS� 쩙��ǛZXG����Q��?�@���=��;�BC��Jݥ�h_�X�:n��s����hu�U�%�B�ؒWm��7@��� �zd4��,T(%�E�t�W^e�W<[=8���˛����2���\��Ľ��ݜ�j��h��:I7����vC@��"�=�M�:�]2����kF�[�W���>����B,I2�IfMP���~���8{����:˼-:
v��y����E�{���{��{�d4�r�h"a���fg����w~�3Ҡ31�4��,}?K��0J��M��r�32��u��>m��5/n��1���۝���r�u�U�\�T�[î�t�`z��{�aw3��l�uӁ.�eX��,���������Ҡ=�t-��$�I� in�R^��n��t��;��hu�RW�V�����fU�ۻ��J�Y��B���[���B)g�`���2zX����f�}[�se�e(G���5�,H���4�$3lH7�h�h�8A���!�G[��l5���( �a�4����8���!���
�)�i���J#�kMfg,��i:lI�������&�>u��"u!��Z�L4�%��4���Ѫ)�ĤL�R�$�JJH�Ya�A[R	c���#���oQou`w Dk0`��֓LN�Mb#��23���l{��՚�iHk��7��;<Q��@��DS�Тx
��	�8>�,('`� �_T}S�	� ?f}�YƁ����w�r�t��:I'������2���n(cn�^��]�Ӷ��i��!�}���t�t��+ �J���F+����ؙ��1��wC�q��n�������	!vNݺ�U�׃����?;�ao0�>��x�I��镀{��hr�R�ۺ�L�b��6��(���� ��i`}�����$�n��U��I��>�L��L������=$��}~���C���n�n��2�� ��n���
1�1�%a
�C� J���'�����U��}�͖�I'bbHwkp�>�tX��t��+ �!�O@eإ"ĕ��յڗ>�#�"�#I�<8lu�.d��Z�7�O]s�U�v��i��ݦ�I&�{�V��!�}~��?]����]ժuv���c�Z�J m�i`z1�h�n�x�J i�t�vfg���LvU ��i`}��5.D{^��Ǵ����de��2��n�a�}~��I�����!�}˕D��`ݤ���}:M�>�p�>���E�*�����$���$lq~r��e����§'mmvC�BY�iÜfU�ۘ�n�]������O��sUdR&��A�"mpjH�W�e�:�:�� �oG,�/Y�<v݂��vf��	Tlq#�[ќ�u��u��]A��s�;kޜtۧb��H��DN7΅^�zr��(���s��(��c�B�yئ.�vyð�wI�d8�\�a�[1������o-kn[��i��c{����}�/`�u�����iWfogkkj�U�um�x{�7Y��û��6�<�˫�V�T�V�p����C@���`{�n���àX�'Mj�;n�w�C@���`t��R^�ж;WhhLI%�h�tXޝ7@��K�=�L���\D"
�ڴ�I]�j���׿X�����,G����I��Ի��]��ZM�����{��� �Ӧ���qRhJ�cnY�9�N\��F�9�p�<k��[hЮŵ퇌�$��M6���Ci��d4���@}��x^�w:�(^kco����5Q��\�8Ͼ�7�b�fb�Ֆ���t��^�d4�r��X]�� ��Xޝ7@�˥���C@��1h�(�EZ�KZ�G/8�f'�W�@g�֖��J����G�1�!+N�+Wn��x��%�{�V��M�>��x���CC�����t�T�/M�:K���x�vg)k�Wn݅�0܆�s���]�LbB�z����+ ���t��^��%�u�!V�դҵgfU��ޮ$�A��ؠ>�;�`}�z��bX�>���i���PvZܒ[��u�P��ϵB�pB�!! G�"�������	d"X������Ĩ$) �&�i�������j+�Ĺʩw�����d������z��:L�b�R�Q�:݋������{�0	]�\Բ�-,���m�<��c�@}��v��e�[�x���A���/mm.�gj��E�t�������w9V�U-v7&ނ�W��<;t2�=�������d���J���_��R��m�9y�>���,�l��Ł�{J�������A������Gb%L̪��v,{*�cw�}�2�{�l-	�LHV�^^��Ƕ�cݻ�7J��|I�ph"(V��H	�H�  �G������:��=�B���i$ҵbn���n�����>�9/@��e`}��r�v1�:�In��[e����p]��Lܞ�y�A1�Z�5�s���v,WW�[�N��Ot�&V��%��L���n����T��U`��0�9/@�t��>�&�tp�%wxJ��%����o^��t��>��٩.%ȏfΔ�;�`{;�����;V�Z
v�`N�t�0�r]��q.(�{j���6$OaJ���g����>�t��8�n�c�3Ҡ>o��b�FbQ~��H�tjW,UY-�}OM�\��i]ۇ7g���B\�8���z��ox]�P�'6d�i6GLgzΣv�8���\�*,#�훷����\�'<�[����x�n.���/F��{i݌�j�g�Ok�gR8�硱D�a;v�z�qc�Gg����.��^b̔��F�`s������۷1��cgPf�F�۩(�\V��Un��dN~ĳl�&��pE��W�@�c\�ڎ��t��Nr\4[�U	���]9���""dGbzL̯�����c�V�woW\�ٻJ��ǤL�Gff{�'�S۪���J�qD�ݻٻJ��ɒ���!]ڴ�iZ�7X�I��n����X�:T��u�s��:��'�ޓ+ ��%��L��$�J�b�'t�Mi:�;������x�����P�
;M~t����x��`�9��Ǐ`������[	֩�m�-
��f�Z�{%��u����{�V�}�X}�K�>��P��J㱑��V���{�9�0��X�)����@^d���J�s��A��l�	��N˖��� ￿�h�}������6N��}~��eݴ�˷vӶ� ��S,{*��v�����nڠ;�?��ؕ�B��*mn��+ ��݁���@f{)��K��r�bg�g��ncsn�9v���OjAs���s�F�@mpX��;��dȫ���m��׷`{�Ҡ3=��/�<ܩ��";*�C�uiZot{�0=｜h�e`'M�$�/�wH�n�;I���{�GUy��p�ר���动P� ���X�������Ϸ�ʺT�^������o+@����:<w`{�YA���!��X�`��{ك�ޣ���U��x�8�������mh��Xj�Z�V�$�*J�Cg����]m���9LY��j�y'\�ѷ;\�6���N�����=�=��t�6�zL������eݴ�˷m6�0��ց�I��t�7@���RI(�<ٳ��];=D
g��36��ڬ���0	'M� �"���i$4$&� �t�ގ��kk��HЀ��'=���U���g��h���V���@�Gt鵠{�e`���u��pJđt]1U�M��C5�v��;72��Y���$q�t���y���;�7e���l�'I6�zL��n�q$�����Ҁz�CK�;U2I2w���`z<�kb{�vfΔ�&ց�. �i$�N�*i� �$�ގ�&ց�G�{��Ռ-������=��N�mh������}}aҬ���X[-�i�m�V�K(�w`g����\�W�%���IC�&/-޺�Z�:V�d�Ӛ�7J�y�3v����X5�L��d:`��4�Onu�8�t޹k:�ߧbȓJ��ݙ��mW]o��Q�:�11!(�����Y���H�k �b�� ����O�	"�d�QD�ԯs1NU��:��9�crVf�,)�����+̓��"�<�wo{�J'*:�f�I�����Bz���F"R�PA��fAn-��-�W�C`1�|��OI.Oe�X]��T'�(�`��ó��Kv�Fv��W�[�t@�b�]f;�`l��Mꡡ��ḍ��@�9�̓�`�@o�± �Ǖ1�#N)�5�����F� ;�ïuѣ���'K�D��Q۫�h|��l�w�Ip��l֭�����K9��%�5�j�ʑ�f��!3$�k��-��ٔ�#&���\�
��e��Hn�,h1%
H�5d���0ƈ�#>��j��3�
t��>W�j]6B۶ͤ�K{[� 5�p��Uv�˪ޘ��=�d�gu佳��:&��j '��!��Y8�E�u�F݅Z��3�܂���IJ3�77f�{;��We�p�n�5=���ـ�)��N��g+��@�m��إx�u�L�^š�����l����S1��v���q��J�#�0i�z65��[x�ݽ���k���u���lv]Σz1�p����j4VN����5�ݞ5������r��9���c������N�۷.q���;.� �uN�r�٩L�v���֝խ�6��y��5lvl��\9�L�B�y�v����������z���4Ҟrs��ѹ��?(}/F61�9j۵�l�l���{r�n���9�Y�]#Q��-�RK�ƛ�B@�;'<�p���0XrM�p�lN���@F�Ԗyv�Q�8U�n���@�rG<��<3��;=%�ɜ6�.����.�����}�(�{p)�����򠚮G����^�m	3���J
:�]V�Ҏl�Y�R�h�sc����{���$�ZX2����)SOO<�O/T����7ΗE^%B��%�n��E�t��=�Q:�8Sq��kp��^�`#9�4T�m�/^աK���eقxm�󰝑9��v�m��w��0F���6����4A�4��"��m&���9���!��F��E�e"�]�@���Om��]�d���mQؚu�ur�%�t�d��cr/l�d�(�"�p�:K�I��j9�ӒY4����[��s͎���ۣ������n��n��b]�9�����y����fY�F�;bG:yt�S�lf�ی�Ƨm�{c\.�9;Z��u��6U�l���u�g�9��T�\�q�Eѝ�0)�P�^E���(]�le�K9�l�@����cdل�]خ;{i	��,��d��c	��V�-�Nwns���h3��1�+�8[�Rsݍ۞�N��R.��ɣW��]s�eթ�N�g<Q��?���A6pG� �< �M ��aV�=\@� س~Y��Fb�����5Z�u�*�[F����JviL�Q��:���Ke��]՞{B]�q[n�"OWc���p�Z�u�Φ��9��Jd��ڼ��:���nWlm<�մ�;�v}k����u`��!q�b�k�:;�=�]��{n�1�x���H۝����I裫��B�f9wb�Ob4�_M�1��toIr�g�\]<�g�nM�c`�Kl\�9b�{���KRKDn�94v����X�������ݏ"�C5�λ�v�2S�m�Wc��!���3?��7vt�m݁���M� �"���i$4$�I@7�݁��q@7�ڰ<�Y_�A��\�WHJ�e��+��@���� ����=9� ���Ў]5i�Cv]��� ����=9� ��n��R^ҽ�,X���B��V��GN����I�k@��J.�K���O ���;�b����G�FuՐa��;�3�c�ݝ���bu�;<U�[o��׷`g��P;V�K(�a��R�Pv\���pv~���,Ƴ�X�BK�p����`y�Py�w��.D� �A��(�{3��3��*�I7@�)/ �zA��ݤ��4Z}�V�:T�m݁��qA���ǿ�V�W�ԏ�U�J�А��wI����~n�`{�Ҡ<� �4����:�t��l��s>p�nJ�=q�`��n�qG	�� c%�ܱ�H��
�n^p�����L�>�t�qq%ˀ��۰1n�;
{���0(R��3fN8��K�D�iPn�݁��qZ��=�t4����vz�(�ښ�ٻJ��ۻ?N~.��Z6Ј?~�?��_~��?��w�<���-q:9V��������� �)�x��!�}�X��T�P��y=�37`}����..㗵��i`��tE֗�*��?�G�&����:�r�@��k�*�ץ+��w�X;7<��i�w���4�L���n��R^;�[c�v��h׉�h��V� ~�۰1��P�7V�EA~�V��&�`��t�����f���+ ��_Et�E���V����������J�������,�ECh��o߷�}U��#I5HE5CM;�OI�ӦVޝ7@�s���˗@���t���Oi�n;,�Y|�f�m;y9.y�vP��gF�n���k�X�Nӡ��f��镀ON��w�K�	ޓ4�_PEj���Dʠ�����\��"��(^�ց��+ �K��-S.է���ot���gI��L��z���J��ۦZ�v��x��f���+ ��M�;�K�;���2����v�LǙ`|ۥ@}�����٘�X�9���!�fO߆��֬��mv�$h.�K�3���"ݸ%ݮ۩�1�k���` f�@qmg=Z����%�+��9��C���̽�bK��i���^�Kl2�Ѻ�[�i��n�������C�:w#G���\�-�NÃ�m�΁�f8�x(���ݸ��Xn�G=�m�"����S����GgqC��UP�r�c��׶��.{{�h�X}%���X�̌skf� ��G�DN��j̵Ӭ�4e����յ���;9�'y;q�:�8R�w�����:��Ts#�����K*������˥�wt��>�e`ߥȮ��eՓ=#���3;�+�K�Dm�ۻJ�����qq%yn�����'��Ӽ�O��&V��7@�]/ �RMyO1�tX[O+@�I��of;�32YA��8���{�i�դ:c��u�owM�;�� ��Z�L�g�_���ݍ�g뱉d�;\�g1���=�����{���e�6s�	���T��$�1!��w8`��k@�I��owM�=W�tE4閙bi3 ��v���8��.s�6�P6���p�;���'v��h��7��}�b�/3٩%Ȍnt�>m� _�n�ut�Z��N�����0�鵠t�+ ��/�!ZV]X�خ���PĖy��|��T����?EXY%��ʉc��.L���z���N�5��m���틌�sG8#��;l�=�t��:I��o�M�:Gg������MұZo+@�&V��M�:G�t�Z��KB��S0��T�1݁��(�r��q�$���K(�S
2C����7{�~룪���r�������ĝ��I2�����1�J�c���`5�u
{*N�HM�� �M���XӺn��L������κ�(e3�L�N����/����Z8�/e�k���F��c7Xqv�ƞց$�XӺn�$�X}�mh|uDT]+V��5m��I&V�t�Z�e`��)hWj���n�[{�I&V�t�Z�e`~��s�uw��RZ��GBWi������w�`n�Ҡ>y��>�\HH�	�RP��hQ8 �>�V��@��)��t�V�a�I&V��;�r��c�X�" R�����]���m�����[�9�����q�$�"V����40�һ%R�؝�hw��s�I0}�!�I&V>�%�Ci�6ƞ�G�t�hI��}��ޤ�J ��.�{*b;=�3��@f=�,ۥ@}����e����
��V��@��I&V��M��qA��8��<�������w�ؕ٘�T�m݁�vwb��s��e`Q�?Ue�ߎUai��c�m9[Uq(S�5��k�M����#Ц�!m�{x�e�ܛ��ut�ыiVÎ��V�Qd6�:�.Wf�Ј�Y/v�.3��ItS�|�p]\�y�[n��Y�Z�kr����k�#��<�n.�j�۰��,�2b�$��j�ۋn�E�3���7S���Ä�n[㣴6.�p�Ɏ��o(ggcon-����Gv�|�.���õ�.�{����O���ݦ��,R�٭vvJ;Sǐ�uaul��v��Ia����u[����a�l�9�� ����z{��πI&V��n���9hLb.��j��w�{��^�$�X�I��K�%T��n:ǔ%J�k^�$�X�I��K�=�}/@><H���n�We[N���t	#���k@�L�N9*%�0V�Slm�$p�=��ڰn�<w`Z���z���L�rVl�9۬��"��I���^��������iӢ�Y�=[�ͷ=��:Z��m���ؠ33)P�ʠ33)P�� �w��սV��9�����τ�QҀ�{*���J����>���ƨ4��V�T�7m������I��{��@�L�x�t�IRBBiX�=�$�+ ����$�X��n���9hTݢںI�v�`y{��$�+ ߺM�$�+ >�Q,�;lT0U��;�ج�c*��ǝ=�GjR�<�Yݣ�$�w �������$V[x�	$��7��t	$��={���Ge;hN�Jʶ�`���e`����I��zq|�\V0v��6&�@�L��{��^y��~�m�M�������{��廅hݣH4Ohp��������6j$6���K��_�������ڏg����-�`�R�u��_��W��75�:�K�b�#sǅ��q;�,0�j�=鼈uBHJ@�BKPUI	����;yg��M?H\����:a֦Nb��mmF�����3�<���O�^���b{��12�Q�15���Ih����2A>o�KRu>jw�UE^�g��^a�w��k���dB B���.��X�)宴x�����z��%�B����<����]�BO�*��c�k>l�(%S_CR�o�|��u��8� �,���WSM����5�ۏ��^^�85��_�K�'ƚ�ĵ6��}0HK����'z4L��
s��:��Ȏu��o"C<*�*�����5�YѰ��w��MV�I������0�6\� k�O<��43TXч9�EA;c{�dy�6\�B�uEs���Av �B�"�Q�=��s�S���A`OAS�H��h�+�$��(�8�[t���݀�8
T4�$ݪI7X߫�����$�X����x��(�ݵ@{ٻ�w�
baL�����	$��7�t	$��7�2�m�~�����[�2�ݹ��̛
y�õk"Ӊ���<�mc<��ق��+�12���݀�t�}���r�$�+ ����1%J�E��M=�$���Ҡ33)P�7w�r ŏb()�EۺV�;N�����;�������I��J����eZt���V��t�����P�..>���i�h A<AK���g*����[
vҷ��e[N�����I��{{�ՠbŋ���Mȿ��&�r�LF���ۡ�X�bf;���эY6�f؂�S����ac�˔�������ՠw�~ՠ{ٔ���W�����`ݘ�(�ew����;2�}��o8�8��7J���wt	�e`}�J���M Ї�h�@_����@{�P�,�의���*&bePj�#�=߬��T������'��BJ�$���>��mҠ=�K({2�cw`Gw�����q��ۄ��3SH=`�a83����\z�3t̝{h9�]v����Ն7�i����ܛʣ�)�{v�/S�;�Z��o&�{&��)�x6�y �wm�ʣǧ&p�s�.KZq<]gD�k�v��Vj�K���vlv ���W�<=��u�m���ڜ����"�����'�͊�o��FQQT�qgӷ;k82sW�eJ� �,���S	5���$�+?]��m�	�1g
��DE+�u�zn\�n�t��h��$x��3�8��^��G3ۻ=��>��*�̥@_ٮ�6�P�pI{���t�E���L�~�.��7J����W���c�1=�JS �{*���v�ct�}����)`q�~ �Wm?�HM��+ ��2��ό~�7@�r��:ui�2�u�{�X����t��{���9����$qȫ�DV��
���{=g3�7;ls��s@%��lR	��.[��ˎK���ց���n��+ ��2����u�j�Պ�[v��wޓz��4�R	2�
���3+ �����O\�T�$]�
���&V�s����oӦ��t����+�j�m:�7�p�>�N��݁�n� �l0�EJlwE��8`����X���f,�Y�Q|����S����R�u�wX�����'��v�NK���ԉ�.uri:K0�؆��g�{����7@��+ ߹� ���I�rTTL�v�?Z{`y�J���Y@{�8P��vP����t$�ݪJ�u�o��ws�঑}V9y��~몿{��U�{���,`;,ok@�0�t�I2���V�^�]r���S�nԔ��݁�������������?�G�1�W��D1�m�;C���B\��[w���t��"��2��ە8W$�Z{�I&V�t��;��l�M�:���7)H��q7\�@����@�8P���mҠX�袨����Wk+@�0��I2�����w��[C�v��m��t���������+��B
!)J�J(&�I
$�.�D4�US����%zQ-�(�m��;OtmҠ/�:T�'
߱݁�%�?��w�p7v��X����q��6+]$���:^Su�qz3�Fp�<X޻-�,�J�=��TfN\K����T��t*�4�V�I��H�k�w`6�*��V���.DBl�G_zIQ�%D�vJ��۰n���t��|`��Z���J��	=�����T�ͥ@fd�@^����*�LUlN�]�N���+ �������m�T�X����RD�v'�UO#;�\�nb��W8����r�~�\�nz�.��v�\T�h냆��0�;g����v��^̹�	v$̤��c�uF��I��Fz��u��B�f�����co�d�=�ps�<n ��kc���*j9�nDɗ.8m�ӆ�۔CZ�p��c���.��Ҏͷ.�N��h�I���0�����٣i7���vٞ!��%�SG������w�Ϻ5����k�2rt�8���v!qٱ�[;yuά���NJ��U2�w]�QU�V�5pnΔ�c���P��* ����ht���4ـl�M�'I��oޙX{���u�[t�v�*����t��*=��<w`5R�ήӡۤ�n���V����N��N�+ �{�@V]۶ӫHC�,�Y@_���@_�,�?8�?�����^�ּ�����b}�W-ܘ��]�C���k��.\�.A�@�ĢI��׷`<n�d���d�@OK��,H��Wn�Z{�N�+�H~ A$N ඉ�.s��8��.O\�@?�������+�~j�bv���u�o��w��oӦ����'�,�0�m6;��tp�7��t	�e`�8`�W�'E�C�SAM6`���2���0�>0�r_��67i�?������{<��aP�TК���R@�N&�HJ�V�m�-[l�COt	�e`�8`�|`����$C)"�����n���0�>0�t�t�X��:�����HC{Z��oӧ]P���i� 5��.�+ ߺe`u�]���ZJ�t1�(���t��*=�� ��P�"�I]�i�:L�~镀g�p�/��K�q<�h�ީ����9ۮe�h1G���=�^��8����V�\M(!6Nڃ"�l�Һdt���r��j�3�8P���t���ʉtw�I��wE��tp�7��t	�e`�L� �뺿.MZC�SAM6`���2���V�όT�:�A�E�m�hi�$�X��+ ���OI�:�.a0PQ�3�D����2��̤�����,���l,B0�P���
B'��{�ϴ	W,럘�i�v��n���V�ό~�7@�L���GE+�W :�3�������<��s���J���Eݣ��6�p;\ONn�S[��s���nY@_���J���Ҡ.#w#��v:D�f;%<w{n�Ҡ>����;��z]D��$R-+N�Zw`6�*��J�����;�=��=��VW�h,X�?����@��8`��M�$镀J���r�%��}��";J���e[�q%����ʒ�מ��S��/�����DU�� �����'����EC���s���((�@ ���
 
@�)���Gw�?�K��9���������~����?���������������?��_��b���. ���������O������UW���AUZ;?��Nc����~�����?����AU^������������!?����'��}�_�?jl��Q������_���ȭ�*��D(�*%*%
$ʉ(��J�B*�R�P
R(�(��*%
$��	*$,(��A ��)
$(���$��ʉ �"J������L��B�0�L�$�)B�B�2�$B�@)*$�P
A*$,(�(�+*$�� �(����B�
$ �B*$$������
@ʉ*�� J�
$
�(� ����H� �B� �Hʉ) �$(�*$�
$� �$��(!! �@�!
2 BJ	,��HJ
���HB���� 	!�!
	!(�
��BB	!��*�
���$��� ����HJ B		 ��� @H��(�J$��@B��!(�J��*�J2��! ������*�@B)!
�� 2��HB �! �!	 B�J��@�BB @�H)!
�� (�H	! ����+	
�HB�2���HJ
2
�
! J$�!*@!"� @ HJB2�(A!�@�H��B�$�� J2� J0���0�H@�!Ȅ!(HH���B@I D� P� /� �I ICH��$A ������$!#(� KHH�1(L�	B !@� D�
�J�g��?�������tUV?�����?��e�_��AU_��s:��������?��?�q���5��"
�����w�����ه�?�DU���U����@�����#;��L��AU_��_s���S�������~ɧ��{�_|�X�,��Y���o��?�U��vdo���9��~0DU������ ������z7E���?�g�{?����s�<�����?�0����*�����������c�;?���{����{���U��z�����g� �������o����~?���(+$�k)h4���0
 ?��d��1+⯰�>�v�J[j�������P P�@
R����0 m�2
N�m��hE| �IJ�@�� [4 Z44h
� P ��@��(� P� v@�+�    -G�P�eTPPA�fT��&��ru�{oz� ���bx �cv=�L�Gp=�4x�=t/-N@ m�j�6��S�תk�U��=�pZ�,�������Ѭ���ws�櫰�b��y�w� to�z	 2k@�2�3� �|P���)J^X l�(l ���
�tR�n�@u� �(�뢗 i� ���  ��  ��h \��l� :\�Fl���
P6e ���k� �`Kw :��)E��   �G� *��J١J�N�)F�r�y��z7{��3��K�����͞�!簹����G�m�t��y�=�  �;oy���Pyxf�M'a����{��G�)x���v<��i�u�p  {����u��@ �
�;w=��On��Aj$��w���9����>���b�G#\ �C�s`;�@��K6��ǈqr�� �]���1w��=��C����  �>��R�4��Jhk�h�T�t9��76��<�ۋ�{��-:<k �N��r�ƕ�ROK����3��   U��9{�g�4����{�z�N�([��n�^��ãs��      ���6�)S@  "{J���T   ���=T���  	�j{MTLR�  ���T��)P  Ԥ�� �OQ>;��C����ן�5'�a�����_���w�ʀ���QT�ʀ����*��PU����y�?���R~�X���1��/�M�����Ф�ݤ��8��r;'��a��Ƨ�����Ԗڢ���2��J꠬�2�����T�d9��I�/����焮h�BGl0��fi\��3P�@���k7�0�!�܏!�FY���᎘a]�t䐤3X�7�4�Ce98�F��!3[8������T��Y��uU���\Y�E:A�YU�l�Y�]�\-��O�������{��U�]o[w��r�'55�Ѧy��p�>�4K���bA��V�7K��
h!t�3DK�7��s�wϫ!��275��k�]M��n��M�><�)f��!
��$	������50��l30r��K
#)�����Rr�JK)�z����!�!*F��K0�'���a���Z߰���S avp7d/���I$�<��޹�	Cq����o	�	����A$��xY��?�6U�<�����g���A���(�Ϊ6�G>��g#�[���Ɇ3L�[����$Zs����6f�8��wo�|��Δ��[��O�jr��oD���+�l9��{��U�V�>,�5\��_=�m���*�~{��ܷ�3b�ަ�r�!p�B��\͓y�3~l�
k�����k^?}�=��ci�V���߾���&P!K��ILHGE�v�Ӿ|wu^���];|˻�̪\�YMe�v��s�y��9Ҳ�u��(U�޾���z�l���FӞ�9봃NH�)[��3�j�X�;Ok++0+╼��kyH/w��\�r�2���J۬����ߍ����{��ٸ�5����k�,)O5�kK�$�����aX�=f��xr/�c}3����v��)�x��ګ��}\y�k�K�Y��1$��{��vO$L��/�����H}��;tU��bF�ͫj�m
�t��q��)4xq�$Wm�5�B���<��9��/5$���FI|�۰�"�;#YsE��M�.D�kr&{y|}I�j(}5�A��h�y6nFBf=�&s��0��B��ω!��d=��p�`�桉@���H�f���t�9i�RZ��	�=��L9�K	d	M�.5��B��]	$2��vy$��d��<'��xK��m�x� �E�.oe����o��.��.�����5�l��&��HT���G!dÃ�!��BjJ6���hƞ����y��'�e-�o˯>%�mhEk\4��h(��3F�)1ӳ���.:)��!��a�a�jӗd85BZC�Rp�8��he�\OOJ�Fa�F�T�5�3[�a�np�0��B���4Ɠ�Y����e�<
B��4f&�����af�.�{�*���b��R��e
�7����Nb�p�7�^{��C����p7y��y��3[�毞s���k\��`J��B��称w鹽�ۣG��B��g޼=׾a�)��7R�A}vz�|ԡ`F`K����L��&��H��<�@�6��ᢰ�ԑ�ӑ0����! ��֣Z���B�$J2B�dIV�¸)����$i��F毆T�e8sQ�J�$*��aX᱔Ą���8M�����|<#~�-�����y���\�vb�๿yޒ�^�.o�/��~!}4x�'=='�6H��L����!sL������75�/),#��#>�<&xr��r�)IƐ"I GЖf��k�׋���yJ�J#�����}b�;��
�3�;���N������+��ڼ�q��
j�Q�$��.���F��f�5�HF�l�����C�G�n�r�R�owJ�y���w�&V�U_�ڷ�kXk^�SgH��VA�xxFB\M��yH���!]�4��c�\ۚb�![y�|S���9WMq IP|^,����[�}�wW���\U5K�v��3��S��G/�>VaXZL	Ys��!&��'�pл��Y3�dڿ}zC��/�L�`�;&k�m����_��iT�[��
��*�t^s�^K�wn�w␞t��g�ҷ�)WE��yFf�W)�;��ͭ�]�:��tR�ΔT�WJ5�T���a]������3�>�j�����ׄ�һUu�����>u+Tp�/�y��M�Ͽa���O8^�_
��f����3I1�c�SRR���.�+��ֳ�>���
W�=��>r���|B}�<J�f�99��lǑ��Hhٿ<���8Kﲚ焹�Og��H����o�'�y<���z���Yb��>>!s[�7���1�H�2�$��3^��g	�0�^'$4l!L4l�
&B6p�2��7�0���dn�
�Ñ�+4�a��7�r�~͞�;|t�<�4��j�^zh���	��)�ɗ����xnmV�\u�|��_gk(W������y��0���=���\�B�e$�ߗܓ������d���,�| D�L5�$)�I���a�&����l��CN!$)�2kA��R��+%<�>�������a���S5�Y��X����IZJR�Y`IJ)Yj��l�������]Fl��8@�
��$$%F���[��.ﵼ�����e��AMש�ŀ�0�D������<|/�����������$M$k�2�0V:|>����C٣I.a	��|�|)���}�9�3g!��0�l*B��� C%����n���s��D���>xF�XF�n'�Mӕ%V�����|hס�q��r}�sSG9l�����A��"�7)���Iy<8i�ML��3^�>ֶp��ב��g�xnSr�_r{��җ�/�t� ��.ꮕ��L8��=�J��ߞ�/�7���,+f�P�fhf�Lnhd����|��_0���I
��@�
��K��ټ�>��]f]�P��kS5�������w����X(�+~��p}}�o�w�=�v�������o��'�o)� /��߰(}����'0.K�]1dp20�!a3�HyCA�=�٢D��Է%Ng���_�W,����33���c.���rkW%4�����f�לp�jrIV]�
[�{g5����uc�x���J_�����	>��8y�!���>��PaHϝ2��T0��N}�ِ�n�z{R0$����D�	�4C�Y$<$�k�ρC�rIS�8h��|��!�B���UyR��E�>�j���=���Gy���ґ�!O&�H@%�)��L�e����iCӇ�禤$��׿}L�9%RK�ꏂ<`��Ᵹ�8��vݭ^l�9��!}&]{�	s!�r_e���) ���|�xK��o���Z�J�|��m�ǥ�'~�u~�/����P�$	2 H�h��(��I=�|�W�a�\d�CՍ0�J�0!q�3ni�r$�3\���j�}�7y�D�B��8d	
ῲs���o_F��K� }e߇��Ӄ��¥9�J-��{���%t}�G�CW����u�<X�r�OJ{�y��K幭1���]��Rs��3\����
��|J�9�,��+���R�e��UWt������=�Bj�7�M����������"�߇2�g�7�����ꯝO�7��U�E�b��{��9>�en�7B�J��ۻp�H��j{�)��=͸y��Ͷ��ޜ�R�&�]�Ho~q�^g��A.k�nXs30�\ONy3�'��%�!pפ.�<�3���eP��\������L�df��Y�m#�n),��|�x[�Ko~�ǝ'����V�ӎ��_a6�u^s��+)��Tg/���K���[F[��D�����<�&�����gָ�~;9ˮ�y"�}���G/o�	�u>�_2��
T��u�
6ov�`����H�0���k�
1k��8���<���8i׳����H�J9mޮf��h|;"ClZ1��d���>8C.�,�8P�%��R����S�I|�h��y�ק���)�
a���6�[��a����.].j\�5�<���G��C�Y)4�����ghl��f��<��.�0�#0�I�fM��Z�wɗ�8�!3Y��8@�/�a�^JĄ����:�3^$"\	�F�dp�5������T���훺���/�5����嘼��̾��y�I`B�W~�W��Wv�u�^}w9޾���=�Kh<֩��Y������sF�h&�M1���
�$���+��,с�)�&��\�Xmb�5)�e�ĳB���7�7���ٛ�BJ��»_#rn�C4f�a����I-	-�ߙ5�N�ߺ�ī�T���	�j��y]N�E�WR��(�>15��%�I�:��:{.�yB̺R�9�No~���'�	��.Y��)a�+24��Å�u��$���lÚ1l�ߎ[7�hzh�[���,.�G^;QÚ�^���}��zo����z��%�k|6��a��טWЙ4��o���O����m4\�r��;�Q��L��=穙|�P�-m�=�s9�ٽ燏�xm&��!�%�ja�-��T9X�H��{�vE�S[)��c뿊���37��B�����(�r�R�Pq/�I�&��r�oy�,%��J�2{��u�ֶy���SN��w~��L��|�T_+Y&��yH�e��m�4N{:���k���	C�P�{�y�d�&���u�<��n `Wo;�鸕"���>�[�wJ���Ze})��׬�6q!�� �V��ә�|�y�kG��y�k%�}����%�k�,j��b&1��<eao������9�ș���{�{\t)�S�����L����7Ẓ�3ٚ��$H��c� ��'��������p��y���WTR>X9��!��9�(��JD)LВ�h+��sF�i�g0<Hf�w��$sͅR7�BRa*K��K�3=�|7́�*F�_7����N$R��.�\u��9痛=�	Ln��IL�B�B�׿z����c���w��_3N��I:H@�����뜧����[!�L#SCo6ˍ���s[��]�<�f���X�ַ��5�]o��kw<�aL	Bk��ɇ<��t��0$7O9=IN3��{�/}��}��B\����׻�L�6�z�2�π�č����6cu dXJce؀FY�J%��<��h�R�[��n�J�X��٢�!R�)��i54a2��IE��@#!ye��% )PWkw�nb�)"��TP�t*����?s�����^�\HO|����6x0��d���G	H1�C.y�~��`S	\	I,�KK&\M�!R6��q�����n���fCs+������9ʫ�3>[EU�7�w(*�>�Ue��)=�#�[�E��b��3e��R��;�[��iS��eQ�D��%��s~j���		!�RH�!��ڧ���^T����2]U����ڻ�����   -� �h  h�      -��� ��  m�  � ���<       �{��x        �     �   ���     !� : 6�   ��l  �h$         jٶ�Ҷ�-�+(�O3ѳMW]WQ�v�ɺ�Hk�����[�j�ƻQ���_S8����	�WCˉ�ܙn�]���r�Pl <��УP�g�.m�殪��Z�ۂYҚD9�C�LtkӮͶ�8`5i�  �:�{c���U2���]A�Z
ZU��U�۱���P�&��P ���ٖ�z�کV�<-P!+��n(Un�H;m�$[Cm�9E
�t[UUUUuF���  V����A��m[@ח�� $ڶ%��%�����b(E�y�HJ�U�$ Y�gc����]w8�]�Cv�֤�  �T�[Q������mWU@P�V����������ʷUb��^+���&
#`����]�*�
�q�B�.���g�yh *ݺ�l��[U�*���]��+�*Bq�mR�J��z�[l+UU;Ö���/v�U[UT�aI�Z��(͘
��N���6���T@!;UUUmJ�K�&v�r;Ŵ9������)m����P٣`���]����ڥP(+��k���U(�-�"9�/�DW	�<^̲�]��`,��T\�f�j�9��uҿ|�v�X�y�4�F�\�n�i�יUۗS���J-�jU_��`u2��om���;F@M@(͆T-����mb9�	E\�(�pm �l{,��iғ=���c Fef�\'g��.yD6_��m溝%L�O23;=��N����7M��Ù�� k������g��ص�v�N��Qʛ�j�>a��&���U��Tj�5T�-N��{���mT��r��4+mT�V�ձUT`��#q�_�k[�
�]U�y٥���mO.ґ�"��]m�y���k�����
孌�ʠ�u� 5mj��-�B�╔�5PJ�cb������G@d����oRlⱪ�(�[$[UU�R�j;��lU��uU�Gh���� o6ݰcrܶ�d�����40R�36+�h���m�� XŵU]ThW��R��UUu��s�}n�b|ck-� $E��κ��{M��MUUT m�uU^���'fU�n�vGq�M	ťM�=������&yZ����e�on��;�eKm<a�HI�u�����һ*�����E�AU������TS�*�bE�ڂ�[�7f
V^w%�g�UF�l����H�'�c[�;\�D3�\��eB&��
8A�
�I�>C�lQev��Gd6�7W�U�H;]���q([��;7J�y�P����!ٳ���<�k��=k�wH�n��i*<�t5��[ csg���=l�g��':^&���t7@+�{U�k�r�tm\S�d�Nxꨘ�+m��}gt�L��C�qڶk;"8�p�,�[[��.��Z�;/m��C�xРrḠ� ]���h���լ=<��#bJ�aڪ����N�뱀�[��q=���G�j�e��K�NL���:\�n�eḎn�>N�����Px��R�kjl��
��T��Uts�M���k����8���!m�PcmJ�v�-���V�*����g6�fz���H3m�m0S[m�,*ѱN��ꪩWj8�Yk�2�z�ST�l��NR@C����*V)Q5�WU�m��6�ʄX\�[����"1�4�95K �-l�*��mr���ޣH;u�D"D�X��P��wh7Vö�4���͆� 9�v����UU����U���"հ�\
�aNG�E)-�PT*�+����uê6�`뷴�R��ʲdsȪ�rJ���
��]UT���|Ϯ��N.�TP�O=*���@!�s����m�V�s�����@+*޺�q�#nz�(�*y��@U{U��<)+�� *�nnr�:�$�S���j�u���cr/j�������7��.!m�;z�7@P!Z�R�/JKN�l��UQB�B]#n2�v�͢�[V, %�BB�خ� b��q�feZ�M�u�&����]V�8���`-��%�
yM����v]!v3�,nG��=5Um�N�,�,;�x"ĠPv-����"Y�eؘ�nޯk�ԭ�u�W]A 2��7u����x�c���K��
���0eP)f�ܴj.��3ֱ��늋r��q�d�BMWY������0V�uh�h|����d��ܻW.�-�)B���TK�l��U���Z�A;��L�V 2�[��;fS0�ωxC횩]�]ty���y��7;�@t�%&��	v8��-�U�l�UJ����ZDt�[R�Ϋ�rEVqsT9jy^]�(�fV|��l�MUK��� ڨK�/i�۳M�h��H��=MVQ���z�8�MU�J��X�����!UoV�[U:�Z�� UF�٪�c�Kjt�v��5V�;4!��@�v��]qU*�Į��SU6(q�l̜]ەU�������j0S(��l��i�Dt�������[�UR/SK�Ӻo8L5.�p7+K�؝XWE[URg�@�n�C�۾�]��
�#Hs3�k��\: �#�;h�t���T�L�XM��'�j�Xw3T���j�[uR���:
g�fX�Y`��9A�e ��V�cm��q��rTL��H�R�Uq���LV��j��i���A�)�)�8�W��)" �C+��PHGEm�.��V��J&p�T�.����� �N�!���`;vgG	L�4�iY%��T<�tv�cZP�ى�"��NΑ	u7X��yR$�y^���< ���hE B F��V{�ض�Ezr�l�DԮ���5lE�Η��{@��f��Z`($Ŕ���U4٥�lEG&�꣄���*��vڕ�x,�ZL#Z�0�]��;(m5U�c7����ؚ��� z:���qO!n�4����F���:&�c�U��:8ĭ�����6�2L�'ft2�+��$Nz�,<��%��]��B���Uɳ�6�m�ҭ�\�P �V����<r�U*�;�v��p���h)Ӱ��	��q4��JNm5(��2:�3�.ջ[�V���5ΐj���kiWvi�6�8�N1pM.�..7plV5ƿۇ8P�71�㑔X+<��m\:Rz�����j�ۅx+/A���&m�i6ц���ZY�v�k��#ۖi�n����wcґd�㙠��5���:Q�9{c6�^bb��qI��o2�n4���r�T���� ��bu���/���K�*R8�a��2i�cKb4��0.�K�r���MY�me��z�UA�Ճ��oE�qq�e����N���eZ�K��N0�\dT$
�A0�ԙj�UX�����U��*�U�f�-Λ [�U��p(���6���L�K�֬m�`9�NƫRry�"˷�鎠+e�\�Um��v��]aq�'F"��
������T�n��m��샂1����*�j�{g�k��K�UF�{,˻.���e��Ғ�ÖWљ66 ��j����\L��J:�F�l�q���UUWT�ԡ+\9e�8a�Mj:��J	5/E�8$���1���=e��ޮ��]��ݜ
��F@�M�Z�`���Ĳ٣P����m�[/ڏ@�fvjB��j�T���j���|GC,	c�m]�M
#��T$J�]]Q��UR��UWmJ�V57��7V/	�Tӫ4�W>�WmUѻ:D�*�z�U\�@ :N���BE��ڮ��PȇVP�s�˰�R�ƍ��`
ڪ�M����v�r�)�UP�Pe�:v �?_sy�����F���Ӈ���k� %ZU�$��ݘ�v�&��YV۶�w$�Y�4*�Uj� ��AT��l��Pm�iہM���m�[e�nU�l�*�[���n�SR�v�5q��%�۶�, @UpUU��Wf���8��r���y[Q��i	�gq��a��EZr!s�;�V��z��9��Uګ�꭪��U�y�I��˪���v�E���']���ER� ˴K����@!�YK(.H��-�UsT9T�(^�em�Oo'f]�ny[�%wew\:3g�J�pL�ݷV�;��j�A��]Ek+ZN^V�&;�Uf�t�x�bY���:^��ڦ9�j�Rc����WL�s-�KP#�� � 6�]']��2�ë*Sٛs6��c�ٳ
?|}�pl�O+N�j����PՎm��5OuUe�"ki��^^���l5UAŵ�VQ�*SrA�un�W\R�,��mAPR� ��٥y6w5Kt/]
3�y���+*p�q�\�,EQZrs�a��Z�CʰVi,9j�1Gj�ՌKW=���:���Q��++�]�F���UPS�«\0�UWBP�����+Z�-p�hК�N�-��Xj�g*e�� 6�,r���eG����O=7`�@+���*�FJ6 %(>M�_�,���s��k*򭌸f�c��jUڬ�<p�J�:*�ڀ���v�5�R�QA)Q��ڕٕ�j���ڀ�:��8�gCe� �I6ӄ���C�� ��Z�ͅ9�N�͖���� �i�ԫ]\˱.�R�HMT�Tm��v�Te�֍Q�ud�U[�MQEc���p�+<�V5-q�B�,�kEU���į�#�)	�ڭ��L��Ld�#PH :�I��b����%��b���{����T�����P6�TX`:����?�b� ���� �`�Az�`��E]�X��xx�Dt�1AJ�q<Z
�QX`�P��S��W�`��p! 0BAQ��?AE�ۭ� x�ĉ�}6�-P�@"2h>
"|#�ǈ>'�|A$��������x(�(:~���B�֐D��HV ](�*�������炸@�w��S�c�t��	�(�@���W@�`l�|Sb+��Gh���mG���'��~E��iDxf ��l<0���`	����� �=�hE� lR @ސ~�A_D��h������}~�$"�Fj�Z��_W�P� � ~H8"��\DG��~P� &��I	$#0&�)Hc"�HHH�J�x* ��"�S�=Si�8�'��|'� x���,@�P�"*J�"���(��؈�=�#	 H��/����}�c!�X���
�x�<L��X���M�P 
���􄾢 ��@���TP�����A�E#�TU}Q������5	dX4�H�3%���N0R��h!B"D���X�F����D�"E#\R$F$K��Ϸ�kZԖ�TUUV�6� Z��Y0��`:A� $-��yPA���{TZ-�ӝ]iJ${r�F�-�%rl�mjKH�����)����3.�h��a��ܶ��m�)8�ݳ����9�Ŏ�b:eE؆����g2�0+\lk57O3l9�Z��֝�{�_*뭶vŹ�q��vێ�7idWe�cB�&B�K�����-��͵�4*>
[T]�MH�S)a�f��h�n�.�3EYk��V�G�1�h�E�Z�X �ձ��[��m���H!�F�ώ��[�.6��)�]�ɲg�@$mu���p��6nxIC����Y�&�a�&Ғ�1��4&���B�2�m�������]t�p�cT�jF�X.NN�.�W:ۨ�$L[;��*XѵS����]L%%q�#��0��b.[n��H�.M�@��	خa5 ���f�bQ�ޔ]Ռ;��͌�8�I��5\R���&�Ҵ�3⌎^Ql�8:IW��!e�
�dN�as�J��(��]dy:�����e3�,]��WL6SK�.s�F�Цx�+�u��
��R;��X�nĜe�����V����ܷZ�[�#�&w�۠zŨl(�:�b@�Yq=k�Ey��.Ţ����eP�Ռ��s����s�0`]���*�ѭ����G��U���u��qm
<	�]��;���ŝ7'���5]=5��<����W�2+s�װ!�]d[g��n3�����=���	P�e8�k��$�-�$�m����T=����yE�i���6�1�j{-��v����=��[vm�l-�i{&AsmGywm��ɮum�d-�G�{�̤K�{�fA2�j�-\!c<��QݕT�v�u��˶��ҷ��M�k�1�5�ԡF�2-I��IdGV0�:�j`�xz�m���,�����`'�����F��������,�s�9�2����F��R�M�öf�E�:씛�k�v�0������0��V�X���k��p ��M )T@6�tM
��D�����
�<4�A
~�|�v�q�\a.�'.փ=�Mc]B����z�b[Y�"�`:gW����#��J�)h6Зu�����&Ύ⸭wl[(��&�@��Ҳe!1����[��N��͎�NL��'a�%�v�c�l���s����lPܜps�n;C��9駮|n�z��#�������g6�gn�*F�`���B[�h�TrJ3W%�Co� ����d�d̋���@ݹ�s����^6p��r�^Lq���WKn雱� ��L�_��}U����7n#�n��v�5cl�8�e��mOe`d��'u� �K��J�B��B�� ���X���	�p�8�e��j���
wV���7X���	�p�;�ذ	�ٕ��JQE�0I�M��\0��,{[2������^�w�l�]�o�f��"�����w�å4�XDЦ�K�U���sR-,��&K�ɜ��}����>�|��;#�95� 9�eK�v�m4�m˚��{�����|"8�!bB"�1)귈�d���xv8`�`�l�m:B������� 9�;�{��{֛M�邘��x}�Ӏ{�p�'tp���wg�6�����Ս� �u� ��� ����'z����_�w��t����G�ڞ�CX�d*b�`#)KWJ$A�r���4V��^V�T�?�M��{`�`]�x�p�9�p�9��]�Ai���-���/ ��;��ﾪ���D�G�E�N�iիo ����9�p��הH(B(�e
	d�h�	 	0$X���_W99���:�%�m.7n���[*�l�;�p�'tp�8�%��À{ԝ�9vG5Zܳ�w�ӀqvK�'c�����9SiݥW>���@˞�Bsq�9ۘ��mm�ҨY��,-F3)�.`�Rf�����K�'c�����'tp�$�Z���ՉU��Э�;3�W���X����/ �ި�m*-&�m�{�+ �Mp��}�}�][�^6?:\���ڤӷX*k����f���}7 +�� &� �s��I�	�����um��m�l��h?;���d���{�+ �n�p��߃YE�+c"; �N3ĝ�ǣk��s�Iٝs4pkS$Wl�R���ԓE�6&�vG� �ve`��UWuo�x^��~n�4��g��0�fV��p�8�%��p�9�ʗY˴\ܵ�g �����?�����J���`��X�mlVݺT�ݦ�فﾪ��o}��;��`�̬���I�uq������B�x7\0wfV�5� �����w4�n��3q0�Jr�f��Z~�ܜ�ק�n�������+�!��T�z�����E�laX�:�U�)�����e�G��ɴ���!8z�ܯ����^xȣ]����X΍72'2��z���nn�§�5�<�\g�1�-�#M�]%��n�u�m��v�n�3��.����{c��X�4,�s1�e �l5I����-e Afa3*�&c����O'99�묕58��L0�[��m����Ξ63�Dsv���{�i�v����β��Z ���>�����w����/ �ɕ�s�ʔ��n�!��V�~H����=��V��;�"�
WvU�;���v^&̬��Tٕ�F�Uq�:WjՍ���z�^��+ ��� �6e`]�x�DZacuM�0w\0V���8���n�`�ꪯ�{���s,��m�#���\�c2n.ݹ�l�${c��B�ƽح�z�l�r�N�Y�j��;R{+ ����9��ꪯ�� ��e`�C֋v��]�v�n�.�ٳ���a�B�d��!#HBF��l�JB$��H��S�H�Q�$*��̐"E�XЈA�B�l`�BZXJi�������7�X+veg�"{�Z��7aa`:hV� ������9[�+ 9ݏ �nB��Ub���f��]��Vړ�Xv^���.T���I�w@ݺ�9[����n�`��y8�oK��e2�S"%66��ͅ�Gr]���a���ښ}sӺ�Ǯ��W@��$R��E�V� �dx7\0�fV��p�5�	�(uwvX��������2�����*e3*��� �ߞ��}�y82y�#�
/��7=�}��<��}7$�y�Ee۱1�[tճ �n̬ �dx{�{��$��M:t��˺-� 9ݏ ;ݏ �ve`���}�����E�V���'V�ã#�x���2�'GX��Š�bp>jvvv�\����ǀs��r�&V s��܅ZcT˦�M��ٕ������������c�9��J�TRv�t۬��2�������wfVɴS��E*M�]$�`;�[�O<��nI�}�f��!��ax& ��@�=��7$�����jj�wV���� �v<���UvL��;����ݏ 䎮4]�팻QN�sz��y�"1�v�z�}��3�"u�����V�O��vة�i���x7\0i&V sv< ������i�mX�[0i&V s� w�<�� ����V5�s�l3�_~����<���$��6Qs��Հ�[� �dx;�;��8�����*�iS04�m��`ｽ��'�߻��O|��nH�H��E��?'�����K��{)Fԛ�y)�lL�CͮS[m�\ղf�4���:���-&͈,h!�Z�ܨ���N�sf�ݢ�<��Ͷ�[n���Qz�%v��q���0�0�Ķ�[ʅn2ch�5 �c	S�T(mqhkun�\�l������;��[p�n�<����=�_վ��e�mn�L��=�mt��+]�b�ͻXo'=��2��6�]��99/=��s�w�������;#�2�FK��:���9#f���������קUն^�:Ě{jj�7ߗ��.� ���wfVɠ;��$R��E�����/ 7�<�ٕ�s�L�ii(�eZ�t�n�{#�9ݙX;��8������q�tU�n���o �ve`�S+ ����� 9�qYJ�5j�M�i��9ئV�ݗ�������o��豃cu�b������pP �F՘aH3M2
ЦJ�8���c��-�v+V� ����� �ve+꯾��;�^��'��}���`:hV�$��>�[=#! �iO�i똌K��r�Ē��˼I%�{Rܸ�#k�j���?y�� �����$�U�W�$��!�$����T�_'WI��hĒ\�S��$�U�W�$��!�$�u̥�$�ڕ�.��J�e�n�Ē��˼K{2�Iw\�bI.w���]�}�rOs=�]
�+f��ŭu���x�nn�v8�<�m��c�h&���F�gy5�1��1Hƙ۰�>���`���\I%��9\�Iu^�x�J^�R�6������P����u��`������ �\�I%��s��ݣg����V���6�I%���+�I.�د�ʨ�{+bf��f�z^5�׼��7C�y�ߐ���p.kq�	eHO�">�$d�$�r�[�n�h�f��0��޳F�IBP�������͎l�t՛B��1(���6J.���Z�:�\q��qc{�tW[��C����eHBVox}�y��rg�F�;�jMތ�j{I�^�?J�4Na�F�2�ٴs͜��ѯ'fk�9�:^�@��"�Z�N־��ϵ�s��x�w���'��,�r��B��%2�3=^,�m�l7���x\���/*R�ǁ��k,ɞ�
D!�'"|@0������tn�{�#u��̮:�3��I�	n1�8\O}�ަ�I�%��¸0r�)+,/�R&))��D�1����bLL`��M������7�����	҅bDw�{Ƒ6^%���f�����-e-!5��W�B����*�Dxzm
���#���$"�B+,HȄ� /� k�O� c�("��Q9�AJ�*W�}��{:s�%����$�jT��)�V��9�w�sx���@�}�׾�?{�l���E�=�sÜ�ߺMi$��M
��$�ݙ�I~ٞ�8�K��n�}�~=}��������WCɼ��heu.�R4�D`b:�-�x�kfV/��[��H�-���_�/@{%�Ē��������^��?�IO_���4A��d� �ﻹ�`�"�I%�d9Ē�s���g�/��`��<09����}�@��׷�Ϥ��/�KIv{���Kj�\g�IX*t�ݘ��}w=�x�JK~$���|9�n>�D�RLHV4%HH!s���N_ˮ���rn�C������ɛ�`y�i��߿}�߶�RJ_��f$���VbIu�z*Z�nM�`:�!�8�\)%�0��=��[����rd�w��_ᬭY%��I/�޾W8�]�2�I%�d=]���t {>�}��ɜg6�g}�~��F$��2�Iwm�bI.lS��z�׿U��[m�ЌL)z =��ݷ�$�ا+�I.똌I%�{��nȎv�63{����}N���}��K��#IsfC�I-�+Se%t��;lX�K��9\�I{f{��I.�g�r�|�5����ꉑOJ4E�=����JG'my
�^K�ks��G�.y��$i�ҍ��2�.�Ј��������e�Nۚ�,�գ�uŲR@����6�Y�Q�	T�nњ5z�Ů������(g@k�jmp:\��4�t,�=�z7��G�n����f96�%�t���^��kt��sջu��ցvx F�By�Ɍ��~�w��"�fK���.��g[�\ݘAÂi9'rr@�=\����ۣ Oi���0UIX�Z���ܮ)�������d:6Xp��r�']�Il~�bI.l�s�%ݷ��v���}��f��ˀ֑�� ��s�%ݷ�$��S��$�u�F$�?OOe=r�t$�o}�~�>Ӡ��9\��~m�?،I%����q$�d���ˍ�l��Ӡ���;��z/I$��!�$�e�,I%�ړ��iմݖ�M�8�[�b1$����=��Io��X�K��9\�I�
������u� l�����ۑM�Wz{me�fzKE����]�kl��,c��� ��z���%�nIs��+�W�֒���F$��~��l�Θ�o}�~�>ӯ$�~�+����=���9m����f��߷��?3��ʟ�?ӪV6\�k�� {����$�똌K��w����$��߅�$���ZV�R����M�8��rg��I%����$�e�,Iz����{��$����6[�2����@~{׷��>��<�K��\�Im��1$�諭��v��:4q�6�f�l�ơe6	m1c���ai
�,�s�������I�b��Y�+Z��l�I)���bI.wT�s�%��,�6��u���O��l�f�%�ZbI.wT�s����K��1$�g��8�]��N��l{>>;
G3+mE����wy7m�����9v<��E���H�a�J��k��lQ��[A�6!0� pH��j)�
 B%�b$�1F%�U	�$N�y�w�״� ����y����crى/}w��x�K}o�Ē\���s�/}[�߻נ�_y�3�Muu�o}��-�bI/}�v/v�Ԓ���$��!��?��9&�Z��Dt�]#kFhY댗g%e���z;I�hMϮ�p�`?^���}����DxW-? {����<}踒K�2���Io��X�K��1�V�+*�$�s�%��#?W��[�����g�� �����I&��m���Kui�K��ߺ����s�:�$�����Ē���$�*J�%���I����9ė��|��Ē]���s�%��Y�o��D�C�� 1Ҁl��{���<���~����֭�t��M�Is�/��$��L�Ē[=�9Ē��$�}���]y���t�Y2ge�#���e�V5���Ъ��CS�,M����Y���9�,�m\�< ����Ē]ِ�K���v���_+�BSż�f6�v�1�R� ~�޽���9��T�o�$��~�W8��ne,I%���J޲��X�V���W�� �����}����6�����$����s�%63�2���P��Ϳy���ﲇ��u���s�/�}���s�9�,K{�q�Ҵ�j�lg}�~���� I�rrN{��Ԓ�o�X�K��|�q$�~��*�|��Ϧ�m<L��r��V���.٣�ztTX���%�������OFYͶ�p�%죪�ض�|}���R̔ -�e5v�lh7Z@]:}�͝�h���L���6[��ĵ��&a���^'�����3�4�ն�' �nP���zۮ���<!Z�<��k;t��z��sb� �����i	j�5%��#�v� ػlu�H�{ǚ�"ˣ��W��I$��I)^��s�E��h�PM`j�.��ǝ��uA7>�I!�=�f�]��?K�Od4g��n�Io�g�I.�q,I%��W���m�ﺇ@����J�#qT9���	w[�g���K�=|�q$��ʼI%ݙ���m�����(��n: ?l���fVKg����y`j�ω��r��������?��}��um�����9.E��ݞ�V<y��L���)Ӳ۬lp�=�?yp�z�ݙ\ �}��7�Q��D��gcVw�6ƻ- ���ԗ/G�挼q�+�\�u�	�i�g ��X&���7ve`c�;��@ęWlO�m`�/+7�ܣ�
� �2��)�%"�`�@�@*��6��`?}]߾ߪ���w+ ����X6@�n�Z�J�ʻI۬wfV68a佷�,����Vܸ�wE�L�'V6� �0	ۑ`�/+�R���`����j���J��0	��z����pI�lp�7n�;N�0�]<���VNa�ֱ�j��6�1+-�k.p���f��KueM�]�5������n̬lp�W�q���=E���8�3�\�߾�'?��$��~�_�� ��yY��"x���:e]�g ����ww����I	 AYg� �)	}B����Wص�^Vݞ��9����@մ*�cl��}T���,���+ ݓ+�U|��g��x�@ęWlO�m`&�x����'�\����'w =�^���e��I����0.Cii.�ÏGae�̈Yq���»4������N�����j�+*�ݻ|O{+ �0�%������吝�����;��'hI�u�M�ﾪ�����^ w���/�<����䜐/��ﵵ�G ���uOz��e�?W߾���������?��>��w�Z��\]��<�y���o �=��I0;��J�>���WJ����mM���]��ܓ�c�e�͵s�=���p���<���~��~:�~�xɲ����ڶ��v�G��e�n0󨂹��9+��pW��u�ذ�$�����]�g����`[%�&�~���g���vG�b���-�U�fղ^z����z�����&���_$O{�f!�ګT��
�X�O[�;�ea��K������͐�4�J���j�ݼ�}T�ϻ���䟻�_��}������	96�����m�}������rά�{����~S�
}��?O$����ٹ'�������$ZH@'�3g��Q�(�d7p��8q�q6����nd�ϒ	\���a�F1�Hr�'�\Y5��Ĝ�T$&p�3A'.j�hl"�"���l`�`F4���C�g9��c�}�׬����O�I���D�g���� ��/���? �N"菹P}1��nݏ����!�C��p3{��{����s@Y`l�J��@����	���T�8k"4���d��iQ�@ׂ�p�	�w���s	�#�,�
&��M%�q��H�M���"Ϣ�2f¦ތ�]��"ryK`RYF&�'�k͋�"�"���FF撆\!�쐹9�K��KHr�;UT0e@UU�͍m�w�}�� :�����Pi�lk�*���7e�rɢR�Iʝ"h�5��R�
#�v0mG4�% ��(�=�Nn�V��j��qZ㙌��f;����	=x
C{F��ah˻:��.�SZ���������E�ln���MIK�B1�����-�֣	U��r6� 4�Y;e�۫۴�;��p�UF2�z:@x�K�J]��%�Հ.̑@@�Dk<�%|�4S��Ά䎶|�	�rAꂹ�,��1)�u�g5y�#ZcLP�.!�b�bg�)�젚9���y8Q�LNhÎ�sV�;j��@Gg]�7�g�g�y�Ⱥ1ګ�G`�>ֱ	;�eMϗr���Udct��m�=.�TN�tw'W\����m���I!��9�/�����뗋�YSNYq�c������Q�w�]���Ãr���C�C� ��E��U�R�/Il�H��Dt��Yj��v�Udc�[m���<��<n���+���V o
�L��A�B`k᥸Չ��EJ�.(ȝ��s�7;	�,e< �������u���Gd�s���P�7S���/��wZ�F�6$6�N�X���b���M��*f�b��0��9X88��v�<e��yհ�<=�!�Ryq��;�]�Ƴk=�z�!����&�4�V��H&�.��v��"Κ���2n���L�W\�b�:aLLhi�2�H-����q�m�wg`O_}�m�zk�7�MpuoH���e�e��%���õ��r�k,8]�.���q�S[	<���k���K��{vږ��W^mZcL�H�T���<��w�P��Z5����҂k�&m�v��;Er]���:Z.�Z����۫v��Q�;[�r���]�l���j'o2�����a�N��S'�̫�e2��׆����v�4�2��\r���x�vָ�A�����A��J�K@�L�2�v^A�)��㒐ͯR�K.HF���pĵ-�0f`��Z�uu�2�b����w�>����0�A���UW�Dp�A<�D>�*�~s����T��%�U��x���XL]���r ���"��BV�,�.�n�&�:R��y�R�-���T&9�;n3�yko �Z�yk6�1�u�y��fʖ�B&�O.�^�� vۚ�x�<�Ɂ�����8P�=sm� p��Cf�k ;�+���xs��zܙ�=�t/8�<(�0x;g�B���ܣ='8�u�Z��ɜ���\�nuٻ�w''9'�'��}���#,)5��xV��^[n��T�p���f-��eM���A�e�����<�l�]��J��8���e�`�e{��O?��f[wn�ۡ7`�ـrl���W߫�=�߲����dp�O-;����VW �������M�~��_]�ߟ� �����6�w)|������W���� ��`�1���$�+ �?+JݟX�U��ـrG�}_vOq�O?dp�=��q�1sB��b�1n����s�+]�^���R3�-�.
�����<��!�ev����m��{�n��8~���� y"X�'߿o��r%�bX���?�h�h�l
޹;���/!y=����r��`'iV��m�U��I "� 21X�D��*DiP�S��*�m �9��;�M�"X�%��{�ͧ"X�%���w��ND�Tș����o�. %k�z������������ND�,K��}�ND��,O>���iȖ%�b}�wٴ�Kķ�����\gj
�޹;���/9����fӑ,K��ﻜ6��bX�'�w}�ND�,�1ȟw�?M�wy�^B�}���n�v�(��f�9ı,O=���iȖ%�b���fӑ,K����iȖ%�b{ߺ�����/!y���*�z��̄crq��sùşL��n�v����rI&�R��X9�s:�����b}�wٴ�Kı=����r%�bX�����~b*y"X�'�w�p�r%�bX��?m��WD�a4fMf�ӑ,K����i� �%�b{��iȖ%�by���ND�,K﻾ͧ ��%�b{�f�\�!%�4S)�kSiȖ%�b{��iȖ%�by���ND��z��Q$K�w}�ND�,K߻�ͧ"X�%�߾�'	�W0��M���ӑ,K? �PȞ�����Kı;���6��bX�'�w}�ND�,�U�=�{��BE<��L��-a�kP̷Y�bH$��}��D|��}6��bX�'~�y��Kı<����"X�%����̶�Me�5�\��v�/�S��d��A����Nm�W�����������z���R0��듻�^B���{�ͧ"X�%�߻�m9ı,O>���h�r%�bX�����r%���/'���ڸ]�`P�V����"X�'~�y��ı<����"X�%�߻�ͧ"X�%��{�ͧ/9�H^B���}�K�i�+��r%�bX�}�s�ӑ,K����fӑ,K����fӑ,K���}�\��B����}��.�lۭf��"X�~H���s��r%�bX�~���iȖ%�bw���ND�,ʇ��	A ��`��i�#�@�>��g�"X�%����ng⚄�a4fMf�ӑ,K����fӑ,K��EE��߼6�D�,K���p�r%�bX�����r%�bX�vM���h���R̶�Bnb\Ϙ5���R�e�:��*7N����{�m�,��Ԙ�[�'w����/'��xm9ı,O>���iȖ%�b}�wٱyı,O{��m9ı,N���8M���l�f��"X�%���^��r��DȖ'{��ӑ,K������ND�,K���6���ؖ%��ztɜ2��i̷Y�iȖ%�b}�wٴ�Kı=�wٴ�K�,O{���r%�bX�}�s�ӑ,K���S�ۚ�e%Ԗ�ə���K�,O{��m9ı,O{��m9ı,O>���ӑ,K�>����r%�bX�g��ɩ��̹��V��jm9ı,O{��m9ı,?(�E����6�D�,K����iȖ%�by��iȖ%�ba�Ԟ���)�@�R��f�F�6;��V�u�?�뢐���p����h�;v:��1�&�q����fy�`�������&�u�lY���l\]�k:��\�/��0u�v%�㎻E�I���z���vl��a�V��۴���jP1tx�^�=sq�Ov�u��+ZE���pn��:��v�UY����0��А��\���g��5���I'�ߓ�$�N����ƚ�a�f͙�&����*�k��lOe�F�����������!sӌ&sAu��듻�^B�����]�ND�,K��{��"X�%��{�͊�"X�%��{�ͧ"X�%���=���Vc6�o\��B���~���ӑ,K���fӑ,K����fӑ,K��﷝�NAE�,K���̝&�i0�2eֵ��Kı<�wٴ�Kı=�wٴ�K �,O>�y۴�Kı/�w��r0���/'������3m2��N�� ,O{���r%�bX�}��iȖ%�b_~�u��K�T�<�wٴ�Kı>�缓Vk)5�Rk3Fӑ,K��﷝�ND�,K� Dϻ����D�,K�߷�m9ı,N����r%�bX��ݳWVTq�Єq3��$��`�J<tz��_�M���Gss���]ul��{��������y����yı,K���kiȖ%�by��iȖ%�bw����ND�,KϾ���'w����/'����e� 2��٩��Kı=�wٴ�7�D�,N����r%�bX�}��WiȖ%�bw��iȟ�"�����ծv�`P�V����/!y,O����ӑ,K����]�"XX�'~��6��bX�'���6��b���}}�]ی;u�³�N�!xX#by���ӑ,K����fӑ,K����fӑ,K�w�6����/!y>�'�K�Z��3k��"X�%��{�ͧ"X�%��{�ͧ"X�%�����"X�%���o��ND�,K�Ӱ0ԅ3&e�:vÂ�ei��#��GJv��*��&�Ι\ʡ��@�7��j�	�2k56��bX�'���6��bX�'��xm9ı,O>�}�؋Ȗ%�by�{�iȖ%������m�/-�f&�+z�����b{����?$T��,O{����r%�bX����ND�,K��}�NE�,K�zvp�չ	u5!n�4m9ı,O>�}��r%�bX�}���r%���U�,@��@v
�%��{�ͧ"X�%��~��"X�%��{������ә��jm9İPϻ�ND�,K���6��bX�'�}�ND�,F���56��bX�'�u>Ι�d�˩2�֮�m9ı,N����r%�bX�/�}�ND�,K�����r%�bX�}���r%�bX��=�~��a������mf)�Ki���5۫:���k��0��Mk��uuA@*�2��Oא�bX�w��m9ı,O;��SiȖ%�by�{�b��bX�'{��o���^B�����7eG\�33�m9ı,O;��SiȂ��bX�w���Kı;��iȖ%�b}����O��T2&D�?~5�'��ɚ5�kS52�Z�ND�,K�߿p�r%�bX��wٴ�K@�,O���6��bX�'��y���Kı>�wm�ɪ�L&��5�iȖ%��bw��fӑ,K����iȖ%�by��8m9İ0�C����"X�%��uۙ��&f��0�kSiȖ%�b}����Kı<�{�6��bX�'���6��bX�'{��m9ı,O�/~����WXeѩ���K�(�a�����K
NgI8�]c+c��X34��Qu�76]I���Z���4m<�bX�'�~�6��bX�'���6��bX�'{��m D�,K�~��"X�%��{�2g&R��.�ֳ.��"X�%���� "%�bw��fӑ,K��߻�iȖ%�by��8m9� �T��,O�ڝ��kY,��h֮h�r%�bX��~���Kı=����r%��X�'��s�ӑ,K�����ӑ,KĽ���PA�
��sz�����I9
���xm9ı,O;���"X�%����"X�%���}�ND�,Ky>��C�j�h��l޹;���/%��{���Kİ@O{�xm9ı,N����r%�bX�{��m9ı,M �H,B(n ��߾����ɱ6��Eq����p��n��"��]6x��C�c[sh���5�<J��ȏ(;��ڌu���뒠bsf��V�m� H���0���I����wv���uM`α����.��ZQ��;r;C�m�[x�ĸ�c&l����2JĆw0	nB�^Ӏެ����Ͱ�M�	 &9�/<��c]c�Լ�����A*9%W}�s�u�.��7*�ü�;�v
�ݝ$��E���z�w;S�͆����O��I"��b�ܨLŹu�M�"X�%���߸m9ı,N����r%�bX�{��lUyı,O;��SiȖ%�bw��:MF�a5��kFӑ,K��{�ͧ"�ؖ%����fӑ,K���56��bX�'���6���*dK�}�ff~�!��0�3Z��r%�bX����M�"X�%��{�jm9��,O~��6��bX�'{��m9ı,O��a��Me&�K5u���K�P�;�{̛ND�,K߾��"X�%���}�ND�,¡C"{���6��bX�'��~'5�3%!�]9��՛ND�,K߾��"X�%�	��}�ND�,Kϻ�ͧ"X�%����Y�N�!y�^C����9�J5������;E��k�][��ޱ5�F�f�b.�	����AL�u)]l�S3�N�!y�^O���ͧ"X�%�����iȖ%�bw�w�l9ı,O>��6��bX�0�Ϯ�5�t)��o\��B���<�_v�9'�:!ťR��f@��p ��N����n�R��
��F6�	E�kw�P�@�,K���Y��Kı;�߸m9ı,N����r -�bX���K�9��Yu.��2�WiȖ%�bw�w�m9ı,O>��6��c� �"~���ӑ,K������Kı:t��Iu�Zh�Ժ՛ND�,KϾ��"X�%���}�ND�,Kϵ�nӑ,K�;�{̛ND�,K�����ud�k%�֍�"X�%���}�ND�,K<�_v�9ı,N���&ӑ,K����iȖ%�cm���SQ1c1,ms�,6ӛ��S�����C(��݇<7�5�9'��&ۆ��m�a�֦ӑ,K���}۴�Kı;�{̛ND�,KϾ���r%�bX��wٴ�Kı>��g�k0�d�$ֵ���Kı;߻�6��bX�'�}�ND�,K���6��bX�'�k�ݧ"~��2r�����{s�Yf�y��z�����b{�p�r%�bX��wٴ�K��Re�|�C:o�7o M��А&Yv|P�Vҁ��O]�YIe�%,���d���B���5��]��f�D��$s�y����ن	x�5�ys͜���`K��9S���ѽ�xjc$8n�є��x�淤6XW�yy��lC��K\�V%2�����y��G+��p��d�k���@1�jZ6�e}]�B!�I+�����c�>o�"S�FkM_q�͞>�XX�А�	�s�aH�Dѻ��
�8�I���0��B�ۋy�8��^kL7B��p��a$�&�G!����zO2��I�aD�q|�����$6s��!&b����,�#P�*D�H��R��Ê$�z�|�ȇ� �X��*��qQ�$�hptE �,M�[��9ı,O����iȖ%����z�o���LY��3�N�!y,AR��{�ͧ"X�%����iȖ%�bw�w�m9ı,O=��6����/!y�߷л	��5!rι;�bX�'���ݧ"X�%�(}�{�6��bX�'���ND�,K���ι;���/!y?{�S}s���qj�0`rB՝d�kr�6����n+����p��I�NcR�7"kY�p�\��B�X�'�w��iȖ%�by����Kı<�{�a�D"�y"X�'�k��ӑ,K��Ӯ��a.��M��Z�iȖ%�by����Kı<�{�iȖ%�by���r%�bX�}��ͧ"(X�%��gv�t�Ʉ�.kFӑ,K����"X�%�����iȖ?�X�dL����rͧ"X�%��{��ӑ,K��{�s2u!�k.d�h�r%�b�by����r%�bX�w��M�"X�%���w�ӑ,K� bdYlN����r%�bX�{ӳ��5�L2�a&��]�"X�%��{�d�r%�bX�y����Kı;��iȖ%�by����r%�bX��>�K�C��j�g��r�����8�(V6�F�*MtV�Ib5�tq������=̳��u|cf���"X�%��{��ӑ,K����fӑ,K���}۰G�,K�����z��������z��Y��&fM�iȖ%�b}��iȖ%�by����r%�bX�{��&ӑ,K����i�%�b_���&j�,�STɬ��r%�bX�}��v��bX�'���ɴ�K K��߻�iȖ%�b}�wٴ�Kı;�d�s�-՗V��.�v��bX�b{�{̛ND�,KϾ��"X�%����fӑ,K���}۴�Kı=:u���Zզ��[�d�r%�bX�}�xm9ı,?0����i�Kı=���9ı,O}���iȖ%�b~P�|��t��s����Vf	�&�.�M�:�{y.y[����W�����>�q�q���\sq��%%sn��"��^*i	[���'��s�.H��N����Xu�2�u�1�ᝮ<���=s]�����ţc��:�-% �,6��%��%ư���inu�#kp,cFCC�0.A��M��^� 8�ٜwt�\��ĳBm5TM��&�	H9�-�D�,�c(��&�\�9�g}�Q�C����T�p�nZ��9�(�q�h�!��y���M�|ۉ��,�h�5�iȖ%�b~����m9ı,O>�ݻND�,K�����9ı,O>��6��bX�'��v���kSY��5u���Kı<�_v�9�,K�����9ı,O>��6��bX�'~��6��ؖ%���;�.��S,�u��ֵv��bX�'}��ɴ�Kı<����r%�� �L�����m9ı,O{���ND�,K�{�8j��$�.����M�"X�%���w�ӑ,K����fӑ,K���}۴�K�lN��y�iȖ%�b|}��.���B�gfu���/!y���u��r%�bX�k�ݧ"X�%��{�d�r%�bX�}���r%�bX������΄�`knTF,�4}������b�'�fw#���mr���w6y�Z9��M�"X�%�����iȖ%�bw���6��bX�'�w�6"X�%���}�ND�,K�}%;�f�.k33D˭]�"X�%��{�d�r/�Ѥ�|A���ˠ|�Ȗ%�����"X�%������r%�bX�}��v��bX�'�N�ö�Z��d���ӑ,K����iȖ%�bw��fӑ,�,O>�ݻND�,K���ͧ"X�%��gv��rB�M�m9Ĳ ,N���n	 �}�v�I�9��f�pI�O>���rwy�^B�{�~��,�i���m9ı,O>�ݻND�,K���ͧ"X�%���w�ӑ,K��{�ͧ"X�%��vHsT�sF�!�5u������# ���l���\~�#���6-zuV����=ev��]-U:��y�^B�����ͧ"X�%���w�ӑ,K��{�ͪ�bX�'�k�ݧ"X�!y?y�݀�1n�<�����/!y�}�xm9ı,N����r%�bX�}��v��bX�'��s�NE[���_~k��N��g\��B�����}�ND�,Kϵ�nӑ,v� ��� F �%pD�v#"dL���ӑ,K����iȅ�/!y��Ś��b�&L޹;�,K���w�iȖ%�by߻�M�"X�%��w�ӑ,KlN���m;���/!y=��N��ŗ#6m�S��bX�'��y���Kİ�~��"X�%���}�ND�,K�uޝrwy�^B�?yz�S Dמ���㍰�m�=���-Z2��yr�K6��94�&��,����[�'��^B����w�ӑ,K��{�ͧ"X�%���f�9ı,O;��SiȖ%�b}�ݳ3�2BS	�W5�iȖ%�bw��fӐı<����r%�bX�g{�kiȖ%�b{����K�/'�7���f�;�^�;���/%���fӑ,K��;��[ND�Fı=����r%�bX���u��K�B�y�^�T�b�KUN�;���V��;��[ND�,K�~��"X�%�{��[ND�,4��j&��{v��bX�'��}���$�.���ֵ��Kı=����r%�bX�^���ӑ,K���w�iȖ%�by��u��"X�%��|^�J�-4#���jn����M7.�N�FV\�HM�FF\/1r�V�RN
��0�s�ι;�,K��{�ͧ"X�%���nӑ,K��;��[��&D�,O~��N�;���/!y'���sU��&fӑ,K���}۴�?�\��,Os����ӑ,K�����iȖ%�bw��fӑ? �ș����u����#6m��\��B����o�ߵ��"X�%��~��"X�%���}�ND�,K�u�nӑ,K�����v�]kV�3%��kiȖ%�%��~��"X�%�߻�ͧ"X�%���o�iȖ%�%��w��[ND�,K���3���Ja4K�Ѵ�Kı;�wٴ�Kİ�����O"X�%���w��iȖ%�by߻�iȖ%�b|�yB0U����#����Y��˯u����.n��7.g�l�E����4�ഐ�=��� ������ۧ2J�Gn�U�vw\�N.|�qgo=V�j�8�y�6uD��ù�)�5;�ڔ�@�(䴃��J�K����ty7��ʉ�v��40؞���юeD��&)4��B$��3�LҶgqj�yqζ�'�߱v5�c��؊*��j�g��8�=cL(Ebɝ��I�rI�N��W�����f�9m��"nq�V�pV6"Ś��J�h���h+±������,�i���MkSiȖ%�bw���6��bX�'����m9ı,O;�xm9ı,N���m9ı,O���u&�L�n�WZ��r%�bX�w_wY��@,K��w�ӑ,K����fӑ,K���}۴�D,K���WE�&atf\�k6��bX�'���6��bX�'���6��bX�'���ͧ"X�%�����ͧ"X�%�ߵ�sR歗D2LѬ�4m9ıD�=�wٴ�Kı>���m9ı,O>���m9İ?��TȞ����"X�%�}?w'��h��u5\�jm9ı,O��}�ND�,Kϵ�u�ND�,K���ND�,K��}�ND���/'��>�C
�Yc�%���W�Ǯx�5ٳ�o-��[�	��^�tKɴþ�wr'?I]���듻�^B�����;�N�X�%��~��"X�%��{�͇�D���2%�bw����r%�bX������).�5M$��fӑ,K��w�Ӑ��"��6(&�ı;��iȖ%�bw��fӑ,K���u�N@ı,N�wd��)�Ja4K�Ѵ�Kı;��iȖ%�b}���r%��"{�_�k6��bX�'����ӑ,K���v��l	�,�e��֦ӑ,KlO��ݻND�,K���m9ı,O;�xm9ıV��{�ͧ"X�%���u~(��\�S�N�!y�^O��{��r%�bX�w���r%�bX��wٴ�Kı>�_v�9ı,C����WA�M�	H�7���i�z�h�..�v��[L=�Ѳ݅k��s�9��E���3Zͧ"X�%��~��"X�%���}�ND�,K�u�nӑ,K���u�ND�,K�j}�ɚ�]�3F�\Ѵ�Kı;��i�
X�%�����iȖ%�by�ﺻND�,K���NEı/�~Ζ��.���Y���Kı>�_v�9ı,O;�����K~�ВX)XF@�b��!��xx �xX�D��}�iȖ%�b~��_^�;���/!y>��o��\�g\\��r%�`���u�u�ND�,K���ND�,K�w}�ND�,K�u�nӑ,K���om�0��MS4f��kWiȖ%�by߻�iȖ%�`���iȖ%�b}���r%�bX�w_wY��Kı/��C����R�i���[�f�L`+ /�]zs7��8�嫆�t�fh�H��e�rwy�^B'~��6��bX�'���ݧ"X�%��u�u��șı=���6��bY�^O}�m�o-ƃ�j�듻�^B������i�~F9"X���k6��bX�'����ӑ,K����fӑ?�95�/'��u�3\���T듸�%�b{�]���r%�bX�w���r%��"~����ND�,K�k��\��B��������H�ř�66\�r%�bX�w���r%�bX�����r%�bX�{��v��bX*�$��!a�U6#�iy"^�w\��B����x��>�m�Zf��"X�%�߻�ͧ"X�%��'~�]��,K�����Y��Kı<����Kı<=;�k3Tն^\va��r�A�F���:Ź�[(]m�y�]�=(�K����W7�N�!y
�'���ݧ"X�%��u�u�ND�,K����,K����fӑ,B���}��}��V�u���N�!xX�'����m9,K��w�ӑ,K����fӑ,K���}۴�O�
eL�bw����5��kS5%ֵ�ND�,K�~��iȖ%�bw��iȖ�%��u�nӑ,K���;�ND�,K���3;���)��5�֍�"X�%�����iȖ%�by�}۴�Kı=�_gsiȖ%�����w�ӑ,K���v�0�#��Y��MkSiȖ%�by�}۴�Kı<���ݧ"X�%���w�ӑ,K���fӑ,K��t�FC�͐�I! B����ۍ�m��dRh��I+�7S�љ�����H@���l�Ff�3)�����1$��!CB,1�J��69D�]���ȵ!`�H�$��u�§|Oq�ŐdVB$�O"@͐N���`�H���!���#!Ia��4'�� ?�JA���#�BD�`FH����C�	@�<�)`�ɢ7N����n�`AY�Ͳ��p!��!1A�E�$B2!f�zMCK�Fp<kx�!�<l!	��4h	$�� KL8f�Ca�I�,
��dIA$����(B�ƒ�mCl�I$�0X%���n���h����{�ff[�k�*��QnQ�c����6�`6� $m�C��`p�\ ��v���W){ubn)t�Nh	1��{[�`���k	1�GRm������R�P7,T�R�B%�ʆo1�ʍ�l����c�"n��n&2@�u9�'��\EACjh�)Cx�*�ݎ�v�gP��k[q�2���G�Ϸ�^r0{*�6�#k����@���#/[Ý�:�A�K�Z;4�tɺ
����9�9��
\�y�S��s(V�����9K0=��Rs��<�>F�N��������jy���Z^�7.݃�|��i�P���ۭ�6��&-�da��ic�Jp��5f=��d����d��	nM5ɮX�D�9̀Y�S�]�a�y��
m���
:W����OYy�i'��r]6�ݸٻ,r��c�g����4��R��� (��e� .ұ�^����@+Q����e���ʆ.�Җw>.ŭV��(�E�vG�{��7E��2���S .����C�xv�Q��k�#WU��v-�.}*/B��̀�4���0��q�cZl8��kR��U�8��]�,�)7���[F:��8�\:�/���;�(񗃵3�67��s �hD̖}�v�s�j�Թ;��i�qv�JM5��Fl���ۇ����9�]'���쐨�P�X"X�7$���f�b	S��,GX��E����\�'�9�]�A�GQv�:����<	7��ˡ��3A�9l`.[����ڞ.s�������G�(i5f�c��|�rc=wk� ��*KƦ�:�0ϙ:
�}�qoM��]K3-�\@Ι5c`�]��Ñ�R�8ٗn٭ug[D��]�Z�z��"�l�3fh�fe(�K�X�T����W{^�h��u��݊��Y��"�ډ۱7�q;i�����A����uŹ�4�J�r�Ť����1/�8���'9ig�7JN�&�^6�a��ѻT���`�ӛ�r�z���Y	o%5�#�B�+�U�n�O~H����x�E������ ��@ODt��C�A������G�t� bV���&��}d�s��N�ٕ�9���F[·�۱<�Ad;��緳�v�1i�K�)-����\��Nn���G3�bϷӌ��\�����9�:A�cc��n޻U�Fp�����ͬ��v�-�v<���9M�x�^{z˷��;d�mwg�{d$^���7��͵�=	c�^]Y8��'mK�=���̜��ɠ��γ����F;4����{9�I�94�$�w����D�:ٻ�� �q7nYg�9Չɮ���+����\��y!�^�f3nK�L�]��,K���}�ͧ"X�%���w�ӑ,K����a�D��DȖ%���w��r%�bX���7�h�,��6�]�����������~�m9ı,O;��v��bX�'��ݻND�,Kߵ�w6���PdL�/'��?��
4�1��'w���K�����Kı<����r%�bX�������Kı>����r%�o!y	���+WM��M\޹;������ͧ"X�%���w6��bX�'���6��bX����fӑ-�/!y=�}t�;(���q�z���X�%���w6��bX�'���6��bX�'��}�ND�,K���ݧ"X�%��߷f�ə,�.3YiL�B(����s����wk6�1nq��\�}����S[�Z�6N�;���/!y?y�_]�"X�%����fӑ,K���}۰�3șı=�����Kı>���Lo�Q��Cf����/!y����fӐ��v� ��ı,Ou��v��bX�'������Kı<�������/!y���v�Kcv�����ӑ,K���}۴�Kı=���WiȖ%�by����r%�bX�����r%�bX�����N�kF�j�9ı,O;�����Kı<���m9ı,N���m9ı,O>}�듻�^B����^��un���5���Kı<���m9ı,N����r%�bX�}��v��bX�'��}��r%�bX���d��Y�Z�٬Dy7azZ��m�fbR<[�y�j�Y"��ny�s*0�Pa4��z�������z{ܬ��;.y`�~k��U}U��������QL��Vp�ݼ��W�I�~k ��6L�)��ěv'I���[Xɲ��������S������ܓ��f䒦�>ʺ-��66�n���6L���/�%�O[�7ǝ]��h�RcBWl�&ɕ�qwe�&�x;� ����nv#f��)mT�yEԌ(�
M.���0$�X�7��>p�;�/]�YT������ݗ�d��s��M�+ ��!]YtJ��]U�� &�O=�$wc�z{�Xv^����+���&���`d���ul����O �آ��$�U�n����}�����`[=x6Jx�բ�>V��&HK��)RFI!$�Җ�HtӚ�$qC&cL�FQ-``Z�H@�XZFB�	�@_������� Wt��!��]��ucn�.�x7`��̬l�X��e_�v�C�Z�|p�JYΝ�ㇲ�t�}�n�1M�Ҍ��V���-�t
�0n#h������;�2�	�e`[%���)e�ҫt���ݙY������߿eaԵ{���I���uw*�&4+�� �&VŲ^�#�xx��V��T�����i�Wcl���{�^ zO �ve`~�^���Y�+�.�U�ӿ��� M�<�n�r���f䜾}�nI��(�=o��Y�kRM<L���QKdƌ��u���IYs�nX���s�S�L�p�Yc��\p��6�]�sz��[�0iM q�S��^(2Ϭ�V|�7��6;[v�a�6zTc�������1k�$�	_GQ�.5�Թ4��M�8�)�e9��tv%��0k�z�ڦ�ц�hM����(�Ֆbd�y0R͝�a�6��l��.1ļS%l�ۛ@Vf��k��n��9��sw{�v��ps�Ee��Ce�c�61���]�֏ Y�m�68�TUQF��hlg܏��r�	�� ����ݰ?{߇�o��W������-�bl�&���$uo�x퇞��{�����aS���11��ڱ���0S���	�#�~�-��;0]U���Uբ�.�}IN���� ��d�T�ZH��V:m
���`���o�� ���}���>��g�F�0�WB&��v�מS�\Q��2�����ذ��ٙqJ�ݳ ���x;�����'�;���8���-���tn�
��r��ټ��.��>�g�ܓ�}��rO��_M�? fOߡ���fY?e�}wn������`�� �엀w��]*ַf����?��<�w����?{��`]��n��ۈ#��N�� �0}�}��z��<<�����Zi�T����)��T�$������u��*,y�;�!+���ֺᙕJ��0�����p�}:��fW������� ���b�0M� Mڏ?U|��=��{|�`���u����k�?�I�5�ʆ�R� ���N�6�UWϊ�K�H�Q�
B�"$c��Da)slLF��V, (�dI�ѥh#$��1R$$ 6"�����x�mG�r�ܫl�I4%v�v8`Se�ݨ�=_UR�3�ݿ*J�|Z��N�]�� �/ &�G�ou� ��;�
Ƭ�n��l����N3�9�۲]oFc�����7��|��1kӪFB�lZ�� ~�g�ou� �����:�z����c�M���m�wM��g�=�~0��� ��~�H�~G�M�]�էM�ـ{|�`]�x$��w\0���Qt�vY�'�������߿~�$���}7'�E`��$#�	RHFD ȡ$z0P �M�p�"�Plmm+�`�� �Jx���l�?����qwe���]�̕�n�&Ѯ]Å��0x�K��&"J�a��.[6�ܼ<��۷=�0:�UO �u� �8`]�~��������ή�V�?�i;�f$p�8���I)��g���#ތ�+=�]���ݍ� ����	$��s��I0b"�S�I�m�������W�wc�I0?W�_.��^�W���Ƶ�×l�p�~zp���߻��I<���ܓ����'ȇ��,$RH�D�1"@��*����@� ���AH�!���b��%{(sT�K���7
Y5���C.�9�ce�Z��g��Y,r;l=���n7>q�]��S7(���<܅1��"l�Ltݧ;<�Ům@��^���l��W&��	�yE�s���v	F-nb71������|�	vP�tsM	��m/n�=��̙+�2V���5s����j�QՈ�g=�+0������s�r�s���h�ำ0u�lc�bh;��m�JGj���70LcM{f�f�V��hM3U?������/ �IW�����~0��V�R:8Y��շ���_���n�wc�I3���G����!���n�/{�x;��� ���������٭�+*�p�~zp	�� ���������z� �uw�I��Iؕ�0	�� ����"�*��~zp�O��b,,1��m�����p��ֻ� lî���u��{��	W_�w��g���2����:�z��J���lp��!+�S�(�xI>��o�:� � @	��V�P6؏T���z�ܓ�w]���~�����_�O��W\�V=Zwc�M�~��.��� ���x��:h*�ա[0	#��ݗ�d�����^�s�����SmS�M7Lv���/ �_W�}��_ ��� ��zp��w�g��n�:XQW�a���t����`��E����պ�7cK��i�~���ShE���n�������H��� �׀�/W����U��vǀsu� �8`[��M��6�ܱ��	�v%v�H�r��ٹ�'��y�7��@I��vf�&MˣU�X�ah��!�Le�h+�������B2ҥ3���
2���ڄB�J\K� n�Q�X��R,�7�CeM��`����B	�64�!u��fE�&͌I5��&M��s%ї	�1 I�6`ŌI��$�1SF3	pi�6]���x���4��竼\Øŉ� FNulu��na��hn0�Nٌ�P� D�\�5��*R	HJM�6J]���R��@�0�@���d�&8D� �$b.% Ú�m�c���c�!H�R��bQ�]�2%�Y�ꐄ�3c� �.� ��d���SQ�i�����b�[XAQ�r�	� �V��I0! 4���D6���`����6��H�q�@�����ä;�=׳X{��j�U)�Cv��m����ۓ׀���n�`nE�B�,�	�x7`�vL��=/�X� ���C�N������A�Z�B�glX�Ʈ�pr��5����\(�Z��q�>]�lW#�����nE�w��`݃�7c��ڡ�CT�U�[0	�"��_U$n���I���p�
�6�6�&&�����;�ذn���p�&܋ ����Ћi]�I6�n���p�&��]���"�DX�F�$4 r_$�y$�����������8�*��<��+ �r,��� &�G��H}���TvѶ�� ^l9���|�^���]v�+;miNZ���4�]�0�;�g �߼���, ��x;�����v%)��\���� M�<��ۑg�着�	��+��;T	�ն��xx;0	�"�;�ذM��[C�+�e���}_.���~��;�ذ=��zJ��$�<ڢ顦
�
ـN܋ ��}[�yp�W����U*��U
@��!k�w�FBP�=aA�d�&�RB#��$����ٶ!śa�kv�`sִ���*\	ѰXB`n�h:����`�*�{=u� ƥ��T�Q��@��[���s�1>�YN��v�)�W�ͼ�;<�ۡ�!�.�iQ��bC�<&Er ��%R�l�1�p�������;=Vmk��Ǫ�x���õҀ���1���d�S��]'at`�b�臧29�nx�v6��4�1�D�_ǽ�ē�[z]�� M
J���r�K-*�#%��Ŵ9T�&�LQ�5�GRqb'Mݵ�n�ŀv��9�2��W�A�y`�#�SnҦ�mВ��n�x;&V;r,��� ��)T��I[eն�wM��X�Ȱ�R[�<��W��#�#4�+��J۬/k���s� &�G�s�e`cV[;]�rm�7�{������׀s�e`�"�:��r�M&[��ڠs����tD7a�vW���9��Iƍ�&F�����:YZk���}:��{ܬv�^������7ny`��V��,.��u���'<����-j�0H'�� ��J{�MNo&,�r, ����m�%C��
��l�'nE�w��`ݨ�v8pޝ�-�[,k�.��~�I/�=��I^x;&V;r,n�L��iS���	+k &�G�s�e`�"�����{;Zi�K1.�[��qL�5s,�ω�[tSCK�GC�����OWE�T�:���iX�C�o ����'nE�r^ŀv��;�;*U�v Ul�u�N܋ 佋 &�G�ove`cV�Je'v;b�n��9/b�	�Q��@��Q�@/�{���>�>��uj��	N�Rh�m� ���ٕ�N܋�����;�?RWi�_�պ���x�fV�諾��\���v��и��;v�Eݥj��ca�t.�-J��J��I���=���5\��А�B�m[�v�X%�X7j<{�+ հ�Щ��4����9/b�	�Q�ݙX�ȳ�_U$M�G��m���wBJ��:�/� 7�;r,��,V�j�*�6��bN���ǀN܋ 佋}��H)P-�6)`����� A�bE�F
��a"�2H������(!$��B���S�_;���w۬�Lѣ-�&�I6�	ۑ`��Xۏ 9ݏ~�''��o������h�Vūe;19�l�la��\^��]���xE3�@����SWm�\�s� �q�;�����~��	�i]]ݞC�T�-[k �q�;#�'nE�w��d��]�/�$���.�J�� ��� ��Lr�� ���x�j��HtӡU�V�;r,��� �q�;#�5F�)�Ҧ�����;�ذ)����3�� 8dO~���au���NM���W"��IˮW %���t�A�š��<�d���4�2Qtl<e�C=�f�yP�c;�
��a�𥕩��G:�p\Yh�秎{.ĸ1���=lv<��LƬC�lR[BX�뜒�4"M΋s4����fm�z7=l��%��4n��	Zƣpu)K"Z�Nz�qr����uĒ<phD807%�6��2Q��
oj�dp�I�U�ww����و�z�˴j4H�n7S�K��+�����6"�Zf��3M��I�6�L�t$����6��9��N܋ �ob�%l����M���ؓ��v8`�"�;�ذ)��ݮ:�ŗ-�8}�����Xۏ �d��	�+�K)��nݶݵ����[�y`R_�����X[%�t�K��*M���qn�x;&V�r,��� �����r����X�Mˋ��Ǎk���u�\p5��7%�q�V��e5�7b�	5���e`�"�;�ذ-ۏ ݍ/Z�
�e&�Yշ�w��u/''	�J��S��g]�X���������wt���v�X;{Żq���.��V�y`on��6�M�[%m`z�]������{{��q`�QNQV���V;e$���̬{{��ŀr��x�����-7O�[p�K�b�ѸqPs��귞(V�1��{���XT�*�����w��׀s��`�6^��������[�WV�v�v���ŀr��x;�+ ��ŀ�ZV�QP��4m����ܓ�{���>Ԁ�#Ӊ`D�F�����B	/{��ܓ�s��Gv�U��Ӥ��w���wg�X۞X;{�RK�&�(Ʃ$]4�Uv&� ݽ� �ob�9JIx��w��w���F�	0�Y�>���s�u
�^�Q3�Ū,]Y���,�	��Ҧ�ڴ��9�ذR�^����7ob�&�ݗ�i[T[$��9JIy���H��e`\��9�س�U�Z~����5�3
�����v�,��� �)%��v@m���f�{��ŀr���2��'� 
H: �aH ƀH.0]
%
��{��7$�y�\>���[-6��X;{�� �u� �������q��eE��$� n]�ou��[�����nR?�<y�j>8U��X�	��Av��^^��9�p�&�ŀs��`�q7Uh��tU�V���6�,��� �G�M�Q�RJ��:]�ـM�� �ob��R]^^��;���9�˻�*c�@��V�X��s� ��������z9�Ir�$۴����J��BG�w�e`ob�;ۑ`O(������鶍e	F�I@��!Fh�x��V�#]�C�ٰ�4¬`kAY>�''��]yq����L�ȓ�����XJi7s0�c hĄ#V�B,#;Ӥ�1�ځ=<y�@b���7Z��,��B�'�B�&�)�7��o������u��w͓4xCEM��OKIISn�����q�h/�qS4ĔR,b�JR�R$0� A�ר�"M�N�	Ͳ�I�}���#������T('5�4� �|'�8�c�t�dB2o{Ȝ $1dCI4����\�L��.O�:��9��ԙ�f�I��Ȭ(Yi ��2���v��-ؙn��{����YwOo�0�#��%IjZ�@ƓAsP��ւs��F�%rs�4B�J�u�+6&��M�vBBc�,a�*�ibI'���׵���cGS~�����C�z:	���{��h�UUңnʰlEUUK��R�T�m��-���Xl �m�]+�sW2HRv�כ�*�l�tn-�� I��]F���X��66*d\l:*tZ���1	�9��On��Ȭ;vm�j{o*��ً��x����ZUgqv�j��ۛV.@��R�:f��V�d"a����X@v%�믖�{GU��D^G���h9�nm,˷cx�1���[�n�5hZ�,dXD��6�wI'g&,h\�/X�2GB�Z�U����W��<�����rY.5ˌV!����,�֩�.XwR����r�L]�
�v[U��2.c����:Z�ѻU,�:x���װv�P�������ûD�j�O�l�ѵ2����9�i�l�Ӟ�3c�@�d�Ko^E���-ܚ�i�^���6�c�s���	m�PŅ��)m%T�!�GB�u�nzUn�j��qT�c����P�ЍqH�)�ϯt�w`CvoG\X뇚0�p��.�c�f�<�R@v��(�:a
\����M�����+��Ŧ9n�m�˴�� qP$�3+�K��@ΗV��.��̰��l6�a�f-e����*%lg]���(�q��̨�q��sm`�Cn]����NȨ��K�؞�şc۵�l���ݸ�e)Z���%���h��m(�N޺���i6:�]��`�v�&u��8�86��k�8=3�+\�z�1	��-cf��΃p�mE>��ظ�t.�q�ld4n'�I��k"m���2-�9۲.�R��ǈn�|I<'q�x{���4���M�v�z�Ƹ�fӭ�Dk�Q�ۙ;H���,l=\˽�-�Km��Z���	��ѥ
v ,\掍�U��KԱ�t�-&��ĝ�t+z�:�ۉ��U�uu���Ez�F�FE�GhݞuM��z�O�"Q�����m�
�"ݑ��F-�v6m%ȋ.6uΪ����1T��k���q���n3�q5��ѩo��E�ֵ%55ur�֣Mf��T�t����)ϗ@���"�< �H�+�P� mc����@R>�/>Ǘ9�I4�2@
��Nz�g��!����Ů!X.��zL�b���7/���]s󳋘�s��"%3/��;m�t�ɍke�+��_MYn�)fR�s�����b�ֹ6�Qq����v*^�����t	����ł��vb�ð���c[���Ɨ��ݰ1,�1뗵��G���n��p%Ԃ���cM��e7jx���Jݳh�h���$��'9ι�N:�-�(Ǖ,U���6��%Ia(7B&�v�s�ö��6:�Ps�vst	p�5�3
�s��~�&%Ȱ��^�������������V�M��$��܋ 9's�=����}�lv�c��W7�w�"�I-��}�޿y`I���TT&*N�]���Kx{&V%Ȱ-w�E�w���o��J��jݼ��+ ��UUW����7o�X�=�V߹'<�ϾE���є��GA�t���`"�AU����J�х4׳�3�8+��v�Uun�pz��w�"�I-��;��V�_���*c�@��V�X�3߮�DG�� #2K���nI�>�f���X���q&ݥm��V� NȞ�ɕ�Ir,��� ��	�]�ucm
�x;&V%Ȱ��, ��<���C��)��Bm�%�X��\������ɕ�{����ae&&KJmW�����c�	Q�gu�S�sA���sS��UWF5�a�-����<�l���^���=�X^�,�'hN�]��l���X�"�;�ذv2YM�_�U��V���s�e`nE��_r�����U_|��_}_W˹{ rl��M�R�CG2�j�uo���$>���o�o~: ��o �d��7�˻�/������6���, ��o �d��&܋ ��Yޭڮ�B�d��m�4�C@�l4�	b�X�	��g����R�J�D�-�����-��Xۑ`u� ���j E�:v6�M��'d��}�UU$z_��H�`���t�'L)��c�6� ��7\0�URG�x����	���"��Z��v�7\0wH�	�2�;�UTU/���惡� �����(�'t'`��;�x�X�Ȱ	���l����4qPh ��^& �թ(�V�j-o�\�z4LJ��wV��ZwW���׌ڿ {}�v�X�p�	�#�7�������͇3�w������ N��ɕ���"B�wg��v��v���, ���vL�w\0	�۲�lVS�o�X;���X�`z����X�y��j��hM���+ �W�g��s� ;��x����ݫm��v��J%���nm�Y̶��T)Kq_;.�,���z<▲m�x4�1���lv{q��+-Œ��]�b�ۤ�[��J'Y��ˡ5�6j$6�_(G�n	e�JcK-+=vW>{D��X�)ȗ=�!j}�s�3�d��l�[cY�V
��9�ID�G�z��+	��#WUш�+f���Rs�A�X��g^M�k˴Bin���M�mFy��W�<87c��3��N"��e���h���n��Лu�7�p�;�ذ{���X$�� SC�V�m6`�p�ݏ �d��9#���F��D�;�;��0wc�9ݙX�p�9�p�9��e[(��];(o �ve`�� �u� &�x��-�*J�n���7X�p�9�p�	�<�{���? x}�;ˬ��)i���	����[(�Khb²:7���8[l��UN�8�ƙ�3��\��{�_� ;�z�wfVɳ+ �{uwJ1�U�����M�'�{��]�F$R,"�#� A	#	a�"� 4(_F����f��߶nI�5� �wY.�իV����x7fV�ɕ���� n�<�u#�[�Uav�Zi��9�2��p��G�Nɕ�e���Z���v� �����	�2��L��mܲ�kE�Ѳ����6�isG�[n�u2h�uk��[�����!D4 ��Z�U8�v<vL�{�+ ���d���_�.����'d��7�2�	���<ld�aWI[-�umݺ�7}�f�{�(#�]tZ�� ` b�{�"�<e��~x'�V;W�]\�-�An�v�`u� 9�<vL���+ ݴ�U�v*�շ�v� ��x�X7fN߾zp�>���v7��0����7���9�#X�f�X8m���\-:�t9\�~��<�.��iӱ�I������9ݙX�p�8����Ԏ�[���Zt�M��ɕ�^���05l���t�ūn��bN�v��v� ���ݗ�rI��s�e`WR�E�Q1Yi�&ف�m�x}�e`������]��[��;���h�Z���'d��9#�7\0[����.*�X��5�0��L@��U�Cۄ��['1ńe�n�_4fU��sh���l���y��7u� ջ/�}��A�{�X�W�/�*E�H����`�e��e`�egꤏK��W�b�ݵ[l�"�׀Nɕ�rGn�`[-Wb�����˾��X}�� ����RO<e���ݺN�
Ӥ�n�lp�7u� ;��;��?��w��4�����KmÃr�)�F�c�%�a�j6�Kʭ2Gh�	bm5���	:�5p�HɄn;ngl�� h�^�y�"�T���2"��㘛�l��;���Sz��b��a��ѱR2���(n_]]ɬU�Y|k<\���B�ok��c���/fx�u����h�dC8���k�1nY�f;-��.���K�n�_��c�����{�H멒����"җ[��8�y��egc5�}F�7`�;t��&{v�Mm`�wn�������ǀrl��}U����'�o�?׫o�>�u����S ;��&V͎�g���$�ׄ�t���P6�����Hᇾ���W�����{ߞ61K��E�l[wn�H�M� ���	$��$��\iR-بn�i��n���y�����r\� �]\-��z�˵�tr������j%U���Ӻ-��4�0�m�ym��]�31[��ǀs�e`��`�`]���M�f4sk��{��r��<�x� b! I��+��G�Y�ry`��`�c��_|���{���;�V�.�7X}s� ��<�6y���ܜ����m�6�vr��$�����?��� �+ 佋 ����,��"ڶ�X����L���,�����t���	��کt��{<��h���תD}q�n!�O-q��U�׸��"�"����m�	?~��9/b�;ۑ`�c�6Y.�]��n�*�wn�Kذ��X����L�����coԗW3\���׀ݏ���ү*�t��Uyg��[��t3S	hk�D"�hI�P�ʚ$��0���{���F-���,�'�FHD�eIP�YI[F f#p�H��n8I��L(&�٪M��8��J�͒H�yF�H+,B�,�������ejK9B�������!$�X�� � �m�����.�3��)�xf�a!$$���F�&�����A�@�$"{�& A0!�iVd B2!B,T� ��	5�$a S&�Ʈ��G��*a�@�ء���X��>}�!�P�=]�UDJ�(��E�}�7$��0	�����v/��WV�k 9��ɕ�su��u�� ���FUۻI6�;���L���{r, ����+۵cb�;e[hX�Ѽ;bё�	�[���f靭��^���`K5�i���u�su� �nE�ݏ��}��' �w��E��1�T���Y�꤂l��7}��\0���J�JQh-�m��ݏ �d���]�~0���͔ԻE?�]�Wt���;�2�Mp�;ۑ`q�G��Q�# ,b�iB	�"H@H�Zƥ1@�׾���f�Yz�2͝��?����=������w�e`n�*�Ui�6���Nқg��lխ&X�m�����C]�CM\V����k�.���=�v, ��x{&V���KUI�/�v�ն��:�����UW�����߲���Y�ꯒ6x�X�m m�1�v� �����̬=�����:�=x�F˷n�ݗi���u�����V n�� �/ �d��9�˻��Suv[���u�� �]�O_ ����|�훒 Bp�0*�����ֵpv&���2[ s ^���T�l��<2ŵ��i��8��������{&�ι1TU��W�����E�]�X��+�KA�v��{�*p�g<��xŵЖ�pj��|�k3�1Y��ŝV�&vN�a���kb9ۍ���������i��q���c��2%�qY�C��n|��طk3�C(�]�4����9�r�[vv+j�V��$��>�8�3t�-;����� W8�i3��M6�4��?�7�R0-#�Qi`-�<3�U�o�� �d��7�2������==M/U��!���m��ɕ�ove`{#�8���6UԴ�|��ҫ����ٕ��|�W�� ݞ��;[W{�s��ˮs8�I-��ߞ���ۀw�2��̬�KUJݫ�ݵt���.�x{�+ �ve`;#�;�jۮ�!GA[�4#��Yhv7dw[�a�;G�t`秥���yL;.�"�j�Z�����+ �ve`{#��A�s� ��N�ڬv�ꣵY�?���ϼ��D���>�K%���rO=�~��y��rp���^�fͮf�98���9��`�X6�,.�Q�`%Rϋv���=_W˱�,w���9�"��G�N�iK�*��.��;�2�mȰ����p�5J��bB%��P�:�t,-��ERv�z;b�Y�	�狭���i�����c	��:����ՀuvK�;��w�2��j��E[wj趚�m`]���U_|��~��7g����Y꯫�:��U�n��nں�ֵ��{�w�rO<�훞=H�FdBd�!$b�0��"�$"��$�?K!I$!H�N�_��+��U
�o� ��z�lWM��6И�M�}��v{��n���8�%�]����%WwiZlwn�`�̬��^��/ �ve`��⑋�y����;q��l>ٝlF��{m�&uXdx}n
A�.��n�/*��'9�9�� uo�xd���+ �ve`u"��*�|[�m��s�"�}��}�Fｕ�n�e`]���}��I�b�*Iݻ�ն��{+ �vea�o�xW߿n����I�Y��;3���<��~��=����'<Ͼ����+�� E ��=��y';������C�,����n����^�܋ �d��;�ذ�a=��3hLf�me�ȍ�����g�6�ɗ�¼��[���E.�R���̒+m����ɕ�w��� ��˱�e&7bc�6��L��ٕ�jݗ�s�"�;���FRwb��ݦ� �ob�6\�W��W�wo�X����v\�ww[W��uwV�X�"�9ۑ`l���}_U-�<�(�*��괩[�V��܋ �U}�Or���� ��,}U⾪�=��e]����j:W��(�P�Q��r�Nn�ye��5c]I� 
=^�R��k;5�oVW��ݎ�'`��q�f�.˷���HYX�lB�B����۶�F|ms��у��2J]
M]�f��+s[X�YG�q��/(����\3	.�&A�u�v�d���͵t[k#$CmQ�'Ob<�"o8�p��:��d[΀�k�,�\Ō�Ig$���NIz�u����M��#n5�Hu���i{+���O���?}�d�O=��`�Ҋ@� �e;����������n�ypz痾�����7o�X��뢘�MӥWc�X{r,��UI�<����;�+ ݫ�V�]�bi[���0	�ذ.�x�̬�ٕ�uM�*vت�v�B��.�x�̬�ٕ�N��>r�e;��&:I��'ve`�̬w\0.�x�����9��GJvp��=en%����{lz�e:&��U�j��0�o
����u�w�2�	�p�8�%��2��v]�혩5��eg �=9��g��H)�T7-��f����7$��~پ��|���`Z���۰V��}��96e`[%��p�7�(�t�ڥwm�ɳ+ ��/ �����y~���p����e��,e�j��z�K�7��ul��rl��=�����.�q�&��I��� �m`[�IK5����0͋]tԫ��M5���31���c�ul��rl��q�[���h�,õm6N���Ͻ�� �d�{���˧v1U�I��ֳrN}��7$���ٹ𚞣1����m���(b��|ꪲ���snE�s��
2��ںl��u�ul��ou� �܋�W�}����X��J���Yl�N˺��&��}�}U��ˀz{�XV�x���g�d�`��y)�ms(��4l��h��3��W�Ԟ<^S�m�v�!�Ӳ� ��/ �&Vղ^68`k.�QI7j�ݷx�2����	�� ��/=_}�RF��^m��t��;u�j���c�ղ^6L��{��J��-��6w ��zp'�߾��>��nN��"b*=�y��s���������v����:�K�&ɕ�wd��&�������y��Q�g�$&^���2%��ʷ"ҍ�IH(f7'��.�����St�����ݓ+ �=�W�U���xvו̥v��vYj��;�eg�=<�`��x6G�v\�wq���;.��u�M�V�x6G�wd��'K��YE����vl�:�K�	�<�&V68`^�ڸP�n�+�n�l� �ɕ�M�VϳrN� HI�"B@cb@aS�c�v��O5A��sXc!(�p��	8�B�iцeF�c�]nQ�H��bĐ��l�aH@�6o{[�U�i�
�Ȅ��K�����)kH&����HQcR}Mi`D�����{�%��R�l�|g���@�6����BEg��ZIM�2�T����C��Y&4L!�E�BD�b��V��6�'7�a������L����F$$$�<�bɰM��6s̀m���Z����Ӆț77	dA)� BE$gw��C�Jf�2d3-�H$�3Dӽ�ѥ F$!tU����bBFɭM̆8CZ�b@�)2R$*kx	�e�j2�w���w�74bu"�`�H���&��/�?� �@��a%������UU)V ��M�������@j�VU��ڨ�}��WmA�U��tZ�,tv�^l�uv�=r����I��;%����]��=p�C>do8̹U���{J���Bv�M1�j��'kn�P�L^]��K|�8B�u40f���e���[=��  i�l諜1���m��f�a��D���I�M\[���2\n[��!9��cA��������[�#k��Wvǜir�Z]8Q�6c��0n��b��V��gLYv����/	����`k�ی`0���ii���6�IAÉ�$F��mI]��A��ZAM��C:1�"��\v���z�-v=gW�k��+��f�Ա.�.�8c���ӑ�$ч����s�piݤ��{\�67G2�������Y{e��mq�|x:z�L��v�g�эX�Yhqf՞7�v�@/=�l
BV���5fBa��cA���G%j� 8���c�C����&�� [���4 \h�_��C$�h�iT�.�%�Lfװ��|r�g[n���TH�ū�02n^��=�����%ݲ�4�p�6�5�Nu��aZ�*��V�M���û0]y���vs�	�<{N�v3�;
NI��\�6l.v3���<�a��r/"�#tX��]ep+w.�;��/s���BEBX3Y�2�fG��KK�w7+�<��8)��u�����r3\��9�>�A�`;�����a"��(ˢ2�p7T�h�Cκ惱v���=���:L�V���Mq�*F�řO &7!f��)q������.G�.es���k��F�aԦ�֩
����*&|7�3[�q��Ԭ�\�Ո�Z�0�E�`�#i.M����!�Z���D���q��{nŗs�v)��i�h�ܛ;"o�k�����-�=b]�H�/\��u���vju�`�9,FwoY4d�������mX,��$j����f�4�#.	r%�r�Pu˥1d�m�t�11�i���P�=E4��D?U�`���$ѡ >U
���#�=�w���-��k4�F{�ٓn(�L�2�lt�1x��ڸ+��]��=��j��Ѵ�#�;u��X`�ʩHl�96���`H�e�b73ʥ��yM�g�{�!e��]�n��\#���a�q�&ղ	^������n]B]aK@���em�L����1lic5�\�b��8䲡��z+��"R.n��_3���sfm�K	��:����ʉ�����I<�p��aU��:Lbv����F:��*`s���G�ë��q�j�f �X��k��������w�0���l� �)��7V;��v��n�	�� ��/ &���p���r���f�ZM]�.������n�&�xv�X�p�lTAҶ۫��v'n�nǀn܋ ��T��v�PV�+�]۲�M�v�X�p�:���v< �n��CV4/^��#����7u�0�QݙW�hY���:wQ]�
V]��.�]�sx}�ӀuI/ &�x��X��gŒ�s&�L�M�9~��߽` m"� ��j��W�Y's����=;3��|��_�����V�R�m� zO<v�,v8`RK�:��H���n�*�wm���`�e`RK���U�ԗ���%/z�֝Վ�ݷwm�vL��Ix7c�7o����Y�f��X�5���:�N��H<�	r�Ǔ����ٮ�ms�h%�]��,v[m��$� ����"��I<��?}��' =��	��U�(�\� M�����_RD��,��e`RKϧ _�b��Ͱl:댽[}=��Փ�~�f��.�� �`�dE�U|�����+�� =���"�R�5H-�����&ɕ�uI/ &��[%���Rϊ�J�C��� ;$x�����>%�� �&V H��R88`���[D�Elq�Z6�.�s쳭ˊY����+L�� �ܫ�	�<v�X���<�����"�WC��ݷ�n܋ ���#�	�%ZR�2�wM��X�p�� M��ۑ`��]D[we��b.ف�K}�< ��x��}w'
5)U�B�������t������(�\� M���"�&��Ixa���U�d��yeS��Ʉ0��u6��=$[�V�sb�q�0�șI�F�ۑ`c��$� �#�"�Sm�-����vN����zu�'9�p/�����y��"�'mK>>�����k �^ sdx{�JK����%�\m���+n�]���l� ݹݽ� �ݰ[.��,�cE]ݶ��� ��ŀl� s~�[�q:�Ci �>��Me�ԤprlM��+�����ɺCK�� jE��ZU�<��Y�5�σ����"ʬo 5\;�$h�ݹ�5�۽v@Q�r�{���jێ'�Ӝ��H7Ly��4�mx
Ү
@�X"��.b�e��ʜl(3i�Υqn�{n�.,��U��=��.B)�o��e�؏en3���JO&M�n�Uu��t1�zLegf鶳E.��=*�'sWSR�C[��y�]�j�&�/%&��U�E�1���R���(.��rC��b�S���ߖ�Ix͑�#��B˨�6���l�M�T���}�WԐv{� ���ݽ�=_W��A��Ey�m�;��lN��g���� ��ŀj�^ݺR]��բ�;,�m�#�ݽ� �$�}�UUR]���<�%�/�lI�v�v��{�Ix͝x��Ӏ}��@�f،�*��˶�r�Y�cj�ꛚ�.E�c3B��y���-�o*�4#����)!�]��^�� 9�<dp�;��`oQ���+wj��x͑�/�U�}U*����\p�;��j�^�ںۗh)�®��x��wu��_W�%����y�U�Q���2�v��ـwu� �$� ����e`�,�%��,v[*ݳ �$���˳�|{���;��{�:�:��!�Ε�6,.���
9��T��'h���#c���*�=����klN��6G�l�+ ���Iy䍗Jz�۫V���շ�O{�Xv�,T���#�"�J]�@6
���m�ݽ� �6^�ꤗ�PUTR--dF��1#�"B+��58�UT3�c�'u� �h*U�A:�I��m�T�x�����su� ��}:�K�K���9� �ߺ���&�`���:��hn�wM+�����Dp{�E���7�� Ŗ��Z|���m��m����Ӏ}��%�����{�j/17V*v�m��7\3�I{޼ �x��j��K�l����_[�`���ݏ �0n�`f�e���e�'n�=�UW�vO<{����_M���{A�$H��A$Y �r�U�T�x�z�srO���٘�Z�+MZm�$��9��j�7 ?��� ﳤ�{���M�of�ۈnAv�Ku��e�ԫ�����4�%�u��v���hLWj��`�p�5l��ݏ �+ �h*U�'WI;��f�d� ��xd�X��,�UW�J��7g�b\�8�ew =��� ��e`�ذRK�;R�n+�|��諻�o �&V��T��=_}�}R�w��?}�;_�Vk�S+8���Ixɱ�$��;Y�����[i�d�92�9�[tڣ�2�s�ƼvY��֛�u�[i���&��sfě4ɴ��v%��q�=�xn���G�::i�:�3��#�A� ����{��YrFXݧ��\�Y�n��6��&lW��i\١�T.�?Ϙ���"��0��%sc���T�i�vv���D�b`�v.���������ú��5�=n6\W"<�����:z�z�.��r���=��ge�1��ñ���d^z�Ϊ�3CAɬX��M�����q{޼ ����e`�p�͢;�v�Ӻl���� rlx�2��`���IhخۡX�ae���L����%�6G�E�)j/�bJ�P۬�|��� ����$� �0	��*S��i�J��M��%�$� �0�p�.���0t��ۍ�f��[#���/�65P�fm���3ȥ�8� �X��#��aKʶ��[����w�� ��ү���)a2kD2ۚ��{~����
�+������D���I�3�${�h���TX�lw�l�� l���2�RK�5D*Ke1��v��ճ 6H�l�X�%�{�[&x����Vڧt�m���&V�Ixw\0d� �n̦ҫ+�U��8T:�g�;=�V���v;��:���*mz���)s�V7XSFl+8׽����� 6H���~0)B��/�bJ�RM��� l���p�5I/ ���.QE���lm��G�s��797�	��!�a$HF0d<���[�O_X�������櫆c�a$>���d$\��q�,�"A�1+��l�����3!Xn�u��K���q!B	J�<��[���H�$��Ϧs�w�0X��s^�.�a��&����������lT=�|ZL�D���٫�|������FlM�H8hd A�I$!-��.$<�2]�͏)m�=LōϾ=����s���.J>iY�w��c�������t�s{_�~����p�K>��<�SHh!���I"4�����FB��ˌ���繻����5��w�>�C�E�<J�y�䓇�34I�Pd	HY$&Vɚ�ٵ7��S�-��e0.|�%I�$�$�5�'5�S�f�*FbA!Cdto��KÃ��$�����!BT�e���sݦȟ.��{��ݟ@��-y\Xc��k����%� �0�R�V�<�/�D5���ICq��᯹��Ą�� �9 y���)s�[y�T�>DCH"a� �~EB��|#�E|�h��<�^v���<�<Q& �����8�~@u�\��ܓ�=��rO�=�0��Wi�j�o �v8`���<��}7'EE�g{�ܓ��_��kI�Z��RV�T���\0RK�9]�� �z��(Yf�VX��$�vs㶼X��zݥ�<�l�Zze6�j��(7m�cl-��;�p�5I/ �v8{︂/{׀v_��]���b�lc�`�K�9]�T���\3�_RA����M�͢�KWpgߟ� ������ ݑ�Se�mӻT����ـuI/ �� n��2�TW�ؿu�rb�:B ȑ �WLF��#zk�y7$�����[�M	]Л����#�9[�T�rI����\j&pV�	���hn���.`�8y��rۗz`�:۷�2�h�E	6RUwV�8'��V��$�UUWvG� ��O�)��+J����x+u�=��}�}I��^��V�y�6�=t� -7EZ����{׀su� ղ^��p�&ը�W(1�m��x��d�S޼{Z�uI/ 丅J�j��+Vʷl�5l��sMp�:���rk��Wܗ���s�<On��Yk��\�M��AE]�^+�8����M�r�dnLΫ���dc�u2��b���&(�ۦ��lx��tp#ft�;U��f��[/�cF��7\�ԛ���ӟ�Z�1��kg�l�M�ћ��k��f^�z���.�^6^�3q�� ����'g�1��5ĳJmh�B����{C����܍4�=tr��Hz��4�-fuOw}9?NrNM����Mm�jh@F�ᇝyڶ먃�ti:��lZ��F�+E�5�^B�j���n�J��uI/ ��V�x�%�7N�RV�WWNـlx&�`M��ok\3��}I��wg�2��]��w���"�/ ��̬ �c�;��	O�M��;�m�Se��fV l��Mp�9+i���ڷ�Wm��6e`͏ ��T�xZHj����ͫq�r�@z^<�N�F-�*r6�^y�=��q�Umå����kJ��w��\0fǀr�fV6��\�ֳY��5����⃴� �� Z$`3���I�o�ܓϧ�l�� 丅J6��+V�� ;$x*l��5l��ou� $ڴ�Wl�v�V�I��r2�[%������^��{�U6�����V�x�`d� �6e`����{��T���X�+FP1V�7k��,Я9N���Ų=����U�ҊWSB�6��-�����`͏ �M�X����0%?�I6RT��ـ6<�6e`�%��p�9*S�)�� �&��9SfV��^��o�W���Dh0C�Z���
��\P˞|�`^�� ����T���j�n�Se���j�/ �I2�	�j ���vӷBm���{���o���;^���{#�9�����;�;W�Ӎ�y����/01]�aup+Y�t\s3�j�p�s�-��eU�]rLܜ�߻�*I��6<wfV N�X�i�m�Z�ě��$�����+ �6^��M�˺�6]�۬ ٱ�ݙX���Tٕ�v\.� �2����ݙX���Tٕ�B�Y"B)�d�!��I#$� �� ,a@��|��^�_w7$�����X�,TՎ�`���?v�=��zz��̬�UR�w�*ڡ]�J�(���'`rg���k�SͲmq�2�32�73*�e��E:�
Uv�V��;[�� �6^�뇫磌�	��we5W뤑Ai�*�
ـj�/ �u� 6lx+����rs���S���Q�ٵ������ ٱ����l��!R��e7Jճ�m��)��v�?���wfV N�X�i��vZ��M���p�$�� �ve`� ����'��$��љ�tRRR��3z�.]D�����\]g�F���4`�tp��ıB˂�eSA5�r��5a�+��;j98�Z�v�/D���Qj����d�hö@�^��Ӽ���&��iU���a�e\A\ApR6��1�)F���
�q�̊�d�`���;�Ϸ�����=/i\��T�/1�P�l'9�5�s�.��Ce����<���:�l1۱$������rrI��䑓�uv��Tj�X�3%  .�s��d��T��B9�F95�S%cX-ݶ؅W`�wM[86�����	6<��p�;.
�e*MQN�i��w�2�M� ��p�$�� �u�JZlb��v� $��	��Kذ	ݙX6���)��RE��v��'k\0	/b�'ve`���*��$PZn��R�`M��N���	6<v�� ��}�u<ۺMXq�ʹ�c������pݺ6;vPg8�A�z4�o5����3�P�K����+ 6lx�k��l�(�JF�"ˮI�g >��y��G�:y<���a�BE�=4�`����;��uz~��fV��b���6�j�T;o �ָ`��`���<Un�mۤ*WM5ut�Wv^ɮ����k��r��K_*v�S��x&�`;#�7��N�����@�f،�W�5�u�Ic����)�Wj9�L�2�S�mÖ����J�b©2���ն*j��p��<{Z�w��`��s��D�v 
��I���k���ŀrk� s�<�֪�:�����![0�\0Mp����Q*0 I��u��$�߷XVВ�\��&m�l�95� 9�<�l��;��E�Hݲ��ճ�v� ���i�+ ��ɯN�<�y��'�`?"��8k\��q�{���8L��W�i�7ֹ��%#�/8�ci���m����V���\0�#�5V�VݺB������u�wve`������X��wW�S�J�����95� ��/ ��̬��+ �u����Vة�f��/ ���X{�+��IU��m�����
TXF��Tqm\RF	2Bi$(�F��["d[���R �x9{��7$��:vژ�V��M��7��+ �ve`��qvK�?}�+�hi�0�WAN��͟.:5��w5�ǒu��:�눲��ul��ۢҠj��b��p[=x&�`Se�︂mOe`��e��'Cm��ឪ��H����j{+ 7�B�#vʶ+M�[�`Se��ٕ�ݏ �� �v�U-��m�M�����Sj{���� ���v^��e�i�]�5ut۬ ��xz�����s�@��&y]ܬ	�TU�PU�uPU� "�U_����EW�_�'��B
�P��T !B
�P�$�P�B��0T"�T (�B*�AP��T"�0T"��T T"��P�!B*���T  AP��B*�U�"���($ ���T �EP�)P�B���T �AP��B(1T"�B T �B(T"$ @T"�B"0T  AP��B����",EB  AP��AP��AP��AP�+B,B*,U
�T"�T"�T"�T"����U��T ��T �AP�!B"�*��T  AP�#B
	P�
�P��T "U��P�*T"��B(!B�U*T"�B�AP��U�@T"�AP�P�0T"0T"T @T"�P�EB0T �T"�B#B �T ��EBB,B
AP�0 AP�1��P��B
T"!P��EB�P�B
T �P�U�T"�P�0T �B�AP���BDB�T"��@T"�P��U)P�B0T"�T$E",��"���@EW�**�TUj�"��PU�ꀊ��TU��"���PU�*����TU}TU�b��L��ʧr��Y� � ���fO� ��~@Rf����� 
#��m;cA-�ٚ�)B�@k-j� 2h�Q��*� QB�x}�Jhh� ( � � A�h � 
 
  �  h�4�  PP4 �Z �   ;IT�ت 6�M �vQv���u�[��{�_w��8�j7���3N��@ջ�`b�m@��W� �j;�����)�^l}�O�>���[��<���=7<�> �ϷA���zy� p �>���5 ��  s�Z�l �ǐ����ݏ����t}i���^�s��S����o��=������w�>��� ���½{���\QG�u��}�����c�5���C�|����4{�z=�7}�|�x �� 
PC�ڰ�8�����}�ϠϾ�(�>{:R��w:R��Ez,�zP�6R���Δ
S��(S����g��K�g�)K��E)K�R�  )��z ��nR����e�8����
R��p�.��R�=��)F�� ��:QJs����r����:R�   Y� z  �- ��6���C���.w:;:QJ��`-���W�Ixf|���C����f�����vk�� �0s��}�;��u�껰zw������-�p��Y\�}��ϳ�{>��x  �>�BZ������0:�����w�W���3��=���Q����41!�������� �z�8   #��:���OxF�t2t�t>vOz�'�������CG���w0�� ?DSmJR�  D�*�%?Sʃ@�3*�i�d�  4�(��* �T�F�Sm*�� h ���ʕ	� ��~��?��:��_�����ק���罞�DD^����DAU� 
*�� ���DAU�qV  ���Ԟ���jM��l���d/����o�������Μ)�9��w����/��R�6��LɭC니�;����B^��s�����r��s�;�$LC#L�|m�#Z@�HFH0�&2�c#��K�!�$��P#IB����,d�c[0��K34˚���$\�J@�)����HR!�)�aaf�8ۚͲ᠄�Yl���#�*���Ǎ�a��CBySS&��	rP��B�f��a(B�� B`J�p�2�+L\I��Ě%I�Vܫ-؞�|����DMB�1EVX��Oʤ�Q>լ�B�es;��_	Ӹ��~ҫ��}�j��j��>(�W>���Vt�k�Mww��a	����ä$>1����̄�
��G�w�y������q�m��~>~Vp������z�bH~���1����,�))�_�}a$!f���2���)dHԄ$aI`V,H��˴����sC��@����ں/3*�㠢��^����3�+��r��]t5r�'yk�CU����^m�sa5�����q�N����[�>Q	>L?��R����rrp�',%�������yƪ�u�V������<�/~4}��^�>����$d�"�����d��{Xf��۪�y���|k.�U��.��W��7��{���3FK���K�H���X\ɭB櫎g��$Xh���%0�\�?�k|	q�3�A��ɼaLxK����Z���q�>�K���e0���˚���ؐ�Tꮪ���AM�iwT��{�;nޗK�U�gh_g�f8�N�g���&}8|��mk��v�q�BO2��w3������J~�?s��}@¤$K�5���2c�e�4h$I��C���BA� ƆC;�?�8hִ��H��Nҟ����5�d���H�>.�@���2�\Շ��s��I�%��7�|�k�I$��H�B9>�����8a��3d�0���믺}�|���o����Cdb�ns���v~7���wm��g>!���s�������R7w�ϳhC��JB�ĩ $Z�p!\CAE�dn$��xB��c���끣x�R�(m#"H� ����"F�1b��F��Iu����=��dR��*@��bF�����a`V�ԶQ/�^~%�^��yR� l.��|h������$�Xh?��ٲc�!p%�eωL�ĕ0鹯�Ү�%�Kw��WM��+Y_	]�+��$xF�+�ߎ�X�hc �6p���K������J�~��.����O�RB`di0͚X�C$��4e���3����?|Nὕ��#N�at_�o�v�3P���I�!��vi&h��L�����a����ӡ.���ו���Yx?�>w9�{�ﶓ��ۆ��4S{ӣA���m�4?~\]�[��~�¤(�$�7�}�}��{u��h���	HV0�`�]����$_�:)��u���}��46�������o�cҤ(�X?�	�Z7��������f�;�h��9��~P�D�j�fr����ko{H��O�/
���q&�l}�� 8Qĩ��Ӽ�>�ʮ����~�'��9���y���~�Ì��ϙ�5Ϥ�ӥڐ$�aH��#���'>n�>&k���O�����)��klE�����t���I��3x�BMxJ����rU4�sX���q��! `�� ���f��*�k7!�&�
�f�b��y0d+����7��˼9��bbѥ�u�o{6d́n�%H�4��
Xj�~���B%�������J�bLҤ�{��}�w�ֳL�7�;��x`�Y/�.y#J�i��;�H����_~?B��|�ύE�7�EZM'~e�ɯ��im-M���xG�/	�~�����{�w�}���aYH�T�p��K5�r�M�T��M����)y������;2���P�O�yh�7��SↃkMG��Lhf]���֚��l`D&�v�e���= �cǩ�c�(0 @������u���ѹ��w��+n�Ska��J#��]8�Н�J�L�l���.k�]n�[!pY\H���7�����9�s_~����h���`��bKD�ZJ�[��C�r����tѦT�o�߻!�7�SGxX������z�ސU�U�}3'2WE*��)�u�o���者������������!�1�t`[��rBƬ�19������~�!m&�
kT��I���YD�t���gw�^�eWq	SڼJ��T$�i���~�5��ZU}�!G�s5�J�G�8�{�٬d3,XȦ2Mˁ�[~&�w9��9�����6��R����0�U�u�8��6��}��H��l��[�qF��oFn�j&��HR�VG��B�mj-�>��L��7>Z��3��ӕ5��������$���\������R��+��vG!�l>Ԝ%��w����_|��w~q]ew��Ӭ��ӎ7�
I�iٶB%pѳk
䆒0۴�Yp��T���|�ur}���S �a���ai7�qcL\
��4arj��7�����g�W>��I�#�"�3H�B�:bD��Ը�f�SB�-&�Oͧ�4���J�:He[��kR�n��樞������	�_\Y񡯓 �c���٭�7n�s_��JϘ38D.�$IrS8k�k]�u��,ۄI�	L�(D��\�F0�
��"����wm.h�{�O߿_�"B?(�~m4��{'�h��g�k5�'��*'�L>o﮵�b��U?g�s�s��ZM���}�\��5�0°��4%�$���ߣ����SC7��i.��W�w�O�^�&����#FC�(l&��k{��`�8����KHI i��������W�xA$)�+�V-`@�\���w���X2^��O���8N�"F���>mcB�S��Ii�X��"�I�2�
���웓����C�����3\�N��]a�ß��\�������~�HG�ie�͖���N�@���1f��b�.����a���g'�>>��s5����$N1� ���?]#܉|�L�L��J���a�3Q�ς�eÁ�!��@��1�&J@�Y,n�o�jo9�}~��>+󠫁X`@���3?h�өMs:	��B@�	F!Hjܭ��ׇ����>��T���=��4}ϧ�`Ħ}��8���R��0�$6�g�bm�;��}�r����r�-��^�_Iϸ�[�9
��f�0�k	��F'MLճƓƢh.�W9��ʶ��_��4�BZM'u��|Z��xK�sgڿ������?H�4��'&V'L�()>
�e�Ww(Z�)w�|����p�6MK������s�w_g>��?0"�˫55��M�ٴ��G�e�!-gĩ�n�$ s��}�g�e���ѣfɒ^�bo�����"�����#�ﱋ�Y��Np��@�8'�Nw�	�o�I��2�!���2���͟��9���z��Ǝl�5����}���3F�)L4M�Jf���f6?,
�6���p���dvB�J?��寧omԒS{
[p4H�%[-1�T�X�q�ā4r�HFd-�eYLa
ccs FB5 Q��"Y$!�0!M�)����Q�]�k37�����LC@a0�C4b��cL�L4�FkLi�(0�c�Ѡ��j��K0ܸM���ޒȚӀ°&`H'�C����a��nB��H��V*�%Rou;�4�ِ�;�<g��'Vj~��:M:���B0;��\a�I6l��s�le�5��3�x������T8s�PQ���[�_ �\a����W?~�>�s����y�?~�d��bS}F:X�b�	V	^�fkcHH�Q��~G��H���	u0�XbJ�0���N����XHo���A� �d	�*�)�
�>S.�4d!���$0�@�q5$k�"2a\t��)��"CԜ41���ˆ��� ��h�sA�1�\2fp��9Bi�uLb�g�qLsW6�h��e���@��#���@�f����q\ک�F�����c��uխnoet|\arD�L$2s�~5s-3�����-�k�J����ӈKIo4����˫�c�Q����_C��Bo�]��4i�
CE)�7D�c����9�U�ޱH��
l8o�Ӝ��3S���sv`q�b|H//{�tU,N��f](M��76�q}7��9���4�I��K�0�Np.��G�����F$9!a3��hĲ�~���~C��NrMh��9�����ĉ����&��l����~.�h�F��CZa3Zmo�9����[´b��2�D�$a�B�Bނ^i7.lѭ�������v��k�.6ɮ-&�U�08o�6B������.@�o�>䚄���q�)�Y��Ba:I�g��a	��'���z5$Y!	c�y��D�ZM"7sM&�/�����������JO�o��
i����L���z��k��5�-ψk��kK2B,&�	:�'MgӐ�;�n\��o�������U �L~?�%��8|��O�h����IF3[��]��"i0Moxq�&s}�����bA�cL������������$�F~w��� �$-kd����ޔ2��>.:C-58萔 ]���4虤�8F��F�%J`�2D�1����Y����s��斜�!B��	��l�c]Mm���KT��O�c$B@���	���R	!:N��
r3�7�	��o�ތ�H]H�kY�)66n���|D�]pֈS4i3�H���b��﷕�In���'��>{�I��l����~HTxԩ��.���O�&���7�K�&>˳�����s{�	`4a`�� ��4��曳4f���sf����, �;5�~��}��s�&�q�bi<Mϐ�'p�9˟k���oW\|&Tl�s�$ΪCa�@s�,��w�w�Rnr[�w/��g�)$+,���&���k��_��?of��RA.h!L���5�O�ÜMg����a!\5��wy4��B�%�5�X���(Jsl���C.�nMl96O��9�W�k04�Li���|7�4[K�*���+�o|�7P�5��MED.h�����h�9���0�l8~ S9 m�!����߹��p%"I7�\�q(��k6��Bh�^�=����UUUPUUWUUUUUT�UUUU)-T�*�UUUU]UUUUUUUUUUUUUUR�UU��
��UUUh��UUUUUUUUUj������������PUUUUV*���
��UU�U�UPUU�UuUUUUUUUU@UUUJ�xs�UU[j������@��܏V����/D����TZ�i�SV�Inġ0*���M�����e������8�	v� ]�cgF���F���UM��HMO���$
��uJ��5,�4ivm �+�J�\��� �*��W
邙��j�ʰ�+��뭹V���Z�����55UTh`�V��*��R�m*jـ�[r�؁��j�j�����U��V�Ij]��j�)�0r^���Pb��U�4X��
���N[8Z$H�(*��m���Q2�{j�� M͘CF!5��b�F�E4*�Y�P��Z��ڪ��`�������.�l/<Ա�UK�!N�թV���@�]*]�h���+��h��i�uTmUT���TUUF��PZ�r�UUU�UUUU�eP*�U�P(��V�5Sk�ک`�j���`Z
���Vm
X����y2uT��z��x{l*��\�:v�ZЂ�W�1t^�����An"L�QA�X�	�p����������]���Ƃ�R�TV�Iv8�W��@mٸ���2�gG��U��8�kj�a�i�*��շ*�p����2�S�M�R��kL�*����v-�U�%ݪ�����U�T
��&F�yf�Gu.�Y`%�ܹeU�j�]����nnj�:\p�[UU@mJ�T�m��M�AUP�pye���kv��7k�����R��Xz�b��Z���*�vڃ�jU�1(h`+��.�U/%���aV�n�^�/[/,��[@mmUU��T���Uqè�� Ҳ��_�jP������jڨ
�`(
�A�W��
� 6j���k�U��܃R�Zڕr��5�����U6���<��#<���a���YZ�pm�Yީr�Rۍ�I[Yo���vSq2�2�7�c>�ؼ��*a�-��U��0�(���)	fcq�K�.�؇�S����u���%6�d\�k���J�p��V�0�����#��`�\�m���^��
˲�'i�����j��V��<#![;�n��Blhͺx�<%�������c���W%�Y�n�U	UUFt5Gir ���5�T�ɨ��\�f��@�m�\�VҨy��C}_�U * ��S���WTJU=3ۊ����������I�l���YZ�
����V���Z�V�PqUUUuJ�m/-PPt	Nh.��=d�AB����n�7DK�C��+FEڪ����p�PUUJ�T�M��u � V��QQW	LSE�ʫ�� YEX�i` �vV
���v�C�����mĄ�C�m2��AnL��ӊ)\�@�F �kV�V�X�f�UU�W(����A�ąZ�a�U�*�ݕj����uU����%�����f
�ݶ���I��ڥZuY3R�������P�ۍ�\�f�t@�N��s`xD�����[L�Z��1N#�86
�Z���Zt8!^�*v�TL2��!UTJ/9�gU\R�Kc
�1<j�,�5O��J�%炪��50+v6[��qmȬ��]U1�Kn�N7�k����4fv�s�/Wnyq�)E*�[n�����Bk=�+-Mbu���������k�<�8���f�݄q#��Y��Xئ�:�<��Z1��F�̏j�T��8�a:Sv{; ����d�#+�VX%�!k�/�+�k����:��{�ɰ��ٶUԫR�,�ԇ\����8/@R�+�ӱ���l@+���US�K��9�jJ�B��GU-!̙H����T�eV1V�*�ѩ�2��+�	��fyP��j��jݪf�UUe����e�XP��J�V�$�T��R�P<G m�7"�ڪ��j�Jm ʷ⟗���*�����`7Hfk�S�:���ʵU\���ڥ&Ic���U̿_|c}�P�cU\Dt��8٪��l���v�����k��퉦ƶꪀ��]��jT�WT� J�P\��4�L�D�s���iuKUU*���ڮ(1�4�@k��"ڨ����7g"� �R��6m�W���c;tW75UUc::����1P]-W ��Sl8���e�P�ӢUvg)Ҋ�<����a�Wv���҆х5��E��T�Bj��U�^LM����IeYGm@U++UUU]Ulmt��ɤ�z���0᝽rc��V0�[&IX�<�S��6��Z�JL����@]tcU� ]�P;vWq=f�j]�U��4t7jB�u���u�8��[Pl[T��[!6�Wu,��O;+UH�V÷.��qKT�F���2�<���UUUUZr�V�UP�l�1����ҭR���mU��N��1�ʫ�]U@�lgQ=@jj� ��ꪭ���+N�&3��`\QUUU� ��mñ"�U[�m�]l�Q#���Z�ni]��ڗ��Aą�s�l�Z�n�P��K�r!�E"�ΐ�����
il�a�Z4��d�ѲZ�{���*x(o�.(��:�u!H[X�cl�f)	��9M)�s���YFtl�P!�r�4�;?���)Gr�7�2%��b�9n��kõ�u׺���X��Bm5b*�Ab�(L��h,�v�x�l�f���'�]�U�U���mk�]���`x��=�%��h�n32�UmU��2�'de%��k����ljv�m�&1KUUmR����m�P�@ҭ�� Э��<��V[DPXӆ��F7`ȵf����U�'l;/XԵWUU�-U6�����.q�ʶ�`�g�kZY� �@�SUU�J�m@aKZC Zڪ����C{�ۢ�@��
�Zڠ����j���(mgi[t�rlK�7+F��`��[uUT�T��r\Ie*�X�kv�����s�9��5UUS�M�yL�[&8�R��!�kk���E���8����'��8�	j��*U��=z�q67+;-�U�G�܀x]W�MP�F�X�T�6уm�z��[��X�t��ru�,��U��@I�L]>�JӐe� *�wi^��r���WNɺv%�y�@s�^�8
�QW�Ф AZ\��UUm9���ԗ	kl���@6������]wNV��SFE��鈛r� P(u�����Hx��][K[V�{6�ݘ9z�힓��q��:��l�6Y����h�Gn�z��Ԥ�c�� �����UU�uvZ�]�ʏtB 7u��4�/&�6�L���UUUUUsjCkcs7J�h��B씝ش�]qv��VIk�ƌ�}U�K���̫U*�uW�@
�˳Q��Q�� QW]E��-![*�֑��!�utܮ��p�|��?J7X�4*�]T'm
WP�n��,��È}���z�ح��ꆪx,x�����'E�м�s��{k<���]�ttp�c��$XW)���]J��mt��#v�F.^:�p@m�
KT�pd�0Z�V*���q톲���rQ�嘳�eX�5�R��*pT���m+��ۏ2�gE�i�������7)��g]UuV�+ݳu\&�J�pU��%���j���9�@�+���� �1����N��
��]G�mk�&�!�� �!�j��V٦�X�T�!�kմǳ�v�{N����ɻ��+�z�]U���Yꪪꪨ^	vZ�8��Zy�j���l�UUlݪ�2o`�s-m*�YG�йi�m����,�ɚ��JS��()^��NԒ��ok�a��煫�*���S�
�TUZ�a���1����V:�VY���i�Z.U�#B�mR�n�uUUTAؠ�꭪�iv%��T������m xث�qU�UB���Zj@���AiV���^�]�j�j�.�
�*�A���!B�uL��U: ���A������.�ݻ]���UUz�����N6�u[UF[��`����5T�W��q�������v�`��]���ܰ�a.�֩yZ^R��n�@��j�Wf�SWZ�´UUV�8��[l�[@U�uV��m�nb���Ucj��1�M��%mRR��o0X܌Um@K��Ub�%m��PVUUZ��*���M��h����mS��U@9��tP-��=/v�h-���=���q,�8^YV����p�����dUYU֖\��0&�+Eʸjj0���ﮭ>��Pq�J�U*��UV�(g�UU�=�99�4�����5�UK�����-��d0@!+=�<���؝�lU*�R�����ܫ�etM��ZP0
��X��UUU@UJ�UU]�P��.fs�2�ѪS�uJ�*�m[�� �*�IDwڇF�d�Ե++U�VtR�cUU@\$-�����kt��UTp؜ZTn��źu���<�n.
k9ʷK��Ӎ6�UT��%���R��ʵN�5�c�9�嬆����BdV��tD�ݮs �t����6ԌU݀ �ɺkP�H]Z2��^L@T�Q���n��ŴH�۪����y`*�������n�s��j�n�.�193T�Z'����Nq���sRc��e�[�mR릓,T��5*�P�+S[\礍G��r�nr���I����ۆYxrT���,+n��7g�0J,F1�@�XԵmZ�����U\�)W�P&�颀��:�n%�q ���t�� -��G-V�R�UHM]J��UU�@AL��UU�mUd���<�E �L�U�W*΀%s-Tjj�P*�X/:،)]���p;UU]m@R��ڵ-ѵm\���	`��j�����U�j�m�� M��"�@���Q �S�0�,H� Ȋ1�� ��E� C����6<A����4���P�A�O����
�`� M��Oɱ�lI d0X�� 0��" b&b0�/�P����SB��O� D^��E��.ǡ� �Av��_�� ��w�qQ?;M��U^�����S�V��Dz ���+�T҇�l6����1?&��A`��8��M ,h r ���t� ���ʏƅ�A;�!�E�'�~T�uU*�q��z��*�A>؊�+�D
�Pt3A	����I�qT0 BE6�M���*|
��~U��1�a�$Qd !"@]�t*&���� ��A��|�7U��Z+"�0�X@� �,%ڂ?"bA���Ux�qP\P�UN�E��z�����D��b��Q>H�TD^����B ��B�IZU*!FdH���Bd�(AP 1R�0
	D��H!Q�B;�wO�����(��j���i]�35U@K�ey��-�Y �.]*�c�h�z��Y�� �z�]R���,�\�$�s����Z%�u�i�Ɉ��UgNI)�G	��+�`<��t�ҥJ��C�0j{L��
�!B���-�vØ^�,���uf�u���u�&���S�9\F���D�I���]��eL���@�M�h,ke�:6�^�K�l�˴2u����.�$�SGp�&4���R��+M�f�D�����X����3�lz��`"�e.�yJÃ�+m9h�.θ��9mQz�2�� .�E#*�W+[�a�[�IqA�G��ha�s��7J�R�-ۂnЎ�!�f�,+�aÊ��r�դnڍ��n�쑻�F���qg-����7nw\���&�d�ry	�Kv4��ME���+re��Ǝ�w,J��Ӫ�`��D��۶�p.��p�q��BS�]n���J�%�L�<��9�}��t�R����1��<G��g]Ϝ֋]l���۠2X��4����m��ĕcBvg\!љ�v��v�Hv:�ց��&;���̶v�6��,�,���ujH*�W��'b:��\b&��jŠ�mۦݙ��vl��Xj�3�6�keh�b�CD!�m�c�+f��h�0�nIi8�ƕ�7k=C�=&YqV�n��6`ݸ����<m���Έ:[�"�:X�6mP�-�PBط.�/*ziP�u,q]�$�l�`����f�f�.vV�Yp�km8
�%�E��0�P9@�.wu��a�gq��d0�p��3U�Ĭ�Q&�Ӵ*6)���n(4�K�N�ue0�A�e�����4����TU��\�$�V�uX��p�k�g5we�� {&�:��nˮ����;q�x��!�;���d�8 l���� ���ۥl�э��+
���%�X^�ރF��)͋0��m�6�F��2��]��x��`���Cp�'`��5�+,H�2��i���b��l��m�B7:I�;F��b����a��kZ�('���
�S� ��C���D:+���Tڠ&��zf��3;b٨�
�a,�\d�v[m��n1�X�`�&W��=���4�u֐�ł�L���i�,m���h��{�ӎݐĻ��j8��»���a��q��s��+5wkɛwv�]dj�hF�W�B7C
1��fF��a�Q��4U������s����)F���͡[&P��>c5-�
Y]O��$��Iibɤ�7 84A��j�u�ـ�Y�֒ٻkI@�i���qq�i�K?�͉�޽8��; �ݼkذ�Lt����>6�� ��� >�^5�X�ذh;�r��[V�7wW�I/ ��,V��vJ��Ңt��v�t�wwx�"�5I I%^ l��v�Jj���豻��H�X$�x�`9+keN�	��um��/@q�hSi��x��K��YBƗK�an{90O;+9E��X�lNȯ ݗG"�;ŀuvU$�!��uwm4�{.�UqQʮew�\��U���>s�}� &�/ �n���Ruj���k�`ױ`݅�Ip�5iM)VZ�N�wo �{ N�W�oe��*������Lt�-]*�n� Nȯ �ˆ���b�=U���$;��^��I؝�VРW`�c-���n��u-lT-�����;���5Z��~|`I��, ��^��[*6*-�Zwf���b�	ڒ����kس�yz���*�d�nI���]�'~;�nk���4"���J�B�@bQ�H�E���\��I�Jcm喕&۾�X;R^�dx�"�;ŀ|�*�r��7N��mӻ�5vG�N���, �[/ �p�%[wv��);�,-T]u�&�R��;�[�+���Z�ͱ׌O9*)�;t��	��-�x�`�b�	���]���Q1�59l�N�n���,�9UI{� M�� ��,�D�Ț���Ҫv�`���엇���RS�y`�<��Զ]2�N�rջ od�cذ�����3�%�s����6��ƻ#����ݼc�`M� �6 ���p�����,�kUmZ��U.�Ͻ}���8x�cY�lWm���&��[�s4���v[�i*ai���^�x��xSc�����}=�M�w�Q�P G-�Kf�5M��"��Ȱ�ǀuvU&�bi;,wwc�"��Ȱ�UR^^�x^����8���'v����=�s��=~��o�x��x7e�iCS�ˤ�&�`엀j� &�cذ
�{�u��
�f5׷��2�64�#�O<�p&��ۜ [���)�!��7)lm�l9�a0�E+n4�RXP�]l�bXa�!qv ��R7���ONL����b�0�F��tmѤ#G\�R(�Ik��q����x�c������}���\�J	�iܚt�B�s�p��ݓ��h0�����/g������vq�l����ۂ;lo/��C���2*�'3��l�����㡗p5܏�!���C�����<���&�]a��.�6l��2k22��_�v����ݗ�l{ N�x���N��t���c�	�/ ��, ���n���E��bwC�Ɲ���b�	�/ &�/ ;6^6��uj�Ue���6�`~��q)����=xٲ�	ױ`ILOl����� M�^ vl�u�X���s��9ޗ��� �����D�-I�&I��y�6���B�b��7���wR�]�댻�%2������b���r�\���>x���7�Ca��tG/ ���n��"%
���l-$%!H�k `XH��D�	!!�[XHɔ�l"D���H�$`H!$	!
[	��bƁa �� ��ą���C��������v{X7e�-"bi59n�'M;���^ N�/ &�uȰ�8k2���^�Io������� �\� ��<ii%�����8Ze� M�x�`vG��K�;�[��0��68�s�N���m��G!����M7*ۥa!;N�p��t��n�>��N��� ��^�6<mz�蹶 ɣv[�=�ק ;�ӯ �:�X�SI�m�Ӻ��;N� ��^�6<+�\��]�55�Xݗ���6JCe$;jڧw�uM� �{�r, ����Mj�7��j�X�� �{:�, �����/ �D��caWmX�gA%L��Gt�\F�zfM��۞���`�N���Iہۦ�Վ�M;��N�� 'ke�ݗ�N�� ��uj�-��-�ـ����ď)<�k�X�`T��wV���
�o �v<uȰ	�p�&�c�7u�Q�E����wx�`��MfǀW9\�9�$������^���Nֺƌ�9n�;�ܮUW����l���v�n��s5�օ���h���S������@oml+�����fjs6�(��Zv|�'� N�uȰ	ݸ`.ʤ�)���t�� ���I\ŀNˆ6�ŀMj�7�)ݕc��u�X�`�l� ����YM)V;��v���'e� 'ke�ݗ�N�� ��uj���vU��0v�^ M�x�ذ	�p�
⣜��*486��avu��{�p�ѡ0��mrh�]�<ջ2�� h5�ۀ��/e��Y7�V��,��q�Z71��sҸ�68ۋ�f��L��m��;��<�wa[GS�as�ͫf�{)`�Inq�m���&�7n֖4�HZFU��&�V4��4���Y�1d3�	��^�m���e\�;��P�v�ư���a��wg�-j�n��X"z�Pb�{�ǹ��ɺ6S4�ۆs�9�dk]��@p%,f��gg�/l��"0�r�W0�+v�(�Ww�M���b�'e� ;�{׀{�qЃ�:�^:�,v\0v�^ M�x��a,��գ��-ـNˆ I�� ���	�p�$��n��6Յ�Jӳ �i M�xݸ`��}Kgܠ�RV+�j�x7e�v�I�)�x��j�wn�r�Z��-��uE�u�&^���cθ6�۳i��|�hV�r���Ӏw�^�)���W+���z��z����n�gl� �������/��H����9��3�< ��n�0�A��U�;m�*ݻ�)�x7e�v�Nɕ�M���.�m
젦���n��&�� ��+ �VǀoA��Qw`[�i��&�0	�2��lx7e���Q��WwT�N���׭�@r�I��e2w!�b�����2�ۂ��.�5�5��8rp��y8T�� &�M�`II6b)6Ֆ�J��`M#�	�/ ��v=9���/~��}ĵn��w >�}x�p��ߥ�Q�T�;t�2�j�,��?f�B�ZL5���sJBB+�']zt�u�M �9���#��&��K*T>����J�:4�d�iZ����!�h���m��7w������O�-7���l&�,�k�`�� 7�麷A�3z��N�<��C���q��,Fgl����_�>0y���_h�9�j]�3����~��T�[�}��E���R�a��|��Fp���D>5��Mk�e�fn�5�{�e��}w��v?o\�8�[!� �~֤�&��^t>��_�`��D�Ͼ�'�p�&��M�c��<�n�n�w�����tڻD�����Q��F!"H@� FX�@��H� �A���A�+D�W���P�W~͗.ԏ ꜕.�t� ��V[��$ۆ;.R�<UW+�zO^��&��e[iӶ�ـNˆ�� &�M�`]Im�Ndd�&�u��9qw7Vy6Azw�N	�&L����nh���v�S�v�lx7e�m���r�_ ���`�.|�kj�%����^�}zp	�p�"�G�oA��QweZt����v�Nˆ�< �������+J�_ݲݘ�`J��䓿�w[����D#"�=+^bIE�oǹ��o��E4܂�I0vS �Vǀv���=� �zX�ݾu� �\i��(�֚��-ⷎB].nq�k�=W�9�8��rݴ�-�������${&�0�lx��Q�'@7vU���	ŀI�)[ I���+i�
YV�t���X�p�"����/ ��XT"M9ęm��v���� &�x�b�&�� �L�v:E���AI*�x;%��z��z9�Mr��'�A~wsST�Y�#i��L!���D��Ά
�F�{' ��R���i�+�fc��6��9�Ab�u�pq��F�ll\���p\�5�}rM�ǝ�q[�vMtZ��H���=�쀼iM��we�u�vh�nE�^xy�k�d]�t�-�m��t��&�,��O�X��������8��8fV���@�{-���]q�S�X:����������h�FV���������է��ju�ں�Z�P,ZZ&�%��!sA���&��Ӻ�Av,{U�i����@�_��	�b�&�Q`엀l��e��V�L�N��x�*, ���	��J�)'�Bi��o�+��Mr��	�/ �.[��R؎7(-�n�ZV��dx�p�"ݏ ��E��*]�ҧ�;����l�`�UU�'��z?W� N�x�r�dV��O�ն�Rt�zL��oL�cY��	R�����0q	�79#0ĝ�&�+mݘ��0	�TX;��	��j��R�7m�j컳 ��E��*����UU�G��	6�N�tױ$���o�{+���I4�~���$�.�x�TX�j�R��nʶWwf���yl��$r����g�{ȯc���[�m2Ɲ�]��U{����l��E�~K3�yw��K#�9IIbj�*���L��s7݅�����!��W�bpo׼����6����}����,u�X�E�7���o�s��y��b���ۆ{���?y`[<�	��W)"/W��:N�'vpN��s� ��]Άǐ���H����b�j���%�BA$�� �FF,((B,(V�lA�Z�R����}��tXd��T�SC�I�+j������s� ���,v\0=�W�s� �ǒn�g폎˷k ��,�ʪ�����Xf�0�ʮUl	^�M�������&k`+�In����ȷf�`��p��\A6�)0����O3-�sR��`�;@���G�`�{�\��{��4j��y��������${~���U�6H�~X����`�g���q"z"��۱�I�cn����H���UU%���{�y`��&:d�*�*Ji�$�a�_y�m�z�w���r;R �Wd�E� �
V ��	�_33^����o�燇� 9aaef�w��z�U�\����,G ���|��"b[��8H�30�7\�T�C��p�t^�ٻM�Y�u�����'+���\��=�<��Ȱ	��+���V O*�2���lV�ݬ �e��ٙ#��~��6�~��-6��Κ� ~�<�t�eFRۦ߽=�i��s�Z��ě���������"���[|����X�s��{��'���	6^���r����~&�}�k��ۖ7l�M�vr,�9�s�US�����^��<I2��xu=��kE��]k5�8��Z�E�n�ի�ǔI�E:�[q�p)v]�z�!m}����\����7�5<��� ��,��x�2��j �Ǳ���n`4����4g)Zz.�G���c,�����@�2��s�G4����N��N�S��ͷ�v�8���\�i���W]�9Ω�}A����퓻s�tNpq�#�#�e�κ��5��=�H�o��8WM�Z���]��M�?&�l�Bw�خ��K�C%.f.�e���.�5҂�q,m�����x��<I2�U_ �s� ڒ�c�4��wN�&��["y���%߿~��oߧ�m�������G<<<�Y���Zm������w�� s������t nqq�ڄ�څ�U����,̞��&���� ��M+�?)>����Ǜ�A�`��� �����ΚW@���o`����m��?wn�]+;*��2��ck��j�ѕ�‡�+H/���rO���i��jx������ o�����;�<� ;�]���w�Q��pѫ�Z�ݶ�~�xs�w�ɅLQ��B)Q*G�уAm4��*t���o�ٟ}��m�g{齀q�U��$����ۖ7-�{ ��� >��f� }��W�|�v���>�!���U�l� ���� ����@���o`yN[�I���'�l ��ZrKw����$��g���RK[�oI.���䒔�S�܉�^=tY�[VuƖc�]w%�xN��S-��p-��I�潼��i��f�$�g��}�Iu���I%��~�z�Z��W�����j�YE\�o`I�ɯ%$��� �}.������H3�[�A��FXYd� s����}��s[��qF�Z "�
�@*X �P�� �M��g��n�ｵ��zOzM \���iR��	-���X�9_}.���mo`I�ɠ<�)';�]���w�Q��q\u�.����o`X�r�zM�;�]��>v] ��N���F�Dc�e�B�x3��,����k5��ۮ{sd����I�r��@����2�߭�$��� o����#�e�$�܀w�����+�=[b�*�\�ɠ ܒ����WhR���I)'���I.�#y��8���'�b�T�r[w�uw�� �9ݭ����X�����4 �����>G:��*6�
�)e�X�I���-��{�h 7���`w8��8Q
$z('T</�l������~��1Lr�d%[��w�h ��K?f+�߿^p�^�.����o`���z]�N���+7#V����gd]D
�]���Lж_zH�6���B��ɰ �������ˠ�s�^ŋ��ޓ@W)�)<�+*���`��eגK2H�}���rOzM ����رfI�%QK���� �{���;�4X�I��]��]�� >]ti��4IZ�p%�{�ŋ�bX��Z��M ?~�w�qs���K�b�Yo���[���S�kn*�\�ɠ �{۽�~X�Y�,�J_/~�������;�4 \����F���`F"�z����!IcHN�z�It�L!	��B���>�}�gv���@�S����Q10h��d������8*�����i�al?s�����h�	�������]taN�p���Ԑ�5з6�)HRFS 0�D���B�%XV���������Y�r⮞FqV�1gC�J��
,V�(��d�	�]���a�E$D��@"��@�5�� �c���Cf�W�0� �8|H2�+��0���aJo�h�f�7����Һ�ÌI�"�o���.��YYJX�m��I4���~���Z��Jܓ� U@UP�*i8ꀶ�
��y���m�S���b��s�؎��bhL8�N�a�XF^�ϴ[t�v�)�Yu�B��n���)����eb'��r爎��U�O;��+²��(j�Ft�i�n���4v��e���5DN�A���rX1�Lt汉f䁻Y�i"o�v����x�)y���4��1��v��['1ד��ˣC���.ȥ��v*t��jq��qڥ�k��([�`~s�̤�Cd�k��N�6�e4>�r"v����F�l.���\�cfr��8��74�mV���0e�a���\�M �
�1�ˮ�z�f��X�m���*\�))-5�@�X�m�tƍQ�	��|��ڴU4B\�P(݉�Dn�YEĄ���0����U�aL����:��4�̫6Ѕ���s�&�{vm��.��D�ݭ�=�t��^�I�΄ȣ�v�NȄƊNLv�spq��7lcn�9��ͭr�[���K��9�̰�=P�v�����N{�z�t�ʞ( ��P�V�a�j�v����[��	h"#�"����m��˻�K���3�r�+l������㜎�w2���az�]�V�9p<{N,(�v�nl�����@�Zs�����896��+��#����õ��	T�@�`V����n���nd������!�lO+g<�:X�[(i��3�cXg�����Xާ�Ε'�q5�u�jG�S+;��{m�o\�az ��7S�!�m�ٱ�t���d�6n'��9v.�C��H�e�px�86J^#m�Þx�V�!�z4tְFɎ`�7#�����g[n(b4��:1�XTK:�K.�:툝�eaA��\c��g{sȹ[���[���;=f��G&̘�	뫨��N����	�a�ؐ��,Z�LM����4�>틲�=���mEz�J�GK��8�'=������w��p˹Yk��l>m��`��j��.�����*�:>>S�P��'�ڜ:�?�G�Ux����:wN��'�o���k-�'�0dӫ���mp�ʜ�4l14*&B	vu,L��V�M�N��/d�d����]��j][�e��Mf�q0t�8�@)r�n��F;-�9gB`���PDw[���6�W�i]8;v��#�^���4\Ev�T�q�]�v�:m��M�ys�ʠ=�VØԇ�3c�}���K�sMۖ�1Z���dmƒ�[b��r��N�]����bX�]���P����0f���o���9w����5��c��� �#A��$fe�=��%N7%�� gW�K���v����w�{����뽀q�4�M�X�+e��9ݭ���~Y������ ~���`��ۯbR@�����	�c��!*��:Ox� �����@�����{�� :q8(�ւF兴��I�{뽀��n��������}�h ���s�er��Yn� �� =��w��}���@�s�{ ���Mѹ�V���m�;+]*j᳸���(Q��h�J���)��o�J)TR�lV݀w����:N�� 󝿒Y��fs� ��~�@�F���l��P�%�{ �;�hJ�kM5��Q0@� 2Ad� �1�@�-$UT�Z����\�uz� �;�����bV�������V� ��Rh 9�~�� w���=��O��mo`'�M /����$�P�8ܒ��b�'|�n���mo`'zM�I>�}w�)�!�I���e��v� �;���yfg���� ������]�@3�0�)eB���d�GX4�Eŷm�AeP�h�ki�K���z�1[Uz��1L�kU��� �=�h 7�v�`ޮ��g�����9�~������q�C �i4 �;w�$�d�yz� w����:Nt���K�:�D�c���Tc��� =���m�����_��A<� o[��l�`�����c9Ԥ��km��@~�I/ٙ������{ �'�I� �;۽��y,X�Y}�(��F����QT(�j����@.���{�{~��]�� 9�wk{ �u:vJ�m�ML��`�BZҤlB�pD�E��9��lݭ��S'��wMK��ap6�� }�z�`�s�� �9ݯb�I}���Φ��I)]��7%�{3��˯,��$�����8N�� ���߳�$:�}�4�M�حRˠ���[��w�h<�$������ ^�� >�\}��1L���-[��$���Y}�~�&���~�� s���ȋ���x��W �Q�����{ g��q��V� J�� �����,_�31[���� ��mocw��@~���� ���G,��Gt��v:��ְ]�\nԺ�5���יBS��Ӊ�&��e�:����;�� �9ݭ���e�,�Ź >��w��I�����B���s�Z��X�����޼ ��^{��W)#k�E�HM֪	j�m����m����K1 ~羯 �{�' �~���"2��^I�Q-��{[�O{��ܓ��wf��6���<��`}��!\� �}�����s���?~����߿~� �%�bY����7S��	�n�d�][��2=p�F�V�]O���=b}�F�.�?����x[�B��3IKB�&"��b5���-��m���έ�=�(��V�sF�h,��������CE�l�i5#�Y���d;n��؜�f�а�i��Z��f��t��eQ&tl<�)b�v���Vӳ��9`԰���Ccmͼ�FZ+�#qCr�Ν�.��](�:���E�[�͢A.�7�e����m���%�ћ�����y��F�݌�v^��߿e`�^ M��U��[~�|�|<��k��L��e-Z`I%��/ 'dW�M�+=��9�H���1�����v[�� ��� &�W����r������z�	]h58�,��Te��7�f���߻�ii���v�bI �}�߽1��R��4�n��	�e`�r����9Ϳ����߿^ {��׀~��Ƽl�K�_\�s�(;c��-���w	u-m[De��W{$�0�kj��T�wu�^�x6K��Կr�\�����v��J�,���Ѩ[�f䓿��o`"��SZ�����;=��6<���?r���*z��$��]��`�������d���\�K��� ==��>ݜCyI%`�������R������� &�x�*�{+� ���ut�n�-]�� vIx��G�nɕ����D;T��s#��á��<c�۶�^�E�[�ǡ9�֩���%t�ř4���5Z�([f�o��� �ݨ��2�ʪ��uzy��h!=e��Pvۦ���5�Ř�����O< ���\��G����Sv�]Qn�=�e`Sc¯���p�.@ *"�b��7��{׀j��<�Ѣ�D�2��T�wu��(7���7$�ｭ�?^�雓�*�{���	�`��*�WV%v�I/rO��|g$����rO׿���('���{��%�gV��g;b��I�E\[���Ź�ڸ�\%�slNt{7"�WF�j��-���I��uM��9U\��{޼�{�o(H�t�j�n��I���UUq#W�� {����%,�_��Y�>���~��`�;j�o��~�m��/r��RS_�K ���R6S)Z�([f��I$��t��'��6���f���	�_��s7$�r���f����j��wx뒖$�XT����� ��'�Ϗ��Tr� ��x��=����98{v�W4�f�xv%�A��{ѭ)	��V�I�j�6�{��-6�$� &�~��r�A��x�+�j�5e]*i���5I{��r�Oz�	����'w�7������O=�$���QEic�%�m�����ý�~X�$��rp߾�pg�|;�]Ve���\s��U(�O �����#�	�^���7��V�L��n��d��=UU\��y���^�䥀:�9Uڕ��Y�Ͷ%�P| E���n)����pl<����)��Ҧ�o�ۮ3��4Sl��y���rEl��h�cq�\c���79N�n�ư��W�;n7�ﶯ�I��;H[e��8yA�p�I�v��K\\�pxm*Cvwg3�Uv^��8�q�cGjgu\q���q6xp���f9��Mi✎�7���⍘�.wcVy��k�,��e��5�:I1� ����e3]B9�;]�Ĩ��[\����e��r�c	g噘����Ur`�^R� ���< �K�7\���Ur�A�{�X�S���q�۴���	$��+�T�#��`��V�$y��*�:�O�WM���-�ۻ�$~�,l�X~�r����y�S�x�����h�;�˹<��w��'��{7$������P�bS�����oˮ~��ъ�Z�êH�s��W����{޿Q�Ix����~{��aYcA��o���VXP�6��6z2݆��eH^�m�IB�ӱm�`�.�jN��y{�x��$����9_ ���n����uY�
M\����8�"$B�t�Qf$+"# �D#��! #h�Ab��E̓^���'���ܓ���׳$����H���S��������N��O��g�32O��ߦ��~���5J��WƇ�+��n� �H��� �\���+��K��� ��y��z�1�����I�r���=���|�{׀E$x��N]�j�:wC\�Hq�c��N�ʐY�MIf�+.�ZC�������N���c5^Q>���{԰I/ �H�\�9Uϐy{�x�ty?SZ.������IxRG�N����'{��w����O�a��(T�;C�����~���I
�,唢~��?�] �0��9.�^�qr���)��$����s�HdB�??!߳�l!�c����@�P����,�H�:tY��3"����Ձ6)���L&�����H���̘|Z"BF�?���J�ҺW-E��F�2e��Bcd4?�N~��d§�;�d���϶�H�݆3x��of�a-)��lÓ9�$� �I!��|5�%���H� Ȳ����k_i~f��͎��9�6~�ç�@�;�_21��|�18}(c�T�����p	�	�hءQT�~>D���A�?���S DU*��@����LQ k��9��I>�}t�����QuJ+m!XK4ߖ%�9�<�s��	�^��]�RmV93��]�;��K�>�I��������"�<T��V��ӧE:�>���ڔg��������;��N�\]&g�p���f%.��t�eAk6�~��tRG�E$���?W+��ߟ� ����E��5vR��"�<)#�${�Iy�W)"#ǙL��:�M��<��x�j,?W�Uq�������~�m��g{j�˖ܶX[4߳0���, ��� �lx�����9TUET��}�ܓ�L��K��F�$�V�M��{�U^~��9�H�����{�i���\��qqȼ^8��x�{��%ø#n�J�� b~ř�::�puv�uut���/O<-��	�<�Kco����{;Zj/)EIc�B[�&�� ��E��^���Uʴ�{�_��m%6o �����엇���//O<��,lT
b+@&M]��UĽ���^���x�JX�Q����vS��"�<��W���9�`엀~��;�|�
c�T̣@�A�c7mRI���rs���E�1��urr��ݻ����M�]�-�JGl	�T�90Z2�څbb�e�:��i��^���+m���n�Fk�Q�C�l�km�g]"u�8�X�8viB�4J��&[�.�B��ۂ�Odʸq٥�#g��P�ʱ��b�:S�jI�e� �.ݎ�����B��6mxlB%1�$�N�����Lvz�ɑ�ЉѪ�<$��.nZ4���j�� ?�y
#1�x�N�ջp��?� �� I��	{���zެ�ϊ���w �w��=I�=x�����	��	�L�]]]����l�)����*�ļ�<�y���>��)Ƌ*�����)��M� �� I���m��JC�n�M�xSc�${�l�)#�>�ѧݫ�LJ�b,*	c��1M��$��{�6M]t�౫�1+���ċ�1S�)4���煀l�)#�"�6*�
�P�YsEܒw���Ӹ���H�D?��|�>��s��>�/{�x�JX�Q����;������M��R^���`�=x��h�R�],�M�{3'��V߽=�i���J�s3����}~�wٖe"�.u]�;�ެ �e�I���Z�ЋE (Me�H�q�����ҳ:���cb����7�)��Ixd�ד�b���zz��� �H��s� �����'�LK�v�Rn� �H�	� �ȰI/=��$o�,��B؛�����=}�f��w�s�(��ٙ�K�����ߏ{�M�/���D��D;��Wo �ȰI/ �H�=������x����
�4�Vݬ �K�=UU��y����H�X��Y�s���y�g�{h�,%y�n�d�Գ�(���s=�JS*vJ�g�Ts�� �H��� �Ƚ\��{׀Dx���)N�ջxRG��RG�����xRG�|�c�UwV]�]���H�X$����K����=��m��:�I܌uUZc��o٘���� ����	ŀ���s��rdŀ}];ۮ����J����w ��>��_�?y`�/ ��h����˦�S��<�d��ۦpx�V��K��2��M�L�"ya��M9��IY%�m��}4ۑȰM���\����J�b򦝨����6��ޚ�ĳ?)��߮��߿M6�w�����ؤ�4���X"������߽���� �lx�E�|�KtZhe+v����{�����<���	��Iz{׀DW��B�]�մݼ)#�?r��޿y|�{�ܓ���nI����E���@" D�d����Q�MnL5��\q]��@��[i�q'X0G<r����=v��'n;��,�rD�;��ew`Cs���m�̝:��u�ݗ>)��N�gVuF7FN*:�����۠c��ԃ�]6�nLnѕ����'v�9:H�&�r0q�	m6�e�k�.�i��Eg���j&�,�[��<���&�Dg�,Q6a�6�4V��K�I{���-����[d���.�ʀ["Wd�Lk`[ݜ,�b�#11j��f������vӷ ���, �K�"�<)#�'G&����.�`�^z����y�^��#�`���F:J��ۺ�M���/ �H��E�Ixҵ\t�wccv���c�`ŀ$��9U�s�OO^+eЏ;N�2�q]��6=� 6Ix�e�� �B���M�M]�EZ��F��0J��5$h@n��0CP�
yuն����@�f4��is�����^ {�z��b�W*��	�<��G��Չ�I�SR浹$�������ʼ{����v9 l�x���T�,��N���b�6=�UUU$OO^ w�����^��G$V.�[�=��� 6l� ٲ��b�;���Sut���6^���b�${�bQ�c.�eճ�鶝���+�&�
��xY��������AZ��4�[��ut���"���X�b��/ �ݸ��$��v7bwo ��,G�`͗�E6<k�t"���L����H�, ٲ��Q�PDA��������nI���݁��a��WV�tݲ����/ �lx�b�${�h���Ӥ�c�V'w�E$x�b�$r, �c�=��n�r�P�&Kuem�I���[/=x+���^<v�jx���"[����m��m۷�H�,G"�	6^��)B#�o�we�.�`9 I���� ��X��b�]�.�`�/ �H��^�X���O�����c�Q�e���w �s�n��w�rt"#����fbY�ֻ��6����Pp�YKS%�G�`����_ {�׀E$x��?%�	pJ��ع�����s�m(�IX9��:��F{qQ�M�H�[�7Na���R��H�X&��"�<G�`(6��.�tݲ��`�/ �H�	ŀH�Y�s��H��Mz�Zt��v����/{� ��X�E�l�QSiЁ�K�4�;�x�b�$r, �e�I�(�	v�wv[���#�`�/ �H�'{��ܒ��߾��;��P:���$059ݻHH f`ѭ��!�$�0 ȡ!$ "~�����,V �7����	F ~�ĒD�BD�I6�Hd�!>��~�a@��h�FTK��`�L�q�IBDB@d��.�6o'zHB#�j�i�"I@$'�k���F!2��$c��,����XBwb�F!$$�f #1 &a@���+��c5l&0�4@ ��.$c]�6JB0 �	7���.��
<Y��SC��R�H	 ;�����1���%8�e�!�F���u'.�:��-����'� ������T�@UV��ea�gnX^#c�'\�G���FN[�-���VÉ���@���]%���MbۆK��.j�a`��b�ێ؏N�m@��,u;"�^|$d�aܩ=x�뛀gm����	�0�YD:��om�R��#m�]gtr
O4-U�`�tV����=�#n�PuJ�ӌu�$䶵8����ؽ��\��J�jN��;�]Ԥ�1enK��
�Ų�:�9IzN�FClom���=mK�@*�k�*��/7
	�dX8��C�YR��1j��Sd��ӮË�z��ۖ�p��5�8�s��a+��iJ�k��x6�����A�H�Ʀ�S0�*�R�a �v��;��^��;	�����a��t�L��:.07�u�����/\nϢ�鲡��{#��v�6���U�^y*,��1%Yx�U5r:�J'fZ�n�#��s�U��.���j�Hj$W'9p��9]Ŭ�ֹ酲�d!�����#+����jc��XWP��,� U�T3�����XV�Z82a�1�1Yh]P	{���i1{v1C oX��F���p����*�.5Vأ�B��]�-�r=�M����⺬7X5�bX��N��c����ݺ ɩ�>Q�k�;6�XŻ%��Ũ�5i��uv��>��Wc	�Ǟa7r�I���݌s��9��YI�`�Nit.���u�<�p�v���:�a�j�vjv̺@��{o��&imL�x�Rk�G�7jzy�r>&H�[g��,��EZ�1����ʎsTlT�f�6�b���GYY�8kc	��j�h`�)-�$W��t�E/�!�o�:��;7%kp3k�ƶ8��i��yzb)�s�'ef�l���R����ʋsȤS�;�˒�KZj���|0P�!HB�l9c�ͱ��I�3��%JGT��],@ѕ0�c3��
�;[A�s��.M�R79�yz=/xtmu�hq�ֲ�v"��mul�浮�"�%Q� ��J�B�C��Dp:"�i����?
'���U�\��.8��r�h(ώ������ֻqv�ݵK�U�<�V�/	ں�'���fXLY[��aK����T[��F�Ҥ(���5��S�gql�[ݱ\����[�m�ϱŸy�r���V��X�m����R2�h��ĺ��o��B{��m��r�k��B�+����B���[���E�ΎeMa�gD�	ET�7�xeѭֱY�ZΣ����x��i]ɸ8nmn"=]�/c=O�ˈUlJр����xRG�H�^�Us���������*j�v��n� �H�	� �ȴ�}�{u噘��q���BUae���y�� �ȰI/ �H��툍'j�*�IݬG"��^��� �A��M+�m�N�n�`�/ �H��E�H�X[�ߟΆ��&@N+
�>'�����W�RYr�5JZ�Ȩ
�S�g��ē�+��"�<G"�$r/Us� =�z����B�K�4��ݬG"��pFlG�E7���������$���X�P�h�*�ڷe�X�"�	$�c�`9�p�K�V+E�X"ݬ �K�69#�`� �tJTՎ��]����Ȱ\��_�ȰI/ ��	O�Qfv({Bk�{vsgsΜ��N��$7�nG�d��CcCJ\��L��]���;�ޟ���x��x����k�!�!�?~���?�)>��,K�����ND�,K��i��
�N��䦱m�!�w���Ӑ�PF9"X������r%�bX������ND�,K��}v��^!�.�7�-�7U	�;-5�o�bX��ﵴ�Kı=���iȖ8*'���0�M����]�"X�%��k޻ND�,K��˞���h ��VKu�o��z{ޚŷ�ibX�����Kı=�{�iȖ%��#2&{�[ND�,K��d '�ơ	Im�ŷ�x��x���Ñ,K����]�"X�%�}��[ND�,K��{6��bX�%�t��b�1M]Tz��eٌ�!V�%�nlZ�0Ԗ��n�g5���D�1�z�4|��bX�'��z�9ı,K�w��r%�bX��{ٴ�Kı=�w�x���=W�g�Q�;��,���,Kľ�}��!�ș�������r%�bX������r%�bX����X���ˍ�׼����KS��m9ı,Og���r%�bX�����Kı=�{�iȖ%�b_{��ŷ�x��x���x�"-���'���r%�g�02'����v��bX�'�����ӑ,Kľ�}��"X��0�c�^��$��L�%aV��Y|D�Fa
JK�-J^���S��"{��ɬ[x��x������)m�v��fj�9ı,O{^��r%�bX��ﵴ�Kı=���iȖ%�b{׾5�o��z?ts�%�H����Е�W(TlDII�qx��pvr�U��\�H��%����v!T]�O��^���/��kiȖ%�b{���ӑ,K����]�"X�%��k��ND�,K1wס<�,u��VKu�o���}v��bX�'����9ı,O{]��r%�bX��ﵴ�Kį����sэB��k�!�!�����9ı,O{]��r%�bX��ﵴ�Kı=�w�iȖ%�f/��<A?Jd�[��ŷ�x��x{��ӑ,KĽ�}��"X�%��k��ND�,K��}v��bX�+���3ըժ�F�Zk�!�!���m9ı,O{]��r%�bX�����Kı=�w�iȖ%�gK;��I$��:F~z���]�Z���b^��j�m�쬰�`B�n0b�X�u�@e�j��ظ�A�9$ј�6����x{cn���R{��<����;�a�qa.`TMclLb�T6E�ͮ���B�6|����0L:��&%� �1(i�u�%] ����p\k'*؄5m��v=%�1�c����������\�l�iH�݃k�*�]C4���wN��/��&+�ԅ�:WS=b�,Z�*͡D2��#q���[�1��N2�]k։sZ�>�bX�'��siȖ%�bw��ӑ,K����]�"X�%�{��[ND�,Kݝߵ�.�:�Z��ŷ�x��x���ŷ��bX�����Kı>��ٴ�Kı=���ND�Aʙ���rY��[`�O$��-�C�<C�����X�ı,O���m9Ƌ����&��!���]� �'��w��d�S$˚M�$OD�;�fӑ,K����m9ı,O��}v��bX�'�����!�!���I������iȖ%�b{��6��bX�'�뾻ND�,K��}v��bX�'��{6��bX�'�$�=��-!�kR�.G��s��j�w�Rn��i����)��I������h(I,�X���;{�X��ı,O{]��r%�bX�g}��r%�bX�{��ӑ,K��:K۔�,�b�*Zk�!�!��o|k��#��W��<�Ȗ&g}��r%�bX�~׽v��bX�'�뾻NL_�b�b��~�W��H�qJ�0�WiȖ%�b~�fӑ,K�����ӑ,K���w�iȖ%�bw��b��<C�<_.7|�8��"�fk6��bX�'�׽v��bX�'�뾻ND�,K��}v��bX�'��zk�!�!��_u�#"%��mC3WiȖ%�b~���Kı;�w�iȖ%�b}���iȖ%�b}�k�X���޽NO��b�-#�V������}��d�b0�����:���\-�*am���}ޚ�צ�=����9ı,O���m9ı,O���m9ı,O��}v��bX�'���ډ��9n�Mb��<C�<_N�ٴ�?±ș�������Kı;�{��9ı,N�]��r'�2 �{��h���If�m�!�b~�����r%�bX�����9���`Dd"HӀb��$X���$#`0��"C(22)$ �J-i"Ab U�@��蟢k߮ӑ,K�����m9ı,K��2Y.x䃬��ŷ�x��x���ŷ�ı,N�]��r%�bX�g}��r%�bX�{^��r%�bX�gI{r�YnK�R�X���{{�X��,K�｛ND�,K�k޻ND�,K�u�]�"X�%�㺽���]���Ѱ�џ<v�r��J�u�x;ۣlHO6H�ʚ����/��x ������%�b~��ٴ�Kı>����Kı?w]��r%�bX����J��|���y�Gb����f�m�,K�k޻ND�,K�u�]�"X�%��뾻ND�,K�｛ND!�/u�O�I-n�jnJk�+ı?w]��r%�bX����Kı>��ٴ�Kı>����A�!��W}�;id��d%5�o�bX����Kı>��ٴ�Kı=�{�iȖ%���A�E�c"���"cE >b��Oo���r%�bX�����KYG[�SX���Ӿ��r%�bX����v�D�,K�׿�ӑ,K����]�"X�%���߷�`���c���6���Õ2�-��e&p��@i�+p%)��S��8�35��"X�%��k޻ND�,K���6��bX�'��z�9ı,K�w��r%�bX�����K�YI��j�Y���Kı;��iȖ%�b{���ӑ,KĽ�}��"X�%����ŷ�<C�<_O&x��mQ��a5�fӑ,K����]�"X�%�{��[ND�,K�׽v��bX�'s��m9ı,O��Оֳ�f�,�5���K�K������bX�'���m9ı,N���r%�`~Ř�����~5�o��qu���Qڥ-Q[�[x��x������-�DK�{��iȖ%�b{���ӑ,KĽ�}��"X�%��P<EaDF0���$U��  `ŀ�B(Db$��;��^K���j�۪;U�N���@9붧�W�h0������b�0�@��QA\D�ԩ� B\0ہut[Ÿ�*�u�v��{H��ų�#Guj���#��� "n�����Z����h[q�I�H�M�rp8q�bή�a�d����%nD���),3�)����[pkd��&6zr f��ݪ�w9�r�,t�u��f�#��c(�4��˙�����P]�DC���9���Û�bbs��O�hWF=r���ݲ����Zl�R5WhR��(G	���Kı;���iȖ%�b{���ӑ,KĽ�}��Ȗ%�b{=�fӏ��{˾���-�nc��b�Kı=�w�iȖ%�b^���ӑ,K��{�ͧ"X�%���}�N5�x��x���X���d��r%�bX��ﵴ�Kı=��iȖ%�g��k��ٴ�%�bX�����X���|�`��lCmj<�kiȖ%�b{=�fӑ,K��{�ͧ"X�%��k��ND�,Ľ�}u�o��^~R	�����kZ�ND�,K���6��bX�'����9ı,K�w��r%�bX���b��<C�<_F������!�s�\�ʹh0��n�	
75����6!e��-J��-2ڤ(�l�-�C�<,O{]��r%�bX��ﵴ�Kı=�w�iȖ%�bw=�fӑ,K<\�^i��+�a-5�o���������'�G��Sh}�'=��v��bX�'���m9ı,O{]��r%�bX�����v�]�"Ku�o��{׾�ND�,K���6��bؖ'����9ı,K�w��r%�bX�����Q�����m�!�.�wٴ�Kı=�w�iȖ%�b^���ӑ,K�=�w�iȖ%�b{�}�V�0����K5�o��{׾�ND�,K�#������D�,K��^��ND�,K���6��bY�x�b^�����ʙR�F�B:5p-�j�.)Wts�tt=�m��nK 37������M�d��B�%5��x��x�~��[ibX�'����9ı,N��{6��bX�'����9ı,Oޚ�Yg��G,�����!�!���|k�ؖ%����fӑ,K����]�"X�%�{��ӑ,KĽ=<d��Q���Km5�o��vsޚ�Ȗ%�b{��ӑ,h�zBK� �"���+8Y�H�� ɬ/&�i�h��
m!5�&��cUMh��aL1XЁ�$��k%7���H�ACP*��HP�	B$����¨N��L\K�)�CI�6���4B�	ru�Gd��a
B�1�d	�#��M��<"B0�I�Cf��Ƀ�̅��I�Q��6*b�#�"`�ne���#EL&i��p��eK	#BL�	K(!�D��!
��F#	X#cX@�B!a�kFA�M`pF�C�U"I-� �*B��
�)�@���b �
E+B����,���J��A��B�]Ge�1M	Yt�a1@�i]@�D�X�̢h`�6��rMCy�͘@�& �J��J�G[��ݰ#)�]�*��6d$,J$V�@_�@�	
+�j
���q~A�E�(�E� �?(&*��>�{���ӑ,K���]�"X�%��x��~e�HP+r٬[x���J<_�o��iȖ%�b^�{�[ND�,K���6��bX�'s���ND�,K���O�ȑ]� ׬[x��x����m9ı,Og���r%�bX����m9ı,O{���r%�bX�w�~�?�\T�k�T%��6�8�b
���&����U��ʌ8��ћB�Z�3Z�r%�bX��wٴ�Kı;����r%�bX��w��Kĳ�w�X���������be.�����ND�,K���ͧ!��r&D�?�����Kı/����"X�%���}�ND�,K�;�Zf�5u�]I�����Kı=���iȖ%�b_�ﵴ�Kı=��iȖ%�bw����Kı;�>���3.f]I��M�"X�%�{��ӑ,K��{�ͧ"X�%��u�]�"X�I$X�@"C�6!�&��{�zŷ�x��x��z���GI]�&�Z�r%�bX�����Kı>��ٴ�Kı=���iȖ%�f#�ﮱm�!�.L�}VKU��X��h`@o�J�Q��ɀٕ���x)E��Z:E]�F�F&D*[i�[x��x����{6��bX�'���m9ı,K������bX�'����9ı,Q��x��mD�2�[5�o�����M�"X�%�w��ӑ,K����]�"X�%��w�ͧ""�T��w�_��T�W(���b��<DK����ӑ,K����]�"X�%��w�ͧ"X�%��w~�ND�+�<_/7[��e�v��-�-�C�bX�����Kı>��ٴ�Kı=���iȖ%���2&w���ӓ���F������[bv�X�ı,O���m9ı,O{���r%�bX��{�m9ı,O{]��r%�bX��H4�Hp%$�ʶ�E���1�,ȑd����>�/�`���n�+t�k ���c���Zå&Daq^�{Ampb������Y����3S 'X0q�ঢ়�v.��7��l��3֛d)�ۇ#\�lmº%��ʽ��ݣ���<�cj���*!&�T�XV����<���m��Z�1�T�IN5�ڐn���u�F�U%z롽f����q�8�&�Ea��#Q�A;��'��{v�}�"3G0F{r���ð��]��J��<�]ԑ#���%Aų�c��4L-��~Nı,K���6��bX�%���[ND�,K��}v�O�dKĿ�����"X�%��?��9�&e��Rj�SiȖ%�b_�ﵴ�Kı=�w�i�TȖ%�{��[ND�,K�����ND�,K�f����u�����u�o��{׾5�o�bX�����r%�bX��w��Kı/����r%�bX����%��!R�Mb��<C�<G����m�bX�'���m9ı,K������bX�'����9ı,K��}fO�[#�B۬[x��x������oı/����r%�bX�����Kı>��ٴ�Kı/����%�t��c�L���T�R�'�N� N�Qκ�[��EY���f7��F���D�,K��}��"X�%��k��ND�,K�｛� 	�L�bY���k��-�C�<C��������vF��K��m9ı,Og���r� O�H�I��"��S�ߢ}��9�iȖ%�b~����Kı/����r%�bX���$~�p�1�mT�k�!�!��wޚND�,K���6��bX�%���[ND�,K���6��bX�'�wܤ��Z����X���ff&�x������Kı/}��m9ı,Og���r%�`؟g}��r%�bX���mZ�$u�Z��o��_�ﵴ�Kı=��iȖ%�b}���iȖ%�b{�ߦӑ,K��;;>L�e�F3�U���B��V �����!If�M�2ն0����I<�C�&�Z�r%�bX�����Kı;�]��r%�bX��w��Kı/�ﵴ�Kı/OOd2K���p����]�"X�%�����ӑ,K����M�"X�%�{��ӑ,K����]�"X�%�~�o��3=��75��5�ND�,K���6��bX�%��m9� ���|���n'����9ı,N���r%�b����R�̣Z��o��{�{[ND�,K��}v��bX�'s��m9ı,O{���r%�b���v(�D���!�'����9ı,?�B>����m>�bX�'����6��bX�%��m9<C�<\\��7܄����P��=iB�e9�YZ�F�*��nnrM�����m�9dLE��K7��x��x�?~�5�m,K����M�"X�%�{�{[ND�,K���6��bX�'�wܷZ�W)jr�-�X�����y��X�%�{��[ND�,K���6��bX�'s��m9ı,N�ϭ�Ԭ�����X����w�X��ı,Og���r%�bX��wٴ�Kı=���iȖ%�bt��,-�E)h�e�ŷ�x��x�=�Mb�Kı;��iȖ%�b{�ߦӑ,K+�@�D�BD
� �9�0ȁH�aB�1��Bu*o�9�s��r%�bX����'�L�*Kl�-�C�<C��w��.D�,K���6��bX�%��m9ı,Og���r%�bX��D���ݿ����r�JŠ�,2�1T��r����f3uu���m�Bge��$���Kı?�����Kı/}�kiȖ%�b{=�fӑ,K���k�!�!�_ޗ	\s(���'"X�%�{��[ND�,K��}v��bX�'}�siȖ%�b{�ߦӑ �ɘ$�������fani7�O����ؒ	"~���7�?�{�ߦӑ,KĽ�}��"X�%�|�x�"c	EIMb��<C�<]�}ͧ"X�%��w~�ND�,K������bX�'����9ı,Oyw�
��eRQY.�m�!�/{���r%�bX��ﵴ�Kı=�w�iȖ%�bw��6��bX�&�@D$��O̹!i�j�F,�����7l�qƽ�Åw#����3�o[DV-ٮ�m�[;��6�SO��z���i�A��6�:�'Fj�\90�	P.W��e��u�s�8y'=\�\����-�Tj[��͓ڳ>�xQ��<��m��c����g���F_`�؀�tge'���"6�Z'a�偘�uq1�򹺅��)]�Q�2	��-b�$.,�经��)�|<=�,؛�JA���	r�G��ǳ�]$v�=yyn�JA�-�\ �5u��~�bX�%���[ND�,K��}v��bX�'s��m9ı,��w^zŷ�x��x��<����Z�\��kiȖ%�b{��ӑ,K��{�ͧ"X�%��w~�ND�,K��������S"X�����B\����]kZ�ND�,K�����r%�bX��w��Kı/}�kiȖ%�b{��ӑ,KĿx���3=�5[u&�Y��K��`dO��s�m9ı,K��kiȖ%�b{��ӑ,K��{�ͧ"X�%�N����p�52�9k�-�C�<C�w���-��,K��}v��bX�'s��m9ı,O{���r%�bX��k��&Fj˸���]�����ب.�KV\�
RǈD��V�HԦ�8qP_�,K����]�"X�%���}�ND�,K���6��bX�%��o�!�!�<�x򅑴�9i��Kı;�w�i�|�mخ;���'{���ND�,K������b�s��5�o��{˺��Z]h��S5��ND�,K���6��bX�%��m9��B"w�_��iȖ%�b{�^��ND�,K��=.sNB�-zŷ�x��x����Ÿ�%�b~����Kı;�w�iȖ%�bw�ߦӑ,K�韼XS�,���e�ŷ�x��x���Ÿ�%�bw��ӑ,K��}�M�"X�%�{��[ND�,K�N���g��F:ȯ�7�۩�kb7�*�9`./NsZ�"�V2�VSLBˠ��H�.��Kı;�w�iȖ%�bw�ߦӑ,KĽ�}��"X�%�����ӓ��y�����`WKMb��ı,N����r%�bX������Kı?{^��r%�bX�����P�������XЕr׬[x�KĽ����"X�%���ߦӑ,|��)	 �� �Ij-P�@��Ȟ�[��r%�bX���[x��x���n��H R�a��m9ı,O{]��r%�bX�����Kı=���iȖ%�b^�޺ŷ�x��x�.��,�:��j�9ı,N���r%�bX��w��Kı/}�kiȖ%�b{9�Mb��<C�<_r�2y�K�� �:l&a`��b͗�YI�뵶�a��X=^zΦ,pS�qB�I+�Q[,�-�C�<C���^zND�,K������bX�'����ND�,K��{6��bX�'�����9$����X����{�I�,r&D�?���ٴ�Kı=���ٴ�Kı=���iȟ�S&!�������j�iv[�[x���bg��iȖ%�bw=�fӑ,K��{�M�"X�%�{��[ND�+�<G|��b�Ƭ����b��<DK���6��bX�'���m9ı,K�w��r%�`i��D��R
.��0|����ͧ"W�x���Pz8z�D��m�ŷ��bX��w��Kı/}�kiȖ%�b{?{ٴ�Kı;�w�iȔ�S�O'��,;�,p]2a/�ț	��Ɲ+�L�[�x�ܘy6��0\9/kx���k�[&����Kı/}�kiȖ%�b{?{ٴ�Kı;�w�iȖ%�b{�ߦӑ,K������̓������!�!���5�o�ı;�w�iȖ%�b{�ߦӑ,KĽ�}��"X�%�|~��O���EZ��X���}{�X��,K���6��c�$2&D�������bX�'�w��6��bX�'O�ܾ�]���(���-�C�?�4�������Kı/�����"X�%����fӑ,K�VdOo��iȖ%�b�{�97Z$dR��Mb��<C�4��}��"X�%����fӑ,K���]�"X�%��뾻ND�,Kn�ɷ��Nb�@��@�A��#`E��bE�$$H��0 `��ge�p�cD��(� @��0�F$a�۽�D���12%�"�F[H�M��$bBw����%���3	�ċ!��`�4,����"��P�D�J	�A��kk��l�Bf�4�aE�jA����f~.IL%�jl	I�\��VKD72!��	5�f_��&a�9��@���3)UtX�IFU�JZ�MeĔ#P�2T"�#�)J-d%����D&H��B@�������iJ�_�	��j�WnÄ0��c��`��t�Ffh+��6��B��a"ȗ3f�s&��[#�	��T�iSi ���H��F�l�'�C!�YF5���HHK�iRjj \��	�M���s�tBh��؎�>C�[Mނ}J�bM}�8k�́ �ZZ��$iE�	�y�&�|s���Y�M�e��.��cS@UVԻl�S�PV�Uhk�f�X:�^:�+��a�4H�TT��֔�)�螶6z-۠ӹ���f�Az�1۝av����kl���n����������m��:����v74s��VL�m�)��x�9��d�Z�r:�ԗ�@u���=��2�;\9ؗ�� U`E�c��٫�;7�L�E���s��Tf{8�>���wP�+퓶���r��,$���;��b!eI����`ԩ���쩫
BH[]̨Ҵ���5=GmрЖ:�6�b�X�*9��X-®�u�8�&���c��GX���Y^m��z�{{�W�-�oXn�s�{u���o[�4�>L2�1��U�nx� p�tr��oo�7gv��Nul�;O�����R,�8�<�z�����ûV�g!I<���5۰��;��WXC��]:�a �Q�b1D^L�m@%̓!n����6�c�E��p-�� ��=�/kaD*b�'e�DN.��h���8<1�ڙ�ƱW���3`�)v�F<Ul���8�c@S�a׷X���./]\ȼRnfF�5���&�<�� �ٻg]q��ۅ�z8��#;Yqۍ:��'�/rN�Q9i��9��T�)�\���uV�xlޫ������dB��E"E�v�m�6��V���&x�y�u���'u1��۱��:��"v��h��
-4�u2���&bVX&C�3`P5	cZ#�M��T�8-2k����ǣ����K.eX��Ʈ�y`VK���cK\ty��9��p�0�5�t�n��٫�;���Z�؈wn�\s���ێk�mZ�C��5����'.�6�r]������qQh_UZx:�w"����乫Ѻ�Mb�R�ŝ;����h�Ɠ���)��WKF�1C9-�Q ��l�T��lu&"��sю����猝�y<!tq���ɯk -�f��ڙ˫Ab�D&�5v�Ȧr0�s�� )%����~b�Po�����F!�DU� �ۂ�П�| � P�d�P����uqR�E�e�U�d24�:9�̋m2����u2J\Ш�B!��|7s�d�u;A(��M�l��э��m'BD��V�.`�m�jZ���M4Iv ãt,͇�v�HDlJ޻]<3�qM^�V�b�[F� ��/���7�Vm �b늝����A��3r� ��\�m��9�Xl@3rd�p�1n� ��ЈT� ���t����_#�F�*�kJ���gH�vt#ŕ����[f�r�uXq�jv	�ʆ��*/�>^,K��~�iȖ%�bw��ӑ,K��u�]�"X�%�{��[NE��4yFا�� �۬[xX�%��k޻ND�,K��}v��bX�%��m9ı,K������!�#� ����h�Ye�ŷ��bX����Kı/��kiȖ?�2&D�����ӑ,K�������m�!�!q��x�F�V�妱r%�bX������Kı/�{��r%�bX�����Kı=�w�i��x��x��w�Ѓ��W0��n�r%�bX�߽�m9ı,?��o��i�Kı?��]�"X�%�}����!�!���/����D��Z�\i�1PJu������)�hnvU��'�v�2�ц,цɫqܯ�O��^�%����]�"X�%��뾻ND�,K������bX�%��{[ND��x����J��:붚ŷ�xX�'����9��6�q�Mı.��kiȖ%�b{?{ٴ�Kı=�w�iȖ%�b{���9��əf�5���r%�bX��ﵴ�Kı=����r%�bX�����Kı=�w�iȖ%�b{?z�禳,��R1�n�m�!�#����m�!���k��ND�,K��}v��bX�%���m9ı,K�B��S<�Y�k35�m9ı,O{]��r%�bX ,��]��,KĿ����ӑ,Kľ��kiȖ%�b}�������C�f�C��H�g��'k���Jm�1	v�̂B��Bd�h)�*��O��%�b{����Kı/��kiȖ%�b_~ﵰ�}"X�'�{�k�!�!�}��0pTʜD��r%�bX��ﵴ�Kı/�w��r%�bX��wٴ�Kı=�]��-�C�<C����RYX�Q%�ӑ,Kľ��kiȖ%�b{=�fӑ,x~��y�v}���˴�Kı/}�kiȖ%�b_�}��aA�]e�X���$�V$����}��"X�%���{��9ı,K�w��r%�bX�߻�m9��us�g�%%rqX[n�m�X�'�k��ND�,K������g)�U/l��==x�P2��l%�BY�Ԛփ6W]*��ʹ�F˯[Z�qũ��k��)6m��g7��޼ ��x�e��E�j�G��E�����w�v^~�s�\H&�׀{_���c��-��(��E��� N�x�`nǀv^�Ѝ��j�i+��N��xݙX��*�U�9{>x]v[�
vr�t���E� M�x]���b�>���c��:)�eق���hL�l&�\�a%��j9ip;�:�H�0��,��T�v�we�G"�'^ŀjݏ %�Q���Ybwx�`^ŀE� N�x�z�7i;,��Սݬkذ�j< ���	ױ`we1�e;i��;E۵�Eݨ�vK�'^ŀMۆ��8�n�V]�[N��엀N�� ��/��4��bX��\��ds�Wl2���/�XF�ڴ@t5�OWn��nq�d�tfM�˷����m�q4`c�3"hV��,�<��g.L����^L�����nk�����@�he�(�a�m]2��B0Ø��L�{��������@�����6Q9��+�ghS[ X�-Ci���ώ
v����%���;7<R��*�=����aU�<�[�厄����mB%�_+)��:�
��$��d��x疽9�X��sv졥j���7n]ڏ 'd��l��]��`v�Eݨ�vK�"�ǟ� �OZ�P�U`:Wv`�W� 'v^v<wnd��St6+V�E&�]����"� �ۆ Mڗ���.ӧVX�� ��<wn7j^ N�m�bK3>\�z^�$�E��E�}j���!��-�����d�d�
���m���[.���BV'v��/� Mڗ��/ ��<��M�eYv*CWf���bAS�� ��E"�,$ S��V�-��v�ut�MJN�j�[b��� 'd�.���9I{e��I��j
S(T�6*�ۻ�"�;� ��� �����t'e��c�xݸ`݅�엀E�< ӱ9v���b.��Is��rp^#'n]s<�p�nu�Xܰpjq�Sp�h����� iU8�}����� �dxݸ`IWPm�l��˪M�/ 'd�-��v�v�uJ5�Ё��ҫ����	�}��?(���U	ሎ!�v�UUͭ�޿���x҇��m*ht+Mݼn�0n��vK�"��vq����P�ա�� &�K�	ݗ�E�;�#ke�ێT�u�p��[�ףZ�W$j���|���O<�t'$�k�9gC������l�.��	ݸ`ݩx�8�2R;��w�E�}I\,nԼ ��;�F�:�Yt;M;��lۆ Mڗ��/ ��< ��ݖ�P�L��+�0nԼ ��x]��mW+�Sfa�}%]A�I��v]Rm�� N�.�x��0wj^����c����Q�^l-�\3kl���F6�X����/#�/bzœ;a�I��]&�b������N�� 'v���W�l��=���*�f�һl��޽8;�/ 'v^v<��I'�+-&$���ـ�R�we�wc�'v�|�N'ݲ�ڴ�i���/l��[<�	ݸ`�Լ ڂ�t&JV�T����dx��0nԼ ��x�r�T�v)e!��LЇ��g`h�j�c�����xrYl u�ݦ\���|]p��4f0�.�oZр3�ce�I��k	�i3َ��sufX��ȍ.�ݵ-G��6:+��#�͐Ęò����df�/,f�_v���O��Yw���A4�˰��#v���Ϩ��A�h�kLŗ:��Q��k���j��GUtr
b��Y�R����N��6|.t�Sf.��V��I�20�:��n�ۣ4s�lRl����l�-���w	�+WV�mݾ��� Mڗ��/�I%�����m|��sթ(9F�Kf Mڗ��/ �lx��3��+�������]�^ }�~xWdxz������xT5���մ1]�dx��0nԼ ��xeT�We�/��m���N�� &�K�	ݗ�E�����ui�ñqc��"�@k�OK��h�I��-PiBT��3";\�nZ\�m�4j� �θ;���#�'v�ut�N1�cQLV� ��z�I�!�@�By�(�U�� � {���3rN�p�	�R�j
qЙ)ZiS��wx]���p�&�L� ��x�H�')Z��cn��z���� ��� ��x]��}ԍt���j�C�0	�S+ 'v^dx��0��7o��Қܵ��S��JC:+)Q,B/�nf��*��RR����n� [�Kc�IS���=x�`�p�&�L��뉂C���i	���b�&�� �ڙX;%��=Q�n��:V�v�	�p�'v�V]�������2��@�M6]���dbF&�d!0��".��Ш���T'	��
flIɨ�)ȑ���d�J@'8ˁkH!��	�Mj31�l��Ѓ�Չ,�)�s�K��	I$	$��`Y	 Fbb�~��	��K.ɆH��d �i��X�ܒ�T)�Bvp!,"�A�-�+#H�6r�.�q#�q�!�M�%���z�w�Wf�^�.���T��T~@�mT>U
�����ߦ��䟻��w$�ߺ�x]'h-$��j��'v�V N�x]��	�p�>]����Z���b�u��^v<n�0	ݩ��{���[
Zk�BD�9���XZ���s�W�ǚ���Vw;�QV�m�;as��������v�N�L� �����m�'*ں�����&��=\���/e`�z��#�
����S���j�Eݘ�T��	ݗ�E�:�, �F��e��N��{g�rO~�z�I߳�n���E�$�X$#*R�THc1Ɠň�/�>ӻZm����6e�QV�+��'\� �{��2�w޼����V�B�Mm���f��5�����r�m�tv�Fܬٶ��1��!(dr$Q
趝���=x�T��	ݗ�N��;.�����j��>��V~��RAힼ���}�"�r�\�A��S~bv�V�E��)<�	�"���K���w�{+ %h�'�7�i]ـN��r,�e`�p�>ZA�`��j��wk ޹��2�͸`�E�Jʮ�.qU.XB@��I��z!6���[��i5�����sf�e�89wo/�]�a�yGs��$a+cv�o#O]�@]h�S�3������(�������6�np[֬�F1͞�om𣣝ȼ����UNDc��-�[��8��Cmk���Y�v�rv#���$�o;g�[���	�t�g��)"g�m*I[i���-b��oܵ����Q��&�[PE�wIl��VRf�b%I`��J��R�b�'��	J�h-����i[1�I�FQ;t"��t����͸`�E�o\� >��F2�e�o��wXf�0	�"�7�E�}5L�z�Z`��v2�ciـN��r,�e`��Ӏ~�7��褵�ܷ��$��߼��/e`�p�'\� �v1�V9�itr+x�}����n��	�"�;ױ`]��wWi���]�-��2V����c���hv���,0+p�L)1_�'l�n�4�'u�uvG�N�޹���^��B���'�'M��ۻx�f�j����r�ɏ�,���XV�x��7L�v��bN�`k�`MS+ �ݏ �r, ުZ��&:�����o�f#�t�֛|;�M0�r,z�X��ؓ)'�J�)$����	�"�;�"�>��V����ꚛsrz�%��U�m�hA˭Ɠd&֘�
����&�HQX�.�InR�v�	�"�;�"�>��V�����ۻ�3e�����o>��䤎�/e`��x�g��s�����>VU�tTsx�~�����p�t!!�Id�#bF,$2@��!B22�bHO�ʉ|}���~�ܓ��?�w$�}܆gc-�,��BU��bXrsޚm���4z�X�T��	�)T�B��;����N�޹��2����v����BzX��q@��a6�8ع^5�9h���oc�[hR�80�A�6���s�lIݯ���� �j�X]���E�ꥮ��eN�Eݘ�+=�W+�[�<���Mۆz�UT�v �T'V1U��;��}�N�7n�+ �vt�wv�I�x��/m�� ��� ��e`v�ʣ��H,Q�� @�) H�F.��n��ܓ�Me��j�]�Bv�ݬn�0	ݵd���{x}��rf��+K�P!5bu��F���[�2[��n72*9��n,	�r+���uvZ�0	ݵdx�`v��e7(wv��]2ڵk ��<uȰ	�p�'v�X�
U:P�6������N�7n{��s���� ��y�-*7H��۴Ɲ��&�� ���E��ʮR�߼�uR�����wB���wK��W����=��X{.y�sg����ͣsE #�`���r�cWmiyT�g�F�!��y��`Z�x6��h��g��K��Jj���}b B���7e��e3�v�֡sq���#ɫ���B{X�*$]��7&w1�\�N�-4.F2�#1��ѭ
K�O���s��&��ˎ�I��(p�dϵQ%c�֗Df+ՃعhD�0�vq�.糶���gK�����m�E�<��6�rZ(1ѵ*����2�`!Ӷ�{=��⽓H�klڱ)6���.H�$����� �r,�����9ϐw�_�iI�N�.�AI�x�g��$n��`�W� �� ���m�V�������`�`MW��<uȰ�G���uwb�0�����:�X{.��Sr���ղ�һ0���	�"�;�p�?��zpo�{�\��%kE���Y�Ď��fF���H�qR\m"�3Jŋq��ūVZ.���m��'\� �e� �j�`]��-)G@7)�n�wk �e�;_Wo�TVs��U,�\0]���;�^Y�|����M�,Lt���+�uvG�N��ˆ hP)9iU�I]�Wdx�`�`z��r�}x�6X�r��`Rn����ˆ�u\0�Ȳ��ww��e�z� Q4`�-��g�H-�X�VTKnJ�0�у��9��R��*��v��>w�� ���z�[_ �p�;��[�n�`���ـ}��`}��X�.{.Wv���v��WV+J��;�"�>�p��U�(�B$Q�A��3�w]���v�XF�U:RЮ��X���}��w��}ݷ�Uʥ�~��:�����i�awv`�`�Ur��1�|����ˆ i؜�N�Rv.�͍�&�8.1�1�]a�n�vչ�tMٶ�V��]��h\9N���u`�`l�`v\0���q]եEYI[��w�b�>�p�>�`=��:kٙ��=��E1�X�RJ`��ݗ����Xݔ7mٮы���8��8��]��O��ݻ�Ȣl ���}��'���v�ӻ�]�۵�}ݷ޽� �e� ��E�u��n��:eL,wK(9E�k�[@��zl<��z�ͷ�$'$�N�2�9�����?~����z��=�;�ٙ�-�����M����Q�)_v��\0��X��q`]����(�N2�v�]ݘ�r,����x�.ު�ȊU��4Z���}ݷ�ݏ �e� ��E�+��ԪN�R
�%e����ˆ�\� ��n,Wy]��]9��~�D��dĐ!�����#"I=�|��^	�`�B@�F�[5!6;*d�@a��}�< �ĥ4��ɜ>$q%֎O��"�WJ�������0:t�9�A�LYR@�T��[����n�)I&���F$bI�A�X��Z� b:66ZK��! ��$#C�O��4�����@�m�� B� ���7�PJ��@akH�F`@���X�FF�XI!xЌ"����0�YSF��6ĀAi�:`�b<��# B!���L3TGG ��Ѹ࿶���l@�5�m	��h"FV$ �Ԅ�a�� j"l ����n�S`�6��l����yv~�8���L^}�ޓgCuvC�0(����9$�BKd�l����O}>牲 R2�3j�TKV������e
'���B���T��Ze���7G1�Ѥ|P�P��s���N�L�q�Lj�me]�p7Ff������m[y�c<x`��-:��3�9A9�d�4S���%x�]vw���,qe�"B�,��0���ʦE�i�fv�x�y�ʴOnj�n6�x�FL�a�'��dۙ�8���k���&{*�#�!�N*�(�2D�Y�b̄Y�uR�mu�f��MJ���(9[=��$t5&o�dl��\���,U`�KDvxv`&�Dq����H�ȎOBn�A��o�x�K1%�v��q�F�����a�-�@��3��웳x�#�9�;!sJr�훓�]�-�ۣ�\D!��]ej��r��m�g#Yz{�6��vB���Omk\�.Y`(�5��Sx6�vG�Z>�T��c���׊)#]��ػ(��o!l�K�٧{�IY�˲��r&ÕgF�f	�c ����S���`��8�"[v�b�"����m��2��s�;ּ �Mf��s#�מ�ݵ�m�tܡ1�qX��`�3��N��d���ˮ���۞���M��\9i���{l�=�꧘�S��+흺M84[�e���<����jD{EF�+[UG�K�� ��uF0��6G�4�p��^5eB���y� Aэ�crz�&iF7g��4�m@�l� ��g�y���v9%�ftX���Z�ܣ-�#(������V�E���9��ݖmz��\�i���S�pXѰ��l�s���n����<vS\���@򒫗�S)�չ��D�i-
��|�o�v�#�\���Ogxy۔3�ݹ`u�)�D���ְ�#{s�Ⱥ�g�<u�%��^�9-�4��*���P�Fi6V��U\��p��rͳ�� y�����0r�.B �X�m-�m��6�a&��Gll;��xC�F8�@�Բ�vF��L]���K��zb2f�Ag�AY�2�#�9�ۢ�I:u�������P�;�ȩ��c�~6|"! 4g���V��tu�0&�ro@\�V�]��:IϞIB4��`t��3��dD�i:����wK\'l��݀cU���X���!ک�E#���ԉ����:���m����+Q7�xm@k�ƍ���q�\g]c�<�6�+�u�\���#����)�v�d��wk��;�'gh �7$��q�i�w6�]B���\3��>�� �'%q�i|�(�3�KC��[k��}��rz�c��9�f[;F�vN��N�a:FWm�v�/����gz�|�p��X��q`]���(�ܱ����ڷv`uȰ����:���l�`wg��&t�v�`wmŀuwc�>�p�>�`�YI�Wnݍ]�n��:�����}�"�>�f��J�J]%j�v���}�"�>�2��_ ;=��:�$�?����I7 -��|���@���ey�!��&lu�\vŸ��<v�Y皶�{��,��K�$� �P�;�`��F�x�{�'=�H�A�'���w$�{�ܓ���7#���5��@ߓ�����nS-��6���e�  �lyXiMH�����17wx��w^ŀ}$yX��r�.�z�o����骻-��Wv`ױ`IV�<Ip���{���cK�ZQ�b���q�[y#ip�k��n8ܠ\���E�%�z/�8�:�۵�}$yX�H�	%����9_P�w~� ���]�sr3dF��>RG���9�${޿�y`IV{�����&��5 ���}���=�?v�|(y F(�� oy�s6`/{� �D�����t��ـn�� �H����K� wT	��*Wt�iݘ�G��z����?���~0ݸ`R�`>]*M!ݫ�j��!�wUF!#M�hWey�Z����`��c��8��t5g.ۺ�>RG�M�wn�ŕ�v�Ԉ�+I�]1��xc�`�b�7�V�<vQi9B�ubWI]�v�ݸ`�ŕ�I/ ���q,�j�M��wf��YX����XR�[�(�J�@�0�v �7��}0����i�t۵J۶`��xuȰ���ٌ�7�r1�#*�۹�t�[X��j��9�z�]KMn��K�1.Ǆ��k��~�Ȱ��+ �vc0��xZF��ꔲ��m���K^X�f���ƀ7g� �ˆ v(6��H������v[� ��ǀ}��vK�	[�Z\WL�[�i�XWv<��ˆ�v�X��� ��ݻ����>�p�>�`wmŀw�b�N���B; �#��)�Y�$!�[d�P`�i�s�Ŗ����JMr-����˧5�n��u�gc[9���J=���99Ƌ�b�L[�:�k��5!#UWL���� 
p46�ж��YͪL
%M�4ս�H�yW���ULgd���\�Ue����6���g݄+9"b�I���ٓj1ٔ�l��N�w:学<��tm�:�7G$�Ӥ�I�'��w��rr.��+!
(�Ѵ�9���OvƁLW�Qe��0���*�����k�o����M���� ��b�+��\0?��*{�BU�T�m�V���[��W9��$w\��;�_=6��/^��@�9ܒOW) �(�V�`�<���`wn۶���(����Ye�� �9�v�}�n,r�U�-ٞ0�y�����-�N��v\0�mŀw�p�?�{��?{5,�jT4�Ʉʱ�k"��s�E��ݎ��������4��Yv��.�!+�0�mŀw�p�>[#�;ŀ���:e���SM��7���W9�UUSgV�x�"�>�ۗ�~��l�҅¹f3�����pǱa�r��we�,o�����5)[X��X����b�>�ۋ �ˆ�<V��'�t�4�eڷk �u\0ro���uOy��b�5j��� s�H��Fn��֧�<�����d�2X����U���\l,tf���<��X��p�	�(����Yv���>RG�v=� �u\0�`-"m0nYN���k7$����rN}��p�D`�A�V@��Hd1�@CB�����r,-J��ut]�"��`wU� �������, �B����'V��;0�%�-���b�;�.{�k�V�]_,�z��Y��〣G��;ut\s�aVq;F����K6�ª�l��?�������p�mE����;�V���e
��xu�Y�H��^X��^�ݏ �$�ʺj��e�Wf�v�X�����Xf�0[�M���$�իX�s��S}��;��;6ea?H�H,�"��I��|�G������ݯIf�n�l9x��,�fV�v�X����i]�5Mf�"�nNɱ��T�N	봔^�g�x6쎷Y�1AlZ��; �ٕ�}ݵ��<�{��Ll'���%B����q`�#�>ױ`�2���W+��"���un���`o����Xc�`�ۋ �Z��lL�ۦ5ww�}�b�69�v�X��r�II�^�J����;(TXYv�`�E�w�n, ݒ���X��*��᱖m�]����ج�V7<�Ȥ�km�2^�%�C,n�.����l5b���J����jA	�����عϬ@3rY��n��v��u ��z�K�8I��k6Иl))a��%�dfݻtG]��;m��KX��u� 8�2w=�L���bgbg[؍f%��m�8�Җ�f����#�f��4 Pq��	�ݿ[����ˮ]����[�i�#t\^G�/w��������3��N���wp�v kp	כ�m���$s�N+y�&8�n���62����>����^��ٷWw�������vӻ�엀}�"�;6e`.���j�Z�t��V�V6[��>�`�2��V���/ �t��hnYW`�Vݬf̬��e��/ ��� �q�m���.ؕ
���^ I����0	6e`
�ԥ?�!�Z-�w�l���������s�c��r�6{u��z	|Uo�y�tt�\���r��ϧ �۫W˻x�8�T�bv�t�oZ�䟾����Q�����L���rN.���l��\�G}�?Quw|h.��wf�Oe`ul� �e�ױ`�N1<���&�Z����^ I���ذ=U��O}X�N&��;��������vK�7�b�&ɕ�E��x���Sg6]U�e�`<s�KZ��U��60K��b�����0t�����V:j����0�e`�x�#�>ZF�7,���ӵ�l�+ &ꗀj�<�r,��T�D�v�%E�� ��^�Ȱ��+���C�a�RH@�a		!$BLo��ޟci>�΍ k��݅!�9l���5p�&�#T�$uh��#���(4��HC�� Q	���F�HuYy�)`��s���$X}�p�K����@�}�[t@�0�B!Xa*��bBp���:�։Sf�y���1�X�<�b:۾�ω���u�y0���XGF��$XрE�	��B		B2,� HU� �vR0!B&����	C	��f���p	E�k}J�iH��t�E�/� �c"��\T��j	XR�����~!HR�%����!�a�X䭡�CZZ��"m��e#B T����ԛ��! D���ߨ5�v}7�RotI�|}� @�5)31MU2+�nvr�>;/za�Z������Q%�u�doBf^I: b�?_�����~*||�ы��b�G~�]�pᩳl$'e��9Y��!��pzB� 3!XZ�A� ؠ�C��?"b��A�#�Дzh T���W�t_��"����_f����ܒu����q>;���ڻ��)������$�Ur��Kd^��kʓln������>Sc��^ wuK�6K���{E��*�ّ�a���Txs�y�c�OlW�ᕥH���	t�kCFᕊ���wo 6Ix��/ �.�9ϐuzy����I�]�$�2ۻ����x�p�>Sc��^{�Hճ���+����U�;�{�� �M� 6Ix���^ {���zK.����T�)��%� >�e�_9�Z�R�(�*�X!�9믽7$��{2��e]Ьiݼd�`�l�d�`.��s���$M��V�:�UIEq֓��N)]�Ɍ�:�$͚ť�\�˛.�Yv�`�KEO�����	%� �9�ʯ�{޿�H�w��TDW���6��޽{333?�=�M�O_����h�҉���i�N�`G"�&ˆ��r�	�E�}6%۲�"݉����I���ώ�E=x�"�>�b�6q����"� �j�x�"�>�b�&��ܓ��$ �U	�gs&v\���4�3Ϧ�p�/OI�� �����m�eD�1��.1���hq��a��ʍ���������������[�]��̏\��kٙۅg���݂��7`��F?Q���W
[��'���U��ں3������Zp�q�b���)��S ¦x��ۍx�L�pr�K�h�x.�F`�q���ւ��l��I����E�]i��Uw��|5sZ�\�qӎ��h�P9'�X����w�㱇י0g�8�V��X�#"�BT�-�w���,��,l�X�V���kj�:�lv��x�ذ	�e`(�^���$ui�t���*m������?�o�xRG�N�� ��&8QeҶВwk �E���� �{#�`�V˾[�:,�i��I:�,G"�>Ql��zܤ�HN�캿�W�%�/�����#��^��^ܴ^3d%j��c�����:l��|ݿ����H�X�-��E�< �N$�5n˱>;V�������ρ $Ea�����(�^��v<a'o*� J�n���e�l� ��5Ȱ��&���0��*-�w�E�<.�xױ`��x�Z��:N�[N��۵�Eݏ ��X�6^5Ȱ��s�\��^~mZ���y�$�]T���hb�������Y�o`u%�g�-�Zm��+b��l���������o ��X]�����_-U�ة$���e�%� �{�Ȱxn�|��i�-q4����N��s��X�P<�����7�g<�����h֊6�M��-;� �{�Ȱ�[/ �.�����.�|v��X�E�z���z�����'^ŀN��ۺi�Ut�lk.	��Sh+��n�:�8�J2���a�4��vb���U����׀w�zp	ױ`9 w��nP��Rv�[N� �\0	ױ`9�e����)Se�v�(.��'^ŀI.�-��I.ˤi���;i:IݬIp�>Ql�Ip���TWTD�P���,ň��H2HH�F BH�	�_��8�ɋ ޸�7R�j��j����>Z�^�\0�ذ��z��~S�7FÆ�ݦ{)�B�m�
$j,D�h�f��mc�ޛ�1���O�N�����}ŀl�+ܮs���uE=x`��I؝'˻�x��X�2�����E6<�9ʪ�$���$ݗb|wmݬޞ��>Z�^���ذ�'o*�T諶���ղ�Sc�'^ŀlٕ����%tP���w�j�:�,f̬��������(Z���V����8B�\�ͮ�����GkӞ��a��86�8y�@�DI��E�%�����sy3�I�[ǳ���i�91w	�ɡ�X�#�ù��D%7\h�n���8ƨ�UQ���@e�4�L+bP~ۃ���b�G���n^\�h3�]����'�`��g%�I�e���㍭�W&���%��;0�dI���[�l��I{TyY(�u�5�p@V��e͙YI��Z�@��6Q��Q�n��u��������7nivD���*N�[�aCWo�z?E�lٕ�|��x���- �1(�S������7�e`)%��6<G"�;j�dUj�`�I]��]��b�$r, ��x�7e�[�X�Z\���6<G"�엀|��x�ւ�
���'˻�x�E�6^����/ ���r�����Ե���圱�K!uk��;�#/yv 2��'B���<�ݕ����m��߯ �H��͗�l{�")��X�r������2I�$��V�F
1 �T�/O^�~� 6l����7(Ҥ��ۻ��/ ��, ٲ���/ �Mj
��I��U����b�6m� �l�x�e��PN���U��;��oe� �l�xٲ��E�ltPl��c��ӷT�����!ԩ�c]��5۝�<���ZOf ���j�N��M[��|�K� ��x�"�7�E��v7�t�j�3����͗�lr,z�X�v]���%@ݤ�>;���;� ޽���p�` ���߻�nI9���䓿�c�ڲ�'L����ov�|�˼ �l�k�`�"��Sb���˻0��w�I/ ��X��0s��'������\`5Hi�\�AR�Z#�/N����"w=� U�r�$�;'�7��m	������ ��X��0��w�j�lq*N�!ݲ�'w�Mr,wn7j^ }$�z�	�R�.�t��X��0nԼ ���	�"�;�4�N��ۥ��ـv��엀N�:5P��B�EQ�Fcd!����lBIj%DR#@Z��l�Z)K$��,$$
�(���U\�d��, �b�[�[V�6�� 'd�uȰ	�b�	��=���ͽ-�D2Fܷ��8Q���=`�u3��8�@���N8)W��32��X���mt�������5�X7ax;%��kJj�Ь�Xݸ`݅��K�&�ݒ��cJ�n�L�� &�W�I/ ��X9�צ���H'PȤQ[aU�~Y���}�^���n�� &�W�j�rb"�$�N��6��ޚm�ؖf.����I;��$�߿krO�W��W��DAU��DAU�"
����*��" ���� ���(���� � *� ��E��D�"ŀ�D��A��B���� *��(��*"
���D_�U|� ��W������"
����*��" �������""
��QU~QU�b��L��q����� � ���fO� �~� _mR��@]����z�n��]h�n��W�de� ݺ����.�kTS���s�@9\����M�I�       @  %)��5��  �
 P   4Ј �(R�H@P��    �J�606� +A�������fzw�<�=�ma������o ���`��z���o@��=j8{|��7���aϷ���Ϊ{�>��>��}�_{�!��T�o}�G��2C��������n��ϱ����w��  7�� ���ڔ ��Z�(��|�=�|C�=�����U|�=�U�^�W�E]���;׭>�;�����u�gW|��KnϏ���ut��h  �or��}�#p�e)�3�7�t;��>����q�]�����p���O��� [��aB!��L�F�|N��k_
]���{��{�����J���}���|,{�Ny����>�[7���{w�� �n���l���͌�z{}w�ݎ�&����R����p��6>C��v�y�O   7=  �(b�l���=�&%����料�C����iJ�pzR��Ѧ�� ��GM��R�M/3�@�:zR�/F��Ӽ�C�i�0  Ҟ� ��Ҕ�׬��ǥ)�s@��Oz� ���ݑDێ��K� l�E���Y�J   V�*���kkU*�( ��ӭ��pt�����@җ�Κ/{�:_}����������`n�#���g ��)�@�[�a�a�  �w��}9���ylv�w�Y����3졞��2p���t;�px_>��� j~��ڔ�M� "{J�~�4   i�R�O��&�@�He)P  y$�R�  �!JH� h�OQ>?�����o�:����2O��k��9��@U~j��UUЊ"*��UU�aTW�*�*�EO?~�p���S)��+��HҐ�M"�i#cC1M,3R�i!������>��V���ר[VWs�[F����x.,�_}��o;�R�ߗP!*�/��v���%_r���[��H}-�߲�m���<���I6�����bF2���Č#�	phZ��xr�i�S5:��g;������\��*�)���2�@��o���E|��Hb]�x��tO�ޱ�|�]�LNƨH#E���|����h��`�RI�s[ߜٸ�m�X㣛���5y'��n{�o�4�F�8��F�M���s�c5/4nE�[ŧ�ל%e��.1�	!B0���!#ƛ8�G�	O@��/�7�}��Ѯ��K��x���[�}��6�!	۫Ȓ)����� |���_�zfhG��}���%�.��~|B眛ۤ$XJsZ�J�n����{�������'�Ms��\��\><�aO]Jh���a��<��:�b���i��_,�[B��5��Z$����B��	��5��|h�����.3=n���s1���֏m!���	�}����sA#��Bh"Q�3�����<�R��y'���3~�OIq8h�#����8��k>�k!���B $�q��8 H@�m�\��c�<8�.G}�(@�	E�!G���0�27z m09��,�	L!�X�Ѿ��cieBa�rBl���yh|p0�syK��&�ݾ��)���j`B�3ϴ±���c��M{�ɽ�HK�rs˷���nw����D�|Q%x�΢�jܮ�����3��oS���}Y�.$������p����J��;:Wkr��"����n��u�W���z���U��5�w��]��߇��(�Fh��ƌ�ňĀD � E�4��Y�ק��|x�!Od H��0���a��1�B�@���"�)��"JbK�H�5!q�B,�@�@�M$F*���$�F0�Y�.F�a�i	 ��d�.d���T�XF����I
��j���n���=�鄐���%L���	s�a~���f�������qё��P��ܼ�w��]y��&������s|�|[_n�����jOj.s����O3sU�����lF�[>}xϾ�{�8;=x��
���$bS4o�M��jHw�So~�=�RqcH]<F1QƁ����v^E�BԲ.Dha � Ĥ��ݻ��k�˭,d�����H<OJow\h���zvM�.Xk�l��Y��e�
@�3s�q5���J���5���ҷ>Y��X�5��ĕ�büO���) @��g���ra24a��m�g���D�}p�����i�q��fU�o(o7/�Zǻ��P���G/�=���6��o;���s�-hϑ[ܥ�X��������}x�H|[��|jFR_��C�Ż��@?����d.��G�1<|��u㼵}�x���/��[��8��}	
f�X@�\\I�i4a��p�
�٘i"��L)��,��k�<���0��BJ�F	�W4Ca�'�P���YB��]�؝_uc_*Y������sw�����+��N<�t�v�"����Q�8k�*\�kG�<)齞觺5�+��>�<�3~�1�����p��� T�Q��h�԰U�q`��i�g���i�>/����n"��@�} ��N�5�5��3G	��4:׌l�)�I .���}����+3!�Y5I��aan�l���`�M����!��$S�pWռޫ�b�_/�:�Yn���}}�K�T��s��z�h��ո�5�K�^R-�ŗq�u���zO	���B�w��
�h��k-��z_X]{ƾ=�0�n���<�7�	vo�|�O�&��OP�8W(B�DEe�4� %o'Wؐ�@� ��"���!w��o�����!V�Av䏽 Nw�§�Op��xB�
����0�Kv	�Bn���x���>][� ��i
��a�������sD��dֶ���
0�,�a� I��oZ��q��*ābˆ=�}�e8���7Hn�,ņg����^��@���nv��Pt49�;��8�b�!7�5�䄧ן5�5���pH�!�����f!}����Ԧ�ABn�d I\�W�'f�B8&���Lø��]+W�BUc��������!��Wp�@�F��!"R�kl0)��S�f���1����[}��vz{L��%	O��#\t]o�˖]y9��fdь	��$J'�D�_&&q�Q�@#HЅ�eҋ���/��<�!:P�-%�؞杞}xp�G$7��BR|�WǱw�#�%I	�W�:����W)"S!p.xL��ﳞ�5$�O7�<a0�y�$���#94zNL͚���`V5cL	L%��y��	<�jOw8h�H�`B�Y���Is[=fo�y�aq8I
fI��dz��u5.�\Bk��uW0�<��<毺���8:3�4��.@��5�!H�����q2Ac## �!$���P��# ���|D�����-a�@��`��D����$HI 343jA*E��`V��<e�[8S�5�a��$��X�,X�!�&phf.W	� �EV����k�/�ft�����}WZ[SZ�����+��h��]���k��S75�k�9��٭�g٣d�1�ۚw	0�ꐁ �3ܓf��f�6O���Z!Fdd� �}��a�Ͽ�e�ذ�!K���B��i�o�ˎ��F`�%I4�1vcI�uybuy��7{:kVN�T���'��F�����g�8&�>�➞���p���4v���{�]�x�M7��I� �	%>f4��#F����)���\4h��X�� SSh���y�|��c�K̗2��1��T�aD��[�~�BH�#RX�����K�b���)���B�!��#�$���P1�X�i�q���e�\}jAivĆ̜7��d��ee>����d[�l$�c2M<���(쌉	�yy��$���a|�3F�I�$B��Xˠ�@���(������>ϑ!���q��b$�
�F��y��q���nkF͞ A���l����1	����S�����>�p������}kV�g���0ѷf�d�����f�\ee5y)al�,�nD�]�����s$�K�{��GWl�f�ѧF��}�!!H�Tg�<U|L���tp�����>��
4���'�77��O�<��C�$�s��3���<NY3�\	�	{$�i�ܬ%JRq!d��kӛ�n��\��o|��nC�=C�gC�]h�x��R:W��.}�s5��Y��p�oa�!Ye�8kX�a�je���y�s\w'&�����<��4XR����<�����^_ik���y���I	��}ewl�W~�F�s��k=׼�^6���[��^���l�i�g�{Ϩ֮�4�/��Ǹ�G���{u��!Tr�:�G|�r�ێ��O/̹gY!\HV7&�7��əa.��lӇ�!RC$/5���nsyf�<��-��3���Y��[V(�3�u�*�e>p_y%�!)�7��َ���rCd����[ϭ]����Ը�b�
w�O�cs;'����6|�굋�:J�'\;Vǋ�:�;�W3�e�V�XѕOeIY�SY���ݞ�1,��z�2�i�$'��4ƞ��/���.k6L��߳�=���3A.�kX_Lw��Sŗ4�+�P������.�Qw]V��*��N�vϟ��H� G��<�%��G��|u>\+!ȄR�g������/٭������sÇ9��>x���ۭ�M�p�ꉏ�w��	����^�uiwP����x��jj>�3ɧЁL/��z���5��}�hF��BF��}�!�O�i7�J�l-��ݼm�r�MU�Ϩ/�۽ߋ�ws��W�	�	�L�\H\1���H�#G�f��	���:v�M�����7�0ߞl���bD��@���������L���*������B�h!2��1�!p�a�o~ՅqW8b��	>*Ϗ�;8Bd]�MS��s��9>��\�s��g�$bHB��S9��iÉ�RS^�/kۮ��N��e��:0$Jr���L�[a���/_:e�ԯ���O~�Tk�U��A߹:�$�p������Qu}O��V�˨�Ѩ)���_s��f�.�GDjE�,XRK�S�H\m�7�a�]���n�7���9��1�]kx<.m8E� g�5�x�^i%I0ַ�
��0�r7[�;��Ym�i��Ś�ў'�#�>�
��ﺍ���f�+���&p�{�μWE��=@�%߃�f}�S�q�E�|�����X���>|K�:|�_�}S�7A��߆��d�������`Q��
%�	��!@�nj���3�Á�_o˯����6�[e���G.�]����n��E_�>ϴ�ڱP�!���X�tI���V5j�<�C9��!�Q����NL��$l�
���ޚ진	���z�|�� �9F���9�z�^����$Yg�פ9s��<�%*J�Z�<����ʑ�C��th�$��9�<vrp|�D��E�
�`0��! ��D!X0�msaF�:B�c`U�T$q4Ja�H��QX�""W�f���,p��J�&1��1�.�4�a�l�YM k��7�9��9&��Mj�Fۯ�G�+��P��tO�������č�
��|vJ���]J��^e�s�*������}�0de���|��Me����ߖ�۵�+E�X距掺��V|���i	���g;V+�ڷE�Ӓs�c��C���}\��D.:m� �K���ϻ�5�q�E7���v�Th��_*��N��u��Ed�d��9�XS��/�+�֪��I�Z�x�C�80�k �_��v��<��3��i<L���o7�8JoO!��MƓY�F ���d��d�gAH�m�f�X[�֎sz�	9	���|���ϗ]>��|�����}��T����۞��.o�Y�w��$�\��=��Jdu��cCz�`h�Sux��U���wx���-�N.v,��v���5���48}'<�!��q�3�9x�*}x��s��=���Z�AۥY[��������s������]�ed�C�]�6�{��}�r�絒���y����vI$�I$m�2 �rI$�T�UUR�J�UT�UUU@UUUU*�]UUUUUUUV�@UUUUUUR�U*�UUUUUUUUUUTTUUUUUUT�UUUUU�������"��J�Xc��m���m43"	5 z��nu���q�2��[R��t[.���mڼ��P1��ZE��d�*�UUU���[V��Uj��j���U)����c�A����l@U�-����*��v�6z�ۑ��Y�z^֖"�|���Ϲ틸���D.dzY(�5R�UUP��UUUUV*��� A����v�����L�ڦ����W�6��*�ں��ګ�j�4jj���ܭR�UT��E@�����*�LA�W*�T�F�YZڔ(�O5*�Q�U;s�K*���[]PqV�)-UBC��]M�ڣ�����bڪ�����Z��*��UuQ������V�MO+m+�����
Q��ڧVEt)!Il��UUmS��6��J&���UU[�r��v�vm�<Eֈ)j���b-�aj��g&��$�m!��=���qcT5�[,7T�5U�?|*��H
�m�T2(R����Cb�-Yت��gn�0TRL[�W�*��1EU(�h�m��v2J�M���
��z��ڀq��=��Ӗ�������W����U�u�/n]�����(�
ڪS�{��U�.���VF5UUUP&��Sa�a+@��ڬҶ�]����
8���
��ҭUS�;WR��I�r�2NH6!i��V]�J��M�I�=��#�ti	�J�����!�������x1��a%K�\Y皪��Mu�lSb����b�V�IJ�N�V;�U��sn�c�1c,�m�ǯk�`�rZQw����{6��/]���;p�v�� ���#�v%��9�#���Z�ъY��n,���p-�70r�ݰ]U��Ts��Fv����-UUjƖ��5��M�#�A��lK0�WqWj�c���[�c��(`�u�UUU����&��Mu*�GӖ���ȭ!����X����U��*��+/6�Tp]�Utۭ� ����P����7M�ꮹ���lWUU�n��P���pc[.h�=���UU��뭶�]Ùj�de[0�4��b�-�4յeW�Yٍ���ʅ\��@J�<��]r���V��B�U]Z���N��*�V֢1B�T�Y�s�UUԑ��#h���.��Tkl�j��U�+�ڴ�K�eZ�+ƶ@
����"Z���*������UH������T�d��n)l��՟^8���)k^�!���*|dBԘ�ku,§����j�mܭ�YO�K�[�
���@H�j�YP9�FW�l��5Jꚪ����=�@���`/���,XUlk�M����-�c�.�5s����C���c`em������K����^Z|�o`x�l�ͼ�G8�S$u��#��-s��,�U�^��J���I�����v�����	4e�ϖ�+�bx4�"�\-�6����=���qۙV]�2@Sn�w\�@��^��.H{ZۭM��qN��SD��P
�
N8�4Q���s��0�B9`��mۉ���OR���̎ۑ�b�ۚ���&����u�q9���i}Qe۷)��'GE�*�T��j4s ޕ�Bp�]U凂��uKT�G]�4A�uUpۗ�]�l$m]�v����LU����������pm�����[񓰍F�P-Vl��i�r�[`e(u(�-����B��2��V���7'c(q](�&@�j���:�	�Yʫk�0.�W����,r���J��M�:{���k��t%��5ֻ�/m�Yy���oSUT�K� qR�R��a��� f�UUV1q2@R;���rp�5-N��yj��^�������۞�OUV7luUqE�U]��%j���:e�8監b�x$
%r�����b9 ���6�-Ȫ��	hڴ�e�g!�H�B�[�y9�ع�W̜܃Uc4uKI������QV�6m�hZ�\b�\i�:&�E�P��T8�x�3n�\�ڝ�UUݰ�B>����eܹ�m���Q�r;-� n���d�b�Z��tΉP$ҍ�Ky�l�Di��L
m5umV����ݭ�&�(�,4�XkȬb�(��-:�F��UUOe��
��m��c����a��v�(���=@OJ�nk�r�2���Β�9��w�v ��x�M���*�$г�;F��� <,�L���x�s��[Nrd

���3U\��ڧ��7G@�9�����9����E
�.M�5��M�;s5��A�l��U���uA���t(��
⊀�C:�\�U�1UVb�-���*@C,�U]���] �MA�3q�q�����d'֪�i^�
wX�<�mUU/-�u��0ձ��  �j�G�J��C�K�O$�ګ����2��^@pl�PlUK�O]�>+)r���ҭU}U�T�@mWO; �T�UUTm(u��WX����[Mۍ���{$ac:�e�Ij�������\t4��\����L��UR�;.P�[Uq\�UZ�]b��*A3��t���&�Q�1��fۅU`@͋�, 
��;fV����f�L��y�eXK`朴�2�GnFj���H=�R�2�g`
]\�K;l�2S�ӓ�Z�?�:��
vx�lE�UU�n&7Xx���=���eϮM�ڬg0�m;�b�j��4.Ͷ���ZݻKu�N1���uF&���E�[��B�2u$ Hf�ùP�ɦ �n��V�ǫt�m΃6+q�쩎!����؀��^X
�]���gg�[i;S�ʜx��ǹN]q� ��V�؞jڥ_VҨ@U�j���:0���;;12������ɻi�v�!�2j4i�p��b��UV*��X��H�ݚ�Z��s�(,�����
	�C��j�����K��b��N#����WKj�lb��U%Z�Y�D�
�UT@80rG#Aї�0�7l����5f����N��Nw�n[B�e�t��о�-�)��#�YW��"��;<�����]c�;���g(3J�I�E�)�ЬD��P1ۆB	Tb�M�m����k�b��9�mʗp�6����#؃.X���N{M��������VCv۬UKTc��Xut�+ϑrK@���H!pO�ն̲�\2�� ��oQmgz(�a��nx�v��:����n�SGKp��a��H�մO'd3�;�GX����l��#�w
ŝ�WhKl���ꪝ�n�OX�| 6���c��Ar]�&��j�O�6��j�W�ɔ:�Rr�mF���)6������������v�NP�ܬsɶQ�Ek6-ö^�e4�U@��l���&�`*��4 �����!�kl[&2�k��l��@J�W+�݇��[UUғ�j��F�.1ۥӢق8:�����[/ۊ����*�U
�(�����ܫ:��j��ζ��
���������������������
Z�
� خ�ZA�m��]��PAPU�F:m�5���Y�U�Z���Z�V���j�S4�����w׼�ly�M,;
�u�!�hw��|g|�t��By�MU[UmUR�T��յ D���*�6A3Ȫ�D�m{jV���{l�����h���*��UU����U�(Z���X����3�V���%#�� ��ܪs�)m���Xt2�UT��=@UUUUWU[P�UUWUv�UU@V�mN�j�GPr�*�PJ��m�z��[���kj�WH�z�k��e�R����(s�i�^��,	X��&C��������qV�m�fWf�jU����U�q� ��U*��T�UUUUJHUU�)��cp6��v�v�۲�O!��	�(Y��zש���j5UUK���UR�UU])�u&�J�5գU҆�]�D��*�PS��Tٶ�Ÿei�ΉT-������W\�땶�U�(*�F� ��j�UU!��]TQ�ݶ55Um�WU[J�UWPU[UV��z��V��Լ�':�(�����s���2 ��Uy�ՌU����J��[]UJ��V�J�UU*�q'+k�L"r�v��*�����Ym-b��ձm&�Ҷ���Z��eeQ�Z�媪�RӘ���ʮ��u��W.Z�
��j���� 
�)zy7i<�F���\UP-ڜ�4J��EUPUUUu@PTUmPPV�[(ۜ���m UUm����*��ڶ��3�W�_i��F�6���K�m��w�ܵJ��,\�\��R�5�UU@U*ʵP�D��=���b��5�U*h�'[�T��1��AU�][utb�U궪�Z���>��yv��.�i�"���U�6�ab�@$��<�-ڪ�������T@�W��t�[W �a���]��x��;[Xl��nG��Kn�b���7j�V�&��B\��$��6w] =u�S�`�mgq�J������[w��CUUJ�*r�j�#"l�K< uJ�V6��.��$�*�\gny�����Z��lJ�F�ꮇ KUR��\��)�UTP��J⪮���� �� �j����UuUUP��UP�UJ�UUPPQ�wT��!ݲ�i���j�Dv*�Lr���j�g`A����VÖ�{�r�T�ɻm��V�N�T�1j�ʵ[g��!������m�n-W�}�lU`�Z���	�pp�.�\뗳d��ޏX�[DeܵU/T#�˞�st\��3�mu�7G�T:�i: ]�۳�KD��#�^N����UmUU�V1Ub�Bw`�*1ƭ�N�������UDU?(�h��T0�m��b�H  2@O�:;X;��������Dبx�R:�< 4zz�!~T�P1Ei���^�m���;�� x�����ҁ�8C�H�"(x���@��L���4&��qEHLxpP~
���>h �P�ٰ�lX�T�����@ z�m#�x� ��H
�P�U~ڊ�С�0�}���k��N�z�	�Q=�N�|W�Q�	�6�S��|�;�џ��z�#�4"$E� }_�A��}�M�7fR�tOC %J��M�*=*'�&�_>��A� M:D_T�EGh(hPx�z��D"�|�� ��M*�<+�B� HF$& �EH ���PD6�4U�Oj"@AA���>*�]�b��V"HXT$�P�I
�a�٠�%O��O@>@o�V�!#*��E-�0c!�6(>
x��"��> �E=`@�@�u �CA�v���@>:|� 	�M@�dH���*���t$��R�Q
�����j� �j�@���e�V"(QlA�AX���@H������Uġ)K��j��r�s�8:냍�� i�nM�g'\uqiCB��ú�N�n	`�P;��.�q{�T���<ͣT�:�4�q��˄��ۄ��<�;D��Ijf�'-h�-�[A�nR�����Vؙ��X쏍�������h�E���e�M� 笤NT�q��͏�2;�kk���f����cBٮU4�oq�J������X�@>�A�xW�1�V\�L9�W;��/mU��9��N�M�l�0O]\�й]VzR͓�u8X�a���a5q�K�I���lgj�j�<�̰%Y���S����歍�ݒꚸ���l����goO�^a�Wf0L.�b���K�y3�mN�U�fqde�Y0��[��� ��ԯ���$kY�m����(�����L�i��+�iYT�0m�&F��D�6%$\�#]r���iI�т��E6�a�f3C7"%\%pځ�ی�;k�+��9;d�y,�:��a����s���8t {Ta6������2e4sm^w9��. Q\�;�� ��cI��vE_'!��x��"�-e�0��3��ePƹԮ�1@��bF�u��2�9ݞ����S��vdW�6v�+Ǳ̎�&�M���;�e���6�x��k���p�f�i��ڛ#��v��w7⃎��\���(G'����q�\��.��g��#�M�ᙰ=�cq��U*��#����
UZByNv�c�s����H����a`�Yh�[!=E�0B�5��g��jz�]2�#��$��FQy��uelm���ȈE
�X��g�Zj�҅s[m��<qp����`5ґ�H�d�)<��5�e�å�Q�G���vDl�@�WP�<� �E�eĶ��.��
�d��%� ڃ��v�;k'1Z�3��P�Qq=N��pX�帡�&V�<�i7��WI��4t@e{Mڸ�G=]k�F����a�d��I?�~U�U�Q �
��������@�>D�׺I�����lD�f�V�4R�y�F.�qk^$�/n �r���Y.�ɹ�{��b]L�ۛ�vi�)H\V���ð59��w�RV簗��6ɡk=�ɍ�e�٤�m�l� ���mmj���k+��ة6��^�6�]���<`@�����D&�"b7�֖]^� �1"k�&ʕe�z�s ���BǬKf�ֲ�u�V��B��;.ÙsH%%N��D-XV�+�r㱶L��}�L��.�Б�Y�6��Ձ�k���LX�vP�*�iШ�ݼ ��xv�<�&,zT� �T��8ꪧ,`��� ��ǀ}6b�7�H�{��	�FbݺwI�v�U��ً ޕ#����:�e`�(l���wB�J��`Ҥx��x^���d� ����l�ĩ�ʆ�y�#�sE!v35DN�IvaQ�R��`��<Z��	�v���x^��ً ޕ#�����n�uc�WWw�<���o�x)Q/��"�z��7�+c����	�f;v�[Z�v��]��vb�7�H���8�ٻ=x�=X�8(��ʺB`2��`Ҥx���vV�dŀ|�eb�j������e�{���&,z_}|����۫e�a�-�[�`�����1�rE��9���5�̡B�iD+7&�`��2�]�������Ԏ���v^&�ƭ�B�Mݺ����q�g�Xe{� >ݗ�wkc�qq6G'��v��)ҧV���� }�/��(D�"	bA$cb)$F$�Hk^���ܓ�=�f䓛��WUV�`���V�{����<�&,}r�k�6wt�Eݎ�U]�ݭ� �I� �e� 7�/ �?�Y>�,}a,�cR[+uXV����Q����D.�0��fjnܖ�	��ሂ��v����Ob�>ڑ��e�����ࣺ�ʺBb��X�.�qq��=xʞx�f,��)v��Lӻx��x��=�s�UW}=� ��<��N]0S'(`��� �ݕ�}6b�>���Nq$�És��.s�%�v�}x�E�M[.��wm���ً �Vǀ�/ �ݕ�������XM@R�e��t�7k�'��[\�k���Ѵ�ū�|���3�s�wVʪ��J��we�������;=�X�z#�uUm�U�˻x��x��x�&,�[�׮4;��V�˺E]� ov^����� ;ݒ�9��7BBT�Hԉ�,� 
��x�;��� }�/ 7v^6�wV�V�:�0�H���x��XI�0�%���t���$��NQJ%��4������� 7+<l3'���&�u�В�
ۜ��E�%	��uɹ�!iE��]�u���؀�\Ɣ�v�j�>խ�[vk��`�b�E�NX�Q˻�u�kmݭ�/SR�@�١/bm��؈���e#O�}�|�v	kRt�/[��/��Vp�	v)���d����MNY�.*Y��&.���%�G��_�Ж�a3��
vZ�)L�,�k��8F�+v�(Q�<l�F���B�wN����� ��x۷����#�7�q�`��9CWx��X۷�R< �v^6ƋWV�C�.�� �v�}*G�n��ݗ�!n���]6�������qZ�A��w��< �z�we�>?��0�uGv��V���˻x��x��X�nҤx����e<��������U�qn�C�A�@�U���l�գ>�H�Pg��=��[m��=x�n�H��$��`M��E<nB���.8ԒY'���o��"�H��l����,a���$�X"BTXJ6��"�$F"� �R�K	Q�)��'9/3�]�'�{�nI>�e��7i�Kt�N�1�1�Y�Nԏ 7v^6M�x�\0���1�]�P��v�<���=x�=x�.�H��v�
��	Rc���	�/ |�fC�'jG�ݗ�N=�P�p�/�x���4��GV��\�B:�:�${R�m!��Z��[k	nSz�{.�H��e������5�SN�:�0�H�͆���$��}��
`U�vձ�Zn��`���;��� B\�IdH�鼜6I���d���,EG*B�q����[��� �앀n��&���(HJpBԒI�y�L6I��c�C��xv�<^��⺺wtE6���ζW�Vex������uחK�Q#L!>tv;S�bwCi��π��+ ;ݗ�n�ǀ}�p�>k�q�Kwwg);.����y�l�S� ����>se`�q�|�J��Rcuw�okc�;�p�>se`{%�5ňB*Ս��U]�4�ِ�>{�����/����(T�i
��=P4��$������=��U�74mK��|�e`�\\{���\���� ��4���B]�4�&�S84��:�A��(��:5۩g���^�h��UUwu�엀}����`=����ՋJF���a�%�{��VRi6w��|�J�5͕�H�v5v��n��ݼf�0���se`���>�)����&�՘�IX��������`5بr�����'e���l�v�<f�0�����G8�(b���U]��YBusڍ�͓�4��]�ml�H8:5�ޑ�69*�b;�����t�pn�,Y�ڐ�&����vA��Ʀ�)+��t�⎎��KT�
�c-���9�8�h�s�����q�\�d�b9�p�6�c��4%���35�l�l$�T�����A��d�	m�B�p)iI��`��N�J�+��*����$�I{�mc����bA焠&	�����k�+u�e�ִ�o.�%�z�x2�;mP�;�*N���@���l��$�\���ňB*Ս�ʪ��l��$�\�����!ljSvQ|t7M�ـ|䕀k�V�[�\0i5J,�Yn�ի����5�+ ݭ� �.�IX_Y �ݕwWLuu�n�ǀl��$�\����j��Uj����;�
�1�v�ŲL���=�[�[<6�N������(1��.0dR)"�O�&$�jG�k�W��>a�/��`�n��n�����Y��'�g�]����x�Z�BF��97{����uٹ'�}��滪�T��UZT��v�rJ�&�����p�'jG�N��m�)S�%iۻ��&�� �ˆ;R<�d��X �`�WM՘v\0	ڑ�{%`v�}��y@�9������t*����]�`-ӷ8c�5�[�&�^q�n7R�:� *��m��dx^�Xݸû. �5��f&Ԇ�VI��c�H�d�d�f�0	ڑ�l�� ��쫺�c���_��.|�Y�3�Y��-s��ײ��'��7���ą!��<�t��<=8be�߂t4���������&��ݑ�<J�Þ: ����Ht¡�5�vn�np5��)�6P�e�.!�7��$H��)CA����N�5��&l�M���@�ti�{9�o�K����f�J�>���i%-�1S~z��@���{�h����I�i�|ij���!�k{J@y
cH��!0ü���^ox���Ú۾���9��=כ��~ќ3�_ uC��9d���5wu����,�b`4�l��k1u	��=؆?L��$��[,����4E�tFC3��[���h�0�.�����NaP�>Zh�A���>�� ����tD��4��J��pt�	"���I8���<���DX�ࢆ�E��K�ײV����x,uawIݻ�Wg�vz�`�p�:�e`{�.sx�O}�ת����n�	�UY�vm�?�5������_�����&ֹ�ubÖ��"������8��Gi܊q-�ig�N�[�R���LF��Mr7�$��'� ��}�>�����8���8����`yK0m+J��BT��d���7�#�z�a�{�~0	*y�}���+����(�;)J麳�=��?��L��T��7���JK��V�[n��^a�$o���q6{�<���<|/�g�Jc	V%dY#]8�� S��ύ�A"GOڏЈ�17!d������=�������'����'�p�{�=���K�5��򭌁������n�'N{>Gd�F9s/6܂�n�6ٺ;B9e'4�fύ�yY�zxI�ݱg@K5�$�5�27����v|���ܞ�,ޯy��0�z�g��]����hB�Q�*8l����/R>���I��Ϗ�����$�:��Q�N�ʎ$�����Osf�;T����~<��a�S��UI��9`��`|�=�0	=~<����~���I�߿pܓ��dV18�K�{�?\�4�c�`�H�vF�#)\��cn�K]����F�kd���7�{e��׆}����.��Թ��h�A�[ZA&���C2X�Y�mx�!5��,0�x[�9%�j���r7KB۟Բ�P�������[Փ�����4h�4������t3�In���x����ڶ2Ү6�B6B�a�4���O;!��/^62YaNM���%��f���?:t�^�Yw�Q��&1j^y�A�6욥��;UP�L�4�r�ґ�0/k���k؅�1��:��������x�/ǹ�	�{��;ǳ���K޻�Ui�m�n���8ٲ_�{���s���l�����$a�abMHY-�<�=��vz�y|�{�� �/��A� �$��GM�z��l�d�ݚw��fM6K�S��i�I�ѭ� ��!$q�l�Y�zl�� 7o��D��O���b����D�n�ʡS)�4X<;9-p%�pte{Q[�1���m�7VNh`�w7���-E��p�<�3U�svi����o�]Y'~�|tqЇ������^K��ܓ��{w����TNr}��,��韏�6O^~\�-*�ڽ�Se?+�����l�ş�'���6K������A���� ���>`U�n�[��Vf/���� ��ŀl��7��b�-@n�P$�I��7�fm�$��d>�p�6m� ���$��y]U�5M^Zڱ�-,Ik13g:�v���z�ў�J'����F�e&�bV�6�.����� �e� ٷ�ً �� ��v�;.��ݼ�ˆ�n{���x�U��cE���ـl���#�B���$ �����@�0$��[�"D�`�\ $1�0X0  �K���f��\V��.�n�� ;դ���)]����0>��M���n��`��|����T��g.���0ڑ��}�>}��w�����������۫es���R��g�a��[Jc�9U3�Mf��Uɽֶ�t�r���]��?z�d�`6��9�5Y'}�Z�&�
$�Q8l��\3��?%�vW�_� ��ߞ�ۆ{�@��(���I4���9�l{���Iq���}��
uK:j�S�VS�0=�.9&x�7��`��}7'�BP��"�9��HTt�%T�H&��u�*�>�Y��t�'p���l��H�)ٷ����:�_�wf,��,�ڭ��0Bd�A��x���tw�pی��;M�7(t � Q�.�g����3�3wn�΁��_� �ˆ�����<`�<�V���������6I�b�>�O|�}��|��T')]!�Cz�g��ݚl��ۛ�¸y�4�'=�N��H�Ii5�����d�q茶Y�l���M�����$�*~�~x���Ϙ��cN��n�`y��x�?qq%�����@�r~�~��ŀG��Ou�� 5�++uWL��;�&�T�Z�&�n�/����h.�4`WP����4��+i�3�\\{�9c��Fn�&ҝU�"��jĚz���Ш�s�^-�.sp�,�v��;k��f*:�;g
6\��0SגP�@�ҰLF����G.̵���ԻF��� ����9[�>쑷�S��9ÍKk��^ڣ��p��֛Vww~�O�]��߁�]Ԅ���-l0).�+�pGj 35p1[���麔�է������"e��Ǡ���`K}s��7�ؿ�9��_� ^a�e:j�S�VS�0����{��X�_�?q���d�SfYV��wt����o��_7�� �ˆ�[��'�<�YMD`�)$Q�d�@
Y���_�?q7���N{׋�>֌�B���-F�N{f�$�n��n�ذ�p�q6l��z�Ъ��Ù;7�uU��Y^�vMZۘv3�6Ca�e#��4F `LCB4��K18���ݱghq��{���ˏv�ռ�X<��s5�7��y��6��'�XX@h! �,_��bȎ��=.��|D1v��������?W�<=ě��b�ě=D��"���buI�v�<����n���;$��ϑ=��$��Un��"bM��7�f�O<}�b�=�����	=~0@t{(6�m�&�Rr�p��{��?]�{�����8���_� ����7HG!Q�(rF6�Ye�\٭śX��a^�"Y�֚43�Z�w�v��[橐��]�m�&,{.�\0�����v�Q�!BH�pY'�Ɇ��l�lY$ڞx{&,��:�O;��j���UY��'���7$��u�� �	 ,!�rʥQ�$����,���ŀ{e��>k��d�j����]լ$���IqV�}� ��b�6m��%ǻ=��:�<�G�n��0�&,˜K}3��n�b�7��}���?�u�˸�'`,���H3g�:�7�tnj�^�Ն7�SjO��I&��ȓ0�'T�wk�7}~0�f,��.s�K��{ /h�=Uu�hE�n�ـw�1e�qs������6{ذ�\3�\T$iӰ�Q����O��b�>옰��?.qr�O���$��X۱��F�q�RH,��]���}�nI���r|�0b[Z���`���WW�煒N�/���̢̍���;�p�?qs�/�-\��ut	=�����<���Wٮ�h�h�Z�Gn)Ȃ�ۡ���zɇ��Dp��L���n�|��V{�Ʈ�vr�wUg�n�b�;�1`vLq�٦�=C�Ei�(�BD���o���6{�Xg���ɋ:��^�VL�:dm̹��'���7?7�����s�Ԫ�~�� �/�!��e��]���֍����s�܄��b�;���~\Is�8��*��� _���Uu�hE�l���w�b�?$�����$�����$����Kx��K$�l����%'��ssY�4vK&�pSIt�L��Z��-��>?�d
� �a��}!=�B���!y�uwu�C�qӪW3 �	}+H�����D2�"Z�`��T)�i~�#�E�c�Ga$C�X p��%�"D�#��R2]9�a���j$a$�/<NpH(�H80�!���X�1�d�#J@h��Xձ��J��5��`�D&��B��No��CN$5�nh�۽��
>|K��$P�7�M�G�쓄
BM��7��G'$������c(@�e?`>��ώ����u���rNx��Qm���	2�[UY إfx.k�mь��ڜWY�ѩkB\���K�
�9x���td�Cj��'����r��i[�A��o��}��]"-��22�[8=��/QXria�aPvf$�IM.2��\LB��;9F�����clr�LP*�'e��m<�pcļP�e1�e�]	�&��v�fsq��[��Nmŝ���.����.*S����cnY*1���m�[EZ�s�֘��@���r�s�v�3 ��3Ξ�=���!��.k �f�z��ʼ�w>{qJ�DTf�P^�p��3J�O`��ː3��]Чj����[p6kcio&�΃��n�I9K������f�x��[��B�Rs��	g��9Ƌ�힮��1g�v21��������;$s�Xq�'.�a��a�q�-��<	z%���(LK�ыc��H�N��j�u�nٝZ�-���A���Y�S�XM�	Z;a2�����m-"q5��T�S;R2n�s��ɶ���6�1��-���E�b\�[]��k�r���h�/<E(p� 66K+�42󳶼m�ͱ,�j��o!�y�R���"s9�kFݏRUڠ�z�c�p=�m��'Y�O;)��cO1�3���v��G+��#td������Ѷk���Sq�����3�8C�F��Ȕ��u����b�C3�y��b��eҘ2�bg�%�mh��]����r΂�I|�
\��/[a`j�M�Q���� 2�Z�XV�p��B ��2���)���vL�hS�ҝ�쳉r+`��:��u���v��^���N�m�9��u�����VB�ͺemV$hL|n�@�|5�x�pL�]��K1n2vIa��m�T0���d';[�
BE��饀�fL�ܑ;m��*�(%�6|;�e;1��ipC�#q�ڃ7�K:���;��"�e;��;�����(v��E���f �A��ȅ���՞�f66�꺸�/c���6��I]���z:R�D,Y�̙uhp��i�lC�Oj���8� qPD�PvF('� �xd��;k���g�����\�"��j���:�*��������[q6�+�Mrʖ���+u�Ƹ�����\� �����������'�t�;Erڃc6⇆��c���.7*�Z����1��1!�wI�eһ�)Z�h�`���z��4b:m���{��=*-��n�V��>�㶱n{K����6n��ۖ�
D���Tﮂ!�P��8Iy&�4YiL%�4�2��͊�i���0�YQ(� 1[kn����H�!�p�����!�'�=�Y'�̱�}$��$���_��<�����U���7v��LY/%Į�O�� ���Oq���D��L�f�rGUk ��b�;�p��/�J���~�O߰}@W$h87cE�r��8,����?ힼ���O�=��:��Su^wW�n���%�\S�\������X{.{�J���
ʤ��Vdé&�k,#k��6�z���na3ֵ�+���&��cH��Tq�����{�vb�;�p��.q~\�h��x����,Um�Y��,ִnI���u0�,aB��i", ���H����E�����k�rI����옳�?$�T
A�ߪ�۪t��'��`ݗ��S�R{1`�{ (t$�5UuN��P�ف��$��=Xｋ �ɋ�_��I�����ɣq�$�Dc�5"�O{�b�:�=����7}~0	�#�	6�9tիMes���<����ě�s`�r�\�f��	�b.�ϓ��b>��bVV�L����b�;�p�$��K�^�6�����y{�ݔ��HV����Ş�K�l����;��,d����K���H"�?���V�	�_��&,"��D040� �@��~ٹ'�ߵٹ'����>�m�ֵ7'�W�J����X�~�� �ۆ�$�IW�!�4�;�J��2����������%�ǵ��	�_��&,���nH�����T)fsơ�c\a�4q�1�n�0�B�� ��;��Y����"�n�ӫ_$�,wn�L^K��q�ͱd�4�j{LF�-�M�d����s�K����� ��ذ��y���	�k&ێI��
.Gd�{vŒgdŇ�˜K�[u�<ҧ� oT��b�E!J8,���_UP��Ͼ�Nf~�w$���ٹ?Pb���	J�E
�T� #�AnO~� Q�?;m��wTpV���e� ������\K��߫�I�ذ	�1`��/w�	/.7JdϦ(��2���.-�x9.7��`Q��Z�e,��wH��YLo]T�8+wk�<��`��X옼��޲|�lY�Hz��i��i����I.�g�����*�~��F6����/�m�6d7���	��Nj�B�a���8�~��m�������..%UO��f6��f�s�$��Ue��$#I���Z(3�{��r�o~��7m��=��9m����	��Hi���1"���e)8�Dي�m��~\Isޯڷ[o��^#�����IAB�*b%q2��b(Z3�����N&1��.����c���_CM�m��Pxaas�A�upt�)�t�d�zM�B�b276!%�qi�[��d�í�\$��8��X�r��kƃ�FJ@.q���e�Ö�B!Ʀ1H��c�NMm��]���x��u�	�%*�lΎ���$dĤv�-l,u�mC�H�8ݜg\;+�1ڈH�:&�;I/n�7,g=��:I+vb�V3��t�Ŗ[q�6{b8hrTV��;����M(	��l���t���M�9n�$3REf����$�{&#m��>^K���i��/��ۚ���!!j����Ig�X6�K����m͹oǽ��{��������l��d��H�no8�K=2++@��S}�|�~��m��-�(�]�  �8�� Sosd��Y��q$��,Ih)�noG8�Dz�����Y3Zַm��>��9m��!�P�s�ym_߿�'ϊ���ݼU_�~���[�%�\ݞҼ9ێ�Z�!��N�n�}��ܲ��t
ڡB+���$(�z�^͘�m�������}ۖ�Ē�ݶ��|�����*�܊a��ni$���s����/9�w���ݶ����9�m�ߥ��P�$��B��HII�)��6۞������?�~�J��z��o����$���5j6�1H��rKI}�Rns~\�If�,I%����[@SoٲZI%��FB�
7)��Ē�b1���n���z�m�z�m�����m�~?�ߑ2'&Ժ�f���v��R�Ea-X1$�:evV�P�_Ν,e�}��AӨ��$��<�I%��-$�{=�W9���s޼F6�zH�Awn�ai��$�Y��
���7W8�[�vM�m�Ϸ��:�� S�_��L3��e
����ܗ�����ݗ���K��	qp"�H��P|@*�>��������U�{�o_�����,1�6#��Ϳ%�ī���1�����6�}��}���BG��\�I!�Um����-���Is�xyĒ�P���'I{�5s�%�d�m$���u6��A�a�7:�n��g���ͳ@�3[=t��&z�gG��"ı�s64��v?��W￶�m���?�m��G�..%�So����Ͷfv�l�dp�%5$��K����h�$^ݖ���v��$|��_�T D����FB�
'	)��ĒϾ�m��fC��ʪ%O;��{�<���OK=�2L[��&v��ӥ��{��r�o��u�������[p �)��?�~*�Iy��HA�&�%���mʒ�m�[�-��m�W����>*���շV��Q�j^-�g�i�]X�F1صc���Ԗ��kfЩ1�OBCT˳#����$�����I,�^6��fC���{M�Ꞻ��nzy�UЍ���c��I,�U� (�^��g9m����[���>�Ӝ����Pu�[=��v�6[�v_}�����U�������}���I-�4�I%�<|x��$�"���IX�U	6�c��{=�>������m��r|�d��Lb##��%�v�K����$�Ъz^x6�ݙ��m͹om�8�E"�`��h�����;��M]e�^F[��% ��u�*n�=��Z%�K=i�U��Xvb
���ա(܃4�hۊǁ��`�Y2P�,iN�dq,��f5۔�=��c<c�+�<kj;Obvwc��$A�H��w��Q�0����<*O��C�f�Zp���fV�&}oge���@n�Z�{-�,6PK�L��J�򲀓R�q-�G�2`л:��O��AÄ�0�0��Ԛ��f@����}��p�,ƹcD��i��)G9���c3�N��,�c(�Z����$?��%���ZI.�ׇ�I%���
��]�ޞq$���j1r�HU���}xy�T	"[�e��og���6��\US}���$MLRq$��lV�K����/�
��9�ZI/{w��I"<��J�y�0��Ci- P�����I{ҭ$��{�r���
�������T沓(��G �K�s
��[B��{7��m���f6��l�}�m�WP��:N�Pw�c�A�Fi^������FL��3M��T�sO&��	�s+��Ga���v|����Ɋ���g��%��i�%_��W�=G�_�v�m�������4�t�eHH��R�Eb���h:M4D� 1Z�#q1��A� 	���?
������-���_�ݶ�<���DD�in��LbF����	�����x9�m�������k_}��r�o{�ڶ�It`�ڐ�.A�q$��K���}�/�m����~I.qr�w����$����Q�!�LRB�$�{���$��
� oٲq$��oO8�]�U�����~)�e��X,��mҚ���^���2�"�-��A]V�f&�ut�;�wI��<�A�2�&)z�I{6KI%����$��澗�~<֭����9�m�r����4����W��|���W��ޏ�����r�o�����? ��Z�������d�6�q$�\��I%�e�����o�m)�5/��P�����nCu���zա ��4�VN!��Ii�b�[ W����C�Ԧ���:�'���m�J�#HX�)
A̅-.71�%��ȗZ	m�cc E��<SR��q%0V�e.���se���e�$
Z�����#4�49�6D�ZHC�e���T5�1�� IP�Kl�מ�{
qe��{��ZC��	"���zeL�@�`�T�4�!�h�=`R!G[Ⓜ�mWZ�BlލM@�0�d��B�f�E8��$ �qa*�� �v<#d"\N����
��P�P��`	=PC��������:P^����{�sWv�{����[m=�[>�Җ�lF��|W��Ӻ�}���������m��O��wkc�͇E�����5wccuk ݗ� ��.s����wk�x�LX����qզSb*�ȏh�5�˗X�t�܈nB`�,��k�us���wI#�T"2��NC�O�vŒyט��옿$��k�8��a'���~_��ݔ�Qwj����ԏ ݓ��Ǆ��L7�@���J0F���
)"�$��`�lxy%����<�^��:��(:������\{�<��w�rNy�}w'�q�DR!PR��>X��o�N1U�����x�In߼�O_���<��:�tjy�I���j��X�q�z�ۍI��ʙ�P':��K>wN�=��B��������	��<v\0����./�o��x��i�*�Z���v��p�;+c�;*G�ojG��\l:/x��R�����>ך���y���To<�U�s�4�$�%�#!��Sp����9S�~������7e� �����Q�We�uuj�Uo ��#�?q~\��}��W�<��x�%<x ��x�l�̻4V�.-nOs<����i��.ݶ6�C����k SY�u\�`-a����T�Wg&T���MN���{�	��	m��̷	)af�R���ݐ� ţFv;Q�����{_0�%x(�3R���9�����ޢNK��8t�Em'f�Z�`��D�j�̫-��:�\�� z��®w6��ujƌ�[��q�.���h��r�u��N��l�1�l��8|l01�<;��:xDf^�x{\S�
l���E��v�g�,���s�}����_vV�R<�ԏ �]�Q��W-՘{[o9��TOU������. �E��Q8�j�wo ��ԏ�M���n��`65��UE��
����ԏ ݗ��<��y����=����
���$���;+c�;*G�ojG�=�>��>���ZPHݭu�N�F�v�T
vq==�{;Y���;K��Y�;�Nz5��Ln��;+c�;*G�ojG�nˆ Hީv˲�V:�uo �lξ�J0���Ar_����w��f�6V oTD���WT�P��ڑ���u�e`�#�"}{-�b���U��x9._vV�u��n��w@�����V`rGXeH���x옰}�P��-��ƛN��Π|����F:	�l����ѭ-L��&���u�:9�a�m��dx�R<vLX\�� ٧,��
V��WWo ��#�7dŀu�B�ʑ�6MZ�Lv���M7T;��o�}�rO>ϯٹ����"�߽���v�� |B9E+v�]��������vT� �ԏ ݗ ��R�we2��V����;*G�wjG�nˆ�-ǀM�R��Z�wm�eq�^۱+Y��H�,�l��B\u���K�z���c�2�18dp2���=��VI��a�Od.\���_��
��E�]�]]]��7e� �R�vT� ݩֻ�'J	�2�W-լ�K��R<v�x옰j�[|�q�V����;*G�nԏ ݓ��s��R�l��	�t�v��WUo ݩ��إ� 쭏 >��o����f]��aAeH;��̤y�����:8���8냶�W��qF���-ǀvV��Ϙl�y���u�"������=̘��U f����S� �ɋ=ĸ�*����ߊ�H�@��N|��d�y��}�1`Ir� oT	j��v]ժ]�s��\��&�ذ	�\0s�I#���d�^���!
T0����=��:K��e� ݭ� �8���H\U�Pa
��E�"�~\��a��;L�Z5.]\	��
�kq1��`5�=]���q'�m����c�y9���O6�;]vN(gn�z�& �u�"\��a(�9�9��r�zt�MV���b3$�+�lF����̙�X;W�p��W�暴mf�S�b��-n�m%�nƳ���Q]�=S��a0@3L����m��S�Wv�0º��j�M��V;�N��>H��ӧI��]>�Q1M����@L[m��C�e�w�]G0�X����)g��Y�KU�uk�w�/��>�`�����X �t��(�v�j�*��>�g�I�J�x��,t��($ssP�Q��P&���sj�;ݘ�	�\0�.�Clw|���[��{��,�S�Xݗ�qs�%�r�g�<�_���V�]����;.[�>�`mlx{��~r�aRI'�Ed�"���'�K��-�Nmb�f픹�ָ��mPv�������6�Ue���ށ=����ǀw�1~U �]d��~��'p|�G#��#�5sZ��s��� O�Q����}��7�=�`wf,���C���_,Wn��ݞŀN��x~�}��Xv��֦��('e%er�Z�������ݞŀw���{��=���m�^�ʦ�����>��Xݭ� ��1`�_������A�e"k��Ё��2�]v�Γene��h٘�bhhm�Ȟt��7l�ݲ�����n���>��XҶU`wf,j���n�X��V������X�ً �����9�wm��cuk �͎����Ic	A((|�Pw�������زI�K�j@`p��H+ �dŀ}���ݘ��v*��.ʻ�uj��P;��}�����X�lu�}��D�P�uc�Օw�Ɨ��n6�љKY��jqӦ�'&�f8k;�t+Aj�E��v���ݘ��k��}�1`�lxv���CVp�]Z�>��<�ً ��ǀ}�1`��[iT�j���]Y�}6b�7���ݘ��ۆ�G�N�,)SN���7���ݘ�����qr�q'UR�A����ܓ��;75l�Ԕ1���ݘ�s��W<���ŀokc�޹T���U�E+V���mt�h�V�\���u�fm�N�PĆ�yы��-[�Ln�`E[�.��<vLX �n�U�.�UՊ�ݼ�\0�lx옰�l��qs�I��'\G��)8l��<�d�{�k �͎��\0�V� �m�՜�uv���X�lu�}��}������P�YÕuk �͎��\0�[�ً �r���@qW�)e�J��h��E1$VA$� ��`�c(oi�C7uy�Hh�x�dx�f�0#1 fp(nf�6d!tIu���g�������A�!ș	M�#0�
�D��f�!7��D��B1HB�F��LE���I !D�0- @	&�H��U���$��v��Y�� 1�D&Ґ�%4���I��8V,X�-M�����q$X�0!4+B,3a�P�M,P�"����u�J�3͞��thg����F��0� H@#��&jHBB7#0��p��sw�Ɣ�*��O.�!�=�����$&6ܩ �I IC�������+,�<F�6����4\WN
C+�F�����z�K;���ꕂ4*��Yv�p�����B֬��2d�dl��������*�Mq6\��w�Mt�hJ�-1jŗG�n@|��mGWv�3�pY�e����nI��r-cpv.�v�f75e�l�DnAM���dؙ�0뮝��7�f{2�Ke�(!.%l��[bۚ�}��:��kPK`�����������`��ܼ���a89�[9�:u�%��¶����Ƞl��YX�f�躌�u�2	Y���k��Z�ͺ�ѥ�Yoh�5�.n�a)�u���Y �j����t�8r;�6^ز��f�V�s�����|Խ���ScA���5�S����J�ш]��,I]T�AsqE΍���@x�e�n��϶w��V��\m���E�v����
��jԞls��%�CQ\�\6a+�]�bjLm!;zi����N�2�i��F
�K�s)�����ZǊK�V��1sf0�����2��ƥ��'�ޛgۇF�
K��֤���� 
�r^�W��}0�7i��2^v萘"���;n#�ci��ur=C��'��;��y�sΖ�l�\�Z�pۀ$e�h�í�7e�󜼞ݵ�*k+yF�$l�X.؉P���Ƹ*��p�b�N��M�M�G��[n��V�i�I�-��iT��n�hjB�)m�N&t�͙�i�6��l�'l���`�:@W� -�juH�Nnmc��%�#(  �Ng!�rcJ�qY��dyznbJ۵�!��`��a��2둋h4��c���u��[9�I�lm���I��v-��pvQ�khqNz �qK�,r^	�!����[Q�D�4dM+K��� y�Á^ܽs)�l���@��v��<��mۖ�����)�p��a7Hv����+ƹ�I�K�YotEƗ�%��K+q��ں,K���5�Q狶�l���vǡ�C �Y��Hk3-˫|�ih��Ƒ4 =�4�x���xiO�O� ҵ�|�z�� �~Ϳc���.�S���+�$놙NdmY�Y�]d�]�hؘ���#Q-�)�+2t1���<�AۈVݤ ��(�R^���3v�%��
����R�O�N[1�,9	F.�ᣯIMM pԇ]��0���4kDذ��#�e��e{U�xìl�{����!na÷�5��a�R����
�� �iIRW]�+3���0��t�W$G����'`5�␱�%H��)����f�H�[]�8[��9붠6 �����$��W���~���}���ݘ��ľa���X���I�he*i�ݘݭ� �ً ��%`Ip�%�s���x���T1���Ob�>��� �K��kc�>3��>��MsQn�����|�o�~0�O<vLX �2��ګ�*��UwO ���ǀnɋ ���G�?��,�l�y=�4*ްuv?}�����Z�#���!�]��m'm�gb�;"]/;M�6��]Z����;�<��1`v���8����d�^$�"Q(�\�̞���78�@_x���9��#�6m� ����v���1� �ݬ�ԃ�;%���v��'�� ��A)utS�e�[x�ʸ`v�<vLXO���x���&��V���wv`v�<���'���;��7�vK�P��:uuM_.��k@֑+�	�fn�
q�;S��9���s�6w]��-P�T:��nɋ �l�0�p��������^��k��?�իWE�7V��\o?.q.&�����S� �ٖ/�	�V�R)$*�tc�Y'��]��s���U8�T��IƦf��=ǺU�s�I��H�p8�m�U��8�.y�{ذ���.�R0T�6�e���x옰%�������v�<wf6][T����&��ҝ���e�낹x�PHl[����g.���4�$\��O ��xv\0�l~�>a��ŀ
-Q�/]��&ª��;���K���<���,��l���a�U@ӫ�0��<�&,<���\��`=~0	h�e���uo��{=��=��`5 IQ4�!! B6��%J[R�!%*R$���,d��%�Hĥ�d$��d,a�~DM��~�>�~|�?Ǩ��؆�u�x�����p�>�lxvLX�	G1�'�Y�2�/H=rkVN�;9{n�l��E�by2(�.�\*YR' ��t�p�����>�lxvLXݩ�oT	UYe��.��۪� ���縛6{ذ�yy��p�&����lv۲��U��;�b�>�W<�{=~0ڞx�O@N_2� T���b�`�p�;���<�{�, Qj�	z��I6]*� �ˆ��ǀwvb�>�<���;�����������5��K�m[��Nֆ2n��ۖԓ�*s�s���n���������eP��L�Zb9���XkY�M΄�)�j���o3��Q�.�2n��j��W��q�5�aii�i]B�X��ڱ�U{4��^B�K5�m���]�l6�����͆��ىKb�^S[��!�۴.��t�ĻH������,���FXo�;��;����y�����k�ؘm�v��� [��׭��h].'r�wd�x���c���@����;�1`wU��0����=���e�v��:��wvb�>��o �e� �kc�$��ּy�*����N�U��/��mH��8�^�`wvb��t:��N�����ۑ�ڞ��a�{ݗ�����U�[���m�V���<���v�x�R< �R�ӵJ�;T�RR�X��@�u���Xf���<�`q�6k�$bm�v�Wo ��ŀ}ݸ��ԏ��7jy����b�`�����g�z@x,_N 9�<����rNy�����Y��%��@�(���ݗi6��[�7����>�lxwf,{[R��<8�v�Z��U��>�lxwf,{[R���x�ւc�|c�N��ݘ�	��L�e|e{� �����Ǳ��6�qYj��ai��z5���Eƞc�cca�lTД�W�60+s)����okjV��ǀ}����e�$�bY��ۆH$q�TqY'�~�`w��������_s��u�q~�Q�3�����`�%"�O����<��ş��"@c$H��!@d�*DB FDb0�@��īR6��"A���$,+ba25�	��k��v�C��d��~��J2�J9%Ȭ�����`�u�}�#�����<iN �vt��*���N��x�����wjy�ݘ��\�-�w@YT�Ӳ��j�֞�>��5G\N�j�ͣE�2�ҕ�Ō�"����Cm�]`mH���<����|��R�X���	��r��4�]���ǀwvb�'kjV��+=ě=�0^2���|T:��l�ŀN�Ԭ�V��ǀ|�qU��탪���{����^�_�� �keܛA�1"��I�ȁ!꯮
�_~�$���}�f���������>{%`��$��~}{���'e�x�D�vZ�tZ��UO�7g�X"�����n{���:.)�V�ݎcnCp@���O|���'��K$�rdZ"z�u�'|vi�r�r��x��x�̳ �앀}����O��KO����\pD��g�?���Y�}�#�>�lxwn �ujb/�@
J9��(ܛ��=��VI����8���g����X&����4���kc�=������t�߲����]�"�� �� P�D`�@H�"1��	 �H��hd�R�UJϦH�vf��5nh�Y,��C%%v{d�,,E[�::�����Y�{N���5!�q�T�΃�s�4Μ�hn3�ys�Y ǅ��pBY���wHY�ڏ6O(]>N����4XMpB"�A&��W�I�u�˞=���D��F�F�/nےۘ����Q��x��v&Ulɰ8�ؙL9�CH9i��uux��N���D�ۖ�&�A*�䩿�$��	$��|�na��s%��Uip��K�����45�8��v���6�V�%|T:��'e��6m�x�R?�\��~��|��C��7&��U��fܧ�}�#�>���ݸg��l<y���q�R5d���VI�?b���͓<|��Q�uHܪ�Wh���V�uo �Vǀwv�lٔ`~Iq�&�Nn�D�C��LqY'��� ٳ(�>ڑ�J�����Z�:��{r��9�	��,���������"&s>t��qm=�k�)��߫l��Q�}�#�>�p�;�p����A<rH�ۑ�$��1_h �@
4 �A	�(���g�W�� �/��fQ���6O{�,j��2�'UV�����ۆ����Q�vT��6-MAb��v��� ݩ�fQ�vT� >�/ �	Wt؝������fQ�~�9������}=x�lx�\Oэ��;]����]*�Yb<�s�"���L���su�˻2���66��4�Z��߿�o���� ;���7kc�6l�0[�UX�;�J�V���͒T��'����R<E�g�Wbwe[uw�n�ǀlٔa���14�X�ÔL���K.���Cl����&�3n���
�M&�A��j蕸���JJ��- �Wtٱp6@*�o.��R�Y	%ѥ� WA���-0$fLp#DIe�$dRf�de'$a	�Ԓ!Yr�4�F�l(B���9t��(T
S5%$�XɆ��)Li��oL]0M�.�[ؘ:U��K�Ja�!(@*L-�Y[ZV�JY�M��l@�-7�6�Tɘ�@$d	�a0c��ޘ��.;�jXT�-�YB�'3&kF�3�;s ��T B�j�� ���r�6�n�F�+n�� �H��#8I#ы�I��L�F�a]2�E*�l��2�	Xq��������S��C���#�TP
�<O�L:��C{_M>�)�"
����9Ë�ڬ���K�;ݷ@TnЭ�ʺ�x\�s��Q�u�z����lx �n���U�ڡ����>se`�e�����2�Y�"�r�� @�a��Ǝ��r�l[�.��x:h��x%R���#��Il%n�����`����2� �l�b��+m;��)�����<��l���0��� ��^��;��v�c��0͏ }6^ }�/ ��� !�a�9.H[�EI��c�I�s%�ov��$�S��u#��\������#;�q���IfD���'�̖I�_�X�,�[�%9�z��Sh�n����ew@;^�/hK���ٮ�E��ڷh
�N$5!r�.&��'<�U�{�ǋ �VǀvK�;��@8ݡ[-3�uv�͙F�+ >엀okcͪ)"G�bH���%"SnFl�չ��}ڑ����͙F6F��Iڱ��T��<�[�V6��ٳ(��o���yDׅ��][UUU[�7����, �l��ԏ ��T�2,����	$�p�X�,	 `@��� ń �A ��k�t%m�rÆ�gs:�Q ѵm�׋��q�۩C��wG%۰=!���e�*�XA,��p��-���x/5Iێ�S6*�5�ݓfIZ���mgxy6�lƔ�=,�ST���� �FA� 6�B]�`]�K�Q���%wbVn����fv������=��0Y��،�nd���솅��B@����r�ma�fΐ��5t�f�U�����c�绻�Βn���������:����/N�F+'��q�,��m�-n��(�NUݵrV&�Wv���ŀM��}ڑ�����VI:qn����$�8dQE�M��|�%y$��&���7�� j���U�N��ݦ�� ��J�7����&��� w�׀H��m�*��ӷn���lxfǋ >�/ ��J�;ݷ@Tn�-[����vlx����d�{[�h��n�C��]���gu�nz�q�\v+����k��g��0�1����F:�i��~����V����K�K�0�CذOy�ST��L�k[�y|��߈����'���K��s��;	� >�/ آp�+m]����Uu�okc�;+eV�����|�%`8p�]lwM��Wv�<�Ǿ�� 璘 ��#�7���5��շV�������R<{[�[*��xRF��#�Յ�Mm_���`�һ�����\
oK�ٽ4�I��� �16�	8�n@������_vV�[*���E���b�i�.�����;+eV��ԏ �m�H�݁l�%N�� �r�}���s�%}�\�}��� .�ڪ�5]$Ӻt�}����xelx����=U�z{�`�q�Z>WXϲV�Ķ�=_���_d�_P�
�7WT�t�]���!,��+4l.a��k7 �dXp��re$q���j�Wj�
�uWX_d���U`}��0��J�#��ꝃ�l�ݻ��;+eV��+ ��J�;ڑ��װ�$�2��'����<��VC���[*��FF�M���U�WXݩ�ԏ 쭕X�7�z�	Z�H��D$Fz��E��I��Da 0B\\����N����S���:�U�.�v�t][�;�p�;+eV���d�u�+$�B���Ĥ�H�i��ɂ^^{I˗��`��!YNzQ��D��ۊ{����T�i�8����������J�>�H����un�U	�Ut�'t��}���d���<��Uf�AX�&����d� �v����X}���T��[j����V��e`��� ��V'�nG�p�*�n��M���`��� �d��ԏ &�x\\Jul��|�Xݩ��Y�j�F���Xk)h�W/X���h�[��hl"��W��:۳f�Ɲ7b}E��n��Wgn��	�f�F(ݤ2�u��a�9�m�p���sm��,ML�e:Q�7e�WC������V:L,quvX��8�������n� ��-v��Kc�h�.�ҙv^N�6���fPV�YsG`�����wO�}n�_ZB��Ǯz�nB&�!�h�����\n-��M�:��x:mƒ�D��% 2�����<���/ 쭕X�*�M���U�S�xݩ M����U�M� H��B��U�-�t]��	�^�[*��J�>�H��k�m]��F���d�
��m�d�[�vI�\� &�x ���U�R��*N���`앀}ڑ��/ 쭕XS��m�����`��"��P	���A��qkR��\�.����Ԃ�b!��u�>�H�l��vVʬmH��T��[j��UUU�=���ė"�9���s���U`kc�>}��E��v�uMڢ��� 쭕Xڑ��%a��n�$���I�$��%)�˪����=+�x^�ՀG�V�[*�����4m�kv������� �d���U`jG���8��T�r('d8����vA�u��"�3v��1Y��{Z[Vl�ЗTئ]n�_ ������&ˆ�앀}�c�.ج�Zb,���;�q�v\0�d�=�Yi�]]�U��i�Ӻ�>�߶nI��߳rя�>`��28E|�X��C[@:S~e��0	ڏՀ}�)�
���uo �ݕ�G�+ �Tr�	ڑ��T��X˻EU:�� �v^���`v�x^���l��):T_
l�å��g����v�Is�ݍ�Ǡ�hӎ��n�.�[�b2�-��!��$�,vI�^b�O^���׀u����ݻ�t�Ӧ���R<��s�.��9�eٮ}���z쓋��^�
H�ը$�
HԎ8ӷ�k�Հ������W� �׼���B�)]ӱ;�uwX��>��[�sϵ�ܘ��*�)�� ��5����9�m�	�	�A�,������R<��ǀݗ�jIv��YvE-��5���fU�ICF��<uD���cuٺ�0��BA��Cs�s�wLz�0����R<��ǀݗk�K��W� �����)�Gʪ� ����we���/ �e�<�=�'㘬e��S�x�z�}ڗ�}��}�����X�M�J2rId�.��O<�<��ǁ�s����5�?~-۴�un�7Uw�~�y�v�� wv^��s�nH�� �0#9K���ZCG��p��] m�����v{�R]� B@�0����J%.�{�WM�ѫ�ӣ$� `H`�b� ���"21"@H�@ӡ���"��#J���r`���R�
�E"�0���a5��hu�&�:���#$�$��$ֵ�e#D� ��$abi1�&�3F�1�ĖU� %)cD��U�0�D����x�6��ׅd��t�B`&��Қ��9@�;�@b�H�e(*�)�!�!J��M�R�c��@5��A$#-�a,)(M.�(F�B!P��l�4�e6p�h�i.�A%���bMJ�9h���Dvʱ�	�E )m+��� Q�%IR�`r�5�C�!�3N�Q�!�� B,R(D��`�"�!!B��T8E����	
Zĥ�-���JA!KI	����6�h� �-���8�PHH��$�A+��W`+���Q�U*Сd����Ʈf�F�����,��b1#-�`j=# Q@�nͶ^e6��m,�i�:�3H����x�h�i�8�ڎ�ؽYN�'Qɺ��6�0ϝ��p��S�y��;���8���jv̢���=�y�S���lg��+��M�⎄�s�*8�Mח��c;Hs�\��i%�殏kq�qA�컆˧��m�!��7`����S��K%��u#g(��=����M��5]QԢ��-�0�v�v3���6�6��R�: &���(1�آ�˝���2�����ҳ!��:�6���U�m�y��u��A�8�0�+�\��N�޺�
7F�6ܷ-���t��r�ts�dЙ��ئ���%m�Dѝm�#d�몴z爣mȪ`�Pr�BUs.E&,.�F�n�m��;;�p�@Xn�Ү%Ŷ�N�d0��vfK���+M�ԛ]��l��ve�n�׳���m{;�� q�S����ڪ�a�/nW�-��t9ۆ�T�)ۮ'��p7A�ۓLne��v�ٻy�c�f9����+HC�&���f֭�����kB+eV�^c�5�#��m�x;h8������[+�#k.q#L.�;G����V�h�n
mn���f�-�6���$ ����T=��r����]�њ<��ዪ�M
��"�2�9�B����)��q-6�Z)�$���n(UT��&u:;D�R��*�K�r�#id�3  ��c�6{�l�gvI2i̍�[m7lMu'n���ѵ��t�,l�k �f��B������I���f��Ov�6�""b�);6��;���Ryn��yLi�cl��(�[E4X�X�=�l[%t�BWwI�!:� =&�EX�]y��N���Ρ��-�4
<-Z7'G\+S��N��+�F���S1m�R��]g����ٓ�0��m�V��D6be��܉Fbq�cQ8ҡC �. ;X~��W@�9����M��}�O�"D"-QKET������ >���P�Ф��h�5t����CiD� ��y]�۞�،�
��mjŅ��:�Q��-�M��he��0I�%�`��re�s=�ۉ֫6&�@�m]rV��v�z�G 1�1��Z�K���J�d"h�\X�1,��+e&�ݰc�Cd����B�I��
�>5�S�cˣ����;%�Z����/U�Q�,��`1�іRYf�WM����s5�m���wt�wK�G�|��ggGAZԉ��u��4��7'k#�vzt��1;�Râ�v6;.��k�wn��	������}ڗ�ݠ�W�+$�|5?�.$j[JH��{�d�5�j^�ԏ ����l�t���ճ��Wx��K�>ڑ�v�< �� S�ORt�[�c���>ڑ�v�< ��I�wj^;%<8��wT��)ռ��ǀ~\\�{'��#�^�\��$�+ʊ�M�[z�/��;p��`۝.[t��í��GT�Z	
��`�k����? =������ڗ�k�V�kc�>pQ�V�]&���5�krOo���ڀ��t��_a����O< �%�=Rrݲ����T���#�>�lx�K�>��o��>'�_XZd�8�n|��lx�K�5�j^�IX�Z� �bF������'ٙ,��B���G�z��[ i��*�C�EN��׮{F��'�tP=�v	H]Ml:��WRp�.
Z
�mj��S��_v]�䕀w���.%���� ��Ī�U�X6:��9%`�lx$��k�˼H�Ô6SwGT����< �&��C�� ��[�|ַ$��`V���˫�ER�V�=�%�đ�q!#��US���#��^�X{[�R�Ul�ݱ;wwx���5앀~ݹ�_L�g8��޼����t}������ݨf�1�l��䕄L�AG%�0��A��,���,�ZAf�#J2cMH[NIt8h#A�Ǜ���Kı=�_v�9ı,K�{�m9ı,O�߻�m9ı,O2{����]���F��O�D��߻�ݧ!��L�b_�~���"X�%�������"X�%��}��ӑ6�e:'G����B��j�ʮ��â%�b_��u��Kı>�~�K��ș��߳iȖ%�b}������:'O���X��4HŻx��bX�'���ֶ��bX�'��{�ND�,K�u�nӑ,K��dM���[ND�,K����ۚ�P�˚ֶ��bX�'��{�ND�,K�u�nӑ,Kľ���ӑ,K��=���ӑ,K����Z�[b��!(%�\������e6֗Ƥ�V�%U��N^I-�IO#O����,K�u�nӑ,Kľ���ӑ,K��=���ӑ,K��>�siȖ%�bw���5K5�i3����Kı/��u��Kı>�~�Kı>�]��r%�bX����v�����t!��m|dN3M��M�"X�%�������"X�%��{�߮�Ȗ>C"dO��]�"X�%�Y��K��A�F�^�p	1��7.kZ�r%�bX�}���9ı,O}�ݻND�,K���[ND�,�@�Cfo�]�F�4<�}�E7#SS5sZ�nj�9ı,O}�ݻND�,K���[ND�,K����[ND�,K��{�ND�,K�>�a�2O��kdSe`.3�%z�mWMvm��^-A�����8��Z:2���M���bmk���!Ō�>W��;�[s�hl66�GF١�e��@��4�x��f��ɍ���b��A�u ��.;c�윚��i�J; ��Hdu��7X����oh,ػ��Vn��l�Gl�;d��@GH���R��"�UKT��1I�\jZ�b�3k�E��gz��g�	���KX��ű���h�yCby�s�#��ł�k�S6]K���~t�:'D�_���[ND�,K����[ND�,K��{�ND�,K�u�nӑ,K���vL���SAink[ND�,K����[ND�,K��{�ND�,K�u�nӑ,KĽ���ӑ,Kħ_K���al�ֵ��Kı;�w���Kı=�_v�9ı,K߻�m9ı,O�߻�m9ı,N����l�e�em2浛ND�,K�u�nӑ,KĽ���ӑ,K��=���ӑ,K����fӑ,K����^KK5�i3����Kı/~�u��Kı>�~�Kı;�wٴ�Kı=�_v�9ı,Oࢡ�����!l�!4ji��j�S���������v��+2n���F����NUݢ�*�d��r�Mh#A�~��p�bX�'�w}�ND�,K�u�nӑ,Kľ���ӑ,KľO��֭NcNB�rK��A�F��oM��8�!! V##�"!����D�%��k�ݧ"X�%�{�{��"X�%��{�u��âtN����~+m�v)���8�Kı=�_v�9ı,K���bX�'���ֶ��bX�'���7C��4��h��0�LE�L�m9ı,K���bX�'���ֶ��bX�'�w}�ND�,K�u�nӑ,K���v&\�a���[��ӑ,K��=���ӑ,K����iȖ%�b{���r%�bX�����r%�bX�w���.���k�L�86�z��e$����#��\=G��qA�v��7Z}��y��Q��Gm�t�:'D�=���ǉȖ%�b{���r%�bX�����r%�bX�g�wZ�r%�bX�}����)\��-�t�tN��:}����9ı,K�{�m9ı,O�߻�m9ı,O��{v��bX�'~����bĻ(+s�O�D������ӑ,K��=���ӑ,`�+���Q��O"f����r%�bX�w]�v��bX�'��N�2&�(��Q9%�᠍h#C}��iȖ%�b{��۴�Kı<�_v�9ı,K���bX�%�t�pd���\�n�âtN�������Kİ�G�w�n�Ȗ%�b_;��iȖ%�bw߻��r%�bX�}�W���o����Y��\C��wb��qz%�N%���%�Cl��.�[9[#f�:�O"X�%������Kı/{��iȖ%�bt���iȖ%�bw��A�F�rz f6c��kWiȖ%�b^���Ӑ�F�$N���&��	���6��H�y��M��btN���'��!��v�âqbX�=���r%�bX������Kı;���r%�bX���u��Kı<����orj��浴�Kı;��siȖ%�bw�}۴�Kı/{��iȖ%��$TBx�q4o���ND�,K���y-�td0�\ֳiȖ%�bw�}۴�Kı/{��iȖ%�btϾ�m9ı,N�{��r%�bX����s�j\ˈiV��
b�IstMu��X[����8q�W�8A�JL��5�,�q��������bX�%�{�m9ı,N���ͧ"X�%���{��șı?}�߯�>�tN�o���?�Z�#b;m���Kı:g�w6��bX�'s��m9ı,N����9ı,K��e�᠍h#A��))�̄!���Kı;��siȖ%�bw�w�iȖ%�b^���ӑ,K��}��p�F�4��s4���)��YY��r%�bX��]��r%�bX���u��Kı:g�w6��bX$�Cd�wC��4����`f6T�C��ֵv��bX�%�{�m9ı,N���ͧ"X�%���{�ND�,K�뽻ND�,K���-�\��w�]X�.Yd��p]�GC�vL
�2�;i�YE�W��v�9x[r��&n8ݠK��nY��3
K�L`�[5�Js5��ikş���y��k�u� S@n%XAmH�V��c6�:�صK�qO3]g�5��SB��u�F���b�M#��i����g���k@�9�.Lq�vw.���f	��x��mh���������:v|�o����0vk�)Pt�aa�m��H���JWA�c�dD�̶�e��`�ݼ���ı,O�fӑ,K��w�ͧ"X�%��u�݇�Q'�2%�b_߿~�ӑ,K����ɗ�MMBZL�fӑ,K��w�ͧ"X�%��u�ݧ"X�%�{�{��"X�%��>����O�&TȖ'����#�\�FL��sZͧ"X�%���~�v��bX�%���c� �Dȟ��fӑ,K�����6��bX�'���r��̚�R2���r%�g��ș���r%�bX�3߻�ND�,K��{�ND�,K���ݧ"X�%��vw�Dԅ$�*G$�4��hhy��9ı,N���m9ı,N����9ı,K߻�m9ı,K����i9�,܍��ͣS�W�7$��d�W��Kd욚wY�3xF��K?x�Kı;�w���Kı;�۴�Kı/~�u��Kı;�}�k}>�tN�����[n+���5�ND�,K�u�ݧ!�*�< �Qb���C8M#�T��ȞD�.}��iȖ%�by�w;��"X�%�߻�ͧ"X�%��ڟw&�IRDȍ"�4��h-��t8Rı,O�����r%����;��iȖ%�by���r%�bX�����kQ�CVR\ֶ��bY�`dN�����r%�bX���߮ӑ,K���}۴�Kı/~�u��Kı<���ؔ?&1[u�âtN�����ͧ"X�%����iȖ%�b_{��iȖ%�b}���ӑ,K��}��>Z�\%��
d.��mGDh���mۙo<k��1ƃ]�Jǯ�tBu�����nkY��Kı<�_v�9ı,Os��m9ı,O����l=�DȖ%��k�ͧ"X�%�߾�w)����d��.j�9ı,Os��m9ı,O����m9ı,O���6��bX�'���ݧ"X�%�{	>�髫�K3%�kZ�m9ı,O����m9ı,O���6��c��_���U-� !	�!��F��ctaF8�d�)A�榐��d#!	$�8岆�L6[�^ZG��d�,�� ��q����!��30�!{@�!P�eHP����U+b@�
�%���BI�i5E��1��	��8�d��ѢG�y��B�Ὄ!5�;�#��0�����
�28x)*8�`D�7p9�7��䞂��*h��͐' ����	�!I$�ɨ�B�0���T�w�2��uw<U���N���~G�6�P)�D�PL4�*��	뭢�=EM/�老W�x�O��� ����o\��9ı,OsﻛND�,K���j!�\B	
9�᠍h#Cn�ӑ,K���}۴�Kı/��u��Kı>�_wY��Kı<���d���4��h{�;v��bX�%���bX�'����6��bX�'��{�ND�,K������Ge���(U�[p`e��5�-��cѦ"F��+�u�nS�ԅ�Z��r%�bX�����r%�bX�{����r%�bX�g��m9ı,O}�ݻND�,K��=9�j9�&�
[��ӑ,K���}�fӐ��"dK��߳iȖ%�b}����9ı,K�{�m9HeL�by�Y~&S��Z���ֳiȖ%�b}�۴�Kı=�_v�9ı,Os��m9ı,O����m9ı,O����SF�����jm9ı,O}�ݻND�,K����ӑ,K���}�fӑ,KkR"H�  �T��I�?ׄ4�!��}������Kı?}���7e2�V�Ο��:'G�~�b~r�C�����i�Kı=����ND�,K�u�nӑ,K:{=���Tm&��Vk�0qz�h�B�y��^{v�ec@f�2��moP�.�-.�u�m9ı,O����m9ı,O;��6��bX�~������%�bX��w����bX�%{߳��5�5MԤ�kY��Kı<����r�6�MD�>�]�v��bX�%�~���"X�%�����ͧ"~U��,N��ͧ�3	6�4��hg����Kı/���m9ı,O����m9ı,O;��6��bX�'�e�3!i� �"�4��h_����r%�bX�{����r%�bX�w��m9ı,O}�{v��bX�#=�A���`��4��h}���iȖ%�by߷ٴ�Kı=�]��r%�bX�{��6��bX�"U
�>�����0����4Z�n��LC��jra]̸Sa����l�?9�m��G���&�,�d:��!&c���<�S�ͮ���1��0�����D�-�v�B:���7\��`֚��·�dx*X�C,�PN���X�Ʉsi�qǟe=kp��M��7`�7f�v�n��ȷ�X����<t5vs�^���,z�t�nl�m���� ���-p8��h��a��x�lY�v@��tnS�t��n�sb-�����ɩi�R[n���v%�bX��7ٴ�Kı=�]��r%�bX�{��6��bX�'�k��6��bX�'�}{l�I� �k��O�D��߻���9F9"X�����r%�bX�}����r%�bX�{���9ı,N���k7CjWgΟ��:'O�o�iȖ%�b}���iȖ%�by����r%�bX�����9ı,K�߿[�.�%h�7cΟ��:'O~���m9ı,O=�ݻND�,K�u�ݧ"X�%���o�iȖ%�b-#V���FE���p�F�4�ϵ�ݧ"X�%���nӑ,K���ٴ�Kı>�_gsiȖ%�gG߰���1��&���[!@׬�����c����ݲ����Od�4��t��\i�ܹ���Kı<�]��r%�bX�}��v��bX�'�k��l=�/�5ı>�˴�Kı<��ΓYu��˧Rə���Kı>�_v�9,A�E<
 t(�&�X�s���ND�,K�u�ݧ"X�%�����O�D���}?C�&�"Wk��Kı<���ݧ"X�%��u�ݧ"X�dL������Kı;�w��r%�bX��З���.kAn�2��9ı,N�~�m9ı,O=�ݻND�,K��ݻND�,KϾ���r%�bX�����6J��%�fkWiȖ%�b{���r%�bX����r%�bX�w��.ӑ,K��w��ӑ,K��;%�}s���$�e�P㝎���xx�S��c��ɞ	26��<�a���Ƶ+��O�D���_v�9ı,O��}��r%�bX����ișı=�]��r%�N������f��Z��\����:1,O��}��r�9"X��k��ӑ,K���~�v��bX�'{��6���A��,K���Ƥ�՚ֲkR��Z�ND�,K��w��r%�bX�����9Ɵ�EaFCB���BH��$I�������" B@�+$���� �~a�������iȖ%�by߷�WiȖ%�b{��2\�[�k4\�5v��bY���>��]�"X�%���w�m9ı,O��}��r%�bX�g�w6��bX�'�5��2�R�@��᠍h#C���iȖ%�bw��]�"X�%�|���iȖ%�b{�����Kı)�~t���f�&.R<˦"��hW�(y�79bx7U�*����e4�%;�:�Ѭ�y׵5��ND�,K߾�uv��bX�%�߻��"X�%��w��ӑ,K��߷ٴ�Kı)������sZ
[u���r%�bX��~��#�2%��~���r%�bX�����ND�,K߾�uv���Pr�D�?~��9����a5sZ�r%�bX�g��ͧ"X�%��o�iȖ%�b{���ӑ,Kľ{�u��Kı>�gI�SFZ&��I5�ͧ"X�~D dO~�?M�"X�%��{��v��bX�%�߻��"X�D�,DI � �X,� '��.�A�D����ND�,K�G�]8d��mHn�h#A̷�ӑ,K���}۴�Kı<���r%�bX�w��m9ı,K綠�������OM%�ˆ	�r�:�q:��Lej�;="i�:8]v��wwC����f��Ԥ��_ؖ%�by����9ı,O;��v��bX�'�߻�ND�,K߾�v�9ı,Or}�r�3V�5�K-֮ӑ,K����iȖ%�by�����Kı=���nӑ,K���}۴�Kı<鯧M\��˒�Բ�Z�ND�,K���ͧ"X�%���o;v��c�PB"w�w��r%�bX�����iȖ%�by�gNSSA�F���f��ND�,KϾ�v�9ı,O��ݻND�,K�뽻ND�,�)2'���ٴ�Kı���RS�7i�]�:|:'D�>�_v�9ı,N����9ı,O3�w6��bX�'��}��r%�bX�w������	JO����L�\�B83��[����Km��1i�lH�:�3��͓p�طK�7$��m�ƺˊE#�Д�u�c[6���ŧ!�$f��!�6@�r<�/�=���m��p��]�P� ����]ٓOc8�DD�VV]��g6
S�\p��7(1��V�ֻw�����J��Þ�t���Y�����wm��58��l���[u&�O��q'����;y���l�Rn�ce�V2�\�J��	U;k�,t��y�j���q�x'���v�ie��f��%�b?k�۴�Kı<����r%�bX�w��Wa�Ay"X�'~�]�"X�%������A�����âtN��������?��,Ow�v��bX�'~�]�"X�%�ߵ�ݧ"X�%�|#�oM\5�f75��m9ı,O;�����Kı>�_v�9ı,N����9ı,O3�w6��bX�PU���""H̅��p�F�4O��ݻND�,K��{�ND�,K���ͧ"X�%��~�uv��bX��짾�(�k�]�]�:|:'D�bw>�siȖ%�by�����Kı<���ӑ,K���}۴�K�'O�@�~kR~�v�l�f�ݨ��Oc���9�;�9���'F�c;n�Xt�cdԳY�fӑ,K��;�siȖ%�by߷�]�"X�%�����iȖ%�bw>�siȖ%�b{��t��hѢK&kY��Kı<���Ӑ�~���!
�wq,N����r%�bX��w6��bX�'�߻�ND���TȖ%?~���d�.kAKsY�]�"X�%�߻��ND�,K��{�ND�,K���ͧ"X�%���uv��bX�'{�p�6�l��ֶ��bX�'��{�ND�,K���ͧ"X�%���uv��bX��N���m9ı,O��?�SY%�֭%ɫ�]�"X�%��w��ӑ,K���ﺻND�,K�~�6��bX�'�k��ND�,K��ߥ����Xv��1�kh4��ȻQqh ��2�8�u��s�zgE�g��{�{�oq��������Kı>���iȖ%�b}�w���lD�wI���XP5�}R"$�(�NH�P$P&�{;��O�,K���ͧ"X�%��u�nӑ,K��o��ND�,K�&f�S�8�r$T��p�F�4��7siȖ%�by�}۴�K�� �<��Z	PbE ��X(D�l�,O"w[�5v��bX�'�ٮ�p�F�4��&�3i�q(���m9ı,O3�w6��bX�'��}��r%�bY���}�ٴ�%�`x�"g�����"X�%��������4M2Yd�k6��bX�'��}��r%�bX~A=����O"X�%�{�ߵ��Kı<����r%�bX�w���MYvH2�m�޻S�s|��yp�Չ���1фu��N}c%ɹS�a�゚�ND�,K����ӑ,KĿ}��iȖ%�by�����Kı<���ӑ,K��~����h��Ku�ͧ"X�%�~���Ӑ��"dK���ٴ�Kı=���j�9ı,O�߻�ND���S"X���~��ֲC5�ZK�f���"X�%���w��r%�bX�}��WiȖ%�b}����r%�bX�����r%�bX��>����5�Ym��kWiȖ%�by�{�M�"X�%��{�siȖ%�b_���iȖ%��AO �(����'u�?]��tN��:=���S��ݮ�卻'"X�%��{�siȖ%�b_���iȖ%�by�}۴�Kı<���ӑ,K�ﺒ�ߤ�3�k3FA��u++@�",��R�ɟ']n�=��jۧD]��F�K��(;_:|:'D�=��~�qȖ%�by�}۴�Kı<�����"șı;�w�m9ı,��&��L�Z��`�)�᠍h(�w_v�9ı,O>�y���Kı>�~�m9ı,O���6��bX�����?��NU��âtN�O=�����Kı>�~�m9ı,O���6��bX�'�߻�ND�,D��ߏŶS�m��-�gΟ��8�>�~�m9ı,O���6��bX�'�߻��<��,K߿o��ӑ,K������%�l��Y��r%�bX�g��m9ı,O;��v��c��DȞ���v��bX�'s��ͧ"X�%���� ���Km�FP�0����C�@1��[��y���B@�������9���=ϊ�rl0��PRDV1X@� ���+y�7��A���hɍ�%�Da��&���3$l����L#	I`g<q�$���!e�sdH�RQ#�DI�$K��v!0��!U%#+5��fi	7f'X��D�a}�ĉP��4���MXJ��Ȳ/��t;�b�*DO����3= 1/�M�HZH@��<>��`Bo�!#��%� �$��"��0-�H�̓cp�ih[n���X�oP���;�_}�F&�pp��_}'�:x'�kb��K��i�4�\q��n��?}��Ii��RAF!1�5�B�"F��K`N/Mߺm	��(�<�XB �`FBH�6�%0{�aQt����[]4�d�$�	 �Tpp�Z5�*��v5�83�Z:L4�Fv�vH1��ǝ9'q���p��* �ݱ�8ԛ�<ؠ�v�׶���3�pʏ;#*�AS�:�㝶��� �9�kAɶ�a��L��6�.O��n��|���KM��`�9� AF���y�~R��G�p�y�g�lx.y���n0�ag#�l���ii�ծ*������c*w:���t�j���"�i�*�s3�E�`��������t\��Y������)F������L���F���5��j��;=�r���m��7S�����#J�T�s��m�ہ㭆Ӑ�����kd��h��k�j������O���WP{Q���l��Z�1q��\iqۧ�醫��r���u�mKa��j������9!H6|�n�+�M��0�n�pt�sQ��<i켳;i���8�]kh��ͮ��>Xu����� @�p�1�E��v!��և���f�Gf-�r�sR�	6�#b
�#A�i�������S�X�sL��=M��'z�1���d�lJZ�#6�%�dIe�ˡӸډ;z�,9�Ǻ���E�Ɓ�jl&Ў�6	v.�����gn��ɉ�gF�J匌��%,���e��kl\%0��d�Ӟt22&��>8�b٪����
mK��0g���Ă��P+M#��Aŧq�ݼ��&vny^��4�E����[V���(*�N2mN��ش5�����˂��v���)3Y�Q�:xH"�����ތ���Z[���h�3�	H�帺�=��q�&�b�<��c����v�4�f	�iv�-4�@lR�g����S�N�@�:/F�h؞���k�A��g�\�����aq��y@����2qAӹׄ*�1���&�.dy��8nxp<������H�����m��GN���2�XS�ny���P���ݕ�Jd��k4B=v%�:Z�m-*�7����I;�7K;�tꊓ�TB�������
~�T@!�a��py����R�sޱ� Ev|�8�Ru�@R]���6�d�n���W7ֶ0��v7���Qh�u��GC�y���r�f]�4�y��W p�lغ;f��۲lP�hJ�����CfcV�`G:�X�Vۙ����pGA�\!�C�Zk�a�ͥ6q�`��T6�B��	mB?1��2�G]�j�[Xl�-�� �JPs�M'ww��c��+�ԡ�Q�0c5]��m6�Dn7k�\^.��7
���(9�hඩ�~��x�,K�뿮ӑ,K���ﺻND�,K����ӑ,K��>�siȖ%�b_���j�֍L�u�]�"X�%���uv��bX�'���ͧ"X�%��}��ӑ,K����i���q���7}�|��կe�a]�9ı,N����ND�,K���ͧ"X�%��u�nӑ,K���ﺻ����t�O}�T�l5ؠ�v��bX�'��{�ND�,K���ݧ"X�%���uv��bX�'���wC��4��'�3jd���ND�,K���ݧ"X�%���uv��bX�'���͇�y"X�'s��fӑ,K�������]\՘��ރ9Ԟ��4�ۘ@Ғ��I�V�2���. gAB%v|����'��}��r%�bX�g�w6��bX�'��{�ND�,K���ͧ"X��F��Km�)��6�]�bX�g�w6��TN(�>EӸ��bf}�3iȖ%�b{����r%�bX�{��Wiȟ�r�D�=�9�cl�M����]�"X�%����ٴ�Kı<Ͼ�m9ı,O=�����Kı<�_v�9ı,N����8��Q���t�tN��:{���r%�bX�w��WiȖ%�b}����K����ȟ��߳iȖ%������nu˅�l����:"X�w��SiȖ%�b}����Kı;�w���Kı<���r%�N����z���e�kaB=��]�d�qi�t���Sh��r6;Gn(^��q�H�[Q����H��᠍h#C=��t8h#E�bw>�siȖ%�by�}۰���
��&D�,K����m9ı,g����T�62�b��y���:'DN���m9���"dK�뿮ӑ,Kľ����ӑ,K�����ӑ> Pj�4���u?�f2��"qŴ�Kı>���9ı,K��w5��K��: �4j&�}�߸m9ı,O����iȖ%�by����]KI2�WiȖ%�b_�����"X�%�����"X�%���fӑ,K���}۴�Kı)�)�F��"0Ò9t8h#A��w�6��bX��H���~�O"X�%��u��iȖ%�b_�����"X�PF���cA��$!H�$B�FCE��ʲ�ӂ:[�a0��y�*�s�ë���Gv3׉)��h�r%�bX����m9ı,O~�ݻND�,K����m9ı,O>�xm9ı,O~����p&��-�Z�f�ӑ,K���}۴�Kı/�}��ӑ,K�����ӑ,K����iȖ%�b_H���]kVj\�L����r%�bX���kiȖ%�by�{�iȖ%�b{�wٴ�Kı=���m9ı,J{����5au�(d�]�F�43ۼC��4,K�{�ͧ"X�%��~�fӑ,K�� (}D,B(?/��h�4/���4��}�4FbQHi��X��`wn��^�vb����o�Λ��E9����k�J)6�*`f���.��e:v ��.��Ӓ�U��]�wn��^�ɋ �ۆ��w�tʺ� ��R��K�I6v{ذ	%��;�p��kuLQ۳�ʢ����LX��0��0}�/ ��bX�+LCUWV�ݸ`���}�/ �dŀn�
e.�i����;����*^�ɳrO}�_M�>V |b�B$ �N�������7嶥�����g1"� �F[���b[4�*�ݷ�Dr���O�� I:)��w9��
�I��]�FՅ\�l�'�j��1�d����h�9/!B���'���ع����n��cd�����\�ZB03B�[)Iٻ[ QV3֗�m��Y�x�@�^[$27��a, G;&�U�6��.+�m��`�wc$!-���+nKWf:��:u�I\��,Z�p��[�Cێ.�Z:�{����ϓ���lX4��k���62��uuo@������LX��8��;���~Iq��D�ʭ���ձ]U]���,��K���<��<�����
	#���NӐY&�O<�[v��l���Ѯ�j���YVYWv��lx}ڗ�}�b���\\{�<��yx�S����wo ��R��LX{[ݭ� ���{�A˭,h�/n���Ʀ�:Pٶ�'8;��j�u{c�wt���GUw�}�b�;ڑ�����ԼwcƐ�[85Uuk �jG������ڹ�q'cڸ����`I1`yt�Z��l�n�����kjV\K����ŀn׼������:)���ռmmJ�>�b�;ڑ�����jpn�������>�b�<�[�<�J�x�=���7R�ך�7�B{���$��B� /<nWN�%��t��r�����\e�ҭ�x��ǀwkc�'i�q%Ϙv{ذ�Q���)J�dqY'�~�d��^�d'dŀokc�'t���r��i;��N�p�'dŃ\Z�s���1c! !#�������y��rO��~��C�n�2;e�]U:uf;&,��� �[;��ov1,i
���WwV���<mlx;&, ����-�w9��n��K`)����{���*#��l�N�Cml��9�q���7H1�M�� ��p�'dŀw�#��lp��c��j����u�0	6b�;ڑ�VǀI�����]��1���ً �jG�}+c�&��x�ybi�#�!#��$N�  �麮I�s���>�ۯ��T� 1�y�� �� �8���k]�<=�jX*��;�e���>���	�w� �kc�<���^�t6ھ;.����g����{L�n+�ݹسٻq�[��B��a���G.���)
wo�=�ߌ� �kc�>���n�ۡ��jʧT��� �kc�>ݸ`�uys�q�l�9�I�V�UU[�7jy�n�0	ݺ� �kc�6x���)�t���>ݸ`�u��ǁ�I'�s� :�.���2��ـN��x�[��ǀ}�p�:��\�Ӥa$:;�P�{��h�F��t�䭮^�0���q�`H����F��Ǎ\�w]B��ɥ��{4��T�;v-v�#��U�u����p�WG%��=/�S�����K�9�-�nяjp�Һ��X}wk#2ge1��z�b�j����X!�s��YIe��J[q�9��71�`jV��4#�w^b�����c2�]�5WY���={j��qh�.&�������;�zz��O���������ɺ�u�j�	�����u7#з&�Ĭ����:K���U���
�սmO<��� �v�s�S�O|}��"��&ґY'��� �v�Eݸ`mlx˴Iv�WN؝۲���n�0��� ��� ��Dq�9J�M U՘]ۆ��ǀN�ǀ}�����6�p���Tڪ�0��<v�<� ��p�)~�]���wN�;`p�m�8�lc��5��0k���+�,�K���A�GT�22��������y�����������=�����R-2黻�'=�~����	�CZ��u�]�<���{��W��=f��I)2�I�x�]y�mlx{[��ǀ��j�[��Uռ� �jG�}���y�L�< �O�캰�n�n���H���<n�G�okc�=���Z�­���B7l8l}W	�t�q��n�o;g��
B���ݨ��]�n+v]ݼ�[7n��7����H���R�S��;�Q������<�[ -�cmS��v�����okc�;���߳�9Ç!�X��CZ�H�|���}&�ϡO%4�	�!��K���.g�y��2��-w�rp��'�]y��\<�P��o�5�K�*4�	*�!�o���B>�����!A Gz]3D��r6MsE|5��io�����5	w�u�	�$�ܡHa��S57����9�s�+
JJ���q9�\����iH҅`��#��$�'_>i�1/#,fJ%癠�(���R8k�C�\=g04o[ =B��9�XI#n�n)�>��Bχ�`H��� ���d��!��T��0��E�&q���a�X��@��l
�fѰ&�O�]s�Y�!��57,>����0� ��xMy�]n�{��K��@D��`a�c$_��YĒ�CB
wO5SyĔ��R�_�Bf:�c���k��I���O!9��� E��0z����J�Xq�q�$ �"	I n���@�@+���/���I��@L6�@����p�@4|�a�i":Q�M���OO����|�Ĺ\Ky�]Ϯ�<J�x�bXRM�I����kc�>���v��\��s� ��晁bv���t���>���v���� ���������R�ݦ+A�dEe��vR���e����P#�bݧ��RGm'Z�U][�>�H<{[�kc���}S��'u`:K�	P��Q¬��b�v�<�[�jA縹��a<UU� ��M�"�O|�U�y��VI�^aVI矱Y'���dH�K��#�I�}���v��ݕ�|�xs�p��� J�R��>�~s�rO~��,��+��AN��ݐ��vV�kc�>ڑ�\Isg���YT�]��H�Y��G���K��-�Z�b����-��L&t�Eeq�DͶ�O�}����;�����~�\���?b�;�����+��C����w���8�ě;=~0	�� ��ǀl�b�buAm�����ˆ�cŀwkc�>����[���
)R��XI9����6T��>���l��B��mUZj��ʧk ��ǀ}+c�>�1`7�rJp`$C�Q�����s!�G��f�Y�˙�� �������dfa�S`�4V��g[�	����Mlk U&�X��;������j�̸k�(��. m��q���y��n���mqkm;��:�S��X��:�F�0���5��j!�YF�G�Ip�Y-�h����k����E�s��>����p..z�6�F��g)��n�h�K��+X���Y���CY���~�k��ܵ�Ɂ�0�b����`��[n���3Pm� �����d�cPD˅�!�@d�&ґx�����LX͏ݭ� �k[�5vhUv컻x�&,fǋ �ݕ�}+c�>��IRv�|
�� ٱ�����>���l�`��6�T�P��T�� wv^�ԏ �e� ��Q�Ꜳ��Eݲ�6ꮰ��x�\0	�uݭ� �c�6�w:!	c�8����Ԍ@̸SJ0�$C��҄�S�5�7]nA�
>�}��Mۨ��lx{R< ��A�X�L
�Uv`v�<���ÈI\�˚��]����v�x�LX ���Kn��J�[N��7kc�;ڑ�I1`����
���j�ui�U;��w���I1`u�0y��}ѓ!� �P�"�O337]� ݭ� �jG�.$���~|�L�v���ĝ�r#��Ț�6�=�j@wmsR��6d�.[p�\XLK"Z�_���7kc�;ڑ�I1`��6�T����T�՘�lx{R<�&,n��ި����wJ���]`�H��LXyr�����..y$��Ü��VG~0}��{4Ŋ���wMݼ�7]� �ݕ�w�#�����ht��UUk ���{�%�R�W@��~xݓ Hk��f�\K	�X�#bLiG��Ue���K��`⌶]��:�y��c��\�hݒ� ;ݗ�w�#�>옰	����&��V�v�������xݓ7]� ;ݗ�/�r��_��Zwe�j�ݗwo ���,n�� w�/ �jG�}�L%L-&4U]�c��	����<�>��Nl�D����	��0!��"�/��E �T><����$=�l�����n�ۻX���[/� w}��&�1`��̥�Z��]�/��,*���[<n�ޘ5�1=��z���χW��Ɗ���$A#�����VI<�d�Nx���ė>`l��wǆ�r�t4�v���	��X��x��y�!B���|I~�&�E0�n$�O�w�, ��{R< �d� ��6�
��L�V�5����ojG�l��M6b���7Un�hwh�N�� �ԏ >엀M�X���xx�ߜ9����h e%�V�4I��e���KSF9#�r�B��^�i���CvΚ'#�Dg`�5���?l��5�ґ�@
3����7�K��m�&ne�Z��Zκڽ�.Z��9� a�a��m���'v|Պ�p�	V,t��I�L�^������Q@�봊�4rk����i�@�M�8��#i���j�.��WuZ[t��R%~�ww�wt�D��M����b��6����8���5��5�S���k[=�؃��X-i�Un˫���xݕ� ;ݗߘv�G�n�B��i�*��	�+ w�/ ��#��%����R�Н;wN��`{���R< ��^7\ŀw�q�|j��Yce���;ڑ�ݒ�	��, �v^��3��t5t�v��.�s w�/ �jG�$����I�b�6�c��LX�8:s��4���p�d��j�GZ�F`"]�Ue2�MҪ�_��`we��H��\0�j�vZ�]�)֍�'����m`��A�>�K��ĸ��$������<v_�n�� >�N7v���VI����H��\0	��, ��z��]�WC��V]]��n�� ;�/ �jG�wJ��]���1*��w\ŀݗ�w���l�`}z��uN�T����ycd������ƺC�G���l��o7�d��Rb]Ee�4Jg[]���~������l�`��,�S���T圻m��� �kc��>�`u�X��{5����,j���v\0��=�l��U�|�C�EM��5�l��� >t���(n�N��� ��1`{%�>�X{.���2�V�ալ �d���+ ���n똰$��'$^��ڻ����@�p�;�qh� Yqf,��\��bŲ���p$��(��Nz����ɋ ��1`{���v:�:�;�wUwXݗw\ŀ���>}��[ӈP�9m_��0�s w�/ ��J�>�`��j��t*-�:uf w�/ ��J�>�`U���`F��ė����k(�d$� �`��!	h�k��[IY$ 4,h�DP1�s��ܓߎ��eσZ���� �ݕ�}�p�7�H���x���@}Ż����Y�[`PU�Z�h��E%��O^x4]u�<ጆ�mu�j���.�� w�/ �ݕ�#�$���wB�J���7�H���a�=x�=Xݗ ���E�`�Йwo ;ݗ�u���>�`O�^b�I�`IIP�Q��N�Iq=�<��_�zT� ;�/ �=���8�r��D�VI�a�K�A���vy$�}�ԓ�g���¨
���P_���
���PZ*����TW���*��@U҂�+��U`DPT�@�E `�E b AP $E b�DP*�P)@1�DP@��
�*��U@Uʪ��TV��*�EP_𪀪��TW�*�*��UU�J�
��@U|@U�b��L����� 1N� � �����!����Q���:}3( h { `�^��� �l����e��n�1���V+������� �,��@�A���!Q��=?�RSOP     � 	*� L  2` I��U4 � 44�4  <��h�5�      �(�MOT�F�i��i���#4OSh"D2���Q�56Dڞ���=5���2x��Ϯ8Ta���P[DA���܄@]����h�#�Y�QP�@�@��`�.�a"FYL��[��'}����N�8�؀�4�L��  ��X�睳 	 �   ]iU�������P      � ��� a$��a`�p �j  �3��E�P  �U�UV�����$5� �  $g  
, �����vQ�YDF1U[m�� E��7b.W�B�|n�㖟��a!g���C$�a�d��lf�0ܑ$ۄ� Q�c�aOu%�������A���5��F��ofU!�����$��3KhJ���Ɍ^ٳ��VxyU��f~?r{��+'�Ǉ��Jf�4��-?8	�UkS6<Pi���KB��@r�;�*���T�Ho-O@��\�{	���B�@�+�4I�RmN,�,�$�!|�>4�1��O �n��}����y<�X�o�O=��<v��2�a�Ϙ� �Cى�#QxE��lJ8��`�'��_7�z�c���|ƿ5��%jm��aD�\�C)0S7d�SF1mI4
=Ce�1-�X�)\��t�,؋esYl�$9�V�m�m.8@�ocB%��q�@�m�L�5f�魣lu��ĺ[�u9-�K�M�֬ۮ�V��άc�HX�LT!��4ʼ	�a�ݱ�ل�2���*��5{[���[e����iV�Zm,[@c�9�ԓSx�����*O���0˂��S�G��Y$=�u>�������o���m��YM+MA�Y\���Y�4�+nج	Xkk�jMBlGg�ilu-��z��Xq6��v�ߦy���k�5��4�P��m`�����m�K�w�`���ܕr��ں]��]��m��m�ںj[M����6�0���îp�R��r��Zms2�l�y̓��P{4�w��e`ٮ+\��ֵs�.μ��c[��c��#unKΦ�2�%�l�T�@�:����M�(��֤�ѽ7a��f�uf�ʕֺ$֭�ժM�i�Z��M��Q�4h0��n6zYz��mf�l]��6Z��,�F]6�~:;��PC��6������r=5<��Co�3��
��D!"rF'�=�(�N���H �sI�G��Q�� �8`F� ! �"�̜�;�N�gHI$�!$HI$����HLLI0I$Ą�0LIY_�礼����������J*j*j*j*j*j�j*j*j*j*j*
�������������&�&�&�&�&�&�&�&�&�"������������������������*�h��&��������*����B�`j��a8+��^����C���	A!\(��T���" i<
��J7�ʉIӠ(�zI���vrN)yZ[KU���<(�i �JMsfp;s��X��ڗwj]ݩwv�R�  ��             PI	$�K)[!Z�+ZkK��;} XD�����{�sY�c��33"f}�ݻ�b!�fffg��Γ�C�	=	�!�	0�1�	1z���H�:�-��c�����x�T�Ԩ�^���v�GXB]6m�!�@v��T2�(M�odYs*:�B���F���LŶ����7wĒ?]��{z������6�6�������h��6b�����Ӷ)���ʺ�̺̓&�81W[�l�������ׄK� ��Hܧɷ�c�Ro�>bp��X2�MD��|��3Oa�v�N�}u�^V�,п�����������g7��Md֐��/4m������l�r�˝F�]�(�������y1�m� e�� A�Vh�[�X�҄.�;�^%��f�p�.��ߓ߻�.=�cϘ� ��=� <6"\�(Ā�� �S-1�>�T���UP�������UY��wwǌ�7�Z֯Zֵ�~DddI$d)�톱�#?�U�x:6�">��y��t\ɥ���0箤+w�J�=��9D�RA��%:z_�G?~:�^�W�z�i,p�!���,�G�\I]�akoh$��9*��Z�xdF�������R! �����/�ܘw|^���v�n�!��fo�0�܄U��M=i��g�2��r�* :�L�@���)�R�����LC� �> ��t�4��E���.g��n>:C|�u���e����ä�2t}�(�a�Ā�hO�!�s1{�J!�q7<]��
�G�4�5n>������5
3�C
s��vfE��L�H 1T�Z���wUFT��#�'^&�͡��)��`ƬQLPD��y&���i\NO_��c��8�ux�0b30Dz�)J׃�9gxP? _iAP�g���iTEB���P�K�VW}�T�*ff��UDDEUUP��}�ۻ�LDt����5�뮹��j���
�E��
=u�Λy�(v�M%Q��T�S�	�m0�IWha������:�f����n��ecJb�v���Ͱ
h�ͺ��m�	�sX��߫?���{�$8#@�����D|�����[�Kb<�Y�Mnm�����lzB�U]@/���+>'~L_��q�o���o8����>b��\�)ex4��k@�"u�%sW�DJ�<������T�x�"�"!&f`�^f~�DBȀ�J�^O>�KI%�3��w)������Q�q��u�b�HJ�;���y��h����x����S�5�'q���P��4  #�p&x����������T���2�ٝ]sU  qƌwu�U��][|w�v�+ڦ��2��*L�=�_��>A
<0 T�r;�j"ٴ��u�4��fԓ;Mc�]���5= �(J@>Wl����U^9���#��{6:�>�R�y9h�4��Y�x��9�GM�E���/2�ffdL�DD��ɝ߽����"T��L��pHbH �X�L0
b��ɂ$ �d�F�*F-x�׃��vDP�r�i�.�� T8׎���f�&�(��7
��)�SN�$s3����)���	Do�GH�lOd���	<$�ǹ��_�����,�2Z����FC'O�PA�4u۰�YG܄��<{���O��הH���\ˉ�ݧ7Fd�����+$�'~/�q.��v��%�`$��U9�cp����N��1�ͮ5M�����sTs7#�2kU�5���ɰE�~0�?S1��Đ�o��G3�Ӿ�H��,�h�I h�$}�k#��Ř�Ug�H����eKZ:ƛZ�}ϗ��������SI>Їy�K�@P�X>f$k0��n����t#JǾ���k�Fa�wNN���m0�ܹ�;�w�X�Ԭ�[��j��N�ȏ3"��އyџJQ��~��(��e��D�̙�x������{۵��":fffd��y0��@?0����IE�ș�|�@i#�	�ʑ( J�$|�j>yVY���]�V�Ym�.\ٌWU�
��n	B�Ir�C[��6���[�V��,����Jl�_?�~_�B��,�AS���@��,^dB;�wwbJ�B��;�r�D��D:I��������m�uf.U�T�Xm("��	����q/�#��s2@����X�r⎞��qٟ'���Z��^[�\5}���R��ȷ�0gi�����'I��@����m֊���~e�L0��g�k[��X�ak�g�|uI_��>��s�)���Qe؟�9ga>#ۮ��O������(<pl,CEw����O�<I=2� �G��S3x�2�I���j�W�w0q��k�CI�����j�h̉c�����;��s%[����K�\�}V�̾+�:l�3�N{�0�S�uX$��`��_�O�w����������1313?�������3333�%�3!�"X !� C���e�U�C���b'�����Q]�~D�+3�m�$B��@y�P��<-���M&���<�� 7A��GL7x!���D�J�$H���H%&&҄��A)"a0�0�O*̞��{{�������7\k\��u퉌���|�| C�gGi���6��m�wf�A6%�� c	&��*�N	w���9b�0t�b��;.����* ��x�`����%�IYy���Qu��eqE���<�l Թ���n<��x��a��c.�E��������χ����D-���'��sx���vys�s�C� <!�CY��Z����]�_��/!�I+Q�>�r	ƃz���db@�_ph�/�3����^7hL�^qU�r���<n���|������
��n�ͧ_� �%����p�'�y�}31b&bfb""^eL�}��?��h舎��s���HE	 dyG�IEm{�
� t���2��	%"@�"3���F>x\:�m������휺�]�"�s0:��U����a��Z�Q�!	���v�����m���$�����<�,�**��:�pFߋ*j��3Z��|��R<>�����e<{a�H���x/Ff��8�1��K �'��ЙH'�#���-���}���T�T}2�=,�33o3}��p��~������:>�O,؄C$L9w��'p�O���Z��m��R�x�~�����o�b�v�Uap}Z~�\�ٽ����s�/�Y����7�x��WR�F,g�v�P�Z+L���C���Bj��!��W����+���@^�w|�q6Ob�x3���yPؚ��گ~Q���}311&fb""f$��o���}�3335�pl�b��	
B��F2Jh
����R���x2-KI=
�aڇ�"�3k� �ؖm:���z���PU4��b���}cw;�$�7������y�� �o�ԗ	@.��L\����x�.R1�>|� >z�sc�� ɘv+7���rx^�S�;CB�S`0"�mk�z�>���韯�A&���2(�.�� ��(h��wX)�·y�Y`�#�3B���c��BPC�:�Ә���y:DiWC]�E^���ǡ����5� q��q��ӮyH��5�L�����8G�R�DOZ+7�0�ʌ������:sM����;311&fb""f$��w����:"#�fg9�#� ��6Q�C"Ȥ�'��'�#�e�H�^�@:@NN �,	 F@��YFe�q	'h���/�8�`uSM���Jn�i��Եɭ��3D�R��ِ�Yf �e45�m����Ï�y9v��+e3���R�>0SUu�*�b�<rS��|.�ɢ�I���ڷ/��[�y�٩:�	���3
�� =�O�ueQ:�k����N"wpOǉԝ`O�
��3�w���]�t��p���[iJfR̷��f���`�~�G،՚�wU�|ᙆ0����̬�?�`'۫��^㛓���_nBYp֮W|+;�.�V>�,` ����|����\��*���f�}���/�C�~��u?��GJ5���0ӑ42����DDLș�����33^�u��c��9�s��6� �D�����x>7	�0�׿m�vf!>���=��;�oͽ��Ƿ�Ż\FV�����^�����"˵v�����M��I�ư�`���a����>�f؞���q!�
�g{y���"a��z�|��77�c�������	$�t��!��Ӣ��,��� �yy�_=��=������3],�!��3+����R~��mUv���O�N`���U{W}��T=|P�5� ~��H�蚪% 0�P=�^��q}%+ I��w�sZ:��x�<X+���U"���(�)�D��� �؉ �P`�fD]vm4MR"D �b@�NC[�)��R%
]�9�����8���Y.H���JMDr��"���%W��l����<�ꈠ��05U������u� ~ 
z��H�[�)��B�G�(� �� Pٲ��P�~���(�ݛ.�X�����yM�$��3��Y>��P��9(�� P�p(�w�+��?E�D�6�t���	a��}�z>?��ԗZb��{�U�����׾�Wև�h��A����� I!!>�@����G����R�+����8��I���Q���Gs���=�?�ւjUԒ'�7�}�*�)�!�MEEP�%T �IBҕR�CIITR1@D�4+H$��)(�hJ���HJ� JB�,�H��S(H���(D����F@(�_X8�T�R���1����Y��G��*��BnX��~�}��>O�$�硷�ۼ4_���=K}7��<�Տ�h��|�	�Oo��}��64d����ǣ��������|���S��ױ@��"(A�����t=��r۽S�9R "�v� ���~�#���c�%R{��'�=`82A}_����p�O�g� ��B��JcU��PP�LUQT��*}܇)�p���t%C�!�J .(�~��=� /w�����ࠨ_w�i���cלSA|�˳��o��������h���;���@�j((tr��l���=O	�<�ʘ0BЏ��E#p���?!���9u�I�ǳmd�͵ N���;�u_�NM�M�����O7�0C��g�/=��� �`�t{�O�6��

�ѻ���\g��A�x�����`=�?E}v'q;���ػ�)�4��