BZh91AY&SYˍ����߀pp��b� ����a}?��@� � 
P
U� �B�
�� B�J�T
 ��"* ��@R��J�RB��IE(R��*�T�*�����U( U@�
�!P��%)T�J�R* �     c   �
  V;�ݯ���Ė}��k;����N� ;�1�ǹ��N,;n}ܨ� 6��}���ӂ�  �N�.}�^��t�SҺ3TP�n�)��V�n���R��h��u(�m֛cW,*� h z�  
� vӷ����t�U���ܹ]{n����p�{ң3�j��ŏ��'��m��=�F-��W� xyzW[�R�p ��C�ݏ^}�H����{ۅ>8z�}�[����a�2u{ּބ��   �   b���%��`�>뼺G����.�M�i˺�rk�.X�ۗR�{� ��Pr}�L��(H ��ɥ��7ҫ� ���˻�ʼ[�]׌��q=�}ǉ�gT�������\ >�     (@a  ��}��0�Yv˟g+��Y�L�s��� ru�9{\� }=�O��s����t��q/8 =<<�olNXt�/s^'�5;���LU�{s�lx��nn��� �       � |���{�.Xtn�:K�7	`Ѵ�rj�s�|���\ZU� '=%�o�c�n }  ���y�=��p� y�2�����W w�y�*������x׈��ϻ����y���         "�Sm*T� �h  ��"jJ���0 3SC@"��UJI�d�#@��M1 �b'�T���J4     ����M�T�Q� d�h B��*AM'��S4��44�����/����w_������G^���`������AAU]�*��AU_�Uq ?�
����U]_��r*����J �������j��������g�oe�x���'c����ާs8,PJ!.Ʊ8�k#x�2i:oo3�W=a?;�]��;����yGPȔs�tI�ŉ�!&��4.��EpTL7�wv	�k�F�y�-OK��;3�7��XS���;����{�|�[���J4��<T�QM}�,�1���l[���]sV�����&,�2�OQ�����.܃3QBw��YrĂ�����F���r���KNP�%	Bj����5�y�{�׮k'�#�W5����Ms�v�s��=PT��k��>����u]�x�;�'��|.��p.{��[9��U�yh��⦾9��'�"���k�츇_��(J��F�GPa���L�5j���M��UV�l�2�z�����7	I�r�ɖ&U��NHfQ�j��N>�c�J�7�����1d�d%hg ��w�2i�䆲�2���ɝ�V�#!��CY	FCd%���A��S޷�#8��C��k3:�w���Hi�kS�`(����7F�����Ͽ\�]�g�;�k� I4ʳq���w�{���{3Ls�ݯ�--�=�@�^׊�w�������rUEϷ�BHSFV�#$tKT���&�E���A�����I�qs⹓^J���5��f��[��n�l#7�R�	�z ��Ȼ�ܜU��kÂ�U�߶o={ ��(�[2q��s'[N�fAb��Ӽ�5}۷�Ž��v�x�9��A����cL�τ��\_p���>ًy���b��-F9W�pX�%��*.�sZy���Y�\��x!w���U�E���q^��y�Ͼ�����7�%����.�}���?�55�X�b��˳i��)�5�[[#p�f���u�����(O*�Q� �����! (<#S�ż����C��0��dC���i5��5jF	�'0��`'�[���6'��$��9�/��6=���6�9�j%jE����E6�朴XA�Bj
���`�$H
�j(�!F�h��0X,1!
I1�3�n��W��(���||���܏]��P�i�k^'2���׫[�H�^��]�\�N��~\k巨�s�|,�y8�<�	F&:���F���A�6j�`�����)՞ޘ<�-ffa�u��AF��O!5�:}<��ꍛ3V��̌؄�D׌\1�I�r�53<f��E��ğ<>n��f&����V��&8�����1J���/�r�'�|&�s�5�g�qL��e�L�tN+��̩����U��-S�n*�WG�Z3H�Ovɋ�&���*�w���z�x�
�հ|���}]U�)�"u+CU�s[��WV���`�j�4��5��*ϰS"�\L��/��K]�ހ��4�D�J���Ъu�lI����&`�[�px��ւ ��9ۘsv����٣��<�k%.�(С1�]-i&��U.(�.Nbf'8�Q9���Nuyhٷ\�NK1�Ā�j��+��A�}�V�'"�O6|�o�7��$��uy|q��b�.��>uA4Ğ7��<�nTD�����855�q����7��_G�� C�+=��榮��(cm�.�ƓW>���U�������"�|�����㈞Κ+�itϓ^�w6>���)�=�M��[����@n7�k0�1i`�]���N��Z3�VwM�Ļ;3�s˵	�6���g��1�ML������2�ߙ�����_cfP=J�T]�b���Y��|L�R���2u�)�l�3�|���(��P�`�ȕ�2c2��v��C*0LI�D2-�B\�K�.���$آU/�k��E���O>硘���I�N�z����C�7˝>�j��Ὣk��_9�{=�uq%W�Mx��|jNF��16�CZ��\�5����.FI�Z��N�4�;�O$�8��w��s�b��FO]:(��:�Fj�i�Q�l���Ԡ��_&��y5";�����.^<�V�zs��6��~Q��;�:��Ρ��5�}\]����m�ŷ�"i�A��gV��D�|EQ �	�� a�8��s��F}�����b^߻�K��?����f�U���1��ɫ��.����J"�4�2V���t�����s��ߞ��U�\2%̑���ʳ��$�&(�!ʢ����/�8���Ѝ�~�{�o���}����7�)j+3�FF�1����7{/��(3�L�*L����.�nrvh��"M�tt�<��lZ�n{$�ܗ/|�׍l�Hrг��߻ީQа��{�ﻫ���;Q��-�|���w�$^4���Sa9���pC*鋪j�	��T�^��d:#�a�v���Q.�Ji�2�\ȅ6����ϛ��*⋼���/��;�pZ���r>��Y�X,i!`ߦ�|�L�q�6&���+ԺGHP�'P�&�;�J���Ǉ7�iC��-�a�7	YENBX%	Bk0JJ4e�K�$�15fb�|/Vq�a�ziD�f�Ow��v>��zn�{��9�0��'ryj��j_d�K��..wT>�8r���w}>��f����.|'��.qV$`��4(���Ir$yV��I�՚I��2�PE&.���b��V�U�dMCj�_{t~�>�9�e꽜Tӱ`�E�k�����\ϖ�����M9��9�Ȼ9�r]�� ��I�.>i�gWy�y|�s��Z��{�+��yb03;�x`��_,��ŁD��9}�WV��b�bJ�j\�:�B�oz<n�4&���5�U�#4{�¾�>�|�Q��.���C��驛�7B��B�Ů5>���7�B�*�����c�s�kUD�j{�Oo����w�9��떴�e4�Dj	��t��-b9��|�����>�y��߸�}ʐ�e�kj��8qC�<���[}��ؗ7�-�S>j{�o����I��/S/�����A�-�/O(��:Y�w����O,m����I��@Fd0xHxP���]��w�s]�:�|��Ɠ�j$�x���ԃ����X��`j�8�7bɏ"���nn�(�5'*��b���;���̄�,@�"h��5pA��W�r�G�]�A)����|��ӭ��!�f5	BP�C���l�,p�C�e�H��z)[ܸ����xcա(	K���%cMf.F@e�� �)u�â�{�[;trxLd�N$e�9S�tkY��z��[xh5�2��pl��(�����h�����S�	�Dy�6gC(����z��\����d۫|��M3��<�'�,F�����TĢB�k"�m�*�Tڒ��M��J�MU��*��*'$0���5ļ�*�I��s�ރ��L��y�ڍf!�����Ĝ�,���s�dԱD�hm��0vcdc�� �:����^2j���i�w�R���'~Z��w�ʯ+k�P�Y9T�H��E�����]��ԓ��Ȇ	�sj߸���=�["hr��H����I�N�]ܧx��@�R:d�nX��c�J��;����T 20�,�� HO7�72���f�޲ߖ�ӫZ$�ZB@f�1�4���ϣ�.�!�gU4�(	�<(�m�@B���d�a�3#���yԱ���!u1��H���O��%IAb���X&�ջ�i��c+Q�r3�Ӛ4�%�9y������g��$7�����L�R���E^%8}3��p�#x}��D�Q�PHπ��xx�MY>��_cK�fբQC ��"2/V��vE91�x⢯6�eI1|dȔ�8����Q}�P*��~Ϯ��޼8�{��=��ƍ���2`���Q,W��m�:(���p`s]���(��OrO�1<N1\��P�kl�ע��q��w�{��&�#.�+�¼ԅ �]Q����F 1��Y��p���&Bd�c�C�e��LX���&�O��b�&D`�s0�n#������gc��a�N#ɷ!�����|�Ż�E�/�S���կ�ӱ
t�>�NB#��!��JĆ�:Z��s�	O8��ME�M%���q�L��o'ph�HEA�k[�A�0i�ǋ�k���p�ο�-�pi����hFJq5�p:��ndx���e\L���>\�	�dI������{��`(,j(5����:�W%�s�EEm��2�ę�յ!˸�x���LB�5���q�ί�Z��5�X�:�D�M�e�~�*�x&�1��&�S��I�VLԔ�*��3�(��TN7#hM��!�b�wʍ4F��B����b%��c����.n�g_'� ^b: mD�v�:�P�&�r��ѻ�W�"9S��6^.ք����q�(�����z�N��M��T�Q���B9Õ(�]��bf0|Sx��#+Oq����G�1�n������.n �1<M�����'Z�������1��N�P��@ĝZ1u	H�%�lbuSu',͂ȥj#G�	��53Unړ��;3C�V�����a��w�:�"5�e��d����}{�dki���jLF,M�Q����!5>�kSk˿ww�	@5�0�����JՌZ��PQTH����H��5m�N�h��*�t�e1��J�՞�w�4Ԝ��BF�Y�,PI1�	׻�K�Jʒ�`���
�:f�y�dS�쓏|�u�Ն�5n9���������'Z� ���FX9�����<<���M�	��*r��GT�s2���и��n-u���k m�S�;nc4/G漼��7є��=�[���؞����ba����u��xk��$4��)�$�X.EC�b���&�y��Gba��F&�Z'D�EF��46��ȳ\�8Ew�;�9Ũ���uΏzLѳ�r:�l:��E�<봍�氊dJ ��i�˺��bV[9kqf&���k5����Gs��$3Y6BQV��Z���8N{�]9�Gx��X�*BZ�t���:�i�]�w��Ź�&#΂3�&�Uf��� ��}��ӹ���]95j�t��փ*�ORd�*2��vM����A&ۙ�<Ȇs����/s��� 4�!�D��>\��\s�U�@�Z�9.�v4ٻ�L[�|Z%�$bc��дj��-L��DK��J���f?���RmD�d&б��s������b��n41��aŝ1&���㯟�=��}o����lH         �      pd  i�m�     '�d  �    �    �c' R����P�  q �sm��N       a���H[im�$�k�     H$�[xp d ��%)������9��2AmUv�v���Mn]�j�X�vUi����\�\� �d�i�eX�^���R�t�6n�V��v�Niݞ�f`ݪ�TWg�Ð�T��4����j6q��^�1��

��>wf���%ݞ���c��jZ�lj��U�k�\ňɗd���X�ճ�n�m���r�_�L܎�z�Z����r��������J�WZ�^(�{Nd���6�MG M���6{/]]b�@.s��G�z�t�ėu�@I����^�l��Z�r�C�-T�yKn4�*œ�۪�]5�m!4�V"��]T���]UU*E[X6�C�U`��P����H�"��:e`h��h.�en��T�=���U�����meӜ����@�<��j�pJ�bu+n�O�U\�p�P���� V��K7�����m��g	��m��J�S�pJp��K��m]U+*I��e�����h�  ��f� m��M� �������b*�`ب-$݀�c����l��ۛ��	�;�\�]tڭƸ��<;Uq�m�I��A�C7]\q��� *��N��٫��ձ&4;��9Y�J��IlFƉ䝯4��<@+K���r}V�{�K�By�pd��f�u��YeQ��g����sm��nݣ9��b�=���=�'kQۭ��b�����s�U��S��n�j�����6ڱ�������  �Z��શ�5r�����=���2;�9�u^�b�(�
d� �i����M4eo-{��R�=W��,�Qy6��r�:B�\��Ҋ)6ʫ�T�R��Q�T�2�R�=��eC����ݹ]�����؇��e�U�jw-J�]]Om��^a/G[)�sm�]�Z��L���UTpU���&�eV�+iI�,���ݪ����RC�80���)Snr�e�Bez]�4�NP����[� �k8']ס���y������&�N�m��A��� �&��͵	x\�R�T�WO.l�we8,t��v�:@R���������K�5�j�o0�m�D趀U�i`�\�J�UR�� h��>7���EZ�����]����buŵ,��[pmpm��9�-궅�0,�'���uU];\c�Ш���6��ckwH��[$t�܃(�6ڶ;m0P�X�m��8rMae��Z�&VB�
���  m�h6ت�b�)܆�]�AJ��� {uC��l�]N��[#r��͛:^���$���� 8��Q¶5Щ�HUP<ݨTt���V���5Mcg+��@I��c�&�6��t�ݴ�j�"Z�v�1R�n���;��u[�j���M�j�1βg�]�s�L��v]�w�ͷ��\��z
�4P2�u��[Κ8�f�*K���t�iKh�WN8�/V�@��v�֘����,��L���Uə��}�ꋳ�k�7�5�n޹�V��
�.Ύ��%�g�3���M�چŪN� �kMME�Kj�q�JP�֩�u9v�;:�V[��'�<�Z�㗚�^vjn�Pj���NMS&�.˳R\��9�[p&�K�cu.h6��mg+�mÅ�r�k��̓D���iamV��#�s>�0�̓�.G��p�UU@mUt�:8y�\��n&۶[���okՀp����KT��+^�J���9��ruuӉ��ꩇ2�k�� H]#�k2�����V�v&ݭ!)��������J���UܫJ櫈�6�:�   �m�4V�]&�b@�l��%fu��A�m�Z��/i[m�L�I�\ԧW2��+�
�յPJ�ևHH^���m� ֶ���/;�щy�<�q[m��Q&(�QB� �r�Ӟt��!c`4Rg.�#!�L����Y�z�s�X���U�ʡ��We|�t���i��\�Up�4�&�]�4W6�D��s�Ѫ-�ܳWRq+�DmU�YӬ.	�U�E �X��F�YpHHm��7+Ars�Uyy��Y[#�C  �]�]Mu���Q����B��j��@v궕j�'�
��yn��m �]�Nն�lu��Uu5%6���8��0��ƍ��M�mU�;���km��-V�%��U��*���H��
�Hm�'K���5���6�  ;ݽ���+��a�a���cb�q�����9n�k�\�l�� �  �$
�BiV�yV���`m�&�6ض�ճ@�ȧ]�cD�q���q��;D�IN�e�iY�
�UL�0 �J�vF &ݭ�2Kd����v�i3l*m��l� - b�@��9��Mp�	$Xd�p m��� �ٽof��АZUt��k�FB9yd
���T�`$p�����f��6I%�@[� -� t�26�����`n�	r�-�n�6ZlpHzz@:�`HI�Ѷ�R��]U!��;�lL�R[kj�������� �[B�;[�L:�*��T�
����( ��vض� $��Ѕۤ�2�َ=m����N������$� ��J��TӘ۷=v,;m̭����U{okk7$�wE�ڷ[(�js�N��6���u@U�zG��&,�xĪ�F�j�� �K�m�]%�^t���i%��]H ү[m�Hm�5� ��ɳ�䍶�aU�㊹V���Y����bV�6= $��\��n��3���k��6�b0V-^�����kډKe�A�2��O��n�g�3\�9y��Wk��$�SeQ4�rdݝ�ғn�xh��Z���k �Rnv96rm��"�2�����uJEF���$U\�-����o��ɮ��*;���8�x�8�7l�nl�
���ls���کV󮒅^5��aػ��t�)ÍuWQ�X��HK��zV	�j�w�䂣de��1��.�\�]U*Ԡ	K����ck�[Tnl���takk7R�΍"^��u��Yр���kwͮ�>����@*��PlB�ef�j��t����fs�&U��+�0�pp;�ڪ�E����m�G�� ���M�d�ِ	;F�L�fibZ��,����l  � 6ڕj�cj]��jBkj�`�H  �*�ң6�yZ����p7[wI[��o����B����j�Rkn��nUk��=m�0!Kr�T��<��-WmU*l l��UJZ˂V
�tH_|�?AKU�[�j���`6�V�`��U����]\�M@J��� [F� m�v۷dv�����K��km�F m�;nX6�:��Sr! ,R��"l�i��������M԰W,��*�+i�-�!4	����N�����%�j������UR��S#���WO�r�pb�CiRY�R�x�Җ� �nͳ[Gt��
�՜9䪔pP����v���げ�f�<�J个�D�!��+��Z���l�\�T�v�㤻G]ѓp
�H�mzNk�0������dn���g!k	�f���h�"���,�����/��N�=��]�4��WUmR��P�Z&��ەjUU�j��Z��7)h )hs�y�H5��. 6�;m��m��V����E�V�	 sm���lpUVҪ��ʧ5J욗���a@p m�I�v��
BUU	�ێ
�;nŵ���8%�*�N��UڪڊЉt/<�֥	�<ǩ9W�Z�&īO9�y]�ㅰɁ���H�� �J����$  v�m�T��ʪ�9�Ҷ�Lj`���B��� m�� ��UR�Ny݃Xd
����mH���`�ғ�Һ��Ь[@ ��R�֢����i �� ���%�{o��`�M:6�k5U՚�V�D�m���6�@8$-�Y��]�k�Q��;Q`��
��fʴ��d���%� H�pڴ����Z�3!�Ev���m �v%�qO+P�Ĳ��4�kXn� �<u�����C.��2�km�UU�@B����_f�8p�m��*�n���R��l�n�m���rKh5�ۜ :���Fj���(�m*��YV�5��Ult�l�d h��yd�������s��1��bb�T�U��֡�ՌH ���ۥ|��ڞ&(�݇�ѳɒ��Q��p��g�2mP� NȭWl���VԾ3tp�7m��[x�l u�@ mZ�J�#�MV��'��ڱn˴��vֻp �]� U~U<��T��U*Ԫ�M��P%j�8 ]��� ֶ����, 6��lM����`t���gn�H�m�  �I�ې9\`a�j���b�U��yZ`�#R��Y������	����j�9u��@   UT��R�@K����� $H 6٩5Pb�nX�E-T��Az�pq$���3fؽh m��)�2-���Jk.�һ>ْ٪��(u<��'m�DOJ�jjT8j^N���Z�jNM��lF�zQ�3�g��ݖ����^Z�������6�]�����ƴ�h H6�fCY��n�\�հ�J�z�FU�6��[�:;R�Wjz[<<�t�����
�U5*��� i(�K��R*��j�s������{��g���
������������|"x�p�4
��������?���)*���п�:Y�I!N���"��:a:T�:�!�B�:T�E�v�+�W�@4��q ��Q0T���� �@��
	�9��2J@ `j _:Їn���ð�p�qI�$G%�\�������u�/� <���N	�=��^)�	�'��p8���'��j��"��=UHTCB��uIȒ�hU<M!�L'��!�;Mx=*�{��a�zDC��C��b/O�p{Wr�a*b`a8b]�i4���*/I�H(H@I"D#�:8��¨>�hC�; dQPOeU8#�4NiPࠞ(��� �8!ꊞ0����$!� %	e"���X_0OGGj/�)�0����kэ���ꦔ	t(;���v�)�� �R�Jv�������ib��Y2H��	`�ɕ
�@`Cj�&���
��OQ{E}}4 i��
��bb�a����i�N���8�a;G�+D3!$�b��������@=U=A�
�H�
����3*eC�9�.X2.J�F���0Nd�f
F8��a��x��.�<�JI�BIB��P�G�)@��	�4t��Q0=�CHBs��ivz`K�<z_ܿ��J ����O������_�dT�*�!
@BF����
�̖?H���"�0�"2��CW�2
i%J$vH�`��k� [@3k͇����m�$��^�[��P�e�JZnۤ�Z�Wl��,��-cq�n7E�ˍ�W/Y�h�5]W��&��.�-'H�C��i�乻cn�c��5�CV������i���x3%�#�ٚ�8����g�1�l�l�t�l[>ê�;���Q��]$Z�'�n�B��̭�ۥ3gƋ�r<����n9�Ц�E�'�[(�3u������LAc\�gpV�sv�Y[I�f�k8�6G�& ��m�+���ěmG(�<�V�\mt��W2�A��UI�&��GD���O9�Qz�:O7lOd�[z�qJ�.�^�tg��q�jK��\�un��i�KE�KC��n�Q8�V�8��m�8��i�N�eܬ��n��U�*Z�����hk�x�2qn;m�n�|*�zҾ��!�S���ѹo-%���Z�JcX7�tq��A�$����m�z\c`:Żn�j]�\m�!L8�s��Q��v�h	j5�L`D6��.��g����g��Nvl�n��$-��6N�V2�qF�4��b<����Y�F4�*TwRU֣m�C��ڣc��}���bݕ��]"[s�uR�eU�S�@�H�ysAݧ�{=��9ۅ�ur���ݳ��u�x�\�3v��e�����H���qŸ��� .��y��$�f�c�m2	��U]�LK��A4�$�ˡIPJY�W�����+��;
��/�ڠ&Ĝ,N��m���W\g��=�tg��S�:SŬKNn+cD�.;m1/2(Qխcb�8K���q���9���z�S�X� l;ջ�[\�\)��j�G q���v:k�pu��eg���m��J��]���ۋ�����E`��l�Jl�ku��yzJa��vyN�<�NҨi�	�@�ml���6Ԩ��n��r�9kl�q�X�����A�����l�V�Ԛ��nP������rU���rYT�8��[l���46�o���w����й����q&�����t�*� <P=P$P� |>�v�i�� ��dP�/��2l��[`ܤ��\��I�Ti^N��N��Cr��ڨ;X�mѲ��7G`�H8�l��c�e9������岝q�ݮ�Y�gl�/n�6y���p�+m-!��:U8ٌZ{�����VSqVԹ�1�f�g� c:�+�,��m��R.�VY'�'�th�.�͌�y��1�Ԛ�1���،'
������`�ͬY�����,�Eؽ�⎸��0�"DFA"�G�����}�x�9x�{�;��J5l�v�C����Ͼ������/�����< �/�Kʥi�]���7��kL�}�� �UX}�u�����:��Hݕh���@=�޺���{����|��9�Si�^�{�t���@�}�Z;>������ʪ��S�Kt������ڴ�}���]�ŋ��s�mDKnc��9�r<���};�c��pS.2/[��m��-5�.�6��������'���>�}���] �}�|���TYGk���-�@�g�{䗌���������1T�}���7��������{ڴ�=��ݶ�MRM� ��� 7�焯�UWs�e`����q�ڪn'dr6�m�w޺��j���] ��z����y�J�� ܒ������� ;���s�%U_Ǹ��m�'@uv@"�%��պ1�9�p�e5��U�]�c\N�;d�:�%v�jδ�����x�w<����=�W�I�Sp�� ��z�;�]���h{���K1�_������E[��l��~���ｫC�8�I�ł�$ah1N����o��>��@�}�؉SUJ��e���j���] ��z�;�]��yL���v:u�}�x��< ߻�@�}�Z�X����bq@hq�*�i�ݼ����K�r���r�[z��7>3��v\�Z4bջ�����v�$��	� o�� �}�Z����Z�V�\�����3�ڴ�����V��j� �{n�yy����R8���ｫ@>��V'x�n����X�mhODR��H�@;߽t�}��t71��>��؛G�����ʺ=ׇ��j&1е7	-�}���s�z�ｫ@>�޺�����1��m:�E�p�C�H]��B*v���ǶoJ��T�sj_n��2��qT�� ���=�{V�}�s���l	���;�):l����;�� ����s��s�=}�\1'wi��Cn��{� w��@��4w�ՠ�?����e���oW껝��_�X}ݕ�}�z����%dVI$m�۠q�ޚ��߿qp������@�&�bOI<K����^���ue�j�6���h}������.~-��{p�������>����+06X.��p�a�O�Y<��(;����<��}��Z�L��z�'f��Y�=�{l0T���v�������5��pf��\l���W[��6���t���:�q͓\�೸�NZ����eW�.q�mkZ)���j���TjR\�H�C�׻ݻ�����1�� ױ�[�%k�ݹw�/]�L�WRey�M[��2u�F�*��Rv���b-$��'I���޺���8��M�G����:����X����Uv�<�� ��ڴ�<����jn[���]����9���@;߽t:���U�T������9���@;߽t�}�u3��m
UUR�@���{ڴ���@;�޺}�~K1fu|��?�pF��zTCu���s��^I��jz`nݐ�t�H�c��ن�l�5�mր{� }�s�6��R��V�}�e`�Y������j�o >���~�B}�5��$l�VQ�[+[zY�K2f'���n����V�s�z�����%dN��#�@��ޚ;��h;���s�z���잰�G 䙩�N�����cX��V�{j���ڰ�;�)?�hTА6� 7�s�%��@���`��+ ߺ��AZ��8l{2͐#]N9��<nn1فM��λ7Z����ŵ�}�ߟ���_�߽4w�j�w�] �/}<�ʠ1S�M&���� ߽�X�{� o�z�O��VЭV��@����ڶ����|�  ����䋥1u|�{�{wn����4�OO��ݦݡ��X�{� o��m��X;��h|����l��n�s�z�}��@�~�� �~��;�����q�5�q��6T���)�]������r�-����2��xQ1W�n>��s�{V�s�z�;���|�����V���I7�o�쬗a��< �� o��쒎r��;�I��6� >�G������x����=�>�%B�e�n�+M�K�����������h)(|� 8�*zh��7�����L�"��%����~��t�������x�W���j�LB+��s�i	S��6�]t9�:���ܝ�mz�v�kb-ӂޝ���7F=�||�ϟ�@9߽t���@9߽t�Oz��$e�ݡ��X�{� o�������+ >��s��wv'm���~��@9�޺;��h>��@����V$�[WiZ��x��<~�e`������@:�/�zC,#��[�s�{V�s�t���@9�޺�yx���ĄdM�O�9������C��k������m��:�f��.ݍ�<S\�qk�u�n�u�@l�W"��S�T���%v�����q��
t6�瞯L-<�����t�sy�u��%��n%Ė��s�ˮ�;y�v�Q�����%)tQgf�p���h���s�v����z:�c$jy�d;g�+���?Uˉ��ZTdv��Hn�3g�mtg�R��Qtj���wo^��ɠ���,>�J�n���iCRe����sx�ͺ�m�'*[����Cn�?̷I��6��w��w�] �~��9߽�@�x�ȉ�t�I&�~�< ߽� ߽�X�{��g}=ʡZ��,��;�����������tx��<�|{�aM���P��;��h;���s�z�;�<�����5i�6�M:�������@9߽tw�j�9ߗ����a2v����m\�wg��mx��K��w[ee��2�[[Pq�MW�m�����>�Ձ�{m����@{UX�Q�J��rB1۹����X�����#��c8��C��~u�||��v����C��~������{s���7��ۜ��\��9��Q�(���s�sy߽�Ͼ���~���~^*���B�%�[��{m������j��{iӻ�3g��)��`���vu@u%8N�Jyȯ;f%�N�t+�<�H��ά��g�\��\Rߞ�����9߽�Ͼ���}�_O�F
�VEQST��{m3��n�|��[�i;���*M�I(�U�.������ڱ�����#��=5(�������u�L��u��k�/��:���ߞ>h��~x}����GF����뗽u�k��By*F���,�b��=`t����4�p�	d�c���*������C��履bbS��pfu`%�q(?��'"��w��0+Ό3��F>�Av7z3
1O9���gXs''��Ȝ�!!+����Cq�#�SpP������zW�x��M�:�6=�z�<	�bELAS�9�y��	�!��Q�f����ɥ!���>	M�|a��l��H*JH4�3����0<@���>��Xb��H���3� j
���ݛD(_��8��i���R�l��]�e�t:�:O&$�����㨬�̣�Y6����h,zIC;�)��+7i��|���=��D��|�t'�� �^s�E�G$,'�qC�<T�  `p]*t*����?��1t��a��R���o�R��w����)K����y�o0�f���y��|R���>��ԥ)w��o�R����pz���	s߾��*�?{��XX�q�����ᘉK�~�|R���=��ԥ)y�o�R�=w�pz��?�W?��lӗO,i鱎z]�Z���v�z��'��������X�M������v��m��^���ԥ)y�o�R�=w�q?w;�;���w`w`vK����jz*I�"����R���߷�? �JP��~��)J^{����)I�~{��?�1~_�TD�:Wk��n� �@��{��R��ߟ}�)JRuߞ���R3���w1b\ί�?E2���Tn���R��ߟ}�)JRuߞ���R���߷�(H��Îhi�1AJ�&�d�'~
~�U�������JS���ܲ��v���ս�|R���=��ԥ!�Y�=���,����ږg;�\şp��o�X�fU<<Zm��65��N�N�*U������Үy6�Ƚqڹ*.r-g���x�����)JP�ߞ���R��Ͼ��):��~��)J]�^֯��a�ʪ�����w`w`g_{U������y+�JR�߼��R�����)JP���ߥ�ĬQѸM�.���3~��w0�)=��~��)J^y��┥�y�ڳ�b����O�Q+Ս�e��
R{�����R���߷�)J~�߸=JR����┥'�zV{��w�Z��Yf���R���߷�)J?*$~����)O=���R�������ԥ)�|J�q!&oFpt��!) � �iTLdMj�;������ΰxf���k�v��&�邭����d!r�l�{]nI��\�{]�����[�vA�n:����fЯbM�{u�\�:p\��`���ہꮆ�-ϵҬAk�;�<=�m�a5����:���z�����[3S�m�n����Y�ђ"�,�9�:�g��\��b���9��b�F�5��P�A�R5�c��um��N�{q�cYk<lxt�^�~�X��,��֍8�a ��,�rK5���tuۭ�r��1n���s��ץ\l-oE�Ӗ�o7������R����߾��)Jw�}���)I��{��JR��~�����~���TU�*4ݻ�8f ��<��qJR�����R�����)JP�ߞ���R��/߷e�홳fV��qJR�����R��y�k�R�>��pz��{�=�\R����r�ꫪ��˖�e՜3f.���nb(}��~��)Jw�{���)I��{�p�A���3���Ӗ[l��71�>��pz��?�I�^��\R�����~��)Jw�{���JR{�^W�d��qr񋋆Ocv���tF㗷1�^:�A�u8��B��u���|�=��`s��}��R�{�=�\R����=���	Jw�{���Ee�J����G�JV�9�GCK5I1D�35Sn�����Ǩ����:6�%5�����)K�~{��JS��ߵ�?��������KS5T�DEU�����ލ]6�ԥ�����)N��~��)<�Ͽj��3���٪�T"��%�s)C�{��JS��ߵ�)JO;��=JR����)JRt}^���i٣y�[.\����R��<��qJR�����R��y�k�R�=���pz��?,Ē�^��H���嵀dR��"�l�g	��X�\�ۗ��'��9K��1ڭǪ�3f̭�z�JR��=���ԥ)�y��┥}����)N��~��)_}�{�U�GKej�캳�b����k�R�=���pz��;�=�\R��}����8f �]�~~N���I%��R�>w��pz��;�=�\R����WDf�k5R�d&4�{�U{�>����)J}�����f Y�}����VGd�v˺��bü�ߵ�)JO;�߸=JR����)JP������R��/�L��k7j�k[޸�)I�{��J���~��)JP���߸=JR����)JR~���_���(ě�4��b�v��m[�;o<;D��*�[a�Ӯ�Ƴ�p�g��7]�IS�Uc?û�z5tۻ�?��cԥ)�y��┥'�}���)OX�{�U� �*��-���1Ͽ{���)N��~��)=����)Jv��鹈3b��~���TV'Qu�wG�JS��ߵ�)JO|��=Hҝ���)JP���}��R��/�e�홳fV��qJ�߽��R��y�k�R�>���pz����*yD�� H�+'���BW��ٹ�3b���ߪ��:[+V��|�)N��~��)}�߾��)Jw�{���)I�����JS�9��V'c���<��grx�]�(:��f-[]e`6�ڍ�	�쮋��=[��	�o����[z޸�)C��~��)Jw�{���)I���� �R��<��qJR������UĬ��$뛺��b����MIbKJR}��߸=JR�g�~��(}Z�������A�
Y�I�$����R����~��ԥ)�y����IX�.�g�݁ݽ�m݁݁�w�	5YTI�:����b����M�A��}�߾��)Jw�{���	�D�$���|��@ܸ���a��������t�(}�߾��)@~%�^��\R����߿pz��;�=�\R���ҁ��?~�b�	���W��n8q�����Km�s��Wd4��sP1u��!��σO:��]��G"2�.����y�G9l�t�0�Cc4�'���mͻj�KL��s�e[` �s��n9��fȁ���Z�M��]9'A&y�L��B�Y)W\���i�W�����7B<�x�*P;4gnT.�+�S���E��sƏUʘH�Ѱ���R{O^8��)3g�b���V����U5X2��t[��iF��T�u���oܜ��y[�f���kئU���r��f �_?���s)I�����JS��ߵ�B����~��ԥ)�^�n1��l͛2���R�����pz�)N��~��(}�߾��)Jw�{���JR{������ݭ�����k|�)N�׿g�(~�߾��"��y�k�R��}��pz�����D3�u�K]��׹�3?�,L���~��)Jy�}�\R����~��ԥ('~�߳�R�?w�oZ�h7tnu��Y�1b���M�A��bfKR�|���Qn���jVσ�������n)2����K^U)g;r�7/]�xUCRe]�CGc�P<d�<�;����v��9;լݫ5�oz┥'�{���)N�׿g�(~�߾� u)Jw�����3b�����Uv���Vp�A���o�k�ȋ��o�7�q1=��o�a�k#XoXA�U0
v�JP��}w��R�����)JO�{��Y�$�`f/3��ҢB4�*���w�(~�߾��)J^���┊�'�{���)N��\R�����^��TN��[�ug��fg���n%)I�����JS�����?�.C��߿pz��=3�?~�c���[6j���R�����pz��? ���wR�vvu˺��w`weTۻb]_�ߓ����#XT[dEr�l�rF�j�&j3���pp���H�uo����3M���R�j���b����繈����~��ԥ)�}��� Ҕ���ߵg����~�g��l�� Y^�R�>���pz��	�)�?}�\R����߿pz��>�^��P)J{��Yk�[�8M�7ug������q)JO~��=H~8�H�]��K�L�a���UI��C����5�}�8�)C��߾���A����_�2�:F�v��A�c�Z�������N��vvt�+g�R�>Ͻ�\R������v��a�՛�5���JS����)JP��~��ԥ)�}��┥'�{���)O?����a��(�*�u�պ��M���������k���n=q!ΰ��k���]|ݞ]�5ETSQn���jVσ��(Z��)JO���	ԥ)����┤b������TV'K�˺��b�����q����~��ԥ)����┠3��[>���
��i�jh������)JR}��}��R���{�qJ !�?�}���JS�~����(�����r���+���Vp�A�Ij��vvt�+g�݁ݔ-Sn����0�D�����åĄ�1�b�hqrt���h�	���o��=JR��ٙ�c��m��d*���{��~՜3�%_����qJR���~���R���~չ�3b＿1���Ți��y��5�4l�)&9�՜����ł��1��7?{�JYu�\Jһ		���ᘃ1~{���)I�����JS���P�(}�߾��)J]�_�j��Y���foz┥'�{���S����(}�߾��)J}�{���JF/{��ߩ%��u����b������)J���=H������k�Fb_�{ߵg����{���A2Z]���)K�C!���߸=JR���ߵ�)JO��߸=JP~X�.Ʒvvo&�t��4�KE\D���)J}�{���)G��@���p{��?~��)JP���}��R�ñ��wbu.d}�5���9�˅Ǯk>��K��֎����X考GZ4���1���Ø�pO5�	0��!�k2��#�+:� ��� �m	��6�r�F�\(z�Æoyׁ2 ��8ns��1�jǦ�ڛ��f���wd�.Lr�[7�HIKEDEIM15A0q�! )bH!��*(�L$Z����YJI�J
�"JiIJj����)���T4dR w�<Mq��������15	!�DS32D��8�E;�� }���$�&�"�Y3 ش�:�[��
nx-�	���YW6ڃ�Ġ����kj2��(��$f$0��$h
h" ��* �A��0�X��ր��q{�v�)j��'@�!KB�i��7�-�m �6��e�����]#R	�i��Uj��: �o�p�خي��;\>�w��n�n�Jm����4���h�'k]�X1�s���v��,��&�&ɯr��<�n���\j�d���h��6���("r"�x�n�snz>��Q1����QK�n�D�n{+D��%4r�ˮ��:�u
�汲G$�6wU��h�'=[k�u�u
p�Z���[�$�����٢��s<�w�sE����Fƌ�������Ia-��h���Bk�7�m9��I����QETc�ޝWmNvmm5���ўǗW��-����:�y8zs��^��@̙�Pp����g��1�8�Gb�I��f�qɬ�9;Oa�n��K���k\��ma�Xy��=hƸ�1���s���7g�l�:J��䐸��tϭol�q�����MPvR]�h���`,��$շ�3�"c��ͪC�7�d��dʓ^�y'p�z9��
��U��'S��9G-UT=���k��+*҇<n1vUZ���2��\hG7+ɨ]��ƒ��}��c��cG�ÐeӀ�����R	f�!:�g7#v��cG�è�甹Ay\;Pu�m�s��,c;�S�5���^�Ok�_�{|'d����Fv�n�h�ɵp*$��-�G#װ�%�v.n���7����݊Wj3�b��A����T�0R1��m��n����4$�譁	�jP��� {v-�wJ��\���r���̓�B�p3�1ND�4�i�l;l���CRo/
ێnv� Y�\�y,lL�����)[ڙBƚ�f<uN��5Q��c��T�vc�;�^��u�4U  �ȴ�,�u��*��^ed-�3*ɰ��ܫ�sexITz6�-�D����>���z�۷R4��E�ݵ�+R���cJ\�I1�PS��mN�M&�dn}� +�U�HK���j��*�U�V�Mn�1�6�"C���u;G=g��@��X��[ ���c�e��8��y��ֵ��]���O?*w�m� ;;��v!�Y�)��{U��
.���QywC���#lCr�A���\c�ㆺ6�l��X4�W+"S�Fݰ,7j%\�j�,mf������vx��a^m����E�G���5q�͎�%/1��D�p��� �l�<�p������^;��d��٫��s����y�k5�J�/5S�b5�#���D��P-cL(�"�y�������t;��&���@t+A�Ql0�.�^F������!�9�9�e��5�d�i������Umۮ4��E/8�j��ɵ�^���">��Ȯ�v��Tꪄ�nb�������JS����(~�Ͼ�R�����vvm�БEED�=Pf���R���~������>��ԥ)�}��┥'�{���B��=�Z����-�@r��A��g�}����J}�{���?�)"�~����)ݻ�[[��?۩L�ĳU�L�]ƹ�R��}�{���)I�����JS����F�߼��R��y�g�?8dn���f� �A�߽�ڳ�aJ���ÊR�>���pz��>Ͻ�71b]��c��YTTU�'X݃�lf�)�k�g��#��FEMk�ݹg�;5v�پ���6�{�v�N����՜3f/߽�V�R�>���pz��>Ͻ�_��W+߿wf �YG\ļ4�%ESX�ԯ8?2�*L!�"%&c����7(obt �s��7RY�%������!��-M-UEdT�� �j�庳ww�[`}�f��d�W�6�:@�X��ϖ��-V��jW�������˖��Ŧ1�ڧ��v��t��wwߵ+�-S`|�V`�erD���������Z��!]�βv׎퇛���slMl�<+0��w�|���,ee�k~Ա�T�-՜��3���w/� ��[hUM�j�	�O+@�:+gv`>[�0�[X��Ft3����#�z$*H� ����=�v`�H�6;���n��֩e� Q�������r�:�	/8�f,x�/�_��@^]|`
=�l5�gx�J�o6¸%��r�l)�}���@ĳϿzh��7@��gW"Ֆ6��4[����Zp�0�c�'jV�kb����:t&���V���7�ՙ���WCMO+@�� ��� �Ҕ[;; ��c`�YU�T�A!US`/-Y��;ޔ��[䱴_�,����z��-�:lL)�Z{�}�J,�Kgf`�{T��V`~�'�W[d��$���bK��wc`�l�0�s�4<;�0�<
,˅��N�I>��I$���z�������,n�]\��S`s;4;;;v���F�M���mh]���bt��7M�Nĩ7e��Ëtgp���n�kvg����0��;��������8>�����];�v��$}~�`{��,K8��~�y��͹p���Y��>�%6��3;<v�c`�l������:�u�n�~�'Cj�M`y,l��S`��%�� �<���P���<�&������bľ{��?~��s@��"���D��k@;�WTl���t�$*�l�V`��3��{�����n��ߦ��%�X~����c����i��BW� ��X��{-҉u��3���.yd��p��;/k���q�Xh:�nN\�������]���ni�C]�mv�!�-m�;y�C9��[��cP/���*^[�M�u��V�i7&�	�a��q':Q����;����v�RR�V�Nٗi�7o%1�ܷ;f^&#�,e˗��p��NH٧o myȘ�
Ѐ����w{��V����[;x̦i�Wb�\�ѩ�N%}E��(���'k�UV5Wy�i���aM�������/%��z=�mݘ�0�T�ik�l���V�m�w�C@����'�M�>�H������[hUM�t�$4����S`/-Y���}Jl�V�Euw)Ka��.�ڻm`W�������[�h����S`|�6DEP�3PMD�`G���3�3rޮ>cWM���f }�a
hy&*(be�<Nd���vp9�;�]�c#\��/@Gn������/�Zum�I5�N��h�tX��U�}~�`_@:*�Ε[.�լ�\����ߵ� ~�@;C���ww٘��6�+Fs��;C��7U�M4U�UM��.���S`�Tl�!�z��`u_)Bn���DMf ��G��V���Sa�;�I'������*�v�I&���k �%� �]8Iv`G��W� �-/;o�y�7m����*�bp���vcv���C`������������r�V���*n���S`n��>�%6���bJрj&M�*Hj�����7wVg3��C;3�����0G�M���0t���v�:-�m؆��_�X�9�դ#A#J0�J� @4�@�
!�D�HRX ~S���D|��>X�t��{���/�Zt�Ui5�����b�h�=�6�uf;43��;�w�l��Q�����AQ1�`�j� gvgv�n��>�%6-V����J)0����QIT#�n݌nK���Μ�ɍ�=h�0����Y��U�7WPHUT�R��>�%6-K�ٟ ����$�R�ݶ;L)�Z{�}~�mݝ�Z�6����7۫3�������.�斈��&f�jfj�����v6��E�_�Uwt��� 7�Im�UM�t!Ym<��Uz��`wt����\�������j���s�ߺ:��Ѵ�����U�ݳ@����~�6n���z=�l����r�bj ]u+.�W��ؽp[��'g�n�HL�e�m���)	�=k[w*���\��>~�7R��=�6�ۺ� ����Ue��4�ZM`�&֕_��� �wV`G���fvfa���
:d�`�bm]���u��X��7O�_�X�I��z�e�N���Ս5�W⏻�n���E�ot�Z��'U򔭴��0���{�}~�`���2�G�M����1���ۙ�ɹ�����a�b`n�ь�k�����c6�ݱ	�X�^z�{ u�;bG���Bss[�m��A�.ע�ݹ�ܽ:�F�5ce�۩�[T��b%��F�˺�-���غ.7<d�n��W������tk���d��t́G��+Q^��:�:�v'=��\
b���S���v�����a,k�8Pq�ʮ؋�GNH㥘(�+vH���f%��1$�{��~���#�m�v�v�m��]p]6����v(ܽ��\&����G����_��,+ML�UT���c`����uc��yE�����*��N�����{��xvxv`>ݵ������h���&h�x�!� ����.���S`ߍ� ��<��R���E��������Z����h�����vfa��j]�t����A�����h���1j�`�o�U���Y�}T���q��� ��d��Ż]e�G��S�]T��:7F;�om���-�W绞��>]���b'�0j�7۫0�j�w`1j�h�]R;����H���;��w߱�B,%A����4�Z!j�U��b�;��@N&�r����&�1����|�P�m6�A#�ⵓ_M���|`�U[�8	kF�i�i��tSl��@��E�l����Q_���t�x�?�@��Wr��l��i�������F o�U���Y�3��}K���n��MН݉�a��U`�����x�JlZ��j��~qs�o�^��t��b'���n[����p\NȦm���x�ny&w�w{�;:����$5DU`-K� Q�M��R����3|˺�.����T�UA5Y�R����R���Y�����&J�����f������������}�Xtd9֝�9E}�Z�*��57�\6\�a�ي��&`$$��0i1qSy�hsR#k��T��U."Z�Ȫ�����f"��9�C�Ib3M���&Ci�{��a�����'0hŧ�0����<�Qn;�tk6Z
0�}�熍@L�Rf`�3�r7�Ѧ'��14��P2X*�I�zxsv;t3S�3�l�I �S!2���p�9�1�pz���ƀ����� &(�J���	�=S�x���ס;AIP�G��Wf!�@��v�`;PT���J m�����ϻ����s�~�*��Q�H)ҫ��v����x��7@��,{�C@=A+��):n�:H���>��UT��`�2:G�}��*�Rʻt��V�t[is��Ͷ��fj'��j���\�����V��wW��m��ӫ���y�K���m`ԫ���w�.��zb8 ��%$Ӵ�&��k@'H���n�N��U~ ߤ��_��M�v����U���Ù�gf���V�wc`�D�Zv~I�m�
��}��t{���]{��tu]),2$��*��xC�t����m+n��=�	�U�3�f�V� �*�>�՘;�����������ly�un�b��L�x�Gkc�5��]��;�Ǉ�����[�*b&����� �Vۺ���t� �<D��*�wi�v� �%Xn��F�6n�F��j���'�:-����n�/�X���!��x�Wъ�M��WMӴ�C�ݺWt�%�� -J��uf�(��X햒m4�v��7�d4�ߙ��gh���.�BJl��ݝٌĿC��/��V4�[+rbp��y3�mp�vH�Ҿ:@��r�]u����=�k86��b^��Z���8�@��۷=�kv���4&ۢ�,�Ώe����A��%umYFH9Ӎ��o/3Å7n����;�-�k�x黴@-�!��.E6�J��`uz3�y�pj�u���&�yv��H�i	�ڃ�_�懾7C�xꥸ�\�q]q(�K��N�?}���Ğ,X��f%u�r�*��Ե�pZ�{�����B�;;9�Z^i�.	������,J]ݵH�+%�RM�����~��K�,}�!�{�JU�N��"�`���}��UW�$��� I*�vp>�&���"�bj ��� I*�3�m��3�wwU���v`۶�Zuh*��6��o ߻�$� �{��_�$xWx!/Ε[����4I UV��3@$���vC@$��b�bN�&��L�j��fr�F�r��%/8��������ܻ<gZ������l-����n�I#�7��~��H�	���m��ӫ��i�}��o�kА�XN��	(3Phxwy���ݛ=�h�IU�����>�ܫ��I��Zo ߻�րI#��To��$� 6u��պJ��������䉁�{��w&��~� ��S��Ԭ� ��;n��{���<~�M� �G�o�t�gv��z͝h�[�y=��6�<�U�g���m�us�L�ȯ�=sǽk�JږL�p$��Ͻ� J���Ͻ�0n�w-:�bt���7�솀I#�7��$�?~�뻄H)ҫwv��br� I*�3�՘F;�48���������͌�%u`bU�0\%tw�4�6	�x�K�,~�d4
�D�<{�(�+m6��i�/�, �U[���@'tx���>��g�d�v�v�B�����S�v�����#u:��,�i����fR,*�j��k ߽�k@'tx���_��v�����K��f���	i��j� �vg=�Y�/JQ`g۫ ��������E��[o �����H�ffs=�c`�U`}�N�DS�S1U�Mf3C����tXj�����Cs7���K}��߸W�ο�T��J��B*���jX���2�V���Y�K� �+�X/�ۻj�l��$��κ�q۬�t�t6Μ�	�^ۅ:qTgv�nuo��w?|]ኗ�J����$�	�2���7@Q䧙ݙ��]����7t��UT1QT���Y������tot�owc`u[_;�����sL�LMML��CUQY�tot��V�n�k�n��>�ܫ��M����+���궰>���gggxv����.�h�i*I������� ^J������|g�~�*��~��Uqp%E�i����h@�&	�MP��Ip(�15�Ҿ��N��v�b������s}�n~pC���gb�v��g�Mڋ��K�ی�In�e盥q�����z��g�1�ױ�m�p��;v���Ya�|Lgs��yɶ��lP��Ph;�8�ͷv��:�[f���4h�i�G7�S����L��,A���S��=a�U�)dX:u��p���`y��m��c�j{�+�=r���T��toϻ�9�����=��ڈ�y選9�6㞞QM�F�t��;��i��v-��6����]�]�\M@�2EMT�Xܖ`gTX��V��d���ja��a������IM�f >��� ��Z~��s������MLd�[)%z��C@�镀}���$X���"��ҫ�bi���e`{�n��$�Ý�݆��u��&�y���ehv�`{�n������;�eh��������KdP�9%�M�8(���.�-��s�M/���=/�����}�~Vd��[4�h\�`�2wL���������f�=1�TQ3U5-$ַ���>��]v� �Q�|?!�����,�k�If�$��>�b�Ьt��k0�;�e`�t�?���}�6��|` iP���y�"�$���v=�՘В��F �����q,�N�CE7I�{�I�_�}˳��Iu������!@�$�[e�pݸ�6`�ֻu�99<q��ۦ�����Y8��-�xS�W�:�_�N�h�m`$�h�e`��t	~�`=w|EK�WN��In�Y���wM�	��L���U/ɺbt�۬�}����/�I�II?fS!�4$ � e�I$��G�z��Y����꯾��A$���i4�6$�@�����L��;�V��7@���%X햒M;��M�:d4�]�2��t� ����n��/ʕ�Uj�L?cv���κ%�1y㛌�=�Pp�q�T�}��l�:��I��hI]��h�e`���IxΙ��ˤ���-�!���ufs;C����>��� ��m`zK�D�t�[��7m��R^���gwv���[X���5	Y6X�1��Z�ס�f#������\��}�|Q:�1e�C��Q,]���z߾m�?H
����I'4�7u[X���ϩ.���OtX�..�^���i��E��N�v9'��t�J������x��#��Y�wb���554�TU5���Y�|�(�3RX������X�)]��i�Z������)E�����v�c`K����fs��م4R�13QP�1SQ`}�ݍ�}�������{V`����h�i�`�&f����wf�r�kn����^UUU=&ց�)�v~i��� ��t���^�zM����*Η��}�/^���dE��P���5&D�d0"6�Ӵ��ɖB���ѽ�A7w{ު�p��uSG1��u���LD[wi6E�	ai��3uESt'�xv�ä:TC߾�	��̇o��]��5����xF�9��%5���#A��x����Z�{����:mq���B�hI�ԡ�7�L �WX��Az�9:<3�Wnt�R���un�9���h�'�\^g��ی	��ڝ�
�l�rk)g6�B�g9�Kω��ʹ�f�"�L�seE�u�ѹziJ6
.\�l�R�vg�Y"��l�P]vd��u�B��=��{F��W�v�c�����u�4aɢƵe��:�4���d���-�ɉ���m�4�P����'�y��nctl��؆��dԗkX#]P���s��(�$���gv]Tv$��Oiy�\�d����
�t��]������V�u���p ��L��a�;����x�
4��\`|�܇݊��%�;uq�㣑ظ(���95��������;k�8uaFV���1u��gm��[��^۱c�v7%*E���3p99Д��"�k̦+{N�k4�nv��Z�"�8iDݴ6N8{kl��;-]Е���ɻ9��6���)b���F.[7"��#T���ܣ{.�3P�2��ۄ�tʁP����[3؈��C�R��=V&ES=�/I��=m�̬���X�t�6�Y'�';�m�v:��ٕ�z�'9M�q�q�:���ĒոθZ��I����]�����M���u^�qX�6�������g�4=���i�<�&�ԧ8�'�9��d̤����kṈĄ���4�SҡQs܍����:2)*���
����ɠH�]���P�k�U�^rĄ.ic]�ش��L���I�ю<�F�؊���8s�]�q��5;v@�)�M=�0i��m�H�k�qO[.�	��i6[j�[W\iY-�ӵ&Ú��6 4��Q*�O[�M*��2QY]�.������zl���z�Q��d��ggb}��W=�]s��m�[I��dG�� �	@��T=�6�l�誗vZ�s%s�^P�b�(2�H�Xm���m�bBڵt�b�r@(��jz�W���q�َ7��;��:�cq'Fwj�=5�>|�&"�ٴQv��!�b��'�:�@��N�\�=QT�������`����ۍ��o�30t<�k�@f{:�v�-�ۇCٛ[I�[r�0�,��.ٹ���nkM��m���3���h�[;qn��k���s9�C�3�V�t���L!9;�[�����dz6���9	N��^����!�y\��mź��  �4�#:rn^��\�G]v�O<譃j�8�3��\GV��ݎN�"ȼm�&��D�y�'36?;׻��վQ���0��`;U���-�8���jzێnŔN�۵�˗;��#�hʷN�CE7��y ��K�7�L����m�ό�����Q��50�#�'l�� ߽2ӦV���yt��a��7M�R������%���{V`ҔX����3	
U&�M��[������t	�%�����+�N镀N�]ҍ&�BT1��� ^���ϵ,ln�k�{V`���r�ˍ�^f�v�X�ۊ�dN�1��ٶ���vʒ.�|Fv����G��5�`��e�HM;�>�����N镀}�t�yIx�zGW�1XВ����N镈�&Q������{�Y�}��X����g�<����&�z��b��{�����*���mh�#�$���)�5m��)/ ߽&ր{�<��{���+���(��������?U� ��t��R^��B1&Z.�]ڡOk���H�s<0tҋػ;wd���Ǳ��d��Mj@�E�V�I'��� ������wv�f��ܯ� �c�闚�y�&J���=��fs3;�4A�=�`}��� =�W�zDX�I����I=�=�}�r����}usC�#$)1Q(U�"j@�/�C�W�u��W��������n؝��넲��,M{z����>�ڳ ��(��j�4�\e�I	wN }���@X��ޙ�{�K�7��J����uj��#[�a9��mi�_3��9C� ���EՖܼ���i��Tշw��V�m��۠{ҔX��C�36 {�U��6�	��)�5m��)/+�~�}��zG�}�t�q��4ա]t�QU{�р�U`���}����?���i�q<KQ �HUI3�`����V��f�JQ`�ۙ�a�fԙ�	b	"�L����9��l�x���pE I>;3|�����_w׆ 'oL<�Q��i�ﻦ�����C@=����~_����n�F:V�R����\�k�۟iZ�앴���]Ƽ��<���w���\��V�HJ�m��|r���~��h�#�>��7@�+:P6��M�vݴ�����9����7{����v`zR� �'GJ�Rb������@=� ��%�;;�{Ӫ,��`�%2���v�l�o �ޓtyt��d4ߨ��<N9Q*���I�I��N��>�+F }�����`��w1f~~��VC+h���D��%�l�\�LJ�im��˕z�Ԁ0
�v�!=��1�{`	^�O��F4�͸Z.�.� Ѱ�Kx�(9����$�Y�`�nWZ$�2.�4s�`���c�������q)�'�;5pC�rOC���T�� � �E�`�w�ծ��M�*�3�&ҥj���.�@����N�L��ݮ�v�Õ��3�L��fgs����9J�����K�4�����F��3�7"h���nor@�k�u�kN"(h&�j�&���%h���X���vu�:�?=�{����T��&Y$�f }��� ����7etX|��9���<�7t��UUIQ5V��f�.���~������#�;�ȱ+���I��g{>��;�{ �߿]ﾓt���n��۷m�M���d4
���������^'J��H�N���t;!Pv�g�K�L"rkG��B��h�ݤص1�5uHv��V'�hފ�{�f��Tv@{������uD�2�:0-�@��~�:�+��5ZO�TXy+F }�U|��@wp��h��I�I��S����!�{��=�I���mݫ*��i;���N�{��� {WU��y,�=��ox�q!���i$� ��< ��&h��}�� �U�ƭ+�6��A4����3�66����u���]f�3��/æ��Mӻl��{�n�����UV�}�<t���ڶ�D��3SU��i�{��� ywU��zMҿ~���n���N۶�0���}uUߟ}�]�(�$
	���X�O���z����z?� >�9A]R�iRJ���31�����Y�{�H������S��Q5��@UV�� ggv����}�� ��<|��MR;G�l��mG[�{r�Y6-���c�͟v9���vNc��S���4R��'����%h���[;;�0���i;
�j ��i��bh�>�+Fs<@{{������>��/��wvgxm�Lt�D�P6�Ok@=���������X���*�������*&���ݝ���K0����,l;����;�Ì���3;�͏�Y���BxQ5UR'��y�;���@�IcY�3������{���>�I�N�dUbj�V¯��x�n١��/E��C*7jq<��%�����n��V�m۶�m��:mhݪ�|��gw�>ݤX�Q�&Y�����Z����wG�}��t�8`�Ս������ji��*�z���@���5ov`�Xj�F |�U�䨮�c`U������w�� ��b0媬9��5ow�pˮ���	�������V�l��݈�.�V�u�^����W���`�BBB�0�)EB�A������Z�$�U�6�B��S�nm�۩�����x�[�����u�`�C�����ye5%�vq��d�麀�h�p��Mg�9�q�K��d�Z��11�T�5��v��֓��`^c3�2�Tn���P��0��l�-y��1�uӜl�uѧ`���%�3���oj��]���Z�,3S�\�qɝpm�Ce�a�j�Я6iEs�&f,�߿{���ݷ�������:���F�t�l8	ɸ�nޣ/-�7���X��Ў#V�7INT��y�{�X�%��i�}�V6�}A*G�t����x��n�~����,.]��n��j�"��m�V��-=�>�p�>��k@>� ����}����[�۵m��0�鵠wG�wzM�+�� ��_KJ��ݱZ�<�@>� ����}��}'d4Wp�R���*wi�գcg��S!�l�*
�փ[���:s�:ݪyZl�ҿ�Ҷ o ����}��}'d4���IEIWm�V[����o����~��'̅O� �A9��3����W� 5%V���fwvh��GC]U��Q5M`{�_��xw���镀w�q\H����
���� >Z����Y�o�[Xs�{�g�nꇚ���&J���7|�`����Wc`�W� |�U����O��������rru�
6�͕l�[3�q��d�bv�3��5��6&Ş%�&�������F |�W3��[ݘ��9�ꩢ�j�**�ji�y%��t� ����{�2��tIU!ڻj���<� ��<ޒn�U[Ew� ��CT!h� a�`���FhgXXX6F @8K$`�`HaRĬ�C���2��3,hr��1��#�0�R�(�0
�&:/��̋R{1�<S럯��[[ﳇk�NC�Fa��8�U��N�Dadc0U�$%TY4��1F	���"C�"��
Hb�`���Kf`m4(�[c�����[D��μ!�a�sg]���L�I�-ƶ����Y�������X���8����i��ƴ�
Q�R�j��bM� ����{:�s\Tό� �RV:6�N��nxF�Ӡ[F�0�i��"��w�"z�z�`uc�@�]G%�	�8қI6t�t�$����F,�#��:00�)ě3,3+*���A�nޛ�VafDDa`F6�f6����0)r����s5(j���%�Ӡc�� ���`���] �	ڪtiC�P�L}DC� N�E=8��h'gR\K�(�qa���uh�~���))�aꉊ�j�Ø����uu���I6��H�����v�AcE*sU5������w����ouX�Kt�ĳ�Ab$6І�WmSt��v�;"�;n�v�ՊѸkn�\���0��4���`�t���#�7�M�=�2��.+��X[��=� ����gw�>�wf�u���{V6�]�M���x�$���+ ���k@>���~���L�*�V�Zy�3{u[Xo�� >Ԫ�30�0(D�	(��3�*v�����>�O�$�����_U2�����h��*�>�%��U�����ϟ}��g��	�6l��PR*1:�L�y���L^\�;"���9��̩��Q���6��+��`������>F�M���,�<�[XI�u+�)���t&$]�k ����;��k�рly)�vvh��47sDM8AR4�L��`˭����߃��,��7@�t*�nՔ	�QT�䳌F�M��jY�3;��&V���2���v�In��+~Գ ����>[���z�K3�F-�������ne��y���k����w��:�'n#N5�K��Ei��3Y)����WU��lA�\5G�:�D$RU{n��8�]�c���T\��ہ�d{=���9��H���q��m�v}��λ+���*>x�Q/7�ñv`6��!=��䶻*{\mڻ<Xd-Ѱ�x�ݼMY����<5N�s�-�0�q��Q�6��8���n"�\-�߿{�{����s�������NGrl�gqq]\�QHC�^x��Ƙ��gk3���u;�U���l��X��tzKk�h�g�67�lI��DEQEժ�BOtzL��N�h�H�w���wwf�wwh��UMSQ3UTT�X\�����vh����w���;���I���(��33��"�=ޓtzL��;!�IJ�JMI���m�4w߿s�$�3>��ڴ�vC@�� �^�$�;�-S��2�������4p��=�ps�ݴZ���,�P����\]��uv�Yo�Ot	�2��vC Q䧙��ywf �\5�D�,��j�;����ظ�b,?f�1:$1��1����1(�jM!�&�4&��hz/�gff�ыf��Z� [�����
a7L�e4��I-�@���N���ߪ�ӦV�d4����&���56����`�����`��� �߻�+�!�]Z�T[{�}�2�w�og������0��lCH�M�c�v�Ǥ;v�v��B��Emzu�[r���ь��\z#�긊aj�n�m�~�����=�6�-X�}䭬��3-HhLT���a�z��`}:n���Š{�{�A��?O�Y&J��A�lں��~못�߸rW� C�- �$�$D-�k=ן}��_g�}�A�y5��ܨ,U�/8%���Š/$���j�vwgf�K��p��5c�	�t�u�OI6���Qt�X%ݘ��k���x㨙j��&h��hztu��/��������wl��6|]��fN/ֲ|�WXϥ
�����������t	�X�鵠PJ���ۻ`؋i�w��{�V=:mh=�o����T��$��`���	�&ց/���n�w�T�۱��i6�Ӭ�:mh��`��t��o���~���a�l�.�Xc��M2j4ڇrė12�C��fF&҅���I� ����c���o���2�%I4L�$�U� �ڦ���Y�}�X� �~�����������1��F������rg.B뎃f�GM��M#�3��3�|ܒU? �/߳ ��H�7�,o����WM����A4�I-U55���E��Ic`G�M��f&f�9�TIH4L�12�������@}����k�0	�+��,_�Wm����>�tX�t����k@=A��M������'t��}�p�'��Z��~�SJ�F$����]m��-mu�v�ݔ��7�=k"���e#��n7l��;�y�#��q��c�p����E;�t8ͽ9׶B�g^x��<&���ӧv���G�:�r�N�s�L�q̮���X�H��j��<�H3��/�:YX7f0��۞vJN�Ӹ�u��Qйe5N}� i�J��\3�ј��M�T�]�*Ă�ϓ�v�Y^�{�{���l�yn@����UM��&�s��N㴻ӹ�.�ե��۷t��uj�
����R^=$��=~�N�t�r6�ci�M�i��;�M��� ��7@��K�x��]3,�T�TLLL��[`��<�,â=������54�ʒ�%�b�f����wfgx�]�`��}�mh����J�b��t�����)/ �t�Z�txӤ���g�է99:�Z������F��K�܈<^K�v�yܮ�D��T�����n�L�Wm���6�����I��R^<u�q�wt�4��m����G����6�;�;C3�{f�e}��}�J,����~B5�Zc�v�x�$��$��wvgh�K� 7WU���!ECH�.�U��{�}�%�{�6�������\�S�n�6ݫm�M���� =�U`g�,�>��3�2����;��p�xmmlf�n
l%������n��v��z�J�鶯��t�&V"j����`g�,�>����X�JWщ��'J�J˶��I7@��K�=�t��{��=�r�@O�Yn�QSU�ޔ����V6	ݞ lgd��G�c ��`����H����l�'ׅ,���� 0�C��S���f��mՁڹf��S4T�S@UP�UE�;4o������`{�V`yIx|z�\n��*��6ݧ���G��N��}�%��I���\��C��c+��|/K1ng$%yy�E/8�Dmn�q�[��ɸh_mZ�#kj�MX�՘ޔ����,f| ��U��f��4�2CD�MT�f��(�g�7�ݍ��������fff�:9G5!$��I5T�E����l ��U�;3��-��}�%��:D�Rv��+��V�{ڪ�����>�������p�
��;"����:��g�n�����[IYv��>���R^�M� ��<p%ۺm�+�,�6V�ݍu=��͓���qԛ���:�J%�	ֈ"{2�?�e�Tƛ��)/ ��&ր{�W��}��t��hc�6�n�}�mh���zt��)/?P���q�YJ�hM����{��>���R^�M� ���Q/�'lT�SU`}�0�)E��V6<F��{�_ҿ��Ch��V�I�����{�Ս����3�V`��Q�t8�پ �bVc���@U�/�Q�7�]X���=�o-1p��%<rI崌V)&��(1qB���\�8X�v�]Q�Rm5�_��r����ż�N����.k|)m���h�G%M@Fhu+dk9��Mބk{���9�V&U��d��FS�QȄ�]�L��0�hr5r:#�ӑdk�"%��-�8p__n�Sh*u�99x����4 ����1�)&xi��2Ӿi�f"��[�LEϾ��'��s�"�.�IO�������6�����l������4%�-��}+��:�3f��kzr�l,8�΅��YOp �_چ������0.Y�'�#�>�ǵ�EX��f�dcd��a�gY�wJb��J��0�8גd�J��Ֆ��Ɉ�dJ��H�����aE�a��Jӹ�I�tp(iGp>�e�a:�6��ît����� Ml`���a�l^���`!]cse�[d���:�Mt�]q�� v�A�wj���s��^A0px�d�
St<tp���Slt��s�� Av�ȹ�܉:���'<Wm�7'Em�Z�8;v�63�1q�H=ɷ��']�4m��j���c\���X:a����,rq�d����=�N�e}������]N8Χ��]�����z	ax�m�����!�H��͇�`���/.�u�,����J�l�#U����]���UHb�f��ܪ��2ve�A�{3p�*:f��*/ Ӫɩk"��8��8���g��
K���y{�Ŷs������=nc=;J�71[�錛q�\X�6ӹ\,	kn�����K��N�P`����nݵ��m�v����槀ݝ�jV�c�� �h��n�<��^��t���xZ^s�J�����^��ێ�']���;��Q�Q݀�`z8����U֎{;fx��ێ9aZ��8C��t+��i\eQCt#�Y��]��Է�c�k�,ٰN.����T䫈�y�a�Ћ/-v�s�c��/kg �=u�q�X�Ͳ=uԪ�Z�v��Pi��0��[�z���<V���@�^F�!6�Ƶ�qŐ�rshw#e��f\�{H�ulH��ъ�XR6�g�=�{F�v�p%UlcS���T�N0�������.�@kt�#ѵȰ�^/�R�Y���X�`:��0�,�i��چ����..�#wl8ὲ��cH���<�>s�cb�L(�c�sd��bCv��p.�<����Q��㝊7d�ѳ<�e�Z���U̫�-����.����*�]U�����`�uX�M.֚�i蹪�u/at�*�D���wH�G$Yɺxx�����-����fƒFv	]ٝ�q�S��`��y��4lpv,�=�n7:��j�����NR�'Ev+-
�����E�t�����H햻9��̻qC���gV��8"p<��B+�)ڋ载��G�l:v/����(�M
�d���A�
p�^�N��t���Z��Y�<m� G=61\ƕ�K�ѝ`^�ݬ��ՌFz�v���9)�l�s��Ŧh�R�⵷�w4qӨ�����l�����h�R���l����՝��m���!Cq�[m�M��S����,��v8su֎��L�ӑ��;lzva��mq�D�:���������6]�c�:'k=��[�[�\�@�JGjU�E�*�'=[l]�]��w������<jz��ϭ'A�	���"�td��%iV�N����u�:a�E֝��8�MQ��uc`����՟�}���'��J�;IJ�yZ�tx�t��)/ ��&ց�����vҥe�o �Ӧ�yIx��6�����\�!v���*cM�����{�K =�U`��Z� �J��RPK��T1Q`{�K �vh�]X��fߧ��@�Ļ����m4D:Z(�܂� sN�kZ��{r�ݽF(S�+��ǲ96�V�}���^4��Unզ�I�|�?���M�>�������K���rn�y����՛��ʺ��~�=��iOT| ;@P�u�z��r������߷��UN���Eժ��Ot����wM� ��<}:n�w��l�v��4����mh�����t
��K��WH��NժhV���{�X����=�`{�Ս�kn��(�g8[��5c�6zyG,����(v;]����6����wU�Ջ�S�]�9ag�3�V`)J,}�cs3?�
�7���?���*ƅLi��>�K�=�I��u�E�}��tp��cC�n����=����ln���w|P����
�� `tX&J�.Aqt����n}7t����=|�4���-�LMc`s;B��l�]��R�a�{���9ɺe����
j�"�lԦ�E%��2_tX�%r���uu�s�vɋ�[Q��l��R�\3���G��ڸ�����q��qݝ�&���덞��R^�!�u�E�{����ʀ�6ݫm�M��!��UU_�]��5wv`)J-��1�ڔ̳MD��LLL�Mـln��=�,Ù��#�=�xI��Ɓҕ�ch�n��T����>Ԗ`)J,n�F�v�ٝ�6���,ĳ/ӻɠ~����v��aot���wL�����I7M��~�{�nS�9$��]��=4q�ӹ��]���^h�̘�;����xP�ʴ]a��6���x�L�����n��R^��v��5Cn��4��� ����=���U� ���i*�Z�����If��gh�K��\�� �����!�]Z�M��C��=��������Ú<��� ݎ��M�nմƛ���!�u�E�}�M�>�K�5��S�8;�*���^n���[��ګ53������\��`z�V:Wq�9=dYC��ˍh����q��W�Mm�ű�q�m���u�7L3^��&�;���D��{Y��P��#�	٠�܏7n�m��ʤ,�{D�svβ�]��盍���i��[��ee��ۗ	]Krv��D��wg�qS�ػr�,��[�"o*8moL͛�.SS%���)m��,I5�i�9�q@����r�v�����燧f�gr�[��.�|R֍+�mGO�}��+(��oͶ�����>�&�E%���+�����;iR����I7@�)/ �t�`���%���EPI-EMV`��۪р����RY�{I*�I����`[w�{��hwG�{���}��wǯ���~*�6�����n��R^�!�;������~��&ɋƉX���nM����i�Bsi0v֏ϱ���Խ����VZ�"��]ݘ�R�ڕ� ;�<�⤨�!�]Z�M��@�)3��`(�D#5��B��
zA=AP���>4t� �I7@=�6m�V�n�t� ���t�t���k��$�����j�v� �����t����L����;h����CI���n��R^���� �Wq���6*T��T��9��ᵄ����yέ���.�G9b��n0�E��a�m���t����褼�L��wtxN�tq&
�I����v���Z3�� ]V�ݘ�R�|zࣷV/�[ݵ�hwG�t�:���~��;�5>���L@E$M(��A-(�"~=\�{����ʾ��� ���J��Ҧ��xI&�E%�:d4���>���Ch��V���@�)/ ��!��Ӥ����ի�PX�m�*:��l7m�]\��f��n��z���$�����h�i[�4��:d4���:t��}���$I~N�&��m�� ����L�>�K�;��{�~�cG��m]+M�I7@�)/ �&C@;�<�=�T.Ӡ��Si7�����w_���1��3z�eř33�??ۼ�x��),��-�m��� ����M�>�"�?�$��5�I,����Q��:�ԏ���8���OG�ۛ��;\�ݸ��K��h��@[����$�� �$��.vf|�\�����L��L��!�Ӥ��,�9/@;�<��RTc�.�U�m=�>�"�:s�����:t�����6�Cm�n��m�9�z���:M��� 7�}-_�4�hm�<���,�I����9�z�W]�#�N�ٗB���K��n�Věs����g�9�"��u�+����0�+���du[�s!)Ӻ����E��h�(�)��n;i;)�8l�v��$�Gq�v�rp��ʭ]����ǳJ�4Vv㗇�ƶP��3�u�a�a
\
�ۡ�t�U�QG�����["d�Gkו�,�k��A���<Lʃ1��h�ঐzQcj(�[�7@�)����eK��/�E�9W82��tn�o��)͑���h]���9P��:���gщ1$���`��E�HZt���0�%6����ff�B]6T����]�PYn�6�{�}rE�t�%����:M�:
JBjڲ�M�ET���� ��U����wf����O��(ӫv�۽ǋ@=� ��n���E�t]"�
��ЍR��T�m7�t�7@���,���{������-U��;VѠˍ؋�nGr��PC�:��mۀ:����qs�T��6��Ui[Ot��,���{�Ӥ� �\��݈M�V���ʽ�^����*|0�ȐL�#�	րLY��C�����fi�����0��M�D
�������Ֆ�OŠ���=�t��,��E�tE�N��&�ةYUV���<.�ـz7�lS�S��G�{��r��2�ƅM�Ot��M��wT����^K0wfor�-�ɻy�&ٳ��n���J�<�x�e��u��nu��Y��><�{={�]�:�,�S`.��p��V�%�������iՋ�c��z��{�;�f�y)��j���<�S#U0CKEEMU���f�y'�?����h?$?մ)_��&�]tƈ$1��8!��Xc���t�.�rxhB��p�Vu���24oi��#A�FیGFh��`g�L9��i
%�q;QdN
88� x��`o4�&�ʌ'f�f+�:֫M��:bF9;|���^t��I0��}Ax*u�`���O T0�.,�=�C�z| �!SbJ���i����0D8_�?��wG�}ꮄc�.�U��{�}~�`���{�UQ;�7@;�'�bN�v�m�}�%������f�y)�?37ڛ���y�Nt�V9L<&6��<5e-ɱ��K���QmONq�*VM��,y�Ck%����۫��_{V`G��wv�g��j�0t�0K�TE�RMMU���Y�������U�Z�����4D�B�e��_�XN鵠���f�N���j�h&��"*�Ý�r���yuX�,��g������q�p9�5�itJA
�.�B�����"����)���Zji����l ��V32����(��5n�. }����#���n�T�s֤��^��X�ٻkuێ����71�ڳ.悮�[���:zM�:�"�:t�Z����W���!�WJ�E��@��S|��.]�����Z�g;;��D��Ʃ����"�(����wc`������;�v`
7�lQ���y)���Le�̽ ���	:M�:�"�$�6����v/ͻ�i�wm7�I�f���Kuc`���5��5���C�Ѡ4xmRY�(b& 2 ʹ�# {�on��㸷f��M!�n��h4<IZNֵ��F7eG��w��O=�9�u�n�QڠS&h�;1ӻ9��[k�F�m@��LG�^]�5p�S�n����z��j����`q��08؉��vb�C ��&�&N���Jv]��r��R
}n@V�;�/ss��z���]j�����e������j��=��1Ş��}-T+�L؎�0B�M�?�{�ؿb[�.��lr�Z��|�=����Ԩ�����*��N�A��۶��c�ӟ OO�I�Z���{����J`���M;��m�zM� �����ޑ���J$��V[�i�� ������zG�n�,l �<�Q/R-UV����˾���`{|�媬�v���Z.�;I�w�x�ݐ�N� ��n�������:n��gv�q�bE�G�ce斑ne��Yy�,�a�T7;���uj�e��XN� ��V�K9�پ�Q��`��TC4�Y����k\��W�{������_��M�>�H��d4�2� _����������7ږ`Jl�gvh�r�� 7�U��M
	j����"�k09���N�M���0�UX��`�:R�6¬M;��m�I2����&�zG�}�R���Ӿx\���f#Vu��v{.7!Dݽ]�u�����s������4�N�_��ն�{��ztx�R� �%\����]|`���OD�H44�TMUX��g3;;�@-�����媯�����>���J��&I���ot�$�6�����EH�̰UQLţ�̊/���hgvv|?O������� [
S�SMTD�D�M��fx�wẁ˪��j[�u�E���ѥT�۶�ݤ�ӣ�;�M�:�"�>�M����߾�f�ܹ�ڹ8��S�m��%p(r=y]k����.X\'[���NϛE����t�H���k@=:<�y�G�ED7!j��y������ě=�ݍ�˪��jY����o���������"*���.�l ��V�R� �H�x$J$��V5Bm4�և;;Do.�j��c�M���̙�ٜ�f��B<M0iLM����i�B���`�68�68�qTY���Ϊ�(=�
%�A����j���jY�s�)���=˯� ��V��QEP�#��#�.ۣf;$���vnw���tp\�Nì\�wH��۴Sh�V{�u�E�}:d4ӣ�;�&��~)�V���i��}:d4ӣ�;�&�~�`�]UI�ݻmݥ�h�G�o�,Ùٞ!F�M��]|`jj��Mݱ7j���I�_�XӦC���#yuX�G1�K�DD�A55�ǒ���˳��7�U��Գ ���/̎$�~3+�e�����X�6�ඇˌ�D�n����G�X�kk�\��݅Pg��Ȳ��t���3���9�s��
��!0�ض���6���_I���W�=Z�;2!mh�%��)le�y͓�#JS��1�1�.vL�<e���H���(l�q����se��rR�t��6D��reI*��Y1���5����8�R�k���4!�eI`�3�M���P��[��>�Pmպ���eU��OB�����{\t�3[�ms[q�����m���?_� <�U��Գ�;���
7�lӣ��h&�i����� =�U|����ݘ�{���n�l o���
%�B��[���;�t��,��6�����+�\n�M��X I���E�};�ր{���7@$���ui�h��XӺmh���ޓt��,﹈��I]�wk�LM�6ܝ�����e��xv��k��z������!'O��vbJ�:�m���V�{���7@��"�߀�N�Z��Wb���j�J�&����Y�aٝ��hvw��=����р���fvx��ls�DMTSY�z7�l��у;�j�~�[�t%1�l*��˶���d4��V�����=;�6ӣ��kX�	����tx}�7@��"�;��o�,I}���G�8�.J�.E�9S��M��xS8��x�0{DxV{ .2�F��eL����Lj']������8_ߢ�>��W�tLx�q�E6�B�B��@�������� ��x}�7ww(���4�5RA$MT�-�GU^y�����#��f������_�X=GT�]Rt7n�wv� ��U��� �<��s33���ݍ�yqPt��DT�T�DMU��$� �h��V������U��o!Ląof�gn�ۥ�nu��.^ܹN�HZ���������n0]�>�mp3~~m�����}/@>�G�{�&�
�e�%���n��߯�>�1߽���%���U�;D�;�zjH%��a6'�/@=����I���<ޝ8� �����9� j'l��f$����f }�U`o�X���3���;;3��,�������fU���6TH�RB����� �I6��tx�?~� ��?)?"���q�:�mJnݱ[dӧNZ�[t�����	���&��+��u�i�he���I6��tx�$��fv���ѫ��;A7uL3M1EQM��������I���<ޒmhtu-_���v����I7@���`UUQ�I6��tx�K�K�E����4�@>�G�{�M� ���I7@���wN�
Bm�wm���c`��V�R�����1��u���L��$!lq3xr�8��ړbsgʫ�K�N:���,x!*~�#)*C�\Fm�8u)�s37����G�V��/�5j��g��A�<8XDFc��g7�`jD��$�c��:��Ż`^c��ʥ�7�d���K�0bѡ�CQ��]2�N���	�q�)�i\M����A��N���5�4���`�ag&�z#5�k ��oeG���� 1'֭N�����ΉMi��a���l���Vh�4�R���.�}�$�pR���3T�P�L�%F0jCGPx��5� �^s ��ŶE�xFP�0ü�&�:���Y��DTt'��aA����2�GVa�3�v�9����S����	I��A��[`���XV�NT\���1�QmJs�G	û|Y�w��'���� m���m�6�!�m��I���K@m�[z����˜S�/n�6�Dcg\T1��T�u1�k��"ll�+�<C[�Oh�Yê�y���0ɞ�r1ʜ��۳�T�6�a�ؠ5���Wa	)�:�ZNF�m�b.�km�iN�s����ɥ;^E�ʏ�g�NM6��㍠���nCcF$\��j�+�Sn�����\^�*��m�k�W�*�Ӷ��c�ř}	��ڡ�-�N6�fps�2M1��iڹ�ez�۞7n]��_YǍ�n�]���ԑ��ͳȖL�Isͱ�ƌln�i���M�{)ۮt�tgukBAm�+�wZP�n��X�=A�d�b�r�j����rY���8g^�>:��'aݞj�ۜOJ	Z�&�<�	��T^�a�*��6�6�g����i�K9-�ǭJS��r{J2���s$��I��N�n;F���t�<v�3�s�-�Jw:Q�`���۬� e�5Қ�Ŗz�n�gBmU�:��f� W\� 8s�l�J�%�]Q���6��W[Kf�h]��W����V�nQ��$ҫ��M��5���.\!��b�z�h跳�����U݅��lz݄����\.��Ǯ����rmֻ<���X��Tp������Hu`��7u@쑀!"�
�S׉.ѡ�T�u!.u�V�8����
HNғ���nJs�(U��k9���[AI���N-�Fp�P%.յ3��Nwkm��d��Cc���kbDw�B��z���c.]��MX�K��nr��']�DK+�9ݫ��K��7Bv�8[u��\�[:�r�-WCbStʛl��P��.ɩR���I��2�{���]�d_�O[�˔�bn+1v����2�l������;S�ی�{Ni�k���L��ls����r�N2���{�&�*�.�<PM�h�8>�q�۲v�m��UU�l�UT���+36�:4q1��y�nS�uml���8�M����k8�N�N.
R/�n�{���D��p��M|���@m'h|!�'�b��(�T8#�<��9��y��5�XVk�������m��#abk<'T\������3��7�q	��+���e���n�9�K������?=!=�֧�F���@]m�ݐ�un3l8(

��rd����C��eS@�"��&��0]�=qЎ���N���n;lf痻{3����d5�]!ɜq�i�5�%bS��Ĭm������ζ�Au��s�X*S��=T��?]�n��ݗ�ȲO�a��VN��a�=$:�<un�;����θx��K7�,�ѵ͕A�V"[-�W ?���t�t����mh}@N���:_��[i7�wt��}~���k@>��]�$,L:�x���H[�	/8�+���jX�s������`-]ـ/�:um�m��w�}:M� ��<��n���}˥�\��D��:)�4��<� ����n���K�>�3��>���{�;P�$�����^SqGJ��n|(�����n9�����a�<��v��ށ:n���K�>�2��<�GJR���e�:�M=�>����E@ �OG��ek\����U��Գ9��㩺���I��*���.�l �ڪ��Գ �˥�uZ��$�Li���?�_����%ݘޝQa������ �&��zixih����7u,�>���I���G�}ި��� j��m�m{(m���c��r�C�s��=�v�k�tl�"�m�Ch�H�+Ot����$��{Us3�@$�� ;�sS4�53SQE5Q`|�,l�vf���`-]ـ}�J/�� �t�LC4�UMMDDն n��}�fϰ�;�C��:w�a���!N�\��k��ʺ��ߺ:��QH�$����������vr���=���vр���<���1�E4ET�`zR��ڳ��7WU��yM�>�v5.۱�?ZNڧJ��C)՛�����n���='94K�i�Y��=��^����v�xӻ!��G�w�&�yIx�Iq�i�'M;{��{ڪ���ݘ�{���-�`|�.���:_��[���;�&�yIx}'d4����ǎ��!�]Z�@��x��tXӽӀ����f�g�f�������k >��jb��*�j�$�f����h���<t�t�������A�"�Q:��(@U*#��� c������;�5ˁ��ҥd��|m�F�&�Š�G�OI7@��K�'s��D�5�TEL�DDUU�����wf�;Uq`rU� �����m�*�� �������G�M��i(Ý��ݢ��`v�v`�V�T��Q54A)�wL��Otx�&���`x��L*�WC����� ~��R�G�M���Fm�[3��0�f�b�]�h�=9��$��:Q7s�v������ِ���	7�{p��:�w�Mq�ln�3L>�לu�Ru��B���/6�ԙ���lS/F�s[��F�ŰWбw.x�z��6:��뭫��n�]	FM�70��<`q�����x�w�B�t[e!�N�^�ltO;������;�+���i;`9jă�1����[���nf�b35�$օ�.�qg��ɝsZ�:�<�vW<sc�g\ku�tX�ɍά��f�\�爚� r[ـ(���Z��{UX6���HB�6DB9y�??��o�K0�\�� �]VKVg;4@wB�*j
����*�j����] ����V`��`Y*K���v6���fe�����Y�(Z�Ù��f�S˧ ��4Θ�6�v�wv��'N��tx�:- ���'�Ki;���U�[�Gj<�=��.G�H������q�ump��ֈ�vӺ�i;uv�{�tx�:- ���$�7@�F��-~�m��EUUX	J�9���]���������%ƘU���t�-o�%����a���r�:=�Հ�GJ�k���U�i�
�D��7@$��{U`Z��|�M��D�UHCKDMf w.��t�WW�˪���{�8��s�%�L��E��'���Ǝ:�-��"�k��,���/Xy�cM�K����n�x���I��Ӧs�;0�� w.��s.��J��j)�-�= ���'N��tx�����D�L�Ͳݤ]ݶ�	Ӧ��{��i��w�1�,���hJ��z"���<������uUܕX��C�5�SY�3;�-S`-��pV���wwx�˾���H��ݶ&X�m`���G�I:n�t����.YWJ�m6�4SO6Z.+�`�^}�v��9�n|�Y2���:��Į���(&9�ʭ�n� {��]%�0��y����t`p0�%�ᥢ����Ij��ggg�r�;��^�t���$�1mҡOpV��T�`��U`$��B6SMAUTUEASUa�������� �uX	$�;���������Z�O<l�����Ӷ�,yz ���If %���%83{���@4n9S��h�ݞ�9�\�����[�%���a�(�;ֵ���|�X�X��U`wwv`�TX	N�8�UX����i;uv�{�t]/ ��E��U���fs�4@�]sU-2�QTKTD�UE��+�pV���Y�j�W�}�BGt�Yj�i�ks1hN� [�f�uE�;;�mwt�p0��K�ҫv�x�t	K�'��iW�{��WD.�)H���IR		S�qY	Hy{�?x�.ؓ���n�9���V2�18��M$��7^�]qL�^e���&6 	v#���5���݌&�l��Wg]-fǚ�a1n���miі|�(����v���?+z�Y�� #�g�7l���D���P����"�@���zz�U�r�8-�k�=[��n}n`��6�P�]t덤�䲢Wn�=�Aau�趔�8E,cu��8�b�Ė/�%�K�ί�i��	I0a��T����cgM�Zųr�2�!nN�s��Ψ��':�Z
�����׀N]"�	:<zI��r�;�ݷm�;�')$��vh��]V.��)���}
�*_��m+H1<Z'G�N�n�"�x�$Z�Q\�L�Ͳݤ]ݷVI,��Q`%))����`-e'=52DLUf �� vd�dZ'G�I�n�u��lt��E�9�K+��v��v;u���n�\���Y\�u��N�	�Pn��Bd��I��o�� ��<����{� ��q��
�4e�ٽu��]U}��o�_UB!eڧB�
`!��;����`-�Js���2�8��)婢�����.���Q`o�R� KUX�%eX�`�Ю�{�H�^���	:<�$�\9J��v��ĝ�����s�>�&�.���q���xx ��T�m����.͹�-[V���Eq�65pl���~o�x�-���Y��I���&�~����>��t����cHWv��=�M�:��`9���N��JX?���i���6=�l[ZY�g�G���a����jۖ&INbѠ�Vf8b5�B�!@Pm���_�]pC�o���՚D&5�'�N㳡��uMk�A�	�\�A���]���)���7<��Dcc��AG �"���̰�2"��(�FH��
���<[�����-�Z���a�YXƴ� �(��8zm����H�#����:��+��>��5.��EIu��6��JFM���\U�=��QA�8I��A!�ǁ�=���	���f���e��p���փ�ir��2Σ��p��
��� < ��[G�w�������g�"�|�j��)���Ţ�0lN��E󲎃	#�,��\HӬ9�C���9���"��<�Ԣ�OQk13��]�tu22U�H��o0�0��.ss�<{���;SO��,A8�呭���E�P#�`�`�z*���zDM��E��Qv hUé�H�)��5:P=�����x��g���U߾}�]U���;N��LlLJ�&���� }��yjY��3�;�B�����*�h&J��6ֳ@'txS�L�%�E�}�_���=Z�1��G\��R�x���Z.�.$=��6�'��ð�e����N����:��o ��n�/�,����S� �UX7�� 
��Z�����G������7�ڰ�Y��(�O�n�۶���k ���<��M�%�E�u��:*��t4Ӷ��� [����`
<��s?�gf����i4;�'x��K�lWm #ǀ��λ�ʼ�^�>�'w��v�E�m���M�*_�Xt�b�7�ڰ9���I3S4ISP�	{��:�����^����ծJZ̴q˴vzL�"hqJ�eIbm�@�~����>ذ���ݲ�Wfܨ��!�&������7����3�D�U`wj��%�E�w�u�cvU�mӻ՗��<Ot�_�X|�׀�]ˮ��U<�4ML�Xs4wj���6}��Q��<�����S����y)�3g���Հ�ڳ ��n����&H؄�RB��%I�N��.gx�l��#�p@��ٓ�cv����:ݪI��6q�٤�{s�q�7g����	5��3���&c��ҹ���{Ғ$Ӛ[</c����{+`̔�ݎ�m��nm؉,���s��ޑ��\l7k �lv�aC u���*�Hݒ��6����@�gb�ݸ�u���nYG=����lP�U �K�z1�����ww��p�ŗ;<-����m�+c��$�ƴt@l7l;7���m[���)6�uv���^ w�� �	K� ��<tUuV�n�V�2�wJ�/j�G��~�l_�gx��ؔUD=STT̑UU�ݫ� Q��ߧ�x��<J'R�
��MQbOt	~�`��^ w���=�t	9�J6?�lT�V�k ���x���H��]_Jv���Ӷ���m�$ctu ��fή�S��z����sq���m��q@���.ۧw�/@'tx������@�g�z �����ʭȪr�o*��=����$Ć0d�s�Q]�!�<W�7w�u��7�� �{��C��2�i;T躻Ot	~�`��^ w�� ��7@�r�;��nڷWm��^�����{�����}e{����wm'M�Y�zޑ��=�4Np�;���������߆���%D����Ia;�&⎕�;P����q��U$<�=��UD=T�13$�U��.����,�{� =�s�$�}JX7ERI�,I���|�׀���{��s��l�ة���3 ��w<2��`&v*'ȩ�L �]�[\X�Ch���H"`����Yzޑ�{����w��x^sލ����yjh�������9��{�@�]/ ;��}�X�P�P�ݖ��6�Wk-�c�^z�1u��\�ٮݳ�i�v�쁘����,��N����@���/u�{��	=�t�B�:wm��V��w��x��<Ot�_�Y@u���WV춚V�2�wG�I�<�^��6Ͻͦ_�Ӵ$�e��	=�tzG�w��x���D)@���J9*=�f+�1f/%��~��>������)%�A3Y�(�S`r�j� [��^՘�f%��͛�Ym�	��VT�n���k�a�4<����kG6Dˣ�9�պz����Į�7z��x��<�{��~�o�;g�,y29����&�i���� [����0�J,�}�|��� �Ĕ�K�M<�4ML�Xڻ0�J,��Ws˥�� ����Te�I'j��Y�j�E��O�,����]�/����CL��&նZf�/u���V^՘��X�ݍa�h�v�"�Lp��Y�k{����Fk��Pf�n���v�f�;=�VI�m�g��A�!��n�]��z��=�Վų�TR8N`�K�^����9{��]�ۈ�j�L�ɝ������2Pv1k�SJx��0��6���ƈ�Ѯxl��Fv�u�"J^��F����\\s����)��G�v7�����5�p5i�^X�<K�Ƭ��q6l�}v9�R���pn$����ffb�b�ŜIf+�uvdM�B�i��cCh㙸G:��ב��K��o9k�a�+P��7_|v�v[v�k3/@'� ��7@�R_�m���x���m1~MZHV[o ��Y�(�S`o�� �{jـI�k̫l���TX��_�X|�ׇ�~��wG�t��EE�M?�hLV����;�� �{�'�n�/�,ﺺXۤYj�n�����	�'�n�<���^��?�Ү%-]������Sӛ�c�2�!��δX�N��u�+8�g�s���L4�IO-MS5Xv���)=ݟy��}�w���4(�]���k[못�_}�y����p��N"oJa.�T6�]Y��9U��{��=�t�B�:e�i6���x|�׀���{���K�:�ʝ
*�ݶ�M%����<Ot��z�>��9����s%��HF;n�'�n����/u���x��r�Lo�X��1�K��cJ;�*.�v��5�غ0\!.ƴA�y�����c-����,�^��{��	=�t	\���Ƅ�i�X|�׀���{��\�`{�W,m�,�Ct��V^�{�o�}����W�'bG���n���˥�{����~h�:��o Kڳ >IU��O�,9�#wUX�����J��:*В{�I�/u���/j�����:a�Zf�&`��I��=�����\th��[���%pÔz�Ψ��ҹђ�cU�|I>�f��/�C��<�{���G�u��:U��N���f�� 7uU�Dڻ0��V��׀}x��U&�hI+��x�������^ {��IR��(l����"	��fgf��wU��:��=�n�\���a�96���]C�ŭ��
G�むlG��s��߸�g��r�,%#��m�9����{��O��t�#�7�R�YWJ��[��Cil�8����v�
=�f"���U�����1���D����1�Z�O�_ =�U`/��0y*�f��:��$�^��	jh����;�j����>�� �{����Gv�;N��]��=#�7�� �{�>�M�:���i�ݤڷe��?�~���^ N����tzG������m�WH�������wf�j�x/'�G*���9���0?� *���������#�| E?��s��lDN@* &��`(a
 g��������*�_�u���?�y�'�������s�<�?����2�W��������p���������Ē����G����?��
�����?����p?������3���(����k������n��g?�� ���������� �`� *�*H���
K(14
R�*D��(�(���� �0�K*$ʉ��H�����ʉJ��H$(�@)"ʉ
0
J,(��B�"#*$ ������B ��J�B�
���J�(�@0
Bʉ
!
$����
BʉB�*B�J���J��,�� H) !*$**$�)*$"�
$�
$�*$(�� 
@0�@0�B2�H�
@��J$��
B�*��H����B����@��H����B�$�@H��H@���! �HH$�"HB��� $���H@��@��!��	 HB,$,��,HK!#��,����@�����"0���!

B(0��@���B@�,�2��A!�HC	! I!	!	!	 BHBHB2� H�	*���� B2,�� J�B2�	HJ)!H@�02�!K(��!�@������	0H!! C!�! B�$ J��*� K�,��$�HBHHL��H!�$!*J��
@@) H�(��� J�B���!*H0�0��D�HH�! �� H������!($!�$�2c1�"�@��(BXFP�	AIAP�%PXBE�!E� V�$	!
 �
A�@)A�aIBB�`	D� �dT�!T$	QXFP@�	XFB	A�H�!$!	! b �A�
Pb@��de	TV�e�a�e�a�eaI �FFB EeE�E!@a@HFU�YFA��!��h@�%!B�P �!@��	FA� B@�@�FFP$%d�@�(�B�
%�I	Ph	�3�����PUc����_��-�?��Y���|�
����g�3��������_��U^������܈
��
 ���Џ��J�����'FhPU�w���������5��^��uã�@UW�?��_�U����2>/�����ߌU���U���2�����?�/;5��_�}�@UW�۳<��`��g��w��@UW����Ur���_�����/�?�1AY&SY���d�Y�pP��3'� a�?UP�J@ E_`�     4    R��:���[*�@Wx�(��@� P   
 h�n�h �@P �`t     �T F�  x    �u����@2� Z������`}�9�[��������Y��h�˳\�:{�pzxf��iW�  	��Uqn-U\���]����6�5\ڹ��ث���U������7���ψV�lv�(�y�  7=�A��c����x�w�{��������.}΀=70�/{pPǯT5�((��E)M�q���3e ��͂���PP{   �M�� ��O�����YJR��E �3���R�s�([�����
R�1��� KݹA@\�P��hl-�(
E� �� bhR��>�^�簯M�47�Ӻ�n���ק=�<�{��9zo��t7Y�=x��  ���6���zh��⇝�2�&��ǧГ��;�����7}�x  �� ��P��;��{>���C i�>�Jzp��W��3��{��-�����w^`��8 !���u����O�;�|������!������{�U���w�]��oO�w���  =���QC���t ����m���������9^� �O�-�@����y�iӐ�{ �>'���8  ��y3��������r;�9w0�C�wg��ky���cshv�@p     "~�Jm�JR   ��U)J~���� ��*Uo�  4 j{MTSĪ��A�!����R���MTi� ��R�� ��>D�����a�Y�������pΏs��u��^����PU�"**�����PU��@EV"���?�x�o��M��~��7��ƞ��捱Z�XB�$�i�����9�C_~4I��h��Xғ3Y�s��[�!I�BVS$�_Ce�)��?`K*�gNP��>��[��T#�}ki`�w>�y��v���w�;G{]�[�	n���T�o�_b�ov�(W�}�xƾ�ՙ�3������ס��nֽ�����g��ҷ�6k�>�4�s����N\��J����eo���չ�־���ΈЁ]�(�B��rjȲ�7�'�~7�\����7�p�p���������j�W�tMm�wt���]_)��V���	e2�Xo5t|ˠ�Sg﷩��~$6a��J�U��]
�u�Eޢ^nV}yiis읻�i���
Đ�5�$����G����UuG
������P�Ǹ.w�>f=�e;{�Y!%�P�7��5�͌���~�Ct�lє�ɶ���Np�B��h�i�\7����Y��I�d"n���2S0�&L����m�����Jf]G�d+��۽s/ꮍM0�a�t{����>��?	�(rA��v:0H$"�)�HM!��H�.���|� �i�#�HƄ
����t�1$hJ@��)����jk�j�]v违o*��ݧ���-���k��'KH���g;��l�	 cO�rZ��w�C�V~�B R���B�����"D����A�R����t��K��Ut��>[����D��ghatꢦP��
�On�ώ�}��ϧ?k�E�0�%!�&��!WZ��__�mb�}g1v�e�Y�z�sh7��PR����3R�m��򫿲�Z����o��4��)�45���0����l�ޟ}h�$.����UV�޿���+k��]:���WW}������~� �)�#�$Hh�X(@�H0`n5�$\C�Z��B�]`~�Ч�ƴ�5e��표e�g�>��}ӿ?��#%�7&r�h���%���d���4��F��w�^��I����ݴ��� �zA��6��&;�ԇ�y�C��i���h1���/�05� L�`��a��s@~`П�g4*�T*�Pg)���'�/�[[��}5����}��n�N0��ky3����?�}~����۲,��Jsn��f�?]���|��oL��H�X]R�4��$XXQ��>�)eKHnu���&��6r���j�&֧������2�މ�u}��߾�}}�χۯ���*m,�WWŝ�o��WY�� ��E²�u�ۼn��x�\�J�\yK��p�����������y8U+G����k���T�I��)��w:L�W����}��[���l����+)����C��P�B�Q�1� D�F+����$DlB3[.��}�,����+����w;�����Ue�[��d�ۡ�Y�Ͽl��u��I���go�;����|y��Տ�in�J�;���a�z���y�[!,�x	O$�M~.#:`�k{se����j4�Ip�S����I��F��T�12:Я㱦�E>�f�����R �J���c������3$�@:�FĦ�0%9����\_�Bsq D�X���Ҙ0+)
�)����0ֆK�Є��HQ%k	SZݼx�KP*�k/B%r��9.Z,��B0i����v܁f*JD�c�G�x�c��iY�ǻ��.��+���1�Dk�)f�n��Jc>/6hԎ܅I.Ɇi��S\ϿSU�3��۸vFI�O����ͯ�kr*J˟fJC6�Y�w��bB���4c`V����.:!F��$`Sf�\�.���p�/6��%#HH��W$.@�O��ޡ�20�@�
i���<#d�
!�L~�i��R�Xˆ���Wc)�FD�E�џ��Y	_�!ܑ��9�ݷG�L�fÐ�#�Y�q�fĪQ�~H4�!+
B�,
���!��l����!$B��)$��	��̄"j%sQ28P���F#i�He$�2B�3r����@�B�Ʋ��
�U�Vt�l)�M�>���!p���B�����~e�������I�!�|���n��f�L��Sf� �A�,��0�ݛ�.H�c ��k�HM��,6G�e�l�E��	BHыv7�
��@��.CF�sK� !�!�0�٤�B�7B�6@������D�����"�[��S�l�!G�>������~�H���a�HI��%��u��$_�+�V�\��B� FJc`D��c`D�5�||;a����ĒF���8�(cVH�I��bm5*I#���t}�����2�\���9����P��Ԑ��	 ���!#�l� �Hp�A��raN/���)���Hh�v�w�p�6o4R3����I�	$�nϹ~�n�~5	�i�����w�L,�/ƿa�8�a$��p�չ�0d	.�\`� \5�%�l�ʃK�.!Ąa�p e��fkS"B`KJ�a.s�{&�3V@�d�5$�X7��C_�@�T��i�!�C6E@���:J@� �ˮY	�1!�4#p��!R  �- �@�(Ga	!bY���_+� ��f��Ie4j�8Yz���ç9���(Q$CD�jX5�F��~��C���R7��4�i"���>�B��m�Ƶ�M�n�P){�$	�ZL4�2��!����������1�i� �`CLX�	�8��D�R�2��L%0�	y~���#s�Z��BQ>'��t2q	b@�LK��$��H�L�$�HJc.1�a)�����p�a�B��U�@čs3�܍�� ]�������dĔ�%2S!R!XX�I/X\��S��M>�r��nvG��#H X��R��$E�ˇ���$XF�����~y���$%5�nkv���8]����063EHP�!8�:$5$:"�֍��+��cV�4{I���~� А��i�$Čdg�M�I���w�\�8����j䑌������㙭��]ZY9�|hIden���v����D$�bE�S�Ȥ�SR�B,`Q�S0�M34f��ɨx�/�F�K�y�5���mܼ�уN�5 k_]�$�~l��Oߤ�ے�d2m��R�y�y�����9.�A	�r����i!�����!W��ևGڮ	8�7��2O�1�ͿM�)���,��fO����P$HpX�$!���Ѱ:Jq�0�K�!Rv!p�ԁ
�H��B��+��� �����<����.y� l�d
N7��`�5���$�~vs?I��tCI	\������ >̢��͹�.�<�L�LѦ!D�֬�O��&R0a��ߍr̿h�R�XZ��@��M��F�� B�������S�d�R�SD����t������aÔ)'��ig�9���}�܅K��T��*�Uuw��^m}d��)/�J�o��N7�s����#,�$͓��s?D��!M�0��5Rn�q��ܺ��o[6t��Eܲ���, doTN�$�:�4 Y9�w$�/����C��,˿ٙ�.��ڻe	zY`�K���������yb�����4��K$�~-�9�K7�K`]�aB�;	 ���\�	e٨F�E��e�����E�0��b!"A� Dk�)��k����#&�@���	4f��v�(y!��_I͆�r�W�P�HT� ����0��$Rz#�S�
c%,��\,�
:�H�ŌCb�oL��e��ӟt��Ϸq�͸M[0��]l(J|K�N+Z୔�B����ߖ��f��v�&��@tM�>��~8�l�����x}��Y�]uC*H�p�ލ��4L���?~8�d)�ۮ/h��\!������N��p��C�g*�,�n�Ԯ��G&v\�p&b2F"�a����I�ln��埛f���_� �I��.�a�5�p��}��$
���������d�?.CY�
�C:p���ˉ1��F�������7�_�!��~:a��>�HA$WE)�7�w�sx_�sp�΂\Թ_>�_<���$��;	�&Vԯ�9�}�<�h�ϧ��OK�2����ޯ��q�����M$��$�0"�0i�ha �'�-����F{wy�}��m��i	f�B������X�	�kl��79L�����r'@�Y�}.�W�-����\��n6�O�%974��*�a�.2�LK��wNM7tty���Y��æ�e���h�P�
�0���d�F�s��-u3Rؐˑ���m�3�D�����ދ:XMI%6i$oSrF���s����k��i���w���$�1��e�\`�4¸0HqbD�� �]�#-���~������"��)����"�Ζ��@bFı)!HŌR�R&���G���ȳ:�*Jz�I�Y#a�$�˦:�aHƸh�Fu � ���n���4k[�_��s�g>���s)NC���3��r��|��,�ѯ��k�2�>�7V�ߦ��[�w��/���J��Ҧl�iJ�s���jY,>߾ÔQʭfp�37�̱	1�����I�����~�Ϲ�m.�:��/��\(��}�ˣ��ٛ�;�������r����vϫ��:l�u���v��}���u�/_4�!�M[����J��*bN�	��M�I.��}	����ʪ��UUU[UU*�UUUUUUUUUUUUUUUUUUUUUUUU*�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU]UT�UUUUUUUUUUUUUUUUT�UUWUUUUUPUJ�UUUUTT�������������V����Z�*��������������������������V����������������������������������������₪�������
�U�&�� ��t���K�y���P֤n#u��%�WP�Z��:��P4H	eT�cm�����#��)Ij�۩����.2!�j���f���V�y�Iy~�yo2(3A	�ↈ`���[�͛a��@ք�s�{���X.v������Y6����U!N�0MUUUUT *���٫j�촱���5s��[��zUuK�p�Vʵj��{�l+UUà��v�Uh�im��n��Z�S�9n������U�]�ѷJ�@]8�U�K��4�PYIA��]�U	�U���ib�Z���Uʪ����6��4ZKU�U�S�媪�ڇx�)�!��[�T�9���NE��&�P�F��s�+��6y�M*�&�*�UT:v��U������86�VV�Tu�U[]VH�q�o�����⪪�@��h)j�)B���%*��v�V��0���la�U��W�M�U�];�UG�8�v9��Z������
UUUmV�U�UPR�����HG���&��h�Z�����j�ڪ��aU`��U�4�UյU]��`�xL5ON�@3�]F�*�3���ڮ�W �P�ڹ[��U�v)V�d��ͪ^73��i6���`&�r&nZ���)=F'�Y^�%V�pE�w�3��k�������5�V��bܼ��ɟ@A�;g[S�-9j�Ғ[�ni]q�9��0��ڝf\Vޱ;9+�)-��S*ф��tr]���h;��9�m-��f�'�b�
꺩�6T.n��Ү���e��u�T��T �UU"宬!�j��K-P�ݞyjT��u�dU�p(-��OYn��8�2�V�<�l�kl�s.�uUG <�El9jکWj���A���-�����癖��
�q�a�u��AȺ�GplrX-3hv�g�L�*�
���Q���UUU�PWf{*�uJ�[[U@�UU�������
ej��j����V���^Z�
��en{	M:㮹T��(J�R��� ٝ��Sj>���PA���|r�P�� ].�j�����乴V�J��*�U�R�T�#
��)-�c�誩W������]V�@6��U�Z����vU٥Z�����-*�U�UUWR�W+� ��PUmU��J�����dj���UU2Eҹ���S啪���`VyUUiV��Z^Z������Ԫ�UUT��R�X�[��UuV�[UK�j�U�N��
ܖ��m�TNs�x���U��UV�4pT��Uk�������>hj�
�iV�ꀛUF�����wV��մ����v�୥Z�����U<���Jl7 2�"��Ώ���j�\fU�l���b�N�.l�M*�]3�j�MO�1�&��E��ETU[UUU@UWUJ���*�s�ٵ8��[[U\���l�X�̛�h��� v�VE���`�j�(nU��U�����z�)�	#):�j���\��U++\�U��UT�a��vMO)�s�F�ne��7] X	���j�Pp�
�<�G����C��ݬ��.l�%%�m�&'pp�e�P�<R>���lr�gE�H�K�V-$����0�p®Xk��UmPIټ[�n6�i�Yy����t�t�Q;`
�eP��:0�1����N+�UPԲ�W R�ە�j�M���V�:g�u��:휗�WU�<�q��c3P7YT�c9�GA���}�,���x�km��9���M�Ġq���F�;4q��w2����Sc�`�d�(p�P�Y��1fk�A���c��AѹӴ������p�\�y&W�-ٟ)J�<�̈́�jcl��"�p�5��X�n�MW.��O�;����Y��\�ݲ�F�֧�[a����E@�M�Q�PQ����&LJ(n�Uk���U�+��Y�s�j�d����\��i�3gZ��=,��r-��H٬vq�E�\m�ٍВ�y��:�*�M����e��!y�A��m�\�nM٥��
r�8k)q��;U���T��6��1�K���p6�ힵMO7��5U�>]�(�[�����i�	UU]:�'XԵ6ڠ�j��y�*k:vZT�׶V�*��R��.�8��UPҭr[�UW��8\CT����o�{�mF�pvү[T9�j�]��ڥZU�X� ��UUT�V4]�zW��nQ�j���������V�UF��{eݗ��ب��,��lcf���YWX�wV1�+q��'��;d�5e`X��.��X^N�o8q�y�)���K�eٷVm�vU����n�z�B9^^����P�nk6�e
vv��)n�{u���ψ����Yl��QV,A�˨]<v���j����Nllj�kyZ�VV  tn�l�mUT誕j��8���UV����S�xS�; �M��bÐ���C��m�6��ӌMU]@ru�Q,��m�*Ԯ�(*�����
+��նΪ�.��¦J�j�VV�P]UU q�Ԫi2�ks��m��UUHH�"�T�F��H	����m5UU*��̭U�5Ʈ��vj�UZ���e2II�d&�ev4+T��Y�檪��Ur�E��j�U.�Ha�H�����U s]Uu�nԼ�UV�[UuUUe%�r*��V��UV*�0�TWEU����r�R�~]u}R����Uu6��G�5�ꪐ�ڮ�vU�����	°UUmmuU�gp�p*�]յU@C����D5Ui�xG�:��v�[�Uwej�W��i�[�
%���^YZ��nا�S%�ʳ",��s."cQJ��P�\�����tD����`UU*�c�*J�½0
��4�˷]���ՑK�U�Lq���6:���SG����=��I�z�Y�e��Ts.޸�dhl=hBj��n�j@Y%�Ey�l��v�M����-^C\]�svO[���x▝��5mR�poU��ط*�p.h�5��*%��\�$��`�U���mѡs�ƭ�i���MU*�K�� U@UU�V���vZ�]���+�[gl5�ElT�5r�MT�,�UVԫX���z
��Z������U[�j�ڮ��Ul���UU�� z�Z�
�]�W5YV����^eBk-UT�i�7;g+U �UU�U]]J�U�P��T�+p[UU*�J�,��UUU@[]O+���으���;ʣ� *�`���>�����V��i\�.�U[UUUUU�"���M����U��Bj�v�nVU��Im���+5�*��U�+���ղ��vPi[D�v��:����SC�V�@-����N�v�*��xJ����\�.qiОB�c�5����m`	�m�f���ɮݘr��a�،��V�tG�:2@�I 
�
��m@\v��k0P�9I�I��2�C=7H��]�Uu)�(�<�mYH�j��UV
�'mP\�.ڐ��eZ���+T��6�T�(q�:�VW`��|}�4p�W[:**���"e�v��UUu]=)0UUHQ��)�(��;mJG��L�5V۵@Isl6�O��PqlszWf��R��pj��g���J�:�j���Z�V��d���UUF4����g�5]UUU�V�^��v�j����X+�:�Z����jZ�����f���*��}���U]UP���dr��UUUU�Um�UPUm�WT����������J&� �X[Pe�bam=A!DYL�L�ȬV�m����h��gi@��fj�Rg�a	i[k���!He]�,a�ev��*鸡5s]J�Ul�xW�U��v	�vU���9�k]U/(UUb�AR��Wnx�SB�W]A�WC���媁 �W���TuFFWj�̪֫<�!vZ��+��UUm[N{K@UUr�[Sf���"Uj(�L�0�DݝT��`*�����Q�SU[H%�pUX��)�N������UUT��tP�U���8��`%j�V�V�G5s��ѐU��Io���v�*�UmUa��L�b�iW!��ٮ�q�jRq`8ݚ� ꥨr��h���v�U��g�6܃X��|��Cc̻ �����(,P)�Ա�ѭ�,#�f��ظ����Arˣ�'`�S5*ݵT���N�ܶ2@ƭ�Ԫ�U*��ʹ��P����i��*��v1�6%j�ъ� ����p#���6X��Z�k����<�ej��U֦�3�M6�(zm�/(MU@)(aQ��mJ�UU��6g[M�j��IdHT��xf��)V�
�̔�ƶ1Ir�U�B��U`�5\�UUT�U�U9J���8��[iV�,��ε5
�M�.^�Z���r�d�P��luUU@UR��U)-�Us�
�������}U�T�P媩�j���b��ʪ���J���V�UUU�,�4�ذ��hٝp�Us���Z��Y0t�-#l�U�[T�u�������U]�\���H4kQP�>�Z�y	��W;:B^�U��6:�jYC�Z��Z�[`t��&Ԫ$tAs�T��@6���ဨ
U�V:�@Z*�U��,�8(.�*�m���*k�SMC0��U�ij�UUK̓��٤�Q�M��>_�]�����gu��UUR�Z֏�AQT҉�&���P4p����!�º>P5!`�F ����l"ŐH�O����SoT���QPқ`'�( h��?h���LR�J8
�J�n��NpGb~����٤r�4
��`��� �J�jj"=C�I1JJ0�dH�@���C�*5w^��v'T*
�>u�̂���� ��Ag�t ��0g±�"��B	�j+��Ӯ�T���K$HBW��>@� �I�����|�E�H���;���"�Ab?" |�DȬT�U�hQ�S@?������ � �Q9�0@��*!ġ�U:A@8 �(@CiB��(#�P���D�DA�/@?X��<P0W��&�(��bA�Tq
���6����A��
�"�����U�p�����d�
�H%i
��J�����@�9�$�W�
�~C�����E:�C�(�a�0�\0@�U����Q࿃�tR3q�YPQ4����'���S�6"|(I�iJ�XVД�! %!"�*H#X,�! Dc`� 
[lb���~���B�i���62)�T�O�u@�$@�vh���`*m
|��:��ꀊ�� ��N0q���D"#! H�@@.(P��R�KK"��HU0 ����'/'e�PUUUU�UUUUUUX������ꪪ�k�������ꪪ����V��콞պS1�7L糃OF7I�Q-�oh� �ue��QN��N�IU�b�dCsU��Q`��eesU5�-�mʻA�T:{"���=;6��jS������L��ϕ�d;g��n�l�7�K*�UŠ35�tƙ$�[��n��Dv��7nq��6ky�r�(w���[uR�ew.3м3b�7�x`�m/c��g�5Kh�ɱ�3��3]�n�^J�Q�n��Ef����h	�L�K��ݪ�ݺ� �̦Z��\j]V�-�@.uC<S˶ۓ#�[����j�+th�K%
J�^���R� +v�L��ƺ�082��I�[������-�A�';�^Nǌ��	4�����vx�ͭ��.8��z{gf��:bњ���k�\:Htg�aI�y��"tg�FZ�kI�$�v1H��k�+c*m����x���8�/X����;�se������g��Y�b�óۈ�9x��{A�;gfv�0��V��\�F��=qN��Eۊh�E+�ڀg�^8��S%q�ۢ���h�Q�r�Δ�f�`�f�@��[�����\U��+`f�AvT�ں����爹X��5�]ZDf��C�yv���EX=�m���D��X��C�˰r���Qg��ϣ"���igr���/Ti5��֭S�X�6Eը�c`5ƈ��kMu��nH�v���N�i���s���ۧ�������5���<����6���F!)��%U֔�YZ���`6���Eq@J�Z�ܜ��s۪w[�zk��6l穲�Bn����+v��vʠm�I:ê�NB2l���l����Ԝ�C�i��%�!���G=w2�"'֓6.��%:���ݩ�)բ�u)�-LTc*�١X�fcY��j�J�  �^V����Ysl�B\�D��N{]#�ޥi�<�m�ܣp�k.�f��99?Og$��v�(ES���� 0E8!�N��_�H� �799y��%��z��6��f�R�"�d�3�<��՝B��:������Uh�<�6�!���wBe����6WHinBG��u�v���!�u���͢f���r���cl�NZ�ވ����X�m�e�1�f^mƤ�1R94q%�i�l�{k�<j
� @��[e�!l6�7X|�rn�(���۰љ4K�����Rf�j���j{�����eX��-lKE��hX��k�%-lX6�е��M泖����� }�� �����r��A=�� ��z�*�5e+�ZWn�nǞ������{|�`����J�eYƮ��I[x�I;0[��nǀ}ݔ��WW�N��n�o ����x7c��lx{��Ҷ��*�Sv�Wv^ M���<v8`�W*Hz�M�,tI��F(�V���1�m�Z��rZJ��tP��|���,сv��i��� zO< ��ǀN�Wv^���m[���A���������Y1�!� R԰ _]���߾��)�� ����ģE]'ce[M:M�v8`�e��Us�H��x����7d���O��$���� ����6<v8`�l(Ec���-+�x7c��lx�p�5we��{�B=t|��\�m]�M:*a�����ΰ��&J�u	���3�ce��!S�8��n��o�׽�ou� ջ/ >����ڵu|t�[v�6��`�e�ݑ��$y�r��=���J۫l�n�;f�� �������P$��ȄA]�A�G�a��[�}�uٹ'����M]]�M�t�n���������/ �l2��V����Ю���lx{��� ��<��[({��e�,Ì���á��p��f״�U�N��S�����2�;JVu$��ݏ���/ >� >���$���O��$�����W*�������w��n���yMYJ閕ۼ ��< ��Ǉ��-��`l���*T��g�mZ����ǀw��|���%{���3��\�$�6������wu�Dr�ex{�˻/ >� >��x{�}��#�I�kW�{T�*ʨ�A�j��SAc��&i��2\�Q�Y��2W3 �we�ݑ�ղ?W>A��}�^���`��N��� >� >����`[�����;-���Е��V���`[����5��V���ݔ�+����ٞ0Rz���ղ<�@�m'b�O��$��V��\�]����=�nI��ٹ%G�A��ȕ�RB*�H	X�Q(I%���߻m�j��a���
^z�v4\wڝ-n�I,"6��Ҵ�PʂJ�H�[���F��%�;�L�ʺ6l�N�������HMn�l�r)R�Ϳ��B�'^{�g38yݡ�ϦR�V��l�M�`�Q�[0i�j�!.`������&��5\mMP�Ir5�Xi�س쳃v��Hs8������3�"y1�a٤O�W���+2��y9<�%�@��#mЫ r9�r���.#���W����ͭ�%p�j�3f2��
L���L�����y�ղ<w\0��xt
�-,�����x�l�?W9ďl~0Rz�wc�>��W�ի����n���N�ջ/ 'v> O�׀{:=e̤�oԶ�������dx�ȰȪrd�d.e�r���� ��w� ��ջ/ �s��-�������F�S���sq����k)��<]赁��7N��!K��A´�/����<v�XV�s�\��<�	��^wk��D�G/ ﻽���@��5�	-�%!f
�~]^ zo� }[#�7vQx馋`���Wm`[��nǀV��	۝��I�HRn%��&�gp?I<�[�<��=�}ۑ`[���*X�%g�����dx�]��/��'� ;ݏ ��S 5H,���Z�u���[��Hn�fk���,E(�f]���Vz��3U.�h�.\�/ ��w��{~�� �u� >����84[v6��*�un��;�p��dxݹ�ݳ��i�AÕ��~zp�����H+�E)~A;��O�[ŀuM��}6����m��V�f }[#�>�Ȱ��x{��m�v�7l�&�9x��zpo�wp�\0������IC*�7�5�Gsttf]��/��V��m6��c���J���i�|]-�8�ﻸ����ղ<���4��E��wL�����g�������un��RF�+��	Y�U۫v� �Oy�v8`RK�;�p�>셫�WWWL+n�;o ��� �^���T�	���	���@�p�y����n��J�"��`RK�=�3������0�Z'R˷(�5�4f�b�U֘t�PH�(�ͥ�p4�X�ͱ��رM6+\-]�=�� ml� ��� �^���X��V�Ql�� ���c��$����4�wk�]۳�˧m�v8`RK�;�p����T�ct��>7t��`RK�;�p����v8`�TR/)�tēn�	�2�kdx�p�:���s���r���,��^K�m��[�
�c�Jp��Vʽ��4X]��v���.�&����
�4�<�P�/����O$����i��:7@�h�X6Z6]k`��WJk0�3`KD|.#z]v�3��\b��\��>���`48�n�p�)�0�6�� f04Ԍv�3hыQ\����R9�U�sS�6�w�nNɜF�&�U������mp"�a�g��5��I3��LLH�zI�úXg�g"�h�ۗz����%˞�X��ڛ�Օ3g)�<y�ca����͎�+8*�Ҷ��W�~x�p�:���Mٕ�}�W���郥mۧm��� �^7fV ml� �`��mն	[�U���IxݙX9T��^���?dU2�.�Ɔ�v6��7fV�jK�'c��$����w7\���3�}~����� �^7fV wR��B�v��+�؝�j#����-�/�9z�)t��Z4]���>kvb��z��RK�&���9��R����{���%�x��z ?������rI9�%��0��"�
��7�e�F$��*K�䒛Q�$��QŻ����2�� ��ދ���Ӿ�)���K�$��I.�2�]
�
��V�1$��9�$���I%��/����z ;��ۍ�6�F�2�rw�IM�(Ē]����$���Ē]�r.� �NNI��Zu����Yb���#%㱃�ևy97�؝�ē��Ip�m��j�`fe�32�� y����`���z ]�r/�I)���dP��][m46���I)�2�{��]�[)���K�ف�$�{%���ʫ�G�Q�ݶ7E%n�$��O�_|�Sf`b[��*�|�_�0��.�����$'YI~���BC�iC��J��XI�H���a��o���
�dNf�3&�>&��"�ւf���ғg�MF3he[�]�t��?g�{���!���!�*wl �j��H��������R��H(dE6U�M��`)����{�Gd�$���) ��REc�4�i�����Ϧ� E>*z	 U輲���YJ��+�>�TF1�&��o��V5��5�('/� 2I#&P�C�N���'���_�vDz;���������+?~��I����Y�"E�47��E�B1�%�r�jK,�����u�����XM�@$�\�H�`~��>�T�� =S� ��AS���%�lUC��E���`�< B��:��*Kn�I|�]�2�$��wk�]��n�k�Jl�I%ے_�$�ۙK^�s�mﳯ�;��}��WL���mĒ]�%��IM���$��9�$�٘^��a��% ���˰	�q��]��"۪�Wc�;N�"G+v�ۋ�8���tY]2�+n��$���X�Kv���Jl̷�rw�o��w���~��S^R9�ۥ�$�iȾ�ܻ����Ē[~���|�����l�����i�R�F6��$���Iv�K�䒛s)bI.�>�w���޺hgL��am������r�{�weݶ���o9m۰�� @�T)U6��X�[7��*� 08�$���[������2�	��J��� ���P� �s�IU3�]�I��$�{�1$��Ԩ�^��\ ��۞e`��v��'��7�o�g����V�q��qaZ�v�n> ]�9�$��px�K��_�$�v�RĐy糩�v8��E�N� �޾�����%�s)bI.�9�z��E^��i�x�t�.: <�}��<����ݧ"����I.�TR���+l�2�� ���P� �����`���bI.ܒ��$� �����ӷJۥ���Ӿ�>�9'<������n���weݶ�&"/�$�
 4B"	R�2w]ֵ��'OJ�UKF��t���+�3�^ڝOn�3*�^�2��S�ú�fq@m���o��#1�hb&0)�'l����� �������6?����ܱ��U���6�E��X�a�Z�0��A��0�i"-0�z��Zک:b��Q_lF%���،]#��G�[՞I��&�mU�8&�8u�K
�V�	��-�AnQ�.j�5���e���C��9%�ަ!ܡ�a{�y�^W��26jǗ����n%��h�dc�+q�i��J+X���Ij�y^$�����%�s)bI.�9}�y���-���l���y���%�s)bI.�9�$�Uȯ?�*��߾>���mr%Qw}�{���t wiȾ�*�����Ē[s޿�I#oj+CM��*�0��y���� �o�$�����/r�~��$��Օ~wk�Xg�f*w����= ��޾��y�޿�KIwiȾ�$��l�E]���ŗl0[�^�taۊ//��܏<]�2l�q}β�/SM��;j�����}�[�2�$��ӑ~�W+�_����D�ߓ�����a���l +���7�C�ʜS��̷}5�^r�gs������������9=�e����Myts�� ����w����=�o7�}���w�C���}���M4ma�c���/Z��'�$��|�]ۙKIwi���`��z�΂�
&� ��%��Iz�?}K�[)���K��+Ē?NI�O>�����R��1B�f��͹G;O��ޖ���0]qӺIB�벖���[m46���$�_��$����>�$�o=7@{�}��|�OL6�l�*�X�K�[���꽊�$�ײ_�$��7�C����}f�pL¨�[�e��ϻsv�y�w��_�a��F��eKE�$�e�l��@9��KIl��}�IE �av>:wv'm�Ē_^�|�]ۙKIwkr|�G���� ���}-���M���ݹ��$��쯼w�$m�'�$��쿾H?N{�J_�;���E.�ڏ,t��X�h$��H�"�2�v�R84C4�30~;YoNo%���E�K�$�z����$v�'�$����?��{�� �}���i�k�b�� ���G���T<���w��o�C�)����o}�$�}�zCe��l5�w�$�{=|���2�%�U����|�_7�@~�{{�Y�mr%Qw}�{����X�KvVx��;{Ė�eQ�A,DW�
.���O�E��7}�_w��M��*�S:X�K���}�Iyk�O�]�{�����z�@�ϼ���!�lη]T1�,<�㞀�az����nͺX(B{=p[1�/﹭���\0�Q�|����= �{>��I.�̥꯮�[����$���*BʹC�v�z ;����}�����H����)bI)=Y���;{�Uݥ�x���&6HAs;��w�C����׷���U_��%��x�Kg��W�$�aAV��^]�,: ?���{{��o=��w�9�o�	����~.�����8\0���(귾���� ���I�Ny���[�%<�b1$�wL��$��h��Pp�[��UU�*�UH��Y��	��;^ag�ۏ.�͐zn� �l�ݺK�&ᱎ]��J6����f�f勁t\T�2X���S��fz�@8R�$XO���CUf2�.ԺELЙ�� �S1+33`���ГƘ���i<��i�+1��Ķ�AkV;Bk�:�qΕ�^��[l���h�e��i�r���[�z����+N���Rjo1�nגrOd���<���'?�q1���5F�XB\������x�r\��$ԇn�1��o߾�����Rg��w`�~���`�>�^��<�W+���۞w�$���][m42���$�u�F{�v��g��I%�<� ��������������l��`R��6A���c���U%������ˀ{�v����Qj�N�<���'�r{��6~���}ۑ`z���[!�0/W�X&��wn�o ��e`�+���/��� ;ݏ �U�mR�c�C�0O6�W�ϱqa�t��'����g��Qk�����&+z-	���΄3�o���,��� w����W�;��V��_��8];h������_r��t���Bar������ęp��K��q�1��"Y�I�P���(Ԟ����;��f����ߕq#���)]��J�N�� ݞxݓ+����Ur�K��`�� �ȯ(�N�j������W*������v��wtp��*�U�%��<��؆�Vf��W5����s�w�rO�D�C����{��>�X����X2�v[l[p�jD3
�͔�� -��)�l:XU�����rp�u:04�,���2wm�� �ve`vL�s��+��������Ս]+aci�6`veg�~�W.͟�e`������W8����
����;��Xw���'nE������`�
� �* �Z�B��U���nk�nI���훒w���Zum�.gV�'!���Zl��Mٕ���w���x�BK�gN�+m`�0s�$����{+ �\� ��2T���R`�
���D�^���E�fa�,0]�Q0 5�j"b�ܒM���K�4A�(�O�;������e`K�{���6A��6{��j��V:ݺ�>�Y�H��X�?�}�N~��i�����Q�i��m6f�_���~�Ur�s�����+ ���V }�QZLWv�
n�J���W*��g�I��ɕ����VW;WH�%����R�$����d 4�b�ʞ���r�I�������n�Cf��+ ����[?~�t��,��� }�"��JSx�����V��mT�x� �jt��;[UkB8��?�y$�#`s[|ev5��߿~��K�`�?W+���\��{����o��_��j���*M۬�r,�9\�r�6A��$���>�Y��W*���Jt!z�e+��J�X�?�̬=U��9Ļ��V�_��� ]�]�L+lv6`~�W��9\�/��������r-��!�����?�������L�SY���m۬�ɕ�~�Us�r������.�'��0ݙXr�9U��룕J���V�L��Ιx~�L���	~j�C2|�Ӓ��Hp�Mrp�z%ֶ�B�m�9��k{	p��.5�2�M!M�h�B9�鹸0�։u�SP�3	(K�"F�k�C��	��$�($F@I#$t�BD"F�K&���A)� � �ʁV�dMb�ĉ�Slnȑ$�bQ�*CbX�XB(A] �����	$�1��A��$"\�D��H���b�4H08P��HI�,03��p�(tY�K��k,���N~�����7�f��ZYM�|�~�B*����UUUUUUV�Z���U�����V���
�U@X��������VZ�]�]�l�CPB�u1����.3��k�t[kYN��G[sv�ݙ^WY`���`l�U;1�"
�߽�u���.�(���	S1#������P��I�t*h��fr,Mf���%��8�
x�M�����g���%f,,�InĸFɵ��Ď^��g�v�Z�>���,ᚇu��}u�:;al�Ė��!��G���e��9֪nkc��e�(��>���!�n9�t��vr1 i�� �(����u�hbc[d��y�ܘ�0���W&�(�Y�k��-�iR!I0(�p��vI��(:\gV#Ë��S�5kD�.���[�i�j6[�5h�J:,b�+��8��%��=����p�{U�뎝����\�m�HM���A���mp�.0�)K��
X��%c`EcbR4�y�6Rӧh�)�v�g��6"��upB�UA%��u�i*��$����8B��������^Yؽ=8�M�[\]q��^��
������;�g�^r]��h֭��%�Ѕ5	v�-l��i�Q2Iv{
���n%�\u�ǖ6�)(r����vڌ�A ��'��έֵ�@/4��
��Sʲ�eC)s�-Ӻ�+	�Q��,0��z׍\��a֜��]�ȳ�Z��m2�y��3#iMي�X�T�7!��ZU�|9l�o�ۛ6�`EDt\Җ:���.C�F��1���Y�[�m���9�֋�#�p(m�5���������a�kh�X(��dSlc!�PT������V0�[�$ͅ�2(��\lJU�B
� �l�ܪ��ˁX�s�e��̼�m��t�֬�]�gm���Y��¼�6y����.�ͨNw+�мc:�[�t<�J���^��r ��Z�|�r�m�c�[��d�����/2�Q�����<j���B[��:k;t����u���%��`�|�Mf�%�I��3&��.��!�T9�P� ~U �|/Ȁ�Q��P@~@P�_��/Q1R*��_�_�ڗn�ܵ%8v�n�/%��"sɁ�d�fh�L(�E���f�6���4�c����ζ*��[��`�$B�{l��v72�b[\L� �ԅq岔盂�E)MJ*�MdfVK�`�v����Ѳc<g�s�9FN�n̸cx{s��i{P<Ykq���=`^�6��	�ь7��iI�{Q�/gCڏ�q>�ۢM�'�3X�a�5Meˬշ"J���I.�)��a`�ZJX�e���9r`0���CO� n��& �bXͽ�����OM���WWV��m��u���׀w�N�f�(,����nI?wǮZj��i��B+w�w�N����W.�O~��6~���|�����KO�M�?3e�LլS�M���>�X~�9�~��Uޯ��x����j�D��m.:wv
�`z�ʥ�{��:�=x�W"��*�Jl�Հo���9p���s8������O'�����&�e`[��ۡIE'tn˽�<O��W�\]n��U��aL��mT�Г���I��)y0��6]������'߾���=�w�͇�E@�"X�'��߷\��B����{���w[�k�F�WiȖ%�bw���Ӑ����,F�Z��a`;�p���,�m�j&�RD�K��~ͧ"X�%��｛ND�,K�M{�iȟ�2&D�;����3h:95e�s:��������}���D�,K�{�ͧ"X*�%������Kı;�}�iȖ%�b}�O����f�]D]�'w������*~�wٴ�Kı?t׽v��bX�'~�m9İ?���N���ͧ"[�^B�}�_ڍ6���L�;��K���^��r%�bX*=����Kı>��ٴ�Kı?g���wy�^B�}��%��5�̪�ٛc�ۃf'����Xȍ�Ÿ�L8[]���4����GNӍ-ƃ�n�b�>_B�Љ߻�ND�,K��}�ND�,K�{�͇�0T?DȖ%���]�/!y�^O��ԟ���/;[�:��%�bX�g{��r(%�bX����m9ı,O�=�ND�,K�w�6����bX�z���&�W32�R�ֳiȖ%�b~�wٴ�Kı?|{�6��cP긡Q0E$K>�m9ı,O���6��bX�'�	�r��&�p��u��r%�g����O���ӑ,K��}��iȖ%�b}�wٴ�K��AK���'$<����]ɜ ʭe���I��wI�$���ﻛOD�,K���m9ı,O���"X�%�߾���Si�K\�ĕ�1�m�����!FLLf��X�JgQ���ص�I$;�<Ѯfq�D��f��"X�%��}�fӑ,K�����ND�,K�ǽ�j��bX�'~�m9ı,O���֡�Fjfk3VkY��r%�bX���si�"X�%������Kı;�}�iȖ%�b}�wٴ�ElKĿ��{%&�f�I5�\ֶ��bX�'�{�ӑ,K�����"Xؖ'��}�ND�,K���m9ı,N�׉�f�T֋:������%�M����iȖ%�bw;���r%�bX���siȖ%����`�� ̣X!%Y�R���D�P#�ȟ ��u?�p�r%�bX����>��j���ݙ�'w����/'��}�ND�,K�`��������Kı;����iȖ%�bw���ӑ-�/!y>���Ж�V���G���qȬF.mv��uv;9ʅd3sn����y�L�6ލ\�l4��u���/!y�}�kiȖ%�b}���m9ı,O��mAD�,K���ͧ"X�%���훙o���љ�3Zͧ"X�%������?��2%�����ӑ,K��w�ٴ�Kı?g��m99'$/!y����jv��w
�S3iȖ%�b}�}�iȖ%�b}�wٴ�K K���{�iȖ%�b~���m9ı,O����e�5�Y��D���ND�,�>ϻ��r%�bX�}�z�9ı,O���"X�+b}���iȖ%�b}����kS$њ��噬�m9ı,O�׽v��bX����~6��X�%���p�r%�bX�g��m9ı,L�l�,���'О���Ucq�շT���Z���Q99��cu�v8�l��%��f���b۸ue¶���q��cs|&j��3{j2��o�ʮ�W��tm�u{&CL:ʩ��+��3R��1ɣ�n2¯���b������p7M�m.��6����� BV8��[���>�<�s��^�j+��mq��֟,�c\��ݸ犍te�i$��Hg�X�V�B��fEԫl�z7s�o�½�CbjZ�b�R�N]�/Z��L։&�!nk[ND�,K���6��bX�'�{�6��bX�'��}��Kı/�{��r%�bX���u�.�M�rwy�^B�y��p�r���,N�}��ND�,K�����r%�bX����m9,K��w�=�
]:��fd��iȖ%�b{>�iȖ%�b_�����K ,K�t��"X�%�����"X�0��}g�[{5rm����N�!y
��~���ӑ,K���=�iȖ%�b}���iȖ%�؞��ٴ�Kı>�'M��,�.��f]k[ND�,K�x��"X�%�����O�,K���{�6��bX�%��{[ND�,K���{8K��kZ�354�!����u����R�k��>��oYE� ˨h�4�>OG��^&pol�Y�'���Jy)����m9ı,Og{��r%�bX���lD�,K�x��"X�%���_�x����ݜι;���/!x{;�fӐ�=A]�#��W�2%�{�}��"X�%�����"X�%�����"��C"dK���������l��������=���m9ı,O}��6��`%�b}���iȖ%�b{;�fӑ,KĿ��_�%uV��2u���/!d�/}��6��bX�'�{�6��bX�'���m9İ���{�iȖ%�^O�����u̌�,듻�^B������"X�%���޻ND�,K��]�"X�%�����"X��S�����-���!���@�vLS��H&��]ڞYb1..�0�6��zIˡ90����fd��iȖ%�b{���ӑ,K���{�iȖ%�b{�=�h�"X�%�����"X�%��C�[{ˍ�H;'\��B����x���?��L�b{����Kı;���ND�,K�׽v���bX�'ޒtٔ�f�u�5�5���Kı=���Kı>����K "H*���E�,�n�4Q�BUE�H�$"H��X�N	��Cb�S�*����ֽ��Kı;�{�i��/!y��}��r[��e�bι9ı@���{�ӑ,K��u�]�"X�%�����ӑ,K��������iȖ%�bw��e�sXk5rh�3Y�iȖ%�b{���ӑ,K�~�^��r%�bX��8m9ı,O���m9ı,O�������P�Ќ�o9������k�2�6�ή��JZ�1=;�,��칱G]snT��j�?D�,K�����9ı,OwǸm9ı,O��m9ı,Ow^��r%�bX��zOd��\։&�$�5v��bX�'���6����bX�}�p�r%�bX����Kı?}�z�9�P��"X�����]��de�g\��B��������ӑ,K��u�]�"X�bX��׽v��bX�'���6��bX�'s�)�]L��3Y�.h�r%�b�'��z�9ı,O�k޻ND�,K���ND�,?��@/6�D����iȖ%�b{�{�Nk53Z˙5)u����Kı?}�z�9ı,O{��6��bX�'�w�6��bX�'��z�9ı,O���/�7�e�
�'�:�2��#n.����kTi���y�"�L�;�D�:)[�[����%�bX������ӑ,K�����ӑ,K��u�]�Ȗ%�b~���wy�^B�y��\w�,���g\9ı,O��p�rbX�'��z�9ı,O���m9ı,N�k޻ND�D ��2%��O�.L��]j�5�f��"X�%��k���9ı,O���6��bؖ'{�{Y��Kı;���ӑ,K��{7�u�hњ�\�$���r%�b'�{~�ND�,K�׽��r%�bX��}�iȖ%�bw�{�iȖ%�b_�x��u.f��ɭI.f�ӑ,K��u�k6��bX�{�p�r%�bX��^��r%�bX����m9ı,M�Dd��/~���6��f�W]	��q)��mvQ�#�8����s��\E-'dTպ��9�ݫ��T�*��1m� ��:�:۬�I��'�z�-֛v��f�MJ[�q��nٲ��L�&
�c��nhBĚ52FW4t1�p6��.�uls.��	��h���\dvsq�t�m��Nj2��D%���ZRR+����4� e��mtͭŚ����c�����Pu��!��R�fW,.,�l5�(����׳�^l�y�آ�qZ���]�s�Ql˵�w�N�!y�^O�{�s�N�X�%�ߵ�]�"X�%���ߦ�S�2%�bw����ND�,K�w�/�]:sY�.h�r%�bX��^��rbX�'�{~�ND�,K�׽��r%�bX��}�iȟ�2%���{�[ۛ�� �rwy�^B�y��_�ӑ,K��u�k6��`ؖ'{�p�r%�bX��^��r%�bX����;��+vZ�)�'w����/'��{Y��Kı;���ӑ,K�����ӑ,K�c�>�����r%�g!y=����q1n�̬v˺�����bw���"X�%�w�{�iȖ%�b~����Kı;�{�ͧ"X�����ߡ�V�16�C��ʏhu�Q�].!��.Ҍ.tg/`���+qjr�ΎEU������������N�X�%�����ӑ,K��u�k6"X�%����6��bX�'{ٿJ�c3f0kvN�;���/!y?�~��9�'�^�9�b~ ZԠb� D�1�M�L2�����&"�� 9���e02@.@�q�|0q�$L�bg����iȖ%�b{���6��bX�'~׼u�ݜ��/!y�}��H�T�m�٫��Kı>��ͧ"X�%��{�ND��"�"{����ND�,K�k���9ı,O�5�3�ɭd��3Z�35���Kı>�}�iȖ%�bw�{�iȖ%�b~���K�[�����r%�bX�������Nk3-�ND�,K�k޻ND�,K�׽v��bX�'�׽���Kı>�}�iȖ%�b}�$�%��jͶf;i�Q�fܩa������Vq�pV;rڭB���'re��i]���Kı?w^��r%�bX�t׽v��bX�'��l?�*~��,K�����r%�bX�����/MjfkSZ�֮ӑ,K������Kı>�}�iȖ%�b}�{�iȖ%�b~���O� DȖ'{�d᫖Lu�5�E�M�"X�%������iȖ%�b}�{�iȖ0���O�[*nɣ�ɩg߹I{X���Ҝ��}��F4��(d�i>�%!NlIl 0 q3��°�쓙���7���Ba��Q�p�t�SF�I�X�肚@5@7�@��I�T�v@�B~⸘�����lh2#��m�d����c&��4�|�����\����!4��ż F}�@�_�S�!O��(D��։�.2�:+�t"!��"&&�ɷ@��p^)��ϑP���z��+��E@���m�"":v��� ;J��������iȖ%�b}�f�6��bX�'���^2�#P�Vu���/!y�^O}~��r%�bX�����Kı>�}v��bX�'{�p�r%�bX���Q]��jb�rwy�^B�}�^�ND�,K����m9ı,N����Kı;�{�iȖ%�b}��^䏀�!+��f�m�4b��&��y��gA
�j�U�b`�C�����L&طi2��M�"X�%��}���Kı;���ӑ,K��u�]�"X�%���ߦӑ,K���^��d�d��3Z�3.�iȖ%�bw���"X�%���޻ND�,K���M�"X�%��u���r-�bX����za�ӧZ̖�SiȖ%�bw���ӑ,K���o�iȖ?�"dN�_��6��bX�'���M�"X�%��C�$�f�ֲfML.�5v��bX���ߦӑ,K�����m9ı,N����r%�`|80B�$$R*.�&dN����Kı=�{�m4Y���Mk5�M�"X�%��u���r%�bX���6��bX�'{�z�9ı,O���6��bX�'�{�ӓ�_,��)luf��vHL���L\R��R0vDtsa�zE��,#6���n�i�%�bX����6��bX�'{�z�9ı,O���lND�,K�����'w����/'��~�f�ȡnkZ��r%�bX����Kı?w���Kı>�}v��bX�5�g��|s�G)�r��<&�ӫcv䙚�ND�,K�{�6��bX�'���ӑ,@�,O���m9ı,N�^��r%�bX����%�\�fY5��35�iȖ%��W"w�ܿ�iȖ%�bw����ND�,K�׽v��bX�'~��m9ı,O����i�W�C5�32�6��bX�'���6��bX��(A{��i�%�bX�����ӑ,K�����m9ı���'w���>�m��+�6�⫗ JvoI�;sj�;�+�GK=����/mu��gp�8D���r!>�lW>��Q�Ȗ3V�X6���,�9竮��ݜ����E�����7i|E�I�rum�t�m�4��7A7V�vM�z����(�m'e�m�NUȪ��i2f3�Ja�$gf��`�f��4����5�]���e6�*�J�R��h�R��AΏ���� m�9,3�,�FL%m�[�,�]��:M��4�l*K��jG�$�������޹<���/%�����9ı,N���m9ı,N�^�fӑ,K���ߦӑ,K^O~�諒�3�ڷA�:�����bw�o�i�bX�'{�g�iȖ%�b{�ߦӑ,K��u�]� ����/'�}��+vZ���N�!ı;�{=�ND�,K���6��c�0L��=�]�"X�%�����M���^B���>�k�M	�͖!�t��bX�'���m9ı,N�^��r%�bX�����r%�b�'{5�rwy�^B�y���R�f��*��ӑ,K�����ӑ,K�}����Kı;���m9ı,Ow���r%�bX���vx���e�)-S���	�mnm�4�,FFl��,�3Ee��.�b8�LآӢ�p�c�w���oq�{�o�iȖ%�bw����r%�bX��w�9ı,O��z�9ı-��߃���-�3c7�N�!y�bw�^��r q~% ��0+�� ~r%�bs���ND�,K�k��iȖ%�b{�o�iȖ%�b~���|�Ff]��N�!y�^O���M�"X�%��u�]�"X��b{�o�iȖ%�bw���ӑ,K��wž�d��iֳ%���r%�d��}�&��	ｯM� �'�N�I�$�z'���m9ı,O�x��.�V�ɩ��f�ӑ,K���ߦӑ,K��g�ͧ"X�%���~�ND�,K��޻ND�,K��ޒ]c���fO�NY�Sن�k4�[7m6�m)�kK�1����}<�x:�YkEV���d�,Kޟ���r%�bX��w��Kı>��9ı,O}��m9y�^B�y����К,�bQz��%�bX��w��Kı>���Kı=����Kı;��si�$/!y��t G,���z�Ȗ%�b}�{�iȖ%�b{�{�iȖ;�����*�)"X��׽v��bX�'���6��b���y���]T֚��'\��B�,O}�z�9ı,N�k޻ND�,K���6��bXb}�{�iȅ�/!y>��}�XmV뙊m��N�ı;ٯz�9ı,�{�M�"X�%��u�]�"X�%�����ӻ�^B�����)x]����3g��Y|��N�-ã"R0�K��ƖU��x��f�,�WE֡��d���ND�,K���6��bX�'�׽v��bX�'�k޻��~��,Kޚ���ND�,K9��1�i��.�����/!y���޻NDı?{^��r%�bX����6��bX�'{��m9ı���}���B�[��rwy�^'�k޻ND�,K��ߦӑ,�,N����r%�bX�w^��r%�^B�}��i���n�We:�������ޟ���ND�,K����ӑ,K�����ӑ,K@x���� o�5�{�iȖ%�bw�=g\)��fkF�����Kı;���iȖ%�b��u�]�"X�%�����ӑ,K��g���Kı;�I}�41�+����na-�5�k�����Bw9a���qvcqQ�{�w�N���i�Xc�Z��r%�bX�w^��r%�bX���z�9ı,N�k޻�B~��,K����ӑ,K��}��n�Mk&��̳3WiȖ%�b~����?�b"X������r%�bX����6��bX�'�׽v����0r&D�?}���F]��s1M�u���/!y�ޚ���ND�,K���6��bX�'�׽v��bX�'�k޻ND�,K9?��>��D�[2�n��'w����G"{����r%�bX�����ӑ,K���{�iȖ%��,r'�7��v��!y�^C�L~5�:ǋ��rr%�bX�w^��r%�bXG���]��%�b{�_��iȖ%�bw�ߦӑ,K����:2$��B DFT
`"")"�����s�~�m�b�hT��PNӠ8a�,6�Q�\.↭��*��1�F]t�Ke�X&������ųcg�vAp��-ɮ>!^8v�;73��>�% �{s�ؓ���L/"'<s���N����!�<��	�k�j\g����[v�1L�.�Sa�����s>˝�g����;��C�M���GjP4�3pj(hA�F���<Vi��<�.�-�;��s�5���If��[&j2�'8[�;vT�%"ۦ��u���8�T3�s rL��2E�������vN�;���/!y=����'"X�%���{�iȖ%�bw�ߦӑ,K�����ӑ,K���OL�m4Ye�L�f�v��bX�'{=�M�!�"dK����ӑ,K����v��bX�'�k޻ND�,K���r�͖ۢ%3z��������{�M�"X�%��u�]�"X�%�����ӑ,K��g���Kı�}>�b���ܙ%Uo\��B�HD����ӑ,K���{�iȖ%�bw����r%�` Ȟ���6��^B���~��
E�&��]�u���bX�'�k޻ND�,K��ߦӑ,K��{�M�"X�%��u�]�'!y�^O����K�ò�h]G��%����x��c�W��
�{IY��Y���WD̙�3D���]�"X�%���o�iȖ%�bw�ߦӑ,K�������c�&D�,O����v��bX�ry?D���h-�Mi��'w����;���i�m�|��h;dK�׵�]�"X�%����]�"X�%���o�i�6%�b^��_fd4�Y��jm9ı,O��z�9ı,O�׽v��c�$2&D�����ӑ,K������Kı>�=�I�Z�e�F�Y��ND�,K���]�"X�%���{�iȖ%�bw�ߦӑ,K �>���Kı=�V��,�e�53Y���r%�bX��׽v��bX��������ı,N�_��iȖ%�b~����Kı=������>f���hK(�I��t$��1.[��ٛ�Y�+�2N�����sm&�v��j�9ı,N����Kı>���Kı?{^��r%�bX��ND�,K�=�Y�e�Z�5I��h�r%�bX�w^��r X�%���ߦӑ,K��f���Kı;���Ӑ[ı>��u����T�W5u���Kı?{���r%�bX��ND��� �F1�B,"0���P�`�#)$H��*lM&�{����Kı>����ӑ,K��}/�5��Lѓ4L.\��r%�g�C"{ۿ�ٴ�Kı=�o�m9ı,O��z�9İ?�D�����iȖ%����~����D�[2�q��'w���%���~�ND�,K��z�9ı,O���6��bX�'{��fӑ�^B�{�e~�
0
�w1�c�Jv�z�n5(��/U��앃+FSPްK���zx6��@�lb�Ao\��B����z���D�,K���M�"X�%���{�iȖ%�bw�ߦӑ,K�����om1�vN�;���/!y?����I�+2&D�=����Kı=�o�m9ı,O��z�9ı,O{վ8�4Ye�L�kZ�ND�,K����ӑ,K��u�]�"X� �2&D���v��bX�'�����NNB�����{���il�.��'q,KR��u�]�"X�%��u�]�"X�%���ߦӑ,K�� � 6� 4�1"��b���M��iȖ%�b}���[y��kR�3Y�]�"X�%��u�]�"X�%�������i�%�bX������r%�bX����Kı>���>NYC��mfZ]un��R[��2���]�]נ��G��5n/8�]���BG=�g��Kı?{���r%�bX��׽v��bX�'{���TC�,K��{�ͧ"X�%���]�SRf[�%ԘL����Kı=�z�9Q,K��u�]�"X�%�����ND�,K���M�"TȖ'�Mg�d�W,֡u��35v��bX�'��]�"X�%�����ND����ߦӑ,K������Kı/���Jh�1v���N�!y���K&��fӑ,K������"X�%��M{�iȖ%�-��뾻ND�,�/'�Y��˻n˶xL������b{�o�iȖ%�b{�^��r%�bX��w��Kı;���iȖ%�b|���<H�`Y��Z��F4%B��W{@����	H1`c
	%%���P�S�hcL`5�8�jAA>�$�0".��SBp�dWih��!���=Ԃ�a�C��>�͂s��57� �ăE��<���ت��������UU\�UUU�U@v�UUP
�V�UU]UUR����������n+B!���c����vMi��d�toj�*W˞�P�sl�p���vƁwb��v90��	���;e�\�Ȅ���(��v����,���sEޥ�<jf7�v��.[�����crqM�t���vIx-@��#�pb3^Xq�-g�`��3ۘ��$/P�:f���\o`�,T���؍��<%�Ƀ�nչg�OS/R�8�\On��'`��%闗=dƝlc����mkxD Ǯ���d��6Ȼ��WK ��UF�Wm�]:����U�VZI늻U/��\�ݎ:����$,�:6���k�h��f�Ě	#,6m�c�fV��� ���uy�i�ʵ�pf3Ӟ'����	�x�v,���w3�l�����C���8/jX������6�K�BhGJ:�.y�4fls�2ƖE�:%*RX�Ss�:Vm�zL��M�j��Gn��k�RP'g�=�<�ݹ#&�Z��.y�s�9���6��G�����52�r!�dc%խ�p��ؤ�Xq�L>����r�����x�r�ñ�mi���D���[u���,M͚y����'9+-�V��c��Xf��*�-�1Wl�n�vӇ��0�nӜ�{,��=��P[Ⱥ�=u;b,��tQq65�35#[UqI��(VXsh�8<s�n�Q���A��T<�z,�X��ԑў\��(r�4	]���!`\��Xm�U	K6 �7c$l;[�7:ѺvN8��mm�nsnҙ���݀;wd2�A�q����5���]ەY(,�D2���&%��ЩQm�j�Ie��h��a+gf%�*j�*�/4/��ɶxn�����/�+�ZIOmt�x�U�L�u�mIDjYj�P���t�.��@W����X�r;qk*�g�v4娕Y^���7�R5؊f헧�x}đ����]�.F�@����$�fܥ2��'$����9'>P ЇGH=AB��&�'>>�T~D�� �A@b��p5Sj��%��֪�'OJ�UU:ՙy���.��N��rAo�C؅��"8㓗�āә�x (��3n�;nnԛl��qh�[�xn.{vXŻu<Xd��]�ֺ�tڬC��te�4���J�()�i�9�@����[2��{\�dO#+۶ݧ���;J\�iC(�p��.�:n�ϧ��\i|�:�e�Յ��`,BXk�m	��-[�#�Y�社��`S-�خh�0���b��m�)E	��V(�a.n�\eB}�I��)XR��U�p�Kı=�׽v��bX�'���m9ı,N���)�"X�'���6��bX�'�����Va+�sWVfj�9ı,Ow���r%�bX��{ٴ�Kı=����Kı=�z�9,K����am�ճZ�5I�ֵ6��bX�'s��m9ı,O}�z�9ı,Ozk޻ND�,K���6��bX�'�����Z�Y5M��n�Y��K�,O}�z�9ı,Ozk޻ND�,K���6��bX-�����ND�,K����j�2]3Ra�3WiȖ%�b{�^��r%�bX��w��Kı?w^��r%�bX��^��r%�bX���C����!�r�dZ΍�0x�&M	zY49�͛R�."��y>�=Z~��<V�e��r%�bX��w��Kı?w^��r%�bX��^���L�bX���~:�������=��k���-�S�SiȖ%�b~���1> ��U$VAF
 �i+��%���ܻND�,K�Mw�iȖ%�b{�ߦӑ?�*dK����$��96�m��N�!y�^O޿�rwı,N�k��ND�ı=���iȖ%�b~���Kı/��ߣ)XR���N�;���/!y=���m9ı,N����r%�bX���z�9ı���{�iȖ%�b{���b])ŘQ�d듻�^B���}ߦӑ,K�O�׽v��bX�'�k޻ND�,K���ӑ,K���N���ckvv,a�gŖ&���)���E
�2��[���rh��`�5a��fr�9H�#��v?y|}�� �7���'?rrk~���������
�ꑊ�]�k �G�\�+��D��,H�um���_��@�O~��Hl�).2`<��p���EK��ʪ�*�@!��������_���ܓ��]���?��z�D�[2�n�տ���No��ߌ}�,�0��, �ʻR�+�ʺm]$ـ}�"�=��r��g�����n����U(���m*�a�Ls�m�˝�����l�%��a���uvn�ZG@6q�tæ\��޽8���p�*��|������#�������X�{~���r���{��o���}.E���#}<���\n�6��m`G� �nE��r����������p{���5����p?גO"��w��,���v�Y]��/UW6�� �H�� �1��[������������0�g��c��M[.�}.E�}�8`��}����{��*�DuqI`��u�e���a(�RQ��YV]�a4K��"D+i���gZ�-���:-�P����?w\0�{�܋ ���,j�6U�e�ـwu�=ʮr�#�s� �y`n�N }ޘ��)4[��p�wݼ��9�%�� ��B��.�U�WV;�n��>ۑ`n�w\0=�r�u�, ����'J�HB�[v��>�0�`v�,� ��'?�<�-���UF�m�j��%6��H���n ��l�R��\1>lT�Q��뱯�QX�R�k�ѱҪhV��^�m˭ka'���R�r�XW�fs��S�3Ԁ�R���qӣjyL�v��U�.:;t��I��3㴝�.��5�B;fY�nPe�h�v�v6���5k��=a�l�A�c)mXKx$/g]3gv	�xyl=��z?��?ۅ��K�fe�����t�%��59)�e�"�°��:M=���\n�[T:�|��`v�,������?��{�^��~���n�[��\�f�ob�>ۑ`wi� ��~�~�������U����e:������ۣ�s�wn�{��픑t+B�V0�/�L����}�ذ��X��le�j鱖��E� ����_�~��>�0�Q��Ń-Y���2�[e�r�+�V�\Z��8�0�
e�6�MC)�?��u`mȰ�GW�6G� ��� �:�ƚ�e�շ�7��NI�y4�ӑ�WgoGw\0��g��~�߿*�buwN���&�{�� ���������j�.7V��h�`~�+��s���o�?��܋ ��� �knR.�h-��m� �k��s����$��wu� �=PY^�B���vU�m������6|�})�q]1۳f]{s{M����p��������߿^��������;��`�^OͫJ���T
��7tp�ԑ�?��� �nE��U�]�_�=����le���l�'��eȰ|���h��\�s���H�$�%���9Eer�]v��W��� ��������mV���o��$<���o���d0?s�d��W�@]��]Xk �nE�~�s����>d~0{���=�B��;x�CbQ��G����$�,Ra�P���X-�zSɱk)+/-�,�Wl��&���	����ۑ~�r�U_ ���x����\n�[T�l�7u� �r,�$�H8g��I$����ߥ4V�f�eS�~����^6S�����X�c���l���W*��v��^��~2I��k�rv�Ad`��$����"�b:P �.f�۹'O�n�j��n�i*ۼl����?Ur���ߎ������>RK�"��%P��m�l5w�c�L6)eٖ}��,�;#re��/AJݦF�l���:��8�|��&܋ �I/�U_ ��?��u�v+*�t�f�r,�$�vS�����\���U]����w�[�uc�n�_�~�IN~�r��?����	"�iҶI[V��~�R��0	#�E$�ܪ]�{׀M��X4]��V�4[0�p�=��9U���?߿_@�����&�� �r��G9\�R1`H�Ed�@��y����݉��4#m�l2�^�ɟ���+�;kh�a޹�z�
E�k��ܤ����S6�y�\�C0rcjU����Kb�4�X0o��1�ر�Ǜ�2�i\S��[�vҷi��5�[�VT�R���oX�{��Q�u��h4x�K��v@�T���b�a�%�U�@!�#�e�A��X�K!Z�6QpIC�6SV��]k���NOxG��O���ֹ�-��rWF$�)����,n:y�Mm�u�����$��gˢ��!�O@�~���׽��M�������=��/Xۺv4ح�]��>RK�ܮ$zx~0۞X[���p/�χ�1�$��������;�ذ���|�%�T�(�	�m�J�l�;�ذ���|�%�`����]+*�i;k �l���/ �����ŀn�#��ѥ�,�$��	��;��ٺ��v�b����(\��tɿd� ��v4à������ �����ŀE6^ vE(�ҷBBV�jۼv���H�$d$�SF���
��������>]���+�ʪH�������e�j�-���,)%�.�x�8`����v��]�wm�)%�.�x�8`{��Urg�,����WGTZ/.�����ﻫo�rI%zx��s� �Ix�U�݋=j�i䩲� ����уm��s�;Exܲ��A�K��hx�߸��/�U��F;=���w��`I/�+� ��z�ϵ�|�A¤Ì\ޭ����N�r�{޼�}��&�� ;!ujZ�2�t�f�����ڪ�s꯬�)�U&ɒj���޴!$	p9�u\��|ʬ�o�+t���͕��a��AB`��3�,(�q(�
���̪M�̹��3z�t!v�٭��I�  ��3��1	�s���~@����-B1���OƃBd���J��"V���M&R�m�%܋ȵ�ZbH A�BHŒH�e�aHRVVR�VY%%e��¬�U0p��0��c�B,HH��� P2�B��-��!6�Ke+HJ!)B�>3@��D�!J�Th�,]R@��f�	c�±�!,c�R�hĐ�
0!�4}$Ŧ��5IrI@�eeIIIH%���%@�F4�LU)I��
`�@��ư`��Ȑ�i�d�ڐ b� P�BB��4��Y4Ł!eP�ŃGI�%a��	!7 ��`B�����А��� � ?��@b"��|�'V(~A�~>�<V~@�)��b���`c�!Rycv]X����_�߯ ����`��E$� �)E����+V��`�{�L��^�� �l��N��K/Q��gsuj�iN'���hckRo���8���F�.����Pc͑����cd~0���|�����A����=�ߥ4V�fY�' ��{��y'�KOT�� ���`�p���=��%��lM�w�u{޼l0�p�"�^7�8ڻ�l��
�����^��7$��צ䝽�sr��TJ1h�`:48�T�hC?_��܇��^�3Jꭚ��,���Ӏv�/ �l��M���?Ur���YBS����+s�#.f�,���^�T�͕���G����Բ�k4�OH�N�j�V9ˠ~_�~��^6+ ��ŀHT�.���.�n����^{��RG��e`.y`I/?W9I��^��Jؕ
��6� ����{���Iy{޼����l��bWE��jڦ���8�s� ���x�Ix�U�s��ߏݬ��^�ԋ��umմ��"�^�^6+ ݽ� [�)
��V�r[�'?R|ݪ�ٌZ�nW�b�l��p���N1I`�NR^W�u�$�����8��� b�D%l3Q�<��.��{�<�������n$�W�3���6ي�9&��8��,`Z�,`fh:Z�i��8΍��K��m��s��I�q�- p6[�z5l��mc���i�sfw��,�ca-�e�dr�;v����Y�V8F���˙��ԑ�{޽����Ӻ�lKhM���������z�]q.<-����3���a�0�����!�`u2�m������׀M���7u��Ur�A��z�Ny?6���(�B�]��&�e`��E$��$��UW+���ʜ��?j~���R`M�έ�}���B)%�����W���=<{+ ; ��J�t˱�V�0?UUr��~�� ���x�L�w\0	
���X݅մ�$��)%��UUr�<{��	#�E;��?�&���^���T6����f.2F2�2�1Z�UM�]s���۩�^�Ő�l��e�m�6+ ��)%���:��^��	cJ�-��Ҧ�� ߾�f��Bn\"H@���c�k!R!-T�HX[F�jK�����p8������;��~���p&�e`K�)�h-�m�]� �Ix�Ix{�ʪK�ǲ�	#�Iq
Rn鱻i7����.߽��=<{+ ����U/_���=9���v�����+�x�L��W$���<��x�Ix�
�����R�:t�u�Ͷ�n^%/E(I�.�GS��)퇝Ɇή���Ui5v7X�`l��|������=�����h�:av1զ�.��$�n�+ ���U${�{�w�݅մ�+n��{׀O��ٸ)�ȁ+ ����je�X��-,��+�.�m[w�ꪥ$=�`\��>��`~�UUR��޼���X�wW�e�t��ـn�ŀz��<������8`�=(�Xxa��&:ɜ��]n���>L�T�Y�bU'��9v�ԫ��:�u���sj]_�,�$�wGv�,K�Q�ln�M���|����$I� �����?q#|W��]۲�hT+�x�~0�ذ�Ļ�XW���%KIH'N�m��2�`��`Kذ���>����UJ���UXe��kc-���0��"C�� ���u)� ��i����۷f�M�2�Gy�J���c����v:t]�WV��{���{��A��7u�ryym����ԁ�2�SF�֛�+<�dk�t�D[�1�;q�S�tF�햠��:����u{޼wGw\0��X���X
خ�e�m��������,�$����W��߿ �ң���WJ�����>�с�wo ���N'M�t�cWl�>��`)%��8`yI3��_����64�n�V��^�����+ �s���4�� `��`?����UX�ͶAU�9�H�܃�q��9P�gu\x8��n*��K^Í���m������#ٯ^�����)�]��e��a��\4E*�le���v�d�4v�D"�d�H�fn��".�Cin%����Tږ	����v#a�K�0�QF<�M V�<�p��N�)mRT%�dJ{e�Fi�͚��n��u�{g�^6t�f�W7d�\VZd������{�N��~FZi�Z�T0�̈́�LXvh��sW=h\l��yttv��5�3�Vwi1B�w�;�0ݙX��,�$�R�R	�WM�V&]��wfV��� �I/ ���?RA����+C`]���n����^�����y8zN�ۉ�Y�����$�����x�~0�̬�{6R��"���[V���8`ݙX��,�6^ M�*�P��W�C��ȱ�Ͳ��,��䧙��U�,���n8A�J���4\�d�{�y8�w�X�Ix���qJi�[�۹�f�nI��ݻ�(��,��w6��̬K�(�li�7LV��^����UUq-��X}s� ���c��vP�
�m�����ٕ�}/b�>[%���n��m��2�`ݙX��,�^�����*��(�z�WC��47$����g,��M��,�vx��E��p�붥r���E!��l��=������{��wfV!R�Ֆ���Z���^�����+ �^ŀn�R��]�]ݫbi[�wI��n�ݛ����`���T-Y�0)b|�b����,a�*����()#X�P�8D�#h�3��n�I���7$�HZX�;�˧v�顺�7ve`Kذ���S�SM	[�۲ݷXe�X�Ix�\K �ٕ�}�ҽ4��\X8k*���½�ͳ��	��57>��۷O���4����Ebt�m`-���ٕ�������;�~��v�Hl�U��~{o?r�6Oe`�X�r,�+��H�/�&�%t�Ubb�i`'���ذ�UĽ�~0	��, �u*����c,.�`��`�� ��`,�YJ��"=�@\�\ü�}�&�����Z����V��'c����&���;/b�&�) �����U��P���8�R$2��[�Z^j�چ\N���q�x�4�ٛL٦�4ML�����uCwfV�{�s�������M�.�l����p�;/b�>�� ��g� �����J�ݖ�ـI�� �G�\K ��K�KI�M�6&�ڶ`*�}��o��X�`~R{<`�I���`&ں��0�q,n�`�� ���S���:0wF]7���{���k����Û�~�o�!;$"W�of��_��:&��""!at��_���XS�$#!�a Isf�_�F��a��_��^�Z��E-@IH~�1L@��!���j��/���L��ŌIHF���Η|���kW_���\�˚S�kJ? lL/1��Č�'�o3{�A���5�5�44������;pm��JH$` $&��� �	��HŅ��@�������z|�D�Ո/�d�C?]�2�$(JV�."��@��0����0%��$�|����
m�T��޴͑bHM����I��Ĕ I�~Ӡ� �Z1�.q��`cKFI��}�)��$a#I�)!!����6�T���#"H�e���˄.K��.�Ho��l��B<!��:<��ت�����������m�UUAv� +*��V������
ꪪ���������bw\<���;v��g�Qtg7\�L�J��ۍ��� ���l���콵���v�1� �.�=vL�۴�vF,�X��2�jke%��%qk��F�]�l@<Qŵ�9�g]t;1�WF�D��5&�4�j��B��۵�j4��C`GA2�n�4�hRf8jT-�\$v�Cb	e@��)s��f<�*ی�Hg�:�ix�7�c$8a�Pfȼ	��8�Uf�l���;d:��R¥��t�c�Ws�=3�H�Ôcv���B3BY΃.���kv���U�9�ƚI���g�jxdm+�Ÿ��p�J3��:��qy	�4�D�w���Ñ�';-N��f��S���6_.�u�i3F�ڰ�]4����+YKm@\��vm&J�яr#�fN6ݑ6bُu�h�`�=r�gs���T�z	6�N����������S\s�Gl���	������`�ֶ�F+��U�eY�`:����{TRt��Y�h�^R�N�T�w/0Fpˢ\��g-mN�;֟rnk@�CXV1S�M��"��ImŽ��&�m˻s�#��A��\�̡��Z��4���6�+���H弩�-�h	�ٹ�(O��;Te�g\��ݬ��+��<8:�cmu�+�ZL�5Ф����YA�(�m��nA�,KR���8lŧ��nL�s)�!k��^³��OI;vg�I��α�3ٻ(� V-��w�M����5Y�+Y:�l�;�`������R`D�v��*vU͐��qa�ݗ�]Yats�Y�"�2�I0@H�+��d]��@�!�"T��7S�5Ap5<i���Q�bp�nq�3;��x�f�K����:�9�p��j�c�a,�1t2�z:z��9�ۢ�py��<�>Yt���I&�y���mp�A��(nP1�enQ��Y�£.6J���`&�����eW��6�D1�	�8��U�tMt@�D�9�O�G@E�tU
� �h�=*~D8a�@�:uL��ff~ֵ��334ꩬflqȨt�'j�l1�jڊO>Xݠ�\n����+�<�ήCM�vrt�M��n9�Z��R��ڃ�칌�i�xnyu��F���b�cOEV�6.Ln��ԽM���*����V�Pr�uGc���v��K���y$�Ţ�ryM�%@� [hR�;��q�\�R�b���Ap��Lm��b�OKu2�n˪Z�;�'9ɣr:���f�Ŏ�*�1���,�2�'���t"�[(m�%̳AZ֌Sf�-�Dֶ���>�� ��0	������� wb,<��v2��0��N��\K �{!�Wyn�����ճ ��f��6�,v8`��-,��+�]Ӻ�l�;5İ	��`��`~^�g���a����Ӻ�J�M�� �U[�<���� ��`�sa��aL[�i��Y8-���(�H��T�K:�I�T�]��0���V�ݒ�C�o�y`�� ��{�ʪ��=.y`��z�m1��t�m`��7�� |�B�f���w.��>�ܓ��,v!�1]�m��M� ��-`ob�;/b�'c�)BTm�I�c-&����&�ŀv^ŀN�v�]���XEt�X���;/b�=�o���M���&�ŀn�#g��F��7h]ͣÖ-3��c��h8Z� 
e����7e\�7<��.V�v8`�dX�ؽ\�s���,OW��e]�]�WMU�f��E�M�� �^ŀN��QD�)�];�T�ư�����a+9UڮQʪ��@B)�J���"�b�������9�ڑ`��`�n�V�bn�=�U.�g���{�����g� ������cM6&�l�'u� ��"�"���>��w�9j�MYNӦ]�[Z�;SI/�l���ב_m�ݛ��9��]���`&ں��0�,.���`���v�'M��WcX]�y�s��$w���=���7�Ȱ���M��e�ۼ��aꪤ�D�`[=x�!ww��ut��'Wm� ��{�]�{���ȨAB����&�w㹑WlWj��Ujـou� ��/ �k�;��!��X�|,�	kR�[�\+1�XS�':̎�j �_mm!�b��uj��>�g� �k�;��\0IJ0O���7x�\3�q#��l~0���ԑ�_��wN�|wl�=���'u�s�yl����`�@eݻ�6�զـN�;{;�+ ���{ٺ���[5u6N�wݼ�ٕ�N�;��P6]��M��6����p&�cj�X���৚�yX6�P����qƶ�=�X^��zXm�q�P�;���N����7N|�8"ݷ�Ey���;�4@TX�z�ŉ��b0F�12F����F��y�\q�Fދ��j��Y4ui��QÈi���K}�6���y��
��V�:��I����Ua��[�jݭ��y�Rʤ\�to�ګ0����YA��)*!.���9^f���9�p�3Է�h�;1�A��6��p�v�.��ʰ���}��N�w\0	�p�6BU��t���t�+v� ��w\0�Ȱ	ݙY���U$l�z�FU�.�t�]� ��� �܋ �ٕ�vk��$-*1�.��E�0�Ȱ	ݙXf�`����t'��Ю�m&��ٕ�vk���{r,ܮU{|,�4��y�%���i���9z�"��:{4�l[�b��%YS ʹ�j�ƫ;�����v�/s���ag��5��W]5T���<a燐�_�"B   ���`
i���%�;��I��ݛ��=8���u��b�j�l��� �ٕ�N�;��uZ]:t;V[��	ݙX�`u� ����zvm�Yr��Ys��;�`u� ��� ��+ �J�%�o����r��gJ%���v�]K�u�F��n��4f�؂:\k���z9}�w\0	�ذ	ݙX�`]�
/(b�]'il�'ob�s�T����=���'u� $����ۡ]�ݺ�ܓ�����;��vnaE�	�ł�HT��"y�4��� ��E�J��J����m� ����;{�u� �(iݦ&˺�m���v�,�� N�x�
�
��4�4�n�I��=�mZ'��HR�E��<���[�c� �*������;����{�Ӏ��� }���N��U�����$e�>�p�7����lۗK�4Z�ܜ ����������`w\0�v�Ytբ��H�o�]ٞ0m�,��*�h�Us8�T 5���[�t�N���jR�.��V�v�,�� �������{����ԆB�4�ȑ��۬�S=j0�P�O!�"�6�1���-�[m������� 'v<�뇫��W�?}������� ��\��	ݏ ���N�ŀ}�ذ�q��݅�]�v��>�`��`v�, ���	J"GMli����^�<���, �������WD.��ʲݵ�}�ذwc�>�8}�v���cnꪱk�h흪�Ӻ`�-K��/*��T���]^#ėZ�R��,_��r�mD&��M��:6�t�ʳ�V�-l��q��T-V�ft5�H<�xô#s��ъ�^�'�ǃ�1'��X6m�Z�=�ڕ��ѽ��N�iFb��-XK,����԰ŵ�%3�!*���b!We��`���R�E��aq0L6ҙ��2K�X��j����d&�w7u��%�*�ݡ��#�M���5�K�V��n0��;;�+���β��;7����{�ӀN����_ ����6{ԯ��V�˦�v��u� ��� ���`�Ǟ�$z�E%���I�E�0m�,���W=�� ��� $�J:I�]��ݥm`w\0wc�>�`��`F�(n�66&�ݶ�wc�>�`��`v�,miIԫ�*��Yh %.�`�4���Kۮ�������-�8ljP��+F��m��w\0	�ذ�{ N�x�/�B����8}�v�y/��BD2�dHH� �U"�1AN�� >Q�l�~��.����w\3ܤ��%tx�lc*�v�ݹ���u� ��� �	wx��Ln��k�ʤ��� ��� ��� ���`�|XMZ�.�E�x��v�,�� N�}[~�>���+NjT��̈́.��6���]���O3.)T8���n',�ǋ��.n�"�;H�g�{ny`w\0wc�>�`�)GI>+�B������� N�x��v�,HХ��Cn��� �����eIo8��0�!���	��3M�����6C�㔉R&a�'j�R[�# �!r]�L5ie��g��RRXI7Kd�۰�����! �A��q�$� @~�k��$e�9����Ϳ���pk������jI��Sh���J;�B!��Nr�g�$SD4���K���͒)h}����7��ӌ���Zʖ�>Wg>x���?|*+�=�� |��b'�� �'Qq@��U]R�*���s:�v��p�;��i�m�]�v��>�`we�w\0wc�%(�phI���1l�"���>�`�ǀ}�p�=UT���K~��F]��mvVl�a�BT6D]elT���8e�@m�ۣf���[w���`�ǀ}�p�9\���^=��w��[at���l�	ݏ=ʪH��� ����>�`�*��Ue�H�o ���Eݗ�}�p�	ݏ ��*�YM��tՎ�l��s�K׳׀wc�������uW9T����`�RET�b�*�
T��^�7@滚�ܒsǬ�N�v�N��V� ���{��^�����`we�+D�%v*�IX	�u�<�0lg���]ؽ@4V��K=�i��\e�+�(�Yr� ;��x����"���>�p�;��Z�馂�.�m��g�ʤ�-����� 'wׯ�$��>)��PZ큰ٽZyl��v8a�${g��� �t�wM	0���޽8�~��;�p�"���$���O���7V�f vlx{���xݎʕiB�h~XP�(-�2(�),Z��*A�k�˹�;�kZ�h��VڪD�ssuyoL6��YT�jXC6	���ut;Cl8*(�qڷb�

;i�x�ѱ5<��n<NftK@(i�1e��DFӕ�(<[;��Q�d��1fb��)�˹�n .��E�֫)��̘��Bz����t�<�[]5
�'`�13�z۱ջoW	E��2b���Z�2n:�Q��tf[n�콖�۳dzs��]f2f��� =9��L��k���%X��^����U�+���ǚ�&�jQ�k3n�Lh�f2P�~l~0����0wc�;�ZU�tq�N�J���Xݎ;����Ӏt�:��0��[��>��X;��w\0�����J����+�k�+�w}�wc�uwe�v�,�k�wI���wBm����ݗ�}�ذ�����~��k$ny����糓�yM�ݍnv�ZnQKn��r��tcN�s�05��\k+�`]�xݽ� >��\�|��� {��t�����\�������HX�A��Az����ܓ����/ ���>+l.��[m� ��<���%�g� ����;�]��e"鈻��=\�R���j���>��X�dx�ڕb����t��]� ����>��X�dx���R����*R��������9�ڭV�;(�t�E�h�*�<�5s8�vN��V� ���`ݑ�w\=U�s� ճ׀Oy�z��Cc��J����#�Ur�����V�^�nE��9\��d���*L-Л.�M��I�����ﻛ��B!$�2� ��"�,#$�T 1�E�����y�A-��;i�݉�]���UR����;��, ��<�� �A]K��L��7n��r,�.��v?Wv^��#�J�.��6W���N���x��`�F4W!�z'�gnէNgpEma�ƻ9��fU������;�p�:����r,�FӲ�|i]�x{��r���5l����� }�{���G|O�e]����`�z��r, ��<��i2�؋�$������~���ߖ }���nI����ܐ``~ �D{���]f�+bȩX�A��ł8@�
0 ��&D'�y䏞H���n�z���Q��]�X�dx�ݙ��5l��v�\�{^�눵��U��0fy���6cư�ik�Raa�f�x�h���' ֳ�+m�.�.�M�����:����r, ��< Лr��]ؚE�0���܋ >� �u� >�WR�����xݹ }��U\��\�]����"��xʒ��|V�]1���X�dx{�Wv^��u�� ��]ZJ����|v����ܪ�\�G=�����`ݑ���9�6؁�"X�G�{�ff�&�rq�����씧�+��[�q��;�S]۝���"JO8xk��gt���p�Lʥ��E"KU0��Y��9��2�T[kg��Q���q27F��(CM���0���}q�v�,�r�g��>�욢T�hy��4�%��[w�f�tc<�m�"�B���]���v��\]���D�4L�m�Kv�n�/�ƙC��Hnw	�����<���9��T��N�B)���V�=�'����B�[��NF��+�sA�ږTP֌��XԦ������7 ��v, ��?�9\�U|�v?��{*ݥWm	'wE�xݹz�ʪ���U�o���y�0���	�Х[M��n�j���c�;�p��c�>��X��K�wE�.�.�M��}�p��c�>��X�R[�� *{��N�uw`����dxݽ� ;ݏ ����=�!o�B��6�y��[5�{>�9,�d��7��ۙ��P4�Gk2�Y�ͭ���m[x�� �dx��W>@l�x�{֯���մـl�>�ڮs�ʣ����a��0wc�>�g�s��'��V���W�j�wc�ݏ�T�v?��<�ڕiWG豗l��\�%�y�۞X���=��R���{O#�V�*��I��
��>��X����������s�>�S�#��q[�c�5E��NE�q�v����V�Ů�U��V~�m:�X��V�] �~�������|�߷D�o�v��a�mԮ^��р}���>��X��y��DT{֫�v[�դһf vO<��v����Q"�Aՙ����?}��7$��feK���v2��m�w\0������_�ʻ�{��=��~�x��M�Vճ >����<|�y�w\0�Rސ;dvb���Tn�`�W��H���X+r]j�4gѭ�m\��#�i�_����u� ;��u� >ݏ �6�Z��tpwCil��c��ʪH��� ;'��u�?r�;�z��'iU��N�Z���~0�������x��Jm[�E�B�l���q.�y���`wc���US��W
�P����"�v���w�r�I�K�t�:Wm+����������{ }�< �t���ڧƮƑnK��k��ڡKh�%��M�Lѹ0�aw\��V�6�uB��Y�m����^���� >�����U��������ut��U�����ŀM� ���ݏ �RZ�O����ݵ�M� ��ᇹĉ�� ����6Iuj՗�;)_�v��u� 7��ob��ǀvR�#*����]� 7��ob��ǀ}�p�%�mUWB�k��74h3�ǕLf����(�^�|�U!L�O�>!C^ஔ>w�8l�`��-�$�������VJ@� ����	L�	;��?�w���sD����,���I���P) �1&��ǀ�;�D�7��6F�BXQ�� F�����&BSHș�m0��""������@�Eֻ4.�v�]!���?8�ϥ4o���%��~A����)��
��p!#c�?F�C���X~/��m�۬�����%ϳ��)�>�CJ(JJ��!`H�X≠��x~�S�z��Q�䤬�d�}@�����hŠO��.�#+JbT�ĥjW4����y����K���uG��m�y��(AUUUUPUUUUUU��UUT�
�UUUU���*��UUUUUUb�i������yZF�9Nыn��z\
���lGKN�vZ��ۧ�l����gf��:-�vN��m���#��#m�_6��#R:�)Z�M ;q]�ćE#0O�99,��A�2��Ɨ���zU�s��4�F {u5��A0�h�B���tx��l3.f�<��>v�.�T�cJBSm�v�s7�U���Vcy8�`=0]���KۦT҂`���u�N9ױr��R�[c�-]�q�<��jud�8�|��ݷ(C�Lvݒ�(�givp�HJ���<�@kd����qk�35��!�-��X6����pۦT����B]ۙi+h쵻>Xޢ�����L��T�fc �D���\<��7�Ź{l���;�ta���5c�t������jom���sEc����y���뛅{@��kdv<m,��)�b���4�p�Ym��H\k�n�R�V�ZL��#�%.�#�u���m�@�է�C�ƹ7Tl�����l2�r�p�esp��S':x:i͢�TV��^�b�j�Ko��7�k���Q��v�-X2%��֝R�U�<��̙S^��M�&�ָ��t�m�c+qc�C�Z5��FV5�+#s��lm�q� ��M�lF\�����M�U�dKݞyr�Z���B�Y�l���^�3��ҺsE*kaY�k�H�m�^MK�Ub�,ᨺGa��]+�PW�=��m�gٶ�oO]p�jU�fiu�Meb�t�����G�8ȌfP�9�G!E�nL�;*K�� ll��Rʱ�6�:��v3�v�C�t>l��!��t�sU�7#��1�E8uC�`Q��m0J�ګ�Q��*��v��3u�!�**��g\hJ�8�Z�$bZrFy��c-<i�M$���Δ���Z5ؚ!<���g;m�T���I�NZ�@��U];�\���]��vwD������;�j�W�غ�wj��L��j[���Mk5�uN�|*�	� �z�� �C��j�p�PS�U�����?#�'R�{���tų��Sn�9kת�n �;5��ʬ|Ĺ%Չ2��8c5�̧�q��S-ηE���f��|��p�7b.��h�{7�	�,��>��q�-ك2�RT�����T�N#u�@� ��8�Vb�F�)4a.pK���S0�\.�$�L�rb�(�̕�ȝv�Z�X�L[�a3:��fY���ѱ�ӳʥ%vح� �4�7�=/K:u�q
��<7m[kkq뱮R��U��B(Y�A�L�T�'�'A�d&tn�o�{oߖ }6<�� ov<l`�6�ӢۡZm`�c�>�`�c�>��Y���g����էJ�v�V����ݏ�ʪ�R]۞X�O<UZ����Z�L��`�c�>��X���?R���E����4�	6nw ��}���{׀}�p�:�����DI��*�v�6puv���>9�oW���l�k;�;�6�hՉ��m�Ս�����#�>�`]�xݽ� �4��YyC�ƕ���'?}���J�������{7{s� >�=U�H��V��tpn��.ـj���>��X�dx���%+�NҫlH����{���s� ;���>�`{�����׀zy�z�MҷN�n��k >� ���uwe��wݼߧ�gf��ֆ�-�M)�ˁ�;M�A��&�#L���S�z����KWn��B�Wm�w\0�����}$��������V߉����Gf�WK�f w�~�q#�s� ;���>�g��Hվ�����`;k�ڶ���,	9����6x�����Қ��צ䄛�l� XQm��i���X������;����c�>��X�
���N�]1�x���T�g��wny`ݑ��Wr�.+(�e�]3�ۜ��E͹+�k�!�a�"�t�=��r�*���-N�U�tpn�h.�����>��X�dx���j^Rv�n�wM[x���\�A���ݏ� w�61)I��[�E����dx�p��F���=�~0��l��t��.�Wm�~�/I�0vy���[Rஔ��k3��䜽��;%�f�R��2�ـ�ǀ~��������Ӏ��x'؝e�+���sc��y�;`�J�P��t�
1V� �B�e����Hv�-�m��� >� ����x͈Ie�m��ҵl�:�%���=#����'c�~�D�����E�������G���+������}��;��V��tq�J�E�0����� �엀M���/);J�m$�Lj��'c���{�_�zG� ;��W���TQʪg���UX�ã�AU�9�][N�݂��P�G"��w)Ů4:�Ls�ܼ�u�:5[%R���ŵ�m���	K���M�덈b�Jc�i6�lՔ�i�˸-���7G%Up[#�%�]��))c�f©	q؅v�:,��q�W�mF�<�����s���iӇ��Boe=F�%)	�-��9�y�p.`�]�y�D�+g�.���'�]����o{�t�l�Ah�Q4�mnޠjC\┰�/���sh��-������1Y*��.ـy{޼n�`{#�'c��=�#�͐��gp��ӟ�y�l~�����`]���:�P�wo��ؙwl��y��� �엀N���ը]ZhC��m�o ����^;��+���Oߞ?{�I`�@�ں�V���^;����	�p�;.�Q$n�>	�v]��(?zI��Q�4�m�M�[Ef��ɬ�G�r�«tՈ�b�ۿ���� ;�;�Wd��H*ʺ8Ӥ�V��������M���� ��;�ݕ/쫫���Lj��'u� ݽ��s�{c����	6aj�6�ۧV��f�#�X�?����=8݇�u��3d+-�����U��{��=���7ob�"�J��:�ZM4���.0]X`�c�iH�r��O@��X�"��8���o.��m��� ��v�/W9ʪ��?}r��:hwi��m�o ��Wv^;�;���!Rʺv�:��Z���$�~�$��ٸG"������Y߻�nI���f4�%IU�5e+�Ywm���ݏ ��UUr�.�y�x,U�tq�I��[0{����M� ��f�&0I�CJ��,�.ef��v��������]��:1֖�&�]3��Ƭ���I���'u� >�;��W+���{��Z�M�v�զ�nـM�=\�Uq#�� �<�	�p��>{�G�FVW�wߞ� ��x�\0]���KmD'v>
�wJ��s�\���� ��j왹?|�>��lu��f䝽�.vhhwi��lv���Wd�{�ٱ���=@CT:���6�Kp�t5����ܼ�H��ژӧ<E��鶁񻤮���޼{�ٱ���`IT�c���-���u� ;6<v�X��y��$l=��*ʺ8Ӥ�E�0}<�	ۑ`�%�u� �T�C��]:I���x�Ȱ]�x�p��+��}<�I�-]&�;t��|���5vK�&� w�<v�X�j�EG8�B$X�$!�B��	�<��n��l����J�u��ӑ�vRvޖ��Cڰ�*i�5��!�	����5KKw�5��4m- ̤�\�P�8�<5�(���V�:u�UX�kG\,�'W;�e}l�ݤ�8�<=Խ:�ݴ��;u]*�`�bc�-�vGr�6Q�A��X�n�v�{t��;3�ZNش��`�pU�%�n���G������T�e�J$�`b���p�I��|�9�<o��%��dV]����S�x���k��i+�RA�M�z�7&�=�Fӛ���t+m��� ��x�Ȱ��.��J!;��]�ujـݏ �� }$x�p�URG��K��c��Э��~���� �����6!*�n��]��I7\0�p�'nE�HJ��V1�)_��o ���ʪ�g���߼��#�2�5�G�\n�t��jr�Q�z��I�U��~��>}Xc�t���n|=��J�YƝ&�.��=�:`o׺�wm���� �Ҕ�I�v�!��;fw�w��6 �,J�C��Q*���μ�\0�g���?{߰�t�t�ӫM��k 7��� ���8}����w���3h�ª�	��n�;r,�w���:�J���@�ں�l�7v�0	ۑ`�G�M�v��	$������u=�/!9;Zt��a��f;s;1��&_<&Q&�hv;��bul�'nE�I7\0ݧf�RYN�݃�wB�k >�<n�`�N�Ȱ	�V1�)_��o ���ӆNP��}���bE�O�HK�rS���B���6Ci s�x���ӄ�b�!�ϳC�g5�h�?F$ I�6R[I�s���������?]���ڎ]M�����?��J@+��S"Ѱ��HYt}��5�n�~�$�d�����j,���8A��V1 E�, � ��ã� ���)1 $ ���G�i�Ba�M�I������Ā��!~@��j���\���E!0(8����a�SA����ÂP8!��P�Z(O�oQI�k_!�)��X%!�=�����cub��C@�����0�h�XwB4D�����5��1��Y��͠ $ގ�\f@aIQ�O�#���^���3N�H�$a�� ���i+B�Bfo��X\�[7��d�8q�w�d$$֔0�?*��
A��iҤ��~^( �SB i"�`5�\��C�PbE#q�`\@���|!��_w5��$�ﻭ�?}D�e*ʳ�:M�]�ܥ$��yo�x���{��r��&x�;�x����m	6�'V�.�x���u� ��y8}�Y֍����J7��W0��,��s�[����8��#��5�겙���v�����G�M�wjez�����׀zQ<�����&�N��x�p�7v�Vd� �H��T��Q�I;��V�V������E�/ >�<n�`��F�C��e[�� ��^ }$x�p��]�U'�5H&U!�@F�C4�l�f��7$��T,��݃�wEݻ��� ������>�"�=\�t���z�N��%b#�Zj�2�T�e�֨AX��������J�ʃ( �lQ��x�_�;޿���I��}.E�s���������)VU�i�cJ�����r�I��� ;�y���}$-e;�E�BM�I�u�}.E�l� �����M�YeҶ��-�B��=Ļ=�I����}.E�M6,�c��	��6����ӆ�� }�<�G��n��+����ź��ue�u
M�{&
��By����.��7�%���qp�V�C�2���۷�;8yJ8P�U)R����s�m��W��I���\ՠ7*JK3A�X��mp>���83��Xz����bL����60�onI�,]��P�5dTӯn�(��w�M�5�:��Q`�^3��fxzڶ㋓�7fy�3b�)Ԥ6x�.2��g$��pӫ����&跂smg��z)��%b=�5F���2�v��v7E�@���X�m�l��`K�`�#�7u� ��%-�v�lN����X�����`�N������y*SUn�񻤮����x�ea�RRJ~0z��H@�)^SL�|v��I2�[�/ ��X����%J���'WM�m���K�$� }$x{��p�	�N�i�f���.����كӎ�H���;E�d#9Nk�5ٌNJ��
��M�C����X���$��_~;������劐����Nw���М��X|���0��@t"!�	��No[ٹ'/�sp6\� �lYcv]�MН	���e`���eȰ�#�>��D��ݧ`[bc�X��/ �r, �H��� ��J4Z��r�J����X���#���ܼ��W}����T��c]�&��4S�^��k�nJZ��6"���_5!�tZv��ac���x��}��/ �r,B�J�e+�wm�ob�>�ۗ�N܋ >�<�DD ʲ��[J�w$���w7$�����p�(�~� � �b��f��krO{>�ܓ�B�j�WN�m6+�x]���#�&�ŀ}��/ ���˥m�l�[�+o >�<����v\�^d��ϊ���.ց|T3+��8X��D;�P����nI�z�ر��N�-�:�6�6�,�x;#��� ����wv����Z������� >�<n�`�)(�V�c�\�һw�E�/ >�<n�`m���6H�%yWc�O��]ݷ�I�nI߾�f��>�����*��H ? �^��nI�Ӳu�͚���e�v�7\0W+������׀��^�y$����#��:W�����B�EͲ=r2�2fn�ٳ�-�Nҭ�G`4�Vq��l�����~�Wd� �H����7�<���/V��t�&�b�w�� }$xe�X�{r�ܪ�$I=̫�-�m���	����xe�X�{r�{#�&�Xݗlt'Bm���,�x�8`�G�}[{QZwv�������x�8`�G�v^ŀ}����(�č���Q�T�-��Uu�3�UZwC'l%���q(��9���z{��у��Z��˚B��T�s��r���Ξpl��Mj�m����W�\�A������N�z
F����X�lz��.n��GN�"���eJ���s%���"���� F;���Ԍ.���.�7"F�+�5��vᱍ:s��B��G���v�M*�3�ap:��$։�4]f�ѫ3��Q�*����݄� M�˕+�53��t��)��32#H��m[������T��F��Օm�v��;<�� 콋 �{r�	$Wvc-N��I[0�����`on^ odx�J�)^SL�t�m���`on^�(�޼V�׀wBTIU�j�ĭ�m���5vK�:�%���`J�|ƺ�����_{��}�^�{6����z�,�]���v��.�1
� 6�l�����%�o:T������|L��FffR\�U��}~��p{���on_�A�׀zE�e7e��	ԗZ�䟻�v�8(�B:�C�DHB�F�5�0�,ਮ�2OK���m�, �H�����N�݅4��+k �on^�� }$xe�X��J4U��챴�+o �܋ >� 콋 �ulx��^Z.�>7t��X�dxe�X��ǀ}��o �t���-��/��M���t�,"ju�4FZ�3R\�\���`zv����y��t�)]2˻o�7�<���� �܋ >� !VU�j�ĭ� �kc�7�"��#�;/b�>���wCb2�uf^���� ���xi�$�ČC��i����w$��lx{*V���)[�I��vG�M�� ;���	ۑ`�DYN�v�[�M��M�� ;���	ۑ`����?ԟ�߭�1?(��M.�ي�l�^����� �j������8�I�+�v�C��7jy��"��#���^�we�i4�30����'c� }� M����� �	f0v
�>7t��`ݑ�ݏ ;���	��v P��j�WL����{��s��������;0�7�D)&U+K1s�,�BQ�d����w ����K91�tV����x�8`]��nǀI����b��s�n��^�s��:9�V<��v�Q%ͱ;�A�nDy��%�x�p�:�%�ݏܪ��^��7exʷE�V�V꛶`]��ԐzO< ݯy��� �ݰ����al����	� }Sc�'c���/ �l���wv�)��E�x�8�k�� ����5we�ݏ �ƒ��;,cN�o ���UTrz��{5$�>���$�TU�TU�E_��Z���Р"��*����J����
" ���P �A��B
�AH* �D��F
�A� �AP��H* �DH*
�D�� �F
�D �@
�P`�DV
�H*Q`�E "�AP �EU��
�P �D*H*X*�
�F
�R
�
�
�
�*�X**B
�V
�P�� *@�� H*��
�QR
�P��P �DDb* �D
��� �A �A`*� �F
�H*���"*
�`*�*"*��* �D`*R
�  �DB*���@*���
�*� *��
�`*���������`*R
�@��E**
�
�"��
� �F�"�@��F
�B�����A �@`*
� *T��b*`�A��B
� *��H",`�B�"�B� ����E��E �D *X
���b*� H*Q * ���� Q *Q
�P`*@����D`*`�D *"*
�P��@H*"A � "����"��*����Z���U�PU��@EW�_�TU�PU�B����@EW���e5����P3�E� �s2}p��AO��R(.�ӣ!lklTي��Ĕ'L
   �"�  ��>@�)PTP  (�
�QJ %��
��J(��BR�RUR P     U	J��    � �  �) � �Nx��w�K�\��s�7��uOy��������o�^;t��nW��d,���J{���4��� ��5\����<�4��_s���{�y}k���wy:U� ��w��#��\�=<��u��p  �   ���M=�Z.7pj�{z�Z9v��� z&���xޯ0����Z��}�G�*���_m�w^ ��zQwg�+��SO=_mŽj�������*��q�_< �������u��yOUٻ���>�   
P  �Q�4(>{�[�|�����` �w{� �]�w04�  �`tr�(�g��� 1   LA�8�� ��`z �`(6 �l� :�g����ӈӦ�A@��:� t  y�@   )�0UX �=(�� �zާ�^.�{�T{�Ӗ��S�N����/m��[n �S�����[��� �|��zo��{����
%���[q��k�7W��wv�ͼ�w�U� �^W�[�u�9�{����ax ��  PPI��Oo���ץo7I;�+�ͧYp��^W�7���}��={}���� }�O���}�x��  k��ڽ��N�\ ����6�is���O,�o�Z^��T�w����-�x���3/y����^   ��)���! A��jf�J����d�b'�UJU=Oj��d Љ�U*M�U@24 j��J6��@ 4 DHCR�=Db���P�o��Q������)����n��(������5���@]"�"��j�
��  *��TU�
�_��H�@�#�	�XRfVP�L�QB@�% S�H?�ַ4O5����������#H��ԕ@��[
aC4��ZJ2�d��rsZ0�&������!8CmXD�!G$)f��X]U��^�mo�k��Z�x��
�ݟZg|������X�HZ�EX��uN~�X����=7��j������Oo>])�sD�,`E���y�|�d��d����@��.ލ��<&u�}˳[<3��(s�m2���nV�]S�*C.�=��5Zo����p��y����ɋ_O��EsU���4�X��{�s��2��@��2�J�(J�j�I�s�y9�}����/�hc�����+nx�_��D_V!L9��!&����s[�O��p!R0�c!��@��5`T�Q�bŀI��	%�dt@)���\���m��!�X@�f̧5�3p�'9"Jɇ<y�o������A�o�IxhѲH�1B�H� E$�o�f��1�	L�<՟rP��s��ѠƔ6'��X)������|��� �@�y�sQ]2���
4��0��/��$8ˆ�T��zkӐ�r�F�*NK��#���!39��Z5�-s�2����R{Sޥ�	j��z��u7�o�+>�Z����ټm/��}���4Iˢe6l�3����{��R$hV�cL��<g�9�>׌�f�g���.����L�.���Z�EY�W,��.��`��$bdw��$+�ެ:�%�SXQ�!hF��D�2�2�V^'����t�Wc߼��`��ߍ���!����eg�VX���-f��xy���pe�R��~kV��(hS/�:��Ѭ�R7S$aB(X0�@���
�G��y���P$i}��-T���_����X��{,K��+~�6d�p�#E�l�@��R2�A�I�����S�3G���Iy��xK��<�9�i�ZS���0!�Ja/��H	�Ȅ�)$l�	�sX���.�P0�K����nRe�<���r�j�}J��:Ck)�g�/��2���0M0u�.�t=g��	��y�8�(8�a��s�]��3�o��9��`@�`��Cc��)�f�t`F,6c�!P�H%�&��S"h�l2G��|ٖBy$Yq���K����x�aL��o7�����
�/���kS]ʑ����Q����	IR��g��=�9��'��"��zL�o.���ݑ񴐞��⩬ݾ�n=�W�/������~�sӇ��!p0ӷix2�].�G����3t�\M1+��1ߤ�ǆy�o���"2��4]�f����f�r���:�Z�$*�Oν}����v��W��׹�w��H���m�sշ���s�g���Ĺ��i�>uЀ@��������ѽ���;�ٕ&¬R,��4� VW 4�R<a�ȿx��y=�c��&��ʕ*�
���HM\�|dg���[�٩|�''9�疟]xk�!��d)K ]�B�G=���\d�bE�D�a�h��T���y�5=��GlHc����>�����+V%}�����g�[�~��HGqk
a����K����ю�W�~��o�9/�<q|��ӏ�-����_g���|=۪=�
�ҾF�ᬼyͻQ�{���﹛�Zs�y0������kZL�i�z��/���F��D��������pq�H,
r�x�ݼ3�s4t��}<r]s�xq����2��4�2�P�Y0�)/�s4M��4[�HU�z
3U�U�};����:_�^,�Ar�� U���H�{���Qu��ĩ���&m����Uw��<�׻��.B�+w*��\�Q�âx|
�"	tm>6bZ�:`\�<�f��y�^ߑ��n�RZ+�
6�'�5垙���)�����q%+K�a�q#j��kY`B0�p�4F�Au�B뛹�Xq�B1�h�5�Cf͹�k�I�D<�<��Ղ"A��4��B$� 8�ָE�.��J��!j`�B�B"VC�F-�Z�X�6������mb��}�u��Mux��������"$�(�SJ�޾�{K_F$"p~� K�[�=�>�|�|�H�A�zE�!fk�����q�s�g�\�,~�������V}�s
���]5��/5M_U��^�)\����m���V���+Ǉfފ��|f������"�5�>����v�ժr���u�IQ�UW�W
╮�V�Dպ-Vq������f�O	u})�	\A�p|
9�&D+��$B&�$�@�t��j�V���_���C��R�W�8���e���g�ov�OsD|Z*�^����HFд����l�`\4m�)��\H� BBs�T��CF�!$�	E����}�`4U�m0>�_g�R�j�ː�B���#�'�3���j�6�nkHU���&ؙ����KB����O�v�Xh�4]nq��7�%`F�L,)�+_Z��W�jm�׵���O=<6}������L��&a��]i���/�o�B�Y"�F�y��8�{��Ġ@� �w��}R�b2YY+���{7�>�:�OI�<�O�O}�.��_Z���ҽΧ�ب���{��M���!BG��@ꇾG�:�'�G!����(pg)}w*�W�Ū��<^���籄��_"����a��{_�z֭���e��&ߖ���h�9�L�-���7vI�CXid�Ie��c�#GP! �D#�,tE�)�+� +����\Q��R�������Ry��)���s�mcpק5�y�D��_]Hnk��;V�}��[Y�?e����Z��������?��	�`F�I����(ĉ�����a =���E� ��X1D� ��H"�!�#"�b@! � �1H,a�c �"D$BA# ��@�A�F,1TB2$H��  @A �RF(E�Q ��`P��kR5�H�q`8D*@���S!�i�r2H0 ��2HB41 �H2LH�)D`�211`�X�@�Ŋũ�32	�1r P��@���R
��`p$4D��CN$
�@����$t��$pt��������I�$t>ġ���lؙ!� Ca�i������0 �CP���H�00T�������$e `i ���XD���FDȓ$�u6�����̛�q�������D�鹖�i�_.sEe���*y��7[�ȓ��\ȳ.�璖�a��xF��9�F�Sv����ٰ��bI��t�
��@��͚|nM��n� �X�dIH�H��g����{���h�ݞm4���m��d�y�fK�@���x��g.)'��o�����{&q�L�̘B�	f����������`�dH���ב�6}��D�k�<<vF��a$i��Jf�5����@�)�.jH�:���y�T֧	T��A����K�3�u��vh A۰�)����������	#��7ʐ��[�M�9�d)#	7 @�$"��K$�X�`j�!cP�>Bm�HVX@�ˁg�>���;q0��a%��ߗz�X��<�ڒ,����<���^Vr���UؾT|��_z�eZz�B�ʪ���Ye0����I����HI�����L#]p���]$$zc,0�.��0%0���{�y'E���q�-������+�9�{!�%�i���_!R!F$c1�@�c��	B�d�Z� D14��,b�P5��)���!#"j$"�����#b�P R1�7�B���u��7���	�@� ��h"��$j�,�*f����l��A��8�v��#ǆ$H[�̘g�������xj@� ���l	�4B"1�j7#	��!r�hf�O�H{�{䱐�@�!�����wB,_8�ja��l��f9!"�D,��Y	�vɚ�ia0�6OY�q߻l����ḨʜM^�<���a	U�!$0���-�� 0d�c"}��q� �&�C6B)��svR�֋+��0#L3f�7�Ԓ!!0���3R�_'�
����!���_���ׯ�1�S��硯���#K$	2V	�w�9R�.�����*B���ڀ����̀�W���{���m��m�Km� �� -�     �` � h $      H��          	   6�l �  p h  H66,gFY��I*����8�(���үe薪RdwT���u��ὮA����)J�ʷ��Ue�mK���j�ln,�3EMҳl�q:ٶ��%lp m ��U*�U)!�-j��ST�.}� h=l���pv�m H�^�̫��� y8iV���m��)�  �� h�H�� �6e�eXݩI����kk��ٛ9��xG���V��
����f�b��!�������7�15�#��,�Z�G5����m��;�g\�^{ On��m���Y��s�&�}g�j!�f��&��p�-�ېMh9N���qCb�j 
�,�P�ב�5�U�mq��H��E�:Nݳ[ֶ��Wvō��PG��*���6��u;@S�+�V��mīd����m	V��<��78�
9c�����r@ ŷi״�I�[@ ���6���ڳI�#6�- ^�qoMf�a�{I��D�����6݀ pIj��[��mV
z���UR4��H��.�Hm��M-�ci�P��sջs��,R�6^���i\�q��P]/V���TrBU�m�[[t��Pl�ul�y6��+e��rϬ�A��z�)��C����1�I�0��v�{e���v�KQ\�����#�L;p琞z�7h7�����b�U�Cs����9�Lճ����\Lۆd���t���V�q-��&���P���6֧d�Ե���RR�czݥ��$��J���t����=K]9�d�ez�ڜI�Tx������vJι�Jw.{ �v囩V��yءV� �3�Y�⚪2�KҼuٗ�Fwf�smu�V��5L�eC��8�n�j�ldUj�b�����r�i� ��Q���REK':j�.iV�ҬF�t�Bma���ڪ�ˁ�BJ��M"K�	WQ�l��gvWkv�T�-0]0]��8ݷ��s-Q��������6%�����U���2��K8˛;��>�3�I�!��B��L���r[ay:�.N�-��<q`S���I���� �kK;Zۣ��i���'`^8�<�xz�Q9ٵ�1��>�u]�U\Ή�������ٺ�m�3�����oQpV�؟��®�V
y�SST����[���[&M�6��LN�H9��]e���N8h-���	�Je��������  !l����(��J�� n^��J���i2l��Lj�U��KD�ZYZ���Q�k�M�R�ԫ*s�;*�d����S�j�˵UUFψ5�.�p*��M��6��T�U�折pzz�
�URJ�9D;v6]�-p�l���{V�n�P���&�Lv���O73�<��u�5pXj��]gv�'����v��}&�#<xS�ظ]���݉�[�Ӷ��.�8�M�@  I$��Md�t��W��Ieh�nZ��
��Ӣ��@j�:��P) ����m���`8/[����"6�R�U@\Z`n�ږL�hz��%��M�XV㓆�*]�8�� �����`��G�vݖ��7�|�am�e�m��Y�$�-$�*zГ���]b��V����fp�  	�U��%���8Yu�*��ꪪ�G9N8P9��-����mn��dkd�&�� H l������� n�6�m�i  IzZ��m�cjͭ�Àm[k4���ԛ���[ 6�  7m�h�m���l�^\\�`0]$뀐� _�7�  $  @	cZ	n��   e����UEq�<=�
�yoll�n��^(Z7���   �|��@��͒�knCm� 9��&�n ��s��[v�)�W.�Oc$G�q�>��\�㟰��\�v���f�`rK	�4�rm���U�h7�x�@7
d����X�cSK�-UZE��T	T�N�Mo��@m���8����+D��e�$��  ְ��kt�OJ�D��`H�j����붖
�.���V��jFYܣUU*�m��]�P�.Z��2��xV�g3*�غゐ���yUvkb���֛8���7<�T^j�����Ǉ甆���+ŗ�V���v%�en�[�v��z�l�d�o�� �Uʣ�i�td��ۏ�<��6��m�Hk'��k����  ݶ q��6xְ�j�ݑ%�l==�,���K�a.��Cђ���`:[S[@���m���mv���m��B�a���[UY�d��Ͷ�>kh�u� 
�]u*�\pJ��� a�  �[@9�P.I�X
��IiVŴ� �h8���� k��X6k� )[l	M���-붓m�`�-� 6�m�d � -� ��@H  ��` ]6 B�;`p����S��v8� �tX��0�ʪ[,���TVж�i0���!�0� �  �lEej��(�Z�ekP�CV�[E<��Lv[�,�A��ۨ��$66�a6&	Wi:;îJV��N��_i�R�1����� ��N-��۱�λW]!:	�z�Ź'.� �����}���~�S��N��ve\�6ת���`A�-�+d&G-�⊪ �d���L�����;� :�ר"����Cmձ(9n��:`*�y�bڡ�"BY�V�L�[wm� imi9gT�fŴ����̗Ζ�v�.1GR1,X��\*�Ω��9��K���kn#����F�9'��vͶ�d8��>��m��j��Q�2{ �����t����5V"^�h
El�6�u��8�L['k� �٥�ƺڑn�`�����՝Q�Cqu�L���0SUO+�j����	f���M�#�X�#����e��9�`e��������2��P� W[m�	e��j�  ��V�XvÌr�[5UPJ��T�m�����m��m� p $-6m�1m�,1�4Pp �m�-�fݦY;^e�� �@ $	    +�W�h���[;#W�� 		�A&�ٮ�6����e�6�:7n)V����C}���|��&0ứ�*�U��d��h�N���8v�ʙ��Hm(l 0q[S�x��%J�mg*�����R��r�\�[*ʦ.�퍡���C�-�.��-��]��i�V�ڕ�WVIn��Z��Z�I@�X m Z�$��햜$[��$|p 6��b��[G m�[N�p�� $kՉ  ^mR��[i(Ӭ`[@ ��u]M[n�6  D��b� � [@ ��` -� 6�[m� �  $ [�  6� ڶ 	  m��� m��ۂ�kY��l��$l
]پ8��CRR��[ml6ض���� m�UR�R�J�����Jˀ	ԁ��  $ֻiWJl       l �m�m�@� �        [A�I� �g���  ��   k�        l�@6Z                   	                          h$      �|                             6�m��[[      �`$�	Hp�}��-��5�m��H6Z pЖP� kn�`���!�l���`dH��-�h���@h���&�u�68 H�b�h��P��J�N%٤$#]��mn���� �H�L�����D��	           �f���(�bE� 'm�    #m�� �6�[|  p$��� ��m[-�ԁ H6�6�8k�l   ��[v� �[ 	��)��
������u/�@ �����HM*�T�R8��v�,\6n� �[p��R����ֆ� 8-�m�Ď �p�`p-�I����M�Vv�m�P849�G�6�&2 $lĺfֱ��� h�� �Vډ�tK��	U]J�]%.Ĵ Y�玦(X�0�]ʾЈ<#I;��˫��3ӫ���[a�n�v�.�m�@'ݮV�vZ�[B�m�Lb�eZ��k`(S4%� kXw[�r۶�[��lH�P-��k� �Wm+7�pw�/7X�^���4�\�%�@ mm��ZM�Wm"�  �ӆX�d�� !%�6�m� [@  �`8  7��� z��nY�Kک�9)Z����8긳9k��aбpڛ�7O&��mm�6ۖ�t��̻�ڀm) 2V�]Wg@#\���c��6��Հ�lfi_��{���w��s�� 8 �)^�5O�� t���a$Ad@!H" b��A�	�@<%�㊧ʮ�P�:U��T�&рx�D�4�� P"A5�x`�T��,AO �F.�N"�A�|��U_�!U`�+���BA�A��]
g�D��aP-F��"(H�ډ�	�!� �0��E� ڰ� �x	����_F��������M���+�xz��E���Hϴz:D6��D�tOW�x���C@)�!����}�L�$����
�����Q~`�&��N">�<OW�QҐD"��I���l>H|-�P�x
�@�_` �v���HB,a��#;Eq����(�{��(��T"x��t`�ȨH$ �� ��%`�1G��=0� ���q��@҇��~���"��8 ʵG��ldbx(| l��dT#)FF($b�����`���
>�j���ʭG�)렉B,!	$d�CG�`� B���6$S��<=�|x�]ojd$H�Gb��	"��|���}��!��`���%`�J4�m F",Rʯ��������f�D�@16І@�@��WH�/� i�C��4kآ�s�������௉�?�(U�"L#C+J ��D#U�Pd�!VQT�P�dE���37�kZ���� -�� 	$p����%D���m�����t��*){Ks�:L��a�Nr�dj���=��PN��׮�7�9�n8����=q��qkqη`L�x�(p�XWI��m�� �6�kƽ�k��jڞ�����^1v7q�3���nh�α�:�8�r��Nb��k�������<*s�cs���q�ۺ��v�㬥�;��tn���$���{�w-ha��	�=\�3���掸��a뉱����omd�tU�;b�nlU�k���Z�i��r٨�]��^7�^}���v�m��s���	zT��FY�q�c�;Nr�p�;Z6��\ ��������b�96yٞ1��X���� ���X���r��,
�imf���j���yU�m��"XLӺ�)FCN�(��..ʻm�	�J'Ovư9���:�Ƭ�R&Ҁ�q%��Z�`���7XS�W/a��a%�\�&��1���ɫ�v	gi��2R7;<g'a�uL��5T����F-��2ܲ�T��S`Hd�୶L��H��0��oFx�u�@�F�|m�#��kv��j��Y^��heu^�fs�b�����UPےc�\�v�O$�ح��M ��u���E#�k8�㎵���m������:6�H
��f�uL�9�Z*�bzDk��������%B��D�ݶ9y㪮K�K��nm�dm��H�[������	�	��-i
���vlk]O<�v��'K�L�E�M���6E�mp �&�ݛl� ��   �`    ,0�     հ /E�v�t�VW��k�wf�\����R�@	2lR�UE�V�@5U�Y&!�*ϗ�l�i^�_�д�<;�I^oUlQ [k�T^�ۚ���Y�3��+8l\�)1΂�p�����@j�n��ۊ�� /"�\�r����WZ���&�S2\�I����؝ (�H��hDЊ�@?"~�/�>(z�����Я��Q섙���9z��g���.�a�m��8_�o��!m��zT��/]�@��l]69�6�j����v�Aܻ-��S&	�2붆s͞��l݉�^z�������J/k��q˹�oe���պ�=!Tl���JBk���I2&�^+q �Z� 6���ܣ�Bx�V�Wg���OUc	ٍ��\��b�%a��� �)��˹�2��-��m�M��*8�3�������^����x9�G~-z���7���@9�ܿ�K����gS�/�� ���j�7�v��l7�� �H�oF�耗T�р]�^Y�loL`{�i�7�L	�.[�S!J��Vax����0&�k �M�08��r�n�	Y<�����7�L	�.[V���0?_���ʹ�Sp���،Nӓ4X�9�v�l�͵{H�,�kG]5������p�˺���;�����&����LN�0�\�S��Tp��ev`>���j����AҠҞ��ks{�Ƙ�`{��ll��`�fX�Y��f[�Ѧ�F��$���d�l>of���	��UҖ�V�۸��:[kz[�Ѧ�����b̱]�&�Ζ���-�����q`Ij�]�Ae�J݊�H�ju>�;5/S�eG�.�Qi�v��FƢs�@Z2�%���g�q�����7di��9r�
�1U,YX��.���07di��6�K�Jy!�ή�	S��;+AeX>�q`N{�߳s�(ADNA�U�0������y��~��y��X�\�R ���[V�!͘��lwF��4���EV�V"�.��Q�l����07di�0x�����;Sr�*I�qR��	9u�a8D�)��X���kb�D�S�ٖ*EU⼬�`{�4�ݑ��Ζ���-����m
�bʼ�3/107[Ś�B��{xg���|��`6��9�Am��Հq�sn }��þD����X>�q`�U�h�J�KfeQ�lvL`{�4�ݑ��%�i���N�3�����y'oI��UuYQ%�����=�w�!͘��l�;��ó�8����&kG�[�>�"c�ե�s p�m�R�zj��lz�p�V'G�vV�ʸ����!͘���y��{� �.-� �+e�b`{��l��lwF��n, [��58�uYlV���m�=�`M���gK`oqY>��&�-%r���n�Հw��X��6`����9��UҖ�V �׋ ؈��|�^��z�`
 ���Ą\�A��"bF?%i�j�g��[�fk52�\�t��;N64W8v9y���In@];uQ��Y��k����@����\�wj� gm��es@�b gjw�-�h�������kIl�@�T�DH�U@[���޽]v8�5�{Cv�\q�en\;K���44�;6�MԨ1mv�����Nm�  �^6�8���&Uh^��m���׍�I3�b��6�R�~ٿb-'7����3P�:�kav�)��c��ݣS�Ե͂��n̂�m��t�s��lv��C{0sf���oF�+�L�VU�̬̺.� sκ�)���,{�� ��u��]$V�գ��Y�{�n,~�ŀ{�sf��ـ|�վ8Z8��s^b`M��Ζ�'t���L1|�m ��'a%0yl�޻�>�^,��0Q�Kz!t�!�����=��[a�n��[$�m�ڷ`��'�ՠ��O'e�zu?͍����׋ ��ű��C����n��|�-�hr�W,�=�7s��O	.�jk5/n����d�tS����Q���*��X�� ���9�Ю�"�3/106ti��:�K`{�4��QEW�v�A��*����""_n^� 绵�}޼X^,uMd�(9|-�W[�`n�T*\ox�w�� �*z� r��e�ct�����4Tn y�n^y�pqYJ����^v��Kvvk��.�e����06ti��u��[%�6�)�YV���V����׋6"Jd}�{X�w� ���X�\6����sv�򧮰��!DU("P�	(Jb;
"�!�"�+ذ>�X ��LVA�%��7l�8�ݘ����>�n,�G͘�q��P����I\� �ti���Lۮ����-��s���i�na��U���b���:�ѣĥj���sm��z4ƭ��F�3�mΕ�1���L�����-�����E�c[`��`�>lΦ�|�f��q`o7u��]�ΦA��º�2����`{�4��Ѧm�K`on�KTj��m	,�=�7��pܓ�2��nI�	Hh��OUv�_�No� 9��=���烕�`oF����?_��߿[�Ѧt��� ���Г�+��"��+���d�庢�*�J����}`��m�>�`q[���:�~�V�lwF�:4�'.Z+ Ӓ�e�`n�����n���q`�>l�7���`71^Ve�=�`l���륰:�K`l$m
�b+ef^b`l���륰:�KaJ��<����-�ʬ̱U�&m�K`ul���ti���,׈�˚�;,�5b7d�i�i��1%%7���,�!x�nͷ��v�r�;�J�-��l�I�*>�<� sQ���mq��gZ��6;r �m�79�����]m=g�hF�i�W+�(`�U��E!�L��rL�2���}�U.xi���mﭷ�Vg���`��GrMc[mb'���ِ-�m� �n��ucT��{��JW=�c�e9�욺�x�ter������h�8�	2\,�Ԑ�k5L�Y�̎]��]<���+ٲZn��U�.d5*\<�*d��-��8�yـ{�n,����9�|ـ}�ڵ�b�Z:��/-����oF��]-�+z[���V���G�rT�*�7�n,�G͘~^7����>��,�_yͣ�;EX�3���:���=�`ztk >_.!��%�vY�q�͘|���W�o;�X>��0��$�+�L9i�ٹ�4��%y��̷��xz��Uj��X(8�H�r�*����I\� ��n,�o�Wi��D/�;:����1*���l�`�wy�s��x�a`�$
 :@��g��}�T�loF����-�ʬ̳3/���6�KeU{z4�푦����(9U�Z7]�`=��߹`v�����;��JW���aX�0.��ލ0;di��}r�S��:������dN�%Lv��V��8�B7�:�<��c-�*İ�T���N|Stq8�%L��@�w��}96`=��߹��1}�6����;V�Wi�lBS#�{X:��׋5(�\Z���8G,�Q�f��ـ{�l����D����z�B���p��<@��
���a��Ą!�G�)Z>��2�����kN �D��!���@b�y�b�nOt�H:�Nj�f��p�6{�Uɀ����Nf�����=��z3��k{�!e&6�9��Fy�p7�ܾ�kWT��N(�2������J���"q�_$0ў�s&�pG�\���!���$J�⬬�i8C�W�g8h9Ć(�	�^x���ѡ8Tj�5�N<C��F���5��ئx�,p!�^�ǀ z��P�6��Nx�hh�P�`b�@4�D��G�>PH�k�QCb|
AD	(Q]�����{[[Y����M�U��~:��x����`��,�NM�lO�������{�+T�ɪ����Xx�,�S#�:����=��{� ��/��a�5#��vG#�%���ª�I�C��A��j�EU�EҗS�>ͷM�am�z�l��>��x�squ/�7��,����s���,��0�=��(�Q׾ŀk�b�;��:�$���ں�bmZ;KF�x����?'׿/�}�[Xl�6�� jp��l&�R�	j�9�7u���{0�7�����_��3!Y��R�(�z(q�D� {y��ܓ�<�0����Հo��f���x������,�r�{k�㬮�m`lZ��.�e��k�0��vmV��V�l1fx�X�E��p��-�v��Nu��`v��m�K`{�+.}�2����WU�lލ0;di�6륰5�6`j��"b$�r�K-X>����u��S��=�`{dE�O�ݶ�Vϣ���ـ{�n,�n��7v����v��Tdnـ|����J^���w �S�X(���=R0%@�`@`0�� D��k.��M	3�m7!̮筘%�jg���lcA�$�aF��E��ȲΗN���Sn�x��Gkp�˙����ڳ�}�U��Mqr������ۡ6��r�+��A�PpdLN���Q�m��	]`�Գ��;�6� �����ɵk�V�wZ0�&ۯBћt�$�]ͳ�  �b�����*r�/Fl�#�yp4KϜ\�5�+��I�����Pw�^oY,��+s!���y��pt�\�	��-M�A�j��t��9SUp�6�VВ�߻�X6F�n�[jt�S�Q�`U�v������푦ۮ��ڝ-��Ѭ�_yͣ�:��%� ߣ�� ���`v�� ժ"Y�eYu�w��Ve��1��Ѧl�0&����j��R��u�p}�ŀyD$�����K��>���vz)���b�e\�%;�sGLr������ʰM
N빧A����tΛ�3��X�u�`]�B���:��;�2xE�Q�im�`��ٛ�^b�ĔBp��~{x��,�ojP�K;����%���� 9���=������q`��ـs�|{"�6�+f�[w�L�`M��lgL`E�r����U���&l�0+�� 侺�>�^,bKh״+��:��iɱ������nF&�.V2�El��[h�k���X��� � ��?e�6�K`{z4�푦�TF��8Gk���f��l�=��� �۸��sl�=�پU,m �N<�`{z4����*b�_ʂ�}HT�l(P`HՕ	)>��{��'�Ww/}������ -�����Yj�=�n,~��0?�� ��i��_ŧ���]�b`M��X�]{_νŀ|��`�%�����L�+�����`h:-�Dy�Vl9�u*�v�<pݣ��xf���f_�����=�`zti�6�e�7c{6EbmZ:��%��sq`�5�����ޖ��~��v��W����`M��l��lލ0����\2����~��0?=�7$���rx��I(�� �!.B�Q�_;��, i��E�EM��fw���ޖ���i��Ѧm���;��P�zv&��ʋhӉ�I#�T�B	9u�a8�͘�xZ�C�n� m�؛�4r&��g�s��X��ŀs��^��6`��@LC��[Ke� �x�f�����ݺ��/}X�ol���P��yGm��Հn�x�هSs�ŀ}��,��>-n+H쨗uW8/��pww��Ł�QJ����x������j�ia-q����ŀz�^��}��7v�s�w��8DA�B@�&(>I�[�Jf�L���ON��+Nnq�OY�:"k�E��6�
e�����y֍����xL:���Y6�(q��ф�ݴ�g7	�6�4F�N�0E�Jf����t�ٰu1�d΍%q�P�dL��t��[v�k�e-jBr��\���3���C��k<���*6봬�l�   [dUg.jt���Zy�����ؼ�-^�{g��D�����jo���4a���d̍տ���c�ng9i�W'.�:m(E��� /,�n���D��W�M�R�Dՠ���<���9^��Nk���, Z���� �]�e)���s��s��Kʨ�[��:��X��ž�)#5j�2��;l���<m����ﭶ���c}JI�w��}m��nA�m��q<{�R��l������
<�߽�2ff{����fz���3�
M����[o�Gq1Z9m-��m���W���|K{����{�Ξ��o�ܦ6��A��*�Q�U%�K"#ح:�h���]�(9�2
������_��s?v3�`*;m$v��m��nA�m�}���[m�����y썿���{�m�`�V7�vTKe���|�����k|�`���T�ґ3#,�L�4bJHV�`�h)@� �z��~�Sm���W����ܣ���II�k}P�F�+��$�����{���>���O�<�I+���yd��������3=\��:)�A-�6����$��ߗ9m��u�.����s�ޠ+���M��kW<��"��NJ����v�O��Q?
���~��m�g��ɹm��߸s���ݻ�vm1�����vv�Em���
H�ͣX,���?~�w}{�������e��+=m����ﭷ���1�߻��uy���{�1<m��u|�X�$*�UY��3<���I(K�E�������߬���>�i�IIz��	�r��i,��o��}^��{�f'���^AR([D� "H���G`/�&s�w�9m��o&��Ͼ-1��Tv�H�^���^N��=Om�7:{�m�7r���O���{�m�`�V7�һ*%�T��>�iﭷ��/{�=m��w��}m�ݳ��E���:��2W]c��p<�P� y��&9���d6[�Us�ۭ����\n(d�
�q[d������r�o�������v�O�/dm�7:{�m��*�2�H��X&�6��y��}�I{�1<m����ﭷ���g|^IkW<��"��Nʽ����ى�m�}��}��B�D]ۯ{(ə���/���:��'�87c����o�x��������'{����Ͻ��9m��j���`d\��0>&�S�F��ߔ�HR!*(l�~��9��K�m���7��U,J�J{�m�7r�o���^s�qs�����x�o�s4����f�a]����g�^�=�
8��\[n#TBz�Y��Ni'���������?v�Vf����������v�6����?%���󜭽��d1��7��ڞ�TvZ�v�}m�ݹG�^/RF���=���;܆6��y��}��$���TV7���*���m���O}m���C�x��I�w��}m���(���u�CehV�%��\Ϣ�D%
�{ܣ&fg��|��fe�yd��GZ�����[oN��7&��������M�m���Ü��ʯ� ���<Ծ[m���Ü��3﷓v�v�/��G�Nv�!0 �(R0�"f���&
4�5KF]���]ks5�pt"�kI�������k�*���%!�$瘆n#갤)�F��c77�o�M�jk&��.��%�F�����L��h"��!���.B��X]5��Z̥g��a40d �&�SDؙ� @�[�4��3Dٍ�"����c,,SL$܋<��r�, Fo~�X @$R1�2
E��@"�b$B(@)��H�R
@�B �)��`�V#�E"�F�!$�#0�FiD�����0-$Xs@��_�)�<��C�h�z>B@|�,FJr �~4`�(���$3 ��� R@]����]���Ԭ�hO�	�֤@�ΐ>����� -�h�e�  �BBE���R��U{�[�K�`���F[�d�Õ��&�eV��[T�[U��a$vڟa:N���۱���K;G'\ۉ��V0�#��R�<�6�v6.
�{Z�+\�N�-�$m�7-u��kϬ��q��˷3��6�b@}�:8;��l[^��-��86�z�X�Ʊc.��eh6�V�M̓:QC��m$�L���۷�}�Ӯ[H���ҧjMÀpEײ��v�Z�cu۠����W�
�-z���npm�6�Y؂�3Ƈ�UJv�ǜaoc�:�<�TSq����eS�v|\��ѧZ����A��a;T��;sxL�3�\�ja�
¸^�Px����p�M=�s �n���`*���g�!<dj=�6����j��y �yΰH�=T9Uc'\Tr��d9�^Xv�Ƴn��ę�ז��Z�Ey �GY�O��rݥ���d�N�n����Ͷ&].�S���n˵ɩ��\!��;{I;;.�m�m�I���M�K�+kRLgl����2�g 2*s��\������m����ܚ�6�d7b�W�n�κ�������;�� ��R��jn��^^d���u1�#��Nܖ�idʛ����x����*�����.i���kP+��C���^Z�iQ��q�m��܎7HsK8�؝��:��n���De�/.��5��N�&�:ڪ�#mvC!1:�ꀠ:�j�
亹y{e�=�+E�.�$[%��[�dڀ�n:F�� j�  m�    m�       �`�`�;]�$m���]�����IH�� �=m�Kp�`.�d�2�N�
��P�B���~Ār�S]5��P{rpܪ��fk�u1����X�WI%�Xy�j3�rP�[�N�=hF�l�8ri⋰��xW���|�� 'r�Rf/\֩-Ŭ���\�˗T:W���h�\�������� >�1�S�W���{���w{ۿ��e{/M� v�,Y)c���[�a����c����٘��Ͷvxމ���Ź������S��Y-��m٩eZ���VI[���u��f�=eH{q'f�s�g:�r�r���N8@8������K�^9�!�=l]�tuzkkJrcYgj�����qĹ�e��`��fŴCpn��G][�x7g\g����n���"��
'���u	'%զh��Զ�qs�v{;E�#���m���L�(�M_��[�����ޥ�M_3-�duѧ%_��{��)wm��=��9m�g�o'Uf[|����[n�WP�Z��v;kn�<m�Ϲ��}�x��(Ww.��&fg��|��fe�yd�II�:���Ui J�Z����;ܓv�y��p�/�_��ֿ~���]�m�����[l�E�c��W-���co�/�{��{�m���G�����W���������m�����𞠥��c�{�m���<����~[m��ަ����p�-��3��=�x��'Iȃj79���{q��\��KKv��w+skR���w����.�z�IP햏��}���ﭶ���cm��o�м�%��Ͻ��'&fe����^��+�2f��ִs��|���l؁R-"6R)mH���,�B
PS�#u�{߻Ü��{�oR��o�{�s������vk̐˚�eֵ7m����9�m�ﵽK�z(9������{ܦ6�k�sm�duѧ%^���B���|Ի�������>�z����������^��}gW�<V���rZWeO����p�-�������������-���Om�� y�ԥe�V�Jȭ��ki5�u�ts�g�ʜf%��w�l�����wݨ�ʭ#�	Un��Ͷ���1���7���3-��S�Q�J!r�f}����fOy��$��il���ow���ޥ��H��u�rffw^���ffx�Y���B���̿��O	�
Y-v;W����߬������9��P�0B������n��y��{�m��z���UIeC�J�6����%����W�L����̙����_}2����y{����;z���
�B[e�{�m�r¶���Kw������{f'���y��}m�B�i�(��X��e�8E;;S>D�\<��j�;*̨�Ӭ,���{�B�\��H
9`�m=m���}^��{�f'���y�����m��cm������G�Z,��[owl��x��I�׿/������33-����TB���#]2��:䴮ʞ6��w��}m���S�^y䓽�������ى�m����5ѭL�)sF�֎r��C�}�����{��Xm�,�y%)%"B�@(ʉ`H��H*��!_|���wi�I+���m�7y��Dz!(^��\\��b��w�5?�m��.�:��Ejۛ�bq98����bg��UP���Uӛ�{��O�q�g��Wsu7k�7wk �^, ��{	D}!��q`w�o��c��\�v�V�׋<��""�;�z�{}� m�ś�M���r��*����j������XjJ���ŀn�ŀur�WJ��J��ɻ�Q
w^����� o������� .�Lۻ�4L�r��X[s� �Dz!%�o���{׀n�q`	$�I>n�6�5�F��:3�uok\��Ѩ��fy���;��u���ۻv��ǎu^w;\xwD�{<��b��gMV�z�N�
��"����7f���[s�'���:�Qcx_��tg��v�ԉ�>�df��n�ո�c�2��']����=���lJ������-��s��[v۰ݶl�`  v_qdYT�I�$탞vyN��Sٻ�꣋i1?߻��~w��wu�������f�љ���];*�W��ket�^��$��yRm���^�����87\��뫠~����wv������A��� ߂�e�Lԩ�W3v����M׸���� o�~�/9��m9I �[p�{� �nqa�B��{� 9���q�D����Uw7Sv�6!D�ݟ��� |ۼP���`դΣ&ʥwW5h���X}x�%
��]��|��b�9����`�"���NF�H��a\:ѐ/aW:2QH�Dճ��]�o�wpeD��(ܒ�]�z�{ۀn�q`m�-���7^���m�	���J�Y�u�nI����x�(	�)�P����q`������DB^���Myo���J)]̩���o��ŀ7׋�Jd������ΰ2˺&�������X�S����������	E{w�ŀ?-WS�.jf�MZʬ��=�cN�0't��ti����s�����(�(�]4z�9�dx9zR��y�hV���&U�{����ݜ6Z&�仫��׸�޺ŀ7׋T(����n���jxLAJ��j�7�u�=�y(P��{}� :����ŝ�x����"�W*vU�w�ݛ�Ny��ܠ�0Dc"@AaR!��F'��A�*t!rw��9��� 㦊�;�E�5Uuw7V`l%
"g�ݼu�,���`y%��W��x�<�n<�ʪA%U�d�� �^,RP������z`�n���u֪uB���c���0�Q��f��O���I�X+�-Q�n[my��9�+p+�*��F^&��N�0l��	(_Hn�ŀ5��e�EM�U�Uլ���͈����wo �ŀ>��,�(K������]�53R���� u�׀|��a�Dη�� }���u��M�Q�;jv�nW���� ��sf����w%&>��
��#ٽ����O	�([m�ڰ�b�;�� �����ŀy%�P���M2-�퍭Dpbb�dy��J��Ɗ�.�C�ۆ�}���|Yz�7e��\]o� >�w�|��l/�5��X;:��(�v�I)���s�6s^��5��Xy�fzB�$��8ۏ'I"IYGm�9���`�lŇ�?*�{~0�޼ ]\]*��U!J�E5V�5N����]�q��>}x�/�Pe-��u�hK*�9�.�|��߳�o������i|���68�ǫ'U�z�X�;a����Y���Kv���.�}}�r�[�:-�,�J贼��E��'y(N����C��?��n�90%ԑ����3<�{s��sq����R3�͒�2Y�����q��-�I��M��zqV�n#]���V�Q�h2�]�Ilz���M�m[ �UT��6ӱ�Tj�D�(�`��v
��������ѩu�55��s��~s�Yy<�9ЗF��Jn-��Y�<'
�]Y�g���^7��@����|�z�'7l��6�<�xϯ ��X�/�]�=��Cn�qT�v����Τ����X�oL ��۟�ټ�`�𘂅��sv�ok ��fJd�wo ޽ŀ{�F��"�Б�VW���׀����x�=	(�BU��W�^DP�cU�ݰ�v� ��ۀw�w{��ok �M�舗���W���3��[�}���	r�y�N���I�'h�T�9,���O����G-����X�]b�)�����wv�5�ʪ�
�W(����>��,��T(ğ�J&CP�&�h��Y� �H�0���bUGqg#Q�qDDy$�:_��� ��� }�Ś�D��;�KTpn�-	eXy;׀����I/(����`��,�]WR��ʺ��W�yLl���Ѧ�0�y�}�޼��� ��E�;]� }�ŀlBQ����9��8 �����ߟ���%���n��K��%+vM#K�L����%K��]b�����~����n�wwt]��oq`:np��J!(Q�J���,�^&|��*��vu���Ҙ�1��ѦI�x�x����~DP�cU�ݰ��^ w���0;�4ƅ�T�� =.�/������/�h��,d�C�aF[������=.�7��7���`ă	#�٭�1`����=�`�ʞxl'�����h�����	Z�x�Ő��P���e�f�f��"K���
ʩa%.�T�a���%!��ԈV�7��-t�$ޙ3�C#OC�	�*q� $cH��� E�"Pp�����8i�qR(���(�#�8?ob���
�� ��x�x
x?��M�>H.�4b����iQ"!�mx��C���y� �&��.y��V) ;%R�]�l(J[{�����>t��[w�
-\]�@��j�U�x�$i��BK�{�����;޼X�s����힬��������6�U�Y���sЋ:�L��'.�W��~����>�>CM�d�Z.�W�8 ���w��z"(=��,t,���8@����y�pyǋ }o�k�sb"&Nk�7`M����Ww�q�ŀ>��G�(��������p�uF���m��V|IN�ߖ�Og [�
�$�%$(DBP�����9�ɖ��*��.�.�`:�TBS�v���,�w��<��5��¢��
��v]�Q�H���g��=�['n�h�9|�g~��}&�>���Yh�v��?w��s�n,y���/=a�f���w<��$N�T�Kpލ0'H���S �&?�|�P.�-���)X�*�;��,ݜ׆�Jd׻x��X\�A�U��"��������IEwپ� ��׀w�x���,�p,{�V�Z�X�+��w�zB�J7w�\��b�>t��~H��X�UQ�`D%U�/{���ߩ���l�/]�l����ح��šy��֌*��;��61���\�k[%�ӹ�� �T;[tt]�v=s�����c�r���N�ݮڃ�]ٸ�.W[d���^ٜ���D]։5]R��i*��4q���;1����ظ�U���ftGit�<��ѣ�k���x���    ;m����Tʰ�Q��c!�&���g��ӆm��7~�w�{����S��3Zɭ�&�p�֝Y�c�k1�/]^Ŷ�5D�X��Un�NP�u����\@u�R[}���ŀo7q`��x�ݸ���S�񊅶�[��>��5(�9��8�v���j��.��Ʃ%,,�m�`vw� [�5D�oq`�q`�:��T�������`��wF��i�����޼�7��X�VKII%x��ŀl%�w��u�8�78�n�,�sg��(�/�^;i�m��3t��QH�������o��onz��2vy�#w�k�ŀ}�np�n}���{� �����ȉI-�ڰ}7^b�x��<!d6|�h���w�߷`}��,y�� �qMUZG+V���� >�x^,5%3�w �[��{�E��Q%
Kn��7{�k�ŀ}=��4�_[���R�&qI�����10'H���:L`l���8�͏�8�4dhr��*�e֟8���&ܼ�'�GX�"Ea6�߿w�w��O�$���YW�o'z�y�p����zû���;��p�V��FWk�	�cgF��i��rS��Q�O�g�X�VKI[������7����y� �V����W��f���n������s]��F�<��*�7��`�78 ���j���ߖ��`��DJImnՀs��xR��{������ŀ}��T5Wk,,��jNnf��z,YMי��45�1�ݶ�d\	4���%�L#���r�\��^ o7nϷq`���
�(�}8W�/�L�a5$��e]��7�6""d׻� �������9�i�7��%��ڰ�7�]s���M��������2ю�)k���j���$�۽x�w���#L<�}�|�T�K���|UK![��Gk��v�^x�{�W�ww���n��|.628��["���n�%wg�Ź��v|9e�z�N&�e���Bs˞EbmRJ�n�}w{� �sq`:�(��ݼ M4�n�ԕ!4�
���>��͈��<�}8��^ �׋=��Q���e�u5H�*��r�0?����6L`M��w�L�V��)r�\�v������;��,��Ł�DyW�o� ���L�X8�-)-���ŀ~K�������ܒsϾ����4��@��LB"�Q� �Q@-h�	�����W����੻a�����~�Kv��ER�q�l]� w8���5�[8�v;ں�<��qۧ���{J�(:����� �ζ�p��g5��iwc��M�����p�v<Zi6J�[��X��l����̡N�����"]�S�n�Z��F�����A��ĠT��6� �jݖ]����v[v��v68m 4nV"e��u�9��j̸fj�����	�xy��ض�ёZ�#��q��3��8Lt�Q��jG8V!�����w>��f�/1h����ے��L`N���Z7��c��l�d�`��y�KĿ*���� ���`�^,ؙ8�%E��u��^ }���7�����ŀo&��8��ny�e��V���{�,��,���D%���x ����e����U#��>�7�&��y�p}˦�̡er��햭07m]���&��lav���p>6����I����g�Q��	I-Qڽ����w�xy�g�B��Pk�b��k�*��f��u�.j�I9��kzGȤTh�����|��0=/�09lDj��A�9iIm�9�.�>�����&��޼ ��ۀo�[<o*%���0=/�~X6�� |��g��:�o��c��\���`�n���?��������L	�Yt@Wj�Z�9\d��6T��ɋ��U]�����ã	vᨰl��+u��#v� �y� ���0;z4��_J`E'��j�(��ʺ��`�L���w���o^��vgS`�����S#<�9i�s��,�g�]�À$� I�ȐFI	��$bH�҆ v�ܘ7�����Q��	d���X��w� ��{0y˦��w���]������� ���ـ~_ws��s��,��l�9�P|���Ez��鵺^Ԝ�X��=�v6��Z�w��J��vT\M�Pq�ZJ힁��q`}�� ����>n����)�x�Qm�˫X8�,��*��{Հ9~�`m��=գz���V�ed%� ��ـ|��a�/(J�}�b���`s�R��
���	,��$�';ـo{�X�>�f��(�*4�H'���BY�ľ�o+ ��a�R�	.���5u�u�� �B�����Ͻ��8�ݘ�{��S�V���6��t盵l�5=j|xD��=c�I��:���*Bj-լ�o�m���u�
<�z�w�ŀj�{�v7Y%��V�m�z%�"U_�Xｋ �����Ϻ�[��В�Z샶`|�k �[Ň�I$�{��Xgwk ��F�m�T�X8�����{�V�w��Kn�<����wk ��bg��+2�/vF�RK`ml���f�_��&	�yHZT���0�� � HI�O- }� �H�]@c	$yn:��d�`BB˽A��_ ����	�!P����Z�20���f�� �a	
) �&���$$���Z��N/��{���� :>�&�	��H��x�40X����h0��x��!�������w}�?ʗ��� *���  I!!"ڶ�L�g/�[�v����q<'P���`�@��햗f��6۷X_y/&6�v�X��y۞�ܲNu톰���E�su�۔���v�8��a�:M��Gi{��8����0�j����m�:Ns�[����z,�S�]Wbz۪	L��i)a���������f	��t8Y���8����7���{(�砗4�x��ؠ��Dz����6�tܻ�N�[[�9�c�`�9��y��1��\b�%��VUWf��C��s�E�&�s17-�3<q�ȇg��ռ��:U�f}�+��H�� �A	��+h�\�R;�:�m�v7bֺ�g�Y�e]���;v4�jg�[X4���+��J�cShS��v�UV	����F��*�U�F�Ηc��7M�p�OO�	X��Gp�s��㡀���p�6��)�&���vN�Tt��Ӈn��6+@�z�x��q�h��K��M]s���[ع�Ii�yE���0�	Sv��Ƣ��c  vI��ᒛml�D�k����v�jBd��8��9'n��W�v�Y�9 �[�6i��pV�gv6��S:n��׳�sZ�N�@��zn&Byi�d��qe90f����[n5�<@�F5Lú"�s�p���s,-N��C��c��m^S7���«���z1�mP�S��ݖ����[K�͌k�Hu:�1�
���^���+l��J0Vյ�[J��u*����*�Wc�n�m&��[�u� �6� � ��  6�     6�       m&�������5+�u����V�*������aR� m6m�  ��lL�1���
�(7X�� �*}��ͩy��Ln�k��V�K9;&r��ƻ����I���%���
��ON��u5ܦi_cU��e6h)j��r�-��.���;v�j�y�ֶ
U6&�J	�����ӥG��R����0����EN|
� B
�� ����{������^n..
)N�8:��պ5f圢^nݱ��N3��n^��8y88�3�yK m@Br����C8�˰���(�i&x8��M:����T����3���6��^�<Pr ����[n8��5�rn��`�ܩ�9M�9�8p��ё玶�7�B��!�[nl@  6� 2�[�'�j��;��4��F��%�i�5�p�h�w^���g﮲պi��y�G��"�U���Z�Y����hWg����{�������,!-_��{0�۳ �7q~^~����߱`�i�
���XY�ml���06������]��ޏb�6YUrZ&���� �ŀq���>n� ���K-R6��ݬQ
{�ߖ �wk ���؉{���5sz#(�n�KUr��wf��[��07di�{�QP��]Y`��u���t���e��g��-ny���hej�:�Պ�r�^�73�BKb��l�>w��'H�vF��K`r؈�Uh��sY.]k7$�߾ٴ�X�H� S�H�0S��N��nCӾ�`ͻ�DL�[�lL⚛D����Z�8�������&M����q`�ѽX�n+]���j�������[Ł�)���q꺊�RZ�����Wx ���^���5�ŀ�ۀq��ZU#PE��v���|h�\�8�wk�)�ΌqU9ẏn���������j� կw吾!I
HRB���iȖ%�b^���a�!�L�bX��߿kiȖ%�b^�t�5��L���˭ND�,K�}�NC�șĿ������bX�%�����r%�bX������,K�ߎ�����IhYVx�<L�3������,KĽ���ӑ,i��"P�yڰ^���ș�{�iȖ%�by�{�iȖ%�by���δљ���]a�Z�ӑ,K?D�����[ND�,K�~��Kı;����Kı/~�u��Kı==���m�h��sY3.���"X�%�߻�ND�,K ��xm9ı,K߻�m9ı,K�{�m9ı,Jw���m��KOs^	{ t!@�q�\�H�V$X퍨
�W.�M�$z�]]��"X�%�߾��"X�%�{�{��"X�%�{�{��"X�%�߻�ND�,KΝ���Թ5��\֥˭ND�,K���[ND�,K���[ND�,K��ND�,K�}�ND��2%���3�f�un��35��"X�%�}�����bX�'~�xm9��"dO���ND�,K�����r%�bX�u�.���5���浴�K��)"~���ND�,K�{��ӑ,KĽ���ӑ,K����8qd�BJK�ib}!B/���<^���.o��/�RB�����iuwE$�E��4m9ı,N��xm9ı,K߻�m9ı,K�{�m9ı,N����r%�bX�����F��$�kY7D�q���vt\���iJ��Rt"�֪�Jܬ�����x��X����Z՞/��bX��~�ӑ,KĽ���iȖ%�bw���ӑ,K��w�ӑ,K������f�u�֍]k[ND�,K�߻��!� 9"X�����"X�%������Kı/~�u��Kı==���m��.d��3.k[ND�,K�w�6��bX�'}��6��`!bX��w��r%�bX����m9ı,O;;d�o�D��k5�Ѵ�Kı;����Kı/~���r%�bX����m9İ����"X�%��N�zNjܚ��MkV�֍�"X�%�{���ӑ,KĽ���iȖ%�bw���ӑ,K��w�ӑ,KĂ� {���5���^����T��WE��t�S�\�f{�����:�;m��/<���tg[������㊣'N9��O����nV�<t���K���@�xc���g��r�3�ȷ%���8�6]�*M�Ƴs��w.��Ѹ�]t���VTۋQ�+���6km�!��ͽ�����5��V�  �	�*�S^�N<��v������S�BrҎة\��/R�o�K�����ϫ�q��(Z1Z��sV�<�y�pr�8�>��n��1ҭ���n5�k٫�w�,K���ͧ"X�%��{�ND�,K���©�&D�,K�����"X�%�ӿ��0����ֲ�ֶ��bX�'}�xm9��"dK����iȖ%�b_���m9ı,N��y��O�1r&D�/N��5�k%��qѩu�iȖ%�b~���m9ı,K߾�cE�bw߻��!-��,�@�.��0��IR�B��pI�/~���r%�bX�w��iȖ%�bw���ӑ,K��߻�iȖ%�bwߎ�\�Lɪ]k5�W5��"X�%��~�6��bX�/}�xm9ı,O���6��bX�%��w[NE3��<]���Ж�kStb��\��c��G�ͻN�f�!��g�T���չ�W��r�k!nkiȖ%�bw���ӑ,K��߻�iȖ%�b^��u���|��,K���ͧ"X�%���?�o�D��k5�Ѵ�Kı>����rD�F)�Q,K�}�m9ı,O}�ݻND�,K���6���0�C���~��i#��Kc�՞/Oı/������bX�'s߻�ND�,K���6��bX�'���6��bX�'�ws�,�n�՚fkZ�r%�g�"dN���ͧ"X�%���߸m9ı,O;�xm9ı,K߾�bX�'O���R�Y��k$��m9ı,N����r%�bX/���6��bX�%��w[ND�,K����ӑ,K������;.�u��ˬ�&�ѡ�)��Ǵ�s�n�K�jRj�������Wn�Km�c����ǉ�&x�������Kı/~���r%�bX��~�"X�%��{�ND�,K����K�i0�Y�Mf��"X�%�{���Ӑ�,r&D�/~��m9ı,O�~��iȖ%�by߻�iȟ���2%���Ӆɪ]k5�W5��"X�%�{�kiȖ%�bw���ӑ,~��? �����d���	�C`���bn'�7��"X�%��~���Kı==�;��0�s2�f\ֶ��bX���{�ND�,K���ND�,K�}�ͧ"X�%�~���iȖ%�b_{'g[tS.���\�Ѵ�Kı<����KİD��o�iȖ%�b_����r%�bX�����Kı���8��8{~�eȘ��!G���]<�mÞVN;&�-q�	
��/Sj㴷t&Ԧ��˗Z6��bX�'~�}�ND�,K����ӑ,K����'"X�%��~��"X�%�����/K4[�fMd����r%�bX��~��9"X����M�"X�%������Kı;����r ��bX�>닱mY-�!�s���g��&x��ΛND�,K���ND�,K���ͧ"X�%��{�siȖ%�b_��;5�k%��pԚ�֦ӑ,KB��w�ӑ,K��o�iȖ%�b}����r%�`qC�""@��� �s�	�r'~��ͧ"X�%����R�an�T��ND�,K���ݧ"X�%��"�u�f�Ȗ%�b~���6��bX�'���6��&x��g����uYk,n�UuQ[�:�!<�W\6#\�eS���5U��&� ����"p�;e��^x�<L�3���of'"X�%��~�fӑ,K��w��yı,N���v��bX�'��'x[f.\�֦e�fӑ,K��o�iȖ%�by߻�iȖ%�bw�}۴�Kı>�~�m9���,K����r�fjL�e˭M�"X�%������Kı;���r%��!�2's��ͧ"X�%������r%��<\��>��$v�m�8�Y���3�ű;���r%�bX�g�w6��bX�'}�}�ND�,�Ȟ����"X�%���3�f�uK�D�Z�ND�,K����ӑ,K��!�����%�bX����ND�,K���ݧ"X�%���:D�B @F��嚟�Y�L�f�.[�d��<�WV����t�9n{vN9�� ���j�m���/M�<�;�,�p�˳�u�ns�9��-��'g�E�8��n�5%��
ƞ��-���;��yK���2d�h�8ص%����6z�>}9���4Xۈ]y�ۇ���q�.��m���+��� l�6�h��q�ˈ
9��P�Xu0�p�f�j��������ww���_n�G��M���ŗ��#��l��y$ť*��]�ax彏]=��5��Iu��9ı,O>��M�"X�%��~��"X�%��u�nӑ,T����k!|B����-6�����e�jL��M�"X�%��~��!�H�L�b~�]�v��bX�'s��ͧ"X�%��~�fӑ,K����sR�ZL-ֵK�Ѵ�Kı;���r%�bX�g�w6��bX�'}�}�ND�,K���ND�,K�|t��t]M[�a�j���r%�bX�g�w6��bX�'}�}�ND�,K���ND�,K���ݧ"X�%���I�ن��35��sY��Kı;����r%�bX�w���r%�bX��_v�9ı,O�߻�ND�,K̞��(�?n�ų�����N�y#�����+3MZ[��E�mP^K�V�eJ�ND�,K���ND�,K�u�nӑ,K��=����Kı;���/O<L�3��:�'�$v�m��tm9ı,N���v���� C갡��8�q,Ngw�m9ı,O>�}�ND�,K���ND� �S"X���u��Y��k�%���r%�bX����ͧ"X�%��~�fӑ,��w�ӑ,K����iȖ%�bt����5-5��f�K�fӑ,K��o�iȖ%�by߻�iȖ%�b}���r%�`~Y�;���6��bX�%�ޟ��Zɒ�n��֦ӑ,K�����ӑ,K�������%�bX�g���ND�,Kϻ�ͧ"X�%��@���~��K�j��-[\ݵՃ����n�qd'f�:P�@j���!p�.�o�X;<-�{�̖%�b}����r%�bX��w6��bX�'�w}��<��,K�~��Kı;�����:.��u�֮�56��bX�'��{�NC�Aș�����m9ı,O~��iȖ%�b{����r%�bX����m��.\��K�5�ND�,Kϻ�ͧ"X�%��{�ND������${�	gڔոh%��C�IM2�&CR���)IB�rԘbJ`�3��`�$�I�BP�Ba2R-2\s3c�q3i�Y��3Mi<-f��2f�&l67����]��*$����$�+!$"�^�Ӑ�\a5�Hc�$���T�$4�ѡ�R@M�$.#6b���s�u�Ɍ̘�E��1��ZD�(D�,H��0# �$D�D��"DJc��<�d��F� �(�4�jd+S�qР���BS`# �l�#��h8)� ڀ�(�B!Hz��(���A׮�‘}D�x��|ӊ�(���'�AMɛD�b{��~M�"X�%��{��ӑ,KĽ�m�E33Rfk3.�6��bY���=����ӑ,K������Kı>Ͼ�m9ı,O;��6��bX�'����8�rKe�U�/O<L�3ż��/D�,K�,���O"X�%������r%�bX�w���Kı;������/R;//m�\�P:�#dװ�U]�n�!��:�q�v:<��nx�.�SiȖ%�b}�}��r%�bX�w��m9ı,O;����%�bX�{��6��bX�'Oz��R�Y��k2]k6��bX�'��}�NC��"dK�߿p�r%�bX����6��bR��7���D���$)i����M�Za��M�"X�%��{�ND�,K�~�fӑ,K��>����Kı<����r%�bX�|vL�u-&�Z��Ѵ�K�,O��}�ND�,K����ӑ,K��o�iȖ%�:�		�X�� ��"�x)�ޢ{��fӑ,K������|�����%3���g��&x�n�g�"X�%��~�fӑ,K���fӑ,K��߷ٴ�Kı?'��w�����%mX2���<��9���y�{��	5K92�2����{�}v��3l7.kR��f�Ȗ%�b{���6��bX�'���6��bX�'���ͧ"X�%��}�siȖ%�b_{�z��L�ԙ��˭M�"X�%��{�NDRı,O��}�ND�,K����ӑ,K�����ӑ?�2%��ߏ�\/(�$��eY���3��<[���<^�bX�'���ͧ"X�ؖ'�w�6��bX�'��xm9ı,N���t�E�k-�.k56��bY���fӑ,K����p�r%�bX�w���K�V���ٴ�Kı:{�gp����j�Y2]k6��bX�'�w�6��bX�����~��yı,O����ND�,K����ӑ,K����6bdHF�WG0������*����4�p�:*-�p�=G���+�w5��.��'��A)��vݴq�Ogt��vÎ ��jQtvh�RYI���jR�
�����ٸ�jW��,���(���!�/���.g�v��M�xu���ak=�8�郭�7F�qp�p+�d��mm��v�cW�]6 m�  h9���#Z���\p�캵3-$�f�hː�&a�W��C�m�~k���ɱId�����m;5=j|xD�t/v���"y�3w�{��^n�U8�Mi��Ѵ�Kı?~��6��bX�'�}�ͧ"X�%��}�sa��L�bX����ND�,K��?IxkI��j�]h�r%�bX�}��6��bX�'���ͧ"X�%��{�ND�,Kϻ�ND��$\��,S~�	���*�7uv]U�����$g{�6��bX�'��xm9��ș����iȖ%�bw����Kı<>�;���2��j\���r%�`�'��xm9ı,O>�xm9ı,O��}�ND�,K����ӑ,Kľ��z�h�fjL�f\�ND�,Kϻ�ND�,K��ٴ�Kı=Ͼ�m9ı,O;���r%�bX��;��Z��kZ�ִdtf�ZG���v��=N1���{�M�m�a���nWPIk�ʳ���g��&x�w;6��bX�'���ͧ"X�%��{���&D�,O{���"X�%����x�~,ѫ��Y���Kı=Ͼ�m9�tv"XYIdRФP�(�i,C)B��m��S"dK�<��"X�%��~��"X�%���o�iȖ%��V�v"�%��;fx�<L�3������ӑ,K�����ӑ,U,K߾�fӑ,K��>����Kı/��=ֵ�,��i��Ѵ�K�Ȑ2'����iȖ%�b}����r%�bX���w6��bX(؞}���r%�bX��|vK�XZL��%�M�"X�%���o�iȖ%�a�c���ٴ�%�bX�����ӑ,K����iȖ%�b_=$��v�L�j�їG^�pR�]v��jN���q�Q56�;7m�;|�%t��S<^�&x��g��~�m9ı,O;���r%�bX�}��m�Kı>���m9ı,O�N�h̹sZ�.k6��bX�'��xm9ı,O>��6��bX�'�}�ͧ"X�%�}���iȂX�%�}�����L�ԗ5��h�r%�bX�}��m9ı,O��}�ND��v�!��#�*���>���r%�bX�{���r%�bX�{������`jZ������n�q�����6��bX�%�ﻭ�"X�%�����"X��@������Kı>��d��Y��Y���Kı/�}�m9ı,?!{����Ȗ%�b{���6��bX�'�}�ͧ'��&x��������������U,,?�}�s����nnۇ��tZ!��dj����㥻��q�,���ev�Gm�<L�3ſ���ND�,Kϻ�ͧ"X�%���o�iȖ%�b_~���r%�bX���=֮��m����iȖ%�by�wٴ�@�,K�w�6��bX�%�ﻭ�"X�%�߻�ND�eL�bt�O�ga,�m�XK��ND�,K�~��Kı/�}�m9�lK�w�6��bX�'�w}�ND�,K�{�K�:��u�ֲ�Z6��bX�%�ﻭ�"X�%�߻�ND�,Kϻ�ͧ"X�g�K&%���Bii)��H����%��� $c�.	$H� �RT�X���j��G�I��x{��o���iȖ%�bzw�o���h̹�֭˚�ӑ,K����6��bX����fӑ,K�����"X�%�}���iȖ%�b~��ߟ���V9�����%�����K�6K����[��@�W�Ė/-�+	a]q<�bX�'����iȖ%�bw���ӑ,Kľ��u�� �&D�,O����ND�,K߿~-Ú�rkE��ֵ�֦ӑ,K�����"X�%�}���iȖ%�bw���ND�,Kϻ�ͧ"Ae�H���KK.�0�35p�P�B:��(@�'��
�<����r%�bX�����K�����b�E��tU�*���_��bX����ӑ,K����iȖ%�bw���ӑ,Kľ��u��Kı/ǽ{��fYm��L���"X�%����fӑ,K�����"X�%�}���iȖ%�bw���ND�,K4��$��JS��YK2�U�ݎ��������=��!�6W<�ڽ��֛az�\����uy����I$S��j#�e/;-�,V%T �\l�h����E	zz��mu�W+��s�2�[��)��Fk,�V�C�C�ޮ{NV��g�un͹e-	�c^lN�D��;l  6� m���ST�Ls�v�yj��͖����앴�qS� 8L��0��d�f�F�sZ��2v�}P]J��S6��]u$יX%���^�����}�I�1,�m�XK��O�X�%�����"X�%�}���iȖ%�bw���ӑ,K����iȖ%�b}�zIy�Vaun���]kFӑ,Kľ��u��Kı;�{�iȖ%�by�wٴ�Kı;�{�iȟ�DȖ'������0�r�kZ�.k[ND�,K�~��Kı<����r%��XdL����p�r%�bX�������bX�%��\���[�֦\�ND�,���L��s��r%�bX�����"X�%�}���iȖ%�bw���ӑ,K���Sq{cqڛ��e�����&%�߻�ND�,K����ӑ,K�����"X�%����fӑ,K=��]߇��P�z���E�iU������9ml�Uv�X��T���q��nn�kE�33Z6��bX�%�ﻭ�"X�%�߻�ND�,Kϻ�ͧ"X�%�߻�ND�,K���gp����L֤2�Z�r%�bX�����>N���ݧ"dK�<�fӑ,K��w�ӑ,Kľ��u��Kı/ǽ{��fYm��L��iȖ%�by�wٴ�Kı;�{�iȖ?�F"_����r%�bX�����"��$)!4���ˤHT��ȉ�2�X�~��?w���"X�%�~�kiȖ%�bw���ӑ,K����x�<L�3���@��VD�v�c��ND�,K����ӑ,K��0�~��yı,O{��ӑ,K���i��!I
HRB�Ow�r�j�lDfúoH�=�����ڽ��N�k�=d��UW-ӫ�]Y��Ͱ�R#_�w����X�'����ӑ,K����iȖ%�b{����r%�bX�߾�bX�%���s4S35nkZ�s4m9ı,O>��6��%�b{����r%�bX�߾�bX�'�w�6��b��g��w����qڛr�%�����bX����6��bX�%�ﻭ�"X�
z|� Я�|��h0���v�J�B�'�bC$
�U4�
��qW@:�6|?xa�D�&k�xm9ı,O�w}�NE3��<\��~�	T��[uIe3��%����3������bX�'����ӑ,K����iȖ%�b{����r%�bX�>>ݝ�jZf��jCWZ�ӑ,K�����ӑ,K��G�����%�bX�w��6��bX�'���ͧ"X�%�߻wl��52ۮ���u�8E�-�t�v�"����h�&�Z�z+��Ve0x�n�����{��"y�wٴ�Kı=���m9ı,OsﻛND�,Kϻ�ND�)
HM�h}E�$*fj�Dՙ���K߾�fӐ�r&D�>���m9ı,O{���"X�%����fӑ?�TȖ%�ߏ��50��Z�jk3SiȖ%�b}����r%�bX�}���r%��%����fӑ,K���t����&x���zǝd��ۙ�5�ND�,Kϻ�ND�,Kϻ�ͧ"X�%���o�iȖ%������n����T}D])G�<D<����siȖ%�b_��뙢���sZ�˙�iȖ%�b{����Kı=���m9ı,O3��6��bX�'�w�6��bX�'�{(~����<���k�EZ��ˎ9Zx�$��Z����kN�ޫ��p��5r�6��bX�'�}�ͧ"X�%��{��ӑ,K������PG�,K��߻�iȖ%�b{��/0ɚ3F���4\�jm9ı,O3��6��bX�'�w�6��bX�'���ND�,K߾�fӐA�,K�ӻ��MKLљ�I�u��r%�bX�}���r%�bX�����r%�bX����6��bX�'��{�ND�,K���٫�3	n��e�ND�,K�{�ND�,Kߵ�nӑ,K��=�siȖ%��*�=���ND�,K��^��D�)��,����!I
HRB�{��r%�bX���m9ı,O>�xm9ı,O}�xm9ı,N��FHI$a! ���/���y>�>^{z,�
�� ��b>�p��f���c�Jɞ�g����*H�����
�|9|���<�,#|YH-	Y|���o�2I5���D&$X38Ù�R^y2��,����6� p�	q����sy��ه��|�X(�|�q��1��I�%ʄ�W��Tپx�,�	s[f����1&��0�t ���<	����͕|�
h!�M&$�q!IS7��{
�|�%%�=)	
B`ʐ��� 	�q�V �0#D)D�n�L�R���1Qp��Ot2 3���:��(hPՁ_i�s~�332�m[\ �p  �BBD����6�=m�D7F`x����xllt.���)�����sP��L�Nk�F��cd�/A]�u�=;�{nzP닳���(�kl�ϗ�1�v]��\����F�Y��ܼH&B���$;�õ:`�q���n��sr����^n��֌�������{8��,5C�R�GC�v80g��8q-�Dv5�0����%�ۗ����P�kfr�9PU���t�1���c��-�M0��9z.ڦ8q�C�w���������ʛb��)�����;�cn7�Y睗r��6���8,3�lt�n��8;-r:6(�n:��p��d��n|[T��lH;��85�7k\1&۲�F�Z.�&�Y±K����,�pr@2�.yiv	�Ď�%ќZ��TM����Î�Ks���`�]�fe�s�b��S�B�	�v�1 E�w.M=��A�avv��SԋG�6�[��rݴk<ι4=�����vw!,�X�vmNr�v�5U�E Ҭ��s���UҊ�ֶUH���r�K�Z�E=j٭�	�k�V�8R'�Bॵθ��8�˛s�N��߾���s�.��X&�ۚ��&B]b���f����%��*�Y�ȳ�Iݺ���s���	���$�ٲ�����M��m���{+Ŏ�=]���vm�W;�b���sg
9��B�^p]s=#c���W�37V˲�v�y�gt�T��.��꺧ۭ��!#��m@"�O=Y�j�k ���@��/�Zڨ-I\Z i�l kX �@  6ٶ�    m[       mm��ck��x�ݶ㜑�k����:������K5�� �6�l #���)�)��)���Ό��6F�J�t��5���S��8Dg���Y��{��e���.z�o!s�%��ʲ.[�.�6A�*��,d ٠6�G�J�9�X�ku'BZ�Y�%ֵe׺ �Q��Wj��k�'�_A!��Q�	P"��W�/����`*x��������o��l���rGn��q:��OE�&5�஍�y뛶\�.�qm�a�q��ٰ���ൎ�tI�u�mƜ�]���[mI�-���ʗmp�p[lf:���n�a#����������;e����-�� �K7�nx�cV�<��Ѻ�Y��=i:�r�]�v��]m�   ��ɦ�h�#��D��@��j�\v�LK�"�����ۻ��s�:~~z>~�t�l��6�Պ	3�t�Jt���{��ѫ
��;Il=\����SZsS�{ı,O3��m9ı,O>�xm9ı,O}�xlD�,K߾�fӑ,K�ｶ��[3R\��kY�sY��Kı<����Kı=����Kı=���m9ı,Os��6���bX�����Փ35nk4e�Ѵ�Kı=����Kı=���m9ı,Os��6��bX�'�w�6��bX�'����e�e֋eֳY5�ND�,�2'��?M�"X�%��}�ٴ�Kı<����K�K�{�ND�,K�z]�:�f��E�f�ӑ,K��=����Kİ��}���O"X�%��߿p�r%�bX����6��bX�'��������kl�U��ݛ0ے:y뜝�p��UFebj�����=����{X9�ݣ%ֳi�Kı=���6��bX�'���6��bX�'�k�݇� '�2%�b}�w�m9ı,K���髚3	n�i�WZ6��bX�'���6������Ǡp}A8�O"X��k�]�"X�%��w�ٴ�Kı<�{�i�)bX�'�������e����f��"X�%�����iȖ%�b{����r%�bX��{�iȖ%�by�{�<^�&x��g��w��'@�[enW��Kı=�~�m9ı,N����Kı<����K�K��y���3��<[ζ�ꍒ���m��iȖ%�by�{�iȖ%�by�{�iȖ%�b{����r%�bX��w6��bX�'��O�{3.O�Y�Zs�uutc0���!��<���p�[�Z��o*e�o绸����+VE��w���K���߸m9ı,O~�ݻND�,K�������<��,K����j��3��<\�ߓqG��۲�ՉȖ%�b{����r%�bX��w6��bX�'�w�6��bX�'���6��%�b}�Kw3/L�&�.�.�v��bX�'���ͧ"X�%�����"X��h0���T�H � $R�A����)UQ4��"y���ND�,K��ݻND�,K�ƻop������FK�fӑ,K?(@Ȟ����"X�%��߿p�r%�bX����v��bX���}�ٴ�Kı/�Ο��h�%�\ӣWZ6��bX�'���6����$����;�{8�o }�mZ�K-n�+��v�т�����pk�ׁz�YۂB,.�w�{��]��:x; ��UZ��{89]s�w���G���, �;�y�Wm��W�}���x��L����ww�]s�ID������A�e��J��{� ���X~�x����`�޼ �u=�J�;e���S�#L�!l��L>>_%�E�p��C{���'�}��2�2�D��Y�fb`mI`n�J`oti�푦m�~I����4���9ˎ��ɋ�DU^�#��U�l�q��e.u�Ŗb��`n�J`oti�푯����|�zL�T:��F԰��#���`{di��ޅ�7o�?����/�_��M����ʰo�ذ_��a�ė��ro^�oq`\���X�Dn�e�&�z�ݾ������+��������<��+���`}8� ��^����ŀ}<�+ Z$�{�����~����8��mֳɋO�T��\O[�(�toۨ��^Nw=vs�S������7f���v�k��d{V�nM��$��q��V��g=�״��γ�+��v:d���"9�:N�Jm�,&��gQ�c�A���&P:-<N�l�k��ݻY��vM�9��s�Dx'e�)���  l�uN�\j���bܙ����gj�7S�r��.���~����>�'&�rݎ���x{H:�7^�LF��t�S�Ge�j�9[�Ͱ�R뼭o���`z��l��L�h��+	eR�嶬߷q`�sI�}���sqg����w����,��e��Հ|�zL�5���n��;�X9�t��D�¦II�}����ŀ}��`l���ST�,mGU�Q�^���X�������0��׀w��l[����9-��ݳcm6,��[Of��O�ϮF[F���5N�N�y����-R!��!e^��;�X��i0r������XM�FYv�QS5VCY�7$��ߦo�S �$��$ E��"6 ~`��'��
_,A����{�Ll�0�"���(�mi0��׀}�7�����>|ޓ ��k�Jݠ��!%lލ0=�4��oB��Ҙ��%a,����V�۸��������M��>��� �Fݩ�Y<���U���5�v�{\Ά��k����)��m*��l4�&��]M�,�����4��N������#L�UawQX�^,¦II�}�������>�{� ���&��7DQ�V�v�ﹸ�$�}�sF�r6z��T��Az��DD�\������
�9��� >�N����r_	\��I���Հ|�zLv�Sw�L]�!�k]U������ޅ�7o�07�4���� �@�slAVJ��Zx8�jYu��)xi�YٜF���v� ��[���~;�y��VeU�^�;�~��F��`z���>�rWk*�[T��J�����-QGwmX��5�s����B����ISR�Kh��`~�q`�s\�>�s^���X�n��䮢��Kj�Ԣ<�Wow�Xu����ŀ�:���J��Ns���7$���4H�AUiiS�`}9� ���X�o��k ���ح]��T��uE������ B"�{lݷk��DC����8��tկВ�k`�&UM���&n�n��,�7� �{�5�%
>��i�����VF;��U�{��,��0��׀{�7~^xٺj�2�7$t3106�?[v�S�Ѧ�F���ꖱƛ�H�,�>�s^���X�o�
yM=��Mʹ����e����/)�����#LW.��ߧ5�����i���'��24�����UI�	�T]���ݱ����p��ۂl����r v�w�{��.��W�#����շ�_Oo[�l�K�/�L�Z89ٹ�+0�/<�9ȩƣd{M�ћ��f��1�WE�1�)dy����js���(A�kn��ǑUy��` ����ͺ���*��g�:���¯��D6
wn���>����쏽.8���ݎ:5K"[���qٺ�½J�Q�n�Ԫ�]6��Vd���Yuq5v�_w��u��W\�P�(��s{����7m�*n��Kj�=Z�[v�S�Ѧ�F��Q��Eb�x�TR�������L�_�B����`��Հ5�I�L�7eM�UfS�Ѧ�F��]-��})�oƭ��1�,�"W*�=�w������u���u��8݈C�T�Vۆ�4vp���Ezu9ln�MӦ$�D�`�jt�I��F�N�mRY�}$���[v�S�Ѧ�F���UE-c�7l��l�>�s^T�Ką�B6T�)bR*0P)�������>Q���y���;��ŀz��f~M�Ν�]���c�+.p׸���,5(IL�{������o�%MIk��RZ�;�~^y9���0:���l��Lލ0=�
�WT�7Il�ڰ_�l�>�s^Ϲ����,�G(NwU܊�ewb�(N��{iL
��.3�v��^ċd��q+�j�׽�h�<PUJ��c���;������F����\�H#
�+2겂�2��`{di���K`n�G��ļl:���Z�m�\�I\� ���X���aH��svQdڤTUi x��ClKAH54���.�9Jb�NQ���@���y.��.�A�2�Fh�3|���9�0��$����Dԁ@�aA3d�K&\q�X��@���i�<I���,$a��RcQ���B@��NNM��\�pe�v ��A00dc����	9�E+Øq��s�%dP����֐1��X��Y$�mi$Px�~ <AO�A=T���ʂE1X��8��*�Q�Oh�� ����>*8}���~JUK{L�`w���UUV�(��LV�[v�S��L?|��?�����S}R�8�v�R�v�S�Ѧ�F��]-�����~[��v:ڹ,n��3�l�+=�8鶮uR������fʸ#:4ik���X��ssW?νŀ}��`O]o���u�� s�AISRZ�m��߷qg䒪6�O������0=�
�WT�u6륅�`�.l����?y�^7�7������9���TR�dpj��=	(��^�νŀ}��`l$�b�A,`+�$�1�(|��X*�f�srO�;�&�ʩ����wx{׋ ԗ���_���}��0ﹷ �k�m�lNWn�\�(�&֎�^�-��E��B�:�������\���X�-q��NZ�$��>�{� �t%�ޘ������Mf!ULՈ���`OX�?D%���׀n�`q�Y�	$�C���gUYsR�n�R� �7� ���Xw�<����>|�ـsx�%v���X��[��Ğ���������a-�n��ӥ����Rڰ~�ŀ~�%�Ν��w�o o� �Bi	*%DD� �Q�P�CkP���:C��#TҔ`��I3Z̶�ۜ�N�qcI���;�If�u�;���)�ۓv�v�g�I���NPw�w>�����c23u�/U��YFwij���3).�2�\�ӫt�;]��;\��T���2n�f��2���\s˜�����#�[�U��� �E=�!�u����L��LM�[l�   F�J��X��\�𧲝/i�E������k�a�[��A�� @��y���s+�]����EZ𪳒�r<4��Ik����j�$��.4��Y�*�ͷ���O�`�1�'F��`n�U�VEb�Uw�+
�-�n���`{dk ���0\��"����!�p��`q�X~���X޽� li�WnT媖J�?�x��{��:�ӱ�n���`w�)��*���Uݬ�� �Oz��u�,�7�6����w��䝳ZF9⪬1�؝��[	H\iz��Y��S���ۮ�BuVe����7zcN�0=�5���z���;0��e���c���-�7�~ٿ�P1(X��� W��d���X�t��s�����Ujh�����.�`q�X�1�J�l�7� �w��~��3!j��eݬP��[^�`{��z�`�`n�U�VEbŊ��R̶��z4����V�����G��p��e/&�"q�f�j#�:;���Y*A	�����������_m�95�b��޽ŀ}��`x���(�����xuv���rʂ�V�۸��%�2l�=� �^� �׋6!(^J��5~C�jm�!�ڰ�WL ��mÁ��B��H����XB@�#Bh�D������[i���4�$B�TW�����SJ��6"��^��{� �����sf��,��W,q�����ŀz�w~_������΅�YK�tΩ0�'*�.�&�#�Xm�%�3��\ڥ�K��e�m4�[�V-6������0%j���L`N���Ч ��j��]�`�[�:�K��@o}x�}� ����%#�&n��T,YYw���yl�~��`{di���l�5r���rV&�m��J��{� ���`z���OJ>��QJ����G�b���5�lE�t� �W�j����Ӌikq�W-�Հ{��`��[��z���ŀq1��b��%�b��9�ngL7��5+��UIm�S�y���߯wu��t�qӭ�'I*���l�ݬ �:� m�X�o o�Z��X܉�d�B� ��m�7�i�푦����VT�ˣU��]+����o�Ň�G���O��� 7{���6
LMI+��,���7� r�u��]�yD(��ߖ�oF����k�ڰz�fԿD*o}|���`q�X丣"�¥~}ݻ���o�W�͵\>T��Ւ7��q<���ġ��]�e>�s�&��C����0p���#�<�D�j��lqGTt��g�Xɮ�)^ۋ�@9�8��j�w@�f���-;9nc���q�CYԕ�<�����N�	���[�N+{s�F�ͤH�[챽N�$� � m&�]4�Ҥ�tuL�sX4U���:Lrآ��۬���n�w?�I��fy��������F^�U�٦u`���ƨ�0:�uҙ�sE+���}xm��>�x������`[�����(!�p�Ś�%�EQ��b�=>^�`9ݸ��[I[�r�m v�߷q`����L`I#L�E5��UU��E�b`J�K`�1�$�0��s��`x��>�cn�$q[0w�0$���#L	Qt�r+��Ͳ�d����.x�Δt�;b�F�GJ�v-�n�[ 6�j�5�Ȗ�l`IѦ�F������t����
LMIk��,��߷qg��$�F)�ͬu�s����g�""d�Z�$���)]�`�7� >��p�L�ŀs���s�n���V�UT��IWX�=���7^��>�x�6!/{M��:�N�a[j7%bhv�gF��`IgK`�1�����g~��Z�\�Rcv���P�K�Nx��mq[��E��l����w�����f�
�ZO��Y���L��	&,�8��M�o�%�`r>:����^,�7�6%2�-D꩹$n��ـ�����Xqx��<��Hԁ$j���R�Z_rn�kLK�-��d�ˣU媼�̫�`IѦ�F�.�[�IG�"*��^ ���Ub�UW6]X]]��>�x�'�/k��������o�Ϯ�J��]6wӈ{s=�gCv��#�j6)��J��P��b�.4��Mxefb`t��lw�0$���#X�q;!5�UU$u�ܳ >��s���L��q`��,�����
d��i�+mF��ۀw��X�n��9��f }�6����RV�%r� �XP��,�K��9<����$��q�����k�rN���3e�M�o�%�`��� ��͘�7�۸�ߐ �e��V;X�<�8f�t���<�9�\
ʵSn�jR�Z��v*����d�;f���0�n,ߵ�Ԣ�"9A���V���뛩-\�ҫ��ʼ��`{di��륰6��`o6
LMIk��,��߷q`�������`����Z�d-C��WmX6>l�>sf��ŀ{��,�pvBjq�呻]nY�|���$���#L�]-�����|!��"��j����y���W� RNk菂���Rsͻ��)L���M���>�h���V�<ئa 	|�y���4�M1eJЅ�O����T���f"�����ށu �N��u�ny;i�a)KJ�|0�H>�Dtk�9�s�2RB[i-��Kw�0�^����%Ē]�������f�}������qD��
�-2"hP�D��"$"�"E��R0D� ���B3%�k^^L���&q��Jx#�����B0�oa��}��tȀmr	��������AO��I$}��m�� �� �Ą�		)-�t�E�6ɻ�`݉�,cV�W��Y�m�;=��6�i�l*.�5��m�ݳ��sf�ۥW%�s�ú�B�aT"޸�!&��BT� ��)&N%�g.r�p�2�:�q�Gn5��-vsg\�<��X�/:�GzvU�nŬ�|Ǧ��z��}$ӧ�id���n��m���ۧW�r����x�o�TB
�#jc�T�+��<��\�M�2rC��dEtwk6�Ա�;j#í�cm>�{f�p�4鷜�#�'0j*X�vH{�y��"(�n�` ��ݶG������8.x�P�B9�:�����8p�� ���'d��;��:9:�.Bg@�.��R��ː�tl�*� MFʖYk*諭�).�T�,��R�PNq���V�q�+�j�W��ݹv�P*�sg��rw]�l7:����=��W��wX˶�k�$ͳ��in,�a��n���e��&�αAv�GY뇮�\8��<K.,=�-�n(���5FC8�ZKZk��J� �;5T��S<�5:%]�8�[I��m�sG�����f4S'm�7��j�������#q��j��U'���R�,�Wm��u�zI�nHZ[@���f�!��̉�nKn���$vۧO'�3K�j�iyyls������w|_\�/	U��t���*��ݠŷ/��+wc`�s�p>d�Weڤ��)9���6��a4���� �VԶ�ԁ $-�ŵ�u�&�v�j*^�F���Q 6J3�l ݶ -�Z��   6�         ��Hm���y��.��^�������܃N�v3�4�vwal�-R�P-��s��%�lj�b�)&[�X����U�&�5OA<���S�,��-v�u���N�Ӻ�̐�,�.Ҍ�֥nf�^�wG;v�,U�S;lV�P pY.��=x�����6�[6�����C��� Dv
U�:�$&�Dt(-��J� ����E�>��{�?��~++�O�&"r/K�lBt�,F�q�m�t��u�v�V�W�������%��K�s�ڞ{k-��4� J|f�] gXj28���Y�7e�y��%F�ҹ3�*�cL�Л	ͷ\9��q�����1��E<���[u%ˮ7;a���^W�)՝m��<� �Lk��>m�  y�$�(r6��q׎�z�<���W@�n���?;ݻ���s�/�
�W_�%$��^b�b1Ư\�{lݷmq=���:F��ѯn���V��AW�Y��oO�0=�4��u��[�0�\�)+q�![� ���Y�d{R���^� �^,ؙmj+�m��j[V��{0��هR^y�oy�ŀ}�� {��ꌩ��d�<�`moK`v�i�푦ۮ���k.�c*�X����>���:��{���=��>sf |}�76�Kb���k�n���7\�X�vm]�8�-�$��W��%MIk����߷q`n�[kz[��Lo)E�C�1���`�|ٜ�?����מq(���:�>�^,�7�5(���UD�8�򨥲7,�8���>���=�w�G͘�)������0v�R���s���ʞ��Ԕ)�u�`�[�)+q�!Z,� ���X�u��[���`l�!-Z��3��V<.�6M-�Qz�]`ݎJ&�Q��6i�O-U��:ܾX[j�7��� �����_Hs����BНM�87,�Gl�>sfuy獛��,�v��7���:�l�N�:�eVK�Z�����,�;f�Di"%9��G����r�����k �츪�*�르��߶�{�����6`��� ��Y�Ov��b�����������	��Ll�0<��+/k�ږy�d�Gl�`˥�8��r��'5�G
�Wmm��R�ɩqp��r�S3���lލ0=� �����"�p֊6�rV&ـs�n,���v��>�7� ��͘�j����\��x�ِ`zY��[���`qs�Q�څ+r�al�|���of����;μXZ�KE""vG����l���dr���6`ލ0=� �����7z+w�b(Yy��1^��b��O7j��.馓6�̢�t�'7U��8�b��d��W,�9�7���-���-��*}v�e�T-��`��L�%�g݆�`|���sq`qk5A�P�ZIL�G]`�u��DB��׸�woLxkf��I�dd� ��͘>���̃�Ζ����R0�����PVe�;z4��̃�Ζ��ޗ�l*~'Ps�kg����0�qB��ų�q&�:���ջv��(hn;M��p�u��v_#�hݺ�[��ۚw\��n��{]�%���GZۗ�|D�"��V�v���LZ�d���\M>���-������|ml,j�\���us�w
�d�Ϯ֎{غ�v�ε��7^�곊muۛ;l  6����|b�c�ST�M4m!���N�C.����J��s'k�����w�;�|����yz�-j���G;D{I�k�*eV4�!M$��}�3�'j�:��[��ȭ𲮁�m�`�9� ��͘>���8�Ũ�mB��|��S ���Y�D)��׵�>�ŀ}�l�Jd>�MtM�87,-�7� ��`{fA��}R��*�r��.������`n�i�����a�/�|���w��I�����KV��`����l��loF�U�)wE������Z��n�eU�z�r<4��L�UV!7g]J��GFyƘ�Z9r��K�v��ޖ���i���U8g����� ��͙��/W�ė�~N���������`E��@���� ��sq`��L;�M�ٽ� ���`ڷT���J�V�YV����`moK`{z4��ܢ1[P��_+%��7�ͳ �����z����=�n�>�c�j�[IV5OF�6[<�=�`����X��Ț���-��8�RD��d�6� ��͘��ŀ}�lԢ!}!���X�mQ�*�Y#���0~���=�n��9�`?�� ����)-t���Հsϵ�ܓ�3ߵ��A��^�S�֙"�(�]!�y��w7$��f���Y����8IL~��`�u��z�`j������ �lɴMM�*�+2�2�[���0=� �ߦ��傐qO$��A�$�;l"j��:Hvڭ�#m0zp�V��=y�B���il�=�7��t�7�gR��7� 7��R��+�[�eX�v�Ԕ%2okv� ���`w���h��R�,V�`�ݳ �ޖ��ti��ܻ��e�U�5j�f��T%	Ok�k �{� ��ٹ|R�y�1O�{Ͻ�nI�����%�:Y\� ���X�m� �SwX'�u�l(���GQ[wj�/#Ҩ���R��9-�6Ò��[�E-Q�A�CIdr�,�u
K]-��z���M�2�[���0=����yV��2�Yw�mɖ��ޖ��ti���tΤ�l�W[:���$-��l����0=� ��re�"�1n;J�� ���X�m� ߦ���<�s{pz��)+q�!���Ll�0&ܙlw�0=�rOM�p����H0H@���;{{ߝ����г��\��^E�]���w��I�I�/,�m�u�.�=���p{���gs����K�n؉�f�.M�k��K�m�@/ �v)<;����c��$3瞹�XgLŞ,@�tGD� xwc��;I)Ӯ̝\n9yj�+v����N�}��Y�L���rMJ�  ��4Y�����J�	�y��y���+�c��	ZA��Y��w��;�����z�����n��M�N]����ȷ���۪�����i4����ۣ�:t�#�N��Z�3/���2��L`{z4���� 9��58���T6� >��Xލ0=� ��}2��*ϧ֮��-�[�{�7��t�7�ɳ >��p-��<B���h9-X�I�����m`9�x	)�^��u��(<���"S ߣ�� ��m�9�7��t��"���\��R- �͗��I��l��\5q���h�P�:�g^�u0�9!Rr�[�z�6P>��b�=��P9�r`_.ThJ�$��Zܓ�=�f�$F1X�� �����T��7� ���r��L�0���R��(8�e�`s���_\����`rޔ�*̻�Yfe���}r��L`n�i�홦 s��jq;p$�m�f }�6��`{fA�6�e��WKW�gE	c���UO�:��m�p=��5&eؚ��u���+���޺�S����?�����ِ`M��lw�09I>)�]�Y�w��ِ`d�`�1��sq`�Ŭ�%qGe�����v� 9λ��a�b���@���!z��J��(�i"�>�nP�4#a�O%6�yu��%)u.�xV��[����l�D�6pp`G0	��G�)Ҵ��g#m'���=�"�c0��{����b���M�f���a8���|͓��=SzHo�a&f������>�j�,-�Op�]���VY��&�IhV�O4$�!�VFi3[B��d%"h�MhuI�ߣLto�{�P�m���g����Bq��!b3�n	3�͚�Z��
��/������LH��<�(|��Ѡ�~
���y�!�L4�}b�g�>rz>	M0���`�t�{'�C���P�B��BDD�N�!5���U��p�&��eg$�5�1�"��5�h�/��Px�i�� �(�cD4%.��z*���`�`|�hx D}P�P��߶���L�ц��S<		j��p6&{׷�q�ŀ}�l��
!L�^��Z�WZ�(��+� ��n,ݙ7��v�Sk��R�i]�)Iԙ��ti�r��A�㞶��"q��v^S�>[*v)T���JYGeX�m� ��9�띄���{� k�ee�(¯>�3/6K������L~ۦ .q>y�T�\�ʊ� �o�0=�`zvA�M���V}sʭ�)��n�9��w�L �w^�'�{�N4�@ 0%T%P��Q˞so k[�p
�.���j�Ӳl����0=�`~�ėz���	kpR�i+lU�6ٺk���n�M���:� :��=�Q�Q6؊ɞq0��9O@;��\ ��ۀ{�n.������z`�FQȦx�-��y�y�D)���,��L��Qή��֥�:2B��m�7��X�Ѧ��`�1�tR+���u�*$���w������ۀs�n,��kF*�B�_,-��=�ݓ 7zc��Ll�0?,I$&��-������?Y^�� ��U��s��v5�z\hWc�9�n<(d��Cn�&�N���Y����Ź�eK�<d;�Eu9��[g����B�>�� 6�E�)b�x���Ý��Y.(�'B��\��<�>x2�E���6��헢���ƛ���
.�n��bc���A�a��  fػ�u��`\��ͼ��|��J�Y�i�KeM�hV�#�I-��~�=�۱�/n���p���|�4i�!��\Zԥ��,�T�qق{Z������E��yw���1��Ѧ�F����5��7ʭ�7ev�nϹ��~�ŀ}�� �:�<�&N-{�U��mVIj�>�{� ��ݘwēg9��7{� ��5����#��BZ�y�`�1��Ѧ�F�"��U�x �/32��`�1��Ѧ�F��� �_p�Z�N��_֫w��+� y��\����N.w�#UPώ���7C�UXQvb�Vfx��Ll�0=�%� ��m�j�R��`U�9��l޼�X��[@#	Y`�U~QR��t/,�o��!�sn�9����kE��(����S�d��7zc{�Ll�09>y�T�\�K儳 >��p��ŀ{��,�Cv`�X�|���vWk���0=�4��Y%�ޘ���w���|�\�lUf:�k;XV8l�s�a8l���n�)-����\nW�t�Ͳ����������-�n���F�x��<�r;,D%� ��ݘ���`{di��*	uV'�
���[0ﹷ �9���Ļ��U��1 �:�PU*��~�vn�:�`���p�;<�:�� ��0=�4��}2��L`utQU�[���+E�`��� ��.��@9���>��� �v�Fآ��Z,��\;��s�dxE놲���+nN�Dݪ4�3c���Z�k�
9|��Հo��� ��m`wti�푦 ��w�^*�*��ay�lw�0=�4����uɖ����T�*�F���]� ����~�i���`�1�Г�����/.�10=�4��r]�ޘ�k��b��<P}h��_�͛�t/���;,!-X�5����x:�,�7� ؈Q�GIյ78�^��H���]. 9�\/f��m��MW�Fqԩv6\'V톊����o �[ŀ}��j���;��� ���녉�����`��� ߹�����<�Ԓ��P�|�����E"n��Z�<�ذ:n�(IL���`o{� 8��Z�B�_,�ڰ�r]�%oK`{di�7�L{�}Z��_,�L ߹� �����@�7��I���ٛ�yFFOQm�e� �w���������<q�k:���ѹ����Ô{a��ebϲ�oؚ��Y�g<���y�8�{s�=�ۗ1ٮ�<��n�a0���l@]=�Q9Þ�x6ν�=Y�bp��\��χ�*oIc���b���N�[r����SY']9rJ�<��Ni7F0�L�r�[nvۍ��۰ݶ m�  knyg]p+*��C����ܼ��U=��\�-;�������� ʀ�E��<35��)Mf�u�"��n[�uh�QיгAK�E&m�E��غs��GX�ʭQ���m�=�w��q06\�l��0:|[B��U����&�F�.K����ɳ�z��Ge��Հs�{& szc�#LN�0=�,���AW�Y�Y�l��0=�4����e�� իj֥�X�J�G,�=�w��~_ݧ�X��X�3,.��u�q�s�˔q��'�:�<��cM�*rP�W����}�'i�z��gغ���ͷ���Xu�9}u����Xպi7]Q�儶��6gW�jK��<�Z�
�@(�H�D� "�t�&bss��v�I�}�k �����<��l�HI|��`�\��x���w^��;�=��M��b�WJ�����4���L���vs^��	�RR��9j�$��e�[K�L�`EKC�ʯ�j���©Z�*��ݜ<�Dդ���HP�R�ܽ��^H�&r���w�?~�����4��Ѧ�P�@��ke� ��l�9��L�`l�K`r�b��-]`yFaW��N�0�䏄$%�򡏠,E����Y;�ܓ�߻����V�	Y��%X7�� �a%�:�K`wH�hR�,(��>˺����d���-��#L��m�����߮in���%ڹ���۪
�)�]����8 ��i�{O��\<�!%�������9�� ��q`l7f���|��0C�$�`��&N�06Y%�	�1����m
�b�W��W��z4��d��&��9�� �f���G]l���j���y�w;��׷�w����NQ))���B�B�|�`ɀfBI"F���("�(>^g}7$���'rY�� �̼2�2�ޘ�ލ07�����ܰ�O�!Sv8BV�lj��֗�!� �6�.ah��N��7�+8Z��]���9�� ߹���{��y��of���8Jȉ��<�U�>u��Q2wkgk ����9��f̚�Ν 2_,�ڰvu�`���0&�i�/rT�՗yW7X���{���ذμX���d�>���Uj�4ݤ�ـ{��Xj�[׼\ggj������"!$���W�j�����
� @U����@_� @U������P��T"$B(� T *@T""�T"(�T �DT")P���P��P�@T"�T!P�EB�T$B!P�P�P�P��EB$B$BB�T"$B@T$UdP��dBDT$B!P�E��T 	P��B �(�DX*��$B
�E��P�$B 1DX �T !P��`�B!E�P�P�DYP�Q@T$AcP��`0�*DT"A` �B
DX�0�
A`��DX�B�DX�B#E�DX�B E`�DX! B(��� @U� ��uPW�
� @Ux��*��TU�
�
��U U����@_�U�U���e5�A蛀D��� �s2}pK� �P
 
(� � �@@  h �  ����HT
UH �

�
�))�RIH )�D�   $P �H@�D

�$R�E �       (�1 ����{��Ξ[�E{�x |����5�1����}>N�. ��[���x x�.�y9�H�cr�/��'����0��G��]�=w��O���z^n�ۀx  S��� 

( �` 1�12V>�jr����� 6�����u�<��u���u� ]a��F�3\ �ɡX��+� 
}�q����W�.YN�6��< (�yN[�R����76��r���� ʀ   (M y_\m�x×^�ۅ�k��U��W8:�����y[�=� �{ϔ���.Yp ���vom��� >��=\�q���j\s��y���W���#����6�Z�ars��^�|@*�  ������O���ʹeͬ�t�R�iJ)`�ܥ)K�r�R��(�1���R�� ;r��M
R�M( ���R�14
P�FiJR�(�wr�R�M�K,�)K Nt�)c4�(�gJ)Ll�(�#JR��  U P(@�� �4�,f�R�ZJ)LM�9>�\ L�������n�7���� =7�m��z�r  3������� h2zN�e���z, =>��q���}�z>�ޛ���1�  !��ғyJUA���hb'�ڒ�@���R�4   ��R�yE(0� *����کJ� 4haF�ԥ4� �OQ?���������R}>�|?h��Ҁ��ow�� 
��@T�� 
�� *��@U���y��}��?��V��!YVA��$����4��k�s��Ѿm	��������l�9�[�/�1��7�(�@FIb�l aA���@�(@"E!@�i�H��d1 ��,c
�$#GC��	$�;�I?��AbI �bH���c$�]@ ��F0�"D��BF@��;� IH()�n���0���r���,���<�������8MH�:���$�H,�#�I�:iB�͆��� $dHT�0���{bT���"���D T�X�����f�َ�� @bH�GÁ �`E�2)]��S['&�"�
�RaYT5�!�1!��F���7I0��,��D��4^B����7�Ɵ�mD�(��V�eЕ��i	�!���`� I�!oF�����Y��,��G����V�~\��%����g��O!�f$`2�
Aф6���,����jv�F HA��" ��ư��B$B@�a��X1"E�@!#$	5Z2I#� ��.��;�l��f�Rjd�tHwRQ���#��$$h#��״�m�Ֆ�A/��M,I8�H:F6��"����V7���֮��8L��D�F��a�W|8���hhĥ4��<'!Â�(�8$��:�H0a.�Lb�|q�`JjCD��h��8,i���];%@�'hMZj�Ņ_�*�<��גg�l!9 #]B%�^>���Æ&�	$�kt�K�"@�Y$I�s�/��D�M�$BB��fM��cC,�C���MӅ%	M�9=u�o��sfXq%�|���oÜ�����đ���t��{O<�}�3e�5���7f�Y%<2#B#	!�y��=�s-,.����H�$|�F�t�D���'���Y��+x&�o�HFC�!K�D�$�4��,�M1�c�F���p�0���W~���4�3���2�i���O54m�.][�C�!��cx%RJwd�JIHy5i�{9<�	���!ͻ�����B��*Q�+�0��ZG�t��w��#�JYx4m���)�DȐ���caF0�@�5�AfYnK�1�p�O4xI��R�q�E4�A���~�y�N�W�!�l���y�]BK��.��d�aB$ �!HP�aF+d��o��65`T"���iZ� 0H`��@�`�4CA�# �(H�B@! D�@�$FA��h�
X�����b`H���A��,@�jM��썊@H�c�E@�H�A�!IH6H!$T�	LjA����e4nX�]$mH H�Te�b}ᴉ#]F��BCK
2���D�	$��E�D(�`�HSQ����ha�,j0��Ah��2��#�זB���-�ZR$4��@�ICo,�w!��$��CMd �����n+�Ԯ��8��!`'T1"b���Bk*,X��ǩa���$���~��%L��m����,�e5�o�ن�)�Ĕ��SN���H���`E�
D*m!U��L0�FaE�M;6�
hپ0���s7��]�׈�40�ѻJy�]B�N2��e��)��a�{���Á�:JŒ�Ga���!���h8�
kxk�^o{�Q��5�!����j�n<!I�"���=!<6Ji6m�p|<��f4 N1B2BH�Mzb{�p�d؃!�dX��Yt2!� �"s�$�0Hmp<aď1JHI�F:&ș!Á�H�`D�H�#JB�HyX���˿&xp��tr7�h5MGp�������4p�[NX�52��<�_.���|vT����ȕ���0u#��i%'0��
D~�&+g�P�/c��,�ޙb��պ<���<
(T�R͗�3<!�7OO!J��Iul٢�,9�vFH����y�����"@�oN����f�Z�0�m�1�9'�]扩��&�y.�:��LÚY�%Hky���Y�����o��(�M<9碌�cX!TT.L�"��E�՗�;q�Ҳ��IBD�$\�Z-Ev(�wL�6�rN>Cyt��3I��"�]b�<f�aYwJ��nhܵe2(]��7qȆ��R����eT�cB>a�W�V��4��l����*BF�!�T)	 1�u�4�M�DMoG0�#! B*V�Ji!�c�R����WH�ܰKF�[V,tȨF�l���x�%�d�o�gҺSf@,/��͔4{�%I[�H��@�=�^�	 ���@�u���v�5"R{�xl����]�����M�zz$�y���L1(C^{�֍�BO�H��g���nl�4O=�
��̈�F]�����j�*nGU�DT.���+f'�H�d�T��P�)�vuL�Q
*cr�j���mO;����ca�s�:��n�so���k��CgBFm�"Đ�i@֌]���|����4�g�^s��hԄ�xo�<��MH@�<��V�jB��	I*�H2k�5���I^�M�!	 Ć��WO��w,>��jA�2)��`@���
`P�Hd@���&�	`T$�-�T�d�$Q!�H ��	�b��H]^V@\.�����2]�&�t8������&��=����x���|z/���燇�$`��M����,��$���0�a��Z�Nmぇ�d���z���!H@�
G�=�i�i�L=�a�g9	d|�7#W���`mk�h��!�0.���t�o�Ki��%;�@��F�Hū#��M)��0��i�&����k�$l�Sb�ĩ���y����G�ߜu�>yq60g��y���8��xB�v���F<$}��u�_.���1�0&_CF3Z�@��ą!"M[��ַ��Wa鲾��p�C�_B V! ��2�0�t�(���"!��M0j�HH� ��K���e�x��$X�I% �U4��<4>I�$��xD���#tY�o��o�!XP��3���� �0�$8a7��!Hh�C7�S8D�.���%�p
H<��IP�Fς�v��(_JI����+�yQ� ���W��"ĉG�Se-�8h<Һ�)��&���%�c2�8g	M1J��2�۪�a����B�4[��5�I&�.�AB%�Ϡ�I�B���%փ�Z�$%���a�	M&��ׅ֧����aXV�|���{���6kF�kG<冈�G�x�kd�����k�����|6�� l==$1��_��[�t�7o��@�R�ZkfK+/v5��<=8갎��Fe��-պ�[!Iu�͕�*hٲ��[��,
:�ْ�3�1�:���Ȟk[�bQ��U0!B)dBBL�GI��"T�MB槆g������j��B�1d�	���O�Dm�QQ�$Wdd^ê���2�bO~ׇ��3��#\�E���bJ���mH54lف�hh6`p60.������G[�<%4K�6��(F�o�.�s>��Hm|�":B8B \Q�L���#7"֕�vy�ϜB2tcn�d�{�SF��6�F�a7��z{҅"�|0�����R��9!u�@甆���+!P�9�\9����BS Ⱥ4S����%�GI,
h��»xI�<=	B�]o�/5B7�&�����!� #do8:b6�p���H���1�J&��3~$�oG� �#bE��îe�0�7�*B�,-�]$����c`�$aP�!u�J��B���j4ƚ�7BB� ȓ{�H�E&���ѹ����YS���FHq�Z�p�d"I"1�H#�5 I[��!u���!	 �E�l!]����! -��P��[<��#t������ ĩ�	 %X��i�qݿ$ߏ�m�l            H�m�h        5�me�#��s��ej�J�݀�%Y;[M�4۲ajF�5����+#��t�x;j2� � d�M���,���sR�n4P2�f����R�هn3-E1�IU���,v�wM�c���c��
�`�7S�Z�+R�u�M�إU�ٗ)<��uN�����n�>�|6��M��m�6�lѦ�l�'B�	i'��j�^���@��6�e����DE�U}��}ʿW@�B\Cp`ͳf��HѶ�$���5&�T�d�KҨ�E��%� ��1m6ݖ�m��K@R��,��R�.�c�Uu��	���5<��V�@�t�ml]�A�{F+�*N�wjUۀ�
�%1��6iVU�-�yn
�@;m!�U@��w[����li�մ$m��ְ��@�`m�,�m� f�
m m��t�)V8%�j��e�[����� UR�ʬ�1��mPij�������+m& q#�-��9h)A��zt��e�zIm���测h  H9�	 ��m�6����9��Y��e���[4η;c�W_&u��l9a����QR$v�  ���N����h���[n��  ��zԖqnնV�86U�հ5��� �m��m��nS\ zĻv��� Y�t�$[g�|�| ^l � -�=�:n��b�6� [%����5�`%P*�PX�����m� p8 �h Fi�f�hZ�ՈX]Fx�T�P��l��m��gX$7Eɱ����U�նܯ�y]�vm����ݶ�[ҡ������o���;l���j`-��T���rҙ��^��m��[�l( �FA��m��ɴ��ēJ�jk5�kX^��a��m�:�Zv�	(�.��ۀ]h�i"M��4��g��h��춭��t�e�\mK�Ԅ�+�;%��h{t��%�Q���ݴja��
��座)�P9��::VR]�*��BP�S��a���H	���[vpgAm֗����@�X�Iz��I�m[mg@puvͶ9�[@ p 6�  �[n[[l���i�`6�H��tp �[v� m�h�Xd i�J���-�mN �Q�aؐ�@8 �m�  �`�$&����k5�� ���%W�Ur�WP6�m�S`����1mZm��^�l8Cm�8m�����6� 6�B� ԃ�E�� �u� �m�f�  6Ƞ -� l�m� �mpCKkCm� p��ڳ��@�e� pk�2�UR*�R�ܵ*է0Č�mBK�b$�`n�զ���   ����ո9t� �[qu]��l�a�6���p�M���V��Z�B�
W�� � �	yWe��V��ꪕiV�6���Uݪ�tUT��MK��2�����  ���ס� �m� .J-�oW  Zl  ��     5���   l 6���m� -���  t�\�J	B���Z�5� �ƶő��K[��[u[��'zX ����e�f�9ۅ`�'EݎZ�uUS�Ä�	�3J��U]t:K�ek��AɃ7��vZ�
����L���}����D���5�8S���J�mG��6��y�V�j��]U�v�j��y#�[�	V\�� p�� 
*���(v�M]R�����g����m�5T�6�m��V�: m[&�E'5��=m$��X#��U����k���$3lؓm��CE���0���É$�6݂U��@˱/0b�h��6�����w�Aq��u�R��0u�gB��[`�]}�z�ݑ.ރq�fP�0rt��٦��H;�xsYڶڶ�+�[J�%�5eY\���9<�a��e�T&���v[<ET�G��KJ�mT�l�S�l���������X#q������I��$�[�4�!g@[N[%]7H�q�Y"K�$��[��h����K։`�K�mg��E\t\Ӥ�8[BH�u�l���6ZH$t۬����ש�m��Z��cj�8N��Ph *.U`�T�6�6 �`$t��݀�kh-���l�UH�HL�K�sl����)eZ�%�^�:Z��۶-�)@mm��P��A����V��j�����YN8MM��m���%��n���@ �`-�  ��� �  m�� mh� [M�l��ۤ�~����� �n���#Nڍ� �p	e�Hګ`%��Sgm%�U�D��N����K�V�,d�i6@�۲��"�(H5Ҷ����`u�����l۪M�Al�s\N��!P��Tb���"�T��̴�,rMf�j�H��_�.��l%89^j���Y)P%Lj�iWjꀪ�xHv%)�(�<�U[U�V�9m�M�5�cZ�`m˳r�Z��"ڗ��s�<Y�ݣ�"j��:�ÌӚ]wF:	��T�]�L���CcuJ��nv�;$�p�퀋��v��S/F�ҳ�`�Iؗ*�j�qs=�����u�WGa����I�I�#�m�vձ�۴[E�R��Y�J��[��Gv��
��]�h�>8��nV��r5cSD�i��Aa%���Hz��[F@[�M��7��n�·����C�CU��r�k'Eƶ�e��Tݪx4![��b�^CizV�vU���u�J; )Ki��� ��l$I��m�"H�I��� 4�+l鲔t���)�Z�6� ��v�Q�z�6��m� 6��rT�M-֨   ��f]{[�m��[��k��  �m����v8	���'m����k�m'P�N��h 6ؗ��HmkZt   H@ n��  ��  l ړ�ڶ�-�h    n�-�6�  6�M�eꑶ�*� mM]�b�N�kf��K/2鈓��` z��`���k��eh� �h��$���  -�[A��ڶж����  @ H   ��ͱ�Q� � Hm� m�v݄��|���i�iK�kmC[F�r�V�UJ�ʵJ�ё�u[;T�Ys5m�ҩ�    9�Ŵ  ������׭��.�^�@��]�IX2p
��?/ʶԫ[uV֠&���\�-�[@� [@���an��m�kX �H�[[Ai�m�h �cm�� ��5l8	 ���h �ݶ �oP�l�cZ� f�[M�[@$� ͮ��@�Y��c^�A�     �0-�[@tk[` ,�RZ�ꗐ�T	C�4�:62@�Un�e�H ۅm����9�� om�m��� m���iUY�jUBj����7|;}��K��XԵKK�k]m[v��I$vٶ�ڶ>�}� �inI�ר������АY�U]P�//U���^Y]ٚ��g/g��W�uJ�cScJ�ݩZx[�h��l�����(��Lc�V�#MڤN���v2���N�y/:��e��ٲ�[�$�e���n��l$m�v��.[x�步X����[p��յm[W�F6�nF���0��n�w5�ԯ�t�ʁ =��Z6�g`6A����XYy� �eԅR�KU*�+WZd�([V�iB��Cu�*�G	��WN.f 
�(�����5��U�T4�����ql���i�	f�m�m�mzK��V��� �)3�r� ��[e����}�>� HX��@���)V����� �٥�;���`@m�m�4��	�  n�� �� -�� ��m�l�-�mv�߃�-��$HZ��V���U�VS�� f�1��68  �m���`          t�m�m�ƊkX8 v��	 T�UF�]U*�AU�l��lh�m�� īU!JU!5U9�H  _��T�c@J��j�yz~_�����خv��j�6�l�	<ݔٻI�YDG)�N3���w-۶۔���^���X�`U�3��JKUUT�&N����f�k��T�m���!��0[GK״V�^��.�ft�I�&�P�8��Z�SL�89��4�4�$��,� H�&�v��8^j�U��*!�V�om�� :Cm��m�'�n �c��j�8k2���pmB�����$m�v������}��UҒ���8��	��Q���,H�4ٺ�<E[}i��� ��慺ۄ�)�텽@8�ڒ�k$d����fqH)K�,�ڶ��I�
�� $���;� �$h�m�i�`��/G`$�m�Hm��f�`� mm��M�l��m� m�mjյ�����%� ,0�khv�L�-��5Q���A�����]R��NQkYq�k��|����*������8O정D���Q��x&���JbDF��SZ�)�(�0�Q&�<2"`(��a�+t�x�Jm��)���|>A�B�!� ��v.�4��z� ��"/�=H�0 ��Wg��LD�OUD0E�}L�(��"�����+�!��S���h؇�O�5��<G�F��SS�m}@O _%C�O ��C�}� ��Ҩ@�0���� `x��x��Q�#ศ�|�?�@C�<F �|�� AQCHn"F@�PGk�GS��~
!�@�Eq~Q)�!�B��>6(z�Q��� U� xhC�ڧ��1UB�q �O�"*���\E�@�C`'�
��x��_�$ �<�}}1��s�0E>�>�E�B*HB||W�6�b���b�!AaE1T*��|�؉�&���
�J�m��}_D^*�x�N )���"�\ 0���L������U)#�)�SHz��X z��� *�?�����A��X$�{ۻ�����v_򠥶���j����a�0��A�M�Zs9��sH��ۢ�t�kf��q f�,��dЩ���SO[F7$%�zs�]�=�m�K��;^��۲�6<�8ȯ �[<d�q<���V�l�m�H@ѱŬV�9;k�ö��E�i]�f��H���/0R�����v��P
���[Tr�*n���k-�u:�����5�Ů��v�g���t2mu	�8.&�y�Ξ���6ܮ��=�\lf�w]��^vV�$]@��΅`��*@-�Oc/n˱@.YU2/1W.�2F�.ZI�%����M��kXc�m�Q,�$��H��8�eg KU\�9Ij���V�vjr�It�]ϖ��n�Ln�1�����Y6�G/���mt8��j��dFm�O����z��Ga���'[���M�����ol7Y�= n�L��.Ɩv�jA��x3t��Y��	��Z�3\�QK�NXH��N�q��hU��J�ڪ�	�\a�*�p�{&Բ��ֶļ��,{Pt����c ��m[I�R�K�76�8-����Tmϫ"�u�73���!g����n�;v�hBܴힹ|rø�����[N���H�:9$�:�6������w��v�=*��i*�U�j�8C���5#cj�g���Pml]ڥJ%�搀h8��:H/U�D��cgMR��u\h�`b�L��7j�m�c�[V�3�d�����j�,��k��u�ی�0.$�*˒�7
d��V�Gk�C��y��m��㖎獴`��u���Q��{��I����;�Y;�]l��u�({rn��K��Ra6t��Wn�n9�ܪ�[ɵ��KUU)�*iR.[2 �5�F]f���J��z��+r�F;[�zKboK����s�^ٰO�=n��Š,=�yn�:q4����ڳnxz:#̇����M�B@�yxik��v�h�6�&^�;�2J���c��75��j����m�����hCZ�8������=�A_@�Q6��*�Q�Nn��}tힺ_\X�pV����si��wۅ�!��n`g�;e�n�����k��X4n8��y�X^i^���ʝ�=ShJ���:Mu��&�ۭJe���5f�s��յ���.��v:6�Υ� �ɻgkQ��vgln�����b ���2D������w/80)��"�{T�G�\��2e���Ԋ�{7l9�d���w^���rm��2/a烜�� *���ɹQیy�Lg�d]�l��Km�ku`ggJ7�q������`4o��7��$�;�)��1#�_ۚ�;�hz٠u�zǑD���Q�@�빠}_U��f���M �=R�dm�62crf��}V�w[4�Jh��hτ��NdM��	Š���Қ�����Zg���=�.]�v��g�7\R��k����G��Vl��� &��;WlNŪ�E��{�4[w4���٠w>���F%�B8h��m����>+��!�CH��Ϩ������f���M�,����F�Ew"�<��^ {��Ò�M�8�:����w�Q\�<$b��&�����Қ�w4����I	��	"�;�)�^v����}�׀uU%�.[<��ܐ��Ի�tUɣV ��5��K�ٶ�"-���Rus�+�cɍ�R<j8|��~Z��Z�j�>����&Y#d��L�N���:Հ�[Vn�,�ڿBC�N�n@wwn2����x��4��"���� �G#���V춬��%�,iD)��t��yڴ��Z�j�=Ϩ�n&���2G춬�֬�ڰ3v�`7���ݦ�&e�6{Lq�3�}��V�����ݾ�ڗ:�՜���"�4�[A�v՚r|����yڴ�Jh�f��Es�<QLQ6D�Z�j��f$^�� v�LͿu���i!pM��S$�@�t��^�i����-��-���<��H��F���^�i'>׿\�}�����V�a��!��;���$��'����hɐiɠ}_U�^v���� ��xU*]���}�%�w,�V�wc.������.���[&�i��͘�4t7
%�F�MH	̉�8������LǾ�����j�y���D�#����M�z�����Қs�F������G�z�����Қ{�4첳��G,	#�/���� �vq�{�٦�^��c��G��6EZy�V����~0�?M��u���;Ơ`�"hҖ�6�F`VPPVD,��!STHB�,�
H�(PRH�L��P�cJ����h��k7!Kӷkn��3�n��l��7/6:�ўL�Ϲ�B��`�ts�]�z5�\��PZB01]��jjܧ2Qy:���޹p���q��79�C��ui )��m����A_�����0�/�(�%U����\�Z[��:�jy ��gh�]l�mr���b#%����s&�zs�c���0�C��؉k ��wwS��jr3�E#
n�H���x;	:P���|ۚ�gP݋�:�$j,M�X�8I��g�@�^�@���@�>�@�h��&7�H�(�p�1=sr!#���`=��`ov�`��bP�4d�q�W�h��h��>W��-��ԑ'1��D��;Ϫ�;�)�|�W�}_U�v{��%"�,�4)���M�z��ߺ�_��IR��{��Is9�����4t��ƕz��ʙ���Ʈ�p�т�O5b�:�6�m�����`c�j��ε�@�׋��I4�r��9r�6�ה��Z��]:���	�D��}�$�}���$�^��Er��b#dQŠw�U�w�S@�^�@���@�^�����H�:�S�w8�?>޼Ϳuh��hm����I%�'�lr9�?,�+{������u�کJ�ڳ�S�H�.͒b܎p��-B������y�`u%�M�Qz��Zy�Z{�4���lIWI�q�8����g�bE�?����W�hg���cR'(��
�XݦX���H�#9��*]r���Zs�(��9�"K$�p�>W��>���;Ϫ�;�)�_e���DJ8��(��>���;Ϫ�;�)�|�W�yv�M$T�r8�w>�%@����Y�K��Mk/�eq=���Ms��"9xH�Fȣ�@�>�@�t��}z������(�Qco#�1ª����e���w��`w�����W�T��w��Yj+�I"n[� ��� ���@�>�@�t��}Ne�@��&BG&��}V��}V���M�=����I'��| g��9���*�r%���Zy�Z�̽w���_�@���@��Gdn<b�g�ۙƚ�������:0\�u�c�����9�Q�H��b�h���Y�}_U�w�U�w>�(�N� Ƥ��`���ꪤ���y���Z{�4첳�D�P2BG*��:Ձ��j���e��]ŀ�KE�,xH�Q�(��;Ϫ�>��>�w4��Z#�QƦ,MŊc��Vn�,z�,�֬��V�w忻�YJ��Y6���pi �Rѵ-k��d����}<���.�Ƥ+XԈ�Ojj&��s&�L�i�_�R�s�\c��,9�y}��U�<p%l6�Nu����l2!O��=�lqbΒ���yy8,חks.�qU<���� �FY�&d�Ɛ��v ���-�6����Ϝv{��f��ݕy+ ` �V�K9�566�a�S֍�0uf3�y�{���׻�{����G���ۖ�d����Zk��p�u�W*�/�x�3a�.�C9�ͧ&%4�_ۚ��������M ��$��Q�&I��}Ϫ�;Ϫ�>��>�w4��IƔJ"qh��hwJh^����� ��\�jD���@�t���빠}_U�w�U�w>�A���5.A�07�ŀ|�U~��}��h��>�CJ�5������K��6��l��<Y%���R���%�LN"%xd�)3@���@�>�@���9*�~��X�_3�ƭ�R�7w�ܒ{�����$HH�`@IX�HH@�4(qO��x�=��>���9�51cn<S$�@�t����M�����������(�p�>�)�}zS@�>�@�t��}NeQ@Q�&9����M����Қ��� �UI%[�o����Kn\�\���6�Gk� �pLhMv��c��#u�ݶh��IƔJ"8|�-��M�Қ޲���
0R7!�nG�~�٦u$�6~�`���}V���䎮�JĜs,�D�4�׋5�,�o#�|�%�Dw��s}�n���y�x�O!$�h9aPb`8�i�a��WlA�q^|���9(T"`�p�X������+�z^%} {Z��"�*y�=���Y���ב ���@�~ .��4b,Z���(ő��!6�t6�� hM��R�� C{�JJ&�6���:S|R	�,�
T���H@�����1�p�tl1#[	iw�0�(c<�t��z��W�G����D�R���V�]�}z�W�
�U(8�[�k�.I<���2B�,��"Q(��D�}�S@�>�@�t����M�ER���)�Қ��4�Jhu�ݷ�������0��-�36RK��:w:�&v9ݏ[�;���^�����X��Ŭ�l���<pr��Ɓ��M{�4u+�8�I0q��}z2�����`=u����2��w���j��2H�4_��w�S@�t����M������J%�4��,��,{L���G#�s��">����'�:Y�}��$������ڷp�-�p�?{�� ���/{8�_��{ψ��#H�O��y
q�ciٍRX�Mr4)���2�[�f�V?���@qț��NH,Y�8|��~4���;�)�wt��}�V1��6�d�'{�4wJh^��=��U!�"l�AHh��=�)�}zS@�����EGS��Q!�ӵp����q��gu7�zq�o�8�K��.�e����%˸`yT�v��T���||�0����?ws��~�
�
$!��#� �A����~��jkz�S�Έ��Z����9��X�n(�`{Es*v�u��ƶ�F�皕�I��T�mh.�k�3���m2,m4)*WL��Lv�E;�p�l��rQ^tk7��b.���{d�.�z�#X����s��C%Ǝ�; m��8۵`b��J��^�N�ьl�nM���x:��N�A��fa��ce�S���]��K4hjX�W�4�|���˻^\��\�n�e��awa�{\3R\۳B���y}[5���Ԅ,�j�H�.�����~�0�g��=ݜ`x����0ރ���r+r�d-�3��}�������g�����uƓ��cNF�p�;�L�1�3܌A���a��'��Xo>�n�˒5w#w�M��g���U/o�8����q�w��X��F�*I�����0�T�{>>��{���=��Ɓ�95dH�m��q�����C;�-����F����>9���KRU-��2ّ����;�)�{�S@���䪕Ux���� �{�-��wv�!�~�٦J�II/ʪ�l� ��N0{4�I$��r��\��Ȝ�.�~�`{�L:��vq�{�8��eC�DlɎD�}�S@�t����M�Қ��ōI�6� ӆ���M�Қץ4��`T�j�Smqݖ��Ev�bM.��q�{#����"��,�:���R�1�8��ɋ4��	!�l�h^��>�)�w�S@��Ɯq�,nD�4�Jhu��;�)�{�S@��+$�
IW*j��`f�e���e���lC�"7��/�C��,�i�zKCU�x���a!�w�S@�t����M#�QƦ,MŊc���=��0�I/ݹǀ~ޜ`��i�r��߿�߿���Z)���v&գV ��(v����-���H�s\q@�f٣U�G��{���{�4wJh�	c��M�2H�4��h��=�)�}zS@�`����14�"p�;�)�wt����M�e4�u͍ɏ4�@�{�4'>�L�s�w��^
���C�	�6��|�kxۉ��BƤ����e��i��i��i��#��5�.�s2��]�8�Y2x��Q�ݳ��w�Y�㠫Q]s��.Q���a���p���?Ɓ��M�Қץ4��,d�h�Hh����E�?�Y��>�)���51bn,S����M�Қץ4�Jh;��p�9��j8h^��>�)�w�S@�t��_p�*B��&I����M�Қ{�4�JhN�Q���mR��B�Is{��I�WC�+�pn� �F�s������$.�$w$��(u��;�W�ь�ݥ��c�|(����͖�����-��2e�էg�uN���	���ҫ[U�w��dW�h��'��v�x�s�%v�uջI�BM�-�A��a5쀪�N���y���j��7��ֶ��f	�/j�y08���sЫ��weȤ�]ޥU�*j���y~Is�䤮�(� yK���^,�<���[f��y�!�GM҉{K���#[-���_���i�=�~1|�ŀ�_��n�i�wn��=���?����ߺ|h��?Ɓ��M��˿~oq9��' �4~��}zS@�t����M�,��p�
A�8�����M�Қ{�4<�\���E�������Q`ov�`{���`�u�h���#q�6���IE�i���s:D&+���UsF�������}���d�!��~4�Jhz�r��a��� ��vY$$�N]�p�'>�L�=��ąB1��Q$WK��u ��s��d��~�$��w�%�UJ�7��s�68����0��� ��qa�$��J���O��|`�`���K�#!n�ʪ�s�E���ŀ��,=��w���q��r��i�wn7.,��f��U/�/���ǀ����@����ֆ�Hأnջ�݆3�LNq�];��&���ښu;	
��I�nF~�Ig�g�˻�仉��B���u��κe��w� �u��~���lr
��7p�<��L�URM��ذ}����L�6o��:+��%�j���'{��O<�L�PO�@�U5HHMR[UJ����|`��� =_�4�Țwd�K��9EHW��v�0?l��ww� ��vY$$��Q�@��hz�h۹�{�)�yS���
E$Q�F�c"�v�#v�����H8����J�Дl�L��F��6d�"p�>���-�s@��S���;�q�r���˖Yn�n븹�=2n��`{μX�L�7��ʷi����ܸ�߽�`�4��_+�~��}��b�??ۭ]�%�.&ӹ	�,�2�Ǵ���,3��B"�� @�.��ְ#W@qJD���9�rd��{~��7(���n�y��0�WԵ}����_��h�M˰\�n�$�#rF�px�b
E����#UR�%�'G�i�7.s($d�A�G����h��.����/���� 9oYN샖)w��f��$�;�q�~�`����U$��t�Er;�r�ˆ�ӌ��4ÕU*�j�v,�vq���q��آ�;�ԕ|�U*�w�>0���X���0>T��UR���ό��ѿ�����Ewww�/��-����}���<��L����V*	A��-JTl4.��������.����XD � � ԁ�1��=� ƣ)��x����XN6Ö�8���夤PN5
�p5�|���Y�ytQ"O$$�a$H�R,�>�HCA[�40����E���.������$R#D"�,0"H�EbA�	$E�@0�BHF �X�"�@$B	D�zmс��0�8�t�n�	S"9�\�k~s�[��i��2B@�$"H��	 �# �HA�� H�	���<�
:4�q�(Q��B�"�I1 �����T�XƁ�bl��5���!�;&�HHhe���RB0`a�U��0�ڂ@,���,V]BRBQ�f�����ʛp�F	�$ D�{�m��a���ۭΚّ#�	3�&2��
Z��t�k7=����u�v�eDp��U]F�<�[q�Z�q�l�������|���6�ڋE�w.��d}\H9��7V����ybSZ�Ms�=GY����댴�j1��0V�RmB��N�m��$ 
wJ���*d�[��Ԥ�Tz�`�]4iď'N��C�z�m�=*VSn����qm\����A=��>ݫ���K@�V��L�̾cSZ�WfT�X�gN�ċm�S����d�(:k 9f�Y�WJ���+�cݞ��©#�4P p,�Sl��V�i�SM�Ѷζ�f����m�m5*�X���v��b�Ѣ���m�9��vX�l��e�ۣV�r����v�m���]��ƱP/I��ns�e��%����=�r&U�<�f*��.�3��)M�)���y�N8�NwV��@��	�B�n�jT���2�0��;��8�:��3��*�ٜR
�:�l�v��kB������ٝ�vUW,ln�q�[@V�r;��t���ml>�Wv�j�qv���[����N��\r�����\�; ����--��v�4�z煴�0���*���Eẙ���c^�r���ʪ�B�� 7V�p[t�¶^m���ym����^�Ԫ9�!�"z�.�Eٕj��V��j�U�@�ЬVS�����H�;n�Z��[*������K�)�J���M�S���d�ad��"�1"O!m���9��!K<-�������lgE�@#�r/b�u�ol[)���u�����Bz��-9l�]_��â�!�^G]�S�-O��nĦrd�ڥ�T�5rk��#UU s�K��;�<򲝹�R�UUUUVVZ� y3(�6�T)j����X��tl5s��[������x�uI���c�㲍Y��m
{w]n����	,-'U���z��@V�*��L��1v���pl�dZ䑍\�W#�J�J�J�[Kԕv�Q6E� ���TO��x$|M�8ܜ�7����C{����̼1;���|�²�.�9�i�Ql&c���/lu���8�̈́���5��gc�I��n�=�$�Wp��%�ּ����+����n��ne2�=W$ڞ^'qE\�6����x�t����eض��%�t�v����YT��R��-O�٩�������nk��-!��Fm��S4�r�]Ƹ6��Y};���z����������q�$�E=4��[<��R.�lnMm�V՘�r/1��;c�
�u�-\fR�2]�MEn���������L��4��wv,_��;�Kr\M�$.�n��?���ޜ`����=��:㪬p����D�N��i�n��ê��7�8�;�q�}̡c �� �D�[n��t��m��>����qIB��������Mٖ�M�YM�w>�?��x��[�4�۵�NN�������r�ܠKn��ǡ(�tujusCQ�6���m��>���-�s@��S@:�2�����&HG�YM���/�%_�/߻�`�L}٦uRM���|�$Mݲ([�`�ش{�4�%]��>���=�뱼x�cN�J9��Қ�S@��SC�ww� ��sN�Gd�i��`�M�Қ��h��-8N�~KEF�8�4���헪�#;��t���;U-�a/<$�:c��{L�n����3��o;!�Ux�=Y�?FA�D��"p�-�s@��R�m�,�_�Ȅ�Ƴ�T�H�*2+%�X��� �٦�ʒ_�T*�Y�}m��.^.�y$NHb��p��O����l� ��Ł�~�4�jT���&I���t���˷4^��-��p:	���4M����ͲM��x��MY:V��qq�XNm]s"��6(5�I�6����m��{�4l����M�v7�Ɯ1��s4�Jhl����M�����D�D�ıG����h^��:۹�w�S@뎪��#�"p�>�)�����}�I^��e���PRt(�� `$ ���SJ��S~k]������d�d.��W�.m���/<m�_W��zI%﾿�Ē�*�I=�f1BU�-�3=+%�L�q�KJEm�;�ovf:�pu�-0�+7U����~�j`��O\in���K��ai$��fbIi��r#&RO��g�$�U~�H��#j8�K��y��*JHϺ|Lm��}���o}���T�ݶ�x-��Kv���x�gl�$���3��Lϟ���I?z�f$��.,�b�bi�2p��K��g�$��v�K[�f$���V�I�5�L��Q[�+q�qy�mﻘ�o�K�[��;Ԓ<��ZI-m�f$��!�4�UMR�M��V�×e�3��;1�N�t9�䛘�gY�2bݵ�r����f�v^}�G9e84E�)eg����Y�Dmq�FR[W��ݳ���{�ru�n'V	��ffH��v�t㓳�����j�u���3�Yf��W��:N�ʜJ�J�Q*�T�`�L.�rq�q�����\�V�p'[������6��,��0�"mIg�ꤲ�`y��vݦ�,�S���;:�&c�����r=�RXδ����>���[3Y�Sr�̶������|f$���V�K[y�G"9��K��ai6����j85.5dvGp���7٤Έ�D̤��df$�����Ikv�ĒKQB�A�B8MI%�߳�J��K��Lλ�f$���V�K%�ѕN$��xᑹ�|�W��jI.�i��$^���K�����%˕�E�c	-ˁ�����<��$�s��m����$���J����|)"q��a���9�kѬ�-�ɪ�	���"�7����j��H�dl21���$����ԒM����O]�{����$���%�W�,����(p��oww��Rj�B�)�!w���̓-�����Zپ�&}I%Uwm����vZj+wn
��1$��v�I�l�I!�2�$����|�]eѤ�"�dmc�7RI6홉$=�U��m��ė��>~�M�ܧ>j������x�f�4��K��6�FbI=wai$�v�Ē�Ɵ���U����e�g���ܭ[�a�t����y��l�%S�q�ƶ��϶�f(���$����O]�ZI&ݳ����gl�cm����6]���!獷��`g�$������獶}��cm���<�+�z��,�(��K�.6��{���Ͻ��ynHC�j��O�_s����9�m���I��o��z�
]��\���6�*�}����}ݜy�mﻘ�����J�I��~������˒�܉��E�m��i獷�$�v������8���7٤��z��������[j�D�p����,\��i��Jd�֞V�MH;MC�j�ɵ�ەB���I'��-$�n٘�C�ez")R��������ޝ��vI.\R�\�wm��i眩*K*H�����}����o}���J����S�5p���VE%)�1$�:�V�I��3�ə���[m���<������B��1�ԕ�ww�獷�ف���w4�����O ����S����鼶���|q�eح\!w�6�������ڶf$���V�I��3K�Ds��s���"r�M��C�k�]D�ml7�����[���R���{�7�c%b�{RT�u$��}�$=�U��m��Ē{wCRI.�U ��a�7�I#}�L�����6�of6����y��UR�I}�ˎ�"r�"�w	������獷��`c|�����獶}��cm��"�pV���獾�����-$����1$��ʴ�[��f$��w�]SV����������?���/;�X�I�{#1$�����Sp�8s�K��z���,e��퍻����D9��]n��kU�O ���\�J8���̝�냇d��=v^y{t�N�x��

�lo6R��<st�Vj�xOK"G]1QisF]�#S�nҸ'3�y��v�Ѳm�y�e�l��D�
YS���A��IQmlJs�Z7/G YQm��ύo�������s��\U��[E!j��綛�������q�Lu��ʫ�����?}����&ai۠�����_Mc�g�����o��A�8+�^����_񾏇E�#���i${��V�Ku��Ēz���2���8���oY��(].[!.mn���處�밴�[�_�Ē�*�I}�T�S"�ن8A��|�W��jI.�l�^���<��ZI&��Ē�[Z2܃��D�����*����<������~�������*_RU>�~m����Y���v� \�y�m���cm�In�~_�6�of6����y�m�J�Z�e��s<��Շt�������ó��l:�I<ܐ�
oMҔ��e
�]l�V$�o���I'��-$�[�}�w��;gm��㖮�+wrӗ�6����&x�!>�"&�����R0T>:���s���r�gvq1�߾������N�ۻ$�.)v�\�������<���i1����T���^x�w���ovk֮n8ӷ.ASFbI�*�In����O]�E���S��8�??Y��(ZA.6B\��w�����# �z�XmՁݖer�S��ZF��m4s`���ܒ-�	�:YE�9��zo��o�]�ۮ���;�� ��4����UR��I~����X'��˗rB�%�n,��,����n�����/�	�̳�rӎX)�� ?wt�=�wM�x�5�@ca-��&�Vq�Y"0%e�V�
�l< C��Г�!
�k������0f��1�y#h`2;�$�X�D�l����O�Z�B�3jB�)�4VB'���,����0		3.�M����5�"D��JЕ� dE�� �n1P�.��B��(�"���Q<ǂ>%4��ȃ��*#���)�G= ���O6�>� �#��D<�T�C{�<�a�O��}0߽���r�ܘJ��w��z��s@�����h�Tx�K�Iiˋ ��^��9RT���< ��� ���XʕW.�[�#n;��i݇m�Q���NC���[�
@q��9�J�n�ԒJ^f��$����ۑ~~�|`��0}���R������,���"��!�0n��h��`{��X�٦r���5�49�J7r2��7{�`{��X}K�IR�߾���}0=�餖F��\!w*�����,��� y��j�J��v��h��D8�9&I���z�� �T����݋ ��^��>UK��~oۇ����r����x��Sm��f��t\��ס2�3/�����;�E��	�����U���Ł���z9�c��x��XeƋ�wdP.��5�q`f�wrڰm���H����<l���#x���z��s@�ڴ�6~��wwb�7M�.��I%�Q�vۑ`|�ʩ_�g�< �ﾘ��,��w4]U���X�qh��0�RT��I}��~_����� ݽגAU8��(EX�
�+h~A�!0��@E]vI��%޷��W�':X�f���>��i���Cn�3�+����<u�9�7)n��H�g�B�8�v�"�蠴-R�r�gF����y.xy��r���^Ct�7V����m�,�+r�N�&����W�X�����ӭ��c$
9啐��)n��|Y�X��u��r��TvѲ��eԛg���aR����n��bʃ�1������z�5����1@M	2��_��KK3�m�*	��B\��r7a�Yr��׋�L������q�_���7r�"��w��74�빠Z�Z��4���cma�nf��w7�b����x������:��f���HڵrI!�`����ݘuRM�wb�?n�ŀ��5H�! )�����0��X���X����@k��Lq�L�NM�w4IR��������n��u����%V-�{a�jE�h;q���մ�b�T�� j��]�<�nh:]���[���S��1�j�[�DG#6�q`>;����$�▝�nE�y���/�F� �X��v#�T? ���߹�����X���,���ڎ�t�8]�+ Ǯ��w{��B]c�Ł�O�����f��u�Y.LW*U{��Pc�Ł�uP>DBO����3�FE�?�1)3@��w4��h�Y�wu��/Z����O�F��R���<\���)���/n�s�u��( �����4D��2'#p��>ߟ��@/���wqrU��ob�y���q�	q8����;���>�]���yԩ6o��q�Ȯ]�-ܘ�w�s���d�O�G" A���U�@�������$��{��}��DF�8��H�Nf��:�h�Հ�ݘI=���wawwrE%�q;�9�ou��'��O ��ŀ}N����%P��NH�䰖d�]���Ĵ5��yM՜AŇ�1�a/"K��(E��PmŠ�f��n��:��/�W������>g�T����Wɀ{��,�T����,޾��v`V.�$dX�Xc�(�hS����^T���ޘ�v,Y��r�2�ۄ���Oޝ� ;��{��,�D�NDW���d�s������	\��< ����:����x�/���ڴ�jI��D�r(�)�'[��C�6�sē����6X������;,v��$�d��q\�dP�rx�v,�:�h�ՠ�f�}�tDl���q�X�{��䪾�vo��� >��`���:�6o�]�ܑIq\N�H�7��+ }�V�w3]Ł�-�ڍD�;�wU&���n�b�<��Ł򪯒��>���>g�T�R��;� ���X�I~�{����<�O����Oh�H��Z$B uҀz�E7fw]���tk���H�'hv�l���~�n��ub�&W��az�b�{qٜcuR\�m�t\�ĕ]2s�3*�:C�C����0[������E��c�6-�I�0bl�@�(ץ4�'nQ�g�n8rD��wlV룴*��H.�]I�aƥٝ��vB��<lWd��r���ݻ$�Z^#ѹ��u�:C=�mu�zz��ݚ��5�6覿*�P���7��W����H�b	���Nm���[ݙ���w+N��U����>�jtv]�6�n��ߋ��[V �����,�rˍܻr�.,�����K�Wa�w� ���X���Y�6�����H��Š��4�w4�.���Z�U-q9�Fɐiɡ�[��X��b�?m��W�]����=[��652)q����K��z�V�u�4�w4
�\TJ1<J1őS�����3��\���M0F�´#W�|o���n�tm�$$s�$c��/����@;}ـ{��/�K��a��}� ߯��5��n�w5�n�}�ov����e��=Kw4Wj�ؑߟ������qܘ�v,�=�X|��z���~��hV.,Q�a�1G3C�����_s��ݘ����`�w�\��GrոF�X�׀|���~�o�ۚԷs@��*�KS�'���oJl��Vӌ�ܚ�St��On�Q����?����qƤq���q�۽0�w4��s@�v��UKdJG2�"��� ���Y�����X�}� /���������L�Cj'3By߯p�'�k�O� @ �@�(���%���y$����{����]��$i���'�vq��t�=�w�$����ŀ{�ϝ����q��� 7���>��{�^���-��h�X�5RdM��0`��՞,@�s�u�7JZ�vo�;\�25�����+�qܞ�݋ �}{� ���}l�>�]VHȰlŎ�� �}{�>I|��ٿ}>0���{���q{���d�E��JL�:���o�ه�/�U]���,߹�� ��ͱ���.9b�r��*o����,�s�~�$WA��M:V�țUID�߳L���y#w.+���L��q`U/�T�����/�w�>0��@���eQģaBL�H�d)�M�c:74v�+����Vک�[3�8M5/'TN�dR�ԙ�}z���Jh�g%T����ذ�-��Ki��ˋ �}�gʒ��*UJ�>ﾘ}�b�<�v�gԛ7�_;���qӸ�n��� �}�X|��U$��޼X��0v�W��B�	܌��L�%T����`�z�`����J�7��0ߘ��2,�X�9�׫��:����V�w�DL�Fd�b�R	��A��H|�0N.Ȥ�) ��xP�Gk؛�*h2����P�R
��ȑ� i �`7y	6f0����VK��!i��5������`�n��I��=��7�y�T E	������h�H�@ф		T�a�JE���F��9��lv��A14�޹{׽������56��UU����́���G���1GA�.kY<rU��� ����lPJtH��7!�Vvxs�anq�){"hV��zlaܢ�]8ZuȻm�8w9h4��H���nZ���p8���%'�QV�,e#����f�ݵ�\9e�Urj���(���i^��\�L�;�lV�շ��j��j�v��4��!c��]�Z�A���43��� %t&rk���� �s��hp0O/+#�i���5 � gAr�!{f��p�Ev�Kj��B�@��Y�[�U��)�<�$��Y�7  ک�v��ٶY{4���	�g�\��2�� �m�iN1S.��"]m�lT{nѳ��q�ٷ�0b�um�)��%��N�!��zw'T�7[87;�����<�Q��8f�]�j���	�0#ʳ*^<�+�F����p�'���&c��X�7M.8J��K9�Yݙ����H�=��I@l�!2�Q�d�3i�V��tOD�U����Q��	X"q3�pZPm��5V�[��[��ɛR�s�"zu�Y�[x���a�6�[�Wn2xֳ�7tA�Ϗi�g��I��d�� lؕ {b7kf�Eӝ�������A������N:��d�EPU�*�T������<��)�B��Aab5r�Ҩ�)v�Y��B+e���`�A�˅JQl#�gX�R��R�Of��%@	^nvػC1�Aת��k�X÷Qdv�x���@kf(.2�NV�ٵΎ�����k�݉�u��Ym�;Ŷc�	�c�����g��t���ֻ%��+���7�9��u�p�r>���k����ţz��*үWT9�>8��$k5��ic  ��M�]���h��8+����#lѲ�:㮬�[v&����O\�;^�K2���G8)���cs���I�7;'F}q���ܖLjd	ڻd#�sj9&"�(�5��ԉ=T>��w��D�&��/��Ѓ�|(&��+�}Q(����ڂ)�>�m)��a��}<�k,�w=vH`��ιfv;Z,�ƭK��{-�\�Kd@��p�%�l�4���h�R�yz�R�d��ݒ�:7+�]e��9Ğ��vA�Ϸ	��[p֐�Ż8�ab�h�6��ݺ�����r�XA%�G�l	��n���;��Sr��v�gg{wV���]q۟[.�ܶC�s��٣Y�ݢٯDnw>��Լ�V���}����\�S'2��K�]q*��|�%�T�۴��P�sF��wv���hJ�;�h�����ϼ��u`k�q�b��n,zZ~qqFc�'�^�hz�h^�s@�����:���["MI�6ɐjj�}�,z����:Հ=n���4��7�85&h~^�?�@�����v`u'����7��c�$rI"�6�s4������]��ߏ��������n�	�T�'�p�n���vã�_��_���M�OV��e_����|sn8��q۸� }�}0w�ŀy���h_U�U�H0ȓ�"ri'�}�"� *��N(�k�,�M�ŀ~��x���ͱ��Idi��\�� �}�ŀ{����;{��݋ ��{�#�!$,.ˋ�R���s���{���>I����`��a�e�,W.;� 7�ـtr!����;�鸰5�j����.���jV�����.�l3�'n^���-O��M�R��T����#_m����X���,ݽ��J���`}�}0�w��w%��p�;����|�U*l޾��t�=��Y�$ټw#�#�Iv���<z�� o�ل�ʪKr)�U�5  �@bA#�@��d~C����2I�~޾�!�޽�Q��-�e�wp��I���`��Ł�jZ�5�e���h�THr��l��L��ŀrUK�n_? ��� _[4Y�pO*�iǍ�Ԅ& �X�F(��)�xh�v��T�.U���nR�`�dX��1�#s4�GV���h��9*����X'���������x�~��T�M�{�0��X��y�T�����:�,�K�;� ;��n��þ��+�~�<�����Ȑ�ț	�iɠ[n�����'�k�H�TbD;+�1�=�Ƈ	�*�p]������*_UUR��ߦ�/���˗q�Y�f�����-v� ��h۹�|��_�v;M�q���E�����S�s�N�.�NZ^W:4�p�c��V]�{���-��5�n9#�M��������_[4m��>�,ZWUo"�R5�1�ӏ 7�ٟ%UK�T�+�����>� �ڴ
���G�$H�����7ٱ��UJ����� ��h�dX�Xc�F�h׫��ՠ����IR}��,��xdv�bq(������޻���eS�U⤩��tB� rK�v���m���ӝ±�0��� y��'�H]h�N@�k�ݰ��	�즊�vIё2�M��YH�:}K����V0j��u4�6�QO�[��s�ah+���.�ų�gkm�8�3��W#�%Ӟ�d(�G�m���pVU4s����Xv���6��.�Wm{nǭ���;�m�i�yg* ����՞���[�ˑ�#�R�⤿*��US<k��.)qւڤ��@���󎱪�4ۓj���F��K�F6�Nbw3[m��wL��q`�����%K䪿Xw��<���Y-�H��dV[�0w�şRJ�����0��x����IR�*Wgڻ��cc�G$��5&h�/��:��K����\�]���<i�وĉ�r9]kV����׮��1�u`u|�y���&�Z}l�?fr��0�k�`k�j��p��)R�!���{@�\�_&�;����܉K�s���hlWM�B�8�d��%��qܘ����7׳ �o�$�_RK������=��;�%���M\w y�����yJ�ٲ�׀~ݘ���ϕ|����=�Qێ8H���0����v`ﻋ >���-|��1���N-��_RI+����wذ����7o�x�kFȑ$Ĕjcrh���?fR�������x��f�뗪��ۆ�-Xs�vӔ�MoOS[�8�$��
�Dmv<�kE�e���.h�aЕ�m���׳ ݿu��ݝUT��;��`�uj]ˑ�'m]ۓ ݿu��I*l;��wob�7׳9$�|�J�Ϟ��_87%�,W.�ǀo�Lw�Ň�K�$eB
���������'?^��5���.hA"��;�ꪤ����`��� ݿu�|�{�0�m��K"j�V�
;� <�^��UT��o? ;��n����u�y.�c�U/Dʽ�wLv�s�m;��V厙˻z�Fl'����=S�$��ߟ���}��۳ ��qrT��x����`׬a�eܻ�rGq���f}UT�gv�, ����7o�y�U*I&�}�e�&D�Sԓ@�����^Vh��@/����uF4�QI"dMI��%I�{_L��� o�ـ���		R��6��� ���7�]�qH'm]ۓ ݿu�/�R��������`��@���1V&��<kȚ��\7lv����T��r� 9g.��3�%�d�_ɘ�iŠ��޻���g�ʪ�u�<��2KM���Ԏ���q`�:��j�[���ȏ�%Wg�m����v&�
;� =��� ݿu��g{�0��X���mGrܵ$��nL�T������`��,�R����� �Ё���[�G#��n��UR��������s�d����$�PB���� N�5�����t���l�!�1mh������u���g/m=v�� ;\ntI��-A��+�r����n��<)�++���u�qš�cO���R�]d�q�ֶ��+�<�[3kv�K�m�/V�u�e�N����W6��t�K�k��9*�Ƌ5(�jb��o���lc:��t���#R�S�ui��*��6�ue;7/"܇5�����}�����u�*����gRNT]ȳ[e��B��˴�M8.�Hγj뜌�ʦ��]�9��;�� ǩՀ��_Ds�z����ݸ�%�� y����M�׼���ﻋ>�M��r���CX�Rh�;�h��@���}yY�U�ɕAG��6�Z}l�7}�X���0:�O�o<����ZXB&�&H���w4׫�������[�#���s��9 �9�l��Z&ۯ8��" �n:�uΰ6������l���X�9� {���k���@���q{�Y#��$�q���y$��{��>  ����b!�\����y0ݽ� <�v�|�*�M���d��܊9ǀ�� ��qa�U$����u�<���.89I�1�94z�hު���h�����R����v��%۷n89#jݹ y����J�t�~ w�� ��w4�
(�x�SB)XБ���&��е�ÙBm1+VF��>������{���l��F�p�4Ԟ����@;��ﻋ�������s�볜�wE��۸��۳>�UM��ذ�k�n�U�U�j$ia�P�"rh���$��߷�՞SPd�m�D��%#Ye	e%H�et��d
�b ��;�22������6$�Kn�%B�
@�,HE���������@h@��/�M)��.�j����R��.����i���bHq63Z�8�p`P ��A��m4D4`͗���GF��M2����0��<������)�j0�Hlb;��N���N��$�������"F�,���v>Q�08��54"p��!Y@4"��)�6��Xy��O��#PC #�!��@�D�Q�x�����Q� 4����G9�3V�w]X�(��"�bjࣸ�>U�*Uw�����_|�}l�-빠\^�HHI�F8�jLv�׀|�*�*K�}���� y��4i�����I���1"D�u�f�f�O:�qf�<g����T��V���;a�U)#NH�Z^������+?b�^0��{�u���E�q]�r���X=N��Z��s~�DBE쿶&�j()"X�Rf�{�_��k�
�k�-빠u-�ZI#q8'��&U*}�y���w�Ł���]$��4+��}{� ���e�I��6�Z^��}�X���`����RIwsO�'U�-,���\rq�t�y)2Ր3��,��ݐ�6��)I�{����Hv���̦��}����z�Xε`5����lk�ddjݴ��Gq`��ٝUT��{� ��u���,�����C�	��!wn\��w^��5��x|�S}�ٚ���P�)#Q�8E"qh|�*}{�xv�, �}ۘUR��7�������#�ۘ�N=޻��T��޹�׼�~���%R�T�]�������z�C��z�j� ��죗�sN�V4�V�k�Fźa��Аj(�`X��iC�8p�=�)��8�[x��R+Wv���n�����lN�WU�/K[�r��-�1�e��sbb���\cEa*U�;q�ԯcX�&p,��]r(n�9�ݡ��\�mS�ײ)]TiXX���Q]�Zn=����
cr[�����w���{�;}>᢮�ې����d�,�/-4�P���f�JX���2���=�{�=��B��P�T�����Հ��VZ������X�܁�%˹.4�Ww.`���nl��X=sW��"#�s��G.��_;>��t1\�w }�}0�wRM��z��{� ��n�Em���F\w&ʩ%I>�� ~��������b�,��1�D��7ݹ�rJ���t�~ v�Lw۹�y*�X�I��q�q����L�Hc�7�V�UsҭV��ΧM���-��m�����*�^�o]��g�~���/࿵
Iq�R'�W}��b���V�
@
��DIVa�{ o��0�f���meܻ%����۹xﻋ <�v�I*������{� ���r;��q;�6�U�\Հ�i�Z��{��s�����7��o��w.Zq���0�٦�%׽���v, �}ۘ��]ܒn�	�T�S�8{7ey���&��g�8"K��w"V��µ�ID�72���s���7��, �}۟�IR�n�0˳��I�"�Bc�Ǡ_[��]sVݦXks~�9��"�z� �\,rL ���0�٦)B�"8Dr��y6��XwILP��%3R�ۗ.`uR�۹��{� 7����IRT����0yoc�ˊK$�K�Xks`{�]��X�?MX�L�?����ؿ��]L��p]����][u���!�z�\�F0#n��ԝ�{��4��,6B6�6���~��h׫�wJhu�@�g]���2'K'&����g$��wg=� �۳>��M��u7�]˻�-8��H`�8�5��x|�M��t�?v�C 7���W �<ML��`5�̀>�V=wE�y�Ȃb��qLA�ĪV�������"����Ԏ����0�$�v���ݜ`��0��_�����.Fyi+Z�WEN�^��[%3nM��j=�weAx���ב�S�ޝ�D�`���`7�� z�{����s��w� ���ڻ���nY�`��춬���7�ܗ�s܎r&OC�!6�ƛi����~Z�� �����>�@���[���M�LN- }n��w%��u�DDD'�����/퉴�"qı�94�����rڰ[��+��"9��PeB��7.�%ǭ��l5��2�֞Ƚ��(����[hf��mZ��嚝�61ŵ��M�3�6���Ѧvv��4�qZ�]�ط��NGmZZ"L��bd�G���a��	S�,���ݞ����[n7.��L��%���lѤ;iwd�iZwkYv6��Ef]A�O���Gf�D���r��i��\��6�;-�Q�kv�p�U���������G$��N��f�n�u�i휐P�2� ��D��wUU$�M�q����Ig�w_s�:�V�}n�޷Y��uBA���8�qh]�@�[��w��h��םJ���~��&؈�@2�<}�ŀ{�w,��I&���x��<ͱ�M����	����T�%�S��˱`?��+\���XwbSo���Q���z��@�mzz�h�V�}k��SI��$ks���,���v�s�5^.�pG�Дl��K߾�wf�MB���6ԑ8�_W�ߞ�޲�zչ�z��@���\���M캷[�I=���3� �|S�P��O�o��y��@�mz�u؛JDD��ղ���^,�ߺ�����z����OƁԷ�["q����E3C���*���;�s�� ���0n�Xys��#rE�,q4��9[^��Ī�IUv����;~���?o�L�}M9yW���I�v�亯k��^F47p�ܛ\c�X���#x:���ݵn����)�w�[��Jh��@���f���j�8"H`��x����g����߿=�e4
���o��q(ۖ��?o�L׻��J�T�^R��U�Є�	�4� �Z�Q]��/@a��z�o��'}��I>�{��%�q]ے;�p������׀o�?^��޲��׋dR7W�x��4�9*��R��wߙ�ߧ��9[^��:��HڒD�jLx��U���l��f� �vu0���QQ=�[75iI�8�47�]F��YM׻��IR��� �;�dr7"��r�"�?~٦|�5�u��ӌ��q�ʪ�9��5"$�$������� ��f�|��&��� �ޜ`��VcH���N=޲��]f�<���2O���v��(/�j��m�sY$����N�eܲ�1C	!�_u[��e4
�נ{�S@�9U�<$��nbnIL�pB�\��
<\c��Y㐢Ӑ=w#V���3�-�LԥT)Uz�Z���{��%��y��;M�c�ܸ����p�*�^��YM����=�)��331#���FȜn&
9�$��;�OƁ}�nh���*�^��wJ�I�H��j컆�J��w�� �ޜ`���*O�{8�7�����H�n�Fh���/;V��YM���@�������x1hE@.(��QU�d�������n��	`T�C�a��`&Fd��>���Jp<�R:�KGg���v�������7�O���.����Y���MMc�u!�k��bB@��HJ���>v+�B�$�����TW�#4�
`�'�V$@@ַ���{�� �M. Iz��4���cm\�{�#kd�a'-)crk�u�*n��$��T.0�('�ʔg.FM�J�=��;hȚ1��^�����vxݕ|�]+��Ā�C�Ɲ�Q'���q�;Lf��bx&VV����=2��s� ���)sSs��@*�mu<��i�zI��5��r�L�+�v���9F���y�y3�-4u�]���4��+nz�rjv.w:�;qnC��3̦e���47@Kɶ]m�cC�����MG�h����Z��EU�Vʁ�����]� )�6M�� �W5�;m��:鲺��+�+�����a˦Ͷ ���b�Wu��a�����Ud�0�p���npD����!�M(�C��M/y%��
���N^�7,rt�&��6�/k׬H���8ۇ ����k�Su���}i˼�Bq���x<��yS��f��Y�J�IH8"��������H��t�8��2�ʀ�R�L�����^Uz�Vw�8��=�l%��+�nwh�6�� pWV�yӷ+;�NtN{�NR�5uks��1�7<[�ف��@z��wNʪ�=�F6��VXF�/b�ul.t���izyRc���UT�i�X��K`0 ���Z�U���j����{hb�Wg[X����ٺ+Zm����IfX��@۶u���X��
JU�-��[��P�ճcT���*�r6�F+��(a ��4�1��C�����'�e���P��Rʝ�un��yA����[�k�B���G=��ٳ�[�=\���y��t�on��M�8�avv�U̹���qX];����f�"�]�mT�T�u'=r��I�m�Ƹ\ 6��7*�4���T�ɍQ���X��k�3�=r�I6��e�q�L���ć\�b[��M��f{3�=a9�#�נ^�c�u�+bQ�I�6IX�Zf�Wé�㊞b��Urb`�W��oA�M�{���z���A���~D�SjpR��~��h6,��W� �U�U,�i~T��#�w.\�]�]�S*��8���(�ڌt�m�zڐ�vM���3ۮ����g[�f4�nVG$��%���:%�u2�El�s�\[�V6����:hKmV��݊��M$��goi�z���N֭�r=�F���tgi���S�9[��,dM쀙K;	Z��ǩ�Dl��ۧv��5�װS�S��B��rne�a�av�uԗe�UB��UU$�o�<��w3�+�m�b뱷/bG�D8r���	�ᜢ�a��n,�	#�$I�p�j�=�4�7���|�J��a�|��Ͼh�[���!��z�h�V��;V����Ϊ�����k�N	ڰWI�_�s@����yڴz�h{���r&�ېv�����gm�<��`}J��w�� �7��B��.ܔ�*�`=�Ձ����~W{-��߿��~��ɿ�ԷC&��K�ѐ6�5�%&�!��6.�t��#b�rV{����I����x�Ɏ	��-�O�_u[��f�R�K�����vs�n�r\�����nd��=��)ʪ�T���3��~��^���3�J�7�����$Q&♠w~���h���/�����VI�BG?��$�4�ՠ~��L{�U$��������Lk ���=�)�_u[��e0}ݘԩu��RZ���rⶣR�M;s�2lnVw5׵��ݷ ]�n���:�ګ��"�2T���`�D����<X��S@/[4���*�`�X�ę"�jf��Қz٠w���}�no$�;M�c���ܑܻ� v�L$�Ϸ�ɞ+�|R��4B��B�*�HD�n����>�d��>��"q���� ӓC����`��ŀ~�f��%�w�}��;/��M�ऍ��#��_u[��O{�vbr%�bX���ىȖ%�b}�{��,K���};��M��G��<.��e�;����É�(:�Э�5m\P�������\̕�@�w����,K������bX�'~�vbr%�bX�{����(O"j%�b~�����I��I�����18G(�㻸br%�bX���ى�~#���bw�߸br%�bX������,K�^��Kª�I��K��s	i�q��s�,K�����'"X�%��~��Ȗ?�Xj&�}���br%�bX���?LND�,KϷ�������Ԇ�M�f'"X�%��~��Ȗ%�b{�s��,K�����ND�,����� LP�&��=2��&Re&R��оm\�������9ı,O{�vbr%�bX���ىȖ%�b}�{��,K��v�e/
L��L���k���ܑܐ��bb�9�v��ԭtI���[)`6kn-㨌\7nz�y��M��)6�����{��7����f'"X�%���ND�,K����yı,O}�vbr%�bYK��ּ�.K��9j+���&Re'�{���bX�'}���'"X�%����ND�,K�o�����"Ue+)2���?��A�$���eȲ�"X�%�����19ı,O}�vbr%����j'����Ȗ%�bn���)xRe&Re-�x]�仑H����ND�,K�w��ND�,K�o����bX�'���19İ?A5߻y�br%�bX������.ۗEq�p�^�I��K��甼)X�%�������D�,K߻s���Kı=�}���Kı8���HIQHB!o~��'v\��� �Y�v�V�R^?���˾��^�(�eJՓn�0nݎ��SBQJ���]*F��8M���ۍ�v���e�[����ȍ`���&ĖĤ��s�':�n�\e�{V������:�w��Jd^9`�b�*=��=����������綶�:�e�v�;%��W��2�(y&�!Ȋ�mv�����\��ŧ\�&���t/R:�8�ٚv:%<��@'3���`���A��[�ۗ\��i��������\~�ғ)2�)}�xbr%�bX�{���ND�,K�w��U9ı,O>�{q9ı,O=�t�r��"%Ŕ�)2�)2��~�ىȖ%�b{��ۉȖ%�by��ۉȖ%�b{�s��?��������ڹw%��7p�^�I�X�}�߮'"X�%����n'"X�bX������Kı<�띘��b2�){�{�8��+��m��&R�,O>�{q9ı,O}�vbr%�bX�{���ND�,T,O}�{q9��I�������r\v����Kı=��ىȖ%�by��;19ı,O}�vbr%�bX�}�����L��_%��0�v\��_m��3��I��3�z��Z��U/iI�rˎ8��]��_�L��L���Ϧ'"X�%����ND�,Kϻ��"r%�bX������Kı;�9x;.\�"��n;�R��L��^�����8�` � �����|��K}�=���bX�'�}����bX�'��s��,K���P�-��(�7.K)2�)~���9ı,O}�vbr%�%�by��;19ı,O}�{q9ı,O=]̿����� �<��I��I����ىȖ%�by��;19ı,O}�{q9ı,O>�{q9ı,O��:T��.ƤD��^�I��K�~�ىȖ%�`�{��ۉȖ%�by��ۉȖ%�b{�s��,K7������?ep�L��m�h��Ԩ��)���q�&�55.t�ΧOS�l��sw��]�nbr%�bX�����r%�bX�}���r%�bX������Kı<�띘��bX�'�>�,�7�����v܏)xRe&Re/�;�R𪥱,K�{����bX�'��s��,K������,K����\�{���-E �<��I��I������Ȗ%�by��;19��6�F�m�<C��8�x{�����ND�,K�w;19ı,O>�-�H�%��K.ᔼ)2���)~�oy�Ȗ%�b{��ۉȖ%�by�s��,K����f'"X�%������ܗw	v�)xRe&Re/}�ۉȖ%�by�s��,K����f'"X�%��^��,K����~�M�!3
�X6o]��E)z�%���a����F�=7T��n���{���w}F�Cf�m��'�,K�������Kı=��ىȖ%�by�׼��Kı<�{�br%�bX�zw�k��d�ڂp��2��&Re&R���)x!$$�<��ݦA$���X��H�{�)aK���Ε��Kzq�P���e7�o{���bX�'�v��'"X�%�����,K����f'"X�#)n�q��)2�)2�_�ͩ"��&�Kw�ND�,��T5����X��bX�'����'"X�%���gf'"X�D����������^�I��K�[�1�$n)qܹ7���,K����f'"X�%���gf'"X�%��\���Kı_���)xRe&Re-�����W.).Z�i�m7h��gY1��Wk�[�VB�Y������g�h�rG]Ym������X�'�}����bX�'��s��,K��]�u�Ȗ%�by�s��,S)2����]�r�Y�e�2��&%�by��;19ı,O5��X��bX�'�w;19ı,O��;19�Re&R�㗃�ܗr),�ᔼı,O5��X��bX�'�w;19ı,O��;19ı,O=��f'
L��L�׻b��pR��"X�%�����ND�,K���ND�,K�~�ىȖ%�����R��L��_�]̿���W\ىȖ%�b}��ىȖ%�by��;19ı,O5��X��bX�'�w�YK)2�)=��)�7q˸�y۝I�ڞ��s�kD*��{#嬠7h1�Z���k��v��d󛦮r����a�Ϋ��&cMÉ�&֌e����l㋡ێv�o;�Ng\.:E�r����恶���{2ὐ�r�˿��}��IF�DTݻ)2��2���p��̅�;X:�<��f�b6��3��"S��㳺���G�2Z��o{�������=��;t�~.\�1kcq]8�q���%^�[�v�u@:�2�	���B�4]�H�!���&Re&R����19ı,O5��X��bX�'�w�0?�@"j%�bw����,��L���+]�$%�-�2��'ı/��w�Ȗ%�by�{��,K��ﳳ�,K��߮vbr#)2�){�w�8����h�&R�bX�'�w�19ı,O��;19��]D�O~����,Kľ���)xRe&Re/w�ߗ%�.H�Q]�of'"X�%���gf'"X�%��\���Kı<�{�br%�bX���Ŕ�)2�)2���7�Kd��ȯz���'"X�%��\���Kİ�*1@=��ߵ��Kı=���19ı,O��;19ı,O>;�E���0f]u��ݵn�1�D]��r��\fW�VR���y/<����fJ�4�m��D�,K�w��'"X�%����ND�,K���ND�,K�~�ٔ�)2�)2�^���]�QHK��Kı<����Pڤ��>H�`��1��}臨q@��X�ı5�sɉȖ%�by�nvbr%�bX������O�����'������FHӄ.E��)2�)2����br%�bX�{���ND��0�MD����x��bX�'����'"X�Re/oӭqqY�ݵ"$�R��N"���\���Kı/��w�Ȗ%�by�{��,K��ﳳ�I��K��E��$���H��Kı/��w�Ȗ%�by�{��,K��ﳳ�,K��߮vbr{��7������xR�W0&�71����KS���i�4ۧGr���%j!�{����_8����@��w�{��7������Ȗ%�b{߳��,K��߮vbr%�bX�{���r%�bX��u�.K.\����.E��)2�)2���;19ı,O=��f'"X�%����n'"X�%����N@D�,S)wv��q\v��p�^�I�by��;19ı,O��{q9�!���D~��|P�I��yX�����4h,RMs��682��&�Md�!4KE�Þ&�DH1 �4E�h��AP�]!�]����7��<cZ<�C��M���, S���8)v�H$7NmB�CB�]k@)��BΧ��'��%}WR�H�-t��	��ܡ,���jB48����0�8L�YXT$gG��|��f��a���󆷌�l�OT�����]��*? �ҨEDb	�'�@O@|�����)�D��bdO�����Kı>��ي��L��]�r�w.[�H�,��Ȗ%�bw����,K�����'"X�%�߾��ND�,AlO=��K)2�)nͱ>���Э\�w��Ȗ%�by�s��,K���gf'"X�%��\���Kı;��yK)2�)}T�w�חn����H�B�U8��U�k�wK}���� 1�Y�7\Z�r�#.![aƈB�R�Re&R�?w��br%�bX�{���ND�,K�ｸ��'�5ı=���18Re&Re/��n�뉑�ݻ�$�R�%�bX��~��'!�R:���'�����Kı=���19ı,N��q��)2�)2�_���ڒA�b$���x��bX�'}�{q9ı,O>�vbr%�6%�߾��ND�,K��_L��I��I���;��q��5m��'"X�~EX��s���Kı?w��br%�bX��~��'"X��Л��衱D:{�S��/��>yK)2�)~�ߒK%܅���ַ19ı,N��vbr%�bX~X������<�bX�'�����Kı<��ىȖ%�b{���]޵����!+gػ+ �`v�b
�v�7>8�&W\�]m�jxn!'\���r%�bX��~��'"X�%��w��ND�,Kϻ����bX�'~�;1^�I��K��^7n����L���br%�bX��}���ı,N�����Kı;��ىȖ%�bw߻�LND�*���'{����o[���oV�w�,K�����br%�bX������K��Q5����LND�,K�����r%�bX���l�j�"��]�)xRe&$�K�s���I�bX����S�,K���n'"X�%�߻����bX�'u߭��l�:.� I��I��I����,�^�K���g��Ȗ%�b~���19ı,N��vbr%�bX���� FAL�`P�m����H$� �NIw��[.�`\�T!� �V6
��.�q�6�=dc��� �q	{v����&ܼ�c�Q�������.�zV5�'0��a�
��������i�'i)u�l�i]�ڊ۪;$zx^.s�s�'k�;F^8ɩ�	eNs��S���-l�΢4Q�6%��>���b6�N8��:�3\K���ϖ��yv��[f��=��sw.�w/)~�T��%�����2�W#n�Tu�+k���z[��v:��wIiL��J�6�Q;65]������7���{�O����Ȗ%�bw��f'"X�%�߾��G�,K��w����bYI��u��9B�)n[nG��)2������ND�,K�}����bX�'}�����Kı;��ۉȖ%)2��w��$�]�\�$YK)X�'~�;19ı,N��y��ȖbX��}���Kı;�{��,��L����-;�]��Enᔼ)8� j'���LND�,K�����r%�bX����Ȗ%�bwﳳ)xRe&Re.�9xݻ�#�8�ܗ19ı,N����r%�bX=���Ȗ%�bwﳳ�,K��v����&Re&R�7���i�q�q�cѫ��;uڄ�TC�T��Z���5��D��Erۑ�/
L��L������Kı;��ىȖ%�bw߻x`~'�5ı?}�߮'"X�Re/�}�/�+l"��\�)xRe'���gf'!�P3z
�dND�5�ݼ19ı,N���q9ı,N�����Kı;��n��v�������19ı,N��oND�,K�ｸ��c�AXj&�~���19ı,O��~���bX�'u�žvIwb��v��^�I�U$�W������Kı?w����bX�'u���'"X�%��~��Ȗ%��[����!w�-�#�^�I��N�����Kı;���9ı,N��oND�,K�ｸ��bX���������MCt���]�۰�r�n����Wn�ז��ȹ۾���I�Q]�"�^�I��K�w�)xR�,K�����,K���n�FyQ,K�~�Ȗ%�b~���K�\R;�dN�^R��L��]����~Qc���b~��\ND�,K�~�Ȗ%�b_{�w�ȟ����)}������\�q����^�K������r%�bX����Ȗ8~")�B���<�w��7�Ȗ%�b~��oND�,K��;�o[HЭ\��yK)3�����ߖR�Kı/߻�x��bX�'}���'"X�%����n'"X�%��N��x�[��-HB�YK)2�)?{zbr%�bX=�����bX�'�ｸ��bX�'~�xbr%�bX��N�����:ml�r�rtԳ�8-p܇��A�u�B.On�ˍ��Wf}1�<�[ޥ����%�bX������,K������,K����ND�,FR~���^�I��K���X�qv-ٽ˫��,K�������$D�K�~�Ȗ%�b_�w��9ı,N��oND�,K�}{�K��A܅��r<��I��I��{�YK�bX������Kı;�ݼ19ı,O��{q9ı,O~o[�$r��R��L�%E+)o����,K���^��bX�'�ｸ��bX
b �Ң0CL�+�n��T��#�"�iD��y��8br%��I������vˊ�,�;�R��X�'}���'"X�%��:�߿oȖ%�b~���19ı,O{�vbp��L��\���.�-B9$vvq96�e��Ȉ֊���<�F��_�}�Crƺ�˃��L��qyK�I��I��o߷�Ȗ%�bw���'"X�%��~��ND�,K�����,K���βK�W�&R��L��]����bX�'��;19ı,N��oND�,K��{�ND�,K���_�E����$�)xRe&Re/{�vbr%�bX������c� j&�^����9ı,O�����b2�)u��`��dt�\��K)X�'~���'"X�%�~���'"X�%�߾�ND�,K������b�I���x�2\C�j2Aۋ)xRbX�'��;19ı,?�{��Ȗ%�b}���br%�bX�����
L��L�~}���T#@ߏ��3`M%��i'��h6u��p^��rQ�jH^n��[l��\nt[���0Zc
5+�qPR�);��A���{)��u��sq��=��8�n������8��u�
zys��{��p��qd�Q�����dV��f��ͧ>3�] �Z�R�FN��ڹ�qʻhM�Is�ч��T�h�-�r��m۳fl���z-68�8����}�����֢%�5�Z��8���X'vp�jc.�Q�f��T/ �+�a��	���{��%���8br%�bX������Kı;�ݼ0?�)<���%�߿g�)xRe&Re/t;���۹#�Wd�19ı,O{�vbr-�bX������bX�'��;19ı,N��x���&Re&R���ڎKr�]��e��'"X�%�߾��Ȗ%�b}�s��,K��w�'"X�%��nq��)2�)2�{�G�9pw७]ݘ��bX�'��;19ı,N��xbr%�bX������Kı;���)xRe&Re-��b� �0-^�w��ND�,K�����bX�'��;19ı,N�����bX�R�{8�^�I��K�[�-�ar)��_Eu>�ڱ��H�Z�5m��ʣx��u�0f�yLݻ%j���w�����oq�������bX�'{�wW�,K����f'"X�%��~�ND�,JR��n�u���ڹ$2��&Re'��;���D<|�6�L�b}�����bX�'�����bX�'��;2��/�%n���K���%���ڌ�]�W�,K��߿s�,K��w�'"X�b{߳��,K����yK)2�)v��,r"A�L�n��ND�,�@�O�w��'"X�%�����Ȗ%�bw�guq9ı)K}��)xRe&Re/ކ�����.Ib٭n�f'"X�%��~��ND�,K��;��Ȗ%�b}�{�ND�,K�����bX�'�|~������{�;'t����Gg^���ڞu��kb�2�t7
%���}���ZHӆ�{���2X�'���ڸ��bX�'�����Kı;���� �$��~�� ����'-㻱KV�[�H ����i�;ı;���Ȗ%�b{߳��,K��~���r-�bX�w}���Z�nI��)2�)2�{��Ȗ%�b{߳��,ttT��!�O�"r&w��'"X�%�������bX�'};�5�nI.
B�e/
L��L��nq�Ȗ%�bw�guq9ı,O��vbr%�`~@�������K�e/��n�}q24�W-C)xRe&Qbw�guq9ı,?�߹�byı,O�w�ND�,K������c���{~~��LR�U��k�hl)�M+��'J[uԮ&�Mc4�ѧ��.t�;��$��&Re&R�{8�^X�%��~�ND�,K������bX�'{�wW�,K���^�R�jKe�Y-�p�^�I��K���e/�,K������bX�'{�wW�,K����f'"~U5���;��v��˒�Q]�"�^�I��K~��br%�bX����\ND�,K�{����bX�'}��19ı,N��õˎ�Kq��p�^�I��K�s����bX�'��;19ı,N��vbr%�`~P��� 1$D|G���"k��y19ıK�ﺏ,n�pmBZ�r�R��L�����f'"X�%��~�ND�,K������bX�'{�wW�,K=��~~~o�uRݐ��+��V��^�A�Ku��ȹ��5��m��`
�<,+���v��F���nbr%�bX������Kı=��ىȖ%�bw�guq9ı,O��vbr%�bX���l�MW.8'�E��)2�)2����R��X�'{�wW�,K����f'"X�%��~�ND�,K���jC��di�.Z$�R��L��]۝o)x%�bX�{����Kı<�����Kı=��ىȖ%�by��v�ԗwb��r[�^�I��K}��)yı,O=�;19ı,O{�vbr%�bX�w��'"X�%��~�楑Il�%�.K)2�)~�o<�Ȗ%�b{߳��,K��guq9ı,O��vbr%�bX��l�CPa�6B1]��������h�@TP^��)����V0,Q�i���B���!s�)�f!�Ui@j��$	l�u4h
j�k~<	s�I�l��B-��C^D�@"@�"R�B<Bkg�O� ��"F2.����
��4M:b�֤HBB�D�!X�	�%�
at��>��(U ��P�~T�t�$	ZQR+ė�|ߍ߲H�,��MS`m)'�Vצ�ՑNq�����cf`�y.N$�ƭ��}�C
&�G�5e��e�'e�!3�) �X&�$��J������[�y�|[q��]�2Y���
Ajs.T�ur@�%31��cK�;*�����fy��	��e��m��[�U���v�V�5K��f���%���u�������[ΰmN��Ψ����v[�\
ޤ-�m����,vxck�'v�nq�i�j7n��6kj��SV��JpS]`k<�B9�$�\��� �2�˳ ��tJq�Pr@��vZ��kh���u�j$A��a��T����UjU�YX�k �l6�Em��hV9�k�YݗSl�Ya&���\��:��]����e4t���m�Kj��X�tz�:6A:�nI���3��zx����=�v�;�}�u:6�Hs����:���j=�9����&+�NVPMƜ��Ċ�.*��ʮ��m{m�r�Z���u�dh�ce��dР3��6�j��J	�k�ʱ�,f�� � K'�m;rN��]s���O�=`��go<:�k�Cm�;.����q��2��n��L�;:�����=z�z�<��ľ�uI-�\�LIc�=�.v#f�"��]n!��Ў5vJ:�V��U������Zt�<�`H��t�n�b�(g�B��8��6M	���I�9�{Zj�Tɔ�.��-΋jN&��XZ+�`+�����-�+�[IX禲�l�����5�d)_��'�n��%s�qŜ��Q=Q�`��<�����&V�s	���m�j�Ƀ���/R�^[��&ƽ��֧qW4��Yw[���X��iɳ��uj@�U�,Hp��;�m�[p�\ U�M2��]��f����x�Y�꛶�J�a۬�Η*|�|*�����%��F��Wn��:����s/�mE�&�t;n\�ӭ�I��@��#����{8-67m�9�l�ݵ����ޮ����u��	��P�C�0�")] ���A*��O OP�����UU��+J�Լ�O#�#�ӈ����y�&�q����+���S�e�t�]D�Q�c�౮��B�fy�OU�8�6;	t���X2�P"�6����jmV��s����5��Xm��_0!�Gume�wn����#��gV��[�F�۰>&�]�(R�J����U�4�n�ii2*룎ۅ%�W���j�]����Ұ��s%��nD����%�"��y�%�2�������}���UuR�#��N6����QNg8�p�]�[��q�[y�IѰ�ۻ�.K�Epw�/�L��L��ۜbr%�bX�w��'"X�%�����ND�,K�~��ND�,K��t],��F�6�����{��7���������bX�'��;19ı,O=�;19ı,O{�vbr'�5SQ,OV��?jK��d�n弥�I��I�w���br%�bX�{�vbr%��T���~�~���bX�'����q9�L��[Ӻ�$A%��)-ˆR�Kı<�����Kı=��ىȖ%�by߳����bX�'��;18Re&Re.�w1߈Dn�88B�K�,K���gf'"X�%��P����ڸ�D�,K�~���,K����K)2�){z��m�;Mܴ���cu8t���9ѷ4ĳ�� ��Q�bs3ͩ��S[t�h�^�o����7���'��;��Ȗ%�b}�s��,K��߳��,K���gf'"X�#)~���+%�]أ$��&Re'��;19�0%T���2%��w919ı,O{����Kı<���\ND��j��X�~��,r)-� �]�p�^�I��K��~���bX�'��;19ı,O;�wW�,K����f'"X�%�硽~;wr��v(�p�^�I��K������bX�'��;��Ȗ%�b}�s��,K�Q=���19Ĳ�)}���%ܸ��,w��I��K������Kı>��ىȖ%�by��ىȖ%�b{߳��,FRe.�v	��q�7i��˪c]��`���K�iy`D������y��齋��p��p�r�R��L��[�gK�bX�{�vbr%�bX������FRe&R�۝o)xRe&Re-��[RDH�A���)xRe&Re/��甼��Q5���s���Kı=�����Ȗ%�b}�s��?���'c���pp��2��&Re&R߻��'"X�%��~���r%�4�~J�P���DZ���7�D�'��?LND�,K���n'"X�%�|���&F�� �$2��&Re&R�۝���Kı>��ىȖ%�by�����Kı=��ىȖ%�by����%�]����&Re&R�{����bX����g\O"X�%�����Ȗ%�by߳����bX�������n��t���Z��ô˧�c����5�WO+֤knס+���gB�{���]�s�,Kľ{�w�Ȗ%�b{߳��,K��guq9�e&R�{8�^�I��K���~;wr��z�6jn�{��Kı<��ى�~Q��j%�����\ND�,Kﻟ�'"X�%�|����,K��{��ԗr㻒�d-�2��&Re&R�۝o�,K��߳��,Kľ{�w�Ȗ%�by�s��,K������R\-�-ܷ��)2�>J����{ό��I��I��������*�&R2�uJ�����ͷ�o��ԑ7L���{��>���>�+Z�Қ֠�����8�r�DH�9R�ŷ5�.�Js�]a�aZk�6�oF��UɄ��޲�ץk@��S@>�Y�r(es�C� ��4�J���s����ŀw_��κe���:�IqvA�%���f���va�IR�M��������M��;��+���{��>���>�+Z�Қ��k�9��Ȝ�޲��ٶ�߽�`��ـu�EUI-�n����u���-��v��r7��l�g��	�����t1.�N��T`3E,2�W��K.�ș�D�	�Y�ջS�Qg=��Mny�Z6���`���QJl
�s�ߍ�_tQ�Z۫�k�N�8�l�6�2�7mѩ��v�=@l�����Ӹ-�z1��d��dܝ���U�ĸs�N��K*�N�n+�n|���"��������x������ m)4Kss���Gk�m��W�U�G#a:��Euu�g�а�a��F�N���k@��S@��)�}�)�}���k�p��Ӎh�Jh{�4�e4�J���#���k��J`L���{��hz�h^����M�-B{�Ań�4�e,{NU���2�܎.�֏zg�'�AAHh^����M�t�������\R�Rb�9�rF����"w-�eR��1���m�`9�u�a�^�k����G0m�JAHց�t����S@��S@���h�u�Ib��Q�@��2��r#���']Y`ov����M��V�H�Q�?��@��S@Ǵ�Y�q-�^,�n��*i51��Dp�>�+Z�Қ��M�YM��_�X��1A��;ݦXݦX�L�1�9V�Z"~q�')h�:6:vu���;u�9;TJl <�\2��Z4:cR�9�(.��I����2�κe��i��r"#n��w���x����]� ���0{NU���2���2�7�0�5�D)R�pr���x���0�%�/iQK�]���SH>����w��'��L��[H�G0m�JAHց�t���t� ���0:��?����彌w$��Hc���}�)�}�)�}l�h�JhZ
�8ҎH���L���`#ú�&�ˢ��u��;�od�ױ�CY���؃���N޲���ց�t��{vq�wt�vK��W%��[�`n͕~�BF�[�u�,����J5&I�Piƴ{�4��4�e4�����Q�G�L���Ԫ���� ��N07w,�� AIH�a�E�X1F"�U���.��P` l	�yɒO�>���"QH�A��}�)�}m�h�Jh{�4ٙ�������x�6M��07k��;��<��Q�ӈ���문�abI��)r�j8���~�� ��S@��)�}�)�|�R1�qb�$�4{�4�Қ޲�׮�@�:��6�!�6����t��������Y�{�)�}��]�9�0Ɏ�@��S@���h�Jh{�4l��8��$n"8h^�%���2���2�κe��|�Ⱦv BuJ�U ���G����]��߷3�ۨ^q-��P)���O7bE��	63�iCu���eͻ*�:F��-�/I��@�j�;i�Þ�Ƣ���2�-����Ɩ��=��dꮮ���'�3׌��-���;:۶��v-���2�2-Z�69�	��#B]m���%m�������_5��6�u�HS��l�;[L�^��4d���X3�Ei��u�"�
��$��kz�ֵf�ڴ���b�^��.^�Y��3��3usW&j�����6�(�7$����v䳀�ޜ`o���}�)�u��=Ϩ���ܘ��׮�����׮�@��S@��ROp�6�A�&hz�h�ܖ{���� ޤ����7!��=��,�=�g�����X�߷�U��#��Q�9��e��]Ł�t��wE�Q��Hv��d���4���h�3U�C�;k��r�C�lt�S�0�;���`n�������ڒ���i`dwRy#�[�+Q\�E�y�f�t�K�UB��>s"9�%��wi�=wn�����I��N�v�Қ׮�������Ʊ%#��D�jHh�Jh^��޲��v��$NL�G��s@��S@���@��S@���)�$�"�e����9�=������i����-�\a�9x)M���9�7Y �4�e4z�4{�4�]� �%C+��	�y���-��=��>�w4�e4W�����FD�4{�4��{�>��3A}P�xF�U$4.�!m6�;jF�o�NF�!(�,�J�2+
|{+���@�sÐ�,t�yY������zg61�
j1!B����Dc�!��6��Xſ p_F���!�J@�($�L��:H�.�.��Q����RA�G���Z��8���d"쁴3NO��M	�tD��F�.�&��>}<�i �g({�a�(d8B��5�R���X<S�*h��$�����<�7[!�4m-�i�!�bc��jy�z;��%JM|1�BM'=��< �{��OjPC��=Q4qD�B*��mT04�8�� �@�!Qr$ 2��WJ:Co�hP�)肼�>��$�y�ٹ�����r��+�n\0:�U?ݽ��?{ӌw��`uRUI�����3�D�o$��c�I�޲��v�Қ׮�}�Ef<ncd��M1��u:�^-�ϵ<�8�r�-��ҌQ��(����q52H�Dp�-��=��>�wU$�a�ޜ`�ޣ-�ܒ\Q�ڒ�Қ׮�����o]��J�=��wd�w��\0�݋ ��S@�݆��t��}��=�	#�H9��YM�v�Қ�pN���B���tw 6@@�jR#A��FR�]
K��$%�@ m=Xr���$��~�()1�j
C@�݆��t����s@��S@>[N���qH廮�Ů�L>��ݜ��N�]3kWG4i�x�j'0M�Q�9��M�e4�e4m�hN��n	�d�UM6�,�X�tX��/ܪ���{��ݹj�-E$��ޜ`۰�=��>�w4l��H��#n"8h��h�Jh�������s���%$�dJ6������`=t�;������9��ß{�?�������-�&B�40u<Di�n�5Oaj�N�p[m��%�:��x� � �p<���M-��^��c{F��$�nqC̝��$^�m��	Q�c��қa�����۰)�x���vv��q����{;�Й1��酑ӭ��n���l�Ҿ6ύ�[q��r�� ٍ���6�UHɺ'sʆ�m{F3�/[n@`^���{��������d��	�p�v惮�=�º��lte�~k�:l���Y+ V��f�J˖��8~���?��M��a�}��/��'�dRLq�d����S@Ǯ�3�L��e�>���
Ly���>�v��M�����h�&�sM�Q�9�t��z�h��4�]��ו�8�q&�1������h^��t���㕐����6��&��mWc^�$\�<.Q����sn�F݅s=)I�	���(�L�n�����a�}��/YM��6Is$m�D��$��߳s8x�����TCS&�&��)�{��.u���%�L�F9!�}��;���}�@���4s�(ۍ���䄎s�h��4�n�@��)�w��b{�I��'�}�@���4�Қs�h��aF�b��Ǌ9n�#`q����6�!}U�`�A��β�V�F�Bۦ�PR0�8�����a�}��;��@>�Y�T{��0I���C@��2�ݖՀguՁ�n�5�w#�n%1�8�wYM ��f�?�� �T��$����9ȎG9�]��X�^,���(��Q�&F7 ��f��e4�Қu��:ثnH��#n"!94WL�=�;�7��`�u`f�U.���b�c���mS��;a��u`Wk��]3�u1[(�]l�ݱsĕ\���@�����e4��h�S@�}D��N$$p�;���w����h^��;�j1=�	$�)&h{��=l����M��� ���W2	1�i���/YM�ҙ$�߾�$�8���B#��s��q��{u`u�"h��)������>�)�^�s@;�f�z�h��~>�m���4Q��JLsm������;��݄�f���X&��8�^�s@;�f�z�h^��>�T]�cq
6d��&h{��/;V���M���[m�smFF;� �ou�o�L:�7�݋ 7��\��b��LiD)���M�����4�ՠz��&�H����	4��h{��/;V���4�?R�I*�f��r��n]
Yl�ݕ�ݭA\��Ў�VY'�7X�8+tm�\۶�n^�e�A��܀�K;\�����L���@;%̽�v��tI��ϒC�Ӷʣ��<�
tr��'�=��O��9��G�g�硏�1�s�jx	6�H��%����Ƽ��P�����lc��\�]mh�4�򺃲'����26�d��ѶcdX�N�訡�Qp0T+nY2���?��эv���-�Q����э�W����s��u{s4�zp�^4�~2I�7V�mX��`=n���#sY��������j�>�Jh�����h�!���27	"�=��/[��z٠^v��.��1�Gq�4�S@>�f�yڴ�Jhg���x��21�h׬�/;V���M���=��i	�kV}�e#��8�a�-&��v� =�.�خnӭ�l=[-Ҥh��XݦX]3�G9����<M9n䉷.���e��RD"�n"@`���Pd	4id"�@%E�$	Ay���3]Y`���z���!L�7�E4�S@>��@�e4{�4첳��IŒcn���u��=��=l���c���1�&8�nM��h��=z�h޶h�b��������N����x�h�oi���v�1��n�sV���,!����H��4{�4^�����z�h��X���GQ����q`���޺e���2���K%��d��L�ܙ�z٠wYM>�6����O�OQ^s���2I��h�D�@NdM��4�wYM��M����YM���[�jI1�4{�4[w4�e4}٦Ԗ��~+n�q]�Q�m���N�i.������L�f���R���l�nwi���!��� ���`~٦�YM��M�,��'�D�d�ܙ`g]2��t���e���Ł�ѕ�c�Lq&A8h�S@��S@��s@��S@�u(��N89�J�����݋ ���0.�H��R
�Q<��}��ɀz�=c�ڍGQ�@��s@��S@�Қ֙F�֤��P�q�����`y��d��E�{X䝧7�� �Y���K$��d��L�ܙ�}�)�n�e���3܌A���,�c�
j)ݸ�[�`��L�l�ݜ`�v,��4�T�lս�X8\�շ.u������YM��h���)�9�z۹�}�)�����M�,���ȲF�I�ɖu�,	�#�߽]\��3{��@U�Ѐ���@U��� *��b 
� Uʀ�� W�� ��H�Q	E�DX#P� �DX"A`�BDX�A`�E�!E�,*�DX�DT"�E�(DXE��DX�E�� Q(� � ,Q*�1DX�Ab$Q$1BE�EdA`E`@	E�DYAdQ�P�DXAdAP�UA� *�� ��� W� 
� Ux� *��@U�J 
��P Uʀ��� _�@U�@U��PVI��U~dA
���@�����l���G� ���kA�@Ӷ 8�-D�j�@�kJvvĺ�B�
t�7�   B�lJ
� �3JZhR �U ��A$�h��٤*Rl�B�z�AAB����P
*��>����o�Z2n�[�=�*���ݝ=�u�o<m���ݍϥ �>���9�x��=��næ��>�5�Sʝ7a�#W������ 

���|{<��CN��y�*�o����!��<�B\o�Á��������^�I��>}��u�`>�ބ���a�F�-������@ B������o!�cҶ��/pp7`6ǾϞ������^���p�L��4�`{�R�l��v9M�G���:[={�v�XV�)��
@I@ѽ��(�E��n��݇a��wB�{�:n���������;��9:�x<	<���w���݃l�wc�{} ����Р�uZ�m���twc�����p�� ���r >� ��J�� [� �9�� �B� Z��� ��t�l �>�94hwo{��   Z   �($�i�I�)L��@     ����R�$�P�  @  ��U*$jz��h      ��U�T`       )) $F�
=M1Fj4z��&=(i��5<�A$�"4��   4 �����uϾ}ߎz�y�׳�����(�w9��R)Њ�}"H�ܟɊ���������ݏ����*�ܑ�1���8:�"�������h$Si�_?�|gן_ÿ�߷��~_��ffv��˻��m����������������S�����u�����������{ۻ��������[������:4n�o��+-��v�nfn���������������r���ݻ����bŋ�ř���s��}���nl�In�����a�����)KwwwwwwwwwF�UUi�������� � @�fW�P�ď9C�D�r���%�>4'ƣ�P�Ɗ|j��"|d���U>2��U_"�ʧlI�v�'mA|j��T>4����^�ޒ{�x_U�J�1'�x�/�+�*|e=eS���s
��^�G���5U=�8��<eu��+ƈ�`��R��GƥZD�ңޢ�0�_mTsA|j����|ju�+����|eQ��U�>��s��!����	p�$���~��~�4�=��*��Sr��%5$��)s"�I�&��>s@{�!{�J�Ԛ��c�N�3���r��{:��i���]W�Ι�Z��n��~��2A�Jͺ�j�,(�	ǨPh��b��<Suu(H>4��-ˢD��J�	��h�����R��U�@�)��;�Cu�<xZ~#�S�2P�`�YH2��d7��j?ʃ��e�mN�2�f�$F�PzU��A�oZ��Ϥd/Z�
<	&X[�A��NZLPc�2�tt�+'7|L��IW���p�gU�V�q�*���
�CaQɜcng:2�cg4�3
�Qi(a��T�����J	R��Y~�O(��N1R�nmn��$V�SE�v�UӦ�I<{D��h׹��f���b�R�#D�� B�AQ&owW����
�J��p߃�5	Ov�aW���OyWR�^�_V��$.Qa�鱷,��8nf��6qgDBHHF��Iɓ|jS���G��;��{��;R4`\%Yɰ��f͑��m�ǩ������P�A*5��֤�(�5XH$#`d8�ٸ�n,Y���qu��0�0b�2���`jklH�bB�5P�%gVf�Zh5�^%D���,��B��I�Y���ku�WeM����΄t���
-�@/bk�*guƃ�c%(��$C��D�N�t�N�\�t!;�)���HO��3q2����p(����F(�m�W,��8�#f��	M�����$FB]��&�%��6��\#$���9c�����z��e�<h��U��c����a��j�{�(��k�@��Dh%P�`F�Wf��\��	0�	Ҙ�e�ɭ���)%F�浲5{sr�5�t�`�2�2��eoU\��aN��]!�kF_2w��S��������㐨�U�Q
��1�NY�%,����߯a(�Qa(%m�7*�
��t1�@l�%[�H$�j$aJٚ�+5��Y}=�Ua�N�	a-L6�W��ŧ�z�1rҺN6��s��\ͳ�F�MfM�͙V���$,Q͚#E7mݘB��E�0Ҟcp#�8l6I�#�e:�AӉ������7efw�np���F8�0ָ�0̳5����3��՗5��- �8L�D`�~�)5@^�Șwֹ�
d`���Z�7]�󺰠�E]��U�ǽt�`Ť��xX����IF�>�^�tj�ayy��i�4��;�U�w�*t�oFRB;IE�"Z����HFh�g',,�k0��U�1�8�$��}k$�]� J�>�3Wo$] fإH6*�3a�"SUz���_eVh�\�;҃��( S���5!��h�����֎�t�X2��I���?K��'��$��]٥JE*��V��byfk@[�W�X�|�Z��հ�cD���
ɴ�ΰh�#E�h�Jj$]�h4��Κ�m���KRB��"H4[�7�&�Ѥ�T$�e�kVڵh운�4O�LXzc �Ȱ"$c��VQe_�r��	0��7�w9�q�@�00��thcH\��Z��%�v���IE�^�GB�.�����ڳa�M����&�7zw7�f�exʼ�QF�e*>>W�e;�h�7�~->�.�~`�~W���2��"Ϥϱ�� #USwsF�9����d����r�ŏA���T0Pd)j�L���zda9G"�2���������L�y�p^Uz�Z��+�� ��12�<��M�6���N�#���4`�6l�rHM;�08FHH�i����H�|���n�	�V=:����Jlt�Hi Q{!¡mT�D/%O"uU���^ˑ��`�>b�ǀ�r	U�;��D7�2��������R	˽Ֆi�/���Zs���T]����U�5�����|�<R{�q�XJ3Enr���Wd�~k�5���?�������BX�*V��M�XQRH»�A�%�2�����B@)o��H�I ��vBRXi��&OQ���n��H$��.�
(�lLY#
���i�%@�ݖ`K(�0�E��P�D	9f�nq�<�u����l�ӛ��J�X$HƅX@�P��cX�sw��w}�V��h���Zp�3�8�x�@J�$!����Z��%,$�䳁�f��tβZ�����6<�a0�DזJ���"2m#*��3���ֹ�qj%�!DY��uF�~٨�#Z�	 �I#R@*�(��ݗ+Ȧ�w�L��^$�kʠ���r�~��
�SB���?
2� ��%���ZᣉV���) Pg.��ƭ\WU�\�l�S�"MU�-Lqn�U�ր�5�[.mX�k��6glqt�xxL�]+�N쬶�9tÉ���7�f���:����𕐂s],!Am�F�4�5Ε$�Ws�6���nFH�� ��0�᪖�n�߽��\��4#���o=�<� TbB$����	E�[�mu����eZ�Jq����z��E�cPD���.���V�%��٩U���+�}B�!O/d�H)$�lȿc�d�y-ᡃ��Ɔ�xa�'N��se�bl�"E�B7N��0�{�8{2NhR!�YUy�eH`5$���$5(��j˰��'�k��C_�@ʺ�,䥁��C�x�\�=!Ce٨HF2S�f�{�l�v��BU�['w���E��1 F�ҋ<)�t�Wu�7���/^�p��N��Y�k�/��6<C2bA�t$��œ�CO�y<��Fv$�۫�Q
j�2��=�7�Ӱ�6�$Z�4�0���Q���{]�Y|���v'Zo�±%���![���MɽFE��l�J!(�ly��)H�1�	w(���J.IVg�:��8���qn4ƌ�6-,p���-q�X��1�H1�Qi�9��B�^:0ٸ�Ya
,�a�7���TI,�ҘoDB*��ٜߩ�32ay�$�µ7�����o6s�K��Qy�[�������DK���rI&p��\볞�񥚐�hH���J�YQ4}A�[��K#ޝ8pѲ�tX����f�g�U����4�[�VK
��L�����M�#�g҅$߈xdP�0�O���'pLX���gt��,�G[rm�9���|�vG��-�(�2!����FұVߩԀfͅF�7zˣ�'�xb�"��H���
�L�s�������C�a�.��(�:��~�t�=}�����������|�� m�� [A��ڶ     [@    h  h  �        ?L<                                                                             �                                                                             `�                  �uJ�6��]����t���9����l������[��&�  ���v�l��ڃ�m�2�dH�h�4&���+EYF��%YV��� �k	 p-:��F��	6�I,�ل�4��-�h�Am��
�d�h�shӮ�H� �F��ۜR7\*��e�cqlU�1oh�
��g��A�&����H�n�]�4�	�<9��L�g�� m�$�l��%s:[Bml��;+ ;9��ݫ6��I�k���@�R�ݶm�$�m�n�		��6���E��%����a֤k��m�t��p $m�Sʫ.�Ut S�j�c��[e��e�	6� <�_<J��dyf
�ts�,� p��d�6�Ѯ :���$�v�۝�����v�ؐ�ڭ�j��e[�t �r]� �0Tnz�bY� ���+s��V.Hq˵3�sr�;[���(����6���)��<��\M�V�ޒ�:�a�y;s�qۜ	�6Qy�u*��q��
��9�()��٨rQ�ls����F��C�)�k��"�*H48��T�1��~��ӌ���v�R�����kp�U`����NG�yi%����!Υ��[=',��UUJ�O<�t�[u�HE �n�A�F��P�j�������}�5����ݶ����on��b�
\�!��gb����\� �9Kl�K4l��CXbݮ�I۷'WXðq�@.�aj�<�1�m�Gm��4.0�C�4\���`uЗ;+�L�8��&-x�zoW�&�f@AQm��n����+KoD	*&׮&��`^�d%�u� ���Wk�K{L6�m�Ma�q�sm�4U�ke�l� $-)UWI�&��TgSD�۵*תU���̽�F���K.$m�j�*��$H-������q�
�F�O+�z���A�7I��4ڭ�6� ��m����K�O<��@Ef�V�d-��b��+E��A�%WY\
B�f��V�Uڎ5m��;�g#eZ�Z��%%��~ݶ~H�Y��mB�� �䨼�e.������	���c�9��J��v6��V7[�Wf籃a�)*j�W�Pږ�ހz�55J�;-�u���]7N��l�8dn� ����Pg��^ZA�)�U9j�jJ�I��6ݖj��8v�����:@6�l  �6�� 6�-�2 ���ى95T$�`�-�^�4��$  -��[dk�ֲ4�=kCm�-�p�m�   �MR�\�ZP�V1������yj:� �l[��mlհ[N��m�vm��,v��614����m�m��[,�v� 8�m�lH �km�m�� 8�h��p�cR�U]J�����*�a  m�  4U�8*�.j�ZtHRʬ�  ���H��;m�������.��m���e�H'��<�6�j�m����6��b�I��m[�������t�[�͙րz�����ko��X[�� �Z5q���Ů��OmT�7 -�K�kV�;Z����p�)��U �ڪ�U� -9l�� W����(p]��ۄ��@�![;����nm�m��h�ۮky'oB�M@-UR��ۍNĽ��E�v�Xd�m���'+=��n0�\�����Z�iV��\ׂ��k�����:�²�չŞ�[�ȈΪ�vX���Wl/,�P�$�6�`�6��vͶ�Z�m�uE�  �۪��wf�7h�,�W}U�V� ��2�O$�3�Wd�M��
��1��iץv���qT��:$�P�/[YRh"'Z��t0�sq!>ٸ�![qƌ'�"�A^���oTQ�[����;gY��Z��J��;�!�E��6�щS���d%���vH
��8Iv8u[e5���{O�<賓�5��N +���ۂ6�*�����<�$
�3�-֔���"�Ԏ[W����M�������/�n/]�]�FgMy���̬t�ͬ[{=�29�;Mi\ml�j�.JVO8�f��W�-��l��Y������5����)�T�R_��u�9��ި��,���C��諸��-�\�Da� m�y��I[�
�l��I�.�{[7,��
kq:zl�6�v�6n�Z�l�aĪ��*��PRʴU�����-u�H*��k1��ltqQ�<u��L�u��S��VU^;N�s
aӷ*��l�����gWU�n�ڹIJ*��V4
ڽ�����	3�l���jhl��  �e�ixᖺ��Bi�]x8�V,Q��E�E�r�$;}��A�����x���N�<tL[M�D��$n�v�@ l��z�ݢ]�bB5�� ���hЭR��P9�U�m�MĆ��	-��Qێ�Nm�݀I��*�mf���U@[YB:Cd�iT�!E<v⧫\m8������m�+(�uUɖ%��[�D܄�U>L���y��l�;2$v�$h�3)r��4�i�R�*����V4P:C�m�:M-�6�	���3%�3j�R���y��-�z��M������d]K'Yգ���V�F�](��ع嫬���_T'@4�X��U�{A��UZ]��j��P(��k+�sﯾ[�S��k���l;��U���/��~�	=_}L�..�]�:p��G^��K�m�m2��
B�z�}�ݟ��"�'��k|G�&�? � %�:[m3�cP3��I�]$�sZޖ���}�j���T�f�I���l^���.�� 6��m�NR�ț8�;����Z�[�t�;` ��m��lO/N&Un�#j͂v�e�H��uVª���~C�⪩V�� ���W�i��Z��[S]������m��sm�gCk�5̓?�vLΟ�*����g0AE>�\���{�O�t��L#�88p�8c��c��'.5�YU˙�1����ŋ����\K�96N8�ss~�nq���g�1�q��㱺��m�Z��XRR�a-q�v<pǍ���{���Q�A�}��G�#��3����2�1��1�G�1��8��1�g��2PG�#�dec<�1��Dw�Ҿ�W�K�;%�/�}#��fTZ5Q�:�;m�Ǝ���:��s�d�S���yK{�y��'d̵a�Ԩ�L���5+�s�r��p3��;)�^'$�mC�v��茙i�q:�e�[EнE�Ƿ���ށ� ��ꖐ����T!���Q���On{U�z��	�S�<��0�Ηu�)�:��N�;���<�� �� �!�� p�"k�D)D�M���G�˽U{��LyS����S�;��+��й)�a�W��ҽ�."�S"бz�\�<�t�d�/���{��G"]��x�@�x*y��Z)��[��3�53�i�rډ�ǥU�<�z�Zb6��=U������Lju;z��Z�4Ͷ��x�.wj{��u�G�����3bn:$$X2�DZ"F��zL��U�Ե2ɚ�P�+�K�z���=��g79�Z�f�ƞ��+�9�� ֍eQ����e��@i�1
U�X�:�^��g��yO3��ne��L�I����>�UJ*	P���RM]c���7=GUN����2]t:ٝ)��\���|x�%/�ڔ��OKn�ߞ��)\פ"d&X[h��n����J���LW��dK�+߽��=z�ٺߍ2 �`!m l              ��              l   .ʆO[^�I���;���:����t LwcӨ�T�ƅrLB����ۙV�$���� �A*�ut���q/,��۳���C�F:�͆���ڦ�i�PxBU�Z��]R������ӛ�
@W76�S�E�5F�A��u�n�]ZPb�u�駄s��4���"7��nz�.�i��E�n@cv�SrSx"�7n�q�M��Gt;m�ځ�b,L�4�j��F�W�[ŭC���wf(�Í5ݺ�����¨i'sv�� p��]umTa�75� @�-e��(�Ygbpl�jeP)v������l�� kA	ˀ�90�җ�4��j��Vnty�]���K��眇E,����U��4��� 3
���+jaH���F��n��l"��(s� Mcx�{rd���vKV��x�;�]i�������Rd ��������ɩ�@�M��ܟ}��9�9M�5ϋ�Ѐ���)��"$���y)���.v�兺���<��￿
������I�ٓx�JD�*QhJm���g���Lu�����c=k��(n�������k�T�<�'q�����L�;7:���4�9�X蛽?[:릖a��-�޵N�oswv�n�W;^���n�}���V0������e����ƨl�t� �V��@��|{@�AǨ[`t@9`�z�$1/K�FT�S�"H�A�p�O�X"�jf�����ľ�w��Ϯ�Y��� m� m��f�ۭ�r��ʠ��,�7�Z�X��v���7!��&�:��WA�RA����ۓ�宀+9���h��T��ŏ��ѳ5��h��H��g�q���]�ET�K�}w��v�Uc�f�< �ApSZ��]��VJ��T[��x<
��3�@2;���J�2�i��)�oTo�x���]�7p�e��hܧ���8c��c�|��7�#,�5p�U���$�j��Ӊ	������Ͷ�g�6����)T/3\fn��lǝk}��uR�N���&V.���(e���U���ļOӛ)���,צ=��/o{2g˔&Sh�����Fl�Q����(uA�'�8hY�u����T݆�HHa��]��c�#'g��d�=]bq(���.���$fjl�5W�7Feɒ�r��F'5�6c��c�z�F�7�m��E��v�Ʈt�]u۳rE�eL���u^����ߴ�z�Ǻ��@�#{���Zq!0��T�1�q�e>�� "����9.A��=�i�a^���,b��^溻Q�W.v9��;�
��Re���BόV��޸���[.R(��U8c=�`�7�8�7P�����m��{mE�OZv.�zIn`�jF�k����Q�rm4bLf��yx�:г�[�6��
ḀQ{��obM�Ww���,c.L���q�hY� A�u�}���;F�IK���Ӱ5�o.o����)!�����h�*z��X�Ӊ�Ѳ��_���{��tq��*�䙕��\����\�)�.���\��jQ,Kp�U��(�,��{��ә�Z$�e68�`�fLV�>�׎F,�KS�&SPӦ*�����q��UM�i��9�Dp t��1{��=�Y�{�6���A̻~��;o��f+��A" ��0xzy)m��m�     ��m���T`1Ј�a,��cm�qnG=��˶ޏN���&�$����v���vj6�j��m['Iؐd�tnҍm�ŋ+�� �fůVfuK�2%s�W��u��W�Ƀ�]%q���U(�m{�������^�UXy�Daz+c��K@�Ձy��t���sM��Yգ9L��,���c�z��7F�Je2�������b�sf���~9�46�HlJl�m�֜�l��g�7���ķ��V3u8�f���z��{�'P�%�)��m1���_v��`� Dst�@D콈��6�u3�m�i�%	��7lՅ&S	xq�wl{��Dm�����,���ｕ��$� ׈�ʸ ��mD	 ����x�����m!��jhfn�eN����6��t!��!�-9Lt@��!�����_8��ѭ�RR�\׎�1�ٺ����f�������6n�.N�̺u`.ݧ1��E�����Ć�hǷu�e��Bό:�'D�
e�R�^�mG����v���:��-ܼ�]����p�H@�z���Z�7y�3ىkfT�MC�t���=���jB�n�MJ0�̙#ۺ�e㎼�O�g={�{�U]1��hh����ݕ�Gk��+�{n݊X�,�әJe��������+w�s2,c.HiKNS��_ 1]�Ǻ�ǆv�l2��2������i�{P�ȱm8��l���=��+5DH`������(]Ըno���+1����:���}�a��أ�$��m��x�r�))4qc���΀�X�\(�q�J�h3
e�^z����н�c�qN�aJFSEPӄ���m��T�Fn�MJ0�F+wX�^8��,���lM�d�(9��/s\Vj�O�=�c=:�8˒R�i8��,�9�s��Ɣ^ĉ=}��ʦQ��       �g]�N���Ym�Y�x����$t<Aي�Q��>��*�K�&{V�f�n�s�T���;[X"�=M���6V8���/n�xܢF0���J%̼ul���$��q��^MɱZ�"�-�aj.���|�y<���m�f��Ԯ[Ut%�t�Ki���|��;��˹�ӭZ8�������.�]��HL&�{w_������"��h��&�dL��5�f��D
�6G���	�$�%��M�d�J|G��m�{��.�ҥ)��*��4E]�=��+5
����ۧ�1����O](��"�u�m��[on�z�gs>��/�q�f� 1�uu�R�$V^�}߳�.��
7 �V�{�Q�{l`;61�$4��)�n��|B���cp�8��ѭ�R)�.��0�vǶ��n��vZq!0�1[��{&��٨x~9��w9�'p���� ��`�^9§^z�t��Qq�h��d���)�!J���bϷP��$/m�9X'P�%�Ӗ�٫�g����W��"�3�qR���T4�wn���I�  �.��ր  ��O|�=�D���*B2J*���c��>Ȗ6����c!�Wk��䖾�jS	��q�u'�\Hv��&�Y\��̯�V��S �:|}��M�Y�	���]�Yټz6h�f��e�w��K%D�h�}����d�F/H�wCߦ��JD��#(�4�U�(�J!|��,"��Մ h�_N�%� h(l��w��0I$����։�"��^u�k����Lb�`���S@�Ah�}�J�cL���s�;������􊇿��G�"&
�?U
�6�lNN;lͧp��ʏ�&�y��N#I�ʸ���A���<i}�����ݸ����d���a�6	���7j=��� ψg���)L�� 4߁�~��L�MwgWI�~� q�l�6[%*�nUș�'"f�M8�#ճ���Biƚ��Qfp�����{~�(��6H�e�8c*�(P�����F���Ӊ	�ъϾ��fn�3�ɲ�~�� �	*ٽ޻�=�a�����l��@����4���qG��;wA���$�_��g���Zs�" �(_���/��cm��
�����+]bW�q��ĺ�5uؼMk�k�s��s��
��=�c�6w����jPP���1��ǳq�m�1�ǈ/�aJd �x�?��gT��hþ�8��D�iKR��=��Ƨ��wc�f��e"��46r}�����߾�}��	��'��F��,X�-��)
%��}}o4��       :M�ɯ,�n�*̀Fm�M��V�F�L�HZs˰u�J�vC�����az�=�V3I����*"K�	��GF����<�瘩�Y{F������a/hLݡ��][��q�:N��LA��W��~�9�vç�U�Gq��J�Lm�yĲS��m���Y�	��Y��g��}�<��{G		�S�)?
���0���weEމ�&Ih��#��a��.�ݬi�{:�)N�^�L<�co{j+�͚��5( �%���a� �����}�y������eUY�i�
�v���8xYB�^��T8�{���i���A!��+��B���x'�� @�g�}�W����K���j�G��� �ք��v��Q��o��������|>a�R)�.|O�L?]�5}�>/�.���鐞,���r�\P�u��8G�8`��9�I�f�K$�bό=�c��" _�6�m���m��2�Y9z�K#Ǵ�<�4K�L����^v~��G��ο��g���;{:�)MC�wvǻ��f�_��6�A	`��x�}�B�u�� ����r�.��k5�8/� �P*�~C�1���Kp�A̵��sO��ڑ�����c.R�&�"�Pf�`
��}�Q_� pD|C����L.�f��s���D�#<vgV��j�꺺�QR�D'6/����{ﰽr=��� ��J&��o����`Vrh���Bd�L��{��٨Y����ʡw��`�h������#�͏�"�E�ňc��7^�:������\����%�J
Sex_I ;�b���f�� 
�����	�%6Jm2����+����h�F�<�&KM�\�!��G�T��}�{����i/nʖ����_w?�m�����<������K���-8���,�v>7}�#{�9�H�e�7:���b�q�� �|��Cu�$���1��y��Ͼ���O���<��HTa F{��4����       :v�]{n��ηF(]�`���C�v�
ۍz1�mH�!��+ӹw��I���~�,�Ű�h�b����X�0NzV��l�hmtm��Յ�`�%�c�zsU�f�np�K�ָ��F��und�=�5θ�����]�^K�'9`;1�u)��<.�NV����iI$&A[K�UB��������D}��5B�_0d�tiUi>A܁[��=ݭ�[{:�(#)6K�̙ d�̯�}�06�Q�k1��BC	L��o��f�a��/����:�hjHK	5Cݺ�=�;�+v���m�ܨm�`�!�{����:�'��yH���M��*T�L�)jZq��c=#��b�����5�H�z��#�G�Q#򐉿[�Vt���BStS����^�Ik{���߽����f�FcN$ wv�W��< ���g�
��������S�}��s����j���n����a�cA#o��� ������ko4�Ͷ�a��K؉��6g�r�+M\�]T��at �-*%����I5��V_mP��*�1��BC�3����9 ������43�=� DH�}���MP߾��{y�`Dp?P@����β�QrI�]���t�%�JZ�����C= {��B�_v�^�a�R)���v z�(Y=��=�NG���| 4˪\���%k��m89���J�����_K�
��#o�����t@d�(�}����)4�ݯ�m�����w��`�-ܷD{y�Q�@�9�}����33��A$f[3C�؂"��}�����*"qZ��Q, H���_Zg�;�!����*d�vwP������A�����w�X�m��(,h��[��~�|}�)��/�C�m%��w|7�=dx.�������1&���� 0"G����ӣ�.RԴ�>ς� ׭��h_<@#�p�e%%�.hvLa�f: ����'��5�9̼j��2���J�T>ﾡ�{���@� Gc�������߾��ȊZ*���׻a���g��y���� �@n�Y(kH �\��	Pd$�$@�����W��$ѐ吅�se��%_�7�4�x�����1�L��;�hu����1�f����v0�q�E��c��,if��w]�\�Ǯ�df��\��(���E���d+E�1����1�06�b͑���wɏl��{�W[� ֬��S�R�Ō!7)� ,�:eZ�c�!�U����B�%h�!Ƈ���{Rބ�5��	1 ߫�	D̓�!�.d�tm0\���F�(
��j�[jm�                           �       �ô�wv������w2�	�g����mۨ�R^Nќ�kZ^�<�sgg)�f
�h�;#"�]�q�O9;i�ԉ��*�GR1i-� �af��t���b�|�ܞ|�{<Y8�8ݲ>ܳ<�im��͂� �i�I�x3���3n�T��x^.V�nV]u]a�=�iVT,�:�pg�84�N�����u��e]�]N=S5*���8��n:��m�u,�4��ൠܮ�k���k+7+.�!�۶�~��|��)j�[l#l|�1��'ml���L>6��P!M�VT!�u�t����UPW@�bIP� ������c���6��>�\�+�e�����,i,�+%&�6�{i؝��&  Ae5=Je�/%��D�6�q���ӽc�BC�b�t�9D_D�l�������,�\�VmR�~'M�v��i�-�t�GՓ�j�˞7Y�𘺖-����ژ		CLIݚ�D:�KR��k]�:6��s�E��*]�竀ݥ^4+� ��.6�l�pT1Ngf$���.y��G7IX�B�;�|�����^ߤ]���ԫT���VJܬ��d
t���V�!�Ar�٭��_W����m�l  @�p        p 8m�Ͷ�m�m��6�	z��S比]��(ܩ�V*��uK�<*���@y�����C�9ɿv���ގ��~e�mUUUU@    :dms6P�)��@NӸ�3����?��[�c�ݼ�ݧ��oU<���Р6�;r����@�f��[c�v܂9�e]����##��*]��k���륥���[�n��[�4�Xӗ[�GL��f��d��������f
A��`�,����v��̎�Z�"Y4qc�����vJ���8�C�I�eSIa��(���#��* �}���3<zPI�=�?���n�9���/�\�g1��II2����u��"w>L����P�@�*��~ �}^$nrS�  �{��785��-KN3�����o������=���456�E諢�����sl��160��w�M�a�R)��òx��v�_k�  #��35�8�K1'	Ͼ�� �
:D�P���Ƃ�pV�z��o�w���'�Q.Ns����R�*��ﾢh��`DE�\�7ݬ]�kIi�)� o�y�����  g�w��͙�|e	H�
��#1 ��T_v�#o�ӹ�km��	�&Z�j�0h���׊�	C"�t�, �a�$�g�ٺ�o���"�܁��45	�C��Ɏ  F�&k&>��U t�ӣC1˺ˬ�}߭���*X�|)� &�����E��k2��-M�"}�] wu���k
Ǆ �w�F��\ӉD�S7P� y�z�V (w��k�U��p!��c]����F�����rIzYԳ !9�^��q��+$x@ �=ݔ=z�\��Zi�h��. �$wc��b #ofw�BR,5B�@��x  }ݮ6�Fn�e��a)���'~������o���������L^�~U�[�" %a[x��I�??9��� @����c��}���3?6�m��m�$�kASr�����vʋM��g9�sn�:�x�_���vb�9}ۖ ��gS����0�Jr��ѿQ�K�������������F,N%��Q����* ��&d�"��P��'3*�D��Dm��$� Dwcz�\��Zi�q��w�$U7�~��5��q��dX��ow�|M��/}w��m|      �7\慽v���WP�ȗ;<�WTC ���r�[6ʥf�9EI�6�R)T�p�//j�t�s���ZJ���H��X�1�g�UIM�bՃ1��`@X�]����m�m��Ix�P?+�;[���333,��̱��i�������/b�H̪�c���k^�p]��N����/wX���@�!�~Cp�k,��,%2��^b��b�B ���,��4u���|F�&��=��'��9R�ZcD��VH��3���=�Q������SC� | �������7w�y<�i2���gq��Һk���8'D�d9��oӸh5I�D�S�9��{7Xӻ�b�@������!9IP�v������Z D04@��Z�x}������K���2�)�����H���=ݯH�;�<���M��^��@*�e��� �o!^ı��J��S#����w�����'�_��y���:��3)Y16�%D�ܧW����J��ʔ&C����Y�w�`�|�l��a�T���{y}��}!�{X��k�M��y�IK�sG>�����ۨ ������u5�O(�D��� �߱������5bp�,9s� NoRf��c��g�����`o�v~(��/*��zɟ�� ��Md����ܱ��r�]��3���r��:F�:�W=F�]��a���LVH�2�D@�@��j6�ys		H�/�� TEfc����� �@>��e9��aIJE;���f� D>ߐ�H�:�,�@��T=/{�7�&�����t��_��C���gA�CC�s-8��q����������h=�6�r�-�N��l��FQt�SN��f-ވi3L0�E3.lg������P #��{$b��"X)��ە� ޽b����h������������Uz����j�}�7�o����`�)4�1���
��[����ys		H�W��*�({�\Vr��3 FUZ�2�      MU�&M/�ol��T��hŻvYx댶�-���U6��` �i���Ae�����5���l�QZ �x���n��S��Z5��\��f����cq�6m�d�k�p g��u�P��+3��V:պk�$��ܒK���:U��Ռ��D�'\�鸱̝��98�_���(�RK	L�6~ŷB�Y`g��>��Y�e��	5C����#W!Y {��Tx�p�K�i�}���c"wc��Q��+K�S2�tFsۺ�v1��	����8H�
`e��B�B�n����B�@�O[m��g��ĺg���ax�w���c��չ����2Bfۺ����Vj�p �>�ܡ�y0A�ĩX�_�x�m`�V�!	�
�Ԑ��u�GDf%�S "�(d�B�L���tܟ������k@�Tv�~K�BR%�.�t�N��DF� �}�T_|��ݲ��$�����b�1�f�ށ ���5�`�fP,$ѢO����� {�D�jfO��zI8�N̶۪6b컵[=OF`�-vjm�q�ar�s��9:���1�Q����Nv�I�Azd�y�� ��� y}�D���_H�2\�$�PY��d��3}����@"�9\�$K��4}3����7{�FcO�$A'j��rB]$$�K���W�ԍ�Ο�
ikŐ�f��Уu|�r��;�H�!����)�
a/d��*�[��h2��0���ej�]w��jF��0{چ'H��t!W�:���`���Umg
u.�w[ ^BB����yG�kG7�P"��m��D�sz���]T:��| ��@�GǮ��<	;W�<Uw���oW�������ύ#�`.�ة�� #�{$ױ��&�n�		�INL��>o��EL��d�b�ϥ\�Mc�`���JtI�ݪ$��KjNyO�����>���~UV(��3���mYħ��]ru뎎�/ܜ��ۣiv����`;�g*I�v��G�!a&��UkWs(�RK�I����$�n��H�����aU��n�3,�BX�n��59�ޢO�:��@.�'>ZY&�_Jp�4fZtN�w>�I�C\���M� ��A�_M��߻�$>���a��L�!�'mI� /$�v��/��9�O���UU\)��� ��^-��l���@Eb^y�����Rp�,)b�=����7��G��ށ g�;�"Mf<<$&A	��>$��Uӹ��>�(��V_�"���%|�.T�D�����f�J< D��,,�}ݵD���J�BR,4������Q'5�I��ʢN_͒s��2��$���D�ե�~  >�u�'���&�
�����T�.	��j�?�g��0      ���]a�-��07-Fu��.vlm��ѱv�	.���EY{F��y�,�򫜻�l�kc���:��޺��9M(�k��b���$�ې:�n:����ܭ�n�t�]ٻN^�cc���ꐽEG�.۽�۽�{��Ӝ�9�ӷn�UtE5���+���*|v�;\��\�63N?qM3L�&P���#�$����Qs�|�����_����{񺶪tvgs���'ӥo�I��؀)"�w���)Ж�z�nqqD��vh�DL�;j�7��',����`�h�s٪�>�ڢN�6OD@�奒n՞ ��ʚ$��j�'�s�}:Q&�vM��y�UVfJ�V�260F�帩�����5Ư���L^�S`��Iʯ\�y͒}:Q'�H�� T���$�nl�VR�l�d��)G�>���G��1ƣ�3����D����������N_k�O�l��{KY	�!�d��w��$��U��6I�҉=Jʹ.L�,$Ѣn47�ɩ��d��I�l@>���Mr��paÕ.e��}7�UT��Ҝ��,,���'f����} �Xi��dҲ�e�r�b�Ļ��w�6h��E3._�7<Q&�Yd�]�]=$��y3�o�R�t�f�9ˋ��<�*�d��d�N�q&O�Y�SD9nQS�RN}��ԓ}�?��~"","�*p >B�R���o��o�d��s����+����|�w{j���;<">�Q'wg�����l�D�N�I ^P�O����y͒k�X�uO6�'�vpt�t6���0�V�n��9z�sd�s2h��o0�>�ڢM�?���M�I�֕�X2��hQ97���DBG7�:��W~�1���y���=�ݚ�g�K,D	�׻�,���TI9|V�H�Z�螁&�I�c�]٭I�w�@��sH�@u��~u_��$4�Q,�s9�I� {7}�{�T�w��Un���Zצ�s�BN�^�L���j;K�$�^�t��6��v����o52I��� rO��d��^�%sL��:$�s} G� @^ss�r�vh�����  H� H�t����[):��D��a�6����$���I�X1��RKHɢtD����k7k}33�͓_@�
Do�$�k
�,AK�3�fo���)� ;��쓓�}���?��� ����vƺ���VJz�=wʺwϫ�:��      k2���t�Ӡ��,�ѓp�=�P3	q6vR�NP������S�b}d뀵�v���8:����Slrp���;��m�\N.�t�]Z���y'���2�N{^I5��E�Ҭ��2��-��X�����ԡ�J��9/9?�'$hu޽����*�$�"���.B�ΫP3J]�Y/_�ɷu��<n��{;���l���Q'�l2Mwd���*��S-K��9<u��������9�ug��w~n�L��9rp��`�h��Ҹ�I�̪$��d��<�ɛ�g�R�Җ|Ho����L��d�N�O� �}ZY'��AM�&RR�����K���/��}��t����U]2����UE�h�tr�.x�n8?L��Ѵ�v���������+��Z�_6I�\9��RKEL�ک���g�~?!"�~G�%s��sz�����E�{�<��w�7�B�^+�]�?����9�ӟ�'�k�$����7��Q�Æ���O��o~�I���$���y317ݾ�I�⸰�E3.]}:eI;��u�6I�w���7�6I�d���m��jQr�U��]��
��>:&��[��oZ;��`cD�O>��ս��^��R���}:Q&�n�2��I��zd�wUx	��͒_��I�s%����z�`ɔ��D�f�Q��N�����Onrf�s3S,b����!�]*,����D�̟ĩJ"�J���&�I^���>�ʢH���5k2
Ih#&��id��ٻvI��w��o���?�UY�h���U;:��J���m��L��`�_8�wXKt%bT��}�]��VI�5;r�;;��a�JZ��r����$nx�NO�7RJ��o�I;��K)�n]}:Q雜�g��W��TIί��+ŉ�D�[4N��8�骙+}���T���}��ÊxGp
a*���ʟ�O�}z��I7���K�bI�.h���w�I��@�{�2nx���[����9%�o�Uvlb��,ێ$��뜪�G��R�V�1e����k�����	���I���B �\��}��'sg�0���e*$�t��� 7;��7��Tvf���` ���/���$���$����M^eQ؁f��t$��ޔI=�娲e�m��~��w��{��}:Q,D '��I�]��a�JXR��&��$��D��e���v����#}���A ��ݵ� &%� [��;4����fx���ӻ���ã)	�0��Дu�Q*�¥%V�(l��(�BŔK*ʺ��Űp�M��a�t!d�a��h��D�j���lm�R!6�!$cɡ�L�IAxla#�����!Û
��{[��%��cT�cVL�"�E1Wr􌼜]*�<�d�h��$�                                    �k��9;��{f��X���ʱX�iY�y�f��3$�`�q�ɒZ�s(^���Ų�є�z��B�GN��h�ݦ�F�����7h��M6���L�l�Bi�����"tt�}(&�ܻ�H�Bk9�x��f��^H�)�����Vn׀�#Q��a�/`��a3�5\h��oak�#B&I4�Ud��n�2r��R:3�۫t�ƶ''�n4Q[8�[��TT��Rz����sY�p�.��y�c�(��D�8l���f�mJ�[�������@�R���j
���.pN�)॒%��a��¨r`ղ�r��, p �鶘�;[�m�k���f+�ܩ�!�KaH^����sn�;ul�99�#6��sCg�`ܽ����ZD�f�M�V�ηn!,N�]9L�57��_����ѷ\6�I�GP.��"R��jMlA����6�jQ�^"-nb���2[a�b��k�3�Wݿ|}���MA�C�#*��"%)f2c�y��F�LX:4.-�U�	��.�(��t�h��[�n-��U�.v��[7"p���*�3UWi{�3�6�d\\WaZ�>L��Ԝ]Rڭ

ڹ������������9�������GGn#,��2�;;:vLٖ}�������_B���W҉�砟B��I���E�y���j�*�8�������P�5]k333      ���z�mrݞ�v�Xy�"-�n$f7[N��m�@(kz|�b���NF��s���@��ٖ�F�R�u����zf��D����ݝ��5�XHUy]����9�3^
�h4G8���6�zE6��33舨(�5N���O1��୭Q.���s�nH>�����o��)̹u�M�Ic�2jfO�����3��2Nr�8H�`�f�7��{2}���&Nn�I�Ҿ }���ì�pRiK>���}�Q's�'�*�
$�-,�C��pd�fS�o���UI7<Q&�0�&�I�v�ĝݞT�Bd(a�D�N�I�ݤ�5��D�^�I�78f�m��av��6;sv2�B�:[$XM1to��gIjǺ�򻦍^0�mW�$�sd��҉6 O\�˙*��kU�rN}����q�A �������2K������+��D����.%"Դ��Ow͒}:Q����d�wmQ'gs���)�j_����L�XY&����;�L���%��EK$f�9��%O���'s�$��G�߯��&��[Z^��oD�����:U�C�>��??U��h��NY�Nwt��M�I���� R&�|Y �Ϝ�%L�tN�o������s�r��h��ک��@l�t�SF�����o-;���B�C���  �	�H��D=y���OvuQ'شk!�����D舉�|Y'ٺ���9́���w���u�%�4E;��}�A� Dު$�t�Myqd�{�Sm��D+1l���6�
�]�s$��k�f�1��.�^���<�l��-(��\{ �"m��zd��<��B�R�nx�� @�.o,�}�TI����7�j��"��,�'5qL�f�Q�&s~uRL�id�Z��D�NY�~ _�u�'�͓��l�& 	�A�	�Yv��a��r��+�_�5������Z�pﱋ�J��蓛͒m��Av��M^�t����U�$�j���Ξ*�Xz.^��fy���"
BZTR�VI���MyYd���0M�I��`�C`���̚$�-/� 	��ݪ$��d��:�ޜS��(K%�����\Ҝ�l�e���?����&�����?}�Zw}(�����̈��}D��ǘl��f\�$��,��z�T�O�����8U\���9<$���E���UUUUT    =OTK��Ō����1�"����+=�Ԙ͛��t��5�@^�͑έ;t;e�.�˺� V����.�g�Vܖ��{k@�d�r�c]:�a�a81�JsيЄcm�:��in+ׇ��΋.�o�w�z�[���f�"����]t�ږ�*��nU�M��cV?wi����=��$�s� D}<T��2�����rÖ�r�sﺫ�&~���Q&�D����]  4po�
�J2�w�l��-(؉���$�vUw0��2��j"|��\��I�v�o9�MZ����@��������I��9�U�2sy�O�J$�o�y�6��Uת�M+#�w�y�;�$�F������s�vh�ٲN}��D��l�S��Jf}k�53��2\L���D��n�""��: ��Y�$��W2{,�]�U�pH���WŲ)�r�I�/�$��\�}��N_6I�C'	,f��k�$�n�����58Q'��C�n��N��}}��n�o?W���(�x���zl���ͷe����7]�Y��U��Φ}�8ٯS2�r��MNrO�q�*I�v�9����yJ	�^7�l�_�����Y'{v��y�|Sz�s(�(��D���VI5��Z� �"Ȅ�����9[Z���4-�6wb"m�7��7>(����`��[>'�wz�>��O�J'����$�?hZ��tus���@��������ｽt���ʪś\Uc,�%�j�Ų��l=��/m՛��M���_[�����?u�;��(��fsy��7�j��"��,$�/����$�|�ٟN��"d׭��nI�-����w���gӥ����Mx^�%s��Ļ�} 9�L�[�L�o���:�hJHH�b�k첄z �3=�tI��:����)Q'ӥ~����T��w�fL��TH7$��� ��ڭ:i,�'6�HvK�5h�r�!�r�gF@�ܧ4I�\$�ٕD��}RO�J$���A��l�'��U3&�[$���I���H�?0���e��D�����S���2}|Ù����d�ϊ�.BE3._�&bmp(��^0�L��j��@ %���&�iY.*X2�o>a�����뿦O|�$��D�w�@�0@@X�b�ZG0N-|�ǝαlץ��jm�    �Z�^&�J�r�ݸ.��Ӥ��'KZ�Kj�]��/�l�;��3�H�����6�e���+�pMu(R��ҭ#3竂�u5@���M��PN줆,�ƻ��
6y��;k�&f��:�7��{��u�J�t35 M�a�9�'4�/<�O���%B	:t��'~���&�$���4�}|�$���	\�d9�N�7����9��9���$�>گ	����~K� ��R�&�''ה'��TI���5k2���i�F�57�A�}�ʢM澩2�iD�=��82�E9hx�}�TI�;�@w}0~�_}⪳3UU6�$^�,��u��0�lm�"�6雤[�5s�{��T;���ϭx�O{�}�O�pr�*Jf\�>헏�s�K�O��}��֪O��^����� �9ˊ�p�RÔ(��������L��٩��%׮��nI�,����TI���9�?�W��d���	i�˙�����͒~ ��$�,��̪$���6�m��I�� ��fۣ� �^�\�J�)���m��tͦ������B}k$�ﲾ��No͒}�F��̠Z*E~�$�n�o9�NyS$���feISI�ݪ$��l��D@#���	$a'뻺
�
�!�Ӑ��?�T	��h��Q�P�e�r� �!V�"0o��Y(6�B@��f$(��t�������5��B�FS)���&��y7|�E�f��C7�vBvt��ܪaP	��n�w*�/!yf�FU�F���fJֹI��PC�k
-
�T�n�޺nvY�v͸֚�cm�sc.kJ�c4M�S4�aP���5d�*�yV��~�{W���黪�*��׍{*��]��/0�������cC�����`���4�n��<���F��@����6;t�T>���a�z:�%<^z�ҽ�x@iN�<'T�zͽW ^o���A}V��	�Ӹ�䉔���0$o}L���1�f�a��,_o��l�\�R��eˢMm��?D;���&�����/��yo�������%lT�h�\M3@n�c�s*\55�T���H�ci1�No0�>�ʢM�>�2gm�I�[⥸A&��D��گ�������{D�Z��dؾ����L�3)�'7�&g<�$��I3˷�3�'�"���*$��a}k$��o�'{Q�
E# {���f	��v�M�`�QrP-"�7�K$��*�7��'<�$���6�l'	�l6�[c�:zB�T<):rk)�b�+]z�n���{��@o5�ON���\Y'��,e�(52�o9��d�!NI���d��ꯀ����IL�r�ڂ$ו�I�X���o7S'ڴ����D�-oWŒsw���9��z'q�K�+�\T�$Ӗ|I�ު$���ޒ{P��7��$���j�4���4��GX�g;���o'�yֶ�    � :4e��l���kα1�Bms7c Cp];K�":Z[(���B�h�R���+�"Wnh́�2�f
�&��l�͞�9��r�`;= �v73��;Ht
��Nr�\u�jG1EQ�$m�43�BI��{�/���X� �ll�4�6�\��g�}�u;ۣU� }($�Ii��fR|I���9h-�>�����[�Q'wD����Re����&�ad�u�Q&���5˕�p�QrP-"���?�$�f�g���33ڂs&�~s�r��<Mx�o�ޒlsڣ�>�a��D	����O`Z˒&PaL�D�sz�4$��2O��d�u�P��7�*���i-�9n\K��S��9�k���ڊ���ؕ))s.]w�&gה'��_ m�u|�'��\��T��
$�./b�0��RB%FTnok���r��7��&�I�.*l8A&��D�^�Q's[< JuIu�Ɖ7{�$��e�E'D���2Nj��qd� O��~�ov��RdO�2�^'Ӽ�$�}}�,�쿪�?^�rM��m��	�v��r�r�UH�X9"�lKtq��L�"�AƳ��k�D�^mQ'׻\#�I�A\�N)�Kh��y�TI���7�"K���O��M�4�裳�y���1g9��CV�����^L�k|��RN�pr�%JJ\�oĞ�%Ҳ�5��~� �}�y�����r�R,9B�>��d��
��ݒ{�j�9�"O��\��m̈́��B���YG�ψ�[�9���l�x嘷�a�ݪ$�kڒsV�	>�c*I�צKN&e�%'D�f�	7�"K�b\�^ݪ铹�g�2&�2��N����a�k��D��l���c!�P-"�d���I��ԓ��d��B��$
����6	%����O���p
��!j��T1�5;� ��"z~Y��t4P.Lx���U9�zu�Mb��id�������m�,����=0Gi���:ȏ��s��M�������ߔ<�$�+���n3���TI��/��))r%�{@��Y'��TI���BK���R�BǫN�T��(~�@��rY&����!&�sD��ڢN��'mI��K$�.2eFIdN�d���9���id�n�Q%�D�9�iʙg�      :ӵ�ZY��&�ˬۆ���̠�CL\G�ܻ��c�`Ă�a�O\P>1[�Gl��C����JEP�u�9	��-p#��]U�L��d�Z{,��N�m�<'WU����B;��P�Kɻ���t�y����uQ};�eֵ�������ۓ~��}�Pv��D����wPD�J�&�ۮ�����k�2��@�T�$�֖I�fTԓ����'�I�̜+!��a����NwuQ��@�>hu�D/���F����蟀��'���v�D�K�$��*�',j�%JJe����v�D���$��W@{�����ꪹ�M��j�v�9x����bnHk��T��n\J�4*P�&�qd�feQ ��j�L� �5儬pe,�,�&����{��t,��Ok��On˒f���}�zdʇ%�e:��OoS$� �������&��]n�O"dM�5L�v�D�J�$�w*���M����p�S3(ʑ�n{^�I�Nv�Q&|�&g�|�|����؍ӵT7�O�Nl�$��$�W9��z�7P�A�e�d��憎9��'<�$���rfqm��9"e�N�9��'<�$����d�v�2w.a)Ir�tA;�\�z�L��H�����L\����!$XDb�`0L���s�ԓ��̒pbÎ\JE�(Q='q��$��׽$�6�9�'Դ�n�.\�4I�ݪ$�u�N��I��xY'�����`4����y���z%qzf�f��fj��[rR�4H\�m<�����Aoˏ�"Wv��;�"y"|i�{_ "dߖO����s���&O�h�S3(ܴ(���2O�2���	o��'m�7=se`eJJm!�NwuQS9��=;�"u �� J�A�Q%( ���tT���L�T�w�H�A��u��:��v�D��0�'�}����ު�]��FYfE���QP�^Ů�_���tz\SS$��y���;��*� '��$�է\����(Q'E�ЧA#{�TI���9��L���V82��M
$�wUv��Ny�&��2M�>2eC��2�🷩�v�D�\�&����T��ȝDȚ�j�;�/�r}i�A7ݵD��l�"��f0A<�R �.t��zw��kz��p�1�4�M1�]�/<>%��[fX�5�����f��rłW�5�A�I ��d"#��,h���4�cݏ��*Y�U;�e��o|���2��[l̑�ĺ�7C(�iXfe�BU�I�@1aE� :��M��TJu`�z@%��.��J�e$:�9������V�Xk4Vڛ��^�W��0=#m����f��s�Ʋh��o}��m\��,d�1���#:�Ω]@w�����0%v��wsx����80	"cmfkw��L��3v�%C�"@&�C��p��3"PB�˔J�`w��Wu{���]L� 2%6^���&�����7���� ���                                    �nݵ���&)j�Vqr#he�\�	p,S��zc�9\mϮ۞(��I:VV��:�t�v�J �O�'j�p�jIg�75��v�����;1@>mh����)��kCπ_�&mw�v�0�z�vH�t1�����LF�NY�X�f�bα��qժMף%Ngbu�`�lݤ��&��<m��A����1ڼ$��O$��u3���G#�6ǚ��v]�lqty����]�&��]V &Qt�k0�Hm��Ұ媵e�(�8�2s�[�*���U��P�ǵ<�A�jk^��n�*�-�p�A�q���*��3� )�Mp%H@+l��֎qD�����;h��bN��H5.��}0�Au6Ѯf,� U���[�A��V9����ڝw;@�ףW����"Cc ����ڻX��%�|=T��;Gi�[��X���C����j8��G+���k����ܫFʴ�n��hU{�V����TU@��@Np9V�!�Cax8�)�ݳ�^v�N�pGv��m��9cX��  �rc���Ӧ�Ѩi5�3F2}_mCP��o���~6�5Fbx����[v�w�rKSƐXZu��fk[k�F�I'��O���&")������S��	ЙI�uJ�XZJ��*���8<AEw��w�ʬ+d���      :v�i�K�룴�Dо��;�z,�v��zx΍�N�f�k$$0v��1���۲�E��Z���.aj��QG#J4i�H���b	�=u�z:���\��=�X��6 c��]����tt�m�Q\0�NI!�z�n�Ut���K�6�  ֑�+�)p�,����fe�R8����O�2��ٯ�I;h#3?O�:V�T������}�U)���P<���|7�u����F����'Fkd����h,��ܪ$�rF�h�RS"[�nw@�ϭid��ڢOf�I��9q)K�(��Z\̟��w݁��)�o���}9xC��Un�G-�u�I�Y�#���y����%ë7�����qZ������tuo�z�wޟ�N4:�| w��}m�h��ԓ��2`��@U� �u� �;j�$�fU)���'Q2&�STNNk�^XY&�r���oU}kF���@�($(��\]̟cʢN�I�AT��{&��ʔ�[��&������U��0[��^���Uff�+vе���`v�<:�]3����E��lƔ�5U�!��(y�73^\z EI7ٵD���}�h�RS"[��g�D�J�$�vUw5�M�X9q)Z�D�Z��>�ʢ�z�t��R��Oԭ�2I�YrL��*�F\�f��DM�w���͒kD�^|~�&��>��#,���O�͒s�It����n�Q$���m��I�
D�rt��db]jܥ���:���1s� u��2n}n�$��i��w3j���z9����3I�Z_� ����UU�'���O�I?\ڛ̠�٢M�r�$�kg靴&���N�X���&Pm�����'we�3W��U=���R��}���|�|���IW�=���~;��:�|�@�����Un�%��ѭ���@3��B�������P�9]�.��;����<󮊙���I>�&���n&Q���s;���٭�s�)�.���C�꣺�'��2�r��'���Nyz&k���7}�������"|%JMU̞�&���O��TO�'���} aZ44ʔeH�O�qd����A=��'1I��tB�-�ڀ      I��kvL�'Y�o�elh�v�#B��71��&೟ھ�<��kY9��!r;k��Ȱ4i�Xl�1�ݻ<;�*TMٵ���\�����9� >{]ɌaE�<et 1���Y4�)jmb��Z����YƳ$�b/]`��6mKӜ����}�}��]�h���TI������Xd��Œzrį#��E��OWy�|��m�߷j�2�q��ђ���KtI�A\ɯ&Y'�ݪ$�kd�V9q)�
&g����7yUE��kd����i6�L�ї,�&�v���6��x��Myid��#�y���UW$ѭL�䖎K,^ו�<t��l����b%��?{y�M���qd���Py����<�=n�����@��D�B*���"�m(~�v���d���N��RČ�ѡ�T�[S"�7k�$׳*���׵$�*I.�բ��K-�铙�TI��.I�Aw�|h����]�C��=��(�� ���{���t���?*�t��R�Q��c.���M-9N@��X�]n-Ͱ^������{�>��*�'s[$���\���-oI�fW�$�kd��'��	��er���Ψ����B� �1�Js�""�=2�e��z�s$�ݰNK!JtI���7�[�o�K$��*�7x'Q2&�-5D��'Ԭ�Mw�t���~���UY�Ҩ���[�)NӨ��ָ�G5�ֺ1ɮ��C�<��:��:�n��$栊�/��h��A�E�D��ڬ'u"M���Jٓ��J�� �iߤ���&�I�-,�^ݪ$���\T��2%��O|�$זI�}�Q> �ݪ�>��I8r�OecWs*��$�֖I�fUw5�M���DM��� �x[5֗��ZX&��g�gѵt�1�Z�گ��2�Ϥ�߾�$��d��8����>�Ğ
�B���u��Nj��/I�n�/�;�"y"h#)� ��'+�}{�D��l�~X04ʔKs2(��ZY&��TI���7�"IۛV���E}{���|�j�9�%���f|�����j      eM�i��w�<鼌��<����][x;;�\�����Sd�\ jm�ۮ�n�f�Q�k�N7RV��]*h,��: �ʫ���Q�vgmUǩCu'B��f�#���Wo�{�<|l�0�mvĊq�믷�>[#'���ޡ�ν�s�r��{�U]1��n�Wt���I�v9ȏy��_UUE��!%���Ng6I�A]-?��țϾ�$�{G�6JR�K���'yB$�VY&��TI���>�r�R-Kb�5�zh�>��Q'o[$� �.��m��2��4Oы'��I���7�#���D�ށ��h�\�m=����`��@�}��|�����6b���t.�Y��j����ƲeX���m�pYz�sw`{�}o]�,�뾪53���rՌ2�%�2(��_�f�,HAJ)�����D���Uw5�zsX_ �d���Bfe�-�$���Q's[=9�"Mys�I���2B6ZtN�����[$��"K���3^��I��0��L�n�9�K$ז�>�ڢN�I�7���cF��Թ%�
�vm�upj�����S��<��,���,�^̪$��ٹ��'�ω��e.\��9�UD����oD�KK�[7��49,�)�'��$�!s��=FUU�˃r�H٫=	F��6lnn79���ۚ�j{�hBPWɣ}0M��=�ș���X���I��"Fffɕ�(�t�{�tM��1��*�����]�T#9��8Y		L���J0��3p�×E�cAd,l��h�Mcl 0��5���/UY,�J+?���^"T
|�*�Aj�4D�b�Q���<(E�o��[�@	��O�bq"XE�(t��W�	"���؎�qV{F����mL���۳�B��y�{�J�m��'j�ɨ�o����Lp��3�.J\i�(�6��4�l5S����x�"���U\�Gp���A�Z��j�D�3RZ��7�|�����	J�Ȗ�6�u6G���=ٮ<3�r�l�����C������?s�hP���4D��-��J[i�b7�b\	��|��x���K2��1��c�@�>���oyS������a0�0��l�V�D�3]%v99���D�9,�*����53��"ku��:���-9Qy�|�'�:b}�}C�b�E�>�F����mL���=yob �j��U��������Y�Ͼc/z�ء����������!�l��~��9߾�j�XE�=F֛CBs����$�I|�[H�N�UP     =-�qɵ����Y��h���%g��Gٽ����!�:�6��wZ��'�.[Vw��/��%0ns���7&�7�;Q�m"�]��6r�5M)y:�����v�u�<�3�Pu��V�p;f5�����I�~���*�Ŗ�'3ͷ�E�.�$Ueص����,��\�1<��ld�a�.w��f����uˉA9j��x�{1��Q��N�m8I���1��c/�y�
>��q'��%��P�� }�Tf����c�Y�<��("ӕ��
����c�u�sm��-������汔lN�Ln�f��#�fE �Aʒ[(�i��b����!�Dy�}��Z�rP!��Y�}�,DDD T�yW�������v�Z*J��;yi���~1�����6JR�2%��"��+ӆ+��u��9q("\�C�:l��ڡW�=z��7��UT>��w�s�;$\�y����2l��[S׺�{z����@z�<9)4&]�\D�f������ @7g��ʗ�[����o|��̌$"B220��Ng��� ��z��ȼ��:���� ��D�����������6����{Q��� >���m��L)M���Y��\K��ٛ�u��������( �2�;7�^j��"k۵�q�d�E�-���K�DD*^�@Vu��8�  ��r�R,�4/���c��={�W�IƜ$̙N:>��ߘ��_��Ya�N�e	�#.�0�e��B*/y����! 	L��p��C��R�mꏯ5�w�����ϼ���UWa2�nV��F��r��؜�+�?�(KFA��iˌ�A���{�X�`Qu�CL�@�&h{g&b�x����C�,D,&�A���C舁�@�ϐ�؀���+*J��ʡf������^sN�ɓ)D��(tD~U߻���~���n
���ij��^��z�|������j      �I�ۍ.���8v��7E���]$�M���M�荷ۗ�m${R4K�&�LvL��ҫ���;�������)]I�cF�%�D<է�;��s�b ���9ؗ=M��d˓g�m��S2���F����97����B����K�a�V����TӥM�h�q)�- ��q)^׬������ '>B�?�8I�2�^|� #���/>�+䀯{�?K�%*��=z��[���^�:��h"Ӕ��\}��'o9�z��9e3)�sB����f,���Q>�6�*�m�	���z�=<��OK*��sj^��nۋk��f��9��=�~i��+�G��+Y*J	˕C�S�� ��<3m�@_�_�D@#0v�L�A�ME� ��>?^|�^�c݀�p�,�C���@ef���6��+���NfL�^s����A�  _����m��,̶���G^]�әc���'�n�w���D���2~Q^�A��0��B�bu ��NTW�~@g�z�^� �̞CYL�@��P����|�lT���Jv��^�]�:;,D�,6ҏ�����dz�Cb ��/�6��+�*J��*^�� �7�{��^|���+m�("�4љ^���F!�I����`uQ�T)t˦�;����>>��:�Ev�%�*��p�DH�ږ:�G�����N4�&eʖ@]��2�E{�{> W���%�)P�@��׫S_U����BE֓��vw���,z�O diʋ���|c}z��������gp�B�ܽ�[��^k�%,<sG7\~�g��JL����t����/� >�/>A��V�r�c�ߟ���_�'��;�bq�(JD�R�m�� �|@�^�"�N6L�a9�V���6�X���QB���p�If]i��1V=yC�uEe�F �Q�UU�����{�$��\��ct�i�L�^�k��J�ɣ_���޷�)��y}f��|"1`��J�5y�h͕�5@�Z�+V���7DI���_(��1�WWH��;�_{�Y("X�/��t!��F��Ü�C8� 5�0��ìG�]�R�-ݐb�Tf�07a�+SAt/!aV�$%TF� �I�����,�9����D�l�������|&�� p��     ? x                             ur=q��r����v�C��%j����۞����lq��M낭W>W�fwI��nEI�-;��s�Su:��Ul��\�v�l*m-��f��-�8[����1S(jLe�#	p������nʓK�l��1@��,�E�n;:`6�)���N�Ӊ1"�:Ǯ<��u��^r���=ء�m���:Dt�%<Έ�[m���&9�v�cK��M:����as��g_���v5<�vئ��v�1�v�sԶN�����l�s��K��'����v^e���1��l:v�e�!�k�r �j���GZHr�$.�M�B,��uم ޮ�ܗ
�.�c8�" �s5(����r��eٝ��6�Om��L�*v"�Oo�F�y�aﭐ!̦'n8�l\;Mk�4p�c�U���;��۸�V+,ٝ��^�KIs0�:��Şq���7Ϗ�Ű��3uРs;]�ӓ������`^/c�Ӽ��}p���#�5YOE�������q�l�gf�vpq�nX�,jL�[���e�ۍqc�eCͷZ9y�����s�m�4E&
2#�����챍ld���q�0����* 3�[Y�&����Rnu!����n�m[�Nrs�������I&���O������#���3���h:���������|y~��߉|�m@      $�
������Z�}�8z��qѶ�b��Ȏ��=�h��Ò歵2�s�9�L;�<h�4�&���f:c4q,e����^�+���1�����6ǧZ1�0�Z��ي��b�K�p�:Y��r��j�����|Pgd�rt�PD�[n˓�ז�9���_�ʢ[M��2ُ{5�e�v �|a��IС�fJT6�\{w\W��U^�ȃ��<��,"�i��}���#��^ϛ?^���!��% Q.��sF3٬w�Eu��6�"�L�1��c=�+m�����v���5����Нm&�9Q�゚�i�<<��N����A�ٍ���l�h�Vc�v��&�$X� A|B�D}�R�U�1�8��,п�n�R�U�ߧLU��_j^XN5.je���3أ݈} @�\Ǫ����3,������=��Q�"���a�3Ͷ�a�gYԞ��zq�ե5ee�%�tX��et��7s����W˘��� A}z�3�!��% P%���  E^kz���~>պ�, �&]<���s}�p��eR�!��"��B z!�{�hLe�	��(&�T=�Te��x׷X�5�d�	Ȕ�sP�X��{���(��d��m�e6%@F��{N��Ø��ո��[6�W�뫮{�����?1��xP����j\ ��dw��;z��f����1^���*��6�uꌼ\k��W������&Ia��� �����XX�	"k�bj	 R��CoMlww�I�'���}�0��,��r	 ���`�	"V��i7�O���$��}绑' s���Wx���[-�����⭱֌B�̠�Lκ��a�b�u9r'����H'���$D����)UD
�e������̡( �J�x� �������cQҢ~�%�A$���`�	"o�bj'�Ts��ل�X�QW�A$M��L�H��|��$
)�Z�J�߱5�O��0I�4w�I����eVi7�N~�LA%Rk}�&��A>��`�	"k��Ȥ�kw��ˬl˕��lI�9���5�Os��H$���i�I�wɂH$�ް��}�6^V\� �    ���v]�6�����sjUVN�<k��n@;Qa�x��>�Ol	\�z�[��佧�<�a�����m������.�C%\mWA�-���� �����x�oU�:��ָ8�-���ri��9�7	�����U���vA9΍v��ka9�����ۀ��>�nW�OA$S�~�A$OwŦA$��&	"�&��ؚ�H&�Ҿ��M2�BH$�����HA=���$D�?~��A?s��|��RD����ϲfw%��M�$���`�	"k}�&��A>罭	 �'�v� �)��{�����A�
����&��	�}�$�H��2	 ~@?���$�H�����YVeJ�&��	���A$Ow֙�O�|�!"0+�� �y\��l6a�̰K�{U҅L�]�l���u��.�����W�������Ȥ�ww�`�	"k}��$�}��	 �&���{1����m9�O�]b���k��N��� ���5�M���$D�~���E7��z��2�Y�JH���w�MA$��`�?����i�I����$D�9���[�2w��A?wقH$����"�	���I|��MA$o�+�*�˙yW�9
�H��֙�"�[�w�H$����g��L@�5� � �ޜ湶�m��R����ݖu�wbcv^k��..i�(�馭��9'޿�	 �&��wI�$�}�f��PI�~��$�{��d������A%Rs��`�	 ��s�I��� �	�	 ����W�(��ʕ�NE$��`�	"s��ȝ����pۜ�[V�-�o�d� x"�m�p���LA$N���E'?x�a*��+3BH���~��$�wwɂH���}�&���`�﵂H$��߼O�������$�o��I|�5�O���$D�~��$�o���Y���p̙d��@���9�WT��	)v�_�ķ��V���w�D�~�PI�9�hI�;�Xjj	 �]�`�	"o���T�%VB����D*	�}����n	"s��$�~��`�	"o��bj	 ��WJ�eT�s/%^��I��� �	��a�H$��}�bj	 �s��H$����=�0������n	'�D�~�}0I�9�}��$�~�s��md`�
q<�&���i�I��ϲ^U�ʆ^U�	 �';�5�zG���A$N��L�H&�}�A$O˾}��@;;\m�u���r�Sb����^���v��̗{NA$�߳�I���A$OD���b�	"s��PI����	UX^]���$Dﾴȕ������I|��MA$�w0O�.�đ(������d��n	 ��~�RA$M���RA?wقH$���i�I����˼lˬ̭/cPI���PI�}���H��֙�?A���`�	"s��'�d��]ޓpI��0I�9�ZdA5[��I�wϾ��A �I�R��������[���     ��i�l�tD\�^0���n5b]<[���tx|F�]r���]��a�4Ҝ˨��mI�Ŝ�%�K�{4�.���ira� ̌%�gilD;a"
�Q�<Ӧ�1ָ��VpEó�-ߤ_}p�4�����~���O7����k���F�\�Pˤ9�ă5�����֖��7u9�����DA5��	 ����&��	�}�$�H��~��3
���+I�$�s�f/Ѩ$����MA$}�`�	"s�ZdA>���/*�L3
2���H���bj	 ���I��� �	���$�H�o��ʢYf\��I�$��}��	 �';�L�H&��`�	"o�}��$�N��ل��/)��	 �'}��E$[�b�	"o�|bj	 �wقH�� �d';�ffeYs*�#��gOj�#vnMJT�\�i+��5�|�?�'<�샭��;j}�9ߋL�H&�N�U�fe]愐I���MC��@��؇(6"��قH$����Ȓ$�j��`�	"o��O�Y������F����ټ^Ơ�%}�q5#!QM�2�I�7�}x��NP�\�_YU&\2�JH$���}i�$�n���$D�>�PI ��k�I���{&aV]���n	 ���X$�Hr<��PI�}�k�I��nD��9;��/J��3D�X��{@M�d��sj�:5��P�%N�NT��f\ЀH�L���I�}�hI�;ZdA5[��I�>��+�2���K��M�$�}�<�PI��L�H&�V	 �&��ؚ�H$�>�3	UXd33JH$��{�MA$Su�V	#����7.ۀ\k��RI*@�T
!#!#!#�'�b������RU�B0����šӪ��BQ89�E��*�0t7Ǚ��:�zw���w;^�d�%0��B	4xܬ�]��ƪXK39��xl�y��HJN%��T��������R��n��y6	����s�)�%X���3:�Z��H�gJrQ��Py4����5\�$T��Sa��m�HJ��,�Qcz�U� 4�.�l�Y�]_"ⓨ_��=N"�bc�O�e�x.�xS���\�k����6�=���t{T�:��=��W�b�>_�]�+QI�>�A$M����cutL���&��	����I|��ZI�O���$���{��2	"������h�*�&����w��PI����$D�~��$�kw��$D���ٙ��6��U$۱���^8s�v8�46�hK�h�X�ܮ�pI�>���$Dﾖ��Mn�0?U�\����ؚ�H�-w�+��Re̼�В	"{��2�Tw}�$�H���bj	 �w�`����z%D��&��&aV]���RE;��0I�TM����D�~�f	 �`^r�ȀH�سAʒXne�	RD�~�PI�}�$�H��֙�1l}%���\`�U�X��*ls|ɂH$����_\�*�2�f��I���*	"w�X�C �z`�	"s}�PI�*~��/�@.��[�1-��)ʒn%�ͤ:K�M��J�:[F�͉ �'��i�I���I|���pI���I�=���cutL�z�$����*Ơ�';ﵤ�I���I��c�3%�bH�]�?OV^4^y�BH$��}�MA9T'�قHȲ/;��A$G[��	 �&��ꗐ��]ޓpL�ȇ��X$�H��9�ND�'.��$�H����E'9ҽf]�W2�BH$��}i�I���I|��MA$��A$N ��V��w��N��ӫu��      ��fX�u��;F=�nضՃ�S�r6ɸ۶����;5�a�C������$�ƥи�\��5K�ݮ˓3̫�f.V��\(�#&|�4B"��k�0��Ca����ֽ��0|o�2�ֵ*rN2O�I$��Eݪ�3�[՘��y�G=6մ���5�?��ci�,���rvNI���H$��wؚ�H'��bH�	"}�ZdD����,ʺ�ʬ�E$M��u�OwقH$��}i�I���q?t$��߾+�EYf\��n	 ���0I�=�Zd�E7��0I�7�߱5�J�Ow'��UVWfU�I�*'�}i�I�/��I[�ؚ�H����hI�6{;'����Y��A9��$�M�o��MA$��0I@(���w"N@����Ϫ����.�۲j���v\ƽ<��u����f\�\���9;�ϰu�OwقH$���i�I���H$�������&]����H'��1zp_��
�nв�!O&)��a�$��ݦE$��s�n�9��&�H�	9Ε��Re̼�В	"}��2) ���b�	"o�}15�O���$D���=�0�.�K�n	"���0I��y��&��	�}�$�H�{֙�O�}�K2���2�&��I���MA$T�}�$�HH�{֙�Mn��$� rNrI��?��UWLe�b��TjP���t�«�re��2���̗{NA$�߳�I���A$[���I{�鉨$�N���0�U�C3�lI�+�2	"����$�H�߾��A>��:l�=���V���D9'o�H$���ؚ�Q��P��(,��{��/
 `���?k�u�$C��z�i�I�,�f^4^y�JH$����~��A=�{ZA$���A$|�LA$Mo�'�/!U�E��7�O���В	!�H/�߭5�W{X$�H���ؚ�H����_�UU�D�lV�I��+Uu�%dk�G,\��<e̼��	 �'�}i�I�/��I{��A$���В9�s�fw%��n	 ���`�	"k}�&��	�}�hI�>�֙��o��fUԘfY4$�H���bj) �ｭ	"�5�}i�I�o��I���z�Qeە+4��H'���hI�>�֙�M��0I�Ck!�AI/�h�^�Vs�5y���	=�O���2�ʼВ	"}�2%Ĩ����f	 �'9��&��	����$�H��ު��333ĬҌ= �FQ�mp�R٭N�$<�ùy�(A~=ߘ$�{��`�	"k}�&��	�����*�A$O~�i�I�l�^4^���9
�H���ؚ�H'���hI�;����H&�y0O�5BH���'ꗐ�t]^�pI����В	"w�0�H&�|�$�H���bj	 ���_YU&Y2�4$�P*'~��"B����`�	"o��PI����$�H����엕Wr�����H'}~�$�H��}��$�}�{ZA$N���A$��	դ���z���{Zڀ      tn�,�ɜ��l��XY�rjJ��i���F���LBTC��n7zL�l�ѻ8�Y1]GP
 U,��j�˃HbF�Vkp�E��eh�Q�Mb�viF#�޴j�{6��]�L;Q�0S����6QS� ,7��ʻ�fffe���ջ Z������}�FpƓ�un�%6SF�[S��H��bj	 �ｭ	 �'}i�I�/��I�}�s(��ʕ��pI��}�/cPI���L�H&�|��TD���PI���x�%Ua�2�BH$�߾�PI�o��*5�r��&��	�}�hI�6{�f9wU�YZM�$�!��H$����MA$����$RDﾴ�$�o�s�/�xVfM�TD��&��	��ƴ$�H��֙�M��0@������|��H;03���)כj�R�g\s˴s]r�raVd��]^�pHA>��kBH$��}i�I�/��I���ؚ�H$�:W�UI�2�4$�H��֙?ѵz�O.�uk3Y��8a�k��>�T4(��q�p�;��
����4Ԡ�6Ud�����n���2�f2�h��f\��sy���62�2a�tN�� �rZ��su�f�Gޘ�n�{9+u]]V�̰\`l�����ڮSJ�+���'E���P��H�=}�C�k���4�\˚s%�^�csu�o5��-8���̧|������㵑�p���V�Ɋ������$�����y!�>�����<��-���_��c׺���vG :{��m��A6&f[D �ؓbp���콋�4)�fK�)ԹBe6U;�>>��>���/9�պ)%��Y���2�^w1�1����$��oouFo)s^�a���퓁�fZ,������/'U�y���΅�N�X��Q�H4�CTJD#P��^�N]^�D���4��.h;ņ=~�6����~��ʪ�E�\q��mt��ZC�e�E8w�s��=��\HLM/;�3����1�1�'����W�f����=sf+��=��L��-9lY9�W��+٬z�\Vd�-�(L�KT8@�\b�5�]���@��{1w�HHp��1��1�����Gt�1����Cl͟vm�f$E73��T��>��t�?w��~����?���<�~���j�$#$d�I# HN9ͳe�6m�l��i���6ٛflֶڙf�5-����3$�,�mC-M�mL�im�NٙJ8�U�-�lSiV�E�SI���[(�d��mJʹF�eV��$�A�D;�@檓jEm�-�����sE&�.x��m*���!��¶�̆ɶ��Ul��U�Rm#m�Ѵ�[lQ��&�Cö䎶�[2jڍ�ڕ�%��%sA[F�lٵ���m��P�f�ckki�sm�m6Y�����LқF���Y�cm��[f�n3�[h�-�m���3ce�.l͆�y�y�61m%��̵�0��)�s�[KlQmRؕm!M���TT�;�� ڒ.��9�QmSb��U6�l�J�2@�%l�u��R��P�6�V�6UUl�R�Ȧ`mAl mJ[
�l���ra"�x]��'g��^����҇��M��;�_=����������T>�O���G�j��������R:~����#�?ė�����G��������T7g��%?�K����O������� @    ���� @ �f�6��P�?����}�U������9�P(�~o�=������s�H�	������j��~�")�L�}ؑ���q�>_㿲����v��o�r~߇�0�� }����>ߋ�0���IOO������O汝�?f����o�ܺ����?���q��?�]��������)/�����מ9�i�{����~��x�Ks.M�%���CjK03-��e�M�l�M���E��)�Tn9)8�[R��M�[�T�U��3T6RmJfJmU�6��)�-��BY�Sh��[*m&�l��ԶM��h�6��LĨm*L�Sj�0�ș��Ve-��1�f&��I3��I�M�fKd6�mB�F�L�6�imH�i�ڬ�)�e3&��3M��e�5�1�26��֑�����mJ��3Hڍ�56[Y�'6����̫jM��Im�+jU�&dM�b�<�6�Ƶfm�cf�j���mk3i��lٛkM�l��ff��ʙ�4-Y6��c�l�V�)/ѩR�Q�!ib�Ԛ��* ��[�@�P��Wa��a�lv�[?���g�RO���).���}�������G�S?���fz�W�t������/�����i")�����S������'���vg�׉���_w��ߓ�g����v����S�|��_���;~$�����ॏ����7�}__�׮���i��/�"��϶H���m��g׻����_N��ھ]���^.��/������Ew�ݭ��m��_���1)ə����.�νy��.���TE�(6��n���n���vyx$E;q���x��~�������a�_��J��������?��N�������s7�����~��+��?W��>~݉O��ύW�����$E<;�������'����?w�>߶}�x���t5����Z�{�|B��?������'��c�[��A3���?�����4W��@��M������c�b���������ߖ��}�7��IO���꺿Q�}�%۷��đ���¿Ç�u��r��Z�1?���k�{S�� �� _��ܑN$�$�@