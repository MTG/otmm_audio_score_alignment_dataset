BZh91AY&SY��	��~_�pp��b� ����ak� (���P ��) U��QP������� 
)*�JI*�)J���@��R �$A@ �B�  (
H�� �@( �� @ 	(��( $Q�   ,
@ �P�(b }��b;�S��0q� {ޔ���K�@�1 � (�}5�3_ )ťQVf�5N iT14���*�P�bk���>�΅SJP�4�f�@8�鯠   �     �R�i@w�_M^^�ܧ����;��� }�>�sK�Ew;��s,t 7R��6>���K,À nH�k�rC.�۾�<|���}�gץ��������U� <
    I�Z ۭ�w���<m+����@/�ܻ��s���'[��0 �㑖��%�� ������ y��GNZ��y>�s}���PL����Ũ��x =�� P  
�� �D�n�qc�.{�C�� ��-�N�{=���g�w� q�Y>sC���y��\�����{���o��=�sn{���� }���d�c�w;����/
�� *�  ( �@|>w`�;W=�/6�5G� �c��ϡ�\×J�ǚF �\��n-���7��u�y��<��r�^����{�s���� Sq�ng��C�|���'��       (D�"jm�R� L   4�D5%J �   �OǪ�J��      D�*��d�F  #  0E?�i��TM d�h�	Th�L	� �b|�����5�����?�o}�u��������� U�����EU��W� **����EU�������������/�_ڿ�o���՜�%	o� ��10��(Mf	�J����<HƄ�)f�탆�6����!�ɓQ$c�ada��2��0�l5!�	��j���S�v8q�D]G��ߧ�L{��'!��`��\��GfY���;4�N���YBje+�1TD�SBw9+�����]�r\�$����`�%	�N�ӻ�rr0�T���#\r<ts��ox���IԛMA�g�
&�(SR*�B�(����tN]�x{�����b�ͻ3�2$��pc��CL�t���h��a<\��):�겸��KX�y3ۋ����Nf's"h���W�JX��҅5G��/o�8U�@Fڿ[w��w�=N��S�g-]ǘW��u\j�U|N�I�P�z5du1d�i�&݌�&�Ɩ"0c'9�Y��19�EELHc�	�9TGR�! �!�R$6��������t�iT�(�S☓�s����\X��fHgz�w�fF���`YYu��㽐A��'K��w�-.��Æ���b�T�M�^���-��9�G]� T�TR� �p�Q)2Ji������+)A$ÔS���:�@\��Jd�Ǣub�FZ������F�4����c�8M9BTF��Mo0� ԝ����X��xw����Pd�Fh{�\��X��-�6]���7��Rq���q�����a��y�p����.זv�Ӊ�|�vt��{k"�y�ɋV�,'Ԋ�$+{�tuѳ���;�5ZW8�y7Yb�S�=��ohq7�&�n�j�ۡ�2&2qr0�7�P�BP�������|��\���f��p�{�V'z��a��v���DѼ'�::����n�,M�{��Y�$螠�N`d94ąJ�e%�r$T���h�6����^_��"�s�Ք�bM!6�&B�m���1�+Yah[�LE=S/�z����ğ0]S��D��E&&�F��bK)���e���JQ�"r2\�ד��s[8zvxz�<'a��%N��!(J��9����;��z���GG���w�g9��]g�e^�¼��n:�r�̓$��:�\��,��zBO�K!��Nbbk,T�:�L�N�:��D�N�:��M�yݗ �V��M�pD��R�Vw+������6��ˮy_x�D����SBj��J��#Οc�9�p��^�ѫi�n��2quJե���P���i�ԝ�w�~�E�;|��c	@h��ƽ�	�L�Xh�:���0���"�������;�]��Kr(���5�S�Y]X�tV�p��HN즔�I����L���wK�N/ 6nC���잨<k�n��3�Q�N��!)�����"���sQ`f�K1c �Y&�!(1��z����d�#��˜#}�0�q�5��7�#�0�A�JO�\ΰ�k,p��hb�m���h�f�5�yb����*Z)QY����Ru�X�Pi��Ɇ�`A�a�N�8��D�����h���L�F�s��}�w� ���.98��5)�)D �(��B]Kj���ga�Z�0��=C2&�2d�LN�)uN��]/vJ�ti�(���}�{����O�ݛ����oI�.���Q}]}V�)�XF�"����G0Po8�b�����+V��H�	)�0JT4����#F�ջl�\�\��
y^?q�",�.!:��C��D��
�P��I��N�۰�X�=��<��<:y��x�F��t���p�o�$�n.�r���ѳ����J�;��r4m���(J	�X�5h��VhJ��#.�C�Ԏ+������	-�$^��;u��Y��P��Y�z6����$�d��h8��4�&8Xhհހ4�٪N��K�켌7�r0�u��uӉ�5�������%�<5�k,���賀��L`�-B�ReO�m,w)u�4�$P�%uT��N�:�x�Ŏ{dw��e�Xoz����]j����Ρ<����n/P�BP�BV�ERU���hzl���W���̌N��w��8�8�����}v:� 0�L�P�׎fN��w	�ֻ9�yv%	I.�ipI�!(���Y�skVD����rfs��9�v���*T�2E	�%	��$ŗ!�%	�u�BU�bu7&`,A(�h�&��N֦S1H�����%:%���nۃBPi��' ��of�Ӂ��L�ĭ`�j�C�g��6	.7R�<��)�s8�y"� �����(O3��d%!�!�`fhJ%�6�`�%�!+N�d'P���-��M����LԹ����Ҵ+ⶴ�'q�l�z����L�A)ZPT�	Ԩ2�B�Q�o֬��]�Z<Ei1:Ma�#�e�u�<<-�8E��Nr�@D�2s,ԇ;ݷ�גl�:��܃��Jz�9�ލ�Ûx����{1F�]�t�tq݆����S��%��r3�0�����Y�,]�̊�vF�I=sRdVfj�P��rp',]]F�b���1qqX�2At�$�bMr�BV!��%	A���`i�9�P�#Uw�J�\@��Jg�-di��S������x�����:�usQ�<��]�}:|�k ��3OQ�kFd8FN.P��m�V�#����ph�
_K:����������u	F8���8vk4�A�&�%�-:6��U�V�\z�F���f���g0<U4���^X�W�pq_.1v���M{�%$��J�/�/'ڔ�M�h�%)�j&��2��Y|\�)����"��%�C��f0͆.�C�;���Y����Ek��S#�3Q�:���Ü��4o��Bo�<�ev�
�]-gr�ֈ�լ��uB���,C��Os6Q#� ��L�BLM$���\M	��ܙVl����d%���i�&A�&��y���U���Qg�ƺ�3�e(*i9J�(�L
t�5.9i5�P��+��9|�(h��\��	؜Hj	�Q佶LHT�;�z2���Hh���$TRq��QT�2\rp'�lJ��pѦ�k��I��S�Q�M"��5w�T��|(�[Rwם�ME_{�ʷ����<  �
5�<�񃆺֎A�@3y|�y\~�5o��Fq(�M!�BB�ct�F�hN�B���X��jR����5��M�e�ֳ�֝ƣt
2��J��v�;üB�|�1N��;�̻�r��1
V4��U��[w	�a�2�X�:�>�7�5�]*.+����5%�MliNR�&�PT��	�eМV� ���ܸ'3˻��ëG��kl����,gN�����d�^`��u�3FN�L���޵��\����}��a�6��Ӛ� �q�'��8@a����`�f	CÆ�|/'Q�9:$�2L�mfLy&V��cw��aQ��mda�c:�Lh�Lc# �Pw�tx���Rbd����0X���uxK�\�,��+��&���U���{�m��'WOg��J��O�xZ��P�����2]>ϫ����L�6�~a��k\
*/��N���yI32�R�IF�j��4�r��3$��J�nHff,n1C�uA�+��b���\��-qs<DK\��ZK���E��|�VRX�	D���YP�.�|<�@{�#��z���
�g��I�:4a�ºN���pa���e����%/�K�y�U0X�e4�!ދAy%�+!P9��Օ��/ ��PT�B�	:�:�00|�i���)��!.F�Ƞ���N�[����Z����YS��
qy,*	��)�����C;B�U�ˬI�[]����Tf��(� 9ޤ�N�ۘ�ηru����Y`Iް45��#A��ƒ�&��M"�"����A��f{��|b��QC{{��`I��V�H5.;��	��7�'Aʅ9R��2	�N�CB`�N(]���Y��#��bB�/_��ଵ�>	Yp�Oc+d�I��rsC�O�(z��49	BX%	LH�J�%�%�c����J�J��ި��)�;�s���X�J�J������HfI���.F�0�
����_���)e5WKc�X�.	��҄g���c�zv�2�=q�*P�M�"6��`�*�R�u�j\rY�r�P�OQ6``�Rd�y	�%	�NBu��{蛀��&N�,0p|��`���j��(��Gr�'�w�p��N�(4EP�'	�J��0KA��V6{�[��A��CZ��-�,M�JSC^|����I�] ����,!����4n�;uW^gk�T�9�be��fBy����$H>90��1NœW�GmB[L!+A��$� ђC��k#-�tnqr4m-Xx9�K�h��eDQy�K��jI�33Td�r�Kֶ�&U�1,I��wA�Jlm4�}J`ja�$g��$��Ԙ�fNUdL�r	��YFp�g`u�Ç^����)�8�ă 1a�S����K��
���:�����O�$ ��9�  |	 �   tHm��Jl   G8  jZ  ���    � @��� p5�H�����8�$   R��)�M� 5r�m�۔����D�a�]� .�P�̮�Ʊ-�ĉ�	9�$dm�cC9n�Z������6�s�mm[$ n�T�]f�2K�q�*��)T͆L+[JHU��N�V�]S���/H��Zj���q3ώPp��S$��L(Ɯa�'u'b���m�ۃ%�h�S$�+j�.�f�m@��m�����cqU�sR�B�1Kv����B�5��i��g��Z�J��%ev����� �pUJ�*���QUt!��LW	'Uk��[:[����jM��p&�U] tn �	������l���O-�)dv���ث�U�[�QfNS5��L���;j+�MY̊n��s��B��am���t�d�8M����
����� ɴ��Ru���qP]�*A�UUW&�H�-�n�#m&�J�V����h�NriX  m���kXm�k�:K���$�   n���k�Ŧ��e o���l횶-�   M�`�C,����AmT�Sg*�b����� m<[,�U4�p�At�Ӷ8~���}�@��$(d})�)�ad  �k��I���GꝽ}�����$l mmh۶�ҁ�$p��t��{һ7U�{v�j�*�=b�'�Ʀ�ڝ9�l�� Cnki	����m� ���� �	 [@-ӥ�u�mA#�m�� �a�[%$�[@?��m�� �lXe�)p��C� ��s[@�  ,16���m o���ձ�m�-����v��UP;J��2Y&*cn��
��S�sd�k��bU��G��  l���k�u  �R嚠A��U@J�mٵՙN` �9��j��)f��m]�l.����K��f�!�trKiz6��Zl�Ep[:m��� �$����]m�� �l��l�N� m�Oi-�z��ڥYV��^N��U$m�0 ��`�i"�^�c�$-�@�!$��`�b��l�C�d�8[@h  �n��  @  ��n ��s�$3N�,۶ -�������	�-���nm[@�    �� [m׮mG  [@ ��  �hl6�  p�V��5��� �MP�P�����|l [I $��H pm  V� �I����ZUBm��^Z�W5��ij���[*U@�i�o��-�� �-�P冓m���hޜ1 rF��m��m����m&�h7d�p�p��8x[���,ge�SINl�հes5�R�W@M���,�*��3)!��V��N�y��mm�ީj��l�ַm�l  ڶSu�Q� � [A,��p������ ��	 m��hm�ö�mFY�HP�U���m�A[n[@�@ݶ��i�PH9#�5��� � 6u�d�[@I�k[% Ƀy�� �    q�-���jI(��;m�ٔxG� 2�6� l ��U�m�p���R   ��$   <�֙$n�m��H�M[��m��k�@�c��k]z♶�   ٶ$8���) >9m ��m���I;K$��`�zMh  8���i5�k�[��N���0!m���5U�J�F���'K�l�ԙ�l  �����$}l�d�b@H�b�6݀3��M�v��L� �۰�f6�6.�[@5�*?f��R�m��n�H5��q Hm�] m����UZ��2.Ҳ���`h� �m��s$��Vm���[vq��m���C����Ӵ�8�ST����5�I:u��kp[Km�����mv�  M����u�-�5�(-�i�]�w���GJ�pO+.�U*�S�z� m[y%�Z�H�#�Im�]�f��ˁ6��T(��,���J��V�)�J���Z�U�s6���ZѶ�z�շ�˃�4����][d�vT��v��8
�-�v��C�l v��&�@k5I��R��#:*U�y�U�H9�����c5��N�u@@m-�6���|���6ۀ�Qm�k$2,�]km  �g� t�$�7fۀ�YͦU/V�.66̴m���Ucl��,��bYd8)�ź���   ,�ۂ�l�%��6�z�[$��ov駡����2I�ڭ�mv¶ v�+�͵Gj��.�E�UZ����cqUy�U�i9|$���G��vV�"�Z�P���=�7sc%�sŰ[�����X
�`�n0�V�U�`z�8���H*U��(ζ%��#�V0�4��n9�w*�U@UJ��d�mp��ڴP    .�mv�F�a������ �sm�vu�I��l9  �l��� �`�� �����m�  �����m��  	�  m���E� $�m��m��Aƽ���� [@$s��5����Y�5����`[B����i�WR����-��D�k�����s� �6��ƻ  h����   �H���"Cm��rD��pմmE4���-����m��l6�d�$A����(�s�6���E��R�]*�R�[.QP�6�   	�m�� @ '@�i�f� pd�_8� ��F��j�m��h n�܀ݶ$ �'+i$�ݮ�Amp��X��l   $�d�f��d�` �cm&ݮ��YmҶ�Ӏ���*U�UP%ڕN

Wefڨ.�e��tT��UU�4+QF��V���@8��` -���&�e�h׮�#n�9���݃i2��ͤ��@X�I)"��e�$ �v��O����k����pԀ6 6���vC)hm̰��6�U.� �;T�-Ү��U*���')�rd2���Uj��eh
�  ��SI�8�� �l�6��g�r.l�lm.�؝�4�5WXt��ݵ�gcC*��.;#�Y5�m����Y����a��Az՜d�8 ��;��V����XЪ[��X$sm�T)���Ъڔܧ��[P"G6�` �-��`h�U�X�; �[i1 ^��� ���lA�]$Κ� �� ����L�5���08m���I�ަ�H���m�m� HԝzԀ   l[@ �h-�	 v�  6�`n��`�@     8m����` �`�K��x����   ��ҍ�l� I��'��U����U��@       0䄍��iv�.��J����5���m- �-�l6�4Y���  p m�m��ӀH$ �e�6� 6Z �-�@ �   !�R�u��A�m�H���R�Hkn �`  ��C��H� l   �hm� [V�  ��m��   �kXm��  [u���m� �m  7n��7Y�kn�i�<�쪎Z���ڸ�e�*�U���
]�ֶ���l��\�h   ��ֲ�D�KU*�UUJ�֓6��r����@D� 7Y*L2 [W�F�-�  l��]��`V^j���V� ۱ �f�i0�%�-��5[Զ�:ڶ��J��AK�T��Iv��l    a&���%�:ۻ[t�m&�ݖC��m6`Ø�����;:Ѷ���rPֈe`6��Z��+��PA�8vey�4�͵U[T�M\l�khڗ���.�H�fU�#M��;/W+c��X�qKTu�=fܥ���A6��vy��2�U,Z�[N l��k^�D�	l ����� ! ��ԫ+W� m�  $     x$�o �m�m��Zn���pڶ�@m�\a�mm�t 9�ņ�l�mְ   @l  m �I��� e�   �iQpp�6Z�m&�n�       vZ  w������`R5��   	�M����Wi���m�� �` m�@�[�D�6�[PT� 5UT�p�   p�[M��m�4�n�ٶ  ��*W����Y�j��c���tR�mPR�N��l�ɀ�I��lr�$k�-� p �``ʃ�ʻUF��U^U��ݛ$��u� 8  �h�    ��6�4���
���_　*�������?��_H��ʬ!
K0��D��S� ��?��T������I*��{8�l��� � �� 1A�ЗB �؏��%$��CB��H�� � �=*��p6 8,�Ѕ�"i�7��7�8�r oh����<@�UFp�:|�"v:�����al{iDLR8���8�@<�x�58���S��� ��b��:�+ھa A �MR�,�� ��"'��] ��;E�S�Tw�G�@�Gj
dM�`GX��OAث���_U�A`� ��p=A��p �TS�]��  a�N�@::A�G�@^z����2(��P^�Da_8v z����h�^��& z*�(&��WVC�x���<} ٠ F�p�d`���(&�(��8�����<QOQ|
@�v�q睫�B�"/|D�S�S���|�!������������?�ӱ_�I$�2�AEC�B���(T��%43%A���
%$HiZV��i8f��uov�{��6_n�����$��h[i��u���m;B���'�'U�u���F��U��1�+�[3&Ӆ�nԂ�͚�r�v��/ke���N��Av�RI�uѵD��5�'m^Xh��y06�vr,3�-�]��,sx��
(����ʛ\p����D�l\�41�fz&D$sl��y-�h8�lշS�oXv\p�um��j��m��N@�x$����s�ZU��kT�n��[���gfv�Z3����x*���fy���AF�b��j-�#m$��i���\]�H&�8%tT�t$Xԑ\l�Ec<��mۃ�[9��W\��^��#��dҽYݸ��u��L�X���h�q�{)U�a�Ъ��1-U�����[ae^�U�(�k��6s6�2ЃRYA+Q9vQ�d������GZ-R���l�Qgd��� �Tڱ�e��iU�6���qқ�F�j�S���A<��(i� ���-���r�YI�L �5���:YV���V&�MGU͜[t��Xh�Ή
��8�>_bH�\`+'s���ckv�Ӟ-6P��'��<g�ѲcQ�������`x)U��۬�5�먖��(,n��Y��^Ҷky�k&����C6p�+h8R�ykju
�"Z#M-դ�Ԓ�ŧ@� �j�NѰ�n;q۴��ѩ�g8��=3�T����Oxc�秚m^{d���m��ْ;u���:{z�y��X�v�ƹm:Vڭ� �Z�
�A�1=2�c;`Tڪ��jJ��VӤ���w�[�j��Hm=+-,�f�P]�Kq��ic��UHu� �N��Bk(ʨL���*mp@�EU]�Ҹ�x�C��jr�A������gkCU������=�:�d�����:�������V��.`.	��
]n�� iV�������I�M��bC�&��l9�e�UUQ���5�X	U㣴��R�邑݆qq��hw5�i�e]�v�m@@T K�ww�����d��@ʄB���5t��6&��@�ڂ��>	�'�k��s7�z֬ը�.��6,��z�yŶ5�`��ەa��k���z��9:v���춓`��88ِ�ݭ�����r�g�^�MVVQ�:��Y۳ �q�ͷImta͓d�J������;bاmɫ�Ql�6��=:�1=��.��+[�
���]�nP��m�s�s �w)�&��q C�R݊����b��\vΪ�gT]��wo{�L<e xE��ݱϝʸ�D%�j��P1�!����՜�n,��vw���y�j�m�J���ն��w-`}ݙ�R�T�I�w�`�o� ｸ��<���hr;�N����ŀw}z`����ـsP�m�۸��ڒ]���� ｸ�>����q`�&+���ݸ�ܖ��ۋ ����9��Xv{^�my�T\��e��mg���3��D����X�cݮ��==����e=��p�q�c�i��>����ŀwg���� s]l��v�Q4�����Œ���I���@�ڛ�޽�9W���U�y�0|жM���"�
Ik ��׀{��X��f��ŀsѶ4�Qq�݂��o ����>����� ��k�5�l�mD���w-�-`����������x��ŀy{ڣ�-���=�uǵ��;���u���N�E�cP�mgQx��8�{Y��
T!G�9���zn�����;��x<���lN��ww	%��9��{ۋ 淋���X�Ɋ�˂�X�%�%�*��=�ʺ���r8S0��.�FĔ�S��eB �Z�i�9��޸r�=�~����qkjՎ������swq`�L����k��{e�Wi�� ����9�^���ŀs��0	UK�R&�V:V�J�J���)?�9��m;`<L�u�}����}`��/.C�+9\Ԗ6)%��m�`������9��X��BG�i�Bl)�l�=�n,���swq`���f�j'm�m���n�w�L����s�ܬ���`�z�u��:�m��0n�Õuߞ��^y�9]��~$p: pQ=�ֻ��^�U��2�N�컶� �}�X����9�^�7w�%IR^��C�9)��W;q�������'ua�s�;�]Um��/>���y:�on�WNݕum&�cM� �ٕ�s�z`�ܩU_q}�+ =%#�u%N��������swr�w�L����k��z�Gi�q�;� ����9�^���ŀs��0|Ѥ��F6Gl������;�n,���s۸�lm�?-V@w`�ـw��X�w۟��ذwצ��!$� G�p�p�q@Ԩ�$\л�`A�C H`X)��Ҍ��j�L?����#Qq�St�,��sA���4X��z�=�8��{jW����-�G9��#��ll�+�ͮ����x}u���[<q+�.��y���
������uv{Z���]�Њv+�1m��nۍ�57'tvϭC��hr��5�^G�J�8z��q�IpnP�׸*�&��6��ι9^z�6�Q�f8��:�wi���v0��@�W2�M��;�&�e�x�T�C��g�+��c�����C���J&L)�ź��{��t�M{ط�QX�,gt{\0{w+ �|��;�nV {��sEn�D�ܻ�v`��,�T�;�۳+ �|��9��D�N鶝Z�� �|��;�nV���s���;�&+Nli��l�[�`}I�*HI{vr��\0{^�;� {v���	S�+m�u�s׺�{^��{o ｸ��ݿ���7jAZ�݈���]7n#�]m�s�9ۮl�r[=v9�[�<lve���뫱�m]�;�Rm�ݎ�{^�{q`��x�h�MW##�	��ʮ����׈Pv�*��+ꨕ,�o�� �f��9�0lm�����aM�m���+ �ou`��0��^��m��ݻ��v˖�%U-�`���k�;�nV {��W�Rci;c�k ��O�zl��߱`��x衮5���qG*PGfEN7Xڸ��[t�{gn�p\Ҽڷ�O�M��nږ�+�v��� ��o �{q`��x��x�Ɋӛj[mƭ���VJ����Ȱ	/b�;��0?j�8���Iww-`��x��f���Kkj��R��˼0��, ��&��wݱ�v�}����� ��q`��x�h�MV�cQ�	n\�;��0���׀k�`���-X���w.��5��v�8a��GG3�n_��{v�'a Ѯu��#V��7��X�7^��ـw|��<�[zҰM�wm4��������}�$E6^��+'Ԑo��]�C;Jۦ��Kذ���׀s�Xm�[����ۍ`J�^���$ٕ�{���}]����y+כ� ��1ZscMKn�,�,�7}��zn�v{^�z��7�g��u�]�;�^۫�6Uݭ��	7���g�:�Ç5wY�\n<�F��#L��9����x}�� ����-Rk-[�&����7g��˥RJ��R�IH{r�0�߱`��x�h�MV�cQ�jK���צ��ŀs�u����lm���%�V��9���zn�ޞ׀w޽0�-�m��ܹ�wq�X=7^�Ok�;�^�7w��(J�$�R���>u|�ݪ�c�49���=^�&z7�ykl��n��3ɋ\�g%�F�5�u��� ��s�G�GM������ �:+�B2�Z���\�;���b)���~|_u�L��g˻���0��2�@�.mrq�]�ԻpU��I�z8��!�.e3�{rܴH�@�`��fL�ܕ��pN^,c��j`S��H��)kn�ch�M/���r��s���=[�[�/r��+�M�ͬms\\(f�p��y���zg�����B��{}�y�swr�z�V���YVӶ6�I[x}���9��X={� =�m����"���%���y�����]7��$fc���o��<���֋w�w-`��x�{o ����9�n, ��&��܍Glcm`=�x�������;�2�z�^k}�eiwp��˖�'vp ��N��T�]l��9ڮ��VC��*v��Wc��+.����\����}��qw^�뛭�j(+�h���_ww�Z�DI�!'BH��?}ϱ{����n/[6ۻd�.;eݷ-,��qx�W=�n.o���戲��w.ܗ��}���n���m.{۸����Y-�Wwpd�+���/�}]�2�}�ex���}��]�)�L)ОѱLp/[��v�ǉ�[^�7[{�����wumٻ������H+w	e˾.��Z^�qx�W7۸�{T)ŭ(�9r�Z^�r}�ƞ�vl�\�k�Ew��"��n؛�2��i��W7۹�/�$��	*��M�`h@�sx}#p�|�؂s}T6���`��;��à����R���@��b!��&�8Gq�L�1f�'��v4Ҥ&p<8�T5qW|'N�`Ŭqt5II2�#Y�[��d�D�fn�Rh���
�7��2��t��DAC���F�N�Lf� :����kY]\V�1 03w�=8 �{D�?  � s�}�
��G����J��A��J-J�&J{׾�� U ���~�\R
�o�}c��G�o7�qJD���~��ԥ)���ÈҔ����pz����������)J����>O򂻶��񹙊�U �]�~��)JN���=JR����)JP��}��R�� �ߎdi����kikKz�Wd��vM�6��\�	�c\��u�8ۭ���nܯM�[��{���ow�}���JS��ߵ�)J���=JR���,�AT���{[d�E�w{ֵ�R����k�~@g%(|��߸=JR�~��)JRw�}��R��+_X�������U �@���}��R���~��)JN���=JR���L�AT���ɚ��ؤ���yy�R��{�)JRw�}��R��<��qJC� �%�
d���$@��}�=��߽��U �Z��d�"��[���R�����pz��$'�=�`����bU\�m�*�|�G��bz[�"���Pgu�n}��>�y�[]��]"˱%/W{��Fmvky�[�����)�y��┥~����)N���qJR��}��R�T����O�r1��5-�̪AT�Ww߾��)Jw��s�R�����pz�����k��l%�@G>֒@�$��PT�w3\��JS��~��);�߾��)J}��8�)C߾���JS���_o�%��ڸG/*�U ��߾�\*�R}��8�)C߾���JS�=��R��R��kr}"j�˻.^*�T����{�qJR��>��R���{�8�I�����JS�E>�I��f�<��b͚�b��]���QCmֹ���M(�闩�7)���F��h��w
@m�ʆ�i����x�q���\�)3�N���{v�u���xǭ��N��N�^�t���z�5To2��X۩ݒ���P�\6���<ݭ�-�q�z}��n誶
��ax��y"�t�9P@&�{dȮ֢��]�#r��ٜeU��e���QŞĳ��Gm�\1&�<���9�]���n�S^u�.h�F ���H��ݎ��1=T����o{��~{���R���{�)JR}�}��R*�_��eR
���L�}.� ��%���s�ԥ)��ÊR��{��pz��;�>�\R���Ͼ��ԥ)�}��(�9ww-eR
�����U©R��}�)JP���}��R���~�ƐU ���(�|��;e�;��\*�)�y��┥�}���)O<��R����~��ԥ){���_n޵X[�;ַ�)JP���}��R���~��)JN��߸=JR����)JRy�|~�2�>���m��N�m��O���M�!c�طOm�8:cc8q���gt�����[��JS�=���)>�߾��)Jw�{���	rR����~��)J~����ۻd��W嬪AT��>��u�Oǈ�C���ߺ��({����)N���S�b��z{�3_��ݺ��˗.�W
�K�~�2�R[�߰z�� 	)�~���rR���~���U �^�G�O�R܊��
;��JR��>��R��~{�)JR}�}��R���߷�)JO{����[�kQ���y����JS�=���)>�߾��)J]���┥�}���-�w�o���?{2�]� ���$��nU�0��v�g��wW<m�pW8����%�����g�)>�߾��)J]���┥�}���)N���R���ϊo�jKm��B��W
�H��ʥJP���}��R���~��)JO>��W
�HߚG>��-��]�R�(}����)Jw�p��h�F �<��S�u'�w���)�{w�ʤHs�m�߂
尸�.k|��)Jw�p┥'�����)K�=�|R���Ͼ��ԥ)�|{����Էnݫ�r�U �AK�߾�\*� � A�{���JR����~��)Jw���*�U ���(� �,�q[�����չ���w����g���V�M�j�&;��ܲ�V�e�x��R
�w���R%(}����)Jw�p��)I����*�T��w����;r+��(��*�)C�}�����~��)JO>��=JR���� �)I��ze�����o7��k��8=JR����8�)I����ZS��ߵ�)J���<*�U#|�|�>�VGd�wr�U ��I����JS�u���)J|��=JPx����P(*tb�h`V�aA�e�8�����H�����)JO<�s=���ky�[�j����R���{�qJR��Ͼ��ԥ)߾�ÊR��}��pz��{�;��~���s�lL�%�2C]�Y�`�#[mG�8ۮ5L�'i�dr��������7h̭�7���(~�����)N���R����~��u)J{�{���U U���k~+��⼹/1W
�
w��pⴥ'�{���)K�=�|P9��y��圎9�}IPUM*Uլ��)JRy��}��R���߷�)�+����߸=JR�}��R�������r�[���U UGw~���(}����)Jw�p�-'���b�H*��oø�����
;��JR��>��R���Ͼ���)JO}���JR��~��)> ��w��hpb��X�n^�����=0c,�:��g|�����H���:�rZ�p�;���[$e�v[�:yd̼]r�'�)[ey��`�Y�Z���-��r��z��9�+��۰���n[Y˸���9��1\k�2<J��e��[::a�W��;Bgk��i�Jp���cC�q˩Y��[Z��IGs�,��8A�����-!���[.�t����w|����Nܜ�Ƿ��}�w;�@nܘ����m˷\�����*�v�;������a�Ӻ#\���p|��rS>�?p┥'�����)K�}�|���Ͼ��ԥ)�x����E\,�Yw-eR
�����U����$�����~��({���R��~��JR}�ә�ֶk[�0ު���R��߾��)JP���}��R���~��)JO���=JR�~؄��Ԉe�L�K��AT�W���z��;�߸qJR�Ͻ��R���߯*�U U���k~+��⼹/8=JR����8�)I�����JR��~��(~����)Jw��լހ��u��g�#ɬ8������](n��Hͷ%�]��n2v�v��j�[�e��ԥ'�����)K�=�|R���Ͼ��ԥ)���ÊR���y}��Y�[��v9x��R
����ė�*�];���04+�Wj����%(~��y��R�����)JO>�︫�R
�� ���(K���]̪@��}���)N���R�ʤI翿~��)J}���\R����=2�v]Ʈ
ݲ�/31W
�K�oز�R$�Ͼ��ԥ)����'� �}����JR��G�W�'z�kZݽ�g�)<�߾��)J{��8�)C�}��JS�����)<��u���ٛ7\���k֫����ݹ���ou�[��ػ�kj7�ٜ';�ٸ����*�����iOs�~��(}����)Jw��p┥'�{���)K�������f͙f�[��(}����� $2S��~��)JO}���JS��ߵ�"��n��}� ����y��U S�����)<�߾��!��}DvrS3�}�)JP������R���s�f%��I-\	-eR
�����*�T����ߵ�)J|��=JR����8�U ��/?�nՄ��ڷ/p�AI�y��┥�}���)N���R����~��ԥ)�ѯ��i����ʕ�k�b7hE�kۏm6��ힶ�u������%�qB;-��%�ʤH}���ԥ)���ÊR��{��pz���ǟ}A��T��D���]��C�y���)Jw��p┥'�����)K�=�|R���Ͼ��ԥ)}�Gگ���7�f��[8�)I�����JR��~��(~����)Jw��p┥'}�g�Zٛ�Ѭ�[��=JR��{���)C��}��JS�����0dII!2�A$AHBĒI�R��8�(��$���	S��0�$Y��c3�����p�AT�=�B�K�F�v����(}����)Jw��p┥'�����)Os�~��);��߳Fl��Ї:��m��v*�ln�v�p��N���
�`�*ҥ�g�w��6�m�V�z�-��=JR����8�)I�����JS��ߵ���.JP���߸=JR�~�?s1�Yn�����U �AK�o�b��R�)�{��qJR��~���R��l�Ͼ���������i�۶&�z��=�=�\R���Ͼ��ԇ�P�)O?}���)=�����)O|�m����w �s*�U U���W%)N���R����~��ԥ��9ǳ�r���8�p����D�%RW{]�8=JR����8�)Iן{��JS��ߵ�)J;�߸=JR�:��CB��$��ce0`I�J@� v2���|��@V�,5YS�A��Y!�:�����0�
t2�@5�50�C$RB�$�JRPK M!�٦hXjC�vq��6��L2B@H@�Qֵke<T�]bA��H:�-�B'@�B���.�NX�'���&Y	��F6��ѣq�hJ"-��	`u�*J�P*
��'1�FV�a��bHH
!�Y�0��d�FKmC�CQ�L���I����+Ю���鑂�X���g��-w�nJ��(F���]u��Qv��C��3GɊ'T�������DH�7 :)m�޴u؝A3��2l62�TO8�ޘ ���I	<D�}�y��a����� �	J�bI
�d7�	�p�����!�`�!�  �@��fBB	V�	�R돽'�q
Y�%e�����I#�f.� � �fdJ���%�V�40��� 3(�/�jT�&�WBE(R�k��j�F�{�k3G[dp�Z�8ԡ�
��n#N�
Vێ{2��kt�m�W�|29Syv�Y:ys� �qՁJ��hN�ʛ	����t�������s�ts���:0���1�:��;��aC����-b��jBn���᪐U�5H��m�/��u�����s��9���C%��8��]�ݮH�vn]���l;;��v��9����j��u* ^�=�H��j�x.�휠��>����$��G���«�q�U۝β�hq�(lTjjڭ[J��;mmra%��vU��U�54�ZZ�68���+�]�ڨ�'��l��Bl9�Qg�]�yƬ������}u�[����Mhth�������3J�G=�PAv�q��5�Z�b�U%C����!�RvB�c5$��q-H��䪈�
ӑd)�D&Qjl�nA�f��/l��K���+��-����	[[E8ď96+�~_7�{eO���za��nѱlt���&Ark�hk�G\�4��dN�5u:�unB��mp�5*������΃�������v�3ݙ��P��n�n�@{(�U�J�i�Lh�,�Լ�2��;��K�i�[5��9����f��������D"a�2�-#�i%�mJD�ʡo �����T�jIh�F\���"�+��g��;H�8�^���$4u͋��h˷�6�y �K�6��^4�8���=[m/E�Ƶ�n��d%#���ͧ����lʕ{a��e�V$�֙��Ҭ��Ytf��lj�L�X�4�`�۵�jN�Y�]B�UQ�Tvn!V�hܧL���6���l�[��6 悽�\S+ܛ�cv������W�9.pݶ'��ޛ���n�h"���ׯ[�n���8�I2u�֖��;��n1��q��{Q'6���d�����V���wne�۶���!�8�����P���m&h��Bz��l������|Ⲃ��K�#q= !p<9��d@� *�>������D��z z
�z�v���;E�C�"�y�j�^׻�v�[����(kj��W�h�7'uK;::/6"�u_��*R�	Xovl�dnN����.����^4����z���G:��[��:ƙHk�)'o=�g1cM�cm�-�Un���w�+��Ѭ�qūuuI�;
8�ҝ����/a�k�S�N� ')��d �W�'%�1����r�J�2��EP�<kp��c�x�ۧDYP��ۭ����w����ƷmqoJmt%y�.��˻u�aJ7�=;n6+�j��M���MH�H�W$�]�_��U �����=JR����)JP�߾���R��6eg�P}��=���I�J�����)J^�����@g%({���R�����ÊR��}�pz��.�>i����mh.9w�H*�*�����)Jw��p��$���~��)O x���AȄs��z��t	��o�ַ�R�����ÊR��}�pz��=�=�\R����=��ԥ)�$��W$���\��H*�R��߱W%)Os�~��(}��~��)Jw��bʤH)n�>�Dn/���ݐ�ot�!��PQ�lY���3%ɗAO���.{r��ੰ��r\���U �Z��L�AT�V��2��UAٳ+ ���p�Ek�;�-Yn�.������IKM$��j�0�BI-+�� vu���w��<n�^�=�D$8�p���iD��������?e`�����/ ��H��`�]��ڶ[�Xg�r���s�1}���y������8��Cj�/�o�W�^ Uiݑ�͙Xf�� �o۸*V��ݍYcb&cq1�� 3��Q��u�m�t<��D<���t�j�˷uv��&�����;6v:�1��"9G�5�g����Z��n��;˼��;6eeP���W�^�����DңHW������n���݁������8*�b��Ձ�ɕ�w��������i�|�~��/g��"��� �ٕ��f��;��$�v[��K��y��0J��_��������V��,�QN�ht�U�����gcR��s�ɬ���u;��vn�
j��C��j��M��c��2�M����/ �����dV��lwv[-۬��9�5{e�]ݏ�vl��z%%�6��aV�� �헀ywv> vlx=6s�&�*]�����T����'��X��t��v���a�fbA��ԛv�D(�V���|Б�PH�������_ ;6<��9�5{e���e�	6�s���z`���[�̔��t{v�m�n�Β�vK�ݫ�O��.�]���C	ʩU���9ݓ�W�^�_�]p�c�'��#�vڰ�ݻC��ݽ� ��/�ݏ �vNp�Ek�;��1�촛X}~�| ��xvI�ݽ� ڞ�D�ݻ�V���|y���ǀ_���d�]>����	�
TO*���i)���cw`lDy��`{'몮�������+uZ3?���������Ǎ��]�+f'm�l��g�����I]hݗPWi�.�ӫc�F�Q�7CM�z�V���6޹�Z�8eK���Di19PU�=�=J8;�E5�6Rv�<PK�R�˨�9��AH��I��@��� +ά]��ז��6-:���9�v���<p�t��25R�R��6���nf��zV���m�7||�3���mD�r�m��!.��I%K)zs��\�bk�[�]�vq.��ݴ�÷o=K��e��F�D��N�7��
�PU!!T����l�]�8��َ�""���݀x֠�������#���@�N77�H3�@��۰>����j"�,M�o/��ǀw[w`}�mtd�s`>d�&虒eL�N��xvI��\� ���|�{c�'��#n݅���4�8}r,�^�} ���쓜�^��V�m3���s���m��Jn^�n��%�<\�F��^�[�K�-�(���N�| ��<�$� �E�mOm"�]��r�9e��' =ﾼ�HEP*�IDrh>�n�z[]�O���s���v5J�"���&�L�t��n��������/�� ���c��$;UUv�-���nl�n���w� ��6f�&R�T�*�]�8�����;�Np��X��m�]ҥ��Ɲ��wf:ǹ���d���l�nq��n�荍�K16���H�6P�x�_ =��6���Kk�{'��%!7D̓*fiT�UW@�w{��9�D$y�����߯�ݏ ��F�E��ۺi�p�Ȱv�%�ϻvm�x�$� ������Li�M�ݿI| �lx�<wa��^�z������S"���a�y| �lx{6s�v^ŀ{��' �IR�>_6�I���,#n�m���7)��5�r]������`;���獸�ڰN��"�aR�X����8�@����� ��䤱�m$�tX�� 콋 �o�_ 7��͜�$TT�wWiSM�m`��e�}������{ s�	ZE����]���s���=���c۰>s�t>�v9�r�]/v�����w�_ ��l{��v��Ii��o 罳��l�����}��Ȉ��&�@�D�4�������#���Z�:'ms�8��tH��qٱ��i1�^��U���,jݱ[�@��?^�������{�9�ڸ5eZcM���]ݏ�� 罳� ���	S�H��ҲݧV뉼| ����l����s�ĵc��-׵`g�	9 *H��M
��7}��/l��M������RX趒C����"���8��V ���g�݁|����Dg�>4�4='9�v��Efs��d�n�s��!c���9눦�u�8)�[n�d�t"�\$hB#�#���m�N(�@��'g�|�.�c��.�v���A4x��v��:h ք�Ƚ]�lmCϗsF��7�Q)��um:6�jDSj�r�K�Y:�W��{iN� V��J9�-r�P����s��	0�d�.��#7P�0`%n�j����+f��1��#[vb�׻�s��A�<�+;�k��{;��v�n:�`���^g�˸$���$:#zf� ��{V ���g�݀ױ�@�uy	-"�cV��1�{c�7}����z����q#a�FꪕRL���I��	6~� ����8����H���Z������6��<���M� ���Cc��{��� ��)*�n�w�l���G�I�s��:���(�eA�cd	���GS�րқ�=/v0��l�uϜO\����N+�՛J�v�[�o3:����l������&p�FE�'t4�������B�O9Ȏ8��c�t�o� �xf�%��ChHwB��8�lx&ɜ*��x�'8�)�i�T�E2� �d� w�<zI�T{��ըH�i;*�f> w� W��L�^�x[�>m������Y3��:�zl�<��i�l`^�](n�SRz̓���~q��;���g��T��IT�t�ݻ��s��n�#�U]@{g�l��~v��v;n���:����d| �x��� �+j�2�Li����-� ;�l��)��߲,ZL���8YG'�u)��C�4wuR�	0�p�����S�B�48�r!�u�S�';�Tt#���&+"N�MJM"R��8>�^���@�@�4����B��`"k��6�.*bv��8�EY�۰�hu�Ґ��  �� Bҁ�4��
�
&�`��b�8NÞ
 `�v��xoh�D;z@U��u�|�޺����ʽ7ґQ��WcN�8�c�}#�$�9�=�ذ����bRƕ]ӻ�һo �I��^ŀE$��� �UJ�/����uզ��wm]�S�)m�ǯ8	��:����\�v���8N9{����)!؋o�v��E�G��G�M�s��P����i���-�> w�<l��޽� �l�U��
��� ;�6I���%����Հ�%!˚SR)SUQIU7�I$� ��b�"�G���]� �ר��VӰ�ݻ��� ��b�"�����t�w`k�;1)O��������ɰm��.k�4��3n����Tہzڭ�B ����e*)ML��X���w�<M��pz�,վ����
�i;�y���ǀI�s�wױ`M���Ju�]ӻ�Ҷ�&���^ŀE7c�}���UB�&ӡ!ݫ��8wױ`M���lx��� ��i؆�>N��"y���@����7sv�zq���G9B��Ь�?�1�B.F d�LBDL�B]b���1HJ�$j�)��+� ���.�]�`2D�v���r5Oc\�8(j��a�OW;�����3���t#[W��v�x��vz�8�RM�x�C,hF��ڜ�|D<q�G��qtqM�@�h�h�gZy�:����B�q��W=���&��$s�;ts��#X]��n�q���,.�n�HQ	�D�@6�-�CyK���]�єY�eE�������#�l�7Q��=<ɑ�v�b��!�e�}��x�?6N]s���n�ss���0:���z��Oi������[sGwݫ&5��:u�uv�^ ��u��w`{Ӎt�c�+m"\�v�V�M&��$���}��{ױ`M���lx�=��le�j�UJ�*��d�] o1���G"8 �n�@~{�`}�ȩh�IQJjII����8�H����^��X��� ��՗N��7��� >��ɜ޽� ꛱��Je��&|�5њ�,`�.�a�ƃ��݃۵m��z�|�m�H�H۶X�,�KnK�{�}��^ŀuM����}#�=ت��i�hl�.�ޛ�Ƶ%\��_���%�����ܫ {��}�݀}��J��!������� ;� �����X�t�Rؒ��Y�>i/l��d� �FG���׭#n7v�v���m�ݓ�޽� ;7fp���J7��@�Rwt؝�{�����ue��4=GQ�q,s�u�����'�s��Qn��Xݻ��� ��b��ٜ �<{�s�{��Բ�J�V� vn��}��ݓ����>k�h	L�V:�h|�o3�� �������H),���
� B��)ا�:�޾�r��7fp�i)I�]�WV�v���9�=�ذ�vg ���G�{�UEr�v�5i�p/l� ��7fp���ݓ��n�"ꥵv�V6![�W��<86����uf���Q��!�W�\��gەӲ�M4|���f�� w�<{�^���@��J!=IID��Q=K���}��ݓ���/ ;7fp	[iP��V�jձ�m�{�s��ǁAٻ3�� ��֨�[n��wSWa��Q��g��������DD/$C��s�{�-��mHݖ��Gwxٻ3�Q�H�����헀v��d��\���f;��ۃ��	�	~�)/K:%�Ū�-��r3��f 1Y-BԖ��ɮ��>�u�3�n�/c��A��X $�l�3R�&�����7vs�w��7c�}����TW-6�BWi�� w��7c�}��ݓ� ���Wr���i��v�USv> w���9�*���c�<����ĕ�V�*�<| �<����������]�������&�@�%Uu�߯�߮/H��ky�ўS��:��!�m:�`�Z.1�nk��ufݮc-v���e㶑����[K�Ql�xwg�]Z�ٹ�������������K2.��ꌻlZ�N����ywԹ�:��⛘���Q; (0�W�[��ʊcQ�>�rv�8h8��t��2�)�/Z&�杩�3�+ъ�uv�N8S�<9Ua�%�ծ���~w�|�����:7>�|�L��;�jJF���s��oW�nf0���i�2�j�hB�m*�8�<�$�Ej��;o �����:����� ;� ���%	�wH�ӻ���������!���`ǵ�3�n��G"��5�5Wi1�vX���n���c�7�'8W�^�ٴ�[�-�cx��U��ǀovNp�l���"#��[ڰ@I��IP�J��J��{�s�u{e�f�� w�<��7�@�8�izq�q.�[{{kc��o���f�hۨ�r�/I\��gߎ���{�}H'[5���^�xٻ3��ǟ}U@ovNp�_�]�vZ)���ۼ �ݙ�Q���7�����U�~��]U�y���@ywKE-���V�*�Kg ;� ϱ��R�ǳ�<����JP&�eڵlv����W��d� ����:��|ꯎ�c�=��(�MۺE���wW`|��z�#ӭ�|�{]>����[�) N��r�i��dP�v��K�K�i&1Ý9�cG]�ў�)�ޮ�W�'�Ljݖ&� ꛱��������헀mvm�j�1ն&s���c���{�s�u{e�Sv>UPo�.��'m��i6���9�:������� X�d��\=�7�߱��#�=ت����RT]Ym�pDG���|�1Հ}�u�؈�D'���n����R��TEL����u`E|w���9�:���	���?�;-�*�:Z����nݻ��pNM�K�n��u�Da���VK#�M˻�PǗ���c�7�'8W�^�7c��ҡIe�.��i��{�s����}H�׳�<��� ���{00N�USS�n�|�^�xTݏ��@w���9�;�fRwJ�cMڱ7xSw��Uߞ��U�~��]WB�$F�)(QzÁ���
>^k�k�zw��S�n��ݦs���c�?}��߀�ǳ�>O1Ձ�jJ&E���;����wR=܇�k�8�;�z���W<c�i]�N���um&��7�Np�l��n��W ;� �b�6Sc��T]]�o���/>��)� ;폠^6��"9	��:�%(�T��������`{t#���v���|�ElbV����Y�����/l�������sЎDY�u`<��M8�eڶƚN��9�g8W�^�پ���߷ʾ^����I��v}��`����<��

@��LJ���^y] ����(�S�ϙ�v�¹ћ�߆�7��f �5�����{��E 8�4	BEH1��q�I�:�c��F6��4���|N��_0�'N�M���	�AIC0C��GZ#�xse�Ý�Y�v7�h�r�P�� oH��XY�6J6LH�X�H�;1lA�S�^$)�IT湬Sc&�Ҟ	!*���y�� ����I�rB��)��F���(h�Ԡ�� hĪI<�ӷF�2\��^�t?#��C[E�@�tS^���l-nY>-��9�&��㦠���ذ�h��'Mj��W��c]pnl4��7;���3�A��
��
��"�ҡ[kH�nn��[*���ɶg<��w���ӯu��RGI۶�d����u�kű��؈�.��V$B�ˬuu�'��/3����l�{C5��6UK�gm��5��]��h]l���K<�UU��F�m�(mW,=]a�vd ۪��Qv�vۅ2QӨ��q�55mT��k\��f��Z� ����rҮ��s���<��^R�B���)ۻҭ�-�8�c�0n�r���&�"i�6y[�ɉ�P4�,��ԸҀ8�����c%W���j��*�9�/T�U�[d�̪���+U��v�� �Ip� �K]+�˴��EP�92d�TO�|�Avl����t���e2�vqGR5�<�ON�)3P�<�ZnJ�۞N��Ԧ�8q.�Ǯl�v���ͫ��6:^�1q+B��kK���gcm����J��B)n'=V�l�v-�)�mnwc�="#�]���=Xp�f��Yٖ��[r´��,�ݧ�����ud��۠\x��M*�UI�XX%���ń��x�ډI�[c��m�8'E�\ԘjW�yJM�02�fF9�6A��u7��7�`���r�ڎ��h�f��P�m�zӵk;��Rg6]��`WC��Tpe��A4�j�����Y��	`�$�i��*ۮI��abŜ��δ6���d �bK�UR�e�Gli��$�@3���X�h�G�TRƷ�����k���ZlѶ�&�n㹕jb�TɹM��-��!�Y�'���� �.��^���rr��.\n��a��%�9]�L���t���\��8���;8ps�B *�UX²!mU,�bv��[Dhep ���vWf�6�*�5� 誣,����[<��#����� J��Q��w{����ww���wA笄>�Рp^��@lS�N!��'����b�;5ѭ̳�x�qT��0����r���Zn��],E���6���؞�	F������9�m�x�u���W���Nۈ[J;m�����7�F��;\<�&��9�sm�n��iY�ۜs@>�ۉ6�n�[��L6�1�q�nZ1���z7mնV�r`n�v��t���5�Rvah.WfPl�9AXA\YEy'dUY&ݖV��:y�K?Y��N��pa��i ���|f�W�6.3�wD�;��E�`B,,-+t[v�����"�/ ��l| �<{6s�{�2��ZCnՉ��<��> w���9�:����IA)�n�ll�����}#�7�g8�{�=�����V]:��m�ٳ���� ����H�O*���
���o�ޜk�y<�V�����6��؎s�ٿ�םr밴�0���Ѷ��M�ΒU],_�I	%���vW��W���'x��`b����7]>m��9��z���XR��[m:�b����G����9P�"���$��������]��:���$k%@�v%Q2���IUUt��݁�N5�<�1Հ}��7��8vݪ��ڻ|�~[�~X�'���c�9�Np���wV�ƭ�i6�-ݏ�_�T.�c�;�Np��,��C�4(��%�Y	v�U�����auv�v���ӍM'-4�u^gHM3���}��X��]�vޜky�A���`<�ځ-�)*�TM%UU�/w`wױ`[� ;�(O*���t2'�|��ߞ绿_RQR),��D/�.�c�������B����QS*M.��8,M�� �=��x�� �b�;K�,�+ln��Y���lx6I��^ŀyn�|��f��P�M���"@�}�\�;l/k��=��
��c[���N�����=���Qn�*j���݁���Y���>�:�hjR�m*��ڻ|���X�����n��8��T�TR��R�]oj�>�:��#���wn�����	]��2�t�V�Ms�������vޜk�DLp��\�À����z:�>�������/�cI�N���x6l� �b�<����>�:��CǻS\AQP��TR.�1�[gA��P�m�VSZ3زq=��;Z7rl�g�d��<�v9bR7%�@�Ͽ<�}�����l�� H��Wr�Wi1�"���<����"9Ȉ��Bc��=���;�ذR�-
J�[�Y�V���@�x��s����Y�u`=-RR]�b��Ӷ���l���^ŀyo�>UTw�&��)]�T�ݵm�wױ`[폀�ǀsf��u^IR�QJ�*��Yd� �-�R\�x�;v��������[�Is/�c�Iצ�c����X����z��7Nŵ<�<����,�D j� @#�	��d7X�`q�#ֶ:@�x[�(�F�F���G���E��lܜ���$ʚ�G�m�.Mnj�9^-��\˰�6k@��n��j�G@�glQ)E	m�m�v�VEѻ8�8Vz���r]-K����(QN"[��s�7e٢�y�:8���@���lZ �6�:ڴ� "�Z����ݼ��߯�{tǎ��s��d�]c7Ch�j(���U�j�� �����BG�^݁엫��c휈�p3��I�����x6l� �����|�����߯ ����H9M6ۙ�%T���`�c���c��={v ��L���rY$.K���~� �*��߯ �͜���X��%*Q�Wbvch��������z�����U�ˎ�wj�W�v��羫&O(V�ZI�bǏ��ǀof�p�q���r���ڰ5��ݪ���-\��]�߷�s��_.U*IJ�l���Zx�X��]ӑȄ�[	Ucwc���<�~��{c��ǀs�o���U����ۄ��I|yOl| �<�6s�u{e��%�)-Y$w-�\�� w�������$�����=��{=���}��B��8��׍�cݼ8����n���9/(N�nf��۞H�����cJ˧V�m��$� ����n�Ͼ�}#�=�n�GM���@��]��k��DG���}ď=ڻA��ۿ�#�"n�!mR���J%R+z�r�߾��:��߾�.��C�<V�����n{���ذ���%%m������lcu�/w`{'�lr8�[{V�)-ښ���)�������n��q��噎��n�n�����V%��6�2lj�{��46�1�Wc.&�t��uqە��m�V�����{ob�<�v> wv<�9�Np��Ȩ�ɔ��J��M�3^�9ă��t��݁�e3��pA�p�5*fݴ�� ='�sd���p�<�v>�PJ���V]:��m��'9W~���Uy��Ϋ��b(v���7#�;=�T�cI�����p�`=����c��xۻȌ�!�0+GHp�y�#������iNkc6q�݂�KZ��w��I,��v�~m����~��ݏ ��9U�:�e����$�[v�WF%����ǀsd��[�z�f:��r"8��F�)n�UUH�SQSIT�t��݁��s�b"��ڰl��	45)I:cwm]�p�ꏗ��@���V���Cy����߬8�D�&R��TI5S�<�1Ձ������{]绷`|����A8��?>Y��)my..r���r�l�֫�/�Wm���3����`��ⷎWt1��s���]�D�3��[Uے$ԡ����*ս���;]��V��c�5j2V�Z��И��#�z;<��G-ƻr�s�/1Y�&�����S���.�x���T��0��1l� �a���5��x!eLn�*y�X����W0:)T�h͚�����E�n����_b#������K{uĄp�B�����%����\�m\s���,��7n��/m[9�����31�ޟ�͒s�un�Ϫ��������TϭXҲ�մ���sd��wc�<�v> wv<����6�l����`�f����]�3X��{V�wn�!���T������*��W@�������l������ǀv��)[�e��ř��ݏ ��9��ǀyn�|fӥuITV��e��oW��WQɃgv���U��!rWh��u��ٵy�QcB̷v����x6I� }��yfc��DD|��{]u�KS��Av]�nK� ;��璮	+$q@�)�	����r:�1Հ}��@�m��G� �w�"i������I�����}G6l� ;���	��;E�v�sc�stǎ���]�X�=����$RRU(��Jj��^<w`lr!y�|T��������>5YiYu*ݽ8��;���1���nS�L%��Z�Nx�a���L̉v[wu$NK� ww��<����wc�9�g8�R�cMڻ�v��o ��l|>���ٳ� ��x!~�."R�j�7Hř��ݏ�߽���@�tHQE!K0�,PR�E����<:@�D͆I�����'[
�'�z�M��$x�֗Aͷ��ζ𓨌���Va���P1p_P�S zQAOp�@P�0Ժs��6cr&�:J)�K�	��,^���s�@u�M�	1b-�Bzk�lv�mr4�jhDo�hd!@�+I��F�`�)S	D����#�G�כ��N��qC��$	J+$}P�t>��t=�oX�x ;�b����"��6(�{۵A=���;��<�� �Z���ݴ���Ut7����׷`y7��<����>ݏ � D����Ccv�o��v_@��!s�k�7��/;�2#1Ľ����=q���y۶財m�H'��-ۍ[=��lu�$nE��7�i���c�wc�9�g>��un��;�A Uۧh�i��c�| ��x6l� �ݗ��l�Po�%:��Whum+m�ٳ� ��x����wc�=��uDli7��wo����x�{�:���~�+ �@�@��Tﯪ��������b�Jm�7wwMZj� ��fp���ٳ��v^��������_o^�d+dY
=nn��-u��m�<6�%́�M)�i۶Q����"c19q7M:1,�΀zO� �͜�[�����&���6��blv�M��6s�}Aջ/ =�ٜ ��x�%t�6Rm+|��ذ[폇�U���I���@m:��ؚi���R�o9	�ǵ`ok�[x���r9��ŀwv�ev��.�j�1�> wu�@�G9�u���/W@Ş�V�Q���߯�߇Z.K-�N{hW4��u�q�+u|N���rb�w/,n�B�"�:;l(c9v˓m���v��R��k;=���*��],��
irl��gy.w%7)�na�Y� �܏ta�u5vzn���2k�-�^7X�v�i�v�-�kF,����;�V���[��r��S��lc]S�&M�k�i���W���%ҫ���������~s�{�����\s��K�;Y��Qùzy�[��_V���Ev�n7w$,��&(j��KA�)�[]�um&��'��� �헀j�l| ���J���64���������b�c���|�������۽���(�"!��6*���R�T�S5=��j�>x릥��۰ǳ������6ԩ���]�j��DGk���;�5{e��� �-Edmݖ�����l� ����[��[폀�<x=*�(B;��5m��U"�]cs�6�����mǉ��\�vM��v;s�!u�j��bcM�jݗ�E���ٱ��g8v��uWbi����o����쏚b�A�h�:Qu\{7vs�j���;6�T�E�v����͏ ��9�ꪠ�헀E������lUwIմ�o���{���=���{X� �㮁�sFƓZ�Z�|������ ;6<vl� 7�[�:�
�T�R��뛶烶�C�ݴGc�������xyɁP�m�n�N���c�fǀ?�;�9/c��xO�	hh�Jh�X�1��c�9&�p^�x�����t�B�j�[����l� �헇��,չ���c�6hjW*�e&�bm&��>�^�x����͏ �9�7�N�2�M46"ۼV�c�fǀN͜�����RUIn���
5����˔^;ݎ���cu۲&�]�hM�ky��}�#���I�I���wo-�>�{���	ٳ�W�^�c���)t2�C�i6�>x�����@k=��玻�Ȏ$fƹ�[TRU\�	I3W`5�g�5��\>��͏ ��9�	�J%7M�e]�Bwn�<�߶> vlx�����~����~�(�j>Z��5ʾ���V�D[I�i�X�1��c���ꝛ3�j���"�l|��ZJ��NwUwH����И9�m�O��ݨ�4���w�v��h�����))����IMU��׷`b�9�g���G ��s�k��X4���*�i��7���/ �}���~����s����J�_~�S$�rJSǵ`fM��˰5f9�<���6�[m]�[�| ���g8���U|E�����)K����[I�x��� n�x[폀�<D��[���\Q�Ev�����Zn�ĺR�ʔ��t^�A[����:)��'I�1g:tLƺ��zq��9p��e6퇞�m���n8�M��U��y���Yj�[h���up+�+�e���Б�ٶGn�e�b���^��%��3���ڻ�U� �]��J9G���Icd�����ٝۂ`%YA;d��Ӣ����/q��m�&�sW(�mB�����{��~��Sx�뎔ꥃy�[gv����{v�q.�g�d�{g�4���&��{�G��,lm��$˷� �lx[폀�;6s�V�Jn����i!ݻ�"�l| ���	ٳ� �ly���A�Y�I~?$�ۦ��3 =�~x��vjCǵ�5<{Va(C�E%4Tҩ��Ut6#��8���������� ;6<f��r�l�i�&4�8�l�-���͏ ��9�$.X����==�6�ș��p��v�lq6��[����j�a,����X�wL�]��� �}���c�'f�p}���A%ZN�m�ۻ|����#����յ���|ד� �G�E�������N���x��� o�<?}�%��ڰk�����@ꢪ�J�&j�6#���r!<{]Sǵ`<u�'f�pj�.S`��;�;�x[�u`ls���8��k�o���{t/-�4���	�i��Q.��ˠ���C՘�����;Aˋ��^w=�������"t�<| ���	ٳ�W�^�c���ZQ�]��Ӷ�m��g8UW�T�c�"�l| �����ԮQv�e�o� �lx[폃����0 �!u�@4 ���vˡV@�dbJ��*	���	��&#� ��BU�*"~S�}u����9��s�o�4u)���m5J�x�!l�{V�{]��݁���|� ��[m[n�-�> vlx꯾��DDDDo��~�{=��:�;ϳ���m�����c����k�\j��H�m�.�ͭ�g�6�{a���8�*��?{���zY�u�r,玺�)|F��T�2��j���$E~�V��]����#�	������XӤ;�x�6~| ��W�UUD����v^�Gv��!'Nݤ�X���G�N͜��e�{�Uk
��$����*��=�_ ���ѹ�%�v;i+o ��9�5n��"�l| ��%j*�%v������MSL��8�����j�gF9��p�m��o��� ��[֓o�V�-����}�UP�g8����b�m��m��c�d� ��9�5n�ʯ��;6���i����7���#�'f�p[���� ���RP����[I�WCx������zY�ua�\�B���@�o�����%�&j�Y�zY�u`cu����|����Nr�.�3U�	�ۂ������I�x�Sx�C�O{l�w�y���a�`ɍ(�<�4&��Z�3N����>Br0�͋�b�	��`$#�����[3��Z̵f�+���*hW�e43�g�0�;�� �1�E7PŊDBP�%�3E5@RKG�X�dfi"
Z,j��gZz�j�RP�`a5x���$9�����d��0΁��b�J8$�M:J&�T�ȅ�wn�-��n�e�� M����������.�n��f��N�f( ���e�ۍ���H�m�5`茔�����y�ge�cp���V�\���|Z;Q 6ݕ�b��:j����v*���-@h��.�J��kC*��^�p��Z�v���i�2��#n��7݅5���r�e��d�k����g���a�R;E�k�z�;l�۩�U,��v8F���g&�΋�AXX4pl˳Gr��@�%ph��ί�H��bc�m)+��:ZSL�ƺ6��|�=��-�J�k���/U�7i�Dûv�9�4�V�m�D���⒝g��笵r��F�!�Nń
ܡ����\�Tڍ
ʦ2�
��V��% �V��e(��$�\J���j�	"	�*��S#(���36���нE6^�2���v�n�&�j�T���ȼ�Ɗ���eV�l��4k�ye97��sv���4es���Gg��
Ռ��U�ZV�f�,l&�v��N�akT�]I�N6�,�'{]f���zw��ӌ�v�WE��<��t�Z�ٜ� ��Bc,irų�
NȁU����viCtJé6�;�7��U&2O1���N�b(�6��Q��[��ع"k�nc�3	���!����(��[wgnK�5[��T�n��j��{%̦�Kr;�H�t��tsUՌ{oFM���3ݒ�\�Ks�5�qmMꗝ��A<�J�e]�^��&�V���Z8\�J���b� ,�$ >e��֣P�!5��{iM%l�$�vɺZ�����ҵ!�m*�Ԥ�� Imh�bCD�鶂���̭2�x�=��3��t䊩wh]�t �˳� �mQ�뵝]s���l������j"�%�k��Ĳl]�l�ʜA�5*�T�
�UPB]@�VJ ^��t�%����t��f �X7f݆W��]�� 6(
�zrYeX�������v�F�[�n�mf�t�V0E]�=��A�*��a�UC�ݡ�����G�<�(&�Pڤ�Um_R��]]��8ܹw�8�u�v-���7�m�:�%�n�K�x��h��2�7W���������x�e4%�{h�q����%�ș�^e���S�Mkg�)Ӯu��`��\�4�%c
�7[��Gf�QDs�s�;lWn�k��ӓ�ŗk��=����5v��d&r7�//GX�����l�=���g#;��:�n����6�6��� g�l�z[ϻ޻�73��ЍF��s��\�*��0ȃ'1�rg�%�Y��Z�6ƛ����wn�]�> wd���x�y�p���M���y8��v'J�c��� ��9�<�e�o�>P�%-+���I��J�vl� �ݗ�E���ݑ�q(tJ���R*)U]��"9%�����ڰ���D���QL����[w�E���ݑ��g8��դ��3�'iڢ�b�2��۶�����F�mZ�k� }/s�;V�{l�k���nݾ7��ݑ��g8���Dr�jx���	��
%B����U`w����IqUR�U�X������| ����e"/�ww�T�΋�� {v<-���� ��9�	�P��n��N���"�l| ���	ٳ��nǀqumBRM��]��ŏ�}��@��G#}�~���g�՛~w{�?W�|l�~vKU�z���]:z�v�{n۫�X�y�M��6�k�8��v�ʸ@�I�4�ET�U5V�^݀{1�@k=���#�6�Ui�J�cM�ݏ �}���#�'d�������E��V��"���ݑ�_W�mE $�=B��R��H����tJ�)��s>���pzG�rm���nݾ7��#��7]�ۻ �c���Soj�܀�!- �T(��IUW@6��=����� �e#�Jĕ�Q�t�5�������ϸ�;��+<�ޓp^;j,g;s��n��J���D�� =���=�u`cu����n���6*��U%�էwm�n�| ���	�'8������hD6ӷcb�X����t�n��$c{]Soj�̔��N��N�����	�'8����v>���}^������G�r�IӦ��ƭ�ݏ �wc�vG�N�9�=�{e]�QE:Lm]5mR�6>�3�m�f�8s	�J[��֙3�x0"v��К(-�����E����#�'d�� {v<�h�1�m�n��c���wy	�ݻ ���Y���""#rt����I*���ݻ ���M�9��!-M�� �n�@��K����%ʂj��y�Y�k�jm�X�n��!o����C��)UL�U)U*j�Y�u`lDG"!{7j��n��W�{��V�;��Q����[����[-������y����Zyۛj��E��MSP��δWm�Pp�E]��p<<'9�<j�2zݲ=s��M����^��+���@�G��:$;U�1ܚ�(6�V���Ǟp���GS�P;*E��lr8x6��9��w���/m��@����m�n�Ij��&ָ�f���F�
��.5��v��!1��x�hUXq̒���4���w{�{������.+l-Q�滱��W]�1�=��ۃ��p��nv -���~%���T���v��~mt��v��]��l|v�Kn1�i���v�;6s�ݏ �}���#�6�JP�մ˲ݧo� ��x�zG���#�;='8�I��h���T���j����H<�k�{sv�Gf:�� 1�i�n۾7��ݑ���� �c����n��Ir��N�����������<Y���5��'h1��q�	s�덍�	�HR�
*&�UU`{sv�,�8�zG�Up�#�=�J%�j�j��c����ϗ�V�T��f;��| ����l� *yV��N�J�V��w�ywd| ���+����p-�x����Q��ݴ��> wdx}6s�yn��<��>�i$��&�N�����9�*����v^�ݑ��#�%wҮ�*,�t�[V5m�Qύڽ��v@�"�W!���������s=1�nwm���E�˲�ڷ��/ ����ݑ����� �e10��v�.�z���^�9Ȉ��ry��@�7��[��	ݠ6�)�i�n۾7��U߿}�Uߟ}�][4����p����=��9��r����}���¾6��թm�����UJ��w�pۿ<��#�vG�{��K�.Ք� ���ݏ ����ݑ����?���u�\��-gL=˒���C���tꭺ���>:v�	q���R�󳏞��w����|�7mZV������#�vG�w۳� ��x����-&�t�]by���J>�����{d� ��x�n��T��i$H�ݤӱ�i;o ���� ��x�G�� ڛ�)V�M��S*��6"#�#��X��@�cݫ ���㈀�{�r�K���)�ݔ$ݵJ�x�G�� ��e��t������d��"TLl��c�kmt��cw'n�Gp�n�sv�!Z�`���NҪT�H��2��ww.]̻̾�{���g�݀{1�@��n��Pm��;�o ����c�:��| ��������e(��]�)�I'o� ��xTݏ����9�x�CvժWM���:��| �������}U_ݏ ���RԴ��ӧn��<��� ���[����~��T�����+�6;��#�+�� �P��)n����&$KS�G1�tt�S�g�˛;�Sv��F�����Ϯ[t�*r�`��5: ��L�R��
s�<ջ��n�Υ�(��r�.�8쌠��0���Md���6����OXrf�1�����m+�z���m<���m��s̸,0�in�8.e��m]��h,��Y�Ȫ��n�ʹ��x�LW��w{��w�����͘�z�]v<][����؛9���Q�k'��q���G77n�݄5*10-;oϿ�������[����}��� ;�<`n���i7L�-ӻ|�[���� ;�<{�9����W� '�-Sl�&�[s�>Z�Հ}��M��B�r"�{v)?^��UϚ��v��y���@ϳ�Y�z����~��&d*HQRP�Ut�1݁��"9̖�zW�?> wdx�ȯ����T�N�nwV���oK�n.#$8Y���rM)�<r\'������V��� ��ݏ ⛱��#�7��� ������V��ٽk[�*�>�߷�N����0�t�z(z vwY���*~���=����d8ٝ��5E2�TuMv��v�}����q#��/�~|v�J"6�����v����owg8���)� ;�<`n�R��V+-Ӷ��nǀqM��ݑ����4����V�M��軵ۯ"l�-�{n���0CqÚ�<썶�4��uص����� cX���M����qM��ݑ���� {v<���L�m7n��> wdx��� {v<�I������ϭUӫ;�o ��9¯=���ٰ{e�; <6$f��5�iл�=]�e��x8�A8pP�sC�[V0�����{J�H�]w�k�8]�1�R*���!���%&Ӧ1��61�!�M#8�b�A�͊��B�T�aت������q�6*ڠ��;+�qUt"���w�=� $��	��)v	�ݢ�N�� =��$����}F��� C�H�M�V������I ;�<3� �c���1<Dl�IB*�5�ϳX� [��|m�F�����l�^��ՍG��8�d�"rՖ�\�c��������n�َ�"/��A廻Vr�Z��JU*�T�)�������A��t-���vG�lԪ:i�ub��+�� {v<�I���#�7d���`)W���)����9'wv��v�cn�.9�L�}������QSSUSSU7U�Հ}��@���{�߀1���I ��S*� Й�Ui�!'�F�v���7mW�b�x�qpn�/���m�2�6��WM���ĭ�vI� {v<�I ;�<o���]�ai�t����f:��G!-�ڰ=�����x�Cvի-:I�w�yI#�vG�n�9�<�e�v�R�]һ[���7��W���vG�n�9�<�e�RH��Dm&�i�m+�������#�8�l[��`y���)��R<ۊ�HAx@ 6��M��SB�RAUJ��>�\W$�h��.(÷\Z5;�:'�Җ������D=u�m��G��F����n����y$칚g�Gy���˨~7r�973i�8jݥ�6Z�판cn�/]��h�rʂ�Mt�F�p���y��pO�����̝s��Wd�\�{v��%�]d	�瓞^F�kG9�Gcs�Pgs*��r	�vɦǬ��m�ت���m��\'!=+ rkV��v�!� �ޮj4�fu�" �z��.�pvn��y՘�e���;]v�������%�mK�۷		i�y�k�����u`y��9�3w`{ 2�P1�$ݴ�����/�� ���p/l������n�V�ݜo/�y����vs����9��[s`?@c;(��R�BSU���^�{���'��=��/�� ��w�˰j��
*�����9�s��#�6�X�n�����L^�H���n9vӴƠ������iҎ78�')3�s_g�']�q��O5�j��N�;�x�> w�<wvs�.�׿~��~�9.��rK�37�W~}����"1*� PL�K
� `OX@ �g���]A�$��l��{m$�#i[��N�S5]��w`y{��r#�K���X�v�a�Q.�U*E$���j�"98�zɽڰ��t�1݁� ƈ	7m!�x쏀� �n�p/l�}�H��?�t2����{��N��.7E�v:cnv�pu��@�������^�uU�YLvڷn�-�| �x{1݁��s��G-�^�X�N�
&*��P��t�c���BF,{=�v��7]�s��=�k�ԁS@�J��8��� >߷����JIP�U
ʮ�O u�o�ʾ��몯��߶�nڻ���&�� I6g ;�<I��mȰ�^�-KI[����-<��� W�U�ٳ8ۑ`ٳ9�������?;E���%��6z�{���kD�[3�-�7��8뭮;(��,ZT�i)��^��䶺 ���<��{R��ڱYn���6�Y� <x�`����������vЕ��f���6l� �r,�����n�V��-����G""#�^�t�{v�mt3��"�:IL��@��S"@��v���:�k��Uw����wI���o ��9�?UUF��V ޽�<n����bR$���t�8�]�97Tm�rt���9�g�����ڜ���	���)/%L��.'e�� �nE��fpl� ��9�	�����M]�Zt�ݵ��fpl� ��9�&܋ ;+�.�[���H2��� <n���vlG99F��] o_���hZ�ƛcM;i]��M�9�Kk�>�jZ�k�n���P����I35	M]��[]W"#^������W����uWG��(�!�2��-,� 1��W�w��E��,��/l��ם������L�.��u��kK�+��-���ϛ���.���kNM;m��.�8;<��8��q�'�h�)��u��.��+TO�;6��`�<�ݝ�Gg��8hg��ŵvG��!��<X�ݷl�=ql�#l�M�軛'h�2%����r��񵱂sQk��]��vm�c����q�ݫ�yzmοq�L����傰�9j��/�U$N�{]�����v�P�2;�g۵�=�G)�t�ZRݍ���q{q��	��%m��USHJit5��<n��7vۑ`��J@۶ջw�m�plu�r �n��������e]����vĭ�o�� �^ OM������v��WE;o�ɷ= ~x�`��B#�y�������C�V;��n�zl� n��	����Ixe�'��bl��:����s+ut����mn�$����x�Ѭ����|N�;�,-�]��e��� ݑ�}'8���ꯀ'����hR�cV��N�Wm�����\����5L���ٜ ݑ�j�q�I�m;.���y6�珶r" ��y���=�b�UrR��HSS���D$�^��$������[q��;��J@۶ջw�m�pvG�zzNp)%���큱�r@ܮ)�P*QP�EB���נ�ݞ�@��q�7$�J2�ӎԩ�	��$�Z��T���S4%5]77n��m�@3�} 1��H�{<����QP��j���ڠ}������<���s��'���v���n���ٜ �I�_H����b�J�2� ��o�wϺ�?o� =����R�q[Gy��m�o�ru��\G �s��<o{`{	Fȶ�STMIJ�SG@��݁�6^ o�fp�p�6��WwZ�]1�t7X�7�봱�q9:�Z�vz76��{v�ODt����4WQQL徾������~ o�fp�p�96Np�(�2�n�wr�������UUU$�� ��9�<���;�Q6�"�i�n���y�}0M���l� �n��PMGĖZ���If$�J�}�}��}���W�{���i('���<�G;
v����x��QP�EU]����@3ُ�y�:-�w`{%��v�\��n����kl��g�a񱝺q��h&��snz�q\J/��f��)��jz��}�3Ι�-�wȈ�#����mz��*����:Yi�g ݎ&���$� �ݙ�=��,�666��ĭ�$���Ix_W�U����0	��ƕ7M���v�w`y6����c�tm��3 �Jeo�v����ٜv8a]}��u�^g�}�U��}�A)�����P/��������.	|z����w%!�p56 b���hD�'�)�0�����c$\���h�L���;�0v�k ���4l����j��� ��L��ҫ�8,P�@"Eم�HlE�f�K@V� ``�>��6�@��
E�N��qw�;ծk7��������m'ArP��E��յ��rX��:W'ZhA�'h!I��q�MU����f�kJ�M�CV'��It�m�l��m`e_7b�:�¥Ӹ���6������!������x���� ]&ᚨ�ζ��[��s��j�2��tH�q֚i����;�7+�-On{6���km�5ێVæ�* �uYY(�nI��n�ӰqnH�\H]�)T����+M8�;t�EEc$kv�1�s�67!q@	�l��RR��ݍpUGMk���Yx�S��q�R��8��`��Y�F�=�O�^�Ӎ��+�w��^t�jt<�<�{��w���Ɔ�9qT��\Ó�:g������Ċ���ԇ1-V����Z#�Yy�ӣj�������8�zpRv���vr��
Д�v����-��B9����pj�C�ΈD���!��ɀ烛fy8��Z�z����j�m�G
����CRQ�ZY��m�a�6�P���`�y���[A[W�1ʸ�3��дnw,�2����rv��6xˬM힠�)!�Ր�	��Ǳղts�j�v����K]�輙bڋ������,�����w�i5Zi۶jli���Q�u�+� �X:�T�J��Pmi�n��(,]h�UR��X2Q`+e)mI���b�h%����l�����D�a�9�jy���z��N^��\k=�גц�n����ÜMnִk�j�{aS4��5UFHv�5�WJ�Ϝ>ץ�km��h ��A��g]��Ӟ��0 �l75x�ƴ&�W�$� *K^�Hen��թ��iIj���핥^����f���K'F��*�v4ܮ�W���(����D.�3 �;��;Y[[&�m<�H���6����.맦�8]��&.8��� +��aej��0���V�=��]5l9i\ �rY� Xe�5�(,�\��l0R�Z�ـ,��p��X ���÷l��Z�1�b������꿞�؈����(�(2�<�$��E���:;WH��7^�3f[�k3z�Zސ���:Ն��7kg�&�f��Z�NZ�ŧ^uu��S�\��,�����j�]�lh�ƭ<F��\�2��9��
�̝p�M5��r�Y$��K�Kc�4�c�컷s:��m���<��F����6C��# �M~W[���2��<�%�5��Hձ:�M��*˚�+Pt���Y5�6��������#��8���M~���{����Ȝrs��fz8y��T�w'�����pN|���@Z��r�����$��m�X�n��r�̒�3�>���@�ۻɷ= ��}���$�Q1R�S4��:�����HŻ����l�L��Dp�r9=��bV�)"�`EU]��wg����o9�DBM�i�>�ݻ ~\1��R*I	��UU= �f>����-�w`s��y6�Zy�G%qL���U����t΁��^���wgyh��l���U%M��y�\�<\m�vS��-�yFh�b�7�}G�Tn�4S(E��v666��ĭ������RK�����0	5K�*�;�.�ܸI|�}���.$�$��U*�DD\DG�)o{`|�i�-�w{�DDr6D�e�(I�i
���?g ݎ&���$��EjR��V�v�-���+�v8`�'8���}�3�zJV��&4�Wmـrl��RK�����0o�����Gi��>wV����ɴq�I�����+�1�F��<p��>c��������6����1�'�-�w`)�$T�J�)���{1����i�>׻v�}��i�K�L�"fQP�9�s�U�o�u��}�W½¤�A�b�b�`	3�E�}���Sd��=�Ф��.�ۻ���}�DD�׻vn֝67���Ӡo�.4���v�nݗo��8`��G��� �֝�7v���)�=]�S���5ۍ�<�1�5W>��ӳH����򐚶�(�m#�m�,�����0M���8`�(�R��T��Tҹ�����t��>׻vn�� 7۳8���W�Ʃ�Zhv��d� ��o�fp��w�9�Nx����UWa����ݸ���s�����r���(�F
�"��<R  �P�!�g}����"�o�v���*N�m� �n��[���[�����@�q�
asI%65kn}��c�k��OU���n�����a8^���^U����v%�<���� ��9�=.E��ٜ޴����v6��BSG@����r8��;������>�7�T�ۻm7n˷��-��g�l؎BM�i�>׻v�#��[E�;i%m`�vg ݎ&���r,�E�*�ڶ���m�� n����d��r, �n��%�I.%I4דֹ�d�Xղ";Tp�״��@�[��G�aź ,t�)�:�:$�n�K��ͻm�(a��i��*�;;�hl��\k�[R��5m�&魄݋A����R5vŵ����p+�C�&��oM@u�nNb������w~���v3�{�s�\tHݎ.ڵ�T���/\���<�<�E-��;�[\���� ��}e�t��[j�)0A�8]�&K�痩RI���m���,�Gf �z���pp	wh[ڣ��,����5�s�f�a��y%���ـ������������-��g�{�3���"!cų�<9S�D
U}`f��� g�l2G�rl����U��I;(T�[m`�d� n��͓���X��V���[�,I�� n��͓��[]���x�{`fJI9���QUUv;Wm��'8�Ȱ}�g 7dx�����RQ�&4���)�i��oi�s�;�ۚ�ӝ���Ί���g#�N�u&-�6��e�� �� o�L�� ��9�=[Z�φҡݧm$�� �l�ք�$�~U�;�߷�|���~��UyI/ ��Dڔ�&մݵ�m�pvG�rl��RK�����(�+�t�-��x�ɲs�yI/ 7۳8�#�;^�]\VP�j��Rm�ycs��c�{��o�Ў{���@�\b�m�^=�vPw��Y՝Kv�q�D��wz^�wbi���f>������"���@��\����[�,I�g 7dx&���r, �n�������i�m��3U�-�w`y�k��"'�9";
9�1�ёrB�5 �,��`.�P���>A�P�yo�~�Ψ���}!q�N�m�i�v]�p
��dp�����8`���ku*�LL��v�Wl�{vg �0zI��Ix���*�:(t�������=uیm��tu���x�G�)һ���۰!���n�VR��V�v�[o3�n��m݁�۝�@f7��5�"�Z�J����0zI��^ {۳8�8`�IW�RiSe;����<�K����ds�c�t�n��s&\�v;�M:I�w�����=$����1����#99�UuURId���y��O��ӄ�7����t΁xۻ���{3l�����o��dM��,�u���/c�g��̠rٓn-��C�z�k��?]��� K�i��t�2ճ ����8��x�ݙ�=�� ��.4�Ӷ�m7n˷���@33lc�tm��H�m(��7t�wi�H�w�l�?�0>�搜l���r,�E�(��V�vЦo���t΁xۻ�8�CV7�h7\"�Z�ET������6���N5�=�����@�ʎr5D�����벐�~󯛰v�����uKƍ�r���ծ�!/e弼[	s=j8S^ѧ��.1����]<3ٺ�7Z�V�^e���>��^�O���v.`�hŧ of��c��M�N�7��H���m�8K&{wi�ݸ�ۡ�'Zw%�ma����Weca'W;TQ-��fR^�¸H��û��<.�4h�"�9�����}��������ܒU�;]n�nd.5pcV��N)hLh;n�v�r�ƽ]�vޞ�gF���s���{v=��T)�����5�=�����@�f;���d�;������x�~ş�$�>�L�c{v�q�󜈈�-<%���j�Yi�b��ݎ;�9�=��`�̬޴�Kv�e�n�+f�Ds��7�X���=�t̬:�2}m�W.��r�%�n������{�,��Xt�1݁q��ؕ�"��=���h�q���<.��N�Bݭ��Ln���p�C�u<v����m���Ձ����9�~���׀wP�-�(��ۻ��/��w~��i/��KԒHIG#�Ϣ����`<��@���;�������m!�-][�e�v����8���ٕ�s���%{e(��j�e'J�� �ݗ�w�2�n�0?/��~��͙�U2Tʂ��it�� ��������~� ݛ���ߤ���+l'Igt�n`j�K��Ǳmm��<t�^v#ϨŰNܮq�
��xsrnG�}`�;����`�̬޴�7X��ն��[0w�9đ�v^�l��9����ﾠ6l.4�նݶ7w	/�^�� ��Xv$�Wi$!(.aǠx�,��TL8d%D�Q5�RE�cO���Yl��c��,�B!��Gf�����q���߾�+nII0Ac��y�DSHI���Յ�牅K��A Q{m�46DfA`F�cI�I9S0W'"��(��i�F�5��*��r�JD7чOSs���g�t�(F��ēC��R���g�@!	9��v�����b��H�(��>�ߛ4�cz7�7;6x���u�Rxv^C ��a��B0�*������%h�fYӣU0������$����`A��$�����!�,�c0��a�M��U=EMC��zU9�� =� 6��p� LD}oGB�T:P^����o��p�Pj��;i��6���@��g@���v����<�k��M��vի|��0���;��8�ߦ�oذ1�$���]�h�"ٻ����-�.�]�<��g��qi�yz�o+�]����i�ljـs����1�@���h>n��77aj�"�O�IҶ��5n��;�X7^�;�����I������'��B�j'h�.`ǽ��y��@���v,�= xz���t��i*����0��9�5o�k���`��bQ�.PK-M��SI33")R��I4��W'�_V�l��B	�v��[0����꯵n��;�2�nޘ��I>��V�q���QHy�ϘG����v��9���N�m�ۙ�\m���
�[m��v���8��x}&V�צ��g8��C�5N�v�����y��Ns���:�{���{��Dr8��q��UJ�UM)SW�֝���p�%��^�I��n����][
�Jh�lDq{�����z�o����}g@�݅�`��UQIMU�����c�^ea�>�����G7p>��pV����p�\W"��H\=e��6��6k�E�^C�ζ��yu�jr��N8I6۷�Θu��r��J������ԩf��NI��M9&�'^'%$��.�!-�����;��m�]��Ѹ�c��uUϷ��"��8��v
5� '��\z3�.v���s���@��ޓq��|l�ٹ�&��Yѻz]��OR�$�v�d��&�����>|~��:r[)[ث��k;g�Fq����}8�v���8%��ˈvx�g�7<]�����ߝ��y��@��g����0�53j�Yt������0��9�5n��;�2�z�Hլ�1;�� ��c�c�����%���t��t�eƕ:��m���ݾp[���L���L���p�(��C�N�E�x}&V�צ��g8��x����g�v㟾��r�����G�gd����<�n�v�W�X��O��۷i�y*mL*�+�vG���p[���L�wɎ�5����r�����%U䐣�@���V���Uן}Ð^ea�7����HR�*�*������z�o��/2��{���qsft�t�EZ'v� ���9���9�l� ׻��}�|I���Ԋө&.�0w�9�5n��;�X=��е��̖�]j��YP�)�:|�:���Lm���wğ��^#��`nα1��m���l����/ �e`�=0��*v6��e�� �헀w�2�o��;���A:Q5N�v�����]���9W^��nXP��=q�#���]{v��=��8�UL�UM]��p�p�9�l� �헀w�2���	��L��V����p�s�q�����@��a�>�,ښ�
�Q����
�`5��cI�d��&�x���^5�2k��MG���\��r�_��w�e`�=0��9���Wv�ubC�ջ�;�2�o��{�����OQ��WJ˧W�����w�����/ ���;�I*6���I�E0V����p^�x}&V>���d�A�CǴU�D��z`H\iS��V�ݵj�8�l���+ ���w���%��/���z� ���{�n9 �ܻn,� ���(Emm�=�\ЛPhqKvբ�w-����}�,����g8�l�����%X��c��V�\�\0��9�5{e���Y�"n�%唪��-4ճ ������^ݓ+ ���M��V
�wn黻o�W���&V��� ｳ� �_K�[I'V$:M[��&,��� ｿs�k��0��T$*��Z}��>ٽ̳z͛ތ��V�9{z�u��oRt���Q#l���^���ٮJ��U�M̇d�!�n;�1����/ZL� �":��LWS�Wjq?�k��;�+7=od�un����9e3D{e�� 狱�7%����K���xۭFzn:MZ�p����c�3�����O0���K��Lӝ,0V�I�=��9�0��[J�h���[��T=D���twنh��(��lj� vʹm���O[d��v�u�duZ�(���l��$�$��V�91p����;�l� �헀wd��;�I*6��,N�)��`��s�j���;�e`�=0��ƕ[i�m����b�9�c}����G��3�{1���(N�N���Ӷ�ۼ�&V��� �g8�l��E�K)4퍶Z���>yL�{1݁���{�t�U�k��G`�e[E۶��7c1ۏb��q;jof�;l���Z7s�f�a�d�j�R�,f=���@��o9�<�t{��f
B�T�LUL�U����s�b3�)(t�9y�>�ʻ��0��9��򖥵I:E�t4���2�}���%��Q��v��_��+�zk��{g8�IxvL�����oi+T&&����p^���Xw�L۵ϰ�Z���A��X�ʸ!Ƿv鵜�ˍp��v�6I�I6�\Ž��S,����^ݓ+ ���w����6���
�6�;w�vI��w|��=�l� �\� ��F��M;cm�w|\�m�`���p�u*�6�Ԓ��u>^�E�l���7��RzR�N��i�������`�e`�=0	�)EV�+�ݵM�ݾp�Ȱ�2����v�U�Wi����q�<��[�h6�l�Q�0�~�$��+Un�t����-e��vR��i��;$��;�z`��݁���@zs.E2�L�B���,<�wy���{v��]�o��9��h٩��u`���������M�r���t<�t�]%�������T��ls��!DDq�n�@���t���~ܬ?!�*|+Ͼ��絛|�uLt+�ۤ���&V��� ����W��UM%�R�+iڡ�rs����n�N�i�.wI��pk�jP��;]�WnR�N��M;cm�����`��s�j����UP�e`�R)�vҥ*�)��{��w�ȈHk7g�{v��g���$k݅�&�)䪢*�j���k7g�}���>�V�{��q9N�i]]*N���
��0}���%�﨩w,WiU�4w��<���9�Ǿ�n����@��G����@**��QEU��O����A_�o9s��
� @D]��(*���*���kGw��EV���?��?�s��������s�?���o�{�?���+���?��O����U�����T��UUW���?��TQU��)EU�1�/����_�L�����g��U_��?����������������:�A\P��	I@��H��Q%�FI%D�Q�HQ!VI	Q `�H!D�Q%�eD�Q"DH�R��e`��BI�"� �
DhD�)�($TI�&��@�
ZP�B�)	!	@��bB� ���B�)f�B	X	YBE�$RB H� B$	VP�` �$H@�!	H	BB������$	� D(�)�B$
��!d	Yd%����# J B�H��2�B�� I RL!B# @!"�(HHHH L!����H�(HB�"0� ��� 2���"� B��)C A �H�$#*����#) @�0�2�! !
���!� � ��) � ���� �B0$# BB3(��B�@H#�(� @�0� �2��2�$#
�2�J���(H2(��  H0 0,�2���2�(���"�+�	(���#J2 Ą #H0��  � � J0(�@$##*$# 0� �!(�0��!�� �D! � 2*2!"�J��B0 B0�#((B���
$�
0! B2$ J�4��$ I(̠AHA R�!(����	(�� @��(+�B #
 J*(*2�"�H� B�#
B���� J����l�����(������u�_�vpӏ�O�x����g�g����O����F���#_�� ����*>?���w ����QEU������?�����?��Њ��٬5���f�����ٿο�z�y�����
�������_����oe?���?���W�x
�����������i�/�3�?��o/��5}����\IU"���������f����������G���]o���t�����W���?��G�����e5��0�8n�� �s2}pM| �   ���@�%  P	 P���IT�T  � *��PP*�D� �	R ��IJA� *�(
@�     TQJR�QQ $UB %�   ` @P*�( O{�.gsS�^�<G�o{�E�����M\f�8�:�nA�@�O\��f� /[���wy � �.��b<����r:���S������w��F9���@{�	|�   
H v� >}T���M
bPd)� h��(c���h4�� DAc   �P�� b   ѝ�     4�(1 h1�  �`ѐ ��@    �  @(
$ ���� �}|�y��{�^�^��Oz��r޳���X�κ��{�co� m��E���㛼 -��\���}�>�kq� �{-��v��W���_}���+� 8��w�<�^{+�x��熽x��@
 �)@ �� ��QŻd���w<���+� }<<���J��6s����q��� �<=��>箼ί :�iy���J�� ���R�w��O���x�s���p �����g-^{�y4��ҏ���$  
R� Z h��Vg}��Yt�&���tw@4�T�_C�C�޼F��xǪ��G���g�!�()@y�zx[ǻ�� G�N�8��q�w�Ǚ���y�Kϼ##ŉ�   O�6�J@  ��T��@ hD��J)�@�dتTJ�1 �?�%�)J� h ���ʔ� )�5��/��O���9����S��ݯɴ�i�zw�
 ���QT���"��UEW��AX�*�����b?�H�B�$H$"������$�?��ٶ6�H�$����Ϙ|�O�W$�$bR`��~y��)��))��p?�x��X$H���P�V��{M0�~���>��4O�Ԙ��*J�����RY�Wi�k{��P� �*JOٵ�gs��\E;���_WR���)�%�JB�I���T� @Ș����eX�n�Q�2"�QK�*�=Dt�j%�'���=��	������cdƺ�������i�(F��P�9������F�!)�)��%�M���ha��f�&�3!0�F6�h���ֵՑcp��;Y3AB�s�V4/b�7	�O�?��i���X1�&�c�g9��2��6˺s���$嬑"F)M.�l���
�"lH�@"��2:�5!Mh*b01 �6p��4�:�S3C�"�H��5P蘛��`@k�`�~4�F��\t�~z��%4�|��L˿�O���0���77�HK���14�"�j��6��K�2�Ri��3Rl�0̺��0��nT�[-��]<aN�_�������&��Ȑ�Lu�ICA�m�a���� E�`M,�B6gf�Zh�*���a��sZ�k7�p�l8�0���%ь!�sD��N����0#Wt����ٯ�z!.k��Ҹ��$`����4h��{�l����U�ɭ�:�ܠ�\�g�H���{
j;b�ԻN1�8h��C�'95�sL�'?|�WΣ��\��9��IQ94�1j���8��!Jlm���k���䢖���s���8˚aa�蕤ZJbb�eav�D���*��B�!�qaYu?h���0�)��8E�>?́��݌�HP�1#A�@��q���=(Y\��g��N�0'�q��a��N~�:C�(BRu=Ją,�Țh�N�*8�tk���]�������z��R����"'��=YO
WW"_ ����Y��9�FB52K����b�ԂD	�`KZ���!+>��A!(C(�6@�!l!�M��w��p�C4a�k�,�*0)��T�Zn�HB�Cd��``i�
$I��1�$2�4����0�O�k��
���oM�K���D�I����	�5$4���
�E�C��'��xfF ��QW
�ʱSS��v����j��JU�\��Ȱ R� #J+�,�"V���Hu�
u4�Ā�I"k�ѿ�p,[ T04�r��b�����o�9�8Hu���,Фd��P����p��@���D��xB����(E�$�#�`SD�$�i$��!aPi!ĎP(t�p}HB���`HW5��@λc��g�����9��g��������Y��� G̈́[ek_h�f��_��!�&�6*j%2;HT�7���r�͙M�'��unn��q�J�)�
���i�ޮ%YX�JA"$N]$2�w����F]� ��U�v��
����P j��'�\������D?���'�d�i�iM����H��C��i?�0��3Fl�@�S��|!YHS��m�ϰ��H��C��'��ġ���>;N	�l!Lӷg �ąS{fR�
b^�껹�\wsL)
B��
�=V!��l�	�5�$�DLA�m<�A�O��g8D9j��!&ƙ�*�!�f.a�҅�[�A�⒐�M��]kI
�,R@n�w�<���f�w���S��U�i��9j�H�9\UJrTOW%q ~q�#B�`H�0�����������m��JB�G����;ϒN?)�&��Rm5o��gd�:]J}�o�Qb�T�� O��W$Z~X���Q�4lѲ~ϡ��K�/��Wk�ۢ QA��"$D�B�Ip	p�5�����Ĕ`�F�l��zM~�!V�߀�X��"T�ӾZf������q?0��H!�$?$���>��ϣ�!�0�?!P�"=�!�<$ Fca���^J�L�)��I���Xl$ln����T��@��B��M��àŎ�?�!
���6�:��N�.$����@���WK��N����U�����|�`|���Sm��F�$��_I���p6�0�k����J�rd�MpS�s�kX���.��5!�pӢ\d��0�l��]�cp0��~E�k/\$�0 F�&9�\��+�#��_�e�XP�1����)�q��|������!��.c))��S�M簪T�)�F9�V8�C"�!"h�vɾ���$�i��CRV Đ�V "%%`@�)�G��LM#�]j�F�7Ĝ% F �|�Ffbi7w��]�F]h�)�&V[��B�$�P�[�����I��r���p�D�P����櫠�n�j�5�2$ eĕa`�S_%��j�7��uԔ�!.��lbD�5�Cl����!��\b�Z%̹.0��$;R1���ߌ8�'����祄#xK�.���`F	sPe�����_~����[�by5B��ĴBކs��W�F>���Iz�����>�ni4l�0�V&5�.`��B�u
*�t����B�!����2o�.Ոݤ.8q�:M:`��ѳg�Z$)����Y��'�\�-���\����N)���J�X�h�}�˹�Eq5I	Bnj�8���+R��D�%�Uѯ߷�}��%WDX���D�VB��VA�d)�K
̬1��	lB�HQ�`��⺪ �J��P�n�V�:*��}���,��0�"�&�Mh��R6f���ѯ������d���w��|�a A6�!C@�� p�[����$�롅�d�0�!��-���R0"�F@���K�.�r� g$����&�[F$0�	���͓��8�L������r��	XЅap$��h�-�.pՉ$��VB3e%,l�!im>>ٽ�~� K�O�$c\��z+m��!>炳���m���U
*�rje*��(-�jm)�Ɵ�"�8�o��>�рȡ�ď䈍t?3�JƓ_G0���)(���K��1�l
� a*K�ZX'�!>	_�{��h�i��8Y��j~����h1`A���2a�!_y*�r��A
8.�ĩ�N�\H D�)52G>&c.1L��.*b��/Z���Y/&��F+�.�"�Fku"1lJ婮%��ռ��P�n�
h!��p�&�6Ư>�e�4�!u�/s�Ϟ��1 ���C��p��9[�\B!��L�<	L������#&jc`A�q)��iF���5	J�H���BP�a����,�@)!e&0�!�P� "cAU�%��!Yr���D��B�L��^wz'6��t˄*B����I �)��5����L�uq�B�J�h��s[��39̛�eԖ����F)3L���0X�"�]Y���V���H��b���B�UHU1#4
ġ���]&���*y܅�5SYds����*�arg�*�w�}��hϹ�oH�d �E4�.¬B�Q��Kg�!�S�(¤��!+��c�HDlB�|l�>�aBH�b4�ʟ��������qѶB0��m�&ɭ�ѭa˒Ϻ�]��w��䬭#X�$	!HR��a#JÅˈR�,�%	L�B+��D%u�p֣��
D�di�B�
I�Ew�!�6F�I ��X�`vO���	%n[��w��?p%e4�++���\5���<!&�얐*B�H��q�I.�u����(kN�F���4+��+�F�
�b`�CFfU�ja��P�7>ȟt��/u����1"O�Z	!

�)�փY�p>N�c�Id��!�2���I����(�����?P#m��    p   	�  �  �       �`  N�� $�m�      �h�` �`         �6�   $    h H        p6�     �SgF�[j ��\9d]y-��B-������[@R�tX�%��n�+嶶����̶�+m�W@��:��vĀ �M�UUT�@,A˳�.Kh< l���N�m�R�6ۜm�RiM�x�j�ڤ�	�0sm���]�Į��Y$5�m�U��^d����;nx��mQ[�@@�ʧL�1J�l�v�O2��A��m��YV����z�U���*�t���U�ʛ��5U�N��Ul��R��ʫ�j��[�Qd�0Mn,�^m�m��䍗�Z[vg��z�U+�eI[G���v�z�q�=9�[�a��]v�I̋6�{-��������:�7mcc�vW����͵������2�V�gC��y}P�GjyV^s�.j��m���j����N�N��/��U_��)^�Djn��ny�m�nZ{'gv�㚀Z-R�Y����*�V^~��>�� .դP��n�`�$5��-�څ�B��4*��cK�Fl�p�%n�4!쎔�$A͵R�k��[��v�@涪����@����[��ņ�,�����e�{%�[�É�s
���J�EZ��p�yZ�$t�Q���ݸ̷AvF��Y�j{mهsV�`�3*�lUV� ;�i���m�6��[@  n�[CUm�[{  �n�I�з\�	�Y2I 	hq:� �mrUr8n�l	p*NhU̫�nݞ��+����V쪻2��Z�u\�!���mz��m�u���mX#���d�$,�U�]�
��U�#-�p���z� 	 8t���#���]nǁ÷m� m�88�� H�vٶ���Z��:���T�l���
��eYy�U�v��I5�{� [@� 	 	���cl�� m��	޶�dm��m'   	ЖP�č�.���`*U�j�� V�_Ar����� 6�6�l�i,� ���ݗ�ڶT��h6X.�4l��֛=&�@��n%���   մ Y.�ݶ  �h8 ����   *��W�� !�7V�P]�nzR@\m��R���ض�I���$��P �UUJ�P �oF+ko`���/T����$m�  �.��-Hm�(!KVP�W��İx
�z�����T�R��P���  .Ki�o�ӧ��Yd����dm�����m�k�m����*�m �f�[RJ��8���]6S\��;vܣZ�Y��;t��Ӎ2h-Z�[�sOf r�m��*�-��vrcS�+��-R��ġ���fـ��A���WfV᫃�Z��V�"Kj������j��,�l�	�C�I0M�Y�q�͸6�v�R�l�[��W�\���  ���Hu�[m�� N�rY@�^�հ[Ku�� f�Z��n t�  Zne����^�+j�@��[�Unπyz��,��]m'��hH�� $ �kM���M@�8 �U�-��D���!m-�Ji(�M�k��Ί�v���G � [R Hp�v�Ƶ�0[@�M��en�
vYV��5ݶ�P��U�=�)-�I���lk$k�I��ѭ�l  [R�� p���m���8�k�\aT�v� �uԷsmm�6�$�_���}���6�d��z�	�=�*��*�v�"� H�k��m���m�Lݶ�N�#i0�=�J�UR�0vx��ol�)k�i�`�]�Y猝��C����.�pq��\�*h��&�V�QOҠ`�k@7�*`�p�lKgJ�\�!�Y:ɀF�fY�� � 5�9�@��N< H��ɨm�tkZcH6ۄ���fm�I%� h   �׾>��v٠:������ 9�   6� +�V��AyV [A ���[sm�h 6�f�9n�[&��om���IĀ��� ��@9 s�� �ˮ.�l�M�  	t��Yڤ�-����>�� [@�@[Cm�  [��4�jvm�۶��[� ^�m{  u\�m�v�v�!��[M�I��lؖ��Yp����,��É�����V�UU� ��[Uu���\�l��)E�¨���*�J��P ��m[:MJ [@�i ��M��� ݶH6N4�\6�$ �� �d�M�Vꀮ�UU����\ i��� ��Z p �d	�$��(WHL���U*�e���6�a! �m�� � ��H�YC�-��]6�m�m�] ��dת=%��j'YBF��p �����@=n� ���i0t�㴼�v  &�L2���*��O,����J�@  ��l�aS�;i0 [m�{m�^�ޫ���= m�زeCb���7:�`l��+.����o���t��.�M�-�k<��(q��+�vN�ؠx�U����m�s�P�U�x8�SAmP�Z�$��E��h-6q��k[d�Xg]3b H      l�1��Ayn����� �ݐ �òY@  ��k��m�D��i��8�nذ�0�$mrIZ���r�pMmZͶm��-n� p    m6�` m�X���hp6�  �g8�f� ȶ�i6  ��cv�:n�z`8h"�ְ�H 8)N[@� �i-�&H�Kmְ ݶ[�רp�` l[dΆ� ���ק@   �  8  m��C`��@ mm���5��m���@ /Z-��	$�����|�  ����  p    �G-� � :ٿ7۾�A��[@I���jݰ� �t�p �����a,�;
���� 6ۂ۶͖��a    m�  �lh   �` ��&�ۍ�`  $   9͢R@  	 	   �H  6׭�  �SZ� А  �dM���e����}���   ����Im �` �ͻ`[AkM�l�N����      ~� �Ә�`  6^���ͷg  ���d&�ۀ M�	4UmCv�p �g6ݩ�N���孶���nڀ��@m�$�5�1f�Ԗ� l �09�n�N��%���7mq͒:@����5�ѱm&�J+`:�� N�M��9����h��Ίpke�G`[8�z�.E�JtJ�v��BCm�ەY�[(�UT �5 �L�  �6�V�� �l��6݌�     ]�啕j��t�UTs�ͫ`�#��   ��m� >ݴ�|[e�������X�(Vj�@�yh
��5 W����   �m�  T��\�X�J�UM�p �Kn�j� l 	������m��:��U��R�*�V� ��� �[m��Zl   ����k�N �bYV��*�V�j���z���Zm ��vs�۵�@ ��6�p-�H.�s���e����n�$[d-�o��ݲ�ձ�� �o
 |m�ڶmmͪm&D�  [�[,��oi2�I��u��R�+���~���@�4m���2ٙy6� ^�$�y$ݛdi�-6H	��L�}�|�㛑ӧC���� �v쬫�ŵN�L�v���m�ƶ奣��I�
�]9��d�>���4 �N����ڔ��M���(���QUT	�'3���������ն�h hu�4��?'�[[I� ^��kz��b�  -�m�� ��uͶm�&�M��� �   ��n�Γi6�v��6�pHH�8m�� � �V�H�P-�lvⶻ�u� O%A[�9��F��â�K/m��W6� X�kR�� [F�m��&�h�'B�ں��6�'4��4m�-����I�*E��͛�:�,Αͤ�\�t� X` u��h[@�U�=9�h
��h  �y��lm�UW�j�wf^�PTŻ^�j������q����X�ev�I6�Ҫڬ���.�`�6��3UTa�>���v�T�j��D�۩C����R�WUWAHT�-�Cp�̫UUR�f׉<�R�Rpvݦ3tum���rJ  [%.�@� Hh�,�� ��ڕ��p �`�#EA��_��p� l lm��� p�c`  �Jp80�m�lm�[jf�@ �  �,��l l� m�h�R�PU���v���l�UFEBA�t�`�[��  Ͳ4f����Z�%3D������b1����?�a����C?��W��Dq��@Ȃ��*|V����b�Au�� ���D���\@P7�~7�?|�ȁ�v)�?�~T�E7��Pp0�J )�,�&�1 �Fr��lυ?$E$F"$~S@.��W����C�G��T��S�|���@���i�&"��=H����'�@8"t?%��t����P�*| .πv� +(�T0 0�P��A�?c��P�/U-TB��������=��� �#����t�� ��054:~x�F)�Q���M���QN�zb'��~O�a��u���Ž��T�)p�(�Wg�Hq��A�T~QE���%^��1Mp����A:l/�z:�&Ȩb|*�e��:��> F �0L�Q!G�pS@�W��Ez��4�56u���_���GH�:/�~W��� ���"��~PWhH;�D?}����]k�"�<Xi�@`@Db!��TT���"���h�U���P ���1(�`!A"��h�h�V+bF��(� e���kZ��l6Z6�m ph��������:m� �-�l%���Ϋ%�5��Z�5�'e��N�Z��uF1#�yZ:/\\>ǁa�ŋ{<�F�g5oh�)؈�S�[���V;;.�2��8�H�N�pL��-��仠���]�y|=\��"��$��=[i���2��5�G`U�j[�(�5)g2�)���vwfV��x�G���ʴO*�[��Z1���룱��فb54�z`��EF�zN��u��M�{k����5-tU��[{,�]��nɶ�V!�
x�'�حpl\fױE�!�W��P 
uh(5�vױ�v܉��ۢ�=�q�)�VB�ok����;S\Ŝ�/Z�
��S�@�m]<uSgm�,�Rt$���S���i 'B���qQ���]d��%r
��X9wJt�wi1A�O�Vf
�n\�y���[Z]m�5��h移`�S�=$v(��639�#�Q�6�ͫ+�-�s�v��2�QzM&ܷ�뚉7G��g�.Ģ�pՐ²�x%�����g������ӻ]a3q�[tvF��GA�]/n�B����g���ĳی��^Gݧ����N�6�k`e�䶸��'>UY!�/[ �c��1jY����6�]3>L��m��%R�e��ܰZ�v��X <Y�	ؠ��v�v�鹜W�v�tm8�-��6Z������۲[҃���F�[ЛU 5��6� ����-�!�;�u�˭�>Lci;e��u�etk��R�*:ݶ F�9�ee2��I�.L5J��X�3�ۚ��孪G��;�r��8z��ͭ֔���0u��
�)�0��T�{Wj�ʚ��*\��2�7Ah����
�;th�vKvѱ��N���6L�����	gU�܆#a�$�5Hs��y��u�9c<���Nʹ���3�-� 0[��\�Su\=l��v����p��ң�w"��[Z5Y���(��0RM�bA��8�~P��D���Ι�.���BD�M���&"��@��b ��|�D?(�����<k��	�;l�v�.��8mt�S�x�����ճ�uVr#�Jr�
�%ӓO)�xe����\a0:W�rGD.��6�w��>³�}���b��	�d4�.p��]���s�WT�,�H������F����x8؀��]#ٚ8�������c�M�N��:���[�)*�qt�r.�hV֘3�t����%rf��U�:Q��Y��	�,˅�2�nx�0<+��y�3��W�`�;l&1ȯ;�1�>�:�w4�� ���h���(>?ĭQ$̒IJ���i�z$��=^�F�\�����1��2�at�b��4�:4��"RI��N����z��Ab�M&�^�z��hޔи�e�@�ۍH���6�mǠ[n���M�.W�ށ%F���YY�%w�B��3���5i���h���.0vA�+�#m	�{'E���2,G3�;�>4l�h���۹�w���`BFbn�֢��V'�h�R�@�cn��/@��k@���6n���|�/W�3(�:�n����R]�!�I2a�y�)����1��q��m���$v<��$�F���w�~u}9jĝ69!'3@����m�����w4�q`)��q�x���0���D]�i҂=��;��{<V���\�=sƣ�t��{"�䆁m�����w4oJh���H@�I����I�d�I6��q�oSlp�c�����m����4�0��T� "Љ�!d�����F�:����ٰ3���*(��_�0���Қ�n-�������X�Ma&&�^v��9{k�/[��{zS@��(6�黉�.t��M�r��m��ތk�e<��}��)m�ʻ�]�CUq�ۗ�������4��Z���EM��8��/[��$w�|hW�ش^��.<�4ī�BNV���3@}��i+�5�/@�M����i��Ĉ�29!�^v��9{nnI����ɏ��8"`Y��D�ʪȦi�9�,�H@�2ҵj򕁑�ٰ77mXܭ,��Q`y���߿�u�~6�^N�z	���܋�q��6JhN�V�3����t;�Wn)�.YWj����rmh>�4�n��? ����;�S�H)�E��hޔ�/;qh�������yŀ��Ma&&�^v��9{k�便}��w�|h�;��e�1ƣnI1hNq;엠7&ց��3@��t�ݼ�4�F�i<��8��w4���߻�~8z}�Gwf�iq�j�iJ�����BۤEG6��J���
b&0�(R��$PH��$г0 )��Q�)��������[;v}/]���%�f^���v�Ґ9i�,AO,�-����W;��`�z�5�m���m�6e^˪w:ø�F��bJ��ɹwF�Ў�a��a����I�����l�M���Ylv��J��g<^s@��[J�J�.7���ݫ�"�:6oE�a�q����m��j���1e-��r����;��6���=�8Fu��I�7V�i�DL$��a��1M�Mtw;��!B�-�F��|�V�eM���쭓Z��s�.	�խخ������;�n-�����s@��S4��`��2�0�;��KJ�W5�/@�nhޔ�/�^�1Ē��Nb�9{k�=�w4oJh����B�Y�fd�ɐ���ܘB	hM!1�{}�`s�^,�2;����u
D�8a1�3@����߭�ZW�ށ����%W'ej����p��OY��5׳�)r��&]��=:'�A��'?X5L<��A�!�x뒖���ށ��ڕ\�~A�h@��?��<��Q7$��
���������KRJUau�j��ei`gguE��1���&�y	q�޻����v��*�נ_nL��+�fP�+BUs���h�%-�����s@��S4��~Y��$����t�	ʗ��v9��7�f��n����;��Nٹ�Ϙ2k�ɵ���&ͥq�<�Ź�wj{j�0��A�Z^��o]��Jh��WR�R(�أ�N=��s~���$G&ր�rR��w��J�u�f%Q4"��Ұ77mX��Qd5i.-�hY-%�.�bk�`ffڰ9��%J�)q��)3@�]��
��@����-�s@�;���8E�b�*�^��빠^�s@�]��Gq��:`Ͱp>u�)��{]Wy���3v���o
qJk>�r.b«�IO�o�빠^�s@�]��
��@�ܙ��+�$��	��-�s~�ċ��h9/@���l�8��Y�,�qVYJ�$��^}�@��z���z���uz�N HƦ&�s�WZ�om�svՆ����	%i6C���_�U�<Šz��4�1�4��>}{Z�O��ے���[�����>���2��t��U!qv��7f�t�m�<�a���5�Β��;\��z���v��*�^��빠y�f�l�&�����VvwT_�I=i!&�CCM̞�_���o�X���R������B(��WZ�oJh���;�n-�(�x�m�BF�z���z���v��*�^��ܙ��J��$!�s4��hs��WZ�{��ff_��ˈ �I��˜�r�&���6Ӥ��k����E�\�s�z��r�/�N�Q�jn�^�ᶀ�u��3�:�;)��b��+�Ƨ�g�R-��q�vX��v9}�X)�s��lp�Ν���n���8:4�:��̧
�b��ɰ<苲��v�M���Q��RD��v[��@]�m���>����]dkAq[�&˺݊N9��'mq�]\m�U�Ҹ����w�<m&��/nz���'������u���Hy�k��q�U	�AaV6'��x�x�ܦ�w�m����>�Uֽ�빠^�s@��&�� �i�Z]k�=�)�y��Z]J��4�1�6��=�q�)/��K@��^�w�J�ٖ�F7D7!�^�M�v��*�סqu�s@�0x�aH��s'uE��KӞ�����s+K
W)ګ�rF6G��Ӄ1L�p���t7b��Y^��n��F=�֝�P���ۏ=Z)$��$�](�$�����Ē�.�����(��Ͽ;~�@��Y?��9f�f�n��3��9�| HRcR0�e�w�i�ǈ�.�����K����Ē�����nnbm
��$!�s<�$�K�Ԓ^t��$�](�$��|�<I/]+��6�Lchq�jI+��^x�Ut�ԒW��<�$�K�ԒV�4y$~�����%WJ=I%�R�3�J���I%z[���� �z{9�[5�IXMi52�ԧ���1�O;�y���m\/|)�Z���D#��$��}�y�I^�Q�$�Kqy�IUҏRI.��n��d������[ok��~U��}�{��-�׺��%�_��<�$��L<�@��&�F���-��$^�����30ϖ/�06�S�h���Q%E '��B��f������j0�"��:���$!���F�C*A=� O����c�?$��������(k 
�Cn1!T(~O��p!-��eH��H1 �r����6�7���lqU�c޽6�7�u�6�]�Z�#��) �F�#���~����)��)��?t������8���h<8M
��V��>L��d��a���O�p�USJ�T0v�Mh2]s����7m���5c��<��I$��$^���I�����I>��jJr�����)~��]P����hm�q��ԒW��<�$��ݛ�����K�[o��v]�m� 	�>��߆{^�B�x�=�m��t<vN�x}<e�S'na��ŲUk8n���+gڍI%z[��H�)5$��|�<I/]+��6�Fchq�jI+��^y�U]�;2�$���~��]�=F���������@��	4�/<I#��RI^���Ē�Q�$�Kqy�IUaR�bKnRU����x�W��jJ���z^rۍ��V�F� ���֡�O�WzU�DDnb������UU]
�~I)����K�G���$��fjI.��7RK��Vj�i���&##��'E�>*94ZCv����r�8E��nҖ̯]��D�dPjDjI.�u��$^���J��g�$��u�JҬ4jŋ����L^x�E�I�$�[�y�I^�Q�$�Kqy�ߛk��cO�D6��q�jI/��y�x�]��5$��n/<I#�)5$��'�V�@��0bs<�$���jI+��^x�G�RjI+���x�^�+��6�Lchq�jI+��^x�R�{��J9?T��IG�Q�$�UmUW���~u�w)v���fp���W��F����6$��&#3DS�b� =�s�m]��Wl{C�޷ng�{;BL��#<\n���_����|sn��in����c���ok��wZ��u�7���l��"��!���n�60;t$�g��`y:�ܣ���g1l6��Tl��W/�ݤ���QT�ɤZ�tbk-�����QҖ�7{�������>�m�;���m�v�����+Z����n�~�����7l�H��ܜF����ܼ�/��jI+���x�]��5$��n/<I*�*NLl1���6�&���o��%�.�RI^���Ē=��RI.����"n2HA�ng�$�t��I%z[����m�����K�ߏ<I/h�'��N0�5"5$��-�����O��$����Ē�Q�$��XhՋ0��I$��${e&���W[�Ǿ����F��󥸼�$�9l�)Q�Y�臭�ܔ��a1����;����gd�3�G��35�X�4�D��q�x�K�ߏ?$�{�Q�!~�7K�\�9��I?g�jI.�������L0Rx�]��-T�I�	�v���ƹ�m���j��o߿o������wT_��~}.�:�)��� g��W9wkJ���J��N��v�u�δ���ũ$��*�L� Hs�L��I{e�RIu�O<I.�w��]nY�%]�I���n!%��"Ԓ]n��K��ũ$�[�y�/JMI%�wcR�Y��p]�9��g����nPM���v���.%0;���R�r�!p�BΫYM�y�I^�Q�$�[�y�I�I�$�ݧ�$��t�Q'��Iu�g�$�zX�$�[���%z]F���a�����H&�<�$�ғm�����s�� $R��ULs3����z]F��^���Ē��b`݃Q<n8�p��K�m<�$�K��$��l�ߒ^��&�Z�K��q����QE��$�{oijI/W9^��x��$��5�Iu�$���O�jM�g��Ly&޼s��Z싨Ӱ=��;%v�xz�<��[� ����x-���M�r��߰ �����~�_'��I%��d���ZI���I%+�*L� Hp7!<�$�VQ��g���bS�|~��Rg��Iu�g�ҫ��*��~����,`8V��������~�;�z�JW9�s�wi���$��B�$�~�b�$m�G27!�/�g���n�⛶�{�zk��߯uٛ��
����-b!�
�?��Р߁�P-�����[o}3�\&��"q�A��$�[I�%�����?I_��y�IwK�Ԓ^:2� y�$h%�;��v�K���q�zҙ��{lC�v����="�L�Y@�nL���\��'�$����K�]F��]z��Ē��A�N� �R'�$����?�?�&b�=�ԒJzz����[j�r��/�Y�|�(�&,��$���F��]z�~��]�UȯRI8��$�����Z8�cC�#R_cn�~��%���z�K���ߒ^�d���5$����Z?bH�UwyY��I|��z�K��U{����II��jI%��Y��I>+�]��­��,inV�t�gn]Yl�md6@a֊q�����V��V�OQ�&��xٗ��c��y�D]Q�U½P����)�c�@��\�!�/a�m��Î�4��Ӥ������$l*��I��nh��ɺ��Q�U�hrE)Ğk�199��ݧBX����2t���6I�\v5�8��=*���n2˚4f��>E@٭��u�Hh����2��]]�4�y:����x6:�s���N�{����ѳ���0� �7���%���jI%�ْ���]W"�I$���_d���4܇�$w;��M6��a�Ҙ=��`f��E�������xj D�"�R- �i4=��%~��@�w�yJ�*��&0�$p���V�ץ4}}V�ؕ�w�x�?��I���@�Қ��_������}_v�N��}�ɮ�zڋ����;We���y���pp7g�˳k[9���v����ƞO�	����`�w�m&��S@�Қ�;��$
)&`��� ��*5ԡt�Mh��2�֖������܇\�h}}kg'I.�V�H�X����4�2_q�{��U�w<�{�3@<��Uue�B)Yw���q�4��Z�ٚ}ܑh�Eʼ�Y����-]��_Z�=��������:���ｕ<TP<f'���g�Mu����s �V���ns�`KR�s�?=�5�,Ņ���R������d��8��? ����>�U�%yu��2�b��*�9�ڿ�m$�!��MU���`u�������H�h���\�X+�-EUU����`s��KI,+��JRI��k�O�|U�w}�X��+TISfe*/0М�_wZ �h��Br��a�|���RV�eYv�e�����')}�3�<�����Zi����ŝ��k����%����h���ٴ��7
'k1l�x�ڟ�w��Н�lq� xۙ< ���@�Қ��W����[�>M8c�5�CNM�Jl�$}ۑh��}כ9ă�ԹK$Q� �����z��i����cs٠OL�~��+��eb��2�+�ЕĜ�� �\�����.ꪀ)	L �� ��VB@��!�&��!&�]����~vO��Z��"ǌ$"Q��4��@�N=��>�ȴ��4�g����N�i�M���v��Zv��-r<j�r�P1ٵ��N �Y��e5�x��a�.�fg�y�������s�_X�f��W�y^�bE�Uї����mo���f�w�f���f�H�6��%e!VU�j�^- rC4��y��ܻ���@��?���V�H�X����4"����y��ִ=�$�h�"���g2�IqX����f�9_nߎ o��d�ŀ��%4Ɔ�V��t�C��|~���'�HM�P���H��E�!��$b$B �(��B�(B�R$f�;���y��1����f^t�<�j,# ����@`���$d��R	�Bp]B0LB�A>>g�%e٣X���0 BH!��2)#P�D�#0"!���4��{P�W��ԗ2�]�4d+�gx�
�t�ZIvACK��HG�A��@�`Dc ������c�hs? W���e���3�F���,��c��`O�aWZ�I�'4��j�Y�$!D��{n��<�]��\w��<�C�[M� H&�8-�k5� ��� 8�*զ�K�	�����n��*���ڧ�^pg�Kb�S�l8�y{Y�|cp�ɽ�]�N
��J���D�F���ol<We�Sf������c�N9���҂��p��BT�`��!�l���Aƍ�r�Z-�F;i%���܋!�\F���Փ��3iᑫ�:OcMm�W)�z�֮ݎ���W=I���C!4�� Q@t�J�c�����uI5�d.z���`�l��bu\���l��\��,���p���� c.c�qN�<�� N'�n���92���I�i%�eg��˺��z]��l]�ɰ	n�kH���`IP�〔mY�]pl�E�[n��ix�%�z�=�˥��U
��5���e�:�|q��l�6�����e���jxSk���U�+ֆ��Vɺ���v��'�Gn�]U����#��Z-͍���;ح�N��uR�M����[[n4�ʎ0��[m)�F�����NG8re��\��x5��ƣ����qu�o6�+���"�*$g�}Y�m^9^�Վ�-'�"�۶ y��[�[�bn��^�CM7K�i�vYZ�ck�V�,�nӔ�0��/[�پ��s&h�#S��kjBN�`-��� �y;j�s8��m���8d��VT9�^����aʄ�.م�ڠ�Z�7;�h�jU�B{m�˱ok�;N���[k��1�s��!z�
��!R��6�7I�g[ 5VӉ hӈx~�|���m#&����*��ɓn���1ĻRc�Wf���ۊx�f�0$v3�U[f��y^��t�N�`л��qʥc�QG�n�vI��z݇�u�h�h�S���.�&��iU���n�.�Ez坵y]9GѺ;S�`�{<��q�D�흲�a�V� V<#ӻ8����sTJ���ٶ�w+6�Skn� *���-m�c�Ƃ&HMe@�W�'$ф���E�l=[����{����p��Ɵ����"G�;A�C��	�'� z���J[I(�*	&L�A �u3J��%��ç)��lW�l/�4[oJMQ�G���9���md^1����ںѴV�h�h5]��\������t] m<�q��vk�9�m=.�W;�����!�\���u#�i�M�:x�n�O*�����(A�v��lvDݜe7���Xr�˦7����A[W��C�*���vSu�zנٺ��ϛ�;�V���ۂ�w{۽��w4�m��u��+b%�&��mjt��s�h�뎉����8[2�s���gcs6�!�}�|h[I�yϪ�:����Z�o�9����4��7�Uď���C@���4�XGT�a!m7	�yϪ�:������U%�y rC'*�_�6х���D�A(�Z�ύ��M �i������j����J�ZY����@���4	I����Z_q�ԫ�6�&���F���)�sc�b��ؓ�`�Wc[�ҙ�tA�����}��c�r�a���?v�֓��#���mW�DȖ%������r%�bX��{�%9�%.R]Y�f�5��Kı>���(�R*@Ah���Z�T4�&�X��ɴ�Kı?w���r%�bX����������ș����fkZq�M[K2���r%�bX�����ӑ,K���ߦӑ,�,K�{�[ND�,K�뾻NF�j�j:b��D���"��&���İ���ߦӑ,KĽ��5��Kı>���K��dk�{���j�k=��2���DҒ��Y��ND�,K����ӑ,K��뾻ND�,K���6��bX�'���6��bX�'�N����ə��&G���z��n�5�n����u��s�n�k`��ww�;OŜ�ڴ
-��r%�bX�w]��r%�bX��w��Kı>�w��P���2%�F��}�V��j�k��L�>�b��S.��v��bX�'}��m9ı,O���m9ı,K�{�[ND�,K�뾻ND�H
dL�b~�ϥL|�&%MD���j�k=����Kı/}�Mm9ơ�d�\@"~���Kı;���iȖ%�b}��rz[�YM3.K��r%�g�L�������r%�bX���]�"X�%��w~�ND�,��>�}��BE>�;�0ޠ!D�"��3TU��4s3i�@ނ1S���6��bX�'�ﹴ�Kı/}�Mm9ı,O��y=v�w���ZN蛳�����|u��.��2�����;�z~��W�@q�c�w�{�K�﻿M�"X�%�����r%�bX�������bX�'���m9���{���?���5)qis[�w�%�bX�����Ӑı/}�Mm9ı,K����r%�bX��w��Rı,O��p���\ѓZ�Lֶ��bX�%�魧"X�%�}�{[ND�lK���6��bX�'��si�����zs�L�*�����*���A�ԍO��궸5P5^����Kı=�{�ND�,����!v�c ��#Ră
����ͪbBQY��DW@��>Ͽ�����bX�5�lL�>�b�%Q
����@�@��w��Kİ� {��i�Kı/�������bX�'���m9Ļ�oq��n�����tn�B뱪�K��ú���9��q��㜦�zd2sp��������=l˚�Mf�ӑ,K��w�ͧ"X�%�{�zkiȖ%�b{;�fӑ,K�﻿M�"X�%��{�'��]fSW5�ND�,K��� ؖ%��｛ND�,K���6��bX�'���m9ı,Oߏz�9�%.R]Y�fh�ӑ,K��w�ͧ"X�%��w~�ND�,K��{6��bX�%��[ND�,K��Ojfj�-�I���r%�bX��w��Kı=���iȖ%�b^��5��Kı>����Kı>�ǽ���DLR�U0MQmpj�j�s}6�"X�%������m>�bX�'��{��9ı,N����r%�bX�@M$@��N��2���5%Ԑ�-��R��肧��m���F�Iy���(�{�\��6.7�N���g�X�6�wMu��'nj�������,/0<�KY��-t����gw<�F�݋$Om���9{l��;tݙl�(�6��]�J���fM�v׃�ӳ'H�ͭcmڮ�^��fx65��\��b�����zǭ�	8݄� �m��v���]k�#�k9�8��$ߞ�wu�����Y^��h��%�z���fg�됋��ss�Sru��3+�<�N�\ѓZ�[��'bX�%����[ND�,K�k��ND�,K���6�7蚉bX����6��bX�'����(S(
�!T��*��5P5_{]��r��"dK�����r%�bX����6��bX�%��[ND�,j��Ad�=5�L�HT��\���﻿M�"X�%����fӑ,K�������"X�%��{�ͧ"X�%�����I�2�r�շ56��bX�'s�}�ND�,K�w�ֶ��bX�'���6��bX6'}��m9ı,O{���[���&e5sY��K�@�N��V��j�\��y{鶰e�bX�����ӑ,K��~�iȖ%�bx�J]�$=��!u4iԺ4�m�uqa��gg�돎ݱ���k��g����6���L�ꀅ�TEUUq��@�@�O��m�D�,K���6��bX�'s�}�ND�,K�w�ֶ��bX�'{���k4�5m,Ժ�m9ı,N����r��U\wq,N�9��r%�bX�������Kı>�wٴ�O�G��{��7���������K���o�܉bX�'���ͧ"X�%��;�k[ND�,K��}�ND�,K���6��bX�'}��'�4d��K�ͧ"X�~��.w�ֶ��bX�'��}v��bX�'}��m9İ'�L��o��k�P5P5���>�S,UJ�h�f��ND�,K�k��ND�,K�{�M�"X�%����fӑ,KƳ+}Smpj�j��z� U*����guI��r�[��1�5˓�8-��k�Շ��y�=1�]gC{�[�oq��'��~�ND�,K���ͧ"X�%�����fӑ,K����ӑ,K����<e�2��njm9ı,K��{[NC�#�2%�����ͧ"X�%�����iȖ%�b~�w��Kı?���s'�-�B�X\���k��Kı;�{�Y��Kı?~�}v��c�5$9��y"~�w��Kı/������bX�'��}fՒ�]Y���j�9ı��w�iȖ%�b~�w��Kı>���m9İ?�T�Tȝ�����Kı?���YsT�a��f�֮ӑ,K�����iȖ%�`����ͧ"X�%������9ı,Oߵ�]�"X�%�������.��L��Vg$�:玟X�+I��r��k��"`w�e��<s��l��S����~����{���g��iȖ%�b}�t��r%�bX��k���,K���ߦӑ,K���\$�T�5�%�fӑ,K������ı,Oߵ�]�"X�%��{�M�"X�%��~��i�%�bX���M��a��Z5Mj�j]�"X�%������Kı?w���r%�X�'���ͧ"X�%��u�K��K�k��VG�STUD�D�Qmpj�K�{�M�"X�%��~��iȖ%�b}�t��r%�`t�W�v?�D��O{}��9ı,N��w$�e̹�rۚ�ND�,K��}�ND�,K�뾗iȖ%�bw����H�����mpj�j�Y�򀏗~�yy瞳�u�y�\�+�5�]���uog���|�}=u�:�w��>�����O���Kı?{^?�ӑ,K���w�iȖ%�b}���`r%�bX�g���r%�bX����sVJXaufL�5v��bX�'k��N@,K���ߦӑ,K��=�fӑ,K������[ı=�x�˚�9��iu.�v��bX�'���6��bX�'���6��c���"dO�׏��Kı=�{��9ı,O��z]f�)�tSWE��M�"X�%��{�ͧ"X�%��u��iȖ%�bw����Kı>�w��Kı;�zL�'�i�j�3Y��Kı>�z�9ı,N���6��bX�'���6��bX�'���6��bX�'Sg*{���?8��;p'r���Ԯ�ꮻ&+��}�l]z�ۃU�L��G��5��I��g@�Q9nK�Ӹ:�����!�- �������[	��T��1��k��^��8˂�r�^\]����h���l� ��۷P�nW6d�wm	/(�t�d]<�#���H���<.c�g����}�nb��=���/���=�v�v�h��=��9��U�	��w~�������n���������k=�U��A�n9���^L��;nņ5�'�_�|�wԙ����f�ND�,K�����r%�bX�w���r%�bX�g����%�bX�mj�[\�����lP�RQ1D̔T�f�ӑ,K���ߦӐlK��?{ٴ�Kı>�z�9ı,Vfߋk�P5P5�/OHO��1U[sSiȖ%�b}����r%�bX�w]=v��`ؖ'��ߦӑ,K���ߦӑ,K�������H[��k5��r%�bX�w]=v��bX�k3oŵ���������5P%�!�?k��ٴ�Kı;����3��XaufL���9ı,O߻�M�"X�%���ߦӑ,KĿ~����Kı>���9ı,O��w���Wl��[��$��'G�yz���X�Ⱍ.�nggmt/i�2ۏ/[����}ı,K�{�[ND�,K����ӑ,K���w��,K������r%�bX�g�z��l��E&�j浭�"X�%��~��i�b;�!��5�i*):�U���H��ȟD�7���ND�,K���M�"X�%�w��ӑFı,N��	�8�T)�4PD��\��������iȖ%�b~���m9���Dȗ������bX�'����m9ı,Ow��OkSi�SD��ͧ"X�%���ߦӑ,KĽｭ�"X�%��w�ͧ"X�؝ͧ"X�%����f���̷K.�SiȖ%�b^���ӑ,K����m9ı,N�^�fӑ,K�����iȖ%�b|~��!9�a���R�e����u\0\�sr�xzuɛ�8����i.u���{������*5�������ow���~fӑ,K��u��m9ı,O���6�# �&D�,K�kiȖ%�b{^��	r��V,�kY��Kı;�{=�ND�,K�{�M�"X�%�{�{[ND�,K��}�NAlK���޹�9l�8]Y���k6��bX�'���6��bX�%�}�m9��6�Q��~ѳ*hWh�"��L�5���!.ք�sG����`T� C+��2� ��A�� .g� ��>$)�*`���kā	��ԲE�#���� `�Ea},���#6P�#�)�� �k�%n���4CW�?T�u桑���"R0"1R N���d�e����f��h�!��P@� ��h��h����(��>l�TF�����Ȉ��&�ꊟ��lx�S�}�?f�{6��bX�'�׳ٴ�Kı=�t���5�4Kdֳ56��bX�'}�z�9ı,O���m9ı,O�׳ٴ�Kı>�w����@�b���P�I4�MUj�9ı,O���m9ı,�u��m9ı,O���m9��DȞ�����r%�bX� t���),�h�9w����Z�����7X(�3�d79�[2���^;vӣ��{"Jo�w�=�yAԄ�k}O�mpj�j�}��,K�׽v<�bX�'��}v��bX�'��o'���4։��\�fӑ,K�����iȖ%�bw�ߦӑ,K��=�fӑ,K���{=�ND�,K���z�5��5.�f�ӑ,K�ｿM�"X�%��{�ͧ"X�%����{6��bX�'w~�ND�,K���d�&[�Y����r%�bX�g���r%�bX���z�9ı,N���6��bX� �����6��bX�'}��=	�J[��V浴�Kı;�x��r%�bX����m9ı,N�^��r%�bX��w��r%�bX��<HJzg5�.��mv�ٕ8z�k����fv4�j�s�'ld�IBg�F�(t�0kb2�������K���ND�,K�׽v��bX�%��m9ı,N�^=v��bX�'����5�����Iu�ND�,K�׽v��bX�%��m9ı,N�^=v��bX�'}�p�r%�bX�����f�L��ueֵv��bX�%��m9ı,N�^=v��bX�'}�p�r%�bX�����Kı=ޞ3!8h�5�54Mf���Kı;�x��r%�bX���p�r%�bX�����Kı/�w��r%�bX��i���\1��MML�5v��bX�'{�6��bX��o���>�bX�'�{�ٴ�Kı;�x��r%�bX���x���8�aP�&"V�1@�B�����dV
'�6��c��ܛŞ�֑��ƽ�r ��fq�92W�����l
��-v:�f�ab��KՍ��ݢMϞ����=���0]Fx9�=d�ǀ�c������/e�Ŷ�q5k=�3�\r�6�%Lg�G=h�+b̜;�mk�j�Ǳa� ��=��t6��v�a�rַ�i�xF3ݨp�Ջ6�^E{�usה��]/􍘍�d�[I��������ю��t���ݞ�0+�=�j�n��nҭьv�wp\Av����D�u��S�,K�������Kı=���iȖ%�bw����Kı=����Kı>3�|a��ܖkVe���ND�,K���6���c�2%��kg�ӑ,K���ߦӑ,K���]�"X�%����_FfR����&�WiȖ%�bw����Kı>�w��K�AHdL���]�"X�%������r%�bX���e��e�$��3.�]�"X�%��{�M�"X�%��k޻ND�,K��}�ND�,K�׏]�"TȖ'���.�˙TMM��j�k�W�E��,K��;�fӑ,K����iȖ%�b}���iȖ%�b~�\�u��5��9#Λm�֧�ɺ�nI���s��!y�:[��ݐ��G�9ı,O���m9ı,N�^=v��bX�'���6��bX�'}�z�9ı,O~���'��榵.k6��bX�'}��NB���'౯�Q��Ȗ'7��M�"X�%���z�9ı,O���m9ı,W�U�O��r��E
����@�}���iȖ%�bw���ӑ,K��;�fӑ,K��{�ND�,K�ޱG�������*f�k�P5 �bw���pI���͉ �'���pI�>�w��Kı>3�|a��\�3V幚�ND�,K��}�ND�,K���m9ı,O���m9ı,N�^��r%�bX���Y
w��#p�َ�?����<?*�=]6��pi˳��@�ӳ?��;��Hp����%�b{����ӑ,K���ߦӑ,K���]�"X�%��w�ͧ"X�%��{}m��e�$��34k[ND�,K��~�ND�,K�׽v��bX�'���6��bX�'}���r%�bX��z�֜3,ԆYu���Kı;�{�iȖ%�b}��iȖ:Ey	詭�bg����Kı;�w�iȖ%�b~�l/*��&�"�&�����@�w;�fӑ,K��o�iȖ%�b}�w�iȖ%�bw���ӑ,K���.BpѪkNjkR�iȖ%�bw�7��Kı>���Kı;�{�iȖ%�b}�w�iȖ%�c�~{���f$Y�\�j��R�1y�'3XۜX�n�3�kv��v��]�ɩ�֤�ɔ�N'�,K���w�iȖ%�bw���ӑ,K����ב,K��o�iȖ%�bx��뙭K��5,��]�"X�%��k޻ND�,K�뾻ND�,K��M��O�H�@�z��[\�����|����2f��s5v��bX�'��}v��bX�'}�~�ND�����ӑ,K���]�"X�%�����HK�Jj�2�Y���Kű;���r%�bX�w]��r%�bX�����K�臈��N�=��r%�bX�����-��%ՙ��56��bX�'��}v��bX�'}�z�9ı,O����9ı,N���6��bX�'y=�Ir�Ė�4OIv���o��1ώ��C���ȏ��:\e9'�+�/�$�]j�9ı,N�^��r%�bX�w]��r%�bX����l?��DȖ%������r%�bX��ש�kZ�KsD�M�j�9ı,O����9��H�{��[\�����{��Kı;�{�iȟ�S"X����\�pѪf���չ���Kı=����v��bX�'��}v��bX�'}�z�9ı,O����9ı,O~��a}�fkSV乆�ӑ,K����ӑ,K���]�"X�%��u�]�"X��ʺ����iȖ%�b����3SY�pԳ.j�9ı,N�^��r%�bXG�����%�bX�����v��bX�'��}v��bX�&ǱU0k >�;w{߮����S��5�ۗ9�@�<��PoWlWX.^ޮ��h�n�s�(q�8�3�E�?v�hn+m��ݬ�#���W���v�݌9��K��Bz �m�8�nŠ.��^�KE�'	�n���t�չ���١]�tX��qκ�Ƌ��m�Pe,cB�Ìl�U]IFnyx��Ȫ���= ��\�>��PήHU��#�ɩ{v֮�$�X�n*�$����{�����{�7bN��ݞ��λW^/m�v�1�<�^�9W��!���s~{������.&j\�3Wi�ı,O{]��ND�,K���ӑ,K����ӑ,K���]�"X�%�����HK�Jj�2�Y���Kı;�nz�9�X�DȖ'�k��iȖ%�b{�_��iȖ%�b}�w�iȍ�bX���Yyl�).�ə�M]�"X�%��u�]�"X�%��k޻ND�,K�뾻ND�,�dOr]�"X�%��k��e֝��fYu���K�K���6��bX�'��}v��bX�'}��]�"X��$S"~���v��������US��D��3T[\�bX�'��}v��bX�'}��]�"X�%��u�]�"X�%��{~�ND�,K��nR�WS3h�Y�k)���=���-�u�E�V�9����=mkų+�{�Z5fSf�S4榵nj�9ı,N�۞�ND�,K�뾻ND�,K���6�"X�%��w�ͧ"X�%���׌.z�I5�5reɫ��Kı>���>E0C�
�O"r%��{|�ND�,K��{6��bX�'}��]� ��bX�=�zh�]fe�R̹���Kı;�o�iȖ%�b}��iȖ%�bw����r%�bX�w]��r%�bX�a���e�	�5.KsSiȖ%�'���6��bX�'}��]�"X�%��u�]�"X�-��{~�ND�,K��oА�E)��e&�WiȖ%�bw����r%�bX"������%�bX������r%�bX�w]��r%�bX����|�����Z�ۮ�\s�]<9;7��ݰ^�7OWg���n!E�3��k�1�`N�gfkSWiȖ%�b}���iȖ%�bw�ߦӑ,K����ӑ,K�ｹ��Kı;��{3Y�E��	��jm9ı,N����r	bX�'���6��bX�'}��]�"X�%��{�M�"%�b~��O�d%��d&��jm9ı,O���m9ı,N�۞�ND��S��I��EZ��ND�����Kı=���M�"X�%��?w��SF�S4d��\�m9ĳ�`��ܟ�iȖ%�b~���6��bX�'}��m9İ?�H�W���\�����U�'�S ��jd�f�ӑ,K���ߦӑ,K�;�o�iȖ%�b}��iȖ%�bw�7��Kı;�OR{
MPv��Z�:}�ٲ���l6E�qJ��G;!��/3���}�i֗/Y���w�%�bX�����Kı>��ٴ�Kı;���r%�bX�w���r%�bX�a���e��jܷ3WiȖ%�b}��i� 2&D�=��o�m9ı,O����ӑ,K���]�"X�%�����HK���C2����r%�bX���=v��bX�'���6��c��Tș�����ND�,K�{�ٴ�Kı?{��%�ܤ��&f�5v��bX��'���6��bX�'}�z�9ı,O���m9İ7��|�B@��A���n�X��~��ND�,K�맳Z�:.���&�Y���Kı;�{�iȖ%�a������}ı,On]�"X�%��{�M�"X�%����n�n��L��є�XK.z���%@�/[XT�̇d3^oc�f�\�9$�{f��j��j�9ı,O���m9ı,N�۞�ND�,K��~�@�Kı;�{�iȖ%�bx����TѣT�5rk5v��bX�'}��]� �%�b}���iȖ%�bw���ӑ,K����ӑ?�ʙ���5�e�����52fa���Kı?{���ND�,K�׽v��b�%��u�]�"X�%��kǮӑ,K���]��ɩ�����356��bY��2'����v��bX�'�k��iȖ%�bw����r%�`؟w���r%�bX�a��3�e̔�[�s5v��bX�'��}v��bX�'}��ND�,K��~�ND�,K�׽v��bX�'�/�Ck ](`H� +�.��(��bD�!�i�kJMt��&?(f�qr@�~���A	@"��ʜT�9�M #)*��l�!)Q�zۥ,GdQ:�j�T�c�8��x�D�R�!$T�@�6~@�;���ʦ1 XY�"Oˣ��X8�u~���M�b�$����*� �H"t0�2A�U�~���MH�v�l�y݊�l�"��~Hă'�;�m�h��"���,U�Xwn�A����
�,*�U[�m��� h[Cm�m,���z�wlY�v�8��TJ�#V�M[�m=�	��R�y�N�N�g��q�9�'�պp��l$Y.��-of��nڹ�B�M�u�Y�]��ʳc�0�lY�ġԼ��LW&�6p=ed;Y���s�%ΰe�]����֙�I�Rmn类�	ɥqC��^6�R�dztT��g��#OG���En�����Q�,��/�G�S�y���V���eX5�L�d2�j
Ÿ_/����;v�Om�m�S�q7[j{E�J�`�X�\l5�a^��b^\��EƮ�6�4i�Ntb�N��VF��6�۰s���GD����D�ь��F�i�<tA�lV���{q��T�����Xu�-<�eڗ6�kp�c����l���<Ó�Z��͌U�#8�n3u��J�I�u:�	Geඕ���k��|9g�ܮŞ6��a1Zۅ��ɹ�2[��m�<���0�v�M�����
I-Cv�;���ͤ�+˓����	�Z�˻0i��M�3/n�;
����G�v:��-z�e����tM�K:�Nu6:���I�Xc��%D1.���V���E�y[i�v����vT����Y9����Wj�%p�H�m7TK�[UV�@dV�1���b�mD�kʀ�U� ���T�y�[j����n�bd�M����d���D��i	��
;kIv���,���<v�Y�n;hN�W2\�[�����['N�Sn�l������m	ё��Hk���6�
Ą��Pt�P�g�WUi�]ȾW�b�<<��Lk��n���{\��M%��Ei�ۑ���<�[�qY�k�|�=��̚i$:�X�G8ٶ$ڶ�h6ۖ�E����5p��O\�J:�gW��])��s5���� P!�0��\sک��`"޳τS��k�nqs˻���
���s�@/���P�*��^WB�ga���b�3E��D13!�"�!����T� ��Tb!���WK�S�pS��hO��/�P^�!m�ۭ�n\I[3$Y���x��W�a!Ҏ�Erj�����Z]��<u��m�f��ͧ���ȳ��v8秷+m��qApS�t�헔��=�c�.���Z�@��͔�N�g�<>w�)�d�����K��wd���G<�Z��ԧd�nv���4m\Bcs�a�|R�G�Tv;C�g�&�����Zē��]պ�p�����v��øz�tg�3Ve�B(��������YN�u���Ҏ��ݗh�ne'��uIooiu��s��\�$%�K��L�Mf���,K���^=v��bX�'���6��bX�'}�z�?�}"X�'�k��iȖ%�Y��LȂ"a�PI3TT[\��b}���iȖ%�bw���ӑ,K����ӑ,K����iȟ�ș�����5�Ӣ躰�k5��ND�,K�����ND�,K�뾻ND�,K�׏]�"X�%��{�M�"X�%����<k5�,�&�����r%�������/�#R5^��_E��,K���o�m9ı,N�^��r5P5^S���E*EJJ�"���ı,N�^=v��bX�'���6��bX�'}�z�9ı,O���m9ı,O��������0����.�G\u���T	�=�7�{���G9ݶ,1�8圪��T�$R(�fUG��@�g����Kı;�{�iȖ%�b}���a�"O�dK�������K�@����|T�T�
j$��-�@�D�;�{�i�~i�,�laZ�/S�UU�"r%��o~�ND�,K�kǮӑ,K���ߦӑ?�*dK���I���)��V�j�9ı,O����ӑ,K����iȖ%�b}���iȖ%�bw���ӑ,K���oА��K��3).�6��bY��2'���]�"X�%������r%�bX�����K��>�w��Kı=��[�e�YufL�ѫ��Kı>�w��Kİ�B��z�>�bX�'���6��bX�'���ND�,K��Iw}5�k��흑�T�N�b�	���z���8���Gt�u��t�]�3�=���ӣ	���{�T��"�>o!�7n��r� �����:���1���MG��t�����TZ��4�:_v�1VVQ��IQ$U��ذ9�ZY)���ZlJT&��-c���ذ3v��322\jF�a&co"�<��-v���M�r��/�c��,q1��7m��7���*-�{��<�{W��^�LL �9:��-������-����j�WQ9����͞�ew�@���4��Z��+�	.E�N̅b���Wj��hۦ�r�#���"�?w���URC�8ZZ!+\"˻�Š|�C@n�ZNUs��]�L�{����;��;̼�VZ˫\2�0��9T����y�tօ�W=�1�~΢#���k��nI����1�D�qhwJh�lX̭,�݋��mug��D(�9w�/VEu�M�t=;s��d)�W��n6{�L�-�J�O�N�M�Ъ�!MR
�"��?��Z�Қ�ՠy�)�wr�q���HU"�&eTX̭/��M��I͞���O�.ɞ4ɗ�鵋�*�\��5L���Ł���ϛI��3�G��=�����ptx��(&�9�ZXݩذ9��I�ۍ��Ɓ�}>00�!F������X��9��n֖3+K[�4���HOΕ2�[3%�rBّ�k3UÜ����鶍қ��[���8p:�=]d|F�܋�l���Ƙ� ���f�3q�k��g�����vF�0N�8:]�0nbiz��W�7XDr7Jƻklu�����x�y�B���֗�-�Nf"P^8yƂ{���3�ZՑ�u��ؑ��<��%h8�<��l�͹�d�D�����<�/Ge�S�Z�훪k���0w����Sv���kY��Mm�ba�[��r�v��rZ��#�2�ZH˻F�N,PiA	5�Q�Gyߖ���,fV�$�Ͷ�]��}S�X�_MG?H҃XF�Z[)�߳��ďm�\ˋ@���[�W+�Ď�j��Ue��!��gƁ�X���ߒ�� �ZX���R��%�m��m���ύ���<��h�d��$���E����;ܭ,&�[�_��}>4z�V�x}X�$m��f<sxc;.S���f-���RVC=������`VD�od"M�@�e4=���jv>i$�I���WŁ����?L2A��V��ܓ�w]���|SB�D�K�S�`s�ZX�Z_��S'�����%6�R��?�{�Jh�.�S@��)�yy%M�_��$�-W�UV���@���4�<f��ymh�.�$s�G�`��-��߳>��~�eŠ}�q���!b�A���Q��=��Nݦ��� ��$�@���9�Y.6�*��g�uḿ+~�߿��������>���s��92���e*B��
b��;�S�&�Qg�Ŝj#}�����W��m%�Jd߼W�TU,l$�$�MŠ[�?���i������	���I������ح,Y�R�j�]��������H��d4��3C�]��h.�R���uwu����h|���rV����hv��=]��\'��)�8�ĴB4s�F3�Vub���r�=�d#��fx�v���m�? 䬆����u�k�U�{2Ѥ����`��yY�������4ڈ7��E����`f�/ͯ�w`�K=�������E�f���@��)�u�)�yzS@����E^$�3��%U[��vVC@������$Jf$�iq6���_"����R�IT��TUn������Mw������yh�����k��X�eԮ�!��wsK^8��՞�rd���� U��+�J,��c��ƂL"LK4/Jhv��;�q���r� rVC@t�˫>N&񷐃nWj�;ޔ�:�lXܭ/�_6�jd���ȟ��Su�Į�h��u����_G�����x� Yt��
��,�C�Uʮ'&�hG��:��s����-ߪK�X���Q��$Qh^��>��I&�������}f�lX��d5�!�Y�IL��Lu����fh�nD�]�mWpV�|p�;N��Q���Xʶܦ1�A�d�����8�0��63v�z$zL�z�1	�n��b�<d�'��o{tn��mOFl6S�[tpg��4]���N�7/m��C�]�mu,��Z_8Wn`�tM�noM���tN;]�������â��x���]�A�cf(R*��R�U$Ъ"*��Eq�i6���Z>��>�	L�k-.MDu��K�,�g@gI{5�Ϯ]�]ϓC��D�L�'�����{'=vsb��ڍ��m��~��@�O��Ŏ(�q$�@�_Z�$71E�}C@�����s��)u��2L�2L�)ߢ�h^��=��S�"���h>���^*��b��Zű#���"�;�q��Us���-�&dW�������:�V������b�@����{���˻x�wj�Fn��ݦ��\�0pl�;�Q݃�'J�=��|}�}��<.bqx�>4�Z��4�ՠ_l� (�G�X�!�wX��g�`�5iE-T�1KBP�",8���_*���_����ȴ��f���>�%5R��Jř���y��Zz�UI>���o�|���v(���k䆁�;�`gr��36�b���M�Ͻϋ}qz��Ҭ/-P�"�1h�����s�T���>�!�u�k@�|�T�,-z��E�9�����}ALD�9��Q0q�n�q B�������}��\]�t6x�E��<�)�uv��빠{x�7x�L"o�Z��7�߿$_��@}sk�����-�&dW��IE3E�������ڳ�Z���v�h X�)�;J�f�I�M~b�	"5iF9���5�@���3dc (E	� ��*��`����bcʡ��ʴ��{�I��	��]��(���{R$�$�bp@�Bi#���1�$b�C�$�&����a>�ic'��N�ئ@!h�>B�Ұ���S�N&��|�������DQv���'4;
=�7�����r,�֖!tQ��%Dժ�J̻�М�9ˎ{��<�/-��S@�۹�_l� (�F�X��hܨذ>i��Ͻώ�}�}V36Ն���q����,Rm�:�n�[�I�iӿ~�N�u|�l���r��҅��� �^<H1�^��@�۹�y�w?�3<A�X�Z֦��9�F(��9!�_m���+�76�	׊-�{��W*�;-��qb�8�	��h�����U�y��/��h���2cP����+4ҏf�z,�Ł�ݵ`�t�!�DRM�qN&�NO߻�rNw���cŒax&��<�)�_mܰ;���vc6l�{��"�Ttm�Ɏ�z��V;i/J��ȹ6�y\v7H㵃\Q��6ݫ&�%̄T�%L�7�X��V;1�63kK���D�*&H����iX��W��mDɍ��9��?|���� ��(e�X�*����Vrc}63kK>i����{֬�����)Vo�L�����Q����;�����j���i�͸�Ӡ�E�2�9yb�j���4���&��������ͭ,*BMo{�'$"��
`���	�3&*b!w=�����6��]�C;#�;E]9�<�q��9N:z�C�c����F�^ܛv]6�r:�����Ge�8�=�b�y�����9ε�8�J,8-U�l�Sfm��s*��ڴ�dǥ�=�x��c`�\lP�70��;�m�����a��g�Ʒ�pL��#�6����Yգf�I�1�z�m�>�=r�zí��Ew�����ug�=\��6�u���W��r��
�:#l�G���L��U����{����q�d��/vd4�i��>��z��ˑhb�b�&Lj'�jנ{�Zy&� 3��E����~m���4ۙ񞫫�*�Ve��k2�=�4���u͇�:�Iz}L�U��%���L�6�n7���3}�Vrcvtz�h��.���lL�����[��'+��W^)/�s!�|�7���Gv��<���M��͑�,�-�mmnb�Nع냟96�l�z�����b�<r�]�hv�w�}׌�>v��s��6� �E�Z�Ŗ��v�/@������2 ܕ���;����.�{��s@��j�jvI#�㉍�yxh7��>�{ZJ�W8�]�/@��w��	ɏ�X%
C@�s@��������R��~�Ru*s2��a�X`���Z�ݓa��&��n��5q,TNĤ���m�
:�&ݪ��r� ��vzu�����cXf=�=�C��L�`����)�y�u��Us��}��Z�	�\Wv�!]a�n�۹�w[��y����e7��:��ap�Wi�a�yZrmh�9�`�(hJwv��;���{�He],.�]�]�hNR�����d4�7���M�����,��Z\$�Ye��7��'ݓ�~�6��Z��4���x��Q"�rDʙ�:�k�.CmI��ų�Ƣ��.�ͧF�K߷��}��I�Lx�����s@�s@�ֺ���h�츜x��(�������H����Kqh�ok}ʪH�ϳ��dơ?(A73@���=�ִ�)/�&ց#�Z�uc�Fb�.�2&�z���<�S@�������`Fh���%�,&�5�Q1�汽�lz����(S虘��%QS1����4s�#���v����ZI�)��z�o0�a5LԸe�CS5|���Ӽ���.{�8Gm�z��s��.͞���$sk@����@n�Ԫ�W>�～4���� �<Px��&�h�]^�����x����|��.�%~k6�P�w�w> ����5�= ��nG��G�iŠyl������}��ք�&�Š4�"⫤�o�i�h[w4x}V����������	&�o��;j@;��]�'E:�Jە��ڻj�n�T�K��%1�6�V��&7��&���\�x�:)E��8�)psb۞�Cݣ;�����`��n%�u���\� .x���aoI�sc�][�#C�{q;5���4v��b�9쾮�u��v�GSk�� n��G��Z8�z�v�@=�k��s�	���Z�F�=��yP��������~��}���֎�gݨ��X��Z���:s��m��}�q�;�>{;0�u�3�;��7�&Lj�i��h��@�}V�岚�������8�,�"Mr-��Z��h[w4x}V�~�UU�ڄ®�����Yv���{<h�{Zz��Yn-�qh*�]��]+�V`�J�Е\�UU���ՠ8\��;�U�yl��yz�Ŋ6�nf����;�U�yl���s@��P,��1A��?̄��Jl�v�z�+V�v�]}�v'��˱|�)��#��-w�yl���s@���h�V�G��Ǐ�@��M��ݯ&��7���N�,�͛;���m��M��n�������M7/@�L����tцVRXi��˙�~A����g}7��'����-��<��hڶbx�L<rBI��#3f��6��6�Ͼ��@Ͼ�Ձ�'6,���z%ETQ2T�p�Rn�1���°qu�씝u�n��cg�o�N4�n3x�&�x�r? ��Ɓ�s@���h���=\~��'�2	�<4ͽ��r�UT�i�疁���r��۸%1�ō����{��$�~�ni�%���?��i
��q���3���Hh��4��O�6�q���Ł��Z�3�Z���#�@��^�岚����%4ӫ��c�G����������O�I5�}�W@���r�@���V��0�'���Y7j��ڪ;v�NB��ڑ��/��d�q�mS��m��M� ����/RS@�ٳ�i��{����yTR�EE8�-]�h��o��]�c��I2����W9I�t��b�Uxe�^M��x�=��9Uľ�mh�!�{�q<����!�z�S@�۪��Ҵ��4��C�I(bI�CK@���y��7$�G�&{,�bdp�<��h�)�r�@��h�{���.	�yML����������ai�1tt{`\��d����2�ݱsŮ�]�]�~8d4�]��g���s�	��b�
��-
���0�?�R��	&C@o�k@}f3}\�q d�]̵��̻�V���I�����/RS@��z��BH�"F�Yj��W9�#��@���z�i�?}�>,Q��QR�R"��QDLҰY��}w�6�}{Z�H�������h����S�̀UVR~�d"�=%���|F��M)�ȩ�>CBD��$H	��P����9�B����+i $v��_����ր��AӴBo��� 8�����?8IjI����<�ȷZ�v�kHt����������,��]66ٷl �i0����oP��۰�]6=e���Q�r\i��H�R�n�fg-�vE�{�)�\�Ҫ��%c�t�-�$��G\�ڠ�q3\��M�����.�z8��ulI���Kg�S�Pm�%����җD��v�Ò�莈�g�˃4�1"+&
Bj ��U[U��ܹQ%E8�pvw+<fa;`j5F�ƹ�c,�R�۵8���;W/��e�G4r`��.�N�ktU�0H4Hl-8��g��]��d��1Ԙ�i	��c<kfX��8�{e⶞ F퍮T�5����];۶7H��a�Y2���n����'�[.�WOlZ3V�A�G��x%���p���#�y��]Y @3��+J���u�A�6㋉۞YHe�l��4o;f��q�LGi��N�Sݮ��u�Fv�㗒`�"�CV�<Á�a[n�%���J�VG�mt�	�uΌ�UN��ys�xk��Ä���pKl#� ����ٞݪ�k��F�$`�\��c�d-pU/-��s���u��;L�Lٷ�DU�ve87F�;7K-�'
��$�j�	c�<]O�M
�C�tv���r�d�8M�c�ݶA�� b����*��mF4V�H�Q�Y`^Zڪ�,���ͱ��S�5^�`A���Ԫ�����
�]�4�ę:Y@n۱���$�j�[��9����q�C9(q�r;v��6�nX�ᦗtW6�D�2]�;`���jWs�z����M���9痘�R��,0��W����q�`W��1J��wcD�ε��A��J�LiQ��CK�cj���;���ݳ��M��G�.�vϟ��vxj3&�ƍ9MA��.�m�U-�{O50K����z3��ݕ:N	L��3�0l����`�m���A�1v�9:�@�n����,<t�c�d:d6�.��W\��9'h0��:��)��:��W�6j�Η��Yu.f�.���c������"~@�E�ؠ~E
����DX�� :��UИ�
��z{�3�ch�����'!2G?Oչi�Ұ����(��#5M[��N k�<�:�6�#l���ڃm�=N�۪�;v���.ay�u�4c���7a����gq�a��a9g�Ƥx;t���7I��.\����&�'6�
��i�j�/6fs�;M�[l!&����
4h����J=;�wb�nl�r힥^mX�m����ƪ0w��y�����X��Ok�l;�7@��zz�Q���ipR9�9��U7��]i�u�O$;�eMGwf�ݝذ7sm|�_6�d=<g�:�W^V�`+�3̽�j�-빠^���U���٘���2XZ��һ0V+�Z�mh��h^�@�ڴ���0J0y���s���(���kA{�Ur9�h�b�
��+V^a�h>��=ʓ$_��ͭ���r��/���˷aܖ�(��5q較��^�o3���9�v���h�a;������S��x�.��޿yh��h��z��_�E�@��}�9"F�D��-޻��k�4�\M�]E�;Qذ;͛vwV����.�F]eeqa����$�E�Uz��j�-빠{m5�cQcŎD�	��
�W�Z�Z�w4')G5E�>�2�"�����2�̽�mh�W*��s��	(��]��?�������ձ�vT���y�b&�4��f.�kg��;czH��G�����w����u�X��|�=��>�Mh>��v����G�6������*�^�yڴz�o��E�jD�)&���=�M��;�d�ڄ�b��B�@0?D1R���")IQ)���'I!�j�'o{j�����0��%P)���
`�����_!&�޺�X��k@m�4%r��~�O^�߱z��2��JC@���m��*�^�m��/r#���I�d�,��?,nv�GM�l�άcF'=;W��i
˒�}��OWj�Y��w��	&C@i�ހ��z���$sk@��uvZ��p�ŗI^O��r�$�G6��3}ćڂ�DW��J���^�$�h��i�W9�JI��"�^��W�;N��WY�bN�w4l��W��2��۟���7;����m-��)�"f�@��h^�@��h���:�.�7��Rm��n���������۶�?[��=]��ܒ+pE�k	n��c����9zo�7׵���L�����qDc�,Y1Ǡ[e4�w4�3@�}w�ʮr�Uv7�U�3^Z���4	���M���Us�ʤ��^�$�h�}x,2��YVbĮ�'�a�5��mhJ��.z{��?��#�����7�8h�W�W*����sk@m�4U\9(�RK�!&����
C�DS&b(*f������s�֎�i�Br�:,-�nz��h�'����!�{9ŵ�`��7v�2�Lvs�l֋m�wV�O�s�y6������˄z�����Uc#��*>]�[��"Si׎5�&.�:�=���d�$�3mm8ŗm���Vޫ�����mq.66��qg3p�l���a�Dե����z۷\�9椺W]���lu=�F0�����ߴ�O��t�e:4�rfrLx�)���k=��\��\��9`.<u%��Ơ��r?����Z^���S��� ����=Y�|���'��	����w4l����z�ՠy�LP�፡73@�e4
�W��
;�h9��w��P�.b�"���4�]��#��#�ZQ͆����_8�1ƣ�!���ՠ[�s@}x���z�\���Kn��WG;�v=���чՅ�.�;����ӝ�#V�̳������q�Q5^������4�]���Gr-�\��b�U����&iX�Z]�Ɣ4�$�$�J�W�y�ՠ[�s@��񱪱���Wt+�@i�ހ�m�=^�r�ޞ��?���Ɓ��h+�@X�r=�h���/YM���,�+���t]^%b�Š7׵�J�+��~������@�b�OZ�x�B��2)����[���'=ps�<��(=u�z!�a�F4G�6������*�^�yڴz�h�"U���h>��ʪ�U$Gr-G6�׌�9UqW#K��o��@��Z�m�-[R�hP�BI���Z�FJƣ��m&�>�W��ٰ3�Q�5R���b���C�\�s��s�h̆�U���ՠyG�
D�bB(&�h���U���ՠ[�s@�q?�w�l�+��d-q֞=�����(�bݭÜ�Y�sWU�,�<�!7�xfL��RD�' �}~z�j�-빠^��{�Q��%�������j�i6�L��P�W� �rk撈9
�e�< ���@����/YM����ՠy��0ʣ(���ۊ��'�m���}ϋ��}6��ņ�����)k�RwW;�`gp���$Hc�C@�ޯ@��Z���z�,�i��5z�*4I5�J;]�E��u��6R�q;i3&s[gDsi�uf���������9#x�!8�������]������˯�@��_B8�r6�PJ8��]����*���/;V��UT�����f+�H��w��G���*���/;V�}빠[�x��X��Ȕ�U�W�^v���sBs�ʥ�h�Ae���`��3̛rwb���ڰ76��6;�6[O3��J̆	4�8G�RE �M�V��Ƚ�R��;U�l�ɺ�f�m�E�W$4l�kVqi� � 9����Iݹ�۶�+��^�53����c�;�V�������2�F
n�F�ͨ�l[Ɯ/K,�3��x��8%��AvKf�zvf�4lۏ�v۟�q��s�+!��hG�<���uv´u�t�맞l��p�l����7^İBA���;/2m[��8��]��=�Տ�n�	�{<��l��;\�!BB]�2����8�8�ژ�G��G>�r�u�����$�k@}x���~�s���;�hveB�X�K.�V�^V���]n��mh��o�U��ClX�B���ċ/30�"r^��m�'+�5�m9���֬��|X�(ٚS
UR�x���/;V�z�����*�^��ؓ��H�h�QŠ^�s@�UW�UU^����S޽��Z�����mn����sO�&�[EǍm�-����>y;1B^8Ύ��8��:�l7|�w4
�נ^v�����G��UcXD�	�@��{��4Ş�&"|
*����g�g�]�>�}��>�f��ʪHl�˥d��R��b�Zw"�:���W�d4.E�r2B�1*&J"H�������S����=�g��mh�k@�ה�bHQቬI��-����4]�@���h�T�Q"��2��X,\"N,��^y���1�\s��q�q���l>ѻ��{��~��x�DĆ7$=���4]�@�޻��)��b��kH��F�,ͭ,�6Ձ������l_�I���?�D�H�iA%!�{�����,���4�c�%�H5#��hM��2���BԫS�%�+4 Cz�CtH�Z
��H��!�>�Nh��!w��,�@�&�j@��[�Ԝy7�r�UJ�,6h�;a(E��D"pD�f�������	SA� ́��>7�h��V
Aݡ���<R�,,"0�hRܔ�i.�ځMi~R�q2����<�|�u�;��ih0�Cʈ�A��"��\/1��q�����>o!���(�r�����Xb�J�&C@������4=����~�FG��汿ÑF��y���S@��^ց���RR��b��ˠ���N��rng)�m�.�d�tG<�� ��']��x�HX��E"����@�޻Z[�Ns�U��]�-���b�U���Ĝ4=빠u�����@����}�)�(�xbks4z�h��3Iĺ�C@��mo�#��z�+P�$�$���É��������x�9��V}��C%���\i��>��,憎���x�yp�=�)��^�u�~��9��~��� ��̵��/���`m�;�ęM�d�+v��i0�<�`�^9��D�I	#m�JC@�޻��e4=�M޲��>wG�U�,��+@����Iu�4�C@�޻���ZG����L��i8h��u��<�����x�<+Y�2���s����>�Z��hz������\i�x�L����ڰ>i&����;�76��3�~P�ĩ��4L-Y6n�4*Y�C-����H[�̹�c������^Z�=)���w9v��'���.7��)���+�D�k������"�ۊNP�v�J�<"ݷ�6rmG-mi6^7���D�Ô�[[�ۆ�tY,kV�Y����7�nd��Y�����@�����ڢ4�L��˻-7bu��>�d�y��\"'j����x�	�\����Jy祎��� �6��LP���W��JM39Enݛ��}���>����k�dt�/c�d��t��ې���Yu� �HYtUڤ�*=��~��Ł������s}j��o�n��bC����������;���*D�<qE��ㆁ�;�j�4�Q��������v�d�$m4C��<����n��)�{l��n�5�cB(���37mXi�����3ޯskK����?�;��j�f7����Q�Zn���nq�����m�áܹxy��vmi�@������e;�g�ffz�96���Wu00T�f,��@���ޔ�'��-b �v�:�m	4Қ'��{}j��N�X�O�<Yq���	��4z�h��i�W*�Iu܋@���EuhYtU�J�	^�+�˓���=�4��h���=����M/�1!����h�)�u��u��-�IO�w���loW:�Q�j�Ugr��y:��+���{'gmۛMv�;������*�瘎�	5=;�3r��3�Z|�M5����@��/��&�bh�)"�:���\��fC@r�Z����W*��塀�H�X��Xbį0�#�x�:�iQG�$D��)H H+��b�v���y�X�k����R�T�B�bNW�h��hzS@�l���(������Ԓ'��}V�*��=��fC@뾵�z���cT]~+�F�����k�!m���d��#ʅc��6�&81�����ԉ��oC�\��xh���{e4���=���<�̥e�t�諴��~x͞�W.��Z��-����$|�/W1Z\�bC��ߖ���Z^��:������*��bB*�J�����i��i�������WŁ������$4����4R��$F�W�h���(�7� ڈ�fo޻�}����d�d$i%RE�u����]�����u}V�s�Dac�L�0M���z��a#��PȻ�XƌNzwl�l��K���{���kw@J��r~��@��ZW�hl����'�U�ȓp�:�V��}V���h��<�#x�XX��E"�=���9�f��s�竗s�<h��-��Ʈ�\k'�'�ȴ�S@�ҚWj��q9�-��P��]]�v���@��3@�8�H�r����7�q�q 1�t���JjL���0�ă8��7hݵ]��N��;�c1k���b�]��mŔ:�������J�f6Cm��͈砃x�cY�v`���i�0�P8�!�"'�F��u���n��t��64%�L7�j��-v�}���Ch	YnB��_8��\�>S;�l�ʘh���6��
����`�Lq����*�Wm/]���nVɓm]{GkkrF��fZ_=V�ʾP�))-MDM���1�6���!�cc�����W}ݎk��;�H��O�Y�J�e���3��?�@����BW+�	C@�7��eX,�T���Š4��g?���O{k@��x�>v���B��q�&,��$������h����v����\nPXǐ$�h����v����O������_���<�0N�ڴ
�W�w[��[Қ��U�c�@U�q]N�����9{[k��c)������wl�qvH�a$D#lY 1bjI�@��zz�ր�q���ˑh&r]��*��b�l��W��KM&;��3�@\�@i���#�̨QYvUي�V��+@���m�=�J&��ɵ�~}w��.�̻B����Cܥَ-&�������~�@i�,�Jc#X�&�Z]�����h��hg���|�X��Ǒd��=��ހ��#��qՈ�ɨݐ�]̳p<�����ո�H�b#�G�_����c4�����]k=I�r`�V*������2�?yh�������W$pܥt^Yy�X+�@��;{����61b����
�V
D �X"'ɦ�Tג�i�I��{~�`gv�X�#lY`�,MI"�hT+�����4=�W�U�[��-���ؼ�4�J&�z{n�}����Z]����Tm�-�5�B�ɣ)	���`��3���ϝ��|����z!�v�|�@&����e4k�
���;�w4/W�27���crC@������r�Wg���?{k@<f��n
HF0r5��jE�|������h��h�b�#�H�")Sa�M4�s��=��vsb�bc`4�Ʊ'��i$Ӆϫ��l����4Ōy@Nf�}����Z]�����U,Y[��)2��̈́�źx������1Zݺ{SX�;���*_1�&I����ȓp�=���*���;�{S���W��!�8C.�U2�8�"�h{���}�4k���ب4�MD�qǠw��h��4�\��]���"뗠}��e���	�'3@/u���Z^��-���׫27���`�@�}V�U��-��oY�\y�~3��sLI��0� � ��v0�C�XաdJZʈ��qE�8�^��T�j	�	��S>�*�5� v�I)���D�M�t� (	H�!�6 B%�c~6�O������hi�cmS�h���=����b��=l�3���!��"��&t� ?qD�p�
i
:ث�S{������{�~���ą�2�6� ��݅�����:� ��M��d�v�����)� ���,SR������p��fv�Y�8�3I�X����D��v�Ql�u^e�,�G.O6����x�q��$��gD\K��t��f�]B��@D�Zsյ�u�r��n$D�)� ;S��(����n�;c���3�OWnvϥ։��A.��.Q��=X���T,؂Э�Y:�ڇ|:}4�s��
��� �ݝF�j�8)��-�9U+�:^4(��'�څ��J��W� ��DY6�����-�euX#�:�1B�mi�n�]���.h�b�Qr7'nx��y����p��8�e���Q�� �.3m��u��x�x�t��JO�rC��l�\IA�&��\�%����@�獯	�+m����cmۜ��2l���ۭ=,�mחn�-r]p���l�X�;M!tQ��ݙv�^j��ZU��Ggs��nӖK��:��A���lN��R���\c�����,�'��H�����h��5u�{�O���8��g0��A�g�x	�O,]�8͓::2�i�,c�/�ʥUT��D�3)N�ݓCs�=�g.�M����T,m`�;;u�1����r�8jU�����!��RJ�o0[@�l�d��6�b	�)gkAr���z�B�� k��t�/[�Yɴ�<

�g�R����;
�&�;e'r�j!۶9���mϗY�)�sl�nk���2ZjW*\�ֲ�Jږq6�ɰ1+��R��-���M��h&1�RdUɝ9�EB��Z:ݳvL�.��ZzGr�F#8���cF0��۞R��kp+���ݴ�o7��#�&���B���#Q��A�R�D�xa��L	�G��=���la���v���/2T�K�����5�����rp��!;��n��ٵ��sW=�y����>�zɣ�=r��/�f��ְ��bI��gO�5�%�ե���5(�ʠU��SH�0�/ b��4�t�P��uǮ	�: ����~'���A�5!m���[���,6[��[=le-mu���9N�q��+U�3�Z�S"\J��k��q�r��q�n��Y��z*H��;[lV���j�֏=��i�ƛ��')�7n�ssld0��P�u�nG�;�����m;.��m;s�nl;v&yP�O�u���p��M�l�e�:: �����"���U�7K���D���cj\�5sXfIuu���o�P��I~�����7W:�:���c��qc7�F���K�t�D���{-��՝��E�������s@-�4��h��8�d�28�z���ޔ�;��ZO���W+�ʻ=��*�b��(�J�zg���������J(��=��4z�1<q�L�@N{}k@i�ށ�����R=���}@'$R-���ٞ���g�$y	\�~@ݸ���R��Y`]=���.�k����`��^[�p]q�`�6H��铣O��ؠ4�MAA���s@��M��Z]��ה���	��).hܓ�w]��q�tU�4uU�-���w�`z3}67v���i(���=Y�C��LnHh���*�@�۹�_l��U�G! ��1<Mf-	�Rۗ�}$����w�ִ}�X)���E�@�۹�[Қ[)�Uz��9eĿ-n0x��X-̦^q5���������m<�g��R�灆A�ƚF9?�Nf�oJh^3@i���? q�4	7)]^Z�ay�`��u���UI7/@q�4�߱#�>#lY�i �d�8h��M�������_-hW-&�=~�4�����ب4�MB6�z^��-�M�Jh^�@���YeҡZ����4UUr���x����:���r� ��#mb��	�������BLO<.\g��E9{D�dNѻ�mŘ�� Ć9$4�)�Uz��Jh���U�8�`���w���뽜�U$H��!�7Қ{b�R0#Č�9�oJh���޻V�U����ؖ44�38��^a�9\�W�a�5�/@i��nM���AP�X"0� ��T�cA J~O�'���M���ى�b`�Jp�9{k�*�^���Mޔ�.zX�iH���q��ErѮe�#čcv������^�ۆ�z�Z�%ݱ�si獙�S_lUz��Қ�)��@�R���i�Fԏ@����bG�Y���h^�@�'VF<X&�r}�h_^i9T�Q��y���f(��$1�!�z����zS@��4
��FF3 ��$��*�^�ץ4zS@:����C�`C�������I%�AIY1�|_�)��DOK�=T�9��z`��rk�%�
�dڐJm^8�tn��N�zr=9�wk�jzkɸ����d�[mݤ��h��.�ۉi��v3���=�<�FNb1m{>-����]���'�ir��J.���Aʅ��ǰ>��{6���甠q���$�؅��Kە�ݠ�.uf�@���[[��=�i.z[�ў/33_����՟rg��Ѧcm��y�'��Q۫gN��9�vk��s��r��s�4Q`2F�%r?@����h���u���r�P4��C�UʥX�%V�J�O�<NC@��>4�Y�Uz��FlH��r���V���4�3@��z^��-}V�}(�c�x��y�@��z^��-}V��\��s4�!J�U*իV�˵�z^��-}V�u�4
�W�~��.;��k��^��G�}h�q���z�r��G�u�={j^T��!{s1���.x�'f��c����f�W��|A��4-�V(�H��I5UE�f���oRM����n�]���gƁ{�4
��FF3 ��$��*�נu�M?�K�gƀ_��@�lV%"5�(���zS@���h^�@�{k�/�;`��Ҭ��˥y������	����d��JhZ��A��G��&9$�w��E�ū�������gldk!��y�mЌd�uZ�x�X�8E19�u�4���J}�3������Q�c�1�RM��@�Қ�ޯ@:���Ҙ�5A&�j���:�������<��w�No�<@���BKѤ�4�P�w�{9�63=66V����@���h�z� ��h/���{�%�YuFZ�J�+�� ��h/mz^��=^�z���w���m���ԛ�;v�1�lg���s������<'gmۛH�N��0���gZ��^�ץ4W�^�u�4��q���(���zS~H������<^��鎻�Y$�����������K��/@q�4ަ�lq�L"���C���������̭,%=M\6	p�Bz��x@	ZX�%���(Q):� �?//��ӈ�5I�n7����̭,�sf��mi`y6�wƙ��N�Y	��L=w>7b��7/a��]��I�.Snw6ֈg�����[���P���}����z����S@�{k�<���4��h�z����<^����h[^��a�J�+����4���IIG&ց����9wU�&`�A���4�������]�{��(��@��e偉�B"�G�^�s@�{����X��́����RJ]�mV8 <��yۓw2K+\�F����}��u&ӫӛk��/����8v�<�[���(l�u�6@���Z��^v4�]nZ�sˎ\*^r��*��^�����dܘ��:��F�;ns��\㘱�̱ԕ=��K�h���2ufE�jČ#[7J\m��+��-�n�5l��Jg�:��q�	�D���6xIM�����nݞ"
-6����5sE�3F�3D�QO�T ��������"�������p��rJ9�k]��x�9��v�]��W��n;<�����z��Ϟ�zˆ���נ^�s@��ٍ�5���S����h/mz�w4W�^�u+k�Pq����^�z����W�^��{��bx��&�H�C��ߗ�Oՠuu��^:4%/��^��O�ƚ0M�9��ޯ@�e�@�wvl��V/6���Ĥ�!Ǝ�˷Z���
g����������Z'	��x�: �vq��y�k&�n>���a ��s�;�d�����[mƚ�c�Ē�rN_���!��`�Zm��srՁ̜ذ76��Q�i}���,DRH���nh������z��1�. x�p���h���\4����h�6c�Ȱ`���Z[.��z[w4��Z�P�,s
O��0J8���c�^�oD�vX�@�5�	��na��Ƿ-�A��B,�����h+��m��<��h��h��O�!��5#�/[��<��h��h.��+�0��M&Ĝ��}U�����i���3�)-�N\̂o�����adQt0�>�����2IH�XHI�c�xO�#)���E�q�9˳�`Ma���꤀��~���)(B$-?4&��B��X��/�bCc�P��!���# }������H��h ��{ �a�<xp�����	��_�	,��F1W�2���%Y�HH04l
0A��P"�U��1:M�*D�1
D��#vk�BD!����"���)�N)O�MS�!�>��#�^�l�E���X5֛���Fq>1H�A��@������;�GD�C�3?RC��"�"������$�|�~vl!V4eHQ�Ft�N�'�|/�T�:��9�4�O��~)TND ��u�� Gmꁠ?ϟ�L^�Dg?Z����s�Z���T�ꌵJ���x�'9��F��n^���ք�q|�Šr��ܒ6��c��	�4uz����}V��e�@��2��#��n�od���![�G��9�tQ5�͞�mԳ�.�@��-�O�o�����ݾ��w���r�	Ү\@<i��ē��yϪ�;��h.���j��m����JT�P�	����Z�O��;��=��hs��Q��R($��BI��y�f���vx���}w'~$0��R�h�A��10$Q-h ��R�[eD�"��Шt>�����?�lk�� �RM�vՁ̜ذ36��ͫ�`y
=;n?[��v�7Z��H�Fmx�>ϖ�[>�NF��<c��a��݅������Zz�Ѡ�^O�;$��>r^�R�0�b�ҍŠwYp߿~���{o�@�{֬d�����qFo����dD'1��h��4m������ˆ���X��j!��7$��31t��h;qh��F�~�^h��@<$őē��yϪ�;��h��VwvՁ�������2B��,�S�rD�M»�ՠدMY;��]�z��m�\���id!���)�6)}pUÛr��l��{��d�k�km�Ѳcn�-�s;���RkO�����0��^�s=	�M�5����Ʈ�p{�F�����Zlg]��QpIN�����Zm���!�}F�D��ɳ��^�YsU�v��nk�ؕ\W:x�q��Z5�r���� W��>>�m��uuh<���ǉ��99�͢L]n��ٚ���'c�m]�ݐ�\�����?[o���ݾ ���w49�Z�Q7�АHr5	&����w4��Z�\7�����|65�1�AƤz�I��w��ZJ�RRL�h(���]q��ʘ�$�'3@�_U�[e�@�^�@���ε��Q�
,15qh�p�<W��-�s@�_U�{�ٰ^{���m\:v��f����Uiy��</nKZ�����D����I����^�m��z���.��ND��E�@����?�Ȉ`4:�?��T�77���'ޙ(�?'�z�J�qt]����s<�-�.��z��h���ȰdQ�ԋ@�ˆ��^�m������s��o���A�$��=V��m��;��h�pݷ��w����;L�0��ѩ��J�U��vQxoP�u<q*��◈|r�s��q��}��nh��l�h+��eǜ`4��bě�h��l�h+��۹�1#�+٘��Xbj6��-��x�W���`���_Rm�J&=����;�1wt��,s�M�4��m��;��h�p�/tW"���IdQ̽���Wq��	&J4���@�~�������썹�e���L���X�oM��dܡ��f��:9A�ttXNf�篪�-��x���m��=�	q�d@II�H�_eZ���@o�k@���R�� �˫S]��A��E�z�o]��_U�Z�*�=���cU� �=޻�;9�`n�-�M4ƥl��jZ�X'��G&���rOǜ�dˇ���܊��_Z�=�1�_��u�����ߟ�����ߙۿE*qб�	�w;��8��!��Om�����u���0/jk���F�Q���ϖ�����-빠y����l�,s�JdZ�ޯ@o�k@������5���Hm⁙�@V^J����$sk@����"R]ϖ�����=�դH�oE9����@�ˆ�����-�s@��%ǉ�@IH�"�-��x�����V;9�`q��4��И��?�[��s+G6ڙ������nd�y�:����w�hK�q�r�s�9�m۰�,�-=P 5�x��f�����lvAjZ�dv	�<5�:u���Z�m�X��<��Ŷ�3<ڱ�7[k���@�r��G�;B)�xхݒۙ�vf�Bv�C����aۭ�6�92�;H�=��{A����/����H�t��M��g7m�=�GA3,՚�3FR�5rd���b(xz+]%ƚ�I,A�2bf*����R�fSW�d�l�,�H$�����N���i��bG���NAp��$��>V�=�w4=}V�m��wO�lk�,m6BG^�$�Zﯭh�th��w�~a�8�1���b���_U�[e�IUI|���I��~��ܪYuB�E+J7�m���W�[n�ﯪ�;/U�(,@�A����@�{k�+ok@���Zo�+�\_2LJ�ݵv���]n�d;oUG'FIť�2�u��W�W���x�:h�i�U�������M���ִ�:'9��\��W.-[5��f�.�e��s��۲!kRC�+��*%E�E��]S�*��ˢ��>����o������px�!#	�Z�\4�z��w4=}V�u1\xӤX8��h�����h����.���lj�M&�E#�@����_U�[e�@<�٠~�*���=�g�z��/�����rz���<[��v��/loR�7)�ͷ��z�������w�[e�@<�٠[n�綽��<�5�Q��m� ��f�m�����@�VȠ��1����@9�ڰ7wmY	4�]Bm�Bi�Z8I6�ƚ\m�/'y�V������"F)�X�rh۹�{��l�h��4.:�&�ıH��h����.���w4-;�wňN��mm�9."���Im�g#s�hkg��\��)��̎]���N���LjE�[e�@<�٠[n�ﯪ��+�����N)&����E��h����.���65A&�y�rh۹�{���+l�4�ݫ��	�Z�H�� ��a�I6Ҍ��E��z�� �wj�m�-CK[Iѻ���M��)0�	*fj,l�h��4m��=��Z�()���v�玣i9y��n��*�Y6���70-�ն���l9#�ȕ8���-���m���hz���.z��$ȱ
dĖ4ܚ��o٘��;��$�(��u�Ď�ed�1,ʵVb��9��gƁm� �����h�-�wC�0���V�	�)2JZ˯�@����Қhb��yL��R����9��9RI�|wI?~�ߋ�'�"��ڈ"��Ȣ�����EW�TA_�QU�QU�EA�@�T"AP��P�T"AP�U�AP�B�T"�AP���BAP�P�0T!B@T$	P�PEDBDDYB$�EB!B$�T @T!P�B0T#BP1T!B@T$BAP�EB,�P��T"P��T $�B,B!B1	� �0T!	BB1B AP�@T"�P�@T"$BB�T"AP�P�P�B,EB"�T"�AP��P��P��P�@T �	 dP$P�T$H����A_�A_�QU|���EW��"��� �����*����"��* ���(�*�(�*������)��(�B��T��8( ���0�w�     �   �     P  
:� x  |� P� �AE(��@   
*  "�P��@     (�   " �   !� 	  �*� ����ũ]�s�w^-/6����< ޔ�w������W[�n���= =׶�9�5{�ݼ Z�Z�{��H�� �JǺ��}k�n�^�͗�n U�{eW'�z���N6��\   _   P	J�4 ;Ҫ��媯7r��/B��Z��}����W�-�r���WN\�k�M����q;� ����S�Υ��ﯶ�n�]͗�W6����m�� �z�tz��˻z�x���&�p |x  ( RJ
Ec  �>��iqΔR���:@���)A�� vf�F�傔� � �)L@ ;3� K1� bh `�1JR�((2������8 i�R����ƀ   0 
� �B��� 4�cJP14�+�]*���U� [��,������彵��}���o������/\��׀f�{�j㻶�� I�����O-OoO-��{��{� �+��.^^w�.ֹۥo |> Q)PJ  łC�o��^�����;/��=ίn���+��)�y�.�i���N��^��9v��@��}�m˾yݷ��  {+�ng��{��\ ��6�jr˭��{n-{W�����V����%嗬�;�NYu�    ���IR�  T��53T�J�41Ǫ�I�oQ&� Ob�P�*�!����S�%M��*��db40���jR��� ��u(_��~/��#�~����Jc��"���""!(�_�5誠��*�*��UPUઠ���UV*�����?R�G���Mm�t&n����M����D4X`!�tE���?��9�y�ˎoD"�z�8�C�1�4��`h�y������%��B]@�c�T�BNs����H7NR�22;`A���tm�Wm"Q����4�]�
Xl�	vI.dB���\��h��$)��� 1J��O��f�M����n}���s�z��e9�腈U�D�#@��4��pt�>i��0$���x��"2 ��BI!$`��v5q $VT��c"�X�NRo�9�c��l�jE*�1MH1�"h`YN:��Ԑ��p�ߊǓ�yi��$ֈf�\�"d�f���<u���X#�!WJ�A���V0��xc����f��*B�$F�hp�aA�h1BьhhX%d��ُ���GDd����d	P��`M)��#��)�i��� E�������7�����H'n��!Q�fB>� H�d�������MBH�$�)�ZR���k���|C�H�T 6<��O<�BF-H�>���Jc]6e�Lݻi$�v�:�AB��2����+o%#��)��caA(�B���#�䄑+*�'���A�+a�I[a��hR �@d $��14����Đ��9���Cp��`D���5���_��!�#I���#%܆��7X�`�]L���f묠T��a��Ml�8��$0�]$�@!(�H1�]kP�� D��J��$`T��b$������� ���"��42a��а�.�6Z����*3$BH酐0�t@��$|xM�?bJh��D"�b"B i0�4c�xm~}��a]
��b���S^ q�$J�P�@j�u!(�.U�Q�T����U�O泆L0�E��&�2��Q<�9�a�)�C��y$/�3{���Ls^@��C���}p�Du,�į(��ğbHB,� Y4�U�	�@�D*�}��_��Bő!)�H�FXMv
$�X#|�i�Ͱx(i�g��B�h܇7#��5����
�C$ܦ�7,M&@���=��t�{��M �!DM D*�H5�^' ���!]�(i"Ȑ�!��Rh+K�M8�
񤯚 �D(�c�!�!��B|�M�_Z0���`51c>���#��1���_	 Rc]5����H�M�m �4�0 W@PÎ��Ml5��d!�\�v�&BH '�V��F��78g��g�9��<M��<|U�0CDX�Ji�4A�E
�ȅ�XA!$ZS�](x4k�) �FOd3�O.�@�M�
���B֧@��u)�!,Û�V3��4�*Ƅ�]�6k��9,�s8n?i�[� >'���ջ�Œ��͐g��D�W����l�#�SBc�6I���`lHP��@c�q�[2X��6�z��aF!a #!p�C�h���ǧ�t��"�R���%�&�4�h�4o~�a$��#<�R2H�P �SC4��{��B%	�f��+�	�|�2YM!��M<���Jj�:�yw�@H�HE)�C��5�f;��Õ�ֳ`p�xMBR/0��8�jħ�Zh�"�W� щ�����E-�"�����J�.���W����C��.�����0I��#��<��&��B�a���7͛�tB�����H�T4&$B��5�==�
����h� �C�Pْm#L�2�L�H�F�,V"�Ā��GC �hR"�BS�!U�TC�\��'�A��0��p���]�eh�f��	wͤf���a*��SA�P�C��n�Z���=��>@��a
�C� ��c��3A9���U�/�	th��	R$`_&�!����7}}9�1&�1%ee�x���n���F�0��<���!y�𔜅F1�I>��&�lK "\�y������K�!u��Z٧J&! � �{�4#x���V$�}SF>��B{��%�o�=�<�z�(Z�$��p`D1Ӱ��߆Aܚq��;w��טf�����焦�ͧ�g���C��F��f�@`Y�B;vs{�m��v�j�@4R<x8la]k
��B����z���8sGO6l�Njlc��&��8��	잰�Ml���F�ߜ,�}9�$O�`�ݐ�k% ]$
���1`�N�}`I ц�)�$�Ӏ@ m}H���9l�$*������`�Gg#%I,�V:�sp1��y�\�p�̆��l���D`CQ*B��}mk�L��S�9�}5\0�ss=6rp��.��h������2�	�_N<0�9M�Ӹ�4zl�w�6���XSo�#���c�D��U�*Ђ�0a$"���B����,����*F8�@� SX�>K4|��y�3W�͞�'<��Gt����
�F�&��������-4�zMa�Ofk��N*E�L��e�B0��5 �a�
��b��Oy�v�׹ˬ���C����߲��	�(�����9n��o��_>�&��B.�f��XEa4s/&�&�l�szB�$U*Ӂ�4etR��d9�!n����g0�ėY̖泇�S��< !Mm2�{$i��u�T�1X7Y����DGL���h9<n�P
E�r��&��5�&����*i	#]!�	<��o�Jk�>��7#���p�'����M��aCBF��	 ��d!]��:�B4�6��78x``��dL$��REdaa H�F@!"ج���H&&���>G�p�ts@� �cO�Ռ!B�g��G|���H�� 	�0�1��*���礔6"�d��oWf�U�Q�0�X%@� z�|~H���$���S7���r��lx�1����pcD"-H�B����J�7�%=�$e�J_����y� �%�bCA+�z�S'�6l!BS!u��L�m߷�quu!�>IʇmBcBs��G�@�t���<���	��fx�!#P��0���M�!L1���.�]s��kL.���Y�Qi,��[[[�u��PB����
�aV$!"��$,��9���F��5���U�쵤��:��Q�&�5���☁�2E+!��P�f�!2再&�к/�4�A�BB�B�H����GщF\}pl �k�r�]rSQL`HB�#���p	t�'Il�܌��1)�4Ji^�n�' T;�xđ�
D�WGIM#Bo�.�����!@�U6��]8�N(K��6�h�a��R#�����>B>�Q"T���\��D��CN�`xC���vq���Ӵ�M5�h۰��� ���      �h    h      Hm�       �` m�    @ 6�            �n�         �   �`   lp        I�6ۂ���-� �5���\�[@8[N	r,ʊv�\�6Z �h Z���  ���   ��*�t�i
�ݞ�N˔U倞ykv����P�����Á�i$���`�[�h[I,09��tZ�mX;"�$�gg�f�@��E�vz�A,�<�q�����v5*��_D��t�ˬ�28���`D�[����Y�+�Yx�;Z���g��md{O�
Z�;0�-u�+-*�`�b�P��6�\W�+��V��V^e:ܳ۔75����A�N6�,��Pb�̆��[-@*�"5�l㤸�l�qkxi6�WAN��$�QE�PK�^����#���ʒ��\�Pt��WOe�S�3�����v�%@TmY@f�p���pt���Nh�l��8�8�l�J��y�D�6�ڨ+�IW�� �mU�U+0Jt�pS�E'F7 �@m�(��mUT�[x6�a��8 t"Y.��m����z�~� n� l�K����  ɯ\ !�-�� l�� ���6�G�.ۋh�Z��k�Hn��H�K�X�Iw\���"Ҷ�f�[p�8G	l;C ��� ���b���m��
������U�k�EubI�n�R��L   	�  p :B�[U*ʰ�U�Y5���[��m �t@*��>W�ڑx�UPmͺ� H�8�['LZ�[R�$6�˄s�� �v	k[��6Z�t� 6�jZ��� ڐ��:��j���T� ',�2`�d�$qʱ6�H� OY�v��`���� �c-7�pK(�:�]��;�U@]R����.��` $�d���,��$�oH%��m�U*ݕ�S�յR��j7�8�h�[�U��v�Q��e� 9ͳ``ְݷWM���m�44(��v�V4,��R�U.�m� 9m���wRmփ�X5t�k�/�W#1��f����wS2:�w���Nign�A��E7�n;t�D�j� #[ug@Uvԫ�g`���V� 5�0�$    n�-��Ԯ�-�ݕ�+H��y��� Ӣ��-��M�d �� E�@ d�Mkm�[��� ���%�M��m  hv�6v����  � ��c�FҮ �}��� 	8	:N�ٶ6��` [K��qmm� �-���   �c]��L$>�}� �d�$at�ݰ�I�M&jC�� ��v��m��� H�x��-�   � m��trI8h� �$ [@ 8 m�    �   [@   [��-�  ��  �c��ڶ� r�   $�   ����l� �:@�Y( 8 "ڐ  �d�  m���	6�`$��k�q�8�n �m���  $� U�hm�m�ݶ ���   �v��m��Pq��m��6�   �p   l�
�R�M�k�@SS]   �   .�A�bA��� �km:e�@6��`6ꪪ3FG���n� .�����I�r��mWJ� �I����UR�H^kd���j�ge�r%�-Tcn�˲�zܣl�u\�-C�CMΩ�Z)�3�Y�C`ᶕjU�8������;�K& �p�-V��]@g�	V�    �nu���&ձ�l		  �i��l   e���ݺmvd
RC�7i��.�� wE�v�f 	jT��Hm8ר m�D��0Inv�l �H i����9�m�`�Z��ɶ����m��m   ��vRΖ���  ��*N�� �pו�b֜I �m��(8[m�۷m�ml ��6݀�bĆ� H�8�Im�[�-�.�@���f� -�6���sm�[V� �\�6�[�6lT�)�lv�@:@  q"EM"ћ@W/*��V���͗`n�Kh �h��)ms�mm ���c�ݸm���Cr���8����8p8�k"(-����f� �z�1
�i9j��÷`�2�*��������^7&�P媍ȰY*�m�v ��o�	�\�E6 �i3v�6�$:�*S�N��kM���I�Z��Z�y��+���c��E��{m��nl H$�Җ��꘰��}���r:��.�vÂG-���8kX��v�m�A �� �y�T��ҫex��)	�4:ąϪU�:%o$涣T�WN��t��d��`�ƶ���AZ��3���uu�����$aG�PpUE� nl�q	�&�q�P���v��{gvn��V�rշm6� i{K�m�[~�i-�� �D�j�l�]6m�m��i-���� <t��ݗX���$�UZ������j!�����-��8A6�:��$��m�7m�d���I��n��� +v�j�4��� Ƶ%�m�鰓 p Y-6�#�  ���Plɛb�ۤ��m�6ݙ m�j��%;:ݶ ���� 8H�@�L����  $ ���    ��h-��}��|	�5� ��v�  �J����$�ְ  9me��y���iWH��@8	 ��q� [Z(&�l$Ŵ �v�ckͤ�H�`  [v�6�m�    [V�K��m�-�km���`  $�F�m��$5��-���|�� �-� �d����l��I��m�lݶm�E����iV�yj�
����\-�vݫf[|p-�I0 6��i0~7��*@6�m	 -��ו��c��jYv�68 �M0ت�;b��Y"�ګ�Z�$��9SG���`�IJ)s��~���!B�8z5�y��&ihyy�Q\�0��H6��6������w�8�m&�N�픲�.�  ��6W[��h96�kto[   $ /Z[@  0$Hm#m�m� 6� h���I��I"�� ��h۫`H�֢����d�� zt /�   ��          f�#��s9� � @t� $Y6孀 m��m� ��mk65Vm��  -�  p   ! �m�  -�� ��pm]�a�����y�$`    � ��V�m����[l$��pA͖��  Hp	3l�\N��`��fݰ��$��M+�D卖N�� -�Hm�����    h$	  &�������$�^��Cm����m�@ h�am#m���v�n� $d���E[R9�Uz�d8�lv�M٤\�H� ����s�� �4�M� 	 ��    8  �,sm� �m-�Zl Kn�][V��UJEʼ���i�n�:I ��퍳���� ���6�XX�-�� �ck5@��Δ-���-��a6�   Nm��d���݀ 6��)!�kՂĄ$[p6�%�m '@v�ڢ��i�%�Kʤ�s���B�����6i�H�u�
�5��^���J�mR�M���^���u��'W]a��E�4�4���dY
�Y�\��[u@v�K� 5Un0�ld�╪����`�4����6� 6�:�0 imCm�ͮ� �:긳���HĴ�@�-�>�` � -�l �m�r � R�����I   m��6� �`   [Cj� I6���f�� l �9��m��u ����l ���� m���d���8��ޠH pi�3lj� ݭ�    m�   m���  ٝk  F뭭� ְ  ��I     m�A�I&���e��m��`���m�    n�d��U���U/�֨�ka^u\�y��������(UJ�+l m�@  ���@  ��hn�m6�I�ph�@ ��R`����Iu ��l�*�x�53���,��)���jUV:  ���N�[RD�@UIVݴJ;m��v� [P�h  ڶ  �h  ��[@�� �  6�          [x��ض�h �H��www{��y��D�TQvE���c
R �! ���()�A�Qh��#�s�Ġ0�!PЈ��d|8���QR�� ��R(�R4�4@-�Q#�U>G���#g��\E 8� j��QO��< ��>�&� q � ��;8�Nz�P=� 3��PP�⧢���E(m�T�@N:<�D<1�?!P���O��
z �@�8z�}4K� Ǌ��(��� p�"n+�n
xpS��Oh�������AX# HF@�E���6��b����#���D'�||@��`A�*kŨ$v ��SH�	�>�� �ا=D=S�ډ���qUP� 4U
|( �lC�銨���T�Hʭ����<>E� P��<u�< �D��'�;�!D�<�Xh A< 0���H��U�~ဪ�"!�2�}`@#���(�(1�@�T�O�)��Q_H�\Gh�(�3H@B*��Q�'���H$"�Y�Eb{���������@b�� �Dd"��E�C������_��o��9!� � H-��  ��7`�d��ki2(��
�0�F�l��1���mUOnWvض��0��)d�݆�����Nv�qEñ*C�xrԡ�Ň�:v�Vܡ�V�M3��T�i�Z�*:Җ{r�;P痣m�t���%۔M�&��f����YE����WmAÙ���\��4�2�.�ulO��N��]*���&�@��q��m�I��Ǩ���у����Q=F�3�w�+vځ��Q��U� 6{\=(�-e�FwX^[ss��SI��r�[Pg�SiH�-{n�흖�US)�8"��������6�l���`J���UW���q��\*�X���X@]�Q��V�B��m#�P敇9�=��,1�=6���R��WF�1�q©pS�8(��ݬ��*���r��T��Y���'N1���!vY�[8�&��rͤ�Υ:�J��R�D�ڧ��A�y��Z^Q"� X�z$
���*��#��x����V���3Ɛ��z3x����Dc��ϲ�;\i��rS�ne[r/O����֯Dvd�C�e��!��f'�77f�jJY�H�[Z��`� ��O<'\Ԏm�BBU�ư��,�6�5Ur��!*d���g��n�v��r��CTo11�A��욹���glw=Fׇ�n�r���ٻ\l��S�[ԧu23ӻA�m�E� W�Nt&O+d�i�#;l��`.���Uڕ�ۓI����2	i�lU����&M�<�k��
�p>hwmֺdWv6����l�Y�4v�흵�0휚7��dD	4�Q�p��b܏I���	f�@VHj�����T����:t6UJ���p�p��&t-�9�6����v�ڗ�v����U�y��hZ���t�n�*��h�N�yYV��[B�6kn�[Si6Z��-�;^��
�ꭙ�n�6g����\%�$�/,jj��6ʱT� Ɨ�����{�ߟr.�iS��EXb��
lN8� ?
A"���G��@~Q�9���ԓY��B�E�
��8=5��`���N�Tӳ発=ƹ�������:I-cD�d6L�j�[R�T���۬8�d�9c���QI�/n��h1�S�в���es��Eƪ��8��݆6��+��ܪ��m��хM�mW]��\좳�ZwHZ;w6�G!�5�f��]y��É��#���3o)�.���f��S.d��2̺4���۩�e>���C�<�>��nNNy@�Ǔ����9���y�b^g��1���+ ��u�*��|� �H�UjF�$�Gm�?}���r"!%��U���׸����u�-M�%�i�)j�;��,�wq0I1��t��t��+,�]�Vf^e0;z:`�c���U�I.,���"p�8YhB9V ~�ۀ{dN��0;�:`yN��R�2��L]����ՙ��G�n�p��'��ː�hɶ��6r�ϓ����d�������0'tt����M��.~���9ye�X��ň�����*����u�~VG9� �&0=�'L�]���Ken�;V��q`�ݸy7�}� �wذ���e`��Q�2�ޘ��ȝ0&�t�����;I����뮎7-�?}��`�������λ�5B��ZUL��E��On
Ka�7>��A�b�T��N�<p��W:Lmul�dį\�8h���ߧΘ�0ޘ��ȝ06tO/�%r��%�������ݸ�^,��q`��0��Tq���rI����sϾ�74:��(�F�TH��b'�Q���P�%s���,��ŀrGT��I����1��:`ztt���� w���>]&�k����[K#� ������ ��l�����]�����D��i�)����[v�ɜmc����{�C�f�p�& ��i��e��䲼��L��0=�'LN������db+�F*�X߻� ���ŀztt����!�\�2�X�`�+�`{dN��1%��� ���=�T�9]�8��]X����;�~ٹ$��~����i*�P��a�t������7$�}��kf���^%e��S���������� �9���}��jr��XT�-r���:����Z���Z�n��͋'?�����ZDԪ8���U���� ���ŀ|��zG��ŀvM��;v�d��S��y�l��ӣ�wGL��0>]6�k����[K#� ���XwGL��0=�'L���V�x]�efU��`�wOS ��l��ӻ� ��vG�ȠW,Uڰ�wn�G;�?/��ŀw�x��Bp�G � �P��#U%!T� ?T(�X�	 S@� 4F�!`� ��M(w��w���o���V�HZv+�{>ސ�����V��F*^]�ld�cx�u�x��i�v�i��g4\��\����+���@'U�w&�^�IsVut��A��K�m���ܱ�����	=G='c�=%#[2�8��`�n�nn�,�NM��AٟU!�m-�N �V�{rU�tF����!�V�8G���㆑�v��C��Y�aŖ0RpZB��_Og`J'&���c��kO����<;\p��u��:�3iv�a3��|�0=::`wtt�;zce��Tdr�q���`���?��f��� �>��A�lY/(����/X^^e0;�:`�1���t��� ��لMJ��,�dr�qr�$��0;��t����]�=LD�)�I"��"��0=:��0;�q`~���{�4g�s�$TMJZuOF�^'�^�ݛ��܍�Syz��aՊ�5��@��%q�VZ+h�*���b�;��, �����>��ŀj�EG-$�-5s�=�߶n��Q'j�|P�1d*IT����>צ,�׋g݉�k��¹`ڮՀ��pN���GL���.��U֫��p<�����{}� �{���wn�Ǳj�2Yc�0N�\����66����o >}e���C�*X����k�׭���h=�yA멷���0rgGlu�)v*<�P�ۧ2�N��}�˺[ ��ӡ�N���-���I,U7l� ;�v�\l>�����b�:�ݘ��kOmCvYU���� ��;�>}x���%J!T$�	CJظ��s~� |{xF��uj���U�v�+1���������0��m���t�Q�G*��� �-�v����1����x�~6�4���m��Ps�Q���j���l�[v�n�Ҽ<�����w�}�|�Ԧ���r����T��GL[����B*�u֫��p��m�qq&Ͻ�ŀk��`~���l��^RD�vի��fVc~�:`rޖ�;zc ��m�7�we`�W K-X�"QN�������c��BH��J4��w�݋"9*nr��Y�ޘ�=�������z[ ��vs߇RY֭���7��d(�{5����%��s�n\���.\�d�/Mf�k�t��k�Đ����09oK`�1��J�^�ӎXղ��w ���Y��Ė��8��B���v\����o >�sx��;kr��Qڰ��f w��`�0=::`o]uڙ�h��%K/-�v���D����U��R��v`�i�X݌��U���g��ŀv{�X�u��E!D*�|��Q�Z�-�(º�+%R�"�F�]�F�yK�ݢ��%7�ǭ�v�Qځ�$����Iu��KApa�uHϹ�&&�<tc����2�v����|����$P^]%/^�!#j��x������lh�"�U�]r�T�#�	?f�`6�o�B7���G���*�V��7j�%'���3�Q��HI�n��2���-��;&J�΋��\��W@,}�����|#�WOF�]r[rl8A8�v��÷��n����v5t�D�W��{p��L]��oL`{dN�b͔E��Y\�,�`}�� ��ۀ{dN��0=:];���+�3,�WX�u���Xz!L�^�����|���P얩l#����X��Wt������J���ww$���>m��5D%�ok�����07J��V��P��[1LW63/Pu8��t<;�)nd�w�hQ�[�U"�U�|�ݘ�{� ����\�����`�=�����-N�5�$��~͎$� �E���:`n�遪t��L&^U�x�V+.��Lt���K`�ۀ}��Z���c")V�wq05N��;�c������b�Y\�-�`=���$�=�O�owLXm��5(��\ ݪ-���D�S�]^gi��{#Ŏ�=,i5����$�Y5&,*�"�
B��Y�?{� ����I05N���'�3)^]�U�U����6�f�D)�ww�׵�9�ـ|�m�+N8�v�:��7wpܓ���ks��/:�bg"�#�D���T9
�P� U���3|�@1S`��$$��S@��J D5���5�Pl�#$`�����;|y�>Q_ ��Z�»R�i�x!�4h�4@�_���@�
+��9⬐P��Q��t�A@4���� �TC���0H	A�;~�G@��E4����{��N/�>��b��K��-���ܪ�E,���Ok^� 6����LXS�{�,�z�]QQ�Ѵ� ;�����צ,���}u�Hy$�(�l��6��Q��l��ѵ�ݹ�����5���4.���GE�=�7lڛ� b:k��� �5���;:��ّ���}=�~��H��&� r�`{}�?�K��G��Ӈ�ɯ}x�ubԣ�n��[��Y\�,�`~Iq?m�<�\�R���{��`>�X�n��*�EQX��k/ ��	�S��GLx�D`D�H XՍ�(�qs��|�>ܿ|���w�;*r�l�;��ރ�R�-�:�&.�w~�������K�&�Nmפd�	*�c9�f�Z��=�ty��Z���ܻ�u�x��2̦����`E:[oA�Wyիm�ʯ$d����x��l	�LN���t�Tŕu�/0+�L�K`M�:`t���_kj�uD�9Ee��~w�p�~پx������~��H�-M�@�U`~I7�{� ����\���wk�Iȟ?y|�B�Ȅ�G���=w�[&�dz�.�2���ã��g6;6e��f�����f��e�rH���\f ��#P�l�'U:���9��q�p7L-f���:��v
}f�Qg���\�r��]��ݚu�<Un�m�卷2�S�^������l/c��4�z�e�@!x���7�JB�v��q�6[��^���r���X�nW1�mh�rۄ.��ۘ��{���������M��6�6�嶦����[��^���S�լ�n�q9Z��av����_����RK`M��0	$��Keҫ2��3,��L����%:`I�	��x�wtQ;*r�j��[0�u:`I�	��0"�[aS
W,�Z�X�2��)�I&0'_D��Il��b�5w�Z�V�;K�-���&RK`M��0	$��ib�߃f{zZ^��YݬvLr)>�W�k�m�l�6��+G=�'<L�X����߇�u�>6�`[w��{8OI.�jj��V�l�7�Ջ=Ĩ��.$�L(����o+\���f���S��I�a;UX�����ׇ��DB�s���(�C{��`�{5r�����Vff0'_D��$��)� �ݸ���"��
��Y�u���;z�I1��t������e]䘻W	�Z\7;�˷m�\Z�:mK�N�v�\tq�ĥ�q"Y�nk��O�o�����0�cT�lRK`o+r�݋fQ�e0�cT�lRK`w�� ��uj�[*v��8���~��߾�[�Lkc�L�Ss��N�����ݸ�&��X�-�B��`r�[���t��K`w�ћ��+��[0��1`I%/wo�;:���n���ZUL��ѡ�'�]m�Gϩ8E�3z����,���U���QH�j@NR������������:`I2+�	Id�����=���wf߷V, ����..6}���'BB�-�X�ݬ�mb�R������׳ ������,��m%��\I�}��wo 侺��!H�!(DD$� ���#@"�Ө���;�܆�^�sУ��jU`�ݸ��׵��{Xx�ŀyGz�S�+�m/v�{Nz���r��������].��{h�n�Q����?�VsX+eRUyk������X%���6�l/����5ҙkn蠱]ԒM���}u��IU�� =��� ��v`�tf�UEc��I��풝0�1��t����-�Z����S��V w�ۀ|��0S��;d�Ltȯ*�˼�J�Www�r_]`K��k�wV, �� Xp֎$qn�kQ���ꤜ�%-k#�)`ê�ٙ�ۉ�N�{p���Ӵ��Xs�P�:5��8�r�mɜvӬ��.�4܇����+��Xq�l&6T�ܘ���R񰕍���N�I�ˆq2��]&� �ף�Ք� C�۔Ω�j�Xz{F�J��2�V�v�76\q˰��^���gc�ۭ�e��sR5��H��T�Yp�F���[�Mw~�������ﺸh,B\�\�2��=�wU��Z�O�]h�ſ�y����9r�D�nJH�Y�=���;��ŀ�v��0���`=~~"vT��-��a���Ր�qs�$�|\��}���m���Lm����������=�:�u��VX�I.�3�I.R:��Knt�y6�7VCm���W�Gm#����Ir�մ�[s���%�%;I%�&{ͷ�z�:�+R�1�T��M��ߒK�Jv4�^���$�)[I%��bߕV���=���gm�uܱ����C�<�õ���wk��%�V�c-�=&�܊����]rS�����Ir�մ�[s���m���X���0����m��y�>��A������y�.Y�V�IKޗ�$�\��i$���x�T�K+q�_�ͷ׻�cm���g���.I6{�!������6��vaP��0��Y�4�[�"��J_Jv4�[����oˉr?nx��o�<�E��,��̴���R�S������|{RI}3�M���]���m��ަ�2�R�U�K1���8ݲ��Kv�f�-ٓyz��c%aS%ЖB�ϼ;��:�u�QaT��o��i��m������]����Fߟ�b��o�{�^_�e݂���Ͼ����w9舅���e�����_���um$��p������I}O2Һ��XG]��m�������׺b��x��f�P����w~Nr�o~��ݶ�y���+�q�?~m�^�����JH�=�S�bi/�]�w�_��Rb����j@NR�����sOߛo�۞��K{��I(�[I%��x���%mY㧒۴n:�Yݹŷ��鷣�9��Ad��OV�"~��MGd��m����~��M$��ɞ�IE ����K�?�y$�}�MB�$��-v׍���o�ؒ��R�����y$�옚I/q.�)*��l��~m�{�)�������$���I$��g��]�����رfefU��[���$���Il��i��zY @`A�D!BBF0B1C�R V� $�*�ߞk��&�7m�ǯ~��G���Ki��m����o��g��]}cI%�=���xe�A��&�)tL�p�җm��A�9�]�:�άFͺ��຤���s�[:g��]}cI%�UUn�J/�u1�߹������+$��ߛo��d3�$�����<~��z��Sm��v���l{(�Uڈ
q�Xcm��sOߛo�w����sܶ�����m���6����pU5���C�S������cm%'L��K�Aմ��Ww����K��["j9"�!��m������m��L5�m�}����߽ϲ��n>)�@0R$��V<	d����a�d��#��6��N:SP�!��$�X$`���HH�&"H�6$�������� ��"Hŀ$D$�\;���4��D�i��ŒGB��!*:A �,��bA"��$���gq;�O� �C�M�$"E�S`4ె��v1����b�Q�,J����@�"E�Da��P�BH�b�dd$$FH��O��X��B$�b�0!�2��� J�C>+��d
|b(i�6�YPyd(���#H�:OO��D~����h1%?q� @�j23�Gc ��u�2�Z$`00���6"&+	D�, C�ً ŀ�B!�`I"� �O� E�"�bD�HA�$� ��&�ۢ\�F@��߆Ԣ@k��b�E	Gig�����vIm��!� �)BAm[M�q���%�m�mN���[QD��)��[�%+Z��A5HMD���lES��#���k��c��[��#�5�Pޘ7�:����;r�\�nv65�(�˵���:�IW��2���c"o��>���Ç��h����(�"��%v�i�d� ��Ʀ�H[l"�N{B5v�Ke��ύ�B68�R�^�Ȳ��r��Qɻ��\��Ib��mֹ�A���S�=�V�s�a���Lcb��w�a�q\3h�]�y�����f[*�l8�U:؄�UU!L�&}�"�(�
��U��ptO=Kɜr��j�ns����IC���9�erҭ�ӭ����(k��H�'*��:X��X5�\��*��,�97;:������G77]���ȦO Ҍm�b�yQ����V)��h8����J��F��ey���e�\2����z2;6�t�eR�(�yUZ�g1���q��L�W1`D�@e̛c�v��w*d.Y�[?Wkч��{vM�&����vx���I��ݓ$9�V�=7h1ˢu8^�݂�8�-T�,D��۬����na�-��v�rj����$���T�CK�٤�n��H�
ۓ6�ͭ�m�i"4��Xݳ1�A�E�:7D����s��,i��vrJ� �'k.ڳ!\���u^�]2��\��ȶ����3Z�2H���k��od��Uڕi]��eҳ9Ɗֶٶ�]���7 *�j�㓪���)@Q�X����k��EY흮�$ԮwJS�(����V��:���볰.sK�3�۰�e��ʦ���G;n������U9z%���tô�����g�j]���W$����u[/�]�8_�i6�C��id+G_S���lʵR������6���m��7i]��0 �e� �k8֕�p���� M�6Iy��a�؇3� ;lk333333ѣZ̗���Q9���A6@}������>��|�X��񻬙�fB�2���7HS���:,���5��Z�Ѹ�39�N����X]!e%��Ӧ��Ym��O;E �x{=w!�&g�f���Ud�'wp\�m! ��n��tWgs�#)�diX�ƍ���3���ɷ���mj��DTc�x
���F�5����|�~S�z�'[&%Gl:٥��f)#�/hmͮ�0�+�,�bt����piw=L����}k�7Ѽ��m���k7�=����\�/nm�&�9�TvKl�7,�ߞ��1���sOߛK�GcI%.t�y$��v,WwfZ�aT��{��?~���=��Cm������}}�����wC�[kNZ��Iu��i$�N��/�~�Ww�um$��sǒ�����o�-��G-���`�I)��=���um$�Np��K�Gf6�����?*����H������V�It�y$�옚I%Ӧ{�%�E��i��&��K�B���v1�]��6;��n�.̪�T9�m6����z$����It�y$�옚I%Ӧ{�%�Sm���pU5��ȇl��ͷٻ�M�j�M@XAB$D5�i ��AGKS3v�����[o�ߌSm�{�~��$���ޘD�,rJIE���4�J}>�y$�t[I%Ӝ=�����cm��zO�r���cn[��%ˠ��I.���$�\�ƒ��U]��}~m���O�r;b,*��o�8{�%�#���]:g��\������ݟ��ҶB:�$�:�6�k�����WaŐݝ�z����9����>��܏e�,�u$��󱤒]:g��\��� ?������Nr�~����5n��Y���m�{���)#׾1Lm������m�n�3��������~UUc��ə�[ooM�ݶ�~�Nr��hF������!����}~m��رIjv���jʵy3>��B��o<}��ϫ}�d���_v��������+m���󂩨��D;e?~m���V�o�������=�خ6���4����N�
-��Q$����;m�2l�Ϟu�\m���=ka�Փp ��޾�0��Y�q�X~m������m�B:ƒK�8}����󱤒�����Uu�m��-���ϴ�W<�����ߛo�}���o�ݿ�zH��Q{#�B�l-�ˍ��۞?~m��܆7�#�o��Ͷvy�\m����t?�ѵl���������i$��}��I1E�%�F����	B!r"���o���ߛo�Sz�YTr���it��I1E�$�Np��J_GcI��v���v����q�&hFu�a]�ί]ƈ��B�;#�.��!��F뮓Z�]���y$���ƒK�8{�J.����}�������b�%uK8+Ȝ��1$�Np����_)�h	���S�n�*�%��ȇl���ŀޘ�="�������Xe���]f^S ���S; ���X���[U��m��-�ۯn����� u��0��KaJSK�&i��<;ffa�2�-��&�f싗�s���eRu�:\�Wm0[�Lc#��s�8s;��ԝZa�͙��.=f^u�;e�z�8ɗ�ض��ǉ"��,�n�p0PW<�E�̎�gpv�n -�V����N%:��kC�%�9^u3����{7H�n�����.�@Y::M����w{;�<q��(:	�gj��&����#���(�c�6�*�Gk��rL޳.�YKrf�]kR�X��V��#�k�;�ƪ�V���h{��kv÷�NXX㐤��Wo@��o�w�� :��������8�9�0Eҩ�*U�]ـ7׋6�={xǳ��u��~��L�8��8;*��v��)���`t�遵!�J�-a����c �E1�Ӳ�0�v���bjZ���NJ��;��`t��t����	��5ZyH�8^.یݽ�mWS��zkp��ۜ�U��E�ղ�NDV�[�ֹ�So�ߟ��0�1�l�1�Ӳ[��P��(�%�� ;�ۚ���s����P�HMv]���`��f�JK=�쥵K��r� �|�p��0;{ �6t���R�̵j쬼�^b�`ṽodΘ�仾~�ڃ_��,Q�F��� �ݺ`��^���;xx�#�d�F[mٞޖ*�$\���l��[%��n����I�qun�kl�x'P�XjD��m�Θ�6r������06�!v�V�;jG%�����s�K�I�}��������?n�X�-R�
�
�c�d{ ���meUִt�\ ��{p۷\(5v���l� ��f u�� q�]�l(�/^i�u�g����G-v���� �z��}�`��`k]EN�jj�gN��]�rf��tyv��֫Κ��<#��Gvl����I\P�H~�����?��d{ �:t���R�̵j쬼�^b�`t�odN��>޽������,�5l���܃ ���S; ��JJX�G��eX\�8��}p����:�l�QiD(��r"""�_3 �>��F��*ԎKp��ۀw{t�7��0�ݸ�������X5K#���:;kԓ	�b8�޺3���c#�h�g�Ȫj�jP�������Ӧ0��0=&Eee*��0̬��/��0�1�n�1��2���,�J8�k����p�r�J!D)�ݽ0�z`��R̤�^ffZJ��S� ���� >���>��'�r
�Y-v�� �����0��0?US�]��~��^��.٦Y�V�Q&���k=�ۣ�J䶽˞�^�&z���uSu��d|��%��mY�:�����v9������r%z�QYW\=%�b�Wn�&Mn���$[�6�q��h�[�a�m���n�����;b7*��9�7$)�������q��w4�[A������^#\�(���;X��gD��=����Y��T�q��$��V���u/~�Gͮ��)dHU9J2N'T@q��#s�+�z_N�n���ֶxy�hx�����ߠ>��0�1�l�1��2t��\qQ�lq�i�ov��׷ ���0:�-�-Y�X��]�0��0;fA�7�gL`znŉ�Z��U@rWn߶�oݺ`�ݸ�7�k��>���MGl��eyx0&�A�l�v)�ٚ`�K�xb=�v�ah�
�n*�f^��[��z��6���S�C����}�q�T�4�EdC��|���������n�~�� ����]D��ۖ��ST����WW����`I�ӥ�>��'�r
�Y%v�ww������ﱀw|������ZYt�ş��3)�����S{��������߲�Y9\��v��[�a-�ͯ��{� |� �w���UlKc��Npl뛺�X6�`��/0�nۮ�p�u��:��{�w���:z9�����ͬ��ŀu�������@w}��=�z�)�]��B�@MYu�s�0&�A�{��]ķ�����YU8;ev�	-X��� ~����ˎh�׈g�����S^�"	�-�hX���0.�D7�Ư��<�DMuj-�4����&�f�1b1��G��Pddg�h������%�����!��x�(�žBW{x�qDH�0���TN|�&"��T�*���>�8"PO �`>�<T����~G ���bI%%�I����}6�n�,�Δ�|�I"�!�ʰ<�w޸����>ގ�::`{`	B��Q����I^f��`�{���q`x��Q���>����M>�K��1�ѧ�k<�q�ղ7bxܽ]v1�����u���7�J��X���O�0:tt�;d�/���?u^�v'`�*rՀ}��L�L`rڒ�::`{e%*�_+�X�� ;���:�[�q��}� �ذ��valv�jG%�e�D�����GL=�uܖ��K�N
�-B�������� ��q`n��:��_O=i�ԒX��WSi!ڤ���n����n�d�=g�F��^D뛥��L9T�v��Z���ذ��f�gV�����>t�7�d�+",���d���CgGL�0=��I���[m�`wn� �{���0;nD����(�X�ݕ�����|�������0;nD�ޙ(`~���GdE�P�KV�wq`�K������F�7� ���j!+��)H(��kJ��
�BD�H�Q"-����"�E�$A�����>[Wm[�$lg��l�ݼF�܍���k���4s�m�VQ˝n[pW�v����s�zpƺ�M��] �F�n�^�;Y�4��[R�pX��
�K��X�&�ܷ[Ñ�x��;kM���|L�kd��7Y�V6�k���i�{hl#bCx�f%dW�?�pim�����s�8w4�3eًl��ǰ�i��<Ԏ��C��xܪ�7iYynO�{�;���ն��m4v����jH�tɎ�xy�m�����u��vs��n���*:3�f�f]�0:_�07�J�:`oH� ����-%���Z������gy_�;�t�ޑ�v�L	�]:VU�WhW��рs���9��a�P������{�y<�v����l v�0:tt��܉����a�.������=S|�I"�!�ʰ�M׀yo����wO�0:tt�+�D�.��2�)�Ӳ���;���7��m�K�p��۞sk��Ӷ.��T��rIUC�ڇ+��i�s�x���^Q�;[��r5�w(���m�9
����ʷ����]勋�%�K�=�{��l�}���4k����V����?}7^\Mﶞxw}� ��or�Y9\��%X[]y���ٳ�}�ڰp�����]7�Ikp�V�rW�w�wf�{�LN���0;��v�*��e�_;tF�.ڽ� W�R��:��9x�n�#,d��D�\�X�8)Ij�R[�����������cg��T��a����`{z:`yt���7�0>�wy&�=��7�drRDB;V�����Y�f�`� D �(ED,D�V(l����'6���;��,���G���[m��-��ޘ���GL>����[����#t�B��Ye�~ۦ���}����[ �I�Ҁ�o,���rJYҜ��8a�n��v];8�m�״.�N����T���Q�i�}��,Wt��>� ��|0$����E�e�ʰ�{�<��޸��� ���X�ݘUe�бV�nۀ�L`l�>K��� �����%ӥb�Uv�qJfn���?o�0��X߷n�S��ۀwv�,��U,f^U)�}� �����٦�6�(��-N�*�B��:���흊�u��\��n�Ǖ��eS��K8A_�_}|]�R��wB-fW�'}�0t�����w���L�C��ܶ��nlL�׸���, ��؅28�)ܤ���0�ĭ^c��:`n�t�;d��{� ��4����;AGl�a)}{��9/v���x�O[�0�~���,p,� ���0������u�� �:�`�F�!Dq"D$�*$H���n��d��2Y2�Y���t�����m�^�m�7k�Y�}���6��I �6�w;��E�x��8A�\R�9ǻiSC�.�n�t
�b��&Ӑ��N7����<�8�Sg�i]ՠ��#Nc\�v�=[J���	�:�~tq��8�r�e�8��K�H��n�Z�cX�a,C�����p�6���]������;��s�^l\/n���{������`��'aݦL��O�յ����cW�qmr��qg��k�jK�!���Y«-b��;g�����w�L�wq`�wf�wb��%%�W�7e���ٟ�(�(J�����;;�V s�۞I.6w�����-�KKm0���`yt��7zc{�-貅����Ki��s���o�0���;�f�/BP���`����U��o33.�2��L`ovA���M�__E6J9kMб�m�ku�:��c��u��W�*�PW�"�ևD���� ���$����忀���~��0�n�.s�����=�$&2��Qۙ7$�g�z�`����z�=͸��ۀ}��g��l��o�Zۜ�e�WY�� ����7�cgGLt�0�nɅVZ:�b(�m��I7�{xu�,�f�2��x;�K��YW�6���ŀq/�����޸�{� ;�6�rڭTn���v�KۗF��α�f��n6)��7���NT�;�V�qX��ah�W�>�_ݓ�L`l����2�~̵wu�*����͈����w^��>�3�q������M�[mn[p����<���na𰈰�ҩI�>�� ?}�p��܃�I
I[$�a)��`ݽ0�n�<�Q-��۫Ă���nPM�i�~ݺ`ʿ)�}� �}���`{��J]��"�]�B�@�.7^q��s�]��X8 Oոf�l������}��]��Uo��~>�wL`l��d$�ee�L���r��n� ;޻�B^��������v��݋ B�]V!T�s; ���}I����`nú�IS�Z�Ձ�q��g� ����$��~�ɚ�$�Ј%b�.���%��I.ǹ� ׽ڢj�I*ɴR��0�n�B^���_ ~�b�7�`>�>�jr�c��Sv�v�����]�Wt7�vz7<[g>���r;�J��[m��n o{� �{���n������ �wD��u��J�%�^,����� 5�׀�w�J!L��^$!�YA�
;eX��� ;�w��L����{� }je�����]M�\�ف�	B�}ݼ ���>�X�������§m�^X�L�� }��� ���7x �Q�6�#M�~ '�� ���f� 6D|׊�1S#)��C���/�lB��TҾ���h-cu�-�1�8D�x"z�������V�� �`B�t�Ƞ{篲1�C�R	�U
��h D��+ 1<�����ȨN0M{����~�k�+#��aA �t���zzx�48�wx�b.UM'��#���ń"�`��	��}ӹo�n��8��l�� ����8  pu�m�m/ZH	6���ڢ�/;*�1cUu�	@�*�E��VG��W�ug;���㢉0B�tۃq������Q��:�qGc!�t�m�;i���̃u���N2.5���`�W�7L��*:m��{g`$��W���j������qٶ^8)-:�Nn�����l���T!ֹ���9V\�*�ɶ\r#�뷳ڶ�����pn6�k>;lT �ey���Pk���صq>��@_m�1�A8�n�y[rnݕa�ۥZ��g-('lMUS�����p/<�m,S[S�+uvm+�X�ܓh��:24�5M�VUyj w�UUR�t�i��T�lu�)v��scc��]$-�J-�S���r��[i=j,9�۩�����8ݏPIn�t��������L� ���������n+bU� ���ڦ�T����	��A1ll���ͪ�Ê94�\�1�.
q��'�&�(�R�.6C͛�8�Re:S-rg�������aײ!�U�D�y��!��Y��JG\1��p���R�\�!I�m�Y��$��Sڛ�ڗF����< 	MJ�]���X'�����F�t-��ĉe3β9׍;D����F:� �ҹP:yb�%@�`W:�㠥(
5m%�*��#Rr&N��4��{iԂ$,�$�A�dt��,R��h8����y��n�މ�lT��*һxT�R%�[��J��W(ʓ�c*��J�X��$�crU��[% ��΍�]S[g�W��%n�ÒGl�u��T�Ҭ��23+;��ɝ�����WgiV�-�s�TOFWdK�1]��ne��#=�3ӼuA�)vmv�ka�]I;<���Ŵ��[�Hm�l�R�@5*�TqSv�m���
�����,kCm�-h4�v�{<������6da�l�1re�33��m�pq�q�V;mf`�՚�K*�.�`'�⪕[��)H���&�|�t(<�N m`/H&C�@�"z����W\�ك^�rP:fn�<n��qE���$�;���m�!��s6��^1�`䰏:�\s�ܝ��넬�;`�Z�.��u�J��˸�m�l��8#�h����3\&.�����N$�rq��3ƍГӴU��9m����95�����r�z�Lm�K��*09C�B��6�Ή�9ےv�����;q�;hwEM��nr�Nj��j��M�v�# _����Pj����a�:Du1�q�����G�ð��ϋA�4�my���ő:��*�`�ŀ>;f w�߾�5���=S�:J�
��V�m� ;����v�ow��v��%�9\�����1�l��0;fA���G&)S��m��m��M���w��X~ۦ���޸�'�R�R�+q^cgGLِ`�c ��ԗ�F���)K"E)FB��"��#�p*	Ȩ�+UGȫ�iڰ�q:���.u��,k2���vɌgL`l����oV[��X��L �۷?.�
D(>�$�����}��7$��g�g������Z��V�m�ߧ�����?���|0	�}�oKy��$B���m��O��~X��� w�ۀ���?3����T�(;eXِ`*��vɞ ��::`��,6�uv�:�nt9������BuX�h��%���<�<v��wYk�<ʌ.]T��bX��{��r%�bX�����r%�bX�����~I�MD�,N�������&q3����ԕ;��[���Ȗ%�b_{�siȖ%�bw��iȖ%�b}�wٴ�Kı/}�sj�.3��L��wD��8��Y�8r%�bX�����r%�bX�{��m9Ǐ�t/��D����q/���m9ı,K�ﻛND�,K8���HC�P��K,�8�L�g�@�N����ӑ,KĿ���6��bX�%��w6��bX�'~��6��b���-�&�����\��+�����bX�%��m9ı,�~�m9ı,N��xm9ı,O���6��g8�����89m�Ԝ�4ږR�]�\^�`4�����Y9�.йu���M]�<u��8�c�e,���r%�bX�����r%�bX�����r%�bX�{��myı,K�{��r%�bX�{�y���2�]�[s3iȖ%�bw��iȶ%�b}�wٴ�Kı/}�siȖ%�b_{�siȟ�U5��S���K�䙩�3Y�6��bX�'~���iȖ%�b^���ӑ, A�MD�~���r%�bX����6��bX�'��g����9]����/�8���'�����Kı/�����Kı;����K��`�X������C��N���ӑ,K���d���MasWY����36��bX�%��w6��bX�'~��6��bX�'��}�ND�,K���6��bX�'�P��O���m=m.�a��.Iζ�ۧ��ٻ%�;����f`�70߮�}��|��25��%�bX�����ND�,K�{�ͧ"X�%�{�{�ND�,K�߻����g8��ޭ=~V�V+Im�ND�,K�{�ͧ!�Fj&�X��߿fӑ,KĿ}��m9ı,N���6��bX�'�t������ˬ��k.fM�"X�%�{�{�ND�,K��{�ND�ı;����r%�bX����m9ı,O=����`fK336��bX�%���6��bX�'��}�ND�,K�{�ͧ"X�6%���6��bX�'���f�ZіMh�CsY�ND�,K�}�ͧ"X�%���fӑ,KĽ��ͧ"X�%�}��ͧ"X�%��yڈ��;���p�Z��.�U�H��E��l�_V�\f�O$c���q۬�V�ػs��h�=v��1�\Wm՝�Z&�;I�0��V2�sت�S�9;p�U�2���5tO�j�\����j=V.p�ֱ�����-;aۮb�'e����0��-�f��rS��2��$v�m�)9������]]��n�of�/R�Mj:rٶH����%JѦ�w�߾�{��>^w�����ˤ;4�,���'^����rgnvou:�s�:��<�5SE���QYm3�㉜L�g���ӑ,KĽ��ͧ"X�%�}��͇�b)�MD�,O���M�"X�#8���>K%-���㉜L�b^���Ӑ� �MD�/�~��ND�,K�{��iȖ%�b{�{ͧ ��&q3������J��[m��nq~8X�%�}��ͧ"X�%�߾�fӑ,h�lO}�q7�	�{�ڒ	"����\lpN�x�\@�\�����Ȗ%�b{�{ͧ"X�%�{�{�ND�,K�߻�ND�,K�O�up�fI��L̹�6��bX�'����r%�bX~��ͧ"X�%�}��ͧ"X�%�߾�fӑ,K���2���i��h��"��݃g3		Nt��Βg�/��D�A#m痫������{�ı,K�{��r%�bX�����r%�bX����l?�<���%�߿~�ӑ,K�����Oٚ�`fK336��bX�%��w6���=1D�"dK���6��bX�'���6��bX�%��m9�,K�~�2fjd�Ham�ͧ"X�%�߾�fӑ,K�����ӑ,KĽ��ͧ"X�%�}��ͧ"X�%���)�əf�3Y�6��bX������"X�%�{�{�ND�,K�߻�ND�,K�}�ͧ"X�%������պ�L�jf��r%�bX������Kı/�����Kı=����r%�bX�{���r%�bX��{gu�E�K-P��-���Ƴ�"%�8|��0�E��<�9�bۋ���nga��F�����D�,K����iȖ%�b{߷ٴ�Kı>����Kı/����/�8���-���B���k#��D�,K���ͧ!�EH�&�X����ND��a���{��ٴ�KĒ�o�!|B�B��TB�kOP��Wy&�L��s2m9ı,N���ӑ,KĿ{��ӑ,|?GI��N���9�~~ͧ"X�%�����K8���-�&��[䤱�+�����bX6%���6��bX�%��w6��bX�'��}�ND�,Q;��~�ND�,K߻n�����a��33iȖ%�b_{�siȖ%�b{߷ٴ�Kı>����Kı/�������&q3��Q�$~�K�`ӐU�,�:�m���{H]�����j�s:6��E��(ӱM�nq~8���&qw۞19ı,O��xm9ı,K���lyı,K�~�m9ı,O5>�N�L�0̐�s3&ӑ,K�����Ӑ� �Q5Ľ����r%�bX�����ND�,K���ͧ"~�����]���Q��Ic�U�_�&q1,K߿~ͧ"X�%�}��ͧ"X�%��~�fӑ,K����iȖ%�L��=��+��m��m�/�8�Bľ���ӑ,K���o�iȖ%�b}�wٴ�K��C�G�✑7���m9ı,N��sS5uu���,��fӑ,K���o�iȖ%�a� w���6�D�,K��߳iȖ%�b_{�siȖ%�b}�g{�e˙&�b���:�F��0��N�4$����mc�{�uT�'!;8$�䥢}��Ou�bX�{��m9ı,K���m9ı,K�~�lT�Kı=����r%�bX��ioNfj��L���\̛ND�,K��{�ND�,K�w��iȖ%�b{߷ٴ�Kı>����r'�Ab.�j%��ݷd��ff��e,���r%�bX�k�kiȖ%�b{߷ٴ�K�D�N���ӑ,KĽ����r%�bX�{�xfe�)sD���m9İ���o�iȖ%�b}�wٴ�Kı/�����K���MD�?w����bX�'���S�d̳2e����6��bX�'��}�ND�,Ko�����Kı=�~�bX�'��}�ND�,K���u�^�_���	�*UΌ�vrb����0��q�C4c�i7��Ol�6��/2D<�Q�C�v��mc�,&��Ki���=����1�ɧ9��k���cg3�c���3�Z��G>(�u����q(DW$�#V�q����#>P�m��J��u6�-1@��q��2U��ͳ�AZ�F�l�!xvJ��;I�����l7���̤�n���?��w~wv���s�ݾ��=����&���{Or{gb�^��.ks���2�=paS�#\��P��wK�KZ��>O"X�%�~�siȖ%�b{���m9ı,O{��6
�%�b3�{��_�&q3��]��z�v9s32�ffӑ,K��]���r%�bX����m9ı,O���6��bX�%���6���bX�'��7���]]k)�˙�fkiȖ%�b{߷ٴ�Kı>����r%�bY����ٴ�%�bX�k�kiȖ%�bx};ٮR�����i�_�&q3��[�g���Kı/�����Kı=�~�bX*؞���m9ı,N�������JWl��L��q3��L�{�z�9ı,Ou߻��"X�%��~�fӑ,K����iȖ%�b{�d���;���3�pRg�f������v�-�,�h8��]�f{]����wu�v���z�8ٙ�ND�,K�w��iȖ%�b{߷ٴ�Kı>����~yQ,K��߳iȖ%�b{�p��&[sD���m9ı,O{��6�� ���ID���!H8t'�7����iȖ%�b_{�siȖ%�b{���m9��j%���Y3,�2CE��ND�,K�~���Kı/�����Kı=�~�bX�'���6��bX�'���GtMC5��f�kS3&ӑ,KĿ{��ӑ,K��]���r%�bX�����r%�`؟{��m9ı,O{��k��3Z�332�ffӑ,K��]���r%�bX~P����6�D�,K�~���Kı/�����Kı;��Ѯ�%�����رt�,�Ѯp�L@�v9�=�:-�n]��Α*��Kf���bX�'���6��bX�'��}�ND�,K�{��iȖ%�b{���8�L�g8�u�O�:��*�<�iȖ%�b}�wٴ�?D5Q,N��ߵ��Kı>��ߵ��Kı=����Kı;ߩoNfj��L���\̛ND�,K�{��iȖ%�b{����r%��5mS
Mp���7�y��(n�(A�X!� ��H�&��t����
0�Fh0<������i��|H@Lڱ
1Z=�R2Pbi��"4J4j��)�$�]��
h>��ZH	��M�Uk�*;�O�u�-�����*>� $<<O G���T�y}@ ��ʪ�QSj��^.mOTh����M��8m9ı,N���m9ı,O}�[�w0�X�FV�f���bY�H:��~��[ND�,K����iȖ%�b}�wٴ�Kı>׽�bX�+��*�N��Er���q3��LO{�xm9ı,?# �s��yı,N��ߵ��Kı=�{�m9�3��OV�~�����(��N�wnmڵ�r�-nk��a�,8p��l���^:�E&d�蹚�iȖ%�b}�wٴ�Kı>׽�bX�'��{��Ȗ%�b{߻�iȖ%�b{�}u٢���,j�[L��q3��L���zg�ı,Ou��[ND�,K���ND�,K﻾ͧ"%�b{߈wSW��m��[3����&q3�����/��bX�����r%�bX�}��m9ı,O��{��"X�%�����53WW3!���ֵ��r%�`���~��"X�%����fӑ,K��^���r%�`|�QP(�^����Or%�;��r%�bX�=$�ٮf�Y�jC.���ӑ,K��{�ͧ"X�%����u��Kı/~�siȖ%�b{߻�iȖ%�b~P@��N����˷`���VѢ���a�X��V6ppA��t��pJ������}H��R�3&�Ȗ%�bw_~���"X�%�{��6��bX�'���6��bX�'}��_�&q3��]���$U>;���"X�%�{�{�NAı,O{�xm9ı,N���m9ı,O��{��"X�%��w�d�a3FRYu���Kı=����Kı;�wٴ�K Fı>׽�bX�%���m9ı,O5>�N�L�0�3Xm9ı,N���m9ı,O��{��"X�%�{�{�ND�,EB���w�ӑ,K��������jkY�f�32m9ı,K���m9ı,?(�u���f�Ȗ%�b}���m9ı,N���m9ı,O�|?��ÿ]���C�A����I�y��{��5�����^�vJ͸Ƀ�f�B��>W^�,r^� ��Eon�۪p��4$��t�۶$�l���K��6ñہ��*��Hn�9��덭��H#v��%F�.��r�9l����ԉgHn��!�UǛ�W`,695v�D����e7E�L��C��Ɛq7`:i���i�nk��28ۈ�8�YU�����m����X��'$��<z��Z�:]v��f7#aۣ�j��]��{��7n������ͧ�,KĿ���6��bX�'���6��bX�'~��6��bX�%����㉜L�g��?~��;h���ffӑ,K���w�ӑ,K����f���MD�,K߿~ͧ"X�%�w���r'�"(:���'O�?����r�C.Is�"X�%�����m9ı,K���m9��5Q/����ND�,K����iȖ%�b}ߩoNfj��L���\̛ND�,Ŀ{��ӑ,KĽ��ͧ"X�%��~��"X�%�߻�ͧ"X�%����$U4�m�/�8���'��siȖ%�b�����r%�bX�����r%�bX��{��r%�bX�����YB��ӗ��F-s���s���񗇎D�aN-��Ol��Z�؞��%�Y�ND�,K���ND�,K�w}�ND�,K��{���&�X�%��߳iȖ%�b{���?e�0�32m9ı,N���m9��`�r&�X���m9ı,K���m9ı,O{��6��b���/n�qz(�b�QGKi�_�&p�,K���m9ı,K߻��r%��bX����m9ı,N���m9�&q3���z7'�l�,��3���ı,K߻��r%�bX����m9ı,N���m9İ�>׽�&q3��Z�x��8�:ݖ�"X�%��~�fӑ,K����fӑ,K��^���r%�bX��w���q3��L��H�5�����49EF�\�ݶLp]��Vg�s��ݶ��Q<<u�������/�8���/o��p�Kı>׽�bX�%���lW�,K���o�iȖ%�b}ߩ_��c���X붙���g8�ų���r%�bX��w���Kı=����r%�bX�����r"ؖ%��K�ۙa�֤35��Kı/~�siȖ%�b{߷ٴ�Kv�M����wٴ�Kı;����r%�g8����+,Er���q3���}�ͧ"X�%�߻�ͧ"X�%��{��iȖ%��&�k�~ͧ"X�%���ҟ�2�a���fM�"X�%�߻�ͧ"X�%��{��iȖ%�b^���ӑ,K���o�iȖ%�b~�{i?y.���jfa[���C�׬nѼN�V��Uҷ���v(G_�'�4��-�T|�I(����.�L�g8�������"X�%�{�{�ND�,K�}�ͧ"X�%�߻�ͧ"X�%���߂O��Yl��s����&q3����6��X�%�߾�fӑ,K����fӑ,KĽ��ͧ"U5��޷�53WW3!���sY�ND�,K�{��iȖ%�bw��iȖ#bX������Kı/{��ӑ,K�-�s�����
���/�8����{�ͧ"X�%�{�{�ND�,K���m9İ"�ß�D�;����b~���m9ı,O}�K˗Mə��˚�iȖ%�bw���ND�,Ko{��ӑ,K���o�iȖ%�bw���"X�%��c۾�%p#�\�䫇�7k��Y������a,nxK4�.5�#^ z�s��q��{�[�o%�{��6��bX�'~�}�ND�,K��xl?O"j%�b~���o����&q3����ʩK�E�ݧ"X�%�߾�fӑ,K��{�ND�,K����r%�bX������H/���'��ҟ�&�Ѣ���&��	����bH$���}��$��%�w6��bX�'~�}�ND�,K��ܧp��4j�:�3Xm9ı,N��y��Kı/}����Kı;����r%�`���~��"X�q3���$�'�[�Yl#�8�L�g�ﻛND�,K���ͧ"X�%��{�ND�,K���m9ış��Ź�d^P�%����I*vGKkt�ݳd���f�;��]�Qm��6��p���Κ�n��nʐ*�h����+!JK�ua��SK�%u%�bEnKl��6n�6����<I\�ޮ�mWn���':�Lu�{��r�2s��n�}�&bH�d�nǎN� r��u���V�ofRt��	 �y��`�l�����6иLX6��K�h苝�U���$�s�Ɂb�nPLu�P�D'u�]����ݛ�uXx�=]v1��N�N�~���|_:n�fCW.j�6�ı,Kϻ�ͧ"X�%�߻�ND�,K�߻�ND�,K���m9ı,OO�׺�e˗Rs%�d�r%�bX��{�iȖ%�b^���ӑ,KĽ�{�ND�,K�}�ͧ %�bX������\�nk.[�5�ӑ,KĽ��ͧ"X�%�{��6��c�j&�~�w�m9ı,O߿~��Kı=׽�GsY5#tL-���ND�,��ED��߿fӑ,K������r%�bX��wٴ�Kı/}�siȖ%�N/����-�,�Ѐ�-�/�8��bw�ٴ�Kı;���ӑ,KĽ��ͧ"X�%�{��6��bX��~~_�^w�ʖ%�=�hn�S�ʽ�۴��������tT:z�%$>��/��-��&k3&ӑ,K��{�ͧ"X�%�{�{�ND�,K���m9ı,N���6��bX�'N��N�dѫ����ɴ�Kı/}�si�xmAșĽ�y�ND�,K���ͧ"X�%����6��bX�'����󭔲�]��㉜L�g��w6��bX�'~�}�ND����MD����6��bX�%���ٴ�Kħ��?~��;h���-����g?�� �����~�ND�,K����iȖ%�b^���ӑ,KĽ���ӓ��L�gz�䟭u�]�����Kı;����Kİ��E5��߳i�Kı/��6��bX�q{w<g㉜L�g�+{�G-���	�&̝��4Dj����H�UR�*ҪpV!�U2�J𻣂��1U��~����{�������Kı/}����Kı;����r%�bX����m9ı,Ou�mѮ�!B�[336��bX�%�w6���X�%�߾�fӑ,K��o�iȖ%�b^���ӑ,Jq3���++��� 2�s����+���o�iȖ%�bw�ٴ�K��]��Q A�E�T<1U�Y\��B	`)�T%@��F�����hlP��|�bn%���ͧ"X�%�}��ٴ�Kı<�om:R�˺&��ݙ����$%D/{�zm9ı,K��߳iȖ%�b^��ͧ"X�%�߾�fӑ,K��߷)�5�tj�:�32m9ı,K�{��r%�bX~T �:�����yı,O���M�"X�%���}�ND�8��s�t���(��v�GK�n��M��{/�\��nc����������ڷ��ˬ���.k5����ND�,K���m9ı,N���6��bX�'{��l�Kı/}�siȖ%�b|}�~�v�Km�s����&q3�ۻ��r%�bX��wٴ�Kı/}�siȖ%�b^��ͧ"~U5�����\���\r�K�a��Kı?~���iȖ%�b^���ӑ,T�,K�����Kı;����Kı=��-��ɭ332ܹ�6��bX�'u�{��"X�%�{��6��bX�'~��6��bX��	�
���͊�ȟ�~���Kı=��Ѯ��ctL)�̻ND�,K���m9ı,O{�xm9ı,N����r%�bX�{���r%�bX��d?<�����HawBb�^��n��7D!������m˞��<R�7j�^-���fm9ı,O{�xm9ı,N����r%�bX�{��� �%�bX���siȖ%�by����eə5p�\�ɴ�Kı;��iȖ%�b}�w�iȖ%�b^��ͧ"X�%��~�fӐ�,K�~ܦ�34�1�ə�iȖ%�b}�w�iȖ%�b^��ͧ"X�%��~�fӑ,K��{�ͧ"X�%��~캚ֹs5�\�kSY�v��bY��k��߳iȖ%�b}���6��bX�'{��m9ıV����nӑ,K������������j�36��bX�'��}�ND�,K���6��bX�'��{v��bX�%�{��r%�bX�z#�O���BS� �� :�l����g4 mYh����iH�+"� (����@�� �ӊx�
���YTH�R�����$�B0Pŀ
B< $!D{h�"� I@B}��RzkY)�|�Q<��x��!���R��Q�:X+��'~1�D�\<$��|}�dgw{�{��~�n[�p��[V점�m6�  8�7��h���Q! X�eZ �V�&�MR�LW	�l���j�^[ev�U�K͆Gb�Z���<�Kc����U<m��c7�HN��O%.KOB��\��1����oR���u��[Q��[5��R�#�P.=�۴k����Q[G��<ff�ؚ������[m�ܮ�g�h]���]W��N;�&Ɨ���Dhw�ӎN�ѽ�����O��\�p[F^�Ӈ\��.kmme+>v�cڵ�q��T76�J�v�WHүTkaZ����ݻv���Ś.�4n͝ʾ��j�93-�� m�'E�M�\�bU��Xwl�`���k���{%p�9n���`��0�Y���`Y��q5���������tk�`]H��2�n �U�E�u��T�1.��e`��Ύ�l��H#���5/.��kn�,����$V�b�;�'9Y�5�����]S���ݵ'�pa��l�݋���Vc-��m�9&yvΰ��%��G��\��0;��n�� �Y���7g6u탧Rg<���3��.Q�-��v�!���\�FQ1�2�vɗh�2NIm�0�VTͮP�T��/B�.���
��h]٧��-U�	������[d�gt*�,8�/��ۮ���b���0*����s0��H������: �4�dݙ�(m=Wr�Q�-c�8�Mn]�j�Uڕh���n�Z�xY$
���g���=��Z�N��c6��]��ƒ˒��zqI/X:�g#�LXq+�ۉ�FRZ^����4t�:"uג�TsJ�[R�
�]%Ö��۳�e2@im����)����e�`���ѻR.�z%W�
�i٤�ջoP�e���U��=U�Anm%6�H-�vͶVׁr%���Dq�5�e�!�X&�mUw8�V�dGV��v�:��F���8s�n�,�@۴����At  ���8⠡���ly�4�� ���
!� R><A�DTW�s�~�ſ3��m�-9%�Wcp����n�n�p�)��M�X1z��F���T�Af�'
�`���q�볉���!2�$���\��*�\�h���g��\S Yܚ���=t�F\ \�خ3���δ�#u��G�v6���-,��/-��[��I�%��l�����δ�A�����E��r���k(�&�l�l'V0��ZynO��{��y�>��+m'"Wtd�kA[>un��gs�9{z{v�a��N��uX:�ynX��f�\̝O"X�%��o�iȖ%�b}�w�iȖ%�b^��͇�H��MD�,O�w��"X�%��㴷�?W"���붙���g8�Ž���.D�,K���m9ı,O{�xm9ı,N����r*X�%����:ԘS5�v��bX�%�{��r%�bX����m9ı,N����r%�bX�{���r%�bX�{�xf�ܷ.�k&�,ֳ6��bY�D�}���6��bX�'�߷�m9ı,O��{��"X�
X���siȖ%�g�ޏ�����[i�_�&q1,N����r%�bX�}�v�9ı,K�����Kı<�wٴ�K�&qsw��8��WmV�TԜ��q��n��cS�=;�r��83sx�?�w�����3N�s\��6�D�,K����ND�,K���m9ı,O;��l?
O"j%�b~���ӑ,K���w��I+�A;,�my���g8����{6���ߪ�@8ȞD�;���6��bX�'��o�iȖ%�b}�}۾/�\g8�ū�'��Y#��X�n��r%�bX�w���r%�bX��wٴ�Kı>�>��r%�bX���nq~8���&q}�Q�I��iK(�iȖ%�bw��fӑ,K�����iȖ%�b^��ͧ"X���{�ͧ"X�%��O�oMs.�d���r�d�r%�bX�}�v�9ı,?"��߿f�Ȗ%�b{���M�"X�%���}�ND�,K�v2v������f�׃/�om���v�۴����ݜ�t,ɇ��ޝ�;~�߽�7�������m9ı,O;��m9ı,N����r%�bX�}�v�9ı��wߓ����:F�Inq~8���'}�ͧ"X�%���}�ND�,K�gݻND�,K���m9ĳ��[5�����P,��8�L�,N����r%�bX��>��r%��tDT�PDc���"#QE4��hB�4�x;7�/y��ӑ,K��ߍ�m9ı,N��r�;�]�6��a��K�Q`j'u�v�9ı,K�����Kı;�M�m9İ?5��߼6��&q3��[���RI]�A�T�myÑ,KĽ�{�ND�,K���f�|B��������_#�����+Z��ڹ܄��hָ�6Hבz��3�#���.ǷGj6-˿����J�2@U��W� �x�����
����j�{�lr�)K(��7wq`}� m���g�d�*gV]�J���Seլe�� m��Д)��� ���X��c�]r��������[0�ŀ�]I(��߳��>����ȝ#C$� ߵ]0�:`N���I&0��fi^fV*b L��n@��ͻV/m�܍�����\aGul�=2+�)Kaaڭ0��X�u� 6��}!��z`��*���T�w6]Z�k�s�&Cwv�n�� ��ŞK�Cvy���؈���f {���>�f�����wwq`z���]i�B��R�[v�.s��j���,����Ԓ�*�{޼����r�)I(��7wq`˜���������`�%؅+U*J)E�߇��T���^zn��s��C�l�\6�Z��k�	��n̏P�c�A��-�����uH=e�<ӳ�� à�4�q4��vMY��a������L���6�;0R7�{uJ�E��u���ړ�z�(����v�����;�yER��������dM�����F;h����Ǉ���õ��l��gX\�b��5�y.p�{�;�Cp�U�/R{��w�w��w>�*�Cc�=�B�n�>�q� '�t]����N;y!���@#\U��WJl���=��`m��j������� ����g,
�,� n���VA�$�0;� ���t��au�jl($���>m[0ݳ������p�����X@��Lu�0��� m���S�՚`��*/R�1���m0��L �ݸ�um�7v���4b7ģ����a��Hh��OY���U�4]Xܜ�P�Vr�n+]��갮����� ~�[xn���[��8ӕ;�M�U݊���f���Ӽ!(Y)$�f�wf n���F�-nR�R�Z��v����P�M���n�\�]i�Yi'%���m0�w^ I&0ISL�V��U���Ԣ�� m��5(�S�շ��z`�n��ݘHݶ��j�"m�/1��㮧V�o
�����n^\rs�Jx�rVΎ�Cv�t�ȝ#C$� ?n����0��L �ݸY�؆��l,��Z��v��BP�^Q	(UF�o� =�z���ۀj�Ѩ��Q��WKi�w��8 �w�,���HB*!� hU�Tj��&��srO;�vnC�׫ak���]V��qs�$������}�	&A��}�\�Gb�Ki,u�m�۫n��L��ـ�� ���>]V�"�h��$��w�n�/���>m�vg��ݻlVU��P{��{�����̴r�)I,r��z��:�݌I1�zJ���\�)O0��Ř��˻0�:�8�"DU�ՀsZ��;���.$����qkU�R2�vY�}�ӪcI�`rޖ�����l�&�C$��s��\\\���_� ��~0�:�"!�"'�x� �s�i�KadO��n��L��ـ�xͧ� �P�Du��o��\�����v���tyl��Is�eogu�[�ɭ��v����������9�!�.c�&fOd�����lt����0'L� �\���2�FR��1f[ �&0=%GL	�!�u��3˜�l�V���u�muز�����`w_D�'I��u̴r�)I(�`ݺ`�� }����uo� z�V�N]�Ux���3-�lwL`zuGL�w���8�[]�j�7 �[*�=4�5�|�U�J�&� ꣁ�w�;��SlN3Ǡ�{s��RF9�0�C�:Uܳhd��9z΍9�M��t�&	.F���
���m�5ssc���Vw����e��*%;Yl]Xq]�[ۻ`�;�/k���mc�4�b�6˱�*����.$Lu�9�l���x����i�l��ҧd�"����Ut\�/']�T-��;�������5X�Ȝ��۞��z���b�Ӷ���!�r�:���Ut`�X;,���\��n,~o�%􃞽��{�j�l��SeJ�1���0&���z[ �������i�n�WU��Z�X��b�;=�6G�(UG�}x}��X\��N^H;y],� ��v`�ݸ�ո���� ;���;lm�:�+����DG��]��������v`45��&����P��N:��N��W=���7e�������fv��5�#u��Bպ�$+�`{��`M��˺[ ���]F����d����wqd�� H lh��DY`Y���D~�)�g/}�$�������t��q&��y�H��E+���eX�����Ԣg�K� ޽ŀry�*�|u�V�0?��q&����>��7��-�lodaJ�b�XZ�3�ddt��-�N��{_��8�I#��XH�eN��/'��oa����.���%Řl�wwpg}�pk�WT�UYVpo�� ���8����.�W۸�Z(�o+��`�:&������~���O�#�r�F�uY����\�z��SK��>X�D>]02}JL�@�tlЕ��Y���qB����1 0�t���$��b����
1��Z�5�:��Sz�N1��&�060Ӣ����� Oo<X�!Pq ��E>D���/�� a�� ���⩪����i7#���Lur����fk]�f0=�Q������&~������=�=��9e����V߻0=��0N���uGL��pbS��i�Q�ݪtuJ�=m҇����>ю�=��v��Wtt�B��<Ze�t�p��x��x�(�K��ذ{�H:0T���J���n����oGLu�Lod2�R�X���X�1��ꎘ�3�ߩ-�>L�o��4թ�]+�Ț��V�8�K�ߖ�Og >}w�jD(�P���� ��{UKE��t���gu�J'�����ŀw�x�p�2�{~SWX���O��w�m�=�����j�qFG�N����Ѣ8W\��Ӑ�n�L~�>��0=�Q�oGLu�Lur�����G]�[p���Y�K����=�,�[��λ�P8�d�������yL	��`{��g�$}��`l��X�ղ9��
Z�%%��9�%�'ɀ}��`{�����05o"�sd�rR�6U\��]�P�B�k~_�w��k�p�9	$�$�(�IB��"A�b�V�^}��{��]���[�x�W�k�{pQY���ć�1�u�FMu�<���v?�����62�:���֦X���b��Ս��=���ˀ(ٺ��=Bp,�'.��Ɣ��w��=�x4��F�ձ�-��\�\�m��gjE�]N�˹ƽ��N���Su#��� Pm�V�Ts�um;�n�g��Ը1l��C�q��]ӵ2dnM/��w�\\\_�%������֒Kcc�U��!z�m۶����!0N�q�����X�f����	���42�z��[� ߻t�?vw_�.qs���\����ۮ��H���̦��0=��0	�1��ꎘ���R�;y]-�����~�6""!L񵸰�0�773WtF�r�Gex�7�����,~�� ���0�]i�F�%���c����<X��Qz�O��w� >u����ߟ��Lv��ȇUŝ���gN�=��9��.ݴs�٭�N��|Ҷ���ʵW������oL�� �+�X���#�\����)-0���*`,�� #�$Փ����Ҿt����z˲,�XMY��w�}ާ�B�J&w���8���?};���W\V(��-���\\I*��^�� ���`�]����6�v�)�j� ߻t�?w�L ߻� ?w�n w�U��h僭���:yǴn�qQm����Ӹ�j�K�qz������Z(����ʿ����w�w�ߒQ	}!�{� 5wvUd�F�r�F�0~���8�a����7�q`w���$��8ӕ;�M�SwW7SWw�mm���a�%(�(��3Q��@�矹�nnI>�\�7�l��Wh�����ۣ��7�0wT�*JJUᐔ��t���{t�=������۫ذ��� ��y�バ^v����i�����v�ّy��6�>{ruӻŭ��gL$+U�R2�9O�����ո�	��`v�A���^%X�WW���w�|��,�IL��z`��������3ɷlU�Q;U� �v��;{ ��z[Ӫ:`J��ʼSw6]ف�ДV����{��>}_l܂؊RP#j4R#3I@�t ���iZ���f�>[�:ۖ8ʜ��v���� �I.�g~_�w��vـ9�j)�ڪ�4��w:#F��5�	�&��SrF�\���ݬp��ܻ��y{8�t�+�ZX7�>t���odoK`o�K$����-d%X��ŀw��0[���GLT����]�X,�����w��`:�=�y$���{��ذ��a!�W�\ej�L����=����0�S��`oL��īdҺU(����>�,W�k�qp{�䜿{��$��$��$��Z�..0��9KPZ'[-������ۺ�^��7�r\hZ�Vvv���,;��ݽ���Z�\;U�0��Z��$p��-j�({\���	q�C��~���Վ�� ^�,l<3P� ]p�����m��A����T��#3�w`�[c���-�k��
Rb70��d�IjI��6�N<ˤ�nz�,I��4A��Hs�+��e����y�e�A8��b�B,�bt�����w��������V�j臫��"]nHռqnä��7+�Z1s���+���V�q9�(F9m%����t�{߻t�<�K`{a0:�F���+B�+yLwd��#W��`oC�Lގ�Wۮ��2�*$n� ���0o������u(�X�WXe��w�lo������>�I�=��|{�z�K+VZ�J��������lo�ߠt��>���û$D��ϓn�s�i�6������ M̒���ut�Y���������lo�����t����j�:�+���?=����K�즺`v�t������?b�WKT!fc��6GL���)�>�}p���$r�Ѧ�������{�>�� z��U�f��]{�J��r֤��`��L ��n����n��<��yJ9h�dv	���!s�F�`0�j��h�#����aۣ�ڰ[���IdV㭹c��ʉ��������:`M��W�o\3�#e_<$��̼Wk31��L����� �'wns��I��<��!m-�Yjqʰ'}�vnI�}Ϧ�,�E���aRE����D��)�E�%���޸���, ��M�;J�n�����{l�޻�9��Ł�
=
!BU��q`G�M/J����.l�� 't��(�6GLwd:[�V�p�	�1;kk�kq�w�W�xܼ��ݥ8�k�#��Z�X��rv1���Q�l����0	�1��m��U]�]��)�.� ��,��!(����o� =���9��ŀ5μ�Wj��Wy�����`{��`�cw�u�o۸�Wۮ�-�n�hG%���
"g[��9�w ��,D(�]q�q%之����0�?d,ds���Y��NQ�l��fA�N�� ��d��Q5j���Z�r���]������7fD����%��gHӏ,�U�:iMMZ�ŀ>;f >���y%	(��y�b������;k(Z�IV6d����0&�遴��֫L�er�L ��n�z�\�\I�w�ŀ{��0�v�el���:�1���:`M��l�0	�1�����䵒�Ф�Հo۸��l�޻�>}�� ���#�uU$zD��@�'ȑQ
hj!H1�0"�F
Ŋ���xT�_��ĈAO��U= G����{�t'�AZD! ��0� �����:�>᷑���u�@ Ef��*1�PYB-j���$,<U&#W�&��A!��kVS^��u�� $8pm�($�h   �t���K(���"�	 �_X3"�{h9�hf��a�dv4�v넀�e�(8��j��>�9�f��8%��5l�Rl��������]��uλ=Xk�q@�X8���^�8���w3��Z�b�g[u�ܤ��	5Pt��k�b
�禲[N{.�['1��K]Rse����؍Ջm�|��]�Z��&۝!ļ!�n���yb����B�Md5�u�MZ���B�X�7���7/Q��-Ց6�EX�L�!�U�[F�O6�ۦ��#՛�˛%�m����4��ly$��l8���K��#Bv�]�ni'�P*���jѺ�R�.�`�"�E9$�͒؜��������~��c��Q�U�8�oh�-��nk�O۝A�,n��5���1�#.M�"ԭ�N���Ǯ�&�V{E��10h����cE�z�;f��{Bۭ��\�j�2	���6	�T��1g4ƍ��,l��Ψ΃�r���sm��/+`ǅȗY��#��*7n�d���ڌ,�͌�-�#�Բm�Im��l=�:!�லvI�R��'��o�ЬJ�7\n�չ,qXnX)J����v�3�c�̖l�;k]3փ�t�m��$mu�����p�PӑV�5T��]R�g�"�)���[wb᫯L۷FqKmVmν���v4Ǘ��O�9��DIA�kj�RKa��'�b�m���ۡ�q@�q�౐kj�v�Zv���si"��@�Z�㇖[q�����c}�-F�����2Um��I�b
��uյ��a�m��q[;��IP�UU���y�i3�sr��'`&(j�+Wv�7\�Ny}[��moU8S���:$�Y0�2;nٵP@Tj����G�1T-U�Q��e:(�v��N�����]�@�d�_�����;-S��,��N���s�*��^W�ز�'��2�w]nx�t��R��WJ��� �ȥ�~=���~}�{�0 Ý:(	Q��SB9��L�сC�/�x>#�CS�T3���34d�dʶcb&Bٷ	/;�:�� ݳX:yk�oWt��.մ.L�m=`�.����~�~ݷkn��(��g����fA�5�#rfۇN��vͶ��s�3�m�i�'9ɚWTJ䎍���].K1#n��U�p;�); ׭���C��
���|��m��q/Q�<�8-�9�ugd�u��gv8��h���ל����yګnK��s�$������~��X����[�agK�G��=&��û;�ubB�;�:����|q���V���'%���?���wL`zr��dt�%l��˶ʝ�������q$�g���X��� o�l%�B�TwQ��(������jf�� �>ŀ>7�(�������n���w��m$����`���� z��BS��ߖ ?/?H�N��mc��`��X���׻���[	/�5���:ų7�dՋXܳ��n���$��r���F�I��=���J��u�Pq�pŎ�ɡ�w�m��c�(�:GL	::`{{!�x���Z�r����Xq,�Uw�\H��Q��M߷��ŀ��z(P��;�D	%��V�%v���b�$��N��GL	]ѫ�ʳ.����T]����Q^��� =���7/��ŀ��tr�*v�nJ�t����:GL	� �?J��)�*R�Gk���X�RD*l�v[�^��]�[F�K��6�v0�ˑ�P���gΏ ��,��^��G(o�xY�;�[I/,���`��Y����m��z����<�o��H�N��m�l���n�ŀ���MDAs�UCK�W�
.�)u��y��ذo��g݃���W\,�R���芯o�x��b�[ŀ7׋ ��n�V��Ej�r�~�q`��^���7^���� �u5J��bi���ft::7&�8ۅ�:w=ۛԥط7]9#��;˛��(��ۆ�^��Θtt�'I�	�����V�X�,�H[V��ş�\l=���=�ŀowq`��]��ʝ�S5V�����a�3�w��ŀ~��Or29�mq�-����O��~X��X}x���HH�
1 s�UM����y�':o�l��^Wk!*�7�����&:L`M�t���t�����$���x��kt��Ш���g�=�i��׌���(���$� ��������:GLF򻻗��b.�h�����l(��{���5���������v��V�VEb(1�pw���[Ň�L�wq`���;�:����B�Z��`��X��L ���~鸰]���+%�)j�� �{���n,��XBO���6j�T$	l�j��m��\1'uY�-�����$�ζkn�St�X�h�È��n�q�M�'����v�6[�MOm�GS�Iq�m�T�c`yK����:j@vٖ�]ګv�`�8��T��-��rl��^�	��4o���_nv}JMnkum�:,K@si\����(m!B��p/1�U����cA�v#��Ď8���q���@Q��ۮ�����w��{{���r_�vm;w�Jmn9q�Dvݞ2�pFݱ]W1��^ ѱ�svz4G
�!�i��TrZh�����Mŀo[�
0�l��D񡓿Qu%ME�������f���%2k�ŀov��׷ �Ӽْ2�[Z��BU�owq`fA��Il	�GLz�$��Yx���x]�0&̃���x��(K�o��,��j��w(���\զ)%�&�0:H�6GL	��H�ߚ���J��oo<�f�i�ێ;]=�՚�;7On)dk\�����G-�7���GL	�:`r�[�έM��euX��-Xww4�_�""b""!.�!,���`>�� ����;����*Il!!mX�w�$��GL�:`�E��ŖJժ�����D����7�n,��X�0=�p����VY�),�`M�t��#��09I-��RKx�.6�B*S�u�E��6k��u�LAGIۭ�ޏ81�����Qze4�7��������`���;-���Q�==� ��m�GiT%D��`��,�wf7���GLF򻻙���]b�Uk �� |��a��P�� P��b��!L�D��.*	T%ĕsy�� 淋 �r����U��E�(�����Q;�o� {�� |o׻� �����,��U�NRՀt��l�������t�=:���S3t�$��v�y�u���[��Ls��g��ӯ�a�6T?�����[���fex��09I-�7���GLWۮ�J�
�UG$� ��ـo�#�I0$���T��-Yu�U�ک�����,5DD��w ߽�w��l�r�h����`��X}x��n�.W@$ �!%���g�}>�ܒy����,�*��/���09I-�6��,�	Ga�&���܈�� ���=l��v���G��]A�X�
5h(�:P�r�����erI��dU�ʾ����`������tt��m�W�����yl	���$t����)$�>�Z�C��Ub��`��X}x��Q2�wk �鸰��ɥwfw�e�ffSN������������˾=[r�eU6� �$��GL�:`I��՟����z�m�-9%�Wcp��]kۗ��3v��p�*�v��Ȝ�XVݢ\u9�F��=��2(��[s���d$6bUp.�nB�
ٹOfx�S�R�F�� �<�I8���ӐSf2�v��8�m��q��kYtt��(�3���v�1�ڒ�G�\�J���q�Y�x��#-�����ݯ���c9��I��E�r�&��{,u %N�pj*�b�Uߔ�g�f�f��Hu�����Α6�e��&��P��۠L�j�;X僋)�NX� �*��ݳ���,���tt��$�������yW�+��(�X[x��S&��X�ݬ~�qg�\�9��wV���P��I�����)%�&�:`t��Q�\�m��U�ʰ?��q=�����|��GL�0=[}fR2�]jªj� ��`�JI�����ŀu���w^�Xܶ���\G%�M�t�[rlZ�^���;<"O.z�=[V́1��;c"�	�Z��ڨw���5w,}�:`mt�]ee�R�ĩ#3�=�߶o@�$�X�T"|PR$"�w����krN}����,�(JUG��왕V]��j��� ���X�cŀu�� �;l�?uu��GF5k%uGl�?oV��:H���)%�7��<��/)]���Ԫ��u�� ؈�O�4�;�X�k�X����cq+��;j&�r;�L㵻H�Z�u��-��v�0\V��n�GiT��)%X~�� ��ـ}��ŀwwq`?�$�m�"��-x)%�;�GL�:`{nD��߿~H�پr�V;��#�`��� �������؄Yą ��Z@�[���P(��s��G��|7�Ȅ*:�c��U0�(�\��a F""�"��
@�1兡BGP���!B����!F�ĥ�	(�'� �D[�M�4����0�o��0��R,F$B����51�X@��e�ϯ��V<��q=ߋ�u����Z�[��6�BH@�F��ւ]C̛�Vg�a�ϔ�@"A����0bI���R�FFF���1d"�X�H��L_B�!�� z��R�? !���>a��! G��Dt��?"IR��BQ�"�n���v{�X}�֦��8�jJ�Xˏ}�~Xݞ��:�v`y=�~�����j����EQwk ����P�:�����,��� ����jr��XV+e
��d�;k����ݐ�"�=���e����pu�|�	��YK+*����'I��Q�t�����v{� �V���tcT�Wc�� �{/ ��,�Ss���lD(�I*���c�3eթ����*�`�{ˤ�:L`w0�P�%�ee��x]�0<�K`��q��'9���
V	�]K��ﳫ ��vG�؄P��d�`�w�zCcߗ�k�ŀ}=n�5�[�
�a}=�R��뮲βrkku�SW���G��\tA��ר�C] I�kd+�`w0'H���[ �&07{[Z�C�8㉩j�7�������Q��z���^ޝx���"d�tܶ�XQ9k �`=�� own�tt��#��2!^#������n�TL�ݼ��,��X
^��o����/4���حR����׋ }o������ �A ����������ѵ@[��!e�Mƺ�F���G�:⶝�N��;^6�x�s�n9���d�g\��}��O�Q�z��")�
|�W��u��v�����L\�s	����v�Zc�D{/����<L��ٵ�VrX;V���c��F2�1�l,�`Z-��=�'c�c������=��xD���s�<� kY�ɞt����ڗCf�r�b�"��kv.�����}��n>���^�\�RƑ"����d�n�v���s�a�QLj���9��e������Ilt���::`ڴU�J�uIG*�?>���6�X�L	�0;ye�2��0.���]� >7x:��a�
&u�ŀr^�7{ ^eZF$�#
�������������v��s+T�&WJ��fSwGL.���1��Ww���nGK!iS��KY�un;m����wku�`@tv��G�}�Ǟ2請u�`��+�exSנּM����{�ŀo�)�¢���J���}����� ?b�z��p{[�L���L.���ʖB�]�Vef+K/1��]0'tt���-�o۷ :��67K*r�U%X�����[ �&07����*����%� ���0?w޿���,{�ŀ����JYm��B�F
�nٍ�M���v$���u��x�c�Y�zC��H�v +"��-��=�z�uwq`�:`n�D���y�k�XW���Ԏ��:`yt��&ɏ��7��/&��i�4ӊڰn���߮�b���X! 0��;��Ͻ���V�,��n[P����rZ����1��0'tt���e���6��ժ*�� ���׽��=��X9]s�	��Bwjf�q[i5n�o=��Gg�>�������'���tb���Si�K#�e�v[�~�n��7�07o�`d����-,2���^WyL	�07o�`d���u�I����8�uZ�꒎U�w�|�l���Ԏ��:`v�˵qb�1YJ�� �&0=�#��Laj">��J2$!��8�s�rw�ߞ��ِ%����ew���Ԏ��}���;�|�I1�ߴ�E�����d�]r[rl8U�uc]���=�%�T��gF]�60����g��*WY�L���ݾ��t�ڑ���7-�UB�Z�+-��N���c�R:`t���H�O��Ve,���j�������}��,=3��� �f���˭;�m5	B�ݖ��Z�`�� �+�p6gwv���S6YT��R�*�7wq`};� 7wnI9���7$��ȂH1A>"U��?F�y�,p>�G��_=�B=ֱ�L��Z�o�wb�5�E���8O={urb�IZl��J�t+��n���^[-�nӻv�g196�t�7K!h�cYX��;R�f����.]N�]�ך�n���w[�^pN��z�b�|I!׌b��嵖܁p0�g<6
*h}إ�g=n��<lGG9�2[f�� ��{�~��s��l�H�@�B��KW8���%��{���~�o�L�n9z������AֽN�؄���m�����k���z�z�Ԋ�UWSV��� m��>�o�/�{��,{���h
Ȫj�^ l�ڑ������?�I��v��[n���n�W�� �����.$�{7� 7���>ٲ-M�%�i�xfS�����0�1��t�����
J�,���N��?�׷� ��ŀz""�����ȝ���I�<�ׯI7Mu�u�ƛ��7h��$�62nnMt�p.a�a��V�J߼�޼�1��:���_H>�� �;�4�#�+	m�?}��ϒ_��`� �GT*�R bEU�&GL	� �$��������)a*�7wq`��L?͞��p��ذ�ՠ⣪�:�!eXod�1���0;�t���j��@b3(U��`$��Tt� �ݺ`=h���-��n=`x#]hۣ�c���Q ��q�hy�v��U�]=�A���-l��\t����{���`v�A�l�.]Ԥ�]�J�T�fVe0;�t���l��Q��{��j����ڰ�;� >m�:�""V(Qj5BS5�.b�7^��>��U�Q��!,� >�ۀzuGL�0��;'Ɂ���e	�(ŉe�0=:��t����0�v����2�eh�+�2r�	N��ts��hm�&�v��G5���L�i@pR�\IR�#v�S��Q�*�ｋ ���X�����n, �uh8��uWm,� �:�g�D�wwo 浸���X�,�W* �̡V,�`$��TŇ������`ݾ0�]�=�\��UV\���lD$��I%]��q`��,���$����%��/ ��Z�NJ' �N�j�;��X~�� >�ۀ~ޭŀ��6���*�:�ٰ�M��[�-�J����u����J�܈^�n�q9Q�P�(���j�;�n������z<���(7wذ��aJh�UJ��(��X�n��"&Nk[� o}� ���Y�&γW�~�6�eV;���+�L�0I1�oM��e%N^Yk�J�?��I��,��, ��x�k[���hM+&���N�;V߻���\�{޿��I<��vnI�UPU� ���UPU쪠�� EW� *��UAU�� "���W�����"*��
�
�
�"� *R�H
�b�@R�
�Q *H��
��""�
��*� * *��A *���D��T`* `����D�� *� *��A�"��"����"�b*��E��@ *P�,E���AU�"�E��A��E(�`*��"Ĉ�D��@ ��"�H
�  ���b��X
�V�"*R�
�H�,�  �� F"�U",U��DPb��U *A�"��,��A",@��Db��`��* �",�A� *��UPUʪ��� EV�*�UT_𪠪��UW�*�*��UAU�J�
�� U� U���
�2����؀������y�?����	�| �� (    QK� � 4�   �	�π  E"�@�$(*��T *A   H����T(    �)@�U
��>�@  ����� ��V�v =���ɣ{�����#_s]>�==����}��7 n����O��Lg{<��s5�˅� q��L��t:��  �(����e37M�N.���p ��.[�����e^���f޵9���:�ʙώ�{�w�{Kɾ��hf`��=^
��Ifϭ:�}�6O[��P   �8=�3}����FN��=r�����st�vwj�Y=��}ܽ[� �}�L۾ܯ,��w^���s�^��
7��\��\�;nf�[�R_p�#-+����z�ӯ]�����|  UP  W �W���V��w7���O�� 0 �@@��Ҁ>� �A���� �� ���G �'AJ=�@�:Q�@��
2h Y�R�wC 7w �@� 6}����� (AB��>�jY�8r{=>�����w�͔[�{�y�v܃^����%��d�>� ���k������_z�GF�>�y� i��s��G]}�|���t  4   
�4jI(��O(h�hjzj�  jxI�(�A��  4� �z�J�� � @  '�T���h4�  �4  5?Q�Ē�        DSDi)D"z'���6��I�F���O)� }G�o�=�*����M���q�� ��fS���Pv"������?܇�����: ��?�����hn,d� �����_��4�� ��H���G��8}?�������������m��m��n�m��m��om��ܶ��n�m��ݲ���333f6�m��m��T�m���{�m�۶[n�m����};����zz�m�m��m�ܶ�o�6�m��""��$ E>���TO��@>� '�l�O�*�U>��UEQ�(�C誟Ar ��T>� }C耟EP�(yD�*���(D � /�G�(�@� �EW��AQ�('�U�*���
� � ����A� &EW耩�Pl~�� 芩� �@S� �AO���D~�{C�?}߾����s�P��І����4���
=@�����D�(J�uN��:;�O\_��n}wI���CI��b�W"<Q	wT���N�4(N��t��D�i~��
�RN�
9D'FE5BJ� J.
B&Af�Σ��SJ*�o! ��#�����-4�(���C`�}�If��k� �nY�pb]�v��5��8ĉ)w�&�Hq���C��33<޷�X��0�[�z���p,*<w��.����L.����c.Ü$BD�<�>��yv��aHP��H4#1$k�Z��]�/<�!!/��P�Aс]3^�9�af�O50��*ˬ��4bD���.��^>1����{��,HÆ�W��{�4�=���y�\7JB�XB�"D�����d1����\�}6 �Z�.T�T�]M�pw���B�H�	Yu�5����/�ԁ(/��aR1�SN���SA��LG��5����� � �����=�k|<��-Px��>:��1^��c���:�j]xˆ�>=�a2�Ya����0���5�E�L�1{�#�u�u�Lu-3F�(o�s���	�ȁ@��5A'��I@�b��Ccl��2Vj��5H��C��m�}|B,#X�`Q"�`E�C�֞z9����B�m�/$�ͳZ��恌J �2�ro! ���K�ٴ�OB4"p�y	Ow�{�M`ŋ��J{.�$�+�Ѕ�]��M`F�	.��h��
o�秦����]��zE��\�.��{��F���!�$+�"n٢]0���u3`Js�,�� HCT�Y��!���d6B�� ���)+,����=�!r8�J�!�g9#$#���"BH�4 i77B2%�,j�@�p1���6�iLI# �A��!bh�d��l
JD)#�߾Ѕ�oΈo�5��t���WH�So�%�m�,���рC�BJ�%-��5�M�7[�kA GNėY���s�3&�7�M'h��7�aI��l�H3A��f�ɦ��J��!�E�d��V2��vx��H��(Ʃ�� �%6��#2y�ѝ�=ȉQ� A`���x��C�BK A�i}N��;�$53�d����㏦͝:�A(h16�On�� �t�l��%�*`�<<x$nq��x:A ��v$� Wj�L�b��� ���}�&7A�!YVB���!a�����ד3 ��
B�K3|��tt���V\��
��O�=�f�ᬇ�w���Rmu{л�9m�0"B�}<���^n"he��RR0`���(L� ���=|�ނ�=e+��f�N��d]u�S�J�7zT$+�H֝��}No���Q�D�j&� �eu���>{��G�T�4�qJ0HC�l=�@�H0!���0�4"�#�P*�,�at��h@���U(@�@4�) ��1"T�T�
Qt!���3S^Fj��'�`I�� 5���@ŉᐮ���x�Hh!uB�vE� h!M�B�HD�X�*:q�b�b��H4MH�
�X��R�ry��Ä<܅��Y"y�:�<!: Pa!	$��x�sP�s|d �$aM1�������!E�<6u���|zS�tc��s����/�\��Yŭ�YmJ QŭP��d�S�
D��
k}�MbŪF���M��`��n��ɿ6'�>�w�ӛ��	u�6����f�5o�S��X �s��������x�N�p�B0)�1��!u��Fzā��38��}�'@�$H�[)XT�XX�(D�)��(B�]Ze��$�(˩t���.�tR��
���0���aB�{�4p6w#<I!	 D��"�,rHV0B,Q�B"VIs�y���9�;��\0��y�s��͸Iz�o� đ�N�әT�	
�L�(B-� �D�E�Hp9ژ�Q��@#P��E1�z*@��w���M.��l!SC��&�vWP�hMf&t0J0�1ˀ�14X��-͒�-�@�&�y�HT#`���F4�����(J��1�]s�2n�;�FOr_��CE#b�D��	���N��CP�B�Z5��xH%hJ�Aք�w�x2��Z}�wz+����s:n�8���tbJ0��2O82J���`�љ��^l	MCN���2�7�����Ӈ��x
Ca�a��8�7u'�4�2$�ΐ�*0� �cSf�ﭸ_}4�Ji�M&F�w��<�&��$�c��3!XR��Z�5
��YYM*�0��X]���3XBaXX�L؅)�$5)�M�!�Ͳ��0ta�K��!��љ B�k��n�<Ä�"0J�! �D����]s��ą��Xa�c�@�f�;�jK��"�b���SX+)	��P�l��>h��y�:z��F��)�B��@b��@�B&���<�уJh��%��D�5bZk�L��]8ְkMa�1����M<5��I�����!M$�C.S`�1.��!m|�9��W���]a�i��GN��ĔHцQP߄��5�}�6N�_d��D
��ѢB4n2�|�/��@�%H�����@�M�xyO�7���$�a�9��Ѡ2�(i�5*���)�2�a!!��ŀ��@>>��(G��$��0�6�G��rz	��@$qv���ټ�w邞�ȕV	��uW9�$�d$G	|me�	]$ � �b@h�V�,��N�y`̹M<S���e%�4ˇ�i5����%e�7M]��Z1��؅�+
��n�HT�R5���1�F�`��a9���S�b�k���l^3F���a�tc
h@�liq"�M!�U�J��0Rc��%���P����5f���љ%y8T��S**�����t�2@��F�2�A�J�+�H�)��m�Q��7(v��<w�}���d|��I�����n\vU�-}�E�kf�𐊄���eU�t������ȩE!0(�*�Q���#�A!$��2=mP$��-|��ϯ5��I$�I$� $              m            m    �P��` ppm��   �` H 6�  m� m� -� ���          |@                                                                         ��,��n���$�5�ֶ�W m�hA�]nm�ֱ�m�w)�� H���F�I��\��*�9�㳳Q�k�l�1]���e^�K�0U�����<��؝���<�#�&Uc�.|�YL1��KU[�E��Nsh�qh�jc���O�vM��W^�6���g`���F���������QE\�:��Z�^4�Y|�|�}�E�M�`>.�}t �@Um[T:6 ڴ� 1���A�5r���Z�&��ӥ�r@�u���
 m�`'W9S0    [@ ��j�V����p��T�Zٶ*krڪW�Ca���٤$M�S0�5T�n�;m�1��d��ݥ���*ѭ�v����V�b�	VRP1�V�jjlH [B�Ҥ6�Z�qA!Ā��f�N`��\ 6��m �*�.��MUu{$5�^�}�@ �e��.�L      p[%ŷ���� �� [ԑ�E�[B�q� � 	���lm� �`�[��B`*�j��+[:�e�F��[%�k�t��m���u��  �m�����Nd��Y˴�`��m�m�=Am m-�mlm���Zl $�kh
��9�&f�*�m�um���@ mp$  hHm�:mr�ڪM�	I��	�ā�F�u��A�� H-�����mm�  ��o���6�ޠm�B:I�u�l/-��J�UR�&�2�O<� 
�*���m���$�m"��cEդ�[@  I��-�ӎ-�ںJ�Z����G 
����q������e�Um � l [A�l�kYλm� �� BF6��[[ltm��aB��6lܛI���ܾi&������5@A ���
��Z�Nؐ��m�����Yy(e�v� ��imԛf�h�b�  �I�RF�a�m\� .�-����r
�mS@,R�+^�0��iv�`��[E����!����*�Ի2�C�����m��� �c\��v�r������Zi�qm�Y�Hmչ�N�   �T��b���\.rʵP�� #ykv���H-�����]Q��eݐ:��ɗqa��gc.�[�N�����<.V�,J����V�xs��ZU���*%�&������Kh�l��8�iʙ 	���2P#�#m�f�h�a�   8�  �*m"��mL�ŵ���i:M��m�z��m�nv�V����v�
�U.���� �|����҅-ㆬ�'m<�ՌX�UU*�v�1��k7m�����H�v��9m��-�H�-yn��дZ8�\��=[lXe���۶�8�4��q 9m lm���ku�z6.��y��宺����86�� X�j���^�8  � m��P V�K��ku� �4�;m�m�  [@��NH ��mYƷ�B�㐝8�@���m� 6�G-�|�v��l�H-�z�K5��v��'���Z��c.4r���/$���,� � kg]C/n�����Ur��Wm����Ȯ+���Ʊ96��4i�e�-��    �K٫`Xd�{}���]4��$ �h��,X��!� H m��qؠ��r�IW 86O  ��ք��v�6�j�-3I&ӦAm+m��6�     d�"�N ���j�n�9����n���%�f��M�  ]6�Z��a [@ ΂%���6�A���U)(
�dڠ��������F�
��	 ��q �p 8�Mk[Kh4PH���äv��ױ��{t���� =U�յ��`8�u�p�Z �$I�T��%�\�� 8Hm��`iR�m	,���KoC8���I O���:�0L��T�0�+�J�V�+��w6mKrI��8����Ij��� �v�(N��cnl� $��W�������sŷq]R���N'��C�������KU ���*�����mNR���y@d�vZ <qm�Lå����` Hڽk�H��[[@r�+rʺ=�zGUUJ��!�z�i�k@H]:+[!5P�[����8:��}�H1�f�x89�ڀt���uy�@�;�1���elݨ�m{6R�'Wl)���U+1�����` �-�0����I ��n�o$�s���͵�Ė��$pm��: � ۫v�`�U]����� ��6�۝h  ��}�����X`54�� 8ת5̍��@  ڶ� %�� $�Y[l�f�l�7En��Ӏ���$�$e�o4�m��8��m�  8   H��m     H  ۰-��`m� H �H��mm%+��$6� �m���'Kh6�mp  ���!�8 q�� 2[R 8 �mrڶ�hm�  8m$ ִ�    � -�6�E�z�o��}-��F�-�  �6� l�����08qm j�$�m6� �F��I�#�m&   $     8�m      6�$�q���n�9��H h   ��ɀ�e�At�m�"@ h  �        ��p  i$� *�����������}��fd�.�m�n[�N�$d��+�ZN��m&$�  G� ��6��  ���`s��p�6Ir�ֶ�t崃�F���kh:A �[oZ�Hl����7&�m HM�uJ��J�����m  ��oj�4��D��/��$�-2� �n��Dy���-�PP�  ���d�g-�]�� n�	  �  6ݎ֤�6�;`6ͤͶm%�u�3l H8� l�   [m��خmn8s���}��}�{qď;��
����(���  m�p5�@�n�-I�/Z �]68� n�CY��: �pI�m۲@I:���� $�h�f�ۀ�1[n��ʠuWUT�"��m*Nm:�"QJ�5밁�qJ����W[d���d�8�6�,�0Ż6�m��m����`2[N X�j�  �X� �ci:M[�� ��*�$�PRE�$�܉:K��[$�i�<k�����U궫��Bʻ��J��� 5� 6�n[@   ��-��"Zcm�� msm&8 hm�u�@ �l  �ݶ�n��Γ�-�*H�  �IYb��@ 	��5���Nh�N�΄�5\��Kv6t8�P5��J2�[��c���cb�����0$��'n�=�{���`�hi� pV� �@VJI������$�:�%j���7�:*"����{�"������
k�VEk��៭,�(�� ��A�DB�  � $A���F�-,$�a$�=����� �¶�6�,���h�!H)JQ�(U��� A�B�!B�! B�!B�!@                        � I$��B@O�P����(���������G��_�^ ��M�Q`"'PE�*PJ� g��@���S� <AG��<8�TP�(1j1C�����on����Pn��@�B��A}Br��Q����t�@6
"�:�pV��Á ��y��H��!�DDꯀpb�X��ǨޥB�*MT<=��t=I����t����O0/6�d맃����G�ڈ���'v!�Ch�b�M
�� ���]/x�����N�(����8�p@�%��j*ꀄy���ԋFW@ ��z�T���@
"�#`��_<
+�A����uE��Qг���ҧ�*���S�T�A��    @    !                                     �Q  �$� �"@�g�y���>���������؋'$h�``"TH��Q`(�B��H�`�E@��U*U`��-�TZ@bR�ڝ$AL�4=,�l��� �Nh6܁� W��h�$    �Ȱmq� l�6�              �+]�mY�l����/j�����-��g�=Y$g��Q9;0�\ڒ�#X��Z���Kԩ�m���mn0��ێ�iT��@������;vq/2���NKcj)T�n������mNb�6+��j��jP�RsT�� �12U�H駁oe+&4ع�n@*5���x����S��*x�u*Q�;�gls��G8��[�쎱�!꣄�s�!ٷla�v���v;g��@�� �l�]-G�l�R�g^�R,��VXB�.U�K�5��k�/d���0@T�zi����I�D�UΌ�'���'�%��z(z�)���_>7F�m����::r5c�����Ʊ�D�˳=7j��J�8m���
��Ű�E�b:����<p���)	��Y�:����'��Q�nAQ��ѴrL��
�X���ѳ��bx1��6����VC�ػF�Ԗs��{b^Eon����W:��z��cO�L���u�V�X��G#^��[d�˱��u�N��BV����
��c`|�F�<D���R�����pd6�MXm�Y.�j�Z�
Z���̹�e�ZCm�� A�lj(�z|��z;��#I�1�đ�૫]���8�V���1�.]��Fg'j8h�D���e8gf��/�����:�9��qI��Pˡ���q����c�����ې�%*2����8��T�J����H��t�����6���߭�o������g���G}������̳1�zqC�*{���p �'4��pM(�臈9Á������c��u��֍f`ְ  ��&�n;cp]76۩������	�Cy������X	�sX�^@�pˢ��P8�ݭmgb7�jq���"'�r�d�.6�<��:u��%�n�	�i���[��t�XL{��摔��-��ŝ�[�w<�nq���Ź�4�Sr��1���+A�ۻ߯w}��}��k�8r�T�=�r86xۄG�l��W����M�ho�ZCYn�÷AnxLA�1se�!�"���y��OÖ��/=_�wۤ�H�q$�2֞_o �ׇ�y��ga���\<�͂��^lk'z-�	@ʌ����݀v�`���ʼ���4�8�F�5�F`Bo˹����f�8�9�ТԄ��b�\�� ����XC3��Oor�z5HL���C�{:Q�q!��q<�OM^���}�g��l��	�$$�
U��]̜�W���ǝ�7�h�P�߶�݄լ<��^�9�)2\�v�`�Xy;{wr[|���
���M�ˣ>�۬rcy;v눺+� �k�c�j-�[Wb����P�-<����� ����̆�P��yW�w2�݃�y�s0���̙��l������tJ��|��9��:l��FDJ(�-�;{�U�<�����8H���jp���������wr}ݜ���E ���TES�nC����3/j؋�8�����/o;�\�Ռ��s}w2���V�w��⍵m@K�;z��Z�y;{�VqH��d0�;{�U�<������wt���"(����ӤU��۷�|���A�y�)�D7{�a����Z���L�Hƹx�\���hssf2 ��{��KH�E�b`�@�ݔ{AN�u�yv��mv�_k��G�j�e7�'�o}�ov��������8K1'
8ov�����*�'0�n����|p8�2֞N�AW� ���]K0�a2F�i���^l��ov
����7��mF������Á�}����9��|�4�%Itx����""Q���i4hX"U�V�BJQ���j�5S@��M0t��r-[��}�w_f�[{w#m�  �ݥ��Uv�[-�x�F�ά9�^�M!�\��.'x
Yx��87�$�8$.�Dvv�5ٝ�r���m����O�fA�B��k�y�G=]m��[c��B�61m\ٮ�m����n��)�1fu*��l��ܹ�:ũ�u�D���7LDhh�s:���}>�tl����tr#�6�ɱp�Vsm��4uŶ�E�:f����U��U�}�j���.���)"(���qi�"�6߶w킳8%����fl��ov
���v,=@�n�JP�� ���{�^{�U�8E^lf�,�Rr���Gm��^l��:GE�I��'
((�y�;� �k�.5.�dݛ��B�u������_Q��;�O'o��<88F_��Kt�L1HF��fzN�/�@r���Y�Z��鵹#iF����݌��u��0�֯b��m��K|�\k3ނ�i����wt���"1	Ioz3r�`����o���PՉ5p���vgv.�e�:D6Vs���c��f��F�a���8b� �b�/���3v�0+�-�E@�nt2���8!��Az��]��w�b��	N>���k
.h#��䜻܁�z�8�o�5R�b��w�:���v
�Y��$JHr(yY� �Ǉ�{�_Vv�+!
2R��c��{]���Xm�vL�+A8xT���V��rDK�;����*�K���Y/#RF@���i]�#�r�<���-jB�{Ŀ��#RJ��	w�W��D]����q���9����+-����8��T����z�׻�f���;{b�&�e���= fnA]Xyw� ��}���v'��q�;m6yɱ�J��n2�TV����	�C���C���+�.��ޛxa�G5��o�5JP�X|9��y �.�����ȻƆ�e�QJe$%7<�܂����ua���܆2cNH���wv��z���ntެ%�ԑ�&���K3q��1���]�֗z�o���z�<�m  ��WP�%F8N�5�]�;bw4�����z���%�o0Rnn:rc@j�2i��C�7��:�+����c&r4ơ$7Z��v�!�,lU��/Tf�:�v��L�1ݰp�ms�vŌ�֋��;�v�mn�W�o&�
5���B�CS,��D�]Q�Tbڍ��B2��w�]�z�u;�k�c�3��@���������6�t�4�Չ�.�بc�n�l�9w��nc�f�Yۓ$�\�c.fnAYy �܂�������m�C%���f�z���n7�`bq�Jq��3r3]Xyu�m��A�F& ԅJ���� fnP�`��.��r��Ip��F3	�n{uV����]���ʌ��ZNa�;���|o�\������[�o�� s���TJ�����l�}��� �	��1!u�`���V��^^P�XK�Ԓd1�7o%������V,��I�%Hъܒ�mi��\���3r��\�(U#n�����۴7��" ]��������k�t������_lM��h�n�c;Y&�u ��L�T	7#L�:=�ހfnAެ<�ۃ����D�'��37'����7kO3<r
�d��u��l8�����K1�_ե�?[y9��kZ�����aY�P5$ +��@��4mBY�dX�HJc�@�P��� /�J�"�M�rP<E���"衉ᡰ�Q��ᄑ�� 0"D��R!1�HB1��`F##�a�ZM�;#1�# !���b�A%#pw�f�-䮔Cp$l(�Sʣk*�<�q��Jfq�Ԃ_45�w�q�����H@�W������^��J���?@~W����T�|� G�Z�:ju�:�����<�i�Q�2�5JQΰ��[�֏~@@ƺ[9�Q�%T�JG`AZ[��5-�B�,��� ��  }�)�!NA8�Q���w#V�ݒ�e��k��%%����Y*Ljų: ���9�6/���ƃ#9��&R�1C�J��i�܃��^{'��Ți8��\?���v�d<�� �+<흵��NH�%���<Fo�Q�-#�!��B��F���߇���z=Ω"�QH�ґ*��<͋�Xc�ۈ�m�V{�d"(�"�B�JF�񱍪e�������9V%�:���[G����	t_��������\�d��0��aqG iȡ��k��݀g}�U������[&4��}�7|�������������m�-6�y�j�0�g���y��/����Cs�9m����W��v��|������$��>/*����(�rI  :s\�;e)Y����tz�����f:y��O8Q�'	�#&{E������DW,؞��#��gj�
�ɲ�Lv{6Q�s�6��[��Z�9��8��s�s������>����9��/&똵!X�g��p�,z��jzp0[�����j�ۂ�m-fq�wu��[�vƞ��w=��>Iwo&n7l�.�m�r���qrD�i���g�R�?7? ���o�Z��n�`�T9"��J�����P�Zy89y�g=� ��AG ��m����\~�f���l�È�#�2֞v��܀^nmķI��$�P�6�
� �o��Z���l4�]��ͭ�G��ݶ6��Ӡ��ح�t�N�};��T��J4䋎>��zy�<{�O�  Fo����28�H�=UR�3~�W��=�{4�w�/]�hCs�9m�����k�;�Z�"�Z�����P�n2�����j�ov
 ��w��3˿Z8ʁ��1�R�*�ޠ+7�Auf�v��t�����u��[���^�)�r�svp3Gn.ٸ��b�c��`bI� ��^n	g�b�onx������p��qW���@f�w�8�g�x�Kt��)H'����ݜ����!�=U�W݃M�\���Q�i�u�����7���߮�q��q"��Hyy���F�����7��1��n(T�I��=�(��]������gűEs���sn���S���|#F(crN�;����;~zy��;�m�9n6�۾ڮ޽6F�N9ȁG-ܗFP�T�*����^Vo� ��o���+����!%�Nd:(N�����k�y��(�G�D���� �}�w�z�*�%$ihlۘȻw��cD��Z�ssaJA eU7�}�}��Uˏ�ҕf.(�M�sts+�n~���J"�)��E)���|o@7׷��nc��TiƜ�q�C�퀑���˽��~XN��r$\��7}�Q�CI��P��`�Z���1�%Z�.`�̡���W�^�ރ���m�3#�F�3>Ϩt 9y�3������@܏SYZIm�9�I��  .䢑��x�PO�u����`��պ)ں��ty���Чm����B;�3ف|Xx�ڛt��j���DmT����ܛ��0)�.���6��m۪���� Ú�r��ج����wk�ɢ�vl��S�)��v��nvⵛ�ZV�K*��Unx���w{����'��^�m����ș��b�ʇ��/<�w�,v�v�^��N���T�TM.�/:�
o���&�-��QB��	T�U .�נ� �ۘ��Cyt:I��˔�hUJH�՜s�1�Cx�}Ku���s���8�N���`��߮��O^�i>�Ȝ�3�
�Ѿ��n�~#�u��}i��"%�^����=�;3t�c�J��sƪ��s�:j[;�����H�L�lk73����wN-EHъܒ�qx����T�#G �$c� ����iϲQ��֚m���*4��on�����;���;61���c%����`fnA}^<���ޫ�@�08�����,�4~;�T��^/��Z
��Il�[h2d��nNڲ�n��E ��/b��@�[��7����������m�\�7�|�@�8�ND�7�tD@� �����d3�z��\��+������n~�<$s��8o�@�A���Ǟr9�G2��IP����-�4��lŧ�~�(��ŝ�:�#F(crJ�~<�ܘпks=�z�\�߮��u±�*�6�
H�3ǶJ�f�b�Le#TfiA)R�HÈ���8�E���o�=x�	�ǡ)]:��w��x�ٞʣv������97}�_VCg�s{�
�ÊD�����tn/�{�{~��T(bD�Eaă*� �҉,"��G�]����,�8_q��fnN^c���d��Ύr������m"ASP&P0v:�-�7;7��Zxp��E2!pD䉐c�_��דs�������ϵ��#Q������g�(�����<o5���sIR4daG#�o���ܜ�����6il��#QH\0�7�#��.�o��3�'��A*���)O���>U�m��y3=�+�qw�n�k���)&�o����@"`5�! �1��Bu�"-��B*0�B��+��kL�	1`�UqX�"��H'�����6�z"D��0�H��1
	#
~0*�"�X$��СJ$��ΈMe/����$3ɯ��b`�	 ��,`7HA� �`1`�"H��"�1�0$���Ap�Q��z�ԀkM75��.���t����vn���ܐ  � �	I!�V��oPp� �              z��V�;l��u��s��(NU����@-�z��H6.m��XG��E�����)�S�/R��#9{Z�=]��r�ބM��_>m�����ې���V�GZU��PFZ�x�Bw*@�L ��6�����V��
5K��4�]V�
��m/@s15�I�a�z�J���2D����"�p�k]
�M����YT�OZ��x����:B��ا��m+�a;ec�:�Vއ��y.l�����G�Ù�^پ�1�c�~������q�@��M�-\�����!j"�]������<���m��#�nUr�S��$��kTN�<��s�cł6�q�m�q��6�)��H��.�n���"t�3vU� &�b^ŋf�v�+�	��OC�f mq���m�(%�*Թ,!]z�'n������*i ��bR��<�Uq=�����Ը�@�x�8g�;�.q��a��M����ص˅�k:)ֹȚ���.����չM��AL���9���F�8r�h-��\� ;����*�R۰֞�j���l\��0�P[�DP�=K�Ғ��m�������u��*�UUe	S�u�XG��򖇴��/M�q�"&�m�˳f�#f��V�K�i�i�:�F]K+�K��xv��:	݀'��[��kim�˫�8xf�v��n���N�%t���֨��ȼ��إh������Cm�(ʲ�In�s2��,��/8���C���Q��MDA�9���A�>��x �P?#��@S}|�\M�j��� �����<M=��
�P�ےI  &�z�r�ճm3�X�s�y�Vb�¨�ls��h�����t���VӴJJ�#��8ݺѱ�gn�n������)���g��X�wQ��9�'���KU��t�yx�c����"{�be�Z��v�Uj�WB��zW����s?l<��F�꥟ �k�J".�l�.�!���%�4L�]�
���n;h�ʍ��s�U��u�qW7=u��V}���ُ[��79Q�e���j��D��-�����7ڎs�C���%2
��Q�x�n�D@n�h]�A��:/O�O�r'$L�8
��{�>]��v�#�V�
ӌ�r4�`�i�f{ �c���d�3<������2PD�5\hP;��^59�;��Z��ػ_lRjx�����˼�������A��50Ӝ�Ep��Z��T D Po*��OO� �g^Kʙ()I)�&��=��/������L7k<Ɂ�!&'E��s�wr�s��;-����Ò����4�uܘЀ��n�9��vd�D.:�%�r��m�qئ�նm���� sC��=���6���$�P�w�4��p��gÝ ���<�?�.D䉔Tu�ϟ���m��s�.ݮ�bM��JR��D�@��O�~�y}�~� ���p_�'>ť�Q�Y<�e*��D�J�<� ���=Y=���-顏0�@�(FQP�&��� �|�܃���	{=�	Ƞ��]��F���'q(�dq0݋��O����R�L7 1��y��˼�;k�Ä�^�v�E!AB�T��Fgq�lü�r��8E�N��#��]9����9y�˿\��	_�o��BNE����|�M>y����A ��X�D�B%�>�A��*� �t��@��y��?�����R'$L���_�s7+���˿\~����n��L�.Ɵp�B�wM�t��x֤��rg�;+2B�$�m�6�
��<E�_=�3Q)�r���r<|/�}��zXJ��B~�A���J(#������BC7e���L��`nd i�Kq�܈���/5���`v�����-Ji��q.e�y�0=���/<��"s>p�����?i��q/,[@  ��p�3-1�F�V���Gn�9i�SBL�3�Y6]���"���K�<�#V�.Q.e�)�Kl�R�D���j4�d��u窿���p�&��І�&w[�/�Ү��5ϗ<X�v3�b�zq	t*r/4�%�jx�G)����V2\f�A�`�o׾�w�v���e��3m�v��'W��j�e�9����ܫL��POm`-<��(l��^�y�Aə��#^�%���,,߃l"�(�f�9�A>�D�k���~�	9��1#�?	���&QQ�$����>0.���Z`{=��#l���������s�y��T��`z0�D�چ�C��P#2|0>\�����?%���Ng�C�_>z5H
��vĸ�ݐ2 �'O=ǀ9�ݮƹ�r��r;Y�ss�s�(��$��A	&�ԏs�]"qφ� x���!-Pg��Y8 �����p�';�'��ٟ�m9���"NF�t|������BM��0�K��j��c�|�l��.2'F�4�.�X}��纘�7�%��L�&�`�M�yN{{$�^�I;Ս��A8d���)�Ζ�VD��$�^�pb-8[�HPr'\��J1�I��v�}�>�i�~�`�r� ��fbh�4��9v�F�b����ax�M�	��ە@eΏ��Zg��T�f��:���ʂTĴ�8i�(*/=I�grX�i�A���Ju�����P���Q-�0��>�`v��v�i��Įp�},Cr�zs��k\z�vs��7�nCv�Dst������5���\�nzo�`\w!���� g��M�,8�j�C��Y�	8/6� g�X�>0-EߔL�\�
\b�Vo�Pf�>������ϡ��<�2[�mđ�M5�ߥ��֘��?���~}F���M�����j�d�LL��i�qy�=J�3=,'���sL8AQ�h�	@�8�c�q�-���$��ѵ�&7T�������ƃ�~��0+1�w�a�e���/��2LKLd�NY@{��
 ��`_|��|2N�0
HT-AD4�f�|�f��s�n��$��$��w�q����4_�`^Cq�4�*�X�Y�DَqH!pQ'j��̂�9�p�4����H\INs�'�m�����#m� �y$ݳ��0���D�J	���1
�S�¢lH���A�;s�'N�-az�d��t���n�`�����c��6��M���l�y6�rsF�en-+"���MP�q�ƛn���B�D�v�a�-��ٮ+`S���۞���\��ݦ�h�r5,pJ�N�RE7 �N�����gH��fn(�gi��gkm7�\sO������K��_��|0;���m�n��s*�b3},�i�۟�5	=ۍ����Ro�D�zI�z`�i�v�,�3,mJ��q*����� ����gs�L
�Mk�!����$W�I=�k�d��I�?I��ps&$��F����jae7t/#��h��2m��nX������t�*Œ�����/Z`v��~ƘٽR�q�F�q��-�P��A� (�~`��(*|�V�P�������?z�$��"Oo\;�i5��oL���6�j�͟��T}��\{3論��!&�=��l8�A��5���BM�����Ĕ^?��a�RܹN"u��3|����e�*�|0/���~<o���X�s�l��X2c�Ɗ#���8��ޙś��`A�
�*��P�"	��Lt���"N�VBs&��"l�M���?G��KR���T��0/1���L����=��d"Z��%��d���$۴�w�y��y��I6��i�wﳝp|����4Е4&h._&���j�f�� `��X��\ ��^x@� ��|�0B3�HD�iU�R$S#"�>*�A���E�Jb@��@	Pw������ a@���"�)$=�鳈ȵ@ ���x>���}H��c����Ez��H�?�z�7T�����7x�r|0/r �@�Kq
T�߫�^���φ�ٽf2�dF�I�h���C�va'��Ҡ/<�������F">`�"%LL;n@SZᲙ�k���.�丮�E����������KX�~����U(��(I�mg�l8�A�ӊ�9�y#�2I�����ƨ${��cR0�5�ɦ�@��L��J�J!E��A��֙'���R ��-�$��I�0���A�/ʞ������	cjSp�[j� ɟ��0����L�i�Ե<�׮���ŎY���\�a��c�6�˱O=u 4�H�i��l��7Z`v��Z�G���`}�����)��6�_h���0;s�3v�D@��d�a�"�.e��z/=R0/'F}ߵ���0;�d�ˉj[d�@^O��0a�^z��n/�0;��s*\5
F�$�3�i��q$�6�2�����I?���=H��*�B��
J�@*�����;��_p[/om�  ��$D[�t��U�%�*`��K-�
�\��H��6�+;�lvPv��i�V� c=�k��n@=E��E�M�����v4����v	5��ծp\�|m��jӠtnHT��Y8]:�`�i�*��2�s;���t2sƷn�,�a�6\���T����A� �p �]�
�DKa)�e9�Jvw0O���k�[��M-=T������/[o�����K=�Ms��q�'"eP�Ӯr#�x�`o���:=ٓ')�%!U$�7$��Q&�#�8�E��02�i�|�CY2D�c��edA֙1����3'�`^O��"����ĩr���0/���:0<��J��b#�	��h"��5=��M������])��������7[�5i��/�eφnp~�3�����C���*�4�IGD�]aHz����$�ϔ�F��$�d��6␱jJ7Z`v/!�}��сVnSnF$���lQ8=,���4щZ�d��y#~��5�q8MW�;��^N���給l�C�K����,�tF�ݕ�y��xϫ�4�2\3�L*gWe��n6�rt`��4��Ό
�с��iN�-�N%���R���͔a����o�$�Q���㍋�9$���d��kٓ����ET��s����`U�L�ߤsI�9�l�2���90��Ƙ�с�j��Y*fX�/'F�4��Ό�}���?�{�K�2$a���I�1�QCθ�9���y�S�;����ͥ�Wni������}�����D��`wL�s-�m�S�Uy>v�/'F� ��q�r��p"����dؽ���̈�5�*�|0x���27*s,�/'���@^O���B�.q)�9�^�|Pg�l�L��%�^m*�Z`V[����;R�L~�}��Z������Ϸ:n�n,e\fk3ظ��ŗIN'n��:I�\�Ws���=?���c��I��k����N4�I���Dfφ浕y��D�_/xc�d�m�%��o���4�uR�/���;��.eH��&%�֘�i�۷�yD��P�[R��r�f���y��y>���$�Ѩ�  p(�`������#ٙu���̱�-���� ��).񕣥ۖ̀�ֳ�-��݉�]�Z�Xt��T�{��	�k9��6�o���۳���WN�Gm�<��2����%�5�9�l�+���KS9:��ۣm�v���k�g���V�:x�mj��Q���ڥ.d��kIX�e�'Va5Rt�d����� s�v�!)�AN@�2�M��J Ԓ�mɔ.�f�+m�~�������%Q����pIOU���h��|2b/1�U�֘�7Q,s#r��2��>��I|�M��`}�i�۷�[�mA�"Sd�C6P�4���#�o�y:030�S�ܶ��T\�o�&�=(��a�9Ó��D$�=���m�'n
$�d��'���/1��4�,��c�.ZĩgDݬ<GK,1��u=��i��l��K�I��w'=����T��Ke��?�nҠ>�k9P�<h���W��8�A��4I��'�~�K�s��.*�����(��?ˉDÛJ4�q�J1^H��W�I9�<w��o$�d�ݸ�Orp�LQ�9ģ7k�{>��a�IE�i0=f�X�F�Cn[Tr|0>��nҠ���~�M�}B�7�O�
"ZA!&o��'s�y��<bgk�MfK���_|�ˢ-b$l��4��cL6/2�gn`͟x{�Jq�䁸(�~���7�4֤w_�$���%��k����R4���6�âO.�G�I� X @�U6�'��I��N�'!ޢ�Y�ḃ7ZfDe������������qDHq��Nn��'�y�(�Yy�I�~0�x9ެl4�BxS��ȃ*�vezs=���q[�A	���J G@������q8�u�j���L��*�|0/1�v��Orp�lQ&�6�|�l��w�i������M�K�ܨm�j�͟�kj!.D^y�Q�z����Q2KCr��C(=�$�}�L�i����ݟ���(2�Ԅ���[��|��ВS�G$�D�f��I�qq^f�t�8��i��Nc��"�n�6���vs��<�懬cn��4�����v����q��dH�i8:I��P�M��	7�גI*���L����Y*[a�y>�"�i�y���U�%����r0�#L��$��w�K�ݡD���&�:��� �Q�9��@����$����'�](��˺�~��OBrp�-�'��
$�=�k�y��ӭ���l�����{��fİdIFHMB���>���1
D�AHA�D��4��z,�����`c ���$��%a� '�הB��ZE��@Y� ��T^�
�l=<�� hH�h�ĉ7�LX	�F�Y �8���B�htCV��� (�j�N��X#R#"0"�D"��	�Z��� T�8�E�LC&(	�����{}5����o�V�  m� H��[l[G-�pHp h               ͳ�l/ͭ�rM%���И3s�tͲ��/l�We�s����pV���ۚm	���0����n1#F)p-f�ô;��b�ѱ �u�c`)���[;r˴쬱L�+Aqg<m��J̑������[[��t��I����RM��t�p��{qTk���ume�����sǝ�3��9���ݴ�8�m���tݮ=vN�8h��X�v�⁥8�WK�J��9۷$@ո;�0���n1�Ea�X�n�㴻d���!\�M+*��u��b�Y���ȱZ�'�;4.k�ڑ�k8�Ȳu�� ڌ�A@Z�����P��,2��n,ɳ�#o� c"�Z�l�#���UQB�ٞ�
���6�'8�\�n�ָ��2skd��8ҥ՘x�&L�k&싷"����i*�Y+��Rl���ad5+�lm^'�9w-i�]m;�T�p���s��.����rmY�rj��և��a{9���hͱ�\
ed�5*���@�O`�:˯B�uTs���Y�q@ ��sm���镝j[`&v�[�0$M����m1n�����ZRZ�h x6�iL��R��J�UUYFyYS�=��84N�Y.J:�_<j�q�Y㜣�����s�Kj�u�d^s3�Hҍ˺�n���{����*�ʫ!2c��1vd�C�>��dXPˡu=�������b8�	�족\��Ԇk1l*����5;r�:�9��/EY��
�Q��d�B�����@�(�	���ZuM��@�u����������T6���4�S�"��� ���@��٭�����[�E�b�  �6���1[����BY�vٲL��%���4�,i̗|��}��UF����Og=���.{��n)q����c���;v���Omj�N.ȆM��ɗ�ֻb���fu-��=�]g8���bev\a[)G����:^|\�"hI�BJ��v�{�����'B6yD���<�7=�;Eϓ�.[rY��v��?��|��"X�Kp��m��~v�6"��P�O�v����Ʉ�"e���9����=�=�������V�DD>Cr�R����02�)P���m0/�{.drH�&�"Z�<{}�6|mB�i�E�:�;�tc�d��	�������L��*ٻJ�/���[]���O�3�޶G���iSF4dmi��C�3�ҝNFP �i�$� ����!'����h�\�y](���s�j���J�]�������@��ORE��*���9��9�.%��S�‟c��77)W�?k&&|��-A2�665�P����Ƙ�i����%�j\��(�_�7Z`v����S���@{|5��䉖�e��0'����
�zP�L�GU��g#Q���1�"�pL���`:�9xv�;�َ�) �q! ^)���߯���m��xP���*��}�Tn=�\�r@�71�@���@^N��i��֘V`��M��[(�сy�yT~F	���4uPR����$��g�rN{��ٗ)��T�1%��0;x��oJ�t`U��2e�r�LD9T���^ei�3g�6#7Z`b�Bdk�6��7�x��Ggq�[..�3�tZ�s�ے�̸��%𖠙T�?��ñy-~�.�f����D�K�Pۙey?�$svI���۹�_s����$�p9�9>������-\S9��(��én�+Bp�r@�O���3u��/'�伔~�\TI���s������e�LM/�g� �i�i8(�n��y:0/1�z=9���$�_o9�>�H��!���h��L�ar�U�Ǯ����p�]m��B��N$�7!�N��ainnТOs�!'�sƵ#`�yyHĊ�
J���/1�� TM��I���D��񄚳c&���J1D��i� �ǥ��K�9���֘���&L6(r��T�?����Ƙ|��M/=9��4�7�>����4����B��(\�9��ǿxH�䑱2Km�  X��+N�5׮��OV�Ug�L�
�u�zpsY��8����)�w2�v�i��΃u�l���¡zlh���$r:�k��wTMmĻ�,S,����ޤy����U���\t�.ઃ�tU.ֹ�r�ɞ-�[��[�6�v�.̏5��sq����� ��͖�n3Y��2��[�Eh�'U��)t�ŧ�=�%;4��Db�.c��ߌ��0;x��o��_$�������0=}�2�Kr�S-P�4���\�9v��&�aD�]��EQs��dT��'wޟ�G5�Ã�n��=�A	4���S,6�l�}� 8��,n��@^|�""��Ւ�-��5<��$�3u�˜�J�iP��T�o�$�maU���2�&ʁv��SŲ�Ӽ�V֙'��?����	L�o�����\�����%ľ\���|03�eJM$��BMP�s6��׀P�q J��O����A���P�%�0z4ŪX�Kp��2��|075�@^y�n�O�^��1��8�x�/5�nߊȈ����̜#K-�mKey�0/ˉdei�3g�sf�D�0�$@���!�m'�g�=n<���mciĦՠ���)��6吥�1����~(�сy8yqT�}�#���F8hPI!T��s6�
� �QyXQ�D;�T��ɭWy�9π��l|$bH�9�(�~o6���s�!}�gP�����h���0�Vlc��R8�I(h��3}\aQy��v �����;�����u��p�)6=�Nnύ{������o����֘��D<L�Hcj8�<���<>+��4�@��]��i���g�z�(Pۙey>����yTDE�?I>�?2�
1�sv	�  +j<�I���D���>H�KCQ⍴�7ό6/2����ၛ�0/��Kqa-Po8�7k��>7vO{�2O�hr	����B_��b" ��ɗ"Ų�T�I	��c~��ޮ����~(��|v�B� �,  MQE�K�t�㭈�v�4�t%)h1v���s�F��������9��۽��s�vcW��GpŽq8��Q�D��A	5w�(��<��*�	���g~zϙ��.N"�����Ԩ��0.�ߚg�3ҷA��JR%%I�"����6���b�s�Fn���/}>	R��p��qA�ۤ' v ���:�o�$�}�I���p�@��y���R$`Cl  m��x��r�V�3qQ.&M��2�n�į�ȥk6W�NT�Y���!LJ��q6����.���A��k�3N®Qܥ�p!�pM��y���0Fkh�rm�mȖ"Ԝ��s*պ��;����5'nQ�G68�f�Ge't@�knu�_�P���e-�	2IsWZ��g{9�86��Jtx����WB�6����o9k��^KL��*#=�8�U��J	ߵ��q#IAD���
$�͆�4��֟���A�嚘ܰ��3-t��0���L�ķ~�@^gԨ��9��Ԩp�1@f�L�6�y��A�������0;�-�.q��q�$�zI��P��Ś��\�+�{I	T��ㄸ�d3q�jb��:�N�^�+bi��n�������??��9le�����i�w�0�g��$h�7uo��8��p8 B�PR!C�EB���""*��D���F�yv�ׂd�|��I�À8���T�'���H#��CC� %y����C1cX�
I�|r����x�Dlo��ˋ�%>�u03'~aB�G�HK��&�'ƍ�����<��i�w��.b1�×-
H�/[<��ч3-Y?�~���!�8��$����w/=}�M�rڙl��Csv���YP��k���d��7p�E�D���M�G3`�D�d��Q:��{��L)"lT̪$����qY���!�٥�^�δ�I���ט~I��   @ :�?O:oEWL$ڜN'�H����U�m��B$%ed���p�{ �k'��s�ct��g�q4B0�bF��TuWHv�mSd��7��w���@�g�p����ݓ�{��Wgg���=�m�~�i]���o�!���s���c۷&qذÇmێݻw���
B� B��SF���������K��+���qvQ�#��#�1 B �����a���@���� 9K�N�$��I�j���E$$�}>�@S�߇D���O.�D�����g��	20���D�[�}��s�}[��J����ʘ׶'ognٝ:^슆��ܻn�����l�ݷQ��$�]*T�R�i�z"7ޥ@f�Lݿ�u�<���Hzt%8�a�Gw=��G7g�|��|���%pq#v�}f`i�a�7_�"�w38�`^��Hh�(��9CD���<�I�{�I<��2O�x ��/�x�G-T��Pr��Jd�T8���0/1�nޔE�0?q]��S���Q���qp�sc=s�֫G:i�hӥ;6(�������P�㉠���}��۹��8��	7�$��oQ8�e�)�Z'7_�]�8��#c=�i�~Ƙ�Y�j\�nT6�Z(��`^cL�\��Eg��%+̯$��0�"D��*����01n���~(q�\K����K�(1R��Х
��&�=���̭:�z�`~^[�%��E�9�[�X�� ��uPꅶ_i[FH]^S�F��.�`t-��L�2&ɸ�p�8;K�`�Z�$�npʰm�òqv�gd�)�kp��l�3\l,'^��4ړ${s�k��ηCۛ�+�.��㥧]�@H�:��8��2�z��l�zr-�%�]�s5�c����ְ>m]���O�v�[g�rE��qp�x�����%�7k�kw{���_|�ɇCl�k�{��Ƚ��4���!&�D�)r$�S�m�Ԓ��"O.�N�  FD@ 
��C�-�Y*b���4��Ƙl^e|h��<�?�8�������Q�'Áqr=�Ԙ���2/�ڀ�֘ٹ�j'!�Q1D�̚}�J����3u��{u3��oS�b�`J��;e�˹w��6����V[rY���ۚFy�\�ԧ-ĳ�l_��y�0/���J��3v�(%�����R�7�n(�i�[�B0`@S�� D@�<���<v��&��P�-݁hnq�Ӝ�
'��!'�oQ�%�(���0+�{J���l�q,�J68�A����63���Ƙj�9���\����:$NI�Hh����P�ޥ@o�i���}�]�6#Q0O�sng���#�i,�v��\��guǐ�[OHp��1��G�}$���ۿ�o88:�Z��{��L(�M����N#�۳)P���cO�I(�=9:�Y�p��I��P��o���`iS�A	9��	7��$�&F��+�}ȉt�u�&�Ao�H�<��N�=�X!,q6��֘����+�ug�$�8�K�@ӂF�&&�XIo�'c���5< �{�������F�ޛ� {�`v�((�����.��(d�iCl�j������̓��f����l�88�|��GR�4Cc>��4��%3�kL�~��/$=��ʗ0C�9�/Z`^cL
�znOG�g�`�v'�j��l�\0>��~^�#��9�`{<�y�����N�򄛼�u#�8��%���x1Hm�#���ˋ�L�Ok<k<tg� �Ȗ(��8��/u��2/a��Y�K�9\�'~���7��20���GR�ϡ���0/���ߊ�Ͼ\l�ҾP|m&�P�ﾂn�d���|h���(M�W0�ۜ�4��Q1g��$��0�2/a����ަ�}TH�%�D����q��i��֘���������u�H�l��M(�rI$� �����6E]ɯK:ۧF�nh���8ajV��1"pX%�LpI�i�r�ڑ��[���[n������^<�rn�M�m�A��y��gp���ێ+lJ�͆z�M��tZI�h%�ɢ,��9��ˍ�nMؤ��B�@�]j�Uh2Ϭ�ğ~�}�ߎ����n���W��`��/ltr�]��9��y5�m|����GL$�6I����M�4� ��R0��ex�1l��ܩs8�3u�o`v��@\f���#�9��l��4�b�9������49ıo�sv~K3鰩���(��/�����@l{�`^cL�ό�Vb!��̐ۙeq�x��}֘�zP���Ƙ�S�"��%�c���9:y���Sٺ��=��-���/g��8��7���Z`Wm��.3�����6�#m9��M��=_� ����ͻ~(Ǿ�o`w��(��Kh�To��#}��Ȍ�4����I�>�	��I�Z����� �{�eDB��*�����۔G�!*�	RUN��o4'� F�@�y;$����Աo�~�{W��""[	��K'm�c���ŧ8�r=X��(�]29u+�#�33+�#7�`U��'~�3Z����ӆ9M�J��7y<kÃ��G�BNf�	'��
Ks��TF(�R2e�#}�i����W9�I(�Z�����ވ��/�D^{�����o�٥�u�L�S�8m���0�K$����qo�$��қs����pQ&�D���  oxxI���s%��g8�
� IB�e�$�4=�<���� ���jɃ7ia�[.H�NTNBS$�3Ԩ��`fc^�K�Tg����+�h�8�Q��p�'V�LH��!��I��4�����|ɒ2�M�cR���Az��h�� L����%��D��xj6�jBEF(�����Iy������$��|�0  >������}잍8c���(�(؍�������0=��TG߾�G=h+n�ƻwe������	JCՂM�O=�B@TF(�QF��'V�BNfA	7~��s��������L�S�8m�z �{Ԩ�i�woȠ23���Qf�iM���-�)I;��n�a��oV�Bqw\�wsт�H(���4O�-�t���ru���B����M�aq	�58qg�OsD���$������w�fu�M����5�B2IIY-)+)-+$#XH���Ie$( A�%l�I��ž�A
+Ā$6�q&��V �#@�,`B0�-�0O��e��D�#���� �n@8@qbE!����C`��E�t����`	u!�6�z�kp>wi���_�2&��h   �k�$m� �ŽN	 m               ��taiU��l2�^G�Kk�Q��8���^�[:�,ᖎE��T+n|�l�1p5U�I��Vm.�b2Bqvz���v�Ÿ.�e����v�����U*ܛ���*U���掉�YY8Cj����Z5#cd��q)�蛒��֍�h���9˱�5XԙzZ�ۮDԌZ�W��oR9w�[�N�+<v�gv��s Z�Pu��"�+��H�
�7��6�Z��7M�7���۴�ĶY]�AN �m�6���J�ƴ����gj�t��g\@&tW)�{qr�qG��t�-��I�DȂ����){q�0u��jс�lq��f]�:3��A�su�u�{�u�y� C���I��\���ٲ�O�j�P`6ӯL��n�ѱ,�A͉��Ǎւ����m���۬Z����p5��^�I=���`ul�OIr��N�N�2f4r�P8�;�n�g�3˷V�Ma˭p��bI�����lt����v��)�-e�/e��wfU�V�
x�#��A�ng�6�J�U@��T�:-�rp�oF�U�b�퀗X�[-��i:V��RL�=��[�m�R�UyV�Mch:`)Ik�d V���)O+*u���LSZ��Y�78BмHca��v\u�Ļ��S�+fIye�2S8�,�����-��9E�3��Ψ�uv�y_�e�OCۉ�%콴y[<�a��=�U"�)K[-�`a���P�tصm���)n1�:�2M[L���f�f�������(>)q^�J��9D��Q*�ڕ�1(����_u��sS��fcm��M��  ���4��Jܗ�}��>�b^�M��Y5�Yë�ם#�QNs�mb:����n�F!ݐ�݃��ރ�z���:�mĀ�ap[o�[G�+�,[�9҃X{�U1mR�C��NHEbR��l����<v���ٺ�~#���}Ã6�=�ӵeظ�W_�����}���vck�/d밽��568��-�Bt�aas����`��v�6䑑G1�3<�]�L�ޟĸ�8�|�򔑼;�Q�nq��b�7~j{o
"��4�ˉL��f�jSp�4I��׏I6��K��03<��`�D89R��P}��J$�97t�': %w���'3$J%>C���P�i�w�7w��՚�'��E��L$���\p1�&�q�Nݜ6��ݞ�ŬMqZ3�?۽��
�������?_4��s*#>��������(N$�APQ&��B�>�N����?� ��`����h�G�_��5#mKC������A�֘��T߶��ƏH6�˘�#��;���a�v���ů|�&�����4�P�t�4���Į�z�LF��
�i������!	�#���iN6h),�������+t�@��RJ���&�I��Nf��qf�I�d)�-�P�һ�1Fp�����`w1�_�`w����2y�*���T�	)�%�T�7oA��!���"� U4�D�4�����߇�$�f(I˼��np���pQ;�·d�� ^����ܜ������A�[j��ϩP����?%�bs߶bn%�bX���{�߲sX��[�<��vD)��%%�4�l��"j�e��ޤ��.�.f��0�yı,K�ߵ��*j%�bk�ى��%�bs��0?ND�K������Kı=��%�L�5���eֶ��bX��}�q,K��ى��%�by�p�r%�b#���s��<�#�����H�p��[�6��bX�'��f�X�%����ӑ,*�MD���X��bY��{�'x�G��>��i@�q�\6��bX�'����"X�%�}��bn%�bX>w�17İ?��􋁞w��޴���`Q�&<R|�H�˓W���r%�bX�߾�&�ؖ%��{��T�K��>ى��%�b_<���r%�`؟�>5~�5��>ٝ{=�'��Ѹܛno�m�n6��gf4�ul�1�[���m9ı,O~�f&�X�%�N{�I�Ȗ%�H��}�6��bX�%�﵉��%�bw�vv�Z�fj�]a��Kı<��17GQ5ľy�siȖ%�b_~�X��bX��{�q?
��j%�����l��K�2d�Fӑ,KĽ�߳iȖ�b_~�X��c�@��j'�}�q,K��bn%�bX�����f]f\�a�\��r%�bX���kq,K��{�q,K��l��K��5^��ٴ�Kı=G�n_��0ֲj�Iu��"X�%���l��Kİ���p��Kı/���m9ı,K�﵉��%�b�a�oϷ��B헯��X�� �Z�����J˵����V�j����`&hw[ ��2a���{@��$�=r�W�鱹��v�K�Ayu�wPmS�#�d�q�����Ck�{l�v�� ۰)�͒����o����fK#�Ss��hyZ�k��Q�I�Ev3ɇXr�u��`�١z�,�����w���n�%�~�ob͜ƶK�g�=�6I��m�*���n�3b�X�-�(O~����7���x�}ݘ��bX�%��{�ND�,K,	�����Kı<�vbn%�bX���MFT7
��:x�G����ND�,K�﵉��%�by����Kı=�혛��5SQ,N��:|\3E3S���r%�bX��ߵ���%�by����K冢j'}��q,Kľ��ٴ�Kı?}�֦�C5u����ӑ,K���bn%�bX��ݘ��`ؖ%��~ͧ"X�%�{����Kĺ��}��55��j�d�O"X�%��~ى��%�b_<����Kı/����r%�bX����Mı,K��ِ߯˚�Z����C�vU6�qŻS^{=��[�GXX�a�55���8�D�,K��~ͧ"X�%�{����Kı<�v`�c�j:��~ቸ��bsG��2�2�k5.�6��bX�%�﵉�C폃��K�؞ı3��17ı,N{��Mı,K�翳iȖ%�b{�����Zɫ�]kiȖ%���_�ى��%�b{�vbn%�bX��=�6��bX�%��kq,K�����W&��)�[�6��bX�'��f&�X�%���nӑ,Kľ��dMı,K<�����<�w2�[��ʋ+.ND�,K��M�"X�%�����7ı,N{��Mı,K�>ى��%�bp����k%�$��57�q��/n��k^|�h9]�HJ�ʝ;�Y�ԛ�4�f���r%�bX��}�Mı,K���q,K��϶bn%�bX�̭5����<�{�<�N#JI�<�bX�'���M�Q�,K�;�q,K���wٴ�ı/~�x?8�g��W�l�8cM��ND�,K��ۉ��%�bw�wٴ�5'��N"4^4�� �|7Q.?kq,K���혛�bX�'�緥��#3Xh��"X�
�b}��siȖ%�b^���7ı,N{��Mı,w5���q,K������]f\�fK��r%�bX�߾�&�X�%��}ى��%�bs߶bn%�bX�{�w�%�bS�/N���!�O�%2���� ��d�Q�q�l,�ҵ:�ynǻ��u�|O�&�K�~��Kı=�혛�bX�'=��Mı,K����ND�,K�����Kı;�����3Z˪kV捏"X�%��~ۉ�A (	"w�{��$�N���HE$M��"A�j%��{��Z�K��&V\ɴ�Kı?}��siȖ%�`߽�X��bX�'���Mı,K�>ى��%�b{�Y���j�f�uu�ND�,�E�M}���7ı,O;۳q,K����17İ?�S��g���>��&ӑ,K��������!��33Z�r%�bX�w�17ı,O|��ı,K�}�fӑ,KĽ��bn%�b"9���K�Ӑ4���	�514�D�a��CgqӸ�Wv!`"ߎ�{���.��)Y�����,K����bn%�bX����ݧ"X�%�{��b~����'�T��p��Kı>�>�4K�!3Y�\6��bX�'��M�"X�%�{����Kı9��ı,K�>ى�⃊.ʼ<��[�����\]8��,K���bn�bX��ݘ��c�5Q;��bn%�bX�y��nӑ,��{��I����M\2�[ND�,KϾى��%�b{�vbn%�}������v��bR*-�{����KB<�9�SP�A��b�:x�E,N���Mı,K�3��ND�,K�﵉��%�bs�ى��%�O���9���-�I"A��1%$�H �7c�h�]#�����VU��}�'j�4�*{9\�G5c6��sa0�X��[UN��B��d���V/V�X�c�;go<1����۞���7�wc,��q����l�@Ek����o9�
�b�PԺ�v�zv����5s <�k�,����+�rwq��>��4����yn6��l���<\���=u:���9���5��n�]��7���x�?}�Ϯӑ,KĽ��bn%�bX��v` n%�ySQ=��17ı,O~�=:\�Y�ɒ�]�"X��{����Kı9����Kı=�혛�bX�'�g�nӑ?�)���b~�����չ���ӑ,K���혛�bX�'�wf&�X����D�����r%�bX��ߵ���%�`��w�th�35���ND�,K��ى��%�by�w�iȖ%�b^���7ı,Nw�17ı,O_r��0���f�p�r%�bX���}v��bX�?����X��`ؖ'�}�q,K����17ħ��a�_�H�A@� ���G�u���]�>h)������l�M٣�w�{��"X��}�Mı,K���Mı,K�>ى��%�by�}۴�K�G��H��Jb7PDܮ�x�G��}�p���"g�{����bn%����&ӑ,K������r%�`ؗ�~�&�@�MD�}�w�^j�ֲ�5�sFӑ,K����bn%�bX�y���r%�bX����plK��{�q,K���k2]jY�	p�r%�`�'���]�"X�%�{����Kı9����K���MD￸bn%�bX���t���Z$̙��]�"X�j�k���&�X�%���f&�X�%��l��Kı<�>��r%�bX���߾pɚ̖�:ʑm.�̇K#wg9{^l7cW=���1����}�ܔB噙��ӑ,K���bn%�bX��ݘ��bX�'�gݻND�,K�﵉��%�bw��lѣX�֮Xm9ı,N���M�,K����s[ND�,K�﵉��%�by�vbn
�bX>k�O���d&k4K�ӑ,K������5Q,K��(0$z�=x;�i�m�l�w"X,�Ȭ��dg�D&�\a�$ Q�%��.��I�@�,����,�
�aᢺkkK
=1�R�a�#I hbXBD���M�K�� ���zA�HB@]�Ԃ��!�`[֎h:6� �����c
���v�p-/6�=��BS��P��_|Q1^���U~��|G�,S�T}dG�L�L�o��dL��>ى��%�b~�ݘ�x�G��xtGR7ȫ���ı,K��kq,K��{�q,K��϶bn%�`����nӑ+\�3��F���#p�M�O�D�<�혛�bX�'�wf�X�%��o�iȖ%�b^�~���bX�'�_��Y���kL�����2K&ǆ[�n'k\=��`ZJ�]'~�>x��r+k��~w�ı,O��f&�X�%��;�ͧ"X�%�{��`~R#Ț�bX�}��Mı,K�����jf��	�6��bX�'����c�6%�b^���7ı,Nw�17İlO|�f&�6%����gg�K3,����sY6��bX�%��kq,K��{�q,K��϶bn%�bX�y��6��bX�'��o髫��fff���K�©Q=���&�]��MD�l��Kı=���6��bX������k�)@с&�`yk̓B�(*jP�Nӑ,K��l��Kı<���r%�bX��}�Mı,K���Mı,K�����-�n��jR�˻
�\�ݽVDǮ�Հ�q\�l�N��b�v��]���ꦢj'�g~�ND�,K�﵉��%�bs���DȖ%��>ىG�x����8Z�����\<%�b^���7ı,Nwݘ��bX�'�}�X����%����nӑ,K��߾$�3Z�[�%�m9ı,O>��Mı,K�;�q.T�MD����iȖ%�b^��bn%�bX9��w�(\���)�+���x��~ى��%�b{���iȖ%�b^���7İ2j|��&�X�%��L��Ɍ2� �+���x��M��`ؖ�H����br%�bX�{ݘ��bX��bn%�bX�î�>�<Q0@AC	:���Ow�6��,�m�  -�Cnx�j%�X�.��6,�l�;պ�4suòƷ6p�݆ܛ
��;9�v�CH��li;N�5A�]�;��p<��u���=�u�N�З�1��P��e��aZ���夂��`�ER��ێ�� ���=��t�z�.�hX�d��Q����ou�w}�}���֊ۓp�ݗ��;�Ʈ4����.y��z.�V�e��e�]��,KĿ������%�bw�vbn%�bX���f&�X�%����[ND�,K��7����%�!���m9ı,O�ݘ��bX6'=��Mı,K�}�u��Kı/�}�Mı,�g��F�c2�榰�r%�bX�w혛�bX�'��{��"X�b_~�X��bX�'s(N
<�#������.d�)9ı,N�ﾚ�r%�bX�߾�&�X�%��=�17ı,O|�f"�<�#�l���-D���#���,K�﵉��%�b�}ى��%�b{��17ı,Ou�{��"X�%�罟Ms!�	��a]hզ�� ڭa�+��:y0��uh@xغY���w�{��%��{�q,K������Kı=����"j{Q5�}ˉ���#���n�^
$l4ӐWqp3��H��혛���(�
^(A�P�'"n��}����Kı?k��Mı,K���q,K��ٞ���&hԺ���iȖ%�bw_}��ӑ,K��_}q7��{S"}�m��Kı=���Mı,K��9��#H#B)#��x�|���n%�bX��ݘ��bX�'�}�q,K騝��u��Kı=>�M�5us	fI�3Wi�6%�b}����KĹA<�ND�,K�}�u��Kı>��\M��U5��G���ۭ�'eI��ov4d�읻dl��<3ƚ����`���f��e��Ma��Kı=�혛�bX�'��{��"X�%�����~r&�X�'���Mı,K����Y����c5�ӑ,K����m9�$uQ,O����n%�bX�}ݘ��bX�'�~�fӑ>���<	���p�p@܎�:x�E,Ou����Kı;�vbn%����CH����Ț�����r%�bX��;�����:�bX�{ߤ/ֳV�&e�r%�e H�}ݘ��bX�<��Mı,K�{�u��K�#��S��<�#���zх�;��iȖ%�b_=�X��bX�/����ӑ,K��]��n%�bX��17ı,O�y��y�B�4f�.|X=;�B����-�'���p�FY�ٮ:�f\Y�z�5��%�bX�k�ߵ��Kı>�~���bX�'{��Mı,K�Ϝ���<�y��%8��ӑ�"X�%������p=�A���{�ͧ"X�%�|��bn%�`؝�}�bX�'�}7����%�&\�]�"X�%���ك��%�b^y�bn%�bX��߻��"X�%������Kİ{���kRkf�r�a��K�¨��M{����Kı;���m9ĬK�����K��	��Z��,$TغDx�DM�D���bn%�bX�k���e�m��&a��Kı;������bX�?_{����`ؖ'�}�q,K���	�G�x\0��H�N9&�ny�x��S����O�V�5t�1^��А�`ڵ�s���.��^'bX�%���q7ı,N��17ı,O<��q,K���⫃����g���B�Ɣ��ND�,K�{�~T�MD�5�vbn%�bX�����ND�,K��#8(�3��<x��%
�6i�m9ı,O}�f&�X�%���iȖ?�@B:��������K���������g��0��JS�Ma��Kı;�w�m9ı,O���q,K��ى��%�����}�8(�#��<|t�N2�Q��y6��bX�'�}ߵ��2:���'��f&�X�%�����Kı=���6��bX�'�;���9���&oY����r6�  m�}�x���/6�0ۻ%�)r��2#��ݷd{:Xqvp�ֶM�a�N�+�����KҜ�\
��Ԏcs�/&��x�C�͚rV�3&�¯�u��8�S��s�ʢ��B�6��H�Fsx`���t髻]z�jZej�X0;\��igX����m��ﾽ�%v�v���."�H���d�o&۳wN8�e{n���K؞l�]���'�,K����혛�bX�'�wf&�X�%����M� ؖ%�����n%�bX��=�4\	���Xm9ı,O}�f&����o*j'}���ND�,K��v�n%�bX���17ı,O|�o�]a�ܺ�3FӐlK��߮ӑ,KĿ}��7ı>�O��Mı,K�}ܘ��bX�'z{�U�u�Mk.ӑ,KĿ}��7ı,N�ݘ��bX�'�}�q,KL�O|߿]�"X�%��#|�V#q����x<�{=�q,K������Kı=�=��9ı,K�����ı=|��뢺��M�m��ϰ��V-�Ft�Uε��b�GrF�m8�pt�#��<��ț�bX�'�g��ND�,K�ߵ���%�uS���'"X�%��=��Z�&�̌�ND�,K��~�NB!��Tgֻ���'����\������l��Kı9�혛�bX�'�{;�]f�e�eԺ˴�Kı>���n%�bX���17ı,O<�f&�X�%�����Kı>��M]\�\�.��ND�,K���q,K������Kı=���6��bX��߾��MD�,O�Ͼ�F��˫���iȖ%�b}����Kű=���m3�5ı;����Kı;�vbn%�bX�k�m��d2�F�y�˞�ai�8-]��g���E��tuٞ�k�2ۚ���6��bX�'}���ӑ,K���oq,JD�;�v`m6x2��!���<$a�p�S��A$O��&D�%�bs�vbn%�bX�y��Mı,K���6��ؖ%����څ���j���ӑ,K��{�q,K������K� �*V� D��X��`�+������O����"X�%�{�bn%�bX�w���W&�.h���h�r%�bX����Mı,K��y�iȖ%�g��~��ND�,WQ>����bX�'{3�_��rj\��a��Kı?}߸m9ı,Kߧ���Kı=���bn%�`Y"y��17ı,O>��3Z�e�0�g�7'N�8��g<mڸU��C1���z�f��,݇5.k.���iȖ%�b_��X��bX�'}��Mı,K�>ـ&�X�%�����Kı>��M]\��s35��"X�%�O��NC�7��,O�ݘ��bX�'{��M�"X�%�{��bn%�bX��=�4\	p̚�iȖ%�bw߶bn%�bX����6��bX�%��kq,K��ى��%�by����2ۚ��6��bX ؝=���ND�,K��u���%�bw����K���y!�@S|��Ϲ&&�ؖ%��_���[5�K�6��bX�%���bn%�MD�N�ݘ��bX�NyBpQ�G����V��KKA^�����Z;�axf�׋v�W3���6:u奻����rR��1	���d{��`e�L�.}��[$��8I����n"�4q��~�i�wo
 �d�31��6N̐�"%�*��ǥ nd���Q��ٍ0=f"%��.&bY@̖f4�۶�v��71=&&Bd�m����.�g���P�e��K~�i�m��l�(�& f����W��|����o�b�TN�+�H��@JYB!�{De@сM��i5⁳t�D�@dB0��H�HBc�/����j���@�%$�� !����;�kwZ��%( �tuPO0m�~�D��m��`  HmrD��$ ���  �               '5��Lhkd�{5��.%���;0V$�$�i[Vݝ�r&�͵�=g�7r ��U-���4�ړG96Ɔ�'m���;���\�6��UN
�V�\��{]��J*�UÞ�&4��k]�m�\S;,ʇ�Ju�����J���_g�R��yquR�v��Wc�N�^j�Ԏ^
�p�m�cݒv�ױ���vWg�����qH����P��nM��;(mO9^]�i�rN$��CtW�ts�v�}d���+��UT���n����q�6��1�p3�5�ft8�U��V�[�����
�EC�V��1U���ey*�х�x��3�<<ٳ�*�SR傶�=���� WD�
��l M�U�ڳU�ʒ�)�;�	�����S�g��m�÷Qi��F�^���8u}��;FTV��<�ZzMn�sg۳V�r�ݵrj0�Fv�c���X봶x8uZ��q6x�l:n���!Eݗ��*v���׫�\�o-�n�������m�R�y'm�ut�϶e��UX)V�fl�;��ڹ`T6�q ��yZ���U�3�]���K*E���6��I�u�N�8�l��=Z�r����AX��7+�=�mI����C�j=DL��6��L�S&Ērrs��v\o��Uf�I����n���j۠���V���ރj1%פ�O%�I�<nx��Y���.�- 6��c!0���κ3a9��5���&�3!5��a�����*�D�%6�
� #�O�#�(@�:���Z �OA� ˵ ���h�!a��ˬ̴�L�  :����j,�;�K\��x'���7W`ݢ��o��������6�}��a���s�[�Ml7n6�8%V��z@�mo9��h���6ͤ�1���vb��y:�u]����5�=�Cl��<�w,��ծEC�y�W7Y(�#o�;��A��F����ؐ��;��M���U~p_889�T�.�A#��� ��.�v�P�UK�B�yAu�z��2�����Mx'A-~7Z`]�?fK3`_e\h5ӈs ڠ31�N 72X�jv�	�ϸ6��D�4"N@���'���31�{�s��3��L�~(�%�1p����{�BN�Fa&��O�\$�/7�8đFi�:I��L���Ӡn��T���l26Ɲ�Nq��㮶�x����nz3���=�]���s:81"���i�D��NfO'�k�	9�$�^�IZ���e�qƜ=$���^�͍��"!�� [����/�҉<�N��������ԤU2�*�s1B�83����e��̧*a��#�Z�;s�����tD8��*�G�NbK!�f=(se���0+���q+��b'�DC8J���×�+�nn�<7	�قn��h����th�tX��������$|�{������2Ɇ���١�Ĺ	�u\�����/�,�9���r�6�Ģ&�M�|0*��G��O9�P��X��0;d�C��1/�,�;��(�e�w80*�F���r@�ˉ��P���\���x��c�ߊ:y5�ƛ�lb�eD�,N�����Rnƣn�v�+��%�M�Ӛ���vp`_g]�(7e��̡Ĩ��!��rPs��_L���P��X�&�$��!-�n@�j������`]�!�w>Qո��Cm,��s��������̝����P��`(l� � �R�آO�{j ��Z���$����W�J��Df��ELM�m182���m��lf+t�ӧ:Goq-�&�쎢߻o^��Ei���&��Τ{yT(�s�����ۘ�nfdľI���J�q%�K�taQq>��1.E��j�3w]w:3������ݥ@{4z#hL�n\�w:0��@wo)Pn��������R�@eΌ
��T������@~BĀ$"�HvI��l�5��ZkSuֶ�  9�mN�a�v1��[v"�9��b砮ZD\m�u���;��o�m�`��zz<K���Y�V�@݌�v�v�N��ly3c����;�'�8�]��'j�p�L�vI�͠�;h����fF����8]��r�\�C[!V:�8h�P�)��jfL�k;�T�'[�Ham�]�Lb{p;�؞���u`�8�c��t\ܯi�Oh��-7-�2��{�� f�+���4M����,��B%$�(�wޖvp`_g����s��6�H�K���сW80+o)P����-�.)���;����J�/vX{�/�7�ၛ1���!�ľ�������#=�;���|0��?��k[�nƜy݇��v��ڸ8�Y�+ ݵc\�-�)�B1�ْ
$��p�V��*�Fwr�v ���&G(L�n\�ܝ�]\I.%�H�#'Fo�J�7�s��8����mN���h�z�`��T�6s���N��i��m��Pl^NҬ�65��c!�]���p���j�@lf��ǥ�I��(Q'0璨DQ�DD�I-�k�l�Y�%�Ӹ��2Ӭ!�:Y:^��ۮH	q@w'Fvph
��/%�F��Ҝ���p�&\2��ϐ���R�63a0*�����8����P��f䝾���z~�<'������:��\0�%��$�-Ũ��k�HcmP��`U�
�����R�7t�&&�2a�s�_��:0+��I��
H:�	
"Z ��L#]�ه�v���n&0/�8�zg��Ѕ�	�3(�����T��l}Ps�� ��g�ۂD���o>�
$��P�V�;�с�[��8�ڇ-P�����P�����iP��������D8�;���80+�����R\�:��aJ�B��&�˒���]j�4ÁB����	=�e*ћ
�p`~K�#�؈Q�i��3�{:�x���su��K^Ѧ�f�ٮ+M���(�z���
���]�q�.f8��j��͆\���Ό
�����10�r9nb��N�
�����R�63a�yk(q1(r52��:0+�����\�w&�I���m�!NF҇���m
&���0*�vt`R���Q����DwٯO�6�G;I6�  *��Y��	8�_	U\v7�ɭW/\�t[�6�MC盧�Y�]!��#U;wd�-���u4&������3��
nz��st��\���J�6b�67%�QYckgp��E����������dm�F�~�N����޻ϕ��e��5K�h��[sY�a�>��@NK���4�"E���@�3�&�g7~�}�X��!"�jm+F�/]�*M��ﬓ�_�HU�
��`Ww)P�ݡʕ
%���A�3�k�-*��CD��z��9��SP�@�4I�l�]̡GR��P��za&�`Q��i�D�4C��@lf��pa�8�}����܍��s1����@z/!�W807����B�4=���x5�AQH&D
$����'cy7n��AV�����xJ���I�d�O�ڳ�0u�z�`dv�}Vɉ��W50ֵ�rN����_F
2 �H�v�q@���϶nI��ےM��L�#�3�Q�N7#b�7��
$��`U��4�ꎫ�ᄎ"[C����`U��~�߷���#ޥa6�q{�K����	=��N-y�H�[��`�O
=���VS�f�D]W�Vn5�b���G<,[��~�`Ws)P����s�\ÆL��!�@v�jJb���E��0*2� &\�plcmP��s�<�������I�m�l�  � �`v)<��{� �� ��h��h�Bf͛%�L R(���Fj�E���Cq@�BI��R$� �`E������̊P�$G^��d�4`�0�%���d�kA�3��{�4�h�y,��$J'���a�
$F�X���Z�F@!U�߯�F#�'yWWO �͆���5�X�IR"ؐ$�X L$"��E��$:�) ��X����$`����I��`��0�X��@�D��`�Hu=E��v �P��xD�A�  Bs��<z�}� ���9�E��P����P6���:��xN%�K�.d�L��T��uLL98�a�s����s`W}���̆姉�0��2�"e��nҠ'����=����\F�6'\�n8�m!÷ �v�qE���e��]�7K�ru���-�7U�ݥ@�,
����m0:��pp�G-�˒����{806�a�Oov�|9� H��RP��P)	.h�����̶���@nC�xMI,��)�2��4���R���?��5T	"H�$@�@�AY$$$~�BE��D�F,R1B�MJB,$��A�"@O7wɓV�����kZ�I3/������d@f�;���]
$���#q �-4��( ��L獺yۂ�V�=�m%�v�e�D)�Z�w�m����
���7-�m�*���dꘘrq�Ṋ�:?q%n�L�6�p{���oT:NC��h��l�e�I@\{B�Wn��&Za2�u���V��hksd8����J&����M /�nl�^�>Z~
 }� u��M6���1%$�@ �����*�F���F��)!��D��dl��2UL�9�E��{���2�tګR`NI;)۲�nb�f㝬�룧S�D�ݲ7X�s��6:q�tX �=P�۱5�c�m���C������/�Y��&�����U�P��7tn�Ep��-9u���k2��NĜ7:����P<A��엙!���-��[���w�\l���b���i%\zu倻�%�f�ݘ���w �����A��֩�qDn(y�g�5����삺����Q�m�8���̀_w ��<��Az��9$$67�}�j�*7/}��K��N���"CQH�v֞fw ���_w �M��׮�vgv��n����ec�Vs��Mnbp]8�P59n�������^����8)�T�&�JR�Cn��p3$DF �(�@������y���p��!��i ���Z�ه���w��`9X�L$\B����Y�V����r�5m2�H�I���ނ�w��;Յ������DD����EA9HpEZ��F�K�=���nHԍ��e�N6��JK��˗w�w��Vd��F�.%!qȹ��Aެ<�̂�^._uazj2!j)��}߾�����O,�@�� z#�}�G���2��I��3p�{�e�<�w ��<�݇��i9$�����?߶�mi�2c��/�Q��6���;vl����t���v_j�IwW��/�f�q˝�>}2
Xy�ym�pf�n&hDc1�� f^A[y ���W��1��4܆�e�V^W=�s|�n4�Q��H�F9��Mf�{�l���{�9}�� N$T#Sb���{���k�Y��̙�',�?A]Xy}�����i��I��H��Wv�cT�9��i�n�N��+��q5�]�nD��s��x��yz���`˷���8��̼�Me�/6
���s�����KpF��4���2�k��a�^zк/�ȋ� ��2��WV_o`���n�͍�E�Lf:�����+o0=�����^����]���˙�om�b� �=έ�k�3��[���À��vj��F3��m��"�fQ��ms�o\:���jg]HF�ZiXR�b{Y�w�b��u���y�Q,�������u�g6��7\�5\�S\�%zq�+�P㝥c^�)���{DWc���/7Z5�kSSfa�����Q�6�'&�n���v6�9��ɱ��W��]�����ˏ�t6�k�+�ȃ� �n&y]��+/ y�ua�Q��f6a��
1������̓����{?I���E8��ȤFo���<��A]܀wsNƓq�PF%��ʻ�+����+1<I0��c%���h��� �͖z�~ 9��8�^�L	(�=�ݧl
�؞��h(1p��u�t�+���Ԥ��[���Felr��ӻ�z#�}C��_I�fe�Y��`y翳�_��o�+RЁ �0"��e �� ���֗�*��+��`�σq@�S�3%�����wr���;k^�.8�M�77 ��@2�eV�w�{�9��Ij	t�7ZYy���Ï��m�	<
rBQC1$��M�%���
�θ�o9�1�J���.H^lՄ��{�����N2!�㡖��v�
��^l���P��2�`�̜�н���|��N)oټ=��s��|pH��4��{�P��/�/��W�cM�K����^k��0�������Ӎ-�E�@�m"bHEI������^%�GF%*0bAD$�	�43Rtv֞e��W� �͂���0���C̼�ػyP��/��ޓs�#*\��݀e��}Xy}�����`�"�p"��A �x�]��_P~ @�|I%���-��y�K�1�N]*˝9��^�/6q�W��-LH� yx7`�a��Ț�v�F���/+�͘��%��'6df^�;���7�Z�ʻ�|pH�nj��Cw��G�#1�s�9�u�΂�nKhm���j�_oZ��Õ��H L���C��_o ���4�l��|�NJ(ҥ"��J0��� �^kg~ќ�O����g�Đ���I$���"(?�������������������?����i�}�!m�d�X�E$�_��E dT	$IH!   s�È@�"��EVAd  @$!$$!F2@�FD@/��D�����H�HH��I�A	!dPK ��S"�d��"(H�$�� �� H��"' �9TD�YJ!H��(
�b �
��Ȥ�0��� �+  HH*R"�$���Ȉ,�*��� �(,��j*�(
H��肀�"� �#"� H�-�)b,�*XXjQ�+�I,0(DQyTĿ�Қ5��'����DQDd~�˚�����w~������iW���j*9������P`)����������A�/��a������?���O��������Aߦ���ʃO����A�OT@A�����?�	�����"��C��4A�	O�~���G�����"`	�� _����O�DP�@�b#��'���O����6��U���_��Pd$��!�����O�y�H8�~x� ��������C��6�����7�~���Q�K�
�*$�$��$�²BH��� H	  0�`$�0��,��!! AH�2
����! "
H��,�ȲI	$�! 	$"� ��  {h�,��� �
	 $"HB$�B �"$�
*`� �",��*��� ��B�H���� (�
�Ȩ �2
#"����$���"B
H22BH�B"0�+"��( �"� (����H Ȥ�0�EcE�DX�E� �B0��B �E��E��E(E,Q*�DX�@Qb�E �X�"B$�DX�P�UX1EB1DXE�Q$EB*�P��`EP��DXAQddAP��T!H�+E��E�$E
��H�a#��*s��~��{33���=3�$?��������A�f�" �h߬{�a��#��@;�=��� @~Ϙ_�?\A����� ����
@� ~m\������L	�����^��}c��|���#�z�� @#=ȁ =�~_��	�oa�����_��H?�AA��������{�~�$�F�~ {y��"#�TG��"  �8O��W�I4�a��TAhBw��L���P�2�AE���=OSO!�F:ӷ�3��?�O@A����?���7���������?����������8?���P����2~�=?g�8� G����>
�  G������@A�0QC�������|y�����>x� �� ��Ȑ1DQQ���}���{��`�h{�D�9�� ^�^#"G�<�'��h}^�s��bȈ H>��06��o��������H0D�������=��p��g�w�  �����t���4��`{k� >�G�?u@h ��G?�]��BC�(��