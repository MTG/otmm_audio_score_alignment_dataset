BZh91AY&SY�����_�`x���� ����a�^}  $   P�  � �҆� UF�EM
^�4 *���C�@'Z�� )�&��R  EŦ�Q�T@������J	k)A "����	J�TR���		D *�"�B��J�Q�D(�)DK�J��  A������ɶY���
��D�O�Ip>��Y���=�6)����yvlt����=���a�X;�"� ���n�k﷾�厷�>�ڛ�|A���M�޳��]={�g�Z����פv�em>���OY[���Х*���z>�]��{�m�|�� {�&s�HUPJ�TJ��R���w��*���{��� �`tw`Ԋ}��v}uD�!�cAk Y%�G�G�/`<�(UQ>����@>ǥQ��3�� � ��;����0��a��鹀zK�< U(� ��y�zUU``	���n��Pu����>���.�ܤ�G�wX�P��>/�X91 ��}���,z�,��d�R�6g�;�{�9�����3�*�U���@O}8�S�Ua�'�;�O���bjz8�����F���h��=���}���T���s�@@�:vA��n`P�nP��Z��7X�hs� 
��x�JR�HT��]��}�_[�d(-��l�#�� ���9>��a�r�g ��R��8=P��X{���nSM�����c�;�����T��;�����';���
 PP   
      
 �� �����F�@ �44�5<ʒ4�`�ф��j�*h�@=@4     $�"T�F   @��J&@�Č�bjyOH���M����!��?Jf�     )�����/����}[>^y�o�o����z��EEyTAS�DEE~b���"��Eo��X�
���)�'xA�����S�����_�_�4�PS@P�K�<K��'0|�>��_�R�}@y:�5&ѐC��I�A�#%�=I��Ժ�R�CSըWR�.�z��.�u+�]O�(�MJ�P��O�CySP����ԉ�MJjCPƤ5#���P��7��`�.���M�u= ���� � �JQCR�j@R�jS�5"��G�&҈�CP���WP (!ܨ�H�E�P(jQ@)�5��Ԡ��.�T� ��j@25 �y��@��y)F��iA�JV�(����U)5 ¡�) =�C�<�C�D<��T<� � &�5"�@.J	�+�(d ����*�B�l �C��R)��]Hd�J�9!��@�?D:�5 {�=���=����{�Cܯ�x��:�Ԛ�R�)@jRj]@j �u!�H<�$9��?���}è^��9	�u��MBjCQ���WR���䚄�Hy-	H&�m.�ԀjBj�@z�%5�^%���ԻɩN�R��l����������r^�2\�ԛ�I� d�@#�K���Hyu+��y	��H��r!2��a�@� d�@o s�(@���B� �!�KB�C���2R�@y���Ө59<@Rm9C��R�R�P���<ːd��Nu�j\��rD�$2SI�5	�5�]C�K�i2R�K�u/R!�mC��*y yI��"jGP>�R�u+��NҺ���_r�5�����@��S�H�eԺ�p�PP��JP4	�P<��<��D�&�B��@��Ժ�uĺ��	�@�Rd;ʎHd��@�HjRd��KĆH)��2cP�5'3N��ɩC��R���B�PNI�� d�@B�Hw+䮤��! 2 h�rG!r�2W$7��i�)h�<�$����{�����<�%rW�!r�x���u'��r]�y&C�K�����&�5!���5#�]J�WR���u j�5j��\�2%�^-�2!����S�rr]�!�r\��4�AAIGs�RR�@T�PJjGPju�Թ.K�B�	�d���RjCR��R�Ԛ�R�!� 2 �����y���ԋ�R:��
jSR9+�� �;K�]HjR�P��#�u&H�&@�ʦ@Kħ��.I�d9!������O$�!�!�.�B��rL��L�� 2�RBd9	��(���O�� yj{$�2�P��Pj5.Й&C�d�Bd9C�d)�	�Bm�P�9&I�sNK���F����RjOS��9&@�FC��&Jd�\��|��$�!�S�<��&I�d�A�Je�&FN@Ò��;��d9&I��HwI�d�C�d.H)�
P�(�x�8�u�3�5!�u�5�5.��Ԧ�@�(d&G�d��C��d�C��.C�9��d�.HdA����2@� �2@�_VH	��S@�CR�R�]BujCR���y��2�_�k���áKU�&_~|7Α5=�]׭b��Cw��g~�g���}<��bt�M�a��ߕ��_����W�kcw�˫֘��z��O	e5�<~W=�m6��s�.��ə��+��69N�S.:B�TP\\OU8�>���oݚ����o��qGU)sC=$B�+�~j�aW=���b��X2b �OZ��>��E�#�����s�L��ފ�m��ɉ�����8�Upz/���+�����
�-��b��һS=���&�`S17>������w�%�O]�t�"��j{�^%]�'�#(���ȓ�a�(��dS�����j�ܳ��/�U�.�>nձ��Rwʙ�]D�sN*=>p���B�+uM����y/J�}}�x�U�sگD*�=W~��
'փ��肋�CT\�]G��8"ɕqp�l��a�F%�{�8�f�p�6c���0�`�o�w�/w�p�La�/�A3)��Ae�H)<ǽ��_3A�n��a�Ǟ�����E���TA��u����ĳ!�hn�4f����1�=�N��t�y��������Ofa�|{/�OR�jP-��nmɩ|���4�5�tscp�/������3���XW��z�(�Z�i�{}�}��/��e��8e��3�"u(!�6	YD�p�ph�K�}�����n�]aR�6w��f˅¬FG�����9�aq�)�NQ��CG���j���ꬿ@����-C�3�Ƚ���X>y��y�1��k�SϥHu!�M=ǅ3O�Ĺ����R�<�O.w"^6(�㘖��ćR
O<~�N=G�n#��
�R2H|�����۱�n�7�9����}�9�C$��=�M�2G��[O��	�<��<n;�;�Fr����<2������<%b �Hx�FD��9Z󏗸�D�Oiq�}���K�M�L�lM�!�
G6r� ��
ì����s�=�������ؽ��.�,�rK�\m�����Li֮F���0b^sƻ������+�,�g���M�c��3c��2y��<>=�M���i�cwq���pDq��s���4�C]�^�6,�'����Z��Ho�Szg<�<� ��\�sv�q���\#���ɔ�s��	:3�d�
����l�\��Ä��L7�Q�<��ǡ�P�=������F�k��U���<Lnw>>�yi�l����
f��;z��Q��YT�_dć�����==n��aɩs��7��t�t�y�19���䰤�/�u�R��Ʀ���iC�J���8s�~9@���b��FqH;���o�/��r$��ؙ7YL�S#]�ˇ6��1)cX+J,��1��^a���'s��1�\�M! ����q�6lv��ĳ��Y�0���pO �0i�eq��9��&%bE�*�3�7�5�\N;�bZ,f!bF
v�s>5�]��8��,�2N�UaP��s1�*\h�SG3�h�5r��]��D�j�rZ}���J$��f2̊��W�&e�*VY>�2/Z3;��|�y�;�z� �s���4Әd�yɮ ��M�.���EÄ�����sݮ��yV�,Fft{������z��Oy��v���q�6Ȣ!�{�{s���
�D¥�4���;�����s�����09�8%�r\�nzs(���o�~��di,e>�&x���J�i�:w�>#1�J�GԼ��dxp�Lu�a�>�ҫ<�
�3���9��
�P�3�f\���:ybs�l��Xh�߃O2W!�q:�^v�>ڏ/pJ	 �q��h$C-� Ġ����YXb%^W.6��Ķ���.�.fd2�����͆����j��v|D5O������i��¤1 �n��ւ0���RDA��L�Nz{�}��y��������o|<='|yP�e���+"�t>����x����2&N \���sp(���y�m�:�8��5��y�<�:�12л��7Q(T���U>L!����*�����������K
�=S�Le1)K{O&�8f�/<�m�8��q
j�w6O�������wEod�����c���˚n�ԩ�;��6D�[�]L����>^����T���U3�%abT�ejk.�p��,��w�ý��7 4��7���R�eN,eDe����Z�xa����Qwr�C��Jqy���T��j�D�2��J,�#�E��e6TVE�s,8��+���"���"��Xq5��%ac��L�����X0�#+Nz_4㼲cC`�TD)7̡��g%#QMD���Ȃ���u�Ef������T�`�Q1Hd�����,n�č�EN��,�J���	A���f��,+DJ�й�oŸEu����6c��T�:�����*��~=7��x�iY���aN�������R�sF7��nЮ59�8{��P�x�.JNM�����|��v7�`��������Y���sbh�jf}u=&�%�̦p�gx��J�%����aZ����z{�3�?dJ�x'�syΑ�\|�4�I�����hFŘf'̗%�n�T�%3L���Y9*������dQ(�4�M1D:g0����rHB����T3G&��i��8n7=�|^�%����C]��!Y`�&�X3K6;��|s����Ӝp��m�{���o]��ݾs���bC�
�R�`_���Q�7�f4��Kib�C#��˝���(1��~�i��N�sx�QfiLg\��0:m/��39MW��|;����U�;±~abq6"w���i��J���2J��DW��Jw��E/]��{ܮ�~�:�_>���|:E!�!�IS��>��ӹu��4�	����]GlPE�=�^hP��4�+�w��;a]�us�e�surF�qN��T+(%����wt�/y���h�Xh��Y��a����<:�e%�Y^����{�o�\�A�������K8�:� ��,�`��Ϗ��V"3�S�V�\e�����\���VǃԩְeaF}Bǯ�uTw��`d|%0C�H(l\ǝ��.>�z��+fY��0���Ы�Q�be������D�k�RVWm��E��Lܜ����!ôA��p���]�t�)����l;q����iєK������)�;�#��f
7�C6s �;��CR�Ԃ�������M8�'mQ�d:�1)��r�5�k�
�����iMB�'S���6�˔��`9�njr`^����MK���w�p�w��}���5���!���L�CZd��g��6��[�揊r��inl�A�'��7���;�Y���V���9q�KYA�ˀ�0.�A�Gw��$��������H��9<C�
Ś(�D����NF�p%X�騔��9l���ه ��#r���)t(��V꣹پU��0�qsɂ�L�K�^��y���=�x�v���f�u��i�o���N'1<�`��p�OG�x3��9-j��R�.���/��C���:��i����w��S�C���xO9<X ���9S�s�1%l{�њ&ac�]�PH3�*}L�1�'���X�6�OA��	���èV@9�D�K�����򾂾.��)JR�W+#J��xp�qr�K�G��d��Y��X=��9r�a�9��P�v�8���]�s�7}yu�xq��}�;�3L��ٜ��aٍ0@����giO|{2��)*V&��D+(��P/��m�y%�r'5�2{�`2�Y�dOYd��#��}e�[)���af������=�R�Q>V>�V�j�������.!L���2X��}�&%v�t���︣���O��xv�;Q4K�J3_z��G%A��+����R@��)�kb�[�<8�)�N�s��0֜��{�<,�D��1
N��c,��&%�v�$�MyeEZ���ި�]���9���m��rq�lLn�GGƂ�į���Q��>�k`���3>�q�q����F\��WSD�$<�brue������|J�C�ÿew�眎gpK�r�-4n{Փ��ύ����b(>���n���X��b_y�2��7��������nxh�jO�d��]e1���a����&�7�=���p�s+�,��38v�eN=L9oa��v�-�P5�������q�D(��
��b_G�-�>��}bvˆ��F��n�������O��}_y�7�NO)�S߸�9���o,	���F3w��<p�s1]�R��C�Hk&�y)��:3r�ƎA��&pe��e�1LJF��#�������&�z��������CK����Q����>4*)��E\u��8�:x�Ni��y���3z��2�flY��Yp���Λ������y����m�g�->7o7o���bwiVY��H�39�\w��t��.�&����[vWs4�������	L��)�^`�֢!V1��	�3$�)*�E�ː�V�Radh� $ZFT���0.�C��*C�.y�w���ߍ�S�#
�G��BP�BAɡ�`�y�0�`$���c�}H)+>ID�I�+]I�M�&7zu�q�=��g
��e%n[Ͼ�������{���Z ��xJ�DaeB�E�@A@�en�iѧ���q�RhJdd�`�BP�%A:1*q+`�����8{�L������Ck-�`��1B�X��KnG2���|�wѼ�r�w��[��^��!f�٥�L�1�: ��+(z��7\ʃs[���z�J�95ܷ�s�y��`�1���W�N5]ύ��L�YM���:��6;�9�����zf�d;@���/�{u�Ծx7��a�*����S[nd311�6�h�6��(�lKQ��Z�s��t�%��0O�����0���|6�8�Jၽ��
�0�c����DO��LN�����5��Z��S�)���80U�T�;��TAJD�c4q�2�[�Ҽ�'�IE�a�<��s�g�iމ�9Y����ݳ~�{�׏ep��_w�c�:r��PS#kx��7,y��禠s����L�0]l_~:�M�T�)����}N�ur�\�&&�/P�m1]9�-i���R�h��s}9e4���YCxW.�i�F�+-ȗo���ee��� �}�%o|��W_)a>�lp>�)Ȍ�]�r:�G�]��ϑ�:���y��<����a�v�-e��ղ��d�Ϡ���:k�kt�/��<� ��u�^jt�][�� ��d:�D<pK*1��T�9�
��9����޴�^M���}R@��Nv1�U��1j�W�0��+�a�j}~�L�4�-v@:��"�at��{�;]噖�wq�\�>���]����/UEEP�"%�1��C��8��sc�;R�a:T2�%غ��h|�C;.�r�.�Պ�uZ���!�����Y_<�y���04����a��L*����u�W;Q�1d�g�6�Z j����ml����/,����<����V�=&��C\e�lmD���S��]���|�tz�N�˔��v�T������iQ��KaC]�/�Qk����_0]����fffyUUUUUUUm���*�UUUUPW*�����UUUUUUUV�*���U^��y�j������UUcUUUU]����*��V����EUUUUU�uUUUUTlꪪ���������������TUUUUUUUUUUUU@�ʪ�������������
��+V�PUX���d�V<�]W�������������UF����c:��՗Q4�K��Zj��gɵV&�U�$���ڪ��cVt�{ U�*��5f2e�p1�>���d6�&��*�KT�۫#�y�h��f��2,��M�օ�n�ݪQK*�mU8�m��m[l�8��M6�,Rr��S.���m��XJ�m�$è*�X�<��i�.	�N@U��5�@Qb;6�R *���]K� Z�^
��nj��<�������V��-+UYA[+R�s Y�����5`[��b� ��T�N
�����-��ٮ�Y6'��{N[{��8v�i�"�[T�p�WUT8�`��TZ�T��[4PU[Sdj��)l���*�`� �K�^�� `TD�]tΌ.݂�6vk��h�*�y��
��UUbj��l�S�{S��U[l�*����l؛ * m36�u7�s�90��qҺ�E�beUJ92cF�W
�*�����j��ʫ�P�D].���	u����MN=���춣��7@�\s0n\���	]��5A�20B��v`�j���������,�	����kn��4Kp�Ʀ,JQ]�upq 2���WR�T�	HUll@#MU�v����e�p����k)�:xl��v]d�<�km[jU'l��uu�N�AU��ؘR��R�O�6���%�L���U@`5�kB諶���mAA��~���]T/TV������y�����sj��ijP�,U UWm "���e��q���qۧ5e毾{�;Z�jTM��mt;�T�;�T�wr�iĺʜ�v֪#�S�e��3�qN�Iޖ=c�f�k������Ү��*�u�����c�l�g���lщ�.��j [�-��
���N�Zf�^�mmuUUWE�GgUI؝�!#2���bK�Ɔuģ�����ɵUJ���r���H��^ܛ[S��<��6�`�N��&�C��x4��&���=8~�Y��eQ7\�κ�bc�*Ca�]SMMxX�Xؕ���iz���˴&�Z�%��Z�6��YYuI���m�ͅm�6�,�`�n;q�#ir�8nV�[i�j�q���+VL�.�Z��Tu�0�Z�=��.��m��*�&.��F��r��������5۶� P[l��� ��{��U�pܥ��* ��jcU�C4�� ��ª��GLbgT�	�Murt���:������UV+U[��q^�����w<�l��_aPe;����bl�y�-e���5���.s��7��7UUU�V&���H�廚��-�M邕
�
���m�UU*�a1h���6��k�V
��Z�jPy��a)v���2���P�UTYfŭ3v�5�j��Tl��t�qA��ctV�;�-j
��z�Gr7I!����"�g�h*�y�����@꺜��X{3v�f\�[`9�B��ǀ�XÅN��^]X��k�6���jt�BuC�4�j2m���4w���i1,��*���6�`1`<6˴0@� je�eV;	s��b[3@!pR rv��G�m�5`�bH�����&�T';mU�Å�@Y[-�l*b<K���g[�q�r�1#ny�TM]U/0t����]F�m���uT%��c�[l�X+��Z��˱�h�����m{�Y˭���y�<����Z\a�ْS�N�m�i�ܫk���X.u�,U@���5V0!if(*�T�]U�ku�,�:�Xͪ�,Ռ�F��p��Ki��׷�����+f�Z�5�e���a��c�+e��6�f-����� �M���D�.�иZ�4j��9T��6�F�*������R���B<�(+��@�Y�@-Ⱥ�)ES�ZK���<��Ӷ���A0ۭ�s�4��;�gV�ۮ��i��ɾ CG�w�UUUMn]\�X!A��[I��4�݌�k1�ρ���͛CV��l�`��6�j�Uv���vY�meP4��fm [�.5�-hL��;J{��5Q]��lV%B\CQ^��i�E�x���km�� o+��mK���m;tPr=R��pE�q�n'i�jCfSqى1,���mv&���AG mUUX٪Wk�l�VT#�iѵuѮJ��IXP�+�U�6�[AVT�#���
��Äs�h�+43�P��y5і�*���Ճ�[x�ڂ��u�N�WEK��W`�+4��u��h*V���m��ꫠ���Zv�4�u��q@i+�%n�)S����Q�UU����uQT�� �Qp	�\ε�����Eƃj
�j�snʯ6�[m6P$�҆�AU X��i�,U�@B�q�æ��-��P�h�t'vĶރTɳ��< /5��kY�m�3���H[��2J��2� �DV\����E�n(��SA1�]����U@�4
`�r�

f�AB��h�'zb����lv6��BL��SJ�l��@6�uЍ�	l����v��*�j� �� t��-��]� ��*����
��UUU]��*�����D	�k�c��U���*�V�j�/*f���!��uR�r�s��p�,61�p�H#�T���9�R��sֺ�Ջem�4ug9vB7�p��,t�#�Ԛsm�M�B͂"-]qǀ#��2f�M�9xLPЭ%ԓt�ex���U�K���}m��k�J��9O)A�2��>�����ն-n�'3n��Y�F+b%��{�EWC%�9ua�m�4#Ƭ�`ܪ+�Ҝ�9t�W ���mP�UUc�[Wl���]���*�:���u]U�.���ê�i�� �8WR��a.����ִgu��w6���LCVـ�V-v5h�V+j �P��L#f�Y�em����ڽUT�Q�UV�t�9X
�+��W;��2�CNV�m���껙-C9�-+�Y��@� $R���ƀٺݻhK':@:� �i��\� �i�WWgi�t�������Z���-�����}�ubnکZ�m�J�(�c���eA-�����+�*�Fe¨��m˕˔3UUx���
 �rشeF�*����)��8W(�pN�s6��ĭ��:��J�Wlb���yv�6eiy�W�m��V�c���?*�ꕩZ���஭����ڠ���� ����Q'	NVV��UUu]h���T�Jl*�m�U@UUUUj����Ry�V�#� nV��V+�U�QV���]�qtX@w޻[��^q�AT�]m�*\���qėe��Ekm�ꊜ2��l�*��e@ �AUUUUUZ�������Wr�Zj�m�*��}.~A�@�ζ�
�ꪫ�@pR��AUT-\�v�1�*L�l8Rl���eUU��2�&��U]�Xl�b�*�)Z��6+n��V�b��UUP��b��UUUUUX��UUt�	�uV+�ڗ; ��A/d;bjaU�eUUUUUj�����������J��ٌ8M��*�em]�W��V*� b��(EUT 3��#VB�St�mUUUc�cn��u���m�'SԎ�8ǰ�Ƨ#X���|��;pnu� BF��;�7B�00��
����cAj
�-���ճ��G��~o)��ESl[UU��We �����<���5U�δ6�_/}�}Uʆ�UUUUUM�8�cc` f\M�T�n�$2-UUm�UPKRҴ͵V(�쪱UUUm��5J����WUT���M2�Q��TE*ԭUU劜�,\$T�*ڪ�iTTUU[mU+��T�����]���E�|U�߇�}�UUU+��8ݠ��[UUV�[+TU�F���m
`�I[)K�Ot6��b��+X6˔�f�ٶ�8.��GfڪT�mi�t�T���-6��.`�+��ت�b����WC�P���D� ,�+�����nJ���jV�άڶ�ۧGM.�j!ǕP$-U���鳦ʪTW6�@�] Gd����P����UR���m�m�*�pAV��#9�
���^^j��1�kX�Q�4�m����s,!�Vkv�U��@�&�3��xn
h{:,U�bwk��C�k�.I���1s,�Yi%ճ7 �;71��l�9K�y��@�6Y�6ѕ43� �!4�;�����0]VHF�V �q%�aÛ���mUt(��T7p ��VZV� ��!U� :��nF�X5A�)�EC-l�$0�t[^T�Y�K����M ��n:� ����ի�K��!�m���"��kKJ� iU��ǵϻ=S�:��F���X� Z\hlMcj e�v�Z�S��v�_��{#Ӽ�-�|]/N6�j��+m�Z�7<���G-UV�[�mkh�D�5ҫX�<UX�lf .��ٕ�E����j�WchU��1A�\�V 6���V�5WJ���TuZ��5Sem�ej�������2���PWi���Tf����'��W[7mPU[ev�+�8�*�ڪ��b�]� � �j�Z��Y��+j젪� �kUTUUUP��(*ڪ��Ub��A U[`r�� +h ���U UUV+�UUUUPꂪ�������j
��*���]WR�UUWT������-��U P����[b ��p���*������UUV�Ul+UUUUUUUUUU+GUUR�%
��m�+�;� �*m:�k���*�$U��EU�(u6�Yp��؛ ��k,�ݬ�,�*��.I�����(����l ������U O��G_ӏ�|b��v���N����L�-��6�DQ�VUQF"(�ɕ�e�-̖�*���Ud*�l�L4��� �P��BQ0
JO��?�3�$j���kBv�H�"�em�
P��� ������*n��?�{�7���ED�QAB �� �� �� �� ��*��(�����5QUQUQUQAT� �����������UPQLPQQDDADDAUQQQQ�DQAETAEQ��ERQQ������Q�QEP����Q UEP�E5E�ASUCeS6���w�O�G�	E�H�`�J*V�����r�D��MWa� ti���3�!�H"�"�o�TҾ�艀�zl=���U9�Aߨ�DU9�D] ��P6�`�}�8�h~���N�^b�)ځڈ�:�B:��|^� ���\7���P� �{�9�!�'Y�&�FR�@����'����"��"��LE	P3%�E�~#�Gb'f��N)ߢ":�]��+��P:��6��*�0�"�
�(	�6�]p�M�����z�Et>��{Y^k�D{�1����*n@;;��==P�@��v����t�f�ζ�8�� �c2���*�߀��@�פ	�0�}�}��T�QS����:G�⠻^�� wb�� �C�6�`����y`�����9 B�h����_FE�� �$H��2�H��&(2,��B10`)�f���T���3k	�6��	�	�]��A�L��$1��'�
e�I�0�1r�*BR$�#J0[h�j-"�b�ČhմIJ,�"�ؤI���a`8�)�Pa�:QO�)������T�C@��m_B��0"w��l H��t�:U]
`x(�����$�B�%   @	���6�B @   i�@0  @   �	Ml4�¢��\�QEQES30QEQEQL��33�������������������~����}�9�9���S13USEUT�˚�����컷ww7�]ou�;��%�E�EjRB�¢ �)fɛ̀�J���B!J"��!14�hф�d
w�)�Z���F�h���y������|Q�Lܳ^�.��l>1�_�����m��*��{��;ظc����x賵���/��S�CU�y�y���P�[�i�l*7����x�㚊�P�f��=�{����P=w���F��żȹ���}<��D8�j��ʇI�̩Mj꠪���5T�}�ﾨ`UWl�j��vQUWm�4��te�
�؀T*�p1����]���p*Fx�FD�[.�rKWCL+	�4~_�i������"٬Wb��N,�Jj�;���y��oHV�[6s<���Lv��'��K;�R��]�"�MK�Ȏ�(��s�r�����7Kj7�.ev3�L[�6x&� ��6ٌ�F�����Kr<4T��"�����mC]j��df\�����Sɚsrv����]n։�0�L�b_�;��(w���f)�-9�X�Z�����3�ZO,Z9���@�t"rč��3R<��:.�Y��5q�`%��?l�Mz|9w~S隻�k�=�B��L�dX�ָ�L$��
{R{ve�.l���lCD.�̷�����R��dYe�����
����8�:�Ľ�R�v�媄�O"�s�zݗ^��p~�ۮ~���T�kj}v^��03�;c��" p
bTLF5T�*;��sSv���;y��B�t���N��<����0�:���&�8�n���l�u�����|r$��z
�B=2�� Ư�w���.�e΄���E_�V]�d�le�����G���p� 7Ooߧ�����F�NU���<9���=�م�˥N�qz�`��
&0AЂ@x�;tz���6ҫ�`� �v��y��ڷM����~g
շi�7�����rmn�)�kÓ�Q<��.Wen��v���^���ѣݮ�Ö3�b%g�-]�(�g��@�3 G$�)�Y�gn��\0,�M���:��{�N�vٲ�\�˳���Kv�&�s[����ԁ�@T�&6��:��d����7�ִ	-Ö� p��!yOj�;r׳�W��b|�6��YK��Ί�-�:��٥�\Aղ�i-���N ���L:��(��`3��;?s�~�~�.v�j�Q�dX����5��5nٮ����8c,X�����F��i���b0ZH�m�Y�,v�*����n��q8ۆN3��ʣ�rp���x!ö�P��=ӿ'�ۻq/�������L��bp[ml�e�gW�A�q<&����|����u��;i�^��5p�`�q�a�Wj�ƥ8vL�4�3`-T�"�V���5pX��.n]j'�Y'���&qB�_Qx
s�ȧ;|�@D��N�g���b	�(m��	�)�P_:��Z���Fl��{�:}4��ϼ��n�f
�m�16 hb:6�n�(=;���q���z�p�b��,.���ּ�j�x����ڑ[�4G�wέ��*������K�j�7h}���y�9{��%�	JT����ۻ�-��&Ǎ����J�GZ6����Щ�
�q�B��c4}7nڻ�`�6�- �Yin�GL�bmUۉ���^{C�����o���'؆۫=���%�Sƪt&A����'9'�9��y��0c�Xc���26�)���ߣ:��8g�G����<v��!�>wʘ��Q5^}���?J�gs2���"%8�!�$LH�sٔ��da��zW{����g1D�&&f%LK����20J��{���s���g��0�L6�a�q�网t��ɣ�u��I�ј��x����f�f\�]�y<�{�W3eB>�{��@ ��OO��M����G5ۃ������[l���]�uN���d]i<g'�	�ɂd!�L��mxG�cK/�������>��4��c/g߻�w}����)�Ē-s�=��.+���){;쬇��C�RD2\A>�����R�s�y�ﲗq�4����	j�""iI�fL��dR�?c�W8�fԥ��""T9�s<���V�2�w2p]�����-K�^����+n���Z�۳�4��^c+܃�Lgms=�����1�K�z�/7UU6�^ݍ9wܔ��zyY���s�BȘJ!L�m��É��z���O;}̮{�j�B�c3Q 7��9�%W=���gs)q_$(�7{�}����is��n|�G�zye�G�"�f�C�)+;�K3тW}����d<�e�bș�c�TD�nM,�q�.������yy�ʢ���&�pq\�	+����%�ͷH�j7qrm�*�x���v�6���n&]r
 �>|����ޔ�;���fL����Z��-
f&*E�̘�s��N����l`���*��p�[���7�32�Y��K���o9�#���]���U�y�%6�������M-�+3�}����;�N�qe{���v\9��߽�y�y��o��,Hfm�Tg�|�>��O_����/w2x��8�]�f��r7�Ys@<�7��[6q�����a֧�����c���ƅ�L�o���ĝ�fR=�8jIｳ�����DR��BQ[���fdQ�����{������3)��bA\���X��'U=729�����ϟ��3s�\�����N)��ݚ��DB��=���F)��0����"[MC��g�r��U/fd�_���Y���/�>��[X���&Æ�A)�f� �&퀩�M�3�Z��a-f�.=ac�����br���Љ�ضv���\uZkP�������A���F��u(3�fٸ�ơmηV3d�o:�z��-��s��O��bsl3��E�Y�"�R8�8����&�V*���i[�T[����n��E`:�]e�,Q�	U�Q51��ܖА(�i�ݔ~I98J�v�-uЇ[hD��FGA���������X\����m�&�ʌ��'rG!G<� avnMqX>_}���^����}�y��b	5}�PKA)×.bi{3%+��R�\���z�f,�#�����9�+��u�����kd�g|�	`���p2D���-�­�3+����[�g.�[~~s2(	���K�eR�fOYܕ�.%��i�2�l���=j�e8�Ϩ�[mB� 0�
Hܛ��<�H*�b�SS�����}�߿rg���R��;쥂�i�eÙ�2\��nÝ������o� ��ʠ�A&���ȥ�X��� �T��ڒ\K�t��6[~9��}K��+y�f���S�
xL9�yl`�v㾢�w&R��e.�1�K�$!�Lˁo8�8�{���rR��ON���uw��PKA)�r���.�(��U��]������y>٦�}ΛJ[�k�EʶBMeЊ4m5nh�b�v0�)� ;��YM�����VV�&b"NU�%_�N2r���/{s��B[�=�0M�H"L�5���H�_�\�da˾���[p���	�J	�+/#2��#V��j<㧲a����/<��3(p�DL@�M*�fV��%wc����W:��B��S(%��D��rV���J����0�t�Þ=�e��\��sFAݫ�g&���p0G3wW�km%Ϸ��Ή�p���,����>���ﾰ��<�|z"S!�I������W+ٙK���Y��V��^���-�S�.\�Ҽݔ�;�uηӓ��W/��Ʉ�LCf�ۻ�����/������6Bj"���G��/e*?<�XL2!�D9�"i{��[đ}ﲖ��Y�r����ߢ��]�V���uÕ�jWMS�9M<ݭ�M;^� MF�M�n:�n.���w�~���d�U������y��L"%71 ә�ffJW��=��}�Z=�B�ʙA.e��9W잝mtTe�}K=��30g�d�
HDD��#e�2���M���d��8�b�$6Jr��_s)a�g>�w�w����:q(�HaH� �b�~�����'9LϺ������*�������.���	Pv�Y�r͎�\U���, ���cl]W���`���qP�^d�9��H�ͰXg��m���un�h۶� �F3C�,k��qi�n�v�`Jb�f^5]\[�V���I/=q���q�WcqYW��W�%��0	��`8x��'uث�x��Û��h�l�Жk�n��p�۹�O�I甽�*;�i��ۗ(�tx��j0㴯����^���tn]r�@�հ�~54L'؊L�	����x���W��q*��J�y�Y
LCd̹d��l�\ʿz��̔��<�IB!����U~�,�d�]���;��z���B���%�C��v���W}���:�9��x�f$Q3.""q4��rﾕ}}9�~�Ͼ�߷���#�6.����%��Q]��69�
r^�5��U��:]wkuuzT�sr���V�����\�8�nliź�/ů�sM��/+�C���س��Ip"X�cJ�1���~뮾��ys��~�v���,&H����M���2;/݌�:{ϓj�G�L&9 �&f&�{#_}��������8u�Y3
"&!�fY1(�{�}}97}�Y���䍜��k�nÖ�yKn��;mDHj�,��S�c��f��-*I��e����9!�1�y�Jo�=4�ْ�}���i��)p�ʔ���9W�e2��2s��}}5qc�-��l�H�̌����y��;�d������Gw�qEUW�uws3L��UU����������v�������{���8�JP?�/��;��Wýt�0?�A�g��ye����:Od��:a�ӈ��e�(ࠥ���	PNL����/�����:�7�N����6�'|�p�	1#�H���AD{A��{l(y�;a:��y铱�B��7����{:��~`R}�}��y|Q��#�6�h�]���� ��2Z�4�)���P�2��i����HB�")�B�h��́b{���
��6㶬c%������oz�|*LYi���l��������TXR��Դk`؈�����^J9����[��"`ܭ�<��4C��e�c!����mG�e��fM��q	H��I�p� �ł
�h�\� ���0���!����w�x���-���7�3B�,A��b�X��-��xc���H�"�0�	A w��N^f^s���F �D&d�i`�.�D�IIP�����S"B���WX{�	�����a"Xؖ ���UIwUrb��|`���E�4�W4$�P���c8���	VkH�� �
JR�~�g�8͉"�aF��A��mgc0���Ĉ�PL�uQ4.K�%	@'�]�D��cF-#E��cre��-L�a�%�0�Z�7��g\z�cn,=w�UH'�^{ �z4!����t�2�֔Sܩ��;�#ċDʠD�,��(�"��vv��m{<�@	 t��@~�x�Z3ծ5͜|�Gr�O�2z�w��B�8��>�'{�u���ش��{��}�ԔD�#=��g��f�ݷ3^,�'�j^{�ג4/���`�4�s������榶B�\��v���Fm�&���0T��wy�u��=�>t�W iN�w�^�h_��\F��
����d�a;==���wn��N'�{q�N�����ɴƦ��MKf���݆:e��v����v��E�Xw�~��:��s��.A�i}w�p:3n/P4�64��	p>��H�	��Q%%���+@�Y�\�@���0�y��<�=vC�P����:��J�>{o���s1�;n��s^�*a������� s�y�pD�λ���&H}�����.JR{��=��fj�e�.;ɻ���'�+����'߷���hy�ߙ��)@���NT�!=��ri(A	��#� �!��ǀ��
��Ѹ�ws!{�+�%���!���$��X!�s�����3����Л(�ֵO~������vBo���q�]�ne�b�E�]�i�ɚgJ��6�����R�[e��;=��h���ww��ל����p�Ҕ�}��H����n\�,<���:��+ �>��f��ۣ�e��Z��)JR���kc��XL���wPw�5�j�)@����ʚT�q�������m��7w�N��g)JRz��~r=JR���2�r�)=Ͽi8�Y��}���.�3n�rAd�+|���	�a�LB{�w�Ҝ�>��%)N��{R��ޮ����Q�9��\��A�/nN��JQ�d;�k��R���q'��w�G��iO`��X�����ٸ��v,E�+���<%��T�g�W�z�v�]�ι��u�w����JY�E�n�ۄ�S9�T���{O=C��yϙ6W��8��j�.2[b���f�&Q�t���a�km�:�J4�x����5ݝ/1�(�C���7a6�7 Y���i�n�.���/<�݌rպ2���gVP�3�$�Y��"��J ��i���]P�ff���K?��[-���M�M����bh���E`�����o���dle�� ^,kW�į�46��\ʥ]�����=�~�q�Y~�M��({�?x�P4��{���d�#,���B�ldدgQg<�䷜�k�h%I�]��2�)O>�\R�����qB>x߯�͸k��j����Xy�~�:����'������ބE>�@y��6���;��r[�Ky>�ﾇ���h�C���ԥf�� �<��\R��뿾��R���6}�2���wߞ�����IOL��3�sJn����Ad)}y�m��)@i�=�:8R���>=��Hy7�p��D�'���{��4�~��)��T�!yH���v7!�Q�W��2��nz�¹�[HB���:j��oy�|��)Jy�v�)I�]���yJy��pഥ'�{��JR����m�K��LKt䂁��������G@)�lzF���4����' Ҕ�����)�~�ڟ�$5�G|/dA�03�B	nf&�,�%����p�%(|��<�<�����ڒa����'Y�����i����v�����)H��y��_Bd�ߟkjR������R�r{ϣ�Pr�O=����p#��5�^��痜��ߟkjP9uמ{��R���w��)J_]��/2���@��Fa�Zs����J��<q"�[)�[�Zd��2
�\�nוD�s��&��ƶ�m�
R���3\�P4�y���ʛJR�ߙ� )�)u�f�@�h�V[y��ۦ����m��'���}���� �
N�){��}������lL��Xw���	��+ ��kf~�6���7w0�8dO}���q�XG�zf�,���'�0r��w�2T�0�Z Jp�L��0��A0�J1P8�4����f�:��]�z�J�&�q��R�J}�~��k�L���s�GY�fҍ��擨E�W��\�>eA��}�ԇq�O�}�G})���g9��+�.X��qn�Tr&�7ָܸ��I�~���J��?=��R���6��)u��R����I��=��I�1[tU���1���TH�\<ط;J`��`�`��L��WW�'tRv���W���3zOP��P�����(E'�}�ǒ�)u��w�ox���矸N�l����w2�cMݮe(|��y��Д�<�9R���y<��#ԥ��o�\��y�)�8n�C��Kp�Mrj2�s�K1&�7�5�)JO{����� 4�{��H,������ ��߯�m4�kf�Z�k\R���>��}��R���w�*R�^�3����>����L	>LE���:�d*HeȘRK1T;י�}���Y�����5�)J�������N:�d�yy�ɯ9?{���%��|�^�u)@���mJR�����R���{���[��,	v��T��
�m�9���h�`�F�l�b�]��N���h�v�A�����P�]�r=K��`m��R�����9��)2�����)Hn2_O|ϴ~��:���ݼ�:�,���f��m)I�w���K̚�9�r� y�i8�yI�O~���3L�f��3v��)JR}�|qz�����|8�?��9/�{�ǒ�ߞ涥'"V�s�ܪ]r�ys��	�AC�Oϵ�)JP�w�JP7]�k`ҚU�xu�<�G�Jy����&��w��WwNB,���߾p?'P4�%��7�JR��Y������NA�h��#��,6�{��{�����ƕ�΃��1��l
krC%À��F��b��Pm�&nЌ��PM�	 �ذ�Ų��K��vv1���j��nmr�m�r�[��kv�p�m@�$;Q��A^w�8�i';U��1f���V�צ��n���<�v��1g-���m�AM��a
.�t���в�f\�����_|}��4�qO �֦�Ź ٳ,���l���~!�|j3���z?����#.$&�%�%nn&M*�n6W�H�ǜ��r��w�w���E#y���uH�{߼��ԞA�ԏ���^$��,_=� ���[��>3n��4�]q�䂄X~��߯	�?ʄ$� u�f�9R��:�y��07�B��ٰ� �����3��]ɷn�ַ��R���߸qJR����t<�R��μ�[����|���){�柷k�p�]�y��p䂓���D���_h(�yߺڔ�.��ߜ�u)A��]o�tr)\Zun6�"P6�J�����;��F@Ѹ'����P4����@�}=�{���JS�g�zբ�n�]�qktq@���$��T�H�14t��PU4ypw����^��k4���fuJ�=w�r=JR�ߜeʔ����݂>]J]�7�ݵ)�$�G~\>w2�v�6�3xN�C��o����d����ӈ��1���0�����& qe2d�H���C:� �J��[��R���~[�����}��C�H���A�����ww3���[��JR���@�=w�#jS�����޽��@����\R����~i��-��*�y��u�]a����\��JR{�~���R���w��)M@�Z��{�ǒ���s~�1�M3V��$���߿v�B(�<�>�\��wy�@ħ^g��,�Xy<���қT�r�A��Le	����nQ6�Z6[��pk>7�{�n�ӫ��:Q���/9;�9?}��x)C�{��)�z<��R���)%g8��F{M�31��ˇ1'�){���q�~B���n޵�a����u��}��R�����qSY�~�����sx6��w7�N��5�)JO}��x=H~�� �Ր �CLe��Z'���BҰ�8#����m������q�*S'�����'Y����˚�v��uqJA5I�����2���w��(��}��Cq��%��l`������s.�-v�6�7^��E���~��/qL�O/w�]��j���-�n���qۺ���L�D1��}s(��{C�m���D�h�S��g�����d�'��J�YT�Y��]d����y)Jw޼��)C�~{�5��ԥ)����|G%)=��m}ݘ�-һ�^f�:�(O~�΁��(���)I�q���JkY��9Rd�>����C��~��9�۵��5�ݰ>����=��R���{��R�"�(����y�n��T�����,����>�>ͮ]M��.��o\O.�)����8��S$��<�c�JS��ޭ�_�u�~��9�~�6Z���H�Ŗ� {���kf��������ޏ���~���d0����7s6���72�ʠ�2h�q#�\��	�f��fҠ>ԗ4݈��K�pK��0�r���`Z6q����ڭ�q��H�C	tгb��I��L��8�"��UUO@^��In�ٗ`}���s�I�M?nM ��K�p�Q34�
@wsv�\K���m*!��7&��x��\�}�BfI �p�1n&j��m*m{7f�.s���Fwٗ`�i�I0KR�f3*��s�8��g�݊��$m��f]��q-���Ň��@g�߅2��)AQw}Hu���s��-�ݮ��oԨ��&�j�92�qwwww337sv�������������ݪ����{��{�;���*���J
�)h_�"�{LTĕ��*�?̘:��Y?�@��ydiSߙb[����Y<�� ����ܞ	���2s�X���$+��5�C�
��]iC��(@��%NE� �ptb>s��!4̌t�O�����$��� y}
CP��6���I�_���8l�N�M�{}��.�7��舥P��Z�A�Dv��b����V�t]�3�H��L����SںR���q[lm�S�=��M��άv��Wl���F����] �5UJ���U�UPuҍWUU�k�3�r�x�;�ו)���
R/	��o��|��l������Z10��9%��l-?������Z[<u�M-
����xK�j�F�&>i��֌R��`�	����N�x˾�'�p鍝�H���7%��'�l�u��VU��۰����v0�9�k��$��3,��8 �fb�--��c狷�ۗJ�s���Ѱ�̤f�ᚦb��i�Ju�^�g[m�gg9օ	5��9�@�]�mC�;x��vJ�Nn�ƶ췑DUY˕6�nkؽ��L��ҝvM�[S^b��9z�m
m;vuQ��J'X"Ѷ�J�٧��ˉ��)4Mh�#m(�1hJ�4[�hDƻ�J@�����ܢ��fD�bE��� ��ll�3kS����B�N���֠��ɝa�lV�m��� ]��a�/�;�K̯;L4��1 ��ۗ&p��&�z�0ܳJ�N�^ݕPا����gI,FZ��9�D�8�UU\�b�^jw[7�8e��K��b{Ym��v�li-���l��2���2��5.9Zn�k�	�;v,2E�Q��\�ji�8�d�η&�,��=Ev��%ٝ�5#�h�Wd���HfҦv�A(ţF�ʀ`��	˺FݑK��AUa-C6�Q2Ѧ!��M`�6���p]�,cmv�a{`}��խ�&֛gWjA�!�:\�e.Ԅ.c��b`2�x �Vq��ݴS���p�VʪHW�-sַc� nY�;=kcR��ƺ��+ɚ;rnΞB%�2�l�3s� ��Љ�NnNᇶ��^F�L��d���6���H<�8Ѹ���Ad�n:��m�Vj�`��h͋��%��L���c[.��zcv���VUņ�%�Sub��%��5��s0[*�0բ�Z�h��ɫ�OJq��l��W�V�j�{b; ���JK�X�\���Nw��'��WnT�� �� ����{P���H#�OPU8<z�z�T���5����{ߗ����5��׷ߑ�yʉj��vf:oÉ���S�	��eҊ�x��Ql����<�|���{vc�X�E����	�w�����K��Ksu���F�r�mSa�|o��:ys��,k�0ܴN����{r��i8;rc��'��i �^�l5�P�5�1�������^�6����i��fA��:��͎2�.	SF�)gi���4��j���f,���6���[C���$��ǘ�_���A��:��w��d�%�6"��i��u�������<��Y��8���4t��k�ᮡ6Q�2��@m��@b�ؑrpV[)����IwruԾ/v��/W2Z�|���l�@�d�bK:��}LC]��ؗ��R&�D����'J�$...l&�@wф�;�{.�|���v����2���C#{oݾ��M��$�ĸ���(�۰;�(�S5�-�M��Jfjl��Rwӄ�;��/z��'Jq.$7�/nM��y��QɄL���(�n݁�\�8�6���rh�x�l��M�"e�@�1uˑ��6�4�#��=�(�n�,�,v�[��9���ilͦɰ=�����@��Ё_cĮ|���.0�ٻv ���=�T԰������=��8��lL�32�D݆)����J+3 �	%D 0� �ZI)��e%|�#�P9.���~.*�y޺�:5���$����s$��9��sQ3`wф�y��w��nl����&���_�%Å�Rɂ�p����� +�&�)B\�	5��h��H��e�݁��Ҁ�8\��M�G�Z{�˰�ij�=C]�[r���լ� ��c�ƅ5�$�e�m-�Ra�Zº]��,N�å�C#{�o�~=�����a ^{2�Ĭ��ҁ}Mi��&A(n�f��G}�t�	�*���V�����_E��y��r$&`p�E ;��v�'J:���}���?s����$s��IbK�쵎���߮�l��H���Bb� �
f�&j�G��\_f�� /g�@�!H\K�'߳*��Ѝ��-Ks3	�
J �z% �..'Wؐ/=�v����x|݉ywnv�yA�J��=j촑�1�������e�a^A��y99(g�X�vwǢ���j����`-�N��ŭ���M����3.TH�)�8���۱r����Ҹ�3۳`�ɥ�պ�6%�&��L���(��4v���$�}�`	,��S1�e1�2�ĕ��ė��(3�٥���`��۷b?qs�{RV����=k�M�@��q)�u��e��~>��&�7U3S`#ٱ#o�qqq4�}���>Y��B.�nՁ��r�i.%�ZjF�̭�<�t�,6W[;��&�n\̮�5���������Y(rȒ"(���@��Ы�ͩ��J�/��@m���I �HA.bff�̘�K����z#ӑ {��vs�@��|�RܨS0���-��ʚ�D�8�}�ŝ�,��ҥ���3E2�S)�V��M���Ȑ+�f]��N�	p;�ͫ�ų@@�)�H���{v��>q/��� /}�5m�~�H��eqB�s����v��c8�\�ōe I�mǖv�3�;�s�m���t�p���&W�X�Ѭ�[Wu�v��IO >7����p���!�3v���K��M�.`��MMeZ/�{����Gjқd}�X�8�v6�X֮[%��lnz��L1�ӺF{��Wl%����+Kv��%�P����M� ��M�b�yu��7ZpI@ �:�@p���m B0!�z q��x�<:8�����Α��#,g�קH:���������b#�3�e�lI$�6����"/l:�~�Ҏ�n7�69�7�.+|�.����j���D��2�"K �3f� �D��}��vs'J�K�:��alJ�b�2�j��;���s:�s���N���j=��
�,jS�"(?����\��������K �w�4\J��D�6���L�.ƢI��㎺�<󌹪�;ʛ�w����A�Ȑ;�s.�E��5�tH���I�5v�� ��k��h���Tu�e�2�Pp�ϒrBM,xo,�5�Gs�5⯿���:����a��e��8�,̝*/�{��Q�)�obn���=_�.R��V$����~&�����ڂ ��w�]����[�q�bv�{�q�$�������10Юu���~�����ٓ�8��q~̊ �x�@wPu��3�)���|-����9���y�{e�y�"�/މ.qp��=�`��bS�#s�s%o��T���!�}���M�2t���{9Q�ɡ�̒"�v�����Ԩ��hk�Q,�70�(��e!5�9�#Yӣ�Q0@���sR��� w=�s6�䕥�&Ǿ�����
K����C�s2���۵s�.$�n���36(���p����A �q#Nfn���Ґw۵g��.J�s�\L��""�$�$" �	0��=0�'_D���=� �nk�J&H���Ĕ.q2��4�z$��.�	%�����y����)�m�M�A���0��K���^r9�� _w&��!��l����꒳�5�,�+�j�m���:d�ۂ�w4<f��]]�:3��m$�t�����b̓] Z�>���#ɨ�F��dlKNf�7$9����uĹ����&�&"���.�Is�M�s������l���8we����f�/މG9�E�9�`nFk�cg<jk)Ǝ\1�uQU6q.'��?nĂ;�ݻ}���?qq�:�ĳ�=�.*B���w'"PLCr�pI~�m؃r3]���4~�Uo�Q���ˠ�-h�Xm�a��-��r�)��l�΃-����'rÝkj[(;L�~[��� �w&�/މ���˰F�CR�b��t�}94s����Q-���v��]}�q./�\Kn�����D�q6�����}��\��3]}ܚGc��&�"[�",(I.lu�6��f�S��M��ĕG�aR��Dd��Ipܐ�n�܌�@|�8�}���옔{��.�����9ūi����M&U9�%��@���0#T2[hP����.��3�̞�pX�z댰����>p=�q��SC8D��Yo1P�&G1	�� �vI�FhSYF�snwK���mpV�7P���98-+�.�Լы];	Q&�J$0G6K����j��.݇<����LvƇ����Ç���f�].\q]���[r�#��j+k����0��V���[F���O���M<�J���#(�M�qc65��^ͥ�MRĠ���jJ�lZK��Nr^f��%�LC	�f\K��:��TЀ�z$����#���}��:�g���>0�-��TUM�w2'�s��}�V �c~t�߿���?z��B��@%v�5���`nFk��q&{�SA���:����$%G�q���9Ż���{�4~�I���q.F���������[q�9��@�ɠ8�E�� �w}�`k�=)��Ӂ�k4P�Z���A�7k�I��{���hI`�Ѓ�ftm�h|�'�����i����M�M�f�s�v�f�%����Ѓ���%C`8&�䈊=���.]����iD��pBM1�665(�,`(Ԣ(DC-5	p�he�)�a��E+DKB�� ˉ��Rb�,�����v�A��d��C�L�s�޵ʮ�=�|�kwߣ$���{~M��
D6v�(k�ؠ-�ܚ>���s����D�^�6�/�=�I1!�%L�bb�7���}̊=�d]����s�)�ߢ�_щ��b-��TUM��d�y�$���U��3b�7��4��=	� jGiV��6�:���w��SmI���ll�qu�@:M�÷���J&�!ALQ(��"U���w��y;07���qqSl�zT���I �����Ձ�3b����ʚ_�*i�ѹ��\\I�Ĥ�u�>��C�Jp�p����}�M��R4���e{�uUUV]�����UWwwwN�������.�.��n���z�	HCi�9��Z���⫞�z�J!�ع��N�6����X�Q,�c��`�lP8H|RWh���;s �`ZJN�R�6�
��
�@ܨ`�42\�<d�83��d-��%46B����4�,p��R��o���P���4��wvn��7LEP&�@ѐ�&��fRQًa�K��m!m�4ky�b$�]HHd�ON�s��b�`o��������F
��e��%)4Jhwtû&#��e��I�pl�wmnw�!���ƌ�0DϦݡ0�CdJD�i2JPEF%���Y��@.�J��O�ہ�)N���c�Q@hV&<����2��ZkHȫ�Lk�K�88�L����|�w��������R6���
��@�D��1�~
���^���@���]��� z��PO�;[_9>N||�V�c��v3���uW��?$�e�o:�7��@�=�L�Ôۉ�Q16�̥ ]�e��6(8�l�;o��c%�	�D����x�۰8��lPw�4�<K.���2=Ӱ�^�s��)Fx�j��^�^�c4��4B[��t�%�Kn~Bk�kӭ�W&�����}�E�/�w��|��3�^�݂�1��Z����T�11@�l�C�<J�s.�י�J�5?k��1.��jlli(^f]��PWѻ�Z �����
1�%��@�����z�����l�~\V����92,@�$��Hj�/li$7{݅�H9B�����y;��{f�����m����F����\^�J��d-��3�SV�d��뇭릷�=������clGgG)��TL��������D��}�a�y�w^�\�2S"m�Lݶ)�N��&o�v=��>O�n�쩡Hο7�l��I�d�k{��mٯ���GP�v=�@_�Ġ=�=�,��@q1�3w��6(����}�#��e�����e�s%L�f(}�E�Hy�(�7.���6)6��\�@�$������fmϴ��y��^s78M孌[z�)c ێ@���:k�t�z{URl��������G�8Ŵg�E0˙�B�WQ%F��fvL3X ����Cu��v�<ƘOnر��knkx�gC61E���Ė��MĪ�Wv-�1�lF��t��n��P��[sZ͇���lkrgc[K\rO=S�wT�1�Ջt�/jb�O��:ԑf�^ЍN����:I��g�����v�q��q�9������-6xӬ\\Y�ޮc��K�r������9��m�L�_�?<� {;�v��n�dY,4�ؠ����lJ��R��twwn�칖��٣[o=�6<�1���B�$��e��� �f� 5�ƨ���c�rZ�vՀx>�E.$CP��.fh��ld�*^k�;��e���f� ���$��@�L�*�L�F��\�;x�.�3�6hA��i�l��}��3YMˮ�kY��[���s�uc�-:2d�[,����O��ۨWjW��72���j�� �f�5��?c�7b�<��.2[��V�͚�����J&&@�D�� "Pΐ���!�滷�~r>~�=y�u��ܘ�Q
b`r�L�3V�_���^F�R�o=캰{6h���^�s�	CsS5�9�s#Hמ˻lG}� ��q:w܊��q�Hf8r8�1���m�������T}@���!�)�s�e2D�qx��-��yW�1�[[�ͨ�ܽ<�f���9���Z�]����~��4��}6�f: =�i����<�Z�	�I4�3*(<Ǵ�;9���٦�f���.!������r�3.ϒ�Z$�+~���P��$��������@y��̆<ɖ��D�neˠ�wwn�=��A���ؠ:_�)�U�� �(���M� �f��}�E����~̻-���O�鼎�9ie��sJ�j���1��^�MmwP�h��7:3]]���:�u�2�IN"g�g��h����;վ˛zٛ�4���q���l!�L�X�c�r�b^f]�wٳ@k��(~ݍ�53a���`o��v=��@M�q@y�9@o��B� �M�&Ss7e6{3g��5ǲ+1�9)����}1��>�������W��,֥�%D'1$LL�_}�@r}����s.���3f�}�_�����x�f#��S8Ѯ��jtq�6!qѸ�4&%������s.bZD�N&z�k�;��]��fl�I.%�P<���l1���`�Q �3������.q��ߦ���v
a��[�)ٓ����B9$� ��&n�=�l�_s"���r��˱ ���T�S���)��T��8�����l)���_��a�\]��ߦ��Sߜ|9p��d��B�݉�Ļ��oz��M F���\��T��\�%@�Ox;�����^;�=�?EJ�q+��Τ��7b��c0�*mcw�׳�# (�5�Bb��(�v�T�7[��_���<�~����m�9�����t�٭�ym���Zk'>�OF�X��1f#j�"�I[֬����J�ɬ�2:�Ln���f^8�eێ���Ә��9��ܡe��Y�b���h8�tp�!h��Gc��L�6
sF{bn�� �]�wn͒p�� _�@ә/���#�]L��Lx<��*R�V:�3t�U�5J�E��Y���楤��St�Jr�ڐjEs߾����͚ Vw2(:�#v(^��
3�L&5(q7`y�͚���̂�̂^v#6sn�������L���̉�fdM6=���ٛ*�9~�^�qp�%T�Xnć[�f]^��SA��I/��n� ��b4�6� �q2�3�ͻ�٠A~ܚ �dH#U�g�{��se�unʴ����5�O<j.Tp�	۵�=�^/^0��<�Y�ڮ��f� wۓ@[�d}��Zp��ۿ]�/��@�D�d�8��@�ɯ�>�9b\�ĸ��.ӎ�o����շbٟM~��|b{�I)�SU67�P��.�K���.�#c^�6>��kC=/�	�"XLBp����w���h�͏l�*o3"PY�H�a�L�q7`��@B�;� ��H��&�/r�cZ��m�1*d���.�wgs�%��gqCr��i�W�F�M;Y���͎�H�0�"fI���A��ڰ݉3��-���S@��k�C�D!8�q36@����~�Z�9�ހg��)��̚�D`�i�9&(��wa^mw�q�[|�U> v��J���%G�HS>��=����*���[�����=�I�A-D�Ն�"7g��p>���͆��ڀ��m�]͆��e��%C�����M�"%����=�4����ui4Sd�������OW�8v�"��ژ6 0lF:�xj@��B�(��L	L����[76$�����͍��}ܚ�DBk&F�I1l�͊V�ٯgb�o}�Bw�D���Vc��(r@�L�pM���P�vh����̉ �}�]�}��.�p��nbb���ۚ��۱(�}�~��G\@��t�k�(c�쭜��}<�����
a	�ӈ��;��s����]���P ��J�}�O}�n��κ-�a�X+e�#�Z��� ���٣	���8.�c�m�x��P""bb�3ۛW��3a�ł�����	�@ޘ�옄��6�fn�͇�-���ɠ�A��]����zT��F��%�"PL��G@w� ��$w�d�[͝) s�-�#H��LD�����܉@w��Z�l���R�١��",R���q11�=��V���m���5��#� �\���uڹ�����Ws33wue������S����WwuUUWwwV]��ū�qp���	"���y��Y"�����l����D�@�S��I���ś)��B��:_��C>Â���
�� Pa�-�fb	�J�	�n�!�{W���6�����a��!%dRNP؁��ϻΖ�w^��������ԩ�����߿J�E��GU�C��B�b�s2�����E\��X�ڪ��������� ����*� UW<�6�5UU�k�u`�v58�Kfq���3rl+۞��m�+������.}��ve�ų���;ms��ss�l!�\d��Z���5�W;X�Շ��g.6�+�kF�����w[A��+c��nl�[>�] g���t�vі�Q�G;�����QÚ���H������0�<O8�Hn4�m�&qZX������&MeS���*sxk�{:g����4�f�J:�2�7��m�X	IQ�$�p�-˻J�0��/��f���l[�kl�
����u%�e�$\v^��W9�F�=;�:���y'B���KN�a͸{<lm��ၬ���ml.��ōc��Gkd���p̦��mtc�>�8*2r������؈˞�~��M�U�)��e�����c�.��Le,�tR,R�-�0�AaD� �۱:�3(p�E�y��&^wlas0؛bNv�SXN���-h&��y�5�JX�L��l�V��cl&J���G�n�l=f�LqaN�����N��tz}4;���&��ȏ`b9�wwZ��e�������gm�;��8-�ڜ���ٱ�r[�m,]���a�m:Υ^$˹�1	��bvh��2����v�jjB��l�jGPAUa��|�wn�8L�FqԶ��X��URs�91!'$�M'VWmUY���3!+�[ \��]�l����X[Z
]�l����"�cX]i3m�,�rd�@�U�]�RZ�mT��v�xj��n�P�MV�]�qv�UW���0�P7cmGr��&m����[=����2���b��!<�N.�؃��,rҩdLp;U���c�pqӑԧ�˓�q�m��@pF�SD��K��n��D��B��X+ T�"�an(��f``� ����]��<�w�=6���06��Z��j�zNYs��L��J,X-�{����)�qǎ��a/�k2U�*�~|/� p*�{9��
"t�B��D�w:�|��AA8�O�� A�Q/�K�Ij\���}��OЭ})��ڟ��uz=o�jK�I��3�1��J�$��PΔ��V��쾷�Un)"IrL���$T48!�Oo��;�~s]K`9�-���dƘ4��;䧜�+0j�)Ś�Wh��4���s�*|8 l��	�f�ifZ\8��Qs��;���|:�Q�p�Z*��mΡ�jy�=���pD�<\c44#%�t�v0��q
��b~��Y�r��禆xp�r]l�u�Cm��χe�s��x8V����m���)��I�{s�<������*�$Ů�7�mî̈́�Uٕ-�4a�R�N�7v��O�k�
�8&d����s��<�ٱ��j���Ϯ�#�}�0ӄL��̔��*��d7j$��Ȼ3gJ�.q4�g�^���
`I�1l�ؐ;��.�Y�Δ��*�����m�K����A�yݻ7gJ Y�y�h=y
@/�32b�$LKc�j�Y�:E03}�Z�n��{=���i�lL��&!��f3'`�����[�J�r��n(�{j2�eR�d�M:����h=�;��E���`7���@Ix��~��4)L���V�72'�8�q$�{|�����S���v~��t����4�DfDC5�P9Nbb)�9vln�76h5�̉)�^^�)""E(j\�"f�A��@�;��`���e؀^F�u�B�n32�&(
y��V�*�W�@w36���lP���r֩��(gS���O��݇B��\�T�ڴ�q��m>3��������ۇɁ|������9����y�����D�?M<��Dkm
\H@DL9(g�뿗8��T@�����7�hfdLLA�Ł�1	�RDč��.���lPo�j��.W).p���h���7����v��b�Ky(&I�"b�37\Јo3"@ﻹv&�f��VB͕	M�5US6�� w�̻fb�T�דA��?W��[tHݛ.B��
j���=z��]�a��V���b�-x�Qu!�04Cj��٭��$�yw�߻f6�fҠ�ɡ �2$��՜�b�˘�"kz�n�R���1��f�7v'�_��]����)6a�P�D�̹�@�f�M̉���Z�33iP����D1�ӈ����oﾉ=��ށ�ϩ]���K�}s�_���2dXҌ��'�0�`��!��H|
ϳ�w�w�����jX4��Jp��f���6� f�M̉���{�`8>	G&�]��TR�홒:��Q]����g���1��9�����9�F�j��m����gc�6rh;���{r�%��V�q<lR�`�beP �ܚ��K���@S����-�ӟ:V�-=���D�)�*�:�636$�3/݈�~ȝt�3s&�/��l�J "Bbf(>��|��m��ߝ�̕@�D�K�ub�s2�D�2�M����s�-�?�&�36$��˰��.L�-��b��D> �ﵯUv1�퍹Ԫ�L��m'�Z���[\��h]FZ!ujEX:�5���"	��]Pr��]���NXkXe��r�-f�W`�O^�Z;VJ͕��e"]J-���֠�!B��
V�v�N��l�\��ݗi������,8�q��NϮn �3ˤ�ۆ�u���n�93׺�q���&��h7frqͺ��n�]��Ipo^�M76�-�::-����j��Yn�9�������3	.ƥ��LC�"LJ�2��,ɠ{ ��ٗ�.�=�:�w�7�b!�8������y��.q�n�w`{c~t��4|����&�9ȗ1@f}�M،~q���.C�̘R��2غ�<�nBDU��k� ^f� fdHW��ګ���b��pӘ&��Ӡ�ɡ326�{��a�vv� ;?{-�oʹl�k�d�3s�V�T����q������ޤN�%�3l���6F�v&�=�ݻh��q[~Ϧ�;�P���% �`r�b�߳�l��~�����=���{���d������Ϣ��l{(��"q.%��þ�-S."@�.e�LU��c~t{��VT)�7v$��˰A�o0f��H��.e�}�$��G�ߦ�>��o=��̜��5�{po]�@�Lq4�&ln�I�\o˻���ݍ��w6h��H�4��if�k����b��66��;8���Pә��h ЃxV )n�h�PC�߳��̌�@����Ć�Z���KS	 �Q,��@�ƭu�8���w��hwb@���x���K[,�dBs��] ��sf���~��\ $r�F�-�/4 ��9ˍj�32�A�F~wl��Yb_)�*��f��Ĉ3��e����ۯE�ml��4�xc
f.f(��ڰdf�Y�҈3�4(l��Db�g�Dˁ�X�8ͭ���X6d�|�yS��W�����O�V�c[�V-�2ʵL�>[/���۠�_t٠̇,;{� �5`�!�C�&%K�t{�ڿ˜樃���H�ٷ`fF|�[ww=s�0��s3`�]��4s3$�H�ܚ3&2`�%��&��mݴ�{�~�Uwߟo|��|l
���irK�H}��~��������]s.n���u������lߛFÔ/���fw�/���"R!�0)"!��6�T��)���C6ɗrt^]��۷��5�2Ԛ�ûm�>{������{{�v�Fk�ZA�l���-�7*��f�̓\�E^f]�=����͚BZ�m<1�3&e�}��ށ܌�H�D�k�k"<��N���H�.M+{#5�{�>��9���s�v�.��i�(jP���13��� 1����؃�b��������(H�,����Bڰ,6E��Bf�Dz��)/Nۛ/tQ��r���(-�Xgyr��3,�*�naq1�v�&��.����&�CS��;DR�O[�)��7�&��ۀ��`�hMj���L��.l&	s���#���Ͱ�V�λB�0�\\2�#[st��E̺ا 8�ֹ慚\6@�B!Mc����V��b�E��%n���ݥ�?''d���/99 	]��j{�΂$���]y�,Z.U����d����{�w�������w0&�Y��<� V{2��y;,��O�h7����D�1�ä{��v�1�5E X�FdЃ��m��ǒ2 㘕����dcؠ�rh��q%�L��� U�v���űT�"""`�s1A�{6j�Z��U:o�������~�k���_B�%�Ji�����5���yvL�͊�ܚ �Ŏf�`%/]%�����0R��KL��m�v��v� !@�j�i�L@(��3�;�wf��1�lm��l�^둌-w�g"&x)�\8���?f�9Ŋ����	"�1���Ā$!�<��qq.8�S���M��9{��`!yXlC�Q2�eLL�C�wf���r��]�3яfhf�c׮��
S"i���u�u�y�n�c�ؤKe�6h�s���j"Z�Là/��v�.(|����5�s>�����NI�}���|����)nQ-�X\.�=�H>9uT,5�S�9��-p�#6�%���t�z��DJ�D�Oְ�g�@�Y�@c*�#.ζr7kA�)�8q0H8����g� f�k� ���V?n�"�:o=��'�K������_��U�e��B�8�W����}UQU35J�""���UUU���yǷ�����d������g�����y�{����N���2�'��k�����ep��$,5&��S\�"�dq�ҌLj�JR�#AFȰ��AT!���33
;��Y&OC@7��)mXa`�0T�'��4�q�#A%��+J%)Z�]���`��,
9�Y�BP���f�̴La#�e�:86R��&�J�mK�.�Pw�5�"`���4�ae(�E�n�6�֎�Q����X9`v0��k\/AT�CanP��5�S;0�fF����-�*ͭ%E����SM��2���]4��Q�v�F,[�s&f��)��ï�]���a���Q�Ӈ5,R�A�D.��0� ��[,�fP(#1,H�� �a�.�}���F�)�����/�W|�=�K�ۨ�:��ס_��
e�{�Uk�F��/�?��'���%��33Yo?Ϥ�0�K��T��˙��?��54Ab-3%���w.׫���(��aD�08pM4�M4Ҕ�L0�	�ه�e�K/W���ˮ�=R�����s3x6�a�l�@�p
���8 @�h 1]����p��4��Y` 0W�r |��Oo�}�����D-H�2�Ҥ���DP,�	��% 9�+���(l�{)�"��K�h���( '}�9��ܞ�ךD�Dw;p���uWr*}^잉�G�i{�K��#��uܵ��(�� ��D'0B�9�t�wwo�a�'b�;�٠1��R�^��DD�&Id���bכQ@8��k�r5�P�s-X���k��q.dnT�D)�b�&�q��,n8�ђ��5�kw����no��>�Q5R�N�o�}>�{m�o�����}��{��ߪ����C���i�L؃}���l;�v�>y�E {ٓ@g��KBh�S0���;�y͊v����~�T�T,��B��$�3j�ƽ� ���t�fy�ky~����H���� @��� ��C �=��f�:���^�����NL	�� w��BO���w&�~͊�N�g6:�k�m'n��ƼH��Ve9P.&X�6�.4LR*�@	tx�u�ĳvp��v��3Vi����=^k�Qy�}s`�?6y{� w[i�Љp9p���ݻ�ˑ�;_E6n}SB������{��[-LD�L���ߺ�\o�H������"=�@����t5a�%�$D�33�;�ͫ^�+�̻����@g�7�>���Dۘ��ocu�^�u��-{�E {36��?s��9�/#�qxR:ē�����>���Ȋ���
*�s�b%� Ƽ6��k*Q��z��0�8;W���<�:5�٤���<C[QF6�&��-8V��y�����Sv�!fl�����Ab.t�طnz��i����s���J�\��fl�jf��PSd̨�d����;��v.5l���\��t��y�$�戺:����� �����S�ӈ{p.��{Y��5��1q��Ywm���I!s�g�Yc�jPm���R�0��4��%�`��1��f���s�On����`at�[�3��	���wwn�X�6) w����.qG�d�������
.	�\�M��>��{�E��1����`	nl=S3)NL�;�٠3J�}�qlG��~����
�����|�|��5)���&j�;��󺦨}��]����͛ ��M ���k�Kr�B�%�T�wf��7~� Ϸf��3%H��z�!J�$C]�t\�&�u�hԽ�<���@ϑڋn��塸�-A(�9s#��f�l��M����"�Y����`C�Z9�T��n��6���������V��:�҄ȹ�H`d�H�@JHh1����SDV4��Fia�88��\$0�-&�&2��$��L��{��7�~���͊ �uf7�\D9aM�ʰ�����̻.�@VFf±��� �1�KGj�1˕A�q.s��L�����5�>� �fM>�:R�:�#fB"�.&�5�ڊ@��ɡ�z��7��v��CB�[<d�iI�%�"�)DŨ�Ǎpm��훃����v�昪���m\��m���^����{��`,y��YB��&!���T]t�����s��g�}V���E nnՀ{[i����6�*���w`c�ء~��i$	+�9K�s��El���ʔ.���-DL�A˕.f�Y��fM3ޕ ���+.�CV$A*�L�s1@�� �s���R���}��V
�~�v��~���Rݴ)�)]U�w=���m/��6����<�������'�9aB&���nƒ{3.�Ǚ�X�C'2h3�2Z8�A!Cq%��f�ވ}��=�ɠ��8H&����aL2�{`c�د6k�ݛ-��In�3.m�9��l�Q�(����&(R�0�6浳v0�A��ʰ��S���	�$�#$�d!!di�ܚ����8��mt�����CR�7UT�́����3.���=�ɠ?s�Yİ����F�eJ�/.���������v�v��[H�òW�<h�o��e-��0w�g�߿]�[��ؠ����}O�y��Z��	&"Ss5`,~�b�=��@w=�����߸��{Pl�À�r�a�HA�B��y{׽f<�ڊ 细�C�N$i��nfl1�L�Y��v?n� �3wvhA��cZi�DrSn$��^����tcc�ɠv0��S�8����d�Y�^I�9������v�W<Z� �Kv��F�5��=/.�G�Yv#:��66u�Pq�%��oT�Nv�lxe筆�͎�uF4ܵ�T�'V���ipNn�c9�����`q:M��(�LE�,޵ɡ��J�9�#M���-���l�12Yt��9����� �ɗ���CC���8Υ����wH�͝����؁�򢮚�l�C-��$�9�3o�N�~:��r�'�,��;t��6�p&[wU�f̫�]R�؃Lk�0D������"u����T�#;O ��˱����91̉�2�32k���H#swn��Fk�lR�HZ��9������i gs2��kN� {ٓ@����r�D��@�qs�\~��퀵��3@��T�0�Z���-LL�e�&�kٹ6�n�cf�ʐ�fU���7i8���q�j9�0�g'������eu��.�
˂�k�sljrʲ��{��n
������k& ��R�����tŽ�\a8DHƢi�UU��nʟ������c}�M*�,(o�۾�M=�m�8���f��n������L}.PD��T�Ͼ��1�lQ��D�}�X}��0	�JnܓD������n��Sy��э��*C"=����eE��`�B\�bZ��bb`�١_^R�=��E�#3bն|�8��ᴃb#s�^���hK�j'�[$V�sR��5��5����Ѷl_��ofkIْ��ة���}��w32��fF|�@^n�Xu���#%��!�U ���vdf��ɣ��L�ֻ�%�!-ʘM����ۙ4~\Mj#���:~���[c��[0�x�6�Fd��ސ�������My_��˰u�k�p�	"eD̺ �,ɠ32T�f�f_�̸M�ֻ �l�Z��'��M7S6�ʐ>�������c~t!�����S�ȉ$ #Ċ�U�:�D\	l ��63��(E0Z����������0'��P��y։q���@f{&z��ʥ z?d�፩��.j�̌�_s�&�wM�weHg�.�q��[��c��s*\�b�{�H�̕ /���`c�ؠ��y�d�r�i�D�X�%Hff*]Ey��m�{S��<�w ��<�]��b��c|��H�5U���`{6c]`�y�4 �zT�~]~oxNl���1N�lt���6E�+��5�a����H!�i�*�=��t�&�o�,��t[ffT�4�J��}�ݻ ^G���S�j&Q3.�fnա��R��dw�wTf�T�/wa�������fKw�*A����qDF���@n��zvYo�>��%���s��n�n�v����P#fE�y�"�ƞ��4�S�bn�_nN���fE��T���e��Ē��q���<�o�Q�����qUT�fjf���UUUUUO;{����N���$'�A!�	ʒ��ȅ��L�D�.�2���foS��/xp*)��nO9I����	�"y�Cv=JS�lߕ�;dl7�����*w걈����p�B�[ϡ�" "S��cmb�C��	��4����8<�l+a%(�hSzq��a�8BҒQ��f;H��J���l�^H>riMT�7.�1�!�T�� �'Ĥ�^d�D�Y`c+��B,)�P��w�`@�f���f&H]/0��%(�I�N@Gò�$w�}��СK}tT��Q���Ӹqr��$B%�*q�e�P:�]�T�����s��u/_�;hy|�����@*���r�Evʀ��j�����UX6�U/=*��UUWT�"�m���UT��L���v@-�p+[����T5B9PW �؍l��v1�|g����G3*k
ڌ��ơ2�!�3�m'N1� ���*`�^�,�wsd�r�scs�n� �˶E�2��TÉ����6��
o.����v급5�m:y���bw�J�K[��m��mҙP����nLr�Fm86��:��L�:Ŗ��R�0F(G1��B�M��f��s{/6�z���c�re�>��x�'.�h�<��v�M1�j��7/�z��Æ&����ԉhZ�������0�Ã�t��aմ�O�5�!���KXC���MY0.ֶ�d��d�6��[�َ�g���4��d�mr[x�5�."SL�:,"t�^���g�k��^;'�LR�Z�p� š/����[Fx�����AS�Zֺ��u�lm���1�qv�
���3�G ;-�̞І��ر6ת�#\��ۭ�7jf��<�D��y�*��6PM1�4�R��<���������ve�Fn�Wu����y�\k�[F�ep�cIT����#m6+p
�g�㷏3�Ȏ�c.����4�{<�#�]���N�e�:�z�&éc�hϴP�.0�9 3�w2�V#'��od�ʀlU��ک{c�8vm6��ؠf#j�m��!�����b�V�P8d���l_ub圦�\v����d;��b��,���6@9��S��9��͎.׌���gN4Y^��6c��B�tӳ/sSkn=����a�z�Tݷvm'u����{c�X(��p�1=�漛k%z�֛`:�H�N�]c6�=��,˱΁%6�@�7��9������\g�����K<�0{r�S�T⪭��i�!�[[����� l��HZ3mC][�w!�ͰkX�.	ʚ�vy�K<��,�n^���[����[���*ST/jhS��Ν�Tr�l�G�Sн�ҟ��􃀨�C@�E��|N�0"!�"7�/9��	����!K������~��:ʢb�R*A6Wl7��^�p�Y��	����ӝ�V��9sUql��Q˰M��y:��5�A�b�v�n��[l��Q�]|J���	�u��ތ��k9�w�7�1��ɲ��<���i�l�ghC#k��z��l6PR���������w[�l5�S��<[F�x�Μ�S��b�K%�2�u^YJ��7��,j�F�4x��59C�6�su�n��@-fwp���M\J�a��ay�|��B��4�v�������pY�exص��h
�6tLbQt��$K���pK��lT�sg:��b�r(A��T���d]�������-����)@���:�ݥM���f݈3rt�1�sf�ce�X�3d�6C*����vCk^�ҏ�J���c��=��e�O?��a����M��ۗH=�3%H#s�˰�j�aʎD�&B&J ��&���\Idf:��m�#�ݥI�}��|�$M�`;i	�y�F��Y�ٮ�@b�.��Q��C^� \�-��:n!L1���6�� fw�v}���$��1��4Cw��e�)��ksr�_���~�ć�J���U�6>�[6�3"���3�y����<��ზLGV��J���8��
c�7}�y�H4�{B��fT92R{�E a��m�o�{�Ʌ���8�ëзe��6�qQU�Z�Z�G���oz����}�E���{K��?<`��J�Di��k�`�۠55��)�]�R[V\[
Z@[�<��ô�o�]�3#u����?...wK���������݈a�l'�P��Ҁ0�(d?;��e�� ���T�9R�!(���_��j�Ƴ�Oj�otT�W~���W���'�:��Wg[�tU�þ��V��p�$Ұ�qq..?�u��nm}քll�@{�8P�Ld�!��LCM�&������l�@��t Ǟd���k�٣*�L����p����n��K�W�� c'�)���;'X��V6�6t����Ǟr����	n4dkR�`���L���c���U�#{�D#��˰}���;	a
!n�	���U;�ᄁ���]�3cu�6�v7 {�@d)!2�tq�����}�l=��j�~��w�8��J����� �އ�TB�s#!L�fj�ϣu�ݏk�1��Q�N�?{��~������-�ŀB熷YK �Pո���uvȼ����������a/|�3*D�&e�p�FcT�<��m��e�65k�{���l2!L"!�
�wM���y�e�!f��=���M7���������M�Lã[�nj�f�룭��:�l1�9@j�lݔ>C���m8��63]���k�5�����>��լ7e���&e7D�H�{]��G�% �}�۱u��N��.O�~��l��C14���Vxyn5�챚Ld��>����s`k������+�vL�Mۿ�_p/�V7Sͩx��ۜ8Vlf����;A�۪@r��ѳm�NӮ`B&�zۅ2bM�[�R����+̖/+ѵ�T���\V�%{7�A��O:�08۶�`;+�֜]�0��e��.v"� �s��[���ܹ�W7\�I�Hxl�>�w���n6j�X��f�И�V]CL�]6j���߻:k�M�)7��<�-U��jY׻��~�,+;�.�����zr��Cy��@=��Kn&�P��v���k�;����"����؃�۰�S�6LK���F���=��6w�����<���$��IA�fV2�|؏fE�A��v��Ӛ����܅�;���$��2n���k�G{��_%��o2M5�AI,s0��U�ma-�sd�t",���N��6仉����T�C@�L4��(�}����t�f��8��{6h|���6(���271^��Ǐi��\@��B,`�1 �IPC. `�I�aJC))
D�5{���	�A';?uގ;4Ps�+����r� �j�q1e�%�pV�'J �}~�~�}v�|�wX�͔K���U
�׋6*"�����n����*l���(P�Aƥ�2DQ��d�Ձ��v���Fk�͏����,S
[p[�qy��,��6ˮF�>=8��Z|띌2[v�Vz�1ȑ��Q_<���~��m����@#�������������NPL(s.��Fk�m�rbA��w��n� �����dDDHT˰fD�g^y�]ul�{���00A�p�.����盔�Q��fu�޾���r��c1���2T!�P塑3B8_������Ҁ�zs]��Oّ g���KdKQ0ۘ��sgJ���v�ȐW�>{�[~�S�f'���,�i5�]-v۝�'eA�:�L݁�tm#��l�>Nr�9���`��{m�=߿n��ϿF��=���v+]�bzd-DLH��U; ��&�|���{�(�J���B��q�M���H��݁��Ҁ�l� _}�E���1-Jjdq3V �\\��'a�͝(������" yȊ�(	��[u�/�9`�g1�$��jb\�%tLl�B����w�v^ܝ(�Z�L?���c>�^��'��>μ�š�lA��	�s8D�$w)�~I9�c�u㡳�v|�G�"QM�g�]�;�:~\Vû�R�;����0�sq�LLQ��ϮЁwrt�[�fҠ�"W8��*�D�6�"mXܝ(�ͥ@"�� W{���>Mm���3�������I���j�;�So���b*>̭)K`����B�D̂q4�s6k[3�m���O2t�c����Ա��](���]ش�ōeCSu����[v,�܂੬:�<a�\u9,�<��e�Mڛ�ق� $�\���M��ع�۱P�؄�2#��z���t���|�-��/b�ҡP�DM���xr�2�6�z�&t������n�q�ԙ�;yy�xVv`v��Eس�;��2>���6�b.����,�KmT�M\�c�.�hO	#$��t�n�P�.�6�.(�vv@��@�B�X8�񼡚�e����,9��BYq��8��m�����������:V=�FV՟�\�v�ؐ.��j��$%�3vٓ�y:���:����C�w�����%B��}2�\
&%�P�ߝ _}kR(�{>�b��PŸc�l(nX�!������"@�{�v�Fk��n��W�י��"\�qSh�_�`.o�u�#��� w��V��A�!�@
H!ȵI�05�q�i�c��Wn&J��͊�$��P�;VsEv�?>Yo�O߷o������ќ����｛v4Z�F�	�r�&e�K����W��Z$�� 8 �*�""&�@�A D��� �T��Ax��%go�Y߮���Fy�k�6	{Y��r��1"�.���3�]�c�:썘�t���T����8��q1��\�\\���]�����]ly�J�;�D�-_�����a<q �f��n�w7k����%���۵�z�o��:n�GZ�3.ݷq��N6c��c�hD�%`��J]
lk��4goZ�I�c���=��/[���DJ��}v�7]b�Ƶ�ja���X7���+��]����c���Q�s�g�J�R�.`�8q2���n�ݍ�E)_��>�TC�����EUUU:�����WuUUUUUWj����˻_9� %�&��r�ʩJ*���<~?�0x8�9C��0`�l6#4�+�0?s�����o��k[�����C� �Tt�tc1����T=n[]�xt�6gu<!Ë��C�XxQMK8X6ĦE"���$H( �"hxذb��RX����J{�=�1���fQ�̊�rpG@�p��Q��航Jh8�,Jr��M��������L��I2M$/]�f�{Я�C��.�w�M�3���f^r� �h ��M��z+�@"�/��`��b������P� `�_}ġ$��8����=��{�>��zW����G8������>�����wI�{�t�(P�\�3-�����Z�g];�͵`�D��]�e��4�Y052�8��1.���T?{"�｛|���#u���b"Ħ��,����p�V�f���%��#c��1�qF����l���N�\��Bs��樱�dH��]��Ѻ�ˢٷJ��炎F$J��DPnc���@܍�D��ݥ@#��L�Z�?=S1�x�G7`nFk��nң��>��6�̺�l�����rB��c�t�r�S��H��n��.{���R�ZƜ/�h���6E��~��Ҡ>^�x/����pB�����P}o�v ]�إ@wwiP�=�6����cr"lڃ�v#�*��0��U6㆗�nJ嫜ϝ�Y�@!M���w26��3rgJB�Α _}��#!�B��Q3-����7�:W��s�⨃۳�B~�D�+�}���s�\nY������E\L+����������_}\B��{�v�3^�%�=�P�b\4�%�Qa��s�{w>�l;����K�r;�_L5��G#R%CN&e�R��>�)��8�߶���7>�T!{﹪��BN�P$��ϻ�/ص~�]N�W`Sg;e˚ʠ��sAug]vޝZ���ӳ����1�WL�R�|�c��H�|�B���9li�Ġ�v�Ò�u"���뀶#��ǔ�b���%t��b�8�wA;]��v�tlu��K��f8l��{��1E��Ulp�p�6�܆����U�c��J�i���!ܦe�bbP-��\j�J�啎5�����f����x�Bw�w�5�;Xc�v��Y�Kmu�m���CJ¶ jAa��Gh�{޲س][IM�,�K؀��2�}��F~t��Ҁ/��K���/s6�A3H+�]�m����P�Ͽ}{B��۱�Fk������֡��B��- ��č�_��h!�mP#sӦ�<�fP&\�	�LLP��b>���Ym���P���%���!�O�n��$j&aD̶�.{~�����T�J �}��۰5`�b��1(�S����%Ni�Uk2mh�����qV�܋x%�C�#�UD&�P�L�s%�~��B��M�c۱s�K�����@��}B��7-i[��꯾�����}�d\Pa�r{۰Fl<ؠ<�� ���BY"%�L˅�3n�=�u��Nk�nD�����b�K�bP�n����;�Nlܘ�R���� ��IsI"j"ee�#���(}�E o{�V�7]�(3�bؑ9��,�7M5�*�0���-F�3sqZ;i�p��' �T�R�pD�T��ُ2#i�w3n��u�#����`�y2�511	Ǧ���������}<��}���n�4P{蕩&���fF�G$�6�&iu���}knj������KU;٭��D�����zLLH��˰��$ʙ�P8��1.��Ē�Ͼ��g��pS��y�{gJ@	i�B�9��!4ɉ���fD���n��al�ùl����a���:X��J�.T�#R��r�ӽ�U�[;mƅ�Ա3���5�����(��Y�w�Qss������bu��NL�� �wډ&&	���3V�n�_.q�ﲴ���/���w2�x�a�o��@]4�eݿ�����^�&��߆������#폾{l<�A赨a0�Q$\�s��Flā���]��F�Po8�B�2�#]wwy��zv�����bsi�����=��LLDBq3�۷`nF�7��� w������Me�}�;.j�E6���ϳ�էl-"lyu�,��X�8,�3�:\�6�&n��l�v�lFc���%���� =�s�D�8���J<��2�Sa��$
��]�7�:M;%�diP�"a�P��U; Y���7۷gˉ	3s_Ԩ�v�,��j#by0���.b(<�rv�1�rt�a���A�I�{"P^�G���	�j%]���uѭ��N�;�D���e�y��s�r�'?3Nv�p�U��5ʂY�/0���K왆w7"k���q���KÉW��0���n�u��3r�;���W��ԍ���x�)b���[��O6��ǖ#s���;(��\ˢ�*��)x��pYp�T�'��\W(ն��t�t�M�\k�Ib�:l���V��\.n��׬�A<��snX0n}�|��e�n3���3l�0���4/-7�D�1��y�L�[Sw����w*�P:���7��}�ҟ{l��N��<�	�i�a±������8�E3nD�[~������}�6߻����s�E��� ����f�(NQ1J��ȟ��D�ͻ�G�:-�}�����}ޱ��+@&O�in��.�[�����3((��H#o�!㘈93ډ���[ZP7���T /=���v�1��bSN&e������J��{� w�{.���Ҁ�����g��{{�oX:��.��8�y���\3��n�f<m���ηd1�waV���ѓJ����ؠ=��v�N����)PC������D9nI�����ߔq.�J��$�/������@gwiQm�����I�����H���<nX�n��6~(o�� _}����f̹"[��A1%�7�J��� ��U�˕�/�lK{����)m-� �lH�g���̝(��J��s���g���ά��� �,L-���1{q����ִgZ� 2�lFLe/�7��7	Ӧ	Hs1`n����N���)u{����ߵ����^)��+���OjM��w֨�ؐ;���ᵲ�y��L��Nfe�K���J�l�dJ1$�R��$1Ur���U��$^�u���3��IU۰=��t ��[Q*!	�"iXKO=� Vg����k��v�<��Ul�M�CD�8	�1���v��qqO�V�� Ϸ)V6���]<�'�í��s�A�靖�Cf��K<�۞	�8��J�Z�:�l˖�M3h�yW[ݍ�@�o�� /w� ��{.�����`d�j"d�t��a@�P��]����I%q�߁��G%7
fY1J�F/��5�n�ݑ=����+�s��ajbG���n���k�3��('�$�BW�R�U�+C�\Hά�s8ɘs�q.쁞�gJَp�l/�D���e��B�5�8F��$Ĥ���4�%,xcmq�d��1q��n�{
����[�SE�E�����'
܉s���$��)��	ms�l/�j"\L4ș�,͉��wٷrث�m|^�"=�ʎ��u��KD�rۙ��w3n�ܝ(;�gm���`�o|�>���$b�W�[~�n��fҠ�"x�}�`���S02Q.��)�̥@�P��gz�gJ��?{_��UUUUDDT���Q3;UTT�MUUUUڻ������������������H�*b����bY�'3"\Le��*"�)r�0U&�7��r��<�?K����Gɓ2�0�j�s}���C����bo7c��64����;���""��HցӃҕ{þ��A�Ȃ�����6L |�]g$`�?}߬ͱ.Wvlp�s[ɽ�A�h��"�s0-.�jz{o[�bZ�����'�t�;;���D�w=����	�ɗ<w8��=�p!��s����J0@w�}��Y�"�=��;��M�h��t�:2qy��N��;0��C��cx�Oz�z4O�	��=�=N~=���D|�����tn��%8Y�ﴙ��������S��~��;�d)A��I&l
WW�\;�tZ5D��f0�O����-?N�x"R�%!$%���R��tAh����}��b'��w��O�ĉ���5�YB�n2���E���ͧ
5Q_�����<�P�)���{�7v�����nR?v;�;�c�\�mUUZ��l�$"�����k�UU`Lꪄnj�UWT� tv�f&ق�h`n�n���<��֠
�Neհ�Zڬ�2���M�N���u�B��g�WO$P�ˬ�^3;,h�)���$y����Zq��z�q��袅��\˴�X.!)��6�,-�����(٨�b33 �gv�v�`��ڂZ�-Y�۳4Q�Jg�������!��5�չ�.��5�U�]Rٱj�"��KGj"1�����]��w�6�`�ݱ���%��.��G�'.ݙ�ٚ�h&�ҁ��Tf�������;�+�A�����A�t��T@�Yܤ:�Ӯ���cod4�1�4"��d@���Nr�k]F �'l)�F�����:�5��%�I����R�Q�.�@tH&ē�alm�e)�y�VqS��<��[������z���^�V+�����M�����w:���v��D�5N&���Z�sahC�Nf7(�:�GZβ����������u�{�@͒PP�x2l���Ҩ���Z�؍s�x�LC����[���=��u�͌�jz�k�6�vT���8����2޳z���"�N�q�6�P��j�uf�'��Rs�3ۤ�,8�$��"D�L;Mg0��($43��z�j���q�@��U�C��ݺ�컗K@�<9\#���6����ؠ���MK���*�
�˭����7ɞ�P��� 	���H�Y��su��:�Q-p�U��&Ȥ�,�$-�����-vz�sr�ڞcV�]Ρ�ӥ&8����D\ܦ;х��2�= D�����ݤ�{����:�8y�r�ץ��k�ɻ��\]2f�]��|�yya��4�&VԚY���[.��d��� ����K�6�T�̒�:��.3Y��%D(`[�E�j���Bv]����me�T����*M2*�el�4��1r�je�n�����O��,�t	'd!�*	\�ت.��e@�W��N"8�:�L�U9�v֧<{����hqlW+���؃�.bV�������9�WiˆƝ�m�K�^���՚��]aQ����n�/|f��3n�Sq�bŏ��m�G�[��kv�+9��`�QҦ�o��T��~c�˒�{E��K���>�K�g�7��~c|�IZb�x
F�ӉՓd����'ݍ<����3�<�ڧ�yv7
��M�`[���8�H�8�%�7Qu����wZ,q��G��R�r��;8��g9m�IА�/7m��̫�7c�w�W^�ܛ����FB-իv�wG�#��;\tɡ�D)D���d�x?���w=��a�3�1�g�2Uy�y0���&�����ۻl���@g�iPs�>�̛��:�r	�Q37bܝ(w2�@�D���e؆ޜ74jbfbbT��32m��n�(ۑ>l�O��nΔ�fd-���r�&LM+ �Ȑ+�]��������)P�(* ���i��V�p��i���m췽f1��g��iT�8�4-�P�8d�ԴJ�D�@�>߮����@{�2�@#��_}�&bf�T�M�ۻJ�9䗹����>��|�O�!z����D�fJ �ȐF^{�?I'9$��������A]E�����}����6�7c�����B����a�~�?}1 v���2~;l�q(����	~ݧ	�Bn�U6���l������}#�72u���LH����y/� &�8�1\���CKp�s,H�6/CB��[�Cp�\We˄�C�9���;�:R<^�҂����qS���u�τ}?G$�12@�J@ovp���q}��ALJo۰;��:_q$�$��_���.T���]���H��]��n>����W8d����}S7m��r��2<�,m��(R�I3[}ŵ�`w#u��Mﾝy������}?�R՗X��YN�f�{�,3� ��U��P�9i��%�����I^ލ�x�T�#��g�Շ�I�[�R�bɎ%j�
�.���{8��d�*k͢�}��X� �7樆���I��(d8�
�� �Ȑ/�����k{�t�3�K����̧�P�b��sn�^͝+�ǜfFӠ��Rw���"\'	��9�����~�� =�?K��D�s�vx�L�F�P�;����k9��U��7�-�&Y2J��&H�V6>����%����Y�;�^Ҥ
_Ӽ��z�Q,r�Yq��m�;Em�A�љ��)]�Z�f��Ý��:X�⢜�-NT�d�S����aH �2���Tv7��R�dB��j˘�ssn��f��J���um���e.�sϿO�A.����l�fҠ3���l��@_��v��ㅰL�(Q3*&eRgcq�fD�~���u���tt�{5Ñ�q2۸�`#w"@��s-X�7]���B�8��葓�=��r~�nfT�~w6��k�������3�m�x-b.�yۛ��9;m�e{�s�w=S�q�����"���j{-NI��[�$����J\p��gu�G�t���z��%i�v��:��V�`�vGq��Y�A��]�v9��rA�[����()��E���-RZ6�-A�I�ox��ӹ�j��;����/m�`uv
�i2t+\����$��Ʉ��$�t��W�5�ιn�;)q��4`���;�WKL	��IqKU�� cy�zsո�;�� O���g�����￟ףl��iGZffD���ő�˄�L' �D�lA�ͦe�Il�'>�)��S�.�s��>4z��"	�D̹q*���=��M����v7�}J���xj"b	!��5SQa�� w=�,�Ts�q=���+�֩|26&��MQ3�͍ݻٛJ���t�Ȑ.�C<o	����C��"	cu׭ۛ��a�WɌ{.��'&�ek���2I����lY:Q��Ѵ�g�%w�r�!��o!F�e�9ls3PYQ�oﳝ��}�{��;S�$0a��|�obA��+:��7] �^��r8��*[u��h�ؐ;�ݻ���qd�6}n�����Tد�$d�&!��=�}��3Ѻ��n����H~g�HN$P�dD�ݦ��n���q������ĀZ�~ʳ���i��R$y�Ff74k���eĎ%5�q�1����C���[��օV�A5��t
�ݭ,��T��;��:�r7�@]>k��&L��ɚ��76&��w2����P�3�:VT(#�jQ�DĎ852�Rٛ�`wњ����Ǥ���pH=B`�X�V��Eח�Aڈe����W*+܉���� s.\C�1v�d�@gvt��̚�9�23��ź����܄����Ĕ�wcJ�{"��۷g�̙Ҁ3���Q!�3 �e�z�]qEF�t�v+l�qRb(u�F�v���:�p}�C��8dL��S� 7v$����R�3#5��%;�G������d�!D("&h�ۿ���c~t�>��fD�D#�f�"H��dD݈;���
�N�V/=�ۗh�X�fG̒�̎&] �%�%Ǜ?k����]z�^u�ZEr�� Ԇ�G �C�@$�}����Y�����a�ۄL��	��`���f]��#u���tKj���RJ��.dS�p[� 4�m���tq$�7�/1�ݫ�Og��v6��G8�P�)�1�a�f��27]=���03=S}��#x9�Ø���`fFk�G�7��D�/�ܻ��^�T�}"	_Kq1��S1*���� ��H��eŰ�f�t��5�4�A����H�"���[ܘ�A�g��ao=�j��qqqG�콧@{v\d㙗D8��=�ٷ`{3iP#v=����dHࣹ�����P&$N��-�S���0L̸�D�L ۦat�ڨ(mh!�n^�M������Q�n�c�9=���8�ky���{qÑ�g�8����c��9�F�7 �
vgj���»Hm�erѵ��V֧���ӻm���ǚ̺m&6ҁP5�k:U�����޸�Ӷ����r�{��m����X�5���uq�vɉfT��np�p0>s���"ݸN�X�
�*G ��c�\���[�o)�@>t��8ݙ�Ƽ�"��qDL2 ��9B���f�����@�G�P#3�ۿwfO�(�dq129��2�l;���BfD�=��]�~��T9�Zƙ��73	�4S�݉��e��ٓ����Ck�r(�$�RL���y���H��N�c{��7��(w��˕��3.&�A��jJ�g%��� �l{�-�s��}���F��\%� J�ͮH�˶x�2a+�*M�z������ ��#s3
N�5����!O���r�}�G[����S���̻���$��~�����3����WϾ���ٻ��MY�<�c�H��&!�W �����d�H��t#�1���͙��S09�Q$�Ո=�:P���`{2'���/�j7Wj�o�Ū>�"f	���d�U6^�c�3�L=�wbfN��%�e����G \�%Ir��:��i��č��\���a[�����l����qQRq*"Z��MM5���H#��e�̟���8}�}�>��
&$p�9&"���۸�D̝9H�Վi�=��F������˘�(��6�ݩ)�nǱ�~����QUUUUD(������uU뻻�UQUUUUwe����oxT��T2՗�v�ք^%��\lU���̮M���(�`��NZ��Hq��7?�&3�d����)a���-'F�H���d�G� ����G,�'R�tv=�s���6թ�D�yɴ0=��w�3%a.�]�R�N'@5���F(.a�v���7-b�UbJֵ�p��R���`�C��z �P�(IE�V2"���%�`���y��J�y������B���&�V>;|,�4S��32<<��Ґ���[YxIH{ޯ#�Ḏbm�����J�=���5,6<җg��Ѹ��r�q�'9�8&	PD��^ONp�*�tif����E��楱�H����o6@�&D�a��e��Xu��^̄ P���Pbj�"�,�&ZK�0q�Ϗ�s;ϫ�{�$!�'�l�����!�P<����� ��v�i��S��:Gi�A{��y rz���5�qy����'7�[�����q&��IU�FĖ�7cn�^�9ZۉpL1��LIH??���@��y|��5.}��j��~^��5.Zss.";��ؔ��)/fn��{�O|��g��m3�Ĺ#u�赚�f�[����1�1^gy�[]Y�.�0�m��I��b�fn�]��in����<��l�>�,�S
r�D�qUp*����k�>E{2��~ܡsV(ٙa22�TLMsu�5e�2WL�ݮw�ݮ,:�9F�.�55�׿}��<��=��q��X%��$�A���g|(����	����wSO�%�DAf��mq�x���e�g�����t�k�t��:�[@��Q&�j�j��v}WS�t��ֻ(��(�@e�!��?���}Yh�F��f|��,����//���M��i��LM#7Ӈ�qqE���ݕ���^ �{6����V�g��|ژR�D��C�8��}+=��\���=��t�o����"&"b����~�yf}�/o�W�%w|ײd� �D��D��]��izm�{;�]���r}���'�}�aR,r��4��=�H�P���in��Y����<�v.���+�=�,ڍ̎�]cM�C������.㍧��]OYS�����qn��wY�&6�� &��L�RŦ2I�t��]�r�m8P�v�O����|��p�y9�ڻn,ع��#JWR�i�.
jk��������Nn�9��1��rp���ٓ�Q�
��ImmO;:�\�7R�n� �I��N
��d��.�����#��b�[��:�7�S�c\Nr��.9KrVXAWWU�,���}��|��ٕ�g��]�ͥ�gv6=DL�������rcZ�n�(3�ݦf�ן��q��OcOE[��3.-x�o�\��ݬ�q�_L�����F�f[��7.ff���i�\�{�E��2k���k��/aǛ�C��̸�u���|��z�{ە��fҞ~����iav�q�P$$,��ae"k�ƚ����æ�Ė6�Ժ�t`�R����nJ}�f_/s6�k�99���P��]�f�np���~���v�$I@A���F) ��Gz9��"{�^�F	Wsҧ�Ͻ�6d�"$%
&'��~��mc�N��DJ�粒�ׁ2L��J��DD���0�/��]��R�������� �D��#PL�	wے���NU�ۻ�I�nL�...�a�
6Dܑu��m5F^^�������8u��`�f��4`sK�VhK6�]J�:~��4�T�Z����E����'��ӕ�����Ѽq$�@�H���s������Ɨ{����r�����o Ȑ-�y�o�����߾o��PЫ+���GL���}���{�-�$*S�̷�v���^�s+�7wk�ַ3�~�	�̃���q1\�͍�~���}����ϟ;��s>y��8c�4*b +2�h]X% �:�1�Cm�3.�og����U!��"bix���/k�|��xɢ���v������&F�%LL""k�׸��秇{���wwj�G�p�5�L�Z�ji�=�r�~̥��������=���CR�9&b����y�<��ft筻͍��BfA������ �I!9:?{�ݝ�f~ĉ&a��e�������'�n�/{rW}߲����Y��o~b&b�8A�$�@��Վ�Z���1�Y���ŚcPE8��m>w�^�%'�D���7��F������_$����E�Ϗ�)�QJ�Sӊ�fl��w2���v�o�O���1�O�eK���q1KtϾ�wwv�5�4�����E�"5\�P�i}��#�}��I;�}����]����^l�28��0�K;�����w������z ���bL�JD�Q����WٕE�{2���� ���c�1ٞ�4at��Vm�UmUaj�D1�Y�;����Y�Tq�jl�\�p�3(7���V��,)X��`��.�<X�ܝ��k]�-ҹ�#q0�Jڦ�6S�	f ��^ɢ�l/vCJ�:��u̝;v8�gv�p�jM����	�1��`�&ʇs������[:V���T>���������$�$�� ݶ�8f��tS8�'vf�k�g�Mbm)�n]1��;a����m���N���b��L'z��>}��e�}�\���s5�:g�8�P�&���T{ٻ\�wwi{^��{ܞv�荂	r�q$DMr�wk�f�k�히������5L�&D8�3.�
^��X_�2��nW}�ݥ����TL��2���s�����/der�۵�k�j��-K0i���CË����q�#:ũQgWl)=�:&.˯��鉶f�c72�1�3������矽���=���������fH�Q&A3�=k��O��{`E��6�-��%�4Fb����*����~��]��*���_pZ��ꏦI�ډR�8�X�kR,��O=��������/s(��J�%1�54�]ܙ]�)/nn�7�3�fG�&�D�/{3J������`�Y�?J�����1�\�0@KiGnV�8cX�om�c�M1H.X%�I�-%6��q*[I�u��������t��J�}�Iy{�Ǫ[��Mĸ����²aw�R�w)f��.�g59�Q
eCS2ɪ��g�y�=�RS���b"y�w���v����3�~�)���8!��LR����w7b�����ۻ1���"ImJ��Ss5��vѻ ���d��nW>I.}Ͽ��6����y�-bT�6�5���҆lj�se�ݓl3))�e���*�f�b$4M���؎^{ҽ������q_�(�LJ�pL:���ɡ_W��E��ي�_���q!w�n�"E�&&��߯�K�;��60��>=�J���\8���\�M%��[Ksc{��K���.BIn4s�L���HH�D���kV�%H� ��)(@�
 �"����@��!�V�f�Dv�j��=R�.bT��sKq�4����矵e]5�ͺ_.q{��ϓ�E��n(�i�9]OQl׭9]���hgb)�LK�X	,6�k�{�~�{�������wۿ%6����ws\d�fa�&%�sُ��۵ʼ�Ƥ���g�=��I�K��	s4��۴�66Z��z������}��Xb�la�����������W}ﲕ��7k���p�H�̶�SO��d�ߗ3w６a�ҽ�<��o���\�k�AQ]�`
 ��?���ٰ)�n7���R�i)Z Y(@�X��Zj	�R�JT(�%-ҬJ  R�r�P��ZTh\� r� �Z�ii �J�ZZJE((A��@biPV�%��JQ�D�Q(@
ZF�J�(@��JA�JP�V�Z�Y(
� ��
 (��B�fP���H���J�V�ZJ@(�D�)P�J �B��H% % Ћ@%2(�*��B�J�R4�HR�ĨBP�%
P��J������� P$J�҃H��L"�*�%R�S@�4��
҅B�BL*Ш�*3 �- D��R
�
��@�%"��	��(�j�TB���(Q(
$�Q�D�@Z(ThAhF�
�P*��$�D���AU)(��)hP�R`Q
i�A��R�(�P�@�f�� R��%#@�L�)B��)@ĭ!H�M*	�@54��LKHR(��� �P�EH�HR�JPJ"R��@"�E�%R�" hZ�����V�b�F�)b"R����	��Z"P(����(i)�d&�)��
V����`���B���(�bD�
D��J�)b���!���B��V�I�)R��iB�)��
U���B i�Z@�hbV� H�
��
R�
BX�B���)� ��F���)h�ZU �h �&��%Z@�
�(B9�д�E�4!IJ
D�JD�D	J% (�%5J"�1M

�4+H��D�RTHP��-� $�#A$	@�B$�4
̀�9�D��PJ��(ҥ�CL�Q�%
0@�A%�ABP�T,0�J��	@4P�M�(P� �I+J��#LJ	C� L�$д5B�2� �%U �)0E�R�0L�" 4P�ȭ 4�� L��	0%"P� ��HES� �"D)B#@�/'���8��T D�@P���7�?�������S�A=}�� ���y�?�T�@?�A�@?��ECc� "���"����PO�������$C������" ���}ǳ�p

����~�����󢂢����
 �
�r�?��y�����Ԉ���>'��������Y%� �T %ah(*+�~z�_�9������n��������7
AQ~a�_G�o�)�(1*1 *�@��C #
��
@,(�
 R�% � �J�
ʉ"��������"�� � ��ʉ0
@ʉ,��(����
J$��J�"��� J�+ ��),���
J@))*$@)"$��J�!
$2�JH)@��L� ��)! � ����� ��H) $�(B�

$*�
� ���"��*$�*$ @) @)"@)@)#
$,��������0
C ��J�
J�

@� �0
J J�B�(� ����0(�������	*�!�
@B"HJ H@ �B!�����@HBBB*HB�$!!	!,���HJ@I	�!)) �B	 $� �!$"B@��HBI!)!)		(HH��$!	!)	(H@$#)�)
� �@BH"�",�* �@��! 2
�$��$�2(��	(�,�)!"HJ�@$		 �H����	(���BB$�"H@�$�J@ H@�$
BH����!	! �@�(�J���H� �"���BK		�BR�BP$�%"ДH���B�!!J���"}�� m*� �)J0�$���*(+)"�
ҋ$�J��,�"²´�� 4�0J�(��H�� ;}���~_����[����p|+�ӓ��xh�����
���۶�?�׿���i�>��}A��L7��AAQ_����X=���9��>B�����

��a�=}~�Q_��}�¨*+�q����v�����q�� �7 ���3��C\����'A�(*+����������TZM=m��9 ���;"���ϸ��$��x)���l_O�������I���_y�\��������|�<����(������������PTW�O��� ����ﾑAQ]���|x?��������V��1AY&SY�Eh�c9ـpP��3'� a�?��݅ >��	%鼘(���h� �4(�k� 	 ��z��Ԡ
Li�@=ut�� 4� -a@:  t (iY4d���a�D�@��5�m� (:�4 Q�� @]��h�     l  ��E�s� ����>�}�ã�{�Z�.�v�6�ys ����x)�ټ}���   ��97��;�C�������{�������r6�Ϧ��{� w}����Z��O@ �]��@����x�Ԡ���J{��AOA{۔�<� �� /$��^�4�=�p 6�zΞ�=� =��c�� <�} �)�c�   6
PO����^ =��Jww t�{� wqJPzSs��; t��  ��)�yg��0>�{` |�@�k�h:�n�j=�����9��{����S6�6���>����{S���w�D�C   C�3k�}�O�g�-�� y������<���� �g�>�q�����Z|P  � _0hź=����6C�� ݀l�^��{��!�����QЍ�@��}��0� �_;:���|����]�O;���l}>�������� � ��E�����`4y�=�f���#C�4�X`�O��vfG�����ޫ�3���(oX|  }�*�<�=Us�����U{�����ö�m#����>
���*�6|��{�C�r��zx    O�iM�)J� hتR�o)  4̩Jf���� �S�j��ԪS@�OѪSM%J�40����)�@G�z����?�����I��g��}��������w���
��T��
��* *��U����~�����C��`MCv�)�nh�嚷�����ofY��a ƄX@�e|�ə���%�K��8k1.�u��곷O�������ʒa�.�!���ya@��Zw�Gz�.�.Cf`Z�n�����e���	˧˽��R�7CK��;�/	|�Z@�S��^�!L)	���	�����8sϦ}�k][�r����>����y1ҙ���9����s��%�1�t��i��\<��;2W# @��Ђ�Ɩa	�%�H�$("�3Y��{�wq�.�C-��L��o�c�����oM X3&�B������\���C�fNFLpޚo��S���Z�[J�%m��)�n�Y��K�dܠI�.B[2�J�����.f�pҐv7����F$����J�n��՞\<�6R��,!�o5f������O<;�:����ӑ������%��0me)�3W8GɆ�$aYHB�v��7~��D�7O� �Շ�xl��p4�0�$�a�)��F�������ٽ,hF�5s�vg�C��vM���o��8�1!@�e0��D��f�Nf�˜��� �V!bG	 ����=y�ݜ����x� ��K�*J��M��O7�O>%�H$���z�	�{��f�f�v2��#�{�(��{�u~F�뺖���5�2:SF̈́)�"BS@���`�R}�H��cтF��L��}���E�A�	�LP��0(��bS>=�)-���IB!I]�I~��ѭflI�����	;�,�7K���hﲾy{		���)#!F��5
f�Ɨ4ޞO��y��5�xL/�I��{zv���,xM��s�� Ö�!�`K%�!�P2��0ѦJ۰��6y�(swZ���B�)!���h�5�u�; �*�J%�W[��6��$M�����`Cs����﷤���Y��}%�	t��w�;�O>��h��%2�$cRJ#(K�'%��g��x���[�\�����F�y�rY!$+|��>n�吻d_d����N��˽���>�����z�� U�X%!X�do1�-��7w��<䝰і�X,�S�����2҅�Y�6�����bep��w~�%=�P�j�֌[����wĿ>O��K�~��'�^��ݪ8r��^n��]	��n����e����9F���������=�+����JD��܏��|�^���Bd�ѐ	fѤ�>i�a.���v��>H`i	O	��H��'�'��Z�/��]�aX�$4�b��Đ����`�h�X1 �FE�!5
�r�޼6�[�n_	&��.`��B���#&��Gs�9s�=+�����wd=ٿ�כ<���!#$��2h��[�l��G�.�adJD��`@
�XHQ��B��2�K�c�H�k��H0#1�ɐ���Mʜ+�.�Yt`JfO��u�y�Ϸ�O3��h�c����Sq��fn�o�S�6����iB�����]̲�%�d�a�*�¦�de�~�����}��JI�~j����S
Q��G��O4���l�l��"fkg�K��'0��\ޤ��>���k.fHX�ۘa��K��3�yυ�^y���������	&LO)�5D�NRג޷���G����a%
34J2�,Ĭ�-!1%��RBD�.B���+��B�a@��R%�2�F0�fX5�q�0,H\.�����"T�>�`/��]��Poy��o�����'���fz>@�� w��xr��,���'��x��r2:6<ay�)T0f�����Ip��s�sd�y垱���3ͳa��2����<��WN��&�4؟y�{'�sG��6jY��Yr>�r���H���"P>�n��7���y�ϧ��n���}�KO9��	�B�&�.�����Hzo�@8�1a�>�&�0a�4�{�͙�*F��ZM�)�+�����K˞���	,��G�(���>��:.r.�H�1�p�,�
��p�|���P�C��I�szHC�:�Zf�����+�#��bHBA"�H�#@�CL�R,C	,b,�bC����f&�R� 5 �0}I���$I����.��&���za�<��xg�.I�����\�\Y�K1�ȗ�v��a�-�d H(Fc���"�"K������]nI�C{%ąa`�D
H�K�F��`\��#1���!)"J�-��I ����B�:�H��%16{�$��"�,#�^L	�{�W	���)#$i)i�{d����48�$��%1Ѭ�kz�'	yf�&�J�;�2�OVR0��j�t������]�tE�||�N��qރ9�e3w4zM�&�<+O���!<�)MԪ��i4��-�8q��a�FT�0�Sr�5�����A�6�z�C����v��i�-faI�f��緜�	&S��d�KH�!�ٳ{�?]��9*�iUٵ����ͼ�U^�x�٫ra���y�\٢ @��y��	����8�H�ҷW0�%�R���j\%8fh�X�FIB�[�m��5���Ͳ�Mn�X2�*�
�io.�����;h��g�e��5��d���7�.kc��|8{.�I���Wy���P��B���y���0��C
���6�ٻ&obv^C�BB��wcb�;ϗ�w��ϥ<��Td�UF�"���ʥ��jH0�A���.|l�]��H|�������4/�g�#	F�$#��=�n�\�t��ㅔ�_2l�[>�o��8f���)=��Rv�e|�F@���4�S�Hj�R3��*b�R���7���%'0��W�&�nN|Mf��$�٩�y�Hf��~\3���p�s��Y��%�e~%��5���Vġ�
D�H%��m	J�!ݓ#�B2����so~rJN�
2$r����! �G�3Z�{���<��'H��B2$bI�ZL K�\3n�a,w����y�@���F`JČ�,D�����߂4ky����z�^a�||��E�,�9
�T�tA ���`@�Y E���$�z��{�68�kf�%0���D4�YY�P$a1� � �.��]����{�y�5�޳K��8��"��^}�n|�9K,ܓXS)	e=��8C!��!V&F���y	�"cR]M��ٰ��P��fm6B߬���3�4#8g,�2�ѩ��.]��{	]f��<2ٻ�=l��v|���	�'t��w���g�5|�{BWS�Mh��� ��ݧ���a���d�����@�BH.��B0$bI"B#u5u�FYR!T�V хB5$	YX�8�`�"�)�rjo��)HЁV�0	~�W�f���
g��ܕ���ܳ͐��XB{��כvE�p��c�����T�+$H!#|�$J����Y.fvL&J����}�P�Ԫ)*�Q��P��������I����{��ӓy���l)�_�ɥ��/�$$�M���������f	t�>v�C��,`|�.ky��c	s~p��r�P'5�V�s�h0�[�}ϓ���S;T].� Q���WFÆ'�)1�$�jf��w�Q���C!y��w�N����ӻ|�p���o;���˧ξ�ݲY�8�D30��o�]3�+$��(�<�1e;�%�Y;�#�-��þ�S6��n��y�%)/�m,8n0��!!�K5�a��C�Ri�c	S�ק<#f�!�{���ҢN�߆m��I=)��뜛�L��^{�B����A�Y��w��5�%���� B21�	��>�=7t5΄����c!Cf�Ϗ.{���L�=�����h\%���79N<��礼'���3A�xJc$�c�.i�
�a
����rx�`Njo�n_]����)<�d7�!!�Z8Ŧ�a8m�SVo��=��<�<"C��əw�Op�m H�e"�
�B���H��[0��A�$��i,$���, E���.�o`h8'$�2�!n$�7Yvm#CN��\�޶��K����Դ#B��s	iJY��ɨؘT����%�#uJww�HK!v�i�t́����K�cK@	��d!߽��>�g��k�=�ԩ���W9�&鳓Y5s2%IIi��f��ׄ(�k\7ta.xI�����y�y���$�B��"J�f�σ��H�0A�cHBA��	_#8M5���ЌH	&!L�#e"Hr�%�0�Gn�/{�޶|�;�,7������,��B�5���Q����&b@���}�P�	O���s�u��l��%��!*�) \&d����с�a���$B0�ô�23L�p�K�|A�>����t7r�)��i�$��_!��~o���o�Y��d�5�_���<=מ�v��0"�Ip����\���In�o4l�Q���Ҝ��[�!���� ��>l�0��4�$!k
Q�Z­,$m�\ް�0�N<.�ɷ�D�򇐄XBz5HH@�	�Kyk75��!%	C���GXk^�r��!iB�L2%`����G��V��"B0��\�m�y4�V�B��j�	B��Z��I�O��xHJ1�*B��c�����_9��HY4F�2$Y�'�@C�R�b��
���,}%����3[�l Q�s6���L��-�̶o���5&����7������o���ɘ�9����)aw�xk�l�Nj���6���B�/4�9K	�y�ߏـ��<"~��!���]So��k��1w2��r���K��p�;��!�_n�x�%���9ƟuUUUUUUUUAUAUUUUU�l�1UU\5UPUUU��z�������UUUUb����������������*��Z����ڪ���h�������U����������������� ݝN
����J��}UUUUUc�UP@��q���VVYV���
��[���;$r�3�*iXK��:��T$fͶ�U�UU@UJ��U�e��v"�r������UmUUUAKUU@UUVܫUU*�*�UUR�@�bJs=�]�헗iV�`q��j��ej�]���IK���ڧ��5[/<������^L%���n�zLwYz̸fLB���\��z!ڞc��O�x��f�u���*��R��*��	��`�a%���clF�X��*�e���膳at�SWUR�m�h ��[Uf�UU)�6B�Z�Uy�v��Ft�(��i���r�*�������֩���-Ҁ��Gj����P@;//+V�9	�ꪝ����FA`l�qpb3���[k��rK�����+��ZSjšٔ6%�IA ��cbR(-���	�V����A�fU���U�}�}G[�J����[��U]�*$�Pg!]�[*�J�Y�HL��R�l
�mUJ��+J�uU�d:M[�U�UPlm*�)5�IiH�j�a�����
݀�P�U�\�ҬdZ��@��Y*���U�Z�����X*��a̻6�V�s��UmUUUUuR��[V�UV��PAZ�båUJU����X
8le�f%ꪪUU��p1b�k�ݢ� �mJəy�ZUP#���tU&EW�j���&������R�6�hh �%QX�X5Z�1AHݲ��SͰ"mr����a�����ĳ �)e�dB�����Y�u-��܉�Y�3i^|��ۜ�!s]�2�P�9�,�ڴ�6s�P��)^R9Zz��6��4 �sm��`9[�[^ťu�UG-�WTh���xgD���h�N쵎8(�S����y%�.�Fj^��kp\�er�ֆ���-�u���s:�	V�laĲ��go��� 뭶�
�d6+ �U^vn�[UuF�G	�*�g�!�ι9'6�@���j�
 D
��F$�@�*E`�kOh�yz��m�qZ5U+�U]UUT2(P��UN�UT��Tj���:����[vݮ��5��UVԅ��[\X��*�\����,�U<@첻1�@uT��7U�U�ZC�%VRW`���T�e%j�N�mU<����h�r�mU]pj��b��9� �J��@j����U��U����b�P*���#A��mUg�|8b��<�X�Pq�«V���k=�����J�Uu�*�ҍQ��)�궪UY�UU*�UUU�]��ͦU��q�*�7/2���٫j+81��v��*��Y`e�8Ӡ j�yڪ��cT�cUuJ��Kr[-n��*�說f��H��St�`X�Cm��[UUgeڮ�/
��KU@U�]�Q1��h5�Z:f�X��HU�j�v��vvm���cS�UW[�����U�����}���)V�*ꪪ���*�#*�
�U�b��R�u�R���-l�&���]�jڶ�ݗV�Fi�W�U��^yW=���HƁ+].vU��R
�����k�Cr���f�*��`��ځ2�Z���Z�gqJʻ�ӎ-��5J\��lU�A�ꪯ)-uU[G9@����At!Zh��Wz�
(��#*����[+Q\E�Xo*��j���ŋ�
�x��Uct���B�*� ƙ���+��J�*ŵ�:�ꪷgʫL�Uj��z�§}��m�c�3m�cŠ�!3�1�Wh���i�nc�R�L;��X}��Vy����m/�$/Z�;&)n��=!���qr��a�k2�Z�XYQ53XW1�\�8��"�\�6/��;!�kpݭ)���`\d�` ))R5��,��H��`��quoe(rZ�v}m����h�4��1�J�Ci]��!je�T\=�3�)�c�)��U[SmÊ�(3�s���B٨���mX@����yS]��� ܼpJ�V���l�l�*���Դ�kbYT�������P��ϷI���N�I��4�#`�-�![�Y����%�^`ۀ�%+	̨�Q�.�vT���-�#k�+���+��R0��m6�h8�M�6��J�4T��M��bJ \�C���u*ܭkb�a0�5�ܶv��s�ʥ5�t+�r�T�Y�Wn���>=%�iS3��y��,��:�w��Jq��)6ʶ�J"@b�@��j�V��k(z� [�u�@��e�Ad��tc�6c��F�e'�a���^(#���P*z=dҸe[uvܧ����az�z�P;k�1Lq��qs<��.X��vKSJў�ŝ.ۃ�Q����-��3���� �j�KC��*���W�D�/'~g���::±�@r�[�T8B[��X0��#]�]v�����7P@����v-�[q�l��8��OUv��^�+.��3�ۆ��竏1�2�v�k�!�i
��b��h�ʠ�R^��k���T�}��|�GeL5[�6�����ت�
U��j��we����Z1M	�볫4�����PGl1o+�T�C���+�k6��7�cI��t�QXM�R'N�Ŵ�dZ��%l�mV0��um�R�<ڙDcpV���6]q������u���mm[T�6�fF�]t��U��"�n�YZ�^�����u�¶�@V]���j��
�m�j�;V�+���J�UWUrd�cv�����k0L� H�U���Q�t�ʮ�յT��$��U���5\�U]*�P�Ԁf��)g	���:���*�١�LW`�����!�.�R�*�UUV�ݢ-r6͓Wj1�-e&dN�" ����^����j��|���t��3�@�2�( ����)�
��imZ]��,�e��X�j� ��ʴevh�6��)�5U8�[UP
�U��]V�+�s��i.=3l*���� ��
cUUA�5���l@WT۶�9@�mgfc��X؉n5�V�P*�A�݀�n�Kh+nƕ�j	v{nϒp]*��a���ca����^ə��&��ЇRzC�xS�ݑΩ������6�X��,�! C!V�	��{g��-8oa�+�q�s��2�@���̛R��vPZc�d�3e���Q�X��Kѽ���P�T��j���B��8DRՀ
�[�nP��i
 *�*��Q(����T;�W[*�TF2嚱��]!��>��:�6ˆjU��;j��.��A7UJ��m�+���=r�3@��v�A��D�U*Ύ�J�;7Y�ڪ۞��'\���ji坬j�ջ5v�R�,ۑA���S�X��n8Q��;ҵ����	�/��c9����m���ډ��kk�]s�z���t��c9kT�nWD���[ueK\�4 ���B���"� ��P1�l0UU��c���� �X��P�]�C��J�R��x� <u�ɍ�I�1���p�N�ˣ�c�jJR7I�p��UW�d��[��d�5�wl9u�6���� �Q��
��4�R�\n�n�Bdɴ�U����M6�W4p@<�ܼk�Smv
�"1:��+ET�UU]UUT���U TUUUU9�֭u��⋪��۰m;UU�l/Eԃ�(k  �U�y�n��/8��E���QL�RR��(��gb��[v�n��Em�-m��B�[j���
���틝,V�=��jUd,�5�5��pfʪq��Y��Ӣ�Vҵ� �n��j�ҍ���Uc�j��SW*���KrOIe.�������c.��fV^Z�,�.�]QE�FV^٪^8�jt�l��V�PUUUa�2�i��Wf8,��j�m��R�Ί��1�m�V�@���ꪮu�������U�V�xu��!Q��6PWj�( �Z�������cRUUUUUUUUmUUUJ�*�]UR�5����MG}<o����j��ڨ�` �qv�X�^&�Qb�vUj�j�vYyj�X𼀡3��UUU]�ʵR�mJ�*�b���U0UUUT�UR�� mVn)U UUUU��`��r�THM��Mh)V��T��
�e^��y���P��n��T�sIns����:���U �V������ C�/d��UҐkw-UF�j� ��U�*�;�V�Z�ڥU[h 6�m��yv����jy^���m�j�S*�U`���l�����m��K]U),kL� ! P��m�/6�o#Pdζ,r�eG0u����n�R[mł@׎��Ij�������S.�U��݇���G�·:؀ꪪR�uv�`7:	I	�*�l9��u���7b�cRÌ�ŃFnj���f��57M��,��P�r
�p��Eє��j�!nd)]<�۵,�:ږ�XF���f�*ꮪ����UUJ�ܫUUU*�UU����Z��� +�z�SUWUUUUR�/9G�������������UUU@U�e*������TUUUUUUU@6�� ������v� ����
���� �f2գL���Pvcv*��������4"�ە�����^�Cf����v���T�]uUR��Ut��UUUK�T��X*��Z���\�R�UU��
�������eX
����Zڥۖ�UUUPUUUUUc��������h
����U�WH�UU*Yj��k��>��j����PR�R�U]PUUJK]UUU@�UT�UUUH
�U[UmU6U�n�������U�����~������Zϑ���5sj���E��]����w�5I��UK}�e���;�T�����:P .�D���(�O�� b?؊1��#�B2F$�#��M��� �"��@
�WD����DC�n"�5]��Zx���*q OЂb
xP6` _Z��"lLx�"��q���'�q_p	P� �Sh� /O�DN��H�HB2 ȈB!A6��=W���>�����2H�$,H� 0��`��!�~M�>�A⦑�G傇|C���>лb�AX"@ �R PCj<"(z�P<F�XG��!�
�6aP~J���� z�$A�Db@DЅT ��|��_QO�������� *mFp�A�B0 ����LW��j��D"�� ^D�E
U�@= !�D��'�`���5��+��|�)@x�Ei!��C��`����Z�@(�J��T�EB��;�C�=AH	T��� x!� �b
x�}!�iX�6ФXD(�d���B`dB��$�im!l���-��!Q�H�da!YZ�ư�cB�J�RX!H�!B�eR�H0���Q���H�
-�Vr�1'��{�>)61Q�B ��EOE��"hU�!�!�� H��U�	�D�@*� 6�:��]��uB0R��F� ���C�P ���q�)R%P"��Tը�R�9/8r^BC��UJKZ3[͈
ڪ����U�����^���9Z�i:���9�T�m۩P%�j��gNCP�V]����a[�ݎ.pO:u�ⶭ-���l6&^d�r�������X�\�)@�Fi#�Rv��2��ҵ�&��+S�m�+[V�F�$�{0�M͹؞.&ݻqpv��I������}t^��"s�>:y�t�J=�*��s)���:8T�.�G�c��@���q8��6�c�l&��7]�F��1K4� f���l��<Y.�m̖z���M`�@2��[z�s�$C
wjkuf���2X�X9���Z�*yɮqsq;���+�i]�7\�z�.0���e#v�	��L��A����pm�5����s��-��ZQ����Mx+(M��q�ktcى��a��G��bNN�粼�e,`uvc�gl*�Y���)��:9�-q�1�gck\)�l�d�� �k�&��f��5ZD.�֕�t�vr��C:�V��5��4���x��VA�{Qoeڜ�rÃ@'s+�`0I\J��n4�a�a�UN52�M�g�8-1:�ql��u�жp�)���z���c�0uam��{�՛��ħ�8�X-R�rc���n���-p�m��9T�Z�g�$��88����,W�)��7H=i�n�}c<�u��j�a2��Ɠ7����]���\X���qm��-t;vNԢ볜��hZ�`ۑ�W�Vvg;$��j��m؛[mҽ)Hĩ0٦#l-!&�l�Ĵ���YMa��PŻX6R�fU��`[Ga�k-q)j�K�⪣`��YK�"�2�B�6��0d��*���9�D�`�@T��"��x6��T�<��:���<={e\qP�&��k]�a8q�78;t�mT�Ui�G\P��B��+�űAf������N�sv3�`9y��Zk��6��`%�b ��Z����j�*�V���)x6%#��%^nb��n���-�&kY��T��6#�D4Ё����ب���D<N!⁴>U}Wk8NI�y�b�:A��@
�3.vے�wb��5��H3uZ3]5�[��0���=;�F����"����l���/i0�ҫ�1�[���^'�nv�j9zw$'�A l+��-ܤ�5��@��&I�!Լ]kp�e��3�t�s�np�v9b뺮��2@W	�D�Я$v�V�������溷�0���E�y�t2���;���9�����������\�yܩ�rm5�Ғ�ړZ1m����5o��M��}�t�Ž��>�̬B���:Wt� �ve`)���&V��/ ��#��&����u�|���>�X����+ �u��)4ҶXQv� �d��5we��X��, ��[
m��V���X����+ �k��ɕ��'99�<���[5�)5rJ�qh�+цt��shv�,9j%����p(��@�)mӠVU�wn�w���>��w�e`���஛w.ʻm2�)ݺ�>��}7�N�A�
@0Tt�{��V����+ %J�eږ�����Л0�L�Wv^�ɕ�}5� 6�[WI][,v&� �ݗ�w�e`Kذ=�W��`�~�,�N��;�i��;�2���x{&V���w�������R_��&e��ױ95'$�;��m�HpS����3�GPxJɎ�P��%I���պ��O^�ɕ�j���;�2��QI)����2�x{&V��/ �d��>Se窹ă��/ʚm�E[���� �g� �d�s��j�F r{����y��0�R��[m ��T����X�\0�L�Wv^ |��Hv�1��۬�{&V��/ �d��}�}�Ԫm��:Z��֣�0�[k�h��Yq3���"��	�Σ��+����N�&���+ �ݗ�w�2���`�P���v����`�����r�I��X}��ɕ�H.�\;�k��� �ve`v8a�R]�{+ ճ׀ot��Q�!5t����c��d��:�����T�\���V�����&Xr�ـ}�2�]�^����>��z�������qm۷ p�X�[Dkj 4j[l8�%Fw6�&":*���֕��ۋ׀w�2��p�9\��;��V W��Ixv��!U��ݎ��fV�ݓ+ ��%�t+`��C�m�E5n���xݓ+W)-[^�=�����VF��4Ӻf���w���[^����>��]@VՑ�V�E[u�uwIxvL��vL��\�\�Q�j(Z�7\�LC&{=�������Rb�j�D,�,s-l�[6�Vl�ճltÌV1<n�u�5ڛ8��F�LJZnd�a�,��˙��r��Oݮ;:�ݖ�!�93��-V؇d�v�Ɇ��CqZɹ�/��m�'&����f�V`�)��t�4;�z���?s���S< 2 l�ӧbvS�l�\����iy �Ʒ7E������I���{-�c��q�������E��ct.sq�Fj�b���ƃ��ΎF�j;�y��ݝ���&V�ml��jL�$ձ�I��>�p�;�e`v����2��R���I+V���wd��>����;�e`mȰ`���n��V�պ��\����~�d�V���+ *j�+�n��Yi���ٕ�}#��ɕ�}��/ �*����Y��8�-�#
%��rjnqd17!�v��벆�qlƮm���y�m;u��~0�L���ܿr�\��� �J���׭]�i�t&������G�E���)%�I��#C��Sk$ֳ��nIϾ���}�"�W) �� �~M���bn�����ݙX�r,d�Xe.�ʉ�;m*����{��+�{�����^�ɕ�}�[/ ��U��DMUղ�'n��d��+ ���^ݓ+ ��>���u�@&rMn��װk��͌i�#�{3��|��{`$m�8���Gj��;�e`v���;ݙXݽ� ;Qm�M4�t[�lj�`��vI��}�ذ�2��e�.[�t�VZCV� �+ ���`ꪩUr���/vL�{ke�t4"�heջ��J�`n�`�e`�[/ �+ %J�wwR���i�ui� ݓ+ ���xd�X�Ȱ�%Z+�㲒�u��j�f��qu�aK֎����G\Gr�0T����N���lM�6ԗ�wd��5l��wd��;�/n��+c��g��ݓ+<�I�<g���M�r��^ڗv��-��M� n���X��xvL�aA�L��!��xvL�TR<�&VW9�p�$�'�!''!޽|�����x��.j��X��x�g��|�{� ��{:�&�ݮ\����!�,c
1���لq)���hg�(��Z�p-��&��t�VZNշ�wd��5I/ �ɕ�E� ���KN�eջ��J�`���H����<���vI����j��5vӷm6��&V�)�&V I#��x�`۰l-���5E#�;$��$��&V�J.Yw�wV��w�]��vI��j�^�����=����|"1`�"���" � 
�U
HAY `@F!B�!v'f��q��3I��7�@tmmˉ&�Qne��������S�<�8����&0��q��V�1�)I�f���A����
*h�f��]��6�8x�%a�	.���������^�@n�`�m�d��ﶾd��u������ܲ7�[�:�8��Qk
ke[QRN���6�k���.gn��J`�Q�OWgjyn�����f�B]�Ĝ���}`K�X��PlT5�)f�hK�Ml���B͎��bGH�Eu硻nfSutv��@����nɕ�DI�&V!Ab؄4�j�ݶ��2��#�;$��$��Ce[V���V�պ�"$� �+ �r,vL� ��,���݊�V$�v��&V�Ix�X�H��D���]7v�Bn�RK�?�=��"=�<�'��o�;l<��+-�`8��a��`f�&F/,V��F�<k�D�	:ʜSX;M���;�� �I�&W��W�'�� �N*'�i�M��l�=�����bT�DY*�
� �"����)�+�5��ٹ'�{�� ݎ�(�e�%�]�Ӻe]��vI��l�+ ݎ�$x{AZ�R�i��Z�M��L�v8`ԑ�fǀHQj��T�E�ݺ�7�� 6�� ;6<d�X��9�׀z��5[�k�y��6�[���P�����3��	h9��CS�sZ0jH��%�$��$����D��*�����xRK�6l��$��6<�URDZ��5c.��h�V� ����&�;[*�U�,e8�U�c	w�69��0��y+���m��Jy¯�<'��|�}�CF�$!B�k)��7)�`r&���y8�]f��r�w�!�9��w=�&��,��k><a�M0�CC��'� �oԙgޒ��|��$d<�53Pp����Ϗ��mΒg	���s���\�y�����vs�DJ$���X�,�}�����]�`�O/��,R�����1<�f��8��Bh����5��B� ����z>y�1*yS^h����ĵ�6l��>rau����(J��D��1�@��Z��*���<�d�(E����1	�$3�;76CZ#"�HF!���XZ*Z���F3���bn[$ZQ��M.:!͓��@��ߥva����6�P�X$ȓ��
V�*H:6x9����x��{�	��!HB)�ԫ�1מeB2�!����}"�����s7���J��n	�F5E�WB�F���E� !���hE� � � x�*5ЀP��<H�~ M$W,����`Eݗ�T�+�D�`�6�[o �� ڛղ^��Jzy�ki<;M��YlV� ڛղ^ l�����#��-+�c��5���5���Q�H�F�	M,� 1m��<�*	�#]��j�Ɲ�*�xT��fǀn�s��+�� ��y?UӺe7V���x�c���$I�� %{�xT��ܤ�ࠣޤ�- E��'�� ڒ<<��{׀���6�l�)+m�6Uݵn�=U�RR��<W�����nL|Y��$a�QB$T� �E!!�,�����v~�]��:|j���Ixk�W9���~������V v�m��twͲ�	]kh j,rK�F�Ԇ��]�T8��Wۍ3�HvX�;�3���5�����6~��7d���#�|�W����W��<�6Xڵm�vL��	��x�{׀H��s�.�j"�߆6�݂.�n�ߏߞ�$� �G�nɕ�}ң���%����,��M� $��l���� �x9V�5�v*��x$� �\�s��������< ����rk��E�;����-%4x�2�sm,�v �e���K@�z���y� ����^��s��Ρ;���������qi��ɺ�d��ۧ�x�Q�ݴbp�����ñ r��ؕm
�BBT�Æ���D�E��(X@p�Qt�"��t/�^�7[	��-���hٞ�s�ЪD܋'aΥ���e�ku�`6��q)�e���]���� lw|�Ix%ɵ���3�W9h���SV�4Ȅ�ж,X|Q{)�%,r�@!j��;H������� 7��|����v�=�
I��6Uݵn�a#�r��������̮�����߿�v��1��v�z���H��U~�W+��������~��	���
�њ+�e_-�$�@�����;�� �H�=Uʤ��� 6�y+��1�X�+V��;6e`�R�=��o�x$� �M�\�4�I�;T�fq�m���8t@6ɶb�a��c	���Qlb��9'l� w�f���J����ߞ�d� �G�r�A�=��wJ�Wv��m����=�{���χ'9�}�䟹��g�6{+ 6<�UU����j _��&���Z�� ?~���vea�q"x�����.���x�9��=�`��<.�r��K�������)&�@�Wvպ��� �*������{� �ٕ�~�r�U;k{?8�ڦ��F��P�����D��Sd��e���D.@.
P���s�r7�.��[HUc�We��?)�׀H�	ݙ^��9>P=�~���}��jL�3J�v[x$�=\�URG�{+ %{�x;�|���@���~6��5��a�����}ݛ�OO��[�/4�,B�X*a1�E*�R�2q*�B�S�Do����nI;����Q[cv�.�n�=ʤ�{�x6y����.�{��;��]ڢ��Ս;�U�x���W9K����w��X*H��[����;vX�,#κ×�!�ss�l7 �ѹ�^��4��q�ӷ�$% �;.ך��9| ����z�0T����W�Oy��b�������	��?r���\�]�����������<�s��s��xm�j��ـ���l�W9�URD���=<�`{�+.��e��wj�m�{��r���x'��	���W9�TD~"�x�@�.i@�j" 4 c0 �%t5�@@�� G�m�_9��ܓ����P����nۻv� n��W*�����, �����z����X���r��Z[�UWy��9��ݩ7#Q��d[?��;c����Yv������ ��"�	������W�����[M� ��K��ʪ�ʻ�������'c�{�Hݠ�R�)z�XӾ2��O^ l����\���U����V z�~���Ejh�]����[�{�nI�{ݛ�OO��[�� �U���^��E��am� -��	�2���?s��W�ߟ@���׀$x�9�(��@:Y��eN��a�w��\]jRm	��n.l81B]���g�����p6��t��D�� �5�ia�u���Mm(d��i�5͌e#��^��v�	(q��P3����i7����j8u*K�xB�j�kvWE	f1�1Y4Q�Z[ %W[��7k����De�/]sm���m]�zظ̭��Ȝ����\�6
&��&�� ��T��0��#�@�ΊQi�f��r�Ye�ۇ@
�k2�;	 �\�,O���hvw�[����v�hG�ߞ� �G�UW�=��V n�����b���v������fI����ܓ�߿lܓ�>��o�	IP�yl�E��m�w����	�2��9UUIy���'� ;R����G:ŗl�C���?�'$����y:���~��y��w'EB�����Ӷ�y���˫m�$x����U{\�����;�+ ��B�K��J݋N�����2��i.3ob�g�kp9�j7c�e�m��rs�����we����� I#�7�2��r�ϐyy{� ځQ�^wvP�W@�X�G��ӁG%qR�"z��B�0+GZEI
ژ-�a!	���`F"�W�F�+Ψ��w�ܬW�����Y��s��<Qr���Z�Hm��M���"�G��\�%�\��	�y��D�����
l��n�=UUK���<���$x�+�^��Հ%��/+N�Uc���m�^ŀ{�\S���z{+ �)�/d�j�����V�֔�ة�����C2���B���Wd�:�_��J��xګc)�n�m|=�<M�XQH���*�A�\���@�E�1۵Mһ��&̬�_��UWg��~��߯ߖ l�竜���js�I_�[��E��u�yy{� �������$�E8
:dh@,��@ B))$@�*�"�`��V
X�S�r�����=�+ �h4h��j��N��[x�s�����	�y�6e`{��qz����;[G��^Iڢ�Wƛ� ���r�==�|��~x�c�"���a�Qv��y�k.֑���,�[�����L�n#kU6G_ӓ���nԥvÖ�z{+ 츥�͏ܪ�9�g��	[G��	ݻtS���u�v\R��
��W2N���nI>���ܓ߽�f��A�ZJ���'Ö�Uݧx=<�����? 	�L���훒}�?_ٹ'����Z*FU��?s���[��ߞ��~���<�>�f��x�-�$`lp1p��C$�ti�!�)��00�04���E��lRuD|�w��rq�/�I/�3��f�Mh���kiȖ%�b}߻�iȖ%�a���߷��ͧ�,KĽ����r%�bX�߻�m9ı,O��K�������z��5��մtT<���)л��Zg/m�=:wv�;����Tԣ�ND�,K�뷹��Kı>����r%�bX�߻�lPND�,K���ND�,K�I>��'fan��Me�m9ı,O��w6��(6%�b_~�u��Kı>����Kı=�{�NEı<=���ߨ�\��.���^B�����>rr%�bX�w���r%�"�%��u���r%�bX�g~�m9ı,O~ ��_ʹ-�a�����NJNI�"�dN����"X�%���~��iȖ%�b}�����K���� \��w��m9ı,N���9Mk5�C2d�ִm9ı,O{���ӑ,K��0��߮�Ȗ%�b_������bX�'�w�6��bX�$C^�0$�9O�ȳ�WVb��l@Ѹl��L���n��٤6.�>�x&�xp	��H�a����,�! @��V�`B��i8�� �r��!��1��!$H�d���H�I��N� #(%ٯt�� ۹����˂����o<�6�C��sa��5��*R�a)PVڪ���t5�UUj�"�~��,���d��	�@� m��  �M�c:X"#hv��miJR�GgMM(X�r\�Ƹ2ZLkceA3¦rN!��eۮr#W���R��Px���k��Z�yf��������R��L��I�dr`pj�����Nr?v�j�,����'`wF�-�9\�b��KZhV�΅6�ف�Н�^n�pű�8��k(�ac��\J�&�����T{kj��{��'*�6v,9U��\�ʹĤ͑����A��/J�c�NYz8Ø�Y]�q�Z�%�#����f����v�#����w;J[&��:!ܓ`r��i�f�XذBPV�Krr�ɽV�Akm�M��hцc2g&-JE���2+�MQ�' ��T�V�\�L��:��q�a[��	D.����I�)X/*C8(��hi��ґÚ�b[��l����N� �֌˦9�B�e=��<�Dvu�Z��0k`܄�����\�;n4�݂'�* ���2��j+2MzU�0i���������`KPj^0j�CGF��2��/ga�媬��S�&�\�r����5	�(��6�]��8�h�=�l�g�� ����u/�絩�ܼĬ��لN��Ɨ�r�ȼA���{� s��v��j��b�l�fH�{��1e\L��l�0Ɗ�,L�WX������;�âӲ�^� �V{pb7HܳrηWD���Z;�َ�:&2ےڶ�d1�+T�<��\�AE�P�+-�#k�mX�[0F�c�u��԰���h�P�,r��ڼ�\���d��#L�H\�I���B6ͺ��mFZ�{`eZ��u�*��FŔ9���eÈd� j�Q�)y뱬��D��s��Cv[�����I���^ob�d೼�M��\\aԓe5�I�62�4x�
���m"� n�0V�]z������d��L��&� RR��)*�V�z"m$#Z Z�e����v���45�ֱ@�O�����=_WH� =^#�W�S���%P ҉��L~S���b�U�Ǜj�Jj���b��e���5u��Xu�Ӂ�ͱͦ��`�ಳ��Ϛ�&ٱ;��d����-�M̼�P�$��!�j�n��q��jە9.ؙ#{gC�m��V�!�"ۂb
��L�te�[��띹R��ȧh�v3&���d�Vv���9�p;���rq;���![f;V��S7l���rIE��f*�a��m�cc]���E������'v�~|!�c�c�1������'k�b6�j�n��@�Z6������!q�2r��iȖ%�b}����9ı,K���bX�'�w�6���bX�'��osiȖ%�b}���况�h��ֵ3Y���Kı/�w��r���"X�w��ND�,K���fӑ,K���w�i�"6%�b^�~��~Q	�m����^B�������r%�bX��]�ͧ"X�%����nӑ,Kľ���iȖ%�b_��w@����\�<�����I8D�;���r%�bX�����9ı,K���bX�6'�w�6��b���}/I����:T��r{y
�%����nӑ,K�/�w��r%�bX�����r%�bX��N�6�JrS���w�ߒ�2�&��j�ۡ0t�c�'mɠ��u�(�t��T�ew��;ް��i��r�(��'Ò���%����ӑ,K�����ӑ,K��:w���_"dK������K�������`�ʹ-�a�����NK�����Ӑ�PجF0�%kh�"֒h#E��Tr!��X��-"��DIq,L���ND�,Kϵ�nӑ,K���w�iȪؖ%��~���D��Blb���|9)�NJ'���siȖ%�b{����r%���b}��۴�Kı<����K�B�w��߱�q6��r{y�EKߵ�nӑ,K���w�iȖ%�by�{�iȖ%�6'���siȖ%�b_;g�c�j&f��fj�9ı,O��{v��bX�+����"X�%��u;��r%�bX����v��/!y�߿���S��D�����p��\�m���Q��]�P�c
�^ڷ�tK�1�L�2�r{y�^B�w��M�"X�%��u;��r%�bX������,K���w�iȖ%�bxw��~���"�9=���/!y>�;��r X�%����nӑ,K���w�iȖ%�b{�{�iȣbX����{l�1��]��gw���NJp�=�]��r%�bX�}���9ơ�A��` Ț����ND�,K����ӑ,K���N����p�Z�Ys[ND�,��S"w����9ı,O����"X�%��u;��r%�`D"('�w�M�$S�wM�Лge<���Ky?��^O,I_���ٴ�Kı=���ӑ,K���w�iȖ%�b}�O����h��J���g��tc��x3�j����g�q�iy8gsp�E��!��6
��)r���bX�'~��nӑ,K�����ND�,K��ݡȖ%�b{�{�iȟ���,K�{�)���M�kW$���r%�bX�w��m9ı,O��{v��bX�'�w�6��bX�'~��nӑlKľv��f�F����ӑ,K���}۴�Kı=����K �,N�5�ݧ"X�%����6��bX�%�Ӷ�C/u��fh��j�9ĳ�"}�߼6��bX�'樂~�ND�,K����r%�`~N�"� ��o�j�D��~��r%�bX��鹖�?h�ֵ���h�r%�bX��k��ND�,K��A���~�O"X�%��뿮ӑ,K�����ӑ,KĽ����HѶQ�Kph��՞c����<`V)qkf-�` %׆������{�?<.���ND�,K�뽻ND�,K��nӑ,K�������Kı:{���9ı,O=��nfgL2�j�n�WiȖ%�bw�}۴�Rı,O��xm9ı,N�뽻ND�,K߻�ͧ"�%�bw�M}p���l���ff�ӑ,K�����ӑ,K���۴�K�,O~��6��bX�'~�ݻND�,Kӧ��fkXW2d�ִm9İ���۴�Kı=����r%�bX��_v�9İK߻�ND�,K���r�ܷE���\&f�ӑ,K����iȖ%�a�b�￮�Ȗ%�b}�߸m9ı,N�뽻ND�,KivTR�i��ل��j\5��K�cX��q�M�͗��O�*7Y���쌱�"�Tv
C;h� ���Xږg[3�A�sJqb�_(����V�Kg(�xi�73�B����qv-��4��"Lb��qr�2�`�3-�d����+�nkM��qms�Pc6�uڕ��i�L�u�-��&X�+MA�5 �*Ip�����1�OM� ��lK]��;Z�u�N�;�'I�>z��@i����.�:�Ͳ����(�7a�p�4X:�	�����׼�5�:)�R0T�'Ò���'�u���Kı=����Kı:}���D�,K߻�ͧ"X�%�;?O���o�iV����^B�=����Kı:}���9ı,O~��6��bX�'~�{v���%�ק������}[�5��=���Mx�:}���9ı,O~��6��`%�bw߷ٴ�Kı=����Kı<��]�;3$��WXY���K�B����iȖ%�bw߷ٴ�Kı=����K�V�����r������ݲ���a��h�9=�bX�'~�}�ND�,K�
����ޛObX�%����v��bX�'���6��bX�'�}/�l���K`vR��npX8�a��3n�(`�3C	cho�T{lJTRo�'I.��%މu� �o�*X�%�����iȖ%�bt�]��r%�bX�����"X�%�߾�fӑ,K����nr�sXG2d�ִm9ı,N�뽻NCZY=�M�6��ș��{�ͧ"X�%���}�ND�,K��ND�Dșľ��r��.��kW	����Kı>���ӑ,K���o�iȖ �X�'�w�6��bX�'Ou�ݧ"X�%�|�쓳Z��Z�F�jm9ĳ�U������Kı;�߸m9ı,N�뽻ND�,�@�=�wٴ�Kı)�Ӷ�/u2jf�m�M�"X�%�����"X�%��f�۴�Kı=�wٴ�Kı>���m9ı��׼��c�p����WD�6)؍eՍ���iI�3GZ�+�,b��;�R�ǖ�]d�f�Z6��bX�'}��nӑ,K����fӑ,K���ٴND�,K��ND�,K�g�ٙ�rB᫬d�j�9ı,O{��m9�0"dK�w�ӑ,K��~��Kı<鯻v���%�by���lc�	Z�Ao���B�������m9ı,O���6��c�P�B��F%X�d��@�	 	Z4��$�+�"l�2&t�ݻND�,K���ͧ"Y�^B�}�����+ &3vo���B���'�w�6��bX�'������Kı=�wٴ�K�lO��}�ND�,K㽝��ff�ɒ�ZѴ�Kı<��ͧ"X�%����iȖ%�b}����r%�bX�g��m9ı,Oʽ���3<�Z��.k2��j2:����W#(��d���k#=��lU���%آ��.�D���zk�^������ӑ,K��߷ٴ�Kı=ϻ��'"X�%��u>�m9ı,a?�C�_���+�7�Oo!y�T�߷ٴ�@�,K���ͧ"X�%�����r%�bX�����r'�Q�$�&9)�g��L�%0�'S�,K��w���r%�bX���ͧ"X)bX�����r%�bX����m9ı,O�>��W;�K�fXfMf�iȖ%�6'��o�iȖ%�b{��iȖ%�b{�wٴ�K��3P�>ϻ��r%�bX�}'�ٙ�r�᫬,�Z�ND�,K��}�ND�,K�{�ͧ"X�%��}��ӑ,K��ޛ��r%�bX���NeǷ�ڑ�!�%��<�V��.�"�XP���r��B������B��֞�jm<�bX�'�~���Kı>ϻ��r%�bX���}�@�Kı=�wٴ�Kı;�gҗ�Ւۗ5356��bX�'��{�N@[ı=���6��bX�'���6��bX�'��}�ND���Aș���������G3)f���r%�bX�}����Kı=�wٴ�KlK�{�ͧ"X�%��}�siȖ%�b_=�-�/tYu��Փ��r%�`%��u�ݧ"X�%���fӑ,K��>����Kı=���6��bX�%=�߰�j��*F ����צ�5����}�ND�,K>ϻ��r%�bX���}�ND�,K���ͧ"X�%�����~�����eI��8�6�"�it��B�ؼ����Ҷ��.*�X��ISp���R@un"cZ0#��Vʙ2�L(s-����V41 4m�ˈ�](L�����J��Su���b|ۈ\Ep\��Y�yf,@mZ\��ܯ�m'z���i����%�C�'�^�H����N6�Y�[��1.�7�4]b
��z��1��[OBi������=��L�.R8�	fZ�1��0��Z)2QCK�Le%u���}$Ќi��̐�̡���Kı>����ND�,K�zo�iȖ%�b{�w��9ı,O}��6��bX�'��nd+�֥��HfMf�iȖ%�b{ߦ�6��X�%��}��ӑ,K����iȖ%�b{�w���O�S"X��N�fd�s!p��Y�M�"X�%��w���r%�bX����m9ű,Os��6��bX�'��o�iȖ%�bx{&�s��I��$�j�9İ�{�ͧ"X�%��}��ӑ,K���M�m9İ?"}���v��bX�'vR�&��ܹ�����Kı=ϻ��r%�bX	�~���r%�bX�����9ı,O}��6��bX�'�>���~��Fk�<�FS�8�s�EN��n�+jã�e\�`�K�SC)�Ƒ&H�p�{����yı,O��o��r%�bX�}���9ı,O}��6�Ȗ%�bm���W�)�r��]�h�G� L�ړ��r%�bX�}���9�I$ ��F)HĄ�d�!�da?,�N��H��I	!$D�VH��"H��e E@�t`P0`��HF0�@�%�d 1� �����I&$���! D� ����P`�$I���� �d
+#`AF$	&!JHI"AdH����B!B$�t�,��,O��|�ND�,K��fӑ,K��ޛ��rbX�%=��4�)͝+{���%9)������ND�,K����ӑ,)ș��6��bX�'����iȖ%�bS��'sT�S4KsSiȖ%�b_~���r%�bX���}�ND�,Kϵ�ݧ"X�؞���m9ĳ���OS�^o��k�i�{���%8X���}�ND�,K|ϻ��r%�bX����m9ı,K��w[ND�5�O�߾�Lm�uV]�u��)����V��z��g��sN`�Nvr�π�����}ɾn���kSiȖ%�by�w���Kı=����r%�bX����l?"�|��,K��6��bX�'���к$��7;��JrS���~��fӑ,K��>�siȖ%�b{�M�m9ı,Os��6���bdL�b~�{)�$Ւ[�����ND�,K���ٴ�Kı=���6��c �$�N���%uekY<�)*j�X�A�~%C��_�xC��۩&D�>C#�H}�h7�6�s|w�2�-P1MwLbM��I`xcg �,�G���Gz�}����83|�%�E1X�`�7d$y"�7�i-̞+�[9)� F$b؄�,�'�pH � h�({�'�n�]0��%d�J ձ��hx�K�I��[�A�� ������3y��57n���5"��)�6$��D4|#�"A'���!�H�Z8�@.ԀOc�Q�:m�>�`B#-I�����<���F1@�l������ό5	 ����=�<���a- �I�R#�R"M��hJx��k!�$��֦��!�f���6 ������6�� ��������O���CG�SJD<H��5�s��r%�bX�w���r%�bX��t�vrK��nd,ֵ�ND�,B��ޛ��r%�bX����m9ı,O}��6��bX�'��{�ND�,K���fe��.��Z��f�ӑ,K��>�siȖ%�b���m9ı,OsﻛND�,K�zo�iȖ%�b~_u�{�Yu�˫�p
��l����9nGۮ ���۱H��Dxn*��vwj"��3X�����%�b}����ND�,K����ӑ,K��ޛ��~`DȖ%��w���r%�bX���S�?f�fL�-�M�"X�%��}�siȖ%�b{�M�m9ı,O3��6��bX�'��}�N�9)�NO'�ӡ1�<��&»��"X�%��7ٴ�Kı<ϻ��r%��dL��߷�m9ı,O���f�>��%9<�8�j�&�]5�M�"X�%����nӑ,K����iȖ%�b{�{�iȖ%�@�H�A���1m��t�fӑ,K���N�2[�;!u5���]�"X�%��u�nӑ,K�����ӑ,K��ߍ�m9ı,O~�{v��bX�'{��t�&���\��Fh��I�9�Fؕ���r�ֻ6�SU����)�Y,��L�M�"X�%���w�ӑ,K��ޛ��r%�bX�}���9ı,O}��6��bX�'��%���3P�̅�kFӑ,K��ޛ��r%�bX�}���9ı,O}��6��bX�'�}�ND�,K���M��]�l�CL���rS�������nӑ,K����iȖ%�b{����Kı=���6��bX�'�w���l�S'���B����}��m9ı,O~��6��bX�'���fӑ,K���w�iȖ%�bS��^��sZ,ɚ%����Kı=����r%�bX���}�ND�,Kϵ�ݧ"X�%���fӑ,K���9'ܼ��r��J�?ܬ2`vMKa5���� L�Хy�_���Y���:���sn�E������qD��[������a�[`U�����X�̇�v���ufM����mU�&�()b�st��vA�aǶ:Qx��Z�fĠi�p�@�����Ա=�=��j��I';��%���68q�8�#s�	L����Hut�z:%�B��:8k����O��ܾ�XۘW���tm�F�҄r0[T&�����3r�b���Y۝f��Y!��kG��Kı;���ӑ,K���w�iȖ%�b{�wٴ�Kı=����Kı<�C�2v��f��i�M�"X�%����nӑ,K����iȖ%�b{�{�iȖ%�b{�M�m9H�L�bx�wy��K�B�k	5��ND�,K�{�ͧ"X�%���w�ӑ,�"G"dO��o��r%�bX����M�"X�%��a��醬�ff�f�ӑ,K�����ӑ,Kľ�Ӻ�r%�bX����m9ı,O}��6��bX�r}���?�@�bUY�O�%9(�%�ޝ�ӑ,K�����ӑ,K����iȖ%�b{���ӑ,Ky�ߣ���.p�Ri����<��%`R9lxК!Ml0�F6ؓ#A]���\ɚ˫�4k[ND�,K��ND�,K�{�ͧ"X�%��{�D�,K��N�iȖ%�b}��;�]]�F�T�.j�9ı,O}��6���6B(��!!+�S�� @���8��U�uı=�}��Kı/���bX�'�k�ݧ"X�%�~>e�;�5�SS4Ku��"X�%��{�ND�,K��N�iȖ �%�����iȖ%�b{�{ͧ"X�%����R�[1����>^����,�ӵ��zwI�$�}�}۱$D�Ͼ�n	"���{�ND�,Kϧ��p�`��D����צ�5��������Kı=���ӑ,K�����"X�%�}��u��Kı/{�fd5+qqb6�M��J�Yc�bċ�x.�.�N�e���W1%��'t�OOx� _Y`�ꚻO"X�%��߿siȖ%�b{���ӑ,Kľ���m�Kı>�]��r%�bX���aN�j�ffjf���Kı=����Kı/��w[ND�,K�u�ݧ"X�%���6��bX�'�����fj���]f�m9ı,K�~��ӑ,K���w�iȖ<� �`&��H�﻾M�"X�%��w�ӑ,K�C����_�5�]R9�Oo!y�b}�۴�Kı=����r%�bX�����r%�bX����ݧ"X�3^����>�L�]p�t�zk�^,O}��6��bX�/���6��bX�'��w�iȖ%�b}�۴�K�B�}�O��{��c�+.��.�f;Cd;��9r9�NRgV������bY��X-΍ML�-�M�"X�%��~��"X�%��u~�m9ı,O��{v��bX�'���ͧ"X�%�����!�֡uu��ִm9ı,K�O���"ؖ%����nӑ,K��߷ٴ�Kı=����Kı<��]�����\���Zf���Kı>�]��r%�bX�{��6��`ؖ'���6��bX�%���ӑ,K������s�53SX˭M�"X����o�iȖ%�b{߻�iȖ%�b_:}�m9İ8�Q��{�ͧ"X�%���^�N��l�5�Y����Kı=����Kİo�>�bX�'��}�ND�,K��fӑ,K�����j]�]�Auc�BQgd�rr�u�\Nqi��7f�#�Wj�^�XK��%���֍�"X�%�|���iȖ%�b}�wٴ�Kı>���l?��O"dK���p�r%�bX�߻�d����F��L���rS��������;Ð����,N����ND�,K����iȖ%�bw=�w[ND�)�����������ɔ�6N�|9)�D�;�w�m9ı,O{�xm9ı,N���iȖ%�b}�wٴ�K��������3rw���NK?+ȟ~���"X�%��>����"X�%����fӑ,K�ȝ���6��bX�'�㻲C3��fY�Lֵ�iȖ%�bw�_��ND�,K����߮�Ȗ%�bw����r%�bX�����r%�bX�
tH�$�H�� s�$״�f��q�S�;e�#��E��mNm�;�;-"P�s�wS����"�;�ݶ,gKk;�m���A�����S��l����1�����0]���\�t�8v���;%����E�h%t��QԙBܛm�c*�����/�l]m�מ�L��R��VlP-�e�r���h�Ж3-�tںv������x��z�nG�v��u�w?���'�0h�(��]��`��^7v��:��nZb��m��ض�rV&=�wv�vm�mqp�gw��,K��u���r%�bX�}��6��bX�'���6��bX�'���sl�zk�^������@�0kh���r%�bX�{��6��bX�'���6��bX�'������Kı>�{��'�����/'{��3@&T�7��bX�'���6��bX�'�߻siȖ%�b}�����Kı<���m9ı,O~;I����:�\��kFӑ,K��;�nm9ı,O��w6��bX�'���ͧ"X��RdN����"X�%�}��a�~��5tj��j�ӑ,KĽ���iȖ%�by����r%�bX�����r%�bX�g~�ͧ"X�%����	۬֋���6�
!e��Ƶ������͝���pSɌ`��t�5�9f3�Xc+�/Mzkŉ�w�ӑ,K��w�ӑ,K��;�nl?�"dKĿ���m9ı,J~>-��2��!��2�Fӑ,K��w�Ӑм���hڛdK���ݹ��Kı/�}�m9ı,O>��6��bX�'�������,2�Rf��ND�,K����iȖ%�bw=����K� C"dO{��6��bX�'���ӑ,K������~�k�j�C#�'�����/�~�bX�'�}�ND�,K���ND�,�ș��߮���bX��vv?�k���e4L����B�,O>��6��bX�'}��6��bX�%���ӑ,Kľw��iȖ%�����[����u��f�J�LQR�xTq�Kx�-��.�m5�2���k5�X ff��Fӑ,K��߻�iȖ%�b_;��m9ı,K�~�bX�'���ND�,K�>���SWa��u�Ѵ�Kı/���[ND�,K�߻��"X�%����"X�%���w�ӑ,Kľ��Y�grk)f��\�f����bX�%�w[ND�,K���ND������)�q6� 4X�������Kı<�߿\�r%�bX�gݲ^�֋�V�ɗ.���"X�~�����Kı?}��6��bX�'�߻siȖ%�b^��u��Kı)��/nY�:�5�&��6��bX�'}��6��bX�'�߻siȖ%�b^��u��Kı<����Kı;��y�Z�t�m)X:���3)�:͊Й�֖�R`�"P0�]X�H6Wi�5���Q�����,K��ݹ��Kı/}���r%�bX�w���r%�bX�����r3^��ק߿~��Q! 0Ԯ{�ʖ%�b^��u��Kı<����Kı;����Kı>��ۛN��^LrS��A��5�	r���r%�bX�����"X�%��~��"X�!�2'����m9ı,K����ӑ,K���W�d��m�fkWZ6��bX�'���ND�,K��ݹ��Kı<����r%�`]���z���)E��s�6��bX�'��Sw'a��Xe�]f�m9ı,O��v�ӑ,K��G�~���yı,Ow��"X�%���w��|�5�Mz~~�@r!����B���1�r��>�n��;+6�Y��6*���#\d2i��{���^��ק���ͧ"X�%��~��"X�%���w�ӑ,K��;�nm9ı,O�B��
�b�|������������Kı>����r%�bX�g~�ͧ"X�%�|���ӑ?*eL�bS���d˙��ִL�h�r%�bX����m9ı,Os�v�ӑ,Kľw��iȖ%�by�{�iȖ%����|�{Ho�,�a2�y���/ U-�O+��y�M�X�fV$�ai���wj��jڼ �lx�fV�ٕ�j������>H9ʢeeQZ֐���!��|fJ���
�a	�!O4D�.�8�T(
�Љ��(���4.�V3�VŁ�j<H1�1�#�)a
��S�m�%��'���I��X���<�<癞}�hѥm��1!�PUUPU�l���U[�L�)]���q���G7*���9��	� /m��ݕ���sg��Zݩ��v�*�/�a3��d��Z�����)�(�-�R�bL���6a�j&�'�˰LJXY�ʚ&2Oan$�\�&��T�Ler���knE=nJ�Q�R�;����������-�f �%�n�:cx���T(�� �9��W�5�Ǯܔ\�t��l�
}-n�e)	��m�11cbv�Kxn^�f��z\St#/8�m�Nza`v�b�mtf����qd��4;�  ���)Q2�C�	�T�ex1c��· PMlz"`�@�nFiUd�YhbdVG'k �n�˸a`e6�V�&ҹjv9����eu��n1`N1h9 ��Ƕ���:����J �:��!L�0�k��^���1��laD�c�R��q�l�v�&)���C+=�kvW�,�:�0��ۙ�ڂ��K�c#�x�1����VP�׳�h���z�AIZ�s
�c�6�J5��m�� ���#�T�cq�f�hi�Վ�vC�.�w;����&�sE�"�ܬ���;�̬ts��j9�z��
�C-�1+�9@�ݎ�ٞ:�m�zն+B��ui�x!�����-��A�S��<�sۖ]�m .����l�&#jċ�����¼��hכ�0g�t���7�70C]/�D�^�`{Y��ѫe4�8\�.�]p*pAKSGe&
Ls��Z�M���T�p�K�������L'lݥ�b;ueͫ�qQU!�m�ό��ӽ�^ei���e�H��:�K��v��J�Jc����6퀥T�7h�b��%Є�ܯZ�^w6T(r)vk��BgK��y�$V�p�D�N҇/Jq=l���Ns�h]uT��:R]��8@h�ܠUT�ʻUU@ۃn�שj�t�%��v���� -R�UEUR�6^*�.T'�B�@�Ҧ�6����&�ߝ�`���|�*i=>A� ���T���� �TF�� ����%PP���5�\_������{0c5��8L�]� z�1�f���"P��[�f��0�R���eK�Me�8���X٥ �5��j�Ӱ�P�\�l:��V��vFKX�� n
�LI�EIP���
G.�.;q��ll��֛E�f�K�!1a�p����<R�#"�$��F���S���D�Γ��F;�[�M��*�lVDt ��Ͷ�I?��rO.�=����1:�5��tg�f ��>�7:k�p����r�y�{m���䁢����ɕ�w�2�]��ܮW>Aվ���Öy�I"ն���ٕ�j��.�x�fVz��=**j����YI�u�E��x˲^�ٕ�w�2�{��j]�j�[�i���d��+ �ve`�!x���J)�Ct�eն� �l��;ݙX��^����[~����ʲ�����P�a3� S(Ks�	U�U�����Wn<'*��n����ٕ�j��)���$��~��g@�>�K/�ؚT��Wd/.��W3�J��>Se��2��̬l�%ۻ�����;�/ �M��}�2��̬ �d��U˩ut�J�N��� ��e`ݙX��<�6^���,��BI����7�2�we��6^�ve`[qK,�4�s:�Yom�`5�,�-!
�l�P�+�vL�R:`��s��2,����6[�7�"�>�̯UW9U���V n�]1��CVg8\�m��w���'$�Gv{+ �Oe`��x���J)�St>]������;6e`���9˲k���r, �iKV��F�"�t[�Xf̬#����T�'���긩qy�|�5E��`��mȰ	�2��̬-��K�5n�Һ\W����lsy�����9GG<���:�i�e5l�E����.��>��Mٕ�wve`�����t&���!6`veg�UT��{+ �7�x�0Dӈ����V�n��̬#�<�ݙXڊ��*�j�]�I�u���R���<z?ݙ[��LO�	���W`)����ՀM�wh�Mp�ջLM�f�`�2��2����Uv��/��p�3bpu!���°��#����)7,��d6kDx�%\�u�n^��r����e`6e`���%���V��[�
m�n�`�2�ԑ�I�E����e`T�h
Q�|��E�n��lx��x�L��fV6S ���Wi]7t�m�yK�z�	��Vٳ+ �Vǀv�\J���S�w�od��=\��{��(�����w��$���ot�Rj(�e*�:��u���X�K�q�Ő�X��tڌ+�q��Bv���fcu���T@nL���Ι� =�}���
fjpqYZ�,D8�J����Aՠ���gQq��)�V-��M�;�5�Ƙ����I�$�h�l�6�<5Æ���d��fuV7u�������7��7Y�dN2F7��e����51&��tŊm��>Χ�9�5�uv�YT�A��f��� cZ��������+�ة4e�6��lr����>�2����]��	�2��T&���O��'m����^;&Vٳ+ ;ݵwj+e�X�ݦ&���^;�+�RSc�Gv< ��#�5E%i��wr�	6e`��]��	��T�En؄&軷Xf̬#���/ ��+ ��g��0�nb��musRq�#ù�����tv��gVb��sۭ׬��\fv� �� 7�7fW�� 鱗�߿$�U��ź.���_�}��䪮w���9ª��%���;6e`��U�r�#k@/֩xN�l|����{+ �d��RQ��ۑ`��Kj�V���`z�ʪ�R��}X����;�"�&���>ݡP�]]]����v�`��ۑ`ve`�2�ӓ����P(L�1t��u��6&�]4c���$.��j<�nmT�����c�v�����Mٕ�wd��";#��Z]"�V\��i���Mٕ��W+�=���y�ۑ`H�"�v픒V�Wn��XGdxmp�h`#`� �`,M�}����ﲰ	Ru-U�������`��ۑ`ve`�2���q�դ�]�����ul��Mٕ�wd��";#�
��ԷJ�:�U�F!�˚���;c\>�}~�lٵ6�vX,�	X�VT"1���t�m��m[������;�e`��[%��� #j�
���u�wd��";#�:�K�&���>ݡP�t_.�'m��ղ^7fVݓ+ 7�i+����c�v��xV�xݙXvL�����m  X
!>��[��ϋ��̶�rʲ��w�Mٕ�~�r��{�W����ݹ;%�YV�ui�V<���Z3��yb�F�܀�z�2@�s[t��[�V]�&�*�V軷XvL�#�ݹ;�+ �*QN�I7��)[m�ݏ �6^;�+ ٳ+ �l�wIv[wLv��l�wfV�fVݏ �t�wQ�����5n�	ݙX͙XGv<s��S�� ��)��%B�����6l��";��͏ �ٕ�}��yÜ�s�*�r� t�������A�Lkc^8���>;�� ��&[mY�c6���% ����u�2&��}>��%��B�-�֬]�<X��y�tB��4x��:S����A��wg	�X�g��Ȯ[��Ng��]lt8Zm/7b�H,N��4�i�QنiH@��j��m�WKn�{���8�q��9����ـ�lV|�`˫n�Mf��D�sxo�e���	N.�٘3���t����7Q���{1,�2��Xa�b�g�"7c��;�+ ٳ+ ;ݴ�Ի�ջLM� ٱ��2��2�Wv< 쥥�F���L��]��N���6l��	]��fǀM.Z�Pv�(h�Eݺ�6l��	]��fǀN���>�R�������� %wc��;�+ ٳ+ �I��Z�F���E�P���&`�yI@����c;a���4�*�rq��b]2�2�����+ ٳ+ 'I����KCWm����n��ϩ���d O!�(� �7 I�l� �@��(����}��`�ǀ6<B���#j��U�m7X͙X:H�fǀn���;�)SUt]0�v'm� N�< ٱ��2��2�{��u��:�n���5M��z�\�{��	�� �$x�\�������J�ӧb��r�]�8�{�;�p�n��q8i�`��'9R��M��ӵWj��{+ ٳ+ 'I odx�r�ܺm��7Eݺ�;6e`�#�� �ٕ�w�)P芒n�h�m�X+�< �>�[���	�
V'��X�0��%eiF,�����0&1*@`� �VH�!`FL�i���ߖ��莳Q�"Aaii���h@�̖"�b "I�JB� H��Jn��b@]k*\ ���wXN#��$&����Uəs`�o�5����krL
d��&C����<��%�)�b���y ��d"�I�\V�$]�⍉�	H���a0ӱ7� 졊���^q#!sZFd��xL��D!@�R`F%H�)l���Hc!%�RY��X�fcX���H�IX�,�u--H�JR����K)#tTJ�	J���2��A�RH1 �1 @#
0�%�q�؄�*��M�p�`CV�����=����eh-4'��D�1B4&�A8�)���| �*lQC����AX*x{�Wb�����nI��� �2�&:.�n�b��=UIM���=��vl��";#�;]R��hwv�|e�x�̬�fVݏ 7�<�Cm%J�5at���J�v͋S�Nl�ZARVLД�a�rSSv��R���LA�� Jձ�_����";���G�N���7jR��⺻�����	�c��UT�M��6{+ �ٕ���.ȭ&��ջv�� odx�fVٳ+ 'M� ;)R�Ƙ�ZJ��7�2�͙X:lx(�Q�$D�	�Q�Ab>��A��+"�#J�RFI�1rr����熾�o����l΀vlx:lx���ݙXdS��m�
�Ѩ�Y��F[�sr;�3nv{!�b����@�X0l*�m��o 'M� 6lx�fV l��	/Wd�Yv[wmR��fǀN���� J�Ǟ�U$mhZ�w���i��m��� ٱ���x�c�5E��E�i!%wlm��fV N� l��=ʥ6{��6W�SUg��qҵjݷX:lx��OO?��=��'�{���8>7E�B+�� ȇ��M� ^�Sƚ#*�-T9�ni��J̛�<6���a���0A�Yx�q�i]�#�E�8�K`-B \O/x����W1��k��<v�tpKJ�H�/!+XKˍ4��"m�+��1k�-m��,�Vg3N�e��o٭B�5,��tj�����cj�svDL�)��[�Vl�-F1��eך
��@,�mܠ�̋I�N��$�O�;�o@�L�2�̀�Xi�IT:�K�y�{���F,u\2��)���$ˡl��۴6�wc�7�2��2�UUʯ��y���.O4�t�2˵v��ٕ�lٕ��ǀ6<t�i��4Ю�`6e`���Ur�'��6{+Ԧ��
���c�n�`}Iz�y����	ݙX�2�	R�pWe�m��� �#�'d��6I��M� ���%�)+|C�u�Hk��͋S]��+(\]��.��ۆۉA�M.�-E�ez�=���l�+ &��ϐ���6Z�H��n�(V&6� �&Vs*�9Ó�+ �r�Z ���2�HʴU-V��!)\��b���",�-*@-P�*6� TVj ��!Y# Da�\��XA"a�a�H�$��ʮr�a�� N�xݙX�R�;�K�\t�Z�m� N�< �#�7ve`$���mdV��unݢ���r��\R��^$�V�L� �$x�Ilwt:v�˶� �ٕ�l�+ 'I�Ix�Nciݖ�\��c]`��6M8[n۫v����vx�=���1�	X�P�]f�\�#.��}�+ 'I�Ix�̬v�,P�m%Vݺ�	�G�$x�̬d�X�g6�EګV�m� �#�7vea|��(�TUUr�#���T�I��I��A0�j!&7�[o �ٕ�l�+ 'I l��	-K�RR���ZLm��fV�R����zy��2�GV���j������MJo5�9Hq��n�sګu`�F�:�CFY����e�\� ���\ ٱ��2��2���E����7n�m�͏ 7v<d�X:H��J��n�2��ݷ���L� �$x�G�I��wj+���m�m�$��	�G�$���~�O2	���!Ȓ-�ĨPZ0��Ȕ�qX�����#�V%Gk���h�i��	�G�$x�̬d�X�T�y]����6��c]���h��`����f���8��]V��w �%o5�0�J����{� �ٕ�l�+ 'I�t"��Z�I���n�ݙXwfV N�<�^Ns�v�Tz����t��=��[������7w�Xݭ�N�uw�Wj��n�t��-��ݙXwfV w�h��ipv:nݢ��>[%��2��̬ �$x�+�EJ
�)H����XL3�ֵ��L�e�[ѭ!Jۋ V�c�]6�p�i�d \P׋0Z�Ҷ����	����=qO-�!8��`�Y�v'8穌m�ܶ��2e1j��#l�Z8ɛ�Si9<���k���rh��&ÛX��0ݝi	H#�n���)��4���j��6ұ�vz�	βg�8�]��ȞA��t���2�m�+`�v��!q�&����{S> �;�+BY�t�{8�v�F����@L�fh���mS�E�E�th��:���۾���+ ����	�G�|�K�$�Ĭ"�m�N��v� ����	�G�|�K�7veg�č�y��G�ۡ�m7X�=�|�K�7ve`ݙX�z�K+�b�i�6�=��+��۞��g���̬ �6<��EI�I��m7x�fV�ٕ��ǀ|�K�"U�ӱ	�dp@�ʍ!˥I�xXi����˴j��A
�i�i�H�N���ZM�� ����	�c�>[%�ݙXݭ�I�(��N���ֵ�rI��ߵ���@"b�_d��ٕ�wve`�mW-.�tݻE��|�K�7�2��r�-��X�'� })V�n��VRlm���s�~����'��+ 'M� �l��I���DWm�)�b�u�wve`��-���̬�9UUS}^�+��:V�]f��:Y�X2�f��0q9�ln���X�oj��S,0�f������|�%�ݙXwfV+oW"/�X�մ����|������{߲�O~��	�G�}]	�I��m�x�̬�=�f�<x�+A1B�!��bJ�C�@��J�[4�)�l!��nLF�������{�nI�s��"�*E
����۬{�+ 'I��� �ٕ�wkiRw
��+��m�X+�<�s��O_�zOe`ݙX�Y���۴�)*Ulb�
q[Ir8A|]�%�k�<ROvJ�=nm)�)3��E�tݻ�m�)��	�2��̯� =[�<��B�Yn��VRm��xݙY��\H���X��y�ݏ=\�q"z vQ��E0l��X����	]��fǀMٕ�l�tYv[t]���`����c�&���ƈT%�0+�Ͻ�|7$��c+�w�v*�m+t�xٱ�ve`�2�Wdx��b��ݎ�]+I�V�D�wgK�WXHC���jm&;(k���*	���Zi$�|v��=��Nɕ��#���>@zO<R�{��+b۬vL� �� M��	�2�ܩi���Z�?A�m��^�~�~z7c����)/l�V {g� ov�ur�*X�wJ��	ݏ �ٕ���T��O<��B�*�EL�ۻ����X;����� TC�>ޡw�pi�CQk䬑��F�#�ɚ�u�}�F0�0C�	=�����N{� �u�bI��bkHK���P�$����#,##iD_Ci�42�i��Dhh��m3��ᚋ��IhH�)���6�z'�]�|&��洺�)��	�=�_wy�W�#�pY�HyƲ$"�sZ���,�\��_{p�p����r��9S�̧T]PI�A͇��mz%
Q��l%�y��r����C�t�%Y�y!�d$#P�� T��˓���'���$�L����� ���T��|���-i<}g��&�ÈCp�ޥ��0�)+V� ����,��ID�UUcPhi٪�����+lm�8�v��".�C�T̪�A��3F�E���é����[\�ʖ�%�����:;M����h�d:3�r��Kb�;4ڠ� �H�*`v�h��m�Z,3v�;h�KI�Y:��E��,��5-F�p�r�N&�`;g؍$�� &ka�mc��z*<�����9�+��X�5�zͅ��n��[v����mI�d�:9݋
Х���9�������6�kD�]!k���g�&����:��-sFI@�2�l)��S4��������@Il,���6]���6R1�N�v�VV/!����|��k]�iE��X�4	���E��E�0�-�\i��M�e ���F�U�۳�^dLv����	���d.�H�x�0�D���9��q�MF-��;�p���-r�nݭȏ�,�yJiqmŭ�M���tx���l���<�|̦����Zu�Բ:8��4�����^۲�.ރ[��iAp�����Ui���I�$�d�;��,�;U��w�v,W%�:���F��g���ej]��j9�!M��(�`����ֱ��-8�օ��GR�-�<�lyp�������v�F:��^�0�+u�]��(�zlGM�W���t�`�0D%�A�elJgC.u��\�k���i
����ػ��6̔eU�.�4x�:by��WRj��6,� r������\nC��D����٪�]�^_m=����]qk�q�vɑRv\���+VaN-����&2���)���,4TK��6�.aVV�j52���.^l9�q�Z�L��Cvs�5T����݂�P�n��g"���b(�oX� ��cL�u�j��T����dr��(�%��T��*3Y�Y\��ic]['l���T�u�rU\����U�Ͷ�{<�e�l�b�Z�SW����@iI�,�kv����-��B�#�(*���:�:��ΝӺK�9���D`���z�G�b)�|�)����������*��?��vd��fkZ�k%��4-kG�L�`�bd��ܶ�;����D��v����yb�Pٚ�Ă�hY��q΋����wZ��<��y݀nȅh՛����z<��#<u�x5�����LJV��3u�j2˂�r;���3�o7l�Ɍ�%Od,=��d��ŗ��^V�tEM�ў=�7�۞m�Mt�x�����Ņ�mQM(U3	ӾN��M��P��`���W-�ٵ\���vx��<!�9�Zӵp%�����х�D�E0m+�Xٱ���� �d��$��v���t1��v� mnǀ�<�&V7fV�#!V��v]nպM� ���M�Xz��Ľ'��i<���A>�I1��oԻ'���{+ 7�ǀ�<R�A#I�lE��`ve`�s��O?�=���>ݙX�\�6?zЋ�L�%%l\h�5.�\K�
,ke���S$��R3.	�:1��V{m��y�� �ve{��W�='���.�K����L� ��}{����WUR�r�bܙXݙX�6<�(�D�V�6ݶ��fV7fV oM� ��/ �RvUܷm��I���`�2�zlx[���fV6�bhT�ۢ�%V�u��c�=��9^�=�=��Nɕ�|�����ٮ�G�x��J�Ͷ��7^ ���L+���c�'����p�\��Cg\�^������fV;&W���W�	���;Zy>�m_m�����'d����n��"��6P��2�n�	�2�zlxm2��\W
�9EIHH���20$1S�)E'׀}�2����;��J��[m��U��q)���<���n̬vL� ��V�P���1ջi� M���\0	�2�zlx�)�\>��N)�rP�� ��cFXiJ�k1���FZP���I�*��b.n^�����'d��������=�,/��l����`�eg�U�H&�� ='�����&���Ip��%i*��� ��ǀE�/ �l��'d��6�5P��wV�.�V�6��e�Mp�'d������W*��W)�x��*'�PI6���� �l��'d����x]�x�Cm%DM�:CBUY[�͌iFn�C:�0#c�j�@�ƶ�}�r�n�J�ڶ�����e`�v<.��+ ���)����Wv]�n�Gv<.��+ �ٕ��h��Z�N����.��+�{g����xR��J��Î�j��Mp�'ve`��x]�x�MW-��Щ�v�0	ݙX��T�g��yl��Mp�s��TWv�C�ZM�1�-�M��Zb6��ɻ�t-��dc�=���h�l�%�#�(��T��6V�c�sڅ;&6te_m/�0���zn�ִ>Q3n���C�N�-��yk�ヱ�k��-2���v �u��=��:�ktGb$�W�P�	e��,��jZ��mc��t����vtr�VLa�ګ�SS'^��8x��m��JYV:I9���H8y���3<)�)�lXX�Ic,�tx޼�>�œ��mlk��q �-��v����L�?�����|�v^�ٕ�N���6�5-�wE���bm��ǀ}6e`�2�Gv<�\�s��ò�^I&����;��`�2�Gv<.�e�E)�J�ڶ���̬�$Dl��<�z���`�Z	�-�ݗm۬Qݏ ��/ �k�;�+ �N�?g��E�Ɗ�<5�4�:��Z<n�v�*��mh�{	�1N��q&[n��7c��[=x�\0	ݙ^��W�"6y�z�<�����-�w�}5ɾ&*X�Paj��m��+�ȐJ��E�Yj$U*@� �⸇*�M���"6G�M� ٩ݥr��B�m�l�7�2��ݗ��_˳{��7��� �Z�.A&�%bUm[�iwe��c�>��ove`[���j�
�WM7x���W}3��M���6�v^�Q��qJ-�ګ���)g��]E���+�W���4j8;;/�)I�BM$�W��}6e`ݙX�v< �lxTEl����m7X�fV{�H�$����	�2��kJ���hWv]�n����I9��ksF	 9�f'���� 'Q7��{�rN��vnI=���"��cc������Ļ���=��X{�+ ��ǀ(��*)�.�&�;�+ �ve`��x�d~[~�����D�`KE�i�\F֦�-�!5�Zh���Ԗ���PhƊ��N]�:�˶۵@��v��7g��Wv< ��<wfV�+n�r	�v�[V� %wc�׫��+�v�[�=��w�遵�5*�t:��m�N�o >� ���ٕ����W@��j�ЛW�m��ꪪ�R��}Xｕ��#�*)����y��ܓ߲�'��.��r���u�w�e`���[��	�2ym����ZƣH�/(�F�) �K-��^YGmT�X�&�V�M�i�����tg�v��Ҵ��e�v��V�� ջ/ ��+�r�������	�$�ɫN�M�T�x��xݙX�L� ��~�9Iz��^Tq�.������X�L� ���v^�$�+���T	�7n�?s�]���`�}����������]й��7B��ڷX+�< ���͙X�L�j�\�(Ԥ.;���C6�P4tQ)��cl��n��)qh�a�k@�C:�ͻ(�YJ��7>�Zu�sT��n�R�[.:y��n�:�XD[����2�5�ˉ��ݭ![a��!E��U��bR���N2���qL[sd%9r�5-ͺ�g�g_}��ͻ��s�%���8	��6��M�RF5�݊֫Hc,T6�a�c��Mb��wI󤗺wtF����J[z�-I���9Ƭ�@Ԍ��ƶ�����(��=��k��j�Ҷ�����2���_�r��U]����=�M��,�Ѻ�H��ɳ+ �I��j;#�5n���\�r�"z����t�պ�;�{+ �vG�����]�{߯ ���+ ��D�N[J�J՗m۬ �� ջ/ �ٕ�Nɕ��R����c��M� �#�=\�O}_����k�<���sD���F^܂�'Q�ůUk�������6�J�Y[4�x��&̬�L� �� 7dxȓ.�z�]`T\�t=��βrNB���H(A���@�)���eUUr�԰=S�< ���ٳ+ ��K�!t���ڷX�� M���2��2���%J���"ݫ�J����W+�������O����I&V mvG�}�*֪J��V��2��fV6L�Q� M����UR�Ea�K�K��pP���t$ҩ��j$f×Z
�,4a6�Z`�-J��-4h�����e`���l� �ٕ�v�D�U-��Z�յn�Gdx�#�;6e`�e`��.�mX�lv1[x�#�;6eau��qQT*��re�SSRA1���)JBT���CXj���-J���2ZjS+���jF6!9N?y%���!Pa��<+Ȟ�YN���7��ic.�n�!20�(I��b������X[�vj�CV%`�RVRB���U4jˣZ!��I�h��!�8��70�3RZd1��h\!&A�d(@դ�+6h1�!�Ɂ�L���XI�[HV_19���f��)e!G�\�4T������� ��4��E��b �| �@ڸx � _P�z�� pP�M!��Qv�� {��(%WC��X�lxR��(�aN��m��fV�L�Q� l��"\uwݫT	�۷X�2�{%� �#�7�2�	�UҬ��&�V��@���$��cv֚����<mf:�\mb�y�eիL�MЭ*��� odx�#�;6e`�e`́��	:�j���ٳ+ �+ 7�<�V�B��������fV�d��� ;�����Av15n��L� ������/�b�EpZD��E7>���p���a��f�[��%n�`�G��ǀvl��>�:���q���Il�Y����4i���430��u�Yf�&��T�[�K�-&W\�N��m+o ;�ٳ+ �d��� +z(D�)�:��ݶ�͙[����ݛ�O��u�$��~��(�Q=�EߒvZ���ݺ�=�{+ 7�<=I���7��X��V
�`��ZUn����� =��vl��$ٕ�o6�EF�Hi��V� I��O�'���9$�~���'�}��$&���X��`��	���&�0�j9���j���o �y�qqc�׋&��Q��$��㫏��
�Ȗ܃�L�����O< �'��I�-�Z͹��ckc�i2s�ћs]C=�7�x�3@[he��+�/ic:�gqs]���ۄ���Hss(�68�R�e�@�!qX���r���o��h~�l5@��8h^��
��m:݆T}ȽFy��,\VN��;��:��kj��]�N[�#fk��%Ƀ�&o=&�sY�-�4�3l(VҥMtwU���~���2�{#��<e�D�i$:�i��u�l�+ 7�< ݑ��2�ԭC���e�j�+��`�G�l� �ٕ�wd��	ݴ]�,v����m�~���R[=�o����X����J�ȘS�6��l��ٕ�� }�+�Z�t�u��>\�f"8Ǣ������N�bn@֭�qCC`v`^���=m���2�{#�����Ur�A���j��j��V�f���=����9'����qUs*���ܑ�K�`�2��Ԩ����	�WM[x�����a�%�����y��r�K��WN��m�{�W=���	�߲����G�Ii%�i]�e�m`�2����G�wob�'oe�v\ۛ�/��'���E@W��l��C #�uX�U��i?��$���@�7~l����G�jݗ�vl��ݰ���6�������?r�"�׀o����#�q#�t��g���]P��m�l���ea���W9��(�9�D���	=6U��%uue&4����s��-���`}<�vG�jݗ�T�-%&�E��i���� �U#dx��xd�X�T��ն��u��Wn���N��6�	���U�4{:�e"L�W<Ąca+Ɩ�4� ���^��d��&V vH��
�*]'eӾ1[x�����F�{+ 7����=ď/ �ui]���� �=���< �dx���Ԩ����V������ܮU%��� v{� ���f����� ��M}�s�����Rc��6;b�����[%��̬ ��H�Ji��5t�|����<�Z�P[E����4������ ��˒���M4A�c�z��ﻠy�ٕ�I }�6U�w-]]���V���X;��{#�"����V�|�MІ���u�� }��R^[=xｕ�NJ�K8Г]5m�{#�"���;�2�=I{g�4
����v];���Eݗ�z�g������ >� �r��\9G9�B0R ��i��.�°Yi�2B]+��ղ�{������{g��Z�!B�Äܥ����y7ޒ�B�̓�Xq3���(�gb�5���UL4���d�m����h�*Q�чux��vHJ�Lg�Rch��lK6��%E��:J�A\��28w��\J��lY��km��<�4����yzj�,���)�k`2@Q�	��쓕e�`%��U-#-�="�Z���:�,���<e#].��ݯ����ChI���v���ۿ��߲�	��vG��W�<��x׫���C�V�����u�M��Us�H;���<��x{&V oV�vJLwWI��M�����e��X�p�'n�
R"�auC�m��E�^�ɕ�M�����5eڸݗV!���xf̬lp�� �d��)�lHV�θ�%[CT	����F+4pd�Wt�rkbP����К
�F�3�yﯦ odx���fV9*E,�BLuc�f ody�g9��ʧUT�X��$��>�ឮ$n�V���ui�;���E�z�	�2��� 'dxQ);)]���ۼn̬�8`�Ԥs� �y/c�۲��i6���0l� ��l�^[s�O����vmL�2��(�46F6Pe�+�F��]�z]�/6������ln�������ذ	�ev�A6:`j�
ݨ.0����m��с����7��dx���K�]ZM:I�x�2��p�UUNWpXA&ȵID	�á �'5�x��X�M� &豦4&���� &�����qz{�V�mxqgc��0�%���O{<|��V�8`v����M��6�h܋�o+W�1���$f�%��[68�G�$���@b��L���j��#��&V�8`RK�"��R�ue�wl�m��&V�8`[%�/b�s�H�佉ӷe+.Ҷ��z?�#�6\� �L� �V�vJ��tU�7Bl�	$x��x�2�=�.W$�$��w�s���H�!��z[��	6e`�� 6lx�چSl�k��j9�!�]��@��ǬF֦�L�96��i.c6i��!�p�}�f̬w\0f���+��l~0�%A^��lcI۬�\0fǀoc��fV9*)�`��ӻf l���p�6l��&��m�Դ��;V�;0�2�	��j�/ � �)՗eݲ�ـlٕ�M�T�x�p�7�!.e�+e�~�'2���p��6� ����=$�⻃�w�aJ]���!	)��Ie%<�s69��h�z٘��YV����Gjo^! ��l��=�h�<�&>�y�
O7���i�S<��:�+!�d�*�	��)5��ߞFi5[�	���| z���}}" F A�B{���>a+N��B�g	}Qa�gr��,RŊL�O#7����C��Ҹkɼ����xl��2Ȼ�@�C�I�b�5�J�o���I��Ğ�
��HS��*b�c�+��T�Z������X��!9�[(,X����|�w[=�5��
����\��5��mH"Z`s��)��t�.�>��D�%Ѱ��}xzd�(����=���� �=&�NL8Bq'$��0Hr&oN�n.%ٰ5&CTy���@g�������Ts
&[��ny����;`C�uW^dE�Pɋ��q7�4M)� ��!HD�
����^�s(V��l��(k^������J��>sӞrR/����6B�a�+.�K��D�i*���10`ɫЉ,�Yy���s�s3Yy�l�g5�O�m|���o�*�P(�����*�U�R�i檪��U	r��ckA��ε¹���ʫ+mB.Xwf��6C���&Nݦ`K����1�)C�\G#Q� ���f���[��vߪM}z-һre�t���iwd�������2�ãA�\��V�z�RKt���:-�gF�Cj3D���9��)1���F&yrbi\"[++��ز�T�-��Á�A�D�ۭ��pZ��Ku=bd�^ݱ�c�Qx����=�4u�����1ۥ�M����I�j�C�-Q`$(SmX��z�x+z-7h23C3��g �u� UW\��K�C6q,�΂��Aut�����s�xԅ rQ�[�\)z8m�u��!�X�f��� ��KcE�켽�����G$�p�����#���9�sv���y�r�η��:[�/#e0�iX+	��5���G`�!|	��7�'ԝ�i4	"F��v�&�J��G2pf�2fŒ��J��a�j�<�Ӱ��U��T�b��⽩�Z�����jͺ�'���y+k�5M��&B9��:�U��k,"���(҆������q�Qu�j,��B�ad�X:Ь$ؓcs��m�&����fTA��Xs/0�[r�,@��Z��M6n�4�^���i�:#r6c�/#�؋nq���e"nȔu9�1�5J�pE%���t�6)�D��C�����l^C�s�F�MB�\=��v;Lm ���`g�a4F𤺢为���!D��UJ��[סlե�h��[f[��c�����ճ=J�괝����vuInI�q���
�87�>�:1n�R��J��Z��.u�@��qm�D-��ʎ0h��������%`�)V�jmiH���V���LX�*�Τ�|�1k7� ��<�ͱ�LδiP��ϑR�U业�>��%zW����*�U��j��.,lI)�ͳU���˒��uj��j��Z��cA����2��!Y@^���I� ��:����TT�>�;��"�8'�~UF"b��PCh����t�QS�pbI�$���_�Z0m��qw'̶��Ş�V)� �՜Ŝv\�m=rJѷq���E�[7)�Gj4�!�u�P��t5�x�\�2�H\ā��,�Aڲ�BK������q/a5����瞱���D�+{:�KU��q���b���x$�x˭���!f !�u�����n��D��´2JDjK��Xţ3��a)pU1�/�rI	'���$��>S��B�"%(�c(�S@�(���1���jmjw�;:ہ��6�a�t��J˴�ۨ�� �$�vL�d�X�[B��wN���ě0�"�'d��6I��M���ꨠU:����͙X�2��p�5I/ �ԥI0��Ri�6� �&V�0RK�;6e`ջE�@M�V��u�l�eȰ�2��e`dE��%o�*�C�j��[��\#�B�$���a�ۃ���
�,�qۀ-�ؐ�ڻf I#�6l��$�+ ٮ�^���`��o[�{��l߿�#�kM�j/�@NG�?o�훒w���7$�}�������U����]���`��V�\0M� ٳ+ �e!	˶��Wwi����������fV�����V wW�]z�]��	� &�x�2�	ݙX��|�l�vƛ�-R4���b3Bͩp<��!s-l.�Y	��I�d%Gh�a��#4�������vL�Mp�W*�A�'� �� N���\IZ|J��$ٕ��)#ޏ�����$���URA+ҭ�&����f��;��rO�����^�������c�~���X�k@��wB��wl���{�fV��(�K�;V���j��7u� �&V;0I�ur�����X����[
�˱�Mn�)��n��x4nl;\*���Ě�t�:Uwb�e�� �L�w\0RK�"���;ݤ!5-�����6�����Ix��vL�V��WR�����&��d���/ �ɕ�}���V���
�
�'m`]���X{0>�*꫇)lP B�" ؈���}��s;�O���T�(��q%iЮ��;�e`�p�;�"��G�w�*�w��œ���@��f�S�QTG�5muo*�4y0H�86��qj	n�c���Ȱ����e`���v*i�i]� ݹ~�H7g�������`ЫZ.(�[���N���ǀvI��}5� ղ^!i�r�.���o �ٕ�vG{r, ݑ��E$�-�����2۬�8`�ȰvG�w�e`��_��	/	x���Hi�b
�b�n����u�<;�Mp�q�p�Nz��ͮ����i� ����\��X������4#v��3�Z�kM�Dڃ��=����0K�h3c�	
ҙ\ՃT��
�F�q�\�s�� ,��s��*��;7	�nu�<�h��lAR�m��v���ѵ�ӓ�S�r�2���:�Jq�0�K)1��,v�V�}I�O9�rI9�O�1p��Iv�B� �#e�%դMY��s�6�LvF�s�t�!l���2��	��=�� l���X����J�@�*�����<��RFｕ�o��`�ȳ�H��&]՞��HE�E�o ������X�`�ذk�`���Ҥ����>ۑ`��un���+����}X��(<�V�ۦ�&����v^����>ۑ`��i4;.�R���չ�w�[�@�Xs��jY]y�����G�����U�.&���e�]ۯ���y`n̬mȰ�fV�-R�J�]�i�������\����8�.�,�fV6�X騦�D��]ݧn�`nE�}�2��\�K���vOe`�-���6��[��k �ob�&܋ �ve`nE��!*P0���0	�"�=UʮvO}_�~��>�p�=�}=Ӹ�Ι�Ů�]ef��r��lո3ˬgWVx��vʡ�5�y�8p����Wm��+ �r,�{6�X�ݺ(+m*Lm!۬mȰ�ذ	�"�>�2��I)bh�N��m`�ذ	�"�s�H��W*�0H*`������rO�Ͼ��p���\Q��V��l�&�ŀ}6e`�"��W*�ٞ0��J�K΋�V$�]��}6e`�"�7�2�	��`_~��ۛu�K)qf�1�\�}*{w�n۫�2fu؜n:�[87!`����cn�	ۑ`�p�&���Us���{+ �R�����j��m[m`�2���8��~��6Oe`nE�Њ 衇.��u�M�����&܋ �ve`MUݒ�P�:N�XQE�{�xnI߳���s�u�ܜ<W�& �|���}מM�'���S�5�iX�I۬mȰ����}��g@��<ߧ���T��Z�YLա˘%�,��a�!2�A�.��s����WZT�c�M����68`I2�	�"�;[V-/��/�� �0��^�W�=/�X�<�ܤ�hZA��:LV�cf�{�Xۑ`��`c�4�SJ	SbUwv�۬mȰ	5� �&V��ʪ^�g� إ�u�6���M�m��M�lp�'c�6�X�G9\
�8A ��a	##$"��r����Ҟ��l��.-W��u��Aã�Mɐ�#(� �`���K�� ��hⳂtj囨�14�(�e@���X<�۲w̫�8,TWD��i��M��kIt�K���ɂŉ4[B�!�4�HܖV��`���B��F�+cc(]\)l��ר(#l�5`J�C\Ѐ�"	b�S2��Q�����yVǶ��YA���[�i�L� �A�թ����9<</�ȉ�X�3�%j�&J��jݛ`�ۄ���+Ng7	�`����F6���.�M���e`�� �r,n�`i�w�_��+M�;0	ۑ`u� ��+ ;]U-۶��ۻI� ��7\0	�2�	��}*"�s,`�m��m`~^��V��v8`�"�>�ժ[|*]�.�[f7\0	��N܋ �}}:g��_����jݣ��FQ��QԮ��r�yB���]<Ir�n�=���M�t��$�]��$���V�ތ]��އ����%Wwi�ـN܋>�9EUVs��UU�8�E$�n�w�rZ{}���+�fb�+z�޿�-�x�Ȱ	ۑ`hKH�� ��i� �v^;r,v�X�)zL�O�j��Uv�+n�	ۑ`nE�M�-���R�o&�^��N&��1��s�m�ذ��p�@��5�t0Fh'��[�&)uht�L}�mȰ	��E�_������� +�YLI��M�n�`l��N܋ �r,��Zۻ*�;v�WT�� �d�v�XG�U̬�\���WN��?^�x�J�CC��ff�0f���X�}C��x+|����P�6��4D��T$��E�"e�
c��t�#Y>��鹱�D�!T�p`Kڂy�JNL���p��K���e��T�ִrx��N�1!�2_-���M��4�)�m���@�AѢ��!���]�.� ��!]�!�`aX�7�P$�8��(�$�d͆�a4dc�!��)��0���Df���#��m�A�G6M��pKF�BEd~Pڜ�&`��df(L��@�|�hA�T�*L�)"�cRE'��GA��Gv@���##<�l��4+r�����l�=9�J���!%2a�.�.D��-�lSb`|����>砠����*/��Gh+�"!�t����������<��}7$�ɑPJ��1�;M��\0	�"�6k����s޼i�SK�V�*��Tݳ �r,�܇�$���I%�s��@>ݏK�ms�m�B���"�htQ����/\�5��M��jP��΅���32��}��=��^�����{�\�+������I$�@��,��H��V���%p�I%ݙ�I)w%� �w��} ;o�&�HMLl��v$��̇�$����IwfC�J(�~ ���C����Θ[�۽3r�|���9�m����n��\H&"�(\�TX�@2+R,0��b�� �_o����$�^@W��:�cv��Ē]ِ�䒊8^$��̇�$����Iz�����>���vj!���`�B 	���J�Kv�ѶNW�:i���C����C�gz�^^~/IwfC�J]�w�r��봖�g��I/B�@�΄��;M��$��!���r�Wv�w�]�H[=�>�$���y�s����߯���6e��b-�>I/]��x�K�2|�QGĒ]��o��|k���V3)���?s��]���>�$���^$��̇�$����;�o�fx�����O���K�2|�R�e�$��̇�$�*�r�ïw�'�k}q0L�k��a����Xu1tr�j͘�:����˭tn��>9���8�������A[-�L�\�a��A��g
C%������R�e��]�S.�d�#��ڹF(�q�,Z�Oo]��eu��v���sȺ��cN�,�yF�i�M�%�+6��(qZv�z�_�W�q(Y4�68wid�ʬ�1�� ��3��G{��~{�)��L噵�	�$`0�6v
�,)-�v�\��҇]�F{8-ų�D�h�ܭ]�I[�Ē[=�>�$��˼I%ݙ/��t��M� {>j�\�0��J]�W�Iwd���$�ٕx�K�3���9'6��t����fR
����	l����BR�e��K�2|�Q^�x$�'�b�*-[�i��>�x]ِ�䒗{.�$���}�IM,T��MqZ홼 ?��;}��}ݼ-ِ�䒋fU�I-�֠�V4����)`.U�ͩmm��mq��G9�Ѻ�vm�����cqe�v̰����@;���Iṅ�$�[2�IvL��$�U�#vܫ	�������������		� �$B@$H�=E���~��y7m��}��9e�f��x ����g�Y����@:}2�II2�Il��{�˻���>�$^��n_�`�`b�����nII'���%�&Y�$�ջbW	�j���-�������}�o��[re��Jvd>�$�\���-�	�#����X���ٺ����(���Yw:[H�� ��-�fe �5٧���g�%�L�ĒS������KI})�.�t�-��[g�$��2�II��I#c�ĒRnC�Kab�r�Bj������I)7!��$lpx��� �fy�����~�fn�o��:Y}�e�رپ�~��� }�Ⱦ�$�lʼI%ٹ�$����Wv�32�*x }�����~�{��}-��|�K�Ʊ$���v���,O�k˧����L�k�^k�v1۷.�YƷ���%�]D���B�{������IvnC�Iv8�$�޹�$���t���6�:� w�;}� ���� �w��@>�w�| �O�n�:�v7uvٟ$����$��d��I-[2���܇�$�*"�s,t�'n��X�Ko�_�$��̳IvnC�Eq�� �#��(��W�}��m�|j�3
teu��.w��}��� ~�>��^�$����I%��/�K��W+��U��1,IKc��%��+�(c����'`�M�;a�4f�;k�W\f�vq�W\q�!N�-��|�[{2�I%��/ܪ�m%��e� ��� �2��رپ����cIo\��K��F$��܇�{��9wh/��߭vͳ3-L��ߞ�=�ݙ��$���}�Iv�e��IT�+cI���Rg�$��r�g�F$���<}�Iv�e��K�܇�$���]"&ʶR��1[F$���!��%�ٖbI.�g�9m�{��f���$g�1�!�Ҭ�0�� �R$	IK/=�yJB�;0B.0�Z.cL���yoi�4XMj[��F��F!�yc*:Xֵ6����5!UK������&9��ؚl��v�A5�6y�qe���Z{s�Ƃ��Zϡ�S��ڎ��5�pp��c��fC�=�b�+�(����b�)�c!3-"��Kdd��èz��ԘLi���"L�Yb�P5l�������tm����ɃK��I�='cޤ�j����`SgYIr\j���"%��ף֕:��5��#��us4WU��~����������=��3I}ِ��6��m	Rv�؛�Iw�>��I-٘�K�̇�$��������;��4Y6��ҋv<�I}ِ���*�$�{��������Ǳ-[�������o����ʼI%���}�InǔbH]�E,��(XG;7�@?�{� }�}��	n��Ē_I����U��6�=b�m�M�j(X�����'n��X�`y���@G<���Z��\֎&y����d����%�3I}&C�H�Ȟ$�U5H���j�V��Kvf>W9A�:�*b�I�!�bhM"��Eݶ���|�I~��7ve`}�wH����X>;�X�8`{#�7ve`�X�IbUut۱��m�����̬��+ �c� mj(%A��Iۦ�[xwfV�ɕ�}#� w�< �l�J��&��p0H�h�������s��B5�vP�[e���`�5H�lX�h�g�n��X�8`{#�7ve`v�T�Ҥ;E�j�`H�� �ٕ�w�e`؊I9e�t�N�N훒O<��nI���r"yEa*��K�e`H�TJFRmU�[��պ�7ve`�X�8`�XSPKR��
VU�I[���+ �G��+ 7v<�9���˯Yn�S��c�%s �5����9�)��`�ۦ��ɰYV5惶�E&M�;3�{�~���+ ;��ɕ��%Q+�v�n��w�w�e`wc�;�2���x��
�M'e�v�؛��ݗ�w�e`.���+ �U˫�":t���M��ɕ�|����L�����b܂4�!�&Dc��-�߳rNxOe�S�-��]6������;�2��v^�ɕ���$���yO�]��RЙ�+�EG/���ۆ'vڎ������و؝�:i��rj�V�
w���V����;�2��r, ��Rq��[��պ�:����L�����+ *�\Cc
VU�;�x{&V�c��ɕ�y|����<�q�]f[��;3���Uqw�<`��V��/ �d��	�,J�WWNݍ�	� �d����=��$���5$���srOʈ
���_���
���Z�����DW���*��T@UТ*��� �"�T" �T"�(�B(
AP� T"�0T""T"�1T ��P��B"��T"�AP��B
)BU��T �AP�, AP�T �$	B+B)B
AP�B"$
��P��UT!BT#B0T"AP��T"T �P�B	B)B$,�UB AP��P��T B ,�U
B �P��0T"��0T"�@T ,UB#B �P�0T $�EB+BB!B AP�T �BEP��P��T"B+P��P�EP�B0AP��T"�B)B!B)P��T �U,B$�T @T AP�U�@�DYP�DX�AP�#B	P��B�AP�DX@T$	P�T#P�T!P�B!P�DT$@Q �𨀪��U��T@Uz�����⨀���W�* *��QU� (
��@U�DW�W��(+$�k,�F��+0
 ?��d��0/�@ �hS[Xm��jG@:$W]wZ�̀h:::;� iZ��  2 F��h��[2  �@  )��@ P� )@ )T  � 5F@ `    d4� �A��8     ; ��� �8�v�]=���U�נ���=9t��I8]� ���G��3��7Y��    !�mu������;g6Xq죉�� tӎ�׹�0oZ�!ɫ�6���@���
@�4�PR��m�!�.Ʈg;���������ͨ�����l� �ۀvg����  ���x�.�yް�{���{��'��mE;0����/G4 =�:J4  �p��@ip ���s:)f �w: �[3��` 0 �tt��]B�� 	� M � �(S�s@ �v4��J �g@�J;���.f��;b�(��悁�Δ�se(
Dt�i�  n� t�m�  ���0�t��
����G ���q�w0:�� ܤ+��;3�� �`z�`<ޞ������z�;��x:R����'c�����ˠp  �� ���
( �f�8�r�U��wo`{������ۯ`c��X�NǑ�X{���AG��.�z�  ��`y{���6m�syv�L���O �o<j�7W�{�:^6�j�p "~�Jm�IR�	� "{J��eF� 4 �LM0�b`&����DڥH� ��U%6ҩP  Ԥ���������k�|�m�ϧ���\���_�QU�5������ DU?����
��D@Ub "*��_ֿ�h�\M�nBnH�%?��o�əpbFSZ�L��Cɠ��I���!Cw#��&��O�1)�c�LtGN�d����d$RH�1�9���h$%3̌&���-�#��60/C�H��q)�����naq �!$i$=t�#���u6]�����$���ĹvK��No%�<��v{�	s	�(F�X����5���I��0�Kr2]�&#	_O��r��BB8z�`��%�&�f���Œ>�|��h[|�(�b��<��Sc����$�4D�&��������l�)L5��/�s��<XP�/�kp���5�j#B#!d	%��b�q�̾yw�y���k�^_)�4�F���r�$�b����\�=�i�K�/2C�7 !"˳�%O�&����a��R�s���Ω��̪�D��3��١t�3Bi5�|�[{���N����ϓaM[ˣ<�Z�w�������ĺ���k�n�<+��}yN�����I.k�/ٽ�.�}�>���>;'̃
@�X�1��w�	$J:�w,�#�ֳmet�i�i2H��,�E��"����y�+����	pK(TU�2��	�h&�D]8���ٞ�L)��HSF�����'#!��e��"Fu�!I(:��	VC	��}צ@h@�Kwʻ)�e���䞫
���i���ߋ�!<w|ۿ����U;ҕ3�\(	L�mH;[ݫ9��7��1�S����g$޸Jf���D�8�]���sE�.k�K����d��a%�&��0,g��!�ɒC[mi#�f��E�yu��+����㼗-׆��מz��y����,��d/��Ns|w�f�L�H�k1�q/���/3A	ޘ]$gG���`��P/��@���}w�aH��ɳf�M$�.p�BF��� đ�F>�D�XFѓL�ֻ5��#p`F��4n]���Ǘ��zB]!5��{�����LK>A��[�a��/�C琬��`�$�h֌%��Ź���.���3=�/���vxx?m���~�4����2,>g99�"k3�Y���io�G
Ŗ���(��\+;��W�(���n\��<q"�!��$���S|%�]�1"��dK���y�;�*ۮ��Gl�N����z$��s����w�3����-����P�RfҰ��io֙o�D)�4a?�!%�A�!a�����n2�[�u�fd�+
h�JE�l�6�!��Ɣ�p�IH�27��Ć���j�t��K�c�J9�L4)�5�oD��;�	�n05ɣۧ~R�V[��c%�cX�K�k#�fr�ѼɲQ�Ĳ�p���Yk��{	�P���wF��]sņg,xg���Q��HF�$�����
T���$��-eXVR\p�abDY3۽��;ދ�Ͼ�}���qU�tR*��̶߃VB)	8@�xa�����5�#IB�2ʑ���M����k.��e��p�h�	D�Ñ��o�����X�5����<'�u7M�y��	-�pd.f�~##��K�ssh䔘B̑�
HY$5����/���XBT�VRFV渐�m��<*c0���2m#V�u�����
�$d�ˌ��5I,ֈ���E!Y���daVS�7v`��Ԕ����@��a3f�|��I	W�"]�	̃֓�<S�h���<��%[��&�!#��4:K�yl��f1�/Y�-�l̐�.Y�2P���MA�"B�@x�,Yԃ��]�
�\4�%�5��!R%�3����2�FILL+����o)�<<1"ѠEkM�)K�lZЁBF�B���a.`sWp��5iO���3������?�o<�O�?���"1VU��t�nbB	zY��_���o�����A)-/!����d&��Åc�a.�3g/�R�9Ky�×Ke�G�����&�!592��pb��$�%Č��Q{ܓ~��{���;Æs�T�ڮ�g�7r$�L��֋\cFSd���G�qB����x�H�����䇧'ń�XBy,ؔg뫨~3������t���@���$�)��)�l�@��͓F��x��g�GB�!%Ư�<��o��_�o4�_/�x��9\�^�d���c��S+�(��<��t� BH��y=��No�a_<�8�O�%�t��B|�٬�[���%�sP�"�E"9
<8�cYC<cm^ᙟe����ڗT�Vh��d5|2��!R@*��i�\�>6���o!��ė�bJ�)�`�0e�\fM�e>������2���o9\�|�z|V�ʄ�y�������m^[��������d8�������'����N
B��[XF�0,�I5��{�I��I4�H�����w9o.���$BS!Q�$+	26��y.�@��!<#�Yp9ˣ�<��B	
��o7�.y��o+���'<=5��3�l�Ѭ<���8���~�H>��	$��R�eߚ浲�|���:}�q�@���/'�s�����v�N^�Uh�Tp�����2V@+�A6o^r�63�n\��!V6H������52�Mn��ր�ff����}|�~�\�)�H�g����5�Z�f�kZa��cI� K>��yÞ����|Og
�v��&ǲaJy�=�!���(K��=��̐������y<��R6!T�\!k{7�q<�R�iB��.���-�YČH073��97�>�,1��wq�0���*sN�&��Sg*�J�(V�����TW(���<�$����� �Eς$A"ċ�V:)Qo�(t�	$�%�K�OK$)+	+,�\,%VX�Q%b�R�C�7��,f�|lf�JD�������H�	��fL��O7,%=ػ�K��y���Qg��>��	�5�l5�:'�|Ow~�\M"H1"N{��ٞd��;y�MJ8¦��M���x��l%��,!�
��x�*�P����j�M�30M�|���%�@;R���a�]Ĥ�5�\&�r3��������~�^;�����5�����Y��5IjJU��y�v�����K9���"�%�4��eIf�f��%���r�L5(K7
�0�aq!u�2����L	`cB���a3R`D�dq��#HR$�a��d��L2Q(1V8�HH�����1fBMfo\.�Čb]	��Vl�%��)%#!Ia�)���0%�۽�F�ސ�.B��!��a	BЙ�Ӑ�,�C� @�=%%RT����쀳eh��V�*���H@��L55!-	��'6�l��a�ĈE۲X�I�uS��ߚ���]v�kQ�(ծ��6���{6N�R�l�
��D�JB�y,W���}�'�H��$���7�=���{Og��ݽ4�i����m��I<&�9u�$Y������۩p��כ3Ak��g#<!	!m�IZ{�<=6��$�F%֦[0e!p%�2\�)�ɽy}��9�j<aOV!<eؤ���c˯]'��I�4y�x�ɗhqw��ݼ�����{㥟(c�M�X�YH�l�!�h�b4Bf����)�����Ѵ��_3^��7�7̗
�d�����Iy�\q�D�����fa��V1�HL�W�4󄉃b\�͘JI�ϯ#	$���BFI%�$��T#U��=Q�p����y�uZ�6�� �2�������D��I��$�&S!V�	�8K6�~�{�Mݒ���IH����w�)O7�k��sd�{c!.���P� ��p�7����p��dvB�NF��sw5�IHR&�9<#$�z�P��z�'4k|5�6���)T�aP�$ VV6І�T��P����V@��P#.oЃ WN�����F��H�B��h�B�
�X�K�<	f�_wx��H1�
��f0�c$"B"Y�	���+�7.��2��P�F�����D�{�3���.�v���ׁ9��߹���.h��\���0���aXQaYjXc.P�%HZ�Z$��)�`�<��C!K$(��F �B@�S�y��OL#C+����fNT��<�~���߿xf[$N�%��ym�����ΞO[����?r��޾C�4"�Y%�f�B[!+i�`F��.�5���\<ވI�m%��X Ȓ1�	8J��#��5=��M{��h�\5]�5H�)}'Ҥ��,,H�ˢIIB:@�D�HԎ0���	���<a ��H�"m9
ʒa�*l���c̌ F1�B2L��rOg��5�mg%�l ��p�8k5��X�����f�<�.���ͤ�2k��&���r4���	��ց�.��ݭ6�QÊ�������(Ho�@�#<ef-�p��8j0��Z��u�a͜#Y�In�p���8d��ωsP���r�V_	�a.�#��R�׌�����盖h��ͳ�
F�M�b�i��y,��xK,4���$/���#p�e.��H�`Nd�%7��G�p�3l�	���\/�O}�<���&���p�g�y4a�8K��~����w�_R�O�)�S�fs�33s�w��C�R����BRK'�La��9�ﾢ�|��1�T��C���:�4"Q��!#�U[UU׽ͮ�.����h��g�U�a�! �C�3a�o\��f�ÙB$�6̒����˭���a6O&o�n_7�����)�b�8�n�y�;�k�����L�ul�B����K�)�ʐ���EI@i�9C��)�J柽��`N]{����`;,�F����au�<�rf�����>�-�kP�F�Cp� (Ġ�)';�Ϊ����������U*�U�W�������UUUUUUX��

���UUUUU@UUUUUUuUUUUUUU*�UU�UUUUUUUUWUJ�R�p�UUUUUUAĶ�UU_|UUb��������UUUUUUUZ��j��J��U �Z���;]*�5T�*�7]h]�2�0��f���&j�Y	P�ʪ��V�U�R[n��j�����֩������tUUUUUUUU]Sŧ�#�aZ]��;��UU����8˭����G��P]kmu+��h��
����ls�mI��x�����iP�`�)�WKn�����-�J@5ʶ[��(1[ �UV�R��6��
�:���U]t�Rԩ���*��g�]�c�+��
�:4	E�ʪz�z���yĶ�ǩ��UU"�e]*�mT�͠�6ݘs�c�nU�RZ��,��@�UR���.�*�+�vP:��?��_,�U����)68{2�t��m]UU*ԫUT�:!V�U[UT�R��!��j��Z��j���rҼ¢pB5��[G*�$���k�ٞ$�G5ù�X�D��'jL��:
�c6+j�UgV�8�ĵ�n5�W��>y뮌ŷ ���X5�["���ZJ[ U -��� d(±�ܬ��1��Z���^��~�����-�]e�Wv{d�<�U=����F���>��̪��U��!��u��Uh�:�����8)��#�8���UuJ��Ԫ�U�����>�(�;!��UU@z�8��CaYWh��fUΒ�	zհ�V�UUR��/)-�d�
�
U�U��*E
�UU7��U>�Z�<�X����啸8�r���砅�K��M�ֹ��QdV���B��uUUQ�����@���*7��m�T�Y��R����N�\I��ķӻZ�H
��23��a�͸!�MɆ�5N��%�{^�+�;;mF�O�R���ۛ;�[�+'	��y۲v�T�Yf ����ݭG]f�v
��e;������nD���{N!�ʶ�J�M���y�)`��s�N��1[]dU�D��:�*z��<�dz)cЕ��RhG@Y��<s���]F[�^l$q���0\��1�lZ����Bm�ٕ
�W$&`@J�ĕ�� ������~�A:ٮ���t���*��kFBih@�9Z1�Ӄ^�)z������f�J�UpUqS�@�bd��᪍7E\ݺ���9F�A��-mVȵٮ����q N�$�X��U��B��,k0e����fR}�xj�B�O,k�!��ҼYw�2C�غ�Ĵc]��^vL�2�X­{V���Mu�v������9mQ���)�n��^��퀹mȵF6�ux�^�n��hc$����IJ����,UVm3�m��qPj7l�mՇ�����ͭ���v��uX𤊜q�Ɠ)����sZ=U�W��cE�ۑpv����v�e��
�+5�`� �Ll����X�p�*���[�
�m�����gm�g4�v̼�P̚86��JC��d�ux�'�Ѯ���[�!L�Ucz��m�U
ݶ-�!-��Y[+l�]Q�U�1�F��Z��&�4�1G��R�m�q��ہ붮r--$`��L��r�P�;nwA��uN��Ӹ�.N�N���3�+����9�2 cl4��/Z뭟UN����y�;h(N�J[3�<���=��W�r�J��UT+�s�S��j@ Qj\DT�82:��nܱ�=5R���w*�(rlѵ�Q�I4vl�,(���/*��1qez��;����UN�\��`YAhH���j��:ͩ�������32�t&°Q�9j�^�ڡ�U����kiV�(��7UTںT�n�n
�e0g��ȳ�Ul���O=h2���ڝ��Uj�m�VRZ��<C��P]�F���<���i�V��R]Oc��/2Ԣ�N��n	�VVVTۢn١�ϣ;#l��R�[nf�`\�X답��-S�*�J۪Z�vc�i��@5K�eV�CM���˚�]l��cT��:�%�`���-�5lՀK79 
M�)���9_/'l�2�ꆼ�PF�7m��sJ������[0���.�Z��n�GQ���-R���B�����P�����c�Iy.4�r��
e�ۜQ���^|z��<�\�9��Y�{&�s�	�Z�v*��������m]j�(4�;`�ʝ �s�j�����4ک^]�V�(s=j[a�Ƴ*���n8�smPU_}u=�J�WUJ���u�C +�6�UU@uUP9�iV�a6���dઞ8�<�X��}\�2��!$�z��I�(�:�����UUWR�+�gM�H*��)EX�k5�֠�Cvw]
�v7��;v|y�
�]&znnv��5�H�pFe[k��a�h�e4�l<�\�z��Xv���Vm�l��+6\�z�.�UU����iŸ!�;UU�X*�W�h���Z�Le��2�T]ٌ��&�\�m�*Q�WB�}��o��ÇnU^\�����!�۶v�j���륜ʻ@Oh�8�9����iYUZ���+vʵWe�ΐۇF��U�UuLb��R=m[U>��F�K�}��[k�� %��SU�I9���j�
�B��5U��Z�U��
ZC�8҄�mw<�uUF��Z�8Y��P檪�j�.Z
��.�V����Hot���ƺmRn5�U@���
���UZ�Z��eUT�*��W:((@�70�kMV�-�
3sU@UUUUTF�V����ҷmZ���|Q��UR�UQ�Uj4UU���Ǭ�X�7d��qz��^ej���-*�@PT�xD�U�Gl�\�nYۚ����Uj����� �UU�j檪����H����g�Z�U�v��Y���7T�tq�T� �u�-F1�4	��x*u�)<�p�5U�]��ゕm�j����08G��[�h
���������e��������V���*�U@UUU���������V�z��V�A(��%TTU*�]��nүV�W�QEUPUR������ʪ�ATT62�
��5UUZ�X�5v�]������R��J��V�;PQ3�h���*�V�t�UR��[U�eZU�����V�R꺹P*��UJ�V͠ %PeCd&��X&��ѪM��V��畀�2��]�`��m�檪�]�Z�HZ���������U���V����(��^�kX�ɹ\q#m���@ʵUTx+�mT5@UUU\�UcM��A�6*�YZ�������.��U]@n�a	j��2\R�d�sUWF�]�lP�M�ꇰ�nU�D��UUUUUUA Ub��(�J�f�4e �P-@Uj���Z�P(
�ୀ����`*���O9ei�٪�VV����	���Tgnӝ5�iv����E�n��Nt��IU��W#,����v�V�mUT����UUUQ�*�WJaf����keZ�<��ŵx��J�������(��j���YZ��5յ��8q/-UUUU�[tUUUUUUmT�]]I��J���X+v�g�����P�-l��ãT�4�θ'��vW��8�\����nSf��Mv���N�,�UV�T�mT�Զ���à���<l6�UUmU�*�	'gm<\���ym*��ꪪ�'����n2�F�|����X�^;Y4l�)Ӵ���cN��M8]�r�mKr�K@U.�W�"�n�@q��kcr2��y[�j�-�[`;5�u��	8�;�R��W��x6;'g�8��s�����y��÷lY��.��C�;B<�mQq�j��X���s+�(��([4�e��5�H�uLE�vCUn�ɛ�Y�Uhr�ٺ��Tq�ݒ���j�n��3H�!7N깮%�7'm��Vbl��L����a{a�;Џf�Ṵ4�ؐ�]44���4s+(��k�ʶ$¦ȯg!r��j���]�M����8Ҝ�/C�q��N�������Xv7��b�yyYӎK���)*lV��e^���T�*kr���5��5u�sWlԨ�rV��(��-F���#UUv�x+Ud4�-X)�iIlk���[e�4�UUT2B&C]Q�NU;u56ڪ�UV���񢫪�J��_�����UU++�\���	t��UUJK U���UGjm��`��MUU*5��e�'�~�
�s��������J�PW�s�ʀJ�@v��8�	
�h��L�YU+�U�jv^[����d%U�gp;654:	T�
�]8�@��e/Pۋ��΄�۶ ���]���*�������n��++T7���7�!�Ҫ� �UUUUUUU[U�T�-u���+�t�UB��G��j���j���Ի+��k\�+�@�.�U�T	V�)v�j�&ݥZ��n��Z����%��V��B	�6+k6�6�U������������ �ꪸ��uT�A+�� ��"�UY�خҵ�UJ�Umr�I�����
�������nh���)Z��nf�UmQ�UUUK���������������V�\�UM�uUTڪ���jڪ
Z�qUUJ�PUU�uPUUUUPU�UUUҭC���mUUU@UUF��UUU@V*��������UU@b�ڶ������]@�UT�UUR�UU*����ʫ|���A�h�SU�͗���B�gH�UM�����j���lR�ԫUg��`f1PUUT����0�Z��]�eZ������3ڞ���M�UP{s�x���Wʪ�U[).ՔUj"Ux2m[tA�u͎MBk��(������8�������w���'E��`$N"	A`U�� 9�!�1" D��H@��БXho`zJ0I`�
����V�`چ��s����8(R��W��D؛Ux�O D��PM��&���6�z(x C�n�� z"*��=� $H�H�x���D�#"�U@6"|�� ����b|)�Y�� $RD�_�6q��+ _QW��'�Y@�2!A��E~^�j`�)���^ �'�/�� ���t��)�$� "�EQd(��(@<Db!�J����(sUF��)�\6 |�:P��� @< �����T E�{��Jb#��5}j���)�*�vV0H�d�I�Et�b��8�����1j�Bz��:�W�
�� �D�nQt�/ĄO���A����xlD������!!(	��a@@��/��V�* QB @`5(�EB `�b)1�>P�T1x�T4��2I* h�����4�������H����	`��0��	
+F���"�)�m�e�BE�HIYE����!,Im���J��R*A�#(҄ @ XHIIe���"`I&�=�4��:!"H��U�Dx�=`�B��U1j*lg�h�J�0"�<�G��|�z*���� *���е��b�b~�P�B�"ȣ�� ;G� �$��XNrr<�HNKd>���UX�D`*��F*�J��J��5���UUT�P������ҮH�쳅{a�9��4���3�06�Rd�p��/���P�S�Cv�넍��Zb ���X��3�xz���3������_%�d	����s�C�5� �������j�ϭS�<k\���q��:mqEV�p����r�[M��:knL�mz��X�<g�r�'��{j��8�0�ݻh.y8��.`x2��zݎ�㣳��Y�:�Sa�M7C ��7%�jٵJ�
�) �,�C@�*�0�e��1͊��6�"!�Q���g�`�s�܆��$�ܽm�ep� H��E�u���6ڥ��iy'q�.d��Ȑl�t�[��nUgT�}WcC�Td�GQ��݂z�ѧf�2ts�d�6��(f�
7CֺxLF^���v=c;8�7KpM���Q���@S�� �;G��OjꝔ�Ņ����+ֺ(F��$��j�n��cUg\ M�[�.�g�Ż�#4��qL�l�mk7����e1����x��k�R�<6�':E4G[��!AVbumf��;�� ��]����E�a6�ٕ�LM��
��6N����v%"S�@<��%��m� 9��h^jtUUJ�d�v��n̡PUB�����]���J������%�y
�`��5�nڭ��2�49UIF1�k��.x�:���W]��.
�L�ul�6��g8�{v��i��v �T)p�L�mYF�b��J��&&�O�5&H
McPq�]��O=	�y氪����q���h mc����n���G�xL����s�+�n�vǍ�3�q��p"=[]� ���D�1�1���#4a6�H�A���*�	�vuAP$��s��\�	����v_E��SܰC�V�PM˝N�1�\$��m�J�M�ӝsdj]�Aɓ-U]FFy
a�����3qZ��`�W�'64g����c�m�ص�-T[�:�����intth62��re�k��:�3O���A���N	�҃�zt6���A|}x�C�>U�|��{����>�i$�0��X�KG��6dt��R�ݱ��O]٭��*v:#��a.b$,��/��ؙ��9\�k^����5,r��i��oWG]���@��4h�\�S�fX"��sǍ[�d��7X�"sn�*Ě)+iW���m�VcTl���Y���n��ȋl�VM�&��Imv�ʸ��ɺ%a�t"G�r��5��#&ToK�᜻pqu��U�T�u�����.�nd�Y0�@��r���(�x���90"�N�1Ǟ����6�ۛ/�H���I%�w_�󽴒�y��@��^��oX&/�3������M���}� �u�x w~���@?v\�3u��E�#� w��}� �GĽ�W*��{=|�D�y<I%���wfl\`��ӯS������~����m߻��߉z)�c�S������O��� ��^r�}>־�v�z�.x��ܝ�5r����xz�c!�ZE��2���F�8w	j��-�h�͔֙߿ S����I%;���ImF�X�J_v_�$��ZG�tA�Į\�� ������7'!YOPb�D�3��z�m�I.��_�$��Kx�K��,WMՔ�}����x ���O��� ~����w��B_.���h�I$���H��OI.�c�䗫�ʽ����� ����ܡv�6������$�]����%��q,I$���W�'O���z���69xĭ��њ��[K�c�0���A��
ӮC�݉�ۗ�=^|�#�n� >��Ͼ�~�/C� ��z���}�x {��������P����%���X�Ko�/�H�<I$������96�w����˨M68eǁm�=�s�����kv��!� p	7''9ﾏ�u�����< >�>���^Q���@/��� ���}���=ǀ�~���>�fML��l�� >��_} �7�q� {��|� ���� =�_��tC���]k t��[\3]M3)N� V۬OE�7Y=��s�d���G/��~��n� =��|�	.��x���|�[�K�Ee����6��� =��}����rm����� -���Kv��bI.����;))��@/�ޏ���u���Nsm��� ������� �E��1�q�� >�����z ��_}�)�g���s���[��ϵ~.}�5Lj�}���< {޾�n�| =�}���NN��.��8u���WGg�q��la>y�l��MݮƷ-ݧ�mρjy�\�m1Lk2�� ����>�{r'�$�����w�����X�K�B����%^\�_} ��z> �����|� �}��Y&��O�|kt�ɜZ햾 ��w{��{��������} �u���߾���03w���$�}��� ���}����˻/ �a.�)e4�
��ۼ ��������>��/ �㣜��O��s����^낵�,�Mquu-a^+�!��U�f��R����i�[�6}j���q�c#ً��<qs�ty�£�{:�N6b��9��@�;u-s=q�!�����R��Sc�C�mf��9�hDK��<q�F��v��m&#������h)h@庮���S�`m\I���u��Μ���o7[�j�S��A��'�n�W8���\��rAa
1[��I�6��<�Z2�+9����[��q��
Þ3��t3���s��˹225];)
Э��k�|�e�R엀nǀ}(�'7WI'M*��f�ݗ��]��������;�p��Ge�IJ/.���V� ��d� �v<���/ &�[`�V�����r��IvO<v?�v^�)���P��銛�m+o ���ݗ�}Jl� �v<ܪ��o�%��gP�ָ�]�6Sf��m��B �{oEŧϬ��v��u���&ҵ�n�=xԦ���c�9\���`��TC,@р��o����}'�?�'ec!����2e���1-HP�P��!C �T���ُ �_��/<���րAK)��U�+n��y��p�>[���M��HVҩb.Ō��[x�+��6g��O^�)������	�M�h�M*��f�ݗ�|����.���c�oj�e��;`&6Wg.S��<䩠]��鎫��oe���N���e�V�[V���U�w�|���۱��p�>[��lV(����j��x��x�\0���M� ;%�m6�Uo����{��v^�_Wy�W+�YX�2< ��UԤ�*-ۻM!��f�ݗ�|���۱��p�;�َ��˻i!]:I��>D������`-�x�t���r���M���=G:�'G��K�({g��pm��G��[I�6��e37�nǀou� �n��>D��	
�T�
�2�!Z��ou� �n��>D������\����$�����U��`Rz��6< �v<{�݌��R���Z�V�[��M�N{��ܓ�=��rl�UM�'��F��o� ;؋P���J�6� }6<��Tٞ>m�,�M� ���������Y-�v�y���7��mɞy����cr��v��t� �� ��l~0��Xț }6<�����MݦƐ�� ��ŀ|����c�7��w�tզl�+�	��|����c�7��oob�;6Z
R�4��[o >���{{�;#�6��X+�2�8�
��;�p�7��`#�< �l{�|��bD�	1E�AI	"A�	�Vg٩�a)hW���b���kW!�K\��gA����p�n����;w�A��'��r��Ę����ݳjw�f�eʶ�dv�h�f�؉���t�=,�\���e�D�9�;qw%�r��f�.��v�N�f��)KR]R����T��F��V��/�>��>��0�Ӈ@]��nܖ&U$�m�v�:�y�t�߾�9f�I��0k�B�&�+q#���Og�zf��l��=��3���v��xGAn��d�1`�&6o����[}�����`v2��U�ݢ���]��|������`�ذlE��T[Wv�� >���{{��e�uV�FڻH�V$Ҷ���`�ذ�ԗ��Sc�>U�8���e�;�l�7��`m�/ >�ٮ�H��b�{C�L[k�!�^3�E��m�Ɍv뇏(XϐxF�	s6�����]�|��R^ }6<�\?s��W�&���7�����n������nN���߻���J$��� �HЇ��m��W�U_a��� �Ix�jK�;
��X]�,��+B���p�5M��}��� ٱ�PD9t�_umU��`���>�R^ղ^ٮ�eQd�l�v��Sm��%���.^ٮv�,˲y���N��6�#C6SX�^�Ŧ�P�%��
z�F��''^��5��ͺjhZ�����w���ջ/ �mIxުں��v��4+wn��p�r�5I��;-{ׁ�p������I [������#U@*O �'� 쵲��������Q�.Q�\�i����<M:CI l*��HJ�P10a1H­�%m(F�*ń��ٳp �6��\Hzz�(l/���>�:��С*J1#!$�#�"�̮��$V��5]&��K)V�ws�ha����l��#ȴ��f�!`����]7�.��*I9�f��d-�5����Ҹ�1��t��z�ݓRJEy�߹5�����09KXAӎ�H2A��V4 %`RځM.yp!���.�b$X��>��B��z�.l<MI�5=���x�츹Y���$53\	��<<��_E8�2���HG_#��8m4,f���`]y�MD���\p���zn��&e!H�%�2�� �%%�StJ� HLhT�u
M����f�ϗ���((�%`:e%HBЩ�
}�!9f���)t��8z|���H��(�B�Rf\#	X�5��!BV,`FH�! >A�B1���%��`FY�b$$�|U9�Mkԛׄ��J�	��=���2��`V��9���!IFV�>��:,'�RС+����]0��9�nXT$!6F=5J�-� b!�$`DcH$��"CA0��T� T�H�>�q4d�H��`}��޾��	,XƋ��>�ނ>�O��č�!��sV�C�E�h�@�7�Z��3G����������!��_�~������L�EGՊÆ���Qr(�b�$"�H�1�� �H��z����`�b;P�>O�~ �x	�W/�T�Ü�����&����-:.�Э����>�R^��/ ��qm���7��\�4"��+w�$x��g������m�/ �Ԕ����ϡ��csσ&�p�IEWWe���㍜�렍-��U��dqyu5��j\� �G� 6lx�jK�ʮW����� ���_�,ԕ��]����_=�Ӳ׽x�O<�L����UvO�U?U�E��wj�m�ֿ~� �c��K}�e`�<�v"�A�c��EГw��R^���7��V I��]mUW*�8s�QB�Q	�@��64 � �;�o�3rI﴿��8�+n_ ����'�|��O�I�����=���׀�l�u�uk���,ZS�n���������
�H]P�f���9m)�n-g�6���u��ҍ6g��z��R^ I��I���K����lJ�v��e�/ $��	$��	6<�\H��pTe4"��+w�}T���������${���'�{׀}�DEj�Y�.�V��{��Հ������R^���/#�_�N���;J�u�lx�������������|�߾����>���C���z�	nPn����]v�Y�/�J�F�܅ݫ��\!�9}t {gh:���H�34�9���6�:Ϯ=�\'76�z*�T�	�9�������>_\�ԷH�M70�;qv����N�Cu���(������5O RIѶù�;; A@F�f[
�!�����I������ilf��yyy4:���Eo&�ѝ���.�e���7Yp]�{��~x��/.=v�[׊U9��,$�3��0�l�3�]���fj@�6��)!�<͂���V6ށ?Z����7fW���zy����^�I+��w�6<�Uq#�{+ '����%窹ă��J�t�I�hM+o �����5����{�/�ٹ$����䓓�O�掹�(ݳ<zt�~������ߵ��x=<�?W+��{��7j�u�4�wm��v���%�������ߟ@��~��	6< ��T���BI�
LV+��M�sLϕ�{�ЖnyBd��S:�6�O{��AYe4"��+w��<�	�e`���U\��k���'����j�vb*�2ۚ��{��7��@�1�+��z�9'y�krO�������[�(�����u߉X�n�< �����>}�%���G��<�����*�IF�Wi+i����W�^���<�	�e`{�U\Kޞx=گP�Z|]�� �c�=ʮsޞ�� ��������t���,�k}�ĺ䖡kc�85��w5T�=p;v��ZQ�f+����:~�&r���v�7L�ZV�@�=�+ $������Ur�@M�x��W��T��݈i]���Ǟ�U$w֧� =��N���UU$v���7m	�i"�ڶ������'��~��Gr '����X H��
H�81
Dl�|޻���'���nI�b\�4"��+w���%�O<��e`����o���aG��t�����]]�X�2�r��ޞ=jz�	�2�ܮzz���1���5b��f���(�K����Y�6%��k��6g�:Iy�YxRaV��4�������"�K�&ɕ�W*�A��e`EQ�����e×�>��o����~��l{���O ��߲��G��UUq �Ee_�5V����� ����$�+W9T�����~^� ��mEv�[�Z��UU�{��O{��rO�ϯٹ9��9VP�Q$T��<��Ě��\�Ai�PTdFT(���W���=ʮn<ݬ ���e*N��e�]۬ ���z�ǯ�$���	$��?wu�?�ݽ�z8�A���q!]D��s65x,Db�ѹ㍴�1�K<��+Z7.Ht�m���{����2�	6e{��y�	�*�hEE�� �ɕ����ʻ?~�� ����v�^�/��+J���Yt���=��V vlx~�UW����׀z~���M��V­�t��������x��׀Nɕ�������������� {/���.	�U�����U��������Xٱ�W9>���[>�,�SbgmL),ZWh���ֵl�(�Ů�z���y�;�#P�%�ۚE�aM9ڱ��cqn��}���_ne퓧lv37��ŐG�����螻3W/M�Kk�ݲ���s��p�ruK�8�X�܉����vx�rcמ�ۓQ8M�����D.'n%�As��k�04�k�Q�N܌��;�{+Cl�����&&�n�Ƭ���}$̕<ǤfA�dh���o�x�>zk�k�y�O���^�I�ûpۃp�<����;���k)*,��~�����Mٕ���\�����xV�x�v[T'L�	7XݙY�+����v��<����2��;������&��.0�s< ���\ ݄xz��U%'���O{�Xշ%5��Z1j���wwX~��$����~���lٕ��W*�UIo��l'e���n���K��rO}�훒tT_z{��}�<.�^+�[.�ڡ�&��F�h�����WX�Ŭ�l��Zc	������N�)7�'cP�>��X�#�"�%���U|�O{+ ��&B/i]n�< �}���I�8�$>�c	�hċ�Z��`X����ж��	)���/|�f���ٹ'�}���V�<�Q(�]
®�m�[^�&V�9I{}� �{� ;"��7j��Z��Lw��R{�V�����ʥ����S֛���N�I��&���=�qo���^�� �&V��Zߨ"��/-�#F(F]�d6�-��X�|ti��༚�fc���5��m�M�����_ O{� ��_���	�{+�9��~�����o}�k��ֱn��M%��r�UU]����X�{�V l����RF�<+T���S��v;�'���I����r
~�A��"0HA���j#�#bิ��F5�D�d ��R�b�6�~z����ܓ���srO>���ؕݬ�*�E���ʪ^��Հ�� �mK��UU)�� ��g�[��@������ꪪ��^������$ٕ�oj�e��;e
�BV�$��x��̇,��]/j�r��,�����	n��=��yw(t�R.���]���^���$ٕ�I�+��UW�zy�������e��d�a�ܓ��f� ?�2~��훒O߽��wIy�Ur���[/�N�&�uc�	u�rN���ܒ{��ks򠟕@��~�~���y< �}��sk��q2]���W9\�Jzy�[^�\0�T����<��#	!J�p��`y������S20�����=��?xnI�gߍf���0ю�/�}����?wN��wN���?��~����d��iYc�'���,u�v���`�I��Ή�n�(�;���Iю/�]�̥�|���� �&V wv?s���|���=x��#��i]�2�X]� �&V}ꪮs���=��~_�� �c�~���q ��u�V�(���u�'���=\�9�%��� ���QʊTB�]�*�o�+��U\�*���������I&O�N��I�I��}����n?AkWR�2e��nIϾ��rO�E?~����!'�<-��R�-��T:UUϊ��RQ�����������eMCg�"��~3��;���Y�5�֙�Hx�nr����fO�.IGD�i��YCd=�O ��20���#����|dX�P�o&���5�#<��_7la]��Aɤ��ɰ��P(�7�4��|P-j	��C�&�vEf���!PjbSݪ}�S��;Ͽs�y���UUV;�Ur���v�5�U]J��WB�5Ɲ��=�}}/�#���b-�.�]l������GWk��aD�Xr�g[N��ݪ��ff%�4����v������*�syKm�=����l�8���E�"�am�����$d�^V�q�.6��bC*�Y�p�pv+�*�M<��r�5I��z����s�t[�n$W��ۮvJ,힞 ^IՉ�ڜ�3�;��V��"��N�n^d˻<p�f7p�_��oy����%0�B��@k$ƽl�<M����h��;n{t�q�5�j��(��b�&��r��!8�����a�z���u��H:�)b��tc,��fR���Yz���+���xm�'��L d����	���l�7N���ɴ[���%a�5́��K�7�/�6�x݉V`uZet�R54��hF�]km��pFr�B�|�g��p[�5�%�Հ�2<zvy���p�
P���/������C�&e��a���\C��h��j��ۘQ]�\��s�xu�^y��-��[���[�̈́4��^P���"�8���C�&L�M����G�iӹ��H͗n��M���<:�u�>�O��]S�x�m�R��RD�mni�Tjj����&�l��n�
�W�U�s�� ��B �:Nϳg��e�2"�W,[g�ڭI��DZ��FSb2�](`��{q��f�݃[z]��dzc.ʰp�vՓ�&�X��F@]u���u�]�.`A���tqᐄ����]��������1ׅ�Y�AR��+5�
�{bݸ�(�xϭ{@��J����PjM5�aј�Wtl�+�v55-�k�ٻl���e;uo@�-p�#O%���mǠ�\/8��3p�v��y���=�r��m��� LAe�KK%0�#�ĭ�+�ճ��MH��Zj��g��3����Z��5U�z��*����UV+]�n�
�2���6rf�X6��B���-����T�@K�-��jb^��R�`B�-�֖bV3��@�W�6��DҀ��0h�����u>p�
��hD����pW��W��g�� ��w)�S[k2�iXM`�k�9�\�<���֙�45=T���۰s���9����²��]����"����b���c�q�Ō8�[�[�r(f�g�k��\�j�1�����6���$61�����i���uX�\��W��Q�
qYն6I0��9�۲�0Yf�\��ND��\��	�y��{v"t�&�B�)�j�1�F|�ߤ������u{^I��)ǜ۴����g�@��d���������痜��L��;�t�O<��R��.g���� �v<.�_��\��w|�`O{���v1]���wn�������)�?_�Oٹ'�~��'�{���m?ކ��V��0ю�/�{�=���a��UW9W�~��������QR����!�v;��W9�]���=��$x�9\�����W�x�c�v�L�E�0	$��=\�r�OO?��=x�p�>��-�]�V:�Z���x��q��7L�ڇ)s�MR��聓D�݅҇�I
���V�(V�Nۯ�'��a/	=��}?��$���훒}bN���0����k[�}}�}��H(0"�FH	#*A"���"��TP�$D����\A��s�;�&�����c�U$Oy? m��VZc�o��M�X{����x�����e�n��`���
ف������ �O<.�^�s�_����߭۷v��t��wn�����|z�w��&̬9ϯ���Hi�X��i�\��Ԧ�P6BVgn�X\�%�S���/�ln�݂�˻m�����;��I�+�>@n�� �����S��E�� �c�~�G�������"����DҽK�^[i�e0�ճ �������np�l�N�k}���nI��ק���O�f�.Vx��I�}��������v8`}^�W*�=�05�Q<J����v��tL	ʮWݙ��=���ǀ64�:e��2�x ֆ+e�0�)�]� �'j��&���p�;��s,���J�Lw��?�2����U_ ���^~��.��Ӷ��m6V������ăvy�^���?�_���i��/��9͍Yr3��� �B^�]�~0O{+ ���UU���\��I?M������{���7$�߾ٹ=�B, =H*UO�
q�矼�ܓÿ����u]�IQt]���p�?s��U~�~��v��{��"�K�>�Ԕ����)�h�J<��ێ^(�����=�.���DZ�!*�g�@���7�k��`�>��}�x���HK�|�����/�+��n�m��ݏ=�$yz���;�?�eg���%�t��]�m�^�z���a��^����g�٪bChlV�e�n�=UK��� ��� ��x����^�u=i6�:n�ӧHM��e`��s���~}��_�^�~��r@�0���F���g�O�U�M)��[FZ*f�.�.Nr�
���#�v[��&�V
Z� ���xH��i�̻gny�qu�aX�����'�ՂAcvM����t���=��B9e�[�(�+�8��\s³�ї�՞Ӽ�@���lC��^aqo`]����^��a�f���G[� �؎3��6�r�ݶ���G���1�H�V�&���&���.��5l�.\ӭeת��7͒����[��66�50^- �K��`�M�����XF��.�묦������8F�6lϠ����Ixݎ�r��{���;�z�c�7E�lWv��/ ��� �L� �v<�W)#�<#ºĮ��J������~0	$��ܪ�$M�x��޼t�Jyv66S�`{��8��� &�<)[/ܪ��]����+�J�[�]�X���I� $P����~;�<�{���7$������;طcl]�sD`cƕ��:q��N��2�/:�f�[�s`{:t��:�U�|�n��/W�x�\0�e{��UW+�����Kä邫��Z��9���o@6*�0��/�D��������rI�w[�{~>�7�;�N�:v�������n�1��j��߿e`�c���W*�IOY�^�����o�1iU5ٞ���ӻ����� ��?~������9�U�{>����llV���wv���/ ��� ٳ+ ;ݏ %wU�.��S ڶ�X^\���-Us5b94�'f��3s�q/5֞���ɼ(�O-�l4����|�`l���c�s�U�z���$'��M�D0l�����'��w~��Wa��� ���~���r��x���Ұ�E�u�g����db�b"�#"���`h�*F"�IH$	x����uG��{�M�;��ٹ'�$�6QVWe]�m�{��qo����G� ݓ+���%6y�t��;O��Ҵ��w�}5� u��=�W+���t�y�l��ܪ^�Q�Uv����o�QeW  (�U���`(C��:;&��%�n֞YY��6�����>��������Id���ʯ�v{�X���+t�J۴�P�� wv<�s�I�'� ����	ݙY����~��]�������6]�o �,���6l���\�^��V OO<��$�J��E���+�S�<`����6<�r꾪�+��{���a^���e�0�ճ �L� ��x�Ix�8`�����vS�:��=hݴp��d:���!L�˹��\u��L@�h~���<�h͂�Y����`Y%�H���U|������Q(���.�ʶ[f%�^{��$w��V�{�X�g��UW��U]���ԩ4�� ���7���X�2��Ur��?����*쫔���I�:t��X��8�=� �?�$��&V |n��n�I[����u�n��r�^�'��;�{+ �fV ꫁P�t;ږ�kʲ��e)��A��!@�EMf�ĨB��#�NZr�v�ϗ�ɧ�޺�a�o�wT��$���d�
�-���\�0�Zp��2�ݨ<�d����k=�m��k�m��;UЪo�R
 <@{m+=����Bn�ݷ9 �m=����["8���%���0,�0���5Ǻ����<(x�����׶6[VǶ1�������+��oK���<��C[q��˙�5.��.��"D\&�y��q���u��"�7 �L\�@�퟽x͙X�2�U�W�'��l�ĝ�IQujӼf̬�s�H����'��Iz���$l+Խk���gj�n�I�f�a���K޸�x��V M�������Z�E�u��s�zg�޸�x͙X�����������r��{�����ـIz���UOO}_�{�X�p�?W+Ҩ��>T���Ù1߻�k�Ec��Mr��$�dk�)u��)	�B��l��-����LP�w�{���I��l�ꪪ���z��=�cv�i�n�	$��ͪ�����6��!�Yc"A�HBKH�"F	1�X�<b5�J�*�, �&ȵ� I�!�($��	�f0�0 C	LQ�L �����,#$@�!�HH�0�X!	1�?+���N~�7$����6�L��9Uă��V�n��[��]+�X�{+ �qK��r�_�Uʫ�O߲�߿~��>�����B��I��&�R��X�e`{��*��{��;��WX�mAujӼ{0r��s������Oe`n)x��l��v��*�� s"P��E�S7kb�-!pmU��E�1���t�R4v�6<NMqV|�}�ɀvl��&�R�\�9_ ��e`�U�xuwi!]ۤ�u�vl��&�R���nI�����T�"��~'�J�e۬������2�u���i��!�o �0I �)`2�M:�o3'�ة�*xZȇ�1"\�$do+�lME�! �xhA�%!��0�B�@����f�C`�H02)
Ѳ@�� &�=!Y9�Yh�G�Ԑ"2p�kll��8ĥJ����f���A�%�|!��\�����:�E�xy��\M���	<�|癸�=p�ą���}�<n�����,d��6y� ltC����'3�����! �"��|`<dM���<���\2�T�|��RRXLT��R�6F0.�r$H���p���Ӷ,ap�Z�` �	�1��!�hC�h�����}2��	"E�9ͧ+�<�XF$�X�9��='��<�s.!.�~av�.�IP�RHB�b������ ��
�'�'�P<OG��}������EÈ����A<��{��";�:���w�7$�g���lI*o�j�����UT���V�Oe`�X��/ �V�wn��j���+u�I�+ �+������������������"X�������<��[��/8
�:�K�/=v�g��Wv=d\�?wI�<�_+�[vF�Ks?����~���|���x{&W��~��������o���ۻhWN�ݺ�'l����XݙX�̬�W7k¯%u�+hB�E��;�{+ ��+s�JI��g�xzV�+,���q��&��UK�{��6Oe`v���UTr���\���� c�#�(�l哓~����m�|[ٺ�!�`�XwfV��W���e`d��'�C��>��a��l��3js����]���Rb]���+�k�ƮɩL$m?N��y�ׅ��Hwn�������L�l�^�>A�{+ &��$�)X�X�Lw�l��e`u� �a/=Ď˩��ۻW@��Vـ{��V7fV�����^���uWv�A�&ZcN���`{���=�`Sǯ �ٕ�I0�E�wm��bI��"�K�?U~�*~���@����`�2��W/�9F�ϧ�v�v��(��u�BՄ�cM����~��6����͕�l�d��]+�M����u��Ռs���-��A���.��r,,�GX�C�YW>[L]�h�c�^���5����m�3�=N�<r9�-$f0 D��������!oq�,�P���i^<��.!q��s�6��M�����q[P���0o�A�����"����+:��R�䓧�N{�ϟ2\c�B�N�E���[��Ͷn���۝���e,!��p�.O�b�-���(hl7�?{�X�� �k��^![JYuw��U�I��$��H��yO�{�+3�꫰ڈ=W��HWv�7l�7c�E����s��Uw���X�ߟ� �UFʵ˥vU�[0���̬H��R�x�	�xm����-1��ٕ�z���x��?[	xt����v˦:�I����[�矶Ӥڻp�+k��/T��/�w.Nom�3��ɍ0�������xϿ�� �a/�9ϐM���5Vʻ=m��L�х�jnIϽ��xT<�
�H��
" E����kܮWǗ|}x��e`G��{.ҵi�v&�m�[	x�fVz��B���`�~0�PU��+hBE�����r�r{�`{�~0��a9\�U){R^!R��,���c*դ�`c���-�/ ����>ӡ���cJp�q V2P��C>�U[�F����s�j	�t������9YYY�`)wn�vπ��E�%�ݙ^�s�_ ���DU�=k�Wv�Э�[R^�ٕ�M��\3ܮRA6/ ����Aj�T��g��	���r
��� ��7��]���<z��Icv+m��t�+u�I0��`l%�z��� �[ү62�&5wJ�0��`�\���	��X�� �l��IN�&Zjղ2�X;��j[-� ИԄqW�C�K� ��{c]/bwn�M�blـE���ove`Gs���`�$y+��>$�E�� �ٕ�I0	�p�"�K�6��e�J�Lj�n�	#�����<��^;�+ ;F�*�N�$+�t��`��E���N����U_*����a�j*���Ք+��I[0���wfV�0wc��IdLg�v� �R��#4�J�"	ye�J4�#QBh�\h�ፘź�5Gx�̬v8`���W9\��j�=x�{�[����e:T+u�n��W) ��<T���'veg�#V�ו�e��cWj�f w�� ��K�7�2���}�#���-�v&�I���U]~s=��x�߲������吏�^J���%ujӼ{�+ �9\�$�x��<���/ �����+�*���(%�T<�E$A���^s��^����H͆�f6;(L��e\��7E�U�#ێpY{]n\E���{c����ɹ�aS3�Ѻ6����ˬ�H�V�C
YtLs�����yu\��R5M�اU�.�8�x���\�u���dL��+�/GQм���[]�+Y6�,�u�cP��|-�ͺy�����\��ryj�Y��)t�43I����s���Q�k99;rs�9$�Ӈ����A��Acfܺ�2aM��E��2���͸��s[:�tn�KA�7<t��[�S������;��ۊ^;�+ ;(���-]ۦݳ 'v<�qK�'ve`��?�"*�=R�����]�m�/�׀N���7c��Us�{g� w�=Mr�lVӼwfV�0��{��s��?O߷�}��߮v�9������ >�յ%�ݙX�(TZ���E�YPW�1�:�dG'��[v�Ǟe�6�^�Cu֘��<�̙����]T�����:���{�+�9U_�]�����~g�L�9�ɭW�?��}��:W'*�[\�*���c��7c� }6<�8��D=j���|WEջ�&�� ��?W+�UĎ�y��{׀I�(��up�F�rx������? ~���,�x�R�3� O
ZK���]۫�l��ǀ~��<�l�V�_o����;֦�al!q�h��"��a�$#.��2��5�����ۍ���6$ �׌��+�m���,{�+ �� ����\E�H-�Z��k �ٕ�H��� =�� �{y#UOz��ݡ��P��������Ü�����pV�{���I߻���>��r�k]]��O���m���π{����7�2�?.��� ���^m��ݧJ�bm���`���W�w�~0��m�O���rӕ%�-�.�4&y�z�6�bN��G�q��qsϡ{B����J���ײJ�V��M���0wc���=x�R��2�M6S-ZV�f�g��]���� ���׀N� J�%-] ��M�f N�x�Ȱ��W��=�+ ��?���EJ�R쫴qYv��r,wfV68`-�RK�R��P`�����>���䓞}�̺��Ъ��m�wfV����_����@?O~xۑ`T�LvS��ӻ�����3��y��8��=�.`�'W]�ލ����P�p�U˫Ht:T+u�M�;��ob�I��}�x�w�����6��x;��#�����'c�~�W;�y�߆��V�餛x��,w\0�I{|�`�y�J+e���tS�Yu��;by߷ٴ�Kı;�wٴ�Kı/���m9ılOs�w6���N���z}��5kT���O8�Kı>����r%�bX��~�bX�'�߻�ND�,K���ͧ"X�%�Eϸ2�D���F 21��b���'�b�D��[ ��pօ$� �8A J���7Zs�ב��C=�vBО��V	2��H!# �&f��%��R�R@օᬶf�Ez�L7	#�l�t �BN`y��0�@��$g�x7j_Mn�)�4p��'dٰS�j!�A��Fx��H����{�'g>���y�=��OʱUUV UJ�U�r�R��U�UUT[R�Ub�Δ�++� EE3�%u�s��k�UwM�&�ѕ��H˥��TU��>.{H�%�Wڦ��!�{N�����e�X�R-ѣ��6.#G���-M+���5J,Cn8S��ۆ:�ʡ�S�Fsm�`Ƚl�	���Ḵ��홖휥�]V1)ջ�ԼA]����܎�;����{j��=�Ӆ��
j��[$�������.;h��	Ϛ��=��9�d�A��g�����\.R��B�,.��rJ�ˌ�x(����
����#;���N�4��;o9�jlhC�B�E��K`֘�ɲf[k���1Up�b�;\7�{\9+Hr��t<<�l�ń�M� P%. ݕ�ڣ�(�C�#��3�ݶXy����كlr%�a�Lr ��}��,���F�Q^�M�)�JE]Jի�5�����P)��L����d�b)�\d�9A�'[P�(C�����cl��'@���/K\zy1���v��t�	��������6��&.�\���n�=W�R�g�� ��]P�Q����W�G:c�U�q��:�YjU��4�W;v���4�v	�����5���T��)��zqe��
�`Wfu�{gPAJp2Ɲd�^�>��im��{��]���"ٔ��)�`�L��/&.�(��j�5��ت]z@��s���xWG s��ưޮ�tdXZ���N�m[.�F�����ꒋ[v0X;j�#�+�:������d��F�d�,PcD��󹮌C����99x��n^�6�]��V��v��\h&��2�ճn�`x[o".���x�XF�k2b@2�QGj�S��h�6�b��Z:t6���0�s�V��a��h�m �vE���wN@Mk��UA�2eaSF�V�ƪ�\��F���X�
]. ��*�+����=�ei�󋂞��{�bED��KrL�[��"	�(UP���Nz���h����S�I�����T3�P�`�|Cf��TA���m
��_P7��R�B�3"X���]<�엞Kvw�R��ܨ@�,tu��t2�@n����{s<�*��J�5[#�-^TZ3&�kM��3)�ɑ���7 B{�7Hs�Z�F�mdҵVx�m�'=v����A:��uֆ�N͗`�:��X��N��c�u�$�����=��'֌ճ�m���AǃF5�9^[T9.RӬM3���$�HwN�ݟ>�1�ݻ]@{;��T��7/Vzq�tg�=�X8�J���g����҆ي���Kı/���m9ı,OsﻛND�,K���͇�>DȖ%������Kı/���'r�̆e�ə�m9ı,O��w6��bX�'��}�ND�,K���ݧ"X�%�~���iȟ��2%�}��?Knd5tS.L���r%�bX����M�"X�%��u�nӑ,Kľ}�u��Kı>����r%�bX�����ִ\2�2��.�6��bX�'{��v��bX�%�ﻭ�"X�%����ͧ"X����o�iȖ%�bw���[��ֲ�jY��f�6��bX�%�ﻭ�"X�%��}��ӑ,K��߷ٴ�Kı;��iȖ%�b_$'oٝ�U�b�u$%��,܀0*��چ�tC��Нe���t/����i���T2[U�å:S����{�ND�,K�~��"X�%���}��,�&D�,K����ӑ,K���?~ɘI�I4�0�Zͧ"X�%�~���i�mT�����LGo"dK���6��bX�%���[ND�,K���6��bX�'{'��S�ur�5�f���ҝ)ҝ>��ͧ"X�%��{��ӑ,K��;��ӑ,K���w�iȖ%�b_��~�}k�f\l�t�t�Jt�O���siȖ%�b}��siȖ%�b{�۴�K��;��iȖ%�b_��K>���r����m9ı,N��m9ı,O}��6��bX�'~�}�ND�,K��{��"X�%�ބ���H�V�F�\m�K�������{�"����su�ܶ�xJ8��\v���g��bX�'��}�ND�,K�}�ͧ"X�%��{�����"dK�����y��ҝ)ҝ?i���W3lT-f�SiȖ%�bw߷ٴ�? �G"dK�����r%�bX����ͧ"X�%���fӑlK��l�˭k5�.�,�fe֦ӑ,K���w�iȖ%�bw=����K��u^�G"r'{��m9ı,O}�}�ND�,�N���{�5��s�f���ҝ,K��{��"X�%��o�iȖ%�b{����r%�`~dO~���iȔ�N����'�����c*����ı,O}�}�ND�,K�~�fӑ,K���w�iȖ%�b_=�u��Jt�Jt������F@*K��z�y���v��v��u�ۄ�V:q��l9�Mf�֡���e֦ӑ,K��߷ٴ�Kı<�]��r%�bX�g�w6��bX�'���ͧ"X�%�|�-�ouu��34\���ND�,K�u�ݧ!���2%������r%�bX�}���ND�,K���ͧ"X�%�~{)o���nf�ӑ,K��;��ӑ,K��߷ٴ�K�ș��o��r%�bX���߮ӑ,Kľ��v[s2ɬ�̙sY��K��"}�y�m9ı,N����iȖ%�by�۴�K�����ͥ���I'?T�[%��������	�Ǎ ��O5��ӑ,K��~��f.��,*�t�t�Jt�O����Μ�bX�'�뽻ND�,K��{�ND�,K�~�fӑ,K������uT�I�sÊ׍.�Z���X�*a%xX7;Sc�EI���L��iD���D�,K�u�ݧ"X�%��w�ͧ"X�%��o�iȖ%�����s��O�Jt�Jt���S]�*dB���Kı>�����?"dK﻿�iȖ%�bw����ND�,K�u�ݧ"X�%��a;�3	3��m0�Zͧ"X�%��o�iȖ%�b}��iȖ-�by�۴�Kı>�����Kı<��;N]M]h�5sWZ�ND�,�@ȝ����ӑ,K���~�v��bX�'���6��bX%��o�iȖ%�b_�~-�fh�356��bX�'�뽻ND�,K�{����O"X�%������Kı=�wٴ�Kı �	��q;��=���]����2�:��[�]�U��dͥ�iV�l��:�b��<lc��
�l],�Q%٣�F���my;z�n��S�GJ��d.а�-�^s�fo3#�me��ɘ�ۚ�E5�I�q��I�X{vwFV�8ێ�v����gi4�ǘ���%Tk[3i7Es�#;�����c�'�٬!b!c���L�sK�Am�r2�q�G\�wܓ���}�&$���F�J�Qȡ2G3�m�s�9�u�.��%���m�,�ηA��8,�m���j�=�bX�'����r%�bX����6��bX�'���6'"X�%���nӑ,Kľ��v[s&j\��Ku��"X�%��o�iȖ%�b{��iȖ%�by�۴�Kı>���iȟ��DȖ'p���.��.�ۢ��SiȖ%�b~���M�"X�%���nӑ,h�lN��t��H����ͩ �'�}���fff\�n	"v'�뽻ND�,K�}�m9ı,O}�}�ND�,K��}�N)ҝ)�����m6r�r�|�Ȗ%�bw�ͧ"X�%��o�iȖ%�bw��iȖ%�by�۴�ҝ)ҝ=���.5�׮öiu˳�yͶ��#G �gt�쥄4s���N1l>ֈi�F��m9ı,O}�}�ND�,K��}�ND�,K���͇�	�L�bX��w�6��bX�'�C�!���ɪj���M�"X�%����ͧ!�<��T4�'"X��w�iȖ%�bw=�siȖ%�b{����r'�A*dK����?j0��)���ND�,Kߵ���r%�bX�Ͼ�m9�@�ș�~�fӑ,K����fӑ,KĿ=�ϰ�t�e��35�ND�,�*,��~���r%�bX�}���ND�,K�{�ͧ"X�%���nӑ,KĽ���2\��L̙��m9ı,O}�}�ND�?(eL�߿o��r%�bX���߮ӑ,K��;�siȖ%�b~����cD�D����[ŗ�y
ß�ع�\�d[�m��ٱ���<�{muN$.�e.{��=�bX�'����&ӑ,K��=�siȖ%�b}�����Kı=����r%�bX���;�fk!K�2k0�֦ӑ,K��=�si�F9"X�����ND�,K�o��~'�2%�bw�w�m9ı,O����ֵ��5��s&�3Y��Kı>����r%�bX����m9�},���"C L� ��O"k}���Kı;���m9ı,N�;/d��䆛MY��r%�bX����m9ı,O���m9ı,Os��6��bX��;����ND�,K߈v��!s�T�5sWZ�ND�,K��}�ND�,K�u�ݧ"X�%��}��ӑ,K����iȖ%�b{�����*mӱ)jr���ܜj�y��C�&��ܾ�d��ρh�nM���[n��m��D�,K�u�ݧ"X�%��}��ӑ,K����iȖ%�b{��iȖ%�b_��S�/f��,�����r%�bX�g��m9ı,O}��6��bX�'���6��bX�'��{�ND�,K�ߧd�,�ur��2�Y��Kı=����r%�bX�w���r%�bX���m9ı,O�ﻛg�����/'������jP����,K���fӑ,K��=�siȖ%�bw;�siȖ%��<"��!T��n'�ND�)ҝ=��ɽ��%�����y��ҜX�'��{�ND�,K���~ͧ�,KĿ}�����bX�'~�}�N)ҝ)�����v��a��e����f۪CP�e%�����+6�Q���G8�vm�:�y��ҝ)ҝ=�����Ȗ%�b_}�u��Kı;����r%�bX���m9ı,O����a�o2m4LֳiȖ%�b{�۴�Kı;����r%�bX���m9ı,N��m9ı,O=!���c_�7.o�>)ҝ)�߿|��D�,K���ͧ"X�%����ͧ"X�%���nӑ,Kľv�[7��2˲y��ҝ)�c����ٴ�Kı?g߿fӑ,K���w�iȖ%��wQ?w�~�ND�,K��$��w]Y.f�ӑ,K��{��ӑ,K���w�iȖ%�bw�ٴ�Kı=�]��r%�bX��� b��H�B���Ht���}��C[M��������՗G�8Y1-��p�p���8�(Զ8KT��@ <o\u닧SY�HGa���ţJ��r�YC��NLv^�G��F��Z�snq��v1S6q�;97\�2��a�q�P��&f#\=�"ki6q0O:n�[3h�x	խ�[��WDR;q��� �j���Dt��n��-��˪���s�y#����Z|N���CL�w�����N$�y��Gk6Q�J�,!�f:ql�;V��&N�a����l.��fcn��d�ֳ��Kı>�]��r%�bX�����r%�bX�����9ı,N�~�m9ı,K�߻3Y.��r�V�&�WiȖ%�bw�o�i�~�DȖ'�k���Kı?g��ͧ"X�%���nӑ,K��ٝ�&�k5rk3&kSiȖ%�b{�۴�Kı;�����Kı=�]��r%�bX�����r%�bX��5�u���Lѫ�2j�j�9�ș�����6��bX�'�k���Kı;߷ٴ�Kı=�]��r%�bX�};/d�2K�FJa5�ͧ"X�%���nӑ,K��~�fӑ,K���w�iȖ%�bw;�siȖ%�bw�ޙ�f��wc7;/�8��%��T\Y��v��g����n�bꍔ�R7I�9V����ı,N���m9ı,O}�{v��bX�'s�w6��bX�'�뽻ND�,K��a0�L��3E.f�ӑ,K���w�i�x������,ddIc�Ttu�z�'�,Os\�6��bX�'�k��ND�,K��xm9ı,K��%'ӹ�����3WiȖ%�bw;��ӑ,K���w�iȖ%�bw���"X�%���nӑ,Kľ��l��.]Y�3&k5�ND�,K�{�ͧ"X�%����ND�,K�u�ݧ"X�%����ͧ"X�%�{;�fk%ђfMj�D���r%�bX�����Kİ������i�Kı?g��ͧ"X�%���fӑ,K��9�ߌvN׍%���AG���ycr8x۬��n�v�κCp����t�zt���Ȗ%�b}��~�ND�,K��{�ND�,K�{�͇��DȖ%���߾O:|:S�:S�ߣ���;Veaq�����Kı;�}��r
ؖ%��u�ݧ"X�%��{��<��,K���ٴ�Kı>�~����-�%0�ֳiȖ%�b}�۴�Kı;�{�iȖ4]�`2�w�f��,1��n��E�ju�]�I�:�&��Z��L��b@� B�$�"BJ����R�B��!����)2�[��-�),�JB�(�!
��$��d� ¬0��R�d$��,�#�͐�HJ���HU���N�3�IBP�V�kY�.@��ٞ�n�i��o$��|?�,�C�a��1&J@7$d��G
�p�
�s��75��ܙ����.�P�ɕ8��Hn	#�Rw)C$)�&dB �։0�RP�b�,��0�J��(R\a+�Q-<N^f5���9�t m����Qe-��сu�	e!	YldB�����k!C�rkT�D5L�� K+,Im%V
@O�����A",�;Tj��� �c>@lW@�����P
���"� ��O"f{�ٴ�Kı=�~�m9ı,O~!�	grsWX�5�3WiȖ%�6'}�xm9ı,Os�w6��bX�'s��m9ı,O��{v��bX�%���aҚ�K3D5�Ѵ�Kı=����r%�bX�����r%�bX�{��6��bX�'{��6��N��N������J�����&�e)*0�q����wSe�f��c�4:f%��]1��sY��Kı;�����Kı>���m9ı,N���m9ı,K߻�m9ı,K��w&�ML��3&fL�k6��bX�'~��6���DȖ'�����Kı/�����"X�%����ͧ"X�%�}��t֦���Z��SiȖ%�bw�o�iȖ%�b^���iȖ%�bw;�siȖ%�bw��iȖ%�bw�wV�Y�3��j�t�t�Jt�K��}|��Kı;�����Kı;�wٴ�K��4Q" *�"H¥�i@�� dS�QA�'{��v��bX�'}��sX���t.(��O�Jt�Jt�{���r%�bX��wٴ�Kı/{�u��Kı/~�u��Kı/����B�A�lG[`iC6&q��HGJ�$����Q�ǥ{Jm��/l^��Y��"X�%�߻�ͧ"X�%����ݧ"X�%�{��[ND�,K���6χJt�Jt���=�/PuT�D�,K��{v��bX�%�{�m9ı,N�{��r%�bX��wٴ�O��S"X��C/�.j�dɚ!���ND�,K�������bX�'s��m9ı,O��{v��bX�'{����Gșı/Oߩ�_�WF�,)�.���"X�%��?~��ND�,K��ݧ"X�%��뽻ND�,�ș��ߵ��Kı/{��K�ї5�us2f���r%�bX�}���9ı,?G����v�D�,K����m9ı,N�~�m9ı,M�Sě�d���2nV0��SHP�a�aD�G@$��]��kV�RPn���^j�ڭrr���Y�`�p']��R�8���M2>��p<�/HNe؃���`5t�����HK*DwUH40��J������E��ѵa"�s�[Vqt�=��n�3���%�pN*�C�.�0��k��{fC=�Э�cu/;@V�71��l�uD��=���n6�QP�̌�t:6����e0���p����'I��'�
y��pb�"\�X:n�{�#fN:3l�աɸ����X3��P��[V�J#��l����/!y�ߵ�nӑ,Kľ���ӑ,K��w�����"dK��u���r%�N����|��\�fb���O�Jt�,K�{�m9ı,N�~�m9ı,O��{v��bX�'{��v��bS�:{�{�ں�e��E_:|:S���w��ӑ,K���w�iȖ?�a�2`@��}�v�D�,K����m9ı������	3	��i��fk6��bY��ȝ��~�ND�,K�����r%�bX�����r%�bX������Kı=�>�I{yu��6MMf�v��bX�'{��m9ı,K�{�m9ı,N�{��r%�bX�}��m9ı,N���grMY�.�e���kUs&�݌�Vy��vwr��c��
�I�z�lF�kvD��'�����*_{��iȖ%�bw;��ӑ,K����a��DȖ%����~�ND���N����������b��O�J%�bw;��Ӑ���B�@��$�H0* H�����$
5(T��\����oJ�wqС�
�H�`��%~�*���r%����&ӑ,K��~�fӑ,Kľ���ӗ����/!���@;(&��w��ı,Kߵ�ݧ"X�%���}�ND�,K��{��"X�%���{�N)ҝ)���}��cfL	vo�>D�,�*�ȟ�~���Kı/���[ND�,K���6��bX�3���Ο��N�����!��b��e���r%�bX�߻�m9ı,N�{��r%�bX����m9ı,N����r%�bX��	��3�V��1`<v\��:W�n�I�K]-Tq`����3�"miU�s�°���>)ҝ,N�{��r%�bX����m9ı,O���m9ı,K���bX�'����%欗&�L&f�iȖ%�b{�wٴ�Kı;߷ٴ�Kı/�w��r%�bX�����r%�bS��g�|��랠���>)ҝ,N���m9ı,K�{�m9�z�$��$ZUS��N�]��r%�bX����m9ı,K罇u0֮�u������r%�bX�����r%�bX����r%�bX�}��m9ı,N���m9ı,K�{I�;-�IL�fK�kiȖ%�bw���iȖ%�a�X����m<�bX�'�����Kı/��u��Kı;�'�l��GYX5
O���ʗ�C��ynL�s��2;l5�9m��q�RcWKGK�N�Ȗ%�bw���m9ı,N���m9ı,K�{�m9ı,N�_{|���N��N�t���Q�;7�ڛND�,K��}�ND�,K���[ND�,K��ݻND�,K﻿O:|:S�:S��~�j��f.���jm9ı,K�{�m9ı,N�]��r%�bX�}��m9ı,N��zy��ҝ)ҝ=�=��ܹ�ΆaMkZ�r%�dP�bw���iȖ%�b}�wٴ�Kı;߷ٴ�K���?�ՈA�!�Qnw^{~s�5��Kı?~�{���D̚m0˚�ND�,K��m9ı,N���m9ı,K�{�m9ı,N�_v�9ı,O�����WXh$�D����)bsD�cx��5�T!���Z�)b�[�r�@.K.L�a2kY�'�,K�����6��bX�%���bX�'{��v��2%�b}�{ͧ"X�%�}���i���\��Ο��N�����iȖ%�bw;�siȖ%�b}�{ͧ"X�%����ͧ"Af	"w��#�ZL,��3I�$�~���6$�H����M�$O�;߷ٴ�Kı/�ﯝ>)ҝ)�����IV.��gk6��bX�'�w��r%�bX�����r%�bX�����r%�`؝����O�Jt�Jt�����k�vnJ�'"X�%����ͧ"X�%��w�ͧ"X�%����ͧ"X�%����6~c�L�bX���!C�0�*���w���pb`m��s����t&�Bː�Y��8�s�6L�%�pKB�� ��Ò�d����i�L�y��Niä����L��oSWu�z�.�p7[�8vj����"�s�]Z��6������)�!������*L�Q�M;�cue����%#(���a�^Q��S���;P��4Ѱ�Մ��O@������9^�M;����U�_w����c��z7DS�=N��5����1��&��	�y���`3%�&�h:�S;#.������^%��~�siȖ%�bw;�siȖ%�b}�wٴ�Kı;߷ٴ�KN���������H,%Wy��҉bX������Kı>����r%�bX��wٴ�Kı=�����O�S"X�}߰���%�M�5��r%�bX�����ND�,K���6��bX�'���6��bX�'s��m9�)ҝ=���=f����*�t�t�,� �"w��~�ND�,K����m9ı,O��w6��bX�'�w}�ND�,K�û�gn][%ֳ�����Kı/��u��Kı>����r%�bX�}��m9ı,O>��6��bX�'��v����Y&f�ïW9��8�s�\ϭ �T���Na�S�P1�F�E��aw���B����g�w6��bX�'�}�ND�,Kϻ�ͧ"X�%�|�{��"X�%�~���J,]2�1��:|:S�:S�߾��!����P'��"y�ߝ�fӑ,KĿ}��iȖ%�b}�}��å:S�:}���F��9��\ͧ"X�%��{�ͧ"X�%�}�{��"X�XdL��;�ٴ�Kı;��?t�t�Jt�O~���ns6GWl�Z�ND�,���~��[ND�,K�w��iȖ%�b}�wٴ�Kı;�wٴ�Kı:{����kY�ɣRkD�Zֶ��bX�'sﻛND�,K﻾ͧ"X�%��{�ͧ"X�%�}�{��"X�%��T=�߿K�)�b|g�Ċ�7b�t��y綂%�͂��g���*�bWA����Cg|���bX�'{��ӑ,K���fӑ,K��;��ӑ,K��}�siå:S�:{�}���:�"��O�,K���fӑ,O�Tȟg�߳iȖ%�b~���m9ı,O��{vχJt�Jt����i������J��9ı,Os��m9ı,N��w6��c�z	�JCb�JLTրZ���U�m�ϴ=,M���~��r%�bX�~��ӑ,KĿ}ۙ)�\5�L�f��WiȖ%�����ٴ�Kı>��߮ӑ,K����iȖ%�b}��۴�K�)����u��L�2c9�t�t�K����nӑ,K��{��~�O"X�%������Kı=����r2�)ҝ?���c���K3ZLZq�氖ib�Z�KYF��G4�Cv��Sl2�c��]d�Mj�ٙ���Kı=����r%�bX�g��m9ı,O3��6<�bX�'��{v��bX�'~�d�f�l��fy���/!y�w��Ϝ����J�L�bw�~�v��bX�'ߵ���r%�bX�����r'�ʙ�?O���[�F ����O�Jt�K����r%�bX��]��r%�bX���xm9ı,K���bX�'ݝ��s2i�Ւۖ\��r%�bX����m9ı,O~��6��bX�%���[ND�,� 2 z�pr'�{�.ӑ,K��O��o$�5�5a535���Kı=����r%�bX����m9ı,O>�{v��bX�'�w}�ND�,KϤ������\ʴ��y]�)&��j��6v���'l���H�g�Z8�7.y���a˚�߈�%�b{�wٴ�Kı>�]��r%�bX����m9ı,O{�xm9ı,K��˖����f�֦ӑ,K���w�iȖ%�b{��iȖ%�b{�{�iȖ%�b}�wٴ�ҝ)ҝ/��}��0U�las|��%�bX�����r%�bX�����r%��dL������Kı>�_���'�����/'�}��1�h�@tm9Ĳ�$O}��6��bX�'�w}�ND�,K�u�ݧ"X��dO�o���Kı?}ٲ~.L��3WS5��Ѵ�Kı>����r%�bX�{���9ı,O{���9ı,O}��6��bX�&�p�o�\��C4;�Vr4D�1Ù��Ęj�͓8�Sn�R���Ҕ���g6m��d�3]d�ٕ�y��i���2	&HOf�so�D���Ё�� ��fb�_���!��l���A͐ٲl��H>0B��	�e�̉�Ѭ;(I)樆��SF��D���o4BD���n&`j��3MPπ"g�<�I��Mlxl���4�Izp���C!�{�G"BB)}�^����X�d G@y���9-���	Q���o-J@"�&c�g�	!��)#��8f��BV���ў*�UUT�T�]UҳO$�oj�UAPX좬�m2�(���B, ��V�-Y�fpt<L`.	�ٷF�W��[��-tLYQYa��s�S���b]h�͔�w*@ʶ��\å���X���ȧi�H�N�:��۳�j�#q9�j�4IۗV�	A��$��1Fm5��n�N��;mU剦�S��Q�6"cE{�DsÃU�;<�̒��fįW���'P�ۣ���:�"��R��m��"��N�*��s�8<P�IG`�f��Z3�;CF�$,��A��񗖠m[��hMR�AeF��9����snqq��v\V+�6n���ȫN��z_"���t�2=:Җڞ;n9
�ݰ�tV��P�#!���#T�X�c�͝���5=;ng.���a�ZYԷ�n݇9�X[b���I�ݞ��pr����Db�1t�ݦk<b��;�64��L�Z�se��̮��̥�`�hprN긺䋮yy���-4.��������A�f�Z�M�ԅ�3V��k� �@�.�g��y|$��'m��Ͱ�Ni�t��ї <�y�X�mh��D�룁t��"Ll�!Ŷ�KU<��y�F)B�-͑��hE�a�UTV��� �^n�a�@_ ��1�%`K�n��駐���.��˲�;66�b]�r.mV�6���r붗BY��v�Pƚ�c���ժ�'�jD�b��ܗ�HF�+�^�+��"�D���k��	�4����e,یm��]���.Hm�qkv�n��N<زn
.q�<���OX�
s�6��c��[��"��&W�+d7b(��%���z�4v�Es�7;<�P�*��҈���ܛrkCb�x^@�\�4�F"�D*ib�B��:b�@+.��Ob����&�C(ĵ���8�W3l���9�H�A�,�j��Y�X������ڎ '(k�&��u��;0EUGLe�2�����
4�7ZwFܺ.�Q��x�.�M�ʉ��� �>>�+�T���4�a	 Sh Xx|"���g4�99�GN�}M��`D�6��ue�
����^�=:�1]:�;�뷠6^.U�b��v��L�[�N\���K����X8�=(�kô�M���su����A-t���[�M-�p#h�v�7s�k4���z�c�Dq�p��ζ��!�ظެW9'aә��OG�,��L�5ͱ�	�\l�N����N���	v�k9�k�l;-���-�ڽ�i�����y��ZqmJ� �ў����3���`�mp��.W��gXݱ��F��:4h��Y�ju;ı,N�]��r%�bX��]��r%�bX�����~Y�L�bX�����ND�,K����	o.��[-�[��ND�,K�뽻ND�,K���ND�,K﻾ͧ"X�%����nӑ,K����I7��ɩ�,�5���r%�bX������#��)=�0�ʪ��z��`����TeՒڥB���M��7c�6�,��X�X�-Z!˧n��-�� �{�UUs|����{+ ݏ���$��/�H�6f��e�mu&ݢ�Ջv���f^<��g[�v{==�n��MyٚT�ۻ�����_��	�2����s��K�X��^M����m0�������}7���E��s~����>�>� �J��ݦ;N��v8`�ذ��}�� ��wj1][�N�t!�`�ذ��}�� ݎ餺�h�v	+J���0S+����@��� ��/ �����7��bG�^i�a*GK�7��W��z�g�.Ѧ&����6cʗ����f�c��0��r����o��`J�U՞��
ڲ�;f�ٕ�uwe�Mp�>�p�:�K��pm��E����ݗ�}���WI�Utr�`Ґ"PMoY����s�~ٹ�[r�Tݦ]�e���r���+��g���� �ve`]�xʦ�cC廷c�l�>�p�>ݙXWv^�� N�J�`�eX�*�7m[��#�%���@��ϮÌ�FXM�
1֒�t���u+�t���ـ}�2�����s��?}Q�W�I���E�n����r�T������ �ve`��2�TՉ+Jۼ���۳+ �ݗ�wbB�1�ZE;m`Mp�>ݙX���W8NUUt��wN���o�}�����d٘wfVv^�܋ �� ����H�&��M]��l�5aI��%Kɚ�c�!���r�G3�"K��p��.��;�wfV��ĩ�Iڻm7x�r,w\0�̬.��Sj[BuCc�	&ـN��ٕ��=�� ���>�tN+-�+�t���f����	��������� �KQy�SaN�
��u��<��;'������ݗ�ߧ!/{�kef�e�.h�gZ��������7U�����|��{[n�wC�L�ϋ�k �)�����%� $��ډj�p����IE��:�\�Og����)�n׉놛t�\rX�(o6��p�m�u*v�@Uq�K��\/)0Hw���<��"+��r����}?��7}�jY��7)b�6� k�	vd�j�f��ng�&E��X�Z���t����7���)t	ζ����ˏAhRpW��$1�trv�+2c�]�5���Ѻ,_@�ze`u� �n��"엀we$�*��%H�f7\0��x;#�;�៹U\���_���l/���v��T�� 'dxv��ėu� ���R��e���x;�窹I���=���>]���[*�M��Wcj���`��|������Ur��R�����v��6.��&�ݻu�4��*ݢ�:��3ΰd�=��0�p�n�tt��!�_������	ݏ��W�l6y�0	�:?YWM�.��wf]jnI��f�m>U�2X$$�,c
R@i@��"�H�hJXAH�%b�c%��ʣ��URa'�<�0	�p�%CfP��Iӱ*eݻ�	ݏ ����UW�]���T���7����%M1%b�o ���N��엀���*]]�iZ�m� ���s޿�=���;��`�Д��Ӷ��z�7f"w�8m�NxM,��m�BR�l9����r�������/�߻�	�ݽ� ��V��._t;���x;#�q#e�,�?�d�-KeZ)���uh����{I>��}76l��b u�|�/P�(�ﺾo��$�~�[�uWa-��"� I;k�r���T�� 'dx��wu�,�Ӥ��'h-� �d� ���d��>�r�m��M؜�t6@&�h6lX��8j�-� PΠiG�9f�84�Wi�c�'_"VyF��E�.ۿ�7g�6L���-��	���%M4�bM�l�Y+��s���z�0<��x��`gv��۫�ƕ���۬��-���#�&��*��6��m�ݥl��9��qz�x��x���Us�ڤ������97$��~�dϮ]Iu���xݑ�c�ݎ[%����n<��9��j�����<��r�+�r�[u�&L�t#�B�
B���k�<�b�2���?{��`��E�_�9�g��U�<��N��wv� ݎ[%�d� �&V~�8�6:=e]��ջ��Qm���� 6H�	�e`#�%^ʻ��ćN�L�n�?Ur������e`#��^��^��^�-�SM$X���M�+Ԗ����=����UM�w��b���2�gu�G*۷K�9�-��(�B&�u�h0���T�Qxf��N��X6&���v�O�]��ۗSj����N6@�9Qʶ�r��͆2��� ����Ӵ�=fu���4E]��)�s�L80�˺v.�+e���p�h�!�2g*R�=�z�qz8�y�8`ᐄ�X��a42Xf�͎�[t�#��ڊ#=���f�������$��4��`�Ko`�W���!g��G�]�+N�k[���s�z-���(��!e��ەsv�+?�}����"�/ 7d�\��l?{��@��W_�LBm��]� �d�V�x�2��៹�r�:�]�R^���w`��� �{׀M�z���˹���`��~�Q�e4Sm�-U��n�	�� �0�K�5I/ �ȭ�'LIݠ��l�6Gܪ�\���"��x�u������zy�\�P2�4Y����ks3�s���,�7c%�&�̄�eq5�e�wM]ـE�^�Ix��l��Wun��N�
�v��߾�7�<�`  H�$���qǜ�W+�Uޟ{��?RK�>��%l*�I�n�	�e`G-�����}"@K�ʶ:WV��`~�Ur�z{<`S޼-��	�e`iQ����[�V�-���K�&ɕ�M�����,�J�F��I�&]�s֒Q e6�l@eZ����+^0���E^���L��m�=�N���&�.�xD[)����Z-��;�+ �8`we��<��"n�v:�b�X�� �v^��WL�R��/�]U_z<�x�S|��6�&6�4E�BFa&�d�d�$aa#@�$�wWP��46�T��(]�̅%�Dp�J��a�q�<��Hf{k�lh=�M+Đ�Ov{��dϷ�9��x0)r��j�r�l�<�7�Y�sf�3c��/��M��i9�f�w+��%�RML������V�r8�
�C��|�S����O9���4*/�i�|U0�z�>�©T�0�/|�}�y��9�l�Kg�Ϯ�}�lv��5e���O^��	�2�	#�;[2��tSv���m� I#�&ɕ�I0�K�>S`���P� l1#�kqt&����rf6���nC�α��[���`nhীN�e`c��~���<��TW��1�%V��u�M��H���x��<vE��}��1��l�V��RK�	�<v+ �3�H�%��%�J�$�	[n�>^��^���V68`r�]U$��\�Nw�������[z^�v%��1f�m��'t�X��E�/ �d�����^p�Ut�6"YI�o���3��q�����l����vśg������W0�cF�K-��zy��"엀E�^;[2�효S�n��wMYi� ��/?r�\��$yOz�m{�X�ឪ��q#�Q�V��V�v+�]�x��� ��2�	�� �v^���贛����i;w�NԙX�� �v^���J�q��lJ�];u�I0W);�}��w��$�ϧ�7$�1!j ��(�H%����-�f�e��.� :�m���m���yԺ-�f��
׉4t
���㎕bH��z���\�=;�8�eݕy��ɱ@֊��5�R7�4݂k��t���.��V����e����O�c�͎L��ۓN��&V���uk��v��㍻1�'`��;z���Ň������ĭn�<����q�(���ݣ��Q�V�������9�㪷�<���N�*�`�R�0T�8�ò���jJ]nCl5n޻f��&�-97g��V7wv�-իf������<v�� �ݻ�!D�:�����<v�� �l�#�j�v�a˲�m��p�$�Se��<��˷M0cI�v!��UW){����� $���O�Ӻ�'��l����j��{}�� �G�N�� �8`I�+�BÉ���u��'����LG�ܳ�[����(��F;G%�0����6]��<v����s������ �X:��ة[I$��'`ዊ������U_9ڪxfG�6^ M��lE��be�� �0���	�<v+ �J%9mU�V�۫t[u�E6^ I#�'a2�	#�ջwuHP)�jĭ�xRK�'a2��� �l�W�JS�7j�G������P��l�f�����`��!G���u��in�ٺö.��=��l�Se����ut��c�)X�:�6G�RG����"����e���F�GB^�n��wM]�7$��{��{}�����gP�S�Q9���Y�Ok�M��[����j�v��z�U�JOy��{,�;#����f*t�$����Nɖ`�0���}��`��ux;wɻx��.ݔ^�xj+���\=��[s����Z����B�Be�:1H(���>?O �Ix�v^;&Y�N�FKj��jݺ�l�"�^{�Rz�o����\3�H���^E0MX��� ����,���RK�5�]�-�wG.ʷn�=�������6G� ���ٹ<_�Z���~W�y��`ZK��j�e+�Xw\0���|�K�'dYX��
��P;ެv渘X�s>9�vwL��۩�hG��  Xa�t	t-x�v[�)�o߿w�|RK�'dYX�`j8]�tS�M�S.ۼ ���n���M��$��:t��.ؒb���M�X�a�K�}��l��>؊)ƚ�;(m��X�`]��wc��K��}��������ab���:�%������v׽x�`s؋P����Em��u��f��n(^�-vY�Mn�.�u���#ղ֦K�Ƭk�r�c�:^��0�j��;�����j.���tᢕ�^i��<�[mt���6`�ЅAɲ�6�89^�^�΀�>M���5��zvvwhD�8k�(GJF1 K.ĳ���5��S�8݉�cp���~�>�b��Ӊd�'d�gUs����SB�P�Wmy�gd��3O6��K���YTa���b�!g�6w����4vNGh����m%��![�r����ߟ ���^;�����W�� �7�j��n�]��o �oc��r�=���5Oz�vG�ut۸�Ut���R�v��&� wdx;#�>]��ݭt%(-�vڧvـ� N���do�M܆���v�����ڶ� I��.ˏ �\0]���~>�G�/6e�m����YėqfX3�گQ�)����X�+u�<�B�Y]��|���	��Eݗ��<�e:LN��M�M�7\3���圢s�����,-f��� ��g�ĉ
�'��+�Wct�;f�׀�<�^ŀM�WV��r��&�J�w�ݏ �"�>��������<��Z�y[G.�J��>�r,���x����*�mQ�O��wc��9��t��i�N4r]��K�+�:8�Κk�eDҶ;Xp����_O �ݗ����;Kb`M��)`��j�-X[f��W{��}R�,�0�[3�vʵm]��n�[��I���ٹ�Q� Q&���l\�y��>[=x�d�WWi'LI:w���[���p�>]�x���K�׀vW��6��]��;k �G�U�����[=x��ذ	R��*Ɔ �X�G�S@Q	�a���.�����c=	�$� V�.&L����X����v^��/ �Kذ��`�K��k��V%v�������� �k��/=\�H�7�wez�uh��Z�x���}5� �l�Wv^���K�e�j�ڢ�0>�Mp�"�/	=�{�nN�Q:)��9����ܓ�����N�j�-X[f�x��v�\0	Ū(��o�����I_Q�2\���z� �1:��������Vs��y[u�[.�鉷x��v�\?wt�C���w��߳іjMF:ц]�N��<��G� ��z�]�x�QS��M���N���]��]�x�¯j��۲Ս�`�]��]�x��\0����.+\umX��� �ݗ�N��}5� ��^��9�Ts�9����4���$�zI�	���	��<OO��$�/��������Y�����$p9�jl�Y�ȑ�H��
T�!���%�9�9,�C�Zy��o��n�~s8�R5%|#LׇT�+�y�o������$My��� ��q��%�h�h����`�VQ��/��3�	�zfh�sS5�+
8:����׾W��eMs4���P"�����]x�y���!xq���7����C�cO��=ܼ`h`FV��!		�u A�t��!���4�ˣCki���&	�)<����і]��Hi�ϔ����l��P7O˓ �S-y�קƴ��=5�Yx�8hxʔ�0�B$b�8�}���@�1$2*xӥ&�%�<�f�d%�}�y�=�P�����>��6nց�R��tw�`Be���y��n��n����!�Yy/,���~�^^H~�g��UU���PʵUr�U�nU�PX좩5kP��3��]p�K�p�]�z�/�\��:6�#�d	E��l$Ԭ�ĳ$���p}c��s�;N;P��.h����Z�^^��^���sW���`h]���h�ݸ�-��ٴ�v�7B5e�4���E]�fJL�e;0H0[���Ilr�M�h"���<l��
����j�g�]y7nC�1<�'���%	y�����۠�Ʀ�q��BMm̤�]a�dN1@v���=�Bz��:k��L�f������a�u�������;s��:��\K![T�uG!,�)��b�����D���Ӵ<ی= ��n�U��h���@M�L��Y����j\�/n8�65�1���g��'R�l�+nd�E�CJFk�\�8��%�0n�6q/_/�_%-�. �lb�V;���I��0!�61��x��u�1�����N��.�e�1�8V	��1c�4�ҙ9 �������{�ZM�l��n�� ��*��X�M��\��K�5��+��������"Î�i��Ω��8ڝmch���a,4�hŹ��!�c�Ż6U���⓶#t�qg6 �U�ce �����cv�m˼�F��N���WՎ2om��5"�Pt��TTZY�m�e�#�",Bi)tm3ʗ ���-[�S�]b�4"0�M�5�m�oET��w*��l�Z}
�N2�2�T�pn��ʱ���㎞՛Mt\�h�0�'c�踃��ck�؆.c�3V�@�S����v�
��g��3���M����Z�,�Qe��)��4�R��c_1���c:9�ѭ��N�Q��inq�����Sfk+s�#jCVBlL #�l�mvx�g;
�k�F��5���k��7��������	��ct�5QXG����-plJ�L�geQ���-`%`��婨i�V;U]p��ù�D��f���$���RʵT�=xj���[l��t]����s�5�c4�~�=|� ��>E:"��;<W��8�mq`����|��l浭K	KK���Ys5+���Y���5�&�+���hM4%�a	��1RM4��]2�
��|�8ח�ɻ��gs��=4� OM�:��6"M��6��p��2'7����mkB�]ck0�Ɋ�nܒ=�@�
�dtJ�D�Ԗ��c 6���&�hl/\s��ª1�iq����5�M�y5���R�W3�-�5��0L�?˝�������[�7�C3h�X[4�1�/�gd�b�n�V�``�96��0�K
,��ݎ�6���������X]���p�;K���մ�T��[M`K�`vK�7u� �֢��J�t&�j�-X6�����ᇒ�Ƽ����I[3�m�ۧV��ۼw\0	�j,�0�%����tՅ�i!�v�wZ� �G.�x�`H���3[�q�	䋮7@�o@��P{@���ǃ:ec��f�h�Y����Dr'��{׷�"�/ ��v5�U�\����������y����Y&�*����z����?�R�+����`����p�ܮr�ʤ�Z��Q~V��ڱ+�� �?�j,�0���";*�ʖڻK�`+f�T����w���"�/��$��'�[I5I�E��X�8`M��n�;� ղ�);L����3��Q���i������%�fK��%�Lbf[��5
�&x�ܷ�oN���7u� ��E��>A�y��=��*��n���16� ���*�T���^X}�� �l��9T��r�΀�,N�Htݳ ���,�0����"�TW*(��� @OE|�W�?f���`ݨ�*�[Ce�i�m5�}5� �l�?s�M��{|ז���#�V�+��lk �{��� �Ƣ�>��vPTS�YhL�ݍ��1����z��Ƃ��{^���9�!����w91*amX��� ��ŀN�Q`u� >��t�wu-�v�.��k �u���p��G�onE�m)�ժm�vQe��ٮ����Ȱ��E�mm��b�)�o�]���K��x�����K�_W+�*�T����ҫ�?(�@������wj~W��LJ�եN���Ȱ]�^ٮ���.�J��&����f	[Z�)�چ*�W�'�N;;:�����:��U%��`╈5o�_����p��� �܋ >����-:�E�L��xf�gꪮ$���	��,Wt��l*���U�J�n�b�`�G�onE��.�S׀zG� ��.҉*t$�V�N܋ �ml�m�X�����*�Զ�.�h������&�ŀj엀E�/	:&Bt�H�%@):t���ѴhKv`��c� ͇��^�F.��NM�3��GEIx֤���jv1��-e��h�Ҥ�XXsR�Ф
	95�u��nJ�[�'�P�8��A9��)�F;M�1"����yZx��ҥ��rm3kA�G�c��s91���\qR읎�k���.3���NWn�spv�kc�H�&.��`�#%�m�qHd�q.�;4����X��U�߽��;���WUpU�y�j�՚��4a���M@"p���khO
�)�Q5l�u�x;q$gύ���ۥ�L`�SV���w�����X��x�Ȱ	���kn��)L��un��5l��⪒=��,�׽x�س��q �Θ���*v��[�^6ԗ�M�V�x�\�:Uwh��M�m�/ �����=ʮ����o���(M�1�j��x�p�5l��N܋ �jK�;!N~v���57/J���f}=��f�QF�;�ݻqnrE{>���r�'k�]]]��ղ^;r,m�/(	��j�R�X�� �n���"��Ug9×��UR�Y�{��=���5I/ �+��]K-�_.��k �ԗ�M�?r�Ģ�������$�n酴˫�)5n�	��j�/ ��6ԗ�mm��bD�Ro��Zl�5l��z�����_���	��|����q�|,V����ׅ���(ў��S[<"k��y1�vq���4s���a��on���߱�x�p��"���|���e�@�k �jK�&��d�v�XRV�
%�];)��V� ���߾��#���,V��Z$x�3�p�� p�}ߺ�ܓ����'�C�8ڠ�un��Z�`�K�$�m�/�s���0�*�W�J��[�Mp�$���	5� �6^ }�/�����؎(���u��K厓�sk�nm���α����]��E��v	[0	-l�Mp�5M��s��~0�/4�t��
���V� ��,�r�"����~0	ذ��-V*R�M�4�ݵ�j�/ ��,R�/ ��, �kE-�5m�V�@�X�r�����z�	JO^%�X�(8����<��}��s��>�i��m�N�����e�/b�>RK�����o諒��x�!tw*��0�����ò��ݵ����f�+���`]T�qf� �X:CM�v���,�$�T�x��ŀv��MRhun�ݗm`)%�����	R�=s�=�$o���.+�SISI����׀mm�Xe�X�IxQ]��V�)r������ 콋 �I/���)��X��_�2�+v���'m`ob�>RK�'c����`���UW
9ʪ��	D�F0%�x� �l��)̪�՚�c� z�qʹ�dئ�99��O�2�����ˍ���բ#���-hw=���]kFt�Q%㚸���uI1<�¼`�a���զC�ktS\��`�૎�V����Py68͗�l���b6��M��@��8����M���gNN�X�kt��x�B/�f�=���
���&.��g4t��l�̺�au>��Ϲ�rI|g�� 8�������x�n=��ZWG]��n4���ج��k]&�v�د���m��?^;0����� ����]�ZV��I���'c����`ob��� ���_J����`���ŀM�� >�<v8`ojR
J�h������, �H��p�6��,aZ�-�V�+i�ح������mm�Xf�`�n��n�KA�&�R[�%u�u[�&-�2����x%@�O#�ѷ+����Hݫo�&���u`�рf����WQ4��awn����;UʧB���T?0rk�דrIϻ�n����)"R��'T��݂�\N��'��l� �6^��ذ��%�E)Lc|j�M����Se�����UJzg� �y:e��cO�;v��l��Q�/���� }�< � }���� %�B� 5���8�(�Z�ugM���V4Uu�M�Wo7����� ٮ������
��(�R�(��v��\1Us�H>�<T�x��Ŋ�#���"i5N����V� �H�Se��G*��[�NsPtP�[I�\H2	#c�]i��ӄ%2D2G ��v�C7���g҉�"m�!(\#`�)S 	�f��.U����:MT�є!����� 3E4���H��D�Ƀ���b�Û�5	2��C"�F��D�"�����f�h1��j�0��h��kAO8J��'��3O2,�w̸��b�����M��FU��j��_h��h����;�!yF.�O�;��W�����0�����426r�g�Cȃ�R���_B����Lf������5\�9��M�*lu$VA&Q�j��xV��F�ɬ�fB���Q�1���A)Ë� �4� ��3�Bń 113(5fnT1+��
�;�:R+�DC�M��T
|�qR�� 4�!�"/��{Oy�Dtl�4��(�"}�O3�_�r��{��rO}����iW\��'_�߾� �%�,f�`{��).��x��X���؅˰��x��ŀl� �H���������wla��ÙBi�n7�J���v-�^�n��.7W�۟afy炢�f�].'m`k� }$x]��\�9U�	R�%ҥ.���J�)*I� >�<.�x��ŀM� �t��ڵm�-��۶��%���� ������q�m;C��������`u�ܯ����u�r��8�p���dG 1#
/ↅG򃇜����O߾%��;��G�Wm`u� >�d���������z���Ye��i���vKp�E�u��t��mb�(3Xj���,sh�J�cuj��g���%������r�߾�f��N��df�L��f7�E�/=ʮ$mO?�?ݑ�T�{a��p��Ӗd-�sY�'���L�\0�#�5vK�6��wn�n�ի��m���^�y`�y�� �lp�7n�-��t�n��'m`vG��<��� �{++�p�Ho��}B۳�J���DIFXX`�-�1�DŘ�L$K'�^�ٱ��h3� ��p�cm���]=��M]��&�H����!���Ҳ�����u
1�����͘Xhq������a�`�\}�D�Wa�`]�G�4t�9�S[q����e��"W��[��m����w.�ő�4����uqrF]��	��{Z:[;��Gb�*���j�!�;��t���'$�By���R(J\U�R�&�<�I��
�6ap����y���q+9����vZc�|M�m��O� �H�v^��_ $�����unӴ;i m	��v�p�;5� ղ^ ody�q"),
^�t�f����d� �����aFӖ�V:VX�bl�:�K�� �lp�;5� ���)K���X�v� 7�<��� �� ����Ex�4�m���?ut{}�,�'SF�Mpi6�`�YV�)uD��պT�%��r��}����p�� 7�<R�Q]2��a��nkSrO>�_M����H@A�d$G�>T���I�y�$�}�<�#���*R���;i	!6|'��{#�;R8a�R[�X$U�V;-1;|�۶�{#�;R8`���<v��-����6�Ԏe�X�G�����}�ߛ[(ي8�P	T��FJۥVSc�u!6��<��ɱ=�=��y��ɔ4p���>}� ݑ��G�v�p�6�F�Q��իwb�`� 7�<�#�ٮҋJZ��L��v� odxjG'9ϹY�9�D�P��(����u�nI<����V�n�-ՉU�ZV��mKp�&� l��� ��B_-���ݪ\VـM� �#�	��޽�[w��k�X��v55�dO6�9�0�ж0��\�v��wcr��{d���sn�n��$ـ$x;#�6�p�&� n��`��|N�m�� ڑ� ���G�okS�v;v�aE��o ڑ� ���G��<�v��Z-.�6�n�`� N��1r�Qß�
	 ���*� .|k<�nI��2[T��V!Yjـ$x�R����%{��7\0r�U[��{��]���n��}\Yn]�7>�q�C����Y�.:�!�t,���Q�@bQm����|��0	���s�{޼Q�(�x�e%V%i[xԎ�p�5I/ 'dy�W=JD�wVӫ�ݪ\VـzG� 6H��RG��x�y��5h�m\�v�մRT����S���o���0	���*;)�;�v�o 'dxԎ�p��<�Q<�A�2XJUB�Po8^NO�g�Wm)��:���G+Hvt;�n�C�)E�(��R�77^zK:���L��^�AԎD��< ������ ܑ�G�:u��gr�v;Y�����f6�WA\2Lj�(˦���P����)ӱeB�s�
nӴ���p�m)<d��v��m�V�1a�F�����;\���.�N����o4t�"�TX�J⌡*3\��S%���M1��k�;9�s�d��7����R��:�mHMf�͕�ʶCϋ;O<�m����r	���/j+%�lh��I��z�_�m�X�G��<�nJ�\<V��t�f zO< �#�	��#��
6�����E+�.��5l��lxjG �c�>�ZR��e��1ݻ�	�ڑ� &�x�����j�e�9vZV�ڑ� &�x���vG�z��'��t��;�j�҄#q����y-� ��Ÿ����rd���#�7h�n�]�n���O��}�������� ڑ� բ��KWl��\�����~�7��-F*��Z��b�W$P�U3Rw�w[���=�p� ;��}��_�]c�k�[U�_ �����}7^�� �~���z� ~���Z�\���@>�9kI)6?�I$�F�$��c�䒋���K��/.�W {�_} ��I$����$��9kIzz���]�Vd�$�FU�p����(���qD�����	�Hm���9�vy��97
������ĒJM��Kj㖱$��c���e���7T��e| ���$��9kI)6?�I$�F�$�l�Z�雉f����M׸� ;ߺ���I� '�`H�A� @?�I����� ����� w�^��]1q� w�u�� ��_ �����}7^������wF�M.���Kdo�S�?�I-�/BSg���m�'w}�ؼ�&6Hl�rY ,���F��/5q�^YUڻy��u�݂�u��Ѯ�Ī�_@���Ͼ�}7^�� �����z� }k��Z�2�K�
���u�<� ����@/۱<I	ov<�$���E�����\x ���~����c�����{� �l�N��[�l}�mȞ$�[ݏ�Kj㖱%�\�ms��/���X�R(� ���5�`�I�3Y\f`�!H �X0QH"y��ߺ�-��>�7[�\f� ߾��M׸�I%����$��Iz�}���1�ұ�A�xU�S[���.��p<�d��C;�����.ɛu�\L~ ����<I$���$����봒�<��$��T
m�M�8eǀ��u���M�{��I/l���ڸ�I%����t�-�ҙ}��׵� ;�����{� ������z�vq+�6<Iz��r�����JU���$�S���_��� �[_�u�-�����Kj㖱$�{���{�$z�[I%}�뜶��"���DW�*"��aDV� *��5U_򈀪��QU�@
/��B�P�BAdBDDY a	 T$AP�P�B$B EP�P�A �0DX	$P@��/�
 *��D@U�"��QU��
�DW�" *��U��
��D@U�"���__�����)��:N����,�8( ���0���C�@kTv�]hm�   � h t*t�Ί F��+�@ ��ҋ���  ��vΝ�  
(ivP�]�Jmݚ:� �  �Ss�ٶ �(�((  :8�fn��x    �  Q�(�
$�9�(t���9�t7{����=����ڃ�n�i�R�h�}�:��xu��v}�A��¼�� @ -^{��X���3W �n��u�!�����
��}�/}�x=�{�xC��Tmw��� �j���@�����z;�|}Qݝ����F i�`;�K�o��]�t:�Xy=��=>���56|���  =�p<���h}o �>@���<�\����{��s���^`8��@�P�  �gZ5�xۺ�d{���0���3��w0���:q��ݝ�7��`|�p  |�۟a��u�Z:�f�0>��l�����H� �����c��� p�)@� .��ǃӽ�t������Δ
n` .���� 3�A@w4Р����
O`����z{ �� v�R�  s`�� /N[8 t�� 3��@�@��AG��s��� � �ws��g@�  =  �����٥ �h=��i�)AL@�3��' >�R}��.`��}��0޽P>w|�}��  =����{���'�;�wc�:g����
�7�\���C by � ��M)��%H�� Љ�UUOT� 4 �~�J�#�T�h��5SS)U4�# ���I7��H  !JH� h�OQ?��_�����o�̓������}��@_�Z��U Ut� ���U U�TU� 
�ES�?��V��Ia%+s�������s�m�<=�}H�0��E�)L��2�)J�}�j�!?hdbC����s�n��Jň0�m-*I �  �$�G!�4D�!�"D� �b1� B��(h�z��0�a7��{��)�|Ǐ���K�������l�xy�Ӟ���޻�;.�/���"D��"Ra�B�%!�H1�ak��h���7��N}��l!H��h�ғ[׿�]�c!Bၽ��p��B0#L���	`X��&�/1�)�,�!�$HR4!p���zg�U�:]�����K7��,�,�q��,�y�5�m�N�2)RU�peĸ���e�I�,�-�CYYtOd-��$�"� �C���24�5�O�<�1����Y�ׇ��VSP�*A�FD��F���d0���5M�����\�ryh��G�Z�!6Yp�O��vI�@�e�<�/f�GD�	p� HL�2Cit���i�8���䷶2���f��ro'5�d��У/��7�������ۖh�����$�YD����)-�y��!w���F����$�K�\&s\\�f��C�%"�<���i���>�8i��g���y��>��>We�ϳPW����0���{%5�M�Ya�K	�/N�(;���.o|�<�s���n�G:*Ě��ɼ�G9��l�̘ʐ# HE�ge3XI�фHkY�1!rW�y�H��)��w���l���5�2��p�Mjq����H�"�[��fb�"O,��]�%��{u��a�kR�&�^ԇ!H��y�9��	|�y�����˚��k���or����e��A,�$!��f���[�/��<���L�\2�����-�f�'7�p0�\�$��,�M,����L{�4���͐!7�9���Y女o��o��P�HB��]$a�f?�K��x���xXZ��޶g�7;י�l����<|�o:��9,��Jd����������XR��JJ]L7$L\;0̈́
BBj�&�¯5��)�r��i�$2\9)BP���� IB�MJjZP��J0�
F�5�O��`R!C,i���9�7�}$!oI)���
`B�`he������hל��xϽ��%��CX��ẅm��8FT��r0�2A�Yo��0�����8Y	w-�X�*x�,ܧ��;����o�����Nmߔ��̼�uNSRA�2d��%WB�GZ}���to�G0[w�T�u&���,�~\���Z#p%���i&��oLt^8|�������{9Ε�>�{�Me1э5$"������HHU�����gƴO4n�޾�	q�"�0��f������!B9�s���e	0��<�a���4�F�02�L�f6x�����l35�9rBT͛	u�.o> C#q#	�]{	7�5�H@"@�5��&�R��j��I7F�ʰ�$�m��I!��}��{L7�����#F(R�nF\���@��.kdA�I$$�ݞy��N�����C˒K�H���\��a)Y�˄�y���#%$7�v���^a�A��B����0փp3Jl�<����JK���!�
��
��2�Ow��I$.��)�a\�(Bk�j�L=!q�J�	�Eա�=ą�j���0�����Y��9||����	8h&ka7�	盧	|��<ނf�9�Z�4Cf��= HE�_b��]�eL��7��	I�)IL�\2�˭�$�0�B�I�%n��K���l�<��	��u�l֘�7|5�&�y˹9y+&�B�(0��m�׾�k g��רp&��y˞m��v��A5m����9�$��. FS�7��d�Z8R	76y�).l�\���ߥ9���'=��46B"}�!�H|�>.�	}��#<��'����	�J����Rf��4'�q~��C	�.s�a
fr$�6�aL���u�R����K�Y��8K)6{=�.M0%�CZ�"0B����X�H��dd�\���	�4�a.iY��䜰���[�at�iN
�hY�]u�E�e�xR�k~k9����BI姦[��owIB�L�$BcR8�$s�$�3!��@�J�,$�!"Ą.ݗ4JK'ބ�}����P,XH���K�}43E)��H$ �2�
��j����	 F2��E�����:�-9s
��ݼ�-����Rnh4S� �I ńH��k�����'5��|�I�b�'���J��B°�1 a	j��f�BH��*ژJ�		�\�e�6&�����/<�e$a#e!�7o�p���Y.���V��}el�>tƁn��>��3G��gK����7������6K��.���3S���k�B (F�X��LBȲ c �@�)H� �D,�i�i��\���O��+�Yh�siȼ6D�@��]K7�~o�m.��6��Lѱ:K>K�˸s�yb����+ǲ�i/f$		ÖssG�x�v\MM)Hg�$R/��k)rߙM!�S&XCBb���u�S�
`M0�$�%#"D� �Ͳ������9�0�±i�e�f��0�ɓ���������������BÁ0���w�5��L�>��)���o�ۆ�Cr��qO�o���fRGEb�J��л������t���O��Cy���}�a��Å���B�aq�ߚ����&��@�Ix�,3.NKǔ�7#�m�A�>y�7e�,�c�:3�}3[�>�\<`H���HF0a}��od��Y$B	"���71�[�.���W�����	͜9�9��N��~���tI��#<���U��<�Y.��;��֕�B@�!�u�oYB��͜8Gjd	Hy��M�s�ֳ�<5Xq�^a%�a�sÞpނW����s��o� ���B�����p���C�<۪��@�"E�D�B禾��,/7R3\2��(K�B�#���v� ��<޵�j��vH�!VMd�"��@H�R���O7�4KB��w
�ai�$HBKNB�B��!IbH��-��#pi��
A�M<ц�$��Rg'3w���pKXP�)M0�B&!.��p��3�<�Z8s��Q����m7.lw��7=��o!&f�c22�e�%�%%,)X@��������;{���;�^JK|�[�����h��D!�� Sz�np1#���G%�����H��HŁI ���<x$X;w%<�����>xWǼ��/�Д��Ä O�B$��eL>$P��[�:]�sy�y��g
�
Ƅ+��#���9�tC1� D�!̅ra��Wy�ׇ���=YZBщ�KFQ���RKxm�	9�.rU�Jo�&��a�}�5=��ra,ld5��5�3A%p��RY%��BF6f���sdl(@�c�d�D�CF���I	.�N�	��<������K$)�5�K��#6p���I1����Bߡę��jBB�
L�5�$��I.��l���3���%ލ��L*Jr�j��F��25��᠃4���)3���R�2�%��)���:Ow�S�x�e/�Xn1�e	Rs��j��=�i��r5���ᩳS|�$�]R`DeJzRZ�$ H2Bk��2i
laam2|��`@ �"9�i��^��l�BE��(�K!!k�=��O �� ƅ5E�\�$��rq2,�~�O+�g�&7�y���c%HX2I#9w�rk���}W�_�B�#Y!H]y���>i���F�3�j���S�a?~I�RB,<��B^�Ѓ���y��XY����)0��w��c��{��Vֿ�}����Z���]mUU�P!�j2=\#�z�w8��� F� BI@􇤺��973d։�i�!.`B��Ͼ%���m�P��x|���HJ�I�e���M�7.1�M�a�u/�������	��6���ٯ_'<���T�!�A"xm�7@��F�,��B�B�����1�XR%�b����$`�#RP�B� �H\��#�ad��I	%�H\�(c9�f�$H%���cR V2af9�P�L�=�����8��!p�`�#
f�Z�Sd+�!(�1��~9�Ğ4H1#F!0�HCߍ��///5�&����L�vi��HHD"B�7L�o����=ٲ]h�X{�|��i�R�n��153�-���HbE�a!$ ��,Y���k\7�'�h5F���@H0k�	tc��2 �GPh�pT���"0i��*ư�Jh��
r䗀GǶ}�$'d>|�[�̙�����I�F!kc*Q=3k �&^{�C�e~g�!�
Z�g~��E
�"���EY�w�;t��h%1����u�I.jl�m���=��π�N��a(Fg��I|6K������ �N1�~`F!V��L�	��fh� Ĝd��N>�ԯa�x]�@���>vX��<�si��ڽ���gIa,P�$�!R,B1�Xg�� C�P��6��f��]���f���436;�����>�y�IVV�3F���ɽ�H��e�^�{��rBRXK4�����'r^��]��\1�2b���C54a�[o�#f�n��YO5�f�)uY	�v�������٘����G���xC5惡�x˄&��Ya��q�EacB>$+'%�4k{�>2��B�$a�]�}a|9��4��%���?��ӿ`���	�UUUUUZ������������������Z�Z���Z�hZ������������������������;SPUUUT�R��������UUb���h���������j������خXud����Tx*낶w5i8U�.��֭-T��+̾2��`j����d�
��C�Ei����6�2��+�y,J�*ҭU�:*�@n�nR�mUT�Z�V�d����W�����U�UWU�uU@UUUU*�!�īj�k[Q��j�����s�
�.�]������s(MUUUV�UK!5UUUUUmR�T�@n�UR�ڪ�����kg��R�*��Z�+�UJ�ڧm��dX	T
�(�W�w^�� �ҙ�^���8�5�9y$��UV�4��yu@f���Vk1���7c�@��q�ݶڦ�8�6�=m�k;����tf�%��u<�*hV�9�mҬ���v,j�-��%����
����������RR���`��(�S�u�.���v�+\��l�yYJ)b�p<J�g\��@[UmUU)b�U�m`�JEP,
AUYep�"�++�*�
�]o;L���gU������^	���8����c;Tn�y	��,���TGMR���UV���ƥW�ɖ\v��=��ꩴ�ڨ���=J�Ʈ0��uFG�Z���#��
���V���mN�C�ytU���Q�u^��M�UU[lW`�T"�<�GZ�TuxOt�� tp�L��jB�*���NU��m��M[��A���Z:���X���ڞ��-\�waH���쨞��H=���hw93e+s�CK�4Z����Y�eB�� {>}�*{v
��÷[UTH�e*�U��*���X��l��PQ�C([UU]U++]n��*�Um]!8�U�x�UuN�:�d�
*��v	���
�V��TTjj�V����jꪪ�����������Kɶ�����jW���P/+UmUuVC�T�u,�UZ��@T	�b:c�ER���U]Ue[��U� �b��XCf���:0ҩ���U�W@.Q�V�U�U*�i�;U����R��=�PUz�W��lj�U��yڐ��-���RWU6���hM�� ��zV ٭�mu�6�4�T���J�)-�*�R��A�4n7�x��}T�E[����&�C��P�7S�UJ���i� �;%!;TL�Xİ[U��mr��=�AES�Հ9SKm�*�t�שii�On\��Q�����(�;�9들�mq5�zZ����8�U�䋵��݋^sr0ް��d�)uFa��H���:۷@���z�`xm�`��[�q��7;Y%a�f���Gg7e"�%V�X�WCM-�����q��3�-��C{	r�[W`�S�����Wkl�6ؚ�
JCTmtjv��f��G��A)m�Qvn��c���GN�̢������<��Pښ싙)�r�r���
ڠP�P���f��˵UV�L�涥��2��s��
��@i�q���:*��W��󑣦^Wh���9�FN��Yڪ���	��D�lmI��Z�%�c��;��"�.�9L��m�*�������v�ʰ_Q�j�B�B�ꤱ�t*�ή��W=��]Y��˶�QH������Yw�6���2�uY�?uM��\���0��66He�;��qU[+)W�*�����Y��[.�T�Mn*�[¨M�a�asUT���8���$:��i�M�;�n��ݙ�Z���*�tݞ��M��K-p����q�+9��N�ʨQrAB�*��vP9�x��8�!Y����K;7Ѷ�*�р0�?��n��Sc;��[�Y����U*�J7B�=PnV�JT�Tkb�f(n;2�[�P mPu�+�^ѮL�v�j�Bj�]l��^���\(p��#f��[ ��+
������@^�l�.�+�.c��僈��@��M:'�
{"Y�<l��d3�h�C����D��<�S�H8�F��j���V�
\�,v�,*�?��ϼ�U3�J��T���������(i�p@s*�n�[jܬ�]T�v�)��RG@=Ѩ��,�՞"�rղ���Z�$�Ҝr�+;X+Qݪ�:fu��dfK�T�ι 	�]Y�A	���A��n���オ:�iV�"��[��U���gt�N�Z��c�YEs�UZ��l�/`IUX�O�7+�N��9U�ym$:뚣z�@�6�������/��Z���`*�*�-�^v�� �W]��k,�=�����Ǎe���02��-�.�kU������Z�u[����w*�T���xrR�U�uT�`���V�Եtki�6�m�]O<[\���x:�e�Nu�iƚ��iR��7mg�
���UUUUeb�ڇ<�򷶭�
*��ʾz��J�`����vUV��y��L6�.ў�F�@�V�����/:�l�*�!ꪫl܅���D���b�� ]���%[�m��+�����m���A�����TJ�
8�V��x6w<�� ��T�V������X�{����;�5x{v�[�V1�8�١u˓-v]�\�sm;��m�R(q���v�ݓ�ޮ�=5[A������ӌ�m�6��ӹt.�78���Gc�pp��v�R�a�R��v�g�Z���x�y�tm�Sj��WeZ�몪��f�m�[�d����d��r��MK���+kLM��'r��ꮁ��*e�.y�m+�U��Ƚ���UUuUJ��ۡ�b�m��R�T�����*�K���c�9iV�����*�Yi�ZҪ�,�R��`ge�,S�zƸ���crD�F��m5�ҭ[,Q�U�U@##T5T��|��#i�PP*F����ηm��\����%�j��j�JJ�QBe]�I6,�HE��)���k�[
���}�*��vf����j�UD8(e[UVcjҔu�V]
��1�*�ˌ#��v�I�l=5cX��,tA�������u�Acjd�2���7j�+Kj�]�����_R�^�ڪ�݇>�j�S*��<5j�@�
q��(*�������e8��յ�U\���,m�ҩmq@UT�q�e%���q��r�W����E�RZ{*�U^����������j��Wg)��U�^j�ڪ�
�����SU*�U@W\��U*�[UU�m�UTsɺPꪮ�ꪵ!USv_5�R>j�b�YP�
������<��
�-mUZ������ul��ѯj�lʁR�UUV1[mUUUUU@UM��������Ub��\���UTUZ�`,��U�lY"�
��W��j�*��T���j��V�n��4�[V���U@uV���UUmW{���TQP\ڶ*��� sgd��M��h
��U[PUTR�WWU�r��۩V��	�
�[[y^j�ʻ*�� �몪˪jU��P��jjH���㞐X-H]uUSj�h�1��j��������b���U���+UUUUUUUUT�T�J�U[UUUU*�UR�UT��1��oz��:���F�"ܾd�PJ�ʷJ�D�UUUV�Ҽ��Bl"[U\�r��U+�O*pmc�[x�UjUh�B�f� d�32ك)Rڪ�Ut�R�*����P�6vj������s��UUUUmu�nH8eUU�@ʫ��Uj�[�*�0�UV�Q�T�1읜!�n��UU+�2�6�ڪ�V��X:��;5U\UUR�mR�UUT������eUfx*���T[jA���U����ڹ�UTUUJ�/E.ň��E��YS�@�n��3WHHP �W���vjءV��{T8�9U�Zt��61e��'�5*�v;�l�V�K�ÖRS�usuU[l�,UmmUJ��+sWj��i��h�5U7\��j�Ðv��W5P݊���]u\���Zt2��Z�`��@な��L��UUU)[f-�s�u�Y:�(�T	�z��.*�LB�PS��[u�\�61NԬ�u�X'�q[069򕞫"ywiW�΅�ɫɅ�N�u�^��^q��^ظ���uۑ�9{`Ӆ�r%Q[�5�(�Nz�g�c]g5W5tH��K�	�0bڗeP�zT���rvƵ��u�7�e��99.�";]�]Q�v���Z��0�;G��v��[�cϽc�ǶU��tq��W�檙L��p5��I�b����T�l�j���v3Z��Qen�(q��-]UUuU 3��vŃ���qƙfHutm�0dm�.������c�]+�T�<Ьe���Ԃ� @U�SՖ:�n.�I3JUT@KHm2UUV�j�.^7hq-]\�<�5�P]U��.�E\&I��m������4��WKH.Q{U�V�*������ q����mc1ca� g �����^(/�ث��j���X+�����b��y�j����e������m��ԍ@*�UUUPJ����������U���B�fUUUUE`[tHVj�n�������[[UGsTjj�Uj��������Z*U��*�
���������������U��j�����*�����*���RZl�UUUUU������ڠ*�NeZ�������U����j�U�������T;#TWUUUp�C�e�U��j��P%C��۩H*�Ͱf�V��l���U������UUU�UR�ʰ嫶���`��j�@��*�yG2��m:*��*�R��R����Pau�$�d����˓Z��UDT����@j�ª/" @�1C���lE?��!(B ��:$$��R� �d� j>�U�H�ҏ�Z�&)��_DB��Щ��
>(��Qv�"��`@Fv�W��rI'�POP~��|.8q�|�D�E|�?*)�M" S�I� �x|������iT'�{E��@!@I$|�=�(訯�����p�)IH��$���!�;U؉���}A��(���/8.�6�|c��z@�Q � ���\D҇���Q4Ч�
qچf� 檞��POE�>���|@}x i��
*�A�.�UH6�A�BX����l�A�	�!���ڈH�AO� ��>("D�C�(=A��� �sڡ�O�ǀ ��0��S H�#�Tb� ���*�
Ad�	�!�P�P� �:�N��Ƈ$b���N�*��C�����F
A��bA��,�� K�F���J�cD�B��IH�b
K
�HJ�@+ ��)F%�%�IIe�`V$�H�Ѭl,�%�	J���� �F4*�Č$�B<M���� ��sB�t���@�c��@$_���y �8��]�����_�=�U��@"m�]H1J#�L
 HĤ(�"B"6)B H��Ro嶂���݄���UV�mUK�5R��F��q���4�7�j�����lRD�����'$6�P�Equ�;5 �e.v��=V�v6�8�2n-k[���dZ�N*�Ő��<�����^+�Z����]��W���`�Ѝ�2�d��Qࢫݴ����ƈ'jnme��x�v����9&�odu����p����uR��X͗�3��E���e֓Ad�Y��ɹ�q9)VٔmUeA2����i�	���r�7t��9ך�J��綛����wa�vܭ�Pc]	ڬj�sc�ȝ�x��-�RWY��A���#D��I�iL��v#"00GW���2)�v7q��M[F[�n��rܥq�d�R��\�U�)e(&�Cld��^XMxWSZL%���f�[Ga�l�4����*;p������&��.p@:	F�
k;W;IZhհ-��(6�M�&@ٕ�-��:�y������A����0 [��V��5ht���\���8ܛF�%��+\�T���4�;3t��5���rq�*�o��1�N�@�nNmkn���g�|��P�	
,65���	@�	&R�D)]hfˉִQ!f�<m���Ns�(���;a���J.-�l��/]̤:]��p�Y�"��2l��4i�E�,TԠ-J�ڧ�ɑ�.�$�ʨ�ҷV����6�KW)=���4�W��8zcѦ��hj��f����dVm��5��cl�S��N�d�ք$:ݚGc[E[g�'oc7A��x�ZR8��8M̠�Z]��Xdֻ�j���	^9l�	�(
������*8������ĉ�g�	�]��ru�����İΕ1K��La�e�!��1�q�J;'8��A ��%�UԖΪ�'mT�b�6nv0�(�G7*�^�鍖�Q�{WmJʱT@*�ki�n���K#T��]�gkZ����G&�6��f�^��	R���.��� ���]*�����D�
��D0AM��>C�_ �4��J5Y8Y�k�+a�����Cm@�vՅ��$],��n�)Q�D�XF�3R�-�S �V��}�p�g^ݨ�u��1�Ɂώ3!���y8ڝchngM>�x@��pT;=�n�q���<��XX�l٪�YH!�d��IMM�7��S.��
 m���ghct��g�B�mخpC��m�k��,�^
�9�vѬ�[u����!�P�w�MH^9&�*�>ۇ�`���9�vÐ^7=�S��Ó�[m��wd���� ����͏ ���Z��@�Cv��	� lڏ 'v<f̬zD��AbQ]�8۶�f�x;#����IOOe`�y�X*H��S[mն� ����2�nǀ6��>ډL�I�մ;co ٳ+ �v^ lڏ 'dx��ʪ�kǽB_&�V$�]]bcf��P�E�n�u�xޥض!��ˋu�j�l�T̮��3����������Ix�2�㠥Ċm�'w��f�߽�k| ��V6|(���z|�������5n��7IL�[�4�[t��^�fV�v^ lڏ ��qXZ��T����Y�H�O^ o�y�{��s��~��'��hT��`�Hh�u�jݗ��Q�K�`�2�W�=e_·V�v;�}usO>���\$����}*�r�����c�\Kq	�C���vwm������Ȱ�2�[��	,$Iv�N����t����fV�v^ lڏ=\�U$vW��6�MRm�cmd���ݛ�{}����<�"�a[D�q�r<��, �t��[i��'v�ݺ�5n���(��Ȱ�2�㠥Ei+@�j���(��Ȱ�2�[�������X�3*Җ6a���kiI��j��:�ʊ&5`S�Ϊ��&��x��F�d٫��w�� ٳ+ ջ/ >أ�$��qX\�]�.�f̬�UUʪH�g� ;	�}/b�>���Ri�-!�v� �ݗ��Ǉ��Ļ�X}=��M"jЩZR�m�[V� >�c�>��]�9��lܟ*�N>�����7$��"K��V�ui����� �l��5we��lx�ʩ�z��t�V�Ĕ�Yt�XWk��h��ʁ=u����q�נ��nU���m��+��ra[��{��>߿e��l~�W>A�_��v���t���N��`�e��lx��X�fV |t��E�n��v���lx��Xz���}=��E'� 4�'t�cV�ج��=\�]����Oef�)�g� �ߞ�������V[��o ��ݝ�?{�| }�缶�.{���m�)NE������C�����{.�틠9�^Y�a�Ы%�4ͱ��x6�`�kB�GF�P�h��4�jƝ#a�������*&�3�7a���9�m��':W&�]��`i�f�h��q�h݀ru`9���r�����A<���� �5�vD�,t���,G r��[`��۬H1�"u��r٣��v�fK$t��엢N�ٰ�ݰȍ�����9&�������LR=���g��-���{���^p�d3��N�瑞�g,�`í���n�~!M��I$�v?�I!n�x�K�'����a1Ho��͈g> ���މ!n�x�K�'���$)��N]�R��}��Y�fv^��{�| ;��vw��߳� {�ߞ��ڔ��]Ulr���rs�m���� ��� ��ߞ� =��� ������.xh;�����/���~{� �ߗ�y��k��ޢ��ԅ���Բ�%����nC�̘��m��0����Em�.H�8�۶�m�鈺��ʽ ~���@loI/�G�W+���^�oI-$=Ʊ�6��/z {����z�cC渔Z���P�B�	�;ޤ�����$��7�$�wc��Uݥ<�
ka��Z�e| ���ϝ �良I$�v?�I!n�x�K�-*�i۶��%���r��O[ĒJl�ހS��g� ��|����6��S�"�6s� {�=�?}�| ���zO}�> �B��`��v��E����j�16Ќl؏(�h�-u���M���+�A�3e`�{�
~��� ����$��-�I%����IvZT��wK*�*�� ��|���߳� {�>t ?}��=���^�6h	�����߳� {�=��,�������\��$�f���$�h)Ee]4�
�.| ���ހS��g� ��~{�
{��� ;{~��a��3q���6[ĒK��|�B�-�I%�v?�H)��}t�]3�R�!����듷i&u��J����0��D�5������Wc9� ;�ߞ��{�| ��� ���� ��`����*헽B�-�I%�v?�I!M��$����{lb��v)��[g> �~�{�
}��� ;�ߞ��{�| ;��ﮤk6/zO��> {��[l�{�kv�*�@~���~�z� ��#VUk�> {�$����z��$�vy��I
l��$���!iu��%��:�ṃ�;��u	�7Tg��+�L��v6��v4E�Bd�ހS�~π��������� ;�ߞ� �}��Y�ҹ�j�eπ	}ݏ�H]��$���e��Iv[Ē��|Y�0j���e�@)���	v����$��-�I%�d|�D��B�>�gRm�� ���n����| ��� ��π~���c
��{�
{��� ;������>�|�ߵ�[o��(�2"D�2,�2�F(�"@��	Üs�gHk�i4�U˚Zi�ѳj��HW7^�,���n�bd�;Nx�+qX��GvYؖ��wW��9n�G#+��(�j�ݡ�։�A�.��j���i!�-̹��۱њ[�u�hوLifC��\ִB���p��ڍG;ũ����u���YB�U�mAD�[.�v�M���M풹W��%ŊqB�r'F�jkP�d$�9�4��;O��9�<8|�n�R���:���8��s�/�t���؞�z1�6��i0�
�+InFݽI$��|�B��$����$��߳���a=����PL��;%�I$�ݏ�H]�oI/�c���� >�YU��� ;�ߞ���oI/����Iv[Ē[�%��M1��� ��π�}��@)�g� ��~{���_����цMr�� ;�ߞ����| ��� ��π~��j7;m5ըd�ݲka�D3;T��,t�d��W2��y�i�-���0nj���ހS�~π�������Us���$����K��4�W^�mk!ff\�kvހ��w\�R��)B��@ʥx� =7�ؽ���$���$��e�I%����Uw{�bP]������� ;�ߞ����> {�ހ{�(˱�~Q�M�s� w��=�?}�| ���zO}�> �O���PL�� �%�I$�ݏ�H[��$�S�?�I"{���0�p٘3Z`����JW"M�dBQ�M	hJYp�`jZ9�Dɜ�\� {��zO}�> ߾��@�}�| ?}�ŧ@nM(�ge�@Bݖ�$�����I.ɌĒJn����'6���_�l�p�&�.| ����[m�﷩�xz�RRG�V�X�R���(@����5]X�l���ēd�����[�V"�[H��
$�*��%c	��M!�r_�h�Xc �}�A�s�fM��-� l�ٰ�2󁆠j�H�G�L�p�iHp�	����ŁP5�&���ؿf�K�0���dލ���D�	�H�4$�ԭ"h��L0�|_a}7|���Y3��3Ĝ$)��4�����LIC�v�8�Ě��R�J�2���BJ�y���r���d	p�P�`���"V�e�B"�).��c�J{���ĩ�+,�@H�m�,c�0�^����b��
1#(D)(roB	u�vMe��l\1�`��)J�I=�xfO w���>��r\��ٸ���,7��n�*r܁�G&bT<T��<9�䤛L5N*u�_�tU�%����!0��eP�P��2��h�����CN����yo�Ä=�|7ﻄ�E14s�W5���J�B'(��)|��'0�6l�, �U0\%B	! �D")IeH��%$!13_y��󇖞3.BF�1�10t
���Z��ֳ(Ĉ��9��Ѕ�����g5� ���޽�z���tCG�x!�CkꈟESπ�E�� �RAT!�O=J��`T~D��|W�LQ4�@������-�^�����O}�`�2�s���m���o��<��$�ݖ�%��w}����$����U��ٹ�ڂ�� ��~{�
{���K�#��]��"(��4�ۧ�6�%.�u��u��UC��O^��N����ΰuލ91e6q���u��Ͽz���I�+��9�I�Ih^��Z�,mU��x;#�$ٕ�v< ����H�ؐ{��2�[v˷m���X7c�ԑ��� {}�}�Б���V5n۷n�=�K�y��<�vG�S�C����b��*B*��+_*@�'�r�U�~�+ ���,Bjں.�m����ʪ��s�O��_@�?~����m��=��.qK�f[ḗB���'��;����>�z���@2;`�+�������VW[�Mһv���@==��	�2�n���W�I�$�"ݎ�.�v2ݷ�Nɕ����y����	�Uq#T^.�a�M�mUؓu���v< ���	�2�	6aV���whM��x7c�	ݏ ��+�^��}6�˽[Ͷ_ ;����~�'?s������ߞ M���*�q(!�����uAe5��%CֱR���!WL�8�Rx�f�U����g�v��E�1�Ms�L��Ɓ;���={b34v,�?玌.�J$]*���C`CP#p���2v�0�b{d�����GnN�t
W��Rq�f+�\�A���uL�8�'X��=h�5r�s�î�}I[�rV��P�����;�#-��Jٮ�A''}$9$�M�F8+�4�L���lmv��X�q����k�
JG�	��X>W�#2��W���� ���ݏ� =���;@���V�m�u�v<�) ��x�x�Y��9č���&��Be�j��l��	ݏ�W��*�w�{�V ~���	�BXe�+�
؋m�r�ʪK�<�l�V N�x�+�{g� t��M;�I�e�n��&���?U~�/߽������͏ ��
ue�Pv2ө\Pug9:z̈V�V������#ȟܓ�>jY�2e&�Y�m��y�� 6l~�����V�OaW`\��l9\� w��|��s�|��I ��8����k�s[�{��ٹ$�߽|�99��Nl{������bٵ���{��;ݙX]{���=�� 7}�N�*�Q�5N��e۶�=�s�[��V {g� }�������� W�16�iݦ� 'v<ܪ�w� {g�����?W9�UmzP{�B�GAl��[!Vݡ,f�U��C��P�iV��,0F���9$�V��*d�v.j��?~x;���{�U�|���<�*�����$���I� {g�~��q#�� ��<.��*��<����I؝�v��=���	ݏUs�ʃ��F xB(`��8e@�,ZD�~���_;��{�xiD�+�U)X����l��r�/I�yl����U�^ٞ0z{
�@�ջE����x]�x�������l~0nǀ~�*{�Y~pQ�]qƓ"��&��a5Aו���u��f��θ���}�xM�eS���j��������v?s�_ ����=�
��σ)շl�v�;����ʪ����~x�=�����ܮUs��h=u�ҷut�v��$��"���ܪ�q.�{׀{c�wv X�����m�x�W�g� ���x�`vr�,b�@�� �$B8)�4"�A���(��dD�A��KaP)�r�=UU]}Ϻ���2��N�����-�x���3���� ��/ ��	{�{<���5Z$���,��>�kz�lY���ن��%�ŭͳR���~�QO�a�b݈��~�� �v<.�W�:���J�����שP��6�f }�W9���?)�׀j��^;������Wm�ұ�.��<�z���?W9����������<KF�]ݪW*Ҷ�۷x�R]�� ��� >ݏ�r�U���7����pY}�����e����~��Uʽ��>��O~� �v<�{ϊ$7��1[r��;v)�Q���f{m��J���Ylt���T\�t�h�ݧ��^<s���>ۓ�t�ݻL��`�s;h�L�Aͤ�ƥH��R��i��v,�v�e�n���Mu9���z��D���L��x�&݁�SIA`S`�W�i��š����G1��8����9��������i��u�WX�)r�2��)��l�>�y-|`Y�д]i`�	�#6!��c��6��V�&�l�]`_}�{&�|SۊЍ���ߞ��/ >���s��~0��K.ݺbav�o �ݗ���?s�v�ߞ���������$v�!z����v+�w����>�ᇹU\H�<��y��t�C�E��n�+m�O��� ׽��~�䓞���'T|���䞔�ޙ���.L�C1[f ov<�ʪ�R履����7�^���۵�n�Ŧ��M��@݇�Z�q`�ȋ���-�0[Úc��'$�E�ـWm�IYm�� w�� >������'o��nI��ffR�\���f��$��~���
mZ�
V�aI�)$@����B��dR�DJB�$+����ɭ�^��;{�srIϽ���$��pY{����f\�߽|`vK���$w�� ='� }�DW-S��RM�+k�UK������lx�Wu�� �RK-�B-&�-7x��x���'��wo�X]�ym��/�m�,ZP(*��
Jh�Ҭ����V�b�FqH�8�9e�%����R�!|n�E�m����{����� ��_�s��vy���撶�ZvSv�[��܋?~�U]��{��	=��vK�UU$j��eߝ$�L�'m`�����=�[��?,b�$"�� UB�A`"�@�8���X��*	@
#,Lr)1�x�����~����y`5��!]�]%e�����*�In�< �xݹ��T�d��;�D��v�יM6�m�۱���s����d���c�&ܫ�V�7`$������N�7e��@����6˰��n�H{''9��,�k8�Uf\� �߼�������UU\��<���=w�T�at7hV� }�~�+����I�����'���nI�3��
��ݕ�BX�J�e��x�<����?
��\�~�߮�����$燶��1�V�TZm��\�Uq.��M��rI�}�[���G�a
�J��Ȥ^1(h�+�F��Ӕ�]4ы��>R����石rI����nVk\#��_ ������9'�rr�W����5~����c�	�(]��1�-1LĎԚjKL�P!�:��k�Y[y��pV�rrNO	|������c-�d��>Se�۱���W9�	���;�_Me��T%�.�|����=��r���F���Oy�0{���r���H����ګ^e4ۡ6� w�� ;���9\���� �y`�
��Q8��M]f��?'�L�]��ܒw�����>��O�/�Us=���ܓ�����ZV�I�j�� ov<�s��\�9U��ߗ@7��<�v^��U�G��W���4.�z8��Ek�D�B��R&}��=��J��H�yCI��=޶3�+|�f�|���F$�k�����<}��f��4��&Y��<#@�|+� ۶����U�o�zO<'8�J�Z�f\�]{��#"�''!Qr����D �H-�|,9/�|[h*���aK�
�����^y����<��l�uC�:3���E�j�Vv2UV�A�*������kv�K��9�p�>���>�DN�]jn�@n��
�.�$a)�/l�&�]�ώ�'��*h�5�o��@˚41��lY��L�*���Hi�H��n�ڇ�U��.�mˊ�Βx�8U��ց�-�1�j����"�WJ�L�Jz8œ{.<20g*EU���u�8����:���d86ó�͞�{X7I5��G Z6tpΝn����킳��k^R���
�!�sY���2�e���I����A��Ҿn݉����*=( �㭮���7Ӳ:y
�]�mʯsb�a�����\��ݷ8��3�W��s	[��җN��vAE���N�9�ov|�8�	�
��O7�y��	
��f��Q�c���u2�s�g�<����Z��-���+g�6�\�t�y�������C��з�1κ p�l�Q�&��OF6\u��E��e\�M�i箶����F�y9곗���ڕ�-���t���%�Wk\&۴m���SH㜽�\�ob�h��x���1<����=v�X ���z:˙���Q�ѫ��o=F�e3�3�v�t�ʹ]�(�Vz�`2�����������
���qnn��ƶ���t맨�.�ܬ��jqc[��];����&�,�e�8�RnKVh;/�l���m�.��eS"t�Z��/<Ǝƚ�Z��]��yrk�]��vU2�H9��e��	/k�yf	/8����T����S1�ye�@j�k�-���ә�0���s)�xΑ�"�h��5�BùGn� �;��a݀�t���k4H�� �ٶ��qH�^�:�}���cNI�Q[���
8.�]s�Qu����8�G^�|�g3�	N��vDz05�VV;#m��h� "�Ll;����'vҭ�ҡ��L�JI���	��	9�<gs���}�Rb�J�粯lAAp�2�*33M99�$~44���) �C�`����=��*�̀|�}'9>�9'���o� �j��]uH����ð�N8��8�sU���H6�Wמ�lK75��\<�,�F2��q�>,؍�g��Nض�Z\�ɚOOe��M+ee�#��i�CF���ːSA;�L�a׷�4u�ۭ���oK�q֍i.�F�C���ϵ��@S�k8�*���9��[��x�n;[��;r�$��Յ5���Qf��[.33�d�ȋw9��e�xfJ\��j�Y�vl����h��ˎ��'�;,)T��%����rLy<��`��Zn��'�~X�����~�r�_ &�<�QR\�e65i�,M� �ly�U�ܪ�.Ƚ�׀�����o���%��}��\��ڣ��_ �����c���r�.��� w�� �Q�^�n�鳗x�I�o~���?��� >���ʥ�'� ��Ť$��0�jۻ����X��W8��������c�	���c��v�|M�J��Z�w�����Ov�P��Iqt� R��d��9�HO]+�V��ۺ�� 吏ջ/ 7��s�UUWl7����?K%�J��F[Q�_ ��~�xI$睖I$ s��2"ы"�Z)F�#l��H@������
��QrN��5�'�ϻw |�޾{�%�{4���fV�[�� �<���Xz��;��j�׀w�R���X*WC�M��=������un���RS}�{j*K���M�����͏ �6���=<���X������R9�i��ڼ4�n�\iv��L���о�j��27�.kQ�O4|<�^l;7N�^�� ٱ�ۑz�����:���j����wWn�� l��ܤ���, ��xۑg�T�=�Wv�V���x��� 6lxv��F���W{��O��u�'��g�2թ˻�l���~�����~x�~��{#���W9W�敏�b����E]:I�;o ��L	��R���l~0�z�g{��`j����u��!��scDWo.C�
%f ���8Pc��.vВn��k�	���'u� ;6?U|��s�?RD��!	^U�V���m����I�y�۞X��竉�\�e:l��jـ��N�Ň�&�� ��� ��*��[t�Ҷ��r�����{��Oߞ;����$v���A�E_<���=륧�e�t;-݅�k 7�<�\��?~����	�ߞ;{!D�-׷f���uz&xI'��֍������Ã7H�4Ӊ�y�bl�a��/m���� ;6<�\=_ &�� ���v�ם���l�͏=č�~0o���p�q#��Iz�E�BM4�}� ����))�~0}<���(�;nݴ$��m��Jo��m�� ;6<W����!,e��I:��o ��� ���U˟���������7$�b$������_rg�Ԙ�Y�9��V���:k0kb�H*���V�,SR���ʡmU�n�L`k\$�fkM dk.e6ƈ�c�8���c���G/A��� [�dҞ�#��H��q����ps!�a������vg����v�电:��Ps���N��62�	=�s�"Y|���UIn,�q���7&K���Kj�gX���2�6!)tLvI�I�q���is�m�ᦨhM�0qGpYp��iK�O#�b(���f�r08��'6[�y��	j����?>����){��}a���a䆋V���n���	�p��ĉ���s� 6ly���H��^<���:�[���`��X��X{��'�����\���V�0��.�����/k�X=<�	�p�u^�*�W�� ��B�\�e�!�[���'�{��$�(~QCg��t���^����>��ZX˧`��E�ư#)@�4�L\�XLǈ�j ĥ��-G��������!�P� ���ov?����{��ʮU|���xe�QU��m4	[j�f�l�9�UQ "� N�������݀o��}�p���?W*��r��=��cW`���w�l�~X�c���r���v?^���Z�EJ�un�t�;m`z��Uq)��wc�6<׹ʜ�}�}� t���� ]�L��|�� l���{ l���%>��eH�큀խ"Й�֎��m�G�$�.���y�rrJ0��]���E�� OO<�ݗ�6?W+��v?�~�QI+Vՠ�Z�o �we���s�UU]��{��6y�0fǞ�9č�V�B�Uk�*�I[� ��x��
,�2 H�`.�F5`# �#*Z H��U{���	���5o�x�*T�+.�v�7v��\�ݙ� '���ݗ�ꪤ���ݺIK�&۶�+m[l����+�U�ܞ��'���������;���P����e����8bf%B�K3t�������N=q�@^�k��aZ�M[�'� ;6<��ܮW�	���6TT#Ք鶓�N�Xٱ竜�Gv?=�<��ş��W9_��6=�����@�bU�e����x�#���U%ݹ��y��Jm:ubi�Iۼr������;/�X�#��r���s�r�y`���E]����e�x�r, ���ذvG�~��l�Yw敺hK�*`;���5SD���r����[aR�2�r�6�'<��Z�W��|
w�	���wob�	���ϐuOz���J�=i"�j�M��wob�W+��I<���^ };���s��?NI6>��Ot?+��nvsk ��~�x�d�=�s�����<�� ui�*N�V�ۼr��]��^ O{� �܋ ղ^����^S����;m`d� �+�[��)�^ݎr�Zr��	�WqS�ʻffGf�o2\B#��K�F1oN�%ۛA���h�ݭ���	�wn-��ds-�(�D+eI�(�:��8�wO�v�<�X�F�v�]\X�t
�wi�'��\v�:���{�> �R��ۇJ0�5%���2�ɫl\���k8��du�Xԅ�u�+�r�e7GT��{6ݒ�4���؀�48[���F2��Y�x��e�ڬ�9'=)�+���K���C��0�)�
�.������X�z幦�.�)NL�xߗ��/6Yt7An�17J��~��vG�wc��ϐ�y�ۥ�ȶӧLv��v���{�<�Us�������,�+�����v��4�bm�<�`͏�Il�y`���7�Z�+�Uq�t�M6�=�%=<���, ٱ�?s�������x�ز��~��F�a���7nE�{��=<�W��������<���l������2�U&��9�2�a�`Z���S�c�(PZ�+n��_ OO<�Ix�c�\����,�=FJ۱R`��ݷ�uI�oZC�a��"`�22H+�P� �`##"B��1Y�������"$b��	��F A��bQ� ĉ A"$c��ab$Ȑ ����b~����~x��~X�c�s��$OW���:Ln�RT6�?RA������,=\�~�*���~��E����7E.�`[�LMһo ݹ l���%�z���S�� �����m���]��fǀ{�UͿ{�����7nE�E!B��=@M��rqeT��%˺b��{�SGn��X�A��m���Nq<�m�m�«M��j����ݹ�U~��T�������zM@�ٿ5c�9� I��ۑ`M��wnE����*�W+����,��?kj���_ ￟ǀv��ٹ�d(aԍ���d"=$�$bpC�3���3��Q�dɘ�a!	 �¦y��Y6F$	���t�HA�p�-X�4�O� S�"��$����Yq}!�s��<�"&�v�6��l�U��z��(hTpÃ ���&�I6B�@ �iD�M�CF��H�����1>H@��A! dD �$A��Pk̉J�b�oF�BX0�WD�+��!	�D�IW���c	Kd���%�Z��B0`�WQl$$0�EZHmy����A!	�B'ރ��lƆC*_���� �	��qh�p��%�����zf>�@p��f)�u�t���0C�>�3�l�Y(��_CL�� ��B���Br�!W$�a���M(�T�_E�`!�"�!�����=���A�h���UU��s�\�^����	'���H۴�!����jف�W��׀j��x&ǀn���FշMP��m[xT��s��9��y��	6<�O]��U�h�*x�J<��9�̮�H�MY��9�iiU�^Yb�	rr�By<��+B�m�@�=����	<�`���9���_�~� ��	~�C���j��7nE�j�/ �^ l���T��GW���j���t����=xeȰ�_����~x��,d�b�Wv�S�U��Է��=<�ۑ`w*��*�!#D�0#$`1�A"+��﷛�s�g�C2�>�f��;�`͏ �V��/���׀wc���~׳Y��U���*p8f'5v ��X�)rg�Q[I�`x�����`��.
��4����j�/ ��r�@OO<��DV����I[v���5M��wc� I��ۑg����OR��mӱ���M���� I���JK�X��TҊ��lN�Ъ�f��/zy�\��$��0M�`]:����]�x��X����x���� I���¹ʢ���Uݸ�{?�}��S��A
�(]+:\cT����n^ԗ3Գ�z`�`�cw%�t�sm�{�a��橺��y]�]�ԩ~7����o\DktKԝ\C��;�tL���F�O+[�pM���n�5��mӴ\�j�����&y9�A��c�Q�Q�i�FY7$��^�uIsn���uc����^U�m㙛Vh\��W!/�y��*�']f�m�.c.�zR����Hw�����:-a��\]��.�3v<;�� �bc(P���MT����yb��\�&7Iݵ�7����>�� 6lx��X�2�@��N�ؐ�f��c�7ob�6l��H�*���e�]���0d� ݽ��s��Kޞ��;�?��hI�.��M��n�ŀI�+ �c� I��it�+�)+nݶ�	6e`lp�	6<�{�]Z�(����e�a�����c��l��0晵 ô���,&B�ee���c��)�u�}�� 6H���X�2��JU�SmXդ�ݳ$�߽�[ٵU�
�� B"�")���M��,=9�]άwfV��*�j��Л��t��wob�6k��.��� OO<n�WR�i�n�	^�s����, ��\� ������N�:I%l�>ۑ`͏ ��ŀl�� 7��-6��jݻE>;��1��]
��`Ď�mìndш �VJs���7trZ�g� {�� ݽ� ��/W9ϐu{޼z�)�`��h��;o ݽ� �8`)%��<�NKO聯��룘Kr�-�}������f�غ�>0н|�w]��7ny`ݔ���j��
n��5M��H���`z����I�^(��1�.�&���	$x����z��l�I'>���.Ֆ�H���$֦|v�xe�%��跦_X�g�:�i�-G6���[C�J���,KذSe����m�VRci�e;wl�$�� �6^ I��5� ٳ*�)%t�t�V��5M��~^���o��K�`ҮXwVB��e;�w�H��p�$��W9�]����*%��;I��m�v8`^ŀ� I����wt��s 6K/�1s�-ʼ��2�M]B0-vq ���051n[[�*����`���	$~��s��	�~0��YWI�NƒvSm��l��W8�{���'��I&Vz�"OR�E��1�.�&���{�x�p�$�+ �6^�?���WY�1�e�=���;�|�{��V�l�UU%�{� ݺ��r퉦һ�i�0	$��=�W���$�{�nI�s߮�_�E�t���*�X�)�R���M�չ�Vj���	�<��㨬��;V�ۋ�����nN@N�7bqқc�p�JD%MpB�f�kIl���ݮt']��ɺ��6�"ӝ�P�H�u���7iy��ѡ�Q�949�+����6k�Sh�G����r�S�7f��)���x�xe�ҫֺe7��pM����xg�q����;�9�]�fkYm�nN���SElİ��3��5�&h�dTX� �̞ża��LE��ˋ��0��m�N���M����=��y��^���m��7�Bj�	��lx�{&̬aW�Qj��;�I;o $����,M�_��d��'�Tz�hI:@�M��}��`l���c��+��^���;G�+h������X�2����M�ܪ�.�<���b.��i;�M[��/ 7���ŀ|�{�����:���JmX�M����5A7Na�ߥ�{8�����=&�rD\�<��H�ݤX���O<� �G��9��=x�l����T:����7��e�*�o*����s���]�X]��wc�;ۥ"\����6Si[X��X�l�=U�W*�&�<m�,wfZAIU���I]��|����ǀoob��.��,�.YEݖy�V�(N���ǀooj,�r,�6^��?���#T5��%���%�4i�$R��(ꦻ a,kF��i
h|��v�����>�� �/ 7v<����M�EۧwwM`H�|���ݏ ���`�+)]5Luvեt� �/ 7v<=��+��s��r����������+1��E�;w��U%$��	���>�� �/ ���%��e�huui��݃�>�� �/ 7v< ���K뉒��+�s�+13[���f�0`F�@)�æ�B�It٧6��.x�f�Z}#��6^ l���`�	$��Ī�!В�k �/ 6H�{�xˑg�T���(���1]�e
�� {�����x{�Ľ�������;�)Q-1R����m��j<}�}w$��߳rD��tD���k����<��{��������`9����ۑ`�9���/���z�{��v�3�tl�\� ��GP��.l
^�G6x��2�gKә:�\�^�k ��� �^ N�G�n܋ �j_�!�[bV1ۼ�Ix;��r,.��r�IU�^���U�[J��[� ����7nE�Eݗ�uI/ �n��%]�t;�[�n��;�"�"���:�K�:��x�eZ��*�v�v^ղ^�6���{�}w$�t�"�li���͚tj���4!���d�1�<�X�n� FqjB���%�t%|�8�xA!��c sA����J$H�6����tDHS�F��o\@�.���8���e�34B1����Ӌ/�D�HxCG$c$�a!3L���2�hf��.V4�I#�i1}�R֨�`s���M#�~��Z������Vꪪ�E�T��UR����ӊz�hKh�l+p�E�e���ۧ��:��UP�ॕ
F[��u�ތ*�r$s��t�>4X�Z�!���]zFE���yݭ �
z�<������!MT��M^3(�n6B *�t�i��`�!��3���3�$��q)I]`<ؠƕ�f��#L	��Y�lE<�8ӻj��zLj{�i����\���<��ӈ��m��֯q�;)���mlG:�����Q�ܣ���YXb��g��N�mR��iD�*([děf�4�eG@8J��� k���a�շJ�W�ܩ	�-��I�d����T�C�,��8<<g���]��pd�0�0Ytֳi�9�i�9WhR˸�ň[��&lWzc�Ǵ���'�CA�8�nMt��y7m�s�ts��}�jn��m�ay�y�gg����Qt �]��@+$�P٧��P&%h۶#���ԭ�4�gs��\v�����)[�]RѼm`�CmcѶ���(�0;��u�ܦ2����&f=jZ8�v��#��q��5�%�A�o�&룎�(خwL��)�
c����x�e�V���H.M��sJ���YqnI�q�
���v�p) $�Nw�ǌj�����&읋n�W�����5�(�+å�vz]�Ɔx���S�(��oY��iz֠�m] @��-*�IK����,�-�m��0j�7<@x�*��RX�֌��UUe�V���r��qKҤn�:���e�k[<�-UtPg2�<��d�lp�KmR [�q{�+u7�lQ`q���gm�j�nw���QGM0<�C.�Xv7bnڃM�I�6w/��ݺ��S�`f�0dx4ր!�Jؚ��by�8鷖ĕDm譣:���ٖ0#�I�Ίk�&'+lU�8�;>&��9��m�� 8�馺tF���c��b�R�*�UT�ڠ)g�`:U����l�ȷc�aj�v���w*���յ��]fa�Ѣ� �4��}@ڈ���#��*6D�������/���� |,PC@���<�=u���՘C3WSeJ��,n��4!RZk��v1J�ns�4�@�Ф�Zɵmj,�����z%�LFe�kXd��p�
L62�vK��vغ3�I�`��\Y��h�Pؖڶ�c�N�{s�#۬����;0�e�8�u��l"3ݺ� I��f1�NN*z�y�t!�ؤ,��2f�el�I�i:;
2	زu���nh׎W����Ae�T�w�s�/'Nv�|�m�jܺ������Ѓ�Lfa�хLKԩ�I�y��gGnu�s����uvڦ�ۀ|�e�]�ݎ��s�l����*<[J��-���:�.<�0[�������8��]%��7��)�`+��	<�`�e��<Tۏ ��+,�SiӦ컦�X[��I�mǀIr,M�|J�)�[���� �G�j�q�\� ��/ �"?z�:���ۭ����Q�`��y⁫Z�Rzuv)#�ݎR�CF��f�iv_�}��z��� ��/�r�ϐ���������tL�r�{ק������FrE�r�%�ŀlx�eǀM�U�
�:I*I+f��, �G�|�\|����;�}�.&݋����$� �l��	#���,����
�h�i���>[.<H�l�� $��بt�e�U�7V�b�<���u�x�s�卆уyk�ʹC����:-�j�v�v�$p�6^ŀ$~��9��T����z��iSj�Ҷ[f��,�UW+��{���:��� �8`mK�WYN鶒�4��	$x�T��+�U�EUVe��j�/ �]���j�i;�o ��#�$�eȰ=\�K����R�V�ݺj�V۷m�#� l���ղ��5HR��4�v�-S�WN׋���s��r���Iһ;iU��h��m�u���mКIRI[0d� 6H����8`�`����6ۢ����<�*�čS��Oy���<����
��[�i���.<H�H�I%�P�i����x����0��� I#���������}��~_^;����)�v�i];l�	$x$� ���$�����yW��h���snv\��먺��x�B�'�	�۬l[[R��m��I�F:9)���{���:���I2�l� �P6��eڦ�v���=\�G}�ea�G���d��"��K�V[�M[*�m6��L� �#��ǀuIq��I�
�wn�=I{����� ���>�2���]
�+��7mһ������9U����������Ԫ��U]"�+�����T��N��5�yr�7�7m��9��ޖK[���"��s�\\	��{����ǚ{Q��*v�����������6����m8r��f�uz���.�a��w%��9��v#���	�N�qP��d�M�v5��&�s<�JZWa!r[tVU�� f�TCM.ɥ� ����gq5r�1��������nǫ�R�+�s�g91��5�¢��	�t�HB-ɚ�,tƜ�����3)�Q�`x�X�!�I��r���~=����d��� wv<K��*ݦ�*�-[x�&V vH����Z�y���6~�X�eӵwn�+n�~���wc�s�j�[�&V��T��+-�Wl=\Kwc�5E�<�&V vH���E�J˵M��m�����=����� �x���BK����EÌ����T��8��u�9�ŉhZ}���9�lQ)3iv�KT����;޽< ��x$��>A�=�H�_�B蔒��ܒy�kx"�.�Nf�<-�W�l��s���RA �^t��N��wBv� O{� �l�xPl����즨Ur�ĭ;�v���r��T�g�O ���ݏ 6H�	-mĭ�t0��L�m��6G=Uĉ'� O{� >�S�=�{ϒ�9�g�l�^�=OC��\�F#a���sL��ÃF�HXL4�Q`�tn�F�9O�$�x�G�I)�G�*_ٔ�ۻWe'm��<�UU$��O ���`�ǀ����J�էIZ���%<H�z����\�U�Ԍ���;����'{�u�'���R�]��J�hv��G ��x$� >�)���\t2ШI[0���� }�S�6G ���V,nj1�h�t�2LK�a�<s�� 5�=�.S�1�6omaz�5t��v�� �#��Jx��jݗ�}�l6������| ���>{�I�?Rz�d� �Y�N�WN�|��x��jݗ�$x���ޒU�1�N�.�m���y$����ܒs߾5�0P��QB(�Vq�C �eK�2��N�P˷x�G�z��vJ��	�?�v^%Ϯ27��G���p�˲��N�=�v�;�usm�=�wWuƵ�@Ό�Xn&[x۴�l��v^ l����Q��v�ݻ�I];�6G�/ 6H���K�7u���$�$���/ 6H���K�6I���*�*��H�n��v��O{� ���� ݓ+���9z�z�	�����Z.�]�un�x˵%��e`]߳rI��}�� �!
"� � 2*��"���߳�Ku�̎f1.&3��D�\$�/h�;���lsHg���F܍ӛ���8iE�n���^.�"˒[�Lb���sM
jjzc�xqӜS�{�l��:�5��M;�Z>\Z��n�:���r��b�'�#m��;vy�·C��� %N�㧂�A�������TV��̀���Å�g��p�� lGʚ4Yl�٬�պ֭�T6
!
kvna��IH��Nݡ:�1��4��P��`0-��!��Z䱰��3:g�l�������]�x6G�|�Լ�6U��M;I���;u�j���	�<�6��d��6TT�f�7b�˷x6G�|�ԼI2�]�x_u(\V�N��i���R��e`�c��<Uwj+H���'mS��;�6I��ݏ 6H��ڗ�l4Pŕg �5�]Y�=������eq
��)�hfg-�s)X�5�5��ņ�g�ݏ 6H��ڗ�l�+ >�*�)��q���_ >��|��$/d�$dd���k�(!���W׀w�e`�c�7e5E�,.���7V�|�ԼvL� ��x�#�$�H�7N�*�6�ӼvL� ��x�#�>Sj^ޒU��M;I���;u�ݏ �+������J���e`��U)9�󦕻G�iS��a��(�FM�_�z8��blJ�,.�&{�-���YB�1h���e� ��ߟ �{�v��2�{��*5).�wc��x�IW�I&V n��@{���"���i��&ڧI۫�$�+ ������DOsCBR����$�K���&�;4Mm��IJ[
JIK`�6D�F�c�ݷ0�Xdpd�ce$h@��,-%% �RH�XFJ�&9Dr��"G�e��-2��F��1�Hq!
@!
�!iP�H�B1�0HĔ�hJ$���i�܉v��
A!GE���pߊ��7��7n�	�]l"VQ��[�a)�����	����#%���̄2�HJ�J��P��32P�cRQR��)
K!.\*��Dn�hV�	)KJW�V$`JBp���LH �)8�	r\R�*��Q<GC�k�MU7v����o0���&`�&���b�u���������Ռ	e �����qV$�@P��v ����� iA�W��� �|EQX�L�<�l��>�Z)%wj�����`%�y������W�l�+ 7T����[��V�i��d� �;sޫ�	�{+ ;�<��U㡶*N�9��Pp;K�+�[�'kt��v	��ĥ�,��1k�K�ћE��������$��� 6H�	,�N��l�V�ڶ���eg�H6{� $�xV�W�n�Qx�n�M�]�v� ;� M����W�}$��;5R9���R�� �����W�Nɕ�<EC�� llP,AB�Q�P��$e�%x^r|��|���߽���������d��'d���ǀv< �)�㑍�n-�e�ke�̻=G^u��κ���u�>�!�WM��.nX*Ff��vL� ��x7c�>[%^�u���wj��YVZn����ݏ �l�x�Y�r��	��*�����v��� �wb�vL� ��~���}��ޘ6�����?��}��'d��ݏ��R^�� �����mP��M%m^;&V�qI<� ���䜾}���< �|�
�抸[	��R��P*�.0���du�Ч���%t�D��0�p �M-�sRj�5�mcY��`�������#u�s��X̜�뱡����r��vM�J�Y�j�a@H�l�)H ؚ斩�v4[�Y]�*�g�N����3�
�n��a]5�P��&�t�r*������y,j5;q{!ዧ��KP�70�O��<5��:�CR��ԙ��55i,�Vd 9�͓/48��7e�P�wm����@`�NM�*�Y�ban�G���Ѧi�j\�1�7)���z�nǀ|�"�s���|���e`��̦�N˥I�x7c�>]�^;&V n�xʃ�b��v�]�V�x˲+�'d����RII<� ��xUݨ�;�]���v��y{}� $�x7c�>]�^�u���Wv���*�M� wv< ���.�W�O����oߥ�۵�b[* ˙��`r�t��%rλnכe�4�c���Ύ�����ӫWwi�m� ���.�W�Nɕ�9'�����>��l.��6m�ɝ�nI��L����`���  ,�* ��@ F!	 ��2��#"@�"Ȑb*��PL2�J�+�' 8rWk��W;��ܬ �� M�����%�V����^;&V wv< ���-�^�IX�Ze��M]�v���s��q-�� ='��݅��e`���2�M:����x7c�>[��vL� ��xQ�U�۞ιG���kl�x�e��(���),Sb;�腙�9H@سf�6e�_�uI��	�2����ݏ �]�'N�m:%l�vL� ��x7c�>[����E%V��e�U��� ��x7c�9̮UT��s��ʮU7�&�wve`�R%˥t����v�v<�6�}$���ǀwe5IGut�t��[�o �n������	'� n�xd�N$]���T��>��'/VC��vwu���g�:m��
���d�4�vHU�Sd��wve`�ǀ|�ax�%b��e������`ݙX���-�^��+ ��H%Y��i������݅��e`wc�>Tv]��ڶ��ҵm�mWn��vI��{��ܟ����3
�A� �����5Wv�ćv˶�:���2����� �n��s��m��_���������N��'E`8�o���4�L$T�5xǞD�iۑ3�|!]��'� n����/ �&V n�"Ut��]��N��o &����^6L� ���j��vOYB��Պ�������t�;����G�H]-��VS�i��x�2�-���Oy�-�^�T�V�ce����`wc�	�<��&ɕ�|��������H�������8��]��٤kA�ƶ��:ܭ��{�/
�q��:��N���������+�������0�W��R`��,ҋ����YP���X���e��5{.�����$8�����c6b-q�1�"��T�`�)�˩q��M�����GB0Z�؆�V��e�CKq���J�E�R1�-t5�/k)5���99'���e�<��b+x�wl�qZ�6{u�-t�$IDƬ�IIX��4!k2��]�N�{�� �n���`wc�:��v*����Jշ�|�axw\0����#�$E[(� T�ݶ�:e�#�ݏ >��݅��®�|��	�6�W*��RRO< �����;���H�]+�I]�:�m� �dx�l/ ���v^�W���-[�eP���^1� ��p]�N�3ٹ�^s<\�킷�G'.�њ�5}��s�Ϝ��p�5n���c�$.�ؔi\ԙ�Z�kZ3rN{�<v����^ w��U�d�&��e��+f�v^ }������U����;J�Ɲ]Їn�=\�]�� ��^��NU]��T�hVZv��+M��U�n�`wc��c�=ʪ�{ȱ}MX�Ɓ�-�V����K������ۏ31����W�7kR���3r�l���������۱�-�� ��
���WR�\�0���۱�-�^�� wR�UuwM%`��M��nǹ'/��3s԰~H�$,x�<�0�*. `���� ���������|��ce��ѕ\ge��l/ �u� 7v< �v<at���mQv�v��>�p�=�$���y�)��v��,)]�M-��!��x�k��[J�ܞTಓ(�YZ�kR�c�Qڷn���e�[0wc�� �M����l�H%Y�cN��eۼ ����ʪHݵ�^����ݗ����}ﺗ�&̦��~��w�vk������ �]�% L���`�J����|���{#��`�A���?������3rO;�H�]�&��6��ݗ�����xf�`v�A�m5m�.������;�Σ������N�:�j�����86��XEE��J��I�M�������p�W*�A%�,o��J�Z.�ӻiZm��v��W���`�"�� ��R��v��.�bj��p�7nE��T�7�x����M	Ye��݂l�+fqv���	��v+��*��g�}#Ȳ��T1ۼ ���[�^ٮT�x*�N���|��d Up	�`B+"D!<����LD��c�jp�����u��Qݵ� F�3,
�X�	�a��Kv���&���'"�хU���H�_8s�|g8as��oc����"O�.k�!���B���������Z�����Q]�)���\aˉ01!(����0O7�%��*ou�YC��'��	���jƺ)�l��R���A�H4��LM}Y`�"k\&���4�"j�C���P�]�7..�7|���aIv@�������9P2����-ζ���MR�v��m��]�\7,�F�#�S��0�FG�mz�jUU��&���a���K��`�\6�gXѮ���Kc`ȍYn{F��eV�4�]����lT�Y
����5"�ؗA�uь[k&�R�+[�Y됸<�J;v�"<���t�nJ�W�-�]v���7��(9w7�h���[[��<�*f�emV�L`��ho]O,=<�
u������������Mɮ"�A�m�T�M'l�īNw�9���K��y�a����ܼ<p�Yn� �وB�"T�Ӟ9{9�أ�[[��sf�c�}�vg �%�g#.�)Q� �+mn2�عV��j�xgh�;�kc���u;r�ԥ�7#����d;=��	��â�&��2�緬�s�����\�+��k�������`�0�T�Q��pi7aΞ��#�����́.�v��V��ANm�*�b6�۔mi����Obnm׮�4�y��g�����j'�(1e�E���c0����nә��`ڼ\�������s(w�vN����B�Ǔ�<�HܗRb��&����X>�9]��v���ՍI���r��v73�͌�^��0�iC�n���;n��b��R˶��s��n*���6�
�&��[�m��cV�5�6a�<Jv���=�U�����焖� w:�l���{pl�z酩�jӡP�MϢ�0e��d�Zc��]��U��\��l9���M��SS�X��8�!�p<��; 9��a�V����ڸ���DW�c��We��p�)��pa9�m;F���K�&Z�h!:�.�*��e����Y\F)ţ�2ڗ�L�n��Cu#�OV�zt%� s�;Q����p��vvٽ��zs��)]e��Ѳ��9Ut+P+��+A�1�-U�@+7�8`*U� J�M��
�f���LUTgv��qJ�x���e�@W��Yne5���5���EЈx"Ю�������?#�OUT� ��`��z���ҡ����%��֥֭3X]R�Jɻl�N��t\�m�dx��,s5˒D�����	4�ڑ���:��薎�;p�ͬ �t���9�3���[Eq��9rV.��������s�bZ��q9��t��ժ�s�a8�ӻ�gmt��I�9S���A$('d�%Ʌ��R;-�\v�`w'v8�ư�\L�˗qX�n8u���xx{f�-�ڭ�$�'&����6`cLױ<�y�A:q��s�-����6%�!.�-F�`:[���̦������ ���l� ����n�)�lV��t]�xf�`Se��G�j݊�	�×e�U�MUm�Wd�ŉ~���ӑ, $2&D�;��6��bX�'߻��iȖ%�b_~��va��rd�h�3Y��Kı/���m9ı,Os߻3iȖ%�by߷ٴ�Kı/����r%�bX�{�t�C�6�vC_9;y�^B�{����"X�%��U����ٴ�%�bX��~�ӑ,KĿ{�u��Kĳ������I~�X��-b��m�("���ry�gB�ضҲHPk!,�������&kFq<�bX�'����iȖ%�b_}�u��Kı/���l?<��,K����6��bX�'ߎ�8a���I�w��JrS�����}|�� �����r&�X�=���r%�bX�g�tͧ"X�%��w��ӑ,K���R�ٙ��u��5u�m9ı,K��w[ND�,K���3iȖ%�by�����Kı/������NJrS��}��6�W�2�]�"X�%��{ޙ��Kı<����r%�bX��{�m9ı,K��u���NJrS��}�=���:�B�3iȖ%�by�����Kİ����ߵ��%�bX�������bX�'��zfӑ,K���v�r�ff�[��\�z�Bn�1�V�|5�#h�DҲ������,#ȍ�B�B�$�y���^B�/����r%�bX���w6��bX�'��zf��<��,K�����9ı,O��~'�f��Ms5��"X�%�����ӑ,K��=�L�r%�bX��]��r%�bX��{�m9^B���~����`����ږ%�b{���m9ı,O3��m9��!��)kHJ+R|��K�s��r%�bX��~�χ%9)�NO�F��{����jf�r%�g�RD�~���"X�%�~���m9ı,K��w[ND�,K�����r%�bX��ӧ3)��̖�R̗5��"X�%��{��ӑ,KĿ}�u��Kı=�~�ͧ"X�%�|�{��"X�%����$�K��xՔ���9(�m՞�p�px��:M�wk�vl^ɒ�lB�eY�V�����/!xX���bX�'��ݙ��Kı/�w��~	�L�bX�g߿fӑ,�%9;�=�M��欭W�O�%ı/�vw[NC��k���b_���m9ı,N�{�6��bX�%��|��rS������{xK�͗hb�W[ND�,K��{��"X�%��{�siȖ%�b_~���r%�bX�ϻ;��"X�%��{��2d�v�Ff]k[ND�,K����ӑ,Kľ��u��Kı/�w�[ND�,��τL��o{�u��Kı<����62c`�����rS����{�u��Kı/�w�[ND�,K��{��"X�%�~���iȖ%�b{�{fݵ����ɲ��.S,!5����m�>����B#X�a1�Z�:�G�pZL�Z�ӑ,Kľ{��m9ı,K���bX�%�ﻭ�"X�%�}���iȟ��D�=�&���٩sR�5�L�j�iȖ%�b_{�����bX�%�ﻭ�"X�%�}���iȖ%�b_=�n���bX�'{����f�K�]jdə�m9ı,K��w[ND�,K����ӑ,Kľ{��m9ı,K���bX�'�}K;fsY�5��5sZ�r%�bX�߾�bX�%����iȖ%�b_;�u��Kı/����r%�bX�a$�}�-˗Z��WZ�ӑ,Kľ���m9ı,?*G=����yı,K߿~�ӑ,KĿ{�u��Kı:��P�A��	36v9΅h�lqCSB�F)H%���
�mOB�Pj�ݰ������Q�![yvLd�i�q�m�I��ۆ${/�b1�`8kE��1�9��f����e�k�.-���u$k�$tګF�`K
���	6��I�~�v��F"�؝� g���8IVˇ�#0U��:�:�4mn2��'�ՐHf샊�Xy���b�چ�X"�nɥ�v9�?�$�,�w�i�it�#3�1�F�cD\kű�Bu�,��8�Є� m�ym2�8��X��=��%�b_�~�bX�%���[ND�,K����ӑ,KĽ��u��Kı<�wa.e̓٨��kZ�r%�bX��w��r%�bX��~�bX�%�{;��"X�%�|���ӑ?��2%��?I����eɖ-�k[ND�,K����ӑ,KĽ�gu��KQXdL�}����"X�%�{�{��"X�%��MR���jj�Mj�ֶ��bX�'���u��?G"dK��kiȖ%�b_���[ND�,K���[ND�,K�ɢ�gsR�ї5ul�f���Kı/~���r%�bX��w��r%�bX�����r%�bX�g{��ӑ,K����w�5�f,1����܄�,����B��SMr�xR�-�!�(,�R4�
�I�����%�b_���[ND�,K���[ND�,K��s��~c�L�bX��{����NJrS��}����9�Դ�m9ı,K�{�m9�P�Q< �1F�
DZ�$��2B �  RV)H�Q0 <�Ȗ's}�u��Kı/{��iȖ%�b^���i��rS���� �零ܺZ��|��%�bX�g{��ӑ,KĽ���iȖ?� �L�w��m9ı,K�����r%�bX�����$�.�5s	���k[ND�,K��w[ND�,K��{�ND�,K��w[ND�,K��s��r%�bX����L��[gl�fk3Z�r%�bX�ϻ��r%�bX�~�bX�'��s��r%�bX����m9ı,N�{.L��kY)��"75q�m���W=���2۲�]n��)	����Z�k��Yv]�'o!y�D�w��iȖ%�b}��w[ND�,K�߻��"X�%����ͧ"X�%9?��{n�D¯��JrS���;��bX�%��w[ND�,K��{�ND�,K�߻��"X�0���V���5e��\�󓷐��K�߻��"X�%����ͧ"X�::?5#J��IW�l\)��b@<=�b_��涜�bX�'���~�ӑ,K��M�&.�5��W�N�B�NB�}���8r%�bX�����r%�bX�g{��ӑ,K��w��ӑ,K��R�ٜ�h�e��Lֶ��bX�%�~�bX�'��{�m9ı,K���m9ı,O��y��Kı=�����vιG�|���2��͑x���U��7#�������fK){�Ia-I��jt]m<�bX�'s��k[ND�,K��w[ND�,K�{�m9ı,K����O�%9)�NO�}�=�-��qv�ֵ��Kı/{�u�� T�$O��t��H$�~�H���٤����%9>��JSm}Ů�g;�ND�,K�{�m9ı,K���m9ı,O���Z�r%�bX�����r%�bX�gN����tXh�Y��"X�( X�����r%�bX�g{�kiȖ%�bw;�siȖ%��Ob������ͧ"X�%��f�;���SZ�Z���JrS������kiȖ%�bw;�siȖ%�bw=�siȖ%�b^���iȖ%�b}�ao��+�l���J
T��He��mmwWJ�C���l>���g�ݏIՅ�jٚ�kiȖ%�bw>����Kı;�w���Kı/}�u��"șı;��g�m9ı,O���f�2�%�j�kY���Kı;�w���Kı/��u��Kı>��;��"X�%��u�ݧ -�bX���Y�3�����R�iȖ%�b_���iȖ%�b}��w[ND�,K�뽻ND�,K��{�ND�,K�	=��2�3Y.�sZͧ"X�~ dN������"X�%����~�ND�,K��{�ND�,P�;��siȖ%�g'پ�{Mn��G
��'Ò���;�w�iȖ'쩑?g~ͧ"X�%��?~��ND�,K���ӑ,K�������4�Eɓ5����	M3��n�s�`��p�Sf[(*jQ ��Ws,Ԭ� 06xM+1�[nh2��,[�[�6ik6�ඊ2�V8���;$����ۓ&�5������Er������\���Ց6�D��Vӳ�O�˩]W
Pdt��V=�j����ɻJ�~os���%`*ʐv*���M��q��wk��$c/m��f�{l� ��@����\���f�&a��N��7g�Ng{k:ŗ�X'���q�<�����Sd�vጧ�Oo!y�^O3��fӑ,K��w�ͧ"X�%�{�N�a�A DȖ%����~�ND�,K�~���0�m�2&f��ND�,K���6��bX�%��;��"X�%��뽻ND�,K��{�ND��TȖ'��V��c�2]]K�f�iȖ%�b_��~�ӑ,K��u�ݧ"X�R&Dȟ���fӑ,K����~ͧ"X�%��f�~%Թ��S3SZ�r%�bX��۴�Kı;�w���Kı;��siȖ%�b_���m9ı,O}��̙.j�kV�j�9ı,N���m9ı,���6��bX�%����iȖ%�bw��nӑ,K���l�e�:IM��0�*YN�+v�7�X��,tĭ�b��ia`�@�i����r|9)�NK���6��bX�%����iȖ%�bw��nӑ,K��>�siȖ%�/'�K}>��5�+.󓷐��K��ou��3�@�(@��"`2D� ���	�Uv��Ȗ'|�|�ND�,K�뽻ND�,K���6���ʙ9)��n�?Spg.6j����%�b~��߮ӑ,K���fӑ,K��w�ͧ"X�%�|���m9ı,O;��f\%�م�W%֮ӑ,K?)2'��s��r%�bX����ٴ�Kı/�}{��"X�%��뽻ND�,K��N�ƚ3)�5��ND�,K���6��bX�%��u��Kı;�w�iȖ%�by�w�iȖ%�b~��y����W4k5.��4]P�6�lgq���(ۓL�<�[��M3H�@n,ێ�f�F���Oא���/!�{kiȖ%�bw��nӑ,K���nӑ,K��w�ͧ"X�%���/��8�L9 �����^B��{��m9ı,O;���9ı,N�{��r%�bX��g{�� %�o'������Q��.O9;y�^B'�뽻ND�,K���6��c���}=��$�cKJEu$�P�R�/�0��P$�YIR���%����!"@�! ӭe��X0���HCK��Y!hQ�=����8��ˬM�D`p�`Ñ>y�<7�%%��#˄F�T�I`f�0�R�bČHG-��@ц��%�$!|%r���+,��B��y��t�CF��ٲRxy�E���B��bD<!�9�Q�L���햷E�!�4e Њb��v�mE}S�H���<�;S�D�>B�x(��^*��MD����m9ı,N�]��r%�bX������kZ�p�L˭]�"X�%���{�ND�,K��Ӻ�r%�bX��۴�Kı<�۴�Kı=�'����Zfk-�nkY��Kı/��;��"X�%��뽻ND�,K�뽻ND�,K���6��bX�'�O�fK�W$ֳw[<��u���X��nTV��f���Bus�gP�%4K��*U��j����^B%��뽻ND�,K�߻�ND�,K���6��bX�%｝�ӑ,K��]�fd�'l�L�˭]�"X�%����ͧ!��L�b~�߿fӑ,KĿ��?kiȖ%�bw��nӑ,K��;>�i�\pѩ�Y��fӑ,K��w�ͧ"X�%�{�gu��Kı;�w�iȖ%�bw;�siÒ���'��:n{w�E�s���%�g�=����ӑ,K���_�]�"X�%����ݧ"X��jKP������y�ND�,K��R�7�cA͎Z����%9)��{v��bX�'{���9ı,N�{��r%�bX����[ND�,K�������^�2F�5��k<��Wi�v��)��Z^��B����P%�ѕLj��i5���r%�bX����r%�bX������Kı/��s[ND�,K��{v��bX�'��a�9��j��.��WiȖ%�bw;��Ӑ�*��,K�������bX�'�����9ı,N�_v�9�&TȖ'�'����KK�̺-�k6��bX�%����[ND�,K��{v��bX�'s߻�ND�,K���6��bX�'L�Nܸj�&����榵��Kı;�w�iȖ%�bw=����Kı;��siȖ%�b^���bX�'�������L��%�Z�ND�,K���ͧ"X�%��?�����yı,K������Kı;�}۴�Kı6*�xk �*�����o�[*�Ʈ�Wl�.J�lg��a2f��&.t~�ǥm��gD,�@]1��6i���lR̺8�&��[�q[�h�B��@����Cs���\(s��x�[���ȓ�B�m�N�n�:��@��\8��nr���r�8�K�d�m�iD2��`,�{vm�X;\F9-˝u�3!
��_npW��B۵!�.2�Q�κ˸<U�P�ӓ��9g'8]��fa뵹�|�6�B9�1l6��W��3מ�N�n5k����t"��v���Κ���Kı;����r%�bX���;��"X�%����ݧ"X�%�{�{��"X�%���Yُn��5u.��ͧ"X�%�{�Ӻ�r%�bX����r%�bX�����r%�bX�����r%�bX��Vt�&��4�j�[ND�,K��ݻND�,K��{�ND�,K���ݧ"X�%�{�Ӻ�r%�bX��|v��.�t]j�Z֮ӑ,K?���ȟ���ٴ�Kı?g��ͧ"X�%�|�׺�r%�bX����r%�c��D���~항4�˼��rS������{�x��bX�%�^�iȖ%�bw���iȖ%�bw=�siȖ%�bw�:��o�:�G!;�l�s�qdޠ㵮� �6�\�8���u��q��a/����bX�%�^�iȖ%�bw���iȖ%�bw=�sa�y"X�'���ٴ�Kı?����Z,�sYu��jk[ND�,K��ݻNB/� F�N�j%����ͧ"X�%��w�ͧ"X�%�{�Ӻ�r%�bX�w�32fa�&jS%�5v��bX�'s��6��bX�'s�w6��c�P�Dȗ�ݟ���Kı?~�]�"X�%��vO�nBf7S+��]k6��bX�'s�w6��bX�%�N�iȖ%�bw���iȖ%�bw=�siȖ%�bw�Vw;p՗���Y��r%�bX���;��"X�%����ͧ"X�%�{�{��"X�%����͟��L�bX������5�$�˓��\ԏ.6��zC]��;��,vƎM(n��0Z7�1��4ζh:F�����%8X���߳iȖ%�b^���iȖ%�bw>����Kı/}�w[ND�,�/'����t�a��K6]�'o!y
�%��bX�'sﻛND�,K�߻u��Kı;�����O�S���}��6V���K����NK������r%�bX���ۭ�"X�3��T1��$C�"y���fӑ,KĿ�}�[ND�,K�#�צL��f]6浛ND�,�(�2&~������bX�'���ٴ�Kı/{��iȖ%�bw;�siȖ%�bt�~v��2�Uʹ���NJrS��_�v��bX�%�{�m9ı,N�~�m9ı,K�{��ӑ,K��w�|�aA��[z�\�6ψ{Wv��;�[�lEzF������wOj�a�ӑ,KĽ�{��"X�%����ͧ"X�%�|�{��r%�bX�������%9)�߯��mu��o2�ֶ��bX�'s�w6����L�b_~���r%�bX��k��ӑ,KĿw��ӑ?eL�b_ߥ��7�2ᚹ.��ͧ"X�%�}���[ND�,K��ݻND�,K�߻��"X�%����ͧ"X�%���l�3�i��5�5��m9ĳ�������9ı,K��kiȖ%�bw;�siȖ%���AD�BEC`�S[�~�/��r%�bX��t�嚷.���Z�ֵ���Kı/{�u��Kı;�����Kı/}��bX�'{��v��bX�'���ú�歞;]aYΖ]qѴ	�\��ݾ�g��/���rth�Ժ���1M,{������O����iȖ%�b^���m9ı,N�_v�9ı,K���m9ı,O0����-.k2�5��r%�bX���w[ND�,K��ݻND�,K��w[ND�,K�߻�ND�,Jr{7ޞ�]�;kr/��JrS�����ݧ"X�%�{߻��"X� �Dȟ��fӑ,KĿ��?kiȖ%�by߮�\��ja�˚�ND�,K��w[ND�,K�߻�ND�,K����iȖ%��fD��}�vχ%9)�NO}�\kuɗ9|�Ȗ%�bw;�siȖ%�a��w�߮��D�,K��w��r%�bX�����r%�bX���-$I�|z�q�Jٹ��Bq;sv#"5z7c1�����F�;<�0ÜJA9�ā6ZT�/��O��-�L��n7�DѭH@q&B'F�qX;�f��1�;;�2Qخ�v�ˡ�Ij*�;nz�L`"%���V7Ri��^��,�q����5E��x7Rn�˫��eM3-�8۰K�͝��U�v��ų�J��k<�	�M�=mC@vْ؅�v����s��/��`��]��䭵`i�]J�r�;�=���\vEn�5�� ��m�qbh��W�~��%�bX��~�u��Kı;�}۴�Kı/{��a� �DȖ%��?w�m9ı,N���?���Manhֵ���"X�%����ͧ!� #�2%��?~��ND�,K�~���r%�bX����[ND�*dK�;g[��5�Ya�ֳiȖ%�bw;��ӑ,K��w��ӑ,KĽ����r%�bX�����r%�bX�������չ��,ֵ�ND�,K�߻�ND�,K����iȖ%�bw���iȖ%�bw=�siȖ%�by�~�w!isY�M��fӑ,Kľw��m9ı,N�_v�9ı,N��m9ı,N�~�m9ı,K�O~��a��ϭ��N�k�Cš}Zۮ��;6ې��/<�	�@֚�ƫ566E󓷐�bX����r%�bX�����r%�bX�����r%�bX����[ND�,K��we�ræ�V�e�5v��bX�%���[NB!Az���Q7��{�6��bX�%��u��Kı;�}۴�O�TȖ'{�߭�2�rI�ֲ浴�Kı?~��m9ı,O}���"X�%����ݧ"X�%�~���iȖ%�bw�Vw,;����kV��m9ı,O}�s�ӑ,K��u�nӑ,K��>�siȖ%�������iȖ%�b~Β������*��r|9)�NJr{p�Kı>ϻ��r%�bX�}�y��Kı=���6��bX�'�~�?~����Ř�u��� ZR�;u���>�ـ]^����mM�K��k-�[�O�,KĽ����r%�bX����ӑ,K������q6	"w�wI�0''�����h�݋�_' N@���~�n'bX�'����ӑ,K��~�fӑ,KĿ}��iȖ%�by�>���Z]k34��kiȖ%�b{�{xm9ı,N���m9ǿ"S�V&��&�^��ӑ,K��w�ͧ"X�%��I�ӥəur]kY�sYtm9ı,N��m9ı,K���bX�'sﻛND�,�L��ߧ��"X�%���ݖe��.�.fe�fӑ,KĿ{��iȖ%�a�V?���ͧ�,K���߳�ӑ,K��{��ӑ,K��w�s+��91i^���q��}��b�:�ce']�����g�Ύֲ��w1��,K��}�siȖ%�b{�{xm9ı,N��m9ı,O�ﻛ��rS������{}0f�m\��,K������r%�bX��{��r%�bX�g�w6��bX�'sﻛND��TȖ%��i?���5�K�ֵ�Ѵ�Kı?g߿fӑ,K��>����Kı;�}��r%�bX�����"X�%�糳��jY��,�!u�fӑ,K$����ӑ,K��}�siȖ%�by�{xm9İ?mq�\���~��ND�,Kﾓ�����v.�9�r|9)�NJr{�}��r%�bX�{��ND�,K��{�ND�,K����ӑ,K��~`���)�v繮;��c�i ��۬���ō�	D���f���ݍ۷;�;�ok6��bX�'��w�ӑ,K��{��ӑ,K��=�����O"dK������r%�bX�����.]a�Z�̹��6��bX�'s��6��bX�'���ͧ"X�%�����ӑ,K������r%�bX����f\��sE��̹��r%�bX�Ͼ�bX�'sﻛND�,K�~���Kı;�����Kı<�w��%��&h3Z���ӑ,K��}�siȖ%�by�ݼ6��bX�'s��6��bX�'���ͧ"X�%��MYܤ/f�Meֳ֭Y��Kı<���6��bX�'s��6��bX�'���ͧ"X�%�����ӑ,K���}P9XB�`�XI	4������>b�ܙ��E(��� 2�!4n�ܤ�ټ/�	'8Pp�L��'G��Nm��%����7�<��y���܌���a�P!�8�.k�Rp�81;�Fb�	L�ɲG�^�U��H�9��H^J�'�$&���a>$y�����1OM0��������ՙ�x���P�qu�{���S�E�R�b�OI������ߜ�o�P�/�ڛ�����Ғqik���5�Duu��@��,%-`xSe!C4o}��w�𡬾�
�5�O<�vm������C�I�o�9�%
�X�xy��	��I3������8���@�]����H$R&�)�l"�g��y6IP�H��dޗxP�=�Z�j_<}�:�[ނ�e�l�����l�.JBc��;#����kC �`�N�\��|��\.atl���2	�1�`���՘���]@���@hBbl��}ٵ���c.x0�8R!8������[.�w�I�Μ��i���/����U�*ճU�UUQ�mUKߞ=��*�mj���Y��<*V�n
�H\.I�)@�Z��cI�4*UR�� �T��ܩ�۠ ��$�kk�,�v<sMϋ�s�M/1�9��ly�f�-�)v��[�z�@꣣W�Z&1ے�M���c��1�biQ��#`Ğ^ݬ��x�e �S$��[�����az źs4�1�u*lۈ괹.Ë�lP��]��WM�f��v��8��S�&]�[��J�p�fw�Ԫ�(���ѭ\�3�@p���#���q���jFݽlN9{:�,X���z�pk<x���8�^TTq�Qe�aw��w�r]��1�\��.wb���J�8sj�@�G�Oi+t���{W8U�r=��ZUH��.�K�L����ud�:��;%�NU	�����Δz�ֻxx@���1��mwgJ�d�J ���$�\�̰��=����k���Yz��3�lJC6���l%W%��GU�Č̊���,\<IV=�wm��v�W��=��se��Es�@m���B�k���5jDX�I�@.�tS��(��ݙ[s��R�^���Ζ�[��R�A��hm�e�=3��.ub�VCck���
���n��4��+��X6�^ۗZ��Nm�;��1:A���̜��r�6l����3���L�o ���N ȦFZn��)e]m[UUS��R�8�H:��ڳ����ڗ�ae�,�6Ő��k�ʙ�9J�C�P�,Q��v$[6�}�!�	�@�7!ۍq���Y͒1v�v��Wx�]z�{�@*��Fb�r�4�
G;-��2B38�凬0T�A{s<'��r� ���;�:�L�s�:�l�ӣ\� �㤎svص��M>�Yڼ��̽s׼[�ooA�8\��{N��Z��&:s�T�+��\UX�Wm=fik,a��.�盀�挐\�Tr���*Bc#7���U@����T�t�K�m�:r�K Ǚβ��z����z��YqwbH"�UڧɆ�Q� �  �E}QT�(�� ��T6;_�NI=�������
�1��k��@[gɣ��.�l�:�vFݐ12S��e�؄y�8��qpV�f�(0\q���B<���q��]V�,��T�Y2s�*j�U���ks�����׷��ܻ;Z���Г�
����v�5���waW�h�'�n�n�u �Cu�����dl�\kP��y��,��فCs���]��V�E��)���`"6a��p�ћ{�ss��cO<�1q�ڬF&}��5nz�WG/^���ͽ��Mud{`0��;\��ۥ6r�?�O�%9)�NOw�o8r%�bX�g�w6��bX�'sﻛND�,K�{;�iȖ%�b{���gěRj)I��9>��%9;��ݴ�Kı;�}��r%�bX�{��ND�,K��{�ND�,K�~:`�T�.�9�r|9)�NJr{��siȖ%�by�gxm9��C"dO���ٴ�Kı;�w�m9ı,O1�ǶvK���4ۚ�m9ı,O=���"X�%�{�{��"X�%��{�siȖ%�bw>����Kı<��}���ت݅��r|9)�NJr^���iȖ%�b}����r%�bX�Ͼ�m9ı,O;�g�"X�%�|~o��z"y��;J'KZ�˰s���\��iS/Hs�����sȝq�Ԙr�\WY�.k[ND�,K��ݧ"X�%�����ӑ,K���vp�r%�bX�����r%�bX�}���)�	�՚֮ӑ,K��}�si�E?E��*Ŧ�tU���"j%������K_~���}~�s�j7�h�Z)W�%N�i7n��ye`vK����~T��&�TZ.ݶӯ��U/^�׀{� �v^�Kw�_V�<�J�h�I������x{"��"�/ ��?K�4xM3�]��R;r����T+==v#�ٺ쏲BX1�,�*L��EW�:�K�;�V�~�|���xW5U�;wJ��w�w�,��9UT��=��	�y�l���8�I^�Wnݖݶڷi��=���9��8W�Ur��^~_��x���V;�
��V�+�]ڷx�#�"�/�Kw�YX��� �d�I	!���'v�x[%����,�-��vG�I��-�i�l�%b�zV�X��:��>盒�k��Y[��;`Y(4,ہ� �PU�[{�﷓ �W�{�����"�/ �
���mQh�m�n��K���xݒ��"�8�E�t�2�x�#�"�/ ��^V I#�;ݨX*ʶ�;.�m�/_���7g�V O��[�j�#C���e
����!��P�#L޾�u�'��(�=MX�[�Wn��b��	$xݑ�I/ ٲ�SV�.Ye[V�m�'[�q^0s��v�n"���+��3:�X�T�۶�n�n��u�H��#�"�^�ݍ��:WV��E6]Yjշ��<�\�H���vz� M��vC$�2�;8�۶��K����� wdx��R������n��؞�r, ���[%�-
������Cm<��XV�x�����x�^�
��q*V�-��$Z	�l��æ�2]jb���Er�YX�v��q��q��[FN�<;s����7m�̊����o�H�8{=i����:5�����BZXB�F�e5Y�˳�i�XqtiBb[\-�)�aM+n�����%�\�+L$[f�qvhM��èѥ�Ja��$�Z���h����;�6^w{UnR0���+��km��*K��b3�$,q��ѓ�� 8�}cA]��y��榶�]�6���psۦ�B� ��l���Ͳ�`AqH�tJ�w:�[�������K��G�v\� �)EB2��N˺���d���A'�<���j�/=Ď�j��x
m���w�yy��"�5I/ ղ^�ڈ.�n��m�i��ˑ`��d�r�T��/<��E�_��.��Wv� n�x���{xeȰ���z9�n�S-�M��lKp�s�IX��T��V2�T�!���V�`�B\�i�m��K��Q��"�ݏ �- �IY)
ӵm��{y����ͪ���߼��y�d� �`�[R�6��]�j�x�Ȱ{#��9�$o���/<�'dUucC�J�0{#�� }أ�7c�6"#*۴컢����G�{��*�w���$���;*sn���u�����`���㎧����<W�r�u�qH�8�	lX���[o||���`�G�I{�I$�!�wm�ݶ�n�x�<�vG�I }5G�ou:�k��]Պ˶�$�Ͼ��Ͼ�[�a�%�A""�×\�9����^x��� �مЩi��(wn��� }أ�7nE����Jo��B� �RV{�]�[������ odxٱ���}�`%wG��vm�7h��H\s[=�z��wYD���)e��H�����.m7�onE�� vH�U�|���y�P��U|��&���=ʤ�}�< ��y��"�$�B���i;.�m� ��݊<v�X���.ur!D��v��\�UU%�E�E'� 'dx��U*�U�UD�So�~�����'���:j�Z��v�ݦ�[%�� ;$x�~޾���zyŶ\�h2��ZWl��.Wkn��=��e�I�N�uދAp�͡+��]�w��< ��݊<T����.��U��aC�v� l��݊<T��{#��ďW�@/���WhV�x����5I/ 7�< �#�$�TK%�n�[I�;M�� l��d��\�%���l=I:�%j����cm�͏ �*���� �����+*���r�+��� ���KEfM�/Թ�+�t٩�m�K@-�Pd�v]��v�<u��?��&{Z�qQ9v6_#�n�&,	��Ua"�f�m�Y�v�[�:�9����F�@w��]�����ڛ����9ӵ=�l��M���kYF5Νʚ�c�q�m�v.۸��4	�����V�w�Y�i�]J��
Y�[�#�q:����ג�Dz7�ۧ�e�K��κ��j��?�윓��{)<��6�bm��jkR�-B�3��~n��Yv��0����ֺ��n�k��^�w�> |��׀�< ٱ�.uPJ"[�v� }�G��< ٱ�d� :n�)�V�m۶�M7�ul��6< ����<{�خ�\J�H�o 6lxݑ��xݑ�ݘ]	Z��Nv�xݑ��xݑ�͏ t�4�U�C�}+����L�����%�BZ`q�K�j����d�ܘ��`J4-1j�]ir���w^��L��vĨR2Ǭ�fkY�r�[�O=��oıQ�C�Q��s��~�r�{|��<��H�z���E��)��v�x��V wdx�� n��	��b��N˺m� vlx�� odx����ՀuT%�z��V:�����lQ��G�lٕ����B�ujٵ�]����A�pn�1Φ�Mu�` �K���-�	.��cr��s�ի�����6l��͏ܪ���^x��,�]����bV��f̬UUT�vlx�< ����'vat%j�m;
��	ݏ >�G�O��U�N�8T`A��#r����1�a�O 2!�1��$X�a�� �@K�o���$��l�DȌb�-P0"(e)`�DJ�Z�eS[��䡧(kV�H,b�i6ko�@�$X<8���G�~&b9͍�f&Ӏ̮Ѹ`yp/��p�����4�BXIt�i��mf���5BZ-�z>��싴�|#��cl�! �,eČG5� �9T*tR3_C����ȅ&D�,pO�/!���L'�$$����69E��Y�y���Pq\�!��#�G0�#��rfi��kO.B��2y��k��.�JJf�kN �"��}�h�6}(BXch����"�0�qPO�"|	�9�>6�֧�i�W�H�|��<�WH�p�#�`���W�w��ݞ��7bC@�bQ��	ݷ�H���&̬�Uħ���b@��.��7m�]��fǀI�+ 6lx�<��A��*��(��c]w'�X�j�^Y�#�1Zh8sm��e�7\�Xd��������< ٱ��~�9_ '��� ��<awWc*��u��� >أ���fV�-��;�մ+M� �b� $���X;#�7j!�m[���mZi� ����X���nN�#�E�@ؖW"i����$���&!�E:�s�y��{ڝ��^L�ċ���X���݊< ���Us� ����]i1Eƕ"�ˡe#r�z�8����㳧=,\9�V��n�1�PKj&gm	����xٱ���J*��s���V���Qi/[V1	ݷ�݉窪�	��o�� ����\�URG�b@��[�6��i����;$��	� ov'�vjw.��o���[o�\����� ��� 7�'�� w��1U�[WI�M]��� 7�'�v<d�XW�WQUG9A������,���� ;S}[����Ӆލ�,�}��+�\Es�.YSi�ܬ`o����V��݂��l���cl4v8Z�`��7�+h��A�j<]�Z�]q<����WAs��{u5=x��Nlc�/�� Kn��f���֋��;�@�lz�j7	M��Q�p�:vq�ѯ!���H��ɭt�Mfk1#`���g�a����'$��?��$�!|/�)biK�i<X���z5fY�ێ�z��3Ջ���-�!�,P�HA�����[������ M���e���y�$�!���.�tح��I�L� �#����Uq#���%uj�<����$���d� ;6 6H��2�%j�cT�.�`� vl l���e`H��TZJ[T����̓��<vL� �#�>R���E�N���.�c]p��ȵ�����r�{OPi�ۇ=�8#�a*�an�6퍶ǀ$x�X�G���ؐ��'vںM��\ַ$�߾ٸȂ$��X,R,Y��$������< �#�<�e/;�v�n�aN��|=�< ��< �G������5Q�ԁ��&�i����H��e`�< �v�M]4�v���� I#�6I��H�f��d�����h(��L	h�Xu�y�gc՗Y|���U�t�ل:�N���T����%i����V I#���H��2Ą���:�[� �G�6 6H��ef�GcI;�U�K�tڤ�����$x{�F B!���� s����7 ~�����Y{{�tȪ����$x�X�#�̓�;ؐK�[v�t7c�m��e`� ;$���<a	\�һMR(LEO8u���3��=g�7Tg�i����g��m��v�t�WwJ�l�)�۬ ݑ�d���G�nɕ�!�DP�wN�C�v� wd��$xvL� �#�:�v�N�i��7M��o 6H��X�G��Q�cV�tXTl\��m�f̬ �#�:�J���E@ŒBH�@}PD���y��s�fUҤ���:�[� �#�?s�۞�_����;�e`�r��=�[����fsuv���%Z�3�y���s�eY箼���(��&
9"�v^�}>����	�<�&W�\���<ޱR����ݲ�n� &���X6G�ul�y��D�$�E[�c����g���dxy-Sޫ�Oy����ceSa�3��I%���_ �=� ����2���������v�ղU�ݏ �ɕ�Ͼ�䞃H��$�����B�NS���7q�4�XFf	B��s��y��^���nݚ.�sȷJ�dC��X[�����b���k�����3����۞^n��F7!��<��Q�۠m�ֻj�t�N+K�sw(<v�TX.ȴb�x��x�3��n䲜1�m�	�-lc�!�[tQp_�(o&4б�c�k��m��fT�5�0RfY��bV!`�6�F���=��f�[��Q՟��������g\�5���SV��ea6�u���0vԔ�y�,{v�(ty�3p78�3j�aVn�w��_ ��{��vG�j�*�	�݂��Upk�%m��wd��	�ղU�ݏ ��ʺT����i�4]��	��d��	��&V�ē���n��wm���w�v<�L� ���lT�Iv���|wx7c�;$��	����x�r��|�@�~�w-�F,-�nز+��n-���Nl�3I���a)e�!�h�uuJ��U~��}��	����x7c�	�Kv�K�q������Fs�{'$%��:]�MB� ,Y]`��5�R�~0	�@�����W����;$��4�(��Cm�m��ax;���e`�ǀ7IN�tZM�t+e��ǀvI����{�M�]
�%j�g,J�wd��	ݏ ���`���>߽��ֹ[�ۘZ�P�n1�s��U�K
u�7e.��X��@ܧu�M�+t�C�i�u�v<�{��ݓ+ �ē�X��M�[�o ���`�ǀwd��	ݏ ��ID�I��n�� N�xvL�>�S�c�D��X� �Aw��}�ne�԰��E8SL�I�lc���X;��ے� N�x7In��uwcN�`�ǀwnJX;���2�ܪ�=��W�Rwv�۠�/Dbmv����1�=��x1!"t�8q�#��+��t;`$�g�j��^ N���X�p�5V�)1ݺV�cN�n� $��R6���$��d��$�]V�R�ĭ���2�	��j�*�nǀwve]*���ZN�ݻn��%�[%^ M��>�W6�$�BE�Ɠ��>�5 ��IF֨bY���,(���'�g����{;up�,^��mq��x��� &���2�	�"�?r��g��}NؒwvS��h�Э(X�u؉�ʛG%�k�� �a,l��*�e�S��|��_����;$��&܋ ղU�mD��I�Վ�����;�e`nE�6��	�< �t�Ui�i�N�;�u�E�^ lڏ &���2�M�J.�i��wv��z���SҼ���x͙X[%�����v閛bn��	� ��r���] ����k^����*�U�� ��� @U� ��PW�  *��U�Ҩ���A_� �ň�"� �� ���"���"��� �"�U`���"�H",(��",b��", �����`�AW�@_�� *��U��U@^ 
�� @U��� _� ����W�  *�  *��1AY&SYԹ�O ��Y�hP��3'� a�O������fV��TY� ۡ�]Av�w#e��-��  �m�U���:�GM������;�]4V�N�u��:*�AA��ֺj�
va����IUkK1�R �]��PPm�����'@  ��     � *Ko;
A��6�s�;zM)J=��A��
;�p�����7M�������;�{��<g��>�s�d��   @kﻠ��W�=�s���w>�U�v�lNں��{�
��Y���}�Y����cٺ����O�=u��JJ���E@�{�Ϋ�>�޳����{^m������^����G��C�`u���_})���π@�}�x  ����� ��o�;g�d��c��`z���]<���q�|��v�=����@�����J���w�y{�'m�����,���}�{�J�y����2G{�W��>y��6����-k�=�x �0��8�{�ן}O�G[�>�x'G����`t��p���DR����q���� {�PU�A��$�5�{��4��=���aץ�� ���{�w�[����2=�p��������o�|�<A�� ���݀}���m�|@;����:w�����m�o�nϠ��N��� ��<   a�!�h��o����R�=m����}�����Kw: x�����M)n��fΚ)��r��=��4�r��� ����4�   �.�Ju� {�^�Δ��� n�
(��R���zR�^�^�{�ܥ)N��(�e(n� ;�Ҕ� ��қjR��  "{JTyD @�MR����A�F�"~MU)'��  ��5Q1J� 4ha!M�)"�4<Sy\�_����V]s?�?�ZI%R�+��6��� *�� ��"*�� ����j�
� U`��dATS�������������T�nM~�>/�٭��Yo��^���HI"R-���/��)��q�'����!߹]��3�4tѯ�N0�Y
�/�pWǟZk���w�LT�ic�˭��oA3Y��MOġ)���Z6VoG�M�g�}?|p��0��$!k�#5�jvX�����=u{�8�֙�B@�$�����MԶ4,1e�O�,���?{�y=n�L�~�	u�k���IK-
_ٍ�k�.�Xd���B匄E�7)k�3D���>�滾n�������(��.��Z�so��*X��,�����0~"� D#L��a�"B	sF�c�����u����L
a@�(�*���j�~~	>�B��
��p������vXHs�!�'��@c�"K����l?]sY�^o2vrV;y�$������otGyJN��~�Ce{��^�P�X����[YmBŐ���D�D���Bc�XI��6��3ء �a:�0�X�Hh$i��+
°�c\��棘\�5�{9�������GB�	��{V�"
� 8q������4}!��#]nс�)��sF�I�A
��,j�J¶��/}��\]�����BY
��;��[��<��/9IH]�߬�w��e+��\�t��Q��Ժ\�oq�
�?��ߕm�K�%{��pTK����b��5�f��]oz#)��~�ȑ"���ɇp���~���r}w[���b�X�n�w�aB̢��)U�9��}�X���l��4�%/�͂we�w+n�g�Jǫ�$N�����~�k?o��R�M�͒��?4�#�1�X�Fw�_����W ���H�!&�	I�.K��B�(}sa3�w���2nn܄�bƥs����{w	Ä�๐X:�;u��L$�9���3Fj��!�S�l���QWt,T�uԎ�mt��X�	��ϱ����O��ΊW�e��������o�f��55������� p����U�������1y�gU �'?k����_���H�����.�O����7)�I���� h���,hZgMf܃�i�) ��5����O��afb}�X[�_���O��J}��Ч I%�{�'������a��q�su N���s��9{�y$�!%�')i���i��U�������^BJ��5L5�Y��%�N�w=����)IB�������Щ<T��ӏ��8q6�w�߶�^^��z�u���VWv���|j��HV"\_����h �Y�o�9��9�e�0����W�q�p�}����7�9��y�Е�R?��&������D5��D�bB20 7?k?�l4r&ر HXb�1�B"A D�a��oƳw�\�l�J0�(\�Y��?c��!?sy�e��M~��%~� �B����M��$a/�5~�����p�}����������1�-���a�P�L6�u����fKy7�o�~�9��H�1 Hɛw�YtA&�>����M������w5n�8�8K��.y	)�g��!� � �;ñ�m���B�B�dd$�kX[ ��F�Re�T�1���L Hed�����R�JwY,����\�l���U±йV��T�aE.p���U�}���n�B|�4�O���r���+�L���7r4�fN�tKIN��X^�
�2���d~��\7Ēf��8�?of�I59��7�s�c���gA�D.8w�rdc�\H�36n�d���
@�H���љ��,!	`���s����-�Wǽ(���%Ā���R�t���S��hҗ��f���P�jI H$$�,�#�d'�Lh��m3�ҲYA������z��3�%�`~ V,�IB�ځ���u`ɧ\,e{au���~�f'�(Hw��*a�y�l��~�'ۚ����F������	��c��ߌ��o�ͽ8P(��%,���,ϹL�����HW�5��#X�n0e��T�b^�|�ξ�M�0�k�6 Y�!��u
��n����z����fy��K;zN2�W<:�N��L�t�l!(B�0!���$+(F���s��o��ȩL9�ÒJa;x@j�A"����)�[\SRHHG�s��9�^���/L�HX!���cL���/\�s�R����wȌ��ד~��qw+����*�B{��>VU�y1/�˪I���oA)�4F#�G�d�n���+��k�I�{��a%��Rc�a�� !�R��{(�����ė��½o�Emes�U��g+绸�
�y�Y���K��.g��.q�f�� 1aS!�v�q��g6}�t����Rl�Yp!���/�ԌI�� Mp%��hM��S�A����Λ?r��=}��8千d������o�*0�f~�����Rnn]�)�7
aun�H��@��/
C�i�{�h�t����.S�;�'];�:$8]�c�NO����Bwz�T�\vcG���o����\��n��̷��5k��Uõu��^��Fv��_n�=F���N3	�&r�a��~.N^%BM��ϸ]m�Y�a���BA�2��{�)ۡ?�����a�_k�Sʡ}[������l�@	xNZ �c�m<���#0�%?tNwi�JI
������&�͌�m$73g!�ӧxƤ���vg�oWI)g|n-�VX{)7�~���`�G�
0�G���̚$aJi��Y5��~G�Ӽ�ak��.��f�?h�Z�� �Ͷ�g�X������{�$�I�^����i�:��8.ל�JCuIV�O�\љtv��'����T��!/�_�iӼF%Bx)�NHB]����Rx�']饝w��ߒ�5w�W*�ehS���_:헴#V�9���x�	!���4������HW-XXB%aB"jg��Ή�� D����4����)
`pa�rZ6q�L᫚�.K�	�!߾n��ٝ�ߺ�c	�!
[�JS���V�$�B1jF� �
�JK,3_������t����4�HP��0`�L�~Ӛ$��p�aXP�!vk2����Ԅ���G�@�I3QJ9 �$K@�"B���Z$"K;Ͽg98���jF$���YR,q�H�cK0%�B!HP �%!H��$���l$�3g�>�\�a�Gs�%3[!������9�d����]n�Q��	B���ވk5*JB�p�a+1�f0���qa���HH�	�f�}�ee"H�n�BS!sd8\����<��%0%�[��ԍ%��0�°
7;0�.9.��4�ԑ!A�,e!���N�1�e.�l�BrM��I�p��K�wza�C�)�l.4h�+���I"�H��!0!� T �B%!H&F,A�ŤY��0��.�W� pa$H��&�#XH�#X'������ot�L��̇-�#G�i�F�;7����|�!�՘i��J^8R�[��)f�T�	���%W+�T����!�M1B��)	$i�
��F@���	 ���*ڣ�o��w>����]�|0���iN�I=렇 r���4pe�l�K�g)@���)N�.���VW�9��o(�o�Y�w�������3�}�,�F�r��:�ġ�3*�I�2c�a�˼������Ϲf��g���|�'5���s�&����9	(K�����
a)��,$[q������5�9��L�9��IW�*�w��O2�Y�է�Q�J���M�2��';�5��Dֿ~�/�J�YH`��Fnї���U��t�k
 �x�w�[?s��t���>��/�t��7;��Xi\OM$�fg%�B]�Xf�Đ"C}�3!&���]@�uh�me+%��$!$6W?~��$n�C��7�<ͤS2=�4��U�h��5�Ca�?6꼚/ߎ$�		/e>{�p��ap����˧�;ٽ����ߎ���>�س�ˁn}��ߴ�2��:v��a���nn�m�s�Q����x��.�v��b�;��Uw��,��|;N�>�K���a�*�oy��w�o��ɟ�\bD�HT�`����� CW\�y�m�;ћp����B�0�N���.p�t�\�LM]�5�݇~���ο�sz7���𱔃�)nd/����p1��E!GF�V\�0��i�\t�ְ�m�RXД%���RR䱙�3-%��$���.F�B��	XH�4�����ieל:��!
ix�]ZC��/l�۳A�B��
��\t����0;sSXf�$ц�,)��d�5�������V`XbF��(K׹�^��CBv�6t�b�4�0�-�W5sC���G�7z�B�M�u3i(a��ƛFJ�@=�un�aJ!dЍ%�ݲ�q���׍]4 ]&�XP�{��%��N�$]0�2��h5����f��7�� ��O����)����<�K3���%΄�B���nI��wD��)�(D����s�p���Vr� ���J[���rw��H�c�?��8~��RR�XF��B!�C����w���?C0�FӁ��	q#�Hh������!��~�l!������� 0)�"H�BD����ۮ�=a��=�Ǿ�4�?�
� H��,�%H���Hi��F�Xfh]=��/P#��,��~�}��/�?2����p%�M����������3��4��hN��lK$��Ɵ�, D��Z�I���������!4�˚�3\Is}��e����澄F�%��W)
a�SJe�ֆ����#6rafndX�L�B!kHjD�dm��y;�|���ӳ�FB�B�B��B�!�H˶��$��F���ą0�RBIdѨk�p�F�	ys��=�;�n��n�:!-�й�#s�;�l ə�nFw�s��a��̤��-"p��fԧ�}���M`b�(��ZqQj�mO��'p�� ���8|~�2�G$Sߵ7��	�����BC�s�!,�)���*����UPUV*�UU^UU��{ʬUUUUUUV���*����j���X*������V������������W���������U���������������*�UUUc��UUUb��U]����[��V������fy}}=HJm�7V7{ia��Q���m�:�.dXZֲ;[;� TV�aU6�*�Z���+\SUUUUJ�I�R����G5J��3UR�NR:Z�v����6��iTw*����U&�%Y�J�UU>�Ի 4�+�j�����t��9Uv�D����@�K���8�^E�
9B�Gb��5R�W�����F�<N���̺�7!UUQt&[��A�*̶%Z��+f��\i�ڗ��nf
�E�lh���.\��ch�{ ��Nl;�8%m�vev�m�*��[�v�[�����m�����������
�`�*�PTK����k(�Tk�ғ 9)V	J��Tэ�v��\ۂ�//dw6㭵������ � ��'n�m(<��V쨛�ד�,�z�H*�rs�����������;Ԫ�µ�R�1Vj� bx@���Z��a:��M뫁Wb�k�T�s]�P��˚��+jl�%$ D+jt�R���8)]�eWu��nxj��5=��%R�aY�i�<�Ug�;��>�����)]�+�3U �
�U�v�B���Z���*RZ�[W7���s�fURZ��V�5�CU*Ժ԰�C3m�UUUTX�d �j�Vw];5UUUUaE�z����B
�h*�ڲ�����ΝU\=�Wr�	^��5��j*�ղP�m���Qn}��UmQER�5UU:�����W��R�̄��Tkc���39�R���g���Z�k�X�V4�l�UT�M.��-������Js7f�mU�3*&�iХp�H	�<�;;V԰T�V��W�AT�Cvy^|�wb�A�[��T A���sR������mS�=@K˰rF�����A�Vڮ�^B^m���P	��n�vUX إ�����ezڹ3c0��q��}[P�gں 2�.�gn]��Λ���]�k3͕mUc )+꯶T�p[�V��7a@j�VS)�28�Eq�M�5�}��<�;�OG�Z�6�댥���炴<�7c\6u[���{�=kqH4j��oZ�Tl��ѕ%�=��$����W�Z11ѹ������ԔMQ*ꝣyk���.2).�E��[m�j��+�,�A�$3�x��Z����mOA��;;��)��/��p����j���]�x7V�vW�q�
1n
[� �
ݧ�-��ת��&�rr�l�G	Jપ���%����lbϬr��ۜ����'#����\�e%v:V�]�t�6m U]U���c�5*e ,c7.]Px��ةI����"/[���w7��{Cn�͋y	o���v�� �B��{UAh��왎;Gm,<����� ��Nxuh�K���3N���1��p9e�%�]n6���e�ﯽ���c=v���ڞq�4�+r�W����J��UUT.t�w�Du@rWf����UcU����ٞ�/9�V[��s[[�],�T��n�ғ��#��ȝ=���V�U{\EU[1����� �-¶[1�D�T��#ءd�Q���:��p�\����B��ͣ��>1���R�)%I�i��ʜ͏p)�6;v�غ���T)r�q��U��ʵӚ��U]Y���mc�]�H�b��:0��:ܵ�÷PuuN �:��5�@���%j����۞�S��hA��wo����yU�%e�S˺��M����[�)�l�bұZ���4����!���[A�� m���3�1�v��F��9��EZ����Ź�.��r
���R%�v#����*�Z�@2�B�� q��@�ݹ�P<mCNhra�Rptw3�m�(N�wHMR�y�c���h퍰����_K���ZͫE6��e%�]���څ�����d-�-l�� u�K�V�Q�f+-���ݤ`� R�UAU�(�V��f�Ɣ�0,�b��v��vҭTRnI�yr�͠N�My0���G�|�;u�<�/�..S �Ԩ2�PUW@=�AR��ڷ5�6��V��ޘ�ݪ�
P+b�<F���李����$L���#2�ň 1÷@ m��9Z�����*��uOS]AUUT�A��n��1��A�K�s�T%�l�T�Ԭc�m�h^�[�(!OX@�ꝺM��Ա��a��(U�ڄ�5w ,2FQl�EU���S(�9ݹ�r��+s8c�=Yy����nNtCaz����5��S��:�$6y�n�)�.��*qF��aL<��W9l݃n˥BP2�t5�*6�K��v`��EA>��K�?x`c��l��UP�(�x� ��yxZp��ke�����j�J8�URXV�H���\G$[j���;e�� ��m�mT��Ԯ���x�\m 3�t�� ��x��U��m�wPF��.&y�v��UhӧV���J�؆�N9��%��8^�Yƀ�y\�B��R=�6�=N�n]GT�E��<ʫk��UUb)ʥjA{tn���7UUUUUUUUr�UU�6Չ �y�*�Z��UM�Y[knk�����UU��W\�vܚ��4�GgI#ƛp��8��6N4�l�$5qvv�B�mh��Ʈv}R�S0Ui�Gd"+ɛ�������[�r�VQ�ȐF��P��@f�H�}�F�L��]WU�Vzmov�p8*��z���>�Hdj�#�p�Y:�Ug���"�KU!I�꺪�Z��6�AҔ�"Ŋ
�j��썎ΰr�s�Tb� UWlS�6����/C������lUU6^Z������[�j����收�eiA����q����Y�6�yj�Z�T�X�٪���]UUUUV�jz���>`{r�mTJ�UU�/<�UUR�Ν�Z�ꢭ]J�UUU-)u�uA8Vi(8^z�^](5P]UKR�X6�UR�d�PuWUAl�UPF��:��)`L=J�F�z�YPj�U��V���A���Wk�(6�\�5A��UX��ꀶ�p��kj�r����??<�ʭU�UUUWUW[UUUT�UU�*�uU)-OcMQθl��@j������rѩ�1�����uT�R��UU��^���������Uɘ*��HEUAX��Gr��t�n��)^^�4)�J���,��kpSUUUU˲��ڞa���� -��Wj�������������)V������>��ҭF:����j�۰Bf�m��	^
��XA����j���V�Ҫ���ڡUUV @")<�UuAUUUWUUWvx�>���5+UU+]J�
�eey�5T� 7���y.̫�+Um��2	���檶�j��nX�.�UUuU]J�UU�U�V��P�UUST5;�{[�*��*�e�z��������F�bؼ���U��@)-U*�S��Vy��������ꪪ��
�����V]��
�Z��V�b�j�Yy�)ʳ�9(y���UR�5@UUUUUR�TUJ�R�����]UJ��@UUT�J��W*�W*��Ƒ�T���^j�U��t�N4Ҏ�X��i�	I����plMz�.�Pj��h�U��P ʮR�9�)vY]�ڭ��^�j��ـ������^Y	 :e��n�*����ݴL�Udz��U9J�'9[�u"��U���mUGطG�Rڱ�40���aW���j/W:����vQ�v�$�k�Jpʡ��[U�J����z�%+��Z�ڥ��䔓Fچ���J�)�@E�!���Pt@�`�p[O[�ڸ��c����m�=���ZȮ�H�4(�� �`,Pʡ:�1����50ݕ'"mW����-nq���� Z�m��J���nljn8����_Evcn�R�.V��'
p�Q	�V�Wf��9����
06�Ɏ���ԨR��	�"H�٨���#ve�ӹ#��K�صص�*�qյ�E
UH�\��+lʯ`DJ�,5�i๨�;t��;k:w����)��݉�f2^]��:^6hw��p [������*�Uջv)�=��>����Z�o�b�`*2�fS�:���N�L��$��6�N�-l�.�� �]�6�N�M���J�i�:����rmS��\ڒ��7D��4-�e�%�̄Ò��(�:�'V�l^�W��#�#I<�Um�în�*�]Xݻ8�j��UW]t�Tkm���{v��j���%UPJ�9H��J�E�N�T6�(�U[R��y�KAA5UU]��w��x��ņc`P��KUPpj:�
�����*��Z\�����<�0u�j��9�	�ej���F�����\�ݰR�T���n�L�UUR�5��Kq�uR���7���L�!�]�k��B Ŋ����*��˻F@U�ڪ�Z����yZ����ڪ�����AdYV�j��������ZU���Ke�-UUU�PUUUU ���K�ʵU�UU^�˝��^��q�U����LT�_U}U-*��@U@TUUUUU]UUUU@UR�UUVԫV�UPUUU�WU�U��Uvj�����V�UUuUUT A*�Į��++@PWUUT�TUJ�;;*�֩� 
��^Z�
�ګ`A�/N1AD��-�l�5��UW�$w�Ejj)��ZU�cWU*�UMS:*�m�eZݠ�*����V�Z��i�kj��:����fQ������Vr�����]s���[	�5c�ˈ� �J�A躭���<r�9,�U<U!Q x��!��S';\n^#���}(T]����A������4g4�k3_�� "����h��qF� D�PЩG�E�!����#���b�A���"�i�� ��	���SG�DT4�$>Mը$ �!�Q��b(;S��uQh�]����*�+�6��>D�P�DS����W��:E�6�"b*�> ��E�� 0i��x	@���b"�� u�t	
 ?"�lO�	!!	 �)�HD�0�C��M��E��9���P��T����_#���(��`�� B H(��"|+�:@@�؇N`�	�Q�ҋ��t�Ep�H�`�8�"�S�()� G�ʣ��~Oʮ�?!�;Tڨ`M (1���H	 �(�&�� blU:�_���M�J|	�*�U�aE�I>P"6 �@C�A���O�L?'��O�@d$�%v��HF ���A1 �@�R# H,-��"�*D�
��D(@�l8�>*.ƈ�U���!��@�pGH��>�,%��"KP�����J���HR���Ȱ�d��JD��m"�#BH���F	X�YB�HYE��*�RJ�
DA�+#X6��O�����A~�"��h�HH���GH�`��@>*	 �R��H���	��_���PU����*H#$A�
� �Z!�Z�*`�J	X��m�!�b5`��X�� @"V�H��Ü�H�����Z�j���A�����]mUUT���,Wnn5���$�N�������'`�Yѷn���jʩP����z�䐮!EA�իmݚ9�76��;]Uӹy�=��Ѽ��0�4%��OM�7lmـ;e͘e�-m��D2��ݚ`��ÙYwd��I�J��8\f��^m��@h�e�b�ƍ��k)��j�\d���H���B��׶��]1XSn��k���9�g<�ӻ=��n�Su��ܼ �䚛^[E\�#A��N�^G��ΰ��<�h�ջ�r��-F1Һ��@�m�;
CP4�8YW�0i82�:ݓ�݌<̚���ق
�,B�b����n�j��W��L m���3	���WD�a����\���n������ (�R�1�[����s]�
���c��n��C��R R��wG=	"�/���A����v0oR\�&Ch{�sh��g���Mx[�Hf�f�E֌㘘}��t��Cc��&zN���=��ܯ]�k���EЉ����&�a���l"��ό�)3��lZg��ʢw57��Qh�e�k��r�U񳖬��\�M��x��[E\p���F@	Y��$��X�5�C[�\wH�Yx�'M�\�6.�zM�ښ.�vsNx�ZU�Pn	�-���-�����T X��90eX.��d�V�9�	����Ejr�*l���'3N�2��8��5Vd��@\�:.RT�73�,95�����I�v�k�ͅ�aa#��X�9���+�p����/�����c��a踸N�Ico9���:����$���r�l��p��J^Z5������vCBbTļp�Ҏ�$\�їM��b��R��q��h�&U6�Urgs�6;i��K/�wNVIUkR�����������c���R�RU�J����b���)4=e�yu�-B�a1�;�9�/gf���;��5?�i�t�U4�!��tU�)�� �BPB���т�"pDЁU
�T�$�O4���e�A�cf��n���1-R�ШZ�t�R��l�{`
1�����6���cR�o
^{E�M+�ͩ�[�ۋg�{ay�H��=�'�k�s����n;p �-���{Ok�6�v;Y��2B:��bT8�9�㬋�Q^��J�i�*PN��+���ɦ�&Y,\э�c�հv,�#�Ө�hr�W@q�֬�kR�a�P����q�3 �_!�(�� �'x�9Ng!�����<w��.�ln��nkzpN�{�� �'߿}��A$����v%�bX����iȔ�%9< =C�m*�����bX�'~�ݻNB)ı,��֓q,K�����ND�,K�����NJrS����{��2�[��r%�bX�}��I��%�bw�{ͧ"X����;��7ı,Og}�u���NJrS���Y��8��gmkZ�n%�bX����iȖ%�b}�ݕ7ı,N��w6��bX�D��z^N�JrS�����;5SB�6f���Kı>��ʛ�bX�%��w[ND�,Kϻ�i7ı,N��y��Kı<"�j2��L֍�����-h�BT�C�Ǯ�@�]��x��b��r!�3�����������b_w��ӑ,Kĳ��bX�'w��r%�bX���ʛ�bX������K��,]sk��N�JrS�ĳ��Dq>")�@tD ?(Ǒ?D�9�~��Kı?}}���X�%�{���ӑ,Kı���-7V��m�V�r��G*vO��"X�%��ovT�Kı/~���r%�bX�}��I��%�b~��òh�5u���L֍�"X�%��ovT�<r&D�/��kiȖ%�bY�{ZMı,L����ӑ,KNO@���K��
S+/'G%9(�%��w[ND�,K���Q7ı,N��xm9ı,O���q,K����e��[&��2CS2e�����:��oN\����1���<͂6�k�����rjܹ�Z��Kı/}�j&�X��#�;'՜��R9H�#v^V M��ں�D�S����v�;&V�&V M���G���9I�� ���[��U�Cn�	=� ���t�T��r��F� (�.O����'~���5E �˫N貓�ݺ�	� vH�	�2��2���A[aV�;�m'm�d� �fVݓ+ $�נ;��c�W7�B��.���z�c�z�{�2��+�-���(t&���d�{6�͖��շ�I�+ �ɕ�lxݑ���
t+i��\���`ݙY��r�zy�g��	6e`�	 �Wt���B�� $���#�ܪ�%�Oe`Oe`Vʘиӧbv�Z�o >�<d�X�̬	���>r��W8�UY����7j�%��i1�N�d�X�X�G��<��W;^���L[��6ڢY�+i1�9�'B��vg���XR!o
�l���4hۯ������< ����W�'��#����V���O��� l����L�d�X�IQH"ۦ&�;V��o >�<d�Xz�������������;�J�[x�s�O{��'�� �G�$x�\�ƭݖ�k��n��e`�<�7�'{��ܓ�*�.�_�-)ޗ�"��9�c�璸s�A��>�=����o&�[6jL�#+�6x��1�͚�{�p.-���z��V�e�����g"�*=U.z����b�Y��v��.+��ZB�RRA�h�i�6���'�y<ҙh��pkV\-9�7k1*���ԅ$�p�d}���Q�����I�5�8z�l<����5��7Xv����Ǭ�jL�rwt�'��^[7��Ḁq�\� 輌=t6炷<��Y3S����svV��n�a[���
����נ;�#x�e`$��>��1�\v�ؓWwj��>[#y�Id��'d��	�<��A�J)iնՃ�ۻm��M�+ �&V M��-���%*1�Eӫ����X��T��� ==�|�F�	$��:��;n�l� �n��	�e`�e`�s�sߧ�wƮ�b��$K���9
��:��5E�읮.r���V3V�v��m�����d��;$��W+����������I��x�0�Rx��Kk$�!������&f#	ճ\�.@�c.{2����)#y�RG}�����|t�u�{��V M��)#x�2���$��m�CM���+�UIz{� ����68`I��}[!��)�e��Z��o �I�&������Oy��J�TUt����`���s$�P��&Q�Zy6��zpn����k���VeGUvUz�=}:I2�l� �I�;���|n���V�I2�l� �I�&� Ӵ�,vS��:�X6G�N^�����F��E؆���7$�&V�)[l�m����7�M�+ �L� �#��	;iՍ+v�x�2��e`����%)͉һ�j�X��e��]�+۳sÎzأ�d�와vW�w��	���u�uv�w�ě������	�<���&ɕ�mw��R��*۬ �#�>]��l�X�Y��;^��n˦���j���xV�����&V M���"K�Wn���mݶ��	�<vL� �#�u\�UUT�UT�)QC���u��;�^��4��ZM5j��;�e`�R����wny� M����zM][�����m��K���ܷg���7h�C��3�V�q�Lk�-�\h�ue۬ �#�>��w�dxvL�TR
ݻwv:b�i6��{���&V M����
��m:��i�� &���2�l� ��#������ݡ��e�x�X6G�}ۑ� M��]�&�;�J��� &��r���w����}��[�@S�� A6֩ ��T��$ d�B+Ba��3&t˫�)�2����]m��i�=S�
�����;�-�H)a.�f�y��h�RŘ�9���/cH��el�6�Ya-2�r��\\�̗�O�[s=A2�����;�����1���8���r�I�y7<��ۮ	nLg&(Ty8�V��k��xMd��6�n@�ŷt����:n�6W�`&���(z�w*�Nմm2a������3SY��am���ՂrCwWc��X]���ţ(�|���x8^u;ͺ�WN�v�]ݷ�}����� l��ݏ �wiݺM�N�n�m� N��d� 'v<��.����6�(mZ��d� 'v<���ǀv��tZN���]��Eݗ�wnGx;��w�T���)nݦ��YlN���#� ���Iv^I�E��v�/M[���E]�����0x{ ���8�S5�sN�r�m�l�m:��i�� &�x$� ����r���ׯ�X�F��]�̳5��.���������)��F!9��PŤL0B�`�mWz|��Xk�"�:���;S��"���**�o �܋ ��Ȱ������sc�ƭ��J��+M��mȰSe�wc�5M��|������Ll���Se�;��Ixշ"�>Z�*]ډ���t�F`vΫo[��/�1��{V�^�[v�8������47J�� w��Ix�ۑ`���$#	+�%�鍷�j�/ ��r,�Ix�%�<��H������c�-�[����,�I��K��rkR����o!8�o�e�i�?fe�fRX@�e�%��ov��I�H�� qb1 ,X��"??��u�H��2��|+�'�P��&3��h�#�J_�8���:���~�f~,�rw�O˼kg��!0�RT����/��fg�U~;�����-���\��o�e$Ĕ��	[T#�(8�
B��R?"i
��YL]�\�MP1003P�!R$
jJZBtͰ��hX�����1��+&�T]/u�����?B|f���ĝ�L+
�#)]����+))2��
�~%	��.hYhPfI�~ӝ3�f��� h�~w���}HзVT#�JJK+,�O����kC���_��3D�A����d�.�hq�1�!X% �%5ł�@�+�J1�,P�IA ňX�#H����[�F4�IHP%e	HP�YF�3���ѳ_����H�X �aX4%,-�%��7w��sz/d���	����8f�L�B�C�K6d���X�����ש���3�4��wk�\�k(�w���p�C��R�fE �d�?@�B�~9�~�c4忥¬�����<%�]ӋgƿY��6����$��M��M�:͢W��:����A�	��D$V���?
&
hD�=�tW�.�ɥpA�@{��}߹��<������{6 �6667������j�!�p�֮�A��@�A�=�f�A�����}��<�����w����$���������O���m����.�� �dx���s޿�ڗ<��%�u}�{�d��2ZZ�2��]�:״�[s�,A`덙{���C~U�z�_�;�꾅��9**�ou$�+��^$�ݩ���JH��rrI'��������y�����K��V��Ē[�2}��Uݤ��7�$���|�Q\����]�[sԏ$�[�i��n��>�$����$���/����~$��{<}�IE{V��P�+��	z�ʪ���z�䒞��bI.�2|���6 �"X�,�D	D�A�l��!�$�Ws����$��?y�ĩ�K��6���I}��˻m����T�������o�����m����ն��~�j���5cm�4�#�k���[��&m㕍u�C�l:���W�wcǽE��O�,�V���$��{<}�I%�7�$�se��]���f$�]��'�;i��]���I-���Uݥ����䒗�f:��߃﷾��'�߿��[�m6l�m��Ē]�����_z�R��I}�I|�F��$����
BⰡn��%��{�3Iv?_��H���%���۾��}��b��.�XUN�����_�$��W*��x$������[&3����$����k,k[�@v�R��D�ۤJ�� R\csdf�
5����������y��끔 �y՜�'N�(L=�v���g1���ڳCY\B�Ạ����
��[�f,��q�=g��\����hø�2�B���Cb�!-0���jR�kz�cP���xN�������I}<T�W]A7B{��8X�S��;�f�mpLŹ:w��=�;���>�^}�͑e2%�ղt�u/<4���\��cnU�\$]�=����gc���Ӻi�r$����x�Knl��I%�c=U��Jk����Iy\���e6����I-����ܪ�����ĒS}���H�2�{�����M�M>%l�K��7n��$�����K{1E������T�=��SĒK߽���I%�n�!�:e�lė���w7<�|�]��߲�$�^������]�{�bI%�	��Pն���I&SĒ_������=Ԓ^���%}��}��m�O7���8U��Nid)@k��r��h�w��]���wh�5��������ށm�ui��;.�>��_����Il��I%:�K�w��'���$�kj�=AHL5���k��߳��M��������fK��6L��$�ݏￕ��W�U6�����s�vڅ\um����n��#d�x�*�˻�~��䒗�e��K��z͜�Yv�AY�vߧ$�߾�=[R^����%�&Y�/s�������$��ϭ5xa [�ǫm���z�ݶ�${�{�9m��g�Ü���{�[���Oz8ϵ�.6�fR�U[��:K�t��7B��#�0It&�A�-	G�I�o��/��7n�RK���Y�$��O��H�2���'{[|�{��m��_��k�Y�-7g�$�{����\�ݢ{�OI-����ۓ,�r��%�x��T7eۮr�g}�ݶ���{�r�@r 8Pr

��.0A�V�����xo��~�M�m����s����]����3��q���I������ԥ��f$��M�W�$�\�S���$��AC���'t�!ۼ�$�I�x�K�������RIO{�!v���%����V�Ա���#�%	f��]��ؙ�r,��4cB:����������{��ff�����$���/��1��Il������Q{���o����3*�v�:9��m�I������6����������*�$�{"����'$�_���5xa�[��V�{�ﳜ�߯{�7o�3;�z��-����:��|=�ة+��n*����$���p��m�}�Ü���{�M�~���� �%A*Q�:4��4�@����R�@(�M�DȊ�@P���{�~����_~�ԗH�Zl�um��=��;�$�ɌĒ[se��I&SĒ_���=�ϥs�0b��6���S �;Y����������8"bа���fc%D�;ԒS��bI-����$��)�I-�Ӿ�����R�:ٝf3�V�[o��E���9wiz{�$����H���UWv��\(��EM��BDٔ�$��'����Uʻ���<I%<����%�ۘ�[�Wj��1%�\�=���^��bI-�E��/��+��U�����$����?��Em�:8Y�v�}���[j�\��{�߿-Ԓ?{�SĒ[��W�$��Wd�H������f-�����e+�0�,ʭsA[c-�q�C*x���3�˖'���r����Ec���Eb��ۚ����J�"���%s�O]<\��qۃ7�T�O]c�5��٪ܲ������8�1�#�+ES��.�\)��@vx�pF�l�3�Ѷ{�V�^ط���hp�����n��h���-���(��v�C�[�v���,f{��:Y���|�Ʉ��GR���VM�8xS��8��8rҐ���-,�O����g�p��M�Ԓ^�߽|�QlʼI%�$��\�;�I/\�I$��^m��J���|�Qlʼ�s����6Ҟ?~���	���[���;��9�A��o׾n\jh�n�Ia�}_|�J^�x/s��r����_|�^��I.�irTU��f�r����
���߿��-���������ݙ�o�Lϻ=��9m�wڹ�]f�X�1��wV�z���m����������$������$����$���+b��M��a[,2�LT�F&�rm�Ǭ�����67;����ܓ�N3I���(���������IwI>��BD���W����9'�M�i�R��@���I���	F!�iRZZ�d��FF�bAJJ,���%dBA@a:?���O�=�z`��,Wv^{��8�I���t����շX}��Ix{��J-��J����wV�-S�QM����K}�<-��v����+�]�����iRm��T�m����s�%{�W�w���:���sv*nN.��	���xk6Dͯ![�uڭ�|��'��R�M�ϧ'N�uˠ]"�6컰?s�<~��|}��I��ϐE�׀����a2���������O�9Wd_�~��{���fVz��#g��(N��ݕe��l�;�����/:�\I �����G�0X"� �1�L���� 24 "�� �A�Q"�a*' ��/�g�����=��znsɉ�=�69a�z����=����V��Us�]������^X��t�v�n��+ �r�U���;���v^�jP;A(.�C���\.�vz�ki^B��v��'<k�c�K-��'$��N����kg`}����v_���W�6�X�k�2��h�!�K��ܓ�����W����x���V;��r��I�%zƨn�	;�t�k ����7t�X~�UW+�*�UW����5~���	6�
�+�uch�n�=�W9UJH{��=�<��������X\O�]"�3Z�2:�h�C�m!�.�m�M�h�4m�! Rna�Q!�~�O������y,���,� jk����,�+�������߯�~S߯ ��X�g&&��S��-@�Z��I_=m{��ӼnE�#��C�������E�Ӥ����F��)+�����x[������䓓�y�����9}� lr� ���e竜�9�_�S���x�?~��6^~�*��H��ൔ�C�W`�����x]���r���Qzz�)=x����9�b�˺��O�9�$������I����ܓ�ﻛ��?�E��ߝ��y��Ui��6$��5M��~�r����U��{��	����;{tW�9��%3�ZX�&os����ZVj�j��%!�b�dt|�aG&�toC�M
s�\�����E�G\�~"�6Gyb~�M�贙�H?�D0"D���8�t�$#���H=f:M~�9;$�O��|?C���@Eh*J�B��H��zW��$��
���"h�@�7��_�|�KK%�>H�#�7x� ��9��?e2�i�ݻj�e���.��UUU�T	��1�R�=^���̺F�0���R샓[V�;�U����X�;s�:����q�-�	�������9��qc���˘�L1	k`7��͇"DR �)��o���Ygz\y�zM8�
�ڴN�v�#�WhȲ�T�Yw/5�����`.��Vve�x76ø��V�70�C��'<r�:�tn���P��f��N��^�H��^:EvGS@l%��3�h��精Ε�6:7n�齌ny���B�,z�9ݹ�[��J��6�t�2����K��e�[�0�򼶭��)��dɭ(�b_��R��Jq�3�pnllN�Gbz��w�Q)x��N�
X��T�
��G�q�	�$,�/o�OA�����x�5Z
B�ճ��l�q*��4�e6�=�4<ON��շ/;�!B�Î���3�ݥ
Gq�7X���F�Q�O+�mH����wI��÷`N�I.���V8q�ٕ�݄��Քz�kHj-�zN4�e�'l�N���;�=Q#"���[q�F��ݦ��[@� ������ɞj\/dͮ�]�*�re]t�ݠ�FA8p��z� ��l��{!e�.%�ĺ�gI��<=
�����A�]��kﾾ�xqۤ^�C�s���N��n��m�\)ES��
0�˸Z�T�C�j�a̮:X�� lܜ�-$�ù��9��|G���d�]��۵3���r�uH�hˌ�m=���n�S�Z�θ!���W�|ݭ��n#v0f���ڒ2e<K�vE.���nT�ڛV86���#On����lV�r�uH����8	�*#�d���ϑN��%�۷.��P]\v�(+�oQ���\�e8Լ�d�I�w-���͹fF.H����6u�s��a�h�32�N��[v���]�u��m�yh0���%��"�;0��nY��j�ᝪ��,�0��+ !����]��gF�۲ѭ�V��	���V�s��,�A�D�ӱ�:$`�rZ�S5qG��I<LD�SȒ�O�&�_�?
'X���!ê�A��"= �*�����S������-R���f�&37��ć.3�P�C���&EsɞݷXz��]^�/%U�^!��-v��&!��-����͹n箸�!nn����bn-��Šk�-#:��(�/rY�f8g���6U�dh��U�q��ɀ{]����p�+����8�؛��$31-��L�v+��z$7W��Z�	+#��	D!6��ܨ��''�''$�'�}q$�rg�)β)�g�M����Vm��V��&%���jL��I'�o�IsYAV0�ց���>��w�N����r����x�K�
���4Sh�n��{5���Q3'�s��rN����ܓ�����E�+���ʕ[tLv��۞XT���W9�K�g� ��xwGWJZ]5wH����=\��߽��<�����/��+�^��,T��ޢ�j��Ev� ��/ �s������=�<������>�u�m��;�ms��ݮ3rgI�T��GJ���c����}�rH͐תI��髻J��	�� �{�܋�r�����퇿_�, ��W�m;t��֍h˗Y�'��]�ڢ|D��T�A*4��PXE���Ti"4R,� R!00�_s���߮�=/�Xݽ�y�RD�5�U������ـE�z�ˑa��%��~�O?���_=���i�J�3+����|�� �~�v�X�qK������vR�)�T[k �܎�W*G�/���׀v\� �s�)9(�[n�|U�d�)���a�5�3fש����^�É���w*Z~���Q��x�1��i�_%�,)����^�|���ְ�y�B^I�����m`M����������y`.��W=R�/W��������~�wٹ'~�n����n&��^s�]��^��kv僱�حYm��O�\���/�ܓ��f䝽�sr|xDw��T{�>\�gl�][��ژ�ʩrK��O^65�-POv��YHmy���:&�At����{c��,
�G�m]Mj;�'v���&p̒�����y{޼ �v<lj/W+��<�����
�en�� w瞽}%G����:���I/<�zK�V+��!�v���y`-�xz����xݞx]��*�۫4Zi����>���rO������N~��܏�	�k����%�@$�8���?߯��?}?�il?�F�S[����\��ܽ����~g�|�����=��̗]Ivm[[56�|�����փ�֜tYv��F���~OBk/����J�Zm�g�<ddXݽ�ܯ����%Oz���v05wWm�ddY�H����	�y����ԑ�Z�_�ӻj�ct����s� 6H��RGd��'��,�i:L.��JƛX�%=�< �x�Ȱ=�]��X�{�북S�E�;i��ݏ �r{�y|e�� 6H��]r�\+��9�p����/��l��c�7.-й��g+�]���r��l��LZQ�
Z�cg��ay��)T���M�����N����}����m��i�s���ӊ��i�н���-�
u�A"6��%�ar=�(��m�㮰��`yIm�"t�z��������qV��p\!�N�W�{�l��1c����Ї��V�%�x3�Bab�0����:º]0�aj�t�I�M��xD.E� kf����*����N��&��on{q�c����;�}}I�o^��a���F~X�r, �#���}`l�x(�*���j����� l��wc�6FE��W$�;-
�:9n[� ��� wv<=\�RS�g��=��%mYD��X�7E�x�s�Kd��'��,�^��\�S���;	��EҧN�M]ն��2,�ʪ��ʪ��~�} ��ߞ wv<��{�w��AԹ-�6��c��]t��D�U�%�a�Rm�*�-͋�};�t��o����NݷH����^ l��{��哾���䟽�z��tkD���k5��}{�����<� �@�( ��I�s�ܓ�䜿����/��9��/����4��aZ��������a��9\�%�=��"��xS���zġ����Ӟ�Ӝ�H���g��^���RK��+�����< �4��*�M�$:�cX��,T��{��#"�6IK,�cm��×V�!i�9L�0�;όz�&�[lv�"%?�<����ٛ�L9��]�������z ��=xwY��ʯ�v\��<�R�Y�C�T��� �v<�Us�*����?,W�~��{�Uč�W�|���M]Ҷ����>[%�u\xG9��(���KF)�Ad@��%����~y���=˸���"���M��۴6��Zk�\�]�{׀v_��wc��9ʥ�1y`�ؐ��&�v�N�ۼ� �\�W9\��ϠI��>Se���xn;������'3��BPǉ9�F�Zczۛ2,�w���ya+ P��)��w	�a3����w��X�l���9ϐ���
��$]N�W�6&����=\�q#��׀u{޼ ��y����Wꪪ���?��U��|Hv[�5~���>RK��������Fy`�ZD�r��	�V���9K�~��<�=x�,�hHGI�
<��oٹ'{���r�&�]:)]�XSe��Ȱ���>�%��9��'��l�k�GHB�nm���l:l� !LF���:�1hW�Q��Ng������ut��+w�=�3��"�^����s�_��t��|*3.Bm��M���W8��{�X6y��ȳ��U̟��I�SY���Ѣ�w!��~��ݏW9�%$g��_����+��WAi��Z�X���RO<H�,�r,�&V T��锸��m��dX�\�����;=�}������T+ >7��̽�)"D�U�qU%�Ԥ�j1�S��	�R�h͛���|�pµ�M�MX����TG��
�9�ZmzЗ�u�PC��*�[�1۔��A�� ^��{q��P��؃����&�ю�GYɛ��"�r�O&�H��Y���G#�b�I�W��[)g�eof��#1쓦R$�lKs]�U�֎I�D���#�K���Υ�{����p��^�=�A���x�J[-v�f��0�Dڭ!��œ`�,��^�Og|}cm�Wc��5�?~��`l�X����_ ��{�j�J��+�	���+=\�A$��W>A=�~XW���r�<�=CI��v�J�u�O<�����K������V�V����պ.���m�Ur�ɞK ���xvL�����r���~x�J?~c�݃�]�`)%��Uv{�W�O<�x�ހ��ϧ�^���hW[)kN��2pu�ۄ��Ge����P���=�w1u�$���m��w���V n�xwY�W9��{׀z����B��!�[��'�}�o����@��ABAXB*E*��	Z4!	���J)�0�!r�j�� �ƅ�l(��f).�LD]Bi�$ "Lq1p"�B��1 C� �0�X$f�Y!��D�G"V)�	�$����ܮs���3� ��~X�&Vz�UĂ���/·l)ڶ���X�r,?r���\�U���� �����H�e1��BN������ɕ�ݏ�ʪ��0��'�դ����gmڷx�&V��*����#<������'���q-�	-#)u�a#M�$�{8e=�g�$����%����7_����>����1R��|$��;�Ȱ���W�s��l7߿e`�z�`�uj�N�ݶ� ��"�>RK�>�2�ݙY��UU���s����£�r�o@y���@s��f�����7	���p��٘�A"D�p�M�Z�B"0��8h�A�R2]�q��1ؔ�7D)W�>��!:c�B!��/�7-��)��h�2,��b~ٟ��&�Y���A�Cu�t�>��ͬ�	$���|&��J�_�`jk��X�f��!��f�v@"E��#�	$�&� �q>HbB"H����ʻNhl�����I��5 2����~Bp�M�k��ɺQHI *��b	r!��WQRAB@C�O�	��"�!Br���S�y�@*p�!C4�iE#��}�L�0��e$�-?��N���o�2F��`X�`� �!�HF,��$aF\��Wc��"!p ���@�����4��@�D���!�vӐ�P�8�]	T�~���J����8�'�@�
� lA*tP��q�+\�?w����~ٸ�g��vP�Ɲ�Vۼs����}X��XwY��/ ��R�:W�mc�պ�;�2�s��a��'��{7?�-��{f�N���)˖y��ױ��Dӝ��;X���]��Yea�aI��Y�'Sh]���(�s?�)\����ul��l�^��~���l�� �?~�2�6]�۫�5�|�%�l�X{�+ ��"�$l�	yح�8+n��;=�vL�?UW꫹�3��"����j�l�Ң�v1R��`z�I�}X��,�Ix�3�p�ʪ*�#$��H�``����U9Wݏ��;Ҷ�4��m�;�n۬��� �so���g���n���$������%`ۦ��k�s��n�<�5S�9�;�Y3�.���j@�3狥�����5l�k�j����l�X�̯r�A�3� �OF!��6&��v� �d��7ve`�dX˲^{���Re:W�t�-�wn�I�}�Ȱ�r����xd�V T�]�K�v�����9K�a�u{޼�ٕ�� v�U��-�v"�-���^��d����� �u�`UU9EUf.rr�ӗ��#�[5���J�U�\�,�[�9�X��aւ��Oo���-��f�R��k&�4�N\�-Ǳ��D��ׁ��	��lT�X������3T�`�T���l�g-��5m��$�zD"���]��O+�e��nNWsu�a��Ea�˛r
��.c�\@Z�ۭ-1���p:����Eٶy]q�smS�:h[���5mw^aM�y��w��眳��Dݲm�98ӓw�8�����
oM�8��#�b:0��p��N^&��8q���O�V�v^��E�|���M���K��wI��ݺ�5we��H�<��O^�ٕ�zV�Z�-�'whm���q`)����\�Jl�V�^��$c�����X��,{�+ �ݗ��n�/� ��vЙnب�k ����=�ۓ���w�}�"�;��|un�e�ݖ���.�\��7hd���'I���䥰;/lM� �n��;�u�un��;��,������ �x(�j�t�ƞ�rO߻����	Հ",B � ��V(�k�����Us�'�~X��Vջ/ ;R\mr�7b-������X�Xo����Nz��6\-$��U�|J�-����W+�s����z�����UT��`l��V�զ��R��`�`�q,�܋ �ɕ�~���=�����b.摻���#�݇[p��Y�M���=2peT���&㺥��h�������r,�&V��Wh���l���;i`mȰ�Xw\0�eE���M	�v�䟾�vnI��ٸ�Li�@�p9�s��ʪ����b�7nE�E�+%�hwV�V� ����E�}�"�>�2��
6�R�]�X��0�,��ɕ�n�����g���%ݲj'���<j�+=gps�3���y�`��V�s�ZC���PWF�?`;ۑ`l�X�\0�,lui%����[���+ ������|���y`R��*��5lT�n��p�;�Ȱ�Ȱ�L��[�x��;bN��v���� �\� �d�����uU�����!���Tƛ;�>�"�>�2���XwY�m���ܰ)$Y�V�i�U�s@��/D�Vw �>�Fr�ױ�S���#)ڭ[-�5J�X�&V��ŀwu�z�\���vG� 򐻯P!�Iڡ�j�`m�Yꪪ����Xv?�&V{�Ă� =hU�wa��m�dg��u� �ɕ�}�ذ����t7Am��k�T��<`g��{��}$����}z�t�ߜY��.uٸ�fV��K����3� �^ŀO��"%?#(� ����(1H�ޚ̷,хְ�2�L��u����k hyb��4�d��2mBjaG&Ĺ�i�uH�s��5���W�^v�y�X���E1�l�v������^��3�g�a� W��»��3.�6X_�t$y��+�P�SA�ty9ɞѸ�HX��v�QWk8��,��v�]��s�t<�p����Y�M,��0X�1��
�̜�Ő{�8H�j�6���(�S���6�k�L�&]ɳ�QKp\�>����v��p�1�{�c8�E[J�wm*v�ց�'� �k"�>�"�7�2�鼗�T�wM��m����>RK�7ve`wc�7h�,v�MSi6;i`-���p�5n���ʪ��{<��������m�Um��7�� ջ/ �ީx�r�v{<`S��z��N��M�v�,�z��H�}��}J�����&up���M%��.�l]�#�L=�,n�W����8�q�v�:�ۍQQ���/ �G ��?r���	.y`���6��:|M�Zw�}��+��9UO��u����,�z���(:\�v
݊ـvG�wob�ܮr��Ke���;#�}�8���]����o �ob�;��^�܋�Iw�� ����6��'wnյ�nީxv�X����Ȱ���huuv�Yi�ƓK���ȣ�D���v�M�{^�r��pmj�Z��P\.��o}� }$xv�X�/ �م�ƪ�M�j����#�>�`�l��܋ �e]ԠCt��C�j��;�rnI��>�ny2�A�G{��������%*6Ъ;WGWm��R2z�ｕ�I�� v��V�.���M� ��� >�<��v͗�vIK,�cm�/�E$ݷ�c�ȹށ�Q[��Ϡ��ŷ"|~Hlq�#֝��g������X�/ ���ڥ�d.�;���x�8`�l�������q#t���6����ӻf%�׀w��W)#������ބ&[v�i���]���� }$x�`.T2�+���ʴ����ϵ�'߻���ɫ��i7IP� �lx�U�&x�QO<�0A�
U���U�!����8�ip!b���
k�ac>9��K�9����R���um[x�`Z�<�0�#�m*�4+V��`Z�<�0�#�7u�=\�q �����uwC���V��Oe`�G�ou� �ձ�G&��4�ۻu�I���Vǀ}$��>ڲ�����i4�4��7u� �ձ�I2��#�;UE_������n���"�)FR�b�L��Ja6r|��?r�~�狩f�4:��&
�O����M]Ɇc:"'��1	#$FA�ِ �Dv�e>?)��Ɩ�~��,T^3 ������M~0������'��@�(?����u��䚹3DUmnԻ-UUYP�Z����[��ٵh�g6���+.�éxX-�-����*�6�u���ϳ��렴�8�]��&0�^&��أ�91+8��aR�#K����H�]t���kl4�����cF���)��-�R�����`�;�������n;U�ey�W˥)�h$��=��w�h�\�+Hq'nC��jm�q����U�Ԥe�;��x6
1��7^p�*F�؞�c���6�Mv:^˨9wP]:�v�؇�h�����+��*��g;	������ zS����Sh0��m�	r�sڈ�ay����gsU�[��tR'l��˹4���C�g�-e��q�ܙ����mf����M��ώ��96z���́ۉ����OSVY��Д`��I�@4��D"7�c@r���)r�p뜑�+/ ��uї��F�%�s�6��� ��;rnF��I�0/�۵���d3��v��u���)��N�K�ښP%�k!�nI�-.��+q��!َ�1�ɭ�SC�K���t�=[c���y�9�l[��"nۂ�ȳ�]���CV�rZ�ָKm��D{rr�]�{t���k���AV��t�z��҅<��qlZܦ§K��:�8lu���\U�zh'����ib���������5�/8ļ�6rB.�a˕0���h�u:%8d݀1��݌p�Unܛ��bN�Z�gl��E���s�n7$:9O.<�oE���	��n�{%�6�3(�q�zАʥ,ѭ	l��1m5]�0��`�����&�`�B�ܹ���Sv��E�ljF	�0�ńf�Z�<!Vј%I�FbVY,��Zf
J�ћ��%��&,Kqٻ���Nn:�69�d"`�;vR"j��!�D�L0�u�EUT�p-F�N��[v�ѣf�U[Y�5]Fvvx����(���j��Ӵ�Ja͵A�r�]؎��$e&��*g�l�[s �rNNPt%��D� lWH���|
�b����G�C����b��@�9$�I';�)|��X9�F�ۣ�+��d�%s쐻'%�l�Z*YsYhK�tP�s��`!H�%�+M�S$V�vx�\�D�̆��\pN9�=r�r ��0T� ��6f��d,�����:9#�5raGNɬ�t�]Z�ݘt�Ǫ` #��5h��;�� �s��f����V�k��u��6љ��
�8w\ڐ����$�����!�����e�% ��b���j�u��Gt�opx�����^c�.�v�˫c�>�e`�#�r�U�	#�vQ��m�i���`զ���+ >����[{�č��$���ui�*J�`g���p�5j����XU���R|,��m��p�:�lxݓ+ >�< ��R[$��[���[��W�����\0�Ө���B
�H�u�3�M��`1VxqǅW������>,��ҹ:T�)���cI[xݓ+ >�<��s��|�TS� �����SI��ɬѹ$�{�oj�d �|WXm��� ��e`��ZR�[-���o �u� իc�>�2��#�;�x�e&1:hj�۶`[��ٕ�M� ���h����M�Hl-��}5� >�<{���� �()21]0v�@	[i�is�i:��7W#����ŵ�!ʇ��r{==j&䫫��h	� >ݏ �u� �ձ��I�;����נ<�ߍ�	m^�������W9UT���wny`�c�JU�*Hm�B�X][;{���k��]��	#� J�iFS��%CcV��lp��ǀN����R��<�	� �J����v�u��;&Vݏ ��+�<瘞�D���B�6�b�s��a�Uπzwbm��4�;([.��`Nn17�n��'d��6�v^7fV }6<�o�v�:l�������UW=��V w�� ���D&6�؛t`�m�vL� �H��*��� J�� ٰ����һt	n�=U\K����� �ݏ����Q��%��Z��ɀ�d���%'Pz�/�߷��䟩��wD-���:c��	������2�{�@}�����b���iYs0����n��s�#G����K1M+jdbR�4)�t��V��ק�;�+ >���g� ���)��IRl+o �ٕ��q ���q/l~0�'� �u(&�M�ڷX�����v��x�̬t��X�մ���N��Se��2�{#�;�qK2��M�Wvݳ �)��r�U���N��krN~���I��?���n������=X�V[��7ol�Y�se��sR��J��l�⳹�T��knxtw#<v{l�^'37[���^��6pp��N݇!v�<���p�(]�2�67���7�sTRu�5r��9��U���d�SR��hcv�=���SsL1��m�Gq��sw3��y7&lt]�g��*\1��3jz�-�/;N�6�9���Er��ӧ��z[=���%����ͺjS^ ��$]��4�rL���ۓ���b��΅]�V�\�w�M�+ 7�<�܋�U�����='�;,�tZ�$+u��~�H�߼�����;ݙY�ܻ<�W�͠J��T�'Lv���~XiM���n�L{#���eՔUZ������o �d��� ��"�"�$�uv4RmЭ��ɕ���܋ �.�x�l�Z��B���WuYX�b�ɥ8S��]��c���N�9�v]ˮ&7=�A�*Mݺ�w�x{r,��%�+����V�U�뢭/Rn���m��܋.��]�}��8USb��/ �ɕ��=\��䖟���}6���균<�}��;ݙX>RG{#�;�"�>�Lk��l��˗trrrr_<���@��<�܋ �.�x7c���	[�$+u��W9Ļ��,�W�,�ٕ�z�y�J���@Z�wB���`��C&]���u뜜�.N��s�8��r�����Nӫ�T�1�ݿy`v�E�w�2���x��JGM�U�U5m��}ڽ�=\�r�7g���<��r, �B�]�ub��+k �ve`���@17_d�T�.��ϳ޻�w�~��:�e!A�iq��M�u�wc�>�Ȱ�W�`�̬�R�R��[K�M��܋ ��{�ve`�����=��t�v��G�Q����p��kGX�kF��X�zf�Y`AfΠ�fun��ݦ��j�,�������v�,��"����LV��X�ٕ��]��ǀwny`v�E�MٔիIؐ���%n�����{�RK�>�̬T��t'v�����1�xݽ� �)%�w\0s��h��$�p��/�>� {�,�����1[��Ғ^ꪮ�� l���w�ހ��<��&͌�,.V�IKs^<=\s�Q|c�b�d��5<��8`׮�7�[�w�}�p�� ���`��^�[)
�M&ڶ�� wdxݽ� �-����+ ;8hD�햝��xݽ� �-���&V wdx{Z�Bƕ�V�j��m`z���z�ｕ����ʥ��׀wh��7whv�2�+�xݓ+ ;�<	�����'�>�u�'�O��U ģT���	�IOz_e�1�؅ҭR]j�9u�]��i�&�%����o#�Hcsl��b���{V��E���	Y9�'/ok�G;rFS�碁�	��u��] 06b�:��ѩ�e;=s��!m���|��ݥ�����9�9��kF!��W[лF"�b5@T�ck�Q��6�Ţ���1e��垭��&j�smFt�x�7	�4�ܺ՝6�)�VY���	���,66�c4P���t�/\!��Vp�S��D���p�kni,�3��v<��/ �-���̬el�(M�uj��
��5we�Jl��+ 6lx_@F�M�2ھ17n��6^�ٕ����/ %�+���n�M��ٕ����/ ������HU5N�mZv� 'v<Wv^ J�ǀ}$��%H�{L�6�l���M�X\�W�wK.�r]kn���67.�Ś���x-�M�j��e{)=x+���+ 'v<v�a�f�nɗt���]�~�C�!/�\�����d��#\��UY�'����ǀjݗ�l�Ex�Z�2�Wm�I2�wc�5n��";��vc-]����wN�.�`�ǀun��";��n̬jVʼBi���i[o �n��?r����<��{+ 'v<��s�W[xU�����<��݁}� �W��{��O$Q�은$�JZ��N�����6lsE��[~R��x۳+ 'v<�/ %�S��ҫV���wfV{��$������A�[=x���*󢆩�m�j�`�ǀwc��r�U�� U��!/�l���Hm�M3 4M��i�3`Kr@̜�%&8�4�%͆l��R�d���C
Z@�n(�0�!�JV��
�L���OΚ��yk�º�H��7�찜� k]��FX٣�R!��id���8$aY�r�`�R��&�F����B��,��Ya)I������D��L
��`!	��f�$���m��H�VX��� ���PF�rM�+(�0�HJ���0���
JKd��%�!d��^L��$��k$! ��D��B�	NB�Yd�bˡ����,&)p�!��������0T��(WYD��BD��aFB!FYBRR��Lڛ٣�|���p���D�T8���I"#(�S@� N��ҧ@SH"�âP8(��%Py�Kw��M�+ ;9A�]�-;�%m��K�<�	Kg� ��2���xݭD�,wt�5wN�x����>�̬�6^ }ݏ �!Wr�*i%m])�]a{vc�ϴ=!t6��\�59�cg�P��"s�Sf�x�\�����:�����c�6�v^7e�+�ݷj��`)���r�<�����^&̬jV�ƒi���wv��^ŀm.�M�X�l� ���G�v�M_;n��ݗ�I&V�/�(��C���� �!@	d"�F1"BX$s��o7$����F���ջ�7x�e`)�����y/�=�ߞ���*ٯ,Ԑ�uWvs ��=-	svr� �����b�?B�{�Ɩ�-5I��ZM��uzz����m.�l�X4��1i������x[%�K�/ �&V�/?W+�H��e;�`髱�k ��z�	�e`)��	�"�$�����M��Iۼl�X�l���X�{=x�}��Qv`�)3�;�{�����~���'� ݓ+ ߩ*9�|� ���p�(Z'����7 1�%,�`���w���Xu���2��G#��)��y�B2��@��v<�۶�������t�]�Cs���ڎr�Z��ɸs�+�F+��v���9Ĳ�Cb:#�止�l�A]��mC�8�9ۉ-��>ņcn�Tq�s ݥg�4���.��/C8������ M��������N�q�#7;��-��=.�\�3e��H)��C+ŨKs	Ǣ�4�2�R�i��K��z��r�9�G�o;kJ<�a�v/' ����IZ)�*�ݗmt�{�[���2�UU�|����=<�+wHw�Zm���e��e`mȰˑ`h�*�e��n�M��&V�܋r�\IW=��iI��>�TtS4ݫ���.��,�~��;Kv^7fV M**��Zn�;�![X�Ȱs��rz��{+ �nE�}ͬxz����6�K�A-�K��B���e��;�y�n\մg�t�`��m`��/ �ٕ�}�"�UU|��g� ����)�v���`�;w�N��ϟ�c*2Xc"iR4(H�`�����%�$j��D�,Z�4Gf,pF�"�h�#D��D�` 1"	�0 `) (��^��ܓ��/ �]�x�"ʻ��t;�	��>Se�vK�5��	�2��{:Kv"��M���rI'9~�{����x��|���
�
��Sn�����w�j;��k��/ �l��� !;v%t*
TK����rv��pb���m]�-�<��c�,�M)y�6�i��x��|���'c� ouG�|�����i�V6��ݗ�Ir, �� �\0�TUr�M];wuI[w�I{ ouG�����FE$B!�P5��Z�ܓ�������%�Չ��ĭ� �� �\0�v^%�X�T��ջ��m�	�o �\0s����_�{�<�{�<zh�)�e]��BT!5՚��F�%�΄BxM��0x�:՗��#���7vخ��� �we��� 7���7c�ޛNP��N��v��\� 7���$�˲^ l��G®�ul�ۼ ��$p�>]�����vDՍ�l�V�	��6��(����� �Ix�K�����2#[�Q#&1B��V�g(\H[By� �E
���7j�۬�{v^ wuG�N���NI���'�Q,3m��Ѓ@��u�/.ӎZ^�7p%gj۰p��S������T�m|��^ wuG�N�ʾb�e���,S��;�����'ve`�ǀEݗ��H�EGj�ҵw`+.��2������v�HG�w�^Yv���;�5J�� M��we��� ��+ �N	+e5E��
��"엀E!/ �0$���&�>�Q��]u�3/��+���Kf�4��X�L��rd��V5��țS@�	I��JMmL�mc�X4��7AP:�Q�=tv����%��WmB9;#A>y'���n3�m<���b�K�0�\ϴyb�'�b�"���*랧2Űut �V��.�@���+K�b\`r2���v�6k%���]-\������!u��pWm���U���=���p�g�	��+�����lu\��yoIrs�p�y�dv��p�p�:nӼ���N��V۾����	#� M��I/ ��n&��]��V���5�I&V n�xRK�>�*,���H�6!�X���M��}.TX�Xe��R��ݲں��oܮs������;��y`�e`�ǀw���K)�;hwv	��>�*,vL� ����e�����]?^�"�m��ǎ��i@�3���u�I�n�z�s���fX&Gj�[b�5ѽ���{+ �n��"ݗ�}��7b����Q�-���{���'s��+�X��e�E�Nɕ�v�k��Z|wE���[�-�x�{�Nɕ�un���*���[T�VۼUqv?z���z���X�)%�n���;t�ݶ�ۥ�E�^ݽ� �d��)`�9����Ӣ�ޗi�A���/�D;(۲�T��;��qۜ\\�aL�2�\�7@���QKr��{����'nE�}�%,.��j���E5l��P���'ob��%�s��<�z���x�4��m�ěX�gݗrN��w70x����٭��4E�����A�@���\�UUQʜ�����}/|�	�i6��J��RVŁ�Uq{_��Rz��ذ�� �vZ2�M;lwlj�l�:�e��o���˞��+ �~מ�c�!���V�F��l������q�n[�\q{\Xrn�Y��KƼA�eڷxe�Xۮ%�wve`�ذzR��UշT�V$�X��s��D��X��,�r,�W)#�E~���պj�۶�'���M�� �;&��t$��T4�6+M�6�,mȰ	�003�p�w�U��9s�`Т��*�­�(.��&܋ �� �0	��`��Ux����F� Y���	�����l2FX4 �d��lcz.��v�+sM�������I��M�+ �{�A�~��=(��6���8�,�� �ʯO{��K�Xۑ`�``얲�SI�Mۺj�[�m�Xۑa�R^�{ ������q�C`5i&�.��|�)Mr,n�l�X^�y`�J��N�PʰM��NɁ�M�+ �{�����6.��2��%3w1SE�:��� nHO���$
���NRBB�_�6�%5HkT6���/ ��'�MO���B�k|&������f�s���j�f�P00~~�ƂoF����4K:�Ϲ�-h��I��B�'�?b�as�5;��Mtp��A?_���:GiS�r��Q�0�q�*u�$�ߩ�����3��wȐ���Y��e:���h��HA�i����3D���A	��9�K�:�L�9�~�%x|�6E�	�/P�!��b˽��N��tr�r����m��[�U��Pj�����\�UWUJ�6m�O�2%��+�<�v[Rl�f�;5$�"�\]<��X4䎖��&�p�9� ��a�yFn݁���.t^i
N}�����r�8��c�mR����4�2�y�<�#8M�I�c���D��49��[�m0���;9��X�rV���)�y���k�<���걖,ug��[��e�˃=�����`�q�VЮK��
r:x.�b{|�g)��l�'�@�n�"����B�a�����΋b:0[j�ڃ{@�3���+��iR�nc�-�jj�4d�rb�$`]��Y����tx�b�;t��
W�mԔ�7B��&�ѻn&I�vvO'6�rc�;xjx!���+�q���\��g�We�h�d���,�8Y*B�¸0����Au��/\����YvR�2�V�)�*��8�^v���i^�q�v�n5�k�vQb�3�+�(eJ焹�듶�nثg����<8�X6x�D��м�x��q��n1��/1�@�t�mT^}��7kyxh�<������đ yt/�`y�ΚG��\A��� F�+�ݐ��O��R��;.��tvClN]v���Mǉ8V�g�u� �K��9h��q�q�'3���%Sx��z�!`���:�� ���㝳���UNq��(J�Yc\�M�Q6��T��7D��`)o�F�xpL�Tl�9��+�-��]×k\�ji�'n��.��"6䕡�X�dY��ڟ�W�jd��ݳ1��X�ʂ7���cn�v��#\Ɠ<��l���l��'�h�]u�9w�B8;��l"=��s7I^�<윙<sOI!�'q`� E���kF�<n��T�-F�L���]Ra����{\��:h�IX6��p�*ږ�Z�Lu��%UmEЎ�H43��N�9���N��.��z�nҜ�q5�:�l��(�m�g��t��L�C��������T��M
;��>��b�T�AX1�`*U ~_�Dp��U�SH�I?d��:U�[K�j2�G)��;5�h�6�I��'+V�L2J7s�L��4g�v�A�@\�#j^0aIt�ĺig1г�q��	�`]r�rcL�㍌���uv�*�4�C
h�6�!)� t��l�q����V�.|b*Fq���뢈���Q*]�!^�4�:�-+�Ʒqnt�mV��Bq�ZwJ쾴s:ru�s����R���{����u�v��72��ɨ�.^��L�/cT=�{g�ʬ�84��S=r�g�M0h�X�ذ	�"�'d��>�R�**�1ح7X�ذ	�"�'d��&ɕ�iE)H����V� �r,vL=�r�����)=xt�R�YI���WbM�vLn̬-�x
��\� �Fį,BCg-��&���=U�r�׳�����;� �W9��@���XU����ET.{\�$�<Y�v�¡8��cfZ�r�ڳj5���ٝ���߷@{�H�	ݘ�*�A�=��J���J�N�\��SY��ܓ��������!E��}3 �ve`we��IB��CJ�[m`�00	�2��e��"�"շUuwV��M�v� ��+ �v^;r,vL�֎�R�*-2��ݺ�&�ŀz�������{ ��+ ����-� EYwg-��L�v8tt����R��hi�B��|y�Վ����P]�����;&7fW��+��K�XaR��e�M�n�����``ve`n��>�"�&ѱ+�
�9h,�� �ٕ�;~���\�IB���%*Ĕ9TW
\�V�O��Xd�we�mF���6;3���NrN_w�����y`I00ݙX��ƕLV��]��}.E�}$��7ve`��o@~���g���k)��1o'�07vH�3�j�� R�;v�/3c��8Gf�j����}6X�̬v�/s���� �_�Uh�n��m�c�vL��9�RDRz���� �l2����J[�cbi��ݏ ��v,�vL� ��KU��J�Ҷ�ˑ`wI��nɕ�++�\��[��NY�N/����~'�Of5Z�7kj���2��2����ˑ`��l�c�m�ʏ9���=�zB�\s�ppʒ�M��B���Pc:����C����&V�ݗ�v\� ���+ ��E�6�&�5M[��ݗ��$o��X}+�X�X�)ƕLE�c�n�ˑ`v���7d��:���jU.�&6R㱶�����7d��5we��"�"�QZ�E�ut�J��vL���K���^�� �mL��FP]�V�)�����-sAq�2K�sn]�Dr�ʷ��ֱGe�j�EUzc<k�Ԅ"�dMfr�S��K��C]k;�8-K��\���Y��0�H6��D"S��=���H��f�uv�R�$2ϙ�W�µ�KR�:�<h��	�j��
�J�ǒ%�n:�N]ǔ��6YH�.M�!44ya ��P.�.q�޸Wl����p�D�Ñ�k@I�t�㻺v��/��\u�\3l��K�Sg�p��Ndv�otg�܊k�>C}���x	��wZr��t���RK�>�S+ �ٕ���
�`ڥwTZ�x�Ix�je`�2�]�y���*�;;�!m��.�w�w}啀n���yU\I-�x�Ix`i6�4݅]�:�� �ٕ��$ul��^�� ���+ ������c�ӻu�|�������[2�ݙX���*^�)x�x��q�s�:Y�nv����Ouɘ�i㝏	���y�)���x��:�v��^���ٕ�wve{�_��j��x�~�?	���+��֮��}ݛ����(P�R�P��T!!X�4�H
	(Z*X�`%a���c��\SZ��{�`jݗ�wnE�E���V��uui����ݓ+ �we����.���l�~��>�LJ>1q���7X˻/ �܋ ���+ �ɕ�o%B��&�+��ջ�:�K�=]�{��	=��/ �m��m��ui!qH-p��!񇥺��1��\&���C��^\ͭ-�I
�Bn�����7d��>[���%�����)��բ��vL��)#�O^����wI��v�GWiۦ���u�|�e�RK�ԯ�E.#D[
�	��"�P�Q��<E �������=���ܓ���ޥ5Jt��l�V��9���݇���̬�/ >�ۃcCT��m���2��̬�/ �^ŀ}	2�F�ܡ�A��Mu��A�=�n��'!�b��E<�qi a�o�t�;ǌM1������M���:�e�Kذ�J��>��I%ST�4+v� �ݗ����*���^�`v{Օ�w��}�6��'l�wTZ�x޹�v,��ٕ�uy绠;��6�\�Z��[V�rI9/���rO��nI������#� 	��r�Og���>������aV��X�ٕ�jݗ�}�ذ�"��;47�rreX��$.i��:��c��:�[���x�$[>��G�Y�Z��t�����O^�ob�>�ŕ��U���V��{��`��l�V� ���`wI��}ݙX�v^~�q �(m45K����;��V����>[����, �V�wN�'O�1����9K�{��:���m�X�����Հv�B�L��n�`-�x~�K��݇���fV UV�����/�ܻ�6��Z�B��V1�:B�j�l�J��W���������<�U�"N�b��T�{lPݵ7a3պLՄ�ɞԎ ܮ�D<�9^^�������kj�cpD��G.��r����Z�T�`ڤ��I�92� �V;g�����[3V��jifv���77vh�5�j�M��\f�pn�!nhѭM9��tkSB*�"�P4f�o�m�2����w�1�(P{YI]�f3w �ۍ��_T^y� �p���m��X۵2��fW�s���r�a���x����e&ӱ�����k �v�V����>[����,�Uʤ���۴��
�h�t�`g����=�����~�����V���p�6�h��wCn����{��L�wfV�^1U�����ݫw�}.E�z���^��I��/ ���˫�v�|�ڽ(kCl耱4i0�Ŕ� չ��f[�c��a��Z)��v[)q��X۵2�ݙX�v^�� vm˷t�݉�ݷ�f��>�����E�X� H`,X  B"�"��C���<��9{�ٹ'~���IϾ���}]����J�M	�u�|�e�K�`n̬��+ �w��&'i��uE�w�����W�U���o��+ �ve`-�x��w)���V��$��>ݙXwfV�ݗ�}�"�?Ur�+����$��2�7S�;s��>��GMv��2���<p{�f�3w�\{�p����eg@�߲�{��v�X�fV���p�m�]]��n�{��v�X�fV����RD���J��`�][E�xv��}6ea��E%ErVg):*�)?wxՙP�#�	��v'#����M��Y��f�c)'���$a霍>>��mБ$�>��o#Ѕ�#4~yvȤ� |�
Q%H��Jh?3!u�Z̙&a)E&�X|���� R�/�W�ὓ��2���t?k��s�)(�q�֎��I�!h��>'ߙ��ٶ��$�پB�1�9����P����t�!|M/��%��tC��%�H�$C�c��e&�(U�I)���T�vp�I����&u�!�a��������u_�� � �����0Z��ӿ����? @��>�5U�~E j��G����7$���������t�l�R���X}=��w�2�{��v�X�ۊ�ӫ�ݔ�m�u�w�2�{��v�X�fV+����F��-�^t 3�fe�q���yU��2{\�f��ú�������&�>�g��ob�>�X�� ޕQ1�MU���[xݽ� ��e`�2����Ԕ�Si�N�U�I��}�2�	6e`{��^ş�UI��.�t�N�)���q{��Հ�� ��X
�����+��9�c�;X�e'&��ui�hm����	.E�}6e`G���Z�#��
���]B�fh�f���Ȑ&-���x�Gn�:�����ui�I'm������	#��d��$���x%-Q�
m���v[f�d��r�\�q"{�� n�<dp�s�U�$%�7t�X�T6�M��~0{���� �l��>�����-S)�+�x�����}6e`�K��*&4骷uV+o ��W*����	=��u�aRET>��Kۆ��K��[�]+����0����]�2�<:c�c���p������2�c��i�so[L��,&c�ۅ�!ƟF���8�x��;ux�N���@L�"���rx�:�n�6Jt"�#�a�4q����ZekmF\K+V�%�[>oozڞ�� '�a�;h9�ç=�k'q��)t���a���3��a�0v��L��/I;�MӤ4��,5�vrv�p�]�����A�c����8���������6��<�7Mf�վ���tݑ�wc�;�"��T�n��
c����`vG�ݏ ���+ �wiL�M��黫V�o ��ݎ�fV wv<d���I;QwI�[0?W9T�=�0�<����w\0=\��%4Q_���塶��<���x����*�hB�k	���s/+	v1��fX�7�C&��	��m��0�\�͐t�W�>�ذ���&W�U\�s�vy��J|�]ݡ�hv�0���Ôp��+��UϪ���p��ǀn���Di�MU��l�>�e`����p�>�`]�w8Uۤ�ժ�N۬ �������&V�jrպWt�m �������&V }ݏ �])pR���I�m��am���7e�6/��`;��0-��#��tծ���������̬ �����*,t�N�e"�;� �veg��y����;���A�/]�����˻V� ;'�s�ٹ����DX�߹�rnI�������o\�̰t����rrK�L�vG� �ve`۱�T�E+�we�9n�m� �u� �ve`�#�>�p�=U�ݕ�:V�.!]i������ȝ;���[��v�%B��i4���@���ժ�uE
��6{�V }�<����{*cTUۻLuj��m� }�<�I���6G� �veg�#|D�wn�n����;o ����=UĻ'���y���-A�ح��6�����3��=��wc��W1]����}��}ߎ�趧c*�݊ـ}�2���x�{�u� ���]_���pv���*�#�Yҁv��i��nw<��a^-�j�U�|b��v� >�ǀ}��`w\0�̬�l�v�V��vӶ���� ���ou� >�ǀ}KM�]�v*g-�ݶ����\0�)#�<��� mt��6:�V[0�`�����X]ٞ0�/e��V��uj��v� �v<� �~�f���vnI��p:��R�B�s�f���[˶�6��yz璸+�lαڤ�<�3�+u����p77	\��m� �W0��b��V�<�s��r���ع��%#c�!	ee��s����Z�f�������3�]�	��u�n.��%��x7�yv"�6�3*90;_��[�+nԎ��0�F ����s:5����v�ٰ��-��q]Mq�6�R�-��l���N�����Q���ԄФ4��.q���՝:�|��a#��':l�b`�Y7Uo�j���?W;&x���{��W��y�[�Cbn���w�wu�=\�RGd~0��x�v^}�RF���J��+Uun�l�>�p��G�|�e��p��
K�B>1S-[f }�<�/ �����64��[���T�o �n��;��ou� >��bN�[�uir�K�L�\�gv��V�Y�F��	p`ho�������J؅L�m��l���� �dx6G�WH�.4�Um�,�ܓ�w�7ÀrH~� �s��[�N�c�;�៩"H���E����	�X��< �#�;��M�+ ��N�vZ�ucm�N��	�<���2�=T�g�����N��Z��6���l�X���l� �I�o8��[x)uPMB*�@��Z1�ka+y��)r:XB�K^)`&�0R�d��*�V����e`�G�dr�A$b�˽+-kH�!�g@y�@7�� ��lp�:�c*�7t;���� M����UUU�S8�
B�b��� �.�� ��R�����\�awm�m#u� �0�#��W����Z�YV�۴�۪l�;#���9���?�$����y�V�;W��7���r�u�6��ӻX��8�]�n��/�Ӑ+�V�طZ��mrtߞ��ݑ��p�;�� ��N�v]+wm6����#�;��wc� }$y�URFȝN��M��hm6�	#�n�.�x�#�;�Rƒ�e5Ɗ��l�ڥ�L�.�xV�x<ܮWj����� O�'bM���L�v� ��^ղ^7\0�XГ($�-
��L8�P�מ�2��^���&��g�6��9�s�V���v���:�K�&�ݎ�W>A����[G�y�v�9m�]��&�z��$��yo�xT��	��K�Rݶ�[u@���p�"엀vGn�`MN��c�i�I	�0�%��� ���p�>�����m�7i$���0	��n�.�xʧ��o�u\Vs�e�>59��a�ӌIb����5XnG��| g�Ä�����=�U��)w�X��c�4Jf�'u�a*��ztt��a6�N#"��~��>3L�a���_��{^�3L�8�f�4!R/9�gđ�.������^���!�4:�S8�Ėz��.�V�9u��?�V-`�_��7��<~�5���O����B~��.��p���F�%�I�ĥ��֓tk鼅��'��>�/JX�C���x��;�����'u��t��
�! >�Hq?
@ A���,خ�3���ͦ���㮑$����?y�F�)I�Q����ĸs�l�r�c�����|jF��&��@����s�wy�x���:0��2�o.���-]h!�3�H�nhOvw���}=Ӂu8�!"� l ��+���d!��$4ith�b�Ȥ$���\� B���+"��#�kc�e���kq�O��w��P�R�d����"�2|s�Һ���~T��t	��*����D��N�4I����B~ةN�B$���;�����2�Wmv�9Uj�vf
����.���H��5��I\��&k(��v�;<�^�y�#tM��.z�N��m�"��
��-0n�0�/��ύ� ��^�/�-�,q��4[��DDh�j��CId��W!]s�[���qj�L�l�6��	N�ĥ<�[k�n��=%�'�EV�"���Md��x]�׉<
7]�6�7ӣ�p�!�h�إ ��J�RE�%��-,�Ea��ڒ�g�|��̎���4`�M���vB��� ;ye[2Kywl�ś������x�����m�&����'0�0� υ͑S׌�MΘ�v�V��a���<_c���B�#Bm����"�`:'���%l�������j��z�8�/m�V͍	Wl���Lu��)���k��⬻���!8�7{l�Y��nɀ�g��ܽ7gr��v8^�Xy:����s�A�Z�&�6�q��0�5]98��kr�Y��\�	������u���,Q�&+
��`!ñ��h�ֱ�ʬ�ݡ����4��یJ��/Qj�Puև����Y�l&�:܌��z�@4IY�)a )����O]���P�
�hŃ�è���-{!��fy��
m�*��v�n3�5L93���H�]�Vib���l$�7&89§B��L�Z��VL�`��J���)TE�%LHkA��fs�68ͣ4J+56�ս;�8�qΐe�S).a�J�N�چ��T���ӥ�5XƗ�,�8�lvŖ���g7*���ķ!�=�&���Ӄ��T���V�����'˻=�����r�u��7�qu�LX�d�N1��B�CTq<��cm����:�����g� ��m�&�c�j��Ln���v؅g�q�2H�c�����s���ڛ����G;��/m�^�hUVUV�W\D�W+�����8.`)�AԲ�:^��N�n��q���-ǻW)�Љ!0�:�j8�d�7s�cb�xCd��f���nh8�b*�D�Ȋ�?  ����"��,�p�@�b.�@��|�{�?\̙�,X�������R۪�f���������ɡ�vEL���$��f獣�뙃�:���m�������cRi�g��"���.�gYZ�܍�,!ɤ�H�bD䣪�j�6.7��ɷc��eZ��m2��I���2y�;>T�ۘm�gۥ��^&66ѧ�b���fy:F,M�gl���ڹ�l�z���x%�˃ �k��Np���:��&v�r� >b�ڟ��Լn:hy|���x�'�C��Z����f6X�*���?�� ��^68`�)cIU���m�ـM�]��	�� ��ڛj'bV��.�]۬.�x���#�{��V�6SJ�wI6�n�ۼH�M� �c�"엀v�mhAշVU��jـM� ٱ�vK�6k�)o6!��(L8U��@��MrJ^�n���6��e�*�j:��2�'@{�@{{%�/b�&����Qjۦ��B�kZ�䝿���}~�p����#�tq�*A?��L)��o=�w8ؖ'}��M�"X�%���}�ND�Qʙ�����gY���љ��sY��Kı=��]�"X�%���~�ND�,K���6��bX�'��{u���NJrS��O���p���f ք�j�?D�,K�����r%�bX��wٴ�Kı=�{ٴ�K��	�?�����Kı;�O��a�5�q�j\��r%�bX��wٴ�Kı=�{ٴ�Kı=�w�iȖ%�b{�ߦӑ,K���OrJas,�\l	e�J�SF]X1wi�a��&�N]#nx��<�fvr�CFa�nr��}^��^�'��{6��bX�'����9ı,Ow�����2%�b_��kiȖrS����￣�Z�V�e�rvrQ,K��}v���"G"dK�����r%�bX������r%�bX�Ͻ��r'���2%��<O���jd,֦ff�ӑ,K�����6��bX�%��m9��0���Xn&�{9�ٴ�Kı?{]��r%�bX����S�QJe�.N�;9)�NJr_~���Kı=�{ٴ�K�XdL���{��9ı,N�{�iȖ%�b~�ޮ�We��[�\����%9;�{ٴ�Kİ��{]��r%�bX��w��Kı/��kiȖ%�NO���Sv7r��Y\\ٙm�rY���ܝ^�Xʸ�뜝��q��s�������zA�e��m9ı,O{]��r%�bX��w��Kı/�����Kı/�����Kı;�n���k2h�&�2٬��r%�bX��w��Kı/�����Kı/�����Kı;�{�iȖ%�b}����SF�U��]j\��r%�bX��{��r%�bX��{��r%�bX�w^��r%�bX��w��Kı/�w/�2�5����n�kZ�r%�g�"g�}���"X�%��k��iȖ%�b{���iȖ%����!	|� eR�AJ$t�B('蟻��kiȖ%�b_w���c�V�y\�rvrS�������]�"X�%�﻿M�"X�%�w��ӑ,Kľ���ӑ,Kľ��12�+�<�fYU�������]�q�r�1�*fhrr�A��
��OqȖ%�b~�w��Kı/����r%�bX��{��r%�bX�w]��;9)�NJr}�K>�Y���y��ND�,K�ｭ�!� G"dK�����r%�bX����v��bX�'���6��bX�'���g��u���K��m9ı,K߽�m9ı,N�]��r%�bX�{���r%�bX����m9ı,O�=�楹����.e�f�m9ı,N�]��r%�bX�{���r%�bX����m9ı,N���m9ı,N����5s.jI��iu�]�"X�%���~�ND�,K�ｭ�"X�%����ͧ"X�%��u�]�"X�%��� O�Z�`�{�����L���umu�]���;1� (va�dWu��ҹ�A'�r��1+cyy(�7<��v�'��{����lE��h���7�6������{3*L�cpnVv:�i���m��h�Gi�j��	�\��\��v��[ �;s��ƒ�MӪU�&��ja�Fp��x·��䞪;$Sԛ�y�v3�8�])�ڦ.�WWQ�'O��ݺt�
�H�P��~�\��궙2t�]��&w�q
3=#�e�=�ce�t�94ɣ���-3}��z�z������r%�bX�Ͻ��r%�bX����Kı=���iȖ%�b_�ܿ[��]��������NJrS���m�!�$r&D�=�{��9ı,O���iȖ%�b_�����O�r�D��>}��1�:���s����/B�*{����r%�bX�����r%�bX����m9ı,Og��m9ı,俧�`���&%j��N�JrS��﻿M�"X�%����ͧ"X�%����ͧ"X��!2'����KNJry1�?����[��Cd듳��,K����ND�,K����ND�,K�k��ND�,K���6��c)�NO'���;Y]v��a�a]�%CT�K�e�R4����:^I�n�X{;��d-h�f�Zff���Kı=�{ٴ�Kı>����Kı=���iȖ%�b^��kiȖ%�b}���֭�5�5r�ۚͧ"X�%����]�"&�"��D��&�X�{{��r%�bX�������bX�'s�{6��bX�'�=6�f4I�-�Z��r%�bX�{���r%�bX��{��r%����=���ͧ"X�%���{�����'����^�crm9ı,K��m9ı,N���m9ı,Ow]��r%�bX�{��듳����%��v�����,uWiȖ%�b_�����Kİ�T�{~��O�,K�ｿ��Kı/�����Kı;��YO]9tL�Ʒ9m���z�]���)۬]n[W''v'q��u�1�9�˚+*�\����%9>�]��r%�bX�{���r%�bX�Ͻ��r%�bX��{��r'�eL�c�~�kC��I��=���/B�/����ӑ,K��}�fӑ,KĽ���ӑ,K��u�]�"X�%��yϹ�nKv����'g%9)�NK��m9ı,K������c���*M|24��`&ƪh
<�Ț�z�9ı,N����rrS������z�������l�;�bX�%��{[ND�,K��}v��bX�'{��m9İ?�fD���ot��н������Ɇ�\Lֶ��bX�'����9ı,N����r%�bX�Ͻ��r%�bX����m9ı,O����e�p�u�d�e2�^[:lH��i"nUcQ�&1:v�cXJnf�l��[�'g%9)�NO}��6��bX�'��{6��bX�%��{[�V~��,K�����r%�c)������;4f\A���'g%9(�'��{6���1șĿkiȖ%�b{^��ND�,K���6��NJrS���}n�(\זmU듳�ı,K������bX�'����9ı,N����r%�bX��{��r%9)�NK>����Ζ̢������bY��"{~��ND�,K����ӑ,Kľ�}��"X���x��,�%�p�O��� T�N���kiȖ%�b_��%��u�d�[n����Kı;���iȖ%�b_{��ӑ,KĿ��kiȖ%�b{��ӑ,K���7|��kY	Hp�˛�w<gwl��Y�Z�#���Mt�B�7��(z����3�)n�0�;��rS���K����m9ı,K������bX�%���m9ı,N����r%�bY��ϩѾ��Ye������%9,K������bX�%���m9ı,N����r%�bX�����O�2�N�������"5�%�Ze�O�н�%�������bX�'{��m9ı,O{]��r%�bX����m9ħ%9=�~�o��fX)jez���%�bw�ߦӑ,K����]�"X�%�{��ӑ,K�DfD�����iȖ%�bw�?���9��$�K��ND�,K��}v��bX��s����m?D�,K��^��ND�,K���6��bX�%CO$��:-S���Xȩ&w��&f�%2[f�[<5S�TJ��\T-u��{v��ԉ��������V�8��u�u�����.a�����˝�A��ֶ��y���Kw]��nv�+8�t�.�
���c4������S=v�4t�pqKA#ϵbb����mm�T��hFG��A���ls���u\r]s�gJ�����9#�J�\��
Y�2��E�/[��*�>���V����$䑝�	gF��Wk:�V>wm#�p�q�1���r�.�<q�b�i�m�354��Y��Kı/���m9ı,O{��ӑ,K��{�M���L�bX������r%�bX�a����V��\����%9>�߻듳��bX��w��Kı=�w�iȖ%�b_�����Kı/��K��jf�Knf���bX�'{��m9ı,N�]��r%�bX����m9ı,O��siȖ%�b}�=|f�kS.e4L�M�"X�%��u�]�"X�%�{��ӑ,K����6��bX�'{��m9ı,Ozv�S��ֵ3Z!l��]�"X�%�{��ӑ,K����6��bX�'{��m9ı,O��z�9ı,H�ǎ˻쐍�Iv�����Tѱf�л�s����w����l
Ն�K^.�a���m�"}�{I�$�}���ؒ! ����n'�X�%��{[ND�,K����=�L�պ�,�5��Kı;���i�~A��Q@�Ȝ�bwz���Kı/�����Kı>�{پN�JrS���y>��v,��E.N��,K��u�]�"X�%�{��ӑ,K��=�fӑ,K��{�M�vrS������~���ݲ�˜ݧ"X�%�{��ӑ,K��;�fӑ,K��{�M�"X��"w�\����%9<���O�e��Z��kZ�r%�bX�w^��r%�bXG��?���Kı/}����"X�%�{��ӑ,K���[6x��\�!&BR�cX:ks�& H�n3M ��v��Lvvߔ��i6�Q3q`�����%9)��{�iȖ%�b_��kiȖ%�b_����� '�ı>�fӑ,K:�ϟ=�s�˱�2��t��Щb_��ki�b���,K������bX�'�｛ND�,K���6��y�5��%9?x}a���T�,�7.ӑ,KĿ{��ӑ,K�����iȖ4���E�g��\���̲���3!���$Y���I�����6gM�,�nB`J˨�.7ń2�Db�ʁ����u���%!��LSD᝸@����@݉��D���&���I��'����r��t���N`h FBJbwQk� ���d��2$V�H����O�5�d��w��.o�ی!&�,~���Ă�c�m��JF@�$b�5.l�j!���a	BV0���C�6�^]�!��_��qO�3IF��!$�{$��]�oxDM��~� H�)�)�0ޛ�Yݙ��2�1��Y ���al��	X4�*���PԻ��ā"m0��M+������_��ß)���9�
f��Sx(oJ@-�p#6��'u �Bu6M�E�mGH5����B0 �4%�hPAM�L�(0^�QWC��DC pA�u4���S�&� N����t����ND�w�M���L�bX�������bX�'N����fa��йz���%?�9�Lry�����r%�bX����6��bX�'��m9İ?��3����m9ĳ������
Wir�u���NK��{�M�"X�%��{�ND�,K�����"X�%��;�fӑ,JrS����/��`������cH�^:se{]����g[y04�e&�!e�VKK4�C6fb�nԹ���Kı>�}�iȖ%�b}�{ٴ�Kı?g}��(�"X�'{����Kı?�{���k4[u0�e�ND�,K���ͧ"X�%���ߦӑ,K���o�iȖ%�b}���ӑ,K������ˍj���w\����%9?z���r%�bX�}��m9ı,O��p�r%�bX�g��m9ı,K���|.��m��rvrS�����Ϻ��9ı,O��p��dK��w��6��bX�~� �jB�����0 �A�"w?]�"X�%��k���sY�kY�!�\��r%�bX�w���Kı>Ͻ��r%�bX����m9ı,O���6��bX�'������f��4^���XRXŦ�Z�]�6,��ce۞��ryr椱{0��vY���z�z����iȖ%�b~��ٴ�Kı>����"�?DȖ%��{��ӑ,�%9=����l�i���;�N�Kı?g}��r±ș����6��bX�'}��ND�,K���ͧ""�eL�b{�h����ˣ2�kY��m9ı,N���iȖ%�b}�}�iȖ%�b}�wٴ�Kı?g��m9ı,O���s��5%5&a�K��ND�,K��ND�,K�ｭ�"X�%��>��iȖ%�b}���iȖ%�b_��C�P֦�n�ə�iȖ%�b_�����Kı?g��m9ı,O���m9ı,O��m9ı,JhI?{ڒf �������=]R�o3d�9�y��ػ�O-�p<�s�r�BA�Bq=���nݕ��&��L%6�a�1v�:x�Ҝ\�����ckTb�l�9����3�-q���@��R"�=îZ�YJ�uo5j��U��$���=nr�@@(�|�
	�;b��8EmX�"WY�c�B�	�t�;aZ�Wt����s��7�j��\'��@!�"��7���c#����Y#�����^�;YI_��%��P����p�@�U����u�bX�Ͽ��iȖ%�b}���iȖ%�b}�}�iȖ%�b_�����JrS����<�=����e]�'g%�bX�w���r%�bX��}�iȖ%�b_�����Kı?g���r'��9$ד������2�i�k���m9ı,O{��6��bX�%�}�m9ı,K�w��r%�bX�{���'g%9)�NO��Yo_$U�e��)��Kı/{�kiȖ%�b_{��ӑ,K�����"X�%��wܝrvrS���俧�o�\�1�ڔ�Z�r%�bX��ﵴ�Kı>��iȖ%�b{���iȖ%�b_��kiȖ%�b_t�&e���3,�h�a�+e�n�擜��^�v+
���dnD��ppM�PJ,&K��U듳����'���m9ı,O}��m9ı,K�}�m9ı,K��m9ı,N��ԸrCZ��35��Ѵ�Kı=�w��>t�	� �� ! �� 'Mb@ND�K�~���"X�%�}�}��"X�%��}�ND�,K����]CZ�%��)e֧�Kı/}����"X�%�}�kiȖ%�b}�{�ӑ,� dL��}���Kı;�����5��֭3WZֵ��Kı/��m9ı,O��p�r%�bX�}��m9ı,K�}�m9ı,O��=g����Y5��ֶ��bX�'���m9ı,O���6��bX�%������bX�%�����"X�%����ן]Y��6�Q��<�e]@n�ni��l���M��
��YU�H�7Eu����?,K��}���Kı/�����Kı/��m9ı,O��p�r%�bX��씗w<��kE-��jm9ı,K�}�m9ı,K��{[ND�,K���6��bX�'�w~�NF{�5��%9/�߷l.�h۩�wIȖ%�b_�{��r%�bX�{���K��bHT6'��J(�7�;�o�m9ı,Og���N�JrS����0���:�i��Ñ,K?@ȟ{���Kı>����r%�bX���ٴ�Kı/��m9ı,O}�ԸrCZ��Y5�u�iȖ%�b}�w��Kı;���iȖ%�b_�{��r%�bX�{���Kı>粒5p�u�k	ne�e��	�k�e���7 .jRֺ��Z8y�14�XŢcM�T듳����'����iȖ%�b_�{��r%�bX�{���Kı>����r%�bX�g����-�9�s�듳����%���kiȖ%�b}�{�ӑ,K�����iȖ%�bw�ߦӑ,K��!=�|#�h-r����NJrS�Ͼ��iȖ%�b}�w��Kı>����Kı/��m9ı,N����è�n#3�N�JrS���y�_M�"X�%����]�"X�%�}�kiȖ%���a,�!!�$����T�Ț��iȖ%�b~��JS~�K����Y���Kı>����Kİ�H�������Kı=���ND�,K﻿M�"X�%������f~��L�2�{Mێv}�g�6��WN����!۸=ɠ� ��tv[MZf:!�e>�~�B�/B�~������bX�'~��m9ı,O���6���2%�bw�^��ND�,�%��������j���'g%9,K�{�6��bX�'�w~�ND�,K�k��ND�,K����ӑ?�f���'��[;�K8�:��Kı;�o�m9ı,O����9ı,K��{[ND�,K�{�6����%9/���|��mM�T등,K?�H�����r%�bX���kiȖ%�bw�{�ӑ,K�����N�JrS���o���e����[��ӑ,KĿ�����Kı;���iȖ%�b}�w��Kı>����Kı1�Z6bH�B@� �{v��kJ�2ك%̲�=�e�����`ܶ�o^�0�	�l�M)���a~F�ȘC���8Lq�s����p�Y���ո{{^F��yGv�"6���-��/`J�[�7%����ks*9�aWCL��`P[�n2#R�q���ꂛ��f�K�ڝ��cmn���n�r/f��+S�E��6�
0<rU����J�;t�&[Ψ����jM�rs�&�kZ0��ݠ�W�-��!/b�7���m�(ݠU=qCs�Ķ&�L�Z��Ӓ���{���6��bX�'�w~�ND�,K�k��ND�,K����ӑ,K�O|}��L��ۈ��듳����}�w��Kı>����Kı/��m9ı,N��p�r%�bY���HP:�ڬ%�9:���%9,O����9ı,K��{[ND�,K�{�6��bX�'�w~�ND�,Jr~�}��,ͫu�-듳����/��m9ı,N��p�r%�bX�}��m9ı,O����9ı)�{,>/�3f�aCe듳����bw�{�ӑ,K�����iȖ%�b}�w�iȖ%�b_�{��r%�c����Kgͱ�CR�P.\�#:6�E��Q])9�e��yۢr�rJ����t[)���u���%�bX���6��bX�'��}v��bX�%�����"X�%�߽�ND�,K��{XMM5��2Lm֦ӑ,K����Ӑ��A���;��R�r�`� (Z��"j%�{��kiȖ%�b{����Kı>�޾:���%9)����>6c2�TV�j�9ı,K��{[ND�,K�{�6��bX�'�w~�ND�,K�~�rvrS����p����c���Y�m9ı,N��p�r%�bX�}��m9ı,O����9ı,K�Ͼz���%9)��3��qk4m9ı,O���6��bX�'��}v��bX�%�����"X�%�߽�ND�,K�|{�����h�e̒�+�쌹ƛ�VŔ��$S�x�ɻ��67Ds����B�46�aJg'|��JrS������v��bX�%������bX�'~��m9ı,N����r%�bS����B�*�u�-듳����/�ﵴ�Kı;���iȖ%�bw�o�iȖ%�b}�w�iȖ%�NK��a��0�5ڵ�e듳����bw�{�ӑ,K���ߦӑ,
U� ������N���6��bX�%������bX�'�w�ɇ$ɪCS��Z6��bX�'~��6��bX�'���m9ı,K���m9ı,O}�p�r%�bX���ڤɅֵ��SM���r%�bX��w��Kı/�ﵴ�Kı=���iȖ%�bw�o�iȖ%�b 8w�}?��:a�"��C����&�ʩtچ�aRq�6���uͦ"�4�~�bX�'�����r%�bX�����Kı>����r%�bX��w�N�JrS������|�* "�m9ı,O}�p�rș�ϻ�M�"X�%���~�ND�,K�}�ۮN�JrS���x�>˕�Z���6��bX�'�w~�ND�,K���6��c�C"dO�^�m9ı,O}�p�r%�bX�vI�ONY3���SiȖ%�b{��ӑ,K���{ٴ�Kı=���iȖ%�@�|�����ʕCB�[�L �U��Lj�H�`XU���(�⡨��?rm9ı,O���&�c�֥ɫr�sSiȖ%�b~Ͻ��r%�bX��ͧ"X�%���ߦӑ,K����]�"X�%���ק����v �i��ٲs0��̘��k�À�<�;��$D�(��j�ӕd�Y��~�bX�'����6��bX�'��p�r%�bX�����Kı/����p�%9)��ϭ4�դm�q��Nı,K���6��bX�'��z�9ı,K���[ND�,K�����e9)�NK��!�L��˳:���bX�'���m9ı,K������bX�'��siȖ%�b}���ӑ)�NJry��O��ʷ9�\��N�K����3�kiȖ%�bsiȖ%�b}���ӑ,K��w�ι;9)�NJr_�=!��j�h\�zND�,K�����Kİ�+^��ߍ� �'�����A'>�u�$D� _�� _��
��
�
�T U�PU��@W��
�����* �H��D*��b(��X* �"�0H� �"("� �"�1"( �� �H� �"( ���F"�1"�?�* *��� *�� ��PU��
�@W� _�T U�PU��@W�� _� U
 *������)��NNoo-��8,�󞳮����0e����[fM$�l��
���@8� �  �R @%H��TR( RI
*�* �$ �"�  ʠ 6
�S�F�6�r[}�+E��|�;���7}�� �       m����������00Wz��@(w��@
PU�{�������
t4�A����:0�����{��܍�'a����V�l;w>�}T P}ܡ�0�f�p�ۮg��b�*�7N .��p�(�yu֭��{������v��|���  �<u������}�|�}4E�;����O�|>��}�L�3Y{���v6�w���=|4�@
 l�V�r�6�m�pW�w{��޳��YcM�ݳ�_O�|��:Ֆ47�>��������o�C    ɒ4ڤ�(      Ɋe?U*J�      OǪ��i M    تTOI%       �� jR�i�� �L 	��!HA$��2��I�OJoRm��i��ԟ�_��>��~��'�O�
{/�����Pqo������DD�@U �P�?�����G!���"*�� 
�B��QP
���/k��"*���2_���R�����j/���4�դx���*(�Pc��Y�����z��&\# �`Y�0�PV����b��j������0���~ֲ!�� 
D.�F͔6&�݁4D�#z��2��voy�3�N�6�<8Gk��ƍ��^��[���$���hc��we�y'26���ț�S9"���ֵ�Ӵ�hZ�14h�-!�ދ���A�r�@��v�� ��*�Z$LAw�wT�-Ks�Qq!;kS�iZ�E�M�=���V'7�dU@dh��^o�DKNEJZ���oHzH��-_�k���"����ֵ�tFOx���LQ��,bbf���u���f0�.�z�T&պ"ǤU	(�D����
�+MK��&�JV��#R�l�|8.�M�����ō�F'�%�f��?8�㓄���=��i
7q�he��V�hߩ1!:��i�J�����T-�J�!��bh��!���YsVk}p��{\Z��Bii�;�q9��(�����F�QB+CM=�Q�oʅ�D��A,������h,���e�fl��s#�<�kn�7�b։C�Bj�ӋI+Z����-i���w9�.ǣB�t&q�H�n�.��{��9��3Zh�Жa�e�sf��t'Hi!���!9-h����ޕ�3�;�0�u�a8h�7��%��/P`L��gx��<wtM^��ND����N��j�)�ЊEa�-�V�H�+9�Q��Ӊsg!�W}p�]n��,��@$$��9�`$�n�ش^���� A�l��4pI�����C�]�j�i��ہ	��5��lγF�%�0��4�G�H>����7�i,'�0v:`�F���z�:޴3�A@SE6Ri�b�j���R�G�1R�	3ۓ��{֗I���5#:kT-w�+e$��&A��7NӻJ� �D$Q�Kv���Q�PRZ�M'v��ޫ\Bbr%{Z�8*Ę����}�;;t☇5�y��1W���&J7�sDØdYd��ͼ"�+���M�g]��M��&����-����Mq�;+]p�������3 aE38�E�|��w˚޻9w�;��O�����p��b;�۷z��l�$�$gO�;�]�ERe�I����I�ĝ8���o��e�޺��&�}��sI&Z0�3���j!ݦr�N+��/wԊF�RRxF�$�l&�e�pזk6�˨h�H���g#Ndj�*�9Ǘ#[#Z��է�7�1�o]���GB�����m9a��Q�����#6�^�!=�wm,<8F a0��"#�+i	�q;P8Zn�HMA5v��%w[��nvW�G�g�s�}{��"��Q�lt��O{���K��!���oӮ�;�;�6.$00�a���������M�98�NNk��^��ѹ:M&LNTHN��!��tRc�ڱ8��u]��%�A��	A��5vk^��\f#7R�ՐdL,�[�������!�11g0'��ޭ��y���׉���F����IF$��̭����#0ь0I$�3$c`g�٢��<l���m,4�2Q47lbt>k�		���֋hTr���Ui�4��75k�������e�K�v��&]�:p�#'�0X�&vPƵw���{�{��:�Z':;b"��z�ëq��֌'4j�£<�����q�`s���g[��X5f)fm�F�ah����C���4̄�8j�0��f�0�hc0H�16�A�Ȃ���2��dkD(�O��!�0�N)&|3ܽ�;rx7����	y�f%��ht�Gw�<��Øp8�?d�M�3�`b�㳰�k���Q�%@A���� �I'%�y�=,�xp�4�]������&'f��\���xBm���|Y��"�0�¨5�{�Z�^���3�I��ɚq��rBBa�6Pd�D�c �F����bM5�kL]��n�� !��*&��ah�IU5B�0��Re:�!4h���E��Dӱozݭ��έ<'z�,vEa�q`�q�	�Hr	1�c	�(�[��*#"$�&f�9�1���X�Y44��d�9c6��aR#��J�$�28T��aTc���6��ChhL@�4��h,��"�D1�"m�hE�1(�C4\5�E�4Xh�ȳ]�1@L�33T���L��L33313315LL���L3 U���EQN���(����h����ȟ���{����C��  �   -� ��lS��    �               ���                                                                          �yn�0u�m�j�[i0 �)@�<sQ�pUJ�\�w)�5^�ֶ�H����̨ܯLةh�nm��#aRB�jkT�UJt�ʆ�<��m�����c���^Zڪ-�mH�����-��m�l�   @  6�!��m���� [@   �@      ll    H6� 5��U[r�m�o$m&��4sHm�cm�BM�b�$��������ľ�z�R$"��$���1"�tgH�d��%ۡ�9�AmH���c�-�T@�*�*Ԫ�lH          v�L  E	i����z�m�K.�m�-�5����]�h�i�Y� ݫv$$��ku�,#%�q6��t٢���K)�����/U�<d�V�/]��Z
駝uRն�  � �`��1u�H-�$R�<@ ��݄�l斥�Su�y�V̅�[��8 �q�Nk�C[v�m� �J�V�V�����?$�r�O/+g�e�\��Xw�UWW<�Nwl4�A��D�F����C�$������m�+0b�����(8�]��M�A/.؎2ҽ���3�^ض"q����
U�ڀ��:�)eZ����ʴ��m�� ���dڲ�!r�.�J��;F��[%�o����6)�F�W�T�5UU	�c!�l�kaZ�����=���x[���^��cɫ�ي�b����Ë�3�vi��X!ٶۋn� N������bk��jÒ::6n�Х�m�:7c���y��ֹV1 H� ��&�I��M@�S��83�e��<�B�b�a �`	6��v�3�6�6�'����!. q�mf��.�ڙZ�(�,��}{N�s��z�S�� hm�4k��$���V�.�j���`,gcdI��n��Gv� �v�H��UCh��U]���j����ׯ@H8'BKM�^ӴC��tL�\�dj��:h
� 2۲ʹw۱��S����ݙ��)Å�Q�EvN�}?}��o6�nFC�kl��G�'.�2ݺێU�w)���c���%�ݮ�������n+�Wr�i���/����\kc��Ʊ��aB�a�q�t/*\�u�<�Zӝ���6��������F��m�:�kh����F��-�B�'�����K�W̓� 6�:s�[[u���[m���[[m�ԋl�l�$[y"���#&�M��;sJ���z��ä��c�lr\W0SK�y�ƴ��xNm�gNM��M�ń�Y�3`ử�f]βؓ�(�SN� K�-�
���kƋ��i���a�Cv0�u�<g@� r�S�,p@tT$���Q����hS2������t���y-�[[iMU�v�s����%�P۰�#�v���l��1j�������1x;e�qibҭ$M֥��8�zN�mK�L�.2O<�ݫg�/@��mw��t����I�U�va�ۂ��[[l�`w[�
֖��Zu�nH�][C��6u���$սܤ�JR���ѭ�����j��Q�i�cv�ṥ�RS�n�:����5��.-�H!�l7m�XHmN� 5��e{[i5;T�[ɍnM���ݥ�`F���6Y[�l�ڒ�-��5����<��7v�����t�.u��s�E���z��d�=�/9���[U�j�D���1�i['e�m�Td����n�`O$Y�]q�6����\;�j���٪B�1�����b�&�aܦ�U��Ş����BA�m���FZ�����W��$�姕�%ڥQ̒�Ŝ�%��g������n����C�$�A�ӻia�MS�U��V�8�I����ݽvM�*J�m�m0��[:p�um�[BI���
��\����n��3��ە]�t��YYj�[L5U�L&BZ��	T'-O+�m[!4�+s��UV����ٶζ�2[@[)��nNĶƲl'���N��<�ɑ�#$� Z3���i	�q��W*��� ����%k�ծv�ɧ���7cwa��:�l+���7m�T��κ�̨s�Q뮗���S��J6�&�R'�kcC�0��ⶣ�$W[�2��j�m��݊ ����YW��P�[m�4k�iV�VV�D�$�V��\Z���+i7$qm,4�8q��"@�z���I���m�����j��iV�st 6�V����v��n�pi,�� K(�&iɵĆ� H�Ib�l�iIeF*�
T�y���v��sβ�pL#YF�+N׭��Uv�iVt+�u/\	j��Nu�-݇����g|� ��d�}��*��'��:P�~?p@�_� �R�;�t���L@.!����<�v*� �_;D� l�>��tiD��{MB���VS�U��']�AN � ��Q�� !^x�2����D�$�F�;�z�:Wh�� �
����uѱ�>�/b±(��/@h�y�� �Q:��OG@�z�Tס�Q�v'H%��C|O��)�HC`�rs�'%Ҝ�LziW���S�6J< N�@��D�x �~���i]�iP�_EL S��"�+�����k�@�O�j.�z:��Jb,p&�� �!�K0����D�%�I�2p0�VT�pd�î�5�N: =N
�D�6�Q�j7Sciԯ{6��ҟ� ���/�'W�������aK�	�]�w�����Ǥ�mn�nm� ��              ��uS-�{r� ��6.��D��+T�R�m� EZ�w[��Y`j	z��7bg�`�p ���kmVce�v���R�w
6�:ԎmS�g䁦:�fG^[�b��U�m==��u���c6}�H�pն�۱��ݰvE�1l�<��!����U'%�;��T��i���`l�E�ŵ-��۔���N�a]�I�{:��-��ő�yJ�/��v���-"q  Y:λ��N�UJ�UZc��������q��a���X��%r+��2vs�3ꮓ<jM�Ӹw�#(h�3\	gdon�G)�u�!��,�[�6#�'N,���6�AHI��$v9��K�ɝ�9�k�m��65�*���NC=�����`����M:�h��n�p�0˰<��s6�g\�0���73���G��UБ�r�D\`enհ��A�Ձ�hUbc^Mou�x}�� �?`M��@��E>N��~ p=~��P�;������m� �rl �\b�U%��i	���8�!m�,T�y����!�;����ƒ����oh�Q�m+�71�s��-�M�HqܺLq�&���Éҧ6��y�;���L�.�EG��ە��M0���v�{Q�!"7��=����U��#���Ub<����f
T�pn�����$Б���ׂ�a$rFs����V��N�t�wQ�q��y��$�D��_�{D���sa.OFJ^�\�wd[b�]�M�b�>��b<���y��7I=��|�	&G,כ2#��пG�1����}k�=�����ú�;�bD:�����j�$}��w��{���L+����eXo&�01��v�U+�� ^���M�}k$���cN��� ��<�d���6�����N� &D9�`��IQ K��'�ܯi�� O�VH=�e�m@�Cx���?�f� �Pݬ�~��X��I�&7�"q�y�5��,�ܬjsu����V�	�@v�A� O����p5����� �d�" ���'�z뉪�T�͌�{����<��2 	ٙ�I;iR\$�q�N� �I�p�Ud��^�8D�H�X�� ����4	�z9�4��! oa��l�,V+��lM%V�. N� ��2A�D@G$`��6ӱM L�d���&�X�E
 {��Oj��� ��0L4	� L��&��������@���Ny L�d�" �s�Mjv��	�@��H6�	��A�I�	F[�$�  %�ٝs�AC5/J�u��Ѣ%2@���nݩt�:��nrsm�x�рET�^����t�qδ�ɱ�x��;u��qp<v��5X�v��L�%>�P�绋}���+����7n�,jݫb��O���;��j�$3ђq MϘ�	�m|q��x�m@7�ڀ&�d��]|0�I N��'y M���<�n<�lZt��@��<�D7# �w���۱M N�Y � 	��	� O�@&�w脙���hZ������M�I;��H2 	�� �D�20���3.e�%U�Ȓ¨���H�#��2�$�<��5��. N� �� �	��H<ߧ����I�P#��$� ��0	� K�����,Kăj ���&�7k$�����Z�v�]�ggi\x��1� j8X�I N��'y M���>�y����^ �P��$P�X�����q�HoՒr$� D��M�}���X�`�ăj ���&�7k �����`�V;�n�H6�	�ܯ�eGX��,��BY�E��g':F����/ M�wy��e��}~���j�$3c$� ���N� ����'X���3y�M�n�H?e��5���w�ݬ�0		�}�]o�B7��j �G��H2 	�əv��m+����ͤǮNK�Ss'����ɶ�ƀ&�Y � 	��	� O���c��A� L�`j ���L�U�`��	�@v�A� O����p'��j ��d�j �k$_������I L���9�<��2 �|U����)�E! �|��  �],�v�� i�n��3�k֪TGr�;S�:^�m�A�c5� �>�ь%��`"Sj��Y��ڝS�Ǎ`�u�o(]!3v۶mmw}�ݶ�8+��7Iۑ�/뷏�>�N��P:�K�8����S	�t��I�J�� Ȁ&��d@v�A��|�cPb@��	�@v�A� O���H�r'�	� N�2A� L���/<M�ƀ&�Y � 	���	ʀ'�n�k)�ăj ���&�7k �z�#Qf0��i⋎nܺEd{W�"��b�k�a0	�� �� ��>�D�" ��}������8!�0�>`��(�
M��<��G��nc${��|���R@62A� 	�ڀ&}y���K� ڀ&o0	� M����cƠĀ'm`��&�d�j �{z'�%$�21�F�H�v^dF½�;*54? M�wy��e��~ѵ�ܑhoՒr �k �Q#� �����m�d@}�$ (pr�&X�62Q�ᙣ	�Clb����!f�M�hJ,�(̉����h֜�	�8saf��.`k�17�s4h	����O��g���������7�مjͻX�A�k��5�$�#dxc����p���C���a2մ#|I4�M[@�M�$T����SBa���"`.��,b"h��{5��$�g5��0�5to��Pu�X,���k����CV�6�g��7@���|�| x�'�>��
����\P�{�}Q�L�+���%�'�� ��T�N�XL=@���y
t	BP�%	�ؔ%	BP�	BP�%	BP�%	BD%	BP�	BP�%	B|��BP�%	BP�%	BP�	BP�%	BP�%	BD%	BP�'^�ݬϚٚ����(J��J��(J��(J!(J��(J��(O�4hJ��(J��(J!(J��(J��(H��hJ��7�(J��"��(J��(J��J��(J��(J����(J��(J��J��(J��(J!(J��9���%	BP�$BP�%	BP�%	BP�	BP�%	BP�%�ݷ{�_���-�����js0�s�sW�G_C�?dױ�w�nJ��(J��(H��(J��(J��"��(J�7�(J��"��(J��(J��J��(J��(J�4hJ��(J��(J!(J��(J��(H��(J��ϛؔ%	G���J��(J��(J!(J��(J��(O����(J��(J��J��(J��(J!(J��:���,��2��(J��"��(J��(J��J��(J��(J��F��(J��(J��"��(J��(J��J��(Nw��%	BP�$BP�%	BP�%	BP�	BP�%	BP�%	B|��BP�%	BP�%	BP�	BP�%	BP�%	BD%	BP�'��obP�%	BD%	BP�	BP�%	�%	BP�%	BP�'^�皳e���pJ��(J��(J!(J��(J��(H��(J�����J��(H��(J��(J��"��(J��(J�����(J��(J��J��(J��(J!(J��>w�{��(J!(J��(J��(H��(J��(J��>|ѡ(J��(J��(H��(J��(J��"��(J�~y��v��{�uД%	BP�	BP�%	BP�%	BD�	BP�%	BP�%	��	BP�%	BP�%	BD%	BP�%	BP�%	�%	BP����%	BP�$BP�%	BP�%	BP�	BP�%	BP�%	B|��BP�%	BP�%	BP�	BP�%	BP�%
���b�� {�v!BP�%	BP����J��(J��(J��(J��(J��(J��(O�y}kY�k\-g�(J��(J��(J��(J��(J��(J����{��(J��(J��(J��(J��(J��C�0 ����߾`�I��$����.ݪ`�6�s�R�z����Z͛�6��U����}t%	BP�%	BP�%	BP�%	BP�%	BP�%	BP�'ϚД%	BP�%	BP�%	BP�%	BP�%	BP�%	BP����J��(J��(J���H����*Z�b�&@=����{��wP#� I�̧IKip {R"��  ܌�y���5Vi ƈc � ��� ��
N�$�D	>G���~����¸�_e�  jd�	[ʃ6��*]�b����خ�\��U��]�܈ktt	�KG*.��&su]p63B[9d�����]����}�p���cv�ڝ�5�;�Y�Nvݪ�ǻ�5/U ;p-[v֋�gf:|1n��ۥb���䌐{�gc�(�$@�<�v��ݷ�A� !"�#3̐d@r2G� @�"�۰� ���b$�:  � �|�������Po��� Q��<�DA �3# ��T�����{# M� �������Wn�v��+f���j󬱵BG}���B�բǵ��{�Y�*��ȷ��[��H�G��B��z�y�|@I	���I�$����o�� _|��c�:��vC�k61�Fv1� H�d��ӵj�	� 3ޱ"/c�Yk����c6`u��خv��-�@Z�I�Z���M����_�B	Ĉ�s����PO��āB��}�2c�9�R»aY�w@�p
 EQ@�5��y���X����v3��!�\�vOt�Y�d�  g���_������Y�C�W�2�@��q��.e$����c��e��BH4$��t���IH� � ��G﵏�^�ϱz�ڵv���1���ވ�Sm�M EI4y�:��G��A	B��`!�p� $�g}��I5�$F /޵��3�x���c�Ii�]�q�r+��]����fܭ��/�\Wk�ݑ��2d�"=���)b�.	��P��|���<w��Uf��1�C� ҹ��O����UI�IR����o�bD>@_}�O��uN�H�����?}�}�?w���   ���mY��	$U�F��s�mZ\];�i�*Ρ|�nٓ�<e�u��q��TJL��C=v}��n�o����sr���fx7W���3��Z�dˮ�^��G�#M�6N�^�����\�q]�[�������ӫ��o�#��>�@ �r10E�M�a�d���nF$^$�C��Ӥ�ʧO�Dy��@"�G�3�j�ث
�� �!o�1��>��I$}�<���R�:\#	����r�<�wJ�WcۅXբ-�\'pI�;��X�G�1�G�@	�UH��Πr�cf�̓�BTRBH�ĴGA	�L��d}?.��2@6�N��fd�m�jZm��]���yS|x@3$ �s��R�ۓA�y� �� ̐;T��5`gV\�.Ir=ׄ;۰7�vd�g9�]厱��Ո��.�v91*�����Խ86M!�>K���;v�O������ߞZwh��@s2��)� ���}��J��m�h�k�|��U�wj�_�(�I�e>�!��@g�,��	u�r�����SDe�zUU?O�; ̻���e�3��@���� �%�wZ2@6��b��j�7&��]j�7�*g�c]�+ĒU�55b��6�s.��doI*�l3$ �w�r'j�ɠ3$��*J�ʩU)���}��R����W�=�\�@y� �$>IUW�UR��}v�H���&��uURT����n�̐�*Ԫ���I�@R��V�x�U!ψ�y�i�E�z����R�*T�5�:� } �>���pzh9{m1�v�x��N��J�jkH���6�@q�3&$���k2�fyM�hz �9�J�$����.�̓�*I6c�:�Km��� �]���T�d�� �M��V��ރ�T��N���d�q��J��J��j�v�q�v��} R�R��=��}v����U��I��T��`�, {ސ�?vv�b�֮8o�f�nb�`"c���ΝӼ�<�Ϻ�$	��0m�             ~0�   9�*�\ׂi���q��5s�k
Ҡ ԫ[r�m�  ��K��Y\he���gv\i7%�d��̀ ְ�i�a` ��EékjQE
����ځ7%�n1 :=��u�x�$����%�ΗC���+su��iq��i!؜�RJ��ⴡ��v���΍A��X�ۧ��6Y@wF��V�vĔW��r�	�ë3P9U9�9�sn�uH ŧ\p,'���)��S�w���ڝ��>)4M�.���I� $�ѻq�U�Uj����<vv��۰�5����Od]�����g�g8��J�qyM�v�`mS����b$�.�*��m��T��.ݸ7;/[���J�x\��Y\���ҝ�R#�q����-^zv{{��sV�n��N�LC�0�K<V��$�\qe�!�식��]�ř'�N#[�s�M�*t���pu:��Я���X\9�Ɲ #˶69�f��7nV"V���6�l��!wiX��+�1��@��A
xІ|@;^
�����Bw�O�t�E��w��I$�H 	k-�/fة�Wl59IX�'n�G<կW����g����{�R�gӭ�;n7��OW]�-M���nv�Y�"��r.��]�I�q�����=N��+�$�e����U��۔;�j��ԧ�
N�4��q}�j$���u�9� ���i����1��h�@fI�d�T�����p�9�T�k8���ӽ�˰u�ԓfu�3$ ���c��惩&� �\2@�OY��9����^�lo`c�}\����� 5��n5vL֠�N��88��:�#	�/(�ZA%����̐�.�3�*�j��>����KM�����J�3 I	 ta�"
B\��,[��p�pvN�{9}�ӻrh1�q�3$��;��R㖤z �������=� ���Fj�zސ�.�;� =���~~T�s���fD��n:��qS9թ�$uz�|}��:����fH��� �3 �ސ��񳙟��n��c{ �� �$-b�T�$��O�v���� ��z���j�����RJO��s�݄�����|�� ̐ɾ[�mݖ�\B���n�0#ї�N�z�����$�c��fH��;��R㖜z ���{�`�k^E���z@5�]�{� o� ^��i�N�U*_O}�����p>���I!���IV�W���Q:ݩ4������]�� ̻{��;#��Ru�k 8�:ݽ��')![��V�zm�� g��H����1�1��A,�1��&6o�� �px�ɾ[��i��9�]�s� o��H}��F��[�A��� 9� ̐:����Ys�.;Cz �8�˾ր��]�}�:�	$�U	��w�_��$���   ��`�sMV��g�g����gV܌�ͶTV��bV,l&ޞ����t��k���n�A#B[\qؔ圢t�>n�rm�.���[��)�v�_9o�w{��ݼ���0��u9�)�>)Zݎ7$�����ɳ�xO����^�v�ϋ*��� 9�,�內zy�`��{�b����&7jA� f8�8u*o2@5�v�>��m��2�M��s�}v�T��p}�PK-���3$�_$�-����8����v�dj�2�[�bY۴]��p�O����������KM���˰u��ʪ�J�fH����K��&�3����R	�D�"���sU|�Z�y�%K�URRy}s*\v�����Hu$�7��� �p�9Q�Z���%O2��n�3R��u���-��Ӛy�`��{�׽��t@V��2�)�E�nD�T���&�� ��3 �2e$���.��~}���lo`c��UU���;� �����9�T���:�Ylm�� �]��UR����4�Q*�TY����ɾ[��i���S�f��p8�v��e�=�}�	v��c�J�YS�z2@/2�7��w�q��O�8+���щ�,wE�<M䋲~������@/2���c�s|�ɠN=�&Rl�;v��qϩUUz@�u}i�N�~���p�6}� ̐��&7jA�i7��z��N��F�7`s3��ޛlo`c�o�y�`�~R[�����wj49"����X���N��=ަ��mm����.�>��*�u�=���p%�ހ�e�RI�� θd�$�z�)����a� �� 9�����@5�v���j;v�y$��pv@�d��E�o���8��k)R޸�߿{��S��߿��6��  @U�9,P-UR�^I\7l��O���v���S�v�^�$[%�=sk���@J�������p�.{cN���;;'��vc���=j���9:ķM�u���&n2�;c�ٲ�v��pW��y~��ⶻ~���>����BDw��Vi�#���/� (}��Ϣ�v~�c�8�$�~���������Y�N�$�C�"�fH��Wڌ�}���;pw���2!��w�M�4�5
����7vc��Eh�.���̕�:��$���KV�Sᚨ�l>h
�$�Hĉ1@RI��Y��+41%2P��A)$�t����_�3���$�����N�M|� ������_"��v*�pw��y�� $���E8���3$b{�ȃ�������|���]�n>Z�a��n݋J�����pX�8�*^?�#�A���$P�1+��T��I$dA���;�� >���ڶ��=���<�F�͉������1)��5����M�xN���p8K�M�J�X���("��MF2��T��a�t�M�����6�C�OA�(��
L'��=��I��x<���p�'bڋ���� �$��z6�s}pv��τڒ�ӚWZ::� �Ȉ�J�]��x��
��Ha�b'������QҮ�*f���M'�8G�C~�=.L�&�Z�r;�=�s���Z�b��=��
�1����&��b::]z̏3Kf�5W 6�������������g��7���X����y��wQ��S�V����u�{߼,NqRT�dG���Ϛ=60C!@-*{��xf)I$mA�Y��y=�z7�GWZ�M��g��6ɺ�1�"l8��Y����ڇ�<��2�6�{��k=���-E?Q�A�͵�����Ȇ4mA�Y��yO�X��3�mg�����P��_=�  e6io[�mJ�U]�nU�EF�����P�;�`q��4�X؀��-����N�MZQ�Z:z��S	�n-���N�1ѳQ�{l��b'r������/�T��wv�/�sfz+�g*u��Q+�E�кWTի	�g�3���=�y�O��:J�L��r3��mgpSWm$�;�>u�� ԑ��d�ܴ�v���<��mC�فɐ$ٶ�܍�;Y��_��@��/<���\��j<���4p��mGyk6�=��f�3[�Z��s��D( �$Ã `�,����2�7���U���3�mg��o#j?Of5T	�c��H����` ��}?h���t�.��=������������δ&��Ԝ6�q�h6a������}�4 ȃ�Y�Bl�#�3֛X����y��wT��ܺذ�fH�b��n�   �s|�z7�ūV)���A�mc�y�x��2#j�͵���|��ﱪ�%����6�	8��c�)��@�̃4u����n#����Mj��&wu���������w��W-�T�~��r3��mgpU;��IP~�m�@/#���Q�b��Y����څ�v&�)2(c�ŏ2@,���xt��n[���g1߀ .F}�c���f�C<��̑�v,�wt*��A���;���ն���	�,ﵙ�xԈ�:)�V�̑�@�yr3	���]'��}��   RV̑.V2\������ ��`M���`�f�6����m۾�NS��P��N���-�H)��Y��ӆώ�%�F���㶡�t���U�ܔ��������uqd��3�觨�.����j�jH\��kF�c�{o�Oߙ��s��5#IbF�'��k;Q��rҺv�n���=�>R!��.�;�d���B$���mX��������ksZ����Ɣ�$7#Bn)�BxB3t�yp�B��:�����{�ʖ��U��쌀8�A��ћ�mG��܁<L��s�� ����޺�qp%K�~G�����k��r$�$mBn�mgj?{�����$լm�i�A�t�'2dS��ۑ)�<��ֳ��7���{f<p@�f��r6��g�}_��V)p��_O�<�����v,���SC���3$fb<�z6�;axm��|��mC���N,R$�(ぇD.��tf�X{,-�څ:L��9���.F{���|�����G�����Wb��SwIU$dA��a5$fy�ܴ�������y��t ��"�oP���b�V�n�5�#"2W���n+A KL�]���Yl���Xx��g�_��_��Y����5�L#j�͵��� P��	j�X��=#9�g��}�U5[b�&wu��;�^�<����\\	R����O���a���"I�tc$3�CUC&l>E����銡"H<�|C�ھ��*q�;���1/��A�QR���v�]R�%P�����k�w`Ur�l                 �˰Йwu]om6�N�tgk�]�%-J�U���   ����!; (�'dPf���a�-ۓ��V +j��x�M�Ny�q� ����WK6vUL�O@�/�����K���6��l`��S���۱�p3�XUY�� s�ԭc�Yѡ��7nM�Mۧ��� �jk7h�.2:v�^c���[;q�.�C���`�,EǞ�Z�	�od���4[y̖Z���ۍ��e�] m�yʎ�` ݥ8͛W$���r�'c��΃q�������Yź-�\n����k�ậ��v5��j�[u�d�p�X���9)��5�k�w� guu�����<X$��:B�Φ�c�Es�t���5X�]\T�0�$��8����Ihm�6ˢ�[���2�L@��K�AkE<gc�n���u��y��E����8N #�m��:<�P�`���nf	��
�[{$m���������0�#�{Mt��l�����H�;=A<DA�a@�v�  �G�~���?��I$�H �4yn�l:�ݗB�l��.ڻu6�l�+�`R�Mwa�Tq�Nb�vwg���p����/kЩf�ۆ�ɮ��A�g��n{vK�EI�+=
�`&bG��f������E
�e^�hL%2<����-�UI��g7 �<��g�+j�S���<��;�kgS�Wt�7l��G����������mGyk6�7גk�ѵ	�f���~��X�[3ӲX�.1m�U��m+�v��U�����y�ꀀ	�����)�fH����C��{������qp%K�b=�.Fwu�j̱M�%I#ju�k;Q���Jc�1xu��|��?��������5vJ\{p4l�5�9^�C�pO�??~�g�~ ����K��Rᚠ C<��̑��U0��	����XCH
�Y���ڧuV{Y��=� 5";��5R�:L��#�����O�§��{q��uv�[;��2�����9�:J��=�/���9�2�7t�$���@��̑��vgrҺv�n�����ڇ�V̍GQ�k;�ڃ �h>� �t���1A/Q�A�Ϳ�?����}�H�)�T ]���rQa�3�N��kvO?�?~�$gq_<��;���;���k�hO#";|�j��t��3���u�{��\�IR��Fwu�j̱M�%T��C� 7�fH��zd���wwwww` nl��M�z�a�I����M�̵MqN*բȂ�U�a��np�e�O+�z����'�8:�=�mƮ�q��+\%��f9��e�������?RˋC�3:��SY�,<�$�t�Lq�/������F�>�[2dL%��܍�;Y�W���mGy|J���xP�o4mA��mf�>�j�d��/�����l�0��Y$2�vG��Ejuj�#�UMUاI��g1�X����/��%K��� DD��!r3��� +�{�)�I$���X�"���#���t��.H ���{Y�FD=�]�v�4����2!r3�����wj��'GT^z.nǛ��p��RK�����c��̕�z-�g�E.��;� +��d��#��V�X\��w͟aI`$�Q�|̰S�ϷY�#����{���:J�N�{���������??g�ȥ�X����jH�t�� ���&�6�v�����b��_�|�ڍ�}ul�$P4ٶ����KY�W��oug=Ǯ�߾��� @	""��/��T�;�#���w,��G��cH���+���#H����Y�9���L����Z�w��F�7���:L��=�wP��y�}�r��IR�؏q���c��,Sv�I#������
Ȏ�g�!n�R����=�wP �	" F�M7d�I$�I$�V���`	,�GR��g����D�p�g��H��<��(\�X�:�a���U]tm��m�\��s
<R���θ:;���w�:9ܮ{v\D��;��)A � �0W��D�&%Lne���=8dG�yt�	0I6wk;�ڄ���k���x�~��!-f����X�904��Ok6�v������ֳ��;Q���2��6�w��	k>��1�Iy�S=l�Y7:�ȕ��t���_+�t�.������9�2�7i$�}�8���Ÿ�'J�z	��;��w����HGb��Y����ڇ�S�P$ٶ����KY�W�M����Q��c�3$cA3+-z�MU;�j�U�j�ض�DQ[7\�2S���2!|�2Fw���j�,.�w�"7�	�K�3$g1 ��c�L3�o��0m��'Y�4C	�c2,3�2��!����i���6�0�0&"�0�+�3�D���Čуod�iz�iK��=�H4H�AfB��%���9�(�p�E�_���
�s��d�$� ���@t@��G�i��6��AN�Q� � ���; ����7δ�>���%K�D{�9��9�2�7i$�;�M�m��F��<�L�I�1F���c\�p���svQ�����w�gj6��ճ� I�mgyP���>�✉��������k�8&�oq���p�:���اP��I+B%�B=�T7�c�{��ٳbᶳ��7���ޱL��E�%#��:�j��[nyꁎ���3��s�A�͛�r�n�K�D{�9����b��Sv�T��޳$gqo{���j�pwu��3�� 
��Xi���fH�5�FD.Fx����ۻݒ=�  �,���W*�j�v	��y��UU!��b�9DRs�;Y�nq�Nܜ�{2�lMI��1��y!&E����rd��&�Ӳ��q��y�#�
6�Dm����܍�׿;��ۮ�/��l�]�kN�,���c���h���)ȃT���!~�  �F3'�&���i�u��g����V�apf�=��T+"2"����)�La�#9�dB�g���\�J�t�G�c�|̑�Tǖ�[wI]�O��b�v��������fd�I,Hڃ�f���~����^:��p�MI,1Z�pY�bX`2 �!����>��C�zq1M�k=�ڃ�����NET� +b9�.Fd�w��M%wh4�̨Ok6�v���؜Ēb��"�L�x���۶�q�1WZ���Y��gj6����,�&m��#����}<.W-Ҫ];�.�zA�g�X�]�d�b�Hڃ�f���~�ޔ��UK����wv��2!*��.��I�T0W:km��tU�Ü�@�p�yM�k=�ڃ�����NE��mGyk6�7w*i)"ѵ�f���_��@�>S?w��C�(�i4n��:c6�{��k?�'�_����o���ۉv��\��Ŋ���V��_�|�.)x�����;��U�G3$��M�m��_����}�M�U�H�s�G�V���ua&���KY�E�✋1�ڎ��m�g��]�<�_w��@   �[BmD2�J��J�� l�Ѷ�$׮����m�&��}v�x6��y�p��P�^����vܣc^Q�g�ح�7kn��lp]j�zL��\�p��:t�\��߿|}}'��\�w9U��v�O%�nC߯ï��k;Q~�U� ��ֳ�|��m_����%�b�2F{�ȅ��߼,Np$���	��9�/1�Y�*��*IP���Yڍ��mF�� �d26Qu�-ۨcr[az����:�~��v�jeק�l�]$�x� �|���~�k���X�~��/�
���{Q4�vC���w�� Wb7�bڰ�Z����{�g�����k����X
FS���N���Av�ӻ�j�h��7+3%o����y�����B�N�{�\������]ؤ�Gu�X�_p �A X�ٸ���ZI]�S��Fs<�u�6����v)�wu�Mg���������nӻ�R\�7�k�W'��ہbs~?Tw���mbf�x4��$wT$
�q�#=��9�ʕaصK��3��;�Q���,�L�Y�F�7HAU�Û�h���HR�؏q���f����n̽@S�d�P�ڧ#j �ȚnA�A�$��Ok6�v���e���U>���}�g��޾��ئ���{�B*D9#>��~I�|>���� �#�SʛIXI�u�����!��ކ�&.p!o|���ѫ0Z�3	\��0��t\�V� �P�E��$'�Ϗ���� ǣ0�7&�5��L��d=w	��:L ��٘���P��3��{Hi�Ͷh                 ��)�]3�n���Y���ڕz�-��b�h���l *�J���#�Ѡ%U+%�9y�<�����f����f��
@*�)�u �g+���`�j�6z��K�[	loVx���l� �r�ݺ�9:��
�'��T2��k=Y�������v�'� �%GC��v�Zh.��i�f��k�"���t�9�:{�b�5� x�@Mr>vG���
M5�����]�NƼ�sI��O`ܓ�V�Wm��WN��{5���ӱ��Цɱ+�)�9�v�G6��V�����"[�˪�k���f����znܝ���ŗ4���;=�aPg8�$f�j��U��!����n�홁�x��&�m�v�����C���=�:�"m�N^g��t&�Ը@���[9�z�-���hZ�\��2U�&�L�\�l׈b�t�b�j�s�E��c!�5K�-�]����c���㆕3/⨜����6�M�^��v(��h�
)���#�zL�������o�  Ilk�Ӕ�cR��T�eqjL�F�b�la<[s�v�eke�]қ����i�]K�gF�]g��N�la�ig`�&�u�>݀�bɹ1h	��U�֪Q;߾�o��2�:�gn;:�I�E!F�`jjb�(�Q�Y����ڍ��1`�f���6�-g��������v#�_�$W>��#1�wa$�2!|�;���G۝�I+��|���G��r#"���-6��J��1A�wYi����Dz�NEo<;�2F{��c�3�ڏE�wB���'�NƎBZ�ubf�ʚĠiP��m��FO�\pE/���ڎ�;�
clS	3��@��2!r3�l�d����j:�Ħ�:�݆�mպ_pX�8�v#�B�	#�ޱI���FD/�gwY���e�����:�{�rfa4�TmB�u����M�  �݌瑑���_����~��!-f���k]#�7�8%��Ց���Z��3ئJdMbP4��Ok6�v�'ڮ8"�n� ���r#".qS�0�;��q�/u�o��9���ӱ�#�,
$��n��o�by�bHڄ��m~�~���~�q�Vp�v�Λ%��a�H�5���#	�"II��u��|�u�6�����Rl����y��G���9�?�;�KY��3V�MbP4��Ok6�v�'ڮ82L��ֳ��_o>}�=����t���   �]�Rҭ[<����K�Ek�@���ku0뢺��q���\� Z�N<�c�9y�pG%uQz�y�<���[n<�7�y���f�8+�����=��~��-�k�fny%����9�ۅ���vx?_���dB�Y��xX��HR�؏q���Mr/z�'Ub�FD/�c��*F�u��x�+��7\$P����Ȅ����v)6w��q�/u�wT�wUUL;ݸ��X}�NSz.��nä���� �E	#�C����٬����n�iC�����0��2:M �3�i�޴��/��kV�R���{�8�ȋ�TıL$̑��;�^�<�����A.���!?~f���Ϣ�3jD�Y�$Ԝcvf�:ޛt�GKQ�	�f�Yڌ��|�)0?���ڍ�\�����6�w���|0� �$�0� @$C��>�?��;�O�6�=���k	�ju�k;Q�۶'1$��1F��y�f9�3$���r#jL��ֳ��;��	��%�b�2G� P�r3ɿ�,}��.���#;��5fX��X����H�3�1�I%�!(���|�)0?���ڍ�\��dqbm���\�m��T��]��Qp�o����Sl��#'��$g�$z't-��#�B�Y����X�Jj���2!}�2F{��=�����ē�,絞�>W�#{М�
�&d���B�w���������   �/P�2
�N��U�=�����4­s=l��̫����m�9���S=ogvy+��P5�S�Gr�֚s���giɧn=Z����#�.{J�`��A�m�hUT��UT��9������v@����v�u�R��Ϻ�����}�����D"��|�|�lSb�RH��޳���W�El^~T�������>{�~�	_u����m�����;�^�9Ѻ�R�-��Q�<�$fH��˴)�U[�Źj����|���*pbf4bP4��M�m��F{����g��^� "A �x���γޣ'Y�М�
�&w��qޱ��{��E��B�G�	#���>�1�ߙ��1�ǖ)1V)$w|�3�k=�~ L���jƝ��.d�["t��jI��-���s%s���u�i�����pcl���#o����������o���QU�E�F�P�ht�m8�ApTʷu	�1�� ��Y�0�1, �&,l,f�P[�;WÚzprw�0��+�h���y��섉#o=��v��� �"$�@<܈С��FXZ�@�H�Z�8 �o�T�'J"|_O;DN�j�)р�uuޞw֎]ax5�A��1;��Y����:�Rf'ᶳ�k7������*D�I�����h�N�i�:���Rgی�#��/u��h���H%�"=�1r3��9���7Ub�#��/1��gq~/b��J��S�� �}�fb v� � *F����a�	�}�g1ޱ{�������+�%7N�Y���H�H�6�<��&7
^6�ݬKY�k�����SGw� �y����� P�;�[iX��H�s��Gw���	܁A�����m�%���_x$1tȏ���'��F(A�  	D*}u�>���� [r9�3 R�C�eZ�a!�ٹ��u�I����mѐ7�uvֶ�v.��g�r[*�v��u�wW���v�Y6�G��6N
�v��gulɗ]:�v����{���$2ձKմ�#��n%ܲ�q9��h�-u��W�J�c7��UςY&�6�{�3yu��_��	6n�{��X�����1�R����G��.Fg#�8�J�n��M5��39�F��껷j�aUݤ��g4��u��[��)R�a>�;� ��fw*�i32?<<A��;|b�Y���7�	
]2#�c#;�b�X��U$w5��f�f�3껦%�`�ᶳ��7����������]Cۙn�Y3u�H�o �G�6�Mc�&���r7Չk?we������k7k5Z��%b�;����	�#��Q��n���ڷV��$���f#9�tPw M&oV{���KY���Oq$����-Q˷p�e�����r� �L�������X�Y�)1V$w5�\�3231س.����;��w�P�Fv1*u�L'bձ�jz3�#9� n�
�<~����y
~6�Ә��o1}��H�ME$�X� LC�dֵcvg�t�hLd���&�6�7�s�+Q��m�����v��ބ�U��gw��!*r1�����	�~��񋑝�b�X��XT��X�����G�t� `�h��3<���t  KK��x ��VCRIe��4��U��vl�����ݶ��'xm�S��NhnўxS�3#����u��<����nX�λ)���:�6��Q�m�\IJ��P�֪�>�������v��EA���Y��'-�h��w`]�����J�wݺ�.�hNF%L~	��Z�d󂇼��b�|����:���9x��]uw*k�7ky�y�ȹy~k=�3y+7lR$��Q8ԁ�blS�n��˘͹[�b	����GoX��{��cҬ!K�E�I6H� �׌\��q�\�ޱI���#21}�d�w~�ܪ��T�wY�c;��X�u�M�HͿ3܍��k?� ~���?&��wWU�`� �vһ�WbºnݧVS��bE�.�>X����1�v����ͨ��X��c��~ A@�Tl����Մ�3��s��7Q��c%p!K�D~U\�m}���fd�Xm�	�$sNȼ�8T�n��t��,Hݬo#n�j/껳2I���gu�p�1�$�Xi5��2����ܯ�,e?Q��Z��G�*�Ƿ^1cK ƍ���6�6��ݱ9�$�m��8��r�5'�\q����n�uf��=γ�� ����5a5L��s��7Q��c%p!K�Dvs�#n�*�7�č���6�6����3$��/Q��mF���_��&��5�-��mj5Т�D��H�<�3̓����e�>����w��l���ֶK��v�@�D@a�k����9���8�,I�kD��0`�ѭ0�����kk˛]�Á3AG �&�f�������.lH؊e4I�+����t%��9�\N�秙��ӄ�`m��s�B]�u���'V�x�ֳ\�,H�S1H�$�5 ���:,:�
I�.�贆��Ӌ)1$	*ة�� t�`�]}��[���Ѭ�p[@                 &*tȺ�˰�B��5 =�c!��}���d��URzU	� m�ֳm6YcV��R�t�Ka�p�ɑ[ m�å��v�[��;[c�����*�vV�핰`E����ƪ��j��л�9+��n�kv���nj+��C۝T��e�xҜ�������ۣ�a��r�Ŧ^��P�T�]�f]���B�m���и��Y�ж�}#�t�Mr�sֲ��C�PFw kg��Kv�����9av%�)��m��Ev� *�j]���b9tm\�~~z��=v5�vס���{3�u�vst=�y�*��Z�8�<(��t�a���uu;etr����
h�]�������ٲ6x���,����Y�)�=���u-�7n��	��r�:,v�۴㝆�v���ED�Sٗ��N�RIx���+u�]�:�"�lq��W�q���E�m�^y	5�j7d0���T%����ӹ�j�ƕ�]n�k{�`kB��T�_@:@�^=��O$;Qǜ>݂�m>|ꋿ   ��٬�6Zw:Bj�@Z�@�d��ɳ�ۓ�KڲXM���-���k�X��Dj���$�85�֡7W+�h���u����s����d{1�k�g-��v�n�����{ޝ'��dxӘ+�v�*y�eV��a$ņ���{�ˌn��r��8�mG�1j6��<bǈX���X�!�l�dE�{M�LCo�Ds5�Q���]��0��m���l�Z����#����cO=f�t��ݻ-������`�_|�wȾ�׽�%W��� X��_^#	 ��"@�ڏw��/���{z���%�"=γ";z����T����Rk9�e�$G����`L���Ũ۬[�"H�n�G-2�8��z�����T��ҫ����w{��wST����@43�̈ˏā[S<��Y��ϼ�����(�`���|�'�?xp!K��G��H��X�[�)��
�;�� �ͼ��n꼖H�p$�	��u�Z�'�^�����f�l�\��,L@�?_��F�Ũ��ܯ��c��Ũ�u��!��� ƍ���6�
 8@`�
#���(�;}F��NZjŋ|�#ݬڍ��{�$ab������,�8�b�kE��=�Ӯ#3��s���o~����B�L��q����U�1��$m�7����Qv��Ȝb��ͨ��Z��Y@�>���m�-F?��p|0 ����Y$   ��^*�l
D�xBTt[k8��n&��҃�c���d�lu�;��K4�3AcRv��`�'��ьN�{=u%��z���[�.�E�hqYs^�:�M��y�y�z��:w�_w{߿����{u#uۓ�[Z�$����)߫�u���F�X��;�U!a�w���G�3"�4;��q��Z����̈��;�֫ub���=�wq�dg���h�I.��G3�w�w������}ܕ��)�$��f��vc7V�NZ��� z���.�mG֮���c�u� �[7���[����H�u��>&��#{C���:\;�c���.��㪤,SGwX�<��̈��v+�v�����ҷez����ucu�i�I�
��u�gu�p�(N�En�]R=��b<���^�����I.��cD
Uld�@!�C����̱L1aRG=�w��R#�z�۰�/ߑ�s6��X���Rd�<�	,i���v��==n9U���b�9��qn�I�"7(O?*	���C��$G�1u�V:�b�4su��<�gusz����mpB 	�̈\�= �:z_#;�֫ub���s��Z���RD�P)#S���x�NZ	-Eq�K^�W�i��Y����ߑ��J�A�1ďZ��>��W�;"�U+v��"<�3�n���⫪v)#���#��! H��	��0�q��uޏ}Ǟ��{Q���Вy�s����  �η����T%��Ʃ�ȓ
�kB� ��C��D���ٶ���A.q�{v�µ��5ѷ/���r��eW���W���n6�92rB��<��Z�eE�uz�Y����}����R763r��:����Ff؎%27��#�X�G��fD{3)���-�	�c;��u��kU��h絞�<�cu��1<,$�L����ߑ��O��1� I#ֱ���f����~O�����7��3����V�]�~��z�~�~~#�c��ɘ�ďZ�$p @I ������йS��$�ݾ�c#��.�v���,4�n��G��!5"=���T�U��"0w=fDy#��j��T�XLܻDX�9���˘͹[J�[�V.��g���K#ϧ�h��.��@��H��b��,SXI#��o!;���!���,�b3� #�h��b��'A����a�m�4�����4��pS�t!"h�����ٵu �i�2B7�%�i:�Ѹ�.)�!���i�(�a#q�"`�'�#��� P���*�dEа&a�rz
DXS�����C�ت����!��P�>�4	��v�1P� z=��N^s�m�Q�{�M]��$E��B��H���f81#�ߙ�F�b�h�z9�4��:�{/3�;�\����R�a&��_�9���(\�r�ʍ�!4~�o"�f�}=S	5�,�����y��2ǐH��Z��6��XАx�HBb�v*|�On�4>�a*]?Ds1�{�|8�~�b�����n5�ղY�4v�xL.�ئ��#$c���E��ުnX"if<HW���u��ԕg'Y�$�dg�����7�޼	����@jD}�1".F.��u��,SGwX�"�Yݾ}y׻�|i~�@  ZtV5�e��Z�y���N��VƮ�>n�^v:��,v�U�H����	T���W�<&-v��[W[���n��n\���;�W݇��=X���w{�������/���:6X�'�n��Evng�n�(y1�"��Ⱦ�'��b��Xv��H�q�cu@ 9�������.��G3��^���c@�#mcyk6�owf$�Hb��ͨ��}����f,i��Ey�����5�6��Ʊ�Gֳ���Ũϲ���jE<>ː�m ���
����y�>c�>h�~C5��x��X�E��ˇ�ی4�T��7Q}�}������
[�j�����F9���ӿ��pRj�+aU6u�֭^��������<~G3�����ܺ��*H�����ک2�vbN4�/Q{�	 �$��Q%�'X�]x��	#��F�b�g�u�M�2OQ��-E�^���~�q ]tGN��!���g�=t��['Rlu�=������y��Q����7V,�����y�]۫�3��{���������$�dG3�H�Q|<@= \�v,��MU�I5���}�nFdG�y�<��V���ٸ�{Z�CV,6�4m!K�D^c2(hI�T��N���=���;��ꂇ$��j���|2#���"7#Z�cUHX���5$c<��̈�{��&�R���E��F�b���F|B��w�I$�I$� 9���-L`�"��Y�c��	HGR��aE*^,q��7n6�N֓v�mS�U��Yc	̗/(��=a�{�\��:Y�n9��u��aT��I�� �I%ʪ�E-�J[���;a�2d��v��iԽ7�Y��i�v��ڦ{#=�ve1����x�|	R��bD^��r馪¤��܋��j6��bNcA/Q}�ڍ�����M�In��Gw�G���zӠ!�۩uF����YF�lS�uM�v�ի��dG3��Ϲ��kY�6Z��}���R���!?�Q ���������y���NU*�Q{�ڍ�Ϯ�c�$Xϭgyy�#<����|������c"�X�9�"�VԒ�,42�\�v��7v'!p��$Ln�2.q�̕�:���1'C���ͨ��>�_L�1#���!�A��EP Ăm8�"/jc�j�ӥ�"<�1��7Y�{Z�I����;��u��~ 	��^�v�4���Y�(�7\u�z�u�0�$���w�n���[n���3���w����~�ģ�J�L��1��ZǪ�3́bG��o#�X�#0��D�q$G��u�1��^xYN�I.	�q��y���9%��6��j�ܒƘ6����0[���mغi�IH�b<���oո�S��.�y���<�g��I��SC��{���Y�oz����| 	��{�fDy��{�m����n��H^�r!"?��:�*��(�P#��P�pb~�����G��?טu�{?~�������� /U"��zmPq�\�]B���ϟ�4k�:O��t���~ېy���W<��{��{k��]j�D~6��A�7���F�}�}o7Т*�0�矋��?0�i��P�#�T��������G���|�����������DT��������pq�'����?���&����Ӿ�I�?o�1��5��_�����
��?��bE d�@B$P!P�@E e�@U�QQ5 .�Et_��9u�g��k���v�����������C���~������@�����~�C��A�?3��/�������x���~S�O���x~�0�[��_����~?��5�������?����O��� �����?o��MO���<���΂O� *�~G��"���O����&��ᇯ��g��4�D���j�vh����� ��:���ި4��q�XǏI���"������"����x?���C�����?��O�����ve�}�G����S���?w�:0 �r?���������}�?��?��������?��f�@_������?S���?/|����1���>�P	�s��>Y�������?�ػ���p�6�g�C""��`��_�>�����>�fh�y�.�>�wI��?2$<�:��]��B@�Lb