BZh91AY&SY�(���_�pp��b� ����ak� (���P ��) U��QP������� 
)*�JI*�)J���@��R �$A@ �B�  (
H�� �@( �� @ 	(��( $Q�   ,
@ �P�(b }��b;�S��0q� {ޔ���K�@�1 � (�}5�	5� R�ZUfk�T� �CJ���R��
&�j���U14�CJ�m� Ӊ���    }� @  
�(��� �}5�����yiO\��n ������1w4�dWs�]�0��@u*��cc��o0����8 ���!�2轻�����=}��\�}z_|��˞Ξ[�e\ ���    �(e� �=���{�{3�Ҿ۞��� ���˺ڷ9�lq�u�̣ �9o{r^{ z�`���� ����t�{����7��� ���a����\Z�NAǀ�|    �I@Q�� }�I��7<�绔90=���
��@����X>V{p7z ���0�8����Eɡy�>�:w�J����<��q�ڗ6��y���L�Kv;�s�]/y�� >��@ � Q�E }�>�����W=�/6�5G� �c��ϡ�\�rһ��zF �\���Zq��  7��u�x���@�=;����:bw 
{ǣs��s�}O�}�'��       􉩶�J�` M0    ��ԕ* @@4hh E?�U*F      ت����  �  �?��)���TM d�h�	TOSS�&�`�  yC'ȟ������_�������ﾎ���{��**����� ���DT�TU_����@�
��� �����_�Ȫ*����*(������_���7VsP�%��A��ba	BP��P�M$x��	BR�a��m��C��&�H�0���#@d8	�a��jC2QD��{�N����05u��<�0r`���a97��k����Z;2��%��9٠�jv���S)]	��$j���]�Uw^�y&&N/3�(MBw.�؆C���E:��՘xAb��s��vk{��/BN��j8��P�7�B��T�h�E�.�2p��8c��]l��3h6mٜ�ё&�;��g�Ӥԇ(cElk	��%)I�U�ĴRZ�;ɞ�\�G��s1;�FP�ł�:R�x��)�=q{}�­Z6���ۼ�#�Y�v���+9j�<�ʿL���Vګ�u"M���ѫ ��1�'#N6�f�4F4��8��b�6i��r*(�bCHMAʢ:��	!�!������0�V��`�H�j���Er�ğ3���.Z��� ��2C;�@��C20�\��0"ˮn���t:\���9h�u�^6/r�m���]m�)̒8��X��
��m�;��I��SLL5=�发YJ	&��p����J�JPs&F=�22�6�͜-�J4a��� v'#a�i��*4dky��������Ĵ���ӽ܍��'3C���>:�4e�l�ﾇp��b��]o�u��'������s���vqv���N�N���s��w;�Y;ξLZ�	`�>�W�![�룮��w�q�9�Ҹ���ɺ�ꜘ��O#x�C��ȉ7w�WV�Q�1����A�����`�%L73�j��306���:��;�&��÷W�2&��<9��`t��p�9bn{�&��v'D��s � ��ɦ$*V�+),�"��m��F����}�z���$��S�N���i	�I2Sm��!��Z�B�Rb)�x�[�|�g$���h|�$W`�)10�z5V�X�MF���-�rR����䆼�����ӳ�ב�;�!(rwY	BP�%	����,��dt���:<=��k9��2�8F�*�8��kq�[��d�d��&����:�e1d�K�"~bYײsYb�	��`]Bw	�'R&Bw���՚n�����?:h�˂&OB����]���	��N]s��ƪ%�$�
�jP�&BP��yt�y�;�'���N�[Ow�A���V�.FнB��(��H�^��C����/uh����<��JFX�`�5�NBd���GI�p��a���Qu���U��W!�z��:[�Eԅ������Ӣ���NbBwe4�jLL�H���f���2Xv�qy�rd%'d�A�^`kw}����0�u.9	Ho �4owy]�7�Y���4�	A��3ս=��'Qo\���C�Q�v����Y���Rx�Z�u�CYc���C[h���o�F�79���@hE.H�V�R�J��Χ,^����:�L�&L5ks��tXaĜ'F�sFНBf�6��;��I���q��n	�H��J!!E��[V���;���P���i7��%�bu)K�t�*�{�W�N�D�$�#�o.�|����o��;zN��ut�������	H�J�5q�?w"9��yǋ���x1Z�.�E IO��P���.�:6��ظ�fb�z��hS����y8�fq	�.�E�$�P&����N0gDRwf݆�\�����^������S��5G(;�<Ԙ���x'!%�qtÖ�NN��5�.BPf�����npĝ@�BPOdR�٫F���³BP���u���q]��f�N�Ih�!"��1۬����X����uu�{ѷP`��]�'%�#Aǽ���1��F�����V�Ru�:\�e�a�ӑ���8w���L�&w7wX��(6�CYd��|��E�H��c�j2�*xfsi`��K�0��!"��(����F*u	�c��,s�#� �3.��{՝/�Z�T&��u	�L�'[qz�����:*��5t�CУgoG��,tfdbtnC��H����g'���|M����rd���s2u�n�N�����˱(JItK��M�	F���S�Z�$��>�3�X�9���T�R�%�i�(N�(Mfi&,��(MK��Ų�0((����3b�DD�5NRv�2��D��Ƚ��)�(F�P�v��L�99h7��{5��F2`�&%h�T��=DQ�Iq���YO˙����QN��%	By�%'!)�� �0��BQ-I���(v	X:u�k!:��%	m��m�t���f��w7���_���8Ì�h3f��h�7�dR	J҂�HN�A�M
��~�g���"��+H���kQ3/���h]��,�Zs�ư�$I�u%#�f�9����gIզpXp��.BS�I���l���^w�{و�5�����c���4�7�����-e���%	�`�hv'����Yb��dU;�6:H����� :�3T:��㓁9b��0�SW�)�����ђ�A$�k�j���(J�N�̪����V���V�S<�k#LMڟ�������G`d%`�ԛ�������[����F3X����x:�cXj0c!�2qr���lj���S�D8R�Y�g�4f��Gv���J0 ���%óY�2��6�.9h�ѷ��������7�&�4���{8��a⩧�����K����pY��e5Bk�i(1&��BVqx�)y>ԦZo8�EA)N�Q4��/����	OnP]�An��-`hr�1�l1uZ�ߗ�����U���+X�������Ԅ���6٣|��}	��+�8U:�k;��Dƭe�����l9bHfB{�������e:bi&W�om��h�M-v�ʳg�7'!,to�NXi2q5γ�_2�W�:�8վ5�I�K)ASI�V�@wR`S�٩q�Hy��@]V9��QCE,��-'hN��CPNJ�%�b@�����ї��ZC@4�@��"���(������	�㓁>kbP��w���6�]o\�Lt���"���iݩ���ʧ�K�GP�ړ���jj(���6U�(��(1�`Q��双5ִrZ���;���q�|ER3�F�in���r5Bt*�D��0��R�P%!��rl�-�����5�Q���Uݫ������/M�ъv�y�Ve�;�����R�����J۸Os��2���|���7a��z�Qq_0��WQ��-X�kcJr�	4����Ms.��H�����9�]��.Z=/c[d�v'��`c:uP�� ĺ��{�t��0jpl�g���o���'M�����^�֠9���<�����2���3�0J5��y:�I��&A�d�k02c�2����[
�X^;k#��h���cGrcXڃ���Խ:� 0ܸ���ĕ�k��\��!g��_ �4'���p꬗\���m�	:�{<�W�<:|��������v!���}\�b`]I���6�Z��@QQ}p/
uek�I����:J7KPd'��K��%!�&&BP��rC31cq�r#�:ܹ]��-����h����"Z痺�\��.��媲��pJ%H"ʇ�pd����3�^V�P�\�<D�LIѣ.�ueW��p���.Ύ&�)|r\s�R��ē)���Xz�-�Y
��(>&�����y�0x����(IԑԘ����Hw�	NY	p�4fEW���t߮�O����Rʜ��S��aPL]iH�T�wU�r�
�&]bMz���r�6n�D���&u.���u�������N����]9t�4�i4%
i���W��S3�\s������3�%� �L5��A�q�&��Nf	�v:T)ʔ�A�M�t�bqB�u���WI��)z��e�q�JˆB{['ZN��4S��Bxf	C�e��A��J�(JbE2V�,�/8�(�̤�P�T�P�D��F^ALQ�����RTjU��ݝl�C2LN�0�qr0����U5%�Z���K)��[h��IpM�6� c>N�,��[ӵ��A�	R��l��K�T
���R㐚��P���z���:�$3�Oa(Ou�r��lC�D�F�2tY`A���`����dh�W��F�4;���=��`�3���w	A�*��8NBP�'Y�Z6��ݺ���`�u:��%	hƁbn��R���块o
M�����D�aw�w٣w�۪��8;\�����̓,��C2ͥ��Q"A�ɅНيv,��%*;h2�`Y	X�7�&���ЗYlãs���ij�C�΂]�EW*"�(�Ȯ
]�P�2M��:�'K��r^���!2���bL\ۺzSci���SSI#>f!$�&��#2r�"d���N��23�3;�N:��o�IOA�V$���N��*^n x�W������fb�<O��� � �   �$��   � �2(0m�   	�  �h  ��h   � 	 dڛ`�ց � 8XH� �  Jl��6�l���]�gnP.��xB1�v���TC�2�;Ķ�'@$�$��Q��-�底j�tN�[״��ŵ�l� -��S�u���.��T�+h�S6A0�m) 5W[m:%Z�uN����"c�!i���y��>8-A�dn�L�֝0�q���ԝ�FM��n��L�ܭ�ȸ`3�m�e�׭�ꂧ�8���W�Ku
��-ڎV�
�פa���ٜQj�+Gh��ں�:��� r��U*���+��EU�t�M1\$�U��Ml�nv��]�6np���UtѸ`'tN.sG��[�<m<�T����[Wb�mVQn�E�8AL�P6�2�����	4g2)����PC�9
�텶�cqӭ���96��H[[l*��� K&��I�^7A�Av�p��UU\p�I"�8���d���}+][�ӳ�-�I9ɥ`  m�o��I�a��M�$�.�Kd��   I�����[U�\8 Hm��ۙ��jض�  6��6�	���[%�PM��$!�
�3�H ���l��Tӹµ�3N�H�8I���%�-� p����������  m�WI&���v���ֆ�p�m�H m���n�wJd��v�Ү��SJ��Vy��V��|�v���������kjt捲����&�[�E�  F7�   [d$m �N�%���	�m��HE�l����qm ������m�a�ܥ�n�H	  �M�m    �����Ŵ8 -��V��l��C�e۲S�U@`�*�;�dxp������+�Lf�͒����V�U�`� m���ڸ�m�I�  �uK�j�oUU*ݷf�Ve9�D�ru��t�H<a��5�tc��oc7m.6��l�	��-��`��qi���l�m��l���mu��k@ 2]�lm�i;` ��=���� j�eZکy:��T���� �탭��f�z��`���D��HA�m�hղII�[@�m p-� m��   	   6�5��� ��;h�n� ���6�b���@$l���m��m [@   �l 9m�^��	 m  6�8h e�m��` �E[C��� H  E5@xi@j�����m�m$ 8���a �u�  m[  s��&�h�iU	�h�	yj�\� ����r�l�U [m���$��hl�iC�M����H[zpĀY�m�ϙ�^�������H��Y��`-����n�k�@���-M%8Hm��V�����K]6�:@�8������UZ�m:)�@�9��z���I�gZݶm� j�-M�YG�Hm�[���� Kh$��-�q���m�f�!C��V����Am�m�H	 [v����A ����8����ɐ[Am'5�l�&��|@   �$���-�$Hh���� fQ�`8 8�[@�` m�p ��IV-���6��EH 8  ��[d�   �xoZdP��m�l �5l� ��5�[Im� 6٭u�f�    fؐ�k[�h����8 � ���i$�,��m��LI�5�  ��ݤ��q��pQn� m:V�H�����sh�V�Tpm*�$�.հ6�Rgm� B��[d���Q�6݉ I#m�h�v Ζ�6��6��2@kn����غmm ׮���y�OJ�lm� Xa ��ā �mt��'EUj�ȻJ�fvՀ-�l 6ٶ��̐mY�6Kmm��ٶ�CUp�NӦ �MPnKl��;
	$��Y��m-��� ց��\  ]6�۶�a�ȷ,� h���Yw����Ν*��<��-T�UN-�p �Im�k@#��%�[Ev��;'.P�c��P�Z��� J�+�U[���\U*��=j�W�����akF���#V�S�.�Ӓ
��Eum��U�PUڪ�8�*��m��	m� �/L����&�N�K�H��TVh�UV� �j�K+U���i;���nhڪ����n�E�[u��ȲIu���m���0 9Ҵ��ݛn mg6�T�Zظ��2Ѷ�s�U��#wl�m�e�ষ뒳kh   ��n�0�^�e�}l�zսۦ����,�&Cj�ٵ�8K
��l��6����@�m�Uj��=��U�@iW����Zr��n	�Z�� ej�B�ct����m�T�[��nʺ.ڕ` *�������[PV����h
� �W7L�:ؖ�0��UX���WU�,��ܨN�UU+���ŵ�. �j�@    �i��m�(h6����6�Ͷ��֝&�m�p�i�ۋhm�N$ ZoǸz�u�� � l���8Zl4P  $l ���tE� �M��ݶ'I��`6�d�m ��[pև\.��f�ֆ۳m�89m
��rÔ��\J��ض�i�HM���B۹����#�  -���H   m 6ۋl��i�i�[V��]�~6ܶ���� m��a�@� ,6Z��������KUKt�UJ�l�EB@�`   $6��� 	 p � #ͧU�����|�@G 	lh�a��-� m�[rvؐD�����v�]���bFHm�   �7m�m�c��M�m���v��e�J�[N ֶ�8�V�U@T�jU8()]��j��ݖ��R��UV�ЭEC�Zꪭ �m� ���t�m��-�^�ȍ����[v���Ò6�g	cY$���`ٗ�H�����>��(M�c�8p6�a�[R � ېk���,L���2ãd�s�T�,��R��J��Ҫ�T���|��mɐ���U�j���*� ��M$N�l�Pl6� C����kş]ȹ��|���bv�� �\Ua�Rgv�ŝ��Tz����d�]�z��Yf�@gC��;-�Vq�8��j�t�zUZ���!cB�nk�`�Ͷ, QP�j��B�jSr�0� Xam@��m�l�m�-�iW Y`�� 8-m�āz��`�gGձt�:j� �  �l� m3��Ϡ������'�z�#k39���� [Ru�R    m�m ����$ �` ��I�m�m�	      ���6�m���i.�m�6� ~�  �/J6ݰ6Ām&ʔ�j�T
/5V6�u       H  Ò6�m�۴�F�*�Ëh׫[@�l������`�dk�l ���m����'N �m��` �h  �e 8   ��Ku��[y��"�  mKA m���m�  ��I   m� p e�� mZl  � ��  ��a��h mְٶ  [E�  ݺ��uM�j�۲Zf^evUG-UUUm\u��Pz���	]�ԅ.�k[@ �m�Xc�J�  	 �Kk�D�KU*�UUJ��I�kn9a�zRC "@���& -��#��  �Yb�f`X���"��B�v  [L�m&�D���X�z��[VК�^�)y�Ui"n�6��     XI��p	m�����& �I�m�e���m!M�0�8 u5�Cj�δm�m�\���
�UR�UP�R� �;2�ʚ	cfڪ���M\l�kh����d�Z�s�*���]������aGV�Y����:͞�nR�ug��e�ٻ ����k��������ӀH�&��ץ�&�F� ��ꪪ�H@4�*����[@� $ �    �m��-�m� pkM���V�(�k�,3m��N�6ذ��m�-��    Hm�  -�i7  l�   �*.��B�����`       n�@ ������l *F�2 @  �����uV j�0ְ� ��� �H�wH���mUJ�UUJ�J�@   [Ki��-�Ɠm�6� �����d'�VvZ��X����[T�ԫ��e���6�` �d�������Kj@ 6��A�e]��ET��*���͒ �v��   m���m�   [@D�O��W�?� UW����w���YHeV�%�`e"O�)����Tڧ���: ��Ҡ�G�C��&�<`N� � �� 	t 	��:$����9�hTQ�U4 @ �G�R����M=�&����bcg�D�P���"������O��DN�P�� ���-�c�!���@' <] ���������@z
x�w�C�=�P}GA�E{W�  	��A�%�}$ ��@��]� ����h��x
���b(�h |��ACb��L�6I� ;p�"�!�㊽ l�N�<{N *�t���9�بGA (8(�"H�P<�S}�&E�jߨ�!���P�^mK���@%X%�0���v�Ҁ'���4��.���МEѥ�g<At9��)� ��H��N<�{�Q�E⏈�
z*t � ��D5�_��EW���o���G���	$�Z(�(`���b�
"$�M�Bb�$4�+BH��3[�5ov�{��6_n�����$��h[i��u���m;B���'�'U�u���F��U��1�+�[3&Ӆ�nԂ�͚�r�v��/ke���N��Av�RI�uѵD��5�'m^Xh��y06�vr,3�-�]��,sx��
(����ʛ\p����D�l\�41�fz&D$sl��y-�h8�lշS�oXv\p�um��j��m��N@�x$����s�ZU��kT�n��[���gfv�Z3����x*���fy���AF�b��j-�#m$��i���\]�H&�8%tT�t$Xԑ\l�Ec<��mۃ�[9��W\��^��#��dҽYݸ��u��L�X���h�q�{)U�a�Ъ��1-U�����[ae^�U�(�k��6s6�2ЃRYA+Q9vQ�d������GZ-R���l�Qgd��� �Tڱ�e��iU�6���qқ�F�j�S���A<��(i� ���-���r�YI�L �5���:YV���V&�MGU͜[t��Xh�Ή
��8�>_bH�\`+'s���ckv�Ӟ-6P��'��<g�ѲcQ�������`x)U��۬�5�먖��(,n��Y��^Ҷky�k&����C6p�+h8R�ykju
�"Z#M-դ�Ԓ�ŧ@� �j�NѰ�n;q۴��ѩ�g8��=3�T����Oxc�秚m^{d���m��ْ;u���:{z�y��X�v�ƹm:Vڭ� �Z�
�A�1=2�c;`Tڪ��jJ��VӤ���w�[�j��Hm=+-,�f�P]�Kq��ic��UHu� �N��Bk(ʨL���*mp@�EU]�Ҹ�x�C��jr�A������gkCU������=�:�d�����:�������V��.`.	��
]n�� iV�������I�M��bC�&��l9�e�UUQ���5�X	U㣴��R�邑݆qq��hw5�i�e]�v�m@@T K�ww����E�O�8Z �T"V�P�U�/|ؘ
'������O8�����]u���ֵf�D�uv��gVK���-���Ʈܫ�=c]��N��ӷm��7e��v��!�̅��lv�n��8�=��rj���!�mN*�ݙx8ˎ�m�H�k�l�&КT���5�ܐ��;nM]j�d�NY��A���1u�Z��W�l�R�r�薨��n��3�  ��N�5v�ڐ��U��[�5��uT�:���{�{��a�(�.v��|�U�J @�(����U��!��D��7.���q`~�3�?��� ����]+m�m;t�Z�<��3�T�
���b�=����{q`�y-#���wv�˘=�� ����;�n,ϻ� �=h��q]۵$�Xwצ�{q`}ݘ	Q�n��7�LW��)-�q۹-�����ـs۸�������|���l�d1v��	��gm�n���ʰ��7�]]�z{gus��{��4�t�4�w�}ݘ=�� ��k�=�n, ����i�-�����%Um$"�)�	-����7y�{�r�;�����v`��l�#jEl��ݛ� ����?n���� �li��C�ar��{q`}ݘ7wݞ׀k�ٶډ���v�[.Z�;��x��ݵ�;ٺ�{ۋ ���G�[ͨz)��3�ki�wm��덭Н��nơP������p��.�=v�B��swq`��x��ŀw���y�F؝����K��s�u����Ok�9���o�����K.K�U�{Õuߛ��p�aG\�8��(��!ʄ �2)�=�sY�p�^{��������6ի���X;�� ����9�^���ŀ�[ ��n(�(�wf��ŀs��0{ۋ �}z`���R&�V:V�J�J���)?��˶���&^:�>�Xۍy��>�F	ۗ�!ە��jK�� ��0{ۋ �}z`���i!#��ڡ6�6`������9���wۋ ��m��Ӷ��C�X����ݕ�o����e`�=B���
�6�M��{Õuߞ��^y�9]��~$p: pQ=�ֻ��^�U��2�N�컶� ߽�X����7�^�7w�%IR^��C�9)��W;q�������'ua�s�;�]Um��/>���y:�on�WNݕum&�cMց��+ ߼��7���U~�{�V zJG�u%N������y�owe`����ŀ�[�Z��N�hwf��ŀs��0{ۋ �}z`��I5\�l��'%����w��X;�� �q`��~Z����X;� ｸ���>8w�`�L��BIZ@�!(�*�� ⁩Q�H�#�w�.��4� ���R�s��B�	�0��[}}VF��H���,Y{�q��h�)��{Bqd+j�ԯ+'�[f�s��,G���� Wg�][Cr���1ƶx�WX]C��w0a;�φ����;�w.����Wlb۵�ݷ�jnN��Z�q�����..k*���;np�`�`���,��pU�M��l#ї�rr���ml��p0u��=	0�a���7��e^�:8�w.&Mv���<�<�Y�Z�fWy�l�5���·�q �L�Su�u�x�Y��4���on��vX��{�0�vV�y�}�vV {��9��e�H�]ܻ0{w~�M�����镀o�|`�τ�N鶝Z�� ߼��>��+ ߼��7���;�&+Nli��l�[�`}I�*HI{�m`{�0�>0�ό �u#��	S�+m�u�o��`�|`��^�{q`%�G��nԂ�#��ֺn6�G���ns�\�|�z�s��2x���;����Wc�ڻ�wb��Z�0�{��{q`��x�h�MW##�	��ʮ����׈Pv�*��+ꨕ,�o�� �f��9�0lm�����aM�m�{ݕ�{��X�������VͶ�N���n;e�X��yȰ�8`��x��e`�=B�j�;I��X���Kӥ�n�� �f��7Eq����K�9R��;2*q���Ĉ�ۧ��;uۂ��ո�Z}rlvԷq]۴�`w�x�ۋ �f��7f��7�LV���R�h�5l�;���UU$w�E�I}���y�T)Ŭp�K��k �f��5��0�Ue*[[T���e�]�o�q`�5�c�&팻��k�`�^��ۋ �f���F�j���Kr����o}��vn�_}� �V޸�j���K�Yw ���7;�	�����:9��r��'=s۵�;�s�\��wf����=ٺ�}�������u�J�6�ݴ�C�X����~�IN��zs���������+��ci[tյ�I}�y�n�q`��x<���إ����������N�X��倫�}UUB)R�W�7��b��ƚ�ݲYnY�n�q`��x������o�����v�;wF&��W l��[y�o#z�,u�j��&��<8y����F���s�u�����צ��ŀ4Z��Z�lM����n�kϗJ��B�@�����`}�b�9��|Ѥ���ƣ�ԗ-���Lwۋ ���7g����g��K�8�ـswq`��x�=� �z`~[6�Q;�r;v�㖰zn�ޞ׀w޽0n�,UVP�I�][�|����U^*�Vhs!{,z�L�o�����u8g����K΍Dk&���6AA��H���Y�3%�6tV+8�e�`
�#m�[���w1]��S˲��8���;vϗv��uE\a�eX�n\��㌻��v�u����q�Cl\�g��h��	��I�̙�;��Ԏ	����tV�L
v�#p嶶�`�6����?���/�g>�o�3ձ�u�r�(�r�����,���5�mG���hk���{�m!4,8w��>���vV���o�0�U�퍶RV����X�vV��� =�m����"���%���@���t��.��G31�@�7��~�
qkE�;�\���zn� 罷�wwq`�� t�j�Yv�F��!��}�x�ߪ�$��>�X�}����N2����B�e�n�7\ ,!ӥn�;W[+l�v��=Ր�ʝ�����Z�wu���.{�i{������~u���5?�ݴ\V^/���-_"$ꐓ�$
�WV���ؽ��u����-�mݲ[���ۖ�{۸�w�+���7�iw���sDYaq��nK���\��qs}��=��\�TZ���+��2K��{wԩw���o�b��l�����u��+hvѱLp/[��v�ǉ�[^�7[{�����wumٸ##��)w"�V�˗|]�~���n���l�o�qt��S�Z,Q�r�ܵ^���?~�q����eo{�J+�C�E��;bn�˻ŧ��\�n���:IВ��
T�v��7��1�W��'7ѵC`I[�vm�=<:�E).t	��""j�w��0s1�iy�cAM*Bg�3�CWw�Ђt�vZ�A�T�� ��5���kfM4HFf�&�,ݰ�{��*!@н�GL�<PtD1�0�	tj���h"�L���ֵ���k �0G{� �ӂ ��L� �= ��8@��{��H����~z 4�ԯ�a�ԧ�{�"R
]߷�U�U �F���'�9�{0��{��J���=JR����8�)I߾���J̿k߿k�R����m���(+�h������R
�߷�R����~��ԥ)�y��┥~����)O� ���F����涖�d���vJN�dݣn�m�ΐ��5�n�]�����v���t�Q�e��n���o{��y�߿pz��=�=�\R����~��ԠU.��bʤH){W��O�Yaq�w�k[��)J{�{���rR�Ͼ���ԥ)��p┥'~����)N����[�����.eR
�
�����)N���R����~��ԥ)���ʤH)o|���]�A[�KǗ���)Jw��p┥'~����)Os�~��$: �QH� �A`���|BD���#�qY}�ث�R
���(&O�,Q�%��x�)I߾���JB}�߶߾��%U���R��ɔyI'��r)i��w\V����s��u��ku�� ܻR�p�����f�f�������?JR����)JP��}��R���~��);�߾��)UHߚ>$��#��R��ʤHw}��R��{�8�)I߾���Jy�ƻ�F�\�s�i$BH��LWs5�pz��?{��qJR��}��R���k߳�R�=���pz��=�O���ݲ[�ݫ�r�R
]���U©'�k߳�R�=���pz��>�߹�*�/j��'�&��qܻ���H*��׿g�(~����)J}�s�P4�{��pz��<DS���h��a�pF,٪�,=����U6�k��+N�tҏn�z�3r�.�m���p�݁\�l��m�����j���=��M�� Ƿm�'Z۱�ǀLzܮ��y���H*7�۳U@��s(�����+q�N���m�#�����7`���`���v����,WL�%j��L��j-N��pb7-ќ�}��UYZvYy��Y�K>�q�ݵ�m3��n㞵�n{F�E5�Z��֍bM����*m��s�N��{���n�翿~��)J}�p┥'�����"�u��U �AK{��G��R
��^o\�8=JR�y��8�)I�����JS����)J���=JR����Q}b��wr�U �AK�߾�\*�)�y��┥�}���)O<��iR
_{⏧��#�Y!��U©��}�)JP���}��R���~��)JO���=JR��a�k5���U��ӽkz┥�}���)N���R����}��ԥ)�y��┥'�����)�ﮉ-�ݴ��{1���ۭ��":M�t���Ӄ�63���_6wLm=|޵�pz��;�߸qJR��}��R��y�k����%({���R���������Kq۵p�ZʤH)s�߱WQ���x��9)�}��qJR����}��R���~��?f)I秿�5�zѭ۫�ܹr�p�AT����*�U U����� ���{����%)?}��ث�R
��}d�-Ȯ�ࣻ���(~����)Jw�p┥'�����)K�=�|R�����/��Ƶ�޷����pz��;�߸qJR��}��R��ߞ��)JP���}��R�����yQs��-���b	�(m�M����X�3q��i�z{gus��'s��OkrZ�o{޶qJR��}��R��ߞ��)JP���}��R���~��)JO���������\D.�p�AT��~��T��}���)N���R����~�p�AT����s�.A�ݱY%�U*R��>��R��~{�)Of�$b
C�!�N�8R}�}��R�G�~��AT�W>��� �[����R��~{�)JR}�}��R���߷�)J���=JR�gǺ�y��Kv�ڸG-eR
�����U©��~��({���R��~oز�R
^�}���R˷��;���[��ɷqѺ;	;�z�ڕa��t�v��c��M�.;�aq��\���U �G}�^U"R��>��R��~{�R��}��b�H*�|۟Hӷ"������R�>���pz�iN���R����~��ԥ)�y���
R����_n�oQ�F�y����ԥ)߾�ÊR��{��pz��;�}�\R���߾��©R7��3�dvIww-eR
J��{��pz��;�^��R���Ͼ��ԥ���((����F(�� eh�Qc�;{�{�ޜR����'3߭lַ�����|�)N�׿g�)_|��=JR����8�)I�����J�����?
7:���t�r\�$0�۵�vb5��q�Ӎ��T���v�FG/]�~?�v����3z�qJR��~���R���~��)JO>��'R����k�ER\�m�����l.+˒�p�@�~}�+JRy��}��R���߷����g�}�Y��s��'ԑUTҥQ�Z�l┥'�{���)K�=�|R�ҹ�����ԥ)��~��)JN�^���q�,.7.չx��RTww��JR��>��R��~��)B�}���*�T��o�&�;�[���ࣻ���(~����)@~	<���R����߿pz��.����JR��H��~��,���/!۪ʑ���2�8#���w��o�͝$�����Ӯ�%�G
�����u�FY�e�c��L���-2q9B��W����u�M Nb�\�)�W�ݣ�����=� �ޜ��嵜��=n��M�ƹ#���,�[�%�ӣ��y�c�&v�Y&�ɔ�mO@v49�����j���Kd�w=�����C���+�Ѣ�8�u���Jn��wω������|{q��Χڷs�t�ɏY0��vܻuϹ�\R��:�n3���Ϝo��;�5�o����%3�s�)JR}�}��R���߷�iJ���=JR�牋�4U��%�r�U �AK�߾�\��*(�H�^}���JR����~��)Jw�pഥ'�}9�}kf����o{��)J]���┥�}���)N���R����~��ԥ)w�O�mH�[��$�ʤH}���JS�}���)<�߾��)J]���R\�m�����l.+˒�ԥ)߾�ÊR��{��pz��.����JR��>��R��{��Z��GP��{2<�Î��� �u҆�\��r^����'nwm����v[�{�JR}�}��R���߷�)J���=JR����8�)I߇�ٯ����aq�wc���U �Z��LIz��Uӱ/�h�B�A�p6��A|��R��}��)N���R����~���U �[�	�ℸ���%�ʤ
P���}��R���~��)��@d�{���R����ߵ�)JO=��/�e�j��/2�3p�AT����*�U"O<��=JR���~�)B~ !��߿pz��/ޔ~�~�w�v���޶qJR�Ͻ��R���k߳�R�>���pz��;�߸qJR����_kn���u�]l�j�ln-۞�>v��]�8-�����q�=��p�ü��8�ے����v��<��qJR��>��R��{�)JRy��}��R�����kxkFa�ٖo5�qJR��>��Q� C%<���R����߿pz��=�=�\R*�*��m��"	݁q^\����R;�߸qJR�Ͻ��R���Gg%3=��┥�����)O~�>�a�[������U �AK�o�b�H)=�=�\R���Ͼ��ԥ)���ÊER
]�����v�XKn]�r�W
�����)JP���}��R���~��)JO���=JR�}�Y��ѯ�[��\�6 �v�\�����k.N��m��ZN�m^�� [w#���]̪AT�W���=JR����8�)I�����JP�ty�����Ou"P�j��i��<�pz��;�߸qJR��}��R�����)JP���}��R����W�N�ֳv���R����~��ԥ){�o�R�?y��pz��;�߸qJR����3�l����E��|�)K�=�|R���Ͼ��ԥ)���ÊP��$��$��J��� ��!bI$�H	)@�Z�ifYN�r�����I,�J1��y�K~�}��U �F���}%�#h�Aq��R�>���pz��;�߸qJR��}��R����k�R���{�٣6krhC�F����v67m;uI�S^�WSЅg�q�iR���;��_6�+m=|���)N���R����~��ԥ)�y���~Q�%(~�����)O�}����,�rIj�Ik*�U ���W��I��=����)C���~��)Jw:eg���P~��^	+��;�lM��)J{�{���)C��}��¡�R�~��)JR{��߸=JR�������n�.�U �@�}��b�JR����8�)I�����J�<s�g��9�q��UR��J�����pz��;�߸qJR��>��R����k�R�>w�pz��4uǰ�$�$!
&I`$'��`�����%�@�eM#��%怬3@Xj���ȲC�ucI�fa�e �(k@ja��H���"I
���($�@"�B�LаԆ-@���m��d����$��j�&�x�J�6ăA,�u�[H�N��w)�]�F���O(L�A�l	QѣF$�LДD[���JT�%4�TNc�4��@�RĐ�C��aq�� ��چ9���%!<��;-��W�]C��#)f�a%�$*�LZ�:ܔKBP�%1)���K���R&�Df�/�N�e�烩�! $$�*��n tR۳�h��:�g��d�le��q��0AS�x8���n�Y��|V):X1@A �Ē)T�od�	!$"C�*CP@A,�I,̄��3:2��zO@�� J�#3�`�G~(&�]�AA�ȕ�14K��
haBEf@fQ(^8	�ԩ�M����P����}�ծ�f��0�f������q�B5�J�F�����e����v����6dr���t��z���Нs�6a�7���巣������k	�t`W#�"cdu��vDg�S0ZŽ�Ԅ�m���U �lj����� _4�aysm���s��&K1�q�'x�q�\��ܻ����8vwM���s��۲�n1�"�T" �z+��f��l�\%��9A�|����I�3 �+�ۅW��\��;�eH�<�Pب�յZ���Hv����KQF�J��ji촵 lqEu�Wf�i�Q�Ok��ê�<�r���B>�2�Y#/�����&�1������ѷ��U-Jf�d�{�*����5�j3��R�l�J�MUhC$�� �jI]��Z�8(��U�6�"�S�
�L:���n܂��Y�^��=d�ɐWa[m5��&���q�rlWT��o��8��	7\�ò=^ݣb��ojL���.��L��;0i�ȝj�u����k��jU7!OQ(7�l/e�e���f=�3I���^݂�<��Q��v���8�4�HY��y�eX8�vѪ�t��kzs����'USU/AƈD�Pd9�ZGd�K�ڔ�W�B�gD5�3��ԒѠ��/ EVW���dv�Hpx�uerHh�Yїomz�A�X�\lu��i�q3a8z��^��kl�]��JGM5�Y�O��ٕ*����ƬI9�3m�X7;d���UR��^� ��in���k�ԝ��h�
��2���
��&�8B�*ѹN�P)��m�K.�n� blA�{�
��W�7`��%�a)ү0r\�lOo7�7K�&��E靯^�tݳ��qZ�d맭-��vqt�c+�����NmU'`�;1mR�Uc
���۷mUٖC`$p`-��#k���A��Lё�����)IeM�����eUꗘF:�z@B�xs�A�ȁP U,}�ϻ�?���� ���;���v�	І=<E��L��w��f���[�P��7\Ʈ=.�pnN�vtt^lE��K,0T�.���ٺ�ܝ���=j]�ob�h=1��&���uKp�*u�2��;ZR:N6�{J�bƛl���$[��'���W��Y&�V��v:q��;;9��^�8ל�l� NS7.�Aܯ&NKpc;�m�� �LeW6���x��v�
�-�N������[vkv1P��(�n��ޔ��J�]ۗ�v��odzv�lWn�2Ot��'m��-��I,���U �AK��pz��=�=�\R���}��ԥ-}:eg���P~��~JB�&�*v[o�ԥ){�o�!������߸=JR�~��)JRu�����R�������⑴]����U �@�{��*�)���ÊS�X������ԥ<����o9"�@G5��$SPRѾkZ�8=JR�~��)JRu�����R��<��qJR�����R���^�l��m\�;War�U �AK�{~�\��=�=�\R����=��ԥ)����*�U �������R\WcvB���܇k�AG�}�f��h̗&]<Jw�d���n6k�����r^*�T��k��2�R[�t���UӦV��7@�W8���Ֆ���`�ﾾD���I,Q&�#	D$�Һp=`g]^}�}��������s��BC���*��Jho^<z���V��M�9{����@�������V�v� �{����z/��Xo#�^׷}�ݔ�mRC����@�\}�=��+ �wM�6��v
�����,lD��n&7 �v;BJ7 v�������9ȇ����mQYv�ҡ�ջ�"����N�@��;�DG �����sP��PX��;�yw���L����7@�r��=�H�Ti
��Z���M�v�}�����z}��s��V,�]X<�Xޯ�$ݰEݻM[��R�^��zӦV�/�L�>��s�8�����`}��R�%��ŀozM�9{��\wT��E:I�ҥTv�ݝ�=J�v��ok&�nΎ�!����ٻl)�v���7i7�3��镀lr�K�9}��=A���ݖ�v� �N��r�K�<��@�t��z���BC��M���/ ���= �tx�t� ����v�Ң�!R�����7�`׵�/��o(�_�P!����Rm�1�-[�O@=�BF�A"��*{3]z�����/t��_�^�'Tn}���L��ku���n�n��mڹ�\.�p��v�㱺��k��^waa9U*��x��n���/ ���Z���	��H�ݶ�,wn����_E�}��K����7�t�Es�;��1�촛X޿t� ��<�n��_E�uOu"Qn�իwwm=y��wG�_���d�]>����	�
TO*���i)���cw`lDy��`{'몮�������+uZ3?���������Ǎ��]�+f'm�l��g�����I]hݗPWi�.�ӫc�F�Q�7CM�z�V���6޹�Z�8eK���Di19PU�=�=J8;�E5�6Rv�<PK�R�˨�9��AH��I��@��� +ά]��ז��6-:���9�v���<p�t��25R�R��6���nf��zV���m�7||�3���mD�r�m��!.��I%K)zs��\�bk�[�]�vq.��ݴ�÷o=K��e��F�D��N�7��
�PU!!T����l�]�8��َ�""���݀x֠�������#���@�N77�H3�@��۰>�����$EX��5x�^�{��6����������|�HM�3$ʙ������I�޹�
=� ����v;�t�{�}�`��K����>�&����j�(.(�i�Ǵ[��m�mעSp����v85�,�t=���7 �����:]�h�!Gͷ��zK�{��>�&�z�XT�R*U۹.�_/2p����ԄU���G&���������>����9	 'cT��*���iT�W@��v�z[]�޿t� ��xH~K���А�-UU�����q��y��j��߬�ٚ��J)R8�itd�s`� ����}�`��wJ�`;���ov'mݘ��7����{Q�ݹ����67e,��3-"��C�i�yz�����vz[]�8���)	�&d�S3J�����ۻ�G9�r!#�wW@�N^�{�<z��h,wn��@��E�{����~�����zI��⺜��1��-6�}~�����|�݆�!{i��7"6&�L��������G�}����,�_���%K��|ځ$G�2䰍�E��k�ܦ�jT���yv���a��:v���6�8{j�:����HSU`{�����]�O�� �tx�?%%��i$;����K�}~�������	.���T�E!�X��t� �tx�:n���� 7�	ZE����]���s���=���c۰>s�t>�v9�r�]/v�����w�_ ��l{��v��Ii��o �{��)��_wG�� �DFhl94��&��4��ET!����Qй;k�I��E��͍�{I���uڭ��acV�����?� ��tz�����n�}
+��Օi�7t[w�j��= �tx��7@'�<T�R*1���iպ��= ����t�?�����q-X�z�u�X�BNH
�*f�B���t�/t�T��Otx��䤱�m$�t+M��^��u`��f{�Ȉ��DFy��OSC�s�mN:4Vg:^M���:�9랃���n'\�5��fM�B.Q�F�"8 "?��v��[Bvz�ɢ��:�r�j��G���`xzӦ�hNL�����<�w4ms{E�n�7VӣmV�E6�'+t�U��{g����i�봣�"�)�	��=�1��p�*�N2�^�3uCV��f�h�ҶkI#mb5�f)�{��
7:��43�⳹Ѷ�Χ��{���n�V��n�q)���J;bC�7�jp^ǵ`��f{�{����H�i;*��y�@'�<����k��Zo_�6�n��U$ʛm4�o ����^�x�:= ��<�T���V��Xݻ��^�x��Հ}�롱��=���C�Ҕ�i�7e���	:L��#�$�7@=�u�7��P'ʂ%D��5%T���7��7nz^�au�n�v�8,���9��p�W�6���:��o3> �<N�t���N�4�FE�'t4�������B�O9Ȏ8��c�t�o���xӪ��c��$;�Zot���N�4��H�	:M�yH�E�NҦ�)�m��&hޑ��M�*�{��>_.BGKH���U��1�����OI3@�{��wH�m�}���|��q����[�f1��;N��c���Cv�*����l�������0k?,NR�U*J���nn��/c���cu������ �]D�v��v;n��@�{��wH��H�	�&��(����-1���n���z��xa�:c��c�~ȱi0*� �dP��Ԧ�MH���Jl$�M�K����N�
��Ȇ�LĜ�EQЎ*�X���;5)4�J*@�D�;a{c�� �0f���
C��t�����������g�n�]��JB��p �� J��� t*8(�L@�x"=� c��m;x(�#���ὢq�E�Wg`}ֽ��z�3߾�*��JEF6�]�:L���}�'I��}�=�A���Wt��4���$�n��_E�E$�@>� �UJ�/����uզ��wm]�S�)m�ǯ8	��:����\�v���8N9{����)!؋o�����H��H�	�M�yH�E�N�4��;k ���@>� �$�޾� �}š,Uc���1<ǠzG�N�n���.�z����`8�Hr�ԊT�TRUM�I7@����"�G�K�_zG�}��:2մ�,wn�v�@����"�����t�w`k�;1)O��������ɰm��.k�4��3n����Tہzڭ�B ����e*)ML��X���}�'I��z�,�ޔ���
�i;���}� ����_E�E:G�w�*S��"��&���	:M�>��XS�= ���6�	�]��@��}�@>�G�I�7@>������i��v��u`lr�ݮ����`{Ӎtr9�:$\V�e�-	�r1 �&2b"`%�N��BU!#P`�.�LD1\��1t��C�'���ӑ�{�Eq�@sV^;2z��-�ɝ]�C�ڽ�+���Ǯ[��Y��R�nk�zcB7Pm����!�R8�,�[���mJ[D+Dk:��@��=�BX�X��6"���wY76�#��ۣ��Y�r��cuÌpu��au�th�B�OB%��n
��]e�쮌��C*.g6ޟg�1-�`�1�����L�ӷ�ē�9�/S�����|����r�C�F�v{��eGq��whGk�.�{N.���P:ۘ�;��Y1��9ӭ�������k��ߛ�ޜk�4�h��%�wn˵i��m�OI�_��޾� �wG�{�Ƒ�-;U��UAUW`{'�y��~r9��v��ݻ�FEKDJJ�SRJM� �wL��#�;�t
����:���wN��v���x��H��w�&h��X�wG�}9)�o�:L��5њ�,`�.�a�ƃ��݃۵m��z�|�m�H�H۶X�,�KnK�{�}��_E�|�t���H�}TW-7m�#e��{�~x֤���K�T�$�v"<�[�`u�@ϱ����p�T��4��;k �N���tx}�n�����<���K�J�v0Uf,x�>�����I�޾U���uz�:�wm�j���6��t��{��`Ӻf�}�$��_��I��bwe����C����x8��iG��eı����۫��I�k�E��Acv��} };�h�������(�v���T�В����3@>�G�w�&�z�,�WӨ	L�V:�h{x�f�}��t���#�b1 ��+��*H@�a
�H�b�<��z��ʮ�w�#IJM"�ں�������޾� >��4�}�����5i��<����};�hޑ��I�߻��uRڻM��ҫۍY�c�^�º�u�j�(�l��+�.|��3����h��?;�x�zG�w�%�����^d�Ԕ�J��Ի]� ���t��|�����3@�֕
K�lV�[���;�t���(>��4�H�uur���m�qU5vȅ8�z�o{`y��dDB�D=�g8�B�>vԍ�n\ww�N�zG�w�&�^�x�ē%����5ػ1�͎����hN�K��IzY��-�-U)hD����S1��j��o&Mw������cw`y{�Z-oj�y&�`����14�UW@ϱ����tx�wG�{������+��l����� ����������� �����N�E4�L�o����@>�G�w�&�UG���/��T�����VbǏ@>�G�OO�������]�������&�@�%Uu�߯�߮/H��ky�ўS��:��!�m:�`�Z.1�nk��ufݮc-v���e㶑����[K�Ql�xwg�]Z�ٹ�������������K2.��ꌻlZ�N����ywԹ�:��⛘���Q; (0�W�[��ʊcQ�>�rv�8h8��t��2�)�/Z&�杩�3�+ъ�uv�N8S�<9Ua�%�ծ���~w�|�����:7>�|�L��;�jJF���s��oW�nf0���i�2�j�hB�m*�8�<�$�Ej��;o �����>^�x�wG�{��:��IBn��-��ƭ���K��p�s���[ڰc���7vr#���dMU�Ljݖ&� �N���tx}�n���K�:��@Je������o����Q��<��7@�{��G��/-oj�y&�a%BU*�i*������N���x��7�@�8�izq�q.�[{{kc��o���f�hۨ�r�/I\��gߎ���{�}H'[5���<�����3@>�G��UP�I��/�Wr���i��w�N雊?"1��^���ʺ�߾못�=�\�/��R�I[ui��ı�h�����5/,{=�[ڰd�nI�]�V�i�x���I���/ �N���_������t&��"�N黫�>^�=y���� �=���cw`y-ߔ��v숹q4�ڲ�m�n�ե�%ƴ��Μ����`���Wm���&5n�w�|�tz��<��7@�{��_N���[�:���������~�;�t��^�������Ap�1;m][I���t��^��RDL�+����{�= �H�}TQ66�J��-��"#��s�>Y���>�:�lDr"����7W��I)DR*"�jz��:�"�{��;�t��^=~����2�����`ήq��۱�k��ذA���퍷\tF�1%d�1\�ܻ��Eyy| ���t��|�����@�֕
K.�v��M'm��I��UT��#˞�@�����c�����:�UML"�������K�>S�=?U��<��7@��L�ƛ�bn�?)������~�*��~����N#@�(� ����}/5�5ʽ;�A)ڷLln�7Ǡ{��?�~UP��{�X�z��:�>MA�DȢY[gbᗛ�㣊G�ې��v{@r���~V��[�N�WV�m���n���K�<�t���tx����M��䨺�V��/t��_�)��}^6��"9	��:�%(�T��������`{t#���v���|����1+m��uf,�z�UT��<�n��{�#��{X%(N.�v��������t��^��龪��߷ʾ^����I��v}��`����<��

@��LJ���^y] ����(�S�ϙ�v�¹ћ�߆�7��f �5�����{��E 8�4	BEH1��q�I�:�c��F6��4���|N��_0�'N�M���	�AIC0C��GZ#�xse�Ý�Y�v7�h�r�P�� oH��XY�6J6LH�X�H�;1lA�S�^$)�IT湬Sc&�Ҟ	!*���y�� ����I�rB��)��F���(h�Ԡ�� hĪI<�ӷF�2\��^�t?#��C[E�@�tS^���l-nY>-��9�&��㦠���ذ�h��'Mj��W��c]pnl4��7;���3�A��
��
��"�ҡ[kH�nn��[*���ɶg<��w���ӯu��RGI۶�d����u�kű��؈�.��V$B�ˬuu�'��/3����l�{C5��6UK�gm��5��]��h]l���K<�UU��F�m�(mW,=]a�vd ۪��Qv�vۅ2QӨ��q�55mT��k\��f��Z� ����rҮ��s���<��^R�B���)ۻҭ�-�8�c�0n�r���&�"i�6y[�ɉ�P4�,��ԸҀ8�����c%W���j��*�9�/T�U�[d�̪���+U��v�� �Ip� �K]+�˴��EP�92d�TO�|�Avl����t���e2�vqGR5�<�ON�)3P�<�ZnJ�۞N��Ԧ�8q.�Ǯl�v���ͫ��6:^�1q+B��kK���gcm����J��B)n'=V�l�v-�)�mnwc�="#�]���=Xp�f��Yٖ��[r´��,�ݧ�����ud��۠\x��M*�UI�XX%���ń��x�ډI�[c��m�8'E�\ԘjW�yJM�02�fF9�6A��u7��7�`���r�ڎ��h�f��P�m�zӵk;��Rg6]��`WC��Tpe��A4�j�����Y��	`�$�i��*ۮI��abŜ��δ6���d �bK�UR�e�Gli��$�@3���X�h�G�TRƷ�����k���ZlѶ�&�n㹕jb�TɹM��-��!�Y�'���� �.��^���rr��.\n��a��%�9]�L���t���\��8���;8ps�B *�UX²!mU,�bv��[Dhep ���vWf�6�*�5� 誣,����[<��#����� J��Q��w{����ww���wA笄>�Рp^��@lS�N!��'����b�;5ѭ̳�x�qT��0����r���Zn��],E���6���؞�	F������9�m�x�u���W���Nۈ[J;m�����7�F��;\<�&��9�sm�n��iY�ۜs@>�ۉ6�n�[��L6�1�q�nZ1���z7mնV�r`n�v��t���5�Rvah.WfPl�9AXA\YEy'dUY&ݖV��:y�K?Y��N��pa��i ���|f�W�6.3�wD�;��E�`B,,-+t[v�����t��yw�= ���N��{�2��ZCnՉ��<��= ���N��|����IA)�n�ll��ǠzG�wӦ���X��G�w�. �XҲ�մ�o �M�>��X��G�zG�zyU.�؛�*.�-��=�ƺ��u`y���n���8���]y�.�I�p�;�jN4�,�%U���t��^P��7e{N%p��nX�Mbw��V-oj�>�u�3���#� ̗��yz��)�
�iЮ�f= ��<����r��Es��Ig]w�=�ƺ��u{H�J�F�J�eMQJ����=ݻޜk�yfc� ���@op�T�ݵv�C�w9��RO�{��7���}���ZC�e���<��=�UP��G�}�M�>��X���$hQ��K����l�,1'��=`����r��=ͳ��NZi��ΐ�g!R�Uڰ����n��8��9p�oj�y�[RU(��J���^6�����`]��}�(O*�қt2'�|��ߞ绿_RQR),��D/�.�c�������B����QS*M.��8,M�� �=��x���_E�}K�
J�7I],�z��<zI�޾� �����t͹����Y�u�D���X��&v�^�]�{u<M�Ʒ6?���۱�{69�,��T�X=ݻ�N5�<�1Հ}�u���&�T�ݵv�@���`]���>�:������G� qS�T!QJjIJ�tM�� ����B_=ݻ�s�`���2�t�V�Mn7�@>�:���zq��1�"5r�^������߿o��xW�$��Ɠ.�[I����t�}���V���@؎r=ښ�
��2��tY���:�r�t;mⲚўœ���ѻ�d�C=�%�I嫱����/:�}��{�@>�G�oN��.)Uܦ��LrH�it,�:���r"!s������g��z�,i}B��m�Į�fU�}�u�/;���}�ƺ�{X�T��jح+t��zt��_E�yw�=����'%)]�T�ݵm�����<���}� ޛ�8�y%J�E*��s�e�܃���Ise��۪�N:^��J��lF$i̼rU��'^��m��Z�G9cO;q�lL.��;��\�#OOX�d.���� �h&�9��c��ưl�Z��9�o8���:���u�J�u�rpr&G��*j�Q��5�����x��-s.�٭�s��� HF5��=D�%�=����Y8#F���Y�2\"��t�.�J�/�d�E8�oGe�hݗf���p���0Gasom�h4ی�j�S`��)jv[��7v���~� }�u�/;ӑ�s�=��t���I���f�W=��l�c��#�	={v�^��{=��r#���@:�'$RTL:��m�Ӧ�/t�=��G{����^��Kb�r�m�3 J�%��l���ݏ�ǵ�>z����(�qI��H\�0=��|RUG}�^͝7@���`�T��Ge]��U���۳���ζ���W�[�V�.:�ݪ�^u�0/;����<�[�i'A�= ���N��}�ƶ"9��DB[�j��JKv���R��r۹w�s~߹�*I|�T�%*�=��.�i�u`{wNG"n�il%T�ݎ��˧��S�����<��~� ��O� �n�%���K��=�������t��^+�P}b�ՒGr�%���}�^���RK�/{`yc�����`|�'ٚ�T*9C��x�=�Ë��-F������v�o[��䍰������V4��um&��7���|�����3�� ��<�:�t؛�j0���d�]�r"8�f����$y�������Q�uij���JQ*�[��^��߹�W~���v�����������n��_E�}K�JJJ�ILK���>��^6���N5���qd����R[�5UIRSQSIUUt����d�]�3X��t������^�K��zm�d�Ո�A�hmn4c���\M��=gF��+cd.
۶�K}}`�_E�ywtz�ty@oI7@��ED�L�E*T��h�Y���9�$ok�|�v��)��s�������S6�{�1���x��t��0.�@��%L�jƕ�N���x��v���\���}��W��D�P�w�vG�}=�T�cI��XYv��w8`=����c��xۻȌ�!�0+GHp�y�#������iNkc6q�݂�KZ��w��I,��v�~m����~��@>� ޒmV��}��tIB�햮�K33@>� ޒn����<�1��s����B7IKv���EB���J���|�v��c���&�Հ{���$��$����ڻ{�~��/c��噎��c���9绿Xp���L�E"��j��yfc�y#������wn��f9�7��q3~~|�5-�<R��\\����F��WL^5n�ۥ��g��S���S��o��c��牃��.��gm����$2I�CA���T9�{-�pv�qv�Y��1�j�d����y�1s2Gd�vy��6Z!�v��d^b��Mu3탬�e�\3��ݳ���nas�b�v@.���.k[&�Bʘ�$T�%����7�;��`:tR��ћ5-�u��zݛߝ���G�;�}\���ᮅg�-��KWe;j�1�ڸ�3��Ya�nݛۅ6^ڶsucM�fc�z<zI�˺^~��˻��;��~�cJ˧VҶ��$� ��<˻��������t�Q���♂I����t,�u`ls���X=ݻ ��UR�f�fb��S5]˻�����7���W��}��/�E�*R�v�WA�3�}��$� ��<˻��:u:WT�En�&Y���qz.eu�6wn�n�uX2!�v�:1�]�ݛW���e��wm&�m$��7���f:�Y��y <��@�`����]�r[�����y䫂JĄ�P 
z��`�~�t����u`cu�/wz�� 8���Ți���r�= ��<�oN��wG�}�A Uۧh�nխǘ���]�� �1�Cc�'�j�y�����J*&�������^o^��t�z�tx��G㕖��R��Ӏ��c���n�v�=��]nѵ�d��Kv[�����ȑ�e�wRD�$��w~��}�= ��<zt� �r�M���]ӻM]��yw�=?�tx���tx��t\D�nհn��3�}�׿{�]^������&B�a�X&���"�)���xt�0���gION�(ON�ԛz&H>�6��.��o�ӝm�'QsC�2�Ã��4�b���=f�@���&&��;����`)�t珊l��2M�t�S��*- X�m5� �F��@�5�E$0b�Z	���׼0��l��i����ߚ6��B��D.V��=H����R��a#�G�5�7�ܝ�� ⇚1xH�VH����}P��{Pޱ@� v	��_UE E�l<Q<��j0�{S�}��]�@�Z���ݴ���Ut7����׷`y7��<����>� � D����Ccv�ot�t����B���ok�^<w`dFc�{�m�Ũz��E���m�eB���Ou<[��{u���H���g�o.""��.�G�wG�oN�����}�A Uۧh�i��ǘ������t�t� �{�i���A)�-XһC�i[o ޝ7@>� =���tx��.���&�Z�v�@�>� <��~�U]����a�H�*����?W���@>�)�4���5i����wG�oN��|���߫��{���}�{񐭑d(����0X��C]����X�G62�4�E�n�1GbWc�������4�ĳ3> ��� ޝ7@�wK�w�f�8����[c��m�Ӧ�_�>]���wG�N�"WI�e!��ҷ��}˽����PwG�l�7@���W?]���j�U.����{V�������#�u�X��(��N�v�V�c���t�s�Ϸ^��r�tY�u`o9��_���-�q�q�����T綅sMϷY�!"�W�鹬�&(gr���-r-����҆3�p�Wl�6�onz��jx�*z泳�+n®@]���<p��&̎�w��rSr���5��=���FwSWg��yq�.�&�R���u��gl�wa�b�QF�b˝�N��%m!Hձ:�*��:|��5�>�R`4�f�f�_n)�y
^B]*�On�n��{ߞ���>{׻���I��?Z4�s�u�]u;�����xe�m`�!��Wm��wrBȮ�b��J����U�U�'V�m�{������]�@>��^�TFƓ�P��{�r�9����b9 =�k�}���b"#�9ȈA�2������U!T�O@i�ڰ�:�}������5}�d�:��5*h*�GW{ڰ9�������^�x.�G�w��6��blv�V��t�����wK�9w�= �H�	���P�t��XնRmU�EF����mWqs�ۏ�%.��v웣��v�v6B��m4�ƛ��t�.�G�N� �N��}�S�ʻM��� ������d|��b�@�Iҋ�����������PJ�cch�nսo1�ӣ�'Ӧ����9{��w�=z�S��[]�um&���_�׿Xc��g�Ձ�r�:�q�1Dli7��
�����^{���G�O�M������Wc�]�j���
V��sv�v؈q�۶��t�v�ہy�O90 �7M�b-�Iݻ�"�tz�����|�"���s�/	��-IMt�f= �tx��t^�x.�G����Z!q�v���v�V��t���^~��Y˳���G�t��U��M4��M���{�����}:<d�x�Ԧ]����[w�r�tz���	��/t���%T��7�I�Q~�.X��,�Eᓱ����&0�]�"m�۶�چ����'��>�_t�������v��c�������t^�x]�@���)K��*[I��	��vG8��zY�u`<uݎDq#65�Bڢ���JI���{=��:��~�>�>�7@'.(��6ݕwM	ݻ��~�������t;�������~�(�j>Z��5ʾ���P"-��4�Y������߿T�t���^{��>�r��Ue�s���G�Ǉ����n�x����Gi���s��|�=�E.��MQIM%T�Jj������@k=��"9G#� {^�@z����V�LLi��9{��w�= �o׀}߷�sR_��UCk�/�Jd�NI@jx���ɠ2��v��=�Ӧӫm�����}$x�t� ���*�w�=z����N�N���}:n�wtx]�@>�<D��[���\Q�Ev�����Zn�ĺR�ʔ��t^�A[����:)��'I�1g:tLƺ��zq��9p��e6퇞�m���n8�M��U��y���Yj�[h���up+�+�e���Б�ٶGn�e�b���^��%��3���ڻ�U� �]��J9G���Icd�����ٝۂ`%YA;d��Ӣ����/q��m�&�sW(�mB�����{��~��Sx�뎔ꥃy�[gv����{v�q.�g�d�{g�4���&��{�G��,lm�j�e�� �tx]�@>�>�7@'.(��[mv�C�w�E��������t����T��Y�I�&6�Eb�Ǡ��� �Lwf�<{]Sǵ`f�8tRSEM*�IUWCb9#�}�n�k�@k=��ӣ�:prW(�ʶ�bcM���/ ����ӣ�'Ӧ�,Y�P�枞ʛF�L�[o8tq�v68�u���lsb�5b��XSyJ�e�V;�K.�[w�E��������t���N���'L��mݽ����#�����]_��U�	�&��<.�G�OP\)(QN�T��M��O�M��G���Ж��j�=�k�{��1����(J(���؎DG9Ȅ��tOՀ|��@�N���qr�miݡݻ�"�c�c���9��{]}�n�3��yyoɧ>��L�L�`�v�(�]����0�N�q�z\]���\|�N��X����G�O�M�9{��w�=��KJ1����v�M�}:n�U����tx]�@>�Ӓ\��.��Z�1��@;�{�����҆ 2.��d^��t*�̀lIP1%@�B10�P�4~$�t�HJ���DO�|���n�_�x�M�;�:���"�MR���D-��j�=�k�?�;�1{��@ t�m�m��y�@>��U��~��׽���������>�Nn�bގK@��6�;��tuq���#�����7g6���H�e�p[�\�`�����w`b�9�g��DG9Ȱ�:��R"�F���J�v�@�H����玺���G"j;ASH��Hwn��:= �H�+�UUQ>�7@��/ �G�Iq��n�tV,x��#�'Ӧ����{�R���~�$�U�%T|������7>V���m%m���t]�����}$xI\��¤�.մ�wVS)�i��gt��mU���=\�M�uۭ��p��7+z�bcM�˺^{����?~��}:n��8u��-��-��"�tz�����t]������@;M����y�@>�<}:n�˺^{��'�.�(ab�V�sU��-����i����{Xo#�����3��j�3<�	r���c���{X��t��v�v#��r9��C���a�p��ࡣ`izC��C�^.��!����6]���D�w�z2cJ��:�	��ք1�өp(ChO���L&�b�X���p"X	ġ����V��`V�-Y����Ť��c�J���M�Y�:�22L{�M�1b�@P�%	D8L�MED���*�A�������(A�֞�ڹ�!M^% �	u�|3 ��+%�3�GA�� تR�	(��N���U1�!q�۸�n�۲YAm'@�aol:�������n�[�+ٹD�0�@���&�m�n6�o+��$�f�X:#%mk�5�^s��YB-X�8�6հ�9�s�m���@�ewX�sN��e�x݊��9�P#;�R��Z�Ê�/�v�9zᖺ��wB)q�L��<�۫n��waMg`�ܣYa�m�2�'k�Y�h-Xp��m�㞽N�8�6�y�UK� ]��û��ɸ Cs���V�2�����k�4�E\.�3��#�X��dJJ�Ζ��v����6�*fy��uҨ���<f���x��n�0�ݶv�;'��r*��8��Y�&��-@����Q�c��a��(ch��*6�B������U��HâU���J d�*��"pClڱBH�uʣz��Ǌ"y1�ͩ ƻ/;�/GM�ת̸�v5��ɠ��.�2�/&񢳲vD��U��3��^YNM�\ݢ�m�\�z�����c)�m��Y��	��k���Z�&�Rv��Ӎ�>���Y��q���G���(ݵ��f{+�#l�7���g,�4�ЅX�\�l�B�� Uc/g`�P���M���A���uUI���e$�+��X�6�����e)V�6.H����dv�Hm6�:j�.n���ے��V��.{d�=��d����s)��܎�l]%�]�uc��ѓe8����d�k�;���Mn�[Sz��hs��O(R��Wj��ƴɸ�ծ�eV�;���6ض�,	 ��j⵨�nHMku��SI[ �I ݲn���5���4�Ht�J��)-��[B�6ؐ�%:m��{ojt�+B̩�5Ol��9�9"�]�Ge� +����5[Tq��gW\�l��&`ey=*���qZ��q,�@q�1��s�J���UT P�P-�����]5�d`)��15��)Vٷa��m�Wj����^��YV96���{t<�����@��Y��*ՌQW_ǽ�h:Px�
�B�=�qP��hu�1}D<Q�O4�	����*U[W�T��WWm��7.]�;N;�r݇Ke��u�vN��l�����:r�.�L���ǥ.'�n�nƩl�3YM	sF^�,�u��b���e�&n�mp=��Z��t�k{X,�6�.�XaM��{ٱ��Q���ś��v4��1e��ayo`z@pGj]�b�	���������;7v�h)�=Ol�������8η���y�M�M��㡈�>^���������Czt#G���W��ʇ'9Ì2 ĉ�k��IkVyü��M��챺��۸��G�t����9�����/'a��an��V,x�����t.�x]�O�rIKJ�5v�lvһo �N��ywK�"�tz�H��ؔ:%TQE)���c������@���X��t"��vd(�RT�cb-��"�tz�H�	���t��Ē�3�N���Qm�
�J�m�q��E�ţn6�v5��>����m���m���m7n޷������t���Dr�jx���	��
%B����U`w����IqUR�U�X������| ��y@{�H��.��5I~t]��wG�E�������tyT%6ƛ���ӻ�����}�<}:n�G���5|���)&�N��]bǎ�>��lr#��׿|��t���Ϳ;�ߟ��>6G�;%�*�E��.�=v;o=�m�άJ<Ҧ�؛]�ۜ]v�v�\ u$�J��i*��}�n�=��5��V�H��ܕFZt�Ҳ��{�� �����#�'�M�;�9S�I��M�T���E����#¿W��Q@ I(P�d(��2��h �]�8�gbϽ��=#�6u���nݽo1�G"�n���v��]���Ձ�:BZAD�QQ4�����m݀{�<.�@>��#�%bJ˨�:p�ɏ]cr`�g�s��F��CoI�/�3�����L�E�%[Mբ]������:����Dr�o�v�qF�TR����ӻ����= ��x�I�����˨\���ث<z�7]�ۻ7���@��ڰ3%$��S������}$� �tx]������^���WLS#�6p�IӦ��ƭ�{�<.�@>�>�n����wYE�1�tյK�l}�gv��.��p�֔�n"7=�24g��`D��4P[)[o �����G�O��Z����@t��X�m�w��= ���!#}��`��@k3^�DB�n@N���T���i%U]}��`�:��9�%���`�����iq9��R��PMU�o#�K1�tM�� ���Cb#�-��� �q3�*��J�*�MW@k=�����D/f�X�ݻ���~�*�'b��1����}��z��e�R��\�"U��X��O"smY�8H�ɪjy�֊��ȫ���G���:�[�O[�G�tpɳ>��ӱ�ct�����V'D�j��;�[�٣jݞ�4������⣪v�eH���G�;�5�n��9��t�hݞ�����i-V����l�6����W��Ʊ�.״�&6���
� y�^�]���}���wowv���%�m���:��v6��
��=���;pt����m���rr�ĸ#|0�*�]�� ��ͮ��x��=��Y�@�m�i6;i]��O�M�wG�E�������(t��e�nӷ����^�O��#�>��tp)��Am��[o ��7W��y��@������u��@cV�nݷz�c��G�}=&��t^�u`lzH��0�t�T�W F ��7Oi�ζ�I�F!;A��K�68K�/\lnp�M �B��QQ4���ۛ�`yf9�9{�?�U�t� �ҔK�j�j��c����ϗ�V�T��f;��| ����:n�T򮻖��V���'v� ���z�H�+�~>���t��]K�(�lun�
���}�<�N��ywK�<����i$��&�N����N��U~����/ ���z�H�	_zU��E����jƭ��9�W�����B���7;��:���ng�:@����趙v[�V�@�|��= ��x��7@� q2��Qi�iU=��n�c��DB��r9<�k�{��<����:�)�i�n۽o1�W~���W~}��ul��N~�G�(�����ʺ�������
����\V������U*;�߹�n��^��}�<�JQ/�]�)�]�� �tx�t�@>�����o����μ�]��釹rV�sԈt�:ΝU�^����Nܡ.6r�*U^vq�����s�wϔf�J�V�ݷ�j�H���{�n�{�<�]JZ��m:t�.�<Ǡt�%�UW����&`��������#��H���I�cv�v���t�����= ��xT�)J�bmP���UWa�Q��B�����X��tD#܃��_n�� aL�&�V��5w�z�H���.�=��lDDDG7[$���cd&��X�k��{�;v8��vC��9
�+0�}wRv�R��D)�n[��r�e�e��n�@�=��َ���u`?@:�sh���ěx}�n�{�<�;���G����U�(��.Ք�$���������@>��t���R6��T��ݷ�|�tz�H�����~��ǻ��<�]JZ���:t���'�����I��t���߯�z�*�"5��⍎���A����� /F�9x�J[���sI�����t�4������2���݀��ѣh�v�s��(
���"y�MN�')�*�ԇ#��O5n�5ۇ��q�"��˫�;#(/i��/b��Y=�o�vCv6����n�}y�[J����[O:8A.�j�`�\�.9[���q=#��W@|3�;9s�*��۲��{9�;��������j��9�f:��]�V���v�&�k�;vZ��~n}�Q��۳�wa �J�LL_�����������Wt��;��߿W� ��x@�)Kj�n�v[�v�@�|�tz�H���n��_�W䎀�T�(I�i�����`cu�b9������݁�O��>�P�~j�m۶�[�z�H�}�����s�-<�V��3!RB������gَ���d���>_�= ��x�H��MP�*m�m7;�plӍ��ݷ�,�tv�9&��9.���]����U�;�@;{�� �;���G�w��t*Jn�mZV�f��o|����~�]:⣘G�0hP��J���	��	�f��|��� �c��r#�H=��fvf�TʩQ�5ڰ=���c�7�Čok�|���zu��Dm+M;i�J�����t� �tx���}�<�w%R��V+-Ӷ�@=��wG�t� ﻦ��\��´Jm�7Eݮ�yg!o+�u.�q�����dm�y�n#�ŭ�=����?�M6R���wG�t� ﻦ����>�P�0v�ݻ�o1��#�;�M�wG�|�������=A!��Uӫ;�o ��7J��߷�f�허`� �ؑ�6h�٧B���v��*������qB8`�mX�Sk�>��*Y"�Iu����uw�|ƑH�RJ���0��N��C����14�ㅋ�6+�E
mS�M�b�? {���Ǡبj�o���Q�UЋ�?g��<�z'G�N�����&Sv�;ot���)$z�H�?~�GwI�#7mZV�c�����= ��xf7v��]b6c�
x�٤��U�km�f�� ����\�\/gZ�6��s����qZ�2D�-ڹ"�w��}�������lD_#���wv��$�T��UT�RS5]3�ԃ��[���t� ��Tt�j��e�Wot���)$z~���#�;���{�0}��\��P����,��ڰ=������|�93�����C�EMMUMMT�W{V�7]W#���~ ���)$z��L��tBg��BOX6�����nڮ9�����݆_Y���ld�mU���5i�[xt�t���RH����.�)v	��EҦ�� �c��8Drb�ݫ �ݮ��ۻ ����7mZ�Ӥ��x��= ��xt�t.�x�W�]˺Wo��N��x�
�_�t� �n���/ �G�wZIDF�nƚvһo �m݁��r9��f�Ż�V��������)Q�!͸�����`jl��iE1�*�$T��s��rA�q���ڲ�;uţS�3�y)n�����@�C�\��m�z�j�����IzN��N˙�&q�p�n�����w.s�s6�#���^�e����6�r����� \�+d�N��nWq�-g����K9z�|��8�!��uvH�Η�l�rXu�@ ��y9��nV�s��v7=ew0��g ��l�lz�k��@튭�9Yvݝ��rҲ&�o{�Wh�����֣M�g[�"	w���n���f�۷��Y��^^���h�<n�z�ޒX!�Ի-�p��������`M�V����1�v�)5�&�6� ��$� ��<ޝ7@��K�>��:��M�m[�vkyz�����<wg9�/c��亮6�3�"���E)T%5]ȅ�׿X�^ﯤ� ��<{���`��
UU]���s��9�G,m����t�߹�<����G_2�r�i�AOmm��ӥnp9�NRgd�,��bN�+<���j3vի��Zwn�RH��H����Ժ�^��`�Z�I�D亻��/$��U]����l�ī@A0R,(b��=a ��{��u���S�z��J"6��M4�3U�>��v���M�"9ľM�Հ{7k�fy��R�RM!M]��r#���g�|�ݫ ���@�3��h���I�i��5wH��H��t���/ ��$��S�S����mԃ�nZw��q�.��s�k����w���]������n���`۶ջwYm���#�3َ�/c��r9h>Z�j�܀zvHQ1T(�*����g���"1c��-{�`y��#���c\N�
�
"W.��<�~����g��JRJ�J�VUtx��}�U��}�]U}�>��cv��էI5n�I�4��N��N� }��RԴ����4i�f�N��~��ӧL�'\� 'N��o�}�[~>A�X����Z���g�׻<nִ۪Oe�;b�S{ks���㲏1��ťJ�����5�۰Kk�>��!G�*Q�ݫ��+{�N�DG9 >���<x��� e&�'�Zn���t�:G�N�7@�r,�J�~t۶ջw�����G""#�^�t�{v�mt3��"�:IL��@��S"@��v���:�k��U}�	�i�]�e�$��='M�?���]n� o^��7]��G1)RO}�N�c�؜��6ݹ�M�s�곆��z}��mN|�t��J����H����}�"���4t� ��7@'��ն�����]�k ;�L�	�<�t�uȰ�^�w���� �O34�u�<�;�b9Ȉ9��5���z��@��B�F4�i�J�t��mt���K^�t�5=JTTԩ&f�)��Kk�j�Dk׽�^��*�߽������C%�0�X E�E��"�s�������������e�1Y:��ɓ��Z.�rmiv�b��e�z��v���]���iɧm����'g��G���:�]�R�5�Wn�[�E�=�ej��Gf�X�l皛�����ZG -�������q�6{g�����-��m�)��sd�&D��BWpn^z^6�0Nj-r6k��N͸lr5��n9{�s//M���;ɗv�\�Vr�-RU�򪤉��k�~�w�n�qj�Gvl�v�g���%8N��J[��Bv֮/n \3�d����*�i	M.�f�}���@y���}r,�@wT��m[�{m�� �w��盻䶺 ����� �Wm��1]�+o ��7@�^ ON���<ӥ��v��WE;ot&�����f7]�py�����ն�v�wi6�����#�'zM�<���},�?�݉����:ή����ӷl���pt��#�ۭ��F�[')�:t�̰����e����#�'zM�<����� ON��{šJQ�[cM;i]��zzMޥ�_�����x��3@;�x��\iRn�N˻h�{�y6�珶r" ��y���=�b�UrR��HSS���D$�^��$��x���]q��>��� m�jݻ�m�ht� ����yI/ ;�l�C��qL(�ځR���*%��&��� �k�ɹ$
Q� ��v�H�0L�)%R�f䚤T��)����v�nz�x�����jFk��������Uv&� {��v�=��@y���s��<��hwh-�w�ӦhzM��Dde ��P� E� 	�x�h��|��}�Ty�~��^_H|��C��Gy���u�-�w`nN�����r#����la(��Jj��)Q*h��<�K��t��0�zU��V�+�:N��C��}v�8�'#�Wk\n�F�Լ�onۉ莓;�&���*)������>�_o��t��0�&��Q�e �6��;���߳����H7�_���n��:^�QDꔋM�ջw����;�� ��n��:^ w��hPMGĖZ���If��J�}�}��}���W�{���i('���<�G;
v����x��QP�EU]����@3ُ�y�:-�w`{%��v�\��n����kl��g�a񱝺q��h&��snz�q\J/��f��)��jz��}�3Ι�-�wȈ�#����uz��*����,��3@�Γt)%�wt��-�cccm݌Jـl�n��$�
����PwwL�;��;��Ҧ�v�nݗn�&��31���t΁m�vd�L�-�I7m![� �wG+������ʾ=�!� %1��X �0���wRR#���\%� ��\C���s�n�2 N��VP��� �d�:�q��6�d��P�-�)���=r���`�y����C�!�P:X �������� c��U{����HH�0����L�ih
֡�Gӂ�h�B�H�I��.��z��f��7����^ �0-��.J�ȵu���[NK�pA�J��M<��)3�."������ZL��iTI�Hj��v�.�m��]m����Y�U8T�w ]�b�3��#s�1s�<�d#������65S`��3U��X+tU{�]�_4��:�M;\�t��sE���of�^�-m�&�q��tڥDΫ+%m� �m�Zv-����e*�C�ñ�ei�#�n�Ȩ�d��n��>A�w���.(�6-�<�J^�[�� @j��ɭv�Z�/J`2n6jU{G���`K:��g������q�tetN�Ι�N�����v�6��غݵ���g.*��+�rygAl�9��W:��%�����Da`�/9ZtmUR\��0�g�NjN�P�N�[`A@:�N�;�3V崓hG66б�RhvY����9�]90�sl�'2�R�U=]-]m�@��S=��Ý�jB*7kK2=���6��Ԫzl�8�CxKh+j�C:��9W�u�Z���FX3p�nN�� ��u�����e$1���1v��:�N�r-Vn�Z^zIk���,[Qr�Q{[�%��=��n�`M&�M �v��A�� uUj2N��b`�RꚩV���"�!�:E勢-��W7J,l�-�2!B�A����0���43�]Ȁ��3�;�O4�8S�)���+�g���Z0ۍջ8��s���֍t�X�Ol*f�ۆ��(������V������m��m pH4P,��zs�{� -�F���ք��J���� �Ik����YZ�<�M)-UUU@�=����u�f���.�N4�U�:U��h1�]
�E��Q����]�f�"w��v���M��y���q�m#�]�OM�.p8�;lL\q/' WK����@�ay8��{EZ�j�r�� �rY� Xe�@PY:����`*��U� Y��"��аs)��n�ۜ��cv�S�.� �U����@<N� ~D�A��	�� @~�/���`��ںD_D���ٛ2�kY���դ�<��a�����:�ut#�n���G���<t��*c98p��Wm-��@��e|�*����i肹�s'\mɦ���R�$���c��X�#��.��ά�[ne�O)ñ@��'g������2_����~C��6�!�s�rq5lN��e3J��
�]>%wVMs�ͻa8;���.G= H�j�"{tS_����s�G}r'���ٞ�k8��8���b<p7\�>�p���ܥ��wIĕRM�k�ݹn\��]�|߶���w`y6����pĜ�&*U
f�3G@�ۻ��#��vz �큘�؈��G!�V�J��E$PL���1n��31���9ȈI��:ۻ�`ˆ:��EI!1P�������1�:�n�s��&��O���*���в����8`�_����|-ݝ�E�7��{�QT�I5�-���x.���;p[���4��o����J�۴n�c&]:�j���[o����n��m�@3ُ�c�t�9t�Mw%ۻ�	/��ﾙ�.$�$��U*�"";`)o{`}�����""9	�_�An�n�B�x:O��;������Ix�E�R��V�v��o3@�߫�8`:M�<�������uj]�cI�v��Γt)%�{�f��0w������C�&ϝո�kormn�{$�,�tvǆJ��qѮw"�O�X�g`���m����=��`f:d�"!�n����9���IT�35 �f>��!��:��n��o��-<�s#��DL�*eW{�1�:�n�q�s�9�AÑCLSZ,#u���Ϲ��r�t�4x�)(�˱���%l���ߢ" ����۰3v�鰐���֝�!q�M����v�{�zG����x����Ӡ[���y!��%!��=]�S���5ۍ�<�1�5W>��ӳH��8XSyHM[y�]���ܶܖ`��f��0�&��� ���uJR�R�USJ檻�1�;�H�^����� �wL�=%:��&5N��C�`:M�=#�~�t��8`z'1)�"�R P���6"9Y�� �߾�Ϊ�߷���碸�a($����H �@ȇ����ު���V�;��T��X�UwJg@��݁�-�����
�8�J�խ��h87�t\\!��5=V��u�<^��V��z�m���4U�[�,I�f��0�&��"��t�޴����v6�d�)��[���9H͝����l�៨�ƕ66��M۲���-��g�l؎BM�i�>׻v�#�����v�������3@�ΓtK�`uz�j�n��m�ht� *�t��z\� ;��4������k��\�\Q�E,j�8��:u�:�+�6�뮑��qn�:Jlμ�N�3۴�����n�v�p���cnʸ���1p���Լ!�[@�ɺka7b�rC�l���]�m`����
���	�����Pmۓ����8�ut�߶������l7c���k0li�W%i�/O �Km*����.n��u�� #9Ϭ��tkm[�&7'vș.K�^�I&�k��W �v�vb'�� �v���:���k� 3[w<�m��{g�^��-�
�m�_���ϯ�<���c�c��cu���D,x�bvg�*yH�B�����]��c�gH��&�����m$��*t�����f�wH��I��ȰS���Z뺷bX�y��#�>�&�r��lD�Cǻ�2RI��J��wc�v���7@�� w�L��!+���*J1$Ɠ�?2���5��r���v��t�nnCts�������Ӷ�I�y���v�{�z\� ;�&ht� �t��z��)��ҡݧm$�� �t��B~U?*�l�����U��~�<���}�Q:�+I�m7mm��4�G�l�7@�^ w��h��آ�wM!��I��_��&�RK��t� ��W��W�"���*M��<���{1��=��@��݁�G=�r�w��qq�<=��x�!�A�n�1gVu-�<Eǲ�Zs�9�	�z`	����{1��=��@���9����Œ�$?�unı'���#�6t��z\� ;��4z�K���6�tҙ���<��yÜ����Ča�d\��M@!�"���)s0�|ET6��[�߿s�>���`��*t�m[M۲��U��� �f>��3�_�w`df%)��C�N�J��wL�:G}$����~���j�:Ln�n���=uیm��tu���x�G�)һ���۰!��n�VR��V�v�[o3@���v�nv-����װ��j�TCT�ـo���yt���t��0�U�e�T�N���<�I����ds�c�t�n��s&\�v;�M:I�w��t��0��u�`x�o���G ����U]UT�Y3~�`}����7t�.�w���8`�M�<�K�wt����w�ݿ��7㤳��z�Լu��۶�o2��fM��GY뭮;�w{��/�i��t�2ճ �n���^ {��h��{�T��m6��e�����ff>��L��wz���U����T;��]��:I�Ɓ��~�ToI7@�\� ����%�j�n�
f�X�L����=��t5c{�E���"�0��*�T4t��v�q�������:�Ts��&5o��T�u�H
ݿy���;q�viz:�%�F۹n{sj�W�����^-����)�h�ۈ������G.���uZ���K+l�2�S�`�vA/n���p;0m4bӀ7�s�B����&�'N���W�pdx6���=���n�s��铭;�ධ����+�����+��(��nt�)/V�\$Xva��xڞ�4ZN��e�vrt�����www^���U�;]n�nd.5pcV��N)|&��W�s�J�^��;oOb��K�\���x��=��nU
j��}�?�tf>�@�ea�/َ��:�>��.F��7r��߱g�I&���:��݁�k��"" O	s3r��VZiX�+@����wM�=��`�L�޴�K��e�n�+f�#�_y���n^���e3�^ea�<�T��m��e����, �߿UD{�,��Xt�1݁q��ؕ�:��=���h�q���<.��N�Bݭ��Ln���p�C�u<v����m�?�03�?��ـ}��,Wn�ݻ�l���w��ƒ��T�I$��9�����}��o.�~��@���;��J��3�2��qK��X\� �{v�c���c�t�VǱ�j`���):V��]����+ ������~��͙�U2Tʂ��it����#��9y��@�����ƺ�F5���+l'Igt�n`j�K��Ǳmm��<t�^v#ϨŰNܮq�
��xsrnG�hH�o��u�X�镀{֒Gs�ڶ�+f�{��H��/ ��2��|e~���ӡq�N���ܸI|��~�}�bñ%*�H�!�"�5�r�*�� �����H��"*&�b�jH��c�)�����-��lp��e�D4�����}�4C�zî=�;��Em�)&"�p��2h�iI!�"Օ��<�0��s[� 
/c#��Ɔ������,�3��i2�"'*f
��TP�a��;��F�ՅPY	H��0�I��c�s^������ؒht�B���c�[��h"-jצ��U�[�dG�͡jM��;�f��oF��f�ѱ��v�O��h`L>×�F�BP�w8�a��L� �:tj�2@�b��d���,0c��К����5���a��� ��1	�J�����zЯB��=\ � �8N t�	����(�@����� ��M�;�A�t;��MT�6���@��g@���v����=(����*�i�ݵj�ց�T�\����~�}�b�8�{̒�=��ьD=�w���9�[�]��ny$7v�[z������~V7H�WI�Ӳ�ճ ߽�tY�z���؋A�t΁��T�
	���m�˺^��e`���7�߹��$��L?k��~��.F�v���@�=�t̬:��۰1f9����e��e�IU��hH�}��n��{���g��1���K��AAESD54��DL��H�``*=k�[��^�����k�&��Cl�>�����ܻ��z}� ���oۤ����n�.��;��� �y��v�ݝ�9�i�m�[s<k���Ym*um��M۫�{�r}�2��|`}w�:�T�wi�Hn��}��9�@^z��}�w`b�9����G�5Ƣ%U*�U4�M\X�Z`}�.W���&V��B|Yq4*	����؈�����M����c����΁��T�P)䪢*����1f9�y��@��à}��݁<�n���~~q�Z3����]q\�h#=!p����ۛ� �m���xt5O:گm��Y�E˻98�$D�n�cO:a�:��[!(bk�&�dJ�ln�䛫�Ӓk�u�r%h_)u�	n.��g�ݞ�{oB����S=[��}�펁6�ľ��Q��8���јݑs�g.��vՀ�������fh����14n�΍�����ljz�a%+�k%>�4߾��|������Ӓ�J��]��Y�=�3�lu��s���h��`��,�v\@s�����<���,�����c�^ea�>���v,�= �=]�Z�V]:��w��}#����.�xޓ+ ��$�\�C��`���{�����G!/f�c�|�3�g�B�J�[m��v�������zL�{��{���:Q5N�v���n��&V�ό��t]��o�j"�Bj|�q[RG-��h�.Tq��vI�ثl��v�h�yu�q�����v�ג�Եj�ց��{�����zL�wɎ�5����r�����%U���@:>@���o�r����G@��ào77aj��)�UDU%5_|M����c�^ea�R���������h�C����zL�{�����^�� =���'�GR+N����8`��n�˺^��e`��c\�l�n�֮{>������#�	a�[����w|I�۵�;������Ƿ`b�9�{c�^z���T�m�m7n˷�/t��t��7���7�t��p'J&���Ӷ���ʻ�߸r���~ܰ�qT�X>z�dG#�����Y�z� q"�����ݽ����r�K�>�L���B}j���-4ճ ����s�f��n�:���yf��TGiF���¦�s��o#zɫ�:��g�W�c���p���ч��R5���������&V�������_��[���&������7���>��7@�z�]�Z�V]:���+@�s����/t��I��}�I*:���I�E0V���t^�xޓ+��>D�*�{ñ�~Q<�;� �B�J��ڶ��V�@�}�2��>0��M�$��E�.��鞫#��^��H)�.ۋ6�.���[G[zg�lW�9�a�#�ғ����?�����oy�}��n���/ ��Q�D�wlv�j�ց����t^�xޓ+?�'u"^YJ��12�M[0wO��9zK�>�2��όt���hW�ݻ����9zK�>�2��ό�{���~�d��N�Ht��x��c�^z��{�����s�".��V�Z}��>ٽ̳z͛ރ�A���(���z����
�gn.������rV�:�zh�d;%��q�ϩ�X���޹z�g����jb�ڜ�
�S���]����Y���{ 8峫t����)�#�.�y<]���.N�t�2X� tus���j3�q�j���4mO[����5�mPnby�-0�ZX�>�f��a��jNY�6�ϙ��8X%*��P8�oFoZ޶�z���&Ο#���3\o|�c��\��6��ǂ1<um� z)�)�͑�k�ݒ��-�ф�d�p�ԧ&.��?� ���/t��+ �֒Tu�$X��Sl�>��n���/ ����7���:J�Um�ն�����/c���7����q/�S:�݁�:��4��;i��>�2��>0��7@�{����e&����V���8`{�n���/ �I��~�J����,��-ʶ��m�5bn���{���P[{0\��g�jѻ�{6�dx�'<�P��J��`{1����z��cy����3�k݅�0R�jb�fj���<��s�b3�)(t�9y�>��>�>0�E�KRڤ�"�:n��L���� ���/Ix;�B�1]�v�W�]�h��}�t�����+ �ZIQ�ԕ�aLf���t^���L���� �~���� }��[�ܕ�ܫ�{wn�YΜ��	�h�"H���I���-픢�e������+ ����>��n��:���
�6�;w�}$��>�>0{�7@�\� �����V&����%�p}��{�߹�iԪX�_RJҪ���^E�t���;�R)>)R�LL��V���M�;�"�>�e`w�����t���mSm�ot�Ȱ��X����{���H��+��D�/������a{v�0�.t�h�n.ؒ'�.��e��,���I�J���� �I��}�|`��n���^ N�.��*��K�3ذ<���r31��'ut��X=m56@v��ـw�߹�1y���B^{����΁��ˤ�T��3U54����s��(��9���{�9W~��nV��>��o}w�W�B���:�m�v� �I��}�|`��n���^*�ҩ@���V����=i�ݺ�F��<\����hԡ��v�v��v��l�Ӷ6�j�ց���r��������X}�E>�®�*R�R�:��w{����vz�kN��z���F��Z�j�J�"���j��vz����a�>��݀|��-���Ҥ�i���ߏ�8`w���M�9zK��QR�X�ҫ�h*�XyL�c���c�x�U~�õz�����``
����TQU��I���pW�w���ƅG� ".���@�A@�����������_�v����������������������������}�?-�����T��UUW������?�EU���H**��������G��<������uEW�?�{�-�}���� ��������W!!RP!% DhTIeD��E	Q!eD�HU�BTH �RQ"IeD�Q&TH� �D�D�EEX$ ��`�)!�(F�J@�
 �`	��B%"(B��"�
BHBP&@���  �(F��
Y�!��@�VP�d	��B� d��	U� @�a	 � BRP��  "@��   ID�$
 �
@�P��!!YV@�	E��0d	DB@Y !	�!@�BYB$	$
@�!	� B@�BD` �$BA�e		I	d	�"Q� �B	a%	B�$F�A�P�@�V�Y $R�!d$!	B�eR�Q�e$FP�A�� dP�!V� � Q$ �E$ ��@�HF�`BFe�hP( i�bQ� F �dFPFTD�aQFA�A	BP�e IE�`	�FA��XFT%�dB�aR�%A��`IFAd���a IQ�dA�$@	F�a�eD�` �$% ���!Q�`� $A�FB�$PI@�UF@ `(F Q�e@�P�aD�aF FD�	YF���d�	%�!	$
P$%R�!%P�d�ea@��a@	@�@%FP$U�	! @� B�aHU�RU!@	@��s�����������g��������8���o�**�������A��������_���**�����a܂���%EW�������TU_��s�B**�dg���4l�Ώ��f�:���=�G]QU�����**����~���u���# TU_���**��g�8���!��΍�~����<?���O?ю> �����D����������EU���s^���WW��?o����������d�Me˔4dX]f�A@��̟\��| i@  *�@ U �� (��Q@�%R�P � 9UT��B���	TI	
$� �T B� E    @���)A@(����*�.    #  
�T�@�1 
w����j���e��^����[������w�]5q�ٗ9��g�  �Ҳ�`Y�� ��tw��@6 >� K����q�V�r:#�OGz��n�5�z,]��o07� P{�    	� � �U1p
&��,�G���w)@�h�   t  @    � @   �:@@ $  : @ D   	�  �@  �(�P� tbh����3̓����ھ��O||��5\F�76����Яp ���n9��㛼 -׾��[}��y�n>�w��^]�맖����r9_p �2u޺��y������i� �� (   R�c� �[�K�/=��ʺ㴡� �J�Ԭ���&��ﻪU��J�ܭs|� n�m'��ϻ�m���>��W.����nz���r�ة� )�+�p�k�ӓK��J8�¨�   R� � ��s}�=<����帍��;Ь|�i�yz�e�m�7�n�9�����q���wx�M㷌y���ǡ���iY=/{���������f��>}��6]��ӳ��G�  ��"��*UA���ha��&j��i�42���R�P��2h4�"{J���4@24 ����j��@ 4 DHI�JH�Ѡh������������������I���u����A^�����"��TU?�DU���"��
 ��@ES��S�1�B$X!A�$IDH��lB�hl� ��$V�BH����>c��+�D�1��t�?<����B��߸�<N�$XT��(c�t����sT�kso�'��Le`%e	R�g�),�����4�5��a�P�`%'���A��K^E�xEгW�� D�Z^�%!B$�Jd*E� d�0�a�j.��t�̄��o�ɥb�D�ъj5��{[�@�
h�a?��1��r��5���aJ�(B�9�h?o�pѾ�HJa
a�IsSf1�f�j7Y�ɴ��L4�Ͳ�4}���B�dX�:s�L�B��\�Յع��|�����D�G��$B-I����}7������8rF	9k$H��DK��904²ț,D��y̎��HSZ
��HtM� h�!��TČ�숤-0�T:&&����&���0Ѱ W&ߞ���@�;�/>�2����� �:)� �>����%M!���M���fE��L��v�l��ԛ1��3.�f�L$����,��yq�D�S���kD6p����1���6�$#Sl��P��l�qd��2�eXK����٬֚)�
���FB什Ĝ֡���6?�>�0%	tco��>1ӱvp�#��;8|;6k�^�K��|lt�$(@�0 `��?e��[41�!�B!rkq�[������&���*Q�w�
��F�!p����Ms��S>���2�{Q�D/L4�贬��DT��
vp����b�ќ�}��39���71 O��Ì��މZE��!�,FVl�J1��A�*B�
�+�w�S��9�c i�XӄX�����
-���+�	*�\N�i���������+빠.UWR�W]SW����(J�GV��B�K�A5p��iY�鐷���
S�C�q>u��7¤Vl�h��ͭ]q�¥��Q�*��Y�����#!�%��`c�	�jA"ְ%�XZR��Mc���!��[ B���&��;�D�h!��0�S5�RH��O�*`-7S$!L!�FH004��$�F��MA���P'�5ą�q��7���Z�"m$�fk|���p�Xԅ*��żLL)���D�t�	N�o%I+��p%�F-�{u��aIW�0!s�{"��iH@�@�(l�8���Zk��!� )���$���F����l�P�҄Xe�j�!��[�}����� m֊~`d�B���B�ZH'��?G��	K�A��dvdn$8H��P���LM#$���FH��5H���B�������FIE�!\�/Y:�q���;? Z(L�g]���?�,b��b¬>�af��"4�HS6�m�	�}�}���~�|\�ԛ0�44�����!R8h�'��~8o6e6\�w]չ�Ck��Ƹ1+��8*�
ċ�ג����j�"hQQGI �̮�$d�jQ�g6�/	̉A$�J��|M���8JD�,�qH��~����$C��� �r|fM�����i��$�Q��?~v����S4fȔ�8����1�&ݜ��T�48��|��Jh��� Q1Ӵ����;vp�HP�7��ae.�%��^���%�w4�)��!�хbLM&���Y�U�MI �[��V��
]w���4���e\ Mn�R~�s���e�.����%!v�e��֒�X�����Dy�)����gu��r��+c�"���*����u)�^�� I�8\e���� G�c "�JFB.:�w7��I��W�)�O� F&���>H8�����!Hi�տq��`�!u)�u��E�R"@�1?a\�4h`i�`XBR~iG ѳF��>��!.D�7�m]��n��D1D��I��%�%�\�$C���Q�]9�l.��5��XG4~�cP#P�SN�i����h?,����� ��x�`���k����>�b��8¤��B @�8�������r4!y+��3P�:a&�3�`HA�t���BRG!S	d"y
f�7[�:0���(B�||l۠�}:���dE��廋-j%\e@���ua����>M��>H�s[�)����i�w���kx�8~S5�k	LR%R92}&���A��5�cp��JK��Ըi�.2K��E6JĮ�1�k�"��.F�#
��.V��H��/��(B��XM��̸��>v�i�~Ր�f1����,���HG>���e#L�_�sZ��bK�B�$U�ׅf���I\^vE"��1$ Ձ@�	F	X1_�~���H�BZ���G�'	H�H�%ğ>љ��M����E�їZ1
c	���.��)�"V�/�).Ra�D��\���!Q 0)�����"۬��Me�L�q%XX7���w�ڵMƤn]u%3HK����!`P� �u����|p�A�0���s.K�2�	�ԅd�;��0����u��a��K�� A`F�\�v|fp��߷���{��Q�v+uܓ��{͓~!$��5��ǩ��}&��h٪a�B�PB��Rk���)��VZ����B��`h�s�7�j�n�8��&�0h�hٳ�-�	p�l�������.k��[���.k�}L'��B%r,�4
f����bE�B���DU�O��r�i\Ц�4�ê����Ͼ�}��,`XT"V+!X�+ �2�I%�fV�F��!	[$(��i
��eݒ,T��	�VF"�0��DYw�����d�Y�)4rkF�j��5����}��p�|~ ���Ӿ\����	�1
��� ���݄�oo� �],�# f���i%0yl0Ԧ:��@"2pu6BXF��)w����9$���n�4��Z1 ��HdH�&�l�n��2e����tK��JƄ+� |\�E�l�s��I F&B��))ce�Ki����k�]�~a#����[n�A	�<�x����m��Swk�uH�]�II�H�BT�QП�"�8�o��>�рȡ�ď䈍t?3�JƓ_G0���)(���K��1�l
� a*K�ZX'�!>	_�{��h�i��8Y��j~����h1`A���?euHo�a��s��\����{�et�!W"@�A�L�ω�ː*�BR��p/fA��(ԋꎫ�L�g�nzs�/R'��^�W�B񷑜w~J��aM ���Ԇ����sL�F��.�e�~y��p� j��ĞDJTIF�H�e�Np��o�k|�D���51�AD҂b�,g;�!JT��.:`�%	`F�`AH���b�RcE�R(!�BKb;�a����(E+�J�L��^wz'6��t˄*B����I �)��5����L�uq�B�J�h��s[��39̛�eԖ����F)3L���0X�"�Z��E��D��E^T
aT,B�WhU1#4
ġ���]&�����oJ��\.�}�8��ʕ�e,��9�^Y�>���1"E�)�$�
�
G�-���IO�@�
��lJ$X����	!����d��	 R@`Q�P�ƻ*~RR2�F��G��F���Ŷ�K&��F��.H>�w�w]�
J�����b�`XP$�!J0J���+#.!JT�Ԕ%2=��!����Z��L)	��
1
)'�ހ����$�Ac�A��>޳t$��n�uު|�����K�����	p�º8���w�Z@�I#ǁ�I$�jH��V\��;4f&��l��L���d*E��	�WQ��C��"}ӟ���0?'ĉ?]h$�(@*��Zf���:�A��%����!A��j�
��"�<zk��@��@ � �   $   �  6�p      m� :6� �M�        -�m�m�        @�`   �    -�        ��` H   %L-��m� [�r���[$�[�9��ݶ���'j���%��n�+�mm��˲�2�j��%]�� А۶$ �;5UUJ��T,�>Kr[A� [d�zu�m%K��npI��I�6�とv�&�H�Ƀ�l-���J멕�C]�ڥZ���Io@\��mV��  l��t�s���m�� +J���^e�h�ng�e[j��H�@mUQ�\��[+�U]T�V��n5(8쪹f���9uIS���Ͷ-��ݰ����%��fx�'��R��Q���q�q>��m���Ӛձ-�85�`�4�ȳi�� ���=�q��ͣv�69�e{On[.��X!��]FW"��l�v9o/�@��O *��{E�Yca㚍�� �Q-@8��a�)�I��e���T�+��M�]���3����Od���sP �E�Z�7pٺ�S*���_�U@�]ZE��� 8�CY��� �P��HUU�#ƅ��q�Ze���V����=�ҁs��9��U�u�p=sN����R����m�#��V�kqa�K���0vYz�vV�p�n\°/)R�V�>�:�V���-�A�D(�;�n3-�]��/sVqڞ�va�ո)��ʻ[USm�Ŵ��h��l�-�  �I������ n��$�h[�lݬ�$���8�h ��\��E\���\
��s*�[�g�h
�k�:@ջ*�̨ tָ�WmHm'l�^�jx�c�i+6�[V�#j�:I嚪�˰�PJ��ec�,3v^��@`m�Hඃ���[��p��i n�m� 9#��m��['Sm�^�E������v�UUL�+/5J�ݵ��Mz���@�� @@�>6��-n i0E����ln�I�  t%� m�#m��!t�J�mUU$
�[+�.U��		 m�oVζ�ʐp �im��z��b�*�,��A��t�f��Zl��-@K5��P6�Ԁ  [V�d��[v�  -����� @TU��=J CXn���,�������%����'��UV�m6���A����ΠA�ވV���k�^��m&H�` $ $-�U.��-Hm�(!KVP�W��İx
�z�����T�R��P���  \��6�O�O������%H��['] 6����.�k-�4U��A��.��6�s�q�7m�,0�l��- �vܣZ�Y��;t��Ӎ$�Z���j��@奶�c��l����IɌ5Nԯ�K��rA�f�1[t�]�[�Wn��v��D��gQgMѪ�]�Y�����`�5N��㝛pm:��*�V�UүZ�8gd F�!�Mm��@ :��eq{WV�m-�� �ij�6� Hq�kh i��U ��4��[T�U:إZ�v|���Id�tm��Zlm� �  � m�6Ë]5  �mV��`	n�4T���I(I�<��6ݮ�G+:+8۔ ��Z8 �hڐC�۰p��5�a�� ��l Vꐧe�h�S]�mU��5Ys�2��ę�m��`$�v	7�z5�m� j@��$M�m�ۊ�s�f���M��i����kn�� ��>�[�d���$�)�t'@�̨7WP��E� ���Kn�	gP$�N��l-��6F�a�{��^��Z`���q�X���R�"�n�p��
��;]t�M��]���c��T�u4M������@�jր0n	vT����:�gJ�\�!�Y:ɀF�fY�� � 5�9�@��N< H��ɨm�tkZcH6ۄ���fm�I%� h   ��|}��@uO+uUclAy�   6� ���
�j�s� �<��A��$s����`� �fٶ[��ɭ�'�i$6�D1  �m&����H�  5�닦��$�k� F�&�l�v�*Khpi6��������`  �M"��`6�7� ׭�^�  ]W$fݶ݁:Hm��v�`.��%���\#���*m��ms�mUS��UJ�� �kj���Zk�m����(����MmR��ʬ��ͫgI��@h�m$� I����[�����ƗK����  �l��a���+��U`((�]�m6�ޠ���@ �,�8d������.�UJ��Yv��Y&�L$$��  �`�	�(zE�5��ݭ��M�K�$�l��G��pumD�(H�Vî ��}~� Hg��`� ��&�v���� �Ɇ[p�]�����l�l�P  �m�l*{gm& m��m�K���{]s�ܭ�&Q6.��@�s���<b���[�q�(��ػP��H=r���r�f�SɌ҇�Q�R�Gd�-���X��<�ܧ0[UUZ����4�嫒H	4^���g���H�u�6 �      ��V�10H/-�U�ݵ� H:mwd0��P  -���h�bQ;2�i6���[�,,��� [BܒV��6���[V�m�[E�p K[�      [M�� mm ���  6��6ٶ�2-��M� $6�ݶN�����Ȱ5�$ 
S��m�&�KsI��8R�u� 7m���6� ������-�5u��   ��    �n���m4P  �[p�hkm��`$8� �֋h:�I0m�����>�� ��m�඀     ���h ��ζo��ﾐm��D���m�l�m�!�]%\  m6v���K:�¬���Ĳ����e�t�H   l  8��   6� -�l	���m�  	   sh��  @@     ��p  %�ִ���$  mk��v�m9���}m�    d�hm[@6�  ee媀��r�UA�� ��      ~� �Ә�`  6^���ͷg  ���d&�ۀ M�	4UmCv�p �g6ݩ�N���r��[V��m@UR�-�$�5�1f�Ԗ� l �09�n�N��%���7mq͒:@����5�ѱm&�J+`9` �f�%mzsm	��c��:)�����l��r.zS�U�Vm�yU�%���U@@MS@I�`  �f���ݶ$ ;m��۱�    $ 
�yeeZ���'U\�Y�l �$u��  �p� ۶��l�\ 6� 84�kj�f�T	疀���RඖӁ��   6Ͱ A� UJ�H5ʵ�T�!Q��  ��Im��Zdm� �[�}��]-�Z��6�[dXl��m�-������m�$�`  ;�[]:p%�k�*��nV��8�[եf:�i -�۳�6ݭ�  �ٵӁm:At�c�Ŵ�-`�඀�u�"�!m8}��햘06��� �xP�o�ճknmSi2$� ���d�{I�H�v[����AKl����/�} �n��Y���ɶp��%@k�&��#L�i�@H\�HZf���܎�:d�kh :�۲����;��`�-`�m�5�
Z8�T� ��ӛ��vN��(��@˴��N��Iq�t�yz���EU �D�c^���ж��ڶ��m m n�&�����ki7���cmo]�l[@ �m�� �n��Ͷ$�I�6�@�  C�@6� � F�]�ЫUVVZ�p$vǆ��$ �ջc�%�mm��V�bθ�	�"�p ��2� ���tV�e�J��b�`k�m]uV���*UU�I�$Z�I�D��m6���'M�I�&�7Md�h-�2R{J�t����f�N�3�si:W&]6  m:��V�ڞ��	�Up�D��  4^m��f��ʵT��/Ҩ�knץ������m�nC�@MM,W2�T��gir�� m��Xm��d��U��r�%����y'��i�=v�P�+g�T�#��UU�R ��hP�63*�UUT�SkĞE��f�8;n��:��[M9%  -��t� A�$4S��Pa�[�mJ�`;m��`�#EA��_��p� l lm��� p�c`  �Jp80�m�lm�[jf�@ �  �,��l l� m�h�R�PU���v���l�UFEBA�t�`�[��  Ͳ4f����Z�%3D������b1����?�a����C?��W��Dq��@Ȃ��*|V����b�Au�� ���D���\@P7�~7�?|�ȁ�v)�?�~T�E7��Pp0�J )�,�&�1 �Fr��lυ?$E$F"$~S@.��W����C�G��T��S�|���@���i�&"��=H����'�@8"t?%��t����P�*| .πv� +(�T0 0�P��A�?c��P�/U-TB��������=��� �#����t�� ��054:~x�F)�Q���M���QN�zb'��~O�a��u���Ž��T�)p�(�Wg�Hq���T~QE���%^��1Mp����A:l/�z:�&Ȩb|*�e��:��> F �0L�Q!G�pS@�W��Ez��4�56u���_���GH�:/�~W��� ���"��~PWhH;�D?}����]k�"�<Xi�@`@Db!��TT���"����	��	D�Ab	b,QJ�B�E,�`�@�V ��E�Q@��_hֵm6�l�m�� ��m7am-Mxlt� �[v�K3UG�VK�k�� k(N�+R��!��bG�t^<��}����"yN���j�ўS�)
�2�F'άvv]le�u�.qR�����}�[m�wA�ɚ���z�!EմIu�z��]tre�8k����8Է0QjR�eS-c��̭y��Ύ=#gk�h
�Un����c����Gc��ji2��uh
����a��e`�:&��TP)�jZ�eZ��Yx�a�ݓm�6�C4��OK�Z���ͯb��Cүt
�@��Pj��c����EX{��S���'\��cLv���9z^�<]Z�Ҁ3�ںx���VY"��I$)��KN-�� N�9C]�⣭�̺.�GnJ�
-T�r��v��b���d���ܹ��1S����ۄkuv��Ov��l�jzH�0Qs8lfs�G��Pl5��VWv[���ˊd����M�oe�5n�	$	��H]�E��!�e��K�+�7o=��=���G��v��f�F���0�Y6���8^ݎ�qn-9N�Ik�g��2���OKU.��m������mq! N|��C ^�A��M�bԳSv8-� :m�f|�A��#�J���dm�`�/�UV�@x���A�4h�Z��s8�T�9���qp[Yl��m#Ui�d���֍&��6� k�m�A�^-W�Z1jC�v%��9y�[�|���v.˲1��2���c���Tu�l �ts�4��e�ʓ�\�j�Uh��gK�5�!�)�[T�exwF卨p�7c�[�)���&`4�37l�S�aE�r����=�5Y�T8���e�n�Ѳ��*v��@��cm��%Iۂl������8Ϋ�FÚI&j��!Z�/�Pr�x9!v�<��skm\gn[N `�%�=�f�ئ6�z�݆����ݚ�G6�E۶��j��E�Qyt`��7Ră��\p<�*���ԉ���3]� ���'��9�LE�����A8L0�^�(~Q��ۿ�xם��v�d�;v]Dp�頧��\;�1����g���G��FK�&�&Sp��u�S�g���`t�`䎈]W8m��;W8}�g��g�Ź�&�i�\���h�8=sv����0Y�(�	U��u��i]�p�q����G�4q�Y���h)W�>�T�����u���v�nR:U�����]�Э�0g<���ѢJ��5����t����e�.Y�2e@�&��`xWr��g<���v�Lc�^w*c}4u���`�Ł����:w�`a\@G'	!9J�ϻX_��0Is�[Z�_se���j���.r�I�d������X��K5���V�+M��["��$�M�4
���m��=�)�qˆ�k��E�1�m`ۏ@����Қ�\4��%���v�ЪUHnJ�5\ez��A� �9؍���%��=�y�m�1/d∲��E��x}gƁm�����w4����H�LM�Bw��I�?�pj��Ɇ� �W{�n�s�j��;XX��)$r�(�)�R,��%���j�M�r��7v��yLm����<��8�m�ߓgw+KwkQ`u��,اNG�69!'3@����m����32Ձ��\����6!I��"�N��ܕ����>@�Z��5���Kؑ�G$4l�h���۹�{zS@�u��B��M�4>��wvX�����������:�0p�c�����m����4�0��T� "Љ�!d�DC�������� �jm�͓q��#��{zS@��Šr�נ^�s@������$��4�ڜ�[��x�}l��`���n�A�˝&|Snܽ��D�l���� �YO�k�gq�[ur���f��\}���� |�,_[0�ڜ�I����&�y	q���ߒ;�>4���Z/mz�SbU�I!'��v��3�1;5q�}ݖ�����i��Ĉ�29!�^v��9{nnI����ɏ��8"`Y��D��J��Y`f�K�R�:
�����n����5�� }M��>���������ۮuy:��&��2�sr/Y�kΚ��)�:�I[�xβ������]���ґ�IS������������9��]��@��b�"AH�2,G3@��� }M��:u��7�p�)R����$��4��Z/mz|���4�ύ��q�̿�8�m�&-�N��3vՁ�v��>ɘ����)�4Q��O!#�=����������ǀ���:�`(KУ%	R�����BۤEG6��J���
b&0�(R��$PH��$г0 )��Q�)��������[;v}/]���%�f^���v�Ґ9i�,AO,�-����W;��`�z�5�m���m�6e^˪w:ø�F��bJ��ɹwF�Ў�a��a����I�����l�M���Ylv��J��g<^s@��[J�J�.7���ݫ�"�:6oE�a�q����m��j���1e-��r��7����[��.��H��/'&��Z�a�50�d�&��695���j�s���p�1{��u[��96Gg��Mj;	�p�'#V�b�����~_� ���:�`���=��+�Hj��T�����1;���}ݖw>��=�)�_z��c�$(���ŀt�u�k� �����S�t��]k5l̗Y235���A"�BB��W|�Հ{�m6� ��^�_n'Q �K�s4oJh�f'`u��,��j�Թ��n!�� <��i�5צ��y�.W��˼�g�D�q�;c����k�)�Ǒ8�D7 �7S�1��,��kR���ZXh'�?��<��Q7$��
��������Ji%)+��y� �u� ���*Sx�bm������빠^�M0;�n-�mz���M���%QB�a�s�Os/K;7S�1��,o]��mL�#a�df&��{3�7�f���wsmX��,�� o�}Y�\:v��8�|��]�M���6m(����-F-��S؛W1��
jp:�`���u� ���u.%"��1�4��=�w7�߿bF��;7S�1�2X}��b��SV"�UZ�7� ���0�%���M%�SW��wsŀ{�h�I�h��$QI�z�ŠUmz���m���1�vHc�1�(��W7X�x����;i�8I�)t��3l\�p�m.��U��{+é9Lݮ���j�[R�ϱ������RS������7� ���[u�=jҚ�<D*���+32��I�;7S�5��>���s��f녉�g�'$��^}�@��z���z���uz�N HƦ&�s�WZ�o<X��`4�F/)I)"�&&85�ه���b�=W��I��q�grՁ�����3�u;s%���<�c�[�G�y�Q|��
�..�c�Ԇ��.���2�3��Y�Pr�k���7� ���y��5�ŀ{Gh�,e"�J*�N�X�f'{Ē�q$%�$�#���׷����ڰ3���ԫ"�d��<��9$ŠUֽ�Қ�w4�ۋ@�J4�:��m�����빠^�s@󝸴
�נw�&bo�"I`�������S�9�� �� I�֚���e#X��s��X��YY�&�t��v�<v���+�.p�TQ�\e����:�M�K�|6�����p��q�On�cS�����8�,v݇m;�۬�9�v��]�N�h�F��^vs��S��{�u��	��tE�N�лr&�Xv��۩"zֻ��Р.�6�y�Z�N|�n��5����e�n�'�f��8箮6��i\M���۞6�m�=[jg��~�����a�$<�������������F<I�t�Sj���~������u�@���h���<�u��"�$�s�WZ�{��oJhs��WR��Mb�f��{�偝�ag�o웩���,�brd*'�ő�h�S@󝸴
���\]l��<��<��A�!�h�3�7�q-�ݟ��fڰ3��,)\�j����N�2�LR���݋s�e{[��>�#Zv	C'3n<�h��L^x�Ut�Ԓ^�_3�J����w���~�?>���� ��.
r�:�Lݷ�g{�|s�� @���$"�a
6�J�ӥ�]]w_j5$�{-��%WJ=I%�������HC�y�I^�Q�$��n/<I*�Q�I+���x�^�W��l?,����ԒW����$��G�$�[�y�I^�Q�$��Zh� H�9�M9��J��z�Kܥ�g�$��u�J���+o�A���s2�kD����je�e�O]g�.c�w��5�ڸ^0�48.6S��	���F�?I}~���Ē�.�RI^���Ē����]���d��!�ᙣ�����wf���������[o�u��K���}�y�Iu>�<y���$MU2�m�k1?ߛl��m��RHZ��$`��4C[I(�����f!V�KS�X�T��A�`EZ�I��Hb#b�������'���{1��؎�P�P~���ϔ5�\�������*?'�p�8���F��HZ��c	�HIEx�������8����^�vF�:�[��	�S�Ԕ�d#v�s��?ZЍH@���� ��blqW���B�T�Mt4&�C��D|�&|U2 ��Q0�]�'�8r*��U�;t��.���r�w]ݛ���U���_�HE$�b�Ē/JMI%����~m��e��{ĒRn^��6�^�4����n8�p��J��g�$�t��v�{�]�y�m���˻m�3��{��k��^�c���a͸�#����o�猾�
c$��7=�J�g߿�%l�Q�$�Kqy�I�&���o��%�z�F����m8�I%z[��>IIݭ*�m�n�_�6�{Yl��UM���g�@c�$Ә��$��|MI%z�3�K�]F���-��%U�J84q�,i�MIV�[�y�I^�Q�+{�]�y�n4k�[U�"�Bp�(�^c/&ff_r��E�WB���r��ͷ��������ܽ?~m�;XU���{su$��5f�F���n"b28�rtZ�⣓E��7nK���7/c�\n��)`�����xD@��E�F���g\^x�E�I�$�[�y�I^�Q�$�*�F�X�<��I$��$^���J��g�$��u�J���}���}4�Co�'&�������%�.�RI^���Ē=��RIyr~ElT�S'3�K�]F���-��${e&���o��%���a�d�6�F���-��%��^�������}{���m�Ԧ4����~u�w)v���fp���W��F����6$��&#3DS�b� =�s�m]��Wl{C�޷ng�{;BL��#<\n���_����|sn��in����c���ok��wZ��u�7���l��"��!���n�60;t$�g��`y:�ܣ���g1l6��Tl��W/�ݤ���QT�ɤZ�tbk-�����QҖ�7{�����}�s���|Z��;U��	b항`v�o�o?y��rsv��{$H��N�`�svn^rI��5$��|�<I.�u�J���$�V'&6�BKnRI^���Ē�Q�$�Kqy�I�I�$�{[Iܑ7$ �73�K�]F���-����6��|MI%��Ǟ$��t�Q'H���KΖ����l��Ԓ]n�y�IwK�Ԓ^R�4jŋHE$�b�Ē=��RI�����RJ���RIy��^x�U����a�(�,�tC֋q�JFn���t�x��`�Ƴ�q��#�����,o{�x�q8�<I%��ǟ�o���[l�Y��.{��i����v�o�U�z(�Ԫt�:�����fZv�J���KWv�����~m�ݭ�m���o�_�}�Q�7����x뜦f7��~��ޙ�5�/&D%hP�]�7�
=���6Ӷ�jǣ��`�
R��W�$������v�x�]��-I$�ܳ�J�
�����BKnE�$�ݧ�$�s��RI.�,��$^���K���>�%�����ls���i���ܠ�;���s�t\J`w\!̥l�!�Bẅ�V����Ē�.�RI.�,�Ē=��RIu�O<I/h�'��N2(5"5$��r�<I"��jI.�i�J���I%�*�G\1c	0�M�y�I�&�m�����-N H� 03���g��	����I$��I�%�p����x�qH�5$�^�y�I^�qjI'��+��߹;[{�����͊=�Jt�J�����fZv�o˜^���Wz�y=^����v�������S���?(�NI����V�"�4�mm��]�����;����=uƣ��|���x뜦f7� ??���_��+	m����5.}�m�V�-�ޮ����6�ITW�ͷ���_��U7�����m�׭��m�3
��R�9Ĥ�����l�c¶~ ?��Ͽ7����[-�\�9�)#��+������[m���b�$m�G27!�/�g���n�⛶�{�zk��߯uٛ��
����-b!�
�?��Р߁�P-�����[o}3�\&��"q�A��$�[I�%�����?I_��y�IwK�Ԓ^:2� y�$h%�;��v�K���q�zҙ��{lC�v����="�L�Y@�nL���\��'�$����K�]F��]z��Ē��A�N� �R'�$����?�?�%Sݯ[-���o�~��9����������_Q�LX9<I+gڍI$�����m�|����]��Ē��^��4~Y1����/��~�d�Ē���=I%�����o�U���2�m�7�(�����jIJ�~m���r�m��I{����z�{��e��}��ߛo8�0a �d�k�4�+U�z��.����6��� 0�E8���`x+Pn�Y'����s���l��э1�xN��".��*�a^�qe�c��1� ]p�xސʗ������n�^���u��=���$l*��I��nh��ɺ��Q�U�hrE)Ğk�199��ݧBX����2t���6I�\v5�8��=*���n2˚4f��>E@٭��u�Hh����2��]]�4�y:����x6:�s���N������ѳ���0�������m����m����j���뛮[I%�V��$����A��<�	w;�ĸ��/r>qq(���U�ܞ�;��,8��Q'�h[I�y���+��s�-�U�T�y1�� ۄ�<�ڴ�)�{��>į�|M���ǉ��O Ԏ^��>]��� ?�������)j���<�跭��qۉs�vX�ל<=Wv{�6�����Go��|i��`�k��o�������<��hzS@�gs��pbj�$d�N�;��]�k�����Mh��2�֖��������֖�N��f�݊5t��(�ITU��v��;��,�8��̛�`�x�>�1�T�P����%Ǜ������`�¬5���v��MR�RDG27!�{��������=������a`}�V8��n�QA9M����^����Iǖ�ޭ���8���������~{�}l(�PS�
tGT�����_�����~7+Os��}ٚ��֩�r��©S�䢬��ʿ%�$�8���7�^,��; �f{�٘c(�'5S��E)�����0ms�*K��˄�T�\\^��	�x� �7�`~�N3'
��M���$��f� ��*�?}ܫ�y�zX5�&����	u)�6��>�;�������ɵ��g������V�b�FL\4K��al�Q�����_<N�O����N�68ܗ%*��~ �^ϭ�����z@}�4~�ɧx���iɠu�K�&ϻ7]�f�`}ܫ�q���f�$Q� �����z��i���!���}�����0A|�NT*�nT����wJ��6��k
�$I
BC (b� E!��+F�H@�Ɔ�I�!FI�is��ɕ[�`ncEiJ��QM�rQV��ʰ5,ܽ?�f��aV���nr6Fr9hc��
@mV��u�K\��\�TvmkxS�.�{��Mg�>�X���UW�3r��?}3�w3
���������E���*�EJ,�L�l��zU�w��`w;X^�Ϟc���&5J8�S��Ҭ��ʳ�ܓ}����M�3� �����E%QV��f�7+K�Ӹ�=�7��M������_��@�Қߖ�� }�x��� �o�B�	A�0D�s�*w���n��? rBlB�WDH�$�B,H�� � D�#� �b�D5�`	B#4�ܿ���~я��D��2��q�cP8a�7G��@]1#$��L����b5	��?a+.���uv��"A8��D7�Ha� ŉA�E���B&��W!��g�p$#3�b�#�f�Р/L��Kh�\@��x���F00X)���0F�3�z}]�]���;p�j��b��� �6:����q%����sI	f��	B$M�������u�������y`(
��-�� $Uѵ��m�N��` U�­Zl��������ܦ�њ��	�Q�p(��xĶ,�:�Ëg������7l�ۅйD�T�j@Ql1�A�kk���vXu6hj�\�q�8�㙋�()���p��%M
I����]thݷ*��۴c��Pڛ�Ȳ��ih�MY9��1ƞ���1p���5r�O��Mj���	�esԙL\�2J��MT��1z�m!lm`�T�[vB�I�f��V�K!WU�]\v�u��ʘ� �[��`@2�8�3�Qϐ��ﱯ�C�+�n��v�\FV{ܻ�<����p��<� �즴�+�4��8	F՝��A���[���X����YG����]�ɕP�:�3]��l6_��7��vʓ`����=�ϡ@6^ny�qƧ�6�;:��[��ha8i�l���p�Gkh�}�v� 5�YY�\�r9^(����ع�s����$��U-��a�������L����\նқjڨ{��s�&Zq����^��^�j:�l�XF�jr��KB+R�Fz7Ѕ��ё����X��xb(M�`�
�S�<���Gj֧:���]�N۲��c]J���g�@�v���$�y:m����2`��925:�6��$��M /Kȱ�T�Ƨ\�n�ݐoUa�'nҲ�Ͳ��]T��T&v�-V�r�ٹܛF�R�R�m�]�{X�i�u��J�\mɌC�gI�8W��
�͹�1�t�Vu�Um8���N!���면��f�T�/�&M�r˛��[�I�Q]�Rv{n)������eUm��e�x7	Ӏ;�B�2�]�*��uE<m���'��vm�)�5�]N�s$� �Ù�VΧ��t�f��v�9�t�F��O�����	��k�vˉ��Zl�X0��N�����Q*��Cfڹ�`�۝M��H\��gK�@��A�K�<m!5�i^T��F`rg���o{����89��. @8�y����Ӧ '蟕��lE�.�>u1@.pԙ3'�5%���3F��n[��:r�A�zF�����b�Z�uv���t�ö�Au�:˘M��Ehƌ�v�U���I�n�a���E��ͷX�f�Ù���b�Us���=���e�ۭ`�GR8&�ݳ��YF��h(�Wl�˶�dM��Szў/�,\�cx�0��U�q�p:40ْ�y��e7]��z��^���x��k���/�w����wsK��ʷ\����"Q�nݶ֧O'=���蘁;=�s��!y78��S� ��m�C@������@�U�u�Mδ���"s#q8Xs0��K��d�vnV�����/�aPcń�I��&��>�@�Յ��%ēfV���V�./�31�<x��Q'�J)�~��@�S@;3
��ef���k"��q���%����5<�ҿ�L�`w;XX#�|m�&���F���)�sc�b��ؓ�`�Wc[�ҙ�tA�����}��c�IQ�7t��gqټg8�r���`}"X�'�{�iȖ%�b~=��欔�Iuf���ӑ,K����Ӑ��H� }�F�Uh3��P�ț�b{��&ӑ,K�����iȖ%�b^�ޚ�r'�"dK������i�55m,�sWiȖ%�b{����ND�,K��~�ND�Bı/}�Mm9ı,O����_�&q3��O�uS�)���$��-9İ���ߦӑ,KĽ��5��Kı>���K��dO{��iȖ%�b~������tj挚��fjm9ı,K�{�[ND�,KO����9ı,N����r%�bX�w���r%�bX�=;��r�W2��	��q����f�v���w�+F�;v�[���%����N��g<v��mm9ı,O����9ı,N����r%�bX�w���(@C��&q=��U�~8���&qn�,��GRᩗWZ�ND�,K���6���bX�'���6��bX�%�魧"X�%��u�]�"$2&D�?t�g��f\3Və���Kı?{���ND�,K����ӑ,j���FA�E��2'��~�ND�,K���6��bX�'���'����ѓ2乭�"X�*1Dș���魧"X�%������r%�bX��w��K��A[���M�$S�Ӿ���K��Va��MlI�9��t��H�b�o�vm=ı,O��siȖ%�b^�ޚ�r%�bX�~;n�&��l;���g-'tM����b� �>:�]�e�_chp\r���?_f�׋�8�1���ı,N����r%�bX��ͧ"X�%�{�zkiȖ%�b{;�fӛ��Os������F�\Z\���"X�%�����m9 �,K����ӑ,Kľｭ�"X�%��w~�NE,K����8h��5���kiȖ%�b^�ޚ�r%�bX������Kı;���iȖ%�b{��6��bX�'�z�y�fMjj�e���ӑ,K?�dL�������bX�'�����Kı=�{�ND�,����!v�c ��#Ră
����ͪbBQY��DW@��>Ͽ�����bX�qg��H��#�⡪�U|_�&q3���w~�ND�,K�����v�D�,K����kiȖ%�b{;�fӑ,�g8��̊Dk)S9
C*�y,wsc��-�ק�r������ۛ��|c���̹�d�jm9ı,Og}��r%�bX�������bX�'���m9ı,N����r%�bX�g�rz[���&e5sY��Kı/}��r�bX���ٴ�Kı;���iȖ%�b{;�fӑ,K�����Ú�R�%՘ff�m9ı,Og}��r%�bX��w��Kı=���iȖ%�b^��5��Kı;�t��f�Ѣ�d��ͧ"X�%��w~�ND�,K��{6��bX�%��[ND�,K�k��ND�,K��{��*�
��UQ���/�8���,�͖��bX��3���5��%�bX������Kı;���iȖ%�bA4��;��\��lԗRB��Z���V��I$�sm�Iy���(�{�\��6.7�N���g�X�6�wMu��'nj��������0<�KY��-t���ֳ��w�l�Œ'���k��An��n̶q�uN�.ǥCy�&��k��iٓ�v�ֱ��W�/h��<�n.Tt1
q�{Fʽcɮ	8݄� �m��v��m]k�#�k9�8��$ߞ�wu�����Y^��h��#�[7T;37c��T�lss�Sru��3+�<�2�J��
�MʛŇ8���'��*�r%�bX�{]��r%�bX��w����D�K��w�ٴ�Kı^�h��B�UCU�U|_�&q3�����Ӑ�9"X�����ӑ,K��w�ٴ�Kı/}��r%�g8�u�H���NB�*_㉜,K���6��bX�'s�}�ND�,K�w�ֶ��bX�'���6��bX�'���&x�-˚�V���r%�bX����m9ı,O��{Z�r%�bX�g���r%�`؝�w��Kı=��'�nFD����fӑ,K�������"X�%�?�������~�bX�'�}���Kı;����r%�bX�=җfId%�]Mu-�շ9�Ň�5���n>;v���%����;l�rF�3�U0i�2QUU_��8���&qv{}6��bX�'}��m9ı,N���6��bX�'�ｭm9ı,N�]=��i�tj�Y�u��r%�bX��w��>���&�X��sٴ�Kı;���kiȖ%�b}��iȟ������;�ow��������K���m�"X�%��￳iȖ%�b~����ӑ,K��=�fӑ,K�﻿M�"X�%��wĸI�F�5sR�iȖ%��dK�����"X�%����]�"X�%��w~�ND�,	�S"{]��m9ı,O��Ro'����Z5M�ֳiȖ%�b}�w�iȖ%�b~�w��Kı;����r%�b����mK��q3��L�ͣXl�Ut�l��;�OO����F!�A�\�x�1�nvCX4v�<���9�B�:�����{��'��~�ND�,K���ͧ"X�%�����fӑ,K����ӑ,K����<e�2��njm9ı,K��{[NC�#�2%�����ͧ"X�%�����iȖ%�b~�w��Kı?���s'�-�B�X\���k��Kı;�{�Y��Kı?~�}v��c�5$9��y"~�w��Kı/������bX�'��}fՒ�]Y���j�9ı��w�iȖ%�b~�w��Kı>���m9İ?�T�Tȝ�����Kı?���YsT�a��f�֮ӑ,K�����iȖ%�`����ͧ"X�%������9ı,Oߵ�]�"X�%�������.��L��Fy%��<t��IZM/���\����ts,��೘m4�e.:�o׻�����d����ͧ"X�%��u��iȖ%�b~����^D�,K��~�ND�,K��p���S4dְ�5�ND�,K�맮ӐKı?~�}v��bX�'���6��bX�'���ͧ �%�b{��6g��ch�5���v��bX�'���ӑ,K�����iȖ!bX�g�{6��bX�'��}.ӑ,K������5��\ɩ�W5v��bX�'��~�ND�,K���fӑ,K������K��ȯ<�"�������r%�bX�1��I�2˙sV�56��bX�'���6��bX�'��}.ӑ,K���w�iȖ%�b~�w��Kı?��������/<��wn��6���z��˴vvέ����ϝ/�Ç��G_��?'ۂݸ#p���>�bX�'�k���r%�bX�����9ı,O���lD�,K��}�ND�,K��޷j�K.�ɗF�ӑ,K���w�i��bX�w���r%�bX�g���r%�bX�w]=v��bX�'���sP�0�m.�֮ӑ,K���ߦӑ,K��=�fӑ,�XdL�����v��bX�'��]�"X�%��=�K�ե3.�j�5���Kı>�wٴ�Kı>�z�9ı,N��}v��bX�'���6��bX�'}�I�$�T�9�Rfk6��bX�'��O]�"X�%���ߦӑ,K���ߦӑ,K��=�fӑ,K��*l���~�~pc���w)�ȽJ�t�S���D��[�:�\�^$zX\Ԙ�Fp�e��A�;����[,r��
kX�!�����UNN!=��/n��^ӌ�.g+�����h^�v�L=��K�ѝͻu	F�sfM�vВ��H�E���8�ȩԈ����9�߾��؆�-�ݝ��j�s��n��j挱���z�u\p�,�w����_~�v���<M���Z��ֳ۵]��㑽��me�ΎS��Xc[rx����q�}I�]��\�WiȖ%�bw����ND�,K��~�ND�,K��}�^D�,K�맮ӑ,K����)�d�˩��SSY��ND�,K��~�NA�,K���fӑ,K������Kı?~��6��bX�'�{=�g���]j̶�ӑ,K��?{ٴ�Kı>�z�9��,O߻�M�"X�%��{�M�"X�%��wy=	r��V,�kY��Kı>�z�9ı,O߻�M�"X�%��{�M�"X��C"~���iȖ%�bw����g-����̙sE�r%�bX��w~�ND�,K�{�M�"X�%�~��kiȖ%�b}�{��r%�bX�����;���!��9��8�+����^�<��@V68�'K�ۙ��]�n���������}ı,K�{�[ND�,K����ӑ,K���w��,K������r%�bX�g�z��l��E&�j浭�"X�%��~��i�b;�!��5�i*):�U���H��ȟD�7���ND�,K���M�"X�%�w��ӑFı,N�ޓ2I�F��sSR\�m9ı,O�w~˴�Kı?~��6��c��"dK���[ND�,K�w��6��bX�'��o'���4։��\�fӑ,K�����iȖ%�b^���ӑ,K��;�fӑ,KlN�^�fӑ,K����3\��f[���Y���Kı/{�kiȖ%�b��{6��bX�'{�g�iȖ%�b~�w��Kı>?t���0�Yu�C0z���u\0\�sr�xzuɛ�8����i.u���{������*5�������ow�｛ND�,K�׳ٴ�Kı?w���(��ı/�����"X�%���{/�%�B�X\�Y�fӑ,K��u��m9ı,O���6��bX�%�}�m9ı,O���m9�,K��z�L���ufkWY��r%�bX�w���r%�bX������K��ڝG�9�F̩�]����;�!2$֖kD��WZa����u�MSP||�U`�\|��_�?������ ����k9�W$b� <R�H������B!�	��&� ��QB��3����𕻇s��_��S��O��DR���H���H�:��M�e����5�����"!A HΞ`|��l]�+���ߗ����Y�G��Q��H?"#�C��G�*~P���%O�OD�����r%�bX�w^�fӑ,K�����f��0�-�Z���r%�bX�����Kı>��ٴ�Kı?w^�fӑ,K���ߦӑ,K��g��5Jd���.����Kı>��ٴ�Kİ�׳ٴ�Kı>�w��K?�"{�_��iȖ%�b|�!���Ĥ������8fΧ��j��3ls��`���\U����l�y7��v�G9x�D�ߞ��{�K>���fӑ,K��}���Kı;�{�cȖ%�b}�w�iȖ%�b{ݦ�{Z�cMh��%��m9ı,N���6��bX�'}��m9ı,O���m9ı,O�׳ٴ�Kı;�n��k3Ym�R��jm9ı,N����r%�bX�g���r%�bX���g�iȖ%�bw�w��Kı>1�<fOa2e�ՙm�M�"X�%��{�ͧ"X�%��kǮӑ,K�����iȖ%�2��;�o�iȖ%�bw��CЙ�����unk[ND�,K�׏]�"X�%���ߦӑ,K���]�"X�%�~�}��"X�%��Ą��r��<m�ٻ2�[�s�\���Ɣ�Q�x�팃�i(L��ݥ�#lFT�>�~�X�%��w�6��bX�'}�z�9ı,K�w��r%�bX���z�9ı,Ow]=fkMsId��Z6��bX�'}�z�9ı,K�w��r%�bX���z�9ı,N����Kı?�Ǭ�R�3D2�˭j�9ı,K�w��r%�bX���z�9ı,N����Kı;�{�iȖ%�b{�<fBpѪkNjh��kiȖ%�bw����Kı;����Kı;�{�iȖ%�b_�ﵴ�Kı=��y3ڸcMh����j�9ı,N���m9ı,?�>�����}ı,O����iȖ%�bw����Kı? �6�C1q @"$LD� b�j�A�!LȬOw;~�1��nM��ZkH�u�c^�N9 H�38ќ�+���G��qy@֖�`3J��OX���ۇJ��&��ZL��j�\��.�<��Rc�]1�y�sgg��b�T����ę�9rZ�]�3�#��]�fNĶ�ȵU�c؎0��[Yx��:v�;I��9k[���<#��8��śg�"��m�����R���zF�F�2`������{�w{��[�:it�n�c���׆�׵m����7iV��;W;�. �Y�qb�p��N�S�,K�������Kı=���iȖ%�bw����Kı=����Kı>3�|a��ܖkVe���ND�,K���6���c�2%��kg�ӑ,K���ߦӑ,K���]�"X�%����_FfR����&�WiȖ%�bw����Kı>�w��K�AHdL���]�"X�%������r%�bX���e��e�$��3.�]�"X�%��{�M�"X�%��k޻ND�,K��}�ND�,K�׏]�"TȖ'���.��jK$�k56��bX�'����v��bX�'���6��bX�'}��ND�,K��~�ND�,K�u���ʷ\��]nc�1���mjq����a:�䘁�;,��3���9����v��bX�'���6��bX�'}��ND�,K��~�ND�,K�׽v��bX�'�t�r��SZsSZ�5�ND�,K�׏]�!@�@�X��(����K����ӑ,K�����v��bX�'���6��bX�'�C^&zk1�Z&��SZ�r%�bX�w���r%�bX�����Kı>��ٴ�Kı;��ӑ,K�Z�lOG*�����%���g�'}�i7�O�{�ؒ	"~�N�7�=��~�ND�,K�?G��ɓ5n[����Kı>��ٴ�Kı;��ӑ,K���ߦӑ,K���]�"X�%��h��;���쑸v���a����n��R��\�4���� d�ٟ�~���S�$8N�ͧ�,K�����ͧ"X�%��{�M�"X�%��k޻ND�,K��}�ND�,K����s��fIuffhֶ��bX�'���6��bX�'}�z�9ı,O���m9ı,N�ǹ��Kı;�t�˭8fY�&��WiȖ%�bw���ӑ,K��;�fӑ,t�� �SZ7��{s�iȖ%�bw��ӑ,K�wk�UQ�%"
�*��㉜L�b}��iȖ%�bw�7��Kı>���Kı;�{�iȖ%�b{�O!8h�5�55�sY��Kı;���r%�bX�w]��r%�bX�����Kı>���K�7���~?O��ċ=���W�B�\F/<�D�ks�+��&v��mn�.�Y˹y5<rMjM\�L��}ı,O��}v��bX�'}�z�9ı,O����yı,N���6��bX�'�{p���Թ-�R�\��r%�bX�����Kı>���Kı;�����&D�,O�׿�ӑ,K�����&L.&j\�3WiȖ%�b}�w�iȖ%�bw�7��K �,O����9ı,N�^��r%�bX�?{~������3)5��ND�,[��M�"X�%��u�]�"X�%��k޻ND�,�x�?A���s�]�"X�%�����nr�nR]Y��3SiȖ%�b}�w�iȖ%�bw���ӑ,K����ӑ,K��o�iȖ%�b~��w���$�!I�IlѢ��.��f9���v�]��6�K��$�%y�.��&��WiȖ%�bw���ӑ,K����ӑ,K��o�a��&D�,O�׿�ӑ,K����O�Z�R[�&Bh�kWiȖ%�b}�w�i�$r&D�=��o�m9ı,O�׿�ӑ,K���]�" eL�bw��rI�F��2j�V�ӑ,K�������r%�bX�w]��r%�bX�����Kı>���Kı=�����I�M[���ND�,�뾻ND�,K�׽v��bX�'��}v��bX�*�'���]�"X�%��~���\�Mfe�R̹���Kı;�{�iȖ%�a��߿���%�b{�_���r%�bX�w]��r%�bX��T �M� D�(4��4vOL�\��R�dɆ��������v�u������V��=r���C��?�_s�lv������̢9=�Up�^-�i��Ý�t�+�'����Ӊ��Z�U픴]Bp���`{�N[����WE�{M��P<h�Mvܑ�U�R�4.�8���%Q�Ԕf痋x����^�s�	)��x��g��urB��I&MK۲��-�:�ۊ��.q7����w7{��M؇��ƺ7g�w3��׋�p���]���c�-�ק�U����d�x�ߞ��x�����d�K��j�?�X�%��k��iȖ%�bw����r%�bX�w]��r%�bX�����Kı<~��		uIMXfRk5v��bX�'}��]�!�ș���{��9ı,Ok���9ı,O����9�,K����/-��%ՙ35����Kı>���Kı;�{�iȖ%�b}�w�iȖ%��L����O��Kı=�x�̺ӣ0�,�k.�v��bX)bw�ߦӑ,K����ӑ,K�ｹ��K���dO�߿�ӑ,K����O�Z�R[�&Bh�֦ӑ,K����ӑ,K�ｹ��Kı>���Kı;�o�iȖ%�bt���_j�fa��5a��x^���Ȗֺۢëg���vܞ���bٕ�竣'}�G7�P1�������ow}��]�"X�%��u�]�"X�%��{~�G�,K��;�fӑ,K���k�=L��Ԛ�2���r%�bX�w]��r"�!��|��9����M�"X�%��｛ND�,K���ӐFı,O��=4f��2�f\��r%�bX�����Kı>��ٴ�Kı;�nz�9ı,O����9ı,O���g�˄ɚ�%����K���}�ND�,K���ӑ,K����ӑ,K�ｿM�"X�%�����HK���C2�Y���Kı;�nz�9ı,?�c�����}ı,Oo�m9ı,O����9ı,{�����{w~u�-Pm�C�9ή�����{Gn�/Z�����{������̘�0'b&L�jj�9ı,O���m9ı,N����r%�bX�w]��r%�bX���=v��bX�'{��fk4�]a5��M�"X�%��{~�NA,K��;�fӑ,K�ｹ��Kı>�w��Bı,O��i�Y���4L�љ�M�"X�%��w�ͧ"X�%��{s�iȖ=t
1 )!<�]�Ȟ���6��bX�'�����Kı<g��[�hѪf�����ͧ"X�"{�����9ı,O����ӑ,K�ｿM�"X��L��^��m9ı,O��_�Y��e�։��)��ND�,K��~�ND�,KｿM�"X�%��w�ͧ"X�%��xߦӑ,K��=I�/j�+�\�:�A��͗^.8�a�.x�U�b9�`�Yy�����N��z�V�'"X�%��k޻ND�,K��}�ND�,K��M�"X�%��{�M�"X�%���|L�Yp�f��s5v��bX�'���6���@"dK�����ӑ,K���o�m9ı,N�^��r%�bX�?{~���)Md3)��ͧ"X�%��{s�iȖ%�b}���iȖ?�EL��=�����Kı?g���ND�,K��{2^[-�K�2fkSWiȖ%�b}���iȖ%�bw���ӑ,K��;�fӑ,Kz1�Ah�$ �����@剜��˴�Kı>�{5�Ӣ�,�k5��ND�,K�׽v��bX��?k��ͧ�,K�������r%�bX�w���r%�bX�������a�]K5�5�C��D�v��k
�9��k��s,�˚�$�t�B��2MY��]�"X�%��w�ͧ"X�%��{s�iȖ%�b}���h�bX�'}�z�9ı,O����4j��&�Mf�ӑ,K�ｹ��ı,O���m9ı,N�^��r%�bX�w]��r'�S"X��W�q�&�U"�I;��q3��LO����ӑ,K���]�"X��b}�w�iȖ%�bw����Kı<{�u��jfd�j���M�"X�,����]�"X�%������r%�bX���=v��bX6'���6��bX�'�~��L�Ys%3V���]�"X�%��u�]�"X�%��kǮӑ,K���ߦӑ,K���]�"X�%��j�CP�Ĉ �A
� sH�����'�ؑ"�BmZ@d҄��]>a	���\��5�߶=:BE�ȸ�2�:�D~SHH��E�� %JTp޶�K�N���+�N"m"@�"ET�`HE	6*���(��"�Fr��H EVVD� ������(�E�_�0dS|��	 A )-Dʤ�2�ȝꌐcCp�)���GR/��!wb��/1Ȅ �_�1 ��F	��*h�"E`H����an�ݾ�~�c���X
U��H8Ѷ��  -�m�`8���U�Z�wlY�v�8��TJ�#V�M[�m=�	��R�y�N�N�g��q�9�'�պp��l$Y.��-of��nڹ�B�M�u�Y�]��ʳc�0�lY�ġԼ��LW&�6p=ed;Y���s�%ΰe�]����֙�I�Rmn类�	ɥqC��^6�R�dztT��g��V7/R).�g.֘#6��Y�x�^`�&06�N�4+2�E ʰk���e��p0�_Y�s��v�֞۠�b�@�n����>����{v�&��4kr½;fļ�8��]�m�h�ڜ�>����oDl�`�q����u��8�ۣ�9����x���ح�3<��n�W��kF��\Zyn4˵.m4.���]>==v�uMby�'2�Ë��`FZxg��6"շ��[���m+D'+��[(
�r�-�]�<mm.�b�����r1pd�OF��ymkdaT�p��6G6�Z���fwi#	�IFW�'kY�����v`
�%:�f^�7hv�׶3l�N�u]\Z���ه�7��	��%�t�:��N�a���W\J�b]�<2�V5�4���Ӷ퍶;c������в6sE[R��%�JᲑ��n������d�ȭ�cW;V�ډו��`A����P�l��UO.����9S`'mp�'i��+R�!<�s�G`�i.��:���]�'��k6��m	۪�K��u�\�=d��٣[��1�6�s6�Btdk��驅��B�h@�I�Ny��yEuQF�U܋�%{f!���qlN[DƺZ��=��ɰ�d�[9�V�=��O�+Ź��ֺW���L͆�C���s��bM�dtm�@��{P횎�B姅�W�u���nr���p9��`ke (�E�.9�T�Y�oY��)�ֵڷ8��ݎ�\�x��`�9۠�aިI�l�
�+�j����v�]�Թ�/6�!����>Q�M'X*�@ mң�~��^*����B~.q
��!
��vۗV��{9�8+��Ht���\���&#3V�v�j��cY��si�ma�,�vݎ9����{��P\��.;e�'��lX�˯m�V��=�3e(�Y�����s�=9�u��4�;,x� ֩�)�-���v���W���A�x�Q�������ɝo.��$�7Wun�!WUn֜w]p��j̼�A��q�xyxy�)ۮ��zQ�=[����+{]��`��ֵ���۶�\qd�N�����7���'�����Kı>�w��Kı;�{�a���ı?{^��ND�,K�g��Yyl�+.�ə�M]�"X�%��{�M�"X�%��k޻ND�,K�뾻ND�,K�׏]�"3"dK�׏�ֳN����	��jm9ı,Ok���9ı,O����9ı,N�^=v��bX�'���6��bX�'�k����4L���WiȖ%�b}���i�G"dK���?�ӑ,K���o�m9ı,N�^�ڿL�g8�N�TR�Q)B�QiȖ%�bw����Kı>�w��Kı;�{�iȖ%�b}���iȖ%�b ww�����I��h*�]z���Y�ڨtz#do@�k'`�s�lXb;rq�;�����Wk9^�׻�����d��o�m9ı,N�^��r%�bX�w�����ı=�����9�&q3���v׊� ԧ	%���bX�'}�z�9�?�X�+B5��~J����ND�9���iȖ%�b}�x��r%�bX�w���~8��|P�gb�z��jStܕv��bX�'�{�iȖ%�bw����Kı>�w��Kı;�{�iȖ%�b{���HMd����Z�ND�,�H���?�ӑ,K���o�m9ı,N�^��r%�`؟w���r%�bX��w�-�ܬ��&fh��r%�bX�w���r%�bX`!�߽v�D�,K��~�ND�,K�׏]�"X�%���$���׵�uv���*]'Y�]��|Ľv{U�f���#�\���N�˷Fpg�U^�ta>�~N&q7�7]��ei`fLX���0�2��;�W�9&<C�0����<�ߒ7f�vٕ���3���Ռ��R(�T\�7f �4� �u�
P4H��"�D	R�
��ѕ�����0�Y.5#x0�1��hwJh�V��t��k�V�r��1��8�$��̙���ٗ��7f�v����?/����)�&�
	�Mu!v[��S��y��n[����ռ��s�׳�=�<.9��Z�Қ��Z�ҟg�>���7�Z EA�Q�H��2b�{ě>̭,ٺ���a~I&���#v1��:d$���fV�d�vo��'wkŁ�O/;��Y*�r�GQG¥U�{����+K2b�a8�}L@���s���"w�������W�'&,c�0����<��+v9�=�l��� ��!j�D�Oȩ/m=Z�K�S�����nw7��>*������sɘfR�&C�.Z�h�*�HR�8:��=���`~�k2f;�{XX�Z�U7uH��E�UR��=�l��Q�IrCޞ���wkŁ�ښ�Y��2��"�JtI(�3&c�?w�����I����Z�ߖ������cy�� �u� �����8%
""_�oƁ�}>00�!F������X��=��pnـ{�ـTG�HQq�?:T�`.�5l̖u�fG5�ʎa�NUUNt�F�M�m���;p�uz������:�Y[�1�AwMB�\f�Z�c2�s5p,9���`�tpt�V8`����+��ln���n��v���-��;�L���b��
; �%�/ [���D��p��s��gl��#��uӱ#��yGNJ�q&y��C�s��� +KOi�y�^���:��7T�Eіf��
n�^S9�k2��[sX�x���Ɯ�]�#\����팇>֒2�ѻ(�b�JI�d�8����̬,��a�=�s��_@��O; �z�*�r�7Dh�*��������$��ei`w6���gq߸����ݘ����Z+����5���7�Ӝ6"gz�`sv����*���%Qa򈈉޺��>�>4�S@��)�^��ETRR(��S�>������If������@��uh�ՌrF�c����K���{;�j��sT����moiŧt;�M�'x�!n[)�y��>�T��$��\��f׋�?"z1̔�[�njnIϻ���D>)�U�j�S����s+�<������n����o�y�}��ț�e4}����T�	5�PI�H��y{�)���X��Ł��,�*c�x]�H�����!�[e4������ݩ������k� �el��]n���{GT��M#��>-�I�;=�s�h�\m�Up��ۛV�m���i`}ܩ������?0����������HR�5Q`}ܩ��������ig�&�v����;ݭ/�9ė�R�+�%"��L"O�Z����:�V�~��Qj�
E�Q���`�m�.sqC�"�*)�(���<��v{����q���v��>}8�cREC��N���,.s7U���kK�2��ߐ,�e��~L"�q���KC�~(�{*�n�Z��wc.TǺ,�rt��n�bx�3R0uG�3uV��ea`w&c�K��Ɓ��%�k��!�{�_���.q6f��`w�ZX�U��8��$��UJ���UU�{����)�u�)�yzS@����1Jmʪv��)���X�U���;]����	~P�gu���I������H�R
j�Q`w1V���������Oy������:����mҺd�G-�]�-x�C�S{Yɒ�6�3�W�ЬN8#���rm]�pso�߯��a`w&c�;�k��8�0��ZX�]<g���6�m�@��Z{ҚfQ�����/�q/s���C�?"z1��T:nJv�׋��c���nV�l�v}�� u��ԌQa����5�nV�rf;s�\y��z�T�ڱ	���I�H��<�)�j�<�\\�_��ro����<v.y/�ZRN�%���,��Y��l�e�ۑ2�@jG[U����8�ӭk�b��2��)�h�m7;tƫ&Nv�#��ݵ���8޹�Bnۡ�؁�:	�s�^��e�Sћ�����9�v4�S��Ǜj�P�bGK*e֗�ۄ�+��u��Óu;ǆ}����lA�i��r�0�9�&Ƨ��C�Pl�ن�����ͺ��b�{�������A֏��FϴBS&��K�E�=Gl��Y�΀Β:�k��\����&�N���N)�E�ݚ�]����p�r��DDB��Y�w̧�qb�F8�rE�w��w��ͧ���r��;�1߹��q6j}�jR�B�5N��36���v��=�ĳku�;����t�Q9MFH�"t�[>ܭ,ٺ�����ˉs�3m�1i�(k��REEJ0t���l�;�˜ϭ��,w�����.�ڸћ���wi�8�#��1�)�w`����no�w{�ov~��YD���/Y�wX��<�)�uv��e0G�<B��)��V��~jҊZ�b�
���$D0Xq*'�U/���],ٺ������l�q�������:�t��+K�3�\I7���[�_- ���9�F(��9!�s�� ��f��\�~���"����`��ʉ�%F�钪��߻XX\�8���z���i`w&c�:��yN��v��V:s�[���#������s;<�`���$�@���ww��v����:�h�9�o�|�/Jh]�@�z�h�%Ǎ�,���5���M�����u���^���O]��M�C\�"���*����0�x��I�N"m����QЁ� b�����Vn4��a��,��#V�c�`q?_:T
�\C6F0�P��!�Bҩ���Ȇ&<�>L ̫J��w���^k��،���7�"A�@"@ W�&�8�Ja#�F!�7��I"k�ɩ�閖1P�p1�T�M�d6���*=+/�8�D�l
�ʪ�
�A_�(�E`?
��sC�У�:艈��:����ݳ ���S)8�R��IJ�y�s�s}�=�O���zS@�۹�_l� (�F�X��3���`{��\�}��|������寶߿��.7��@=e�M��Vm�-��4�߶�N�u|�l����9|�iB��� c�/*����n|���`�x�$��>��@:����?(�XG$4��W���ϳ6Ձ��z���a~\I��*>�,��`�Nf��~��/�X��0�������ڵSe�.Jr���q'��z������fZ�Ir�}�nS������ܓ�Iq�pǋ$�&�ME�y�S@�׋ �� ����P݇�!U���ұu����I�]����d\�E<�;�q���(�{������|��Z�������X�<X���`�l�6c��S)MQ4Y6]U�{�,�DDB�7�^�������e��M��v�����R6ܥ`}��e���XY�.s�&��������{�%*�M���I�����fޖ�ݵ`}���K��w-鹿{���+���Ɗ�TXd�v������~���l�<�	B~�}Ǔ�UD0ɊLRș��B�{&-���mے��vG:v��sy���r�t�f�;]��ڽ�6�6�r:�����Ge�8�^^b�y�����9ε�8�J,8-U�l�Sfm��s*��ڴ�dǥ�=�x��c`�\lP�70��;�m�����a��g�Ʒ�pL��#�6����Yգf�I�1�z�m�>�=r�zí��Ew�����ug�=\��6�u���W��r��
�:#l�G���L��U����{����q�d�EJz�kK�Ǚ,�����û7V��.��/�dơ1p�=�z���g�Y?{=�'��^��Ȋ�f��(��D�R)�8ꥁ���`}�1��m���{��_��Cdmӎ:(�Qa�s��8���;��j�����z�h��.���lL������,�Q
;�������5�s�Z��3x'���ch�0c�OJY�[N����>��s�>rmF�p��Q�]���x��M��=�z�e4k�g�u�mX�7Z�8���*G*Xw+��ɑ ��-u��ާ�g��~�nh��ZmN�$�q1���� ���x��(Q<�~���O��}pNLx��(�Ru���d�>̬,5s�O���V��V��&5	�B	�������������nh��h�W�D�LJH~N6�AG\u�۵]��Y@�.�N��Yy��kǷ �SO�dԏ@��M�m��;��^K����5�-6�5��8�����=���;�ŀ{J�8�l�\�g_0�H�������`fnڰ=�s��������x���@�N����JV���<�`wv��?}�j��'���Xwu����tۃ�J�ٕ���ww��f����%��q.b� f�~肪��Js�v�ʘ���!��]Rh8J�V�.�/w��}���$��&<q�@�����w[��y�]^�k���\N<xڍ��LR���ܵ{�ϻl�7fk�?}�j�ēg��ռ�T�����J�����2w��o��ڰ7smX}�X�*�D�2&�z���<�S@���^��`Fh���%�,&�5�U��%�]�1�Ƿ,];B���TT����+������܏6X���.quf�k���DQԡ��c��(Y�;�Ay.�籛��qf�G��G>�r���A-F���͵`}����̝ǩ/.}��x��}HR��R1�J����%��;����XX��W�����O�?5�i��;��;��{s@��qUv7#�G#Ǎ4��<�a`~��V�'q�o̬�`cŬ���j7�Q4�4-���>�@�|� �v�b"�%���jd�qQ��S��t/4���(nW��j�`}�P\Z%/O,��h�rHZ3���R���3��s����0����D��m͋nz�v��'�ku�L#�]�����zs�psH ��8k�i��&͎�un̍�����nN"<��DKʅ��������;q��yM��������eh����� �ծ�Y��&�ڍk5t����Bz"r�w���=�������ϻQs�����{s�t���;D�4�jwn6|�va��<g~vnI�o�2cP��#M̠{G~Zs�-��<��hܥǉ��d�hC�hϪ�<�S@�۹�{���^IHui�(��%2)N�uN��^,ٙj�.7�&k�3&k�>k��	�N(�C�r�K�I)�{�+4�����h[)�^�1b�ō����{����h[)�ym��.vT*ŲF�PF����cO�֞\iM�.��]vb�j����K��n��w��v/�e7�hL�n/ �ߖ�岚����U��[�I27<Hn=�e3a)�_(IV�n,YO��:{�`�(G#om�h[w4x��g�Ǚ���v��?'���R�����7�j� �w�~���y��X�+�fZ�33�qGNQU�QWs�t�:�?(��D(���ߍ���Xt��`{�o\N��!Q'\�cs��)�`���):�p�9b ��X�'�iv؆��M$���~��O��n����9wW�z���hOd�X�2��qq$���&���},-��<����)�,m4������?_߻��|�A�i%A��!�B�){)�a�੡?"Jp�G/ТQ>��s�� ��R��h�F�����9wW�yl���s@�IM ���dr�Q�ć*X�XX��\�\I..���|���4]���s��&��6�G[�HwmU�M'!l����H�q��d�^8Ί��8
F�4ې�o]��%4��&���Ŀ0�����=�j��!Ӯ:*9)X�+��R�6X�ZX�2��8�;���⎜�"!(�1�l�32���\��n�sJ�����<ySQA6B1��l���o ����PD$$��J`I2D4�
�Mw��rO��}�g���A1'�n�z��.��̬,�}��k�\qS�$���|�9��K���7GG���{�N<^-�.k��<艩���+Kw%���������7smX�:z!��TcP�EQ`%�sg�7v��3;�����s�����j:䪩Q�T�7v��2���/RS@��z��BH�"F��9%Qa��q���V敥��;��W������Ł���N��Ht뎊��̶`_:�v��x����?�C��??=��y��s F���>��Il-e���SJC!�*}ϐБ1�Ii�#!𸹎hТ�F(4��Z@	����t�'5�&�t�����0� }ut���DڃCD�p�x�5�-֤����� d r������~�ѵP�Yyj��m&��#���-���v��k�Ǣ�s�4�K�0Z�WjT-���,�%��ȷb3� s���UA㓠��r����d�aѡ��{Ts�&k�;i�W=v��؏G[n��4v�il�Jwj���R薻��rQ=�L��pf�F$@��%d�@�M@V��j�[ۗ*$�����g��"�lF���x�;�bE��^[v��j��2���L��������v��i�3��.�˲vx�jL`4��j��5�,QlS���[O #v��*c�Ppu���m��Iu��,�u��7v�lkg���Z-�V+�'�-�q �#�H��f�q�Bq��<��.�� �땃%q�V�:���q����,�2煶s�}7��r�8�&#�N�׷U��or%Wt�����0V�M�!�v�a��V0��]��kk�c��#�ݶ�]��:�FY��v �<���<���a�v��%���	 N�{u��n�T��c�O0\�.[�g�Ӳ�*�������f�:���P�l��"*��2��u����n��T��������Ƀ�.����t&�j��;F�j�S�2m&ر��� �r�	�Muup@J��+	E$s�ج�/-mUT�@\������)�M�U� ��kjU@���TU.˄�zbL�,�7m��GL�KR��J�V�l��8ۡ��8�9�lܛC�,qu�����H�fK��l�5p-J�NqT�i�]!��<��jUU���"Q*��9xN5�
��)W�.�h��ֶ��2���V��*<�(iw ��mV�6Gpt���t	��H���N���3S��Fdڸѧ)�25� -�J����iᆦ	v4W�Fss۲�I�)�Ӧ{�v1�,����6F.�g'XHm��7�%����v��Cl���ڹ�*�9�'$���Y;3GJ��Æ�M��b�s��9�eԹ��x �S��O�>@{�ȉ�u�b��+�*�bDO� ��WBb*����{�3�ch�����'!2G=z�-9zV�9c����f��c^]q��ug�']uf�dm��9{Pm��ǩޛu\c�����/3�.���q�Z��4�X����9�6S�#,�ԏ�n��4���4�˘2�Q���d�f�P��=MZA����c�i��m�$������AF��9�{I@�p.�[m͛n]�ԫ�m����q;XX�F�����||u�:t����S�st����M�Ɨ#�3�݅Sz�֜qgZ���C��]R(�0�n�����(_�!}��X��E�t�TU�X�1���Vw
��ǝ�{ēg�t[=M��(prS�7smX�+����V���܆	F#�C������ǹ��`k��`fL�`�Ĕ���X�:z!��NP�EQ`c��=Ż[���������Y������˷aܖ�(��5q較��^�o3���9�v���h�a;������S��xQ�T�z{����Z�3�VK�~a����;��d�D��Q&�@�����DB򈴵:w;8������M�'��TT��q�C�����|�
�W�Z�Z�w4m��lj,x�ț�5�U��]�@����=ͷ��έ*@�*:#�����d�v{��%����ܧ��ǝ�`}�w,��b�	0m����'�q�"i�NF`r�F�yL��7��Τx�����|�p�8��9)����`gr�;w%�k�h�]�`�`�<1�&�h��h^�@��Z�w7�h�����NP�UE��se�������& ���$�8`~�b��E�DR�&�R"� 4��ZH�P�O��;f p�p�*T���*Xw����97n�����̬,5q/)���X���R��2F�DҐ�-빠[e4
�W�[e4܈�A��`�$K11���6(5��:�����y^�d-�+.H^���u=&�� ���}���*�^�m���?0�͵`n�QHG�G�U:��E��;����wkKw6Ձ��������Q���PI�H9���O�޻�{���owkK^���_ G����Ĝ4z�h�M�mze���"�V�)��o;LD������M��-��W��-���w4��pq��@آ�o8m�u,����ݿ׭�ݶ��ަ�����^�[�-�XKv�;�UQ�{�,̬,���~a����W���(�r%�&!��l��ײՁ����ם��s��Hfz��*��:q����o�X�����%�.,J���@��Ɓ�X(Fjc"��J�x�v��1�l�3&c�ԗ�7��iQH�r&�^w%��Ēݭ����VfV��sP��_�B\��a��P4(u�F�*6�q��浣��hМ��v[�����0���?�|h�} ^�qmkX7<%�MƝ������5��l]յ���\�M�q�:uv���y�C/9�X���tʏ�u��g���u�qɋ�ꎩ�`�p(�.L�[E1e�eq�$�����"dx�\K�����Y��;[=nwz�5in.�r^���:�Ny�.��`����OgQ�-{���w�|���ʹb�NXl����Sq�]��{ȹ;.���r�\:x�K�(D�PHqH9�}_-�]��0�������-���r89)hz�h�M���]�@��2�$�#�Bnf�z�h^�Ah�&�7smX�FV48�)�����1�r_�lܛ���͵a繷��W��_8�1ƣ�!���ՠ[ܵ`gr��1�rX���w�-t2���GN�ݏo5��a�axK��*ht�n�ծ�s,���]�#�Q�s&�$��m�������V<�Os�ɺ�����S����)��`gr��K�|Iu%X�T��9ڴz�h�65V6
U9�<�K;3�^\���s@���{�Q��%c�A���ՠ[�s@�e4
�W�x���bDR������ܵ`j��ޞ�����ՠyC�Q��-�}eB��2)����[���'=ps�<��(=u�z"y1(ƈ��Л��^��W��/;V�o]���J�C_�bC%UQ`c���Iq&�ɺ���Vu��9UqW#K��o��@���x�Ő�#�$��/ʽP����t)���������:�;]�
��BT`��R�����8��o�`nm|h^�@��Z�}`�O!�"�nf�z�h^�@��Z�w47����pq���`����u�Zx�����,�Lxs�v�s�#��3�������|�����0N�����ՠ[�s@�e4�(�A\J	5	#�/;��o8�9��Ҡ76����q$��~�pO�&&��?��4�S@����hz�2�Ǌ<14I)XjK�\�S���,<�K;3�����)��޷��'�K5�K����rHh{����@����3�XX����X�P?5'�u��IGk���N��f�]�&H�d�kl�h�m:.���{3?fȷ�����	��������w-Xܬ<����,���*TH�iA(��/�w4�S@�ޯ@���~\I&ϵv�T�i�QN�%+����*���/;V�}빠[�x��X��Ȕ�U�W�^v��ܵa���OsoK�Z:�6St7	#�/;V�}빠^��^�z���\Ŕ	��n0R��c��m���je�^ȩI��㊶y��s3K��"㫒6C��8��t �onr$�����{ǋ��/\��{r�ر֝˫t�KC��lic�7[�p�f�l�-�N��n��<gp�m��%�w=;3l�6m���m��7o�<���yq���Mq'Wl+G]wH��y�b:k�֥��ڼ�x汄$�M��!�ջ���u���\��&���.2Ms<�=Q	w��xss����jc����y����B�%?�n�Z�3�XX�<��s�ɺ����@:cN���`gr��1�2X٘��e���K����Q|`�_�bC�����/;V���./s�\���Z�=����y%(��<1��@��Z�w4�S@��z{bN�	#i�	G�{�j��I{�$�����<�ޖvf; �ӕĂ<O0$d�r<M�r�l5� d�n6o<l����	x�:;+p�8�E�s4��hu�@��Z�w4x�ƪư����WZ���i�<�1�QP6��=�=��C�͵`gr��.q$٘h�'���QN���u���Vj�{�ZX�}w$�N�Jt˅̚�%��ܞ�T��{�`{ޯd�vd�v��,
$��Ĝ��)�{zS@��;�fZ�<��b�֟� ��1N,��^y���1�\s��q�q���l>ѻ��{��z���x�DĆ7$=���4]� �� |���]U��J�n��]UY�>v�w�,�`��9�Fg��D��"A$m�����=�����0��{��X�o�hHG�.�|ʟ�GR�OȖ������ /�h*� Y"Z����9�Z���#�u��$H�`	 [�nRq����;]U+@4� <٠>��!��1$!��y�w�K,K�c|%Li ,36�# ��9���X)wv�ۇ�`�Hf찰4��1�KrS��?j5��H	���|����W��W�@5����* ~��'�q���߄	��ٺ��+K�l�Dɩ���QN�uk }�����0?B��y`}H���7�r(М4=}V���,�w-X̬,qn�m�n��!S��帝qF���S
�J]n�h�x�8��N �#fx�HX��E"����@��rՁ���y�$��ܛ�`u��k����Ĝ4=빠u�����@����}�)�(�xbks4{������o�mi`}��W����r��86Aʪ,?.s��ܽ,�֗$�߻�ry�W��?�q���6���_�D�<qE�<�8h�����s�������`~����w�������گvޓ�^�I�ۣn��`��&�{c�F%�頺�ڥP�o�߯����`�ـ{zـo;f �+���U���I�J���X^�&ϻ��������w7�>����X����p�7��`�ـ{y��5�f �ɸ�YACN:�U(���fޖ�͵`{l��篪�<^���eƞ'�$�U���,�$�|�Ϗ�O��;f䟸�W��J��cD�Րcf�3B����2ٙ:䅹\˚��g��yx�<���Ja�6��]�l�I�|3˅��8
y��J�4��a"� ሻ6Ⓝ��9݂��O�m�%���Q�[ZB�������eQ=��-���v�\��X����7v����%� ��j"f�F���.�c��E���)�-�r��D�X�g���O��"^F�9��ڸ�1v�^ �B�8W:99F撞y�uG�t@O&(]��+�}%5��TO<����G�ڮ��9�GM��:�I�@�L�]� Jn�� �lu�i�K@�z�`��8�l����,�Md�/蘐�䆁�)�{l���w4�w4
����5�Q`�8�zݳ ��ŇС%2��b�7��`��dq�F�D1)�z�h��h{Қ��h���cY1d"�Uـw7� �Ds�><}��`�٠{�G�Ʋ3#�BLrH#�����í�gi�8��C�A�����\�<�û8E�4z�h�)�{�S�f�b_@y�j��ME"�
q�:�E����f��?QkC�Ӱ~q(P�DB�	U��_��?�`���/O�<Yq���	��4z�hٖ���o�7]�����ϲ�EE�!HەE��s���w��X����h���=����M/�1!����h�)�u��u��-�Ax���l;���΄8�mڽ�Yܽ��N��
�筞���v�Ó]����������9�#�)����S�p}l�;]��IB���-����cq����@�Յ��\�fwkK6f���{�Ĕ�|�����5��Mʢ���x�;��n�ED�� � � �򈫇8��XOI����ex�3��di�1ȓp�:��@���@�Қ{e4)E7�&��8�k��Is7/O�gv��;���$�}�;=������ٮ,���i��4�*�r��t������GkR&浽r<.���^~��@�l����Z��Z�e,����B��*��ea{�%���;=7���v��&ϳt��N7�lHc�C@�;��:��@�Қ^��<]�RH�`�k�ԋC����?{��o�|���Ł��aak�G8�,���(F	"5��D�OAEٿ�D��3~�ܓ��WT�T�ETm���`w2��=ś���_��-����#fI�iY9<ެ�XH��2.�V1����9�$���ib��Q�����EAT9T~7+K��h_U�u��{�x�5V"LI�@��Z��Z[)�w�S@��Y`AbjI�@�����eag�9�s˒o��X��;���O\k'�'�ȴ�S@�Қd�v\y����ih�N(�B��TX�������׹���eaa6��� d0 �[{�MI�/N�c�y�hSv��U����#��=�3�ݞ�-�ё\�YC�X(*���ī�cd6�n�؎z7�F5�7fI�ƞ�s����"p�h\�X����?���Ƅ���-[�E����]�m+-�V7K�Ջ��gsm��S<P�2�v�W��	�6P\���[����X���y2m�k�h�mnH֚љ�=6��|�)%�dٚ�5)�jm��9�֘}�8�ls���S�ﻱ�c\<�a�	�)�K3�H�T�n���?�7���ٹ���Zj���w+K癣���@uQ��S�1�r^���Cw޵`{�^,�f;�H^خ9$Ő���R=���ޔ�=�ՠUz�ˀ��J����ޔ�=�ՠUz�	�<�ߕ���.���""U7�,�eZW��;���-�M�e*��̉)ѥ8ѝ��חD��D�H챔��t��q�;�K8�:x�Q�+���p�Cm��;���s-X��5/�;�u�<9�B5eS�T�;��W��K�.%×fͯ�>���ǝ�~l��KD*�RМlr�������&c��M���`[�ۚ��ՙG��m��ػk5��6X�2Շ��no�,y�9"S)��5"�*�@�m��/�XXd�;Wك,�TӄB���`�=��ހ��#��qՈ�ɨݐ�]̳p<��y%N[�*UETM2�J�����>����'q�_�c�:�lՄݡ���@���[f@<��-�}^��fZ�%�����8�B!*���w;�'ow7?�,A��P �@�
�H���D�DI��hO������?}�znR��,�k&��H�*���2Ձ�eaa�q{�s�={�`u��H?M4�J&�z{n�}����Z]����Tm�-�5�Z���є�����0V��z����W>NF��=��t?�"4��h�)�{_U�U�^��۹�yz�Y��FFГ����s�\\R{���j�ϲ��&�V�)!���'�����w��h�)�{_U�{��@#ĈJuR���\I�w+{����N㰮1�H��O��l6 �9��s�7$��3�ڎB*
�r���ea`}��hwW�w��h�dU,Y��):�f�̈́�źx������1Zݺ{SX�;���*_2(�1<0x9bN��Zw%�߳-o��{����iRA�� ��)�W�^��۹�޳@���@�z~���M4�J'z{�j�3��Y�q.7ݙ�����`}�R�1� HNf�^�4k�
���[w4-�Vdo��$��&�������[w4޳@�����9�$�a��_�I�R�;	Q!�,jв%-eD~Ї8��`/Ut*_���F)�s]ː�b����N��"G�&�:� ���Y�!�b1��]'�WXJk��f��4�_��5��������׫ L��ç�~~H�t	�]>@�E�(���B��*��{�����O{�I�t}�?��hd�m�AKi�im[xlth l�Z��3]��&�Gf�Jl@ +��KԬg1�s��;k!�E���E�y�3��i�35t<&6:�#�l�u^e�,�G+oU�ͳ�Eny�,i���f����۴n�M���P�lP<V���mz��`ܨ��[�v
l���J)�v[�����jL�7:�:M���^����˔l�V4?8�Kv"�巋#GV�P�O���v�!Q�6�[����W
[��mq��q��R�C��B�N�pn��[�ԯ]p� �ltE�a�x���VWU�1���.f֚��خo"�抶-��#rv�,g��Nٞ��
��6X*��͐��6ݭѷYnW�W��K����w$;OV�\�Ĕhβ[�.i��1�1�x��0�¶��ɭ6ݹ�(�
�&�+�����[�yp��r�%����ʵ��$�Enٗj��Q��p�X��vw;m��9d�s�N�)����6�T��u*��{u�>��^A���y�d��O��W[g�����
��:�s(��y'�������s��3�� j���0ob�,�UUOX�LS1���-�47<U^hԛ�Z�r�*�:B��c��X�#� �Xw.���%[]AY�yڮ��RJ�o0[@�l���l�5�'l����s�5�D
�pKT���8[d�oH-g&���WUAW��a�U��<�Ga\��l���@�mD;v�0^�m����3E<��m���mt�[FK@MJ�K�Z�]��[R�&��6%x٪UU��{)�R��1�L��3�1��ȨT�kG[�nɞ3��2kOH�](�g��h��s�^2�nw[��������d|��ڸۨUr�dj6�H ^�W(��O5<Ɂ4�YǴa�]0m�5����X6%�J��v^4���f��:^ NN�X�'q9ӎL����&��÷E��>~~�^�h���f�	���XSZ�$�賉'�SSF�n�in��D�)�P����v)�TD�=�PR&�n�
�Q���4�@!�8���D�=ڈ4�F�-��ƶ/nSvXl�O2�z��A(��zzۢ��P�QEj����qkQ�dK�W�mb�:�N9�Q�9��o���~x��8y�����;��u��l��n1��p��n�۪��L$���!]t��w��k���E�ˣ��D��ۛ݉�T#S�u�v84:ySg9�qΎ� ���zex)�iC���s��Q.�3�,Թ�j�̒����q��@~7�%�����7W:�:���c��qc7�F���N���#k�ߞ��6}��bi^&�_�z����[w4޳@�}V��ج#�H�##�G�ym��-�a`w���yܗ�����=����R�7)X�׋���g�K�M���`}�����t�R�N�n��,�w��;������<�{�zXS�6şF�	�I�@��z�g���~w+M\���2f��fS�:�g����s���d捊�Ws�/-�.��m$[���Y�F6���j
H�-���ـwW9��:�5�b;�kSE%�K�7$���f�_�n�USަ���ܓ��}��s����
�����1(~ �I���~Z]��[w4��*�H�$98�uN�x��͖ۻj�ϲ��;�ڴ}�X)���E�@�۹�[Қ[)�Uz��9eĿ-n3<>�`�2�y�׋Ү��tdX:����m�C�1K&<C��%�4�r~#Ĝ�ޔ�;�XX�7���7+Kw4�N)Q�U7Cr������$ٯ3e��gƁ}���$}��m�>� ��GE��3e���agϊ5��B�Ĺ�{�M4�����ب4�MB6�z^��-�M�Jh^�@��s�D��D�,���K���z~^������ŋ�0���I,3�k�"��q��S�����NC��<Y��yqf(�1!�I�Jh^�@�Қ�)�Um�2A�9DC��w%�l����������4��`�`"G�r=ޔ�-�M�v����=�,����㨜�,7����w/Kwe�v��srlD=�

�"���V ?�S�*�8�߽�X�|]'�Ӂ*��r�������ޔ�-�M祉��km�֭�F���#5�ڞk�Uz7nm�qk��v�ͧ�6g=L�W��=�)�[Қ��4)��Pi���mH�oJo�$}��{女U��+�a�udcłi��3;XXs�Voo^��7+M����Q��Hc�C@:��W��:���oJh[T��fA��IɠUz��Jh���u�6I�C���!����m�f���ܤ���~/��Δ��"'�힪p��p=0V͹5ؒ�K2mH�6�n�'Ka)ӯNC��1n�q-Od��MeX�l����s��nv�t�ĉ���;�N玞�P�'1����t�n.�M{۴�s��%j�h��B����\q��q�r��P8���x�B��m��ʁ���H:�t� J�C���[�Ŵ�=-���t����������gܙ���4i�Ћ�Փ���ճ�OJË;5�ڌ9��9`r^9Ι�q��ĔQ���ߧ�[Җ��S��V�w%��\I�
�i���'�'!�}��׬�*�^�ץ7䏾�1<q�L�@N~�M���zS@��Z�������1�RM���zS@��V�y��`|��9�Gq�R:��u�M��h^�@��z��n;���s��z�.���Z8�v~�^�����u�^ڗ�3��CF�^��u�l1˞;	٬�|�� 9�η[�n��<۬���"�T�E]ݘϝ娆��P�.]���XnV�w����3T)���1?�94
���zSO�������;��H�D�bJ)$z>�`��p�;�=:�`EMر���O�<NC@�{��~W���W}��:���媭Mdx9�c�]�{=^�Z�hz۞�v�F�l����FHwTI��b`���z׬�<^���)���r���>��G��I�8ǑI4���Jh�z� ��h�Jbx��i�F�@�Қ������}D3�s|�ƈ�^�.���,��{[�v���ܓ�y����k!�z����Y�~fKy�zXn춓��Q��tۏ@:����^�ץ4W�^��w�b���r��OF�M❻W�3�\y9���tum����͇$l'jb�Gvz���rh/mz^��=^�z׬�/tV�f$��G�u�M�#�]���V��d�3�L������㨜�,���`��Y�7���3r��/u6cc�b`���zߗ����6{� ��f(jL@$A�B���� J��Q-�,!B�Iտ�33����@��7�RG����� ��u�ou� ��u�{�� �D(?��g��;Ed&�10p\���݊&�ܽ���9v��&,�M��h�Z y��ww�]nO��j���￿�4W�^�z�h/mz��ucc@&�����Z�;f��� |�,ͺ�Jn�*4ӎ��,�V��d�S{���]~z.ꢑ��H16ۆ���2X��V����8�6��72��`bp�������=^�z�m�[�T�E�$V��Ș�}����;rn�FIek����{��N��uzsmu���vZ9��g�kv4����u.���"�+\�K�Ɲ��\nyq˅K��^��[�U�zV�r�9�rbnX�;1V�;ns��\㘱�̱ԕ=��K�h����^�ȶ�X��kf�J1�� ]ev�%�mӦ��Q�L��Y��;a7(�Z���	)�]�\۳�AE��i^��3u�7c��w���w���z���[�Ox��.hWh�.�jU�Wp��rJ9�k]��x�9��v�]��W��n;<�~q�s8W����/Yp�<^����h��1�Ʊ0p�br=���[��x���X�uR�Y�Cq�����נ^�s@�{����h��5pCI�8���8�7+������b,5?�we��L��b&4тm	��=^�z�.��d�3���
[�%�54�P� q�q��r�֪/a���vӯ���w։�nv^=��@5�c���'$,��o������w=��@<^{�@�]ն�i�9�[nh��r�������(�];T�,Q�`���X��� ��F~Jd�ؾ�H����")$z��4}}V�zˆ��^�ޘ�<m�LRs4��Z�.��z[w4z�1�dX0p�cr-���z����z���(S9�1^�a�QƇ�Cr��z%#��r��8N8��s.�=�Y�W���(�v�m�?����m��=��p��0�\)�R�#djG�^�sV$yϪ�/Yp�<]��W�`	���0M�9��\� |�p�8�;a*22TUT��:}B>L,�j.�������5�I)		5B C�`��	�ae;����: �9vq�	�?=T�OԐ�%%A������@! �~�~o���0d�`���b�# }������H��h ��{ �a�<xp�����	��_�	,��F1W�2���%Y�HH04l
0A��P"�U�� ���j�S�!P�G�A-��[$"R5XX$R P��c% U	�)���~�>6'��a��'q�6���~��. ��	��H2BXH�S�a��!��h��H|�g�HrԄZ$^�VbC�@��=O���̈́*ƌ�
0(��.���S����*��U�:�����A�*�Ȁκ~@�!�P4���ר��ߣ��������͖�u*4ӍԔ�7�����X<͖w2Ն�q�e�h��7$���X�1s��� ��,�\� �vрkAC^��nz�e��M��#�c�:(���kf�g��Y�ˎ�s��`ۖ�����ŀ{�����>��V�
� 4ӂ��I��<��h�\4Ͻ�`}���y�s�M���ҊB� HE�Z�O��;��=��hs��Q��R($��BI��y�f���_/Hk���=@�">��B�Uh�A��10$Q-h ��R�[eD�"��Шt>9���_�`n�a!��$�Ӫ�[x�us���F {��������q����;�A��8,�F3k�i��|�݊�9�l�r6�������(߀���`w�X� �����;����v]$�$Ti��)��V"���M�ٛVwvՁ����yĹ�6u�4�U!!��1��h��4m������ˆ���X��j!��7$��S�}����Ӏw;h�w;�����d��8�s49�Zu� �s�[x��D}QI���EQ*��۳�N��ky7
��V�b�5dp�C@v]vY�{]�f�rn���������إ��Wm�����I�o7���cɭ��Fɍ�Pl������BuI�<g<k��n�hÓ�{m��&L]6��866�����B����i��Yv�E�$Y:^.��Gi��7�i�q��&��e{e�=T>qۗ�͹��bUq\����75Mh֬-˯���_ |��������[\x�^Ó���$���]��n�v:��ݝ���.�Έ�9�����l�0�;��-�s@�U��x�	�#P�a�x���-�s@�_U�[e������c_!cdjG`n�ڰ;��;5q&�v��se���`4�/�6	��;��h�p�<W��-�s@�{3y��MF�Z�\4��m��;��h�vU�͋#���cIGL���u]�P��/6Vg����k]>x��<���wc��M&���z��h��l�h�+�9cpYr=�w7��OȈ`4:�?��T�77���`}�Z����=�l�D���p����h�p�<W��-�s@�x�6E�"�$ƤZ�\4��m��<��h+�cx�čr)&��[n�޾�@�+`o9�n�dh�M���8��)�{6�p7��^�<�OA�����8����#,cl��H���s@�_U�[e�@�^�@�.<���$�'3@�_U�[e�@�^�@��͹��^��`��Q��m��z�=�� V&�qqz�9��N=��Vݙ�����dPX�c���na�x�W�[n�޾�@�ˆ�{���nIS�U,��V�3�������??���9Q�\ŉO�N��M�M���yu���(ޛ�5x6ɹC6���tr6�Z�dP��y��l�h/z��w4{�\x�DcR-��V���� o�,v���= 5���~�K����@�w�=޻����@��U�{��Fƪ1�A�z|�`��8u���P��I�P�'�O��M{f䟏9�ɗ%M�9J����;�ݬZ���l�3;w4��C|0����"n,LĻ��q�YL���c����T��:��q�5�JC���u%?�n�Z����3;��=}V��z��Ab�cIL�@��:�� ��9��Ns�&Fݯ�H��K�z�_�4=}V���Ů���6Xb�0��*D�j�լ�\� m�F��u�6�,���'�$A#�@�ˆ���u�6�,�\� �(�D(JP���n �]nö�̭�jfk�z�4k�U��y���{��q�}�.��]�m�L�%�n�س���9@ ��lG1���G�k���5�k���'<��\����!hF9�v�c/��۷�t��jƈ�m�b�m��ǍL��a�FvKngiٛ�	ڱ�;gŇn�\����:p�m"<��e��Sp���/#[k�6��K�3L�&MҲ:;)�Y���Ý�ϻ�����=���� ?}��\˭f�d���[%�͛�1�SmV���von�u��n83O�ŧc8�Ǎ9!�'�@�[��m��<��Z�\4?��?Q������	q�}�ۚ���@�ˆ�����<�R�
)54��j��s�7���RM���,��V�%�N�C��&�n-�.�ޯ@����_U�v^�dPX�d�I�������o�\� m�F�B��u�|���!�K�����5�'�{^'�p˱��m\89_���٧��V�vV��j����;3+����ͫ�Sf�l�r)M�T�)X���h�B�kRC�+��*%E�E��iӆ�1?��WRk���O���h۹�w��V$a#�@m�F {y� �x�ms� �)x�H�"qI0�=�4m��=��Z�\4}����M��Gw�6�,v�� ۶� ��x�*�	�yy���Y�1	�NOX��g�uS��<e��]&�5㙶����\81�6�u?� m�F {[���`�^��aŉ�ۋ@�ˆ�y�@����_U�v^�dPX�c��Ҫ�`���o�(IjDF!BJv4n�!�o7�;˹'{�]&��ۃ��H�2bKnM�w4}}V�m� ��f���]Q"D�8�+�&�`��pݴ`���o�*�PQ5��cS�Ez��n����ɴ5��l�w[v��tfG.���miI�H�l�h��4m��=��Z��q�<��p��$�@<��͉��x���8n�0�LUEM�I�"�ɠ[n�ﯪ�ĭ�p�=�hP|~�\LI�!9��
���]�ܓ���M�'>�u�(*����BQco��YQ7IR�J.��pݴ`���o�\� ֿ����l�x�6����
��]����k�ns�[nxN�{fÒ0�܉Qc��np��0����� ��9�vрv�q�2,B�1%�7&�m���f${�5��Z� ��r�[:������j`�9��gƁm� ����ڰ;�LD���U8��=��N����`ffZ�3���	�Ŝ�J)�r�;��`=�9Ż���'����~���rO�EW��EW��DU���"�TA_�QU�DU��DU�������* �D���� �D*���@��
� �ET��*
���"�*`�B
���H*"� ���
����
�*H*��B
�H* �@��B�*�`�F
� �b�B
���H
�����X*�� �D� �@H**�X
�B
�",b*"*!  )",`�B *
�
�b**
�@����E�� ��DH
�
� *��D����
�X��E��E��F�B"�����A ** Ƞ H� �H��AA�"��uEW�* ���AZ���QU�DU��EW�A_���*������"��"����
�2��Z��((=J�����9�>�w�          �   �  �h <  >D�(J�J��QER�   T  
E� ��    R�  �`   ���  P ��`\��.m�R��,�4���o+xx :�ۋz�9��]=��rz�{���X����� ۷�������� ����r����'��M=n c��g������o�x   �� @ �(�����1<�C��ޝD��U�}���}K�z�ם�j���qgYp �һ���9n� -w���YN�>���}5��N���μ�]9r�{� =�m��w��׎�%�wK���W� |���(� ��N0��_NO��<���gJQ�#JR� g@)�`t�,��&��g`}=)���٥4�e�
R�  ��ҔR� � ��X JJ3��4� ч�:8 ��
h���Δ��i�� 
P P. ��bP=:\�(���}Ͻ�E���en-N��v��s�\Z�`� ��>G�,�n3O;t�� 
wJ�ܞ�x�^��r�;x�R��}@��VmO��t����u�����o |> �P �  ��`Ql}�J޾�־������mK��,��� �����Z�=�yܼ�{�y��ۀ��{�W7|�r��x z�7t׭��w�m�@�U�}��s���^NN����w���k��gZ���ԫ�   4�&Sm%*��db41?�M�*R�  O��)�C& LMD�*��梤   ��	Sm*R�  "�b�� Ѳ��{���p���c�s����{��{��� Uz��� "�� TU?� U�P EW�TX������)C������c\	�C���"h�O��K� "D#��>�������g�.u���d����`L ��5�d��"�2���(`�k�2�
��"�7d��0�������$�4���GL1R�:j�J40��i!CZ�P��ɢ%�$��B�H�\.t2�!G<	
d2��"��z=�u�j5����`�c����`4Sx{�
��Dh�B@6
8S/�@����B���1bFA�uI$$�9CQ���E`%H+F2)�I�CM������##���H�\Q T��A�! e�d9q1�!/I��_+�c�Mϡ&0C8	s���ۣF�>q���.2#�0� ��rk��j��-9O���H���&t`�!R�09�7!�ɦ@�eB��40,�b��ɗ�gg�E�#�2XJ�`@��h�°
&��G�ILKL���bFB�#$���w f2M��B?'�G��xl>�#q�;�-����ISZR���M��~C�H�T 4;���>�BF-H�<�d1m$�0Ƹl͡L��4�M:YK��Iֻ3]HXP��r��b�I2�PJ0��l�H��*9��%b@٤��C{��R�;�l!��"c@h64�@�@A*C)��G7�t���x�l�j!r�J��P�1X1+�p!�F�;� FK�P)�걹`�$.&l!GYL��� �3�gU1��ژ� �%p�! �@�� � ��!��� D��J��0*a@2���&uy��~vm�H! ��H�rF�fH�.��pA��4F2�@�dBHᅐ2E� T�?;&���ޟe%0dr��SLB@�@�@��&M^��a���$:0� �X�"2�c�����V
NN��fe��8`Ϋ�4��S;32d�E��&�3{�>�9�2e�B���3�!~�k�ϳ��o<�C���x���\rҫ���ԟ"HB,��Y0�U�	�@�D*�w��A0,Y�h��e���A�C���b�o�i6��9tm6l��,� Τ6}��$����kj*�ɩLjj0X�L��$�����2si�4>�G�0��a D�8�6d��
�!C	D�h$e��X`"\8a�`+���`���.H��E�����H^4`�����w!��FL2���H�X�rCR1�B�Ṧ� SC!��M�0d�k�ֈC=���~L�H '�V��F���3��C���:���i�w��A�e`F)�
`�L�+K"Ja��iNJ�!C���H1H 
2rC9#a>��*`�E�U� �;jm�
`���	fM��g��a`U�4��l�#��Y�;5�i�n&4`@>~Nɋum�%EѝgвD�Wl���tH�����2�aF0�0	
�1�[�fe�,C@cg�(��, d.M>���Ӈ�p��"�R���%�&%0�h85���BI�s#>�R2H���T���{Ϯ��d�
J93��%p�"u���C2��a@��Ja����Sa��˻�BD�B)Ld7�{X�q��ލ��u��3�6L�������Ci�Jp�LdSj�4�H��W(�)m9�4��?w�Y�\)����9���C��.1�B��LL��>���Wa�đ0.$XBG[#L�z5��6:H5�#	P��H�p1(c�p�U��ϱ�"A�E�Pљ4��u�SI���i�b, �H	HDp0
�"- > "X%D>e���}0�9�֍��!�f��5����%�����!�A*��S�P�C��j�ӻ�sf��0a�0C� ��e�����\e�mK��0B����0/� ��4��ssF��ؓI�����R T�d4�a\.@ B4��wd�:��V��òRn�a$�9$��tİ%�'�rF04��\��I�1��i(�B>���4F�o�eb@����0d��@��'2h!\g\C����� B�E��Jl�#��ˇA��k_$��0��.�:��c�ƶ��Y��Ji~�p�t(m>��r� LgP0��޵�
2i��t�j� `�v�6l�¸�ɤ�B����x��f�7�o��h�f˥41�u����:��rN0�L4FJa#]��N�*o��;#�����p�+�`Ń\82�$P�WM` SI!� @ ix���sh�$*������`�G!3��RG!�$���3�d��8�ɬ���ѳ.G&tn��b#eH\�96��357����Ψ.��;�������Ts*�9U�r������D����U������H8h�u������XSO�#���e��"P�R*Ђ�hAl0�
�F@�
�!S�f��%��uA�EH��h1�˦�~$�`�o�gg|�9Ё7�'$u@�Ŝ�8��``�ni��HH�>9���>a	�d!ge�r�,	3��˘B0a��5 �a�
��e	[��7��V��3�����C����߲��	�(������ێ��5ä�w8M0"�]�/&2Ea�o7sI�����+b@�R�6�3�5�H0HR��JB�Aε��y2���;̷8�͑��C���@�0d�eƴH�����eX7�XQ��#�HG$��ϛ����dԹ�0	�)LtC.��*a	#\!�	?\뗙�1��������r_����M)���#qs@(`YW�&G(F���m:�ό�D0�"d�@#II��dd��"E	 ��b� �L=4���yM�G.��B$�i�5c �P�C\Y��[��đ2� 	�0�1��*��� �	(hE��	#rkF������H`�,��C�ԋ\e&�ߩq3�u�wl�2cC�y�/�ִlcD"-HߌB��M}�J�5�%8�������O�l��>bP�$0��t�ft��(Je��	p˄�n���������NT;j��#�X�' �p�Md�l�Բ!2��s�H��B�`��Ѣɖg�]����0�\V������w�=]]����@�$,7
�aV$!"���,��w�Rك"�~��Ń�}�-i<�+Σ*V7��Lrbpڙ@��"���T�U�a3�L��`�2d.���`1(HCBi� U��bQ�W/� ,Z�.`����1�B�)%1��o`K�P76BKf񈆤d`�ٔ�`�I)�v2A��;M��u��#����%0����\d����!@�U4���.��)�%	t�gL��`��b��1�0eFuT�DZ������cp�#�8�0�4�8B���F�|a�:H��3��6��  p ���     m    m      	 m�       l �  �  H �             [�����     @  $   l ��m�   � �  i6�p[@A���e�  ����hi�.E�QN�k��f�@�- Oپ>  mm�   �l�J�]/ZB��g��Ӳ�y`'�Zݩ�v�T @�-�,0�p�I+m��-����Kq����[VȻ`I&���٥P ����j����K2O'F�>~ž1]�J����'h�2r�;�$pkX-�����|'J�^9lN֪j8��[Y��-�����<�DK]u��J��6ث�<k<���*��9U�����N�,���aŵ6�PlS��: lT��!�q��PʵH�b�8�.:[+Z�M�U�PS��	-TQl����0c�H飭����W&�*�U��q��������*�P[VP��-�k�#i6Ӛ-[%s�mD� m�%ҫg�yQ*����B��U�y$�H����UuUJ��.��Iэ�,C�e�/;[UU$��Xm-F �K�0}���^�ߤ  [�������q�� �k�  Hph� �!mH �����bK���8ֻ9���R���9,���9R]�-�h�l H���ٰ�j��;m� ��B����}�� ��p�1H	���TK	�UWX�*յ�"��$�7i)km&   ��  8 !M����eXU�É�����\�-�D�� 
>W�ڑx�UPmͺ� H�8�['LZ�[R�$6�˄s�� �v	k[��6Z�t� 6�jZ��� ڐ��:��j���T� ',�2`�d�$qʱ6�H� OY�v��`���� �c-7�pK(-�i3����Y/���m��>�K�d� 	"Y(�$� 8	6[�	g��pJ�erT�m@T�xZ��&/Z-���p#]�Tm��m�sl�5�7m��v���[y
69݃k��+t�UK��` [Ae�(]ԛu���]%�������p5���u�]�̎�]�"�9��YۮA6xM�웎�4�:�H��Y�]�*��9Ƣs���wLm�  � ��m�u+�i�en
�,n^k�t�4�m��@rF�Si�$��� �m� �+��Z�kV��� $m�Iz��e�[@ ������n� H  p �i6ݎ 	J������� $�8$�8f��cm�pm.Jŵ�����l�   ��v�I0��m��m� �A��`v�m&]4�-�[d -ڻ`m��8^� H�x��-�   � m��trI8h� �$ [@ 8 m�    �   [@   [��-�  ��  �c��ڶ� r�   $�   ����l� �:@�Y( 8 "ڐ  �d�  m���	6�`$��k�q�8�n �m���  $� U�hm�m�ݶ ���   �v��m��Pq��m��6�   �p   m�Z�V�ʵԠ)���   p    K��kؐm�2H9"��N�m��6�	�����ё�j�[� m�[zMo$�9E�`��WJ� �I����UR�H^kd���j�ge�r%�-Tcn�˲�zܣl�u\�-C�CMΩ�Z)�3�Y�C`ᶕjU�8������;�K& �p�-V��]@g�	V�    �p�:Ԇ�p�j�ݶ�� [��i�   ����n�6�2)!���n�m��  ��ѻk3 ��*Sm� ���� 6�"pm�$�;m� @$ ��i�h�6Ͱۭkh��^Ywa��� ��  �m�)gKasm� [D�'Yv� E8k�ͱkN$����l�-��m۶ʶ� [@n�m�bCl�$m�H$����E�H�i3l 	�X��9��-�h M�m�`-ԛ��M��ڶ;e� �   8�"��h�	�+��IB+mb�f��n�Kh �h��)ms�mm ���c�ݸm���Cr���8����8p8�k"(-����f� �z�1
�i9j��÷`�6g�IjCax`�m/�e��r�F�X,�s�6Ԯ ��o�	�\�E6 �i3v�6�$:�*S�N��kM���I�Z��Z�y��W+m��ċ%���m&�6� �Iw�-#��1a_d��u��]�&�k�غ��ꐚ[�+���AT� �ԩٹ�V��U@Rlhu��T��tJ�I�mF��*����t��d��`�ƴq���,�Uf2���C#>HX����X@��`�dM�㌡g�8�<����uUV�rշm6� i{K�F�-�m���C�I"@5V�G.�6���m������ <t��ݗX���$�UZ������j!�����-��8A6�:�l��6ݛ���P�H$��P�M�M�	��l5YYMU�cZ�۶�t�I�8 ,��l ��  	@
���T�A�+@K�;m�6ݙ m�j��%;:ݶ ���� 8H�@�L����  $ ���    ��h-��}��|	�5� ��v�  �J����$�ְ  9ml�[r��]T4��QY�@9���Ĝ| ֊ɵ��	1m #]����i ��6�  ݪM���`    մ��t�a�j��v �n�  	6Ѯ�m�	i�z�?��E� ml�t�#  m�� ��ppn���7m�l�md�����U�^Z���*�#�k��۵l�o���& � �m&o���EH�-� %�#]���8,ss�]�� ��Lv*��ضyVH�v��V���<�T��lcX'�FҊ\�|�|�i�]��=̼�W�4��<�ר�Cln4knl�k��n��		���I�i��Y
[l  �p �+�����\��7��   �-�  $����6� l �mgj$�i$�[u �	E�mհ	$NkQA��}���[l�=: ��Z   �n          �l ��M�9�� H  :@ ,�r�� 6�m�� H
嶂���6ۃm� �  8    ���6�� �� sm�6�Ͱ�vU�N<�0    D��[M�a���xh��Ku� ��KM� $8��m��'e�v��n� �m���&��i"r��'R� �$ ���`�}��    ��� J�Ԏ�~�O�m�L�!���v�i��  �ݰ������f�
U�m�	2mfs"��۪�f�vٶ�f&��.M�H mz��9��r@�[&ؐ�Z�      �9�� H��ӭ6 %�m�][V��UJEʼ�����U �v�UQNEi[���� ���6�XX�-�� �ck5@��Δ-���-��a6�   Nm��d���݀ 6��)!�kՂĄ$[p6�%�m '@v�ڢ��i�#v��Ij�[N�UmK�l�f���jkK�9٪�nڥ�*�V3���+9V`�kvN&��5a��E�4�4���dY�p
�l8�����n@j��av��Y�+UJ�m���R��L�  �`��� -��	�6�  p ����` 9#�E@���>A�  �� ݷ�@ 	J� 6�n	$   ���`m�   Im�` 	$ڶ$t]��� m� $�6ٶ��� 6�l6ͰF�h����[�r@�lz� H��Lͱ�`v��   ��  ��pn�   fu������Z� �[��$    ��E$�V�m��I��m�� l-��  x  ����rT�U��^y�Q�¼��M���U6P��[l m�@  ���@  ��hn�m6�I�ph�@ ��R`����Iu�KU6U�x<U��U_��k��{rv5*� Np�'f��"v�*�ݴJ;m��v� [P�h  ڶ  �h  ��[@�� �  6�          [x��ض�h �H�����{�����?�`� (D���T�1�H'�|%�? �QH��(�N|m(6�T0"'�D~6���"�L���R(�R4�4@-�Gj�u��3=��(�XT*�u��]�v��H@�'P@�.��+`�`(� 3��PP�)�N
�4
)CH*�E6���a���z�B&P"�C�l�)��8&�%�0K� ˵P�(��� 6
l5�j
|lS�9D8��,Ad�0�d$]Az�m���ܨ�	�~@�Q	�?? 	ߘ�A�1��:�S@)�p ���� �M��(�A8:���EP�C��ظb�,G`� �t��>��D�(a��Pzd��g�4��Q/�A	�T�A�,0��� A_�v��DzU��fAU4(DC@f�x��G�D2��i��*tb��+��+�t�s�!�� 8��:�b	D�B)�M�V'4 ?� ��G�:�(@�FA,QH�Q@��A�+橋�c�1��9�s�	 ��Am�m�  �t����%�[[I�D��Tȑ�z6�lѬ�-�TU=�]�b�V��;����v��z��9�x
��ĩ���R��$��q[r�m[a����4݌kw{mE攳ۖI�Z�<�hg@[�go.ܢh6�5�c7gv�:��-pF��lڻj̗j�'��a��!t೨�b| l:t� ��U�,i6r�s��[n�2O��|^���e����V�Δy�C��[��nJ���������@��k(��3���ۛ����M6땺ڃ8eZ�H�-{n�흖�US)�8"���������v�cu�j[� e^j���c9p��b���av�F[��u����9�a�t�b�qe�@U<X]�d�Q�
��N���L;v������˧�R�If��t�8��\��g�l���Le�6��:��m+�UK��j���8-�=iyD�@�`Z��*���d��P�.�E���Z�ڤ�BCt��e��e���#>˰�qq�q�NM��mȽ<r���Z�ٓ�m�k���;]��T��E���)f%"045mjx���� tVJ�<�sR9��		V#��L����U��섩��4R�M�����-ۮ�Z�ʶ�Q���5^òj�[m����^kͻm� .3l��&�Xi)<m{��74��n8r/ ��s�2y['OU��`͔ �v0mR�ԫJ����4�]u6�2��[��L��x	V�i�H�|��ۭtȮ�m #;5V�P�ph�5�;k�a�94n1)2��iT����Ź��)��J����+%��Щ#]�t�l����uS�����L�[s&m�;GEV�/�wP=�	6���n��mS :0X�Vʯ#B�&ӮA�VU���*�ZY���@��J�@=�[v7=n�-���&n�t3pCR R�k�����H6C$�e)�m  *&L��)�".��S�DQ"�1RH?�4&ܣ�@Ch��؏�㢀�Fl�0p�]�L��\*j`���n-�Sc;�SNϞf���8^s`n.���$����3)��mJUPRv�n�㵒L厎Z�E&T��g���N#Bʒ&���[x]����Gkvx۬oX�g�r���ʷF6e�]v��s���s�i�!h��l�0�\�)���u�o$v2D�:�`ͼ��.f���XὍ*
iȎ�MK-Ը���-Ŧ.+�ݜm���o(x�w|�W���@nC�������n��P>����z�þ�b�7��?UZ��I((���>��؈�IlD(\ỷj���`�ݸ�6E���r4�7i ۊ��T�=$��RϺ<��XQ�[��Հw��, ����T�~��rMT���#*����st0�ͤ�&�=�Z�n*@6�,���E�Z��1�Z��T-%��tyv����2p�۬�֌�ks`�.,�8��ٹ�{f^�= #qR� ��p�I��䤩��(�*�7��-`a;L���N�ѩ!�n��ۯ ~��ln�[+v���� 	�j>��}j�9���ǲ�Ev��]� 7���?}�� '8� ۊ�L��^U�{{z^]���%�@?��H�T�'=���zx��mU��Kbv�@hMϧ�Pzػ�/7��<�4Γ][=1+��]�8�r�W�>����q`~���ۯ��^YP�%r��%��� �j�%�@z8���#)�Tq��� ;�v���x���#�(Q���1�O��B1�p��~���z5�wq`3y�=�6�eN�9n�햩��n*@��S2~�y�fٺV{HG qR |����x�%�ޥ���H�$���X�h-�q��6��F��m=ۡ�۳P8�ӓsr$��Uj�����, ��ۀ~�u��?ow�gc�e���U����5�� =T�m�H	I��@#��8ܷ ���ŀ~��,}�w w���>��-RD�v8�	�TҰ>x�X��XwX8�9
a
�H-h�:p�M^w>�X�w�,�V�en�V��q`wXu��`|�ڰ6"(��d�����]�\Ak�f^��vװ=:՝�Z��ctvnlY8��Vo�w����㛑6�c#w@5����ͫ�סD} ��VY�y��Sl�T�#����x���T�m�H��dҲ^^��n����^���H�T�9�t�� ��%$��Tv��������KT��qR�S̹��X|�*��XwX�w7g��׶�'9��ԓj�A~��D��BV�T��R� ��DH�ưH� ��)��0Q� @*aJ#�&��q��䒷�*B��^8���FG�o.B��Z1R��c'��cƷM�Mô;M�S9������i\��:�3�7*��K����Z��^{m������n���hI�9�;�)��ٕy����pl��svIg2rm\B���Kim�qڰ�C�뒭ˢ5�wTG!�:�m��<=m@g4��������K�,�����V��{;Q96�]wLk�x�Z}<e���z㇇����ה,Y��@#��8ܷ�n�,��q`�w w���>��-Q��lq��R�>x�_�������ڰ>x�V���V�ev�Հw��X�sP�
��*@z9�ʺͬ���R$��K�x����Ձ��j�����`3y�=�6�eN�9n�8*@z8� ۊ��5�G������Q�=�x�n�z�vn�[r7iM��뱇V*��K��8�0�cV�:��O� qR |����|*@�r*9i%�j�Հw��X%�s��=UC�A	0�Ѥ��^�� ��� ���X�>�O�]�&���ݤ ��@z8*@z8� ۊ�Ӵ�)b����r9n�{|\��*@6� ��@t˙R�2�ܱ�'m.�{��qM�����}p��K�o�m����eu;J����un4ټ������c��3��:ɔ�x�f�����{�����v�� ��@� ���X���"jU$l�Tݲ� ��ԔL�u�Vu�'1����i�n�*���p��m�?owJ)��@������n��jHo��|�j��+N9cV��V���R�9��=M@�2�Gm��v������ݸ�z����� ��kwe,��AKx�&��=����v��a�*�L�D����ӿ���G���W,N�? w����շ ���X_�ـn���B*�u֫�ʫ ��u{
�;�mXq�,;��ɳ���yI����ڭ�>�� �� ��@���'KٚQ�^�Y\�,�`{��rm��`�����XWbD%P�R�];V6����U]���7sq >sP�P�*@u�ݘ �3dZձ������7�
7��q�>'�sp��ۗ6�8���͵tvL���Hn�U�� }������:��� ��ۀ}�U�Zq��[��M��ѯъ�R"93���� ߷� ?}�� ~�;�j��ܪ�^� �1 >sP�K����v.���FKFӲ� ��ۀ~�u�@z8��~�Uo���zM�˽�2�Ҷ�/7P�-R��Hm�@�u`}�(�ș�]%4�UR
$�c6��^h��h�o)p۴];���X����J;P;����!�=`�.���h �2�n��4$����v�p�fSns)������ڶ���v(㡢��$mX9^�s�7�,���*�W@�:�`�PF�~;�m��:�o;�܏O�U|�/�n�9tJO�63g�g��Ɛ�n��ev[�vL����&���x��X����w�>E���\M<�u�=mɰ��Pu۫O�^-����M���e^��7,cdC���~�b�:�ݘ߻� ���ŀo���"��,�@�Z�ۘ�9�t�������#��-��e�߻� ���Ň�8����X��L�oڇd�Ka���s���"�[snj�D��ӎ']���V�wq`_�U<�����@{��H�s�]m��evų��sc12�S�n� ���7CùҖ�Npz�u�����n�m�����@y�*��~��O�T��*��F*ܴm;,��ݸ�Pq $��$�DI��Z�;��X����6�eQ�r��p���wLX���q�@���s*VfU�nYve�HI :㘀sP���ۥ�DX:���V���5$��wy���۵`jQ�����]�~�Wbjvk���>��dx��'��&���8ä���&�ŅZ^���Χc[����� ��RI :㘀�7��mNY-R�]�`�ub�s��l���X_�� ׻� �t�'6V�qMMU"iR�nՁ�x�gaWg�	Rgmc��c�3�T]*��T*�
�b]�u�d`@c4	��BH��0
p�@h�"�@5C��P���C� f4��FH�3�L���D�>ҝQ_���k�%t�di��6!�0e�B��� +���M��$>E2
5�G� �C�f� U�t�$���EG ��a�����TM�>��4kh6ώ��,-��U�YV�>�o� nﯸ��x��a�9�{�`k�kjiqQ'*����� ۚ��ds�R��*@u�3ߘ$���g�F�md���r�.n�mc�nuz��1�u�6M�;C1��u�a�6���nWZ�G-����,��o�/�u�}0�f�}p?>��E�$M�a9JVu���s�����
d׾����/%��>������er�Ձ�J맳`|�BR��|��`|���?wvaP��U�8� ;�v���V��	]KP$BJ#! XՍ�(mK�?wY��'�}��Nʜ�[-NKp��b�:�۳ ����:��@��ver�НvD���9�^���l$�����mj��y��7�kl;�dR	�
8�u�QaV w�ۀogu���0��b�5w�Z�V�ܪ�K37P㖀���HG5��������h:� ׽ـo�� n�n��׀j�[Wk�&	�+,�`�tŀ�ۇ�����<���_�wc�^RF9jl"j��I�{v�|{:�}!�����v'��_+ P����ow{�������׃e�k�\�;�W�xt�ҙ�K�ɓ6��f�����f��e�rH���\f ��#P�l�'U:���9��q�p7L-f���:��v
}f�Qg���\�r��]��ݚu�<Un�m�卷2�S�^������l/c��4�z�e�@!x���7�JB�v��q�6[��^���r���X�nW1�mh�rۄ.��ۘ��{�����/#U���5��m�m��mM�sۣ��	���˦���Y�ݖ�r"�1��$�`Vn�����& 'IJ��\�wf5
��l���v`��HI59hX�+*�6�73v�wL���)R �M@G�Z=ݘ�-�saGN�j,*�ݚ����& '8*@J�JEn�;K�-��w^�wf�n�X��p����k��K�%�*�n�7�X��R}�n�۴>�8m��V�{4Nx.��-�u�^�wf�n�X�ݿ��پx���<�j��V�l�7�ի�J�����@�v��5́׻�=���~��H�mC	ڪ���`<�9�b""˝��У���k ��|�`Ӗ;+���{;� w$��)R rM@yɈ����f��f�n �1 ��R rM@u���>{�ɱZ��1�Z�j�Y*.wG�n���^t��Ν��@��㗉Kr�D���6f�f��
��j�9��v`tZ��H:�� ;�5���& 8*@J�JEnʝ��;n����:�va��+��0iD�QL���7٣RI�{��I�����8��k� ��ـw�� 9&�:㘀�,�M���+p�l�`��b�<�I����o�׻� ��zx��mU��Whp���>�h�n�����sʊ,�>�K�g�&!z痵T0���_�7���>{ݘ^���wLX��r�jK%���m� ��>X-�X�ի ��_�
&N��Y��!I�0~��߷V,<�I�}�\���~}z��S�KW*��W,6%/7W���Ձ�x�a�,��P0@`��8�q{���߽��7�����u�Q4�Xq��63�����y`g[V����-Oѯ΄�� ,E�T��M��ێPwkpvv��t��E��YFIg ����}�}��������5�{�`=���n�^������ ��ޯ[V�1�f��|�y$��_��X�z����#&�UEc��If߷V, �۷ ��v`=���b�E-M��v�� �M@u�1���)R�]r�jK%���m� ��v`�v{w� �uZ��u`
��!7�y.�w�"�/q�KZ���X0��vfw6�`Ӷ��$a�4�,p���#N�v4�1���[rg��!'�M7!�ab�J��k�	���07&6��T�l%cxx��vr��L��GAd�CɅ��8���5e3�����zڭ��ѴҺwL��ն��m͗r�/1��+�����tYf�\ԍ`��:�)�7�\9��*���]�����k8ݾ�����%�ɳ/N�Z���ۧuX�u���uі�@�[��=}۾�.V�����n|��r�ζ�Xu���N���o��Nʜ�Z�����n��{��I%#��$�{�_ߛo_��cm���g�ͷ�6	�A�$��ڇU�6�}�v���n�U����#��]ݼ��
����~u+�Gm#����m����o����m�n��6�}�v���{�7�#�"�,c�Lm��������7VCm��柿6�^�)������m��㨈q��vv��]��.:�>���2:.�:�:95v��=R͝TV1X(�~��}��!����柿6�^�)����ݟ�6��Ŋ)mCH\��&������{��A�h�00g!������ތj�oq�;���y���� ����э�Yf�~~ ���o�����K�M���cm�����ͷ�ݘD�,nJH�iq���]���m�6����?~m�q.G��m�����BT��-���~m��Ր��~�}���m�o���}w_�ͷ��kz����O]G4�ck��v�c=-ۭ�l�fM��뱌��L�BY��xw�!WWi�?����柿6��ݯm�����ѷ���6���痗�Gm$-��Ͷ��k�DD(��US-׽?}33���\����]��ޒ?z���:⣖XG]��m����{����hƭ� hth!������Ͷ����m��3g�TV1X(�~����}}��1����ߛm�n׍�rN������ݯ�b������*��o�4����=���6�w޿�6޽���}��GGc�-"j�V+�DӧiRz�d��/i%z(,���ړ���_�IfE�S�m�o���o�۷���׺b��#o�����m������IGZ�����o���3.\��Wwv�P�����������������e��~~ K�U�������wwq��Www~�7޻��v��A�$��ڋ
�6���柿7m�3��Km�w���m�s�,� � �"�!!#!��R V� $�*���c��d1����=��Q��,R�~��n�U�����������8,�ݾ�� ��ʹ���z��p4�u�2<�J]�Wq���u��M4%Y2s�:�n��vU1���{������m����y$��6��ئ6��7��UX�`��[��m�wL�y$�����g�ߛo_��cm����ߛo�b���QN9Km��ni��m���߸��{��7}~m��������
���Y[�v�~��}��m��{�����6����x������MB�$VD2�a�������wn�b�����wwq��Wm�~S� ȤI>�|�	NB��0�R$:��(Gm�ȆCbI �H�!)f!$$b(� �΄���X1#@�{�H�R$�XDBH����r�4�>���$�eF$BTp�A�Y!ĂE`�0I|�e=�>��DѢB$X�`��4 (SE�0� c��F#�%��r�(C
$f�Ba,B#��f-B,!	"E�E��HHD��!#4|	:�Pr��1�Iń`B�e1`@���zW$�
~b(a�4��(;�2�R�Xő��d��Ϥ./ 4�P#ݸb@FFl��`��0FY�D�I���Y�!2�$,���fVA� 2�!��H�$�P�c���bH��"@�tI"D�0 ā�����"�d��|iJ$�F @ A��$H! �P�(B����ߝ�HpH�JP�[V�m�m� pIk�p[S�����Q ��m0��IiRMn���Q,�q��T�h��m�Z�+��������n7��θ��s���ܻ�3���d
!��i�θhRU�L�d�Xț�����%��偧&ūn�f�:�Ⱦ5�@ݱ�s�/#�����V����Ѝ]�R�`�A��iP�� ����r,�:㜩;krn�� �D�X�(G5�nP}i1���pU��v��خ���c�mW�.bj�6vg!Y�Vʥ9�N�!0�UHS8ɟmȽ�:%����yGj��R�!�Z	���v�,:j��%*��籕�J�JN���
�L��I�]��tEUu�K�v��tض���dɹ�םgt�F����"9����8�E0x� &�cn;Sʎ^w>ڱM���A�6�(��jT7Z45{+�T�'[/:ᔝ��l�ёٵ���*�G+ʪԫ9����+���g�Ȣ��$�.d���v��S!r�R���X��<F�۲n�5�>.����V:NN��!�j���A�]�����F�01�1j��b&����dldF�s�mf#���Tl^N$B��k����m�I��t%���iwI�̝;"O6�4��mv��,n٘��"���T�lx9�k4��;9%R�J���mY��z��:�l��My�V	U�[v	J�x��!>��[UZ��&0p#]����]!���N�,�A�Vg8�UjBU�j]���7 *�j�㓪���)@Q�X����k��EY흮�$ԮwJS�(����V��:���볰.sK�3�۰�e��ʦ���G;n������U9z%���tô�����g�j]�5*]lR�Thu[/�]�8_�i����We�
�����2�T���5\����uU9��m�[F�+�Cr��U���լ�ZW�a�Oc3Ё7I-��d�J�j�pdm� ��lJ��*&�u��M �|��(�b*tplt�!���Nޟ\���ٳ�9�4�=<tY7:pj	뚵��qfr;��&�{ڬ&�ڌVb�������v���$�z�C�L�2��k���ɬN�2���BA�1��K0���FS��Ұ����q�f66:;;���o4-u��;�-��������ҍ�k#k�}�w��N��L�l����f��]���Խ��6��\�d���݉���wy����t��:��}�>�ϖ{td�[�_5��������.\�6�X��rKS<�?����U����j����
���G3޻��҉�A�$��؋
�6���i��������m������6�������Zr�i��m�n�1����o�����^��1���sǒ�����o�-��G-���a����}~m���cm��sOߛo�w!�������ʪ�b�R9-������)�����?~m���^6���?����O�/��ݦ���].�
��l9��Pmv���-���3�-]6W+�<ڝ�()�)T��}�柿6��ݯm��v���z�LSm���pU5���	s�fov��w���4��0��"D@2!��0�p�3���s}뻹n
�]�ۍC���Ufe������IIe�6�{�������b�����wv�E����p��/*��m�6忿6�_t�1��w���ͷٻ��ߗ�o������=D����!c�"©�����?~m��܆6�}��������)����@wg�㴭���evųy�,fV7�u]�Cvv�붶^c0掋����q9k��O�m���Cm�x��frq���I%�U3;�}33�W��RXjG;� ��������-r�fe�>�fg8��z��\{��y�UU�V
G%��6ߟ��Sm�{�~�~q�#W^q���X���{��;ݶ�رIjv����J�6���q[��}�~�����m������o�{�{ߔ�����ú�Z��)�����F���x��o�6���q��w���Ͷ�p�S��U�VrE��v:۲d2��<딸�k��z�Ó�&�A_�z���<y�[gS;�m���_ߛl�M�q��w���Ͼ��M�Cm�����9j��m�6忿6����璒7�����m�o��m�{���Iy�/c$q�X텵�q���s��ͷ�����${�������?K���s���"Z6�����ߧ���1���o���l����շ�4֨VH
���WX﻿M��}ܖ�Ƴ�\�[c���m��v���g�^������?~m��܆6�٭c@���2X�)3B3�
�uz�4@$�mqة��u�a��7]t���-~~ o����| 8�=�.師��ێo�ww-̥Y�z���NZ��o�����)#��b���o� }�{p۷\M�mdC�4@H� 㚀=%�@8���iT��(�!l� ;�ۀ�^�ǰ@H�l*�ݭ̼���L�*���Ձ��ޟ��Հc�Z�T�O��QL.����|z��.B�l�M\��/n��X�V�-�碻i�� Bcq�ÝyÙ��=n����l��aq�2�1�-��1�L�vŷX��<IE@�1d{v끂���,�dvs8���Kp�n��H�Otjq)ם�8�Z�-���{���ݍ�(�ٺ@�v_�>��t*���lW-87�s�݉�ƑA�N{;U�q5����';��%33f,����/Ƶ!�3�g5�഼+��K�jݸ�s��vv��\���y�c���nøv�n�"�4i��`�ei`7�Հc�^�����Ձփ_��,Q�F��� ����q6������ ���~��L�8��/��@9��\��`�q�X�t�LMZB:V�r[���n �� qR q�@I&R��ݫ��V�ʼͽ��`�q�H�5 yǷ >�M�E���#���ȝ@�ݽ�mWS��zkp��ۜ�U��E�ղ�NDV�[��YE��	�`�sPGsP{t�>viP��(�%�� ;���l��0�'Y.9{�I;�3ـoݺg���g�@=���c��cw�����@>��@�s�܅�9e���p��L~�� >����}����`�v�UUUQ`gr�`jS��� �s�`g]� ���ǰ�("X�Y+��G]S�olcd�r�,�`�v�n:M���p��[`es�:�z/7w//ot@�����`�߻t�>[��bj�Gb�H� >�˫؈J!)��,�ZX<u`|�ŉ��-઀���ۦ�v���ʥ����p����?n�p�Խ��v������ 8����8��s��ݞ�j7%D�� �����`����~�߯���~��Ӣ�m\����]�l:5��t;%�� ����%�r;l�W5n��������`����7 ��h��,q�+-d�ۀw{t�'=� q�@�@y�;�j�ܬ��˭���9��j ��j��0����+�*9m�ʰ<��q�׵`{;V<�X(��Bqk."9�N��`���e�8X�R9-���{�@9�����j���Jq�]h��I��1`o]�g�a��틴g3�^��W5ۮv7|�o�s� �������j:�-UYL~�� >����׷ ��t�>l���drQ�KSTX^:��˫5(��^mi`>��n�rGjn9m�6����M��� �j�t*��r��
�ݳ7ou �l�� tsP�׷ �K8�~�dZ� �[��n%m�q�,���3�/�9�Kkܹ�u�B`��:�}q��U7[lGʫr\�՝��YN�'c�����L�"P�5�u��^v!�v�d���,�E�sl�Zv��6��^6�z�(C�#q�����rB�:���l��g�'sIմ٬�l/ ��5˲�yݍc����tH��h�9ŞK��=Yn�n��+��Kߺ��k�uJYNR��ظx��]��cnz�v�K��m�`Q��7m'`�-����n���n }�{p��L�u7��㊎[c��L ����M�s� B\3(�*ԎKp��ۀw�`�n���n�wb��-R�*�9+��}6	�`�:9�?�Wo�j���SQ�+�TIe0��L �{�`�Vu�,��3I�T�\ջN���̽;��c��'U�mGj-�&�^���?Ϲ�M<$�|�I"�!��> ��\ �5 �l��#�bͽ��lm�p��ĵo�\K��~�g� ${ 㚀��
��ܼ�·7l�*j��v��S,��dǻV��� ��z��؝����V߻t�����˫�������۩U'9\��v���� ���=?��b�7��0�6�h7��4ܲ�gι��5�a�v
]���V��k�7Y[��/�q����Kc���#���y����1��""�� �������+S�U.U"���7�T����M@K�M��6}�_8*���`�����jI7��:�ع������y�jS*Dp[~���)��d.7D5��|!�)�&8���WC � ���a#�fwJ���&�55�D�xd1d�����)�G;W+~���� �&&0(d�ϝ}�M�u\�QAڪ}C�%o��T�B��U*!�x�G �E٠ �����'����b�>t�7�d�+"l���~�P��؀���*@{�p��QGm�6�_�l�=�o�/�o�֬:�XQ	(Y�&uL�d�EW'����hӍm���z��j��<n^���XT�q:�Ux19`�AYk����w��Xu�H���w�& <��V]�U����7i��H���w�& :8���M�V�'+�X�� ;���:�[�q��}� �ذ��valvǆ�m�e�n��R�T�q�H=��7f��'j��^DYUx���*@;�1 �:����>�uu�l��3��Knэ����G��t۬zϜ��-ʼ��7K熘w\rU��~m���� ���玥�:8����]��I"�!�ʰ��f�v�0��� �����h�C��7,�9͔ :8��EH�%�=�2�dnH+mt��Ͼ�~Xw�ŀw����Q�~���GdE�P�KJ��7j��IfV��=�E�޷j�0ȡ��)H(��c
�
�BD�H�Q"-� ��"�D�\�%ȹϔ�nIKPZq��p��������������s�b��Ƃ�{m�J�9s��n
��N�rv{.q�N 8�\ɹ�aڥ�HU��;Y�4��Hm�V�B����6���-���v�:vN��h��x_%��&Ħ�sՍ����1��t^�ؐ�.ىY����\G�n~�>,����"��vb�=�q�1iu5#�{P�5�7*���V^[��j��ĸ�\���ҖZ�H�D�#��&;�碝�:���m�-�λ$����VNW,���Vݞ׀}ݺ�t���T�uØ��7n�ܭ���6����_���T��"�vH���X���
� �� ���Xq�Vz%�s���M���M��:s��� �`��,��u��կ����� ���T�%�H��d���$��>�__�n|� ㊐x�l�Z�,�B�`Ik�C���{U�`}/���s�nyͮC[NػsmPa	���cT��O�=tl��;V<v����7g ���?dnH+mi�W�}�wU��-~Y�
KЗz{;�V�=�`c�k�;���0Q��ȝ�`��,��T)�����Vx�]Ԫ�r�e�J�>^���@�m<��v�ğw��`]7�Ikp�V�rV�}��������y%�0?�S��i���#Jm^ݐ+�)v�n�v{�u�U��2i�ࡿ{��}ù�]��نf�r|��qR�$���c�n�����R�im`Yj�?}�ŀ~}ݘ�}ݸ����$��z��l�JH�Gj�>{�L�}ݸs����  � `�B*!b$����JQ�}	j�:����{j��`d�C�ڛ�`3���;��0�n���g�� �=�~��$����nn�M��������>��&�>�@wfW]�W�9쎐�>J�0�7N�.��v6����y'[f�VWkZ%جV^����[s���zç��n�7�VNW,�¹V��vg����ڀ��� 9��&#ksv�Cr��r�wP�������������nŉ�Z��W�6�ˋ�G��ŀ�}j�3�Շ�[SU.�X�6XKd�X�S ���X�{�z� �}�}��`��l��m����u�ܗc��흊�u��\��n�Ǖ��eS��K8Ag�̸�-��Y��_�7����M@t{s��31a�Yy���y���&��]���s�H�۞�f��'��I
I[�[�w��s���5 z9��C0�f��Q�*��{���|�ޘ�{�ˉ�w<`�&��+'+�X�YU���|�<�{�k�1�����`J��_�"�}$Q}��G�3����k^x��qq��zM�+��f�{K=cO�|9��v� ����ut����ۇ3ˊP�8�m*hb�Rۭ�.�T�]���r�����@�1u�G�l�m+��Di�k��.ڧ�i^�S�!9gB�Ύ5���]L�'�ix#�vyC�۫Plk��%�hs^�u�خ��Z�k��qX�3]3�u\nr�+͋���z���ϻ���m�v�d�����][Y;9M�5z��)`�|��F�6����{����X����%?����o`�|��Ɉ	�e*�	Ij�M�n�{t��%��.%!���N�ܰ�^��L��7Up&�Ue�nf����� =nL@�j�ۦ���u���,�j[Ls��x�y`�Ձ��e��/BP���X�������m�Kf }���>�ls`���1 ��+&f���Wzg�r����85� �\L:�S�:WH���:,/J����w#t�B�V����K�t� ηZ�#�ڰ5�Ӝ&2��Q�i�~��2$�ԗ�$�a(���YN���V^S/R�2n�7�-m�W,u�m� o}�w�PT���L�mnn��V�IUUa�%3��X�mXc�XjQ�����>�)\�&�*m�p��Ձ�K�oO�nՀw1Հf1���j���-��r^ܺ4�nu�%c6.{q��N؜9�ݖ�r����W���b����6�׀��� �j ��:8���v�|�9"���m0�n��8�ww� �ذ�ۦy.6w�����򪪦yUV��XyL��Q!D�B�DD)G:�`u��w.�ML���In���ߖ��|`~ݸ�%�7����W�1Khܠ��TX7L�<�K�����`u�2Ϳ=�?�T�v�HUh%���0�s` �=���	�ڷ�-�X���<}�tf���n� �� 6�:=��]0�vaU���,U���{ݹ�	z��{���3�Ձ�[�-��bLv���� ��t�ɳ{�\ ��\��V���-�j�؉���`7j�31Յp�P�!#HD��Á��1{���{�D�,�J:������p�%�������Հ��g&'T��U��u�!�H�������/��n���nx��}6r�vnn$j���o������v��Lߤ��`8�)��5<�*yʙ9ʫ����p��x�~���v��\�l���!R�PQ��V�֖�n��[ڰ3^ڰ7��Ֆ� ��;%v��q.&����oj���j��w6��;��唦��u��+n���@���*@N����u$��:�E���^��E �]�#� 6h����6eS+���!��9	x&�(�W�A ��X�r��bŃ�*��h��0�F�F+PwJ�l2�B$\. C�s}ǒ1ȡ�)�A�*�T��0"��b��v����ȨM�Ls�6���5��8E`DtZ�#$"�5�8|�09\:���2����ۦq��# �A���~23�I|���$�B|G+y$]�[m���@-�R��ڶ�l� �֝���i!V�KP�E.^vU�b�IWR�l-��w+����U �N��wc��E`�d��7�;s�g�<�)ru�6��C����4v�s{��=e&�d\kAî�<�T.n�WPTt�)l���I�u�E���=	�;���l�pRZa-i�$�ְD�r4�y��C�s��&/lr�6�vU��l��G��og�ml;ӎ:��m�h�|vبA����ێ��i��j�}Ѐ��,c��q�݀60��ݻ*�7-�J�e��
ZP
Nؚ����)kg��^ݰ���bCvͳ��n�b�{rM��64�h����6�YU�8��`s�UUJ�ӭ��
�uP1�Κ�Iuscc��]$�z�PT�=������OZ�t6�nq��.y�7c�[�#'�E�,'6;0S+�"1{crG6;pm:��ؕpH+j󶩻U)�F2�BE��LD���u�j�p�B�:W6�j˄��m�I鉩�-T�d�����f���<�N��\��b�g9��u�`�s�9G)�v6�gk҃�� �u1\0gh��&� H[2��V��v:��4�5ө�M�tm�q��S�r �ԡX�ڨ)��yYY�j��������Jg�ds�v�oke4"�q����ʁ���*� ڹ��G)@Q�i.�Vn�ۭfݭ�;���qZ�mF�I y�Y$!���6�+���v ����uU*�J���:���iV�-�*�������J����.f	=v��Yڀ�n��R�F��<�,��l�Jݳ�$�ِ�s��	�Y	�dfVwm��;a�[;*��ҭJ[\�(�&�����b�a���@F{j g�z𷙵t��v$��C�Zg��� :���
����R�U*�J[H �F�Ca�j��<��*�U�U\�[A���hm�e�m�.ӯg��v�� �\�6�w4��\�zꉙ�;l���Y��ƽX��7mfie����{{���w���Qq�s�DR=@�	���b<hX��ɓh|��N��pMg&LLb�bLfٗ5�@険����sc����f;5� �lkA��5x�!���<�5qϳrv�g���;`�&��
��9*�{.��y�sD������L�p����Zv�8�B�����7BON�W��[Χۘ���sk�!˹뒥1��,�ܨ<��1
vP�g:&x�nHe�nvG�H��8��6�=��[kL��^b�I�;(��g��(5tlu
���:���wz�|#���ld�Š�k��y���ŗM^T�m�{}� ߶��v�~`{w� �����IYaY�*�7�@�������9���s2�o0�7t@����@tqR�m� �z\��N�-����9�{Vk�Vu�,6&^nՀ��qK$qJ��-�>��,�m� ;�����p��F���)K"E��u�s���nr;�k�|����'��m�iڰ�q:���HB�e	+vʿ����v��ݸ��ŀw��Ֆ� ��;%y�f���w����Pxd
I%�ˀ}��X~ۦyq6}�zL
����R����׵`u�g�^mi`���?}ݙk���!^T۶�'�o�R?�� >�Pnj�9W(�3S�P��`��0��߷o��v�ow w��R��"«\��C�oI����'U�v�kAr]�ͳ���n��qŖ����BB�`q3��}�_�&q3��y��:Mı,K��h?$�&"X�'��_��q,K���I\o3.qq��9͸�s��Kı/=�gI��%�b{���&�X�%��{^�Mı,K���t��bX�'^v���..f�9�Γq,K��{�Mı,K���4��c��8�Ģ� y����K����&�X�%�w�����g8�����B�����YfM&�X�~@�������Mı,K�����n%�bX��ﳤ�Kı=��f�q,K��|[�������.q���3I��%�b_s�Γq,K���}�&�X�%����4��bX�'y�zi7ı,Nz>��ĸ�s�)�Ҝͧ�����ۘ=�'0��P�lN�Y.K^:��e�^�>�~'��u�����t��bX�'��l�n%�bX����Kı/��gI��%�N/���m����
�ݷ8�L�g����4��bX�'y�zi7ı,K�{��n%�bX��ﳤ�OɊ�8���{�?�u��+,�8�L�,Ow��M&�X�%�}�{:Mı�1���gI��%�b~��l�l�g8���ݞ"jH�v�8�D�,K���t��bX�%���7ı,Ow�٤�K��X!#��"|��}����I��%�b~�~�~�囉���ߛ�oq���^{�Γq,K��{�Mı,K���4��bX�%�=��7ı,O�������������������l=�y��ݛ�]�z��6f{!ss ]��＾/�73q�ً��I�Kı?{��4��bX�'y�zi7ı,K�{��n%�bX��ﳤ�Kı9óؘ�3e+������g8�Ž�x�/��
#1,K���gI��%�b^����7ı,Ow���n%�bX��~�Z�P�X��L��q3��LK�{��n%�bX������KlK��4��bX�'9�zi7ı��|��������m�/�8���^s�Γq,K�绯M&�X�%��{^�Mı,lK�{��n%�g8�����H�	hU7e����g�b{�צ�q,K��=�M&�X�%�}�{:Mı,K��t��bX�$�!�� B
��c�"�42z�e���,dp3gr�j�8��6�y#��uc��g�@v�ۘ��sEY�طmьr�B�n���7l��H͹�vڱ���T����ۄҬA�@�%i��|;V����nn�Q�	s������g�i��sI;,�78���OYmk7Ohے�d�ԙ#��lAI���od����ؽ�v�{0�8�z��kQӖͲG..�͡*Pn�5{�}�;��/�����-��j�v�1�n�:�v����X�;s�{��k���gZ��Y+�:�4"���}��ŉbX��}�&�X�%�}�{:Mı,K��t����1ı?{��g㉜L�g��O�'�`䥲gI��%�b_s�Γp� �LD�/{��t��bX�'�{_��q,K��=��7Kı9��}q��d���s��6�9Γq,Kļ罝&�X�%���^�Mı�ű9�{)�$�Os�Δ�I�8��[.!q-��j	 ��u��Kı9�{zMı,K���t��bX�%���7�&q3��Zz
~R���k�����q,K�����Kİ���t��bX�%���7ı,Ow���n!������m��i��h��"���gKd�4$%9�k�:I�;v<]�Y61�yz�.P����.q���:Mı,K���t��bX�%���7ı,Ow���~"},K���zMı,K��n����4�g&ifs��7ı,K�w��n@����'��zi7ı,O��l�n%�bX������Vĳ��_w}���V*Ъm�s����'��{�M&�X�%��{�4��bX�%�=��7ı,K�w��n%�N&q}�kɅ���QYm3����+�;�{f�q,Kľ罝&�X�%�y��:Mı,K��4��b���/�u��[���YVq~8��bX������Kı/=�gI��%�bs�צ�q,K��=�Mı��&�u��Qy��T%,j��8�ﺹ��f�p���a����y�6s�ŷgk��
��7M��.3��9��v�D�,K���gI��%�bs�צ�q,K��=�Mı,K���t��bX�'^���&qqq��͘��t��bX�'=�zi7�*G1��~٤�K�������:Mı,K���gI���f"b%8�W��)�KhJ��i�_�&q3���k��n%�bX������K���p�'�"n%ƾ��&�X�%��=��I��%�bw�-��31�\���f�q,KĽ罝&�X�%�y��:Mı,K��4��bX�&"{���i7ı,Nw��O��3L�rf�g9Γq,Kļ�}�&�X�%��w^�Mı,K���i7ı,K�{��n%�bX��̽q���v�q��Œ�Wm�8����i���[mVNgF��pPȷTkOknx
��~oqı9���I��%�bw���&�X�%�{�{:ı,K���t��N&q3��o�^L-eV���i�_�+ı;�{f�p� �1ľ����n%�bX����:Mı,K��4���Rb&"X��}p~�����qs�L�&�q,Kľ����n%�bX��ﳤ�Kı9���I��%�bw�����g8���hz��Wc��m��s��K�,K�w��n%�bX��u��Kı;�k�I��%������#�7"kZ���7ı,O>���X㒵-dr���q3��L��=4��bX�������%�b_w���7ı,K�w��n%�bX�����_Ȋ�C�r��uŝp�V�kq�t�vr��״K۷u�,�8I�N�	/9.sns���Kı;�k�I��%�b^��Γq,Kļ�}�
��bX�'=�zi7ı,O{Է��\8���q���3I��%�b^��Γq,K��=�cI��%�bs�צ�q,K��=�M&�~"�&"X���=T���U*�%UU���$)!I	���Zn%�bX��u��K�D�Ow��M&�X�%�}�߳��Kı>�}�[YF�����g㉜LI&qs�צ�q,K��=�M&�X�%�{�{:Mı,�$�N���cI��%8���{�5��Z�J���8�L�,N����n%�bX+{�{:Mı,K��}�&�X�%��w^�MĲ����J<���W��<��P�����.�Mȷ&+۹����t3F9gg�ٷ��&�v�t^d�$ݤX]�:C�%�$����-��$���ڔ�#&��7a�޺����B�sΕj���bֶ�n�uġ\`���[���W<��C�-���-*�m�8ڀ��	��6x�VP#\[6��h3��=�`���(X�&:۳/i��T*�2�i�����S������93���ɂ�z�ܞ�ت��v���n���\T���0"�*�AY	,vB�o�8���'���]&�X�%��{�Ɠq,K�绯M��bX�'y�zi7ı,N{����ㄑ��j�������ow��}�&�X�%��w^�Mı,K���4��bX�%�=��7ı,�{������c�)i�������d绯M&�X�%��{^�Mı,K? �ǻ��t�D�,K�����n%��&q|����YJ����q~8��ı;�k�I��%�b^��Γq,K��=�cI��%����w^�M�7���{�N���|�)b����{�KĽ罝&�X�%��{�Ɠq,K�绯M&�X�%��{^�M�g8���8�����m7ld�ٶ�vp��+���k�':{�qY��f. e���|�ݲ�m�-U�[nq~8���&qv{}3�q,K�绯M&�X�%��{^�� O�b%�b_w���7ı,N￿+k
۱Cv���q3��L��w^�M�`U]���v��!9<�蚉b}�k�I��%�b^{�Γq,K��=�cI���S,Nb{�Oœ9�&s!��8ɤ�Kı=���4��bX�%�=��7��,Nc��4��bX�'=�l�n%�bX�v��VBK������g8��{�{:Mı,K��}�&�X�%��w�4��bX6'y�zi7ı,N�P�	��m��-����g8�Ø�}�&�X�%���{�Ɠ�%�b{���i7ı,K�{��n%�g8�7b����2�R�1���Mѻb��Ѯp�L@�v9�=�:-�n]��Σ��)c�Kfq~8���&qw���8�	bX�'y�zi7ı,N��4��bX�'1�{Mı,K�	=��72�C7\��n%�bX����?D1,Oc��cI��%�bw�~Ɠq,K���Mı,K��+��ls���%v�8�L�g8�wޚMı,K����&�X�~S�2lP�cg�Ot)���gL��(`0�O�dC
4�� ��;�p���5�F ������f���p@��$ �iX���R2Pba��H%�U��ɔ����� �� Y�I!ġ��%V�vR�����R�-��� ځ����G��
�'�#�	�T�wx�&@�
c���QSJ�D�\�N(<�:���ND�5��&�X�%���^�Mı,K���D�rg8����8�n%�g� �'s���i7ı,N���Mı,K���4��bX�'q�{���g8���wߕV�[v"��q��Kı9��f�q,K��0{��M'�,K��;��4��bX�qv{ޙ���g8���o��,Q�j��<�n�wnmڵ�r�-nk��a�,8p��l���^:�E�my⛾�~oq���;�k�I��%�bw����Kı9�{�Л�bX�'=�l�n%�b3���爟%��Ƭ���/�8��bw����Kı9�{��n%�bX��}�I��%�bw�צ�q�3���/B?��m��[3����&p�9�{��n%�bX��}�I��%�bw�צ�q,K��9�cI��%�g��?~��;h���%����g'=�l�n%�bX����Kı;�{��n%�`u�>��P!*����b]o�Γq,K�/.���?Ye���g㉜L�q=�k�I��%�bw����Kı/��gI��%�bs���&�X�%8��ĸ��h{�D���!���;m
�R]A`\l;�t]���n7������	Y����p|���%+�J�q|q3��L�����7ı,K�{��n%�bX��}�I��%�b{�צ�q,K��;.��s��`�[��Mı,K���t���bX��}�I��%�b{�צ�q,K��9�cI��%�b}��fs2̓83Hd��9�n%�bX��}�I��%�b{�צ�q,��9�cI��%�b_w�Γq,K���)�ɜٓ&\9�M&�X�%���^�Mı,K�罍&�X�%�}�{:Mı,EB���Mı,K8����,��5d-�q~8���'���t��bX��B8��߳��%�bX����4��bX�'��zi7�L�g�KW4_�~_̶�K\�d�d.�L���s�-��-�7
���Vm�L0�6�v����c��X��+{v ��S��Y�''P�ݱ$��g��tj\�ٶ��mQV.ؚCvA���7\moZA�Xm�(�6�p�/;���c]���Z��{7���UǛ�W`,695v�D����e7E�L��C��Ɛq7`:i���i�nk��* =���6���w��/w��n��\5�.��rH��;�ǯ`͵���n�vcr0��86�e�����ݺrc�A�-��nqt�g8������s��%�bs���&�X�%���^�Mı,K���t��bX�'N���&qqs���͹�s��Kı9��f�q,K��}�M'�ꘉbX����:Mı,K�����n'�"(8���'��~?Lo8�����̗94��bX�'�~���Kı/y�gI��?����{���7ı,N���Mĳ�oq�������ߔ��E,U��~oq��A,K�{��n%�bX������Kı9��f�q,K��}�M&�&q3��]���$U4�m�/�X�%�}�{:Mı,K ��Mı,K���4��bX�%�=��㉜L�g}�����XԶ&�ntbѷ=N�q�9��޺xx�Iv���Ht���(Pv*�A�[�_�&q3��]��f�q,K��}�M&�X�%�{�{:��&"X�%��߳��Kı9���?f�L�2��s4��bX�'��zi7�&��
�&"X�����n%�bX������Kı9���I��%�b{��.`�s��a����i7ı,K�{��n%�bX������Kı9���I��%�b{�צ�q,K��Ob�cw9�%��s���8�n%�bX������Kı9���I��%�b{�צ�q,K [�罍&�X�%�ӽo���\\�0�qsnq��7ı,N{���n%�bX����Kı;�{��n%�bX������Kı;Н�5<g=/�vu�B�\���c��=b�>S��v��Ѝ�������4���o�ߛ�d�,Ow���n%�bX��=�i7ı,K���Ю�X�%��w^�M�7���{���Ӄ��)6�H�}����ı;�{��n%�bX������Kı9���I��%�b{�צ�qı,Ns��z�6bL���q��Kı/��gI��%�bs�צ�q,y�~b`�MD���M&�X�%��n�.�)!I
H]ǿ*��T��Pp,��t��bX�b{�צ�q,K��}�M&�X�%��s�Ɠq,K�������|B�����=�W��4�e��g9�Mı,K���4��bX�'��{Mı,K���t��bX�'��zi7ı,O��'������C�׬nѼN�V��tZ�����$�Oi��Z5���b�QGKi�Ȗ%�b1���Mı,K���t��bX�'��zi7ı,Ow���㉜L�gwS~	?;de��m��Kı/��gI�%�bX��u��Kı=�k�I��%�b_s�Γq?����bx���x����sg6�Γq,K���k��n%�bX����K�,K�{��n%�bX������Kı;�O>�󛛛�L��\g3I��%�b{�צ�q,Kľ罝&�X�%�}�{:Mı,����>Oc�l ��?g���Mı�{���?Ã��ȇũ�&�ߛ�o%��{��n%�bX�}�{:Mı,K��4��bX�'��l�n%��{���~�~�~�%p#�\�䫇�7k��Y������a,nxK4�.5�#^ z�s���3��Kı/��gI��%�b{�צ�q,K�����A蘉bX�������bX�';��2c38��̘��c9�n%�bX��u��Kı=�{f�q,K��=��7ı,K�{��n$�PI��ҟ�&$�����SPI��~ѡ$D���SPI�K�w��n%�bX��u��Kı<sڔ�I���9qs3��Mı,K�﷤�Kı/��gI��%�b{�צ�q,K,Ow}�g㉜L�gw|IOηZ��b�:Mı,K���t��bX�'��zi7ı,Os�٤�Kı=��zMı,K[Q;����Ę�s���������t�ٲWX �q3p���ݨ��z\θz�IwgMy7Y�7eHN�X{n�y���%�hK���Ē���ʱ"�X�+vѶ ��.��J�v�v�h���v��9��`ۮ��7�ɓ���u+��3E�&��v<rv��۬@�^"�{0���x&��H�ͷ ��g���q���b��j\�GDJ ����bIg01���*V�1]�{:w[e�n�ٻ7U�����c(�t� ���w���|���M}��oq��K��^�Mı,K���i7ı,K�w��n%�bX������Kı8t�}��777�̸�f�q,K����Mı,K���t��bX�%����7ı,Ow���nX�%����7������78ɤ�Kı/��gI��%�b_{�Γq,D�O���M&�X�%�����4��bX�'1�[���f$n	�ٜ�:Mı,��ED��߿gI��%�b~���i7ı,O{���n%�bX����q~8���&q}���al�dN�Lg:Mı,K��4��bX�'��l�n%�bX������Kı/��\��q3��L�ݾrEBH������p�yW��v��6�ܺOZ"䤃�������E�.��j�{�7���{������Kı/��gI��%�b_{�Γq,K��{�M&�X�%���ԧ�b��1s�39��n%�bX������>4���&bX�����Kı=���I��%�b{���=�����ow����5������X�%�}��:Mı,K��4��c�a������l�n%�bX��\��q3��L�ջ��б�mu���t��bY� �������Mı,K�}�f�q,Kľ罝&�X�%�}��:Mı,K�:O8�󛛜b�̸�f�q,K��;�Mı,K�)S���t�D�,K��gI��%�b{�צ�q,K��$�[0Ba	�'n�Xt���;mos�Yӥ�v���guƶ��tp]R>f ���n%�bX������Kı/��gI��%�b{�צ�q,K��;�M&�X�%��s��Ǳ�P�&Kfs��7ı,K�w��n*�bX�'��zi7ı,Os���n%�bX����q~8���&q}���ev0v"�%��s��Kı=���I��%�b{�צ�q,b�t
1D�1"�E�P`�>ʫ�Y\�c��X
a�	P!�Q�C�?�����:�bj%����&�X�%�y��Γq,Jq3����ד+��u@��g㉜V~B"~����q,KĿ���t��bX�%����7ı,Ow���n%�bX�=�J{&3�.r��g9�Mı,K���t��bX�� "��?~��:O�X�%������Kı=�k�I��%�bE�'%��!��*9*4�9gngY=�m��ݤ�WM�u���y�=V�V\9X��L�U�����{�K���t��bX�'��zi7ı,O{��� 	��%�b_s�Γg8���-[�~�v�Km�s��Kı=���I��%�b{�צ�q,Kľ罝&�X�%�}�{:M�_ˊ>(q3�uyܓ�-��Wh�q,K�����M&�X�%�}�{:MİRı/��gI��%�b{���&�X�%����7��`��s�ۛ��i7ı,Oc��4��bX�%����7ı,Ow�٤�K�����O�T~�hT�����M&�X�%��~�1��7�L�9�Mı,K���t��bX�'=�l�n%�bX�����Kı;���I��������?�Q����HawBb�^��n��7D!������m˞��<R�7j�6��̘��c9�n%�bX��}�I��%�b{�צ�q,K��3�]�X�%�}�{:Mı,K�z��!���:�;m3����&q3���zi7ı,N�>��n%�bX������Kı9���I�ؖ%���Ԧ=3�8-�\\��3I��%�bw����q,Kľ���&�X�%��w^�Mı,K���4��bX�'=��Õ�)w.j>�~oq���7s�������7ı,N���M&�X�%��{^�Mı,U�;���I��%�g��?~��;h�������g8���u��Kı=�k�I��%�bw����q,Kľ���&�X�%���>T������T��M\}4l~@q�x4���WUu0�k�r�@
4 �m66b��@>0�O��Q2`��D�U(��8�. mI$#� Ra�!
#�D�@J��	�'c2�2`��
��5��4���Nq(	�����9���z�i�O�"�ڎ\*K��.p.|H�r�m��8jݔ-��  Z�඗���
$$/Y6ض�VP�d�I�U���5���-UK�l����y���A�D5�s:7d���4^�Q�(�uţ���.��K��иop..m$el�ԭ�#]fzV�c�V�kfԼ��T��t��곳��V����.��6&���G��#����jw+���ZG3;;�U�,yӎ뉱���Q�㓬�oj�����=gW3�ї�����"6˚�[YJϝ�����r�@�m��ͱ�����4���V�=.�y皥���ڪ�3�s7f��_n�"�����kp 6�n�yE�īU���٦�5n�/��J��r���i-\ �Mf�e����q5���������tk�`]H��2�n �U�E�u��T�1.��e`��Ύ�l��H#���5/.��kn�,����$V�b�;�'9Y�5�����]S���ݵ'�pa��l�݋���Vc-��m�9&yvΰ��%��G��\��0;��n�� �Y���7g6u탧Rg<���3��.Q�-��v�!���\�FQ1�2�vɗh�2NIm�0�e�T�����/Z�:�;[̑m�Ln�e�v���k ��q�l�l�[E�����3��u�C�T\��R�zۻnf��)�`��RGB�ƒ���8����V�2E�u�i�˲�]J�R���q�Ѫ �٫[@���쬏n"�V�S��,X�M���N��a,� �ק"�8�pbr>�Ň����ۤe%��N&"fVuۋ-���:�dʣ�V@"ږ��Wj�.�l��ݘ�;)�Km=0��H�d����;.��WN�ڑu#�*��R�\�ê��j�z�#-�I�����.��Anm%J�Uv� ���JuT6����Dq�5�e�!�X&�mUw8�V�dGV��v�:��,�9ͷ`�l��6�bLY��7�m��h"�TەAC��C�!�� � QM���9�(���H��N��"��o���f��9�I3��0���n8:����\#Jk��nV^��D�Q�Gg��,Y��¶�'�;p���C��%`�L�I*��&�
�W=Z;2���4� w&��A�vO]$�� $�+���a�ó�3ň�g6��]���3�K+w�g��#�iIc%� �tţxs�6�v�>��<�q�l��6Z�<����	ՌA�薞[�S���{��|������:2rӵ���:�Y쳹���=�v���'Aú�
��J��ʩe���8���/��zi7ı,N�>��n%�bX������	~���%�����I��!�����8?�!z�PE[�w��ŉbw����q,Kľ���&�X�%��w�4��bX�'��zi7,K��9�pc�3lq�2S8�n�q,Kľ���&�X�%��w^�Mı,K���4��bX�'y�z�7�&q3���++u��R���[�_�'�� 1����I��%�b~��_��q,K��9�cI��%��%���_�&q3��_Oz?42�[T	��3I��%�b{�צ�q,K��s�]&�X�%�}�{:Mı,K�{^�Mı,K������g��e�N���/��q��n��cS�=;�r��83sx�?��=_c��>x+�j�������,O{>�t��bX�%����7ı,O��zh?
O�b%�b~��_��q�7��������6V)w.�{�7�ı/��gI�p���P�'�,O~�4��bX�'��צ�q,K��s�]&�6%�bt�a}��1s���ͷ9Γq,K���צ�q,K����M&�X�%��羺Mı,K���t��bX�'�:O8��r�UE�&����
HRB��ޗ�ı;���I��%�b_{�Γq,K���צ�q,K�����r*[mn�i�_�&q3��[�|��%�a��?~��:O�X�%��ߵ�i7ı,O{���n%�bX�����r��`���J�A����wU����yŻtm�|��un�I��d��coN����>�bX�%�����7ı,O��zi7ı,O{���n%�bX��w�8�L�g8����v�0�'H��c9�n%�bX����Kı=�k�I��%�b{�ﮓq,Kľ��s���&q3�f�y���[��L�i7ı,O{���n%�bX��{��K ���;A���D�Dq� 	�
�P�	���Mľ߽�&�X�%��:k�I��%�bx�u)���pK���g4��bY�X��g��Mı,K���t��bX�'��^�Mı,��/{��_��$)!7^�Q�r����1�3��&�X�%�}�{:Mı,K�xצ�q,K����M�g^��9=-NZ�b-PQ�+
J5�0��5�^�*��H�86����ڍ�r������.�)c��o�>���n���;����������}�Q�e��,�,����m�VNc�6�X�S/�2f�i�,��B�"t���w� 7wn��L�j�,��Vg�I�sD�W����XmՀ��2�m�V	%�%ϗ���������@�'H��.�'J� $�R<r��j ����� ��LD	�[��ݹ�j��{�������+�)�wd��nk���Ѧ�uQ`6ݫ�1̀6�l}!����<��j/Z���t��{;�?�{޸��0��Y俤7g��NK-���Ү\�X��U���L������ŀk��`���܅�;h����Q=֯KwvՁ��sa�%\��U�����'�S�(�(�UE��v�(���w����`>�L�%BK��k�(�"�կ����F����M�\�s{u���ݫVtMu�;^�ّ�,z�7E��s�v5�����vq�CDt"ƚ�&�nɫ"���L3�s1:i���f���f
F��n�WEs[b�&��u�י��+�=� "r��?ߔ�'|/(�S�w1��8yl���q�ը�mP�8��Xxv��c�5����]����%�կs�b(n��e�O{�����>���e^HlvG��Vm�"'�9�$񎋵\[��o#d175(k����I�m�:[O�{o��� ��L���������$�l��"��� 	$����I�@6�}��ꮑY��[�~�WLwn�{������p�����X`f�n�	&� �� 	$�~�Ｓ���Qz�Q��WKi�w��XmՀ|�u`6�䳃$CѰ�,]I��Hh��OY���U�4]Xܜ�P�Vr��QS���E?���XͧVn���[�Xi���u�m��ݷ ?n��q.,�92�@ۦX[|�۫:b]V�-�,�ʭ�7v�w��a�qq6{������}��7�-$�؝7t@7�Z �M@���$�?���[9`T�e0wv�K��{��������� �{�	��X�[/ �bv��յ�·p>m/�����-��V��r����:F�In ~�[PM���@I�c�(�6���\��R��t��BP�^Q	(\������U�|�u`4�\N�$������3���n��K�@��	��%��TO!PM*+��g�� �ݾ0�^�����uX�a�Q	$�wwj�;����2���7�~��Or�-���ݷ ?n���`�v��$����*�l���z�vmk-�s��{vA|����n+�<'=N��b�B��ʃ߾����}������7W���֖Nc�6�XͧVZ�S:��E+���m0���>^�8��H�� �ڽp�t�ˉ6|��Z�lT�6��7�ϵ z:���l����۸�G[,��P�-��\��(Q�g�z�{�����>XDB�4DD�]�ۀu�k�4륰�'�j� ��e����`�Vͧj��P�Dca���.��j�J�:�{^�n�ս��-l&�.s�ڟ�~�8�{���=�X�-nLU4UQ�z}�ܰ�Ձ�iڰ:f wWY5;lm�:�+�`�v�6���X9���"!)��9S���%�Q�c���y{�ۦ�������;��o2��\�$��U�<t�3���c����uo���/5�ZH�v��-���v`�X<NՀ�ݫ興S�+�T�(.���vzikR��;l��L/JA�Gp�9�w[X�؜g�A���n��sr`;F�t��f�Ɋ3�r<�N볞�g�Sf��#d��Z:��I;XvvK��c+;��{a������.�8�.ޭ�ݰZٗ����R��όR�N�e��N��a@J�&:��6nt�<e{x�i�öl��S�f�M��⪺.U���*����������Æ�0�z{s�X/PQ��SlA��vל�d6.R�EL�q�X⮌#+e� {{�`|�;V�v��/���XǶ����ȝ#C� ��[� ߷q`wf o{�?�.6u�{�ۮ��dh��)X������6G�(\���U������ ��wU9y ��t�����@�����9�H�vM/wy3%)�\*j�`����Dy(����W@��b�:�ݘ�l�I�"�n��b�K�˧zϫ��Y}���J���z�3;C�����Ӗ�-���9n��]0��� ��v`�ݸWQ��G,��Y)$�f����Ѭ&Q�@� ��� �����`�证Lrn��ƀ;���?wK�s�6w��zG��)]�'K*�5��`�ݸy.7���0w}� ���HkU��X;,���9Į�s�@s�߄� ��=��U��hc�����o۸���� 7�� �[�����I����n-���p������r��P��R\Y���wwrl�,M��]VDԔ���b�?w���=�� t��t���m鹴���- z9�7[��.%��|�����7S��� >�}�I7���Ʌ���c"\03;JL�@�H84`J�Ĭ�pm�P�a&0�H0A�0���R	F1HA�eu��v ֱL`�1�%��2a�� �!1P����0k"PO��R�>;�b@�A�? �`:
)�N��wk�ʂ��qI� ����SΊ};�{�RM��ԓ|:�܍�Kh���-���n,�wq`�;��\o�o��A�_Q�,��f���H�*@y㖀=�����������[0Ba
#"��N��Zg��P���[g�1ۧ��pN�s�h����e_��f������z����K��b�5�!���R2�I6�����u 8��Z��V����#C�[�~�V��;�w�l�< ���|�5jm�J곊W*�R��BQ/���=� ��R!GR���Xf��.U�MTT�\�`}��6����kmX�v�||7�
#m��Gl��U�(g|��sٯ<�ƫ7�dyD�����=#�u˫9�ڼ�3/so�9��<�EH	�*@~���WZ{��Imu�� �ާj�%�(�=��7���u`<A��G,��I(�`�n������6{��}��� պ�G2�!K\�(�Qa舅=t�lq�Xf'j�v�|��$5�𬊧I+���p(P�u��/��u���s�$v�P��E��w��C�T���0\�cC�3kp=��^(���Z��VqE�m��F1!�m�F� pAѓ]p�$��ݏ���5����+=���)8 �ظ}�ca�j��r�
6n��OP� 	˰{1�)x��b3Oi�"dѳulzn:d�6�9F�t�Yڑv��S�2�q�n0S��h��H��@��ՠ��][N�۷YŇc'�.[2D���\n�Wt�L�1fq��2"'��L:��&󙅤0��<Y��nݶW�n�	�uۏ��^����{5��Z�ZYZj��t��ށ����r�`}��?��Q����MZ�uһIR�j�7��0ݝ׀�v��ո�_n㊩h��������9�l�Y�
g���`n:��5}��r�F�r�Gex��w� �+�H	�`��{�;��.��ܨ���'�U`}����D(���O��w� o�ۀo>ٕ�+E �#��\Yѐh��vt�s�nS�i����G<q�������I)U�VKjU�oݺ`�ۦ o����0�u{��/H�W$)kqJL�jI�s=��@XP?@#���Hn=���ڰr�`vN�psD���T�<��qՁ�bv��(��߻�����~�w]�����Q�J�U��(P�\�n�U�����2�`�v�3MZ�uһI�[�o=����5 y���:0���Xgvx3��q��b�T[v+s���8�f��F������w�t�\�炼�W)|[�,�XىגQ	}!��b�.��VKdn�*$n� 7��^�%2mmX�mXfS/ВJd�Z����o$��-�����7��5>�E�P 'j��F�?��\��~�� >�\�7�l��Wh����[�	�`��{9�@n��[��R����U�~�n��B�ǵ�mm���ѐ�s�yÿJ7fv�b�U���ygx^;Glȼ��v�=�:�݋b��̳�ˣ��d�a���~�'ڀ�u '=��� =�a��u]R���[�~ޭş�$����ov��5�ݙ���o��۶*�(���H�߄�@K�1��*@E��x�r�G�EMTXlB�%׿x�'��~Ƥ���Ԃ��RP#j4R#3��`<	 S��Jqs�{s<`�}�[r�S���`9�>XI,͝�|�,�S,��?���\��{W;��f�k��ܓ\L��#n�{ipn�8lqn]�{���_:L���ͽ37s�s��Rs� =�_�ـ}�yv�)iej�Y	V�wU =�_9�t"�*J��idu���$� �ݺ`�w^����I);���,���X����֫�2��� =1�@{� 8�����v����U�b�9f��7����]^׋�x�`LD P� ��$��t������{���I3��lur.r�:F���I�˹.4-[+;;t�g�l�N�荻8�m˻s�F��8Dp�[=�I�w��!��?e�v�j�p�/g�6���N.�`urmn��W����J*r��ܻ�q����[s쁵��)1�vd�r$�$��h'e�i
�=R�$�p �a�9˕�b���NҼ�2� �Bk1H![�:}����w��������}ZA����<�u�#V�Ż�xܯ]h��㇀�3��[M��z�l�j�C����o��ϕ =����R�H�*�U#���U�~�n���ϟ�� ��{߻��Wۮ��2�*$ot@z㘀�2*@>qR��h��(�m�K+�Kf� ���X����$���L�=�=	]�����0ͤ� <���b�ɋ ���<qV�q���":랂x9�mَqb�7��pA��z�	��T �x.��M3r�Lͤ�� =q�@{�}_����,���C�W�\etr�罘�<����"�� =���K��q:F�;n��7�n���$��o� ���;���Y�4��J�����Xi`1ՃԹ��~X�w����ܵ�!eX~�� #sP��� >��,��7bғ����!s�F�`0�j��h�#����aۣ�ڰ[�����D��B����X�K�`>�k��2�2wQ��Q�ۜ�W#���6�w���)� �_�"S&i���8UQUR��Jy<�`nnڰ>̦Y���� ��aRE���D���)����˟��I7��hԒt�Sz�NҪ[I*�?w�L ��n��VP�Т%�?{��r=�<^�W���ͽ/4@���qRt���ۦ��f7m�n[ʜn��x���ҵ�8�;�+�<n^P�nҜn�5��i�Q��̭�ˢ���s��:EH7���v�3wTh���М�� }n����B\�����}V{��`�����֤��`�;� #sP��� 	]%��n�z��9<�Qa�B�3��X�;j�}}ѩ?(�Ϊ��t#=��jI�I�}����[k��n�z��n��7�`��p� ��d��Q5j��v�ql<vWu=ury�ّ<�y�	uB:� ���$-���-N9V�n��7�`�lG�P���3�>�`[�3�T����ݣLͤ�@��GqRt�XɟvkU�R2�]� o{� ��Vj�J��ݵ`nmi`}ܦW+evH�Q��ۀ~޽ŀo۸��n�����;�Q��k%U�I]�@N�Rt� �����ԅ*�8c p�	ց��D��SQ
@@����)PC!B0V,T_�'Ā�b�_�)A,H����r�S���}99��N�!i��c	�� ȫL�~��A�M;��M��G!Q�Vk��� 1�h��1 Aa�2|�_(���ģ[�K�������m�e��m   ��ぶ�e��dQ! K�d[om;M�Z�-�M&ݺ� 1�i�9vڬt���dٱ6	g��[;���ԛ,ez���tp<)We��s��V�P+�8:�תN#�8f]���uւ�X�Y��d�)<�MT�=���X���鬖Ӟ˻V��u2��T��kg�(Fv#ub�f'm�nV�;���Hq/n۫G>8^X+s�h����ɵ'Z��$�^6�cp�X���E���qb�g]dAD�铤0ʣًhމ��;t�dz��e��U��P t������F۬;���	�TZ�v񹤞�mm m�գuY(�Z��m��:+�������Cpl�������s�{�8�oh�-��=&��V��:�dX�9�kol/:cv6F\��E�[Ν��u�1�]�MR���m�b`6џ���Ƌ(��v�U ���[���նd69g�lƩFpb�i�7`X�]��Q�d�'�5���kX^
V���.��R0Gm�Tn�P����Y+��[Gs�d�v��e��{t<tC��]d0��c2�}��Yγ���R�%���r�JU��uN�ӷQ�3�d�dZ��5WN���8�Y����F�tk�!CNE[�R;�uJ��\����kIm݋���a3n�9�-�Y�:�V'E��^�>d�.�%y���I-���L�U�]����n�m�q�K��A��Uڕh9��[Mͤ�*��kc�Ym�@Bʴl3}���~ü�ڂ rN��U�VY'�+km�V�/	�e����l�%BiUV������u�ʞ������X�\P� �s9��na��T�O[Wh蓌1d� ��f�@uQ��:��:�P�n�[���\��q;�\�FPN
RZ�ڠ\�L����}Q`���C�[u'`�X�Ί�h
��+��YF�ݙO;��<Y:�LF�Yb�m�)N�� �dR�M�)�S�r	� ���%D"�L�h)�2+�B�@P���	�2��UC;1N�ȖE[1�!lۄ���\vƴn٬<�ʷ��{Fj�&y�E���tZv]k�~�~ݷkn��(��g����fA�5�#rfۇN��vͶ��s�3�/�wf�u�g�rGF�֎q.�%���]̑�5T�r��z܎�t<�p��8�Z��I7����S��c�VvN 7[M�M+:^�Ŋ�'�7Lۗ�.rfیg* pCyݤ����K�k��j7c��m�{gԣWvwX�0ą�&w&u���|�������z�>�t�9�UK ��x������V�v�Wۮ�-���hG%� o{�?�$��;�vՁ��j�o��J���3Q��d,ds���vۀw���b�7��VyD$���֖��Xa�4�IUG9Q\�S��+��VyL�����BO�y��������V�:IV �;V�(�{��ݝ����C^���������ѹ7���m;<�'p��k��n]ӝe�4�:�X��'X�ٷ��� �M@zK��ȩ#�`��ҩ[V�+QA�[�~�{�4�N(�ʣ�SV{���I9�{F�����...6|��Ik-U�I]�@}>�RG �����)�q�j���k���`yqr{���z���j�xݫ k��ʪ��J�C.�6�rjt"�r*@N�L �l]B�Qb�*�pv�����/n����n�u+�����h���q[F׮��r>���L�*����v����G�; �����;����m$���BU�o[�~Q2n���5�Հ��j�d�;#�;k���U�{��X�ݸw�:+3U�Ҫ\2�(QpHհB�P�{uGmX�ڰ:��p�9�`��<+��5(��^��=��X~=j��EH	T��=��݆�[��E�ʫ��Ձ�J5���u� x�`l{����ڍ�·�ɱ�6�z퇎��v��)v-��NH쁿�����J��T�O(�_�vՀ�;V �7�7���qZ�c$�E!mX�;W�Q2�j���mX�`u����S�#rU��ۀo�n,?�~�{��ذ�]i�B�G9m�7yUa�P��3~V��Vx�X	.��")���9�S@��7���?t�=��m���BU�G"��*@ɨ	Њ��3�f`�����5 �][�*�[u �A{s�q�����=x�����5�e��$qR �M@N�T��EH���&�>�W*����qs���b�=��,w��?�g���[UY��$����mX�g�L�nڰ{�w�ujv2YUhNRՀowq`�� G&�'2*@Jn+��·%�)j�7�`��}��wOb�7����O���6j�T$	l������Z���i&ȤCcf�'3��ۻ�&�#Z7��2rj����o��~듪X8rOm�GS�Iq�m�T�c`yK����:j@vٖ�]ګv�`�8��T��-��rl��^�	��4o���_nv}JMnkum�:,K@si\����(m!B��p/1�U����cA�v#��Ď8���q���@Q��ۮ������q��������Yw=�U]b���N��<e����b��cml�
A�c&���h��,Xj�\]r-o�����X�;V��B���,?�DOZ;�29�mq�-�=�=�?�$����`﯌ ����N�fH�imj�Y�@G"��@;�bs"��Wu���Z�U�o�t�:�w��Շ�%���{��r=�s��T�6̭��ͤ�& '2*@9"���� ވ�,pF��KcM��n*�z�v���vm֑0[]������Y���t��F��U�V�mљy���ȩ 䊐�T���ـw�ujl�[+��')j�9��F����UC��5��߷�RO_��L~鸰�{��
�[H[RG �1:R� 	]5��]�S��ܕ`y.=�������*@H�����L.��ݽ���@N�T�rEH	T�w$��n��핅p�9#j�	EU#�uٰ�\�s��b
:N�mv�y����n���)��MT�9J��ݫ��VKo�^J;���ذ|��ۊ�ҨJ�I*�7튐䘀�ȩ 䊐g;�̛R��8�yS�VKo��՗�����2*X�F(�͢%Ar�(a�����ѩ'��tjI�};��ک؊V���.?wO~X�� 'H� �I��:�wF����nQW�n�� 'H� �I�	�7 ~ޢU��*����1��w^/E�M���;��q�/mm:�\F�eC��ݽ7�Յ��	j���b�:�v`�Mŀwwq`��]��:��IV �I�	̊�H�#��t�r8EJ�uGl�7�7��Ň�9���{����;��6d��T�U�'R�1�j�o�%��
��AYIH�Q )�=���, ���ۊ�ҨJ�I*�7{����,�;V6�X�J2�xO9���vg�5�Y�fw���<��c[n��ۓ�nKb(V9\�Iqe2�$�Z�*�e_��{���v��ڰ>]�7-S�
�9f�i����,w�� ��ـ}�:�6�m���')T�mڰ�jͅ.ww��k �7��+aE%����`��XKo���D���X��jfyEp6ͭ����@;�bt"��*@n�q`�����z�m�-9%�BFa��]kۗ��3v��q;Dm�s�w�n��D��VLu9�F��=��2(��[s���d$6bUp.�nB�
ٹOfx�S�R�F�� �<�I8���ӐSf2�v��8�m��q��kYtt��(�3���v�1�ڒ�G�\�J���q�Y�x��#-�����ݯ���c9��I��E�r�&��{,u &s�I�d�g8�uTS(�T3��sg�;cX�gn���*�M�خ�&�P��۠L�j�;X僋r���B�:�QpVx�C�*@9"��*@;�b�>l�r�h����`��Y�q$��nڰ��,�;W�"!L�4�fx�v�B�)%X��ŀu���7�7��ŀ|Ϻ�m`"�U���D)|��X�m�v�x�X.�5�S*v!UBG,�;��� ���I=��|׶���,	S�r���*��z�{pRY4�q�Oe�&Ů��؝��$���յ�(�c���C�2)�������9�T��n���S�^V��\c6���&���;�X� ��Ċ��E"@�".�Z��,�Ձ��W�P�$�����6ԥ�S��Gi�y�L��n,� =�Ν��e�e�홷����GQR� =�ܓ���T��v�ԫ ����=�s�Q���%��؀� '���{�^�m�)�u���y3���"�k����2�ڠ�qZ裭�U�R:���`��Lܓ���*@u��̛��[W����w$�n��*@{��˜�>]��-Ec�
�9f�{}�RNw�ѩ���Bf�,����܋$b@�?��N����u��*8�c��U0�(���a F""�"��
@�1݅�BG���!B����!IBe)bBJ�0�� D��b-���Q�� d�k�p	� d��R,F$B�S	�11�X@�����yA��;�C�5��8�J����-���p!$ F#�}�c.!�f�J�l��E��T�@"A�sO�`ē%��R�FFF���1d"�X�H��L��ɘ|9  x)D�!�����a��! G�H���� 0+������P:�ݘ�kkShv�q5%v���w�`w9�6Ko���;�:�nڅ`�嬄��`��� �\K�=���$���*@u���ڼ�/{N���N̶N�����m��-�ѹ:�&^ݬ7�S����S��k����32]��v�	}!����iʝ��E�Zmf���n�w #�RݒZ x�^�B�$��W��rf��)�EMT��+��Z�>�o� �3v��ՠ��Uc��IV��v`���3v�>��%��@����� p��k����q������qR��*�`�Т��^�����>ծ���NX�6ݶD�i'9ɳD׵���ì�����<���3p���k���r��в�u ��r*@z������7{[Z�C�8㉩j�7j�Сs�N�ܰo�Va���s�\�>�e�
�Y-� ���b �M@68������Ͳ��N���ف������7M�,zݫ�	/B\��{�j�S�G+�2*�ͼ���@68����& ���p�.ħ����R�ۢu��[��k��on,t{�+i�lt���lg�g;��,cJ�����6���'
�EY�DS�P5^5�wڲGd#	1s9�&k�[5��i�U��:n�0�2�f�Y�`�Z�s��ۀ!�r��m���h���8�,@�Q�cY�6�
�B2��f�3m���1δ��gG&yӂgGj]�]ˑ���٬�U}����?	�~�r*&�R�l���!�/��6O6�7jL�y�>���Ƭ�s�HZʜ���IW�?���,�������;ӻ� ;�Z*ݥN����`�ɋ�]���!>T���H���XB*��ـ���>�������~��,���>��BZ�em��y���N*@F��Ɉ?�?������m��&�VՀo{��ϻ1 N�P��H���zna�\Ok\���V���on�p�v�X� dG`����|yL��mB�rV��~����5ΜT���H	��U�n�y2c��5$���θ��� =ʪr"!*IBK˴_W~�`n�ڰ>�o��]i�#�6+U�7e��]�X��R���:M@��L��sj�m鵙����H[��5ΜT�;�Z*�V�����`�wf��ݯ�ƞڰc�`~I�l��(�UH.uy6�P�v�n�m��L�'u۬�Ɠ�γ�&�J'�ў���Ͷ��~��t�n*@wc���{7k/L��/7P�R7 =nL��v��l��H��c��`�N+j�5��`w��6UD!	BD@�!$�	d(�(,yn��7j���wUHT�Qy�f��H�r��5� 7��Xw�aS�C��UP�W����<�{����}j��y�l0s;����\�+m#F�����������spܽ�����p^ΌV�M��Oi�D&��R*@F�v9ht��:�9��YT��R�*�7��X�N���v��[���6�^n�Q]RR�i �O� N�P�R7 ;�]��u�+"��%x�n���wF����s�:�P��ʋ(��6��Sj9�w�'�s��$�s���u�m�p�-�X��{����< ����G���l�v[pn�t�����p���ƻui6{�Kn�3Ό�HlaU�6�,NA��VՀ�ۀ}�� �����w��7-�UB�Z�+.��� 䚀�T��H�.�����
��]UBY^ o��~�n����{�ŀw�|���֝Ҷ���]n�p�-�X��,�u�y�{޸է���,�K�)T�`�����s`�V�Mڰ�����!.-G��O����TP�������G��_=�B=ֱ�L��Z�o�wb�5�E���8O={urb�IZl��J�t+��n���^[-�nӻv�g196�t�7K!h�cYX��;R�f��Ky�M�:Aw^j=�Dzwp'��oT��Ş,��C��3�k-��aR�xlT���KN�zݹ�x؎8�s�d�͇� 'Kb�&c1N,��n�t
�+I$�s�q/.bY���}2�e�nA�'�����VP���p-��&�m=��e�\�w2**:�DuIc�h�� �ݶ�M��%�����'�5(
���u��hI5� �R�y�&��}2�6V۬�n[�}��b�1�j�%	L�q���ڰ:���Դ�r4�-Xwwߧu�w�p�i����[P�(���j�3��6�����j�ǎՁ���������ʪ�;5��Ԝv�쉬k��7S�nї�I4ld�ܚ���\�Nî5AÓTt}�U��X�X۵�_�ov��>gy��Cdr�a-����|Ȱc �8�T�!	%P�HK�7NՀ�� �u`.�͍��N^YK	V��� ��L��ɻ�VsM�`�0�*&�Q��30��@>{�M@z:���ŀ}�]��u�+-CU�`ۻpGQR� =��]/
&�-gk��F�;��r��ێC�c�lүb����>{?Ph�U����J�R� =� �&�:d̩VӒ��4ӵZ��wߧu�ۻp�ո���-�Vr�B�j�3��6��Y�%؈���(��)����X��ŀ}�ܪ'
���hB\�@$���� ܊�*����>f�4�#��� ��[� �v*@>�- t�P����sn�0�>�ͺ���g���ܛ��cEӻb���x�{V�ù��CT��ݮT��uJ���b@>qR �&�=EH�P/+K�H��YV߻������}�\�j�,��ŀ}�]��u�
�CUڰ���>x��6)��mXi`f7b�hW#t�R�m��9Ē_�$��{�����XܦXT$�duDD5	Ff�ˀwgdZ�NJ' �N�j�;� =� �&�=EH��y�L���i�al�q��n[,�뷃��;��m�����\ݖ�r�e�Wn�a`uU�`��2�:۫���y%	.�7w֬����'
���Bʰ����\�&N�[j�m�;���)�$keN�&�,��c���j�,����;�w ~�ۀt�lvRT�喸ԫ��$���+��V�n�==ַ�`|�*;i��j�;�w|�J9�ݮ��JT{ܵ`~I$�DDG�I ���UUW�� �� Uʪ���T_� *��Q�
��*"�*��@��@��@b*� *T��@V*� *��E���@��A *"",��H�� *����D�`*H
�A��EF� �X
�@��B� *���", *"* * *","�H
�P
�B��"�P`* H
�X�,DX
�H
�Pb��� `*",H��H
�� b*��@� *F(���E`��"� ��P��@�"� *P� b*�EU
",U��DPb��U *A�"��,��A",@��Db��`��* �",�A��*��UPU� "�� U� ��ª��� _� ��� EW���*��T_�UAU�UAU���
�2���y�+u������y�?����	�| � �  ��    QL� R�4 P4   h�   j*�� � (�*��
�$�E�"Q@   E���J��  ^�� R���(�ۡݾ�C�#�x M� }��z�� 0�t��_p �Gѐ�>�� zs�ӡ�$2h>���  P
( ���I��ئ�ɧ�� pdi7wA�EY�.�ܓ6�c������2�8�x-Y���MG=�{�^��Y�`�nFW� >�� � ( a�
{���9�.�n���w�Y �q+�Omyj�w�4�A{���NY}���ri���W� qԳo�W-Ef����E� i�L�I�^����sd���  UP  VwpP^�NMw;�7�ѐ�� ���vt .ƀS iJw �f�FM�A͔���z ��d �Ҋ�J&���P�:� �)FM(g�}�|P �  P�����U���d2.����YSv���ۙ�������Ñ�� 0�,�>�u�pH�4thi���x��w���o`�f�� @   )@ i4�IM2��0�42dLh4I)JFMdѡ�24ɓ&0�~=U*4�D   2   تT��T�L	���0��A���&$�)G�0 &F   ���D�@O�G�O꟥7�h�=4ѩ�:���|��az<1���	i��w(�����7i������<AEC�A�����#��o�������X�4��џ� �qS�S�H �����a��7��>�?G\���o�     �   �@j��@9� � � @( �6p[� � � ��` 4    � � � h :Q��DCp�V�IC� O���@� �@W� � 	`�A� �~���~�
?EP� � T� @�*��>��� � "H ��U~�
@�@�*�� � ��@����S� �� � �E>�� �}_���T~�� 誉� � � ��A� �>��y� !�@O��߾����z>,6��C�?���<y�~���W�~�f��	���7p�3]��1��27�<9�WNc�Æ�a�1��P��n�m4̤�I���#�������s���^$�a~�������\yL�p��bjP�'fë�Jt�g_����˗1�L0����	f��a�f+��S��d}�:bD����7*�+�6a���3��I�Is�s;4#��C ק�������ޗ��ap�3�9�5���A��H�S�#�p;�w�.�)
���c�I�g]�i/]������Y��с\fy$�:'�a;ɦ�B����SH��8ˆ�/Olja���7q�$aь+�p�2c���M9�eӔ�(E�*B$H��5�f�.p.�>�'����&�����;�3����!R F%eλ�e�w��O v0�
0��jc
����{<�ΐ�j=�<I��q!X�L $4��Y�KJ��!#�ÀER��+�>q�tF!��.�0iS ���)����`XGLYa��K��=#7��c"�&��֠�����۝d�%��(D��޻��'�"4�:��	;���)H�plm��+2��D�d:��9��`�@
�d�� ��,��;�w��P�B�m�/RJ��!ü1(0�����ẅ́.o%4��#@�'Dtt>u	O9�<�`ŋ��;\�T�6�'A3B54Ir�F���=9<<2�|���� N�[��8�wd�y9��<�7��� �X�%!��%���Sx�]�f!��R�5�J���a��P"`�:�@AH�X�`�`E�$z{_$���!�t�J�CB'����0u�!�2����,j�@��=1��m��5$��L�腉��'�}1�))��=��<��3��!Θf����{ᐮ"b��z{9��7��`.)�Hu	+�(�(Ah�
c�a��4�����x$��V��vq#z"bt�G���u�{H&���% ��4!Vr�;��Y��\!�A�&B��d�÷��#���ă@���������H�B�	 �oD=�����А�Ā`�'�{r7^3���aف÷_==@ �058�'aǌc�`B��p�or�U0N��	�=\яC���`@)��p4u�hL�c�����+�1�n	��d4�$+*�V��$"CB"�0�i�gsw@����]�7�{;�3n��:�e�LeaIp��Ox����y���󸬧����S[���[y��=��w��e�!�XHU%#	������p�DT�;<�ޢ$;$E���}�}�2.��Z��e��*ԤkNڬ�.���!�(�,Z��@�0Y\ӓ���i��Ib@�T��D;���$�A��x1�]h8���@�h������2=eJ0 �� ��$bD� �$���$ C�nL�3,{�t@;��m��������X��
���ÏA
�.@��<"�0!L����H��Tq�5�Ŋ4"� X�2E V�2%*S���C j���q�=G��D�(0���BN�N���cw�2b�0����Gc��B�vp������C��<`�xw�u�1η��i�B�-m��jP�-j��
QũB�*���s�S5b�#[��'׀��ng|';�v���q�lSM�'�J��i/��T�ʹ�5۫!��{g\�č�;�Wt$B0)�k��̝ap��<��AOD���= �"D��)J¤b��āB$	H�!B �si*@�(J2丌��.�HZB�+(K�桧 ;N�t
']����p �������"F��"�,vHV0B,Q�B"*$��v�%����(�����ܻ㤗�_z�`A�#ƞ�����
a�fn��=Ig,'&E�HtD8��Ӫ:P�+��5�} Lӗ��L\
i��L\Ivq�r&n��p`�a6k�A j`QcR��xK�l�͙�z���F�!+
0�i$))�
!��(J°`�.�]������Y<�{Fl=���\%��0����A�;�P�aB�0�	gf鼖p���|Ђ�������Nl�P}3���M��x�IsH�pԔa �;�d�LQ�S��͹� ��c�T�]z룙�Θ� �\t����C��t�"U�ނu×$��bH��aP�����0�xۥ���L	LcRx��U����D������I��	
��+/�Z�2)����@�D`�8B��Hu��!�+���E!D�Jd�!���2摤`ᦛ.n�4�%0ݐ!F5ӓyx	���$F	T�"Rp��B�]$.����+A����d�C�E ��Ǿ�S4V R0CÄ�X������@��D�%XS���X	�CB0�5�S���4`A��L%0���"�1�-3��0`h�h*�k�qk��8n�����tǣ"jv�m�k����$�]� :�u.W�5��78�^���	sMcLq�B��5%0�h�s�y{�מy'����%��P��	TÑ��u�{�++� J��+���vwN��9�Jd$�a�:��a�2�(c
d�,jB��b����bF�� `������HIYp���>c�vu<	��@$ux�v�p��˧1��Ln�Cw��tq|a��(J��tۺ�� @�E���^�d�xI�k�{V�˜i��� b�E�Ei߭&rtޭ�V^�	�e�SKF1#���ā
°!�v�$*i�)�Y����#X0
w�4�o#�)�^����P8/L�CKK
X[��zb�5�4
 F�1u"�LCD�*��H5�py�ZK��#�*����ffݗa)-�d	��5,\�<�NN�˦^�3%��^�z��ӭ{s��ݏ^z�V��י�$���k���;N����A[��c��2����O���v֭�m^^^p���z�ex����*R���r���&��]�^^��ߑ�߇���   @              �            �   �M�  6� -�  � �m�  6�  6� �  ��         �=                                                                         BD��E���� ע�x/Z�u\���-��5U2���ʩwE `"Kh6زZk�[%e�R�3��;;5v����غZ��U�亰c[k�,Č=�ߍ}���8�eV8B���5��/ce�'NT��]/dYT�L~>w|i�nȵʗ�U��l�, Xa����ۉ�/#\ڳl(��kx\��e���%�#!%���V���V�-�!�C�`�H����[r�!`�ӯN�����[�l(�m��H�Հ   � �f�lo;���Le��b��-��y�6L���BAT�.�e��M�]�$8v�cU"��m�����A����;R�\ۀ�k�B�m[[e��.��m� mgJ��5k�� H׵�i9��mp ڶ���|�H�ź�MV�k�����$��o6]l�      �J�o-��$ -@��#l������ � �}��6���UT�T5�!0J�#�z�&�I��6��,��\k��$m�l[�m� l�H���s m&��]��$�m�m��zh imh�`�mm,2�` �&�[@ [v״ݬ�d�g$���m���@ mp$  hHm�:mr�ڪM�	I��	�ā�F�u��A�� H-�����mm�  ��o���6�ޠm�B:FX��v휬�UU-�m�.��͠��l�h�pm���	$�i��(6�&�   H��Im��qmH6��U�� ��8  �t�V�Ę 볶�m � l [A�l�kYλm� �� BF6��[[ltm��aB��-UԫTe��S��I����8pm��k[�n���6��lHmp���A�fݩs;�@�R�@T���Q�Ŵ ��,���Êڸ5�2@]6[Kk��� ŷe2��{x��Y�UZ��@KE����!��2�m�9.̭P�&y@���j�h �2ö;[�s�۲����Z��]@u&nHmչ�N�   �T���,� 6�ioi�m�uр ���qt���T�.m��v]��nl�qW8-�v2�%���)�n���mr����i�enIW�:
 U�[����X6������*�����
9S# "��SfJ $w$m�l��m :8    �` %M�^�-�����U*Իv�J�^���f۴��`-�P;Y�V���Z�]W@ r�)"A�Nѵ�Ż��	�դ�ٷʖPV���1��
L�*��8&�/]���[m�h)K^[�l�-�&� �mC��m$x��)M)vH[@�mm6؜���%q��5����U�x�աm�e�� �kև   s� m��J 
��rt�n��w��gm�m�  h ��I� � -�8���]r�H�m���H彯�N�p��m���j�A�a��m�+�UHMEs\����ɲɷj�V]�  �` 6�u�&�9�4��er��Wm����Ȯ+���Ʊ96��4l�`*�
X   	4�ݚ��H��}ޅ�I��b@H���M�� u� �� ��p�`'�M�-$�p�d�� h�hH	7m��k֭��4�m:dѢ�� Hm�     �J�-�d�h[v����m�l�X -�^�h��ۀ  ��k%�� ]6� �"Y(-�m�ݷ ڶ��Tɵ@mU]U!n-��A�i ӎ$ [N I�`�im�	ޠ:B�8t�)�s��7-�N@x�3פ[m��{����$������"M��]�,���m��Cl�� [H0���hIg�6�[zŠ��I}=��zu�`�l�m,�J�ҭU�J� ��Ub�	 qm[C�V�ݳ* l�TQnP/KUZ  �(�mͮf�UT K�-��`ۊ�m���q?T��=]U�=��-bZ��yU]��6j�j �[t��N�@�-��t�\�`�l 	 [W�k�m�$H�ʴ��*���9�UU*T�k��e��UU��l��@J�r*�WH����� �Q�.989�ڀt���uy�@�;�1���elݪ��9���\m����[V��l����Xn���[Pa';YT�@�	2�R�l�sQOY���)`s�f��N�������j�y(�WM��%�i �����@ ��ﾸ�������n�Q�dm�(   շ� �-�� ��f�6��`�(�vN� ඖ�X`q' y ,ky�h�Ŵm� �   �@���h    @  6݁mk l @ m�D$kh��i)\6�9!���m����:[@	��k�  ��I��� �ڐ� k�մ[Cm� �i ��    �oQ�J-���~���[C��v[�  $hm� �	�'`p�� �XI��l  	�u�0��&Gf�L   H $    p;n�@     m�I�8� � ۷n�I� �  � �[d�m�ޠ�l6� �  �  �        �H8  ��l  mp-���ޭ��ϯ$�]=ڶ��Nv#%[U��
�bݴ��@  	H� �`   rZcm�Γ��D[a��J��@V��iP*��kh:A �[oZ�Hl��c�nM��m�kYÆ�L�m����f����&�䍧d+kj�cյ�1���v��VW5�6��m  !�v6��m�k�  [���@  �� �c��$ͪN�T��2�U@V;	�ej�H8� l�   [m��JvFd�d�x����s�.���UX�_k�ԫom� ��� I�I����`.�	�p 7k���\�ۂOnݒ 
I�m$ '[jU�����ثvvVU-��l�cr�J��[N�b��vN66)T����V���2@�֛lu	bݛl ����RۻlKi��m[  $��V�n�-�uPQt@�U(
�
kmKֶ�z��e�O�l�dv�@����P�2��7D6�"���p�� 6�n[@   ��-��"Zcm�� msm&8 hm�Y{  �`  <���u�t�mwT�m�  u�H����Z  Hl����/6C��[Ӆ�2U� �d��cgC��\�T�s(Rs���,�h;�sʘ+/RѶ3�)��*��� 8�r� M�VJI������"�R؛Y�{��?o��<�;�8{�n��UA����#��Eg���-,�(�2B!"H�KK	$$d�@�l�,���K�$I,�a���� XV������R R��))J4a�
?���$$IB�!B� B�!B�!  �@                     �I$�I$�B@I	?:�(����!�������W�P=T�"�
,D��X��� �` c��8�
<F��Ҩ��Pb�b�c��y��ΐ5Q���uP<�OA|�uy�(�"<=<P
P�zG��@< SD����D� x j �'���QъUbON��P���&T;<�Q=��Zx8���N�4/J*l�ǡ����#�8�,(�C��G�T)��؀!�@./�= �C���S�T��E�}A���/g �0��<Ȩ��8�Z2��^���@��z�� �. A`���瀁Eă�z��`Q�g����O; 8��SЂ�w_T��7P �   �        �                              $�I'��� AD�� ���������UT� lqu3
&P��R���`��P-D��R��� �T"��O{��\��tN8ǖ]�߂y�Ye�k���y�ώ��ߧ�    	 -�E�h���	 �`-���             IZ�#j͛mkeŎ^�۩٥�Z=vϮz�H�-��rv`8+��%LF��mص��v�%�T�:-���mn0��ێ�iT��@������;vq/2���NKcj(mh�^-�]5l�iOb�6+��j��jP�RsT�� �12U�M]4�-�dƛ6�� ����S<T��bU8[b���gR�%�Ӹ�v�:�4q#��ŻN���n�8N��;"�v�p�j�:c�z.)4 ���v����z6�%/u�"͐�Z�e�@T(��]���Z�ֱ��2�H�ɳ@N��oH^��t��N`�U\��"pH:9�y2ZA
碇�r�,�6x;moq�ӑ��5���5��&V]��A�W&:W��H K%�^��IwR�2�C�Q��s���
ڝgv���%e[�؍������d\�W��h����p�#����FҲ���7n���/\���+m�����z��]Z�Rc�Li�����cN����X��G#^��I&�m-�؂��:�[U!+U[ud�Gm��>g#R�!n�-�r�u����)эK�m<�MT�V�KP�����'j�e� b��S5�5��dt��OLuk�"4����غ�0˷h���Cg蕕1#l����fݷ8�QS��c�M֢��]��;��6�n��n��.܄1)Q��8X<�q�^8�b��UTL,�Dlw@�J8
��6�鱉�	�����/M�\Ͳ�ɻ��ftsT<S���z P�xt��	�"�!��@t�<P <A��=�n�a����k  :��n�㤳�s:��'��Y�IF M�����m�k6.kK�NtW�j۵���F�MN"v}ؤD��B;����y;pt6�9�J�݊.�[���v���3��#)�3�[[�,����rGGG玸��M�������������{���m}�_
����G�p��m�;`�*����<)�3�ks�sٯƷ5��g��D_o�f�;R.[�����(�5����熻��^��h8�N�����r�ᬼ�3-�	��3p�^l�xB9y�]�5;�l�JTe��sv��_VD��Ք���N$Q�B!��ǲ�h9�8��7Ne4(�Iu��z�: �&:3������ma���'�܀f^�R!��npw�J='I��#�(xve��:��7%v��v��&L���C\��9��^ �{�w��I�`Q�m@K��l��-a��{곑��q$d0� ���yoN����@9�Z�AQZ	��]!���c�����u�]�[u�:��5�L��^ʢpw�����܀v�`̶p&�8�Yʼ֫��.��Uq�*��:�jH��|��ovtU0+B�b��i���:l��FDJ(�-�;{�r�����ܔ3w�Ӂ����-5;y;� ���g�� Tr/��Ȋ<Q�� �4��{V�\Q���I�ȊP��0�d�$�P�s};� ��`塆��oqFڅ��%�޽5�݃�V������9$(�an����Xjv����ƫ��K�T�BM��}��ߚs�s�~dR`�1�t4P[�v���j �1�r�ҹx��ov��^�*�gm/-���t�0��i�vQ�XU;u����Ӻŵ��}�O[�7}���f$���zU�[�_V����tG	f$�G ���}Xjv�^�7q=���������<��r� ��9Գ�s0Iʼ֫��.��Uq�;�oqFڍ7!%������;�K�w��"�
�J���v��DD�*!���&J�J� :@HA	J0Z��D����L`�*Uصn�S��:��i��v�  m�U��:!l�e�]{:��9zY4��ap;@L���T��V�����&�� u�#��ɮ�월� �3wce���:�Y�qз:���u�k�m�+d�ŵsf���Wڭ�v��0řԫ;�i�z�r�����ֹ�Ol�1����p���X�)�v�]����l\/��p���q	%�Xq3��!FC�����+[)gG)- ɥ3UR�SSUU��H�5�̓��]�`�bgd����5�̓�̀v�`�5˱a�*Sp�|�4��{�^{�r��������E' -�;{�tv������@8]���ۯcA�lN� 9Z$�ԻU�vn��E
���	Q��n�j�qi���;��
#/ރ��鈘b���C\���P�T���ID�7 �5}6�$mrDK������;Ն���z����$(�arU�
K=�;�MK�A��%��/IRE��'z-5�U�����`/�`���'�1�.2
�������!������.�V�̍����Kp�Z. �2 �[��݃;�vų��M��O�/^�U Fg�qi�w�:ߑ�%'%���9kz8(dK$��m���a���ʜkMK����"�v�Y��$JANEs3D�xj�uA}Xj����)�CJ�(H�T`!���l��f�yZ��§5$R�ɍ9"%����vZ�R�`�VK�Ԓd05 {���֚�g����x��T�B#��8/�� �᫽�2�e��Cp��f�g]w�G�����T����x�Sp�w�E@�n0Y.pwq���9Ն����`��`*:)$&2�	����&Ǒ+<ٸ��QX��#�8#��	N1��7 �V�ۃzm�n�֢a���ʇ����U ,UT	��=�;��:Fg��[��"R@�qCY��s/ ��s�_M��c&4��wv��z�����XK��$(�!�8f���j�o8;��w{�}�>��o^G�-� �^
����	�f����lN�:�[֤����
M­�NLh\&M1cWv���Y�v�>��d�nF��8��k;m�,�h�]�V�L�mQ���g�3��v��tm��5�3OZ.����ɵ��_=���(�v������2%r�"��n�n�����{��p7�P�S�6�:�=\�	�oVƧup:]�y���f��c�o��&]�j�1����]���\�c.�܃�y �܃�Xk�;gQP$ی�K���f���W{p�7�`bS����f���W{pso ����a�����Zk� ���l3�zp�@�h��T[i���n{uV�]l��m�<����\�����-3�<��܃��fno�ј�kp�ͅ�cNH���}��C� H*B@�$"o� Bf���Zj^^pf�%�jI
2܊�o%����7 �,�[�'4�#F(crN��Wypsm���3��2�p!��k3rb�U��z�רUU��߱����`�_;=q��؛n�0��8�v�7c�;P�!	���&�i��E�{���;Ն�������)�#p���(P�n֚���9�� �{��R8.�q��tg�Z�����8�s�]�����_sP�@����B �����̀f��������*0$�I@X�W��A�b@�� 3P�\(jv`�p��h�i$h q��0#�@��a��dc���1�B,�L3���d�@�X D����F t�JF���!�-�WC�$p(�S��k*�;�t�ꒄ�5Z�Ay�����#$ F+����Q����&%Uj����� �⽟�� �@C� E��D���X�?���w����+t�\JHn(G��}�;��ϲP
����߽dƜ�3�������㖴�g�A�P  }�'�!NA)ƣ"��9&�얻=@zV���+�2J���D��H��lՉ|��d����撤h�jE8;�uU����y ���>��􉦓�9e��7�z�솯>�;��]�E�rF�.qkaJ��e-rF��t�$\D%)��(T
���Y�rA���DC�)8��V�o�{�3_�^}�v���K!F� �`�Ry��6��3��_�W��X���.�8.���t<��j�E��]�;����a[���@ӑC[��|��w�-f*홺ɐs�P�׌��K7��\`���A~XN��"��8�Z�]��?v�����}�!�����t����k��A�#7���$�>S�$1!5��  Nk�Gl�D�v��=zsb|C�<�b��(�����=��@���n��0Q�6'�$���7ں¦2l������͔{�Ͷq���Z�9��8��s�s������>����9��/&똵!X�g��%K��A�Z����[��ה�窊�\u3��w�����[�vƞ�'s�ہ3��v�f�v�b���q'+�͘�P�'�֜�߯��?����3~�9kCw�2�q�d�K��Ҽ��,�Ӎs���J���Ji�Jq���a�����3F�p�l8��9����o.^��r��	��$؊�܃�� �܂���ެ^G��pٵ�(���à�f�]k��j���J�f�y�9��#m(Ӓ*q�^����<{�O�  #7��XN�N%BH��f����W�{}{�ۼ�{�Ni*F�P�$������ܟ����9TFo���m6[��n2�{ �s ��r���GP8܆2\����/7 �U���{�~Q�u��[���^�)�r�svp3Gn.ٸ��b���#����AG �ܖzV*�����@;�ѱ�l8��8>��Uy�;씍�x��I�C�$2 3}�s�<���!��>*�^��=��s��m�ZrEN>|s>~ f�`�U����VN5�$\I^nA��uf��5@f������
��L5���$�Z���E��Oi9��vmɱEs���sn���S�rF)4F7$���U���ߞ���A�̌�ӕn6�����=�{���Agqz�Uy����q���;�y��[�٠P ���3�:���قZq��#EPw�t�y�{뿼���V�e4W�xK~�@�}���A��&H\���U������a5���ł) ��L��\6>�{*����V�6�\Q��)����W�.����nf#�uS}]#[�4��Lleۚ��4䊜|�l���8o]����vF�"�Iw��s=�v��wN-EHъܓ�}��V܃��J��^�ރ���m�fG$����>�� /=��}�8l��@P���$��2Km�  X����9��n+��]g�;�13�n�v��:�{;�w4)�f�<#Ў�A��`_5v��'uڭĆ�WR�k�rl�4���s8ۖ+E�n�`N[4;��j�9�J�b�Ҝ..�ݮ&�����r�8YM�[����n+Y���n4����aT�N&N[���\͆��Y7dL��1e�C�Fw��};ۖ;rs�����u�8��Zvo�~�ߥx��`��XFg���f# ��Q�3=��*��=9��=�w��Ğ��:�I���l��o��������)f{�ƽ�(C� ӆD<}��/u�w��e��>�v"rD�1�g��w��ߍf{ �2�"�D���Z�*���8���;=
Vs�zH�s��Z�6rC��ȑp6���9k]�ׇ�i�^�Z���1�d��/�/�'0�C��Ct�@0���4��M]���ׯZi�)�e��7}�^����o����M�e@�r�s�=���/�M]��ޫ�`bI�ģ�fnA��zk3�}����V
�$@RED6T���rv՗�t>)��{=N���*8;�Hgՙ�ω߶��Av�x��8�95��
�@�`f{>��/����	�\��(��;�`]���x�H�������W�����~�^�RB����n��9kfg��}�[�6�#F(crN^��܈��ә��B���}u����qW9�8�0P�GD��=�W;4�J`�-���dq�m[��U���gqx�>�X����Ԅ���ή�ྯ�۞7k<�@�08������W~�W���7)IRB�7�g���y���b8�"�X@� ʴ�)1D�UpG����ӿ�τ��q���ܕy��3=�w�*������m"ASP&P0�:�-�7;7��Zxp��A#$IB�NH�>U�]v���q��=9�H/�e쑨�MM�g�8ma���]�u��o	R4daG#��5x�f�ߝ]���ǅ����B����H��W~�;kƶ�7!����^n"���V�6㜾R�`א��g�ъuTk��������4��Hl��q!=F/�A�!ۂ�P��F!�! @����f2�$ Ń̫�ŉ$P�1���'BO��"ćQc�B"��!A"�`AO�B�V��1c!�D�2o�6�����Hos;_}�jh�	 ��,`9HA� �`1`�"H��"�1�0$����3Xuf�:p H 	d�K!�
b�gO9V�  m� H�Iڵ�z��  ��              ׇ�tI�[�������(NU����@-�z��H6.m��XG��E�����)�Wl�R��#9{Z�=]��r�ބM��_>m�����ې���V�GZU��PFZ�x�Bw*@�L ��6�����V��
5K��4�]V�
��m/@s15�I�a�z�J���2D��v�ET�ֺԛ!]]���Ξ����8#�@6t����O5��W�v��u������\&�Ws��\��#�29콳}�c�����I	K�㨁�̛Z�1i�B�E��=o/Y3yIѮے+vG.���'v�YT(Iv9x֨�vy�����mp�p�p�袩X�t϶�/BV�(ϥ�'Hs7e[pm$��T�5v��W@F"����@��W@��@f�\b�K��׭rv�	qn�]r�&�̆%.
�Y��[eW��O�ݜK���s�{s�p ���=vۤ�m��m��\�Y����k�����1<���J�8����r��f���ZN[J�UK�UHu� �l .ۙ���-� �i�X�ۍV��c�:r�u�q�f6��A��<�%j��(B�iV���(�J�c�#�CyKC�Nm����W6یeك3v�Y�+F��4ȴѝ�#.���ڥ�ۣ�{=�A;��T+s�mm-�9us���n�b�m�qS۩�d���[����������ԛ���m�eVU�$��f]��s�;=>4:I�l�Y�ۗl&ۛ�����Cß?���P?H��p�_�|S��(?��s��o���-�|���l  Ug���n�7����;�c�r��^F�c�f�K@��p��JGK�aj�m;D���:lӍۭ�6v���i��v�ٺū����0�ϡ=]�2Z�Eˠ��������."ռ���V��.����B�= pQ���˘�4n�n�Y�h����{��{��w��?�����v�&ۅSt��m�F�vй�Ӫ�x�1��bI�&�u�/��;kL�g*�ι�a�"M��
H\��^?�37%fy�߬Ad��t\��CY��r�5��Pw~�3��Q�O�O�r'$L�
rv��]��v�#��{ ��e둦��M�g�f=5��Fg�V�{����ֳV��A�Up\=�@�=x��@,��k�lN<�&p�#FFr>�yi���4�y�3=�{5�L4�D��8k3�?�:�"�N]R�E-�z}�%
����2�R�D�.wH���o.i�_��Aޫ�& ���p7�Gw�b�W~�>��Hu����sU3�UMMU<VP��2�������p]����4�d��)9	n�v)��m�f��y�� �ô������9_n�@YC\��/�(KI�:q�􋦱U8�&QQ�>~�����x�`�O�h�K>��"��	.�u�}�;k�� thLU}T(sޜ��󯹄��h��kX���E�gem��XYD�����B���L˃���	e�.� �5��e���M(aP�n�5���M�;�9E�#���@�G��."`����;Y�a���/�� Vg���=�8�$#q��u�}�9k]�fWo_��w�uH�����Μ���ܕy�W~�8*�����I�BNE���ʽ�W~�?�\ �F�,X�P!�>
��`b�J	="� |8�����r'$L���_�u�����\���H�9�8�J�t�vj�ϛ���-��n��H	08��!%�[n�7 �5��s�_�׻�4$��G��^?y��/�,ߚ`{����e��8i�*��'|� ��`v���>��q�D��A�"7},�`���ߚ`w�z��M17.%̹�/5����`~��\�R�ٳ����X�� -�t�v��ct�p���[��ݞ
r�����C"gn�l���ft{A�ޞA�v�(�2ڔå�@�R" ��q�z2B\���_���_�z��Cn;�ٗ��Wt��˞,	Y��1r�8��9]��)E	l��1E��Cb���U���6m�K~�������e��3m�v��'W��j�e����ɹV(�N��������nB��'��$���I_�������Iг~������s>�}T'3e�ѻ�&d�0*ϓ�Kq-��r�3�������������D��[��Z&&h�i�w80<��=J��1g����5�j�[�@fO���)foWO���U��L�Qk����؝��%�n쁑9:y�=��n�v5ͳ�G#��0�)jQ2��4���E&�����L�����!6A-�HKT����#�\\��c�kꀿ|�3Z��I�����EQ�	;�A	7x���0��qr5fıľD�KTd���Ƙ��s��=��г|`��A��g��͂���	=��o�L$����O �2CFu�>�Tbmn�Ό�� ��5ɲR^������w�����Ƙ�с�֘������(���&�`����m鄛�A
����ax�M�	��ە@eΌ�4��>$�&�����Lw2��1-1�r���0̖oZa�9Ĕdߡ���P��%�3-P{g�@^kL��0;~i�A��Q��D��ӝ�;Z��s��Hz��7k�G7J8�n�a��Kd�I̹r����0.;��������I��Ñ�ÎRb��'�O(!+ͥ@�oόQw�(�-B���D��TY��������C�jx�n%�AU fl�;x�½P��]S��b�P��tBO=��.8�p�13G��4�Y����L��U�4�D�DKE�p%��1�97���RK��X2cu\�����4�ߍ����� ����2�ZP�z��1-1�9e��0=�4_�`]φ���#!I
��8ZG3\>H�k�R[��	9��	=�j�9s@e��Ŭ��4�.�X�Y�q29|��%�#6�n��3=,&��%� ht@	U+�FĆK�F�  ��I�f9#�`<M�n�ڔ=k4bj�q�Dؑs���&v��N�9�RZ����5���[H1��T��y��<m�����X���m���<��ZVE#5h���㳍6݃΄9��X���[��\V��9��"6糺s�*����wi�q���~������]wc6���}ý�p����]�l��L�1u��Mm�\/1q�i,���K��_��|0;����$(6�b�����r�I�I�d�ݸ�Y
N \&��N砄��с~Ƙo����1�ԩp8���сy�0���qF_�0=� �jRM�\���?���I�֢'2���Oq��O�C�T2bMl��p���m�e7t/#�ƌ�S&�N��ܭ�n�ۧq6C&�}�r���L����3��	�y��.3Q�n>�s��@A�x"�T���Uz����~���N^@�$��ͪ�~�DَR�	9��w7x8~�Oo~��'������	��$i�jG~�L�i�}�L7�(�~��\�r��
cf����i�`\�2��y>�i�ԯ�CpBp
H�$�L�d�m�G��wY�8�;n�q�X�׽޾���7���i�ۜ��k��Υ��ߟG��K�p9nUy?�i��֘�i�%{5��D�#4�n;���b�i��;_�����X��2@˱FVTkԤڕ����J��V� ���:
�B���ῂ��� i�� D0A��a��M���@�!C{��%X�"E4 �!2!#ګp9u�"�%5 E�A �<��D�E�P4�Us�0������{�ӈ��@ ���=jj��� ����䪆h�`�������b?���� :��%m�4�ܟ��A���(��6����@e�L��`_��}��c*Dn4�$��Ļo$���o=$�(V\K_BD!Gs��5�)����9[��K��t]�<��>��P���%�}?�i�����A
2�I��\g�̩p�)nbJ=�0=x����!'��f��p�ljF�� |�t�4�̽T���/'�=�0;�s�8ґ�"�p���!'���M�A
?%�S������	cjSp�[j� ɟ��d&oZ`_u�uJ���M�E��,r͇j�����ѷ�����]HK�i��l��7Z`v��֙�"�|0=����[�Pڠ/�4���L����ݥ@<��#�rሇ[n%t=������0;~i��[f@�L����KT����Ƙz/=I��7Ԙ��9�.�#qP����8�W�J���L��`~H�Z���pD�$J�P�+�R�
�1@�@9$Y	�>����6�  �^�rDA��LuX�\ҦW%�m�D�tRfGv;R6�+;�lvPv��i�V� c=�k��n@=E��E�M�����v4����v	5��ծp\�|m��jӠtnHT��Y8]:�`�i�*��m����N�:9�[�7]K�O\.m�o���\��f� )�e�y�4�x���ˆ����22�`�+FH��V�x��F�bIiFŒ{�ʄ��A	=����{`���F��Ԓ�"��'/�NUDz/���ʀ��������n�m�6p`^bi��\�Q�ၗ����L�2���Y@g�iP����x&��`z�����ĩr���0/���:0=Ş�T��c^�"��L�%��DF�4z��N��KDb��ͮ�����f5dH�B8�I�~0��y��H�*qn(I���)��3�M�� �B��*����Y�Hݿ���Hg��ˆ�KsP���y����Ό
�r��r�nT�9�A�2t�?e�(q$�i� �c���-�D��"b�s��80/q�m�P�`P�a)�.'�E���y��xϫ�4�2\3�L*�uvm\��E��w'F�cL�������$���'���A��L*/��ܟ��`o�`��ɗ.eD��3g��83��z �U=N��3�l�����_f�#�rH�1�Ce�>�Ɇ�4��ΌŚ�8�J��9(�сy�0;s��oJ K3c[�Pq<��M�6�8
(y��6���=�rj:z�h;��2�m
[����֘�80/����,��	=ӛ�܌I#(��&���*��@^N��i�ݷ12e��%8���\Ps��[�I���`^4�D�̍ʆ��(����Ƙ��0�!P�8��$���P�0��L��%�f���cL
�zPǦH��x	��M&Zf(J��oH��s��F��Pu�f�0T
0dp��i)I�	��O��pp�.�MK�������b�=�N�ߜn6�K��j�nk��3g�/`v������a��ÒRrs_����i���J���Ҿ�/g��2�m
bXᢁ�?���ǅ�f��P�[R��r�f����V�	ߙ��'~y�6I�Q(@@�(�`���M����7ll�n� ��).񕣥ہ�����lf�L������ä� ����$L L�Y�uѵ#x���ݜ୍��w:;oQ�n��.�Eݒ�q]6V5����KS9:��ۣm�v��k�g���V�:x�mj��T��y���R�2CE���N2Ɠ�0��:zd�/?�A�9���8鰹�]2f˘\f7j�]M�1���J�qP�apI�Ir4�NJ.	#�	;�O�۝���A�֘�7Q,s#r��2��>�Ē�L��4��|��o�"#�ڃ�D��p���}�x�`v���/'FfJb!�[�ڙj�ˑ����ǥ۟>\�>���	;�~q��u��	7�><$�ޖ�4���iP�bp��B��.tM���t��m����6�^�g-��\JOmv�wr��}�J�ډl�3gၼY�J�����̞<$��#(r4�	9�� �@U]P�װBM��{o�|(�p��F�N8�IF8I�zx�y�O<��=0���BIﭴ���\	�8N�Fn׊�|0/1����%3���i��c��nTr|0?�.f�*$߶���ϸ8Iϟ�^�DKH$"Ef��P�C�s�y��<bgn�Q�M�d���}����"ݩ:��0;���̯ع������	%)�䁸8I�lfz�7��jGu��Nn�<�Ys5��m�R4��3u��/'F~H�\K��∍֘�i��ey<�Y*[j%���5�UT���03�i���>�/g�=-ʗ"!KsP���^m**"�=J��~0�EP�V6x!4S��QTE�2�9��zw8�٠��*���~}���}���c�'��i�ۼ�C���
�i�ݷ0�qD��Z�eP������ɾ����0;0a��麉c���mP��y�mD%ȋ�4���R�=�m(�%��C�����Jo�J��֘��*�������!=@03��ɰ�{�w�$�9�7	��pB~DP�y���3g�E�4�� �DKܸ��w����s���J��懬cn��4�����~��}�,1"nbDK]7}J����גI*���i��^[�K%Kl"Z�/'����Ay�0/<�יJ�$��������9g������!ڤ���s_����8�.'A��Ծ.qF{�Lo�J����s�/2������│��	>��o�I��+̷�]*m�F�����.�S���|KF@�dHA�����c�B� Ra �"|�!�_E��Om $0�CX%2B@�1��V Pt Ԉ�=Q
Ai)d�0���E�|��@0H�a�#$�
j�M"4"���hj�!ك� $2�0��%șE=	�@pP����!{�L3 }�Ԋ#����O!d��XI�	
e2Kd�����  � �	��m�h�ŽN	 m               V疩�:�(6���4&��3l�;�[�JvY;,L�m\E=��͡5�6������1#F)p-f�ô;��b�ѱ �u�c`)���[;r˴쬱L�+Aqg<m��J̑������[[��t��I����RM��t�p��{qTk���ume����֛��3��9���ݴ�8�m���tݮ=vN�8h��X�v�⁥8�WK�J��9۷$@ո;�0���n1�Ea�X�n�㴻d���!\�M+*��u��b�Y���ȱZ�'�;4C#�R#x�gyN� <܅��
�F�G�:���a��d����� 1�V�w6^�����*��a��C�p�UTK��N.k�Uk\av9��\G�iR��<i���l���:ɻ"�ȼ�6qZJ��J��T�! �c�YJ�[D����]�Zu�[N��i�®4R��n��������!�g�ɫ�WZ:ۭ���VHͣ6�ep)�9��ԫ[+��=��.�
��Q΂��gu� Ͷ�Gk�Vu�m���0#�&�R��z�S� D�c=���� �ZS%�T�*ҭUUVQ�VT��H�&���%�GV��T�0�<s�tRݵ�=�timPn�L��fcu )Q�wZ�� T�\cr*f���*��Ɏ�l�ٓ�l�3��aC.������Kìn5���@'c���UrF�R�� 
�n�9�Nܠl���\�Yx�*҅��ffr\�f哟����
H���p�-<AS�~@��H��*�?c�T8��@�B���Do�DJ,���/��i�6�Ŵ  	�m��
j�A6���V3i�f�2�J�hӸ��2\E�pR�UF����Og=���.{��n)q����c���;v���Omj�N.ȆM��ɗ�ֻb���fu-��=�]g8���bev2+b�(�ѵP�6��v����aP����]�[��b6yD���<�7=�;Eϓ�.[rY���U��8�0�AE$�	;�G�wm3b/>j�@{wiQ؏o���a��&(�i��Ƙ��T�鄛�pbIJR9 a��s}$�nҠ/'��m0/�{.drH�&�"Z��{}�;�>��a�y�L����Y)��e��|0�^e&�`z�)P�������)4�G���iSF4dmi��C�3�#�|�c�b�G~�7�M0;x��̥����}?��>��6���S|����A?�te�YI�������3��rI�y����˂~H�셦�5%-��V�����Ƙ�i����%�j\��+"�џDf�L�'��^(o���_�2�,�3u��v�WoJ�t~�6.##_ÔK�@Ǵ戼&`NG�p��;n����n�N���/��*7�0;v�/'��U��0>�{��R�8nb%����‼�����0*���%��mL�P���w�|r��D���9PR�u~��d=�xP����r��%KsP����0;v��/'FYi�&\7.T�C�@^k��y��@͟،�i���α��tm��n-r��Ď$�㮶\]jg���燷%$C��#��(�lp�y�Ǆ�Ǧ�x��D�zI�Ӛ�@�AI�y>��3u��`v�����@}�k�0��c2����A	7�>(7����N��aԷ^��8	r9 n����uP��P����^�~�\T��"�����ׇ$���|�ͦi����j�����/'F�e*=��kd�� ~z������!���Lͭ.q��h�t*���GK���m��į���}�u��6z��e�����4�����oJ�Aiqk^R1$e�#L���� l3},���0*�Y5�*b!ʠ/5����>�q.L�φwZ`w��0�q0ءʂeP��P���a丸����*ѦhKq*\ۙelA�>�����~*I��
��!�RIK.gۻ�l�v�m�  ��B�鴉�=z��8�2`�X Wumv[�+Ӂ�ڈ�kq�vp��;�x�]��ygA��6qv�aP�6�{NM�9[��M�x�Kum9�)�$������Z:yʵ ������PuΊ�۞6Ɯ��g�nV껞n �U�L�2<��I�gfn���{������֚KG,��g�����lb�����y�74��t�C���g�4���Lݿ��I|�J�i-���O��x7.G$��M��O�P��ɧ����	7��>B�SgW��(9
")Nwޟy#��a�In��=�A	<C��)��l&�'��K�E�����_T��2"/1�P����@���<$������P��P��wq�S��P�I���n�:�-�v��y�	4�/S�c\���ey�0;v�/'O��_.s�vC}>��O7��T*�����_���*�\I�}?.���/>j$��F��K�n6�Y@^φ�(�4����@͝���-K�9(<�o�������Ydφd��X)n[j[(f���\K#+N��>������MDC�J�	���Y��[�(b��X�q)!������,�$���=(�сy8yqT�`w�P�7L1H�@܇�R�~3� ��?yT���s��̟5��U���`��#FXr4�	9�������UW��U�������=s�`U��j%C��ʕ�A��3}\`^cҀ��>\s���(����bq�`���NnϏ	=������?	���0/�C���$�=f����vq<����gtiāiڻ]&�	���\�<7
s,�/'��p�@^y�Uy�� {}>�"T5.#e��?��I[K6I����M�3�Iשhj"%�m�-P�i���V�l�`^cL��%��G�KT�f�xTn}6Iߞi�~�6 
C�
K�Ux*�
� g=4C�Z���#mL�P�07�K7iP�i�۷ㄗ�|w���qb�&�(�����:Qq��I�tM�����t8�4ݹc_�����䘳�۽��UԒգ���87�&8n\��s*���O�m�*#=��~��(6w����p��[��g��*c}�i�w����R ��8O�UP��|�'7`���4��s�E�}�@�O�T�j\!��P\f�i��/���ﺺ��U��C�~�Ө2;$��ܹ����ٹ�  [z�E�^;;l�r�V�3qQ.&M��2�n�į�ȥk6W�NT�Y���!LJ��q6����K�v{.�k�E��Ӱ�H��R�8�8&��<�^x��#	��J�6��KjNSm��j���wmwa�jNܣ&29�œ0�;);�s[vf�����N�z�d�r�X�T����̜vqͥ:<v}Zӆ��	�sk�^r��k�_���yJ���G��$�@f�L&�[��n#FH�P.kG7}��%��Eym0.����\�;�51�a)�jfZ�67��c7i0>����y�R�;�h�SR�����0>��T�z��..r6w�����L�n\���r��4���R�23a�/1�|���i!.J��p�,�b!�mt2����N��d�Lnٺ�ߏww����2V�屗� f��@df��`]�L=�A�20����N���U@�@�(5"T?
*���"	��}�0;v��� ?o��*T�q�s���'3`�P+̟
���C1cX�
I�|r���'�s"��Z���� ~�tBNcߘL�ppm��@^c��>K�\[;�3u�ߚ`w���˖�$J�L%>��a��VO៾� �e�&�I<�������&릺e��</}�i�w�^�����½d���È��I���A#��s��̞<$��(I���RD�i(����xQ��K���]�'ǽ���{�l$;�I��$�$҄�p��o}�«�$�:N���PfR���F�a����on�@� �T͞�c�����ΓF��pH�xU��x�qS��!?o�P�� B3��?���$&c�����vv{q�Ӈ��ߍ+��?m�Ä3���v�;}�{v��).˛r\��!�`a
B� B��a��������K��qz](�H�:�� B �Ū�P�N`�� ���W}:�'}�BO�sb�-D� E���o-)�{���y�0.�i���[��#FF��zIz�˄��W���z:��#�o�P���9�EݑP�ӻ�mۛ�8:͜��1����y��5����Ԩ�i�۷�yΑ�zQ�S����"T�9j����W�n��yO�9��
Hݼ��F d��8C7_�"����`T-W��r�N[R����IF�z����9?Aڃڀ����	^����rI�y'��d�T8���0/1�nޔ��BO�s[=�*H�
i��lg�t��h��M<-t��b�����}�����r}ܴՠ=��0;v�TE��i�{6�5�\����Q9�<yڪ "���03u��`_�f!�r!�Pۙh�2/a���֙Is��#=�0/1��=z֩R��n!��P|��o�I���BOn�_@U=y򄝽0hjS)�|r��֘s��/2���`^c��xmP���"AC)��I$� �K���M���;e]^S�F��.�`t-��L�2&ɸ�p�8,�`�Z�$�npʰm�òqv�gd�)�kp��l�3\l,'^��Rd+�&H��ד�'�n��7Wl\c83�KN����u��(q��e��%��4v�@SX�]�꬏L��svy�����{��;���je�{w$\)�99��Rۅ��Eܛ��������n�T2a���&�����2/a�y�0/q�B�&�[i�je��Ƚ��5��A�o�T���+�@P�UP �����9)�ƸI��D��Ƙl^e|P�d��{�A�!Cq4J1�}@
���!&�&�q_�x���!':��j'!�Q1�M�M=��\\��E��0/��{��f�:[p[g�C�[���q�ۡCkN��e�%�������8À��&F#�8zz���݂_����A�����<�ކ�R�K�CUU9m�(y��Qi@�*��B���<V�BO��O	8�������6�r���o��`v��5$�����-��@]϶P8�(p��B���R�2/a�o2O�UPY��BOU��'$�(��z�?o�J�߼������/~C���V�wcc�m��ُ:�;��M��gdlEs���է3�.T��C��t��`^cL!v��U
D��)ďp���$�IC�A�{��y�Ҡ63!��Ɵ��	�ǡ8Tp��*"�	9��%�|�?��7��I϶I��ǁ'20��88O�T���%��BN{`��*�����>�?�K�CM��3u��A>H�d��'VyBO�ib�P4��m�%�$�������	�jxAx�!`#������F��LK㖬}�L���C��HݿkIPp���Ǟ��Z��@fl5��֟�qD~G�pܱ�je���ϡ�w�3�F}�0;��@^H{A˕2ܑ0'1@e�L�f�9�{����>�~����������H�-BO�gὉ�Q�lt���0?s����@��C�`}�%d}���;s���!�̎,3��[..�3�=���ў�e�)��(��&�g�	8�T$��f��.W;!�y��J�"e�7*s)�lF�}�i�~Ƙv�V.}��c���I��$���8�w_ў�e�!L�㘘%>Kj��k���E�0�Q���s�Z�Gq-�%P�~(��`^cL޴�?�B��@W�s[�̍�ҍ�  	,n,ݳdU܉��N����+%�p�ԭ�X
-(bD�O9c	�	1�;.W;R1��au5q�m�2�Xp��ǝ�M�ɶ�b��]����5�;�.���q[bWfl3ւm���s��M�A.�Mgu%.}kAr�c��) �P��-WZ�UZ��n(�3����	��� �$�4�^�̓k��]��gg�����.��m�hx���z%�]�L=̯؃6Q�nT����P#}��i�۷‵���${�4�6�'�&�	9��	=��xU%�~P���C�Y�M�H�p��!F8O�]S�{�u{�J� �������C�Ù!�2��6�`v��nޔj��Ƙ�RVvQ]k�ձ����<��a&�OW=tX��{���/�!��p㽈7�i�y��vߊ�yBM��)�*6Ӕ�$�̓��0\]�Ļ�{��������L�}���������'��O<�žP��If����0*�#pܱđ�؈�K���%:��0)-�R�/>i�Wo��W��#F5�O�}��O�(WhP��tt�{���E,[򄟶�{W��"-��g��Y;ml��-9�a�G� ��E��G.�َ(����H$���'�s	?cߗ �֥�]�㘖9lQ2��*���⼸��D�`fkL��dDnxku
#l�!n�qo�$�d�?ʪ��fD�?E+؈���Q͙�����@~�z(���q@n�L���љ����C��3/�fbe7	9��~�*��  ����>^�MH���*�`����"����K��cO6}��H(n��`��y9��槰��5�����R�23a���yq$��@fy��OP��D�G)��N��Y�1ߚ`]�zW�.(��Z= ے[��1��O��!'2���UB��2|xIվP��7���R�*1�v��-�p�'�y��I<�}vO�}S�1� ����q}�Dԏ�OF�1�Bn9Tf?�#6���A�����_��G=h+n�ƻwe������	JCՂ��t�	(H
��j(�<Ԏ��݂w�.qr�31��=�~	�J|�M��D��S(�i���Ƞ23��� 9�4�ܨ�-�Rw}$���éj�(I��$���`�
&$Ĳ��IE���������֥���������Z�^MĹsZ"Y@dg���cL=�������r8��w��ﵴ�����[�:�$�$%H* X��)$)kB�"V�
4��^Ζ�ԂW��$8�u&T�=#@�,`B0�-�4Nȁ�&"8����� -���@��"��i�;8(j�P*(vr��aKx �<��1��ۄ��xH:y�N�c�7�U   �k�$m� �ŽN	 m               ��tk���t�a�z�>�[\(ꎧa��D������qg�p@Z(�ЄJ�[s��eA��y��X�N�:�iw����o/S�-�v�.��c��-T��Z�V���1R�֗4tN������UXԄ<
ѩ'.K�ODܕ`,��l�G.hwi�]��Ƥ���P��r p�M��B�$ޤr�(�)���4Vx�����@����;�E^W���Jtoo$mʵYn��oA��i��l�����:2� m;M��+�iiYq`�����g�θ�L�S����
���[�[����^\��S[m��^�%�I�̻Vtgm[�P⹸�ν�:��� !��ͤ��A^f��	q��5\��,0iצWi7Wh؎�K�y�>� ���Vր�]m�xR��`��m�de끯N����I� ��f:zK��*v2p���1��u��!�kt+8�i�]��Bk]k��#LG� �sc��nS�OaLqk-�{,<û2�J�PSű�jks=��U��%j�Y�m ����x��6r��Wl��*�l͛IҶVJ���ei�
ݳm��j�ʵkA�JK\�! ʵUU9JyYP��s(g]�zb���ι�����Ch�ೲ㬎%ئ�uڜ�[2K�(��*��n�kJ��'g�`.�Qv���s�+�]��W��YaS���g�{/mC�-�{�vB�A+UT[e)ke��i���3]C�^mZ���m��ѷd�i���7&���c舿��
j]WD��	� ���Q^��P@
 g��]���#l���n  ��v2�sl�]J��ؗ�x�hmVMd�p����I@�j)�v�M�A�X0V�����c��;��;�q�;�q�Rَ��q j\��-�h�t�T�i�i�]����p���u���X��e['liS�;I��l�N��pfا��v�8��^�G�w�����1�Ǘ�u�^�lp�WNܷ]	�Ʌ�˪%�]%΍ �D��_�'����x�@w��"�_�8��z=�0��7݆Ӊ�)��$��$��0�<�'��O
#��v8�PB����'j�@v3a��Ƙz��`�D898T���Ak�(I���,�'�A]��({���O��i�wZ`]�L�w"��͆ �v/0!�ʙ��������:읻8m)c�=��X��g�{����}�oiH|�j���Q{������������D����CT߶�~Q�*�:�վP�{�A�"m��P�����ne�hr����`VcL�z�w�@v���2�!���֘x�G{{J�ˑs��qs�f��NS|o�t���!'��=��N��BOs �����PB�G)�Ҕ��qVH�^h�x��@F�c��y�z�6r�t�n�I>>7Ԩ��`w1�޴���3T�d����2��cL
�|`w��9䏷�x6�J	"�R9�A	���?F�`B��
P�� � U0"%pa�,���zw��}����(I��p$�djRpp��KvZ`w����e��.~����ݝ����r�CT�}J�/vX�i�%�bu��59ı,J�N��݄L��[�<��vD)��%V�5t��i�6�Hك�9�8n�ݻ������%�b_>�5;�D�,L����bX�'^}�C�u"X�'�{����%�bX�{�		��f̺m��uı,>���"X�%�מ���Kı;�Ϻ8�D�lK��٩Ȗ%�bu��ޮ�ݹsd3-�8�D�,K�~��U2%�bw�{���%����/����Ȗ%�by��59ı,N���nne�f�n]8�D�,K�=���uı,K��f�"X�%�߾���K��?�=��hrL��h#C��?|%ݙeٗM����%�bX���٩Ȗ%�`��5<�D�,N����bX�%�>�'Q,K��<�|e�{q;{s��v{�O'I�q�6��"�ے�mظ�Ɗ:�3&�Zn��q:�bX�'�}�S�,K�^{Ԛ�D�,JD�y����%�bX�Ͼ�ND�lK�<��f�w.�\Ӄ�Kı;����bX�%�=�'Q,Kľ}�jr%�bX'~��S�?C*dK�w��l���n��.N�X�%�}����u��,K��f�"X�șϾ�Ȗ%�bw��ND�,K�;?4��H�eI9C��4���y�)bX�'^��S�,K��ϸju�L�`~L��s���uı,O=���t�3f]�.g��%�by��59ı,?=��F�Q,Kľy���:�bX�%�����Kı?F�y��'wϝ���]�����  7kT���vX�Yv�u#�nUn�Ƭ,���f�u�	c����{@��$�=r�W�鱹��v�K�Ayu�wPmS�#�d�q����!�5���[��mb�m��f�k���������Y�����ZV���;�G]'\]��&B���i��%�B�2Oi��jow{���,���m�Y���ܗdπ{Xl��\�@Us7�Lf��jZ�P����[�oq��O�����Kı/}���:�bX�%���jr%�bX���ND�,K����e@�q�Pr�Mh#A3}8�D�,K��٩Ȗ%�bw�59ı,O;���"~�S"X��m��M�M����%�bX������Kı;����c��"dO|��Ȗ%�b_<��x�D�,K��}&dܹ͐�ws8�D�,KϾ�Ȗ%�by߼59ı,K�~}�N�X�%�}����KĹS�<��̙��˥�4�wı,O|���"X�ʙ<����%�b^����uı,O>���"X�%�����o���m���n{u@t��;*�`qŻS^{=��[�GXX�a�L��Ip�;�bX6%�߿7��Kı/�}���bX�'~��@�K�����S�,K���>&��ۻ������%�b_>�59�����|b��Ȗ&���S�,K���8jr%�bX�����'Q,K���ys���3f]6�q:�bX�'�}�S�,K��xjr%�bX����x�D�,K��٩Ȗ%�bu��ܽeٙ�i�n���%�bX���ND�,K���o��%�b_>�59ı�{��h#A��q�QEF���%�bX�{�>�N�X�%��~�59ı,N��"r%�bX�w�,��Kı:��z73e�d��d���%�'��G��y�e��6I'��N�L��:�t��͇���b_~�59ı,N��"X�%��p��Kı>�9��:h#A���8<�N#JI��ı,N����"�ؖ%��~���Kı>��{8�A�,K��٩ȟ���,O|��K�&k7.f�t�uı,O���Ȗ%�b{��q:�c� xt��zh>�= ���6%���jr%��TȞ~s��"X�%�����\���0�N'Q,KQ�>�ߎ��D�,K��٩Ȗ%�bu�59İ�:����bX�'I�~O��sv��칼N�X�%�|����Kı:����bX�'^}�S�,K���=��KĲ�éh+Б(�P�"�$���r\(��Ѷ	�iZ�h����
����˹��ٗM��N�X�%���p��Kı:����bX�'�{���%�b_>�59ı)��sZ�B7A��c��h#A��>��D"�	"{��r	 �ߏ�D�I����?a�dK�}���ܗrݛYt�uı,OϾ�θ�D�)ľ��jr%�bX���NA�,K���Ȗ%�by����wr[�\��N�X�~D2&}�����bX�'~�xjr%�bX�w��S�,K�*~���7�3��q:�bX���贈|�RH�(t�F�4�{�ND�,K���Ȗ%�b}��q:�bX�%��S�,K��(����?G����I�i�hF���v;p�l�:w���T۳�R���I��̺\Ӊ�Kı>��"X�%��s�x�D�,K���j~N�dK�*{����bX�'�oޓ	p�M��]8�D�,K��y��uı,K���Ȗ%�bu�D�,K����%���x|#�Ƞ�B�<��A�F����jr�bX^y�S�,K�󿹓S�,K�￹=�N�X6%���/Bc��PD�(t�F�4�~�ND�,K���Ȗ%�D��}��u��T[��٩Ȗ%�bwg5��qDiF9C��4���pjr%�bX����x�D�,K��٩Ȗ%�bu�59ı,O��
����B��-�Ŵ  �<�Q��gYõ�pBR�+*�rL�ʓ�5\wH�=��Z#���{x���h,\�-��nn�V�mӉ���2�ڹ�n�xco��?pp����e���4vU�퐈�u�ù�C<@-�9�@B��lT* .��õӵP�.��Ж������[\M#�SȞ���X�iۍ���m����)nx�oz�u�5ps:�.�칒�ЗN�Ȗ%�b}���W��Kı/�}���bX�'^��A�,K�L��}�g��%�b{����wr�nM�.��uı,K��f�"X�%�׾���Kı<���"X�%��{����O�ʙ����8_�.�Cr����'Q,K����"X�%��~���K� �"y��}x�D�,K������bX�'��Ҙa�1�pr�Mh#A�pJ9ı,N��}�N�X��}����Kı:����bX�'���>&�鰛�a.�N�X�%���׉�Kİ�X g߇�juı,N����"X�%���59ı,O6~���v�`�8��9yݘR��κ]��vL���^'���r)ȹC��4������Kı:����bX�'���S�,K������%�bX>{�>$�#p��9�4��h_��p���țڞj�|��X��bg��s��Kı>�>���K��/�}����*dK�'�e�.�ͻL�.���%�bX�{��S�,K������%�bX������ı:����bX�'^y�����K3B]8�D�,�������%�bX�߾�ND�,K�}����K��P&D�~�8h#A��Dtx)`��Ix�D�,K��~���bX�'^��S�,K��jr%�bX���{x�D�,Kߍ-��M�����˲m
��Wci�n�9:ZnƮ{5s�De����3���J��kws8�D�,K ��jr%�bX�w�ND�,K���o��%�b_}�(p�F�4��7JL0�ځ89GQ,��ϸjr	bX�'}��q:�bX�%��S�,K��xjr
�bX=�It�M��]8�D�,K�7��*dL�b_~�je0�����ʥU@��jIH�H��$w�H�û�;A`]�"��bs u�Ѳ�}!O�!t���W��{�B!d��0bXBD���;%��*���AȐ����RwP���QlW0� �/0 hrd5�Ra�x�t��#אT(C�w�t%�/J&+��� z��|�^���T����?bwϽ�Ȗ%�b~w��S�,K����-H�p"���F�4��(�Kı:����bX�'���S�,K,N�߽�N�\��2'��߲Kѹ�2�3��JD�,N����"X�%��~���Kı;��{8�D�,K���jr%�bX��{�}>�a/���ŭ�ۓc�-�7���z��T�WI�*�([���nA�h#A����(r%�bX���=�N�X�%�}��4?��"X�'}�S�.Tș�d��l��N \��A�F�g��஢X�%�}����Kı:����bX6'���S�ı>�g����R�ɻw6q:�bX�%��S�,K���xjr%�bX�w�ND�,K��糉�Kı>��Ϧ\��.ٻ����%�g�@Ȟ~~tjr%�bX���ND�,K��9}�N�X�����s��������bX�P��}�r�M@���A�F��jr%�bX���=�N�X�%�}����Kı:����bX�'G~�~6뀁U���W8����&=v6�3��wk<P���T�`�9C��j�4����x�D�,K��٩Ȗ%�bu�59ı,O;���"X�%���<#���	\��A�F��y�\)bX6'^��S�,K��jr%�bX���{x�D�,K�Ͼ$�!�����q:�bX�'{�S�,K��xjr%ڙ"w����uĲ�4�\��A�F�sޕ�6˛���%�b{��59ı,O=�=�N�X�%�}����Kı=����bX�'~M�>̓p�sBf�N�X�%����׉�Kİ�#�~~f�Q/*dL������bX�']�p��Kı?G�:X��	�n����ݻ׮/��:��.���P m��;u밭�T���v�ŗam�B�a��V��n�vX�6l�[��6ctvs:�ֆ0�:��v��j�.�h{v��0�!n����ܽ�,Wv�Xk����/Cõ��]�jB�'������K�$#n:�p�+t�Cغr�s�g4,G2N`����R&���n��66�n�X\��Gݞ5pq�H�d� �3�=p�q�&�����ı/�����Kı=����bX�'��p��Kı<ϼ�g��%�b}�ӟL�wIf�n��q:�bX�'���S�,K���xjr�bX�g�{�N�X�%�|����KĦ���E��Q�(t�F�4�{���bX�'�����bX�Ͼ�ND�,K�<�Ȗ%�`��y�Mͬ�nI�q:�bX�'���L�uı,��٩Ȗ%�b{ߜ59ı,O;���"X�%��I��sf]�7L7w8�D�,K��٩Ȗ%�b�p��Kı<����bX�'������%�b{�O��m��mq��:�� ڭa�+��:y0�󜕠-�{cM�ܷI7o��%�b}�59ı,N����"X�%��}���w"X�'��.�"X�%�ߞY�K�7w0˗7N'Q)ı<������(�1zP�� N�r��}ϳ��Kı?3�n�"X�%��p����,K�&����n.hL׉�Kı=Ͻ����%�b}�}u9���M����S�,K������bX��y<�K�奛�M���N�X�	b~g�]ND�,K�<�59ı,N�����%�bu�{�q:�bX�'���s�.�,�6���uı,O����"X�%ڈw߽�D�,K���s��Kı>Ͼ��4��h!ci"Thڎ5N�cFN.�۶F̝���1�i�.�zg�{�/�3�7�'Nn��Q,K��ϸjr%�bX�g���N�X�%��}���u"X�ۼ�h#A�o��$A$���uı,Os�ϳ��? H�L�b~g����Kı>����bX�'}��(p����F��wO�8Z�9{���%�bX���~]D�,K�|�59��| �EP�C�u���럩��%�bX������N�ؖ%����B�Ɣ ȹC��4��{x"r%�bX=w�ND�,K���s��Kı>�~���b^�dO<��Yf����)�7N'Q,KĽ��jr%�bX�g���N�X�%��{���Kı=����bX�'��}!o_7[�zl������
b�����u=�o6k�ڳ����s]�s��%�bX�gߟ���%�bX�g�]ND�,K�|�Ȗ%�b^��59ı,O���\ܵ��.\��'Q,K��=��r-�H�'���g��%�b^��59�D3C^�P頍h#C�����a;wr�:�bX�'�{�G�,KĽw�jr%�bX�g�{�N�X�%��o���A�DV��E�\ ��E��:�bY�*�L��{����bX�'��g��%bX����S�,K�h'��Zh�,$)�q�@11�'�~p��Kı>�|�m�4�l��7N'Q,K��=��8�D�,K���Ȗ�b{�59ı,N����"X�%�{��o�Cv�ui5�s�[��B��ݿ�~�����1���v��,V��H��\���wı,O����r%�bX���ND�,K��8jr%�bYC2g���j�4��#|��"7RM���%�bX�y�NwS"dK;���"X�%��s���%�bX�g��8h3A��Ži(T���N3��Kı<����bX6'���g��?���r&D���˩Ȗ%"#C��	C��j�4��f�iB�p	�q:�bX�'�{����%�bX�g�]ND�,K�=�Ȗ%��̉�}�(p�F�4��㺏�N2�Q��͜N�X�%���{�q:�bX�'���S�,K��8jr%�bX�w�>�N�X�%�����~�W��n�0��  ko\�����:^m�a�vK�R�dG)�n��t����5��u|��f��i�=�`��<W��� U&�^M���;�4䫞�L3[�_*�5q��=\籕Ed�pm�mȑ6��4����C��5wk�^-KLI+k���,�;���m��ﾽ�%v�v���."�H���d�o&۳wN8�e{bW��f ڎl�]���{�Y,K���o�jr%�bX���ND�,K����8�A�,K����r%�bX���{.]	�7fk��%�bX>y�NC���,O|��N'Q,K����˩Ȗ%�b{�59ı,O;�/��.i�ݹ&�N�ؖ%���׉�Kı/�}���bX�'�{�S�,K�￹&�"X�%��x3�F�������F�4��Ȗ%�b{�59ı,N����"X�&3"y�<��:�bX�'�C߲�s7-�n���%"X�{�D�,K���Ȗ%�by����u�L��,K��f� ؖ%����}�m����c[y��3�/k�}i�IP�u\�\ι1�iZ�p���32����%�bX�y>�Ȗ%�by����uı,K��f�"X�%ʞ��F�Q,K�L�ﳞ��2]�.�fi��%�bX����x�B!����؛�����"]��2'���S�,K�����bX�'�y=��7!e��乷��Kı=�}�ND�,K�=�Ȗ%�bw��59ı,O;�N'Q,K���}2�݅�6�7��Kı>��<�bX�'}��S�,K��9��uı,O~����bX�'�o�ˆK.ܻ�4�uı,O|���"X�-��~s���%�bX�}>�"X�%��o��A�F���q�dT�9s� �8C�-]��g���E��tu�趸n��.i��%�bX���>���%�b{����K�,O|����`�'����I�|n��swff�A$O��b}ı<����bX�'}��S�,K���}��u�,K��d.�ٍ�d|��A�F����bX�'}��S�, =�

+Q"AT,Uh0����Ac"y��>��uı,E�k�8h#Aн�k�B�Q��q�'Q,K��ϸjr%�bX���l�uı,�@������%�`tE\�=�tJ4��hn���[.T��Ӊ�Kı?>��'Q,Kľ�>�ND�,K���MND�,K���Ȗ%�bw���nf�.�.R�p������獻W J��f6�ۏ[l�<E��������%�bX���ND�,K�=�Ȗ%�bw��4�Kı<�9��4��h{��i��$��:�bX���{�F�P�"#�6%������Kı=��~N'Q,K�-��P᠍h#Crf��@�B���%�bX���ND�,K��糉�Kı/�}�N�dK���p��Kı;�O)��6۹�]É�K�����}8�D�,K����Ȗ%�b{�59İ?G����>�
s�����59ı,OL���F"�HyC��4������yS"dO|���"X�%��~p�᠍h,��-"p���	�Q(�v3����
=��خgA��lt��K�p���d:�����`e�L�>\�����zX���p�L)�r��`]�72X���'fHd��ȕ@fcҀ72Y�Ģ7u��`z,�DK�\LĲ�=�,�M06�ݽ(�OI��Й0�s4��˶��Ff?��`b������[M� ���\&�k{Cs�-4�!0����J�z��v�@|P��)e�G���ʁ��9�3z�����$   � (��P� ":��Ǿ���18�V
'i�蔓TS� G��{Ф�,%�.a(B6$���[��O���ײ    	 -�H��Ā�8$  [@              �[I�l�-M����^͓͑��ke֜ �c�۳�.D�L�Ş�㛹 m�z����[�d�I����cCv���Jѝ�W�p.]�[	q*�T�s�.H[=��T�m���m�Qj����6ڮ	���
eC�R%:ۍ�V�A��%Y�ԯ�өJ�<����L�Yf���էG/5h�G/L8i6ܱ���J�،�rv;+����k�Fָ�����|]�(m�&�X�6�[{�����M3�q%���Y�u8WG?gh��Jٞb��UKѬqAO9F��:�[k<�W=��[FgC��[^�nŻ��l*��TQ�;�j�[��W��1�[pe�S,�6l�m"J�TԹ`��p��52@�/�7@�UUUV��!�I�2b�|3�����n`Xu;vz�۶���A�f|Q��W��uE�F�m��ѕՅ'��;��[���Ŷ�խ\��m\��j ѝ���,f�c���i���h6�"I�\��]�0��4�T<�.�E�g��N.�0pt0]��U��BV���J�䝷��ҫ>ٖW�aU`�[-����k�j�P�g\l	��M�j���V��dvX
RZ�-��� 4ڒY$�uv�p����j��{[=b�ܯl��&�n��5��Q2�t�'3Lɫ�D��������!���z I*Ȗ�<�4$�s�sէi�w�ڌIu�#S�nm��;<�ij��KH�DҬd&���(q�b�Մ�s����E�m�2�v7)�l2�h>���"'�%;SEE	�O�� h��Q���]��PEU� ��>���9"A`Ĕ�  u�sq��YlӔ��as�>^�� ��x|������u�n+���c��ܒh�a�q���*��#�ky�o�Em��j&l�����A�^N��Wn{:6�e�c��<��=��8k�k�Pㇰm*���F�nM���\�z�lHqv6T����ߟ{��������u3�[v��d.�v�P�UK�B�yAt�i�Q�'9Ęh�J3p|I�����2X���*�A���C����J ��`fcL{2��ͅ�~0Љ9NO��̂PB��2I����O�n�&b�7�C���{}J���L�xP�%�ܼި�Ei��'��I��� �l�@n�L��#Y�Q0��v�u��Ō���sќ-������ܻ����%qdo8���~(o%���0+��b��S��q6�<$��������J����$��z�n~v�+�9ĔA��?��R8�K���I�^I���@����N"T��F���:0.��@�,�i�}�q��e�1%��3�����Ƙ�с�(��p�	���P$K,��x�u�^�st��L>֦�|�GV������m����@v������>W�������r�-@c|$�=3��k���M��M�\$�(V^oTq�"���C�K�������,Kй�aC��`{�c�O�fHdľ���c��ݖ�81\��ز�.H9q3� ��`~�K�Y�J.|0*���3�x??�]C[U��Il���{��!���j;=���� !6#hNbnf�̝���WoJ ��`w3(q*!��hj\�\��ĔA�ƴ�����ǥp�0�i�L�����cҀ3t������Qո��q�D��˜\\m��d�y���Y<�/��?G 
�V �P� ����}��'�g��)m,�|q3@eΌ����ܡ�OVn��YӼ�DKa2�(�m9$�[%�2��di9�;x��jk$\��	����E�}��:>���T��������s0C&%�H�P��U��(��zXs�
�����e���r(8m�T����ўIqDnN�v����L��2a�s4���wׅݼ�@�,
��s3�CMKe�:0+3)Pn���Ҁ�����\B8�5.�<���t���-�]km� Ӛ�����ץ�u��݈��b혹�+��d�g����AB��@���G�}�>n^����,�Vw��D7c ]���.��L��u�l�P��v4j���9�i2A�Q'�6�0p�ւ�Fq���<s��v;q�qr�l�X뚼�aBإ�f"6oǽ���w���}�\�1=��lOK�h:�\k�Ձzs�˺7CEq5�.�UOd�����Nn�I�^TD�^�O���{I�4�Cm9��}�`Wg�|0+o)P�\�Q��FТX50��Ό
���[yJ�/vXw�9m9p�LL�eܝ��T{���IGq���1�1�C��|	ey�J���g�4rt`UϢ�Q@Ȗ�C�ō8�=N��=�pq���VA�jƹ�X��wYtڠ���p`UΌ
��*�A���-�����{�L�:( (T d�za'����$ߵϪ���n�I�8D4ԶP��]̥@z3a�W82M���4��7$�C�Oow���ձ@*�2�сj:���N!���T�l07׵�^N
ﲕ�g�*�[�e��u��f���#N�Ό���J��b��n�����;���84ws��u�P���<�AQ��v��`Ws)P��s��cq�BLK�K(��*c6����9�+F'}Vz",@�g�7:�$���$��\d˙�8p�ڠ>��`U�
�����R�7t�&&�2a�srt`Wgwr�����.R�^�&�H����a�0����]�����b8c���9���j�#R�@v�Fw2��63c�w:023$򙖛����2���iP��������Qո�#�m�r���
���(��`v���jݚ�a(Q,�C��:0+���{�uo��9����
P�� ��P���5ơn(�L8<$���`Ws)P������K�؈A���[�fL��θ�2�2!�-�'�-{F���sf���0�M9D��I7��	:�$��I�^�Ԏ���Kq�QE�p��50*�vt`Ww((�6���(��srt`Wgwr����YC��iC���P�с]̥@lf�O�R�M0�1�3�ۂB���I7��T3�����сK�|�"�H&�"�^o�Fن%�ܒ@ x���9��ҙ_	U\v7�ɭW/v��O)�y�9�j�׋]!��#U;wd�-���u7k���<n�C=@�P��n��WR=���w��^�`�*�cr\��6�w�t\�ډKnv�v�n���^��)���+��F�r�q'O�e����{���� #ԝs���7n�d�a��z�x�
Ƴ��l_|�63�H�Tl��i��r��h���@�7a�W80+�����R�7Q�C�*KC�\P�6�80+���Vj��T���k�B�Q�P���!%w2�輆\���'qC�%�ľ8�%�ݥ@lf��pa�qG�)0=��.f861��E�0*���`Ww)P�ž�yLy�� ��Q"|@c+��N���f���[`�v{<%mnD��Inb���L]i�^���`_U�.[�]ɦfm��=��7�>}(�A "t��D�@�O}���y{�BO-�$n����p@Ӎ���&�ޥ@l\d�*��`uGU�p�G-��T~��f��:0=�i�]�R�7�P�J��j\�ܝ%�gm�or� �/!�]�ciĩHj��-��>A�Ee9�n�4E�qef�\l͙͚�xe���0+�����`U�!�w1���8d̾2�;{�%���{��;���.2e���6����m<�t��n��v�*�P p�N$��{��H��@!1�]�a�ú��8p��4��Q#�܌�!r�/iE�BIC�w�)R`0"�BB@���b�3R#�2ӄ0шi@K:�F2@31����S>^��xD�	D��0�C��	�!)4wƨѐB�rsǶ#�:ު�Ǡ::�`�8ʬJ$�lH{��	�ǚi�	[E z�нW�# ��gCГ�k�C�R,BA @"Bx0c����z�`@%^��$B@�	�`�`v���}����u�"��(r{��T )��?�]"$��%�K�.\�{��ׄꘘrq��r�(?s�/_��&��e*љ�O�a�e�D�(�i�5�ή��y
���U�lcbp��5n���ۀS;H8s���e��]�7K�ru���-�D��9Tov� ^�*���ꎭ��	B����@�K��v�;{��˜I(���D2TD�Pӗ4��`f[M]�R�7!�]�&��Knp�w`Ws)P]��3d�?;ʠH���FH� �"B
�! �#��,��"$�0`�b��,H*d�"��I  � �$�D�C�^u6e�������s$̾2�.��U�����N�˺�}��~O��`����x��udNxۧ�� U��CsMIם&&�,������O��%�W807-��t�o	�10���snt~�J �Ƙ�m*�Ap}��������P��n~��0+/*J��k�r�v�Q2�	�xQ�y��택XF�
>��.�����I�Q8�� �V��Aͼ�~
�����j��M6�
�F��)$� v�Uy|�U�ն�L�y�$<<�L��9�S&�o�dt���z��U�0'$����X�1q�
q��Cu��O�;v��b�����1���`l�C�n��E���+�i��[C̾1fK ��WkGV�i�n�ݮ����09u���k2��NĜ;s����E��uo	z�d��m�����d�]�Iq�B�vخntIWhז�PC����w����A��G������x�iD�Q��(kv�e�}܃�Xk�kq�܌��8�����/��s�nw3�5a�"rEFC"���9Ն�;�so ���4�f�R>��Y��9����I�yS���ݹ�ۣ�%��@����-��Eۘ�F��R*�C��kv�e�F���m��k�����G��̓�;C�B��  x
�]�  �$�Ƴ��t���̙�R��%�p2��k<�y�)+.�jC	���v��s2n<5��A�ő�rDL�ow`�c�]������3ش��DKi�(�T�	Jk�]�/T�c]���Ԩ����6��JN���*����XD:� �Vr0�qQ�����;Ն���sU�Յ�i�ȅ��c����s�7����'vOP1���ߺ�G���2��I��3p��ve�5��Aά5�݇��i9$��ws`�omi�s2F�~��
��,1i�i������ݖ��ٸ���aJr0"�E������܃�Xkyy6��3^�	4"1��;kMf^Aͼ�_o`��x�h8�0��^l��^�������8z����1�.p��=�w�u�����$T#S�U�P�g��Td2)*�c���W��9����B^�A"r E2glj��6vM=�� ��;"�[�\�����I�d�gE������/��oL5 q�&X����e�K/5��a�s�Uw��&X�'$iN����<{kA��������r�/=:����m�tnln(.c1�v֚��Aͼ�e�>? QT�0�O�3뻻i�6�Ͷ��D��eRS)�Y��!�5ۇr3���툌g%�ۓ�E��J8m�{m�[<��L�؋M+��U"�Ok;�[lS����7"s�;�����\��ʧ[�q�j*Ѱ�u�;9�U��5�bW�b�:Ьa���3����:^5��$۳�c��i��˻���!��Q����l6əd]���gh2lq��U�d�i�t����9�@
ƣ��h�5���9����:��8z���cj\����2�`�V���5Yx�N7�@2�`�V�����@;��cI�B��N��\��9���l��$�p��k�^�;{����԰��Wr������2h�%&����=�AA��ݮ���;^���m�qiĵ�������w��;��˗���E������:������=vEjZ FDR!���@�$J��	�Kƹ��w�`�σq@�R�fN��W��9��^n��ר��7
q�nnA��@2�`���WzM�#&(ˁ8/7`y�_V���ݰ��0�+csn��Q�\���PuG'�θ�o9�3�ř��*.d�e��}Xj�{/rP�$�"��>���o ��@2�`̶p&�8�e�k/6^d�*������T9T��3�MN���m�"�H�&��}�Ks|��0���գ��i�
H^lᴰ���^�0ޥ����\���D��g*�;���^%�GFZ�[��㛊P(̓�-i���9{��̓���0���CYy�r� y�_V�	��Q�$e@����^lՆ���wU��$@'2J�
�Gs}>;�Ʋ��7�4Z t �@3��>���LpӗJ��Ne�W����|��b��Fɶ�a뜼��0����Mq�g�L`P�����2��0���e��̽����^o����w��6��6�I�瞟W�C�ߠ܏���Z:��1�%�6�e�}�����rƼ5�{�H L�����Z_o �uᬼ�9Տ�A�↲�Z߸����=���s������N( �2�������T���?�TQ��_�g��_�����0C�c�dM�#"�D�H�?� �B DD`0X$�P��i d2 ��� 1 ĊH"�`�U�J!�H1�E	PRTr X"���,0"����b(Qb(� F �����`� � 6"�b�*HDa :�h@�"�TԿ��0���?o�TO ���:�����9�����%w�*��G� �����8��P`)���'�� �������(3O��/s��ޢ�������?�Py�\?��AA������Aμ�=�����'���5��@G�r�@@G���)���y�����Q0�I���ڄ�%����kç�TG����x #��S�_�O���0�^���:�[�?��#��?��V�������w۽D�?w�?䤇T�̲H���?��ٽ"��Kb�"�VE@d����$� XVI	$BDI $�	@�0DDD@Y��@����	d$@�!	 aI@�dRE���I���	�E �EF <�QEUY I$�	!	E$AaAP �Ad@FAU�P$�H@�B0�P!U	 $@FADg��"����$���"B
H22BH�H����"Ƞ H H�(��  B"�(H"B��0�DEcE�DX�� �B(0��B �E��E��(,Q*�DX�@Qb�E �X�"B$�DX�P�UX0EB0XE�$B T"�DXT"!E�QYB EDYT$$A R!BB
�b�B Ab�A�"H���0^��Nv���Cɻ�ٯA��C�����䠈��� (g�<����_
�;��I�]�ȶ��%��oaW�|����̽J" �=���`j�?�O�?���O��{
�������o����F��?�����������u T_{�
!&�|O��=���W��4ϕǥjQ�"�s�� A���������i�_��懇/�b���  ���Fxd���?�s� �4!y�蛡{?�@P� 6�A�S�x�&=C��<���a�Ҁ#����O�?��#��?�_���?eU����������+������?�������?��EO��?��� G�@?�_����@G�����8����;�o�����~߲0����X`���G!������?��_Ԟ��w���=��E��PT~�����?o؁W�xO�������@�R~����9�O��������ف������� (n�zD��Η����~�T���C�o�b�B�|=��rE8P�7b��