BZh91AY&SY�[��J߀px����0����a�      W�� (�� @ 4 ��@"�((  +� QE �  *@���    d(EB�@( (	P�(H� � �I@� *�J �P���B�I�!�     ��leM������F�-Ŷ�g{�;��O]�n�۟|�{_O}��7�D�[=G��twg���ӹ��k��{�r $73�s5���US�p�n�zs�ꇡ�۩T��ր�T��9�駽�����Ei�3�(��
�T��y�*%! �Q)P�2����u���|wZyt�˓u���7UU�UI{oz�]�{ڗ��^>����n��w�U}9꾜���׽�{���HQ�W���V��ʪ�G���Uͽ�W�g^Z���e�U�B��^�Uw���d�ū�n��&�}�(�|(BH�
IR ��wRM)���S�n�i\ڻerj�w�7ԯ��*�f��U��e\�|l>�u=���_=�UW��ݵ<��+�ξ�! �}�w�ɥ�{�ԫÏJK���-�e_y�%nΗ�w��.uU)�W;z�6�m95\���*��U(�� ��JQ*��HA+�iE=7�)Y>��{:�k�n�;��KqJ(�T������O�N��J�Ԧ�*���M��ꜚs�� ��-.{���/sꠣޔ�ڕw}ޟ6^MNg}��{w�"Y�Www�Sɯ�W}�/���W���J/R�*���*�(QG;�TP��)�>�}/�n��NM=�u*�RR���Svﶥ�ξl������t��z���J����w���H �����˽�O3�ޥ=碊�ޕ,۶U�9�w���nl�w��S�{�Kݟ=��Z���^��.              ���6T�$�    i��A%"��  4� '�JQ56�Dz ` &����T��*OP�  �h2b'�I6T�*�     �A
DJPD&����Q�	��4�O�'�?�����?��N���l>�����}����(��j�B((��@@U?��(��
 ��
��� 
*��r�u�J�u*������mA���i�����O�"�� � }����CR"�T��AC�O` N�=���U_aG����r@H ��!�T�,�@��!w �H��@9 ����<�>�T�S�QB {*	��H!�� �p '  y"�NBr@����rA9(�!D� '$���(�D�� A<�G�QO%!|��<�� rT� 䜔�p���!�'P�A���C����5;�9/$9����H��Ò����y#�y/$9<�� 9 ��O!�_%� 5yQ�#����r<�A�@� JrJ�K�y� �rC�}�ddO!|�J}�#���9"�����%9#��ܯ$����!�$�!Jr@�C��C����<���伇����!B'!}��U�C��_d��NA�9 rS�r����r^K�y	�C�y�^HrD�?II�(}�} B�)�}/#�%��������^@r������ �T�^��;��y#���S���<��9�9<�9	ԁ� �����Q�!�!CP��9
��=��!� >�(�*j�!@�伀伕y/ 9�C�@�� y�y/ 9�9	�y"r���/ �<�@��������	�rG��%9#���^I�/!NK���rPS����H�U��A9 )�@C�!�w)� JE� ��Q�(rDH!�Q9%W�"��NB'$��k�>�혞��N��n���WVf%j��QfeRl���l��E�f� ���:�Zΰ0Ә&y�Ws�x<�|��l�k78E�����)�&�aV`j
<��!�秞�����U��/+�����v�]pO`�7Ֆ̋�|����`|9�X�eTB&�a� ~	t��$O�=��d-�2����|��=���E3��YVX�a�A �!� <9��a��]�:#5��K�F�L���K�cp�%��R�����bWw�I�=4ڲ���`24iUI�R�Bf���$�&�!S���1[��X Y�]��&�C!QcV0h�3M!�!`����^SV�w �� �,�@�� ����V�0�K�f�����0�|c8P�c����	z�j��ѤyIXSp-<�b��O � d�V]���wh;��ı�v2AU7�1D��m�L�W�A�@�`]IӨn� ��0S[4D0�NM�f�pV��WEp]I�R@��!�QM� �L'Pg��SsB���2�ayG� �����H�@���`î�=H�L�#
�	�0c���W3����Y����g�aFI�/�Bd%	BP9&�iݭNe��@b��҃����B�ce��+	w�S�veA<�=p@Ah��7�IAD4)0Y��ذJt�Ih����gΣ��m�	G�)���AL<�V���&�"L0
�3��1��Q �2ה��҄�׾o/����$�N��F{���3���)i�F���}���� ���_��XHxX���M<��_�D=���n���Q��!|�E�N^;�4O��B,p,�� �3PL.��*���J�����BF�b�)�I�{�1��)��Y�5�❛�����bc���0hf����E"��,�5�9U�c��jZ{n��ޱk�f����OoFﱛ��[E�*�SA��71�
DU�2�y�0�x�(0��'-��+P�t�s�%�X	»/i��Xn�W�\�7E�Ad��ea�IS'_|�h�9�PLJ!�
s	�y�ewv�k���6���@Tb������0qR@�I��;���^�S�������|�wwX�WUxt���;�K]��R$t�l�����e�E��{ӛήs�6X�j�}~S��{�̡v��c��Xa�P]�[��m�!ڼr�xVz: �U �(&�M״nY)
A�HpA8]ٲ�6B������6l��#�'"OgCT�DD���ZQy���<�x|e�	�B��A��qE�+��!+gy��ɹ���B��f<�, �	�8�yy{ү9��<U�`��{|t�HZ�yEI^F�� �w5\�o�(q���Ɛes��$X!@� '/�	5&i�]�%�(+W�m�ڇ�8xo���V3|X���]�$�Zc,�y�Y�
@L"��X���+

,��(�C�����6����
s��֝uGy��2�S�#"h��p�91���`�G����ᾷH)g֧4lt�ƍ���+�����U�P,cE,�L�q�o�2/��h[�A���0R=tXd������@�]�owO`Ӟ*�wPn^\��	{ۅR�Of�߰&h@jX:�n@BX�]"n��ĺ$CH]�f[:� J�����$�8��樎��Bk(D�b�C�Ab�KS`�Y�NvPD�H���7�zb�bI��ц�zvo�T���	2<������.�d.�/k�3hYNJ��:�ҡ��]�3t7#�o��`<���
�&���U{�7�TNV2,�}&weሣ���ael�Uӻ��/�Y M�;��>�/���ݦ��p�#��͙�0��(�p�¡e\t	|��9��ŏ$~A�B4�2%���z���j���_F�����0$n!Yg�qj��J�<l��h*i�Q�i�8�w����}k]g�Ly���b��܇�hCý|�����8�Bzv�3}��@V,<}^%�g)���'M-sf��I�Pzy"\4hݭX'9+�����eGP"��F��7-����� !L�Q�6A�-$}��f�8�5�Ke�� ��1Ћ�Rb���'n$���������8�:��*ѝ�:��3YGY�g06A�����蜶�h�٬��w�7hg'0Ų�ü�5�U�4�!�����P���7��iE���xt,����4�r���z;���^ vq��&wn�0vΧr�1/rd�O �	��$D�Nd�&d+�j�4΂����B; \I�xcF�q˺VA��K:NRV,��Y����V��"@A@ֹcd͎XfȷQ�dak���0v���A����<�j֏)����sCA�4���S���Rł��#�Bt@aDܺ*Z
��6"#���跐<X�*.���e�yh�tW4�Q�d�*Qcc��Gh��0ǭw�!r��!	`��&&�. Itw N�N"�V�P�'xP��͇1��g٣��ww�ZG�Wy��J-��H��O$ӿm�7E1��[λ<��c��DF��3M ��;@2(Bt,�g��Aˊ�jd`����~�"sn\��J�V���zxV߱�	N�X mM	I Q!�[�,�����>z!�2Ɛ�"*	/��K�nA��tl���:MVh0Y����sl����w��oG���6��Y,���^��0��h4��d��M���+ج� ƫ�K6q�H�+zH��E���j��EQr�q@��:s*����$!�2A��J`d*tD���dv:�,ӆ�!�@�ϨJ��H6�e��h�33X�a �'@r8��!�M*Kz��	��{���_����n�~�lX�������J�(āҌ�i�a-C_�a	���,%D�!��@!�� AVh�)��^b<md��)HS��)J��>�8��hx�����V��/�n����˼�A-�}�f��� �=�T�w��ӡ�[��
i��"�,���v���kLM����~RN���Ѝf&l�$�f��-	l	*���5�w�'��1�
�l�	AA��dE���6�yc&P�yD�P"Q)�}�vo��Y3�4�Fy��͈+m�%�p/��� ��7���@:߈������c��34X5��1���������H%����� -3�X��|.�lӶV��Y7�I�`�~���,��C+�Y�!�:��u��A�Y��7M�� [�T{��Z���Z�Ļ��ʴ!G��	>�jgA�M;~!OD*AF1(�P.a���\�R8"pѤ�,�}EOg�;z0좉,�X7iI�&�����J�w��JJ�����fp�K=��b�� �pP%),*�P�@%^\cM���_	~�����C�q
C�����.�����Kr��(�|�!oz^h�#��p�1�}�}��A8�C�B�wN�� G4�״{���gYNQ*��sD�n�
��F��d%	A�n�;ߟ�~y7X��J*q�
��}��e ��吝OtE��:z����"X�٠kb m���f�k=/Մd/X�� �E.���ED�>�.*#��R&�Bs
b�T".��A�����65�0�S�7�u�r��}>w-{���g�P0���fH<u�tPu;��YѤ�QYoـ�sՄ��V �@pR���n�Bn�_x^۝Z3q�F�΄�6�z/`7�6�8i�wJO ��2���q�!S �bpA�4N�DAE�Ȼ����v=F^&DEDso�tia��wh��Z���W�x�8����2װ��$�����E;���8&������b��B�Ӵs1��80����D�1a%�w��,����eca�pA�F��V� D�R�m��F:�f�޵�gU0E.h����r �DP)b��(M�`���uE��.���s0et	��=n��Dh(q�)��0!Z����'�>���e�C��ƪڥ�Oا�M��$���|x��l�C`������  E�b���hZ
���/���sM܋�Y����ԯ�W�ZÜ�ȍ�j,���-�.A�� �.�B�o�B�5�7�,.��T��(��Kg�ҌD�#�L��N^CH�1��BʿQD.@�%jcF�(3}���y�dgS����2p�Ni#4ƴ�v�4���>�M���S�����g�]�^4#l]�K�r��]�&�$�������x���zq����|%������:ooZC96�%�A�����c.`��Y� |45A���靸��r�Rp;�zZ,�.���5|44�.6h�aW�o����(C@-��T��n]��IWJ�A�S *��6[=i�
{ڃk��+N�m���ь��i��8�6QN�; 'G0sA��ez��2tB�NQK5HR�E��h"�
� �K`����t!�@�`! &�b��@<)��!J���#;aOb,q�.��A�nf� �~D��8vl����'l��{ڑ��Â�����{��Еpfա)V�h*�t�(:�� "�� 5J�n�0oL�
�o֮��NU�n�!יf�*�+w]�ݢٕ��q�=����[�����
oJ�vQ}�ddw0 4�0sd��i�F|N>��hjk5a�P��SPB�,K~�gD^��5��wy&�]0��=A�1�,3)��tv!��>����#_�o���2ﳈ�t�؂��� ��+����鮸�j�X�@��K�7-�@�0�*��☻>)�F�eT0�Ʌ1b��j�@Ł��@@�:��� �`\������ܸ6�4M%24�R2Ocy��J��~�#B|��Bzm���rH!h�|������k7��/�$`!�A�'�l
-��f��������4���5`F�tS �E�0JPZ"�^`TIk[��o���X�8`oFHu����78z��݄���ڴm�܆d�i(ӌ�h3Z�Ѱ.a	�9w��h��@@1)x�Bl�<s�^㛺"ow]�C��a�U��x�x��!��!��6�
:Qg������1 �$�DULAtM߬�a�D�Y�E��^Bw�:��=�"��woϰ���p�a��������"��2��ʐ�4�b�41 +HTHb��5)e� B9̨8v��%���b �:pyC�	��� D�� %���PP<�h`'bE&R0��hk�8	*h�I7Г��/é0��輍f�]��˳�G^�5���Q�D�,�nS�*)�6�!�[��uYM�L�	�`�����Y��0�-���������df7��� �n�YQ�����<@�ˤ �7��hMt}D+]ح�>�-���^ݳ��r[&m�_�v��U���$�"�L*ʄX��k (0r�k�5_g�.�ˀ�
�掫��e�@��f��`<�H�D� ��h:�;^ǃ,J�E������-��A������"����U31-�6�a���p��73�2��¯���N0�8�w]
re��ù�%!�Ц�<4��ڸ��`��,�Sn�����}�;!,!���P�	2�[b�gp�q}n��z\�@b����%�t��j�Zt�Y!���v��OM<�9�X�#O$����(M����74Ptm�-�A�r�tA� �9�{�/���5��pX�`$�	2�P���X1eD#���W��,��>�<��ݿf�!�A��L�~M��ŕ�Z���=�l���V
�Dٻ�ĈF�8y�\�m8Ha:���xs�O@6������~|�9z68��_�i�q)��M����Rǚ�ge��F,U�S�D�i�_����p!,�Hp�MڵdY�-�T`=,�e�����ɚr�$}����檂��������������y������UPUUUUUUW7ULU]UUUUUV�UV��UR��T�VڥZ����������Z��������֪����V�T�EMUT�UUUj�UUU]UWR�UUUUU1UU�UQ��Ov�Gi��7��9�2�b*�N�ƭ��T[�����[g
�5An3�N�[�۰'W[uu�#�����g��t۞����u��̖��C��m�;]k5p:Ӝd�tC�u�������Z���M��n�F��T=!�v��m�)`��a��S�ή�7g��I�=�W<�X^����C��un٪�)���@]tƭQ�p���Ȉ����p�jM�W��k�S�����NZcf:���	�$m�./`:%,�[jW���Z�Wv�U��UR�T�ᷳ<�W,���uUW�UUT��*�����T���p4��W��l�9�Kl�UU�f���l۶������Z67���?nԋ���\o'Zx�rVz���6����6~v���mq����vz�A�;3�g�"`�t�(ú��+��kгh*�ml���L�����v�#��T�ڜ��.�vݺ@�t�A��ϙ檱MJN�9�{%����G`�l��1U��m�:�{�"fv�P�m�6�e^a488�U������Y4�@r9���Uk鯉�2g �9�.�UMoc[�6��VN�����2ٸ�+*�ֹ�T�G��Ua�4k�ۃ?E��\Y���U]-+��()k��r�!��\V,��)zb���K�����z��~q��5�v�:<V��T��IM�����(�\� ݝm�04ԝ�m�*��&9�+Wnq� �k�,�W[���X�/]�{.���5�v�2�F7�ܵꪭ��-���:l9���8�8!�0��n���l��>Z��1���ݵ�v���M�Oc}����r��An�Ub��:�����۷km�ˍ��%��B�ۄ�Z���W�(4k�@�a;h-Z���Pl!^WV�!�ywA��Z���v�M5�[>M,m����f�3�ѥ����y3Sy�v��{m���͆E�r�;q�7"���nkAbۮ�R�x;s�کT*�h4����kv:����l6� Z���2���g1�3�]/-ukVT/~}���x�ݫ��v�::�V_mM�E9��*5:Nj�i�zș�c���ԇkW-��͎����
�*�%�2g�+�
ꢝ��z��C�Ѵ�n:���7u�]#�҉��O)ѓ��^n��	v$淂_Hku��v!�Ñ�{S��.]������r�1��raR�P�*č�d1�nV,�ۋ4�z������Q�ѵQS�Sn�Fݶ�j7]1T\Ycz�S�,]�N�U���õ��5u��d�V�vɺ�+�@
��]�\���|�����jt�!���^��w��nx���}G������)���&�v�ҽ�ڞN�q	�iI{�՗!��:	L�`}�9�u*n�қ!ɇ�������t��m�Y�]�]]��^b����Ո��h��:�r�.7=�Z(y�7g8�6n�������b�ml帎�i�>
�j�8�S��8��㎞6�,�EWn����)���k�׆��$�)ˋ��k:Ԗ\6�V��Z�n�8�Uߖ�7�Um��q�,�ϊz�B�2�1òNիmUK��ppR.檝��ur9V������8���yw�d��]��ω��Zh�HUW;A�[-�qc���ݧ<�V����m���^x�)��ٷ6Ճ�b`;��Ԧ��;q.ɴ�S�=��=n�K�&ͣ�K/-T�U�v�UT�қ��>�[��R�F��$J��[\$�8v��u�i�!J�����D-˶e�U:"�ֶ�S�{v���CW.K�{g�c��˴��3s��U���n,ͬ΁X���u����ҽ�g�B�]�O[UR���a4��hz�7��UUJ��W���`�U:�bW m��7J��U���r�WbLEV�ջ	��Y�Z����<̵*�:�q���X����(1_�|�-Um��UVd�9�][���R`4���4۳��[f�.PfI}Um��0�,����u��\V�W2ʻӸ�0m���f^�&h*�J�d�+AUA�]b��pcj�Cmۜq�PkmU����v�v�X�&��mJ�(M��9�����b�J�VD��
�NԨ�"�]�W��A�v��G�meN]h�̪��Z�U[&-lه���UU�����M5P/!r+��RYA�+̮�����[ps����0n�ﾸ��;��粼��*<k�\�����[^>��mɚ��-���\��͍�*y��a�j�s�7*���f����5Y.,��V������;�
��Um��Vڭ��Rҭ[j��$A�ft�-�#���z��vNxmȄ�xN݇f�:��ꪪ�p�Wj�J�.Uev�mV���X��[f�	ýr���0;���j�u�V�j0]n�Z몪�3UP��j���-�:%L�wjU�AU�;��\�]VګlTq�4���'�z����V���]��[pj��j����	����\U����<��)�Ζ�����*����&��Z�٪�����"�Ãy-���Wm��-Z���Z�W�u�$�=O�lg���r��{�q����V'.:��u�UY����j�M�V�i�N�kl�AK-���+�UU%���,"Mm��U�`���	������\v�MT�Z��V�@q�^�l�֨*�n�^�����~���n�Ʋ�&��۶UZ�f�8�]<i2ZLʡT�:]�{��zf)�:�n�<��Ҡ�1�˓5�rV�\v��.M�:�rŵ�QUUK���<�O=Uֺ�M�݀ ���j���T-�����n�+	�-U��l�n9���K1PW]AUu\����i��n���U�˷'+�)ej����$�m��6�Ir���)��rkQM+�z��^���'5UQ�s�Ss�"�m��c�g��l��MUWUVͺ��������/,(.�r-AU��1�P���hq�X�nh+��8�Q;f��u���ָ]Ŋ�O����5���]pvݔU�xI�gV{UUXQe\��v�k��v�����]�)ky���ii���]I�=	l��	h�6݂�m�@҇KKV{f����5�y�n��:��՛cv�m���w\d+�gqCܣt0*��\+F6G�j��y��7D�Um�յn�"�m�����ǥU���`,�	��d˙f*�2�h�6�6vPMOYf+��7v�l��\��^@�U[��b$��.x���4���ǰ�n0j×}'ݻ�)�*��d����#���T��r�n�
㍹����Oddt�����Y]�CUlmr�s�� ��RݫjL�pP:��6>�_P�!xښvvp����)Lb��3l
�����ݵm�Sj�o0�Um��V���K�;��~z.�����nCc��|�/���el�E���v�@�u���U��-��ĵs<Z�jUȺ⛩m��kl*fXG*�9X�mq5��[9�9�C���4mul���ԩ���5:ؑ�U+^(���<�;c��x43�Խ������nN�/[m�d�onʄ��{#��:��]W2�QHdہ�˚��i���Zv�9�b܋:��p�P�\�+�45�U�0��ܒ��g�$�F�']s��W*�C��9�..LS�o�ګ�s%vƿG'G؁Wg�Gc,��Ld.���+�i�δ��G�	�D�@B�	/��m)���ڶ��G��_�u����RĮ[,ڸ8|�!=�3��j�x�G]�9���Y�;' �LOK�Ϩɻ��Φ�::�U�>U�ݬ�T;r۴��ۨR��ݹ�b�eYY�k�7S�;F�fֻ�r�*�8j�n�lm!��G<�XK�u�u�x���m�l��|��":;(UYU��V�UmPz��PyYNfZ��ٵ8l�l���� �UX#u�����~v2x����*�R�ڶ��;5���y�M������V���Z��ꪫ�R�UWUUT�����e3UիY�A�jU�^}����+tRP$���Unە�>��f_j��*j��S<�N�UV)��[�U ��%
BF�$Ma�"%]ؖ��Sh�����)�UmL��u�=�5UU*�J��UU�ۥvڂ�ڳ�D�ejݹ����Ut��K��ƕ�V�U��⪢�l�f��*��]+ͨ2GdTcZ�UG )�3��f��T�,+�*��rT���;O�V�l���.��H�jȲ�Rm�V�������*--�UmU[*m֥�9��J�ڨ��Ik��j-Sض�;as���.E���l� U[�,;sUU�-J��[��]�e^m����դ���GYZ���-:�����V��	��Clն�/��U�ŵU(&3��������U�r��Uճ�Et�USͶ�+7W[j�ͭ����=�n��6�IͫHJ��$5T�ApZ��qm���R���ͳ�j�G	Ckn)λɩ�*��g\�Լ݌��$��sqL�g.��`�/@rO)R-s�(*/[�l��+�z˪�d���vʆ�/A�="=�94�n�/19���l뮘����p�`�۰�>2r����K6�s����S�-%��v]���r���2l�֫g�뮱�8�܏=����i�vܹ»�M�A�6��m*ʵr��F��M���I�)e[ME�Bʂ`��\��fjm�l�����.͝uO,���]�_#�,g�>�Ϲ<�`�ꗮ��S����u��UR��\���ÕUx���U�inj���[j��j����6��Ƭ�u�)C%Um��������Knٶ�n�O-����o<�<���U�U�vt��o��S� ��mE�l�յ�*��;&&��t��f�@�m.�c����n��]l�+���8u:W��<�)ɳ�u�.ܕ��f���4�7�g�؃h����1�GTOl�pje�f��e�p�PT=���p��+��`"������b�?�'� ��|�ISS�H�Ƞc,��	�0$�L$O�"��4Ș�̬�
D*D A�w�����X�EZ��E�)d\b�E�)d\b�e�b�\�)e^1K*�YW�V���Ҽb�U1K*���DڵP�VTL��LK���)��;��Ԧ)��n����7R��w����;�[ݽe���?����/� �����+��h�%D0T�@: �H)�� h	S�_D1P�*'j���U�W p=A��О0*ti@|U�Qډ�Yb (�JE$�d��E���C����"z
|RB�I ��4���*�0	!(T�U>U6 ���GJh{}"� 
zP>�C�C��� {�D��}zvUKJD/�h&�CK�S�P� /��I�С��*�v�t��.
2��_ ��O�@��>Ԅ�D�� N�~e�<AqUvPETE+��="(��,�x |�򡂦.�� �@|TW�Q6�
�*�����N��I,a	L�2���3DQ@���0�� z i��C�����_�_�
��ʘ`��������(�������bH�j�"H���
$�&�H�h=%*�	=����|��t8;eĒ$��K f�$�)��F1*���b"��"f
#"0�*���@ث��uE*�0@'ʿ+���?|��X@ae�c�8VXY(d+&N�L����� v����t"R�@D�@{�DH��v*�D��U6����4"h@��=�t
���������������G��UEMUW��������s��?��� �2h��H�)��@�&��K���0A54�i�B�3 )�5��AcE�����ۍTq��a�XQ�H�WLi)rI"	Ddr^�wʿVG7j��UV�A�r�]V�NoD����ܵg��������p�E�#����&8�2��OȰ�3��;�bWRSp���km�V^T�A����K�>���󔘇b�펬����w/8u�t�p���8$6�����q��]q�;�"�m���6"����w�N��M�K��ä�<���,k��#F6�p���w���/|�ܺ�&Η��#�Jn�n��ەn�ŧ��b��˘��b���w�3nm��Wl��װ�Х�*��F�'mu��Gu���ӕ۴Y'�<����wg7.��X�����������h��i�d����4������=��k��Ep��WX^7�7���ŏ��g�ǵN��C�׈sn���.4�y�},��qwc�z�G���]r�z�+�T�:�pn-�
¥<)���vz�p.6@C��ӫ-��	��y�oS2풰�fY)A!D�"K�h3p�J��v`6�w�����t��=nͫ��z�[�d�W�#�dw�Ťm)�ݮ�z�� �%�&0�q-XTa�ZЍ���#x�X��rvc�Tp�k��0遹�,��v5F�E��3�6���+/�Td�[���1Ǵ�S=W\lcu�n9/6(�i�Z����<9P�z1�t�u�;7^n[,Nc����!Þ���@x9d��hݺ�-��ֲ�ls��@>�*�URt��h��3�y�RXM�	n	,���u��$��GX�z�g���H�<�C4/3��[*�knH�R/{�������v*�'M�̺WT�B�	�&�ϧ���N�B���Y@�Yz�W8�#���7��c�Iv^�k!F�@�#r�eG33���$,�Ȝ����*�Wk�<]a����=�7a��!<�vFX����s/����@ꎹ�κ�iǦ�e�+�li..w`h�V����u�� v�+�l�Sٺ�Z]G.��3#���}v2�b�QPF�E�@`�,�ktp��!ڬ4��V��y�u�[����8�n[0�E��JC/~��B�  *�H&	�P8�x	�B�@੡C�	򯀸��D6 h�X�5�D�=�k�k���H��B9��#�;�Lr�c?}���|a���mݼ��ϑWџ�{��l�^^wl��
��p����r�\�I�v��<g�A�HI��'GG�mD�(ّ���j#!�a;y�{1��:l�m�V�E��Ơ��[`^��@{)��u��NL��h�<�}������^���Iip�y7<�s��S�T}r��:�����޷�l@��z�U���2��<��|�]3�)t�^|"'5�0HH�R�*D!�?yY'�r��[��
��Ż���]fʒHD9l�+N�X�j�N�X�j�ۨ�-:L�)�Cq���;����+���"�@�U$��m�u,���<KR�#ګ��[��**��J������<�%��j��Z�C∝A���8�3�[Yy��4��5])ۧ^�.Q��ȗ�{E���m���0n.z��MOM�#ګ��+�^�SdoOmH ��nB�i9c��� �4W�T(:a��r�����໔�p�<��AB�U =@W
� ��}�lv��w{�ZwŃ�A�P����u�]�7��fn�7ٳ���,	��i���ɯ��ݞ�����{{ޱ�C�R)rETUYW>!m%���xB���o�)��"!���]O�&���Mtx{6�m������Iخ�s����k�<�Dq�)���Z��*��֝�{R��JS�ҥ��⩅ueL)�MH�7���ܽ{}�]o����+�V�5����#hnIu�[��b�ν Z�d�H�V���T��� ���g{�N��"DH��V��Uqn������G��L���]T�^G��qjK#vR���,��q�l]���ĥvtl���a���{C�g����b�Q����k�<��G]M]qjK#vR�-I`xIW=�Jj@.[h�7L�$���b�UW+���n�x��^���w!�f7�5#H�$Bo{�8������o!l�<��"�3EIquS,4S�4���������!t�&� �Q�J�S�.�OA�3�����!�&��q׷���yW���>�0�<3W7������4م�$�:.y�
�K�A8yS\رɵړ^�zsRid�	���K��U��x��������������J��H�U�\Ͻ�u��^�{�;W��<w���7D4��t�Uĵ,�)O5jY���R]Qd͖]]]C�r9�	��7e��K#ǒ�{��"�.� ���zR�jԳ��I���˩ʮ�<<LV� 82D��O�X����u�\�l�[�[����|���^jz�c�if�sC��M�R8���&�[L���%<uE՘��ۦ�����U��ݫ� ���\r[�)sCveB��А���+a��[R����=J���]*(X���"s9�UOn�.;�֋nݻ����6yӽ�H����e�\�@kt�j�ʁ�7!�
�P�-(H@�$ʐ��HBF�m8o.zu�q�ʱ_��w��qo���$EΞ���(dN8�.Ioo�XӾ��{�7W�����dZl���I�w���D�o#v[�jԲ7aT��ˢ�q��~��Խ�\=���;�ux;��D Ôd)%���*�w�cN�λ���{��Y-�$)�qW{��w�u��z����|(P�~�|����%Azĝ��r��.��6� l�n����b�ld�:h�PP$���� ��=�λ��L݋��� �o�}`o�M|,��@c�:�wM�j��D�� �.�H����Z�b�-�F��`��X6V�EX�SD��D�DT`h�[S[�b0CF������`d�ӊd�o{os�AUPB�
|}��Vo���;�:����4ah`%���[�����뇻�Ç_��D�6T�!�
 ���q�u��w03����E��Q��E�,i�y�{�9��{���{��H�B(�2$�t�G���Z:����m.�qg�wW��j� " ����W{�9��Gw�u��J��4P,9E�ҎƝ��ow�u�ޕ���X�#�q���
���kz}�߾���~ٷ"��T�G�(B��a��[�y��Q1�ف�Zr�w�+�9�����=�8[(X�F!NI+���w:��zƝ]�Ƚ⸜$I�;\Tv�M��ےri�IED�9c4l��&B&���i�d���η���=���pY�τM�1�Ѫ����R������û�ε�D(i�L&�M�w��G��g;�ow�u�<B�Z�Jq�:�{���μ�߾�ڑ�k��PeA�^{���G�Qp4���}�_
]���{�= ��+;x�Q���1��d��ޮ<z���v�0�jy;a�r7^�FVN�L�-���GR9n��cN��o��Y��Z8�⼒&&� XNXӽ�{���ʷ{ް7ܼ�4���
rI[�t����i�Ig=�W��E  �,���2X�^����i��<��^!Ϣm��1��r8�w�����}��w*@Pʥ%�r�S�RU��Z�[��Yz�>�qմۈɛl��H�B.���M��;#�v60�G+��prW&�Tk�`rguy���m�_��>v��%��Q8�n�ݳ�޸�ϝ�}W�,v2���S�h'�w$ż��;�.�	�94I{Z܇`�Q�V��� �Ne�K,um4vdٵ��r����I��;���z�eM��jݸ=�Wi�Ÿ�^A�[�� UЪUT�*;&Cp�CU�^f�vv����v���{O��;�C�ur�ئ �3bH�a0�nh�^�V����U�����|��&J���n*�{��]ʷ{ޱ��ʯ�r>h�Xr������*��z���*�{���w;���n1���Y�~��;�u���ܫF\Q>�؂KrƝ�:��/����o��}s�z�n�^n��I��0u����`&+hxBݸ�L`�R�>�r��M��[k߷���;>�����Ds��v<ju���`ɫy�f�y��w�{�x��CJ�U���v0�y�w��9�D4و�h����ޱ�}�{���U��S/�DdI��-�cu.���ż�w�����nQ%�q��������U���xy��U�@x������I�R��9�c]���&���㒸N�u/@vvK�ű5�F�9�(4\��mG��/|����w������a*4ӌH��ow�U=�{���^�����y/�&��Ӗ4��u��AC�?��I$AI$�I$����Ͻ���vz���o���bh`����!��(��^���z��a��P�@�@�,�+�9�Z���!�;����s
�8k*�A�2�g)�ii�(���R�X�d�	�mCN�, B��Д	�P�2����׬*�0X!���;`�944��a�+nꟲU�+Fy�Of �`�7�7q�����Pd����n�l$BLQUY�,:���@bT�JSs�_ iRmP (B�3@�u�m�]��'Y�&��]P/<i��`ap��!4 ��tɫ=hTNU��$������t�W�2kĀlb#]`ڛ�n.��
0@�p��d��`����X<��k�u���V�	$��Xđ��x{��H҅%���~��JJK0Ţ�]f��K4H�$�5.ܘ���-�[0ҕBG�[2�${t�yr�Ly�<�vS��h�@�h�(�3�ݞ���~E��z@>T4P��Cz�bFI�	��A��~dt���t����S�{����O�%7�^�Δ�*��=�:�i�<���3,�fNH��#��MP$W��ґ٪���o]	�%(y��s��R��*��o���JR��~�k�o2��y�f��,뭏r�����gJR�>��9��@�>{���)@���}��R��3�ϋZ>&b���p�H䶸�nJ��|C��ն����ں�:��:�9Bi�n�}�py)=��s��R���}��JR��s�����Jߵ��hO�{�V�oX�4�m�,V�MP�~�]P$
$W���R��~k߳�)Js�s;�i?#J_r��kl[��������JR��=�6=JR���~Δ�){Ü�{��<�~�R�����e�e��5�Vlη����R���}��'%(y�s�p4�����JP���r������$јD�@`�1r�Q�(��$z�?�<�5��y�Xj� W�G��-�$ur�5@����s��R���&>�����sh�f�����2�a�!(�AD�'u$�Z8�l۬m�eֺ��j���P�,��.�9��n+5����)�{�5д��s�R��~{��JR���s��{��o�C�Q�����[��MP&�~�������~�)J�}���J�+���|�b\�srh�� n�c|��}l{��=��u�yJR{��·�C����Ҕ/<��y=�R���^��rD��r��
�+7sn��S�u�gJR�?s�lz��<�ߺ�T	��}�_Tf$�eێ]��T����3�(?	'?~�ǹJS�~�])JR{�߳�r����ጙ(a�*DI�B��Y�^��GZ��\�[b���շ��II;f[��v�#���Mͷ�-���-��tk�e�x�5ۮ�٣��禘�<�f�:�[b]-��a�cqJ:a]i��]�q�\�Mi��>t�;#���8�^�ˇ�7t����e乺ӧ��J����ۣ��y�r�1����޼nz8�j�s���� C0�
��K�q���	m�GA	��@�T+�T��<1��|�I�^��J��ݣf�Y�v�-���vN�^#h�/CY�e��y`Ƶt��[����P~��ǩJS�5��ҝf)I��~�C�)����Ҕ�'|9�4fj�kn�f��[�ǹJS�u�3�)JO~���{��<�_s:R��~�>��)Jw�{��P��BGQG���P&�w���aR���}��Jh
_y϶�E)IY�<n�T	��ǐ>_2bm!�o���������JR��9��`�C��=�_g@Ҕ���9��)JG��C��P����BH�T	��}�*�4�E�����JR�߿~���)����MP&�����h��Ē,<���n��7��p"�J4=r)��+��Ťn�]�Sٗ�aE�ce��r�5@�����t�)I�>�:�)O3߹���˒�>����)O=��syZ֫[��̵��y�4���:��#��S���;��s���R�Ny�6=�ҝ����S�*�ZR�����k�o�h�e��Cܥ�}���JR�Ͼ�cԇђ�{���R����s�r��/!��6 j1Q�\��P$
$V��lz��;�^��)JR{�s�r��ٮ��R9�WγQ���r�w:��=�P�^{���)JQ����]r�����JR��s�lz��?*��_h�vӄ�m�w4���8�Ws��%7c&�ܛ��R�Ru7�:�V7���)JO��ߺ�)O3߹���)~�>��)Jw��:R�����侄 Ђf9v+P&�j�|���s�R��~k߳�iJO~���p�Y(���>D��II#��]P:�2^�϶=JP=��~Β���>���fcG�Fj���4��4M�X8E&�sDAZ�a3�bqP=��w�����R���}�:*��{4{D�#c|����Nr��O=��Δ�);��s��R���}��JR������9!��͟k��kZ�o{������JR�?y�ܺ�)O=�9�)JP�9϶=JR�y�~Δ�)�T*� �G�>���j���i�c��1Uf5�Q��5qvָ�u����e�<=g9��nTq&�m��
�T	�{���P$
0��c�)����)h~����9]a�@�j�x��D+jH%
H(y�}lz��<�^��@�����Cܥ)���Mf)C��>��`�Q�v%�a�����j�4>��s��R��=�5Ҕ9϶=JF�o������(�P�㋰
F�C�o��{��<�y�t�)K�s�R��x|�HY���5�@t���ŹߞgJP��6I�+?Y_͖k2�n7���=�R��߿k�)J<���6=�R�����)JR}���Cܥ)� k������ی4kdZ�F�N�*�gg8�9�����6��3�h��N8Ź����U�֬���:��z�JR������)Jy��:R����s��R��=�7���P$Ww�/�E�ce����5@�����3�?�I�95�ߎ��JS����t�)O&��=I�0u)�����ҧ$B$���r�����\��Q���J�߹��R���_|��T	�������n�R]��J����J_`��Ϻ�cԥ)ߚ����'>�����)J}����:����o[�t�)K�y�ǩJC�/���gJD�'>���CܾA�����JR��#�ăM*�1,@�"14�ĕQE�����֧3{�fVf�Ĭ��p���ƫi�Ӻ{uvMn.6�WǞ��䅺�z�T����q:����+��h3m�xt�<'k,��XTf'ͦ�ݶHU48���!.K���:��+g�ݒ�~闾|�<ݲ�70�.T��z�9�p]a�P�-E�tlL�b�u]��&:8R��৴qqW-��n�!Ǭ�ɯO3��g�a�_X�#B�����A]�n$�!Qn%��Gcq�J���a����2��m�ky�������0���l�F���<��?��~�t�)I���:�)O=�9� R����m�j�5C|G��"��(�WT	���s\�{���=�9��d�/>���)O<׿gJ�d�X�&r�9�Y�e����f���=�QB{��~Δ�)S��cԍ)����JR���9�s�9A�Qϴ�P4F&��Q�|��Uϴ�/5�lz��=�_s:R��2��9��)A���k���݄S���U��LF�u���Zj� Wy��Ҕ��s��{��7k�s]JR���lz��>��Ϩ�Ίޭo[��Z�<ޗN��2��V�\Yu=>;:�Z������B�\�Q*q�R�+�(*����t=�R�g��R��>�ﶛ��BhY�ݝ�u@��Mw�P�5I��o5��Cܥ)�{�k�?�? >��e�.TQ�������{@�s`m3H|ەu�Q���Q�����t���<���6=JR��_�Δ�)9�s�p�)����f����fkQ���Ҕ��}��R���{�t�	�I�s��{���,����j�43G�G��0����%����Ҕ�9�s��R���s�Ҕ' rs��=JR���3���ݼن����t�)I�9�:�(�����߳�iKX���l{��;���]P&�+;���M�SF��`�6;<^g8�݇���-kZ�f8Ү��Q�{���$��jD�b��hB+z}򺢔������R���w�ҁJP��n�s�9A�Q_iY�6�Cl�q����R��9�Ǩ �<���t�)I��p�Cܥ)��3��G hs﹭sv�LH�u`ܸ+PĨx�����P%Js�s��C���@�FH��H@�Ie� J"ު�䦹���:R�������)N���N�� ㈢��P&�H�w�_X�*R�{�s:R�����cԥ*y��r����{7*��I��6���:q)O=�9�.��J:`C�s�p4�������)>��s��R��9���\��sN�nX�����m�1]�<Uu�\0�˸:��w{���ݵ��l�MgJR�'>���)O<׿o]JR}���I�	�)�k�gJR���s�~	�$j@���a����+�C��&{�9��)@����J����U���F�oy=E"d0 �S{Δ�)>��s��R���}��)�
������lz��=�_s:R��o�y�AK�Fi���T	���k�)J}϶�w�P�{��:R��#��6�c��5hg'D'�.
�����7��{��)AÞ�[���%SQ�|�9A\�܃ԥ�!S�w�����)9�?~�{��<Ͼ�R���C�Y�7�-���%��綝ʬ7�]�`y�1i��=��+E��n4e�B��i؍6�R2�Y�pVHr2�γ�(O>���{��<�y�t >˒�?k�m��R���w���$8�(�$WT	���{�V�iO3�s])JP��>��)Jy��B�����_|�PD�-��i�,{��<�\�t�)k�9�ǸU�d�~k߳�)JN��g:�)O~��3:�Z1ٙ�F���JR�P 2p�͏P4����gJR��}��t=�P~U�~���Ҕ�'��_��o[գ3f��[�ǸS�u�3�)J?
��Ϲ��C�)�����JR��s퍚�MPu�i$�H$�E"�A$�������6��ۍ��4|g}����F���k;֯,
[&�����'E�T[��\-�0�S:�+[�q��/p,��LL�Q3%�*4o-Sp$��4��G(^H#�I���q�Db�FL��fT�TDE=�g~=�[�f���uXk��U(�[\@E�u�K+�5fe�a���DQ	0E��o����F��֨!2�(�ɐ�	�0vy�CD�LDxk}��d`�MX��BEeHUM�jt[
�r �X�j, F� ��o�8h�-�l��[�E���Pź���K��`Q���0�[i��`�qʒ<	t^3��Ջ�v�{:���E�6^�ACf��tdg��rc�X�+	#AB��C&�!�գ&�������ao9 uҞF`��:���h� @���zMv�6��UQ[�5��đX0����P�Q�OoB �PdP� U)A12QіY`e��AdadAY�u��4Z�AG  z��=��9�^��74�'�\C|��Ф�(p�A�R��bSR �q�! z�溳D��#)���&lL߆PU�|ﮮ�UH��׊�f"<�!Z�b���$1��j�[j�9�EHUWUT��M�m�k5o]�u���+����ٱٴ�M��kv�;B���/\�HV���d7[;F�A'��6���a.Γ���m�p;#�����H��=G9�g�k�;f����^K]��%���u�g�g��^'[���	�s�V�����V��Y��t�ZB4۵�.ks���\�WR�Z�v�դ�cK���kk�kcz�s��Q�ls��Er�P/J����-b:��yD��1��p�f۷�����Wf��H&.i!�h4钭�-��L.��9��bA�bg�������۔gmg�h��Z:.����p^�a�s�w%ZZ��P=�܇c�g;�ٳոbl���i/<�P.������l���K�\yyg��Y͵\cy��a�#�����~۵���^�8al�=]iU����a�ib׃L�+v�	���'�6�ͣ63��N�v����]]t�v�,Y2��x��y��榫��m1���I��N:����$�뉚�v����mi1��x���][p��Ӯ�=e!ŞgP6��vj:^�S��QM�0��=���g��^��I���kp1[�m��l���鋵8Ƿ!Nڝ�~�6�޵�J�[�n����J���k�=m�ŷ����j�k�dl���ջL�&�)�h89޻n<ʛ�Xӛ±��Q�S�b��rm-s�[u��)���|\	��$`�4Y�7/�c���3���5^��[6ɶ���p�2]�1��N��nf�p�_-ح��s>�c�U���
ݼk���^��'�Mv�t�Bm�\��f-�xٸ��N�M���Kc���Px�q�]��7�N�)g����=�ûvM�z\�rjiw��m��3nu�1�Q�ym���U~-s�5;mr��l�O4t�w]�Qo8��nz78b�q���n���K��vlnkh��rvt�x�:Yh͡4��kcv,	k1���p�*r[h�A�m�sPP��F0��j�4���������]�a��y����i��i��i��i��i��i���kjB����
���:4��/�Q� �j���"����F =�Ü2��M�̓���!{bz*���e�Ňː%���v܉�r=�t9<nG���L���*�����.uq����}�����_���ݺ���TleNbLm[$��w5-�+�Ŵ�ًE��~����*ѓ��v<۝%䖮�۝����|ۆ|�nI��nn�`���Iq˭ώ�]s��7$�A���I�F������\���(l�u�h�k[���ja�R
��B��
� ��-v�����5�[@�t�Űw7Bi�(C�Oq�#�k(j���~�o��q�Eۮ����9�r������ND��� krW+�~~�`}�c���5��4��@��s�Ӝ�H7���Np�}���_iY�H�B��q���
�ۖ}Z���D�94��::��8Υ��l#-�b�˘M�oO|�����G���9�j���֩�\]ҧ)ė�ݮ�����@�+�y��w�ߝ�t���{E6!�E!�v�[�����OY�fV�7mdD蚎9�M�>j 9�K|�qD
Tctӗ�>^�v�5X}Z��r9�������0>�&'! ؁�Q�d�^���`T� e(S���	�6-!�8�A���bL�B,�� ��u��uW~{��}��{�k��2���iRh�1�R����ndخ��&�ӑ��[�Jj�j���0L��I�XUUp�f�z�ۮ�Ż���"8�w{�_s:���{�#��ј�C��|���`%UUU����}��+�33w��7a����P����!@\OU�Ճk\m4k��f燑���n���C�w��}�E	��8�q�Q���gR���.��o>�DDD�r<������?E�ۡH��e˓�+�y�꫔�������`����9���|r�S��qȬ�w����	�|��?@V�P
��ʮUC����Ǹ����=)�J�Pn�s��UW*��UQ�o�
�����z�N��G%/�`����&*n*j(��� Kj��r;���@j[�@���{%īcE#%&)��SV�=&n.����@uWKv��nk�1���2}�u)!:W.I�=皬�����u�Uy�
�����ةc�:%
"+����7S}�����[�m^��V(�2}����©L���$��wX �W�Ȉ�ޭS�j����xՆ��(�p|j8�?W9\9ʮ#7�ê�}��Ϊ���������E� % '�pD�'�!����� ���K��锑#�.�@��j�>�r"b9�k}�e}�`9��Z쁰}n�d�DP�sɃ�!6]�v�^�u��.�;*㶇�Ue;4��;��������C�s�:���1L�J�@��u�	5rG"#�{�5XQ��y�9@J���4�zӭ�}����(���7i9���>�UW+��n�W��iӉ��fnI��j���r8��G@��t� ��&��QJI�.��w��9̬{�3ٻށ�n�#��M^�L*Ș
��H��Ȭ�n��~��s�s��~����ޭS��Ds��,<���f*��%bή|�u��kW�wB��v�fumVM�Z�=s�3�aR��W �{�1@�䛢��v�cbx��@���S<��oN�M�5�5ׄ���KHqchX�6zs�(�5��h]2����-j�n�.�,箞�a;[Z�f�ƭ��nm���*�����nM�W(r��N�@�"�H�EQ�n�T�ϝqC�!�:"��ܴ/�?}�:�Z�m����'J�;���ul����80q��y;�z9h֎b��grۇ5�t[�0�R|ܮW(��`GM8����<�� i��=��9��9 �7� ��Xj(B$��' ��%�
���8I���O(��s���\�B$c|��΁~��]�����W8}�zX��>_b�
��JTIT�I��r Z��@��fq�� �9���Vi�ku�R�A�6��z}��?��G"b"9���@ݤ� _<������Ȳ���;q�摅Ԯ�7#����HzM���d���vն��gvi������}�eʉ�$���KwrX��VD�ٻ�W*��ei`z��ؒt���t�-�د}��ο��E�sZ\D;P7Z��>�ސ���0��?s��O9?������NB5�Ex������nK�Dm^��r �B��L]X�H�jN�
�r���,srYE����a�W(�w�(�$j�QBJ�9�ل �W��Z� Z��@�k�`���|������^�i<��/���&�6x�����&(f�����α<�~�w�o���wu�{�偳�� (��tkx�s� �ܖb��yD�*%A*�K�jo�9�@{]� j�z�M󜪪7���j IƠ���A��z:��=�}_�:QL Q@D@��U5
�,u���C��Q~��y�^fy�s��W�EσVI�q�#��@Q#�}�d�Z� Z��{2Dr#���0F��DȤ&����0����Y&�P�=����36��7w%�G��,�9*GGM[�:��{w\t֓��Xq�b���.�7����^.Q�`Ӧ�QB8���w��ݸ�ڴDs��v�N@�)!�AEL���n����9 m��=��+ �����9�UUT�����(Q19�\��9���w�{Ԕ�""�Ͻ 7۷V��R��IJ>Y.�KK�\�}�9�U��s��W��W�qw�!�*���!���^y�����)�7�����n����x�Ԕ����?����V��Z�u���<&m��5h��%箫��^��g�����n��;��|�Ͼ�׍Q5y��� m��=��9�s�I�z��Z�����j�r��7w%�{��uW9Ϲ�u{�tu��L��~��	4!II!��ܞ�7����M��r"��F 4����B+"j�r��R+
�r��n���ݺ���`}��+�1aEm�0�H����̞��dG"%5x�Z� ���꯹ˮUW��Z�J��6�M�����N�ruG+�/Y���4�6|h�l���'3p�=�p�keȞ6�
����qe���˺�0a�9-T񓮮#�9�͂�Cgks!K���(��<y1òGd�t����~�?|��<hۤ�<S�M[��՘�w��Fq����;O�O����V��;[X��u��,��Ls����7��XR�On�:�@�C��d�?_V� ~L��!M)"� �0��A	q�7u1�˸�p��8I��u�=�s��bO��w��>�%9�q�V�̖�?b�3��{�UW@�۷V��E���nR��fe��Ns�����=��`M^��YX�ظ����Ȭ������F9�6���j���=�uq1r9Ƞ����ʪ�>�n�] V���=�[�:+�*��g9�߻��\����%4�
�r��w%�UʮW�5�vfn��W�ɥ��U}��q�%H�SX��rE�y:L����s�,y�5��n۬FRiԎ1$�5I�֮N��<�`-M��{]�9�G9���P��5D�!fA"�}�}����T����T,0�Ϝ�-��'�6����WF#��-��K.͆��ٞ�0L(������]bC@�6� ⃯UU�.��0=���j����" B����JE4��@��4�5�J���T�������9��u�Q�/�x��NF��p� ��KX����|�ʮs���4����G��t����^e�2wm9�r9Ȏ��tk�`Pn�K���*�FID9	���sO�u�\W]S�Z�Wc?l!iL�a�a$�A�*�[r�#B�$"#�XQ���w�}휺��9����
�wE����_s�҈�*r���I��x٥���=��8I���s����G9��N@O�eRHp�O��祒w_y+j	߱�$�H$�D��I �����y{� |� ��	���@�1��(<�բ���Ο<6g\<
d*$"�4CKr�!�Jȸ��Yo^��ƈ���3V��� #ނ��2�#F�P@s�"�:!�ڔͅU�O
 �LQ	�;��l0h�)"AD�wcҢ�
��s5'��&�	����fa��][��Ψ
cT��,5�y�P��3E�z�,�0�B��!� ���TH�Q4-�R2{��/s;0t���S�&-1��~�	����mN�ɍ�:튂�A�a�Դ�J����
Y�����$P�u*B9e7dzk��0��h2f��:�:�FoZL!""����!�#;Ӣ47V�=1QD�&F��� "���3�[��[4����A���6I������@mN�G�E��M�����/b'�_�D�=6�h|N�;�n�g��x�#ʪ����߶i`̯%�	�(�5�9w�9�DDjW.p�}��l� ���`W���N馁�S��R+$�z9��=�ـ�Y��j�7���p���*45)Q!@�E]�0uV�S��\�&��B��%NqeP�H\��%8P�i9}�l��7w%�����_���*^�ﺣ��2���oz�W5f 6���V��&%$�z�lȡT$�{��	B�J@���e��A�i� �o�>��#�DG9&��� >��x˹�j��$��+$ *���ϳ*�o�U\�>�����P�!(MpUQU�q�j�=�k�F��q4��Nw��&��s����`V|ױ���ށ�ʪ����Tq����'MAJ�s�x��R���YE���Gv.��t�`����w6�w{���thr���HX�߶U��	/�y��#�G��`��P为��.
�ʜ��i9�$�z��`�����W*������lT�)�Q�'	���_w�y�f)��� 5x��N z�1 ��'SJ����r�+�U�|c$��x��Ne%�w�\��CH�!rS��28]������p�s�ݼs��}�}ށ歘���s���A��Mì��Iu����l�<nX�x�9�'#m�-���gZ닮Tۘ��(n�9[y�zĎM��98Ld�n^�3nX�����Ԫ@=n�lnz�x3Y��E��[<u�N���
�-1&T6-�κ���G-	7[�W-��׈�Y9v
n�j�&�	n���
A�H� Q�d����+��(ɚru�̋k���ِ�?�P    �d�JTs��dx
nֶ��G��.)�L�v�v��]V��UUq+���(��,W��/�:��q��[0S#��|�5
R�B�;37{Ҫ�A���Xm^��U��r=�K&&��I�6�I��nm��7w%�\�W��`ff�z���芚��:Qʺ �����U�y)o�9i�`g+Q9�J"}j��R1{5�+�[��t4�08�W�/
��5�\�C��^�Z���\�i��E�!��l蓊��v
��q	�4�u�*G`���i�`M_"#�ϵV���Mْ�!��a$h��X��~� �W
!DcB8�J��f,�7[�	>��C�����W���k���׽�}[�Ф*�UP�U�nnJ�6}��d��A:��@�O# #u1ؔF�E9t]�Э��s�[3T�����8�U{=,^�,#c���.(�.����z�y 5xϽ��ݪҪ�InҦ�C��S�D��-�w���޷����af}�;i5������x�+H� PM�����6��7w%�����*�Tfn����0֗C�T�I��\`[W�l�TV2$�΁�FW9� z�V��'(�۶I]����u}��s���Q;�aH�B�jb�F���W�C��Ͽ~�� ��e�����SU�9$��-bK�t�Ԝd`m��s��j� �f0�:���Q
K�{v��+��rn�mj��I��kۙ�	�y�ڋ��D�E�%c�<n��U�wN��y�7E4�a�Q� 	"S��H)*�7wo =�W�Z����9���# #w?/�J18��,�'@��k�UUs�S�O�u�� m;� ��E�q:���$����oz�ݺ�*�Us���n��?b�3|$�Měi�����9����d9:���V������L���9��~��@#E������'Q�VZF�vXW9U���1X��{�>�۫
7�<b�U�
�H�h$t��aN얖t�Hfv֡��륫:���1��{��J)Eԅ'(�۷'@�j�3��ށ�G��#�}�>_}x ��sW�&��)�"�3�����s����+�͟������'��N>r"r#�!�n���j��*&�z�w�k��l�;瘬3ٷ�z���	N6��%Xr�\z���Jp��zG"y�6��`�7�MN:S�2����}�uX���i?��� ���?>Do3�"9�1K*�0�&T�`�,*b	
�J�W¸��xr����6��Xx��+�:�v&ղ�Ͷ�/j�ɞl�vzxH8컁��p�Ȍ��uQ�,<�m۷f��3^���~�۾���}�mnC�>�V;]�/]�8v�.���Sj�1���Wv�6��� ���o:�vg����^�n�{��q+exV:�h��ݞ��Q*ar��J�m)\��N�\�ۺ;s��3����TQ)P�� ��>�1ƂXbM��]��9FW6�v'n7��33h⦔��6�d�́0��B�ܵf)N8dp�d�+$w�̤��5xU%�y4��$�L�w�fM%��b[�f�RS�-��9�p<��謂f�⨚��� z��T��u>����9�{VQ�����QKv��5��W�i�ڟz�l��9��G"s�����`{tZ����)�"�=����U� n���8���*䚂&ܻ1��|��Ӷܽ��q�nm͹�z,q��H�j;��+$t\M!���:�Iu�3�4�4��T���DG;�G$o���7Q���R�gp����y_���s�DG"=�9���׾��>Z�zJّ��=��[MJt��2������V -I�O܎DL��� >}x ��l�I(�)�$V����ޔ�4���ޠ�+�b��wȭKe%(q��h&��E� �"""[���t��������f�c�#J��t�\���c��kA;�����N�n��Vp����k�ɹƛr�D����e�Ob��f��g�i`z��(�I"D*}v���I�DG �>���`@CM�U\��#�&*�C��\H�fo{��~�.���> �R������C�S@�Ʉ E�d�S@S@Oy�����k��7`}���>�+N�%'zr"�f 6�y��N -I�@+��F�J:F3�8X�첂�ʮ��8ve%��j�VI���s�%_>����b���2���j��]K�����v��n;v������}o��З'��]��M� �'ހ�[2 n���Y8�"#
rGX���r��:�DE;�� ��� �S��d�3Q��4F44��@�d��svY��¹�qk�V������I�|I�br]ف�4���Z� Z��C�`�)�he`dBI��UW9�w����X׿/�kB
p84�ۗ�<�9�S�9�G9I���4�� 77e���1�P�rn��
'����.m��]�s^�dh��p����mC��9������ޟ%�&���9U���~�V�f:5*���T�D��@Z��Ȉ� CM��Z� Z��~��s͇��@��JMq� ����dUj�r#�I}ހ�[0V�w5#�
��%��>ܚXQ�����XUs����+>Œ&���$
r+� Z��}���w��� �р| ��4�I$I"PI$�*���v�����02�(�#�+2'��4ff`YdE�a�½(.@U׆��ݙ�K�����C����w0dQ���3�7>�1�ĭ���������� h��u	�Ew�6��Ѭ�c��{4[������[��&k���&�A�(�F�HĚ_��6�DHF`Q���2�Y�ʐ��h�[#7�-kZ�Z";��!��(ߘ���q���Y��>�9��`���A����z�f
Y1a�sm�iњq���&����M��5D��,�3���h"AiA�� �]�(m8�"��!�:�[4�Ģ�\���7q$�e��(A�?��I$r�ն��ds`�����b�KU�m�L�ņ�p����L��/U��Hw��6]��%�9��1�76����;iU�[CF�W6����Vkv�WW��s��H��6{\�m��]��R�'z���t=0����rޞ5(������2�V{=��Ȯ�%�u����\�D��joY����Z�U�w�{���k��杸��6:���)yLc��1�m�
<�v�&�E���7kh�68����;�{77]�.��!�aۖw��{�"��R�x��x��6�{c��v��^y��R
�Ɯ�{D��`�#n[yh���8�������ʡ��O:����E��x��у�略�1�y 9��:�.�!���{@I�Q��CC)�;Ud4Q��䁀݃�v^���n�=��W�8�*-a-�v���Y���%#�7\s�1�]Oc�,��K��umU�Đ��R�{V�R^9�l�s���������n4>8��]f����Ȍ,���6�8�7j�o2�O�+\��g�dז���PM�v��9���t���y8���u�;;��&:�wN�!9�e��痛�����dw�6���׬7v)-��/t��L�5��35�{5��GUEGa�qV����ժA�tL�LΗ��fxq�lM��Ny��[�c�$e�<�Om��t��J�签�m���N]ѽU�57�ܕ����O���)�W\��98�{r��(	Jf 7b�ڤ��ga�]��5���=��^v7	A��9U��i�Ӻ�oq���S���<��Y��%��I����uY�����{\郗��b����m�E��u���E�r�S�Y�ӗv��<�t��V�\=;��5�v� q\�ͯ9��T�ڇ/=��}j0��n�3N���j�F:%z�׫;7������*;��Ң�k��O9��v�yg�q�n���q�l�x�u�����Py�4].�un�ȇ�������N?�����00�	�mXAT����j����@��ҁ(���x�v��W���Q�Љ�CN�?�`����E�$p��CkvEqtr�ش��Iz������,�ˢ6c�c�v�)r�VϚ{Z���g���e�5ܕ'k�v��V�[��x�iS��t�ϵ��s�JsNuL>ҷjd�gr�۴�4G<�b8�;<a7/Z�ݜO8��\y�g��@C���VC�LV(4�bD�LD�q�RI����aM��.R�7��1�=^{Gf����zP�8�lo_� PT(PD�`�&�I-�a���b����eu��%�!rtqխԙ�0]vԧ�w����N���bLR_�}��K �ݖwժ􈈎�r"Ho�����A75�q6'Q�]-#w�,���1X��Ӻ���tu��L�����k,7�ՠ�����@�O��I��f|�������X��4�9Hr����U�Y�>��Τ�0:��#���� �:5*��T2%'zP}��V��,����'@����@=�Z&' �:p��uv�'p��7��gcG\S��f�աisՄ�/jK�s��]�YA��&��ʰ��d)��R]����ށ�O# 9ȍZ�D�S��(eܕ�>^�w��\�(�p���7�&�xY�s�}��߿tuF�nn� �رĩ�r) 29#�3ٛށ�O#��H�w�zu*��ډ'�bLRw�W��۫ ��ۮ���k��8nnok�fn�I��8�&�qsW ۼnc��j����Hj���3ر=�)0�	Jr:aR��5�(GCқ�1�Z�`ĽqR�����nmq��"�*k2��zu:��u'ށ��?G*���7��`{M��ĝN9L�e�{R�����rd������� ��UeW ���_� R
5C�%'zٛue^��o���6�4�D��%r��#��ϼ���X��>�d$�i�JRj���p+3rX/f;+����@�lҬ���Jpi�R#+/*�Ħ� 9I<�����Y����U�T+��(��I:Yy�%Н�q�+�t�(X���۵�^�<�����E�J9��@������ݺ����9΁��t��F6����R�b��k��r2" !6� �ԫ ԓ�t74Bb�*���ҎU�f��g=����LDO\7�z����65ʁ�:T$�\�����)k���no��uy�9��O���X{?lpH�)��q�-i����Zq�"��k{�&���ʲb�[`JI�h7WY�N�d:�]l��̬�	�͚M�@Pa	��oy�a��F�H�6I8F�S�4(1^���e�to��S%1(�2]d��z{S�t����j���_��>ŻEg1: �S��5r]i.�ӫ���ݙ{=��6�X�D���۫��ݛ��(������0�[΁���$�g�s~��W9��4�%)�'*}�xs���U�����<��������FUڹ:�3]��{7�+�fmՀ}���=�%�7QI�G%�����{SȜ�<ۼ��ګ 73)�4�JhS�29}�f�X��l���~�Uy��s������~Ώ~����G�iRj�9��M�l�ݠGlB���Ǥ��cuױ�29'iN�p�k[���n��99B*Oq�z^��]���V�Nɺ�3���:wDYQ��k��R��H���Y�!�"�Mm�){#ծ:��c3+κv�8̽��K�������C��2c�G��Q[l�>:o��.��]����x]��'�F]���+`�c-�ܐ'h"���%�v��k�m[ݣg���K�]��	�&��fm�{,;�c���l�<À�\��kF }_^\���Y o���� ����XX|��j�~�)2"��mI:�3]��I��y+fM�}�O9"��dc�I��'L�;ۻ���ɥ�UI��^Ņ��{J鶁�n�����0&� ��U�s��N�����#T��1�B�7}��#��ɏ �I��F�l��X�@�f.*��4#���^��u�v�v^͚��mq���hn�V1~o�P��F�ʹnN�T|�u��7�(=�4� fn� ��'���E)J"�8쓾����xR���P� ���V�.�� =��q�vu*�܎D�����n(�r�5)&);҃j�Xf찂;�d�����
7sZCQ�P���8���<�o� ����I}ށ���`�Ł��&��6t�%t�f� �ؓΐ�N�n��^6���]�0#��u����|�� T+� �,m�=�mg�Ն��!�%)���nSJ�rXff�u�S�쀵��0��7��"�MEqU���ٮ�W9T�f��,�͖���ހW�8��%)&��ʯ~�7�W~�������#��0+(Ȃ��!b�����*��\"21Y	F":��9�DG9����΁����&C|���H:q���b����vX�f���3]��W),���,�3��ԔID)�W�/f~�@�<�aA�ݖP�d��7i,Ѻi0D��Q�M�.7h�r�}�]Ɗ�r�[�sD��7 �����]!��}@b�k�f��2X{3{��*J�TBJ6�q���0�J�jO�u[~�G9Ro���>���2�l�W����`}����n�ـ�x�J��*&�����M����Hj�`M���}@DB�@dQ5Tʪ�p��͖I��|G�M�
j �����Jـ~�DO����w�Wٙ��炷{��m�	��U(���3֖�ˎ9㱙������٭���<v�7QEݝ�&���%x�P�ٓK �ن�����)˖�����fO%��R�`Lw��SJf`�J AH�=����Խ�X�Xw��a�����P� �(LRw�jV� I���W��G9�p����P�ʭP�El�B�T�ٲ��})^��t�l�?(�F� �s�p"FZe��dP�a��
F	� �@�>��U��|=�n�bk-�^ݓ!���I�켥��������q��hDHن���g:Ӱ�.��@5�Z�.y"we9ov��Fu���G�l'(���N�7�-�$�vI�͘[�{]n-�J�A<�91s�N�F��5W%�^�ma��o��B�@�n;\+�7"�m�q��Ƚ�l0=J�v̎�FTF���ܛ�L�m9z�a�r6
I�!]P��P)�h��M�Y�v�r�ۭ3.�	>\��kw���EKQ�0�jB��������$�zv�WY��U�.l	V]]0�.�u]�g���g�PH�ߓ��Ԅ�~���%�^�+�JJm20j�n��7]� R۬ �(�설�z^�*Zp��!�)�������}��ـ�]��W��ˮ�{[�RN��5+f ����/�-��Q�Cou�v۞y�@69�"ѩ�9�mџ�x'�YE�Z�ω�0L]��@^I���l��y�f�;��e(s�rSb��(=��_w���)v�~>G�+_�������K"Y���@�ͤ���B!i�*r��� ;�����#ڞF���l���m�v����,�f��{۷Vܤ�o������N�BcR�˫����{�'��#���ݎ�/���;�d�6���`~������JF�T�9��xdd�&�yG�,o1��bT]��{Iյ)4�j(��:H���V�ݖ�2~�W+�33w��s3U/�	)NR˫� �x@G�9>M�@֟���<��}�a�a"t�r�:�n��w������U=�QI"QE$J	$�K?s��~����+J=x%�Ö�]����2P�k=��ލ�٥�@"� ��!eN,Hбq��j�P���!B�����=���X��6���n�'t�&"޵w�f�1&��km��a�6��a�gz�ٌ���� ��,�� �:��:�߹�@�8V$F�Ɓ�@��E6] @;r��H�\��b
GA�������Na6XYct�5�1�v9ӹ֚���j6J�dŅA�����!+�K΄�Ԕ�Fu��j��t	#5��30�b"Bk04&S���q@j4,�6���@ف�|�:��f��)�9�6��n�Cy�ٌL�̜l�j�3�X8� A �TUZ���&
*�LV>��@� ����"̈́�7���wǻ}��I��{�l{������ ��Rh���#�'��Ƕ���S՝u�]o:4tlٻ{&zg���!��:Cl2��Dh�A�A	�l��4h ن�0�/O�P �����B ��b� ����/�iU���A��e��P���!⇊	��~����9������U{�o�}�$�ldtF ��a_�s��^���tM���[� �x^����WqqT\T�z��7��w����`}��ށ��+j:t�j��!B�Ӝ9]b�Y�I�g��[^�/��'�E�̱�l��Q��9V��,�=�fK�������ۅ�en�5D$9(�j��@n��rd������0&� ���*lr�S��,�3{�>��Ձ�vX~�d�31b����Q�73wށ�O"r@I��{U�~q��|�A2IM(�S,�(�Ҡ��!љ�?{�Ty�0��Y�ʫ]�U� -n���x��ށ�[u`}�#h�6�:IU)�N��qێ��x��a� �$ݜ��m׵��~��[�B�.&�s�} jw�j���=��bH5�`u|���6��I,�O��=��`i�2wگ?DDG�F��ϟ��s�D6G;�=���w6X~�K{6t��Ė��T��(�e�E�ܙ�����;�-_w�{S������M�I@��N�A�ۖ	jq� =��`@6������CeUH����k �5R#�Q"H�� bL4�!�)�4�F"dPTTJUL�5TR�&��v6�&��I�e�n�1O�s�9� QB�.�.�	�k��׷A�W6��W3���Y�=����-�m�t�J#�]�����C3���g�b��x�#0�kW���m1>[/�&�(���-�N���=���bWYv�89�o>�*��,j�ڀy�T���u�=��N�7Xl:Nwnr���zz���7B���i� ����e@\�"�+� ��ؙ�>tgr����ŭh:1Y�n�כ�$>�W���-'M�EP*7&߽���>��Հn���r�]@}��`n�Z�RC�Jq6T���z�<�I/]��:� K^���� �"bQn7*�7��aA�j�>�"bZ_}ށ��0�P�]܈�D����N�^��_u?n��}�۫���,
�ycy"CDb��8�V�o�{�����7x�Z� � ���߱�r�+�k���Z��t&��s۵����tڪek����<[D0�7�l)w}��78 ޻�L���?Ds�����z�_��t��(ӑ)"��No����d��)�dt
`赥`r0�30�aM8�"�t�k�u����M� Gc\��P��I-�u:��U�����/n�
��`w���Bl��
q8�?s�-���t���� Kj�z�N@�K��H8��Iށ���?Ur)_�E;����K�ށ�"�uϦ]����N��އ<O=g.ݣLm�E�tݮ������뒎:m��[��yY�������j�(_>����l��� �{t�FF�*�;}��櫠33w����`j��`|�X�26'R����M��zu:��y�O89��r<L�p��FO�_v�T����!�J�D���(���]�Z�q����V}����%Z�dNJ�6�B���b��G9V����w�zR�t�yb{P�JD
!E)�RCtu S���3��]u����i�&�t�^W�;��[���C�����Ifn�@��םA��;�f*v��䊠8�V4�&��2l�u�L��x�j���26�Z�I8�G65���1n�v���X�n��_{�PEN�@�n���m�΁�Z� I7ނ�?~���̳>p23 �s ̒04��f�1�`E�ZG��?=�'�[�z���ߵTaQB0��Gs�}�5XP�o�ғ� M��>�9��DoD�'���Ӹ��a�%t�Kw^Qe��"M��}�����wk�΁:��M�NF�J�d�E�>�����қ+6�0�j�<Բ0Ӕ	D��@�f밠�ܖ�y����f�k��cf�J�ڤ�j &���ݛ�ֻ���m�
bu�gR4F�)�F�tc�U`{ٻޖ��n����%����N�
T9N(
)s�n���6Su�ڼ�IN�TG��㻿o����h�W2Lg��c����*���k���P�[��tٴ[���1=��懷�Y'/S�*��l
49�xs"����m,T�-�	��8�wlXT\�[[+b�e�p�-����l��tv�$�}\%����#*lxI�;#z��8��;M�(M�O/i]�-�\�u���N�m��]\����xث��4#م�ɬ񽤣��w��|V���=v�&�r)��:za�L&���(s�}��
m�;���6ka%����n���� ��� [W�{i)��u7ހW��V���Fq��v^��]ޤ� �M�:�n�;�nb� ����v��(=�uY�f�z�n�
��f%�7��IҔ����r�Ȉ�M��t/��6��BOm�U�{uV��n��$�D���F/n� �7y�&�%8:�~� ��Gj��*h10��g]�껛O7q��˚�'5��q��m$r�P��g��-:ف�Զ� }}���=�����t���@����f�Y����;����G�k�ο��^�1؎����������� �F����r�"�"�=���@���g�3�����=�V������dP�$�t��`��0 �RS�n��ӳ0D{ؕjR�j�6Ԏ�3��`_�阺%���l�u�}�>8�&���fn��2��It��v���ƶI�y�z����9)��EWH���7���x����A���@���[W�vO*�DԦ	Ґ���`{՛��W��]��}����դ}����c��LJ';��� �mV�"9���L9�\�'9%�<>M��ϙη���������ҮH�TԤ�v�Ȉ�+��=�����ށ��� gզ�n��iS�o�����vg�{�1{5�Q廎��z�Sv��:F��{�����y<\�7[��F�vC��Su-��
��"�!')!E"�=���@��k�=K}����1X�ŏD����n��:ΧY�Dr&E?/� ��s�o���s�ă���~��D�rG`b��V�RS�o�Ͻ6u��ﵐ�	H��.��5���=���@����Q:{m F�d�a8����T�U|�:�9ʪ�����j��')�t�2�nN�_>��n�u�p�����~�ɹu��+�O,l#Vv"�I֚�2�le��N�!�2�� Փ�9�D�rw�Ek�ۮ���ڬ��瘮��ٻށ��ZS�H*jRm�#�=�ڬ�%8�7ށ�۬ �z��3E�T�LW'�s��� �&��6[u�{_�Xa�T�HNRB�E`{���@���jp�5[s�&)u��S�FP�)$��͛E��{�ė�y��^��9�u�(�(Pپ��YffVa�$J	$�I~}����h9@���Ҩ ���q����)f����X���,��-�󬏊I�������*4Yt�vhI�ٙ�kIMgf�04��}.�g�P`�w]��=	yMߺ>�l����jGC�?(M��#��������s�Б������(6�H�TA���	�(a�	��'���ui]6F���a�I��&�|�Ⱥ��,��Ŋ�l
��Mj�Y9��m� �[ʖ��"�!���0�f`BAL�N��p�Ţ�032:��)/^����BO4�-����l=߿��rg�>fA�M�1�e�^���2��>5�փXi6]o�
�̣K�M�d�'��fk�3:4}���o�ADX�Q�䓁T�c	�X%�c��!�7F���I����y��$e�q��4U7��+m�+Ұ5�Rb��h�T{�AV���;p:;���<���7�;��c]��Ѐ�/4���E�۰x�t_������$r�f쌲 �1z�_��Pw.�5�{�vP4��}����[{�]��YdZ��6�4��cX0�L�P!:��@�,B��]�ew݋�,B� � !2U		�s��V�&��FU�@�i�]S �F�k�$I�,,!=�P,*�A7�`'�ۣo��$��� ���(�U|�'9�m��XM��%�+xv��{KaNѝha�]��E�K�UY��mVGg@�Z�U^�֪ꭵZu�9��n�w�;%]�8Z콮�Gu�sݔzr���f˽��+�1��L��9U]ÝZ����:�s��9�7=m�NԽ]����x��k�9h]e.�黐]��W���.t��ff�\kmF��|����eyr�i84>Gq�8M�=quk��t\I���W�5�#�NSooO�t��uv���v��0=u4�V{H���m�'p��g�z���
nw]W��s6���˸6ƺ��4�m�.��^{vN*F3==�����K=u�����wS(�`A��O(n�#��g:����vk��wU��f{���c�]��Mk��s�<pe�'v��ze�xd�ūm�{���]s��砃��^.,�qs�yVV4�=e�p�/(�Y��)��[j���hl���)��hCNW�夋*��i��T�+�m�v2�~��_��Q��BQ=�Y�f�β�WDB�w-���m�_���Y,aq`ҽ'k��bj,�6���ը��'b�wMԧD�c��;�tY�R�b�nl���^�U����N����
�id�ָ� ���C�%��>R�ϘR0l�<�m�T��v)����*�l��Mi0N��u�e�4]>�lc#���ۇvvv���y��v9<�&^焱�ġ�� yja{����qO)�u{)��mr�k�����]Z�ۭ�L=qp$�YM�u= 2��v3j6�E�[�y|�y{j�a�#�v+�$ɫ�n��'V�ڸm2S�W�5`֞)�q�5ܚ1�$�S�t�f���ݨ]�:�&�\D�u�k��dL�+"�涎ߩ런�{j���lhy�Q�2;pc���d����Zs�\�x�7c1��8^�<�ʛG�vL\fe4������n�8p��{^��v�uH�@�(��9`^)�w3������(2�%�hv]=�y��%.c��=mwm9��\�b���5���n��憠�`�l�k6oZ�÷��8*x�h��
 ���
� �(A��pt�����h*��}D���y�6a҃-a�t��{3��]��q�ɾ�OAu���j�p2r�T���~r��d�d��^���d9�!����ck�N3��W�L�vy���؃��҂�/�̖���s���KF�g��3Ղ`,�ջ��^��\]#J�m���;���9��c�;VC�u>��0v��Naݣl�듴ڏf[�-����s��=��h�^V-Z1��"HE��U
�T(9d��i�6Z�7-���n���5�@�vD���N�V��=�������aۿp����N�������ȃ�'��vHO
� (� o��k���
=���@�n�X׸��<�,X���C�S$n�.dK[�@M<�]58@n�S�5��m	��"s�#wn�k�n���1X�n��f`���8������0 �MN�DF�NzO��<�i`~�9Y����T�%�*k����#۰nw=��n^N���QY�N�vm�<�Q'6ڧ����+����
�6i�����j��p3U;��M�TiF���������`�>��{���~�U���VZ_y�����J�	�鸥�z�Mwl�]58d϶+T�	k}^��Ԫ��A!���`W��+=��p��z��`@G9���Awq14EY=TRs��o���,(���}�הӤ��l�M����tp2�a͝��Y���r���crbxX��Hu#����Y�/f��@�6i`{^���+�@�<�bK����Q%$�@TT�5}�N��jpmj�Rs���cG$� �Ci�*�#�{��^�g�����l>� ��!7�,s���zo�g��<������t\YEQ%r{Y=���N�ӀJ_}���y���K�����*�qX��z��Ft���Jp�b���d�eM��t=*r��t�\�,��p�A�S�	��.\�(Ap�p����B�U�8e�Xv����V�o� �Ƶ6�%B�����q��s��z��M� ����T��}��`r!(��v���U��f�z���w��|�`� �2�n+����ٙT��-����ه�O9�/]f����~�IԠ��G;�=�5X�q���Vu/fo{:�q���:h�ynwC^MSN�D�ά:�Z!z3�<Y.T��Q��ɻd5-5������`\�m)���7�����bd�r(8�>[v�y�����7{�=�4�1n��Ϸ��(O��qH���������� �RQ8��F��� �(��b��u`b��`o�)��9�O���t��MĐTL�D�uq�)mM`�Jp��z��Ŀ�~�{�W�
$���*l8��9�:�]=Y֣aҼŶ�
�s͸�8{nް�O�ź�/'gt]��٠!����2vՎC��x�[�������4�&�Rw��~˹��U��p;sWN�5��6���N���;r�/#\��^�M�Ś��ۃ����U�ޒ�N�j���kk	lpm�=jiQ;
ͫZ�s�3��us�]6�]3�1�_�o�}4�?-��[�%�8��{i���B3V<'Z��)E�v���?�}��Z�����.e�_���7ކN���;-��6OJX��I�	
q��fn��{2i`b��`w�1_��$~���Q RtJ	Q��@M���)mV���� ԛ�@K��j(m&ӎU��w����Z�5&�R� o���wwQWEV^O@�� ԛ�@ԭ�d�t��'�
�KG��e@܂!E6�h���רPݽ���f\@/)v�WW8����C�m�rs���9��f����̚X�qX��V�=��R���MҎI�t�~�|���BII@��%@0�0�0�3�@@4�϶ *��CK�w�Z'~}�m{{���I��4C��I�9Vk���y��խ��jO# ��M� \��L����Ѓʛ�� M'���䭘
|�b�<��cMJQ5@�n+�����ۅ������b�;���F�DԵz��ú�ZM�F���N��>Gpk�C�̚�s�#uR*$�M�DA�@�f�,�\��JpZ�z �&YSu`F�m8�X�ڬ�K�1X�n��{3n���զ�*Ich�ۍ����Uw���}�4~��J�B��T@�0��M� (b�`�%��c�Rv�qvt�;���+��;M�)��R� �Z�z�l�<��=ʛ�F��*���*n�nw�{3n�k���;瘬}��ށ��樔e@IF�v�:�̄���wI[inK��S�[t�w;^�
���ʔ�L�U��~�`g�t� �&�� �̌ ��[�.nj��d��˞��M�z&M�� I�`O����q�:)�rF�>�ٽ��� �Z� ��R�ꑻ�0EE�DH����:��zX����y���9U�ms��Uד��|�D�mG Q��Wv`/]`��Jp�o��[0���=㍑��$HA�T��B��B��U�);��vӏWd���s89Η��j��Yu�<�9�7ɾ�*NDs��I?R�{V��M�Q)r'�����yRs�l�u�v�N@�*seEU̥M�H�z��U���gR^~�`{}�{�}�ֺHj�"�������;��p�M��ySs�����X��!��;~�ǚ�f��c�W@yn�?��g����*�Ug���ɶ�\<�mY9]��wI�����q٩�����uNc��Cs�����=���U4��õ`��N��К,u<�m�ඳ6#C]x(��gl\�F�G\��XL'=�үeV�v/�η]Zb6v��<vl�o:<ɧ>7u��9�>>9�$�˲׮}���m��L�P9���{^K<֘���v��ܶu�DMz���w����z�{���v��7U�(�)mF��Y�(���Z�\l߻=�|�u��7tݝ�:���ʫ��]��O��K������ �MO��r��=�5X�~@>AӐI9��T����=��p����-D�*�n �i���{����ج{7{�>Ǻ�>�գU���>+v��Np��]�T��vv���n�����qX�n��}�uX[�������M�*66�B������S���R^yt��y�	�۵���`���۠`�V�	����QM�H�zٳK�w����X����j�W�kX�&J��٭�y�fs�k����T�i� IaM/����﹮w�UϿn�uP}�4�꤃ٟ��J$���N沺u�ӄ�o�� ��� �f(�h�nS$Ry~�USy���_��mV�V���HTY1n!""7;�=�4�>[��������ܮVlH�M:gꃒ��&�4[e�Z��'�v��E�.�=d���$�y+ch�F�#i�����v�Ʌ��g��@�l��3��Zʎ�"%1�۷�5Ss�n���2'V� �mV�	LN6�:%1�5"�=���@�=�g�|t��"��$�!	^�����:��T�AE�DK��ee����YaUFfEQ&2��c�N�hzx^&��;�ώ|""�kz֜�b��G�͢�2vu0AL�3QW��ִE��h��}Q���i:萀���C�3�Z�f��Ffv6���jѪc:��;�}&�J�En�@�B�(�4�X7l�6�։s�2�1�rZ&7��;�ޫF�10vNS�	�
4�k:W^�;ٹ3�Hh��,H��S5��&b��'�#�FDδP�.G{�NF������c�������/��F�3�X�V1.��~[�N��YaFI�$M��b3t�*�����f�Q`�* �i)-ق��&��`�K�%�d�h�]��a����C{��F�Z5�g}��8*>����D�T��qӠ6�v�' �ED:�4"B�3�����s�?�f��V�� �A�huT&GCI��>�{�����`|�f+��������T&JE(7��ڬ�IN���M��M� ��A߱���7A];�=��ע�X���u[��/��)�<�=v�e���ݵq�����S�`���N����DvAO�:��n�#�(Nr4�`{��{���r�3~��O�:�=�р|�|��&��d�.&��S�`-��=�рn���30�v�EHĚm��k��e������߹������$I���s1� �9� �F�8غ02�&���4;����ݤ|��p�>q2㚢���d�ճ �#�?���O�0k�V|��V7N�@�
P�m� ��r��}�qs�l�.�r<v��۳Mӆ�8�<��	Lc�8X�n�����k�Vٓ��dt�QP�G;�o#>�DDȾ�����_� �O��9U\H+s���P�mԧE()*?/�� �V�9��92������#2G�,�	GIIE&�n�@����ｻށ��ue��y����I�|�JB�ݘw[�@I������Z0��/Ɗba��!� ��_�����]��I�\��ve�R펮��=*қ�68����\F]�[v��\pu��'/7f�c��h��������0�X�v���b��[�Y�[��۟nieشU+�vON��t�[��@���7Wlcs�6���1�3b��g�v^>����n�r.�9!k��'��ӭ+sӮM��sb��yx�-I�hQ��y��1����߷��q���s�ƐP{K�Z�lt5�=� �c��4�ք�1�6"$r����0�G��Q��?��# �� �W�;��z��*������*�>Ś��&}^��@�ݺ�=�����ț%1�u��ݲ0�ޙ2�y������ƛR��$p���r�Kٛ���Ձ�=�`}�V�=��I�QQ��z$�F�M���S�@�@���)�1�F����8�'Y�%�vz
���s������ɷ�07g*��n�*np#�%h�=��~��E����F ~��l
m8M2�.��۳K�U�o9�r#��r`}���w�y��78�{1IQ��A������ށ�y�ZԽ�j�>�&�x��R���sSu}�~�s��Kv��]}��Jр{�����(J��NJ64�(�)��z�#�{u>�@J��ބ�0�\n��ri&yrK�y�\ۧ���W�r
.�����n(Bj	
ޫr-����0I>����<�� ���-����@���o{��UU�l[_}8��� �V�q�&D�:���*K�,�.��������0���.AR��$̕TUu�$�~�^�߻���~����Q��*�n�*('��Ur߷�n�0�����RX�8�c�&�*j�&�ns�x��;f�������>ܚX�����[M=@�T�M1)\����m���l)b/��9y@>n�)
�R�S�
P�8t�o��c�VۓK�d�����F�D(�QIށ����"""dK���5;f {�}��9^l��BU���$N��ƜVg���=�р{u}]�\�� [��Ls5EXPE�n���%?�� I��z�Nr����Pq����M�LE���2N�l�7�~�:���[c:�n%"�>�?o{@{j�<��v|������q��Q�F��c��&�̄���z�tɲ�ڮ�N,H`� M�*@
��;�=�4�2�������0-o� �뙂��	��&�j�O��v���[�@�푀�٦|i��ӻq�̛�������G9H���0;�Օ2�J�� �I§�%���}�{�=�4�1}��?r��fM�`~�k����%D�Ds�[�`DDro�W@J���~}�����Q����!V$�࿊��L5U��]`8H���%�С�ty��]z�ag���o-ѣ�}��}�|!�D�y��c�
nX^g]Gj��fZۋ])8n�Ḷ�w'97 ���l�&\�mun&^P�/;�!�����j{%�7&�k/s��76:�á���5A�3��!�\W&Q���:$�H�=�ѧr�����)�7*ʕ���vMs8�P"m�Ǥ� tۮ�����ak�n{޽����wq�v���/e�1�:zz��wnH���.�by��\r������D�!����GQSbn�|���y�+�����r�����~,�����h��®�>��79�9ɓ_���}�|`
|�`�,*�IХSq)��nozu/n�,�Z�-���J�}��c[N�au7}�n�N �u�ݤ�����Wۈ��M�JC�$�`b��=�J}�	M��nـ(�.���`us�`�C����Uv�uu2%�b'�:Ě����FS�%�pD|I�E7i���vp&�z��0:�� {e*�*nဤ�'�{~���� �(<�}��܌��`��?s��&Oͺ�n웅*6��������;-/fL,�w{�Ve6������5�,U%8��zs�����v2 ݏ��V�84Ԧ��t
�{�����zn�Ձ�y���\�9Ϟc�rT� �m��=vv��zA�vѶ�z�Qks��ٞKǭ�Q�t�t�eD�I�9T܉��3��߻�3wn�k�]��{`fl�(�J�U�z�q`yV��حs���z��@
�T)D���y���?�ί���!%,RʐK$ww��Gy��{��ھ���9vIn�NP2�V�t׺�nn��f��\K����q{��V/�A�	)%' �� ߓ}�r"!��ݎ��Ss�j���g�+�ۢ8���u�L�h�J�mps�[Þ�rk�%3��f�!��bz2��n�]6�Q��If��]���`f<ŝA����P��s���r�N�JlNJ�=��' J���z�zM�g��Dr&E����%C�MJaO��.��?ߕ�������V����䰫m*M�ʦ�e^N�}����_]�=߹Ȏn�� �?*�����_�Ni?���#P��)E�Wބ���u�S�$���a'x�}QH҆ ����Jq���0QBs�]���۞�#�-�Ix]�ڃ�`v��D���`t��	+F�'߹��X/߿]XP{��~�#Bj!��t�7M�)�#o��m�`t���2j��rqGI)8��V~��ށ��u`w_�X�1X�c�(jTB�I)/���0 �S�%J��>�kr�jNS�Jhn)VuױX��pz�zi�d��N�@ 9��Y�9�����P�<�$�C���D�-5���Ơ����f�z�u�xF�2�*36堩%&B-�FMMS�",H�r1�*|33Y��3Z���xr��]		��A�@@��c�yz�0�+
�3CA���i�44%Da$�E��An١� �= �Z
K����V1�a�-�lB�A��Q�B"���X '%U����gy�ԽF1IDD��2P���k�����;��4:�*jF)�b�b�H(� �B ��ZII��L��;$5��C[�' <� � �EhT��2���/� Ihf�W��du,M��@xZ�&�FcPaP3,:es2�Z,�!ݨ=���ca��7~��N�f��ϵU�����J�<TA�i~�̳���0<=�:ma��Ņ�8tEl��1`�
A�j��p�7���$����I`� �Y�&`��ffF�j:���u�`m�*���	(H&D� �" "�
Vb����N�"  ��E0�F]Z����'m��}EdFN�3��5���n�:k�3�"���H`����{�EQKP�1Y���^py��q���筵�Un�.���QT]H5AuU]UA��4�U�Ԯ��[N�͟gL��J��6wF��xd�Ez�H5�s�ܸo#
��)�bm����#�7*����+�u)���ԛ�a�n������p�dx�Y����־��d-Z�V�"�lg7s�m�Kڵ�==�v��*l�<��ΰ�uk�g�n��'M�Lxz8᧮.^w7!�\��V͍ÿ�.>o�X��F��������jzGG �I�돘��۟��ȑ�Fΰ�t���V�2==r��k����i�XAw��*)�:�s���1�;�98���1�/r��n6S���=g�<�귋sT������-K�2�k�Nz��n��:�n�y�^�U��7�;P��nOf;v�]�o,f.�̐�%,�P�];��\a<�v�.N���k�3�q�W�E(B��8-�M)l㱝�[I��M�jUT����.}��9Cs
�3��\γ� 6$��}h��ɺ�N6�h2��'m��@邦��{]<-!\���F�4Y�RS�o*�Hz,ړ�}�M,[�Z*��]]÷c,l�ma�N���y����A���8�y�N���/F�U٦��;3���fŹfUֵ�����֩�t�:�ҭ�����n͘�9��Um�ι�=vwmb�x�m�S��CӞ%:�IV�<	nӼ��ncB��
��56��!v��X3[Z�em����<DW��]�u�fM]'m����6�]��M��뫧��훨��$=�:9ڻ{Z�;T�bs��;uRK���R���Z�8f<\\[J�l�z�>c�j��q6�lL	�����2m2"�mʸ��@�4k��ͫE*��"h�v��X��E5�Mc��ꊹ�I�<glYCG7:ۇڠ4Zr����y6鵫m�V���U]ƦNռ�*�����G=���	���
;H�uե�I��AڻY�^��\IJ�Ԣ�R�g�d�!��,�m��KO*V�Kv�p��vNH�xI��K䙇�N�œ�tu�c���H!���H&�uy-�*/��O��(p?%�Ch��  Q8�h�(T�(W�C��24��1�[���9䬜��[�kG��\F���A.Ys��Nwn�:kXp6�����ȕw�l�<�\g�����⎍���Nc�V�lH�����
����v�.sb9T*�J�u;9����ۖ�A�ŰXli�y�9�z�+�ہ.]/;=�a��ݫ�H�s�z��:5���@��wZA��s��	:p�3\��أ��-�k���2=������i美��j�%���o0����0[\��c�r�x�ݑ��ڜ��/tPE6\�����5�}���Y!�Z��/��(��
D�Rn7���ozi�`�ޢzU�'?�9�L��]Lt��%L$Nw�~�������1���7�:�[����nT%X��0�)�7�>�ݳ #��.�GI7ʎ;�@�{������ݚX�f���g#j���h�q�tg\:+�<�K����{/���K�m{1�k���&H�%TR.��~����4ޠ��h�c�V[�e*q�
Tm%��s\�u�:A���$�'j� � T+���l����Y'w��f�Ur�����iD�:����,��~0�)¦}��@n�����p]�MJaRvu�ﶳ{:�u��\�,�ץ����(����R�7� ��o�ä� ����(�S�������yw[���(��5�ݫ�J�$�5-�i�s�.�]��V�֕��\�*F������N����l�5V����;%��߻�
�ڀ�bmʂ �V�;f}��s�ș�� �����)��ϹȤ��������J9RGp�������9�w����#	�F�`@��B��� I���+@Qb�p<����w�-/�l���u�P�FSJNA8�{�}�	�s�{�ـj�S�?l�(�JU*&����5X}�Eh=�تΤ������6:�9)9@�Yn�fJ��m�zP˹�-�����[���7��
訉�4�)M	8��٥���������@�{���K5��JI�L*�t���fOSO��np��0{ZM�6���E`}����n��Vw�X�ج��ٴ�n�*Q�ޚ�W�7�>����3�Y�\��$=D6�w����wTy���kZ֜��Aȭ$w�X�ج����ך��;���PJ"�&��D�%Hǵ��w%n�G]m]I̕��N�9���y���o�mv�ܖE��Y�Γ��i��7I�߶i`{�Y�J8�4����`}�������s�'�S�po��%Z� ��-��*�Q�9;�7^j�;��,�UU�X�<�`{߷�zz�h);���%6WX=��`U�py�ހ�X�r�kq�&�:	>�@�����4����  ������Gч"$��}�깒�+v����}|���j$����r��pf:����]�{O���S����g8;;�����KYo3��F�+�^�����n;WM=� �6�t��X���&��:h�.�[rJ���2ہ�]��u��7��}s	�=4Zvy�mӤ:x�x܁⼼���������ʻ(:b���ؽ�ڇ�pm9�`�C^����f���٭l7�e]*��z�2=k����:��r��mB�e�3=��-�ܕ.��]����ᓦ/�J���{��z��`� �j�
�"�f҈�EDT	�t[�����s��Ϋ���Ө�=��~����r>��>�66�6��`}���`b��v�~��@�٥�w�k�$�$�D*8� i��=�z-<f����~όq��u4F� SJG`}����@�٥�߶i�A�w]��e%�NJ�	���6����=)ۛ���=8�&�g�t��]�q��"�QM8��lq�ޤ�ݚX�`)*�=�z��j`��j�,@�M�d�ߧ���� *�P����6I`wn��}�4�ݥ��#Hn1�]�5�s�7S}����&_��y~�����E��I��S��V�{���$�Hw]� � Zjsst_*H�������0��y}�]6�������fޅ'|���d�D��{���f�Sb�a��l��6��p{W<HSc�6ʂp�;��,��b�>�s{�������
����ԔhND�Q�vt#']�8�o�'l�;�l�7]fGD��4ʒ��;�7�w6����#L���b�A�L26@@YM��RS�P dG9�5__���N ��݅V�eJlrIށ��J�;��,��Vܥ�W���@�߿R)�N����M�8^L��`U�py�Ӳ�f����}��F��ْ�pP���|-*�l9Ӷڧ�� ���7B�l[�%V؛��_���� ��}��g�쇷��� �[�#b���Ҧ�#V�~��$~�������0JҞ�o�5}77$�.���������G��T���o� ��ҭ�6E$���9V��\����]Uϵ�3����9�u��@��J���A"3-
�;P�����g�R��5"l*+�@�y��Q�&��=��`�l�?s���
\T�8T�==s���^3h�72m�]�mGㇷ����U�;��FГ��:#J�i�UD�����ހ�y�^3�)Z���e�*d�R��lq��@�n�X��,^�v�{w����s͛�~�S�D�Q�$p�<���2eN�2gu|��#�[0�-�I"H��$�:	k��`}��{�V�����>0P�T�TUIE�L�U]]`zOoϽ�l�;�ـ)Z��]�� 𖘊
!H�����}�c���=�m*[�e��$���s��/U��.���A�e|���皹����J�9���8�Ӟ�%�մ�tu�I���v��j�Վ�*N�U*��z��]:�ta1�j�2Nv��s�u�J:z�7*���G~��'ʞ�nP�$�75������0n�n��Z�.M�A��kz��;$:�v-[W����'c���c4i��[OH	�X����{ߧ{�ߏ����z%��c�|gv��uЦԕی-��n�&�(tb³�3j�$���]߾���v�J�X���� �ܥ[
n%#�����=��.$)Z� �M�:�l��]K���&��h���:��`�o�S�o-�����:̌H��6GTG��ٻހӶ`�l����)�D�r)RR�q�ށ��K�l�����`}�n�uײj��l���j �q���(t�\�MA��;B�L�ts'�&8l�\��!�J!�dR.����_{���.�Ͻ1�r�u�4$�t�Nás>�5�������W�Q�}���[ށ�K��7�ٟ�L���!�UUZTے9h=�����{����4�1{1�x��h��FS	���u��l��U�{��z��vE]�㉪�H����=�����zk�W��o��P��)0p�h�ۡ�&����6���Iv�:)����]ks������i�6�àb��`}����f�����Ki��	
S�4GTM�`A�4����py�0��eL��,��%)D��i�'zY�5X���v @ ِ�����p��� ��z�fM	k#��8P�ۀ�`4	�c
�dE�|��t��M�Sa�Y��'��;d���u��w���h�"�� �jֺf�$��P*j�a0���"�!F 	A# ;���݋c�"�ǒ�`�av.g'  ��B�0:
�憎��h����an�
:B�*�@� �3��S[w��c���d+S�����B��)Mæ�P�/P��:���Ή��ۣz�!CJD�H�U}�wa���}�.��z�R�Հ��c�!��c�]<0���7u��[�bP�R�fJ����e���H[�Ek5:#�5��*��Fe�T��eQ����G%(�#P���z��&-v����H-���kf�ua�Y�Z�M
E�Ic�>מ���酑UC^�яm[KC�� F�RH�`�����.�y���c��u3���Gv�ޑ��t��W#f�f/<�V�hZ��Q�6�ݖ8"�(��7�4��̹�����<�q����ǜ���Q��N��>�=ᇘն̽-zz`�F{&���;���\U���.���W��@�CJa��4b��T}C��!�����$��I)"b
=PaC�U�@�E__Dy�=�US��~�{���\�]U��}���ۛH�V�)"S��R+��oK���M������%�}8q��QwVL��RY}��)m��&���N�|�U���Xܥ$�'*$ۢ����x!6ݳБ=ga;&B��v�Ou��Ny	�Ӈ��T��cjG`}�n��j��`w�v?��r��W�]��(���Cm��J��@r���7�78�%X����fӭ�Ӎ��j�N;�{����U�{��zJـ��qS$�e�uyw=ɭ��4���V������1̳`�L�Ѭ�oRIH�N>�(b��Q����uW�����	@�%6�#�￳{�72i`w纬_f;�s��n���6� ���8��V�����ݭ%<Y�ܵ\�`wj���dl��5v�QJ��c�$����N�;f ��W���vCw��z��EQt�$Jt�ӊ���4��ʪ��^�v�����9��ۢ�$.ꦂ.�΀�[�*g�i��=�� ��0��1P['R�N;����@ݤ�  S�U�yjsE�UuS�����s��N�f �Z� �����U=�GĜ!�7�M�6o3e�#�	 ��f^1�V<�cp���(I����� �o>��^�<�k���t���]�8���Oi�S��N��<�ܓ<��"��[�B��]�O.��r?�7|;w��*m�>�Bpr�j�a��;Ƹ5q�v�pyh4\����v�u��1���5�uu�ݺ�2◩�1:]�#�}Xw�E�R]�4n8���m;�۪���̳�T�DQ:3O]f���{Q��7�u���J���:
���r�7X��ֺ��\��N�J�Ԩ�Q9#j��X��|`Ԕ�S>��ށ�+f��mӊ�H��*8��7�uX}�����zYA�l����$f�F���&꤫0ߟ���f�;fTȖ�0���Q�FJQ�䓽ԅ�4���m� ��р{�>�Ӊ"�ȫ�����&���v�n�0{[�E2��,���)��
)ASC�*�uۃ\�N�Ҳ[H<GV�[{n-q�|���ܟj�]T�E�]�@i[0��z�np��,�Y�-��I��7*����{ߧ�]�-$��XD���G#���9�*q�`�ٞ�%��}��T�i�T';�5n�;�X��V�{w� ��:6��nG$Q35u�Gu�0���=�o��n� ;���4*R�eF����4�����9m��i��s��D&(�ɐ�-���\S�O�h�b��s�W��	��z��rpP�AJ���TN/��������VV�3&7=�Z�Dӂ��c�N���-$unk�3�0�=����f� �t����վ�]U������0��LP��X�R�C�����*��D��G<�}���v�}8�2G7WEDF�
����V����׻J���k���1�7I�M4�Y�����9Ͼ������}X��`�~�n�]w)@�S��< 8z�D�#n6�L��l���w	pŕkc���e��Wސ�s�uֹ�����O� ��3QDm�#eF�,練,�v�ۯ�sf��{^�B�o���΀�7X��ޝ�j��۶��<#���P�v�noz��]Uߜ�.���T(~{��d�R���Z�$���X�
&����!���{���>�>��8ԒB69$�|����l���x���t�ȏ�����jf���3uq<L˹S��d{Vg���okq��I�jN� ��H�5 �h|M�t��~,jW�{�'߹�G�>_� �||}17|�*��$��OB�� ��}��fߞ�ܮU$}��J����*44�rod����6��|�s�	j�=�2�jbn6��GN}�k�V~١�Z�0���}�(|&.�n˩�&�p��0���i��9I��>13"�Br�C�Bqt�&�V�ˁG��䋚�<���+fb�v���5T�A�Ogqr��;<vg�A��n���;l=��K7lG�u�an����.��~���<��L�cҽ��'A`�d����R&SAIDc�1�8�g�|;O�Ҥ]�m۶���q��p��ꮉ��9#���,f`%�m�R��U竡Z�X�-l��̣#�8̑@L�����[B�]
���/���8�[<�]�}<�����m��(:���^G�sc�׾����/.��΀{ﾛ�=�z�n����|��jzp��"	��X����9M��;f -J��-�Qv\U��UE]���9M��;f -J�y���{wQL.�U(�47���j���|��@n��l70�.��qST_r�� �w�o�}��s�z_��f`�e�F���%:T��pXZFyL�η7]U	���j�ŸSOc1��)�4��X�w{�7^�>[�v,��`w�X�aI�ڠ��ށ��W]��p�h�����`�э�Z�h������b""��r#���3+ N�������x�$����>[��`����ۻށ�w]�}�kiECdeI��] m����1��Kn+蝯��h=�MuD�IM�#����{�5n�;�uX�1���M:M�46��ͭZ�x���WZ�g�N�Q�:^v֣)[L$ȣ������2Iށ�w]���� �%X�o�6��D�q)�Cq���V�1fc�3���@ջ�� �V�uTr�IM���@ջ��U_{�9���b�Jx���B'Ynj�HX�U��Vg����4ܒ���z@9m� �M�DJ��`���D�MF�rN�[���ݛ�)*�M��}�G��!�T�]�F*�܉39��n���ٻu�Ԝ��ω��[����N(!9Q��8�ߟ���Ē�}�}�[u���R�nB��fl�/2�9m� ���@r�w�&w���r��=�Mu@Jt�HM��`[�}����X��X��`N���SC�����R5n�:��v/g���z�LXbÄaeZ��W��a�5���Hj��"c�p�`9���4kU�1�J��mVPW]k���;��j��*"S���5{���<�`f�w�Vn�k��K�J�jB�D�:��u˹NC	s���vw�|�1��^�&�35����J�]����i�n?�չ�����z���\��?fl�>�nұ��%5Q�U]��[��{�r9ڣ��� >m^ �f;��W7�����nF�$nw�~_}�`�w�%BU�/6��j��"M9SM�a��T�<���ջ��Ͽn���݆۰�q�JR�N$�
��]�np�#��4/���>����^���̿��7�O�f�s�UQW�����PX��o]u�����Z�(�@�ihiThAh
��ThE�A�)T���F%Td%Q��)A(E� �@(H�iF�F�ZA�iF�PZAiQ��D�D�h ZQ�TbbPZ�T�)iQ)F�@�F��hD�)bD�U2JR�A��P���)Y�E�Z�TD�_��R��V�D��T�D&U(E
�P�(H�D��
hbQ$ZThU��A)h��BnB� Ui��PiiDHhU�B�Z�Qh@)�db)B�Q(H�V%��E
AR��H	�4
������J�%
%(��̨P@�"�G$ ��� �E 
@
B (��Z^�\�J(� �P�2�B��T��V��Iw�@H�H	�H"P�B�J�H)�*�-��1"�HR�J�%R+J% ���C@	B0�%(�ЈP�J�"+J4(УH��(�@��( �R���B� ���� �㮈7���"��J *��k���?���xP��_�J����2�� &	�'b!�t*��?���E4���(8�դ?���hP�Ѐ��(��U?�(?�����(��(�h�(�� ؀�����������_��*����O��?��Ȁ
*�������������� ���� U�������}�h�C����� �����?�����I$�J$G�?� ����L�����L��K�������������kApUPB`@	�ReD�DI�R"TI �Hd�$$�TI�VTI`��RTII!`�`�!D�$��%D�aD�$IBHTHBHP�R`�%IA%�RTHFTH@`�Q$VTI�RU�P	T�d%	RT��e!	Y	YD��d%RP$%VE%%RT $VBDI ��d$I	VBD%%BR@$!Pa ��Y $$@��X	A��HU��HU��BIBAII��BBd%RRD!%P$%@!$ I��Y!!@$%E��BPID H��I	VB %%BBU�!E!%B$$ ��HI ��``��@���!Ed!UHIT@��BU%%BDQ��D$	AYH	P	BXIDa!A�$! ��F �FRHE!	@`%D��P�XT�%BB%%�		� P!	@��I�!BB	Ea � ��D�!Ta 	PBF���V�FPHBd%P�IB��e��e	�%	A��e	�		T�$�		P�  �!VU��B�F IBe	D�!P!	� H	P�dH��$a!� `II�BXXBaB@�� ���'0a	e$H�!�$�&P�"@)AD?������W����r��+B7��O�y���ӣ�G������g� QW����_�ZO������S�� ���}O��`�����:��R�(��E_�ܟ�?��(���niU�#G�����[z���;�r��c5��u:�ݝa؀(����������?��A���l�����E_���E_�q��;6S���0Ο�\�5�xw�=ߺz?��{���?�:4�{������~�� ������ ��}����������?���(+$�k'+��`�T+0
 ?��d��1����EM[��@=��i�@h��[Kkblо�\w+U{�9��@�`۳�-��M�될)���f}>�� 
 4�P @�  �J��� �:4P��
�T @H /     ήg�u5��۠��(��J\�+�|6���w���wUyn-T����D�P�[�Z��c���mZ�p�^�>޷|�w@����  y���=�� ��u��>m�й�C���}��+����|`}�:�������_w8�>:�N�݊���)�<��l���@��z^c�@��p t��Q��p�v��� �� ����΀�����m�N�s� i��@  
{��s� t{Ƕe�m�Ҁ;��
S��� (0 �s��+ֹ ��6QN�w{�� <�@�{��  �B@�z�@�2�]䭛�w�����9�r707�`;�/����FN������z|����on�6�vy��h ���}��ǟ{���
]g��}��݀}��kp�}��G��[�p���о�dzi 4��()m�[��w�kڂ���	��|�u��{�����f�����6���5\۹��� �@��cC���W�u�����q���y�=�m���g�x�sL����.�m��wT�Ph�&�<@�����3��9�4y�	�շ ��ް�v۵��r���w�>�@�À�}���=��Я������s`������6�<��`��`      O��Fԥ* �Ob�J�ު   6JTRo)�� 5=��)�J�   =�4��S  ����$D 4x���w�����g��n�ԟ}�|?g���`W໿� @Ut ���� @U�U� 
� PES����{�nn��o{���A��3���n�l���x��p��ĩ���<���M������3<=���͇��+$,2g�:�6i�0�c���|�p�y>ǯ�7���_>?ӫ�E�y����+/�S�+yӷ�ʱ_D���t�w��ʵ�ߨ�n̬�F�=�D��2�M\Z�-�<H���u�f�B��Յ��v^�k�_E.a]��}���v�6��g�nr�9G6��{E.�b��WJ}ݮ�V�����TUߋ��f�c�aJS���4s�<��H+�N��OW+F[�ߋU�v�j���gF�.h&f�KLM��m6u�'3N�^g��X�X�g� �!.J�!������o�t,*��l�r�7	q![�9�6��ŞF�|�t.x��\���������.ƐW�Y�{�YUF.3s���U�v"7��$����.������7�J�����g��i� ���6au͓���92]����ٿ}�2jsYX��۫�~�`�b���Ɏ��3��3^��y�KJ�$c*����F�C��⨢��+y�7�����b��)�J@��S�he�2$�3�1�@���A�싶���^p����o8�3�Ĥ�9!�ϳ��}��K���6���y��=�y�|��R2����K�}�����06���yÛ)�!L����0����XV#��xh�9/�w'��I�K�3��Dm�=ys��f��\�\e��&�'�3_k﯇��|�0�����lJ�S(Æ���5�oH���i����Ϥ�����M,��H��v���m�Q�>�_K�yu����S�o����{�'��ef�fdM^r��_>w�a�����O>��|�n1:��̜��g&��k����~����V]�v�!H[��&���73�G9�0Ծ����L�)��aIj�dKo��7�B$�Ďh���A��8�p��\�|#7!ɗ�L,Z���$#�"1�D HJa���$p�.h�$���%��5����5�j��y,���B��sS3B�Ӭ��e���a�����	��|秐�ᴛa��Y�i�%�����|�s<FO �o!η���z��6$JL����M�a�{,�헜%޷+��R��yM��|���5^ B��!srW��Nkg[˪�QK�*�>�������]���9�W�5A[��֧N�;�k�����2�γ��r��|��e���v��k�|v�]��W@U+xr��O+��}�:\��;U�O9�Y�W�s�+k9{}�k��g¿�x��/�y_o����
��b�^�͌ިq#���ޛ���������.u�.�e��Z��Iދ���9v�3⯼\�����檾����||�(���9�W#g��y�}�V��xy�C� R�ѻ�g_����`}�_��&hy�i�Y=�93��u�k٣���{�釴�����a��0�4M���7��/�����_|aC	�e�yLx�y㭞�5�!0�xa2�߆�Չ|J�1)��/<�����'�j����������10(l<B%��ׁ37�&{
�ɪa.X�����$�9�x|)L>#�P1!HU�U�p��r\��M�9�kSsLh}w5��BT��6
�J�U��V�vC0�$�K)	
��H�(FE��7癩}Ӭ׎�I�2���$��B��nIu��$ nX�eK�e�Sݰ�B��!B4�� H�]��B��Iiw�8{@��f�R�08�H2�'��dJ�{�<!X^>���8�6�8���sG��zK��f\��껪�*�|���]����|�v�9�~q��i�an���]�+�O<��I�8R,�>�AO��=�>[x�[�*+��>�b8�(��\���\es� �l�(3K�Y�K{��v�7�>�����kg�v�6𭯇�u����T�:�f�D�_�ßg�f{�D5�%e��y>��!�9���׳��0�7�S5�S���B�X�f�#�7�! �%�t���>�'��+��V>�~�OvzO6B�B��<ݰdnBdg
�ˆ�4�
���
h���!�.�}w�9y�����3�!,=�>������C��ˇ�K��!�̜	rZ���r�,.$�� ���֡	Lc�#Z`˖q���˽��s�<����߲2��'�34��=6�>q6~��+��ڦ+[[ׅ�����W��q���Ivg�nRfk��Yt_)/ �r��y�[����PJ��\�S듅�x�	^eY��6w2����J�Z�<�w�4e�0����������q���-���>lϝS>�it��m/�]]���Q��km]�gi�f���g�u���K'����|�Z���3������rS>�\�T��o�M���]�.w�V��gx�¿����Źx����u+�y])6󚫼��W��
�;�ǻE+�����|}ABh�BWN_L�oZ�0����
��O6l�M��Lp!��2W!If��5�_�}g�^8�^	�L@�ǿ~7�ӗ��]�af|#y$�&��sj|'��}[�/�y�O2�@P��)|-�{��|8��m��>��Oe=�f3���s
Ue�/�F�
� �}+okJɽ�Sx�V:i�e�o3��
)Gis(���Wwʻ���r���WX��2��2����q��t;��|�k���w����=���l)Y��Eq� �	a����@�6i������/u������Ȓoa䑮�m��S<���Nϟ�BK��<����<=�2i/RKݣ�,��2P����y���5�5�*�����L���\���g{:�;��a���]�[\��b6�\���W��<�Si�L�����˼	��O$������x��t��>B�!%�yIe���Zx���;��|����]�!�z��f��C|K��E�dK����ɭݶz\ԣ
���_�S��_r�ǿ�GV�7
+��k��6����)L�º�T�5�Jq��L&o8a�[Þ���.�E�3��|�S�v�x;�s�fqG|�{��{�xm�y�;�l�g{~�z��L]��|�}ޔ.fStW-��2y<���	I���^6��wC�����}�u��������_7��]��Y�K����焗�����=��>$<�	�����<O���J���/A��6Ѭ�HO7�9�Z=OpX�����ܚ��+��8ZIq�l�7`	K�q�ݮ���__}��k~xxa�+�	���8_<9)���9�7��La.����r��8�'�c.k|����:	ym���������V;�13f�P�T+j����Q��s�O��7)��R�x:w�}��K���Fl�5qԒ"S���@����Z��K�&�tC1�$��IL	`@0�5���)��乗~��p�͞��1��!��P!8�(Ŀ��)�w��6��U�.N�/�������Iw��n-��;o;z�fUU���;�j��yܢ��ǩwC�⿻TUVes�YOM>��xR��C35���	���#��N��w�Jx�1��vp�Y��w����E
�;����\���]��tN�nf���'��o<٭d�/!��u�l�C����_a�&�K�����:��yI_n�x��dԌ���
bD�B
��"dH����S<ɠ����Q����3D�����\A���O�Un���:���f��xؓ�=`�<S�5#����B���������B�\aIaᒤ!(O/��'��2a��#0�.H �
�+�IK+��$�l-�HF�$bĩ�K$)
k~��ߌ�x_I !����It|������M�����Mǌ5�9u�f���
JQ�&�@�J���%wt9���|��R����ox���]3 ]�;j�ߩ=��^��'aH��n��H�*��6�߱ޯ�7�i*��*ۥo����m�uξ�Uڧ��gw{Օ�!=��hK�ݽ��]H]��_,��WC�E=��kWv�����}1#;\~B��#ާ�L7��w�����>�75���52��F{���\�vy�������	�M�<�o���g5��<���Ç���k�ߓ�5��ߔ۳~�sa|&fcsF��~��f�1��k�����,�����gْy���}���;��;��vή}E|*���>W}�u���:��Qe�:'4gJ-��I�6�O%�#4=�����#�}���g���;$ǋ]�`kcw�|����Bs9��6zd=ǝ��k��{����se:t+o�ԾB���3�)ͳ�kS+����=��/�Թs�]��a��!BQ�����9|#|�(���[���. ��\t�m�(̭�������~>�)ׁ{羱�	�Ͻ�Y��,Q�Ϟ�����y�v,#���l9pi�kG�=H�w�k���y�p�饅�j$���nH���˕�nMxx1�֟R��Y��/���q����ݬr�������TR����T[���;\U��s�W��Xf�<�W$=��	&�x|m)� _|7�$<�n4�Vf����Z;�se_���
���+t���ɅP�]����ڵ]��Qok������{�+go��r˱<�^��J��;�o��I�k��}�
a��<}8���S��ïrǆ����ʟmr��ߨ�y\���Q�'{�;.L�T��m+�� �BB$�$�_���}��6�j��>�s7o9�\�^�[��v\�һmr���S9�˺3:�;�a���w�]�|*��n���u�����]�W~��������������2f��'-�/�ߚ�=͡Ja�����{������L<�|�e�e�	)dK�Ja�EfX�P$��q�+��d�GI��o>��3|,�2��)�%�s�#��y��L��~֏���i��B��xxI:��H��R�lSҞ�]����)��J�~�bOp��I�����>:�RJ2�aFz���f�,M; #pf�Rs<�zy�S7xgRo����^��,�cۧ����Wk���n떠��������+�.�������G����he�<���|aLѳ�3[�0����s��m�Mg���j��a�a)���Yn��_K��F��Di�\�٬'=ޏ~�����������d�̹�WT;�_uk�.*ͪV�=�OBC�M��o���B�WN�x���6�c�^�5�i�
��JYJ�4���_8�oE�0�f�C�Os|!�n�N�<�I��t�ST��2P$����]mܘ���P�!L!V�m��ǆ��[�.���Ф$Ky��9[K5��Ro�0/*��b���r��,0'����u��w��%����%0tnk��6{,���y��B��G�%�iG��%e�:��z�Ja�IJ��\%�Og����=�+�/J�T��t���E���6��FO.ow6�Oww��5�d�ő�i�̌��X�٭�V]e Nx{��W8�p=Rka3D�*Ca��K����9�5a��0�3͞_7���q'��5���}������=��ω-ᴓf�<��Z�m޷r5��K�\2d3�2�	�Va3.�q�1�)�Ԍ9 Jj�F{�o�J�0��
�'�L��o)M�4g7���\$��q��H�Vk��+[T#���Eٜ߉5��r���ǁ$#IK3F��{< ��$�/��|����]������*��r���]s~*����|������?��)[�>��ˡZ�m�K�����%������l��xB�E�@�*21��2�G=�=�4���g��μq/Y!w3ϟ�y�Պ��������������UUUU@UUUUUUU*�����������*����������W�UUUUUUU��������UUUUUUUUUUU*�UUUUUUUUPUSU�F�+�ӻTF��UG+`z˛I�X=�[��W��P.�-ZzB�9tU�� u�A�v�/-�[x� �(1��s�v�M+R��'@mUp������U�0�����v�]Q�T�l͋��QG���:jU��i���yݚ�����"je�C��UU��Ux�q�]S���m��ǰ��g�l��c7Bñ��.�]� �bi�M6m��hҌ�ejz�ޡla3�n�J�ndx+��53T�s;�m�Ts����,	;u�NvCqҝL.|t��	۹x�>j�w��M��m�ea�Y�hF��i�et{�t�\��]umhB�;����ܯ��v` ��Ӱ�;�y�-�����V�^�Pv�4
�����8���0�NVAq%�ݷ����ZB�nv2И^q&�[-:x��N7���w��D��V��nV��ّ�囊g(�=�v�j��*��X��uܺV������Hk`㰼��<�:�B@ VЭ&�t�-sSQ���I���*��:2t�k"����<�ଡ�h[����]�SѨ�
n:��*T�
�d�mx8˵��#�x2�KǳJ�U�h^�̪��SV�M�<�P�s�Ւ��UN7`� {q1�Y�ւ��.1*�v6�u��\
\�x���Q:q��g`�*�t��@��Su>���J���ylJ�O>�1X���W�rt;Ay.]���ۀ2�[�j���v:@�eY|�+��s��4��sTlu=$���S��U��+�]�jj�ۥ[��g�5[w.[�ۦ�be@����EK �UU@�q#e�������>����<]4Rj��*���q��K\EK�Um����ô�*F�P��6��쭈�lC0.,Ԡ�4b��b�l��7�2 �v�6��ݙ�댆��Aݱ��=���&��5W�-`�:ݶ�j�����_:lk��MV�=�����c;Ի*�K2��'U][ 2�d&N�e�BQ����2��3�n��Cv+��ۍ�:��3"��'� �,Ѻ��ʩҬ��j�(�.
�wj[��PqR��8�&�n�0���ڳ�lUt�X:M��6��j����N�2r5�U��YV�œ�G\�lU�JQC�Ӳڽ�A´�xc��U�8�'gjv@��o1��x��qK�E��c�K��Q-:^�M]+J�Wmo\�ݧ��=reȼ����t%�����lG^��vAb����ƨr�UT��#�j�M��Wd�5Wl�p\�j^g+WR�=�sԇ*юTJ�ʪ���m��ݧEV��Um��jsN�����.����U�V�m�V5AU]U�U�R��W::���U/-UTUm�R�P���ZU����*����p�vk�l���w�M
�-�>�U��e�ک�ڗf�u�֪�}�R+�Rv�P��%��WH�U@t ]��,b�!m͵���RV�;V�\�Ѳ�6ˣ��#QX5�A*��s��Æ�b�*�Ub����K�PX2����͢X'�F��t��=���UF�gE��nں���Gc�j����6a�tj�U��b��K@��^ԅl@\6
s�����W���c�UV
B42��m�R�g������k X�X����f�J���V�j6�I�m�Wo������T<dx�j�e�_[����: z���q�*Wg��۶ݫf���ު��9qͮ��,P@�ͪ�O;l��+p瞵!UƦ��VǡAF����7X�du�j��7^N�7V��P����w��j����5O1�wp�*�uJ*0��p�R�UV��һ2��8��n��-�q۵�QZ&���$᩽g@������Y紤���p���κz�]d5[�Ks�Ocڛ�nݪꁶx��xj��aڬ�#l�#�V���$l;��ŷ����F�*�8�y��l��\�S��V��[]Qu'm��B��SqCO��Q����;���{v���	�͹��ʥ�֕������j5�W �]!�� T<�Q��v��&�[j(�۴=-F��/$*���l���^�4�P��aB�ֳ<6�ů�@u׮^�]mŵT�@[q�����V�] �#`�U½e�XK�n�z����g��8��J��i�U��ۋv�f�!`6bAu��-�P]�U#Nu�c`��y�#tV��U�U��mKE�� Wi�핍���t�
��yb�56�(�[;����UQ��Vxk�F��h�+4�����e�bbZ���*�{v	뚕gnM�Iy����9�C1�nAy,Q�fe\6���a$�ئ���������Y�[i�Y�	�Yu�B1C�O�sp@�!K�����J�cAĜs�M�L�킽�^���lA�:ܝ�y�1��w�S��,�W�p�W8ۉ-:wMS�ŭ\ô�ۈ���3�L�:��۶Z��69ڑr�Uxs{]�۷X���̫Y堶����8��Y��pq�SSg/Q4z��fm5�knt	�@/Z��5U<ڹ��N�4���WR�2�f3v\�,�V���>V9�(��Yu���$��Ի*p�F	�Z=�H涶�N�3�0�HfU��UQ�=��\OVQݕ�iZ�8*�s�q��MU\�[J�����1N� ���d�6��I`*1]=t�&�n�e�6��*�Wc�-j��UuR+wUR�&뭢���\��F�N@�Uy�^�����)j�8yw��v5UUP�UUUAL��I[3u&��0e��UR
��W*��U�q�jVr����S�/ �2�m�ʫ����/�<��*���cfUUPUUUi+ĠʨNW�M���S_K�MD9e��2�6_�eO��M�@5��̊K�a������j��5U��y�Jj�QVPU�6�i^��]��J]�9��-�����`ӹ���T��T�F���)UUUU�eU�ab�eAr�Up��S+A]pT�vM�mU�jCnk#�vk���Q�UUv1UR������F�:m�c�m*[V���[��AܕSj*���Wc"��*�R6��l��U����g��5UJ���V�je��F��U ��S��ۨ݁��;L�ۙq�R[���GZ*�L4�\�4tg��֪��0(m4UU�t�sWn�`<��2�]5�_��}mN1ʪ�V�R��^9��rY,���v��������b�f�d䰍���N�N�v�z�@Lы��Y٭������m�c�tS��ܴ S��+a�c
��Ws� �� I�5%��5a	�WR�pZC�BĖ�"�6�a�tr���3J	Fk�.���Ԩ���^�î6�����8e�EU�����h\R��w���]Ń0�б�Ƽ�5m@Wl6��e���]Uv+;m������������U���[:��V����̻����g��ХD�0kk�Dq�%��v�cN:�SH-�Ӟ}�kv�[�l��˜sAsWs.y��^7l��btT8��6В���떢�5�GM��铭�-��I�%X	KͰd��j�v�F�u�@4tpKQ%��a�S�$#PuUUu[/A���Wm\�����+��$:�\B%UuD�p����U�ju��/��U��V��`��KT�Mu!?]g�|��JG-�B�u��#�/-Sv^�r�#�`��C<#�WMT[��=�O(5UUUU&F७���[ ��:�V�lS��p9+��UVX�'\��PNƪ���
Z!#.@ �-YV *��-�j��y���ꪠ*� �ڡc�\�m�2L�j��H;�J�͌W�KV:�m^�*���;��v`���2UYqOc��᪪^Z��V��`�O*�d�mp5l���nxbeH�"�۪jڶ�����R���ubH*���*��|�[Y�3UT�Uҧʷ6��O�M��O,�mA���yUeN���m5�F�����R�Gh)j]�J��;/t3��j�Uc�WnV'��>'�����L�1�Sm�������5UUuURg1� :5 oeݝ��	��m)V��ni�h,�qYz���X��:�z�̶�h��n3�ꗰ-�&V�j�rT��Tq�dy[t:��aG�"�Gfw�N:b�gq���<��n�
V��',�USlz�}��O\f�m�a�J	��z̀kM֜�m��4�ۦ�jp<3��d&`
&��j��X�6�a�j�%q؞����s�v��e�cf�0VC�יt���m�)�lǲ�u��K<�m���]t>�Z-�c��I� 2�je@e�U1�!WV3f�TR�[mdR��ڬ��%�K��Qt��n�t.�;*qV(�n��M`������f�pm�tQ�.�����w:����5/e�9%��V^}���Ux
��qt�:3�������O]n�\jrE_�_����qV�*�����Z� ��p��s5 ��[�v{f�UX��UU&�Z��T-�/2dY]\v6ɱUUUK�=U����SR��;��yLU�k\AS�6�]\�E-�6}kj�2[9�m�i�����$A�"�����t�`!Um ��j���j�0TUTøUV458u�e{<�O5R�Ak:��5ːv��U�ɝ&�떀�0+�v�����!����ݤmlPl�[�V�U]��w�[c��,�=�U)u�����zS�������y(*��旞9��C��Uc����PY
^�Z�y�����,l�jk{�\n�፵�V�ӆil�=�c�(1W�n�wIӻ�b�� mP4�q ��_�'� ��"���"5E�)�('���(��/�P
�)T]�'C�@}*�@V��"��)�ؠl�H�Ut
�U�X��Gb
T1= Cf� ��@Ox���"� 6�/�;� �Q��� ��	�|`'�x�>��D�j}�S�E6���c���A~�/�(O_�4����C��EM�`PO=�<4 �ঔ�C�����@��1P_@���"Ԁ:pH�m��$Dt��5��.���Y�TA(�ǂ�+� ��]�*p =UW�A4*
s�$����ȄHĈ��)a ��IAc#H1��		$B)d`�d �� $T" � ����$ �*��E4(@}W�_AG<��F20�!�IB`H0d!	H���$��1��<J p`����1S�C�U_�<QP���)#a@�P��!-�Fʕ)%X���F1�B6�Z�j��I$kb�:6栋 b	��|����Є�Ŵ-�BA��%$�6�z�OLa`�@=���c�D��:���#�E�CJ��Pb~Q �S�����^�u�~*(LH�DB+X�LL#�Ts-�޵�kZֵ��ڪ�V���U�pʹ2u��S�v��ۄ#�]����뢔ԡJ�T�m����3�t;��-0�+XJ�Fݵ6JB�Z")ԁ21uSAl�וIsB�X�K��u�)j��i�`�싮tGh�s�b⬜�F�y�Y�ؔ;rg���ū�%)-����e�*!�b�m�F�)aY����s��n�̳��\-41��BF��bi�B`T��z��V�@�⤛:\:膔KMq"�M.�S#��fn�� Ɖ˦��	cX]	n�LX��u�B,�CB�]f,�r-e$�m5��P!v�H�� �F�F�f#��c�Cb�7gy���S;V!,��0��k��
q��&�* L��Ɲ�S�q�c,�H̴��E)B#s�Mt�D����t٫�!���3��1�Y�r�h�ζ9YG,���iZj&HD�e�<���vs���wf���]f�XP���6�@#6rݵˊ�͓=�Mm&-��ap9 3Yln��jg<v�x=�=���TI�H�m�c����9(�'.琰���Obۃ�P����"Yf�Vʁ��A	P���],nq����]��cvB�V���b�h�X��'fIi�QN��T^�c�-�ЈGY2.]���h��8tm�F�'-���������\l���N�*�5՗��q�\rF������8C9$.�<���;ry�O\�Vڒ��x��Ys���HE��,6b��؝��.�n��lc9���[vX��h�V뱄|���Oh�v�H��0\ Y�i.V㓜
-mvV��ZƖ��������̑��m՛�Wn:ĺ�q�\��ܤ�ʕV(F�D�ij��bVlUR�c�`E1de�`�FK!��9�Y(Vۥ-G������.;\n�x�nf_�����Nݗ�ŏ�&q�`���=R�ͳ���7�tf[�e	ͨ�7Y�d�]�Hc��g�C�ݛ��U췤�W�z����CX�[�]V�X�XL��MjkZPM	����� !��!�U�`'���
|��(x#U](�F�Rω3>�P��x�+�Ʀ�j���.aSXc�tg]rmV��KzQm�,P�`�έm�8Q���\n�d:�Ǝ`x��]�f�c`v��ŝ����*4��5�8�f��K��OR�`���u�0�$�nMu��<�n���7�4{^��`�#�		<<a1^X�m��B�nڅ�۬	��^.�Ra(Y�L�c2�M�F��;�����t�N�d}=U �Z1�'��$�D����ZJ�c�4�m�tض�M�V�������}�`f�u��UW�A�=��"��z��WhuWn��`[��KذmȰ�̬��J��lWhv��m�x%�X6�X�fVջ/ �+�k�U��)���w�x }��}���� =��O} �ݮ�4�Z�����bI-��W8�Z�b�I%��.q$�q� ��y�^m�f.K�+kn.ӹ�ݽ�:��7d��k÷d\�ishx�(V�c��p����޿t���Ē[ݜ�q$���C��Ŕ��W7m��k߯9�� ��$X��$%$jZ��B�pQH�I ��5�$R�+!,�_se,IV�Pv������fn�o�{�} ��t� �}�fy�]M\�)�$�n9kIovr�������+�W�$��=�{���MڷClɲ��{���$��دIr���K�r]�I/���wLٵֲl�����6_8�]��I%����K�}�Ul����a2e!3J�(kn�&�/B�,y�"jK	R;Y�M�ΐ��qۙ���s��WĒ]�{��$�n9kIn��s�%�}�x {����enX�������$���W8�Z�b�I%˒_9着��������kR�Qvq������[o�=�����E���wnK�K�r]�I-�N�m�B�;f{����� �w�����{���}�g��}�5i1�X-k�x\�%�%ێZĒ]��W8�Z�b�I?�{�2\��T���r�2��L͂L*%tM ��V�/[���;p\i��-�G��V�8�]��I%���s�%��+���ޞ����u�l-�l��I.�g+���UWv���x�K����$�n=ǀ�N�6��M������^$��\��^���o�ֱ$���+�I�,%����qf��� =�{��B�>־�v�|�߸s����@H1	�T҈xb�mS;��\ݶ�~՟��ی���c;�@?�� ���s�%��+Ē\��|�II
ʼ�m�J-b8����\�cW<r���#u��ݡ�Zۗ�����h�Q����W8�Z�b�I%��꯫�����%������f�K
l��@>7�7�$�}��Ē�n%�$���s�$�fX��ˬ�ɼ =�������Ē]��9Ē�{�I.l�Mڦ���`����~�NI�߼�w��w���@>7�7���������u�bg�N�/Iw���K�-�+�I.��_8��:�� $�'��}}ٰM�f�g4t���&�]Mù�nv�]���A�w���`�D֢��ܴ�&-�Z.L)p�l�')<Y����r�!4(͐�F��e̥��[�t��+�x��Ժ�=Bq�<���g@N��Aj���xnd�(3�K���)�0Vi�in\�B���l`�ն��HK��3m����
Jf��dR&؁4tI-��.�;/���wI����dc�����U[u�jMzPC���M�:.+�m�<��nM%��E�M�[��M��� �}ݜI.��w�$���s�%ݶ����j�Ś*�x {�����󓓜�m��� �vg�q$��e�$��Z�e�lH�m��8�]��^$��w!�$��دIs���K�(q0��`�mX�Ē\��9Ē�{�I.wr�Iu\�� >���tj���+|����K�܇8�]��I%��C�I/}��]k��Z{<�����0��aU6���G@���=�+t��B���S*Ӭ[uv�ⵝ��$�����$�c��$���{��������x u��9�.n�\�r�|�S_e�|�	��X���ISIH��J8$3R2M,�30$4�H,`BBB#.$ ���H0� F#J��XA�Y!&� hjTN ���S2ۭs|���~�fn��}�o��||���b���� �;�q$�k��I.u�\�IvX�x�i���E��`V���9'9�����!v�z�%�ڗx�K�܇8�]_6ۺg	��4\�� �}����ً�|I%ݙ�BZ���$�f����%�Ř^���цr�8E4Knl%�&MkA�۳ۘ�g�h�76h�S�Ē춢�I%��C�I-Z�x�K�ݗ�$�nP�:��am��&ŉ$���s�%�\/Ir���Ē�7Ē[ӷ΀�]^�o��||�� w��g9q@�	t��BM}˺�\��9Ēݙ�Bt­&�b�^$�����Jh�KIsvr�Ēծ���{<anh1�=��#ܱ$�7g+�I-Z�x�K��.q$��+6���WOd9�v{��,�j�� �I45�������7��[M й6[ˊa�$�7g+�I-Z�x�K��.q$��p� �>�^���Y63�@>>{w�����.ɞ9Ē�X�^$����s����Ak�M�e�]7m��$��<s�%6Ӆ�I.wg+�I-Z�x�K�h�-b�)�mp���vg�� ����=��}��零��B�U Aچ�	�99���:��۲���ֶ�H,X�K����K���R�x�$�]���?�>{|��zz͹se�W�,3'��uz��ޓ:��]�,K3�BZ�7Y�5h�`$��'n��p�wc�9*8`�̬{b�����ـݏ ��sve`��snJJ�ΐ[E�;o ��sve`��ݏ ��IF˲�Z��iSl�9�2��p�nǀrTp�:�v�W�ڡ�]��������J����r@@�U<)��>��3+5�W(NF�DN�'c=���3��jk.���ZщJ����8����(gh l��2[j6�i�at]�h��
˓F&��ұ
��,2��eT���Z�24�8dsF������x�T��hW���=$�eG��$��"������/�/��cD,�4a��tj�2:���m5���1JŖ�k��`�G<�Y���mQq�̸�j�Uؠb�ݸ]�5�Y.��P��̌�F�'��ɡ����i�|䧫0�1���Kq:5vv��r� >���|����ٕ�n��ڭPV���i�ݷ�rUȰn̬w\0���R��?������t�0n̬w\0����0�#-YwN��ݤ�������J�7fV��4�?���wc�+f sv<�)� ����;��n��Sn����4�ͷb��������a;FN{#1[�gas����5��a���߻�7fV���UW�W�@vO<di~�\k5Re�)�>���y�>q�C������P��8`�G�oe8`U�V���Y`��v� �� ��x�S��ٕ�qvZ�MZv��WM�f sv<{)� �ɕ�vk��ڭDV6�i�t��x�S�͓+ �� ��x�����T���!ի���Q��ՉiTi�JE���Nx�#EŶ��+h�!�E�ll���O�{�����;5� ;����w��Wv]ӡ+��I��;5�=�W�RA�y�}O�͓+=_}�����O�'un؛0d��7��0��\O��m�]�$�[�,3�9�7�<�!p0I벃�nki&`hN;)9�c	�2���-��ݙ��L3�&�����F��R�IYXa�f\����٘�`��.�%%�s�Yo$ϚO�K��=YL0h���ћ�h� H��&�8b�;[�\��|�L�9���٬��ktp��p�8�]yO\p/f�i�@�7I�(Irx^\���y�X�CS��#cd$ �R}����/9�B���|�8s��ێxkG��a�[�0y��{��B��ߺ3G9M(@�D ��\�$/1%.�2�f���)��Xx��B"$I\ǥ��Bs7��75�k�ʺ���ɬ<4�]y��8xa�l*@�Ji�,1 TH�c_��f��6��B�Z9�7T�%n��7�\���C�iԦ�Ȟl*b�sFe���eKuqn���.	w��ϸs\YIv��8�ф�K	/��JQ�F�BtF����))��W
�G�$��� &�M��P<U������B	$aG`�����H�� �j�D>E��7d��7�� �ܔ�:���+���7��0l�Xf�`{���<��ح��V[e6�Sf͓+ �� ��x�S�ڄC#��pM�g��%����Jtg(:�d�\� r�k=riňnw:m4�;��6�����ǀݏ ��p�}��A��e`[�׆�v�®��� ��x�S�͓+-�������9��}���j�Xac��}O�͓+ �� ��x���%].�mS�l�9�e`��I���ɇQ�ĀP�D�1.:!��U��j9`t�����<߰?;���0�m�V��p�9^��� ��~0�`i��>�����u㤺��K�eJ�R��-q�h8�WA���[mV.�`�:�O�l�5w���vL���,�J�1�.��]����7��0	�2��ذ�e�ݘ��N��[e6�Sf;&Vٮ[��� ���Ur�.�Uؕ� ��-�x�S�;0.R�c��
����-�x�o�<po���{�����a[B�"��f	� ��$�bQȩ��E��!��6�NNxk���h�wk{�^C90�3n1�䵮�m�ώ1��XP�'��/+��&͹9j�3����q�Mgi=W;��Aڎʎ�m%��a�k�r2�=ms��=ӭ��]�;k�̈́��u��C۟��.#�\�
����/���ҷhk����PL�@*0K8�����T�mf���m�SV��J������;3\��,&R�kGE���l��e��#J��p�A����jE��\(K*������ܵz�R��J�g��O�ͽ� ���v^�(�)`:���tـsob�;5� �ݗ�oe8`��)ݫ�t%wwe���p�8�e��N��,��$����ˤ�V��fV���oob�;5� 䒲�Ltˤ�Wm��`�N���k�\}��g��o��{S2�m˶��-66�l5`bd�**��,��h����%�IF��鱖Ҧ�{{ٮ&̯W�P,�{�]��C�ϊgq�at�.kWp;5�6W�Uu_}uU�Pne`�N[���~���o߬���\��r������v�,�\0��%���V��wv� ��p�7ob�;5� �+ �T���)��;��v�,�\0I2���S���Y��b�`�%���V.�Y7��]�{O�z���Dt�L�ꜗ]��J����k�o��rI��oe8`��`�V����2��� �ٕ�oe8`�ذ�p�9$��ch��:�e�X�S�������UR���(�$(��-I�0���J�������q��9�e`ݘ��4+�lv��� ��ŀvk�ɳ+ ��p�
�6�\������J�Xf�`�2��{{ﾯ���W���	��ˆQYfņf���lmbcn܁ٔT�:J�st`���n�JL�sӶ��Oe`�N��,�\0�(�����V���[�{)� ��� ��wfV�(�)tS��n�wM���Xf�`�2�����JN˺t+��Wm��\0	�lܓ�>5�ܞ�x ���|Ls� ݎQn�V��˧lV�wfV���N܋ ���_}�~Ve�+�Eњ�b��p��%`]l2[�mb-�;]�.|���tQ��v�p	��� ��ٮ�2�`�E�6]�)�`nE���"H�`��V�Q� +v��\��V'��Wm`��Mٕ�rTp�'nE��R�'Nӱ*�n�0	�e`�p�&܋�}Kd�}e�7a��	ݺ�9 �{���~��#�ܓ�~�f�}! "@�! 	���I�E ��@�$B0�	Ad�$!'���i��	"��e��s�-�W[d5�r�hAz;����n.ӱ�sx�� >l�M
p��ǭ�%e���U�g�e|�gB�����HɌ��ed��ljKf ���,u�+R���Q]�%�d�[�0�@uf�a5l��|v�P�Ep�����1U�2�l���f^>�����Xfɚ7#iT݃w2v�S5���u� �F�'9��䜛�l�[�&ɥ��z�c^[KW&m�����u͍	UJ\3���6��FWGJ��~��_ ��l�X$0��4Jv+�E��Uݵ�wu� ��+ 䃆;{���J��;b�`�2�H8`��`�p�9$��V�j�0V�;n�?U}�.��x�=��,��ݙXw\IӤ�.��P��v�Xw\0	�2�H8`���1��3cP��0戶]�M��1�,�mU�`W�&��ޞ�|��M�ˀl��7fV�q���O�����.S�?����y�@�9 @H�N��#F0M���b�!
cB�e$���@pȊ�"TP�g=��o�y`�p�}I�W�/!�6��m[���?%�X~���]����߲�(�%Җ��n��0=_R���6G� ���������� ��y���WN�+B��X�`����U��ݮ����r^ŀmv�#S�広g�ח1b�tOA�V�UMLDe�pR@Y�����o�#�������X�-��M���9 �r^�꯫�6G� ����ղ�][n�m����I��,d~0�̬��I#�N�&�]ӱZ������wu�_W�_A`��E�D�}���rO;��f䒷�
�_�+��f���[&x�&�e`�p���R�x���v'M;���v���ٕ�z����w���;��vA: ݪB���N��H�M�%Xv�D�D�����3�3׮H������w�ݯ��[H��N�j�p���rk��ٕ�� �=��uxIz�z�t;m�;Cfɮ朗6Oe`g��H8g��H������ZV�cl�6Oe`ݙX~�����W{������`�p*���)�Zbn�=UT��r����ܓ�{����d����4�� �@�Y�pܓ���]\��rf�[���9 �~���U}����@���{�+ ��V��ub�n�
�Dڶ@�m.Q�т�M�9_'�.�N�p^�)7���؝��U��IZ����G� ���ٕ��︃���`�B�~TR��6���諭��&�e`��� ���UURA��W��cN��]4�0	��X$0��}_%�\��6G� �=���f�u��&j���@? ����?��~XwfV��_}�_��v�_�_�~�m��hl�9/b�?}_W�������=?~��9 �W�u�������섄�F}�{���O|̥�L����2,B�.Ba! ��f0�!A�a@�4B�"J��S8s7��=��{&���\<i��e3ۋ��HT�L���n]]mĥ"B�/��c%�nXsFϾ=�|��}�{�̫1#��0��/}�ϝ_�XR?`@t�RQ+�`�R�a�O|�<=������:Ba�f�$�0-�����!I��\�!	 FF0�� Br��<2�!��!�0jy�g�h�6a��l�4�y��g�3*_9�����GL��JJ�y��aN�.�����m�h��\�))(J1̥�Eֹ-��R�IN�2��s'�z��e��I�����R?payM�c&uמ 	.[���;t6��Hq�����i�eK!e����R�����IraI�0�ZT�LB2�$�3&jSZ.K�OL���@���r�
�O߾�3x�ܲRM%<G'y��a�7	�q� ����P��6o{t�l[��H���ߴ�4P�l7��32K����d'"�f�^%0|>�o�=��ߜ�=��<�ߟUV*�USUUUUUT �P��+c$�g�ج�(n�1;���;T�J�v���\�nr[��fꚹ��bq�z{+If`c&��RX0�ZR�Y�f��[���5��d�.7@1�Ӈrc6���K��rAt����؄9��M1��8��J�7����V�l!��B8�}g��1�/A�O[	��:Z(E�5���s��qS2�Q�KYQ�Q�Ĵ�&f!+�`�`�5G�.yk�s۝ Һ"!+��6;Km�tL��4a�\��NB�2}�`x�ճY�5,����rl����j��WH�84�8��t�u[.Alԁ��uhB69Ef��S$1�Im�T������t�e��vw�e0�mI��ð��Nm�mn�V�����u����m�[sS���K�F �ܙ�WK�c)u8e��
��j@�f0�t�q<�]���rta8&ca㰁��U�ñ������l��n��<�RX3AN�KeCj�0���ףq�/�.�i�v�+���34�"���2��V3J�B�Ճ�Z\�Zh���;�Z'��ݼj`U�9u1H��`�eaIcuf�盶��̜`{Z��]��ۗj��6U,c������}&�u�umŌS+���M���YCR:Q)n�2�+��UG
˹���uZ�NU�A�KHn��l�@ҩf�ˁ�-Ua::�E+��4/1��mm�h��>��u������l�v4�v��mp���e��Xh*�d�}��2�]�Z�m/�Q6�W=���-v�3�z��"q�����4s�l���m�nRF*�MtJʺ0 ��Ӎ�ƞ�!��M� ��J�l�u=\,l�n�=;��V���9�[@�s3�m� :=��
]��͂½�u��B(����x.F�d.����~��s��l����\q�q�U���y"�j�Gn���"�vN�>�m�,n�,���hNx�i�<�������q1�VݍO[�X۵;����])��7a��d��
�pYm0���M�(]�33�wI����W�0Q�<H��O���
�����T�>g�&4��j��f;R-�Zh��	�2SX$����1du��麏lܶzcv�0�5��#��G�I���=}毌����%�2��-FX`k�+�^��ƑݷV�Tq�v�����D��"@�s�wc:W
�*�.�MR]�I���@^|�f�v�]�p��6����-��<v�	��KfYmЁ���5&ʀ�#��@�I�D Unqa��m���\�$�{$�y�I�o? �?=�ە���עy1�p��vy�qV�{�;�ck`k������Ɨǯ�#Irf�y$��߶nt�,O��xm9ı,O;پ͊�%�bX��_v�9ı,O;��˩%�FCXLպѴ�Kı>���� �,K��o�iȖ%�b{�}۴�Kı=����r��������j&n��m�*�9=�bX�'���fӑ,K�����iȖ?�T�"}����Kı;�p�r%�bX��������5�4e�]Mjm9ı����iȖ%�b{����Kı>����r%�`��{7ٴ�Kı/��-��!r]]SZ�Z��r%�bX���xm9ı,>����r%�bX�t��6��bX�'��ݻND�,K�������b�%�u]�N�W"�.8m$��4�ci\Y�1�;H��wJ�]<�Fmy���,K��߻�iȖ%�by���m9ı,O;��v��DȖ%��{��ӑ,K�������dզ�jh���ND�,K��o�i�\R� �@����EF�T�ES�$EҤ���'��}�ND�,K�~�fӑ,K��߻�i�����Lt�Jt���/��S`f�;E.�6��bX�'����iȖ%�b}����r%�6%���w�ӑ,K��wٴ�Kı<����ܗ3&��$�3Z�ND�,@,O��}�ND�,K���"X�%��{7ٴ�K����"{��]�"X�%�����)L�%�f����/!y�߻��iȖ%�`����fӑ,K����iȖ%�b{����r%�bX���g���B<�rR��o)E���[��rB{v̸�dLQZ�s<�{��ﯴCgBf���h�r%�bX�w�}�ND�,K���ݧ"X�%���o�a��DȖ%�߻��ӑ,K������LTcu��å:S�:{���v��bX�'�}�ͧ"X�%���w�ӑ,K����lK�C�v�ߴ)U<������O~�}�ND�,K�~��"X�=0U�
$�b{��p�r%�bX�w_v�9ı,Os�O��Mf�.��m9ĳ��@2'~���"X�%������"X�%��u�nӑ,K!߾�q	��K?��U3<���Ky=�o^O,�@����iؖ%�b{���ӑ,K����iȖ%�b}�im�ᬷ.c�f`f)�¶��c7j�q�6�1�EH��lu䠺�ӺCz�{ًn��f�t�O��%�by��siȖ%�b{���ӑ,K����b�"X�%��N��ӑ,K���v�/L�Lђ�.eֳiȖ%�b}���ӑ�,K���"X�%��N��ӑ,K��;��ӐD�,K��}���nhդњ�Z�r%�bX�{���r%�bX�t�xm9�Fı=����r%�bX�}�y��Kı>������L��je�k5�Ѵ�K��1DȞ�?~��r%�bX����ͧ"X�%���w�ND�,ʫ�6ьP��������;��ӑ,K���sS:�T�K�:|:S�:S������9ı,?!;����yı,N���6��bX�'�;�ND�,K�~?S��[ڥMr�%�´ƌC$�����"��&��������GmE<J̦�Tֵ֬v��bX�'�}�ͧ"X�%���w�ӑ,K��{�`"X�%��u�nӑ,Kľ�ώ�Mf�3&�����Kı>����? �@2&D�=�~��iȖ%�b}�_�]�"X�%���o�iȈX�%���K��qPl�eh��Oo!y�byӽ��Kı=�۴�KlK��fӑ,K�����ӑ,K��e�u��4e���Z.h�r%�b�b{��siȖ%�b}����r%�bX�}���r%�`)byӽ���/!y��e�y���354���99ı,O��}�ND�,K�EG�����,K������"X�%��w�ͧ"X�%��ƞ�{�Mv���%r�ۚ�# ��,��\� �b���2��ԢR�����@Ȏ�jQ!���cu۫��{��ͨpX]�m�[�ٴ۲rchWn��]����!���7��ٺMi��k���B��N�Mr<�ٓ�vc��:4M�� `����A͙�q�vڠ|���>.���� ^e{q�.�k��F{H�Ƅy�pi�Ůc�'t�gI#[��V9��	V�c��P�7 �T�jb�������u��=�R]}Uw��t�Y-�4B3V�ӑ,K�����iȖ%�byӽ��Kı<���؀r%�bX���/!y�߿~�չ�����<����bX�t�xm9���,Os��ٴ�Kı/{���r%�bX�}�xm9 ı,OO��Lѫl���SY�iȖ%�by��siȖ%�b_����r%��b}����Kı<����r%�bX�g�d���p�k5Mj�f�ӑ,K����ӑ,K��߻�iȖ%�byӽ��K�����iȖ%�b_~g�˗F��fd��k[ND�,K�~��"X�%��V(�?~��yı,Ow�ӑ,KĿ}�u��Kı>>>�~콆^�W99#݌����(%�
�U��E�	����2i�a�o1���#��'�n5��]Mf���,K������"X�%��~�fӑ,KĿ}�u�D�,K�{�ND�,K������4e̚�Z.jm9ı,O{��6���@�i�&�X�'���6��bX�'~�xm9ı,O:w}�ND�E��,N�~��[�)�3W5e�\��r%�bX��w�m9ı,O����r%��%��N�iȖ%�b}��iȖ%�by�ﴷY-�4HMdԺ��r%�`������"X�%��N�iȖ%�b{��iȖ%�����o�iȖ%�b}�{�5���)sD��kZ֍�"X�%��{7ٴ�Kı=�wٴ�Kı=���m9ı,O��xm9ı,O�����L��i�l�z�;��к�fz�J"J��#��p�!��$�Ͻ5v�K���]�"X�%��{�ͧ"X�%���o�iȖ%�b}�{�j�"X�%��{7ٴ�Kı<Ͼə٢��j�՗Z�ND�,K߾�fӑ ,K�����ӑ,K����Kı=�wٴ�lKĿ|ϻ�5�Fiə5sZ�ND�,K��ND�,K��o�iȖ8�FIF��(<L��=�wٴ�Kı;�wٴ�Kı>3�~��I5sW&��˚6��bX�'���fӑ,K���fӑ,K���ٴ�K�������ӑ,K����/�م0�32kF�f�m9ı,O;��m9ı,Q=���m9ı,O���6��bX�'����"X�%��ݳ��<��mc���sfv����9�n]i7#�d\��GhJ���]dl��:�5���ND�,K߾�fӑ,K��߻�iȖ%�by���گ"X�%��~�fӑ,K��o��Ym�4Hj�Ժ��r%�bX�{�xm9lK����Kı<���r%�bX����6���&DȖ'{��&��5rR�sZ�ִm9ı,O~��m9ı,O;��v��`�b{����r%�bX�{�xm9ı,OO��"e-�s.�L�:|:S�;�����}۴�Kı=���m9ı,O��xm9İ1U�!��!�K��w�ӑ,K��>����.Mf��Y���r%�bX����6��bX�'�w�6��bX�'����"X�%��u�ݧ"X�%��@~!7��-͛��qN��tg�(tM��6��)a\G%�뉉�M����{���q]�[�k�7�ı;�߸m9ı,O;��ND�,K�뽻�Kı=���m>)ҝ)��o������qȖ%�by����rbX�'��{v��bX�'�}�ͧ"X�%���w�ӑ?
�"dK�ڒ����D�ɭ՚Ѵ�Kı=��߮ӑ,K���ٴ�KlK���"X�%��{;�iȖ%�by���:M5&MkYn��ӑ,K,O~�}�ND�,K���"X�%��{;�iȖ%�by�w�iȖ%�by�w�-��&��u.�6��bX�'���ND�,K|�gxm9ı,O;��v��bX�'�}�ͧ"X�%��v�y~����`7�c^l�:0T��Yڢ��k�6��N�н��h�
�L���Yx��Tl���V��6M�_���E���`�T%%����ˊ�T�a��	����#Z]!
�N|s��H�v��2��Pv:��\�6l`6�c��J����CT 	jܚ���O�����Z��a]���F�3�CD�uj�`�c����[�A51�k��bZa`��N��I����ړ:�(�����.�OL6�<Zd�u��)��i�Fn�п���<lԲ�K�֮��iȖ%�b~���ӑ,K����iȖ%�b{���گ"X�%���w�ӑ,K�����Zɢd��Y��֦ӑ,K���nӑ �,K߾�fӑ,K��߻�iȖ%�by���m9ı,O���0�5���f�WiȖ%�b{����r%�bX�}�xm9�ı<�f�6��bX�'��{v��bX�%��w�3Y��NK���ND�,TlO���6��bX�'{پͧ"X�%��u�ݧ"X��`��?w���"X��N���~��ڀ�ɨ�3Ο��bX��f�6��bX�"���ݻND�,K�w�6��bX�'���ND/!y�߿Y��ݢll�Qͭ�\�-Zf��q+��@10��Y�ikf��m=�M,���i�Ο��N�������9ı,N����r%�bX�{�xmD�,K�;�ͧ"X�%��o��Jͫ5W��r{y�^B�w���!�&$�р� �"�ICD���Sքtb�d�d2)����ȍ$�1`���	62h�H�	 B�1pG$$1P�*&�T<VD�,N���Kı<���6��bX�'��{v����%�by�wمԴ�Ԓj]e��ND�,K��ND�,K�;�ͧ"X�U
��L���~�v��bX�'�߿p�r%�bX�{��kY���K��殮kFӑ,K��N�iȖ%�b{�w�iȖ%�bw���"X�"(؟}���r%�bX����E�\�hEO:|:S�:S���{v��bX�"�w���"X�%�����"X�%�ޝ�fӑ,K����~�b-�e2f��	�j20����z����r�R,eF���G���$=��a�L��]j�Z��r%�bX��{�iȖ%�b}�{�iȖ%�bw�wٴAyı,O{���9ı,K���rf�W.��!��6��bX�'�w�6��bX�'{��ND�,K�뽻ND�,K�w�6��� �
df:S��~?n�c@b�[���O�JqbX��~��m9ı,O{���9�T��V���no,�7#;����F5�Č3�����	C@o,�H��Fdi�l��RB$2�p��s%$IB�	���.����5`Q�56K�d��M���H�$���H$"N��@��͌d��	�-x��5����<`@�Xy+5� S0�[�98��g9�/̰�ZI)+
]``�4���`�&r�&�foR�(�N'��{/)&4��.R�H��%eii
B�)&�&�`�Z<tf��F��̄�#A��*M��P��a����n�HNB�31-!��4kP��a$!e��S�.�$�	l�af�
D2�n�M�D0�!��Q�j4Č$����bBׄ)aI	.��Sc6�5+"<r���1	L��"�b�Q �W�P�	�=�:�����t���'M ��8��C�ٱG���N���bo���iȖ%�bw����>)ҝ)��俷��!�իGFӑ,K����nӑ,K�����"X�%��{�ND�,K����"X�%��ӷgl�3&��ֲ�e֮ӑ,K�����"X�%�	�{�ND�,K�;�ND�,K�뽻ND�,K��N�WY&un���r���E�ў�T�E�+��ݢ 5�#)���c����z��%��u�p���Kı>�{�iȖ%�bw����Kı>�۰� ��&D�,O����ӑ,K��߿rkW3Y�MkR\��f�m9ı,N��xm9ı,O����9ı,N����Kı>�{�i�"%�bx{���MdԚ�4k0��Fӑ,K����nӑ,K��{�ND�� $ ��;���ND�,K�����"X�!y>�vc�v ÑIU<����� X�����Kı>�{�iȖ%�bw����K��P� 0ȟw{��r%�bX�����S.��!��6��bX�'��xm9ı,E���6��bX�'��{v��bX�'~�xm9ı,O�����~��=F5�;sQ����I�7EvI[s8PM�؎Y�9�U~t��-��,�@f�幣i�Kı?~�?p�r%�bX�w]��r%�bX����P�Kı>����Kı;�K�;0��˙��֋�ND�,K�뽻ND�,K��xm9ı,O��xm9ı,N��xm9ı,O~��;f�̚2kZ�u�Z�ND�,K��xm9ı,O��xm9�D�,N��xm9ı,O{���9ı,O>��0���Z�CZ�5sFӑ,K?
12'{���ӑ,K������iȖ%�b{�w�iȖ%�bw���ӑ,K^N��������D�<�����bw����Kİ��@>��߮�Ȗ%�b}����r%�bX�}���r%�bX����fZg욳!�~��E�>11]�X8-l����v��j^^�����m����'�U�g�ݞ@yqT�7h�׫TVˊҽ`uU5Ű �s5�I��V\Y��H8FB˫��eP��%�xz�:�T�2p���E.T�S����;rs�B�5��5n!b�R�
���V'f��5
g5��5;Fp�`9����źy�^B�5ժP����1�h��U�b��syx榮�ѓ2kE/gp���*nGWM��z��61e����ή��Fy�j�m�v�fy�ӥ:S���;v��bX�'�}�ͧ"X�%���w�ӑ,K����K�B�wt�'� ]��%V����/!R���ٴ�Pı>����r%�bX�w��6��bX�'���6����/!y�����l�0��r{xX�%���w�ӑ,K����Kı<�wٴ�Kı=�_v�9ı,O��_�L�:-�s2fh�r%�bX�w��6��bX�'���6��bX�'�k�ݧ"X�"�����"X�%��um���Mi�33Y�Y�ND�,K��}�ND�,KC߾�fӑ,K����iȖ%�by����r%�bX���i�뫅�3:��5�=B��.4���c��CB�09U�U��k4٦ֹ��O�Jt�X����6��bX�'�}�ND�,KΝ��"X�%��u�ݧ"S�:S��߼�,а�.���å�bX�}�xm9
: (�$S���D��]N6%�b}����"X�%���~��r%�bX�}��6��bX�'�����,p9�WΟ��N��������r%�bX�w]��r%��bX�}��6��bX�'�w��r%�bX�������M�hG3Ο��BHI8,O{��7�O��]�A$O}��&�� byӽ��Kı>ϯ�7�6�T�)�'�����/'{�?_8r%�bX�}�y��Kı<����r%�bX�w]��r%�bX��l�m³Aȶ�u����t�Nj�]�öf��-�=n�`Oi+�u}���w<<�9 <���kSi�Kı;���ӑ,K��{�iȖ%�by�w�`	Ȗ%�b}����r%�bX�gԿv�rCE�.fL�m9ı,O:w�6��bX�'��{v��bX�'�}�ͧ"X�%���w�N@�,K����v�Mi��3Z֋�ND�,K�뽻ND�,K��fӑ,p
A ��$d $D`�A�$@b�$�B$a�dU�6�
��*H�'�w�6��bX�'�>��{y�^B�}���~n��uW�6��bX�'�}�ͧ"X�%���w�ӑ,K��{�iȖ%��X�w]��r%�bX�}��V�	�$�����jm9ı,O��xm9ı,��w�ӑ,K����nӑ,K���ٴ�Kı/�ߎ��Z����
6]t.�;1xG���<v��dt̫�Ol#I-6�3m<�a�ߛ�ou�by����r%�bX��]��r%�bX����6���L�bX��p�r%�bX�ww?a�Zӆhְ���iȖ%�by�w�i�bX�'�}�ͧ"X�%���w�ӑ,K����Kı>ϯ���L��]ְ˭fӑ,K���ٴ�Kı>����r%�(%��{;�iȖ%�by�w�iȖ%�b_�os��欺m�usZ�ND�,�>����r%�bX�w��6��bX�'��{v��bXC�#!"�!�c�A�@��j'�s}�ND�,K�����\!�ۗ32捧"X�%��{;�iȖ%�b����{v��bX�'�}�ͧ"X�%���w�ӑ,�/!y;������lKW]]n���!���l[F���[�.v���jrl%������{i��]�h�Ο��N�����nӑ,K���ٴ�Kı>������&D�,O~��m9ı,��o�y�T�����O9=���/!߾�fӐ�$D"dK��~��Kı=��~��Kı>�����O�$��,O~��ڷD�LԄ��f�kSiȖ%�bw���6��bX�'����"X�%��w�ͧ"X�%���o�iȖ%�b{�{ɖ�5re̚Ժ��kFӑ,K ����Kı=�����Kı=���m9İ?	 C"w��xm9ı,O��yu�W�]��å:S�:}��siȖ%�a�#�{��i�Kı;�߸m9ı,O;��ND�,K���HD�@IQR$� �"BO�����1���]�فp�ߖ[�jzMn�h�v�2[V�k��d|kQE�v�����j���ri�|\�q��u͸D���E�R���llSBf������.#v�1�O->�(Ma�N�D)c��YX��Wm��=K1��guq2�e=����K��#nu�Kĉ���X�^q�l�l��s�:5�$��R�عic��!F`4a�m�l��rs������9�~q��Na-(0V���0��#�D�fL�u�]�z�.�fЌ��=�������MkXe�fӑ,K������ND�,K���"X�%��{;�iȖ%�by��siȖ%�b_�o{�[sY.�,˫���r%�bX�}�xm9�\��,O~��m9ı,Os��ٴ�Kı=���m9ı,O��^��p��n\�˚6��bX�'����"X�%��w�ͧ"X�%���o�iȖ%�b}����Kı<����a2@���Y�O�Jt����y��siȖ%�b{����r%�bX�}�xm9İ? �DS"{����|:S�:S����|����+����r%�bX����6��bX�'~��6��bX�'����"X�%����ͧ"X�%��O~:f�f�L�j�0����xͼ��l=q���h��n3S�ۋ����q���w�y獬5��2�t�t�Jt�����r%�bX�w��6��bX�'s��6�"�"X�'���M�'Jt�Jt�~���n�qtR��t�ı,O;��NCB y�J!�Cl�bX��۴�Kı<���m9ı,O���6��-�bX���yu���q����>)ҝ)���ݻND�,K߾�fӑ,(C"dN���6��bX�'��M��ND�,B�wt�7�5�f�:ݓ�Oo!y"���o�iȖ%�bw��iȖ%�by���m9ı,N����9^B�����(�aKsr�9=�bX�'~�xm9ı,?���m<�bX�'�����Kı>���m9ı,N�o/d�-Ժ��V��x�s8q� �e�4]HlJ��K����}$�w�kꌳ@Ut�O�н�'�;�ͧ"X�%�ߵ�ݧ"X�%���o�iȖ%�bw���ӑ,B�������fo(��3|�����bw�w�iȨ%�b}����r%�bX�����Kı<��xm9$�$/!y������FCUp	�iȖ%�b}����r%�bX�����K{� �"�$dP�V1$C�P ��HH�H��� � "��0��!! u8�l�9��9�iȖ%�b~�_�]�"X�%����u5��L4�Mfjf�6��bX��'~�xm9ı,O:}�ND�,K�k��ND�,K�~�fӑ,K�����CW)��pɣ3WZ6��bX�'�>��"X�%�+�u�nӑ,K��߷ٴ�Kı;����Kı>��~�����i�a�ە�YN��hN�k�Z�;wG:���3,��t��z{M���Z�Z6��bX�'}�ݻND�,K�~�fӑ,K��w�ӑ,K�����Kı=Ͼə٫����3Y&kWiȖ%�b}����r�R*��2%�����iȖ%�b{���ND�,K�뽻ND�,K��/��e�+)C&SΟ��N�������r%�bX�t��6��c���Dȟ����iȖ%�bw����r%�bX�ϩ{;2�ܹ�34m9ı�����Kı;�۴�Kı>���m9İ(����iA=h#��ל6��^B����kg�f�*�3�Oo%�bX��]��r%�bX~QH*�߻��i�Kı?w��m9ı,O:}�ND�,K�}��9f�����'\��/G��٧g��#��x.ŁT�v�T��8��,.�֭�å:S�:}����Kı;����Kı<���ڈ"X�%��u�ݧ"X��������.�і�dٞr{y�bX�����r
#bX�'�;�ND�,K���ݧ"X�%���w�ӑ? �S"X����桫��̹2h��֍�"X�%�����ND�,K���ͧ"X(��b}����Kı;�{�iȖ%�bz{����5����h�r%�g�D����m9ı,N���m9ı,N����r%�`'�;�ND�,K�����\ԗ5�.��ND�,K���"X�%��{�ND�,KΝ��"X�%�����ӑ,K��n���VX����j�X��;��+Bڵ��7��	�,����R�aK
J'��l��*KR]a,��	XVV2P�am�ۛ��X����m*B3>}+=��� �.�N9f��Ya�8BA� �2 $ ���f��ZD=b\$��׼K��9hF�e%!BT��p)�
�Y���<���
B��80$�Zg��D$i��!��{�.��֋@ˁK×7aɄ9$M���6��,�Sa�!1��(<#	earY7ZoM4�y��:�>���U�]UU�T�UUUUT��P<�+!��GVܪ��c%<v䣃p���{7���MŮ���Y�����WS5��bc2ꁴ�;����v�'�f֌�ǎ��<L�"�Ύ�C�-���maMf!wl�x{k-��%�ɮuw;��l +Q��-t֖�F&J�Zf�;�R�	.h0��Ѳ偺�\�]�,��,����;q���R8��,���<���YN���룚�����9�8��/�vܐ�C��ېݰ ��^='�=��8n�Z�{*��� &�K ;Y�Uqr��:Q;I(.5e.�����&�4c��m:�hm�-5ue�wJ���^�U�F=v4�N�*rGL�v����s]� �2k��㘖��q�N^��=�*B`ki�3u���Q����[��8�kU�pM$F�Uu�;+e�Nw&:	����Yc1��fkA���T�i⭮���'���c�i�9����2���kX<��N�� ��V�1V�A#4Z�ۗ�+�vV}q��Б��t�f�� h]��Mf�nٝ˞���F�y�0��4<0H�;VB}\݂��e��-�������%�H3�D�Ge�ӄ43*�E���U['��Z��铍��I��m���Y/2]��[���w�ԫY�x��e['G�H鍠4�k��_k�W9����
��eVm (7sKl��#3�%�7Rfj-���bL��ˮ��Gfq�t���> ]�v���A�ep�,�cY&��u���{K�\�<v�Zb�5�ڡkcAc�*�nA�eX��m0M��s-�(Z<����q�3���ݤ%n��n����j7K�9c(�k��l����lk��2�-V{��Ѳ���9�z�J��:6h��9�����k��\:����Åll3�w�X�j��,[�<��M�ND���l���a��ձ4�"l��i�<a6����m�Kee�Q
rQ*�J�RPD�2e�V��k��ΰ�K��D�h�w��M��
 �Ex*��/�|��]�C��
>6@F Z 
� mOQ_��z�%CL�t5�T7.�p.6�����y�L�^5v4�ٰ� �@6�@����tڴ1H���[��u�s�S�q����S�x�Y�-ۇu��Hۢb��k���6̗s �^Δ�\���C�N/k
�В��p\h�[0�)X��JbP	��7�5��(��H�,�	V��	�˨�XT���z4�֬����ͻIfk	�%���SJ��B]n̷5�����b�r��:�R�!kklRZ�p٪	Fa�ͿwI;��W�2����d�r%�bX�����r%�bX�t�xm9ı,N��l? Gșı;����Kı?gi��.�u�5��3Fӑ,K��{�iȖ%�bw�w�iȖ%�b}����Kı;����O��A2&D�=�5�@�L7��+.g�>)ҝ)�����v��bX�'�}�ND�,K�}�ND�,KΝ��"X�%�������T�W[Z�Ο��I��X�}�xm9ı,N��xm9ı,O:w�6��bX �'}�{v��bS�:{������nn��å8�,N��xm9ı,O;��NF��y`'����T���e�v��ڀ��,�uv���Ћ$�	���m�V4ݙ����K��y0�b]�Fl+>����'�N܋ ����&ɕ�v����[��٫�53F�{�}w�m&����{���Ds�X��e`��X��]�.��V�[����ٕ�M�=_}_%�x�V�y`wJJ\�WNӳ�l�u�M��*e`�"��}��-�ܬ�*���WE:N�n�m�6T��=U�}�~��'��	��Mҝ��ҸU�1���b�#��lVa����vx����P��t� ��Q��;r,��+ �����W��v�}��e`����'n�����k �����U}�G�~0�W��	ۑgﾪ���� �t5m]��=#�seL�/�qbF"�|b-��B1 ��SH_��s7$�}�rN}�&��wh��v�}U�.�ܬ�~��;ݙX�p�6���#��U�M1��X�ȰUWջ=�����9�S+�>�����700ۜ��
��51�X1\�i�O] ���
q��RnV��
݅���fV7\0vS����m�� +aB^�;�X��[�n�	���ꯒ;��� �߼��fV~H򊗼���N���[f��?�Ȱ��W�%�=��zG� �-j��YC;v���W�/k���=��M�zy?}�� H[ń"�wq!�D�)�B��D� ����V[C�u�D�	�\E!BdN���V�b]�Ê/��i
7��o� ����X��J��hi��w�e`u� ��� ��^��#N��ӓ��xPٻi������vtH�m�� u���g�y9�ߧt�_<���i�Gg\πzG� ��� ��^�ɕ�r���cV�ݪuv;f٣�{����<�޼w���&�����G�_;4fd�{0����R^���7��V�pwl.ݖ��{0	��vV�`{꯾���z��(KާmՎ�E�m��p�;,�x]�f������U��!�C�όou`FkT��j�j����ݥCU��H��P��I��9�X��1��p��]��0��9n�:���`�����ű����-)UB�׋�l�����ha�A�ǎV���J;yuqZw�e�]&��J�E���H���sa�5��e%�uу��y����:�^�+ؔ���Y��fM�09�#�JͲjȉ̹fY�.fi8+�W{�䜚�3P�r�t�f�sGG`X��n�7���e�K�G�m�����h!]�� ��߷�Eݗ�oc������}�}U����J�g�]���i�m�� ��/ ��w\0�6^~�����UW�]�����m�e�m����0	�pß|�e� {��_ ���\Bi���~�N�wre�����`��r���`즭RI��V��͗�z�������	�~0	�p�wmJ�ݵi�j��.��W]�8D��l���읺����㐼 �s�����+T�Ŕ�ի�.�{0	�p�}U�o���T�j�7aWl��u�ܓ�>��b$"�-�y��f��"����}U���½���S�uc��m[f�y�0��/ ��/ �c��ۅ]��i��l��UW�|���[=x{0	�p�;R�UtK(`'m��l�"���=�}U����=���;4p�D�]O��VS�f�Ð�
u����%2�]PZF:��띂�0�İ˰Vl�X�������`�8z��� ����;�~.��R�ui�n��'u�?U}UI�{+ ����;ۑg��U_]�_�~���j�$�]�l�'���	�ذ���(+�>��	�E�� �J��!!Bc��HB!"��vUVϾ���I�����=�۬���YN�Ci��X���� ݿy`u��U}���{��E%ڿ�Yt�am����諾&x���e`��<���ڗ`W8YW6U�iC\�,8�Dո�m�bS�<a��<˥�Mخ�2�`�(��e"�m�$~0�T��8�������v��E/�+�j�j�we�`쩕�r\� �nE�n�{�#k�E`z�	�m�c���y`�Ȱ�p�;���2�D[M7NƓk�W˺��I�����>��dd�	�A< `��Fd�ŀn��C��ui�n��7u� �}U���?~;]_�� �nE���aBX��A#�Mev\6R�1�qh%�ф�$�B��K�������r�f��e`�"�9ۑz��	#�I���e;j�MX� ��܋ �������}�߫��޻�����]?�v[k ��,w\0�C+ � W4�)MZuc��m6��RL�n��V;r,�W�}K���yE?h�:��O ���������w~����/��M�j���}�W�I�I`����	A��M��x�w�����)�Nsu]`�iUI���=s'n���h4�'N��'mS�չ�B�����k�E���Ŝ���t�0gr��-�S���X[�cm	��h$�W��srs�S��,oM�r��:sO3���.�A]f��;�ip��K��4>�s�iq��{u��{\sN�s��]s�q�.3��vi뷏t�w mG\�!�i�f�5�ָ�=k��/#��jC�PaWG@�����ͷp�͝5a�U��c)tؠEM	���������,��7\?}�n��V�y4/�f��cCU�����|�wI���?�e`�"��I�~�I4Uպ���m�X�~0�C+ ��܋ �l���M���I���{!��r\� �nE�ﾥ$��;J�O�ʶҦ�V:�'nE�s�"�&���e`P���R�e7wlnһ+�@͸X'ckG��t�cy`�}��EQ������U�G��-��w���?��� �ز�	ۑ`sJ�+bN�vR/WZ�ܓ�}��"8�*
u�2g�+ �߼�v�Y����=-Ax�mҤ��-� ���+ ���K���zG� �KҮ�ڣ�J���v� ���0	�������U���������I/Ԛh�������0����zL��=�z�	ۑ`��l��U�+���oVol�ls	�l=�4�K�p��y9�ػX&Z���G�<�ҍ&��G�=����L�v�_���� �y��;^���t�4�'J�l�$�eg�m�� �y��&����R�򲭴��I7X�Ȱ�pÕU���UX)^�&��M�&�V���o'�"�ݸ1!ZF]��m�5q��5Z	�A�A�BB9��&�����uHڽg������N��Y,��D��xҒ��h1"B���-<F͛��f�u��`�k)��q�-ܺ1�r�4��"Mηy�(3F��)Ԕ���K%�Q��R�H�I���@ֈI%Ik$�	�XV�L%�2-Y+��m3h���	�	��1�����S0��G9��IsBL��4��g!���e�GR��S2����	i� �Zx��g�w�9�$0��,5���IrX� �	o	|��5����-#&���ֈF�HЉu%%��ˉ�覆ݺ{3`Fm��2$�dL�(h�2�5���3S7�o�#Siy��R[, ę�p��y�r]���O9�7E����|�a��\�MR�HC35����g!y!d�P�J� ]q�̈́�,M&� pG�S� ���E$cEXB2XD�!	��HDHBAHq1��L�'�������
| m��G5<�kٹ'<>�f��}˻#h�WO��]��?}_}����s�~��� �2�	ۑ`����h[�*�j�0	�p�=[���\�s� ݎ�=��?��]4F70`���P��Pl�X0؛mb����}��OG$1S�*����jۻV[g �W���N܋ ݎ����k�
�<ڣ�]�)�X��Y�����<�`��`�&V~���]#�t�ݻM�O?�`�&V;{ݎ��WV���ݶ`z��g�}^�V;{W(�ꪪ��A$A���ss�}������yttH����7 �I��N�ŀn�w\0�}]{��Xb�lq���{�mk@�KD(!F�6f-�-pҲ�5�7��=����X��Bn��~����N�4�+ ݽJ�6�WO�n��X�p�${c�z�V�{~�꤂iSº
i����� �?eI���K�~��$��M���&��v�V[f�꥾�{��{o�X�p���&x�7�mQHHV�U�X�Ȱ�rnI����'���rM���H��!��A
@�f0H�LH-��PM����r�Rmsu��6j���尤�t��mW\���:jܫ@U[,ҭ!��B�uaIyR��l��&#e��̕B��Yf�m]�r�uBrJ�hɰ��X7=<k�z�;�����8���x��ʽ��H�r�`Jf� ��9ڳW�qv�Y��^��%C9��i1X� Q%�Y�3���7�ke�SS=�TKt���rs��3f�-�GE����R�fKۨ"D���li�%pэc��FPѰ߸��k�E��pj�����ǀM���e~���=��,���7V�t�]Ӻ��n�`��+ ���ꤎ����Ʃ�t���l�7�=��r\�}�U%7��$~0}����%a6e���?�_?�_ ��� ����e`�Ԯ�n髱�m�m�{0�p�;+\0K�����!��P6G!�3"6ep�h1�S8��l��[rЙ��L��V�6rE.�b�-�l�7u� �p�9.E�꯾��&���$��ۢ�ݶ+/Z��y���F# � 2�i
�$d!IT�A`16}�V}U��8N߸���V��azR�6�� V�U�0K�`�2��%$~0�S�rA���WM�펝������[��+ �?{)��R�����wN�m���p�?}��}�����y`�Ȱ�ح31�pM��] �Y����4eV[�r�6q0�ԃ[6X�L3CYU4�H�\\90�S��r,��� �?�a~�e;
��6�����X{r,w\0�S�{䍗��n�t��j�֮����ܓ�}��p!�w��0�ذ�V�WC���[M���RL�n�����X����<`Z*/Zv�l�-� ��{꯾����7u� �ҝ�v*
+q���F�Ѻ*!��Jms�[�9J����5:SY\˟�)}�	}�, ���Y�;������`��0H����v�N���7u�=T�$~0���`�"��U_$w|��;*�컧tSm����9%8a��K��y`G� �l�uo�J�;�ـrJp�9.E�n�*�}�QW_3a�%�	ed ���E� �9���ܓ�;�;��)�SlT�j�0K�`��I�8���9%8`������{�͍[���1ͷ=H�O:�0j�,���#G��Ҵ���͜	Si[m�4��X�-��$����$��Ww��,TU+��v6"˦�0�p�9%8`�"�7u�9UI���tYwIc�S�ͽ�^�{0m��QTP�nƩ� ����`��0H�?�7C��6��p�7u� ��� ��}_}��k�դ��qc�]����fb2�k
�up�ێWr�e�������>�:�N6�a��B.#+���ģ��f���4�P�ts,�.�:���Q�p�)�Gu��n��N3�l)ۭƹ�����(%���sF�0&�1�i�O!G'<�&�z��<\��rɳU�1�I�D0k�l��ڒ��I�S�1l�s�b����9��ǈ��n�c�mIIVrH +��ƴ$C���׵���|�7�\h�::2��%ƕ�1̥XW;'e*NҺj��k�I0�0K�`�ȰVɁWc�Һ�X�f�%Ȱ��X�`�	�e���&0cf�r,����ek�ݽJ��`˧Lm���_}�U)��X���;+\0K�`�4�e� �e��m`��vV�`�"�7�"�$.�A�+�	I�mcE��;[�16ֱJ��%4�ۧn�t�k.X4�����T��x��� �����e�T��P�-&kYa�jnIϳ��P`�T~����D����p�&��r@`G@65lT�M�{r,w\0�}�|�����y`��|������@۶��p�&��r\� �܋ �l���ΕН��l�&�2�K�`ۑ`����)۲�%v�w^�p�0��M��'o�=��wa]=u���j��Vc<,n3�>o���}��`��M6e`�Ԯ�n�*�uch����^���fV�r,Q��]��;,�M�� ��{>�f�A���B���E�+�!7��n�^��ܓ�rϡH�*E4�.�l���}�/x��X}~��5I/ ��T[t�2��T6���X�%���l��_z�^�p\MVR�� �U�لb��8X7m�R���u��B�%��A`��bm`���n�����r,-������фp��o�|����A��� ��X�%窾��;S��V���'e���y��9.E�j�^���1��X�blv0�l�9.E�j�^�� ���>����$BBIE�������H�D�BJV�D�$c#� o�osrO}�m���Z��Lm��5l��n��Q�-��w�����;R�s��+54yۃ<J�<r�\Of�1�I�l=���y�Kh��8�5��lhe�i���$���Q� ��0�D)Tm)��v[f�Q� ��8`��j�mFS�J�ݢ�� ��0�p�;*8`�D�jة؛X��'��$~0ʎ%Ȱ�w>wj�ںhv���eG��X�ȰWUn�EQE��А�I,��~�y��ѩ���׋c1��~K�ba"2B!#%)IF������g�fs�� U �9��\�a7����a�ı��پX�H�2���.�q36J�8p��:3���7p5��͉vE�c�e26R�*McrR%��+Y�D���̇�J>����Ϲ�ǥ��R\�~]Ms	���59���|�T�����5ag����߾&�&p�2c�'�"h�4��HR�a d��-%��v|S$a3��4Ѿ2V9dJB0X��a۶f�i�7��,��_�_�2��|��k�΁�[�I��x$�2��{���c;T�p%��.Ͱ����aq!@�a̌�2�����a"Ҕ,n������G=�k{�.x�n\eŉ>��	�k�!H7L��zϝaפ[8���6�B롃ЁD\M�m�6���f"P��C�LNOe��͐�,��6O����=�k���.�A��%~/M��_Yz�=$�N#�t��|ߚg��m#P��c)�)y�k�M���?��qHb� '�yFE/��En���k5�2��	g�xp���$HA�e%%�����)i���m��%4�i�$�A�3������ebn$��`���6m����u�5Y�C>�s����|�UU�����l�UUUT��Pp<ˀ��S�����x�CHɁ{�)�j1�sZ���s�R�.�P����7�њ�`h�����I�@�vIn�WL�i�3\T)a4H饆�g��X�+֘[<����&�Z,u����jn1����l�s�/.&�t�1ԡ-*h�gF�����#8d��.lg;��fy�[�p�X���N�ah0��)�6�@wq��NW�n�qn�Gc"ۣ�� [t&Ʈ��W��V�A�k[oCF[�YP�Vb�)��i��
Y�.�E��bG]��lb})�œ�8e�M�M���(/C/�'��Qt�S�x�8��v��c�ծ�fF�qI�����G����rݕ�����!�y�u�qq�Wg�܊���l�XM����f�)-W���VR��8�Ԧ�u�7�)3'R��[є�0Hcmph+	h��Όط2���ŉ��<+�E���V�֟n|ݑ�Q�=�ғp����6�G��V�0Tv�p.�n�S�@��i\b�rN��48�J�rz�\�j،&6i�6pr��[Y�ךE�0&�����d��s���Nb�ڜ\i3h�
U��{�*���u4�^R�pBl�l�̮3�g�i��ܸy����v��]����e��`a9ԣ�u#���a}(ۑ<��GI������Y���2Q������X��&��ª��)�H�J�M+Y6�\�nٱ��t��m�������pWW��e
0����շ^Gj��zcX,�qaǖ�6�Wu�p�U]F�;��lJ��h5�l�j����	��;\�L�\nc�%B^���VYcp�4%pˡ����P!#K�X׀���p��e�"�CGqf,�X޲z�,��`�6�F��2���s>��׃t��:�=!9��r�˽��ۣZ#*Gm�� �X��v�UHU����#��0�%�A�m�4ڐ	��,-��P�Ź�9���n�é% �OT�h��/�? 'D�vb�D��*UJ��8m�S�f�$���䎝���M��]��[M�v:wF�<捹 �7i��.b�5�m�,�j�)e��:d%9����D2�+2����Cq���xl���:�D�C@�Bf�q`X���6���q��C�]���^��j.uZ�NAT�3��#�I5ְ�Qк.N�{R�F�y�i"��.�a�-�73ώ�tn�q�
B�G=N�5m�`R;��Da
�
.�Db+�:3��c��3ka��ljA���#)MetJ�\J�=��)y"��G�6��N�v6�l�'k\0K�`�"���}�G� ���պ��e����%Ȱ��n��Q� �ޥw�V���E����n��Q� ���J��	՗i�ـn��Q� ��0�DF�"��h�m�eG�Uw��\K����������ݕk#�.�:k:�,k�>���t��u�qZ�@ͭ�R<[u%��oߖ�r,w\=�o����xG���j�Ԧd��ܓ�s��@qW\�H�`�0K�`��)�`�ݫ���m`��vTp�9.E�n܋ �Ʌ���:I�M�l�&�� ��r,w\0	�1�n�:��c��+f�r,v�X�`_�������؆�э��WUev�M[���v!D�����n'��sw6�[�j�����X�Ȱ�p�;*L�}�q}~��"4��n�`[�.�-� ����e`�"�7�� ݴD���E7v�wm�el��9/b��C�|����DZ Ͼ�7!68`Qm҉;�𕻶�Vف��w�y`|�`�p��-�L�w��ut�lUv&���7\0���{�wj}m���m4�9���"a�t�:�t����1��F�2��.ӳ��-,Yu��m2�<�߯���O��sob�7�� ��Yv��M�m۶��ek�z���#��7����wf;V�Ӳ���)�`�ذ�p���]���7��m�J�nժn�6�m`��su� �rnLP��T9�{�ܓ�<��nj]d�Yv�m�7\0���{������7��Q�����bnV�կ'�x��Oq�A>W�j���b�0�mV��V�����v��=�X�{0n�`Qm҉;aV��Z�6�Ż/ ������,�_U|��߭���vҫ���o�����[/ �ݗ�scPj�]]6�n��ـsu� �ke�[��=�}��o����e��l��E��m[0	��^Ż/ ����օ��Uj���(�e��,6��׆��l�#�v�ܴ뀍���捽n�Z�l�\<l ,څf^9���U �z���2��T��ƺyϻAbxO�6�	�Ja���
�sg;Y��XD�5z�n�u�)=�T�K�CNRg�1�غŖ+c���$�6p����:μ�2V����=Wn{x�;j��
J�\�OmF�����I�	��^x���3i���re�Z�4��������⬐z۔�ؙ�)YV�Fk0+�f[0�;���'� �܋ ��6���&ޤ����tXڴ��ۑ`�p�&��x����z��Mo뻶�w�vG� �ke�[��]���DJ������vـM���-�x��x7\0���-�TZ�&����[��Se��p�6Y��}��}USЯ_e���v�����'n��%�q;����/h�ɦ84RU�=t��8���R��m�?w������Ike�[��lj��T��,U�������x�B��А0"� ��DqA�$�ﲹx�%����9�,�[eWE���$���)%����7ob�'d�wn��-:C��i��8���j�/ ݽ� ����;��W���uj�V��T�x��X�6^�?���}��}��9����f4�����Ema�.[���l2��w\R��Xzc��ݻv� ��e�/ �^�l�v�EJ6���E�l�6Y��K�`���7u� �ܵE�J�[V����"�5M��ү��܄ �F!�AI`JD��Qb�D����u����/ ��ui[v�)؛X����p�6Y��K�`��):�Cm�t�w�n���b�9.E�j�/ +���;�ue�����rrJ��9Ga�V�2�J�6;MV.�i��Z�v�B���[`�0�{�r,f�`��svawn�i��*�X%ȳ��������W���ЯKUwvݤ6���;#���e^ŀr\� ի@�N����ݷm�v�,��b�9.E��}�}[��w�b�7m@�n��m`�{�r,{r,v�,HS���!Dx�x��٢�H�E�0�����l��x�Aqq�6��l���I��K�`ۑ`��z����G� ��뻶�iS���{r,v�,�G�Ix;�,����un��m`��`�8`RK�;ۑ`�3�ut*�Iջm`�8`RK�;ۑ`��s�+.Ӧ��[C0)%��Ȱ�p�;4p����m��0�b�p8��Ú��\�U�r�[��
y�gv�k�E]��ұ��pۡ���c�x8��%�R�H[tKQ[,ҫe�Hv��B�u��f|�RŮ�1έ1+lЖU���nM�ʡq�cy͹;d���h*t�féh�7�	�u��3���F���ʚ�y��|v�;.k0��<��iQ5ʘ�U�MtsAXYK�����&���ճ[��m9���Ef�M���GCK�@�F.熌���d�F�E8��� ���G���qW���5E ^��o뻶[k ���G�Ix{r,v�A�ӷe�l�;4p�8�����o�X���:����튒Vݴ�0)%��Ȱ�p�;4p�9%P��;T�&� �nE�n�٣����ym����t�X�*;ZCG+9{lr�C��Mu��k�	�0��������@۶��p�;4p�9.E�w�"�9�g�mڡUէc�v��G�ة�T��}Ю �O>�}w$��`�ឯ���7g�wn�7J�������y`�Ȱ�p�;4p�;��+��-[mQn�����|�_��	#�vkQ`�"�:�h
˫I�]�k ���Z� ���zym��?~��?%j�.���E�d�f�ܜ��F:��
�@a�M/��K-LˡM;-[g �F��)%��Ȱ�p�:�����b���m2�k �^��w\0�j,�Pբ�'c�&� �c���*���B���Y"Hh��a!2o@M`������W	n��4U�L�qe0�&�!q��� f�6xyXM�Č`SF���C6�)	��'%+�,�"&�"�ܨd(�)20����Ñ�M:%%��C2�2a���%�a��	IILq�i�	Cbs��51���-�kA�A ��`��c��Ѱ�x@�0e|�X:i��K��N�P&�������	�rP�R$�<��
xs�x$)�d�L�׾�$���&Yܸ>�U؞���F���Ќ�I��N��$�@��H�)���Q= >J)���W�أ������)�� �P�@�޹�۹'�v^ޑ��WWt�n��6�0�p�&븰)%��p�9�g���%WV'C��0	��/ �^��w\0RHi�@��H*�>���۪u�⷇��^v������&�,�hjt����7Wn���{׀w�� ��}U��\A�jz�[D�:�[e:�cm`������$���jz�K�`�n�Aݢ�v�l�7u� �ke��"�7�� ݴ|H���7bVف꥾d����� ��ɵ>�R(RJbи��E�|hM�5�ou�ܓ��>-���m4�7x%ȰW��)���G� �K�D��Jc�E��LE��ÍA��z�1�9����3��Hrka���wi0���e'e��vG�n��r+��"�9�wr���4۫t	�o ����}I����_��v>~�I-=����M��b�`����y`�"��}��}�D���$�����v��bm�&�k � n���p�;.E�uv�ՠ��)ջk 7dx�`�"�9.E�%�F�R"R�"H�b�		 FHA �F�G㰽�	��`<�����X�4{Yx�8U&�'g���qw+��Y�0�u��N�#ԉ�v�X-I�Lx�5����׮2W�d�d{r� \-��]e�s�Q�d3���1�c�6͒��!g�۪�Z�z��뒻p��X��P�����D�ld�����5�P%�ɀ��w՞ǽfm�vV4��*�{��ُ��m�F6�;�N���ͽX�V��-5��ý�c�fe�6�Kd��I��t<�3f����w������i���*;P���5_@����<��X%ȰvG�n�>$BbCJ��+l�;.E�r\� 7dx�`Q(T��I]�I�v��r, ݑ���v^ŀrJڗE�'c);-���ﾪ����<H�`��`�"�7�j⻱S�l�@����p�;/b�9.E�6< �Vԥ��/`��A8�u6��V8w�7�vi�����-׳H(V�U��J�ְ`����`�"����� �?�����c���]r�[}��O=���|���u�v�V9� ����,��)n�����un��������`�"�"ݺe�i�+��o�}�W�R�g�z��$� ٱ�����;���7bVـl��Ix�c�7u� �� .��.�:I�uJ4lvڼqٵ���N���n�o::B�u.Bj�V�Xge�[};�� 6lx�{�'��wޡ2׬���2��M� l����U}��G� ����$��Wԑ4�U�b;wN����$���\0�h���(���(H� E����4	r�]̀OO< ��ա���wht;f���OL�u{޼ ٱ���ov`պuwJ�)&��0)%����7u� ٮ��W�Q���i����iۆnon�άf�Wo[3^(�m��<����+w6ڂ�\�r.����o-�}�ۀl��Ix�ۡ(��E���v� ����UI���;����l�~�N�qe��g@����o~�V�r,T���p�5D��n�.�t�ڷX�w��X^�� ��&䏣6Db@� ��b,�Qr(O!%@�CD@���#
$�4�H�"Z���d���&�Ng�}�[���q�r ĥv[k �$�w\0�e`�"����vW���c�!L�2��n�.4���� �D�������$�:5�z�@��X�`�e`�"�5I/ 9�5ht�Iݡ���2�K�`.E�n��كV���+l��bn�K�`.E�����䤏�=�e`]Ԕt�"���k �r,w\0�e`{���w��X[.��ME��ۻk ���}_}SӼ9$����=�=��IӢ"a1�D"$R1BD$<�~�7씳a0Pf�T��C�ʳ�4�7gtq���U`^�'�3���;cֻPy�l�<�-@*��R�`�*푱u]�[D���]4�`���0]�����y���
s�q�:�u��qn�eÊ�cv@���<�t�F_0/a��*8n�[CGR�+t;2�ɞ��H��α�щ�t�
�ey��"ڎ��۷�qod�rs�21�I�mc�w{ӧ�0��DɁ��8-1��b��d��6��L�9�Y�3�6oU�r�J;Aa��K[�~�~�e`�"�5M������	#�t��?Z�.�͜fym���<��p,���$~0͙X$�2�m$��+��X��X�`�2�K�`�5R���n�۠v�w\0͙X%Ȱ]���#V�7E&�'C�`�2�K�`ۑ`�����;Ӯv`��m��&B蝫)�����Z�e��CT��(�q)^Ujf3hf4�v;u�r\� ��/ ݽ� �ٕ�uwRQӤ��t�k ��/%z����5>���rO>�훒s��뾊�E%�뱢���I��$��vl��9.E�j�/ ݵF��r�At���r\� �܋�_U)��5y*��Wv�]�M�%Ȱ�Ȱ�ذ�p�=U��Wސ�U��/i�u�����;4���f5m�B�pt���Le����v�1���8����{ٮ� �D�ޑ����;wM��k ݽ޽0	.E�onE��d�)�n�v*t+k$�}�s����+��T�g�MI|��7��w�0j�-]餛��X%Ȱ�Ȱ�p��W��R�9�jؒ�HJ��v6�����3� �\��9/b�6�V�X*02ch��Z(Mj��b��.����&�9��*�j�M"i*{m�Iݕ�K ���r,��,v�X�6+n�b��j�0ˑ`��`�"�7�ឪ����^J�*�1Ѕmշm��w�<�ۑ`�p�;.E�rh&"Ym%m����X�Ȱ��}7$����: b��*��|�� ��U)?�v��C�m`�p�;.E�r^ŀj�/ +��&;3��n6���K�;��!��!vxd�:���5���
�`�`d]Ɩb��}m��"�8���5l�諭� ��v{���ӧbmm`Se����ou� �r,Wu)n�X�]?��i��5I/ ���8`Se���B�����Wm]��7��l��x�%��(ح�����l�6G�l�eȰ�`O�0��P��&� �0�!y
�b��(B�c#�D�I�V1R5ӱc�E
x������FH� �M8�m�f�P�`DD��� �*J�o21&�]f�o	�����RBP5���D"�@�+	$$H�<��r%�si�)a���ʄH1��#$"��H!��ҜB��o�~�p�o(X���l���d���""UeR�K�i�jdq~��x�J������[y��78g+���79�i O s�_4��"��Z��{i�E�����h��oD(p����<-���<"1�	��i�sFEXD�)�#CT֭vf�)o�V�B	�!	�#7� �vd�`F� �	 !$ E`�P��e$$!@�X�� ��)tC��!��Z�����������ڪ�����T�UU/S��"�3��@\G'd cz��S�/j��.�^b�(J���������;M��]���N3�Þ�v
�7g��'.�a<ex�Z[;��ca��A�5B�JDъcxn��+k�,֘ �F��`�F����/.أ���К��E.�ئ!Z���̓m�W
#X��
]6�6��Su�飩������,YS���_#� � �#Mk([b�[KԄ��Z���^ �i(&���Q�k&��)W�r�!Eu^�b6�Ĝd��gH��sn6aa��إ�|o{�Ѵ�.U�z��{�[Qd���teͲ��	}B����m�[�7]f��@�N�2��.��[��Xm�] &؍�3kfb.)[�а4N�����j�ĉ�e5��ۃ�U�9^==n�LZ{��p������0v��޺R2p5F��C����c`��F�{�H�북�n�:�M��2�TFko�+-�ᗶX+c���.ě��^ �Ú�`�L;q{v;ELms��U�_�g�w)���������+�k�v;q�ͩ���y���M�*:g��%&�����V2�{ 7��*��V�%=��yi�.�=]����X��e�tn!1S�t��n�ʪ��ő�;�g�=luvNC����@�h��7\s<	R�C�c��99�6]�K�X�[f(0�*��s��4sa ]����.��{X�u���8��4����SP�ke����������z��ƻ.��B��'�Dp�Ձ��&�5��TpVxt[Z�s���ܸz�c/)��q�K]Tr�z���|-���G+��gy���)Ӎ����4��ۚ�b^{X���n� sH���aƮ[Xlt�V�CP&:�f�D3l�I���2�#.�iD��	��]�j��uUc#�v�gf�S��8�2��])QC����m*_z�c]���D�]�Ŧ혆x��C���8c@#eØ6�Z�;9۵R�Y�Qˏ= �I�-˔6m�sY5�}S� �"C�W�
b�����P��_`�@��>T<��@�ǖ��y�[Z\�im��ZrL۸n�q�b[�]��9��@�Ŭ�,ή�<u��>�8U:�E��v�|�0c�сx��k\��^��u�<e��,�:ٗ�v�7K�Vi���)Q��4\������E�yQ��&2S��nI��	�Y�O��:�:ʺPA�q�5eC�����YqP�-.mMV��	��Q{���n͵=�B���<����6���7kpպ���M�nW�E�k��!ɞu��[p;��V����%v�&�������6\� ��ŀl�+ ��M*�[Wwm���7xˑ`�ذ�e`Se�꯾��5�TS�uv�M��^�L��l�T���-Q.��tSB�իw�lٕ�qI/ �6^�v^�ٍ+v]�ն�C�X����`�e�5� ի`Sam�wv���'��j�u:�LQ��;(a7 mr8V늉t\�&�.�ym���w�ߍ�xf�`RK�5wn��M�ݪ˙�sWrOo����`$c$�$ �ЊhF�x��ߵ�&�߽�7{r,��_$l����ҺJ��m�x�?���p�5n��:�_ER�`��t��ـqI/ ��V�}�Է�<`��4�]�.���]�n�]��[���p�8����ta�D����0&1+�1�ѫP�n���Zp�j�'<���ɨ�^�2�MN���e���qI/���\A6���,<��t�+Z�xf�g�����#����o�X��yꪤ���b����;t��f��z��Ȱ�}� Z4dX
RD����) ʁb�`�(�+Qd~S@����3rO{�7$���:t�Z�ݴ��ۑ`�e���qI/ �ݴ(�V�wj�]�[X��x��}3� ���x��X��ΰE�\�M[���F:���9���`����I����lИ��!+rl&���ٮeȰ�Ȱ[%�Q/��L�J�M�l�;.E�����,)�^ٮdҥ,e��+��X��X����p�;.E�}�z��m��q\-��ܒs�w~�����r,����}_|ꫵKvwdh�ʘ|�]:I��;5� ��������Hh����v�@�Ѹ����S���)�l�0���2\ni礳]����̳4T�������V�xf�`]ԕ��-X��ݍ��oc�z���䈧�x�?eȰ]�E(;�[�Uj�l�5l��vk�������_��	�~0�T�p�E]6��ٮeȰ�Ȱ[%�Q*��L`��t��ـv\� �܋ ղ^ٮ���$;w���5�2���ik6�j���%�d% � �Yvr�)���v�^#���z�_Z����nqۉ]�K�pk��jlR%�#�)@�sV�G�����ExMk�0���3P����k�aGTnS�J9"��UF�<t]��AR8W����b��C{S���m�vTg$B��Z��՘��kf����C=t�t��<[U�Jh���l(>��	�I�%�x)|i�����f��L�F�D�z���.w0lZ�6ͩ��1��P�J�7j픮�m`o�X����p�;�� ޑ��wt����v;v�ղ^~���H�G� ��� �܋=U���:A������:I��7���;�� �܋ ��/ �vc�]݉ۥcـwc���ݹ����徙� �ؒ���e����ـonE�ul��vk��0	"j����e����Wr󵞄�{,�:&�^��Y�����]�V�^3Cb����E��zw��巳\0��oc�ݲ���E����ݻ�;5�
�������`��j�/ �B�Je:J�6���;#���~�ꤢ�������DE7Wv�]�m�{0[%��e`�"�7H�ʻ�T�C���V�x�����+�o��X�p��߳�]�i�Va �b����:��c���<XtnʼZ�m	���u���^�p:J���e`�"�7c����� �{׀n�c�[wt�ӱ�n�ˑ`�� ղ^�&V��I\]��4U�k ݎ��xX���� HB,"B0�!�R����<R��P~Ϫ��9��l�� �[��Pj�۴��bl�5n��;$��9.E���(��iКTU�m��;$��9.E�n�V����\J��vっt�6�� v�ݗ���{p�u�d�ݪ"bc\c7iA�nT�� ���X�p�5n��;$��9 ;DSt�ۧv[k ݎ�H�O^����K�`�j�Z�R�V��;M���xd�X%Ȱ��w�2�&��M�D�n�����}�wٹ'���nI�k�>|�D@� ���������=����.S.�����8���n�V��8`P�o���K%��ո�]3ږ���Qlʌ\s]�$�X���Ĩ�S)q��p��jݗ�vG�Ix�ݴR��V��V�f�v^�&V�$�v8g��ꤍ�Q^�n��m**����{+ �^�0[�������N����.�`RK�7c��v^�����{��vz�t${��]�N��w�oc��v^ٳ+ ���rO�H���7��͙m3�+]Z30VZ�h�MpFjY��RZ�i�u����um����;p�`v#����sN+���%��z��l������3��
���hѱn-İ읞f�����Yw��jC������O+�[�A�ŊU��ŧչ)ލ�v7eL�\��7�e�k(��L� ,%m��ϴ�%�s{+�����hL���`��6$��S_�o{޼PG ��w�ֵ�Y5��F[4ʹ] G����4�ۍWW���	��BИe�%�[�Hfb�-������������8���onE�w�2��)
�t�w�vl��8���onE�jݗ�se8]�;v��v0v� �^���v^ٮWu%pwj�-�]���{r,V��\0)%���h�v�;J�&;k ջ/ ���Ix��X�6�{aV���E<`�l3�;ͽ�|c۝�3�Y;q����3�χ��HL����&��������wo �ތ��o �D��S��٣Yu�ܓ������*���������ۑ`��XT�x6P�t���M����{�6^�$�zF�;�J���'i۶��ذ���)%�ۑ`�̥���
B�	��uM��qI/ �܋ ݽ� �v��t���e��؇�^��'��CNM��S�M	K�N0l�ĵ� ��VЭݥt�-7x���Ȱ[�������J���Z�aWi�� �܋ ջ/ 콋 �^�����V��V&���jݗ�vk����3�2�)����ɶ�gǵY�LP�K`Pu����H0�&1)���oH�F���M�.K�s04&E�0A��#��m �i�q��-)bd�2�0�ݦ�.>��i����cHD�M��Jh&Ќ�%*R�y���y����ǜ��w��.���O�����L5��<d"�(D�"R�1ա/7ra���.�m���	~��y>���>���Y=}���"HI9�v���H�̙��X��x�$��,啒�^����8N9q��O�z�01� �}�1�{�p�I
`Ҷ,�n��r�|��<� ���	v(G�2�1���F#%��K��2@�	����A1�#x����|ޓDB	S�
�m��i���f̦<FDd���P��|Iy�{�<�y$]�&l���XB
R�40��-��a(`K��I�YH1H���[Js,(�tD8���W� ��@ >�m
��t �X�)�RH�!!$��Y	c�E$$!!HHFH���BDXDXD�H$ � I$��P�D1a�z�ڨ�ϻ��;�6�X;���[j鶕t�n�?-��}~��7�"��U}_)rz�^K�Q~�hV;�N�w�r\� �܋ ջ/ �/ ��J�Ƃ�iI�ِe�@��28y�8��`H�;\�]�[�'Gg���8���4揶7�"�5n��:���UW�q}~��&�k�;(�n�	�v�V��l���X��Y�Hݞ�LC��|'IЭ�W�� ����{��MZbV;�l����"�7���rO}�~��=>% %	@0m!����A��i2ĪS2�0�LIB d�!A�Q�/׾y��}~�۞ڢ��R�[f���{�{�0U}_J�r�VMպUi��E�d.��3�Eռ�<q��n���$��h�6����3�Z�0�Mu\��{��ǖ��b�9#�������݌���ںm�E];m��{{�������~��7ob�:�(�*����-��rG�r,v�,�{̀������m�6�X��Xv�,�8`�5(vQJ�]$�M�X��Xv�,�8`��UU}��v�>�1�ib,Қ����xN�u����e=�EjDIv���F*X��CW7f˱4���4��Ɩԙ��Wͅ�v���7m��Y97J;6xld�&�n7��e�W\��q:5	��1O]��t�Ppu�g6��y�g�� !	��9f�h�.#f��Q܆�!]��vǖù�	�b�p������%#�īP�Q��YJ'h�0{;8&%*B�j�;��N���'��򣡦RfXvWc;8Q[�K�uTX�(��ee�8�z�[e2�t��6�ƺ䭬e��0lp�7ob�;�0N�1]ӱ]&��X68`��un��;��gﾤ�[^tՊ�[
�V����ջ/ ��ŀsnE�j���Ҵ�Ue�6`[����X6�X�8`�en�6Ң��m��{͹��V�w����:^�ڣ���Є��,�[7����yݺy9�e�v׶)ݞ�������st���9�"�7�� �ݗ�v^ŀs`;�JR����ݵ�oc�w����pP�]ٗ>�nI�͹�#P�U۫��N�fջ/ �͹�0�̦_��aHT�Л���X�x�p�:�e����L��v+��]��ql��n��v^�r,�US�>��ҬDK����f��K����D��Z����\��6�r�\�uR�P���-��� ���ջ/ �Ų^���%Dv��iU��ـun��;.E�ql��n����#M�vҢ��m��r,�d�=T�������b0����%bF$�I�l(�"C��t�@G \�y��:�=xTJ%EϘ
�t�m`[%��� �ݗ�v\� ��LR�j�.vO-�}׷�o�s�O�����y`ۑ`bKc�|�����gt�c��@h��[��v�H87;sw����TjbY�4-���}�w����ŀsnE�n�wf1�?��$�ӡ7xeȰmȰ��un��9ݘ+V�wl���av�͹�0��xeȰ��t�S��"ڷm`�� �ݗ�v\��__P$$� !�Rh��GUȰUݱ*#��wj�M&��v^�r,�r,v8`���u����v�P��3,�FiR5m�9X��{VWuуn$̤al��:R���z`��Sn���Ų^������5I��5y/%E��E+MӦ[k ��/ ���v^�{z�������z�j��m���7��ջ/ 콋 ��/ ޑ�һ����&��ـun��:���8�K�7�� �ٍ�����M��6^Ų^����f�+�|0$d@���r��vw]]��,Sg�݀z�i�$��n�t���q�ysj���>����ր4��ێ�F��۩�p���m�5cc����!����y�,m�\c&c��l-\�r��q�/�i��>*㎚m<�u	��w9�;��XE.\un�L..�vS�зe���Ҙ듲�rfç�L��E����m���4�͕k��	tK���0�rL��*:U@��}���K4A�RŻM���T�������^�뗚��Y���kHdˤ������ۑ`[�������t�Run�m7n��Ȱ��xT�x�x�ݰTF�-'���m`[�����-���ȰwZ�.&����w�uM��qI/ �܋ ջ/ �D���ۧJ�w�qI/ �܋ ջ/ �업�ޅ/�a]L[fMM\�K	�����d�n����P� v�Y�id�h���M��܋ ջ/ �엀r\� �H;�]�V��	���X��x넌R�$��"��Ⓦ��$�6f)Ad"�rN�%�^ŀw�"�;�2�T?��Rt��]��K�`�Ȱ[���f��ۻH�[����r,���v^��/ ��\��V���X{r,V���^�r[{�J޶��0�"V�i�!$i��A'��[��v3�ۧ�$�z���@�Uۻl�I��8�%��"�;�p�9��Gm�v�t�n�.�x%Ȱ�\0[��(����0ۧJݻ�9#���_v�����着�W�}X����]�x6���U�!�n�v���V����0�e�:j��wm���x;r,�8`�`����R�WG4�+D��b�mB`.��=X���Wt�Mi���Jep�=�;l�+�ݿy`�� ���v^�م7j��v*�[�v��0�̬V��r,���pn�v�V�m�wfV�v^Ų^�0�ݰU���X�K�׀uOz�}�}w&�-٘3�L%[L����B��Fe
�
 �$��n� LSY�lܓ�}�!r�t���m��8�K�9.E�w�2�[������vQv�T���Qc� �0���eHFkH�9�bB͂°\ZV�أ��i:�Ct�[�x%Ȱ�fV�v_������O^�^vt��!�i�M�{�+=�W�$E'� �y`RK�7�MZ�Tة&���X��x%�X���̬��,O�Rlc�x��]�XT�� ����:�e���,vS�wi�t&�Ų^~�����v�'���}ՀWꪤW�`
��E��*�+�`W _� ����W�@
��� �
�R
�T��������`�E"�E`�@H*
���`�@
�D��b�E
�Q`�DF
�H*
�P �D*P��H*��*��*�� �D*�Q �AX* �� �AB
�T �@F
�Ub�DV�X*V
� �E* ��"�E*B
�P�� �D*@��D*�`�@V
�@`�@D��X*������ �A �E*V
�P��Eb�D`�D �D*
�@��@**���`*P��*�� R"� ��E�� �@UX
� Q�� E �ET� X
�R
�AX*`*D �EP��R�
�`�E� B
�EH� *@ �A��B� 
�@��`�D
�
� *"*��H
�T* �@V�*�Q
�PH*E **PH��A
�UV� �EAH
�P��Q��A �@A��E���X��`�DV�*��ER*�A`*��EV
�
�b*@ �E@��A��DE��P��@Q *A*�P"*P
�@F���E  *@b�EA��E��D��B �_� @U� ����W�
� @Ux  *��U�@
�� @U����_� ��� �����d�Md����f�A@��̟\�|A�ʥ��g.֨��� �$��@ t :�ʫ�Ͱe��vw)hA� (   @P $�       P� T     @   
       6�� �@($��(+�C;P���3��f�0 �����z��=�{r� K�  �C2{������nxx�9�v��WO=��uB����{Xܲ�s;���  nA@@P U b 6���6���#sk�W��yw����Vl壳�����R�R����]�� c�C�;R�h�WG�[�76��s`�F���8������9hv�ک\ 8 ��U   �jA�+�� � @ �!L �4�6R�)f 6R����� ͔R��   ik  ق�����	� � Q�  d@ƅ� � � 4�  �    �(
 (  ()�j�� iK0��7Ysz�t�E]�m��N�s+˝�KAkw��͇ vm��&D�et�Ɔm�Ş�oY��ޝ^�EE'hV�6]���t��ƞ�  w�P
 �$ 	 `r�mu��ny�-=g;�[\ ����\��\�Ӯl8�6�wuJp3��m:�  Ӽڧ�;)VAaFm�9���s���֗P��֢���3`��CN ��
m�JT�  ��R�Q��P�#�14�i���`"��E57�US@22 j���)=�J� �@�HSeJP�d1O�����鬓��?���׹��L�s��P��N���� �I��H�@I'� I?� $�$��Cߏ�5� ��K��W�v��ӽ��]�߾S��ς�:v,�M*B+���γ3�}�+�[�����j��辫�30��Ŝ^��_|�٧�v����V�w{�z��z�n��̦��z�����N��quq�@�����������9�4�~�w''*��ޢ������ʓ���Ѵ��i9yB\�*���m_s�X�>�;k�$n�eR�s4F�%���9A�*}��o��r���2�nϵ��d����>�ZW�uc�K����Hj�� ����T�9fؐe2��w��s�08}�����Q|X�%�����w�/>��C���^��}4N�(�S X��F�F�K�(2,
dVJ�"�sN�n�3��$q[i�Eb�>�G�����'��,Ț�cf��h&�a����s�ᕉ�����b��7�4��߿Sr�Q�ĸ_�1�.8��Ĳ��`�+V"E2M�3�I�����u�k\��O�d�^;����{�0}6)m��e��~5��̕v���9�������~�3���tg?~�V�B����������_�����UB�)���[���Y�k����W���>����x��ҕ]g�+F���+�ݓ��7�/��ǽ�^q/��w��d]�[Ʃ3]�;�ݮ���N��9�6�׋8K����+���I�����!=_w�'r����:����ϸ�If�<G���45n���yK�7�s�CtVj.���#M��y�7VǑg��sb�)���>��19��r��ه4o���@�r�����ֹ�r=?~�8Sxs[��WjS�����ɉ���ıF�����?p���)m��Q_�ĩ΢��ow�q��r�k��wo���!��8E������3�w�?�U��o?�%"d�LĲ�-ȕ)�]ȗn��A.M	u��3�&����7��ո�~)�w���噬�h�i�����|��7>�������? ��|���,D���VZL֍���٨ֱ�X�����w�W���lK�(Y�}��un&���>�����r<1M��lBۮ��;{����ub�Z�ff}��	d�PL��B�����������X�!&��X���6ϋ��.�N�t�N�7I��[
��l�����Wܵ��Z�Bw}ew�r��lK^ҷ��K��~�Ķ�m����Szn��E���ǲ}�ҍ�h���_�QYd�����4�h�5�DxFl6i�,l�0��	
22
��c��w��w���*љb��̻��ee�s��}>��鷵����{����c]]۬�k��I�?���ޫ��KP�ق>+���3N�R�U��RT��8�
���¾���V�T���f���O��Bw|bu3�V^J��^�.�C�ܗ_^R���t�HN����϶���}F;��r�0�"JpJ%�.��ݚ܎��-�d�adaA/#��ё
�:X�/���X0aϪ�����5��ܺ�tl�sR��B\�p�-�d�Ѩ|w�Թ�74�p��u�7A.k�.h�ei������WQ�k���GR��~��ˮQ����󾂧��B��8U�ٕ����K��:���Е����~�[�����.��\.��Y���2�7��#���b&�D�%��̓p�k������wDY(�0���`�ȯG>���Mk�l�џj^j8#6�J%Дo�de�*,�a���9-sXl���4c���y�?g7�ߡh�.��ں�����*�������G���N��8u�f�ًqgN?�u��[�L�¨��]���;�4w+>ۮ�U��ܤ�G7%��zF�f��6��:��MlcFQ����n~0�5�m�e�A�e�p40��i�f!j4�	"Y�P�TQ��F$P��E[��nDn�N���w����'0�$`���.
a20�4Q�L�Px'd�W/`����-��4]bQ��X8���~���#������޶R�/��b2FP��,��.��4�+t������p�YX���֍�^^~h�4d��������4�{��;-1�����.m8�At�ۑ+ɢ�Q-)uf��2S���dZi��\��*�kg�޹ʱ��r��{��'%3�Q(��)I�`۸�2�*
1Kĺ#LbS�J܂\#L���Lĭ#V��S$JF�����5�L��I!�p�&X!c%�FDn#o86~.7\#�km�l��5���Y%"X�1��L57#Cc"
���]������:��F����j4�r�B�Ż�y��`�F(�65
r�7w��ϕ��e-��q�q+�]Q[ԋ��>�Z���Ța(���f�p�0��W[�MV�`��Q-#%�X0�%2��쫮�f�#n�E��8d�\Ѷ�{D�nk�8�s�X�[�s[�i��0nn��z���h�乂�7�ps�8󜹤w�C3���Ͽ5��IZ4�-
j�����o,�P����#�ծ�Qu��;��uw��+�*��m&�󱹭�n&�VQ��9�G��ħ#�4ֳ5�,�a�*��U�����P`s�@����bA����4�R���[0i�Q(Սl3P�8�X�����Ț�]D�A�S��'�f�i�i�`ۇ�kM�c���Ӕ�s��~7ƺg2������ssz���������r*�[�p֌���
^p�R�w4@A�D&Ss�IpU�4�t�r8h�,�:�.�WvSF� �sf�`�Cx%��S�Vє9�tmPG{@���*A����%�# �&lټ����f��"_���� a���&�2���dfV�)�#dl�3A�B�`���%dH�K%�j�7t�[�F�ld&.�%_!.�u�����G�>Y� ]WG ��lpЗ"]���<�J��1��X��3[_�8j75�	M�	L��s{İD��olF�w�NU�P?%�-��&�k�L܆�۽�Ò��kH����k�2�DԺpL�ɂ~��q�"Ze���#L�&7WS���Y�'�R�ʖ��62�5�˚���n�WZ�8�r���jR5�ḭh�#r�l��ݖ���+`��܆��涜�L��o9�3������T�~8F%��7��ё�N���㟁�l"Pa ��������I�D���Ɗ��lbL�u��/�4�˛ϙ��ſs"z�1b5k��`�)ϯ0s�j�
�.f˘6��m+�Ѽ֮�M�(���V؉\'87z��ߵ��f���H��o��L�XŴ����f���`��0ց� ؕ)�m�܉A�Dno�O�ώL&�U}�����:��{]�u5V�ھ�<��L��ԭ>�ϕ|$ ���˽]Ծ�&��f��r��Lv����|������so�����~�3�i��knM""eەu�����N��q��5������j�A�X��(�Qpe�K�JAA��P�R̂S�"R�S ˄Jd�2	p�F�A)rF�DW �>��խ٭�[@K�����n�L�`ۼIfo���y�K�HK�y��}��?����'&���Q����u��5�����0)��W+�����I�5��1�	cR�P�R�Q�d?g>�̉�9����e�x<�:_اje/���M!
H`�v��To��M_�5x4��y��`��9	s9y�`?gB�R\�~�xL��}߻�1Rw�X�x�x�G|u�fSu���f/���u�_/�x;���|�]]5�w��Ϻ}�7j�1>�ҷ�f��P�o��7u7�e00f5Q�Z�i�|��\�����X]f�8e�ުW+�u�ʱ�f|�>I�����f}�Bj�
%,�`��`7�#a������U{����w��>�����?�>������$��B�.�c�o~� u}�$^r�83��C��^>���>|�9�C|����~�N|����5�x�:r�l���w����뮾��|r��<�m%��wWW})o>�����Wz�Z��k
��[��]k���C��t��><��t��WK�:��T��gKC3��@�#�WڬqB����Z.�M���GP�\����K��qs��4h�k��35I�����ĭ���hy���ד�:���n�s;�d��g��YC�O��9ܼ�*�ߒ�sw�դRu5qp�ٿ���!t��c�|Pb&�����5/���bTn�Ds�
~�����)u����~�f;��(,"D�ԛ�ni174�?	rH��IFRL����(�R4�)a�1�\3sM�jkc�Ԍ)0n�9iw��t}�)y˧�y%̔*�]�})GT,e����d̑�B����Ž����:�!:�p���Y�y�<���}�������~[���Q.�p�=�][�64�ޟ'#]�����w����HK�m��M�4�Ke��nNY9ub�a�C�<JC��+wz����V�V��)�3)�
]h�Ìf ��E��n%A`�pWm��2�J��	�_[A/>����vgx�VR���HpwuV�7K���5����c*X��4f]%#k-�,��˟���Ff��1���V��n\�����
��wK���Oߵ�u�����y��?�r����7��X�Z����7?	*�$5��T�>���@�4_��o��8r���ۈS5��W|��9bj�����8:��/���6%�i��G8S�?��������܃)�	l0Ѿ��W���m橭󔍿L�rF�ܚ;���FH�I��혦��&gRpVUǆUw3s��[�Z.����}ߕ��>���Gʮ�WiQ�����#�P5}��Ƭ��2�~��%�>ɟ)	�J���?��4�[�2Zd�b:ϝ�>���ߒ��)J��2%IL�>W4\�nnlnodr�ߦE.�r%��7Sz�6p�fb�ic);�!�o�s{��:v�z����#3y_}�| ����}��_�]/��Lξ�/����|��/�.�+|����[�ߓξ׻��}�0��kR0e��\�	����#�|UB9QK��<�
�|�5�7���|b��C��n��
q+���L]�كD�(����-
��f6��-�����E9�m�	tA�ˀ�4�{����K��#�[�k;�J���r�4�Y�&j��{����p�Ph	u�P�[�S|����%.���kg쌽�r	
`���~��ãL���Zt)��6r�{�
���ҙ�.�Q����w\v�9H�ba"Q)�XȈE�Tc"2ؑ2%�!�J��S�(�Y��(���S"`c7%8ictj_�f�	�2���sP�N]�{7��7���?Z	��o_����)��5?	\�;9�ۭ�;�n����dȚ��瑹��qF�ϋ\�?%��C!u��럶�3䥩�%0�sF���-3[�������>MMq.����f�Is�݁���=��+���J�f�׼��BN~;��C��z���������UUUUUUj�����������UUUUUUUUTUUj������������������U������j����*�z�0��ګ�Z�04����ݜ���ڮ�,�������{�;j]�U���Z��Y��iG<�����yP#���m���y���(@�Wg�m��av�YWc�r�õ���(��ufm�\KQs�eUX���� p֥t�Tjj��xX�p����{HT5W_�sc�?:�l� �mUm@)b86civv��j(��}���_���-��R�UUJ����o=d6��U���V۶�X�X'�0/��4n�UUQA�JJ�/U�cR�(�j�tͱ/e��p�{u'.ԥ���n�8]*��(ca�6�к�K��^�x���i��˰�(�YDѨ�*�.��谼$O6񮱞r�����xw#���z��v�<�^P�r�F7Jvxx�%\��nçcvml�d�]T�M�*�"�]u���E��&��puʝF��'�US����m�}��x��r�
Wr��p@PRpl�p X���}�9B�8ll��x��@�أ�ncL�T��W�
��z8�ΐ�UU`s*���0n�6��Q�UmN�h��iUV꺪��	�R��*�{N/r����ZW�n
`��V�Y%���.�����n8���d9z�]���n�m�j���n����m�Z2����������m�=.�l���8@j�+��blldDy���ݶ+�\��:Ӧ�ݪR�nاY�L��=��䗲޸�����v&�9�ymn��+,��::-�AܣE>7GTn�]��5LL�!�T�'8�n8Y����Wx�JԤ��*W��E]]��67�ö9��m3Ui��.XMWI���]�K�SF�m��p)�-�EYSge���!N�����V��`�k��,m�v���#�-Hl˲�.�T�9f񋭦�[P�-[LuG�P9�bZ�)�:�U����G
����E���j��j�*8s"���c5;�Z�(���a�� 5��
gdۊ]����G5K�je��v]��YĦh��ݷ��UWJ���	}��SeV��K�@R�f�n��J����)Z�"��f�]��0�gI�K*Yz���;�,��F�=�`6��]i�Ol��r=�xZ�n�X&J�)m.0mUOl���oY��6Wg��{n9��w=8ī����sٓ=Z�bU�*xؙۉ�&��MPR����������L6d�Li�L8���67#2���%��S%myĘ��	�v��r��4�.��C�T3l�+F�Sʼ��\v�]P
Pp
ˋ8!�������(wl��w��Z�j{ENdXqnU��˰��g(	r��.pA ������"Y��nUڶ��R��U.˸!��r9j�	�ʂ�d�h((�j˷9�8U�8عVBS@jW��0D�'&̰�UT�V�O+Wj��뎶�ym���-T�t�5UUR���N�V�gkds&Nm�j��l��@*��sb�A�T�WGON�C�-���socg-+�_QZ��hLʬ�og��^�uk*9e�V��i��tR
���UW.��ʵ@f��L�����r88��m�^��J�g��]�����4{娶6
��';qn*�'n�@��W�v��mU�/e#�Ij�r���3�U�2t	�U��G!s�=4=v�7m�(ۍ�4s�`�%Pe�%Z�m�ђ�����<S�]��슬�����=��v�����nzʭ����jɻ(�T�:��;[UX�(��-�eeۚ/C*֝�e66{m#UUT�K!�ET�Oj��]r���(�UJ洍��=s����W���Z��g!y�p�e�js�U+\�q)[�K+�q��Ǯ}N�u�h+>]���o[3�@�w�Vw�)Y;v�Q�	�z��Z�!J�8�;0vl7m�/4`��=���=zݚ�on[f	�\[l��g�B��Ґ�x��'
�\�Ud4��k�����gq�	]�ȆŞH��A��<�R�rEj���)���K畷Ema��kn���NwnGkQu�ޘP2U�G��ls�f�D�ٍ#��vI�>y	�/�|�TjٯQ�((��=��u�7&��i�3�������9H<n��T�K[]TT���,i��<�ƶB��!<q�=�.�ȭSm���r�WlP�����;<�WT�mG����Й���n�d��n�R���ju�N�U�W��,׵���wl1m�P���w<��[�u��Y�pW<%�s��kv��x<�\�5;���ձ\`�f��eܽ�Kjj�Řؙ�M�q�wkU��vK̗sݱ�(r�8����j���Զ�kc���͞Um�cMۜs$X�B�u-��X��ᳱ��a��n�{nuJ�lں�' s#Y�-��Nm�aq�	��*��8�h-�۪�ī�`x�R����5�;�t����ǳ����x}eL+.��h�f���\dR%ڊT�\�"UR�H���6���ݔ�8��T4��ϒ
ھ�mw�GGt���`뙓�{�C�y4Gnc0&ݲiWvim
�]K�qbu�V�[uH�j�R�uonϫ U�p�R�j�N-��Z��lm@Tl��JN��v2]�=�	!�j�*�9��B�7.,tS�+1�MUY6���,�P�"����Պʛ`�R]�j�u����*ճ��l�U�j��u 8�v�lUB;�8��#��ڠ*ꮂ�KY�����UUUUP���Vx
����T��\�J�@UUTQJ��%�����:6w��oj��[^�Ȫ�UUUW*Ҭ�M[��Fۮ�S���/RF܇P&EV��n1^j�ET�UUNWUV�+1���Ѵ�[ȵ���61��Wu�A6,�:�D��Pqʵ�V��R�UT�J�UTm���0�F}4�UU@U�WR��#������[F��MUN�ڨ*�EtUUPV6`H�6��ع�<���Z��$Z�
���,�0nKn��U]��k۩n��U٧n��ͳ�h��b�
2��PV�,ڨ�V��$��vʴ����9����[L��2>݉V��]�����(���Eն����� id�m�i6���gd���@T��	V��Un��Z���u���,�WlOu�qT��U��y���S�Ue�Z�e{1k�T
�����ꪪ�v�
�Z *.�j���t+k�S� mKQW@�;�̫�u�g��۶�j�����0t5p�0pV�@���������ks<��^=��nG��t�p\7��jYո ��ڀU�\�+����� ��ѥV��u�L2���AK�Q]�b�]YeUn�VV�8j煬v	��WӤ��tkg]�����M�ݳ.�������U�<Q��]���nݻ�uí���r�=a1:�Gi
iY@ڕC�ժ�Pmu��������D+l�Dx[8-�vڍ���+��`s��V�)�P�^m�떓;']ͽ�y� Cȱ�)��s���G�B�cMy+��}_U��E�@�j����}}r�+d5W7S��m.�ৱ4E.��ڪ���GQ�x�2�K]R&:y^��f��ӌ>f��z�a*Y�b��UU]���t�̲��T�-v�uUIPL�t���&�=�dvݭ�"j�svsi��LC,pQ�<a9�T�8㑦�UpqVyك��E)�f��`�*��F�T�Nr$�U�URMUlp&`A 檝��U�*.6Y|�V5WUT���bڸ�F�\�����s!5[.���iv%�#uTڵ[m�.�ٌRg`4�1[K-:�=��m#�ĝ�P&���﯀��u˱,�Wq��Oɷ���Z����tv�.�`뭓�ب�+A��mO�ҽ��#l�"t�v��ʫ����օ �!����|���v#M�ӄ�ݶ��N�Qy<qt���(vu�:a�2�U�tsV�l+�Z)�Ÿ��3�ݵ<���ma�a�@*�T�n�bnڶm���\�����f��띷"԰l� .�d�l�=WZ�77\���f�$�XRͺ�c�R�!�c=�a휢�Ħ7Kl�Ac �ƈ�Uӏ C��ֵ�lҭm�qUT8�H����q�S�g����*�[:*�欻   (����B+nV���c7Fd7LJҭ*�@E�+� �2����R�Tq���U*�TܣUW1�b�*�;(+�UU: z֤]5UU*�T��r��5UUK�-UW@WUY4�lUr��\5R�jG�N�t*�:+j���UT�]��������X�YeZ��ۜV�̣U@sӋqu�[t������l����$��&�[UU@Uej6�c, .R������������+�W��������U��uUT��UUV*���k�B[hT�kV�T�[��V�j@v�ꪪ����(�ɺ;G ^����Y����.Ĳ��}q�֩�Z�ST�*�UT�kOݪ�'[-[�T�{N�1��UJ�Uյ*��`�@��V�]z�݊�c�إ���eOe�C��S(*Fx�����ƭSA����9Lm�g�i	y�+�a�*��,�U���-R�T�u����\��B�)z
	��!v^�ug�[�@crp�J�%!�̪���ݸ.%Xi@���$==�g�G+���fy��$�J��s�D4i�R �Ù�3�!t����>��i��z���x%wo=N��N���]��rq;����Uۣu AN�Fpf���Iq2���Y�,�X�j��b����e`%T�;s��T�J�*�,J��o(uP!�T]����[[Jʡ*��Qr�\��ɳ��)�����KUQT-I��4kh���8j�%����j��93_����CP܇���dd ������$�Y"!	���?�H$�'!?��%� �I�	�rH`I8H �% 
ЅO��~�!!��~��$���$60#	 0BAB�H�|
B�!�#A�$�u$��(A�RF��N�)	;$!� ��I�I?���$섓�	���	�&�� �`vI� |B6�F ć  !8I'd�$���Hn ���jHnB�� 	@�O��@٩!a	 0���@�$�j@�$$��L��$$��l��$���Jt��d���I�$&��0���:�V���$`$�I!%��H~���X�!��j�	8vH}$� 0�F(�DH�A���b�$�*�EX�D`T��d"��"2)�	�	 �H��8@BI ���(��,�"��"�R�e ��
A `H��� h �&�#" 2:I:H||M�Cq���
V��5Z�P�$!Y����JM�D�I"2|K��9 J@?BI; j	'Đ#N�p	��P��NHL<�BB3� �����B�@<���I���Ȫ�����j������8����w��(Q �Z�+n���,�UF�lv#t`�W�'��7a�=	Ǭn@�`��5)b���N��tX�h*#.�is�q�x��$ٟ*;'�F�/�y�]υ���l�)�5h0����P,ܭ�hSyԜ�Cq�C�pl���]�;%��^�vz�l�G��Q��csg.Xxسϔ�M+��=-��.����[�(ˉWK���k�քm������Ź�:;��r/q��E���(�oS�6���lv�ʝ�{�м����ݽ`��X�l�l��vJcnv�n\�a�k�s�F��8���Z��t�$q����X�A�z��i+ls��N��]��cH�ƹx�A�Fs��rֺ�1�ɹ�d�]�C�L^��qٜ;]@��9��F���a՚����s��O&��j���W�g���p;Z�׹�v�[�
r{i��u��Gl�)��k�VG�P�5�knPV�f�8vCbA�t�3{\	볗�ڳ��ky�:�u���'�9��Ջ���uaj+2�ç�Y�^&���㔬��Q���vӒi|*����5@�
���
�WIn2r���S�xֹ�;��2�&˲F��F��#f�M���n�N��-�����n�jK�i��$mB�x���V��V]]8w� �l�TzV���l�Y���^6[j8�8�z�u��hKf�[ll���ڱW0�t�z&xqp�B��%w7a2k�Uv������@���6����v�b������4��\6�v�@X�-��!�R
�Y�]p�)+�����5�T��M&����md�j7mlv�`a^���6]q-��jv�$�ܶ�o)s��l���5��yn��ʰOm"Ϯum�0Z)`�M��A�1зe�X���3�xm��i�;8�c��M����tp��n�m����a%a��jx�3�&���u�`�����6`5M���VRk+5�!�NܻWW!��ĀM����4���D!��}!2 C�!�I�IBM$,�Bj��2��*kZL'Z*<$wx��e�SɇF�;7i �n�uՂ�`���v��t��z�6XQ�������CKYj�H��
��;S�����7.�v���98��*�15��MX��)Wj�M��;Lm��Y��P��8hq��ln^\��gn�r7DqGe�s���I���Z-�r�g��q��JݣuW��*�������Ͻ���f)C��,� mv���˃8v�M�)���2�y�<�q@7I���n�.��Y7n�ڰӻ���9�V�NR�v���햝:�0�J�	��G�+ ٷ^�X�ǐ�bdq�$�]��*[+ ٷ9%`�h:�[n��W`�*� �l�v\0����e�]��n��Z-Zn��	6�G6V l6^�X������uES؜\v��{���q��������i9qq-�cB0�+cP��.��~��~� �l�9��	6�
i%SN����c���Oz�����yK�����*�d�M�`͕�u���դ*������#�+ �ny�=�� '���;Ң��wL`����	6�G�+ 6/ �vn��}Ӳ��[��l� ���w 6/ �vV&�0%Ĝ^	^T����h{��麹��x�q��qVG�NJ�39�� �.�kV-����׀G�+ ��>�X�E��uv	����e`��G6V v/=�$�5zte6��e�իu�ھ���{{������FH@$5Zs�������6��[))���v��ݘrJ��e��+ �� S�nqӶ�5j���]`a��䕀Nˆ���/ziT<bK���m�����Ŕ,�u���'��1���������a��6,����䕀Nˆ����x��C���4]
�U��&�3ˋ�&�?OV O׀G6V���Q;L�����*��9��a����I���}��u����]5�+b�`�e����$ۆ����q.b�IIj\��ٕ�[��Qm۫uwlM�w�v^&�0�%`�z��;,gJ�lM�T� KK���{�~w�|�ӷ-���=	Ͱ�H����gn�S��� ܲ�j����=�~0�%`�e����@�����w��\4++�p������#�+ �n ���'N�Zj�]�������#�+ ��9��k��4;���*���$�~�OV����#�+ ;��oJ�9ʺbl�_���'e� �l� �6^�Xw�`��uv5CH��eZ5]�nYtm�;k&8@�pƍ���We�ks8?x�ﺐ�q���@v��υ�X�d�GnMɝյ����#��NNY8'6]ˢ��;m�G���3˞��ێd���,�l�D�@-��w.ގ����3�n���pP��X"�����E��u��NY��P+�^5�]�pe�bG�ɴ�2�z3a�\���kp:�w�����z��s�>.K��x��-8p\�v�{m���œ��d����L�UX;M�������sҰ��x{��	�p�	��*��jꩺn���y�����OV����#앀���z��W9m��xo��p�\0�%`a��SG)cmժe�զ�� ��>�X�l�=�X�lc�nհv���wf�X�l�9��	6�y%�.���r�n��{^�B���G,F8��Y�mێppq���K��q��z�k����<O^�X�{���>a����#[�y4;���E�t�� �l��ԁ/��pi�E������"���d.8�t �F4����Н�h$�|����}~�sj�V��7�ER�ݶ��W���	�p�#�+ &���G6V���hv��Yi���s�I?W�� =��͕�Nˆ vIN�\*��P躺�	�;�#�+ �n}��{#�Rh�L�X�L\��[]�J6f1�F\�r���R)��p�Ƹ*"�V�p����e`m� ��V vIW�j�9Kn��v�T���M�`�J��*��e`Dlcʧj�Nӵv���#앀�*��s�G$q!}��Ԯ����}�p��(eJ�V��[�� ��W�G�+ ��9��k����X�V�uUWW�G6V7nse`ݎ���=��V�ͰO,̊i'U�\�vɥ���t3�SER� Xa *XXNH+ױS���ݸ`͕�dw�G6V����t�]�'Wf�Y�.6��ǯ�V�UĒ��ǍG�!29X6Gxse`m� �l� ��p,��H�M��J���%oe\W��w6���2}	 �]wf�����)cwTݢ�j�uu�I.������%�g�9�
�k| 7�
b���\U�9���:�q��߿���]*mt�ܙuץݦ�"\�j��Ե����?������ [���
�k| -��t ˗%hN&)�L��� �l� �������
�k| >y��(�X��Pc�&�o�� ��n�V�[� [��t|��,���y?"H� {ʷ@+}�� -�ٺ[�o��u"`�q�)���o�� ��7@+}�� ������I'@�"X�I��5fa��p	1n��Y�f�A��vc��fC���7i���y�3jU.1Q�Iټ�2cJڔֆΨ�<v���#�R'&���h�+���n��/L�y΋nSg\gv�6ɮ��h(	n��c�(���{b�mN��ݰ�̍�o�.����ܧ�vK8v�h�����źADkq�j�:��mi�7Hc����|��j�s�\vט�߯w��>�{�ﵾB��\��������姘6\��0�������h
G�=��I�������� �����ʷ@+}�� 7��A�Ԋ������ [yV�}�� �l� �UHg�q�1Lx7��ʷ@+���ڭ���[�ۋ��l`��)#�n�Weg �훠�[�oyV�����LS�� �;f�n�� [�U�]�� 5�nY�������V�Ե(�ݮ�7ͬ�N�����]/\V6,�X�(1�t�k| /וn�V�s?��s2�}Ӿ�9m��x�MWZ���j73Y������^s�! ����8V�� �-���[���]J46�4ҟ�"� ��� �;f�n�� _�*� >���D�d�@o�{���
ݭ� ���t�k| �w
�lƤR4�$� ��� �ʷ@+v�� ��f��?v�Ŝy����1���km��I�]��V�����`{G&#�JU�ͷ��'B6�iLS����yn�V�o�{��t�k| ;s�X14� �$�t�+9�Ͱ=r�n�y�y� �ʷ}�31���@�N&(ԙ	� ���[��,���lL�3��FSO�W��ܳ��BYϧ�,�D#3[�,��e93E1ct�/�W[����a�e�{��I�vY��c�\��h�5������2��dO�a�]g�:�o ~ٷ(��8r��D{9��ˮ�4��fjY�ަ�z�&nC�hszK��Nf��2d�u6�]�1>фȂ̐�A1�	#2G"���dd�h����x0I�&e�D$a���I��A
HZDQ�Q�r�
[��0\�
1���X�sQ!�� ��4,��Ð�jC��ɇ�6L����t��q6s���+%�0&��T�cx����Fs�1-���~�f<�`]�&k@�/ ��O�͟k/7xrj9��'3��g�~����F��KD��6�$�p�I��>��&��bD0b�
��Nä��!`ja �I>��t���f�}�����r�u�ݩG�b�c��ǎM�
ݭ� �[��]��߳?f6�r�n�tk�{��8�!�� �����Y� ��ٺ[�� 긫��u�Ki�j}�.Ɗ{u�����b�9�uk���d+�ql�l[	ѭ�w��]�� �훠�[����[���7@�y�	�H���� }Wl� ��� �����[�6�����#f71���t���� �[��[�� �v���T�p�nD�)�F� _��� ��� ����u�[w8O!@ID�	���i,�#T"H�Г���3�w���� v�|ѳɃ�9���[���g�ٙ�z�����G��{�Ř�z�����U![�Wh�L������rrQ��v�#a]Z�����n�x{Qp���7� �]�t ��� _��� ��� ����1D��Pc�&�]�� �[��[�� �v���v��pM'1 nG��n��vVp >��n�� �:�&��D�ṛ��Y� ��ٺ Wl| /��n�YX�1L2D��7� ��ٺ����=�� �}���
ݭ� ���>0�D"	$��^�k4�sN���3kZIvn
�b�.�1)��K�����-�l��Lr�&�6ʽ�w]�#cU��;� �l#v|�xἠM�1�,����6`������%�� �s�����u�j���ϑ���n���\m�z�0�&U-��Z.;.:+����ӱڮ����\��oU�4�/�gZü�[)�M���iGj�n�cCq���a�5u��2'd�;y�%����Jd�ou%L���tWr�8�H�����>\!k����E#��c��$��%� ��> ��n�V�o�{��t�U��86�L��1G�����
ݭ� -�ٺ Wl| ;s��ɍɃ�9���[� [��t ��� [۹� e�+�jG���7� �;f�]�� ��st�+8 |����F��Lc�&�]�� ������߽���<�<� ��7@���N�^6;���KI�f���e�ƥ��m�[�����p�A�lb��6���فF�| -��� ��� �l��߿g�0?z> �����D������;����O�H�����-���� [n��?~���O'��(H!��� {��M��c�m����Y� ޮ�\���Ġ$� +�> ۹�]�� rٺܶq�m��&)�D�� ����
�� v�ٺ Wl| =$��O��Ԏ��B� ����۰cc�ݼ�Iɥ�"1�.Li�ޮ|�Q���t�u�WwV����W��a���#�$ً �j&7Et��һ�x��xʑ�lŀl�ֻ�ۤ:�Ъ�.� �R<I1a��]I���K%h���jY�2	Ekd�@H,�#ȣA�0$�75	�����{�l�KL�D�R&���7$����6T� ���l��+j�WUe݅�UV��#�6S���#�$��Ē�/6����M�S*��ЗEb�KՖ딆�v#�\�Tt\�l�ͩ?��(�-I_3�|Iv�N$���\0�5J��m���V��� �R<I1`*G�l�����ڕuN�T�����lŀl�����6T� ضRQj���i��լeH���V��x����D�C� �����xm^��W��N4�HL�C�.�v�$�]�I���x�\�in/*�5N��=c ��P��Bs8���nݪ�׳��秕l,#��M�6d1n�߀��� �f,eH���V�[#n�h�t�uV�	6b�$�M���<z����w��~����rG;(2m��6T� �Oea�s��<ޞŀN���L"Q��Iv�����v�IMً�\Nz��TC��ӱV�T�Uu�l�丹���~���_�<{�gsj���"$�"��`�2
HE�>�[��9��3��ĸ�S�>h�7j�Տ4��i3@�H]�rx1�U��3�i1��\��A�oD3��q�)m:��M�Oj����jP�a�.;w�M�>.�UѲ��zTm��.��r����5�J��/=�����Y�|�8�x���\u���ZJ�1��vvܝݶݻ3)��a�aXs6�-�Hq:W��+�N4��3����S�v�Ӳ�	�B;Л��f9nL�u�&�a�e>Ϳ������F��&�Svy�
�;pl<���g�ۯ����e+E�c�~߽�ŀl����{����}���;���Gr��eH�ɲz�z�	���7f,��>�v��ְ�Z�-��w}���<=��'�`��<�wbe5e�V7UWXԒ��*�������ذ�#���Nz��`j{ͻH�e;@�U�M��qO_��z��`*G�v�����d���ያ���٭�\��2�;��N��lë��(l}�sNS$WeJ��|�{� �Oe`T����=��gW�S���c#�]��|8�Da?�E�j+����(�%L$Ԑ=!�}�?~�W��`T�<�\M��껻v"��j��u�{��<M���8��߽^��=�'ۀN�i;�nb�4�xy���/ޞ�`��<J6V�I%�=~��'�ﴷ�8��r��������y��9���] ��߯ �f,�1�J�#ӽ"��v��GTju�� �L�@؅%&]����)\/�{���|�������D�`�/ �f/.qs�0��y��� vSV[UaCt�� 6Iy�ēg��b�'��x�rV{��l�S�n�4c���^��}��=��o�B'�B�Y$�� �I"$BCP B׿��f�}��kj������jڠɶg��^���������^�ğ��|�o��I����vS�uo ���ys��{�������w��_{ݑI�_3�Q D���\=G-�mvX�6I��H�5VEM6�/�g�<��ӓ�.jF�K4-��߾�����~Is��Հj���C���"���&�Y�q&���� {�z��{ןO-;����8cF2��p	��� H�^���/˜�=����?~�����;6�vڱX���y$���[U��m^�������"2P�2} I�$���~���j��{��K-�V��J��d��~�I~��_�{�W@������e���ݔ;t�ђ�s����j���l2�p��ERU�>�y<�&ymC��v_�}��,eH�E���.q|���� �+�O��Ժ(y�g ������<��h{�z�{޼M����8���~)1ͫ⦺�� ��ߞ {�����O%���,z��ժ:���庺MSmU��ė?..r�߿~���~ŀl��B���ǿ��zc�������u��$ً ���/�%�����������^ Чs�Э��S뾾b8qV�?\N[�������7w�P��S�����7D�>�5�+�Dl�s�5�cl������aJ3�Ս+,BX��V}��iGe~���]��7c���d�]s�8<C�I2e&�98�`]g%ERn<���[�ɒ��K ���怛�0ݤ�t2,��+U���H0��� DC9K2L�+0���$� ��Ob���p*P20�cA�U�DQ�k��SAX��6UDa�&���DDb�$A�<�y�L�5\�57��!u
1�,�liAd��C��亊(�H��2�\���j!"(�����s+��h�$��#��|9�����Oʪ����m�T
����m$�M˄{]f��7!D���C�w]��`h��u�öu�:7b��sS u�vSp(���l�eW#�.�^��@�є4�0R���q��77h��]���'U�9%�2`�e��p�ܜ@�f�MhJ*[[4��� �ڀ�Y}�1�\M�緳�{]����0�vn�Ɓ���s��5��n�.n�X<o`���g"捣�=�hWl�	�;3����"�9g ��vk�g �*\`ī�H���[�ִU�6����K���h��E�7`��qV��DO3ۥy��^Ƭ{8R�HP��/:s�+�ڞ ��gt�>u�������+=|0����8�)���z�����N��u��.����/;�EۓdH�ɇ�]\��>mr�s�Fu��p��0nwV����pm6��(��;�9�9��8�g���t���}�Ts�JJu�;u*�ݫTư��"ҤBͨK�'j�nQs��u���;`ۀx�ޗ�ێv؜A���4uq����`h�'+@5"^k�tz�C�ӽ���ȋkc������1�:�ۖ�����k��-$S�+&D�h��Z�w��[�K1�s��5)NevP�y@smd�wSg�va3�Y�H�8�����C���筍v�����Ls�YQ7S��'���[F��b��KvAg�rK
��WT�8"ih[����ܨ��������5��6Hrz��k��+v	i�\6��c��ग<��̱�
�ܯ6��1B�0�N�,7&y��n���U�f���\)�v��)��^�G�T���6�Xh�V\9��6CO*q6j.�da4��$�7U�҃ �|�uR1s��Yp�8�]���������Vs�X�x���Z� �Z*tN����O�c#�� �����<P��h��ls��s��g�dA��R�z8;9�=��g��k���2/j�����m�U��V��S�h�箜o���(���5����WY�@��O@��$!�6a		�􄇠t �$p��� ~�����3��kY<�wg�l�:8��u\lsCr/s�
{�VcR+�x8��f΃DV��k�m��n{AgYm�Z[�ʹ�{h�3&���}��y�{�Y6�x�9�n�t���`�����T3���GN㋛ev0�4��4p�n�$���M'BmӴSՍ��Z��%�*�۫y�n3Ԙ���<[On����X��Bk�,+�cK�]8h�u��4d��C�!�p����[lfY���eR�Q�]�f��W�E��Jͷ\,g���Z�1�w����?=����u�M߀���~x"���#������b�=>���kv���sx�����Ii=^��=�{��y�٭l��݊ڥ|�)]�=^��$���\������������?Y�aؖ��Z�k�x�8��{�OW��E%�{���\��6/*����]�*����<���sǽ=S� �&,l!N���ӌI����:ݍ�#n��[��6��;b�np���:��6��y���,�g�B����=��6VǀM��q%�.s��^��ޟO�˗x��f��������	@�b�`�H
�Ydd,��r�I<��{ذJ�� v/<�f�*��umJ�Zn���{%lx{��f��<�~���{�yF.5c*�3�����\���=x���~����W�����O����QM�b��� t�� �K޹���{%lx�u��u����0�3[�F�$TvV���csZM�X:N<�?���?s}�<v�Jj��z��;�%l�\�丹��x����v�Wn�-Z
���N�Ş�\I�ީ��=x���Ĺ�OO��-�1����ۿ^����m�I�$�5�{7�}�}�j��]u¥35��]:�]��?�'9[��V��{��'vb���K��{���?���l�rQYcs���D�q.N��|�<��=��}�M=n��A48�Y5`+Zk��R!3�N�Av�|�iWW%�ϧ�I�ɹ�*6L�[����X���J{+�$��=�x~��R�8T3-�8{����y�8��S��z��;&,�Iq6y{���H���8��|���v�^��\M�}�X�{� ��g��[B�l�WX�?s��������?O߱`*G����� �A���`�A%�^��{XZ����m]ۦ���Uo ���s��9��{�~���O߫ �S��w��w6�Y�X2͢ۉ�O:ru�̓j�ui��]��J��s\nE�_��{�����ٱmь�f~�o�������}��o�!�}�{f���u�
���KHv]��;)�Y�.~�8�9T{�{��?{߱`+c�qq%��t��wv�j�����=S� �&,=ĸ�����o��ՀuE[��um�U�c�x\�I?O{�OT��;)�%�$�y��}�a¡�X���������K�8�'�~�]����Nɋ �ۤ��k]�v�<�t�⥱c�ks:c���D�%������HŃ�Jk��6����u�6ugvw>�
=�b����9�ܝ*��ڂݞgW�(��I5m%�p$�g9Ea����3���
�n��.z�G8qk�v��ݭ��.��Fښ�n�s�y�Şs�S�������ݮN��a�<��#� �
Y�u�ػek��m�JdZi�vy$f�NL7b�潷>�I�k�X���mY�c��N��ڮ�6.�~���o�UٸF�l6�~��ՀIR<wf/.$�a�W��ޝ�%f�Й�\�����	ݘ�	*G�})��8�ֽ�-�V�'V��U��=� ��x{��o��߷ ���׀{�7�t.��h�K��y%��_���9��$�����}���%����Eo ���p���_����?~}���%H�L['Y��v6�LI���*P�5W[Wna4g�#&�VHRU�]��xs�'2�`�6M�]��S� �ً ��?.q|�_�����s��V�j�Z�;��Nɋ2I� = Ǿ�r�^߯}���s����O�I�����vf�kZ]h���h��_�<�mK��$���y���Xg}��b)�������<�߻�x�{� ���Nz��F�zʦ��
��:��eH�	�1`*G�u͗xZ�Ԫ-�I��b|l��,�=�81�:L�-�Ɋi�]�_T&~��!fxk`��k��{�' �����l��\�>a�W��ꨫ��;jӰ��U�J��l���z��7f,�\K���/�&&��C�;.��_���kj����n�I# *Ȍ"$��$I��� rI&�s�I/��{���.��찻��ww��%�q�\��='�`+c��y������/ �}7g�M�ұ���	�1`\I)��ޯ^��>�;=��#���%� x�m+*��$��Z�	��\��s.&��t<"�R1� ����Z�6Vǀu�R����s�/�}�~��O��m�u�΍���eK�qs��z���Ob�6Vǟ��~�&��}���Cl�L�v�^��}��M����I��x�y���b�wm�t��[WUv�=�.'�O|�	�x���[\��M' !�I����v��x*�Yi�ZMլelx�^��<M���^T���,�Tժ�&3U��+�cXX��I:��Ў[�MuNl�yW�<�p�R�WCB�������<elx�1{�I|�z�� ul^wV�8�A
���{�Ϥ��O��ܜz�� v/?%�~\�*��*��;�Z�l�c�x���ʑ���f��<��^�ޓ��fr7E3\�������� o���6T� ��'}�]�v�k���{׀}�O_����b�6T� �ė�k�Q�~�3>Ѵ������ku/%�`��m����j���\����[��cے�.�B��i��<-�`�d툘�iCjk13����r��.n�W<�בM­�N8�ggw�qv����8���Շ	ඃͺ���x� �-�c�5�.��ZY�8�5 ;n#�+�G��F�kɸ{���ӷ}�fg��S�hyQz�g�*��]�=�y<��9o?İb��s�zzݸK9w �X1�J�ku�*㧌�ڕk�$��5��:!i��������b�6T��$�a��`I��;���WJں���Nɋ<�I�z���z�rJ�7�l�S��PZN����x5Ix{�\M����='�`E1WeН�
����8߷ǯ ��ՀI&,�I~Iq*����;��W1V�-�Z��=����}�%�O|�z�� N�^��(�ʥT����m��Ŭ���3/7Z�܊WX�4��2.��/�f%u�R���~�~����v�$���~���Az^Fg-�8�ټ��{y�����i&�4Y$��s?�	��0CF���2�1,$B Ysr�,���H�B5��8�kj��w�6�{������Ii�������]�Q�֮�}��kj�{�so� �Hg��{�x�����l�޷hm���2/ �6V%lx���=�s�.&��=|���>�B�h�컀w����s��%=s��O�elx|�*:��1��z���]����f4WLK���m��լ˙�[X�&�������#�pԀ��Y�wo�'�y��%`+c�\K����^��=<{q��V�*˫xz��elxڑ�+c��I~K��UA�O��9�R̶�.�����;��m��KMk�2�%��;k"�� d&�d��i����t~�h��~���ɢ��'�>e� "#G���9�?D�����ߟܤ0a�����"�u�'�H��9����0H$�XF�9&V�K���6L����da"�Ȋ*6#&##Y6hnHe2�a�5Ȕ'䬒#L	@������` ��	H�ңh�Vr�,@� R*.4E>��H���%u9�Ej����*A��Fs�	�Ղ��(�%��ɨ�'�?_����X��>��$�� t�!!�@!�C�'H�I��������N l�&���l�2 C�!3���~���� ����Ѹ�sSh���=�ē��� ���G�%`+c�"�Q<�EՀղ�uf��<ˉ%���W�OT��&�� �b ��b�;�v�y����躝[��ڶ�����i�Ț�����w��}�E�Tn�h�`���V��<n�?..s�\�;A���׀v�}�Cl�������w��Mۆ��x}RV{���l�S�ɖ���vݺ�x��ʑ��������s�_�_�V�����7�l�S]�n��;�ˉ.q�_���{Հl�۵��H�H�BL������{�%����W4�5v���^���$�w����OK�l���$������YTT�zp�����Ukn=d.U����nz��P%����'�x������5���W�<f�0���%�%��ǫ �}7g��X��hҭ��ק �����	X���ˉ.6yH/'���V![(�V`�<�}��<��n�x~���;;��!�ٗms�x��s�J�s���~�~x͸`+e����]�t#4f���w����s���}���^��}[+ ��s��</��C�w'7�b�y��.����4p9�A-[p��V���D�`ݱt������Ȥd�ne{dĵ�M�M�n*lYM��\R�B����"�v�����*�5f`�1�*�PՄ.�j�g`m������;v7F.W��r�������b��j�����l�b| qJ#�7$GgRBݗ���W����[�:��[��t|,�	�T���.,@Mq�E��1Fpc��unq<�����v�#ZX�{���n��q��V��:�p�?_��6Vǀk��X�����*��Zcـl��=Ēl�W�X�{� �ۆ{�$����T��|���Yuo �W�Xʑ��ē{�~0	��� uv�j�����M�wXʑ��p�6Vǁ�$����n�>��ḪgGh������y..O\����elx�L�N���p�F����Z���ﭏ���+G2�.�\%.h��ܑm˵�Ft6|�O<_t��l���K���}�b�>�t>��&���vo ��zwr�L�2�4��P�
BĆ�!�	�}��.�����j���n�:wIt���`�R�UE�%lx�LXy.$��O<=�� �[L����aN���ˉ*���'�y�����$�����K+�&�m����X������eH�	�p�'�:qnTi�rYK*E֒4�l<'����y�S��5n9l=/F���w��}�1ѹnaV]��=�u�IR<Ip��K�}����އ�fL��5�n���e� ��<>�u�I$٫�O����te�x���������"H 2H� I� �o^�߭`�O<.��`�R�Vʱ՘����c�J��<�O��� �&غ���c����{w ��<����?���~0���|;��;����l���V������W]u�J��<K6��*Ci����5[���ǀI&,el��\����=���{��e�+C���N��6LY��q&�����ΰ�#�>�U
Lv�-17V��#�#��Xyqqs�������b�'ap�ƭ2��
���/�B����f��޻W��vmP�!'��{���oj�K��!�r���x�\������<�R]`����2�a��0Z�S�<Ɗ�{>&��<Yu�v�ti��O$�����mj�[�luo�=�_�eH�	ڒ��D�*���]���Ϸ�JS)���8ʑ�������?J��� �����I�?qs����U��ߙ��:*�U��Wo �+��eH�	$ŀl� iއFm6��ѡ�����^����}�b�6T��8��~��~���X��ߓn�
�N��6LX���������w�ͫ�s��W?I ~d`P� ��H����ֵ�f�3sXb��0:�m�\���4��!B�
Z�f�2J��'cs\��5�sh��s��]`��y%�ɟS�`{i��pW0���:ggd�᫮Gъܽ���.P��e���c�m���<e��J�lC5��C(�ق!�-��T��!��yt%����\B�nؐ+8q��ٵ���,��^U��ͳ�BN{
�^u�A��*�1[6����HO�B�v�5n\GS�F��dY4����I�Y�'�y-���b�x���CW����eݴ�n���_���Iu�l�6\0	�\)1��ul
������Y�.6OW��O_������%��N߮nŘc�1U�z��M� �%�앀v��8��1��7���K�~�� >���X�s��%�����~���xV�+whMZueU�$��G�V%H��q%r��y�~�1ł�!�5�)��VۀR7���v���D32R����nr��cR$����MIx���K��q%{d?%Ĺ�qv���߯ <O����UR�]+e]�`*G��\KWV�Ē�$ɋ &�x{%g�l�^�wH�հ
���z{ذI/�.7�=��=������P��eݴ�Z�����g����`T�ˉ���� &��R�VU�c�0䕀~\\����{ذ	%� �}jEe���CV��9�G���i�˴&�s�h�+�uf;s��m��s�/6M�0�Fb�߀���׀w��,Ip�#�V�V�j�����jձݼI1g��d�����z��;y��Z}=��F�Fe2�߾|�^����p>A`C� HD�b �2H���^�n�^{�����e᮸c5�AT�������V=^��$��LX�`B�UUJ�t��Wu�l��./{���'��XrJ�:Љ��˺T��+B8Ӡ�ut��S��Gv.���td��a�{5�V��;����!Zn�������l�=�p{���?{7�t���t<*�d�g�s��*��߿V�����&ˆ N�Q�h�Un�;ـG�V��x~\\K��������=���0�VZ�n���(wwX��8��x�{� ��]v�!�B2`AI �I%��<r���t��٬vf�F4wo �R<������s߿}����~�eH��И�l��*�ꘃ��UM�!x��;m�[�ݰ��F��Y����A��p�l�j��V��b�#�V��~�9��C��^����۵c5�mvg �IY�.&�����W���b�˜\�:{�|2ͶB:4�w ��� ���������z����ۺh���-�[�$��\0䕁�Kߟ���ٻ7Ɩ�9f`A���\0䕀l�%H�s�����7nC�d�H��X��1ns@V��t!D)n8��O��AX"+CSiM�(��w)��Y�n��K��:e9B�c2Ќd�䀖F܇�ѡ0�HXoq��a9 $�VC�H%�ѨR��9���,���2cA�,�������K� ��,C9�Sm���ƈ�Rc�q�,AGlȰI,�����úֵ�kUUUtUU]T�Aı �&D�ݹ��JW����+�r�=6�C6��E>=1�&ry��ؖZpA�:�ۋ�NQ���t�5��ܭ�JF��n�!n����[������0t�5��97O)��;nͶɋ�(v��=�f��n��sQm۝�9�k9��s�_%����KGsp]��e�4�ݭv��`�k�%kfX�a�]h�s\������ {vs�1�99�]�'���� n_<]�����r㤕u��ۃ9�cte��Xcp�9�]ɞl��x9x��u��<��W` ʫ���0��ɹ�ŧ*.��n��䎹�lF+qū�'/l����CA��`�)���FR�ma.��g7&z�P+n7\�X"n�#��I&�1��g�������1���1q�T^M�7[�&�dp����n!�
�L�3nG;�Z�i��Lu�1(F�:���������mཋ�7Cz�n��D�mQ����U�+�	SW����1.����c�׭�y�vRs�U��%��A�Gj�Z\#
u��`}X�Ϟ��y�e�-G��mr	j�[r*��A�w"ļ�w&��̻�6<b�؍s�5�Y$�ní6�b�ܰ���
����@ �WOm�F\��tD�&�J殻m�ٳ��d{��ce6KA��`6bG�v���pO6�u�3����m�:�0��ƃ��{�V÷��=R� �����y��(�b-͓������Zz�ږ��wb3�������<�-%��'�2�%���x���U�-Ɖ��$����v��tΩ�Jg�l��eri9� �����׶�٬���۷S����B\�l��nî�KkŎv^��!�t�[gmi���3�'���Ju�r��%�6Wv�u���D!M�}�9�*�Cqdr�MK�Gh=6�|4C2��t��vG �3�e�����
baU�ؗd,�v��SP�p��hs)����tPu��\˧v���8ͷ&%ðΣ�;��䓞y<��H2r~$jBvHC���Bl2B}8ܐ$� 6C��BH2I!H �:/���4�֌�et���;�8mP�\�=�����ⴗ�����v�v9�koi%@�����T���7�`�k.]Ip̪�s,������p�-��$YB�S���f�"4�:��f�R��f���w%�tv{8��b��q*�;c�Ld�ў�r׭dK�Ȇ�l���JZ�r��7,ؔBݻ��:�stٮ�{k�X7� B��hٽ�h�C�]i̶�Q�ܝt=���0�m������Vɦ�疿=�w�Ǳ̫V6�vt��`*G�IR?˜_��A�߯�z�-U7N�wV:��eH�	*G�l�9%g�_��lw�o�͕.Gҭ����� �.rJ�6T� ��Ⲭ�l�j�ʫ0<������`*G��������~/M���kT��J�6T�<���&qzL�_L�l+���q�aXV�_{٫������xm	ݍ�F�g��]{i�
��ڒAf���|ڼ�K8�N\c2��5����+
þ׽w0�+
�����aXV�}���8°�+g��naXV��>1t:�у����8°�+w��q8C��i��V���p�
°�?g��naXV�}���aXV�~5�<�u�f�E�F�N���aXw�ߝÌ+
°�}�f��!XV���q�aXV�w�p�
°�/�{=cjf���M��V�a����Ì+
°��]Ì+
°�{�;�V����V�aߞ�g4f].��M���8°�+�]��8°�+	��~w0�+
þ�naXV���{70�+
�����R�(�z�x�u-�=hհ���ck`�aE$���,=F�)�J�E��\�y?Jy)�X{�ߝÌ+
°���V�a���͇�'�°�=����q�aXV���w�Ӛ�Mh�i�Ӹq�aXV���p����V��f���aX{�_��p�
°�=�w�p�%aXV=�߫\ˣF]c�usF���aX{>�p�
°�;�{�p�
͓h	�>a����p�
°�>�}�p�
°�)ߎ�a�c���]�k70�*Jþ׽w0�+
��{~w0�+
þ��naXV����naXV����5)��]:����V�aｿ;�V�d���V�a��}��V�a�k޻�V��������F::zei:2���In0֮\v�<dpWD�g�0��j͞�����;�V�a�{�70�+
����70�+
þ׽vN0�+
��{~w0�+
�����\u5��74naXV����nd�+
þ׽w0�+
��k޻�V�a�{�70�+
ÿ=��h̺�u�t�f�p�
°�;�{�p�
°�?{^��8²V�}�p�8°�+�{��8°�+�맵n����F�֮����D1�������V�a�����V�a��}��V�AM�cY$�;
VlkF_D�A��{�d75�� f�;�c`���T,�JH5"�a(��'d��I�>���ٸq�aXV�������p�tj����aXw��Ì+
°�w��Ì+
°�{��Ì+
°��{�p�
°�>���&��1�=�͝��ـ������z3��睵�뤂�����<��Ռ��F�s���S�O
ù��70�+
ù�{70�+
����]Ì+
°���V�aO|w�aSZMWU�kY�q�aXV�wٸq%aXV���q�aXV�}�p�
°�=��p�
°�/���i�M�h���k70�+
��{~w0�+
þ�naRV����naXV�s��naXW�O'���3���(xU9��y)�+���q�aXV�ﵸq�aXV�{ٸq�aP+}���8°�+��4�ӎ��3F���aX_w�����aXw=�f���aX{�o����aXw��Ì+
°I?;�m�e�]c�t.:�k�:U�L��Yns�KQ<�3��u��r�v�3���(m�Wlt�����7��	��=Z�ݞPn������)t��d����Y���q�\��(B�,�����#l*`r�
:���F�1�A�jӞƺ�[+nk�p\ V�+��Ζ�Y3�n��#s/El�ab$x����W��r���I�U�����'�K�9���;V]6l�s`+�V���j��k��XvĊtn��sx��������k[���aXw��70�+
��{~w0�+
þ��l?�0��a���naXV��x�ut��.�5\ַ0�+
��{~w0�+
þ��naXV��}�naXV�}�sp��I&Xc
�����]kYm�ѭ74�aXV�����naXV��}�naYI+���6�X��r
Aa���v[��r桴���/��kp�
°�;�{��V�a��~w0�+
þ��naXV�;��b��MtSX�5�Ì+
°��naXV���z�aXV�}�p�8°�+����8°�+��L��3�E5itڵ���.��z�Y�vvv�ݱ�B*�c�8Sr�V��覍\4`幭Ì+
°�u�]Ì+
°���V�a}�{[�V�a�{��8°�+�;�<�sY�ӭ,u���V�a�{�7'�0���a�����naXV���naXV���z�a��aX_��9���u�3ZG4�h�8°�+����naXV���naXV���z�aXV�}�p�8²S�O'g�/>f���؃j�<��%!_�!�3�����8°�+�k���aXV�}�p�8°�+����8�)䧒�O~�F�p&f�j��~!XV���z�aXV�}�p�8°�+����8°�+�w��8°�+��_<ю[K�Z�.7U���NJ��b�q/����;B���=��u��W.�v4�f��Jy)䧓�����p�
°�/��kp�
°�/}�kp�
°�=�o����aXz{�9���8���y?Jy)䧒�߾w'�@�1�a}���naXV������aXV�}�p�8°�+%��w�	��ʚ�y��y)䧒���}�Ì+
°�}�;�V~����I,��A�[
ŋ�,	0��B�$��%(1H�@a�e��
AY2A@`
HO�Ig��{���70�+
������0�+
��~�n���34in]k[�V�a��~w0�+
þ�naXV��}�naXT?��3�������a_'�O�o�Å
�<��%<��R���p�
°�/��kp�
°�/}�kp�
°�=�o����a_'���6��an��6R�x�e�%��9Lv��E���d�NxLT��$�����G9�3F���aX_w�����aX^������aX{�ߝÌ+
°���V�a��y�.���YGV�Z����aX^������aX{�ߝÌ+
°���V�a}�{[�V�a��wɫ��u�6�Z�8°�+w��q�aXV�}�p�
°�/��kp�
°�/}�kp�
°�<w�m�]b��2�Fi��p�
°�;������aX_w�����aX^������CRx$@ d�`L3��Ì+
°��U߅˭k3.�a���V�a}�{[�V�O� �������+
°�����Ì+
°���V�a܉��}��f�&���mյz3��n��K��Ʈ�j�s��i�xw*�L�M�FX���'��O%!X^������aX{�ߝÌ+
°���V�a}�{[�V�S�}=����1��!�W�Oǒ�J°�u�]Ì+
°���V�a}�{[�V�a{�{[�V�S�����G-eb����'��O%aXw��Ì+
°�ｭÌ+
°����Ì+
°�u�]Ì+
y)�w�}�Tj*�K��'��O%aX_w�����aX^������aX}�{�p�
¡�!8����ߍ���S�O%<��ߋy����*�6��aXV���naXV��׽w0�+
þ��naXV��}�naXV�C�$`	2(�!��P�0FH�" (��������љq��u����Q�0������l�b�����c��8k�5v���װ�f�:�]GSk��-���3�kO�oy�0�����x���:�Wl�u<�zk�y�\U#�,0М�&��kdVa�=�l@�v��GVt�N��NF���Fx�b�(  �v�@��ٵ,�u�c(V�e�6Kx��Kר�ۂ��[3�x"%_*E���O'�G�<�![x7e,j]�vV���ws=���M/f��x�K�R���E�����+
°��]Ì+
°���V�a{�{[�V�a{�{[�V�a��o�ut�atf��]Ì+
°���� �a�+����naXV������0�+
��׽w0�+
���W~�f����usF���aX{;�f���aX^������aX{������aXw��Ì+
°�~;��]WN�h�f�p�
°�/}�kp�
°�=�{�p�
°�;������aX{;�f���aX_���m��h�.��Z�8°�+w^��8°�+���q�aXV��ٸq�aXV����q�aXV�]�3Nf��o\`邘�Q<�哓j�5�n.�W�>�<�\p��i�L�5\�V,9��~<��S°���V�a�｛�V�a{��[�V�a��~w0�+%<��g����.g<��%<��=���p�x�"�Bt����58Ì+�{��0�+
��w~w0�+
þ��naXV�O�6��"�r�n]�'��O%<��^���<8°�+w��q�aXV���p�
°�=���p�
°�>�Z¬��m�y��y)䧒�O��>9���aXw��Ì+
°�w��Ì+
°����Ì+
°�������-p�5�3Wp�
°�;�o����aS�H ��{��7�+
°��������aX{������aX��O��7V��5��MV���1�z�4m0n�:v3p���mtb�9/E�[�ۛ���hu��i�?0�+
��=����V�a{�{[�V�a��޻� �a�+
�����w0�+
�����+L�JkK��Y�q�aXV����q�aXV��q�aXV���p�
°�=���p�
°�?a��V�fsF�YsZ�8°�+w^��8°�+���q�e$�y
�������s3����P)����h��X����¥n�m���[MT�$���������E1�������7.��ku��A�L�e�	v���f�p�2]ƍѣc[�ѹ�Hj��2�8!5��*��ЊĊ9��"Q!C�+$�1a���B�F��[Pl�),b��5�Eј���+nŌf�L�`�C(��8�U�&�0vn<C$0e���S��hP5�X��j0ƶH��	",�9I �� ���D AHL���! ?@�!&�I�@'��'d$����;���70�+
�����0�+
��N��9sZѦ��5w0�+� !�=����p�
°�?���ٸq�aXV����q�aXV��q�aXV�|o�
����L�<��%<��S��_z�aXV���naXV���z�aXV�}���8°�+�;��[(�%��)4T��������H�M�7\v�W��h��,
��]����P��֮���aX^������aX{������aXw�ߝÌ+
°�u�]Ì+
°�y�<��u�Z��ۚ����aX{�ߝÉ�$f0�������aXV�����w0�+
�����0�+
�����n��ѭ74�aXV�}���8°�+w]��8°�+�w��8°�+}���8°�+�'���V�p�5u�p�
°�=�w�p�
°�/}�kp�
°�=���p�
¡�X���,� ��L��߸�aXV��Ӿ44ˣZ]WZ֮���aX^������aX{�o����aXw�ߝÌ+
°�{�;�V�a����{Zхs7�m�����܍sec�cN,Z�1)�9�P��L՛B+B�����-W�Oǒ�Jy)���o����aXw�ߝÌ+
°�{�;�V�a{��[�V�a�N��.cr��n��aXV�}���8°�+w��q�aXV�ﵸq�aXV���q�� �d�������Z�ɘ)���䧒������p�
°�/}�kp�
°�=���p�
°�;������d������}5˶j�uY�'��O%!X^������aX{�o����aXw�ߝÌ+
°�}��V�S�}����B�ٖ�^y?Jy)
�����aXV�}�p�8°�+w��q�aXV�ﵸq�aXV��d	���`�D�dK����	 �0d� ���{o{�w{������oĚ�Mj�(�ڕ-��$1D���E�۷GSϛ]#�4#�GT�p-5u�:�v8�\�l� +dh	�v��]XB�l�p��y�J핯Q��h88��lkfy�ڵ��f���>�����;����Qs���\GAF���Ѷ������[�����p�j�VI������s�R�82��/Hr����N:�j�N�fpP��j��$��O$fCrQ��4m�XH��G,{]P]cxs�m�î��֊��K/;t۪�=�И]�sO�|°�+���q�aXV��p�
°�/}�ka��°�?����p�
°�?���O�:�պ3]i�8°�+w��q�aXV�ﵸq�aXV{��q�aXV�w�p�
°�/���i��Z]WY�70�+
�����0�+
����;�V	�1�����p�
°�=�p�8°�+'����J�8�Uy��y)䧒���o����aXw�ߝÌ+
°�{��V�a{��[�V�a�N��-���i�n��aXV�}���8°�+���q�aXV�ﵸq�aXV��z�aXV�_>�t�L�t��عm��l�U�"��B���Z�b0�["WG[-�=�\��i�i�8°�+���q�aXV�ﵸq�aXV��z�?�B?�c
°����naXV�����2��[��զfi�8°�+�w��8�� ��K�R`�`��`ad��FX��ie�I76Ì+���8°�+��p�8°�+�]��8°�+����N��ְ�humֵ�q�aXV���naXV�}�p�8°�+�]��8°�+�w��8°�+c�tfѢ�5��V��1������8°�+{^���V�a{��[�V�a�=�f���aXx�x����V�p���Ì+
°�u�]Ì+
§�3=���n�V�a�f���aXw��Ì+
°�oc����<7�}��u�{�.H�/JO.R0����.R���(��e���naXV���naXV��k޻�V�a�{�70�+
ù��70�+
��>�n�k*��Ѭ��naXV��{~w0�+
þ�naXV�s��naXV�s��naXV��5�<��ֱi�U�4�aXV�}�p�8°�+���naY�M�I� �l6ù�s70�+
ÿ{~w0�+
���9�R��C�nh�8°�+���naXV�}���aXV���~w0�+
þ��naXV���y�����5[�'��O%<��w羻�V�O� 3����~aXV�����p�
°�>��q�aXV�����\���ZfU1n7���q��8�1�d:�*��"�+3s
�.0�(�*�\-֯!��aXV����Ì+
°���V�a�}�;�V�a�k���V�a���y�:�u�]f�Ì+
°���V�a�}�;�V�a�k���V�a�u�]Ì+
°���|����c��f�h�8°�+����8°�+�]��8°�+���naXV�}�p�8°�+
~��8��GZ.���aXV�}�z�aXV���{70�+
þ��naXTO����H6�aHєV�iZ&AdX*�FLd(�
Q�(� �I�0������V�a�>���ӭeV�M�j�aXV�����q�aXV���p�
°�>��q�aXV�{ٸq�aXV�$�����?��5��Yk��[u�n�U�ຩ�;V�(B:E[��Yu
�<ݜ�f���[u�C�
°�=����p�
°�>��q�aXV�{ٸq�aXV{�����aX_}�=�[����u�3F���aXw������aXw=�f���aX}�{��V�a�{�70I- �����V���s5��o��� ���{�m �����q�aXVg}��8�O%<��_~;>5��[��'��aX}�{��V�a�{�70�+
��｛�V�a�k޻�V�a������5WF:4:ַ0�+
þ��naXV���{70�+
þ׽w0�+
�����8°�+4@;�������;���A��t��<�@]<u����9S���+n�ڼ��@c'oc�h�&p1�L HظX�e�x+6��h.�n�yv<��d1��}b��x��:��D�(�b�a�Opd1u�5�����8��s&��4TAYa� �4kZ�-���ej��a�Λ&�i==x3�m�:���۶;M�z�Z5����Mt��w%�ؒ�1�s��d��U�u�1l�`v����,#�WJ�S�,pt:��S+���?C��aX~��ٸq�aXV���q�aXV{��q�aXV���p�
°�/���L3�G4�k5��V�a�k޻�V�a�}�;�V�a�{�70�+
��｛�V�a���[�WV�Қ.�k70�+
���~w0�+
þ��naXV���{70�+
ù�{70�+
ÿ=۞���Z.:ҭ��p�
¿Ѐc~70�+
ù����8°�+���8°�+����8°�+ｗ�L�1�.�4�h�8°�+�}��8°�+���8°�+���naXV�}�p�8°�)��ﳥ��v�t-�`�*N"���Y�6��z�Of�Rl�s���m�f�h浛�V�a�����V�a�w��Ì+
°���V�a�w��Ì+
°�y�Z֮�u�m��5��V�a�w��É��I?�M��
þ������aXw>��p�
°�;���p�
°�<w�o3K�к0�Z�Ì+
°���V�a�w��Ì+?���{?���p�
°�;����Ì+
°�����p���j�Ì+
°�;�f���aXw=�f���aX}���p�
°�;�{����aX_ϯ�0�3EӪ9��naXV�s��naXV���{70�+
þ��naXV���{70�+
���_����]�f	)XmF���U.���GS�9-F{�sX�V�㩀{>�e�NՍ�&����C�
°�;���ٸq�aXV���p�
°�;���p�
°�;���p�
°�;�ݹ�m��M�Z˚�Ì+
°���V�a�｛�V�a�����V�a�{��Ì+
°���|d�bfit:ә�p�
°�;���p�
°�;���p�
�=�@E����� $eB�0B�$8B�!��8�ٮ~�Ì+
°����䧒�Jy?��Ko>ƆAr����
¿��0�����p�
°�;����Ì+
°���V�a�w��Ì+
°�y�Z֮jꚮ�KsWp�
°�>��ٸq�aXV���p�
°�>��ٸq�aXV���q�aXV}���k۫�֩v|�ZN���Z�-�vL������q�ڲ�i���<ņL2��A��w<��%<��S��{�70�+
��｛�V�a�k޻�V�a�{��Ì+
°�����p���j�F���aXw;�f���$��°��������aXw?���p�
°�;�{����������M�j��ե�f�p�
°�=����q�aXVg���8°�+���q�aXV��ٸq�aXV�����WZj�)���]Ì+
°�=�f���aXw��Ì+
°�w��Ì+
�$�7 R����� �(������q�}��]Ì+
°�϶籴�Z�N�#�5��V�a�{�70�+
ù�{70�+
þ׽w0�+
������V�a＞39�ff�^�;pgv�Z0ln;S��X�p�4��\;'R894Pݒ`�ϋ�n.Me��w�{�
°�w��Ì+
°��]Ì+
°�=�f���aXw��Ì+
°�㥷~�4��kV�kY�q�aXV���q�aXVg���8°�+���q�aXV��ٸq�<��S�}�����u�!sy��y+
°�=�f���aXw��Ì+
°�{��Ì+
°��]Ì+
°���ј].�Y�q�aXV���p�
°�;���p�
°�;�{�p�
°�;���p�
°�<y=��ֳL.f��naXV�s��naXV�}�z�aXV�s��naXV�}�p�8°�+���{�����xu7����Zy�g67�����B%e��(݅���T�P��&��3z���!��r"I4��4C��q�0na��[~��F������1X�#���d@E�R:kZ
`��E�@5wI���a���`�i�L jN�.������Xdn��-96� �0"�+�$�~?\���j0Ƹ�PY���7.�٨�(��h0�? �$��F2*	#hH�'����,#��H��hНܳc "H�JZ1 Ґ����a�
�X��c!��A�DE����±DD@bH��ł0ZR�1��-�AQ��$H��DF(+���`��SZA�
�0`������>�?
�p�d3aa4j�&�0͹�ֈ&��QC
QTpjQ��[!K`�&��C[JHbb1���Df	؉���9'қ�4HL�c1!jq����cX�����A�DE����ɪ,g�
%�0C�PI9 c�"ȑ#A��0�"�ѥ\!�@�`��q��`���ɂj�@�d�V�D��e,� ȱem#���F0b"� \��",�a���33�UU*��UPU�KY�e��m��h�%�)LF�]�vl�Umv9�îua8n�w@ơݞ�Ѫ[,���6�0y'�\cDs����f�L���c�p.Rf�a��g��
�����`����݋���� '�J�-܌��$u�� ��v�ٗǑ�;<�{+ړ�'m�Wl8=�u7�M	l�7nP}F� �Η<�v�6
��^9���bv���V,�f�-�v�.H 9�������j��P��vI�×��u��g�UK� m"����ѷ8.��Y�;�N��;;��(.��6�ˋ�kggv��6M#ö��;%�ua��qs��6='`��7e갷�=9N1HOa9T�6�-�W&�w��9�-����nç�����v��u�([ 㰻�t۷a��.a1��\q�Vj�#Nq`�[�Zg�6m�hMO[�*�3ric�1�E�[aF�e��2��R-���Ǎ؍[͹�c���E-y��3t���l�����\�5Ss�z��\q�n�����[f]�K�-��r�B�{a!T(���*�8�;��v�r�\T8�֜4�,��-�L��Ѯ��j�遜cWZ��3%�;hဣ0䈏vV�%�y�i$;�Ih9Q����p�b�25�u�hE�FCP�:�q�K�ڀ����x�`g����#���Zzl�x�N����ήװ��1��3ɉ��o����[42�ًh�X�.�!����z�\��u+(·�sD�5Z^88UvPU����ű�Q��7�=m�C��'a���j�h��=��9�3(��ݓ%�᪘;ynPqa�^�n2�n]V��qU�T��K��"�����H��[�PvL�˦xy�l
q�Y�Ͳ��n
)��	��,�����lj�֛]��mnJ��'����嵶(�]Of籱B@�q,��Ն��֕�!�k�Y�G�V���.��ӻ����Zy�q\+"\�ӝ�܀z����'HN�!<B}	a8@I#$	d��8H��$���~�a�}�<s>�3WX]]J-i��W2ԛb	�MtVe0L����,6V4�_(L)ͭ���c�X1�l�g ڦs�@
��䡫t9�Zwn��S�ܼ�nКX��Y��s!Z��`�]�笹��\��vT���``�d�"���;���m�%K��5��:7��ݍv�i��F�V4�l��T<�4�2�ڎ:٢����kgV#y���1��x1w~��ww^�u{}�?[\��юWj�����g�y������;Z�ZK�U 5��.����ۗ5���
°�=�o����aXw=�f���aX}�{����aXV��f���aX}�}���WF��U4-֝Ì+
°�{��Ì+
°�}��V�a��}��V�a���;�V�a��s��7Z˧Z˚�Ì+
°�}�;�V�a�����V�a���;�V�a�����V�a~���o+6V�lܧ<��%<��S���~�Ì+
°��ߝÌ+
°�{��Ì+
°�}�;�V�a�}���w<��%<��S���s����aS�@g�����?0�+
�����q�aXV�wٸq�aXW����=�����n���@-T�Z�z��4��m;v��x�d�pC�ۉ�k�h��Zt:��C�
°�=����Ì+
°�}�;�V�a��}��	�aXV����Ì+
°�?����:.�L���u��Ì+
°��ߝÉ�BO�p$��a�����naXV�����aXV�s��naXV�N���x��������w0�+
ù��70�+
���~w0�+
ù��70�+
���~w0�+
����&auGN��sY��8°�+����8°�+���n8����{�{Հ|�IM��նݱZ�0���옰����p���ו�v���MJLg��6��\�k�ne�C��/&�pf�d���m�3�b�۫UU���ײV���K���V n¼��Ӫ�*�n�`䕀}%� ײV���Q6�*�V
�`����Ӏ{}�w��O " ��g�BM����W���6������W�+,�ܜ��y����n$�,�l��$�)qQl�|��M�����6V�V����OggNbd�L���ۊS� ͝=��&�[1[s7��/E)�c���:��8U�ӫ��X\�XҤx��X옰RZRb�e�Iӫ���y丹�6G��`{ذ������ۺ�h�+Cwf��V���=���ק ��z���*�r�;�wvb�:���>�p��K�!r�Jw����]�Z� I#7��K��V�ԏ ��+ ��ŀjd5�t1��^hv+Ӧ�N-bT孖���1��k�m��H� ܦm��v�m�{%`}����X_d� ��:���Z��*����:�%`ݘ��ɸ��{�g��ف�1���ݘ���X�._vV�!H�EӪ/����Z�>}���\0��w�%��}�p��>��Ȧ�l�ݗ��+ �ɋ ��J�>�7�����r�Oj�uä�nl��g�_}�:��� ��át��u:�#��66m��ƫ�ݷn�!Gn�Ý�<�:��q㞑�-'6��Q���l�Ŋ.1�y�o��h���t;�<�m`�6��)[:�u�7��ݘ�6@�����F��#���T;�M=�wX
���lA���t��.A,K�ƶ�7k��g\(��f2�g|���r�ҏ�wm�=��&��=r9՝�|,��n"�̀б�fl(H�A����E�J��|I}�x��d��.�M�����:Wª�옰�d��._vV~�-���A�ܛi�vg ������IX_vV n�xb����]��wv4:��:䕀u�e`엀|�%`a�[�n��vZU:��:�%`엀u�J�:䕀ys���//{���g�s�g���\d�[�f��<���[=\��h�Tc0G$�30K0�l�Z�����se`rJ�5�J�;�4�٫���4�Zڿ�~�m0a1a?� F2A`F~$r�9;X���I/ 'Y)N;�B�.�N����J�:�%`�/ �앀G%WE�n�*�� �앀d��IX{%`�ʔ67Wt�_
���	�^�$�=��~���=���&��4�aR�]�c���U�r��3�׸��Y���Yc�L�=����UUWwx�IX{%`�e`���ݝ�����2�.���N�vV M�����CT��黲Ш[�5���업+�����<��I�� d������>.n����>�SQqP+��Zn����x�IX۷^��
(�[��_-U�uw�|䕀}%� ײV n���(K.�s����n�ӊ v��+qb,�3 �
h��حl�4�G[T�[��M.�����k�+ 7v^�$� ��aI����t+VUـkݕ�M���$������7����ܦ��w ���0�����`�e`d�)�D�<nEĖ��Ė�*�K�{_��?~���wW[r�x�i���X�\0{��ݸ`9%`I89��v��޻P����m}���ti�e�q�t.e�*mQ��[C)aug�G'� �ۆ�W举a�z�`O��Q���e���}zp�IX�\0{���B3�n�ЭUջ��|䕀}%� ׻+ �ٓ�ݾ�݊�#Wp��Ӏkݕ�n�ŀ|䕀u�;)�6�Qj˻x��X��X�IXһ��=��ݻ��Mjk���vȸq��Dŋ�]E��KR==-�\Fօ�q�@�U�g����w4Iv4heR�����n)�Q��m+n�Tf:��=`Y2��빰᭜�+bZ��E���9��p� �{uѝK*��A�b�m.��g/M�ʳ纷���1z݊���{ҝ�����[OV:\g7G8�l�xQ۟$��a��2�J�i�I]3�'�O$��ո~�%�!����[���غ�}9y��z���r��7�����kT�������,�$��R?�����o~�p߾����3�ɳ8��{XҤx���ݘ����U;���Wu�}*G�k�+ �ً �V v������eU�^�X��X\���H���,���T�:�i���7vb�:䕀}*G�{}�w ���%ܾ*�|+6���xz(V������3���jL��aV�������:䕀}*G�k�+w���$�]:PnB&�2<L��%����BB2� ����?HB�a��ՀI.\���e�1�����`�J�7v�u�+ $�xz*�R���ۺW��]`yq$��0~�� $�x���vS�T�K�)�;��o ����d�M�`\I>��߭� n��\�
*����7��)OFe��˦�9{T�D������V��ڮe�[���}�o���	%� �� v����5WChuu�G�+ �\0	ڑ��+ �5e��;j�uu�I&,v�xZ�ϸ-�ݤ:\MjC�n�C"���$��M�XS��7	M
#����pȑ��&̆��i�22&��m�fJ�tY� �(��O�#iJ��s)�5�Q�f� 0a!�B�c3�30EU��b��"B,�DPF",ENi�e0`�+2����%A��bh�Gp4E`�Dc���Y�),�B��9����L�P�AT��5K5�1@P@ѥ�jC�U�R0c�
(������t 0!5 �4B��d6IЀ��B�M���q���rLre`���$B�U;��i�[�X�H�I/ �vV$��{)�V]�+v�h���Ix{��	$ŀNԏ ��n��Cv��eݠ�պ�:������A"�(���k�Є�9m]J�imf���v���$����\���{׀n���P�n�:��I1g���������x��X����c�.�:����V I%��e`I� �`9���SwwcE]� I%��em^��ٵ�?+B2*,�jH�D��0�	$���@�!�I�;�����ϮWK� ���5���<��z{��~�� $���P7�t�E��>=5���]JV].v S&��lkƲ�jȚ�^���=��qu��|��b�>rJ�	$�^�DB3*�_�ZuWuk ��+?$�l=�z� �OV��{���犢��t[�[)�� {��^�d�<�9�$߷�ŀo��x޹)���cwʵC���5앀Nɋ � l�� �EZ�Pڻ�UwhUu�Nɋ �R< �%^�X����k�S`������$�a$؆�ݧ���43p٫��lQ��v����J�BLQ.�`��6�5�<��`h�P�\җ`��lf�Vq!���\rZSֵV�>_\vc��5Zg������9"IӃdi(,��1s�aFf&��5�9��&t�Љ5���F��Z���֌�7Vݹ��&��5����]6"�k��0��אʆ,�(7{����w������.��n�W��kOޞ���v����V��籩9�̥5vڳ$crgK�s=�o�prK�^�vLX[�m���wv5N���x���	�1`׽���OgnWK3GaUx�d�vLX\��rK�CS�)7F�n��E����I!/���m_���mse��vV�B�0*��*V�]�Z�>rJ�5͗x��X��X��vn�Y�,KiIUX\�]P�N#8��G[UV|]KWAus��-�[6g����)���l��5���'vb�8�Ϙw��< �}��e�m�i�ʪ��^쬉qo8����qs��3~���#�5͖���{7qlU�+ �w �����J���˼^� ��"�嫺�WiՎ�`ys������V���^��4�se+��]����9%��d��.\�����]��r���#�B�=<]��lPKlp��@�s���]�B�F\MƐaV� ײV���IXrK�C���Ѭ[���nk6�;�uߤ��ӯ��`~���{��˜��;�C�����F]�N�~���;{ޯ�>�b��1QE�A(#�" �0�# �DA�'ĀO��)	!�z�_�j���j=��U��U�����������>�b����;�����۵E��� ׻+ �I� ��V�N$���p8�������Go=�p��/5(,v����x3Aa�\�n^�Uݠ]���d�9%���$���)?F��s�s8��־z-}}�k[W׽�m^w�ٿ��^� �F�$|Ix��'T�e`Ip�#앀��U�T�ݔ�huwx�O�'� ��X}��u[$���@K-���)2D�d��}�y�kj�����ѣ���]`M���%`͗x{��ӽ���d�0��JK���`d�^�wG�M�m�r�oR��WGj炃���j���;��� ��V�w�G�V�ۆ$���u���d�&�'T��q%�X�n6K������m��2�UWw�G�V�ۆ�l�{� ��ߗ�~����Z�X̰���\0�K�#�]�y$����V }�w�_*\ˑ[��޼�$�{=�k\W׾�m^w��}�� @�	�y���]nf���)��5��\a�m��n.�`�V}�
����4�j���Q������u�qK���Q�8 z�3oR������]%�Kl�$_�ܒ�>�W�f6iJ�1�!f	Tۤ�V�'-s�X-�n^�k��%�� ;�ȅ�F!) ��d�7��S���1�͛3,hv�����;f�o'+Щښ`��]C5[�	��G�d��p�o��\L���a�T`]dZM�m�N�d�]�C)#���]%jFў��]�C�z�����#�+ �K���/<�C�߾� �}�~YI�Tl\� �d��\�g}��y�z��x�S�)7j�Nӵi���>��G�V�� �d��DX���ӥl��V��J�#�.��J�>��~�/�Y�m�31U���W�G�V�� �%�4.ʕueZ5���Lv��#\�8�:2��
�뼌ڛ `�����X����l� ����� ���˼��.��Wv��Wª����3���\�qqr�.O� $�� ײV{��\�a�yU�軱էV;� 7����*�{%`M����)�VSwTXU���*�{%`M��=�s�o}�^ uz7��Un��������J�>�1`d��l��=ė��������C��r�ggV�pؕ��^�Ju���\�H�&'�:�f(�ʎՖVV2�߀���rp��^ I%^��G#�>�Z"�U]��WE��Z�ݫ �ݫ�5앀}$��?^���YMX銯 ;��<���6��dd�HDa$ ��\Ĺk�*��}0I/ :wccWV��1�Wux{%`Ip�	����y$���x����r��𪫬��%���_���^����ӽ�a�cCKfά�4y�1���{sK�����qӴ�֮����bL�::Wn�Zwc�0l��l��#�+m쫉+򵏐#�ӌ�L�q$���#�+ �lŀd���M�W�~t�st�� ��� ��{��	�^ I�� �k"0��i�iڴ��`M��l��l���\�$���7�g��W���c��V�kf��`�/ $�W�G�V�ً �to[��bJ顳n�(hVWGfb�ݶ7���t�ѡ.d��h:-�	8�uJ�wx&ʼ=����^I$�`z{׀l�m�V��1�Uux{%`M�`�/ �Iw�w�H]Sj�c�\���zp��� ;��8{%`�NU���h���v`앀G$��#�+ �K�do.�kd	V�c�J���%�λW���6�"N�ǔ�h"������Sp&��D��X����	��m��Hl݉hȂ�E�vXVA�EH�Q��{f#6;��7�؎k�#�����i�߾?�jnR�!B[\��)�k�{��M61f��6���o��8�Jg#�|�q��U�*��.�R������.w�0��4r ���P(P���R�$F�`�DQ`����MlWEN
"oz�5"�1"F
��E�ю2���nI7�@Lf��%%J��
�&�b`��3�)rC, D��#�F0c"��mB������d1F �ALQ9�e`Qw?�4��IJ64ԓ� "E%�c�VTj���"*��{є�D�kq#9�]C$P�B/[��@c�0`�ZDA�@P�	PaA���I5�#w8$A&��c"6Ĳh!��1������R�9���m�UUv�YmU����� 깔���ѻv;�bS��%ۣqë��9�ф�1����
�W��R^{M��a��nB����gl��N.0v6�v^j��㳹I@:"�8�RU(E��y��L��.��(=l�=˃���gm�e�X�9��x��u��S��`��u�^�Z�d��ុR����֜b�Gm��S��Ui6)8آ���gM�'	G8�w��sXȷ/#����o/f{SŜ��v1��4s2&��!���Bm*&��Ck��Tn0xP6�l �t������Ү֋y�X��2h�q��v�� B�lխ����c�\��pEF�%p7{ �F�7�pR���]�۵F;n��&+;rн/]�1�Z�(��tm�󓮶��6�v9��q�m� q8���E��aKt5�l��,���k�L���XJ�WK��F���ob��dN���+�j��g9�1*Z�����s���{(f����L�q{;����/[�-.}�	�8�^�!`��`۷�����b������J�b̘�T��i�ڳ[TC\	�kt��H�K�-�b&�HS�����mcF�:m��#�ڣ:4ܖx���q"e�v�L����J#ui�h�&�e���v��J�ls �6����t��)Ů�h\ڽ����ۘ�d: ��S���onW��E��n>���.v˗��n#!�NH�Wku���7�{85�`���]��k�(XR���n�km�W����u飵!��Tp�[�B�I�wTn{oMe�5Ԧ�9�.�B$؃ahF1���bB��Cl�M�B��2���$*��q<+�a|��'7=��f�`��\J�ά�/��K�\�Cn�3q���	q=,Q���9�W�ul��a��ضn�e�1?K~^`PEک�e�2�z�f�8��'p�:��<���Y�j�A��g�"���y�꬇c��i�8��;�s�0�;7�f-��mZ�8����.��5v�Um�O'�<���'�y9!	�t�@h�BI� �$�	G�H}��s.�Z��4�Jl���y����^5�h0�{D�Lv�q�ۧ$x9�l�%{lv��K�d�����y�z�7=��<:��7�yv��R�gq�c.:\�W������i�a�>i��W���Z�W�˒��g�"I�O5��݁x�턶]�{d���s���*֟4�%�`���ͬ5.n5��kd38уsmh�8{'��u�ų�b����][���}������C�P9��e��b&|_�圼��<L�%#X��nu��v[��Н;�(ی����]����� �����G�V%Iu�l5�uUvR-Zn�����J�6T�X{%g�O-?��_��L�,�Ý����� �RU`앀}$ŀ|��C����N�ҡ��%Iu�G�V;&, �%�N��eհC�i�����X옰l��l��X�V���4���ڞZJ���<Y��N���K�JB�F���c��R�\W*�t|+��;�� M����� �d� ���X�ms]���޼'HI<<�y �d!�'��koy��j�������{�ϧ�yi����k�I�Z��;�O]`앀N�ŀG�V |����N�v�Zn�� �d�wf,=��=ĸ����]`�~a�:�V��j�wu�N�ŀG�V����#�+ �������l��º�B�]�\�L�V͌mD��Ye��"�M�G��\u�;���Z�#�+ �R]`��Ē��}�b�:�8���b�j��� ����qs��I��{Հw��, �%縔�==���9����]�>����y��f��������`���Y	!��{}�s[W�Ͻ��~s�H�8��y?"8���o3�%{l�J�l|IS��$��(�1���8�3 &�x�%��X�\0�j�'`[C��g ]Z�6���:3���ڜ:m�jl�5���i׵��]�#d��J�� �vV�� �����P�$H$��*w��%��`엀IR]`q�,��V��j�uu�}%� 'd�9%���gl�L�.�b�N���� l����\�.+\⿤�0�
��F2?̑�$�m'T�k�Km�q%O�|Ii�H�pk$�3Ļ��ku]����]���ֈ�A�GO���xzkm����2�� ������zp�%`�U��R�v��J�U�����9Ĺ��=�� =�z� �{_V�y��1<D��*}k�I*��~rz���� �T�]�@�a#�I[k�IS���-�U�;����@�cn��Vd�\��e`Ip�#앀IW�N..v�hm���ҥ�V�.��4�M��6^\:-�y�4��.dI����c--ڹ�k<����<u��m2Fwj=c��t'nB..�ٽ�75{u��k�� ޥu�u���m͟[mA��;>c�<�q�O�CN6m�rT�ac�"K��m���]�����|U-�j
lە�]q��tN�>��^�A+�⫀\�����Lc(��1�Ѣ�F�2����!4@�v;���r=5�m�������mt��WSݘ�|&��y�<[/k�umy�����炮�	�_� ��V I%^��;a�sCM+���ן�y$����� �Հ}%�<�I�_�
~0X�(4I8�W��8��{_[l� N�xӻ�,`���:�w�G�+ �K� N�x�Iq7=�;�=��|\ٶ��Wp��Ӏ���d���J�$�L��*�_N7g΅��/R��^{�a��]�u�e��H��srk��xA�nb0q.$��%�#�=����`�����*��7wX�Gyk���%ʢ=�Xf�8o����w��WA��V�=����a��q�9�V OO;�6�,����Z-Rn���0�J���앀}�@�.�UAj����=��.q9��_�y���6K� �����@f�4�)��
�.�a�q����:�Wjg���]���1fx��N�wJꮰb�x{���p�����Հo�����V��һ�=�X�p�#앀��w�H@��,�W�����G�+
K��25@`# �#)�S�]�K�#ݕ�M��[m:�CWV�ـG�+ 6)/ �vV��8��� ���k�:è��w =��\=�X�p�#앀w�h�A�[�ݙ���z`�wS<;<ɜ�[���\�H�\uP����T�������G�+˟0'����b�˧T���j�uu�lۆyqs�M�{�V {ǽx{���4@x��N�t]�]�}��BK�#ݕ�l��������L�����5�_I$%���kj���ͫ�{��^�PH�~&�@�w��6���{F��慺�.� �d�d�`앀/�{���NӍ�e�Fke��W�]���g�(<3q��nnx�c�*�H�v�81Y�`����6m� �d� ����M�;�[٢�ҩl�*����pBK�#�+ �.�ě=��O-][�E�Swu���� �d��\0�J�	�+l*�n��񻺼=����`앁�9���z� �;I�m���4�w �޽8o���	$��#�+ �s�.q ��$�C��-�&cy���j:�6��k)h۫�W	O�i$\��&���͋K
�2�:�Ʋ�u��p�=�n��v,P�.,n�B�QHC!a�cѹ��N�n��D�θf[���q7�[Yu�U���+W�x҃2�$��W���7I�MM�H����Nw.�v%ݪ�B^%2��Y3֣���t�ذ�Ÿ�Z,:��ay��-��hf:�[l�Wk���y?��>?��ؕ�mF�JmF�]�Ģ���ڈ[���C�B���Ψ��ع�õ��٠y�J�	$��#ݕ�}%� �[-��MawJꮰI*��e`Ip�#앀;#CV��cuUwW�G�+ �K�d� �J�n���N�Їwu�}%� 'd� ٱ��n۔��;��wc�0vK������'v�Y}��حٔt�c�_�����e�>qt�ut�6��s;����IVD�Qm;��HU�����7�j�7���	���V�|[�=�Y�9�> ��!$`��s]v������;�6�0�uAj�+T���v\0vK�	$w�G�+ �(��x��MR�Wwwf N�x$���e`��u����������� 6IW�G�+ �� ����}ݕ�]��<�؀��V\;��a�r��Hs��v�Wn��Lpu�^#E�G�+ �K� N�x�c�
2�Ir�]�?wק ;�z�f�xse`vܤ]��ݖӻـl� ٱ��q4C����Ő�3Q$��D�1e���lx#���z��Yv�ђ~61�3fk��X��:��" 1��"����9��+Z��<�o8>;�|c��ϾUs�����	��.��CJs�h��h����#xjDDB,EA�� p�nkA���rN���0� �8�-�*P��T�|D~�;$�u����eF%� ar"Lu A��&��F*1��%0��O�u���HĈ�D���la;T�d�,�b%�cܘ��XP�C�7i�#�K�@��a��e�J�S{$PIa���O�l�v������h���[H��b��""4��A-�I�h ,QE�z��?~���	��Xd���~��ႰDXk�
|�1��)̙���0��];��޹-�~͜䆒/�L� wB
���CBAA�t$M()�,J�)�
��5Ʊ�O��@!�&�4��$��RI�@��}&�h��4|
�	 �HBt�I2��\�qZ�\�Ė�\�n�0	���7���q�Ē��'T���'v��.%������=�c����_V� �l�wn&��	6W�~�ӱ���SmV�yYv�e�i(��q� ]h�����	.n�鳣uiIڥj�uu�N�� $�x&�~Iy?P��߷ ����o#�Y�2�� �e���͕�N�� �[х4\�/ ;�{^��{���0M��������V�UUV� �l�� �e�Z\�s��9@�$� |BH�}��m^~3�R�v'WhC���>�p�	6^ l�� �l���\�p��&��We�M�b�8nȴ'=r��2��cq����$m�vss�ay��1�vseR�����{�k�#�+ˉ/�w��`��O.�ҲꕰUuw�l��qs��g��� ����޼ ��;ؔ���!-�x\�X�n&��	6U�SBVU�M�jզ�� �m� $�x&�<���p݇��^a�h�UN I��M�����>�p�)s�O=�N���q�f����� ���\��+�ź�2��(�ǇH��0����y�uf�9�\��h�7N s�Nu���[��+�|��N������������ۧ��pD���Ӊ{	�� �$mۓP���Mj�sDtu��$*�i�6��%h]�R�ten�-�KT!�m�<X��y퀶�J ��-3n^���v���I�C[k�u�܉:���~�������kz8m�I�8 px�áh����0u�x��]�A��Å��T�c��ae�YUw�	���e`�p�	�/ {���T+�T�U��M�`엀-���8���U�v��UX!��`��&��	������~�_t�Geli� $�x"�����$�i%<�w�t�U�� H��9��	%� $�xOy�e؛*��wMU4X{<\f����{2A��:����e٫(e��ӌ�Hܭ!f_�}~�ۀw��8&��	��:���n�ն�V[�ͫ�����~�~�H��I�$;!!�/5��j���u�{{�sj�F���,T��j���� ���E���e`m� �Z�6ՅS�UՕWx"�x{��	6��^ .�A��]�ӫS�wx{��	%� 'd� �Ix丗95_��Jι�B���-uAk����c�ř랙3q��,�@��̪�&ـUw�=�_� �e��K�#�+ ��ڝ��쭃�T�{�^ w��xKk�J�*�KnZ�H���F�q��^���ڽ��sn�H04B�I ��B�$�9�s^v�߽�mW�)���ꬶU�U���	6�Ix��xT�q�m�v�5j�wu�lۆ�.q?Oz� ����#���?�콡�K5v�).Kc�e��L��-uh�V!�m.�]�N��]j�b��A��r��j���� �%��e�앀I���T�N�WVU]��e�앀I� �%�N���Jګ
)ҫ�=��	6�d� �l�r�B�eUZ�]`m� &�x"�xM$!!!.p� ��E��1�� �ȣL�����{��j��av�����廳 $��E��䕀I�˜}�תꓥuJ떙a�+m�6��ZK���6���`�;6-W%U��Gj��"������ӿ<����$ۇ��>`{���`��V貙V�5Wxse`6�l� ؾ����Ǻ[�wZ�F4[�ͩ=/� I��b�xse`��y��Y�*� �}��{=��:���6m� �Q�L�媧l��*��Ce�앀lۆ M���I�$����	��۹�+SU����)�JΫ��%p��mc�
�i�cA�l�� Z\�#��k���m��cua�9p�c�Vk�E*n��;�����ی��G<�/!3V��3�*�y�s�X0�k6h�{<�l�hZ���DD@�ۈ�8��;>'��L���Mќh#����m�[���t��!S��M�-khc��x���U�NduS�G+�rΰ�B} �	Cz�4�5�k�Z�P��&/k�Ёl�ӭ�'&����e3N����p��X�Y�4f6گ�}}���w�^�$��5��>�QN]�N����&�� $��M%��+ ����Mڲ���/��� �K�	4��*[__^ʸ�ۖ��$�$���� ٤�9%`�p�	$� ���^��� �!p������n$��6;�'uAc���U2�&���]SF�2�����űQ���Շ%�<E�eB�.�݆[tc4c-]���pI/ 6lw�G$�荍��mP��kZӵ^����VF,X�v�@H�B�a �$֗��w�u�+ �m� ��֧�l��WVU]�͎��J�'v�G�V t�Pl*Ҷ�uV� �d�wn{%`��uTS�ն��@UU�;�=��fʼ=�w ﾉ��mp��2���� ���ۭϞ���b���N��u��Sd�b���z��6��uv`앀lw�G�V����;�w��
���SW;��ӯ �IXݸ`�+ >�X�ӴU+�BxrJ�;6�s�qsx��˸�e`�����ct�Z�j�uu�vm� �l� ٤�9��ŮYVա�V�����#�+ $�^�Xݸ`����Io'�Zk���ێ'�R���I�3,g��L��t���g��C)sY���ķ3��� }�O^�n�0�%`N�ª�j�,�T]����&�� ��V I���*)ˢ�m;��Wu�Mۆd� �Ix{���OiDݫ.��[�ـG�+ $�^�sk���l���-��f9e��p2И2X���bƀ!<�Nw��N��w��
��e�����K�#�+ ��9����¿��8Y�0���!:l.��V�	M����:�V�7����)գ�Gv�K�9%`v�G$�%�z?^�|ߌcwE�h�i���&��<��<��V OG��#�Vص�k*ڶ�J쫺�0䕀5��#�VٯN�����,��,vw�'����x����;6�G�Vֻ�C�HUaeUS��#�+ �.$���ｚU����m_���O� I$�� $�� $�� $�� $�� I?� I$���BI�� $��@`���@@a$�	 "@P�0��@D$��I"@da$	 (I�II$�	����O�B I?� $��@I" �I� �I�� 	$�� �I�� 	$�� �I�! 	$�� I$� I$���d�Mg�H���~�Ad����v@������H �      6V :@H	���J0 &��-P�CB�i�i�T�6�J��R��Pd�� �`�hd�� Q��	 �	΀@J&�h�j�� �	�"f��z�*(��0&�a4�49�M0	�� L  )��U&�5!�� �  `Ld0 �  I�@�$�& 	�LM0���V��e�  )ϬJ�  ��)�� �3�����p�X�I�$�JCdChC�S ��%��L2�eȪ�P{6X�:��!Wq7˪st2�w$�/"-���%A�4U`��hPU%�ՙ��Yg�*2�!B(�(�R�QVaU�e����{���J
�ieJ�+s{���SMf��k"UkZk��%��0�ʼ��m���)�#dJ`U�`��%��2 ��Ē��L��Vh�h%55(� ���R�U.��]���I0�hK�@�ouxUP1��5p�w�P0�j��*��$r0�2�����\�Z�B�D@
�K/�^@���IWx�K�aq�$D�Xي��i`���W�$�*	@�	LR�&�ֈ�	R,"T�1������q�'���%����P��߾��w��                             ?\=                                                                             �@                                                                            �=               -cK�6i�.'���]��/�[oz����"in�@X�v�^:��ם�m5�5�۬\K$a�x���9l�n�3iR�v��sm%�V��H�.����޺��`�ͭ��$v��n��hְ[M�l�Ktͱ�8ۦm�@��_Wצ�m�b��m/i�B��lm�L+i5����-�]�]�$�mF�,t���p$�dk��km�,l���hv���]t�sm��m �[.6�5�st�5����Ė��:t�%�]wM�l�䁺MZ��)�K�\[�$6��6C2���6��[���Ku�5��v7En�D�����M,�ni:ČImr�,�%�qmm�i<����z�I9�U�-����lݣ�Λve^^f]]�g�B �e܁ �R�p�a�@�� 7�@�@���X f�D�@�U/آ�2FvBd�5
����D�	W&!��TII�[E2�£<������߃��    ��              l              ��  ѵ*���;I�v�Z�k2cH��o���V�[.�nk�K�]�\��f��U�fm�sI�kn�/Kk�4U�Zi���N�ӵ�]�^XZ�YO�s��\��6��   m�  m������+^�%�5��P����ubI%K*Ҽ�_�w_�T�ߥ�־����I#o��7r{р Z�HF	cyy銪��f_��=u$���&�o.x� Q�Ċ��{ѷ�雩t��罈�Ξ  �XRb���[�ʮS_}���Ͼ�ڽ���s�4 ���Y������/$�e���믽6�s}         ӛ�m&t��:KzƚI�� VQ���[y$6�s��m�zf�uI���*��c  .�,Xb����箧���I6[y$6�ryH wH(�y�������7r���e���_��  �T1n�e��Cj�=�F�y�/L���@ ��YbX�^I���{箧���I6[yڬ�M           N���OSz�`ӭ��k[U qx]�.�I>m�zf�uI��y�b3q�  Uଠ��ݩ��I6[y$ݻ���u�   f�7s�Lݮ��j�0!Z xA)h�g߿����{��+������u'���g�  �P]���I7n�=�F�W�n��O��{=4 �10Źw���^�I6[y$6�s��  �         m�X�֫%����2��$� ��W�]�f�uzf�^w،����}� *�V�{�}��m�ڽ�{ѷ�&n���U}'�  ����,�ܯ_��>2�[4���;�fӌǵ�4�al���O]�y��u���H��ξu�z�����q�N$�z�i4������~�� i3]�alĶw�kٙ���Ve�b��3i���,��Gl1�}�>tq�i�՚*�%����8�a�^�33     �A� ulH����{Y�Zk/GI��1�y�;���������ү�L-����|�3i���o�u��W�<� X]�1 ���+�Ğ�f�
��[;��3�ė�U��]ӾPr�����;���@ �(���fSf�J1��}���N'X?}�Y��XBY��o�G�ڇR�������:�Y�t_>��  ]�
�{��Hu�q:�H�=�\ۢGl1���{�È~@�%u�J��I����&�Hj�~;��R���w+�\��� h�\��A�6�f�"c>����נ:�nB ?}Z�P��!$v��{�a��;S���P!A��s��*ʽ?��>�f                               �=       4����z_J��䫴J�ͭ�v��y��W,�<�m`ӭ,j��Y�ѳ�IzJ�܏,��R�ۉ����I/Z�:�*��W�;����G��`       �k���ݴ���ɳI5��x���n��	Yy_����yļ��f%�K�=�fӬ����&�[=��Ύ0�-/�  ,�+B����mҾ{ޅv�pN'g}W4�al�wՆ�m��}�e+�t��>� 
�
�$mv��|�޽�i����h��Z{՚�S5t����]�v�ʿ  �K F,\�i����Va�ZU�酳�^�{���q7^��f����c3������Ŭ�s0��4q�i�խ5
f�����q�N$���i4������-.�       t͉��ךJ5�F/6k� ��.F����S���{��q�N0}���&�[=����0�-$���V_6�_3ݐ �����o�8��깤�g3��6�l����at��}������  ,,V���g��p��e��Z�P��&3���8�I}�\�i���﹙�����wY��֎0�-*�t�ىl����m8���C4�a̩�g�h�2�& ��0����e�n����+�Χ�>��m6����Ն�m��|�y�x���m���       �l���/[׮�6�Hե�� �r�9y���q��^�i4���{�4q�i�Vh�S4����Ì�q����333k1k32��L-������ү�L-������fӉ{X�I����� !ZH�H���+��u&Y����[;��3���<�r�p��v�u4����k��-:�u�����Xf]��0�i-��w�8ͧ>��f�L-����Gq($m=��5
y�J�="L ��bY�k��uۮ)1M&�[9��a�e�_.�[1-��s�����w��i��       �4�Rk'.�ym,���S :S�x�I��{�ᣌ8�Oz���L�]���+���v�L\ۭ�R�?l� +�+��a�ZU���i���w�Ì�q��k�4���{�4q�i}�`�ʳl��Y��y�����s�s��_�W4�al�{Ն�m��|�alĻ�� W�B ����v�W&�|�i�����h�2�ެ�P�i-��|�s�s��:|����mw��z�}���}�a�e�_n�[1-��9�fӉ���śM0�} ﾾfffff       �^��d�bŒWS� #!��w��<�s�;��u��Il�{�3��c3���M�i���÷��v�]E  ��Z1,�;����Vw��fӌįz�3i�m1��{��o����Lgլ�/�<� ft�8ͧ����m6ͦ3���3��bVz�Lf�Y�v�q�N3.��  ��X�W�u��t_2I���m8�Oz�������4Ͼ��g���O�q�;�/��� �X$+Yu���q����f���Vo��fӌįz�3i�m1��{��3i�bQ�7��>�                                        e�77V��.�cN�(餕6�Vkm��^GW�Mf\�.�$��Փ�,��]X��jӥ�;x��Su��u���GGfWk�m�[c,�۬ߪ� C��D�B�o��fffff      5ڗn��i�L�W�mڴ�l  U�x���_>�����z~z��:�f3>��m6ͦ3���3��bVye�n������� ��k�ͧ�^������<gSL���fӌ���ޚ�Kf��{�g���~�feݶ�cU��usi�o��?'�Vx�u:�%k�L�c4����ף��r�]g�:�;��;����  )
�%xh�6�f'�[�Sil�c=�pÌ�q������l�c9�z��8�f'�{Y� ]a@��_�|wE�H��|w]��^��f�L�c+��fӌ���zo����ry��ׯ��       �n�6��I��F�Yt�9�C $��]]Y�l�q��{w6�f��{Շǂ�ڦi4�&2�����6�f2��I�U�Z
�;��;���ӵ��㳌���6T�[6��{�0�8�f3=�\wN���{d  
��mv���J��3I��c+9�ގ3i�bW�{/��o��d��mv��|.�  �+-�\�¦�ٴ�{����1��Uͦٴ�s^�a�q8�J��3I��e��� x����|w]�Y"c6�f�^�h�6�f'�Y���ٻ��$���n�|.�r�j�  	$     NYP��M�<�i�t��f c���YWW6�f��{Շ��1+=t�&3I���;z8ͧ�^��f�O�|'�  ]� ��������6T�[6��{�0�8�f3;깴��t_;�a]�v���� ]�b˻��s����v��ٽo�z��Q��deA�(���J(�J"F"
�F�$`��5��J�D���Q��H�hhQQ�
�h�T0F)�D��AH#"H�# �2���D��H��hDj41 `�`'��H@����������O�� QH�������]$�ڵ�j���=iO �bE=j䎞�$<jH鶺zcm.�h         � �[�-�xض�&U�vL�D$&��k��Q���׽֯�=j䎞�s�  (� Wx�xԑ�|�U5��k���V�3M]��@ ���z��=j䎞�5$<jH鶧�` fb.�1cֺI��k�4�k��z�$���]�l �K (AOZ��5�6�I1��&6��F         k�ZѴ�u���z�y3t��  .�V,�j׽֮H��W$u�+��s���|:xҋ� .�PY��SֺI���Lm�]���]�ֻ�� V,B0�)�W$t�� ���:m��cm_�  ���%�Z�=�j���=j磧�\��֗�� *�$SƤ��k���]$�ڵٚj� �5.X� "�Wy�                                       0��I�Nۋon����r��ۖη�ꮖ�i�:r��u�]�]xӵݭ��l��%�΍_.E���\X����7nM)�t�����^m�<�;�<��<���       %ɝf���Y�]j^�F��0�U�- )�W��t���:zԐt�#��\�z*���� ZE�,��x���o��7�Y�o���^!�������N0&��	�	�{_ffff	����^�8��`N0&0'�}��8����`L`O���@�`N0'�����	��cw^���q�8�����}����ź�̻˻�@�`M0'��V@�`M0&���p�	��q�1�+���	��c}����	l	������3330�1��5q�-�8������V@�`N0'��Ր'�	����Ր&�L	���� M�&�l��=���{       �Yj��u������i� F���޼�q�6��`L`J��j�m�8����}��j�[q�1�>��p�	���cw^���q�8����{>�fffb���m�֠N0&��	�	Y���o�sڭf����֯�=j�  Q�v��5$<k��6q��L�j�fi��}� ��,cW$t���:zԐt� ��S�0 �1if,z�I1��zf��?f��{Ξ�0�         6ݣ��v&�%�v�X�,�` �@*S֤���IO�鍵�Lm�͚  ^^�ծ���\�k/ǝ=j䎿9������5�| wJ���A]ί�m��cwڬ��h�P����7<���^�솫O��S��� bĂ�OZ�#��IO��5��j�H  $��RŏZ��j��+�UXvc��t���GOZ��           m��:\�[m�]Q�-�N�`n�,ň��IO�鍵�Lm�^�����@ .�U�V�5}��ڹ#��IO��5~$  �$P�%�Z�&6ծ���^?g�)�/�=i}� *ř�h�S֤���IO�鍼�Ur�T���g�  �B%�j�fi���:z��=jH:x���       ӝ���n�p��u��˻=|�� QE��Ws�Ǧ6�OLm�^���]�i�N�  �HOZ�#���_HA�Ƥ���t�jyF fPY�,X��]���]�i�w=�OZ�#��\�� 
2�h)�RA�ƺI����j�fi��}� ��,XƮH��W$t�� �u����7[���}�6Y�a�T+2���k4� ##�H�O't�t�<�O?��          ?z                             �L����Iۣ�_'/F�*�V��2v�IK%ۭ�\Y�Wk��5��ڵН���:*�4��i&�t�U��k����2�
���*4`�cJv?.{����       u�&k%v�t�nʶB[� &HK����o����Z��5Z�MW=�OZ�{` !`)�RG��XԐt�cmt����٠ e`Y`��Z��5~�d����)_�|��RG���  �*31<k���]$�ڵٚnUR�~�5<�� 
�1`Yb)�W$t��#�xԐt�cmw�`         ��Vk�٧l�v��-�D�� ZB�1bǭZ��5Z~�5\��=j䎞���  �+X���o���ǝ$���&6ծ��S��� ^*����=j䎞�jH��5$<j�H BX�ǭt���K=�i��f{���q�9\��t���>  �X��OZ�=��I�������}l����Y\�]r�SѰ          �5�㭕W�cmvX�7��<��= KB%�5k�4�~��=j䎞�${oy<� e�1�:�zcڮq��&6ծ��U��'�)�  ^$ �S֯�:zԑ�\�r��\�W+��U}ʪ�r�r���ncP�cmO(� ,��a�Z�ٚj���j��:z��W$t���� VY�[Ƥ�m�]$���&6ծ��S�         e�k&k5(�������wuP  /
 1,cW$t���g�}���}��m�RG��� ��­,z�OLs�����ni��}�j��:z�s�  ) (AOZ�=��I�̪��U;��[t�OLm��f� ��,cV�3MW�y�֮H��r�UT����K�@ �T���"�5�l���鍵k�4�k��5t�/         ۲쪘m��%��U^�^z��<�[� W������:{�H鼒W��z6��@ 
aF$�w:�3_*����j��e��=u$����d  �� ���Hm^��۪��W�n�W�n�s�� �x�1!bܹ�G���[�$����U)&�^��z  QI�^_W�n�T�����}ʣU��G��j��I	&�$�0TIH|QUD��R��{=Eޔ�Z���w�Bؘ��XE �:�$�B	J����T��T�늪�s��cu4Ϻ[��y&��ܽ)Z��:%f꧝�2.��ʖ��B��Ի���~)�n�_�N��� UQ>D2  S�J>���S�8�6��g�.*�EU1����.JX
+�x?������W���p�����p�!}3�B�����9�M�" � j ��
��n�4Q��9L!Zצ�����>��DUQ4����c��4:�b@�q���03�y�.�<�wέ�yUD荌B���{��o��O����ۿǉ]O��=����hzM�� ��hw�v�w��}Ǉq�>Q�/H= �
p:�UD��c�$7�1딢n���9�11 ������ 
]5�bT�k��! $*"Y�B�fZ���j1;�Q�zS�����`p첚X*��>�p�y�������7��v���F�Rpӫ��v��x'߫���v�s��qUa����/�����8azj�h\z�B�!N;ޕ�8e��W���_�0UQ6��6�t�g��-Yӿ(L-��,Qr���UQ?�cW�Wb��][�Ui���N<h�)}e������u�c�_���"�(H[0$� 