BZh91AY&SY?�3���_�pp��b� ����a}?TP���� B��M�q4� �٪(:  @�P���P��P��T�E� �@   (   @� ���$ U *
!*����      @%@��(�       �

( � �E����Gz��Y4�����}�p<��A��;� ��\�_'#8� �;�TV&��`����8��LC@Y�N����R���N�ӭ����� �  �(  � ��w�OG�w^����R�k��J� ���Y=�NZ����j]n-R��7J�[��u��z� ��J�s�Ծ����R�{��R�Mu���/[��ʽ� �:�e��rk��{:�Z��+� z   �

 ��JYo��W�w^�x�.g'UL} �=�U�w��y��eɪ�w�ҫ�}���b�3UϷ/>�P����nm*���4}�+�rk�\��^6�ۤ�� {�\[֕ɯ�ί}�U�y�ʯ�#�    � � �V{}yW��_Z�ZUY�J���Cv�6���Zr���*� ,�o��e^,�� ,�ɥ���W�T�U2�ڧ,��hsn-*�� ��bԫu��K��OJ�(ID��    � p��}���e9j�J﷉�����L�t�Yw�<�u/����������3�rk��r�a�9rU� FS'vS�]����qe.�}��+'�������e���^         �?P)�J�` 0  #S��R4��@2 �E?��T�SL	��0#&4�=��)6*�4 ��  S�	�R��@  hh !H@�"�BaO Bz��4{SQ�<���'���_��K�_ӯ���=���׾���(���j��EWJ�
��AEU���*�$�DU[�Y`��������@QUw�?hEU���/��Ҥ�!)�h$�������o���?��E�'-9��B�,D1դ�ܾ3�Ciesrꓔ8bb��R(H�C��M&F��BL��%��y��UH�V{���T�0b����g�45a.F����A�v�8�ZC,(r���2FCs�05.RF5�����g0[��,-�ƪVVڭ@��P.њ�ԴE�o6p��-�40j�0���(%��`�V��|��d�L�['!�4��c͎I�����-ᎎ̰!S�X�m*"Q��՝��<پT"\��~Iv]vZVs�z��5��yk�'��V�E/�7�W-�}�.���ܸ���8z�q�7).����I|EھB��׃���K��p巃�ZGk�mr>n����k����]���y���/Hg����V�,�>m�k��,㵸�JÒ�M�&sV��o��3��C���TC._o�FQ��qb0{T��Z������
\�YNޡ��!	SX��#�劕I�]{W4S1a��W���0]��=���ڗ�����Yo@R=�lx�S[��2s���ܴ��v�%hd��hb�9x��k	BdN�e��9��w�,�	�h� +^����i`�\�!�K���f������J5�kP���d%�	�9�e�]w��W_��.�-d�>�_X<����W��'<��~;��Ļ��ݞ��E�i�T�Ӣì��G��u��j�ɶ�C��՛���".�T A�CZ+�ԹJJ���2ҐPe�,Io2&�����x�{�列�z�W���]{�w���w��^Q��NBX%m��M�F<;m�.��Ոu�:9'S*1ٔZ(J�Ӆ�R�YB�xB���ӜݾP��w��ލ��tx�m@h�J�]���{',:�!;�3n�� !�:!P�|��R�ўTm24�u�5$G�z��;.Z,lv�+�	��<���Ćl��I��N����5���}�fwugJ��=�G��-[�9�	�!��e�1]uP��|\X�֚{��D2�^ܻ2X��s����\�/V����z���_��M]�j%Q1Bm�4������І�q�I<p	j�r�pe���������d��pC%��^�[A��	B� ��˾!>����F[$��2�8��D���W%±\�h�3_�ūLw��7�_l���E�#y������p�@��VK<�d �pqBSN���O�n��Qe��o{K����"���� Z24c��)D��$7yM<�aa�����"2q�)w��9�w��R�2���ka���X'w��S���.�2^� DW��"�S��w9�!*�����kw�v_5�wri�sno9{�q2��Q��TՓDQ;9�כ�!���G)͹i;�ZJ��q&J��j*r�E��%��uc%������Jeݢ�LH�4���Y�{9z���DҪh��8!(�|q��1�U�-��y+��}��[����Q14xf��UQEYm:9]�W�ɫ������j�x���C���_�(J�w��.s��c��!��
��$I��tbZ�T0QD�Tn����5󦚁K]"���v{�摥��qZK��ۂ@�u.��C1�����8[<=9���%����%��仼4P蛵w�K_W{��b�9[J��:��c1�s,�2��b̬-yj����P�{�<����N���)R��F0�a��ĥ㑉9ѓ������軍�1)�wLB���ԋ@�9�U��h�]���[��ՓZ�%��W=S�Zyj��[��&&�������;N��c�����������ú�.��ʚsP�	���7�3vB�bݫպ���g��M���Xaz��[�4ƳLh�Z7MN�9c�oV��Q�~:�V�q�5�]ov-e�UY&����v�_}�s��qjj�K���5�+|���1@Q�D$�d21�S��>�ol�G>���n��E��^��$�s�7&��м�P�Mm��Ӈ�V��b�M��I�Ӂ�5�̷��}z�/�A�oX��M����G��C�3�3z��yh�u����I��E$4����%w�R�UՌ9l1%͸�	X�T&؃��B�SNͨ��D���*n�J�s%1q*����7����8�w�5\�&�Q���_+r��9�#��pb���읷�@���PI9���
X�s9��+��ɦ!��!K3�Y�o���5�����HŷiȩZ�� �&!P%Bi!�	Ct�I$�Rx�oe�%t�V��\��OPy�~��*:YB�*��RǕ8�@S�l�¹X��u��N�	x���aE�&]�R�V�^��������f�D��J�z���Z��ދV��8�!ngT�{J�"%E[ǒ�Sf���>�1��y���g��Vc��3|`���0���{����a��y��Ok�o1��=i����ۚ��uz�ı���NTx�0�oy�udZ���swm�_�����z�n����y�M^�[�t�I�7+H�9�X�;���(H�%�W�8�W3���blT
3�����Zm8j��A��E	P�5VJ乺r��oJ\D���r2\��3#NӸ���uY�z�jA_����/r�]fg1kC�W� m��V�4
�4x��ܡ��7d�_U�]���!b1U�����f�}7	BR��9��4o���d�,�����n�ݥ�����#MjTEQQ"�D�PGZ�DՂ�̸"�(�N&���J)1o8������e�5h���}�:Ko7Yj�]�,�3װ����.m`%:=�a����/�(��/>b~��G>A<$�K�g2�f���%c�U4M�%*�M���I�K�K�2?f:�og3�"��)����ldR.+wwک��~���K��!�j�d�RI�
��@�*BmG�7:�G\����x�G�'}�M�Ú8no�B��<�y�K�YąXI1�ɫ1[�L�Kc�K0�Q�5D��D��/R��c��o���O���Yt����W�N��{��}�Z����A�����j�P�3U��{�qӼn�G/�e=�f��Q�(�Y�ʿyT��x���P�{j�w��R7^j�qAf<\�=��9���~�d�s���te0j���-R�VwY��wfR9V�Ǻu�$	$�Z�.Zg���ģ4��Y�Hk����yC֋Qs���(^�ӛb*�b ��1ƭ8s�I�[΋�뛮�!�
����iÈFbFmJ��Q�zzDs7�����#8o��p�=���aF��'z�h��q���,�F�x��<ل��K�\�M)g1��&�^[��k��|,G|m�<�P��u��,�@a���P�%�����0�!(JN.N�$��x�L��$�3�3g-r�|3V���:ua��K�A��Ld�Mj��os�sC�ü�!(MN=�X�\�!��	���X%	�JCy	Bw�!)�'3 ѐd����;*8n��j����'rj#%ۑ�:�	�i��%	F�d�w��H�%��ްdÌ�v�24Bn�Ad���4�&�p:����q0.��v�!���P������oa�'�bV�K1���wH+J�$������^E�ok�j�E�d�\���Oan�9���b�槧xw*C+��;��X��}T�Ѽt���&'Z�xXl:wbb�6A�jL�6�XӳG�gU���c���pu	BP�۱�9)BP`��7	J�y���Xw�[�R���������j�K�pc-�Q����SN�s}�V6�w��ڲ��"EL������'Cd��n8zh��g2�a̓!)1�[��F��)���1Ҭ9˻���,��C"f�!��Zu��@�2R�ue-�y�3�0K��0JM&Br!(�A�	���n��R���1w�ox���KZ�8�#݌����l�NY=Xz������%ٸL��4sX��p޹�g�i����8�.�`Z�����:�'$��JN�!��"� Sq#��{��v�R�\7�3P��t� dĳs|#����z��I�A����:s[__!ܺYhKA���C.A��2$3�K(�,��zs��7�{+0�������fʱ:7�C#��8���5�y�-ǫ�^��9��0NV�#���P�9���&�{�jph1�������MS!x^u�y�=v8`l*��26lubh5��H{ޱ��4����N3e�e�9D�����0���İ�/,�8RqF����(N�@��C@C#͗���y�aX��Bq��|(x`c��FS�y�:�ƅUh5J�T���]�l�i�#X��j��f����f��o:���ts� �h�@F�KI��J0 �dmf	�'�CS�9i8GV�M�PcVBQ�oX:�����`�HJ����e��f`�My�rq+"g$3 ��u��E۽�zr�R�O�r]��V�E�<��~�ü�1�c#8dc�R���2���%&��N,��$P�[��w�z�Kق�yu����N�)\D�u�sz��x1${N��Yt(����t�ޏ��'%�gZ�f��ug�X%�`5KE�A�]�j�M�`2����}�밂��'KBS�����AӴ��UlA��GC��R��,TnŌ�'*���2�F�s�\�ɳ�N�0JMA�`����;��Ӛ.q������a��B[z\�`�LN�1�:�>��,��:�s�!��1�N�{��7�����kA�d`A���\r����t��F��98�5l4S�I�N�����NBPpr��EN��6{�؅.���"
����%��2C3Hfhɍ���84C�Cen
���1�T5I�ʌ�$��ĭ�c��OA5I��a�b�����0�F6j�ST�CZgu1r2MV����Ӓz��.A���a�\CYʭ��]I����Vs�Yd9b�A��Z8����惆��P�%C��� ƇIT�3|�7!I˳�v��bj�r��T���zN�F.�Da�VM�h��WEDQ�d���%8��a��'����vG,HU;m�g'f��	4b�!�)Qt����W/t�J��)+�����+O����� �1*B&�a9.�'112LL�S���nI羙�14�pe���$ �" �g��V�s���Ν��=�G�����_�����{���a}*� $  $�  ��} ��l	r� @ d  l@   m�W �h �p�    l :x     %��ã�6ٶ"$�����f�6uv�:g7Pu�.^�c���*�'J�+���H�C�ۥ�#��H��z9�K8<ET��:�H�Eͺ�,/�r�0c���ޙP�[�d�m�ݬY2E֩��[&۰�6��渲���h��彪t$�N��*�-��B�r=Uc{U��[ +��d����-I��`*�쵶�s#mSh�� ���;�q��v�\>��+Gj�j]�f۬�r+�xY꾯�����tβ�U\y!1`�mzFK��EqR����W�4�g<V�e�4Qf�;#uAѹ��v�OU�P�=3S�*�67)[�����RóP�WuH��뱎Ȝ�#�)�n��8/m�v�:��1Zvh���B���kD\8ʫ����Ö�t��*�X ��W�C� ������c����ʻ�ݱ�\m�h�դ�C�Uc��!����Xx����Kw#��Od3�ݸ��̝x�e�,c�`�s� s�bg��>;��v�q�sRn�h@�)��V�J��M����	Q�v8�<�E��Y�-���`�C+��x)ͮ�;ij�ҳT8�m�z6�S�L[����n�6��d���x�	�����P��	���4�gɝ�1�$4\����3Ԫ2�Q�z뎵��&�I����c=�Y�l]Bi:,6�[VQ�t�q.WFۥ�U����A�ӻU��ci���x��+�9�ޙu��!v�6�EY��8h��1����f��\t:骫�P��I��3p��wm�T4���u��m�9ٍ	��mUn�t��:��9ܫBm�Qfv�*�����[�v��@<�6�m=+��uO�=����㡷Tc����Nw�k��<Cu�F�ۨ�3=�v�����<�6s�A����\�9�e![W*�8��h@����^������5�ɠ�g8/�g�^�9�z�dUڶq�1�c�t�˴�\{�����n��Yv��G,�#s�f+�켨L�n�c �l���2�KY��ŧhjڪe�� ��g�v���;-��jcI��[U@�P�PYj�T �{4�{g�Z݇�*ڕ`6�S�U �R�!��U*Ԭ�N�Վ��v�-�ՈU:[j��i	 �#�WmS8e��ن�&�+�ƶ,�o)s��MT����v�1v�zT�<�� g��չ���y'���㦌�ɢ3�z�B�;��'Xx^��7�q������2�M�.�g�Ե�v�cN0Y6��)-@j����O;�W��%K<����\�������5�3F�����g�r�+�����Tq;�q�ft�v�W���i6��PF::�H�M�F�5]��#��Fv��\aݔ�vh ƃCɵpn�v���;c��������	Jэ��q�e�q�D�^vz�U�Q��e����Z��ܞ1�9��p. �:^��ޙ��t!��]G����l�YA  �m�pvҎ�f�&�T���@U��9m]�ڨ�֘ ۭƚ��WiV@x�N{�gFΎ�յH�*Ѱ�����ș��ݰ[mUJE��nEsN5���pZh�<����Rѣ�Z���tv�̨.JpŲ��V�V�N���D��5�n�Wd��6;5�
]�9��b�UVڨ'��*���oa��8BN`:��h!���amj��Y�rl^��P�p�v̑!2G$]�Bw[^�^;U�t�Y�z�d�-������FT �V�HT��[m��i0R��m��$�v	 �v�-��K�ٶ���[VYm ֤Ã���vٶ��m�@ �Ŵ���N� �f� ,jXSMc
�UJ�������d�9���/P�$  �h���!vE�� k� m��ʵmT��J�Y�	Hڤ�21����}�  [A&�H;mٲ�[@ж�[v��b@���݅WF�Wg��J�//]R�B���9�'���ST�q!$��ҝ`I;Y�dΣ���< v� m �6 ��j��o5�_m��t�{�xsm� ����`$I�  � HM�٦�6i�6�'@�6�m��a��: 	 �i����H�f���	e�i�  V�v�b�j�gN����4�k��m�n�N���� �ڕUv� ��Ks��S�(	�[%�6��m [v咤6� [Rʑ� 4���ӷ2�: [@$[@i�*�k@���m������cZ��&�K��v��k� pm�d�p mZۆ�f� H �&�f�-���-��[x8  6�m��q�@y��-[v���  ��  pm �m�  9��d���ѭ`-�!�mt�i�b&4��tv�U��z�z�dmThU�J�-J��mRXR��&�8 �bڽj���iV��W��<U@J�a� 86� @�յ�$�@Ht��H�킳�P��I 	 -�8 p  $p [@  �+U*���/�V����h���^���-�(� h�K: Hݴ��:ND�l��>j�~����i�����*� UU�ZHU^6�t��+��-���lp���j�5S��� 	`%�%��ԝ�i0  m��&m�YmkՀ$ q�m���i�k�m�T�V�jr�^��r&�	�v��%,U�j��Pm�m&�7k�  �%m�mpm�	�\[@��I�vں�.̫]U�]Cv(	W�ymӦ��f �\�eU��T��*��u���œ��nd�*�v�PٜV�c���m�
��Ȼ`K��l�L������燂UV������]meÎ����e��0I�pIVF�i��W�T�D;YE"� 7j6
���ʥ��Z�'�nи�� 8$K�S�gÏ} ݥ\L�<�P��k��V���p�  � �cmؐ G����$�iYia$���j��e��G �I��кU7��'����`-65��`�Z�*��S$�J��$  @h     ��  u�   kX�m�  �� l    6�z��n�L�Ž@5�Uf�h�s�m�  �m�� �6Ͱ y��m�(p��-6ݶ�l �+�����8[@����6� �   	�6�  	�+m���   r[�     ��   ��5��շm�      � 6��  6�  	� ��	6�@   $�i ���  k-�� l�Z�mͮ�    ��u�fՁ�m� �i�����m��l���h-�@ ;m�m[q"@86� ڐh �`m� m�R.  -��  $  Ѷ�p �ۮ�	�` $    ���Ā�	�l6� � � m�����k�H m p� 8 [�����H6�m����  �m �m��m�m��   ���I���k3 ��   �Ħa�� @$ �m�F�p����NP۰m�Ā��ݶ�8     ��  �˦�v����5P$�׭�ހl�&�5��m�L T�mͲ�.�o7l�"C�r�t�� &��m�c��˰;v��޹�çI ��e���I��W���N�l����UA��UQ)uJ�t�+�S�� �N� ^���8��  ���[�n�.IrM�  N[l��i0p�8 [\  h K��/[ �h�^�6�F�6��!�A�mZUT����!9J�#�� I��v.V\F7랶dmԴ[m�A��K��ȶ��3O����m���]/�uH [[������r. /Ml�Y,�6ݤ���� Q[]��� g9���B޼ 'I�m��Z�j,���m�m�� ���[�N�T�A��PqmUUa;*;������H�m�%����A�m��
���wN�aU�i�[4��Z��m�G�� $�.iRi6���Z�,��ZI��I+fC�)l��6J��`"h��-����� ���[Æ�N��E�g P��l=�+��Vԯ  #�okVu�V��8��jd�_���8snͱ ��[�ۣ�Ʒe&�,/��OFו������cm��`A|�q%�vͶ  �u͂EU��T�U 06(� ��@�m�,�M���l  Q�WP��������@][ڹ�@h.�c�UU�Uh<m\a���*�]���� l c���:�gK% ���.� �d���o  l�Z  [Cm�ضJ�k(�ܨ.�-@UUU@     � 2�"@ c6Z���GP�Ò6�	 mMI��H N�4�U��׳�$�h	�;k&4�٥m�$�6��c� �I& ��$s�h'N �m��$n��� 6�ܰ� p
��������刢������������������3�������{s�IC�*��*bv�i��R��v� ��!$�R���DB@����"��=A�(�N/��GH��D{!0�Ō]�Px��b(���`"r6�"v";�:�h�v���C�����ګ)R�%0YLGp��@Ĉ\��\^*; u(@��+����= �(�Lp@�D6!�	��xt�$, & >�'�� ��ҝ�@� ��
;����`� �& ��:�E��@� t��;%�c���}м�=^�ti�(8���B���v��^�/@z��؄�8>�x)Є�{����oH���@p}Pv��'�z*#�t�h��z� B�b�� E��E/Hl�hJ�|B.��%E6��Ǟ��<S���T�p1��A�`��`��� 
��0Ď�Cb��� z�H��@��}Tx��p�$����� ���$�BF����j XH$OSxqb�	E�A�p; ��h���蝁(!t�j��U�@SF ���pv���>����P{TE/K������C����(30�*,�%�e�2Q�̘���A!3qª�"I2	�J*����_N&T���S�$A@LL�ؤ"�y�J�D��>"%2���� yP��3WQ�G 88#��:�.�؁���
*vE���h(���G���5����������M)�/���b�hL ]F�14C�Z���K�0���b��-��)p	-�B:$р頀�$$`*T���D��&!�!M�{��?Կ�U�����nUT�B�EѵT���R�J�݅���uA�#�ܖ��n3ԯ7��.�8�F�ӌ[�mg%i�jxM=v���� �ņ4��0��Q΃�x�4Wl��cLݥ����;=���p6�g�S�R�y���p���m۰�u+�rk����1���v���q&�=z��M�����#*�ִ����N�4��׆�["6�5<jEɶ*MK���h�n��qT��<D�}[�糳�g�m�Z\��v�˪�@Y�ՎH_N�W]����iŝV�{tq������У� ��6"m��ײl]�;c��c]�v���֬��nz�e��	-�s��������2�Zw1e���ۖ1��.��+kt��]�9�H�m��d���rE�q1��X�u�N�)vxv�6K��g���<��Rź4:I^T�6�&w=m�d�:�3I��@�f� ��T�;[��HS����r��i��3j���Om��pG=��v�� m���ZI��WfU�%x�.�\Ra��T���öѭn'(��Uv�j��ү��ɤ�0D�$ӯk�-�&p�,��Kn�Xh��3�ڳ��8-��t��gb���7&q���:�ӻ]�o^z�3���<��FS`��!���SSl�!�F�s"���z驷l 9m5R����V�N�/7J��0�m��N�ͻ�-F�cBL�WM�� *l���%�Uv[�!4�<�V7h��e�n����%2��� ���3R�<�@+g�uF��r	t����Z��\�V��"ՖSr�j�)v�S��>KfQѵ�`��;��l�;k���i7)[0JM�q(젪
9@��h��s�;��g`z2ζ�i��e7����l���sv��&;K���%�(��鍰tj��t���٠��q��C�Zm���:\.���#�}jKj�^0n)T�����`�m	�^7Y�գu��"^�I� �Ku�t�^��U�I'L�vHm�Vdf8;���GH�� �����8Z�`qQN�J=�=�O�<���}=S}��dý��33��l�7m��4j1ܾ8ͷZ�Ag�h� �wh^�#�ňbkK�2�v����Y��(5��@;��fb;��:�N�'z�m���N:��h�WWn��F�s�ѼpJh�q��3V�N�m]����Y�A�V�9���@��,�3�j�YZ\LCخ-��nn-�ex��ml��=�.�$��^��zp�N�!�PB�n�wn�{�{�1�ɇ�&�`�U\s���1�y��vxۜ�x�Ӧ�:N��M���GC:����T�����UWunk��~�Ԃn8��)���]X�L,]�;�~�`r���j8�#��ӕ`s�0�1w�������]X�?<MS��HE$�����`w�ج����<�`{��H9(m�MD��y����]Xǘ�]�;~�:�c���z�v.@%�[;���#ە"/���cv���ۣ�n��&-��5u���m�mՁ�y����c�=��VϺ�e<��zѽj7���U׺������J��aޢ�R9e�C��V�s\�:�U���]X���Ք�MG$Q��^�7�٠3#5�M����j��>}J(+����)$lHq�`w�ج�&���<�v��ljA7I����a`q{1�^�v|���گ�V�6���H��*�nD���;)N����뱛$�DVp��r�L\�[B$q$G�8Vn��َ�X�L,x����rJR$�:����@}�:P����gsp��Q�)H�)7#�=�5X�L,ϱA(RTqS.����U�y��]�不n(�%JI��;�X^�vW���?b�}Տ)�R#u>$�����`u{1���+�Ʌ�fx�ۚ�`i�E��0�Ʒ��G-��v�m ��R��<�웆�]�z�ܓPl�����`w�ج�&��v�^�GR9i&���^���W�͚XY���̖�ϲ5 �R6�E`w�0�8�����#ٻ,c�V+=��ӍƔN2	HX^̘���1%����Z|P>Q
PUO�����,`5�5I�ܔHD��K���\��$��_�$��ޘ�����V���������������+'<����bӻj䧔�5�cW2ٻ3qN]6�rpc�V=��ُ~��� =����#QAԕ)&����a�-}��$�;�^$���<I.W='��F��G�َ�;�d�~��/c�Vsf�~�:�e$5I�v^oy��uM�����Ҁ��ؠ�<`GR9i!�%��?b�6����Ϯ��=��r��}�*D4\��h_H4�QGB��h�����DƖ���t��*�������%��$rLQ���z<��FR�xbͫ�M7m�p6i�٠3;5�{e[�qu�u����s�pq�Y6av�5�a��]y8gJ�Եɺ7Fn�m����<�&6�h��;oh�N5��a�b:�5��֍�{&�p[6��ۍ�.f���9�Mq�³	ft�s�}�X��$��N�+�m��rs�i=��(�0���܊YJ�g��l��>ft~w��y﬿m�x�]d��ѹ9����o���K�^�����ۖ!���C�˸^���H�m���w2i`q{1�]�v|����w+���4�q�JB��b��$y{u�ǚ��&�4��J��r�$"�:�����������b�=ט9C�R���&5#�����f���K�y������`������I4�V3��y�]|�$���<I}UES�}'�ܻT�\�֝ٶy�HCmZ�f�z�l���W�U�`�u�ۜ�6�(�4�0�(ȓ�8u�z ϳf�̌�^���n-�P��$���n�qKx�]�}y�	�i_VC� ���@�)�;��o�`{va`qfc�g���I���CnK�~�`w�0�9�1X{�,��dq�8�m�Ԋ�k꯾^�ޖu�2����`w�ج���\i�#N2	HX��V�U}����=�5X�L,#�m��6(�S�G!"C��z-�V�Ņv5�=�i�r��M:�p]f��
TEG"R�$"�:�����������b�=��(q�R:�H����G��K��U����`w=��"�(6E)!�������<�w8R���<Q5սo��׾�(=��d��B�$0�`sb��2X��+�Ʌ��}�ʔ�8�)7�w������X�L,,�vW�P�i�#JP�)B
M��-�B��$PVѤ��El9�����`[��U-��CnK�~�`w�0�8�1�]�v�P��n8'���X�L/R;�uX^�v����#ٛV��(�H�"	HX׺��̖�����ra`�̦�I�*H
E`�d��;;�.s��8�P� c�RR�pi�h���&Q)D���W ������>���`f<�r��Rpi�Q�$�;��V�{fj�Ǻ��̖:��ʐ$7�]��Ӻ�݌lMV�q�����7n�[F��pt��n�� h�عy>�s��,Iog��$����%����Ip������h`���b�����fl�=�5X�L,�ި��I���qX}������a`sb��ԱI �JA$�����X�L,c�V�{%�s�,�$�
G"nH�V=����w��`{�جA�'��P4�y�zsZ�#z3EmD�fٰR�:n�˺tqɹ��m͵��n �O-��\���E`�N��7GNz�//�q��ˮݷS�v͜c6r�4.3V��<��V�N{a��;rv,v�۶BN���O6�#���m���0�:{=���ga���܃�y���� c���$7	�8X�[v������y��� ��td��ۛ�n�6D�V[{1rfь�j����w��{��e�lh�I��˥����v�um���K��}V�nn8�L�[
J��,e�i>d��k�ٛ4df�y������T��J����;�d�;��V=��y���_������F:�4ܖ|����a`s�1X{2X�e%M�j	�%�N+=��y��;���X+�b��H��� �[^>�����Vٯ���ٻM����hD������y��<�OX�Ӻ��E���ә�c[��R� �/�Q(@�l��_s��u�/b���f����\����ｔ�G"rF�3Y�������Ot�e�J'���fs������;���<�ϲH�r&�v�ｆ��ι���s��u���v����M\��7w���ι���s��u����z��J���*)Ⱦ�}�u�/b���ˮyf/�����h��Ԃq8蔄���^� ��;F��(N�9��k[�����7$�'Q�E��{j���ˮf<>�}�u��6�PN
St�q}��e�}U����w^�{ٻu�/bگ��׌�)2�Q&$�^���s��A�ʟʸ|�
�����k^k����$�p�N���6EǢ]QD3ZE�,�F�1j��
�W��pGmX��i"C���(����Յ����h��2h�Rç}��ˉ�m���񵓣ìᙘDSeq����;.(��o}�����"�`6�ѻe�jz樻��(.�z���nc�fir��ЅBT�2��kYLBu�p��J*��"i�����	u�'[7sRr�+6�F���U=s|f��4i4�y����P���e���˰뽽r\˶;�E���s�`��\-T
�V^Y�XC���0kI�(q�
Ru�Tv�5�iwkq����7��c������e�E2��#Z�LM�%���3HRgk���4;`4���I>��
�GI�]�d���!g�t���6 vv�M�i�<�Q? ��Ї�"x(���O�P�E�@;�|c"$�p��Ё�!�Ț6�����Q��e>�]y�R������ԥ)�����e����z�Z��R��y���JS�u���)JN���=JP~A|��߳�R�>{��Z��὎]�-�//Z����z{�BUBTs�}��JS�����)JO<�^��Ԥ}�~�������ι$��nAD4����]X5tp8�N��	X��i��[��u�Q��z#�ݹj;����	U	Q����+UP�Q����┥'}�����w)J}����Q*�*9߾�+wv��&�[W��j��}��)JRwߚ���)O}׿g�):�Ͼ��'��%>�Y�}����,�wj弪������+UP�'�k߳�R��w��pz��>�^��RUBTw���,�� �\s/Z�����{�qJR�����R���k߳�P�����P�,�:����@|�5��y�ԥ)���VRL�Ӗ�p�]�P�P����+UP�����mG�=�߰�|�j=w�y���ƺ�#[[�xV�7'�p=49�r�.��Ŷ���y��J�3p�1s`M��?�)O�׿g�);��{�R���{�8�)I�~}��JS�_Kɥ۹r[ʡ*�*9��|��T%T{��s�R��w��pz��=�^��S�T$W;�Ï�ۊ�.ۖܗ���UBT�~��8�)I�~}��JS��ߵ�*�J�s��2�U	U��}#�ݹj;����J�����R�����k�R������JG߽��R���}�,�wn��W-�RKµU	U{�BUE��=�߰{��>���qJR�����R���=�JiRGFP�)el@��SV���݅�o-o6i�4���׫�8�vt�8�J������ݺ�ʆ�
��kcdn��f�F�-�-ˌ`�]��'pt�u�ݹ����P����;�&�z�맷#Z�v��WV�v3��*pG��]�����I^3�:sm-6�R""�P����>���8�� QD�!�/d\�vFUJ�6�`&�aeR��v��c��m��ږ+P�����PVe���c%˄s�uBu��۰i)��b�t�p�1��I���^a�N��㏾��X�UC?{ݷ����׿�z��=�^��R���>��ԥ)�}��┥'�����k7��սh�۵���)O~׿g)JN���=JR�����)JRw�y���
�>��$ԓ#����BUBTs�}��JS��ߵ�)�W$�����R��ߵ��┥'��{��cZ٣yk#,��=JP���k�R��w�����JSߵ���)��<��R���}�=�IR(�6㿾�����Y���R��H}�~�)JRy�~��)J{�{���)I�kݚ�}�6kn�״����Sh+X+�c(]�y�\n�G��G�;�L�j��Y,q�ۊ��ږۼ��V��*��k߳�R����pz��=Ͻ�\� d�'~g߿hz��/��>kY�7nZ����ʡ*�*9���+Qex��`�{�z��}�5�)JN�Ͻ�Cԥ)����⟅	rR�����Yf��f���7�޵�o�ԥ)�?}�\R�����=Bҟ}�~�)JRw����R��`�4j����)"q��PU}A�s�>�Cԥ)�}��┥'~y���)��[���>�����Z�P�#���o��)O��~��);��~��)J}�{���)I�y��hz��?(?h������vmۭ��=mȞ�hۑ�.�^ǣ�"��v���z:��l��}��ࡶz9�[��)<�߿pz��>Ͻ�\R�����R�����k�R��w���Սlލ�іY��z��>�^��R�����=JR�g���)JRw����������2���oZ�ַ�R�����=JR�g���)O�;$�H	�}��PРx�������;��U	U	�=��n+���[���懩J�>��qJR��<��R���k߳�P Ru�{���*��bo��ۉݸ\W�̪������)@~I��~�)JRw�����JS��ߵ�)JO���5�}�޴f�����u�{l���sr��[jD�1NL��0��;�w|}R1cJ������}��)JRuߺ���)Os�~�
R��<��R������Q�ov�k{�o7��R��w���� d���ߵ�)JO=����)N��\j�*�*>缧�ܱH��wq��񕪒��=��qJR��<��R�)��o�R��w���JS߾>������[��Y��qJ��<��R��}��)JRuߺ���(<�b�wE��x��}ߝw�R�����٬rٽ�FYf���R�����)JS����`�)J{��8�)I�{ﰭUBUG�*��|��]���.on|<��6 v�J�\�U�T��GO;�;pƒ6t"kVl�[��7�f�qJR��3�ߴ=JR���~�)JRw����JS�����(z���Y�����3[5���9�hz��=�^����)I����ԥ)����qJR���߾�Z��*������Gwd���ݼ�)JN��߸=JR�����)O�W$�����R���k���)JN��գR6�Q�Fۗ_p��
�����U�JRu�{���)O}�\R��!*�I����ԥ)��,>?n5����kf���qJR���߾��)@~BA>��~��)I����ԥ)ߟ}ÊR���P/r���@e���?L��eK]Fx�v덽�z�	lj���˷�>��\f�٤:P�p�W=���˯/�����LOK�"`�x�CE�t��K��e�q͸�x̯$Kj�A�m�&�{m��v�l��b�k����;��n�K���=�Y8�̡H�-Đ�VNgX���M��K��jt;T=���8�1�][�]wcs���ο��ﾸ��)���r�*<��{���������D-H�Ѣ[V]��CHi��+Q���+'/h5����;OK��]F5w������6).܎�q伅|�������YT%T)<�߾��)Jw��p�R����{���T%Tw�|��+�-)jIk*����~���!��{��)JRy�~����JS�=��B������S���-�5��R��~}�)JRw�}���JS�5����[.JR{߿~µU	U����Gv���wfRR�9'���hz��=�_~�)JRy߿}��R�{��qJR���c�n+#R�m��̅j��9���BUE#�~���JS�=���);�>����J����p�ЬW���N�i:��C�W)s	�W0�����Y�q.����o���qܵ.+�嬪�����aZ��S�=���)<�>��ԥ)����*����߾��)v��v����Z�)O|���$x��(u��h[=�Hk|I6���mH]�i@���ƤpGzn�gAod6�xU�	1�S"	�����`�P�`���5)I�3���)Jy��p┢Tw�}��*����]���K$��޶qJR��3�~��)Jw��p�� L��?~���R��߿p┤��{�}����j5^2�U	PW>��R�����ԥ)��ÊR�����2�U	U{�!E���JZ�o{��)JN���=JP�Y~���R���ϵ��R��{�)JՕ���D�#PJ889LU)T���'\��\�[\Cq�b��8Վ�n*�����|��j�hՖo|�)O|��R���u��=JR����8 R�����pz��.�k>>,5���[���┥'}�����? �Jy���8�)I�����R���~��ZR���ߣ��٭Z٭�o[�9�ԥ)���ÊR�����pz�ڪ�} ߰��ba��z�	t�J~��8qJQ*>���̭UBUG{���\�ݩq\{��)J�Iߞ}��JS�=���);��}�R��������)I�ۋAȚqD)6ܺ���P}�g�n��){��}�R��{��)JJ�w�}�j��<�~�.��j�%˸X윎���,YZqa]�l�%�f�	�uu�`��W9͘p������٭lݛ��)JRwߺ���)N��\R����>���u)J{�p┥'y�}kz�o[�kv��5�hz��;���p� ����{����)O���)JRw�f미UW�W��չ�P�J���I6qJR��<��R���{�)O�� �<�>��Cԥ)��p┥'�����;�޳yhՖo|�)|��R���u��=JR����8�~��`y�@	���D	BC�%JEL4%"�T�G�/j�Rk����JR���E�L���pE��*�����=>������y���R����~��)*����eP�P����$�H&�Ւ�nyǅw2��n��W2�� H�N��U���Y8�	�UQ-c�c�+�Զ��ej��{�)JRw�}��R���~��E�);��}�R��~֏���k-�5�[�����)JN���=H*Ҟ���8�)I߾k�z��;���pk�>��Z�m��6ܺ���P}���ÊR������Q)N��\R����>��ԥ)��0��{�{��lֶn��g���d�}�~��R�����qJR��|��R��@������y�͝��8��bbI&Z^��`�)Jw���┥�Q��~���R��߷�┥']�����R��[�⾬���$$�0�AI JJ��$y�� 4x�f��%6),��I%�S����'���N�l�E�@Ӱ�o�z�K}B�o1MdD'5ߛa�H!��U�t�k�[-m�Xspx�+��9�g���ɦ��$�"l��]�X�٠�b;cb�`��&@��CI���C �i�� k`rh��i@�D�������I���bXs�<])��捉Z4���V��gP��P�3)P���I	�㙙m���ݥwv�*�q�ۖ������ڥZr<���c�����?u5����G܆S���ˑq�=d��U�6�\	ű���0[�Vў�����Z�H{�X�����fH�#��@���\�v���]��Z�����wm�mٕS�/��ɍ�l��2v�`B������ہ;An�n�����<!�B��n�k���4c �׸y�Ƌ�;�]v�Ga�?i1��n���L��S���7��q����
0�7\ԏ;�����X�<1�8Ě�[��o\����>�_i���ݎC�{XO�V�WeP�E!5f��Ev[�˳�����mÎ\]s�8➶#�]�U��v�N��;l��Rd��2nت��M�ѥ8�Gl�9��kX)�@MZ��>��ڹ�Z�vm�∖�:�N%�"�Si�k\��m�����˚K<,�NWn�����탐^Q���]�f�ٱl��6͝�s����mD��oW< �4�@c��]ۭ�$K<�J�ʫ�'	ŵ�鴼� ��i�+ƽgl�LE�9�v���+�p��˳UJY$�ib۶n�l�Fۗ�۲�ۖ c��ݽpW'B�ܤn6���=;lU�	<��Z��]�x�c��Շ$^�.�q˳��h�綮h�u�d�s�l�' �f�mLx*�W�̭V1R��m�$��|��d6x��>
��r2�d5Աa*]��m�U��-i!�Ӓ]�M���lm#��J��s�e�&�j'�Je��`'P;n���U�Ph��3�'�i�M�`�[�v����p*���� x�� ��J5�qȷ���q���vGŸ-�] ���77VbG)��rk������rב.yI��Qvx�9�E��kn�Q0��3֎�1���u6�$]ldK�Zj�nqv���vYܲ��5ڴYѦ�<��3�����ڙ�:���Iţ6H�Tc��//k�(���MUT�-R�NgYfw;[E�j]���,�2�|}|wy�����/�����)��@:��<C��x�O� ��EC�z�ҏ�8���yY޿�gsz��RL����tiֶ���c���v9�	Þ�_6��`ȓ��㛛ll��sN{��x��n�Nձ����/
����6��W�ӹ�D�w2-c̪����lƫtR�Kg�/��s�Ng;�n��vw`Jͺ[Ȍ����\ T�J����h���+��u�;\g�V
ݗ\Fƛvn�$���3�U*ƨ�sƎ�[e��v����L�r7q'`��Ci����`�ڤ�q]����������i�ƛxM�1]}��q���珵�c�k�R��~��}��R���w��)JN��_}�=JR�y����)I���}}��7�6k#,��=JR����� R��w���JS�=���);��~�����{���Y�޵����)JRuߺ���)O<�\R��
�¹'����R�����ÊR�=w^���q\R]���y���T%UU���YTR����pz��;��qJE��{�����}]�{A��H�d�8Z��'~y���)Q�Ͼ��)JN��_}�ԥ)���R��}y�}��O.6��X�#������A�m�N=N�ksm�,N�o�������p�id�+UP�Q���T%T%F����Z9��m�38b��`%웦]�fH���vo[9W^���ζw�x��)C+L$���2�H���D ��2@�]s^���䒻�J���33y�;]47D��0�/2��=�=������U����}�SP��j���:VH�M���y���u]��%M@^d�{���fm�\�6��s����a�f��*j o{�k̍O`fF��/��v�&�`n:�љ3�{�;�=�u�j�^3Z���-˺�s��s8?;�����o��c���E��\��=Iw��<Is������AG�]���Հ{�f���nA\��3#S�y���U�bT��JO}_R�������$����)��}��>��.��V{XChl^
&fI�\1���[I�M��p6��sy�����l��j���{25=b��{۷`f:U��*�A�9P�J�9��<I���ė9�}���}���W�����ԃb��n1�6
���vڣN�"�v��#^��Os�|w{U�ٙѸ�,UO`}�����W`}����fBJ,n-���)�Si�`{ۻ��}����Ԣ��#Sט�(d�y�%ҍ%'8}�u`{�7_
�����p��1�B����)R�U��{ѩE��F��>ĕ�w��7����g�{��'Q cg�.*�t��ޯ�K�*�7�~µ��F���v�����o{�{uwW�f�SPd$��{M5�w%$��Dӡ0N�t���:rĵ�8j�ni��.-ɭ�I1���g���H����X�n�w۷V|�u�p{&���A=iț�A�9�>ĩ���7�8f�wE����3R��0�����D22T"r�����͔P7�fjW`}����4"&%��e�Z\.���fo�ef�v٪�������cM�⃀���`fjW`w���c5u���ٲ�a1S��&=��u��k5�޲�����M��Pke6�۱�v�;���Ѹڻ=�9�0m���<�n���p*�Vx����k��cm��O
O"�����z�^��6���0͕y����z��]{��c0�^�7Z��E���p����q�[��nc ���<�v�Y�.��V�7�m&Ĝ<puX�-V���*�Z����7d.�s�4����t�\�Y�d�S�UaFaij�.'b�O��v��L�!���Vs�	�[�B�m(S�X���˩N'o��#�(JK���u`w�R���G�8n��maA�;DC���	(��;��x�7Wu��m��zQ�+P�	$h��wo�w6Q@fjWc٪���!%��cd���r��aG�����mՁ�=�|�ɥ����'�r(��m˰>�T�33f�wG�f���Ԯ�+����5�@�R�!P��h��g��'Ma�8ͳ 0^�:�N]�ks�}'SmN2S"r������M,{7y\�ͺ�;�[OG�BE%D�o�wٿ�`��2��N�|0����u�@fꦠ>�IE�y��g�˙��y"X��"$�7Wu�f�jd$���i`s���ϛn'Dm�����SPd$���6QA��a�Ϻ�����6�HtR�U��=�|�ɥ��f�8}�u`ovd�R�QP"tG�Yݚw���M�
�L�Tu`�݆#��t�'qɝu�u_U��>�!�GD廷�;�P���f�j����	(�7a�ׅ$t���G���s�/���߮����36Q^f`��w�<D��1,�Ԓ�R\��a�.v}��VV���C�!V��P�Iؠ`�Y��X�n�f�5R8ԩL��Py�}���3ef�v�y��{�V����BE$9r� ��i`;�jU�bT��	(�9�d'n���9<�{gױ�u�cn�p��c����\V��Bm6��s�S��):lr(9C��ۇ ���>ĩ��Q�k3e��B��n)Dm����ݺ��;绯�{6Q@fjW}�o?��mn~��p"fZ"gy��3c�����E���Ԯ���XzQ���8�'-ݾ�W����^y��u�]���9Q��NÈ}u��=�_ ��K~6H�'!$�U���]��%M@}���3U5����������'nh�]n����#���sr�u���S�ty�����{��Y�""k�3{���Q`����`=��� �)�lj�p)�R��`{�R�=�`35M����R����Ǽ��_����BE$.\����,y%v7�b�P����!����ZZ$DD�y�ĕ�b�P��� ��e���j{>M����jNp�v���%��hĕ�ޖ�7��|c�p~�n��vݽ�ݠyc\�6���T����퍣��G9Bm�od�Gn;S�J��W0�ì���nY�.��k����/=C�sv�l�_���w}Vh�{^rt��k�\q�К7
�'i\�*!A��棰8�E#nګ`�i4VN�X��.��r˴��ڍun�:#j`�k�5G�>K׺Y����/M����ݺ{&.��B�g�߯w���??6���C3���۞rs����Ѩ7C���ʳ�����cI��^��|}��m��"gy���J,3T��+���n�Xz��b$���v��f�7��I]��%M@fBJ/��fwû����g"^f^Zffh�]vؕ5��^� {ٲ����Ԥ�6�h�D������3�IE�fj��y��WԳ?o�pҞ�#u#�D��F�X�$��f�x��4b�vؕ5ٝ�7�~�޵-G�[x:��qu/+��^^���l�2�>r)Ӭ�����SV8�����7WM��]��%M^�{�}����k��+��:�朖{���*���C?h2���M��f&U�0���v�%	kJ��*b ���(ǁ�o�p�]�:��35M{����gͪ!O�!�f	��Q��Is�}�$����=_�� QM������`cc'T�L�<C;;̵�d����h�Z�����f����C}���cW �Gr� =��`o37�-U`}�Q@g�)=��u��A������l8N����?9�����`�5v�۴�J8؇����{�F����5SsL��ˮ����ϲR�=��ut��_�5�)"�G ܜ���,�%'��S@}��v7����i���v�j�]�o���+�8�̐٭���h�f�o����8�(�2��!��S�	&,�@�-F:�]��i�R���@�
i��>�Î>�'�Ό�Cp��ތ֛4c��k�^bF]t��5��" �y�b8�D�p�K\͇dd�09���Aj-���9̫���]b�8oF�@]eZ&�!
Ň,�(��-m�ĨJ�Čc͋_ ��Z�������w��</4tx9	��:!C�ޢ�!��(���Q��p�mf�Xt�9�N�d&6��)Ep����]����A}0��&�M��p� ���⽈x�
x#�؃����T��B���H�J<Ҫt�N��{�:���Ձ���R���RG$'˵�1�TP|�]��%M@g�)=��&��W%JpT�n+���p��,w�up^�vꬬ������F�A��%�v{pH:��C�td�:m���y�q���C�;_*�;�:n�REC����6~,}���	�Tw����]vp��$��*I���}7W ���`w����ͺ���C�=O��Vˁ�\��樠>�j�9��a������s��J[I�)9"�GaTw����ϸr�;�}�V�IHUXs��5���Ԥ�InnNp�mՀ6}���	�TP|�]����F�y�{~�v+K��QS��weyp�\I"ˋ
��#�z�g�t��qZhCq�t#���ksg����(�Z�����g��G�BE$'˵�5{5�|�]��U5�d��3Ԛ�^I�N
�JG`w����ͺ��=�M��5{5��ul��u"�*4�8�����ںڀ���{>j��>@��$�B�prn�ėy���/�y����@fr�j��+�m���.��N���N���ƌ��D8��i�W���ŷ]���5�q�A;lc�Hs���{:��v�ؗ�R��'e�����J�kqv�H��/s�؁�b��n���c���h�m�r�.��:="��ۮ�h,&:�n�$vZ[L��nP�(��wIle�8�H�[�={=�m��L]��D�@n`��t��cO=V���a!���w���}�w����W:u6;��'A)�)�@m����n��W2���	�)�v���yz˓����||�g羲��E%�\W��v{����۫���\��%�6�!�$UH��Z��f���̔��>�S^�x�X���� ܜ��mՁ��n���a���j�39u�H50�1 9NSr�w�up�͖{����UW}�u`s=��N9Du"�
��ڰ�T�3{�o�Z���5SP�JO`f=�t҄)4&T���tg��Wjަe���$���Y�)Ȯ�IJ��R]�K���n���}�$����2���}�,a��|麄�* 4�8|��ٯ :d�&�bBU=^i��3g�����Y2���S@}��|�6�$n�t�)*��}7W >�SA��|�]��j��/�b5e���$�k������\���p�%@���;3 ��	V�jRrER��4�-W`}�����ҧ��T�x��6�GHU)�
*i�Jq��) u�L�!�tc[��n�bu+~{���嘦8���f�X���}�/����p���T��)NSr�w�S�٪h�Z���5SS3{�DK�GR) �>]� wٲ��w7�9>���4t �|��G�t����w�up��i���*S���`}��v٪��ϲR{��c��4�]BB�����ԗ;�Ē*��:�W ;��`w���짯i$�7IvK��{<��q��YŶ�¼n&�s��C�:�s��I�$�	�I�&�RN���$��}x��>����)UIw�_�.tĵ���Wwi�%%�\ �e�W���o8}�K���\��%��r�#�*�$���w7��ɥ�}U_���}�,�-M=�8�q�7'8
���bK����Ԓ�}��^��A*�R�!�߾������z}���I�%���bK����ԕQUK��׉.wsy�;�۫�0��	�EN :��׎�0V�ti�Rӹ-��Ӫ�"��{���v��w��U���7Q� �;�\ �e���U�f�h�{���p�=�`w.hx��Yd�Ɣ�x��>�ۿ��5�}�
sg����5��31�fp����h�����9�=�����}7W ;��`w����-�i�&�RRU���}͞���@}��v�����W[X��_�K�R4�d�-p�͖y����������O`cy�!���HH�`��M(C�J����ݽ�_�����v�!i඲�6]�'2mog���Nm�h:ɰ�v��8���mm:�qG;�[�@��b�x�pZ�������͜��/�t\�%\�8y��T§M��<�cm�	^A�v�W\��s��RFh��̗��؝���kvN]�b�z�b�d��9�l�Y�b�����s�j��vz_n.�eݝ3�TFa�m�%PdN��F�����U^#���wZ�k��6��^{H7a����Wn���[��-r�J\x����&?W���m�L��
�$��������mՁ�ɺ��f�;�P�I$R9�H�v٪��=�f��{ �]6w7y���el��p��A7*���I���4�R���M@}�(�m���II��p��6X��� �5SPw���3�S��.懀z��rS���`wsw��ͺ�3�7W ;��`sp0��إ)M(����Iy�:M�Ù�q/`�t�'YwR��.���?^y���� R_ �n��M���6y���᜻����D;�D�H��｜��=��g]"�ȴ���>�	U�����f�j�a���ݦ��q
2K���f������/f���76~��� ��m�d��T�$�G�R�3U5����>Ħ�ߵӍ���(AG9�=�۫���ۛ�.�{?~�w7y�
�u��MTq5��c�d�pk4o0��rt�`Ͳ�0��룯��*�;��S�R���r��M���vX��� ��n������I*	��.���Ji��jW`fj��7�7W
��i���Q
�7%��Ͼ못�߸r�$��	)'�P��
/�]}�����߿}�U׿:SC<ϥ�Fy�nÝ�W[PT�=�}����9w}`n����&$x�vw�jse'���T�-J��UU��钜�|EN���Q�A6�Fu��GZ�;l�Χ%�M�ɺH_;&u�+������~z\�B��� wٲ����8}�u��76~���5�ԣr�#r*I%��Ԯ���󙫩��{��>�S@oص���8AG9�;�۫=�u�������@g.���a�f$��D��a�}_U웫���;���]W��Bd@(�	_ޯ��N���*����C�9%����v��%47�����l��_������I�Ҵ0[N7*6��:*|*mT�1�B<+v����ʵ�v���=nn��ƞ�b��rd<D��Ԯ���M@nl���7���vX�[���I�R�
Npf�jo7����I��Jh��w��3��F��iS�	�HRU�������SA�ff>Z���������۴���K�04�M=�y�����@g.�37n�>����d�\|�oiF�2F�*T���-J��T���O`bS@t�>�1�{41�/���fY��<HJJ����IXJCB|��Æ����!�: �r�|���J�����v]C����NH��C�q�x��۔qߖ��b7�T5	BR�!H0D�(EIٴ���@	J&�J⯋"�1A���s�Iy0�Lѽ&+ ���"\��U�UĒ@�y���������|UuW��Q�@j�l�)��ڥZ��W�q��`	='���*���nӶm��n;U��ݵ�q�uˑ����͓k�̚ݳ��ݷb�"=�u��2Y;���s�ك�鵸��Z�z��;�Ů���F�2�n���<`�-�w`��	�������C��k�1ɤ�PO4Y���ԉ�+2m���g��p @�:� c�zc��Nw0�k���}���൱2Mɷ&�yDgY�8ٷOs�<����
���Ú�k�]M�c��]���9s�lI�P{�\�c\�cL�Q'��p�GO�]�[;z�eѶܛO�v�M��x� �6��a8�l��v0,z��\q=Q��e]c����d�h�sq�]���b��xK����v5rd�y�|�	v��d�=�'5�ё�
ϵ���p�U[ںVWa���m0u"Ӳ����[[q��4�ҌuP��;*����[R�KU�Xl��V�ёs*ø;k��v�ػ�&��vNSu�T&����x�n8�6ƶ�J�����;v�!"zv�B�j����X�z���'9Ր�*�E@�Q�����Δ�l�<YM�����9rV�y�*�ڑ ڪ2�Ъ�\����-�؇��j::z���qٰN�Ol'g�G�l&�XF��<��Z�,�p��e�c�m��4��	�b���۳l�%��:9sn�+l��.*�v��E�7 2�S��j�Ifs`�i��݋e��)V�$��!*�ZlLn�5D<�R�U���n���/2�P$�Q������ں�
�2J�lꬠ݈��6��Z� ٖ�\RnA4��m��e�ݹ$�N������B�aL���6"N@[��'�ln�0�9�ny���K�q��Kkdl�u=�I������Ȑs���GF�2�P�#��(�/-��\gj`�\�=�z�:؜�3���eT���n]��lV6+#�KQV0�:-��n#�d�s�s5U/.�l�#��' ��ҝ<l���7M<����{���w=����'A�6�OT_LT0D�C�N�:pzC�}��z�ٴك���"pEژ&	�; �3����oz�������c�A�Ha�}/ng��˲Wds �덢w5��Uű���FNM��^77j�2Z7iά�JC�t:V���6��M��tF�z��I�Z��]z��6Ge8Gm�d��<�ݏ,p�τ��V۝-��2�B�V�\�`�v�v�mA�PQ 69�̜t��˧�s��7S:%�j�z�xBu�Y���(8r��*�}w�rt�9�qu�e�g�J������J��b+�E��׈H@���#�&���rGH�r�wv����I���9���_���˺��F���H�5)ʉ7*��d�\W�]��Ԯ�Y����y���3z ~���v�x��.��}]�R�f�js&�����\QG ��ª���jW`,�M@nl��7���TP�Ҙ%��f��n�Y���媻��~Y������p�5V��D�5>3�y�:�fL:��z�:
mju��l�[�vḇ���������(b�(�!IV{&��	�TP-J���p�]M@f�:n�v�1ˍ����ǩ/�}�ͪ�B��@BE4B����@� ϯ�����U�݀�*jse'�F�F�m�d��@��`wsw��ͺ�����=�up�͖w5���RH㩗y���>j�jj���T�{������8�������b�*Dܫ=�����1�j��]��j��3����P�ѹ���<{I�̼��#v�㬯le�a����+.�q[�������;�\��}���}���h�76~��o��!Ҹ��"ARjE`wu+�oy���j�jj��>�������[����!#*@���mՁ����ui;{�3 �;zD�����33y�;��"E)���A�y�nl������jWa���5u���0[_�K�n&�eIr� �j�f��Z�Xf�jse'�5�]����	�֗�8��e���8��Ίk���v�"Wn5;�DQ��g�X[�nu-kD����v٪����I�����5E�f�f�Q���s�wٷW��UP�)=��F��>Z�����hЛ��bR�*Dܫsg�ˀw�5XW�}Twsw��ͺ�;�kb��'M�����9��f|�\�r���M@��Zgg�5�a�#@���)�8���O=UK��oγ����ٙh�7�G)H:MH��n�wٷV{&����V�ۚ�B���Bp��ɷ���>LҼ��.1i�@7��Kq�؊������8��S�(qDT`)/�wٷV{&����Vw7y��:a�~�(iH�a�Ǚjj������0}�������f�X�^YZ��]�db��.Z�djz�]�o{���f�jse'�7�{I�)�7!	�����8sU5�����7��������;�(q�ܒJq�p�6���d�\�y�����8��V�HZ�(�NJHdE�<�Z�:	a=���l�p��ۦ娍@nC����׫DD�[�3��N��8��4�L&:���.�N�,%�ݱմ�q7t��e��v�맓v�c^�
�o�T���g]�6a�:^�4e�S=z�k&�
D���%h�����;e�U����u@W&Vӫ�c�:�I�uչ���u�kq��=\��2��d��:����`�Ԡ�E q����v��:q�ggv&i�jQ��D�6�qG��Xh��Ԝ̀��������djz�_����7����]u`w?k��7)��B��;皬��v٪����H�{���ꈉqȢ�R�i������8}�ug>�,�mՁ�<�`{�J�?�;�>�y����j>ͤXdjz�]��m����Hܔ���=�zp�����#S�$��f�j!��K����.n���^s.mֱ�u<.�at�#�P��yl�*�M����]�d��wg �j�>I+�>�T���y���H�F�Bg��"���v�Is��wk�� T �C�P4U�=��*��~��Uw�5_����W�:��r7��B��5u5���`}����J��<��pIJR�Mʰ�UG��-���6=�I]��j��/�8�e�B!�%؉�,�5=�q�͜����]M@nj�X��'0�,8�㻴�.���ƻ�<Yx�+�oSJ2�s��n6����LWRR4�S��r��MH��~����ͺ�33oJ���|�U��Է[H)q� ���>�T��ffw]\X������U_U#�i��AM)Q�%$)��]\Xdjz?kߍ�kif��� <{Ty��?������r�����Qq]ۺr�����*����������5SPs:K���u�1-�D��2�/@|�W`y��o�U5���`w�5X�����9M��e�{cgbB�5ն�M��l�����ϮKv�X.ya9$n9%(�'8}�u`ffޜ�y�������o�y�Lq����"Z���H�>����%v٪�����s��$=�7Tۊ�9g �j�>I+�>�T��E���TCK<$q	5"����������mՁ��]Wg��4	�D9�w��ʽ���~�BX��hwJ��}�$�U(��x��\�ĕ�kB�����'d��lK�Ƴ����й��$1���.�8����`6�.��7}����`}����+���`}�������W.G)���ݜ�y���n�8٪��[��}�����o3����f%����f^%�����M@-�H�;皬�M�NI�IJRRs��W�6j�j�����#S�W`,�d�(8��N�D��`nfޜ�W���3f��;{���U5 ��oy����~�EP
����~��y.1ڻ�R\V�;Tu�ƪ�w 7��y�'Z��g���{�=�I۲�7��`N�ɒ��ݻvܚ�u�=�:�Xk�-��kNj�C\�q����K�'%c�0�����&(C�W<���cz#e�um��''t𑫴���ӹ��0l�
6Ա�ygN�&�ujp/2h�܄�3����=��f#�z9��:�-2����\d�mʵV߻��P� ��Vr).㻶��r��7�l�b�n�n�u���Zq�D������y;4�����t��8u��`o�w��ͺ�����ͽ8�v����!D�ML� �%w��fgs5u5�uq`}��]W��կZI�J�)����m� �U"��#S�W`}�j���25$���X��� �j�7ۻ�_UW}�u`fa�[%wr)M�T��>���ĕ�f�jn�E��-�/}�zk��>q\��u��ۣ8'V�ͥ��{]���"]2����/�Y��5��x��$���5SPuR,�5=��m=i�#q�)JJNp�6�����uJ@QC2�E��)Mldz}QOU �.��|X�'�$�����w;H;�^H��w��iw���9.�,�5=\��mՁ��)���������}����+�>�T��fa�.�,�ߪ۩I��H$Ԋ��n�8��6j�k�����#S��y��@�hn	�)�ᝂ^#e�B��9�y��N]9��V����3�l�Ef��#���3��j�jn�E��F���z�;{���O��E1J�G��X��� �j�7ۻ��f�X�j5�ĥ܉�qƙ����#S�Wg�{��>�fj��7�x�G����Y��f��6g{oT8�ѱ�	�Ԝ�k$�$7�8질bh��Uv�̵��##���p�F�ִh�n٭�`c��#LV����q�։��r���c䙫$�Ff83\֫4d�6,s{�s4fw�tg4'd��\����VK���gh�7ey����4�Af�msZ�8�Z�j(�!q�7y��RTT�(���zNXdN�v��rr;�9uk]�M&�60�b��P���'
�	���P��'!��E�4��E�!6I������8�:Tx�&�ShqO�j|!��:� �T�Ta`t��!���ڨ� tz��@�.��n�o����h7�"�9�A������vj�jn�E��F��3���ؤ�7$����� �n����(�>���ĕ�#t��<�5������۶f��NN��p[fzИ�lx��c_1TPq�Q�TI�V�m�`fF��$���ؕ5f�;�f"`���g��,�����7����7���[��g�3Rj�ig�d��&G�y��$�����j�X���{Mz�N��)"��s�W�]��Ձ�{�>���5�����D���!��^�N�W�ڡ�>���ު����1QL��G��X��Ӏ{�5X5+�>ĩ�foynҖ�nb�xz��:��u�ml]mpH\�ɒ�l�S�u�E�nn�W_W�KB�ZR�D�����3�jW`}�SPuR,�>�x�*IC����7ۻ�U�}�u`nfޜ�ٮ�UU$o�~��E$��$���n���Y�����(�w�<34�81ʉ7*��WԿj���݅�@,I]�y�����>��k�RG���t���ٮ��n��K���1%���|�%���U@�����i��(��5}�"�5�g�^^[�=w=��e6��m�r�9�Wql`Ӷ㱷#hn�[��A8���=!t��s���{��cG��wn7RBn��,����1Ló:x��-&{d�Fս�m�C��-k�UدXD���[�����	9�����r�iY@g���c6S�v� �Zz�w+vɹ�\-����8�ؠv���G&,֭oxk{ֵl�����P�/,����Y�G!{<b�c���t�ʭ��:<���kv�]��.�����������������>ĩ�������pś��������&9REO�� �i���>j�bJ���fo3��P;�L<đĵں��1�TQ�����R�3{���u<<ͼD���DLô�U����Q@,�W`}�SP��Ӏj�=Cd�n	�Tdq�����{�J��_j�X��(��1��sͺ�=G�/c%q{b�G7oJ�D9eb�e���!#&�Z�Z������J��[��`c樠-W`o�nԎ����D��`n{oNo�w��9!��h	�a�(�1+RDځ�����}ߚ�^{����۫��S�JI"q�܎������(�-Wc{�������v�II2B8����K�~��������y��Ԣ��N�<;�<-3.�癛�3uSP�{ܷ����]�`o�7� �b��ph��}H���[b�hڅzrsb�Z��6F8���ͯZ��E4�D��br��=�� ���`o�w�U� �f�X��mI�ܸӦ�g��,�R�b�vn�j}��«���f�d�n	�B%#�7ٛ�Uw�p���CI0Mg��oN廮��f�{)I$nG%9I9��fo�U5 �U"���TPw���������~'��$�F9Q&�X�����o6B]j���M@b7G"�sv����_v.�A�5���}e猥�2�/U�Y\����羝��AsN��ʢ���TP5+�>�T��T�7v��Bd�q	G`o�w�>����ꦠj�X>��7���N~�xg�������M��SP5R,�33Ϲ���f�8p�ڴ*)�*%$)*���5]�Ϻ��Y�]�flff��!F9���j�3I���iv�L�-iL�4ά�ٽ�!ʧhS�A< �o��Õ}�0_�N'.�'I��F�� w3e�W�y�jU`}�����7��y�"F��ٵ��ۯeS���O}o�s��ss\.�$�k5��j8����j��|�?�����`nj��j�35��Q@^�Q
)I$nG%9I9��ͺ�7ٷ� �Z������3~{��oG<D4D0C<xxif���76$
߳n�媚�_f��JI"q�܎����j��`s}����uaFw�zp�m�(L��
A�31@Z�W`%���߳iu�(-���LtDA0$L�۸-T��'(r�ET�Hj�E
8�]�vN�ݣmnf����b��uqu��`�ȝ\��m�Q��C]�5��-�/]��tqt�7)c�!��[jͩІ8lg�3[C�磍aے05�ǁ4niѷ��ۥ�6���^��;p��wmM�m+��l��X��=L��A���ך��]�'kV�b��p�����I1�SS1B]�ͤ�ggX�=���ߝ��{ۯ������]��ս[Ox$	�s�!�278Ŵ�;M͓��#Rp�U�[��#��D�X��73iu�(�n�w
ͱ%E4�(7*��{-u�(X��	j��fffa�s[��b��j%�&a��*���Ek�9��;�.���,Q�� ���&%�%�f(9�����v�]�ܺ���ͽ8��v��k�JI#r9)�79��M@oٴ�:���v��\7M�۫��b݁�i�h�ˋM�,�u�G���Xh�����}̭]���"Z�߳iεEk5]�������])$��Sn:�r�չ��v�E�������몽���p�����I(P��
A�H�Y��͔Q�o3y�f������@^�TIҒ' �Lrs�}���X�e��:�5��f�w
ͱ)� ��vw�(�6�`w�����ˢ���w8{&�꯳@���J�pm:r��v�\�Xstz�5k�+�ɓU�d�wf�z��VQ�ʋ�KM\�j�wg@��������8{&�{�zp����d�����]�b���]��{�͔P���幮��v����HێJ��p�MX��{��j����FG�Ө+��-�C z ؠzv���oy�z���ڮ�X��4LDL���-#��A�ffg[���1�tP�+�3�4�7��l�'$�1�E9g �Q@s337���f�ݫ���‽ͭ8s!�))$���9HEJ�(�i{=BqlWfު;:��Ny�O/7�y�3v2�u�FRdw&f(��v��(��G��7���v<b�Q'JH��1����M]�3��%\X���j��{��w=�o���R%QҤ���ݿ� ��QA�o1y�����M@g��M/n�Or�q�ӻ8W�]��{7��ͺ����B�@��@v����~ݾ��JB8Ԁ�Q�`^f��35SP}�H�>|J(�LB?����qlp� �#[=[k��v�nD�.�g�x�R�du�.�q���3e�n�,������تm8ےQNT��;��Ӏu{u���y�=�_�os�8䑉Ĺ/7E���Q@^bWgy�uOؕ�8��!$D�qr;˹�����j�ݤXw����#{���	��$�I�C�99�=�۫�̽8sϾ�*��=��������Gh@z�Д����𦿌�E����w�2�w$��Du���<�r	��\,�7�8hO�n�؝Ƽ5kX��|.��M^xiN p5�TI-���Y�)�(�;�/\�a|su�i㡭(쐳����Œ�����N��׾p����.ø���=��\�̪.�Ax؃��]��+ǚjT`�.����Z󇐫���tnLe��0M�H1��:v!�Bv�u�֌M�:�xi�5�*�y�ߘ������ �J9��vA�F�\�:!��C�s�t�n�6[m�E�ڠ���ev�V�S���@��`�˸�,� �kcȽ;tl<q��ծ,�q�2�q��pmM�r��ݹ.=�{
�c=Yѷ\�m��;�m��̛ ]����ʉc�ygH��ў��<�A:ݷv�T���+�y�ri}Rm\��Nn���͞5t���	��.(퓱d��:������ �˵ط��q�/�q�V�7;���'e��!Cs;�p]�
8�]��4�!y�;��'����!�����h9;m����і=n�l4�q�m��%����a,y���4f���{*�5��Η��n�ٺ��[s۲��@�8v���j��y���8�u��<״71��Q���-��J��<i��)WC;:n6T�*��[��Mayb^3�815KJ\�n�O��Wlk��m�2��<�^�b윷9����=V��PjYn
V��Ԗ٪��k��wm!;�H����83�n�;���یΉ ��jb�{n�m�mƩ]B����;�8�Bl]M�0���Q�@@��W"v�LfBjs�8K] ���v��=�x���mn1[����zj]��:J\��f��kG���Xʶ�v֧*�"�S��7B&�]��q]����ix0������-8L�v�]���&�Ӛ8�dCb���eej���ٕ��q7^�.΍��Pt���kpӆv�6�-�I�ۀB]pp�][����[1��Z�TRKs�m��M��Z�4��x *�y�����@QÙ z���iӵ:�U���Tʲ��tԍ�蚫I�2S���fM�W��W[c��݋��u�`fwez��s�¡��A��ʣ:0>�X6����k\n�]@��no�C͕�S3�j��dj�����˳�qAv{DE58f�������OA�m��j�Yk{rX�瀥If��:�MHk�$lR�c2W))Pb���fЮڪ�:c ۶�å��r�,�gu�ӈ�*�[ݚ�����{��{<KJ �m�*�Р@~����� ��]z �!�")��T}��:GB��	����睝�c񓪧W ���tvG*��	
��p0�W$.�n�����sY��;��+���]�\0b��nz��-����&Z�q�{hv��ݨ	� ��>M�����]���g�n���Wu��&@���Ncn�۱.�����E�.̕�P�*Q2�+#҅�r\Ye�Us��F��aԝa�m������.�{m�.g�Hn�������ݟ2:Y�w{������}���k�[��s�'N�%��OmnSĆ#3�-�%��@5�w�m�6:y��e� ��H�>|J(�����n���3�_�Įӷ)��;��u{u�����T���H�7#]3��LLLK����j�3U5��%\XY��7����NIrIR1���j��/��E���Q@��j�f�&x��m�A��̽8������ߢ��uu��(�9���Zs��ZbOd��qx��۶hmk�F��:��ҙuI\v�]��M�\�{�d���S�fZ���$�W{����W`fl������%\X�z#�w�W,wiIw1%��ݠPmS{���f�4�f�(ĩωE0���i:Q���Np{&�;�zp�n���o8|Vm�AMGQӳ��P�m"���(�-f��=���U`{�1%v��NH�F�����`w��]��n���7��E��Bp�+��=]�l��;�z ���.��Rsu�y+v�:��[�p����;{�޴�*��k5]�����߳i�y�p���7�����9$m�%H��8��u`g}��djz�j���n2vL��-.�q�rB���/N�y����+�ܾALHh]*�C�h�{��8��Ks�딩�䑉��)�,9��es�v���(9�o3:���p����"�"B9JB)"�9��偋e�m"�܄����)���3���ٶTN#a��^xu�6�[a�ɪ��cu��[�������3�9��0b�E��H�7!'�7�����3�?X��pPtp�3��ӟ���7c���{��Ų�>�YԖ�R�Q-3�1TX����+����w�S�����=[B��RS�0�R+�%v-�P�����{ޡ���K7���S���yɼV;[K7�䑷$�#"&�[(�7�O`nBO@Z�W`v�a�z�duJ%T�t�J'W;�L]9^�t�]ٝX���׈x�w��b��0�2P�m"�܄������Ų�sۭ�G$�m�QNY�3�uX�U��Q@oٴ��y��w��%!$�RE`w�o�pnM,�_}�y�f���[�@^!B��&	�q�h"f�[(�7��E��	=3?ݫ���i�� ���������^�qJ(Y��[(���S3^�D��7]"匕�x�աK�BS=�����{�v4�L�ڲ�V�S�ݲ7l���Ŏ���;2�{qׄ@��y���K��͜_��o��=�P͠�<Ea���,q �-���r+����]&�u�E�ڒvp�h-�[�ï���E��Yy�B��:�K- hث���m��w>t�S.�5d�i4s�tF]n��eF�i;`�7P�=w��w������7�ٺ�I�[�����p���`��5e��e9��;)�rnnb�u�������ԝ/�o�9)‵���Ų�o�f�,�KhR9*JrF�����7��ۓK;�8{f��W���[��䑶�1D݁���~ͤX�(I��[��������n6�RB��}�� ��`w���Y�4�3}���Q�$�m�QNY�;�uX���fd���}�� ���R�����RB�N|�[<m[t��-��:<��������-�ur�ٲ8�RTR�.�~����4�=�T�������?G@�ĸ�3��}uW����`9?0����%-D���h|�;:���9��]����U��o8kض� �G�E'"�=�m"�̄��ffgoy�9u������g-X�\�j4���=�`w��� ���9�m��3�IH�)�I��z�U��6d$��*E��	+s0�E��F��IP�O�i4�%t��p\YK��Y�r�Ipr��n%�]ɞ+�L��Ti�9�=纬{�zpy����p�b�V�����F�9�m�g�3!'�>�u]��	=�x����Iێ
r����`w�����UQ�	�(�����ߺ���ʹ���pܚ�d�AH��>�����vd$��*E���E�k�P��Q$JMI��=�`{��Ӏy{u�����C��|9��G\�`�Vٵ�]�W�#��8��b��s�]w��R)cQ�����X����^�v{�����V��kK��WW)����<���)#�ݻ�{���ra`��ID�9RH���;��� ̄���1R,�I��Y�3��LC�̴���݁�����`fBO@��^A �K���ԗ�<�I�r�N�Ix����R,�I���W`f)E��^��aI���&����I9����ݻBq��wcuM�R�i��狤Z�EF��`���n�2z�U��Q��{�3����ퟣ��"BH)9���U��Q@gةd$�|�B���(r%&�� ��i`{��Ӏ{�uX���v��lb
��D�Rr=3>���`n�s�|��2z7�ֳ��)܃q*Mݜ�{���wU�������s��i��b]Q��1��5m�� Y��ǯOm���R��M�f�ݔ��Lp�`�8����wW�Ҟ9;i�K�:�]�@���n�s�8��E�h����v��a��u=s��KR�WX8�6�&�����m˜�:��<.�a";n4�S �`XI�W=��2��i-�hu�ueH����-(��Vkxm��e�։A��U�����lB��{X��{�}�ǽ�����;֭��E/lr�/�7�w|�ܽ[��͸3��t���Z�.���Qy��6Y���/�λ2z�#�����z�9�|܊7��M9��=�`s��Ӏ{�uX�y���$~�������LD��oW>%s7���������X��d�n9"�ێ%9g ���>�5]��	=b�X	l���f^^^fG����>�5]��ͻ�Ł��_����`{+jh�)IG��E:R����0U���7'e��y#I$ZrN2u��jN뱤�)C�)5'8��K��ޜ�ۮ��sw����t�J�n4��ʼ�Ϲ�ք�aHP]���4�A�����I]�����7����]|�ː�%M���f?ߕ���o8��K��ޜ ��ͦ�n�%I71/A��7�1.�������T�2V0�[����$�Ns�{�4�>�"��֨�>����(cW3��3�LpRZNx|'<�]=�q;��@Gh-X�v�6�/�9�bi���*1���ͷ���Ł�Q@}�j�r5=�#b3M��u��s]���o8y���ޜ}�\��(�r% �����ߺ�|׿g.O�)Z$e �X��+_|dW�{kz>����Нl�gE�q���0͞�JFX��fY��1cc���[� ��H��l�KE��V�d4�e�5DX�M�Ś�]禗!��g{4E�adgk��Y�E��f�Nζ�e���V��7���
�3��&���+0�,��)"e,1���n"I��6�5�q�bt����T�����,�s5c2�7Zַ2�XYYae���	M��ٔB� ���̬a1�L0��fb�L#6w�n�� �Ăf"'%�̳
�X��1����3)���.�Kx]��a��h;� ��\ȋ�d��3�9�dl�N��e������Z��f���d�)^k�c`a�Z!�6��A�0�g;����#;6dT���0H�	�N�@�z�{E�D���dW�� N��*z����)�}Ta��ѥ}2}��jK���bK��k֒t�J����<�U��{oNչ���s7����鲕�4�3�����εE�۪��������h[_��JD��TTb�!���ծ֞F8�h�YM��t���ҭ����ç[�q�ӻ:�����ټ�皿UWw��� �3Sm7NT�F)��٪��[���7�� �j�Ѯ/�8�nI%(�s�<�U���oN wse���7�ެU��I�q��z�3?ٽ|Xr�>�5]��0��ݑ!���bH��������g(�~��6���N?�9g ;����U�f���l.z3"����2����+&�F���8��ýLp�"�z�����n6Q�2�s��{$��I]������H����7��;��NPӦԜ�皯�$fg��p.]�$�����;��OK��LD����/@}��Ł�QG{�o;�%�`-{�X������v8�cwg ��ؠ>�u]������R,ٚ�"!��R ���y�3�5X���W{��Vh>1%*B(
B0� �)���L�g�����~ϋ�Z;=��K�;n�W5!����˲m�xI�cZ�.9�<X�-�;]�k��g�2K�-��NF�N��\�Y"�0�]yv�H��W�ܶM��w9ӵ<m���7��Y���ڦ%��7��vM�,�=�G�E�	�m��'P)�#�����
ܭ.&]6'���z}�B�9%ڷwm-��`��\>��yg.x���yx���wz�_#��+�����vyɵ�ɫmp�F��6� g�ݞw�Ե�0�����gl�s��*E�|�M��U����)"MFB7���oNչ���w7�<�U��ܡl����N6�����֨�>�j�r5=�b�X�6H�qEu*A9#��>�����v�[����H�>u�(9��t;�3��4�'x����罷� ���`w�����x���#j�����e&Q.��ĸI�M�q!����t 7;�] ������4�Rr+��ޜ ����$�������l.z{PC�]LH�$Loy��s�U]����;�<��Ǿ�8y��ٚ��kٴ�M�� L����J����w���zW=�{���;�[����$�Ns��ﾦfu���ޕ�`-S@gڕ�6iZ����!���f� wse����8y��2�֝9Q���#�z����m�MʝNض2W�L�h�y��z�R����tӌ.� ;����sv������kp��\�rꙙy�yyw���&f(�%w��{�gql.zw�.չ��}�F�?4�4�M�r��6�݀�=��S��݌����o7����f�z��TP	o+�>m�S;$<83���w����K�����@g�+�3�5X�`5�8�أ�$�Z�:�|��r5=��S�$� s�r�]�	p�Y�\s�b�F!�YѬ��Jݍ��x�u�,�n+��Ӫ%4|��_5E��S�:���[�����$�Ns�g�j��RFg鿕�g.�>I]󹍨i�y�ra�%�y�zw�s��T��J������Xyh��a��a�����3{��˦����7#S�����S3	�ᙛ텊B@������LH68oL&jC@``�*S*�}_Q��s��{2mIqEu*A�&h�%v�jz1N��>u�(M�6��Zi-s�tKbS�l1����u�7i�l=�*�&[lf�V���.���3v�jz1N�����3�����J��M4�����f��Q@g�+�5�TP�B4�̏T<�˻�M=��Q@g�+���y�����`f~��p�ᕴ�m��"DjG`g�+�5�TP�u=�3>G.��9��&���$�Ns�b�k�?UU{?^�|Iu���ėy��It�Q�j���d%V��Y�Ͽj̳�oXouQ��"�<��kwN�v�;`���)Eb���S=<H<0��6��Rl�w,jq�g���nvv��_���g�.�[�c��h��f��F�z�=XC�{'���#S��up��f�����jT9Pv���
�Fi�n�5�etMr��zr�amOw�<�\���N�m�&㓇��n��*�isF�WM$��׬��ۋt�*�on��~�~�N6�[z�������7�x.��U�5$��![�[���<T�N�T�!919Pm��3����[��w7y�1{5����rBb�d&���֨��7�����vt������=��q�QĝJ�NH��R�_uE�)��Β��'x֒mJ�(��jNpY���fj�[��w7y�;�լe*"q4�S�b���{�IE�jW`k�����,�qw��6�p��:�`��5e�i�.�X��x����7*u�u���q4�M=�󤢀ϵ+�5�TPb�O`{Օ��m��"DjG`{���eN�f7��z��NS3T�{�IEw���~��jF�rJQ4�8�����f�ջ���sw����V�`��-$<LPb�O`|�(�3�J�;����v�+S��)��N@��\�uE�jW`k>�:���7��Θ[w����� �붽���q���'��;[ɡ��]��RV�3���f������V"fb��Wu���(�gS���'�9�Ԟ���R��6�� =�pw'�p��v�����)Q�������r���~��U�}�����ʆ�_���;����5��xVйi˥"e�z�{�IE�jW`k�0����\ �3C�&�r2H����n݁�o(K����\�Β�a�B���8^���`�rrԇ`�.,�׈t�8���]G�˹�+Oj�Q�? ��Q@}�:����Q@gڕ�6"u�H��r����f�ջ��ϵ+�5�TW{��w1k'�:��&&.��~��R�_uE�l�\�ͦ�4�&�R	�����8��k�w�����j��(eJ�,%Pzz�~ى-����ѷݢPӦԜ��5�����:�u��n��O\N8�RAJ)�M� C+l��b�zrs�����l��n)�\y���㶒6�
rG`w�3W ���`{����u�����V	m~��ӗII��\�IE�jW`k>�:��=���m9#�ƈԎ��sw�f��ٚ�V���-�SR�$���� ��Q@}�u=�󤢀ϵ+�>l�$&)"#MʄR;�ٚ�V����n����$�-ڡ��B��Lb��*p@�̌L���Hs(��0��*!��)R�����5���Q,O�8&�8�	R�9W%S=����R��u����kgiبHb��q�ui\SWEDV_�R �,Es�]ܤ�|�㔬�(S����^h4N�8��Ul�M�IR�[J���*Fu�j3F!!ZI��uߙ��r�)�2��F���LB��	�����ۤ�6j���F�I|�q�T� g�;�:�t6'B]���14��B��
D�5�z�E�*�j�TQpR`X6<���@U1G]�Sњ4d�4�����
j�*F*�8������Jm1�D% �ؕ���y�C˩UV�o��(&q��F����E���"[��J�%�XV����nZ&���}�_;'/gR�Z�"G:6�~B���D�c��7��>LE���BjT� h|^D1�1�_!ZQ+Z""	� 'G�9$�6����@q1pA� 2��,2FU�
(���. �e7%�H9CӘĹ��j�h&S1rD�șdٌEUt���=���rI#�I#n0�U#rl�*�W�h+�=w1L�{t�.5��� ��W�Z;g�\ǖA6;Z�$�@�A"Gb��ZuX+���oCO�p[���k-����T��X�y�M��鐮9�A$��q�P�lc������ܢ�ī�s��Ol[�Q���3��}��˄;��&�	�/`n�V�[�T�=q�v��6I��jR�p��Q5�`n;���w=F�ݜ{7nss�����>�Ln.Sgs� ��{��(8��]�ݱ�]��M=��M�qդc9� v�bmQ�����8j�݊��	�w��`����0��u=�;<7�]Si��@c:�pb��`@9P��I/[�BI�]$g������:�غ;�=N�.�
���Jn���{2DX��ʀpD��� T���j�W��}J�Kn(,Em���럕���R�抽�)4����X8UR���Z���h��z�9�U�DǱv�bk�.��k�`��솜��i&3ny�Ԭ�5s����7�):������b��Y�<� ���3tfv�|�)r	Ä�4s�=��9�z�N��.����t*�n�P�v�ˇ�m�qOm�=����5Ȇ�M�6�c������cY���a�0\c��f l�m��jcv�:�r��`N)S��Ch�媀�l�6�6�E��n�:W��s	l��e��"3�a�:%�:B�V�	�WI5 ����"��Mj�Xζ#����
y$h�q�I	�[��V�R��]�U*��PTl��lVpiӵ:�aV�Qэ��A/&�t2GmKU@U��Xt�a�a陱�[s(Z�d��r�P���-: ��v�m]�Y�<q:�lm��V� �ݵ���F�um�co����T�n5K����!���F��EP���iU!���8��N�..ux�=�I+�Œ�"# V:��V�Ʊ�!"2U9����pplJ�5UA'\ m��k]d���کU�=F�kn�7�z�����of��g��� 
����6D> 
��?�"|���=U�C�%��A��s� q�]�\�֬�٬����V.w&�`��Q�q��w/q�]�1nb@��۰vհv�s%��Q�r��u>���f��;n#X|����7��8����8��H	�c��k��2��9�\5۹�;,q�@���/]��nM̻a���m��;5�����mԔ�m�z����z ԇ--� )�<"FS�c��[s��e �'k\!�b.���]�זּ�2Ms�N▭K�#�r�Uʪ*��1E6��6��������,��nӝ��y�:��1rY"��q��p�.�װ�&�#�{���}���ϵ+�5�TPb�O`njh�yw��*A9#�=��� ���`w�3W ����E}T�����d���8y����>�:���7���tP����V�R��6�
nG`w�3W �εE�jW`y�_5E�6�Ɉ�n]5$bW-p��v����ށ�7�;홫�j37��$萕t� �d�}]��sOOf��]Z�[l:��i�`ظv��Dӕ##�#������]��l�\�s]���%�j�ABI#�'�����ߵ����:,��D߆ �	��gM��	�(�3��3y���8�x�
&�A����o��:�5����g�j�;��OD�9!9)˵����r�7;���������.{sSn��$%H'$v����皬{fj�[��׷5��O�J��מ�bɪ�N5qs���W$�A�ݰM�gn�ԜM4�m&I)JM:mI��y���S���j�f����<3�*D�AIȬ{fj�ꪯ��/�����v�jz�3{���h����&&]��i���3�ؼ��{���Sy��~j{{�������]�ĴL<�D���J�������+��9o�`s�Ioڢ�R&�"��p��V7��w�s��t��J��bNDɮ�fQ�l������q[\C�ڎ s0�cqgX���$ӈgY���:���>I]��z��Ų�t�`�T�.� 73e����3��vlw=��S���"*�%� ��"bfh�%v�I��:������I�I8��)4�'8�睊~��zw�s��SA^f�3h���3�X�%4��P�N"�U��)���n���}$�Į�IC�/@f)�� �T��J����N�����s:5t]/N��s�����ӭ�����zP4�9�n�ꀞ�.��/�fh���>I]��J(�:��=��xx����H��>I]���ޞ,��. nf�����)D�D�^&��Q@f)��w����r]4��߹�;YLݡ�$B��A��ٚ� �T��J��Q@}���\�g��ȩN]� nf����pܚX�{���.Ui�@4P�}?'-�K����n����t�y�ǎ��=<�2+����0��q���z�A��h*��9�Ӻ�;lp�%�`��۴�v�\̒s)�xw3�N1��c ����1u��p6�Wh۬W/�˧D�S�x�ά�D�:Uu2d�A�<fM���;] QP���<d�k�ֲ��m��4�j�;�+=tF4��\6���#Y�-�@��P����k��N��w��q�m��̧h��wZc�f 8ڭ�a�z�R�=+9�Yuՙ���;�9]���(�:���4w��֒rH9J'M�9�7^j���3zW=�w.�>I]����O��Lđ��3/@n��{ KT��J�ך�Wk�����w-8��k���%ܺh��(������s�����M�N4������8��V�L����`mx�=q�PD�'�^M�`y�Y5v�:5Ά��D×�u�η��u-m	�R
�"���� �ݺ�72f� nn�{������В�!D�%���U���߳�3jx*;UE_k��7ۻ���K��3T��I(p����%4�%vsyߒ�(JW? �f�m]8��R9%����p̚X�3W 7۲�����I&���yxh���n�(�7�*\� v�M���p�V7�9R2�c�)Jl���3�rq���X�7)Ć.6�����* wL�D��'s&j��vX�J���f�Ò�(��t�õ�EQ4�M=�,Jh�J��(���~ t���4۔�2PBI,���}���AЉ�	
<�����jEG?~��Ԓ���^$��	��v�
��Ɯ� �ɥ���5p}�,9�������Ms�0<�L<L��Χ��Mi%vݔP�cH�mֻCdLu��n�1����4ܩ�����C�lIiR��iw#�4ۨ��!���bS@^���[��ffkp[�`{3i���C�jT��I`s?n��s��(����n��gw!�%��N�Rs�nd���?j��d�9������R�G�
������fu��� �)�/y+���7�����Ia i�E�����(;T��V$�é?����3��[��Mz��n�(���6��w�:�͞2��C�eq�Q���.��v����8=�o.�C]n8���i�mjfl�w]��e�bz ߷f���BϵE ��(�i�p̚X��V�̖3wy��$z��~m5�Q8�<̽ �7��7�٠/y+�Ƨ�;��5Jn��)I�Gˋ���`sww�q����2g�`{3i�lqJo-2D�L��+�F��3#����IxA]TPb��G����K��]�Y4��*v�Ư9�;�'<D�v�ˇX��2lG���2g���W�ѳ�]����:��n���o�_rY����κZ]��.�/.$�
�N[�.۶x׍ںwFɬ����ҭ��#:���	vhٝE��1�+L�l��dzY@ۄV���uԲ���h�ynM�:B�n4j�ܰv��_g2sש�:��X5d��r+�w,�� ���
�UU-8��ܶ9��k˶�،� 1�#ە)/'����JF���nsu���H�2)tk<e��ͷt$�}��7�٠/V��1�:P�R�G�'����3��`sۊ��(�3�!��*i�b �������Z��Y���1= X�ϛM6ԂnPB9,{sy�7�4�9��~y���T���燙��y��y��l����O@�l��U���ҏ�s/i����l	�c�<7+��cRI�DVEQ��/0�99��*�N!��8W�@s��7�vw���1�M)"Q>\\ �f�ڪ��4����G��@�ν��s&�<���UU}�G�6�v��d�0D�L�r]v͔P���~̖wƷ[mJ����� �d����O@�l�w���o.������q�8�	���?j�w2X���{ri`��6=�GRB�m)I�>�Xm&t��A��.Z�+�;�d��Ch�l=P����h-����9��� �����?j��Y��mH&�#���Z��Ų��1= g۳C�!�}��D�D�Rs�{ri`s�Yݯ��Q��Ѱ��6w��� ��ę�	��n��&(;�<�A��a�Y��$Af�E��g݃,�v��QY2�u�O<̲�1C�蹵�&��y��� �# ���gT��kt���:�07t:F�[��b�&dQn2��(j�&K���� ͦɈ+[ܜ@�|��tu��Eއ�,��8�<N�pD��<Á@L0p��+|{}<�l�Y�`�-"WY�]��&)����s���7��ή��ͰB�J����c�z@H�N���c���4�C$z��p=4i��M4�6�֐"��(()
V��i�!�2��u�{<L�(qS�N*y��f@J�͘�kU1��10:�N�A�@��A�G��x���<�(T}D	�SC�B�J�x�=���B��T�x(�����|��~��0�M��Q8�Ӑ�9�ڬ�̔��v�7��ʸ�>�d�só�˼�K�Խ�n%4��v-�P����`V7�$1��rF|���G
pܜ����ɳ��g��Z��c*8��q�,{sy�=�4�7�0�U��W��`f���"mJ����� Ų�|�J Ϸf��Z����w5�;��q�����$�;:Q@������[(�3�&��I�&^�K �JhŪ�[(�;�x~J������:FiM
�`(!v�Mк%0Oqw�B	#� �V&��UB�T�λ�ʯ#�Ǵ�nHڐ7%������ɥ��م�{�����3F�|D�TI*s�^��9��\R�5�ْ�E��舣���A܊I�R
�"�Ƥ�@��?�f�n�7��%�`kjn������a�d�x�(�Ε�fgp�Jh�u��i`s}Z��rAJ"�v��͖w3y�;�4�9縬����R$�ļ<�31A��7���w�r�(�X�.����֨�I�D��i�p��j�� _۳@}�U���7�{������~ѓ���.������o}���Z���ԩC';��m/N]F�=�fM��ƨ.�dso=ϩ���ݼ��Ju[�x�lT=�O��N�%Zq����.�p!������ma��M�&w�2\.�t�=؆6g�۞�*�v]�欦n�X�*^L̆ ͜;ź7P�b�KGTp�N��V9��'�����BT±�^4td�U�{��w�����xo�?�6����n-�v��[fף5���c�λG[ �[���S�k)��̄G��[@_����f��~j�Ϝ3�SP���;]T�PL�T��橠>Ū���j��w������IʊR�rK��s�wri`s�w�,�n8�%!#�I���E{^�3�٠>Ū��5��"#NB4�,c�V��%��no8w&�<{JOaM8��:k�IH���69�ŕ���s���>���sV��H��C�j��&��� g�e����p�M,y�+=��5"N6FD8�W{��u���R@!C�؈��"�h�/!k�}�4-Ӣ����Jn��ށ��?<��{��`ws7���v�)8$�Bp�9��>͚庮��l����@�z��%�D"�{6X��� ������?}�e{.�����Ƣ*tx^2>����5ں��u�Y���qL��㋆;��I��E)J9'@��?�ܚXǸ���K��-�[�%IHH�Rr��l�����@�l�b�v͚�Vģ�F��i�XǸ���K=���� `�F�G�3�ү����`}�<P�G�O.�32�4I*q��s6X���w2i`w�3��n�R$�uԒX���~��ī�rz �͚��4L�����0��N+nɪ�N5�:�Wn��$m����n�B��FF�F�')Jn��� �dҀ�ak��l�bJ���gP��	?��,��V�{%��n�8s&�+���W���h.E��l�;��� �d���=�`+=Ym9QJR�H�;��� �i`w���0y<D�/�Y�{��Wy~��RR8Ӝ���,���~O`����9+�9���5s�ĎKL<=�Q�^ʻ�a���:F�ch�U�:��gP�ڷ�`��#[�m�?O����ٳ@}�����<P�t����#Q58�p�͖}�����,��W�������n�R%"r%ےP��vإsy��G'��S@n���NS��9��l���=�`�X���w��k���!�J�� }�l�bJ��J(~|�
J� �g��޷���LӬ��; �ݪnp�m����I�3�qN����^�n��ڴW�u���庶�����nJ����&�d���Y4����]_�;��E��cX�>c�GN]G]X�n�j��ݮ2�:^N��1xZ��]��>]ҥ;n��L��.�5<�9Z[c4��li(�uI�	U�/�Ol�ct;9%��F�;g���u�a�n�g5f�Yo7��e�V���(iS��|i'�G3� ��3��%m����w^�Ƚ�s;�iݭy��[��9�;V�c����YM�e�.S@f$������Bנ+=O�r�(�G%��n�8}�K���w��`w|��kqĔ�5"����R��-z?����4�.����%t�q�Gr5�+ ｒ���7���K=���9�#y�y����S@f-W`}�Q@Z��`~���z
D)R)R"|�?�H�D�`��4��[�ֲ�H@�Mư�^�n<�-%�F7$�3��� �l����`��X���R5���I�p��.�H�:R���IY_�LB�����������y���z Ż4gj�����R$pI���`s^���,{sy�;�4�;]VVЫ���h.E�>|�b�vٲ��-z ����NQ%�H�=��� �i`s^�8��v����RA%۔T�ݗ��&��p�k�@�2D�1�u��Jֱ�HԂR8Ԋ)9�;�X׸�.���no8k۠+��(�di�(P���͚1j���E����R�IRN;\ �e��no8mTq�A����!��$�qCRH� *�(b�0��� ��R"Z�*$��" ��0d��!� �p�C��
@�D�G�����;�uX�e;�7�R�i�,yj���Ej� _ٳ@f����jFJi��8}�K���s��@f-W`w��I���1�h��ihgm�
��rq������s�Nv�v���1tb��zN�c)5"!8p��X;����R\��\�<|6��̻r4�����4b�v٪���^�=`��(p%q�`{ۛ��f�X׸�.����%�ljA)i�����3>j�j��‷�6(%�������J��QJ�w�5%��|�xGr�Dq��X��,.����o8}�u`{�Q�bnQ!RR�'PiB��l����c.�\�;QM��n� ��8|�L'��s��^�v{����m�ﾯ��;���`nn��j9J0nG`}�j��w3WSP�<P��4���G���4IR�i9����V{�K �}���ww� �y,ѤRjIQ?���y��f|ή(��4�rW`}������em%���6�W wٲ�����;�0]- ]��@���Mݛ�~oy��Us� QW����#���M�9���Py((k��ED$�������QUk�w�����_��_���������|��������������?������o���������U������fw�o�z�EU�_�t(�
P
��g�~#�����������t�x(������i��o�N������<xW�_�>��������G�����[z�@T�D�JUBI!D�TIQ!%D�HI$%D�TIeD�Q$!D� �I�IXQ$FTHP�BHTHQ IQ %D�Q aD�THD�RP �� HYQ$VTHUeD�	 BH%D�eD�THQ$!D� ��BHaD�I%D��HTH!D�$IQ%aD� �%D�HA!D�VTI@BITIQ$E!D�A�YQ!PeD�Q!P�QI!�TIeD�BHQ!D�Q%TI �!D�!D�%D� �!D�%D�HQ$E�		F d%BP !T�� ����FT	$$	Y	e�B$$��B��HId$��	��		`&B��&@�)
A�)����B@�!!BB ��$ ` d
���$ Hdd!	BRBFBB �Bd"H		IBP`E$%@$!U$ `EI$%I	HFQ!��!)	�"�	���)bP�B��X@	HBE	 $VR@���@�B � !	D!%F �BT�VYB$$	 �!�(!����%	��!
�(B` %	�B@�P�!��B@��P$ B@��	D�!BU�$@�!��B ��a�!	E	UITVP�BUdAE�!	��	��%�%B@�$�P%	E� D�$� � �XBaD�$HB F�d �!�
@�V�$�%$$	�e	P� V �HB$P�!A�aD�$FT�%@�	 a�  �aR�)�iBA��A��%XFEXBTRA��!Q�`��b@�F!(�iP�IE�a	DBIF`
deB��$$  �E!	@F�	Q"@L�g����G��DUX��>��gz�e�?����EDU_����]k��?��������q�����ފ"������o������#���
����
"��q���?ۊ�*��3��QW����;$��e������0�QTQT�=��_���_�EU����i���C�����1EU�W����EU���?a��(���w����������������u�����掿�H�*��?�������������u�� QW����������g���Ϗ����f�?�?��0�������e5��q  ^%� �s2}p�y��d����k6Tl3m��v�ڥ�))��M�{i%t6�G(�mb먭ڨ�M���[5� u���4�Y�V�8=��4�j� J�t��k Prh �P(P*�����A�  �  �]  P��etr�      �=hݲ ��8�j�o�U>>��{�<�������=��*� ����t9�����O�x/�f�޷W� } :��t��w��/]�Q��Y�Usk�w�U����Vm���_[���7n����}�������f�{k�Co�� ��e�����;� V��÷5�=羠^��� t{0>�K���=��zR��%�M���t�{�禆��h�z΀)�z��x t�� t��p:� J/{���S{۞�M:.��=)s�Js�� ;� ӣ{� y��Ú�= �{� {��J]�J��  �u�Zb.���� v�أ�����y5�<� .�������݁�݀{���ͳ���v�;m���U��^ﻯ����{�׽��/S�}��ި{���!��������|'�w0��9hr��   ;���J�
�ݹ���U|�s�����7�pzw�����硽�|�u�C;z}ls���i=�3o���   w�p=���<���S��f�`w��<�)��n�c�v�kPY�����0 :>�O�/@6Ɓ���]�r�㲎��_ �� �o��<���_R>�{����|�ӑ���}�S���N���{  ����G|�{^P���á�`��`9޾�S���w�ψ�G{�N�S�     ���6�%T�F�"{J��S� d ��)MT��T   j{MTLR�  ���5Ji��@ 4 DHCR�"4 <S�O��?���l��������χ��_}�술��w�]*�����_�DPU�"��PQT����a#��)�I`K����?��s�_B�I4l�i4Xf�]m��/!�dk�˲SaJK���̉q"Id7��lݑ��u9�5�߇��;�>Cy����߃<{1��X�Hq�,���,�e�d���Y�w���m�vg�&�i4��P�\��������a�`�ۧ\Z��t�2�\>3��'�>����~�w[��*9�W\.�O��w�_y~�J�)u���u4���w<�iM����hC��2�7�5�d�%j��HH�
f̳[�ĺ�9�����"M����ϰ���O+���*}��Vﶻ��ݢ��7����.�F�S�g9]�[�V�&�56��R�e�l�K������������	�=�	��gWk��QZ���8�:X�wY�mU}��%�{���ɂȻ�͒_'D��e���1�!A�.А�wa��I�D���v�w��;8���2������,XF�k|!L4�lBD,H�%4c���ŭ�į��<��[U����4�u�c��8d}�q�9�D�eߑ��Z|�6�=�/�G%�G���Mn���m�ݼ�޳����I�GN����W)ax��.0d*H�{��'�ח۲�d'3�� F�a�u�y�G.f��B}���5���I3y.kn��~��fh�[�xf2���l��O0��Y	 Mp�JK^��R�J`�<1�9���-��Do���#������0ŉ	% Rp�'H�����4s���ϥ��[��r����|�G\uVݜ��k)**�_ſ�V �vV|U������J_r]�V���
��گ�{�y�g��)�ӕ����f�eK˰� ���a.��B`S���#�XO!�Î���3�(���	v���S 7�!����I���ኸ��	����6U��!���U��Uߊ)������w��g��V+���8@�*w7�!m<���i����>C5LM%%���CACDI�r��s\�r�%M�9HL�/.l���!7�|혶�^�B�}�c��p�>?Mk~(�		�8r�5�`��~�$�!��f�Y��$���	��i��VP��ߏ�/��7�;䄞fy3�ν�y;:rXί�7�=��rM�Q��n�s���|[������Uq_1��{�a}Kc6ZS&�k9<�k��%	!:%c����+�l�7���a�4HC#�Ƽ7̆�������4L�Wz����Y7���3�4���<��>f����|�χ˽�3�!�^ig���BG|��%��G@���GΩR�҈X�oa�Q�7���J�~����)�WW߶���ГN�9wFO,��gq,�����j�}}����N�Т��-���b{:�ܮ�/�~w�?^y=�o�k�f��]��es$�;]˺��\��D��� ᝰ��	���ф���'.�O4x�F���7����H��xO7�{�� ���/��5p�0Ş���ˆ�xFH��ˠ6K$Z"�p��I�5��s�BHqbW�G�`@	�hC�<��hq!���>=�A�~��_���t�����}��A�$"η+���>�s�Z��V�HUv�Yeoyt[�8!i��9f�>�e�)+}g|���3E�ωY���n�c�j{���K���}���Y���K⨷[��NY��IP�0�3f]󛅒ߍ��}����⸖
������ߪ��\��u�4Va醶�_p���=6K9=�������BD�j����|��-�8L��gQ�vQ�8젫��6�&$��W���-７p&Ye	RY�r�4�a#��a) R�i�Uِ(X]�9����}�q��aᐄ�aE+����$V�R���%�wj��uE%S�.�����������͕�Ey=�ݳ�4HGg\��I'�5�)��ir�(���]u�s�۝ڮ��!)�v���~��,��`U�����++��3�
<=,ӄ��h�q߬$[T'�OJ?J�P��%%u��\޺&��+|��eeeYG�*D��0̒GF�My?k�=7��$���m \VD�4ϋ�������Y�K!`^����6v��yu&���o���	#B#}�<�!P��W��"��f.eҫ���|�|�(�R�ں�y�1Q��M��EN�+<ٲo�$0�ϭֽ��5�3sXr�M����m���YJMSq&!M��-���� SXoX2��{�[�%oX]Թ�����c{գkRS���SQԲ;IH��\����lѯ}��j{��Y��VVѵ`�\�i�'��)-��>��R75k(R�7!52�ف-�uC&JL��9�BG�ܱ)@��ѻ[f�R���3Z���==��Ώ{�����_C1��	s|t���	$a�p�4͛��޽��itf��)}���<���S>ܜ�~O!iI M�f��A������߄!= I��]d�:���4m!�	Lܦ�1сHԔ�3�^ �����7sY��r��9�F�棨S7�x�h#":40�H��cOW�6YP���~���c��+v�;߶v���;*Su�ғy�3�iz�� P��y�!Ny %! F��ff�Y<|�.��R���������WW�J��9wܮݔ�2;$������Y�\�&�z�ty)�c5���>��[�-�������v>|��~�t}U�G�U����N�x-Ⴍ����߫;���h�I�7��y�J�2OR��'��Y��/2Ņ�˻w�K1���}����)�v���7(l��mٗ��|k��E���N�j���Ä����߹����y�r���.$#	  �ﳯ;[���l���P�(p��j�f���Bq���,~#A��zkl��n�y'�x�y�]rYw�f|�s���5���8(��� K���2W�����'�S�7��]���6���)ef�E/��
{�0sb��\vF߳��<���¶X�95�H���[�O;}6�꼧�u�>}�q�_8(U�o9��W>�/�~����Fhw��~����'FS�)���������??�ܗgw�J������y�G�_�O>Y�n�3qz�!5�Of<�'Nd��y��2�|��b�� w��$���$�c�H	��
��]�C,cW$�K��1*@���7y!�Z�a�~$�2J�1��aI�8M��6�	���a�4WV���[8�{��i7S5M����<&���\�ﵾ�_nƊ�z8z�Gٿ�����s.�g7�X��ʢ���Zݔ���oj����\>���Zݤ,�B�k��������P^bi�;!u�a���1g~'�;�6�"���N��<���]�y�.\��fo�.˴�w+w�JYw��]�s+��Ϭ��:itΙ�x.e�j������F�c��@��a<�F2&82�i	sD�zq�8�jo��������%.沚۹t��n�����z�,#4i)����Cj�5��2�ti�G*='&'^Bv�7]ܽb�q�9����w���Lk��j+���:qVv����3����K�й��Y�o_{:|Up��]���w[8|���V}�7���AA����]4��0ɣ윒i�/S�^�X2xr��%�NC�d��a�ݣ�ﮞ�S��e�j�<e�x�)�&�YuIa�Mn�wd�<�<v&���&��^h�n8:��Gr�u��{�8I�Mf�+k)).l�]���p)��0,�3�߷�o����q�5��L��#oZµaIK��&НFi:s,������w�䟏|��O=�眞%=�P�'��&�H@ ��xOO�;�\\c��~H.�i.����lɿs���:S��_�Y������.��9��&�g3z7y]��f[����7[��r����|�]s�y�Bk�S�6L�U�����Wv�o:�yr���CY�/���n��qT2�w�{癭�|�7��<�َ����i)�0�.noi�r�@��#��zL��$Ԇ��s�ͭ!�e3�6U�o.��u�ýWT+Y�jO(��̸9�so9E}n�|�]���Yt�Wr�'~�n��{٨/�l.���/a.2�nI�4�~l�!d�:�^�o<�o�!��;�F�RS��BC���B�2q��,���j�����,�W�z+�.c���/�7���1���z.%�G��[z�/[����4�{��1�7�I������Ww4k,ܓYf�Mo�s	rV�<9�d�����O`jl޴j��	FH�XK!m%�#i.K�i�� pGb� q ���������D�Xt�qc��RZE�ߛ	dBR��aXg,,��Y�]4���AX�yA�YG{��T$�n�6{�<��4\���m޷�*HP��9+.�F���%{����<|,�9\X�����c��u|qqB�r��zܹ�$��o���>u�xM��p=����	�?&L�}dܙ.@���F1aa!Q��I|�NaU�B*�׵���u]Nв���g���q�! '夙^�M�Cwv��C�y�߼�l�o�^bJBg�W[�[�B�@O�VSL)���-�j�a���Ç5���9JY��K4eƲ�U�VK�0�ԓ͘WrL<�q�c��7d�-�Gý��>k`e�a+��0 2ܦwXV����{6��y𗼗vy;��Jkz�e���d�$���1�oT����<�O�O��vśχJ�}�Y(JR���>�YH��l�'��}�'�Mr�C�=��<���+�Yq�2�1 c&��s���\=��ea�|ߐ��&��#~g/%�����������V+r������e	��Qu<ݰI$��d+,�!c!7��b��n�Z��:ft���l�^�9i��
��Z6۠���B$!�L��#a��W_s>�;}�uq�e`���e�<�Ǿq&k��0��ux�	��'3N�	�d+
��Y!X�In�,ń�x�U�!�=��c�����{g��ėlaR`@�5�{���{�8��!m�/�:/�P�wIa��&�}����Vy��y!�0�d�-��d=�I �hȑ!L<��05�� �eH�"��<&����1��9<rtݯ(w���ml��.����f�5>c��9��).�Ff��9��y��Bo�d�,��r�[��x�؝^ws6oi��R����[ꇚ�uܹ��	��Y�e��}���|5��B�t�q�OY�$�8l����2���%�4�-�����gÇ��kݓ��;-�����7aQ�	�ʼ6E"B�[� �!�1�:��Cq��@��l��%����ܹ�]�6�BB$�p�fG�)���sf4�r�Xi����٢!湳Z7�K���j@���)���tWD���e}ay�ͅ����w�&kZ��X]v(IB���JKe8�y.�3�k�>=�>s���:ݽ�y�3Á4Sq�~��9�M���Ha9��N)w��R\8d.c���;��';����sC��K!����]}�R$Y$�`E��w�U�'�;�'wǎyJ�Kd���ِ�=[y߹��n�>���g>��6�̻dӾS�����w��	X�ך�a:p���^�|�BenX Hh�����BOH�HlR�A)5�,�!/��onh��J�ư�M�@�,m��̓.�/�=F!���}�|k���k���B�i�f��5᤾rg��A��5��&��%1q7R[e�g����d)����ry�!��_����ꪪ��U)-UUUUUUUUUҪ�����������T��UUU��_UUUJ�UUJ�UPUUUU@UUUUUUUUUUT�������������UUUUUUUe����ڪ����j�j�����*�����U�������UUUUUUUUUUUUUUUUUUUUUUUUUUU[UUlL��*ر��yze�eD,��R�K�(ec;g@)�9�d ���cnrq��Uم���[�V��,�F1�\jUkm�-��4c��oJ�u�@V�/F��4��R�0�U��\%�9�ez�O�TZ9.�d����t��.�Lm�l�!�����)����ۯtgZ9�9����r�ju)AU]�{td����T�yN��mU�vͳ��N����˧F�%m�ѳ������(0�]�Ƽr6hV�nҋN38�3CS#�H�P2��"�6BC�[�-l@��(�	f(2�4CcA]��c��
(�l� Lf4��3TMs�xCl�M�Pp�V㰮��c9q��R�ul
��.���g�;A@Pvl7R�j*{]+� �u��iW��@]�+mQٙV���������|���V
���܀k��X�M�&I�v �g��������Ö���6l@*�+�S�y� ��d 7��e���lpg�����FF]�j�m��E�����i(-�R�d��	YDv坛������x�\����<T�y��>yqI,��6���6�x�+˹wL�zI畕v۶j�����hK�U��L*��
���Y�-���ޗ�uPq��ۣ� �#]uV�[r��l�e�
�n�h;QYW��y��3��B�m���3ͷc��T�3MC��*��&n���������PG�ڭ��]�Tf��m;�N�z�0�٢� �yW�m���yK!�C��ai��%Ƹ�U7-��0����}�4ہѰ#�ERU&% �G�+�s�s��bU�Qi�}�����Ug��U���J�R�-V�G,Rƻ	+QEeV7�TV�[7S���٠6��MW^����� ��d�8��j�����`y8�n�x!�F�n!@z�fw]�i�ȣ��dz�t�<m������Y�n� [ �{�=N�˰��*g`Z��)�W��Û�8�=gQ��Q�^x��D�\�μNCY(��eP�L���)t���YL�H��K�]����dL3\l�f���`������V�LK@�ţ2X�4��MBke� "��^���ѷ]�Ȁ$��Rghsz�uq��e�����6.c&t�q��������F�/��{��E �J���sҠUFtt�i�����!�g�&�E/Jѭ҅Z�e��򲩳��	�=�c�Wd��k���um�3�
�8%�`"�ALc9�N��CH<�J�vc��
�*v��{6�ri7R�L�U���8��f������z�
ۑ&*&��� ��ݲ���J.4��ip
��Ғ����kU�ËGcnێ LgF�k5]
�<��H�dr�z�p���x�=��/`���BT��#e��ڪ�	K�UVڮ��o.b��WV�)YĻ;֞h��J�Q�yڬ��g�z���4\�il� UЬ�뢄#M�xM�����{XH6WTx*�דv^N��:ӳs��G��@y�kj�ѳֳ��k�e4� �s�����-�z�;�J�r{FL�c��g��z�2�,bZPP����VN+�hLH[�n\���k��9$�-)�	˕A;i�֌6y:V��2�r=�ct�]����"hS+��ñUv]����q�m÷d畍��f�07l�bu�t��s����,�L^�A�j�r6��=W"�� �m���j�����hw@hHY�N&m��9���9��Vֆ�,��K����[h���C�*�L;)��9��m����b�/J�;�n�gm��MF�]Z���`m/����k5�������{ʅAm-��Br]pq�E�b�T��quO{m��r��k=�lFn��� j0I%u�8�����.>�MոӞ2���*�<1��0���mX���԰˶���b�����=��'�iL�2��@�]��W�̙�� 97kr��I`J��W�[���nj������n읒5�	�K���U
�Z�#��h ��2.�
綪�&��@�m�Hm��*^�y�Llp:r��K��v�Ö�<k(%���.��<�U]Uͫ���-�4�ͭ�+R���.�� �km�,FiWM,5KÝI�(x籰�	F�+U�l%��@�TL�^B�c�{g�F�峞��c����b7MT��iW��ɥT+������\mq��YR�j-��'$R4-$��VʬXW,`�0�ꩪw`6�Lk�X���!���m'WL�ݍ5й���]vY�����5A�(r��O9���.��u����ܨ5�^%�Yx����6�d���0�i�Q�lh�C�%c�zs�N���wlee�7aCI��u7W v�{f��
T�$)�K�Xs���˞4�:ܽY�Ѵ�l��Lt�ܙ�@���u��ͻ"��U�Y�z��j�� �v	@I[����ڮA�̭Ԭ��2�T��e�[R�i��MCWA»�9�<rɗ����*�C��*�ĥ��J�\�KY�vD6��K=��o[����HM%��+"��Acnٔ5�B`0��ٴ7U:*�:�EV��s����Q���Fy3�ۉWe��T�5��Z��ش����͎�!f�Ѷ�v��5R�\��:�[��5���{b�f�j�K�R�q�*���e@���ʢ�3!��7Ӥ9�b��Bk/
=X6��U�yggr���u���yYP1����V��"cjD�u<'L�J��&I k<��:8�ګ(��j�UPT�����)�f��wPlGh�YN�UUuU�uU jU�������-{j@�\�K$�x��-� `��c�����e�z�2PpU� q-�@+i��"�i�mJ��&�
��UUV�4S�:�}�\�d�	aM�ʭ켱[��{,�ꌝ�`��~>S��"m�jl����nYe�v�*�[B��F��$���5AKe�P%y(�� �EmUYF��i`��̂hi�m�U�qEʄ�UURdGT<nX�c 땽jfmI.��b�V��N�ջ�U���]2<�5kƧ�R�9�n�8��{Rp+�q��Z���M.ܴj@]�y��mّ���n۪��@��4����P���l�#U#��)b�� �vep���W,��aİKj6n�M��P�2��ƴҭ�A]D�
���k���m�V��n�+&��땎)j�89��ѩ8:Æ�{7Y�n����1���/���!�C8c�cK�l��n��r��<;KQp˸$�!��.�u/KD�b��J=E ���z+�	���6�d�{s��cfH�m�1g�&j�ƴ)�=OR�:�.0�)/V��p��v�@� �Л���;�����\=6�u�����������*����؝ѵT��*�m#/��;vz���<��"���2(K��$�5G�WZ̑$Ѹ��`��vXN��1�:���:�V�h;s,���ﾗ�<�&�vM����R��������B�����`�'��T��[��Þ�����\�g5�38e@WC�tZ�X{Q�hZ�A���%�v��j�B��)�KY�:�UUP���.ڗx�h+Ѓ^�-m:�.�)�ͥ�Nݨ��X�͇
K;k���3'�e���0���$j$���у��C�'wt S��Ц�����X�A�{T��a-����H�%�o 'LX�,�:\�Y�v�V����.�fv��j�s����$���t�n�,]*�>�DN@���5���<7j�l+�R��UUU�����=���'c�ku�ŵZx�Y�Lde��:���#v��ۂ��e�ܐ!����{�/�F���,aN��Ī�I�sR7�:h-i�.R)-"�<`W�ŲlML�s�����+J�"Y�&n��N�����a��@�l��1�ю69j���]���itm]T��Sʇ�6�_.QBj��������sv��2nr���tUl�qs=�-�M�Z��:��k@�\/^,��eYOHlA�ԡ��uP�W��ڔ�j�fki*�Y�I<�D閩S���4�U�Tղ+6��l�U�-�ڨYYZ�۞v�Z�`*�
��N���VV������
�S�n 2�U,�UTPUV��5�[f�����f@WU�ηnZ�	Yl��k���y�n�vֲ���K�*�UUPUun6�*�W��
�V! �.P��6@iUV�����Yj��U� ��WU��@U+rʁT1�j����K�.S��UUuU@UU�*�UU����Uu mK�μUT��v��V��^smHP<��t09�\����	T�r�V�`� w����↮���P;z�j�"Y�j�U���+�=[D�FР�-#m�0��כ4Si��`*�+��uTЖ�Rdyv�W��Z���c83�ɴ��A�N�Of�1�SQ���
�k���3�E�[�M���}|��1����X��b�Et4����f�j銪���UUUUXʥy���8�eZ�u�RB�D �]X�@UUT@UUU[[b�%bn����Ӯ�P/ �������e�
�ye�g��Ҫ�(�keӳ��S�m�
��6�6^0�Un�n˲�[y`B�#�l��]��Eq*��R�UAX��m�*U.���UUUPqR��8���R�UUML+U�UmmT*�U�U �˰� l�9��v�;��mmUQuU�ˆ����2I:wER u�	�+�)�}��UM�8��`�BlP��$b* ���D����H,,(�4&�z!/-H��"'ʔjr"J(� Њm@(�d����@S>Z(��`@<A*��W��#“O�"��U'�� �� HŁ�X��I 1�-j?�U��P��		� �C�%��0B�$jCa�G��� 0��D>(��|E� `�@�#a$6*�{D���J
�&��N<�X$�`D"@@� � ��!�*�|��
|�+~�M��$H�Q$X��$d�� ҡ@�|���D��B�!D*��h	hk�'�> %A6�	��!�_M�BA�"h N f��@�TߢH��	��_P_ W��]EH�OE ����F�hEy�~L0= ���~�)��O�� D"FnN&�(�z"1j��(����|����>*�? 8���l�,@��G�@>��(�HԬ@�(Q[P�� ���D*���2	"� ��;G�>"ʟ ���"! E���M���-AC����D}E� <D�&�0CH�J��D�>G�P��m������P!B�$"6�"�F�J�ѱ� F֖��!,�H$`�$)!�am�`�H�a,aBB$����A=��xh�		!��B	�$"�	#"�1��$ H��@��@wH�>��J�Dd�@8����$�#$�"" �����" SA�<�!�!@8!�8
������
��=��Z!%*� ¨���� �\�"*��H@ؑjE(
։A(AR��a(
B
��Ԫ�C+0 1)H�P �։�k��UV�T� ���Um@UUPm[U��UUZ�v��&&Fۭ����i攍n��cm�>�R��L5����ŗ��.��\��&��c����c�.J�EN�i����˕і���Ĳ�2�Rnk�QH��5=�=���ZY���y'k6<�d��ŵ�\�B�A&;:�`cj��Z�k�8�B.�ȱ�x�&�*��[Ԥe�n^V��Ĝ��T��HX1-���Ґ�ay�1��2��t�a-x��ĭ5wr�=g�c�Y,'9�C�k�-Dcl`�oAh����rrd�Ay �,�[e�,l���s���&ڒ,�!��uۆ���lV�dA^�iuO
Cc��\s&ػX7[�>�i�u�<mPO8�d�B�;��rg�&p�yDx�ZӒ�l����%)C[vܙ�dV�Ȗ�탉�1f]���̶�-�%��BTj۬���=���c��c�F�M�[�e��v&���xɥ�P�8���s�m��3��<�nƺ�M�x[�m���=��qõ��g�	ƶܨ���֯n�&Q�K,R�Qh\P&���6���N��(���V��\��� B/m��[�=��W�[v�\���r� uf�ۏ%[��m�;��mu��:�)	��s��kLv+q�;	N���;":9i
�,MtCG$q��\���CJ��b��U��+�F%�]��l`Q6ǄЊp�B��ctj�TC�i���l[U�'��)��'Z�HXF�L["�6��m�[Hg��4feK**�ۣ�@6ۭ�b�u,�e�ekft�E!�{��F��WgQ�؀l0�H�YSi�1h$u�c4��C�Fv�$��fᨁe�bЌn�����#����rlKʝv�lF��ʭ��@�u�-�ы��r2�e��Pq���]��nB�&6h������`�fnݥ�І�{V�.ӝ��PA�)��U��6ж
��4qx[��i�\�X���F��bZ+v��$��L@�?#�W�G�)�q'����
�#�� /�>�V�	��s��⨚�$��lz��."��M�]^��v��]��9��v{Q]�5um���0��iJsp����Y�݇N��nn��L։`��toYa�l �J�4�ƈ�͌��;�ŉ���*�HfP��i�=��N϶ݥ�*:	+�<�;�v �r���"y2(�۳v�:�X�^�C���yvc���V�#K,�{k���i7��(�5]:O��t���<�4[��ȼ��v;ÎW<��avL��{9s��s�\.���^$�L��u08�����U\A���e�:�v|�m�`]�y�vj������{��j*,M��4���[�^������/ �IHMGhBbi���� �u� �c� wdxV�W�uJ�Wdi]��_6�ـw�� ;�<�v+�;�� �U}SfIݯ��&	����qȖ�H�d�H�gESX�p�z�8ta�M6���͔�L���|���^ݎf�`�,�]�E�	h������ۻ�<8rC�O%��B���>���˯���'�{����<lR�m��Z�[W�n��\0��|�����W�qT6�]�;��M�f�g� �{� �O+��)=�0���t'���I�v�0�G�j݊���vk��9$��S�~�3GPؕt�QS��9�쳓���6�`8�Qv��	lM�6b�V��զ��o�E'���� �c� vH�We'�i��.ڼ�0�8`vG�أ�W��F��I��c���`;�`G� ;$xm|>
p�DH�$ 1$A1�b�=QNrk^krN�8`�ē�mһNЭ��0�#��Q��"�7u� ��VR��E�
�lv�x��<v8`���<�i�+Wtm]�����t`G�nFń]n(���.���5f�[��
�۷I2����x�Ȱ�p�� ob� �m�V�S�c��N��7�ឯ��H7����/<v�X�wr�vP�ēC�m��#��(��U%'��l~0��+Tc(I��MQv� w�G�n�{�yҡ�P4�/PW�3����'�~$�4��Lv��M��"�7���< �b� ��}^�)(�42�.�uaU�5�f��X9�P��֭�a��Ldn+i5�\:jVf�ηh�տ ����< �b��U_q��,���۲�:�[V�0�G��Q��"�7���ee]ݺ�t����6���<v8a�� �{� �}���S:k���^����_}���@�� ��{x6喝*t�v�I6`�p�=_-������{���nIM둮����(�R&�y9��oJ%.��n�Y��֩vlR�2�h��
����:v�9x����js�ާZ��q�枹���ͬ!F(���5�hXABA���[�c4(SC:�X�n�v�֡vv؄;V=��kvC-GQ�d�m�ۭyI0�)ĵ��9�k&�r�Q����ր��v\8��yb�� ��jF�g��Jl&���}4�^�=��B�&���Z��R�T�m�]��ԭ�oLjxk@6�������4������;C�JS��t�����bGJ���v� ��x���v^�������CcV��� �b�?Wԑ��l~0�G�r�PS��BUv�n�4��v^�� ��{xej��V��Z� ���杖ٞ0��� w�G�jݗ�rGN��ӡ��m� 9$x���v^����}�W��x�ʴ�笋8���s�us2`�s=���5۱$u��+l�[��0�nG�mU��o�<��v^ vl~���靖��x���厈�6�C#շ��=�ye��{���a�Q�K��
�x��}U_{堳�x;�< �؞��*Ӥ���nݷxٱ�$� 7v'�jݗ�w���C�uv�n�]��=U_W�w���	'��5n��͏ �kb�F4*��Ct]����5n���G��<v�X
Uӻ�_!7@�؝�cz9�Mtl��{9�͛�a�S`h6��.��P.s�l�V�<�um;� rH���<Wtw-�.�J�����G�H;�y����[���ĕ��;B�&��I��}��sv �҆��߳`ݏ �$2˴軡]�Ӵ�����[�����$� �����I�M;4���jݗ�� 9$x�؞΀kWbWWHUh�STy�즜G���n��M�۳K2b�l��ֳ��.���r�y��^�|��^�sv'�jݗ�w�p�X�Wwm��m�$� 9��5n���c�9�حQ���lhn�����<V� �v< ���)�r��-۷J�jݗ��ǀ�<�UV�"P`�zS���5]��x���v�]�ݪcHM� w�<��Ի�y�d�x��x���2vU�=���E�`p+7A <�`b�866��ݺ:ܛ����&��l�o 9$x��<V� ���	�T��.�i���o 7v'���H�O^ n�� 9$x��m۴��Zv:i[O ջ/ ;� rH���<���M:V�t�m۶� ;� rH���<V����H��.��x�#����[��y��krOY�`V�b�e(P�#$ ,��{'ۥ��&�.e�eգ���y���ZGM���B]�R�0ٜt���`���x�s�a���������˹���r-�\]l�GMf����ny1�r�0f�7Ɋےwc��i����M�Ye1���B�5�iK�p�j�Jˤ��6��^�p�B�v����s�V[20���tm	�q�L
�6��K�3�k]����35ɒ��L���-�ߏN�I�,�}m��?�z�h-+	]��,1W ˸f��Q�&���Rr0�e��&�P��lhn�������[�����$� �II�Wr�Ҵ�J�jݗ�� 9$x�؞+���]��Z�4���{#�I wv'�jݗ�l�J�1Rt;Jح���< ��O ջ/%���'I��:��զ��M��$�wb|�I%�ĒK���$v�OIv�A�n9Q�^$���i�OW'ci.s�ca.�{��<�<�������gY����q$�^�x�Iw�>q$�nG�W�̀<�߇��<��}�eb�nT۶��{���z�V�B��H4p �V0��A��[�}�f��6D�Ē�{�I.�����I+-��|�I.܎�$��dO�I-W�^$�?y�}�~�z���R�jU�ez ;�>q$����$���|�I%67�$y��Ѷ�T5Xl�}�zo=7@��ձ�$�doI.n��%��������Rb	�[.�q-�7���Pm��g�zΠ�4�&�\ൊ��X�\�WĒKd��I.��$�\݃�KM�t y�� ��k����`���UWv��8�R�z�^���O����s�`���vu�`�\��o�}ٮr�}������-OI�T1?h�)��{��QԴ�M.��1'����
�sU>=5��7���(��n����By�y2ZY�4K0��a@=�����%�4i�u��5�1�aaG�|,��U�H�d6f�]Ը��}����x0������=���{ �LCh8����7ͥ4��@�~�9t�f�<�d߇9�M�M��� ����yn�^o�ԻǑ��Cy��/7�����<���WH\���l�ffj�9��NL���7�L��0�g ���!%��i�'�s�,���q��"p>�S��ӁH|<'(F�w乢�	�7�s�=D��=c�H�(�.`a2�-��f�I$w�H�N�cS|9v'#!&�!E$��sV�l��1�BJ�_h�aHKˎQ�L�Bb��y�,��l�)��A5Ek)��D֬i)i!.�9���s�VD���	2n�l�BBI*kV�uO4�Up3E�W=�"�y�> >��@� <A�'�|��	V(	��"����^!���#W�x*i���|�I�-�I)��q�whn��t�m>q$��e�$�]ݏ�I!vKx���'$�����=��>w�[V�dT���$�]ݏ�I!vKx�Is��G�y�� I<��_�(`��j�A�E�k��8Ӽ�{S�q;��3�7��\�hӴumZ��Ε����}�z �y��ؒ۽�~����Il�|�Il�b�F:)�*�g= ��{�ͼ�n���z��?{�z�I6���]���s��+��8�R�z�I.���$��%�H��z=�}�{���iX�P]�I$��8�B��$��v'�$���W�>$
U��&�^����37m|���u�:Į�U�
~��� �������ޤ����ĒK���I.V�?!1�E �X�X��n�ٱK��N��W5�9�Ό������,��0�n�$�\���Ē۽�x�Iwv>q$�����<�o\��:��}���e�$�]ݏ�I(�b�I$�݉��x��m[Y�[�۠��ߟߒK���I%��O�I)w��Iv�B��ae[�6�Ē��+�$�;�>q$����$���|�Iwj�Uu����J��۠���M�`rI'���v�߾��m�3߳7m��� �}$cd�>��as�CR��2Jb4��v�*����i0k��2V� ����6��C)x�P.�p�q�g7@gC۷kͻ0��u���g����Y�F5�6�1�4��	b�F���j;���� ��,Bؔ��v4�vKbp���s�4샥���	������k�v�b!�a5�2��ۚs����o��:�1���h@��bh�dӞrri�9;������N	~�iV�e�%Fu��-tm88�����P&�����'�v(��ts����{� �y��`��W� ����}�{��-a�����I%�����]�Kg�ĒK�<�8�]7����}��F�C<�q�r�� ���I$�݉��w���I%�y�"����]�v�D�˺��=�{�$�\�I$��8�K���$��՗��: �P����y� ?ɼ��>�$���I$���$���M��n�6Q�b�j�0�����b8����v�m���Tl�O�YӺ�(̙nT݀%�y�$�{�I%��?��}��X����� �e/��j�:VT��`����NO[���ϻ5�[oٝ�n�������99?����?�,�ul,Z�e�= ���=��o=۠�}<���H��'�$�I��J1X�[#�`}�7���t {��}�_��]�I���~� �_��mvb��hP�x�Iwd|�Iz��;�I%�<�8�]W�����rM���;�n���^S�|	�-�JKu�&U�"�q�aԌ1P����9^���\g��4ʾx {��w@����Ē꽊�_UW.�Kg��Ē����r���Jl�팻� ��~�����+�W�$��y�$�{羯��-�K�v�9�2�G��<>~�����w|�@��O�5�BA"��H�!�� # |��U�W������ �}����z�c����9�[��Iͼ}���`�ߝ� ~���`}9'&�������R�>�M�2ʡ��`����'9$�y�����{��P��}����7�MpO�,�:ps��5�P祛��s�R̖�i�#�*���f��>�I�'��!=�Ů�(���l����Ē꽊�$�od�U}U�w��[s�t ~��~���
��6G��?߮o�"~TMkV�����-�����ݶ���=��rrM���}�����AU�H[rz�$�{�^���]���đ��� {=��H�&cH�W;��{���\�I$����%�{�I�j�Ȅ�d"cd��hCA�U)�_5����ϻ{w�3Ff�ö2���z=������v ����$�{�I/�U���!�Gn����F�2㫭�ꑈ⥕ BH�Y�[t�V��8�~�N�<�U]0$�S|��}�n���=�� ~���'9�����������2�G3*n�/���g9�P�����~�ߵ���~��������u��I�qPf��oѩv&YsC;��7�;� ���G��������$���������w��&�&�u�ũV]�tӒrm��߇��=�?S����f����P�~���rOzw��V�ր�̻5�y�����NI���Nz����I>�?~��O<���7�O 
Q	O}�Q���"�浅T%���Z�N��T#��va�1���
�µ��[��;�9�	�D� ���� ����Q!)�i�fB4-��5e��(�sk��<˽M���zӴ�� � �ͦ#.ِ���S���bXˌVk��a-�B��ۗ�L���S"������ڜCe]��I�OC�V�b�'l�FM��9�u�V4*8��\X�a$����ϳ��s�/r���	6����\2݀3�"���6Ay���8:��6���Vܲ���ӏ_x���[������\���^�܋ ;ݗ]Q^Y=�;۹'�;���E�hԦ�Q�x{r,�����UUvE=�^%��������'9��M�JGl*�5l������KT�� ݿy`<���Y��vf�f�s�9?��S���,W�~�������m�z� ���o�]3V�eV�/�}��$��_����U��Ȱ�$'Wv�s�&�\��WY���5�ٰf�����H:^)�C}9�H���F�ؙe���y��ul�x{r/W�}\A�O^�^h�~�)h�ٽ����w���9�N�ijnuJ�ZC*��&bE
�(9!JD��pLHz�D�����	EbX n ��@۪�Ab�6"c@�\@�@M�1t�(hX(����N��Rw�{��'g����Y���H�YW�]��i�m
�x��< ��x~��W�Wr_�� �<~�a��e�vЮ�I;�����_}K�{��n߼���<}�UU%��<z�]�V�j���� �nE�~����W�^��@$����2���B��R��WK��\ۡ*1cpu���ax�<s�&�h!�ٴٴ�������%��v[w�?R����w�x6L��}�}\A��e`��m�wM�ݿ�]���ﵿ��W2{��ٹ'��߳rO<�s��QKO?~o��f�`��ez�����y|�����=dj5��HJ�JI(��� �ТP�*r��������;]��)�j��[�`z�����׀wn/^ w�<}�I����:���&��R(�$�;�s��^磌ꥻ�>�=��uvK�4�{m=�Pf��4���ڎ�MN!������6bkT"�be�ep�vB~�N���{�vj�N�jէ| ����ٕ�uvK�Ӝ��e��ޟn��}��]�Sgcf�ܶ�n̬�UW�|��}��;�� ;������9�Oz?���K�5r΁������=�f��? ��>���nI�~����ͳ+�v\�9�Ӝ��_}�׹�$���[�s߾ٹ*�b�0>�!|^�6,�BI	�p�T�tPdSP0OP>��k~s7$���kWk	r�C�� w�<��}���������@�~���oo��|���l-�m���<Й��XM�DmF�ZFӜ�ҁ`�=�ǘ������;�z�i�4r�_�y��ݝ�䗀w��_����� 7}�mm׃���v��[n��������Hݸ�x�<�l�Y���H�4]tXƚ-����n�^� �v<=U��Iv{�X���ͭ�R��N�n��k��~Ͼ��nI�~ٹ$�}���@O�9$�����t�����+n�S*�l�X���_U^�ߟ@�~�׀�ǹ �|,�%�a!% KD!F yR�B�"M��ߪ��1�C%��e��q�P��4A�A�͕ ��� �@$}���8��"�F���6�>		Iu`'	�|L\Mz@4��7J��e� B �##0!f��j-��R���`a]�H�=�!7���� �wRh�T�Q�[� L@�0�$��M:�+��D	��|�1�n�S`B]Jozu�CX�͇6d/A����73k%�1qۋ�Ou��8�],ӥ�K���K[	t��Ѻ�֤e`��X�)lI���n��%Ӻ#�#���ܛ��[U@uUWT9@���*��kk(�uUUUV�P&����oNm�5�:�{���p�4��pɖ�kU��˄�k;��d7Nm�9�瓬f��m qȭ�Bj�Ol�����Q�<;��.��%`����u��wm��,Ĳ�
%�$حr᷅eYQ�S5�2�E����e���X��eƫn�;M���ǃt���L�j��XY��9���[Κ�H����[���kκ���;[^��p�u�cx:gvܦ�OCT�ѷ�j��),Ơm��К�E��TѦa0�*R���Z�^.]�l�on��k����@g�/СÄ��N�^poZ��Ѻ��h|a�����Q�w�Њ�W�̀�C.5a6p\��0F�ԋ68��8�����4tA5�K�y��:��ka*.ȸ�%s[G/���bE���&�`�
����qk(�l�c�r6��uۅ�nyv�t8r�GA5:Nq��%+q�p��`*��\�I�*l	�����fjűv,E�1t+
h-`��KAz�6�m�]=]���6@F�k��n��lH��[r�t�e`p�;x���qGA���=�����.�Sny�ݖz��ێ�ۨQ��&μa}�u;f��m�T�6�. �̀k�ͭ�lQ�GX�:s���<��GGX����	�u�����Gl�&�vwή+!���6� [b�"�f��sҩ�D��U�݇Vf
�v��O�*U�ub���ՠ�M��A�@�k�FL�[�E:��
v)��E�!u����7� t���[n�μ���٤���y7"�9
��M�.ٹ�m�t�<�[,1KJkP����u`6��l��n3cd�U�<Yh ��&w�n(X��h����o$iJ9gou<'pS�˶6��ݣ"�C�U������<ch�g$�>�g
���p�E	�V�u[�n#]
Y8\����4�g1Z�=��k���ɕq[���.<"e�˰�ӆ-L�VYw`��ۥֳX�`"�{�"�@�"ix
� a�QCGT�Ҋ|�"1W��8��/��& �EQ�����%��$��	��X�#��-3�ܚ)+�i�A 5��Vb�.����z3����9�d�cS�*�;C<u=�3��B�h���N\jP�6E�i���ݺJ&�D�8�wV��4��Y�M0��BR�;Na�e��Lr�gk��r{;�l<hq8J�9�k
F��Vu��Q��v����{[��I��Ͷ0]b���-�/>k8��Px(&!� yx�0ˆ[.[����\����j@\8����SF��q60�2�7�b����;�h<�g�#Ug��������Q`{��꯾��;=� �=�.�]��;+3��y���{�rI��Nrl��� �~����=�W�|��z��,v�Ƭ���k 7g�͓+�UW�����Oߞ'���9#W,��N��-������]��+ 7}�w�8`z����}�mm׃���v��[n��������݆x����9�e`�}�;cB���ٚks���3��f3<^ۦ�lq��9�2�6Xe��}'t��t��`X���5m��O� w���R>�}J'�w�6����L�bX�߿~�ӓ����/'����vQ��r��:��Kı/���m9
�y��!aTh)H4H�) "�Œ�X���# �a�F$X��B��H	���T�(Ȝ�bo���"X�%�~���ӑ,K��߷��NEU�,K�va.p��R۩�ֵ��Kı<����Kı/����r%�X�'��wٴ�Kı/���m9ı,O����K��f�55u�h�r%�b(6%���[ND�,K�g���r%�bX��~�bX� dO~���i��^��צ����J�6U��>D�,K�g���r%�bX�	}���iȖ%�by�{�iȖ%�b_=�u��Kı==$����nN��ځ�%���^�8�KтTlD���u�k)���wO�=���k��r�t�zkŉb_}���r%�bX�}���r%�bX��{�l? ,TA�&D�,O~����Kı=���ڙ�a�BjMf�3Z�ӑ,K�����ӑEı,K��bX�'��{�iȖ%�b_}���r'�b*DȖ'�|�A��d2gy>��%9/��~�ӑ,K��߯xm9ơ�="��.�b�2&D�k��ӑ,K�����ӑ,K�����{sFd5��1�ֶ��bY�QV".D����ND�,K�����r%�bX�}���r%�`D"�X����7�g��Kзh5�2ū;9r'�{��pI �}�iؖ%�b{�{ͧ"X�%��^��r%�bX�{�!w �%���nd�����񱛍��B��CIՍԷ�M.p_N�;z{Ԕ�n�3vڙ�k[ND�,Kϻ�ND�,K�{�m9ı,K�^�b�Ȗ%�b_}���r%�bX�u�}��M˚�52�ZѴ�Kı<���ӐUı<�~��iȖ%�b_}���r%�bX�}���r*)bX�'��{�3A�9�9z����������|���Kı/���m9�,Kϻ�ND�,K�{�m9ı,O:v��Ld��"{���^����wI�O��]�"X�%��~��Kı<���ӑ,K�a ���"@�& �)h������AdN��s��r%�bX�����Y��F�Ԛ�Z��r%�bX�}���r%�bX~A"������yı,Os���m9ı,O}�ݻND�,K�߱SB1,T�c��l��mҝ��xյ�
�(7K��f\2���=$�oSz�Fױ��ɫ3Z6��bX�'��{�ND�,K����bX�'���݀<�bX�'�w�6��bX�'��M���l5��0�\�m9ı,O3߳��r� �DȖ'�k��ӑ,K����p�r%�bX�g��m9�,K���wRh���e\�rwy�^B�y���r%�bX�}���r%��by�����Kı<�~��iȖ%�o'�O~�c��mF�L�듻�^B������"X�%��w�ͧ"X�%���;�ND�,���ٴ�K�����{�֐auJ�Y�'w���%��w�ͧ"X�%��D �����yı,N���6��bX�'�w�6��bX�$8�B�{�3g������n�޽F�m��Pb��.͗Z M��v��C[�u��dһ!��hC/���]6��V����۷=��5�=���,�p�vq��W�(k�Sm��s'!��hĠ�1>�uՇv�p[A;<�I7�G����Vʼ���{puHEX���m����`���Lm �	�k�uat��Ml�i��9��,�$tt�s}'''<������,�!��!ѹ�YU����minR�[
j��=�"L�,\�g�����
7X�uf�Y��Kı<�����r%�bX�}��6��bX�'�w�6���,K��{�ND�,K�N��5���˫�\�3Y��r%�bX�}��6��bX�'�w�6��bX�'���6��bX�'����m9�,K��y{����Rjf���iȖ%�by�{�iȖ%�bw;��ӑ,P�,O=����r%�bX��{�iȖ%�b{��t�4Y�)���5�iȖ%��'s��m9ı,O=����r%�bX�}��6��bX!by�{�iȖ%�b_>��|R�tq��'w����/'�wٴ�Kİ���?M��,K����p�r%�bX�g{��r%�c)����;,�Sb�bh~�4;Gfz�D\hmڌ�x�YVu)NP�5�ͭm����]4k�(ƹ����%9)�������%�bX�}���r%�bX�g{�؇"X�%��o;v��bX�'�>��w2\mFᢷ�N�!y�^O���s��4/� d :�=U8�<P�%�b}��ٴ�Kı=���ݧ"X�%���o�iȟ��"X���=��W��9�
�t�zk�^���>���ND�,K�~���r%���b}����r%�bX�}���r%�bX���{�SX�Z9���rS���8X�{��iȖ%�b}����r%�bX�}���r%�`~��=��߳i��^��ק�߷}��$�p�Q���%�bX�}��6��bX�'�w�6��bX�'���6��bX�'�����wy�^B�~����85�H錘�7l��d�WnP�x!�g2�jīLի�����{��,y�	�e;���%9)��w�ӑ,K��;��ӑ,K��߷��U9ı,O��}�ND�,K9<��}>��,��T�ι;���/!��{�NC���,O��s�m9ı,N���6��bX�'�}�N@$�%9)�|�ٴؿ�a�4u��'�,K���}�ͧ"X�%���o�iȖ:y���le#`�`�H�d�R$  @���
G��DȞ}���r%�bX��~�m��B�����~��Mj;(�G;iȖ%����o�iȖ%�by�{�iȖ%�by��siȖ%��X�=�}�ٴ�Kı;���8kV�̗Yn�kZ�ND�,Kϻ�ND�,K�;��ӑ,K���}�ͧ"X�%���o�iȖ%�b~G�v�!�����\����'	mˊ��ͮh�)�	�)�c�A���Y	�j��i���D�,K���ٴ�Kı<���nӑ,K��߷ٱyı,O>��ι;���/!yޗߦ�\B�9J�iȖ%�b{���ݧ �%�b}����r%�bX�}�xm9ı,O3�w6���@b�"X��?_��ff��Ւ\�5���r%�bX����6��bX�'�}�ND�ı<����r%�bX����fӑ,K��{�˘�N�I���u���K�Ͼ��"X�%��w��ӑ,K��߮�6��bX>|��S�'ț��}z��������_	��6��P�h�r%�bX�g~�m9ı,O}��iȖ%�b}����r%�bX�}���r%�bX��S߿^e��̙O��Bm`��,h�A�m�Wknu�Ix�QvC%�4[)�Hy�{d.�u"a=��zk�D�=����ӑ,K���ٴ�Kı=���yı,O3��m9�����~��v�v���u���"X�'�}�ͧ 6%�b{�{�iȖ%�by��siȖ%�by�׼6���P"DȖ'��sZ��\�u��f����Kı=���6��bX�'���6��c�`DȞ����ӑ,K��{��iȖ%�b}ߡ�亘]K�3XMf��iȖ%�6'���6��bX�'�����Kı>���m9ı,O~�xm9ı,K���3ZM���R��rwy�^B�~�߷s�N�X�%��}��6��bX�'�w�6��bX�'���6��bX�&��]��.qt���G�ZL�qM�VT �3j,@-�A��WU����a;n��٨���CB�FV^.Z��<��[�91��Nta��i�����Vd�bm���:]ح{r�7/n^5�r�^��xZy[����4�.}�c��.���4p\Xĺ(E|V��54nQ=�nZ�25�x(Qs���
¿���Fʁi(��g;b��s����z�\oҩ�)V{V�9���{UQ��9�'f<�%Sb�cj�h��9ޚ��V9 �<+�6��bX�'�w�ӑ,K�����ӑ,K��;���yı,O=�s�ӑ,K��{�˘�N�I���5���Kı>����A�,K��{�ND�,K�~�56��bX�'�}�ͧ"*dK�>���4Xf�nk-�Ѵ�Kı=�߿fӑ,K��߷ܻND�Fı>���m9ı,O~�xm9ı,N�vL�&j�55f˚ͧ"X�
X�����iȖ%�b}����r%�bX�����r%�`~AD�D�_�~ͧ"X�0��O����6(�g��:�����b}����r%�bX"{�{�iȖ%�by��siȖ%�b{���]�"[�^B�}�r������#5;"Za&s��7V֋�$�9[�1�l�]Mu3.d��u.����Kı=����Kı<�����Kı=���.�^D�,K��fӑ,K���g{�M�2J�g\��B������}�NCb�����I�B�|x�*ƕ5�ȊH�Z������#$�%�1�9%Z��6 >���,Mk_���r%�bX�~���iȖ%�b{�{�iȠX�%�ﺿt�֦�f�3Z֬�k6��bX�'��zfӑ,K���ٴ�K¬Uș����iȖ%�b{��~ͧ"X�%�{����J���.Vn�|9)�NJr{��w�"X�%�����"X�%��w�ͧ"X�؞���ND�,K��{n�pA3L�y>��%9>���ɴ�Kİ��{�ND�,K���3iȖ%�b}����r%�bX��=�)֦�kg�k6���1��D��H��<��Y:�A�����%�{�����(5��4m9ı,O3��m9ı,Os��ͧ"X�%���o�`�%�bX�����r%�bX��{�S2�2j���\�m9ı,Os��ͧ"X�%���o�iȖ%�b{����Kı<�����O�ș������fe��"���'w����/'�}��듸�%�b{����K �#��IH��a�vĆB��80tG���ߤZf�ܴ	&�	Y�+$�)�53!�A�6A����Q.�������V���"�"S�g��jKBĢ[�綁=4��ل�9�� l�[`�B��e��0����Q�Ɛ�8�ɹ�t�`�ff$��Ó��2D��s���$&c3Z��%�0�6f��d$')NR!&�as�8>M�ļ��GN���ۡ�#��r���9$!L�zG�oDiٳy���֭#Yii�6UB4wˆB�xy��2�@���.�	j�d�(Fh�u��&����rRe2C�$�Ԟ�>�ۭB$�эL�"m"c�����"A! BM;�[�f�l��惇/.���%Ԅvy&��I\c�����B,��	���pF��D���Z��f ��|��!����u� UB%8�E~@q ��mSz�	�ãbdNf��6��bX�'s��ND�,Kߥ��Ƹ�\�4V����/!d�O~��6��bX�'���6��bX�'��zfӑ,K���ٴ�Kķ�ߧ���GJ�ul��:������'���6��bX��}ޙ��Kı>���m9��2&D����iȖ%�bx������f9L���je�3E� ���\�Q�%%�S��=:�c�'c�7-8"�*����צ�5��~����r%�bX�}��6��bX�'�w�6�'�2%�b{��~ͧ"X�%�|_�,���˕���JrS������6��bX�'�w�6��bX�'���6��bX�'��zfӑ,K����f����o\��B��������r%�bX�w]��r%��Dȟg~3iȖ%�bw����K�������x�1�g\��B�����nӑ,K��>�L�r%�bX�}��6��bXa�H��H��m�����"X������ji��̃�n��'w���%��}ޙ��Kı~���m9ı,O{��6��bX�'}�{v��c)�NO�$����!��e�WKu��5��h+�[��#�Κ(J�"�մ'�G�/v��nȫU�����%9?�~���Kı=����r%�bX��]���bX�'��zfӑ,K��J}C� ��Eo\��B����}��6��bX�'}�{v��bX�'��zfӑ,K���o�iȅ�bX�u�ye��F��&�����Kı<�����Kı>���6��b�%���o�iȖ%�b}߷ٴ�Kĳ�ϩ��ښ;m����'Ò����H�D�w�ND�,K���M�"X�%��~�fӑ,K��;��ӑ-�/!y���lʦ:V,�rwxX�%���o�iȖ%�a����y�m<�bX�'�����r%�bX�g~�ND�,K��'�ޙ�a2/����eGGKl�l����oWl�ݗ
���/V�E���܏A�nmvͧ
\FZ�q�3�K+j4�88z����y�ĝ:T�v�-qظ�:1�l0�َ(4:�ds��q�=ez�'V����{QU�\�m��Ӱ��OX��KJm��h��I<��yts�u�V�kf�e`fd�[� �@�<f^���+�V|ۏ�p��ՙ�d����Ch'���5�G����:3����Rs=s���i�$��#��9����cO�p���ɥ��c5fkSi�Kı=����"X�%��w�ͧ"X�%��}ޙ��Kı>���m9ı,O=ՇN��չsZ�sFӑ,K��;��Ӑ@�,K���3iȖ%�b}����r%�bX�����r"6%�bw=�r\3.h�Z�Y3Yu��r%�bX����M�"X�%���o�iȖ?�`��2'����ӑ,K��?w�m9ı,O����5Uso\��B�������6��bX�'�w�6��bX�'�߻�ND�,DlO~�y&ӑ,K�O=�S�� fn+z������O~�xm9ı,|�����Kı=���ND�,K��fӑ,K9���K���c�p�њE��OU����n�#�T��%���ך;3��5�kFӑ,K���nӑ,K�����m9ı,O��}�END�,K�~��"X�%�纟t��ְ��33Y���]�"X�%��w�m9
W��-�T���v���Q,K�<�fӑ,K�����ӑ,K���nӑ,KĽ�iw�]�bJ�m�;���/!y=�޻6��bX�'���ND��,O;��v��bX�'��ӛND�,K�����Dl��N�|9)�BHH�'���&��	�s�݉ �'<��I�$����o�iȖ%�by�:t�)S-�3��JrS���~}�{��%�bX�{�Nm9ı,O��}�ND�,K�~��"X�%��d�NWZ�ᯱ�x�fz1X��E% �,u�xwbt��\܀����'t���yuJ4��%�bX����6��bX�'�}�ͧ"X�%��w��yı,O;��:��������y���m�٪��[ND�,K��fӑ,K����iȖ%�by�w�iȖ%�by��9�� ,K������Vۆ�eԺ֦ӑ,K����iȖ%�by�w�iȖ<i�H=p蘩�G�2&D�{���Kı<����Kı=���۫�2��I��ND�,K�뽻ND�,K�~��iȖ%�b}���ӑ,KlO=�xm9ı,O����a��!����f�sWiȖ%�b{��8m9ı,����r%�bX�}���r%�bX�w]��r%�bX���9z�d6TJ2z^-3�Y閘K0�@�����R�-��x�ӳ�\%81�z7�^<�bX�'��xm9ı,O>�xm9ı,O����?�D�&D�,O�����Kı?g㿌��,�jj��nh�r%�bX�}���r"�bX�w]��r%�bX������&D�,N���ND�,Kߵa����f�n�kV�Ѵ�Kı>���r%�bX����ND�,K���ND�,KϾ��"X�%���{5��DA����|9)�I�r��~����r%�bX�{���r%�bX�}�xm9İ<�����"}��˴�K9�^O���)��6j�Q�rwy�%�����"X�%��}�xm9ı,O{��v��bX�'��o�"X�%��vB\d���3)�$��X���ٰB��f��(W$u�9�LM4� _t�=.��J,�]��'w����/'�}��iȖ%�by�}۴�Kı<�{xl?�<��,K�w��"X�%������[��a�5	3ZѴ�Kı<���r��dL�b{����iȖ%�bw����Kı>����r'�T�"X��S��a�S)�����j�ӑ,K���߯�"X�%���w�ӑ,K�����ӑ,K���nӑ,K��>��;��0��4ɬ�6��bY�9��ӑ,K���w�ӑ,K��;��ӑ,K�
C"}�߯�ӑ,K���P��.��L55sW.h�r%�bX�{���r%�bX~����ٴ�%�bX�w���iȖ%�b}����Kı<jm>\�
�
� @�&bB2K'��{���e.�MV�BX�g�K�L������2ޘ��K���sy{V���l�M�)[	cR�M(�#h]�%�
B���עJ���� �冻%Xj1��-e�el@�A����H q�.t�i�n�vvٝJ%�!e��@�<����;q�n�@ܗaA�4�l̽qڏa�iw"�1k�ts9�G5�cT#��K��瞸�c�n ���Pu�M>����HO�w|�}+���37Uf�sֆf��n��%8��)�MH,bࡆ#F\Q��$��1,f���5�nh���bX�'s�߳iȖ%�b{�{xm9ı,O���6��bX�'���6��bX�'s߻���5f�ɩ5�WY��r%�bX����NC��ș��߿p�r%�bX����ND�,K���ͧ"X�%����x�E6j�Q�rwy�^B�{�w6��bX�'���6��bX�'�߻�ND�,K߻��iȖ%�b}���K�l�h˩��ND�,�{�ND�,K���ͧ"X�%���M�m9İ?+�����ӑ,K����,�Y$�E�&\֍�"X�%��w�ͧ"X�%���M�m9ı,O���6��bX�'���6��bX���{����\KB�pn7B�qx�\Ŭ�g2�v�v��\�v�\Q�������y,mˬ֦�Y��Kı=��ͧ"X�%���w�ӑ,K�������<��,K����m9ı,Os������a[�i����r%�bX�}�xm9�H��z'D�q2%�bw\��"X�%��w��ӑ,K���xm9ı,N�P�f]C,�jj��Ѵ�Kı<����Kı<�����Kș���xm9ı,K������bX�'��N�3E����֥��iȖ%�X�g{��r%�bX����ND�,K����ӑ,K�>����Kı;���Y�K�&�MI����fӑ,K������r%�bX~D�~����,K�����iȖ%�by�����Kı>�N�JL]ﳡv�f��)��ᬻY��vW�z+�tc�� ŧc;��ot�"l��ˣiȖ%�b}�{�iȖ%�b}����Kı=���r%�bX�}��ND�,K�^�g5	m�L355sFӑ,K��߻�iȖ%�b{�}۴�Kı<���6��bX�'���6��bX�'�u�K-�Bf�]Bf�Z6��bX�'��ݻND�,K�{��iȖ?�< �RF��H�)�E`� �A	�	ŀ,ND�߿p�r%�bX��}��ӑ,K����6��0�L�rwy�_�K'5���߯�ӑ,K��߿p�r%�bX�}�xm9İ?"}����ND�,K9>���T.��#��rwy�^B����6��bX�+���6��bX�'�߻�ND�,K���iȖ%�^O�{:�pf�Y�9�L�#�0���<"6xn��ţ��ZCb%
ի���t|��S6���֮fh�r%�bX��{�iȖ%�by�����Kı=�n�6��bX�'�}�ND�,K�����f���5���6��bX�'���6��� DȖ'߿]��ND�,K����ӑ,K��{�ND�,K��׺قD�mڣ��'w����/'�|u��r%�bX�w���KʄUș��~��Kı;��~ͧ"X�0���=�{M��] [�'w���,O����r%�bX�w���Kı>�����K��pv5J;h�W�A,"U�S��{"^j�iȖ%�b}���s�5&[��˩.�m9ı,O����r%�bX~(���߳i�Kı>���iȖ%�b}߻�iȖ%�b{��ɷ���x��l�qq�+��b�U��/Nڮ@�g=s6F�rz�`��9�fk���bX�'�߻�ND�,K���iȖ%�b}߻�j��bX�'~��ι;���/!y=����h�֡�-�k6��bX�'���fӑBı,O��xm9ı,N����r%�bX�g~�m9�S"X�a��~��Y�X�i�]jm9ı,N���ND�,K�w�6��`�b}�����Kı>�n�6��bX�'{�w�.�a�&����Ѵ�K��2'�����Kı=����ND�,K���iȖ%��'{���r%�bX���>3�h�SWY����ND�,K���6��bX�'���fӑ,K��{�ND�,K��xm9ı,O�{$`A`D"E$F@������������Ca1M�����4�i����	 p�;�X���J! �A��] G"�"���p��0$�F)���H�2B��}��<�$��Þ8W\��H�,ިL�L��x������3��,�g���Y��l">���"�j� l��X���*� UUc*��UV�UT耨�V�]<�$9�F�۳�:nw�j-�9�q7;�tp�L]c�z�2,n�\n��]x�y��R�!��`"��ƍz��Ҏ���WV�d�:�!Ӛ�p��h4����N2������u��n:��s6 ��-��i��#B]4^G����Y9\{kI+�ز����@n���+���WDƭ���א�gۂ�.R-��r���,���x�-Y��F*�d��b�Ga��l�
��Ҳ����@I���6^^�$�iu��a�=�y��C�<vM�jL5�f��ۉ,3ۑ8�q�a
�.�3�����v�!`ZJ%m��D����X-�Ôر��XA�`Һ�
ZR�iS1�V�f�g�aӛ"e�����yGs�cN��&W��.c�f�H�֤��@��e�K���6�13vm�FBj�JԘ�3�6VX�W��5cd���Q�zS���c����.�ie���n�Χt{o�#�z��@TcL�6і�F٩�Lq�n L6�{�I��.ރ��n�X�t�6#��Z
���:-�d��&�۱xb�	�۷pZ�ۧ$�Y�,�`4��Q���9�l���3�W���k��>�8�=e�8���g�&����K�6�tv�C��{5��>�m���mqp��>Ma'Ji#gul��P�q���0��vǱ�Ew��T�il)Lb�*B�H��5�%����2MR��n��e����Pe�G�I:.r#�0����T�R�8%�m�����eRV�<ΩZ���@]���%�3��j�g��W�7[�c��^�a������+�lZ��n3��z�z�1��r�Y���;
��00�3ϭ�T��9w
�ۛ[����2nDb�y�[&�	��g��Zw&2�-S��h7J"�7L�Xp�2��l^�K�*yg%��)���������j�jM���P#���Yh�B���d&����"^g:qˑ@����pD�E*&����
!�}P�-
�TDW��P|��<���ꠅ@�D�#�h`pO9$�c�F��k���կ,�mt�nh�uu�W�m�-�X���8�l�R�s�xn&�Vf���bU�f�%�ɢ��{B�ĥ������"c����z���S����g�G$4��n�XQ��0k[m�W4hJ[`٘�,B�sx�x�G9�����j�]�c��He���9�Ѷ�C
0JKe���3-�͗v˃���KP�k��1���䓖s�g'}��1�\v�JqO�������_lݓ�MX����u�0-��$��z���1�k��OJrS���}���iȖ%�bw���"X�%����6��>DȖ%��?~��ND���ק��~�����O���bX�}�xm9ı,N����Kı<�����Kı=�n�6�����2%�����y��F\ɬ2�]f��"X�%�����6��bX�%��bX�'���fӑ,K���w�ӑ,K����i-ә5�5�֍�"X� ؗ����r%�bX����nӑ,K���w�ӑ,K,O����r%�bX�{�}�3Lѭ[5u�ɬ�m9ı,Os��u��Kı;����Kı>����r%�bX��{��r%�bX�������$�"�s1wR-�ƍ�^]tj����m��v�<Qt�>�����X��}���%��~��"X�%�߾�fӑ,K��{�sa�Q'�2%�b{�W���O���5�O����KP�#��g��Kı;����r >H�� ��>8��M��O"X�&g��6��bX�'����iȖ%�b{߻�iȖ%�b|}��:曭e��je֦ӑ,K��=�siȖ%�byٮ��9����w�ӑ,K���o�iȖ%�b}���k$ceGv
dOt�zk�_��^��}��6��bX�'߻��ӑ,K���o�iȖ%��'��{�ND�,K�����LX�f�z����������iȖ%�`~�}�ND�,K��{��"X�%�|��u��-�zN���ڡl&�i�,3R6Ce����Dv�l�.�[�Vմbʷ-+ 6i����?�L��)�������l'�~��7�^���'�զ��l�7�eg���H&���7��X�p��URGv���M���CNݻn�o�<�fV�t%����A��߿}���=�߶n]P�m�N�*ۧV����R�Or�	��`�2�?}U�SҼ�	��[T�j���M��\0�US}�W '�y��X�P����I]�tƋ�mp���`�-*V�68�!��O1��\I����l�&�5m�M�{��j<��+�}�OG� ճ��:e����0f�y����ٳ��߼�{���=^˲�����-�����e`5����n�� '�y�Q ��v+EӴ���X��ꯔ���~��O~�����rHJX�\! F����"E�����x�* ~�����y����	�������0�\0{"x;&V�8`��[>�����Ѐ�u|���f]�}6\�Hm�(�V��RTmv1U��T��.>���̡�i�iڻl����x;&V�8`�`uB]��:_+�]�c�9�2���_��������R��������%�I�jݵ$�`k��ɕ�睊#����7}��/�ʷI�I�6��`�X�x{&V����3��e�:YCgή�i��H��;�2�	5� �d��3�w���{uCVQ3�d�f]�l�G�`3"�W�4cq�f�i��Z�hK,�
�QX�%�A�P��-��b��(s���[�t�������\�{n�N��2mq��[���p�a-\U��wh�-�����/D�-f�R:�ֳ�V!��.v�b�6�S+]3�k=#n��h[��5!�&�l���kn9��͹p�7k��	v��ϓ���wI�ܒ>y��5�e�ٳ�⡵��BGu�-ͦ�G��-At�)����k�s����
�}l�V�\0͙_���������������v�itKZ�� �����{+ ;�z��ɕ��#������Ƈt�`��V rIo	��n�L�� 9�������]�+��.l���{+ �0�L�.�Gm��K�v¬m7�w�e`�zg���e`6Kx:@Nұ+�������F��m6v��`�,5���Rlj�Eu%�Ɣ��i�S��v���u�l�;&V sd���v�O~��6�z�2��n�a������o��E��D�
 �p3$��~�����7$��u���~��Z�������uv6�� ����9ݙX�p�9ݙXt�1][N����ݢ�o�U}K�=��7���;ݙX͊<J6.�;-Zi��u�l��ٕ�أ�9�2�n�vRxr`��?\����0�sF�ڍ��c5Ѭ*�Pmo-#�yrf��[��t�fV sb� �d��$����C�:v��iڵn��(���|�����/O^����$E�ů6��|��U���ｕ�lxr���PW���H�D�)$ �J [(��i���UWҚ�L���Q�,�Z����ݵt��`͏ �ve`6(�=K��r��J�;L�2��V�����MQ��X;#�;йQ
�[�?����Ϯs؂��$�s��f���]���srDՀ��\�y��!63V| ����s�e`�G�w�2���eյvU�v����vL������<v{+ 9أ�$�bK�+V�-7wn�{#�;ݙX���ɕ�w�l�]Ran��m��ٕ��Q�'<�훓�5B ,"Ğ
I�;������{�f�]u�`;x�����{��	���;�2����Y�&��Sk��(J� ����sI	�t��mY��qӧWk�+�m!ٙ�Ǉl*�i���+ ;��ɕ��G�j�"����W�M� n�x{&V�� �d��%*�ԧi�N��wi�x{&V oI�ɕ�un��:��t:�cT®�i���Q��X��x��]��V�%x�c�������i��ٕ�}R�����V ob� �~��(�>�ꪭd(�-pʾ�L��i�m[��f��#�ܻT�s]g$�D�B�6k�m�ׄ����]n��C��!��sz�Nn\n��l���q�;K��''�F �b3=�ד�y
�%��9T�s����P+���PҢr5���t�44���T3
�m Ԝgq��Nݍv�Pd�*׷XG2˗��$b����pC�)Ղ�cN+��bh�u�f�`��S橿<vL����Y���\T��X���W���n�)KӍ�2�r�{8���qn���ٞ���w@�d���Q����۞X��� ˪T�Ӻi7x;&V~��� ���n���5n���URGey��I4�CM+�X7�� �ob�5n��9�2�-P-F�]/��e����ŀjݗ�w�e`�(�R�V�Hۻw+��]�x{&V w�G�w�"�o��y��v�if�.��Ä̡�Զ��R���ɝ&�L�mZF�1�#�ۼ��+ 7�G�w�"�5n��:����i�ƺl՝ ��׾Nri1T~X���$�YF1�2I H�+��	BK��ϫ�U}�9v��5we��Xa�/-��Ci�.�V��9ۑ`�e��̬ ����PK);t�j�V��ٕ�أ�9��w�l��ݟ*t��4���ٕ�~���M����?��x����&xv��>[$pV��-:7��y��v률1B󀸸[jqQ��E��n�vìd��\ ��� �c��UU}���XT^^����N�U���v8`n��;ݙ^�zz�=g��S�;�n��![0����fV�����Eĉ�7�4��B^x%N.EB�X�����I8H�aH%�12�բ�]a+
��wX1CW0_�B&�xQ߄`��9EK4G��;0�C|�@ַ��� /��`����d\�嬈����p�'$�� ��Q�e�]Mz$�s|���k�`�OQ�G�&a�\���+In��H����-��HF����i�� IS�;��!��]xfp�\�a$�)&wNh�@�d	�,a
B�)Y���q5��*K�8+�I�)��;V�� �"�b(pAu
�h����'��_�C�G�#�x�Gh��s�,G@C,�ט�	#��/�Wc�v[)�m��;ݙX�Kx;0�%�[��b_[�P��n�d��Uw_����׀w�2�l�WIZH��]*����Ŷ�sԔ�Ƭ=6Nu�:P�-7F&�������V�v�MSwbB�o�wo�X]���fW��@I�[�'���ST]_�wb�k ��/?�����#v{+ $����ȳ�$w~��Ҥ7bwM&� ݞ���G�s�"�:�K�9*8RV�һb-6��X��)y������f��*D DdV �`�de!I�$! րx#�$��}��_/٬�gSr�	����Ȱ]�x{�+ 7�[�9�L�&n^\g&X�1�Z �B�t�5��B%x��4�ѕ���"~�;ϱM���F��[=x{�+ 7�[�9ۑ`����X�N�e;-ۼ�ٕ���H&������ �ݗ����5Ik͂*��
�� ��^V�܋�_%�^�=���;�z��-cwV��7Xv��jݗ�w�2�=��_~������X����˻t؉vnV��Ͼ���{����'����rNy��w$��_��<+��tF"h���*�J�8���S���ƷR�k�/W��[J%U���������$u."P�UX�2a��rs�_K�軎��;d�Uэ��ˡ���t ���d Ҩ��=`3j��k��ܛ�*��]��l'�V��c���c�8dEܽ�4����@{d��ur�n|��I�`޺q;�N��unp�����B�	Kk4D�(j��xJ1!oRۮ�-Ҫ���t��?]��I	' �P�Q�^.X6cM�]q��])�9��+�(\!�A�,s>��B�����m$�V�I�vK��;�ؿ}\�N�}<��շϧ�ԦcM�TSl�����;�ذ��x7fV{���rs�_~��%76�gV�>�P�엇ﾪIvOr�����;�⫲�5v�T�m`~�ﾥ��׀vOe`ݗ��sob�9�R�c��-����ݙX������+�v\��5l��y��u.�4�57��.e��u��%�S��e���ǳ5�H�IC��Ra2��X"�۬t�+ ��ŀul����;#�n�U��ڴ&����v��ͽ��J���!P���H(��� +B+�-ń�ma"�1���ih�F(��2	��+���}��3�3׀n�� ݒ��ة^P�.wb����^��=��II�^V�s� ��"`Pݗi���j��~��]�<`{ו�sob��_R����7���
�1]�6��`�^V����sˀyzz�	�2��+�v���v��M�6�����f;r���;���Z�(�6f�ج>�m���`ob�5vK�'d��_WI�^V7ɞ�)ի��v*e���Ȱ	�2��/+ �{{�H＝x�h��H�m`�{+ ݒ򰯗�W�W�`"T����rO|Ͼ��r���t���lT+V��}T�����z\��7��`�e`tT�m+B�]Z�v� �{�����ypo���obp�9(�%R��ZJ��]:�Q�%� `U����x:�)���s(�+�Z��]ح��n�ŀNɕ�obp�&�ŀM�D��N����	�2��RD�'� �\��7ob�;��B��wlV��&�`؜0�ذ��I~��&��X�Stҿ�l>v�0�ذۑ`�2�'�]*��*@����$l�!$)p&`K$h@��hHF��H$$L�0�cXؤBaK-KhBH�%i
��j�U�D��RH��a!B��P�,� SLK����mK���- ��T]$&��R�����].v�i��=��^��V���ب� ݽ� ����\o��l�����=�����Bq�9�r���s,�/,%�\�l1�hİ�
��)]aV�
�ء�ce� ����؜0���I~��<����%M�بV�۬v'f�`�"�6l���߾���͓����T��~��`[������7'��*��N�V�e��V�v�Xd�X�N�'���)�؋m�T��;$��7bp�7c��s�%��E
��?y=��nb�˄���g��000,g�b�u�َƲ��/9n�;�; ���Ú��m�4o&�D5�b\����5��xfqYᬁP��,�Z��,E��Iv�N�ܼ խ˝�)�8�D��o3 ���!�˶�x�v�Z��*3o�;���n:)b��Wd��'�����Vm�6�֞�p�b��M�y�q�u�[�7F���b	t!�������I�m1n&��)�[�Z�:��dk�`�uv�ۙ�^�sV1֛
B���˔��unJ��=���v8`�"�;$��'b�.��j�����i� ݎ�Ȱ�2�؜3�U}��|�K�M
�X�l�$�y`�ea��JC��'��dN�;-�i�2��m`{꯾����X���v8`ۑ`M���6�B�i��6D�l�[%�$��<��� 1[�CJ���^H�u�wt����n	���X�����4��N�M�ڻV�=�� �d�d�XȜ0i%�yM�utʻ��rO������4D��Y�sf����vGwi�;�N��TZ�x�X�Nz���-�~0)=x;{��)ݱZj�������0�~0[���Xؠ��-�/��;M�v8`���~���߿e`=�����N~翾`�M�1��7mǵ�85C� M�q��b�`tkk��y�tm�6�6�ڶ�]�t�z��X$p�;�� �e���&��v� ٳ+?}�$w�~0	��`�"�"�\n���m]�Xdp�7�� |"���S4Pa��$
%9S��P��DKj츦F˳�bf�(�"zsC�������}��ܓ�}�Tڎ�,��[�$�=�[|7޼�fV�ɕ�wM�e�`�]�
ـuwe���UT��ݮ����{0݊�W��WH�k.�R�aØ�Yͮ��v�s �u�]U�	�t�\&��WIۻJ�V� �ٕ�s�e`��{�v[��n��}���s�viW.VuC��+?}UI��,V�^����W���$zyxF]Ze�`ӷX��,��/�%����ｕ�I�����Wm�w����ŀs�e`�X����h+C��L���	mҌo���.����k%ֲ�]��˻k �d��9�2���,���ށ��}���G�6�;yE�ⲅ�熳�S�ѻs�7<�W-�=.�K���MYwm��wg��v�Xv^����&�8�WI�t�]�۬�����:�z��fV����%M%�m5i][Uwb���ݗ�w�2����]���~��&�Qbhv6Z�x68`�̬�{�꯫���~�~�W�!�T�؆�v��ٕ�wob�8���lp�:�U\���QUA�C�Ar��Wٔ��!��<d$��i�}����&��a=��	��!	e%e$��j>�x���	mf�1�d'�I����L4�6��ꇑ|�##YhP�HNCd
g&�F B������Ϡ��Rxh���-�P8�B	�H0`ɢd��Fa�}�i8�_�q,���3��2Y$|����17���H�������F��F�s�p��$LaHC�C�d籁��Fpn��@��@���CG�q�da��!�ߏ<MK�M���ty@����0$�D�&ɱMs�{!3-��ľ6/���Q B1������$��Ԓ솛-8z|f�h���aH��F���xL��BBB@��k�����k*q�Lḻ��Իi
S0�9e7p�F@���JR���z���8�K��Z%]<\I��oA�s�C|��[���z�_=����#'��=��H��� ]oZ>����	׾���1ظp�2}O����������(h4�0��۳��UTZ�X�j�
��J�UU�X��N�]UUUUP83j�[�K��\nZ�RGg&YT^3�&�kt�[nÚ ���`�m*(˵�[B)e0!�DQS��v���WN����d2֩�"5ǞΞ)�
�4�n�����Lq4X1-l���Cp�HbAK42�9�, d*�t��X��Y��ɦ�JE�(K;v�*}�1�*�ۮ�yf��8�h�q(����RB˘���xA�«�Q�]<i�5E�e:ѵ��:��5�y2nys�糆n�]��q<�/cL�%O6�m��`��Ub�̰��k�$�5��d���ݧ;M�'E�"\l/C��m��IzD6�G���h^�c2`ym娒�aPt��D�G�c�-ٸR�v.L�ذ�K��ծ�eer��i,�ȺÃrn���	�`�����' ���l�txNG��5�H8.vz��%�u�Z�XFÞr��u�,�X��s�u��m���5�#n	D`��i[
s�DK,R��ٔv�ؖ<;+�{���,cv���Kg��y|"���Dv�7m���������B)g[���)����n4K�l�l��v�7��c�����б]�ݨ4yRӄ��({.�-�����W;G�BV���w�͵�f�E&�T<R;��TQ�*r�������w;G;�Xk��O%:��W@H2��Q��n�����.T���<px�蠏"M52��Y�A��d�p��8·���� ^n���c��V�Ѝ�W]8�v0��J�P��d���t��Q��ez��*99��q�)�wc�稽�����r�L�R�r�[
<L�鳬��)1-Λ�4�D�554"�#���^nP�@��R�e�˱��)+0� Bڬm��36�mq��b�0�m�;gb�*��kX��m]ipr�,i�(V��%��X��Ն��Ƶh8;)a*�ic�2a�=,s�1��3%�hV�d�3a�j�1�ea�����d�A�lp�3[0�@W��H �
���>D�Pڊz��t b�H� V����<��qU �C��}<�,��%A�Sk��Ip��sk�a�Ób��Zq����Zے��Z�H��Aʭ�b��Ʋ�d��#�=l�*A��ga�v*V:����ڐ�ʉfJD��z��L�x�9&�*T����)�`q�2�z÷q7�rێ�1��2�tM<ݥ�:�˫i
N��<x��(�p�]:�V7�d��{g���������).r�0���ӿ$�B{bbR�>���n[�;5�M;���Ѓ�Q�Z���0ѕ�j�c�Hi�g���W}�ݹ�ݗ�sc��������~�N��NݗM���-��qwe���s�2���Y�H�D��:�����Պ����� �vea��-�<������Wq�U����]�v�R��r��<�.��0	�$8�+���5Wcm�ݽ� �UW�}����;<�`Ny��7$����ɖ�!l�&���^���9�a�`���/mz� ,�,�A ��ʔ
��ݷbh���ݥm�ݞ��9#������_Uq�<�OR�2��]'bd$���'>�_M��� l �-Tc7��7��`�g�$���[�N�n�wl�;��X��X;�$p�&�$eկ�_��4��v�,��$p��W˳��`؝/Zv��ڻo��Xw\0�W���� ���um���V߼��o�DlP�-�#CT��hK�I�HY���,΃kH@U�j%���݋������uav΁��?�͓+ ݽ���W�Wl��ݿ"��Ћ�l�Wv]� ����;��`�`�៫ꤏH$׆���cUv6�`.v�I��鹂(@�f�Љ�
�d]E�
F"�kH�T�?<��`�e`����mV�;�[k�}_Rݙ� ���s�e`z�U_����ߨ��b���S�:(u�rG��+ ջ/ �ve`���wV��ةY�]�e�#%��<�k��	p-!���؎(��&�H�uդ�dp���ۻ�e`�e��_�� ���x��$eة���Ӣݺ�5n��W�Wԑ7���:��^ٳ+ ��d�ai��7x�L��Ix{&V�v^�.�D��C����u�qI/ �va�'��~��ψ������>ٹ'<ϩq�uv�]v���;ݙX��x�̬�IxݧV�v�j�]�w�-�p�s9`2��]Υڤ�����v�����ւ�Z`��X�]�m� �O^;�+ �_�{g�����x��m]]�;�v���2�)%��2�[�������y�~��L���n�_�~�wfV��J)=xw���7nJH�j���ӻt���w�2�[��vL� ��I˻W��CM��v^﻾�+�����fV U|���ӪGM� �]5�ˊ�Z�2&���YU�pۺ�k^Bm32���f!��\���aB��`�ZЊ� ���h7�cL�B�x�f	��M�a2]b�U�k5ͨ�OsƸ��㓍�dsω������Hmй/k��[1��OW:vy�v��n�e9w�u3e�"�Xխ�8�����z��Z<���V�H个���7X4"�U(:ܣ���|��MB�a������#;\b�07ny��<��*=n����ٹ&��mUi�+�������ﲰ�G�w�2���"�׀l/��髦:v7VZn��G�wd��5n��}����������M�F�M��hk��6{�X��x~����e`^�� ���ձ%cUv�X��xvL��Ix����`��z�۴�We1�ڶ�ݓ+ ��/ �ɕ�ݏ-�ܟ{*X�}��Ц�,��f�V���&��z�-��"��<�+��쐒s�Rt|	��g���̬ ��������=/ޤ�MS�j�;��n��̬�M�@���F�V+B@$"A�5�Y<��krO<�_M�'=�<Wd��v���j��I��ݏ �������Uޯ~�x�ߞ7]�t�N��ۧV�o �ob�8�K�nǀݏ �.QM_��Cue�k ����.����� ��ŀw��<<
e���l]�+�CP�,ְ����K��0,%νD�7����p��5��Yv^sl�nǀݏ ��ŀsc�;���:��cUw�o ;�{���;#�vy��nǀr�*]崛B���ڶ�ͽ� ��.�:������}Ͼ�8E�I"0���? �B������e�y�=<����ueզ�K��ꪪ]��'������"�&܉%ucv�iݴ�ـ$x����"�9�� �b�x�l�'!sW%�`���Ҽ)�Em�g�@�̮�v��#5��3Qo�'���X68`�٬��s�)��^��{�����'6�}~������"i{D��:n�V����� �#��ǀj�^����i��m1�t?���߿= �<�RK��ﾪ�UUV}U�_fd0	�Hq�t�j��Wm�wc�5I/ �� �#�9�'�&6��QBv�&1�q���4뛦�+��_�q��)�6��3�c�ۻs�7qk�����۠sc� l��������� ݨ��n�+�������� 6H�wc�5I/?|��~=IZ)�M]�v�v� ��� n�x�%���J엊�v�K歂-�����<���^͎��������y]:v�JէN�&�ջ/ �� ��wc�9^^I���asn����EԮ�2�E�乳g��r)�VL\gv^�Yt�q��pi�R����aM/h:jYPc`3��[nX��l1��l<����ap�]�oE¦�[�ȴ嚴ѱ���:[/�`9�Du
B�R	��lW��p�L��e�nXą��R��.mMj��h��К�SR:^��`E����<u�V{�v�Y�qIQ+��$X;���$�I:��0@,5�7����H��\��WlNuJ�C08���δu���e�j����ub�� ����< ���}_�}���=���6�˝�i���� wv< ��x68gꯪ�$��uc�cUv�o 6O< ��xz�}Uw��������ʊ�c%n�wv���ݏ �� ���������-]������sc��]�����un��;�����U�W?m7Z�GL;�\�r3�hu�
2sGnqR70p��Xݫ�]��>����ǀun��9�� �엖�4���Inf��$��~��!$Q�UJ1��SJx�f��w6�~0�#��$o���i[.�V���V��O^͎�#��ǁ|�w��14�Y�˺��rs���y��?��~x���[��v�q���[WE�Yv� ��wc�5n��9�� �U��*���4Ӡj��ei�+���#�^H�����%q)Nss�#)������7V�VӦ���O{��5we�����쨕��,���n�[o �ݗ�sc� rlx����RF���y5h�*�M��y��M�&�P�HD<�I�$!H�$�!2���
 A��B(��BBa��D}b�AtO�@�F��,	-�YP�)[Y6-4�a��aCFJ�'�GR,`Hb���H�bJCV����Ĕ��.k � �P�9ZW
k�# �u6�)��)vI##"��b`H'��-�%��"Y�@�HC(�g!�!�f� B@�F�p!��r'
X��i��{މe%�B62aAsE�Э����@��!	F}�)��|��E�!��H�e���n%-���%�a
���h�+m�����B��;��	K	aH$����T�"��Ę�%�XQ�Z��4%���&�BZnd�3R������HIKBT�!	���������!�	�!2��*�%!i
2�+k#+��ɪD�meid��Ér1X���Q%([	li�������Yb@K%�	,�-ɸ@$5Oࡂ!����D�|<@�N(��E��j����/P(�~@~Z��!�ڛ�o�u�'/�}��}�B$��I�Wiݴ�� 96< ���]�x�]���+�^�v�H_5lM� ���]�x$p�M��rOy���hnk�v/�ٕ��ֆ������@�6C�L�2V ��7�+k2(9K���m��z�H�������y�/�#Ν�]4:wWwm��3�_$���	'���/ �oQw�tՂ��n��c��Ǉ����;����=��n�جn�m�s�)�� �g� �ٕ��?�K�惘\
���b��Pd��$�{���g����k�������X����{���y��ǀsu{���̀�iK�m ���&]XS/-��3.l�,՜!��C�qu��i���7x6L�Wd� ��xT�x�����&ò*έ���u�9�mM��</��x��U_W��E�N��K�V�+���y�[���UU|�V�^ w���9*�ڿ����m�~�K�׀ul��$� 9ݏ ������bN����w�qI/ �K��|�O���ܓ�s߮�h*�B��4�ai,*�"�B@� y|���{;��F���V�� �)Ų��u�h2on.,�R�S��X�C5������9��6Dw5�d���PN��%8�[R\�)�4,щ��̧2bW)�Hf�\�
�M�kY��Ժ0�v�G<�"�z�u�H�t(���%j�0XW��gs����{]�Y���D\m��H��e��JcXj�*�h���4��GFfĦj[��4J�f�?:N��S��Ϟ�:��6X�R�$0�{k1]��g.'WT��=�ڝʙm�Y{*6�@$�x����ؿ����� ���?��I��7t6� w�ݽ� �엀��*A
򒴮�V�ն���Xd� �������g�i�D�r�uo�9�!�y�۪g�������XۄE]!'N��i�M� �������>�����ӫosُu�ㇸl�q�h���8�&��[k\]Nc0��Ѥ�ͩs�:��K��Cm�;��\� �����'9;-�}��V��M��L��vZ�3Zܓ���Dv�E(�AhGV�^ s�< �v<��Q\.��:m���.� �G��ǀIr,��E�V;��]+�ۼ}U������{��$���/ �&'�t��Lun��o ;ݏ ��Xd� �G��7g΅wj�]�+��%M[sضy����:�{P�j�]b�54���~�U�`�yIZWL�wj�|����`]��Iﾪ�vy���v�+�N��m���^z����H=�y�����}�������_��|�fW�g7$��{��'�{��8v @ 0�!�� I�0�F���$��X� �I$! HD�84kH�Q�JtE��*	{φ�z^�S�����!��=�W�|����=�?d� �#�;*�m_��ltҶ��� �엀$x��xۭ���7E]���d���;�J�^�^P;���|�me[�QA�X�Ѻ�
�SKVt��}� ������I2�WoQwՊ�-v�w��z��� ݞx}=��|�{���99%������Ǝ,Y�eo 7g�ɳ+ �엀ݏ ڐ�
��|��[o�}�|���Vս�nI=�ߵ��ɋ,� �q�e��YH�+�1��v���}�R-M�J���`]��{��{���e`�q�Wuh�|�%d���K�󚠬�uIٮ��;It�k���^x����2韶ݏ ;ݏ �+ �엀v��b�ݔ��[6� w��&V��/ 7v<��IN�۲��ltҶ�I2�.�xz���H�y����:��*�q���t�u�qvK�ݏ ;ݏ��W�R��V62�����.˻M��ݏ �U|�g� ��	���f�	�c�� �BPaE�B4	�Y�K4[rۙ��L�=�C^hj�����v[ Z�a���&�F�: QL.6I��}�/��sڃge+c��y�ؚjskT��m��KB�NBhC��O	[����Q�\�G4-ۊϚ��!����s�$��	��ru�>'jb��@au�� �WRY�N2�g��
����uj�^�9��V�6ՙc���kw�����6�lQ��m �w$'����f����J�QŷMT��ڃt�lp��[���-�ͤP�]�1�W�{N��#�B��-��| ��<�L���_��W�@I<�	^��Ic�c��m��L����W�[�^ I<����RF��t�뺴6]*v�u�qvK��ǀuwe��2��4��%n�v��ۼ ��x��x7fV��/ �i2ۻU��&�x��x7fV��/ 9���9��B�ڰ�n�%�1lnY�-Ј�x���s��J���-D�:2ᖨ�gUۗ�}����8�%�d� ;ݏ ����j6�	�SW)�>_=�w�y�y�NFND>�~= �v<v8g���H��E߁Չ�uwi�x��� w��0.�xf��7N�7ah�m�{���� �엁諭��-���	S�䅌H��wj�x�p�8�%�d� <��@��$矠Ҟ�)�;�Zק���[r\3��u�t�sیH�ȃ9�����.kt�]���*c�g ;���� w�+�7c�zGIҵv髴][�����9���;�p�vG�vjSt�X��[��o ����7c�G� �"���|����7�� w�<��j��t�v�t��x�p�8�%�d��og� ��҇�v�N��Ӷ���^���[�y�vy��� �oQt�
�Wj��(N��CGTX�e�]@�Z2�mѕv�$μRD�b#��V$�E�ݦ��d� ����6G��/ ٪����R7alm���ǀl�v^ l�羯��%zH�iR�V1�ڶ�=�� 9ݏ 6H������:QZ�$�S�`]�x�G��ǁ�����{��MM����V�?_��̦�ڭ� vH�.�v8`;����{�5֛k��n��Qt q�f���t��[����T�N�EK,��us�8m�6������ 9�?W���q����Y.�Vպ��LV��0���d� 9���ilI�t��h�� 9� vH������ ��V���ڲ����� sv<v8`7c�;5Rj캔�M�[m��c�7c� rlx�>�䞜�F$#@�V�	P%�B6[F$�$�0$�+$,�T�0&̹��zp�a|�ƃ[��IP�:o�}&sn��wT�H�C���uֵ��z�>	<���.��'!f:6Z�&y�<ǟ���
�+KI�9�S�*�a�M�C�]�	�� R@b،�d�B1*R�X�mX�Ȱ�[�$>O>Y�	��K�K=a��ni�\����m��bOL�G��	���Rh��yl��M;�=��@	��Ӳ;��0�kq$0�+��{�ٚ��I�r��a�y�Zn:Dd�-�Ɩ7��|%�y��%�c|��4�s���&����c��Ƥ�6G�YIr=�^�z�o{�I&�d$_<�Ȟ9,�Y����~�5��$��E���&�MG�be�F8\#))�����Ͼu)���Iy4����s7���Sa��08x��C#MBkRi�v箈��d#�߁�T�ɾ:`��c|5��,�y�'��߄
JP�|�!Mn0�X�W �q��8_@2[��y��o���anG4D��C��p��8��ĸ��$�d���O�&	��Y����f�'8$�=-�����a!,�S��יnVk�Wg�p<5�;��UPH���U�kUjU���-�`*ڮ�������X���ZH�۸���n[c	��l��/�fɩu���c��OqK���q�}����a�LG+��:�Zmf5��C]��#J���+t��)����V�wp�RYƼ#�mƁ�`�r)rFFǂ[r��L�v;Sp+����r;�(�����7d���2֖gl8^� �ytH'n����Ă��W9�M�������)Í�'B���:ԜuJq��gv�hm�<�=v�7��3���9IM��6mb��6�-���S�Q5����0��ފp���m��p�kEU�l{���&�U�i���=�8�+[�������Ǟ{9��Mvɢ;��=v�ՙ�A�Q5c	�!����x�c��1�	�7�ε�9���lvz]ƻ�������w�{t�:�ݦ�;vLW'lh웗��D\�����]�7@�Y0�&��g>�]��� �T$U-����n.�]`͞U���v�n_ �s��2�]���l�v��͵ֺ�2݁�ps�FM���2Ɩ�#F���q`�h[B/4�m�a-4*i�\屓ZD����d.|�9��회=�6���ʇ8�]GcL�ZXj0XV�LL����x��n��Gv{��EQ�s��N��=)bE��ȉ�N��m���밹���*�}����]���Sn;-�]�uZ���m��n�.�2�%��YD�v�5F`na���JR�.��Š��jKՋ47E��S�#	�1X9�̣��@��n�gA���l�;<�����"��I�ax�V���llDυ�\Y��Y���T��22���\��Ea93qB����3��%\�����Nݏf��6�!�m��%qk(���5��}�n�Թy��ڪ�yN�<U����4��^.m.�b�_h
]+��M�ƌ��e2K�G#�&m)cf,����7i��g��Tx�v9|ˎ�7�q��:y��.�"�f!���Q�sZE���
 ��C`�PD���#��8&� ==G�
��B!�}b
x� ��I�9&�M���0{)t�CV(�t	OZ9���e�*(�iۣ5�i�'E�v�� \2���g@�EKf��P�B�#��3N1:y-�u��Ǡ]W/(){gm��l��+�1���Ɂu��4b].���IFkMy�$�a�%�� ͷ�1u,��;s�(^��b�;[��ci�*҄��+����꒭k�鍆�m�f��]e ���������'~ws�}-��15��#�,.��7h&�Fչ�V JQ�3V[�`f㮭%[�Ucݶ��;5��M� ;$x�����"Yv��:T�v� ����G�ݏ ݎ�#�G擱	:t��un��������ﾯ�)<�`d��;5K1[i՗V+`�m�7c�6G ��x�G�vY�r��cV۫��l��vO> {���nǀn�Gv���ʺWq��m�<Sq؉�/J͗p�$�c��80gJ#b&l�RlI�t�ӵbm����d� 9��8`ۊ��m�m2�ޮ�Z����[� �ĠB����iv���d�w������ sv<�}�ԑ=uw^�7al�����I0-�x$� ڕ�`����Ӷ�=K��x�:����<U}�]�� ݨ'V�����ة��0-�x$� 7�=��������MM5)�ө\�������.&I�̢ΗggA�	�1��ؓR;7[\Q'N��.�n�I ov<H�����e����um��O���3]53h����羯�H�������<�T�Zy������K��{����s߾��@���)�1	��_S�u������j����'j���Ų^ I#�ݏ �L���pi[N�m��w�H�}Jl������� W;������F�QIIᕂ��q���ܻk<���u-��l[��Ieј��^�|��נl�+ 9� l��R�X5o�X�n�J��6I���� �x=�< ��x{PN�@�CV�LM��8�e�� s��L��#�'i!��;Eն��)�y����6I���
ֈB�`�$�BF
mb�&��q3W߼��y���,i݊�+am6�����e`;#�� �K�.�Z*�j����tq=ld�y��q�����6�xn�j�y�\�6���l���2��fV s�< ������	۩E�E�Ӥ�bv� 9�{� ��x�<��2�v�.��M�h�ӻo 6lx��xz��)�� ��� ٩�:D��`�V� �v<M�X����#�6�H�)[��U��wv��ٕ�� 9�< �v<�+�TG�vs��8�X�Ě�q�i`�CK�
�:}w�B��!�������#e6�N�-]e�6�LM1u�[x"�f�t��k[4�*)V!1-�ώ4��u��J���vq&;!�ۜe�;u"f���6'r2�2�pZ̔��r+���S:iEsmy��-#B�ƯcS)B]3�L魱0,������a�h^h�)�R8��yq�.�5����њ��QT<C�P��/��ef.�,��F��JK��B1fnj��nP&*��#gr��:s���Ҥ���\ �� rH����ݙXzGN�CC��V�x�#��W�vy�g������_RF�%�2�;�����������7�2����nǀr\J616&]�n�ݷ�I�+ 9� I��z������� �u(��]�:N�V'n����M� 9�&̬�]IBiP��_�� z��.�+:Tݮ��y��[#��R�]�ڝ6�ٕ�di2��ݶ���=[o�y&̬��^;)	�|�V�p�f��$�����P=C�Qn��~ٹ&��x&ǀwCbƮ�!S�M�wv�&̬ �dx~��#ޞx�<�w�M�eІ�L��`;��� s�&̬�5���*t��un��	6<�U}�.�����V sϾ����{�u ݒ�L���a�5�̩6`04RQ�n%�[��ړW$���;���������ǀMٕ����N|�~����>���Ä�6���zݙX��x;#��c�:�h[�ؓ�jڵn�����}A���jPV,^j�����E*$ < VY�7��$���rNy���P��7hUm�m� ���{���2�=_}�R]�y�}H:|�V�e[������2�����G�<��vŚm54��v�	[e�t�1�����mְ�n��{�v�p�6bf�v��n���fV s� od~������� ��&�"�CI�n�����U}T�M�� v�y��2��S�줩��v��v� l���ݏ ٳ+ 9ݏ ޒRʺ�	[�������kg�X��V s�Ȟ$�P�E^.����H861[�ݶ꒷X͙X��x;#�9]ٕ�N�H��wW��@�Ƌkj��a6��K�V�ly��j��L �9���cU�Z�\�s:�ϱ�� �wfV7fV��Eܡզ��V�v��	���̬n̬ �v<��$M� T��)�We�������7�e`;��RK�;�%�M�j��T���7d��wc��_��7'D�{�xnI�^�HRt�)���6� 9ݏ ��/ �wfVݓ�<#��A��D��A�$!EH@������u���lpY!N�c���=�ަ˩U۰�瞰[��.yji��te���&:�N�-�/<�l���g��탴:)��'іY�Yt6<ݘm� ���r��La#��Ч=dK`�K�g;��m�kt&���%���Ґ��m�FX�lɌ:��m�����F�l�lMA�fwN⮇\-��te�Y�n�:�nY�v:��*���g�Ns��rNNL���c��3=�N6����׫�1l�c���z���3���R�&�mTKP�M2��{|�׀v��+ ����/ �6*�lWt+��i��;]ٕ�wu� ����8�K�;6,����V'n�+u�wu� ����8�K�9]ٕ�ut�J��t'Nջ�l�������S޼�ݙX��g��~V��:i�E*���w�qn��9]ٕ�su� �������٭.��B��I)j5���YU�A�XBh�qc��B0��g����$��K^SlE۾��<遝�� 9ݶ.�o �l���v���wmRV� ��J�b"��j�Dd�����5vz�	]ٕ��_}���DЅ�][�"���`[=x�Wve`�p�;�N��C�Z-��8�e���+ ������.���$'��`ݫ�.����9]ٕ�I{ s� I���E9�Ww+���Iӻ�8!1P���x݉����'Z�s�zVF֣���ө��n���%n�	���ǀv<�ݙXV�-���tڶ�ـ�ǀv<�ݙX�p�9۔�F�n�J���� ������Ù�!�7�����4��`���1l���v��aa��揣�L�&0Ō!1����!7�z�n A6@�Y��$!�r{d�͐���p�	*H�!�Kl a`H;��� C������&Y|vr���2A��������!++d�-%$%�*��e�8�,L��5!���g�u�IdXX2e�4���[��P�$���$m�+ ��Jh���T�"��P��)�S̃��}=nAk�d'����
@�
0�+#�oi��Ӆ�Ф�y�=��ja/8ƕ,.�2�4 A�HR٠�C �����	��ܺ��O=�!R� �H�8o�!������$GEȲb@�e0!�&SG�ݞ���燎j�$a2j>�"���1H�\oN7	@��:��:��$���u�y���@�Mk��0��T�q��x���%��n`���)��!	#�iK#����^CnHNF��8�A4�h��6�ظ��Hkm)�� aCo0X@�ZA+����T�r�+�Ɏؚ@�@�JƐ$�hZop#]��Ԍ&��B0�	}Qh���)��GBD�G�t�E6�]��}8(�<1��Ƞ`���:�m1��k��C�TVkY�u���C������T�Wn��eZm�����'c� s����/I�O���W���;�vP��;0���nǀr��+ ݢЅ�GI�M��ի��cr��K��h�ax2ꡡ��
���1�D�`����NЮ����ـ�ǀv<�ݙ^������� ݉��N�C�][���c�9]ٕ�r^ŀ�Ǟ���;xK>i���wm&�����{ s� sv<���nګ���'n�&� ��ŀ��� ;'�I�����0$i��H�"6+	" �H�lV�s}��'�+�)N�
�n���wc�	���̬m�X���	*Ջ�9�݂�f�{���w8�v|��S���py'���7$JCG0��ʨXL�e��}����̬v�/UW�@wg��O�O�	[��eZ��Wveg����H���ul���{��"}=^F6�m2Ʈ�&�`�~0.� �������>��a�кh����rs�_7������9]ٕ�oc���p��
��v;w�� r�����qwe��������im�(:���N=qH��wZw�Bv���jXƒ��	�V�su љ��B�Q�HT�m�G1��i݈���ګ�.`!e��q�n,��$�;#6��+
)��	l!�	ie�3�񷃹�5�H�����W<k��F�\�.>-i#;[+�t7Y��i�.��s0r[�րb�� жQn���������_��X)��N����w�����A��������+���r쑐�s�%[Y�p7a��[2cK��^�����V���qwe�wc�;��v��T��L���lp�8�e�wc�O<���䓁|>��O��Mр��oT�� ��x�ݏ ����Y'IձR�v���fǀ����p�8�e�M�U2�Wn���-�����lp�8�e�wc�&ܤ����({l>��DQV�my�j7=1v)Hnɨ���8����/릋�,���o ���v^ wv< �nǀr}��t��[�Wl�8�e�~����HP�b�"�� F�R0���
D��@O���y� ���sc���p��[���.���wc�V�x68`[������j��j�դ��V�x68`[������=���i��T�ۦU�|���Ż/ ;� r�c�=�۠.���tQv���(����
W�a4�8Ś���el��]���::�c��N��WM��I6p�=xݑ�+v<�0v�dt'V�ةU�Wn��G�����p�8�e�;¢ej�4[(V� r�c�;�����9@O@�'�� 3��~� �'�wIR��Ci�5V�]]��n��v^ vH�����N	&ChE6�ـݏ �����kg��0��*�+��iZWws�$��C,���81�M�ϷA�U���f�G[�t.*�Ī�e��� ��}z�nǀn� ��x�Iay��]ҵt�ն��ݏ �� �v< �dx62�cv顖��2���;��ݏ ;� r����R��n�]6��'m`;��fǀ��xIX�̨?�������rO/~��Bt�7aj�� ��x�kg� �~��wc�=_W�K�� �4�Cq`9x�K6T����X�Yʎ�vG�=�7E��nN3e1���ap-�͔W�m�<�� �܋ 9ݏ��qV�^��^Wyci����V�;���x]�x��Ǟ�����6W��IS�h����`vy�vK��I��x�~0n�4�6�vݢ��o ��^ mnǀM� ���Kϭ��M�w�]��	���~�7$� ��cB�A�J�T� `e*�	�J�)���+�m�� Kf��[��E�d
WkX�HfЋ)2�HF
n��O[@j4Q�A��%�C�=�ul�̰���;v�ѵ�����#ٵ%�T�8���:�:�/���n��S�
������5ٴ�.r��X9�'c�N����p��Jb;�
'��H-��j[B��h�B4�L�	��;s`��H�f�r�Y :�x--���x�I�)���)�C�s��9�7|���&)�@.?X�MrJ������ϴ�i\�x4v5@�Z轎uQ��݂�����0�c�"엀]���[��MN�Ӳ�0�c�"엀]��	��ql�:�umR���o ��^ mwc�&� rlx;>H�e*���lb�x�ݏ �� ������v!��n�ڶ��[x�`&ǀEݗ�]����s��=>�SK	�1fӲZu�6�,�D�lf��8h�5�k���Vw/v!�8���	ҵNӶp��x]�x�ݏ�A����N�[lVݢ��o ���o;��Z"8�Հi�`M0
��$�0*%H��)X�X! �G�@�~��ߣ�?o�� 96<{%�2��WE����w�]��	���d�dwj2ݺtĮ�L�v�	���ǀEݗ�ݖ��R;VX�t�];-� ;ݏ ��/ 7�-��2���JHb����]�:j���h ˴)+�0ĭ+�屙(�Sq�	��F��
�����wt�m��yl���e�wfV���Z$9j�Zlh�17x��o ����.���!;��V�Z�o �ٕ�s����� "H6��E�H1�X�P���E"E�	��
(�o/��nI����ܓ�jZ���4�+)۶� �c�v^ջ���wc�&X�c��v�fv^�6+�'u� �c��s�y=}7�7�tD���T+�8�LOV��y�f�#50���H"cR���]v6�� �'���2�v8`we� ��tݪ�v:�� �obΤv��ݗ�uM���;��"��lN��9��qwe�>KU�W�s��`[�GB�`��}T�{=x�O+�9�p���}��Q�`@��)�C����3��`����Ui��������x;�&�`]�xꪩ�U�v��}�`]�w�vcj�
s<��1S�m/;�&5���Ye�M������"��7v��G� ����/��WE��xT�Z�,�]�t%M��`��H����"�����$l��Iڲ�4ݴ[�m�V�^�lW�s��`��y��z㝍.4[]�տI�s��}���;���95� ����;"Nm�mU���յx;�z����玁���I9}�ۛ�_�"(*��Q_��(*�AU�H�
��DPU򈠪��EE_�"�A��F
�X*E**U
�P�� "�AD*Q
�E@�� `�D��
�QX*Db�D��P������
�@X*D`�@ ��H*R
�B
�����
�H*H�X
�
�
� ���� �AH�*
�P��`�A
���A�D��*F
� �DX*F
�"���
�R
� ������@"�A �E�� �AH*B����� �@H
��� �@
�D"*E��X*V
�E��DH*X*"�E��B
�*��F *�����@������A �@b*
� `�@F� *��@�� H
�P �@*
��� *F
���D*"*`�@��@D��`*
�@��A���*(
���H��
�* *�"�� ��A �E"*�`�EB� H������E *B� "�A
�E��E*B���@H
�D��@*H
����
���_򈠪�AU��
�_���
��DPU�"���_򈠪��EW��(*��(*��1AY&SY��A7]Y�pP��3'� a�_|4@��k����b���ѨDB���EIH� 4쳮�����EP�B=d(�2�{i6` Y���h*����(4AF�4  4	 @U(QD��6��
4i�(�$P4�      6:�Ͷ�����eP��;(	=�U�^�NL���*�{���o���Y)��/����}�r����W����}�}�EK�R���ҽ��� $�c�������/}�ޤ��H7w/,}��O�����|=m�*�۾j�޷��j����lm�ە^� �Ԭ�b�$�����êj�ޫ�W.�U˾�qn��z�|��«�y$�л��5]���������S_|�
��T/'ô���񯁣D�����O�������^��6�ew���.�����ݵ[��lҭ�>T�Q,���uO6�ʧ 8}���֨V���w`�z�G;w�Q��}M��}<�P ڠ�, z{��(���i�� Z� 9��s��g@�)��)@  �ٚ Q�Δ�1ԔK S�� t�7w t�� �A@�t*]�OJ���)s:(�3�M����(P
U�}kk	  R��T�gm��.S��(�iM�q��zj�Ϫ��g�}�h7�R��-+�wW�9��e9���ޔ����_|� : נ�w��T�kͪW}��-��Www�Uͪ�eɥ�ruK���b��w�R���������&��=��J�QP���W��� M( )%*㻄���*���e\ڪ��������zS��e��>/��j���}2���y9n��n��NO�*����  
e�iq�6T��$�N{�/���i}����޷+���w�G<�>��>��o|�)�ۗ�O{:^۟a��  '��R�  ��eJ��)T @��R�F��I� ����5Q1JT @��Jf�*$  Ԥ��������Z����?�_�3��}��>�>��EU~e��("��ATU?�("��Ƞ���EUb��*��޿�'����)�I4[�	 B��$��]�hXd�-��:�Ӎ����B��fX+�������+���h^n�R���\��D	��Dq1(1�*�E�a2#9��O��{��Q��΢D��b��$D/
P�G���&l������r:�����r!/4(�S�Z}��cgT����R)�ҨY���Pɇ~�㩳:���"����>�j$�|�q�!�c}�}�ݱ5� ]J%��{�>j�O�:��ǟp��{�V�~�$3��]gh���1]�+ݷ�(<��x�����*�.����\D]\�_-�V���\����w�����O���,��nĻ��ӈHA� ����Vǋ�P��{x,�X�����>	�����v��qy
�m���!L���oj�_M˞	K������&N�+�	
��������Ro��^Z�����לuyAt��N��\�W�>�}i�t1H�59�7��Q	�(�6�Z�ۊ����y��G<�KW9��X��g����k��7��N�먏���mB8���k��DD�t�P�}U\�:��	>(����>_u}�^��Hm����'�O�VLB��D�ˉ��(���/��ϸqO��R#�xG��p��2��~�&WԇW��q�Վ*�cM���ryo^ßq��N!�M%�Ś[���Pe޲ϼ{�K�^�-�Y%Ў�F�BO�E��w�幣��!�I!��e!cX��Y_5ri����c���S$9�}���-�_{;C^_'��Q��zy1�Y��'���{�K�<��#5����uLA� ��D,�m�8'/|�:���{��0O�#�+��߹��##�*��B~j҉�S3��TI�Ϻ�����{��C�Q�X�T7�!/f ���0�1$�h3��Ԅ#9氆���#捘o�k|e�Ue�B.�)~艝�"8�� '7�W��p><�>��|rIWé�WR�I�B��!L�!��=7�xFƜ��.�ޢPŐ.�!�2��n;HC�Q��K
f�bP�9QTU|�w`��ݑ{��QBA�ĺ��$�FB_|�=����	uxfr-�.��V��C7w�_
B��s&'w���q|N숿p�\1	�w�g�:%WC��o,��������%��LƝYJqw˽D.B:H�.���f�+�ٺ�C~Wُ�[ħ�3�-1k��'<�u�F�RL�㲚˦H8^��A�������l��4}틥�CAbMaD�^l�Bl��·zՖ�2���#$&��\�� ���ԑ>MbY:Y߾"��ɉ���v,MN�3:��ݷ�έY��ϖ{���y�u����I����:�������7Ч�=�)uN�kJO]��	߷
1f`3'��E�	X0D<�gu�x|�����쐉�`�8���wR�GO�A�/�'�%|'�u���Q-^,ũ���|8�3�J'[��,Ň��	��O����j���V&Ω߼����6%��8�'��fT��xM��Y�N�T�������JJ<��ޝ�%S�46�O2D�5��Q9�B[�+-�S;~���~�/�;+��9i%5�6�)�.VZ�|Y��[!�c��ane�֋�66H�,&e=�&0��鴁rꛔrɢ�
d�
�( �a\���Y���l ���x�,q��ʸ�x&�����S����⧜��O�S�!de����#���ޞyՀ.�w�X�p]N}��R6}�S�ڻ8uA{���Ʋ��>w�|�~]\ֈm��xTB9o�]���±%��W!�T80 l b� �(�<�+S��Ϲj:��7&'�����B@�IK�.�!,���
JXH�##RHH���5��i���C|�����g���]���0��i>J�`F�ĸ$XE\|��Y�Ǌ�?=k�WY�������y�Ph�~x�������PB8.ܟe*�R�RmpR��$���3��2mx�)�2��	jc�g"E��4��\���93�x�Lߘ9\��7�}�S�7OYsi4C�U�|L{}8��Y�}���9�ݼ(��'G�ᯣM6Ђ���=����>�J阹���y~_.���S�8R�;'�DP}]���c]K�hm���6F]o)�	��ts4�s�X��=�����OQc�PB��'��媡g~���i��x��cx& >q-W���TNo9�{U]y0j�珽_5��œ~�g��RU��3�������4鰔h�B���%0cH�,#`E�q{�� F�>��A���ˌ8�5�R>��ɾV�@����5��y����x���?_���˹�B|����8���U���S�[�xk/{�]]�w<��y�������O��J����nGsT�0�IvoL%��c$q�Bo���,ߕI���76r�j��.��]\���4?7M�@6rq��^,L_.��P[�s�B7�D�	��)mi誏������i��`�QN!���q�	B�QŎjfI��^��9��ř�N^�u{�/��bo���'G�+�Gٝ���.��{�ג�w����}6��{C�}d/��T�6�z�3�O��L��I���Fd���N�s�}��躽�c�E�������M�ÒdJ&�+��8!o�:�=q������7r�L��p	!H�&�I#a,!
a��J�D�A��8E�"y���>�k>ϖ�qJ'��<��5�À��T�V��JpM8+K�@�1]@�O7K�r����X��&z��$!MHN�S�g��^T)᥌yJ����7/��MF�����A�27vB�-�!�B-�����G��č�'�s��8�b�޿�/�t��ܘ�s�`¡�Gp%����`pb��;	���.�8��q���y�\9�H���gO�m�bi�8&q�� �/��JOf����lb5�b@n|�s�{~.@���$�>�#H�+f�Ϙ\�!M�>����"o$��HK�4$��!#Q7��#���ӵ��K�x��q��G:���"CM�on�����\�oM̗�������4/���9�7�Np�}�{����~�o�%��ηx<;���bkpެ���+�Ú���\�5n�Yd�Y�nϻ�M�{�J{תd��za�g�W�uw��@�]��8�8Ϸ���³>����Ԙ�2�%�����HI���{���|�ɋ���
�\�1I�S1>�����GK>���^77�y��x��9��ѾT����]h����W{9�нL˝\LΤ	�9�.
+���FD�.G˟\Bk�b㻶��Ƙ���Չ	bώd�>�	�=�*v|b��D�cS��ϪB��r�r���tI�
yw�����9x}�~�]�1��O�E����V}�^�ǿVe�UR���?�6s�����|'`��ľ�W���{��<��ȃ,���-N��)^S�1t��q.yJ�y���Ա�#���q��@�t$��׹�:F95�Ń�=<�O���p�n:#Sa]�ɦ�\zK��$�oGמ�����"DN-B�7��ľ_p��! ��$2T���v���^�����ulP����S=5���(�$\G"y��޿;_u���ɳ�}���~}U&&�E��\��D.JW�*H�0,�\�ϑ�Ł���l���G~��菲����x?��κΑ1|�"���
�quvȒ��q	 u��&�[����><!���䧴�)�C���o
e�t�l�HF��n)���;q8�(?�s%��F�G�u#�z����Ͼ�8�Q}8��rxg"Mw������>��SH��!��&��&��QW)߁	���lz����۱Dӥ%�Z�/,��?����Ӛ躭��!{�wx���w#Ә�,|�c�us��;D������Tׄ��2w�a�O�L���||eB�V�>OF���NL;��|�P8|uA�'��Q��8��'�ȧN`�ѩ=�s�;R�>2ֲV����������,Z���{�Dq���X-O ]�<�8�	58��� �|P�4F��&&��W��x��}W�U���h��u���|�X��ԅ/l��5f���G�������^Y� �_h#m8���M'1z����	8�&EUq�,�i�o]�q&�yT$I�#�k�Ϗ�؝��o\��FҲ��c�s��N� G2;�J�)��x{R�;}�����?�`;����!�:����%���ry}��X�/~�����5�����q	ED�,|&�5B��ܼ�Y[)=���	#�~������)ytRp�h��]��;���}~~�|�\΢<=�w�RG�k���'�81L�U[W�ݑFrD�|�'�������8W:�C��}̊��q��"�Ǿ��y(� KK��A�BX�a�	ie-%�$m՚�zy���z\��|8���C��萱�M`6��1&����}��^ָ'Ə���/��ÿtk3�噜BE����!��.g-�$̒ͼ��R��gş>
v"�!}�'��n@!%#%��BV��	HI2��7U���Bo�E�f�s����wA3=�s;�ϙ���1|V��4Gv�l�x!
�����s�\A��ӓ4︖���g6/	�>X�	,��H��$���x�D�9 ����#���Z�������(�rg�uF�@���  G884Az���U�o9~�
>��~_9�Q�u����8�s����5yP�.ZX�YG\2O9xI8JK_���h�Y�'�a�lv��R0$VX,R�#�ˉ
ʑ���bK��42ʇ�C�M�˜�pL<9_����'��nN�!���7\����γH��3(�x���TNǚ����I�ͮ�E�ۇ���Bli�'-�]H���f�H��jZ�0t����
Dc���>�.��(K�a��h�{��j�\�m���Æ���|g�J���j��g���y�����#Xהݬ�Z�/���+DP$򏘆��}��q:{*�N|���cB	�ZrI�D��	(2A��O��kߐ�J��!�]�XF���ۺ��X����*���y�b;����5jN�H�T�[�޽��.k�9�9o��P���$^K�������L���}s�{��j�� Ĥe@����qD�]����}�냈;�M�_<B��R������9�G�*���D⒉��S��$�4}Qr�2�M]2�F�[e�Ԑ�ac��h�����t����DkDйb'��5n!�W����֜�p�o����/(c�x��w�J�mdB+r�������$��ߟ�TM7�}2U��>�%��Z
����4`�HN>	��)kE B����17h"n�$�-�y�����8��>"�s���2����eG�8q|%>��7qY�����*���U���ǎ�:�Mf?�Vv��N��g[?��r�Ӂ�),�-��׍���u����|k �B/8�x���ʈ�C���<��wV�xw����	����\��b�1b��h�S���\��5J�vC$�1n>�W���}:���	�L |8�����4�&�a|̮,�TԒ������\$���ߞ�n�O����2@Ȗ�-��s{�X$FW�Կ��Î��}m�ڪ�����ڪ�����UUTUUUUUUUU*������������UUUUUP�UU[UUUUUUUUT�UUUUUUUUUUUUe������������ڠ*TUUUUUV1U@UUUUV*����UUUZ��U��������*UTUUUUUUUUUUl��
���j��UX�U*�UR�UUUUQEUUUUUUU@UUUUT�������UUUUUUUUUUUUUUUUmj%�m^V(�n�B`뤖��m���<rm��Lg��Uh�a��츞�*�ʨ	��g�9#1UN���c#Mm[d(Z�t����@�:�����3mͲdr��
v�T��\�tQx�L�؃�	�ޏDp\c�G8���]`�����zZ���X�vg��#��{���c%�;l\���7IZϒ\�t&��A��\�/S�P�iImn��Fα^S&�+�gj:�It[���*�sѴ��&�Yef�kr��@]i0Ka�*�pUl5��a�L�����.�c������X��5v-DU�guork�-�%(�F#��n\��z@�s\�Ț3�x�����7nmΰ�m�\�s���mKZG��� ��^ĝ��!��-t��G�
	���ۂ�g��)J�Gj�������TXإ���Y�;W[Tu@�WZ�Fݵ*�]�j�Ű�nZ���e��6�r�����B�/T���X��/*��K5���8�1�\v�MB�յת<�[O ,��d ͆t
��a�J�i���Mq�Τ�n����fn��v�Z#	��58�X����{�"@���C;�(�Fe�of��1���$Rm�D�.�K�Y2�&��E����n;jΎ�"s������Ƃ����[e��F�um���8jk��{qٵywY����;[ *��<�v҆�J�97f`V�Z΍�ϣDtԻl��J�Pu�P�6����JK��֚nG3Z��N�kr��μ�б��eWB���B�]�M׳��-��j�4���L����*��Vg�q�h�L��v��a�͘^���l��ϵ�YC&�cBc�'U�X��c���WqdU��'Y��KTv*��q��q<��OI�غ;b�up�Y�8Ͼ.@���Kڭ�A0�l����i%j���Nsv����1���`9+��[���k��d�j�!�j�fvZ��6�i�
�B�B��-Hqr�t��*Xqn%���"b\�`��w>�wW�="&�&�v� �-�<0R�֗S[UGR�m�\�5 kgOU����Q�A�at��tU���[�$���{@�4-d���u5̎%݌�#N�.5�L�m�Mm2,u�^UVe�6�F;n8ڬq0'�H��t����G6ր���4��K�J�B�fҶ�]��ɶn��c*���r�1��j���`�Z��if�'���`���VD�%�Cn��y��j
�خRUzI��t����]������m�*�uP@��\Wn't�m� ��HT��gY%e|�uE����sk\���[�n�����#�ݹHSmmK`������[�]jR�� �Mu��#��@q�&���
S�=�՛J|x���>3��ۍCD���!<Ul	��I���ujB]5��`e)�Q��6]�2[��vݏz-vqB�cZPj��[�q�Y�;v�uVcd�#��İ��b���*�YN��N�V��"I�TxV��Ŝlx����^/e�A�ݹ���T�#�� �����V�X��i���!HJ�s��;@s�aؗ�m�Y�JJ���whb[ ����/l��@ z����Hs�:�
��_R��5���t�v�+/�;Ƈ���7��Q�KF��rtCT��	9糡lZ��:.�=��y�(��k��C��f���-�騜4�i�.�J=�7��v�{T��`oD��P�`V�6^�Ƭ�cU`JU�c����v3�t��
fh��s�ڸ�k,��f�5��v������`�:T�M9�A�06�ڀWI�;A�ћd�3صݤa��� ��Pe�e�*��#U��,�m���k���m�,I�k>'�E\JJ�XҨ��vF��i�+ ,ms1��k�ai��"�Ze9��VlG �8���J�]���&&㤸MWgq<;s��Yl�ٜ��K	J+F�xV��Z��6.��҅�Ha��k=@.��nb���X]��H���%�&�гKָ���E�
��!��:��;��b6���Y���%�չ�T�Uʏh�V�s[UR��ۖcy-�aYU��j�糶�c�w���x*�VMJ��C�9Y�R��m�v�J�� 9���t`�5k����:��m���2�@��3��lZ�\^�籺�i26��}�
���v�����b��,l�vլ�ι��1�v��N��\.��)�\b�� P.�]�AHtd]>9�K�����a���ܚ�'+"t�[S�+��'=��r��`ʺ�x5��'V;cj�30��Kv�75�����<��w���z�m��@�����6��HD�Q����*ۧ1aI���<nX� �^uJ����b���G��b	�X�bx{;�q��̮is�&� 'n8�7�����6�f�]�b��v*N{v�8¨Mu]U�1�J��q�ƃP��7RD�B[K�@��]UT^�EN�`j7��������p��3ʋ�y�7	.T��5����d���IU(��-�=�{ʨ�ڄl�� ��SF�Un)|b�v9��g�մ��qP�??W�j�겡A4P�HmK*����e�m[c �����,�r�Nvl�9���gH�y��m1���2��*�Q�l��f^NT^.{0��v�Q�����un��Ӟ��������j
]S�T 7��˳D�rql��7k���u���K�7*�]<�fU����l����⃊U�h�P*�X*��&x&�����:��=7�-u���X(�2� b�W\�!����[T�i %�`��#�m=UW\��rP����j�{	ZZ����[]犠e3\�&]�NR�x8Y����Ts��;OA�d"#N�'�A�U�F�Cp![��S&�Q6��X�mQ�i�-���P�A�:)��X8(�F�b[e��6̀��v�V�En�]��@�Q7-3i��j�H�]iK��sr��`}Z���i����@u6�h��H �ų:X�@��������VebU-�WZ���2
V%����<�2��V�.P݆�ۭ��C��Y��x��-��Sm�P��b���5�z�/^�[;1#ЗdY�����
m��8��m�U��Uӗ���K+]N˷Kx.�U�ړfŲ�Z�*�\��FUUU�5��
��� \�6-���S�����>�bk�&J�.Ԋ�@���5mUW$%vFf��SJ-�`�������؄�\��0��ļ�T����55 �T�U�EUK�����k.�&[���]SǞ��«o(�u�*�m��Q�
�J��ɗrm@[:7���n"��%�5�CUۜm U,ݐ��N��k��UMS;%�r���Wa��Ǟ:5�+��WA��R�������V`�h��%Լ����wN��&���6����ת�i{b�:���+"��C��ͽ��8D���[J,s��IP	�Qܐ�ê,�h���p��vN0[X�ŪL�Y�l�^����Uh�J	݈@�mr�d&�vX�����;CD�gLk8U�SD���ī�UV8��.���6j��X���6��쳵Q����PS��mn԰�1,pX�UU6�X�8�:�ks���,�e��(��SJ�qJ��P������v�S�*�n�ͣ�v�)���`�y�����k�sZ�ԧd���I��fv:w�R�A��΍�5���,K!����V<]��x���n��UA�R��X6]b�U�4��6��׷!<�vCm�j��R�'\V�hݵu��B�AU�l�U�6iA]��l��']��[h���k+-��!�[�k��U]UUM�I@K�6J�R��%E��F;�X��Z  �ڈ�V; l6�2�u.�tN�XخX��GJ�^��왋��]�G.�3L�� �UU��c�.z��8��I34�uT� ڪ��iaHF���;T9c
;TYZ� ���	���U��WR��R�W��62�^*�
�
�5UUTq�I[��^��꯮�U�)����	�@KV"�@,����2�G%(;Z��Ӑd;v�lm[@I�u�]u��d��T>~���aq���ktPX�d� U����Y�!�[V��PSž���.�8 ���a.��UVX�ff�����*�`ݮ�V�8���ma�Q�.۷-=S؍kvA����B((k+f�69�ܽJ��c��r��+<�����aȼ�V}�&�Z��Sk�aF�r������z�4Q���=p�'	q��f�T*�?k�=����[@\�&��H�����
��[)0���܌T�e�U0�6�qZ�ST�r;A���Zk[�1z���oI��.Z��+�#Jg�X^@|[:Bڪ���e�
@6��R��9�(�#�m�T*�4`ʎj�6��\ɵ�֊���H�V0n�����N� �׀�l���UMH�]�d�l���%����WGu�76�q�;y�MT�i.mո�J�
�ڥM�y���V������b��]-@OmM�l@�d��[iѵU4���UV�]*�Uv�*�[*�
���HAye�h�[�*�N$
�Z����I�q�` �������uE#v�UUm�UUU:�دP���������`=�8��},�̲��I9P�d:%�h5o=�mMt�ںt3��Vd�Mv�ۄ1[+�Vj _i,n�jY5�UATU*.�O�D�����W)� ����b!� $���@�H���J�:0 b$HD|��b��
~ !�}�����U�H�" �Ŏ�������E�M
�(> �D��!�I�B�!���"p��Ê������"�cU�T�Ac"��`ȉ�� �ڡ��X ���"Ă4H�_ S[ �QZ��T��B*@I�ڨqA�|ϸp�
#�!Uv��8� Ĉ�#"0��dc���=G�(�"�����W�LD�	��d��dE�,� $g�iP�6���p6��$�����|���V8 	cO�}������|�*��=D��*A�"�"*C�8��/ʣP� �<Tj?
?@�)Ux*��5d�E�b����U�pM��:�� !�D �8, !�ũA�d]�Q��8+@!��(��-�)�C��R�� ��	 �> <@��#(E�b DH�V6¤,$PH �<t��w�R! �	0O���C�D�@�Uh�� B!(x��� 4��b�@#�����o��'�}@>O�'ej�D��OX
B
B z������W�呏$%FV�*F%#hH�V�0,-�B�) ZZŶP��$�!aVKF�D�l�I+Z��B�D��H�[bK)2�x/�#�@�!!	!#@�BD��R�X!��d#Ǉ(�A �Y$<G`�"/���)#!$bH���"H�(i' � R��A0pZ.�����tPEW��~�J(N.�1�@1(`�b��$�Z�Pb�B��0"P,q1*��"$@"LC)��*ңE+�bL fX�6���i
�� aj��S is�BJrsO_z[UT@Yj���UU�U\UU�Զ�Q��6
�H\�qUJ�m@U�UU�`^�v�͔�	W�����`�2�ڏf[����n�m���r���me���H����V��`lA���k��l"D�us�sh�݄�m%^ԗv��7�	2UH$�u�.�50V6�y��@�����Э,����-�u����^ۮJ�8�`v�K��e�[)eji��+%��Ѵ��c�E�ؖ.���-׀��u�[��@˃T	8�n�؋����+H�36ڙe����͸K�GmR.X�c-Yf! �[�3���wg�3Yd��N�S��61��1�[��+3���z�P^��x�n�
���N�J���/l����OO �.��g�Cp㞭&��Y�;�n��q�L���)����5�v8磋����X�lq�=U�z����c[K1c��xGBcCE�$B�ж�Tj�u�G�A�WkˈZ�a��ƶ$&��4��rl�j�.�&�vmΗF�"�E�Q,&=m��U��)/%�pnQF3W(h��sn[�-uv�N&���M-��Y�C�E;�ø��i���;��]��ri	��@�8��<6���cxvmn��YF��+!"Vh�ѽ��u5�#,w:ch����\g��l�8�܈vT��.ǖx]�V�5�#��8M6
�e�I�-�	�06��C/S�C/I���%Hp)�͢A#5@���$ff�s.7�y��s����n�<��X˭ѳ�m����LE͞���1U��e��pB�lہ�3\A��1���M�(�R��-v�4t�Z��ְ6N�s�]�lk��ne�,i���J��qW9}��D����n�6*�D��.ە.t.�����,$\�.�l �k]��eS-��]�Ӱ����N�ǚ;Vlj��6;kFҸR�̪��0kT����t�ԙ@7VR�
.�N:r[7Ra����&�K��(��+n�<]�;\�줙���SI�VY3B���O���
~EtVm��(h����(�M����� �g�T�PM�N�Ӻ���Ri���[��W�[B��Ʀ뭻k�b.Vs�`�n[�	�Ԝ�J-j���Pt����Y��ێ.Xm��3��
vO�@i��e�]�"BU�8]l�9�l���p9�D]@�8l��<N88�;F���܍۬���xڻX�����hɷg�+u��,�$io�z2�[�7a��XY��p�\�#[3X@�X����3����t�{�s��Sx<���q��=�A�{m�� ���T���G��=��'ڟة��ـ}�y�;����\��ǵ`{G�	M�	�JJ���l�Lsy�H^�q`�u`x�������N�4턳 �}���{n }�ۀ}�{f�Oj�1T��	mV��V׎�������,���,�6:���n���{ŀw�y��!��� ���9 �������m&6�)+)��Z��s0�J����AkcE%�nI*��-���L1�,��V��X�j$SrD�H܄���ۦys�m.>p\�q@� X$r
�����7����'��p?zm�>�nZ��ڕB�\��w�Հy�Vo9��nv����5�g�{�T�5U�� ����٫�X�ia�Ľ�j�z�W7�\,��g}� ���o��wv�����n&�_���n%
Q�>M҄�s�A�99z68w�]�p���Q�@n�����v����8�-����o��wv�g}� ֎�o�Q���׎�&���c�1�/b9	�j�-�0������1n�������}���h%��,
$�,�cbC f[�L �}� ��=���%W��mUM���X��`�u`y6��}7Z��dl�����L ��ۀwf��<��� ���@V$P�a���[�mut�Pf4�ّ��.�fAbۙt��F�;ZqT�jU%r���� �Ձ��X��`<�iȐ�B��&**j�����s��$5�v��������A*8H녍�f��.��L�yďcڰ1n���%=P{F7mq�-�=�`���	���rp;�*��6o/��䝤�� �GTE����� ��ـy�c�1�,��4	l����(U$�c���l�chݟ��Я��/]�k�S]�-`�leBiY[LuV�
�q�z����y��n��r#����X6%��)�&���JJ�l/,u`f:e�w1Ձ�ۘ�7����2�#�B9n�m��;��͈�K6wU��'�`u�VPh���j���ߤ�?{��V�>�|`}~ۀ{�t�7v��#n�
�UEMUXrڰ68��t�����$Є�� �Y
@��o=�ku�5�8�ܮw4cB$+��ZC&N�s��V�-��ث�����:zh1���������7�Ʃ��% {7�vE���:�F�X^�F#	ȇ"�r۶a�,)��S]ai6x[2�+a�$U^y[U��.�@#�y���2��e�e��[F��:��K2��(�H�t�n�ls�
�n��S�ݴ���e��齵k��װV.��w{�����O���},L\p� .]���˝��G��9Ph�lF/-��+��Ô���nv��L��Xrڰ3�JN%�����8����3���@���=����<��>M���C�(�T���V�w��]X��`y�$�	ťIO(T�f��c�7w�`b�;Vc�XsX'Q31*���YmX_}6��]0�{n�>�f�S�����&�e���@�9tb;�Y�`p"c�y�JVS1kr�.�maicn)h�8��$���M���{n ���y��9��=���p�T���hـw�s�jo��+����M,�:4FL<T=�#0��.,�'�`5�s`6��)��*�U[m�7��X__�����}� �}��IU�KHX�`~��r!d�{V�{6����w�#~Q��El!d� ��l�??k���{���gj��fB�
*d����kb,h���sr���������<
4jM�!���r(�GTL�� ��� ~�q`m�`5�s`u�$�quS�)IUU�����#�wI�5cٰ��z���9��+-� ��t��>�{�n(!�1�<A�2g�ް��ŀw��7��Gd���c� �c��Ł��S`wK��X������� ��q`=�s ��l�>�&�X�����UF5	���l��B��i`"�NaQӻ\p�V੸H�ªUS��{�ŀn���f }�m�;��r��)ke���X[j���l����w�������lU�\_}� >��X��,��ՀC�	LĪH)D��}��ۋ >���Iw�
�!`$�"����b� �T_vPϵ���IϽ+lOS�k"N2�p���>���]r^� ��ՀG}�B�(�*�D}�,�	���L�ِ�ņ	`��He�)�e����9�����)*Ugv��ϧ�V��Ƭ��V�;�<FN�ÊxL1U`?N5s��$�Ձ����>�����o��Z*��;f w�u`c�q`lu`c�j�x�W�U3%T�)m��ۋ >�p=�� ��� �wTKcKc,Nڰ��V'�l3X��XDE�琌�
Z@�FX$bB�Y%��,��'��l������yam֥֬ʐ�R��D��wl� ���吤rT�e~��ާ�������VFS���b<����G��R]e��T3e�Cj�c����x�Gx�,/0����K�/ �1��枻A����{<�D�6.wd�JGd��'Y���6���nFz���K�@3��(�IF�k���3�:\7c�Û0m�DAϻ���N�՚7ε��]��-�h٭c�b�;\sc[Yb��f�#U��;ڞ�\a�6�D�����jy�`�����q`uf��jvAؚ�&[f {��`y㸰�eX���#	8�R��(۲���ŀo���wf {�ۀ{�=6�D�/�#�`ی��� ��V�X��X����WÎr��ip>���$��������:�`8��r&�%ML$RvmP�*�1D�m=��ݹ|h$�ѕ8Y��99��QР�U-�0�����ŀx�؈��vl�ԯ��f���Ff���<�߶m��D}b��"A��r�͆I�����_}�`�������V���X��`q�V/76�c��ŀ�.F9��k���{�����n��������Z6��dB�q�lXsX�4�,��Vy��x�n�� D�q?;y ��!9k�mM�!E�I��oL+���Ιz��m�t��)���n,��Vy�� �c���T�D:��#�`ۦ���Hy�q`�Ն�׽��BF`�B�)�q��)n o�~��{nW�M4F�W�C�����$��$b�p�[�!�s��;Mqt\����-���|-!��H6; �$7	�D%Ѫ0�0!	f�&���1VG�������n�Ȍ"���A���s�Ç�"N;4Չ �{2c1OP�&FG*��o7�}����ݢk��zV�S�B��\�	�@;B�.s��u͜���Q���RC{�2��b!q�����ma�hHe��r�Ҥ/,�P��z����>TɓǑ! �0�&sG���g	��j�6���MDs��w��� G���h�(.�<q:��]�g�n��.����9o5���~axo�5�w���)u���ndne�)���
����PI>%>W��v-Es�Wq��h�e���p��.����J7ѬV��xỷLf�����t(�ﳄC�!�N�>}�ӂ811gˢ�`h%)"��&�d��#�\�%%�� !y�Z�Gi�m�����e&n��y�!C����Ӟ
�@��1�Pچ�<G"2B
�"B)-�H�h��	SB���
%v�|��T��<�l����}�1L�U+U,e����<w�c��r#���nՁ�tWɚR�ED�UXx�,��V�n�3XȎq>8�`�@�)���,�X�-u�Z�%{r�u3��.����x5�f[.
�+;��=���<�Xf:�DGPf���K�
tP��	T�6�n�3X�x���ٟ��x���������*"�UXoj��c��:��l��p�j5d�IdTu�m�;�n, �l� �7V��G!G�\9�H0�ڵ!jJ@=v �y�����߹�µ%W�CvՀ~�]��~'�z=Ȉ���= �{V�*(��^�I
ob4H�^�j�ڷ6.ݳV�n�z��mq�:�
ͫb59��QbspܪUn��~��j�;����c��:��l�����*V�X+%���� �}����I�wv����߿%j&�*����Fc��@���6�7V��V�q�+U��Yj�>{�� }�ۀ{�p�ۋ ބ=Ѧ�cM�hV�7V�G"�v�f���9���˹$ȉ�=	0!���t-���>����ɚ����vPUͯls�XCF���9� ���Tg<Ţ=vM���E��v���8E�rb�Pcn�Cs,LQ4"KH�,�[f�E��8�r0��DI��,�����W ��۲�z�ΞE�`B���Q��nש�{5"��cs[��6���q���0ҶX�Ա�+�CJ�ͱb�@e(B�d�:�m�)��7]�հ����;�'�zwt������Xj�5����h�JV�Z�Khб5&���tu�⋀֧8��B
����V��Ł�Kb�wv��P��-	+j���p�w��Kb�y�����1�˚�
&Uy;-X{7G������p��� �O!�ꯓ�p�n����� �n����+iD�0EDMD�SUU`�:�>�w��=��
�>��˾�lO��k��"�dne&���\��61�Bk��T!("��Kq�	N�V�n�"�In�}���i� ;�u��u ��X7b`Sa�QU"*U;V�Cvg���s�%�,�ݽ����{�ş��8�=���7��J��I56�{V �%��q`<���:�����$��P�UUa���ڰ=��KNl7�{^Ձ�6F���P�L�U��c��6#]j����XmՁ�G"#p��[�@�򠓒��,��;mvրק��Bq�3�*5c�P���5�̗�RJ�"j�j�ߧ����}� 1�[�GP{�Xf��[�<S©J�S`�:��s��ڰ1���3&���q6~�ߛX:J�F�V�p{��rO=�훘�&� }IXDA��p(��s��"�T�%�� {~����I�����%MU��5�bϒݓ��nՇ��r�ݫ��L
l9*��J�UU�Ss`}�"9ȝ}^ }�Xx�,����>B2�4׍e1I��d�B��i,�p�	 n�(�M���9",��w>��oq���PR��5> ���cu`{1�o9����L���ƿ"�BJ�ev� x�_��s�r#�#�����o��`���s�&�����喑���In���X7l�s�Kۻq`��`6��&(���0�UU��ݍ��֖ ���nN#B-�H� �b�	���!�!���|�ܓ�gH[�y9<S©QS`w2�`o9�wk�y���n�s���=�RD�)&E6pkv�2�v��43'.�I��+t �@��c�_�wL��L��Cd@o�m�~���ӹ���i�s��9�n��1��3;$�Z�a�fk[�s�~ٿ§�T̟����`f�|X6��"69�rd��L
�J����U[��`w2�g��Ds�r9ȉ�~ߪ�׿\Xr�rT�$��*����G#���K {�V����W��Mk]�?k[���v����f��aV���{�� NI���$��߿�3I-��j�Iu峽I)�z9��	#�|Y3f	�bn��H�v��J�TXh��Z�6��(Ѵ�����GYmr9�n������;���pp�%�\�JV���ǉ�Լ;�aW��!�u��Q�8��sk-�zF����uǫ��V��|�͆x�Ph`��[p�bSJV٦��!������`3Y��	Pݢ��a�\D���Ts-g�䃈�v�Z Ĕ���I��=�5��99?I�a�����JR���B�����/o~���P�w`ܷ���`c�leBi��wOL]��CdcD6]�����s����ZI.�[7��9�JH�z��B��oj5�U�4%��O��s����9'�n��z�Gӿ*��]�}���"#�3)�A%�trx���*���I/7zw�$9ƪ��DG"f|��;ԒK\mU���m.uE�,t�.3{��I?��H����^���RHO!�ZKyȎDϵ�N�	=��Z�P̷6ܹ� ����;���ș�UԒ^�zw�$'�j�I7X���A�6y�����1��`�G=�vx4�d̲r&j.ol�ϝ;�؞%�e횔�UG��Ik����]yl�RHO��G9��{�w;����]1>�mL:��m��{��9Ҕ�9��|�ґ!Hb�xP"��)��D�i(�0��LK�Xs���q��f�u80�u n�����J�3)"a��*k|�j��D$L�R� �QEy�����m�ǻ��P���j�9�r"fR�5�A�D�J0��{� >��� ����;���ܒr*�[��դ�϶�;Ԓ�0B\ԕ4��ez���M��߿N� ��_��$���ޤ�9�Lν���[���D�J�4i�Z9�m�ϧ٭�m��~E=��|f$��~���Ig��;Ԓ���*!)P��u�5,���d�C�-�6�+G�v[��Ɍʴ����Kv��x�s�F���K�F}�������U�%����#����%O>�g��~�9�.�+�q��`$�M����URZ����$�UZI%�|�￹$�c߾xm֮�3-јQ�I'�{�I%�:�HPAk���8B��aaH�P�F$Z�F�%���$�_~��\�~��@�����n�����o"""&g4ګI$��k�I!6�%��Nso|��Ӿ�/�Z�Ho����V��I.���RKy�"�ٮ���{��So�{I1�ޯy41����"l��EV�heDW���搲��5��l]TҦɊO�ww9:�@/P�\a
���O}�=K=��ޤ��r��s��ve$��k�I-�$>/K�cYv6�z <�����N�e�3㹛��|���9m�\�߳[�(�ly�>�Tfc�
��(xog�n�m����r�@C��:֥���[��߻�����h�ԛ�� h��NNs�3�ݮ�$��f�$����ޯ�w��9�)P������FE480�2�A�$R$B0�N���R"��| ?(�3��37m����d�4���^� �o=����s��7�df$��߉�I$���z�^�	C�A�·�(��<�joZ�c���5�p�
�4Vi�"��:wo�/�K��Hĩ�]I$��c�I/L�&m$���[Ȉ䟿`/�߇��~�^��Xj�WAY�`��{�]�s�rI�*��=�|�UZI,�>�{���̧ ���)JP�n������?y�z��Iͥ���z�Y2�fm$���Ij%!T(UW������I����z >�����`_3=>�ݷ����Z�߿~�9m��ڥ�tE�kY\m�� y��;��NIȈw{L�$�}�w�$/c���UÓ��a�6�?<���\|��8a&�������H@!�R�<�B�-�D,)�6�"K�i�h,�+�}u�ak)�Gd��|y̭�K
6����
�����m��2p�-�8D""�{���S��KI F�	I--�"���l�^&�p�d#�b.]�3A������&Ȑ�o�����g5�j@�	e
�p�A�v������ւ%C4D�j).��+�#�B�bSI)@�H�u�`��-'�����[����m9�л P4��B��f��4H�f�r�lW��//4y���UPZ���UV*��*��kK�g*P ��6�V��Uʴڨ�UU�k�h������6�{n�,tnݞ�3�; ]yݑQ=��?B�!7�j=�0����ЗJF�(�m�T<����h���Rݡ[4b0��"b�!�WC%���-�:�=ZPn�)n�2�Q���S���We��K�e��ڬ����N�F�q��(W2��O�x�ݺe;m��C��X��Yr0�t�%�z�ֶ&rvxlK���dx����0m+4���Ԡ�ڲ����@US�;�����u��e��nv���YA�$���޷<j���5�j�{�QL19,�`�j�.�S&ގ�[A�ch�7@s�YfpY���dی �gke�'$�d蔞w�kt�1-��I`��Vi-�hܪ%�����)�`�,��k=�Nݜ#ۀN�3=Z�8�`�xe狞����q�ɢN��=��أIm�-��aP�X��Ϛ!�m�k���6�o�vJ��lț�%�n,]i��%ҙ��- �8����H����{Q�n�F�;-�p��tA�s��K�%4�/e�a�ܽ��sz�t��6���z���W�����{m�6wLZ�V�g8�T��4n�l�^j��Ռ�0:&Z��i����٣��r\����m�u
F=���*���=#��R�Y)���7kR�E��v�O��WC͠t+�p	�s/7�؍u��i���6���^h�Ce�d��:�J�
����=*3plY����9�Z�<�����	��!�9�v�םc-��4psicX̏81h( Z���,�'kj�G�S��OD�B�� �;�6�-a��۠;�M2���g��%Q�¤���*.�p�¼��1��]A���Y�X�į����V�J�ۥl�\9� Y97iɱ��k��dr�3�X�X�G��[[Ax�m5q�.|����q}�cf�I]eu�bzY�r6�ղҲ<AWznY;FQ�X�t=Y�R:��h�j������B/vl|U~�"��E�: >
�#��/�����q�8黺ww������X���,)U�ͷPl������8�����qe��]Ev��wd�n����X	��;nl�8'B�6��3�kv���&�vm�͍X
i���&���`��,�g�ݮ�G2���h 
�E�K5T\BX�qx�<sŶ ���v��:Ś�OD�\�k��ǋp�&�˙cW#+�-��;11;��8[����ɛȆl5[��4�y�;8���P��Qa��ղ\��,l/�֣�����.��i�c(kL�,f�[��ŀ�ZO��Hu����Tfc�Zeg� m��۠���I!{��#��̤�w{�Id�P>��7�@�۠�����$���NURߦ�$����Izg!���9əG�{�s�]Q�W;��=~N�/���r�  .���:~�ݶ���߳��<���ש���n��)�I9ɷ�����$�e���HNq��R[ȎG%c�*�g�}�r�SU�3\�� �o'���[�r#��{��$���U��x�c�I������Q��;-#[H�6�@�kZi� K�uѣ�U��z��Ӽ�i�n/�nJ��� �߾{���z= �����"{\������~���f��.�Y�kZ�-�y��u�4(H"��$j����"�X�	�H#�##JBA!����0@����j�{���$����I$���{�}�UR�>�?���s���l�@�w;��b�Ky�"&ecݮ�$�/UZI&۳�����W+:���sy�~��$�ǻ]�Ib�jm%���#�8�}�IxY������n����}{�yȇT�g�$���;Ԓ��2f�IVI�S�}�.3���mε���#�]h��rYz�m-�K�0��{䓺tϝ�������/� y��m���}�w����~P��kV��~�9m�w�ә6f �@Ս�&6��~_}�s�s�H�&�&m$%�v�Ԓ�8���G"9�UR_F��G-�5[�5����)� ~��^r��#� G�:�����ݶ߽�xs���L��$��e�fh�v�Ȩ?�Z����\���\ݶ�=�����''~�P�{�R}��u�UZ�RK�pT�I�s��c~�y$��l
�M��v��m�n���D�j [����uf�ps:�:6�p1�s�4m��H�ϒt�о�GD�r�J�l�`���s��?{�`V�I{���9�zRC���$��������\�����N���9&�K�w�$9z��I{�w��D̬D} �t٭����n��~���cUio9��D����w�%�\j�I%�]���*�l�ߛo�:}�N���ϩ�m�w����s�뛶�h�I�$XE �C����	�u_S�s��u��~=����\�����q�ݶ�=����G�}���s�m���_�m���s٫CM*���GE-0��Bq�:Q�Χ�nݼᱦ�tF�#��7���Ƴ*�,H�%r�U�~��`���:��G":��Ł���5M!%SQS`����9�r"&L[�M���,��s{�G3�5Adҕ�P����<�ٰ=��Y��%��l����j�{E-�V�$�Kp?qr=�Ł��l�������{V����Al����-� ���f������}�x7~�1��9\9A�,���L�5Ķ�Nja&x��v�QU�5]��x�"�9�ga�w[��[Hnu�j1�v�%l�.mf@�c+�)������e����]�4�!p5��1lp�j�d�^��r�jP�F4�lY��<���O�}n|Kb��K-�X,6�շV�D��2F�U+��RX���3kI]\/V%x���A����-j��ֶ��A�T����@r\��w�;��]�?��ӇY,-�9ţ�9m���6��5m#5ѥc��0�/9����M�=5�3�T!LT���� �c�1��Ȃ9s������߷�71\PUD����� ��W�BC{� ��Հy�W�9ď{_�(�J�U��0�߱`�����D$f�Ձ�f�1�rMU	
J�*��j,7���V��VS�6��&�{ ���&'h��%Jj*�ͺ�>��D�DFW����}q`��zz�ӒJ��N����,n��t��}����K<�Y�`��X �YZ�'��c4��kpM2�o�����n��w�o�.|���߮�H'��%R�DI������7Qb�P�z�rO���Xn�X^:����G܉����e@R��S�5U�c�cuf�#������b�>�ߖ�Q�"�c��n�XZ�l��,6#���8ۀ~����ȯj��K%��}� �7q`�V��X!���P�)��SD�Z1��ʅ���/m<���ф��+bF�
�'$��<�Sh0�pgwm�߶��3��ͺ�Ds��Z�l�o��m��7U�� ��m��丒���X�ߦ��7q{�s�H�1�Q0�QJ�㴷 =�\�كIT �JBcb��	���	$EY�
����?g�ذ����;�h4]UBT�-���qzu��{������s�s�o���~_�����D����ݸ��"'[^ �ݫ����7Om p%/q�1fnu��k�'6k�d��A%�X6�6�&���Vj�\K�MUG@1��`mՁ������Pc�ŀw��oW��`⣢n;p�ݹ�#�Z�l{�������r>�rd���.]A��IQJj�_o�`c�qf󐑍�� z��{�3q3	L�"��)���D'�{��� ǎ�/��������srI�{�u�Ki�j!UUME�{1:�x���x��ǎ���ė|�ڟ�x1�(*T8�n��I��J���j��P��ɂUs���a�g��=}|m�LԉUM*� o��XO���o9�6�����TMB�L�U�����"���mmX^:��$����z�~�M	B���������=��Y��G��XZ�l�a��U5T�UMTXlq,mmX��`u?l�7�����7�ѡ�WEv��:�69�׳�n�X���|現if�=��2��;c]C��'	���٬ѳ�����V��E���c���m(3-�\Vְ�tNI�`��FDBN�]�=pgU+Wq��s�vەW@Y�qml��]��Onn����L-[�-�hf��eH�˻7X��//\�9���aNwl]���zq�cz�g����<+2��͘�!��&�t��l��!�h�=u�6�x%6����\��t�;�t�ߟ��6ؔ��)��ij 5���[d��aw0�
�+	�upK�!��F�2J�SU�>_?���7q`�N�#�����h�rL���S- ����7�H1��`�j��x��9�r�ݙ-�m[F;m�`�_�wv���	ykٰ3�X\0Y�艒�JT���؎q/f�XZ�l{Ň܈�G#��#��WދY�IH��
A0��R����b""3�:6���;�� �^�-M���֔i��B%U:�sH�Ѧ����S��@ƌ�ɮ01��upB3^��X&�K:���XW}������_0���� ���	�^[%�C-������p�D>R����Y`�"P�� .���E̅`7�I�sq�!$�k@�X0��e `�S@�A�d��z���6�;��G9	�ħ&��+���`���|��s�s��%&��\X��Ł׍.]UJ�*���3U`u{�x�,{��؈I��X���$�Z�GS- �wۋ ���3{ x����6n�	�J$�8t�3�.Z�h�JQs�f�"����&h��Eٳ� ��;P"���gv��{~�Xf:�:���DzC>���4[�֍HX6�%X�{n���`n�,���Y��_˒���i��B���p?߿�����>�%xqh{�Q�q���9a��{��(�$�j��'%]HDC�j�Y�3�! � P�IjELb�z�&�5hAvE�����jRR��tݱXa�B��������D���{|���@-�����$d(,	]VW1����Î ��8!�fQ� �[��+�B�YHH՘��埦Ns�������	!�֔����A4[F�Ee<f�$�$-֍����3T�2i�R�+�����gD&�!8bU_T�H�$�Ő}�t�P�jB�{]�& R�]����ev��MS�=�r{�u�k�����M���a�ލ��ˁ$!�>"!+-���;Z��2"/���e�1��8�8$!���CP�f�%�1��9�/}PL@C���О
b)�T>P��G�@=W��^�ȿzp@��AS�W��f �(�5����rI�~�$��9�5Q*�L
I���ՙ�ذ3ۋ �n���`�hq㼖K
�;mE��bw�{��<�ٳ��X�n,/g�ϩ}�<��T���pơ�J���̔�,Wm��V�����6wטoC�c�9TLʪ��	��W@�of��7q��Pf5���.UU���)MU�՘���7q`{؝ŀ{��#3M�ʵH�u2��`�߱`����$��G�}V-ߦ�kc�S"J*�B����^�ob�1���1̈́�s��9� 0`��b������䜬�zF�ѫ܄� ;�m�?s�w���ۋ���XG#��
(�� �������r��N��$&��k-��H�&�b�!3J�*Z�&*N�r[�<�~���ۥ��`�6:�����@K��TL҉�I356q�,�q`�������#[��\���**����f�X�uf�^Ovl���=��%���R�fUTX}ȏ�e���`b��l�L�>�� n�[�V�ڂ��n�NK��s�ooN�����<۫���/nv	"p��%�5U�l��Yzڎ
#�ƃ��*��n���<�M�ӱ�Hrf|i*0��b�6�p�&A;ַv {=n/�(:�d,u�a����68�&���%�yЖh0&!5&%���<�<)�����v�E��O:�W&�Ly����k<��L`��v�]��z�oF��V�k�TcMr�is(�J�� �Ֆa��ܵ��m�[�k���Ao�޾��[��l���&Fԯu[�8ܽ���+X��C������/�7�!s-["���}_sŀ{��1́��y�j�1�l������n�Xr�X�L��8��xi�
��%A)L�X=ڰ;��Y�Ȉ�9�L�������`ZmmN
�H9-�N5`w2�~n��c�ı���J��)4J�LҰ;��`o9����tڰN5`�LM ���	?�g����<�Z��-Ѳ�\�j1v�,L�y���YA2���aP�l��~��ذ����_s��������6%97�(Jy��Y�ѹ$��~�����]�TZ��9�c�!�N{?~��w$����ܓ�7q`�����nT���{^�t��Dsv��1�����7E���%)�a��佽(�ۋ ��(o�_k�5�k_�\հc��K��� �n���X��`�;��� �TB`[����se�6��YM�(wn��ո*��	z����zZ�Kr�!�f���f�Հ�q�1�7��Pnn��<���~P�t���}7^�t��w�n�b#����+cj
E�1�9k�=��� �n���I�����*�=N���w�nI���� �{A<t�U
���`��X��X%�a���=�,�ħ&�E	O)IS5Q`����G9��W@ǵ��7۸�q-H��lm�D:��+K-W'/m�]�=�5VU�=p���������Gmr7*Ur�}7^�m� �~�g��y�O����$�����6k.7*������t�؎r5��X=����s��6ښ�
Q5"J�����c��6�Ϲ�^s������ �Lv�"�27%X�I7�߿\���ܓ�~��rO`)>����W�~X����i'E-�ޖՁ��ooN���ŀy�Vq�)7RBh[,�^"��a�]�)2a����\�ץ��P��|/���[r�]���t��X�w���#���Py��� ����PK%P��m� ｸ��� ̓��~���?~��O~��o��?�d|�%-�������Jj��7~���x�ݸ{�ŀ�I��nTQS5V�svl7v�y�����G�O߿������(��X�`|�XG#3w���ڰ<����Ds�@h�:�0b��h�J��y$�ܒ����L�5Ip&�Z�e�;�� �.�K� ۘI!I�p\�;��nf��d��c��̓-��/U�V�1��m8U1 ���4�j<�����S]��C�f�퓵�X�n�8�$Ů�7���Z[�(� v1��a\�c.�Dm��a�9m� k.�@���.��P���ƭL�k�t�0�a�Y�l�VQ����/�;[Eի�`���N3���rs�k{��$
k���T���O%1���\�9ݒ'
��e��v���~����Q�`ۮ�o@����, �}� ����w�pv ׭ت��##�U`x��8��7f�=��n��H�d�	Kf�L*"E3U`b�ٰ�u`w����ݸ�k�TU9\�u��M�fc��n��:۫��'7f���_����T*mW-�;��X������ =�m�;��E5�v�O�+�Tv,qj�I��\v����#�����_?��*�Yƨ��prZ� ���p�[V��_s��>��}q`w虘*��Aj�[�w�u���s�\Ĝs��s��Gh��`{��Xq��H���sB�bI���%U+ ���y��>�r=�j�̝�`y�&��PLR6�[�w����������$��\���j��;-� >�mXr9��� ��X��X�CP�nݭ;�ۂ�+��I��ڭI��#q�3��鈮Eq��h�B>ަ�ĮЃap�@̝�`���=���<�Հ��d8�	�&D�)�V�n�x�fnՀf�Ձ�Kj��H�|�+U55DTR�UU`��`m՟EG9�9�8pX+#!$H$IHU`�V"$�Eb� @��	�C����s��.䓿{�nI��)d8QI
yJHS5Vr!,�ڰ3]i`�Շ�={V ��A�P��J`*��UX�`}��ov� ��X�w ����O��+$m�H6��X+�0�%�#����-�y1�Dl+Y�?�{�-��f$�$�
����Հ?c� �n�ﮘ�笘�8G`ۮ�n o|���G܎D�=��>{_��VPǳ]*v����n }�� ����9ȏ��ɻ�U��߮,ǥ̈�ID��)���G�zXoj�~n�����@����Ea䈖
|m�LG��s�ܓ�ɖ�[
�) �r[0�����/�.%��������k1̀��B� D���W
��n��)�6m����05���ڑ4�����UZ�[�w������=�mlG#�@6���I�HS�R)����u{Ȉ����V��\��ş��l;��h�k$�u�YU`f��`x�Ϲ	<ݸ���`n���a%P�+��w�pw]ŀg���9śOU��T�(Q3*�IT�UM�ה� �n��S,Y�ٹ$F�r�_'�����<��8@�)���HŐ���j�<���M#�}�D%���H�@��Ja	%�x�5��P�R!H��d�6[6b�8�Q8�0@ qJ֜!13Ep�����bD.����.��8l��D�(������$�!�x�ӡ��`�2`H1b$�#��w��3!0�o�>ִT@W[UJQ�U@UWGUv�Ò*
YP�4�A[:⪕jڥZ���������j�3�m�3�CN7�*U���m֍��Hq�ۣ�q�}�%��^M,��*���Pl!�����ZA��U��tel���2�tζ6�2�틮C[kb;;r�"�X�ә��"��ԕ�ҩ-5��$��QxNZ�N��s��m��Њ�v��ն�,�`b�D9ak��K.��W�[�"֑1Ő����u���4ԍm�[��Z��2�Z� �ML٢Q`�`�)Yלs�E�ڶ^g�.*�+հ�����8���eŅ��y�$�9�l��u�ll�'����헶�6d8� �k����݃W����*ո����MV�|�����9ȏ�Z���n�����ˍ�58�]�r����B�b� gQi�
�:1�mu^�-L	�
�Ѽm4�p�Ц�_#�s�b�]�t9��CM��2v��x%e�Y컆x6�Y�������*j�VY[�]6�H�Ô}n {\%�غ�T�)6v���z�� 2�c{t�AĻO��{k��c<,��K���3�#�v%��u�ttaR��й��-�����\=r ai���#kJє2ʍ�&"�F2���m��SN��G`��6��U�bMYnf��bv��Ã����\�>��0��k��t���Ѧ�:��Me�;��8�lޅS5v��`m��W��V���^;g';&li�q���y�uEC0i21^z�]� hٛ��[�h��ޖ�����!��D�yB�(I�3�ݮ[�ֳ��j�ٞn��wkMY�Q=����ZX�����I�Ji��c���]>:h6�.�m�u�]@�n����qͷ.#m�軪����NH�Q7[���=LuaN��l�9g�V�6��6)��/^���ٓ]e 9�g=&��f�@���g�s��L�g=�p'6��J��Ս��l�\v�a�\鲷`΍�����k�W۬��ש�Wvxd��F��P<E>@CB"g�'�ZUh�>�/���OP:��E��EA*(��WIALCb�*y%��1�cm�<k-�
���#�+=m+=[ulΨ�j��U���	uʞ)t8��I5��T�bʄ�̄F�6�䘺��)tJ��,F�{@˹���7eC<m���LpܓW#�d�Q�&�O�gq ��x8�����m�9R�k:����z�F�B9ꉚ#�@��b;f&fL�V0��3�ᵛ����MZm��H��N�I�^�wt,���?�vǲ�Z6��dK'/Ys,�Kp��mm+�Cde"[&^�Ӹo���X�pJ��SC �ݫ=��7?r9�D}�?���ߏ��o��}4�Gk6�X�X^�6��W���#�s��3�"���SB�E*���i��`y�i�|��0�ۋ �����U\�56�r!y��`yf���w�DB�ǳ`g2%-�������SE������c��<��l�L�=���@Er�D��..1�3��P���v1���xp.�b�5��$�=���}��2��Y����<��l�L���,ݛ�����	*��vS ��dB �D! ��H��)b$�qҟ����>{����׀o���[��GQ]��,y�,�76lG"̝�`bǳ`i�M��ڬ�;���=v`�mX^�6��!fm�`lf��!��DM%56�-�y��ǳ�36��:�����r�yl$+P�j��<����2=��&�����;n�"L"�s[�#ix�c�����\��B����o~�m9ı,O}��6��bX�'��{�¢�Cșı>�_�]�"k�^��������f�������zh�%���fӐ�ș��>��6��bX�'�����r%�bX��w6����bX�zjޝ)�e�W&�����Kı<�{��r%�bX�g{��r%�C�Á0&!= �xn'�3>�3iȖ%�by�wٴ��/!y�}����A���\��N�X�*'���6��bX�'���ͧ"X�%���o�iȖ%��BdO_߿Ot��5�Mz>�����¥�ֵ�ND�,K����ӑ,K�S��fӑ,K��=�siȖ%�by��siȖ%�b{�v�욙2b�x)e�ucWa[r�C�F�����^G���v&�6��vt�Z��O��^��b}����r%�bX��]��r%�bX�g{��Ȗ%�b_��u��K���?xc|�*�m�K�����/����nӐ�Aș��?~��ND�,K���kiȖ%�b{����r%�bX�=�yfI�դ0�Y�����Kı<�]��r%�bX���m9�ı=���m9ı,O{����8���.�f��,��n�m�ND�,��������r%�bX��w�m9ı,N�{��r%�`~f����JD����]9�2�I�@���P������}�~�v��bX�%�޳�Ym�Kv����g8�Ż���/�'ı>�۴�Kı<�����Kı/��u��Kı*v{��55p���-���p6�3a����6Ҳ��v+V��D�a�����0���J�q\��r%�bX�w]��r%�bX�g{��r%�bX�����r%�`~���?_t��5�Mzo�~M/�&��2���r%�bX�g{��r%�b_���iȖ%�b}����r%�bX�w]��r%�bX�w�}�5���K�&�jk5�ND�,K���[ND�,K��fӑ,DlK�뽻ND�,K��{�ND�,K߾�9����Y�̷Z�3Z�r%�bX�}��6��bX�'��{v��bX�'���6��bX�X�����r%�bX��m�\�	����-&kSiȖ%�bw���"X�%��w�ͧ"X�%�{��[ND�,K��fӑ,KĂ��;w�ԥ<k<�'�It��v[ZXh�ĳjh�-k)���������lͶ�G:�e�� ����32כ����	���i�h;���n7'�`M� U�A�n8�yN��F��Y\�4�j�o@��v�lv�rk��!�\�K�gm��.�q�j��U�� �A�;�k��;���F�K���
��B+�	��1v�5�5��G)q�?�$zN��wtg��G�>u�T����vV�K&�u��[�nX`��3fј�ƨ�,!�j���Kı=�{ͧ"X�%�{��[ND�,K�~�f��"dK�����ND�,KӳR���5rjfKu����"X�%�{��[ND�,K�~�fӑ,K��w��ӑ,K��w�ND�r&D�/�3�k5�f�5u�m9ı,N����ND�,K�߻�ND��ű<���n	"���ڒ	"|�I���%r�\�n	 �؝����r%�bX�w��i�Cʙı/�����"X�%�߻��i��/!y�{�����A���9ı,O;�y��KıV��w[ND�,K�~�fӑ,K��w�ͫ㉜L�g��O����
ZՒ�\.�"�FZ�%� ���t-JU�S�1�mE^���- ����듻�^B����z���,K�{�ND�,K���6)Ȗ%�b{߻ͧ"X�%��~�9�����i�����/!y��}�듺{�b� �E�T_*�q �m�Ȗ&gw��r%�bX��{��r%�bX���u��O�șzk�?v�o�z�Lh=���צ�b~�߿fӑ,K��;�siȖ%�b^���ӑ,K��~��"X�����}0d%�n:��;���'��?k�fӑ,KĿ�~���"X�%����ND�,K���6����/!y>�؇��2��rwı,K����r%��*d*����ٴ�Kı?g�߳iȖ%�bw;�siȖ%�bS���d�3���?�,n�8�SF�ԡb�f�m�-ȣbR�ȷ���3%+�:��TT ���t�/Mzk�^�~���iȖ%�bw;��ӑ,K��u�n�yı,K����r%�bX�zj߻-&�����h�r%�bX������?���,O߿~��Kı/�߿ka�'�2%�b~����"x@$/B�צ���֟e��e��{��Kı?~���ӑ,KĽ�{��"X��O֔�F���I	$@�! A�����y�)��L�����ӑ,K��>��m9ı,N��7��5Kn2k&��Ѵ�K�FĽ�{��"X�%�����"X�%���{�ND�,�2'߿~��r%�bX�~��g5.n�D�/\��B�������ι;�bX�*����"X�%��{�ND�,K���bX�%�N�-��z�i���ύ�17%[��N뜤��aj��9K�t (j�u"�v��Ȗ%�bw���"X�%��{�ND�,K��"X�%�����wy�^B�}�}ء�HL׆�Y�r%�bX�����=X�L�b^�}�ӑ,K�����ӑ,K��{�NAlK�����n[��l�5s4m9ı,K����r%�bX�}���r%�bX��{�iȖ%�b{���ӑ,KĽ���7Y��a��5u�m9İB�����ӑ,K��{�ND�,K���6��bX
�T$X�@�Dc�P��Ț����r%�bX�:MK��	�u�fM]kFӑ,K��{�ND�,K�O�~���%�bX���ߵ��Kı>����Kı<��_�!vi(۱2�n��/g��ӓ�9йF��0�bLL�F��D��u��Ѵ�Kı=�{�iȖ%�b^���ӑ,K�������Kı;���ӑ,K�����3Z���E�ɭf�m9ı,K����r%�bX�w���Kı;���ӑ,K�����"~ fDȖ'�v��[sSkWW3Y.f���Kı;���ND�,K���6��bX�'��xm9ı,K���m9ı,K��/r�6��\��sFӑ,K��~��"X�%��{�ND�,K��w[ND�,�"w���ND�,K���ź�3SM�3Z6��bX�'��xm9ı,?��߻�[O"X�%��߿p�r%�bX�����Kı>@�AN����D"1���u��Q�f%�KEDᵶ8��lA�-�d�6KY�J���`�nIt�4���c��ƞ���L.ځg,z����#Y��)ʬ��0%F���b7W%V�꺔���a�X�u�e�q��P�Z�;3�t���P<l�pv����Po`8��yo���@����lV#�ډ�x{amaډS�E�-��jV����zSW[� h4vq��N�$gt����l�� pf���ac���X�`-�n0l�&�]��Q�Yٮ����]O�`atz�D�,K�����r%�bX�w���Kı;߻�`r%�bX�w�w:�������?{/��p�P*���m9ı,O��xm9ʱș�����m9ı,O�~��iȖ%�b^���i��bX��|e�Թ�fM]kFӑ,K��~��"X�%��{�ND�,K��w[ND�,K���6��bX�%��v��f�.�5�sFӑ�C"dK��~��Kı/�����"X�%��{�ND�,��xm9ı,N�ɓE�a�SY�]h�r%�bX�g{��r%�bX�w���Kı>����r%�bX�w���Kı/O��vkV�i����ՋI�6����ވ�9"m��tVL���Hx��x}=�>�a�p%����x�,K���6��bX�'{���r%�bX�w���Kı/{��i���������"��3�N�X�%����6���!�FE��	��`E�B���@��	!#D�da�]�ڋd$���?��~蚉by����Kı/�}�m9ı,O����r'�2�D�?�����f�5�ι;���/!y;���ND�,K���`ؖ'��xm9ı,N����Kı=�^'��A�
6g\��B����{��iȖ%�b}���ӑ,K��{�ND�,Ȑ2'~���K�B��~���U��Z�W�N�!y�'��xm9ı,? �������,K���߸m9ı,K����rtצ�5���I�~�}�g�0�V�k�<�;���s<�C�BZF��1�4S5lt\J�B�V�z�E��?��^��ק����"X�%��{�ND�,K���[��"dK���߸m9ı5�}�>��.̵EY��5������"X�%�~�{��"X�%��{��șı;���ND�-�O�>�ߛ<2�HƢ���zk�D�/��u��Kı>�{�iȖ4^������IC)({�j>fk]�>l����1�$�.0��$%�_L�&�s�\	L��5�kf�lf�@��R{8�IxBx�-��M���T�Ĺ H_ ȧ(H
�M kd�%5���H��67��O&cNQ2�����`�Iԏ��X������l�!��;g5�)�؉GP`@.�
h�&��#Bi6\�IN�k3� D$2�C^HȥL���9	�dO	��[5	��=!X@Ȧ�ZP�&���|HHF��;L�m̔�H�,��.��b'��I-4,��I�a�xE����## �M��d#��n��h��Q0G`��U �Uj ��������z�~D�O�0�G�U�*>.�Q��<����ӑ,K�����"X�%�罽�[q�U1��_t��5��!z|����=ӑ,K�����ND�,K߻�ND�,K���bX�%��e�Ԗ�Z��ۚ6��bX�'~�xm9ı,C߻�ND�,K���[ND�,K߻�ND�,Kú�Xm��ڌ���� ������m��XE`�j� q���h��6͢;�=ӑ,K�����ӑ,KĽ���ӑ,K���o�iȖ%�bw���w����/'�����D�C�듑,KĽ�{��!��L�bw�w�m9ı,O߿~��Kı>����[ı/��I֛ٚ�5�jK�kiȖ%�b}߷ٴ�Kı;���ӑ,K���w�ӑ,KĽ�{��"X�%��Ʃ��dչ�fL���ND�,��~��"X�%��~��"X�%�{߻��"X��" B	��Ba  H���c6x��t��N���m��B�����}>4fc-vٝ'"X�%��~��"X�%�{��[ND�,K���ͧ"X�%�߻�ND�,K�:�?y�&�˒ja1H���U��mi�XK(��^�1+�Z�g��x�f�h�����^��צ�7�����"X�%�߾�fӑ,K�����"X�%��{�ND�,KϽ/_Cd5T��z��������߷ٴ��,K�w�6��bX�'}�xm9ı,K߻�m9�S"���w�����p��N�!y������ND�,K���6��b�b^���ӑ,K���o�iȖ%������}A��f��g\��B��2'�~��r%�bX���ߵ��Kı;����r%�`~A`�D����6��bX�'��5{�kWVi�-�[�6��bX�%�~�bX�'~�}�ND�,K��xm9ı,N����r%�bX��wm��P�Հ�BT���4�	S-����-����{n�3������f�3+QB\��iML\AoYp�i]yWMm��:Vga�ٸݬp�q�l4�\�%��mi��L���b�
q��s��j�vMg9�,]�wY�#�[zx� T��lx�q0�f4ݩ���(]��\˦�i��sHg�\[<�ڃ�p�tg��a�+ۓ(���Z2���VV6�0R��S�δ#�B��u�J ���t�v��ջ\�9��I��͸]�n����ޞbwbPd
kQe���4�N�Os/��u
���O�X�%��~�fӑ,K��{�ND�,K���6�Fy"X�%����m9ı,OߍS��5nf��33SiȖ%�bw���"X�%��{�ND�,K���bX�'~�}�ND��"dK��O��WV\��k33Fӑ,K�����6��bX�%�{�m9����������yı,O�~��iȖ%��>O�bG�֍�PY��5���{�ߵ��Kı;���r%�bX�����r%�bX�����r%�bXϽ�u���ڪ�l�rwy�^B����iȖ%�b����r%�bX�����r%�bX��{�m9ı,�����i����l�2�pf�s=x�;l�v����kk��Q���l��豖�rRX][�kiȖ%�b{߻�iȖ%�bw߻�iȖ%�b_��u��<��,K������Kı;����Zh��je�k5�6��bX�'}��6��P��%	D)EF�	�%S6#���rk*$Ic��Ɛ`@��#$MƳ4ɒ�	d��_D"yĺ�=�ӑ,K��=����Kı=����Kı>;_~���MC!��'w����/!�|���bX�'�߻�ND�,K���ND�,K�{�ND�,K���~S�U}���צ�zId/O��fӑ,K���p�r%�bX�w���r%�`ؗ����r%�bX���:gr�&��7%��ͧ"X�%����ND�,K�{�y�m<�bX�%����ӑ,K��;�siȖ%�^O<����m�3��,�m���-֗���e�5۶+�W\T��b`II[\��*�f�I���6��bX�'���ͧ"X�%�{߻��"X�%��w��Ǒ,K�����ӑ,Kľz}�L4�sRjkY���r%�bX����m9ı,O3�w6��bX�'���6��bX�'���ͧ %�b{���e����ֵuu�\ֶ��bX�'�߻�ND�,K�{�ND��H@"@��q7�w|�ND�,K��=rwy�^B������k���g3Y��K�,O~�xm9ı,O���6��bX�%���[ND�,�̉�w�m9ı,O�j~�KMjc3SV]kFӑ,K��߻�iȖ%�a�Q����ٴ�%�bX����ͧ"X�%�����"X�%�ސ��o.]�6 ��j31sb��:oS�������[�jO���� ���{��zX�%��w���r%�bX�g~�m9ı,O~�xm9ı,O���6��bX�%���Nܗ5Y���sY��Kı<�]��r�bX���xm9ı,O~��6��bX�'��{�ND���^�~�O�\b��=����?/%�b}����Kı=����r%�bX�g��m9ı,O>�{v��g8�����B'UN@�
�g�X�H'�}�ND�,K���ͧ"X�%��}�siȖ%���B��B�
�$$��d�h��XRR X�T�$�k`F2�YH2��0����c�� ش!R @��r.KjK)@�Hѵ��%�	Ih�E����$#��Lr��kR��4�g�e5�?x���/>�O��6��bX�%�ӿ���L4�jkY�h�r%�bX�}��iȖ%�b��}��r%�bX���xm9ı,O>��6��bX�'�S�o�췂�vdս�F�E�a��3Z�[�ζ'l`)�. 5"Q]3`�ͮ�J��)��?^B��b{����r%�bX���xm9ı,O>��6���,Kϻ�m9�B����{Lo��g.�\�;��%�b{����Kı<����r%�bX�}��iȖ%�by�}��r$��$��Oߩ,²䔗4��H'���A$N{��M�$O�<Ͼ�m9ı,O~��6��bX�'�a�}��]�5�3�N�!y�^O���{ND�,K���ͧ"X�%���w�ӑ,K����iȖ%�b_=���rf�3%�f���Kı<ϻ��r%�bX���xm9ı,O~��6��bX�'�w��r%�bX�v!`�B ��P�C��|�)�[�Y��n]sc�����ɸ�f�v��.G����wbj�v���z�����I���S�Ʊfc��F���h�\Re��3�9��A�2�Kmu�	��xg�c�ð����	���@���W��m�R�����+�
���x�p�n�8m%�/5�9�1�[G\6�T����X�k��)n�_6Zn��x�wG"L��3��'I=�;�d/�OB�����7��CG[��JfX���c�)���sqQZ�M!s5�.6�%^�]����T�,O}��6��bX�'�}�ͧ"X�%��}��ӑ,K��>�siȖq3��O۫�#��p-��Y����X�'�}�ͧ"X�%��}��ӑ,K��>�siȖ%�b{����Oӻ��^��M��|�Vb�ժ�fӑ,K��;��m9ı,O3��6��bX�'�}�ND�,K߾�o�~^��צ�>?}�!q��C$�siȖ%��F.D�]��6��bX�'���ND�,K߾�fӑ,K��>�siȖ%�b_'����.]L�kX\ֵ��r%�bX���xm9ı,O=�}�ND�,K���ͧ"X�%��{�siȖ%�bt��rɒrZen"T�ţ�6�RQ�<��u{;�x���E�3�^-�Yr`2X���Q9j�/�&q3���߷ٴ�Kı<ϻ��r%�bX�g��m9ı,O~��6��bX�����uO���kr�rwy�^'��{�NC���H��;G�2%��k��ND�,K���6��bX�'���ͧ"X�%�}�I;�%�%ɬ̷Zͧ"X�%����iȖ%�b{����K����=���6��bX�'��߳iȖ%�bw�T��e�&�֛���ӑ,K,O~��6��bX�'���ͧ"X�%��}��ӑ,K���}۴�Kı/�|w0�9�E�3�N�!y�^O�{��iȖ%�a�g���[O"X�%������Kı=����r%�b[���'&�[��p%�9�Q��h�F�R>��=��n�t�L�.T���!��Kk�ѩ���kSY���%�bX������"X�%����iȖ%�b{��xm9ı,O=�}�ND�,K�����.9lv�,-�/�&q3��]���8����*dO�w��"X�%������Kı/�w��r%�bX���;M��7G;@�N�;���/!y<�{�fӑ,K����iȖ?ï�]ڬ #"���Ƀ�h
v.!\E� X�5�FRD�̒Tȹ� �(�*�ߴb	���<�u�?kiȖ%�b_����r#8���/m?����R�DԵg���@ȟw�?M�"X�%�}����r%�bX�߻�m9ı,O~;�����&q3�ui��F�l�E�Y��Kı/�w��r%�bX~ `+�w��m<�bX�'�?~��Kı=����r%�bX���嶘�.?��U�NN����2��VnP�Thͯ#��jb��a����%��
�2���zk�^,K���bX�'���"X�%����f�ND�,K��{��"X����bC�ڑ*�բ�;���bX��}�NC�ԮD�,O���ӑ,Kľ���m9ı,Os��6���Ur�D�/���2�2�.sD�t\Ѵ�Kı>����ND�,K��{��"X��b{�w���Kı>�}�ND�,K��fN�3Rjd�f�����r%�bX�ϻ�m9ı,Os��6��bX�'�O��iȖ%��N�J����u $��W 
 �y߻�&���צ�5�����!�	W"[��ND�,K���ͧ"X�%��ӽ��Kı=����r%�bX�߻�m��B�����}~�l�6l�j� ��ke��%�Df���eWv�&t�6��R��pqQ@����{���Mzk���>|��Kı=����r%�bX�߻�mD�,K��{��"X�%��NϦf,����֍�"X�%��'����i�Kı/���[ND�,K��{��"X�%���{�i��b�ź�X�Q�2�$c��/�&q1,K���bX�%���c�HdL��N���Kı;���6���&q3��x���B;nq|qX�~`dL�����r%�bX�t��ND�,K﻾ͧ"X��F=����r%�bX��M[��̓.�kM�kY�m9ı,O~>��"X�%����fӑ,Kľ}��iȖ%�b_{��iȖ%�bh�o�*sS�f�=6C�A�	$��_V�S=���;�,��o�x%�� �_ �w��������d��'��6G4n�4�t��8y!>�H>��5��19���4��CY7� X!% �@� BB�ը���Q��	�c�"HH9�����/�Ěmf�xg��Xx|ޘA����D� �BH��C�@���-$%��"�4eX'����c
p�+��OB�6�$d�9�c�� ����� E���2*�L�3�Ϭ����Hm|M{)�0x|��rBRFHD�/�䐎0���H�D�G�/�!�$Ry���}9�9���y�y�c�q!!%R+X���|��X����6q�W�9�!w�^�=�X�@�̤����G�,&q����
��^��j��� �|�9V�\�8Nk�q�eR�.B;�u3˅0��)4sI�)�=��Y�S^oƳ�\��g��al9���sy��YO?Kzx�����-����PUvʪ�5�Ue�9Yh)e@PB��V�J��WT�WUUWZb�̬��RԣvĢd�lQs����4�,մ8��gZ����5I�{s����e��j���E�kl�:WN�8��|BN9!�v0�v1n	���&@�����mu�Pzկ"�3�PFA�;s�U�Gl���ڞ��n1i�G[���`�܈���%^ M�5��z�M�I��Xؘt�iod�dǭ�w=cFR^�Y�0��F]�Ʋ�-�X`i��i�J�XXq���.e���[5�]`�W5��6�ml�*Q�7&�lggΙ�l0�s�%�#o8���7=g��عv6n7 ;��T��u�&������E�،D�Dl��n#m4-֘�Y
�K���#�l�9��Nr�
z�E���r˘��8s�Ѯ���"k.�l�K�����#�md����l�l��b�ޅ�y��:��\�p���oi5:U�lq��rȦq;�{.�{0!��/nۃ\��O�c��*jzɷ5$�9w ;�i㜑��n.��6%5��=Q�)X-�[�d#�+��b��6�Rk�Ҩ�0b�m�4q�B�r�,�۳s)�9�[p�,.�s���:���f'��u���xAc�;t�8�hQ1�<��b��n!�V�Vqa!��d��`��V6���p��,t����"�oeĂ[i�;�1�ǚ7q�9s�=���%P�]i
�t(��ؓ+�<�۶��,u���G;M!���m�)�F��B�S;��,Z����Oi���n-�{�����vLq�0�-�I�(۩ֳsG<��n����^�BZ�����(����;:��("��Q&J����\6ұ[�5�x�|��q�\�pD��c5�����+v�ln�s$�bƝ��^���;���3�4��@��b6�;ۭ�I��'GT0`ۖ�����^�M��*��Ό���M{��-�N�q9��mr��[[S��j�����V����Mp=�t�=;I�l�|N��O�=z|#�*'ʇb����#�pZ�O�OP�N#@;��t���A�K�e&+��-1l�\ԅSX�K�����K:ڃ���^g��lZ���/`ezv��V�(�6�`Z�(@Q�%��,"P]`M�[JfX�E��+4��!�<�$�wBF��r�X Bb��Q����eɚ��&�@���\qH6։)�����	[Vᧄ^Ԋ�7E�̗6\�+���q�3	�����m9��M�n�����wOΝ̏���mf6���e�4�A&�V΋�˸UN,sʷ'Um��"�P
a�:�:~ޚ�צ�?��=��9ı,K���bX�%�����L�bX�;��6��bX�'�o���f���Z��O��^��ק�w�ͧ"X�%�}�{��"X�%������Kı>����r%�bX�y�_GLl,�9�2u���/!y�{��[ND�,K���iȖ?��Dȝ����ND�,K�����9ı��?_I��Wh��v��'w���K���iȖ%�b}�wٴ�Kı<�۴�K�������ӑ,K��;[�'Z˩���h�r%�bX�}��m9ı,?o���%�bX��߿kiȖ%�b|}�xm9ı,O���By�4�u$�mnm��v(z�89��FY�<�(�]�������u��k��v,�3{��y�^B'�����r%�bX�����r%�bX�}��)<��,K����iȅ�/!yg��%�e�!�v�S�N�ı/��u��=P�9���mȜ�baϻ�iȖ%�b}�wٴ�Kı<�۴�Kı;�4�Oā��pV�s�㉜L�g���6��bX�'�w}�ND�,K�뽻ND�,K���[ND�,K����8�Gy\S3�N�!y�^O}��6��bX�'�k��ND�,K���[ND�,ߏ��iȖ%�bw�����Yp��"ι;���/!y?}���9ı,?�W_�~����,K���p�r%�bX��{�iȖ#8����������K*q��Q���X�@
CJOQp.S6|���'9�k.�5�.�v��bX�%���bX�'�w�ӑ,K�������DȖ%��u���r%�bX��>����J�/\��B�����}��ӑ,K�����"X�%����nӑ,KĽ�{��"X�%��v������0�����g8�Ż���Kı<�]��r%����*�}Z�A�Ȑ#(� ��b����K���m9ı,O{�ND�,K7�L�uq����O��^���,�����nӑ,Kľ���m9ı,O����"X��dO���ND�,K���4UZ�rH;^q|q3��L�}��iȖ%�b|}�xm9��~��0���<{��7��k�)B[!��R4\�y�`c@�M����VlPڷORv�!B�lvq�Wm�<��ŀw��X�7^ }�ۀ��ج������*�=��/��s�s���v�dc���׃�)y#��Z��7^ }�ۆ�,p�������~�h�3E)*f�Gk���p�{q`��\[�_>�] ff��ܒp�}��X)J݈�9n��n,����>ٺ��n��CZm� Q*����`Ռ�B�3��Ր�.4�X@�k�J�tL�GFU
��X�D�`����׀{v�^���=��.�j�db,���:�`�����w���"! ��j���d��R�=ڰ23ś�BX��X��V��jbJ��ギۀy{ۋ ｸ��n�^��6���EM*J�U�R�5�ŁܖՀw�0�q`v9ō��-b�p jUW-��^1��U��,�AV��bֈ��/�-�Fs�d�3��vv�]Vn�s��6!��=0�9�W5��@e�R�T�nK�'I�rFlx��<�5ݒ��t�nn`i���'n'��s��P�j�����1�g�p$sX�tt�7&�tb��'�M��/i|�W#��X��5wMs
a�#X�fњ��Gk��<_t�p�j��3���,�G͵��-#��׸�i�UZ�m5�l/f�6o41�ЭK��t��03\�,�m����og�� ��n,����7���S�Ȭ���T��nl�Ł��q`w%���.q������V�݈�r�tݸ�=��,�nl�nlr�Q.	±FՀw��X�۳ ��v`��ŀn��aUtj��e�`X��X���;�َ��؈l�0�{	�\9��we��Ė֒#ێ���rhԸ�sv����n3���ҡT�'�6a����c���'�6��X�Z��8Q�0�{qa�ũ ��!HH����E��%�� x#�����߷͛�y|���>~ݘY��\N��Wx�j�`�wV76}��{�`bp�l�YM;�9T��`?n���ـu�{f�{q`�Vj��8���Z������1���<���h
�q�`��@EJ�v�+�ݭ��	�!aYiL(յѴ�:�Q��oO!=���Y���c��=�Ƭ䶬�5��5�b�jY�w��Y��ޗ����`uz��pZ���EL��,����׀}���/�Ďj�,`���0I�	�0D�ژܛwŀ{�#��\�(��34�>^u��,�ٰ=��,zq��
=�9j��8V�xϫv`����k�>��xۼ4ʅkr�5#+�q�����lEI���.nM�=����K��xY����xa�N��Wx�j�|�b�;��xޛ� :��p�i�T5x�A�]� �f�Φοk�]ݸ��T��^W��a��9^��k��������;ٺ�?1i��H�u0T�4�6��ڰ1���<���{�ĹW�S���y�����)B�(SU`{1�X^nl�X��Ձ�V�&¸�8�2Z���&t,ug�ka�u/K�:�4&���--�M>�zWz�$qk0MMG�n~�X�L���?���s�1�������\��Tʙ�Vq�,��3Ł�N5`w%9r�e�p��`zn�����;��x۷L ���q7UED�,�����,zq���,����m���j�H�!*�Հw�u�n�, �Mۀ{��XW8���X:X����); �x�[&Vp�Nǐ)��bg�1v�dkd.����-ƅ\�)��4�,��Ʊq3�E��������{��[���-���]d����u2����m���]`����,�[�؀=qqGX�v�����89���<G-��Y�ˤ-ět	Ɵ��nJ�V[U�F�U%)�ǝ0G`�F�P�k4����ڊ���^&�-�r$pY$�;���1�on�pC�\�m8��OM���v�s��Ɂ'K�-�h��<�RZ�Ed��W�=�����n��wr#�3%��4[DT�T�"�-Xޛ� �����{^�����I6{c?4)?'�JA�[�k{q`{ӍY�{wn,0ݫ=��U��� ����׀}����7n�Ok����)XIdrJ���,��7k�7/U��N5`�߷�*0�P�]�h`֨#����
�9�����z��c�rN�2ETX�7Vd�V��́��ŀwƭq7UU��,������|��_s�,#R��(���K���y|���>ـ{����7n~\\H�ݹ�ErR��&��Ұ1cٰ:۸�xn��Ƭ�T:ILTTT�RҰ�r""�w�`��X��`v{^ wE��V�R��,rՀ��Ƭ�q����y����>�ֶY��-h@9�q�4ձ�.
��u�.$�[
3c0IP��jk%��u����`wӍXm�X�c�=�.�B���@;eXݞ׀}����=� �������Z�J㍫$�W�}����=�Y���!����#�ÈG#֕*]i1!aNwp_Ij�S�}��"�䗫���R���	������J��K	���|w,n��`���$#�x��!o	�2I�i!"^0�$�1�Ҕ�� d5M���k��BV=��M/��-
ZJ���K8W[8��B1`F0�(��n@1vVP�b����FaD�ml��@�Ip�S	:���p�5n��� Z�#�R�W��@��[��������JJI9�JsA�{k�)Qm����t�Ku��G���!�I�Y����HX1�Ќ%o5p�,y��j����)�a���0l		IaHZ�)*@���������֊J �K#�]h"�XV�r� %%�$a1�"FHŕ�
K�.Kl$�$���6�m.���VNk��6��u���A�I ��! ���@9���+,�ZԁYA�.�a2����Y	Kr,\��JS�YB���A�0֣RP,����s�=AH*x �� z��E��+�H���qD��S�H�� |��>g��Q_D��~�ٹ'�g�]������N;S"u�V w�\����>�����ŀt��uUSR�UU`fc��;�Ƭ��,��uv߹���N��K�5�kI�PrV�%c1Qr^n�s4c�
�������q�D�55Q�3%�:۸����s�7w�,��W��J��Z�)�}����7j�m�Ł�e2�<�b�ՊYE�Z���� �����n�[w��F9F�%N�AE"E
j�:�{ذ36��:�2��o9PDG�@�,&@!�\�� �ą�s������ ���un������[V�9���@7�`<���<��lS�2C[O�*�0NM0x�ո�e.�XrT͢�²�Q�c51u[�qל��T�I*fET��֖����y�����׀}�5�L�&D�e0��uG#���X[�6�^�r#��?8�������In�w�, �wm��B^ݭ,�{Vn��&+�Q$MEMTX[u`u�q`�:�31��7�*���*vZۀ}����l{]��V76�A���P����y,��nss�H����`��C50*d�7(�J�� !�7�t��c���Qyv��&�vU���.�w�X�G"��B
6�\rqoj�X�l��q�2��.���n��
�1��JN�v�6^�j��]ڗ7=��u�Y!w.�F��Gu��q�*�l��ܸ70�׵�{.D��=I��5�[�Z����w�n���KTJ�X�+5R$m�ڬY�SV��rf ���$��2Α�֛R4�d�)�T\�,����V�r[`��r���p.k����C���"�Gc�� �����=�n,��ـ}�t�=��܎=�
�J�3ŁՍ́���u`g���e�l� ��v`n�0�=� �������Z�[d,�*�����%�ݫ p�Ձ�����m�ϺV���d���&������ ��q`u6��:۫Ǧ2%�\JGK��,������F9�����܀���HD�V������⒕�	x[T�����-� �n���������Pa�[��4k5�rN}�}w��W�s�\�2�j�;�:�31�XyR�!:쮧%�;^ }�� =��p�����ŀwg�� ;���U��8����lDD$�����X�mX[u`{c^L���+
�6Kp{ۋ �ѵ`mՀ{#X�Aj��*RHۈ�f���\�y�ZS�����wn4����$!ة$�-eMVQ�vʰ�7^ u�V�u����m�ŀg19�xMD8Ւ׀y�vg�qs�M��o�{^�X�m^�"9	d�{Q"&���Jp�� �7��;��X~K�$�D��I$��NJ����I!ňDd�D`Ȱ��$��6�!P��Q'P�>��y���ܓ��~��'���q[U�*�����K�O߷�� ���1y���X��"�b�L�B"�*j���Kj��Jnl0�V�� ��-l�㥨��F�I�:s1I�Y<i�;f7Q�ʂ���wƌL���lv�ϻ� =��p����M׀���]��YEd�`�y��Ds���Xs���^�D$o�֦D�:ج
��-�7�<�M׀o���{n�y+��A��A55J�y�G!y��ǵ`�:���6�H�(Oa�e�����`�4�@�]�&ƄM"P�@������.䞾�e��(8Ւ׀of���{n��׀{v��B�9��@AȪ��(��lS)�M��ջ�9��ձ;JDں�ORtd�2�d�;)����n� �۷ �{q`��n�j�R��[�?Kj�;�Հ�ŀf����LUJrUj�W�{v��n,?qr"Ձ�;��h)4����n��� =��p��x�K�M�~����~��Eeq�`�c�b9�OW@�{�`?c��=�DD@�iRP
R1�R�"�e�,%������~����6jg��1�:.ۭ�XHgH�ctvMUT.��[Z�e��H��
��6R��T��k;�����,�q�s��#k�M,b Ѵ�@�K�⒦���Ak����h>���C`�n�F:Z��.��k�l��D'��۶�0��ŋ��mZV�J�Xf��qm��Z8�;8���_��ܳ��&�&�����N���[W$t`CxW��4L�T T���7Km9!�:��k`G���&3��V��т������`a���Geb�K4p �Vj/����y�[�~�vz�ۍ�":�l{V��TM@T�)J	��Vr[W��G!#q�ŀ6o�og�縛=�K���Ed��X��,0�V��Vr[Vp���D�e��A-� �=����훯 ����{��S��K�JI���j��Հ�;� �1Հ��[�
�!��ID�P��	J1���`�1��]ͤ�A��jP������Fik�Xر5+�-���Xa����;��4�ln������y��ĵs��P���7&n}�nI�罻�s���ˉ&�z���Y+�� 7G�`78ՁܖՀ6�X�F"&�)R
�&��n[Vr[V�����9ļ���o�n�K���\n	��Vr[V����X�sv߹�$���
ie7{�i��m��YŜ��s��V8�3.+]]�[ix��^�R�b�dUK�wj�3u`bm�_0��/�;�i��"����!G-��s@yfd��֬<�Xf@�-�N^�Kp����Mׇ�\b&� D����Q��O��u���߮��u��
����Yf=�mX��s�a���W�wf��j��R�*�T�Q*iXf:�7�Y���^��0vn����MH*lٸ��SSnM���'�v��np9*�˖��lE��	�����N�p��� ����=ٺ��ݸ�~m����
�U`ycs`���ṑy�z���HϾ���%�]ն���`b���<�XM��=��S	�N���t%� ��������۳r@�E��?lz�S��g5�ߵ���_���p�d�`u{n�M׀{v�~ݘ{�b��A��wh�[1��S��K�H5t�*r͘��(F��WU���x䰖���x�n�,n~�Dr#�ǵ`{��@T��,U���n��7^ {Ƕ���x��^��c�:���rڰ�X�ڰ�u`bȇ,L-�8Z� {Ƕ���x��n�ۦ��dZ�\�ePl���ڰ�uf�%����c��`v(S��\�J���y�Hx���)��6d��M٪zr5�	�x���y�)�����N"D҈&,O���ŋ��{�����BzR��!'1|���@�����F��]v��IR/�ɬ�q�B`4a�I���w�ɣ��K�y�l�|H�9/��l�@����B$7���ߵ�y����SՀ̷R��$
h��� \9�����z_MhCA��ܤ�<�H$�
����e �5H@#��%���T`�r�e4�"��ie	��NL3s2٘�O{�D P%d�8��/�y�.n����h�b�s�\�U�J�n��ի�����>a��w�P�4�l���<�ݻ��/^�w؃�!�ɹ�%�}ԣ�.�q>���3ׇb]��&y=�G(����|�uLV)9���Eժ����\㿎q	YN�)nf\�/8�.,\�b����i��Խ�����	A��<�O�x�L�� f��"M��JS��9�{������yͼ�Bao���1�YI�ly��h>����e��&c��^}��0�hI�r�+K���Ub���N��^���{
u�F�; �yr,K9p�A�+����X:]��\��Ӕpư�7ty���r�?I���ߖ�V�P�UU�4�@UU��U]�Q�In��TL�6�c��W,Tb���(���57[�-g�ϴZtcx1v�I�Sh�I�	v�/��27��8�v�=.��"���]��xCr ��������퉌�`ٰ1��T�44e�5���-�\H`x�n�WF�������������ƗX�9�ƫ6�בԠ�؍������	,%h��ۃ�n��������q\�ήț[1����`y�%k���猇1�#eѦ04v�L��`r.�&;w��`Ѡ�6��c'[��=��d2�� 
kf�^�UO:@�����YCY�ݶ^�R�J]���֕���g���61��/ *.��Zn9��8�ؗ#�a���A��<��b՝�jM09��x�U;��q�rxn�(b��m�ţ�ͮ�Baۍ��T��t���s\�G�f�-�6��@�d���q�/M�gm�왤:�aB��O9*�8�$�4�z���מ��MM�Y���cI1.�	)e��X��{l豕���;O)��=[,�NS��:ֶ�-�wW%�����.-��S�ux�+��Zzv�۱�,�s�v���Fx�TF,�̸3*�4��`�w&�ͥڣ4\Kk��y���7F�&�Jᳲ�۰��2Fě��g�y����;F�D&6-W-��;g+cm��;8�ʛ�/�g�{�m�'�K��d��v1�آ�t���&(��
�5���/s\v�fy6щ�k�r�˻���q�8Ƨ���Gg�/l����N�����]�L7<k�F)��b�ڄ��L���������A�b�vssV-U�,�9�m���e�5��������㫋����ʗ�K�Ƃ\j�61ז6(KHc).���5�cM���Q-����!۝"�c��:M�X"��]pkq�+QI�\���$lDV`�s��c�#KӺ��h{p�ey+a�I/.d&� a�HIA1u�]��{x���ZCo*=�S�1U�SAur�҃a�;�N�����PR�� !�X ����A�*��x��*�ȧ�Q��x.�O�����}�h�%�uۖ�\�$!����ʐ���{&�zs/G-�*���8s\�6-��m�3uʄ��j�bX���%��t��p��u��`5ъ���6F[u��K���m�4�k&��ç)v�����<n8m�plY{�]�e��Z��أ++��c&�Re�
B��ζ�1Ҭ�E��.�m�zz랉N�J��4!T�0��ն���m#�3p�m�CR�;[�����t����"\P�M�\GcrFA�INKH�%qy��,6���̦@��lY���ؤ3 Ō�*JPMMR�{�Xn�`��Vd�xy�7Y5Y䊺ۀwv����7^ {�� �n��l�xL	L�`q���mY��Hy�V�~�� �x6V�;!U� ��j�3�Ձ������t�$�J^B�\� =�ۀwf�����ޛ� �}va �&�v>VY��c4�JMi,s�a�m&L4���i�]��Ÿ�����q�Q%�vn� �m�=���ݸ��ݨw����k��y������ā������,g,3鿕�w�`y�e�Ȅ��C�'��eq���������;�t�����[Z�j��F�,��<�Xn�`q��7���n���l�/�uN9]	m�;�t���2[Vz[V0�A"*'�ҁNq���8,f9R��+�=�)��`˗��bmJ�v��!�)����-�=-���s��DvC7kK �0ؙH����ۀ{�u��$�f�~��s���1��Ds���kj�$IyUr��?~x�n��y��G�#�s�q��z����Xx��V�Uq�v7+�7�u�|�����<�uX�#I3\P��d����dc�c]n���;��k����|�6�v-Z]Mx@�i��mF�/��el���e����n�5ǴF�9�1���UU��[Vd�����8n����*�2��%�����?q��{�`�v��ڰ;�Ċ����U)UM��76���y-� �7Vp�LeD�U%�@%4�69Kn�rN���ܒy��krx�$]��8�q�HBA���h8C�q���3���������Z48����� ̖Հf7V�����V�FW�Yh���r�#A�4�Eޤ��v�]\�� ���.�����7fW��ými�6M���u`7-�*r��h:��J�,�5����q6��������s`bȌ�*f��ML�@���1Հܶ��DD%�wf�ջ�`w�<�MQ����)f�7^ f7VM��cXä¡D��S)A55J�3���������N��}?Ny�.JG@^8j�RcM�D�3eZ2����b����m������+�l�(䖑�]�	|Fu�i�&�ۧܛ%������z��'@3p�xX���f��Ӏf�ʹmF4[�x0��usM��B0@�KJ��ǫTJ/[U�L�2�)�FlMr�@f���Z��wCl@Wn����R�n�pЊv�f�Aq��4¥�G?84"'�� ��̓
�s-�7Y���l�2~8������sm�4e����jb�HG䭒c*$�W\��������pٺ��ݸ�{�U
폑�L������r9	����ڰm��8�ۍ�!qB�J*HRT�V�� �n��s`�:��u
(ayUr� ��n n�� ��տs�N|��շ߽~���2����XmՀ{��n[VVc� �-"�h��U��RX�R��8�˜v��Fܪ�e0���r	��=f�2�L�U�w�:�t��1������jrC`�VT�Kpݺg��s�9���9�b��`��`�X�SQP��F�-��>}�� ��V}�$y�j������x� �*�SJjeUM�6�XsVn�`u{6`�#�t!]��0D���� ؎r9���@�ǳ`�V��D�H
���n6�l�l�V|=.(�E�*p"�v��H��+���T���e���s`�[Π<ٵ`o���j@���v� ��ۀ�ۀ{��_�f���;T��FJ����v�����.q4qDF0AlP=��H!��Qs��K�s�?;�� 7��p�xP��a,��In }�p~ݘ������#���ڰ1�l)��A<��P����Kj�;���7V�`���5n8T��e�J%�K���4ܰlI���B6��4-��ܬ08�Uxã++P��	�V��V�������s���u�^4N��`�W+�[�wf��܈�$�mX���:���74����,���n����w�n�۳ �y���݌���R��^����I<���rO��}��^,P ��8`&S)T W(8��Ez o{�w[�{�u�K��ȚuQX������_�f }�p��x���$o����j��兖�Y��
���UU�ר�eA�:����u{Kv�hXH�[����0�/m�7�u������P[e�6Gc��%�܌u`<������Ovoc�Hl�aJ��!5
TUU��wU�wٷ ��ـu{n�tZ8YdmK^ }�m�5�v`�^ہ�%���o�� ��D��V'r�\��_�� �Xcs`�:�;���I�Y,	 H,9�8$�b�H�.��5lMIdE$	k��nkWa���X��d��ݚ���C��G'��[\���.���X��=��86R��\�!�d�nn�b�A�qlR�>9Մ��=[���V�M�Pc^��[z4�Ɇ��V�p.���]�T���MQ�!��M��g^�6�Gm���`������q3��FG����0�3WϠ�9��p+��iH`�.�]LW�Ns��^\K�����Ё����EY�-�^�g'gF� U�v��J����SJ�`��T�J ����Ϫ�k� �c�_�f��OLu��q��*��cs`�:����;��Vx����"	R�Y�{�p~ݘ������0}���Z5U���nl���y-� �c�ޑd-�Ȇ���9,���� �M׀{�p~ݘ[�֛mh(�7Rb���Pjŭs�
n͝�84�ƅLV�Q�tc�Mu
T㗑�YSL*���k�y�ޘ�|��=�y��5T�dE��ֳrO��}���OA��q
r#�1�yX�7V/c���9Ȅ��1;��r�G%�M��|�n��l�5�v`tDݵG]��Vv̀<�����s`5�͆�^�{6��_���2�eV�ݞ׀k����x��Cu`g��D�X�4���]��h��L-K��l�!4̴vX��1E �q��,*��7k���p��l<7Vzq��!�I�T�H�j�-��}� =�v���� �nV���m�DE��f }�ﵹ'�g�]�8z�| Q��ʔS������Z� ���of�p(ٔ���>��nͺ��p�bȐ��Ḡ�#���JHp��s$5�fh*aj���M�Zr2a
{�lX�p��쁽��ĐWfU2&br�km�#1e��	H%�BfC�)n�F[@�$�E�c!v�ǚ܄a�B0����$x^?�"��Jc�!� ��$�	��_'����ĸ�J����F,>m P�aIR�0+e�B����&2��б$��B����1���_����@�!>���Z���T}3��H�� ���t0#��c53L��1X�"I4�i�Ѹ��㖻�KB>zM���j�m�ZHK�4��^�'$-�ofg-C�kL!*�t	79<�K�9����K��hᵔ��d$a��eˉ"ɖBs['8��s1��HCR�ĖR$�/#H�=09�>%"�a%��f��&g�]h������!$�c�<9�`h��	���%�1I�9ÿy�HI/�6�b���)�mo��݉���j��f�8yx!���d�n�%�0�$ !IS[!&��8[�6dk$!N=+� }�?(�*�#����;j����$"H���kf�f��!���d��_��N�����|{�9?q�)*i���ݞ׀���:�9��s��ٻذ7e�AQQ2T�!
UR�cu`5�s`{!���q���ob�IP���XX�S���&8zKh���E�1pɁJ�W����u�1��B9\�9n��ـw�w����qq|����p�D�����xT�`��q`y�2�;�Ձ����7uEE�:���/S�`���{v�}ݘ|����w]�Q��+)&� �7V/7;@���ï��`��&��U�(�$	a���`;#%�P�#�Gc�kFC��*�QL����ٹ'��\M�Ŷ��j�-��wf�G�\�V�n��נE��2��d� ��:���qv]����5���N%Rr��qn�����s��؈�[�Yk�����;�����lG9@�wU��B�PL�(T%U6��W��G8�y�Հ�wV�G��{R*�K$N�;^ w�=-�2V9�<��;`���9%r����s���� ݛ?L�=� >���>�f�%��xT�M��+�s�Xq��1y������.!rzn�F[JV�M��T�c���u�%��4jFѳ��F�͜�՝�� ����1Gl8� �:�i�R�p��u�Z�a���c;��Fa;�*n^�Ʒ d� ��\��In5�ɲ�XV�Ĉ"755��������,�nզ02��Y��OX����{��d��a�x�D.�y�)b�,�5˔cf�`F)n(k�\u�i·G�r]i�s�A��{I���-uf�l�Wh�Xw%;�{M8M�8�h��`Ŏ7V��ml1��
���UF�%����wn��ـ{��f��밤������,�n�^nl��s`y�2���H߽y񠩌��1��m��﵁��6�S,�n��q�UR9[��ۀu��f��� >���wv��mB*-�M�0�S,�n�<�X^�s`w�F P�_�[�@�v���.��tj?���i�K���ѣ6.�m�<#{k�^+���Ͷ�nՀg����l9Ƭǌ�i$�W� =�ۘ�]���O�0j$BE
0�V#0!
�@I*@��=~@Ca�G�<���nI���n�wv�h����[l�Ui�n���s�X|�Xy��j&��"uX�#� ��k���p�n���{0�ķ�矛���TV*�.�{7j�:۫�8����X<�ߋgv�jj	Dv�AKN�i�q����fB�:"�wk�8��Ene�pҪ*j���ڰ=��́�8Հw�����h��5��m�}<�`�Ƭ�n���\p�Jp$�
mj���;��x�wn&���8T|����1� �#��O"'��V��`c'TR�R"�;^ }�ۀ{v�}�w �t�;��f��э��q�p�nՁ�,oUtn��y���쐒/�(4����l̼�;�k
�N�C��-���=�8&
sR�UܬH�[o�ƪ��e2�=���;�Հ�\sr8Չ�B9+�}� w�� >��������ʪu�0w���S =����Kj�=��X�L�1�4�mn�V[p�n�ޞ�0{�Ҁ�$vU?/�A�M��pl���NV�Z�z{jl̦X��Xrڰ>���=�����[dܽY�>';d4tc�ˍf�fk+��F�Əl+l��r��4��%�-O@n^� �����;�r:��{S`o�o�
��e�v� �wn�ḿ�8�l�Ưy�D$dcP����ĕ*�L�X[�6��s`fN5`���>��:[l�et��}9�3'��u`u6�����ܧb�e��f�Ok�wv�=ݘvـ���b�Jq(����L�����V�ƀ�w������]����^-��XR��\����,H6��e]�Ӟ�Š�]�Mط��Ӎ�[�k�U��*��]P7���C��c5���c��\7�>�rq�e\]*)�m�M,���k�����;P\lu� �df��1�N72I�����f�]��Q�=bR�y��炲�Fu�w��u1��v���`�q�ŲƲS3?��U���|�-�d���f��5-�qQ%��	e��V�u2K�`Ƅ�43�2Ĭ�5�2{m�y��շ��́���Ƭ?nށ1S
d��i*����<����1́�j�;�ۀoOi�2�N9[�Wm��l�=��X^:�;�ڰ;���$�E�F���`��� �}� ��u�}^ـ{I�@��J@��׀n:�;�ڰ1z1́�j���6sH'Ki5-	~^?�t��j�U�&��qC�������F}xs�^�.�xնI�tP�v���`b�c��8��@{^Ձ�"^�)2��Tp�V�?k绣�}$���kNQ�P�$vmLLvбXp
@j`�#N~\Dr"�#��|�������lQ㏎�����`��� �}� >���=�{f��ʫ*�K�YG4��Xq��3Ӊ́�j�ǷDE\$��V�[�|��0vy��;��x��� ��"`��D4mF!Mm���6���`v�V��\չ���QԤ���e��f��=�}1� �n�䶬���H�$���H)R��3'����:�`{$�0i=���Ԥ+���^ }�ۀs����4Hi @�B�4B���H@�AeR�D�@�0��V�5�d�ٹ'�Ok�>^�L�-�qH��-�>ٺ�d���̜j�;�Ձ�"r]!I6�����x}l�7����n�{7^����Z��	�P���%��L�akW:hU�"YejS; b�\a�Vn��h��S��2�[�7,��7����p��x��`�ܪ1�FԼ���]�w����`fNK��X&<l�9h�mUe� ��׀{��fo�n��wn�7Rng RQ�;5J�c�M�{6ݭ,��X_#�{�Kl��0���4y���wrN{1�(=���hӣv�۷L �۷ �ۛ2V9�69��=67ЦUp�B��;d.��]�v�;v���Mv�';9+5r, r��r�c`�Dдs[o�y���s`fJ�;�DGP=����6�t�B�Jj�M���Hi��`=���;�Ձ�9.�Jf��J ���=�c��X[u`bm̀�cj)��	��[��q..=��?�ݫnl�Ls`u㛨&���j(���� �c��9�[�>6MTI�=�f��PEW�h����DPEW�Ƞ��EU�("��QA_�"�*��@�� �B� 
� *��E
� `*��D ��EV"�`*��@B�H���A
�@ *F"� *X
�
�B"� * ��@�b*H
�B���B"�
���H
�"*��F� *��D *���@�*��F�"���@`*��"� *
��, 
��"�
�`*�"Ȋ���0�*�"�
�`��"��"�
�@�"�R� ",Ab*D�"���D�"���F�"��
 Ȁ�H*
A?�U��("��QA^��*�U�����PEW�"�*��U�(����EU�("��("����e5�>P��"`-��?��������=���ASꮯ���Z�Zk��%4Ӑf�R֡@H +�Zh2�R��i��P�� ��5@� s�[�   
( �    �@ 
H
    

  P        υ!P(�R� rwG�=z�1 H
�)R ��E���A���=��0���x	� �z7�⻻���)�[ٗ6�����>�m��� w����Oz�{�9����O{��(��{9w�����g�}�}��_v����|����HT(��N�zo���{�o���{ʭ�n{I�x��g�]g�9�=��v��D�7c��=��*��g�x��}��{�R�͞A�hg�}>�������&�#�a��������| (�T�@((�2�|���>��ۢ�@�`;u(5�F���y��� �P���6ǟ`�X{�(C�8��=����A}o �>w1�c��xk�ް���� �=�����t{g �G־�B��I"�T�ERTP���(�|L�v#��7�Ҋs��R�.��)Ҷ������ܲ��sK��m�}������E/�yN�ir�li��޻���v(*�t��Β������_{6�ªl�ҥ[8�m{4�gEᲫ�n����t�]��^JJYҔ�wu$���i�y�)GN��Jh�=�#��EH�RR
 n,F�t��;�����N@{ܢ��-!�2[�n���OA�ǯl ����Cx���<��k�d�����7��^�ٟ{=��ǽ`���T    �  "~���IJ(�5&  �  ��R��Q$�  i�42i� �EI�(# �0��L�@��S�22bh2h�L	��4a
BMJ����h �4�@Ed� h�T�OI�i��<����e���3���bO'���s�<��Av�?�O���U@O�*�������`���H������y	D+�AD2N���b�EQ�P91** ��?�*�G�*'���s�����{wwwwwwwwwwwwwwwwwwwwwwwws3333v�wwws3333wCwwwwt7wwwwu%�������ww{����$�n���wwwwwwwwwwwwwwwwwwwwwww������������������������������-�����ݻ�������$�www���������������� �` ��ث� �@� �@ } �Hت��	� �Z�9�{�l@O`�� � �*�� � �@� �@
� 	HJ�} � ���@� � ���� ��
{*��{*��	� �Ҩ�H䪮@�ү�� '� @	� ?@	� ``� ��b ��D�@�U�@�W� >�� � u*��� }*�� @�� 'Ҩ@� �@�ү� �@� �J�� �RԪ@v 'bv*�`؀� ��~��9*�� N@� �TQϐ�g�Hr���C#��Y��\�r~�:~�(f����?Y��k|+�9�pᛈim-��[��pY�Ë���ħ�of�h���v�n�������.6�N�(�ժZn��V���5�����l��fi*
q%�\��a�@8$a�8��)��&s*��tW�	�P{`��.���k+�<���<��46W���a��]�W~�t)B�:����0���B0B���<�I*� ���8�)�F�7�[���I��#
��	Ùn��L�e�F����m�<��f��9�D����)�A�2QJ��ȡ�}�(�}R�g�*Jh�N�ۡ1˘a�Ѫލ��d��u�d����EQH�\0Uӽ�:�(R����8����!Ǣa)aj�bJ�9`�x��ŗ��p��[����|���iŪ2<�}�BM�rb�0tʱB볖2��j'x�]�q9J(�=]�7r�6��ȜqB'7�p���E��� sT�z�D�z�ވ篵9��~���i��>a���w���Y�+%	|T��j��u�gX�*��y_7�<�byŨ�<#�: �0�[�����2·�爫��+v����8QTU3�y�Ш��!�D����ri��ú���2�M4�G 4n^��r�~�w�#� ��	wE<钳#x<�
���įK�u��xyT"���l��[۲P�H����I�/�������[ׄЖ�,d֌	'p,2L*��g�v������g`F���형��on�7τ駔U��%����j�^��jr�f���E'A��>���o�6m�1����t���-��{�[�ko�=�F�l�//JR�^N�ieO�$�R7��B__j��.����^f�fn��UU��U�+S�{iP����rjL��wia0wmL�	i;gs}��3M�Z���Ou�=횧7Nq�wI��.P����Kj�WڟU�D,[�FK�lr�sq��s���NF�87�����6e��F6Gw�������w�N�Gd{�J�$�
4�ӽ��˜�S��g6Z��|Ǿ..֧j]�]�}Qg��s��-�{Y�h�o����o����SMl44����f��w=��r!�5-KFS�6`ז�<f's�.MN\40�&�m�)�R�4�8�hÃ�֦˱�2�Z#�|��Ls{���+f������ɚ�♲f�	��8�QS�qT��f�����Y�VB�Y�&�8��2ɴ𗶖L�#zn�E�����f����IKw�-�2��浦��sZ�&'suN8�5�=ѝ�)j��%]��߫++]�8!�\�_/�vu�]|Vv�����:�{+V�4b�����&��k�M-�m{�N\d�1\L��9��:e����	
�;�{����'���**��io�(f�Y1g%o�֟S����=�L�ow{�Ҵi���=�Z�Әv�{�s�<m����Y��GL�h�3W�z��m�	��4;��l2�Wu�^�Z���*;�pUAQ\_J:��J�g$v$I2�!��;�o�	䎯An�H]d��n����6�s	\[���-ޗhԇR��VKGH� ȭDZd�Y�7�v�/uU|S�)r�������`rC.�m�V*kF���k�K��cU���!�4CC%}]@�f���|�{����<=}MM]�2��Bm��X���X4V4�#Mp�Nq῭��/��]�	��>��e�\��*��&T�1փ�u��r����� (�>J;X?���H���ˢ�ɨ�0�,m4En0`��i�GF������9n���t�&��Q��ݖU80n
��E(*�U��<�KG����Bh�#��2�_*tU�$�\�2Xs=�Z�wL�9̬�|l5�d��c�3�qʰG{�zH�w��%�w3���2a�kqt�L�kKy���C�kxg��*�L�"s{R�����x8�N�;wݧ9���s�	S� ��pb��/oN{F����{�ޥZ-�]W��P��	�+ʿ�)j&Ӆ�nRil��<^)#�&��J�DA�IFS�S�ze����Ǆ�&�����萶{��!�X���k�Z[kk�fjVpd�S�S�����M�{L%��<s255���3E�'Y����z��~�b�u��*OB����T#�Z�N����r����{��r����c7�vM��22n�2P-Ǘ
^R���&�����J�9�]E��I���r�W�RN�ݱvw�*���EP#���D9i9_Vj8Z��Ĵ��x�����Zr��6>d���DLX���cR�&�7V�@kF������ǘ��4�t]����*�c�A	QR��������7FL2ZA�
������>a�`�h�4ѽ>i��P�a�̓;�=���O5�n+"��,��L�ea�h�Fo>nT�f�E:�@Q�+�v���������뿥��]j-}GL|�y�'�8v��Ʋ�����9
�y�\d)}s�5/:˽ŹP��ʖ�C ɾ��书���֓���:k��ۆ�5���"�tÇ�O���Pe��6���G�1٭�6���o)�xnN:33͢3�s��'u�����v12��3�͌�˽��kZ��chWy�T�2,�u���҅��\ޱ�A����w]�i4�i9�f��^�cOH�;��󫓪k]�}��y��cִsɐ�oy8���8�z��~���;q<m6���M�zt����w�p��������/��E���n���mޅ-��q�Ch`�2!�'3Dc�]�Kv�����`pL%;�sP�p~ש�9�j���iRx�޴���u0y'7L"n�m�
��#�Qk���^��V���h�Q�B5_O��|��S_E(���}��dͲ�b|���)��T�%��:'+�]r�6i�L4��6�e�*0�L{�ØoP�{�^Vv�0��P
�f��f�kW0�w*�����rQ�)3�3�CJ�{�fH��<���Ȇ��+��SZ�˥��L�2��pmFIT^��\�(��P�T����s�X���1s��:���O�1�6T�nŷ���D�5J�R�[7
f��7�{��ð�5S�75Q���S�W�a3:���1�cDAFD�BV�\�#����9�\2xu��<,��ȏ����ucg��L�.�|<�gOs�z�Roٗ�n`�w�<��F���4,͘��AD�bs�\�6�z]��Cp�omJ�7����bw�{������Z�)y&h�D����ܠ�4�
�q5(b{aݚ;���{�d��k|�y֢89w9z9�5��W|&�4lp�q�}s9���޸�s7�#����H&D0�QXp.BIi�s�u��G}1��NVu�9����s���k�f�z����wlz�5��zM	��IWc��%I3�P`0`40aɞ6�w�(�h���%1k���f�N󆹿�"x1�<Z<Z�HY���v��"����.�B���TT��w� �����i8?�ֵ����lg���8�Q�Mv��"��j�G�:�\��!�L=�|跲��i>��]�i�x�]_0yBuQ��y�5��>����-�O8���3{G���[��w�Q��0�y�Y������r�hy��ﷷ:9]M�5_�ߦua�ޛC�����k&����k6���E��.=Ij�r��-�lɚ���\���w|N�k\_fh��5Ѵ$��Z�w�K�Q>�&9�`Iu�0��,�!��nd#��G`���^:u5/8�䙮zu��a[�z�7�`�U�皚�/b��!�f����s�V;�E
���b�7*뽹z�4��h���ɢo��}�s�x�)�ug9��5d�9��9�0��!��J��*��	Ieʻȝ0Wi}Ѭi����v?f���.�/=�g���{�����f�I���o9��wh�KpS1셚�t�݌�ù�1�*�;�.�g����ݺ�����M�؄�˧t�q���޷�c��eAA�N��W��s\����f���5k��!$Z�m1�#��42Qځ��Pt�190�ر�S[{���j���������7+T��>��ޕ}���EGݙ�¼�I���:]��{o&�r�ji��;��rr��;�eg
^F��."s���[���18��jr[v=sJ��A�o�z�o���9W,m�z�Z�F*��nCN+}�y���ĜцhZ�5VC\�Lh��<�]���؎�1ӦH#1#�Ō' ��Nխk��Q�N2f�l��8�Y�
�880l��Ǫvl�B��ҝLnW�2��9������,4)��y�d��Y�7�ΕM���8�9�dM�2������M�&��>uޥ�y�t>�ﻈ�b�,�tQt_r�.�&6��z����UH�B<O[�����t�Z]�ZǾ��xy$��E��]�<D�^Z�nt�ʳ�S�G��NR:0���G�]�t�'0�4ܐYRB1anO%=���!�&Ubs��5�e����R+�&��yG9r��恲Y�=�&��8�k�JO�.�]��+�"��mkv��V�Tlֵ�4��L�@,Xv��e�\��W�N&��蹚E	��0������CHc�F�=����@����i���kvpWW. ��P�$��W���g61�3{a/��-]���q�My!w��\��9���a
',i�c�"bwa�W�e43tp6f�`��aþ1;���0���[����<��%AuS쪲��b.��E>�	� �6��:f�)�.���[��8�o�<lס$��{� voh�Ko��x}�ڭ�%�*ߊ¯j��Z�hAP�<>����yƷ��d���]��-k+���?�ݣ��Td\@
�2�¾T�`+�W5]`��]S/�T����jX[�K�&�7!�\�>$�v����.��~�Rb��˛�٭����o��>�k���cv�7�2�s�{�$2��޶܆ѭ̗P}m�4����!�_u�����wk\4����=��X߷Ѵ�3|]�5˭A���1���3V@�ы�.k4*�;cH�y�O�������o�����RI����^����(̥���[��i�3�6ߥ+M��}���"~��T��v�6�۲�9t��X����'d�fS��V���`FFY�N�!��m�Xij�
��R{a��X��Lج�b�j�ݮo��\���H��2(�g��a��6�;�(Fԕ`��Ku�2�sJ����KK.��If���uv�U�h��0�������#v�q��E��T�C�K�������M���DL��k��������J��J�Z��K��\�$�J�����U�������������������������V�ڪ��������
���������Z������U�������������������U}PUUUUUUJ��UUUuUUUUUU*�UTUUUmU]UUUUUU]UUUU*�R�UUUU@UUMST�UUUUUUUUUUUUUUUUJ�UUU_U}UUUU[UmUUUUUUm_U��UUUUUUj��j�
���������������Z����\�d��<��+v�z�^ &+������J�mu+��tY�{����+�0mXћe��5֦L�Y,��k�/�ˊ݇q�nm�R5�cdke�"|����=U�ܫU��ƹ�.زd�=T,��&�k��沬����pU[�+��n®Ʒ;�R�Q���`���l�-��
Kn�A,��Ƥ ##�-�����+ֺgr��WX�V�,�xΩ�[�-"��DU�c�`��v������V����v��ڮ�ҙ	�"㕌j2m�1�ӵ����dҝ=+���a6--�n)
Ա�>cR��F'^�.���͊��@&=A)�h���q
�D�z2v���!q��%4i�v@�`΃m�7A���e��K�muE�`(�u�wK���ٙv�Wl�tuu��%��*�֮A�\u��5�V�99ٰ����h�5n6�o\	��k�76���R��΍��G�K��|m��u	��Z깵!����Z�GV�K��p�v�Me�WUp�m���X��n�b�Z���<�<)��g��ȲH�Z�jN;��󴫰݅!W;��孼EV�skؚ�[��Cv9f���j�vۧ�8p�.l�=<�硪�=�e����9�43�T8n��͇���1��q6�����j;1�u,A���G��w���ymJ�?��~��s�t6B�K]��d����nv��ݑ�Ӧrb2��)!��B8�W4��d$�W�nx��.��8!��(�a.!-�%���{gۣgcx���7;G��	�Pug��N����H��1�[/P!F*^Z�y*ݸ���[��gc��l���`�3[/��n�Lv�Sn*zP{m�6�*���n��Ö�vZ��N�l��ܯ�2�ǋ%�D�Y7g5X7QRpz��ȯ��/k�.wQH���dx�o;<�v�4�Oݵ���e݋�fWy���-<�������V����UUUUUmUUUuR�UUUWUN�V�j����d3���v�۝�Z�n)ح��*����R�.��	�7�V��Lb]��J�[��ڛN�X\+�:Re}�Е�����	�30�%khjjM2%���c5�6�v�N�Q�4����3����u�lc�6�F��*:Xvݞ���uc]��i�.�C<�$Q��^�6�3s�,�����[��j��l1�Ș�������.(G�v��w)��kK���8�[e��gG�fآ�`AƝӮNp��#��t�u��Gl��1���x��i۷�X���* utq��7mݱ�9
�Z��
��Q��6��I��^ۇk�h)��Se��2Y ;�ͮN����;>؎M�<��w�5��u�=r���d��M5��з�kvg����#m��f�J��`<	ӳۍI�岕�E��-˪�����e��'y3(Q��\�6�y^c�W���6նpB�0@��L]vԁ��m(�wV
ն��M�#^�d٬�s�YA�dƈ�;)���<��{	J��6�/r�..���C(".�v��4�@T��9���kS�Z
�֨�r=S�Y`B�YlƼ�.�[4�u�z�0u����^�����f7Hm;]m�b�Z}]unf ��H^��;p�ŤF 6�Ghƞ�h㶝Pۅz�wR29�n��ݖ�rM>�τj��;]��U]�E��ngn*L���rJ��ڻ��G��9U��n��X����y����ru��F���c�be�o<pU�G�l��*����*f����pBK�Lu�{����t�ܪ]j��O`	xr�-�Up���B�w�~��ʜY��M���6R��*���ɷ]�:�iVm݂�;U=nU��*�����WK,�3v�\V.��T��6�aM�h�.���9���X.��;Xۈ�l]NY�*˃��cQL�C�IrX��.�qn���L�f�Yk� �����ݡd9�!h��D��)E���uJ��b���2n�C���<�yƑG�K|v}���<�u�dQ�r�ꭵ*�f��+r�؞m�;�c�Im���$�7U��%μ�Uqm�`�6�qR`�&��,D�y���Ĥ�4ꃝ��Q��&��PM� ���ݵ[S��L�����iJ�';��f�xnsSkn��ezyj�� =R�s�;l�EB8ib�;��3f۪�G�7]��x炪�!*��vlv���lm�әl9C�㦲�[U[Um/+Ų�ӵS�:DwX�!��u���k�b����k�>ح�V��[V�j�yf���m
�[K�N� P�n��D�sCmع�:昝���\�s'2;l����m�enȪ�
��j��	!���W�j�� +j���ݣ G-@;�Q�rwT�UE��b��8�����ه��p�����R�QB�j��mmQ����2�F�j�ջs4�S��[�x%��Yq�)G�F���x+��:x=�q���B�d��:�8Y�-UƑ#\��R�2�歫v�B*�yMtuؔ�v����k�,�ԜK-����
�� ��ɱ�յJ��e�5��m�q�8�k�Ʒ/���@U������y
�[j�n�]T]�ʶ�UX շM[V��%�����ܷ�Rf]�sv �ڣ4F!�d�p�S�n!�دXv�ժU�PM�tVp�Uϲ�a��1��HM�-���i��ܨH����;�v��s�J�Ud^��57k�-�����җfF��6�� �6�ƒ�<���*�k�kv�(��|��|�Ԫێ^�g�U��d�1��Z�M��>�eɴm�n�j��=u\�^Lm��#n�!Z9�A�<��n�,��/X�m�2�;���r�ҵE!�g�d��H0"�Zg[_�Gn
`]v�R�o����j��%ū��6
駵��h<E)�p�#U�v�8@GTTt�Ԅ4�V��+] gg#T7��=����v�K6�U�MT�UJKt;�-�݆�3���S��m�[E��V˳��Ō��9��m��m�.<�6{aT63�Z�p㪪������������^[����m����ںe]����ѣ��8�X*ۙNW�[*f�u%��r�[uGnښg��W��ܴ�- S�nط+�EU�q�� �N ")�cVܔQ@+�0��*��:��u��612Z`�q#j%r�(����w�_ie�nV�w,�q�D��:ͬ�ui{'������{�Ľ�X�^Y��Vf�:eۮ"��h��@��<ŪO��V�un1#�A�%��M�\����}�O�«ʹ��c���b�U�ię�j��`$sUR�6�[�:�H9�ͳS֕�G6�	q�s;hvA�Jg�l���9�F��g&�W��s�dkVr�m�6Gtk
҄7�s"����Ni��1�nM&�UpTlmuR���g[�ǂ��]��B�<s�뀮yZ��˄)e�Y�������H��u�k��++�s%�يFX��΂e�f���e���ڞ�;�h�U�����s�S�fK�#lWo"���2�c] 4늱�S3Au�n�KZM�͋2��it�砥3g��,�%�.H�<TG5�Eo�z��On�Rq��֪��Ɲ�M�9FX��Y[��aj�3��[UG/l�����k��[�F��q�U��
#%]1��٠NtU�U�]UD�X'j� 
u�J��UI������*��k&V���ڪ�[k���u��sm��T �ìWA�s���8*�D6\���l���)Ǯr�n+Vi�ʏ]f�`m۵���A���-��ۚ�rΞ�R��j�ij@q��Ul�]\ڞZ{�\ <�sZ�c��|�\p �g�U�� ���3�Ti���m �d�iy�@�����O|I� f��;0�s�t6�3�l�u�E�^^U���kj����uUu�OV��PGA�����A^Z���k��E]�媡L������N�Ԭ�VU��w`�n��˲�.�n�*�*�Py��U[Tvu�5U�K��E�GYd����H�᪶�
X6��=*�n��6��mݳ�YGGk��w/\�XŻ]P]5`��n�ƔkW���ڲ�F�\ѵs�m$�ʄ]0��J�qO�i�=UJ�K]c�UͶΜ��)�v'��X7YY����<nư��U�� /4����5&�9��k�����D:�%�n^�v��u	������l�UF��P��n7(�պG<���\�wu�4J�y���;@.�\[["�6P+�͢_=uQ�����q1�Z�x�kTոڇ�r�/-���}nUW}Ⱥ�1�����s�4jG��
�?���*�/��U ?j~����*�CD�K�Ha	����$&V���f�B�	��f���Y��	�d&ffV����Q�+�DH��@WJ�P��A�@0�\_�BO�
iU�(nF�++ �C�av�~�LC�+� 8�% �]�E��	�D
hW��
*�P���%�j�B��Dڙ���w���}*�x%ݶ8 v�ʡ��>��������x��=> �=GP��4��"ʰ	��HeBz2�'�N#�$Y�"�M�Q�>�.8��,����1ར'��AD�^���B���ބ��8(H fHa'����"z��x!�N)�����xi�����L�#*A1\P�EP_C�|�a��		�1t��N�"!�"I��r`x �����z
�
��M��@6�)!)b)��G}������$D����!��={%3A�v$���'��1e&H;P�ot&*qD4������z# C��i��mH�4�8�>t���t��=]��s� ;Q���郶0CJ,z�)ٵ:A�10�#��Z�#�S�6�PM/�}LP§��L����x��Tr�@t�z(��z� ��OD��.��e� A�Q%@�x(CJK�x�$���@�Q⧇P^x �x���*p��Y$MF�� }�8�e �X�gk�h��� t ���*����^$�r����A��JD���P8�&��T=T9�
t�����DDP�S��'w0UU�`��(���G�����s0d"��2
��|A\F�AQ5DEA(��`h�	e�$����@"���DIU\3	��z�}:�ge����Q��SH�xiN! D��g���|;T]+�����
�
�dS"�+jV�����UU@  ����������������TP@U$��%��-�Im�K�?�@��&����C��;�ffbY��- ����D�h�ԁ�h�І�iM,D�T�8�� h�X��% !�PhM�U���b�JQ	�T�[V%4B�%(�݉��S���Ibkx�d�afYR�㕙I2��ѯ��j���V������������n�@j��j�+�� UUUS��j�e&\M�<QtC�=�`;����9�8���D��B��7#A5�m����s,(ʛT���F:YH<�Q�bGLinJ��q�VUt:��P�.�X]�B��Z;�J���=����:ͱ�[���Nq��̇��>p���'Ls�ۚٮ��l�W��Ux[gF�i��ZqV�^�t7T�l����IyS��Pnn��3�S����dȖۄ��ڵ����� �sn)E�\LU%&��[��)c%O0�vpo	uvƕ�H� Ptγ�;s�ک㦪�ɯh϶G���t�:mӭض�<�c&r<3ȸ��.b8�GT7o�E�{�\^��1�fp�^I��j���6�L.��*�H��RQ
�AFl^�Щ��V6�n�݂5[��9�=��֟[�n��m!1���|u�U��Hz;/��n�sF�a���Jx�^��Wm8�:w��NQ��P�Ls��i��YWrt�F��Aj6��\�i�{:fg"� \jpJ��z<�9#v�&'���}�����igs�M(\��m�6���$1a��=�����\u�a���]�紮ǦT�Et�ˠ�ـ!�֤�^�[�F�k��m��`&��h��=+�ҷx�q���(�9e�Svt ��lPfi�7l�<Q�vIrca�9�ܜ��u�%�D����ThF�ukk	K�:��f�ۋݫx��I��f�ڀ��C�&�-�Ќ�K0�R��3L��N$/�V�Ƥ��+��^�9ڗ1��5[�ol��C�õ�E�j��{��Z5u�v�<�Z5�̩��͢��6���(e��:�9�\�B��.I�C]��=l�pC�ø�N�"�i�Zݖ�5Ц��<�-�,����+��F���N_�4��d�@OE�EL����Bl؏���b� ���x��D�U;Ђ�Q��M�DG1N#Èx$Tj>,*�������囂{�.�����r��mәNW)�q��1�v뗀;5����Ф�譁�l����Z�f0-v#f�3�(b���kp���qN�[5mY�A��R �R�i��*e��#�{g��nN��{u v�ufy.�`Y�[�G<�3�y�r<�u�����]B�\��è�.�"�f��	�4����2�-q�e,�n�h�����
�e�qh�R�+J�	��-�i���������_|��s�������{ԕ$��6�T�vY���� /��`b�ݗ�A��(�R	'*$�`gvT ���1wu�ٮ}�X�Snq)V�f�)wu�f�}����H$��D�1wu�$5����fK�\����O��)Ԭ��!ۦ�[���m�k�۪Cf;f|^�(/;�\��������JT�#�}� ϲT�����5�I����ҍF��s�d޾���= {��H�.4���:;�����I9|���n�zRHi��Ě�VVf��Řk��ʪH�k�nl��+�%QV8���v.着f�}ܕܮ.��;sǐ��B��#����7\�����>]�v��x����M��C�u������c{����㔚�×K2mn�2�0L��翚`=/���]�� ��_z�*S$���R���w]�wu�3�=U�q#=X�k��(�M�`j�y�y�fm@�DB$�T�������y{�1���v鷹�ί	Ԩ���)�fk�g�*k��`g^�7�҃���R�QXݕ ���%�{���f������Io��v���z��7��M����n�2�چ����[��wD)JJ�pq�Q��|V�{����U�����ЕEX�d
�q�׺��9�U$j��{��.���H�x�d������V-ն�{���U%�w]����`w([(��un���˽�,�M.��s��-Q����4�owڸ��:�y��`ۜJU��Փ]��s7o���8s$�{��|��F��Y��kX@���ɤ�����/�Y%λ�EC�i�ۣ�87mW�q�n�����]z��� Ż�dK��^$�Dn��� ;���*��q�ǚ������7#M��*��q���RY�|���{�w����`�[\��o�������3\�+ �� �d��L�G�q2P'��y������n��uo��R��0�O�C ��BbQ�g�Fo�p������{.0��4�dnhK+.�d5Z�xL�v�V�t�t=ri쉷nn(\FyN�&�l�;p�黳l{�k��dr)m�ɼ�4u�/@0E�����qN�:=)�#���46�66��q,�v�9�I�{\m1St�V1x&�Gfq�0�U�b�]n���^6k�ؘ�`��U�Xm�_��'2��q/�Ѹ�ts�gK�d���r�^�C���K�s�K\pS��Ұ�T��m�??m��P�����<�`w��P��6�ݕ=ă;�,׾V�� ��R&��N�;�,�Ů�7��fJ�^�TƒJ��a$��r�l�R� ��b�U ��c�;�y[M):�dB�X#5�31J�Z�q�cͥ`z���Vr�T��[�M:��9-Ɨpd�h7,�]��y�|�ݞ���]-;�fl\�qf�7b�}���L���`}�<�ʮs����w�6�R��2[m��{�s�]{����"Ń���BP\B��c����;�p̕3�Zj�:�F�p$���u���� ��P_n;V֍�E�RG���9\����7vT��ˬŞ\̬X�Х"Hr�N�w]V��V��\��������9�r�\WN�s�&T�٭�G:q��	�\^=cmj�Z+��TT�II�LR��7n��f��gvVf:��}��TT�)D�]f,�ꢷsҷu�N��uެ�:D��Q&D)3;����a҃� /D���T�w�ݣ7�j�{��$N�$����u�Z�{�u��R=\������f��I�8�U�{n��5s3�+�������@8*��)n\�뮦r�fSe�]�E���R#SP��c�
�[E�J�8��}Zf��gvVwT�u��LF�Q�%Pr���w�=�s]U�ۮ������R~$�*�{~�������~����8�;&Q�0�����s�{�w��qĐcB`&p(��-�H��#bK®W9]W9�]��*H
'D�.�z�����=�P�s��t�;�S)�#�:ě�qXx�F�s�^q��(�0� ��W:����KB����%D�(�>fweg��{�g_=깾�)y����]�����}�g�3;����%En�N��7n����gvV}��k��B�����N��a�3;���uS�ܺ镺StDL��ەw���hk��tu�ޫ����00  0`� p��q:��ݞ��r@N�9Ɣ�u��2��긼�s��"�������h�fZL�7�x�P(Bm��d�n�v�8&lΛ1��ؕ����[˝�d�ɜ���4e�.�f�h�pAM���a�Щ0�,�KcH���isɻ. w��Y՝!7F9:����;��/.�XL����vy��#;���i��K�G�.MqcF�[AZ]�7��/wt�'�7lS���Җg�Ndݜ�krh�� u\�ݱ�z��a)l�Z`\�#�c����s���_37e_z:ƣ����9��3v��fnJϱ�^�fF�|r��I.�����+>�Uwr����h�ƥD�(�>fnJϱ�_{�u�w_;�emH�*�2��[t{����{�l���U�����]�?S�;sP�\[�\^�]��rd�\�V�!�W%��N\%�0w+�YC}｣���]��UU]ou�����F�mD�p$�F,��z�C+
vBS��2$�� F����s����s�����2ב��\�.U���w}��߻����Y����x�@jQ��몟}�u�w]XfVʾ�)M��A$��i�U���Xw}V��a���ˢ����W�<�k1�e F�{=��v��n�upnjKNr��76*UQNA��9�i�ޜ�3ew�uSﻷY�����fHW��ʷ��>HI����s=u�}�ܢ�3|��QH�7 �׳Ϊw��[��Rg�vP  QwwvP  9�s�UU_��붜L�I��D�c�_g�laX�ܖ6�f�$C Ͷ�4R��5~4JVc�l�L��u&o��dd�l6�[�T1��(�!�ޝ�B4hq	��*s�T�a	���sm��13�Ƙæ� ����p:��$iv������ۺ�B��	"<�]qw�P�:o�)*ǜ|fƃ��աƚ �Y��\**
@	I�0[�q����ف���%U1��SUIP���(��4������\��� ��kto�\�w��9�e��L
&u\|b������E�N>�a	խ0u����>��ߤ<�:
�7�T�Oh�����};p���Dbɦ�F�5k��p�I�xB=�xpը�%��
�щ�L�ѭ҉������xFD�kZ�m%�"i��6M	�a�d�!�xhf�Ҵ�)������l��g�4�D�[p�$�l�JR~��`Ȉ��vgu��1Ͽ���D�����dX~A^�w�  WjQP6���%%H%!�a�s8�@�<�}h e�ث���D��U��������0�D�7���_o������a�,��l�������|����J�*��{��ݣV������	kZ{<��껾�{���y���$w�����!�Cr�A�M��'g����3�v$�fr�0u=h2�Zd�ut�׽���9���U�{�r��������o�|�?qԁf%�ϧ��������߾����|���K}�)I��A$��i��3��]i���{�+>�U4�dm�)�
'%��|���Ow���H�&�~J�0 |�p&-�)�G*����G��ɽ�O�ee��2B�2fE��}��~K�=u]�����שs��V�kBQSP�2S�����D�f0�����Կpɺ��g��ySj�Dv�F����uW}̺ÿ�����n�{I����Uw��^�g������7�9v�Z��"�$��i���wr|z�6Uw�^��׼q��t8�4���ҳ�|�.�f�i���
�����T�Ԩ������U�U�Uw��{���~�����C�D�d�cI�����}�a����y�NȚz�x���������7�����̼u(�[�W�n
�{m��@$\�9�����d�;�,�ᠮ��O�
#�f�������F4^w=&��ɖ3��s©�Y�<]y6��v�Y��suZݭ5�����cb�����0���ٲv����$�P����v�'il���Q�kœK��+	.�����"H4]��ۻ28�7җ���$s:��eɱی^%6�v�Oh:�q�.JiIr�|���7�Zf�~����_8ou�_�ݍ5J���pR^�{�|����;�ڰ����������̐�1H��+;�J�㬪���V{~�׼���w7ʉ�N���U�:��ww�_W��ʮ���fm{I��#M>o8}��]s�����
~�~����S�E^����nV�e����u�vS�1�0P��ʖ��n0W-�‪%)H�m*Dr��s�=�eow��>s���}��ߟ���ˎ9��f��'<�u��vU?�EC�T�_g���{ݟ�������Ν�������R�j��{����f�׌����ow�u��|�e2��[�@�ł{�~�[I���sk���fl�Q~3v4�*r���慠���_s��{�ʰ��P�����A�I����fo�e%�u�F�%������ҩ���s<m�j�e!���]9'M�O+�Z�¼y.bо�ߴw���]��lk��٥E}�y7�B
E9�|�yʪ*����{��+s}/�3��&�CnG|�9���x���r~! t	 /��a�L �1S��U Ťͱa��ߐz�����Q�k���o��j���06���P)�˯��}�eowү����ʮQy�m�M�x�َ�yl�&f.��s��"!${���H\��}��w�����?~X[��\ˊ�36�^�]�Jq�2n�{���f��]f��řџgt��/��jB�jT)���������+=���r��V�,���'A��Sr�ʳ����\�>�8;��������}���R���s2����[˚6��}����k� �H�W�V{��u����n�r%L�NJ�UPs��=��������
�A"H���!ڃCB�����Q�}���W���7�
H�#n�}�U�s������[�zUn�f��][�������GQ6vՆAxn��u�l:=Ʈ'm�+�&�sWV��N�<t#�ۂmH��W�~��~��wӞ�{yUˢ���U���T�I�J�$��w6r�������������gٟ�yʣ��=J�$k�f��u�_{��.��e����A=��������+�h��S��*	�}\�;ܙR��ѹ�;ܚ�F �߻�2s�|��1�0�#��$��{���H�%�~�:�C����y�a�O@�O����6QT�P+�"f��WB��uՄ��и�(Kh�0�v�Ґ��finI�0�1l��hh�]H��ֻ֡&$㗂�������7�N�ȫ5ۗ��~�����۲��#r� :&��9��y���Hm%]C�=�d�S�Hܰ3kjpn�&�nN���Hr:�SHt���͹b*��"�n1#Rn�nPI%�|���7��ۏ�h���B�e��.��&UtC�'�z�
��ӛ�z����F r�(��s?�Ӟ���Y����=�{�l��>>�m%.\n�MH�Y�����\9�s�|��nn����Ef����9\���k}$��R'M������ky��[hg}�HC>��a�xj_K�L����"J}������:�;��&�p =�C 3�s�I
�Mr
T��ͭ���r��}�隙��z�{UT^im/7MT�7�z����,
�&�xyOfۢ��S�=/�����Ҥ�QB�i��s��M�*�եx��߄����}�{����S1�I�9tw���;x$��D�	�!�z������\x=b�W@��1�"���Ai��
lHʄ4ՠ��m�%�P�CU�HYq�2m�*� .��;]����Ww�Ү�����W*�Gw4��*FY���M��������� }���U\���x�ߺ�\N� (�G/y�$Ag���59��&�����Ҩ��~����`�na�BO5���}������U���S���Q����f��̮��!$Aζc�i��9T�.�35��,�������z���U���I�D��S����;���w���W9TV�+;�-��TF4&;��{���@�;߲��}����Q!�OU
�I1"S �_3wӛ����χ
��`t@ �X"���	���M&�T&����� �9U����{������Ҥ�RR$�q!9; X*�9��S�^G~��tp1�9κ��0�^��*	�f��B�U�}���t���f�ni��ܨ�"(n�U)>����h���u��LF�6�R=�3.�9v��wN��)1�0�#�4!s���8���}�	h�o�,��[��H�l�_�L�2��	)�=﵇;�����������&Q�3,1ח*��}��ڿ$�| J{���~��o��ˏ&\���m�����g~w�;����z�)/ŝ�"��8
�
H"	�(�k
��@�1 �UOʿ~*�컯�`P����Q���껝�}�~�s�B�2}�^�������HK����fـaZj����q�Y��9�lSM��m݆�(l���<��Ԗ�a^;se������g��u*��»��_3��T:^���"�nl�*��G{�����׳��s�V���|���$��9�P�7����G�_����f�z�V31��[��_�>D����>�q�y�y�v|�5D�8h<�����31�ps)�3G�����? ���~��z�w��~�?������� ]��,  .s��ʪ�����a��A�Y�� ĚB�z��pٚ��4���������4ظ`�e��a�5���e�.��]=��耡!��ZCA'h��I�A$���GLg~/]�C�-��Π�mw��dp�	��&`��w��6�!��n6��8S�N7�������f�$�ζpd���N�L`�BDȒ�6���d�Wd�ή	qq-���Κ��e��L߸p�QPDA3�p�p��Y��}���y��7�'`f3d�)�࣬��zڔ8R�ʍ������)��	���,tp3�h �sz7u�_G��삪��5��QDS,���*ꪪ�V�����������ں���
VT;�_}��>���`.�Ѫݕ�Vk8ob��ye���\�V�.�0�r��;�"�1�{0Kڳ�7;������U��a�����"��l흹�c�m9�۩���iƩ�t�;�9�7]ru�n0�G ˈ��+u�Lka�"��aۺiiL�#��m�v�seӧ����D.LC�Y�֑e�&�E�$��8�&��;v�L��� v�M0��')�a��p۵��e#��ڡ<�T��[��<�݋@us�Ӎ�IA���s����󣃫������3[�B/eӔ��,�����ҡv5#-���#,��C:��7<Vҡ�t�ȑ�����h��HY�s��cZu��6�e���5:����9ku�����j:Px�'����Z}�ڦ80 ۫��b��3��uq�`WM�ć��K��i@�����g��g��a�#=	��8v)9�pwVb�u3I�>vuVۧBZ��qf1�1eإ#-ry�ו�̚��� �e����t�T����b����]-1���lm�5sN�g�r�O�\�9{X	H�*X�u���)l�Ny����o�v�H�f
7V�`��P���;�=f�&�v����]�L�j{S��)�c�v�q @��xLu��� ��Wj�+�9�����p,��a[Z{秶 �/.�:�]]^�;v���Muօ�\��f#K��i,�������q����Y����1H�5ζ�wd��7S�sms���n��qb�Y���Gqv�lʻ�c+i���M�	����KV��.�;�i�>D�2��3g�o9�θA�;�-�	�i�-�|vw*�L�c]���/*�g��㎹܏]<�z��1	W��j�ʹ/�g=;#;���Vsm9�HLd�s�!��%���R��?7U^�GH��U2�����D8 ��:G�� �� �_��hOE��9A�D�AX� h�~�"�z�f)��%�K0�L6˥���"�[ `v�h�K)�%j�C7j��h�/Q��6 ݴ��,��X^v�	�ri�7%�.�T������;��i�>;r�u^@;]�g@d�E�.��,�v��*j��g���`�!��31n�\rh`y�uб��$�h��[�t��Z�
�=mp���l`�3�6��7���[��Is�H ����4}����@ [Z֘۴��g[Jy�;[�kn[r�����k�N��ʮ��j�;\w���o��wu֕��ߪ�U_W�_�gq{��sfd�7���Q��BT��}�G>��g�{}/��+�n���@إ:���,��wG���a߀R
�����s�!�LE
��IQ6]s�ܿ��W+���<s��J���k��p3;����i	0�$HJD���}��:�!#�����ѿ�|�=�����ڂȽ=��j���l�#h�( W��w+��ѿ;��1sg��L7ף����w6��k��?W*�J��ߥw��tB*��Zټ�w�~~��>��ц(��	D��1$!. `)�aQB3�H�����$�`?�v��U�O~���u�>�d��`�N �|����\g2��	�).���:��K�����ř���}ﮎ���&�̴�d���I��w'9�~o���������}s��ٜ�##���U��UVw��ss|�7�����yvP�N�1��L�-��i�.�nm�+��Iq��.Km�I=i�4j;^WL�YC������y����� ��<Sü�ޟW�H?	���B9|���W9UUE{=�W���;���9�Up��m$:^�)9�����p����C�n���
� )C��;w����s4�h��@���UUq>E_���������߲k�+y������iB.H�*&�w;�����U-ݹ���:����j>��v�[�(�,��q���c��yvK�8�OU�n�5�0���$�ϞJ�t�ۖ\����}W���w��� c��l�Mg�JTN'#u	�����ʪṮ�w;����{�\��9A���QG��Ǝ���=�C�(_{{���y6��nx�%�+�[)*�b)���������'���BB1�
����`@><2�a?�k����O8C�ZI�x��r{�ʿ� ^�����������x^�wVL�&Y9���m��ru��*���,MiQpm31F:���X�t��_ D�I8��A�?͕ ���6���r���n���:/��9PL�$n��?r�_W+�ٛ�Ł���X�I��Gsf��aR�R1J�Ձ��Ł���g���-�� �ڕ =_,�i�)��8���򸻳|��� �rT�8��~,͇�JRnH�A��a從 �����Wk����@�z~5$����ԓ�ۤ D�*�����c�Ln^ ��<�=�0%j�cnsWGg�a���u�<g��j�&x�M�;t��Q�.�KuRm �(��t�m�&��7��&7O7mn�m��T��3��!(w;�hB3*OOi�v=m��y�v���t��h����AJA�K��\r����ok�u�<\���<��X�ʵY��K���[��]�s�
2��l!P�L��t�H�spke����+�.U�L]T����D��v:�����:�>I�)Cr�g��zT1.��f������ҹ��WX{��@7<QG����馝^�f��w��M�ߕ����� ��S*�#2�pЫI�JS!,��+5�r����*�<X����Kj�N+iz�K}���P�,�����,ɾW�F��	�|� r��`g�*��U^�S��N��}���Hy>��Ou���ճh��Ҏ%Ҥ&�	�ls����s�.^�e�n&�ԓ���Кb��˧��zX]�vk5{�����ݕ =�ަ�r��7p�=�7����L�$~�K��|)ί�滷V���]@�l�W9U^�r�7ދ�t��mH�A��>����;�*�UĎ�~�,�;�tku���Iܨ�a�r�K=뫴s6X�|�?s�UW�_�����I��鱺��~��2lVk���P�z��7n2A��v�M&'B�871�N���aK���sp�w{ܵS��ZM�JA��3�;5�%����ʫE���K�Q�Ht��AH����7���Ϫ���1{� f��`w����\H��:/�4�*	�/}�����s?�b
D���a�)��+#��8�L���� -���>�����m�����޻_zJ^DAD��6�7�T�n�X�|�פ��T�{� ~��S�9Dp�rK�y�X�V�x�:�TK�����=�>3��u��Z�(�]�4u��\\�َ:ռ�x׬"�ڮY�Y�\%�Y�?�����щ|�(�{���ϛFc������r$I"�;_ ��S�U�(lUK7k�����X��~�r�^�*�7�
�&B��4��"�{��3vY��8����|�Tib̯p���&���I*��r���O��S� ���qUsk�?�UT�<�8`C�]}��6]Y;,�l��	9,�f��q�2{��1n���=���ʮV׏��e8�$�j��N�k���z���4��e6�G�����yM<[-ȝ6)PL��~P�L��g���>A�~ kݦ��%96䍪��ܙ�~�����o���uO��r��n��ި�a9JH�w��`f�=k�����5��tj��������R(S�K�R����@:�T��H�۞�`��ܐR R�D����ʮ{�̛�}� ���`o���D?�]ߧ>�I2�Ie�����[u��WykcK 4m�Y�њ���b������\�n
m���u�^'�VU�2wNه�㭓٘��� ��)�V�v��6�B5.W	Pfu�q1�n�����J�+  ��c�#�n:k�<�=<f�NkvoI�O-m�5���ݴ���j��"q��Y��Z^.U!�e"����)>�t�t���~z�~YnCkv0�g6���[��`2�����l�	q���T����};}����O-&�|���~���037Ҭ��y�U���P����&��Ȕ��R��K\���U6o��V�|��;��U$~Y[M���A)%��~!�.��P���[�w���mՁ�f�N���9j$�����6�;�]I��}�m�@������b�z���I�M9#j��{���}\����|���Z�(���s�o�M��6s�uz���5�"hawcm3)U5�݆�*R$�pVR���a9��f箬�z@-w�r�V��3��H�^H�5CR�P�IV����?��%(��O���#z����bH`���� ��H%BW(`8����fZ8�D��K11���A�Uj���=.�/��~_��wvOy����
H����R�47R�g� ��(Vf�?s�U^�W=&���X���
�bu6�V�.����%����7����_<�V�{�{� M�)�)�(�w�U��r�}4��z�.�������n^ܗmZ笺A��oJ��I��	f62f���u��۬�X��w�J�>v2Gm=�~ .�|��?��s�Uu�f�~U`~����r7NF�l�:�T���>�mՁ�OI��_���2���6)���Շ�_�����Ւ�?���ʰ��s�ʨ��s�ʫ��������٬ɪ���ل$��37�n1��0cc̫p��"�+,�M��혨�8�7�Q��<t��<"Y�b��033�ΰ4��Jxy@yv��̽����\���dw�p�p�`e�B4��8�i��;ð��c��S��t��jV�E��>q�;�"��Q�'���-f��-]�r@���M���Ho�ISX��PU��0�i5�Բ6��ލv^�m���$�S�j,�: 1П��'�fQ�㦆G�e�䊴cz6�����-�䇤5ѧ�&@zl6��w$�1U�l���:9d�c�e�?a���"z��E(p���WUC����4�0�� �/QPǠh_QSܠ*��c��q"�����P�+�	�6�z�W�'���<�������\��^g��7U�P�*&�����;����`o���q@>]�<Z�Q�R�P��W䅯|���V�3�����}H?ҹ]�ߗ�_�k=X-�k�i�*��i+�˶]n'�轶�1��6���T����l�����5{�]/�����_��Ur�s�s�5{�{��V�)�I�Ձ�^~^��>����F��>]���SFVW�|hM%)�Uv寀�o��Vj��r�q�Y� �=��˵���o!IJIVVj�n�����O�c��b �ֽ��4��c�JM\�˖D�Ͽ45�(�������Ձ՚�|�����o�-�-q&a�E��n��q�Y�JC����z��o��7�O-�Ȗ���5Ư��OŘ�rm��#V�]��3\ �v�m�8����s�^���uf���~>�)#=��£�8�����SR:�T.���}ݞ,�mմ����T��R R�
+�ʪ��y=�KH���.������U ��V:�㕕�-��6��ߦ�� ����5���~��{yۜ[?��2t�Hd�9�l��[��n皼�-�jc[�&��YP��̸K�2�[�����dsp:Ƴ�ރ"���p�%NĮ \۳�G$%̍���a���!�	��u�:��^���l�[Itm�yĲGc��iu��U�ρ��ی�����]]���Y��{���$&�(r�#p��8K4.Ke��mvwlv3�cTy+s�~PI8o%���vwS+]�R��ܱ���gu1I���ʽz����@o�U��Qi�R�JE�?�˫�!`�U�՚����y�m4:^�"	)I+�;�|���q��o��������W����?�n����_�|�A}}�g�r��M�׿]}����`{_��I��D�j���f���n�Xywf�X}İ�(�-�#j��A�$[����ϒU]پ_��j�ɚ��~�����������.����:�"b�z�!���Jf�:ǲ��٩6�vK��5���U�՚��]���s}ua�YY�)"�)Q��`b�(����9U�8����p�c��B!��=_@��W�&�<���RO���V]پV��U����i�Ձ�<�`}�۫=ʤ��|�
�[� �}�FQi6�Jq)�kj���7��_vo��bцUq]�����^C��B �S�U��<�`uf�����sn�7���~�p��3m:NsGM2t�q͸M;��{]q�9�'��yz�F��ڔ���[�K�ǚ�Iw7�^���w^�Xֽ��cR86��l�w�`w7�V��U�՚��U^���-�n�N�G`f�n���=���U}G+����ȈwB&�U�w?�8�~}���Xg�i'"��J�>ǚ���[h>ǚ�=�s��}�ϒ3y��$hn���žP�r��ɚ�5,��_c�V�20m-��ĩ%q��%�6ƺ�DxƐS���fM֎2�U�ێnH\\��f���{����h���o}?$��UeV@����տ�� �6�R�H�����\�r�;�|��[� �jߐ��R^�TT2S�U�%�{�`b��7��U$��ɚ�3}u`n��Z�F��(�V�URǞ�;�|�Vg�tu_�̦Y�(d�b��������k�	�Q��N8&����*��V���׾VV��A��"{�m�b:��RT�q{R��C�dGWm�lj련�́l>I��:�-��6�|�|�>ǚ����U\�Z��5�*�F�d�9*ė��U������Oߦ6��鍊|�h��!!~E�����%)
T�qX���������V��U����SP�M�M&�.��>���]Xc��%�ܪ�
��ߔԏW��Ui��9J%"�;��ua>~�����'/�\�5�<��I��	`�1	R�=H692U%C�9�W���&�ֈ��k��M�+�n�1�Ӑ�c���N�����n:�Tv��'�^Ͷ��I�(r�7��<V�E],s�{$r�=�sO)Fۛ�l����]�$��6`ʽ��;#tRQ��V2�Ql�T�d���!	�볊E`ڃZ�m�/f��y6�Vݎ�egFԜ�q�\�cM91YH-p�&zK�䕡 Hu1���wf2��Hh7-6�٘/mu��R��rsJ=���t�^����u|�\���������[h�f��#3}u`{�m%<��6�q_�1{�_>ǚ��7�W�w^�_��q�u����"�����`w^�{�j�~��;�|��� ��la)�d��K:���}�X|�&�X�嶏�r��������~t�4���A�%|��+�u@/2a`{0�}_��o�߇&�	�ruI�tq�n)�=8^�wV)7V�����wrEyʊ�,R���*A�@žP�n^��|�7�W�r��y���^��M�]���j��?>|�?�z�IĄ������|�n{�tjI���f�帽�-$��j�3�N��#nPfo����E����b���٥��w�^�**��廷����(�L,7ܧ���X{@�$Y��D������(�����:�]X�۫?%�v�����%'F���t��\�G6g�m�X����قݴu���Ba�dgB��߯ߧ�35�Xyf��U�KS��]��a%@d�V{���Fo�u��1{��y���yҨҎ&I�J�$w��q�^g�f���!�`!"��@,2�I@CHȶ"x��)�z�T��q��ԛ���ua�K�HJN*�RIV�ŏ�P-w&j�37�V�w}���h"z�r���Hi���U������仾�Հg��*��0]x���%$m�Q��`լY�:ή�m�+H���a��X_}�8'�S��t�������}Vw޺��P{�3W�w�%{�(�dMI*��7n���ꬮUZ��ߛ�>��~�{}�|�R^��O���$*��w�p��v~�9U��~��=��]X�j�䉧F݇��c���,�{�7=뫯Ǵ�t3*A,	#� �c �������(�ߙ���>�/(�	 2B9���]Y�����UU����������c�3�&Ѕ��ڝ�p�΋t�3x<��f��o[��t*�ڮ[{�ӑҨD�ܒU����_����>]�{U��z�`��� �8�R�G%X�9���)��=�`{߿]X��sn��8���"/S�T�8�&��������ug��fo���^ �I\��%JP�;Գ{�37�W� �k�W�{��ڙ�;k�`J� ��7%X�mՇ��k�|�����`g9����pyQs���9�pyT(>hc0��LifbH��l�$�x�1��@�%(I���,"N΂;�%,́�n'�cCF�[Q�{�6:��Ji�����vI.�)֐�Kr�uQ�-��3�*1!E�:�r��qo8��*���l4駷����+��EDU7]i;������P�r����̰Z䁸���.� #!	���v�D��99��ĭ��d�G�6z�UTAUE}e�DEa�1AN`�{{���o�ŵUUҭ]Uu[K�UUUU�W��P*�r�V�mUUUUz�jڶ�^kT�T+y���<V�#(���n��A�/qb�ix*�I�c��2�AOY���ܹ��ڞ�6�ϩ�{��GYac��㒱���w=sMMc ɺwcإ�s�8ɮw2<��<F�<�x�q;��u�S�:���=�ザ��r����Y��4��]�E�l����e:�c��w:��8}mlYTpe--�#@�j�l6I�9}�b��ڶT�P���);�^t�A����E7�7J	31)s7��[����������DJ��73�ڧ����|�	�u�͑rT*N;g�L��ԅ���'.����\6����n=];��e���9l���[��A���a733 \���4��Ɣ�p����i^N:Cx鉤E�]M)7Xi]�J���&:�J�sD`�[��E��H:�����o$6���A��ы�z�jk�:��8kq�n^��t�[��7I֡�^�<twH]��[�D�g\��F����vŞ��^
E� �&9��iv�S��`贾;0%Vm%]/S1��D�u0n�����51���A�Ƅ0Z�[�ln�)�����&_]7<N�;�4h-�[��YS�������ˡwC�H�'A�iЃ�N8I��,�"��oj	x����k����n*���k�ɶM�k���;Q��լ�臮z���ۭZOYͫ��R�\�e�0ff�8re�k���.�;,�e��ثm�j��]�4����c��y�4�z��B��!ڜ˥VÀN���һOKu�tp[��1s�]��lR�`06� �W\Kp6�9�Y���XܡYz�n�Y|Z�)%�-�s���$. �a�mu�����7+;m��]�͇1�W:Fk���\�������5�.q��������c�N�`�5�ֱ�EcZ�k�c��C�:�'�E\�� ?�W��j�D*�?���`k`!��_O2~�ػM)�OP*l4 z�������ߝ�}���`�[��t<�ї�kk����s֎�^h�;��Vlc�c'@��.��q��َL� 3�c�t�[��MX��4�X�i���H�)�j"��Wh�ظ��M��::�]A�w��Je��F���f�=�T��qf�p�x3r�ƫX��9��7f�.^�		@�	�s�feU�2\���I	�A6��m�Y�\���7F̎��\W��rl��u�sZ�@��a�?����T\���kuv�@?���-}���z����*�¹U�y{��Ձ�~^Bu��&�`ے��wu��۫�ͺ���?W+�+�ƍ�h�M�!$���{�Ձ��mՀf�Z�1��]o5ҨD�*9�`��ܮS̭�kSv�w�̓w�s�����{���������:$PmԨ�e�f�|����iu`}�۫ ��?��庌� �b��F!;��ܖ'�۫��̫����ⶑ�{�y�9�9%N!Ɓ7�1o�;I�۫i�m���B�m��뛑�	}������6gg7�uW������Ǹ@����ep!a �� ��9 `�u����:�N��3$�ߞ�]@�͢��! 7%Xyw6�X�\6�UI|����z���BQlJ�6�p�������h:�|�|�}�.�>�Wfߋ���g�Cr�$G`|�����UUn��W�$w6x���P}���Є|ۖb��.296���]�ډOd7^���Q�H��G`ug��&��<�Ԓ{�q�(�>E�2r�ﱭ�:y��R�H�A�I�����s����߼�Y�{�[����9č��OQ"�n��� 7��|�5;?�+�s�*v�������T�?.5�I9Ù������$��8�&�?�ʤu���-�;�����U%��#���EQ��Qv�V����>�UWso�u��k��;^if�*t�"u%1��)��u���+��Ѯ��j�u�C=;-�q�^u���#�>�M,7\1/�r߫�U�[�v�5	�M����,7\���Qʪ�ά�;W����ri��5������n6���1o�;�3]��9\B���`�����$$��~�s����{��͞?|��y�����0C���RYq��l�8J��p&b&�����ȁ�Z��(���7�'��;�̙�iH�M�`}�������َ����>����ߖ�s.��k��u.]4u6\���ʶ;B�2q��-m��;�J�C�y͙�l��@=_�8���ՙ��w&���su*J�Ԓ��H��%՛�����Sg��ߝ�����
�5�H�J+95(�2qJ#��ջ���so���U�RF����k�;�W�h2Q���ri`n�������s��M�>���*��IIF�RU��V�������s�ԓ�y��a��ES���sh�%�X�۬��]]�Ԙ�:l��5��wr�m.���]�P΋�<�v�\���N\O�^Y ۤ���;Z�a�^ l6��JCF��MB\���q���X�u�Q���{��pĴ$�n7M�{vN���'EŪ��6V�c�q�H9v�r�$ \5y��湫��'%������K���ؠd_�G�1���N�t��uËg��S!���5��&�b@�m�],�&�t/,�?�o�O����w���sn�W9ʯܪ�u�������
:%8��Ga�c�-��6�͞,}� ��c�s�W8ٵ�ߩҨE#�Q8��7k��`yo���8�V�vw�]6��ӪW\�,������/n��3�������=�B=d��J�hv��ܮV=����}u`���6��c�**N&��j�˻+�z�XzQ��Q#�6�8�y����v}��u�nmՀf����Ϙn?xV���S�2Q��nm׾��^�QTp G�aD:p(�9'ۛ�d~���i�6������$ � �����/�MJM��J�~���vf���XnmՅ�v)
���GM�a���Wꪧ�~V�y��]�ߋ ����;�uF:%H�)"�1nh�"�r���������5X����T���vr���s6˒;l\p��;c<�fy��d��"xn45�t�'q�׺�7\:�����-�;��4
W���7R��Y�����r���z~�+���,��M|��"�?~�8�̷���v���_~��]����~?8�� �bb0RT�aH��R���(��B	���D�]�ֿ~V����ژ����Q
Ea��RY��`{�Xf�>]�;��֕B j*����5Y�IW8��w>]�v��K-��?!8�Q�(4�y���fź+y���+�����Vb��Vf�Ыl�a#q��o����v��Os� �{�`{_��"TQH���w]�]h͞�`~ݞ�� �y�{��V��R�HI#����,͞,7_��{���Ǿ��86:��,�&�bB�p�&�|U\�Us�B�bD:)�"����]��3�'��)
W�'*4�J�HXn��9\������@7��,�6����F�q�E-��6�d(j��we�09��2�=�7V6��g1��j�I7~I�箼XnzXw6��������(ʚ��qʍ��3��`}�۫�}�O��l������g�ꟚP��dT9%X��u`Q���ݘ{�n�X�/%B�&����9ķ�p�s]�w3���+����Դ��~�u)���q�Y����~�W�{���}���3u�?��ʢ�$��"	��
("H��(%hC�JF	�����\F��Vf�6h��0X䭗a�A�9G��W�<����;\��/-�y1ωǰ�c9��S�����څ^8�ϟ	�'\�(�i@��2v�����(�S��*�1�9� ��Q&6�D����px'uG;��5�$y��5��vݭٻp�����̜u�Hn�EpF�LcR������2;�� 6A�M�->�T�<�+vu�U����Irl<�����=lukgRX�KaY��m&�6��}�}���x{�u��}�|�U��wu�U���FTD��q7�����r�I�����:�<��9č� ���'#Mԩ)��7�p_f;q���c�+su��"u�H	����`ufk�;�۫W)R�y�H�4��z��qȓ��Ż�`}�۫ �� ��0�>����=�ݭ��X�G�ȣ�mdZ]AXJE��Bj蓑z�E�R�hU�a#�����3v�����;����բX��F��J��s����@QQD�@��SDQS����
��$�=D�B��A���gsRI��w:�o�y�����#�����:���lv~�� �f�=��o������8�śL%H�iʰ�zXwv��3u��\���y��Ձ��z�6�� ��R|s޺�?UUV�yX�m������`z�$�=�~b߬ʌn����g/n�=�9��d�]p��2��Y��.ƿ�>PG��79m����
����}ܺ������a���Ձ���~m���$�&��FVo����A��K��_����A�
2j��MN9NIV.��X̚_�r���y����E�s�T\�9��_�6��OtX�J�ڭ¤�Q��Pp�cC���Ei�
��x�
1�R[⑛
�h@�T�bMf�DHR���l��u1�#���t�,ȡ���-�ݘ�5�U0T���@M�km0Lhs��In���ލ!-]j�!Y�(�"��O\I^�Kné 󘯝��t�$Pczz�x<�T�-�Vw��X��ބ�vYG�#�k�lGD-�Z@j�k9�b�e"L[2SK48.1x��B��Ebk�T?���d&W��������:fq����8�:pa�pq�x�v�ۦBgl:gN���n��i�fB�g�x��:qӠ}�� �B��E�HX� \ �`E����֡T<��i]�(���C�*� ��C�)�/�+�@}�� h8 T2��_E"?}��.d��ߴjI�p�5EB*TrKk�����Ǜ��k~A�ߔ��u`w6X��@���tF�rJ�:�T߸Uf�ݮ�f���;��V�������5Af�G\�A4�d���`g�-�����H�Ji�L'%)q(���Հ}��x���{��� žP��a�Y�m��	9[���������7��u`e-�>�۫�������9$�Q27%������b�(ۛu`w=,��u�I�6�1�Vyŏ}J׾{Õ]w���~>�A$��$�E2BIC0�AI$��>��WbD��|jI�s��S9͔�	#I�?��ﮬ����>�۫嚠���c�Q�A�B'C$Ù�Z����Px.���qa5	��,Zf��P献��8�I%v�3}�_�;��1�sn�Ļ�@%�ED
�I`}�۫�1o����^�GVo�}���4~��|"�YDm����~V�ͶY�ĺ���Vn������'A*�(�#�|%���f����q�&���I�@�\�~��^u��m���iʰ:�5�w6��3u�/��u~H_�ݣ�R��ph�+H�Q� ��8jC�e����c�����G��9"�D�N�:�hNg����.C��8Ƹ����[�ˣvtv��<jςq{<�Z: 9bE�c[��Ļ-���lL�\�F�����n��e1sn��_nnms��n8}I��0���7W/p]�
ѝ������U3ۮ�%��h)�vϘt��;�:z;e�MU����ز��%�m��n�$zt�6��`��#sv���&V�[L52�L���F�]�h����`�z�+�vmrߝ���g0"I)�L���7?]Xn���u���U|���K��B���n�7%Xn���u��n�XY��_�W�Sg����[r�t㌧���~V�͖~�9ĳ6x����A���"6N'M�X}��M�r�������y�u��G� �B* TrK��j��c�+��`w=/�U̯�Rm����v*�:�,׶8*����g�N�Y���M!%�Q�p�1o����`w=?s��#����,�k��2"	@R&�tg~{�~>KܕU�`�Ah��$�Fmb�h��M$f��#N�jKA94SU�4����}�{�]��=��(��P�]�u��Q�����$w7�Υ���w�M��(-����:��H�*�*���,?������`b�(���仛�X|���׸�%&�Jm��žP�UϞ激;��X~[�~,~|������𸮹vam͉�K�v��j^s���1�d4�ی�>P��b{1Q��W�Η����7}��4P�4��I�(��bq��������`uf����?�UT����"rQS�ɾy��\���u��~S���A�EJ �S���~^{�grC����m�H(ۍȋ�A���ۮ _���;�M,<����PB�9$����\�*����3?z��;���X�
_W����k��;Hlz��l�*�Rn�FZ�SciB��*2�ݚ��ۖ{�u`�{V��W���u�U)H�%Q27%���]w�4|�漴�3��UH��~���һ٥�O��=��p�~�X�����m�F(�NF��$����6X�=ua���:���`�f�&)�-Y9d`E8kA�b	��0K#J�a2L��!�Y3",�l�#�p�)��ǣ!8^�0c�c�Y�Q����R��g�x�D�C������欛�}���7[�8���o�@��w�W�$�ps\�t�z�r�����ժ�ɫ.{M�n6�[���	qF�L�R�B�HL����1v������ gq��s�sK��/�B,$J4�rU�H������M�������\ʐ=�~��!>4% ?{��� ���uz�~��-.��J[N�*2M�s},�[�� ��8^��~�8uѸR��"U#rZH�����o�(�p��R��p�T`l��F~}���s0ۜg7`؋�n�I��ԡ-*2\�+��]��F0er%Bb�A�+�豷S�9��Yۑ	�<W��c������M�e�P]�mU��K�#��gduj�pIO6`.l[e}�pgz����FQ�,qm�ؐ��Ő^�n��p��:Ѫ���v�vnH�k�-���Хy��6H%�0X�ƥm��r�`$��4�4�5�n��n���WX��;]Y��� ��WX����X���{J��\����m�6�9%`��� fu����f���!w5Q~qT�88܉G��� _��m#3�u`f�����\l� ��")�2; ���~H�������~pw��∫!L��|�Ia��9_�������`���@n�fzX��RI�8�i�$���Ǯ g����,��׾A���JO-<����k��<�]��O5^{CY����@H��kc~�*Ӗ��N$���5/lp�ܖw�u`��]a�N�Dd�q��g��s��>�D=C�z/���;߿]Y�F{����*R�$T�&F�;�� ���W+��r�3k�p��,ifb=WM�m��SrU��r�M�8��}��`w3�Ձ�q\U 8(܂��3u�?UW?UWw}:׽���35�?r���s�YJ��p���&mW�K3-������=(��v���V��8P��*��?�;��x�׻u`�{h�[ ��A25�C��G`fn�_��) �W���P���T��բIU��F�rJ���J�����"�7I	���*I�|N�:t�2�DqMHa��$�l#0�I�K<]�D=��@p����5����R���Ձ�[��jD��R7a����]@?cž����� �k�]u�d��&G���ۍ�w�]6�$>���5����ݕ�H>���Ң��JJI�s��I�s�t8W�'�㳖@�<d�s���F���%Q�G���]Xw\�G�l��9h:�?�A����I���JrJ�{�g��q��{�?[9y;˩'=��<��*���U!�7"Q�������k������ �y�H��mЇ�	Q�G`b��=��}_ g��s�+����C�d ���L���L�:H'⚞�_�׵�*~�2:"H����]X{����ײfֿ���b~J�"%=��gˑ�z�'��S[Y�l��/`[ru���hxS).@�(ӎIV����c�|�^�W�%����U��A�(M)����� ����w=�����H����M:Q��X�|���ug߹������wg��?%DG$�Tm��z�K����`o�����u����Ϫ����������I��$t�%{�%�ǈ�z@>_w����۫<��nU�ng�rns���ns���??J��e��}�@�T�B��9��{�@(Z,�4�W}\0˫5�@QNn�kd� [#�"(Ɏ�*��l{7�e�Twz���jq��N�µ�8u�fI����ED��&�3Ɲy'}�F'ey3΂�Li�s�Ӽc�h�d�oN��[��#	t:î���C�`���tu��Q�)�)�!���0}2�ǼDZ:b	:��n,Gp[�� �vp:����Ť9���d��7i_���� �'GDbT��CjX�a��~ 09�IJ����[L^�Ei��S46���ܙ)(��(΍h�ã��(�r<�I�X���u��g�5��PZked���1��M1�,<�h�i���iM���'���븉3\�ף4l�1�m���6��ɪJ��MH��G�8�wH̴g�4M��&&��)�c5�nh�m��j���U�Tcq,M�����ڞ��f0�-�E&DDfRt�8"�q��>y�m��`��uUV���J�U�][UUR�T9wj��j� �����ڨj�e^�T��u��HH��a�q���*5�KlIhmL�Vg6�:�����0Ia���Yd.RGnf�s�n����(1f��:<��㪬0� �D]�`.�T�0j=��1�②4F��[�E[+Jv{n��:x�loi�x0�ݺI�q�@2���'�Ǘ�[��wn��[�v���c3v��n�yݘ�[gm�s�.t3Ӻ�Nwk��Pz�r�/;�\�����"���s�9y������y�8̊jX�^��S����U]���.�C�:��9����z+$[��=���kW򜛮�Uǅ��JݰOg���3�[N+��.�E�Ƕ��Y�wK�!r�L/;n��rjWi�wA�v5�l5�YM��������j��Jjۓc�=��epnFl�aldc3�ҧFqu����^�J52�4F;�����P��s+<���J{3L+��JlS�u�yϑ,�n]���]��iWCJ�1�]�L��s��s�L�m ;h��ۦ�<�۷Zs�p2��5�����Z�F��ݼ8M��1!;ź�flA�!{b�1{x紹�]s�u��y��`4�ݣ��R�B�#f��,
�:/&m���q�]�H%�3���s�t�:��[h	�W.��Au�@.֐T���M5S$hѷ0��K��:��F�'ނ�`'Rܗ*ѳ��Xvݮv��f<�V �h&�[��qLh��6v��R��\�SL`j���]��.��Gj��0�k��g�a�pa�&)Lږ���Qsl���	5ɁbѲl\�xX]Q�U��]n�U���.�Ϊ[�`§k35����Jd�6��H�U]��vt�x�\�r�M���.�q3�r�b�J����Q4����B�Q�1���	s5�������N����
_U�;T�lu�<�"��#�'�j	F�Ĉ+WhQ8 1���p ��ԗ�/!K���̗+��ba{�%���ɔ�����v��6^7!��3���ԉ�E�Ot��Ǘg0�4f-�
���&6�7�p=���v#��B���V�;�3��s�2qpk�ғL�,�4#���(�t6��.��=��T��v#H��@��v�N�c�ܻn��Zy�D�����u�bn��^��gA DM�1F�V�ʒX&.bQ�+k�̦:y��'�ŜT潴�:<Ռ�2m�l��3���EQ�T���^�䄾�?|���]?�]�����Eo��j�N�q����~v��۫�Fy��}�4��2���L���;>K���X�������w�?��Ԅ�ĠF�qI�?%�~ k��ݞ,6��s��X�ՏВQ)�9#e�/�� �ʮs���������Ձ�z@?Ur���)�g��eSg�yyK5ŶZ�/�;��e�A��U�v���J���&�(��0�����>��Ձ�z~�s��A�= ,3�r$�3$2Y���o|��5�>ItB04��@+��ׯ|���$s|ν6�t�U�Jq�H��*���_���w�<X�}�V�����iI����_d����Ɨ�ݺ�1wT��9]�+5��N��������UU�����վS�D��j��?��k��,�6��m�=�����Jd��CPprKK5�]+��*�9C!`}]��X�TV����+��fO�����|�qʒ�=��A��P��u`}�۫�IW]{Ǔ��J4�7`uo�@>�2���
�9B��0�|pSHK�Rd��#�G�!�]o��rs�}a�N�D�M���\�,�{�;��Հ}��z�q�o��O�܂U#J�jG*��������y�uH�!7�y2��bX�'�w��&�X�%�?g�|�~3,#.���k��BX{$#v����u�u�>
ެB���}�=󟼕��f����*b%�b^��j�bX�s=�MD�,K�9͙�|��&bX�'���SΞ���:'OߟϮ{[���_�2L�$���m9� �I�2N{���n%�bX���i7ı,I�~��4,Eh��g�����L3�g�Mı,K��vi7ı,O=�4��c��1�ϱ��Kč�}f#M�4F���6j�����\�94��bX�'����I��%�b^��e5ı,M��L��X���EZ1A�]���+�L�ϵΚF�#Dh�_y��E�v��K�1���Kı/}�2��bX�&��&SQ,K����f�q,K��9��Ξ��9:'Ow�ğ�Y�4�e�c��F�ML01f�5�#B��GkuU�;����&�F�#Db��>x�4F����sf�q,K�<����;�Z#Db����Dh��}���Q���^����#G{��4��F�����vi7İlK�{���X�%��gٔ�O������b{�˫�Ǚd�-̸f����#}�_��q,K�=���n%���7����̦�X�%��}͚Mı,K���h�f;���q�h��4N|}���X�%��sɔ�Kı<�4��bX�0\D��o��Kı�:I>�WϮf�u]�ˮ󧣥:''���.SQ,K���Ȗ%�bs�k��Kı/��2��bS�t{�}��w��ό�� $�K�ֺȵ���u�����_.ݼ��]web�Wu'�1c��<u�Ai��0
#�\�0���.�ONA��u��b�r�zؼS$�'��6}�siJHu�(v�j�k
/gcTKql����Kg(F���y��jK�����LBt�ڬ]r����@1v��>okmLݛF��l� 5�[��S��#����w��������V�t�Ơjzs�q��wi��z�s�#�o!���q۩�C<]t3o�v%�bX����٤�Kı=�5٤�Kı/��2��ؖ%��gٔ�Dh���>m����0u��0�7ı,O{�vi7Q#���b_{�e5ı,O;�L��ؖ%����#m�$X��>������f<�\�f�q,Kľ��2��`ؖ&��fSQ,Vı<��l�n%�bX����y�ގ��:'O�>|_��5]��n%�bX��g�)��%�by�9�I��%�b{�k�I��%�%󽻧�D���x?}�J��%��7ı,O}�vi7ı,O{�vih�h��}qh�X�F��y�âtN���I��<�j�31�.GG	\W%�k�_o9�s�:�-�׬"�'f�,�K�ۦ\�\ˆ�ƈ�#G�}��H�DibX=Ƿ��j%�bX��}��@7,K�u͚Mı,K���:M��ɆL�nK�B�Dh�h������ ��O�T�Ĳq�����b/��z|��2M�ɔ�Kı=�9�I��%�bzw��y���:'D��ߵ�㙭Е�l��7ı,;�L��X�%����&�X���LD����I���bN��qh��4{Ϳk�����8��n�bX���vi7ı,N�<��Mı/jb&s�e5��,O�a9Vr��G)��|^���0Sɤ�K������5٤�Kİ���)��%�bo��2��bX�'���4��F��8}�|BR�<W#�K����Me,�	��1�+�-&n���yܿ�:y|�$�ɔ�v[fd�8�#Dh����Kı=��e5ı,O<�6i7İlN�<��n%�bX�`�gn&c0�&2�#m"+Eh����,K�ߜ��&�X�%��g��Mč�4N}��i�4F�Ѿ�{�W[�&#��m�4F���ih�&I�����u&L�4@]B`_���d��"6�R C�<�'���4�9b+G�φ���:'D�����r`�ʰv�M&�X� X�����7ı,K�{���R%�bo��e5��,O<�6ih��4t^>�E�^fL�2�I��%�b_;�e5ı,:}5ɔ�Kı=��l�n%�bX���oH�Dh��V���X���ji�Y3-�f+5�e���K�,�n�%bi�5V;[M@�uK��'\\xf)\��l:�����t���L��X�%���l�n%�bX����C�1ı/y�e<�LD�,N��[Mə�)�2��6�#Dh�~�f����!)<�߶���/��[B�6�w���K�*�<t�3_e�d�LIs���n%�bX�����n%�bX���MD�,Kx�)��%�Z;Ͻ�H�Dh���{��o2�vY��:Mı,�"b&>���j%�bX�c��MD�,K�>��&�X��QH��/��LaNu&��8�F���߾��^c0�&�1��ı/��2��bX�%��Γq,K����f�q,KĽ����4F���y���7i���̄�з.e�U\��̄#���"N=a�,�7W���}�V�G��%�H�Dh��{�}�F�,K����f�q,KĽ��2�
%Ԛ�$�3���Ӓd�'5�����$�sm%�q��&�X�%��{��&�X�%�{�q��Kı.�=�SQ,K�����I�6%�bzp��%�6��l�y���:$�����wO,K��=��5ı,O|�ys��LD�,N���n%�bX�{9�{3L��kə�e�6�#�5���LF�X�%��g��Mı,K�s]�Mı,@!���;���X�%�΅y_�	(���p�W�)�r�\ܞ��K��;�k�I��%�b^���Iԙ&I�w�����$�2�4?���{C1�@��l�ָ�vQ�53�5ƸP�w�����n�9�yь=�3���n��Z�u8��Dދ6�ׇl{]hS�ĝ�h���20�À���]�k�.��\��c�y��wFZ��
�.�4�7v�cm�\B;
�!˶%I^�?�v��m�B��m�ՖeG�n^\4���fd��A���BǍZ��.Qؑ�H�`�R4i�\`�CtzS���#3���K�ۧ��]&��!ü�B�ф��ƭJn:~��������Kı)�{���X�%��gِ�P��������I���:'O�����mu+[�<���j��b_�MD�,K|ϳ)��%�by�{ˤ�Kı=�5٤�O�"�F��ߤ�)�0�&̷H�DibX���̦�X�%���.�q,z��LD����I��%�b_~�MDN��:z��߸�Aɥ�m<���Y�D�5��&�X�%��y��&�X�%�|�q��Kı9�/���"4F���g[�5��2H9r�M#m%�b{�f�4��bX��>��c)��%�b_}�2��bX�'�g�]&�#Db�=�[�d��d�ap��ڱMk��x��W��<Gdu�����*�����.˗%Ǥm�1F��>���#mq�/��2��bX�&���.�q,K��ߋ�|W�G)�a�~D�N���33H�Dh��s�\F�@K�%�(�E"-LZ
"��kđ=�by�w�i7ı,O=�4��bX�%��SQ>D�Lv�"/�~��@�p�;�|r��G)�l���n%�bX�����n%��0�LD��q��Kı/��2��bX�'xߙ�<`��u���ж�#��Hi����y���Kı/��MD�,K��)��%�b{�~��n%�ct�����9��[�<�������qh��4M�����,M����7ı,O{�vi7ı���t��>�t-n�-�5W9Ǐ�	��λ�Bu��cU��J��������6h����G#Dh�����4F��7��I�6%�b{�5٤�Kı/;��i�4F��������2<.I-Ɠq,����i��Kı<��]�Mı,K���#��%�b]�ۺxNN��:z�����)��������bX�'�9��'�Q�Kļ�q��KT?O����ֵ��kZ�����80Ffv�~���,�&��#��$Q���X� �:Q��	ѐ`ø�㉔��XHq[�W��ӱ�n9dfe&�����f,W�1�!�:&j��F��J�1���,M4��;�����9���xh���`����4��&#���,3�:�zg�UG��������EĘ�H�G�y�;�Ȱ��(�������"(�J��"5��;�cW&#�0�r���q��	�	�E�l��^� ���Y
3����o� �������C 2kCM�Nw���p�����&/il�U���'{,5�Ӈ4�%�z7t͍ �'"31�������[������5���NH�4�ip��t�Xb�R��&L�7�g��O�OO@<�Q{�<C�ڇ����[�S"F���)� (x����ԑ�!�N�S�t*x����b�jNI{��e5ı,Nc��Mı,K�>ղ�f[��S%Ǥm�4F��9��2��bX�%�=�GQ,K��<�1��K�,O{�vi7ı,Nu���o)��s1̺F�#Dh����i7ı,O1��Mı,K�w��I��%�b^{ٌ��X�'qS�������)tnm]WH��,i�)��ga����.;i���4K��󧣢qbX��yۤ�K��O{�vi7ı,K�{�����JD�;�yr����4z���d�����yeɤm�ı,N}�vi7����b^��e5ı,N��\��X�%��s�1�&�4$�Eh�]���6�=�2̲����6�#D�Eﾸ��F��7y��j%�bX��=��n%�bX��5��6�#Dh�~�O�3<��n[�n%�g�1��)��%�by���I��%�bs�k�I��%��h����2�u��LD�#F��G �(��R���]�MD���:~��=���L�L6��ގ�щby���I��%��S�X�����yı,K�>�SQ,K��<��u:'D�������3n3-x4�H�oeq�� ��Gg�8���������ir�M#mb+Dh����H�Dh���;���X�%��y��j%�bX��{U�9H�#��V�z�5�H�RJ�7�Mı,K���)�|*��H�&`؟c��MD�,K�s��I��%�bs�k�I��"����Lt��2�5��.�t�tN��:}��;��%�bos��n%�E������i7ı,O�ϱ���X�%�Ð5^���E|��R9H�#�ן��7ı,Nt�4��bX�%��S�d�&I��ͧ$�2L��������]y�.����#G���zF�X6%��q�~�Sq,K��=��j%�bX��>�t��bX6&@ί�	K+�I�LM�����q�1��~�َRܹ��FX-`^[u�V����Bs$�ד�����/l�ݜ��A�yyC�m����\a����z;X�烯���qn�"{S�̇��d�\�n���X�ل��h�NX\�7E�'�����H\H�] �չ�����B�;71�乸���=�Zh�+e���-�灅c5���e�-%
a�Ս\�Q�fy$�R)��ݗcw1�0�s�5ʽU�v�y^tJO/���-��69�CËUS3��k��>��tN������4F��=y�1h��4o�ޗI���bs��f�q,Kľ�}'Ҙcǒ�.e�F�#Dh�^�b4� ���4s���#m�V���w���n%�bX��wMD�K���o�2���1�l�6�#Dh�y���7ı,Nw���n%�bX���2��bX�'1�)�6%�bo}��L#��.[�H�Dh���D����I�6%�b^��e5ı+G��x�4MDV�Ѿ�O�H�Dh�	������:�;i�n<���r%�;���X�%������n%�bX�s<��I���bX<���&�X��������ߓ$��2`�Mʊvn*G\��*�\=��u��v9��u&���]#lQ�4F���x�4F��7{�]&�X�%���]����Lı,K�����X�%���O��-���#f\zF� �#G/���c��1����v��6&��ni7ɒd��ki�2L�$���m9&I#GO��'�o&W^F�ˤm�4F�';�vi7ı,K�{���X��+Eh����Dh�Q��߾�F�2Δ�?~�UOP�r�Mq�OGD�τ��w�e5�,K��)��%�bo}�i7ı,Oy�w���Dh��q��Jare��n����ı;�yr��bX�&�缘�n%�`؜�y{4��bX�%��SQ,�����Ş�kT�ݵ�Wn�5�n:8��:��3=����5l�Pڠ���7ı,O=�{t��bX�';�vi7ı,K�;���|-�&bX��������#Go���9��� �3���7ı,Ns���n(�A�K����&�X�%�{�f2��bX�&�ϼ�M�� �"X���X��&W�30���H�Db��w�����MI�3���Ӓd�����!�&��	12�e�f�����d��T��L� �i�(��
�,�����N�:�Mı,KϹ��&�X��4x���Gwc�d��e�6�#��������#G/~��h�lK�}ݚMı,K���)��"4F�u�ɯs28��ˤm�4H�'���Ɠq3���b���f�q,H�'}��i��4N���DV�tN�d����n-��i�ZMW���m`��i��n�
F[�J�T����N������.�#yr�\h��4w�߶f����,K�;���X�%�y��j%�b]Ao9���ƈ�#G=��Iǒ��Km&a�m�4F��9�#L�$V&"X���D�,K�{�q��Kı<��٤�O�P�LD�/���٩6��v�Ξ���:'G翷N�Kı7�9�i7ı,O9�vi7#Dh������#G}���[dy�2��-�6�#�M���߮�q,K���}�I���b^{�e5� qCj�tgR���Kݝ��7�٤ē@2�A��Z%��#M�4F��:�n�ܬ�9�4��bX�'�;ݚMı,K���)���b_|�2��bX�u��f����#G�����e��n�P�)����M�T��5�a^G.T��Hu�X��Aź<6B��f;���ˆ�ֈ�#E�~�SQ,Kľ��e5ı,M���M��,K�yݚMı,K�o῔�wYnc�t��F��'~��5��,M��sM�,K���wf�q,Kļ���j%�bX��',׌�^A��ۗH�Dh����}t���2L$��~��uO�F�ԗ�����X�%�}�q��Kı<?t����,¼��ˤm�4F����}�I��%�b_9�e5ı,K��1��K����ǿv�I��"tI�>}����le�mt󧣢tN.�c�{���X�%�ʌq��MİlK���Γq,K���}�I��%"X�8�Q�
O"�0���"�F�Q���11i�q�a{f��.�$�H@�]- (A{Ok��@n,��Q'7�6;6�ϴ���ܕ̲��V�/Vb�q�ŢF,k4���b�;�in�ƍƔhu����]��]�wy��s�B5&�
3Vl�ʶ����7A]a]�ܷu�l����3๷kvnG:��ˣFfY�N�;]ۍ���]�f���m��[�zN��˭���fƇ�fc���D�Y�A��n�(Q��$��f64�S6;����[����:1,K��1��Kı.���t��bX6'���f��'�1İo�wMD��4t�7��[&<�t�ˤm�4X�%�߻�&���G1��{��&�X�%�}���j%�bX��sM4F��?s<��U��8�ff��+ı=��٤�Kı/���SQ,Kľs��j%�bX�}��t��#h珴R�e����F�#Kľs��j%�bw1�v�)��%�b_=���n%�bX�����n����?��%�Ǖ�˙&H�Dh�,K�{���X�%�w�9�&�X6%����&�X�%�|�q��KΉ��O�~�}���8"l�v�Gjn���WM)$�n.�xd�M�-ֹ��g7.���4F��9߾ˤm��F���yݚMı,Mb�=���j�bX����i�1F���=%��
�W3��I��%�LD�;��I�D(|>����B�uq,Nw�e5İQ��ۈ�Dh������6���X��=��?Ka���;s2�m�4H�'>�k)��%�b_9�e5ı,Oq�cI���b{�;�I��%�N�ϟ)�l�FWy���:'D�;������Go;�m�4F���yݚMı,�b'��yMD�,H���o����a��n����#G1�>Ɠq,K���wf�q,K��:k)��%�b_9�e5ı,�N���x��Y�k�l�*��FԺib��.DIR%�e�wB�'�k�쮍���n�f���%�bX��~٤�Kı;��)�2�$�<�5���%'����LCb9�죿�c��B��B�s�a3�,K��c)��%�b{�=�4��bX�'��4��bX�'�~��v�+yn7sH�Dh��w�;��&I�y���\N���@��9
@J�y���U<��3ݚMı,K��SQ,K���[�;���ˤm�4F����;�&�����b{�wf�q,KĽ�q��K�����{�duı,O���+>$kM(&�����:'G<{�>��yı,>X��}���ؖ%�}�q��Kı=Ǟϱ��K�N���_���-a��g�u��Y�ٶggGs�Ò�7�`}=�+ӭZ����bX�%�{���X�%�|�1��Kı=Ǟ�Mı,K�yݚMı�4Cޏ�ψ���n����X���MA�,K�y�1��Kı=��٤�Kı/y�e5�h�^����rc����h�%��s�cI��%�b{�;�I�1��/y�e5ı,K�{���X�"4w��~����1�r�ih��D��wn�q,Kľ��j�bX��sMD�l(?�!��x(�S^D�ߙ�n%�|������W���mn�Ξ���:'G���e5ı,K�9���X�%�w�y�&�����b{�wf�q,Kħ}��h�+�,�Ųr�x������bkI�p���B�P"]R�G��r�v]|���,K�N�)��%�b]��gI��%�uS�xw�A�Obb%�b^s�e4�#Dh�[ϥ���\��.���%�b_=���n%�bX�����n%�bX��wMD�,K��c)���4F�����),w٘ff���ı=��٤�Kı/��2��bX�%��SQ,KĻ���I��"4F�����w)��s2�m�4H�%���SQ,Kľs��j%�bX�~{��7ı,O}���&�X�tN���=��\�L�|����%�;���X�%�w�3��Kı=��ۤ�Kı/��2��bX�'����Zֵ�5�kZZ�=>�[u��?��ˡ��1�㵯T�6=,�5t��5�p�xa)%$�go�*�qM�9FJd�(�j�����4A��އ&����7.�U"��oF�pl��ٳ{A�FM:��G��Hkh����ì�9M_�@�g��c���&�l8m)@L��X�!����t�H�:�y����a����N�DL�Ə0�a����l��؋�3��C���P&�r=H4B���6(Ҽ^�rM<Wj!�c��l�?.�1cY�h���De�0̻�^�l��J��]3k�����^R1����@�`نe�n#�t�cI1����zl�<%���&`fpȃS��1�9<|�x�8������v�4��c�F���0Ҋ$Ph�͖�ok�d3t�6ec�&�i��3��j�@D��㥓cZ+�u�YǹeV��,�*�#!�b�c��f0�-�xc�ջ���YiaFl�G�>��Պ	���a7�ݫ9
�GQ֎��p���5Rk�A�1)T��X�p�cAU'��:��sllU�)�s�z7���UUr�UU]/2�UUQ�յWUPP�R�mP �UUUP�PN���h9��e��S"6\�[Sxr0�T	;�2�;s��2oW-ۄ��ӌl;R��Ɨ�^�Z�s称9����v��oH�uh�s���k��n{x��-\)�.�[;G$q�N��\ev1�JbՍ
���� Җ�6s*x2c�l򐱌n9���E���\��\!�Z;u�.uE��e��jڭث�;��q��]��!�M54�6�HM����e�lZOA�O���n܄!vɅ��\��H��9H[�"p������..�ԭ�>}ï��[pO7nK���:��C�<#ZJ<^��lmu���;v�e��0����lR81AYZ!	�Eu-��.���l��n�0�R�-�k���@�m�a�|��Y�z��8w`5���,�u2[)iE�ZJYUB:��	\�ɚB\��j�i�1���&�ʜ�tV�mW���Q`�Q���6DBWk
���%�����׍�l�Բ�hzL%��2WO�����yN�s&�nM6t�G7.�{�m�kj8���b����<��k��&l��F�]��7d�NnQ���EۂkԺ�p����6���h�O2w6�y�8=�P]O3�,�,X�
݋p\$�T5!j�B���1�]�� -D�+��v3h���&{��M�x^�鲷gv��S�8�I���Ȝ����ŌvX�����������ή��]m��7��A Gf��bͶ.��ά%��/��u�z��5xv8杲c2q:^A�.s��:��k�:N˵y���]��z3�C�2d�}9���[L�������ru��<nܻ��],��۴�ڝ���Tw�n��Ï$�9�5ۤ�{<s�U���j�D�c��r�c��^m���G\�HU�oR���c�n\�ka�8$�IHI�|(�F
�O.�
| �B���L���a�6�P4��"��*�v
`����`�#�
�6/��u���W��\ɓ����e0���ʹ<S�eh 뵱2��Ӄe�ۮ�<$�үPOl�χj8SӹNZ�:"��I�ػf�ݯ1��9[�~�
�/ez+f�[<������	���ѵ�W��ms�%%��\�D���H͡Ƹ��Ʊ�5l.y�|A�U�b�ۖ;�`���Ê�ᚨZ:�<<J�eP�: ��u���[|v�\yln�f�c��%���X͹B��NL.��6�)֊꽍�Kf;)��o�~h�������H�D�bX�����n%�bX��wMD��4N{����#G~�~Q�o3!!r�i�Eh����ih�%�}�q��Kı/��2��bX��7���F�?����������m�s0���ih��4O|~��4F�؊�}�\F�#_ eh����ih�,K���Mı,K���fe�͙k��d�t��F��'���i�5H�%�we���]Xٮ���T*JHr���������^�� ����rXR=�M�J����qJQn��N�p��B���gD�;�k��[����AR9,�6���w5��r�/��`nbU�1]B&6�r��s��8���?*B�ȝ�Y�5��{�e��g���\�$�K�����9QF�w�����g���׶�9�+v$ȇN("; �fʰ'ٛ�|��ꪪK3\G�0�$�qRT���3�V�� ;�p���*����z���w�ڪzV�� ��gBX�Sd����Wr�"ܭ��R���_� w����=UU��V�X�������35�r���}��`}�� �k��s�H��W9���B�n?�3}�XfmՓ��W�T�)�b]D"��o���ݸ���6���i�aRI,�=uaA�� ;�p���s�i�u��qʰ潴�R����>��Ձ��z	�*W��Q��1��j\�\$�MiD�ت�i�[��N�i�"�9QF�3\��fK�ͺ��y�+0�5��8�����q#������ w���v0�&��$��%��f�Xs\ �q���,��Zc�jII�%}�=U�%�� 7|��ݖs�9T*P��0�.8.�
lAx�����k4�N5#r%�5� ���`ff�XPw5Ƒ}2�K#*:B[�4O3خ%��NA�n��Ϯ�¸7L�nBtD�R���;��`ff�Xs\b�}[����r�T�K36��ă7��u@�����R��u�Lqʰ�Vb��Iw=,��Ӵ�o%$�Ev�庠��d�;��V�� �c
�"��E:q��}��`w3n�䃹��u@>Ha��B�@wY}T�s���F�)kr`��ihk�bŰ�nDn�GQ�b3Nt7&wq*����c�[C']�N���DmYl��֥�t`�fƀ�ѹ�1�F��f5��Qw=>Pn�WV;z����0O��G\��y02�c�C8��ð��Y�m�n��X�q�n�]�����&��M�hR�jіٳ���1&�5���B��sܒ;�D��MZ�)����d����ܼ�pj_aQ�q���]��	�Gp�=����m�BrX{߮�3\,p�ݖbXص�l��RmIV��~�r��p�b��;���9UI�W=�:�IH���Q��� _{���g�����2��tD�QE�}��`w3n�����\��u�;^�M�m9L*I%���]Xs[��8�{����[C�&��&Rj4㓰��Fȕ��ʻS��`��9��m��3�ӭ*��� �k��p�����u`:�F�<��-�m�޹A �K�+�P;�r��3n�0� �3��"j!ԑH������ug��H�o��#}� �VF�M$BrX���� Y� }�N _��`wZ�6BI)6�� �� �s��S�y��ݖk3�VԻ[I��m��D��ġ��*[�5�t��ι��u��nwSȝ��1\�r%�f��rX�۩�UU|���8��W�F*Q"�?�;����f�X�H�� �oh���H*HI`w3K���s�ʪ�ª��19 �����lG�U�����(~̎�{��el���&�#��;ܚXn��ٗ,��Us��o�� ���W��r�(� �� /�rX�۫�F�� ���UJ��I6��<���lu��p�N��:�Vr��t����Q�"��ٛ,��Ձ�==��9h�p�da�aRD!�%����_�U\H�~ n8}論��/	��R�qʰ3��� /��`w7n�Ė������Dt��*��K}� w��XǞU�Ȝ��T*� �E�Ғ�����T���|!΁G�������j����R��(����`w3n�Ǥ �c�o������l�����N��+�+rY)�J��kH���j�%�˦ڊD�4�!6�|�����zH�fc�}ݖ�Ek�8�m6G*��z@�� _{�����W�s���םp�JR2�3|�|�ݙ,����3���J��48E)H�v�f����XǤr���]�p�da��|�(��������Hw ���ƖT�]�d�1<03�!��eXfK�Ӭ�޼�`����^��/b&��5�ǭ�h�Y���2箭���jK�])��YV3ɲq��Nyd�ex��=�ӗ`��F�6�[�:%/9W�M��0`e����ې�֒Ʈ��&��T�[p9�I�ΛY��v.��[���K��|�v�M4t����s�볚U��4�e{5z��y���s�pT\j�\�l�<2F�&H�V��*#��I��?漕�-4+���KY��x{1d�ٞ�u������|�C�E�SaJ�ͷ��� ��(�論�so�kK+iIN4GN��w5���,�s]��z@3�fV(��)JD�v�se���k�;�H��P�LE"�hjR
�J�˹����� }�p:�ݛ,�"��M62G`w��K���>���>]�;��
�OTj9
}<��J���5!�w&ސ�J#�	-��4\�$���*8π3S �}�`|������G6�D8E��`fl��S3ډ��`T�y�^�{潷Q}�=U�RGs�=K�E*'%�՞�3�����e��h��NR��4�G`f= �/��@}�쿒�9\�o=�z��U��	)GN��}���{���w]��z@>Gk�3�:.u�q\��{ٜ�α��tk���+7)4J�JiJR*q� �����wu�Ǥ ��}�1����H*9%����;�H�����,n��k�8�m6ӎ��= �/����� �9�ps���7,��EQ�IA�"��|y�Z6<#|�4�<��M1͛�oXc�p��-%(8͐FC��bƎ%0� �"�XG#,�:A��,��M��ġ!Np��fc���Zے��ӂ�u�����HH�u,跙�;�	$�s�0#����"e:MSt��A$��P�h7��b.��K�i鮓\뤉
�v�f��Q�L'6�l)	�bx��f䉦�fny�0fP���ݯ
�)gg]�/d,3�$2fgol	o[�q��b�d��!�:�8�k������o�ad�5��.I���� m� Kh�]k.t�B4����k�R]r�D�VdD�A�Nftj-ip�=�(m����4�ID��jf�j�#U���i��l2�`��(Rʔ�g��r��f�Y�GY�
��L����h�'�<g�-4�Fk�<�")H�#9�P$WzF��Fi��)�h���]oX�a1�W-�A���c,$&�����AyC@���`�L��t�����h7�P�Re�q�n\�/��x(�A�rx�^�eNC��?�<҉�6����6H/���KT ��� D�	��*d<;DEg�IH�~��i䜜���#���OB����5a���w���jn�}��V�qw'�n�%[R�j(�))�N��w����`�p���2.�~�<Ԛ��Z��M��`L�w;���ƻ�US��1�)�$K�E�H��w]�A׮ _q����A����y��u(q�4�v�k��}��-}���s]���H�k�H�%% ���8����w<��� ρ�YQ�CR�������?��yZ�>If��+���JM�tCAJu�V,&
�M5SV�!��-T HA�@s��6��3�E�JBGH �vz��`�l��%����v����KԼ�)�Q�*t3��� �ֵ�Ny�t K'�7�au�83�x�Ή4�/����`ugT���~����3�XƫU*����*6݁պ��\�8���,ǾV�k�H���ZJDME��VV{���^j����P�%���)U8E�H�=U�,ɾV��|����`}��KX۔8੧�gu�>Y�k���'�c�]I9�:Z!�x��p�/��O����x&4��l�׀%�+eyKq;2b:Z���\k�.�I��� Lj��kpY:ث�ˈ�j�ڹ#L�1���I4�7-{@��zٱZ��@kXw�ň�:vx����^yg^]�+����ٻ`s�����^m��UV�8��)Źۋ�q��.����it�vٰͣ����� |���)�-������7�;2[�敶(^]0�Վ:��:��6{l��mܰT�p8��6�������{�ǹ���^/����8t)�m%"mJrG�>Y�vz�U�w�����S�\�H�i���REDn;[['��}��=���T�=���bU�wGNH���|��w�޼�`|�*�T��9Q6��� ���m#�y��35�>�0�����Z�ׇ��4Og�A��z3��Ǭm���Eug�pD�QN&��>Y���^j�
��|��MQ�*S��Ĥv{�N@�@T/�`A�A,c`f6*�C�̌|�|����Q y)��\�����z��n�E�:Ki�(q�Sn�u�>Ǆ�w��Y4�k���#C�Pr%Q�{��R����7]���ŀgu�>�)� �r��Ƭ�n�3&��� �f(���g�i��P�B����p"F�p�e7h{[S8nn��v�8�i�pN�NS��k��>wg� ��b�P��,�J�n�	"mԎU�gu�1eb���`ff�X-�J�����-�m��ޚm�s޺|AA��|�z�8���}}Õ[�p΢V$�Q�M5`f�33UՁ��p_b�}�0�	 �L�I`ff�X����UnҀ����~��ߦ������2v彐����n�x��ٲ�NN�k\�v���M���r��l��,[��1@�r}�ɶ�ЛJ�M'�㍫V�@�2X�SKV�(�;��cR���mXf�32i`�pY��u-ƣQ��`fd��7u��y����q$��J"������h�cwR)"mʒ��׺�3=,̞,W+�����	Ɯ��q��ѹ�zy�I�l�bx�)2�U�lLZIl��Ll�u T�~J w��`fd���|����n"V��Iȣ����ǞVbY�j��pI�s��UU$g��3D�E�qX[�w��p�$fk�wyX.ם%�۔8��m�`��{��_uX,�vt+v�DTn$��Q� �k�}��V˹��3tn �r�p����UE�Ѥ0� ��4���_z�p�bu�ve�����P#�Xk�9��ꄓu/:��g&�:����^b�wV�tv�]��P�[6^�'et\s�y�3�����v�h�:v��`��᳍��=P�X�;l��-��|�a��Xu�J�C����*^(��qb4��m�e�F��J|�����[z���ː�XeM���#0MT�c�o�sm_�@m���ݲo+�1���i:(ںm���Ѷ��uv�Z�m�d1�R�4�	�o�~��U���k���Uh�pn*�W��Q���y�`��v��;��,��ӫ��7�Xۻ,�5���,��V�X6o9�r�M��{م��y��7u�/�V�Iȣ��n��ɥ�޼�`Q�� }��:I���|�)�&�hmr.�k�kG��������sr����[�Ҁm�ĸ7��{�`��ُ�h>̞,��:^M5(��SN+ ��?��W*�s�H� �$��Z��zp4�F���iA�{E1$hy�~ˌ;�0�;ן���n�d��r$�"Q�w\I��Vz�U�}����P��CBm�u�:�U�gu��8�GQ�q��Q7�1w5�ٮ,U�P�{��I����Ά�n�˴�r��wFz��x��x����}gc�m"-m�m�ۛ��҃���?_��@/縬Y��
4�I��ӔTM�Vj�w�̢Ė.� ��_�B��N4�8�Vs	�����ͮ�H�@�Q�1�q&��Di)�.L���|�\��v��VA�ƒ"JJQ:�������p]� �ݚX*�kEk�H�n; �� ��P�������`~{����߅	+�\$ώv��Gj�G0]4GF�c�&�u<��.����sA?���{�`_ϸ�]�; �� �uyBCTP�N���:�k�1w5ޤu�1wzWP����n�Q��]�v�� ��P�}�`wwi*I�I(�m��v��RY�8����\��o�R�Lf������N�ߺ��O��r�M��T�}�`gw]�wv��κ�Ҙ����d�tof���g�+ԛ	�/n1u��˳%�"Z�4DT�q��k�3�X���s_��U���P�j��$D�"N+}���3]���� ���r��Օ����EIJ�#��8*�(/��V.�pݫj6G#�)����W8������`b��f�z�e%M�T��M�K�6��~�r�g��$�y0:�������?��p?Ԧ�� AD1�(�
����� ��?�1P*M_�a�������%xxb)�|шu(d l 5*�� �` 	DF@_�Cq(.�AP!�`�( ���ҏp�+
��� �)�X*�jEvf ����PS��H0EEG$D A(�lt2�'x���]1��
��� ��QY �:������<��x(��DS��
��"���p�߯�G� G� �E_����`P%%%4�EQEU	@P�@J�*�P�@P���������D���(
{��`�!��EO� 7o���Ҝ������*h�7���"�� o��̟ԟ� �*i���؊G?�UUUTUUUUUUUUUUUUT�UUUUUUUUUUUUUUUUUR5UUUUUUUUUUU@�"(y���>?��������8��
 ��c���(��x�aO���2�w�?���@O�?�z*�PQ�?�Y��|O�	��h��/��C�?mO��1��)�����q����Z���k^x��Q���?���	6C���������|��������K@�д�
*4�P�RP(�H"D�4�-+@�B� �����!�@�(%%"� �J �"�
��
� -($B�@��Ҡ% �H�4��
*�R��.�ҨĂ!@����4�@��(�R*
%(P"%�@�
�D!�HR)B��J@�H�-*ФH(P��	KKM#BD�J��4����@RيdEHL14IJD�LCI@�@R
�B�2�\�\��	�h�(��i��&R`
B����B�(T��B ��2�J��H*1
B�B!JD(���-(!@%	BR�--3-,KBDP�!4$AC3ALDCT�4�AII3!I11JD�B����#�!4A,CD��(�J"�
�,*��,�
,�,$($��,�(��(��(��
,�,*�(�J"�
-(�H(��-*����,¢�(��B � ��B(��,ª�?���
�:0��3��l/A�d�������
��A�Aq�MO���?�?�j��~��8>?�����ҟ�B���?�����"
 ��%|p�C���u�?�������gŨT�����ᬿ���FW����������_����(���Ac"~�������������6N�?��O�TA�B ����/�Շ�?Ń�%-_�C<?����"~��?̿�ArO�$!�`�(~���}UZ0�����ן�Q����iP�M�l=��3t!a�Q�� ��������A���"��_�~����?����?�����o���~�X���i���1�b��?��ߧ�z�A�G��?���`AD�Q�ƃ���~�����~�����������h��`� ����qN�<O乇��n7������p�~��AD?�~\���?b~~@��h�Ӊ��_ "*��X�н����`��W�~�!_�0�0�8��{?j�/�����_����\'��Qѓ�l���y��!�W����R%u���]��BC)t�