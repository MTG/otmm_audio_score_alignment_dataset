BZh91AY&SYp�_��߀px���� ����az�    �^pj��X	PZʊTڙ$R RJ�Km�L�hQ@R�
m�A( 
�#G> �HT���
� �QJ�%@H�PP*�UQT��PIR��$%R@A$�J�*�RR��H�   � a�P=   
�=�
s�s�{�j���֜��^�L� �6��|���� ����z}9  ��4�+�ܩTa�WU�U*�R�LCB�wn�R���)N 4)V��J�rԥ*�
P3jU*@ �y    
  ��ѣ����۽7;��s�}��W�|Z���F�z�cw�z���[�1ݶ���R� M��nn�Oux�w�]�-+��r�\��w��k���Ϫ�i��Z���^��� y�z緽ix��nn���t�|}�       =�uZ{W�W6.���}��,���y����+Oz��˾^�yn<�˝�������W:���m�;x �{�<ڗ�������{ʖ���r��*�^��yy\�� =�R���qk�99�ݯ3�mo �@      �` >�jW6��m���ns��rwe� h�un[�z���V�wJ����p�gW��k�W|(������^]^��=���8wKɯ�_�-\�]��} ����˪�[�,��{�[O-ڗ��>�     @� ��-���vם�-qe��ꕀL����K�\����U�wŽ�n >��z\[��,�z   ��zw���+��O=�W6�m�,�W=�_[�������zks۾�����﮻���g����            S�I����D      ��dSeR�@ h   � �z�J�ѡ�L&&#M�2i�&"{J��(�  @ 0��J�M3A1� F`  B�T�L����<���S�g�����i��~�P�����ǡ�_���_}���׿�QU����QUڠ ���QU��E\(` O��E[�YV*�*����?�:�]�o���A�ɩ�O�C�������y�$Ns�=@u
u�u�����!�(~H����?��C���!���_�W�(C�P? ��?$�C�!^@�y�^@�H�9/ 9r ��NI�NI�B���I�����_��$?$S������?%N@r@��C����C�Hr���?P���!� ~@���H�� ~@��)�(��!�G�<������C���9 r���!9�^J�9(rP�*s���ɸCr�y!�W�<�� ^Jr^BrW�r��C�@�_�\�2����@�W� ��^H�9 r��^J�W�$y(rW��%y(<�� 9+�y rC���ùp��9�S�<���S�������9�	��'��"~J�H�H��C��)�9'����'�О����#���_��H���䜔�'!NBrG��K�^K�� �<�伅�%9)�NJ�s�RB�)ԧP��<���JrC��B�����rS���$Js��%9)�Oe=�=��S�}��G�>����+M�	�S���b.�. ӌ~��*��a�AI9a[�`@��
`!˷��ԧ���?n�֨��e��b%.ʀ�6ӒT4�hT�*��N�׌˪U�������dUFOՒ��P����D�)W2c+$?A�y�B��澼(69���\�2���V0�Z4�7n��ͻ��&�4�8��,��>��<+rF``�y��4�,̚|�f�=A�h�f�u:\��Y�LO�U�D4�pv�� �O�9e8(�L6�����`��9`j��N:��L�ΐ�	j��
sګ��Y��w�6f� �F���A0%Y�ǩ�X�H:� DL�upkm�y�,�B(�@k~$j4F�X�٩05��^�`i�k���՚�2��?!"�
%!C���h?A�?�Lw�@�Կ�2�r��I���0�u����0��v$FF%I�j�b�SN��B�;��a�����w-K�� �_�。/�P`�mMv���� ����h���̒s�#����hF�4Ĺ���]�8�Ջ������"�7C���zw�� � ����A�j��cO�dP'B�J����|�b�8��EQ�x�C�B�{ד�˺�ds�~�'5���7h:���LHf��C!�PI��u1�h׽fuׯː�%�����`m�"��ӫY%w�l��)(0u�C�p�`��qF�@ej���ө1Ѩ�2ă-9.�e���ke���F��)!���ffkwvZ˧�7RAIT��FZHp����	`��!�-$
pB
���;�@������d12%�0���[�nbsgC���Fà$'r�P	U*F������}�I�� �P�u��vn2m�������Z�!�a�3gTV�Ѿ���(4G���1�S�&2����d`�����6kFiud�rq��2LL�̌���Y�Ud�!��
���#�;t�%�N�uI�+P��^��n�r��z��ɀ��AՆS�F3L��Wwy����8[�5�8�b㓔��c"'��iѤ	�O�g��ә2$2�)�T8�y]���G�F���f�t��2���"��g�黎;B�X7-V#Ub��Rm��S.�ǖ�q�T�"Mq�B�&�ZgL�6� ����~�5������DJ!���`��
�|���
���R��@"�(�A&�&�)�@l�2�$�a�@[@T����9��f�'F��iu�PZY30JL�!(
�(��0֣5��4l$��BL�D�J�K)2��J�4!��)S��f*��*�b�Ͼ^
��:��~��R�1��K>�p',��x�)�@t,Q�]��-�9\'�|����5t�	H2�F���DӁ��A���:�E������D�̌8���lY�U���,����T�EE��-�P&�#��RZȆ�#LaF��3X6١�����g���r�c�T�S����A���<�2B(K�"Z<Yv�c�ֆr����r�v��iP!b���|�^�B��� P��@UDAwBz���B�Fh #8����zeCHtKf.93�391��π�0ۨ��3:gN�����`GVQ���r4kf7A�5�6Q�`�)U"RE-�H.:	J�`((Mf@U�I����c�|u�g]$��!3WV
ˀU��d8�.�e�Y
�p��AX4����+c�w�Y�����;7�dh��Μ�a�%!�e��`Ƶ�6yo���Y�쵽ˍ�2�il����"�IE1`��>�o�����Wx:�@j1M��QL�`)pt9vz]�^+��Wl޿ �,\�<u|U��B��#)_�����-�p:�ݔ�X5�)�	�J�� ~���N:�@��$���Pt�H0,��Tc�3I�)�jLL�0nۖM#`���& ���A�,� )�A4�T0��u�2�֒q��t��k
m���3F�0��F$�4��bk6Tb�,�����'�� �jAevs�"�9Q�S$�(q��Q��1s	j�0צfn�-�r]>:�d��@!�M&2�0G��F]�.��P(B%NY�����hN!���,X�B�C)��Y@<:P��}D� �5[�	�X��9|xF쳭�Y�u=�'X`DyaQ��E�a}��z��;���G��<W'�
�J�
�����
�� ���G��y���؅lu�+�,��]��M�U0͎Q�ǆ�9�R��̈��}y����5=BVP@g����|⁇TX$�HqU"h�2:)����|/�c���E�{�g}�j5G�'���(��^LS*��� ��O2/�]������B��:
�Ai[� �H���UM>��l�
�=��Ϗj����B�R�a4V��[���
�ݺ�*) R�Ց��A�,��A����;�h{�>�eL4�텫a�6I��2�PLfA���,�-"��'32q##�!#��E�FkE�����1��,5aZlֺ�x�Ŕ W���2-��7B�ʹ�sEw��V�O�S���fq�Y�=.��RS�x�)�|6N>0,��6f�ꂠ�W$5H�O�a��
�(����wߚJ<���&&BjMA��YI�dc&a�;��	**�Q�)��#k!IRE*B3�0�D����Z9�u	o��`�`A�d��Z�[1҉(~��U���(��Th�V�)������I������Į�w��Z���E��o:-}���tQ>X�S���X�2��0 ݁jL(����3(��:�$�r���t��%Aa���]Z�L�	�*�/u��4�������@�%���t��1����@+�0�A��h��{ه��:�Ǽ�`T����@"�ZT|A�h����!����,�a�AXn# ĺ�}f��DC�@N�"I`��i�p0�rٿp̈́��1+VB9e��R5J��H�U�X&�3��I��N�(ugWϝeh����.����&�����p)���¢*����p2�58Д�Qi�dDcb�g��с0u���O��Hj�̜(2��7	[C0J�M;�b��4k��:5����D��I�����Q�d�	B]�Д%	��MB�~�Vd(]N�r��v,��ؖ���h�F�F%N0d%&�(Jy�5�o7���S���uA�hդ��M���-��G �c<�8lp� ˮ
GºC�F��,�Ĝ��$��K01`��cI-I�Є��	�	Nb�\�Pz�J�e���u��o̓#
��X��PjC�0r���e����u�}�=[�N��OTA�2�[	�ˊJ����&���IN���]�zcDJK��QMђ�%�ui �0�3��捄�pf���ă�6w9u�Q�������}>��߅{�Y��Z���'�rK��b:	��4 !�0Z����Y�1|���F�b�ϩՕ��o�3{���̌�\�+[69К�-0�D�OŚڴS�X��0��<���?~�,ǩ?[�f,�k�r�(�#)tp�i�'(���3��j={���oZ(�(�j��!�#2p̰�X�]f�F�橵�Z�3vnp�fg�F�,X����Ĩ��j�YX3�����N�h����N��+,������R�����j$�,)3��߹�c�a��
3���Z�3}bDySub�d�P6�Y3]��f���:��O}�э|��l�3���T!IR,�C��0��B�DEGz�}���UL{x�!��r1(��&��n�:�!:����kv��nDN+�u:u&���}I�-k��4�֪15�F�32���c4�V�1٨�Z���h5�S�X�`�n�k^2}����vhߝ|z����9�v*׀������'@�!�ȥQ� &E�P�`]�A�8�587�
0�T�t�`�%w�{��g}�mٹĞ����
0�;�tx��3�uD�L�l�o12�n�mZ2�Y8]a�e�2E-���w&A���E-N�r,�LkS�'4B�&�E2(D&K�('�.�Z4Z�X0U0i��MS4�f�#]�l1խ�N��A��䘙�0����&L�V�39`�i�t�*t��dp��Iv�$���-%3,J
���L�!��S�˲	rPI��@�^tpc��\D۳�&@&���\��W�C`p��VTLiRᄎ!}g���OG
 �4A�	vŐ��)�­5~=|�
�Hۜ6C��^D9T�����a�)��
�9�T��
��}K����Д ,��Q\
b�g�� r_~���P��P�`�%	BP��'PgAj5'��|{��h��0���!�	v�40C��1X�i�y����c�:׌k{vFhٽ����H$�O��)@�nLL���d㦬C'���N��j0�j�)q�r�\�!�N� ј8�R�+�֫����yַ�f��`�m�(J� 0���15	c��i���ֵ�`�	���3,d�r��Q�n3ӳz�l�����Y�Vm���ѹJ:z8]�SB$9b��{��;�@�l�d*�@�)�N]7�Y��㒮��s��d�еP�*�D$�D�By���K�\��4H ��"h�]����@�q{�q(�G(�P���c�*4_o�]�b�K���0�XL�jK��C��5�t�r&;�H�����:�1ߍw��:X�H^U�@���5^9`jzFk��7�C!(�����剢5:$�L��I��ڝ$d9;��h5V���Q���u�D�V��:۔�i�>��BR��ȝ���)�%��;��3��[�����Q�Oa<���{-2kQ�F����0�Z�4Fj�:�tړI��k}�F���[2:�
R4�f�,��1�
E����m�����d�yhܶ�,fd�)�ƀI]��7	�D][M�l�2eܴ��r��UR���/\�
-����pK��Ď�d���N'e�؜�&�Uq,aw�:�o�#�.ѱ��K��sg�V�~�ΞVa�.̌�$�]V�z��`� �`Cl`
����Р5�*�nӏ'b���`�� Xz ������m�p k Z��  �      ]ypm��[Yf����Yr�$  6�ڶ�R���` t�S��       6�  r���ݎw��uLj�u�Ăڰm�mZ� $�`�     6ذ�-��� m��8�arY�H  �� 	��A����/i��R�	25\�8j�	
U����Y`�P )T
�:�����	 m��+5����-�-�� ��[Cm�$�h-���GY.Z�7|�}�v��vU����V�[��N.͚�c�T!4��[�v�q1s0p'`k���g�Z֮��v�  lmd���.B�j�ZU�`[@F�K5�+6�-�n5i� 	 6�m�n�kZ�6���W�G)�v�@mP�vG�$�e(  m�lH9�[vݎ 6���6�� �)�  z��5��a�  lԒ`.�y,��#������t������^��� �����[�V��UjB�[VrvrPMJ�C��v��U�;��\�/5PkĊ�t�4uc���;UM�8-��VV�d&ԅn�qǮ�N�R�hiL��U8�b%����s֐#R�ח���e���J+�g���o���n�xW�Ũ3 5V�qWU�ɑvi�h��K|�p(�����l��U��]@Ht�*��:%R@�� �K,�mu]�e�6'U<�C��q�46�A<�P �v骔��t�9����VH�3���V)j���W1�r� j��Ά�t�mm	����6�(�9n�D�[v	 6����I�V�6�`��Uj�K'^[RY����A�:��X�k�'g����X���jn�6��ڳ���]U�j�e�n��m�������:�OIv��(�?K9O����v�b-�q�v-�.�	�jڸL��lT�Lb��e�Hl��n�V���g.���k�nv��P���ص�g�j��zڠ:��ƹ��(J�fX�ڀ��������i�#��l�<`�XpmҒ�J�ؔ��k��dYl�ڇ�����vY�����t
�����1�x�k(�Ϊ���d�Q�t&���<���µm	���,DՋ��Zv�)��8�&Y�(�c���h�����> myoZ��:�oSe�4.֩�a����@A8��,*���$����Wl��P.��N`�r�ʹ
����<vENZU�%���uz��]�65/\n7H}+F�j�Q�r�U&���qaM�!4�դZU�.���)y�u� $l��L����� �P��;;Hl��q����
t�j�f����v�ӏ\8 m�M#%+�$6�m �8 m&���ڤ�UYZl��UHX ��E�l�[A�մ�FMU�v�zN���"��<�(KUUWP�u�� $�ڛA��mU]O+VѩW���W�FRWkh�ڐ�ZkXI��-���h�*W�3J�P*쪤��v݀[v݂G[!����` �  5��e�T�ʠQ��+�R��UU�J�� �J�QGV;#��l�lkʝ��J��J��ύ�ۇ�ڪ�CK��-��m���  �    �h ֖��&�ж����l ��d� �n�' ���}��v�6� l��p�g3K���,�|2zT�V�L써嗶�=q������٠�
�h�	 8m��6I��m�	e0[��  $6�d�i�нh����|[�u�6r�7�]�ks2�l�l@  5�m��u�qa��+WR�瑶U��U������6�@$M�Vk��
iM״P<T��5�Aղi6Ը�l� m���KN�h�-�sd�i��ջ�mZ� kn	wK�C 6ۋz�P-��m�6��d6���m�@t��shn��[�Hqb]'f�m�� $l m��LVҴ����gF�U�Vѣ)n�M��! 6�,�`Tv|����U�E�*gK�c��0�Iӝ7$K�m I �� �Hn�H �  6�    l��	;E&����Ӏ�n�j�lt��Z�� �un��R�^���E+m�� n�[v�F��q�U\�P�fQ���U�  �6ͥ�2۶��UU�x6�W��Ŕ�^�������2/�Vی�is��R��[mD�al�C�� m�`7�` �   $[Kh��)��Ԙ�� 2@*����TP3�
�M�[D����l��H����Y�^��y���dY7[�K�l V�BL��U����V� �j�G��pr��h4驶Ҽ˔�C�f��d�#m�;k�;ei�O<����
B m��Nkn�����jN�M�YƐ�S�n�m�� ��q�Q��/c�Ĥ�sEF�A5���2k͜9j�5��)(��U^m��j݋*�98N�����l���5�XI�u[W"�v���rj�ƼcD�N�����wN��j��WL㱳��W��i$  l ��[@ ۶�	�\  �{��   
�
��B�6CV� (	{�W����ؠ�i�n�iV*�xNKڄ��+͔cB�VQ�d��mͶm��HUT�%�@�6�jx.j�mm��u�������A�`6��Z2m��������[R�k�IB�dQ|�0��eS��i�8����,� ����)l������AeV��	���[R2�m�  8  p����ﾂs�D��J�eR�Ҳ	خ3dä�]�v�@�u����@���u!�e6ͻ^)�=�[����yM�jm]U�'@m%�N����(��\8p��]z���\Į^��y��]s��k2��o7b�Y��vM�t�[���Z���Y��J�t^��g�U\����`#�Y6����gq+�8��(r3�沁�p���B�l�f�X�"%�����m�0XݤY����s��}T;v�X�L�Ջv�`���d�$���m�$	��B�m�`��U��ysMUuR��T�S�����۴�a�I��n H�ɻ^��� D�ݵm]J�:/<!/2��U���<��K�/2��M�EiK�q�һ�T����U�U*���YWD��i�v鱶Ĳ�z�-�$p��$r۶�]��XZ�����Sm&�H�5t�-�d	6]��,v��[�v�VS��[���6�e� l��]n�\ �n-��Y�4��g���vQ;F'��*��e�8�k���6m   :�M9��G4��f��  m���Y��k� 6�`-� [%m� [v�  -�GW6��:��� ZN��  m�8����F۰�(n۰m'l[@�d�$ rާ	��` �$Im�E�mm� ����.  �m  �U�UǻC�c�Y�ʳE�`-�l$&���iYf�o� -�p 6�m&���L < �ۦ�	6�0 �o\�f��$R�N�M�zڮP�[�or�R(M@�+�HS�UUQ�ŝ-5��t�� [@�� � ������WR��WM�-�f5+ J��T�$��*ˮ�ݛ�ذͶH$z�m�J���5X�At�J�*�����N���U[�j�K@��m�C  l���HpIz7i��Nʠ4�pԫUU@@V��9����*�4ɻY�k&m�d�ګ!@Ĵ��)g,9٨�ȶs� h+Em<�N�ݯ/;�ʫ��X\�'d�1��V���!��u4��[ն[Di�[@�-��.&ܑqU�9p\ʿ�b��� �� ;j=iT�0h�u��yoK�Y���  ���&�����]T�ei6�,T�=$��=#*���v5�h�J��q��i���ዃ'Y�7��0�C���ݗkP]@�J��mUs����#l׮����*��6Z��U�c�mJ=���h6�̀hӫa�%�����Z�� �8�u^���3:kմ�Ӷm�ؠ  l[[l8/����8�)W�[��򴫧��b�%�c��geZ����6׫m����r�'`-�ԠE����b�Z�-UU.^������՘[[V�h  .J��-6m��9� ���[T��U�N��S�{���Z�SI���e��v�u�� [x�{[�E�
���nU�Wۢ'7J������  � ��*ݶ؝-�n	a�6ۀ"���@�`6���"��pP��$S\�R�7U.��@WZ�vB;`�z��ن� m��M�.֥ ql��vHJ\ m����$ $���� m  �Ymm�	�פ�g���@[@��Ԯ3t �u!�t�^�������R/9�e�6�m�$ �k��N��sr�l22��UUڎ�����s��mr��k8����b�B�O(�S��C
��diI�wbd:�& 7cm��m5.Ɗ�ݧkc`�yk��R���kl�۲������Z�����W����Q  7�~�h ���P����kaAUIAE�%�T��f%��d��b��a�h ���b ������fՂ�T� ����_�UQUTUUUUUEUQUTUUUUUEQEUQUTUU5TR�UTUU �UUTUUUEUQ����c�*FDO�	�`/B���dE�q�T?B2.�{��0�'����lE�A��<= 4"�@��8��CB��N��N��N���!���H� H`h Ї�thS����F�%{T"�U^�O�Lt|��
��#��;�� �<�@�� ~N��޺�C���UQ<���N��QBH�` `y�G�@�ID��&�e���ҟa��zj \�J��6�=�^	�� �P��QE�E��؁�B�`7��vߪ.��	�H&��ͺ����6���0*h_@�)\��@���z�$�II�=�W�U��= M��n�)�`�i=P���>E�q �A�]O _��C�=��T�>���E�6����(^ ��O и�x|	��"�����*��� 3m��a��l6�m��|��ʼ�ʼ�ʼ�ʼ�ʼ�ʼ�ʼ�ʪ�����n۶�;�{����*�*�h��?�
(��k��������J?����?��Z̬̬�����z�d�Q�4�QE5�4�!M%E%4�4�D�P��
��$�H�	�!1�(hh))R
�������"iib"�U�+��pJ��b
@���\��bb��3�s��%	@R�U	�TqEa(ZV�,�� �(
ZD�J\3&�@dPk
4�"X���MQED�U!�
*���&����r��KT��ve?�6-��}�彡�<��ӱ(�T���ۍ`�Uyj���2���=�W着������C9�� U[���H�S:ֳF�qduJS���!h&+-�TUA�+ %���F 2*����C�(�)�=R���,ceiW.�J�%e)�$���_����n.1�ve\�v�TFy��#q7UI�TӅ�nW؊���[dh~o�_F525h�蔳:��;o���;;[�#�%��<1�tf�u�u��� m�6n"�5�.�8�J�	�ݭ.�Z�7���0������#��Fs�v�u㬲ٛ	�ͱ�6y]�n�K��!ۍc��vϗ���!*�8���a�I��<r��Oh�.�J���2R��Gv�*�A'�ٌa�j/�9���k5UP ZBT�ët�Я�-4��PzF54�;�y����\�x>~TI�t��[G.��Jj9�!��J�WI�W
ٹ�Iv���F5�.�Pm��؟7`Q�MM*�շl��oA�:D�X�s̳���N�K[��VBs�TAfxYT���`�ڤx-[ʬ�TMI�I���\b������s���ٔ���ZZt��C2n
Ln�ӓ����imM*���:5�C�Mx�E���Q��5v�:��Z�:�\P�sk�hv����ƛ=�8��v��g��'Ny�3�]��-�;8ӳ��5�x�2��qkw�ߍ~?�y�R,�U��`r����t�ݭ��pn#a���ԛ�/0�;����ω:��m�	%�����v��#�E�d�+d���Wj�m6��4����@jΉU��������?R���+S:$�zc̮om� v(�g-���z���*�mpWn���Q��$t�	$��4a��>t��-� �rv����%�EZw����K#��(s�;�͢�%�����ux�r��� ����wrp-)ёl\�2�:Ⱥ;gY����%mB:8h���>�I���9qj�h��h3���ʹ�+����BU�wQ���ܢ���K��+Nāѹҏn<�;n;;��8�#�2f�uΌ���N �)�ڀi���4 ��|4�H �ạL���!(�|�B�n�0CE�d�5�w��[Z��G�X����gW��]e�:>��6tҪ�^�:�q�]��m
�R1=�,��:x��������d�	�
����Aa���ꀟD��ut���\cr`жi�Ku�-�ض:v��N  �
ݿ��o���ڶ�ip���qf��@�G72q�Җ���v1@uؘ���%�]eݖ�FF!�	�ʈ`���Vp:��gj�pe�6O"�r�1�\c�M�����>s��{(��6�WRAD}�3(>o�@���Y@��8�>���:�T:$B���i�J��H��`w�H�n҂�r�:�"9!.�Ϸg�A�ɥ�>��Kw�K Ͻ���F��"�U`%���;ݮ)��E�������(%&���VI�}0�'3��I�s%����+$誠<2 pi���ΣY:�����-��^��Qv�{pUQ�c\�����9$p���M�N �޸���V�����E�
wUG(�P5Q����d���K�U�EU
P����0��n�Ƭ����s3,X�c�J��UN��*I`-�f�y//Lvv�%�ͱd��j�d�fL�R:��R�I�����`��v�
=���=XV�Q"ѐW,�W��\̝��,�urσ����W��������&"&���Ӵ��8��LE���,��ѻ=s	A��r3+Y��ܡ#� >�t�=��XW�֯�۲�>����q�RI(E9,[J�橰5m"�3�U��&F���~�Ԥ:#�����U�{}4�N�H$d DLR�5��`{�X^��9U�n���2z�H�2�u`j�E���We����S��TN�jQ*�,=���K<��b�zi`m-���%��Ug9��L�ܔX���{h�jv���5�TT��D�P����"r��Ȃ8�rT����i`gޚ+ڽ4���,��� ېn��R�r�U{�i|���X����K+ջ�d�:$@9ڕ��}�y�N��uS,�6��ƛ��$���Ͻ��϶i`gޚX|��jO����ڰ�誣�8��NK�l���zib��j�3��`j�KV��UNT�l�*�&[�y₉�.����0��*�&��ho
�z�TS�m
:��`g�4�j����=�*�#=�M��Ӌv��A"��(��u%q`��z� f�T�^��H�E)J*�8�%k�vK:�9��'6��,�WU<#�*�n'�$V���u�`����}���|�e��~�7(�өR�I ���f��9v!�s%^w�tv��&�"
�(J�"�e�c�lD�RD����f}��\�'X�� �K�	GD��ܽͪi7�d$�893		r����^`�2��Y'��t���n�̒���e{s97��v�;&�.J:��.�,�������pR�al\3�ܰ��;���7T�z��c�;1í�f����GkE�'D��t���J���-ێ�.n͸�G��� �VӍ[�6��2m7j�m�ߐ����i��n�$}ۀ��ѱ������<̽S+�v��'e���Ӑnڐ�!�T���ݺ�s ��,w�ث;�dl�Jn��T�Z��v&{}��y����e��{*9��$����2�z����̺�s%g�<2"T�aB�RX�
�皫��ۮw�+��e�>Y���.�6�p���e��Vs���6�څ�t��G����R�����
�M^�
l:�³����q:[-��g���R]w۲���X�|��
 
�k��ۮ��ILd$hn)#�%��m��T�`�$���5�N�;r�A�Cz���m�=�6�Q����Dю&��=���]�]sْ���X���(������#@ o�n���^�����z~����(%&:T�ZY��^�{,{�x@���8����D���\��^�i6��g�y�)C��Ѱ�)��{��d"�DK�ɸ�C�H%9+=���-w�1�5��%g:<NDR�S�(Y���;��]s=����X��$R ��h���{.�罐J���^��X
��c�熳���ܢ�!��
%�;��g��{熻��X��̒'#eĚpE$rJ�wX�W�P�w]s��Y�?��~�1�W��Z<n�W�㱕�^t���k��.̇n5sRp�H�\ggT���_��U���\a��UL�%PAUS��R�����ޥq��R������I�A�Iu�f��w3����;�e��-	Q�*��j�S���۶�{��-�ߺ���S���6 }�`(k������aH�Hq��19c���Z7}�3���?^o�ׅ��A$��	�N �m��V#�Q�8#*� ���&�WmzQ�Wr��$�e���(D��u��9]Y������c�a��4\��!��E%�3223;���c���,s3$�ȃ.4�I����e�{`��]s3%x{�ƃb�NH[�K��!g1�]s3%fw�c��0��b2�qVg}�\��^��e�������u������'��V#j�h���38�A��u�]�\��u��I�v�����j�+��@��=�N�vrrX;v�#[.9Mɣl��vV�.�I��W�D��d���g�;=�lYwg�D�裠�I���ծ�w1�kv��]�<�/ghΌ�]�n��ek�n8lk;u�8ܘ���6��ny�Jƙ��r�Ͷ���qs�qr����b��۴�Q3"M��H��*P�� ��{|ƌqQ����jp��R��ۇK�!��ݵ�Eh���o�.qu��n�\��ϱ�_^-W��cD�]�-�5�"J9 @���s.���U��e�32W���$�$H���/b��s-��̕��e�q%�14���@�i�9��]w3%g{�c�^�C3��L��H!����fJ��2Ǽ����̱���0�(of�M�tK[NS۞xf��ۦ���M&j'^rŽ��l�rST�=�B䩫߯������/b��s>B�r����ff����[��kQ���}����EPB�U@���|���egs�c��x�)H�"�-)g��u�̕��e�{�g~�)�U #�_����s}���=+=�e�g�"pF�N@A-�;�32]��<5��e�30A�(�e��p$ �2�0Ŷ�>�qy��{h�לu�<uu۶jyn�z憻�.��ĥP���=��H��}�]��g}�0�fD
p$�A�fw�z �(�݀n�6��^ŴF�������B19u�ݕ��e���u%�$IF�I��N]��*��( $�j(�����\�^~�}�xFV�kDc�&��#X� Xf!�q�79'g����JHa<H���ç]ya�OM;�H*A,�1�MQ:u���]Y�E	i��P����3[?��¬��)��*�vJL��Q=�»�2�c������3ĥ���N�;��=_��Jm���6Y��y�=��i`���94�5�S`����,Y�b|"��z�:`��o���������6tO���C�CoK�.J��P�J��J��x�8E��A�P����!�Ew�纶�>"�QpƿNH�ϟ��DТE~��۪��]�ۑ�� ���#�XHM�d҈��H?{��Ҕ�u9���|���
� j�g�K��j�no�"(�␤�[�,��D�Y��
&�+}��p4�s��HҔ��������?����87BI.��]nzZ�8�F�V�7g%;�x��1l]tL�ED,�^Q�U�޷�JR��y·�JR�����������T�<��9���R��Ep|sO�')�FLq���������|��S��3�)JN{�9��'⁘4���?+�o[��M��%�j�4>ş|�p�j�g�s])J����s���(�s��HТhf`��D`��
cwdWP&�����JR����s��R����7�4$���:%g���9�$����ܟ��o�=�R�~_�u�E*��(��H���lWP$C�}����/~��گ�{��};�/��T�{M#�ER�$e��s�� ܦ�1�n��^M,eD!���p��>:z㡾�JR�s})JRs�����Jg�n�5@��ͱ\5@���͹N,�`jH�T	�$En�f�\5@��Q�׿s���9&s߹��)Jy�se�j�"�g�ZDQ��$.�}i�|��>���)JNs߹��!{�@��|�JR���{�4=�R��k�l�ħp��r�5^�4���w)J^s��JR���{�4=�R�}�wT	���f·#!�\��+�JR���R��� ���\���C��Nk��t�)I�{�:�(���
1�p�ZC��q������굮�8�zE���g7g]R�r�( m=U�3O	v����OY�f�&WYnl�'H�'m����X㲼�:f���&gIj��0�uI��1��m=�P�v%'E��"^�Z��tb{2d�77m��8wþ^������,ʕ�J��Ò̪�e�:x6��B�nM�'THGn�ӧ:f��؈���F�Ͳ��hz�{06�$���PB��Ŏ'.ᴉ���`��G:�n��ܴf��ځ� b �2H$�w���s�ߖ^���0�v햿��m��Òsߵ���JS���k�)JO����{��/9�o�(N��Ɲ\3f�i����B�j�5C3&� a�j�4��:�)K�s��R�����Cܩ5CV-�j8�U h&�(��M�s��R�����JR�?s߷�{�&�g�i��MP&�����Q�����o��R�����JR��s߷�{��>����JR���}·�JS�}ηR Y��ԑ�.�T	��3&�\*R�{��t�)I�s�t��)y��u@��MyjZ݈�I\�"
|Zr�jϫh�g�za;\q�e�ع�ܝ���p��22��Ir;�+��T3�4�P2���>�Cܥ)yϹ���(y�}�"�j�5C�u���ĩp���*Rs���q�C�]��J\���JR�����u�=�R�{��t��!���n�!|$E�ɐcRX��MP>�s�})JRs��|��JS���*�CwslWE#T;�4�.���$Y��(Ns��5��R������9JRg=�:�(:%�9�o�)A49�OTE�-�1\�+�����7�Ҕ�>�9��){�g��[�JR��s\�p4��ܷ2�ݫYYkkr�c"!� �s�[�]<i�x8*�Ƽ��ڱ*���wx�����=\�����o{�������{��/9�o�)JN_s�گr���}�])JRy�ﹳ7�6e��ٛ���=�R���7���9�l{��>��|�R����g9���S5@�sd�HM$c05$rK���^s�l{��>����JHv�=���£�B��f8�� $K"�����<8 }�I�?;���R�����JR����i��iIf9��T	��l�R�~�9·�JR<���J[��j�wf�\5@����=��"B`�f���JR��s��{��K�|s})JP��7�{��>�_sz�JR����po��1�l�M�#e�r%N�&T��t������+�h��f5p����w�Q�b@�2',W�P$
9��]P&�9�s|��R���}��Q���׶+��T;�4�hȜ��%�'=���=�� �d�3���JR���s���R���9�� �*��,��Ĕؐ2��"�j�5Cf�)JN{�9��
�2R�\��R�C}�4������8��5N��o])H�������)J^s��JR����o��)A�C���=Q�tP���+��hw��l
��(�o[�Cܥ)y�s})JP��s�=�R�}��t�%)3߹·�2��
c����p����)�L�Dv�[�G��g����l��&smmx���'nJ�mA��9T	�$E}���������˥)JN}�9��)J^s��M@�E`�Zr6�NF���vEp�
S��.��I��$�����Cܥ)}����R���3�懹<�%39�g6a��f��6ff�t�)I�9�t=�R�����JB$�?5����)M͟��D���;���1�)�"��ܥ}	��o�)J��s��)O��|�R���6������Cܥ)���&�27N2I-�u@��Mջ�r�� ��u�t�)I����·�JR�s})JR~�Ї!.�]��?�T�=���)���r�S��pV��<[Y�_�m=�����;p�ղ�&��p�{rh��qH��v*k<���ʜ�Գ�*uD)8� 9J��m��Y:�n�3e���Y� #>|��ʼd]m��ǫ���n;v�;Dm4�^���nQTxԯGV.uR�KR��:�`��JiW�[g�]Fխc/n:�
��yw=N�������ݰ�s��ۀJ�^9��dus������,��4c\�ڰC�z��͋Z7�U�u�r���~s����)>���C�1JR�\�������k����X�dA�	Ӂ�[��5@���s�r�)y�s})JP�Ϲ�Cܥ)�{�5Ҡ�)IϏNk�����3ލ�����)J^s�o�)J�ߵ�`�(�R�g�s])JRyϹΊ���m�T��mA��.�O�(B�d�������R��5���JR��}�t=�R*�s��@�4<<�kNI�2��
��̚n���O9�9��)J^s��JR���{�WP&���Qdi�i��h���M���]wi�n:힗8f�iYJV��[�ܤ��A	�B���j�4;��cܥ)y�9���=��~��s��JSC�ɦ�5@���:��"�����R�����@~�x���ސA�5��m6�qLWpg�@�z����9)C�k��{��=�ɦ�5@��ݱ\  MP�h�r4�i�H���T	���c�B�j�5C�}�])@��߾�Cܥ)y�9��������-��1ܴ+��(}�|�R�����r�����R� C7^Mb�@�j�u��"�l&�Z5�n�JR����t=�0�YG>������i_����Cܥ)�o�J	�����F�`��F̈&�D۷"7$Yr�t-;��%۱0�M�Y�Ѹ�������(�mD���J�y�غJR��g�懹JS�~�.�iJM��خ�N�C�v�*�*��2�ΐ�2R�/>�����߷ˠhO|���{��<�������z=��RjB$j���\5@���d�`Ҕ��Ϲ��!�!�Ђ�� 3�c�v)�\�~���)Bhx��~��j�5C�ε�D�r(C+z�t
���Ϲ��)Jy�9�Ҕ�'�g>旸As߹���);籍L!�H�BE%����v���*/>�\�r������JR�C}��+��"��i��5�(�i�S�r�WmH�=��@���Mtlr�^��2"q�����d��Ġi8�D) ��MP�y���0{��=�~�R����� �)��s��)JO��dl�ktkz3v���}`�)Jy����A
O��9���Cܥ)��GJR����s�WUP�G�6D"���"�CҔ�=�9����O~�::R�J}����)O~�|�R���ǿsb8�I&���
nX��H]��T)J}���)O~�|�R���Ő�Qߢf8�!$�' S�H�����[󾇹JR�����vl��Ѣ͛���l�JZ
}��^�(�'��_�JR���~s��J{��)JO�9}���kYoq֍gO�/,�p��w2�\�q���5��M�[@���kۍ~:��8J&�D8һ�+��T=�6�JR����t=�R�}�tt�)H���B�j�5C�[J2�2�IHmJR��s�t=�Ҟ}�tt�)I�����R�R����tJR}��f�܁@�,��+������X@)K��9�ܥ)����Ҕ�'=�m������@�qĈRAuB��H2O�}����(��~k�)J{Ϲ��)A�$��~~vt�)H�>�|

 q�1ܴ+��T<�����(� ����R�����ґ��ny�\5@����L��I��M����a��B��* 8T�4FؠD�3ZD�i	���+��'0�f�N.I���j0�P��ѐ�6d80��R���@��H]`36 $�ߖ��D#��rB	c,]T�E$�QLQ1yHvA�1�!��))h��f�����F	��m���t���3�b&�η�y�FZǥ̞��/=�я��D��RM�G����B�<�����z�|U�D1Q0 A����J@�R��
M�]>m�Y(d� �wí�|)=v��""�'J��ɕmVW�~/�q������Ǒ�P�h ;PV���$�i�` 1�^��H����J�@l9eZ����W�]�}J��` �IWm�=:G���p7��*%�]H:5KPu��KT�)�+cJUd[l��;l��d9��:"w�n�IW=n�;Ps˴�G�h��xpaj]�a\�V�gm��v�:�gsPtA��xp u�1�s���A�W��:׌LU=H�Z3��n��5�@�R����*�y��H
�k��i,�̝��h��Ї9omnǊ6y1WYa^��j\ݭw;L�#�F�P�1���K���k[`�x�m��2���/���Y�`g�PYJT�6�ĪS�q���2p켂tv�� 2��DE��KZ��ͳ��`um��nGUK֓�d3p�H&a71����ݰX:H �:p�!�+�j̷i�T�+q0C0$�m����:�Κ(
�]�\��m��n����s�$Nz������ukZCY��6-����eT7XW��6�E[S�2D�`AW'0��\;$�Ke"�:��5u�Ӊv9��Y펶:��vN���T����cT5recv5�E���nY0g�#�����!\�.Pܜ��mCi6"]�(�''J䬫��Ƨ���gp��[\V-Gj���;s>�+\�wM�v�+ q�.ї�����t�Bm���wm�s0*0f����M��[+r�쪫u�$˵�'sSm�
�':�t#2�LAaV����"c��{IĠ���SUT���)kM�2.��q�f��)q��N!tYQ�:Slմ��ԝ8qTKW �^&�'A�k�s+�ᗦ�rn:��mN����w�`q�-E/m�0ۜ��i�6���-m��
z�fU��lZ!��c����>X�q�;�ƯHޓj-�ޜ�q���`�q�Vt�gE�Au��d�Q�Rv��b�.���Q�)��D�ax���g�����Z�;m�ӕM�<��u�9�t���j%Da�d�.� �IA�T����<�D�A�C�/��{ꇪ�����(��C +��"�o�LR8[&KWvLl�.;y�WTpS��ϳ�3��]=����~�p���1Y78�ը�Î���{)�� �rvV�[v��j���8�O�S�.^�������>!p�hy
aA9lB��5q�A4qU�F9��"��޴m����cGT�o�G���:mm��g[�,�;�)+jn�=�Istn	??w�<}󪱛d�k�v�S�=Y��2Z�Ѩ�2�3����b�#��C�Αr�	�h�<�\=+�l	�߯����f��IQNr���W���u��g�{���o�9�:�)O=�::R������{��5C�ٮ�5@�����#I�Ke�g[�]r���9͝
R����s�=�R�{���t�)I�y�:�
hwvl�@a��TF[��5@���9�ܥ)�{�5�_�L3���~w�^�ϬY$罏c���,�D�wk����*e����u;����Ss��\u�q%m�e@���'}���'��P��� ����J�`v7��|��&bk��=&�X�������m�z�<t���n�@����e�ė�wj���4�2��/ �w�,=M�ԩ�}�ё�D���� �g�m8�)a$I��ݜ�(
���)�(D�b)�0"��~�Uӿ}0�'���8I���)����((`��,��k��n��:��f���r%7q`f�np;)ԤG*lQ6��X$�#>����j�7ս��K۳��{z*NF
�	R���T|��Վ�I~H���۳�7�ـ�WR���l��³[^�zw	OcU=��i�I���=��6���I������7qڐ�I�0��(�pY's6˜R�X�yﾃ��"":�z��>���8	��1�v�|��'=�M�*�" ƛ����jSl��#���]θ"�2�E��,��������C���l"�犢#��ob �����o����}ܣ��AI�T9Rs�����
T��,��Ϳ�	�8�U���(U
}�۲O7�q8XMH����7����DA�ک9�:��`OsvŒw����f�2�q@�=���
��Y=�\�us�F��$x�-����wwyk����TQ8�A���`׽Vw�� �7l]U I#=皸I�� P�P3#���(�u���� :����'8�&������&�*T�����'��Łմ��}31ԩ�V���G^=�(����(�pY?P C�wq�Ӏ����V����E@||PDQ'�?HA�>`ߴ߹�I�}����o���[�k���'69�DDD�D/<��o�V�s�o��~�߼7'!�e�L�.�:89�Z0Q���Qg����Wmj>�������
�'2n.	/�8V��RwW7u���$�{5�-s}��rI�Ȑ.MWp��/��A����k����ju��+�ټ᪠N�j6�q��q�NAd�\���wU2�">�=Z�`���#~Ѭ��PA
���Z �[�du<�:۸����i���N�&�T5U?Dڦ�`w����HI{�����|�I�d�d��UU@�}���T��IݵȖW/V����O����	Ғ�f�Œқ�5�a@�H6'�̏-o&ֱִe���&:3��֌ q�8��ٓ'U�m� ��
�*l�ӵU�n(�Ҝs>�y�Χ��7M�@8�nݠ�.ڶ����Eeq��1*k�seE5�`*�����5v?���v�go�5����U���2�|��)�΍�7n�(\p��L�  W*�uHYF2.<G�ꫮ6��IS�E�m��61l�W���c���,d�E��w|s�}rї��v5r����ń���:�2�" {��`mwIR�%)Q��`wޝӟ�&Mn�XI�0��/��uq�)�˂�M˺�>ݜXo�����w�Xo�u`\��(�UD�"����ﾈ:���:������>I}�8�3OoC��	J��2eRw��~���\���ju������_����k�;5��-O5�ps����9Ӣ���uUV�ӞUNپ�ww�����Q��**H���u`�l��+�}�����O}�b��ݛ�����S	�"|�Y�^{��u�&��������;��$�g�,����\�@R� G�~�F%*�n$��߹�O}�b͠(,�u`�X\.#�9R���d��5���v���S,>��S���IR�5	JF鸬�[��s�7U2���� �N���J>O.'�Hi)^�u�n(-i/\�9�;k��D�L\GeR%k�#�#�%U��e�˵X�+f��� �$�=�}�D�K�� s���2%IPp���zky��}ԝŀ�]� �T��">�\	,8b	�'8I�fزI�{f��US���+�&	}��}k���uW������;��5�DRNDRAd�(������^��G��N��m7\���)�p�o,�>��,�_wi׀wS���>�~l�=��rBNW9P���P�6:ݸ;y^P�ű�1�ī��rE�S�M��0�����>��� �{���>ݜX����ƩDQ��}�֯E@v��2�]y�}VI��o9�R�s_��`b�P�$m7���_��S, z���;�-ޑ�%SuU��c�� K��Ł���p��ͱd����U
_�N_Ǆ��rx��
�����j��o0��,�m��'��M�G�ѿ&��q�3k�3�0�;a��V���8���igd�u�<�)�G@�V�҉�I(8b
I%���}�ŀ�v��S=dG�^�� �����8�**H�����/�>ݜE�K��w �N���DDH?yϣ����ک#yf ��?�����~��۽j���_�:��p#EO�6������i�ԝŀ��fԩ�j��q:mD�ʩ3 �w����s�kt�^����2>�� �7������Q���]�Vښl��� ����n��1fr��u�t�m�4$'XHaOn9b|�y�ݕ�E��nz%46m����M�l��n�厈&:į)�mvPͭ\�Ƹ.��Px�G�jKC[�RS�㬽������ٟ=��M��Rq�Sۦ�lэ*�����Ѵ��î�4��k�m��n��Z��:A �ˉp�9Ӷ'������{���~N����{EȾ��̝n�Ӷ��閰tn��`{zj)@/Yk3�ʾ����Us��Wwk�� �T�c�S�# �w�Xn�.�� ���wM�ˬ䩗��y�u'q`.�l�5q�O+鐨	*��j�Od5����]̽+���M6OQ�i���(H"DI+0���,ԭ�R�X���"{�߹�O�o��m�i1!@�$I gW��G�}���=��0��,��Ե7�bS$�mR�q������q�v�+`Uc������\�-Oe��ݤjZ���&r�p�X�<�;��_��;�5p�5b͐F �*�n���>�}�ɧ�����gc��E`H8Z�GDĘ�$Q�9����e�b��ѥ�HeN�D�"�Н�
�Z��GU~��~�	=̚lB�$摛�7e�r�q�p��ͱd�������P"�P��gŁ���ـ����*q��n���H޻f���
\���������$�,{��8�U�K��t�ـ}�8���!���I�X�`
#a̾\��i3lKO�D���\'�]]8�]��n�������X顎�wx�����ؒj���fԝŀ���G�R�X���C�@ԊU
I3 �{�X���R�X	�3�}��?DI��O/�UT�R
r+ ������{vqc��g�d�%��m�[������4�
C��~^�6C��7T�G�]2�E�v vR@c#�EӆՊ�fQvp����C��x�o@�4;b׊$�o��Q@R��1.��w�?/x[�<:��M1<@_�C���<볈��~�"�C���,���y���4���������'�b���MzMH�r ���<$�T���F�7qa�o^3 r�t�FT���&�nv�f��oZ�;��� �����n��JQ��8CF��
���Zði'�;�vϵ�s�	����H��1�nD�9��޵`w��gS��}�!�߳ #��=D�*`�r�n���ﻯ����`{�{0�zՠ=�ޒG*���.U�%�0�O���a���q`}��)k��R#*��R�v���۽j��woO	���@�$P�1���'s~/�j ����Nf��Z�7���ՙ������\�$~�*���~/�"�N���#<�h��,�[��]{V��z��� ��oJ�bQ�ۉ)@�$$����<!�I��Z���:����jM�r*��r'"�o,�����3�{3��w]�w������D܈��&��v��`��,Ӷ`��,�S�� ��j@�q���n��d��o��}[���wf�ӥS�Rm�TN9�'�����>�5���{����j����� K?��,!*��H$v�mR���b��8-��RG1�磋a;]m�0��+=����p�9����k��X%��������Mt��Kpq�2YJGm�\���u�ZS��-�m�b��76�0Ѷ�����*/<w[��=Gz����fv�T\N4TT�B�U�T� 8n���bS��:8�k�E��3�.yU�����LR���n�n�\҉ҁ�e��k5oq�VѶ�)�wa�'e�������r n3m�/*&C��I"���Ul�N��8�/�`-i�ԝŇgZy� ��Kҁ��rQEd����G��b��o_����%���'ɨ�E#HrNp��ͱd�o����(�
n��?f ��9tW�f�f`������fԩ�֞`�}��Ru�{�)T�G#$P��۳� ��}���Ӽ�;� �Z��C�UT���k�Pxӻ6��6\��RI����tܱӗ9Ib6��#TK��e�����kN���,z�}��}`�L�f���M�mG9�OFfؿU��D� �^"_�: ���8����]z�g}�X	�� mө���UTԕ��'�z�gS�X}|&��`��V��Hڔap�N���\�T���M'�uTPD|l.�F������Rr!9N;{w� >��{ـvR|�;�Й
~%�T�1+u ��������N;vˊ�7`�۞�6����a���.X˄��ԃ�I�/ �u�X��e'����o0��fӢF7PT��z��=]����� �������܇UR)RJ$P�%�|�]�{�����AU
�P�O��~]�6p���-���S�mG�on�`�X^�����['s�r��n2B~nD�ʒf�S,�l���|�0'�f ���~�{���6�s]{��1��c���S�ũ���3�n�jDZhֱY�*�f����|��|�I���������Ł���#a2�8�u%7r��
u>_���4����l�3���"�?k�>m���rwwf�te��{M� ��X�㢤����	&`�K��ú���T}�8�y�����HA)�
_����������J�R6�E$p�'u���$VfN,�����Ł�z�㪩)��n�-p=�I`^e�6�֮�����sٚ����%���̔��Q�(�B[�x����o0�L���=�s ����\��Urb7P6p�'wwyς,����G�?���,�^�� �O�m��F�G i��V`�W� j[|�N��m��{�G%P8�DH��,�t�Rw=M����}��`=o�U�����(ٍ��o����I�߷��O��|l��{��I�Z s�g��mJ�7��t$�Q�g789�F�p�6`�tR��$euj��mG	g�E�s�t�[x���{Ȳh\^ݎ:wi���uvl<lQ�w����M�U�n۳��M�v�Wm�Z�f�[S�5g���%�q%�n(yr/n�C&!��D닍�����V���58�&�E;����D!y���V�k�Gnm��ZL	IŊ.˄FH��w����ww��w���w{���]�!�KpN
.Dld��$
��k{o��������Mۜ���o�E>L�)�P*����������Ł�}��6�޵`{�.@�H:U�`s�Xx�� �w��a�$(�HJ��D����>�x�z՞��ـ}�8�=����E
˗U�}��S���m��S,?�G�w��>�p��4��b(�n�lI �Nnc�u�,���u��~��rb�l;f6��H���[W��>H :�8��^��X��p�E�8��jϟ �tŒD��s�n�q舏�$=��� �����E�H�R|���?�����������,��}�s��{f��v��5���GD�R��{zՠM�����gW��܀�����ɑ���)Ԁۊ�����>�N,{{� ��Z�7�~ޕ�"�uA#�d��L��w�kN��d�r�`K�������R=�.ΎY�����t���G,Qj�k����o����sR$��� ޷x�wi<�;��`{w�$��R��E2�K�}��zՁ�n�`��ŀo��x����#�)��$I��o8I��i�����~4$π���B�?_	?}�lY'txf�M�*D�m��`휋 ���x��Յ׽��`ۭ�I?mTh�T��m� ���&�`�2�T)w�)�(��n&�)�q� Frݭ7�v�d�:m�8.��W��۱\���n����IWU˻��q`$��u�,w�� ���m��S��E�8�owF>�q+�`�����w~L�SJ�q���n���>��?�������V�f�}Ъhr7D� nJ, j��g,�y����o��@��U������f�?}�娶�1��*������,Bk��@o�����-$����FZH�p0�F�w l�:�m�ز���_U����R�#=T�5)��Cq�����zN,����=]��ջ�5**�F��0�L� OUX��,9:�}�D}'����$HM�q�)R��������?�v`oN,}��EN�,��U����,�<��Z�MՀ��:n�m��Tr;}�ْ�~�� w�e��o�����ñ�m�m�[�������EO�7F� ���J��x
?��LA2t,�¡ @���a&'DLQ	t�:���o���}��B �8�T��	Sɉi\ 0�̩���M�Lǋ�mÿL�0����3"t��-"I��a�a"$a�CB�tî���Q�=���V�ε������������0���V�$�0���m�v�  ���]ڪ��n���˲�[�$�����BAڶ�ز6u��4�D�\�׆)ݮ�FRX�&���f��,Ѧ ����Uj(�m�	�U^�6�*q��N-�X�mSV�s.nnI�GmFŷs�Q"���=3;�+��+cu�1�\X#3����s��v�M�p;5�Z�m���]���{v��-;v��ܦxT�ev�\�.ҦR�,ٳ���M�&�;�nAR6nn9�sٱ�=T�`����\�GW;!��F�N��D���a۲�=�����U�%E*�d�8�L�n[8�;mk��)Z]�e�9�A�+�i��pA���:���W��iLҵ)��[F-6ĵ�vwX��`]X�N�*��/;Q�c9�D�- �+fNɳ�g68�t��β�F;!��5V-�:�!n��P ��8¸��8)V��l�nM�[�/e݂�tb J�.��T���&v]��b`����]�#F�W��SN0K�
� �!RL��x�������.F�e���-)�E�R���*���O%J��..c�[��3P��ڎ%�뱬nGx��C(�+�@��L[��Qi`%nWA��GB�/�(=�r/S�)y�;j8Ί��WR�>��'������u���n:۷��e���әd�4� h��hzp)�C��9�/@��6�ې�u���n1Ql��s���\gR⻆"b�\���$�n$Gi j��$Z�d2�Y�Sk��T`ݩ]����񶝀�v�Z-Gl�F������c������l��]��v²��z�'"Q���ɗ��[�6ns�����ݱ���Z�6R�w�Ӹ�4�7��v��=bi��;	V:Z%�u$j�4�qf�����!=�ͷl$��@��f,,Pl1�\nr;XI�v��M��VݧA�(�85X,��kK�+-���l��8�8�Ny�	���\O]��^ �ݶו�g<�/��=����?�v�o�ݜp�>�PgY��BFD�```�?�v��!E?eO� v$����E6 -�k��@��hG� :�KCJz/¨X��K�,΀Hª-���F�	"�D�
ǩenT���+-�,q�2n��8��aq]�����c��r�o="FW�����d2mi�eڪ^p'0^�)W�h	�(��0�68�Q���Eq����T��7�@*��;���g;la�f�v�Iˮ�ȻK�����z��D�N�^Z��j����ے4q����C���Ә�gf�Y۰b�Z��L���a�S�I4�iO�@k��Qш�%���p�q���Ge1βY-rXt�h8���j;�M݃j�U�:AT��{g�`���=��_ѠW*�'s��	?o�3m��cR���,��,��j˪�wv`N�M7�4)�����eHS���%ܘ��Ł���'L������N�N����M��,?~H��ݘ��9���%�hP���+$�H���"��6�&`�8���Xj~ڰ;�f󄥌i+HOK)F'2�۠��α�<VV
I�ծ�oMC�]�gV�[�w��~ژJE:N4DI �{����eXx�7�P�TQ>���I�3w更IF�-��7s��ǚ����P���4(������B�*v�]��w�����'=�/���*�k��9���Q$�ݽ��[�XG�D -n����Sw2n��A�$U73 �t������ ���X��#���`��Dt5*P��� ���">�uR,�O0�2��^.��
�ʑ�R�H�TnIn�s,[�0�����k�z^�v+e��X�˻��5:e�թ���=�DdP�I���q#ի��M@Xm�	�X��`�2��VuR"�� k��HԨ�E�ӢI�����;����F�(<0����s��uW�߷�$������T�A��Hl�K�u`w�4�&ek��NʦXZ�T��u�n\�V۹�{_uX��}�׀{zq`�lVV}�k���S�v-�����g������J�z��[Բڝ���M�6�4	�t�P*�C�;��0oFX�U�?G�ҤX����G8L�8�+0N����@��S�{%�w���#�}>*"d�D#��/:�5*E���r%o�� ��,��%��pE$0>]ܜ'�g�_��;�����W�s|�������?}>S���͡A���I��쑵�،�p����t�6��[�:�2�߻���ߧw�x%�C:@N��r��aۈ:��-��[�v�k�s��q�������S��H�q:tS��n���>��`}�4������ߗz����0�'�*�,���#ﾀ�T�u7�N�`f�t�(��.;�R�����|X���}} ��X�����o'��W܉�P3TX���5:e�d5�V@P�a�N{�5��$�d0R��S�X����E����'��P ��%�A��$E���(f������k�����ݻ�hn�tcz9r�G�jnH�͸$��vL��kGc���U�sՑU7#�'R�`D�J:7\�;iȼ��>[-m۪�p�@p68��\����'D9f��u��PT��)�-�n ��{b���Զ�j�YkJ�'jQumS���N�V����k+�H�+NQ�'(�i�;U�1뗵�:��wggn$����e@UDh��(��1��[S\l3ٚ�D�����ƌ���l1tZ���n���JT�#��}��X��?}�}�}��t�^,i�)J���!9.`ޜX��fTsc�d��ܖEB����쑵rډ�ۅ�����=�8�?~�=���L6I�cm��I��-ݒj��Ɇ�:��uR,=�JO���sޯ��ʖ�T�PI �v�/��7v��{�ـ{�q`gު]]Hde�����I�3����rF��bԺV���;����R8�er�R���n��˪���0nM?p^,���e���cL��2��h�e���^���;��zt�(�!�{��
)��h\��g�����$���,��Ɇ�
��@���Oͦ�'�}�D��f ߫�6���3U"����0��uJ���JT�ㅇ�J����������;$�we���\�@��O.�L�Ӌ ��{��x���� ����nJp*��ip���h�`��u�ò�\燛�ݭQ���O���F�Sr!�i�����<�2�3����}`wU"��̍n��Pr�8i'8I�٦� ���;$�vi�O{��9�
�#���N�a ɌE��$��},�%�1Y�0 ꨊ�9D�2J�1�bE`�9�DQ��{� Ҫ'�����w��uy���>�ޑ�qJ��r�Uӹ0�-��v���n�a�g�^�gW'���&�EF�=���`%���� ���$��avI�k�Q_�D����<m��4\=t�v�-�.5l{s۲�ɋ�1��N�mE%3)����$��E�Iޟl�\�R�/���`UD��2LTԐMW(�z���Ħ�޴� M�." ����Ԩ7"j���`]������q�ݚl�K3nY'�������� �+�}z��[�X^���q;���,@� �`���@Pdwd�]�~���Fq"�4�R� I�.�O�G���w}���Nl���Cڰi�FL@�IP6�J%2y'�L�:Kx��ӻg j��\����EML��n��%6z�Ȉ�s� �ooH�N][Wt�շr`��V�O0N�jdW]�}�G>����:S�H�ETr������?����K�{�`|��9��Oͪ�+2�O��e�4�X��a�">�����Oٰ|��Z(EH�I�{e�~��7l�����	n�`~�l}��~�㻸�����ˣ*��e8V��8����n�և�[]by#�M��c��@.u����u��Rյ��{�=�y/f�c���]��Ҭ�:Q�Kg9�tcpɷ!J5A�cv�Y�z���T����
-����,�%�w=8�1��9-;���:rO�5]�4v��N3�x��Z�*�E��ɻE��jc:㇎� �"�B`��z�n(ܯ\q���B�@Dv��r�u!l�#rܣ�V۰Yiյ��r���NO���	��ն��f2E�E�D�����{�8�7���{��;��`e}^���(���(�[y��>��^,ڽV�H�?�{zF��J�:tT��ot��Z�*gR�X	6� ��q�U$�O&��J%H^��κ]˺��٥������N,���j'U�w!R��s ��֞`	:e�>�Vӟ"x�8�؜2n�eōN���;*Vݣc���Q@�ۊ�E���{�1˖뱊,����`�W�}���3����p�ٔ�JI�s6i���{*� � �?�:� ��O�VV׋kO3�G�2yzj=ʮ#,5%9VI��}��N��l��wf�Ӌ
����"*:u"j��uX�L��30N�a菏�F��d��X�4�-���n$����#�!?_� ���
�`8��{�3&xہ*�t��yƮ�
��ͻ^`:�;u����-�?>�x��,]t��)��'7��I�nKԏ�f���k����s�UI1R��%MQ`Z�>� ;��`R��z�L�11tmFaw.J�m����U������T�k ��;��ZD��N���(W�@�9���x�� �_ڑ!2J�I24d�#^y��k.N	0L&$gJ����xc���#�`�<�k:k���f�������Y�w*�����N�2��םgY�Ҕ�n�75QR�A!�ǥu��F`���G
ZP��4��j :�(�Z��D�S%r.�m_Y����迫���/��[Հ���{����3ێ|�\ra��h6hѣF��#�@� ' ?Be��*�;��؟̧�UM=l_E5ا��{��G�ˉi�c'~�" ���;^Ֆժ�]�O#E�YnJCq/�U����y��}�^,��V�H���v��xri�l�2�Q��;zq`�����l������>�(uGRH�MF��A�H�3hs��b�ӛ/I�q���X�ݯWS׍����2LT�Lʪ,ّ���i�,�y� ��ŀg�WD�t�D�\�� Ӧ_���&F������`�>�����:��m�������;zqc�;�e��l���]�*U�)�$�V`�e�6�r�T�ѿ}�X�d���`H�;p`������+��o��@"���B�n�
IZ0��g&F�2���݅_�=��p)H9r^{nf��<�;ncl�@���j�����
���t�u��������@��^,�y�u�tXL�iU����t���ېU!`n�vb��q`�V�i�R��Q1�8I�Us0��ŀkm� �S,�y�N{T�ԁ4��NAd�T���`-T�/7���w��Sqࣕ�%I"i�&��m�wf�oZꫜ���W���?�tD���P��EU�RQT���FC�Q]�k�۾x�����1Ȝ����vm�k�<�cu �ɨ�Z6�d#�]e7i��.z�m�>�V^���VZX���]��.��tA<��28՘؄����{4�����"r�]I�渮�*s�6�n�N�,v˶��+qu�qjʝ���mΎ
)XvaA���VU�8t��]z�+Lӗ�<�˜&d��|)k���s<�p�4�7��w�n��~/��p�قR�b@�w@�Vr�E�4c^b�JSdJ&��봹m���;�~�����iW�$�Z��)�z�R$"��qStS��}�֯�T�e��4�7{�7����(�@������E�6�XݤY��""e{��`?��Ձ���5"˫�r:�m��7�p��`)���XLδ������"k�IȞU5E����Zw�)`{�M,=^��i��U4Ȩq��:{$!�:�!i{T՝q���:��ȶ��u��^���$FJt��s0�zՀ{��`}�L?�N���s���}mG�"�5��Uy�>����OЄ�ǊFsI�?������~,�<�:Ӹ�15)�p��U�;��g��� ���X�vX�^���ڈ����Ͼ�"#���w �?\X�����"���ґ!(�I6�s0�zՁ��}�J�u�-T�|�����c�gƋ����'Y��lv91u��k�ͣ`{xZd{=x�;�%�%�"�Ī�q�QV ��ڰ7�H�5�� �N��Ɠ��W �����J�r���f��i�֝���{�t�Teo�5���j��*��m�֝�����HQ�ع�.��`-�����-��#%:UQ��ݽj��w]XԮK��O}�{�^��z�T�fNMD�ʠ��u`z�f�{���q֬Z.U��UHS�O�B�͠�O:$W����f����:����s �,��n�r����QVKw0��,����ݱ��"Nf}/�6~ǭ����)�l�(�7u��2kwq`�����"��W?|3_�8�e�$	����'=�X�An���;�H�16� m�q���e�4J#��Po������owf�~�*��%N J#��䄘b���F!C��Y@b&8(�QJ �� �&���R�(�-y￮���<�~~�pj3.���%��0�ޫ7������I��e�����(zF��lcO��:o�~��o����h��%�����C���;<(����2�L!$(��'߿~��z۸�.w�� K�M��� �
�W��r� �n���w���K�M���� $sN�i��Dؘ�1g�g ]�(KVVH6�ŀc�#
*���8���w0׽Vwof�wZ�}���{\�ʕ%5�)ʰ3�<�/�����Ձ��6�G�� @AK*q��h�\�k[ֳ{��Vw<�.�N��v�Z��J��=��q��M�-p]�0�n��N���ۣn����6m��6S\ Y���7(i�&AT���B�c����cDm��.��̆W&Nص�ٔ��yz^X;��۲��;��A��E�<��uU�NU9Bk����]E��l�cC�N�YΝ�g�Y�Kv �E���,���o]�k���;j��۷Bܡ��6�m�Xq�H¼�W\���T�{\�=��H%n4��ʐH`�;�O��b�&7y�w$:ݼ�!7\�&� �h���X�F�۫�Fwwf �}���{�} �0������$��L��o0��,7uՁ����EN��*5U!`gwv`v�� �����ޚX��~�O� H
�73��,w]Y�橰1�� ��B7���T��s�AP�vr��� [�l5u��{�uw�s�R���$m�yU ��w�-�s`bm�2C�;����r
p$%H��ws2��=�߶>�";�q�F����sf �w����W�Er��Q�NU���ـ�m�?���ϥ�s�5Y'��[r3?H�T�)��>��V������Vwof ~ӻ��tD�Ӎ�⺪{�S`ci�֝Ł菾���������Ë��7�d�ur�v��3�&ln5�Z�q��hٍ��./972��w��9SE�UWH��66�`i�M���`z�]=%�R��QʰG��يd����7�U\������A� c&B���p�{����O��/V
|� Ȧ6��(J"QP��9��VI�s��	9�	m�"�D����?UT���t�;9������Ł�j)"un&�K��o�q`gv�`v�� �ݲ�ůղ���u�#�#� ��9b^e,����֞L<�n�Vz�^(M�,v#�G)��MDF��h��� ���X��,}饁ܻ�9����E����'���_�@ �'}��$��4�'��o9�
����}L)L���c�`W����"˙���0I�X/k�Ww*��#��u$� ��q`g������yΎ��[(!�P�S��h  1C��{e�|������d����X�����X�����zv��q$�R	���0�9�r���n�$튷�=�R���z�0���U�T�#DG3 ��֬~�K��7���Ȯ��R�N��7"��z�X�5K��O0�w��0N@un&�K��U���X���}_�77�g;y�_	;�w\B(�62O*n�D�~�w ��q`��ς3��x]�:�����mU9����X+�� ��T��y��#ￚA�9�Γ��%�JH�� �_��H��$�b��$��j����!�����X����o�ݔ�.U����D(B�� λ ��`��>H�� h���8Nz�DŶ�l�OV�^O[Q:Q���^� �"$���aꔤh�	�����ĉ(��`�k�� =��D�������-FIZp�ƾ�Z��
�#Fڱ0Ľ��l�}��i]�1�E>�0�w�4k;�f�h�V$vY�E%ҏW���4�6�gm�+T@��UUn�4��-6KҀ ��=�jT�ӡC�SgP�-��W�:�-��rZV`tEq��ۚj��
B�=���[��;4�dقMЭRN%��P
�c���vŚ8�����뇵����e�V	��u������l�����n��i$3^\ݰ�r�v��n}�d�`*\GI��6�ˇ��VH[�"����&��F�ˮ�j��[]��7bț@]J�Z�w"�S�f�r\q2q]8�����u�p���2��ō�q���{&�q�t�s�y��'����H��x`�(��m���!��NumF�jh��졊Uj��k�cEU�@a�r9*����+g��d&7n�ˤ�y�t��و]m*܇a]U��,����iK����[J�v]���m�-Ȫ4�Zt�6���C�����k�@�MUU�@�{{�kX ��C4��*�>��b1�#<���UY'y��Kk��=��i3���SF�c@$v���bD�,�B�ř�HUKթGmҦԝpU����Q:[vc:�2����*��K����ճ��o�"m�����Ǟ��1��:����`�vҳ�56E���t��u�ˆ�v��˽�V�y�8cZ캍���vj}�9�Ž�	�v|GC�ulU\ruĮ�h�,�ɧb��g��;��!-�zۜ���%/��n���۞vnS&X���PRk�H��36DZI�(V�0�n&�:)I�=�~~w߁�km��V�X��{!ė�gme+C"�5Ll��v/P�&�GBӮ�dM&�7Z�h)z����h-��E����X^��B�:3������m��Vջ
i�V^t�[lv�� spv�%�`�r���M:�im�
�4��!
ĻW���KhY�,�Ի�qٲu�у=1��u�۳�(W�+��)�gnV��bv�J}�IN!��8��#@뭌qN9(P�\�Zi��RC.�EU �P�b�p
� )���qtҪ%��j��_C�N�Mv���
�)p�rH��Q%-�+�v�����RV�m)ُk�CI��)���][$p�<���}��d���5cI8'Y�Ln��e	J� 5GQ�Ku~�����۶�Qu;;��S�\6��Jm�\��m�5\�A��!ݭn;�X�ە�99�h�-\�zc]9Qoq:�h��7=��Vg&ˮݯ�o���f,f���<a玝R��74t�R�uʁ��s������>�>�A����n�ynV4���\�U�&�OUm\�'vΣfZ�&�j�M��D��_�gn�`,��j����Z�����$�3_�r;D˒96�Ua��s`bi��n���H��XV�:{*��IM���U�3�{0�����}��"��7x���� �GH��f���X��_|�����هUv�U�T��� MȬ~�U���"7i9�:���u���}�|���R�$Dr��q(�J�e��Zڑ��/7W�Zջ^�m]�!��ܶKij9����	q�lM��;��{$���s��R$�mE�X��ٜP���To��tuW���請��j��]���EM��3 ��֬n��I7yJlm��&�9<�cU"%JqX��_S�Ձ��{���۶,�h�n�j;A��9�eU`�NlG��{��@�^�Ņ�����^�@���5J�lL��Rm���3Ү���]�y��
, �7����v6õO9�*lM<�;��X@.�}�d�������W"@S$t���`��s��̂�u`w��\�O0�iA.��Ӣ�� �Ԋ�7�tV�?mYiP�yU ����Ȧ��Os6Œy����$jہ�Iw8OfM�{��o�f`{�Շ�U]��,篜�(�:�⣜�yS`b�y�2w[���E�Ձ���d���4Ɨ%��L�Q&)��2���n�VG\O�����:�m&gv��w&l1���6����wZ�����_W�_�A���`��E#��i�R"T��u�����W���ـjn��3R��� v���)K$� ^��Voog�I`߾�d�7���OV4��%��PU6/'�jN��uՅP
� 
�vL�d���f":�UG3 ��Z���/�Q�������7���P��R5M�t�n�O8�=���[�=���<��Bn��3љЩEQ&�V�{��>�ݫ7�� ��Z�3ݫ��%T��Iw0��, ���Sw ����D|H�����(�b�r;$�~߹�O�v�t��_?n�x��9EFD��ܙ��c{݊�3�t�>�n������hW���2cID�%��'{��Υ�O0M�XA�7H~w?�;�&^X��kk�*�X�� b0���%8x`SBitc�A��A�.K�?��>�n�gA�H��n6^����K���@�صIy�&%�p'M���۔��\��C��v�8��֪[���vV}��r�������m�����ڪ��Al �� ��]��H�c��y�p���1��7�Z��z1�KH��D(\e�C��� Uw<�~�F8�N��P8۹�'�X�p�*\�s�=�*��v;�5������m}���*�����a��t� ��ŀ.�՞i�Q�MH��vH<���G��ŀ-�V@vu._�Cwރ���31¹�	*�0�� [��Υ�1wv`��(�)T
R� ��^U�uX�5M����u��;�S �TA�qE�]��{�`f�v`{�Մ���d�����j�"QR'��"�5���R��EO#�F��F5�"� խ'��$H� 1��\$�~��q��}�j�7�t��3���rގJQTdZٚљ���^{�tu�CU
t �  �C�����s��d����y����wD頍�"�Q��~�K�橳�'_��vAsދ� ū���j��n�)d�a��ޫf�v`{�Œ��{e�z��`0J)��VCo0�w uՁ��T�ݒQ�;M����ې鎜�
��9��Ga��ue��vճ���h�b�v�8:�lMUf�n��1l��;�j�o0�FUt4R�P	��o���_|��`f�v`{��e���#Tہ�Iw8I��j�O3wy�
��WlUP(��ذI<��d�ƽ����U(����7�� ��֬}�	=��+��761"�6�q6rb�Hjwq`R��橰1CO0��{TsqpK���͵p�zwn-7k�Wf����.�+fG�׍ӭ�GLU�����n�K��g�u�b����o8I��֬=�|��]�r��I=�o��L�m݁�n��;��'{��*�ƪ5Qʰ3w�0��j�=��X����t)�U*�"eTnf���y -�V{�S`��܈�|:�y��Eъ�i��r+ �ݲ��y�l��`��,��A�N����i�.�1pi��8�v.9:�S�Yɳ�g�̆x��*�A��v�-ԧn(�Is�7x��m<}��N��}}��:��r�'QA��n�r���{0A���XJ^�p�.��VIݭ͌)�(	�'��Zw��V@oy�lm<�9�v�p��IG��Y��Y'<��������޵h}�k�Cn\���*ʪ������o0�w��I��^F�E��q���Gi�ӵk��n�n*y@eL�h!f�̅�h[Œ��`�+ax�s��&ܽ�����'.�]_��}�әǜ-mq��(�W��U*JsѢ�cm[;�]pmS�hʹ��zefe��E�b(șW����\e��c�6[��i�f�R��Ug�r��dX�m�3����j鳵j5Z�N�w\Y�7h��l����4r=��������+�����ݒo�����3�ky�[���I-�gg�i	���ʨ78��@Tqa'g߹�O}�b�'���⸉��j�O���8[�0���J���Ϊw����y�lm��DPH�}�@�-�mK��s'���ڕ68��o�~�S�ńv:��R��)E�]��=�3�{3*���Հo�e��k�݊6�qB8��nM����[w%�.�{�Spg���6c8�7 d����8�	�pu#��Խ��՞ܕ\���e:z�丫s)sp�&yY�w[���u`gy&���	M<��]�6U7�Q�QR+ ߽�� )�*{{��v�����8I��ؿ�
	�k��MN\�Ȓ̒p����`gS����ŀ.�Veo%\&g�Q<�T���zu���@j��, ^���mt��MH!���;�eku�-�s`u4� �}�ls{�o��p����V,p`(8A�gV����ۆ����]6��:I�m8��Ln	����:�#w�������;���Q�yps�rJN7X乀{�z�֛���\Xw]X
T쪉����$�*�X�ݟ}K���ڲ���ߛ%�JH����G���6
F��Ej�.��d�GZ��<;`4�M��n��
�s��dVjQ�c���A:��0�ę�L,�0,31��fl��캪��U��0�v;������)t,�DX����d�8�`XI��c�ӄ&F�aJnքi�<�Z�I�.�7����+�2Ȱ0ֻ�<��j�lCBm:D �:=:�0���+��*zBx������PЖyE��u����,|����^�ʤ�GU��EI�u;� �� 3��64� %]т�o�D�8��{���i���;���K�8M|��,y4���Гu��q���D����N)Ǝѻk�:�rncmƣ�R�u%X��NL��X�ݘݽl���k�l5DEO�PMr��ƛ��ɾ~��K�`oy�^�[>�|ѷ�!���	>�~�p��V����]O�-���8���`ԩ@*r+ �n��?m\�F{�����C�`t��	�����s���y�ϗ�3��u)��H�� �=�?�����w�o��, 1k��ԉ9\���U�r�P�.sۭ����b������n�+��^���s�"s���W\l�����4� �q`�Ձ��T�@�5�G((�P8a'9�Ow6��TD�s�d���VI���>H����'a'HFQr��#�z�ٝ�R�G�L�y�0^�Ł��|�jP��Gb��I0{zՁ݆�a�n���Ů��7�U�L�D�QN+=�ـ}��V���{�GUiH$	��>�����Te��y#n����b�fU���^٫,�h��A]��k�ls=��z�ۤ3��,�6�r�Fk������SM��\�-��W4�v�G6�������-s��Ͱ�8D��w��9Zj��nf�7Y:n�7Kx��"^����ntt�T���:�)�6�X���m���>��cOvf�y�q������h�#)������ǉ��n
��Wl�فv����˱�i�l�U�%ñt�0���7-�j���7����O��]X��q`f�� �#��*~�I"��o�X{�j��v�`n�� ���gT��	R&�˹���-̝T�`I�X-qVQ�H6��A%H,��Aw�߻�O��Z �{���������*����O�3��:۸��K�wU���y���S�B'�2�q7 �Dr�Q��rm���f+�kO!�T�U�ڟ^N��+�FQ8�O=�I�}�,����}UUB��������5��b".�GdIq98I�l_�z�U�겨�Y��{�O�6ŒO}��H�^7��!fHb[�a|���5'q`�u`f�q`u�TtB$�J�R���U��ح y/U���Ł�M� �qtMr���S_L�TXu��25+��7�@jNՁ��w�!��!�d���~����&휒j�]�*��ۗI�؏�$�#rN�IBS��r\�>��Vݽـ{w�X�����I�kT"�(�TqXv�fz>���7� ��5+�}�������R���E9��Z��l���"�"���<���;�~{�`w��ـw5�Q�E6:R!�n.�=[�T�۫?z����`۸�=��ӍUe]��R\�&7{�_�=᧘��,��?}/�g"Gʪ�����܅�#�gr�R�����ݸW�`(�Q��Z۲�tV�:S�3��o����`	�qW uF���KUŁ�\H�pD�$	f9�}��/�D�n}V@�M�X�O3�G�$y�p�+�L�:�H��q�,{vպn���ـ{��X�\
�I*7X���K�~��싀:���`۸�F�>"H�q3hR�  �U���I���i�EO"�bk�ko0m�XV��7VX�O=GV�8�q�$aD�bg'm����Ѷ�9�}��8:�m.m��/���E��Q8��U&,��j�~~���ou�=�ـ�_EqU:uJDJ��`ծ��Wko0����. ��q��j�7b��&��`g��0�����o�X�I��l�OfF�R�c�������R������ �j�=E{{�Z������ uHu$����-̞��U�Xjo#�7�=�"�~T\TpT�#����{�gq���fڀ�ZW,㫸�ƈk2�u��\�:gǻ�(N�8�s��v
�
M��
1�Ef���튲�k�/��فD���Ar�Me^�㮍��Z�;�֮����3
�׵��U������Kٗp9�|�V�{�qu�1Ys��`�	!	
�Ce��ӗ�f�{�)mųt���^��g�lX95�.4=��\b��7w����O��5�Ͳ���d���$p|��;ʋ���sA�v.5Xo(0�k�L��L�UUB �w�`F�W���Tq���Y'�f��e�[���c��u�F�7!~��"dK��`	�����6*t�UGT�$V��ـjn��:ګ��ŀ�uUTψ�Tڪ�0�޵`���{vՁ�wv`{�D�9��N�H�R�V:ګ5+�7[y�jN��P������ю1��Y(� ��3I�7�:�Bij���k���\fA�q�����{㟾���5X@u7q`n�� ԝ��8���Ş<
C�7��}����C�`�8��m�$���K$�w2��(RG�~�T�P��L�r�� I���:��}�j���ݘn��p�*)8�j�, ;���7[��:�y����,V�W�Q���n(��.`�֬��m���� �j�}}|��J��X60�a��e��K��49eJ�[.�Ll�#�y�`W4nv.]3��5v���[�q`A֕dd��*�&g���H�
���URf��P7}����V���0�sUWQRmR�Y���gU^s�o����:�C�R%R����L�y���;�G�s���}�ގ��K��R��*���֬֞`��Xz&{�:�K\�>���&
�������y�G������0�}���̱d�bX���H��J�2`�'�\JJ�j%݂�9֒�:,��N��ENj)Q@
uHu��޵b;�Yٞ�+��	֞`)rr椨�TL�,Uk��ݵq`n��2wV�_�>��G�ZqDÂ7.p����u��vgx�ŀcj����pNF�qELrE`{ݽ���j�3�e�� p"��T�V��b�?w>�8d����M��3 �wZ���`{۶��v�`H��$����8��N@�lvtl>�pmOn8�:��]�V̏&��յ����6��(ER�8�;�+�ݵ`}����sﾱd��ھ��
��R!W\�V �w�CSyx��,U`f���Q�ڨ�C�qX{�� hnn, 15Vf�q`cM�T�S0UJ��fz���`����{u�{�� ���v�UUH�R$�XomX:�,�O0.vy�����t���fVfVk{���E�]�� ��Q�̢��BfM�RS֌%���Պ�L�1t=2���Ę"�#*L����4b:�4h�
xO�3@^�8���A�4XD�a�3���EBk��<B5&�f��k t� ҫ�(��&�6C��Jh�;�M��IDH413��)�c���&v�К���%��''Q����l`d� �0��޷�K~��$�3��ـ�u)�{��'��#�Ĩ��,��z���</o��wk���ߒ��>\�l�K��[+mUU%ġ ʵ��n,���� %fC9�h *���u��g��k`�)�ve�ŕVz�p���Vڭ�!�y�I	��&j���̪Ծ�iV����"�Iv4�H��Ҝc�-WA׀[�Xg37)�6���� ����F��0N�Xn@.�i��׵H�]$�N�yܲ����^� M)t6�����t�Ѯz�ũ�')��v ȝj璌�k�P6[=l�xn�r��畗��ݶ���-N2�l�c���.��F���G�Ɛ�M���3g����L��m�2Z=t���`��âv�\��ƣ�	P9;-T�kV�e!��\�q�wrm��MUP [��q��Sn{u�>�6��vE������7Q>Qe���4*�,n� f�L�@#t�dU�1�S�G]��ڻU�q��A�;-۷mG;��2(4I��Z��]��L���c�U���:�p�?_v�U7��L�Ud�d�K-���	I�5qcv�d�� H���@��1�b8�q�٧�g�m�v	�Jl,֕�\t�N�Mvѹ8�@Bij)V�9�Y�vK��;�9aAH]]���΍����s�ͥ���\��U�8�n���ܡv�B��k��]6�s�/;�9��*�<�}��9�Z�%�}v���^i�`DU�Uڶ�1���sHGlN;3�v�mJ�b �A&��P�ck��)Z���9Y������Tۛ!H�*�RF�MSIYU��nʚ�^˱J�	P��eR�D�f�f l��Z�dnS�PU��c��YUjj�v����تTb��v�v˙tv���ۯ�����튃9�*v�S������\D�����N��F��
(�)ٷ`�/Y�l6�Z�i��M٣,₱��`]l�*πɟZ��tk,{1�[9���4��SH�`M�Lڋ5���:���)ӷ�2�jՊ-�B�lexٟd�i��v3��FE4�n5FO�_@UP� �t� �)�:�O�N � W`tt29���jمq�\�8���?��lFɊ֒є�5 �nD�Zx\V�R;�+b��m�1�����݋i��7=͗td��c�.٧�S�lai|ͩ�m�=�i�Blvtp ��.���inP�یF�i���Ԧ�g����9�������W�s�ᱣ�Gf[&rpXj�HB�@�Ն틎D�L[�s� �z;tU&�L�0]�8���}ﶻ��+,e�u˶e�tͳ��BXBK8���n�	��a
m�0��0�ԐF�
�H���'�k�I<�57q`��a�������&�rI`���ه����Xol���f;�?g�}��R�	�S��'7޸�MW.}Ӝ�O9`-��`[�:��7B�Q��7�XW�]�J���׀ooZ��oI"uW�t�)u�U`)�Xi<�57q`�TXa�eY0ȣp	1?!,�O��S���ɴ[���:��m�紂78:�͕K5��%ʙ�U8��f@���֪���t�g˷�B'(ET�@)�����H'�"�"�uY���U{���,��no9���ۿ5b8)�A���_�Vw�M��i���� ���Ќ�m��.`J���G���p��ݱd� ���l�Ni;a0���*'�&�l��S�X@bj��+$��N�A�HƂE(1�>�7R�U�<�5��L�]�MnWmu��S��m8�􊛢��˺q`������| ���}�s����v�-�A��UTX��U~�>���	����<���٦��T�4+�f�����v�B\nNw_�+$�s7�=�D�]�B���@{W��,�s��Y'�1��8�P���M�֓�d�g[������fwx����)#hu*P9���Ձ��DE�Σ�b�s`w�<��7ɮF;p�j�k�{����-2�����v�k� ]y��t�h��N�Z^8)���MU��Ħ�;�;�5�q`b�`ʚ�2H��0��V����5�Z���,�6&�:{�n(����֞`���MU��K���r��N�)�p��B�o�pY$�~�d���+I*C�P��w�so���͊���(�*7�f���=ڿU}����Ձݽ��JMҡU8����S�����%:�E�1u�VB�v���K��u�.GK�dwRR��U{guXv�f��`��`{��ʨ�$��+�ʪ� �I�zdO޸��:�;�[VoWQ��:�(���j�1�U��9�����7��P�G#��HrE`��`}�V��ݽ�������G�Cr8�����F�;�<�5�q`��c�}G�L���
��#cun*�Ue�]ˋm�=�������\-�"s�ժ�Ь<x����b����kv�X�v�M������\�X�y�JfۂGt��311SÝ�� ���K���v�d����I�"GR�n�z��d�Gq�6z�vcZy�������F���r��Q����K����۩���u�5=�ծ��s���^-��A�1#���(1���
� (K�R&�p��]ݔ�O�Y�.{4�*OD=�t�v���ݚ��}}۷޹�v��T�D���m:��of��`]f��u�j��w>p��~qSt��[w�ﾙ�ά����O9�H�C�����i!1(�I�|����Sd���<�5�q`g[u<���d�)K�ɂ2�guX�w� ^��b���Iw>�d�Ǻ�1@T��"����;I�rd��ŀwZ� 7x��M�����܈��E��8M!Q��v�9z�V���t�W[N^�θ< \ꋴ��-H�D�{�n�Z�A�;e��=ڰ>����Uu���E2S)H��e�P��
���d^=�|$��w�$�7mZf�rGR��qEX9s ���;�<���s��� ��Vj_r	��*����v������j�3{b�>�n����¡)���T��`��,DG�~u�l��`w��������۵�v$n�jtv6���+�{k,�`���Nƀ��V�pL���չD�⦹ʋ�����r��I���~�� �����U��EӶ����=[����`���3Z��7�K�QPL�m�r)�%홼$��;UB�D  ����P >)��,�ՙ��&v�r#�A����f�^��V�Su����j������<*I�mR$�X���W�]�>�of٫lY'�wV�%ƣp	�
9	F�щ�<7G;l8S1�;!ۗ��I�M<�m��ӽ�N'$n(�S��k��v�`��B�����4�'4�������S*�`�'yﾉ�?z��S,W��O@�2�`ʐ&�Ns��M�X��`w�K�`u�O0�r��8b����ni}Ts��Oq��Uy������Wԅ� i7���g@{��Uݰ�m��t�XoG�f����w�jn���j��Μ�y0�+ch�ۡX9^����Z��aE �`:�^��^8kn02u[��Z*)�m�i<�SwkWgR偍9es���PH�`��V�vڰ>�n;$�ۛ�|)"~�O���Q�HrH�:��,Υʸ���kw/.]
�F�QR�1`[�����d���,=G�Gӯ�"����K
�hr;�Py�w^��`}���/f;$�U�^&�wT:�g�ѐ�V�T�U��kv�f0��72=��2h7��O�r�����q;n��l�5�/a1X;KQS/;�:��e:.Z���
���p�x4�l��k[��C��nȨ�v������p%�R��ɀ;�67B��Ƴ�x���k�;U���V�e��Ikw@K�<�$̬�]-A�탘 ʲ�Yi.���-��iD�n��)J}�ݶ��:~��$��1Y)�E!��V{ V�Gv6�ʡ�n2{rW�����:�A����[qH�Q�)��D)>�'�g�,{���W�]��ov, 㷢�ER��JR%TqX]}��V [[�vݽـ{��X#��wH:�M4KA��X�o�ZO0M�X��`ox�rb�%
G$�RJ��#����=�֬�M,A�{u�����UF1��$��jn�ə�G�gR��m���p�:]#ِ[���m!ƥ�F� c��;k,r� nm���7�p�4ݮƫD�ʪ� ֪(��yas֖0�\Xw�p.������&,ս���*�T0
� �����6�{vłO��b�ձ2��OэF�#�>�wf��`}����ۮ��r9�8�Q�?9�I5Y�jn�ʙ�j����\���ӫ��������$�Dl�U%6�3y\Y�Թ�=��v�M�X�@�k�/9�Ю�p�H3*uH	-����v�U��M�p��tqM_k��>rt�.0��,�O0M�\�¸�7�ڐ"�Hە �v����=��f�ڰ��]���K�6J�R���f���w������V\�rbs2�[���ί��BB�r,0���b  �H�!H'!��D$?q] �����)���,ݧN/�d	�E*af���Q-
�B���j7hΐ;&&d%�;�kIL!�IE:�((Ӛ�JJJ
i$fQ��>�>v���Y���>���2ϣ�9�$L�P����v�vL�!Bd��c�D�zSl0K2,�R�ERT���	b�����c)6xPa?.��M�g���S���f����*�v��ԭ�d3���
I�2R�2Z��%z�)٥�2$&L����;�L�	� 0$:CA��__��2�DCE%%!@R4*n@�u�{�����a�dᓙAFl���T��MJ�4��I�(� �u�j�2̰3�,�Lֲ����E���)�AM4��EѤL��ZB����RR�Bj���{*�n�H�:gZX�L�8��@d�D(L��DG��w���)�/~���v��=N�Оx�+�b/b� <�P�;��h�]��)�i�Y���U���v`��䐈�H*�$���DO_���BW���� �G�����������Fۊ*�˘ �|���� ����&��d;���qr��ū�]�8�	�n����󖰆�inѵƹн������^��K�G�q�i���� ��z>�#$�s`_|�R3a�p$�N_-#�ݱdG{���%6u��=2<��T��y�*����E�uyՁ�Ħ��|�`�Z�����[��ult��$�7_vuW���w�^�����G"a6a�u����T$�,Ȇ�^�7�Ph�I�a$D@A�U@j��	�kbA%��NW&���<�#Sw�j����\�o�w_���_�ڕR�����+�s�<��x�w\p�Zt�nћg�[�v�eW�`�N@UEMWz~�ŀgZ���s��q�Ͼ�	?n��!H�T��'u~��>�艒6S�Y$����:�Ȱ3up*�RH6⊖\��{��ԓ�`��� ��X�Trd�_W�\��j��=����	���Ձ���v{���!#�JP��m��7��U��Ր��l�[�>����#�]��o�b���!%���kUe�ػe�+r�)�[7(�3zU�{U#/M��l��gu��Z's�/�n�	
6I��^�L\�Vm�*N䛜�GQ&v�s�	�����6�ͩv��+��6�a3�G�ʨ�S<a��Ǿ���c�OJ�	�Ͷ�[P��S`UP�u��%m���-/zyQۛ����[s���0�Y����cn��]!>������U
���<.ZI bpDS0q�Q�6�c2��犻p�
�g��7:�V�*l�O�ґ�qx�����{�`}���0ou�f��q�x���`\nl ;�n�M�Xku�艑o�$"S�Ƥ�Ed�{>�� �{6X�U��`{�Vv�tm�TT0�B��f���MՁ�Թaw[��;v'ΣT�r
I�+7�`Z�, ��q���,ߴ:$��	��rj �у`�l���x������G5p��N�����RERFۊ*�˘�[���[�[w ۫�RB��@�e6�l�#�O}��s�Uh �"��>��芢;������Թ`=m�D⑴�M����wZ���e%���d��ۼ�$������HHJ�Qa{�w�Հ�5M���y���,f��ΜE����C%�$�7_uXA��y�kn��3[���6�g*h�q.n��p	����6�trv�V�R{l�)�RI�봎[���⊒�m�3������s���0��ŀf�Vn�)�1�.�<����R�'Rf=�֬���n�mZ}����bo��UUS��
I�I�nK$��1Y��t����"�UK_�W����wu�7ˁt�����'�u�B\nl �� ��ŀbj�*�=Q=�TS�mTQ�`}۽��8~�F@W�X�%7 o�7S5Dу�Ͷ�̳����s��6#�D�u�㒘�]j�v�2�k��]��>|���ŀbM���7�7�<���r���H�Q��=���n�>���w�Ձ�w>t�YQ��C%�UXl��`wu���W��MՁ�kn($N��#��y�f���꫿y��] '�H�@��u�k����GN�&0�B��n�Z���#���޴� �G�D;������ޛ�Q��ґU����j+DV�Jn�4:���U�y5�0=�aPz��S�5U���� ���,�|��Dv$��V���?�T����(�r������ۼ|D�n��������*�H׽�.	DS�mTT�`{������wZ��t��f�{��$��b��D�>O+0=��dXW�Q`n�Ar�� �ݼӐ�t�
(ʪ�k ���T��i� ���X��\}�h��7v����c�,��+<�W;Tvù��:�tJ��^�\XZ�v-�iv(��\�TI��z���>�tY-n=�������v���Jf���e���4���Kx"y��N����,l��5� ��GfG�q�-�-qs�wC#/23
��=\�n�Wv��%��t�p�^	�ML��rZ�V�ٞ�m�y�`mK���N8�Qy�c_ێ�����̜2��$)��F����˗�����b����q�F�����g��v�YPZ62�i��'�d���w���`���٩�p)�\�����u��n��3[��:����\��t∠qr�j��V�>�t�*���Ձ�ݽ��عIM�MF�!���<�첒Y��{���w�Ղ3��)T�n8�N\X�o�w[�&�/	Su`���_��=L�쵊(�8�k<9�`�F�un�0j�f�9�#�d�Kz;W9"�<mל�j� �'��57qp3�j����l�wI	%T��M�nf��|��v�"mN)u]{���Wk߳�>�ofQ�ou4�(���"F��u`wx���O0m�X���~ʖU+C.�,u�U�����X��Հ���`}��q�2��S�������i�۸��ηV�XOb"��5��CR�Rrp۫b�#s��Uk�ە��mһAO,��N�����
��[w�n�� w��`n��8��ԡ
9�g���5*E���y�&���L�jd��+�28"6���N�f�H��w�,P�T�(U5L�P�H�(�@W�Pf�ؖ�<��	�%`h�?ThQԧ�ݘ�u� �wKٓ�k}��F��R��i���	#wŁ��n�N�`u����}�����3���b���@�l d�(Y�������*\9-��=h�#��݀^u`WuZ0 �jxd�jn��3�ϣe�
YM�$��$�=�8��=�{0A��-Xolܠ�s\r8�$C�ӒJ�>���{{�Y���,���X�]ߥ"B��U�I� �wZ꫿9����u���u���&$`h�(H���R�f��'=�hB(�:�!G"���X�ݫ�{0wu�gwu(�J��GD#�ӕgu;���u����Es��)R�mzu�ܡ�/[R�ER)$�e9s �}�`}��ŀ{wl|
�$��l�O��SԠ��F������3�'��q`�:�U"�����G	��dM��ŀv�Z��YVD��j�,�Z}��GvT��}T�$��Oª�����I�l�d���o8I�ɦ�K���	��զ�.+�J�)�`��%�n��<P_R�����?�QU�� �
������1@��e�u��;(Ie�
DJiQh��\%�E(
R�B
�JҀ� �%(� %"�AH!B R�
R��"RR* 	J�@ � �H� ��!B�҂ (  �P L��J+J 22 ��44�*�B�@�H-
�@�
9#�����-
-�*M( � �$ J(4���P�P�B1 �B��$H��� -*!H"� �#M ��(�J�P(
R*�"�"�� 4�H�Р�B% ��u��Wr#��H*�4��@�J	H� � �@�@	@���GP�
$�
4��  �B�4�T��1� �H%	H4��@�B#�P�@�ģ@�"2)J�Т�H� (�"Ћ� �@��P	J��-"#MIJ-*�#",@�Х�"ШЃ@�(P�D *"� �(4�RЪR�B�- �؂�dϳc���h
��(� Q��}����|�l����b"� �}�_���?䊒�����*���*�?_���?������ �� ��O������@Q���������o�U{�d��?������U����P JPDT�������!��?���(������������# 7���*���_���������?�������?�����k��'�P�����������E eD�RIQA$AF�D�D�IJJD �Q$!D�HTH RHeD�%D��aD�Q�THQ T	Q Q! !D�HTIJHaD�TJTIaD�%D�aD��RTHRI IQ%HU!D�TH@HEIQ%@!D�H �@��$D�&TIP �Q)Q!�RQ%!D�
BQ$%@��X	��		P��$%U�� !%DHQIP��Q��X��		BBF ��		Q��$ 	Xd  $$%dFT��	 ��Y	 d!��  %		BB@���$!I��T %		B "B��� Y	I	��BE$! 	��" ���� ���I	PBBA�!E! @��d! 	�b@�
P��
A�	��d%�$��T�$T`%� XHR@���@����  %%	HH  B !	%���
%	d���EhDh	@��"@�IF�  F@�YBE P�%BQ�$B@��!a	I�$IQ!	E!I�$Y��@�dD!	� B�$d	HB ��%	@��%�! 	a	a$�
Q)B$	� �$�$!BQ�!� �P3�������
��~����9���C�����pTQU���sZ����?���?��:����k�����_�j(�����S��D ��_���w����B����U������EW����5׷�p����~�ѳ�����0����nU��Ο�:�&�����:EUn���?����QU�ô
~�~�: �G��qQU��QU��P�����������#?�������E��������������c���(������צ���4��C������������U�?����"��o����E\��������0�������d�Mf�l��f�A@��̟\�޾@� P*�H  P  (�P�) T�Q�I
 
 �^r�MH$@����JAHT�QE "�E@�TP��
�� J�**�IJ����@��'    4   @ �C�=�����csj������� ��b�6S�JOs����^:� �Ɖ�:as5p 5��^��������2�����}�o�U�y{��>�PoOZ���w��{i�,��o=�<  {� >�  $ @��}��������s:R�3e)J0�;��(͔
S)@�&�@Ӎ���@t�JQM� ���P 
F�������G4�(� z�J ޳���)Jtp�O`�=7��E(��R���1JP�U @@��GJS�|{���wo�O]����{km��l�x�^n^{����\ ����}q��ŝ� ��M�y=/^���������=K!��ũ]�� �������^���K����� |
   �( 0�k�}m���\���'�ۈ:g�A��{���v8�L�� Sz��'����/ >�����jo��t�}[�����^g���#��x z��:��{g�gN۟{�� x�     � ���c��=a�7��-���{)��^�z���z��[�{��/��
ٟv}<��P /sˣ�m��-� lsA����1޳�w�x�zn>�A�{������ˌ��=ү     OPT�ҕ*h  OB��T���C<z�T��  تT�(�j��U?�	S�T�R� �"$)��*e G�l(O�_��������K�SP��w�!D$�D/B���� ��PAO�E U�E U�U���x�D�b� �<��kF��E  ń7h�@�O��@�YR]~���FA�d����XԈ�Et@k.���aXЅ P�F!X�4!HA����lXP�<hc��(�D"nf5/��O+
��!%L�7?3i�oA.i��u�Q�Ϙo5�48�5�0�ca�(�@���~�q�P܉��.���d���(��B��j��2HK��If�EĆ���l%0�
�
���!cJ�����ů����qv�/n@��\S�Ip�CS5"!�4�jE��+�Z�(bŀA����`��I�U�vq%�n4A��,X�ac�$���0���rB�P
%"�*FHv��i�X�P����4�$e3Q�cH�1bVԮ�S	L�{%$��̅0�3F�p�v�(B�p&���܃p�+�T1���ˁtL�!Y���1�7vKp�ӸЀҖI D�!�I�w� ~OҬ�p��?��'���=�Ѹ�$�|�B}ikq
D0�?�	���{HS *
��H@����$*a(D��+]D�Jh&&RR��P��2�,�Ja)!�4�~�.?I
9J�48���a$9��a?�͟�~�g߹�����V]�c,.��췜������y���9�Ȟ!�,!�K(�0�,��2,ϧ�>�j�!
! j`�c����kM���ZCJ�+	��$뵄���5�}�j�i�'��S���ĢU/���ii8��i� ����P��4c��$�m�lnq�$4o�RM��r�	�8�0���Nh�!I3[e���g����;��&�o{ؚ��{N�!`�L��-k#�x�S_-#�!#�p��s��,�L%&O��ݴ�%?K��~���˭��K	1���$�1�#YXR2[K����bDn~�,�٠�M�
JB��B��1��HS ��Ƙ�4��uw	�a�l�C@t�#8<�FFY�H�"�G�\�1��$IIƻC������5������1���
�)	�B�$���bt��
0�\.�nt2*a	.$)�
$���)w��"�$`Hb�6I !�7>#L�#A��R>`W�0�5!u.k�a�0ᚂD�t�HR\9ĉ�$B�F��]˩!�bD �ő����f�F��"B1F�(±�ŃƇ74j��R 6��J��w��O)-�h�ρ��'�y��6
a�LL�� I`�M�H$	FW\� @�2��Gt%�D���..$5K����&�C�&ͤlH�8F�F�B�b�<�	VbX�	H�F�R���Dd$��/{���~/�a��5�D�ALL�ZB��D ��+B4�R1)aK�ki�f�FUĈ4>l.h��	���D��MXĎa�㠐`ԔaI]0�!�Ԭ.N��%��rW��Z�~�0"�#B]B$Y	?n�����
bB���5��L��Жp�\c����HX��9(L�8ğ���ϴe������i�3 ��cR)�bO�i�e�L$9*te1���IT$P�i�p Gdk*�	�bF�L����)P�e-�5��I ��!�~��Á).%�f���)�v�D����$��M�����5�"(DlA�n��ߤ�BF~�~x��3�����p8�cB5�#$+-�,1��?���]iO��"D�40��B�%0�	#!�|c�W�}�J��L� �f6q6$!	�5��W噬�-pR�s���0��	q)�?B�D�JI#"D��9ˈ��5��rd�Lbi�I
K�9t�0iM�F&�W
$&%��Z2��a�*��B��ŭmm��V��BB*��������!Ĝ��y��}��[��G��)����9v�j}��т��)�e���7vK��`�.�ܻ�ς'��뷺۷\hlf콷f�7=�pg�t�b��Nrv��<ps.ݹ総y�t�Ć�b c�[27�m<U�6���s����4*�E�C.��hS�-�6���2f��f��5�m�i�j5:#k�Nw����	$�Lȑ��{#޷�:���{ѢS�LC����O�؎MM��7�}����R�lh� �q�:H6%HE�I R(���X�XQ�H1�H�`\�Y��&�u��S&1}�F�[{���bF##$ F"B1�r0��6����a.j��7d(H���!"HH2�X�S����r$d �6��.J�r�$M�.��	�:�,N$ED�F�u��Z�h������ͽ��F�+  �+��*X������������D`�R$� �A Ba
������h���$��~�1(`j\u�$�a�H@�k	������D$�Z K�l�$�	���	>")aJC���>�>HQ��5�]c�߾��6j�XB	�����B_c��0��Gv�k�N���^��:���D��k�k�|��m}�#iMk�u�bJ'�o����/�}�&iz�s�֛DY��ʄ�ȕ�F4�#0c�S[ԛ�S�)~Z�Z8�!&i��k�2q|��ш��4��k4���.����	�����}�H�B��lF�#С��!>��ݕ����v/D5���B�K2�v,@>H\�.k��o2�H�Sj���bE�v-�&�h�.j$	q" CA +
�57�$p�cC!p7#.F�0�@�#��.I
@�s�Vi�X�n��P��A4D�8l��._�g;�W���R� Pr0�$�}������-��/�K䐌F!b9�8����B�"!+F��SB4d4��\�>��gu�� f��E�λQ��{��I)�
��
F��h\�]�����/�߭K�4���w5V�iJ�bE+)'�	H�Qd���+5��bh��	V�4��w�Ȟ.����'z-���O�������7��"!B%\��'oE�B] BH������8�|I���O�XD������d!I7��o!��s|��Z �$& x&���Z!L��"Hd ��6{w��B5���9&K�F�
ۘ��V�Xgs4M��iur�71�ß^��<�<�ۋx�ﷃ�0�,-9�X�|���t�����0��A90���U
mi���i�*�Hzj��M'5F�C��Z6�˜�r�����}jM%��p$	�/�^^dީ��H	p��p"�H��T SRBe?|o�oW��_�7��!�pH�J`�F faZ�\�ԫQT�;����%�?L1�mFӐ�N����ރ�`E�A�L!R A��H�bŃ ĉ�@�I�+u�Ц��9! H@q�4�l�[� �������/�j��?�S5�2�4����
�A��
�F������3A+�6��M���Gߚ��~a �B"FX ��H��O��hdc,"�R`",�!"�H���!���#"�d`ՄBIE�R, $aV/^i��k�1bG#`�#L���%$>ه�y��,��ĩ�	������ ���@��F�Y0�RhͲJ�b��i�"Qk���H� ���|~?��̮:a\�@!�$K"��`�f�J ��
}�}Ɔ�b�e��7���&��@$�),�#*F�d�1� F0"�R������7$�&/R*�,�)(���,$d�c0 }k�D5$�1lJ!��l��f],2��Z.�1a��i! FIM;!h�s$�B�aCy���:HW �0��5
a�4�eܼ͜��2��F� J���)#�#�c�$$f�l���R�d3#?q����|Օc� �$c(��n�ԅ��Z�0�S!E� �a�$$!B%I �-X|;��b@��Ɯ��bOSb��D�H�c
E�k�$�4�h!XP�٬6M�7�\e7e�]�ݻ�a���Z�4#y�������2�������Q Ѐ2dH�5bBF#B$5 ���h(	ˮ�G��Kn-�B�P�m��kn�� ��  ��n������E����h�=#.�]�Њ��'n�*y�cs�9�َV��mV��%��Z��f�O^�"6� �T�	4��V�#i;4u;^�0�q�&�P�A�����]�����a$p [j��F��oU�#x�&�=�\nJ]�5JEj ]�����[����t��CRpu�uB��v�ꯨ���m��7�;Im�k^B@H��h�H��ŷ��w�¥���=md�JKԵ�0v�OR�d�zy(���6��%�R%���]����e�d�l��N-۷�U�e�+[k�h$:I��m�$l-����n�F��K�)�V����jl�5UҨ��j�l*qg�`'Et��M�Q�W�v����e�Ku�V��� m�!m��� �m�@� �sn�e� �E[�Y�l H]6���@[t����ݖKmmx���&V�}�}��Vԫ,���vl�f�%�m� �h�-�`&ٛI�@�-��3l�6��G� �l����m�� I�N��`�� �6ٶ���I  ��m�� -� p  m�V�p  m��� �  mK�R�*t�WJ��@�͹M�l6�M�m��3k&����D6ۭ�m-�	.ؐpM��ж� I���j�$���)UR�m�+ҵ�*]�j�����TҀ�����m�� 6�(RD�WUJ�ʡ�t�`aZ��U����e@�n�mK5�m�D H�� e�ph��XZ��C��U@Xp  h���6�$�� �v8we� ���`�k56�
x�9�=�ej��٪�[��d��$c��;K �h:KS^Yf��j�ڣS�T�l� ��U�G[W�Y� �   ��@��m�Z $+F�[� h;r��.��M˲��U���͎v�ƶeC�AƩ���N��6U��#ȗ6Fr���UYr8\�7�Es��K���a�g54\���ɳy�N�B���׬ܗ����T���[@O��.̯J��;�nآ�����~>�Zy�ԫ� �p�ZUlֺIe]�lB�˷&�`���n�R�m�]��H �p�I� 5�@ $p6� %�kp      lzEӖ�n���6�!c9إZ��Z��y��!��۪�m��%L������ݶƎ���'gB+9�-U�W��*�W��Blv+f��j�m�
@[PL�]ʵV0�j�� v�X�1�,�ľ���h/bۺۛg
 :&
g�B�UR�u\N�!����:۲�֜��e�m�)C�H�}M����
S�5R�\���@ ���z��l��jf-�t9��Kh.����ۮ����Ŵ6��M����n�"�T�v�\�pUJ��ҥ\��I����`A��l'sm�m�a���&�Hm�@m�-r��9U����j	6��m�4۪��� ���-��m�m�p�\Â�X��6e�Vvcm�`�P.    �l�d���H�ݐւ5�6,�%�:�Y��i�Iu�.�jK�1��.ʵ�����n��uG]2�����5��pI�u��K���%�Q�<��!��ojv����ٷ�|c֠ㆤ8��9Bn�^�B���`N���fQ��;�Uc�R���
J�D�KR��P+ҵ,�9�c��J��"�9n����@�$	� ?o�m[hڳ]rDL$٥�F�	�\�T�Z���P1�n�A5Th��e��	T	Yy�V��j�V���I�/C6�8-�R��w�}� ,��I	����g`6��mm˻���Ed�)���3����m��Leʁx)`BV����-��cm���cOM�� �۞v�2�.]��*�]U*쪯m��ꀳ�U�[v���P6�k�r�X�S��Q(��`�h�.�ιn�n[�ݳ������m$�i^P�kN�^��>]��m�A!�	�bA���WX-��rq5lt�cԫ��	[�T#���[
�T��n�T =��Iж���n�{Bj��U�^�W�D�*�i�q��k/QR]��m ֳe�MB�#�-�ѭ�2hL��Wl-����"� �hd��;&�� ���[p�m��@    	/ 8��P�`�x[���i4�8l��l���U*�KJ�J�U'��)�bWU����lp��v�e�X`���*��@mT�RUV�[v�Im�Λ\��	WgH*�Ut��ﾾ@j*��F܃�W�L�$�yn�$�ٴi3"��� {v@W��:���oPH2[Kr� ��uPR�lV݂����y����V;p�%�n6���ß�0��UN�h�.��6�m����S&��⣊{h/*��#�URZ'&U���{la�`sq�T:*���*��r�:�f���hԯ,I#NW�[�ְ6�$2���j�����z��!6��v -�^���ق��:�T:�^�lK�b�K�^�4^��n�� �3���m� �� ��Iͻc��Yc��!�
�9q�����ۭ;`��  �6��$E�n������Z��.  �i�� � ���R����(
Kl�R��UU�� ��OK)��mN�h��[�m��H 8 �ȵ��֝m�d��[KV�mH � �{{t�i���M�s��m����E֪�8ڀ����� �� 6�R�R�@�ù�#]�1䆰�6��VU	���e��`��d�� Ť��#q��6��
�Z��)��B�ݍɮ������Y�pB������l�{TcZ� 
]�Z��W�jV�T{k׬�,�:
�� �W�-Tj yj��d�F��l�d� ,K��j�(�i-������Y$�U@�gJR����gl�ʹ�g%7]�,T���ےH��b���}$���l�222��Uƒݔ��\S=�t�z�F��]�UV���Mu[mJ�,K��V���&G�97�r���v�u�<��<�ü��[2����U@[T�uJ�v�T�*�
�U��+��LŭSIKҨ��ζ;K.v��`%s���\ �����ٻ`t$7U�*ռ�l
�Ɛ�rYډxYd��Ņ�,��s��灪ں� �˯M�m�,�J��8��v�t�T����ߚ�p�-6�V�F�n�4V��*�A��6���^�^�yu�� t�V�ʽH!��	�����h  m [r��eT(��R�V�T��:sH ��@���-[f;�7Cm����f�9��֭�m�l x�j��P6]�Y^�g��    �+���mG@R�3);J��h��6�  �`m���K/  -�  6��mٶ6͘�3��rA��� dְX`8:Ûb�|��m���m�N�l�
�ʵ*�UT�u�[d�M�B�@qm E�f�$���l��
\�6T���C'C5rl=\�8*�V�*�[@    .����l����!�'m��]k+����K���J -��	 �l�Qgݷn [R$�vmE6��+��mR� �� �۶ZLѹ�'��"j���c��:I�9��]�8v��
�m��66Y�Zi��RWE@�z8�U�"����9�r�ۯ�iV7Z@��m�Q�S��d�����,���h��h�H�Eٳ��86�U�!UUV�R� �6�_mG �����uT�����cm�[I  l��<� �uR�l�]u;6� ;j[  ���lh%�cm�H� m&m��t���\$N��jWf����EZ��	��M��    m2 8 8  �-���m1m�d����`�4e�,��` � %�Cm�!m  �$��Z��TU1[�xkg\Tͪ�eeZ����5Rz!^.�eZ�մ���{�N2tmU�19YM�S��HUO��C�'�-�E�KMm���Y���uU+̫ /)�Z%���m IoS�D']����u�:ę.z�H�.���Uڕ^���TU9�#�[mJ�ul���R���B�yz@�fհA�����;N��
�69��U�o����q˃�Ί�n�j�)�PI�p��j�j�۫ey�]�hԪ�UV1p8����M�		:�ր8,�+�;*��V�v�Re��5HR��qJ1t=���;��;Jښ��K =�0����Kz̹�f��ݶ oQl.m�n�6`�Kq�p�6�TuQ�6�͖�7��c�EH[B@�f�8�m��Iv�m�-��ڶ  m�m���-�2q�����[An���[�A}hHp ����jC��UU�������`�e�ʸ �M�� 햎�F�;Y��.�	�j�%��`��I��6�ٵ��7,�q���Z�<>ۈ����D���rL���E8�N��&-���6�3;d��	�Xy��U-�J
@���uR��m���#Q��Mf�̘t�)$�i(m�m�	 ���:�Z֤��ˣZ����*��Q]�ب� �+�Q�R/�A40TdP�!�� ��E��Q08�A*��C�(�4�B��pW��T٥�QqUM��F�_�h8�H#U^
.!�� ~��䈛l$hȪ�_�@�*	���:��`Ca>6.�^���`"�EAٱ�~P�T�|��/�x 3��Q���A����
5C�H��Z�F"�� �Q� �^��"hy>TH;E��C��6����pq���U�"���: �Q�? ��thTD���T�� �� ?*�E�O��>U�S�N���?(�b |��y�\j)D?*�ȜF������N�B-�	�(�³Q@��"����R>,J�� |`� "���M���u )��
	�� Rb@�����O�> U�~�p62��Dؠ`�B? �����T�H�^)1,I(����	�@�"WA�#�� �Ac b�@?�E��p�� �*�z�U_�PB�"� �� ����Tv�"��E� ���#��!�V.���q.�$ �T~տ٭k.L�Db�N�0��+�'v����!s��Ψen��_�:�2�/6��t\��:�X����l� ��p���$���\쒤��F8CGh(�`�gB���.�ݠ� H9�U;J����t��$�����Ij�)��f�r�v�Z����$�8���M�'X�W�P�m�CV�^7%��m��gJ��1FpX���H�H���e��nKȹ��x�75�m���h�{�|�1Ļ-Uʸ��U�j����0�콳��]�Ի�V\=-;���6v�W�-�;I;�I����d�j)�m�n4�BW�!��*iӸ��2���Sb�X�ɺF��B�γ���s���'�K�Qh���g`��'8�G�xʔa�ݺ���,U���)��{�.J�b�=�qi���t�	���k�lMV���8�=��g��[���4Տ�3���X��bH�,ԁ�.zݍ
D���s�9�Cj%�S�<Z�7ii���q���i����ݩ��)xC�Bɞ��K��e�Ŗ�ط��`n�4�E��dl2�U��%J��lK�]��PI]�v�x���$m��I#��d����֎d�uk�9&�S�v�qN��{M�q:�̶�]qu����V���v+S�5���Ycv{��-�E큢`�@CvqS�HW�f���]=�<�0	�nW@FB�1���U�W{I
�Y�0�Ym*)�&�#[V�e� �n�������h����I��%�/V�XBwfV��"�n��öF��Z��W>7n�+��ۡ���\�BZH��n��bR��u�U�vɯ`�`kԭ��7�*ҫ�:]uȄ�҈k�Jsi�on!V�Y%���&ɷ4mbb�]���vG���۪Wz�;�܁W<G	!����5=�%��
��כ���]*8�bjPQ��%6C�6wa栲&�� ���ttk/���ٮՊ��
�9�.Y]Q�����A!�!�A�A�)��"���B&��t��z��ҍ_=����cv�u�p�IM͍�e݇l��ζM+��cv��+An:�t������������\5
']7=qϬ�=�t2����Ԏ.�0�ԅ�Zw�]F���z��;�:�z�VW�ݮn����ؙ��-��[	�[d�+��T��[l��8d)ݛ���1z�79	���&�lؼ��捎N�k;��l�B�~�������@��G�<dym����n�M���n\�����Ü&9�>�@�l�?/r�o��_�����[����Dच�Z��w����M �l�=y]R$ɋ$i5q����{���٠yu�@�wD�'1
8�)�@=�� �h]k�?z��g^y`Bb��2LQɠ��˭z�Yb�u���Y��u3�����B��%嬽�˂㴳�/���>��3v[�'On�]���&ܟ��~���e�@=�� �h��W��1���]w.����!$I�4���ǛI��������h��n�����('c�1�&7	#Z�Z���@��^�޲���^�D�bɎ1��z�٠yu�@�YZ�<�נ�{���&8���<���?k�s�zu��m��-��<����S5Ӹ�ͤ���/Ohlnms;���'3i���wl%��r݇NRM��_��h]k���˭z��w��0���$Z�Z���@��^����oؐg��>`ɋ#�Kdv٠�޺���h�,�fg�X$��� �E0���뚻�}{�sr{�������NM˭z�Šyu�@:�4�k����F��܏@��X�.��[f��ֽ�s������D�����N��oQs�r��+�޶�z����g���pӆ�c/I$Z�Z���@��^����h�ζW-��G]�@�{u噋�#���z�>�@��^�ga�<U9Z�R�tϝ���ok��Ēo������MזK ��	�j&�`�۹�=:�`��DDjH���� Y��5�����Χ.7����$Z�Z���@��^�޲��{��.�%#h����6�"z��Eu��n�us��{h��3s�nm�ƣ�k\ds!#jH���@��^�޲��bY�}���:�'�TJ4夎[�<�נw��h^����@��Ң(G��٠9�oc�?�٣٘�~��yw�=�q�cs&,d�⻺���Q��� w^�|�`���vz�D�IiF����m���t�o|�^��||��m�,Ŵfb���4���v��	mJ��w=s�����cl��6��P�8�fv��z:�RǤe�#i%s6��1�k�R�ԫhll��`4x8mb��ꐍ�z�s|����kV��K���˺��m�n-�+�z�%]]�cM�X�:.�hm�p�<u�Ԙ٭�`K"�DGE�$)���5�$bIK� 3�lu4U<<�{7
ஒ�n�tJ������ݽ}��$Lҵ�D��t3=`B���=��g��:��f�;'[.ʻ��v(����pnM�I%�}&����l_�$�.��RI.��ߒIR��,np��rMI%��ؿ~I.]w��]m��$�^�MI%��N�s�&�dRcNH�~I.]w��|�{w��o���6��;�׽��u���S��RY�M6�f,K1I;�z�i$�}���K�]�~��\��=I$�ݜ��p' �r~��Iz�5$��b�����t��m�w���m�1uU�5�nY�띶YZ�nz���q�â�i�V	�+e��v���z�`���sҞr� ���om����M6�s���,K�m���5$��4O鍹�2bd��$�_��7�� �YP�a	 I�F3�	��{�s\嵷���6��;��߳31I�)�7[�$���s��]o���K�ɩ$��i��Ir��$��yu$����"N[�����I�z�6��=��m�OCI/^���-Y,�� 7�Q7Ԓ]���$���jI%��~��B��j �{A����Vy+8#��0�=x��)�í[��)�]<u>,�g�1�bn&�](6G!��IwK�ԒK׬��$��\��|��齶�v.�V�����k4�Iz���$��k��z�?~I.�w��Y�����q��'��$���Sm��M��X�śXk\���m��;۽���2W�cc��crI�$�u�~��]��-I$��g��$���RI~�Չڤ�DԬp��{m�rwI�������m���t�o|�om���@�u�r8Y̑u����v��$�/�\�����Z�6�;0��
BԨq� _���?$�^�MI%��i��Iw;��$��Uߔ�p�3a��� ?���������=��m�ﴮ�m���n��$o�j���s�i�rMI%��~?~I#��MI������m��{n�m��s��rʫ��NC���$���~��Iz�5+�p
	�pB$A���rs��/{�XR��uV�e�4�m��;w����X��n�m��׍����A��ms���uc��H�ӞN����F��ٹuK1	IN�n.�gj�޺d�Xr��� ���RI{�i��Iw]�ԒK޶~��V�U�cc��crI�$������ڷ��ԒK����$���RI~��b�UR�����|�u��m������I/[&�������.��H�!m��I$��g��$���RI{�i��Iw]�ԒK�r���LJG�A9?~I$�l��K޻OߒK��^����ߢ��)*$"!޷���gr<\]�J
(�c�=���Ύ��&?�}̼.>��]y��-ӳ����-m���<s�&�zV뎭�OE�`�g5�'�f��� ������X�v怇�U��ڻd�vś��ӟ�S���M�ݻ'y��C�����,]��H�r�ʶ�h��Tֶ|�/��;5�rַ��W �(+���Tx�-/s<kF��-$��$%_�{��������Kz�hN-�v��i�47+��pŢ
\��n�uH;،���gm�Je�,���'�I^�o���$���jI%�[?~I$�l��K�غ�a�H6�r�$�u�I%��_��$���RI{�i�����]aJ�QUnF[CM���v�ߒI/[&��������$���x����Ĝb���$�^�MI%�]���%�wCRIy����I[�%p�����[n�m��u�{m��;�oa��|�����m��ۦ�|�uܹ	$�(��qZ����<�i�i�k���v1x�Oeݖ9�cqdncŎ!�IߒK�������m��{o�bX�#o���om�y��	ar��m�>�f��bX�U  2 �
�M(�S�V�5�t�oﻮ��m�փM�����cRESuѼ�Y���w��߽v��$�u�I%��_��$�,�pcQ7$Ԓ^��~��]�t5$����$�^�MI%��]qG�,o#���$���jI/?Z�~I$�l��oﻮ��m�g�tC��n���2�=A6�m/tTZ��1.�Ӽ��ش/m��SKшL	���$�$���?ߒI/[&��������$��sC��#�n���om�����,Y�H�9�x��o���Ԓ^~�����cm}��8Lhay	-�M���k���|�u��|_b��]5R��,HA��"ȤF���H1"@����6��a�]2DB�������	!H���*��W�2		"�[ �������A��P�I% ���ccB�,aKRZR��1�i`@�V��Q�?$!��BI$T���?8C�L�!�sP�H��H\0F�]n�Z����bn~�1!#��5�\�A$��4�!$D��'��:7��t�T}�ԇZT�����"B�&�(9΁�f�HVP��BB�E� =Gx#���W�O�A6/:!U~DJ�l_�$Z����h| U �
�D "Aٛ����[m��[{��Z�j�H���R�om��;��m�>�f��m��ۦߖbII�{~7��/ؠ�pd��4���$��k��$����M�������o�wZ6��yo��h#�:��i�+tg�r��z	H���t=���G9�nۉ���X=,�_��o���m�ϻݭ�����K?�/�u�� >�]�����4U�R�j� �7�9D���g�V ���>�B�Tt�=�3J�
�]U����z^�áb�oϝ��罥�8��]aJ�B�T�v`tB�
v��`k��7����PD?�~��D��E{���ʤ���8�7��W����B����}��>}�vl�躡M��ZL��9�[�WT��ۇ�pj:�6mh-�oj5\tt쮷�����W.v��u�����m��뮏�:��;��#s,q�Hh�)�yzנU�@������Pu��`�I�@���@��^��YM��4�w:�ɉ�K���W��޲��Jh^���ń�$�1�4�j� ��� �B�ל~g{� s�y�$_��!�Jme�55��{[P�;��"f����㵊Wm����u�\gq]�t\	��V͓9���2{)r�H��Z��j2�q�Ku3�6��qȖ�ރ��UY+6Ĭ1"n̺�6��nM�V����jH͖�˕��J�N���泓{nn� 1aT��S�{�T����;n�v{�6�*dpt�8[bl2:i�vn�t�� ���2��I�U-g�6�� ݱ����./*Y����z
�1�p��U$����Z3Z�����<��9�}~���z^��z�h��*LP&6��R��z}�h���/�S@=�د�����c��z}�h���/�S@���@�9J�Lla_�	#�=�)�u�M�ֽ����� �ȜǏCp�^��<�k�9^�@�����J#"5�x�P�!r\����׍�N�\8�k5�g���֖<����88���N��z��X��(�� ���n���M�F�f���;5�ϓ#9;th�)�yz׿$UO�$�7I2U�����m�tL��u`����\Q�ĞG�7��hzS@���@���޲��,�4��Cr%!�yzנu}V��[��u�M٘���l*�I$���tR�-#��'�\��f%��{ku�-��������7��SUtR����>�Ӏ{��`�����>|�����뾙]Ccȋl�}���Q	D����{� �z�9$�d޸��y���n��/�|h^�74�����0F�H�Q�(?>��8wv,��ueZ�,cI8h}�����=���@����y,��w^4��Sr��W.�u�p��	&����w�����o���7	��(�*���gR���+u�}C�Ќ�Z��#WL�]�[�����u�Fd�9i28���4�)�~^���bY�a�N��r�N�	�Ta"�V�{lϔB��BQ���}X}]��}��k�,X�M��Z�����d���� ����5ֹáB�S;�ذ��ƀ>��9ܪ�%�RK4�X���p�ذ{l��
?D$�
!)���<�L��ٹ'��n���e�Zʂ��\���X(�ݜ~ӽՀk����33�{�A�;GiKo"�C\�ػz�������`m�[/kW��cg_��爚��TQJ�(�_�߯�@m����ھ�������}�"��"�jf��?O���BK䒪;�����`l���x�ߓhjbqA��z��Ӏ{��a�P��
����0��Հg��&H6�#�C��]�}�4�����У��g}8j��ST�.��jI��`�ـ}	%������8��,�Bi@�P$
�kSV�a�W�ݞx�`]�Ai�VS"d
 ��Q�܄��v����L=�bIX�鳪�����õ�*n]�C�+A��N�M˧5h�,tZ���֑�s����\��Bԛ��%�[�ɋv��.��:�.#�SuLZ6Σ{Q�k;��a��V�]�i�VU��$-�N�A&ue�.T�wI�t]�d��.�n�2��q�_y�����׵���Q���rȭŞ�ڑz���bo:���h����Bn��ͳ�?�wo��|uŵ�#@�������`�\���]	/������eVX�-"�Y�9�ν{cg9�ih���?O���!)��'7�j�.�PR���u�,^�0脒Jgӽ�@�?�Z�ȉב9�8����Q$�B��������5�s�В�O�ﶴ��RzR[V$�@~�7XB��o����`����o��	K;6��\9��5g���G	קi����ئN��ˀ��~���[�}��p�UE�]~�>��׋ ~���!��z�|}C�	&D�28�{������
@#����M��&��+��bI_�K�)�>z���h�s�^ŋ9�zy��rK[#�r��]Ӏ~�7X}	|�"���p��X��]a��B��נ�,X����ΟN�kŁ�(���� ݑ�tR��SUtR����k�侈���^�_����ֽ�S,n7�&=��ڒ��d��f��v����_Vԕ;���L�b�5�2�[(���s���������D$��u�8됺�Uʢ�IGj���^�,�ى%!�߾���p{^,�P�)��E��e\�+k�����=�;�޽%RH�_��v (�"- b(�
�BI}
G����X�_}8�F�\���+VL�٠�ĒOݾ���}� r۬��սՀ]�tR����s4����=�x��	us���{�@��ZY�X�Q�d�dIc�D7�{sq 65�z�=�\�=�[���W�wwv�G���y�����~^��ֹ�J?Hn�ŀn������]TՓuu�~�7YСL���8��X���ٟ�D���x��xۏ@��~��׋�"#�U���Հl���SG/^Z�c��ŉ��ր�����r��srC� �(E`�`t��0�~�9w$���5���h̓UVM���� �D(��m�������@}�;��;�wO"aP+P��Y�GE����u�c�\�ɀ�{dV�y��s�H���`���H�9�ۏ�]��@���׋�"#�O>� ���h�WE]��
���\�$�(S&��XO>����΅�)�b�*�������.�p�ذ/]a�(J&};�Xu>��T�̕J�j�sV�>I/�%__��`/� n���$�IDS}�� �Ҿ�����v*��Wu�~�7X�>�����W�o�ŀ9m� �8ؒ-bb@�G�:�,�5��i�Z���C]3p��C�?	��B�E��9�m#$c�H$`@�A� I�(�h�!��c	  �DaHHBD�@�b"��x�ֆ#!1!�X�!B!�F�9��
ƄbK++[YYIYHR��#$��$� @���F
1���F1������D���H�b�H� $F)", D"�$�	h���4�H@�`�����S0C2P.ƫ�i.��b1�����>+���AHňF�H�O���+�D�X!����
*���TS���%�Y��m��N�2¶�(W"˓�۰������ )b�;����R�kc"��T	��S��˵����i��3�������R�֗�.Ú��Sƒ܀��l�8��9�\<�t��]��ۥfL�6[�h�qrL)����X�6�WfT�m�g(��������G��:$,�2�X�� N�dCU�m��8�ڔ�cJ!t������;*��kk�1t8bX8�yۃ�v�q-���=<2�۶�絷c���nܿ?f�;4�A��V�  6<j����*tIۦY�ۧ	�Y�n�{{�݋9���g�Rg���U��)
(��髇5��e!s���[qcN��mI��zm<E+�&7V�Qr���ո��k���$޽���v6 �;�|��ngm��z���8w��ђH�AH�2���SKVۂ���2�G�� 旝�V�ͣ��{{kYn�Ng',N�u� 6 jj�V�(h�b�i�8��f�����W` CF���/;���t�[l=ɷ���N��Z/�m��m�n�bl��Bc"6N�^WX�������@B��㮨7`��ӭ���@�T�yZ�7
��s�4Iڲ�<����Z�v�f��� [�z���Z��L��d����d�ջj����@m�v+k`9��u�x��Q�-�km�Ɍdڼ�ȷ[��h�5 [#��W�ҕ���9�g8kw��f�2r�g�,� �o��]�O�!�^�묄���LҪ���ݝ�U�v@��;jnG	pl<Rl;+��c!3GD��5�[[]3D�u����3k��t�"��c�{Zu�Y�3`h �
ۯ%=V����M����'m�[e�cO:�Nt��5U5+f�����e�j�&O�'�}벐��;7]m���R'%&7���fڎ�ݞ41SИՋlײ��gu�b�8��6�ׂ�Ļ	�#b9���o,뀣u��GU�㘪�5(9��3;[����<�`�i۬���Z��6� ������b�kpd��0u�uV��������+���6���@�<E���)�����S�_�C�E���2��f�Ir拚�u���{qD�Wp݁P-�yT,��%]Wm��������xϤ	n���;qW����ŷT 	\�8S=���=�{;]�j粢oNPMM�ˌ�zgY���vL:q�����Ӛ�F��;d��bX�C�=�����T��5�2�V��5�m�ʍq�լ�]lNځ1�&��W[z5���cx�pR�`k��X]eķ�,I~�ƵZ4=�h��Aĭ�H�a�=���5�By;k�#]$v"�	N�N�N�H�����eVX�����l�߿M��r��D~���u`�w�j�.�B���p{^,�B��Q���V����-��{ܰ��i�x���4
��Br��s܉c��r&D������r%�bX�￸m9ı,O}��]Lֲ��S-����r%�b؟��{6��bX�'��z�9ı,O��m9İB��{�ͧ"X�%�Oӽ�fd��)sY,5sY��Kı=�{�iȖ%�b)����"X�%�����ND�,K�}�fӑ,K���ݤ3�lbwTtwKk4=��"�V��n�u��͵��Y�����������t��9ı,O��m9ı,Og���r%�bX���{6��L�d)!}��Ӑ���$)!6���d��SW��3\Ѵ�Kı=��i�UGh! �O ʋ[�
���,Mgy��r%�bX����Kı>����O�DȖ'�O��7Yh�"%�X�bf&bf.N��4��bX�'���m9��,O��m9ı,Og���r%�bX��ޗ<��k�ta��ͧ"X�%���}�ND�,K�}�M�"X�%�����ND�,�HdN���ͧ"X�%���~�疨���m�ų131}�o�iȖ%�`��{ٴ�Kı>��ٴ�Kı=���iȖ%�b_�T#�)�l1&��Ja K�g�-�]�kg�Τ�n$vf��˻��wG�i��ny2h�&f�ӑ,K��{�ͧ"X�%��w�ͧ"X�%������ ��&D�,O�����Kı;��OΒ�ڲ��%�X�bf&bf.N�ٴ�Qı,O{^��r%�bX����m9ı,Og���r �X�%�~����2��d4d5sY��Kı=�w�iȖ%�b~���K��� I��{�ͧ"X�%��w�ͧ"X�%�{=�h�ff��։3%�m9ĳ� "��s�m9ı,O����m9ı,O���m9İ"F����&�)���z2J	�d��V� X�{��[�H�r��si�%�b{��6��bX�'�w�6��bX�'��-�3�l廣��G�ײZ�aR�����[�4 �'���S����vuų[����Kı?g��m9ı,O{��ӑ,K�������Kı=��x�bf&bf'ξ��U9c$��If��,K����m9�,K��ND�,K��{6��bX�'�����ؒf&bf.�k�-Q�t [n��Kı>����Kı=��iȖ-�b~Ͻ��r%�bX��}ͦ�L��L��:#S�I*�!T�v�aȖ%�ʨEȟ����m9ı,O���ٴ�Kı=���ND�,��8��	�����f&bf&b��SZ��%��%R2If��Kı?g��m9ı,?��k��ٴ�ı,N���6��bX�'���m9ı,O��'��=e�,�u��,�vx�vW����/@�O�qֺ�-�n��7X�MX��N��
�f�l��N%���}�ND�,K��ND�,K���6 r%�bX���{6��f&bf'���Q�-Dv���f�l�ı,O��m9lK��{�ͧ"X�%��>��iȖ%�b{��ӑq3138����('e�r*�ZŸ�%�b{=�fӑ,K���{ٴ�KlK��}v��bX�'�w�6����������#U5T�V��IȖ%�6'���ͧ"X�%��k��ND�,K��ND�, ,Og��[1313�޹�*���ZE35�ND�,K��}v��bX��C����i�%�bX������r%�bX����6��bX�$r ��w{�����L���]J��v*vxma�r�jg����)n:�N�� �Y:����]�۾�X{];]Iy���$�U�{It��萐QW�s��䇷���p�*shgr'f�Ʀv��L�l�On��2[�v(�Z�9�
�e'�8^�4��@�Nc�lj�0��^Z��M��j@؛���'��VQ'l�b���!n�7hl+ے�6�-O4nPo�۽����{ݾ����q��KBs6�\[u�V�D1�m�JO;l�-u\tt�,�{���է�����i�k�-���������'"X�%���}�ND�,K�}�f��`!�&D�,O��]�"X�%��|�S�X�J;V�l��L���{�ͧ!���,O���ͧ"X�%�������Kı?}�p�r*ؖbf/��֧�%���#d��bى��K�}�fӑ,K��{�ͧ"Xؖ'��ND�,K�k޻ND�13����p��b ��k�N%�+bw;�fӑ,K���}�iȖ%�b}�{�iȖ%��X����k�L��L��wު4娖T�-�r%�bX���m9ı,?�"�w���i�%�bX�g}��ND�,K���6��bX�'~���s$�i���l+ys���k9de��������-ԓ���w�����MZ�����d��V��ı,O����v��bX�'���ͧ"X�%��｛ND�,K���ֱl��L��\�u�)Uh���5v��bX�'���ͧ!�Z r%�bw;�fӑ,K�����"X�%����]�"��DS"dK���?�.k�՘fkY��Kı=�]�"X�%�����ӑ,�,O��z�9ı,O��}�ND�,K1s�{^j�[����f&bg䠙�����Kı;�����Kı?g��m9İ��}v��b����΁��I*�!T�v�bى�bX���z�9ı,O��}�ND�,K���6��bX�'��ND��oq�����n����\RmEJb�$j����w��9��=n�ڢԥ���_v�����ڰ�u�^�l��L��_Nw�X�ı,N�{��r%�bX���lyı,O���6��bX�%�;;��Q§k���٬[1313g{�9�,K����"X�%�߽�M�"X�%��>�i�bX�%��Tl���S$�Y�[1313��m9ı,N����r%��� i@/6�"~ϻ��r%�bX�g{��r%�bX�}o=�f�K��d���h�r%�b����~�ND�,K�}�fӑ,K��=�fӑ,K���}�iȖ%�b}��d�TP�����-���������kı,K����ND�,K����"X�%���~�ND�,K���Ć����\խ�u�Y{Z[k<Y���C`�j�s��Cy����|2��yg��q?D�,K�����ND�,K����"X�%���~�C�,K���w�X�bf&bf/tk�Z�`آ5�ͧ"X�%�����ӑKı;����Kı?g��m9ı,O��NB�B�D*!I	�+鲪�h��3R�Fӑ,K����6��bX�'���ͧ"X�b}�w�iȖ%�b~����Kı?{���f�kYi���n�Z�ND�,F���wٴ�Kı>����Kı?}�p�r%�`b���؝���Kĳ����p��b�U�5�f&bf'�k޻ND�,K����"X�%���~�ND�,K�}�fӑ,K�w��{���?����HW5X3RD����8f��V�y�1]��g8XJzN������7�'�K*d����&bf&b�}�kX�abX�'{��m9ı,O��}�yı,O��z�9ı,O�����KP屒E\�X�bf&bf.���9ı?g��m9ı,O��z�9ı,O�w�6����S"a����ڋ�*(KEl��k�L�bX�g}��ND�,K�k޻ND��V Dȟw��6��bX�'�����Kı;�{o�.k�՘fkY��K�@,O���m9ı,O�w�6��bX�'{��m9ı,O��}�ND�,Kݒ{~��au5�,0�ֳiȖ%�b~����KıE{�o�iȖ%�b~ϻ��r%�bX�g���r%�bX�P~잾�O��X�nغ��6�Lp��2���ٌ��\���zi-@�K�ۯD�6�n�OFx5�v$�}�g�.u�̼R��Ww�}l^�uR+�ucywmX*�)k���p�d�K��gV-�g�,�A�<l�q٭����ce�ٔT��@�����6��Y[X����[.U�׎�ه��|ڌ�b�@�f�4u�C�\mA�fyn�lC�M9B=���Q�;s�G�Z��&�8��4u�WC�n��엱bY� �MY* K	(�Zų1X�'~���ӑ,K���wٴ�Kı>�{ٱ�Kı?}�p�r#131s�Z�zR[VWvZk�,K���wٴ�Qı>�{ٴ�Kı?}�p�r%�bX���l��(�C1>=?X��NWI]���Kı;���ٴ�Kı?}�p�r%�)bX�����Kı?Nw�X�bf&bf'����D�ʙ&�k6��bX�'��ND�,K���6��bX�'���ͧ"X���L��fӑ,K��a�������c$��V�l��L��]���X�ı,DS�}�fӑ,K��{�ͧ"X�%�����ӑ,K�����E���e�}-k��vԛu������z�c^�^��h���Nt�N�ݭ��K.jm9ı,O��}�ND�,K�׽v��bX�'��W�,K�ｿM�"X�%��;�}��sX\�d�3Zͧ"X�%��k޻NC��"���lX� �#�FaF2�z�P��~@Jr(.
�vH�H!"�			�*��� ��bX�����"X�%�����m9ı,O��}�NEı,Ox���kFY���a���v��bX�'��ND�,K���6��c���r&D�;���r%�bX��׿�ӑ,K����O5d�	a%�X�bf&bf.����Kı?g��m9ı,O����9ıDK����"X�%���Z�zR[VWvZk�L��L��>�iȖ%�b���]�"X�%�����ӑ,K�����ӑ,K�w������.-3�aC�5����N�R���oF�̽�1�-����ˌl�}��q}����AWl�-�����������LK���}�iȖ%�b}�}�a�@�2%�b}���m9ı,K�_j��KUnB���f&bf&b���ְ�Kı?w���Kı?g��m9ı,O���m9�D	�2)���_��d�[+�k�L�ı>����"X�%��>�iȖ0��2$"�l�p6$F-#��0�]AFz�n0�6��	�hң��N@���!
�4Y	!BEm#))D�ġ(R[!ZB���QMK!!!	���ȔfD�0H˘�(��e�bH�`�� �] �9	%J�t�	)$I!H0�i	�RR�@桾`H�m]H�i��X�AO�;�$�$d�����������p]Dz~D>A���N�hS��N��.���q`#q���_�!��H�'s��ͧ"X�%����6��bX���wMz�
�h��v�bى������wٴ�Kı>��ٴ�Kı?}�p�r%�bX���p�r%�bX�ý��5�����ֳiȖ%�b}��iȖ%�`?��m9ı,O���m9ı,O��}�ND�.����]����+ֶ��.�j\>��%i����V�����_{gI���a��k6��bX�'��ND�,K�}�ND�,K�}�f��'�ı;���m9ı,O�=!���%"%d�v�bى�����ｳiȖ%�b~ϻ��r%�bX�g{��r%�bX���m9ı,O�鸧�%��K#vIV�l��L��_Nwٴ�Kı>��ٴ�K�H�L��}��iȖ%�b{���6��bX�b���G
�%q��f�l��L�q>�{ٴ�Kı?}�p�r%�bX���iȖ%�T�K"}��ٴ�Fbf&b~�]�eD�%��%r�bم�bX���m9ı,N����Kı?g��m9ı,O���m9ı,O� ��V�����0�[]����㋷f�@9ͽ�O�ݪt�zis�qs_�&�f�%�r��
�Z�񉘙����߸m9ı,O��}�ND�,K�k޻D�,K����"X�%��{�y��
�U-��V�l��L��_Nwٴ�Kı>����Kı?}�p�r%�bX���i��bX�wE�����an]�ֳiȖ%�b}�{�iȖ%�b~����K �,N����Kı?g��m9ı,O.���V��,#E�k�L��؄���}���r%�bX�����"X�%��>�iȖ%�b}���iȖ%�f/�tF���X�VIGj�-����bw���"X�%��>�}��O�,K��fӑ,K���}�iȌ��LŬ��.�����r���VZ��r�1Չ7f�=�B9 .����F���t��W ��1���'�PC�f�9ĺ���d	wY��&!4��$�ƽ:�mպnX�����YQX֭�׎�������c��6�A'�;=nB�g�P�k%�s�6n�S�uآ��#/Z�\�,�%dݱ�NdU�׋^ӑɪg�K��������%/�,Bǉ+��U+*`��6�n�ŵ���	�5�H�8�4��ۅk���t��e�Y'�}��oq���;����m9ı,O���m9ı,O�w�6��bX�'���m9ı,��_}�VH�r
�f�l��L��}�{�i�-�bX���m9ı,O��p�r%�bX����6��ؖ)��E����,R�!ezų11,O�w�6��bX�'���m9��EX 9"}���m9ı,N�_��X�bf&bf.pW��9j�8B�Vӑ,K�����"X�%��>�iȖ%�b}�{�iȖ%� ؟��mk�L��L������Ж��ۭND�,K�}�fӑ,K���z�9ı,O�w�6��bX�'{�p�r%�bX���'o��]C5ѡ��]"ь�v�jq�B{7cb�u�N�V+�[�rs�%��qI��9)�����{��'�׽v��bX�'��ND�,K���lD�,K�}�fӑ,K��a=�S4aMk%��WZ�ND�,K����!@� �?"� %0��H8)�^�D�,O����6��bX�'����m9ı,O��z�9ı,O�ݦ�{335��Z���5��Kı>��iȖ%�b~ϻ��r%���b}�{�iȖ%�b~���ӑ,K��zn�����K��Y-�f��"X�@"-���{I� ([��8����w!%�'�=6��bX�%���)�&�3Z��W5�ND�,K��}v��bX�'�w��r%�bX��w��Kı?g��m9ı,O���-!�?�L����e�Ǿ[Y�3�pN	��&y�g������N�x��\G!v~IZ֬"$UH�NB����&bf'���siȖ%�bw�ߦӑ,K���{ٵ9ı,N�]��r%�b�����Nڇ%���]bى����﻿M�"X�%��>��iȖ%�bw��ӑ,K�����NA�3'��R�BZR�[Mbى���'���ͧ"X�%��k��ND���"�)�t)"X�}�p�r%�bX�����Kı;������e�5�3	sY��Kı;�w�iȖ%�b}�}�iȖ%�bw�ߦӑ,K,O����ND�,Kބ��rh�k%,�kZͧ"X�%�����"X�%�}��m9ı,O����ND�,K���6��bX�'s��[�N8]�.-ڴkm��e��؉���*��dv��N�˻[����*�ڕ����D�,K���6��bX�'���ͧ"X�%���}�����ı���!~!I
HRB��R���]�awY%�]�"X�%��}�fӑ,K��=�fӑ,K���{�ӑ,K�����ӑ,Kħӷ��e�Ypְ�j�iȖ%�b}��iȖ%�b}���iȖ �%�ߵ�]�"X�%��}�fӑ,Kľ�}���4f��j�iȖ%�6'�{�6��bX�'~׽v��bX�'����ND�,m !����}�ND�,S1s��O6[P�2ʵ�f&bf'~׽v��bX�
~Ͻ��r%�bX�{]��r%�bX�}�p�r%�LL���5sֹkj�����������c*sx��=t�v�j�d���*b���}���N��2Gl�X�bf&bf.N{�X�ı,O����9ı,O��l?�I�&D�,Ow_��iȖ%�bw������Z�Kf�l��L��\��Ӑ�b�DȖ'{��ND�,K�����r%�bX���{6���2*����{_�*�-�L��^�l�ı,N���6��bX�'~׽v��bX�'���ͧ"X�%����]�"Y�����tZs�I%V"��nU�[18�('~׽v��bX�'���ͧ"X�%����]�"X��#L�o���_�RB����F�VM]aw�%�]�"X�%��>��iȖ%�a�{��]��%�bw����Kı;����Kı4�N��(����;��{����J�[��y�z;ƍc���P�ve&Q��M�������c��su��s[t֩��̈5����hg�֮�0k�&x�(T�[����gtdK�D��ۭӵӱ�c�r�U��rw:�0�d�+�{ m�rn��,c�.��M��n8G:�"Ԅ����e�F#V��蚰F�*��7.m+t<62��W��c����"��_��`�"_�!/7�K�CY5�X曀ӓV���(���r%^��Wy��yW�t_�����9F���f�l��L��?�����Kı>����Kı;����Kı?g��m9ı,K�{�ՙ&a�Xf����ͧ"X�%�����"�bX�'~׽v��bX�'���ͧ"X�%��{�ͧ �b31}��/Z�mC���l�X�bf+�����ӑ,K���{ٴ�Kı>����Kı>����K����݋̭T�Nђ;ezų0�,O����ND�,K�k��ND�,K��ND�,��!�\��!~!I
HRBo�}EM�RU�z&���r%�bX�{]��r%�bX�}�p�r%�bX��^��r%�bX��=�[1313��jyZ����G�	���ֺŐ���gF��c�[@�����j�::wbW���V�n��Dհi�Wk�-���%�����"X�%�ߵ�]�"X�%��>��a���2%�bw�^���f&bf&b�|-9�)$��[�捧"X�%�ߵ�]�!�Qz��4Ȗ%��w�ͧ"X�%����ӑ,K�����Ӑ�,K��h�%�t-��X�bf&bf/�=��r%�bX�g���r%��"0ș����"X�%������9ĳ15���F��NWc�W,�-������}�ND�,K��ND�,K�k޻ND�,D�?g��m9ı,K�{��r��F��3W5�ND�,K��ND�,K䏻����ı,O���ٴ�Kı>����Kı;��˗-��3�Md�.f����A��S�l�1�e�;]v�����z�Y7au�w.�5#e��#��bى������{�iȖ%�b~Ͻ��r%�bX�{]��r%�bX�}�p�r%�bX�g��R��uV�v���f&bf&b�>��iȥ�bX�{]��r%�bX�}�p�r%�bX��^��r%�bX����Gi-Z�l�-�������k��ND�,K��ND��W��
���Ȋ|��F ��N{_߮ӑ,K��{�ٴ�Kı=�;�5j���&E]�X�bf&bf/��m9ı,N��z�9ı,O����ND�,������r%�b3{��褒�lr�*�-����X��^��r%�bX���{6��bX�'���6��bX�'�w�6��bX�߿��w߻��D�K�%5tҴ:	"�ui�駲h��ĐW�ưc�tq�b�NjL�a.j�9ı,O����ND�,K��}�ND�,K��ND�,K�u�]�"X�%�Oӷ��e�YsT�d5u��r%�bX�g{��r	bX�'�w�6��bX�'��޻ND�,K�}�fӑ?���,K��?��f��4k55nf�k6��bX�'{��ND�,K�u�]�"X�
1��>��fӑ,K��{�ٴ�Kı?de�[��U�[13&b�����r%�bX���{6��bX�'���6��bX@��M#�@1wbw^��"X�%�}޾�jh�Eѫs53WWiȖ%�b~Ͻ��r%�bX(�C����i�%�bX�￸m9ı,O���ӑ,K������~�p$���<�U��^Ջ�����OCH��h������u�f������bkZͧ"X�%��u�]�"X�%�����"X�%�����ځȖ%�b~Ͻ��r%�bX�:N��֌.��afZ�m9ı,O��m9,K���n��9ı,O����ND�,K��}�ND� ��,N�����RIS�l��U�[1313?~5���bX�'���ͧ"X�%��u�]�"X�%�����"X�%���Sy����	a���l��L��_N{�iȖ%�b}�w�iȖ%�b}�}�iȖ%�b~���6��bX�%?N��5�r�dv�bى�������]�"X�%�����"X�%��ޛ��r%�bX���{6��bX�'��,�`����D��&���D(����+��ErbVX�-��vA�(}����7 ��:nҍ��M�%�D�
�R3x�H, ����ݬ71�fE:l��>4��fMU���]�[�p����3B]vn6vdqhY[�k�Xa�{vR��n���+��T��xm�wV�6�iY�ѭ ̷9�  N�n'�v�I�r�yh�Ŏƒ�p<���cfj�Ӕ2(�f�ע"���mw@��酴$��|c)��Z��Z;&	���ѕp�
�\D�Օ�m��`�0�vj��ٗgLZ7)v[nWaZ�"���9�#nN�msydt/2�MRO
�ƢZ8n�]'*,]U�  ]w���n��ev}��N�����n�l�l��ь����|`I3�0YU�^L;;,��R��Gh.%ۥWm����m2���B�&��^��q�8�|e�]�{�T�.�u��grk8�cn� (pFۀ�ݘƤ�m%���0�Z�1���e��Ep`��g���2���;hx�sԄ*�nuU���puH�����P�d:bi	L�W�mr�g[���; �Y�U6ٖ-�p�]ppl��%�ɱ��f6�:6�3X�7[�E�����o�.ͻ1܎�`0�A��+�]t�rn��i�9���l��#�e�^N#�ϣv+�
�.X�r�&V[�t��c�p˒��v���5�:�Վ+�-�^�U,f�i�c�9�6�HA�z�ۃ�v�#Wm�1�s�1�=�([f͎v��§v,��;�!`��iӢ�2`1Y+��Ax�Z��;��g�3����=�t�������8T%EJM���VV�P6$6��i �p�*�
d�i�n+#��j��$�s,s��LecMl8N�JKâ��}�C�r��6� �Y��d�ԍd\.�D�fy�AW�6 @�j�Z�m��J�*˲�Ҵ�]	c��d�n��#@�c[!�8�稞��/=^5�ؗ�46�gv:Q�QZ��fų�]��ͷu���%f_+\�ɣ@\�����[0�o{ӹ�э9ծ��p����h���A��gZ�M�Z[]��a�;q>�y(�PLPtD6� �T���?�� tC��� AR��8*��@¢O������qWe�ٞxZ�J�]jt�48�5;�V��^�!f��E�'VMKӨ�;�z����3�#�џH&܍��P�=�����i(�8ֱ��(����onƪ�ݗ�[�',X5���
z��e�m��%�ì��7	e�[���p]��]�%��� �p��0�m�뇩�˲�N��Е����^��Ah�m��I%�0���JH^�ϒ�b�b�{��?�8$+��:lxmsU��%�xk��#[��p�	OA��#���o���^�m�s5sY��ı,O��m9ı,O��ߦӑ,K���{ٰ�D#�&D�,N���ND�,K���fY���)2��h�r%�bX���M�"X�%��>��iȖ%�b}��iȖ%�b}�}�iȟȃ��,O��g�
T:ʬrR�ų131}���ͧ"X�%��w�ͧ"X�%�����"X�%��N��iȖ%�b����Gh�-ʋl�-������}���9ı,O��m9ı,Ozw~�ND�,K�}�fӑ,K�^�ך�D�a"�׬[1318�}�p�r%�bX����6��bX�'���ͧ"X�%��k��ND�,C{�??;�v?��.�}>B��i�X��Cq��x�94IӼV�sخ���	�p��~yV⚺˚�4m9ı,Ozw~�ND�,K�}�fӑ,K���]��?DȖ%�����ӑ,K����j~-�ЖA�k�L��L��罛NC������%���!~!I
HR����;�|`�l�ӈ_���@����빧�ؗ�|h]��@)�X�cp�6G��u��-:S@��W��K��<�}�H� &�0k$s4N��?+��_U�w��h�K.�L��N��^�\�N�=u۰�;�Ѱ��;X47]��m�e`�E	U-��@m���]k�}��Gޠ��� �־��왥vբ�� �Z�>P�D���,���6���~l����V��,&8��p��`�l¢hR�"�$B�umנuv��q�:��(Epn,S�<� ��Հk�s��Q/{�,���?�	"Pcln-��z�2�/����s@��M�u4xD���˥θ⠣���OJ��|%�g���
�
�>��C��p�DřC���������w4G�h�w4�ΰ&����R=�n����ÿ-��ihvs�@m����nT�q��ՠ+\�z�a�/���{�`}�.,sd�<C�h�w4���O�}ݛ��ґ�S��$X�$2! "1	�q��ţ$��W�t��W�_��fcŋ�O�=�ƀ��j�+�n+@r�f���Z{��iҚ��sC����@[�4q�K:"�\�z���#��f��v.�]���n�	�������W<u1'�ȿz���Zt������:��@��dN�m��F���Zt�}	G�
�߻�X}]���x�=R��BH�	op�?^�������I&���K@y{�ƀ6p|�q�`�v��Lլ��8�^,����
1?��mh�kެ��U%(�-�@s��`B�˞q�s�Xu�p
��ՙAp'JBdd��YcB��&�&�]P��P�N�D����;<ͻ)��:��8�nlk���J�"7:�4Z��	*�I��)�l�[u�sI���NjsL�V�n^�:�W Pt��%����^��d:6-��6m��k���x�ݞ����͸��G�`nsMXĪ���+�;m�3�hى�6�0k�s���\H�-˶�z#�pO<�n9���w����3+�0M�{�j+��"�t���v�E�3$��n�E-mK(禗;'41H��S��Hղ����_}�t�{Z��(I%�}�, �����XU�E�������h^�@���h/Jk�噙!�z�Ԯ�H��VZ������׋DL�ݫ��ŀ{@��I��ӑ��,I��;��:���@o��������D��ۘ���8h=�`	%�����ϫ ��ـo���(�:�I@��Nc��7RC�3���#jw���.��q�b���ꚳ ���`^��=�rQ�9s�4��&��R
�������"���\\v�`��U��8�v����>JG�*�����<��2&����?Ɓr�����S@��z�jرI�1�Q�I]ݘB��%_/��������u�}�;��:��:��%T�d��v� �K��W�7_b�{l�Ǆk��œ���]"ч�rS���]���g:q\{��9��l��F�m��u�p{^,���Q�C��� �
t�V���8�����t����/v|h�Ɓk��ďu2'�ƛ��[�Qڴ��|h���C�ş$�IE $���a�l�#�Ю�P�G`!g���ܓ��ݛ�~��4�$K&51�i�C�����h|��@�����%<�����j蚵6U"n���Xۯ�/�r�|`��4���/�f�ɬ����i>$ӱ��9\sqO���� m���.�vY��s(���f��;|h�����/Oٶ/��@�5��b��cx�Y#��\�)�~�)�Uz���s~H�a�,s	������Uz��빠\�)�{ϫ�9�s#p��'��V�� ��fQ�Q�B��
"Q6�]w|�ܓ�ϧi�%��JiM���kŀ!B��_/��ǀ����@��zeh�%SQa��d&��B-tN���'m"N��D���WY3I�m[���]oFcN<i��(�JL�.^��?z�h^���;�ۚ���(G���4�~���-}V��u��.^���$��M'��`�4�w�{�w4��4޲���dD�<��2&�"��.�����YMٙ��׾z���V�r�t��eZ����Z����>����=�x�����r8��	P�i����cI�r�vW,Ȼl盁L�^��w��qVK���J��-է��9�[5m�i��l=;6ط
�q\q���iw*3<�\�ڪ���lk��\���؎.wc�����q�m�R[���v�yٞ-��u��kvۄ�H�s�wX�*��6E���\�����q���N��Ky!x�q�6=ee��ɫ��w��w���R���'7KrL��S55f��r���h^uʎ����-X��亮�M�I4Ŏa̄�����e4
�W�{�w>�����ύ�ߘ����E�*���u�)�u�,�S��?y�3��1��cDQ�RG�w_�4��Z�YM�����Iّ71�%�I��������U��>���w�Z���-����E����S@��z��s@�_U��`�C��{Q��p���<���vsiv/H��i���c=`wxGqt߾�nO�D�i���<����XN���� ���*-�����h}��k��b��! �2 2�&�~ث�?.��8�_u�s�=�=�J�*�7HڶU�<���@o�ޚ?$߾w�w_�4y�ˋ$��	��;f �k��׋�(J�_w�����H49F�F�Z�����/�r�|`���Ԗ��ڵ��Pj�i�x.:1�F쾴�ؗ��c��c[Tq�מ�;޾��}���D�h�ln�ŀ4�ـ~�|�~��Ӏ{Y�?�4���n%&h/Jo�1#��ۚ�;��=��#���,��R(�4��t�{9ף�I/���� ��"�C���$� ��-k�J&8��� �?g�4 j Ԩ� 7&q����K�7�:|�(�B(� �~T��R��,��-�2�J��HHb�!6|�0 @	�b4A�	���F*oY�1����hJFD�$IX�B���$$� I6�uCvl�ă���$�,a	�
��$�
2�)
![1$B,I��V(p���c�2��$H0Y�I�D�"�`#	pQ��"~X�łdB@�@�a�Ǣtv�D?(�|!�>8��!�M"�Cw3�vnI��/M l\|�q�`�&��Zً3���p��XOm��7� =����7��ME�{�)�}�}w�����-}V�ݝMX��M�-L��h�IR�`�,c��de�d���}���KH�ʪ��F��l/v������-}V��u��=�[.(LH�2�*����şɓ��N�� ӭs�{�+�����S#�4
�W�{�w4��Z�[��u��cőDӎ�4�s�Z���zw�ZY��)d:*��*(�a Chib�"���w7$���.9�(�JL�.W�h�n�k�h�]���Y��J5EL$J(3VU.^�Փ���\N�l�l�][��]\0�b��g0��F)��n/�{��s@��Z��s@�_U���զ��Q��,� n���kŀ4�\���,�ſ �7��ME�w_�4��Z�[��Z���5lI�	15*��`t%<��N��ŀ7Z��K9�x���S�V��Uc�����,��8�M� ӭs�4��I���h ]�T#B���f$�X��p�H���jv"�	�����
ڶ��e�%I�a�l-jոWN�l�K=�����=��ɛ�f��K	����a��M�����^�� ��:Z<�f�ɢh���E�xa�kt�����aͬ��I.�E$ƳN�x�ՠqA����Ul
kf�� hzm飲VΏrY)]���cq�\�7c�:ӄ��C��"7".r2��׽����c�'�]i��u@���h$�<�\ٗ���2i�F�v�Cy��<:�djF�rmL�L�/;V��;V�S�s�
?Hn�b�"�t]�SeU�SjH�yڴ��Z�n�U��{�GVF�"Q����\���?z�Xt(��zy�`����L�*�PiLOqh�n�U��{��r��@?˫M'�8�x'3@��z�Қ�������=��%�R�DZ�:a�r����^��ܗFz�ħe�KI��s6{-�mȑO�o{m�N��������|`u�ԊܪU`�j�M��޽&,3�@��cZ&GK ���8�������h�Jh����&F��NE�~�����h�Jh��נ>�����㖃��e�A�Y����8�0[M�����5�&�D�%U5]�@}�/M�]]���s�nh[^���L��q���"�K�\ק'k���&�N[����]�v�i�@�@ő9�n$�\�ՠ~�S@����a��Pr
)��n-���Vנwt��kV� ���q�4@X����ڴ�ajD		B�IKu-��� ��ꁃp#�dqh�)�Z�u�~nف�__t����R��UwS%L����7R�`�����>���;��h^ZF�rH������e���u۶�oMp#բ��m����F�Y��aS#M�jG�~�S@��Zw]�֭z�ұ�i�	�17��h�w4Z����߳1#���9��1H�Z���֭z!L�����u`��]9WwwR�ɶ�Rf�kV����+k�����`$v�@�
f��
i_�7���P#�Y�cJbm����M�I�wW�}� n���>Q�B�������Ev��u����ֳ�Zz�t���k��l��'��l;�ٸq��S�\�����wm�u-��/��0;�~a��	��zs�G\���`-��I|��vwT�B�bi!����?��h�� �����Z����ɊAG��Z�e4��`��p9D�\�V��˲�r�LM�@�mzwJh�դ��uٹ&#�X !�WWZMX6�"n�!T[S�5��iy ;P ��,�{x�o�����;nN�.:�ٹ�5�x}�"�e�Ͳ�R�z,KQ�x�C:D6��U���c�M��b�2��f��ejvy�=8xF-͎��9ѓf�Lm؎�3�˦̖�Pi���bZK�y�l��T6y�����ܩg�7:��Ia-�zN���s�a獁�.��8�!�:��w��W?V����U�z��z���r9��{A��TZn��t�k�������nLKs�L|����-jנ~�S@��Zw,���H�I�D�4Z�����6[u�n�>�*��"ϭR��&����iǠw��?Ɓ�����-j٠�;\nXT�"Zh?f%�?N������� �ݳ ��aɄy"M���;�S@��^���M����D�U1$���c�З95�VU�g�=�wE���7�"�vN���~�֨ԹS���ղ�ޏޚ}��9[^�wu��y��	�5ov������b�f|�K=��~��@��@��^���XE �(�6��6[u����%3�Wt��0�����s����%m�h|?�Z�e4Vנwrȝx䑬�n�����)��>�~��ǀ��� 7����I.��C����uZ�Tٴv�f�F�k��n8v궍�@��-����ɍ�6�LM���}���9^�@;����Z��u���L�xUـl�u�%27O� �}X��N:����D��Ǡw>�@������?#�����3k��1B�)|�߳/� ����)�%]��Ucm��zؖ$����@}�_���Ϫ�?+�.(LS	�x�w8��%����wW}8u-���u�TH�!hVȭnZ�m���q�ܜ��m֍΋�
��rty릭�V�Lm�@�mzs��ھ����}8�;��j䛪�UWX�k��(�2r����� ���
d��s\�"Y$m�G��|��@�l����_}��-w�~���ɍ���Jbx�\���`[u�nֹ��T�)	JoJMx��˹$�	�}n[�ɓ�<��U��Ϫ�.Wj�?[)�_>F۸���6M�$f��ږA�M��qg�n�X쒬ʜ��-�r�g�s[Xo&G�!����ߖ�r�V���O�l<��M���A�kC*u���z�v����Vנw>�@��0��1L$#Q�'"�?[)�Umz�fg�V���>ϟ�-�t��A�r�mMU��)�����Ӏ4����}�����cB��#�@�}g i�s�~nـ9z� ��,�D"�����!E�H��!!��b@�#�1���!�	!٥N:HE���0��0�$��c�"��
�C�VRbI!��`F0$*�2pT�� H�(�m�B�h"�Y͑�0a �`� '��~~�C���#�J��bF
7�"��2꣛.ѣ��	0�a!E*>T��I�$x|/1!��x�ĉ��&���O��9����Cd;kـ	�H��$f8�$�~�Ym��s/�/J�,0�Rt��KzD�ZM٧��x

��&�yd�9� q���d�c�MM�d��ٷe8v�t�p`�����ݬbŝ��k`��! �&\�**1����6`��Pp���R�m�ۯ%���,&F����UMIpgll5)J�̙K�a��lU[Js��.�W����6�BY0L�3�
q�n�v�Y �I���@�6hx�\C5&7@q�����r�]����
�*[]��m7��s6ʺEB��Z�\�sV�8N7Fhs�Z���$�;<�u�!2�����F]n3g��6�X�Y����V�.�.qΡ��v�Qڰ�R�[�4�1#!aեۇ��
R��z;h�q�k�9L%[l�8�*JT˰��rc��\�k8�Q�9�DS=���g��g���Ts`�q���6�@smB-���v퓇-!u4��P��g6l�(eʸ�c\��ζ�UV��c�̠%��2�O/l8mnL�N[Y�!�M��3�=�.8��Nyڗd�X\{W]�-��f|'
WF-����w�u� �b�ٮ�ih�f��DC�i�3�m.�UF��0�L��l�n�T"�kL��c�Z��0I=�����n���	�s���9.k�$λZ0�@�����_konMg�4bޙGHmq�vѳ�;Dg��o�,m��W*�`��i�G&��ɤ#�ëF��nR�1��x1	��X �̣� #y�p)-]+l�L�U ��,C���K,�4�ʻs���0�-��F��B Ԭ�JR�vI]�m�ʶ�P+�tr@�띸��6Nr;�Z�."1D�Ŝ�dV��s�,ٴ�3�UH	,�5���U@ JZ�*f����u��[�l�b�)�1a�NHeǪ��n7����XXx�{[vl�sm�]�vzz�C�u�,y�{g��'N#��N�M��dr�9�2*�؎CV�܇V0Jk���ۚNm�q�99&u�<�ѷZX��浗��j��L����+��px���U��?'E*0
��� � #Q"'�`!�G�*��B"gD�8]s.��j:̖Xds��O'��0�FT�B.'���-�a�2#�-ͅ,r��6�1;�	[хK��-�����5k�-�8<T�.R�<A��8"��a0ơܮ�& ���\�ε��׍��N�FC�$��N�C�n.V�`��\odf�R�5�N�k��MH
ܝQ�ӧ����(�*hN���>�x�|��o6-��f�[�]MbUqE�6o,ܶ�����]�[�v�%����ҧ��!nig'.�ԽR�����܌�gR�&>�}�-���f �뮈�� �>�y͓Y�Ɯ��jcxۋ@�l��U����h+���R�8�1�!�Uz���Z�������v�	V)Y%v��b}���ߖ���M����;ZD�S��WWs�4�\�
����t���9�ν�Y����4��ЊʬD�kE=�x(���Pcv�\�t�unx����\��	�q5��r/�{�ƁU����=	%�C�S��<���5e)�����%4_yٮ�$���x�N�ݽܮՠ~�S@��o��Дs�#�;�U�\���?[)�Uz�����F�IdQŠ\���?[)�Umzs�ף��1�1���UU���f�
:��� �>��M� ��-i2q<CDƈǄ�ʣ��gmsD��7O[���K�Q��v���$K��4
��@�}V�r������}>4�_�Lɍ�n'�����}V���M����;Z��ȝm�e�@w㷦��{zh�śC�f�E�{{�f����ܓ�ϲv�J�K%�$���I?��x�}�=��Z�e4���'��E1��uzs���h���m����~|�E���ksLC�q��5؝;������1�.�ru�+��r`��d��Ϫ�/S@�l��˭z����c$r4ȣ�@�YM�$�Ow_��X�k��e\�+sƔ��$4��h�ק�Z��@��O� ��wT�N1Gı9g[�v�� �v�҅z�D(�ŗ����8p�hTH��%Q�l�Ϫ�/S@�l��˭z���w�m*��[dz�u��6!��a�m����J�Yhh����p�n�!�uƺL2/�}O�Ɓ��M�Z���h��P��$#pQ�7���.��Ϫ�/Sٟ�����' 5��4
��=��Z}����|h���w��Lhs	#�;�U�=� �ݳ�D)t�� ����$r4ȣ�@�YM���.����h�g�UP�F�A���x�� ���wn(�u��Ъ����gqke�K��&�u�A:\�h��c��U��B˞�y-� ���un�m�8Z�v�!#�ᱠ'u�Olj u�z�,�:��ТL�h�&4�
����Ϸ��`��/2uˏd���a�,�v�qB��[n�p)��I�=s�3��b�����{[���M�%[���O��z��I$�cF��XJ�7j�i�h8pV�ۍ���Bz���n�\�2�Ĝc�t���ncXҘ�$���|h���;�U�_S@?a��(��Q���4]��Ϫ�/�)�~�S�����q��@�7��s�ǠZ��@�,����M�uz��ֱ9�&0K#�hŔ�?[)�r�@�}V�~����a ����h���7k\���p��0��"g$�Ͳ[�9MN���P�p��\PGU�.6S�׮��=��{R�hd�[\-��Uo�@�}V�|YM���pйܵFJ�K,���^�I%����� @���"hO��,,�w�S@��^���#����^���oM�����X��w�@�ߖ����<�#�kS���?[)��f�����S@?a��(��NA�X���z��s��YM������bRI$���jF\�Ѷ[��e�m�Aח�Q�&e�A�g$�&���D��s��YM����[4g��!̀��ƖH�~�e4��h�Y�wt��w�
#"�<�~�S@=~�6hT�RE ��Et�Y�&bğ'/M���4�9�W,M96�&��f��Қ�,����M��q�Ȃ70xۓ@��M�S@�l��z���gU�o7�1��Mj�u��N7��8�MR5���:ݦs5!�����m�E�[sH����o�YM�����h�)�~���ב��cJbp��e7ؐ^��Қ�p��j$��7��h�f��Қ�,����M ��[cy1B8G&��Қ�,������g�gl�������jܩ��4�G�S@�l��z��wJh�u#"H�$`���p��uѺD͸�wi�y��`*����ah�h�WD52
<�~�S@=�f��Қ�S@�Ϭ�$Ӑj&��f��Қ�,����M�v��Lh#s�94��=첚�e4޶h�U�ǎF�)��)�~�S@=�f��Қ���y��1I�C@�l��{�����@}���>ĳ;ӳQ�dUF�R�O/j�A�nF]���Pr�� ��������v:Mg�D�.�ոluZ�]N[y7W��o:0��*Ʒ5`��(�Gm	n3u��ti�e�i�;�Ƿ\�Yx���5j.OXi�sN��n��u��=�m�Ӹn��O43�!��%�o��<�"�t^����}p(7���r�]z�g�U1�nk<��roV�]l4��U���if�h�����F�� PQ�h�ڵ�'7;N+wV�z)�3�s��x!ƢR4���NC@;��h�l�=��$�H{����]���x�PN	ɠwt���e��?[)�}��{f,M�g=�5m�#j�M�>��e4޶h�)��"�d�L�8�����M ���wJh�YM�>�28�N@M�5V`�����?����?7l�;9����'�ǒ ��cq�OS�m���7GQf]�,�q�S�=��\�Kvq�&������)�~�S@=z��ꠚ�����(��?qe5fg��X��P���6�	'�ֿM ��4��o�ٙ��('21���BHh�����@�}V���oM��:v�[�Ud��M�bow����~�����������PN	ɠwt���Ŕ�?[zh�۠=��_/wL�7T�rG�9�]'.���nW��:�S��]�s���
Wl��uW$�[)�>���@n�M ���wJh�ȨY&"�<�~�S@���@��M��)�~��G��6���@�9zhjbW3����+�tI�!_�mO�D�"!���c!�I ��A�A�� �"2E���&���K��ai%�F,��	�l4D%#A� B!!		 H�B H�
��@�+B���#FZ�J�������^S���͍L_�m��p��S`�? ��u^�u�+�=\E��*�US�Ȁ��
uWZ@:�C�*�X�3�7��4>��8��ܔ��ncCNM��4�,����M ���x�dM�x�i����Ŕ�?[)���@��M�V$�1곦L�ܒg,�����WXX�_X��.`均lF��,�NN�z�o�߭��<�k�;�S@���h{
X�I�'26�9�ֽ��1"�>4q���?[)����ǃy18���@��M�YM����l�=歂�!��(ƲG�c�@�l�ܒ}��[�J)䀌6(�"�ōk31�,ߟ�� o��t�Һ�#�����M�~���l��=�:�س�ryP��6�K�%+s�m�cS���kk�A�x���_Iڥ��`��l�<��h[f��Қ��V����@q>Ȫ�VJ�$��s����)�_]t��0[w�
!BS#��dRD���)������i�(Jd}�xn��7vB�͕v]�cy$qh�^�呂_��h�)�{�uh{�%q�̍�9&�u��s�������@�{t��� ��0s
��[��L֦�]R�kQ�A��d���U��]��� Z8m��X@�(l�z�<�ِ�T��]Y��up�l=sH��ɮ2���*�iE�:e�G#��v�	�ɐ�^-� �{^Ƶcf��k�:�=����vh��-�2ة;�5��&�&���iŚ�Sҹ�{H�e��F��D69Q���}�z�U�٩��f�;�n�9�Y�9���j�1$��1�X��\�oZ�i��˙�'v�G��s;�G�᦬� b��m���/m$��o&'��x�>4u�- �m���*���G}�I�0q�d����~�� ��h�)�wtj�2b�"R&�NE���@:��}���|h~�E�~�$hn@&�uWx�/�^ ۾0k�s���@;���<�0Q9��4��>��}�s���x�]��A��?#����9�Pu��b�G��:W'*,�̜��I�+��N���v�4��(�=��� ~m� k�D(�K�n��:�'�A�F5��$�@?[f�!%
�J*í�����=�X�
��[�8�$M�9&�u�0ݶa�)�}}s����7Ah�V��������B�D*�����Z��4�Y�y�$I�0q�d��݆�~�� ��h�)�m}�DHu
�ڪ)S��� :�������K �Jv�Qk����'��{�1|a�МN<M�~ ��}4�Y�wt���a�{�+H�N@$27&�u�y�26�_vY��w�芠�?�*�늨�-����h���7�?��:"6EIf��krI�w�@s�)ε\���$
;M�;�~��{ﾚ׬�;�S@�q�X��#ɍ�C@?[f�u�4��s��4�c琛=��R���Ւs�N^KV�a����ܚ�h��9�X����J$��6�䟀/��wt���a���@<qk	�y18���wx��3�%2k�� �w^ k�7�H��?��$c�Y#�����Z��4�Y�wt����T&LX�D��rE��b^�呂_��@��ٹ4A��)�H�4��P�f,�7�}^��y{���@z��Jh�,Z}l�={~�a���)c�bHݮѬ���ZX	�D�b�Q�'\�1͎�=s�=v:jh�S@�Yb��f�u�4�k:����E�
C@�Yb��f�u�4�)�{���1�F�ɉ��]� ����w�(I)�n��5���a�ĢN1Lq�5$��f �m�����g��x�Iܪ�ES���Kn��9zh%����^�=����'���ܓ�;`!�����p$A���:�>g�����nf7��\�98ci�l�y�m95��q���q.�]-��ے�Uj��nJ\�u�`�(���0�+v-�&�jø�ۍ�z�k�p�l�@[<��a5c�����2�8�v�q�V�8���T�t@O�J[�ݹ�˝�]��H!�HS��rvNQ�).�Ŕ�N���s;��}����ű�_9IݎSRK�z�H��"���;���{�~�~4��	���QX���Ζb��i��t�Y+O��}�`�	����m�JʩWug�;���,��� 5���!�ύ֯�L��̍�G�� ���)�|��n��=���m�'"M9&�G&�u�4�)�{��4߻۠|5��UA�]CV[t��=��4�٠z��ί"rE�
C@�[���f�w[4�)�w��7s4�O�jFʎ���[q�G����֥V�/l��
��9Ռ�H�!1<��h��@;����?z��W��bQ'�8�����n���%�J��J���4�v�� w����16u�O�MU"��*�#�@���~�,Z}l����˫�����H�w��h�w�ۼ��o8�Ծ�h�*�[ �#Z}l����Jh��Ǡ=�1f/w�oM���7Un����������;r�GWV�4 �\��۞����3�H�n@i�������@��M|��{[`w���s�P��+�wL�o�tZm�@:�4�5��(�M��p�?u�- �m�?#��d$� $�B-#!aYsKL�۠>������s�Uc1<�H���hu�@��M�{�ߢ�aK�Q'�d�89&�v�xDDCo8����p�n��m���R�H��e�)� ��f�y{A��A�s�йw��-������\�t��d��;�S@��,Z��4�٠yyZ����H�~��- �on�9���s����Y�����d��P� ����{ﾚ�l�;�S@���h�J��4ېkrhsw�=�f�;u8����Z�Q,J'�w^� ���܊��P�r�y�Z�ek@/���l�?{-X#�䘃�=��B�mb��"�<b0���UK�cI,�ק4����IK��m"2������w�۾J?Hs�Ӏz�"6'2<iLl�H���oؐ_��h���?u�- ��Z"r&8�$�����Z�Š��@�[�&78A8'&�������h�l����jؑ&@nY�@���4��h[f����n䟍��mN���	�!P���sK�h��`@�sA�@�%ǎ�4�C����Ȑ F@�"���0c��&�����VE
]�BHĒDY!# a!&���A$����5�To���8��9	6 �Hr$%^�0I��� ��VHA-!��� HdBC�y���t�F�@��d���#ac�e"�,"��B0�f�R�~�LӅ��b9y�����9��'GŊ�n�1�kp�t�c���l��۬� i�����Ӧt��͍���>˥�ݛX����e��jWm�� �HaBP9A,p�؁)&8����A�PR��洫+̤�i�k:��k���PNΊtU@�AB���G)�v�m�p�ձ�Z�c`[EC���ګq��=+�m����q#�e��A� x��e���v�������(/�鶮�5q�ϷU��촲��j�j�0���θão�]$ؓ�L�ny�sׅd�&�Lf�ţ�-ڴ/h��IV��Π\ci,�9ڠu�*	�ʄ�{i5�f��b��]]
i ;���G@�C�Aݙ:܆g�=-�Ʊ��;l��:��l�0��	Z5��6r��A����$+�;����*�c��j�2uFJ����V�x����ZL��[; �-�����QJ�b���T�ژqq�����=��)\Q����S�̝��l��uC�@7/�d,z��6�j7Qƻ [y�8��[����n0�Kt��;A�i���1�Yl՝�`��m��e���\ur�[@:��WaۨA�����`"�: j��zXe�'�A4�v\�1o5�[��6(�0��YN4��0�U��b���5��EtqY8����ʍ�9;��ў�+s˘/&�qn�ƘC6�enT
����u�S��hn��Q���n{4��� ���D(&U�R@h
/$A�"8� øض�zr�Se�j���8�j0*����Glpr��6Ů��:��9o4�ٸd4g]$�jM.v�X+�l_|�W}�J5T����u��U[ �UKm�Q�@��k�SlIk=:*d3O<2uq�nh7����\��𑗫Fh�p���g݂��]�ˍ�;��Ĺ���"����HNP�j��R`�ܺenv�����d�K��:Xc*�˻\M�nz[sF���K�sYMd�f��N�)�@8(~6������,1�]���U��^$Cj?���6��o5��s&h�.�mz�㧘��qϷ����66�K��mx�zipi�������c�i������&Ɋ݈��D�V�`�uuZ�GGdILk�����	���=}n]��uŭ`��+�G`�aݴ�5)�si��8��)y1�z�\��䇵�Q^un�@��i�x)���:����7N^�N���=��s(�������v�,�\Qt�Ȇ�\�yq~]�[�S5f�k30�@c�c8z�ՂW�^s]��
P�����D��1�liH��b��8�nC�>�}4��@�}V����h�J��4���ܚ�٠w>�@��X���g�%2IO��(	��J����|���� �m��٠w���ds$!l!Z�Š�� �l�/>�@��dN�'21���RF����9%-�_�9���=�n� ��Þ�D'b�6К�B��غ8�s��GX�r=�*�3�w!�l=�ɡ�u��T�@;����h��� ��h��ޫBJR�Q�ty9ׯf-�P�Ua$FE��D�	��J�O��^�hu�~����"L���Y�@�}>�@?[f�w[4��h�]P��&5<�h����w�nֹ��P����8�����4���ܚ�٠r��@��X�׬�9g���'�#ɏ�L.��p�j{l[�g8��C�lM��=ڸ�wi�:O����,mɠr��@���4�]�H�� z�O�]�R�ꪐ]��`���9$�"&Cy�����8��f��,M��Z�zAʬ#U8[-0y����JTt�S.B��×ߵ��}��a�DRD�B6���٠r��@�[��^�@�[�p#��rh�k�>��}���>��m��t��`�ci���1t���\ue���u�#j����3���m�"�$���
1��@�[���f�u�hzנw��c�I�ヌ�h�@;��^��������!#M9�&�G&�w[4
�k�=�+Z{��?.Ë��@���Z���QսՀn��N =��r|�������S�*�M�ĺ������Qv+S�l� �Z�޲Š�� �hzנUn��Jݘ�ր���X�u�q��/�od�� �^Ywa�G#.�'\:��^�4�٠U�^���X��_s���[V�Ic����n��g�}��=�O��^�@�[�`�����/Z�޲ŧٙ���h�}4/WX�L��%�Ǡ~��- ��4�٠r��@���c�ȱ�ǃ�- ��4�٠r�������fffs�R$M9�l��\lS�헣k5�����M�v�BPaَ���@�,�ktv6�����p�������v 6���٣g����h�7V����5	p���]�*���X�K-fX0�OF�u:��#�\��'nɜ����^�]ki.{�8���W�P�m�
�����{p�'��T��+���snم'u�h�a�盍rk!����{��wws�}�]��@��6z���a}cӑ��Hu��Q��Vw��x�j5�!��k#rh�}4^���e�@=z�����p D��*���6|�gСL�޾��o� 5��yf$�=�)�5J�Kd�-���}>k@/u��٠U�^���vA��&'�� ��h[f�W�f�ىc�=�G�!s�l��ڶ�jI�m�^�����^�4�`��E&�ũ57�M'�;J6��๭�#kqRח��Gn����ʒD8�;n�87'�>]��@��X��Y�m����y'���K��?u�-k��z����x�n�>n�z�n$ɒd�88�rE��� �l��%���ޚ���� s�s�)X;Uj,Qɠm�^�����^�4�Ë��@#s�94
�k�>���}�E��~��l�?sXp�m����71����r��7	�X�E��"��ۧY��OnX�\��{ji�m���+�^�4����.��wUH72b�LL�H��Y����Z�޲Š�=�")"Y$M�ԓI'�w�ܓ��{��M��#��Gň^�נ����;�j$UI'��*��@��,Z{�����?��女�?��8@PQ�`�z�Yb��f�u�hzנ~�d0l���՞�<�#͢���u�Q7T��H"�B�⣳4�h�{i�:���ٞ�F =�x������(�!���8�vz�*j�Qi�n�9����3G˾����h�@�ϒE���b�ܚ^���e�@/u��w�@w�)εjs%�@V�f��f,���u� s}x���5DBV�Z�Q4E!�x���w�ܓ�vj��35�2bd�E��� �hzנ~��- �1"��D�ȰI��
Nx#�3�]�[F��a�=2/�Ӌyƚ!���өQqM(ԓ@;��^���e�@/u�#�[�`�LmŃ�9��7X�;w8 �]���ΈQ2w�_�8@DQ	`�z���Z{��;���*��@��Css8H�rE��f��n��ֽ��?����- ����70j,�ɠw[� �[�_����� y��Q
."#8�����A�dU��Wh7�g"Q4���M�U�Bu��z
����l����m�]���8�\��ݤг,�i)c����$ӈ��:l��n�Cb�3��7� ][t���c�;����kt������y�	�A���m/nǷ\����Nb�����rԤk&m���mJEk8��lH�L�)ihz���qp۵��1n�g��3�{�׽������N7����/Z!�����g��il;b�E���[�N��0��׫��&bmɞ��^���X�׬�;���;�>�$���m<2G#�?z��z��u��/Z���"u�ncLɉ�I�z��u��/Z�޲Š�=�"(�28�PrM��f�W}��?z��z���X[�`�LMǃ�9���Z�Yb���@�����)�vUc"u����#Cb�j8I�x�ͣNgus��?���;��C@g��M���^�ѐ߻�������@����N`�Ǌ<��'>�u������Ae���6nI�Nu������`��g�R���Ց�4�}��{�U�~�]��~�f���$��&ě�4s���`�n�:)���`B��+.�T�<?�qh��a��٠{���=Ϫ�?{���1�&?�RF	��i��[q����)h�j�]�&����3�9Ս��+s�d����~�f��s@�>����=�톀{���J(���jI�{���=_U�~�]��w����Ŗ9���[��Z��u����5��Ņ>"� ��T�I�&А!G6 l���+�"bA$$Aޒ�R0"��! ��&�ApB��kh ��	@$Ӥ	�a���D�@%�Mǂ�,b�`@,�
t*�
�:a�"a�4������!�b@��`FF�H�a#2@���XA��K� �8D�W ��fj	F,ށ���d$u��4���G����j��?,:�E�B @#1��`B�FB,��!�@�(}\b,,�H�b�H�c&��T8�T�2(�D�P~W:��*iUN�-�v~P�Q6��~� v��)��?/8 m��S�ޥ���rN}�vnI�c\�m;UN���נ�O�wۦ��^��f(��;��p�s\�jФǊ<����@�t��������;�	D���0R28.m��څ-�����OF�K���6����q>Y��0Ȝ��X��@�t�������uO%�`}�z��:�~�Q vTܒf��}V���v�������1"�5~y��<?�qh���@;�����������̘��Muv`���7[ŀyֹ�"���J�"H�)$1c H7�P�$2� ib#	��7��G��%���l4��_��E�c�I4��`u�p�o,��w�rIk]ߪ�h'e�u�=�ۙ�d�7h�]��w<t c�`�-���{M�z��g�����p�o,��w���ŀo�]�m;UN���נ7�{�k٘�Ă��M߾��=_U�wtN�N`���܆�w��[w4W�h�{�h}�g`)PUc�;-�yb�}��`��p��Y��� ���8���0snL�=_U�~�� �����{��1oČK1,��b�C�HD�����lw�-Å�0��N�6�6Ta�غn�'v���l)UnK��֞�!�̀W$�֍��T��1��V�x���yS@sH66.6�n��qp�m�=i�Z��xi1Q����ez�s\K����
��$ʲ�*HnJ\	��ݠ5�Rs\p̿毹��lf0=�#��iKKo�l�v��AV�*�����,K�|�Y��+��=���Y�ݙ�B�m�K��u�#x�0Z7#=!u�Zc�Ƹ{<]�
zӷ4�ަZ{�޶h��h���?{�'\�1c&&H�4�l�;���>��^���ؖ&��/w���A71��h���������h�h�u�����	��=Ϫ�?z݆�~�f��n��k:ıI�����@��v���u����ZXy,H�n!�SHL����X��Y�wEp�%��n�p%7=�l�ZF�l�ı�G�r���u����Z�[����Pc�s#QdnM$���f�< �J+��y33���~���4�w�@m���ܵeNIj�Ϫ�?z݆�~�������:�d`�F��ӏ@��v�[4�w4/Z������Lxɉ�;� =�� �o��u�~�yf��w�����v4$�I&�hMh�WG7<h�۱�u΍�ۯ1�@Y���a܆�=�`�V��6�䟀-��yzנ~�� ����A�s�bc�pNM�ֽ���h�l��f��1��bs"v��u�f�����n��3�B�x)c���*?���#�#=��t�����+�Mʭ��)k�� ����l�<�k�?z݆�g�vI�)�M �h(P���~�ݖ`�7x��\��<s�]uH=�z�n:���R-��u%� �=nwH�-���X;*jIn���ν���h�[4�٠_cY��#4��z�[��޶hu�@��W�{܈�pNdǌ��#��޶h[f���@���4�e�(� csQ�&�u�h^���n�7  nb�z�!/��l�+G0o&&H��rh^����Y������ �y�RTt�� 1�8Y!����@�H��:܉���vl�\]��:���p��qbrEO�m�ݖ`�7x���I~���Հk��ؔ�#�c���4����٠z}����Y�	(IL���] ��
L�x��@/�}4/uz[.��۠��R�Q@vT��<�c����/}��@?z٠m���ᑃ	�cN=�n�@?z٠[���u�JI'I"��D Y�~�߿}��Ә΄���h��c�T��X��ul�f����Қ��gd�Bތ�:Nd�&J�ON,�lk��	�駌:��K��F��b�Vn�\*e�%ۇ��9�]']E����ZnH��Ӹ��r����[m�,�ړmث���P�U�I��z���8�m]}�Y�$�d���=���<�U��n��⶗.��I7(7�߽���>�w�ￊ��5<f�b��;V:5r�͎ú����c=H2����wa�FFl7\�LN(�? u呂u�h^����� ����S9�jI�m�����n�@?z٠�QLɉ�!��4/uz�a��l��f��e��2b��j)#�?z݆�~��@;�������wsq�p��܆�~��@;��������S@~IfqE�zC�rYm�#���GN�ܢ�.���a�\��s��6Ӵ�ۛ��+�o"��d$c�O����<�����Y��@��^ F�Mt]��f�E�f��'�������?.��ޅ7F��	J��?DB�?s�0ݮ�u��/�gW�H��q��n�@?z٠����^��r"u�9�2cy#��޶hu�@��W�~�� �����X�F�jI�����^����4����	�N�'�l|=L��=Om"Nn�����]�l��u��&1̎`dN	��LLq	��]~z�[��޶hu�@��%�1̘�(���=���h�[4�٠y{��;�'q'1��	�h���nI>����@:@B?4b���W)(�Jr�_� ���06�9��d$c�M �h^��޷a��l�����I��(ܚ�k��o(�ͻ��� �""#����y��૨b(:�\[ۑ�ۧ�i��k4A��`h��p��=�ͺ睩_�&��w�k4��hu�@�}V��r"u�9�8��f�~�� �h]����� �)kQ'�c�q�&�w[4.��޷a��٠g.�x7�C�rh}����Հ{{�� ������RI(�D �aD�T�X5R���w�7ӝԴ��S����l��yf ~�� 7[�Ӻ� �Jk>������l�kr�fwc=t'1�f����Qk�"ݵ�89��F�nJ^mN�~ �����˺����h�;XR���V�e� �;ۯ,I$r��{��E��٠;9;��	�AF��<���?z��~�f�s�����eS"�<����I?���- ���@;���Z�{��UTP�Em���w�@?fbS����'׾��o�k�]�?�@_���*��A@_�"�*�U��PW��@_�"�*����#�� �B
�F
� �D"�D *�� *
�H*� �� �� �AU
�T
�A��`�A�*`�F
� �F
�`�D��"�DX*R
��� �DH*F
� ��"�E�`�E
�X*U*D
�F*�TH*��H*X*`�E��B*���
�P��X*X*�"���
�`�F
�
�A��E ��*@��H*U��V�
�D� �A@��AD�� B
�QH*H��U
�EA��DH*V���**�T��A �E���
�b
���",b�H
�X*���*��B
�
�H
�P
�D ��EU �D��A
�A����@"�A��D`�@H
�@��b*�� B�*R� �EH���� *V
� *E��A
�E * �A��AV*� *V� �@
�"� * *`�D��Eb*V
� ��B� **� *��2"�
T ?�� ���U�tPWȠ
���(�� U�U��PW��@_�E U�U�PPW�(����
�2�ή�� �>�����9�>���g�4h()Bm�P �( ��t h��P	D� �١@   
�W�)JD*TP�J�I Q
�	*(������BP(�"�(�H�Q*��TUJAT!J���( 0    ` 4     � zR�﷫x�y�;/mq��g��
�������j�s�����R� >��)g���x�� �o;u^O.�ˀ �}zѹ��Y���-z�W��:�����r˖�mT�5h ǥ P   A@�` 7�K-u����{7�� �h^�� ��V-2�C,}-��F��<�ͼ_my�x �}�ﶪ�ݰp ���u�j��ݱ\�r��׶���{�e��e���ڸ���[^x @�   � )�}�w׽��N�)e��,�� ��LMOGt��YJP0=��
Y�l  
1�(M((0A����)wnR�3JK0=t ,�)KݹA@���f�QK,�)@ `�  $   8@�i�J �)K1���n��}��}��.� �R�|�/��5+�� m�����t���x�=��O�˾��� ��mͽj\�ק^m�mN�<>���>��msr�{�}���s���}   ��   @t����YW6�뗘o{�﻾������VmJe�o]�ͺ�ۼ�ҷ �Vm������  ��y�e�w�u�{�>���f����{{y�z��^� �sK�����y�y��}�S弟]��  i�
��J�A�F�"��2����   ���R��&iCF ��U*&   ��$��)H  A1J�H�c��Ǐ��L�������vw�W�;��AU�g�\�����A_�PU�"��PQT�����B�4e?�����7�)��?����G�Z���n��t/o��}YcNV������ev�Q��e�|1,�3w��w��:�E�c��7y�Js������>FAh��r�޲�w��!��;�kH��b�"q% �% }��Mp�a`B�bF��P�rc3n!B@���X��b�.�c�o?&>2�	
��_X'�o�]нWD��u�Ҡ�*�u
D�.��δ��\�*bbH���>�� �w�~�pwg�֘T�b�Ɣ�xK���!����W4-�#���p��b�u�J�ԒQ�Lf����Ƙ�)�0!R����h�Ǝ ��$p���ɘ�1H�W)���rK�m�s#��4���	�&� K��kl��)�O�h1�yG(	���y�߸�;#�I

Ɓ
h�d"�1�S�D6p��F,�G��d����9��>Č
$j�S��pΰl1�\\d�0��Y~���# 0q ���'��4M��f�h�"��� Pf ��M�%0[Ki���
F�BH%� I�ĉ!#��2	Gܩ�ߗ��.��qZs&7��V0��T� �	 �ͩ��.s)p�%%3���(�ޙM�cA��F!q���7��F(�+���(��/���
N������W�Z��U?���?g�s����q\Q"~���t����=�4����_�to�߃��2��@�]�$ά:94.$�k�0r�%q�v�BJH̊$�i# I�&3��L�F/�4��f3� �T������ː��b14&)|0�m�:��!6d���g��l�̉>�7����r`0!�$P%��	W�*��UL��M~)*ym�j��4�s�*� �	"�q��/�l�)|fs)��P�H��Xݳ�IM�����2�Fw���˓' �Ł���as��Sy��q�2���L	u�Hoy4o=��c��cHH��d�@�L7�	�؏.��A��r�N�BK��0F��H�ap@�ɢ\f]���4>�!T�Յ�!LF�aL,��B`�
G���$�J��%b@$IMB�0��4�u�$�C`HH| gƿ���[�(��fmw�:�.*��Aw��1U���.$X�*S�S��i���:����w�!�Z�@���%MЁ6�I1��#�~�E~3��*��:�.̗P�8�]d�Y	���B!w!1�B@�35
ċa"Ԥ�R1�>��N���"I>�}~�|�oni��h�z��H�~#A"E�� @�!Y�!XQ��y��K�#!�^g�.�40@��P�tƌɀ!d2C9��L��"�l#���1Ip�zbM��
1�egZ	q�I�}��È�#��B�ad��dr\⒔�e�_z�j�����I;�IK�#6�H�$�\
JB����7;�ֲ��jd���D����n�'��EӸ+�$.`!�aK�<2a[U
)iRM���H ��B$2�o#	q>	Le�"����k����4эU��@��Q�Cjbd0����(K(�J�!�S���Bg)���l��Y��B,8}�k�IӐ�ƙs"f�Z2�.	�'qdlٕ��@��.;W$H��BR�2��&�tsx�$5H�X���8�2$1D!���r�Y0B��(bBF4$tf�sy�A�@�b��$cF0�����i�7#̆���0e�$f\i�5\H���CϏ�J[��$�R1�~��3z�f>w�8��
$(H1$I$F8�C�7�ؼ�9��@�|��oL5&��M��^nm#�c>�L&CS��/��yk(�	�v�Ȇ�bC�m1��2ڸZM�J�c�J�����D�R%B�`���{�f�n�p�bB���+Ɍ�e�U'�<���u/�&�CStN��&��ص 4��`�GpLH�2���^����<������Umz�Ϩ��%0�9��.p�0�*JB���1	�Q�P�0�����)�� j\H�N$1M�X�1�� ��1$���3� @�����&8FL!Y�����)�`&9"���,�"n]u�i!C�HX�f0�T����7��t���@�&���#�C�����._ܱL����l0h	X41�T��L$��dH- �
JB�IpI2�2$VT��VV2�0�aB0J1�#.	5�0���^�������NV�r�ζM���H�B���0(F�U�c�(`�I �	�gY��p"I�Ĭj@�RL\{Q��V�%��ߐ�K�ӕ��i8�$HF�,����$$a	$�� J`��p��
H2���f6�(D��$H��'Ʊ�X23���#1����{�a�$`��\�BS<�\0�$6Sr�	�k͑��g����`q�\@�7j8XP�3�/��)J�������� F$��1�1����j�|�V���R��~TX,�)�HIIr�T>἗3)��S1	I�E�ľ���9Q���Wy��SD�X!$e��!	�q��"�q������Uyb]��HHɈI(�(E���F�0���$9�٬!�@�c{%�eae2)cH�J0��	`��ذ"@���B@��H� bI� 1��$��!������~`\�S�h+����"�R,!HSdگy�%������6G�34g�ĳz���\']\���-��4&:)n�Y�j�׏>�`4I&)�6~�g��|z�����~&ICR�$$�&�7s�;ÉBƐ�,)�p�G?w�
8�HQ�	L��3�\9`�02�a�.�L��+��k�cB4�K�	a��.3$ƾO��>��a�H��FSL;
4cI"%t�4	`���#�8YF!L�BĪH�u���B"R-t�S A�$����B�#\! � aaT�D�Ƙ�H%���&;��BC!���B)��p@��
�$ �"0��q�$�3��)�"U�
�@B��u��f�¿Jc_�'�@:$�2�YRg��|�����*E�lR�c$�`@�!�XũΘ��2"�ԛ:.�����!	$� �$, �fXb���\339�2K$k,d�ll�a�HHT<CE�+�@��b�\��S�mt��Ǖ}��WW��%v�%���	��͕�J\8*P��,)bIVL3�X\��$	�$!Ě�acm�."�B�*'�Oa�VVV\R��bBBHĐ�l�Nar���B�cb�1"@�B��1)$�ckIJC&�L��.p�1����#\H�>�8\���4��l,$,�!1 ���!
�BJ�b\2�%�.#C!2ļ��Ò��0d��.Z�5��{�� Lk|�Ļ�0�NW��F��]9�Lb�컊�ĸ"�f������^�JA�v�	\R4��'�ae�Be�i
$HJl%	��HI�k"��ЦR��H�	
aP� ��F%H�"Q�E$���V%�F���@ �� �̸΂c&���*`2B��$"���'�H�c �#	�a$�l����
�q\�$HNl�*c$!,`1H,R�H��JaR�M}��e˘�ØS)�7
��.2h���4�
�cY!L�.s�}�;����?Mp�с,B ŉXHŊ"��K���4�@�2�"@"F4�e��P0��L�,�� P�0�B�(J0��pk�WK���bH��lH��!A�!>��eX0`&0,X0�A�X2b:6q�M$�!V$cq���
���Yu�m���B�e@��NG�
L
D�H2BR��`�d+
B�*BD����pA���� �����!�,X�
R� [$c$����Y��	%@$B	 � �H�F"���pU�Χ�K�r�JgRÕ����X_��g�0��� ��ᨨ����jS�<X��HB�'8��#�3�_�e�<0��!aX���pK�%�*\�nd�5���A���p�K "E1�.u�B��s�����;X,2�T�0`�ˮI����B� �ԁ�K1��e�ʜHQ)D_�m
$#��q�Dse�Zt�P"LS8%!I�c:�  ���`  #m�E�P ���.A�9�[Omz�ڶY�Wog�pl�Ͳ�tq�J���룃���	tۍٟ5֡�n�U�^4,�
�U'�u����t�&�� X�7MG[mk,��r	ɸ.k:�,�Fn�Y�bͮyD,v��$�0�e�%��Y��X�fA�̭UE�b�V6r��T�Z��j�U�
VhͰČ�e�HZb�nƵ��u�뭂�	�@l����Z�u*��Z�Z�壍�C�T��9Pz�ٛU: ��8�m�R��R�@��hն���'2ʴ� ����l�m>�c"�+���<�e@�kh�Ie��6Ͱ  m���h6� �!6���` 5�Li�6�4T�)�- �	- �e�M�L�  ��ڶ��� Z���nm�� 8N�"N:,�m�d$�b��n�T�\�'M��),�d� -i�m�ڀ��[����W��40�:h�� �i � h�� l�M'm��[u�dA�^��k@ m��   -�]���a�f�Z�$	V�IN����v�赝m6�j�L ��ڶc�� ��� v���А6�,R�i��RY��5l���G��a"F�p	 �f�۶^� �`h Zrִٴ�m��Pl�f���I[Vm"o*�T�mU.Y�r�fj�<�; @U�@ 6�� �aώ>� X`	�zӀ   [�"d�
��I�mU��r�pU�����6��� d.�����mzې&������r���T�r� ?h��巀[B�*�Ft2��qr��h�����Ÿ.lG'2�F��.�f�c��<��*Ʀ�e��=Y����N�Fx��tW�q���gm�&ӧ�悶�.���%w#���n����y'D�讖�ۂ:���h�$l��H����h6��$ж�UR��i�b��T3��������۶�P�7VH6��n���l�  v���N�օ�$��mCi4�K�� hO��|�m�$m�X��@ /���m%�rF��2ۍ�`�'Ѷml   �n	Ѷ� �cm� m�h�[UJ� e@�]C'K&�mn���   6�0K��v�f� m�%�I�큶�  m��검3n�m]�ܹ����U�5WW3�6���w/rn&V�H�:*��yeiZ0U���5���niM��QbO;q"u�AvUn�:��mʗ��R���ɖ6�lT�]'a�q����rnf��t�0h׍�:@��9*���l�����lG'����.��m�o)�*�j��悬TOʀ�G���*�:&�S�,eAG+UR�ڛ���U�!5�)tPz��\	#�٨���������m��m��V��@+:�ҷ/n��MJ�Lҵ�)-��R�;R���T��].Q�&��^d&E��m2�JH2�8d�[�n������H6�'@�6�H�P��x��N5�H�ʻUR���2��T��nI��J�^�� HI)m�=+m�� p^�ݢ�e����` �` H ������In��m�2}�D�$M��[@ �m� �#���PK�qYKt��e�& �s� ����Ƙ� �ݭ��V�ҭ ���`H.���v�
m���M�'6fXʳ����[H�x��)�"� �[��(�壏$ZF�.��˻l=R�l�&�x�y{Z�n��Q�Ϳ��m�j�GnF4j��������-�,���%ls�8M#�o	}s5N�k���v� 9m6FD�U\�Ѵ�zr�� �NŕU^`8
�I�Z�D� %��X�}z����lUW_Tq�;�ղ�1[O2�I���;l2��h�@m��e�iװ֜Wa`kl�	�w]J�Ұm�Ҥ�6��Ͱ8  z9z�[` -�mm����b���US- ��R� RöZ�j��* [@-���q�H �F|��5�;m�!��	:�Hq�Ͷ8 ��@[@@ms2�R�9��v���{`�)����R�+Ui�d�ڛvi鄀W-T�@ҭ\������g $�Y��&]{^� 4-����	  p�6ؐ�`6�5[V��b�ق�A���t�	/Z V�h6ٻl6�@ ڶm&��6� $��   �5�^���[#v��m�j��UJ�A�J�Rd@����[%!"n� ���@CZm�� rm�d�)ӷ4�T�Ԥ�˲�uUN4�@U���m�84�l�A��:��U�ޖ\&FH��vێ8�tͳ�8�N�[Uڐ�ڀUU띙�$��[dmӒJi�N�E�m�8�`$	-�B��+�>u���7����ζ� [Pi�RKF�� �����i���=cf��	q��i�I[a �p,��n������n
��U]N�D�ʵ��շ��s��n���0��nql�����EG6[��*����WU竌9����Q������+�hi�F(�,�V$۶�K&��&� U\ŕ�(\�<�H5�~..��q(�5qU�5��҃Ř3�@��*M�����F��d��m�xm�\�	�H���){Y.��Zm�p  � �i�f��"��H�H`��nH9%�4����e�m� }��}m�  l�@ �Y�l�m���Sm��e�Mm��J�  ��6{[8�c�5 <��
��p�k�uQ��Æ�;=7l���k�d=5Patܺ��\��٬�n�ss�/�ȭ�KV1pXʹf;#ke�+U^����1Ĭ@U�q*��H�]������U@�]n�M�FӔ�U몾��~�U���� E[X�&�Ƌ\����\�t���$iЇ-�8���t�	��n[H�z\�5UU+�WI��.I/�E���[p�v�N$Im
V��ͺ@ t�ඒ++��i�Cj�+mt�)8p�8-j�8)�8�v�����ة`UTk;v��d��'�U��i],��P��J�ĵ*ͪe]����R�UUZk"�Ѱ�t�U �UPPT^ Q� ��	޶�	�_c��I��D�%ݵ�p %� �e^ 7KDs]�̌�%��U�yj�h��ev�[�
���սv�k49z����-�iT	�@@�T����[@psmm���m�&�al@�r�;�v��i������d)\�j�eZ����� ��n�,$]�ڠ*�����lv����v��6%ۤ��)�Vk�8ggH[d^�-��b"�%�  [@ %%����85p�	vTci0�Ć�>����˻P:��㡳�9r�o9����X�u��6�X���LlE�G������#ar�ù�m[�Uka��\�'A��u<�J�w���˶�hc^�`�6�֠j�8r-9�J�UR{w3����/;-�@W�Z�j��`A�Ch vݑ����pHe��V�X��;L�[J�`���)M���3A�8�l�E�N��H۲֐�j�l��@�ۃu>�n�F�lIӮˀ6�   ;nٶ�   6��ڮl�di��+�� ʝ��Y:9�bn�K���,����^H��h�%Rmem�U��KStu� Aw��aՓh���*�V���l�CnX붕������MH�\��e_W2�v�9$p���[v�bL�l�,HV��HN����-����ߛo�ȃ [C��-�	 �[m-� t5��m�F��n�Kh l   ѭ�٤�+�{"Lt��U*��p�� `�:*�6����ܷii��*��UV�j���R�ڷk���;K[[nHpq'm��[%�v�p�	з�걼8H��gZ����oj�Sμ�m�����V�PR�K��@.)j��
�:�
S�����8�vmL�ղ��(�Ul�`8F�nx׷2��_Ix�Z��t�+lU�,=�Bvxv6vM�+Ү�9��xW�{kiVm�U�l�:�xi-t��J��@PKT�S�����6�m$��rGHI!�p $7E[I;e8*�U���f�j�
�a��V�����v���U����;� ��     	9"۶�p   l�l�ꚛ�� 5�e�pm�l��v���l+� H ��Ñ`m�d�N���Xg��K(�U�$� �h    ڑ�i7m�mkYm[D�m$��a'm�rj�5�h�A��-�imm���oR�M� $ ���t^�ZL�Z�J�m� mH۳<;n�t 9�nݩ[H=��-@]UVԫҬU@j�j�� ��<�K��@P��� 8m�m��H����m n�e��R� �$m�� �D�ۛya�� �km��:X�t����	�ݬC�1ONi����FK%�ޠ�i����m����� ��6��H%�@l -�t.� �@��/ �`  m�� ���� hz����  ����  m&��H��R�l�m�i5��h���B� ٶ���b@�Y�  q Mk	ll�D�8M�]�;[��6�p��m�qm1���*
*�Ȫ~V&@��H���*��TEI	r#�_#"l4�"� r��� n�D�UO�B�
�]sA�	���TM ҮA�b�6��$�DWT"(;A���@����mE�"Dɬ�R��G'N!*M�
8t.���\�Ąa ���z'�U@�P�(���D\|Sa�_�W��
�����p!!���!�(A���DCA� CBu�k�������`�C��j
u��h��pA��pb��x逩�L��x���8 !�jaj���@��"�8h!�v|	�T89�|���x�r�N1��P��� Pڄ_�@60�].r�eGGˎ)i!�E`X $X<O���k ����<G�$��@i6+�S��:�:Ȃ)�I��-W��E �W*hqN*uD��*�H��R�.�$�>�4qj��Sd�B	�2L ʌ�C�#�$F��E$ �zPbh ?�	 D���
|�!DL�"�^"e@6aWf@ �*qM��^��H@<�R(��"��#DRZ��G�@%aAD�)@ ��T��������#��h
���r��p��+���Z6��E��۰L	���yb�Ѯ��5g�E�m�'s��dV�nA���v�Sj��X��m���y	��^LF��������< �A[p����*�&�m=k�ɂշ�	7jt�B�M����YXT�6^�"�U�s��ԛ�ٌILv�.����.q�S�vۮNbkf���\��&JX�0Zx��f��N�@�v�L�T"�ȴd���kՂ@t�̛q$+@��p�[Z%�{���!ÇeW7;Vj7X-v�;�me�%6�]�]�{wm�ѷK{;��rY<^L闌m�'Mp@�t�'FqkK���� 4�qa�%4�JHN`yZ�M�y���[�۴f�ِ�;��ڶ7Z�l����4=�{Xݍiq��NM��\ь�.� hp�+�B\�1]��p�:��;�n��lp���&բ���g���*��e��j�p����:�B�Xۆ���C]��8�sMv���8��1]�3�dчpێnκw6M��5��6��/S�!�չ+(���q��'6�$�# �;l���j�ӻS��u<���Vq̳բ��vM��2G,&sY=&ܞN�u���N��x��bT��3nڅ��W(��2i�Qh%�My�u[I6��h+F�m��)�0R������'s��,�	KOKU��j�eg�[^�ҳ�i}�ZE�����a�[��3�,L<؍��y�R�ӰE�dRm�=&�p��<)DZ�Qc$�R��{kI.h����5��g���]s��[�sr�k��3 $���8*9���A�H��Ąc\���%��$��`6���/�۬�'+�n�p��eQ�9蛮 6��k���)v Z�VIi��.*.�e�F����Օ�m��q m�iyM1<��5+�6rd6��:�e���b�fHݺk�ư��`9�*���8 ��6�j�ɱ	�]b<u��U���Ͻ���<(���d*�m��C� ��W*u�1`p�@�i�{��{�{���>ͥ1hl{ivi��U��St!��2�����_� ���ٸ5��k
��6шz���5�C�Jb���F���m��È�>��@�J�����K&1u�v���ͶZv�mb�W��ۅ�ݠ��m!��&�A��á<u�۱i�hg��jz����Yz9��	�[&6���m6��Bs�:�x}�l�<Ϋ/a�^�=�>�z�ݾLq�܎U8�NC�����퇹\v�	����S��3�����=�06�� n�/���'�}��I�D�m�,��}��| �0=�06H遽ҙ�(��@����"`ztt��#�nt|�Χ���9eMJ����p�:`v�K`�&�K(R�.ե�XZX���GL��l�D���� ���O�ע�:U*��q��K��*og�wk���]�Rg˲F�m�=wWiۛ_%�)]�,IW������ӣ��0*�Vd�a�ʳ����\�酙�$W �$F+RBR�~J�y�b�?6�`���ײ�|���1#%�����d�\=���پ| ��� �v���Q�ebYw��$t��gK`�&����|�}��I��m�,��}��x����^,��,�J�W=<�����h���C�kE��bb�]��nL��NLۇZ�qu�ݰv�km�G�$��0=�06H��Ζ�ٝdJ�WY�� ���$t��gu��ݼ�ēgz���"Gc��2�8ɩ'=�hԓ|�;u8�9�D`�H�X�J)	(P��B���{���B����1e+�ŉ*`{�������d��u���²b��e%l�D��tt��#�nt�+�A��v�,J�Gʤ$�ͪ��rݤ\�״[4��V��BB[o=up�K�M�(*J�����x�������l�D��&+I
��YX�]��?�f̟��I��`{�:`l�Y$�D�m�,��}��| �wo�
g���݋ �u�*�Es�W�[ �0=�06H��U[�ȳS���������#�T���=�06H��t��.T�v.����ӑ{k��I�n�rv��;vq������9��v\�j�]���vRJ�q�2��v,�v� �n��"��b�;�"���Y,U�,����Ӏ쉁���d��u��ϰɊ�L՘�����a�D��v,���u��7+%�R�l��<�Ğ�����߿:`zE�"`m쫘�*J�1YX�]��0="� �2Ns�ѩ&RPg��x����?5��'b%�My��<Ŭ�mr�������j3�gHr�'>9v�����j)+&cWO.���Y��6�4��Fv({p�k�%vHfp ukd; ��J���1<�v��XN��Gv�Ѹ�鶓yj�vw�:Pv]w����=�:�;N�)�׭��[��Hl����vx~���Tlާq̚:����
�mmg�/m�����F>���_�q��>պS�=<�w7@^���va�ڭ۴\\r�;q9�E�=lu�G-ln6�r�U�7�����D���遲GL�
hW�+�@"j� �n��#o�`�ذ��0NW����-*V	$���遽#��P`�&���W(̵����M�Z�舄�S����>�0�n� ,.|�R��ZJ��A�oH��07�t��Ur�%�����/6��u��*U�n��X5G,K���J�q�l���6���X���`m��5�^������%
� }�׀k��*�K@���+����s�Y��!	 HO [�0��F�ЄM$T(
����oذ�w��v^������)$�R�ܫ�v��zH�t���0;ye�=�M��;����$���^ n��07z:`v�遽 �j�/��-bL�LLގ��:`��<���n���Be�j�`KNɅM��<�q0)�k+����sճ�FY�/)]�*�b������#��0�-p�u��D��mBi�*�����l��oIi�����u,.|�*�+�� }�v��w]ᘸa���j���[��X=�XҶbZUNnAY���LzKLގ��:`��ed�]�@%j�,V��0;dt�=�&�&&]�+1]լ�
g�gɯ3q�p��Q6���Ü�,\�^r��dn��ZI+���\��x��0�107z:`v��˼�v]�hw)e\ ����l7}�x{�������bl��º�y^Dv[���֘�0;dt�=�&�Z�j�̬Ŋ��X,V��0;dt�=�-I8��P*� ��#ت]�Z�� ���z�+�ڛC�U�;�w��tB���� k��>�^,�L��s��Z��^n�sb��B��mӡy@��1L�'6[s��#����t���,�a���;����tL�0=�:`m�_�>�&+
FV$�`��0;dt��H� 7���:�j�S����VUm�tt��H�t�q�0=S:�#��c�R�ܫ�}��. ~��xޝ��?~���w������m�,��{dLz�&�GLt����`���R�Z*� 0{���?Q�#��^�im��C���݈�Q��i�4����;k�ks�A	�`ƭ�"f�ۭ��)�$n�%�s�m�<V�m�v����٩�Z6"S��V����ҟnvtm[�I�q�n6���:���5�9�鹰�@��Z�!;�ݺ�	�l�C';XnM9�J)^\צ�㬽�j�DC�bNH��]���\5��X݋`�u��)��Fa�Nn��=�w{��>�B}���xۧsƫxX�E���;-#�vb�g�Xn�;�
�=�G��Ř���?T�쎘ގ�Ή���ٮ��$��B��8n�p�v:`:&�z�0$��J�V�%WtZX�����l���c�F���,D{d�V9]�p��o ��*�$t���������1X|��bI�7:U�:tt���� ���ڣ]�Tݖ"K$c���S�	��P����3��Mѫ�6[dyA}�8��-��%ҹ�ີ8�x���X�]�B�Y�vo������Udu�[*�'~�th�A��E�  �Q	@e���s';��RM���]I;�� ���͍����Rʸ����V����7��N ї�+�@`�&��V�ޑ�oGL��x��f��<�*�,����)�7���D���*�왙�| ��=��Ym3�qD�(�v���κ��k���$#��[/ck\�u\���m���t�:H�s�[�����e{d�V9]�p��y�f,l�f�N �� �׋:S#�i'EUtt�����|� ��,?F�E�^ڥ��g��K��HEH�-�>���C���Cj�@�b���2bP�i��1������R��̒�x|16�.�c��ܬ��É��Ʀp�`\��mӲ�{/��#*P;Пe�!��0�pg!���1�n�h7�$n�DF	#!G�:A�$�_��FIa���D���`�BbTd9,Hɐ�۹�*�$x����+�����m��&�D��LB�d��0�9M"k@+�C��aD4&ÃcPP��J�:�T�;M(�����=P�9���ѩ$�{��I9�K�*uUZ��>�wx����pu����{m���d�Q*��M�X���z:`�&��V��' �~�I<�@�9`�R��Pj�,�'K�Pۣ��gnl�J�V+��6���2	(��.�~ o���kS�|��r��~����ͷ��k����0�K%�.���t�����D�www����]��H��,ĲH��k���#P�USh���ͻ��'C���ޞ�z���F�ww~��_�v��U�RWU�6���m�������o;�fj�n��t�ݷBD��*y����S��}�j�oxp�	1�El��[m_|�o���m�<�b����m�x�6����\�m�_��b��ذ����e3��۱�j麮"���e7�u��e��s!l�2�,��m��o|�޻������oOW�ww}#C����J"
�UV�L���ͷ���pm����������_���}���o����F�R±Ka%6���_}�#7��m��~�=����{�s���}�o�pjD��Rʾ����}���߻}���m�w�6���ߗ�����x��D��T(�Uշf1�k�.�m��=���'��b����l��/}�ն��)Չ"!��,��IONO�k���A2�nrOf�CQ�;]6ݮ؞��E�Z-[�i������;�V�(���]"���/Cի��՗�����v⛝�ܥ�9�b�s�X
�i��c�1od���w:�nz&�:��sG;vٹКǷ-�pַ&K��VW4p�ʫ�p�d`i��a:y �#!�����q]]���d5�k���9�J9x#���d�RU�X�FbH�>q��Q���;vV�F��G>��9n!�J�lE���9�(�5"���ʟ�m�����6��w�/b��6��q^6��=�o�������ה��mM��%zH߻�|�����q_}#o�w���o���������'���*�+����I��)��~۾O�~�}�����$�}��Ͷ� ��������s�I���|�}��侑���z��o�d��}N6�k��y*Ԗ��\vT�����s�q���}��_�F���q��}}�����o��O;�CN��֣t�vv�#�hi���p���s�T�4�:C<���H�V�X���������{����}�e�3�U[��O�!}�L�w����fy����0�4;�v��m��w���w3�ҟ�f�n��~.�m��w��M�m�=�}��3�+k���cǍP�F�m�_yO�ܪ�y��2ff^�~\��T��we�m��o��
H⪦��v�?ߛo���8ߒ�ow�/�m��ޗ��d����?�m��"�yI]V��,�Ts�$��w�7�m���3�7�[}�������tO����s������5��Օ��v��v y�-��;[:C��T�F:�D)#�9:�r�9G̶X��ڻ������K�m�޻������x�$�>����|�����'䧫�2̎Yx�oݻ���رb�?o���~�����m����%�H�_���U�-
�p���ͷ��8m����/�q,�� �J�^AZ�)�'|^r�syέ���׭��νrF��:�-��8��%'�����m���s�m����ݷȸ�}�ɫm��rz���l�e�m�(���߾����Ԛ��߹ݛݶ�p�k��q��z�v�෎�jا)ub�]��tU����$"��R%����`�5ATH��m�����|�}����{����f$��ߣm������o��
H⪖ɜ����y��Rk�*�~P5�[�^��{��{��s�m��u�w��8�/{%�Ȥ��ڛE�Jm���|������o��,Y�I?{��|�~����m�������X�v��Ϳ%�I�z�|����k��v��{Z�V�0	�|?(|���Y�w߿�}�m������e����n��v���q�=�o�}m���ov�=ݗ��7��Ē�����1��Gl���IR4�\�m����`ۋ��sF*�t�s�˹�C�S�F�h�2Z�z�����վLc�}�{��{�c>Gxŷ�{^�{��vk=ԪK[R�,��m�������(^���I��^L�����zg�fw��L�U#{��#�Љ���YW�6������}���[���g�ֻ��՚���{�Ͼm��ӄ|`�����ߖI��߭��ϵf����wf�m�+��=��^6���?�x�#���E���m�wy�٫m����}��9m��߱�[m�{���ͷ�.H%���uvE3�l�ٺ峦�Н��#t]tGK�	-l3f���TK��㓵�N��X]lQ�m܎��2z�����qlc�����D�Wm�)B�@�����h.��e��m \��}u�Oѧ'�I󫚤r����J�fv�v�춐ǜuvZn�"�`�a���N�1��n�E�=Gi��k�Brb�\��5���tlfYrjw���w���n���ø�T�M)r�hݸ��Z6�?�~��:�J\!l�6�+�{Z_�p��I%�ڛE$��m�������ͷ�7}/Ͷ�{��~ǂY��m���g�H���ro�l�V9]�}�m�w��خ1�}�k��v��gڳV�{�;�{�H�H٩OG`*J+e�����s���m���վU�1�w�7�m���3�k}������Z-�)_�6��I$����}f�����l�ﱌK��շb ��}���Ϳ�νg�*��Ե�+5m���ov���������׭��w�q��_~o�Sr�FY"���L��W���[a�M��l�]
;qB��u�=_�w��y"l��ܥ�~��m�޷�����[��������I��/�m���#�B5����9έ�����{<ҡ��#a�#�?]T���~������j�o���f�m���u�Ÿb�mo����
8�&����7oo����߹ݛ���9;��9ն�����|�}]��E$�;jl��8��1�w�ݶ���9ն���v����N���q�߷Q�	�e��X�v��������L�ϒ�$���=;�3==�U�33������ƺ`h@b�����H���c�C�`5X��ur���g<������j��v ���[����;��.�׋�"��u�t�]DJ*�.�j˜�t$����, |����=�6��O(�dp�-�ʸ��ѩ$�;��~���68jb(A
�@A	r*����~����RN���k�96D�C�K*�yff.a��%T�u�����o(���������� <P����[��B����/�v�ŀ���*n�꺬^�<���vk�\�Om�.���'���4H�]m(��N�ȼ�,X��'-xQ�Q6w3���X�^, ׮�$�Hv����a��;�W	j�����\�U�׀sw�8�x��&M��~�e��������n����Uw�ذ>�,W�HҧSt�ʱ]��OogL��b���`[�	JԒ0��+	Q"��`�U0�D�}}���I9{:c�!B����&��pm��<�>\>�� ?{׀o�� ��7Tj��n�2:_kɯ7V��ĺ�]h�礲<�`��������wNx��T���]��=�� ;�v���[��;�� �|�zȣ#hw)uk 7��:&N޾��7�b���g&��O�W��q�x�����׋%򊮧ذ���?}MS���RR�jfB��p:�Ew��,Ͻ� 7��СDG�y���pʞ�UW4���\�wk kŀyz�~�����8���5$��	������q�1"A%Q�`E�0*A�"7I�_)�-E�$K�6�^f-���fGi��5�\4��!2j:`�H��Z	!q�f�6ɜ?���&2�w&2�4�|F5��.&�ʝ�	�RRRVVc3�ńM��BdB1"FH�0a H��1�1���
2�ŤR).��8��"QO�ᵤ�
sk�F�$VBHE	,BH3稑��aLce�#$IB:f�,B2dXA�Gp]�!B	`�F#I	��FF��-K	[B��!YHAaM
D���	�a, B���'��i�XR�,�������ң�X�bK���';j�>s�����5�{mQyf�W)R�9y�9t�{a�s�v��q4��r�Y��)e����a�3��K�Nf�up,����V$�Snc�%^U����
W�U�+nN����v�bi�vzS���t((���%���M:���be� L̴��.0�V��q�3R�v;rlֱ�y9ǴnZ����	3�ngv~CsY��mjWfԅ[�����ҫU��0Jhm�4����++�/lB�5뎶�#T[���;ikҐZ�;\�r��R�םƃ"oWt
�8裓�i���Pxwa�Ԏ[�1b�t�<�â�f�+�.˒ưΕVPU#����|j��%h��ʴ�7����M��I��mvTn��x���Q'��Tk�u�[�ݠ�l���J�@�:nwLJv�n� %)En���/i墫]�CZ��d"P�	T	�g��b��� P��nB� �zU'5R���Z�P
���v���uΠ6�ӻJ��#=��+�)Y�;p�0g��m�v��iI�����+�"=�E<��5t�u�8wW.QuF��ℊ6���Q�'�|���r�m�F�7T��CM���S��b�0��&�:1��֝�1�YY�հy�yӍ�r,��dq�Q�(b<�z>z~��}7Ź���v����	�t�Қ��B9�+�qR��Q���
p"헞Z#G4�nLTOT��"g��0��]e;F/ClY���m�⒞m��HP	u�K���t��E��HL3Ĳ�+7�Fv���9���b��y�\�$GWN�r[�m��$����T�J��/\�TP�Sۓ68ƛ�������E�K4�1�Zy@��I�n�J�69�u�v��]��k	�[��[��� �j5�Qu�p�D�Cm:6af���ˌ�F6�*L��nUHW�m���F�kDj��v��Kl�Y;�kN�5n;@���=�U\ql��/ 5@U��V웱�kcv���A�Q�,,�%�ŋR·�|�W� �p8�|�PS �G�? g�??
� &�@���fb��L�r�j�n��:q�ciGr�A���@\l\�Dk��}S�^5�qFG���u���tj�r�ˆA�b-�f�s�sq-؞4v?{���]
���@��t����K]u��ϒׁvF�W\p5�sSd�{�z3��-��	<��gz�'	8l��A=+���<�GRL�$s��M�x��N�h���$�f���\!Z�=�ǻ�����z��_��4�n6R��6.�.u4�76.3���Z���-�:wܽ����"|��B�Z��ڼ����mٜ�׋�~��}� kh�����Ad��[�7��o��bRC���\߷�\ �{��ɰ޿)�cD�
[�Z� ��v,����zQ�޼��� [�=���8\��e\f,~�����^ �v�p9DD��ߖ��sS]uJ��(��.�`��9(P�
.u���~����7�w��}�t�kR�F�ջt��sƛ�y�jlk�$���F��S �Ϋ����b�bH��׃��U;o�{��o�~m����z�%��9�׀k+��Ǒ�*�a-o�~��X�I!"0H����B�{���I'9�g�o��?��1H{�?���WU���n�`}�X�7xr�qU��p�ظ��v{
Yj�r�j�{17������8ͼX���+Ͻ��9u�JGb
J*�m���������L��`l!qդZV����S<g�9�w;UW]�=%�u�jb6p�A{F�{e�|O�Ɖh������8�^, ��~���!B��]�g ����	%dp�-��p����fb�����;z�g ��ٜ�!(Jd�鹩�YR&�r�U������[���D���@P�y�gsRO��hԓw#.jQ1s�M]]�z��%��ޙ�7�~0��X�(�J��U��޲x�#�"�������73���|�?&إ� �ٙ��B�!b�=c`�T���݇��NE��,c[u�0�2#k�-'}����#�I]V*�q�O��w�\ ׮��3�G����7��@��K-U�W-\ �wo=�6{}㋀w޾8����5v�S�؁Y�Kp}}3�|ݳܢ��� 7�x��R�E]�e�MYs��P�z)�߼`�{ n�xG��B !��Q�!)�������N q�S�*�S%�]��ـ?�ŀyz+�޿��W�N��Ӏ�荶H�dd��8����[̎{uY��6q�7o>g:��巛;W~��U~�(�M����x�wS���O/������?vyx�<W��r�x�֧=䪇���� 7��9$�:��?�y$U�ʟ ����w���l��׀{f�>��T�7\V*�q�N�I���ˀ�z������}��� ﵖ=
Ij�r�j��]�Q	��J=���~}�� w�5$M,� ����Ɇ���`5�eˁ���R0�IZK�,NENi��v�o)n2I<m�����6�y!�{]��»uִμi��ݗ�^��J�����gnn6��:�RR��3�����BWv��t��C��K+��/h�8-�q山nU�ι�D�en�s����)�[�t�����vkl�n��j�K��y��yxwG9�XD�M������MпZ/nQ,X^���E�v���>9���SvF�.؝����؋?�b�
�Jr;'kU�z�Ox���f �v���">�9�� �G��E]�e�Mݓ�~{l�D���� =��6NyB��_wL�VtwWwf��� o���BqU�W�����6���"��C��S��I%2���u�N��fB��{{8��<�<�
�[�7�t|�D(�%
��x�?_� ��x���S��p۱u����Obwd�uA�x`��[���ˎ��<�r�?}��{����O'�늙.��}�|`�l���JK�z{��������v�*�$r���*�1P�J<�Jh;���u?)�>nٞJ"=���I�Q�,��W$��U���^ ���âL�u�{��8�R����m�%����{����	D�}׀>G�D�
[�ʟ ��t�%��8��������\��q85k.�v���:���N��]N5l�]�1-�s���*��!�Ð����-R�O��}|`�w�=����;� ���EC�'#:��8�۷�Y�=������,���>޳��A1u�5ww�s��p��0�"�A	(K�%�B�qY^�, ��� ���67�d�P�-��{3}��� �}�. w{��噏�}��o�~��]���R�i�7�� �I=����{����8�X�}��!#�UP�t�;P^�q�9:$ݮ�$�-���-�j�{r��GZ�V��V9\�|��^����7l�~���ŀ=
�䫪n�)��wWx�֧9TUw_}݋ 7u�z!G����yP�v�q7vN���`M�� �0'd��
��L2�)�.*�U�ف����`o� {M����	(؏$������A5�5VZ�ZT�;�L��Y`l�避�x���I��7ǫr[K��෎�(N�y")5��%�=�B^��=g����K�p�'��@q�����>�{�\n�{Ϙ�z���I�I�EB��8�^,�Jd��ŀ_^ ������Ĥ?�����7]��:�쫀y�ذ��:!(S<븜���z�JGj�r�j�_f$���}p��S�~�x��x�Щ��:��
n�U�� ��' ��}�~�� ~�� ��*㧦�]�V+�E�C�+��X����tJ��
�Ɲ;�A�����\qx�1�~�wG�WS��Rf㕂|��^���[Kmk �MŎö�Om֓�I�x���C��.�[�Ɲ]ni"�W�8]׷v��]��.�{IMa��pZl�n�px({���f�{q���<�cD2 qZ�vډ[y��e��F�u�bG2�e͸N�F�n��qqrK���LSʤ
e��:4bkj�]�nIk�j5Z=g9�n����}�26�)n;h���o� �ۼ\ ���ٟ0��x|�{�e�t�R�.n� �oZ��u�����׋��6{�z�=br0C�Gj���� {M���ηذ��X�;sJbbU��%U�(�v�N��,��,%�QU�޼���ULUX��XQ%թ�>z�`
#���� �����>���*�U���e��إ�7PF��!��g�������t�-�f�7g=����v"�J��Suk�;��X�7x�֧�,K�����{V��H�U�Z�$���ΰ	�}S"aj$L:��¦�oA� F�"�"H�o `��-��VF�
H�!����*�"��0# �p	G� *���_��|�� ;fr��%26/�OGbe��������p�X�B�D$�Uy��`?z��ZT�b@!/�b�au{:z�b� �0�Ř��n�> t���n�KT�v��`�DD���s��p��. /���6��f���v$E,��r;u��Ґm��X��J!Eڼ����wz�f�~�*h�MœV~ {�x�֧ ���س�﯎�����x���=�jp��X��0~n�Д(^�����<���P�,�����w��F��O�`�$H#�KoA`#0@�ƀ�h���H1�j�,emH�&�!�%�jH>qfE \p��h(Y� �0\b:H��Cz*�PȒ2	C8��4�6�v�z9���\����������҈}P>B�c��o0�T�� � p�v��]��uN���:�8�� �hl4�iQ\��8eSb mW�t����ݞ�|v�6�[*q7*���X���~X ���kZ�����7�ґګ�Z��۷�ts���� �v�e|9qD�W�d�/3K�y�F�IƳ�r�f;fu8u���I��(��7R���
�+e������X��<�ף���x����ax�%���`l��6(0�ݼ{;��͝k��XK�*��sv���X�7xyB��WyN ������C�"l��ܣ�p=��}��9��8�^,�DZT��0Ϸb�<
��-���O�~�� ;f o���IBM��wb�L�����k���s�\�;�5a�˵nҀ;��+"��U��IJZ�Q�T������?7l����H7O����k���iQ�w�����P`�&vtO�~��<��ۡb	�R�Uq�\� =�v��â)Uo>ŀ~�0Щ���&���WUw��	%�J���' �w�`�l������0����*�໵8�^,���/?~��>��kZ�Зh��%�UZ"毱�.ԧf��y� ��]iV̕��i�L혘�˷/l��rOj��}�Gn]mq�y<>�*���Ǉ{\�V���n �8�)�r��{etY�n�Ϛ�:k'[�ڸ�٥h8w��W��JnэN���O^�5�͞��4�� ՚�vcl�mF=�X��b��IKpt�r{7)	u����6�n�Ę"��-�vy���������v7��.�K�Kc�m��(A���ց����y�b�ɒ�m�����8�7J��Wj�?{��8��۷�ogu>�{�\u�sdNFv,����w�	&�Q�]�p�ذ����,ě;龊��x*��s��p��X
"=^~�, ��_ ��m5ǒZժ��YS������������IBS��)�;]��Yn�69T-��o��.��Ic����=�|� ���.�~��p��N�z�G��͜^��t�����nu�qbsasn���c�!�X�Z+KUq�;W��z���8�^/$�$�Hv�b�
��ab
J+-�{;���b�wG��	 P�A�@�"~���b�>�{ o�� -�-+�5v\�v� ��ŀ?�Ň$�)��u�پO�~kwJ�`�Z�v��bQ�Y��X�׀}?j�
'���`�&��H���Qʸ�۷�ogv�����ؠ�ݮ.�)%B�+dUx��c����jm$���m�䙮�:ܠ8�{Wº�x*
��-�۾W�|��������u��}uS8�����.�R`l��6(0� ��U�(�C����+��6ܪ��X}�� o��/B"*"T�B�BK����x����.����WTM+�� 7�� 7u��>��X�w�\��%�RQYm�{�W�tB�����݋ >�]����U7}ڮ��;g�Nr���&��[mS�uě]@�\p�'ۆ=-^�6��ܽq$��>�~?&�`�x��ߢ�/(���+�:����\r��K-��}��\�ca��׀��x�ۼ\w��sdM�Ц�ɫX��� =l�:"gw����w{v*���*����M�w���ذ�`l��P!%�$Uk���V�<�J�j7�^�{�\�}	q����׀u����E߬�%��-��m�fΞ�5��7d^K�utz7N�4f�F�q~��}+��J��K��ذ~n��~Q�Cy�,}�ٞ�#�Y�����y��@�w����X��Y�<��;��|��(��L����gGLH��;�v�ou=J��*��^K�En�|�޾0(��(��w������XK0n�,R�W ��t����� s|� ��ŀ~U�(5J��!�Y�Y��es �
�R���4&S��;v�I��t���&�x�Mֆ�
6Ͳ��<��j�=K���*�np ���n��������}o��kjU��K3�����0J�T�j�E�ۖ0n��Wkg���c�4:{Ͳ���y���gk+���Z�rv#^d�	
��4������v�b���u��s��9����8��$��: �6dT��)����^�_���Lbm�!n\�1��l��s'3d�N��n�����u�a� �����wf�P�"��!;�v��7�޼ ��R`l��6(07b�J��/�R��j� �W��ɼ���� o��w�=��f�R�ʯ ��\lP`�&;�&�,̈W�j�L��h����)�����u��������E?w�X���=E7jn��R����#�� �����6������'>C�Bax4�
�A{.یc�ώcS6�fv�� 7Tqcwg�,�
�K� Wv��� 7�^��l�?7l�Iy$�_Pk�zp{���d��¦˂j��>�m�I(K�J!�_�K0�v�{7_ �wx�y,ě:����n��T�TUY�v��~���<�B�3������7Bul�q�N���3���po�0�m����{8��櫏���!-|{��p�wy��=�{��}�w_ ޮ�[f6�:���\����
z�Z��Lh혙x1t�_�>s�N�R�H0����� ݑ�۝-�;��Y��1b�˴�I$0&���Ζ��у��N oz�3U�;Uj8��p�N��'9��MO��$Ȃ���I)���~�ذ�T��wE�����;z0`{yA���������|� �����GUM��%���0?�����od�loF	}Wu�� ��M�{4n�:]gTt�S�aX⮑��n�TmcIE[��+W�8Z���j��K$G�ޟ�0=���ތ�P`H��dC��u&�\�Ӻ��?w}�`oE�`{z:`wE.���_� �Ew8�1`��f��B��}�X��� ���7$Wh�@�-`rQ���}� ��78��	GГJ��YǷ�ˀ}�l�k�K*��J��`�׋ �BIz!%�=��~� ���N ~�׹-���2DJ���q��g��r=b��ؤ���@-�f�<;�����'�[0J��Y���0=�%�=����噋�������?%�K+j����6b�J"d�w���ŀ~����$�l;��(ԕT�.p�o���x��DL���8��b�������V%X���C���ے[� ��������I��:�v���-��t������_}�ÈC��$0�ZD�a�@��hD�ZR1���AK@\�/�8L3�� 6@"������5�Aȹ1�f�G ȩM���(d2&L�Aɒ.��@�X��^w�����X��Sd�
q}���єH�H.���~L���,�/ˏ�h����m�4�e��z;4�(�����Æ�^�{�� ^�2��5�%����(�]��M#1�C��##�CT#����Q+���B�l`���)�i�Tsd%���l"*Z��sn͵qn�7�vt9�d�&ۓshTlE�����j��3��j�vB��l� ]�C]Mv�����uF!�A��[�s�7!���G	Ym�fѭF���JK�f9.	,�%64f���H	Q��३u۬��@�����pk��>��=�m&���.г[�>�ݹ��N�;4=	� i�PAj\�i��i�KL��B�Qtl�` ��� !D��W+���F�N�����c�nJ��{r��8{=t�˺2�-mv*�T�s�/[�Ǡ8��؇��+61�QڷA֟Gl�wf�{�Q��s���y�c(h�d��+Z�Jذ���X�AM&���jM��e{[fvڏ*�q�d҅��VV���\2
�b4�(�X�N�-�2M�����l�pl�5���j�@��9��4�vܘn�n��8�x|�OnP�d�v{N-w6�m�v���p9u3Y�s�.4�e�j�HđmҩFݑx89K�u���{Dc�5p��2-�����P�e.���r�����������<Ҳv^��]	Th�rj�ن�$��v^xZE����u��s�K������K�V�3���\p�-�XZ��ʐ+�h�Ț�b^�q]�f՝�OfvmU�Y�@�1���a;t�]]�Y�'S�b���Z�U�l�Ӂ%X�fv��wXXz��W��x����4��������vB`*�p�*f�����X��'��c��m��f9�f{[ڌs��&皔��դ�<���4q����5��&2���eME˒̓�V�ԛ(ʺx�\��f9`����U��%��ٟ0F=0PnJ��۳�0��9�c�ci��9,p��Uiճ��J�˛iz�+d��B5���ZNݤ��˜f�xR�DO��&Q�T��4�Gj��E^���:���X)�«�p��T�E�N��3���d�a���s�b�]ٸsl�H�E�kB.lUv�%��.۪�
�tN��ԻR�N ���pb�i��;2�y�s�m�w���8�u���Yx̖�:$܍�����:��g
q���}����8�ٺ���w8���r:j)+$뙹����%�yt�g%ZQ$�q�N�\��+����$� ��e�qn٢���R��N�|�2��Ԛ�x�\�ێ��`�&`Bv��V�tVz�%n�Y��jố�/s���r����*�I_@�� �������yB�	{�u�N��M7$�Ta`,07yA������-���Ӌ��,���X�v�#v�[h�������-��t���5BB�Z��Z���x���\���8O�w�.�l��ij+E�e��A���ގ��%�����������B��3Q,cr�:K��6�e���M�D�1���~����q�;�K�3e�4Z��_���>���D$�%����. wZ������j��ԓs�5� G�@6� F��DYCuߧ �	����_�RB���{8��Kı=���g��,.B���n%�bX��}��Kı>�6i7�@�,N{>��n%�bX�s�٤�Kı>������3!��3t��bX�'=�]�Mı,K�Ͻt��bX�'���i7ıDlNw>��n%�bX�w޸����&rLK3.1�I��%�bs����q,K�T����&�X�%���޺Mı,K�ﱳI��%�b{�&�\�9�9z=�e��[�.U4nN��$�8gS<��͔�]�;�1�ڠR�P�r������X�'���i7ı,Nw���n%�bX��}��� �b%�bw�����&bf&b�y3�?�$-U��%����%�bs�צ�p��1��~�4��bX�'}�߮�q,K�����&���bX�9�g�L�g$�&33���&�X�%��{�f�q,K��s�]&�X�`oM�z�@ٸ�D�}��Mı,K��4��bX�'=���S&Ks2ˉ�I��%�';�z�7ı,O��l�n%�bX����K����Nw����Jbf&b{�����u�-RK_1|b�,K�w�4��bX� s����q,K���=�I��%�bs����f&bf&bk�ݍy��B�D�%No/D� ��ٍu�)E�����L�j�=/k�n��p��I�W1|bf&bf.�㉸�%�b}�٤�Kı9���@��bX�'9�l�n%�bX�{���VV�̘��n�q,K����٤�A�,K�Ͻt��bX�'��i7ı,Nw>��n%�bX�{ǜ>e�%�c®b���L��]���I��%�b}��f�q, ,K�Ͻt��bX�'����&�X�%��V�z�%��v�I_1|bf&f(����Ɠq,K������n%�bX�{��4��bXp�P>�g��3�(�L"�:�O�kܺMı,K��!u���L��.ri7ı,N�>��n%�bX�{��4��bX�'=�z�7ı,O���s�&bf&b�Z�y��n+cd�Rط2tZ���j��.+�K�Z��V��P}�$)��p���R�k�/�L��,O���Mı,K�Ͻt��bX�'9�l�n%�bX��}��Kı9�/��2d�3-�4��bX�';�z�7Bı,Ns�٤�Kı9���I��%�b}��l�n%131>��yK�:ꖩ%���1X�%��w�4��bX�';�z�7�lK�v{f�q,K��s�]&�X�%��ٞ-�q�q%̥�nri7ı,Nw>��n%�bX�{��4��bX�';�z�7ıQF��;�Mı,K��^��ea�3	q�g:Mı,K�w�f�q,K��s�]&�X�%��;�Mı,K��t��bX�$ǐ�����=�sܘ7'p�a$��"ǷfMY���u2�n��T�]�����xɶ��ìYigmsN���8��Nn]�d�g�۶��C�{Mƛa�jr�ԪY�d��ʍur8_v ���j7��p��6n3�Lv�v�5թ�n�-�0�\���S�	q�i
�W+�l�9���(�;:	�Aj�P���e�h���tl0�93����������>���D��[���p���u��3�t��A�*�j �p���GF����[3qri9ı,N�����Kı>�}�I��%�b^w�΃��&"X�'?{�٤�Kı;��	�	-���Go1|bf&bf/��l�n%�bX������Kı>�}vi7ı,Nw�ޓq?q,N��u��qq���1f1���n%�bX����:Mı,K�w�f�q,h�lNw��j	"s�ѥ$D������	�Lc�SPI OD�ݞ٤�Kı9�{zMı,K��i7ı,K����n%�bX��gLx1Lc&Ks2ۋ�I��%�bs�����bX�"}��f�q,KĽ｝&�X�%���=�I��%�bt䙗��ۢf�R:[�ʗ��������5<�t^�F�k���L�v9�����5�7����,K���i7ı,N����n%�bX����iı,K�����Jbf&b��<�Kh�:4�U�_�K��}�M&���@HR3��� 0���eD �bb%����f�q,K��s�]&�X�%��{�M���1�LD�9���q��ᕎs	1q���Kı9���I��%�bs����q,K�����&�X�%���^�Mı,K�{؛�8�,�I&%��ɤ�K��1D��~�t��bX�'=��4��bX�'{�zi7ı,O��]�Mı,K����c��S�v�I_1|bf&bf/��|���X�%���^�Mı,K�w�f�q,K���]&�X�%��{��;�Jf�,�n��],�:���y��過��	�a-ܸ���c���Z���Ѵ�%�bX���~�Mı,K�w�f�q,K���]�X�%��;�1|bf&bf.�ў�XX��uK%�Mı,K�w�f�p�c���bw�~�Mı,K���Mı,K���4���!���b_޾1�1Lc9��̶���n%�bX���߮�q,K�����&�X�~Q$>(��V���Z���Q(]��ȟ�s\�Mı,K�~��\�񉘙���u�򶱂��mRc9�Mı,B�����&�X�%���^�Mı,K�w�f�q,K�0B~�zr����$//Y�}WVM�u!rۜ�Mı,K���4��bX����I��%�bs����q,K��;�Mı,K��[g�bg9��;j��y�v�7sgzh�1���m�$�vn�ط��.�#3�{z��}��oq���X��}vi7ı,Nw>��n%�bX�{�١�Kı9�k�I��%�bw��&��#��K.n.M&�X�%���޺Mı,K�w�4��bX�'{�zi7ı,N���4��X���][�=#��Qv�I_1|bf'�����&�X�%���^�Mı,K���&�X�%��g޺Mı����b��2Z�Q��W1|bf+ �;�k�I��%�bw��٤�Kı9���I��%�@`R�@�$E ��K���I����L���3��Z��d�1|bbX�'}�]�Mı,KȌ^����I�Kı9�߶i7ı,N����/�L��Lź�/�%���dl�27[���t��9��ܻk͝�vO��m.�Z*�#dv�t��us�&bf&bﯽt��bX�'��i7ı,N����n%�bX�wޛ4��bX�%��ޥ�`�u[T���_��������4��bX�'{�zi7ı,N�ޛ4��bX�'=�z�7�b�"Y��_1�[)u�:�%\�񉘙����k��n%�bX��6i7ı,N{>��n%�bX��}�I��%��_��=,�`��@Q�s�&bf&'��M�Mı,K�Ͻt��bX�'��l�n%�`~f"{߷�i7ı,O߽�8�nrI,�8�4��bX�'=�z�7ı,?<����O�X�%��~���Kı=����n%�bX����dA���1��ɗ96�鎫9���!HP�F�yu\�1�Ū��=��:�Ξ5]icK������7�c84�cn�L%��"�r��l��jFQQ^K�쵻�rI5�^��ic�D���ux7kmͬsȎtc�R�0v��&�-a�Dv
2������4Ʀ�e�n�=��֋���6��݁�q֭�T�l��Z��QZ
'j�~��LLc8�Ĺ����j �)�
��{"��:vnۮ���F��i�%ŠJE���+�w�{��7���s߶i7ı,N����n%�bX��}viwı,N{>��n%�bX��X�3̄���e���_�����{�zi7�D�K��~�4��bX�'g���Kı=��f�qlK����<��8&i��9�34��bX�'��]�Mı,K�Ͻt��bX�'��l�n%�bX����Kı;���q..L��e�&�q,K���]&�X�%��w�4��bX�'}�z�7İlO{��4��bY����ǩ,+[�����b���N%��w�4��bX�'}�z�7ı,O{��4��bX�'}�z�7�f&b~�4G�Q0x�VJ�;i�d���'VH����q��Vإň#�ڻ�n-p�4ɋ�arfc4��bX�'}�z�7ı,O{��4��bX�'}�z�7ı,Os�٤�Kı>�=��f���d����n%�bX��}vi7 &���Ȣ�""� $x ��q0T>���'��n�7ı,O��l�n%�bX��}��Oة��'�޿�ۜF79ae��ɤ�Kı=�?�]&�X�%��w�4��`*h�"b'}�z�7ı,Os��\�񉘙���n��V9,�@��In�q,K��;�Mı,K�Ͻt��bX�'��]�Mı,�D��{��n%�bX������b�&i0g9�M&�X�%��g��Mı,K¬~����%�bX���~�Mı,K��i7ı,O�=�}��m�:�7iNH'�1�iώcU46(�mv]�)"b�E�%�2.*��;b+A(�.st�D�,K��~�4��bX�'}�z�7ı,Os�٠�(O�b%�b{�~�Mı,K؝��~q..rK32ۋ�I��%�bw����pVı,Os�٤�Kı;���I��%�b{��٤�Lb�"X��}=ssf	3�rf��1��&�X�%��w�4��bX�'}���7ƋkK'D�(�P4AT�Ċ���Sg<l�E&�ϝ��B�c0�f&	 L�Dp�!2a	Z��h�lO�!\��ĉ2#��0CI��m2�\l
�D�¬P�8@\d�`0cA�%�V\ �M
�LPO�����	��}O���?T�:@�q:��L_�2�ѫ����L�� �{4+l��گ1��Q±�*��3"�P���|
�ϓ)�އf�D= �; �AH� �D�N{f�q,K��s�]&�X�bf/-�c���G[��U�_��~B!������Mı,K��߶i7ı,N{>��n%�bX��}�I��%�bs���.q���&Hf�3I��%�b{�}�I��%�`�}��Kı=��f�q,K�ｯM+�131{���/W�4�U�j�N��K���k�̵���b*S�.�O$�ۜF79ae�q�I��%�bw����q,K����Mı,K���4��bX�'�w�4��bX�';٩�c�[*�-$��b���L��^��f�p�,q,O~���I��%�b~�{��&�X�%��g޺Mı,K1~���P�q�j�Gm�s�&bf&'}�zi7ı,Ox�i7ı,N�>��n%�bX��}�I��%�L_�U��mE�1��j�/�L��V'�w�4��bX�'}�z�7ı,O{�٤�K��E#"�F��!��x-T�'�g��&�X�%��$�L~s..rK32��&�q,K���]&�X�%��w�4��bX�'}�l�n%�bX���l�n%�bX��g����3%�!���.��vz��z�J�v{R��]%fv�̀5�v�==a#Vϵ%<�~=ߝ�7�ı?~��Mı,K���i7ı,Ox�i7ı,N{>��n%�f&b��d���%lN�IW1|bbX�'{�zi7ı,Ox�i7ı,N{>��n%�bX��}�I����L���GaD<2��\�1|bbX�'�w�4��bX�'=�z�7ı,O{�٤�Kı;�k�I��%�b{ݾ7nq�兗%�M&�X�%��g޺Mı,K��i7ı,N����n%�`~O\���߾\�񉘙����\���$�UZI.n�q,K����Mı,K���4��bX�'�w�4��bX�'=�z�7ı,N^�ҧ2D�,�U\� �R%� C���PŘn$�b�2ZzQ4��,=jQe�ا$��X�9����y���+���un4vX�\D˪����Sv)lH5�d����x�6�A��1�m���!LQ1[7m���,f��ۈ�R�p��M�K�֮�4g���n��X(�q�p�����b����:v�I��j<����V��3Sfݭp[/Brq<�㫗e��,E��׽޽㻯��v��Qr�]9�օ��g���%�mc��"�m-�e���ܗg�nu�8�U����131{����bX���l�n%�bX��}��Kı=��f�q,K���|zc9�3���q��&�X�%����&�X�%��g��Mı,K��i7ı,N����n%�bX�Ĝ��e��d�0�ɤ�Kı9���I��%�b{���&�X�D�"b'��_��q,K�����Mı,K���2И[������&bf��{��&�X�%��{^�Mı,K�;�Mı,K�Ͻt��bX����~�+),buRJ���13���^�Mı,K�;�Mı,K�Ͻt��bX�'��l�n%�b����~���b*N�[�e���Z[�ջQ�]��0�u�Q��3���$�'[�������n%�bX���l�n%�bX��}��Kı=��f��>���%��~���Kı?~��n��0�9a�r\d�n%�bX��}��/�h���qj%���;Tx󘘉b}�}�I��%�bs�צ�q,K����f�q,K��;�<�jIl�����_�������l�n%�bX����Kı=�٤�Kı9���I��%�b}��'v��v�W1|bf&$��O{��M&�X�%���~�Mı,K��}t��bX�'��l�n%�b������ ��)�_���b{�{��Kİ��G����I�Kı?w߶i7ı,N����nbf&bf'���B�㈶�9��^�q���h��BݮvM��z�Ƃ��B��v�j�-*��b���L��]��>&�X�%��w�4��bX�'y�zi7ı,Op�}t��bX�'1��B��[������&bf&b�o�ZMı,K���4��bX�'|g��Mı,K�Ͻt��bX�'���rz+T��uY-9��131n���Mı,K�3�]&�X�Cq`�:��Q5�Ϸt��bX�';�zs�&bf&b����]x<*`W)��Kı=�=��n%�bX��{��Kı=���I��%���������Kı?w߱7nq�兗&q���Kı9���I��%�a���|i>�bX�'��_��q,K�{��1|bf&bf/����RB���ɏT]p�4d7�:ݮ�?��}�Ik��n	�H�ٹ�V���������q���X����4��bX�'{�zi7ı,Op�}t����%��g޺Mı)����{�$��(�v�b���LK���4��bX�'�g��Mı,K�Ͻt��bX�'��l�n'𘸡����������+c����ı,O�3��I��%�bs�ﮓq,��;�Mı,K���4��bX�'�''��0��Hfaɜf�7ı,N{=��n%�bX��}�I��%�bw���&�X�'��F �#+ ��b�a �� �+���(gE0L�(<& � }Șɝ��Mı,K����`L��UqI%|�񉘙�����zMı,K��٤�Kı=�=��n%�bX��}��Kĳ�Ė%��'�S���b�WI$�b�jO[���"͋9I�At��KИ���9)rg�v�D�,K����I��%�b{�{��Kı9���@��X�%��w��n%�bX��|_ff���̈́����n%�bX����7ı,N{>��n%�bX�s�ޓq,K��}�M&�A#QI����*�M)����
�w� P�����j	"~��{^�Mı,K�W|���131ow��JՒ�T	U�1���Kı>罽&�X�%��{^�Mı,K�3�]&�X�����k��Mı,K��̞n�3�3���:Mı,K���4��bX�'8g��Mı,K��}t��bX�'�����Kı7��X��P�"D��nw�l���3�u�� ��Z�Rm�Ҽ�h�u��ҍ��s��J���6�ͫ�3zy��u.�A�x,a�;\v�ݱ9������\]�;��c<M)����l0�s�f��֑�t�х��;	lkn��&Gi��kH��K�������!�M��yBkr��n;L�)=�OFMp-n�u�!�GX-����r�ÎҷR�D�FN9t_$���+��8�����c��۲�Ê��Ojx�� -����uer��9z�6:�?=���I3�X�ԭ�JsLL��LŽY���q,K���]&�X�%��=�Mı,K���4��bX�'�Z֣�Y,B�L�����131w�ﮓq,K�����&�X�%��{^�Mı,K�3�]&�~H������i�����eU�$���&bbX����4��bX�'y�zi7ı,Np�}t��bX�'���4��bS1ym����T�N�쫘�13��X&"w����Kı;�>�t��bX�'���4��bX�'���i_������n�ԯ��b
�9�q,K����I��%�bs�צ�q,K�����&�X�%��{^�W�&bf&b���?"���Gcp'��̏U�ۭy�&�t�,�W�xtF{et;2Z�c�����131w��Mı,K�{�4��bX�'y�zi7ı,Np�}t��bX�'y�b�JՒ�T	S�S��1313����M���؆v:��K��^�Mı,K�3�]&�X�%��w^�Mı,K���O7x�ř��fq���Kı;�{f�q,K����I��?�b&"w���i7ı,Nw���1|bf&bf.�/��=%���ly�M&�X�%��ﮓq,K�绯M&�X�%��=�M&�X�%��{�4��bX�'�;N���c8!��̙�n�q,K�绯M&�X�%��=�M&�X�%��{^�Mı,K�3�]&�X�%��W�����̘��3�TƂ狝����Y��`�g��b�]�E��laH�Ϡ���~=ߝ�ı,Nw��M&�X�%��{^�Mı,K�3�]&�X�%��w^�M�L��L���~�Q��u7m9��%�bw�צ�q,K����I��%�bs�צ�q,K���צ�q,K�������ea��	�q���Kı9�=��n%�bX��u��K����`���\\@�?
FQ��5���Mı,K�~���Kı9�Y�q���$,�3��&�X�~"w����Kı9�߶i7ı,O��zi7ı,Np�}t��bX�'��I�kU�ژJ�r��񉘙���w�٤�Kı~���Kı9�=��n%�bX��u��Kı>ǽ$��
1�)d��*�I:�$4v���WR���,8�A
kb��9-Y�&s�I��%�b}�k�I��%�bs�{��Kı9���C��%�b~���/�L��L�ޗ�g��V�+�8��n%�bX����7�!��&bX����i7ı,N���i7ı,O��zi7𸩈�'1�}$�)%����[_1|bf&bf-���s�,K�����&�X�%��}�M&�X�%��ﮓq,K��s����EFYUqIm9��131~����bX�'���4��bX�'8g��Mı,��B2�J~ �A a�B~��߿o����L��]_�X߬�Q���nʹ��X�%��}�M&�X�%��ﮓq,K��{�M&�X�%��=��񉘙���n�8/HݴuJ���,I����U9�gmi#;h��g���m�;;O��ex<+W)�_������W|���bX�'=�zi7ı,O��l�n%�bX����Kı9�Y��a�� �겾b���L��]��Ɠq,K�����&�X�%��{^�Mı,K�3�]&�X�%���jyX�p��%N�Nb���L��_��l�n%�bX�w���n%��Hb&"w�}��7ı,N���4��bX����cA��$�����b���L�IP�������Mı,K�3��I��%�bs�צ�q,K��D�~�Ҿ1313��$��,U�
�e9��X�%��ﮓq,K��{�M&�X�%��=�Mı,K��^�Mı,K$����r�{ބ�!1��	&�U!$�*���p`���!	Hđ��$ D~g%!H���"1��21� ����ɩ�RL��I]�t������1��9��H�"�1�@&p��I�	�z]�$&�$�H�B!��9�Ҳ .�Y	`�6����a�Bl � �`0	!@�?UZ�BH��	5�m�؀B*HF(F(Ȱ�I&���l �5
��s-6��KS�#$R1HH@� HŌH�X�1`D� ����N�ˋ'�1��=�${��MrC	!$
T>��:t: u��uц�0��~�w"#دM�# ��`�#�Z"�j�d��r;tg\�����0��{^w��c�xrKȷ6�%��&=�P�`�Xİ�ɱ� ���Ҫŭ
��5@W�v��4�r�]tںkK^��xtD�6P۠�[j�*kd
��)5l�s�L�dL�V��.��5%�����b���L�� �VV��A
Sj��r�l������˄�\�J�rW��.�e��JgbI�vW+� �m�����J�U"����Z���ڇ8Pڪ��5�v�a��v��gG�x�%�e-[��5�@����ۅ�A���6{!%Hc���"&�lc�v�r�]���ݵ��v[�`�+� ͖��f��)����:m�$h���vStRoi�y�v�&W�[.�"s��B��t�t�[![
n�v�(�^�ڷkv^jδ�6��Ɛ��]A�6��۷a�,��)��A�Ӊ�룘�O]d�Ҍ�m��W�[Q�+NR���h������j�o]�&�$ �2,����۞'�5D�ٳf���$��yy',��n��M�K蝦��]c:Sz�J]z��,.�z�pX����;��b�e�f�v�(�D���U۵��9��9�^�e�
�x1y� 6Z���q�qZD@�zڶw�ã��PMO
�`6�z���Q��۰6˵Et��p#!�����k	9�ag����$a��Ѱ++R�5�w&�<Z6	v�\m���d��=��e.y��s��;Nq�^8L�7lֲ�]�W<��ZII�m��)�������U�a�3u��lX�g$��\��.��u���3��P�J�) ��4Z�S�;ZweHx6���g<u�C�)�i�lA�ϲh�dò��co=�t�OWP�]�+�l�F`���Bk��*3�r*�U(T�v�1�$�[v '/[���M�(.�+�KP��V.�tʖ�gٞ�����-���+[dٹ-��Kq6�>�S�N�U�ZB�vZ�cB��� �g�ݢ6�[���jK�$���s�i2 n|+σf��ȺD�OP�;�ڀ!���Ŧ�	L �x
PE�(&��'���u�Y�ی�	��S��T�58-�Z�@�]�&"\��]�'N��b�2�s�l�imI�U���ؔ���ݗR{;[������JEkJ�:�^%]�]@�s;1�[�Z��s��t�d��Y6q��*Ll���&�ktt�rlb`�Z�����']�F{[<��f@XLpuH�z×�ObfMu���g3�m�%� ���p�\]I��3sq1��/#�uÌ��okf�5�t�ngk\=��q>�C�e�:�Kjy*��b�13���4��bX�'���i7ı,O��zh?��&"X�'zg߮�s131o���K��*�)-�1}ı,O��l�n%�bX�w���n%�bX����7ı,Nw���|bf&bf/-����Q���nʹ��X�%��{^�Mı,K�3�]&�X�Xb&"w���i7ı,Nw��Mı,K������p�a�q�fi7ı,Np�}t��bX�'=�zi7ı,O��l�n%�`bb'y��i7ı,Ns�j\b1ǲI.L�7I��%�bs�צ�q,K���~��}ı,Ow��M&�X�%��ﮓq,K��*�;=|Y?�������X'�]�8-/���u�ݱ̚��-�nn�-�r:�6n!�����bX�';���&�X�%��{^�Mı,K�3�]��LD�,N���M&�X�%��ߋK?��3��1fq���Kı;�k�I�y�D��8�Pt�&�X�ɟ�]&�X�%��ߵ��Kı>罳I��%�b��܊9���[�F�1|bf&bf.p�}t��bX�'=�zi7ı,O��l�n%�bX����Kı_���{!-�)r�+�/�L��	A9���I��%�bs���&�X�%��{^�Mı,K�3�]&�X�%1w���-�Te�W�Ә�131X�s�٤�Kİ�	w��M'�,K��L���n%�bX��u��Jbf&b~�֚=eq�8GdT��o{�0�v�p���ٻf�8g�f�p����L�\��4��bX�'y�zi7ı,Np�}t��bX�'=���7ı,O��l�n%�bX�c�=s*όϯ�����~���ll���A��,E�dTYj�+`l�;u$���f�v�Dİ_˃A�^�����~�����v�R5�T��7Us��)�}�`>�0�s�}��|��4���ꉩc�p��N6���7���&�t�;n�ȕ��·`,�X�ʃ��۞�ΝZ��<]��/`�}��:9s-�*ڥM�N����{:[oGLtP`{r�WS�]�Yqj�� �k\�DB����,��� ��w_ ���m+��nʫ�Ik�z:`{��mgK`ogK`J謹6ڜ
�uY%\��Ӏo�;��~�9۩����Yʢ� �9�|jC�"b-g�g��x��Ζ��Ζ�����y1+0WB䎝�׬����i��u��5��32��Rrg��F�B�92Z�LuY_ ���|v:`v��Ζ��Y+2�/1b�Uk1[oGLؠ��Y��3��l��1��>B�TMK��o}|p�s�L�S��;_b�>��R��wK)]�k��Y��3��&�t��{�x���ה���ʬ��~���z:`v��Ζ�ꯪWZ�y5�t<�ۢʊIb�I4λv�!��<�ق��0�t�vŧXݳ���[�#K�K�p�s��%��z'J�����ЉQ�:��'!��p��]v�f��I�הɓjG�.��7YS��v���v�4�J;O7�V.\������D�n�V�mr�`�7i��a��m��ͷ�ƒ��vms�u�7h7F6�t=�cq�����v���aK3~�����}���M�g� +���1kP�s�m�Y�j-Eۓ=#=Z�秥y�.=�+G���t��	��-��:[WEc�m����U�U�;�n�)�|���������M���zQٍƞXex����$�ގ��A�6l69a���겾�f������;ݺp��u��u�Q��T�ڵ�[oGL���Y��2K`y%���^i�iU�Dr2�aTp�M�v��OX����kL�&F���7	ڸ`;g��]Q5,v������7���?l�|wx�߉�Q��,U�J;)�7���¦�1R (���`@hZ���0�,��7��ޑ��(0=�d���ىQH_*���>u�p��Xt$�^��v�}<���S�%[���Z����p�(0&�t��Il	W%]�D�^P��T�1Sz(0&�t��Il	��\ ]?7�n�T�E(InI��fɤ�����&�F�玃ո5	{*���7���͉�'_�
E�<���Il	�07�Ӏo���
[�c��pݛ��M��P`M�P`N�Y//��ŕ1��-|v��?wn��g�4��U��58*�H
U�.�� �g|��5�53���R�)�7��mr�{:[o(07L������R)
�1	�����;�N��t��{��E,p�%�XYmMi�nчkg�P(��ظ�9�{u��-�k����RK�r�i�?vn���t���N���N���5�ҭ�UqI�[w���voEHV��8@y����kq��)T�U�>�ۧ �~��Ilގ�"&"�}w�,)�`z�t��Ilގ�m}�Q�|asL��Ӏo�f��2[�eR���%�;z:`oE��L`w|KߩK�z��]8���ƍ��A&�����?w�rYͮX�k)�v��t�yZnqs�+����P`z�D��}U��?[���{!KU��#��wn���D�����A��eL�̅,J��!]�C�:,`ogK`N�tP`m�*��Y��*J�$��Ζ�����Ή06��E��+����fbV�����Ή07����f~Gk�-m�	�o�vH�d�,.�3�2�4�r݃N�ܗm�Sy@qk��}F��JZM�0r�ZN3���_F�eNI�NH�[Ŷ��U�t��V˕�j��K4L��@=�ڲ5���Zz��oH�����46
���W%��k�����] ]��j2vظN.+9P�c u�9W!u�X6:uA��J���BS�h�t:��	�w]����I�R凲��;�k��mk��;= E�Z�Mˇ��ۙ���6+��K1#�l��\�{:_������~�W�Gf7y`��8�u��m78�l�>�l΅�S'o3�r�`��&Ke��wg���n�z(0l�����W�f%���e�%l��ފ�&&vIl���j�rW%U5,r���Ӏyg|� �wN���M�R��C���]�n�u��6���G7F0��4u/�`�� µ6��H�e���[�����|�$�tP`l��%_��3�E�]V�Z�-jQ&�(��J�&�  cr�{ѩ&���jI���qu�gv/C�"��'%��n��\�뻽�&vt�L�̋�e���J�I����~}��������p�k�Gf7y`��8�{�0;���'H�����ޤ7�tޮݚY'4:�hWU��lj���M*�:�������6��3�:��u/&O�����(0={"L�Sly�Ud���{���>ݺplQ[�:[t�U��b���YiS�(0=�El�u�T}H�^��12���Xń�"��(U0�X�;I�"��$dI�Q� >#eS12T�	�f����}	1YCD�d� ��'��4{���:H�I$�A��)� $�m�	GhoҰ"$ �"͐H��l��S:�!6� a؁�L�&�.�D�sb�x�G��T*�h�U1 :��p�D�Q	%*���ͧ��=o��-�U���R��+��`{b������A��zJ���f$%K-%l��l���lQ[�+.��������$�h.x/d�����gK��DuKc.��-�le����".����;�t��lQ_�XI���'�����mG^7U�U�>ݺsٍ��}�x��>��Ӏ}�[�ݘ�i�+�0={"L	����A�6(0=Ў�a�X%�#V���-����w��Rx
�х�?�#` ��(u0����y��{��/�3r�T�R�k��� �fb�}������ogu�����-��K(��s��]v/�B݋\;WcV�3�a�Yq��0��N����e�MK��=�_��u&��l�07L�>��Rĩ]���Y�~����D(�9����ŀ~n��g{��d$��Z�mo�n����هDL��|`��g �iKe���Z�J�1+`wE�P`l�.���ݝm궲����J�۶��Z��7k\����"?D!-��J�d
6��%
�!�=���s��~�C�g�=z�.2��J*��vM�5H��� ���=�zAY�6�6Ѷ�v��n�K۞�/Z^;k�I���:m�c��;�����a��N���&��̪[����L;��a��{)�s��V�Fx�6��mZ�N-v{!�'C��Y����"x��Y���RL��/+�p�RP�Ay��W[���c��Z���=�������B�vX�����w���cS�x̂�>��r]ŭ8�I�!�X"�&������6����qI>��aH�G.w�����:`zE��,>+�
I,�vt�oGLH����`n�*,���ZU�������	���P`v��;��|��O�2�H�-�����8�����Z� ߵ��>����PX�+��Z�0;b������8�۷N�5���Er7!*�gmr��.������L��v��ԥ�]��,c��v�6��}��E,����vt�oGLIt�ĳ3��_W�;�?(����T��8�n����ѯ�>A�S�]jg���R>�m���ݝm궲����[0="�^ȓ�:[��� ��l�Y�
e����{��o ݛ�`{�:`zEoR"2��ľĭ$�����%�%�0��T���I��QB��h��^�hK�c�[���v׍�����2�ZG�<���nĒV�����[��$��Ζ����v
BʬD������$�L�-�� �>��tL���1SK�-U���_ ����������4�t(�����F���=�&�Ӕ���X�����'�wπww�\훯�~�;�p݋aԬ�T��J��0=2K`n�E���l�b�{�֜$��ƭ��UCR�����
j��ї��{a�MuإƇ:ͳq�	�l`_
������`n�E���l��.��6;*x�X*I_ ��g=#t�p��`�79�&O��:�D%�#V��'�`v�t���-���v����G+�E*��_�D�}�`uwN�;w8�>��EB�!<�bBIso����u�uBB�IW�I*`zd���+`wgK`{�5�]�B�Ycj8�U�m�K�օ���l��{$��ε=;v�]�v�s��t:�ϑ�L�]���+`M�+`wgK`v�t�����|�k�*�V+���w_ ����[�(����0ʹK.�*vT�����p�n�ŉ7���|vo� ��oev´;�R�U�?:np��:�7k\�tD����>������X*I_ ���o �$�m���ذΛ� ��Q
TB�(IA������ D�+1�lT'��L��)z��x�}�V?�Y�۵h�avm�v8V�Ƌ���|r�˝�z��yͣv��%���74�@䒍-M����[�쪮5us�nU���)��c)����n���dۙ[m��qm�e���Ӌ�uΜ��z�#[�;\������z7!!Ύ�og���uZf5�������vF�pix�v-�Mά�a�$$����ǟىb2��͜p�B���.y����ڙf��:�:�U���Ƹ*�瞣*�HZ��KR)-4���|���s����o;�깊��TӰ������s�f&�ޞ���_����>Ӭ�ʢ��ڸ�Il����Ζ����t倣�+-U���_ ���8{;��~ގ��%�=|J��^$,�$��ݝ-�ӣ��Il�����(���nwf��;<�OMLA���aa���U�.�����WZ�/j��7CsR�N���%�:r��:[�#{k+M�uJYW �f����Աt�PD$�aO�� �s�|���Jd�����NF�`�%|{��~������$��TywG�bUEX�H�>��8�^,��s�Д��� �k�μ�K*i�Ke|��x�ݛ� ߝ� �k\��(I/���ER�S���sl�k��Y�����۲a�0�L��v]�x��8�u�T$�ʪ��ھ��~�lP`ogK�z�dT���L����*Wb�J���ۛ���H��f��>��l1�@MG%|�gu�I�y��U�VH��ƻu$��L`m�+2����^*I%l�0?m78���(�v�pu�=E��Zn�Rʸݛ��{1,[;�O���������޷�B�Uc��n����L���L�Ά�g�j/j�9z�Ғc��#B�T����vpݝ��7�:`{�K`{xD�(��J������ �^,~�� n��t(��^�<��%v���[+�����w��|_���?l�����T$�ʪ��wk ߩ����`:�8rJ)Dv,Y��ˀ}�=�����B�_ ��cft��%�:��kM�`96�.�j�c����H�vzԕ��)��њ�g��ۮ卷5�3�:�8ۯ�SsВ��:�_�)�(RU\��k��n�����l�|����ٯd��V���IvIlH���Ζ����+����]��f+`zE�t�w(0=�%�=���2��Ī���$07���;�A���-��J`�7�7�Sk�U��+0���ϕ�F.kH�qtgr�ɯ���BE"�����`�$/�>>!�� q��6�ר���m*�f�1��TD�B�|�>����tnjc0d!��|��\]��� }�@a"A�2,X�@�LdI��*�z*|EC��O	0����U_���H�O�o ��0�"2(c �&� ��"�D2&\$H	�$#&hV�� D��J�J �Eb<}�Y�q�_b�.o�օ��&KI*""%-��۫��;�����m�� V{���s #�=�[2��p�����8�֭S`ҙk.$�C	`����d#r3�(���!.���Z֢c��$�v�\7+S����.���I�D�r��u�r�T�utc) KM ��%�yV7i�
"���_+��u�/eko*&+8�um��0��ذh�nZ��N4�_�}����l��6�����vT�:iX��j�!m� �m��:'ۖ�ђv��<�쮬�V:��7c�y���{�.�I=v=l �e���ҁ��b�n
't`�w;X���h��ɰ�cD��28��U#L�!%ظÃ;p.
{m��5��<LƱR\a-�f���+e;5��[p�4x�9H�s����u�Zg�d.* rm����Yx���9{[*Ҡ6���ũu�a�a!�5��Vɬ�C *vk�V�vH�UBj�{f�`��Y%��F��Zm�)�N�ևzs���3��x�����u	���eP��Q�F��
WYy:M�o#��ͺv������aUCPp�Fج�+��`a���l�J�ۚ�ݫ��sM�ۇm���{3�\㇁�)wk{;�e\�����ϳ�m��(��J��8�dɾ�#6g�|貆ݭ���@��ݝ�@����VA���6���b�4��vY���6R���By�pQ�{Yݙӝ�]�v�[�>p5t�=N�.�H:��(�uq�{u���A��[�#N�أF,u� ]r�n��V� �cR��^�C���ܜ�k���ͰԠ��й-*T8#�o9P��h�e���gt�%��ǋ`�9��=s�a�ǎ��v�%u�Y���{e��N=�Paѻgv�T@j���g��ϟ]���6��6����U��ە�m����s��D�5v�%�ں��|����\/=::�؃�H�9��
��ؚ�~>~D7d~&��+���b����.��q*�8G)��Q�t���c�A(mЎ��~@*@�(�?'��h�W'����,7nJ�E��
�G��f���m��	�9Mm�7��7/$Gm�8�hS��u�.�ۖ gk��'S���T�����z<.��|��c3u's�Քm��+�C�Z�<\�02��K�r&)��XL��{p��u�:�m��5z�ʍ���GT\]=K/i�D��'<��zM2Me"u��v���el#�=];,C�������X��9������NF�zt�� �	�t�l��ﾂ9�%�]�c�o.nΊ8쮼�Wj�XKe}�}|p�$�lP`ogK`z|)Vf%��U�$�vIlؠ��Ζ��������{�qR�UmJݯ�o}|p��l����d��8فRϕ��#-!���-������C�~k���%r��V�_ ���pP�����k�p��� '�7j���$��ōs)��=u�5�:^�i�;�"��s0�Ժ;�ͪ�m��%�;rK`ogK`l��%�Aj��hV
�W�;�n�{k�3H�@E�U��@щ;�owR�o��f���l��� �-He!%l�?[g(0;rK`v���9����b���b�V���vM|�����O�wπ~�X���-��Y�K���-��cft�w(p݋�
�P�����n��B�:�y|͛6� n͹��ݗ����m�u�\j����R��Wi[�$��Il�P������> i�L�2���(����7_:"P�Nn������ٝ�%2w�z�J�%Uʭ�����w�v�x�F��!a�U&���;��o�|p�׮[d+U˄��������-��(0:r�{%�Yj輻����l����A�Ӕ�7_ ��:��G0ʢ�A���z
�֔�]/G��˗�&u[K:�����Ī�)b�l������3��7H����JҤ���L�����-�Ӕ�A��K(R��K1b��%�`od����	�A���Ӏo�k �Y,U�+v��fdK�`���5��Q
�D�2">�'6pDC���{�RI���	XR�W�b���(0'M��>��N���٪�؋e�Օ��vݳ��u��g�hS:�ƫ6��\��)�Ҷ*ʵT�f*W�������[d��ۧ �f�r�!Z�\rZ�8�ns���z�Nϯ�~v��k6��C��X*I_ ���8�n�9(���|`�p{/&�"��$��,`N�ؠ���[nt��qe���� J�C�(0'ds�=w�=v��!$�5�W7r+[g��9���s�B�8�Gj@�;v�8n ݴ/S�<��������t�5e��a�D-�����H�.Rf��7��I-iR�7��t�v���$H�u�[ZgӉ�wC�p��=�6�r�DV�V��۶*^�6�(���n�@R�{�����vMٳ;Ži�:��0����b���SX#Y ��O��|vU�	w׷fz嚋9��)�L��DEp1s������:�E<�ɱ=xsמ�����[]���8���98��o�#/n�댴�p�~�o�?��-������(0&�e��[R�k���N�$�������� ��u���t��%)S�(!�'�Θ�A�;$��P`u�kR,��r岮��t�ٺ���Ӂ������ˀn�?9m��*fb�H`l�-����:`v�����m
���I�����{��4�M�X�5� l�ni�kb��ۛ>T+�{v�#1[g(0'H���K��7��a�Ԅ�� ��ӜXj���rP`{�K`l��-Ew�]Yj�b��p�ۧ �����&��8��� ��X�Gu�Z�,��vIl�0'EȠ�����Il�V�n��;��.�ė�����������n��i�P���v��r��]��-6A�]M�p�R�.�^����R�u)H�KSrU�7�t�n�0���P�H7݋ 5���.�Uũ��I�A�;$�wGL	�A���׮YdErJ�%�Ӏof���;�S�>!PBb�0���q�g�RO��qp�����7B�T�����`]� ����B������uG�ؕQe
�S�(0=$t�ْ[���pݏ�����`TJ��)і�o�Ks�9[�=q����
6���W�/k��%X+1$0=$t�ْ[����f,���﯎�Z�_c����N�*�>t��(�26� �_��,{лX���X�r�k��w��ov���#�����]�*�
��35k��}�`�ذ���$�"!ZAr0�w�{��N�����e��^/�H`l��vIl�07�t���↱GkU5e�WA�Rz�޸x�9�/6ٻ��DFqK����v��� ��Ufb��L	�%�;�t���w��ov�'����+I+���`]� ��� {M�r��9�#x�[�d��{}|pۻ���o�=��7w�\{�ݭ�t��)-���� {M����D%<�8�7�����ae�p��|��`N�I0:��������Yx��e�.|#��4��<����Нt�k��}g�Wn7d͋�6;'��v����ح�w[dw�M�`�q�]��]�=�WK/I)�3e��Nړ�#!�ۜ��p��ɫr��}k=v�-���۳f��g&�;Wi���|���=�F�*ɵt:�DÊܲ�NѫX�8]]rv.$�S[��͵��̙5�͌Z�ߏw�~{����&�]����ٺڰ�#��w/<����Y�mQ;�]�㍷&�;-�mL�
�b��ݯ�{����N�I0'd����r�U�Uu����L	�A��#����0�EJ�f]/���,T����vIl�A��λ��,�`�Č�T���[����P`zH避��'����+I+��w��or��GL	�%�2��J�u33���k����ӵ�	%��.�a�n���`���=c�uH�-vF����W�of����ݜ 7w�06WZ�_ً-/�a��f�I���5�z�Z��;ۨ��.����䱳}���KP�uuk ���7u��ֹ�?6�`x#T�RX���+������uk��o$�Om�N��"��WY���T���-��#�ܒ���. j��RL$��6d��ݍ
Qԍr��]۬���9z�e���]�ѫ���u��
�|��=$t���-�����wg ���{+��+��U�?l�����d�����]��ve���f+`wtt���1�ꯪ}�SN#���`��! ��KI D�,)1(`-+�\&��P8o �M�fW9��k�n%B���!� �`c���U�0d��9�w�:CG#ĉ �I���2B�L:�LI%�/�.7�� o$���&���� �!�j�U�8�4aAC+���`3���g8�`�$#%Y2
�!�%"��Pv �ޤh"j�V�`2�AL h ����"˔�XU��T`��^9=���3@��:�N$"��(��L��|ސ]l�0�T�08&
M�0� d��P0�`�
$YI$��$�k��Gj�~�A��W,��A>b���T�m��tZ�C)~�H�2��`�6	FA�x�T�m� ��V�$�����,~�� ײ�n�f&*�%�v`t%�{� ��ŀ=����fbO��<pn���$��R��-,`n��;:[v(0%�����kD�GrB � �K[V&�l����� -j�3�^�eط����K��2Ӛ�P�b���lؠ���g��꯽a����}�{���e��+v����0?7X�7� {Z�9L����
���i�߿cvGL	�07b� �\���@��x���#��X�;fB��a)@$�F�B҅Å����iZ`�A�(q"�*A���j���?�{��~�k=-��+��U�7��Lؠ���cvGL�U}u��_�-��YX�^��6��Y"۴F�Vt�5��Ŏz�(��C��W~0n��9���>��]	G�o�`���dm�R�)-8�۳�KXٻ݋ ����f �K�71UeݫE�2��l���:`l���p����Ic����*�{1'��z��/�^Ɍ�06KUff+��R��i*`l����:d��;�RM�lH1U���#���o�=7.�60�K64 ��g��<j��]곮���´x�g��w+���4��X�n֋�;=�C��[���]��s�ӎm�D5�`tm.���@ȳV�f)� �s��i���euu�Y%4=�݃=Cȓ���:m�����WIU�v��i�����a뱅��cg[��H��	�M�;�geK���s�@em�q�
��Ia(��%iw�[��Ibj�;��=�R�'>ݤ�і)�-�n:ґȒ�����j۵��(#���qG:�mq�ؐ�������0'tt�����z�j�PW.7,�����7��.�{t��n�f,l��G�]��IX�F^*`~���P`K�1��#��]��]#hN���~��8���:`N���*;��/�/��e�0%���H�;���(0;�6�h%��(����-uPu�!ò������}���]ͪ�ev<�<ݬ�]4�C5���K<�ߝ0'tt�����p���$�;jm�W ��x��T>�`�O
���Lg��jI��{�{�t��,QU��RX���+IS{��L`{�t���� �޺��R�W�b�L`v��;���n� �uR�Y*
�����x��x���0?7XB�]�ʮ�K����Ǚ8�m�m��P#K�dpZK�<:;m͙ڢ�.X�VF�������06r�^Ɍ�0'���ʼ�(�_"Ҧ�P`K�1��#�eGk2�����Yi	{��RN}��ԛG	<�#�**�^G@�p�=�jI���MI>��m�#L��4�v��ۼ\{���9A�/d�ПZ�f����eݬ�XB��~�{� ����;؟`MP$�7jI%W$B�;w��ڔl�ݛs�J嵶ź�9Q�S4��ZJ�ܠ���c�#�n��*��������c�#�ܠ�;�\G�Yx����0=�:`N�遽�	{&0;�CamU�%b���\{������jI��{�I>j��E����g��=�p��=H��Bw(�\��f ��� �����ŀr�v#���a�랸Mۧsנ�kOj�V<vZG��$ĵt��)P<�0���n�Iv~�{� ������С~������ּ��	���p����7��X�m� s�u�
"!D�ڜ��&��%�v�T��'�L�P`K�1���a)Eee��b�Wx�%L�P`K�1���vGLN���T�a�b���Ɍl���:`o��f��-F�����w���s2]מ7J��v�PR:��XZ����kbH%e��������I��Rdإ�:�Ku���<s*�7aGFCl�vd�;�A�]9^��#u����N�v��d�9�ǩe�r���>�9�:"��tR��ܷ-u�E�a<�m�qy�@gtF�W9.6��T!s1�ܾ;\�yn�^ll�����|�s��^l�u���e�G8�v�����qY,�G73"K8�,��,�\��U�{΍�=;�wi�8���s\t�k;=�f�<�	�ܜm3[5�r7m�g��~��:`n�遻���"&e����e$��07dt�����8߷x���H��ԋj������1���wGL��YW],��B1!�/d�쎘�:���N�Χ����	���p�o �^,�����與��A��n��sUC�؞�9���m)v��9������r������}˶��LZ����w{�� s�u�P��!��ŀw�e�b�e��[��W ���9��b)	H�#�+��#*T��A�
�D$BU
.�����X�x�^�\�V�+�Ć���0'tt���_Jȏ���+�_e��I0'tt�����""ŋ),3��˴��P`K�1���:Xfed�����G�r����D�E`��z��l٬�[-��sI����D�lr���>�n�^Ɍw(0'H遽ҙ�*�륟
�����c��	�0=ܠ��β%+��**��ZX��r�wM�,��Z%�@"� @ 	 ���m�8��Ӏ}����2�lM��Q�;��o(0%Θ�����Yv�G2�b���w�n�^�g ����׋ 脒|w
���TD���U���q3ʁɛm���=N��WM�Z�n�LM/1�\�FU]aKS%��y�}8����:`{�A���W*��3R���,X��tt��GL�P`I�>�v�e�+T��Kcr�����;s��$�-����N�y��w�`Z�0;s��$�-�����)�"FXpF��*����*��WP�Ͻ�RM��51�����J�rL`ztt��#�N��������JԐ�;=�����֊c�[���V����K�.�Z2��Uy^9jd�Y�������.�Ӻ��a������~$-��;e\[x��I%2=�Ӏ9���?=x��yAW2�b��嫀w�� wv&�GL�:`Uϰ��������
z�����,��`��_ ��SԈI(*ܹ,��}�� �@=�{��'o}s$�}�gRO��
���_� �
��(*�AU��
��PU�����PG��B
���@T"$B)P��T"�T $B(�T"�B ��B(�T �U �B"�B(P�P�B$AP�@T @T#P��T#P�@@T!E��T !P�)P��@T "�T"$B0EE����T" A`�P�DX�1PEEV	P�� �
���(*��AU�"��A]��
��PU�"����_�����EW�DPU~DPU��d�MgPX��f�A@��̟\���t �h(PP���t   _{�
  ( vv�4 fiv�vPl z �i� �
�4٠   @t  �    ����M� : ˗TgAA�Ph     ���  p  �(@ �@�ܠ;o��3��:��w�q���3��y��v:U�{��>쯀پ@�{�_ 	�>�@��w�h�;0	�}�us�p(+�>��������uU�s���p ��  =
g�  ��CK�}�w�ڪ�ۏTyuNkt�o@	n�����F��}�����;3�T>��u�w�u���h���z�>O�������n��n�������C�vg`נh ��  ��{�
> ���f��n�ת>�x	����7OC��OO=��Z{�g۪f C�70���x�z�{�=<���[�����>�s�݀p � ��   @��O|���<�� }/{�tK�M�m� v �ܦ�AҔ�� ��]�����G{�@�K�� ����R�zts��^��zS�K���JY�����OA���i����t���p=4��e��͝4�X�� �   �  ����F�t .g�@�: σ�s ؠ�K����}�p�6S뼠z�o���l|  C������B�w�H{�ްtݍW��}�ow|��m������O�iM�)*��db41تT�~��  4̪�x�T   5=��)����F�OѪP�JI #A�����)�@G�z�������_��a���'�������@U~j��U�*�*��U�`DW� *�AO����W�:C���n�/J�������܌��%�	���.��^.�
�zJ�E	qr�`��f�,J�ƄX���BP��f2�J�f\eH!!XXP�eIYX��%aYF0a5�1�#H\I��^FA�I�XV��-�1�!���`B�B��\#RE�,��!HBI1��I8��(�J�)��R��&$�+� B��X D�B0d+
��9L'������$ 0��xm�$�HLB*HOt&kA.��2���P�%d� D�!RaB�4��.h�ə�p�BJY�d��.����r%s���K�7v�ɚ��M�i�	�W�x�\u��)%��Ř�扄9svj�)|7�<�s��xY��C�c�i�u%��۬;yx�t�0D)�
A`F��_My�GFFkZtl!W��"��n�s.���6���HabA��@ě�������\Ըy71�a3{.��p(�R�#d�%�%�);��~%ܕ��%��o�I���7�&�ٸCDZF�)*@$k��ӄa5|��r��ni�U=G�p���{�p�C�+�A�Є!LW4�(J	��k��X1�s��^w���ϲ�-���eo��Z%�<��7�:3��5��oL�5J�X��!$$� �$B�	@2 �"�RH�D.�8A��!P�F��%��S\e�B�sA��$�
񅝜a,ga��"2P�dn�4Jb@�)��m����N�J��S3y��ԅ==S@�
�)�ԒHZ.V!%��9����=�'����v�����w0�!45tE8��W3D��s� s��@�.C!����\\��H]������HH� �
H�e2�F�4o��3���!׆����\P���sM϶�'>}�4F�r���,.�q�\e���	Yp����2�sd��!�������5�I�	�$��FcrbD�+3�Yq�e��c΅FP��%�3L˪fnoDּ��G��J�8�g5wu�95�e��P�D3	RRT��!�0�P�BP�57�4�l�"W�?�AlX�Fd�B���0c���I��d���+%HS	r�e����k�������Aϩ�޽����������xB�P�e8±���,��J0��c��0&y��Ƭ�0���hD��I ���4�� ��澆�9�%�P����}ﯬi��H\L\	p6�.�W43D��IL`FQ�FP�Vrfټ�#D�� �HR�"@��
�A&0��n�$�+���B�$D#��'�(@�*F�)$	���c��"@�\��d�G�� k\]}sD*�\%�J}�<Ռ�������0��E h�4�bR426%���VA�@b[ ��\L�J�
d�J`ˌ����8��*y*�!
��@���k~lvo[$�Z禍ed����fi��<w��쐈���!d�Y$n$�(F�a�5"�`2L�R!D[�
�[�}��Ҙ�9>��^�(��Y
���a!	ny�sd�������3Di���&�JѢ$*�F!�h�֦��4B�Pp��d���P`�H��LeaR*��Q������G��_P'�'�f{g�3�G�I�7<Y�a7����FL�K�U����>wÉ��i��ab2]0��uJy�&���h�s[!BH���F$),�{~Ͻy�>��N��#!!)
BB��m�������lXƱ�� �Y�c76K�[B�D!B�ޮ��1�%K��	r\��U�������)�
��*�@��-�n+��+� �ZkE�2Rda	-'-'����˙
�������΁��.(K��!����F���ʓ)�,,�߇��G~�e��.G7�5�s1���N�/�+.����Yn��I��˚.i��50�|�qXD�XM�]�}fp5��3�sD.j1�1�0���Ӣ莭�l��c�!H�7�Jd�jf��G6J�0Cʅ��̖�����Y���9HF@��-�ә��frm�p�̅�&�0��� J��3�G"B�A�����:�Ņp�L��
o[x��Hr��9H# Ĉ!�Ih.��Úך��{�i�!t���HPi�m���#SLJ�8��Q�1`A��$xC:�����p.����'4��h�A��.�uϗ����	r\�<�ów�.�8��##�P�a�IF)��	��!���!pjdp��$�bH�� ŌX �	u�|<�o�s�+�H���$H�@���=7��@��'���J�$�#$�B�	0�a��W>�����5ߡ+�a�q�,���4�|�~�!VD�L.g�ާ�4r���'���|���I+!�o9���gH܃XHC"HV!0aLeM�7�\�xC�>מJˌ�Bۜ�\��J����	A�`�$��M��6B#
F�$1�5�:<�!%���D��֙|Ѹ���Di���ܔܦ����9g�����2
���c,2�%0�`�IRX\��n�Y����n�rt��Vp�/+��U�������5���y�|w'�̦�)�$��XnS��	(JR[���)���wo^�g�O��������]�o���!?�������s\��^k�Ͳ��71.\������p�VD��B!ȡ_L��o<�˓�H���Ń)I$�)��	<8O<9�a�І�Ofh��vy�aJJ�3e2!p�`L`A��!H�c`A�1��L�]d��Ѽ B�����z|ӰX���zN��0�S(]zsf��)CB�NL��7�o~�k3��G�:���ܬ��j^p�	!!Kr�d< W�!I@�bE�ИSZ�ѣ�Od"dj��{&�&䌛�4�Ʋ�� �`Xxp�G9��bɱ���bԅ�eֽ�	Iq��6R2�0�Y0���Ԗ]��
B��|w�l�.;Ѩ��aH@��!yÁK�[�{���oS�kL5�,�y.�z���
H@*�$�#]�>�B���"�	�H1���^������w%g��/���M�I�T�y��.��n����w�hI!1aH���,�i�0��$�@�	
`B�
�"J��.�2��a�|��w��$I��HY�K��g	If3��ׯ��Yt\	�.	sDp<C�޵x�\&��z6^�I.�a��iɪ��\��|*mg{�zb]��s_|o~fUQA���
� ��R���Gs����o,��[90ѾZ`] HH�����$is&�!`Rc�!R3�cǄ��$N���R�����wT�D֫$
f$hB(B����yw6]f�$ܺߜ���j~~�q;468w�����m��.�a���&���zg�M��饲X��u������Fy�m��. Li)�w,���M)t�`nR�ѹ��̆[��InB�(J�H���ā$����fz�jS��9}�[Z���ŋ�|��
��\6p�_�s57-к��ڒ������T������K�]2��i�d�+�ŅxC�4�|�3D�:@���Ie�\���;�?���'&�I<��f�>|��x���a�h��h�`�d!B�h҄)8\0�4�!YLap HS+V �2�&R<)��eȤ�V����p X�E�HE����.�C�+�ZHIe�B�Le��F�od�F�(F�I��7�şI4a���$9�M޸�.�ˁ�2oy��5W6LR��%��	_R���	��oճN|�px��E��Ė�YogJ�/1%��SIat�%��H�k�27�W�W!@4B���hX�dBI����H��H$7cB�HL��yy��3d7 `�5�a

F$�d�c"�B���8>�'<4��bB;,R81�#�ZL��c3�]��Mnxk���������������˚J���-q 0bЂ��#@�� ���F^�Il$ﳪi5:��z6E�@I9
1�
B�h#"VFB@���i��Q"BE1���p�B024	� �T�HG߸BHp|`�%!E�4)��B2$P��"H�՞�͓�B鲴�����IV5�!M��Đ#�	��������9�6f�,7!�*��&�f��d�-$�����,�B�#9�!E$1c0�+
��j�B��M$c�$��4�2�:�\u�1%:���eL�t˒�3	B��3r�������n���,�s�,��^�<�&��ոa��C	!FH������
�X0jh"�A�I�{��0�H��e/w���ׯwY:��z��UU UUb������{ު�ٵ��������Qb��PU UP-"��i���@-��-���J��UUUF��8��*T]��NY)jU�i"j�6X�ꪪ�k�EUUUI�e�
�t�`*���]R�UUU!5��U[TR��v�e�k��V�6v窪U���*��/R��T�%��[�l5N��kd���T�K�T��PmWU�S���tP UU*�mUmU��݌UUU(��UV6�M�炠�{�| 媥vk��n���h�qUT�*��B�ȏ��UJ�U�UW��Z�A
 �iCa�����Gd;m���A�Vؙj��	��X���M �4�nt˴!�ڻ$R�ut�^iV��B�vZ��U�*�UU��&�z�\�0��������� vf��&����UUUtpO+�U�R�U@WWUWUU��� �Z:���j�UV��e%eP )YUe���\�� U� �i
��X��V�*� ���2�Z�	���u���ꪪ�&�袪��G˷�6��ԫ*�e�
�U����(8��a-�U⥃����U��j�;���V���mJ�jD�SEr�6����[,��(k�
��Jlɭ�ԫ�{iRꪪ�*u�Վl�g �Ac�*�@uUUT�����K�\bަ.69%�s�QE@.̭��mn�UuR����J�5�[T[�M� *�����V��Tʡ�[Uld�j��Z�k�Vݠ@궥�gv��]UU)-)hE�h�t�\;�T�l"%lt.䗪�	��OMKɀom�j��EU*5T�!sUUl�T~����d�j��6*��S�Z��U�������j����x�NВ�U*UUU] �����U��W[+ �	���L��T��+���mUX�T-UUR���c�T+5U�U�S+U�E�*�`6��S[UUW*һ5WT�N���X�j����Z�
�@6+�V�������V����3�uJ�=���
���j��;V1�\D�M�UV��U�UJ�ʵUUU~�ﾠ�j�����&�����e^�X
�U��檪�����U�n��6�`*����uK�e�ջ�@T/�e����UR�UUvʵmUm�UJ��UUUUJ�UUUUU@TPUT����e�Tr��AP�Q�U�Y+�j�U� mֳWh��{M��v�UUuR�`�@j��X
U��� �������#/9٫��U�V�+��U�U]UT�UUUR�r�UmJ��T��*�[U�̠l�gK�T���,�;TJU�T*�b�	 %t�F�B�6dVN�ir*���������CF鬣UUUTU@V���/��UUU[Pm�,횪�e )�;�B������v_)�7r�-2��s�S��7F�6��7ei��K͡��q��]b�o(�*�J�L������歩��=��-U���=y�sp\�p�UuU�Ԫ���dAX���Z�m[���U�t�c]�0U�Q����l�UUUJ�0R�������P��ɷ@5U@E�\��u��%J�R��@AK:���y�ܣ��N����c
N�h��������+m�WZ���3\ RշUU�ȷJK���+���h͛h��F�Z��:�����u����Q��3G�xc�S�U\�R����Gn����S����)nT)�Z�m��sШ�k+U���8�%d�r-��ܗ�z��nV����`���Ak���Ǫ:�4��n�a��9ClmN��5+��/� ���@SsQ	v�uEskj���
����V]�^zl@UJ�T��@&�e�-U���[J�n><s}³A�v�m���<�Ƥ�hn�[�v�J�\9S��jT�ZH��]Oh��:-�X6A��cj�袪�*�ꪣ�PST�,��]+�T�WUO+URA�]d�M�˝%�eej��(1�:A�SEN4�W�ڷa+����sJ'R������ ʵ_}�}}v6*�eA %�`vvܵ���'=E��kU����u��/��`��t��%T�5Jҵ��Wq،��ù����f�HZ���N���I�R�R�U��yh8��V�yZڪ��z�ڪ�\7f%疪���B������8j��� �UR�J�үe,TVa��j�����
��<�����S��������
���&UtQ�w����Ik�N��G�&���ʭ@uUuU�s�AJ�+^�ֱ����鲪��m�*�R�UUU,�V�A�y��������Ĳ�e�&��$��UJ�UUҒ��!b��UUb����UUj�kP�UF��ڪ����U��U%���1I�.t:ӡ����ȴ���p�յ+! 1EU�@U.�dh8(�����UZ����U)�n��Q���dA�&E�gwnUq�l�[�g,�c,��/4����+0��Ф܈q���2�յ]U�^y��WT0�
���\J�R�U]]PTr�-mOWU@l��	�3$uWUE�P�s�T���c�3l�`�v��ʂ�BZ�U�L��6��<��|��C��dѡXD�f�-�A�k���-�.����!FH��
U@ٺ�v�����1�a��Iv��okm�B6
g����.�B	-�����ZU��r��<	cV�k�6�4��k��a��=2�B��K�e(&�j�twI˲㛰S	��� 2�Q�8���O=����U�����6 ��ڜ�TnN�i힀����it���a�*�\杳,��X�M���<�  ���;ex����V�bK8u$gI�ʠT��r�PWqC�/GY�l���[�����kt�	�d���6�XA�`�c,�MA�GUt���_WP�<n���\���*HK� 5WUHb	`E�@P��a�,�%Bۊu�v�cP�-R�9����Ԯ�UU�[c6Cvt�!�����R�5Uu:8E*��[��� �vӛX��ð����j�����$YC4��u���PۢQ�E����g����B�Tj�MrW*�S��*��*�P�!��U����;�8 {, 5�/<1J�=�%L�r��,��-UP��تڪ�SUUP��[TR�P�몪���A̅UUP�����*xb��Z`!h�b����T�e���n��7�=���m�m��]�e �:l�PA���[1y�:��U���Wd
�U����U��UX���~�����=�AL�VԴ�\m�ۭ�{U[��[������jU�������x&�4������53;<�c�We��TUUUUUUb� ��TY�ʪ
���u!(R������\à�D�[U]��W,�L���������H ��
��ڪ���\Ҁ�K*�TiEV�UZ�*������6ЭU����U����UW�R���
�����Uu���V�R�Q�s�Glu&�� UUU++SUZ���r�n�UUm�GC�%Z��e�Z�P*۪�n� H��U@.�Hm� \AUUWC��Ж��5�\�*�T�hjV0q��V�u��.�5�UTUUuV*q\�̕�0(6�L�j�ȧr��%���WmN�)V�Z�*����j��턠f�[Oh釸1�qh��j�������5 R�UUPSUUUUV*�0SUW+UJ��)K��Vꪪ��U6;b����@���U�����Z��@jP�,�uU[UT��{8��� +�RԨY#h	 UU���/5�rEqAV^]���3ضـ�j���US�&�8�'gEu@WOK5E#evR�P%� 6�-uHl���Y��� ��f6�M� c�X�UM�� D2���WiZ���j��n��ڪ�m*VV���ڹDXj���ꫝ
����=�+���umR�
�g�Wh����������聈+��3d!#+�Q��ɔjf�\�؛T���&���Su-F�
���"V�Vq�ek5T�ɘ:;<v�@�r۲�ݝ��ΞJ�j�R��	ݞX
�\��,7A��Ǌ�����vg��qD�M�c�U[Q���WUUU�\q�T�u9Q�VԻ`�J�m(Qġ�R�UT�aI�Z��L���*�HB�H���)<��]� U�Sα�ԫU/[Dd��>��]��PU�;J]�.j�A�f�
��cY�9۵6�Ch:Z��V�jU�..\��˻WU@]��i9m��muU�[UH�� 9۶��Y�"%����1wE�m�&��B�v;tl}��H
��1:*�Nζ *ꌏ6�P�EUUP�`��/�TUUUUmQ-*���J%[�U�c��t[T� �X 
��2��f���Jq;s�	Ti�������w�i8�T�(8����zڬ	��T�r������v���J��@V�Z5�����6�J�[PUU@*�Y$yZ���P��UU �UU]J�UUT��U,V�V^L�U]UUUUUUmJ�mK.ܴ��]JKUUUlKKUUUV�MR�Z�����Z����U���3ԫT�`
����U��k�U�
����8���O;Zڞ��7�)�U����[��Kڶ�T��7�':�Xપ���
�V�h�WIc�������^�Wv������/��q����)j�j�A�dZ��V�����j�����U��h .���PB�(G33k�"�AvΗU]U�j�UPe��T���������UHu* A��UUUUJ���V�̧5�i�I�
��I@���Dݕe^���UkjU���u��LmUUUUU�
��,*���9�Ul�UX���))vm�)����N��8U?�AO�G��
��@�D�?�U�0�ீ" !Z��T��a�qU6⾢"�� )��ں6��lx*D�LO�'(�(`D#�)O��O� 1d����OA@6��A�|(�������/��x`��ؐ0�0��Pb� D"�}UN &�����?�A��A���\] z	�U� �"������!���W���D��D6 b����p��C`���r;� r��UJ�Tu�6$~�> 8_P<@�� @$	����� H��C�_�����G�N'�z�� B�B2D���|bU0�8�>>�}O@_��_�#�����lEl�B�� j
*��b �}l �P�x�	�	�"@UW���pDW�?
=PdAF(@ID��
�b����t�N���z=�FU^�q	�$�jc<Xʠ$G[O'n8$�5�ҫp�6�H���Bd���*N�;�����oOnyU�E]�v���B�ma��g`�5���J�mL�d�OD�)� 8//#�C�ܻeՅ��.*݂G<d�K��;[	���#z�����'�Tx���z���)Cn��Z��j�>T�#���ύ�V�*��j坌1r��.\ �L�me�;<�P���� 	*@JU�6�Du�Y��[N�5� �V�EɎ��A���M����\v炽A(�$��b�5���r��k[�\�̙� �誨�\�a��񌐀�[q�m��-�%e���8�V�q�9!1>��D����8��n8O],�xD��^K�&��)��ʠ��4���IOfx5]�U��X�"�.��t�hm-e�J��P �-�9('r����f�0N�r�q��l�M��V%!�-E<�7;lh�
��M'l�����@���
�2��e{`�͡��ӣN�\m� �b��f&����-�df�k�9Nz6� �m�]nާ&��ɀg'`�]���|�=����lf2�����s���Lm!I�q[r6Ru�7�`Sog؍X
�1�\y���q;Z���&y�%Jvgi}�-.��ga����&�(�cm���v��dZ�fX�z3*�)5�MtBK�����s��v�1l�u���
�\�5;��e�.����^p-R�΢�T��� ��$��t�roQ��\R��pB�qv�00�L��w0� �)�.� 1w<k�7g��U���-��b�旁R�氙CE�����lN���h��C(([8Ӄ�w
%�]���v����$�e��JtR���Ά8v��nG�{p���e�Cv��Wvin����� )�Ү�D�PR<dz�@�#"���o2�좓r�\ε�EҪҨ 5�2��.ή{Fy'U�¸٤"ݱu-ȗ-�p���wO�����I��6)�N�~Ew���!�'���('���奓-�nd��Fa�kVV L��*�t1��s%�O�m<[Ty\��̕����ِ�e�
.��b�@�,&�J�\1�T����Mv��N��Zk�mw�)ϓ mn�;��7f�3��L���oCi�hi���K[(�D�lJ8�6�r��c{�S�(��ӣ���#h��P	�L��װ��A.V颢C��t�ӽ>��Ը& ,.�MNŲ�c����#��*��/���.ʷ��e0�� �����ov��_ ��{g�|Ʃ�բ����;�NT�x�{ odxۤʴ�4�'m�cl�:���>�"�� �w\0Ȝe�Yl��� M��nE��ޗ�`Se��(t�T����k 7�<��c�:���>��<���s���'}`�cċL���7%tv;�$�N�3�7l�&����/%�Wc��t�ʻ�i���O<�l���ŀ�%�	�(|�i�n�ܓ���f��YD���i�B�щR2�*�H���Mk>�ܒ}6<���x˻UE�&��Е��>�� 7�<<�v'� ����>��H�J�]+����0{#�>���6^�\]ٞ0o�U�XS�:�E�m�Wu� �/ �����$��O߾�����Df;��e;ũ��m�d�;`խ�X1����e�L��W$SwCt:n�6���=x�� ����&V���VU���h7x{{ odxzG�l��G��?P��VZ����k &�� �mIxAG���d- ��}s�f�{�(�� �]�v�x{jK�:���;�ذ{#��Q�J��M6��:���;�ذ{#�;�/+ �	��ҧM��L�K�eq�de����4zvb�q��ɢ��[<���j�h����[�bM��Is� 7�<�����x양F1�EۻM[Xٱ��H���+ �}��7ob�%waWe`�.�6���yX��x{�\JK�X��x��V���ڵn�l��`�%��ذ�c���V�B 1V��^n`H�v�YI���@���ذ�c�;��,Wd��lU��)���h� �:Xj�b�\����:ה8xY7U��vpe���-ٔ���߾�w��^��/ܪ���;�<���ܼ��X��w�����^��ŀ� >�l:��-4؝��w�"�7��a��y����`.�TE4�%Jݻ�X�r��G<�w�xd���w�"�;�C�c)S�EۻM[X���ȦV�܋ ��[�b�<�Y��+�p�D�3VY�WV�>�՗�&���*����ۮ,�4�UN�!��ec�S��k۲�89��1e �5X�:�J�i�If���g�B�d|l[pPV�|&�=��{m�y�֖�^��!�<�<�zpָ{��ˠ�@��@1p��q�y%�핪uB#�Iˬ���J����`�;�K�^��Nڌ�)C�!L��ɾL��H�a8h��)���d5-s����`q�����Ze������T`J�e�s�4�]Yw��z}����%Ȱ��y���vjع+�*��t��^~�H�����v�{�'�VRb�@n��r, �������5vK�7�r�L��*�ʶ�X�s��[��nڞ�Wd���ŀwe��:`�m���T��5vK�>�ذ�c�=U�y$����mu�m\�mHa�*�A����\v9b���2-J�.m��6E1�����x�� ;6?r�����o����uIU�S��B�����$p��p�9��$�� ��2L�~���� �܋ �uT� ة�.��wl�͏ �ٌ�5vK�&�:l)r�;c��]����[����5o�x��X���	!2�m�����[l�:�%���`{#�;����?}��w%嚊���sF�+v�j�-л�B��&�}.�<O6e��̡R^q����.����`{#�;ۑ���/ �H���m�*�m`{#�;��,����� �vP����:-�o �d�������|t��y�?o�52�me�f`�Ȱ	5� ;6<�e�`-ڨ�t�������&� vlxd��{r, �kn��Q|.��.�9j-AVV��� R��(i�띮�A��e���K#e6_����ـ��Ɍ�7�"�7u� �6�x���"�m�R\y��8�6��{�~0�c�=��ҵfA�������{tH�� �$� �#���7��v� ݎ���Ԏ��Ó�)��۠~���
shٕ��S�� �UUm{���5o�x�Ȱ���K5�VVZ�;2���9mb��be��˥q:�M�e��v9�v����n�xjG��^�r, �dx�v
�t$�V[�mـuvK�RG��� 7}�v� ���R�t�۱�mȰ����.^�܋ �$(���	:j�V� w�<�K� �nE�Ir,t�R��m4�]���I�܋ ݹ�y��ܓ�^
�`�"�X����s����V��b�����mqt������h�]�#�ޭٶ�B�됒Ziᑉ�!'����f`(��J����E�4.���H�U�(ưZe��9���:ݮu�-�Ȟ�� ���<��j@x�Y�1��F�h��޹��O76ʘ����}Of{��h�1Nҍ��p���1� g%�Tb��0lA����D�nx�����t2���X����fu^g7l�b���<�Ձ%�a�	eIta���nD���8���ݮi6զ�@�o�XeȰ�����,B9e�T��6��m`.E�� ���|���M�r��Yl�j�V� 7v<�� }$x�� ݒ�W�� wV��vD�I�8`�ǀ|��Rn��]�um�M����G �����z>�����MB�͵�裎��"�!��==j��n-�X����j�BM6��� 7v<�K���r�<�{��<��δ���ֵ����$��~��>@J 0�FW9������g� ;$xv�X��.^;���w��xV� }$xeȰwc�6Be]&���ت�h���^ݹ n�xknE�HG,���hm]���Ȱwc�;�8`�G�{��tx.��MZ��cIm�	��ViGL��I��N��հ��c�i�Y�9����Uo�{��@��8`)%�nE�n�B�cJ�uwV軶��G�W+�}�<���o�߾|�99����� ��a�̥�p�{׀M���_QS���ES�PV�Ot��+�a��l��`2L�8>1�Bh��P��t��Pخ�gb��`ŉ�-#"M�z�d#E&��!��3�ŉ�!��`ŋ� ��g|uf���En�.�ox���� Y����j��V�ܬ�$oU���e#�'��&k��M��$�O� ��\ s�N*���T�� ���Uj�AR'�*. l�9ꪪ�6lxkob�>]ڨ�t��c�6�ۑ`�c�:���=�'!���w������	V�@Z�2yhov<�K� �M��Ir,��ʽgi,�Ft��!-����i�MgK�@�ݠ�����"���7
 �:��W�~x�Ixˑ`�ǀl�ɥn�ڸ��\ހ|��������ǀwc���'I�j���U�o �r, ����� �H���P霵|wE��m`�ǀwc���#���*R��2��ٞX�JcT;���]�o �lp�6�U{�_�l�y`{���4��
������Ͳ�fLtz����|mG�pW���q1�J�Q�q�S�Yjґ�ٔY�� >���z��|`�ǀv��xݽ��S��-�$�6��p�ݏ �6G�I�b8�n� N�ۻf n�xQ�< �H��p�>r�:Ul�W��xQ�< �H��Ȱwc�6Be]&��t�v��0�#�?s���_ I<��8`�*�L�s�Uڪ�zt�wK�_�ƴ���=R��շ��3�4��6Q��|m+� 7c^֚v�Z�\��Qu ��k�ldgr���d:ژ�s�{3����q�z�@�'�.8m�aǈ�;XwW]�_��qFꁔ¶�F"Ф�v�Tj�9m�mn�X�D0�̩�]��6���;'/78�hn9�]6�݇�L7r#¹C�[\��mKfpV+��#�d���k+6�jݞ���scvmb�ܺ����3�3�d蒈�5�p�ŭ�7�=��, ����� �lx��C�I����m`�c�;�Ȱ���"�7�P�6Yun�wm��R^ vH�ˑ`� �I)&Њt��Hn�n��c�;#� odxvԗ�n�K(���|iZm��� �\R{��5E�< ����c�ݲ]V���� �s����f�mmД���mvL�ڧ���(<v���|�n����Z�x�����9\��{��,��.^'eҧt_m��.^M�U�k��ۑ`�Ǟ�������Ӷ�Wv�v� o�ߞ�{ n�x�'�$�2˫wi�����{ n�x�w���o��C�RC-��V����ǀ{�=2�� ��E�/ ��{��]7G]-�k�WGo�%v�h6 ���������tA�#.��-��jez�Z����� ��/s�\��	'��}�J�J�"���� �H��\�RG�s� $�x�[/=UIc�z�-�[��զ��_��wc�j���Q��A� ��+��e�srI�����qP��T��i���ݏ ڑ� 7�<R�~��;輩r�v$���7K�`����?~}z�~Xٱ���o�W����+iիvһtuIㄈ��`y8ݺ�u�٨R�X-���G'�;��{5l�6ڨ������=��Xٱ����W�=����O��ڢ�\�^���޽�99$�$䓛�{��?~����z�\��D��t�H���1;�x���%�/W*�$����z��),C�CMU�շ��<׽x'������r���s�}��씕�]�Cv�w��<)%�d� �jK�?r���9�z?A5sP�mR����i���=v��?b���l����6���N���_N��P��@��~�x�#�6Z��vG���Tڤ�˺I����~�$O_�׀{� �d��l)r�wJ�j��m�dw odxz���/)�^ o��6*�Tҡ��]۶� ���	��`fǁ�Jze�`�$��i��;�i��o �v^����s��>����~��'�}��$�,��!$��99rrI�͞٨e�c���]Fv��sT�͚A�t6c>�Q0����ù�NȖ�q�;q�@A�2�mȽpYÔy�˭/:.��u딶K��OI�3-\VE���l����&��F����[�<v�a��(ۯ���e�����AV��6���]�#�n%^� �Cuӽ[��lO�A�f!�:N5�*�β3� T��҅��v��z��O�A;�;t#9�pqZ��k(��ѐ�ٺ#������j.�ZU�Xe[���N��@7��l���{#������ �{Ԗ&���U��o �ke窩 ��<��׀�{����_����*م\���߿w���M������RF��x����7u�%���wcV���U�UU_�����	�ߞݍE���r���y��y*�X�J�CI�����+g�y|7�x��X��T��LtU�.�֦�e���!h�9�c�X	i�B� �m���v�m.Y��Rv�_m�g���� ���W����;�=�hcJ�V軻z��ܒ{��k~#,b�|AM+�3�޼ �O<�Z�=ʤ����N��Wv��6��5o�xٱ�����W��~� ��~x�NP�Uv�ՠ��xJo��KS׀���)�y����z�P�4[C�m�Z��-���{�x�����I$��j���
J�&0��vU5!�	�9�ձ��$v�Z#�+�/`y�5��k�_@}<��$�ɌĒK����]�柭bI.�e��SC݌mZm��I-ٌ�ܯ��6�S߿?�I/�i���$�vG���9�����BxѸ���� ���亮�uu�]�1~ �T�	"��)�A�DE
�U�~U<�/}�\��s����m��g��=qZn_}�Nrsw�;� �������xd�m�}޾����Ɋ�u˜�g ��}���9ʸ���Il�|�SZr�$��l+�f�	���l&q]ʷ����nU�n6m��4;Y6q��rH��xˈ�͵w�ޤ��<�I.��JkS,�r��������ecxj�f�)�	.��UUwkѯe��Il���$��q<��߾���n�MV��ߚ�Y�$�vG���~����c1$������������ۭcW"���~��y�m�}��n�m�߾�9mʉ�
Z>`W�
)˩���v�|����B0�1ڴ���[��$�r����{�纒_���kI.�>I(�T�CaW��8ղ�Y8j�:�F����x���P;&�A���%b�wy�	�	��k(�� �{��Jm�ĒK�#�w��%�'���^��{��m�}���~���3-���뜶߮}ۛ��|���tQv��|�a"�vJg;�� ��z��Ij���/߫��SmO{�����_���>|����[LFU9��m��$���+ĒJ{ߟ�$��S*�%���W�q������I~���eU�1:�-6�I.����%�����_�WԒK}�����&U�ݻ��K���> �n#���H�"$b�r������	f�O>h�R��IIQ�ya���i% ��_�I.�-!J���-dȚ	�B�[+CZ�%j(�e���� H�!�&���[l!2� L"ȁ�Rh�a�b#,`0��d�"db��"� ��F�#jB�sL�H���S��!�1�0% V���H�RRV����$$�0HklP�Y$�!!R�1ddY�����c�	<	 B��)xT�"AȲF�32�ƄX0�D @�����7F"I�B!0 0HCj/���=�N ST���XB BFZ��^B�Є�a rr=����ݑtR�
�|�hA��m�IbRb�ZR!,��,�����)	`Ql��)�Hg�4E�� F �y0�	I"�� �FFH��02���i0`,��2)F	}HE]ǚ@�jԈ,6B�m7������##�R�]@$�Dc�QHI�|�<��b�v؂3�X�Q��a5�dS<��K�&�q�۟g:�ݥ�j����|�5Lw����ۍ��@Os��1-�!�mD>� �4(��
����;(J��AC�\Za��h�1u�L��&�G�k���vE��z��r���-@V;k�T69��t�o=8�&ݶZ��j�#~}!�o��WK�ڳk�Ҭ� BM�՘{�b�#J����lK֡��Z"�ZtUզs*��Ӛ*Ue���vv���WiD�U��vA5�D���Zkh�IbR3���ƌ$m�W�s��n���k�)� �'�55�T��N%^PA��h�mF�n���L���g���͈��E�0�5(R�*�NZ��$�;3z�Hb`7j�P"`j��v��(���6�|��6��g�Ȯ���V��Np�Ɲ�C�����٠� 4 j�h�M�Wm*�	��p:`yi]�xۮ��-�U ��k$4��IV�vc,�=���O1�1Ps٠ὗ;[3D�F`@�*0�P�\�zs�6�)HXl1L���lxK�f�Me��� �7.��v�A���,�Łʶ�V����ͣ6ƁƵ�!lgWy�G2;Km�^UI��է�@%�yۇ��t�r���>�ٗ�UL�j��YC)�]�C�f@Be@�zЂ%�$eh��b����lS�,+�Ss؋�`�Mɵ��%���+J��G�\\@N��S7by�+�'�Y۩��i�b)cf�z�U��	���8����$\#<Ap�Ñ�gS��{R�U Ơx# 6������f�^l�N�:� �������z8�)�%�a�4�z(ᰝ����h��[���c�ь-�9x��0M����+OV��F�a�#�-`◶f�S����k[� YMV��UU��)Zر��E+*�Jg���A��Z�p�d���v�I�′\���J�Z�O\�j�%g0iE{ }W�~F�L��%[��h���$zN��+���a�(!�� =|J� +�G�0����kYn�NΧ˞�6��v���%Fi���ȟ_0;x2�SD�"y�Ӗ�!��;N/�I��G^��*�vv��X#�1r�s���9&9c�I��+iI���	F�W��|��v2f��9a��WF`�k�[/����ϰ��m����JM��A$����0qўj�l���ܺj�U5bz�^��%�1��u2�]���I'��䜞3�%�U�t�m�1.z2n�}�K��.�mW ��F�اF镧U�0:kc��+�~ �����Ivl|�Z�ʼI$�l|�IvTWJ���������>��\���)�I%=<��$�-�bI-���YM ۫\a_} ��?W� ���};96���� >��}� ���Bx�L.���$�ٱ��IM��x�Il��� �������y���6ܹ_}M��x�Il���$����I%�c����}�5)M3�9&���t�Vj���*L�Z�̶�pn��Xq�bܑ��Y��l�I$�l|�F���$�ٱ���`;�;�� �K�rX�i�.㵭s����~�����Q� �)⪪���Kvu��IwmL�ĒK�c��W6��g|�6L�T��l�� }��}�$�ڙW�$�se��Ijٕx�IM�K�;[7W*��߱��x o�}��$�lʼI{��U�����$�=^F4"�1�j�< ?�߾������x �͏�Jm��x�KovR��.�ݪ���nz�]�F�6u=u��uI{d��![�j�,��R7;��hlF�+����cԒJn���%6Ӆ��s����W[I/�����z�Y|k��Įk� }��Ͼ��NM�߰�� ����@/����NrI�߾�כ��m˕���s]�v�o�}����(DDw����� �}��@��g�gd2��Ի��Q� kZ�����-����3v�O�~���>�y�#��h��K�s(�H%S�W�@)��������?����� >����}u��خÍݽ��ύ
[�m䶳����5�[\�q_�L3�-Ѽ�eK���z ��_}�-�bI%;�����J)�ĒK�ޠ�v�h�e_} �����l�<��$���x�IN�}��ݢ{�ƈ�c��i� w��}����yɶ;��}����< ??�>,`�SM[3Z�9m���Mw]�零�w���[o��������W 4����>~��W~�}�_�!#|�R�$+��o.�߽��s����"��9���m�����s����k��~�O�tM�흍Y�����uKO��stP�f�B��Ĵ�R����EY��sͼ��WM6ܹ_��߫�� )��$��̳�U_]������6z����nk� }��Ͼ�I�>��Y�$�����${�wi{�Fz�� �'.W�@>��� ~��Ӽ�^������u���3�-Ѽ�c�[Ef����� w��x ~�����y7��ﾁ�HGM�.ʿ�I% �X�K�W/�<�Ԓ$~$�>����Ns�}g�ox�m��EG\�tV.������aۛP�a�0p�s�I62�4��D�J\t��LN��IcJP��mR��֎z���KWc)���r)�u�����hk��&kbL�yNG�[�ѓc�T5e�뤜u����3�.˜O�(�jn�o=�'m�m���2�0Yص'8k�gû
M��\�I�M��mm�e2��t�սc#��f���|�9$��{��S-(gv6r��m����۷A�HG��97e�xmش�A��nux��.� �㯾�_���� }�c����ZI~�_��I/G���S��wcE���$����I%7c��SZ��$������ #.��Lt[k &�x�$x;#�;��`���;;�W��x�����o����X�q/I�wc�$�Z�0t1�6[x;#�?W��W��������t����=.ݶ�����5��m��{�s���v@�v	U�h�WV��N�Ϣ=��k�m��<�nǀ��ܜ祷����o�ӽ�H�6�6��O(v<9U]��W9V��� {}�n�ϻם�N�-���M��f�ʂ�������U%%�, ��x�Q�$>:e��M�{����x�<�nǁ��y�n_<�-�;��"�x��X7c���vG�~��b�:;%�j�d !r�(�SLB���l���M�J�6a����ێ�c�\�ۧE�� ��x��� N��_ �s� ݇�J��V���t�� ٲ�~�Wa�~�����`ݏ<����Uit�wM[���y����$e�&��ss�s�ܒy߻�ܓ�~��|j���k�m�z��g� ��x��<r���� �]J��]�T�ąv� ����S|�� ��� ����}��놄1��3[T���Q��Zu*oe�Y�ے�r�rsB-p$v��N��أ�	��{���y���R�hT�2��M��=�H��y`����G�H���SMRT�۴6��~��	� l�� N���M��tն�P���'� I�[�	��/�\�r��窹����O++Z������vKx;#�7�e`ݏ �ʭҟ�N��U�UL]��D��tx$m���-�v{j��7��P\�'�'l���T�e��v�������2�n��U|��޷�zy'�e'I[Uj���x�L��9\�A�<�O/< ����s�W+�Wg����wL੾+�I�X����v(��r��ďo��	<�`�)+MQ­�t7m�s���)s���y��"�	�;*R�Ĩ�鎕�o 'dx�U�T��_ zO< �}��$�9�����wҙ�Ս����������a�8S�S�FCU�s�MkB*�ؕ�v
0��7B:@�vR��<n7X�i�ɦ$��{c'�&��6�mګ0	s�%�iS�lܙ:N��ΰ���.���Q9�����Sq#�L� ��AE��{$�2&�k�r
� 4�����0�Ȯ9�3�j�f�f�F4��x���@�-��v'�6��X56�߹�ս�
��������
 @#�v��%�1��U��[l�U��ၯ㻻�?Y��暢�;m4ۀo���� vH����|���ui�*=���� �X��窹\H7��x�{� �u�?�7k�
VV:�MU��'m��޷�I���)���	'��u�HcNĭ�c��m<r��w���&�� 7v<��+�*�W{�ߓ�?~����Hum���V&� ����UR�y���� �}�n�����]9�t��[��C4�t�3ڡ��7m���[���b�*������ }�� �I/ܮUs�_��Oz�V� �����Zܒy���m��P
���H*(d"��*A�������F��E0$��	0Y&P�;�P�8��A>Ex���N_����}�~�w$�����Ag���X�J�>'Lt��:��^�s��� +�;���������'<ɼ��I�T�&ݦ� ݹ n�x݄x�r��T�~�� է���1���l�ݏ �+�\�]����z��\0	�Z����T�N���ƻ��3��Śh�ے���4��u���9�$	��tΖm�W/������/��ove~���s��=�~x���Zj�unڵct���)%��X�������}y:O$�|��_X�F�t.n�	??� n�x]w�*��ª�9�2?	|��J�5��l"@���C�'�:Dt�*�A�)��x#���(�)J:Ц�M2sz�x(b��M"I�B����"��n�F1�����Ӥ���@���$t; �w�`�1��6Ln5��jь�o�	y Y� Ne(���S�TM+� S�P�.�S�+��#�/ҩ� 4�G�8!� 0 Cj"��9O�nA�{޼��R���];,M�r���y�vxx�Ix{{ n�B���-���m����s��{��۞X����I ̐�b�pѹ��.��mX�Vb���YFTɯ4D&n�Ƚ��y<��-x1�L���{׀}�ذwc�ʮ~��lCߞ��s�)����&ݦ� �nE�� n� N���H�Ǹ��1���l�I��Ǉ�W�r�����o�?��؄����WwLN���q)	��y�lp�}�+��U�{��hct��-X�;i�T�x���g��'�� n� �\�r�Sg~�Gu�V�P�5�[s�H�d�y�WD�>�W�kX��A�K7�L�b+�+w�6_�� 6lx��?r��zz��u�vʫ����	&� l��{�<T�xݽ�=\�A=�P��n�Rt7m� ���l�=UIwny`���'eJE�>��M�{�����;��, ٱ����f��Q�.�w@��������&���>�{�_��6^����s�=QV_��Ȱ�UR�������ʝ��nh�v!atbYՎ6�e����Ϋ�܏(�m�JQ�9��{�����{F��<�8Atf둅��ܮIN��kI$��2�*��kL\��&���t�5�Íu!a� ,[�jh�b�H\i�V]JB�U� auA��4�W���o]T�#���O7Ug��-����A0$����6�m5�B��I'I		�͌q��q��p$kaܜ�{(:��<��u�say�uN�P�������}�x,h�;d ���� 7uG�uM��w�� ��0�;i���m� ��<�9\�F�O^��� 6ly�r�\H����n����;n��� �����?s���]���� ?{���	��㪷i��7t���ۑ`͏ &����NK�����>�����i�\`���͏ �*���R�O?���׀}��`}<����;!3�lT�Q�9֬E�%��,��	���ȗA��ĕ�݇F�>�:�� oM� �ݗ�}�"�+��s����<���+ʵJ�@�N����߳t��T*�D�'�Ђ��E^y;���ܒy�ߵ�'���x��j�)�i�v���ŀwc�ܪ��U%��wny`�TT�:a��O-�vrNI6��sm��}�}�ф�9\���� ݞF�m;���4��5ulxݽ� �ob��y���}�;�63���m���R�<b�%�!��Nѓ�e�o(F�/�����>��&cv'c�v�w�۞X�r, ����ϐIjz�	���YIڶ����k �ob�����ۗ�}�س��)#�z�|����ՂI����os��7(��`|��D�ϼ���I��ެ ��B����'C�m��ۗ�w��`v8`z��w}�zz�ŎҠhC�;J����ŀ{�U�s�����w���>_~��a.�V͜[�X�S�]�T�rà(G��y1�vn���ŚxT�>&��X�m`v�, ��<{{r���>A�s� 7ު+�S��[���[X�dy��+�n_� ݹ�}ݙX�A�16�ҥwM[x����v�,=�r�����Xݞx��*�4ӥv����UW9K��ݞ�����r�+yV_Vǀlғ��;�i��6���ٕ�z���ݞ��}�ذ�[F:-�n��v���Gm����[h�9��;&�je�5!��
/d�6g���]]7v�vπ;�� �]�xݽ��>A�Oe`�(^i"�.��m�x�엞�ʻ6_�,~�� ��z�#���!�$�1�	��;�<��p����K�^�+aIS�[V��v������V wg���%�~�U˓=�`�ު+���]��]
���#�?W+��{�_�n���;/b�;���wQh�=��b���~+��m0�]�jDT35̍��R[�qd�i��[[�je!B�Gt��Ue\f'm!�8�΀H�l�N��*�5�; ���0�����;��k�5f3WfL�x��98r=q��p뮌�b�7��m����A����1��̃taɳA�Zۉ�Kp��qf�G�W /,m�B��Q�qtZ�V^p�]���.����L��DPh���ﳣ:s����˟Xm�R��@��˭��S5�Լ��[!'g!� �7�#Q��rG�-�1;j��]�V߀�-���>��Xdp�����\��iӥv�!ۢ���ob�W9č��, ��� �]�y�s��~�l�WZ��O-����vG�m.�w\0���m��ڻ��ܪ�R]���	�<� ��_M��D��9����$�ze��)3VZE�m�{{�v�,�����=��|[ಙ��h۶��̿����7�u,�uMIM�`=�j�#���6#�E�'LlV��/ߖ�� ����s��;a��~o ����������i�n��;�ዕʮo9U�v���0/r<���{{��*����,.��t;f wg��v7��U%ݹ�n���7�(Tb�&ںT����r�J\�o ����;�p��UR]��{ǟ�Ճ6e�dr����נ��fx���<Wdo �*RW�N�k��[=n+d܎ƺ��sS�g2gt����ᓨb�2���LW�[�$նb���� �v<.���ݗ�ouԫo����vv� �v<�)#�g��:����Y�H7ҭ_�*E�*�oZַ$���u��9}��܉'�A�����#�P����rI�|�	��#�C�'LlV������~�O��nǁ�������T�	�5V���Nݻ�;��~�]���I���v^��d��'t˶�e�k[{QRW@7Nv�ʺ1ͣ�(J��hB1�0\�L�+�r�y@e�WN���l��<���� �n��;��w�(Tb�&ںT����do?U~�]���׀z~� ������������fa6��z�v^������˳}�� �7�l������նb��Ns������>��ܓ���k[��`@D��k����wL⻦�]����nǀ~�r��W+�\����}W����8`����kV�1�LfW��`�)��r�s�P�K@�͗FQ�s\:e��^7fwgm��M�������s��+���y�z�H�"�t�b������r���Gw�� wg��o?r�\�H��J��V*-۷n� ����T���;�:�z��(YWM];�v� ��6�;�>]�x�R��<`}�XSI��*Wt�o �v7�|�e�v�, �v<�s���p���
I0��H![+5�p8�I<�� BU|�	儍f(�olt(pUٰ(0#�p�C�a
e% ����,�x�P5�!�@6�6�n��@0��s�3y��j]Wa�̆�5�Ske�pl%�,�[Ec��������Ui	BwEa݂�1!z��i������Fn۲Ԑ�IeR�YH�Z�f�PDU�&�ykrc
�˴�(˵���v�����8�n�L��q<g`d�\��E�vۇ"9�V�],t�۶%"�h@1F<V�&�=��J�Q+�WZLh��pA��U�ꊃ
����ّP�X�n�*`��X��q̴�i�]0ei��Q�,e5���9P�7+J�K[mp���NL���l]hrt�yy� ����\�Ь`�I��X�� Pv{.����RTN�@JN7D�p�ѽ�3gv�\��nx3ƮC�v�<��ڤ��E�.f{on�`�k���t��b�hB�����4���c:��-i�T`�0�]�x�)�YK�	�`�3N��Ar��8�����e�+�C��n��OZ6�����L��P��i��[p�(jh��
iM�+���6�|
<@3$�qҀOƽq��R{;�,9�ўx4�M�F6����:-c�`�\��m+r:4�jPX�L���fQ�u���.&�gr�9u�'Um8�)�cu��fjqP�8.�-�v)��`
�-m���m-!έub]�C<sG\K91-�؅\�N�WT�e�mq�T�U�W1en^$-�Uu��+#���0)�z	4�F�R��-��v��j�2�j�]�Ȇ�p��n�P�`�By�ҫ��L�l{[�n*�)ʎ��(�j�r�TWm@)�"�T2Fȣ��X�VS�ѫR��6%i;VV�[���ct�e���pl�k���"ku6����÷�P��\)��a޶q7\�d:�s����Q���u9v�T�#��è{:ˡRr�"BM
Fؘ��tCɔB��v���;P�\�Y�=�@h\B,ѝs�2�uW[�9��I-b��*�)�cU��6¼t��'��(�Iv�(ۇ��$�p�l)�#�`:	25�8����$d�^�$�>ɸSϒ(�Q}�D<�z� i`@V�����<D$��{57�Ř�����-Af��;f8��m4��8�����%���Q�Aۗ`�\#ec��"T�A�'-4�P�v�it�Z��84���Ԛ��&��`^��u������=�z]��P�Bs��M�<+����5��ノ�\m��ܗ݄�(��YAp.�=m����1ۥ�]&�j�'���l�-��\¡X/e�E���:t�����Nxmr&nL'e7&�Ͳ�px�m�t\�]k�q4k�,E3?�ƾ���mUx��^�ob��c��s�����=��߿���C�ubn��{ }�v7�|�e�ꪮW�$�Ԭ�R���]��ـ�~x��� �n��>�p�ͫV�T��Ɓ�m�n������ ����R��:E��M�ۼ�$��� ���	���6',j麺v�ci7Ez�f�8�x��?��c&�k�ӷuRZ ̍mAM5MP�wn�v��w�� n�x������Uϐu{޼ �@����w�`��#���U\��]�w�uI/ ��� �d
U�7v�tU���o �{��%�v8`fǀN��ܹ�cm����������נ�;r;�>�)8��Ӱ��ue�x�{ vlx��� ��/ ��l��xL�4:�-��m�s�x�6��=�z��㔕dj��\�^]��7��6�w�j���g�� ������cJ��&܎���)"-�� �����*qe'H���i�[o ��/ �c���ʬ�W�8����m�$��R��M6� �c� vlx[#x��x�� �Uӻ)X;f vlx[��{&V�c�6�ңiR�M�eZ�ӄ���nd�-�܉l|��wZ�s���H��EX�%�c�Vm6W�z�������Xݹ�����=�~�E6�Zt�l���7�eg�RGv����E��>���&���;���`v�Xٱ�n���Xw]J���X�;,�Xٱ�we��2�>��|�iК.6�+�C�ݤ#�Ц��$R�"&�~�A���w��rI�ߌ�g�Z|Li[xۑ`�2�	�� ;7�@�����v�V�:�ZL�<�l!l8.y�gb�^��B���Դ�6�f��{;�v0(|t�lV��&��X���6�X�{�0��Wv�n�	��=T�o���~��7�e`�@ʺv���0�c�&�Ň����{+ ����;��cT�%m*���m�n��7�e`�"��W+�o���#�[,n�e��ۼ{&V;{ vlx]�x�'9ˮr�TWNR�4L�ʷm;Q�C�t���ӬD5"�WN�3SQ�%
��R-��a�e�"�౲���f��<f1�����M[sM��hv i 7�q��7��u��lc�VfT�������z�3΃�`�N)K��Dǰ�θ�s�7�6�hٖm;�{��.�H�	n� ���@�pt:yYyl�'.�i'�cqQa[��rrI��t��Q�`X�H�mAYe��e��3E0�E%Fg��p#�噅ؕ�
���6V}���� ;6<.��_���s���e`?:�We2�n��M� �������X��Y�������J��h�T��>&4���^��+����;6<�[�E�Q|�v+L=�qod��	<�`fǀE�^��bT��Uv�6��68`��O?�����2�z~�<�m4� �L\U�ܦkICMf�B���c7�4r����ݧqӵ<�;f vlxۑ`�2�U�O?���i+iU���o �r,\�s�ȁ��_��'�k�7$��~ٹ$���{�rrKO�ǟ�b��[*���M�����Xٱ��2�	�x�Ҏ����`z��]���`�y��2��Xݎ�_,e�j��	]� ;6<wfV��+ �G��W��6�Q���ּ�o�hn�[IlS,��6�Y���g��5�ru��[x�̬{&V�ٱ�d�/PŃ�:�Vt�}���NI�%�}�� 7�� ���W*�"�	0���X�i۬�����s�^�*�"�#1N��Q�5���ޓ+ $�EK)2��ժ� ;6<v�,{&V�K���n��J��v�i�Ҷ�6�,�9ɾ����?ٱ��%�L�ӲݧWv���Wd��j��.��H�KH];�gkX�嗏C	s5lY��eU����{��{��`f��W�=/�X�"��>[l�U�Wm��&� ���	�"�7�y<쓐/��gf�bd&.��7�m���M���+ �0�6��)T�&��4��W9T���	��V7�}7 ���`�E��}��ܓ�=%"� |t�m+k �ɕ�~�9��UU���ˠ��<v�X[%&0E]��1��GO0]��<��D�yY9������t�#�t,�-`-6�F��߿>0�c�'nE�|�o�����+�R�t6��]� �v^;r,vL�m�Y�$n����t����һ-��=�<�	�2�	��E�/ �5ʷi������i���������� �v^�qzL�M���v[N�V[uv۬v8`�9���~}~��`�2�$�H#
ϥ'�}�[��VI�� ��T�M6mU���5������Y"�IM<��ʃQ0Af�p�M�1�zn�	�닃+D9�C(�8��q3���Y���n��(
^�mn�l�M���ƖDv���w[�@�K�Lg���v�cj��9������AA\ԙ��鈁W�ͳp.���Ե�R4щŮ�\Db/^Nd�ȃc��ʕ��g�t|P�9�l�Rf�ֲ`�i��bQݫ���n�'jC��쪲�`b�Ktc��f�л'��y�f�`�2��p��ڻ��8�&ZV��{~����V7�� vlx�H��()�i���L�v8`fǀM�� յ!I6!���t���'d��͏ �r,Ԧ��V��TW�B��eZ�`fǀM�� �ɕ�Nɕ��ۨ�S���Z�k=�%�X1Pe�WK��e�ݷ&�k ��5�"����ZK�442��{.y`�2�	ݙXٱ�Mr��E+���V��}�Μ�9$�s��'+��U�Us���t��nV o��6�,�'%���Ŀ�f3e@c��΁���ݝ ����Uʤ��<�	��V��R�M[��]	�Xٱ�.�{&V��ʥݞ��kҮ����V���|����S}��;��Xٱ�߉>��Z5�����u�\��wAz�2�"A(���^k�c�Ir$���NH]st 4�av�z~���}ݙXٱ�s����:�z��{�%n�*t;'n���ٱ�.�{&V򒨨�4�*�]� ;6<�ݗ���U�!��r��R�-ϖ4��.��Q"{��"�@�!MMO��C�4��4;AC�P����F�i��xy�*��Q�>(&���[�p������H���1�0!5j5	G
l��y�,
D��`��<D�0�D4��E؀���{\�Ns������ܬ����
�wI�ݴU�+m�z�T�{=x�{+ ����4�*ݻ�`�R��V���+ �����ob�;6�!��Z�cF�鍐�.�����	lU���q��z��;IY7s���yf� ��2��c�>��X�L���R�2�����6� ;6<��ŀod��>�̬ �M�dEP�ګeZV��ob�7�e`wfV vlx�TG/ ��V��{&V�vea$��~����@���DX��k��c�LXWjB��I!:N�I۬�ٕ����ŀod��=U\�&�߾�{9����Y�f�Gl#K��\6`:f�(`L͋�eR�
&ˉ�[u��y�m�X�L��ٕ�w���i;MwJ�x�{��+ �ve`fǀM��&���հ���[�{&V����͏ �we�>���1[ff���΁�����c�:���=���� ݎ�J��+�i]]
۬ �dx{{ݓ+ ��~ٹ'��UNh�"��"0!ES `�$ "���)$B@ amH�R"�֢�!��.��5&d�5�]j�Q�������$ły���Ӄ�ٽ%�t[�sG�E�jz]�!.��v��&�] �Z���tr�u']���1m�s*������0<k=l����� ibbTr�/.�`m����+!�X㱡�v���mclOc�f�vz�%�3�9+�s¢��tm��������(朗���6UZ�(n;uS�56m)�4��wK�V,ҩ��n�K��cz5�Z��., �Sl6"��EX3�j��$�i6�ˑ`�2���+� 6{� ���9xQ@�鍫V�ݓ+ ��2��#�>��X���S����>�̬ ����v^ݓ+ �ITF	�wn�Zn��#�>�ذ�X�{�"IQ��t�4U�+m�-�xvL�� >�����}�����lŷXK�&�Hծn��;n���'���M:����+�j�S�aWwb�xvL�� ;�?s���ul����>+N����46�rNy��w�1�E��"���kϵ�����X{��*m"�մ����Xݑ�v�,�&V�ob���W�Qm*)����s���y`=��� ����Q��|t�իk �ɕ�}ݙXݑ�v�,��W�k4u��j���Pf������g�m͠#M����:�ښz ԍ$�୻������V wdxݽ� �ɕ�|��#�cvR@۬ ����{ݓ+ ��2��J�wN��t���}�ذ�X_0����ݙXٱ�u9J���M��]�ڶ��X�ٕ����*�u�,�����鴓wh�� ��� �*�Kg��v�ݓ+ �H�-��ݶ.M��L�wkF�	��̶�l.�6d�ʃ
���M˕�e�]�.�d�����>��ݓ+ ��/ �r�aI��m���wd��>�p�� ݕ��Lm]�0�X�ٕ��$l���~��$���cE	��.�`ۑ`͏ �܋s�ʪ?#�B+�����ܓ�߸cv��I��fǀ~�sc���OOe`ۑ`��\�*��^�l�������#;;tQ=�CS�<��6��.��� SV��ɥkʹ�_�~����f̬�r/ܮs����=�?R�n�an���w�lٕ�wnE�6<�d���ʫ�OR_u`�
�/�X��`|��x�fV��R��:�MZ+k 6lxV�x͙X�-��X��?	R��q���xV�x͙Xv�X�c�8�\���I���9�~z�3b�qc���h����U29cqa��]��ڳ�:ԅ�v���P�Ifۓ7d���I���\c;�nA�ɲ�����m;g%�ZsX�藖PJ�qdL�p�v�p�g.m<rm�q8ۡ�B�ǸQƖ�j]�&����bڌq��8ȃ�{p�(@{;BhJT����jD�5�ѐ�TF�>Cs���GK4a����k����l��2�*%b�[6��,�d�KIsnvj�p�gi1��6���Vݎ�c�;�"����"�:t�.�`��6<�r,f̬�5zp<�l������=<��Ȱ�2��p�;*A*1�]&쫻����9�~�.{?~X�{�Vݹ l��	�\��j��Iҥwbn��2��Ȱfǀ}����>{�}��b�5�.��T<�lX4��΋�ܠ���ҬUXG,^�Ɛ�:�uh���6_��fǀul��lٕ�n�J�P]ۺW`%m`͏%er�������Vݹ��I�*\n��2��xv�X͙X~��_��zy���*�Tp|t�1&��fVݎ�c�;�"���uN�)]�j��Xv�X�_�{������6l��?W+�ʥͩ^�;h�[�r�\GFi56�òJ�u�e�4d�^�tDr����rզ�$�L��o���ݹ�fVݹ�R	Q�R�M>]�'m�ۑg�H����6_��fǀN��_�ؓ�J��m`6lܓ�s���H/��Vr��9ʥSܧUŝ�<����;���V�c��U�۬s���9ű�� '��ݹ�fV��R��[wt+]� 6lx��_==��wc������L�`��tJh��n#eqh�ЄZ�d��,.Pɛ�.��+�YVj6%���Ȱ�2��p�W�	��I��"�(��i�6��2��W+�I<�`���;�"���uN��e�0�u�wc� l����Ke�� ����:�����|H.ـ6<�d�f̬��+��UC�p��BE�$d> {����rO6��*1�C�l�WI�xv�X͙Xv�X�c�:������tݴ]��ɐS���y�6��@��3X3S�6�,�lb9k��;M�;+�I��lٕ�wnE�6?W�6_�����h����V�n��ȰfǀwnE�lٕ�n�WuL-�M�f l���Ȱ�UIOOe`<�`���A@7��e��=\�U-��X��Vݎ�c�7eJE�"���LI��lٕ�wc� }�<�r,�_s*��h�@�����#E`��4��G`�P<$����N !���D٤�I����_)�����v+$!�4?L�!%e@��P��6�� @d]"�=8����	����d�:<(Ėf��3J�,f�l��7�l��O �^�
B$A�<_B"'.��	��	G�S	 ��C���k�<�l���㹈lS�Ϡ� �":�'�����B$"H"�����/��m�e2"�! ���*�;
���V�'��Ào`�@���!!F�ўl!#�C�r�d�O(9���5@�4�M*Y�-�A\X0m�,�k/	��k�n��5��T�(�AI7&�9.x���M�k��ѝHR�*�X�ݵuQ�1��8�(�%�햪�[@Q�Yy�+#,���6��(d8yӃ`���V�F6�ʊ�-\>�n��.wj7��]�ʇ9wI����*�my�7�k�¥2���t��a�s�R͹ݍ�fAC��!.\l��g����*�q��VKqO:5�.`c#�ķ+�Q!IZ��2[C����B�s�[6�J��i�� Cڮn��pk3.�(��ɱٞhê!6��2�l=m��x_\���Ͷb�\:����J�8L���rh�5�K�Mhmm!%XqhΚ���=Ѹ�{Xl����\�!3�1�=g�jzݤ8@��[��z�3�r�L���
�Vm5�7�F�F{k5�gvY&�ݶ�+����[D�ȴgʒ�;F�n�v���.Q .�\A�Np�1M"��$3n8�݁�B�+�lu��9Sq�v�M�����y�G1Z���Z�w3Ɲ�sV鳳n�6�q�o�
� m��j;5\�mόL���c"�NɝBi�&��A��sl&^G���Y��m[�vpky�]��,�/2�J-�1�
7P2���C`]��
����{-��y�͸�m��$ZqP3H�۶A������h��U+�g:��=/-,��(��:�NByΊαh�J7a���b�%)t����+'[pmGli%Fv���kmV�&��+#ϔ��M���سv�1���Ɓ��N��[G�������,�'a�n�M�:u;���C���`s
g�#�j��֣g0fܼ<\��Nض ¹��g�)�c
;h�u�n�
���!�LZ.�*�;�5M��-.��nDWi:��T.4�* �uU��9��8�}���)���X���s��*�[�S�-1�/vҕ=�5ʹ��Y�UIt]+ػI��u�&��z��"�xh��D�6	�P�> TC�<G��3�ڻ"�lf';j�]�y�����'���mAd��3r�ԭ�[0��A	X�5[�<�� Sq��m�� �<<<Y	/c��
p�����h2�H��S6������/�n�:�b�-�kU�č��k]#�٣�&V��⍠�vu�p����2-��K�z9!6�xݙPۃ.�Fy��+d�<�b!3�+kuR�<����'�B�ʰ�i�M9&�\^�x+�Z׫���v�'I=�93��.8�9۶��Z���ˋ2��-5���m���� >�<�r/s��W�$�����=e.+t�$ـIݹ��+ �܋ �ԂTc:Vʵbv��r,wfV��%���w�~0	�\��j���%E݉��7�2��Ȱ��`[%�kI��17i[.��n��ȰUUw�<|��^�ٕ已rI?~���z�m���*U���u�x�����F`�K��/��/``�`z��t[j�*������ղ^�ٓ������o�ߧ{;-İcar��d��|誻6�e`lp�>��nʔ�b\O��`��{�+ ���V�x����Tؕ;I�ڻu�wc���ղ^�d��ͪ%��ZvS�`�`�����{+ �� ���JU�t�ڦ��S��6H�i��-HUq�I�˺�ݳ���ZCIe�	�Z��ـwnE�Iݎ�`��WN�7C�J�f[�_�Ȗ%�by�w�iȖ%�b{�wٴ�Kı>���m9ı,O~�{v��bX�'���WR�Rfjhֵ���r%�bX����m9ı,O��}�ND���Hz+�:�<��Ny���9ı,O=�{v��bX�'�{��TJEH�7���JrS��@2'{�~�ND�,K�����Kı<�۴�Kı/�w��r%�bX��t��Cd�3.�6��bX�'�k��ND�,K�뽻ND�,K��{��"X�%���o�iȖ%�����wO�E���V�R������u�!�a	��H�ЛQ�ReК�׳�5��n�v��bX�'��{v��bX�'�w}�ND�,K��fӑ,K���w�iȖ%�b_=�;��Z��f�kY�֮ӑ,K����i�~c�2%����ӑ,K������9ı,O;���9ı,K�~	܅.k3X�&f�ӑ,K���ٴ�Kı=�]��r%��a�2'�����r%�bX�w��M�"X�%�ޟvZNjSVj���\�M�"X�%����nӑ,K���nӑ,K���w�iȖ%�� ��U1@�~D�|���'�����/'���;4p��j`�9ı,O;��v��bX�'�k��ND�,K�~�fӑ,K��>�w���B�������ҍ��J��U�6SL����gl8��Ƕ�S�CGi+%�D��k"z���צ�5����۴�Kı>���m9ı,K���bX�'�߻�ND�,K�{��V!�3`-��'Ò���'��}�ND�,K��{��"X�%��w��ӑ,K����fӑ?TȖ'��?��	3P˨f]jm9ı,K�����"X�%��w��ӑ,2&D�����ND�,K�w�ӑ,K���,�&�iѭ][�kiȖ%�by�����Kı=�۴�Kı>���m9İ?*�"g{�����oMzk�����4î�����Mı=�wٴ�Kı=���m9ı,K���bX�'��{�ND���5��/�C�u�6F���:��][��HW�M��q8��fm���2�e���,�/3��rX��l[�SJL6�iR��8���^�Rm��o�7��-��cE2�T�m<��3�K��#��\�b#
��ׂ`��a���)��S��{Jɒx ����M�
Sbm8��⍺�t���8�o׉.������eh�JDZ�L�2���t��zW�f��8R�::���p�l��{^Ӽ�Bq�ٺ�;[��
W�]v�Ř)�L�Oؖ%�bw��ٴ�Kı/�w��r%�bX�g��m9ı,O~��6��bX�'~;�l��Y��tY�����r%�bX�߻�m9ı,O3��6��bX�'�w}�ND�,K�~�fӑ?��2%�����0֮���eֳiȖ%�b{�~��ND�,K߻�ͧ"X�%��o�iȖ%�b{�w���Kı;߫�a���-�fպ�m9ı,O~��6��bX�'���ͧ"X�%��}��ӑ,K��=�siȖ%�b}��:SF�3Pљ$���ND�,K�~�fӑ,K��>�siȖ%�by�����Kı=����r%�bX�� �w���mn�]s��t�:).�dgex��PY�u絹�s��Y���؎���4�6[��%�bX�g~ͧ"X�%��{��ӑ,K����iȖ%�b{����r%�bX�}ӭ�Մ�N�j�]k[ND�,K���ͧ!�!�b$H
�P/Ϩ	�P�mx�ؖ'�띻ND�,K���ͧ"X�%�}���ӑ,K����ge.�md�M]f���ND�,Kߵ�ݧ"X�%��o�iȖ?��2%���kiȖ%�b{�~��ND�,K�߂w!u3V�M�\��r%�bX����6��bX�%���[ND�,K���ͧ"X�%����nӑ,K����9�5���9������Kı/�w��r%�bX�g��m9ı,O~�{v��bX�'���ͧ"X�%������3	7o.�v�E��.y��S��^Yp�#
�j�ِ�J���a�G4&4¾r{y
�%��{��ӑ,K���w�iȖ%�b{����r%�bX�߻�m9�B����Nw��[�X���'���bX����m9ı,O��}�ND�,K���ͧ"X�%��w��ӑ,�%9=�vG�c�V����D�,O��}�ND�,K���ͧ"X�:��b�_�s
	 "��)�D
�>��&�]��ND�,KϿo�iȖ%�bw߯NRh�2�e��˭M�"X�%����6��bX�'��{�ND�,K�뽻ND�,K�~�fӑ,K���o5��tkT���r%�bX�g��m9ı,O~�{v��bX�'���ͧ"X�%��w�ND�,K��w�-�s�t�M�:�%5����כּg�\b�c"HƎ*NN�Tֈ�8�7�:&)�'�,K���~�v��bX�'���ͧ"X�%��w�ND�,K���ͧ"X�%�|�Bw!u��5��.j�9ı,O}�}�NB�=���7�O/��m	�9��i7�,K���%���2��o���B����w�ND�,K���ͧ"X�%���nӑ,K��߷ٴ�Kı����a�EBcm��Oo!y�^O3��6��bX�'�뽻ND�,K�~�fӑ,K���Ļ��fӑ��/!y?���}�mW�P]�'���bX�{���9ı,O}�}�ND�,K�u�nӑ,K��=�si��rS���g���Ń���f�ƣŎwR@C�[S�[��+�)���n��b�u3T�kRKu���Kı=���m9ı,O}�ݻND�,K���ͧ"X�%���nӑ,K�ｽ9MY2�a�3P�]jm9ı,O3߻�ND�,K���ͧ"X�%����iȖ%�b{����r%�bX�}ӭ挴������m9ı,O3��6��bX�'���ݧ"X�%��o�iȖ%�by����r%�bX��_Y�K�i�Rf��WZͧ"X�%����iȖ%�b{����r%�bX��~�bX�'��{�ND�,K��Bw!�ѩ.�l�5v��bX�'���ͧ"X�%�|���iȖ%�by�����Kı<���m9ı,O{���[S�7=�y�6�6'�t�����6jTq�]�W%��y�n���Y�l���G�+PW@q��hakC%���em�����2���n4��CZu�MF�L��Z�7%��Fuż>_��a�܁�!_<�ɭ�L���6D֫Tp �O���'c���"	�qk/2%fs$L���l�!���M.�4v�Z�.nk�p6�R��=gFt��cI�+D0.ͺB六l-�kڶ��ղ�S#f����KWA�f�dپ�^B�,K�����"X�%��w��ӑ,K��߷ٰ�șı;�w�m9Κ�ק�o^M!�@
	맻�D�,O3��6��bX�'��}�ND�,K�~�fӑ,K��=����O�;�7B�ק����٫l�۝e='"X�%��߷�m9ı,O}�}�ND���"dO��]�"X�%��~������%9)������������ӑ,K��߷ٴ�Kı=�_v�9ı,O3�w6��bX�'��<����������g�%�]4ٱMjm9ı,O}�ݻND�,K�u��ٴ�%�bX���߮ӑ,K��߷ٴ�Kı=��gJfd�֮�JG),�.�,xV;5,�Am�ht���1��fc�f������'�����*y�����Kı<�]��r%�bX�}��6��bX�'�뽻ND�,K9>��v�ZI��E�r{y�^B'��}�NCb�(D=��
O�*�b{���ߓiȖ%�b{�����Kı<Ͼ�m9�2%�~��'�a���ə���Kı=�w�m9ı,Os��6��bX�'���ͧ"X�%���fӑ,K��~�_P�)�1������/!y��~��iȖ%�by�}��r%�bX�{��m9ı,O>�}�ND�,K��w٣WhA=t�zk�^���~�ͧ"X�%���fӑ,K���ٴ�Kı=�~�m9ı,O������#�H���-Mk�49nGh]p.�De��a�e������ֆ:�ϙ�7f�#��k8�D�,K߿o��r%�bX�}��6��bX�'���ݧ"X�%��{�siȖ%�b{��:kST2氹�K����Kı<���m9ı,O3��6��bX�'���ͧ"X�%��{�siȖ%�bw��Na�2]R�3P�ֵ6��bX�'�߻�ND�,K����ӑ,b}LJ@�H1$�)��ler|샥��0 M=$-]���FN8`d����ጋ��l��H� ÒBT���R��&8BJ��1��P���`Mv��zz>
l؇v'���*�>AD=�� �08���Q!���M��>�siȖ%�b}�w��'�����/'{�������Eͧ"X�%��}�siȖ%�b}����r%�bX�}��6��bX�'�߻�����������:K�`�r.m9ı,O��ݻND�,KϾ�fӑ,K��;�siȖ%�by�}��'�����/!?O��W�J��5Ŕ�H�[�JK2j�M�v�nc��AZ�F&CMd.L�,Դ��]�"X�%���o�iȖ%�b_;�u��Kı<Ͼ�l?	<��,K�k��ӑ,K���ߤ)�[&�sP��u��ND�,K�߻��!� �DȖ'���ͧ"X�%�ߵ��iȖ%�by����r%�^B�~���q�X�&��r{y�bX�g�w6��bX�'���ݧ"X�%���o�iȖ%�by�����K�����н�A,�`$��y���/���}۴�Kı<���m9ı,O3�w6��bX��$\H���@UB��K�}��r%���/'~m��x�Zc'���B%�by����r%�bX�g~�m9ı,O3߻�ND�,K�u�nӑ-�/!y�Ľ�c�M0���\JA���6�&�Ug�\n6+�m'�9�a&X�y�m��Ma��55�M�"X�%��w��ӑ,K��>����Kı>�_v�9ı,O>�}�ND�,K����N��G9wy>��%9>�{�w��~�L�bw�w��r%�bX����6��bX�%�w[ND�(�S"X��{?�nf���\��������������Kı<���m9����/�~���"X�%��w��iȖ%�b_��N�)r�!�i���ND�,KϾ�fӑ,K��;�siȖ%�by�}��r%�bX�{��v��bY�^N���[�`�59�r{y�D�<����r%�bX�g�w6��bX�'���ͧ"X�%���o�iȖ%�b{�xp�;����Ԗ�Kr��{Db�&1�C,��rgt�} R�h������#1���(M ��.n�W��n5�\ef�2��r���hQ�Sf���AΉ,,����`.۶˫��4)u��V�� ĥ*M�NGL��l��۳�r��˷k��u!4%�A.�;\���1��#"�+_$��(����d*�U"�^VѸ�E������w��1�sr��;k
��Rt��{x��]�m�]�w]nhQ:j�reZ�k�����Mzk��~���Kı>Ͼ�m9ı,O>�}�ND�,K���ͧ"X�%�ߏ�}�Km�&Aw���B����o�w6��bX�'�}�ͧ"X�%��w��ӑ,K��=����Kı>�vu��ؖhc'���B����߾�iȖ%�by�����Kı<�~�m9ı,O��ݻND�,KΟv|`�L�GEN�|9)�O��!&�~���r%�bX�����ND�,K�u�nӑ,K��߷ٴ�Kĳ����g��Gumr�9=���/!S����ӑ,K���}۴�Kı<���m9ı,O3�w6��bX�r�:vԱ��s��5��mՄK�U�K0:V���-8u����$:�3Oc=3�kڵ�]k6��bX�'���ݧ"X�%���o�iȖ%�by�����"(O"dK��;�ٴ�Kı/�~	�!nSYKL���r%�bX�}��6�����M��D�K��}ͧ"X�%��}�siȖ%�b{����r%�b��w�����q�Q����^B�<�����Kı<Ͼ�m9���"dO{���ND�,K���ӑ,ay������	7��y���*Y� dOu��ͧ"X�%��{��iȖ%�by����r%�bX�g��o���^B���O�}�����ND�,K߾�fӑ,K���ٴ�Kı<ϻ��r%�bX�g�w<��������������c,\SƧ�WCa�tYvIgsk5�;l�g;nye6�h��g5,f��맻�^��ק�����r%�bX�w]��r%�bX�g�w6��bX�'�}�ͧ"X�%��g{=eHU��[[�'�����/'�u�ݧ!�#�2%��w��iȖ%�bw����Kı<���m9��eL�bw����4Ki�,��f����Kı=���m9ı,O��}�ND��������E�C��y���M�"X�%������9ı,�������F�s����%9(�}��6��bX�'���ͧ"X�%��u�ݧ"X�%��{�siȖ%�b_��N�%�k!�l�5v��bX�'���ͧ"X�%��u�nӑ,K��=����Kı>�_v�9ı,g�:C�ݼ�\�%��l�qv� X�+�܃�ӣr�:��uCD�-�f�"�u�ѭd��N'�,K����~�ND�,K����ӑ,K���}۴�Kı<���m9ı,O:}��]SWSY2�r��ӑ,K��>����?
�"dK��]�"X�%��{��iȖ%�by�w�iȟ�ʙ��ӳ��7Wj��P]�'�����/'z��]�"X�%���o�iȖ%�by�w�iȖ%�by����r%�bX�߻��V�XF[�����M|�d/O��?M�"X�%���~�v��bX�'���ͧ"X�ߞ@���y�"kϷ��r%�bX����4M[�ٙ�L�L֦ӑ,K���nӑ,K��=����Kı>Ͼ�m9ı,O=���9=���/!y?����4e@X�wY�q�a����~~���9����������X�7Y^���,&,YJTf\��'��/!y
�����ND�,K����ӑ,K��߷ٴ�Kı<�۴�Kĳ��O����s�;��JrS������iȖ%�by߻�iȖ%�bw=����Kı>�~�m9ı,N��	�B]ML�R�.j�9ı,O;�xm9ı,N��m9�����=���9ı,O��]�"X�������7X�*�9=���,N��m9ı,O����9ı,N��w6��bX�dN����iȚ�צ�>y?z�9�+v�	맻ŉbX�w_v�9ı,?"G���ٴ�%�bX����6��bX�'s��6��bX�'��b�EI	'8rNBI�L��[�M�utS��뗑��9���R3��g��5)��-W@K)�Ύw9�f0�5ZGS�-����qs[q�y����|ĩ�6���
����c#�hBjqt{��L[R�vuv̏a$��+S��E$
�4�5��X9JbJp+\�[-NuG��stT��sCl��^����N��˞�=PYL3O1��'$��{;-�L+���-�ܜ�0vsk/[2v�����ڋ�D��V�S:��U��O�>ޚ�צ�?���fӑ,K���w�ӑ,K��{�����șı;�S��iȖ%�bo�xxѰ�yknS�Ow��5�O��xm9ı,N��m9ı,O���siȖ%�bw>����Kı��=�>0e���6gy>��%��{�ND�,K����m9ı,N��w6��bX�'���6��bX��}���g�ږ���r{y�^K���ֶ��bX�'}�ݻND�,K�{�ND�,K���ͧ"X�2���O��a�r��y>��X��_v�9ı,O=��6��bX�'s߻�ND�,K�k��6��bS���g���飡�1���l�89scq�o]���ihl�JF��&��ђ���l5-��ӑ,K��o�iȖ%�bw=����Kı;�}�fӑ,K��{�siȖ%�by�ݹ�'2]K�֦�W5���r%�bX��~�m9�Gp<QN�n%���{ͧ"X�%��}�siȖ%�b{߷ٴ�O�eL�5����א�Ib�hE=t�zk�ı?~��ͧ"X�%�����ӑ,K���o�iȖ%�bw=�siȖ!y������s3�b��>r{y�bX�Ͼ�m9ı,O���6��bX�'s��6��bX������m9�Mzk�}��ƍ,��V�r��{�X�%��~�fӑ,K��{�siȖ%�bw���ӑ,K����iȖ%�b~Q�������Zk&�h�5��EΉH0YF�*r �lk��c�؄�mf�t�P�(0���)���NJrS�����iȖ%�bw��9��Kı;���q6	"y�{��A>���M�m�\��ݜ�9�߽��t���bX��_v�9ı,O>�xm9ı,N�w6��bX�'�jt�kRMe�ֲ�kiȖ%�bw�}۴�Kı<����KO�>���zz�g�<���fӑ,K���}�fӗ����/'w��z�ݣB�'��Ա,Kϻ�ND�,K��{�ND�,K�k��6��bX�&D�����Ow��5�O���o�j�1G+��ND�,K��{�ND�,K�������i�Kı?g{�6��bX�'��}�ND�,K��]�Ԛ�I��ܱ�컰�Ǟz����Mv%�cp����m3��e�t���z����,K�k��6��bX�'sﻛND�,K�{�ͧ"X�%����ͧ"[�^B�w��w���+��r{y,K��}�siȖ%�by�wٴ�Kı;�����Kı;�}�ki��'I!���7��4K�m�.m9ı,O~���iȖ%�bw=�siȖ%�bw>���ӑ,K��}�siȖ%�by���jLɖ�h�$ֵ6��bX�'s��6��bX�'sﻭm9ı,N��w6��bX����W�ߑ5�y�6��bX�'�~?Xg,�Bi՚��ֳiȖ%�bw>���ӑ,K��}�siȖ%�by�����Kı;�����Kı�|>����(�2d�m��=��`�mb{hD��,U�f��э�R[�f��fӑ,K�����iȖ%�by�����Kı;������șı?~�k6��bX�'���C53WնK��ND�,K���ͧ"X�%�{�{��"X�%�����6��bX�'~�ݻND�,K�~�˄�X56fv��9=���/!y��_9=�,K��u�u�ND�,K�k�ݧ"X�%�|���ӑ,K��w�ӭ:i�I���Oo!y�^N����ؖ%�bw�}۴�Kı/����r%�bX�����r%�bX�w�y���1G+�'�����/'z���ND�,K��{��"X�%�{��[ND�,K��{�m9ı,O�|����1a� ��T4b>Of<%XT��tnm؊��]�>e�6��H�bP��
�	" ~c�Sd'"�1<ϒT��@@!#tJI$.�a�� ЂKI!	�s!�ЬB7ZS��.���m�x8��!A!R2 BF!P#R�,ʻ�L�a�J�@��#*�� �KBX��9�FA B$#!B���B2BFE�FEB!H ��8�]�l|,��ņ��|�"�q3$��$	!NB{���ζ]�%�ؙ&�7����mlpZ��ӝ�ٞNb!3����H� 7*�6&M�����]'a�Uz�2v�G���N���؇u�v�	��*�1�F�+t���ՍR��{.`�B�Wov-�J�ϊC���g����������ˣB!�(i��-r'm�4�ԱKT��*Ւ]�Cө��[Y���U+�"k�9����<�$ڂU�zM1�����T�2��[Z��ylm�bclc])�i	��8�`*ݶ��\F���6��ɓ���{-��Ҡq[vp�ץ�_�@$c/:%bu:����-�5�5��;�Ͷ����&(E]��.� A��Q$��&:9	`���M���a�M�%Q�tu���fs�; �І�2��pثa�٩w�q7δd���]l�r�m�P�$�бa�+/cXh�v
A�������*�檺���+�ɶ{FR6�%[)h��
���[)rS��M+Q% �����d�Q��6t@e�&�M$�a�FvB:�n϶"����y�ռ�خ��Q�T��Z���twm �\�n��	����ȓ㧢�)ބf�c�b�4P]��b�Lh
Y:��K7$[��("�*yeu�*D�W<m/-�6�S���q��̔�x/;�C�)%����Ƴ�m[�c�m1-�ok&��g���ɥ�n8�3]M�^'Z�t�5UNTAn���KM+�wX3S#ĕ�n��*�h��V"�TZ����Dz]��:���mm b]MJ��ٻKۮ��p[1՟6
�ے]�B����ܦ���͙.Bzc0<N�"���I�׎��8:n:[նV�k��;J*�;vq.���tɋ�;��f�pٌ-�aѽ7{)��f6f�������.L�U������+txu{�wU���:�f-��d�����s���N���ʱӫ;��L�0�)���N6uF��NM} ���*��K��i�����Gl�;c4�¦�vV�%��w��I��4� �v����']���z/�p��hN z<���8��ְT^�4��n�P��-ɰn1ĭت$]�:�L���r��Eԥ�bGo��>��Nƹ�,�j�,�a2;*35��C=BA�S�]��zs�ƣ����e�u�f�e*f0#i�61��\mx�<��bJ�f�)	���.IY��jG�U�����#'d���1�5����6��u�6�ud�k6t�ZK����H�fTj;
~��t�צ��El]E"i�v�J9C\��/:E��-��0W�j��M&���[��G���ı,K�{�[ND�,K���bX�'s��Z�r%�bX��۴��NJrS������6ԴbMj���Kı/~�u��Kı>��ͧ"X�%�ߵ�ݧ"X�%�|�{��"*dK��~��XR�՚��ֵ��Kı;���e�r%�bX��]��r%�bX�����r%�bX���u��Kı>ώ��3R)2��S5�]�"X�%�{��[ND�,K��{�ND�,K���bX�'{��WiȖ%�b{�_���d��Բ[nk[ND�,K���ͧ"X�%��9�����yı,O߿o��ӑ,KĽ�{��"X�%�����r�L�ƳRd�P�2��U�If3v�k�R�(�R���h��Q=t�zkŉb^���ӑ,K����uv��bX�%�{�m9ı,O3��6��g!y���w�+��D��2����*X�'~�����8��r
�d@T6�8j���ND�.���iȖ%�by����r%�bX���������Ct/Mz|���g-�Y��n���r%�bX�����ӑ,K��;��ӑ,KĽ���iȖ%�bw��u�ND�,K��s�V�#1���Z�ӑ,Kľw��ӑ,KĽ���iȖ%�bw��u�ND�,�ș����ӑ,K����㚓Y��2谶浴�Kı/}�u��Kı;�w�ͧ"X�%�{���ӑ,Kľw��ӑ,K��߶t�fj�h�-Hf�a���f6t
%шt�fL��.�"`�M��Y��#a�4E�����N%���}��r%�bX����m9ı,O3��6�y"X�%�����rtצ�5���<�i`��TZ+�t�Kı;����r�X�L�b{���6��bX�%�����r%�bX����ӑ?*.TȖ'���C�ְ�Y356��bX�'��߳iȖ%�b^���iȖ?��$Hu!��	o�@>xn'�5�����r%�bX�w��6��bX�'���0ÙK����WY5�ͧ"X�%�{��[ND�,K�w}��r%�bX��wٴ�Kı<ϻ��r%�bX����u���kEɘj浴�Kı;���ͧ"X�%�����߮�Ȗ%�b}��~ͧ"X�%�{�{��"X�%�߻�a��ծh����6cqj��(��i��A�-6��Ƚ-3u�M��J�ubg�W�)�r��G�/���z�I%˗��q4쳅�J����Ix�e`\��	.E�w�%cj�H��� I#�$�5�E$��$�vTFP:�0`�m�~�W���WrN����'/�}��*D`�
��SZ��}��<���R�5D���-�����|���H�{ϛ�	����1����ѕ��֠���a:�ձ�Fˇ�^�vI�b�ʝV�����6� BV� �l��H�	�ư	.E�}$V��-!�Wc��v� $�竕�H���X�~��>[%��0��[WN�]�V�68�%Ȱ�+��%�=��{�x�	�HwE���ulv��$��^ I#�$�5��qZwh墚h���$� �G�M��\� �9ʪ��W*�b{֦���3r��
��[��[2WX�I��W���\�K6�]9ѕ8۵��V����:�.\2��p�`�KE\D�5#�L�r�FP!	�6x-����u<�ó���f8;6�O	�["������-N�c�;���u$u.c6�lp)�� d>��IY�T3��q�FЍX0�#'b��x{9���%-�k�
aX�m���O];�����W&�����rE�ݹ�`6BDn�������޷��5Ѓ��Uf+S��;
�} ����&܎�	.E�|�K�7eJX�I�J�Cn��"������ ����<�W+�J�t�h��0����oN���o���ZH�	�ư�j��EYm��	[��^ I#�$�5���)z��^����-!����lM� I#�$�5�E$��$� �V*e��4lŎ�l����(r�����k��P��̳.X�T���F����7�E$��$� �G�}�L�MUݣ)329o@�����I�I�rqKw�����G�츭;�q��v �� }$x$�Uq/z��x����;�J�U�j�v���I%�� �Ix�����,�i4�SC�۶�	.Gx�%��G��y�߳��4��˜��K�1fw,�J�;U��<Q�u��+�܅�8*F�K��4#
.�lm��5I/ >�< �G�Ir;�	�U.�U��$%n��#��<H�X�%�l���SWB�J�� I#�$�5���ܮ|R�F �
B 2�A�' ���>��nǀN��v��T���$q�)%��#��%�{� ���MU��V��6;m`I/ >� l��\���"���Э�������
�Dj�dlK4G�D��f����K�Wm�f���(���{�@$��I�9UU_ ���x�OV0�Rc�V�J� �G��H��x�����G�nʔ���CIS��۶��F����l� 6H����,�Fq3�U��9�_o�����y��9ʣ�*��Y\����Gx��T�TRi�|Hk >� l���L�T��JD �ں�6�l��2k�XӋF�Kc�\LYY5�-�݆9����7Ks6G;����x������j�^;�
|v��7ae�5m�e`I/ �$� �G�|����l6M�m5g@��������H���z��e`��R�`7VZl7x$� $����X��!���ym����X�<u��<�ߤ� �ݙXRK�>RK�6�Q���BՔ�a �R&�-�m�2�vvn8�s),�(�怹볥�����52�Z�V�5�#5HR�5Ǜـ/mΜ�q��!�ӝ��6b�C�9m�]���@��+q���\�6�FywY �{��ɲȶ�f�����{	�%�vI��.�~����rZJdV^-��V�D�31pY���� զ�#Q)�����{9��3���I��Ǘ�5�u�t��0.1�7�7)��X@˵h���XSR(���Eac+^X��r���߲����|���H���R�V�|��uwn����|���H��fV�Tv��-�$%n���x$� �6e`I/ ٰ�ˬ�SV��i��	$x�+ �Ix�r,wf�S��Ҳ��fV����X$� u��>���B�����Ġ��nT��yH�eغ8;v�:wP6)�ɩ�:[rslM��E"`|��x����Mܬa�U�2�|Wn�I��wnE�r�U\���Us﫜�f�׀v��+ �r,i���HISubg�x�G�mn̬eȰ�Ȱ�R�S-R�c�۶��ٕ�l����RS���?�����fj՛ft����K�`���2�	�'*���WP�&��0;>*w.�O���n�3�p��m���Q�U�dv��M�Z7�|���@6H��ٕ�l�$�k�Yie�J�k 6H��fV��X�r,wf�2�]5V����6�f�{�}�������vtX���=q[���(%3�&T	0��$�0]JZB!�H��xe�%��T������
9D�H�$U��!�H/���6�����%a"��1�"$Ц��~Y2׏��HE��"$4���+�FR�U�@���	��_�C��Wc<��~A�2b�ZB���٭�"��6�*����i�NC�� �h�:Q�K��o"H ڠ���&0��6P}E��Ag$<��ZA���Q�,�Oh� �kE_�R���hS�v��1*j=6�@�Fz��ݪ� �lx:��=��I<�ߵ�'7je[,wv$�զ���%Ȱ��X$��9\��'���#�>+�`	��>�"�	$x����"�^4�`����7MU��N�v�聫4��ۣne4D��ea�h�\�\TЊ�R�o�3�m`�<kob�"�_��W+�^�� ���YH|�-:v����`I/ �I/ �^6͔�U�(t�M7I�X�������G�mv�X�j�ڤ��v�HJ��Se�d� ��X�����9��Z�tHCJ�B����P��|�nI�;�+���v]��n��G�mvL�V�xW�{t�w��*��&̲�lAX��9�V����.����`��5`f�9�QX\���WWm+.�;o ��X�������m�������ӾL$M0�p�<��r,�UUU$j�����x�ٕ�n�r�T�i՗n�	[X����#�6�L��r,t�Yn����Й����#�6�fVݹ�^�*R�X���t2�x����;�"�>RK�� ��r���*��W>���m�9M���l(bpl���h����B6b�:50ri�P��4�*��T�n&cLG*�&SMKK�W
	�1�1�V�b��XL��:���y��)��' ����طG �b�l%��^�N�p�*��OgwD�� ���1��[0e�<]�>���\�by����X����й-g�Jn��뇛� �.�lp]��QDZ����?�I'w<��ﲒ�u�)����rl̐uf���N�n�B�WK�h��`��8�j�F�qշk��M�V���?,�ݗ����2��j�ڤ��-�H��|����#���xv�Y�T���U�]e�T��i���y��Kxv�X��vLT�ʺV5b�N����ۑ`�ذ�G�}�S*����v�۷�n܋ �ݗ�� l��d˫e���j�RV���V�F����ǜ��Y�uw&4��F��A\Ռ)�����+w�E�/ ;�< ޒ<�d�dR��TYmۥl�M� wdy\�Uw��9\��M����:�K�:�e���,e��t��[o 7�� ��/ �ݗ��6�J��MZ��n��o ��/ ջ/ ;�< �� w�Z����`����v^ wdx�)��ul��{��r���]�Ik\R��
���tIXj@6�,�P�5������eAKB��P���n� ��<{��:�K�5n��'d�N���+�]$��6j�XV�x[���#�>ݩ�t���Cm6Z�`ۑ`n��x�Q�Ts�^�@C�!�(�+�^��>[� ��r�gZ���V� ���]ۏ ���M���wI�+l8�w�wc�=U�{/��;���>]�x�]JUj؛��&Qt��e�+LL��H�s(fzP�T�\&4YuJ�U1aTnW�~�o=���0�v^ }ݏ �d��V覊���v��r,�ݗ�� ov[���TT+TƩ�m`]�xݑ��e��r,풭Xv����i��� 7�G�wnE��W(��� ����y��7$�}�h�L���]%m��(���X��x����1ӧ|*�nݖ�Li�0�H�,�,��'�]2l��Y��g��yuhe�7i;i�wm�mȰ[�����m�/ �u9Wc(�Ch��V� ��x�qK�>ۑg�\䜖���?���;L��s����p���>ۑ`����R�;4�R`��m�m�w�ul��j���� �d��V�h��i���:�K�5we�wc��#�U�Wj�9�_�{y�Is�[���L���P���ٕ�^94�,��0r7:��FT�v͸ƥSc"�C�zM%�\м�T�Z�[fH�26��e�K���q�A+�XYU�A��8��狳/�}���Ҧ����kF .L�Y�t��N�A���u�ͪ����l��Du�!��kl46�D���Q��7�۷e��y��mJȚ݆�r�����gI?��t��$��t��᧵�
ե�R����� �NRf�2��Fq�D+qX�GSA��5E+Lj�!+w ����� 7�G�uM��w�U��2��t�ݦ�X����.<�l�V��&*�E�.�5I]	��j�����[��{#�>�*���ݵwm�Se��e��G�onGxdNYn�,N�N��x�� �����w�uM��~��yוk֛�0�������M�إn�`-���4q�3��Yp��sd�pr����������:���9U����OW��������_-��������K,/%��!HU*��(�K����T�"�<��_<��}́�ߢ�� �d��V�i*��i�w�uM��}�ذ{#�5ulxݪ�*c�J��m�X�����xT�x�J�WF]��B�v�m`�G�j������ذ���y�S;V�� 6�&�8$���r%ŷ�fxWogm7n�N���Ơ+�t[o �܎������X�����Ԍ��]�;l�����@ݽ� 6lx����6D�]�谤�h[�V� ٱ�|�r�s�G*��8r�yTs�����RK�'a0Y�t�;%n�fǀoon^�l��ݗ�n�%c���I��av�{ke����>[��fǀ{��W+|�?o���Qh:������ˋ�YSQ��a�E���Y�0��R"�d�2 <ɦ�M��E���>�ذ{#�5uH��UT"ڦ�B�xv�, ��� �/ ��V��CV�v�4��� ��`Se��p�>�8��SV��"���y~��ܓϽ��r^*��B)
�R�9���������ݚ�5���UU�uM��vk� odx{�5�z���;{k��a%jK�f]��A�\Sɷq��e��I��)8���Եn(�m�6�y���˞X�����w�uM��N�9C�Rc��*����=�s��F�����=x�{�(��
����av�x{{r������, ���	,�H-�$�;m7n�=�r�ߧ� �����ܼ ��E'|v��hJ��m�X����B{�^�I9}��ܓ�"���DW� "��`DV� *��U� �
���_�� ���U���
���_����U��
� DW� *��U� �
��@U�"�� *� *��1AY&SY��'b �wY�hP��3'� an�� �"
(  T*٪)@T�(�QE
��  � ���� J (�T� 44 �����@.�  
 5 u@�kl��  �DI@ $�@.�  �   (�@=y��Pӝ)JZe
Pl�P�,���� ��p��=�f 9��^���9�  ����4�)�d!���	� k����r�M��   =� @P( =�:���@�C���v��AU�S��E7n�WwuW�޷QOx�P��z�mp*��n� Wz�1�T�=��3���X��‽<�=!���ӹ�8�@ @(  ��Q��9ځ�	��r�T��zu�P��,�w�=+j�l�v�:w0�A\��ـ��L�t=⇢� ـ�C���݀p n 
   @ =��(����2�; �	=nn� �2 ��{�	0	==�{O{�9Wf�p��G#v�(� ��X���=s��� � =}h �  ���@t�k=��{�y�M���� ��)KL�,��6P&�N�RӀ ����J  N�J6R�� 
l��( w0 t�����P�e)N�� �@�PQK0� "~�Jm�IR �'�T�)��@  
��T���  ���MT��*Pd ѡ���T�iJT @D�6T���1 ѱ6��?������,�:���:��J��2W#�m�)E\?�**⨈*��**��(����
#�肢�S���O��h�?�m����LM$���$!�͡$JJ� S[��M	�g�s��h�٨\eB5%0aCl�g$i�!\H%�"`�p�c!$�VR$4�R��!r�²�B̙.C3DlhD��!k���f�>m��B%X��!t5�%dH�S&L��%bă6���$�6aWK#���0(B�8\��� A�
m%3M�0H����~�gC;Iw��2�4�\,}ӎ�#�Xu:��CȚ�^�Btn$@���:�C�d�П1���p�ĉ,"S�� P��dp#B W��#��T�'��0āRV�@�$d�XV�g��6nd�\%����S	p��"G"�%aB]Kt(��+�qt���`X��Hd)��5�Nj�X�71#0 F���C'K���~m��W��<���?qac�%���"�ϜM<�����x�Na/B�MƟG=k\�>}c$��a�~�$
}����~�$	!8�A�kwt���
0j��Č�y��sx�O��F���h"�hHI cf���h��d!��C>�!��M焥!b��i���IR�4�F�3�T#�"i	 Ȅ��\�C3�4M�2�$>WN�L	\��IL�.|��VF��XF$H�$ T��,�58Z� BM���O�JD�	*K�FF��� �x�[4��4��n.��M������l������;BR4#LIRS�1n�!\$4i�I`G�'��	?J|�p%0]�@�K9�����c�u�|�u�dd
���!A� �F��浓g�ߺ��I
�+��f�L���SF��č�l���!i�,L�H��&81���(B�l�0�*j!@�Ԑ���XZf�]��#�~S5���%�5�]�}�����k�@�3�p˪�oI9��|@���)O�Zi�J��Z���.B��8�$I#�R�8$
�.VZ��`$�I��4̦���bn-q%SL��׽�����B$CF�j7N�k{5�&�Ԋ`%k5��s\�N$��	FC�R3x�"B����� CVfR晚�ޱ����H��q,!�B�A.9tM�$LcI�:�@���}���!`Q��!R1"�k�d	Fl�!ll$�a���2�d>�q�Y4O�-%��
D�!�Y#R\4�� �U�P��B�b���B!B��$���#�HHp��c@�\!Lee	C%�\fY���%�/�.x���2V��6�S��ee	R6�H%0��%�/b��,������z�ZB%��r��w��l�
�������~\�Yp���	������$�������$`����#VX�~e�\����I!e����,*��i�k���'��W�O���/�Ɣ��x�`�8��M]��8�Y`BE����,�����F�W���YN	$�),���D�%���j�ٷ$�Sm��q��?ks�������#��I2�0��Jg����!4�M�$a$��cI	�	�B!&R�?h,�F����FK�r�&9(ZIs����	p.0�
l�vp�����*@�+
��áY�3��!z@��K�f�{�;X!���p���6I[!>q�P�6��]��[����}�_/�P����U����>㥣��͛7�RoX_�.B!	.�@#
���+
������M�.D%%��!8��.a� Il(L���4���36nJE�&i����W�<�Y�wq.%�K��٧D� @��RH��ą�$H�	L��S!L%�%�fka.����W���$$.2�R���d,N sx���9淏�۩�Ӝ?J���ټ6��B`H!�'Xuĸ��M>sRϯ۷�^nof��d��F1�� ��p4��@�c_��S%���+�P�12H�?�6		\�n��C3d�$0�ܝ*l�H�"@�ʚɘ���
�ˉ?b�2! HB� X��)&ɑ�	4�k,&x�d,%����XX$ �p&j��Q�7�JIx���C����ݬ�ݮxEB�&�n,���|�{�_�a�H�Q�O��G�	��I"����H�4`V pas�� �0�q��J�	CT�`D 1 �"E���$�$�
F��$a��i�LM$X¸�7�!,c0b��F6�M����A��4V�CS3r�R�	�!�SD�o�3{�e!�ܻӺa.4!K��u!�N�  �� @��$:�Oĩ$�@/Ĺ��C �Hߝ���O�
Y���%q�>�i��LcЕ#L��D�B���A"F� ���@! ��"�1��	p�D���w>?�FX��p��	Cy�|~a�E�~���$$��cM�af�N@4������P�|�D�+�l%!p��*Z@�S䥚LRq��7Ϛ<Cvِ��@����.��r%e5���ߢ\6��K	��Va�~9���g��ް�~��&��	-˘Z���@Ϸ��D)�.��kf�	4m�0erF��&81f�m�WJ��� S8~i��?aJ�$R�+	J"@�5�퉥!sFfB9��>��%��@��:c6Ԇ�b~T9�a�ԊY;H��L4K&$(F$���"���Y KY]�c
��		��B�.��]��U�u��Ja�����A�a$H,"H^kPNB%B$x� B�8�cYK��/N�Y4,`$%��[�@���~�>ڰ�F������(@$+ĀI���H��"Ƒ"9
Bb�adrO�.�B��
Y!P�+��rD�)��KKt)���L����B�� B�(�B$&?�D5���XI!y�������� ���Cϻh��4�.�zg�P�����ߎ3:c*B�v�(���)H�"@���aF!u!�B��0��:!��0��0�$�e%�p��V�e�9��2��������H�D�$	���XT�����a#� Y`Y�hK#�#Y!��q m	f'�y!ἐ��K!�x���C2��]!x��,��h7.�P�n�GA0�	�)�,��Ú{~�k��߄������!�h��Y�)�$����~��\ѡ�L�B7A3[o&N�8F�qԁ�" VY$S:����K-��D�Б�>K�n0e���-V2�{�τ��u�(D�$Ӆ��a��\�0�R�B�!j��i�,��0�ız����rM��l~x��c��
aB��+
J�rrm��@Ű'�%�Z��XI�ѻ��m��A�cR����&S�s����p��	n�r��>��':�$H:"0�bɽ��Y�Ai
##����kF���5�2@�u��"�"B��5�p�/�֐x� z�O���¥������%�	��Ře,���6��.�g��xݴ�p�sR�L���n���i!���dbԍX��Ӡ�����HNf�������)�4�K��T��Wa*���$�B⑷M2j&����*�v�,����\��q�&'��'�~&���B$d����bD���4��T��VR�._�1c���y��}9���z�+��rV$X�)�6Il`X�$־�>�9��3D���������7�7����C�`�ީ���g�_���%!HBV$.����	l��Ա�!#�B$"�%�c$$1+?2Je�\�iF�m�,a��a#Q��(`H�5J�.aP�Hȅ#D�*�@+�Ĉ@#�e�Ӛ�FB!�l�,jB6u�{�;y�?Y�0�������'�����<ItBJ�d
����dJ�
�H�$T&��<?l�5	
B��(F��(BE�`�H����@���>��޹�T��<��7�Lw$�X1
B��!�Iҡ+ � :��Y��?�qr�4z���	LF���l)��rY�h�l�#X4H`ЅHQ��B���X�t)qaĄ'����5I�bbF# �a��(@F�)&�C�כ�>a�af�Ed�%7)-@�4��He։7�	��m!Y"��h8�c@���Q�X0-�*��`$��I
P��$�4BnC�wB�S��=UU@dp �@ �@M����<     �Mln#H��p���� ݳn[j݀��
�	�������> ;�~8L/6ʯJ�J��� �U�+,�K�0pnһ  ��9���f�ں����C��US�mU*�m�pO+Ίq�Ͱ�cjVƕej�B��S@uUZCy���V���[@M�jx:]�j�
��l��;q��RZW���RR�L��MT9�*&۠)V�]��F�uJ��v�Y"����*�E^�R��&���:�M�V��v�=�����O��9�դZ��S��y7�`*����*�UUU[�� 6��N݅-Uu�UmI�dnU��B�5�k���UR�[*���AW� ��u6�j�V���@��\���AZ+�l/-!5�R���¥[V�[UuE֮e��+��ۤݠh���>��k��8&�Uq�gf۲��v���7S��4 ��V�UwR�����wc��9��T��dS��>��s\ʹlTY�c�8�݉�]�ݗ�����U�j�t�����ڀ]���#3>(B��Ұ��AT�dm�v��O;*�mUUUJ�X�@��1zP�6$Z�Z�k�x/AL��ʪ��ۋ!Oa�B4�K�^ �*��UUJ�ʵJ���u�=^��q��u�:F�$R��^32�HR��Һ�Z�Sz�� U w*���A�[��][�[j�v�ĵZ�:Z��걕Gel�Z��]��%j�%�yZ�����@�w<� ��U�����)Y�Z��݊�up��yt���ꪸ*
����i�����J����W��=�~�Om��iU�F�R���M6��w�y@�A� 
��6ø;�U�UUT�Ej�W�SrSkm��������(v�jh)�����v]W5TU��y�-���T�L���`�bͶ)T��W�W"�m�	eZ�e�Ҡ �UJ�V���[M[c���r�T��l;++VƦ
팇ki��%X6R�[m�W��VN+���Ij�Tb��p$� ���U!J�R��U����Z8�R�KV��U��
�����P6.$]�[m]H&خ@ڎ
^_���w}����z �p�6h���y��N�V�j��j���*pmeAj�j��h"UU��Gp]
�1U��*Ҫ��b��mB9����s+{m�eZ�.�+��*��vj�j�W*�Hj4�iV*�5-@e98 �U���tU���f���^ �]V��g@�Hɭu+�U*�K@��(n�J���w&���w�5�/"��v�M�T���_o�U�h���-uNRSjz�+��GZ �V�:4���eU]6�8��L�$X��A��ࠨX5��fV�Z�^]W=vX-�l�8ЗfwSҭ�8iYy��U�^�=Tm6������v�����ƥݥZ��QUU6�WvB�1m��)2�[V԰��BBbp�v�5b�QjyAy�j��d��UU � ���+�eh	]��ɚ�m��Yv�9JU�
ZmU+�j���eIJ���Uh��ֹ�UN2�0R�H\�T��*���^]����m;'?*ԫV�5xU�;�T���UcW&�W:t{2��kUTQ��5WW�^YV���Z�؍ ��mUT�̯8]�j�T�F�U��K]����R�t9@��[��y皺�ں����f@X��U����aB���O3���@C��������J����y`j�Z���8��n�лl5Um�O+)r�F3�R˳�[U<��U]/-P��m��Q�ʵumR��' �T�UUղ��@Ut��UTU,;�(y��Di�~]pw[;��+�'�U��F�YY�l]�w�ګ���UU 說���^6�� y�P=ڠ���UN�J!���ﾖ
'�����RV9��G30ҭj�j2r�UuN�P ���/s�N��    � �      {�N੷��+������J��@P$*�;iPy2n�4�wB�T�P��]e���BUde(�@j�Iۚ�j�B3��iꡖဠA��$�i���j�U�tR�ڀ�����.Z�v�XGq�9�X�n��wb�lx �m)�UYj�ڠ*�n�M�:*m+� Xw�3!�+�6�UUj�������@��ͤ+n�LU+y�ܱ�7�*�t��m�n=jVݕ��z]�tQHm�JM`��klV=ta9���g�=UU.��{AӵHq�җe�I�{v�&i���z�T�媀���+G���v�^8�&aR��f��h�@9ˬ]���ȉ�IDUU;�^wY4���
�@Ѡ-��yk,�aݮ1�U��dB�x����t�lЬ�@�����u�ps��AT�l*�M���&��\���˶��U*֬���z�jTlSP
���UK��*�p�����vZjM�UyX��t�S�b(մ�m%�p\����ƕ窩]�j�.�U��"�r��jnɹ
�Wt�ͮ ��y�komF��A[U���Z�t-&@ 6�Z��������Ue�R[���AUq�Tp6¬ 6�	vkl��  Y�3G��a	�ce�����S*�Tin6���[��8�UUVҲ�UmU[v
�ﾮ@gP*�jN��m���BqWl�����`*��p.�ْR�Z1�K&j�-����گ)@  �� xxV�+�U[UA�V�� {{�ݎ �  x �x6ʽ ��Ԭ� �m��\UQ�URs��yj�����mI�Tձ�Z�
�iWm�м�Tl��8
�]��m�TmO<�ꚫ`@�<5V��2 �SJ��ò���vT3�(+-���Ԅ  5UmP[e��Z0ʮ�*��%H4<ϟ}m�p[��>J�˰*�g��yj��m��KUR�˳[UU[UJ�z]���C�k��
�
�v�n����V�mU)���U�p��
�UmJ��e �{�z��<�6����x
�S�a�m�UR��Ut@�l���0)pUU[�We��<�@T��	P�Ř*�����d��\�ۘU���(�mؙZ|p/�Uu*�UUK̻c9,nX�+�m�p 7�x]�Wm�T���,@ j����pR��n�����1�P��Eۉ���@m+�]��@K	�� UU1� �
X%���+.�Yv�y[��.�v6���U[*5�J�,�uҭ[NIô�ڠUݷs7i���cc�(2WD�J��-�]N��)����h��Xq*�n]��o�n^����Ʒ=��v{5�T͇���ViUh)j�b�D6j]b�����X�i�:<	��.3fZicY$;�T�V�f��.�i^v�3�.pAQIe^W�k5W������V�T
�5Zt�gYKM6V�UPX�*�.Οl�Y�\\/[�u�3�+[r�Zє��Q���j7�v���Ʈ�A�9������v��i��n:��j9YU�������N��؀�V����[�un�4�*�UUUJܬ������ɷ��U�����6�Tu@UV�J�UPYV�% *���l��&��,��:���y	V���ڊ*��U�BN[�y[����1���UUUCݛ[j�>���������'�L�PNR���,dUj�v�8�?Uѹ������Ќ�v�0�`jB��5g�ƵѤ򳇞�s���$��Z�"vڪ���ZΈ�����D�VAs�,�	&�UYR��<�m][U�J�!.�d�F�TU-uA²�Tt���n�m;܀ ���;v7 b� ��;�t�i�T#serb�+���jW4�,
�UJ:�T�T�ӣ(�UU],KU*�u���ٺU���s��ܭ����unʥj���<��r�]�(� �Ll��W����
c*����UUi��{���]���r�     ʮ� C�wp�qs| *����SUU++UUUl��@��N)>�����u�uU�Ѻ��@
����;�P�5�T T����   ���j���*��v������66۪���� �  5[UmUA	4���@Tk�)nUtUmR��q��)@�eUV�ں+8��j�\�e��"j����VU�<\�`,�P[r���n3����x5lˌ@MZZ9V����Ӷ�b��ت��Ik�����Sm� <       Tm���Ų 6�]A��  ���������� *��P� w �P �7�[�� �;� �Ik�Z��jU�vj�%%ꪪU�j���^^|_W�[O .`<�m �pݯW� Q�V���O����w2�;<@UU(�Kv�n�YZ۔V�  *�Vژ� � m����R�V�T�v�pP �[UR�=GP������s'U��p%T��R&�j�کV��쫌U<�l����R�m*ԫR�K��UUUUUR�� �ëJ��N'pT�n���������]����   T         �
�  U   m���l�;�;���'����      y�V�`v�VW��m�yUUuӣ���Z��<5��vm2;m�\��;�t�;��:lT4�������"��R��"j"Ȃ:��_��6�S�(�P:A��`�nt5ôU>�tA*���0��]����8�@����O��H�8����:��8����UD�C:�D �?~9���D8s��p@�t>")�F�"�X2 �z�U?(%�*~��U�!Á��#��U(*u>�)��H�K��"}�
~L@U9�*����~����T�Q� ��A:(�H?�*�x	�pEQ�#���u�� ��>D���@�B#�T�Y4 ������o�� !��" .�$0X�b��Iê��D�tP�bX%�Qj5� |�NUx�~t+pz�Pv�Ղ��~��?	 sH��� ��0�|���TU��|���;`�U�����+P-R+�h�EH���'�����V���1UT5T��Umm&�۝Ԃ�J�v^7\�"��C��-TꦙwLܐ�3����p÷e�vU�V����+�np�q��&]ZE���ݤ�a�Ո�z����j��`�ii]�2����ٰm��l�ˑ�����:�gт�*�Zv�v�kX��Zϡ6�*: <�S٦^Z��jr�I��mQ	&�{��.�4�j3��cOVį *[�L��T�6Mȹ ��[X!�Lh�W�vi���Q(�x��v�Jm��Y��t7�\��U�vnP�A+s���)��\�m[�#�f�q�v�up����MV�u\�ʪ��#����`�\F[d���{qv���h�%5�2���QeQ���� ��fu�۷;�z�u.
�W�͛gjʛJ��@��YhUj 
��an���8C��JQ�c������X��鳃(Z�%)�d�7^��
�鱞�$��m��khE�i9�K���.ѳ�r`g�hz9���0'�ܚw3�TR�Kt0�\���W �X!����@H�n�R����&�t<]h@!�����!���r�l�qeu�R���"�q�`�,��$�#�{d)�v7Sj� �-���$��4��n�pUPR���HI�[(4Z\�u�D_8zEhK;�6��˗�1���G��LɷR×���8�c���	)�M��%!l�Rꆅ]N�v�d]q�9:�����5�+	j1�@��W4s��vna�s;�RcZB�v;��T��AEt˲�-@4m T��%����㍬g65�2�t 4�8�.�LY��8�J'c�5q��r; �YV��P�V�\�cPt2Q���X�UI�L+ Ф�(�vc1:Zk��cV�)���bf�l�UI;���\�F���J+(p�#q�p�&�����D�������n��L<M�%�6�j�K��r�Q9�r@ `RT��ST�sS8"��5��j�� ����O�~�hUA����~���N�^u$�����]��L�Ƀ�@-��v�	�h.��A�1�F��;%�CZS��ۧ-�&Mh�Q��k+5ͦ����j��+��[&��:U.���݃m@G����â^q�c���K���%2���mv&2���t������.U�q��7������NZ���%A�a���5dJM�[��V��q�VU�K�tUF����I�z�B7��]�nc�{�3�8L����{;q���e<y�"��p���L�v;�o@n	���	 �'���&��	�~���	�ı=���ND�Jt�O���R6Uu�5#q�Ëı;�]��r#�2%�}�f�q,K��{�m9ı,N��u�6t�Jt�Ow��p��\��%��"X�%�{�sI��%�bw�ͧ"X�%��>�&�X�%����nӇJt�JN�i}��u�J�[�秂X�%�߾�6��bX�'L��ț�bX�'k��ND�,K���q��N���{�-��$.G>t�t�,K��Mı,K���ݧ"X�%�~�sI��%�bw���ND�Jt�Oӻ���~i~��فs���nN.���.i�vݓP�Ґ������"�]#Zg�%Zt�t�Jt�O޿�v��bX����&�X�%�߾�6��bX�'{5�X��bX�%�;g�6դC&�|���N��I���p��b��\��h4$�U1T��4b-L]�㸜�b^�kiȖ%�b~�wz�7ı,N��{v��bX�'N�u����5s��)ҝ)����_:|ı,N�wz�7ı,N����9ı,�{�Mı,K��0Z�������ҝ)ҝ=�_Zt��bX�'~�{v��bX�s��&�X�%�{�{��"X�%���wf��5-�RXh�kV&�X�%�ߵ�ݧ"X�%����I��%�b^���iȖ%�bt�]Չ��%�byAG�|���\v��G�oX�!�m�4ҝQ�b��5�YY��JQ�#�9e�� �[�m�K�x��X�%��ﮓq,KĽ���ӑ,K�����q,K����Ο��N���4=�ظ�J�v��q,KĽ���ӑ,K����k"n%�bX��]��r%�bX?��k�å:S�:}����Ǝ�!unk[ND�,K��wWI��%�bw�w�iȖU8�
�U*$@��"T0��
�j2&A��v�7ı,Kϻ�m9N��I������3���.�^�X�%�ߵ�ݧ"X�%��>��n%�bX��w��r%�bX��k��M�S�:S����i��n����,K���v�7ı,K߻�m9ı,Nϵ�]&�X�%�ߵ�ݧ'Jt�Jt�i�dQb�c,�Z��%=���<�Q�p�m�kղnF�c17 l��l22��ק�Jt�Jt����Ο�,K��wWI��%�bw�w�iȖ%�`�ϻt��bX�'�;;�`�m��ܾt�t�Jt�OO��zxOș�����ӑ,K��;��Kı/~���r%�bX��wvjTq���L�zxt�Jt�O�}�t�KİgݺMı�0ș������bX�'�u�]&�X�%���g�F���c����ҝ)ғ����&�X�%�{���ӑ,K���]��n%�`~�RB@X=�?����v��bX���]�]e�7wn��	��\k �� N�x�(�k)�iSUcK:;�u�:�)��<=��c���9���G���l6�a�ۻ��4�o ٮ5�N܋ 'v?W9U_ ==�{h��E�h*�+��6�X;����\k �)RZ@��v��e�� N�x6G�l��&܋ �t�r�%v[*-�x�r��/Oy����mȰwc�;�	
��튑n�m���`nE�� M��U�U«�ײ~/��b�n�$���mP랸�Uy�\��#Bs�T�q�8��*�L��g�6� ����d굓G6����m�h䮁�
P�j��-�lwn������Y͞�u�mp�fF��&޹\� ����f�VNX^ܺvg����&;V�Y�̽\VzW<k��w"ڧ\�B���L6���D�Xj*u��C����w��l���m�B-�(�nlם�	x���Y��.�J���&m���尗��r�w3�Mw�	��C�p�.��>��� N�x6G�N�ŀE���M]���t�m`�ǟ��Oy�۞Xۑ`R��˰���v� M����`nE���h)e�E�;(M5m�{��9K���~��	ݏ &��	�*J�H��6SWm�mȰwc�	�<v�,�����v�`�ІR�aƠ��wbB����Ƃ��4�hd
ʹ��Ś��iZ�ժ`�i���y��;{��T9d�s޻�|}3��33.HkF�L�k[�N���iç��@A��Ȗ� X�gڟ���ܓ��޻�'v<�RF�x����튐��o ����&܋ 'v< �#�>�֊��J����kܮqz?y`�y�ݏ ��� ����v�n���1[X;����<��s� ���z�z0���k-.2�f���ԝvui���M�n4u���5�.��l�^�0��	���ŀN܋ >� �4�ڡ�N�M6���,v�X�dx6G�w�V��+�)���6�X�dx*�*�#�;�ذҕ%i]��eզ� }� M����Xۑ`��.]�h��t�i��dx{{6�X�g�v���o�_@X@Ω.X��U�
�o[e�яNz=~�3�a��xS����͟C�X�Vi���<�	�"��#�	�<�Q���˰�N�.�mȳ�*�����x{{{�H<ER��n�7`�1[X��� M����Xۑ`*�+��+�T�v�i��dx{{6�X�WU����2�#�5wAK-���4շ�w��`�9^��_ w}�dx��-6ݫt��-�jχ^7�U�ͳG<BM
#���牶sg��ΊT�H���e4�M� }� M����XiJ��q]��)�t�k >�=ă��x��,mȰ�K���vU��:T4��	�<��� �r, ��<�P����m*E������ �� }�7fV���R�j�T���ݵ�N܋ >�	;��ٹ'���n�D�1���1Q��~��[m���n��)��F*@��v�����]Y]Fx�̮X�V�g�m!�����{[����/]Uy�v8sv�.���n^8����Ml3*�f��[Z�IvK�lJt$�Af�њbhn��w4�$]Zv6
ʣ�R홻)&�Zt�eֶW�g��B��m ���nEk���pk�q�e�[&"���0��EZ�ad8�)�,�N����UA�8Y��t�Ҝ��ki�s&
d��6�0�V6m��"ĸi�^v�t'S�LsB`��frT�$������&���;�ذ	ۑ`*�+����S�v�Mٕ�w��`�"��#�5M.Ӣ��vP���;�ذ	ۑa��;���==�����V66SWm�mȰ���	�e`��XiJ��r����j�4���#�&ɕ�w��`nE�w�˸�;���,ZAkjr�l둋���L. %I��
ƣ��.�vM����:T4��&���;�ذ	۝�A9d�}�krO����Z,ɪI��4nI��w�(?��D U�﫜���v� N�xݙX�Q����];�l�k �� w�<n̬��R5P��m:-ӵl��G�I&V��/ �8`*�+�R����l��x�2��d�Mp��c�=\�݅�]����Qn��-�1�q���p���#���aƞ�<�n�ĵ���'v�um�&��|v��I0���	6e`v��Ą���l���X�ឮUr����{��V�nC���t�}>>�1�f�g7�m��}��;߻�s�@�CJ��t���R� xA�ތXTb@���hZ�c��6p6�賁?eq�� 8!�`^�	�X�28�H!H3X �.ca	��]� \@M�( w@�'�'��s��	�7Q6��)��H���d�Tf0�K-:���Y`)����&��WD����XD�⮍ �7��؊h"���8
t(�x����@����T�Ͽ�4 �6�E^�?�`�� �5�]�<����ｿM�<�����{ޙ�s2Bk�Y�lA�lll}����A��������A������6 �66
¬ ��￵��A�A�A�A���?��Ѩj�k%�y�k޻y9U\�������;6e`����J�1�m��|��ÐWŷAQ,��Xf:\Gt�#	T�:T�1���x�x���1o;;��?� ;ݏ �ٕ�ϐuo�x��D#�c���ـ�ǞH�Oe`[�^���Ewp�ۢ��n�v��&V�엇�JK�� n�<V�Җ[��+l�[u���)w_��	/޻�O߾�%?����??������M�����!�VS�jۼv�X��/ �+ >ݶ����F�LT��kSXc��X�4A���x��ږ�D� �=�[2�]+�E;v:���i���ǀvI��|�%��"�;͓,���
�J��xd�Xݹ�ٕ��ǀN*鰥M�]��`v�X�̬ �v<�&Vݨ�Eݤ+��qݻ�7ve`{��M�X˲^�jr��:h�V�� �v<�;�{����� ���r�U �J�V[|vp����K�b��,���ƺ��h��j�R�6d߇�|g�ۍb7X��tčr�免�K��Vb/a�CE�0H=�KAmJ[٘'M��˱��7D��Ƶ���%�m*"i�f�ij�C��2�i�ڭ�9,g(�mʂ����d;�,6�42�l��f!�5�η��v���h92�؁�^V��;�躣�2�v�.�D�3��s	l(Ė'u���;���46�	��˶��grW��G��H-��_uc�������d��� �v<.��R�Ct����6� ��"�>�p��c�>ݙXݢ�$�mU����� w�����>�Ȱ�NDK(�VSWwv� �v<�ٕ�}ۑ`n�`�ɕt+
(n�*m�n̬�;��_�� �v< �H�5i�
����hqL��d��Wsu@+�՘,�s��Fge�d&R���H��[���߼��\0���r��r�A�=��l��i'm�*m`n�g�I�� �d��'ob�"�[e+��-��_�0wc�>�2�	�ذ�`-Ԯ�m]����X��+ �vK�;���ǀE��IFP�]�RV�n��d�����x���{��R_�I;�͸ͽ=�h� @�����l���e;g��I�4���F�Iګ�Wm��=��X7c��G��*�������@y(�n����۬ �#�W�y���,��+=T��S��XQCt�����}�nI��������ł�Ε��Og�X�{� �*鳊�v��m��"�;$��	�������|W�ƛ��v��L����<� ���;r,�r�ʖ�ݶ��\;�����]�۸i#8P7�d�[R֬�4^��t��Y�%�pƓu�?�?����;r/s�U�|�g����)�f����J�| ��ﯟ��t�I��Wf�߿^=��0wc�Ur�T��)%�SvZ�Ĭ�m�^�� ��=Uʤ�'� l���(�0BT����k�ų�� $�xݑ�}U\|�8{�����;Kh=^Eڢ��7wwl�ݏ ;�<�$��0��+��;ﯿ�,TtR�l�.��6ئ���]�kxtSLf��r�Nf����?���~��.6�uVZm�{���<�=��y�����WE���-�m��?URF�?�<��#�ԑ��/�ڦ�E���g�� �������vO~������#�����[CE_�0<�������	���g������N�/�t����#�?W9��{���'�?� M��*�U\��\��U�W7d`�ά�ݮ ��.�[u��R{L���5����1�p�8�m,���iz�n�*�ς�i�8��p�jŶH�u�biYWL.�(�+~\}���.����)�Vkť�ϝ��v��\%*��f�m-�$&!��krָ�+S6�0��T�j;a.�7
A���;\������7��Ű��6 ��v�9M�S�8r�]I��/�i���d�d�m�i�������c�ϝ����`���Y��C31�v��h��5j��<�����d�� 6{� ��y���I��ݓ+=ʪH$�� l���r,�9\�$m-���J�]��wwm� I�< ����W*�Io��X�{+ �T�,�ذ��1�����t��m���������,�&V�U\�RO<qV��
�ںE����r,�U[=��	'� wdx
�TM0V����	��e8:y� ��s��ù�p�[��tIi����{��μ��i�M[����� 7v< ���$�o����a�]�T�tl��'�}�o���"tUhdh�˾�{� �_���p�r�:�y��[��M6�g���Ȱ���?U]�~� ����v����cao�jշ��]������ n��=Il���Db^�vP'�wm��0)=���y��"�$���v�v��\Lf��U�g�:�z��5v(,���iV ʙ����wш2�Z�N����u��� ;�<�r/r��A����6���Uڻ���VZm�vG��\��ʫ���ߖ=��V M����U$N*����]"�V�{���䟾�vn`�銡�B(��
(� ��"�_�����~x���}�h����]�X��s��{<`�����ʮU/k��ժ�G��մ4r��ـv<��s��{��=��,�0�5-����J[b8�`��:ȓFX:k��3b]��ASL�����i㜮��Jܿ l���r,�=Uʯ�O<�`%w���|V���r,�r�6y��	'� wdy��G���+UhO��M]����V M���������������
�-:�wwm��Ľ��[�O��krN����Jt �P���(N����ύ�:��,�C$�!Ֆ�xݑ�����������'�~��ݏ ��$��I7�Wl.�ZM�7E�"�M���v��e�*���pOj�C��G͹�"Le�-�m�}~��;�e`���_ݰ'�~x�y��[�EӺv�˶��Y�W*�	'� l���܋=U\H��^�z�m�CE_�X��< ����9ķo�X�{+ �`�\m[uwO��4���U\��]�~��	/��wd���N���}�ݷ��m��̣�p��X�������� Tr���ܮȌ"���!1��B$"B BHBBF"�GY�B�LBF NE!���8q��`�`F1�H�"B+,�HD�, �b�H�1 Ł0�~9�&��P�F�VV���d���0"D�B�$dV$1�&c ��`B1�!$�B2�ĀV0&(o����6�!�B��@��5���2�
0�X--�9 B �(aH���0�&�d����6!H�A��� F$bD�@�!�B"I;�3A��MT���D�H���00����e�0�;y�>&�A���hжV@�]�m��T���̅`*_�� ����I�F��ؠ�ƭ��$	��4Đ���#!"H�0c#D�Y��]���JQ#
Ţ�	L ŅbĔ���)23V�V�,a�b�����<9�%�,I@XG��i�+1U5��e�R��~)&�:����<����+Sj*��i�z)r�n�{���6�����P�Wf�#�I�j4-I�sV�`���ȍaR�;N���N4c6�L�2��������;�e풸3AŤ�*�J���-�ƺ�U��N�,a 6�U��v��+��s�����<��YIB��#V�¦юwE=8���(�C�v,m>)m�1���.kIS�X�Vs�ۊ
��o5�c���аٸ0vY��W\Ǝ#%�V�5��[��ؓ�v6�P�{�*���L@��Y�G*i�lc�S�{[G��7aH�-u��ŷaI�[,s�X^иs�E�vd�b��{f�,ge�dU�-�����{uf[N��w�J�n��q�4�ߟ<�\l6pI�l�U�Y�&Pfb�����s\�&řzz�Q�fWi�ʹ(��rJT�UUV��'GP��1�3���ZM��k��0�z�	]Yܛt����j�xN��&�\b�l3,q�j%8�Q�f��X�ձ���ܜ�uil�d�YL`I�7 Ԍ�њYVk���뭠5� !���V�,�t��<o�Ȁm��)q��"��
4�M��G-T9��U䫮�{[ĽWg���
P��� jmU��h�6�O��-�v�jn��4ږlm� Km۷�wݷ���ⱋ���]�l�.�f�; j��:��,�L��,�D��۬�C�z%���m��(ӹJ�6�zm��'
3�����;��r60��%�)�ⲅ�{	�	�P#�	����5�U�VΡ����tn���	$+i��r��4ĀA�yA�2�[�^���[l����)�m����˲�ۡ����{(A��P����*�G��UnC�e\�F��Vړpf�ʪ%��H�M�!�k���UUN&f�pi�F�d�������Kau��)�s�>F�ـhY�
�Ϛ����,6���l�Oc��Xp9Ӗ�������HH}�c�*�x&��,5Mk1AF��E߁۸@�
����~ڠ���\=u$��v�Cl,"�u�P�W4�����ٝ�"�t!l��ai�zuɴb�-;7j*v�t��ڶ4C鎥�Ck��8�`I��x�e��e���]�{ge�� �����d�-q4t��5��I��.Ŏ7Y�y�S��5�m@���v+Q�<N��89{v栥��{e8)x��7n��b�
�h���5Av׍���H]Rt�q���Xpd��T��kj���t����y��ga�kђ̶b�k�љ�u�iݷV	�5�e��xr:8��Q�[.+��uwl��߽��� ;�<�\0��D%J��U�wm� ody�U�s���g���~0�X�]��
�[-6��#�;5�r���]�~�����<x�J�N�H����徙� ��e`�G���y���wt]۫i� �ɕ�yn������;��l���e��0���B�Ó�ӹ1�e{/b����8��[s�Q�m;Z�k�i�մ4U�[u�� ;�<����U���V�g����n�E��j� }���>��$�$8�@�Iݏ�ݓ+ ;�z��#�`%w��$�&�ۼ}������ >�ǀNѣ��i>v�զ��ve`�G�wc��r����<`��<��
��U�wm� odx�v<�\0��+ �DSW.�t�I�tRWFi�*g��,�shA��@M)�.X�e�D��:2^fX��V�ue�����vk��ve~��W��;`z~��qC������n�����9Ď��V n�� >�Ǟ�+��H����weһmҴف?}�lܒ~���s��`��Pu��w��.��A�n��|V�`~�9���r�O~x�ߞ�c��W9��敏�ey~EۺH�6�����'9�fC�;��X��xd)��m&V�7'��蝜v��#<�\G��v6{Zµps�5��e�-����g����￟ǀ}ݙX�����ݞx��O���[�ڧV��ٕ���o������l��Gix��]�T��U�wm� M�� }ݏRZ�=xv{+ ��IV���B-���x����~�/��x�ن�?�,P;]��ߵ�'[�w�Lc\t�ۻo �/ �W������� >�ǀH�D��^4e�Y��ͱ+����O	,N{-���kfA����ڴ��&�����e`�c�����o�Ͼ��~<'�dks���0����vy�[�^�veg���ey~�V�$>6����<��d�<�v{+ 7g�t�0�wi�V����d������G�wc�'h�9iRl��N���wfV�UŻ�?�;�� �엀e�R�U*�R�v�A�m飀3Fi�P� ��i��rh<u�2Atj%:�/h9���R����[���pX;(�@့kp����\�H�0��U+��x�۬qٙ^W�pg���;zVD��b+.�e!fU�[�)��v�%yWmbN�x��;<�$[gm�
U˸��H۳����9�!��r���}��nE~sn��@�C���qs{-�֧4��jy��Pm����Vն�
Ͻӻ�0x�����9У3%��5ԵGK�XP�CE)\[>d74���(�[��k�&��������������~���u`���M� ��z�5o�xv{+ ;ݏ;�wjr��Hi�1��컰���8���p�>�ly�<����v ~�ח�����U�����9{���$�����]��Kܻ��{s�o��v�T��k�2ð ���^p�7��;����np�3�; 9����\�
<��l�5�:��<Ah��b�z�2�1ϥ��	��w�>,��x�B5����۞w�$���|�]ۙK���In�?� �z�}�a�.%0�w`7�}��9ʜ�Vf)��)bI%$���]����T뭰}�������j�F\�� ���p� <��8m�7�;���9��{*{5������|�� �c�I%�r/�I.�̥�$�6d�v�d
�댼��y� <���� ~�{�; ���� �a��s	g��v���r<��Z�k�����a��,�Z�nG��ѐ�0�4�Kb�.�����3�$�����$�oc�I%��qq�wo5���� ~�>ӿ��������ߝ����Ns�M����o��0��4� ?}��8 ~�z���y']N����g\�����e,I%�ej���t­�Le� �o~w`�>�s��������� {�m=�%Y� j�v$�޽��K�s)bI%$��Iv�;� ��O���u��*5 �ȅ4�V�X4�W���a=�� P�崊˕cF�u��ڦ���RKe�)bI%$��K�gsNl�?|s�M����Цd]��KI)$|�][2�IH�_|�]��p���P�����[���mֹy���*�$��E��ܻ���,I$�=����o+�f�Qqc�3v�}�|s�_������{�{�rۇ�j('���=�݀��ݖ|�\3P�T� ?y�jĒJl��K�L�ĒS\��K�*�~����6eؼ�6��kB%�]��Du�%�R5P�J�4Bk���I�x����@�5�|Wl]I$�{����%�&U�I)�E�I���s�; =���J*�=!L��$�T�W��r��v�����$���,H�=��>�u�]M�����\�uT���v }���8���p�>�N�Rm���� ����� ��Ӏeq���Q���/r���/c�I/zy��Iulʼ =��Ӝ �7������v�a� {��I�S��ܛ��>�s���v]�m��@H� E�N��w��K��7cvg)�n��/:'���.+�e��9�Ʊ�������7do3;4�8�e`��+�b�[0��M�f��p�mΠ�KbxM���^���z3��㍿>���,�-��ʰ5lM\�-�T4�#�k&�!ۂ�E�l���nϓPI�mGk��z1���`nC�U(DӸ(<�]�܆hɵ��wV�ihAU�E�^ͻ�Ԝ�f���n&F��n���n��uzέ����^�v+�����W�m�l�P�U������ʼI%5�_|�]ۙKܪ��i%�O?�H=�{_���5R�f� ���Ns]��o�ĒK����$�V̫��Kg<w�ȶeu��8���������u��x{�sv }���8����oe�wF�;��Sm��|���݅���{y�o���!��ߋ�m����
�p��y�Ǟ�7`�I'�w��z�[-�X�II#�䒕.��>���>_���Y��ʙY���{aƷ766��tC����1�˪���f� ��Ⱦ�$��2�$�Rl~�r������������.0њ8�%2s�����T/X0���I#�z�m0ۡ�T(Ad# �B�UT�"��젴��#�4�P�1@�b��+� �Aʊ�?�Q;�m�s���-���홻m����yT���5/��n�ɝ��; ��� �y�sv�*���*�Z������-���K�m�{�y)�"�3n��� ~<��� =����[o�]�v�
 ���{��-��vz^�J����݀���� }$�u&Ǟ�$���?�I#c�ĒK�R�}�O����%����H�e�J̀�7�a�vf&X�D�ӧt�o$|�ٳfY���Ԓ���bI/�I|�F���Us�m�?���3]��6�e��f����$��I#c�Ē[�E��%��R��_�Iҡ�͟�@��g�8]� _���5�m�}���l`?�`}�]_Ii��5#LhB+�B���죑0�d$`I\0͍.cP1H#�Mf�3)X	YT���00�M���u�� (�	�7)	�i[mG{y+���sc� S��Ƅ�A�!�В1�H�rऄbH(DU0O��@��
.�X�S��| � @�)H(t6�Up<>0�
���������{�� {�e=�sV. :��^���=���%=~�X�IvH��$�=}�`���~�ah��)�� �s)bI/W*��y��$O?In����f��fk��8¥�ԗg(]���dv��ӎu7bA�M]s
K7�!��xkIs��wwm|�{� 6H��ؿW9_�a���� ��~��
��%l.�n�fǀn�ŀl�� �\�=�$Nl<�7bv>]	��$�y`/b��W껟���y~���'v�e6�M�V6����X��, �c�\�ے^�b�V]��IP_��ۑ`������^%�X�r�U�J�W�h*��izĤ�S#c.��s��
2���gR��=��n*^|?<)��������׀uI/ ��/U|�K��펅�n��v�&Z�xT�x��`ۑ`�;Z�E�m:Tڻ�C�x�8`�"�ԑ�y��=xv��D��[��f��M~���� �엀}�� ��fR.�bJ��؛X�����W��{������7�=���v��٩��m���@�6�"���ӡ䱷u�:�e3J�������!��9M���e��!��}���ݭ�%]ũ�8J֐�n�F�Od<�G "V�/n`���pWR�En���E{7r�6�.L3v�9�.���ʁ�i����|��,4��Ȯ�3�WG9�B�R��nF���g/0���7O�.q`�^���t�ҵ@Q�5��\7em��w�7�Zy>R�jgil���fqj�s5�� qv��'�����&�A\`�f"V�9��	v��c��(M��"�߯ �c��� wv<mU�Ҁ�I�nۻw�}��=��7o�X�y�]���ʮ$wb�V]��v�AWL��v��ݏ�!���������>������C�)�&c���[k ;��6^��Us�ʥ5�,��������I;��|���=�W9U���x�	����ǀ�w�E�i����R�U�y�b�e��F�a��{��t��5�ԂɎm]ӡ�x�0�`wc�9��9�|���׀l�q��X�[��m��	��ٺp��4F$Ҫ�U^��\�9U������5o�׀}�� ���H�E�H�uv]� ;��엇�ʮr��g��v��w��N+�XS��P�x�s��9W{�[����ތ'*���wc�<�<z�Wvwn��8`�Ȱ���]������оƎ"y����rX{7<��Xu�����.���:t��ǆt��[52�>v���ǀuM�ꪯ�w|�`���j��V؟e���������0�ȳ�ʤ���S����>$�o ��z��0�]�p�p�Π'��=�߮��{�ܓ���;�fV����:��>��n܋ ;������^ݔ*h���Um��0ۑ`�)l�����lp�;*-��q��glGA�˞�c B[h�M�
ˬ��P�2��#���o#�4l�ˉ� ��xT���8z��_������-ؐ�K�o ��/<���� �~���ǀu4�-]v�vݻ�>��}�"�ܤ���j�׀}���-;�N���[f����vy�[��;]�8`�V�U*Ҷ�O���X��x�[rz���� �nE��ln����tU����Q���=�XC6[=a�H����%�gM&�+|I�v��$���v�X��x�Ite]�MmZ�E�xݎ��U�%���{ߞ�6^z�#�(T��E۪m��0	��, ��xWd����@��8�t�X���O<V�׀}���U~�?}��''��-ؐƂ�&���/ �\�Wg���n����ǀP�UQʢ� �Pڔ
,V!@"�Y�~�m޳l!��8��M0MV�Ҿ:�u�J�#c��v�hJ��cu��n�^���5/<�n4FZ)c,q�����\��g�A؊lzv����n�8��+m��s���M�VʹlY�dvӹSOV֛�����r��_�үL%����2�J���h;b��ŢQ�.� ]��f�ʶuJZ���vl�b�U�ZU��$��:y'L�xn�c�����N�u�+�[.�]mX�Z�4)�؁�j�2�"��q��˨Wi��j��7���������x��N�7t5iժ�e�`�p�r� �<�[=x�3�\��m��_�iSt���`��}ۑ`lp�;�p�>�e��&Z�Į˶�=UUK�����}�p����W*�s��]��� ��Q�14+�g*�V��c��u� ;ݏ ���`�J<���-qM���V��@�L6[pH������v=�i3������,��qxّUV|v?��xݹ��\��Wl6~�y+οQwb)��ұ�0����SP>�t������}�vnI���g���W7��ܴГ
`��s� ����wny`����j���X�Yum����U�]�g��s� ;ݏ��qw\��;"�g�:�WL����ŀ~�qn�?�����>�}<��I�ֹ�ˡ�*�l�*H�U%uԥJ��.n����fղ�?�t���m:���-�����>��X�\0�{��RZLN�+|J�+f�ob�URG}��s� ��z��'��WWN�4Uح������Ň�� ȁ�l
�0�D?���`���hT�V.��۶ف���fx�&�� ��"��\������y�=�Wv"�.�*�l�;�p�?Uw_����e`�`-�����XO����\1R��	���.%͵���q�8k�C
c��m-�!�l�hV�#����� ��e`��Xݽ� ;��R��ݱՊ��0��+?���\�"��x���}/b�>�W7`�v]2����/ ���a���+������ ���X{eDF�O����&��{���]�<�'�g}w$�ﻳrl�!�T7�k�����-���J��]��}.E�~�~�Ur�}�ݮ��y�0��,iI`�bG�[�����an4AK�Vk��.!̶��P��R+r�4f�8�m�|�ݙX�`n�{��s�����wҋ�i`e;+�� ������:I-?�~0��^������UW7�S�j��J�Ҧ�d~0��x~�*��v{+ �����Z'm:wl���۞���{+ ��ܪ����yD��[m�6��wfV�{I9�>�ܒw�w[�|�!T"ӝS�;ǰ�	������Rl�I�`�*�?~u?(@�����\R�F!�H��b.�3cO�M is�@��q���-,���09�]�B  X�XRa �YHR?+Q���N�t��|1�����4�VX��G6DM��4�8���0�m:{1��E�b�G�'b:w,�*Ջ���^NױUJ�%�(�&wIL��i<j5=)1h6PF!OIjz��]��c��rQ�'6�1UQ�1��və�{Z��W]��gE�,=����\��V����ɱ͕H��#��K�h��Y� �yM���O<�J�$��G]�퉃����h��.�!%A*�P���h��bQhQ1��CgZXPy��+:1�oc�m�fнL�c��g8ƭ��xS/�����hv3]�	۞�х�<=�c�ؒ��#c!��z��΍�B=���]��V��b�q�pA�k����n��M�� �g���mnܰ#����-� [cb[:�J}�"��l�;2�)6��d6���GR@9�.�ݳ�WFBE42���RZ�� �vABtnȦ˚�2�l j��H��� -ڻ
�F�S#�Hm��.N���%��I��9�֝2�Y�즸��,5���f2�ی]��h���S�[xS�oJ�����&��K�M�.��v@#�������hǛ.ch�1�;cX41�Sk%�`!v�,�P.YU摹Z�8ف(�n�d29{�yT6L�-��b��i	q�5�n
sg 7P�@�ut�/��q� ���ڎ;#�n�����6���WL�l���4�|�f�K(��Fy3eЍ����΋b]�Xw'e�8�94���07]tD��5;@������S.��WKڀ���t6ٝ�.�53�jB�SM���%�����)��Z����1�̹h�vA�"�����ˡ�N3V��pY���lY�Rj�;.f��/jy\p�Ike�Ř��"��U�� a�S=�P����خ$��躎#]뎼�dj����1�^J٬�@���VU�;y��B�l+��t���[W]mNtksQ���Vc Q#[hqڶ��UUUUT�*ҭ��eaڎhY�H��@��Q���Nubm�A?(�~C����~��l����MK,�ڹ0֌��SrF
Ԧy��!�8�5R�/X�y�zs��J2�$1�in8�Z9�rl*���Y"�l��ʲ������
�v�PFGp����e���K�;����'���%�,��k]�,�.	N��A��c٪�X�DC�Kb�d�Ճ:�H��9Bѻq�։h��n�r�]�6ren��+)躙�����k������טW[vat5*�$��n��:���H{m�Ezp��2���'zǻ�[��%WL�u�zG� ���`���N������￿�O �{����9Dy��f�ob�5M��}ݙX�p���N���_?�����]6�a�2wm������&V�\0��,n�ȇV�vq��%m`M�X�p�7��`/b�>ݡ1Eh����۷n���ou� �{�ٕ�~�KJ�n�=n�vf��%�u&5ӊ��t\D��D���6�6�7����=��R�����~X�ذ�&W�s�_ ���o7��SR)�y������=��I��wJ�Ǯe`Kذ��,�A8Q	z������Xw���6^ŀw��`��}үH7e�b���n��ذ�{���ٕ�N�Q�ݴ���0�{;r,����&���D��'j��VZ�j��̦9b̝rGH-����u���站��f�Y�we�E&
��"�/ ��2�	5�ܮ|��s� �P��tX;8�L��}�2��H���v\��"�/?$w҄ҥ�
��[nݺ�'��oob��]mW70�1�I2�y�-U�,�wN���,Wd��+ 콋 �v��U�i;l�]5m`ۑ`M�Xe�X��,V���M1+n�rne�J;yu�i�\�y�p�1��ͭ˱_+Bv۱����}6e`��`�ذ�Ȱ�U���m���[��\3�ny`o�x�fV~H��^E_�M�@��m� �s� ��/s��W�]��~��'�?����#��j���[X�ذ����l�ٹ>�[��HI�0�M_l܁���1�1�j �`�{�*�Tء��=����ܓ�zM{.�2Md4%N�������l�v�X��o����3v�6��ݔ����)H��Q]�	�/]K3	t�%.�� (��o![hy���۶���OG� ����,��y�X��]'tյ�M�~���U����� ���yX�ذ	�֠U�lV���V��\0����ܪ����y`��,x�[bR�ct˶�� �j�Xe�X�Ȱ=\��U)��Xt����;c�,NҷXe�X�Ȱ]������g9�V�r����Ν'��j�:)����kMl,��V���U뜑'.� ;����� w8�y&`ס]¥�Z��ĴҨ�6��R:3URm�A�V^���<�������ѸS;mɌg#�Z�7V���ev�X^�W;&-�;Et����M�����68n�Q��U�����&Ś�cA����H���F�vG�ˮ3˃f�b�@����yӧ�;�>y�.�f�s���nm��s���^Dݝp����hK�=TmZ�uH�f1T�S���~��vK�>�S+�W�s����O��e���wM0O�m`�%�n���vk���~���U]����Ҳ����:.���/�Xf�a9ĺ�Lfǀ}�Bi �vr��WL=ʪ[7!�w��,�r,��yX����1���ˑ`��z�w}{����A=�sP24&�7C�k-\��ZGWYq��7�s����]���#˨�š�}lV��w��,��2�wc�_ ��X��H��B��1��k �M�X��)����1rO���rN}����ȳ���H�p�7v�[abv+u���}/b�5vK�>�L�vʔ���ݠ|M+m�z��z9�E���H�V vlx�Ѷ\C);��B��Se�I/+ 6lx�"�}=0z�b���18��f�b{��E���cuq��m��¤[���k6�D�+k �E2�fǀI{�\0�hLE*�E���v����{�⥳��z�I�w^��s��ٿ��y���IZ)�]'cV��\��6k�=J[k�~^*����}��l� ����:�\tյ�}�"�>�L� ��x��)�<�s��	^��e����2��d��	�X��x��������j�-���W=8��v,��^k)��#4��F;0��f4Zam6�liҷXٱ�/b�5M��}�^V��6�q�۴������X����K�����6ˈe	��
��5vK�>�/+ ;6<K�`�8�]��`�E�0����6<K�`}]�9�S�9\�w&N�`���.�R��R�v���	���ʯy���=�~0�����q�mm�L�U�ns�@R���ol6Wf;[�r>��
�N�Y�ΎN���;��	.E�I��K��	6<rV�e�tհ�:j��$����	6<Mp�q#��t�W�;e1�j��;�/e`��Jz��\��7�0���n����+u�lx��`^Ł�W8��/}X�����n�HWm�Kذ~��=�vI����ٹ$�~�$��AH�d �=��lKR�u��\:v�1��X�ZLu����K6�v'dR�Cm��3�D=[���0q����/k+b��W�I�2�ㄉ�wm��J�B[5 �7�Kn��up(l�y��m�ͦ4㰎�&�aD�����a9;#�4��p�^�ͳi�pi=Pwom�<m�f4"��v$(���1K���b9i=��t���gH�|���a)shJ���Kb�S.%����IA�cuFf�%�������5�Y/k�����}"�X&ǀj엀n��wj��cZ.ـ}�/+?U$}�I~��;5�?q#��k��[�wnӷX7�x�Ȱ�p�>엕�J]��R��e�v;��ۑ`��`vK���8��y��Tk�cV����ݵ�uM��}�/+ 7�<v8`��U-�W�E/����5v�U�S�mb��c�3��v"L�kR�F�A�I'�F&���t�]�v�@����`� �0���� �ӫ����nI>������ ��c�B�>��7�p�;�Xݒ�	ڳiZ�ݶ�>&��x�������\�).�yX�O<{tl���->Wn����>�S+ $��=�W*�J^�׀Iy�WN貘"�V� ��L��{���"�z�	/b�>��|L ��^��[HϱV��f��[�y[7�^�@6�����$�ѾB�<
B�GgZ���O<{r,KؿW*���	K|/RUvr�X'cV������ĉ�X}��{#�6�9j�]�t�l�f6�,�ea��qr��*�v�� B$�(��1xp>�IVġ�Ҕ��ȐB� �*P4��1��Є$R�E�~"� ��T%�1I���4�(~��bh����
C[�?-7~�����b)b&& 0C ��@�$C""��l�*��w�	ο'+k�\�WGY���ۑ`�WKP�wle��V��s�9{���k ?~��l�� ��,{�6�6˻IҷX&ǀz����z���2�Z��ֹ�ˍn��V<���몜uY���xG�deN�[��Ty��Z�ZM��}��Ix��`ئW�@{�� �螢��jğ��w�I{݉� $��RK�7tq;�l�VS������ I�����l�� ��>DpV�۴�� ����"�?^��ܟ���"0�]�s�����`��*�V�SUt���eȰ����L� ٱ�����fXO��>b�Y�+�������u������E
�uɞx���쳍��أ�"�����X�c�6\� �U|[DN.�v� 7a l���"�5M���H�<[t&�դ��cx=<�RK�5M���� �՛J;lm����o �$�e�X݊<r�IOO<K�z���|Wv� �l� �b� 'dx�&nI�/¦Q@�� j�QGLE
X�T`�Aa� �
�� !j�F���P VQ`X�T �@"� �e���d��e�Bu��n����TR̓]nH՚�r������0x2@+G��u��3q�kq9ٟu�:^-sõ�,�]�����6ٙ_'�6���[v�v��ۓ7m�0c�y�y���c����WFaA�i�[pK����T����hKR����2�!P�;K���R���d]�����vR���1	b�f�jM�Z�j����y����-n�rK�٪�j8�ƭ��7A���B�4A,MF��[�S4[.��Ī�V���(�vG�j�_�A�=��o����T���7��<T��	�2��w��A*�]'cV��d�M�X{��JO;��zy���+�vS��ӷx�2���, �c�5I/ �U|ں����۶� ��q`͏ ղ^�fV+jZ�i̦ƁV��k�YCEf��G�✅e��w5Xƺ%�oY��+r�Y�p���|��^�d�f̯Ur�A'��`j�K�QF��U���}�='�!��$+���9�����ﲰH�� 7�<v��E[vՉ>	��� ��+ ��qa�${}�E�z����n�]�)*t����Kg���zy�����{��V�� ~8 -�'n��X&ǀl�&̬�ŀ|��J�ӦX�z���ÈEt�D��n�tp�s����+hf[�����r��w�� �fVݎ���zy��yԭ
�+t�؛X�2��w I���K�$��m]\V�b�v�`��X&ǅ�S�]��/ ��+ ޚ�n��V�%NӶ�<��<���x�2���,{Vm(��&�ⴭ��j�/ ���W����O;��	�����@�5���C�]��p�6�Ƶ�XK.�8-�������uq0���v�ݖ��pM[n����VݍE�v<V�x[�)N��.锕4[u�wcQg�ăޞxS޼M�X͡P�E�J�U�N�w�lxV�x{��^��V���x��*�]�L�an��x���	6e`ۊ^�
�r�s�EUA�ႀ|x6*��{[�OsP�J��m�6���$ٕ�~�s��_����:�K�?r���r��Z��tj{>W�<jg=��9�c7l�n���'V���Ѧ�u��P�Sg,��u��lxV���s� ����	�h���ۤ��T��� $��[%��lܓ�����W��T5��d?���.6[�`y{���>�t����o ;�c�7n��
ݖ�[�m+m`�2�ۊ^ vlx�UR�~�����t�J���`�� ���.E�Nɓ��N�;��&�R�}�P4q���$A�*[s�vL�/5Fɛ���N�%j��p���^['��h���d�!��H)6��̛d��5�n�̽>�c`0��n�Vwm�R77V�����1����On��p��X�v4f��S�j
�u��-$�!)1���
�Z��)s \b�n ŉ�;98�d=��sM͸(_V���&�4U�/P��w9���ٝD��%n�틫m��ǖi�(ج�Sf�j�7gb~���K/� ZJ�U�'e��	��v\� ٳ+ ݲK�%.�A]�m��XeȰ	6e`�Ix�L��_�����~C��[;
lM����v◀}�e`.E�wj��WI+�r���u����������^���+ �r,��+ �Mj+���V�&�w�}$��:���ove`�Ix�bWd���-�Jv���Ų6\)ڴ�mf�"��HX����[�8�2��5�����{�+ ݸ��ve`�
�mZN��m]�x�YWWvn�%��XT����Zut˫�e%MZn��$���+Ԗ�{׀o���ͥI�- V�bv[�{&V�$��fV�d��J]��]���an�M��$���+ ݲK�>�e`��:~���CL��*�G��9xj�)n��N��l�.���~��Q.�w��z��T�)ۻk�{����vY%�I2��%��Wͫ�+��۶� ݲK��$w��V�����2��֢��M�E؄�n���XT��|�Wy«�M�R��"��"����;�k�6`�?~�{em+�+Ln���v��W9�Uqm�޼l�V�d��}6e`��j��I�m]�x�fV��U�a������XT���J%r�i2�X���bP����Q3�`��hlO(E�T���i��MU��4�^KcuY�~��v�ٕ�v\���s�Oe`�J����4��x�&V~�s��$o��X��v�/ ��	h��w�L�m��r,wfV�\�JK=��;�{+ �ȇV�5t�)�6�ݙX�d�srNw�ٹ7���3s"�� �� $:h/����~�ܓ�m{���T���u�n�%�I2�ˑ`�2�]���F�M]�ݍR�K	�ѕ���◯<�c
b3c����h1�Xր��mӺ�E؄�n���XeȰݙ^��{׀M��YJ��m;u�v\� �ٕ�n�%�I2�톢�M�Ҷ���+ ݲK��R]�����y���պu`���m����W)H�z�o����</I� �JT��j���Z�;�� �I��$x�̬v◀*��r�U��$ ����0�s�H�M��$X0bČaH�wjɤ�5�t-FFK�������"�i2B\!��J��Z+ �/#�r�!3�a�h6�%�d&}rBb#�� �m�FbFa0�	����ɤ�� ?���͢
��s�](D≥ �چ�`��� B2,�c�(P�"�k/���hg�}��#�4�!#~��6����!K��{�h:L �`wU�S}��hC���|����G9PV���TSJ��Q�ܴ%=+���Zl���`}(su�tR��:`�v��Þ�@s�p��ű;xͩ�8�0�݂�F'�6���ۭ�㚋F�q�J�m��˱�s@��`�ݰ���<�LY��!A3=�D+���r�ͅҔ�98�gX�=-;=�� �P��fzmJ�Nk��c���X� ӈ�ї��2	r˩(L!�R�v�&s��v Χ=����Z��C] nP"�n�:����f��Nm�1����E���|�y:��<���b�[�p@&�m�Z��|�s��X��)�'���[+ZnI�+�KFښ)�n8G0���q��[][]Y72�A������r��-:J�k�K��쳩�j78v���T�
����܂�X
UZ51�!TU�k�3�pe��:�+p]�]�2d���䇲X'�Gi�[��m�p��J��w\�	G:vf���8���h�sҰ/O\a��Ƕ��c&0ѹ�R��v�]���ŏnWI�ЄZ�re
�6'N�c��ɧ����7��$��f�ك�A��p*��ؗ��v%��$.�)�W�� �B��qT��vx)�Z���3��� �Ř��R�s[�-<��s"9�ʕDMj�Z�h :�Bg�P��TLv�.�q0uF4�{K�9��4u2B��(�X�a�v4˜�0�R�A�E��錘G8�#�oUP�,Ԛv!Õ����A��V�<�e��Qn��H�N���:�]�h8��S�+��b������A�Z�N��[[^6� �\b�qٝRSj5�n���+p@��l���s�#+v[�]�&�T��(����g���u\M-�Yk���A�+UUWA�@��-��=QJ�&E{n�\耻U�+J��q�K�4�`�m�3��V�Mf�[Zw�l�U�
`������V�^��r��8c� (��w$�Nu�zs�$�Ώ�Ӡ�*<+*!�p��(o��)���!���wC}�<��cy�i�y�f͛caK��������n\��h��4m �+M!)�g`�.b;C��N�5Gq�gm�ije��Xm�4�m5Wq1,��bY�U�鎼�mh��ݍ�uk��ɱ�	�Nmp�e��ܥڅz�F`Ӫv��ymrTV���
m���u����J�WEu�Q�5�Ǳ�����;T�5�at.S�3�.j��f��Q�ʅ���zwf>���<��hf��N�Yv���ks�!y��s�(�txl\a���R��	6<wfV�qK�s����;�{+ �sɯZt��W�4��7ve`���+ 6H��,4�%v�R�m��d��}$���\H�{� �{+ �Mh��I���-���w��Հ�y��2��$�{f��iU�m'�m;u��<�ʒ{��	,�� ��+ �r��K�*y��t����9� ��XF6:�.�,��j�pg8I�dE��.�ŸA�\��Ǉm���}����$��&W��@o��E�zն
���`�Iy�aUv)&V l��ݙXfҤ�U��n�Չ�n���X�#�7ve`�Ix��)HVZ���u��<wfV�d��}$��6r!�U��v��ƛx�̬���_�v{�X�#�	��}]\�'��xy�mA�&�y�.d�]s���%���m-4�A��KX]�&�s�����z��L� ��ݙXzkD.�B���n��L� ��ݙX�^������v�i�6������+j���9T�UV��%��2��Ѷ��ZHt�'wm�ܪ�����	,�� �I���<T�Z��T+�4[u�n�%��e`d� ��+ ��+嶐P6�y��h0g�n8�f�nw J >���ۨ3.���t�]&�B�Uj��x�L� ���2��$�R��+��5Cv���z�$���$�޼�+ �Ț�,;�W�4��;�2��$��+ ;$xw�J��	۶� ݲK�>�2��G�ڕK �A1U޳��'�O�ge5�d՘X��� �d���<��+ ݸ��o�O��ׄ3.��.�̡�[-�ױ-]�r6R�V$�&�$q�6�Έ�J��n�d� �ٕ�n�%�l�Xv�n��I�|V��wve`�Ix�&V vH�ԑ����j�|`�J۬K=��>�2��9\H�{� �{+ ��T�K(J��-���yw��Հ�y��2�=U�R3޼�.X��J�N�7`۬ ���2��$��+ �؝�Zn���R"L՜ݜ��!�������k�-��T�1���n^�m��.M���ӯ����e�WY�U5� f�q/V���"�r/[َv���E�õ�<�sb}��܉T� ʸ��^���t�@�����ţIp����fp5)���2���̗l��P�b�=q����YʵT��-Q,�;6����T�^���:�w�v�0�&Y�0�4H'o:��v�/�WN1�Ĭ`���+���{S<�5n���������n�%��e`d� �冖�q�N�۶� ݲK�>�e`vG�wveg�H�F�
���N�	�������� wv<�d��N�[J�m��-����� 7v<�d��}$��;�[qZwISB|V��o 7v<�d��}$��� �r�ʩ��.����&(���ոI�J��4u��ܚ&tg����j�9[�բ.4&ղ�P��o���۰>�e`vG��;R����چMh��3Y�';��ޅ�X R �W����O���rI���[�wl����Z�V+����`vG��Ke���}�B��]&$�Cv� vlxv�/ �ɕ���gR�[w�I����^;&V wdx7c�"�aN��dN1j��D�>�*Y9q���Q7'[T9�D�bm�Ʉ֞�x.3������+ ;$x7c�7l��	�+Qq7t�-'�M7X�#�	��d��Nɕ�wn����������o	'~��ܓ�w��N��+4@Gբ�/¡�(T�˞���'���պ"6+�e%V
��7n)x�2�d� 6lx�m;%��m7E�n� ٳ+ 6lx�c�7oe���F�ht��h��V���I�$q�ۮ�5��JĶƍ�^m�k�3�ŒV�h��v�n��c���{.��X�Z�)Zn�,i���}I�`od������v�[wƁV���.��Xٱ�fǀw��A�:���E�w���)w��Հ���ݏ��US��}x���\M�i���M� }6< �����/ �ɕ�z�SO{�li��)�z.�/[��l͈l���1Q��w����,�b�0z�l�����7l�x�2��#�5n��������[x�ꗀI�+ >� I�����R�+h�7E�ӼM�X���M� ݽR���%Wun諦��`�c�	��z���e`J�9JИ;t�i;w�v<�����e`�%�rO}���m�M@vf�Z͓]X��G^4\`��3`�cmk��l��nH�1��&�m�h�:�.��0�v?Q���m� ����6v����1g
nM���Ӧ������nvx�Օ�)ʜ&n��W]'eu�󱴃��;0�Ů9e�й��ݐ�mt��>);v�v��ۓm�#mS[$�i��nhKJ�i��W"��.�@0
�P#z���$��_�Rn��jnY��Y�ҙ���;��48C-��[d�K�$�3[p�mo.|����*Eջo �ߗ� �ɕ�j����y��<;�v�؋m;�7�e`�%�ݏ �n)y�W+��*"���Վ��hm��׀lx{qK�$ٕ�}ۭ����t>&�������R�	6e`�%��DGMX
�P����◀zz{���޼ ٱ�{��v�Ю��Me��U%�s��3��/N�C8��	=;�<�7�=#傷gt&�w�lٕ�j엀lx{qK�6�(��+n�tݴ�7$���sq@�"��C$C�B���Ur����� �ީx�L��G�ȫeӻu|�������;ۊ^��+ ��/ �A]�K�|ut�V�R�~^�o���j엀��5����jՖ&�w�od��5vK�͏ �n)x�U�ؒ/�݅1�-v#v�6� +N�K����-Z��������L��a]�L<֬������͏ �n)x͙Xݺ��6��t�I�Jـ6<����6e`�ذ[��Ӻ���%m�v◹'���7)��XO�I�u�UNE�hD�D�H����D�I@�aBb@����ѹG[�aA�Mh�.�M�IXY$�Ѝ �5$�^`H ;�:L����C[UJ�b��~��~p4(�� pW�? ��AV����x`�����+������wx�X�Ȱnǀw�%����D��]����`�"�	���R�	�2�zJZ�][-
ݺ�k�ͮ��;�b6G,�|l[�|���L[S.��u��J�"h�������}��ݷ������e~�W�&���=����w�`�V����竉��X�?&ǀ}h�n��v�m;�$ٕ�od�����R�함��(��u��7���zy���/)_:�!����Pa��7�';���[|*�;)[n�fǀw��f̬{&V l)D�U���*�N�(�`5e%*�q��4&1{\J�;J���-s�p�ؚt�`�ebV���R��X�L� ������r躶�ct[M;�7�eg�&���I�n���'A}��u/�!�lb�wm��7c��nߗ� ���XҵR-�wv�񦭘7c�;ۊ^;&V���\�*[w�J��o �n)x�2��X&ǀ}U���U�����N����)52�[3�
4��B��a6 �i�3vܬn#L�߬�| �kU�l��t��7����ي�sjl��-"it؀n��l@te3U/9��Z��R���]z��K�ې�YMI�mB%�e��7Vr�L�i�$�fݲ����"cpv�J��<8�dlu��"[�dۣF�\�Mw8J�;`�Nn
�����j�@D����k熻Ž`��H�#�^N�!�#ҳd�l5n}�^�a���U�`:�Vm�E����6o���X�c�;ۊ^���@m:-��Cn��X�c�;ۊ^�fV�n��V�n������ ٱ���/ ٳ+ �ɕ�j�-�EЭ�"�[x��[��׀{}�{0nǀl�e�@][e1�-����e`��v<����4NР]�`�U��2tqks� з�{5���d.� �0�b�\��M$Z�tU�v�n��p�	�I9�;��
���{�{f��;u|̚�Y�1���M�'~���&���o�����{+ ��U.mi-��@�M�xݹr�	�2��UĻ��`�����֞��rk��.w����M������o�?� M������'l�E����|i�� �k� M������7�e`¶7vƓ�k�[)����9�N �N�*�Z`�9ۚݓ��P�ל��{��}X%lv�v���|��xv���l�X�\0SAKi�t+e�V�ݽ�y��U�H������ ww�����g����) ���'���ٹ';�v�m��� ��������'޿_� �^تRWv���`��`ݏ 콹x�X�558[����:���	�����9[�/����V;{�����٤W歶R8�}�� ����� 4r�/t�*m��fP����p�l2�/3��
1r���~���l��'ob�	6<�#QR�بuh��v� �fVs��RG}� ���ջq��${l�Jׁ�j���Ӷ� ���ջq��2��u��Țg[�[�~��;����� ������+�(7��s��k�"�"��Ut��!����ۏ �d��>��`wc�;�Ė
�n�*m*����TG#c��5�783u���
C�-	��)sӢ��<��J�)������e`Kذ���]R<a{b�I]ۺ*��`��X�����;&V�i�r�l�&���l�	���#��9U���~��O?�*�'6'M����&̬���{�� �#^T��&%h��]��Nɕ�{���R~������u����0Q���j�n�TH-gs܀�����b�=`�\����Y�i�Z��C�.��Z����r;���ș�	����F����1��6ӣ��g���E��pf7+�2�.��S�<i��sOD�Gcn�ʣ�&�!�\�ڴ�q�6�#��z�Lj=U�K��џ��d��VƷ+
���T��uۂG�q�,e5�`��3�������9�k@k�֬G*b�2t�t�:O<�S��\B9�Cka�P�:Dv
<j��x�E�^��I��D�q�3n�KBK�M7PM� ���]R<vL��u9m������0nǀuuH�	�2���,�{I�Һv�BhV���#�5we���X���	��9B-�V[Z�������, �v<�[z��O,U�V�ۡ��m�.� �lxWVǀݏ ���wWn��W�V7�ݶ$��k�M��
��fQ��t`�P�ٚ�jm+)��+`�6:-����x��� >ݏ��:�z��.NO�M�7m�][v�ʪ��\�8�^�xV� �v<�H�<?
�جJ�cv�� �x˻/ >ݏ �ml�v��W-�I�.�M������c�;�[/ԗd��;�׸ն�؝�7Wm� }����x��x˻/ �*��Sǽ47�\�$�Eؐ�hإvF3������m�����ڷ�j�:���_����7b2����������v_k�v[{Z�
E�r�i[� �v���� }�<��%縑�Uʵ^�]��O5���ܓ��}��Nw��r�#��N�ʬ��U|��ݵ�x�r,���[�$���ۼ �v<��%�m�X��*��x�.z�~�n�C����%��U��Wc�_�g� >ݏ�}���{�D.Sh���.$S�<n��Lg�ԛ�P5��3�k��vGU����M���m�XWv^ }��ڒ�	�+iZ�wv��˦&�ջ/?r���M��^�ݗ�����7c�q�mS�;(n��x�<���/ �n��:�e����\�m��Э���]��� ;'�ջ/�s�ʯ��נo������=�k���Ս�hn������ �v<����?���omc4h�Gg��n4F��Y�J�H�aمB3vB9`��3i�e6�unĭ���/ >ݏ �mI~�*�v��{��%x?~ĭ'`�.:-���c�;�R^�ݗ�un��>�U���m1�C��{ke�-�xz��׀�� �B��O��J�m�� �n��:�e�۱��R^�+������c��I��:�e�۱�ܽ�nI�����"�j���"A���g!A���p�P����ad!1dP�;�i� B2%�~ �H��FR6�":4��"�Ċ$a�آ@�`1�H��ʦF	!	$$!#aF@�H@#$�ү┒A�s�qCI�<B��`r�V��	�#D����h�Hy��"b�������"H��g�T�w��Dbu��8�o�1�&+BI@��D�e4���lDB	�!:.�4���Xh~~��0��<	��H�D�K0r�H�H`�Ɯa���iJ�P`$Q\����f���h�IN�l�DJ��*�*U�Zeo�W8*�*E`&E�*��g^j�v�1�T䖮��Ӝ�bVB�Īy&���m\.qd����z�..Qi�����V���yv��Jco"�Hu]]U��S��:���`cg���{0�MٙҌn��k��nԺ�Vx�t�Np=�q�q,!�r�	�$t7,2����j�*�mh��R��[j(���6h�l�`�;��w�m��p�l7����W�e6���e�YiݬT�3�i(Xsт�<���K�s��/U1i�a^X�C�ɕW�uiK���Eóg��*�ӆ�S.���5�h�\O;ex}nz�;P��k=Nݎ�Z�v69Wsdq�
uԜTE8n��ˀ�mR� ~}}P
�1Xeuے ~~�_eݜ�G�;p]�&�糣h3·<� ր���g�)�-sc��v��ڜ�HǞy�&��:떫nTT�'  �F:���<�ɍ�:�+  h�g�[��-���,Ye���L����	����[�,u��)�T�26���F��#��T�dr�Z�
�<ím���ўm��\���u��#j��L��BSnvٹT�rL�U+d���eݴ'lFHʆn4J�t�i��[l�{��d԰���Q���i�E��H���m�6���e�9��-�dLඞ�'[</n����	���{Wf�L]s����&��:Dn�8^��\]�91Rn3<Z�CT�E����9z��v��F�W
[gm�岚1)H�C��ښ��x�3�=�s-�P]t����B��u���UF�nI�j��8��F ��wa�yv �4��S���Y�<���r���<��n�u��sfV���#iV���-���K&�e�84��6���%�/m���V�`���54L�RnLU��eq��x�������jU�n����v�F��e55d34D^)��_�D8� ?$ � ��6�<#'�u3��v���f�ڥ�?a�b�WW�r��<�x�cA6�5�68�6˥#u[/lw@bK�#j�؛M�j��l5/!;g/Y�h�MakGU��cH	r��'jrR�;T��v��֍����.Fݮ�� ʹ̇W[d��@X�,Wnq�M��vL�;�Y�;�/��ާ�.a��q�<#wf�m�C��dZg&���S����sɃ�2*���/�u'G]I��I�ǀ(2�y ���Rd�d�u���G�t�q�Ԛ���(����_<�ss�u��fW~ ����}�Ix�v^ջ/ �%���tݔ�m�m�^�ݗ�un���c��s���ډ�$�J�9v�����'� �n���c�7��^%^բY`����B���� �v<{ke�m�XդNUؓ�U�㡷x��x��SZ�����|�e�/��qw�Ֆl�
\���I���G�9;l�ts���	LǶ�Q&5�n���c`���{ke�m�X˻/ >ݏ ��W��+-4YM�n���,|ৢ>���@
�4A�p�ٷ��G�w��^�+����C�.��X˻/ >ݏ �ml�� ��NZ��b|-��w�nǀw��^ }��og� ����C[e$�[x{ke���X�v^ }� I.�]�nմ+�4�&諹R�Ҷ�R����r��d�������aa#1V��X��`�+w�w��`.� ��?W�7mO^�Uʴz�lj�wwv��ݗ��9U�s�w�x�S׀w�ឝ'u����_�L����
� ?����$��_����T!� �!�>Z�r����0]���.v�6��C`�{jK�:�����x�dx�p�lJ�貛i��:�e�ۓ��g���/ ��$GWu|cՆuH=c��*PK,V��ٶ��uh��e.�A�,�wm��o=�v��bX�%��{[ND�,K�}��r%�bX�w]��r%�bX��G�]���g��]�O�Jt�Jt�������bX�'~���iȖ%�b}�w�iȖ%�b}��iȖ%�bw;����e������^�z���{6��bX�'��]�"X�%��w�ͧ"X�%�}�kiȖ%�b}��y��i�ɐu�����N��N�	4N��ͧ"X�%�����iȖ%�b_�w��r%�`~SH"D �D�����y�؟��߳iȖt�Jt���?c�!����å�bX�g{��r%�bX�������bX�'~���iȖ%�b~ϻ��r%:S�:}��xm���`[u>����Ѣ�6/]�w /�Ca�Z�؎��]��2d�a�&��kiȖ%�b_�w��r%�bX��}�ND�,K�}�fӑ,KĽ���ӑ,K���5Y,�I�k[ND�,K���i�(ș��=���r%�bX����6��bX�%���[ND�,K����T�5�[��O�Jt�Jt����y�"X�%��>�iȖ?��C"dK�����"X�%�����6��bX�'����,�a5qі�Y��Kı?g��m9ı,K������bX�'�j�ٴ�Kı?g{��r%�bS��Y����<,�w�>)ҝ,K������bX�'�j�ٴ�Kı>��ٴ�Kı?g��m9ı,J ��=��-�k)�f�ur�`��c!�,{n4�츧X�ۮdy��44C���m��ݍ���>W9wP�լ�ń�)E{qְ�0`Wb%2�+�e�tOe��=��ǃ۵�Y�c�#sG�(f��zܱ��v�OGO5pV�XY��nؙ�-����ūE��fr)s�\��@�vpX�m�N4Ҽ�4����@x��QW�C��]������ΒIzBN��"Lۜ:�ZaL�WW���Xg��Y�x���h\�;�;��Bݙ[��ir���ҝ)ҝ?�j��6��bX�'��}�ND�,K�}�fӑ,KĿ�����Kı;�{/��ř�E����å:S�:}����Kı?g��m9ı,K��{[ND�,K�{��r'���2t�O��?���ͦ�!����å:X�'��fӑ,KĿ�����Kı?wS�ͧ"X�%����ӑ,Jt�O�����L���Ο��bX�������bX�'�=��r%�bX�g��m9İ?������i��t�Jt���ݿ�HЦA��O�Kı?wS�ͧ"X�%��}�fӑ,K��;�fӑ,KĿ�����Jt�Jt��O��u�M���΅��Jݘ�nK���Jh��b^p�2�p0]pʀG%+6&Qw�>)ҝ)�����Ο"X�%��w�ͧ"X�%�w��ӑ,K���O{6��bX�'�����%Ԛ�td���r%�bX�g{��r�Awq,K����r%�bX�}��fӑ,K����ӑ,e:S����k7���g�̮�å8�,K������bX�'��{ٴ�K�a�2's��ͧ"X�%�����iå:S�:{����5�RR��"X�%�����m9ı,O���6��bX�'��}�ND�,K�������N��N����7��g�aZ.�9ı,O��}v��bX�'��}�ND�,K����ӑ,K������t�t�Jt�Oz_5?cj�WXΛ=�Y��e,�����m��9��Gh���W!�9��0�,�H�m��t�t�Jt�O���6��bX�%�����"X�%���O{6��L�bX���v��bX�3���y�u*h[��w�>)ҝ)�����ӑ,K������ND�,K��]�"X�%��}�fӑ,K�����g�ե�5&�Z�r%�bX�����iȖ%�b}�w�iȖ=��l�6�o���F������:D:'�;�{�ٴ�Kı/��kiȖ%�b~�C��5�WT�3!��ֳiȖ%�b}�w�iȖ%�b}�wٴ�Kı/~����K��&D����ٴ�Kı>�t��ԙ�Z�t��u���Kı>��ٴ�Kı/~����Kı?wS�ͧ"X�%����ND�,K��例�d���+r��.��;�qd�8�VX�gv�d�z%�Q멆cY���T�fWy��ŉbX��{��r%�bX����fӑ,K���{���U��dK��{���O�Jt�Jt�~����Xe!u�Z�ӑ,K���O{6�����,O����iȖ%�bw=���r%�bX���m9ı,O�:o=��\֦CZ%՚�m9ı,O�{�6��bX�'���6��`ؖ%���[ND�,K�u=��r%�bX���.]j�5nkFӑ,K?�����iȖ%�b^����r%�bX����fӑ,K� ~�~ r&��|m9ĳ�:~�O|v�:2�f��Ο��D�/�w��r%�bX����fӑ,K�����iȖ%�b~��ٴ�K�)��?����_�fԏ��<�5֗-B�]p���`m4�9�2nx�.�]q~��}?y�����ֵ��ı,O�����r%�bX���p�r%�bX����m9ı,K߻�m9ı,Oݓ�g����a0̆kS5�ND�,K���ND�,K�}�fӑ,KĽ���ӑ,K����}�ND�,K�C�;=.���S2kZ6��bX�'���ͧ"X�%�w��ӑ,K������ND�,K��ND�,K�tze=�)�f�	���m9ı,K��{[ND�,K�ڞ�m9ı,O��m9İ?�Y�;���6��bX�'}��[w��RR��å:S�:}O�ͧ"X�%�����"X�%��}�fӑ,KĿ�����Kı*���~ܖb��V���a��lf�Oh8��ϱ�^^KQ%rs$ �g9n�І-��;X%��5�vzN9e�b�V�v1k�n��`9�h�eײ��t��g��Ɏ��k��s�!���U��	ch�	d�Fjr\&�IPl��s���d�4��ܤ(�H�F�b�ڰ�)"��7]�=���6>�a����!>�{%�b��V^��VXf�S.0C_���%�O�_����ak�n�t�YC���`u5��K�nR�Z*R(���m3�E�՚�u=ı,O��ND�,K����r%�bX�������"X�'����ͧ"X�%���k�?�d�sV�Z�5�iȖ%�b}���ND�,K����ӑ,K���O{6��bX�'�w�6��bX�'݇w�L�5Mhц��m9ı,K��{[ND�,K�u=��r%�bX�}�p�r%�bX�}�siȖ%�b~p�z��Z�[,�I�ֶ��bX�'�=��r%�bX�w���Kı>���ӑ,KĿ��kiȖ%�b}�������Xa����ֳiȖ%�b}���ӑ,K����6��bX�%��{[ND�,K�u=��r%�bX��K;��uJk.�z�-�c=#9�<Ղ]hV�fiUa2�k���*�3 jan�J�i�����'�ﴛ�H$���[D$|w�M��K�����ӑ,K����{FW0֡3F�5��Kı/��m9�p
�@(! (��@+Ǒ?D�;�S�ͧ"X�%�߽�ND�,K�__:|:S�:S����/�tVj�.��Z�r%�bX����fӑ,K���}�iȖ%�b}�w�iȖ%�b_�w��r%�bX�|t���Յ��]Y�fӑ,K���}�iȖ%�b}�w�iȖ%�b_�w��r%�`ȟ{s��6��bX�'���ڙs.j�$֌ִm9ı,K�{�m9ı,K�}�m9ı,O����iȖ%�b}�{�ӑ,K���v{V�s\w����˹fy%�l�9{MeK�MЌ�L\��f�Ҵ�����3�Ο�JqbX������r%�bX���_fӑ,K��}�ND�,K���6��gJt�O���i?Dˬ��2�t�t�%�����m9ı,N����Kı;��iȖ%�b_w��ӑ,�N����~<�Xd��̭w�>,K��}�ND�,K���6��c@�v t�qE"~P<P`�P���dQ�D��C&(����D�?	�S�I0� ���j�P �E����B
Oh	�P(��@_��&�	����0"1�% �U6$]�
��|��G@�Y�&�xlpsQ�6hO�� P�nCg�)�|~F18��r�	D��'\��j	�^8�� �À.��ʿ�b�AJ$d��"��J:���@ځ� ��<X�5r����CS�,1:`�@o��	$ t�Ȅ��QC��ʊ��
T�o�8�`k�����+@O�I;�1��ڪ'����D��}�ӑ,K��u���r%�bX��'�z{ZˣReц�kFӑ,K?�D�����r%�bX�����[ND�,K�u=��r%�`(�ȟ���ߍ�"X�%:~�����fݲ6�]�O�Jt�K������bX�'��{ٴ�Kı=�{�ӑ,K��;�fӑ,K^��_~��Y��5B�d[6"x9�"x�����xݕ�P8��!m���
ޙ
ĺ���m9ı,O����iȖ%�b{���"X�%��w�͇�O�2%�b_�kiȖ%�bw���?�0���4K�5��r%�bX�{���Kı>��ٴ�Kı/{�kiȖ%�b~�ND�,K�5�{F��`Y��t�t�Jt�O��o:r%�bX������Kı?wS�ͧ"X�%����6��bX�'�d�}���֚
�:|:S�:S����ωȖ%�b~�ND�,K���m9İ?��A���*X� O�.�D'����?���siȖ%�b|翬<�ֵ0�Z�u�m9ı,N����ӑ,K��}�ND�,K��}�ND�,K������bX�'������%��fiŋd-)�g��.��jwFt�"únw3I�3=Ō�A`.�X��O�Jt�Jq���6��bX�'���6��bX�%�}�m9ı,N����ӑ,KΟ�>�Oߚےњ&Y�O�Jt�K��}�NC�U�DȖ%�������bX�'����[ND�,K���m9�)ҝ=��ſ�\M�����:|:X�%�~����"X�%������r%�bX���iȖ%�b}��i��t�Jt���5��GV�B�r����%����v�kiȖ%�b{���6��bX�'���6��bX�%������ҝ)ҝ>����~	�ғ0MW[ND�,K���m9ı,O���m9ı,K���m9ı,N����ӑ,K�؃�E�{���̴jf��^Jq���3��a�@r���c2�J�L+z�䝛��]��c�J�/�2My1�s�6nv�uʹ�w4�ia�۲Y��RzA&�b�	d�(ڬv��%�9���@+X�@Ļ]�[����@��b���Pu5��F�u�nQQ;rn1���k=��v��	�Z����9<��n�W�"�%O[6�yiV�
��.�����]f�Ym֜�h<
��]��Y��k���-�8�Cv:z9�*�ZU�lp�����+*�ZK�ALi�AfV}�,K��>��m9ı,K���m9ı,N����ӑ,K��}����N��N�g����m��uq���r%�bX��{��r%�bX�ϯ���"X�%����6��bX�'���6���!�2%��;���ֳn�2�Z�r%�bX�����m9ı,Ow���K�!�2's��ͧ"X�%������"X�%���zo���[�[�)��ֵ��Kı=�{�ӑ,K��;�fӑ,Kľｭ�"X�%������r%�bX��}I��e�Kf�53Z6��bX�'���6��bX�%�}�m9ı,N����ӑ,K��}�ND�,K���뢙5��zwNp�H�DYU�ZK���l�`4�ne�
��eF���P�fWy���ı,K����r%�bX�ϯ���"X�%����6��bX�'���6��N��N�޿��~Ntc�V�/�>,K��}}�m9��,�CȪ_m��KZ�8m9ı,N���r%�bX������Kı>��w'�0ն�4ML�ֶ��bX�'��p�r%�bX�g{��r%�bX������Kı;�_{[ND�,K��<YMiԚ�5�ND�,K���[ND�,K��{6��bX�'s��kiȖ%�bw���"X�%���;�d̹p���Lf���r%�bX��{ٴ�Kı;�_{[ND�,K���m9ı,O���m9ı,O����>��4�M@��F��5�;-��(2���Zgڵ�lZ��|��w1;�u�O�,K��v�kiȖ%�bw���"X�%��w�ͧ"X�%�����ND�,K�d��u�)�Y%5��ֶ��bX�'��p�r%�bX�g{��r%�bX��{ٴ�Kı;�_{[ND�,K���Me�Kf�u�Ѵ�Kı>��ٴ�Kı=���iȖ1B��(#B*��<(�(�|(��9����[ND�,K���p�r%�bX��D���3.f�5��5���Kı=���iȖ%�b}�^�[ND�,K���m9ı,O��}�ND�,K���]�D�Aĵ���å:S�:}�}�kiȖ%�a��������Kı>���v��bX�%�{�m9ı,K���l��4�r��e���Ńmc�Vx�4���5[�2�8K3Y�3Bh�v�:�L�k[ND�,K���ND�,K�u�]�"X�%�{��[ND�,K����m9ı,N�k��e4�P�Yu�ND�,K�u�]�"X�%�{��[ND�,K����m9ı,O���m9ı,KӲwڙ�3	��F.�v��bX�%�{�m9ı,O��絴�Kı?{���Kı?w]��r%�bX�=��9�&��u����ӑ,K��>�����bX�'�{�6��bX�'﻿M�"X��r"�����[ND�)ҝ=��O��hі�5_:|:S��b~���iȖ%�b~�]��r%�bX��ﵴ�Kı>ϯ}��"X�t�O����)���nA��1׮��JlWgbݙpY��! M8J��6e�&�j���l�f�q?D�,K����iȖ%�b^���ӑ,K��>�����bX�'�{�6��bX�'�辰��m��&�Vf�v��bX�%�{�m9ı,O���kiȖ%�b{�{�ӑ,K������O�r�D�>�����-eRZ�WΟ��N�������ӑ,K�����"X�%���w�iȖ%�b_w��ӑ,K���i�C,�]YӢeֵ��Kı=���iȖ%�b~�]��r%�bX��ﵴ�Kı>ϯ}��"X�%�ߣ���oe8���t�t�Jt�O�}v��bX�%�{�m9ı,O���kiȖ%�b{�{�ӑ,K��?I>�	?
����m��n�8M���/gq��l\g56�k+p�M� ��@HҝY�+�\ةw~/���\l����;u�v�l.��\�Q��6�p��v�΂)�r9v����f96���i��d���-�$�pC��]�ΰ�G�"z���Et��u�����ӧqC���eP]ì������P;6��6�d�l�r�g�#ʧg�
��.7��P�Њ@R?e��V�2�ջ�z�1u�I����]�˧��x�Q�U���b%ƈ9�j���t�)ҝ)���kiȖ%�b}�^�[ND�,K�{�6��bX�'��]�"X�%���3��lf��F��å:S�:}�o}��"X�%���ND�,K���ӑ,Kľ�}��"X�%�����O��ն��._:|:S�:S���ND�,K�u�]�"X�%�}��[ND�,K����m9ı,O���~����,�å:S�8��w�iȖ%�b_w��ӑ,K��>�{[ND�,K�{�6��bX�u?y|b|�cB�)�S��^�z�K����r%�bX�g��kiȖ%�b{�{�ӑ,K���w�iȖ%�N��t�~'���ڠ�Hf�Â��!�Ƃ�P�B��:gP�]=��a�Z�v�k��c���kU����N��N��o��O�Kı=���iȖ%�b~�w��	�&D�,K��kiȖ%�bt���2ۚ���D˭kiȖ%�b{�{�Ӑ������DJ�b��pD�@��`/D������iȖ%�b_�{��r%�bX�g׾�ӑ,K��ƼCƌ��kQ�S5�ND�,K��ߦӑ,Kľ�}��"X�%��}{�m9ı,O}�p�r%�bX����&f[&j�&.�v��bX�%�{�m9ı,O���kiȖ%�b{�{�ӑ,K������Kı>}��3WSR�kSW5��"X�%��}{�m9ı,O}�p�r%�bX���}v��bX�%�{�m9ı,K��Ը{Y[9^m<ݔ���v6�H������w�gn�ۆ�̛]��!HڹݓsU�å8�,O}�z�9ı,O�k��ND�,K������bX�'��ﵴ�Kı=�S�%��!sS)���]�"X�%���w�iȖ%�b_w��ӑ,K��>�����bX�'�׽v��^�z��~�0���	�=e.S��/Rı,K����r%�bX�g׾�ӑ,pP����DH _ �v~��'?k��ND�,K��]�"X�%����K��֬�j���Z�r%�bX�g��kiȖ%�b{�{�iȖ%�b~���Kı/��kiȖ%�b{�vx�[sZ�a�tL�ֶ��bX�'�׽v��bX�'��]�"X�%�}��[ND�,K�����r%�bX��*�����-�	c�;h�:x�fh�u�+-le��-��](X����5�.2��d1�kxɪߝ?�X�%��u���Kı/��kiȖ%�b}�w=��"X�%���]�å:S�:{�{��mvѥ�i���9ı,K����r%�bX�g��kiȖ%�b{�{�iȖ%�b~���Kı>s޾�jkWRW55sZ�r%�bX�g��kiȖ%�b{�{�iȖ%�b~���Kı/��ki��N��N��g�R~�����1Wy�"X� �"w��iȖ%�b}�]�"X�%�}��[ND�,
��P���Z�M�߳iȖ%�)��}�����+f�s|���N�%���{�iȖ%�b{��6��bX�'�}�fӑ,K�����ӑ,Jt�O�߿��\��-(Ź+��b���I�G<�w��:��gr>��]xL�H�U���j�֯�Kı?���m9ı,O���ͧ"X�%���]�"X�%���{�iȖ%�b~��FY.j榳[ND�,K�>�i�	��,O�����9ı,O�����Kı=���ND�,K���2�sY�:f���r%�bX��^��r%�bX��׽v��bX�'��siȖ%�b|g��m9ı,O�x��m3H�MV���ҝ)���c��w��v��bX�'���ͧ"X�%��wٴ�Kı=����Kı>?�~m��i��Ο��N�����6��bX��5�fĐI����M�$����A$O�TU��TU��D�Dj ���(����"
���"
����� ��TDF@	 ��E_�QE_�D|�**�AQW� ���肢���
���**�� ���(���������AQW�&(+$�k4
�{� ������+Ϩiր>���u�����[� � 
 I*�$(7π 8 Y��J�w��wc�� ��yX�w9nBR�Zt:S����@=�w��*�)�{�Au�4R�c@wP����&�E�+��N���r�@��+��n�)�qJ�l�QZҐKf��҈@�S`�WZ)�z(R���Z�؄��Nƪ���DU*��T7/���Yb4	*T�      ��R!JTh�2 dba$&T�?MO�h�L��@�O(y$Ԡ� �&�#��h$M4)�z�P�2��z&A%I@  @�4�0��;����wI���.�� �O�����+����Ƴ0 @��"(��Fi ���uڸ{q X�ż~�~�?_��������G��V$�
RF%6B_�y����NA�p
- e6F�͕X�f�����U�I	ZƷQ��8��@��ΐŊ��',(H	���s�E4j��	HE��U�2�^�Vdd4[�`$ S�IP�[��w]�7Y�N���Hv!V��Y��Rx��ah�B&^ թ���+N͑R��4�+l �)d$r�1��s�'LJ=��1��F!"PHB�C׷��U��B���a���Ǎ��P��	CB	���( G��ab�E�D.+B��d���@��i#���!��$	a
Q!L������F�6��c
.�
$d`�R7�A�6 �.9q(Yp�O%��O�/+���I�E
2�/�t�!� X��H����kr�7��,�9V�˕|j�a)9��,��|B<0��C΃�z���8��p��0!D �����d<%����N8	�	�	���{']�Ph�2c�i�Q#B�������9Ҩ�h��%�JBD�)�-����U��ޓ� �RE��#RJe2�0�k<9�8�%{���^���#�C���$��o�z�	L�/%�y4�HA6n��Nz��D�k8�LN�1�����J�Fsq�pB0���c�0��/�f̚_%��y�t�ԅ����7���H�#xl��G�x/(��!��M®d��D�$��C�#�FL2��2���G��A�H��H�2'@;ϗ�|Y�,��d۶9)Iw����^��Ѩ}������q�����:,z18�F	A�PJcL��q��^�ڝ�gz���D땱J݌��Ur����0��B�q�FD�	�+�p��َX�g�����|��Y�[~�{�#�d"FXFC�@�	H�Ж3�D�Q����I��#/�]����,�%���2�!o9�I.�a��Ą������\sg���=~\E��P���4%�����'x���Z�(CPa:��N�1��UP�(3b��-LȐ��w��K,����{l'-��bvC�,���g�Q�5)��>7�φyi}L�9!�2���א�w�#׏��Gl&D\��[�P���谉5<*�A��"±=S����;��㥬����MZ�bLZ�"WK������6w��������Bo@�M(0���M.	�����e��5D��S&���X2��
S�SQ#��|D>��.���{����ލ�0c���.L��X]]��؈�����UUUUUUB�]W]�e6P 0����*�Uv��ƷC#´�ck�ث/�i`�@!��ڻa�ٔ2@@͇��p(f���@!@L�AUT�&�5urڬ�E�@V*��-,��v�Sd@X�h1Uو���������q�͍�����X�C+" ��(m�3��6l@P ګj�� �1AUV.�ښ�!,�mlmTЫ��
�����n�m�]DHj�º��r�Zc0���l��:�R��dC���5�+u��Ne���.z�Uv�P�l��ܝI+�^%�Y[ٚnn�ڠ�V�u%*�1��\���͓ �@Mjm�C5P �P��mv�����ڽ�z��)P�Eŀ���V�Pt�L����l�ۖ�y�T5!��@T;`���� .�Wl���������
���krͲ�P�m�I�EX�QE�l���H ��U�Z�[Cg\0R���42�Ha��"�ڻ[��Q�{����R�2lJ���Y��ll�� �U[l7"��@��Ŭ�ڪj�̣H]F *���0��e %���cu�r
� �]��t�l����!G"3eUP��n�l���*����U�^1�mnUUx��#�ʻgc,��*������ ��m� �ڪ�������k6�QE��C 5�Z̪� 1h`�UX���*��j3a���cS<��M���T3�U\f5�B׀.�0L��в��L�Ƭ7�iT\J�Z TG	L�.�knXF�;F����ڢV�[r��+�У��UUU��6P,T]UUPvv�Ri�nqh���l �����ɴ�j�7EMkb�FU�Q�P
�b�����j�m��QK���^�6ʲ^P�h3[m�K���w���0[%m�l�B]�ˆ!	�]�V�v-Ϊ+��B�+p `v�UΥڹ�4��$��(��DX�V���ͮ�Vյ�L�-��UUUV��&-�*J
��������UUU�*ŵUUUUvͪ �fҬ�ƙ�u꫶�q�4�Sl�
�\�Ʈ7��P-1l+�UT���m���,��UUh[��qu9]��\��]n��Ԇ�iJ�,�ۦin\���UM�ZƗ�(f���2-��춑���mش�*W;( �j�6˜��q���T�
�1GL�nM��V	`���%�e.��WM�
�U���5Q�Cl�����lT��m]���f��3@V�[t�13�F6��R�Y���
4kj�h�M�U�mUTU��� 1����P	��@���UT2������e� @UUUUUP2�v�"���IvV댮��D�؆ɐ�5�ST�]V��3L��X����UUUU �3�33.�2;��Ԑ ��S		��Zـ�`�6DRs$OBG�f��	�'pQwɽoKzb.�;@'HeXP�6;!5��^�#�ҋ_:��C�b�E"v��z^��ƃq�')�20`C���D��!�C�{�h-U��FA}x(������<������A��"h/���mz�y;�SG��@�{S�gߏ�:�9��-�� x:"���x��2BP�B	N��x��(����H$tp�<ttg0�mCa[P�Rm`m�H$�
�4X��O(h!t������B��4�M�:��M��f����<aш�����19�B!�"?��P @��
�
��"� ����S��&w��e�QG0�vNj�J�m�lCdSdPj��B�)lŎJ)����MxE�ec�g-���3Y�i�+�X��W*���i�i��X&vC���eʮR���*)�m���C+.ήf�5mU�m�Rm�ɑ0�<�6J�0\�u&�u��jGS ��֔�l��L�5�n0�[Č��E�n2,4r���V�#�k�DE@k��Ř�W
�[���ԉPΨk+�JL�,S��I��ݡ���lZڭ�ep5��#@���<kjmUwxK�nP8�H�D�"������ґ�joRV�d%eu�Tl��{a�ź.B�-�h(`X���6�[�Ѯq��ҫ�����
�\U�Ԓ|I<�z��R��Q�T�([_���*�5�'9Y�1ަ�f�P�]9��<������$�}�_���"�]4�m�5�Թ{[�ϽS.�"�<4�����D�����WS6�Mw'9Y��L��^V��%ZL�!�i�}_�������,N��n�<@A Ga��<�%�f)��A�|o߿K�]��+Lݙ2�K̬{�]�E�CʯM���V��J��cW��"�RI�y�M_6��5�Bb��I�'{�z_��2ڷJ��4̙y�DD@�Q��� �^���� � 󔃨������ysT�ȃ���׵W��C�����|NsuZA�iQ�'<�rN{�>�M��ﺋ�):�]t"�q�-��ip0ZUQ��Ům���qF&�ʛ�ݒآ�3���mA܍�6Sgd��rS9�9'>�I���,��ք��y�1�M�Ni�МqdD�e�]�󔃚�D�l�O�4�z�y}w�A�l���� � 󔃽����ԙ�a���i��"��Iϗ�s�ܓ�>X�$��T&�nv��hM���Э�D��S��
� � �`����ܕ�z�u}w�A�7|�Wh<�:�<� �t��=�fi���~ޓ�'Y���qnZţ��%ea�2���� ���fv{3H=� � � �t�z�W��A��$]�0��}�	��	�sί|f���R{H;�7��U�H<� �'=���^I���n��q.�	��ʓ�Y35+H=� � � �t����e]��/�7{�A�)8{�fi��{�A�A��\�ڏ9H9�A�P��R��A�n{3H=� �� �t����$�3.��d�2�ea�,���A�A�A�){��˼�`��H=� � ��ڬ�A�)5H<�;�=�9���{H:�=���H>��+*��Q���'<��>�I&��LJ�GV�:]���ib�Q[��n��j�c2kZ�k[[�@)��j5����`]v޺t�	$�_.����R�R#0�y��y�A�A����r�sT�ȃ������� �����������/)�"9H;�;~����v�����F]�	���%�q/2k<��fڍ�2@��A����q9T3.��z�؜��ʧ2^W�����KV��:���W����ݻ�M��n����z��CJ%/㠅� a

0@�	`�E� �#	 �"B2B"�+���7I^(�'&/�0���̑7�qg\�[Q"]�9fiu���A2��*Bv��+[������'�|�(��� �u	<��99�s�����L�iIE�����zQW�E]�{�W{�sg��f�U�UAU3T���B�MP'E ��gZ��$��a9��HoI$�j�m���9������r���r�7گ�/4Ƽ���r{��ߟ�zh+e�ιոȫ2�j[�s��:kv^m��Y��w��!ْ<�6�m����z�؛�7$������0��15%܊�eh\˛e�q�fh�ʄ8���ţ�,(�kjͰ9����t��y�.6�Yf��e5�$&\O}�S�f`�_���*�j#�/+3��߽�/����'2��%���VP�	��_�3����j�%�wd����#��l8�~d�ݘ�wﱽ�e�o�� {�*�A����݁�r߄����ٽ]+��������t��vͿ{&^٪�b���f�d|4| �@�`���Z��}�'�$��u8��>|�������9� ��,v�����c�&װ?�'w��.�f��{���s5c���[�
$�p�����w�lwd� N}r�4�a�S1*%5�C-ľ��/��j,n�l�ٞ��7�^ɾ �#�w {��ߢwt���znl���X��	��/L�50�Hm�ˊ�,мg��wK{�4t&�6�P��UB���؃,YK����ˑ�ec�V%V,��ϳ��M�>K���i��2͊�Y�ޯ���~�fC�W?�{`ݒ.�� ��dˢ6�`#���}���j�w��C� 8@ Ox-�Q݄[v�j��<�9�9R&Rm)�[j'l�/v@"�߽��"UD��%�f����7��r����뭢 ���|ݒ�I ��]��`$:ٴ����V����b%�L9
S��*��_7ݤ]��Ľ߇Vv?|���r �@�J�����N I={��۾����~|�O�����A�h��g�f����{UBG��e�TU(�;�w>�̽o2H 8,�G{b^���h���Rm+)�A�U��>?>��=��χ5=����%߾��&�����5?�}c.��|��eW�����AT��D�0D�#D*;��s�`���'C���;�D�\���D�#�ܝ8�w�>c:�(��*#eVGF��,`FE�!	�Bh��B2@K��Ȑ��B�XBB��;$
O��`B�&�<@�d~.]�H$G��q��b)������E+
	0-�QK��vͻWs�,�Ѻ�sj�T�p��;h,HKE� 텙R툎t��mZ����ݨ[m��m���;�� 
�mpl��6{zW�Ji���ƗJ�]�:ck��n[V�J10�l�#6M�Sf�����;P�����cd ��!�p�^]v��e��]���+
f�V+�u���l���0ª�Pu�A�-�Y�X���.U���evT˶hch�MM���mh�3ʆ���)Eج�A�qrj� ��\j�b� '��؄����:;��c�lIN1!'*б�<8���`P�y���m��2X�-i`��6��l�yq�&���q�܅t���\괋M^5���ݽ:�0��Or|wyM��.t-��J�s
e˷����\���$���VO��̧���Y��u�W��1�c�˸�:�D�gk�n08W�{��x~�~<>|��{��v�tM�7�[�qV�6�<��~��}�����:h�e٢���Խ{2�m���8�{wh&��O�>��v��  }��}�����뺲}����}���OIL�e��ʕ�H��{��P�z|�z�n�߽�/[ݮ�~r�-�� �d���Tv<���E��r�R%�2�Q1��r�*�����̨�Ns%�U	���VUC���v�@	 @Iַ&�8_�4Rs1*���b�Z�#շj�e�.M�Z�h	\@�L����Į�ˣ�n��Nqi�Ҫ�lfs
;A�~����}���
�f=wӕ���fUMo[y�J�o�e�JF͔�\GAO}|�y�|��߉��d�Z�y���ws�\���+|>�}{�|�}�g�W9�&�3 �$(mFcʮ��Ng<E��������#@x@ xj=9�s���T'W�̬��W��Xx[a�5�B��+�}�����e抭۫��/2��o�m(��[�@�( d`=�{}����w���ø ��,6��8�����>s�������[l���y����#�"�G�np�׻�����U�q ��G��4ND�D�r7k�;�6��Ȅ�Ҭq@���V%�A�)Mu5u�	R��PX�bW� � �jQ%�\Wl�?�p�z���i���,�Q��u�g�sS��̪������h����s�����g���J��6�i�-��M���$]�Z�y���Fd�,�ET�X�e�ЈqC��kAϾ�/[�H# ������@��y��s��j7t�Mm�ۈ�0�9R&Bm(s�5.�����A�w�c{�����;�}�����_7��2of$�w�A(*� ���$hB�5܆�U�Y�Z"��r�)q_&݃���GM�Q@�'CG���yy�'v��(�7�{�}��5��3	��m��{�^|���w�<O����X�[��A�����Afچw`R�n�����b��!��[�G��:�UI݁��@ H�t}�2��D��R�[������*�6��@�q��A�(����ڠWt��72��\����c��n��{#��?���Ϭ��d��0��"c���6��xM� �� J�l0�є�mղ��4��1����윜缙���1�m+)�pϱe^����;y��<ܟ��1CW��`b�wc	
�Ӎ��%��5[�,ޥ�����\�i�ٽ8�+T3|�pw`h .���=|�CQ��J]��E.U��y�>o���9�9���y�f����<"�{�j�j>���Cvdp�C�m(c0�G	�1B�;�_�yL�F�݃w�Ϳx�������=�ϖ������j�j6��+ɷv ��G�@���]���|�#hn�����-�A�����)��ܴ.H*a��0G����=����M>Y��ݑ�@�q�3��S3CQ�7`��������@�Q����l�F��u���(�Cbe��f�Q���:�}2�Q�7C��CzdZ��re��UA݁h�1^n� =��lGP�
�3��pu�1� ލϠSIL��L��\\�
�\�U�*���r�#��h"sT
`[��	�ipkB�٫��)�^nw��gP�maV��1���<<���w��rqx���^	{�c��]@�m���p<@!n��u�$� ��r�#�m�7p���m��J9B\D���j��e��UA���G�����I@8 D@�mq+�,�P��
GP��>�j���G�n����<�Τ���c;�6�r����į��z�O�w����<�?&���V����ȏy����IG7�6���[.B��G�����{6G#�Fzf5Jp�JdD)m�ˆ�@l)�P��
GP��>�j�����Cރ��>W.N!.��F~��sC������Md
�6��m����d�C6�tGҒ�������Mn!��j6���_M̶qyU�݁��C�C�n�t����2�́H�d��z�f��hn������K�p*'��B�b�KJ�{����u
52�Mp�����KK��rIs���h�� �b�bV����I��D� U�vW:�NB��V �\�.�9Թ�c����A�v-j0�ˮ.�q(*P���"�ر�l9�X)[(�9d��)W���*Z�՛�����ɍm2t� �Qԙp(�M�m�1���[�]j.B�6�	G1�l8(�kk1Twc��!��CD5����[�%�"Tj����D6�(K�-(���B�عT�L��5q@��W,[WLCR�mV�lu���]D�B�\E�����FjL�˪2��.�˪���'�A��[��|{��y�#N"�.�^B��߱H��L�m&��\l�k4З\ƈ�
�䕮�q��;��攳k`%��W��S^ގ@%qv��51)˓�73��E��c��]@�mq*�W��v#�]����t$lCvd˛���Áh�uJ�S�55fq�H�����}����,���-��f�tp�@F��'bň�>S3C��;������ �����47���{;�>S�|X�Pc,��@\kci˃���03 �������!�2�f�qPtP'b��ǭ��k j6��Y��d7P̃�`ɎmC�BQ�e!�>^ygϛ�y�|�m�q��@�gpt��݃U ����9p9w@�u�1���'	0f�O7C��7`���X����-H��
R���s-�A����m�ݏ ��G�v�́H|@Z�d�~39Cv
̀�/cl�UI݁���$�|���t(���Z���rR��P� ���1f�<V3ut%B�@X����݇k��ĩ4U��N�'9�3��z`�t��ƹ3>Ͽ�Ǻ/�rI�=B򇜸;�-B�>H+tG�7C���^F��#�jpw`b=�zۡ���	���?{>u�V�H���>ŕ��gv#�2��t�P���d@J�r���R���� �����鹡�?y��C�!x*W��݁�l���?����us�BP�!��
��m��3 e�re���
��G�����5�<0�� P �GP�����H��%�}�fhr6���+������jK.2�S�ػ��������j�j6�Xr�[9�-B�݈�n��hn�����@�ӳ-�C�sϟ4���~~�y���I��v3�*�n�����>K2�́H�q�?o�L�F��2��[ru��@�9�G�f�t����@<<7�LM�"e���
�`t�e��lfZ��1�q�L�t���Ѻ*��
J6*�`I���{N��a6&M�-�+ 9q-���!wn�{�����n�]t��gu2���[t7`�@�1b<���3���.�ͭ�9̶�!�%�3CmL�F�݃wU�[rqbHd��� `��/`b<�u��݂��hU�=�́H����w�����o�'���mt��<��������$b8����wA������ͷ�{F�֞�B7��2��MU�м$�q|����U��,[�T��-~�sDӑ����{��(i�+�ā`R!!j�T���A�;��@�E��.������ߩ�S�a�\����3Cv��1�S�-���!wn�o7CQ�7`���鹖� �d5L���r�c38�k�/��ͦug��,߼�Ve�� 1���N��gv��]���Xۡ���n���g��B���<���W�е�W�^c�Ѩ��=TCƔ��d��w���mh�V��Ά-��QFԄ�[�M� �YS.)��d�4!�����3��ݫh�]y����]HfZ[6Sh_�{7z�Ϸ�Y���,� e�c%��UÁh��z��݃Y �J�q-�s,���q�>�-��CQh|���>_����+��Xm�8s0q
ps< ���h�L�
���v�%������sv7CQ�7`���鋖�!U2�<�cSP�1"&T��Ø�r��C6dF�댧��бC2X͜����ld�A����d�Ps Z<�t\�݃�.�r8���Aژ-��a0�]�r���;y��2��n��hn����錖Π��F痮]�5�5:O��v�q�����.�� ��܈��0�%.DJ�L6�L!3*,r6����ל��)�́j�\���-��u
��[9�)CNd��#������(�#ً�t������(Er�hV��ˍf�e��jYU.]��]�7 ��n���6�`�@}���H���]��2�a,DD�&\9l�Po�Z7:�r�n�����=��ܳ���.���Ț&��6�t���`���@�`{":�D˘m�3 �
0�����{���,�/Ѱ3#�"8��9r�O7CQ�3`����-�B�dF�W\��k j6��I���Ϟ^�fP�U��paa����.���6r&���̓w
u�˧��Q�@_�	�M��z�C�b��	#}&�#�U�+ͳ��=��7>��_>[J�2�[vuJ@[����n�[鋖�/�����!�W�S���FЯ@ʘl�@�q�0`fQ�s��j-�7p���L���7���.M�l��a=��ߓ�Cv���V���dG��7cy�CQhn���u�ܸ8�T���@�0-߁8�E����|H>;`.��fv���v�c#0$#�՜�J]ɐ�EI!4���H=z�M<HB�)���t0R��i�5 >��b��]nA�2��@-����F�ˑ�u��v��\�-hIQ��B��(1Xڕ�����U�f+��-��]vUZk���[����:c&�γd���d�@�֍�	����Y�nJ�ui��L��U4�Xl����.��m�U�)v4���V�Kn��,ʹ�W�&��b�$nk��q�֕�ն� �nq�1s�#�UV���u��nq0!�����-�V��m\U\�h�,�:�n!p��1��]`&Zۨ�E���h�[�P�m�¹��bm_>��&���x���ݠ�w�|�qщ����I�N� �6�h�J��ޮ��%c(�8�[��c�M.m�h%э��s�e�;6R[h�1sŚ]{��;��k�͔I�0vp�ܻ�k r��1��r��G���b��t5�������Z���բ�f��P5C� {fl9�JA6"�d��*/>|��ϖy��ݎ�n�� p��t�^V���)��N�\��]��m
�R�́�pv�/:y~��vK�����5G=��C����s�s R:�u���g*����yt˟]�g}F��-���E���@�;�\C���2!�q��0���9�)�]r�b��5XB΁���
GP�}֣-:��!��MJ4 ��ow�Oa���;y���yI��"���V:tb2�b4��s�2s 4q
^� <��ۡ��5������9�<H7ߗ�{>^>i��l�<��UUs�؋)���kn]��h�H9a���B��Yn�k�X�ܵ�Zk�3+er�$��y���+3��*1!�E�Ϛv�P�{�FZt1X
C����9��R;�);�����!��L��l���Iϳ�n�R�e�V�st��m��CU����.\H� d4�v�b56����]��i
�R�́H������"��j�MjRo��WCU�.��Ht{�s坼��)v:�hb2�b4��s�2s 40�/Pl��	��#[����E���@����q���J�a1�0R�:��T{=�|����ߐ:�����)/-EE���@��̏�-�A9Ղ�f�#.#V~�����v�`%�9������)�<�F��j�Ml�Kg�s R5:����]��,��m���=���d'v��Z�h���
�Pb�e��eE2��KB�f1����x��L���7L����y�kzn�e�	�ĵ�X@n�|�l�K<���C�:�#����`�L��e��i���24��
GP�b�t�t1�'��<�����vc�U%ö�(����9F����w�9<#��x�4L@h��-�r�݁Hp.B��b��P�Z�Tqk���)����,�DFmц��!��x:|������́H��U�n�#j����@{T&"ːK$c���r��'��RQ�T�0�D�a
H���M�;˪s	��3��I{���hԛ�6D�f/,����Y}���ry
G2#S��]E�F��k��k�8Q� ��}ӷ��$����-�45hB��n�!z�}`���
G��\�F\A�'��:�J����;y흼�߽����̸5m����C�#U��9pqq *Gv�Pǋ�.����HW@�Kg2#�R<:�Z��C���@��(q8 �uKEM ��vv�w4J`�aȣK�ؐ��J�@��«��[��J�ZUQ��p��z�fa���䃨R7�);����u�7��'2#�R1T#y�����@��\C�*�G�z� [p�P�D�b\C�-����]����0� b�d�{� fG�;GP�~�֦�"��j�y����Z�����뙡�ˁ�����L� �ms��JE�|��o>q ��f�Ey��b��|@Y^��:�CU& Z7?/�]E�F����-��$�Bѩ��T�1f"r�jd$(M����1�q~�0qx U�����뙡�ˁ��a����|��0�C�=,�X��������yg���i��t��Q?���?�
�Ur���t
F���.�"�#HV���d
C��r���]jhr-C���mWX���o�W�qf�pe[��A�'��]���t�u�-�:�F�u�A��ꃜl�7`v�%�]���ibWm�,�35�EF�E�ڃy&�����И�B-�+rZ�A������<��s#�#�Z1v#�n�#hb5P)���s x�}�t5��#���s,�.�Ff��^{������ط��5�@�hj5�<�r��)�`Z>�깡��B���+铻�o=���9$��=��ކ�K��M ��
t�x9C�!HS���)�>A!��ܻ���Vh��xLҵB�*[;�)C�>$䟇�{TP�x�����4���1�M�Ұ"����s�s R>v=s41|B�j6�%{EJ�d���u
F�?����iC����@#Fd�y1�l��d
F'����IB�CD�Z*=��w�{y�;�uD�9�)B�����P�Z�Tq}`��d
G�������!ȑ��E�Lx@���ڤ_q66��O�i�����	! �"Bf H�摨Iy	HIHլP�	yA�du�DK�>�qCd������\��V�ZL���D6��c5]j�����6�K�Ȭ�6I���4Ҫ1]��t�,Ɏ5�K�����:�i�r��
���8��:!f]QEt�P�8�m���m@k�� 50�[Q˵��jP��*�ۍB���5+��Q�3Tъ ��3:�,�c0l�\uи�,*lW�A�* � ����]p�p��
C �T��*��@u��kS
<���e��Vl%���F���
n�m�4�� �W.Y���[33&]�]�ʀx��t��b��ʀ������S�*�V���vC3V&3iM.X �)kƠH( �T����[�[b��3D�$4�Vm�GG+M�v޻�w�%��=W���5�3,9Nd���u
F�1��F��j��
�=-�B�݁H���2�b5P1Co}�]�}ӷ�������R�]�RC�&Z��C���/��H �/Um�@�#�Q��:swz9��!���9�)B��W7C�1s������Lڌ�)�L��y�R9��h���e�ՠJp5TA ��k�̧��p� |�q-\�;���QC�hb5P<����)��r����	�mur�3
�{x:{yHm�+�Nd~��Z7a�y��!��A����,�(N�q�h�؛>A����ϗ���vϿ��E˳(�����ˆ��@�q
G�Z�SC�R��8��2q
CV�Flw�����!��L���!H x�C�ѱ�*���Ͷ6��̬p!X�۰��Evl2��D���6nni���j.d�	.0,�s�v.
�d�nƣHj5P)��˃�4s R���t5��!]�.dG����/�ӳ��g���/~���l4�Ŗb%��N!H�@�f���C��H/ J8��9Y2s R
�-����F��j�S�C�h�@�t].�pl��J��U����Oo;g~g����!H��Yjhb-x��"w��r��q����̨c���v���}!JA	��jFh=����s��_��m��G���n;�e�r�	&��7|��ߞz�?aw�r��Mc��BSjnm����r�1���v��D�Nz����x�d����D��S-8M���R:�8ʻ�m,b�V�,��r&ٕ�&"\��t��m��Ƥ�J��my�n]���!�rE�?{��￪e�v�k藙x�u+�76�O_C��ƾvm��kpA����U�>>�N�Nf�,�E�f	��[p�;��g����>/����ћ,�6�"�L��+t������s��$ �Z� $$�ٺCD�!|My�@�>bb�H LC*�#$�1I�}��:A�BB�(B�A��* 0�0D�D�	���K�rY�D$�M8J��L�m����d ��h���;��k��D��?U@�J�E�K�� �#|9ޝ������{�2�o;�%�VG� H@�8I3��Tl�lg*�b���p�r�9���f8c_7~Y[b{�9���#�n��s�z^Vc�H#���Q�Q�f�Q��]Ck1D�P���yq�&���2���6�5ئ�Kj�".���C)��-�` ��DfƜ)i�310�`&%0幗��{����X����ɰUz}��;Y������D52��ع�m��J����'߫���y �F�d��K��i�˶��X�NNn�ߦ���J��ق������~�_��Vc�7���`τ��AP;��|�}�bF���o��r��q.#�.c���}]��A�|}��Cy���R�Ssr >'I$�'�ݐϽ������]�5��c�.a_4����1��5A�y��m��=/����~��|_�|�6��Oؗ$��:�Q�[`��,E�۵L�68r��b����I���lQ�ɮu�\���D��w�r��v#�v�X�*�_�k��R�Ssm���s����n�m�	�Ǿ�����=e�\˱pWX�e�cnw��y������` �{���r�]��~q/2���WS6��(�9�9Q����[����}������x��}�9����ْ&ץ�������?>�_��V��э�EP}W�?D���í]L\�}=}|@���(�@ 2�w�����:=���Hq��		��1�'�K�k*�w��x��z�]˶�_D����@~��$�K�I$�
�>Ho�-<g��Z"~[U�y�f�U{,U �@j
�)� ���@P�Ac��)E��.���������  �4�8Ż�ojk�����/���b6�E#�^$%�6�����������H?��U�}���l��+�v��'� ���'�>G�Ķb�<��w�RT��?[�%������moE/Q��j�ŒI	j# T# aB$Ԋ��P��T" E`FJ�$����	y�(q�l՜���>k��� �^Ӛ����������M��^us����W�_��  Ō�Y�Xo_����NP��r)^yX��լ@ ��`?WA��3����m�0�KրA��g�)㟍+�j�o>'7�4�v\���@A�4��w|��@(�/q
&̹A�ܞ�[3h�S^��=?�p�
��s�����N#p���gM�GI�F�e#� $��ϴ2  -/���2�ݞ���D��0�/
z��e)KW��x���O:���� ���Xq���V�՗���y�╎��CɈl�) ��{W|�D{�  -/�z�&jk�&� ����p62G�]��BA��� 