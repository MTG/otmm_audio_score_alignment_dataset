BZh91AY&SY2l��#_�pp��b� ����aj�"
� D@(J �D �E����IQ)��������Q* ����|
%*(�@P( @   R�  (J�P	U�)" E(P@�Q@�R!*�T�� p    �   ����,f�b�Zr^���`�om+�*�ۤNl)� �V-�ˈ�CJ��N 
�VZ�)��:��=�t(0�gסN- �!�mT6�  ��
 � ���:;Jf5|��.������x�um�����'p�N�j�2�qn�n�u{���\|w����]��-� �;�c9s�^�N��e'%X �Y�ݕ�k�rp���>�PQ@JP �@ {�J�JX��rt�����N iL���g^,�i]n,'����}�/>�� ��M[�Iy� 7R�n�:x��r�N.�� >�yU� �>9�3K���8 K��J�   	���)�����{:���� L�6�)�}ŕ�ˠ�� 0����k�����N#�����1�m'&8�ɇg� ���4���\�^�]��T ( ��� �F{��>��*VM=�#� �FKw���K��7� 7���\��    -\Z]�G*� !�MRŒX̹nmI� Oz�ͽŔY�w���\��     Q􉩶�JT0��##&   ��)J��50M40�LjǪ�R      Ob�R6���0��bdb0�T�Тm��U�@� A�� �!T�F��b ��!��'���_��/�����x{{}�^�4UW����
���TUT������AUq ?ނ*���e�"�������TUU�������_������J���M�<��m��s2ʄ��آ�Bvz�4��]o����:MŮ8��\�&��1Vzy�w��f���!���F{��A)s(���-�%n�U�)gHO��wUq����yk����!լV�"mk0 �'r����λ��"����(ך��f�vh�Y��Z�Slf�p�ӳtGFiy�4��I��G4lÑ��Q�Z�3w]�uE���$�Q�*(t�]�A:�I�yh����"5B6j�jI����-J��N��f��f��Yo������@�;_��gc�D��Nk-�TK;p���Cf��@Egv��B��ܝ��q6Or㑋dzC�K�)p�b	沥�gΈ�h�.�&Y�p3���NF3�`JTY1��:<�p�7����JK3d��K��MPT&'!�yC�&�L����aK�a�NZ
���fy�ȓ�M�����2R�`�[x:�x�I��!!�g�o[S�ל�1�XFR�&��r�I���9	�tl�k\ᑙ��:�]m��a�.9dn�4ZL���(JWA0CT�d�NfYם�6�wްJl�0�d�e㐖TV!��RF8A��&!Y�<.�xF�%8�.>C����24��p:;7�:9��]DH)�G!Ew3Z��[�7�Q]�F'X^{��#���2Д%	HH�'!i�"i���BP��Y�k5&�A�KI�rr�\�,8a���w�0�"2L#1q�MZd�L�!����Zƅ]��ޛ��;�k
�h~�d$$�3�z93ʩ�T,��`��c���x#P���B�&P���D<�,J�	��v�).m���C�M�0��4˨2L'�J0F�r���y��9�#����M���$�X�a���S�8�֮5�Q8Ry���u�:��ց�B��844�p�MU�&j[��Gp�ν�c�3]�o���2$��9��dc�CY��������Y�[p�ªr���)@���J�Р̞@%)TĮAS��p�t-�N�uY�"Iv��W�U)z�h�h;�A*`�0�$���.܃&3�$�,����:My��h�2�=��S�QTFL�Bw���s���A�Mf����%�2�2%�c&A%�14[1*2�9:5b��oif�ۮ��ѽ�:�ѫxtS��<,3[�Fn)��KK���	Ѥ�B� ��Eݱä3���='�G|��|8ҕu�a������d8FG:����ug��=c�Ck:��d�# 2� 20��# �0,�C�kQ;u`��զ��(r��2d�NZ;|,ߞ����D�88i)d��ķ�]8k��$��n����hHg�V��N�#q*Q��ڡ:�d��՘9��n@���BP���E�ze�J�R�	�S�Ĝ�I��J�4�ˮF� zla8�n�P���:���5F�7�0	Y
�P�R������Q�Q��Gsvʞ�SO
P
DΡA
���!3F$��U��p#-l�&��# �a��3�!��������p(t�0�&Bfb�!����FNa�jr�¬�F�"5�ޏ�ӛ
	f�3�`��Lc��"�&��)�C3�){՛l��_xwuOI�'3	�$)�q�����L�d���fc����G�4�5���{��<�z�BV0gR䖶��a�Ȭ�A�a�ubk�X�q�����b�0N�\m�R);:D:�lE	���D�@�=뮨Bx�r�2[ys���pah&hK!��%��1U�V�Xht��/��p��.j`e��
� e��^�:Ų�Ss@��c��;C�����FRtT�T�x�n��)��ia:@�K�h,)$%�2��ԯ���@R4�`���Oe��j���F�=�c��5{g3�=�a剢f�"`1����L�{���>�'ʷ�-`��#2���*��GT:0"#��(�C�r.q܇g|�B�صj�ox%	C��۰���<w&w\�7��2�
,4����6�C���d
bDДC�Hh�+K&%0D��F%�8��Xb�<:���4�b'I�A�j�p�u�n6r`k$;�K$Ĩt�M�pR�ߙ�,���r����4h��2L(�JJ�=�5�;�g]Q��N�ɡ��� Ŝ3B3��d���R��BU���	Y2L*{�IY��<���5i�3I��X0nd�A.��Đe�j�������������w�:^h&�<�i�6�(4A�ᠵdV�A9��I�lBhRDN�C�hy��OW7��ˁk�A��r�������#�f	iq�����MNZbl�-�K�o�k�s��h��w��6�鈁'hC;
 �xv=��~�	��g?c��4�Bx�
$�����vi�TD�-Sr���Z!�9�\��&��6IO0�=���-h�b��Wb�R�֎�8�]�q�$a	�C�
�f��#C���t�����!D(O�u0�Jmb8�Ic+.������+t�b�R�rVÂ����!L�|̚#�N�3!(�h�[��G��F9f&!�ѭx�Cs��6�Ykwry��'���ᇇ��u�}h�3{�o0N�r������t�P��'���:�gK�.����6�;��k��B�4zSܹ�͵Lf����[X�j���cm
D�(�HgP�q409Pp7����h2!(Kà������ǝ���(7�WA%:]XÖ��(NC�� �q|�ʍɉ�)c1�"�[V�fr�{�gU+S��@����"r6S��.`6�'�KBV����)�)f���0`��'Pa�����4��/LY
�,q�@�	G`h#{�i
�P08��h��������k�%	RC' �I�U<3@���K��*Z&�(O�2�c��s'9����N��bE���<VY�v�nLO5�j���d�h��f�����b:�i�k30��yO��<'.�OS*��P�I��k��/R�G ���MI��P�d��݌:��5S�vD�8�;�&��=s
�a@�"A�N�Y=5�v�N���BY1��8�@�r�R�:�I"��K2X���q�O$�8nh�	@a�j*�Pk!(p�BP�КД'�(s��'Qߞ�x懸��v�s7%+H�I䆘Ckʅi���z��mk��;��1
(����U3�B�� ��b�����ڡ9��I>Ɔ2��nC)	��-�j�g9��,��l[Ѕ����owc�����y�sA�4�g�#^gw�dq4��� �:���L�	���\rk%޷���{��qFh'0�M��u��c���ɤ��f����Ն��RXDA��� �i÷dj4af	A��'Q��E��F�i��eJ-H�9�C@���O(�)�T��e�x���86��0�j���X�D���8@��ZwPf���F�3�mJ�r���8����F�TL�wt!�207nMBj5��>�/��<u�	�5eF��7&��Lٮ��:���t&�$��2q�Dg��.�0.�5�����v$�8ΐ�����@=R�p~7xu
���a����d�:~w�C�Dy9�Dn�ǻq{�t��ۺ����M�hzw�O���y�c!ţ��	A�#{�*�5�e�1&NJ윊��x�T��AN8�M���zk-���Rj�7�w�y	�x�b���9	�O-�	խ秅	�C	C�q3�::f� g%D��5cĵ��M3�%���q���!�Hz�q�.ҞR�T�H�D��5���e�K��ֱ�C	�*M�f�(J2ӳ���u(Z�~۔(�R]fړTM�Yˉ%A�d9Fa]��[15�]�:���چ�:"5d�LՕ�ҩ]��|��-	�'q���o�M]�u�Ik��#Ԝ�>��;(	BA.ҭӪ�芗{�4N*0�S��[�ÙZӆ:�]>f���<����'�z�`�@�!9���xR�+9��Zᛩ��:r�(!� 3c8��P$�d:dA9�I�T,'�%s�y�)�92��.�K��*R��j�xwQ7{7�i4�-�q�K�2��=��FLw	��f/v�:�G�rb'�a�E�FȧP)R��yivM'C\��	:ѳ[ȈH֜��vG
�tn�@�1r��ZݽyMLlM:q:}ۊ�Pώ�<JN�	�[��k;r�~�W<���ryҮ�%�'����$�L�J��[!9	�`����M��p2���ܘ��;��!;�4�M��=��y��������F�=�ƷG|�;gQ�nq{��(�x�%�N(@�u
���+"�r%�ӨhB~��}ݑ���0J����Ǚ�)R�� L�+Y��5r�	�W�L��{��Z�f�
�)4�c�12Ǉ��[��&|�:�ɑ��9�}�3:�12���*;z2�4lˌ9	���P��(YX�UB�V���&D<Zɼ�}zQC���]<0��?(Iu%:��u�����yf<Ma�KQ#���)h�]j�ܺ��bt�njJ>���&BP���@h��r�q�I�k1F�����Μ]���Ru�l��w&�'!(V	�R�Et��԰�'"rrBF���lyimju���:#r�݌1�x���e�٦���\��~Hg�&Rd�R`Z��[k�}	����OK��ٝ�:�~-���+�N��f:N�, -�K�,x%�3^7o2��wva=i�S�ڋJ-�a�%*e�ȴ��(�����������﻿?����_UUUT��T3�� ��h $   8  n�  v� ~�| m(V��`�lH Hp8$�	��Y[e���R֒�\�j:f�%M�;	L`	� >����H7m�m�lm�Ž%n�i0  @h ����۶� ��� R�����^���9PU����U`���j���f�`5�l�ͶѶ�e� �8�` �J�I��x�5@��RZ�mW�^Ln��酮^ۣ���/�U|��#��ٴ�$��"xej�y2;�8��s�UK�Ր8,u]���nQQ���0ę��k��+�2�8��Ha&��Rnܷa��$��jD��}gK$�41�H�gD� ,�:^�sN#6���Ii���Y�� ����6�v�� �e*���Uڪ�J��$�K��˶��O������,<ձ��
�US���̀怩V]�rԴ�����2eAUig2"0�T��/<qwn%ݪ�v�%�a�jP��j��-�d�Ɨ��� �Cm���6�i8��-4��m��t��Ǆc��+�U���*mVԅ�p�L v>����ڜ���W+*m��m�_N��%�tu�R�U!y
ZH���ڙ9}�(��V��۲��q®�E������nZ���}?v8M��6�gפ��	z%GrN�,��v���h2Gb�4D٥���Ql��!c�p�K��q��7Z	�1�l���=PuRmݖ��O�L�;+�+��p�R���1!4���
rP��Zy��<F�ظPǡ�F���ݴ�p ��&��Mk��	-��e�:'��r�v���^|�/'��K#R����a˰��v�ԡ=U6��U�-.\�Z�C��i��0[MT0ko�|�  -�l
�P�j�vZ��UR�]8 v��(�jQ�m���Hl��V�"�g[C�� ݶ86Sa�l�0kΜ��p	q  �k�[q��6�ֱ��m,I�l�@.�-�g�bIӰ�UR��\�`r��$   �`�h�%�y�j��=l��+M�cm���Vā�   Y����8N�ӍM���� ��F�V�U�U��`$���l.�`$�d�״��    �e�%��d���e�I�5�x6�8	���m8m�  m�6�@ 	 �v����-l� h�6�ޓ`kZ@l�p  ��ɱqr۶ݶ ��"�m�l�\�`    A��n��-� �8E�6`;m���> [@h   [@���l���d�����p 6�m����ۑ��ɫL[!%
B�Z��R2�0�`u0  �f�6� ��`���    m  m� �aԒ�l0A�hR����m�-���Ͷ .�  ��t��t�� �  ��S` $   |-�� )'l6�m�l    i"�l  �-�@ ���e� m       �( KAt�i-�Hb� � ��m��m�[@ H ^�ݍkH�6�  m�L� $��m�   �����HH��{l   I״ݒ  k[l�݅��� ��8 �� o � 6�l�    ����ڐm��lh�6�  m  �5�H� p I  ��zqm�$ �o���#�-޸ ���]���@Di��V�h�
�'"�:W. -� m"�H�[R  6�m��e�j����j������� ��`�ㅵ!m�[@&F�      &K��cN�&��kDd�5�%�T� p m��%ӳ:�����   �;i5�An��Iu]ͳl[@	��ic���I � 
P� �p�m�N�i�h� p M�e(����\�[lh���ۭ�u�H
Tk� ����$�\6� hݰ���}��o�nnͻ8l�$�i��	    ���( �?mO��  �v��6� �t�h�l   ٶH    Y�.�-��d�/���ֳJأm�kimm��+�UWD�<A��֎�Y����Sk�l%�ڷ���8Z[�� ���3k@��l�B[Ku�� �4�n�kg�j�<H�l��k�2N\�@J����V:���t���֔�(歉��Y�i�л���mZ�l$ X�m8H����͟<����p֪v���q��];s���
k�Ebڛz:r��g�K(X�����!��>��闒a�9�����xuĳ��l�cY��vd�,d]f�2<�G7.�*�����;��F;���0�ɘ�FǦζ�F�V��=��k�W��m<���+UvS���ɦ�v���>�L�a^y@��J�Uc���'�yܐ���ڻ�!���Ĝ�ٰ��ؔ�VC�,乹z�ʫqq�q���j�(v�:���z �	-'���̨~�7��ʠe�� �.K!�q'6��]u�lR��Ji^j��o��|q�6ݒm��	e��e�� �J�p��3�d�5�p�؁�Mg�� )�8MP�pMqv��Mwl��m�-�����T�':� 6�e�={v���-�HG��:�ީ��l[@��Vܐ�m�-��&�f�y{M�۰�g[v�Y,SU[@t����7 �� �i4�$BL�N�YN��th��pif6��@{[oV� ��p0�k���HX5�z� ;0T9`����nj�8)x�J�t�8��n���l�m� �a���n:��^A��z�N�v�C���n$��,�-�H����� �U`6�:m���=R��@�q�X� ��ڜ�v��!$كmm���K{U�l6�Er�p���u�*/p9�n�X`=-ki�Rtuv�������1� ����j����+*��)-O[�%:@�yM��U�;��j܊��\��t��}[�A'�^X(�7 V����s$�&�[�v�q;ƻ��/�'����f�`���㟷�+&պ�6�v�WK��NՍv���Y^�<=��e'\)H�L�;Y.��m��f����	:@��[�lܥ�  y�bޫj���6��4��k��:�v��lm��&��h-�g^l�����@�uT݀��- ��jD�m�Ά�H4�@ �ٷ��8� ���l� �a�6���V�-�/-T;dM5K�(A�l��$��'  ��n�v�h� ݰ  @��@m����l[@6�:m�%�q��M����I[7;^��#ZͶ���l�c�� -�  �K�  �n�� 6���߾���b�kn�η[�h ��m����
���J�lWT�[U(Zl-�5�v�d]6���mU�   $X�ao[��n� m  ��a�m�$m�M�   >_��ݭ�6Y(  ��;i�rIl����@��ӥq��[j�4I@kՁ�����$i:��zX���ɉX�U��P9�y���3Wg$�hZ�=�U�V�(v�d��؁�����z궐' ��{&�|ڻj������'@6�@: ^	6��d��ڬ��UPO(��Ӳ5U�e��V2!��UR��H�|�04$�V�d`��e��������[D��sn�H�����m��  [@�mHඝiK��^�xEh
��7Zċ%6 ���I�LpE��N6ͭ[�i5� �-�m��bp HK:�$�g1mh m� �-� }i�|�m����Z��{*�UAK�n�m���D���   
-��splu]J��*�p���ME���%� x���`$ ��T�ڗ��gnXm���@�]����@[Cn�p�6�
l���,�pgt���S,�*U�5��(�[gs��'8�%�*�򇧪�e�@�l��cm��ͳ��0��M��[V�
�sZ[���;i$� [Rsk۠m[3��u����Q�;5�lŅ�e�����Ievj����L�a���i�Uր*���R��Q��-��I�T� �����������j�(t��?��w�]��`]�m���B��Ŏ� ���H�V�3V	K��.��C� 	�HmG6�H"�Tܭ�M[J�mU*�	�h�`�m'm�lZ��Z�M���U]A1��%�c��������-��u�
b�0������HMu�]��6�FZ�� �b۲jK]� I: 2��KLh�ԩ��3g���9ĺ��[kN���n �jE���`^��H���k��  �y�@�w[I�t=%TMωHx�T��uvH�r�N���0���V^�6i�sfvg[�HH     [d�I�  -�@   6�l      		 � �d�-6m� 6�n�  m������g���m��8�m[�K?s��w��{���~mU_��;���������]���� �H��aG���A+�C�J�rD	{Gg �ؐ���H�*m��B))�x��:P9��8΄B&��YF`Y%Y �p��h�h=���dR%4��`����+�}v�H��v���b;'�O�g��pU�T$�A$���;x�:�����h��z&��{S�Bv����WB
��!�~(��DӠD]'�Q䁀��N�G}��j	��.�\�v�> /�=��>"�%"D��b�R���(�`  &�I:g��C��*�ҡ� �"�@� ‧�קX�8
��BH>���s��6�\E{�` 1ۚI<�ïu�|�����@j
=Ҁx�mC:@��0�����_���������"� @�0@�H�$��B�DP�@
���D�`�(JR�$)1�L�0G	q��L�ɉ R �	�&���aZV�i
Z �����ip�F�
P�R�T�D����#��{�?�|�9�ovܷ�#m�����K��4]MF�삤����c�'E�㶠�eH4���r����ط�Շ/�.�ۡ���j+v�6
�A�^��.q��7'6RQR�V�"�f�Ńj6�X��=C�_�8��H�]��mv�p<��\���D[a�[�1P��I�c���e��,\��� m�x۪��9]���]��`��v��s���x�{hN+�m^�8�ڵ��2���WR�[v��]�i�fy�n���2d�j^����ͳtc��3^�\ك  8m�&�������kM��` 	 �� ��cl��U@uUT$$i�z�P*�v�cY�!W�ؤTf��J� ��$Z� ��K*�Rl
��V�s�歀 ������GUD�SL��I��9IZ���6\Y��e�5���lcl��Pqukq�+cT]6��)�#;bR�i��h������	�eC�vK̼P���r`-�8\N�׬E<�X��p����g�V��Z�3����^2�t&x��d�3������tg�c�m��G	ۥ����2�4ͺ�G]����C8G�1��(g`�4�5C�k�2�O,H��;g�т��t���%Bq��1۶P3��V�
�c��x�ώƹr��������Rp�9	�ж�k���;%ƀ}����nڗ�t�+q��F����wsP!�ET/*S0�JH9��!�V�U(V`�t)�fҲ%�dU�vv@uL��U�S��H�,n�h�ݭ=���s��.�y�<1��r��ւ"�؎1rAӵ���R2�$6��q�'kn!4>���L�m�iC����'�K�4 �s���l�iy��@B� r�k1j�8�*�<�J����p�3��D��k\gn��u����F��(9 ��;!q�qW,[��s'3/�A��w8q��-4e�7%9��Rf��u�f�m%6�8�ړ��l�;�C�������}���z����ꠞv$;�}A�H=��F{R#2��g��X�H�n�p��C�I�V�t-��_z�G��]2��:�FN�^ink�U���U����(J�9mmJ6%`�z��ѻn"��(�;uz.�vr9�q�;�憣�ی�J779nC�%n���pj�8�i�m�/=!�氯�t��Wg��������=%�� �o$�n�ʮ�w	�Zzx��i�/E���o�[�޵`�	��h�3�լ���7n]�;.r>���q��c��9���;l�W���U�sè��R��@f�_7c�V�o{�@_`h+Ʊ�G1<Ȝ�w�����ݽ4��4�*L%I	�f�T?wE voM wwM۽J��`c��Jaǎ8��n� n�����8��|}�1cbjC�D�P�t��Ԩ~��{���~�~�������t��Jt[9����f�7���2�{;�J��]0��+�K�L��$��}�M8�ۯ�u{u��n� }��lqd�%Q'����r��2���Ԓt�s��Pf��{�N��j1F9�2A�9 �����3vx�1��(|u�3&5��1����ݜ�zi�>^�| �g ߰<x�8G"O1G' �vx�5��(��h{�h32d���~~b{4l���d�g����p�"]�ݫ�������ٮ���1Zt{j��P<�`s�ފ �� ��3g�y�y�l��dK8��~�� {wg �4�׺�s=�y�<m�5#k[�*���ʺ���r� ;Dh@
@"I�� �[5�����|���q�9��M9&�������-�z(��h�j��G���'�w_ ��u�wvp��Ӏ3��=M��")��ݴ�qa+�v���:9�[���6\��{;i�t�
~r(�O�d��r>�������}� ջ��uya���1�cNG�����?$n� ���V��`x�d�$�<Ȝ���Ӏj����Ȉ�_'�z �u�/�Y'R�H0��8��|�}������/�DJ��ҁ���ʽ��浭&�{�pX�� ��k������N�w_ 3��jz8�F�$��X<�kr�s�I��@��y&m��C%nUs�"�ۛ�61�B�ۏ����=�M8��_ ��k�[��&Lp�$i4���>�Eo��@��@�]�rd�%Q �8��_ ��k�wt��<P��S$L�%�D��&f(<��>F���7����<P��V�<�8cQ)�D4�| �����<P���wE�탁�s
"^�/N`gbv�v���K[i9z.���jwA��`J���{�V6 .1��eݣjn�5H�6�H6`��nRƚ�%H��5�C�����I�B�S�5���I�[s;n�����{\��sj�9F�1Y��G>ݟ�~vc'�9d2�Vu��ӓ��]�z;Gtgf|�u��t��N9�n����3f����s;f��u~���i>~�諱��.ݝyk��?A���J�qk�'iFn�zFbx�ǎB!���=��[��wE wwM��ʝȀ&HH�!�5n���G�־ [l�}� �ǈ��z�pX�� ��u�wvp��Ӏj�����"m6��ˎ�1@3$���������@v�r�_n��OrAƲ~x�NI�36x�9��(|� ��ɛ�x66��Zm�\�6�% �!v�v�U����'8s�M��;v��(zk��tX{�@[�tPwt�2L�2V��l� ����$�	?,r��W~��w��0I3i4�ւ	K��fL��˚�g����@Z�����1������|��@wGs��t�����P�d�!)x���3&I>�������z �� �����	����m����=�u��h{�h��z;]�rc�\�3���tg:rq�����7,V�=��q�3����1�.ۑ��S1�c<���/;��7���̍�5��(��^&�PDŌrN {wg ���\�w_ ;���-�{�c�d��F&ܓ�fF����S&��d�Bd��bwǎ���vp��'�9�86҈cqp~��;��7���̍��s���9�2A�9 ��u�ۻ8�?j�[����^Ǭi��y&)�������m+�p��ٌ��нd�nP�i����Jd���r!����vp�~��5��(|�����P�`��.N��ڹg�V��>^��ۻ9R=�	qxcH������ugtP�t����������rIwP�b^������1�z(1)P�&IB$�wEs���Ц"!�^G%?��| �ݜ���~�����:��|�<�%��,l$QE���8���1i3�����v�.�e����=+�Vu�VKJ����fh|ފ����;������۞[S"m�!���7viˉ/Z�m��}��� }���ƜNb�x8��:��| �ݜ����ݚp�/	���r!����t�����O�wE�ڇɰǎ2&��I8�?j�=e��|�k���83�bｱģmD�!̙�ћΩeEI�9x���k^#�;��㭩��BR]���`w98�+U�)��7J�����tF�2��J۰k{)�<b؋v��$���$r��l�<g�R��K½�����kxv�����W׌8]�k0V^�EU�.���E����9������C��l�P�Fsr�Ȯ�����[p��"c��/#]/@f4^�������w{�����Z[��յ,&�(^NI6{*NQ��� ��Λ5�`��`�@��"ǂ����7�j�����3#y��yhx�㜒]�)y�������3#y�ݚp/�5�m��2b�����@fF���<P�t����<L��ZTL3@fF���<P������ۚ�Qj1D1���f�>wE owM��@j�� �r��[�N�]�vZ��չ���zu�]���5ʚ�w9��{\�R�Cq��ٛ}�;��7���̎����I[�{���jщ�X��܈m� =����?g�$
)B�	 :Q�ד�@ot�@c�tP��u="��a��L�����O>wE owO �}��@��"ǂ����=�4�/������;��\��~�hI���N�K̍�������{�K{���W��??�j����Q�jm(!�̆a�@�kj����N�@t.�Y�@�=*�@�!�����^�R���3z���P��*&���j���^f�6�t�2��^y"BQ�ːDM.���^f�&_F���W��+�&�7T�⎟�g]`z|��즑�C�	+@�����p��0��6�͹�$6�1=p3qoF�j��XP����z`�u��lW�j	ܮ�A���,I:�C,���uG�0C�*4/�f01$��) ��1�,�+�4YC���1d_x�zd�Du|w�":{<{�7�t �c�	>C��^/�p��0��R�߻��)=��~��)JKw�<�䩈��0J"bJf@� e�����R�����)JN���=JP~Ue~����)JP�����f���z������Cԥ){��o�R����pz��=���qJR����Cԥ���w��￀M��4�O�"q��E^#dh��`�=�ӌ*5�n	�l���c��l���Fo[��)<��߸=JR������)I�~}�����R�߿~��)=��>�ef�ٽef�kz��JS߾���);�Ϸ�=JR��}���)I�~���Sﵑf�W���7���)JN����R����}�)@�w߿}��R�����)JG�6*�TU4
)�H��96��)JN���=JR������	!���*f��������R��?fj�5D�\��U5�r���[�����C�߿~ڏ����@�{�Q������m]6\m�\Z��m6��\�<7V��� ]`!"z��ݬj~��;��7-�5���JR����8�)I�����R���� )JN���=JR��G�\�1����D̪f@́�{��f�R�����)=��~��)J{��R�e��2���(���Q10D˒����)J}���qJR�߾��P���}�)JR{�����R���l�>�W7�z�Y�o|R������ԥ){��o�R�����qz��}���)J�[c� )���`USJk��9�ro��JR�������^�)O�~��)JR{��}��R���!�	����Gm��4Wl���	���غ���W��q�]�;�6۵�M����1�}��k����d,�*�gD��/+�� 9(�W7OV�;���ݼY�B�������F����b�Y�)i`f�X%��#��Kmۗc���<5���hE�o=E�u�B�`��P������k�u��6�u���Dz��&�t�i�Av�u���{�����|��X����;mլ�:�>e��:'�;�;��LX�E�֭�s�MӲ#��˧{┥'߼���ԥ){��o�R�����q�)K߾�|R���~��٬�n��hن����JR����)>��~��)J{���┥'�y��^������?���uh�Yj�����=��~��)J{���┥'�y��^��3#��M3 f@�;�^u32��$J��Fk[��)J{���┥'����^�)K߾�|R���~��ԥ)y{r%D�Jp�%1%3 f@�7{��b��N}����JR��?~���R����zf@́�-~r�z^�3�D�/;�!����s��]��{m������>�n_�&;�B$�"e�fi��d��{�L�)I�}��JS�u�����2��)��d˻�;��4*�Sy��)JRw��}��<��}�x�Jk���┥'�y��^�)Os����)Iߗ���U��f�ov�{��)J}�_�g�);�Ͼ��)J{�}���,��v�Ԛ�d˺]�<y92:����┥'~���^�)Os���);����)Jw���┥'�������.�$D��3X́�k�z)�%'}���)N��\R���߽��ԥ)�L^�|fk�Q��e���N��8r���x�$�l=r�x���ah6,�%��+$UIRR�M)SUUS|�9�ׯ{��Jw���┥'����^�)O3�~��)?�~�~���Z�kf��Y�k}r���~�ÊR�����qz��<�}�\R����>��ԥ)�e�ٛ�ʳV�[��)JR{�����R��=��qJx�3킲��-KS����F��Ƞ��MH��AC,RQ���9&}���z��<�߸S2d	�<t(w�B$�12�4�c%)�{��┥'�y���)N���R����}��ԥ)���e���Z�Voz┥'�y���)N���R����>��ԥ)�{��┥'_w�����6�=m��V��]m��;S�������;��zv��m�s�VzvI��IF�[��)Jw�p┥'����^�)N��~��)>��~��)J{ֲ��k��2�[��)JR}ߟ}��T�;�=�\R����=��ԥ)ߞ�Ã$�nwy�H� �H��k�R��~��)>��~��#Jy�p┥'����^�)N�ﵯ����F�ļ<D���2�{w�I�f@̷{ԩJR�����/R� *t1���(��hg����JR�����Zݭ;����f�[��)J{�p┥����^�)K���|R����=��Ԡs���Bd`BժJ��T� K�$�q��3G���M��=W����.��:w�я��o[3z�V�oY��┥'�=���ԥ)w��o�R��y�qz��=��qd�^x�P<y�$��%C���5�ʔ����?d�'�����JS߿~��)JO{�︽Bҟy�ڵ��Y����e��{��)<��~��)Jy��p┍'�y��^�)K�~�|R��Wƿ��PL��$�M&��2���qJR�����/R��y��k�P���O}��R�����f�ff����e�٭�R�������ԥ�DB|׿�k�R�������)O<��R��������0�$ ����{�p8f7Z����Ƚ-u�Q��.9n֍�sŪ�g�\�c����d�Ӎ�{5m�O5W[])GHM��������۞^w�S��N�Ϋ$�@繸tTq֝��m��:�$n�ur�@�w^s��6�TQ�����gZ�1��rog�WFqp�{j�c�Ɍ��n�9z�;J�]�Gγa.�N/nv�9�8�vޮt���X7�q�uk���w���~��|�]Q��G�,�[���n]p�'0���"V��8���S���6+�ȖnSf�7�p{��=�^��)JRy�����R���~��)J{��=JR�絲�IN<�E�߰?~�������)Jw��p┥�y���)O|���2d����DD�1)�`"i7R�����)JP���}��R���}�qJR��>��R��{������kY�+z����qJ_��������R����~�)JR{�����R��߾�Ő3 My���x�"I�$�/3L�3*S�u���)JO|�߸=JR�{��8�)I��}��JS�M}�����{6fcv�^gnιn�7\��&����F.nɼ�%���K�7��Ex{�g ���m�v�=��~��)J}��p┥'�y���d����2d��{��$��fo|�)O������\qQ��,V�:4萈(Ј����2R�s���JR�{�~�)JR{�}��P�<�_Fi�Z�ƭ�2�oZ��)JN��︽JR�{���)B�'�y���)K�~�|R���}��kY��f�a��7�/R�*�{���)JR{�}��R�����) )�{}�f��24�Dy�yr�0�gy�)JN���=JP?g�}�)@�w�}��R���}�qJR�ߏ�����C�[2Y:P	Ӹ��`��k�r�D��vS�c��C�mX�_v����|Wfr��R�����)JN��︽JR�}��� R�����pz��#߬��_;��2��fo{��({�Ͼ���G%?~����)JO>���R����}�2`f@��G��Љ%LI**&��5����kﳊR�����pz��x�Uv)K��|R����=�Mc2e��AB��P���̩JN��߸=JR�}�~�)JP��}��R��>��qJR��k�L�|ƶh���7��z��/����JR��|��R�����k�R�����pz��?��1�2��B]���˓g<���������ڝ��,Bն���ۓ��=����r"&i�2۝�Rk�3/?w���);��~��)J_y��┥'y�P;�!��R��&i��d����JR��=��R���kﳊR��y��3X́�w��C�3����f)JN��߸=JR�y����?�2N����/R������┥'������X�Z�Z�k|�)O��\R����~��ԥ)�{���'�5| ��J��I����R��}���Y���kfV�o3[��)J���=JP�	��~��)JR{��~��)J}�p����m�����~���^y��ʃƹ���ە{
\a�{!a�fZ��C������:G�N�a�D������X́�y�ފf@�I��{��JS�}���(}�Ͼ��3 f[�zxr(��.A��3 f);��~��")���ÊR�>���pz��>�>�\ZR��+�L��8k6V[�o5�R������)JP��}��E)O�Ͼ��);�Ͼ��)Jy�̭:3Z�#{̵����R���~��߸=JR���߳�R�����pz��~���qJR�����}��޳Z�٣�޹�R�����k�R�~@���߿p{��?}��\R���>��ԥ)�����|L�5����8�c�L��� H�Q,�(Q���+�hY� s��ZQ˨�`@���%�@�	0���D�$L�Q�ٔ�QCa�a�A�f%P:H fH���)d��d�, Ğ��٠��'zI
���	I��D11!XI�Xa��Q&)�"΃X:������t���O|y*�a�eB��QГy����fm����!V�KAYTMDA��\ti�C	���� ;M����b��6Xm]`QQ@L�6o\��-$M"��8G -9eg��(Y��bB�^�ߗ���O����W-�.��\�F�]ME�v�(J�Q�g�G��J�$�d-���Y�3���cs�t��팩ɏ���K����ׯeL�� �>M�K���A�J����q����j��ŝ���ў�u��\�9�뭙��;oml�8zsz��u�`�r��m����������:7�-�6q���$7DHV���l�=�"��)Z��m:{`�4�̍�Lcz�'=SmVÓ��F��iCM��ؙ��+��6��F{1�H �qi�6�f��lp[��陬S<���*�lL���h��,�*KR��*�r1oR���A�V�*�U*�j��
�t��TTY@e��ڕU@�Zx\V����YL���ƥ�I�-H:��b���R���9ӄ����@u#��l䛖�9�C�ej�2:ܔ囗5O%�C�m��J��U<��`S;����`]j��[��8mTX����4�U�4��۶�+t�W�\wQ�s�i_h��tm�]����k�
�9-�t�"W���|����7<�/Og�6޷Z�q���/�\�zh��n�B�|s˼Oi�����8[=^ݻa:��Ó=��]�q�ɐ����Jzq7�� 8�@9~W+�RÌ�u^9�S<&���:V�<:�����
h���-�r�#�Nzlwj#��q�����\�W������D���zf�.�g	Ӟ�S�j����l��I(�gF��-cEk�nI&�Ф���i{-]E�uSh*
X *9�;+�O*�d�*��m���D���g��U�+^v�z�[�7�]�y�G�{[�"�֜��#5��:�;`���ikh�R6�$�MK\j<N`9�姴�*4�6��8��Udqo5�ʠ���ɐO�F�MB�YS2��©�<U�;8kЩTÕ����a,ՍI�v8ܻ�3�B�q,Y�����e`�6�L��{��8���;���yƉ̑`ՠ��E:�n����| ����&nݭִlֳe����#���0��g��3��WJ�(�	�� ���O��"`���:PAM~�ߣ�o$��V�nB���&�ZLLf�ۆFO�]��pc���[m�5nqi�����s�<,�	�����L�l��4�
�8��j[��M�lYxr֍�.�i��;v��N��G�pg����Z�d't=8�\]#���p����E��<�-V�/f�,�Ν�M���bAvɘՀ�v�v�%�մ�b�Kc�s��l�ţ��+L��o�+������ &&^Q2ᬲq�,���
�.:�n�4�b�݉�E�{�3�;Lnp�����{ݷ�������ԥ)���┥�y���JYc�́�.�yyɘ�����r��=JR�{���JP��}��R��=��qJR�����P�JGY�C����S�A0�S2d	�wޤ�3�y��k�P Rw��}��R���w���(�JRw{����~4f��5�f�����)B y��~��);����)J{��┊��y���)e��C�D<Sˑ2�� ���d�f{�=JP�/����)JP��}��Y2���́�+�s����3/.�'iY���!:�e�d�];����@|�%N��k�oU̷��췻#7�o5�R������)JP��}��R��>��p? B#���~���R����Պ�|qD�D�2Pn��v��P��1#+R)- ��A�&��2s_޸�77޻���|a2L�3sbCU ����&*���^�@�<���s��S:�y������<<�'���d�#;}�;c��ۭ��x���#ӯg�<p�T�JH�P���<M��>(�2n������z(����{=��U�piH�"NC�%�\Ϯ�3l�ۭK���˞�\g�D����{ݫ�#s�(��q�p~���+������"#�r9�����&��\�<��T�UUU����S2L���{�`gGy�پ�X̓&L�n��<A�LNc���m�@�=��ù�@Ш������3�~�*�Ƚ=̾6[ݑ�޷��]W�TPG�w���ٻq`|�9�8#�Ȉ^�>��u0@�=.�%�y��/��Pɐ��l���s��3c�������L�㖻L��K&t�mT��y�ZѮ�N��_i5��Vu�������*ʺA�5�~����P��]���I�s��VWZk�#$N&�&�����Oٟ�6;�@n{�j����Rd̀�㓼G�LBx��n����P��Z��L���{뷽 ���G0�&")U=����Gn=��<�����~�����-�A�@��~�*�}^"��$D�9$�t��| ���?�>���� ���`}!!Oo��qa� �pZ���l�&�q��F��u;�}���ܟ|"��l=[:�������zh}��fLɕ��־ߌ3٩_��b����wl�9��k��[�=����Ds���ʲ3Cv5��rpo��|�s��Ds�?c� ��]�1��P���𮞪��d��?��7�޻v�~���m��t
�Zku�5�fjz?c�y"9�N=��=ǽ�>^���ܭ��d���H�aՓGj������Й=�q�غ��&���<�o��aaxν�c��JM��V[G�jR6�6������UP܀;g*�7�cf�qs�ʻ���Q��9�V�n1�od��8N����\uc9���G�2�tv���� -76�U��b�9�i�u�L��<��ݘ�Մ�;.Ӷ���e�I2D��m^IZ�g�������|��,�vy0!mf0��;����el!5ˏ`���d����5?߻�8��YC�LNs�j����v�|���?f����QZ8���E �| ۻy�>^���[ށ�������b5�����ns��/c����ݑ�@{Ӎt=��`?1�rI��"�#�~����{�=�����X�>��@_\��
Q28��Jj��8�@����!�n�>�� ����/�Z��PqO�1���[s��a`HÐ��85�<�\g��t�u����g11&��q!��p���t���������l� ��k�T�,J��7��`c�z*��O�o�&JRT����:{��_�#��Ȅj�(�L�"J%T�3S�=��vٔ΄D����>Y�z��S	T(�)MH�SWa���z��n�X/c����v�q.��2b"�q) ���΁����/޷��{W �ˍ,�&��4�#!���m�<�{Gf�\��69�r=m6��݇đ��&D�΁�ݯ�_�oz���f}�΁�Z�Ԁۂ�"�&b��o�v2`Ύ����Z�1���9�}�7T��AT!P�k������ޯ;(d�.IZI���k�z8����г�i���q!�$8�z}�l����6���{�L��m�M	�#I�|��/Z���}���ޜk�|��u`j�A�)�K�Apn˳iչ�+�팾�$�`z�&�n�T�t�AM�9b �c��}�����y�\�����~�޶p�҉� �A8���z���g�����y��{���9��DBi�*v`���E*�Q54t�{�����DG ��n�kڸwؒ7(��	�)�qtL͏��P�޻z;�@)I7�&e��c���]�/�pY$B�|��;�1y����Ձ���@؏������9l��Nv���sŷ���.��̩uӷ'd�5�T3�׽���ݮ��z�ЄUT���Y�=��ڰ<�9�#����n��kJ�ͳ���G�3#}�&d�����P��]�Ͼ�W�"9�q�7�D�*bUR�L+U�Ձ�^�@��7vDDDp1y���}����ܘ�Pl�18�xۏ���3�����k�}�j�Wk��iF�� �N1���@�����fg�yں�mtf��`JJ�̒�G��yxre�4�X�rXѝۍ�B��PwQ��kf�^Zct�ɍ]�2s0uu��`� ѭ�k�R�kBUH]�[��J�y�L��M	W��prd��X��vZ�$U���������'?od���kx��y%Ph�y�W����{6M��ʯci�]��=&q�����ֆ�g��ي�0�c<�9X��]��1�[���k���X�/;��˽���+�v�<���8��āA�q�<	ұ�U�)�q�G��ӺJ߾��X��p�ƊNJ>��u���7=���",d�] o���^ ��<��&*��~���0���G�17��=��`?C}&�&f�2�D�P��]����L�fϼ��־���1�� ��@��3���}�>���y��o#���{�`c��a�-�*H��U=�y��Dr>^nz�cw`y{�~jR����,�{�v:��/\���ӵ�1�u-�n;sk7X�=�<f�}�[l}�����z�}�E32`3=�����,rL���m<m��=���^~�����D�$ft�A&��&d��2kL�%%��"��ޯ>��L�3$g��2D�y��`�v�������ş&I�&d�|�w|��@>����18
%$Y��}���@3}�7w޻��In�y�ݮ9�/��<��&f���zh�&m���@��S�}���@�Ǫ�X���۵+�ە�[l[����K��捲f���=���U��9/H߮�y�>'\�:����߿����`{�L�|�Y� ���@A������������e3��=���`{��=�7w�s����&��2-�*P�&&Jw���Xw�4y�Z�BC���&J�p2�w�Gھ�=f�Roz34.�]\1٫1��0�l!�,l�펍�sqG}s��;C;�D�.��P���ᾜ]�͆������:��û�&p��͘�ځS�'eqd� kBP��$�V"�Ԇ�u�M�v|㧁4I@yP�	Sa�H�0�y��d�C)�^z�f�'H�?'���b�K�O�ڎ�Q�E�}:Pn��ɔ�I%�)~�˰;}>(���&��B6�C���?m��}���@�� �޼�@��G�8��(�h���37�v�O�3}^,;ޚ;���vɿlPySuF�0ŝ<���'gs�us
�<����jx�n�΢��۫������{�������O�2V��f���{
j(*b�RUT�jh�|������݁��g@�H�0	��*bbj� ������z���!�i�=�}��i�q%QQ*�T%3@no�v�O�3}^,�I2g_m��}C��pȀpB��ݔ�}��2�>��}���b#�RF��N�v��fl[;�;s��/>]6'�v�`r��Χm��.ہ��c.qq���,{7�X,nz��w�)����M�lC������>���@�� ��Lz�yc�&8��i��8��{�=��~>��S�z��>���d���bi���{e8�[�t��|����ԴM��pH�F�) ��yN���}�g ��]���]y�Lq���4��j*��F�hw���
�T�΋n�4p��D�+j���v��ʊ���ˋv�e�`*C����7&����ʋ����.����N� ��d��^�;��̇kvݻ]h�����"n�V �3�(��O�^ɏ��3��Q�n2�����0� ��]ӹg�."{F�<"8�+m�0u��v�v�,�u��ekffl�|�� ��3fsE�i)��ժK̖�6�t�ob�y��g�%��jEDԯA_��}|Fw|gC���7�f�����ｎ�/c����:�䌲$@Lx�D1����������t{z�X��E$��#yx�("S�����<���gYg��G�ݞ���n��I�$M�B��������,���������G���@��	��0m��I����_ 33���@����>���@�� ��G��H�q�!�ɓ�ۮc��q�.�Ŵ���o4��{3��k��1ąOq����@�ݱ@f{��2V��M���T��#�'��ȉ�_{�P��*�:L�BL��D�E��u^����uW�翵ʺ����Sh'?D�H�G�>�w��1�ފ�2b�}�7�����:�&E�P�s�:�?~���j�wޮ�/b��D~�p�1��*��)&$"�|����׵p���:�m|���i8�i�6چ�! e��8�v���䝨|�:b�g���n�����_y��B99�]�\��嶾f~�z��k�~�*�Qby$����W� ������z���=&@f[�D(&��Iw�@>�g �޶�y*وd��.I*I������S�yz�x��M!D&7' ��oz�w�����ŀɌ�zh��.��F��8�ӝ�ݔ�g��}m�@>�g ��oz���o�\D�x�*�'N�rr;��eRr�%�7Ev��z�ɋh &6<���"�k$p�~��|�ފs}�fI������~r�"]�Q2�jjj����z)�L�fo�v�ڸ��[:�EZ�7���D�7$���]����3$����Xw�4��i�
Z%8�L݀��-����Xw�4�fL���]��vvxP���S% fo�VfLg{�@}���@����;�P3h'��H�=c�4� e*;jEޥ����Og��:]�2n՝f�ff~�'3�(��Pn$��9΀}�g ��[ށ��}v�m��I'Q���!I3U�=�7w��DB1c��������wy� �!�Ʃ�4�B��N14�z��π}m�@>���{޷� ��q7?$��F��>�ف��}���t����"9��c���|�u�����Lr"r>s���l�߳f���^��|��lr!s�K���wD�X{j�&ks�Z�$��]��u��\��X69u]��x'۶��ZĔn��P�Ͳ�Z�Az
��!��]:5�q�Ib�H�۲�g��ZySq=���k������wV1�7Jͧkm�<��J�6���\s�cx,r��\WF��^��z%�\�0��np�gh(Ŷ��GUH�ny���*�&��c�I��4dF����iz7M�N�>���w{�}�|��QV�nm���+�YvC%��[M�6)���˚'���~�3��L��T������v�q��|��l�p����a��lRw�yn������Xw�4f��bL���#�bCYF�x䏀}�y����>����yz��;�m�*$p�!.�9�X�7}�3w޻_}��3$�2fv�7j�{�;RTL�$�W@���^nz/��X��tlN���]�2�vAѱQ�6L����n:3\rx��ӆ�I��cS����'��Ƌ���R��`yy��}���=��yȋ�� �Ƿ`ֶ)UL
��R����@/����3&�fV�fUA��M�������� �n�i1Q�DNNs��@=��}�c�68�d}���
s"�\�S%B����o/f=�2wW@;��΁��־ۺ�\��d�F)5v�-��������b���{��������o��ЯR�+�E�z��gb��c�]Y,v-�'!�N�t;�b��}u ��L���qp�m��^����{�=�j��=���A�ɉu�s��^n{��y��=�mtﱾ�ک
�A�k���������py�?Jz��H�9�IU4D-'ȯ9}��yΪ�����=�ʫ����,N14�z�yڸ��o:�[8�����U�7�&(��a| ��z��>����־��Ɩ[1��)��ck�P�1����Ϝ�v��)��� �)�e��ۧ�8Y�B1�d�9�s��־����/Z���y�/�	SMOͼ���T������7g�c����������T���B���1c�����͂!�v��݁�%�Ġ���A0L��p/�o��n���w`�:eBBZP?~C@���_��(�˿�i�1�8ƺ>s���k��ȅ�f=��b�������"<�M53�ڮ{TͶ�rډ���J[>�k���I�֝R�ҋqc��Bi5�;F�����;�<������Ȱy��󆫂���bi��/Z��߶����f�tf=���G9�{Z�U3$��y�tLLPo�|� ����$���ށ��_ ��=k2��'9�s��y��{1݁�����7��2+qF1�dō�8�ݽ�^������zhnft؀d�0$˸rE�R.�٥r`�dД��Z5l�NPp�4��h�8GxZzn9A�I�XZ��1��K���)P��JeGVD��U4�H}�4HUA$��i���	���
'�~?���o�n��E(8D���9N���t�k9�[@��T��;F��tenZU����"�s���K��q�%�s� �6[��v=�.,F�@�h�)b�s��%��c���Y��m�\�:=��s;����u�sn�m�����Ϊ✶�s��u�m���{:��t�N9�R��O�$TUk���/&+Y�n26�LbR5�WN]F�͂�n`�'��v�e��l�Q;m������jm�����EE�j��ٹ�f�j����K�uխ�+H	7.ҁ�n���݀��4�u�`�mR��*�ԧ*�K��l��� ڶ ���N�mm�h��Cm���K�����m+�`5�� *veL��R�b��C �l�Z���;@b���U�Z��=�+0��nl݄�w�va�V��jE7$MU!�Ny�7�q��mˎ�u+a;#ɳK!;i�;l�6�N1��n��$�o!�H��.�i�[W�x;+S�]7`S0�,C��I��8��μ�[�Sm����atCl����`.���At�G��g���g��ODF��s�D��VKWܻ�oc������mg��]�mK;ZdO.�Ipbۓj�eb�	���au��U
�U:��T�e�3�\��l�Z(rYk�xX�
��ϓN6�+����,�V�k�<������+%é'TN�M�.�r��ζٹӎ�B9۞۶Û��1i��d@�b�-(��%�l���Xdt�MT�+RnD�\���K WZ��9��s�[����������V���Q�>� �;\����g�F���qۏ^���A�i���� ɣ�Ç�����'a����8$��V	EFU�Mc{*�]<-]���I�],���)���L�PU���'8q��<T�˩�pf9@��������RQ��I��P9��Gq��m[OZ�,�=*��]ύm��ˉ�(S�dg��+$pəu��FuL��l[N����e�l�v�D�����g��y�{w���ǻ��yC�|EO](����C� ٶVEvm8�j��º�Fk{��6��T��%�iֻ���|My8a];A�N[c���m�q�α��ɲKV��:J�9��\�ٹ�nV�[��萌͌��̕9��5fg����'�%��טxf��w�Wh=f)��L%F;nzl�n9k��]&��:�Bƣ�{v��R�yݚ�a���c�gt����ݞv{�d�n�'��鱳r�^޴MgK���{��C��]0kn;n��V��s���۲6kJssu�q��'n*��W:*e��.q�?�I2`#��-������=���fc���$A8��Dq�������}������v"" �歀D�TUQ5$�'��l3v�٘����s��o�:�
��OXD&7'�v��yz����΁����޹UpX��C�%3W`yy����{�f�t�1��~��D'RA1��YSډnح��N{d<��Wӗm��k����t�}��}��!D����wm�@����}���ٜ�,ݞ���u)JF�R**+��{��^���ٙ�!�m�@ջ_ ;�o:���$Cc��ɉ�G�>��ށ�����l/7=��d��D�(��F7'z��| ���^���v��{AՉ<e�&,xۏ�ݷ��O����ۻ�㞁~�R����g�⻪�\��닅ٺ�<B�x�{;L��[@��ۛ��������g��������f;�<�9��7�ͪ�sP��)
&f��}���b1k���������{�sB��UTԉDM���E��E�K�&d�Rj�<W� ����}uJ(�Lr!E#X) �=��^����ށ�v���X�k+k#b��s�}W�|���^����o��IG"0Ar1�t6݇�/�}���%�<:utmלv���2��"#&FLLr>�}����v�����/Z�s�m�`��X�!J��'�zo��`b�s�=��݁�RIbx�2LX� ;��΁��_ ���ށ��_ ߽���#xڪ�+'��l?""9'7g�7�n���s������3�k���}Y7vu|�3�=J:�q<�D��b&(}�w`yy��������s�=�r��p@jܗ[�T`�!b���q�^�R��]؎��۳s��䫅�.�N����9��7����f{�<R���9�,$���o;���[������{v,{=׽�*I��˓UUUV>��@gwz�}�E _u��w/&H�2Bdd��#�/[��1f���1����s�>����@�$�1���@������΁��_ ����~�����<���q�RC7�q\v�ջ)��kF_c%�`�B���ܜ�s��U͠��Q�v�����[��T^6�Z��V����[�mjϨ�ٞ�Y�i��*�����6X,]F���r�9�p�]�x��5�;m�d�)�qX8n�e�x��s�@�J�gC�ڮ�n��^B��<0u�kpa^�մq����قb�	넟L�k�U�jCxnhحo߻���>�k	%���jwnE�%� ��Dh�uk�j鵳x�ɢ으� q���I�����^��wv��@>���}���FEԌK���:���@��w`y���c��G��`HX��!�ő������޶p�ߒ>ݳ�yz��=��KA���I�}�] ���`yy������"��y	��"$�wv�j���wwoz�p�Զ���(D�L����;<�G�+�>.�� �]�n�e
r�����O�ﾑ�q��"'9�Ns�j���wwoz�[8�ݼ�ڊ����#&&9��/��wl�%I%ɒe2�����������{BI*BS5\��� �{] ��}�>^nz�c�2����c�����wm�@�m��}��� ��~����Ȧ%��UX��E����zhs}�;��6���C��z�3
Ze^D���ն�û
�f��ax;cvi���%�U�A�1�b��|����l�����[k��-O*?����@=��~���H3ٻ�ݞ�����G��'h�C��ԍrp}����m|7;���D1CM	RQ PA
J,0�,K(�D���{ ^g����g >��I���'�(��s���������ͺ�o!'�{�^�l�i)�D�IP�������=m� ߽��V���j+IUNO�k8�D5\��l����Y�1P���TQM�xۙ1�����FI'z�l�}�}�1cs�r ��w`fC��<u౱�8�{o:����m�@=m�����q�#��LK�rs�,nz�c� �n��{lyP�ȱn1dn>�������������u^�eBa��0qA����2���Ħ!&�m9ހy�]ar��~��=߱݁��e$?�]n�s��l���K�EN��b;	������2um7j�;7k�#snmp��SU����`b��[�;�,��t�{ZL��ȞF�'9�Ns�ym��w뷽 �� ���Ι���D<����|��{�m�����@��_ �]ې @�B29;����=�������@�����$���&�$�W@3�7�N9{��>w���}�M�k2C!V�!�T`߿~<��[V���nWu���]m{v���x<�WR��z!�/O'����\ml�6zsֈL �� j�%�-�������W����lT����ɝqK��oAt�cr��I��CBM���c����'q�=9�����3%�3f��i%z��L�p&;$�l4/D��E��%��m�:pmlN孋f%�-Q�fx5�����O{~���~��q�T��U�һel��n_9������Ɂ�j���ŝf�nw.�Y������l/7=�1݀y�]� ?���v`	�� �#K#q�����~H7wk���7=�3�1��*T̍6�JN�������U�_ �޷��n^8��ԍ$�| ���Z�����m���jI�[Y��D�9�s������{�*�_ >�m�@���%�7qH%`�!� A��9C\d�i��ױ��p��-]@�y�>���1�d��#�{���U�� }��΁V��r���c��!��]U�{���¨D��R��I�&�U����ޫʰ5�ފ7|��9	��% �H�M$J�U= ���l���p��n����|�\L�T�m��9�t
���>���@�m|���o:�1	5r$�9Y��}�7v�6^����{`5��@�r;������n��<u��h1�<�ڨ�%�Ɓf�m�'�=�,ipNn3D�ݧ&��]�IS2�)��Sݞ�}�o�X��9h33v�h�{5S �%R�SS��m��k�����cs��0JHs*)L*U%w��{��nz��wg����@MǿƏ�u��ܷ?Z�-�^A\��@7�2\2eڬ1Q�P5 �R� "@����Cbb�z-���I$!���-0@��X&k�4�rm�Cp��{Q7f�ѭ&�vvfX&�:ᰍ��4��l䡲�tc�3�"���V7��"<r)@�{ְ��`']��^����0d�f���(��F���Q�x�?�
>����#��7εʫ�[΁�E��q��2bc��?����f������>�cs�.�c��#�������t
���=���@���m��8�#i���V�:��&���*k��[���Nrty f.i��fO�$4ԏ�}v�]v��z��
���>�k���##Dx.ʮ��X��c��>�ݻSݞ�}�m�@�f �rEnH�F�����@�v� }���@�־�e)T�m�i��
�k��n�t
�k�c/	��fJ�2it���7Ǘ�ffr"0p��H��۷��Z�}�n�y8�@�r1Ѳ�n�TQ0$T�$�� �Á�i0��ol!�у�S&WW^�t�4%$uT�*U%w�����7g�_��z׵p�o:��V��(���jE�;�[ށu�\ ���΁|�\�s�	Dn��(��"I��\�] �����7=��w`fCT�)��8�0r. }���U���޷��p�ช&8����:X��{���y-��_;�DG>r�=�b�
6!���N�0 jBJ$ᎀ�"������|�+:�����G4�⅋tx��˕��=���'��</-�f��m�ۭm�J�C�e��g�K��*��.ҍU�Y�6�M(�ukS2�c1��I5�lm�b�޳�N��u�͏]��m�OR헗sv֝7h�9�;r/]<���[%�[�x�'u��u�vɃq�j��:y��ce�3�;���\5Z�:q�mg�I�~�뻻�s����t��W����+m؉��<�>��n�+�>��Ԫ]�uȇCnl���������������7=��H<Li��Nw�]v� w��w�����=3݀��UU���D����΁V�����]���t���LD���'9·��{��31��cs����1�NR��D�11�����m����΁V��~�V�JH7�,Ġ�9���0�^M�L��K��p��;lR=��ўK7^s�G�%&!���m����΀�7;�A��n�n&6D(R���P����ʮ�����Ҙ9	@�`I04B�<��3{�`y��g���D9�<G9�t
�k���{�.������@���!�m�(�����B�1���z��ُ�^u��)]MǓm�i���j��n�t
�k����@4�CF�$��3]Z^�!��D.XG����4�&�SkX��{\�7g����ѬQ��_n�t
�k����@�v� _�J��Jc$�99�s��Z�}�{�*ݯ�|�ݳ�o�ʚ����#&&9{���~�E�I��_z�6��|���V���Lc��������V^nz��f��q(��
Q&�R�$���/�X�[���3��.���w�I�f�Hɹ��h�.�&��a�ý�i�ժ�lX�v�I�Q��v>rt�j��[ށu�\ �}���y��'�&�(���[ށu�\ �}���ڸ��WV7�ƛks��ڸ�}�t�j��[ށ���#ɒDP��@�g�Հכ��y������4�X��i4�kI�`:`d�d�j(a(�r0"�Xوfa��Ё1Y�8ȸ�bad4�b`�E���ɨݽ�boB�4,:�'P�b��\��:�5�E��ޮ�o�5IJT��rj�T���Հ�-��y���y8�@�g�Ձ�Ȏs�������ڝ��v����g�sm�����D�]qy�y[�=�I�k;�&cN�t�O�{_���'�,�:��s�/��!��Ĝ���9;�.���|��e�כ��y����#��[$(JU���X����̻6q��jY��$�&�k��U�_ �����j�����F�����ۋ#q���@��� }��΁W�|�d�P�̙opx #�2����̄����9���n��ط�z��9��%��n0�LN�]8:ׅ��6B̻;2�ٜ��\gD���O/^y�m���/;g�7=k.��e��nP���J��m�c�T��iŝ���K>�]y|X�]O#�̎�؇���&�[�dqn��k�7mm��8r
B�*��G8�ŋ���hXv�e̫�uqb�u��UW��벟l#񛳉՝��(6�l�/]��g/��۞��'�hf�Qcq�����Ɯ�@�^���ݼ�z��;�[ށ��
�"�Q<FAJ] �����7=����y8�w���T�J���MR+���{`j����;ށu�\ ���΁��ypM�1FT*&�zȅ�f���z��ُ�^����q\'1��N��j��f>�y���7v�1�H&�G�v��]���2���18,΍�1Ț�ݓ��ny����;,~���{V^nz��݀�q��bQ��$�&�k�s��U�_>�������oz���>_n��.�S�����ܡEL�������=5//7�`j����!0R�
��3*%M]�9��^���������1}��v�0�aR���&�T*��>Y�u`l����>y�v�ƺ�K	��(����/RQ�ݎ0���^ѫӒg�c;��qvP9�=�'��np�dq��Ȉ���N�W�|��{�.���|��g@7�bo.	��#&6�|��{��]{W �o�΁W�|���Ʈ ���c��^��>^����>�B�x�à�\�P&�}j��hJB�(JS1���X&�X ����91�E�Jwg�f����(hH�R�(RJ����9��/Kǵ`j���������~Է��Ȍx�c�%�כ���
>y�߀���@�g�Ձ�w���_�Uqb���Mej��Ԓb#Z�s�F#=�����i�1�f�Y�-@v����(���[ށV�|��3�_;W ���p�F��Ks������G8����X���盻��G! ��P�y!	�<	��y]�Ӡ_;W�����n����V��?�R*{��j�~��@�y���s�9Ȉ�2���Y�b�a(> p������ڰo*I�LQ�"r.�z���j�/�l����>��ڊ������ ��^���r�a�)r���g�*(�����vC��9�]��q����1Հכ��~�w`{	FT	�j�Qb`�\����Z�}�{�.���w�[�A<`�F0k��ڰ�s�/�n���t�َ�6��@���j�3S��_fn�`kw�p�۶t
�k��1\+$����cnw�]{W �o�΁W�|��zꮍD�O
ptM6�:�ox�SX�+���OR�#���"Rc@�c)Q9�YD�)��z*�.��`�I&�\WDu�ZR� .�섖B-�#����x��:�3�J��`G� Ǫ���c�f�kGy��'4�hD�h�h"*�R$;(zKZ!$�H��2+�]F6`��h �a�aY**
	�H�"pLֳ3�D�	Z���oP;�x��RkQ��i��,��ǅ�2dVVVy4U�ޘ-�K�k�	(Q*���	�QV��́��vPk0e%��c�	��h��,��@��T� �H�:��n��'`88:L��m�;d��]4��#�-��Z
^0m�H��5m��
3p�xGv{;�����������u��v�9�Ζڮ��.���xOY$�j�� ����u��K�k���x7I��gn��np�֊����v�׋� ��]rh��hwm�n��4�l�M����F��/�Ӵ�쁺守�5K�� �u�7Bj��[u��&�J��q<��� �]<����e��j�G���04��͐*����`U�U�U\lh�Y� Z�RZrβ�!��&��`dcm��4ݫm�#]���H,��m���(.���G*���X� �)֦��4J	����VBjٰ ukSX6�-�M%�ԫ���M(ԯZ��t���H��I�v�Л���GM$��i��YFX��Tj�"I��[zm����q�rm4-�m$�k������t�K5�gJ�fc��V�ue;�v�Ń�rp,v,�v�G��K����M�:�իB�)�)�8��ۣ�.3�	�vL���R��v2�/]+ݸ���%�cu�91�Av5�������l�N�
�LW 2��{ub1G:��3v�x5��g	�nL��2Θ��8�(��]�����.�5u�3�:7.��1v��K����]���5�u�X���ɛ,���\'\@{-�����t�m!(��[e����m<��ZUj�q�jJ��\b��n���@��W@�U+ ���$N�Z�p�5�)�P�4�R���,�r������ڎ�oV��/o0:!�͹ku�������z�$��ثUJ�;q#R��P/*��l�v�mA�f�gU`�I��Gg2�$��Erڒ���S�6W��C=v給�{e@�G$���Mm3V��[Y�`��l��-���	�V�쾵�ě��^[�W���6]�omq'7]��mP�R:fn�u�K�ŷ$�H i6\�JA��t��'B
z��<{������2`��`�qUOQ{;���������k߯e�:�$��t�1�3�\*r-�n��c�:���[��e�[<�W���5�U�v�<��GW@l������Ҹۘ<9;{Xݲsʈbⱀ����5F^�(*�8ݸ�h/�W�)��,Yg��3��e�ۗ��vڛMu�R�:��ە�%��/hYĦ�y����������񡝚B�sx]�5�b��K�ٝ�n��p�� ܟ�x����'/���
˰Ȼ+N-�cGj�*p;���y�LWi�����i	�����5	"�j��:^�����G�5���x�Rj��ĕRT�{�Հכ��y���y8�@�g�ՀcĆǗ$B�1�#��[ށu�\��:^���ڋ�����1�r��y8�@�g�Հכ��y����a�x���b`�\��:^����@�����ǉ�bR,��d��B�/h��Y�L�>_Jn�gg����A�;�gC�%2�@�'�v>rt
�k��7v^nw��Z'�j�z��P!O&����w����s�cc^��-ݳ�U�_ ���p���ٍ�ހכ����c���=��݀|��d�c�$��|��g@ջ_ ������p�$ʒq(2FG��{V,�=~y���{gut�{Xo����8�^n̯�en��q ���j��`7�nū��pm�=s�[)Q35S�/<��9mt�{o"#�7��>�n���5I$�]���@�g�Ձ�1�@��w`{	PC��WLnG�>[�U�_g�˘2K��fN2L��s+���݁���/}��*�����0����a�Ų��@����y��,�:�1��"�
yPL����w���U�_ �o�΁V�|~(��Dmņc&�j0j:p�wIs	�.��'4�X��4Wz)�5<�p���Oٍ�ށW�|��:[����@>��V��&�9#�k�9��BF��z�7n�~��@قQf$�PqFH��q��j��[ޟ��-��]�q����	��UATTK�����]��y����Xcf�&�l�}�\w)^%�,nc�'z����>�6�ƺ��݁��(nUs)+�	�Scv�+6юMo&5Ú�A��ط�B���H:�87<p��9i�ޟc���=��݀כ��~�9
�%AUD����f�k1�w�y�݁�7g�}��s`c��T!O
Dʪʚ����w`b�s�R�{6����)��,Q�LF&�z�Z��cj�<��Cy��x�~�8i-��UU8�&G$|�v��]��o���^������m�ʞ�����js��Y���wo7#���,a�{
��Wہ�mr�)nV�F�[bQ�����ݢ��b%��@�`��X�ڝl��NͰ�Ş�wn���hv���I��}�}�Y�uڹ�mÁ!v֞�b\\�r��!;Q���^-Oj�g��ɐ�3xWok(��spV*��N,��<4U�Dŷ�ƺ�Wu�8�b^���v�ѧ����ŵ�YO�l�uĆ%�ڮẌ�綞���Jd��[tۧ}���\'��2N79> ���8����j���|��:�k�q�R�Ǎ�'@�cw`b�s�>X۫��=�H�#�Q�&j$�eU]��7g�|��V׵pn�ށ�($�4_��"�G�>[m��ڸ�m�@�־����BG��'9:׵pݶ�����6��؎qsq':��#//iN;�R��ˁ���v}�6�r���2�qvs@n%1	�@mH,M��6����s�>Xۭ���z�C�-�GQ ��v�}�'I�o&iJ#�Ȟ�>�V^�=������$�`#���&(I �z�:�p{m�@��_ =���1	�A�'�� ��]�������|�� ���h�<J@s&$���{�5z��>[v΀z���tġ���v�ƹ����SD5�En�ϳ��[����vt��#Ĳ%��s�iN�^���ݯ��g ����PypC��C�I �]���po��@��_ ���1��G�4����<���<�Ͼ�g�R	!�p;C�����e|�{l��_1	�Ԃm98����j���|����|}�˃�`��M�;�7���>M��㞁������D�T70��!�&�q=�B�	��f^�1�;r>u�;��i�rv�I	�(����>�O��n�����!ˢ�Q���9�t+�󸑻o8�ڸ��� wLK<q(�ɑ� y�݁�N5��1���y��}�7�.X��jN�y�\ �۷���z(5�7ɓy�ODϮ���R��!6��"rE���y�>^���m�@����;�$5�Qf8C��x�(2��,0�\p76�$m�p���j��b�=�p�E���'9�>^���m�@�����G"����n��J�
B)J���w�oz��������_ �SG���ND�h���@����>^ݳ�|�k��m�@��P�?H��M�E�>Wv΁����n���y�\�z�#���2w�������3<���mt������)���x9�e��ͶHۑz{v�uzh�gH'U{N��[.zMĆ箋���t�)��XC�J� fM`���uF6Z�ԙ:��L*�Wmu�,��\9;������twdv�u�s͎N���As����Q�u��C��Ϙ͂���.��0����v�Q���3��X1�Q��1u��c�Md�X��d�ɓ]��q��4z��]�h�Η^��ߞ�������K��s�t�����|]�y��qutu�y���a�z��$�n���>���vz[]��:�9��>@f������6(��L�MU��������<��@��wz������TL�\�U*���[�j�<��M�o7n�k7_ ﭩ�����5��󓓠�g �����k�+v΁�KȔ�'���D�����W�|�n��<���7�������1�hq���%3úWd�t��W=��	���;C�\� �R�~�`�s�W�|�n��<���7���B�b$i4�1BH�����:�� &,�E��Qv��I]��wn��^����V8byQ���9�t�l�ݷ�W�| �wo:���iFd�9�}o��`5������`x�g���h��ci�N��p�ݼ����/1��6#3u$D����IJ�eNԬN��p�"hK�nL�z�q����0,��S���@=m��@=v���{�7���;vԞ&�$o#2>���l�t}�݁���@>���ݕ6$ذ�(���' ��oz�[�\:;���٩+�2i�=�h��D��AQu��cV���j`Zp��>3xM��c��1�'�	#[��vh3�5+�u�KRӖ��h�L"1)�mf9*L�Wy��ˢ��8�c��X�deV�FNa�Fc��6f�0{@���DCF��^v����H)������1� ( �G�=���k��k��O %5vz[] ��l'�z�����sQx�H4�h��R. }뷝��|�m���j�|T�*X��,�@��r"k��/����y�9�n�[y�qr;�u�<"qE#�'�B5;�s��@�_ �������-�o{`�3@TTME@��z}���rN���_�:�p��-m��H���'{��N�����y㮁��w`zS	�*��R��]�D%�{`b��\��|�@�PIa�"�S�*:��1x�=���^{�f�4NF��G;'9�<���=���W�| �n�t�TY�c���rȫ�:P�
7gu�p�['nE7i�>=�:̅-ODB���{�W�| ��y�<���7�5�#Ē��C���5����큫^�@��w{�r#�pѽB&�R�S�U.�fn�l�9��Y��vY�=>ŉӆ'�B51N���@�_ �����k��m�@>��aq�&9��|޶��o��������|�������?����d�F��z����^��0�^�u\���4u6�ueC��GY�b19Z��żv��ȯ�9ω6ә�l��h!�*e��,��gN{n�E�.��C���]k���Dz"����ۤ󓴸lV1�f��G+����=v�Y���n����YF���X�fٹEk�t��ѕqe����	F5�H*Ľ�)z)d��7��>��0 ;7�]k3:͙���ݭ�S���ε�����S#�qmṽ��pֳb��UAJ�(���Dʉ�������;y�<���=�oz��ˏƛ���� =wo:����m�@��_ �ݲ@s#Pk$�Rs���|��ށ�־ _m���eom���!B�5=�r8���Y�=�)��<���-�k�G�
a���@��_ ��j�Wk��oz����d��;e.���I�0m�( ��)u�.^� Wn�k��n֐�rjQ���͚��?e6�O��n����DA�DzB���}U_���F�)���@�>��s�S�>t�� m�i�C�����c����ڰ������1̘'#��oz������{6�U�ֽ��Fd�P�J����5Wa��r!9׳�7n��=�-�@�]�q�SS��#���΁��|�m�@��_ ���.68мOAۺ�%�P���a�s涞}F�}Oo���Ckv �8ҒL����A���9�t+���W�| ��y�/���4�E)!B�5=���G9	f��q����x�Ȉ�q#w#t���LM!R$�������7�7�� ��dc�M)R�QDL�DP�TE3A0WE~0��w�\�ϼ������I&)�1Q4UT�6"�{��1k���������)�pH��)�w$�:�����ށ�־ _m���Ib��A�(�$4�%����W;7���s����e��=M�0���i��1̘'#��oz�Z�}���g ����13�ck�����DDDBA����3^�@~m��DG!##]hL%P�W*�U5US�׻� ��]6!'��vY�=���$L*����5g{���b�{]��݁���r��4�W�CE�u�}�|���&��7�!di��=�oz�Z��[y�]��{=�nu���n ��d�i:�En�CڜݮOb�0PMNSV��ڟ����,Is��_����q��y�}�������db)$���x�C�H���|���o����)�7�Ѱ�?L�DN�|��@>m�@�6�͎G9��u�@37w����y1(�<s&$�޶��n�3��o�Ȏr���@�ѯf
��)��ʉ���32��6#�3w{��v��ۻ67����=i(+�&i*�j֌�v���h��}���{��l��9޳��:����n�fn����\�nɱ*lmR��`�K�J.n{e�wHK=�؞3lA��aīn������qc�71�M��&Y�����XV�;1Y.��U��U�=�+���q��>u��&͸9�xq��jۺ�㝎�sf�N�ۮ�b4-Ԗ"����n ���~{�������ew=��Gk2�̓.cѸ{-N�v-��P����3l�Fu��9����������u�3ͻ��|��Zt�n�0UT�D��Vv{��ͺ��ć��v� ��y�-�.	��F�D,�98��ށ��� ��fs�[g �sr�����Т��@��N z�����7����5p��x�C�8p��΀}m��m�@��N�e��Q�, ���yS#j��5[=fk�c��!^�]�����j�;���ϴ̍DNc|��@�[_ �m���)���΀o�el�)!2B`���]��wʓ�!+fI)r{�� {7ޫ�=�Ds��H�=v`���R��*U]�ۭ: �o�ɷ=����8��@D� �c���o:��p���؈�Bm�N���va"aUT�H�*��]�|ۮ���3)� ���;��w����a����(
�kt%�G2��`o.
g���P�\�n��QɗO)H�
*T�Xwv�̦to�>@z� ��ZF�����nw�y{ ffgl��t�w`f"RW	����BH�m�� ��8w����B�2�iBR{��݁����3��1�rL�DN��rt�l��{�7vS�Um���ƫs��HLJj��6ۻy�s���t�5n�Հ}m�n����L�Ŋ���Gƍ��X�0t�l]W%�l�;����u�3�n��N��䚟�X����)�*�l����.�{�=G��!�R!�p
��V�n�����L��H��[ȑU4�I���{ڰn�t���7vS�U���-�����DҀ�E5=�n�̦t��V�G">��N�S��v�p���k����_w���kP��L�Q�;�=�)�*�l�-�����
�PB��Fҏ����J'���������9�읶9�c���N���S	����d�.V�g@�m��<m��G">A�^���������:�I��>[k�m��׵p
��:}q���Q�|����V�g@�m��w>˵�6�S�k�����V�g@�m��]���z��SLd�AI�H�Z۫��@xۻ�8�@��\Gc��@�=45K��ހ4�0���0�#�m�@���#��������@: 0�������X�uf�ʎ�
�88.�Fx _DEl]������w�3�r�#�}�y��w��<��0�&���1���%r�S1E<4�j�*��L��,"(����a�9ތke�L�IDI�Fe��bPa���Fj���f1f=o���{�}�~��V��6���qoK�Y�q�[7fc#J˚u\�) ��'CHF�C�F\�Or��nާt���9��z�.���Yy�S�3����E�_o��#"�Yw7\��=���1ײ�\�ٝ�pf6��-۰��z�qǣa8)�c���k>1�c6��yݐLgK��0���Єl5nM���Y9��HdyZ&ٞ5J��vT��Uًb��;�1[E��v �6�[y�HyR��۴�/;���Y�$���wa��72=�͐*��p�
�щVba�r�T��f� mmB��F�S��4��i��m[ �a!�/Zl��f��0�n��Ae� ����o����$k��k ����`�V@4�d8�A孚�d�ю��&�6]`&��֌i�����4��R�YW�Y[i N�r��͸�%ZWvz���@��۪�(ղ�hDn���8��[m�.@-��%]7��G=��8m˥�҆��d^x.��m�͜t�l��L� �{�?>��;c/<�G����{���ż��-g8e��o.��T����&�Ckg�y��:.Ll�O=
i�4��E-p�iݍpm/ԍI��-�u��lh;V͹,�[ƪy�T|)���=Q��#����'f.v��SqWa=Ǥ��tuX�:P��gI,���ץ�i,�����75+Y�6ܙ�6:'�*hj��gg��� ���V�]�PMm���<��ev�U�mKP�tɵQ�J��ԅ+\���&v#��0�@]@�mU�����۫9yUV�wCd��귎�|��͌u��ݘ-J�h���x�c*i���J�u�U���y��l�Ɍ��;+l*�摜n���Y����豪UL�j�Ttk�]�r<[3�@�&��w(l�vl��vPZ҃P�gH�&��Md��z�$�)�����|v��	<���*���I]}]%q^��YwA��w��/3.t��Z%��]&[p�v̀ ��h5�7]Z��H���<�}��{��W�'���=!����*��6���W�
y˫��^�-�l�5u6�l�\�9l�%��C��ok��gtvۣu6���(�iv��[@���h�B��;[@6����*�R��[+�nwd�3;'8�L��"9����֌�5�\���v۷W�h�3b����¦Fv稍0��+Ӷ��Ct�����u{=���(���p Y��\�=������0�C�g����r��)�m��͞�w~�0|����f�e�b]�ۏN� �4c{VY��j���vܛ)r jt< ����������p�oz��\��g@�o46?�4�/�8�۷���\��g@�Kk��#�H�{:�J*�E!J&fj�r�t���[]��v�E��1
4(�I �n��>���.ݽ��j�o��r��G'9:�ڸ۷�u�\��g@��ߑ��b�z�.������c�?]��y���Wf7#���HӤ�M�Lm�M�2@�&j���^݁�8�@ku`|�@Z����D�;����7�|V3'� ����xz�w��k}y����5�6��!#4��U�UB��5G@��v��[]�n�fS:mT�5��'��rtϵڸ���̦t6"#�[/wj�{�#�d�ȚP(�|�۲���΁��_ ���F���FLcibdJ��CD�3n3�=�d|;n=<��>�΢LD���G��m�ށ��NVݳ�|��؈���A�^݀yÅ��I\U(U%Tt��W��Ds��廳�5����)�>�j�c��&)�rNN��m�@xۻ+y�"�9Tܽ]W��VUkM7qH�		�9' �m�@�{W �n�����}�]ȓ�'?$�UU���t�����ۻ]��ށ�Z�8�q��?6��i��OX
�N2�t�fM�'��[�.6��݄�t�d�Hd��. {}�� ��8�v��{^��.�ƚI��dƱt��@>��g���ƺ�����ظ���DҀ�4���oz��\ ��y����>�U���Ȱm$ۛ�7�����z�;ޚ	I�4�2Qk���ۗ��!:J��D��T��"��o:��8��������~���w8F�n���+gC��u�����[@����}��v7&:�	���[�9��'9΀}���m�@�������U[�6�GP���p����~Čr�t�{� �������eL�(S\IB���32��-fc�7����[��=G�#��?AH�!�:�v΀}m���{�7vS�m��ǉ�ӑ��.��N�}m���{�7vR����M�lړ$�xw��KôWc̬Tz0�E�*�qJcZ�ף<f8#tJ�#C���,;l���L�����B�X���U/\dw��݆v9��;Q�	'8;tv��'@��$��ƍ�Vv�FĻ<��:�༡��xN{WF��ԻWi�A7�s���~�[0t`ۧv����7[�UVۃn��쵤�=[�xz��ݍN����Ǎ��o�幮�^���M�;u�l���)F�m�ώA�ϟjN�UB�D���@�R���n���L��1Ձ�m�C�8��NQ�M
y42�f���Zwb#����7�`�����w�H<������*��(���>X�Հ|ۮ�~�w`fN5�>����b$}C|�����;����L�o"#�I������Iʐ�RbNI�>���l� 7v�t�g �}�kI��Om���K"��M���X�|��8n��pm�=�.3��e5V�~Ib�w�[e8����8�m�@�6\��0jC ����m�{��<�[,��m�@��p��68R�3UJT+��� �u�>x�ټ��B[�Zt��큙�GdPR��H�98�m�@��p}��Um|�Օ�q��dCm(��@�e8���Bׯ{�����7v����2Vz�g8ƻ%=���u�m�-�d���n�����NzDV���{<��a�m��7��nzͷv�L�{��J��*fP���]�{`j{��>m��]���o:����Ƣ�"&b��{޻���d�I�+�*@!�JX�BB$�I����!-� s�ݷ��m|�f�U:�	?$�T������o���t7�^�����;��&9�
@R ��y�*�_ ��{�7l� �����Ӆu��p����ϵ#��.�մt�Fӽ���5=z�/C�$�I��7$Mb��9�<���}m���S��o:�x�x�J&��T��6���HokN�6�{`z�W ���.Lq��"6�rw�n� 7v�t��p�����Ȇ�URS0*B���Cy�G!&��l[�=�����I��dDc��~!s��r"�7��a���EE*�R*��]�{`|�s�>m��3'�f7�6�;�����j��x^R����O% ��#��m��@��\��j�L��ٶ`r`���}���u�\ ��o:�����Ĳ�Z�OͬnN�k�p��}�<���6���9�$f���QP
�"��U4� �����@��w�=���>�j6:�#��]8��t��t���8�Cc�ȈI����ke��J�%@��MW@��w`n:z�����>��z9�Dr��Ϳ;�p8jZ�d�6�Vz"ټrΈ�r���wh�[3�GE��N��l��ʪ�q�DΣ�^x��LѺ�)�c�>8wF�v3�{l�� nyMq:؂y�*���37����	��Z�G�6�ێ��B��C%���c�[�H��ܽ Uc(_�����e̴�v�F%��1�k[�'��rސ:,^s�v�zme77��տ]ߜ��n���=��bۚ�a��N�wT(1M�.n��7�P�ӧ��y��fz�����>s���c}�y�������p�ĎH�x(�6��[o:�[8�oz��p|{J��DDHt'9�����m���n� �m��UV�ǈyC�rN��ށ���U�΀_[8�ˋWRQ�cnw�_=��j����cm݁Q���es��ؚ��R�8r��k3����=�h��l��[;�M`����FpM3�NH��������8�w��=��=�j6��Ğ%uS`o�����$�&dئH���`{���n�a#rwTĮ$�T(EM.��wn��Kk�bm��<���kwE?(�MG'z�ڸ��΁����m�@>���Um&�Q�T�&۫y�����݀��= ��Wq�2DEY��ƚT����&I�V�ǁ8��痷=�YӍ��ظ�GB{�Հ��]n��9�@���X�A;R�
�D�D��]n�
���5[l����_�P���J!�cnw�Uv���gO{Ǳf!Z��)
=V�	sh���X�S-0�%(YF�46�q�5��qFDw"}�$�)
 9��L�b��
�V1QA\��7�L��A6��a �h��T��Jbh5g]�k6{���6pz$8r+I�̬q���İ:��J&A�"
(h*"(���&��I�.ME�:��E%P4���N�&����(J����J
�,�)�M^�BR���"��"��
b�
��j�sDLj��	��/X����-�V�I��ƽri���
�y vQ8��aˣ��*���)ih�0<7v�N�h�Y�[�MEICMSE8CAKV�&��1D�Ny���I�FR�Z5���'�;x��aX�'GAh!��N�.��1t���b���8vu���[�J���4�� ���.v�'roFf��6k7���К:��h7���$2h)4�*w�Ă�l9�S��q���Z%����W��L�#�S�0�@����5��oI�iE�TS�
ͧ[q��M ���:�;���0K��\�w�u�T
(Ԁ`�:��(�s�,�#xg����h�*��A(�Fԛ��B�)$�Nw�5�E�^��'ڽ�]��`+"�����@q�õ �޽��p����{F��U��ٌR)5S�16�X�5�1���b"ν��P6�5	�gx���-{W �6��i㞁卺�?W�<j[3�L��qͩC�mn�ƭא��K��Ժ��G=[���\����O8��&?[o���v��9�Xۯ�DG����3ٟ��<��Q��NN�Wk���:�ƺ�n�b7�BIL��3U=���`c�k�y������@�ht23	��9:׵p[~몽���r�Cv�����i��!v绵`jj�ڕ*
��j���]�n��t��V��]b9ǘ��Un;�sO�7M�4a��8��E9�s�]��;;���WY��ɎX��-�t�k�y��@ku`y�5��^�݁�	�Q�h"d�R��:Y���r#�Č�z���݁�t΀�1		8���gy���=^��/����j�m�t�^,(<2$�LX�q�?�k�߬���X۫�㞁�ˆH���i���@�;W ն��<�9�m��+��{�G"#���I�m�������������5�-��a���BY�!]�wZ�u�$:��҇�]�@i�4hK[b�,C\l�6Ht�Z�=n4�;85 8���]�*[=�.5����m�֭��㶗o/��n�G3� AK��8W9��Ƴ�uGc�3͞,�ς��K7X��¼k��0�
�f�Kb��-�a��ȗh��Qz74�vJ�����j{����������?@~�`Wm1�h�}����b���8��:^�m;�hnѧh�^Kj���>_n�XO�6��G�N���4R���I
������`y<s�<�w`g�3�b��^�$j������Q5P)������`g�3�b��XWk���,V���0F�z��p[m���|��$��&b�I �m��j�_ �m�@�v��䐅�H����o����v�Iю8�/EΫa��{VY�4�1�.ۑ̓&�$P��w���U���oz׵p
��:}^,K*?A#&,�r��n�� 9DG9�]	��]7g@-�8�U���Ɵ�"i���@n[]6��n��n���ڃI7�@�ȸ��΀[�p[oz�j���O��?)]�NNՀ7����v����6���G~~w���ڲ��OGL���N�kx�%#��n]t����Nnӹ��)�����uD�B����{���v�t,mՀ<�8�pV���PX�G;�/�� ��l�ݳ�{m���Q�+��QBR��]�u`1�E��9�q�DDF�ܞG9d��݁���@~q��:9$i����m��oz�)�*�_ 7�<Y�,Ȱ&,��t�n���9S�`j�s��et7���ٰq��:y
%f,� 8)�ն��b���g�'FGûc����ݫ:�
�)�2&����[��
����vpݷ� �б��F���6�|�u��̮�������ش�l�Kj��U7IW{6�ݮ��������m��:�����&ɎLM�8�o�uWy�k�}���^*��(�"	�A:P]�.���^zU�^���Ɏ#s��{W �n� w���>�n��DDs1�H�S554���"I�Cb\�v�ΉN^9J��tF���v�ͪ]�.wg:D�)0��)�.�U�����p�5��#� 󗫠6��S��***^<�} �v����kڸ뺹���"8�}�@�EP�3S�{�`}��t�Kvu����s�>��M*��c��M1I;�>׵p]��:��|wm�@>�6�J6�'�����z �����5��7�jC7��{�{�v]��7eh%���GQ�b�b�����j�vݶ��g�x;���z�\�re�g��B��*v�ݕ2;R� �zݝ���b-�Q��Q켣\�vu<�$���wn��I�:�z�{np͸�A�۰u��Tw\�zP�r�)l�:6�F�rj�$;��t��F/�A����ӕ)����LtGY��v�&v�ju��n�[m	k�q��Η~��@�/F��=f���kVk{�Y�[6yA)�O[��%��q�CЉ��{�c���(5EIQ5�EQ�J�ٰ1{vz{��2�V�|�凞��16Lrcm��>�n�,�=<��kٓ�3��ڔ�c�f�ށ�_ շ_ ������ށ�X�U&�(�R(�|�y=׽��3���d�]�`7c�!�ow�>��ݯ�_[{�>׵p/n���۔˒d�'�!��q�������[�����]�˻y���Vt�f�TȢ
�r�jl׻v�8�@����:��|�m����"i��n�Ύ��-�7:R�2N�OE��π_[{����	�$m'���^�|����/���kڸ�U�E1�s��!֔�@�n��/���kڸ��_ ��a�$��D�&6�|��v�q�������2�������h)��-����t�k���ss�;�;.�G��Y���m�PV�w�߫�8�@��d���]�n���,���y�(������n�n�ށ�_ �j�A�$��#x�rl�n�x��<ȉ��3�t_f� w�4f��~ A�8�oz�v��ۯ�u{��֭�88��M����-���n�����/�w`o9��lͩ����TJ!JT@2w$��
�q�B:^�8�.���Y�K����8�#M�m��5m��u{u��[{�=�j��V�	��~X�:�}�����#u�݁�֝=9��Z�a�O�4Lp��q��oz�e8��W ;���7��S��@g�x��7�|P���{�4��:��4j	�E	��No��]UZ�#@�iHp��\ ｳ�[���}��UJ��&$�kyڒ�.��)W��H�]�є��<��R������Cr9"F��닠{l��n�����h��@>y(�D�P
(�����"3i�Kk��l�U����M�����py� w���/����7�(Glp1�3�y{u��n�}m�@�����v��~L��Js��[g@[����x����}�O@���$�?�ȄUU�� �������)��A�w3���`
(a*�rEC?�b
&L�����̒d�������O����?W���m�����������������PEU_��������2����UV��?�����������C�H"����o��?��o��O���_�o����ԡuQ�~����$�d
$��@@)�P
P�P�D��"�@)$�$�)2�L(�B�2�D�*$�L*
�0�K*$J�B��R�D��
$� P
P�D(��J2�J	
$(ʉB�
C*$�D��� *$"��J�*$ B�(�*$$���
@B� B�(�H,��)*$��
$�����$���HB�� �*@@�! �!�BB
� ��� ��2��� �HH)! $�0��2 �"� �@@(�@! ���@��� J�H���2H@@@@K!�$�@�H�H@I!)B�H��	(�H��@����!*�!((! B@�2��!*(�H HB
��
 BJ!�H@HL�H� �!HHL!+,$�	!,���@�
� J��H� H����(��B@ H�!"�!"2�!+!) B��) H�J0�"��!(HJ�� D!@L�� L!����P D*� ��%U2@��%!	� �!�%� �& ��Rd
@�!V� H�b��)!d �Q%!T�I�	�	Q%%D�L��g�o�3�"����N�����?��W�"����?˘��I�����c_��UU��?�����f�UW�AU������������UW�5������3:?��l�뗼�]p��UU�O���AU���2>/��7��~1UU�;��UW�.�����>�ޗ�sqE���+�2L�������<��`v�g��w��UW����A������O���������e5��s��}� �s2}pI�" � ��@c`��UZ�Z2h=  E��J� f�/JR"�(!UJ��(*B(�� U  �J@P
��(HU U@QH �$
 �J�A@R    ,$ 
�T(0 ����u����s��uŜm� N�nl����gfrܶ\�J�} �TŽb��k�išٹ�� ST��ca�Û;�s9{�<x Q�W\��y��}�>�u�g=<�
��  �J @��������@��l�PX�(��R�o@ ��JceJ(,f��Y�)J0 �(,f����� ��`�(�Ҕ h�� M��
&�R��t�)e��1�
lhM� w*B�� �@   ��&�R���mO}�/���V j��O{&p���v׭�ަ� z{���ލ��  �q�齞N�w  ����om�YWo���|;y����@����ZU�ξ^�L��yr��  ��H�
� A���:鸷jۋ�_Oם� yKuϽ�������ʦ]�W ��A�o��ys��ye{��oq�p>�^yS/}�t��<��.:��6^�� ;���m�;��W�}��[���x�@A@�@&X zS'�i�;��������v�����ۘ�w'_-9yv��^�� 'Jd�מ;��  7�뷛��].@�F/vS��z��{��{��@��O��O&�n,994�x     zB�)P  "���*��   ���R��@� "{JI�%   ���j�*� �)���N"t����G�������̝�t{��������.��U\� 
���"*���U�
��� S��?�$� S�¬k��#!�$+��02� W�D�1�@(@*F�0h��`A�DM	(B���7qi�e`�Zw* �T�_W��@CC���S>��fԹ�g��y4N+P'*�J0���7?�A8�H,b�<e�XT`Ri�Xc��
��q4�4��	b�m-��y��n�2��XHQ�9x��c5�T�!˽���'��;bB}����ė	a�AR� ��'w�}�}�6� ��e �ѤR�i�LAH�>�LFB�2�:	LSHHjaMB��$7j�EҸ�Z�)�����.\�(fƄ)
�H2��%�L0�%0B(E��c,.$(B�X��s�jjb��BH�U���l�@*`��ԅB0�0�
��aX��æ��Ìѭ]�g%���`%!!YvCw��3��0�*���e�I�[�#/+����#h����Mh&g�����Z5�ωq� I 4
a#q���^b�m�e"Д�j`Ȑ��y��s털U�Da��8��>3�0$������5.s�� T�A�~�0_[q�p���Lb�|ɜ�Ro2�d�0�R+`i�L�W�K��<���������0��0!� ��\�����q��:9�.�6�i `1~e�j���
l�!Ih��!J�L�L��@�nCp
�2&�"U`E�"�g��3���.JcT%︝��um�����F�������]�h��"!BS���3�o���~I�I��2����*�����H1�fT�n��ɦ�
��*I*G��+j���R��þ����W9V�U{��L�oa���\�a�ˀ���L
g���e,$	�I�ّ�LS�p��_�M9J�w�X8�W���a�C���	+�>p�qs�T�R	�BA$�"�$�H�IE�l���B��`@�H�`Bvs?}�JbC�@�Jʆ��W#�5�$>Ʃ�Ή����rA$a�N�2����p��y,�Xe1�ep�!dH\h�d�R�<���5��.��k���1A����O�����@�(�s�o9���	
r�����J)D���x�f{f�{�d�ּ��JcA�._��.BM��,��FL����VR���	R���	RD�����rh��5�����H�-��d� 
�Z��#��`�p�. \V+��a@��h�t� ��:4"VKF�j��������*"k)K�?)�?+i�*ߤs(�~$"R�����}mP���$ҩT�����?ZW�@���^Е���r�����m��vU����Q�i�]Q��,�.1󫹯�c�Z�_�ۃ�B,a!H����s'>�d56he��t]�y8ƛ3  E����4h�Hh�D�ѻ��M	�@��� @� )
��J��Юv$�z�����_R���C�+=4��2FB�*��+��H���	$)��0"�"VD���&3Ґ�%3�$��B�+�!:�o��p��NЛ��ŊUyc*��u�v��1�S&;1(�4�	4���`w�����1M�>����Z�+P��z M(��$~���HX��#�B1�B0!XQ$� D�*�bM_�`�Jr���~����Y4�q���Ħ����/u�u�*B�'s���"!�U|��{�n��:ܹݳpŲ���!q$���Tr�Bƒ䘗L�RB ��@c�@i���$�m��0��2\F�zO�3�q�����0���a��H$�����'~� @���RF����ʧ�[��aEod
��m*��������j` F)B-�d
ih�2T U��V�z���n'���`Q!u��^o3Ә�I슖%�}����z�j��U��{ٟX3�o��w�ޝ��4�!BXm$51��X�	�#�	f0V��`4`fI M��;��2�$)����ה�JaL�0@�2@�0�L5
��F�HAV�%�1��l�� @��c�0R�a�51��0$*X��� ��V\f&��aB%��1����vS:���d#q�M���H��#���UU���G����W��u}Gwu5ͽ�vտ;w]x��ӹ���yt�]ﺏ�1�����|}���m�'�>9��j`S0L���b�r�R�P(�F���$  �"".�� ��R(�Y�%	P�0�B�@�E#��G��{���]x�׫ʙ���]g�g���[[�f�B����.��I��W�|^����r�$�5g��Sdi���8��	�F���R\�d#�������C�"T<�JJCI�C�T�$��aɒ����Ȍ�4 �&s�����f%�֓D���c��bF2b�	p�X!%�y�J�&������,��"b �NJ盙�i |c[�&V!V%gw�d �)��!����@CZ{���3��L�y���Ĺ��}��-�D&�5��٫��'�5Ԕ.����\d���k=M���I'E��;e�ć��4��
A��K��Z-�g�˩_��B$ĄL��3ݹ�>�y�5�G�,�ۗ���Ґ��i�$f��uu�\���3��ڲ�r�B󟷫�ʪ�ꪶ4�7��A� �$0��Nc��d��z�w�!7� קFH�q�n_��=�v7��g��C�g����!;!B;��$b�$*H��Iw�l����͙�~!�A������`�e�
�0����XS)#Ӑ�Fc$'��!D��F���M.3�E`) ���BE"	"Ā��b4� ��`�e��s���U����H�SX�a!�@�,@��(LZ䚘�Y@�B�c$P� �a�WB\��s�d! �!!,��a0R	RHP �!I"�"�Xєѣ&�}��ܽ�ш@��"`�Q�,,��0�Al����>_�}w�Зr��|s��)�P�*��!
8X����ɭ��́����!)�w[���٬�	A$Z�*2����~H�b�rr}�LB�vHjBՠ��HV�	�5��Ե� ��E���>���)9x��bD8���_��~z$j��S����h!B\��.2��22�b���$����1���m�y7`ޥwt��.�^9�%�.!�"IG��$bĈB�)>�!`XY�F�9#��)�"`$�#$���bȖp�,i)�B�&�k�����p�u&d�2�+ï���0V$# 0��u��'Nu�ͥ�G[�
�4�E
}y�PW�*/�U�)J��I��`@#3���~頁C�r5�A+ ��(�$0�DY�7����S.k0�};fqL�	�He!L�)�9,�	��J�"i "k���� ������c�15�`M�d9	��\X`��u�|Є��0��)�yl(W�+=�.�r]E�i	�,������60��^X�
��F�H���HnY��7>����.uV�z����|@��HT�9�!�\Q)�1�������e<Y!B<!tF�1��gP�J`2I	.>Ʋ�����>�m��zHR�J�H?�CF�$�SXu�s렌~��
c�5�+�bc�"�R��:�C����{����
!�D1CD
kʤr��ju|3]z��ya7j�S_E�J`#�D"�RHB	$#L1+�:��a%`eWrG@F�)�7)�ˌ�HR�aX�"%��>�Lg�1���B2��A`X�cT�R4$`��@��2sz����Ⱝ*�ŷO:{׋Ծ����R�����s�WQgZ�)é��n���S����ь��+B�'
J��������x�q��p�K0�(c���7츁R�2B2�rh#L4�� WM$)��A�����B�s#$(`"!�� S�
Ct�4��D���.2F0)���\g{>>e�ɤ"S	
&#q0
0�!1k�j1��уH�k�F5�˩q�D $Ě(*ӵQa�y}1�%R{�UQ�   p [@ � [I     z� l m  ������ؿ|��]68���i3U`8 m[6�u�jv�n��nm��0 �tUJ��l�ef Wn�ά6�����e�6ط�� 	f�v� Vԝ ���[qmp[vȽ)$�\tI.��W��[��SVQ��Gg���t  �j�m�o[@���   ���	$m��-�K�Z���Z��Wf�U�W �kF��![�V� ����R[�&uI֫�	UZ�e�"�n�'D���T%�2�*ҳ�ڪ��H'�l,�T;e�I���Il�m $n����Pe��i�i6-�X` 6��[�մ���(ժ�U�Hm�    ��:&�&p6��      � m� �    m� [[l��ۀ:˩5     u��l�n3��� \�m�[�첚��.��MR���UU ^��#m��j���f�` ��`� l�P�`��N.��0�,`�3v�S   ����O�~���V��e��K��m/l����*t[�y��ڥ���i)WfV\[��[T9i�T�-*�m��ɀkZ@[@	�`llv�*ڦ�<F�r�LPpv�[%�m6`*�"���%Z��U�Ub�m��ۆ�-�M���P���M�: 6$&��V]�� j]�,�bI�V�� kR�W�; ڔ���[UJ��j��r��-��BAín�mE',
�V�U�˳����J����� ��8,L��A
��u�nx���&��zJ@�@ �`-�  ���u�J�*�
�TTW8  ��f�ڛ\j�v h�l  A�       	  m��� �|�@�6�ٖԘh6 p��k]���8�m�f� 6���ۤn��$ In�U۱�w,�5�Us:�Ug�y���k�r`�Lg���{p�S�(���ӤZ���rn����)�\8Ԫ�������s�y?�Y���\d����R%�h�{7���+T�QnE�N
�����xj\s ��Rvy�Om�)[�4��ՒYĲ����ג�uGF҄�yUt��:��f�1m$��n��:Ȟ�H�k^�:��[��5*֭�b]u���jtLs�m���tp���T1�'E	��ԇ[�ݺ6(jBj�MJ��<�u4	�� $jM�K5�RΛM,� ���F(U���h����˙ ,2��@ �\ ��Y���-���-q�l3k����H2�Ͷnݘ`2�sc
��U����5��Vą� m�   :�ְ �y�#g���W�[[uC02��p�w&H�L��۶kz]K+ 6��-�6��M��@m�`h-�y��K�/�6�&�m�;i+fݳ��j���Am[[Rѓ�X��k�i���yņq6��Qm�` � -�i����/P*�P�@�d6/.�]��8 �[�� ���i�i.Ůu�@[@ n�4� 	1��   ya�� [E��A� 9n�R�����go-]\���[b�]��h��:Cl�$    H��  �i �M�%�� k۲F����K)�l     (m�|m�6��lR���N�A�    M���-��   �m�   m�mm�Ę�l -�Ym�i0 � m�@   v�[OZI&ͶH�&ݘ[o m� m�h@ H l ������NȠ���`	��IX $*�%5+�O+���U�� m�� m�   ��v�[@�A� ����M���p�#PI!zJ��������>�|��[ �> &� -�Z�L6K 6Mv@   M�Mm�m�j�D����    �6ؐ$   K( ��� ��$�M���	 �~��6�0�m�[@� �8   ���� 6� �bIn� H  ��Y��·:WU[Pv�Ĳ�MPm�� �l	<6�   6�76m���N�5i�ѵl ]5�@   p	+�U����,�K���� -�m'[�� �!6�ڶ  m�ga�n(���j+`r�Kj�  tp8I �l  m�l�,���������dH�۲�Iz޷{r��h0	oX ��k� H6�5�n��m����p�ۛm�2u�F����h"���*�iv@�@�  �k�.؃l���p t�dH�m� ޽n��*G-���h �9n��p m4I%�ְ[N��'o���pK([4�Z�$kj�P���H��Q�/5Ti�t���l� m�Fհ �l��r�� -��h	Ӏm�      �i�km�t�['�M��t�|�         �6��[�-�E��Z���}���rG s��z���$�h��ۻ�J�S�m��J�m� 2�&֪%CX
� �n�Br�F�T�~U�|�P�z��@'UX 5*������>���ls�Еv��W��eA^�Ʒn#�cnm�4�-�x���7h�a���u-S���ڛD�UR�^���U@e���Mh�$CHf�`�I��b�t^�t�[r�,��c�`<e������u��9�Snl�
���,ѣ4��qՔl�iM�=����c8�8ZԄg19�Kg]o,k@p��A$���t�u�MA��m��)��n��@�6n��s��z2 �j�tZ5I��.9�<� b��g|?t<��\"�UUZ�0"(�&�2E�m�9,��`�)*��iz��\V�9u�1F�H��m:�k��Z{<����Uu��讃��4�Q��Y��\�8
R���ms��豢�#���  ��0  p [4Ņ��V�+��:����lUVҽ�C��3��[mr��vx<���Qg��uT�p�if�Kl�:n�g�V�HH&� = qκl 6���Wf�"C�M����N���m��`��^6�U���ށ�)V�tHl;.x�k[s�����mā���;i6$��\Q7@u�� ؍�9���-��S�i6�f�Yg�Q�Dy�kl��]�[��n�3�v��m�,+үz�]��v��+[;R�//+W<��^B�bs:�Px��j����g���[qm�k9����wn�P�F��!"f��#j�`���C��j�)?$}��:�'�emRΉ]��u���]��Jn��@�B@�`k��n���	*AnU��Yp�u�PV�mT�����,?K����nIl	���	-/66�(8 �ln�   ��m    �.�z-�  �Ziq��M��kN� E���o6olְ $�  [-�5�n ��$t�l i&�J�p �l� -��l�Z�m�Jmsm�n�p��[E�׭R��m�F�<��	�Āiͼ3E�.��J�-��Y�,� m��F�l4U����I�K!���� z��`�
����`%W�J�Jv���gi��l�M���A���&�t�2A۶)����v�S	%���sm�ֶ���m�9�l��h��4]kHYƐ�f�8A':�Kh�(R�5A�U@Um*��! �*�T�l�[T���Ŝ� ���Ŵ��m&Ͷ�`�SH�`6ݛml�@    8<�I  [IV͖�KZ��"�` ���.̇]U�!Z9n��z2ĸ�`�����u�ݓ�ڢ9F� 4Q�ܽ�]n��-���9� 8��,P���C뭣n�[@2� mp�`�`�����>��)�� !�6��X���kN[@ m�K$,�lv�,3+mU�g�k��]�s˘�Z�T�r��7%�q\Z���F@I�kR���!m�l� [r3Ӝ�&� 8m�d��nx		�����W`9$�H 6^5��Wl���UJ�@R���T��8�U���0Ă@ޓ��l��h7b����j�9V��,6�  H�[B�dHk� :M�m�m�Y�pnB�P妘m�k�ە�;U��2�Uv�*�U\�.M�Uj�Y�V��M�NKҭ�gJ��t����-��u+;��[�*�
��4(ޮ��L�����W	����i��Y}�����0��e�����2���Ȯ�iz�N�غI��[����lԍ�v�V��1�-�t�q�=nW���@u´::�Ux;z��Lw�-.�c�Ks8���f�-Z��
G=U�`�ٞ)ͱG]S�'T�[s���U/<҄`9���H���v�8��v�GvҨv�jC�X*�좂S���ʼ�tuu�J�$�Ҡ�m���v��9m�h[d$H�� m�l     �p �h     �m ���}��!�g�� �g
��P��B��U�A�U�\  ��UbEUr��vDwD)Dt�(�@ºh")��4�P��S��@�.���e��ѱM &��ʢn�@��($P $ Ab�b�"�B @B$E�z�e:���/��UN Q*�����t l: :��E�!�*:D���!��D6	 �D$ "CKCj�t�&���qQ���~����v�>�d ����@4@�F�� 	�QȊl�":x:�lS�]©�W ?lC.��	 ���`�0t��(?
���J	�6,P���F(��/¨u����*qT8�8��@��G�b�D��Sj�TH�DP�b�j���rdQ>AO��XAZ*aG
H �bĒ"0"�ʇD2�ܠΈ��(�/J�� A`1"@R$1!> ~�0@a0�G�z�2��#��`�����b�F��D(���5DEWj<�H
���4����DŨX
�+�#����`�D����'t����w�w��8q�l$n�/@�6����6�Vw��:k*<֭�s�$J]/d��s�	�A0cvѺ�4� u�ny��lҫVR�6` �$�kd�ֵm�m�5���]�4�'l�Q���mrc-�Ph�gs���U�9�P��&y�c�  � HM���ݎ[�uƭ�Oz�9R�/�v��֓*̀W`f�Ԫ��J���Rk\6��v�o<�s<�n%�"-&܋�5ZMV@̘e���N�l��g��Y��kZ�\v�t��['1�)m����"(�]ێ����5UP����a9�����Q3�z�6���Ī�kv��r<��n��8l9�R]�ͶF��.�^��f���i
Mm Cv��W nRv	q�j����h	R�Ui9��BJ�2ʵ/;ldv���T�ӝ�,��Y��'�
�Z3e"���ӎu�D� �fJBBgh;����N;L�*3F���E��\"�4��)`x&4h��)k;�뉘<�� �Q��mz؇P��ۧW-�Wl�fz�7MvܙU�����l�6�  ��E����$���k�e悜�a�v��S���=Zٸ9�Jv�n�v]�3s�,�y;���cs�'��g��n\��;+V�sp�vy�C��fQ��V�p�6��ܦ�����̓`�5�g��Z��B�� En�YiF7g�e�qks7ls�V�<���麶|�]���v��Ԛv;]qr[ӗ&m �v���tl^�S�+m��5�K�$�ב�r��t`(��UZVl��i#��6�N�GO:�E���n�NC�u�m�ɈZ���ڳ��9�l�E�v����*�����:�:4�]��W�6{r6�I<Kۖd�:v��I7V�݁"�-���W\��k���on�Ϙ�8b��pҪ����٭���)�Fv+�1>���qY-����vӛm�nCvL�C.���z�udR�s�v7Bh��v�@�p+�H��-Ԇ汵�S�FKi��uX �n�z�:�]�� }��@N�Qz�|�G  -Q��b��:�b��j���q��Y�@Ek;��k�;\Çm ����G���N���K����g<>�-�v	.�^+oM)j@�畭�7�:��Kt�dȼcR4c����u]�۸v+vz�V���k�ōI�C�.��ON��#mv7/X'ӴR�ݺ�;Jv��C���c������7�+壌�J	.�5�k��fR#�/��>�{�/s���Dq��*�898�n��>�¢��<p�rl��(�?����?c�>�:��~a�=�������cȤI�C@�}V��S@�;V���h���m�2�Ʉ�H��l�T�rl1�@J�ᖨ�$�$�m�f�޷s@�e4W�hԻ��K�#�G��&��hv��=����6Ձ�ݵ`t(��]�����٪��Q�İS�;%��z�ɺ��e�tg�\u�s�޶���e���Q�쟭 �6�*@96vF3P�h)L�T��6����(��h�!����w��wZ5$���f�����U����7�5�h�T�rl���T�:w5��Q�Q93@����>���=�-�Os{�`n�����SuM�UM+����T�}"�� ?}��}���?~�y�b�o)ӎfKv��ɵ<L1g���f�غ��dФ�Wuּ�W{��;��ʐ�T��"�\s4e�G�0��ƒ�6���e4���sf��q�����QH��S#s#�,��V��͟B��� ��  H�4E"D�Q�SZ�u{�RNs��ԓ��	��q��onf��z����h�� �EHv�˔]�ٵ�Ee���.*@>����q�@?�߾�cX	54:��;cKr=�%��n�`��6Y}\��u�$�������d��@>����q�@sw X��J���2��:�,�6��D$ُ�����֬�֖b�m5*�a.���uJ���ٰ=��՜�$��W��Ձ��6��R�TMR)7U6ٗ M��EH)W�_w��VW}T'ezR�orOJ4ړ4����*@u�1��*@>r��e���e�q���y��.��m��gd۠��5@n�sm��b�����p.��zH����EH�*@J�Fմ�,q�m�m��<�W�w���z���n���.q�R"cxcR;=�ڰ3�ZYЛ�wZ�1����-����KT�*�u$Ұ與��Ł��`y�l��6ՀbŚ���Pm�y{� =$T��Z�"��������_�jDH�l�������l{�yZ�U�]nR6��\�q�#@\G2�T.ki�q9ӳ]���V�nQÚ�W3�{/-!/��X�C�7	�:��@ն�^yy��.�9�Bjg\�R&#R�z���}ƨ���9���*{fxB�b��m멕�k��~��}ۮ�͎��]̢�k�GD���V[��K/F-�O�΍�@�8�b���Tz����c�
c<��c<��!���!����.��!����kRXx�.tEuӺ��h΄;$�?�8���}�.�޲��Қ�ZO�b�90�)������J7;�Xݮ,l�<a�ڪ�$�$�m�f�޷s@��S@�}V�����֊_�&c��A$ә����ꯪ��E�@?�?Z�ȩ �EH	��D1�X��Ɣ������qmX��Vٕ��В̡lOU2S��L�(��܍pݱYjU�J⵹�mŁ�v盜���o�)�R"cx`�_��V{vՁ�ei�%�Ӽ�b��̵�*��T��&���ݵ~K�CdB1�$�C(d� 01BT��	zk��VXӚ�{���ΰXC�"15$���M�9h� H�J%��.�0�nb��a�(I�V�7t�V{vց��M�W�'�1dF90�)�͑R��`��Z�ܩf���ڄ��vȻ!�u���x����룫<�T�M��:�\k%���$� ��HG�@zc����`��.���q�H$�s4�JhW�h�R�{�4�P��qcR!7�����g5��u��B�J��D{ꪤ�݂���ʻ�e鵵�E�hn��*@z=����cI.ic�ѧ�����;�w4�JhW�h�R�������f-W `��H��	
M�Yn����n̘깢7�,X�̋ �"14���Қ�9hn��*@GR�Y�K�����sE���k�P��7_Z�77�XnV���ٽ7-�Rj����T��~T�|�G�@zc��|2�&bX�$��3@�t����M�9��K(Q�F���n��.jY5Cnf��>̭,��[��=��Ձ��M��]G�ш�䍸��':Ohq���]ע�vx:���Z:x:냪|�����M���l��̽��������Қ��q�\�ɍ�Hhn��@y���6ucV<�yH�!�{�)�}zS@��S@�vJh����$�M7�l�@w:� ;�T���ST$����?�8hz�h�d����wF�����ԐS�F Eb�[�|tӺ8���틯m�`��m��4���KZ]Ԋ�W�ne:�7<�61nNi9�:A�i���ؓ�G6Ꞥ8S%��Jɶ1�C�� f�[9w����]��s�a����ųn;��u�i�+le�` 2����v�7[�l��d�٫a�R�ګ@���83Ym r��#��}l}���!'l�E��Ջ�ژ�����۞�ԭ�>�,mf���׽�|~a^û�X��p�q���uju��{��ݵض�'_��𝱹��2�:75��6�����|��l�`���LȘ$�cx�w��hz�h^��=��M��.�Ƣ��I6���@z=���T�|����ˌ��b��>�)�{ݗq ��Ht� =�ӻ�A�{[W[F�l���T��M���o���G�wGLe��[<Q�6行�m/<�[��'Y���PZxS���g�5GM���]홴�|��l�a�UU}��-���\���Ĳ@h��pЛ����ʉx0@	J�����M����;�)�^˗E�a{w�� =� ۸� ���@Nr�n����m� ;�����{��,���/�Xf����6�ϾI.�*Z�K�v��K֫[��y�{������k����
t�*>�k.M��cu����sɓGh��7:�f��n;q(=n�}k �����~���|�^�QjI.�-��$�s�Z�J���1�q�!��R|�^�Qo�m�{]��ͷ�5ö�{/O��	L��H5�/�F�dœ	 �$�����%���տ=���p�'H� � 
��H��0��dP̉�u��!".1 �!�����0a�k�g�؍;��uϾ��K���Tg
@��Y�͉�0�$�� �
` g 3�R)>�q����\$�.#���"@	�U7��@#	x)[��Z	�[# ��Ҳ]#K.��S(���.A��`S6&pc!�!*u<N*�!�Q��L� ��+$������t^�(AO���b�=��{I/W(�$�݄G"Ȥ@�&����6�d�m���^�|�~{ZM��(P�1��}���W_��a?��M91jI/��O�I/+(�$�����K��Š���>��T/�.��T�n����/H�Z8Vں�vz�qƷ�x�U���O�8}�IyYG�$��/���%����I/�[~;>���g���K�4
jQ2'�$��/��߳j��qjI/u���$���z�K��U|,d&"$(�d���%���Ԓ_{��|�^VQ�I/���}�I^�ni���A$ۘ�$���������cV�w�N���z��J����RU�~��ߗp["�U)r�uG�6ߞ֓m��?(��o~Ř�}���Z�K�N7RK���fFŃ�#8����m�L(&삌�=m\�ܸ����GJm��[���@�I�u3AI�T���߿i�/�m���N�m��9B��������~�S�̾U,%Tˢ\����̝��!%3-�6��������m��=�}�DD(S2�Ǘ�#X$H�rbԒ^뿏�I/=�&�䒅3;����ͷ�=i�m�ͽU0�$uL�*h���(����m�߷N�}�m�N�v��>����m���.m�ҕQU(�Nh�m��a�/�m���]�6��m��ͷ絤�m�H��@�,�vߩp�ZKm�X�8�4�\!��ɹ��X6ٶ�4.ۑ�i	vyꃳ���vS�wB��Mr�.�sn��쪜qs�!e
���EVR�v7Z�k\��]�() �fx�gU#��9sn֝���ت����b�/q���ض�u��;��Z�v�kڱ�#2>͹��C���>R��pv|WI!��Vtmڭ�G��f�;�[i���D�\7?Ϻ��{��w~v���nژ��2^����9�,O&�dG��u��d)!�ܸ������}�}|��p�x�&w$������$����$������W���}�I~����7�6�&�N�m��>���������{����ͷ���ԒW/�Yq!��R|�^{ZM���cߗ�>S3�=i�m�f�|�^C�+�4�,Y0�R_���~�}�IZ�n-I%��i��%�������<�����r��/�m�ɭ���B�o�{ͷ�5ö�y�{����œQ�H��������yر!��\�e�ci��n1s[�8��ۇVu�ն�"��{/O�m�l֎�m��ˢKޖ�럅�$����b�bq)�G�I/Y��!b��Q-%S-�[ߗ�6�d֎�I}��}���m��_��Ճ��d�&(�$��}�|�]�QjI/��O�I/W(�$���^%�HȰi(��>�%��{�|;m�����o�[l��D������%�L1�Q<#M�-I%��i�ͷ�g_|ϛm�k��6�d֎�m�I~������G\�b�x�Gu8\���D�=ўL	t�Sc�z����;|n��Q��C�$����K����|�]�Q~���m�6�����-�T̺cMR&i��o=�~_}С%3/vk�m���|}�m�km��&e�j)�g�d��r��/�m�ٮ����z}��B�J ��.�
�����P�X�"0�+	c@ B	(DzD��|�U9�ޟ��J�?}�|�K��`�	)��������o�}�m�W[-�߽�~_|�������j�g*n��G4�ASG�6߶��m�����^�m��p������o�y����
*���9؊8�Z�qܺD��+�+�+�&�׵�\B�ٓ#��Մ��d�&$�<�J����>���&�v�o�m��	D{��ή�[m�Y�)�)��č��%U/�m���N�DB�"s�y���7�m���՚����;�{�wwwyS�����nBӀV������6߶��m�P�g3W|����g�=I%�x7�4ˌ��b�����}�}�5m����ݶ�n�t�&Q��n����o.))9��1��4�m��bߗ�6�d�m���ޟ|�~�ے�m��I{l��4�r�2i��b'�0Kr=�C��x�GG��]��3���:ݗR�Kc)�45NS
SK�m���Nۻ�tP����lV+���u=^��ݺ�Jְ��'�ӓ����i��%�.�RI{ݗ����wqjI+���jHN��*h������-�߽�~_|������e���u��ͷ���v�4:U*�sI�l~�-�}�m�N�v�o�m��;����V����m��o~��|�L۩�J�M��y�wEն_�����}�s�[������n��ݚݶ�qQ�"�E	
;�s�l�ۉ��\�9��nx�X{,�2�k;/��SӜ�)�L�y����ݼ7�cp��i��Q=S�%���AۭdU�����Wv��Gh���������K��zօ۰u���Y�xi�+sRtuL��X�]gŤ�gط=n:N���Y��Z��6M�Ԫ�%�X����kGdU ��nk�8c���;�T�l�zӉ6�;8���qD63��q&TD�� �:���bL��379]�6뮅��y[�`{���W�\pp��r�7�n��{�P�����p
� ����|�~��e����oˢ"=�m��[-��.иr��%S&eHꏾm�l�|q�~�Ol���}��m������"�f^̴4s�M�)4�"f���y����ͷ���v�%�f}�|}�m��Zv۷|&oqq;rRS7�7�o��������v�o7��>���V�-�В�3���g�$����dLD�GԒ_{oO�m����'�m��;��ͷ�ٛ`����y�y'�ݼ�'r����ڇPM���M��uv��T�;D�=���͸t�8��#���V�ۋRI{��g�$����I%����K��*���Ĝ5$�9{�]�(�>�� ��!�%LA�P�J�"��)��6gW��j��oJn-��H�L�UR�<�l�����e���{�~��/�U�cXړbMG&Ò������޵`}�[já(~���[u�\�4əR:����mX�QR��b���T�&�W��hbBܪ-pLU��ּ��v��u�1��&vݱf<1��!"y�d����컈_I�s� ;�T�󬻗u+t*�2����@z㘀�=���QR�6�}�f�[�A{��s��I9�;�S@��D^��P�(��R�V�ޛ1j��ʩT��v���� ��Hs���b��M��u�d���LI��>�e�@z㘀�=���ʕzx<��	L�`D�[��\������'E�LlP�M��:�]�z� C˫��~�b���*@z�& 'K����1�1ƒiH��қ�/_ۚ���|�W�[�)�4ˌq�b��3ٶ���l����?��lޯŁ��pf�NU1��4�9&����>ޝI7�3٩66���4�/u�|jI�o��ڧ#�Ҫ�>{�6��(����Z���j��q�P;�U;���3���E��Mafx���Ѧ�z,ݙ1�fj&(�f�-�� ���=ָ�3ٶ��b���>ޛur�t5R�KuL�*h�3ٶ��D&�٫�����>�V��(���ѳɃ�*jSUR�74�٫����l��"!&��\X�֬x�F�Z)���53%U��IB��%9_����_�=�jÒ��i�h��_�bM,jLq��R=�ui`~���.�����?U���ٰ/���m
	��b�0�B��F!B`E� ��(�"�H22u���D ����Q|h��>��nRRaa�W��	�8�ƾC�$O��ݡ#�!�92��ϒ�򫌔�e�dA$A�TBL�*I4n5�]h������.���V���GD��O�0�&����7~��M*�a�e�T-% �@ٷd!��)��0���[Ӻ������wg~������+�Gd�;`^GV{x��D�mJ�r�)��!A��K��*�t!Vtv�5�����.z�vҴ�d)]�j�U���@H[5T�U+d�WV�J\H;2�`�F����M��3*dN�7�7,#a��͹�Sk�(���P����]+,���7[s��7M{qr���Z�;N���ʳ�ΫHs�섪��*�_�g��q��� X<�m�*]�nz��)z�1;��=�.��M�s�\q�v58բ�u���^�(iܘ�d:x���rF�@.��l烂 ��׍���I-v�̑m�<�]dc����m�{m��'�}�����$�&�Ċ�lѝ�7q�δZ��{m���]�������`Г6�`�%��V�u�]�l�S���.�l���+�� �-�U!J���7��}'lDZ���$�6k��Y���d$�G$�5^�=V�D�p�K�r-�OK��@Ԇ��='@mT�uesX��T��v��c/�k��]�қp�����M�_'��Q�]�-R��G���A��.ʨp�`�j��E� �	��y{K��$��.u�n�\�d��=l���V��1�ƻr�/�,n�nUzsBɞ��7^��Yt�c�	��]�	��rܛ;/�� ���.gR�����n6y.'78�`:��n��[<��G*�<���N����,lNR��&'����Cq�ۯ'hڳI��qJ���N!���,�ә�N��^�;8t=\ݫ�ٻa� �a���9�W8;� s���UU	v�٬�曝���z�/6��m��{g�\�섲�U�%ۣet����S�'6�1��!n�nm�%�Uvy���sہ뎅����gl��dUz��J��a��[9�J�k��ƭ���@���s.���s���SM�;1�i��i�@S����t��έ�N��-Pq�#�:h�2�vy6Tk���;n�tCȬ���%�.�\��]N��K�
�q��$p�� {���������}��w���2A�� �6�So�T��G�/�@;��{���~����Yc�9��$�!ۋCU]@R[�-�y}�Igk`��m��5Ӎ3�9R68�����k�}��Mt=��h�-�ɵd$�(S�g�D��el��ۨe��cv�r��lS��lĠ*��h�&�����\����s�Mn�\C�i�N8莀�.N�<يWp��H-[VT��oE�f�����6��e��$VH�9�Ofn�gBgn��-�k��s������������c��ԡ;���R/:M�8�q�]�=g&���-ũ�.��������	�4��8��1H|���� �r�@��l�{6��5�5�r��5H��`�{W�Q�!L��w�3z�{6��$٩�㥺�M�a.J������>�V�~��&{{�� ����f������)�u56	?g_��� ��mXt$���t����ST�)n��M��j��
#'t��<��YM�������a�8E2���֌�ᶳ�=v��Ƹ����u:sۍ�������j���Ĝπ�i��/Z��s��Q?(��;�~ѩ��,N���)]��KM�Ne�\/�L��L����_�
����Ȋ�� JEzAC�(���I�&�zi7ı,O{�٤�Kı/y���7�Pq,O��bcv�91�[qs��I��%�bs����Kı9��f�q,,K���gI��%!2�;��|Bd&Bd.�m����sf1��3I��%����w�4��bX�%���Γq,K������K��,AD�}��I��%�bw��?ΪT�4�"f�����L��O����7ı,��{Mı,K�w^�Mı,K��i7ı,������Ve،e�#S�r��ލ���h9c���k�1��]�����o���{����42Z��$�*��&Bd&B��t�/��,K�w^�Mı,K��h?(�U>���%�y�O��n%�HL��ŧ� U*&d�1���/�L�bX�s���n ��%�bw���&�X�%��s����Kı>ǻ�i7Rı,Ot���e3�&-�l�3��&�X�%��w�4��bX�'1ΞƓq,jCFU�Ȃ"&"s߱��Kı9�k�I��Bd&B���Z�d�9SU*�sW� ��$P�Nw^?]&�X�%��~��i7ı,O��zi7İ"PK�ﲚ�H�v��\6fɊ[��pf�I�7�{��D���f��,K��;��7ı,O���w�!2!rծ���)�
��>�y��t�,�v6�M�`�۞�M��u�s�M��������'�tdt�rd�������,O��l�n%�bX��}�&�X�%��g���q,K������JBd&B����/�fT�*eI3J�|Bq,K�﷤�ı9����n%�bX�c��4��bX�'���i6%
!2!d�N��U4��Lզ�X�%��g���q,K������K[�����&�X�%��w��n%�bX�1��Rgm�1I�\�f�7ĳ��D�{��4��bX�';���&�X�%��w��n%�`~(.�"w���t��bX���ŧ��J��)�njn�&Bd+�{�4��bX���|i>�bX�'}�_�I��%�b}�w��n)��	��jێ�Um4M���m�
V-�b�<W[��m�n���K��I��~�{���M�)�R��U2����|Bd&Bd-���&�X�%��{���Kı>ǻ�i]ı,K�w^�Mı,JBܮr���.]KT��W�!2��{��� �,K�{�Ɠq,K���צ�q,K��{�M�I��	��f���SU(aCt�f];�q,K������Kı>�u��KRı;��f�q,K�����_�	���_O�R�rT����i7ıA�>�u��Kı;��f�q,K������n%�b"�^��	��	���n�t���Ng1.s4��bX�'{�l�n%�bX~�<��]'�,K��?~��&�X�%��;�M&�X�%����=��Z��k�=v���b^%�Zm]4�;i$��%�e4``�y���a 9�E��ӑ���-�f�o����S��9�ܻ13H�������ݓ��-����8�5��.]=t������B{N��qכ�ݹpو��v����� ![+���K#m˹惛�nݞw7�"GLv�s�R\rն��d��Ju/4Ys2�r7?�����������\Վ�m�Lp�t�+L<V3��4^�=Nm�%�=<=[�7eם�w�ŭ���k��2b�&�q,K��=���7ı,O��{Mı,K�w^�Q�Kı;��f�q,K��_zٛ1�\�+�f��7ı,O��{Mı,K�w^�Mı,K��i7ı,O��_]&���bX��f�bHf� ���9����	��	���|\/�V%�bw���&�X(X�'��q,K������Kı=�Ǥ)��T2Bb\�p�!2Bd-��X�%��{���Kı>�=�i7ıR���צ�q,K��3�3(�II��5I��p�!2!2�nz�7ı,?� 3�߱��%�bX����i7ı,Ns�٤�KǍ�������E3�����rLdDy$O�\tnN����g��.��t;E����}O�=d7Cr�̔��L��L����M���ı,O��zi7ı,Ns�٠ı,K��S�I��%�b{����T�rT���SSp�!2!2�o��p«�!0
2&�b%��w�4��bX�'}���Mı,K�s�Ɠq?�@�b&"X��z[���9���8��s���Kı;�~٤�Kı>�zz�7�lK�s�Ɠq,JBd/n��!2!d�o9���2`�I�d�n%�`6'��O]&�X�%��9�cI��%�b}���I��%�'9�l�n%�bX�1��Jf�g.%f2f�7ı,O��{Mı,K��^�Mı,K��i7ı,O����Mı,K�:��%����6:�I ���oF8�kl��t��.���q?w��|�n�]�3��ı,K��^�Mı,K��i7ı,O����q,K����p�!2!2w'|�	�T�$&%�Mı,K��i7�Dq,N{>?]&�X�%��w��i7ı,�����|$�!2!fW9jy�]'3Y�Kq�I��%�b}����n%�bX�c��4��c�r�,P��M"��,O��zi7ı,Ow�ڸ_�	��VoO�J�9�NIr����&�X�*'�罍&�X�%��{�M&�X�%��w�4��bXb}����n%�bX����m-�.p\�[��gMı,K��^�Mı,Ky��f�q,K������n%�HL����_�	��wN_R�T:��A�c1�w[���;n���>}`y [�p�3z�ci(������~oq��K��i7ı,O��O]&�X�%��9�c@��bX�'��4��b�	��MC[��9���"f����ı,O��O]&�%�bX�c��4��bX�'��4��bX�'9�l�n'�""b%����~ɋ�pB�.s3t��bX�'1�߱��Kı>�u��KlK��i7ı,O�m�_�	��7K] *s@���%��4��bX�؟w���n%�bX��}�I��%�b}��z�7İ2�
��������Kı;�>�Ԧ����	�sE����L��\�}�I��%�b}��z�7ı,O���Mı,K��^�Mı,K�(���	R��.X*�J�Le&�N^�H��"���Eyı�˱u�lQ��-����~��2\c9�Kq�I�Kı9�j~�Mı,K�s�Ɠq,K���צ�Sq,K��;�Mı,K�����9�NIr�&Jw�!2!zs�t���%�b}���I��%�bs���&�X�%��{���O��D�!I	��o��|��]Ju#r�jn�X�%��{_��q,K��;�MİlK��S�I��%�b}�{ظ_�	���F틩�:���T�U4��bX�'9�l�n%�bX�w���Mı,K�s�Ɠq,K����p�!2!2I�kz��'4��1��Mı,K�秮�q,K���{Mı,K��^�Mı,K��i7ı,M�����0���Q=��+:*U(^,;�Z4 �q[ҏ�)iY�FD��m8�9c���u��8�W��ɭ2�[Gd6HJ����짮iG�S�v*z�(���U�ڹ]�cs(
f��Ƕ^��>�mܸg����/�{�N S��::���f��������M�4c;*�*���V�z��G�gӲgF�Krp��;��3hò����w�]���hD��F�g�0��g�]P�G;�Rq�2%C�����z�����1���Fm�i��ɛ��Kı;�~��&�X�%��{�M&�X�%��w�4���%�b}��z�7ı,���ΐ9�URR3Up�!2!8�w���n %�bw���&�X�%��g���q,Kļ�}�&�	�
HL�߿'���4USh�LL��ı=�߶i7ı,N�==t��`��b^{�Γq,K���צ�qL��L���K�luT��ST��W��K��O]&�X�%�y��:Mı,K�w^�Mı,��Ow��&�X�%�����.cq1����\�Mı,K���t��bX�����I��%�bw���&�X�)��+W;��	��	���ܮ�C�L��XSd���竃���t��b��烆�i��m����K[�����ߛ�ou�b}���I��%�bw���&�X�%��g���ı,K���t���L��[�۹���SD�L�n��_X�%��{�4��>�]��L����Kb)!PkJ�! ��-����KFF0X�$�q@ؠpdK������n%�bX����t��bX�'��4�� ،��Z����9�Nh%�"f�����,K�秮�q,Kļ�}�&�X�@�"b'=�~�Mı,K���f�q,K��_��31��!1�7I��%�b^{�Γq,K���צ�q,K��=�Mı,d-ͳ�����L��Y�l�S�)���,�3�&�X�%����M&�X�%���w�4��bX�'y�O]&�X�%�~｝&�X�%��;�7��� +������3F���x�s;�X�㗞)`:��ݮ2���'���wۧk�$t��&�q,K��{�Mı,K��q,KĿw�΄�Kı>�o���	��	��g򦊪nf��C�M&�X�%��wS�I��%�b_��gI��%�b}���I��%�bs���&�~D�"b%�����nc�c3��Mı,K�gI��%�b}���I��0 )�·\`A�@��7��- geH���*h ��!���������?�|?}�87��8�xbKG���v�0���L�Vh��ц1��	�¤$ B�Ӂ�d�	��H���
"12�"k
G�肮��;� �"�	��@"@0D��� ��P�Ai�A�@x�� v�Ah��;@J�V�J���`(�M���G̉bc���&�X�%��{W�I����L�����u,�������|AbX�'��4��bX�'y�l�n%�bX��u�]&�X�%�y��:M�L��L�����|QD�AS*[�.�,K��=�Mı,K����Kı/=�gI��%�b}���I�	��	��x]�D�R�f�ә&{��k�j�k=.�<ɺ8*g�z�r8�x��ra���T�A-��+��	��	��v��I��%�b^{�Γq,K���צ���&"X�'����&�X�%����S��))����Mı,K���t��bX�'��4��bX�'{�l�n%�bX��u}t��bX����ΐ(sRڦRUUp�!2!X�{���n%�bX�ｳI��?��&"{����&�X�%�{�߳��FBd&B�\�P7?T��134\/�V%�X�罳I��%�bw���4��bX�%���7İ8�PY�|\/�L��L���-���7RVpd�4��bX�'{��cI��%�`������Kı>�u��Kı9�{f�q,K���O{x?ɚ�#8�q�`�&������r(��z�ͬrce��m�쑺����qo%�p$���d�,K�߿gI��%�b}�k�I��%�bs����X�%���W�I�!2!vq�&UMM9t6����[�bX�'���4��bX�';�l�n%�bX��u=t��bX�%�}��_�	��{F���&�
�R:��q,K��}�Mı,K��q,ı/;�gI��%�b}�k�����L��Y'!����h��ri7ĳ�\D�u���n%�bX����:Mı,K�{^�Mı,K���i7ı,N���c�ť�XLd��n%�bX��ﳤ�Kİ�����I�Kı9���Mı,K��O]&�X�%���v~�?g9&-�si�TK'�Dl�^�U����W%&���r8���P*��1���4�q�l���c:CFZ������^_���W�F_n�F�ɤw<�g�Dl�5��Y�X��.m�[J�oDs����rfle;Z�����s��O5����t��*�r܆�ƺ��)��F)�/[���ƍ�z��Y-�m�ѳ��y�mxc4�����{�����������ĶNZ�:�x�
�gM��8��;K�;.
�yn'��ٓ�<�lG��ˮ��Aպ;]�����%�bX����i7ı,N{�٤�Kı9����n%�bX��������L��[˗J��$�R&�q,K���M�Kı9����n%�bX������Kı>���@,K��;�[�%1�ۜL�Iq�I��%�bs����Kı/{�gI��?°1����I��%�bw���4��bX�'9��8	�˙q�b���n%�bX������Kı>���Kı9�{f�q,K ,Ns==t��bX�'���Ɋgĩc��T�U����L��^ξ.�&%�b����I��%�bs����Kı/{�gI��%�bw)o|L��PֆI�D݄�F�����>�{E�ꎩyo'4��b��E���<�o�ߛŉbX����I��%�bw����n%�bX�����q,K���צ��	��	��u���9	h�34�7ı,N󺞺M�B�"�0�����r�4C`*�1ı/�~��&�X�%���צ�q,K���Mı,K�9|b�_g6�e���:Mı,K���t��bX�'��4��` �%����4��bX�';���7ı,Nw�G��L����,�s�&�X�@" ؟{��j	 �｣BH$��9{��@C�/;�gI��%�bwǏm�����&c�Mı,K���i7ı,Nw���n%�bX������Kı>�u��Kı=�x�l=rm�A�[8�gnn�s��ݹ���[Җ�}}�ɍ�7��?������q�s=r7|�D�,K����&�X�%�y��:Mı,K�{^��Kı>罵p�!2!2f��Sb�u3CS#%�t��bX�%�;��7ı,O��zi7ı,O��l�n%�bX��o���P�,K����nq��K�i3��:Mı,K���i7ı,O��l�n%����Q 4��dK<ϱ�i7ı,K����7ı,N�A�.N���3J�|Bd&Bd,ｳI��%�b}��Ɠq,Kļ｝&�X� 'y�l�n%�bRI�f�yL�BZ)9�W�!2��wW�I��%�`�^s�Γq,K��=�Mı,K�{�4��b�	��w��$M�9c&jf�e&�5�g���ͲE�rJn'��]�p��s�/5)s�f���7ı,K�w��n%�bX�罳I��%�b}�{f�����LD�,O�����Kı;�M/� �R*��9��_�	����f�qAKı>罳I��%�b{����n%�bX������Kı=�ǌ�qpc2d��2i7ı,Nw�٤�Kı=����n%�*X�%�}��7ı,Os�٤�K��'v[�CR�$Ԫ��+��	�X�%��秮�q,Kļ���&�X�%��{�M&�X�B��q���i7ı,N�v{f-�1�fR����n%�bX������Kİ>�u��Kı;�{f�q,K������Kı:t���&3�%!������Z��b�ko&NK��{dٹ�l��cm����կ��E8�X;K_{�ı,O��zi7ı,Nw�٤�Kı>�zz�?>���%�{�ߪ�|Bd&Bd/߸�$��Ԣg��n%�bX�ｳI�~@�&"b%��g���Kı/}��t��bX�'��4���"�"b%��O�g'?���KE'3J�|Bd&Bd,���Mı,K��t��bX�'��i7ı,Nw�٤�Kı9��eOR���K�Sp�!2D2����n%�bX�w�٤�Kı9�{f�q,K�19��~Ɠq)	����?1:�U�1�U���bX�'��i7ı,? G����I�Kı9��~Ɠq,Kļ�}�&�X�%����T�����&uYŦ��Wb�o j�V�#�ʗ
vc�F���v��]t�@+kC�XN���gsͳ<;l�H�;��h�^����G�4���ݎDA���1�A<n�I�$V�˻k���g��Z-�Wh%\s�cs���z�$��[ɒ���ֹK�vx�AG]d9�4�U�ѻi"N0��Nr��E����vǃQ�3��9�\g=��k�5�W��ۻ��{���{��q������Gd�6���@#HWD:3�Z�@�����]I�=	wn��1������]�&����Ld�q���n%�bX��l�n%�bX����t��bX�%�=��7ı,N{���n%�bX�c�Ÿ��K�T�R��i\/�L��L��N�_E[ı/9�gI��%�bs�צ�q,K��=�M�[ı9��m%"��A����&Bd&By�դ�Kı9�k�I��%�bs���&�X�%�y��gI��%�bs���S2T�t6�UUp�!2$�;���n%�bX��}�I��%�bs��t��bX�@1�{�t��d&Bd,���I�����3T\/�LK����Mı,K������Kı/��gI��%�bs�צ�q)	��ܷ��TD��$�J�����;#�y+%ۭ�R���V�\�o���si�NA��\Ҹ_�	��'_uZn%�bX��ﳤ�Kı9�k�A�Q"�D�K���߶i7ı,N���Z\~��8�I�ۜ�I��%�b_{�Γpڮނ��
�dK�ﵯM&�X�%��{�4��bX�'1��gI�)bX�'�3��	3s�g0�%��s��Kı9�k�I��%�b{���&�X� �"b'q���t��bX�%��߳��Kı>���,�.pb��I�8�f�q,K?*0C=���&�X�%��z���&�X�%�{��:Mı,Ȑ\D����4��oq��������h�F�Lw����ı,Nc��Γq,K��{��gI�Kı;���Mı,K��W�!2!fu�2���B\�j��qN�e���	Ol�(��r2�\&�N��v��u֦t@�1��Lb[ns�&�X�%�{�{:Mı,K���i7ı,N����n%�bX��o��&�X�%���M����hmUUp�!2!19�{f�qKı9���I��%�bs��t��bX�%���t��ؖ)����ˎ�U1̢ff�����L���;�M&�X�%�y��gI��8� ��i���,B �!Ӏ��Ce��K��~Γq,K����f�q,K�^���s�d���uE����LBļ�ﳤ�Kı/��gI��%�b}�k�I��%�b}�k�I��%�bp�/�1����)Ld�q��Kı/{�gI��%�b���4��bX�'���4��bX�'qӾƓq�7�����~�y�p�dgM�r�m�[����[�c�c����t�en�'Z�p�������ET"��f��|Bd&Bd/w_M&�X�%����M&�X�%��tﱠ���&"X�%�}�:Mı,K����]���2L��34��bX�'��4����&"b%��x��i7ı,K���t��bX�'���4���Os���������aїSp�����X�%��x��i7ı,K�;��7�ı>���I��%�b}���J���L��Y�w�LSB��T�556��bX"ؗ�w��n%�bX�{�٤�Kı>�u��K���B#�� ሒ&"��x9܉��ױ��Kı=�Ol���6c��9�s��Kı>���I��%�a�"�����%�bX��?~Γq,KĿs�Γq,K�������s�ZQ�j�՜$rg,�;���Ƿ[�
W;tg�t�]��m��r���a{.1�I��%�b}���I��%�b^v{��n%�bX��w��n%�bRw_�!2!zN�O&�ԧd�.s4��bX�%�g��&୉bX��w��n%�bX�����Kı>�u��O����%읟�EUI�:�H�5W�!2!<��W�X�%����M&�X�bX�s���n%�bX����t��bX�'y3ӘS5*�)S�j��|Bd&Bd/w_��q,K���צ�q,Kļ�ﳤ�K�lK�{��n%�bX����Xϕ��"��h�_�	������n%�bX��o}�&�X�%�~�}�&�X�%����M&�X�%���>+0T08>"a�BA�����RF[)$r�ji�c#�ZӔ�	BDX�AIHŉ:�r��c�A�$FB0�F$HC$V�0 BA!$����Pa�A�$T�5�2� 40��h�I��n��V��{�W����� m�����h�Wu����@�\��V�<N@�6u�I�i�$��3�<H3��p9B���i6m�`� u��T���-�6��( �R��kJ�		d���"�V��3ہ��=[k���{qnKX�q���Ҽ�1����(
�*v��%'J���L)�]� m�"ʲT�*ͪ�@�!���M������7�J�r�����ݫ�V�N#[\���������!�;-��`�ֲ �_&�eN ��Pw��P�up�Q�N�u��me�;_�$º۵��x9묽�k���y��ױ'mtCp���F�N��h�=y�j�*L���� ���:�T� 6I���Z�ga�������
gh6�^`4�]
드fZ��v��*�n�#���3�pԄ�P��jU�����ٕeZU�@I�gh�w-�	lse2�RJ��Ci9������wF���K	�X��D�Y������L�Rt���S���nܳS���-����r�
��k�9m /F���� 6YoI,vD�${:,F��\T�!Ȧ\��t��Z��\h]���sh6+coc�=�\�{q�k�&��7o�˺�Ý^��9s]��Rn��n�vw�l��v���u�էl��At,v)�V[*�DQUh��5���	3����[�|tG/kgԞ��n�W� nQ5n�����d�S�-��dҘٔ �eZ����llsW9�&�'*8g�]���s��V�I��R�6˻wi�����aV�+���d��h&�FL=�1\��-��.�\V.F�� �0EHp���-��͖^�[*�������ؖ�'4ڻc/Gf�e˲FGr��3 tP����gq�s����+�`�0m�R�ێy��F%E-���M����,��<�Sd�u�:͢�E�m�6���Uė3�[�IRZ��؝l���$:�.���� nC����9�ʆ" �@6)��U	�T�T �AG��� :��G(1��pA��Uz�C߻~�����4�6{\n�3H
=Ld����6�j�G��B+b���-�s�l�P��'Wl���+�n[�{8��[v5<�C�Iy'�S%WULD�Տ;b��L{O6�ƮN��6묦G>�h1�T3̉�f�{	�[�ٶ��Zڎx�wh��;��3	�N�!����G��6X�7L�����y� �N՗G��mg\Lhڒ��j�����������{������&ݦ��:H]��ؑ��a�[�s�k�BXc&��m`�=��J��v:�Y���q��'�,K����t��bX�%�{��7ı,O��zi7ı,O��zi7ı,Nw�۵�4��f�-�q��Kı/{�gI��%�bs�צ�q,K���צ�q,K��;}��7��"X���~ݖLʒ��T�9����	��	�����\/�,K���צ�q,K��;}��7ı,K����n%�bX�{�]bbD�U1̢fj���	��	���|\/�,K��;}��7ı,K����n%�bX�����Kı>����`ԩaHuE����L��Y:���n%�bX~�����>�bX�'~���Kı>����Kı>�g��c���t��<�z��dN3���G>F�
^����Q�gK�s�h���PYΓq,KĽ�}�&�X�%��{^�Mı,K�w^���Ϣb%�d'�~�W�!2!v�߂�Jt�U&�L�9�n%�bX�����09C��S.�X�'=�ni7ı,K�g��&�X�%�~�}�&�X�%�˗.c>Je�"�fh�_�	����^�Mı,K��Γq,Ŀw�Γq,K�罯M&�X�%����6*N��3N��uT\/�L��LK��{:Mı,K���:Mı,K���4��bX�'��4��bX����4�)�i�`�UW�!2�y�{:Mı,K���4��bX�';�zi7ı,K���:Mı,x���������F��&4�8�j7b�^��;ƹ��<�oc���l�u�5�ӧ/V�s��Kı>����KĤ,޾.�&Bd&By��|��V����w�D6�6�4�SٟىR�����4���*<	*�$e��{� �9�I5
�(_|}UbI2$!,�iD_��K�mi`����&8�����~��h�,ݭ,?BM��`n��S�y"jI4���-���:� �l�>^T��Sx0i��/���Wsɗ���u�ϴ��/M��;I�f�s��^�Ic��F�u���-�m�@���Vؑ��&�1�NC@=��_$�woU���Ł����{3r�0�bX�$I4޳@����)��٠^�Ԗ��o"0UXtD(y�|X�\X�ݫ�)����0(��)�ȑBU$D�|��P�ߵ��I�zK���"hmHh���{�f�[�h�S@������5��G&<o�n����je�rk��.��xz��(�I��&�<h&
C@=ų@-�4[)�[Қ��qԓX1H����ڿ͙�\X�\Xx�j��1��dȰyJI�z�M�JY����VݽV�Y�v�
RL�**f������=����3ٵa�?n��@��Ac"I��9�Hhy�@����|�k�����q^�����3S�Uɲ��G4@�کUH6�v�iv���y�:�e%۵mg���c���{�����v-[�S"c�G���N�t�Ռ���;�]�>�+�S��T[����x�s�t�J�e�y&��+	[�꓎wk�J��y�k=m��wMp��2)v@�v�"�S�l�l�Gq�oarXc�<\��X�v�5�i�m����d��go�ww]���w���{�� ����9�t[��Cq�÷=��nma�&����lnɮ�1��-�&V]O���`}�ZXnV��>a�}6����%$j1���I&��t����=�\X���`�ھ�2~��t�KTU'�CjC@����4��W������>̭,������,r�9��ǲ�'��Po`�����ed6��,��@-�hwJh�M�>U�VٌoFO��F�!-�{1���n-mǷN|�5�$n*�XS
ht�ֹl�YY�`�8���Қ�S@�ϕz�٠vvu5��&1�����@�e�� Ȩ�0*��*c�c̀{wj��2����铿O~T2S�Lj)�"Hh_��z�٠}�)�u������b���,hm����?���~�������>��^��K�$�MF7��@��S@�e4��W�m�Y�\$�&�D�!���Uݳ֣���6�L=:��U.�a�yxN�I�!��Ԇ�m��>��^�[l�>��*<	sh��Ǎa1�������	(l;����mq`n�i|�6��RL�nI���MIS`�{:�o�g�S�I �d�D"���A�hac"1a�HY# �#H� Xh�2�RT0ȆAȨ�g������@�^�7Z�����MI%�������޵`|�f͇�M�wU��r�5��&6�"1�������nj��:%o���J����
1���O[���(:�;��Q���Of���}���ݜ��s����1���]���
�����T�9��f�[d�SS`���6{6��;;�X�Z�pC���RM��ȩ9�- G&�t^�.���Cm�����B� ��i'�X�$R0��D�.��@��$sĖ<k	���礴�����T����sk�[u÷I���&t�q�p�n��y�zz����{P�ͱn^p�Dܰ/0��Z95� 9ȩ;%K@uvF����0x��ɠ^�M�n恾�5��v����勑�5*A̹�#�u��s@��������,d��5SHh�)M!�+��]ð��7�ZXt'������ʢ����w7K@���@>�R};��=�� H�(����uR�QM)Ӽr��u�I^V�V��l7g{]J]u�����5�Z؛K�������E�b�7t��u��ݪ�^��y��J�2�K����v�E�w�@�[��F�Ph��fPU\G����ŵ�GG��ɹ+�k��U�m�m��v�l�=vy�ʭ/l�G�qW!�yC\����u�u��Kuh7�ŀ�;@Gu�&9�n+Zs�\ɝ)�hL��qw!s�&s���N�s�'���D;N����Y6nn#3�e���$9�ȜĘ�
I>��4��};��/���`orq-ъH�m��n�|��@=z��Jo�H�V��X�bK5�m9���h�5� $qR �:�!���Hr@-�4�)�[�s@�}E�\��(��"d{��� ܊����95�7��� ^l�틶�;H9��n9�rm�t�3�.oQ�����|'}�
4e��ߕ 'c����o`�ܝԆ���%MLsJ��Nh�b"!@��U�UZ�@ȒP�"C{�Vv�ٻj�=��)�*�A*�U5C��ڰ72������֬<Ӧ��i��UN��n��n�<���"��sP~����~�~���j�6�ڐ�/���?�$�M���z��kK�.ż}J��Hݷ-W]_0�cP����n����q�N�+���}���y6�,��w��ڰ>ݭ?%���V3)�1J������73j�D6{���;;�Xbͫ�e�4tUHԲ��5V۵���ݵf�lB�KH��!���J�P"M�0�7��m��5LDp"C&)vb�����wF2��A���E�0�2��9FZ�A��T$T&Q`�:z�b&A�%R.��R�e�0���
�#c(�&q���"c�E�P�$��"�1H��,a+
FH0 )@�1`�8���)���!�$ 	�e�?1, ��c�Q��1$!h`4)�+UҢA4!@��i�%>��G(�����4S �0�W	�Pt�QT�@� 	�D ��6����8(��Px��Q���D/D$��H\���=�V�X�l�7.e�6Թ���$��O~��Vܻ�X^�@��M����X8Lq'T�1fՁ�BP�w��=�\X���������?q`�n����)b۲	��|r������<d��6��
���[��V�Y���~��� =$T�gY�{Ի�d�"���M�e/�%	�{zՀn���ڰ=��[�!�H�o܆�o]� �f�[�h[)�v*��\�I0h#��9�j �&�=&��������D�@�y��ԓ�>����1dm ���l�>�S@�s@=�Y�y�u�!��ț���Œ����m�z5��Pi���gF��)u�:����t$bƈ�rM�e4��� �f�{����˭��M6�IcNt��1�@�5�6��_]�u���X7q%&hR����P�`�m�H��2��J>2������&�=&� ��H?UU]�_�@����X�y@���4���8� s���.�U��:�����[�
.�� -�0p���������Q��v�0���̭����[VKe;{y�q���@��I.ª=��Y ��yV�6��{�l.^� {&M��ٍV���+;6B7c��]%�W9xt�z�s�ݎt�<��J�;m�	��]�X��l�M�5������#ţ/�{�Ԩ�[t����Q���{e\���1�g��Ļa���!y�hzȤ������n�������G��d�$Ҭ�71�4j,�ݝ]�S�tg�5�&�����b�[�J+»�t��1�@�o������Y-��pP��)�	�V�3j�>�f����w]���U�:�ŉJ6��@rj�l�T���`j~�.	�S��e9�Xr~�,wu�,ٰ�ڰ5jʹ9��2����s@;����@��M ����J����,N?�6�g�5×jе�v�Q6%i�Mp��\�����X6D�I��q�h{��>�S��=�֬3y"��S��)`55V�s��C�bX��J"|���	�p�ZI�{ZX{6Հf-٠{֭����8%��M��h�*@Ԛ�<�����Q�����e�e����+^���6�[)�^�Y[S",�Nf��Ԙ�=$�I�@w8���^JL�\E��������V��Md��C٩���8�:��l��3ێn��O�t���6� ��W��'L �&'&��e4z�h�-z�l�.\�pLY��	��� �MG�_|U|I��a���	�@��Nf�˲נI��`��EH�σwo6��K�T���X�3�����Vs-z�*�)�ěRA���,Y#�#^p�=���'s,�)v�r^8��n6m���8�	`��@�����hv[4�f����B�mbm�hک 7Rj }&�:M��.��&D4<Y�� ��f�w����@wH��u��	�WWWza����ݫ۵���nڰ؍�J$@>��c!a��Y!�@���0�`����BBT�����%Z�¦�=��4ؽ�౟�dQ�D�rh�R��ݵ`�v�76���q����9;#�6��J���N��،�b�1���ޠ����c�Y�N"G.OĆ��� �[�`�����,�y$��8��hv[4�l�:M������n�VYY�e�u��rj�f��� 7Rj��&��#����>�]� �^�@���@��R���b�ۚ #qR �j_I��`���L�@3"H�Z4H;;�;9{4�t��7n��jpJiF���[s&r4ղ��S[VQ�u�@���1�a-�q����ź����8�.�H5��Y@2��A�s�v�a��c�jG���m�۷N�M �l�75vj����
��:𱽕�:���v�&Ez�z۬���*n�H܍�A[����&wO6eDT�zt��7�;=��g��Ǧ���9m� j�g\ͪ��s��5�Jv���$���Fx��͞�,u�[�.����rܭ��]u�4��F$0X�ɑ@R�f���1 �l�`��:�eٓ(���ߌ���@z�L@>���U�4��<+ɂQF%7#�;�Q�{������T��+/AU������|X.ޫ��@�YM ���$�0l��9������@{���`O~�G��-6OfW����E�v@bݲ�95�����v�rk�-�r��ɹ6:������� ;�� :nj�t����1I������g�w=� t�����s��Q�י��we�� ;�� :nj��b�Jh�PX����
C@;;�@z�L@zM���λf]��1bY?�2I4������;�)��6�J!FN�+�(ULqN���]����U�k\鄲CcW��\X")��mg�Ƥbq�E���߿OƁ�t��vwY�|�W�}�-�1��QH%��� =� t���9�I�@���Lsc��r��f���5>�0`�{	@
��� �G5
�%"��S �%�;�M���=���/�hI&��������uq`fei`�6�ͺ	I�$D�D�z��h�����-�4���,�U���0�ki9��۵k��率Y�{0Zr\0�U�w�i��9�1�&$!�h����4������=�Q`��-��,f��(P���w���uq`}�Z_%
5<6Q#��4ڨ&����O؀���� M�@<][iU �Q�5�H����>�jI8s�Τҭ2�JR�V�j*�*X �R!���5$�{-�1�E �F�4w]� ��@�[^��YM�'�MF��&�v4�F�km�����s��1�oN�������wƱ����1'?��FLD�	173��M�$��� qR��[ZV�՗[ee�������� 8� :n���K	�����@��M�͵g���z�<�ـ�QBd��ld��f���5n�X�٠}l��y�,,�DІ��Nf�:nj �&�=&� ܊�[��Hg�$!$���U��!L� ��ʡ Ġ;�*��b��l$"�N�32Fl��-Â�[�T)#�]cY����S��6I�H�#���1���� �p=��1Ѥ L+�&�H8��VL�!qA�0h9Ȑ$�-!�v�v_���|��	Ά�~��g$����܆�<T��>���k�83�$B$a�Y0��"XF�����%6��k玊�h��_�	 �0�B0�;!�;��N,�mѼi>R"� c4�,_���19(�=�,I]SLF{3���c�Zc�gs��,��'t�;��y{�������	  ���{;9.�D�G��Q�pG�O/E��TI�m��Ƈ�ղ�c ʭ�0��%��i�����$���iZ����l�m�[@l�׶iURm���f��� 9\��j�47h���nsT�;u�)ni˷KN;a�/T�S6�ۡ�D�l�e��0id�\Lv�rUT�Q�@�Ā�R�T��UW;��r��k�5�򱆮�t�nG�rd�{mۜ�na�'gl.[��m:�&���q�d�a尲g�h� ��mЫ�]������3`Н��d�5;\禗��ڭӞ.2XCc����t�>��)�>�!1�m$��_'L�ۛ�N�l�����L��u�]��M��Vj�[%$�b��L�:{)� ٪{�l�nYڡZU����j�ݥ��K���
� ��mSj�ڦG3��
���h�iZ���8�v:��Kt�5A�Ք���r�ݜ�i96*�o�-�6*�MhJ�WsOG;�U����(ZId4��pItں,{��v�r˳��88��V 9Vt^�Z��u*�KP�ޭm�4v�6�K��E�r��\t��6��m����lnz$�p�ۄr�ܚ@FKO�y�pv�ļ�λz����r��Z�ѭu<�(�iyx�p�zF�7n�`�.�����ڭr�^�Xj�Ӫ74��-�ݬ��Г�s^Y"zv;)fuc��m�v-���[�=�X蠵�κN�����<�ݳ�20񀤶�)eZ����!�:����WHHu,�����(��^U��X�3�8�t��7;(�PY��6$��9y�84��m�v�4��� ��[���f�H�1�=��d5��!�[a�Xꋖ����@8�Ձ�	ϗx,�Y��&9�Vۋq��h���8�R��3��V��3��d�v;
�v�nō��v6�ʃ�(�n����=OB����t�%]L<Y;Zh8�S3��
m�1SuĴ���`� n�����Nw�w����{�ǽ��'T�U*��r�T4)4*'��~E~UM 9X(�Aљ��8�Lb[q����|��#V���VU��j�M��ے�<;�0-�A�Z�yn�è��k�`��ַ�m�2�M;�v�d`����@��$A��=�4������y��j�9�v��\�Z����:C��΋`�3$q�G9��筌���W�b�ql�l;\:�%��#��zK�xk��s�V��� ޙ+�pW8v��Ϋv,�˸��E�zP{���wz�}���/];p��tdY�V��g��`����=�̓ӟeם&H,�Ӑŋ��$���@��v�kN���]�V����)�a_͉6��@�ڴu���٠�f��\�7n"�%��Z���[�Vr�M���`{���=����̅E)��L��&�ouX�uX&��l�2��Pem��Au����P&��l�&�'?g���n֍�y^�!�ҏ8�`������:{E�ٹ���]���-�W��1� �@����S@;:������߿Mւ���!ɑ1!C@��_��U(I5	f�V��V�j��8X7q(Ć��) ��f�I&�:M�ɰ@:�.�������������hl��vu�@�*��5�8!dCb�h�i`rKw���5n�X�v�]���#����dPu���\n����n�w2�oQ�����ܷ]�Ѻ���j���͛ ���D/�{v��:���FLP���h.ί@=�j��$T��ᕗx����+m�UM�fnՁ�eic_B"�"T(�W�*��ڜ���� $����aw �0UXt(�����������͝ �h���?�y�4Y�@z�9�����{u ��D��5I�@=Y���H5zF7XB�y.9�h���a���qÛ�ѓ����o�t� ���� #��.�\�j��PJ�lsv��$�=�\X����>]�^�تV�䈣m�Dksu��	&��t� 	$����i	Ȕ�,i8h�M���Ƥ���s�8���5S���ԓ�}p�aDd�	R�gW��4����)�r�I���&��{gEF$����H^���� ��d��i��,�q��뇴\���������m������c�빠[e4�gW�^�b�A�%nM�s@��h]�^�[l�/p)H �����@u�s�j�EH��]�B!���)˳��m��n��>�,z5���T��h&�T���X���|wW�,ٰ=�w�~�g%�b���x���@�Xa�J�K:��_G!����Ҕ�IZ��-��S��p�akGP�{m*?�d��c���.(���K#��A��k�=�Nss>P�ڸ��aA�u�l��j�9ח	�͝�C��2��`Wpnxn"x�Xq�m�D���	�J���m��:`�ݶ�qv�*�����։����8��ڜIA��'g@��Xuy�����}���hʜb�gd���ѱ��\A�qլ
����k����ϭ���x4J�	&���~T��ln��$���:pK!#�D�,j9��S@�����f��[��{�\0X7�1BFԂ�Ә�$�Pr*@I6s��6�O"2,y#����s@��h]�^��\l��b���7Pr*@I6�Nb �M@������?��u7��g�l��Y��Ņ��,���'N[�킶w<q��m�b�ݵGK�π����h�uzz٠}��h�p��;,�)ݏ�ܣ�E@�~�C
�5U�|X8��H� �� ��xd�<pkd�h[f��[�������u�-�T��HnBL��7"�EHs`��X����ӡ�d�D�D�8�����?�{%�� ���ݵ`n��k�JSD��Ƀq��X�������۴�P(��x�7:0��:	�0�`�B&(I��h��� �&�=$T�nln^]�,��h϶�̬ݴ�M@zH� �� �uhڶ48�X$��>�w4���{52`G.F*Z&�'�:�G� J�'�&������!ց�x�����h�uz�l�>�j�=��!'a�Cœ��<�9�����qR��@z����A	�"e�=�l�\p���d��6����N���u���q�]vNy�vթ��M@y�� �� <�sV��HnBL��'&��[��Ď��s:� �s�n{=٪4I��,n=�I�@s��@$����y]���!�Ĝ4?ˬ/�����R
�|}_R�������wK52`����H��٠}��h�S@����[UF��ډ���8th�NŷNV�xwot���]��� %ƻ2��i��K���n��e4.ί���|����P�ATQS#M�4������@$������s$�k�14<Y1)������@����;���w$��wX����������R��@u�s��WRQ�$�	7�@���h�A�t� �j�U�g�&`n�[gZ�l�l�;�R�ɶ:��� �'L�����&m�q����̛J��W+p..V*��)(z�n"���`.�jB^I�&�F�9ؽ�v
t�m�y�H\��i�9�eP:���e�v6�AΞ�:x8�0��;v"�]=���u����D����"�h�뺧�. �-��W/7�.я,^��\��nۤ�[>���_u���wx�<����[(�A���N��2f�,+Ѡ,��5u]z�,Y��$�,pKRf�o���>x�f�=���I(����Ձ힞B%�D��p�=�����@���`f�i|�D(l�o9��L�T��2��_߿M�n���h�������%�Iɠ}z�hl��oB� �l�:��"m���u���
���@����|c���&1�dj9	�S���)����Ѳ=�h��u��<v���=;�2����=%�$��*@9%4^I#9�����	���@f�Q#����p}V8��6	��V��M��$rD$���]�����b_�Ý�v�U��i-;�tƦ�ԓT�9>޾,����77j��fڰ>ݩ�!&�L���_>ʴ��h��h^��S���� #MFԏU�ٞ^z8;GQ�.LXĜ&V��-��s������׍�8<�XcN/�/_�@��R��H	�%�qa[��u{F^�t���T��qRvIh�D(l����ET��ɚV�zՁ���e-ߒj�T(jP�D@ F$�LK�*:`̇C�m�!c�&����hYXE),9��"�R�Y0BHH$,s�L@�k5r��S
 o�Ɇi�waQ0a(���
��z�T�eHC(?G"(�8����&�<@: `&���gP;��h��&7��(��#��_=�`�ڰ73mXr�����V�X�X��ic���@>�@��s@���h�ՠyuQ<��_�I"F-�9��m],tv�*��Gnk�.���)���g�JI��nA&�rh��hw]�};��Q�z@���`~\���D�mM��T��6��P��=��=��`ou��>���I�&(873@��U�}��g��n��۽j���\�&b����n��ݤ��#qR��H7�)"� �0H�@�{�wF�wu�dO1��,�ē�@��s@�����|gu���`c^{�T�N�3���^6݅�c��۞�]n�y�=Nƍ�K+�m2g�ƜPO�!ؐ�!�}�w4	�*@{��� ��x^>�d�T�iX��W�l�N�;v��>�m��BP��7�K�#%5R��`y����ZY�"&��֬����^H�Ad�!G"q��S@�qRt�����8P��2��4�����*@N�R��b7��"B�kf��Ԋht�Sr�Ẁ�Q�%q@N��G6��p����R\;(gR�m��F;q��&���x�z�f^���x.��&J6|Ѫ��l�.�Z��E1Yz�0��ݪ����.q-Sjv�VNZ���ꆲ&������k8ƽ\�ٰ�nԜ�"��*�9�M�� ���^�4m�knM��[q��h��׮��&��l��f�;��:l4�J]��w~��=����%\$�q�:��"���n����'c���������Mq(�n�S13&(8���g�@�^�@���h��5��I2`����!�|�\@y�� ��H7�@F�²�j�6��p��������T��{z�h�)@	�"��nf���3>��~� :Oʐ͂��HuM��X�A�5����u������n��ج�y"���3��a��k�����m��{Q�'�;r���a�!����C@�s@�u��=���DG�=�\X�4�z%�	�&���5$���m�"�"��]}�����t� �R�ӗx����D�D�����u�����k�4I ������$�%9߾�X߿Z�=���n����=m�G2`����!�u빠}�w4�S@��S@�lj�)��D�m�%ip�DQ����-�����T�?ٙ�ۤ�q����d�����`��{�*@Ne�4�luN�F�LҰ3r���(M�ݮ,��Vٕ��I&�j�d�k�jj�h�.��=�\X����� � DB BF0����	I!$�$��BB��
�!$�����7���>�cfH�%5R�STXr�ٽ�=�\X��>��hb��]�I�1�I����y���� <��@z8��ﺤ���u!Í������E��gB���c�=�Ts��8�*����sq>y��[v�@tx��x�=T��{��s2����RrMMQ`}���DBM���V�zՁ����(Pٛ�MˑTҤLKD��;��j��3mX�ZXs��]�926�Q�f����~���Ł�Nk�ԡ�
��JuC
�a��tjI�p� �BqDĄ73@��hs�h	$T��qRu8-�үsCr�i��YN��G96��[��
yq��Z3�y݆�a���?�ra1��}V���R��H���];.Y�u�Gۻ����R��H���Z�x�.�<Oj6�hw]��ե�	DD7��`{{�X�]˪�LD�,�I���4��Z�n�舄��{�`owM�R��)�*S$���;���������V�+K��$ � ��%�ni�YR:���زf��� �Q���u��i�s����d�KAT���W��,Gg4��xK0[<��n��^��A\�JYy�(+l�S��jP��k6ԥ�yX���F@�}��A�t��=�/\m����r��V,�8ݻ�\�]��-�dI�q�s�L>+] R�m�X8��؎��f��\�u�K�`:4l��\���T������{��C����
�'-�)���;0�^��O����*��Hn�%��Nx��fW�u��vU�͌�߭X�m�ٕ��"�=����zn&h�����:�`{ٶ��6f�~4s��hu����1$���*��ͤ7�@{�K@yȩ���Έ��_��XLjC@��ՠ}lT��{o`��e�NˁVe]nQ��m�=T��{�@{�KF߆�=���ۍ4-ͤ������[]=�ob�ѱ��0O9ЗX�vƞs��A�<4^w�H�@>{�@z8�@�é���ȉX�n{�7츘���k+Kۻj��ei}
I6{���[x84��� ��?u����i9��� �������}�EL�ۛj��ei`g����Q�6��?R�{���q$ڌC�4��3�ZX��vۛj��D{��rk
�陁ƎR��Ggq�wV{v �uv۠���w&��[Ӹ}���9�q����?O���K@{�T��M��=�W䐋	�Hh��~�nh�������BM��Dj}$�SU(A�f�I����w��N�����S@�v��^H��%�Bx�Q9�`nfڰ3�ZX��v��
"w~�h����Z�XcD�,Q93@���興]�����j�����>�p9F�=��k,��A͹��.v
f���r��Og��qe��D�6����f'�N�-�R7�@w=����t�R&%�K�vۛj�Bl�޵`nmq`o�u��M����@�J&[�//v������	�%�=�*@u��,ā��$�����S@�|�ԓ|�tjO"���"8�P�����ݖ#�c���4ϥ�'H�;$�o`��?�a����!Zpr⮭�,��,U�TX����#�.���Y�F����6��G�qh[mX��vfV�
!|�:w������BOj$�h�j�>��/>�@�u��>�u���
D�(��@z=�<r��T���ZG{  �E�$r��h���`��2�*��3
.��ݴ� 'd���{x�%P;�0ؘؤ�� `�&`I�����╥R�Q�.����4%#�$ 6�	�KI� PɁ�E�0jj�3\e�d�%$RQ�v鋘T��Čd�i�c@3��2��'֩!m&ڐ�8��2B����k)I:@�3)�a ���
4�,HɁе&���-IZ:��V�$L��`J�4�Eg�^��gw�s�'���8� 6��U�6�K��'e��9B��^���uy�:�٨���iP��yV��hx��ݥ���Zp
���2���[r�a�j��� u�����*��|I����7.+J��{[ U����c�-�m�gX]�(\��tM�\r��m��;����t�dcb�=(�[��^
;6W�@-Yˀf�Z�#^Y�FԚ�Ps+n�F�h�n�8���66�P��pk���-���0���&���c��۰Jv(�ڞ��:�L�����*<�� �z�n�m�=j�5U*��S���[X��sZ��j�``ێݸ9#����v=�㎮۝�^��HpmRNYu��:�Ƚ';`��65�Fu��U��7D��_��>HTn���5UZ1� ��j]�ی��j�iWi�&p��U��,� ^�ګ�h���V pN�dn{Em�TUɒQ�F�wP�l���m�ۢ�-��vka�r'Z����N")K���Q�;�:�<������N�:�V��kI�E^y ��\���QU*��WCv�j��mS�t��M���M��F�n�f�V��%�⭞bɜ	�7�!Gn��.ѷa�rlp���[�ru�K�֪�kv���X+n�ƍ��M���Gwb�g�f��@�9�f5<�N������[Y�FJ統��O-��(�Y2V���;����n`vav�y���m�se$t4Rui-��\��T���:��qڰ��U����q�p�Nȁ�e%��f�7K�-���`�m��������
!��78Z;E��'��|o���?=`���b%�9�`%Sv�n��.��\�r���	�ٯKcG�N�w%&���N:�*FQi�Ukn�-mU�T-[!5]m)�*;6z���ɈإE��sִ�:�zGm�������E)Q�Vm�R@����%e�0�w6�W"�0�8�1@sз�h�=�U�P�K���ƥ��Ы@Fk�#$���]k 7e��rF=��~{ߞ��{���~=͂):'�"aW`���r�è������/�H^O���%���F��H��t"kf0�cj��^�cJU�]��\���9��;���\��`ؼ����N:�@H̛[�]e ۠6g�q�Ϧi����,3�+�0�^I�����f��D@�1�u��;��iN�S�B��]P�ѮhY��*֭�w7,=�ks�5��)6IJ�k��-u�v��5�\kE#s�������7w�2�ƍ�^J3*������8�.W`w�v�7G�-ǉ7��]�S�&<oҌ��>����:�M����hh��1 q4ŉ(���x��RvIk���c�~!�H�1d��4���@��Z�hl���hH�I�<X�`7-.I�	�%�$�x�=Wք\���4�mɠ_;V�m��/>�@>�f��u�7�Tx8�$nG1ͺv��ܸ�rjM˝�KvmM��nIq֩��.&A�2�%�5"�=�)�}zS@>�f��Қ����I�g�ԓ}�{5��1�V�J���jlޚ���\X�Z_(M���"t�H��*h�=�֬̭4��>�S@�Ϋq���<m��UR�32��32��>ݭ,9D(O���3xu��l&��luE������6I {�3�׆��7I�7:�m���˨��j�s�Du��[G`���G��X��<���dœ��>�R��smX�Zt%�a��Ł�,l�ebT��6��nھQ
6n�q�wY��>�S@��+IX�1<i�&iX�,{+K9%��8Q󪸰=�֬g���I�j��i��Ѐ�{�� =�*@>{t��{���������M�u��;�)�}��:�J<Kđ���u =��n|ʼ��c��|l��M�������ڃ,�Ʀ9���빠w�U�}��>�)�z�T�lI�����@>�-�{�� =�*@s��,ā��$��@��)�}zS@�8� ���Q�SJ��6���j�~�,ou�=9��R�JE�,Un�d��ԓ|Ŗ�U��}��u�wy��EH��;�U�}zS@�h��H�ܐ��EPZ�&wm��ch^<ݧ3��[A�n6��Y���(��ډ�h��h���Jhz�h�eUE$��%�5)����������Os�3Ӛ�uU��$���cNE�}zS@�z��Д7�;��̝�`}���[H��.�74@z�L@>�-ݎZ��hs�K� ؚ�J8����r��`��H� 꾪�,��z��V�#D��m�mN�(S�ߏ��Áa����<7@K�+l�=����r�
�oj�s��Ƙڤ)��3�A�]�%h�Ga���
Nʼ�/�,pFvn�\"�m��u�$q�C������5Q]��ε<�#���-�����x�tu��v�)Н�ԴDZ-���wLr1�(��8�:U�N�f�BE�i��n=����v�m�[0�n�ɩOm�y���۞Rn�0���nYG]���{r͆��apm�����hG�@{�T�}�Z��6�3�T�MS��`}�Z_�	���j�ܝ�`{Ӛ�6f��5S3�5I�� 9��� ��vIhG�@u_$+����x�Q'3@�>�@��ՠ}�ZXr������5�9����5�wW�{����-��� =���*'�P��KQ���> 8W{Y���Vכ7����������R�j�W�����;����EH�`���-�e�yu6�����4���"�_Q_U�@wd���{�.t�1L�Ժ��`g���=��v~����mq`foZ�=�:�l�54���n�@{�K@z=���H�`��a�������JSu4��+K�%�����~4��Z���g�y�H���5���3dLd�d�	�Pym��{Q�tt�n�a�'����ǋ&$�4{����M�>�@�����ƒY���iy��|��r��`��H� w���6LY#Ib�8h����f���B0T ز�P`�
E"���M&�
�������S@�������#sr-�l�*@6�?\{?Z�/m6��&)��׮��Қy�Z��h=n���Y$I��O#��V�N1�R����]>�qM��^�S���1F�0J4���wt���}V���iВQ�v��7�\����m�zw]�6{���3��X�4��!��AdC�ģ�@������H�`�}�Z��t�/&���)�M��áDBO;{�`nmq`g�u�O��|
�Ĕ��)%]�`n�m랩rR��i��`>{���`��"������痍�1v��;s����3e��0�c���ҫx��.'gd)6�sd�al�o$��@wH�9���m���F�8�4��>�]�w6Ձ����I(l���32���)F�� ;��ʐ8� �� ${��E��	(�$��)�[�������(��O���`f�낚hjiӑ��TX�ZX�����;{�4l��q粴�ͱ6cs�6�e��s.[Fҳ��$k9*�W�X�u�����Z�<��/.���aъ .[�f���(�I���TV�P�v+��6�1/�6�N��ͯcs�{K��Gjz
�`B�O���g?X�]=�^ZMq������Ն�۴���ckeU����On�]ie�9�VV��
�F�n�Xjn��ltܰi�c���pj�ay^�?��{����Y�ƽ��6j�Qv2����N�k�ݮxB�]��&�7n����&�H�2!��nC�?~�)�u�s@-�hl�����<x�bI�@�EHI5$� $�ueݼV5���&h���)�[n�m���
���b$"1a$��*@6�	T�=$����l��iF�8����4z�h�٠[�s@����	�T�@�6���Ϋl��F��������Nʡ�ɦ��.����d�r�y�L`�`�<��d ��{�@=�N4�qF�$cXВ��LԒo��u�b�"0�w��I9�Jh���:�\0��lJH��$qR��@z8� zI�	m��Lj(���3@��M�[��}���?$�7�V�J|�&���T����fڰ:����{7�X�ZXo��������1�x��C[&.�r���u���ڃii�ϮZ�	kli7 17a.r�i�Z�"�oa����ʐ�?�x@$1H��n����*@zd���/1fm�{�Y��y��m�$T�꯾���(�z����b�HE�b��po�A�LAD�D�2�K�nh\�q�@�2�! H@G���A0)�'�˂��+���6C��	��z#ZHH��'�B��J����RN㴁��Y��>���p�� �A#�q �$�Ad�f
6�jL�&K�R���0 ���B�@#��8���F(:�0�`DXǒ�L�Y(cHcL�[��@�4�$`P��3��Y�}J\�A/�ٟ��	��l��%PH��1�b��.��0.�-C ġ˷���d!�]�]�J<�A�ک J�`k!�5q���jV0�13�!�4*iC#��-�l �0�5mΗKX�ݘ���c.�r�PZR��B?d�ό���S���H3M�)R�3X��DHD�bB0#F,@!��P��� ⁑Jh\�R?)�(hp��@㠋	������=0&�$��J�͚�`g�mX�t&޲�Ґh���âww���Os�37mXrJ�����4�Ӣ��Ku-�R�=rL@7"�o`��"�Gr��rk��K�ٳ���;\㳮�>ܧ&�q�As���7<q�������q�M6f�3+Kٻk�">a���`{�Db��$dc�ә�wt���Ձ��ٰ=����g����IE&���wD��*@z�L@s�R��4��%ԉ��#&%"Nf��^��;��s�g�Ra
D ��F 
QQ��U/;�hԒ{�;|g76\�U�������`��"���f��l��C�,�¦�5�6�t�/k����n� ��RXx�7Q��Ӻ���@Ƣid�����?^��>^�z!|�{zՁ��9ܒR
R�	�,ܭ/�B�I��;���޵`{�ZX��X̘�%Q�@�zנtqR��=��^������[q���w4{�4�)�|�W�{�LU2<��x�s4�Jh=����*@]Q�UWξ��P�Zx�:��l;��%�x�Ը?�a~��k�Y�c��(VЫ]!%����[y�����R�^á�cҐ�sfݚ�m�Vԝ
{Un�'�QC�]���4���n�Խ���Y���]��ҕ�y5��mzZ���QYLn=[�q����Ţ'��V������t�6ٸ�]�n�l�ڞpB�ge���k����}sU��\�߽��w���O���~QӲ��+1gq��,5�"N�\n�xy$v�˒ы�<L�9	�L	!�~����9�	U��XG7��煗?PhIO�'�z�޻�{�4zS@/'�&7!�#�@����@H�_I�	\ɖ�~JD���{�)�[Қ��z�w4�_�kk&��@��4����)�wt���Ǖ疌�щ�u6 
t�����n��:����1�ɼ�q�5����16�m�[^���M��4�ՠu�)C7N������76��DBT����EUWV��v	�%�'d��}(ڙxH
F)��4�)�^v��ڴ�S@�y��MȈLX���#�-;$�s`������r<Jbr-�ڴ��@�Қ�j�?g������ܘH�I#�,�����˽v �t崑r�/C��&:��N�.�q�Dj2#JE�����/t��yڴ�j�/Q
�47�D�E$4�)�^v��ڴ�S@��E��<7�h�զ��<T4�/���}�����z�)������iŠ_;V�z�h�S@�aV�ׄ�&�M26榝������Dv�����~Z���9xX�ys���AY��e5���0nQoY:�mi�.�8g�ڶ7��!�4�x�!�^�M��M��h�����,�&�P��@��� 'M�9�@F�sK�d��x��2C@����)�^�M��M ��HQDDb�8h�M�Jhܔ���P�UB�`@�JBa>�J����яb�SS)�7J�j�7�@I+`��6���ꪯ��?p/��p<ͮ_p�$�F��8@�
�5ض�'Eϛ'p�j�r[h��i	�>��q`o���76��
>a۳�~����IF7���@G6�����UUU_}vOз\Ct詑�.��;���7'5�ɾ�UŁ��Ł�ڊ�M:��:���㖀�V�:l͂�0Y�SQ�LX��h�Jh�`��l㖀����n��*�w~l,.�\�p\�;��7���ԅ9�6y������B��Wh�����Cu��{�$�n���U�;S��9cn�Լ �;u�rR�<!J�k����XBֺx�vϛ��ˎlvL6�Nzxv����`�8�F�n��u�s�y
���ۧ�ܽ���`I���B7Hm͝�5�%����;6��tNݖ�Nu��acY)9�Y���Y�\#t7'����;�����w~{���0�a��+p>��璖{v��9Z{p���]N� mІ�׭���pܱcRH|��S@�e4Ϫ�:�)���"xc�"#Q�@�e4Ϫ�-���}e4�B���H�Ȥ��y�Z���/���z�hmmk�j O��`�Z�� 'M�9�@G�Z2WFkǉ�J4�p�/���z�h�U�u�S@�eyʯ��L2"���y���g�[�mqd��h�=��g�nYNn2������,cP��&�>��?��h�S@���g���2F�#x+��I;�s�[����,�T�p��u���ե�������ǲ�i�,�E�z�)�_YM�)�^}V�����d�ɂƤ��'M�I�@G�Z��� ��<x�DDb�8hl��y�Z��M��h��TLS�����dU"EC���v1�w6�^�������K������O�qቊD�H�>�w��=�Jh�S@�e4�Z׃Q�?��@[���/`��6&�9h	
P�,�`��6�4�)�z�K-8����u�7�����V{[�F&8�6$���=l��y�Z��|�Zg���"1���%!�W�Z9qRv9hs`��W�U]���o���3�g���j�jw��2���Ç�����ٴt�v�dv9	ҽq���~��� 'c���6	��:��E1���RHhϪ�=�S@�}V�z�M ���Ǎ�DDb�8�u��/�U�[T��|�Zuf'�pR%0rC@�������N배D�k�%J�*R�(@�Ĥ�lB������͛�pjc'�
E�[T��|�Z�)�^}V���3����nE	D���Ўn �6$���[WckdX��3�3��S��41��"��$�M������^����hj��;�)�FH�6$榝�������;����\X��Z�\'�TQ4�F�
C@����R��hl����,��G���(�7m�^� �$��`�����U��Q���!�w����IF�}ǀ׼�����?DB�
�(����DU�QU�����DUʢ"������U�"� �E
�A �EF
�*`�E"�@UH*��TR
� DB
�P����
�AH� �DV
�U*��
�*P*U�X*
�Q
�H*T�� *
��� *
�@ �D*B
�D�� "�E �E������
�R�*�H*H*H*
� �EH*R"����� �D*��
�"�ED��  �DD`�ET��� �E�� �E
�D�� �A`�EH��U��
�ER
�F���
����*�� �@��D��*��"�
�`*��"���`�A
�R
�"�*E *U* `�EX
� ��`*X*
���"�V
���� ��E@��b*P�� *
���D"�`�@
�E�������D
�
�F�"�
�B������EB�H*��@Q��E ��`*
�X
��",� 1C�������"*��QU�"�E]�����TDUҢ"��_򨈪��DEW�DU~DU�b��L��:
�B
c� � ���fO� ��� d�@4   0�@PE��  P� (��@b  ��|P*��ET"B�	J� $  (   
@P
�BDBAD)
I*(U 	
IB!$B��  � A@ P �� ��XϮ�w�O'����}��� hl�ۛ>���ӭ9:w������=)�Ϸ�y�� -w�u^��T� �5=Ͻ���������y:�}x 0L��:lm9 ��:@ � PRJ� �V0 �����ç�ص�C���;� �yd�_w�{ּZU�wT�� ������p _O/v�q��p }9����v+���u*�glw��{ҷ�J�ξfy5Uc5O���(R�"UP( 
@���Lv�X�Q���4 �M)G� t�)�ΊR��(i�#AJY��OM JiJb��J )e��E14�(0= `t�14)�4R��
�cJҋ� gJPX�4ҌM(
bh�JP  ;� (�   �@e:R�٦��c4��Ş���Ҙ 7*X��ӼY���Wm�gJp �;�u��Y� 6���#���x �<�}9oZ^�y��[���&��y�����Ů��wt��w��� ���P  �( ^Ƿ�m���ź����nm�MϠ �{�:�ru���.�{<��� '*���__O��  ��]�{o7M�@�y�-��ů����{�i�w� zS��\Z��î��/| =!M���  ?�M�*T   D��R�=D` C!ت�6�)   E?Б��� ��	�T$F��G��O����9��_������;ܮ;�w?Њ"���/��*� S��*��"���tEV
�
��_�H_ߒ��FYI��H0�%����0�7�o�G�'bC�) ��J|I2:��p�R1�$�!rw�V�$7���4g�C8rCA�50�*�@���T ā2J������B*��#$h�����H�!�B) Eb
Ƅ	�
D�h�$ ` 4 Q��F#D0D�A�1X�)�
HF�Q��_�S����#Yr�����Q�&�)A��t�	��8��L�def{(��R52�������q^Ԋ���������*(���s�jW�[�)���j�f��Ϊ�|��s�������Y����ɧ�([5����u�&�j`sHr�`r��榢08��pl�c����o���I��(�$$����9�)TUB&�!#!�&H����h!q��r����f]��c�$����`jh�F��#HB�)Ns:R;aI&c-��K���X�V)	1.y��෽�0�&JD�fpũ
(����babC�.�_3�p�!�HmL�R0#�0H$@t��` b/�D�0!�#
@�� 10e�P�Ѓ�1B)k��U��E^jwU�̘�����zi�k;�B�ɒ���FHQ�1.9iLH�F4F�HԒK�Q�\n7����N���R|g0�H��˾�>��Q�����q � �d#�?E�;��t�����A2Ȑ#,ZÆI�fkBAD����H�ﻎ��u�L��kԅ!E�X�)��.�)��}�J�0��<�1��P� `�0�"e`2HՅ�2�,�3
�ű#��Q U�T�O�5	Z�-H��֤%�d#n`�1��sItl��H�J1��zp7ݰ��n��2f�dH��(�)	�~��f8t��|{!F�s��s�8H�I�V�D`0"H��X2 H!	V-R1�H��0�r��3����0�gN5ZM�!Lb!��X�&�B�J@�`0�l��w�7i�8+�bb�{>!���?2L���0�a
`��$L$"�),�ֻ�f]���!3Mj�5��2�!^�S�L�B�,�`�u���@��A�B@�K)ص1	,�ap������sV:�E�ir�Ȑ�R�"dJ�*�H�S	�᱉��&��+�SP@�T4CJU"iX,�!Z��� �CV�����"	~�X�	g�<>��ØcB<�s!�	��@� �E�d�"a�V Ap&�}.�I���HJ�2h�s���e	"��]c�fXF$$I��B�#`@��-pI��jr�ۀ�hh�ݒ�S�
K|�!GL�I����2�6[�wߴ��ֳ��ֳ���ZQ� � �ab4	 ��L9�$`��ߋw��jd����Le3
�d�0dHSJ�%a[����Me�O�S�"QX�B��.��Ig��cZ���
-	[Q�8��V���M�hMZ��]��s�M`��b��o�y>�w�rF��&t2���J`�]����p��~�Z�æFHB1���YA�	F���Rf�#L\�k�iBRġ+�gYfL��XU�ط=GNB!��|��i�>151���H�2\Զ����W��@B� Bİ �E)��H@�Up@+!=6��.5��%q�s���c�-{�J���i{�`��跔��	�R�}�$/��B1�@c��P����B�::}��o���F�@���H�R	"��X��[^���O���?�.���ή�����UPÐ!�0�aH$r�и2nv��"@j�F�2,A��l�.��0ö�$�f����ipt�	Li�0"M��$aPb����(c*B��,�Θ�C^�Xg����B<�X�ҳ��c	v9!q��
�C�s�L,�Mi��2B��0�M�`E�� �)A�s�u�&nQ�0K��Ln�*aH\I
�&(H�s9�Q�1 |E����+�,$S)�o���?Q�^Ju�kѵ��]QW_��JBiMT)�U�V������Z�U�$ƶp�J̳3:�3��t|p]H�"H�, �b!LeaGW�8K������0�Θ�L
H.�������pБ�F��B�$h�+
t�\���1�w8� ��+SĦ!�`A*ũ"By�;��������j�[mƳ�.Q~i�0Ёj¤)��|�����϶o3%�Ɠc$���
ci8B�$�;��s���(�;��3���id(RʑE�Mo��x�~��}��XBD0$������ ���B��}�]�~��c��:�vB�h:ˮ'���w�9�f�qӻ�=!pe$�XL$F(.7�.�\}��.��6�,�����������%��w߭�=��;/�4v1`?���տ8�T�Pj�DJ�-ycI
�r�ώ}��gF�\d�l$�p�"�+F.L�3Xs%ѲP�1+�F���� p`X�i���f1����f��.:�)X�XS�
�93א����2s�'s�$Jg��.4q9	�EZD�������.��&>�=	p����;���u�dM$.�6�֌dN�= V��v�d�a��
� 0$0��\��j��
>Wc�ՠ!�aC)��$�K�HXnә�*A��K+ ��Z�Ԣ�}��U&���c'2�:>4��l�;�;xH�+r�`3cC:|1�Di��������Ùpf8s�aĚ�;�}�a	5��9�E�V5#w��L��&~�6�����4��
0 Ē��>���B�	�i���Jҙ�����%�!a!BC3��{6	�b���&V4 RHԃ`�aO��K�k���)���C��	"@�� �� ���F	)#
����\K̡
�+��2�����6r�U��M���־�s��A  NQ{ΈI�l�V;&��5��1�����K��[�_B��Cx�����%��	�bP�b�s�p>>��lT���«��Ј���t�s�ob�9���{��n�0��ϭ���{��Oϝ�.���5��d�XH�Hp��8 �Q!YYa@�L$(D&	!H��XV�(VK���T"��V�2��F���D<I�C��5���L���c����<8sq>�du�%1l�>�u��1�Jg�c��O�7�P�p�|}��U� @�U0A�o�b�	L�u��%��S Դ�3̟vֽ����^6�=?o��n_~�UYX����5��6��e�Ρ�hɈ�4K�7;كX!i�\ƻQ�5�k:3.�'S#ÿ|c}�(D����y7q������7�C1�}q���#L!)�醓f�3۳�3����%)�x��s�n����	\�H�$B�[��@��m��%$1	
|�/Lު���_�I����>XMQ)����D')�@���U��"!A S�B��4�&fXWL �B$Ru+�\��FH1$� 55
B��!B�&1�P�,H��B���H���*��D��!�#$�	�����T�8bR�O�\�_�ݛH5GfV�`�K�n��e2O����zD��h!L%0t�
h�L�a��)��.a�[�P�d3�ޮDH���%0d�HR6�0@&HS	
c:�,(ƜXS	+�5Đ��(D�B�(���	!
"D�Y�q�SY�wD>3���(�r�A+ ���먿l���n~�.uz�,٭�3�c����nmơ��a2�5�w�H�Lj���v���	4��Җ�"�:v]�r�CWHi@�%ܡ�b�4֝G!1CY0$	��A�D�WW�J���jU(�x��*�@Q
X�Mܯ��E j��ý���*�T�  eL�IHV0L���bE��ȵ$E)FĲF�����rꏃ�TU S��I$�  �  �e�@   �$  Ŵ���   t��N����kg�rt**�H��,�֋o�Ԃ�� 6�+���\���1K�z��6�/]s`�%T�����J�L�S� *�j��@�ZP\�SJ:�N��Gb�6S"�NJ�j���Al��N��������Rݑvܠn����R�h�{6N6�e�����ʫpI5�M][lZlej���
����j�vSg�a�Ƶ�   8        �6�   5��m� U'�ِ���PQ�j��j��*�Y�1��n� ���o�>��f]�t�հ@KHnq@�n��m� s�6ݒ ��� m��h $ѭ��h3E�:,k\R�N�amÀ   [@|����; mf[[
�*�J�U@*�[*���Awg����2 �q��MƭBlʁ+WM��� [% pm� p�l m�IU*���UU^j��ZS-6Z [N׫Z- ���Ե��t���GI\����X-n�I���  ��U�i��]��؛l�u[ͷ^� ��J杧����^�N�k�W$p��Sm��p�Fg�����3��x�T�Lc�К�1ș�r���E6�3�8��<�mTc��(.
�q������;=����c�i�m ft��z�M3t^8m�kXŴ  R��l�-��ݭ:^f��yn���Z�iN���@u�
�e���]&$�[o 6����`�l �fH/Y:�m�Xe������^�m� ����r��M��^��Ut��b���i&��m6#�B�-��[�x���;Uq�AV�3[A�&�L�z�vR㬺K������6"%r����FH&���� lj�
Fn�2�Tȕu;h^�b��Zt��̹�յ)cg8v`$��s��n���ؓ[�	����Y�᭺[��4��:�j������;��plE8�Fk��	ӂK4�U���D$��kNZ��9l�;VQ�v�(ݻi^ۓ�B��,�J)[�˦_V��UIݛ�4*�V������m�M�N�X�v�q�wf�6
��;+��[@���9@6����� �   -��/���M&�Q����]�0	 p�����ٳl[!�@HI��m&m�H	lr�[m��%��y�[vۭ�JGm-Ba���n���  �[���p  6��� ���K*շ~/Ϙ��ejn�mUV�n���[�jcMNʼ�۶А5�X`uf�id�$�$� m  m��`6��nz�V�	`?�o��� 6�l <$p���ki#l� -� -����m� �h��k��kjvI�l�6�/�@pxH     $  @   � m 	 ����m� ']d��նY���,�` �l`�mp$ ��j�6ۀ    �z�#m��$-�-��l˓a��n� $��m�-�Kͫa�@$m�ے $ �ݪ�U@
�[D�K[R ���N  [Ci�['` ([��     -�   M�  ,]�Z�"i�  [Ku� @pH9@ � ��m�6�    �q��6�e�$      ��&����m�-�m � � [@v����i,�m���m�8 ��vپ�}��p�'�����     � $l����[@  l� h�$� l �� p �adZ[`���zĚv���DޓpM����  6���m�    �I#��Ͷ8 �\���P[L�N�j�RIC���   ��     n���  m�����m�ո!i�-6�jI$�  �  �   m�I%7mr�[������ �H���  8)vӱ�mHm�[%  ��n�   h ��ڀ �Gj�����m�8-��� �;`��l�I%�l�Yy����pm�` ���$6Z[��� �b�N��m�m���ѐP�  � �`v�e��l	    ֛cm� ݴJ�J�R�(
�1-4Y4�P �p/yzHէl�gKb�    ��  �bKh܂�ekA�� 𓄍�m���:˃ �۶� �I�Ͷ�5�[A��@�V�����j�g���[@m[  ��m��vZN� ��� -� %��ݶ��I&ӫbޫM�� �`-62��I"iX[`����F`H�N[D�mW�E�'C[�`���i��@$����äe/-][·+Z�d�K�d� \T��;t��k���]��.ٜ��D[@4��;v	t�L�M�T
�T�m)fmUl� +����kj�
���;,�%(�8!�ݻ=�@���m����	yi�Gs�o���W�Pl����R�`�9˻X���@@�{L���n�C��>�:*���6�6po[I�Ţ�(�2�;��|�^�D�v��J�m�mp8l[@8o6�t�8��[�]�m�]��M+ N�jU�&E��u��ܵ��m��e���Q�+���j������/]!2�T�*�KT����
�~Q�@��z��Z)� ph&�����Ci7N��$	'I.�[Eu!m���d�T�«�UUR�ʢ����*�Ij�n�m�zAm!��	ݦ̖�l��mjO���9�lU����wWe1���7)����v�cl�����̪e�=�9��zQ�Y�B��7K��;��%��m�0�����Ӷ:R�l��lKt��]T�[[e푧6Ĳl�N����e�,@T�J�Uq��y��yU���n�m�35U(�f��F
ڴ���K(i�-�ɍi��8  m�     I7n����`:D�K��[]R������J��5A�e��V�j����T�T�j�   ���������7"���t��4���n�� C���ѭ^M�m�\�8��[n/K( �^Я<�mWU��VꝶP��-���\�a';v�e��n�@q :�m�ف��a�ɕ9�ͺwgP<��յ����L;�3�6�v<�B��k���*���Rt�k� �UÛ�to`�Eѱ�Q���V�e�)VI�l,
A�;5QEvq�c+�iT8��e`��m�v��D�i~�no��;C�]\	�7����y�մ�ҭTkQ�C����%m���k6Z  *�.k.�l��U�.U[	��E�V�
ʁ��Hp�l�[lI  g��  �6��u��m [@$q�Ĝ j��]���Ƕ��]��cz�e�U"L -6 l $��#��a��l�N�
�톨gp��J�UK�9iVW'e�V��y]�zU��n 6�Im�큶��m�l	6ۤ:@lR���Z��UU��v�6r+Um+gpgn..m���@rZ��d�V��.�s(v�d�%Wm�`9�sM�   ջ �f� Hh;6���U��9l��jP�i�d6�p2��@�l�H��Y�tι�!%i�x�[���l�Ŵ�ְ 6�l� -�m���Ŵ ,�RK&�h�7�o��|:�d�9:8q-��+u�Z���Χbن�5�I�l��L��jYZ����ꝳ4�tz����l���ݮU�(��Y�̛/\(�Y$�.ԫ���﹎�`�7��F�P(�{l6����Khn�!��m%l6� �kj�u�[O���kn�m�	�M�YF�@      �pm�h��n-�����l  �R�  m�    :�- m��� m� 8[@  m�� M�z�� |k��m����������D�Qms�ba�n�h5�Q�-uQ��Gkӯ"4�.��(�$��d�[F�,�������nV-�9�l֛�v� ���l�L�(
�-t�UUT Zdu�ăZ�"L�)oPY�[im�mz@j��c`������ꪮ��9�iBm%-=��I�I�e	6�m 4�e6l�@�mWJ��(�H�]T�*�hm�E�Ӭ�m F�8	 ��e6��.��m     @ h�Te��Z�yj�+�]�T#6�� ��.�l�V�Q+����*��UV܎���� h&��S�km�m���m��۶�0  $��ur�Η$F�u��C�cz�v��#t���J�����^vm�u+m��*H���w�3P k,6�[wl(5����q���@+�,�UJ���ڕ�[]!!=@ul+ �[T�;UUA��$�5��a���u���w�}���h � 8m�   I��e��H  ����t�u�@Q\�P�@ H�   �cm�$   -h kV�Ce�A���pֱ�`:۶�l    ��* *�@P�0"�#DB*$���ʪ�ÄG��(�H�H�qB���CUD��cH��M�Ev�o�P\(�T@���>Z�L"�a� ��7��X�Q�#�S`瀶(;�!����/���z�p�{Ci�(�Nh�U�
 mO��E�@�S���� �P��"@�'":�h#���C�c��*<�����H� x�K�4�l�|��D᯲��1� +�U~@"��N(qzC�
mP��f��x �s�W(�������J|.p�I��EI"!�*]�	�� ;����G� �@�t��%A�@�"T�� �b�T���D����
/N*b�T&2^,�bD
F��u~r����;V͐���; ����[�b�Co�TW��&��V�E
*�a�>2���	����QEW�>�,�10�E����F�� ,D� EP��@�F��X�F�
R�;�����S����	�4]K��r#���3��E�K�������ct,�t�Kuٶ�m  ,�k<c-N}xyݝwg��5�GN��T)[gC�Rӣ�UeQݰX�=b�1�gT/l^eh۫�� s[����\M/:ٻcm��I�`��es�x�r*X�5;@m��O6�kl`���ձ����i.�D�@qm>�u��� �:-�H%�wml�[�M� \�Ϩ�4��{sV֣Eu����r�U�r�E��F��)�
yU���իo)ot(e	j@��
�6�m���-d�^4��Pl�]6�4$U�u�'d3j�����g��� ��9{pJQ%�w)UT����jy%��`��]��UT��+0mu�ؕZ�j�ڹ�`�� ���6U-6 ��#�����#J�UJ��]���Z��6�rmmv�iW]M+1��������2�"�M�B�I�l��m�	�<W��a��`\���T &���k/r�H㖞�Nul�"�qI�v��8���G/jnG�-0�M=!�;1�f.Қu�6��δշ8���U��)oX�"m�,�S�1WKr8�<��mg'r��̙k�����[;�b7dӤ܂����aޱ�z�Z���V��69��G��b�e%ˍ@�	����ոtʪ� ��0���8�Z�5Ź-�S����gM����'I�]u��qA
!����o#3[p�wGg��t��*�ke�`�tfB�&Z�����L"�(2�Q�$�qN�1#�P�fOl�6�ŵl��N��D�i�*�<� ��@qG��:�ib��U�1���W�a:��Uj�`�M"N�i,�m��p�#["�W΍�]nݚ�x�4����'9��v..m��h*�.s�Sgع�I�*W�u�*�\�U)G��v���.��T&�A�%���=	�Baݛ��6M�Mϖ硍]�fܬnv�iW�*��Pm�J���ꢸ��\ww�{���������{�)Go�����Q~9�W�"i��D؀t��ENS��q��7|mmJUl-����r@vnyJ��
�����Wb�K��8w��ݫ!ϝ�r�]Ċl`졨]ViU�.#��:yUkc�d�jZ�۶Z����
.�V����㎏<��m-� *Skϱ�J�M>(�b���{;+{{v��cr��x���rQ�@;l��	� \d�J�-�`��:��^ln���s>'��ػ{�wu�w�|y=�g �p3��1ܹ�><�U^T��P݅Ɍ�;���o�W�o�_<�{�s��Iu�r��n���q��c�n��^�;�۫�ɥ���6%�m���drL��$�s������e�=�PF�OQ#i�A8��6���d���<��c�V�5:l5�n'JL��@w=���@{�K@w8��w{��]����fy�g<��vs���my� z��������k��X�ll�n�p��Hp��7`s�uX�mՁ����ŢŪ
����$������O�#�2��X�\X{&�`n���$��F)BNH��6���s�v�������-f��ېq�BR9V{�K�ɩX;�,=K3}ʰ7���r��n��6��`{�˴ �M@w8���W��������ד���S��cX���4.֍�V,p�r��Pv}j*�p;<9N9��w7L�}�� :=���`s��#�Z�(���K�ͺ�;�4�8��; ����$��6c&i�uRꕁ�;����4�<�DD)�H H���D!z�Mjwz�u$�sn���jRT�$����`qw!�����qR�9hp�W7/b�A�$��wvX�mՁ�y���<���*�N�)!C$�КIK6���ɴ���\��kغ��cb9�ʤ�%�P��K�ͺ�:�5�ǚ݀gwe��ժܓ�jP��+�sf�6{gzf�7;����mX���ڨ��9(m��9�5� �wj�P�&�7�X�l�t��&U'L�H݀w����sn�������S]GZ�1���}��g�
��3 ��@w8��6<s1 {۵`tD(^��,��4���z[�-��,��]�,[�Ԍ���׭���G,Hr*�6�lI��q:R5%t���`sL��&�;�T��p�nmn�fiw�����3t���qR�l,�O[Q�� "H݁���`w��V~�K3�Ł�{��]�blRINdt�UUSa�
<���Ł�<���ݖ+uj�$����RJG)�6<s1 wI�� *�O=߿��>]Pj��58ێ�{i��Ѽ�z��6vy.v�h5�'���ѭwg�X�働Āu���z�5���4�����Ĕ�v%G ��\L�Ńk�w&U�&������⪚�Bzܽ˛]m����Ŷ�ù&�n���f��x:�h�ia�N0pO\�*Z��2��ţ FF�C�D�A�%~.��C,*J]�ɺ.9Qd���_��q�;�̼�rf�2]��3��mɓf�i9�\֞^b�I��8oV{�e�ѹ^k�S� �'و�M@w8��6	 �Z��&D29#vWw]�����Ձ���`qw4v3Ut4�ԫ�(��@w8�ݒZ�ܼ@u��`�fT��z�朧U.�XtDDDZ�UU�����1 ��s��oE���r�(
B�������V��j���i`tj�\��屩�T �L:��r��ji5�����j۫u�sy��y�^#`�SQ���i(
G�5g��{6Ձ��ӒJ!B��y��oK�LөNdt�UUS`{ٶ�<��1	�@�I<a#"��$¾R�T��ꯋ�����7������s�pr�n7*��=�9�5�w]����X����Ti�Ӓ���Xt$�C���́�;����mX��v�"%�L�""r%`b��;�T��b��]�'I��wr�ݬ��2��ZE�<�e�+�q�qǜZ+==�]��5�项
JSm�X�m��9�s�v�I�;��^{@�N��IVV��ɩXwvX�mՁ՚-$���P��`s�Z݀g�jȈ�������.�Ձ繮��u��ڔ�J4�ԉXwwP�*@t�-�{.�m��̟̽&�(RI����Xך�w&�`��`��=�J���#�4��xq��n�,vg]uF�uVj�H���#�֯H8�9M��`w^j�9ܚ�������sn���˔荦�8���X{+[���lם�`foZ�<�6l�Q1	jU$"r%`b��;�۫��U���Ԭtң������ѻ���qR�9�v8Z�����*��(��w�I'y{q1��$�sp��]R�<��6B����?�;���sn�����j��D���P����c��g��.���5�s��m�ݹ�pO#�i�E �IB7 �������ͺ�:����YM-��ID(
)�;}&/�U���R�7��n^ :ۙ�H�&��(RI����XܚX]����������
�j�m����� =|�����qRG���Ө��q������;�5$��wF��w��ԓ(� $pǸ�{�{����F@k�1n [�nk�WiG7N^nf��=9��:Bѷn2�ts�ɪG�'It�s����ϕ�;)�%+��
�ql�J�%�=�`:�g`��f�(�b�vֹH�����me�L�k���P6�c��Q�����M:��\��{N��u������'J�Tn��؜쳎��D�c`��zlV����>WR9#�[�Ny���j4�n�V�ڇc�����Ϯ���~w�(~�v.8��k���@��u�����=�)�=	p�ua[	jH�
j��d�D�}�,�6����`qfjv:V��齅%)���4s��1�@zۗ�}& �*M���INF����U�ř������6����դp�p#�&� =m�����*@t{]�V���r������ٛ�W �=�8�5;w��ENs�Ð���a˱�iM��jw�j�7V����t	�`�q�4�F����;�ͺ�=����f��	B�����ϋ&�TK�����LҰ=���!bi$D(PH% l�s�ˍv�RN^w���sn�����F�
���q����/�L@w8������(�5RA2I"v.��ͺ�:���,�N��lt*oj	Jm�$���qR�9�[r� ������鲝/P��J8����'-�&7DŊ^��m7 ��Ev8�.�\V;r�6���؀��/�L@w8�՚-$����&F�9�5� �۵`{ٶ�?f��6s��m��1��m��S� �wU��fڳ��LF����o�ɤ-��pH�%-�)b0�� �~tJ"�����XBD�����ѵ0��Q-�!���G�� �cI(��L |�>0N���9(� ݤ�@��$�1��9	�vK!l1���tL&	P�� C+	\D�1 Lk�`a.e4[�;��Dj�j�/�!i)��m )�Wzx�S����� :2�������E~K���Q��w�>�`k��6<͚��i��4�$ܒXyfo�Vc�+��\�~ID(�߳��q�4�EM)�3o6����f 95����?{����:�K�67Zu�M77��k�n�Iȓ�,4�m˛ZV�+.�k�磨�qÀw^�� �n��ͺ�W߫�7ޟ���)M�/�mT�L�H݀}��}��֬��v�9�7�/�d��?|���J6�"rX��u`ufl���gzf�=��`�Zc�5�Ъ4��}T����׾n�9��`����p��X� "~O��~�'/����R1AG �Vf�`e~�����US}���~��8��yߒ��r&��V��8Ui΃��::�5��xuq��;f��N�ݛQM��e�9B����������͵`{Ӛ��9��^�9UN���t�rI`nf�_��3�XY��s����$wƓԆ�J�m��Ұ3'����M��3;���޵`n�
��Q�M���|��~J�ǝ�`nfڰ�;o�w�)���MS�橻 �nՁ��_��yx���Ձ�ɩX�V|Q[��j�"���ں���{P���m���.�Q��J[\r�֯qkm�H��>]���v�A��ݺ��h7
�L@@���*�¥����[��)Ҏve��9��+�8ݿ��_�{p�qc�B�@� ��J���ˢ��k�;x�*���<���e��t�͇���F�e(��v�g�xS6�d&�|��5�Ѷ�@��ͣv:y�jh�5R��Nv!D�QW�̩%} ��g�l�v7a�Ѻ�l�<Yxn������*k�L1h�/�չy_���]~�߷�X��V�+[�k����1��Nhj�����nھl�N��{�;�ɥ�զ�rT�PJI	"�>�����ٳ��mq`fwZ�5�k4�I(HN8+�����ri`w��V:�E`e.ᮤ�H�F�f�����*@{�˴_I���c���EN��eeW8-�kK4��-�����,���T�ы}(��=����:�;L�UQ��֬�sG`y�vB��м�}���?~���\i!��H7�`s'4w*�ZJ#W(��w����q`{۶��/�&O�Τ���"r�rS�������o`��R�-��~�RQ�����d���wn��sGa�7��V���̊y�Rkp���"��6|_���@s{��{��m�s�jy�l�v��lU��r1ؐ�Z�!��_\����v�n�e~}ބ���F(F�j	�]<��V�����NQ
#��֬�a�"W�J�U `榇�����DDCfn�������B�l��G�䦩���&f�����>��s��J���XD�6r
BxQ1f-+J0)i����
�w��]I'=�f��D���5)�2HX{廾�X���}��a�7o�{y�2�LT�A�$���E`{�}�N���36Ձ��Vt��)S"&�����$���il���T�Ɖr�etrqGuM-ߟz֣J����I�I�����;�4�33mrP�a�����=B'�S��2S��ٕ����(�;���:{���ݫ�(��v�hs"�E'T���5V������С&�wuX�|��5	��Q���'*��U.�o�=��`{'5�y�Bz��8J>���F¥в�y�����eQUA�y���I5��n*@y�h��U}��z�<�����8�i��jP�k���GuQ��Ӣ;�N��V�LlG�� �T��JrI�3^�X��V1����,��$z�J6Ԥ��"�33m_�����{����Nk�3sSq��n�DӒU��y��n�YС���v���sL�=��L��᷻��I5�����_�G�ξ�;4����2�JsU`{'5��!(����y�� �wj���,Q�*�1"�BP�zf�E'A4ꪛaR�UVV�v��4����P���-x��Y�i�#r�lQ��c
;]:��lm�NҘQ3f�&�IM�#_��!��4J+�W�g��(�탶�=��v��G�m���@in�q�j��Ng��0=x��@D�tm�E���|^��!*�t���F��\ ���c>�/c:P%�=]�a�1m[a�؄�u��k#�6�Z���{���������p7#h��l�.֊���d����^�ۃ[��y�N�]ftn�#�4�Q�u!^=���.�`���_Wf��1x�i��ERTR�4���\��J!~P�C?~�V���`ffھQ�/k��L�*�H:uNl��V�s]�	(owzՁ����Kb��r�������$��������֬�9�6�?OwM��4��S�Fڔ��VfmՁ���7���{���<�`fejn��*t�ܐ�\.�N,Eǉ5��Ky�\�O1s��:�Y��=�j�)q�CtB&���q>{�6�s_D|�wzՁ��2Pt�dC"r&�$����s+�W�VUU�&�Z@�*�ZPB�<�����Ϻf�m���_|�~��&o�Sm.� �g�:m�)'8�Z���I%�����������$����$���'G~�sՊO�}��{�wݮq$���ݤ�\���$�_}_U=�~j�Ic����
F���	��K��6�o���g�߫1��z�K��y��/�`x��~�e��q>:��n۰fP�۵[z|6�l�u�f�y��p��~�w�o��g�T�*`�#O�$�}�Nq$��֭$�fo˔$��m��t���x��j[�ES`ےNq$��֯�ʹ�wܮq$�\�N�I.n��K�ie���8����s�7�m��=���3�A4�pk_^���w�m�;�غ�%���.J`&Q"M�%s�/S͗杤�]��9ĒǓZ���ow}��K}�Ruct�"��i$�7vs�%�&��Iff�Ē�I��I%��o�J}�v�`��.YNL�l���A����Ƿ,�^�V਋c�h�ٻh�SE_��KM�����s�%ܓ[v�Iswg8�Kv5I�3jHԥR
A�I,��W8�]�5�i$�7vs�%�&��B��S��)"��Pܮq$��jN�I.n���m���$�����$�[���fq爠~�W�����������-�9���۔���΂����������i$�O7΢E8#q)�s�%�&˶��(_�]���cm�����m����8�Gk*=�A�Bn��R���B�F�y���x(wUf��z���Y��������jc�62H�In���K�&��$����UWz�Z�y�I%��&�L#I�9Ē�y�w���i.�ޜ�Ik��$�f^�窾���ވn�7N�S���;I$��zs�%�&�i{�m����K5�4�$�;PX�ҭ�E)�sns����W����غ���{����~�&��%�����Ē=��i�?Q#R�H)��Y���q$�U~�����>���߿l���;�j�n\���@L���$FR$BFI�KHU�"�L`�Cf*�2H$P�^�!@�	�V1��K�����.8�Xi�8U1pR @���,��H�}
�ʥ�!�C�a	`�%	V�ѭ
ev@�a8��bAH>H@�$�t$d�E E	I]}�!`DE�a�  D# !�	F0#�1��`�HI�F��$H�B+$H�"@"����$I������xe�I$a ���!rJ�0B1��$$�@�$B"@HF0���$$2��(�5�A��H <��?����U�i�`�#�l��W����H�]�Z����	א�+j"�U�j����U�Qyx݋�ez�#=׮�v�.�I� �Wf.f��6s��م�r&ʵUP�ԛ��˦�N��Ӥ�]+$�����N��v��E�v�1Pum�c�D�[#i�;9X-� ��Λfws�Ϩ��pX;�h�,l��p���͖�{v�ZI��R�:���u�՜��@Y�0[�熶��-���&�?���|%mƚ���˄���3E��<�U���{dS�Ч[�.��EPF5`�k`n������]�$� t�Cm�v��	�
�s�&x\���MWb$�ٗXlJX�0m�ۗ�LHn���� m�l 8f�>�����8��'��S(<V�X!�5vq4<��=��ݵ���  �VYwK*J���UT�ԚeH[�����[^���vQ���W��+UY��h],��V�̪���x�i����(.�j�#Km�^��yZ.�C�v�{\Y�'Y6�n�	خ�9�{A�YH��ɵ���mQ�Ú��%��T�C]��c�kc���F�P��v�0��Ϋ�J��C,N�f�%���w��	h�f#f9k�nC:)]�i헆��Ӄ&�C7��a,�����?r��øyp0L���4�]a 7��1��5J���>�Mb\�V��ٹ�2��Q����kz��1��O:��n:����l�gF�a'(��[{I�>őᮀm�ȵH-��x85ɢ�Ij���<l��[���'�����&���ʳ������U2�rh3�V�Tj^�qs�%��&��n-tu�S��j�vn�z
��\���2p�*�^��֪�( i3M�u�e2@ @ �Wj�Y,Z�j�qU�W�8�U�ʋ��I m�����x� ��k��r�"�w�,�:��#�F��n��7a��D�d�nv�4����@0k����2�M5%�j˷�&ӛ��Xxۋm*�h��%�o �α�Q&�Ȋ����>Q�C{�]y�8S��.�� � Q~��QPf���a�mH-���]���ev[�#`���kq.��a���ѱG	��u+�kc�Nu�l�`t;q�&�I��ѵ��)���q�09�v�����n�ms�qj��_N��8>vS�x��wT)k/\�B�L[v���g�u����a7oJu�=�cl�e�vlnR�*;N�0����� ��rZ=1��S��l��6Ck�Q��=��{�������|��;vyݨ9v���TG�Iˉ�Hxt��o���Y���t�β�㻙�.��R��{�%��~i�I.n�+�I#j����Kw}��H�lg��)b��$�sm���ߗ�Q�!US:{�m��߾\�Iw֝�����S�^(�8QF�m��H׾R�In������m�杶����~P�^���*e\�C�"dr�[o�g��߼����f�\�m��ݛݷ������:���w��3���9����ͷ��sm��"%��^�m��ZI,��W8�X�������(��kɲ�r�c��Ӱ��Φ5����6�����{�|3�Y9�m�5#� }�l����q�m��{��~s6�߭�G����� N�q��KUߟ�m�9��Y�(�� "H	 ����!�*+�V�6��sf�m��y�i$����s�UUSm�i61���J��Gi$�}�W8�]�5�iz���y�{��$�׾��I-ŬMl�jF)Br�ė���l�4�$�{��s�$�sjm���U���/�m�~��M���ӌ_:D��i$����q$�_W�=����Kw��s�%�sZv�K3k[�J����k��<�Z�쉛u=�;X+1�RZ�m9������w����m<�n� ;�w�ƭ������~�3�\~�H��߿r�Ē���7WN$����F�m���vo~E1�^c���5m����om��sjo��P�D̷���%|*�)�؛nJ�K�&�$�ww��.������ y@Q�w�׳�[m������y�̘�n)�
c&&n3��j��_ʊ�=�����}�{�1�m��{�{�����I.�[e$�Hj1�	%s�$��m��!-IBY��������3m����W8�[���tm
�t|D4 F Vuֆ����x�J�j��Za�w55�h�_��w��s����r�9o�$�}�W8�]y57i����.��^���gzf�m���9}D�F�b�'+�I.����W�T�K=�r�Ē����I,��W9������6D�_4ԉ�I%���\�Icy��^������r�ĒǳɻI%ǘ�
�
,�L��M���Oʆ}�{�1�m����7�m��n1�o��SJ�x0�Lw����8�Y��Gr�Q�P��#v$�w/Nq	{��m�7Ē[��+�I,o5�I%����:��FAE��̦zɡ���e�	y��%>:��Kd�����5�p��UD��rWz�X�y7i$����q$����UUU�B���W�%��t��aJ�D�I�I.��+���UU�mw���<���6ߞV�7�BP�e�aŪI�z�Ԧڄ��Ē�]��W8�_W��͓�;I%��r��$�cM�OA�m�U��I{������\�Ig��n�Iwwy\�K�_4�|夒^�曧�b������$�vMmؐ�}_�����p�-�^��3�m�w�ٽ�jr�Ý?�����lq���t���ѩa�FI�2$�Z#�#xrtmCָI�	��<KR Im�e�ն��H��Us�J������>|���8����I��w�������u��ڶn��-�j�B��F�ôMv����aф2��n\v�net;tW��ؠ�Ä�{x��0�R�i��Ѝ��>l�8�4<'<]	���4��+��{�ϑ4&��+
�m��%�7���䎼q̊A�s�*�xq:��V/�������Qq�R��%����|BB��-$�ww����i,�������~ɷ7hb�q-ߟ�	w6KI����K�&��$,��W9���k<x��"6)I����I%���\�Iwd�ݥꯚ{��+�I$�}%����l9>D5I�\���瞻�n�m��|��fՇD'���3M9M��H0�	���vf��
?B���^~�u`s6kV1�h��6e
l��(Yɸx�ۥ�<��/ŧ,�=�]��A0�V�/�|�*$'Ut��6�$�����;��V3f�靖7}�}��c~d̓HN�UX��Wj5!%��K�.ͯ����֬=�W�$��
d?w�e~��H���=�~j��ݺ��|����{޺�7�&Ȥ$�"H݇��"{�~���V�vՇ?o_K�:�{Ѡ�DL����`��`wdT��2�ȩ �˛�w�S�ڸ�	ϷY�f8n�n��V퐆&i�-��S�B��P�#b��)�' �{�V;�Z�37n��q�����l�Ј�J8&���w&��6o�~��5{ߝ��ݺ�?W����T��8I	���V�f͎�$	Bc�[
�%I8��<p�ꕷyyu̽�̺*�X~y;�6wu����s���X�F���c�Sq�`n��X�����zՁ癳`~K3�ʙ�\�7#��Gl��ծ0x��lv+[���[�u��j\\�V%%�՜P6H�w����\݁��j�����0�����8�)���(�J��ͺ�U$b��;���>�V˿��Тdַ��)��n�J��:��`k��6�V�r�o۵�������k�C������v�D'ݷŁ������V�BIL��;��6�i�h�	�8X��v���H�� ${��uJ�e��<��]���ڶ�X��:�v���7�ت{<6p?��{�3�|8��m]��i���~�`y�l��Zt$�|�۳�X�ڃt�xԦڄ����w��Cgv��k��7sm_���DD6{���`�_�����;������ekvt%	&���X�zlsfI��Hꛚ%�*��tB�O۷���֬��v��V�kE-dR#�J*����VBP�wz~�{���ekV���W;AFk8/�ܻDqH	�$�ڽ����X����.�p���Σ�l���s�웗bwN[l�]�$ma�����ʖ�;�7j��J�����V��	�-;4�ud*5�s�gs���_v��
1��B�&W��v�z�Ol��J1��u�aڶ�ݛtN�æU����g[�F�"�����m����U�d���1��� �G��O.�p����%��w�M�2]�^���U�k-�s:�n���N�I,X�^e_m��ߞ�{��}������!J7+@�������U��ɭ��;��X�N��M:r�iL�$�M��;��(��n�7`wwZ�<�5��#}�L��4�GƜVwg��7wmY�C~��vt�;4�d��D�
�]S�nÒ�}��+�;��ݝ�a�!$�BQ������ru29_���Lˢ�����5�	.�����V��Ձ�w�t�#���$�Ci��Ɠ����]�0=p`[�8�:���ftn�Q����Q�Q�r.�����X��J��ݵ��P����v��-��R�Q8ͷ6g��o����#�T��(@��H� ��� �aB���#�T? �������=�����BQ�f�q�-��j�:uM��֬�9��Д%�Q
"g�������_��<�n�nSu)�*�:��`}��v�V�����:!BQK��r������ ��&����͵`rID/g_7��֬�9��������1�.j���'���I�N���.����ħ8�����s�O����a��yL8�I%p秒�73n�u�}��q�޺�7ƞe�>M$�8����j��Ӛ����mkw��IL��.�GI��q��I*��~����Ռy���re*�B ����0�"F!8&�<8*m >�tȿ�H�4�ɧ�rF����5Se�$��D�u�i����v��#2R1bBRA%�m�'�	���C�g!��\�4J��&L��lK	B01$$���`�ql��)��;��T0S
��v�L� @�!	 �� �0.�}~Ew�y�4���D\U~Ga�C�T8�k�� �6� ��v���Qr�Q<���ϭԓ��]X��i1��M�Q�r+|���R����s���r�s0�&���Q��X��J�����p��+s&��[�5��l	N�
.����e-ص�>�'6]��Ş���gq/��R��JF�T��]���u`uw5��Z~J#��UŁ�N99E4抢�s6�|� #{�V�:EH�6�
F�c��%G`nd���V�tD(M�wZ�1�����m̩ґ&%"�9݆�w6����k��}\������ڰ7�ˌbhdQ;ݼ6�H���b9�@{����������({�sd�h��	l�SƆ��m�ݽ�<��1�Qqώ�����J��|�׺�wa��{��Ձ��I��169G���׺�wa���ݺ�;ך���͉�9	%
28���`n��Y�K1�?yXs]0��F���"�����������=�������k�<�hI��8�E(ܫ�y����ש&��gn���;�RN��e 	���{&]�jآ&S:.��4����8���bYF���SIzV헓���=�sV�k<�e9�4�g�kc��H�@΁��L,�ĸ�$�{Q��d���^��2��$�.�uo9��\Z�;nG(S�N��\ۣ�b����n:!�
W��F0
B���)G#%��M�F4��j���ҳ�H�˞5k����f�� �����{�����wӾ�t�xD����*�Δ�ck���.���-�	[l�#�w1H%�>|�|灻.r�d�E�w�ߕ���5X�۫�y����N�8�)n)���5_Cg�zՁ�;���Nk�I�xӤ��4�ȢjDȬ�}u`uw5������7�~������egʦ�m��q����@u�}�Z�4����}��Ԁ�j��i�ԥ7(����ɥ������v���ٳ`nmJ��M9w�2�fm���8��%�ӟ�o���oD��q�¬.n�b�\�6���޾��͵`{Ӛ�BQ0�������UNf��N��,�6��u" ��DR��C� |�.u1y�cRNwg��ښX�	m6�r7Q�%���ٰ=�,�
!$߲ys�guX�-�(sHrM'2QUSa��""wo��<��ٓA��'��l���m7L���pN��X���`��<��6�fՁ��Z�v�JR'D��avQ�Kh���Ϋ\�	Wk�!ں���M����UJq[�6ґ��n��o�����l���]�������&��641:�I`uw5��M,u�j�wv_��H�j��i����Sr=I9���RM�����e ����rXY�v��bhr� �IA^��d�h�&�:��A��"�@f�j��Q��O��X7vX��<s��M�@{����&b���n��k��Xܜn0:Ӧ���ض�m6x�	��l[��{��[J�EI�����?��`fei`}�կ�~��G����X����%(Ӕ�!$vfM/�_U}I����=��`y�6l��6�b] ӑ&�p�9׵��9���UUURX�|�͞,���:WI�$����Ô(�߻z�y�6{+K"�(J�;5X��$D")���I%���ٰ:""76��gQ��>�ڰ6=-~�M�`�v�92ְ�Z5��U0�闡Z�n���Il4O���"켟;]0܏�nl�`s�SK ����\A�7��=�~	�MA)IHX����~Q
�g��V���`g����"#�(J&M�C��%:s4�:j���ߪ���1 ���[�	F����H�G���=�WԱ����,wjia�%�舞���l���s#���sI̔UT�ܭ,В�r�>^wM���ٰ=1�TB����(ڟ��5Tʥ�u�c���:�޶!���}ͧS�m�2N�헴���ǜ=�y��XY	���w':���`ì��9k�v��+��6Ɔ�y9�D]�; xU[��Zь�ض�޴�4Mɇ]�����	��v�`�Xս����u�<��/�k-��Wi
^6�'�Z`��y�������VZ�X��Js��1�ؙ6�>�T]!{!�绺{�}�ߧ������!��К-��v�j0��i���A�9���=Y�s�Y9Ȕ������|�ci���i������ ��_9��*@ewE��V�crș�������|ُ7��������F��P�g�J�L�E4�6G`b��;ݚX��U����`f�i�LzȈ�܎á(���Ł�\�?n͇�$�芯����`�?�H�i�MA)B��=�*Z���_9��@;��sI�1].���gv3{h�k���ώ9�֞�Xܺxq:�w+���g[������OS�y�6��f������#���~v�?����u������]�vR���F����
Y9u���Z�?n���#<i��$�nRl�����,�:���!�y�6<ޛ��mܹ��$G���<��_���o�����k�����}�Ł����M����G#uN���ٰ?%'7��;6��>���`o^�醰�N�Nm�r8��$p-��л��ٹ��{/k���r��.ߞ�i��)Q(Ɖ#��|��M,u�j�5w5��cLO`�NI���M/�6{'�;�oM���پ��sg�q��R��JB��?W������U�#:�-�T-`��d2R�dU�*'A�&���{�o�����
zӧS5S10�S��_�����`k��6�+K���s�9��#djD�G�������w�~8s��1w5��Ţm-M!��*8��2q��W�5����q�h�W]sն�'��/��Ed.�$�6Ԥ�	#���:��X��������m���B�9uSE���V���%
d��l{ߦ��vi�#k</SbWL��J9��y�6��f�IG脦sW��͟��9� �6�DTJ1�8�=��T����ή,�:��b`��EB�KaD8���������{I4����綴�?$�K�P�6�/��k��6��g������<��湢l����7m�P띬�m����'mָ������3�&����IJjB��^֫s]�������f��V�y(��2�R��V��j�(Pُ7���mq`}�ծ�D}UUIU��6���MEEF�,�M��eig�7��9��z��4V�#q��&�I������^֫ �se��X�|������"JF����K@�5��b��~�������_���b�@1 İX�م��R��e�c�xF���q�|k!�]� �&��bB+!"@�����D��
o�4�kE\�
��_Ws�R߹��#��5�i�,v�b�U�-�0g���	'5�t�1Y�4����!Ǜe�Ƽ��@UP6�m%ݦ�<i۶�v۶N�U�F� �K.�r�m��L���nW�Tՠ`�������3�8�+�v��{lr[(k��(s��@�;
����i�у���-[�Pc`�I��:�s��g���s�"����g�mն�\�us�s�e���N��R�*v�Sڥ;Q��ۇ)��݋�.z�Le[k��.�ǳ�g �26�:N�'Ur��t��؎69���m��*�9���[[*���-�mǶ�[  d!�[[GHlk���Z����ʮP��{`\D�+";��ge�U (���tT8��!˔ s��²��A��B�5t��5UF;[AKRݔ��)���!��Tk�nM ��1� �6i8�Ͷ�� "�ͤkf�V�I�$�2kw+����::�)q�/;<�)�ciV��&v۝�ɛnՋmX�-�%q�.�M��N��)Y�wR���
Tt�Zt�2\NY�G�BLˤF�Wj1�h�Fx�w���k��z'Q�[ך��9\q�k�5)N���6Z�9�:3�h�b��!�u�p��ιWlp�sTs�]��d�:^3ؠ�gkk����mӤ�/�6$ j�
Ŭ��a�m���۱K��b�M���ݵ��[K��6�'��95"�S�X�xv즂��t��%(ְ�f�İTm�"�Q��vl��UV%W�/E�J�B�C΂u8�"�Liֹ����*����18���p�.�pZ�$��vF�%�a:�5��7$��h��=����x ��s Y����\誥UU��CmUQ�iT��;(=FT�8���Z퀣	�m-��bf ���1p�gx�06f�����.�^��Г"6��n�����;0̈́��������m�̱�k-5GRk<���˛�V��7iVy�F��8v�
��л-�[MΊ�����{�׻�=��	�v��T�E
�2������|�E�p���%��w�������e���C�5)/8�Im��0#Э��a�x�5s�v�m�K$���T� ;]X�8����VJ��3ų F��:�c�˰
a�;-v͐�a�"Ns��YصGc���pF�0jwWF4��	њ��84�ps�� o$k�
�ñS�H���Q7�%���r��{!E��.S���mץM�g�����;�y@�*��w(S�%HM��L�L0j�`]��0�R7mM��FS���5���ܘyAJe7"Qș@3we����`w2i`s�kU���Z�"���iԎD_9�����R�����_�Uپ��hb^��r���X�<X���`��`w�5X�N�q�:j
����Rb ��P㖃�rE�`f�Zj*�9Ltc��9�����wπf��`sY���*�l�4��-Pd`N�v�m��L�L;���c�1qڡ|x'��wχ��BGn��ͷ���=�ZXl���"|���U��Ǌ��	��G`w2iw�}S�Q�"�wuX�uX�vl�X�'"�76�p�6�� ���=���^^�����Ł��ZƁ]1�D��SU`f�X�vlfV�
|����U=)�����i�RKV�B���q�Y�V�nՁ噲�f�]����N�9�V+�#t��vr\���0K\l)ڴƍҖE�����������5n�X�ݮJ>!2!2OwM����L��O���J���*]�.s4��bX�'�=�gI�~8���%�~Γq,K���߿cI��%��Y�|\/��Bd&BͧĔ�MM)1#�s��7ı,K�}��7ı,Oc��4��c�0B��Ď���Lg���n%�bX�1�{Mı,��������JhH�������������&�X�%��{�M&�X�%������K���D�;���n#!2!g���}2:*�GH�(���_X�%��;�M&�X�%������Kı/�ﳤ�Kı=�{��n{��7�������^]��+f{/��	,��v�4ykj���!,5�.sղ�Ğ&��.�&jjh�_�	����t�/��,K���:Mı,K����&�X�%��{�M&�X�%��z�L`��1�c37�Ɠq,KĿw�Γp�D�K�?~��&�X�%���_��q,K��{��n%�bX�w�׮ubwD����w���oq��_�~�Mı,K���t��bX�'�{�Ɠq,KĿ{�Γq,K��;���b�_�1�79�4��bY�������:Mı,K�߿cI��%�b_��gI��%�����J2�	�ă��G�<,Nn&{��Ɠq,Kľ�}���\�e�͸�t��bX�'�{�Ɠq,KĿw�Γq,K��=�cI��%�b^w�Γq,K��~=�ݘ��$y��C�r�v�/f�-Gg<����7VNl�t:5q������|���Y��������Kı9�~��&�X�%��{�Ɠq,K��;�M&�X�%��������oq�߯~�r	�j�{�ı,Oc��4���"b%���_��q,K��c����n%�bX�c��_�	�������U2:D�Eg8�n%�bX�s���n%�bX�1�{Mı,K���:Mı,K���_�	����m�:������3I��%������~Ɠq,Kļ�gI��%�b{�ﮓq,K�^ݾ.�&Bd&B��9��-MqYq�i7ı,K�{��7ı,?1��^�t�D�,K���M&�X�%��ﱤ�Kı ��g�\&r�l����u�]�иȦ��V�7i�u��ڮ6*sZ�[f�ݰȍY��X�]T�n�cn�v�ȏd	��� �<Ö�*�Kcm�k[!-[v�����	[dUv����0=�6;vѸk���q����n��׭O ]=�kʼ�ヒ�[:�1B��� �h+`3킶�㍱��Z��9y��5i�p�6���C�nã%�G�tR��>�J��;e�E�y�nΕv�nB�O9�q�76B��ۦ;M)��n+7:'/U_�w�{��7��w��n%�bX�w���n%�bX�1���蘉bX�����7Ĥ&B��$S2��S��8�Up�!2 �>�u��?!D�K����&�X�%�y�~Γq,K�����7�L��O��JsN�L�47LuE����X�'�{�Ɠq,KĿw�Γq,h�lO{��j	"w��Ғ	"}�f�ffP'��V(A�^�ޛ��%�b{�����bX�'9�zi7ı,O�}�&�X�%�{9�b�ْ��Ӧ�SUUp�!2!2v���,K��;�M&�X�%��ﱤ�Kı>�=�i7ı,Nx�{3i�y�ە\)��liMX��&�6�N��vRjD�[����u�����u5�����K��;�M&�X�%��ﱤ�Kı>�=�i7ı,O{�ޓq)	����m��:mӪ��U4\/�LK��w��nr�	��A�]��K�^�t��bX�'��}t��bX�'9�zi7򸩈�'����2ffJ�s09��_�	��'~Ɠq,K����]&�X�%��w^�Mı,K�=�cI��%�b}�
�*�Q4R��&�n�&Bg��?~׿]&�X�%���_��q,K��w��n%�bX��{��n%�bRf�(S"�T�i�*f�����L���;�M&�X�%��{�Ɠq,KĿs�Γq,K����]&�X�%�￿~<�{}���a�u;c�C���۫ɺ��3�����U����&���ᵹ����}ı,N����I��%�b_��gI��%�bw����KĤ,ݾ.�&Bd&B~�ѯ���UR���n�q,KĿw�Γp�8���%��~Γq,K�ｯ�I��%�bw����q?b�"X�����b�UN�4*�����	��	�����p� �,K��4��c�O� �ԑ`���E �a#��^��G��l�ND�����7ı,K���t��bX�{������#2�.8g��{��7����^�Mı,K�Ͻt��bX�%���t��bX�b'��߮�q,JBd,��l��UL�uJI&����	��K�Ͻt��bX�%���t��bX�'1��Mı,K��4��b]�7���{���+h�^����&�gn�rgSF�pY���r^.�aV�`���S��&1�q���Kı/�����Kı9�w��n%�bX��u��Kı;���I��%�b}�B��9�2*t�eT�U����L��Y=�7�~C���bw����Kı=���t��bX�%���t��bX�'��cǌ��6S8�s�&�X�%��w^�Mı,K��}t��bX�%���t��bX�'��}�&�X�%�}��Lg7H�&i�D���|Bd&H���/y�-ı,K��{:Mı,K�{�Ɠq,K�d���UjDAƢ�w�.�&Bd&B��t�5TUUSŘ�n�q,KĿs�Γq,K��ﱤ�Kı9���I��%�bnm�p�!2!2��g�J��UFC�.cۓ��"��Ńi�
6�L���q�^�<�$�.��E�����=�{��Y��ﱤ�Kı9���I��%�bw�צ�q,KĿs�Γq,K���w�]:�jGI̒9��_�	��9�zi7ı,N���n%�bX��{��n%�bX�c��4��bX�+��l��e˪RI54\/�L��L���4��bX�%���t��bX�'����&�X�%���^�Mı,K�{Γg)�i��7"p���ԏ��(�Ls߿gI��%�bs�~Ɠq,K��;�M&�X�����{��q,S!2w�_�U�T�Lʩ����	�bX�c��4��bX�'9�zi7ı,N����n%�bX��{��n%�bX�| ��	��Ÿ�.lŹ��U��=\`���ewg�R�6:�BE���N����;��t	��wU8��c�����Ԙ�B�%���ApV�g�Amc��N'k�����n�3��d�H�,�cnX�mgY�r��<֗.�Պ��y�q���ۛ]c���ӬH��U!Wk`XQ�qԒ�����%�B2 �Y.�.M-d��!���u�շ,4lfc= �5`�w�o-�Ĺř,��rf�����0�:ci��e�m���f;
�r�n��t��=���7���'y�zi7ı,N����n%�bX��{��n%�bX��{��n%�bY�>��~���X%o����7���'{�zi7ı,K�=��7ı,K����7ı,Ns���n%�bRO8檊���aӪ.�&Bd&%���t��bX�%���t��bX�'9�zi7ı,N����n%�bY	����4US*j���&Bd'��{:Mı,K��i7ı,N����n%�bX��{��n%�bRn�����*�t�ȥ�U����L�bs�צ�q,K��{�M&�X�%�~｝&�X�%�~���&�X�!�߯��E���	ڔۛn؄�vЛ4g8tq;qs �.�u��캟#Da0o6�1���.3��&�X�%���^�Mı,K��{:Mı,K��{:Mı,K��4��bX�'��`��ك���q1���3I��%�b_��gI�xD�:�C���O�X��{��n%�bX��u��Kı;����|Bd&Bd/g	�9*�R*t�eT�gI��%�b_��gI��%�bs���&�X�%��w^�Mı,K��z��&Bd&B�۔�ȧ�n��ә�Γq,K��;�Mı,K��4��bX�%���t��bX�%����������oq�����sY`,�M&�X�%��g��Mı,K��{:Mı,K���:Mı,K��i7ı,O�����ߦs����I�9�2����8�w�����c3��[��k$/9�ӻnV.\;���ո�?=�����{��%�~Γq,Kļ����n%�bX��}�A�'�1ı=�k��n%��	��߉�ꨪ)4T�U\/�N%�b_��gI��%�bs���&�X�%��w^�Mı,K��{:MĤ&Bd.�L��t�dt�ȥ�U���bX�';�l�n%�bX��{��K���j��U�G��3���|Ddp��_��RF@�;� Utg���'� O�@���U0E����Ҩ�A0b4�*>0�Cґ[ ��kB���iu��@�$�"��K��&BH�� 6'��4�	H�R�m� �@0?}P(�	��p"�@�
g�: !���]�	� �ȃ�@�����ﻼ�7ı,K����n%�d&B�sm1\�5P��U+��	���"{����Kı/=��t��bX�%���t��bX�';�l�n#!2!vwJs'�T˙&����;���bX�����n%�bX~c�~���>�bX�'}��4��bX�'y���>!2!2��ʐ�*IaSI�J�)�y�`�hIp4�k�.�[V�QG��Uw4�銝)�U5Up�!2!2�oU���%�bs���&�X�%��g��Mı,K��{:Mı,K��LL�t�n��ә����	��	��w�V���V8���'��~�Mı,K�߿gI��%�b_��gI��%�bO�p��i`�����7���{����I��%�b_��gI��%�b_��gI��%�bs���&�X�%����*�UH�2������L��W����n%�bX��w��n%�bX��}�I��%��=j�BP�@�U����5�]&�X�%�{;�bV�MME&������	��	���z�ı,K��i7ı,N���n%�bX�����n%�bX��}7�;=�4�#ɩ��]Yit�4+���I�e���h�Lv'[������w#gI��%�bs���&�X�%��w^�Mı,K��{:Mı,K�����&Bd&B�sm6�𩎪�˚�4��bX�'{���7ı,K�}��7ı,K����7ı,Nw�ڸ_�(�p���_�w�S2|�I&I�&s�c7I��%�b^{���7ı,K����7ı,Nw�٤�Kı7ky�/�L��L���w�52�R*t�pg�t��bX�%���t��bX�';�l�n%�bX��{��K�����;��_�	���u��2�2��nng�t��bX�';�l�n%�bX~���~Ɠ�%�b^{���7ı,K����7ı,M�D]�@ ��H ��b	b�����H�0@(�D���q�����Ms��Ų�q���ņb.�o �T�Gbchçz(_K��Z���h������uK�r�j�����T�c@$����˓;-Qd�\�:[�Y�	�Td�^D��9}�ɸ\��;k�	=����Ψ�S�D�l)dۇ9u�ڶ�4��d��� �ƒ��<��\���pg����5�LV{>.M��;=v�Yve���������|�;�Z��Mů//f�YcZ���Ʈ��;v���H���Ѡft�Xng4��c8��bX�'���Mı,K��{:Mı,K��{:�O�b%�bw���I��%�bw��/��L\gkss�i7ı,K�}��7ı,K����?*T�K���f�q,K��;���n%�bX��;��1$�QTRh����_�	��	����}ı,Nw�٤�K�C1��cI��%�b^{���7ı,O{��t�*�'2)sUp�!2!2n��&�X�%��s�Ɠq,KĿw�Γq,KĿ{�Γq,K��ޭ�jN�,uU\�R�_�	��g7��n%�bX�����n%�bX��w��n%�bX��}�I��%�bt������g�6��vX��mjw4t=�*�/fↃste󈧺s��xR컓3��Mı,K��{:Mı,K���:Mı,K��h?>���%��w�M����L��Y����ԪT�c3��:Mı,K���:M�Y;T�hE1F�6[��w;_��b%��͚Mı,K��}�&�X�%�~｝&�X�%��wX�&%��%�&2f��s��7ı,Nw�٤�Kı;�w��n%�bX�����n%�bX��w��n%�bX�ݾ��rMQ5ST�!3J�|Bd&~��V���n%�bX����:Mı,K���:Mı,K��i7ı,Nc�×�MU)çU7�!2!?oui7ı,?,q����'�,K���f�q,K��9�cI��%�b{�;�.�y�*�K�r1n�f�F�u�%�����́���'���Wj���u�&q��:Mı,K���:Mı,K��i7ı,N��4��bX�%���t��bX�'��{y�%ɜ�\��.3�&�X�%����4��bX�'q��Mı,K��{:Mı,FB~��_�	���ͻmI�����M&�X�%��s�Ɠq,KĿw�Γq,u� =����y�o:Mı,K��i7ı,O{���?&�Rɩ&i���_�	��	�{���Kı/�ﳤ�Kı9��f�q,K��9�cI��%�b}�Ms�n�)��'3C����	��	���{:Mı,K�,{�~��}ı,Oc���&�X�%��;�cI��%�g���߿^��Oe�
�yӸ(ۜ�����n�>q�����s-�L�Z�+Lh�)/938q1�fc9�s��%�bX���l�n%�bX��;�i7ı,O��{Mı	���z��&Bd&B}��]Pꉬ�9��Lc&�q,K��9�cI��%�b}����n%�bX��w��n%�bX��}�I��%�bs�x��91��Ü\�:Mı,K�w�Ɠq,KĿ{�Γq,K��{�Mı)	����\/�L��L���x*���2R\�9Ɠq,KĿ{�Γq,K��{�Mı,K���t��bX_��f���VQak
Te $*��h$ "���b�Q+!$��J���E��c��� ��� ���5����&�X�Bd/߿��IҪ��"�5W�!1,Nw�ޓq,KĽ�}�&�X�%��;�cI��%�b_��gI��%�d/С(��_��S>cNS���S�R�x��s���n��u�,G"�K�]��˲�s��	�常�s��%�bX�����7ı,O��{Mı,K���:�>���%��{����bX�'�޿���ʑ6MI2S����	��	��;�7�ı/�ﳤ�Kı9��zMı,K���t���LA$Nw��1��S(rL�+ P��ߪ� P��;��D����t��bX�'�ｍ=�����ow�����&� �qf����bX�';�oI��%�b^�Γq,KĿw�Γq,KĿ{�Ξ���{��7���}���hò�=ۉbX�%�;��7ı,K�}��7ı,K����7ı,Nw�ޓq,K��e����� /�I�'}(��X�R���m ˰&t��ԳV����	�%�4�[�L�5Ț�n/���1�H!ywkh��"q�s����r�*��d�g���d��vsY����U'i�N:g��lq��;�n�\ٝK�ԖY�vyẹ���.�������y�rw:Lv�[����/mgу��6Z�J�4���h�j���e�l�.U�qud{X[��:.���N�;6���4�&\[�n��dưr�V�$덵l���<�(��8���礫��%�bX�ǻ�i7ı,K����7ı,Nw�٤�Kı/y�gI�!2!<3_1�USC�I��UM��Kı/�ﳤ�Kı9��f�q,KĽ�}�&�X�%��;�cI�	��	��{E�N��U#��IsUp�ı,Nw�٤�Kı/y�gI��%�b}����n%�bX��w��|Bd&Bd/w>���EPJ*�9sUJ��K��1�gI��%�bs��Mı,K���:Mı,K��i7ı,O{��+����c8����s��Kı>�}�i7ı,K����7ı,Nw�٤�Kı/sz��&Bd&B��s?LӖ:��UJeinɕ��g�s�al�ō�T	�{Y����a�,gunK��?=ߛ�oq���_��gI��%�bs���&�X�%�{��:Mı,K�w�Ɠq,K��ۗ0J'�2M:�����	��	����f�p��m�j&�X��ﳤ�Kı9�{��n%�bX�c��4���oq�����Ե03F�����ı,K����n%�bX�c��4��bX�'�ｍ&�X�%����4��d&Bd'�kd9:����Ī�UW�?C119�~��&�X�%����Mı,K��i7ı,K����|Bd&Bd'��ܪ��Ҥ�곜i7ı,O{=��n%�bX��}�I��%�b_{�Γq,K������Kı? =��ɏ�I�L��;xx˧�m���ml����;y�5��!�;����Squ!v^�?=���7���'}��4��bX�%����7ı,O��{Mı,K��}t��bX�B�s�RO�%T�����|Bd&Bq/��gI���bX�c��4��bX�'q��Mı,K��4��bX����(q?�5$�N���&Bd+�w�Ɠq,K��9�cI��3�äD��DmO\@��� ��C�ͫ��7��_��q,K��{��I��%�bw���n1�b��&rK���Mı,��,D�{���n%�bX����i7ı,O��zi7ı,O��{Mı,K�����"h�&���MM����L��Y�|\-ı,K�~��M'�,K��=��4��bX�'q��Mı,K���ϗ���=�����݃e�v�v�M3Ѻ�v��=f��=�V=���aՆk�س4��bX�'��4��bX�'�ｍ&�X�%��s�Ƈq,K��{�.�&Bd&By�l�&ꂪ��L���n%�bX�c��4���Uc���b{��i7ı,N���4��bX�'��4��� 1S,K��_�c��ܙ).3��I��%�b{��i7ı,Nw���n%�bX�{���n%�bX�c��4��bX�'���f��RM'3N���|Bd&Bd,ݾ.�%�b}���I��%�b}����n%�`a ]�.n��du��}���	��	����d!�C*�9sSF�q,K���צ�q,K������Kı/9�gI��%�bs�צ�q,K��x�צ.e�L�g2\�.���X癈y�
��g�k�fe-z��9[s��Ŭ��fr�m�������ow�ｍ&�X�%�~�}�&�X�%���^�Mı,K��^�Mı,K����sR�4�EUM����L��O����n%�bX��u��Kı>�u��Kı>�}�i7ı,N�sm�MI��*��\/�L��L���^�Mı,K��^�Mı��D�Nc߿cI��%�b^{߳��K�L��_t��Ujf��Qp�!2���צ�q,K������Kı/�ﳤ�K��9���I��%�b^z�0x�9��3��%�ɤ�Kı>�}�i7ı,K����n%�bX��u��Kı=�{f�q,K�����,���L��7���H�$���P�	 g�&9\#$R$�HL@a�$!��`�#!�/a�'��Sf��xB���H��$�H@ ���b�7���L��ph!y��,a%w�e�����'d)bb%����&~��t�L�ń�"�B	$I"B-U�p1H�, I�4�f��)�D��RF,!�@�@�:���A�҆	1���� �A��\@ʤi��s$�,a��ia�� )Á�*HgT�d �@䈴0�-XL!ܵ�sD�� 0�NobbH�7Fy��sm$[%�4�D�������%�S�Rpkl�*�E�[N�m:��&J�rb�m  u�H��](Fu�vŽ��vE���;MT��5I-7'Kv5��4������I��.T��G���&ҵ�ۦ�F��9.`�mۨ<5x;q+�$6CC1�<���䭃jۥ�GPe�hw�I[c��s���7��{�]&�����1�a�@�3۰�Tְ�Y�=�@�9�쭻kl�r �u����ѝW������у
��Υ��g@�ێFɵ�t�v��2Ja㐫k;�.j��yl*�a�U*�Sj���mֈ���@U��Uj����v�U�Y<��.����m������Z�k�R���	��]��[v�*��Y"B��M)m�����W[u- R���I�� �͚V�嵢����Z�������S,���)k4S�e急^�5j�)�j��v�P�밽aJ���l�6 ��v�cg`�r��WU����6ݖ�r��M�"��6�M`.���Q�����W�������㞇h`�/�NTl,z�imں�p�s��C�0���\�f�'ۣ�N]��h]�m�v:����g���"����B�ɠ�+����ζ'�ї ] 6��Z�^��]�mp;`�T�W,'mX!�Ŋ#G.6���nۋ�]v��TM,ں�w�v^��á;<��s�Z�i�,�Z 3�0H�Ρ�8A*�R2,m�4��n@ȱ�1̉����S�	�u�P�m�,�F���W����q���vkI���a�棃����3ý�O8F��]��K��6R�(@�[e��%�
d��e@۵WUTjV��c��f�u��Mc:�]��S"=�L,�vu�u�َ�*�F{�n�gSxl�Z��wI̡UF��Q��.�(k��
�UU�8edq�̉R{=��a�U�s�/V��r�7p[VY킁Q�v�&�S$��gYyw,vJ��w{��d� �6�SSh�' v��
Aj��JP�`�qS�@�"}Cx~��7�[�˚;J��T�l�
�%�'��.xt�t:�V��n�\�Q�T.0��+��lm���Qʑ�ɛ���ٰ��Q8�UR�l
iH��[03��lF�&�4t��g�ޚ�js����Wf�S��[�a�UIz�5�[���^���y]��*�s�6�n\fp��9t䩣�"�����a���:�s�ݤ�O3 &6Ĵ�S�����St������� �nj�8a;���wf�Nsѵv���l2l���;O�w���oq�_{�Γq,K��{�M&�X�%��{�4�},K�����n%�c��}~���Ui������{��7���4��bX�'��l�n%�bX�c��4��bX�%�{��7ıL���� �%�mT�����|Bd&%��{�4��bX�'�ｍ&�X�R������:Mı,K���M&�R!2g5ɯ�H�$��eӪW��g������i7ı,K����&�X�%���^�Mı,���j�&Bd&B����R ��4�EUM��X�%�}��:Mı,K��4��bX�'��l�n%�bX�c��4��bX�'���_a��-�c8��.JZS��!���y9���gi����u]��v6'ʠrM9EMWмBd&Bd-��I��%�b}���I��%�b}����~Q�D�K��;���n%�bY�?�O��9�r�-�����7���'��4��������O�X�ǹ�i7ı,O���Mı,K��i_�	��	浼Rm�SSQI�T\�bX�'�ｍ&�X�%��s�Ɠq,K��{�Mı,K�w^�W�&Bd&Bxf���Jr�Ҥ�檦�q,K��9�cI��%�bs���&�X�%��=�M&�X�%��;�c^���7���{�����n*~&�X�%����4��bX���;����%�bs��Mı,K���_�	�������G���2PS��ׂ���I�\����R��x}\]���[O�n'),X�p�]���oq����;�_��q,K������Kı9�w��~R},K���Mı,��]�����L���R�j��p�!2�b}����n%�bX��;�i7ı,Nw�٤�Kı>���K��w{�sN�J*DM!�USp�!2�bsﱤ�Kı9��f�q,v��B�@��C�X'�f'�;�k�I��%�b{����KĲ��'Πs.�MMMM����L�;�~��n%�bX���~�Mı,K�w�Ɠq,K��9�cI��)��	�����S
�3Cti\/�LK���צ�q,K������Kı9�w��n%�bX��}�I��{��7����?~�l<��QKl���r���=�͓����p�����;��brZ��Y�8�2丹��n%�bX�c��4��HL����`f�q�/�{:��3zT�&�R�Ҕ9���<��7��fn�s�Łś����Ҝ�q�۔��n��� =�`���1��b�-n���RJM8�`s�4�8�u�~͛�FB��Iz����71��v6)ȓr7�ś����k�;�4�9׺�R�N��9)S��(:"x�WY�:�6K6�x�1.�ݙ�V����0��0)(R�#�:����M,u��7]�����F�M����`s{����Ɉ�ss.�ĉ)�%HX]�vn�<�,�;7g� �k��ʎ
9'ҔR;����s��߫�U�}>� ��7C�QE)М������M,-�vn�*�:�h�QA�HN�ڶ̴����D�a����Y�x�{�݋�l�7�q��v�a�°��/��
��U5\'b[k���:9���XE�`<��8 ���u�5>\ƒ���u�i�"4�n����	c�#C&�-�髇n�t�
���jitn3���#��@ݨ� �p�g�iR6筺��[Aīmp�๶h��ի�[gɞ�&]�vս�w������|�����V5犸�Z��c�J�����6����][�1Dm�
qʑ�۔��H�nO.9�[���@wIy���fm��yy�����Ɉ|� 9�������/	�M��9n%#�:��h|� 9����n*/n��!M9Bd������M,-�vn�����F�M�j�#�;�4@z㘀��1 ���U_�����pW-\a��
��+��F{s�Bz����b���8��$�عlŧ��}�[�|� 9�� �mFTp�����qXY��R���U ,H� cS7\�5$�9��Hs�4���lt�5�BrG`uw6lfm�:?�L���Ł��~�_�H��Ɠ��RG`w3n�nM,,�v.���M���6��NIV�� >�����%�� 9����L�[>\�e˜��mN7�C�������D;<�ۜS=՜����2�������_9�n*@{�� ۊ�d@8SnRL�;�����Fn����zx�8�u����q�ڢ����fڰ>ܭ,�u�" P��8$��	�(|S
���M�:�5�洵� �)�%8�9(���|X{�6��f��fڰ�ݍ��_:C��8�u����n*@z=�<.`L,��,�t��ぺkm�ny�v��ۑ�tv��e�j������{�|�+�mtE�a���~��� 9����[��B�o+`�Rn)#�;��W��Sfy��w_���⟒;���.?�`I)4�`w���@y䖀�c�����p�J|&�Ir'˻=�`w�X��V�(�\DVU^�{6�jh�Y��w�{���c�����������j㎆�	�A������w(��:����.c���"c��u#G,��e�;�
8�mAH��߮�w&�n���}��A�{�`y旛R���i��[�x�9�� t�n������B����`sj�;��V3&�ӹ�Ӥ�ࣔ�Y�����-��H�A����؀՛��"t��E`w3n��&�n��{�������Ɠ�"���eZ�O�Q�v[�e�l��9A&�9y��7����<��B3������XX6�������f��g� +�٫iKa���`�*��7l]v�Ň�k[��J���^�[����}Y�(�V�uC��_Fֺ�f;��#����x)I_X	@-!�2�<#)&�5ņx����4rqk��.�<!\-]�Ḫ
��{���������.���h�/q;��s��Xۭ=Oa�L�r,Ma5���jM�өѰ$��rJ��<Xy�6ޝ��������֬�ߙ(wP4�ȓn'�7]�ν�`w3n�{+K�
�����P� �)7EUM���`ffڳ��3����1���l�B
��n8�PR+36���ri`qn�9׺�FkK[R4�MD�e�����& =�%�qR�w�NC��<�R���m�$�;�n�阣��[I��v����pWob��r�U�i���sm�b�Ih�T��Z ��Z��uj9R������yϾ��]�
!o�)E�=�`{'y�=ݛ����8D�$���ͺ�:�����1�����yKs��e����R����w��`c����y�6fmՁ��C�\�b�"M�8���V[s���Z��y�0�/oc�+k��BΧ�H�v��y%sm�؃v0�r�k�R}�p��M�9�pP���w'؀��H<�������)l�q��N;s6���=�`o^h���w�H�o��������*)�`{g������zS���v��u8Y��D�@����9� ��
X��2i��s�ʁ ��JJ�"�d�XF$!1YH�ls��&(X�$H;0�\A��a"F0�R�$�#1Č!!��!�S$L��ˉ!!h 6���T�qG*��H�N#��Uu�A�����@0=^*߄QU���ˍ��w��I7z[Ŭt䦜LT��7�4VVf�s6ՇC��s�3�]*Z�uR�Rni��& qR�Ih\p��mFl��S
`�t�6�*H�n�'�^{��ۛ�I�\�����͖s1qw����T��Z�3���+�%���`g���vG��Rm�*��=��=Ӽ;�M���j��f��w@���&��V5�����g�Ks}u`f�yX�������H�<ݛ=�����a�D)IA
YR#����vf�8��˧S2麩�3�ZX�3k���{�`y�����O>^߽����Ьj�1¤�*e��ۦkM�3��\6G����7�*q�e3kot�g�Z�-���o`��j���t��j�$V5��U&�{�6�k��;��(�Ìэu24�%JR%`b�y���,�W�_RY��Vc��`qw+G
p��)I^n� :=��Ih�e��Ɉf�N�'ю���NIVq�������M���j���A��4L�ߡ��Zڦy�:�2�������nn:�l�v^�{^���dBT��$m�yƹ�!$Sb0h���fl
t�f�f�]�BΞ��R�
]j�Y{[�݆�(��ův�wq��6��#vݨ#�7�Y�v{g��\ڹ�g^q�3ۮb6b�ݶ�m[��^\���
�ͬ�u�==&ٶv��̶��+�c��U3pfb��s�����D?�O좇�����p��bu��63�u>Z�{���vp��کY�]Y�[8Yqfw8�m�Š{�?%`uf�;�4�;�uX�������I%+�7]�ۊ��K@zd�h�݅m^K/#M6�R;36���=�`srjVVn� �֩	�ND�B��_|�k��ޮ�`y����,�hOhR9"�I��٭XY���M,��V�)|��$D����8��,�F77I�QȻ�'=�SN�����<=���Q�*P��+�7]��ɥ�ܝ��
>P�wW7`y殗M9��U�-��s�I9�3٭|����u2�ID%)D*����v��7`y���n�N�r����܎q���e��x��lͮ,�l���F����Ӱ�
!~�Js�}�]���~�=�K��U�n��)��9D$��nL@>{<���e�ߣ��~��T�����N�/�#s)�-�I&n��ܗp��m����(���DmD�|sg���U��٩XY��sZ�'�Hm9�G*��=���!&�oWK�1�t���W�
!��Z+]z�)��S$���?z;�7]�N��R!$"FH ��u8������1�hԓ��w�NO�޶�IJP���l:"�ޫ��Ձ�s]���c�8����D��
RNfn�$qR�s2M� 㚀������ă�B�z�gd��R�эlc��\��J��`�MX�u>E���3\��MYy��Hq�@t�7�jG��9��.|4�ȓm'��{�ߪ�(M���X�\X���6�ĩDԠNQM��n{���ɥ��y������ �Mji��m��}�|XӼ�l���?/��@U
�k��Ԓs���b��g77o6��DLr�2M� 㚀��,*:�G��5*$�1�� ����	���gtY�<���{+��U����GL�+��c���`ovi`f��`w�Z"n2S��r; �sP�� �9h2M���L�ʷ)�)'�������y��UUU|�������v;�[�*I������N�=��S`y���r��g_�|�X�)
��6��3^�v(����ή,d��oEBJR��"�	}��I�j��Ze����<��d�=z����f��d��n���(���y҈�.�X��c�$��18�D�TZ�:�Y���u.��Z��'�Zl<��c���%�-��7f���m��{bv9�7�pb� Yݧ���c��)�#׎�ʶƬ�60��U�t3�uP�ݺ��P#S$��[\��T���tk�����v6m�Qd���SBJ����UnSV�MS
U![0s���ۉf٘�Ƈ6-v�Xli�nz���iv�⨤caQ�SnG�yw��`ovi`w�����G`{t�t�4�cs4�T��/�P��6{���=�6Vn� �-m���TiȜ�9Vq��&�����T�o.��n�I$NT$���{���uX��Vu� �߱h ���E8�vy%�'H����&�<.]���X��玚9�`m�ง������>ֶ�qv�Ӽ�OH�i�pMBG :c���n =nL@{���(�G ��rJ�:�5�R�+��Т�vojl?ń��j�ICgf���q�M�6ґ���7`qf�7ri`ufk���) ĘT�&7�8�u��4�:�5�z�����v�P�*�7i����۫��d��_I��~���n^��WM��-�NI���s���v�˷G7�Xۥ8�rD�B^^[��a��x�}h�L����^��mh�*�dNI#RSJB��x��3�#���`�8���Xm�ٕ�a�S6�۳`g���Ram(�������[Y���ν��]��Q�Q�J����@>{s� <�L�����թ�u�A�)����ɥ�Д$���3�{�6{+K<�I�3�p�G#�{O6��kg�uk\aOc�/nY��nb�J{��v���+��6<�L��Ɉ�`��Z�KE��aQ�I���,�vw&�rs]��N���D$�;5�)7<ʗR�n%#�76x�9�5XǺ݁ř��;�[��������HXǚ��n��>y�6
B���}��X���#�F�I):dqXY���ř1 ��x�$��f����R����t��9ؒt�3�LՇÛ.�˦�WS�[�6�R�QD���,�vw+K���B_0ܞ�j�e�TQ)BN8��M/�׾V����8�5��N��8�%&�p�9��d��[s����wN��ȓm)��{��Y���M,,�v7vܕ!Bl�%r;����@zۘ�}�n =^�~���d�%̤$V�0#
�V4cu��df~ i/XD�� �P�gf
�@��-*d��+�"�9HL���cZق�-#)la"1�b�	kj���l��Ķ�B֔�.�avL#�dCQ��VŤ]+jD���!X�qLHHD�I0$##0J���,H@���8@�	����[��6�r(8� �D$&���$)e��~��%���&a�N�����6��lwnn]j�;pč���7]����]���A�(6�  96�n�n�ER�)���p皝l$A��vzj��G�ȱ�;EֶI��Uv:�&v��ɤ��VW��B���0�-����ȼn���K��O:9���5�z�E�n�^����m82��������rkծ@ysa�[��mw���:�к��f�s�n֑�[j��3���C`cS� Z�ax��ZtR�T��N˻8ʣE[O%\�l�ڐ����'\���6��KUH�u��pl�R�h�iU�Dr^��j���z��ĵ����"ҭ;��~_*����ԜK��eK��ݵ� �3b�z�d��[���]��%� ���᝕>]�h>�- 
\�� *���R��3���*�k��l�(�2�se�n��v� G��Y��%�:��L��k [T� z�y�y�J����ZA�l�#�s8����)��0\j��s��.;n��F3pgtb��t���v�Ƞ����y�GnwF�-��y��K���sۣ7@�GN_Nyܜ§6�c�a0����ɬ���\^��o<�7n8�I�"9�:Tګ�����j��K���	�0�V͓K�y��j�y��4��H�&)Ij�W|�>�r7NT-�[;�]l�6�C��1@����\\��/tm�k>=�'��\�r��ju5�f���)"ޜ5� � ��1����b�x�v�vS7(RX�\��M��[N�X�9��?	^��n��s��C]jCa	t\�ȸ��N�H�٤�3�Fθ��s�-��N�I[�c�؈��Vj�I��	)��[%&���[�cEUORˇlY�t����
���� pӵp�1ݎ�4��eKzv˺N��j�R� �ش�D��@R�@umUV��ގsu�Ӳ`�\Qu�\�R���a���K��ʔ��Rm*�]^r��f������~�w���i0m6 <0(�<�� ~���U �˴�^	�kr��rg��<V���[�E��jC�[-��Z�d���m�>ݪ��:З:"xīV�I��ev,����Π[h��Ϋv1�tKqU��s���i��m�n*k�Q�cu��ebU�w]nb�m��]��ώ�q����%97�(�s���V�t����9���[uͮ.n���v�6����U UA]�]I'R�/A%��$oI�u�9	R�������V��B�Td����U��|�po�U����1Վ`�%ڻ\�-Ѻrch�p���3�����@zۘ�}�n =m�@�f`��pNG$,,�vu��`qfl��/�BP��twQS35*��9R^耏>�q�nb�� <���>�[BDN(��r;�3]��ɥ�����ν��]�և���Jq�`gri`{���n?z;�����~w�����g%Aꃣ� *�!��6���1�!�gi�'sճ����n������&���b�X��j�1S�&�Nu�Ǯ�����0��@�
aG�_*��]���,����I���n9I6Rp6�vVo���ɥ�����ν�����ƙ"m�n�l9B�Oo}��7z��sT�~P��^{��3W���)	%7#�z�\r���1 ���L��߮���5[qTWl%�FD{N�X�WY���n۰��)�Fe�y�/![��!�_I��a�~�_�`�߄��$z��n&����.��U}�l�����������7ɳ^j�e���R�����<X̚Yꮟ}Kc�D]���l~ޛ�5뛩��u!����h���-뒦 =m�@6��5���*r$�����Ѡ=m�@>{�9hre������%���1�^��{(]Q�k��9�v������^��,<��z�(�����1#��x�%�@NwwEJI�M��I�`n��Xǚ�[�;�3]�w����IH���G% <��@K����1#���V��"��t��5n��,�vI��5&v�r �rE��ι�`j�m$�I�Ҕ7`qfk�$qR���!�	)ٵ+h�ܥ�v�p������<H�n�T�y�koP����K��`�:�%%%)$���ͺ�8��@K����1�K��s�ỀꔷUJ��'5�D6s��l=ޛw6����hv9m�E`j��l�f͜�(o�zՁ�����ݹ��T�e6JCi��Y���۫��KV���MT�	�`�m6�Oq#���@K�V =|� >����{��q��N¬d*��WS��+9leH��:�7�k'^f���&/�̌�vG���G9�)��H�=�=��M1mn�i�.n#������M�<ɑ��6������&x�p�uٜݛ;��)���Xl2��r�r&z��>r����uYc:2p�&��#t=Xݮq��<���y��c�V���Tb�F�Ìb�Q,M��~����~{�w��ϗo�zNe���팯b5�R���G2�W�7ϟ���ޖ��*��T�\QBr���l��ͧ`qw5���Vϩu��y�nJjD�JB������&�<ޛs�Ձ����J!�^p�Ԣ�J6��q�N����3sn�u��Ӱ1w+ZI��)I)SN��͵`}��v=�SaТ'���3/7r?�������`s�5X� =|� qR�ʙuyܢu��ٶ� u<��o.x�M8�s��]>������V֘��7gq���ͷ��������*@zۘ�rE�����e6JCi��ǚ�U}��76����k�1n��t�JRn��Cn'U6nm���g(I&��q6�w��;���)�M287 ���U��Hb���*@z�f�f�t����*i��t��DD{ky������<�`gu|)��)�N�ʅ�P���a�)��/c���5�\�[�����Nxv,T�7*&�%���ǚ��۫��U��wG`uw+[j4�F����m ㊐x��@y㖀�5m�#�G9)�IV;�K��Ȇ�-U�E�la"%$@�"���ٰ7۶����t2�9m��`bݭvs]���já�6��3���t�2'%&N^V���b� =�`�뒦 ����/���B�û����C1ٍKsv���4룴k[N��{�8x^Հ�s4��@7"���rTϿUW�9��r��N)�jJ�9ܚ_BQ���M���`fnڰ>f�mTn��C��Ґ�9׻J��^j�;�۫�ɥ���*ߣr�	Ҕ
I)XtBO�[���޵`}�,9,8�_(���O�}�z�u$����13��Q1JIH�;�۫�ɥ��ɱX��V-ƛ�(�&�Pm�I$��#=5Ga.���\:�ƕl�9"�<{M<�5�L��?�q����`s2i`grlV1��ͺ�73X$ՠb��dp�=�h<r��T��{�W�}�+mDƛ)�R	$����;��V3&�{�b�;��H�t��(3Kݴ7 =�`��{6�}��ꪥכ�`�?6�"JR	�9*��r��:=��?����=���W����׽��|���v�vJ��
�PX:��e����xv�7iК�<^ƻTƮQ�R7HI�!�[�7a���vԘ��l6�{d��e��Z�X6ݶ�k�ۢX9Ӹ���7l[;�\��[Z�h3�\�F}v���E<�V��hΪ�,v!#%u�kE��?خ~Q5�"�`�t���yƕ�'V`��,�X^n�gFHB�d�ք�Rv9⸑99�t��ؖ����Ues�q]rH��NP���cR��N�獏\Ok����6˫/9yř��V.[i��]p�m1)z�°8����mՁ�������ܩCb�
G`qw& 9���"��8Z��&a�曚^���������*@yㅠ1fk�7��n�t�r����`sdT���@;nb�����2��8D�jJ�9�4V,�vs6Ձ��i`R���*Yҥ�MMS
��v]�Ժ��f"��n���t�J;N�#�y;����c�D�)2R$���pw�u`s��
��R#-bJ�3ns�I>�;�_(�qDv�oZ����`f<�X�5�潒GI�QH,�3v��`���@;nb���[���J�)LjB��<�X�6lfm�����+w9MT�*�(�
�ř���}���p�}u`s�4V�$����Dq�C";��Zz�y6�iyn-���m<b훧x&6!���
E���;�ͺ�9��V:�E︃Vo���<���>��B�����qRݎ�w�b��H	�0N�؅N4�r�u�����s���a�w?&\�
� �E$XEd �1$S;�f>�~��FD� 0�R�����bG��Dt�AddH� @I&jԈ���LF�Ĉ�$�@"	�B"��C� �G���)	 0)�:�s��>AF���
tQl�v�n�3Y��"@��-i ����X�~��@�B�hÊ�ʡ�F*T�@�>S�s�k "�~C8�.#J�H�w�.!TGz�ɐ�j/�C uH�}�Pp�ZD'	Y��%��9��.����L�z��R�r1�kBG	����*p�#eDz
";v�b��qL�riHd��)�DY�C��v��H ��G����RM��X�ԭ�6�E6JD�AXך�{6Ձ��ڰ�~�������)SՖ^�fi{���qR��Hv8Z:�U���n�6D��D�O�IB�䝬v,�AZ��l<a��kv�>\�W9"t��R����NF����u`s�4Vc�}�|�3zՁ��*��J��\�y���c���-��HI :���*7*4���X�5X̊��*@yㅠ=m��(���0����ʹ7 =T���A�U����0A� ��w�+�1y[�} ���$���u`yㅠ�-��H�~�*|fVa귔��ϺkZl;���͡�8�.mO.b����8oV{��{1xU��E+�6�����vd�ٛk�a��`ow2ꜱ�RL��UUC�3'5�DB�����V��Ձ�Nh�l��i�JT�%:	���m ��R�EH<p�x��od��1E ����<��{�`vd��y%�9��� L����ۼ���ͤ�8Z�$�7 9����%
҄�J!<��ٙ)�4:�j݀��g�Ķ�+g��(6]���餈��A�Μ���͸$c9m��ڌ�����Sn�ME�jH9Cv]����4��.��8\lqvDq���ftx�;�7;����8꼺,u�b�iv�U(l��)Mk���J��xp:^����$ȵA�mm�V�L��y��L�|�����]R����6�6�έ�@g{g�,�k�
R���w~ww���X����c\(V��ҳ���^�v랆uy��|�x&�	R�ܨ4Ӕ
G�3��Vs6���d����׾��4�e7!e�]���9����<p�����U�G���$�(�Q�c�U�������@{�K@sqR92��)mԕN'��E`s�uX�۫�ɥ�����S@��$�V�$�7 ;������V?(�6���A�)�{�wϝ��P��������r��{N�	`��.y�{H%�v���H�@yㅠ=�%��m�1E �����&��WO��>�,:��
oszƷ.��s�ԓ�f�X[���7R�NG��9�4����7 ;��-�ɠn�闗�A{���=}& 9����c����j��1	�I���qR�� =m��& ?��~�1��U̇"2�Y]�G��r9��GE�ݓuG4����\���9��W��M�m��M�@zۆ =nL@sqR<�E'j�ۨ�&�Nf����� 9������˽�̠�6�*�����ٰ=����J�8��GD(J%
����i`c��l�ց��uI�)��ͺ�;ך�,�����`��{$$b�A9%X��>���d��:��b����s�o�l�ڃ�e��\��.۪Ѯ��Zu�/Ot�l4pJ.ť�H3.Ţ��1�rb�����@Kx̀F�i�ヰ8�u��۫��U�ř��{^���#d�)J�7wO� :ۘ���@zܘ�ޚ�\�}���!�*��<�`qg;1�&�;�jN �`�� S�]s8�Ձ��t6�ۨ�&�R;�3G`w�{��3w�X~͛�(�=���Oػt�ո,k�rv��c����7Oh�:��զ�)ԁAm�n]�r�ug���mՁ���視��wð;�����J���)��ͺ�<��6�3I�>���Q
"a��2�7���A9%X�|�,���.��������:�Ah䔜rF�3m�}�|b��� 9��ݎZVf��$����N8;�����fڰ=�,�f�`��0i'pi���*��xs�	��)R�[ڤ����ϧ�:V�82�����(ɼ@�<�<%n����*���r͝�EP�`�,������,�i:A��ީ�:N������My��t�᮷e�6��ݧ�PQǳ�$��צ���b l��l<����v5[8���&�-YJ\�hv��.@mR:���Y�n{v�sk��ɡ�9�Cحų������������s��ߟ�\�<�m��d�x�>���<[&���5�n�(G8��h�ީn��K���ݶo�H�@zۆ*ݒ+��U��������U��ɥ��n���1��H	$���^fV旙��[p��Ihn*@sɥ���=Q��e6D2G �cݴ7 ;���n��WV^ѐ2���/v��T��{v9���Ӻ��-�2)g&��"*����ӷc+�֞����k��g������W�V�\*�t�J��A9%t�����^lvw_����Ձ��W�T�rF�SN������
!�
�"*Js�6s6���d��ՙ�&5#�m)@�zZ���7 9���-͉2$�diJI9#�;��Vs&�1�����`suj��5(W��Ho`��{.��& 9�������?gi4��}D�5�/J�n�	B����>D�][�kn\�H�����zmy�nh��=�h<���T����(�FP�)S��܍XǺ�n*@s{���@{�����^@ډ��)��ͺ�;�4�>ϝ<rkVn� ���45�	�p��`wc���=�h_I����됲�cT�b���V;�Z�8�����V�9����9���nSum�l�X,��m�g��`��/W�d�RqN/t�T�7jI �(�k�ug����,����E`n�ؓ"MFF����; �f��Fc�+��°8���n�V�E �R�'$�;ך�x�h_I����rK��lun7���֬.� �se�X�D8��T$�x~���ٮ��_��8��Ձś��;��`wk�>̭�`~IB�ۙ����s-���%�=��h�3����nCA�;:�2T�4�N����6ڦ�Ɯ����q�3},��V3&�� ��y����$8F�:�5߾�#���X[�; �se�պ!'���JE"q�̚��rb��H�s#���f��f�Y��h_I�� :��@skv�͉��p�1JrG`w����3/y�{�4�9���(Q
W��(����EW�"(��DUȊ"��Q_���*��AQ��ݫP�B0	TIEA	P�@T$ dE@AdEBAaP�	 dD� ��DU�U�(���EV��*�((���DUȊ"��Q_򂈪�ADU�EW�EW��PVI��{:(���` �����\��T���)%�p��PS= 0  � (  E�4�� >�@��*��R $�T�    �)@ P� �P*HBD��EJRQU
D��*�8    �h 
��� �O��v6���^,�k��l�ݵ.m�s=��D�` ,������� ��j{9=U�x��}�1��b��z�����wS���G:�e�=���y�ϱ���U��J  P
  P�@�oB�k���{�����u��R� ���>�T��]r::}�HLL*�{��� �ϯU�M� z���{��ɯ^��wmW���� ��}���R�ws���*�ܚ����   ( (�� ӥ��J��+�;5sgW�w�t�� 4�����۶�[��kť�\��p}���K6�3��o �x�綽�9}|����K��yu��9��{y���< ���s�X����ռ�ͽ5�  x   �  �n������C9�u��ԥ�R�� ���)fJS}gE��R���R��Ҕ��r�R�M(�)K,�(� iJ0 )JR�(�)e��)e����R�X�nR���iJQ�()F&����h� � �@
 PP; �)J[����i@,f���l��׀>�=y\��W6_>μ�]��,�X �i{n���[޽��   �W�G{w�z�\} �R�}�\��Nc^�o��K��9�+�gT�1�x��� z�꧶��P  "��2����   ���R�F   ��R��MR&  4��D�R�  �A1JSH���'�������q���|bN��=���� �*����QUʈ����QU�dEW��*�PUO���C�B$ �	 H@! �XƄjBO���w��P�6���B��JS0�
�B��"P�H�P��k8���c)�\P�R���q��3�1)#"D�g���($J�
��;,d�T7�)z�[h��4��S��l��ˬ�˩y,f�u�MHF�S���#{F��F朋z'��޾��h#��}��8D��6A�0�1 @�7{ۢ$H$�4�s2lA��(n 6�9���i�]Q�ES>�4�D�V�n�ɽ$ք"�H\"P�2�7�Dț`T1�����mMP[��zr�@E�A]�"�������z�iZA�u����*�}��G;57�[��Cb't��}��wL�ַ��Mf+a$L&F%��I&	��2�?P�!B[M\��Ǡ��N� �HK��6gp�^�.��`%YLo[/oN���ǝޗ��[�dx��22Yo{\w5.���s3�bb�ZB�Z� m|}�̍��k	^�bi���{6�Bn�����P�BDR���2��G`��a�S�+ 2��L�o��0�j��;�}N��ӯ^���vkzf��w2w��x��	��\?_�77�oW��E�:��+�x��t>\g{1�V	q�%�������F+��"q�����{Ӓ�9(�	$�����bo\��wDW�I�r`>>�ɺ���BF� �E+ g0�)nͦ[r�ѴI����ͺ�������ڨ�s[!kU՘hZ��B˜�s�)�S�!pJFcfˌ�aLI��9v�M�O�|F�z�	��!�3@餞� ����.���.2j�B%%�#:}�O�|�����etg[˭�(aƱ%��%i��i�D�Hcސ���ˡ4wss�<���}��o����7&��4����#-ʋ5���U�*2��Z�Ŧ4n\i�3btΡ!�Ƃ��	a54@�!�4eR?P� �ؑ J"51�)Bb�(�%%ƈ\0�
2���%#F`�pԙ	:�q��1�X5bV$���C�9�z��L��|���F�1�
ˮ�}hF_l"g!�fl��L�F�81i�l����5���6/P�8$
a��4h4� CC�V���e$��"�x�L��μ���+Jضl#y��y�:�B�H�f;ۇ"l�M��H�-�&5��
� #�Z0b�0! 3.s!�gY�T�'H�*B��d$L͆&3��:��6��WF���$a�_r���ᐍ0*`��8|��_�q�>�6�I��U���Uf�4�"/���(3@�)�ٱ͠z�_/�)�7�5E���3�߭�>����T�0p����gx��Z������i�HCLơ����>���$ ��A.�C�}Μ����М�}�f�z���m���t��3(�Mu��eÂC�,���M�b1��`AH�$a4�g4D1Lj���_o�N�A���:�u��'�L��,6�@��	
5(��!3k��W�P\�P4�C�����x��%�h�)�h�0,�!�c$��Y�c1,i
n���\���m+$ҹ{��c���b�:���}g�QUE�}�E�O~�}��M��b�ŧ���uFU=�]{j�ǳ�����H��a�����lP�0f�\71�!XS&��gA
��R��I����������A�!q�t�1~���ݜާ]��CZ�K��<6��-"��pR�}�����#O����3���d#�$��b�a�BW8.kb2&]M3Fos����t��&V���ZUЛ����<��.}P����C�HCY�!��SZ�l��.�'>�dvZ��рaF0%�9�w:�8:k�����<�|�i����UV�Y ��5Yq|��΍�9������j8H-cR+"0C�Ɣ� �:�Ƅn2B�%B	~�,��*u#pJd�ġ������H�K)�]3;ր�@ߍ���s�8}u�H��Łe����w�!0B�l�(JĤF$J�ZB�tfI�'x($F�� ����t0i�#X��)$Q��h��%�v$5����š=]������'���\�I ���'�1=[���ki��X���II	vr�X��s#\5U4��S�hm�Ms�B�[ͮ�>ಾW{�� �Z֢wq�]�]�YVk�w�F��Q�
e	�k��%�s7��|k�@�a�|�ý�уﴖ��(]f\�Ɖ�witZ:G���u4`�%4,d V{�!�����.���XSMɢ�4p2º�JY5�k��8J�E�X/�n3�W`J@�IL�$�.B���q�?B����c&	rJ�\`���(2@��\�]���ԗ�oi�o0�#��H1`�V-L'��	~ٽ�"`� �� Eh)�i S��8��$0��a��L�bCe����.�����H�N�e�B�-�
D�k���>�:���Ⴤ%i$u�	��� ��B50D)��L7<!�o3�%1�K��-5wg<X�#0Ď
e8��3��إH��rb�������R)fO��l�'O�����F���)����q!�d���ˮ���?m���$c~Bqں2ں.EV� BB�|�N$L�2_�;܁����y8kf(J#00�2|�&f�$f�M�z�@����N��D��%4�>�M��1�S),���ɱ�ύ��B �wL�d�g�,!`-�# b�d��:&�����,� #H��X�bEbX!HT�A�@"E$b0�`�� I	3��a2���E���X4��BI@�B���\}�}�ó�,{�WP�����.�"�M0(�$��c2��	
��VM�f�}/Yj��~����uG�D!4$���"D��H+�_��vd5�:��5!�� (�
H"�X�� BD#FQ�!��
gR�\�J�2��`�cE�f�L��kr�x3���1�p�!>η�0cG�q�U�JoX�G��r� R!B�*���i������@9�W$BB����\� �L��9u�������$/n������spF�#c�bR`JR�x�1I���<����RnY'��5��Hica6#� -�9)�b���Hdɢg�f3F�^0�@�l�F$!���6�#1� �E"$ ȅbnH�c;�ŢD"Dc�%`D�H���^�:���!"Ak
�K
�%pB�!B4!R,a]l�p�9���XЍHI��!a���`�$�:�z��:��%�D��HЍLJJ�����3����C�-.��8��H��	�Y�3�4�M}���Ѱ E�C_}	q�s�7 �8���+�%� HjCD�v}�SS����sZ�v���h���	 C��}�;	����;���X�	 �������!�',�	���K��k�ߴ�NR�a�!	|�k���;62-��lF��HF6G+�$��!.#%0F�em��8����iBJ˃$���BH�HBfhŚ]H ���+6$�=�X9V�4i�	�N�V @�!2��1���Χ7������BBB,XP���3
C[��u��?=Ԅl�$*&Ƙ�� ��c!
�$��Ja�$��$i�\,��F�$	�����l$$,�����dܰ.� B��`�p�Hs��wIk9:.���,��n�rCD��9�2��8�X5�0��F�H1��onO�d)~�9���s{ v�Cp��H�ҙѧ$R�%�n]i}��լ�7�_z�%^+�u�W�:�g����M��b�`����4�����>�9�' �P���P��D�VEjF���8�p�	
`Qc 1�p�!�dV4$�X0��bFSI"@�YC�oP�ɐ�)�abD$j�(�<{�����[]�mQ�V�m_K�:t� B@$!ZR��ݝ$��E�BR��!cqJF�+X���^��˽I���"o�SW�dـ�/$w�����H�>LA$��
���5"$R+� �01K�r�.�pe���p����I��R5��D�!YB�P�1!�Ѕ��0�)�I\H!RT!��]	�คA]�_$'hf�TT��׻h��WU���Vt�*�*�*o�\HLwyM#D�wC�����.���y�7<�/���$�
d%1$)3߯6�zv2!�˳Q��=dϩ�?���0�2F�&̱�ӷG&߮>��f��W��(�o�E�P���_^��75�Tʣ3�=����z��˪���_ٞ�'}طh����*��Wp�XWͤ�IRI$�    �      m   ��m��m�  �        8mm   ;m�8 $H [F�  M� ���h   ���Zіb�4ݍ��)�U����*ʵR��;`mm�un��/I��c�lT9j�I�55@T���݁:`6ٷm$��-�p��J���'�����r�a��Un�U��$���WIe�6�BN�������t���qmm� �)��   $��m�[��ݪ��-U�@ 6��-�e�[#s�:�e
Z�w��=5�gm�I0P
�Jۍ���6>���0<�]+�T�I��8�H7mh�R��U�m�eXA�着 ڶڶ -Hm��%�ȍu��  m �H�m� m�5���m�m����ܶ��l �L [@	l��M���V�@ m�    �  �7���[ J��/RUg��-�H�٥k9���L�J�u7d�+lJ�U]@  m���b@;m�m��	��Wm'H٪M�h�m��� m��#m����6����ꪁA��ƈr�]o�U����!4E�4�WV�<���P%L��S�-����U��W�����m�:@��6s���K/  ����$ �i��ۢȮ��&ͳ �����ʫ+UR������0�k������5��8��-���V�0����W��
�8�2�UU5��t��[%$[A���-�r���[mUK�F5rnJ)Nl�õ�29b�Km��5����/N���ǔkrpYv��F�U��]]1�ݔw�ڇ�Mc�w�X�z<L��0La�9�UyvmԫW`�
����X�\�t�*۩�d:n7��75UP  p+;Mזv�Eݛn��[]/1�S��֞ L=��Н�	���]F�n�j�j��|6�]�	V�`=)�QJ�U�+�kS���������ι9��7j�������E���*��iWvj����͏m�t�����mA��g4�����C�i�٩�5�!u�;�E��^6P8��X�
�v�N�J�PڗJ��I�'B�����[Wh�U�lT���w9�I�8�I;y����N�B��M�n[��7E1����n��}�[UV�*��AU۷,�q�$  8 m��m�h۪��H�|�X�$zm[@gm4�Ȱ@��5ą�j�8%�-^���$ ��R`K�D*��)PA��ͳUT�*5@\�,jg���  -�m����K�
��*�e;3N�XN�\�� �M��pͶe������U�U�B��V��8���֒l�>q+�Z��r�@�	�Am�$pw4 ]��'ۣ��   m   �l	-�i�����A�U��!�ҭI,�a�i�[{  6�mm� .�I7k�#��[R6n���Zd�Km�%�M��m;n�  �`   �m� l   �`�`  OH2E�@�k��m&�F��m  `  @h��6��I��� p� $z�t����.ٷgmm���k\ m�m� ��[�am �`l� H���   |�Y���;`-�� �6� Bޭ�ƴ�am����m�$�rہ�lK����[l��m�l ��Ꚁ�`m�   m��j� ���� $h m��ͳ�}�>6���a�D� [d  �� �� �`  N��6� �;E>�}m  9:Y�` -� 嚩[S��Y�,鲀�a=-׮�  �ؐ@  ��aժW� �� ��nݛm��k�8����` 	6��޶� $I!m^v��u*�U[Wɖl�AU��]�j�R��Εm �yۋֆ�� �m����Hk�l  @ ���j��m�	    6� Kh  �bI��}�ߗ�	ء�q��j�V��ۖ� $�i��m���ۻn�[M����UF��r��m@ �` �`l�m� q���p���M�@�i -�8�m�  �,�^KZG���5i�rS� [@$��5��[E����l�� 7m���h   m�6�m� [@� hh�֛9t�`��6��`�  @m�mn��8+��T ]���m��؊�X2F��Q����m������m �s�`$ ��Gk��� 8^�Im  ?�[u����� K/Hu� 6���i\��M��-��9V�3d�QV��tm�P:�q  -6m��vQ�kRC���2�l ��   �߾�"E���6�V�I:Uēk���kYa��m�3�p5��] �u�m�m��m�m  .�ۏ��s��$�ݐ 'Z`��ZM&6�l��Z�M6�@ ��=$���˭����:86�8�.ˉ�{n�n� :�&�p6�	)����s����۶2I]���k:׬.v�rU��;Y�'�DL���@W
�]r=��kk5@鞺v�;C�-��9���K���)�]WO)�N��Hq[<K&����g��ӭ�y������[sUSj��%<v/�]�����T�B���M9�HF�&���H�m���LV��z�A�[�g���P2��֌��z9�cq��Ԫ9z�D5�n��n��R#UuV�j��<į2Y�`.�>
�e�5n���lX�*%�n˹����J%=]S�J������FBR�B� fGn���j�Ƕ׭�j�	n����(�qtF�lpD��3�]�D�� p�U`�Vp��r-5L�,`*�ڂ�ݰ��r��E��ʯ@R�۔`*���Pm��-��6�gAe��l���d�m�Y��- ��]u��� 6�N�6끶�m� �l�d��-�E�&Â���z�-I��g�ܩ,C�nv}e.��e��m�5��\M����p�,覭;S��;iUX�@���v�M�#���\ݥ��9:V�Y� $�N���.6蓦��W�m�W�I#]l��\�Om��u��gO=����՛�Yc�,S��ᣯ4�tny��0����	���o��fͰ �m�-�$t�'mdí�Ó�a��kkDɮ�[� m�i��kp 	:�i$8�ے�UR��7>� #M�[����eU�j�(9����Ih
Uڪ�ssmJ�[WX�EjU��{mu   �[v��8���6]nmd�m��-��"ڇ6�-�m[ �Ű媀j�T
Xy�4�j�e�i��    h  �����I"@_�2��O� mR��:��C�ڪ��J�t�y`-�ܪ�x��z�1S�o8���3��fj�r���4�V�Ʀ�з���&{wd��`�����x�VV�����r��ͺlP�W�����B�=��@�l�g7m����m �M�p�ލh		5Qev��j��U�j�%89'7m�l�(����8 �` 	-��襶K֯m-�  �m�i6�l��m9�l$m��]�c�Ct��U�B�UU�  ��K-�o[�Y�tU��Ž�%�����{9�S��@Vm"�"s��*�� R����-��C���$�X�Zbiu�p�S�l�:K��g�66�|?*����J�U�Y��dN� �EŀN�R�6A�I��Uk���m��gY�Ӕ�������H �Z�VNtF��v]�j�!��a��6��v�m��ce�-�M�  VPk��ÝM�U���a�[@ m� �Yg�>���H��6iCc<lʴ���kR�VQej�vj��6� ������ݱ���^Ռ�v|���<�i���ȋ��7�:jX�!awenV��I����J��,6�g7I�y�:���&�*�m@  x�6��5
��KJg*�0=�뫠� ��Z֑���j�mh��H2rAJ  l    8v�E�Xgm&��]�g����;l`V�E��E,��ʐ �P�m[Knղ0 h�h��-nÕ�z���Ţ��N'.Ö��j�V��VvV�ȵ:A��ۅ�*����:Km  ��6�K��n�����-,[vT �M%U@U*��������J�HM�s^^il���I��_���SRKKF��[UJ�6yٶ�ڐ��,���<��7�շ�s��n!��P��*�:��B�:��g^����s�s8����<�s@t�g&ڃF:(Ѕ���D��m�+�m��l
�:��4ݜ-�4����۶u*�s�s�g�U�����$�[�R� @   [�җx&�`�	-�kt��&�W 4U�r�w$��]l��`52�J�Pr�.�\S{]��    kZ�oSn�p q6U5s.ae@j���В',���]�%�$-6�
L��r�m<�͠bv8*�We+)����o�$$�[��6�� �6[�Le( [����3q�TQAU4)U "��@ A� �` "��*������
H  exMF���r6�A�P�P@��)�	AF��L�+�t��hM��+��3J!�*mF!H+��*�$ �)"EH#�/Du���9�4)�$�~H$ *���CGPع���I����4��A�@~b�O��#�z|D�@6!*�"��M"
0b-E��:�Q>N�����hB�� m"�t��d2A�$j�q �=�Ml_�@�B�ڠ� x���Sk6�U��DC#�̀1�����>��D��>A,R"���D 0��(@�����)P�"�P*���T�9t�����@0#�B b"���� �D �*b,�c�.C�� O��Bh�U9 �A�BEbF)	DY�N��@�!��3`H$`E� @����H p ��O��pB��tV�PP;�*|)TZ���.P�+8�h �tEWj=���1V�bր��X
�ā`�"����b,�XD #VE(E"�"�	���ǻw����{_��UP�m��e⪀���O7 9N8�ګ�:�R* ���1�Z�	q�����ŇHԪN��H��!�n����P>9jUS@,�I�Y�S�v�Wgi0 6�`֖�{��Y�үL��$����8n6�F��ۥZlQm�U@ZRT6��h���J���t�ē�9عێ�$�}+zX[���բN��!��G���j��8x��y��j!灍n�+sV�mXcys�[=��c]�h�`�����;�x�����ۚ�a�ҙ݈ �-r�fS�c�ۆpm�mm$[<]V�P���C��\5k%tJK*��wm8�Zs�V��Fn�̃i]�9��R�km��Pv��C[�M5/��P����ڕ@V)	nVy˴�f1���i��gU�q�P"C,��1F�j�U[�Y�P)I���r�e9c�.�Ċ�hU	.uV9�]�:F���m�����Y6�Yv[J�\����Ř��,rD�[���R":��AN�n]����۰��j��epH�0�63L�;���7m�6�͎��!v]�I�a�j�;Ɵ=����{H���U�9���s��;:�c6Cp78L��zy�ݖ�pn(y왌A�l]���፛\���ɥiyyNd�z{]���ûO\��*�.�a�\A��B��C��&�$m�ƽ ���rY%LA�Ԃރ	�T�P��Jɐmم���T9{j�6f�����"ee1�*��z7*���N��@ T��*��U�\�C%��
��H���\�gwe�Z�`7f���� ��Һ�n�"R�p;�U@]���@K�y��I�"��W' ��"k鎧-�m��aBk�h�Z�xKb�!�L;5��s�l��1+ī�e^^Ai�=�m�l�y��͝�q�}��ǶՃ��t�}�Ѩ{�S�p=:�5h����p��mݫ�u��6��jlQ��s��
PuP����/z�USmv���E�ǘDڊ��F�;ی�2�!�-�L�9PC���&\�+�=J�cn[�тq[t��*�/Dw�h���m��c��A�ư��������gh^�낖�3��.b�Ce� �H l�Vx꺌���ۛv�m����V�u� <B��m��:k[nm��V��M!d�{u��B�[=�'u�,ٶ�l�/�l����60\(��<����{�~�Ͻ���|�9wnܧn��"��8�mό(;��.�+�^0�v�T�y�Y�fu�/����n� =�������ｵ�3�~�r����B�YQ�	�z(0&�遽��hN�U���^]Z/1&�P`M��{.#`���<g\�VB+\n[F�07��0	�z(0=eK���Y@�AJ�Sz)C ��0=��`OH�j�Kt��K���.��Q�]t�<���6��=e�"��n��V�i�m%��٫��������A�6GL����%����-�w.�ֱHZ4i$i"��1(��/x����؆���nL��R��3Z�-!�6GL�JΉ�wH�}}��ı$	*�)^*`l�P�6tL��~������|׷]��ԕ�,���ܬ�Il�0='b��U���?8��=tæ���ٍ�u�:L��x���Y� ��ݺw�l� ��qeļ���0;dt����N�x��yA�+�-�>����\F�3�˰�2��M�1{�Oі���]��0$��̝g�U(���$��0H����D$����䌎&ޠ-@-g�)#�*�dt�ދ�>��P�M[��f���p�dt�ފP�'tL���]/까#��մ�����C8 �n4�uOl�c�b�h����팖�lsHY[�B��m�����z)C ��07��__d�Wk-*�Uʶ�ˈ�䖛<�=6g����fmlw���E!Qu%u�:[ ���	��f�I]�n���ɥ�司F�mҧt�۰3�p��4��̅��P�
BEUq~��~��4��7�̈2�,$�t�0&rEl	y''`�ԷDn���ź��z�װ�n��x���V9�Q�gX+$�����s��x��۬�tW~����l	y''`��#L�7�A��r��1�2l�nt��rJ��{GaP
ʺK.��;�0'��`L��j���MV����`w�.1�lrJ��v�$�������?U�&�K`zr�\��x,Xfe���x��۝*���������ͭ��Z��5�����|Q�݈4�.y�&��	�õv;;�������[-��;g��W���y�.驖���G3۝Ϫ' �zy;;/<b@W
b-�:���ɸRwY�`EέI��x٪��X�F�4� jB�ܫsu� ��Wru۶71x㡜n� �uss�];�6�w:5ڷ2�Nc� �����$�E���q�WO��c��s�@�\m�K�1��@�|�����\\�����gm��h�^)`#[�n�Z�q9�1���r�X����ʋ�+�;S���=�ϲ����遻�*���eڻ�J�ˢ�r�ް?d�?���rkL����L̻�b�fB���e�nW�3�ͭ��ΕlgD��r��q3
�e�)lmWj�D�����>�������`{�A��#��0�RT���Ŗ�6tLo(0;dt���.��Mt���
�Gj��qT�H;,��N:��<�AQd���qO,������컭�g���/3��~�:`{b���꯫K\a��zl^���v���S���rO��tk�{H�
�d,��`�BXd�#�����s�}�b�����������'�V�j��x������������w��w� �
��+��c�{Z�O��zl�ގ���[ �}v��Ҳ��E�����0=9L�ٓ`u�Ֆ�EI��ƂW`9Oٗ���e�籬�^�帋ǡ.��c�t�����X���Cw���)��������i�e�̴˺V�0=;����������F�`+��;�JA�,{��ɰ9�n�ER)*��^���m�靜����@e	e�������GLNR=���d�Yېp��%N�KM����Ӕ�`z�L`{yA�����Ϊy��5�ɸ�9��9{S�(T��&�3�E#�-�.�8ac�um4�1SӔ�`z�L`{s��7z:`N�6�աQu-v9,{��ɿ-$�>��=��綶>ˍ�͇���M��j�X��?[w�����`z�L`{p��w�^U�e�/�7z:`{yK��d�^��UU�U}O��1��aܮ�$�lmWj����֒�wޜ�3�`}�sk`s#}������KW�Y�-�u��l��=����<عlY��8���[v�	�\Y�0}������ޘ������.���uaR����31[w:[w�����`{rK`wӑ0�bY��e	+`n�t���0=�%�=���r�%ҵiP�fY���Ll���Ilnt�쎘�^�e�BYx�Lܒ�ގ��:`{d0.���K@�Б�kDk؂�$�JG�� V���Y�U���)ڴ�x`�7Fc4��x�%�®Ş˙ტ��c8F�s��R���:�9�Ѵ����T�/޲���v�Ȭ��ֶE�5���Ɇ�{e�%��㡕/:'��8�	n�s��%��>��s+��c���Aѝ��ñx��:���,���mt�`g���2V�a��Z6-n�kd�۴�������~{F����&;\�;7m��f�\�ost�ݵ�kgZ�i��,��Q[��C��g�s���ٛ[� 遷�cۄ̺�f,�-U�T�ݑ�� 遷�c����i�
�3˺V�0=�����P`n�t��P�yn���2�ZHT������w���A���A��J���V���w���A�ײc�q3yHĹw^gA&�d.��7ST�7`۩�Yp�[8��\9��Y
���I%��YM���ͭ���0?_��ʪ���I�p���Y��\g8���&����4k��T ��R)�J�I��d��g`���ml�n��.���j�`q��6���0=�)� �t�Y�����j�Ōw(07z:`{�S��d��%�d0X��e��J��`~�D���N0?fv���Z��QuU�ds�]k�4FK��<����W�ms�%����Z�v��h�gkR	W�6OԘ쉁��쎘V䛏V"'H&�W`}�w�6}�t`fn��?fE׵J�̬�D��uΜW��3`l���ݑ�6�V�}�}�Ԭ��\J��BЗ"oY6�s��YRD�r�C����H�I��I F��K���;���`h�1�2�,޻��[!����	$T�C@5�j���S��Hf�;܎S��b������Ȭ�"�i�|P��$ChbD����D�HDd��`D�U�X�*�*��2d�;j-]k9{1�>&��p�ڗ ��N�H.��6�C�D
��m! ?�p R'PP>M��d������5$����~��yk1+��K�%L�0=�0zN�ԩ*J��o���8n��U��̳-f*`{�0`�&�\6�fmlw ����di���-�8�^�&؞5�Vt�rm���.��Lf��E�9�j�:˩k��C��v;��ϳ6���w���:fz�$!
��h�Ęؠ���遻у ������m�B�UV&X'm[;����0l�����V�� `�!,/b����O����`{b�%?k�T��M{߷�'���.�����e��}�vW�]�qp�=��9�hP�~�q�ۮ=:Y��Ձ�{�,&�&-C��Z��wD���{qd��O�z�Fo[(�)+������k`}�sk`s����a��6k�O9\��$�Z�ަ�����]��X0=y���di�Zִ�g������R9dq�J���`��~���I*����2kL	'`ڵ���Z���{KO��zl�=����4�iU�M��n����ع�텬�ŌwGL��?z���� ���u$؟0�A�!#��G���"�j*ܽNһ(�7l�thtE�yZz��"��t=���.�`�Bm�c)�@�ճ�Y�!��-[��SQ�s6ll�ܱBݤ8���gn�A�N�Gn��e+��v�OW��۳�ZJ5�Z��dLVW�݂Ζ���m��p�� ��n��u�9���f^��I�WwfU�;g�(zی��4cV��V	iE�ii&����n�����r�r�C��aq{Sg�;����jő�vћR��}`�����4�Z��������0`�'X�#L�)�.]e�@���Y������0&�&e��t�Z0�I �Ș�0=�0=P�'Ҋ�J���LwGLގ���D�ߧ"]bV�����b��GLwF^ɌwGL}��>y[�܆񶱸%�@86[�k�����oQ�E7�gl��aWљ�U#4�r�����0fN�?fF���$�Xz{�[���q҃�����6�{��Y�IR��mƘ�4��2>U|�!�����q���`�$�`w=�k`d��m߶k�����`z�%��/��D��-[i<��Ű>�{p�y�6�w=Ű>�k��8�hB�0����d|������Z`d��Ԗ�?���D���.���U��I����8��mF������1�U����w�[��ڇ���N���<��}����I�U���f{p��1��R�q�X�F�ҪJ웺��k��2I׺�fk�OX�*��j�U�3�����9�bjb�X�	 N� ��6�AbFD0B@H� ��:A�ZD���kK�Z����������c�	#��i]�رS�U쟽� ������釒O=�ql��Q7Yu-v9l6�N�5%�7���֘�#���z_�<~t��8�,:N��UH+��N]фNc1������qs�������J�(�j�s��|��L�4�̝��I%\`g��1��pq�]a"�����$�?�*_$�R�߻�m�����`g�5�i$��&ϻ�p��]Mհ&ow���$�5*�w�5���L	��n]:ۉ��k�{Z~�����3>��w��I���� �w�8�Z�^_Y�}^��3��IK\VG0=ܠ��GL	9El	rL`*�����7����Ҳ9���B-+qXh��&�a�m��I�5��˛��k4t�Y�ˢ2,�X�%�x����0&������c��c�B�AXF��l��+`K�c��	$t���%��V$;�c��װ1�d���{?--7�{�[������3,r%c*i��`e�`I#Lޝ��T�y��`m��������m�33k`{I-j�����ww��'T��QJ���T�$P@���#	ޘ;���6���M�m��eX�[)�ݗ�q�@��iE�ڋ#�����q�6�Q�89��\e�A�́�:�ۣhJ���Q�������"���.ƶ{yx�ۃ�BMv�:y�I8����\��������/5���ك��q�籫d�]ڴ�m��ێ��=������s���q]c����rS\pi�,p5���9u�d��HL�0�-�[�f�O ���ۏ�����-֭=3MG9�;r�ݩM�er(���"�<E��"�����w����h������`u�d�ɘ��\a�����XzM�HӲ����^���-�Wʒ�~��7���읝��Zl�S��
�VYRJ��{z�ɑ�mU%W~����y6�^�^"�U��h[n�����ikIO~���Ͼ�ݶ�'Xm$�]������\k����Nʶ3.W�=�<�z������w6����A!��؈��p��5���܄�e�̘��:�b�+�z���Ի��ݵKGul)d��=�� ̑0:tt��+`K�e�]*�U.e�3�I'{��\"��) ���H��#dD��q[��Uz�~��1ﵦ����L�`K�%ԳYa�XZ-$�::`zr�l�D�&Șܺ꼹�	��]	*`zr�l�D�&Ș::���$M�t��#�W��r�N��ӣ��Q[ ��}.��W]pd]�I�˻c�8m�ݸ,n �6�.�\�3M�%�iʄ���*�-�w"`t����+`:&}��(�Wbe�KB�vs���ɳ�z���g��`��`udǊ
[%�Q�e[	��=�ԓ���5�V$#�� ��w��o�ԓ~�tjI�w=&s����_$�Zĭ��:c �"`t������r>��!U
�(�`$L�0=�El���TH�_gn=Zܹu ؉��j"��/=���nnJ��T�4��/��Gk&ݥJHt���+`uΘ�;�Ln]u^\�) �Z��%LlQ[�t��"`t���-�bX��Y���˙8�3$�5R��5��{��1|�LM
�+�*��l�̻�����gm�.$�R��'��q����x�(�n�%�-�����I%������?��6��]���I��K\��\	{e2�iU΃*(V������}05�����Շ���{PR;JƝR'e\�e��.d� �N���l֘��G{jt���Z얽�םɿ$��a�{Ձ6kL	���z��+�o.h��9`��u]����ww��f�T����c������!H�"��YV��UU�R�ϧ�y0>�w�[^d����������5h�S+�l�.F��/�/���<�}�L	�`q:J��Bf3A��W1�H�B� HH@�;��j��'�損�@rb9 rdpd>"Ș��ǆ�-"p� �.���2���6+�18K!�D��2e�B!�B�2�B�ق0�mj� �L�F%s���B �L4�;I��l*䂘H�>w_`�##R�K���/2�O�(��+�0pD4r؉�3����0A95�R�s��uݽ���?����J�Wr�oP-� M�Θ���p�V�ޞ01�˷9J���Y�K	�닡]�&����mI,�� �9n&c%�>�#k�%㊐�r)UPTMI@c&n6c`Z��P�����h�P#��h ��G%ltqiF���NY\h+R�[N��H�T��uh�v�EI�,��&�x���ou�\�l����[<�x�UƁܡg�׷u��v�y�1un� ��{�W;s�^�#�s��Y�:s�yz�8�F��mD��g8[����6i�T6A|�} X�k����±���֤*�9�jr-Eъ�ڪWl�Շ2�UR��r�n�k�j����WM�.F�)T茶�Vӓ�:�'1��}��[F�n�U�]f�C�nw������T:)V�ݨ;�UV��-���]=<���
AeY�OU!�;� m�@��4�I�UoK�)�mRp�旀�jX���$]�V���)�=h%F�\�ўZ�8�������8�IZ��e6�\m&�:�s�l���`�eR��;viq����n��t��9�UF�8�;l�2t�X�jN"ᗢP�3����Hs�U��*[�s�+[��y}�9J��G��s�[�m�LwJ8���i�nݜ�����b{r�+nͬ�GPu`I,�ۧ�8fN�b��*���sk�2WnU��6�lW���!�8����B�l;I��P'����,=���t<�)Gv֋�kn�o\ʺij��
�����h��lqH;GV6U��vyk��Zu[+g����8��8� �<@T�Ҋ����[m&Ω��nmr�r	��;�.�6���t�͵d�J񕕪��f9�Ci�c��Umt9U��lLl#�w9��VE��F�@�Wx�Ť+g���u�s�:��	6����U���S<9�9:G��	�@��k�1:�Z��z"�"���Y<P��iOl���6�k�'�[��W�-�Ԅ�Wm-��&2�m��u���s�F�Y��*���9�Kr.P��(�����؅E����"��� 	���õ ~ً3����0
�u��tj�wVZ�0*�3@�a76ʒ��5�c�]������r���!;�3�� �3�cb�l���VďD���&rrm�Ό<�1m͵QR��=n��-V�B'*
4���O�=�c���Ri� ��0�YB��K��f2Tzx��Q�8כ�<�ܧT �(�:�9��^�{fF�v6��x���9�8.2��2��P_˽Mˬl��9�9㍓ӻ1���=��d]��N�����6�q�+�����Pf�A��B%�>����q�$�0'�kR_�77���Ň,�ɡV�rES�́�����-~֤3��ml߽7�:�̛�I�5ُɹIFYd�[j��{k`fv�{?~�R���`~���_��v�q�P�uH;*�}T���}l�7�	�a�J�M��w��c�J;�U��W�gr�%���{��gs�[;�c�̦X�e*8�M�R���ͦ.�vn<q��ڱ��ָ�]R`ڲ�%��{4�D(R���o ��i�=����/�T��R���߮����ߑ#�c�A�l�`g�ͭ���DF$�$NAT�C�DJDA �����I�$�;���f�������aAU@���vu0&�`�:ͪT���֘�Z���O��l�7m����o�7�	��0'�4���RU\߾��������J슷-�33k`{ZZI~����?~���oD���d�E�(K�.I�rvɘ��KrK��65�s��ج��s�����w�����͍2Ӫ��ɭ0$��`�;�T�Ԓ��p>������C��7��A�V���m�R��*�ɽ`n������I*ZZl��|W
��Z��[�{��N�ѩé�N�U�����ލ��m��G��X�B�6�v��J�ԕRK�o�y06o�0&dv0��kZ�R{=(}���TQƠ�U�3���2$��2~���ް&H��h�O"�V��H�bv�B�Yf5�E97f��י���9�4ݲ����[����u�W��u�㲮��m� �w.���m{Z�K�3��������B;Y;mf�?L�z�$���֘&���d|��i6}�@�גvE\�݁�{�[���5U$��M|�oXS:K�;�Q��KU����k_��Ҟ�~�l�~�5$��;�I�ǉ� �7�~��gOߩ�p�bqH;*�}��6����f��7Z`g�4��vv���se��A�Ӷ�d�l�[���÷gtm�.�� 3�b[_���z+�Ϧ�>�e�{���oX�`g�5�UU/����`gc��ʣE
T�Ym�w3i�U�T�W8}7�w�c ��שU*l���%�Uj�e[��ml����J�+�roX7Z`K�!_"� �S�ʶZKO���6������[$�~�{�`}Ռ^[в��{c ���ʕ|��o�yx�����6̀������2 @��7J�F�Z��ڷk�e{K�H͇��=l�rz�	��r�u���8�G�m�tH��.��`�uVvp�.�qn��l�b"�\��-�F���H�����������z��.�s��|Ym�1&˶��Q�g5�����'�sƚ�j�@��랼��<%�]t���S����u;B�8���6���@[bΝ�s�0��ƺ���>���w���=��>��u�=�[N�
�;���U�.ؓ8��)�м��q�q��--���o\Hu�n[|������ϻ�[��6�$����]��{)�+r�vKU����w6��M�ｸl��]���mo��M��{��8Z18��l����Od�6�Wrn��ܚ��K�j�J�mZ������&�����{k�6�v�ٶߵ�I��}q��#��t��T�;iv�o����o���I{���6��{�!�6��\.�m�k,M÷^,l��w
�emu�%�6���7�N�t{%D#;���>�P�g8�n�?��ٞ�6�o�w9q�ϻp��䍿g���6�8y	�QHu��e��m����otF���\f��>�ն�w���6��3p��ֿ-[[���n~������s��{��v�o33��~RN�{p�m�w��9��������E]��m�kR{��˜m�����y�g!�6�~J��?m��������lu�J�\㻽�������ܠ����'�޶��w6�J�qH�" +�a"u�G���i:܆w<���	I�E7��ٸ�d]��>c�y�ݖ��u�6�����m�����fg���6�=��m���߁B��Q��lvS�m���]���j���߿qs������m��f��<�q�_�W��������������������~��j�Lbd6�l@?�}�{\�ݶ�w>�Զ����er:�A�,�|c�ZJv{�Sv�~���{���g�����{���{�Q�ʖ����]�m��33��m�kJfo���f{��m��f��m�٘�}d*PtqNշa2�J�x-��u��)ۃ[Q؍Y�1`�"�9�u�j���V��m�_W��}����6��3j~�\�����\�m沅�<���E]�׶�}��ٽ�1�^_{F5m��w�7�m��{��ʿ-+k}׿l�e�:�m\�m���jm��3���?i$��2�����縹��a��b,�F��uʦ�~ִ��{�������n����wf�m����kZ\�/>Sm���o�
Y
F+U�Kk޻��������������u����:ys���i$���UZ�Te�U�j�����g;E���vx�FN�-�:�X��wwo��8P��������o���\�m��6��m�;�^��K�m�_cm��y��B���ʹ����mM�%�jH���ov�{��7V�w�wf��*������s�ڕu���Sm���~��m��+�~�ZZRO�=��6�_��6�o�Xd9S]`B�[W8��Z֤�߫�m����޻�ۑ�;������}�J��E]�׶�fg8�~I%��qN6����s���ە�9�����E�w��
��|p^�벖&U�Đjv)خ ���H��Y'Z��\m��W������Ԍ�0T���Zxճ�Bq��l]:&��&�c�v�c&i�jŇ�w46zex�s�U����De�Wų�f�re �=�q7S`.���L�[Q&n�lY/�P�qv�����܆�X������ɴ�5dnJWH��$������K�h�����h�ŕ6INq��GK�[C��m�"\L�v���?ik[[�{%��H�m^����mM������m��+���$m�=�-����vY�[kh�G\��ly��9�$�������o�������fnm���w�
:J���%9��;ۅ��y��\������=�66߳���6��3drP�������ߒԞ�{��6�_}�����]�ݷ�
��s���um���?�0�XB�e\�m���Sm���׽�x���}����o33��m���_>ql]��Z&�M��Xfn� h�Vp����	nq>b.l@���!�U8�o���s�������o33��K_}}y��yx�'��`�vS�v��3��|0�����C V`L A ���dʦq��DP�))bB0���a+�Q�~T;��������_{D�m�����Z�>�(X%�]�+s��7V�}�{f�m�s�uo�C� ����o��6��_����;��,���#I
үz��{#�www:8{�ww���v���kJOg���m��{��Q�Ɗ�nʞ�m�sxs���i%���)��~�{��m��3i���ud	�ElEѩR��v�*� �ׯUas�pv�l�WLG/P��ܒ���n��X���)�Ͷ���6��vov��1���C����ߵ�ov��~��7h�P�OM�i���\�m�2>���G߮��dk��K��{w{����VR�e\�m����m������E��#�颤0`��Q0Q�Z���T-�\��H$~E)u"m�ݎ�~9�,�������I�XL�v�it�r�b `2P����dt�X�e\�(�BgB�`��L��)�0C	�WDBdu��-�l�I�$��-r�&։�"D�O�q�� ۭ��xP4�H l�j!��8�� !�:�o��S��� �P4�Y�U0�}�����m��{��m�Ɏb	j�-�M���'����6��{t�m��g8�>���m�b�q���R�Nq�������ޭ��^���\ָ���dp������=��߇�0�.�^�iA�-;�;���u�Dq���q�a�¯��x�o��wE8��Z|�o��~��o��ڛm�����-~�km�n�m������;e���m�{�w{}c���#��ww{ѡ��ߦg9�$}��ڮ���"*��*�m���^�ݶ߹�fj�§�9�?~��{���~ڛm����#n++��l�8��S﷙�m�{�ٽ�oםэ[v@R����m�37E\����n�M�wrI������:�wwrGz����C�m��Z_f��N:�� &���jA���؋h��z�b�jJ2V�f��8���,!l���������m����m�����$m��{��m��p��Z��abX����s��ww{ѡ��ߤ��z�sjo�F��'��"�YX�vS�m�����|�3��~JIמڛm����s����YT"5\�*䖛m�R}�߶�뻾���;����z����C������0�[]lv�d��m��sjm����{�Nr�o}�Y��ۿ�ݛݶ����ߟ�ڶ�ݹڧ,<��^�e�.���<�lĻ���\��[��{l{u�r�\DҚ��ug{t�s��::��v��y4�{[�-RЭ��E�^�	���̵������C�}���;�eg�xKu��S�x����(���rN��x�-���k�[���=k0�k�$$�P�vB�Z�d;+���ݸ��O/A`�v�^]�ە�ȗdkhru����w��?׻��O�~�i�E���Xݎ�4���M��0;r����fCnP�q����?�����*�m���f�s�������o�fqs����mM��x����QYU��s����n��֔����qs��מڛm����絤���{ۃ�r!UJ���׶ݿs�ٽ�oםэ[�P?
g9�}��{�מ���m�߱��`Y���W8ۿ\�q���{�#L6��~ٿ����4�Vʁ�`���v�=���d����~t���L`v��əe��O��fXwcC��8ȡU�Up�s�e�V1N�v�S�WimECvS`�s��F��2sR�U��I�BY��F���d�݁������I-�� e0 �T����}�I;�/�w���E�W�%���K�T��~�����*UWy�Z`{wZ`s�w���PGU��f��KIO{�]2kL���JJ���� Փ���fZ�EZT�,Cw�������6{ۆ������ʩX6�j��%aAq��k�n��llo]G��lˆ6��_���˽���UB��$��}������2l�ۇ��w������:YF�bT�������GLN���M�{��IY��6Wl�ܾ6I���L�����F� �G��{K`y�=6b�'�v�TB!�)�=�0?L�0?{�[T��G�(c*�hPc�ɢZ�3���<��������ގ��/.bWx�/�#]Y����^�d����<��OW9�:;r0�����1RM�m�_���lg��`L�֪I%���5���uuw��EuX�l�ۆ������w=��7���/zcWr�Yu�H_ZT�w��`~�f�*T���o'|l���v6X�T*i7j�{KI$�ٿ�nM�=����%T��9<��35�������ld�=�䒪����5��H�]��p��Ƴ���E�n�YH�K�7���.�)��jտ;�����v�l��L~�ٓ�03�`~�}I~���m�6CT�$��dCvS`w������-kJC'�4�Ϲ�[����T�Wԩ.p��l�~h�c�ȭ������k`s&c�o(0;z:`l�e+�J�ݤ�f$�U%W���`fN���di��J��{�[َ��WB�]VG-�`}�n�*�o��f�LӒ[��I	#�	�ED���0)�j��,��t�z%�'	0��:ˋ�wiT8�)%��ۥ+B�gu�IW!�F���v
}e�1M�u����1�g��`�n��臮��v z�6XNH�����)Ń�s-����<>n�e�f��m��g ��1��ϱ�KfcͲ`�9�ۥ.q�W(�Y��&V��V�ٻ$<H�Y�\ݤ�4�ۆN^�8冺����;s�N�;�eɯ)k�J[Ľt�����Z�[����ܧY��������Ȝ:�g�Ѷ�V��]��K[������r�,���S��O�ߦ����`~��l{;���5A��P��ݫ`s;�[��I��rm�&N���di�$��b�wo�x�2�RISd�l�P`v�t��w6�}�����	,�a䖮dz0&Mi��di��%_$��=���x���-�Q0n�l����9����%�;yA���/1Z�̬M�[y����ڈ9�ˠM�[u�# B���ۈ���ImB���" �e��*������-�����T�/�/p7w���3����Fݶ;*�ɘ�RZ�kZZQ*��*l��{#L�#On��}�R�Z ��#�װ3�|l������{=��>�������5mbv�����i$�˛���'�4��9%���Jf{�����ۃT�U
�C�l}#L�W�������0=~���y��;m��{ke�ԯl�T�.�<Ϟ�6������!1���@[o�a�������~��(0;z:`{dt��bŒ[jnP��Ie{�pߴ�fw5��u��̖�RWf�m2��;��s����:0$����i��)!*@���T�J��0�����!O����P.��k�RN������c*�b��ج�����-.d��&}Ͼ����3#LL�\�]T*��l�U�9�1�%��7�fg��>������Ԗ�D(�o�;x`3��-f���۝[����m�θ�.��Eߞ�m׽�
�^�Ud�[8{�����4����%��of�gl�N��b�uv��t`I����}J��'�4���߹�>���l��ۃ�:�Du4�j��֘s%��Wy��07f�����������l=��$�{=6{��jI��5&D��#� ኛ@�r+�c�٩'��Ӹ�1��̜����;�0=��*�U�T���yx���[�;�`s��ݕ�+,j����ネF=�@�{j�p;�˶����/҉�J!U���R��M���ml}���}�}�����=�;�c*��Ev��.�9����4��������o�`d���`g�ͭ��I$��������U�oy��S ܛ��rKg�IR��5�f{k`g��E#��D*�[m��Lǰ&di����������T����ի��T�^+`N�遽�� �"d��;۩'ԑ��Ç;B B2Fdu�c$�RP;��0���D���>��������X$H@�/JP#d @�A��r�b(B0�B8֭0Jb�vA6ԸV]�U�O�0B��]�:F��`��#"��F*n�fs�
H$�Nw{���1�ٶ�[A%*��9�T�mP���mV���-l1ź�mT��.T9�N.���v<��J�&�7y��2��:.��.�M�M��2fj����*8$�
1�[ +���T�.!B�2sTl\�����li���p�!2��,[��L��< ��ҭ�n�Eګ�Pcv�NƗ��SK�쀩�;.�nrz���Rièݧi��ɭs�v�x wn�ܖ�\O.�����Ɗ�9��n�sWY�^�.8x�wm��[;P���]�8 �a���k���cR�]�ɹ6�8*Y�ڎ�������`�B��n�������Էm�T���-�R���Zgy���&Z��m�EspT�T��A�d�̽W! ���a�]��sm�	��n*B�(��DnYِj�6�J���ո#\`��v��KZ��ڶ��t�6�76��aA@l�
ʽRY+�#/c�͓��^�h��cbU�
u�X q��v�u�Yڃ���n�UV��f�]a�6j'v�
m�]Cay�Yvso]�-�	bp�-i�mPi;y8
���=���jz��p�;[7��PXd�wkX�]t\�
�6�;�Q���єތ�;�p���]�)ZA�N8�Y�]���ioN����5Ĉ7a;M�-&��9-����Ӛ̽6�(�kO7k%�.y�m����I�����۞�Y�<��ˊU�.���$[{E���HF��1�aQ�1���K�
��!:�Z�V]�g�5̂�d�s6 Tc����T�vŜ�;n�;C@E*�.���*ѻ��t���t#(f�筜���[��nZe&�����l�@�#(k�����M]]+�,s����`��!@C
��K�V:4@���m��xv��M�[8�V�V�(�s��#>�ݔv1q�`Ld�u��H{`����n�u���va8���h���.�!,���Q���c���n�SV�`�v-�4�݈Θ�{j
P�.8C
UM l��RQE�Xh*�"=M�AP� (dS'C�9��RK�7W�*��NX��5]�Ϫٌ��.��XܝH��q��k�����]m�U�Z����⸮y���Yvr��7�v�f��� \!Ӯ�����]�s�Xg�ɞ��]p�s׸8;G�Pc��զw��3������(�K�v��K&�0�m�YzA��%8�2��v�Mm�v^'�t��=����������J *�@��k�-�Ҧǳ��#�E[Sn��vPM�k�5=0Y-�5��v'�Xn����%w�ZF��(�4GSHv��g��='X��^���d֘ME��廻J�˵W�S �"`{���'tt��{�[���~RȿO�Эʪ��Ye�7���&di��24�'��zm�Wj�N��^����s�[��ml>�]����s�`w��U�Ӧ���.�y����`}Ky�y�NM�̍l}��c���7-[dQEAkU�D�B�P�:����q��k�0k[p;��m�\رm�ae_����`s���}���ikKK�>�����q�D�.��*�Km��s%�V��$�ˌ�~i��5�w&�řZT��4�U�k�������/d��:[vGB1e��
��������/d��:[��3�[|��6X�����-[Ɍvt��0=�0$��*��h�ζG	�x�i�ݹ��#��Z{{Aǫ3�q>n"��K'f碜S?m�[�-�;���GL	{&0'q)��IP1�!�k�����kKI����[Ͼ��};�`}�˄ӮX�V����~���I�>$�EU TQH����W��^�LN��06r&Y�+At��%��c^Ɍnt�{I���-����D�.��*�Km��Ζ�������^����3-����D*#����HJ2R����MO#�C&�v����J�6�K�;f����|ގ�ގ���0=����0	(�ȚMڶ>�mo�6y�=6ݙ�3�����1w�oț�v���w����x����l��rkLI�09ػ"��!TU�l�a�i-'�\���Z`~̍0�U��%m,E�����R�I%�U"$D�\%�K**T�_o�}��n�����wwӔ]�V�����#�����l/��ǩk�����䢠��2�PGcv�jL��cn7Dq���5�U��aW��&����,���b��������l	��[����q��Ym�J�?��{vfrm�7&����`Oe�qY|�D)J���f��gq��������{k`y�=6/�Z	�Th�W\�`gݍ0=$i�/�8�j���37X����Xi�V��;�[��;��;=�3����z�5�&��B��;)��!��Γ�їGRۣ�����e��u���ؐ)ځ��m�f�g!F�2�M�$�]��:l�@�q� ���뭈�N�V�b�v�l����BMX۷!�]vl�Mp#pLs���iێ���q�j7`܎u"v���E�b�'�t!���nm�[=C�]�&�!�[�Q�ݛ��}Լu�k���=y�vvIv��{(N���G�ID���ۼ��h���Ԋ����Tv��X�VN
6�`��u�`��y�O��R�;H����<�=6~��`gs6�q�}����Y"�e��W,X��ے[I06���$����y{Ɉ��:��ە�g���>yٌ߾��%�;rK`n�gw����yH_oc �"`v��ޑ����e��X��*`$Lܒ��07dt���"�v��Uw�i�v��H�u,t�lۇ�8x|M����ۭ��g�������J��[n����~�ml�0N��>��`�.Ձ�Z��ԓ�s�5�D]��T�@
��S�������$��T��ɬ��9wj�
�-*`w��� ��0;rK`w�ͭ�����I��+��U��������`L��324����ֱ^]�+E�x�IbLܒ��#��6��f]����d�v��ep+Ӭq�ۮ9�<j���w�yl�lڹ�7]p��\�ek!j�CnW�;ՙ��>�ͭ�l�0;�K`n�,S.����X���Ę�4��*J�3wz������Y��v�17]pvX�`�˰9�;۩�<[$FF	$F$$���"�R(T$Y$�A-VD�B�h
��to�5$߹��w����mů��K1bI0;rK`wq06tt�ɿ���˳�(�օmu��wKt���� ��0;rK`N�/>��k�Y1E�y1�oF%;f��X'&��Z�Y:���g�*
q���e*`l��l��%�;�[�WE����[\U�m�l;ܻ;3����0'tt�뭫�J�Y���`M�-�:�t����N�03q3u��i
D6�{
�ή���H� ���*��@��*�RII--h�BIi%;��{����Ie��IVb��GLN��۝-�%vml�vd��UD�U��莻Z�p���m��{ �H����M�r�w=�1+ˣJ�լʵ�b�Ӣ`n�K`t����0&�K��/ؐ�f%�&�t�����#�'D����b.�RUbJ��0$�:`zH�N�ܠ�푕v	+)*�0�L6�ۻ�0�z������{��Ɂ|�9${,�n�m[ ��.����0$�4��#L��UBH^Y;�	���-؛��	�t�U[5`�m��8�v��!)ȗ''�lѼ��m���ٵ�z#�vv�Z���m&���:�l�\C-Y��k7Y��ICE���0�l\m�7�V^�j�����\��̑]�z��s����k���շh��6�S7YӸ�����is4-���#3ֲ��h��g�wk�!����C�z�V�9�͹�$�.~Q��Cf�]cB�9x�v�e�wn�m]O��Q�m�/6]ͩ��	�6���&�ӲdgIW����q0:H�N�꒬u��*
D7e6gL�ߓg��mlٞ�3.�]e�\�UnUj���$��N��$P`t���˴��4�li�Bڶ��]���N#��:`M;�R��YKX��I&�A�Һ:`I�� ��03 �˨�jؚ��Lm��(p�ݯg��v=;n��]zi۳���s���ƥib8���:`:&w(03�͍��*�Z�!*��ͭ�ZT2D# �  �e~F����EN#�Vʅ�fc�0Wj�%LgD���N#��0;�땔4ve��Q�&�P`t�:`M��l�+�{�V�ʙe6qw6����� =����n�/�J��ۖ���M�^܄�-ur�[���-��"��t��*$C�!����D��Z���[�Z���?{��.I���}T��a�����N�_bln�Ӳ�ڶ>�&����`ft��$t������U�%��03'`���"I���b���!N���R�
��BGA�,`�i�mL%ظ�8�*'��oĲ��a>�f�i��E�PL�S9a�F��������76a��E$t���u�^/,#���a��P�T�A��㠠����� �HgA��+h�A`�����5�a�
�[�
����. q̤���Ng�`j��8,���G'ȽXɱ\�@�Ű�� �R�	�I �X�$R�0�C��@p�'P��Q8��`��@��m�Bs���L�����V!e%X�ե�gF���s���&��`K�N03'`�ݑݗyk����T����w�7����с3���r�#���8��6l�h7F�@��Eah7��M�:&b��&����s��m2�&���?��-��;�#Z�Xf�����#t�奵��{��֖�lά������N��]]�M�l@�S!�6�:`oH��1���,S��
�%Y���0=s��I7��RlA��6¡�`�IkB�+Yϖ�����؛m�ZvUV*`z�L`zEmtt����.��(��dR!6@'t�J�u�k3�!�r�͍��m�nr����Gk��tv�,`zEutt�����c`EFJ���$Z��,C��:`ww6�fM��ˆ���l�s�ln;����RU�3��Ǚ�`w;p�����e@.���-,���zI���030�0Ԫ�f�L	��n^[T]�/%�0$�w���tjI7�w:�u�R*��ƀ�J�U��*�m{H8&C Ǽ_w���v�J��5���
�c�E����Ǘ�n�N��gpu�{yر[��	�S��ѫ�N�R��$j�ہ0h�ه��ٮQJ�qX�9f4u`�n�`#v3�{nruL�.�礷n�x�pn�dɍ��vN��nF��0T�\b�D<S�-��+�s�Xʨ�2+�]ɍe��t��JX��`��)���tz@�ΜRVu�<�O����z����k�ctq�۟[wQ�qp�d ����.������lr�՛g+ۑU��;x��tt�=:/ް��/�������T,�Z궲U�3;�[ �2wXn�����1gB_mr��%uk�0N��7���!����ml_wUL���
��rٰ3�07eGL	::`m���S-*XV$�V�%�`nʎ�z:`mΓ`gݸl;�*�-�j���v��{ �V�4g=t�uڸyg��%����V�����"���w6��;�`gݸ{\a�������/ �܍�B�ٜ�ԓ��w�l 	�)Ga8���H�z���9��#L	�`t*�ʲ��1,`M��GL	�:`mΘ��N%���e�Y�,�:0�J��&�֘���	�p���f�Uש]V�J�w3i��9�y���0�0���MO���<����{=:A9¨$Pnջ'��;���)�{a[�jNP+X�Ew�m������02a`L���ظ#"�.ЫE���;$�N#�oGL���*2Z�RċV�+J�0�03�gk�*T%�\�����-�6A����)��0�L�06r�ft�N#�V�F���GB�X�[�ǰ?-k޹��3�{k`fw6�t!�e��*UJ��5�@�<��J���vM�}��ԅm�^'�خ{Cb�a���H�Ć���N��tt���Ԅ�]f+.��e���&�0$����	3��=8.;-I+T�-*`I����gK`M::`wW Ʌfi,�ަ{;��l	�#L%T��!􌊄cE'X�B*�!R ��B#*FJ���B�$ -Q$P��Ba�@"F!	 @B1@"�T�1R�!�V0�Y$��	2	D�����q�I9fz7�ʅT*���M��;�`g�si�&F����%W��W9˳mc�i}�`gv�Ÿ��1q<��p�k��d16��ju�%�u�+��t�ml�07yA��:[w�����Xe#Xa���ӣ��(0:gK`n��[�i�q�6DF�*ݝǰ:���;�0$��^ܖ�Xe�31ZX��$�i#��Ӹ�zQ�V6DԖr��ߎ���F���-���-��J�
��]�^�o��_��:=�]prD�pK�]E�$��7*7M�fH�%&��]A�ۦ]f&ҋGF�3��{U�m�g�m�m@F0磈�{����m�ӍI�9�Q[��8���l���P�p��yk���gavCg����x�78-lv^_[s�Vѭ\F������%X��K&��zUx�C��jp�g{�{�*��K����d���pr^�on�f��ςG�۶��:El�ӻi7n�=�Ѻ���b"��9&�\��$ttW*�b�Ύ�����%�7eGL��0����-bWiSw$�vIl�GL�:`K7�fR�P�
�H�K�%�6q06H遷��`s�3����ev������l7�`f����N039%�'���f,�)��0�L�:`mΘ��	����}2�I,�>�����vǲ�KC���ד�n��c�-����nS��;-I[r:��rʶ_{�`}�p�񙵰;�ͭ����%���Ih���I�>�E]T�w�w�d�0=fM�Ř���QIa	)�>Ι���F��yy����F������H�V��=�����g��gn�]ͭ�ޮИ�RQ�%j��Il	3�`z,�0$��j�*�?-�ߖ��ݺ�4Mf0� K3��y�!g�6|Uf��1��t��Ybܗ�$ZK<��~+���0:�L`oW)K���b�V�%�`l���tt���-�'(0&�;��Ŕ]!��YV���ml�3Ȗ��օ�9�B�V�b�P�����U~UN�U)�w��034֘� ��\���,v���kZO�����_��-��GL��Yb�2��z+�{l��06���Ǘ�������ǰ3#y1��"�����*�Z��y2q�L���Jl�����y�N��X�g���(��Xa����0=�%�k�=�6�1�����¸�l*`I���UU%vzsv���0=�F��ִ�3P��	kU��j�y�q�&v�]�խ06n���$��:]`*�RI����ޕ0'tf����VB$ P�IU�D�>�ｍI:w��q3�
�+��b+��I0:�L`w2�1u���V�26��7c�yN/V4�l����NM���G]�4��W&54���Łt��k*Е0:H遷:c�\<��=���.�^ԛ��En;eL\��I�02a`d���vK�z�v��X+-�=��`w:f����y�{k`u�=6p���[E�JҦJ�遽���t��F�0:�§#��q[*�l��ml���ޑ�\Y8��U�~�J������{�J˒5�.E$@����T��!)����&逈@��m�J�V���,���p�$"� V �g)�L�7���c �����d�Y�#Q4(a
b1ػ0�HB��BIb<1�3*���bF��)
���qHSD������
��N�pɒB	�1B���PO�$\`���ME �u;�@�:7���1�7P��z$X1��`N"ʐ��
d!�a����Ѭ��(��$�\E�SA	�dK��s߃��w��3Bp��&B-p��/�8�z�AdU�!$���dCD�I�	���q^�rD$����Fv�n=���������T�X
�� sU@Up+/OA ;��&.-2�AGN�%�.{Z.塼�sٻR�q� ��u��ӓ���K!��k�.�+P��V�pV�8��vˤ)c�ԫ)�K���3;i�a�'lG�� B\	S�EǱl�Y���Κ�&�Ց�N;a4i�Y�58K{vI˭�g"1���x�i�Q�ҼR'gx�]�ݱ#��3��v�@sV.%G�u������s�=�v]#��k���➡ݳٵ�Ղv<lc2�����X3��:�L�-,i��l�Ų�į��-]�K�����m·Y{m������+��UV�7n8qɞ9� hT��m&�-����|s#R���R��fٖ��`ŀN&�4n�p9gm�H!ΊU��fv�j��E�se`���5<V�7U1d��sH����Yʆ�tj�z,���*�Hl򦫭:�MP,�4�4cJ�iev�L���s��W�� �EO��]��Nf��G$�C�g<�R��E��G!��XM��d��+͹� �듷4�S9��Xc��v�b��r�Ucmİ[A<�E�g�dy�˞-p9�`�Y���B��yݝ^p�{;>��.;Nժ�g��`�B�!����[�ϫV�Cu��s��k�X���C� 	ʹӶ��0��ix�YvL���rv��(/V�۷�gvK���y푥�.��&MR�Q)(��Hum!�5okKi��=�Ւ]���y�2����n�l媕CX^���j#��Of�٫��l]��;�8pH�6v,�Jf|S;�lB�ը#͗�vyz{�ګ]lD9NCG+��U���r�j|��J��M���^�j��u+�l��1�*%<�p��,���궚@l���W r6�R�uR���44�A�5���N-����*n��^Z۶%��E��;Zq�T��t'Y��\��;T�pǉ����3б Mof�$iXE�77Scl)ق�[�z��
^R����s�x�2�S����s�(9@��:Qz���P �x+��|�%@��$��Ϣ��nB�R���r3�=�av	8*պC�/)%TWJ��:t�̬�^c=�=q�=�n�Zˌmm%�.�N�՗�FU ���-R�H惹C�.z�q�E��N�]���
;y@�n�x��LK��c
�m	r�)V�����7m�WhѸ�FVs�ʻ^x�@�2��Qzz5��ջk�Ȕ�����k6��V�1i0��Z^�=����So�l�H�r��4@#k��ND4��]�5�\^��N���b�Ù�.N��Ӑ�Z�\��c�#�\��������?3?~�Q�VB�m�l���`t�P`�&\��ٵ�~�%J�䬮�[V��,�6߳.���I�~�M��e�3��i�WY#�ѫz�zN�2�N0=3�a����8���kڛ��GQ[��݁Ǚ�`}��l��`��v=cŎ�b���<�ܹy��
K�[�-���y��Sfk;� "5
�,�;*��傲ٰ9��ly2&�"`m�1��8EܻĂ���qs���I'9���WiE�!T����LL��"��:�5wy�X+�V�!0�[�(0��ݨ�h��0X!^,1$���-������D��əT�>V!+e�װ9ܸl���g��{���;�`}�eʣuZ�
�h�Z(�!��V�>7��o;�7Nۢ��=-Fcvq��|��Oi2�+�i� ���Lw�`z�L�k\a�}|lw�6�%u�R:�N�.�7z&�:[��10;�LQͷ\q�V��`s����3υȱlȁ���2�c:�N}��`c�̕T�L�Z'm{i-?e���n��X�:����m�=	�/�-ʩ�5�`�� ��]�̝ǰ3�1�/��m�]d���J�����݃��;V�;W96!6�i��u˼qv�mlpʶ�VE]v�`fe�y3K�\�ލı,K�Ͻt��1ı/�����.L�f�4�y{g�Zd��)\��9�n%�bX�w=��n��&"X���߮�q,KĿ���3��K�f��s�z\4���&i}�$��Y5S���3�g7I��%�b{�צ�q,Kľ罌�7ı,K����7ıL��.y�K��4���,^��c���[l�s�g�Mı,K���3��Kı/�����Kı>�}��K��G�)��N�_}4��bSI�_w�8�%u�R:�M�.��i3E�b_��gI��%�b}���I��%�bw�צ�q,KĽ�3��K4���.�c���嶪���լm�;V�+��!Bɸ��$;q����t�9�xs�V\\�6�K��I��%�b}���I��%�bw�צ�q,KĽ�3��Kı/�����Kı9�wɜ���r�;kޗ&i3I�Y�<��Ȗ%�b^�ޙ�n%�bX�����n%�bX�{>��n%�bX�����U
����{���&i3I�{��n%�bX~�9�߳��%��D�N~���I��%�bw��i7ı,O��׊�%�We�ޗ&i3I�W�����Kı>�}��Kı9�w��n%�`~@!����~��n%�f�4�y{g�Zq�K)\�In��i1,K�g޺Mı,K��}�&�X�%�{�zgI��%�b^��Γq)��&i~�~i���AF["%��)���fn�pg6Gu��ӝ�\��My��p��\8�۶ �5u{nqE��k�َ�u�����nj�҂fɥ��?�|��w�R�m�78��`}�C���̈���n�ѩ��lkq2Y�(�.竷]^�o&z����z�n��\��ݜ�ɱ���K6��}�y�k�n\Z���1��݋r�kIhWo{QY`�$Bp�B,n�A�Y�c�C@�İolWc�C=�&���M�-6�*�u[-���a��&i3K���ɽ.N%�b^�ޙ�n%�bX��ﳤ�Kı>�}��Kı:w��qq����m��oK��4���'��z\ı,K�w��n%�bX�{>��n%�bX�ǻ�i7ı,Osޛ��W#��IK�.L�f�4�{=w���%�b}���I��%�bwﱤ�Kı/{�L�7ı,N��1㉸�
�l�z\4���&i}��=��X�%��{�Ɠq,KĽ�|gI��%�b^��Γq,K��=}�E��r�;kޗ&i3I�Y=�Ɠq,KĽ�|gI��%�b^��Γq,K������q,K�� ������#�V&R����K�nUC�m��E����kGX#V7/gi�Y����8��3���,KĽ���n%�bX��}�I��%�b}���C��%�b{ﱤ�Kı>��.�f\�d�L��3��Kı=�{f�p٥���mJ"���(i�'�,M{>��n%�bX��;�i7ı,K���:Mı,K�Ԟ�!-e��VYV��i3I�L����{��Kı=����n%��8������gI��%�b~���4��bX�'�;�N��S��e�׽.L�f�4�3=�&�X�%�}�{�n%�bX��}�I��%�b}���I��%�bp�O(T���m�׽.L�f�4����t��bX�	���4��bX�'�Ͻt��bX�';�z�7ı,K���~t;��h:ëɔ�%�K+�f뎝z[9�ۛs���r�'�=l��1�g�n%�bX��}�I��%�b}����n%�bX�w>��n%�b���������&i3K3�̒I�7I3qss�I��%�b^��ΓqBı,O��z�7ı,K���gI��%�bs���&�X�%��z_{��FU�Kn��i3I�L��/����Iı,K���gI��0�>X� ��l � Ѹ�����4��bX�%�}��7ı,Nz{�y���ɉ��)���&�X�(X�{�����bX�';�l�n%�bX������Kı>�}��Kı;�:]8��E������&i3K���ޗ+ı/��gI��%�b}����n%�bX�{�����bX�%8I9�g3�~>��<<��@컎ƌ��G[M m�.��sמ�""vn�v�K���퟼�l�+w��X�%�~��:Mı,K�w�Ɠq,K��=�&�X�%����4�4���&i}���I@U:�F�Ѹ�%�b}����n�$��w�)�$�s���!"�';��5���"����ۏ��$���m��oK��4�����~��n%�bX��}�I��%�bw����Kı>�;�i7ıL��=��m�P�;]��K��4����{�Mı,K���t��bX�'�ｍ&�X��>�\�'��-�p�f�4�����s�6�W�&�q,KĽ���&�X�%��;�cI��%�bw��I��%�bs����i3I�L�΅<����Q�T=lC;�������)�=����H����<�4=���P�"��%�z\4���&i};�cI��%�bw��I��%�bs����},K�����n%�f�4�x��� ܡ
���[7��I�N%��t��&�X�%����4��bX�%�=��7ı,O��{Mı��,�b{P�+����V��i3E�bs���&�X�%��s�Ɠq,K������Kı9�٤�K4���/uf�yJԪ[e��ʷ��Iı,N��4��bX�'�ｍ&�X�%��t��&�X�%����4���&i3K�OO�"�:���f��iX�%��;�cI��%�bs�=�I��%�bs���&�X�%��s�ƓqL�f�4��]E�$�?@�:�RJ�����!m 1�4M����˫�n�y6�<a^(�޾Ϗ��8����du/���95�l欣up�R��1�O[[M�:���'s;�QM�9�Qi��lvn�v��=�n��V�n�Z��i9�q�v�9\eƧ������2ܝ�`-�@�g����Of�'��	p�|nx��p"n��7]g��C"���6�ڮ��I�mc�j��Z[a������p��1F�=��'��jV:{'G�/D��#�c�������q���������&�X�%����4��bX�'q�{�>���%��{��i7Ħ�4��ߐ7�[T-N��z\4��ı;��f�q,K��9�cI��%�b}�{��n%�bX��Ol�n'�%��zP�f�����n.�`�KM&�X�%��w��i7ı,O��{Mı,K���Mı,K�︷��I�L�f��g���T�,�9��I��%�b}�{��n%�bX��Ol�n%�bX��}�I��%�bw����i3I�L��=�DR��N���s�&�X�%��t��&�X�%����4��bX�'q�{Mı,K��zoK��4���,�'+P���tA#�n۷4�9�\˗���:&�t�N�ת��7<�i�6E+Q�QڭuJ���I�L�f�{�l�n%�bX��=�i7ı,O��{Mı,K���Mı,K��z�5*�Y]�Kn��i3I�L��s�Ɠp�h�!��$ڡD˸��bsױ��Kı=�Ol�n%�bX��ﳤ�Kı9����"�GU�7,ޗ&i3I�_O{�z[�bX�'���Mı,K���t��bX�'��{Mı,K�:z�G\Nѫe���p�f�4�����-&�X�%�{��:Mı,K�罍&�X�%��=�cI��%�b}�y�9�US���z\4���&i<��t��bX�'��{Mı,K�{�Ɠq,K��;=�I��%�b{����z�S>8|�$�2V��t��uN]mu�&��mz�^�sۆ㱺��� =`�C�Γq,K��9�cI��%�b}�{��n%�bX��g�i7ı,K��]�p�f�4���X�u���K
�3��7ı,O��{Mı,K���Mı,K��t��bX�%�}�.L�f�4���r����S�2c9Ɠq,K��;=�I��%�b^w�Γq,b�	>!H0�JHX�c	� `� �HX�LF҉-]#BSA6 ��֕����rűa#!F��H�! ������\�˚&��׍8P/^c�9��D����)�`�h*�r���@EЇäz
���2 ��ar ��D8��&�#�N��ک�3��t��bX�'1�{Mı,�f�t1�S�GGj�ʭ[���+ļ�}�&�X�%�}�{:Mı,K�s�Ɠq,K��z{f�q,S4���^�e��K��m����+ľ罝&�X�%��9�cI��%�bs��٤�Kı/9�gI��)�L��S�;\�Q
��֤�:�3+Ŭ��m�6�y�Ξ�	��t��ƃ��iG��cU���a�z\4���&i};�M�pKı9�Ol�n%�bX��w��~F},K���gI��%�bpǧ���(��V�%����&i3K���M���LD�/{���n%�bX����:Mı,K�s�Ɠq,K�/w�Pq�(+]E���p�f�4�K�w��n%�bX������Kı>�=�i7ı,Ns��4��bX�ig|��o�M�`�r��p�f�4X������Kı9�{��n%�bX��Ol�n%�`hJ"`�(�(�=��&1�߳��Kı;����:�����[7��I�L�f�g}�i7ı,Ns��4��bX�%�=��7ı,N��4��bX�'�߿��v���;WR���i�N�m@&ɺ�w<ЎJ��)�:��իm�1���4��bX�'9��Mı,K��t��bX�'q�{Mı,K�罍&�X�%��I�5�S��n2b�fg&�q,Kļ罝&���"b%��w��i7ı,N㿿cI��%�bs�=�I���1��������Z�;-ޗ&i3I�^���ލı,K�罍&�X�@V�������&�X�%�{�߳��KĳK�^zog�lU�l��7��I�L�bs����Kı9�٤�Kı/�����Kı;�{��n%�bSK�a��(�v�[,�oK��4��bs�=�I��%�b_��gI��%�bw����Kı9�w��n%�bX���kC�4�ߋ���qS`�x9nA��J닮��V�΋[g��2���:%]nA�/f걍�:�V��''/CZ��X�Mx��d����lp[z�e	�P��v�h)5)�3�2�cr�V�6(�<;Y�p�=r��u���ƣX��\s��<��ډ�%��1�w�g\u�¨W;��Z��Z<��[���q�n�q�ܑ��h�y�u�M���v}����]��z�cÃ\㰖+��,���f0�7mսp2�]�7SU�(㩊A���zXi3I�LK����&�X�%��s�Ɠq,K��9�cI��%�b{�=�I��%�M,o��nXpn[�.L�f���s�Ɠq,K��9�cI��%�bs�=�I��%�b_��gI��%��/�=��+�RXXKf��i3I�V'1��Mı,K���Mı,K��{:Mı,K�罍&�X�)�Y�<r�;Pʜ��[7��I�L��1��~��n%�bX����:Mı,K�罍&�X�%��s�ƓsI�L�f�t1��dr&Y*�ʭ[��Kı/�����Kı=�{��n%�bX��;�i7ı,Ow��i\4���&i}3'����Z��U���=5Üa���q��rb3��&ׇdݎ�ay�
ʥ���d�z\4���&izwޛMı,K��}�&�X�%������U����%�{��gI��#4�����mo�"�p���oK��4�K��}�&�r��ȁ��bf%�����&�X�%�~罝&�X�%��s�Ɠq,K��O��(�v��vK7��I�L�f�����q,Kļ罝&�X�!��������7ı,N㿿cI��%�bw��Q� �GI�z\4����ZI!������7ı,N~���I��%�b{�צ�q,K��z{f�q,K4�����o��q� ��w��I�N%��s�Ɠq,K��=�M&�X�%�����&�X�%�}��:Mı��/My��nX"B�JPq��(M��B:����kPm��(0YX�x��:�=mj�����[7��I�L�f����oK��ı=ޞ٤�Kı/y�gI��%�b{����Kı9��M�B\�`��.&q���Kı>�o�i7�*G1ľ�gI��%�b~�~Ɠq,K���צ�q? �*b#4�����V�dUG-v��p�f�ľ�gI��%�b{����K�#! �$c#���		I# Fu�`F1 �HA$�
�2f&�w���i7ı,O�z�٭.L�f�4�����"r��ae�Ѹ�%�������߱��Kı9���4��bX�'����&�X�%�{��.L�f�4���~���eV��3�&�X�%����M&�X�%���}�I��%�b^s�Γq,K��;�M�p�f�4���@�r�,-u�Ug���r�p�l�X�C�8�e6��۩�ق�K۰[�"�VQD�i�7i�.L�f�4���l�n%�bX��ﳤ�Kı=���I��%�b}�k�I��%�b{��RN)�R�Q�ս.L�f�4^w�Γp���LD�?w?�]&�X�%��~���Kı=��l�n'�ZIG�&i~���-(�\-�n%�bX���߱��Kı>���Kı=ޞ٤�Kı/9�gz\4���&i}^?-L����[�&�X�~R"s���i7ı,O���I��%�b^w�Γq,Kg� D����( ��Oo^�4��L�f�4��<r����Ӷ����Kı=ޚ��n%�bX��ﳤ�Kı=�{��n%�bX�w���p�f�4���<nxl��H��l*w�8�/��v�����pbkv��>1��8���97sl�nȬvU)�/�&i3I�O=��I��%�b{����Kı>���Kı9���n%�bX��/N5�+��ݷz\4���&idｍ&�X�%��}�M&�X�%��tצ�q,Kļ�}�&�X�%����)'G�ʭ��f��i3I�L��=�M&�X�%��tצ�q,��C1����&�X�%��w��i7ıL��<yG��4;Zv��oK��4��'9�M&�X�%�y��:Mı,K�罍&�X��T���~��٤�&i3K�~���#SNV�#%7�Ȗ%�b^w�Γq,K��1�{��4�D�,K����I��%�bs����n%�bX�E�S�K"�KI!$�y��T݅�16�1��e�vyP�z��G63�����s�o��[��mN�sًbp�6�v�P��v{^f���z�o�\cʏQ��e�.�g���s֧cF�ۡM�]7-���^��ۍ�F{`p9�n;�r'=�(pr��]lE��t���vF��y��qm���5����f��/D�$܋�$��9�]ۦ����ew�"qx$�"�Kߞ��{�����'��Aɹ)��7iTy�K5qsc%�]qbh���q4i���S��!WK{���4���/����z\4X�%��}�M&�X�%��zk�A�E�D�KĽ��gI��%�bso���BFB�9lޗ&i3I�_g���?��LD�;��_��q,KĽ��gI��%�bw����K�f�������4�,���i3I�,Ns�^�Mı,K��t��bX�'q�{Mı,K��^�Mı,�f��b`�<��vEcr�����+ļ�}�&�X�%��s�Ɠq,K���צ�q,K��=5��K�&igAb�8A�K�7mޗ&h�,N��4��bX�'���4��bX�'9�M&�X�%�y��:MĳI�L�k1�ʫ,	#qCUY%�m�m���
�v�7m�v;v+{]����[N�L+�L��1n3�&�X�%��}�M&�X�%��zk�I��%�b^w�Γq,K��s�]&�X�%��O{_\[tIZv��oK��4���/��~7���m�+�13��{��7ı,O��z�7ı,O��zi7�"8���4����������2Sz\4��ı;�~ޓq,K��s�]&�X�%��}�M&�X�%���5��K�&i{�^c�V��U�%����+��s�]&�X�%��}�M&�X�%��|k�I��%��@&"w������4���.ş�~մ�����W�-ı,K�{^�Mı,K��צ�q,K��;��7ı,Nw=��n%�bX��������qn.k��99��ָ��r���xy�kkthՌ��P)�iKHԲ�4�,�4�4���&iwߍ~�Mı,K�﷤�Kı9���A� �$��=즠�	�ΖK��CE�XݪSkH�i}�r�l��bX��{��Kı>���Kı>�zi7ı,N�N��M�B�gg9��Γq,K��s�]&�X�%��=�M&�X�DVWhd�M��|k��Kı/�ﳤ��&i3K0��NX&�VZ��F�X�%��=�M&�X�%��|k�I��%�b^s�Γq,K�LD���z\4���&id??���%i�;��&�X�%��|k�I��%�a�H����>�bX�'}�~�Mı,K�{^�Mı,K���<f��8�i$ܻ�Q=�а.a�ncf���-��[j��;=tRn�Ds�g<��w�{�Kļ�}�&�X�%��羺Mı,K��4��bX�'��M&♤�&igqy�9-n9b�8[�.	bX�';���7ı,Os���n%�bX�wƽ4��bX�%�;��6i~Ij=(i3K�g��WKH�Z(�n�q,K���k��n%�bX�wƽ4��bX�%�;��7ı,Nw9�.L�f�4��<r�[+���n34��bX�'��M&�X�%�}��:Mı,K��}t��bX�G���5��~�Mı,K�O�p�cV7j�ޗ&i3I�O��]&�X�%��羺Mı,K��4��bX�'��M&�X�%�O����4��93ٽg�Ws�6�;�1֓[���x�u�H������[ce�Gi�T�ZMı,K��}t��bX�'��zi7ı,O��^��*O�b%�b_����7ı,Oz~�`�ݐ���3�����n%�bX��u��Kı>�zi7ı,K�{��n%�bX��{��Kı9���zK��Ɍf�9%�f�q,K��ޚ��n%�bX��ﳤ�Kı9���I��#4�����oK��4���,���m����sffs�L�Mı,K���t��bX�'�Ͻt��bX�'��zi7ı,Nsޛ4��bX�'ݝ=��cy��X�8[�.L�f�4������i8�%��w^�Mı,K���Mı,K���t��bX�'��$U�&ýV	il�J�D32o�$��(��HY�$`Mk&B1Dv�h��'�H� B ���@�6�E�ӄ�c���2Q�hV�	a-�!iH�&&%G�d2�j���r��(�k�����.
BՁ�T"�! �O�Y0b�,+b�͒]	� Ҙ&�x��ЮpK�ȁ�HLB0�%���H�Ȕ�HM`,14[�o}�q�T�[j���qU@Up*ݲ���[�S-ۡ�����ɻ6{:非���c<l���$�X�nP�ړ@F��Q]
�؞��Y�K�5T���K���%r�*����,����R�]mF����v�>�v��D�!�Ya��jnp�}��M��b�b%O����z����G�ZR���M�εn�nǛr���F�yѸ@��� n��=��������ɍAu����r�n]�ɭ��z�n.�*���g<��^�\	õ*[�`x�L�q`ہ�Ut��gaxu/0�4v�w��S�O;�(/kn��.'�l�UJgc���p-�-�f��ۇ6A��Z	Z �+T�:�WJ��ⴼ�iVⲕ)AR�ZV��H� "#j�n�PmũV/�%۳-��@D��"ݕ��:��UR��+'���Sٖ�.Ѱ��5�) -��` )�s֑�nȢ�n�#,�6�z��� ��h� �G�4�����U�ú�Rಬ��d�x.��
�9K�!uÞn��6��f��ZԶ�a3 �R�#�UJ����kB����*�:j	ofˈ�k�o��m+Lq�ϝ������]��\��}gk���y�Td0���l`���l��.��$F4�[ps�vgmΰ��d;a��
V6�A�v6:�Ԯ���A�8D�o��&8:�j5�c�s8�����0=q�:䴽`�P�v��OF�X�J�[`x��g�z��*��A��[h��ot�ԵÄ�R:���#���◔�����B�$�T�ۺ��gUNvTy2�];ۥ���H���Gl��n���W�m۵<(R �"̀�#�t��F��:���V��ۛ��
����'kvB횉l|�]�>tZ��f�:�A�����&U���5ٵN�b%AN�WH,��z�_4NR��|u�	6	y+cḈ�ջ<��N�=���C���S9��b��Uj0���[��s����մ�ztJ��$(�ڈu����!*q=phڈ�_
Z�l�N �U
� �d�Z�4��J��Ϣ�%vƥQ�,Wpu����T�ȯ2Wn���,��n3R�N��˴;�;�榥���kM;��&m�`�NB^���������������|G�\������˨G�c����	G���8m)�2��v�v|k���[��tl`l��ۣ�Pٺ�v�D.oS�Vgg�9�L�Z�n�\G&�t�@닍�tv;[:�[%�7i��{�����`��\�TWc2:������ۏZ<������4=���7]��Y������Kı;���4��bX�'9��4��bX�%�;��7ı,Ns>��n%�bX����1��W)��M�p�f�4���/o���%�bX��ﳤ�Kı;���I��%�b{�צ�q?�b�"X��<X=���E�XȬ���i3I�L����I��%�bw�צ�q,C1�k��n%�bX���k��n%�bX��=���j��2���K��4���.���Kı=���I��%�bsǵ��Kı/��gI��%�bs��4���\���i3I�L��;�M&�X�%��zk�I��%�b_s�Γq,K��}�M&�X�%�����5bV[SPM8=W.�����r�t���r�LuC!:9|�s��U��&�\�9�Mı,K�=�M&�X�%�}��:Mı,K�Ͻt��bX�'��zi7ı,N���e�p\�ˌ������n%�bX��ﳤ�0�Ԋ	 0b����O(i�MD�1���t��bX�'���M&�X�%��צ�q?.*b%��O�I9]�X�8[�.L�f�4�����n%�bX��u��Kı9����n%�bX��ﳤ�Kı=���
�2�9^��i3I�L��ٿM&�X�%���צ�q,KĽ�}�&�X��P���k���K�3K��ߎRH펑9a+�ޗ&i1,Nwƽ4��bX�%�;��7ı,Nw>��n%�bX�{���n%�M&iw����7	H5�@1֚�N��Ί����N^������UWN��H�q��(��řɌ�&�X�%�{��:Mı,K���4��bX�'��4�},K��k��n%�bX���W�@�Dv�ݖ�K��4���.��I�~ 8���';�_��q,K���4��bX�%�{��7ı���~�jۡ[U���7��I�Lұ>���Kı9�Mzi7��! ��4�15����&�X�%���k��n%�bX�������ŷ��e���n%�bX����4��bX�%�{��7ı,Nw���n%�bX�w���n%�bX����9�s�.1�s3��3I��%�b^w�Γq,K��}�M&�X�%��}�M&�X�#4����ޗ&i3I�_fm�@��L0�g�w=���ύm+\��g�;�u�n:��������E%G�&����~����%���^�Mı,K��^�Mı,K�=�M&�X�%�y��:Mı��/E��
�2�IM�p�f������&�X�%��zk�I��%�b_��gI��%�bs�צ�q,�f�4������A�;V��i8�%��zk�I��%�b_��gI��%�bs�צ�q,K�����&�3I�L���oҵNƬd����%�bX��w��n%�bX����Kı>�}�I��%�Pl@p � �8��z}��Kı;���F*�,+��mޗ&i3I�]�}��Kı>�}�I��%�bsޚ��n%�bX��w��n%�bX��<8����"p�I	(�u�Qd��6v�,��:{(>	�Y��o6Z+�j,t�c9��3t��bX�'��i7ı�������]��fc�O��-��+N�IV������&�����z��ގ�Eq��*_eb�X����\��jUT�ߤ֘b���#�n�+���%��;�`s�ͭ���l>�&�Ƴ��[S,���x�0=�:`t�P`m�L`uΘ�Ե��$��{cz���V��F�w��D�n�����r�d��Fj�N,QOY����Ժ�ڞ��� ��n�ZiX`���Hj�BP�`�=�'��#cH��N�:�0��8H��<q��:��k�i7[d˶98�[!��9�s٭�:���,&��
��xX��	�#1�M�[�d�4I;S�]�ք��ק��zZws�fq�Hs���f�nV�Sn�~�������旨ʝ�qey�(ط6㎴�bq㎼�y�ԍe;3���֭��PN�Ie]ߺ��`|�ܛ�;�`s��[�:�\�u��Ռ�Jl^d��RUvKټ`zn���C�z�Vϱeoʎ�8�+�vY�1�=6;#�l}��F�Ie],T�%v�0=�:`t�P`m�La����O'��`u?~���ە�i�`t�P`m�L`uΘ��tt�ڒ��Gc�y��X�����g�b۷GJ>�ގ�'2�:oXn&��r��-Tݓ�'��c ��0=�0:u(0���!]vW
8�,�s�w�(��Z�y<�өA�����8��+VR���1$��tt�킃?}��U�ܟ��O��`M�00-"����2ҦmE��c ��0=�0=�U�x�F:Ec%%6{�`y-k'�Ӏl��0;`��띓*�QiP��R���z�r)��8�nv\��	4nG��{Ip����u�ZY+�yܛ��:`v�r���lӥe�^R.�*X��K�\��:[�t́�xc��l����V��v��|�;u>61�  
1!�(�B!��*BB+ �T�T�*WJ�Tܿ���#L�wn�m.�����vw������sk`w;L{ ��q�㲸Qŗ��s�0=�0:r%�=���O_<X��u�ъ'ZUƥ��f��^ø�7N�6㋛9�X�s`Rt���\�x�0=�0:r%�=���W�UW�1�=6�������;V��v����l����<�t#)e�`���Ζ��1����`w��3L�Gb,��W���*���lI�03ӷ-���B�U"�@yEM��߷u$�g<`�5&2]f*���ŌwGLخ[ݝ-�fw.�����U%�-�tU� ��ل����9�uh6�n���=��nl�j����G%\��y�vw�$���K��J�h��=�������ND�������8;+���6�g�����'"[�zc\���*�3ēӣ���l��?W�}�&�����=�)S��N�H�[ND�^��'D����+J�}YX���n�ș)(Y��<;5N��	�VnW��f���͡3a,sb�RV�5��]�F5�ɡ�2��wS�h���\
��HK�&q��[�2;[@j��z|�=A��@�$J%.�3�w��}���2'G�P��1RN�3�ٰ]����'<��sۇ�v�7F�mm�6��j&N���1]���4��,�y��sPH�E+�
��+VV�}ִ���o��V��G맱Ъ���wnIiX���� �磴�t�g�i�[���_8�8��,Ŗ�.~��N�����lW��Y#n�Ym�Y��r�gGLخ[�zc�zUძ,���J�0=::`v�r�{�s��'�;U��٧i$�`w����N0�:���������wޮ���iR�����׽1�t��0;bx�ז\����;(&ک��f�ƶ̸\�ܽ���Dr;��5=Ɩ4ڱ�v�"�0E�]�� �?b��nh�>��{֚��"��[v3��UU/$�����H�Il�d� ��]�ω���j���ڶs��`u�L`:&�GLwY`�]��WYK,Kl���D���釴�{6y��`{K�1؋m�K6�'XK�7�������N0�/$G]�3�w]d-f���&r��GhcN�æ�ҹ:4Xs;f
�v):$���0=::`IȖ��ޙ�����`rxy�ڭTv�;I%[3�ǰ:��c ��`ztt��E>.��X�IR�s�m���`d�=�iUP~U�T����x$�,�J�rȓi]b�aH��O�����Bg$��MjPv@CP�ee�����4J2F,d>QHp8<�<QO���2ZT4e�����XP�k�	�#�d���t��ЁS�XF
F	!6?\��e�S))M�v�	��\0���  VRD#�!:a�- �`"@����.����og����p
h�!XX0>r�+H#����`�?#0��	���i�jl�B#1��B&��A2�����&PY�*ł �HC������|�B+��A"d"��_�#�1h�_T0B �4�У4\'ʡ�Y||��6�-��6ET�V�ɚ8�P�>.�"��� 	2�oTw�}�ٳ��i�'@~u�� 
�?�+W��D�#H$�0��@M��ص�ʓ���g/��L	3�����V��/2�0	:&�GL	9�=��y;���=�:ZF��K+I0=::`IȖ��ޘ�$�ǵcqւĭ��"������s�7+���ӟ+�[[�\Vw/$�d
s�=�]��;2Ҧ��l��N���_W�7�������U�
�Պ+l+�w# ��`ztt���-��n��yY��I%���ӣ���l��0:����BW���b$��ti�&t��?fN�j�*B�*� ���R��8:׽�gRN��gnn%��դfb���l��0	:&;���Z֟�"F�V�G���Y���,�Bjي}x�pW<q��Ml1���r��N�]%�|��k/-_�6OɀI�0=ݛ^K�=�W���8&�u2��`d��J�%v{f������ �w.�Ǚ2F�-VE%��[v3���;b�l��`:&������b�N�H�[<������ �w.��fmlw���)PՊR��`�:�2d����L�-��I(�]�K16^]7`2���[42�;����Ŝ
��û����&���Y5��3]�lr�Kp�y㽜�.3��y��YLhk�I	4BA�����V�Rɹ=jE�7e^6��ڸ��>: ۳��]s��l/�6�r�v��:��oj�\��Gq^1dV�5�kxqWuaW^���
�MS��u �W�+�����;&�b�������F ��n�뻻���_�_���&{}�Z��x-Od��ެ`Ѡ�ѯ=8��ڴu������H��f�� 7﷬�F�3���K��$ް1w/���;-r݁�������;�����{��gز�'c%��WV�����G�`��t��3k`s2�V�7umU�B��w����:[�GL	9�BL�2�1U��A��L�lwGL	9�>�]���0���Q7�Zޚ�UerW���ۮ�clz����W�:ioMY�c3��V%�/1+`{z:`IȖ�=�L�liȻȰ̤*-$fZT����С�#  �	�Y�ֳ�3'q�ff���ty*i؝ %����cL�lwGL	9���J�],E^%K�L	3��=$t��#��06�)F^%`����V,V����d��D���1��i/b���4�FV�"�9g&����O����\𻗄�:(mٱ�ۧq��c���/�#3x�����0;�K`{�t��E(*ҥwy�T�����0;�K`{�t��#Г(�J��G%����`s��[&�׵�@��
��T(����jMI'>糰:��X�]��[�;^��s6��0ݒ[�"2+-�夎հ>�͆�������^�z���f�����7\n�S��Vh���F5cm�������汍onl=6:��x����!`��V#��0$P`{�t��F�p%TR_f%K�0$�t��H��ot_��a�ߗ�r���S�%���=������D��(0=0�]+�B�����u0$�� �d�I�0�J��z	  |�P�'^K��jI���5K%dԥ����{ܻ�g���	��02N�05*Y��o�}�1�d��4v^�V���c����y��㶶o֜ێ���
vs�.s�+_����{�=#L��J��6oXf�r�BH�-n�e6~���̸��L��I�=�UIU]�[�|����h��l�����r��o=��`{�����qVJ�mV� ;*6֝����	�`d��`yx嘪)/���Ę"�l��"�`2u��Y@.�ZX�@�Ye���a�����9��5�i�/Sc����m�0\�se�<������7��v�;f�e���H�*���W>��J��d�aW���ӱtf���i7�{^Mz��1�2��zJ���m��ݍ�vƃ��S��mгb�ft.�vJTNݣ7l�&�q����ܶ�6�u�v��W z��Ġm�BcY7n���v&U�ŭ�^�Iif��\I%�q�\T%f�<	+��tg��cfؓ>����}��Y��$�q;*�Q����� ����H�wD����r�Ax�Z_ZWy��"�0	��P`M��t�r�ϖ+�I%���;�`t�	�:`t�P�7��Ta�b�Vah�Ę"�l��"�l;ܻ3�-�,M�cr�)�'�i��v!�L��I�0>���}߇Iz����j3m]�^ �/mm	��b��6�Vek)�&ji�܎�d]�f��?~_�`:&H�����(0���F�T0�}���*�RT�J��T�cs�`L��3.#`|��Ԧ7!Z��er݁�˃�GL�JΉ��r��*̱���$0;dt����l�̸lvu�D��ۧkrU�;�J�dt��%�YX����=Cn�P3;�z��87F:=.������pS�Yb��N7&h��ft�HN��A�6GL�J�ܔ�̼�j���y�0;��l��%�l;ܻ3�e��D걹m�`M��dR�g���߾H��`v���,x'��*%A\�`}�q ��0;��l���@)����b0���`�&�A�6GL	2�6�ִ�w=u9%u�e�j(k�ۋ�{]����n×���@y8��؋���)[qV��2Kx�=�3�ͭ�����r���b�T�(��+�l	�:`l�P�6tL�&0=��r��x�$����0:E(`:&_I��0%l�Q��t��1bC ����'�4��&֨�cH�p�`]�~�5 �7�Eq��S�:9-�y�6}#L��fN�6�S���l/�wn,nMn��-t��N������|�p���r�: m�hgi����?�����Z`d��`2wi~����`zŷ�y��e%\�`w2�7��{3�`c��6}���6}�@_Wc�E% �C �7����	�`zN�0<���)���RE%����`gٛ[dR�;�`v��e�v��Uk0�;l	�`=I%��� �y�=�g.���U_���*��U_� �*�EQU�B*���TU�"����UW��"1�
��
��"�",�"Ċ"�`��X"," ,H� ���H���*����U_򂨪�QU�*���EW� �*��QU�*���TUw��U_�EQU�������e5���۰X��� �s2}p9| �UP�H(��R�$P� 
JJ QB� �)J �tJ $@R�UPH (H( RT�*B� )R�����A*�*AE
�
��@�   !� H*T ��Nh͚ ��CO� �w0t	� q�e���m*c��\YK} �[|�S���  >�]��z��x zW����,�-\��yo3�K��)ޤ����ד=�qeu��W� ��  @  
���b�}�^�������S�qjU� k{����jr˓\�����\ jU��wU��� 	��J���]�@{�}���ȱ�7f%��l (ͳL^�{��{��۬���K�}�@ 
  P��S�Je�`ru֜���һ� w:\vuF�zy4t��� 8c����  ]94t�:\p :{��@��=�:��I� a�9:�rk�n���' =�   }�   
�P����ŝ�kɥX�Ը 	ҙw{�<Yu��,*��w }���'ݞ�C�i����z�� ;�7��zy|����ݫݞL�� 3��6�i˗���K8��� � >�� �C@)Ͼˋ}���渲�n}� )�A�1( D 
$R�Se�AGaT:\)JD    � D41�;2�R�  �Jt D��:)4G"����i@ D�AM��� =A3T�Q�F@hD��T�@  Ob�H����F#CS�BS=J�� ��	�R�P@x�%	����V�%�s�e����N��qݾ_� Up�U*��U����@X�������-<z��5o��Yƌ��7��n�\��#H%L)��Y#��eg&q��F�6`&07$ْ���"��c##,�@��A���:�Le�8m��r��9��$�Ν�;�� `�P���R�ő��!m��RYq�\���[���Z�ũ1&e �B�1$�,	$2|�&�cq1�Z(b��p@!��&[#*Ro��a~�a%�XSM.�[�4V^g�D���TR�B�`!$�ī$a����I���$�;3!��@�t�7�C�Wp�֧ K�D��x���`�B���M�E*�~��%��0�|��3V��0�ۂ\u��:H�&���B$�%Z�I��$
,��R7�K�[���������@!�!`}�����5��
T#����CK3�@�\��Ԫy����/�Za}ըH@EUO*	3����9wgs���G�0"S	%TÍ\'��ֺZ���2���p������{1��ټ6?! $(��=W��u�Պ�.�dҼՐ�!)[#D0g|$�I$���ͼO����s�S��K`�H��9�LcaXх!q�B�FÐ�!�)��W+$�����â\9HS,� P����C�B�B���cX�-:c\i�IXSpLa�h�r�.rkR�RB��)M���WyyOe�e4��^� ��
Ē��#�H��D�uۢMh�Y�ri>H3�٧#�.M$�8�Uţ� �M("%	^\*��
E�śW���'���$�E./vY��Ḡn2h��\b6��˲��Ɍ9��T�V�  W
A��`V�%ń��lb�	*K##VB,+	��0�3�����/X�B�i�R9/䈚W!c��W���M�բn�L�LX�n����:����綽I��: �dM��k�΍��
`ri$��0�
��M��H)�I�sf��q�B	%
��R@�BH��B�H�R,�BD�9�R4�D������&{��yr&E�Bb�!�HBe]ȱ�HU��1�$\P����O���H�*ĩ�G�!36}�paLc����\{VyZ�S��ϥfeν^ܑfԕ�|zH�� �%�V��K�$&�¸8CD�ً�`Y�H�J���~3�+����CDF߶����^lꊄ(�	��ʠqt�ĩ
%kH� S��3)��Q�jHjReٍ�� �)7�!XA�@�Չ"�B"EL�c��XWɂB�`,0A,(����9�#*ʩ���K�o��?1ML]_�O��;pߝ������n�v���B%R�a���j�bi
�r˽TB��:�d�,	.Ͱ�	Y��\c9�
u�m.�2	T@��#�H`�H�"1bȌH�\C,)0���dnȌ�&�a�MM(G��f�"����j\d���	o��S�l�3�l���U#���	 T�L���$"��-��,HaW���`4��\d"�I�sٸ;��s @��TxM9�B!,7,�Uj�J"D!��3J���m��]��4���唳Ե-�)@�(DHs���@�(��3�֎�ԋ ��(bF02�X\p�%�M.u!&��AU^A4�d!Mf"��RAx�U�$�?>jj���r*�۽)���*i<��y��Sӝ��%uW����N���łRE�`�UZY1�""�_�:J�[���ʻ<���s�Y�Om櫲k=�Ƌ�>��t"Xr\nS:6�JH��c�s���k��8;tV5���NP����0��}�McN�%��E��L�9Ï	C�3���oג��)�7��o�M�Z�%( %_�bR@D��^]��{_o5�c�Ŝ,zH�HP%)���~�i���M�H�1��,���\Cz��Hd�Ӳ��cH�#���Ѷ-�6��Z�	C#�Y�O{ZҔ��J%R���Nz�E��Q(R
%����^H��-�&4�0HVt������\���y�s�i�n�ez����*R��UW�U/����{�}�w:�3��iX�H�#C+�%����H���X�F+�BB^Sg0���;3��B���Ĭ9�"��d �E`��g�N��w�Ϛohi�D�eS�#�4�B"S
dݐ�Lo<��d �3�d+�m	]�Ԧ3��q��"6T���
ʡ.+)p�cXV�̼Ƥ�[#H���)�pF�)$�9�Ne�U�v$	-���^����k?Ip0e"0� \ ���*@�LL`%%H�%���kZι��tL����`˜�m2�$�)��}�0b��cB���D�d�`4��"�!}��0�7NHb���S!�sÌ��_O�od���_T�k#9�y5r�f3���i���LHp����`|CB7:F�}5L��]�}h��n�!�Z��pMuY^�u�Q+[DƤ�i��&��Ҩ �����\k���$au�$0�k�ci��)w�"	�K�Ys�}��K��E�S�E���ot.%�nn7��Q�w� �1�|d����6���A��2�}���D����7�d�.���,JV)�j��YY� �#ʵ�*�VT��1K�$�!p�)���)�7!�e��d��LfB�������>�B
BD�H�F�����[��>�7\.X�D �$*#pʒ�(��s$�\�)߰FI+�!H�!B@��9gPķ��Ʉ�!�P��5���w��ɤ�
�����/7n�k�;�w�Lg� ����>�Z���S-������j��2U�[���Ă�ˡ~�|}���T�#Yt�������{6g'��$�0�������y� B!�	�b�W�8��J�h�
kע�Qx��!���s�\bCW43.�L8�0�L1��C�p
< Ap���.5����NC����0�`�!��!��(]�8�~���
rdE��gU�7^'2�/����-�e�.�]��6�5x���N�0�P������'vn0a ��,>�%��;�7jc0DJ.q$2C�B��H,HD��!B@�H CI)�L���SG�+�C;��c��aX ���8�BB,F!�H�q6B0���'pF.ܴ#1�X)���e�$���B��fh`�+	
`��v}ܒ�H6D�F$H��Τaq�%Ŕ�����A�m�r\|��e�@� ab0R��%q�*S1��36����4jT�Ml"�p�Τ8B��(Dq��}��vCfZ`�ĸɐ�GD.l��1���k�1��Ie�BW�5���f15���'1�l��������L�5󸤸ΉW4Isu��&�\�ΆP5��$I.̬�*ܽ�"�$@�)gk�5�	%� $C�c$�BX �"B�"1K$JF D �XH�@�b �`!@�I�
� �
� ;�"�C#��������^o�$:0!�f�{۲ٸ\o��F��jp�R�(��2�c9����Z��4`�0�h�k
��!�&,@�GPb�k,%y �U	-QIqB�I��q�E�l� Zm�1��X�$�0*aγ�����Bnϔ��'���䐑������"@�X�!T/�n�a.3�\:4k�8�3Z6�Ӓ�#i ζ�옵
v֚"/r�AS� ��J�~8�Ԑ�5��0�<��>��`���%M�q��@��0He4�58o&]�l���(@,i����+��D��ϯX��,xnH!�!L9�P��ʌk�p�~�S��FP���!R�Mnr09(� qL�@�0B)H�9�7�� l�,d��ӄhaɳalֱ��X�ٜp�1�8HP�@�3������
a�@�6$.5�N��2I$l-��p0�v��P�9{�3מ�g [�B�Pm�,7-K�)iH����E�V��f��{4D � )�J�A51��M�$��hhcC	�#\M0�)�	L�#1gP�HF�:R�DJ`3����	��P�C���S(@��
`a4pZ�V���d[,@�a��2m���*B��>�o9�B@   �6�ڑ�� p ^�    ��sm����l �VGI@�5�{s�Mc���f��h�� ��ס�6�eB�[���j�*��m� �a��m��[[lp,5�� N � �a��,��� mpڮ������ҝ6Z8.k�6ܗJ��:�K8����H[׭$aA�`�-.������H ��YI.���H$pKu�Ih2 ���]���{l���.� ���`   	6�$8 ��~�| �����hkXp~�� � ۶�h`Z� �Y@ �m�i�����m�@�    �[�:i��-� �b@    5� � �$�Mo\��b�����N�vä��ҬU[�cP�U[B@� �� m�kh�l ��R�-� 8 �%�   [@l  S�3�4[�����Ƭ��a^���R@�����m�RpJsC�z�m���k�@ $�Ep[���J�pR��z��8h:қ�g���:�.���`Ӛ���u���;���Zn-A�En;6�Pv�燃�;��۴/[���0���+u`q��m�ڊ�tb�B�����u�%�v^T�>/��|BzW)�q�1bE2�C�UҙP�Ҽ���ť�y��,1ɶ/$`�$-���ζi���H��@��z�hzV�&�2��p,j���mV��i��RH ��絲2�*���8�!l �UTm����8Xnt��r� 2[G�Ă��Z��(j���UZT�tˮ��nݩh 	 �km��6��)A��FQVb��r�Pv���I6ؐ��-�X�����^zU(ر��f� �`� ���J�U\�n��ƶ���ۚ�m�GPS`��@���j�mjJ�m����� ��ml� �`�7���m��Px���:�`
P m	�  ;Y+�m@@]UQ�K�,�T�v*�.j��Wi%�X� H �i� m�� ��[w�vT۰ �l����2Lm�   V�a��a [[l"A  m�   $��-�  l*B�����j�`��    ʹ�u�e���I��v�n��  -� m�@ p ��m�   �m֛`	�����j������c p 8�)@ ��w��VŴ[E��l  ���6�� 	l ���	��ҥZ�� �[T�e�*�We�iWh��t��U|W��  6C Y[l�6 I�ʽUm6�   ��ɸ.�   $[N[��d5�8 R�ԫUJ����4�/0a�I�  ���p  �;l9&� Ӣ�~K>���m��-p
�9�v���P���$8:��\�t��Z���KI���T� 
�j[u�nܻ�ԪR�vok���m'%�/hCsCUl��6&�Sn�uul�.K-k����S�r�ة�V��n�A��xn�ʫmU�;����ª����(5��we��ư�ms�q�M�%���C`�JeQ9��Z�V�c��|��~k�p
��a�3��2�K�;A �䦰���k��]�Ԫ��:J�T8r�aU�km�ꪫk����󲴚V���| [��M��'E� �p��nݛt��-��(jk�2�A�lI �`�	6ۆ�^����M  ���L�r����WP�z�؇�i0���R[ƙ��X��&�Z�]��uכ_#�+��Q�n�˰9���֍��k��鶍�N�2N��,��+��3��֦��-�j���l�-�a"JID��m�+ 5*��<�V� ���	V�h8�	V�����0��-�z�NUiJM���-ۆ�V�Gl���+Etl������	x4= E ѹ����W-r�v4�UF�7c[	x7\-ic��ݮP� �E�h-����[m����S��Wj]��%���z�ժ�]]*��m�yZ��:y��k�B'n�:Z�M�et��&1v԰WV^����H�`t�$�l� zG��#�� �8p�\� �I�@   ��t�	 ��` -3h��$�m� Y��9U*�U<� �*�uE� ��������m� d�n  m�mp  8ֱ� 6�� �VM�۶� q��l 6� 6� �   *�V�BU��*�UJ�@UP����U]*�n�H��v]�8-�   l(� uʹ�V�!�8H)c^��l�� ��m� U���-��V]��UNu�Hllm��i��Z��݃m���p��e�+�NIvٶ�� ,R��Z��h(MT�5V���  �R���\9k�G=J�i*�c	5��9���s��&8�K�2%��������Wvv.�v��/A��n��Ym�8���uvʠn���`e)Î�	�A]� mջ��7nZC#�nwFU3uR��p!A)�"�@U*�媀S!�O<�lQ@Xl5R�U��]mU�
ʩ��<�hmm6Zlk[m�Tt��E�1e�T��6��=eej��X��9�Ks)tP  �)@�6�Am[G��[���l  ���������,�{6۶�l���|:@E�m�t��m�[SJΖ]44�� 8m�����=6�,jj��V�&��l�   H� [vͤ�6�*���A���T��U��,�!�-�m� V�a�l ��V�����ϊ�ԫ@J��$��V��U@ �` 'Za��섁�h�m"@km�$�NZf�˦�p���� ="E�^�+��ڠ*�CaZ�]���� ��mK��8Ȳm"��$H�kn��v]��U�djt*ԋmN�UT����ڪ��P	;Kd��%k����  � 8���-�mt�,�� m���m�[���	��  �{(Nyf^\ax�[0
���J6�M�[�6i��,���랪��>@	 ��m4�u���`A�VҭP [��5�T�FE����$L�UV1Uob�Tsngg�[nzvݓ7n�F�y�o��q�ӷ��V��؎s�I������큷kd�5�:��)m��`��U+ѐ���P�6��5J�����fY]��^Y�͵�9�	����� ����Vu��ق`+k�p�ҒҭE�������  8�[^�L��mH\�	�    8lm�� �9�t�.�  lf  u��3��5�Y]�YT	Z�V�J�@UR����C �[t�݀i2�ʥ�]*��Z�X���h �����cm��Q�m�� ��    @�oI �c� ˑ}֪�U��y�:yUUu*��du�U��k����G�Olm�T��,MʪӾ|��|��8�󎇖�,e1�4ܣUUR���,D�Nw@n�m�B� ���*�a8HklhMQm�}���f�s&յ�	��ݴ��mU*�UH �O*�T�չ�a۶�t��od�@��k�^@٪�<ʽ�U�z9��P�8e����	ǹ��8��Z��v�r5�;<���5T�]�	�P�]�I���-�'$���G$6���U �9���U^�K3Ӝm���v�wKX�qo/EN ����G(Aq�9�W8���UV�nˍ�;XQɸ�e�
������l5Vѣt�VR\�.�%Yyl;�vr���ۥH�[KUT [@�!zKe��Y�F@�C�kd9���Ғ�[P�YY����V�fb�S&�@UUU*	n�lY.�kQ� �j���:a���ǌi�L�mgi<uR�<�<첼�Q��J:;]��p���U�y�^[���m�r�Zm�N��Kd!�ȹx�K���U��~�     p��.�ѫb�C�
���j��PO+mǌm�쌇J@��xr�/,ksv\sY{j����ʻ�8��8�3q�m�yWnݣj�Wll���ٷ-�C��M�����Ms�V.֙�z�%����3�]�Y3ٰ�t)ᤗe��R5��oM� BI�ZXl������8�Te�U%�Ò6ͭ�m���i&� �͛n�h�n�%ĉ�J5��*M�l���L�ͪ���nʄ  �� ��d�ᨢꭞF�I.�l[M,m� m6�  p  p�mm�7]�-�> ����K-2��l�*� �M�I��&l܆ Hp>��r� � %T�M�V�<DԫPګf�   Hm�  8�H:EY#����� ���  ��h��[��)���L�U�(	-���vŴ �[�$�8����rSG]�Bje��m����Im-��H � ���   ٶ n����C3mm r���` I t 	�     ��Qm�g     '��mm������&��<-����K�vP�����{��*�:G���� TV ���� ���$E0@G�� 0�� '¨|�X��DT�Ɍ(�TàLТ�Q8���Ps�T�Tɴȿ"wv"��Q>C dRH"1��b+��1:}4�M���=!�����Ad�GB��4��@: ��g��t�G@�����aE���NA] V#�V 0"�D��:�P: ߔ�V��O�48�>� 9b����.L�j��EL� �'�xh� P~��
 ���: #���<��髤AڛUR~m�"��PeT+W��
��N"$`.ׂ�D��"��"����
(��M�gB�#� 'A"�`3�~Qp
��Q�QW�X�L�T6�t�\(B
A�TL�"	A���u@� :@��� P'��P؊|��@���	]��F�Q��Ӏ%[@�
� &C���D ���h 
��(��F	 
T
���`�������� E��!�������S���#�+�v��N��52:�ԸW@��٧���8Kg�s�acd�8��c��j�j�md3li���9J�r� +��ּ��U�Ňj� y�AUU�ݖ0`��n�[@�h��\��:��nbcv�;R��l\Wn�Mc{X��h;f�6�o�i��dݶ�#ι�vݴ��+1F}=��L���e@�N$��t�@l���,[ROciO�vWH��}e
���iL�:����n�jW(��Ue�Q [���J��l� ���)`:�ԧ5�P3W4;#�iY�@sR�C�ۥrX�*KhD�$��m�6��e��]qn�9��)�#�Cl�)�;X�8���͝�e���m�#�ƌ쫱�iN���Z�z��,Z��0�8����)�O-뭺����'f�r;R��u����6y2�
u���d{/��`�v�Oul�u�6j:�nu�nke�9�.�.�N�[R�	�ݪs�ӕYsv��)t��P-��1�Hf�6�h$ڲBi�f���:����Xع��K���e�n���"G�vN����Y[�\�=0���Rgc�� <N�.����YA,�B&�jt=9C��#�;ʰv�6�P�]j:v�QȬr�n6��=��P�;��p��R��lx�X��=�����VH�O+g�vWiU�8M��I2H�ޗ�Ų^г�#��zܹ�]�-�i+�X���%Uԅ��dYD�*lF�	Itfѩ�
�KM��C\9keZ�]Oj4I۞G��5J'��nz�5�Ѭ���OY�tE�t��.ِ�8�s����m�.��ո9{Bm�R�]h۰stmƨ|B��������S;+q�(c������`�c7����G4lΚy˰lv�v���Лq��g��鵲����	Et����(����:��r�Zu@�� �ce#�k��V��`W�{tgN�!�1���;4D��KR�ڱ,�@C�J��\ff����Rc�E�&W���G� �_� o��8b���!Pt  lh�~�O��rA�tp[����Nd�@ n����2h�[�g'Ki ��t��&ɴWI�^B	�lmv��U�l1�&�k���*j9zY7E�M!�\��n8�{GS+��]��-m��"��&F�ɞN7�-��qU��;������񖧃�^:�#ל�o\��v��N�[mʃ1e����
�Dє6��X�a��b�3q���.҆��n�ň�\q�
��ϳ��=��Gʎ{n�m�۞�Nɸ�ϗ&%�V^ZK	�L� ��o\,�H'9�r����LD�,O��oI��%�bzt,ɉ�d��1.1���Kı>����n�&"X��q�SQ,K�������bX�'{s�SQRB�����pZ�*�f�U��ِ�AbX�'{�v��Kı7�{�&�X�%����T�Kı>����n!�����{�o�,�*^2����X�%�����7ı,Nv粦�X�%����f�q,K��s�ښ�HRB����*��*�]������bX���eMD�,K﹮�&�X�%��w�MD�,Kw��n%�bX�^wRz�Ffm�ĸ��b����W���N�4�N�v��]J��5z9wTa�E��H����&�Ʌ����$.���bX�';�v��Kı7�{�&�X�%�َ��5ı,M�<��e�N;JB6�����{��7����	�h�$Rd�BE'@���E�bA�A��ќB?D�K}��4��bX�'&;ۄ�Kı>����n%�bX�N����12\&sfnsjj%�bX���٤�Kı;1��&�X�����u��Kı=��֦�X�%��g�&c��9�L�d�n%�bX���nQ,K���k�I��%�bw��mMD�,>���Kı=:d��e���f�5ı,O��4��bX�'{�v��Kı7�{�I��%�bvc��MD�,K�
�~���gjr������L�u�U�n����y���E�#�I�Z,P��Ͱ\���f��%�b{ǱSQ,K�����&�X�%�َv�5ı,M��d/��$)!u&����TUT�IX�1�T�Kı7�{�I��%�bvc��MD�,K﹮�&�X�%������*�TB���*�]US2Uɜٜ�&�q,K���}p��bX�'�s]�MıT�dK�R�X��)�U Z�F�,LD�9�⦢X�%��;ݚMı,C{����^�7=�\�-����o'�s]�Mı,K��;���bX�&��vi7ı,N�s�	��%�#�w�h�q�im
8o������K��;jj%�bX���٤�Kı;1��&�X�%����f�q,K=��>����a��Pʕ��n��q;z��mۆ�l����{����θz��l��mMD�,Kw�4��bX�'f9ۄ�Kı>����n%�bX��q�SQ,K��3ˊXc��9�L�d�n%�bX���nP��q,Ns���n%�bX��q�SQ,K�����&�X�%����&'s	L`���8��j%�bX�}�vi7ı,N�8��>Ea����=�Mı,KӾф�Kı9���2�.�KUW3wfB�
HRB��55ı,M����n%�bX���&�X�81XV(@@��G�gq5��I��%�bsL`sUj����*���aa
HRB���,Mı,K��ф�Kı>����n%�bX��q�SQ,K���{�1�x�X�� L�F�p�u���9�� S���N��Ҁ�pP��fW��g8ɴ�%�bX����&�X�%����f�q,K��3������%��=�Mı,K��=�d�q$�1�Ld��2a5ı,O��4��bX�'y�v��Kı7�{�I��%�HL�eB����$/;�\�Ԋn�B��\c3I��%�bw��mMD�,Kw�4��bX�'f9ۄ�Kı>����n%�bX�N����12c�32f�6��X�y b'���4��bX�'�;��Kı>����n%�bX��q�SQ,K��3ˉC@]�HV��RB���\�a
HRB�oc2�U��<���26��z~���:��m�sph'[J���)Eu�:*郛���a2�l2�ո��lp�{d����ÂÂ�8��V9ܲ�Q��C�.�	��']:�O�z���wv u͚��糜�lm��r���@�k0�gǞS�7i�t�qÎ��\Wnϴ�W!�����	���������˦�\�t����a�av�y&�.�����8� �=�~v��B6�ul�5V�۲k����v:��
��;G N�2q�s�����
?�o����@�v��۹�^۹��U�q��1����/]��ff$s�ۚ����w���>Yh�m�d��qh|�`�ŀv�� }M��mV8��718��ff~�Ǚ�����`]�`=ΰ>x��Ӡ�Wh��c���4�{^�����>��~��.�3�A5��N8
<A=�,&i���\�2�T�6�<�tn�i�ƒ$b� �F6��V��^�����Q
/H>w�k�W�X��\�H��11��RM��ѣ�Qp�j�D%�-`IrH�ո"��HIF�Q�M&�L`��`	�RR�l��q`o��l�:ϒ�'+���?a���9}���즁��� �� �r�-QN&J�R�f���	$��ό��� �� �7���U�\N"b&7�{^����o����I�K$���cCGe�I�ؚ�Z��l�=��
�=����t=Li�L�#0'�2'�����=���;zـl�:�=��ʺ�&�-�8���۹�w���8����n���eǓ�F��15&h�e0��XLE"�fk~ŀv�� ��b�$bm �F&�^�V���ŀ>o���y�uX����7b����<���7� ��f ���6�}�}�X��;D��\|��	���׵;��Ϙx]�q�틴��O)�6�NW �y�m��`-Y>�)��2U*�����v��?(���/��s�ۚon�s�Veq9H��JHh���>���on��vS@��B�8����<qŠ}{w0|�`�l���.��1)/K�s�vۏ\m����q9�on��P����� �� ��8$ujӦNҺolO>^
.,tR܉�-�h�h�=�g�{����5�Q��+�m�������`|�`�ŀy����&�	i7��o�9�������;��h�Y[ܓB`�AH�|���9�� ��f��0ur��O.D�9�k�h�e4�)�}{w4������qh�[0nـy�ŀs�� �	CDR�������߻}��`�N�]��WV�#]��r;:.i�օ9�۲];FGl���-��.�^�� A��@|ݠ-�.]�iФ�:�Eknx��k��c"z6F+��5ڿ�ϛ✙�5��:ɍ�乽^N<���w�]�P\(I�ܽ[vTx���%��1��q�=.���3s����ۜv��Sv�u�Cs�������u۵��Z��k�*��2=�}�wn�r���6����t���L�ɩ�%�DCj2�yϜ���c� �ꪇ\!)�1(��RC�}��׷s@�}�@�;)�qe�b�����ڎ-�۹�^�ՠw���/�@����bx&�C�f�z�V��vS@�v��۹�[k�O&90���bnE�w���/�@���h��hW[t�H�I�h���>�����Zy�M �hU2`Ʋ<�LqG�d�H��i���d��{2qؼ%��q٤�\n�*�٣Dx)��8��n�z�Zy�Oʊ;�{�����w.)f�8��.rjI�c�����*! �v%���n��w� �78�<X�̈w�Cx�IH���h^���ڴu��W���1���0���|�`����l�=*�1LPM�Ѧ�@���h��h�e4�j�=��2���(�%�Srj8-8^G�{1�7a�=���
7�93j��gZ�EZbp�3��6߿_����l��s�y�ŀ=��+SV�m<sn-�즁x�Z׷s@�}�|��?6�E��$q��4u��RM��ѩ>07���@���n�ݻ�Ǹ{g�m�p�Q��<f"�CxO��a�1J`"��0S��C*�%ьCa�1	���*�1~pVm�M�`�<��1u6�� �3-PځB�iqYFB�����:W;�`327��@7�@��D�Є�(��`��Dd!����JDe����x0Hx6�2
C���@4�&$�12�gQ�eíTҗ_\P�F-�;-�q]ă3�1vB�h)�R ��0���df�E8� �C�&�	E$Y���V�*�<7�J
���U '�E�~�s�z�A�lll{���B��`�`�`���z\o9���K�36�7B��`�b#`����ww=�Ѓ� � � � ����B��`�`��R� ��~Ƅ���������`�f���g4 �666>�{�pA�A�A�A��צ������罍;������hA�lM�������q�#KF�+[gHĸ��vU|�(�6�&�/��;B��{���rX��`�mbj���f�z���)�U�}��=����~�Z�?�3�D�h��आ���V8�:���v���F{ܪǣ�z��&��eU�]`߲0����b\�x�=��-�v�Q����w%]\`>s��D��R�`	RS�G���RD�yB�����I?{��)1)�Jb�C@�;)�s=��������޾�}�Q��!cx��/�F���d�s��6#��ۮ9�7;'T"�t���Lo͙�k��ȡ�8�nk�������-���ϐ^��@��X��Ga7ʹ���#L��f �[0]�}�#��Mb{"Q��$��{޶`ݴ`�.Ru�u���%��E�
<#p��f+۾4+|��VF�r^�f���˚��.���n����s�i� ��0��0%I"�!Hk��%]�%*.��U��9�����L�dX�=T�{+���|��wY�u���$۪{`�AR.IKBe�l`ٷ<�V�Q�7�o�v�/V�e&��DӬ�9���8h��K�v�[���d<�ɍɹ72d����Yn�:����yVy�Mu����pӭV�;t���l;�gk�7n���Q�j�1q�^^�G,�Zf�Wv�.�p�Ws�{��w�o�Z�ܩ�b��^��;4]�k�ݣ���u�K�oWe-�����ԦD���������ۚ��;��{��<���9�{R��O�D�5uq�.�F9�j�`Ru�|�dcH���!I�L#m�b�C@��ƁW{^�K����=�O���ȡ�uu3Uf��I:�:���U��^��^�,I��O�N=�ۋ z�o[0=ΰ�t������]E㝹tWK�t��C�ۗv��<�Q&y�"m'r@Pȿ~M!��H	�$��琉{��N���s����~0y�)]�Z��UUf��̈ԖDDU
oU`Jр.�F{��C�I���K�&���0K~�嶌=ɗ�ـ^��@��JFD���������\��`]� �� S�� ��eU\]
	2"D��4�)�w���*�k�>��h߿g-����%I�i0�[Pu٣u�N�F���Nݔ=�3�)G6xn��������u!I�L#m�b������U�נ|��q���0r!z�^���$��.n�䪳���=ȎD���F ������1"��bOr'��'�>���RN���j|�'����1!��� @a)D�� �L�P�	��{{ֹ<h]����_qC���`93AĽx�%l���>Id`	FəC&&�l��@�{)�{�����F ����0uq7rU��eUn16�nz{u�!Ʈ�ݧw[�vԯ����t<"��W��Flȣ��������z�,�-�>r9H$���8nn��U�.���� �o~��BI%T~���0����U�#��s�'u�����l���������V�wm8�re�N�{���/mԅ&%0��9��~]�u�'���jI���5'V(�^*¨D*�80p�U���{�MI9���2(dlDQ���Umz����h�7vрz9��G[s�.�ɹ�����<�.���<��E�[�d�ۖ:�NW�q��ks"�bo?H���9�{s@��h�e4
��@���f!��H	�E]��l�;�ـ9m���,�/쌤X&�lQ�@�{)�Umz8�L����6�Ѵ��qsu7SvBpRC@�������SC߿b���=��m��B4��[w4�s���|Jـ)IV r9QBcH	 �I`N��������=�ա��%k�z-�0F�n�+h4W!n��v��덋n�.�U{un�%vM������5��Td�nw��V6zr�sEx�S7ny��M{Ee��֚ۮY��N1�ݸ�	�ջ�<��ٴh�����9�*��F���D�5�ǡ��X����s�/mF�ay����OFN.�WŸlNr�(�<�x�� �&�ٶXy3�"�����};v�6�6�Y$�Xܩ�$p�r�c�79�%u�����ղ�l��Y�Y^�����4�l�7vр)IW�}!��F���{��F�1�!�w����2=ʣ��z�����$����ɭ܌�ё�G"M�@�������{33��<h��@��bWr(A7���UWX�"9�r9[�{��{޿��09�%�n��SS�*������ m�0�`[u�y�� �M<�]s�V����g���5�ض|=�����e��#hNǺu�츛|�{����`m��v��ND�Y73u7s*���0-�ΈP�t�P�6�GV�H@�������q`�� ��f���u2Z�SS!q�������;��hvנ}�V�i@mLr4ԙ�^�M�즁Wmz����ʅ&$�UAWwv`�h�<�7_��F{e4Ω�eN`�DЦ@�d���[eqHm����½��p筸�0a���f��M���(�I�hvנ}m��/l����S@��bWr(A7���MǠ}R���s�Ty��`��)ԫ��J]�(��d�TwNـn�
�@���� �=��EN�s�=�{�ۚ�_�1�ŉ�#p�|��3 �� �%���V�f����ȔjD�����V����o���ـn� ����QUwt�0�3�l�g��Y�[<;�]�y�x����u:�^��{���'\8n���~m����# �� ��C��C�����f��Jjc��jL�;��o��6{ޟƁ����}m��~H������6�9�K� I[0�j�=��V����w� �uW�4b�Yr$�4=�s��h���RN}��jD���_"�����W���;�,�{�B	��r-�VF��9i��6���S�uV��ՊW�>sݯ�qxrhN5r�������ϐ��y�T�����}�v��mץ;� ӿ��0�j���C���("⩕0T�T]U���1��L�t��m�`ݴc�s�2uS�U�eu7d�e]ـ9M��K#Ȏre�l�-�ƁՕ�����1���C���DDEo������n���z9^��=��E��0mFH�5&h�M܎G��m��z_�X�,��2.FE
a&��#�l�������,ɀ~H��*A�FL���� D��B$�#4�LHHȢ@���Ȱ��W��*!��BI�����	�ML��5(�!�S����dfpf���#�4�E�Đ�bbH r�$� ��SW`hM�bn� �@�������	�86d��������r�4g*��g�1�d@+Ơ<"�l����a	%
	�#�.�� �#�#"A�������F E"E�@����dd�`D��͎��^��v�{���ʩ� ��WR�@�9�-HRy�iZ��@L� �<�'i��V���:D).�Շ�)�]3SZ�l�-���֤ � ?�B~W;� 
��<m<"�h)Id ��a���ԝ�jѻmJm\��<uu���͞F�#t\�̈́Q.VS���ln]pv�6|�y��Zų[�m�u�vuL�����s�������u�6q���)P�?3_��d6N�.�t�<F�{ڨ6䌝��i^�UiN�[���յ[Cb�V�X�&0�!�Uf7��j�^]��^�0n��~c|�^M���x衐@C����X;�P��4,��V5컍v]���,򦕀 �탠��u<���Nx�v���mJF�n��컱�@�C�)�Vۧr�����E��@ⵝ
j!]��N1��[Fi��L>[az�A��45���b�3��	�6;pp#�z�Nnbg�g�c�v���ڞu�]��M���v�G�%X���t������69$Xe��	�	(���iP��	��sZ̉[*�=[b��wϖ����n���iY���m���*�v-�ޢnZc�Q�����v�;&�}HY�,�]ZBm�1�Q͜�a�6��"�L�	�9f�ɂ���m]z��<�f�5;f6ύ�x�e�T���rۨsc���O0Z�`�1�m��e�r���#��[&G��I��kC�)f㍪-���&svu���X�w �cE<�X�28�K��ڶZ�Uj�oZc�]���Ol���8N�E�V����`|�r���a��l �T�-M��;�֣!�V�l�U��Z�K��,�.�bz�g�p[l�ؤ�ނcdw$��u��D�$3HǄ4cMUjX�/��y>i��Jv�nom���� �Sr �ɒ��a�����;���a�7uv��t���zN��T�l]n��2�P\�P��anVc�U-��#��U
U�af�� �1ju��1���֩e�C\��HZӭ�!+fg��u�U�a�@v�w{��Ez*�QѠі�{Ǘ�t�> qڂ|�;G�Q����ψ�|v�Oh�.���m.���E�F랗T]ӠFn�7��pD\,�-#�ݑփXE���;"���]��<X��NA���h��0�W���N�f�R���n�`�]S�Ϊ�ٶ8��Ŷۮvs\��B�������Eō'c��st��c�yn�;j�<bw[�l��\g;;�3�����c�;:Tф�WGZ�8+�U9H?wϟ>`���6\^��������{����`���:}�6�m7)���3a:m3�g�[׳ƛs�F<���yC�ݾ|��
�<#i�S����ƁWmz���g�{ޞ4��g�1F,�9�)�U����Q���0/_�wm�"Q{|����ħ�7��{ۚ�a�s�M��z[�z"">�����]��Lw����x�V�OuV�"z��0�QL����&��wm�rku�m�`vр(���>���2rvy��g���\�)�dN|gsV�v=�]�#���u߽��x�X��e]��u��>Id`v���"9������U����k& nbN'��{��#��`0�$�
VX2!��%0�����(�"iݷ�w}�n�脦M�A�Gx6�!ԙ�z��@�{)���L��� �o# IZ�����.������09�JK�9�� �%���s���r���0�����Ⱥ�����$�� Sԫ |�9ζ���i[0ݴh[B��1�%1fL��Fڅ�7Qy`37�87U��fԗX��g����q��ݮ*䪂o�M]|[y[h�7v��Q?
)�$�{�5$���fd�L�9�j`����F>G#��L�+f -n�}�tkȢ%��;c����`���qf ۿ� �n����DB��(I%�zp�-�Ɓ�;�YcQH"A���G�	ES�^�}�u�09{��߳���
�ȾC"���D�����<���׌�� ��x��ݾﵤ����Һ45�h�kj�;�G\��]x]ɛM��s�������g�0<�U�e�]Y�nـ}�h��V����-�4מG�D���ɏ#��>ݴc�DD�$��Jـ|��"9����o�Q,�97 ��hwm>r"&zݳ �V�{�j����*������r9�{������o�~0&���jO�d�]��ȃ�����M���B!F�X��������F����6�x۶�e"$Wv.���8�s�N��"����gr��ѓ��~|�9�.�z�����w�ݎ��|��7 �%1�5���� �v����s��l�;����bQ9��rC@;�پ���ɓ�[0�l�>ݴc�s���L8��d@Ә��mɠr��@��M=����l��M�XY	�m�d"��09��x��[0wU�8�"-�k�#�"ai�c��4��F���s��m���~0��`P�DB�V!�⬩RZ���5�H0d�"T®�G9à�90�s5<�����m�X!s�/ω�9� ��b2�6�8+q�����O`p^���:�c=�j�-q/�GcG6��{WF|(����0���g�J��m!YvzJ���tb4�Z��l	��՞�\h6P櫞`,[Jy�Y�:8xS�������ul�X�;H���IӴ�.�m�������F��j�%U"j�U��\ܓ1�s��t��m[��f�ɹ�:�Xf�5�s�ߏ����h��K	b����hw����>����`�骪�Z��R����� �u� �;f��f os��g�ĎW�B���i�RC@���}�h��G92jN��l�>�L�ʚ�**jj���Drz�3 5'x۶���9=O�n�介��f�$�*�� ���#܈�#[��@���}��hg2�5a"�k�m�)�Q�,��c��]nؚ-�����q����m�}������2 i�dj6��[<hv�hw����߾@v�M��<�H6���"����P�/b脐��	{�c�� �x۶��G9�DG*��z����.*&��[����q3ԭ�=��@�gUym�#�Cp���ܙI;�:�� �+F�OR�`���s1�Jf(��>�e4�n�@������h�_���<�dxG"Kt=�qrm���"tl�.����g���s�W�\w�3�a��hm����Y�}ݴ`�|��:�� �rIL�C�ԕ53Wt`۪��#��EP6�x�~4�n�}�?$w����H��N~Q	ɀ�׀{zن@��
���I/G�!%��~�0����6S�L�S�8̃�94=���s�|h���@�����~�K��h���`ژ���0 |�wV3�i���@��{�Lj%I�i<��uǁugn�n��<��<���,����\έ��dB��g� �����������@�t^N8�&�E#�Zժ��9'R�`S�0��Nz9��?6[�����	��S27&��z�VI��""g��� ֝�m*\�	� Л�4=��f+�r����+P�]	B�!%�O~0��I-$�ߔCM7"4��V�s��@����>�n�@���Z�s�q,�Lh]�C�x���q�ջ��6fFx(m�����~��k���H���' /��4�m۫$q�Dr>��� ن�s7X!��q�&��;)����31#��Q�oS�p{����$�EP��~�
�����,���0o�&�kT���r#���}��v�;�pqPoɕ7r`}
!D�[�p���o[0w]F���*�q�M�Lcp�w�`(�[�><��I�{zـ%�Q�{Q�����0'�1�9G�b,����/X7��;�N��8-�������y�w���G[�>w|���\6ч���%�^�BT�)�ٺt���r;U�{gni�!�w$.��vT[��aWc[&ݶg[�gQ:N3;>��47�lC��	��D�W�xQ�m�ۑ��K�����K�gk̴n+lp[�]�Ĺـ�/�V����{��??7�~h���)ۋ���,�����]��[;�n[��ysǥ����{�݊?9��/�-��[0�VI�}ݴ>G9�;�9_��C26&�G���7��3&MT����߯ �v��Q$M�Ԥb�i��F�ξՠ�l���~�K��Ɓ�_j4��U@�B69��mŠ�2�w�u;f�Ւ`z#���G3��-���_�P11�c�@�U� |�s�\���6Ru��� �����.5]ǰ񋶎����q���vɉ���.��F�.z�B��h��0�/��� 7y�Т!zC_�Ɓ�g�(� E��I�{^�|?t������A�fEf'�4D������@BMZ��Q�����Τ���vVF>DDG92k�K����������������l��Q�$�1����F�W����U�s!Ħ"ʚ��=�ـ{[�0��XDB�P�;}4g����#y#���-�0�BQM�^ �^�v��j=�{롯.�{����nICf�7m�*�[�a�����'�w��/��	��F*���<KV {y��v�пDBZ÷��Q�z��_�jDئ6������s�`��Lg��~���M�g��?�0��8��@￧�}�{�5*o$��$b�"B8�qd����I���۽ m�&�9�2Lf]�"F�J!�J�"࡟��W;p\
(B�k�)�NCI� $d `��ÄL%eh1���BVB
�R�!&��[ qނ�,`�Zf�7&��!�HɃQ����y�_�4�j�02]���]
(:�#i�M��nB!5(�M��b�PC��l��)$Cf�X���c!��I3M1��F�U�&P
ci�����a7�QeN��V� �|�⪘�	��r��)�(�\��Og|Τ��{�ԓw;�fPi�ɑ8h{�b�}�M ���@��M�ݙ#A E	�����0wU�"{���u�f�-�h��YS�5�5YLy���c<Pg5���2v��-[�`�>��7W�w���|Ʊ��`''����>��>�'��� ����>2�j⋚	�4��>��>庍 �{f�}�پĎy�~`H?F&�G����=�r9��5?^��� ��3$�q
 lnDhyu�����>����El��0�j\�YWeR/Hn= ���@��S@���4.���3����k~I�$" �I9�����5���.�ݩ�l����^/M̗"���|,|��F�1�ܜ���Ɓ�-�h]�z�;f��s�v`���L��@��d�guV }�W�}�ю&D�ˋQ"@�#x܈�:�����4�e4�n�@�}NH��B(�I�`9��w�u;f�R�0���"s0 ӓ@��S@������4�}�p���D/q��U�|����v:����J�,$�3�egW�_��V�,򥻃�9�ݨ��l������d�B>�hЭ��K�!˻�6�s-�v�zz	����&�� dk�u6�v�K���m�˖�sI����au����n��à�/h�ͷ;S��%��,���;U��nQދ���7Iݹܚ�ʏ�pW`�:0�\k�Q=�lU38�R	�]G�)a�{����w�ܗͩ��/�+�'_��x:�v,/1r��%�`�����1�N�t��������n�I�4�q������0�j� ��� �U� ��ɍ7%67"4u�� ���@��S@���7߱"��2d�xLU2U]`u;�>�h���r=�EV�{$�*����p�꬘��(��&��>��>庎��]O�=I{3���{}>�$��瞃m2~�2'Ԓ_s��}�I{?ffW/��$��o��$���I$��~��[���X%+��j�;��,�T6�����z���= y3��z:jڳ�h����6ov�9�v�V�o�s����c�/���.v��}�Iw����m�QN\��m��w;ޝ��(D�y@ ��Q��r��ެն�{��>�$��jz�K��~�H̉�`@�_�33�o$ə�������	(����M�I%��O�I.Ww��$��x��ԯ  g<�5�m��}s�m�sշ�����ݿ#RIs���7��F�ȏ�I#��MI$�����%�˸�$����o��{��}�
Pȝ���+\�L]�[���rrg�,�m\����Y������E�L��o	�i7�$��o��$�;.�RI}�ߑ����i.�|�����"�2$��q1�ܟ|�\캍I%�;~G�$��ORI.s�}��g�m�f${Y�Q2c��1�f�[m�������v�V����E��'�7��k���m��}�jI.���$ dPYmHϾI#��MI$��g�$�;.�R^�����>�$���jrF6��(�'ԒK��}���u�ٻm��}�M��g��num���ݾ��;���skB�Z�f��"�t�t��N=�j뇉[�� ��c��/[U]��3;��L����~�ޙ�6���K�(�ܑ$����|�W��o�H217�H�I%���Ͼ�f~��B��Is�����e�jI/��FkW�S6Ԑ>�$��l��I^vϾ^���~��l��RI{�ߛ~~ ��N��K�O�?{�Ɍ{<ﱽ�o;�j�[m������
�0�lz�Ip�:�"I�Y�8��$��u�K߿g�����I%�}����������������%�����mA��`L�v�Y�=[g�veAm��k���w_.���X�2q$��o��I%����W���9ƒ��jI+��c��,t�Mߟ��������{���{��}�;ݶ����5m���q�{���7���c���{DF�i� ߿����˨Ԓ\�k�>�$�lz�K�U�8�f��.\��7{��(�{����[m�~ܛݶ߱����q�w]���Ǵ���v��F� }�}�ߝ����{�e�$�����K��Q�$��?eY�ʤ����Iyq��3��khv#�.mN��Z5��%�Z�E�9(�wm��-�N�e:배{ '2�A��Uv��YB��x���� �]l��ճ��3�[��P��ѥ50��u����hy�SX��x����ß|��a�8�Y{n�-wu:�7k]� �-�i�U���a��=���4��#���Y�(�w=k�p����fth���� �ٓĘħ�-t ��7�B���L�kr�zΦ3�EՑG��vc���'�[���sv�GG��wwc��o����J��$�����I+�ھ�$��u�J�߃�Iu�:�A���ۍ�I+�ڷ�
��b���ն�s�ܛݶ��s�Ƽ����P��������u���=�ԒW��|�\o��I%{;W�$�{1"�c��<q�jK߿~�ߛ�}����}�j�oq�wݷ�(/�U�}���$������2(�NF)�K����$��k�����jI+�~�H?���~����"'n[�v���N�լ�p��"\^'v^N.nz����w�|{_�m�Q'�$���|�\}��I)]K��s��DDn�̪��&fR���f���-0\�g��m�^wF5P\�:$�(�D(U�L�=�{�L�W:���e�;������O�����ڴv��\� ��}���j�UdϹȈ���i��L�짘�$��ˈ�b�ɊccnH|��~��{�{�1�m����;ݶ�{�շ��1�{��I#�����A�~LM��$��9�ov���=�ݶ_s�ܛݶ�㝸ԒW�g{�B���,0�LnFْU*��YY�����-&v]''V\�6-�����k㠦<����|�Iu���I%yo���%��SԒU����Iw�.� ds�QH�I%yo�������U;��$���|����{����iw�=�B'�"m@��%S�ORI}gj���3?~3��ĀE��� !B	
�B-�VEX!`�M���D$$�w+>�2ff|��zfe��}4���Hp2����_����? ]^��Ԓ\�o���%��[Ԓ\��' �Bǎ~Dq��Iq[��$��ffw����J�|��������$u�Ex��f�k�nͶ�ɶ^�m����
���;�������{�����غ7N���	%o������}��I/�-_�8�]^��Ԓ\�_��/"�i�&L���}�����\�6��}��v�����j�o>�M���wr�������,dׅVo���O�33��*ɟСDUS���ޙ��o� ��v��5�ڂֶ�������{ǽ����wۓ{��y��:���"@6�Y�ȝ
���5�k�{���E��(�RcԒ]�o����(��ТB���ՠt�߫ ��:�9����H,�Nɡ�r�pN��s�Z7f3�`y��������'L7fqS�n�Ц���==ΰN�X����
!%�����=��#IG�R1$�z˖�}	$�M������`����P�!J;�yf�r	�,x��G��o���u�X~�&���=�Հ{�Ȓ�6�E��$z9ۡ�us��qڴ=�q����_ȌO�Ħ66䁠us���ΰK�Xo<R^Sr�-���S{��&�42�Z��+�#6�`Ce%`I	B����b' `�0�A�#� X��H�H�����o }���$HݡC H��	���� �ʥG���h.�Ѝde"A�(������\��(�tU��7��=�߳���e���m�ܐ��.����T���eb�qn�ᅛ����E���)���%�Ʋ�g��m��6�`%�[v�ڶ�@��i5S�uH�)-W,�1*�j1uv;u@ :x�:Sb����v3��F� 6v��cT�V��opc�����9���`�x7��G�D�δ����U�
������h�e!�)�Hk�f;>�μ��mmH!)���*=����keW�BC�Zlmz�Ke��PmV(yccm 4D���N�msZ��6�e��)�j�(*y&��8��PmlXz�E�c�u�Q�N��vNS����qݝ�{t�^����Qڮn��/Zwd����rԡ���z�[�g
��m����
�Ŷ�Hʝy�ά��B6�%�x֖��1=��Cj��A��ޜ��s��q�yw5Y���t�y��;����e,�8���Q�(\m�>O=���c0�A'Q�d�M��m�b0�ɓ�K.ʭfplb��Gp;����e���]��:�U��On�=��c��S���G1�v�;��Z��GF�&�ٹ�l�m���iM�)4ѧ�z-S��\�kV�cl�JKsl��p(@@T���\�ms0�{N�[�q��$����D�e;PQNgÕq���p5��mk�87��A�loY.���`ڤ7O7�fɶ��&�vxx=�� �һ�0�jAX� �;1=8aW��PU=d��YU8����1L�Q�qY^ne����ܫ��A;rlqbM���w's8��Iۤ�n-�H�$*�lc�����m�bl���P���.�sb3ږ�U뮺�۷kb�����!k�BU�x�i�l�wVk�:��'n��u��r\q�Wî�7mQA��dݳ �`�.G��6�&&V@Ij�b5��09Rf̆n��i��ڀY^w^���5n�bKR1�[mUVջ�\��*�Uɜd�fqqns���"QG /���D�A/D@ h��T6<T6
tU8aL�'Gkó�?&ʚ�W2�5g�l����n���hL��ɹ:��܂�gJ�qe�s�73y8KF�@g��5�ɖųl�k�ut�cw[��Y�9Ύ�㊲�g���7llVa�]i�)���x��g��ķ]��L9P: ��rZ��.;<{]4t#�<Å�u]Cv½�3N��mv2q��gb5�1rk2c՞9�;[n��ek���L��6�vS��0��������|��;���XU�'�j���Ֆ5������۱�jTٲ��Īg������3���5���T.��@�^נw�fg�9]����A)��B�Ǡ|����c��\� ���>��L�ԦG�@G1
%�@��<���V���^���k�/]b�1�ȢDm��us�g����� �v9�8%DhQ�0ĜZmz�3����;}-�}�@���U�AE#o&\���02�(��8뭄��ٰv��˞=p��I�$��kHX��Ѥ��/_=�V)�7��}��DG�)��:��MHM��]T��� �v9�Q���P�	궴
�����{䃝�!���S��h��h]��+��v­����A�����MŠqvנ|���v­��/��^�^dx2d!�z˽�@�o���W|�.��ږSl�؇$i,Ks[�M��^^cA��c�KZmʀ{c���������ݮ4s�����Z�}�@�����8���=_�����D�%�hm�DDL�)���� ��F�ԣIF$��@���*��I� DD�""��E۪9� �s��w��pX��~�'��������� J�N�v�u�6�D�݉dbo$���Z��/��u_y�^נugN�Y����<I@�P��3ׇ���8=�ZC]u���p����Ǎlt�6�dZ��h]��^��v�Z����8Ɖ���@��U��#��`��p�T��56����!F��*��@�l*����ާ���z��Dȕ\It_$����s���x9��� ��U�DC�!�B-$0#�L B�@� Tq�1���H6Rd�B���e H�����	B��~�Xu:+�Y3q7S(���h�ՠqvנU{^���U�y��y9�Y H8��������vs.��w+�Ŭ����n�׺����6���ma�"N>W����U�z;aV�U�z�p��ӂō�dI8��ڷ�"#�B~�Ӏ9��`�J���JH%���G���U�urק����;�|�������"܌�C�9*���6[u�uV��7U�p�ڒ�F�c��)���^����_/����Nӭ�)/C�!t��V]Ѯ�Pڶ,���M�\	r�V�`nH��>���ٱ�&zl��.g��F��{b!!��퇝s������88K���×�����z�+)��vt�]s`6b#nx=v`5 c8ݹ���y��6F�.�@����X������tF�-�D��vWCXH�!��i:s�l��x����y��g#f���o^����<�IjĮ�;�������|��j�0�)�:���7E��;N�݅4#��S��xH�E��.#s�Z֖�o�����uX� ��U��h�z��D��D���)"�9�
��*����=����bG�����i���=�Հl�u��S:����t 0x�i� �s�z�v����@��@��D��8,X�FD��@�\� �v9�:u��6y��s�����̟1�����mɛ'r�d1��Ort��bu�p�d����X:r��m��� ��U�vu*�>�r�����,��	����ꋜηYi%���/D%
J��aR�� �[�y��>��?~H��2$�(5�)���y�{�`��8�n�v��-Rx�B�ǠU�נrت�*�@��@��H�fMOȊ9��b�@��������� �(,�d�>�;!�F�#�t���-̇s�U�tv�q�p��	��\͂�!؈�>m��@ⶽ�����V�i���QD�H
7#�8��}�333<��=��yh[^��w"NƜ,n!\��� �X7r�B��Q� �	!#D��X1$Vlh1���W g�;���z˝��-�¦�K#i��ǠjW*p)*�;)*�|�r]6� �_Ȃ^J0n8�ZVנq[^�U���*��b�Q�'��x�xa��v.ōh��y@O��kWkn�,�,�GL�F��q��$�@ⶽ�k�;lUh[^�e��؈�x9�,���JJ��ț�s�9m��V��G|�//c	�����G�_z/-�k�8��@���֮:�1F�(�E�Umz��[^�N(Ȑ� *
@Ps��W�R�v�%QD�8���Vנ{�����E�Umz�hU 4�M"ۭ�y���Wk\�m� ��x�S���؋����T5�G���@3�m�����m���k�8��@��*LȈ6���zm���k�8��@�����9���K��F��@����+k�*����V�Wz�I
*f���"����۬�n�J�N��ru�s�F�*��
�*�e�������Z+�hVס8'�@B�`�`��\\\c��M'G�7$$ڪ�e �k,�+{@��pi��&\���y��ђ�8%���(��m����8�n^��|�����-�����R{;�6�nѶ۶��l�sP �����A�<OPBU�4쫌1��m�ŉ6����O��7kl��W�����ºlP�b=7c����p.:�^5x�rPp�2 �^d�ss���D��7&�w���ީ��׫)ո���`�E�&6��nq=��\�ͭ]s�{L�EΌe׍O�m���b��ڴ+k�:�k�/Z��	�i`��E���Z��]���Z�;P�J(�G��-�������­�ڴ�NȞE�a"YN=������@�v������
�$6���zs�����e�XO7X�����cB�a�1�h&���y�
.I����r���_ ���=/��=���#e���5�s�})*�6u*�7U��N�H˲���J�Aww8��Y�P���d��:��D����^���T�Wj���x�#�̄#q�]���*�Wj�8��@�ʪ��m!<��r=��V���Z��]���VWي50M�����T���r"6�u�
Su�vت�=���L���XОN2,n��ǟ0�[�
ܸ6��ݛ�盓0r���mӉ(Ҋ%��'$��:��=�����W�g�;��-��?H�E�a�4�zWmzm���ڴ+k�;��*`L�#Ho$���*�\w�Sk����ĒI)�K�s� ��	r�hѓ���hW
�r��V������
�E�SI]`�U�2� � 0Ѥc��ԆCX0YujHL�1(@�
µ,BXPYtJ5�k��f �"B����F�P��0,i����uS,H�F-�L:�@� �fAX�!���!D!�S	X�L��9�0�
���2�p�11�.���p�	��_�$�� @#1R���?m ��R �#b�" F�&C0&U\����8R>>:*�P.%D>��5�jI��{��gpK Q�J0N8�Z��33}m��۬gR�R�S�)ݩScS��$�hVנuvנvت�9]�@��ID�8��%!,�s�Vr���]9�v�{vO�Ӻ�.��#m�Z���1�X�B������Z+�hVנueU\j6�6Oɥ� ���L���6Su�l�U�^�Y\�(��D�-�ڴ�mzWmz;eK@��ܨ�(�YBrH��mzWmz;aV�s?frc��
Z�����Z�~�-��NȞkE����:�k�9�
�Wj�8�k�/3����5k��vWN.���=�.��{�/��tx���;|��u׵t�5ʹ�=,�m��c�@�v����������,�C(��#"�9]�@ⶽ�������~�ď+Z��4�%X��8�n��J��b���N oKq�h��,r�zW-z{aV���V��_��U�U{��M��jnn� �V�p�ӟ��� ��U�� �%pH �*!Dp
DT�`(�1
�j# h+�RL�����d�.�έ�EF��|��J��r���܌�$��p���.�v�#�v^H���m��v�Vk�R�@��Ԟ�77 L՞&F0=�7O6�9P��8B|�Of����ʓ'P��S�s�7p�6���I=n{=�E�Z�r����r�ڵ�I��n�v�n�����(0T�2�Xh�;���eY ���k�˻[ �?����{��v��H$	:���#rǄӇ�\�cv�7'fQ�З�[�u���bx�@�qȗ�v�V�����|��d�{è�"J �Q	���8�k�:�k�|����;�|��܉��EF��@��@��pq����I� ��X�n%MLp#M�����}�@�v��������gpK e��M	ǉŠk�� ��� ��� ֫��OAۆ5�X(<]x�n[.m�c��cc�b�ٳn���!�:�e�+9�S�����R�gR��+T��>��M� 4_c��CĐ��5#�:�kՙ��1�@,`�b�I4�q9��ԓ�������*��F�&��4�����V���ZW-zWmz�E�&�H�)��g���Oyhw�zWmz.>ՠZ>�X��D'$�@��@��@��ڴWj�9G�*� ��O&,Df5�i��E@���Z�h�7/j1�eTǣfϧI�ba��̑7���^�ˏ�h�ՠurנw�&*��$6���z.>��5�s�t�u�t�u�{�"eX'7%)��5s�k�� ���I(�QO����j�*�]1�B%1)��$�@��@��@��ڴWj�Ӫ�ڈx�$2H����f~�k�N~]78��X�:��2*>���J��{�x��tk��h9���741�m�y�����硜��,n�6�y�Z+�hW��]���n�9�f%�qbqh�ՠu^נuvנv��Z���(�!BrH��ΰ�n�j������:Y.8�Hx��̎=�v��j�9q��I��*�(�!�"��l���X
X�`"ZJ!BВXJ�,j"���R�!�B+`A��=�L^XɒOqh��g �M��������$��n�_�čq���� n�Z\�-xMp�pv��f���/=0v�t�6D�u��21��mt��+U`:�`�-��E�<�S��RH�+k�:�k�;ے�+�o߿$Tv���&�&����w���]Ӏz{�`)�t5X6Oͥ�@�nJh�ՠq[^���^�{��jL1(��7��np��`<�`�[0Q	��"���tK�T\��)T�m\��iN�V�6�<��կG8�t��l<�Y
ɩ�f^�r�ր�.��LK�+��pW�����=�V��u͢ ��N�u�L5n#eۇU9��:�nܓ�,�n{8ݸ�ݣ9K.�VޙW����%�
�(9��V��tu��Ξ:�z��\��=�q�t�n�� z��+��QVv!m�l�+�+m�x��q���po7`��x�0��x�%��䳸od�{$����<vNG^���b������.W{^���^��ܔ�9]�@��L�x�3zWmz{rS@�v������LE$K�O$q���M�ڴ+k�;;ΰj�&lr"�fiM]ګ0>��'�Ӝe�X�R�uE� �z��ڏ�1)��#�@ⶽ �-�{rS@��@��ٗ�����!!��Қ�u6Vp]0A�xҁ����5�l3��n�.h^!�#M	(��''��4nJh�h���*�cQ5��~�����9�lʕ	
bWB���¬n�Š��@9�f���:��E������� �i)�I^�L��� ���@��",B�a '#�@;m��-�m�M�}�@��ĶB	�3"�hܶh�%4q�� �h������0m�ֆ	�{ܑq�Lu	�"��/'\�qR<��=t�S-��I�2!&I����?��}�@;m��-����J2!�nLp�;��9�dn�����Z0��&BG�dǓJG�v�4�[4`':�V� `���1�'0�ER�a<
���sFMI;�~��;'@�m�����]�~J""&{����g���;V�v�4���ێ�&��UIswX�B�ǒ�zz ���qrנ�PY\��G�F�`�c�u����8^��ح��ѝ��PP���&���",�G�<�@��@;m�R��G�n�C.Gq3ArU���\���=��G&M�n�7��ڷ߿f$__b[�Hl��Ȥ�g[� ԡ^�93�M����{�_�Y�0���= �nY�s�ՠ}y��R`&�FJ�DB�KRPB�#�|������'�x���b'�L�@��@��@��@9ۖh�H+�yُR��R�f��Z$��ܹǓ��շG� ^*�f⚺E)�LM)Zmz-z�ܳ߳�����WQb(���=��� �nY�s�ՠqvנueUV�mbl��DR= �nY�s�է�b]W�z���@��F�",J~��$�9�j�8�k�8�k�v��u�Y�c0�p�Šqvנn�s��;�7i��-t��R�]H��:�ZBM$q�;*�@B�.�j8�T�i)��C@���w��&3�K�Ĉ�u�IMY�r�Gtb�@��3iP6D	 2�`%��!�H��S�� �58���/1��MJ<!BY!�ؤ	K!VHc$%4k&s��0���� �zK	m0@����)�D��Y�d.X&��I�^fn�>�&5�%9Wg�McZ�ҁ��q�-�DL���t��VFHM�����k���C�D��@$d�X[R%�5��Ήk�	L0i�in�y4�M��9�j�����\b⩦�"�H�L1,��t�fB3\&w�����^���w~~~?j��ɰ�J�UH��k�s�s(R
ٴHl�����)qp�b�v�Dq;���V�䞮IIj4-j��	�nugjZ�`�V�B٥YUV����`�v�H)Ij�#��[�S��Q �1&9��O2�t2���;Uہ�6�Z�u�ʦ��E����vn҃`z�z^y���^ǓM�l�؟.�|�WUs��kn��(=�)���۳D��Ě�2&�A�AI�8���w$�E��U�n���-u6��Z���$5T4���m]<����E\t��*Z�I Dt��Z�H�v���ݨ�n�м�{��z�Q�.]kv����gz����b뵈�C�뫹�rm�ɯWl�lC�/s��$�M�&p�Y�.���:U�����9ؐu������.���`�]tN(��6���ر�oc���G&�k)!uãz���"{m/Sk�v�C���e�[k)�M\lRʚ�dǍ���n��3�S�]�Ey����5�����ÕV�F
��v'�0�6�,�[���3Q�s�����2-��М8���%d��>��Z���»�h���\q*�v쬻[U�t���<�Zӌ��B�-�ڀ��Z�܆�(��"+O��^�*�ԏ54��qb�-[FB���8�N6��{���GL3d�Alg���|��Pˀ� M� �^�4�٤nk`�h�L�k�u�g�ְ:��UZ����Q���%+ n����fI�,�,
��T��������1����Jb���͸W8��W��V;g]���X��c=�'(&jt�ö��]m����İF;�,�rl���I$wF�-�jl��q��Us�{Z�k�g����9�<<:Oj(�ۑ�ၼ�;��]>��h�+I���X��Ss��gv[v&:5�p I�#Bٛv�Yyʖ2�K��zꭍ�vp�U[av����g����Cb�(	�](m��ڠ,s�US��79�o�Qtd��Lh"�D�QraȀ:��F���PA����~p���� ���:�*:u,��\�`K�@�z�(���
;e��®j�;���싍������m�����m�52�󹋷��c�]8sQ���!Ψt��޴"n��g6�]������p��/�:˭�ݣ��j8��^��:3����s��7D�����uϥ�[�W�vu/m�wg�/=L�kإ�ss�:W�����k���q�R�~w��ǽ���|�+dq��μ;�$ػu9�n5 b���R�֜�����V��fb�1wf�Xt���N���?(P�!�����d��%�a1&'Z�ܳ@��@��@��@���B �0�ǉ�$�9�j�8�k�ߒ�_�����|�K!�b��8�=��]n����uB���S�l�Mਔ���8��[4b��z|z��^���<ס"�2d���U�\�� �ʉ���V6�bt�m˜M��d�w]OCQ�X�'��JI�o��@��@��� ;�zh�3�p%?F��Wx�79�ĕ��8���`ks@9ۖh�蕘�<0�pr-g�� �n�y�x�78�S7H�X�0S�8���h;r��v������鈱Ac��#�L �W�>n�s�)���+�>����LhX�5bSp��e�y�2��N�"u�������h:��G����՝�rg����7i��;:�`�J��} jp� ����2	���-��� ��� �nY�s��h\G�F��VM�� {[� �i�	`
IE�lU=���wWRO�9�jI�v�V�mbl��AI4=�?g�}��z��^�}�f�{���DX��U)�Wx�s�g�� ��x�Ӛ�v�D�4	����#"\�Κ�J[�S�����ўnLەj�n�gX+��t$�8�Zmz�-��ܳ@�j�/;�]��E1��IǠs�o�J&C����7��8�7Xo
�ԲȄ���;r��>ՠqvנ|������%
���ǒh��8�����X�8���BKb2Gw,�:�j�� ��k	Z;M���u��;�=��po37_x�˂�uʹ᧠\s��(=`����7Z|g�X����gYmQ�g�q8$%֖>m�'�� o4� �W9�7���:S�����1���z�ܳ@���h�h.�����"ĦA1I�`mj��IN����`��YD�ƘD�C�E�s�ՠ}��`uB��s��L�'x�T��ȹ�����5s�n� q:�;����9�j�>�΂+z�N1HL�H���b	U�A��dK��:�2�4k�A��Q�.nd����QC=�6̫�8Xi^{/]��7�[�C�0�U�sܽ[s��A#t̸z:�Ң�FU��n�oVEŷ>��\���.y���c�EhNi�h�e�hK��ŉt��3ɶ�x͈��[N��hO;u�K��	��r.�b�;�7n7l�#�C���]�n����wq?��7h�:5q�^��s� ��-����9;t�h��:��o����n�g�:�Ę'!�_g��}m�:�Z�즁�3���X�Ƈ�<�@>�l�7���=�l�����>�e̵��j94��-��S@9ۖh��W3���%�ۋ@�u� 7�w��w�oSs�t�.]7��C�����f�}�٠s�ՠ|���f~��}0�g��D1˓�b�K���ke��ᗁ�N��Y��Er-�71�$q7"d�2�L��v�h�J����� jp� L��.�f�`]�U�����UBP�P$��D�DShTZ
:����Ƥ�}���I7�٠^w#j�)�D�z˽�@7�w��w�l�u�v�r��&F$Ƥ�@9ۖh��:�Z����t6:Dک)Uһ�w;�;f��f >i��v�N�b+{\�m]0��\�3�㬎�<pp�nh-�w�v��!N��	���5�m��� �u� 4� =�� ��;�)�	��>�e4���{f�{e4���یi6L�1) |Ӽ ��xb��F��B�$���$ �%b�Q~D��X�I([�nـou� �w*�\�E��ŕD���舝�Np�� �m� /nY�r����h��ȴ����ΰ�N���8���:�	՛��w�:,��.\�`�ѭ��n��C�P�`�l�Z���������nW��+���}X ��x�s��78�ԧ�S#&F&��#�ۖo3ٙ�����@=_���:����;�3	�y&��>ՠ^�V���@/nY�qs�� � ��2(����������:_�Հ�w���J����;����,H����@�rנ�,�7k�����?$����z��
h���.-�kq�8�5��#�^$��i��ݎx����7��f�Zیi6OѬ����g��;��8�J}�r>�7[�S,�vYD����JL�@�,��z�Z�[4�������zD� �"$�������^�^ܳ@�,��y�6� ��?E�@⽯@/nY�w�S@�v��;���ɑ��#�����ـ>�� }\� �BGw�?�˝���:��˦�u4�]s�=u�kjݺ��==��'6.6
�6�cƶy���Z݊�J�(��1��;ŭ�mn�B�� \u�d�3W��Ꮝ�km�-��GJcҥ�4C�z��d�Z��;s������S9�d#��۴jx��{&Qy9'����[-^��5��Rz��zѡ:�5��y�����=o9�ƛ���i6�ݔ��j��������|>7���mN������i��sVy�˫cM�Oe�n�sy}��<�W�v�m%8��?�Ȉ��>�z�����D� ,�ډHh�h���-�X�l��D%'��|J�8� D��Z��Z�^�������4y�-���یi��A�G >i� ��0������<�ܑd���&��4�)�{�����z��@/nY�Zĩ���2(�X�f��ƀ�Yۊ���'��%s��p���+�us"�H���r"I!�^�V�{�M ��f�x�Z�cj�"YŊ~�8�n���3ٮ�A����W��i��� }M� �tڗt�#y�{r��ڴl��Wmz�?J���Oy&��=^y�N���)IV -P� R��Ԣl"c"�-��h�@/nY�^�V����F�����q�CP]*�uZM���`��Ϊv<�8zc��4/�نj��x�	LpRC�����{r��ڴ�)�U�U[sjd2F��{r��ڴ�)���}�W�Ɵ�E��S ��$�=��N��Z�
#��&�ʒQ10"�csp�0���d;��t��3�R@�5�� 2�j�������-!R�$�,d�+H2sMMF�!2�I3P��G�Jd�y���h�q*�l*F�HB0 F~�Hl 0(����S�9Ҋ|� �����E�"|�T&��(�����Y���4�tY&DH�X�`{�`�N����z����,S�p�/_j�v��h���hU2`��l�su����b7\�b�x͑�ڞs�/%���.p���L�Lr$ɑ�27> ��zh�ՀwU��9ȏ��� � ��D�M�C�I�^;V��Go����- �nY�U�'LQ6	La#�@�l���e4��f���ZW;R	�ǂ�D8����~^��ho��@���RqL��@h�B$`��|OsƁ�U���ƚ��R�Ӽ�`޶`���;W��Γ�&�Ʉ��@[mA�>���1�b�y�獎Qy��xz�(dn#���� ��0o[0��`�����,�ŀ�C�C@����g�H����v禁ye7����H���䂉dn&&�W5s�5I� wT+��G92��0��-��銩d���DI�s�w�n�f�M�������U��
C�I�w�S@�v�y||�Ӏ�;�+�&!DLD�F(�����*Mu���NgE"92ܧ�Zz�v�q����p*۫Xp��J&�;	�d��h�������{9�j����g�u�J
���|�������6������\o[�3���Z۰:v͜�h000m�ع/ I�΋���zڕd%tt�"��nN�ґ�\�(���s/j��v�F��E�S�/4�V��%�31��6���y����>A%6	��\��\:�n,;��2w8
�Nܯ�2�j75�8zĩ�΂�ݷ�;�vV�������]� S��
`��D9�Hh�l��ܳ@�v��vS@�*���6�!�4����W�.�S���u[0�� �����Y?%2	�2M��g�^�������@/{f�}��z2��Sŀ�C�E�}��hح�� s�=4��hօ�!�,mFa#X�Q5-#ۢ�-�6s;v)���nM��ۯ&-:�	dm����v� ���4��_߿~�ϐv�yh���d�Bdco&9&u$�s�s��d��aP�kS;g����@;{f���Ԍ�����G�h���9]�O�ߒ���@-�zh��b��D%1�9g����E/g�8^���^ �IN ���,�8�X"c�I�{�M �nY�^;V��e4��F�$Xb���C����/[�@���.�ۣ�悩���
3h�]�d�~���5E����d�A%!���^��,��,����t�N˹V���Y7uj� {M�~��	)�{�`+f w�
��s�芡��_��.*	����� ���,w��~] �I��0a!$� �)�Ϭ�M����ݒHH�F�b��n9=�Np'��Z� �V�y��Y�%	����)�w�,�?��|����s�h\�2L�"'"�qɶy��j�y�_$�;=�Y��q]�'j���듭�J"`�2H�
C�I��Z�`���sN�̞C�75Ajb���p�h�܎r#�Pj~� o��s��o��٘��i�d�ǂ�Qݘ�n�uB���'8�l�ʺ�nc`�2�94=���{�?��{�~��}��RhX�#Ɗ�1P�jP��y���{�Jv]ʵU5j
G2M�}�@�v���^�w�,�8��V+!cā�� '�d�8y�ZBN9e^{x�^of����ܫ�Nn��Q�:��7���Z��� �nY�}�ڴ{tnH�YŊ~q8��{^�w4� �Ss�{[ŀwt\�Ws4Z�&h�*�w����~�P�g{��@;o���0�,H��$�=�ـ{]� 7��Д)�澼 ��#��#�4�n���]M�^ �k��=�ـ5�BV�rK�w{�������ǫ����tK��˔Z�j��C��hA����v���q�[�kvK�&6�֎5�e��u m��,�J�&엋��n�<���<��\uW��5���Q��oH��Pݸ�C�d��;�魻.���7c� C�E�-�u�����+��+�^�5٩{e�n��#�O4]�H�{s�x�Ѹ`�[�1�PR��u��qcR7���w���G=���ke���D�=p��e9m�۰��wn5��{b�y��Ԅ:+�Z˻Q�0X�Lss:^���s�f��YO������Ɓ�^^m�Л&2n< �P�G&E�ـkv�mj�U�E"ɍ�2
G2M��h�S@⽯@;ۖh��DɆ�I��hW��{r���s@��F�����NI�+�Z�����,[�`�"�&�.nɍ����s�=�Zvx=bt�8�ۧ���r����=u��1֝t�t��m���~�0w��h���|����@�¬D�B�Ԕ��]��lƲ#!D(�;� �Z� 7T+�����u̸���XW.&ʻ0�� ��u������hw���HY�'!�|�k��a^�Ց��=׌�Õ.���51#q�9ܳ@�;w4�e4��z�f~�ݰ��A��I�J	umm�|�9e���MZ-g�j��j����$�(�qc�ә#�'�^�nhr�`�εz@�N�®j��ա7t]���=�j����������g�ߒ=���G�5�#19&h]���>��s��	A4E�q(J����,��X�sF]�U�j��������N���`��`~�В�o?~��?J��Y ��Ji]ڻ�7y��?(J"7����oW�N n�w�o��>��F���u��\�V9m�1�qֵ�����d==���4P���n,���{[ŀ{i���N��x�
����Jc`�1�܆��;V�~�ؤp� �o# �V��9����uU�mLD�zo��@�-��9l���{^��j�\N,hc��#�&��"V��`��:�T�z"#��#�G�{�v������T�T�ݫ��X��0u�pw����,��{����'\S<�l]�a.�da�*|����� <��kGMr�[�8��5wk �s������|�"?B��������OT�d���R- �;
��"��0�yUj���S%��bl)M+�Wxkx�kx��3�S�h{s�@>�_Ȫ&�c����[�`��sN���`yOJ2�Ll(�nC@�}�@;ۖh��ѩ'��{u$�hT>�B���aYZ�~H�FFC
fq�4�l���H�"�2"6)��	���h"$�,bRhXa` �R*�����`�$��H���S��M;Q<�r�`�	�-B��[�#$�!����K���"RґCt&��8�a�3�.$r� B�3���xf �0CA"c0#CfR"$*49C��͕	D�8b�kNQ��U�A3�#@���
|.9� @���t�PÑX�"K
D"����]�  ]��g9�i)�ZT�U�Tv�M�:�d3MH5�z�BP��mn�nN�x7mu�x��U�aeG�T���KS�RZ�p��Ut�jn�+<:$#c����fX*���u��V�Lv�T���<Z��.cf���Rv띸f��i.���e)���id��1�-�'Օ���y�%�I��f��7���	�^Ivj��
ZE���h�`�o�n>v~Y��ja��T
�[f��f�P�I)p�a���I��-�U�Axj�Uyv�,���g�$�R��8�u�]��bӡe��N�������yP��<�[&��^��E���f�s�Ѥ:�Lun��t�zع�.6�t�۷7m��j��:��܍��c������#��N���;J�$�bym�J�#�c��� �c�,C��G .:�*�pO`�aHУ
Vm�Px�2���:�j��|�l[Pk������-�����3�%�'F�{okK�4v��i`�G/�ϕ[J��D���r!��
gnmU=���g H�Y)�sJ�5�!��Zε��ᛄ�:�A�[�ɋe�nv\.�n��ӳ������ ]Vm���k����Z�^#nR%Z u��ƐYYJ�s��ZU���Pdw����+']n��'	v�U I,b�/��A�Yri<m�U@s��*��V�;s��*wN�8n#���"��⢍�5��8C�g�s��J�UKp�U/I�5��RK�� �^�nT	Z�<-���W�ۓ�Q��>��謹H;v�:f��W���������9��K.���[v><���U�>F^���\��J�t����5�@]�x�ǖ+]�pj�a������R춑�9'Z�03#U[�*i�X콁5�v��ռ�ݱ-z0�m�$�CI��Z�W�#M�n�Մ���i�P�bq��X�=�T��%��6	����"�J��#N;u�4�d`6��	���@C�Ը�d�ř̅��)�E�!�EMa]�$�yL ��(��|@�6=0��Cc�U�`���\��k%؞5[[Ue�=u�k7�t�7H�9�]yJ�HNHx��wl�/ll%���e�.��{�q�4�P�vg���H�b΍9r���2WPT�������R�@.��:ڷמ:��ʽ�ݶ�Mpƣ17m�p���lóeݓ����\܎½�W��� �۶	�u�=F-�qt�s˛���H�y��}���`l�T;td{.����_��?9�6��N���m��r���j�X�bs�ݎy���_����|F2*\n�Y��o���zh廚+�hW������ős�s$�;�w4�n��{^�w�
��#��=ʣ̇~�����$����X����`sN���`�\nH���Fc��@��S@;ۖh�n��e4���ȇ 67,��� ;�w�n�ŀkv��홶��{��J�D�\:�sxk��5r�&���v�X}��e��^��Ѡ��7X�<*j�������0k�`sN���"��ɏF8'3@岚�0�$ � b�Y�AC;�܎r�������T� �udg���ʚ�21�X������Uk�@�;w4[)�T�b�mOȄ����N��x�nف�Q3���@�o�$�E���$rh�n��e4��hZ��9B��7X��2��7&^4*�&��t�Ц{W�`L��W-��u�#��n���}V� �j� �P���Ajyj�7$P��XFc��@9{f��~��ىN�[��:��L�S�˻�n�&�Ț�� Iüz�F�|9���IFg՗�w��, �AĔՓaRU�+���X�l�5�ŀ�,�>��:��,1�9�-��<��ŀ�;�;[ŀn𤛧R勢��j�kSt��L7j����Ǔ�ly��uG��.B㶘�1������>x���xkx��l����LPm��s4��f��[��s�ՠr��h�n�$��S�L�@�o�M� ��, �i������ɉF��F���v���s@�s�s�4�T�(�c��3>�[s@��)�F�ȚƔ�@�� o4� �o�\� s7]��ͦ��F�
ȱG<f�wfBr>0;���鴺�%��M��\S��q.��o�;�I��;�{f�q,K��s�]&�X�%��w�4��bX�%�	;,ǉ�s0\Y��s��Kı;�{f�p���1����I��%�bw��l�n%�bX����t��bX�'�Ϝ[1�c2`��1�q�I��%�bs�ﮓq,K��=�Mı���LD����t��bX�'{�_��q�7�������ߣ6\L=ߛŉbX��}�I��%�b_����n%�bX����Kı9���I��%�b{z����.-�2ْ�d�n%�bX����t��bX�'y�zi7ı,Nw=��n%�bX�罳I��%�bPG1���Ly�6�q�8y��Ms6���Msu�� ��w=����A!�x6#��x�H�����lB=��1�l��2� �>ヹ����[M�.m�]�����ո��g&(��H�gl�iOm@��v��ڸ��ʎ]aԶ�E�2�]�X�I�n����[N�&gvb�[�r�b�Ean����o��]�iu�ܽ73-�n���ջ2�;�f�1g�
/�
���7�����6�謦sQ������&��n��2!Ѳgc���9���;U%��~_w��=�%���k�I��%�bs�ﮓq,K��=�Mı,K��Γq,x��{��ߦ߭��%�n���w��,K��}t���D�"b%�����I��%�b^{��:Mı,K���4���@�LD�?~��fg79�3�Zf☗Ɠq,K��~٤�Kı/����7ı,Ns���n%�bX���������$/��>�����M)��s���n%�bX����t��bX�'9�zi7ı,Nc��4��bX�b'{��Ɠq,Kľ�'���I3&I�1���t��bX�'9�z�7ı,K����n%�bX�罳I��%�b_����n%�bX��}-�p_D��ٵ��.dظ::�
vGY쩷��GRnW���V|ױs��^��;si�����"X�%�{��7ı,Ns�٤�Kı/����7ı,Ns>��n!���������͞M�ҵ����X�%��{�4����uO]��K�?Γq,K��s�]&�X�%�y��:Mı,K�z�����Ÿ�[2K��Mı,K��Γq,K��3�]&�X�P!���{�~Γq,K��~٤�Kı;��y�3����Lb��s���t��bX�'9�z�7ı,K����n%�bX�s�٤�Kı/����7ı,O{>��̖�8��ɜg9�Mı,K��t��bX��#�����%�bX���~Γq,K��3�]&�X�%�~�����N�����Y�7W�W�������A�9�-����ъ��Xl�;��33��:Mı,K�{�4��bX�%��=�&�X�%��g����&"X�%��:Mı,K�}��c�q����3�����n%�bX����t��bX�'��}t��bX�%�{��7ı,N�٤�Kı/x��1�6d����I��%�b}���I��%�b^w�Γq,v$`� $d��H��>�\*0H�D? 0@���*��J��GF�D�N���Mı,K��=�&�X�%�����=�0\���3t��bX�%�{��7ı,Ns�٤�Kı/����7ı,Ns>��o{��7������6��ɸ�V�{�ı,Ns�٤�Kı/����7ı,Ns>��n%�bX��ﳤ�Kı>���X���i����f�5��=��A1�|]m�kv4��5�v%n��·gFb�ɌK�e�2\d�n%�bX����t��bX�'9���7ı,K����~@�D�K��~٤�Kı=����uPE�[��u|�~oq����9���7ı,K����n%�bX�s�٤�Kı/����7ı,�~�ߧ��C<�sr�|�~oq���/;�gI��%�b}�{f�q,KĿwǳ��Kı9���I��%�w�������u!НCO�w���o�� b'�~���Kı/=���&�X�%���^�Mı, s�O0�`�&B`¿��T_���ƞ���{��7������ߋ2݅k
��ı,K��Γq,K��}�M&�X�%��w�Ɠq,K��}�MB�
HRB���ں�.j�J����ec#Ҝ7c��9�;>.�8��/��=��D%����h���W~��)!I
H_����&�X�%��w�Ɠq,K�罯M&�X�%�~�gI��%�bs��S��.if\�i7ı,Nc��4��bX�';�zi7ı,K�;�:Mı,K���4���1S.�����aHx�&�����7�����k��n%�bX��w�t��bX�'{�zi7ı,O���Mı,K�z���2c�-�1��i7ı,K�;�:Mı,K���4��bX�'��}�&�X�����k�����oq�߿��Emen[Eu�ݸ�%�bs�צ�q,K������Kı9����n%�bX����7ı,J�R��}q1l�fn3�]��s�d��Վ����4�n؀wNn!ϨS+7[lg8�)��dظ��8����'G�[g��5�/�ɗ����Az�A:ܳڄ�<�,�g����Վ�]����s����[6�uk��*B��8dicI$��q=��aW��q�^� muO�-n����'c]u�+�m�+t9�q�x����Xw��K�� JM�VG1�
X�(��#�46T֫$�	���UrM��5ڭא��8�������+���ܜ�����M)�(��wWc��
HRB����d/	bX�';�oI��%�bs��I��%�bs����q,K��s�L��9�s�I�C9��q��Kı9�{zMı,K�Mı,K�Ͻt��bX�'�罍&�X�%���7�]]U�j�쩫������$.����^�bX�';�z�7ı,O��{Mı,K�����Kı>�{f!ff̘�72i7ı,Nw>��n%�bX�c��4��bX�';�oI��%�bs��I��%�bw�,Ԇ=�0\�bf��i7ı,O��{Mı,K�����Kı9��٤�Kı9�k�I��%�bD?����ߟ�dN�$��e�N�5�Ѩâ���޴[��%�y����N:�xx�� X��3�|$�H����MA$�s��	"��r���%�b}����n%�bX���w�1�bc�lɌc:Mı,K�M����<EO��
7n�}�ﻮ�&�X�%��s�Ɠq,K��;�cI��%�bw��,V�vV娺����7���{����4��bX�'�ｍ&�X�%��w�Ɠq,K��|k�I��%�b?o�����[���������o�}�i7ı,Nc��4��bX�';�^�Mı,��N���M&�X�<ow�����s8�;�Y�����{��'1�{Mı,K����I�Kı;���4��bX�'1�{MĻ�oq��~��?�)����h�#t��B�e:H�胁8�屏_��V�_��u{r�Z�%�1��K��i�Kı;�ƿM&�X�%���^�Mı,K��t�'�1ı;�~��&�X�%��g����C6dř�3���Kı9�k�I��%�b^w�Γq,KĽ｝&�X�%���צ�q,K����Xc����!�˜�&�X�%�y�{:Mı,K���t��c@��S�@��F3�RGlQ�6��������c/��5�\��m�)���$���4!�2�PL��>�*t�oxL&���x<��T��>6(f1͠���"g$&&q
�(�>w� ����p�#�!!���$IL�-s��er0�~�b?#�LD�0.^J=�M�z����4��>�;4��pB7�"B!$� 21���!4��$�$dr�C�a�H��z���Fh �@�$`�",b)� �W�X	�X�i�$`ndS���a�
h�!,����L��>���p�!���GJ"H`�a�JQt��E4�"�pT��"k�{G�.�������(��s ��ȑd�`��ȠE�:�G�@� hQ\WǢ}���&�X�%��{^�Mı,K��z_K�����8�3��7ı,K����n%�bX��zi7ı,N{>��n%�`~�������7ı,K�~�ߌc8���3�Y���9�n%�bX��zi7ı,N{>��n%�bX��}�i7ı,K����n%�bX��a��1�Y7��;m8�]OV�tn�|^.X���г��М�c�V�a|�tV�vV���=ߙ,K���]&�X�%�y�{:Mı,K���t�},K��k��n%�bX��})d�0K���d�s��&�X�%�y�{:Mı,K���t��bX�';�^�Mı,K�Ͻt��bX�'��{��q�\�Rg��s��Kı;����n%�bX��zi7ı,N{>��n%�bX��}�i7ı,Op��s���̗̓�4��bX�';�zi7ı,N{>��n%�bX��}�i7İ6��B
@$P��X�耩x�������i7ı,Os?��Hc�Lْٜ\�i7ı,N{>��n%�bX��}�i7ı,N��4��bX�';�zi7ı,O�=3����:1gi�\�K�\�*Ûvz�ظKF�Śz�oC�]���4xיz��ͦ�O�X�%��{��i7ı,N��4��bX�';�zh?�&"X�'g߮�q,K���K���s�pf�c��s�&�X�%��s�Ɠp��q,N���M&�X�%������Kı9����n'��LD�/���ߊ�����W7u��B���������q,K���]&�X�%��w�Ɠq,K��9�cI��%�b^���rV�r��U[��{��7����������bX�'1�{Mı,K�罍&�X�%���^�Mı,K���'�f�%�0\d�q��&�X�%��w�Ɠq,K��9�cI��%�bs�צ�q,K���]&�X�%��W������~����4�[%�=nMի���v�
�"^�:�2�v�h�ۄA���=Z�I�c�u�=ez�ԎÅ^{a�i�Xۮ��Cv�-�/`m���~Wo�ىE�����Ϋ�:v�Μ�3�h���M�	z1c��CI��\�m<��v�]\p@\�掉G�p����qĠ��������sm9�x����c'mu6�	@0v��s߇������}�;�K�G��f�:V���2�ѣc�ɜ[�  �N�zi���3�ZL�b\�'"X�%��{����Kı9�k�I��%�bs�ﮃ�3蘉bX�ǿ~Ɠq,K��{߮'��Tݩ�5vU�B�
HRB�?��q,K���]&�X�%��w�Ɠq,K��;�cI���T�K�ϱ�H`�Lْٜ\�i7ı,N����I��%�b^w�Γq,K��;�cI��%�bs�צ�q,K����F=I�\R�m�n�q,Kļ｝&�X�%��w�Ɠq,K��}�M&�X�%��g޺Mı,K���4��++W�w���oq��_����q,K��}�M&�X�%��g޺Mı,K��t��bX�':���^�W2��B��Qڧ�u��s��H��/g]n]��FnYɖ7:b�4��bX�';�zi7ı,N{>��n%�bX������Kı;��������{��7������FG�n���i7ı,N{>��n��/TP<�L��'�,K���t��bX�'���Mı,K���4��bX�{��n�v��9�+�u4|�~oq���/;�gI��%�bw����Kı9�k�I��%�bs�ﮓq,K�w��ߟ����.6/%_=ߛ�oq��N��4��bX�';�zi7ı,N{=��n%�bX������KĻ�������:�᭲��w���ou���^�Mı,K��}t��bX�'1�{Mı,K�罍&�X�!���{���?v�M&��:����3)CW<sۯ6<��<��]�w^���*m��씹�3���%�bX���~�Mı,K�ｍ&�X�%��s�Ɠq,K��}�M&�X�%��y.�z�\`���.3t��bX�'1�{Mı,K�ｍ&�X�%���^�Mı,K��}�&�X�%��v^��q�����n1��I��%�b_��gI��%�bs�צ�q,b��}�>⢏��j&�w��4��bX�'1��Ɠq,Kľ���1��`��q��8�s��Kı;�k�I��%�bsﱤ�Kı9���I��%�b_��gI��%�b^����g6b��s��9��n%�bX��{�i7ı,?�{�~�t�D�,K�߿gI��%�bs�צ�q,K��;e�_c|�-ۜ�\f������vip{���^��9�ɂ��E���Ҽ�B��v�X�%���޺Mı,K��{:Mı,K���4��bX�%�{��?7���{��������s;��!G��bX�%���t��bX�';�zi7ı,K�w��n%�bX��}맿7���{������N�����7ı,Nw���n%�bX��}�I��%�bs����q,KĿs�Ρx�$)!I]�)_ ]�����!n%�bX��}�I��%�bs����q,KĿs�Γq,Kȧ�EFE@ L�B��T�b{��I��%�bs�K�ٔŗ&&3s��Mı,K�Ͻt��bX���{���>�bX�'}�_��q,K��{�Mı,K��/�?Ú�[N��3\V'M���	籐��u��xBk
�U9�ɋ����A,���%�bX����:Mı,K���4��bX�';�l�~A�D�K������n%�bX�����L\�c�9�qs�g9�n%�bX�����Kı9��f�q,K��s�]&�X�%�~｝&�~  1S,N�ߍ�9�-�..2bg�s���Kı;�~٤�Kı9���I��?��"b%�~Γq,K��k��n%�bX�w'i=�4�3�c3���Mı,�	;�~�t��bX�%�~Γq,K��}�M&�X�%����4��bX�=�����5��'	������7���%���t��bX�';�zi7ı,Ns�٤�Kı9���I��%�bqO�a �>�E�si�,�dKjc6�"%��]qf�On�[��.�bK"�<�����1������WR�`;l�˲�MͲHu���#�л����j�.�͆m���;��5�?4��vY��''2��Ƞv�ɸ�Ō��[9Q�q΋�7�LӍҴo'M��2
����ܚK�����yS4���^��p�[e���2����+WA������bgW��Av;>��3rd����]�崠�*qz���`˧��}�:�y�=W94j�3,�S�닊��_����ŉb{����Kı9��f�q,K��s�]&�X�%�~罝&�X�!I~�U!���*K*��^!I
D�9��f�q,K��s�]&�X�%�~罝&�X�%���^�Mı,K��]͸��`���q��Mı,K�Ͻt��bX�%���t��bX�';�zi7ı,Ns�٤�KǍ�?C��n���h�����{��%���t��bX�';�zi7ı,Ns�٤�Kı9�k�I��%��{���?\���*�����{��';�zi7ı,Nw�٤�Kı9�k�I��%�b}����n%�g�������������Or*��du��x���M�7<n��s���<պ�zn]W..2bg�s���%�bX���l�n%�bX�s�٤�Kı>�}�i7ı,O��zi7ı,O����ɚ`��1�����M&�X�%��;�M­�$x� ���D�KX﷍&�X�%���^�Mı,K�ﶲ�RB�����Uګ�M�(�.��&�q,K������Kı>�u��Kı9��f�q,K�����&�X�%��{��s�g%�s��1��I��%�b}���I��%�bs���&�X�%��;�Mı,K�q��G�"ND��9ڢ��a�T�U�i7ı,Ns�٤�Kı>�}�I��%�b}�{��n%�bX�s���n%�bX��{-�ql�1���[��kYp�$ظ;;g��#���s�[ԉ���v�<�����mĶc��s���n%�bX�s�٤�Kı>�=�i7ı,O��zi7ı,Ns�٤�Kı=�ϯ����A,������{��7���}�i7ı,O��zi7ı,Ns�٤�Kı>�}�I��%�b_O���䜠���O�w���oq�����zi7ı,Ns�٤�K�13�׶i7ı,O��{Mı,K��o9����$����&�q,K��;�Mı,K��i7ı,O��{Mı,K��i7�RB��NQ���H����Ywk!x�1,K��i7ı,O��{Mı,K��i7ı,Ns�٤�Kı?"�������q�JLX���%҅l�울��`���݅��n���8m�du:c�*�wN�n��7���{����~Ɠq,K��;�Mı,K��i7ı,Os�٤�Kı=�z�q��L�ɜ�1��I��%�b{���&�X�%��w�4��bX�'��4��bX�'�罍&�X�%���Щ
�]�H\լ�����$.��Mı,K�w^�Mı,K�s�Ɠq,K�����&�X�%��y.�z�Kf0C�3��Mı,�1���M&�X�%��{��i7ı,O��l�n%�`P0��'kxF�ZR"B��0�҂f%�}��Kı;���0�L�`�nLc2�9�Mı,K�g��Mı,K�w��n%�bX�{�٤�Kı>�u��Kı?��~�����i���c[��5�c���l����71:�\���Ukt�[md�Y�+x�L~{���oq���������bX�'��i7ı,O��zi7ı,N�=��n%�bX���^����EZ�ww��B������i7�D�K���M&�X�%���߮�q,K�������bY�7��۾��]\��st��=ߛ�oq��;�M&�X�%��g��Mı,K�{��n%�bX�{�٤�K�q�����~ӗq8�:���w���O�=�{��n%�bX�����n%�bX����Kı9���I��%�bs��_l�12\&sfnst��bX�'�����Kİ�~D��~��$D�}�)�$�w��n��I�W�H 
��  
��@Z ���W���*�� UЊ?� c@���  E ������� 
��A U|�*��D  
����@_� ���W���*��U�� 
�� 
���PVI��f,E���1V` �����[��  Q
	"$�� @"  (H )*�(P� >"��R�*��� 
T    �     A@�H�$�D� �J�*T��	HB�X  � �A* ( m���m.3�w�ۧ��S!�p R�Y�(���L�ҩW���w�
�jP�-@ ��` � ( (  =��  �    p    �T�áW-J
� �B�z�)�(����L@!�Z�� �A%U@@l uS 0�J�5 �,(S� z9�q��LQ�P2hW���O#��}� C���8��� �=��q��U�7J��A��U��
=�+q�J���k�MOmr�W ��!*@ (��H��-�uӈ73���� �K3Φ�����l=��yv�x �;�*r{�v�ۯ ���޷��7� ��.>}�v�&�\�<�oIs� �]7&��ܽz�{.�wy�� |��H$  � ϟM�o{.���ɯm�l��xCyK�����;ŕۋN� �t����n,���iu���\ :wJ�r�ܜ�oy�W��,��π��..r�;�띺S��y_ y� P��� �A��ϧӝ���<��qezrz�� 9�n.u����.^K��ޙ� iΤ�v����  7���on��r�x([򗹽y[�����uw��{�ӀM�]ˮ2��K��uswax i�
lT��� "������)S@  "x�T�j��� #��R�yIH  *�J=�RT��d )jJH� h�O�:����C���������y����=����v{=���"�*�3P�������QE?�EPU������*���(���<��5~��a�/&����l��o����bl	���pѱ�41��o����f�Br&�̖�)�^�M]g���g��F�Bq��.���R���K�H.��9𑆶rq��	�LV���f���'�yyf�Җ��>�9��h�,��l�ּ6���Ç���3XoϹ�f���4p	P�Ke�ML8h�����o�B�g��s\�l<燱��h`1LL	ϞA�CB0H2��N����,�$f��H �Mf��$2��cC�C�1R08�2C�	%�ߛ�A����1�}��a��<�hᣛl�INjq�8jͱ�`�p q�#Z�M��%�BA�@1]w�|�i'q1a((0&�2%�hϵ�p�>Go��C�H�H8�� !*��3Y���9�����ku�y����ҷ���=>4m��i�`�j	!�-�0g{��y����B��k�a����X	�ɇ͚�c)��Ԫjs�0{� EڤǑ^CHQ��7�g6�c:��=0�uK��'C�њ��͚�5�B0�8h�֍��<,5�=��c�%$/[�����,M!ځ�JN&)]N{I�ڤ���PԤ&�!Y�'7���t�
��Q$4��K�m#�]�h��j��Uc�w�]#��ƾ;�����D�F���4�jip4d6��<0��
4XA��g[4��p��0э-r�EZ	�69�M�2��8aw��٠��#n�RXfߟ���=�p�~7�=�G��!>Bq�)',�1��/�{���}�l��D(p�	�C�Q�۟/W�n�~{GѠޟM��N&���=�:����|�߂�̃0�|_���U�1���vgΛ]r<8��x�&����{k�/D�JC CH�
�<"�������$�}��y����)�7�� �Rݠ_?���zo�(s��h��@�D׾���~�N��n]v�31��!D�#Ąz�7	�Ǻo��Ė�.U·v���(O돦�sMO��G�u}��c ��b���"�����+f���-4�/wt5+Q�F��Ni��=l5ÐDf��ѳ�J�	9g��[v��޽�z�<!�8���o4^�/7����1�~y�`����*������Ziy�&ܥQt�%R�(j�u.��ȸ_o���xǇ�8l���M�p=%� �$�Ya#�1a�'	)"L�3��������?f�ğ)M����O���ۆ��K&&k=�o}Y�E����G�B��j�� M�T	!5%@a:����j6�[tc�޼���$�Hd~IY�j�
�N&)!CH�-{���۵�)��>s�0#���ä�E{Q�Y�7�Ý�|[7���˜g�k�Xk�0ǭ���S9�6sܞ:<F��_Y�JN��o���|1N#�g���9�k��=��8��N,�&���FY�<2w%�?z�$���K$���b5�d˥`�d%5[4}�Kw���.I\���7�g��^�9�a���$� p`�\d�����V�=��7�,ѱ��E;cm,�ƜѶ4kna������a�_7����;�<n��;o��VR$H�a%����	H�hCp#(�p*1#C�Ii�i��C:���"d%�p٘k�0c�Cf�5���������Anp�K����j�#o�a����A0r)�a��o�k����R��!͊���r�ѫ$.<e�8�%"$�52LLJp�V���}58�khxq�xZ5������ߓ<�m�$���'mc I�$2h��6ś����T���zoьtma�4�t�`�BZ��H��0��]�S�K�Fe����N$�I!�h2p�X��`Ƨ6���僢235��/9�}��k���x�=pg�lf���\֤MYܫ��K�߮�����5?�_/җ�sv��sW����$$�q+�e|����ԩ|@H�Z�f��##4�fϣ���f�9��]����;8F7M����ё��*(d|ONi�o\�ٳ5������I�\��5���a��o4czAX5Z>�7���0�Fl���}�<#����3l&�4I����ba���f��9$Y�XPU#[�C��[���b���L#��p�j!�O��0���������b��	8�H��J`��Y���fE<	�14l8����di �i	u4��#<d�j���HD Jq �u(D$��J˲��&l��OsC4Nh��L�aMI�A�T�1�$`�i#dÇ��}�O��[瞚�/�4!$�/�L�ɈQ$�g��ϱ���&���4Cs�	��I�	�5f����4x��Bt$RV�����ӷ�{�	�[��֤�Y��꽏x���}~v��PF�C&%�af��"%���N��MN���o����_�[~�_%��VQt:��W�P����i�WPy��E�Y��ʝ�����I����
&VbS���L�0�h=I�#
ce`$�I�@�ɼ(�u{���<y��&�\�1J-��%�=�[�L~�{��z��SA�:��v1�C� �p��[8F�|��~w<��θ��(d��1C���`a�T��K�#5I�y��# ,���lR��JnU���s;����/J�
�ߌ׍Ϭt�mk��bF1D��a���&���RF$�"Bb� 0���<���fk<�_|��<�$��vF:��4a��(yij�_�
k����^��i!8��d(���9�JI����J1$�.h�>�I��՚�q��s5�V��ٰ�15A�e������s��6�a��CB�nġ*	4P��f9�Y��c9���s���P�����	4fo��֭���5�Bֶ �4j��><���?9�o	�І����L��`��h�#�IT L٧v��a�NȈ�Q&ﯵ˧۲:�f�Hp���b|y�c��`$�  R0�f�����i�h,4�ӹ������H0�8j����*^X�v�_|ק�
���W���ǑA!	03,�CQ��}�e)���~a������K�O�)xK�]�O������؋��
�����*ARC�VB�}�69��W�%��8xއ�@����r��<���o}+vvZq
T $@��`�5�]�2��m���5��t�N�*�0HD#�fP��	%WI�rq��^����0�	�Hp$�d!q��ѳ �0�`t��!&4FFi#�h��iw����C��4Z0�h�C&N0`F:�1Б�8��lb�@dԤ�� U�wc��U`��hv<$���z���ze�LbK}�Kb'�~����ۜ�V�	�&��*Vg�)����-�edRXT��$�����	0�Æ��=֭FӋ�!�J��f�5&
A�L�0A,�������T�N4�΍����N$
�@A@&A�Q�p�up�ū�����QW�5=�"<4xp#4$㤳V��Fv����3�"��N7<ϻ��+��.M!�J��8�CR	?{4~��e����2D�NL�K���:p~#Q6��Ol���2�d�q�e��\HL(�
v�i�ұ�,�* �a�،�HB!&2j�>���{���jij�`�R��N
2)�2��"	%P�
0a�	%�'N�<��n�k�3���ɧ�3X��d�$�b�Ow�N�{��N����8   	 `��_�  �  �m� �I   ���������Z �am���^�MF�n�`��    ��         ����t��m�M� p  >}>���m�     ��ᴛ ���%�6�V��7[x 	:A�Ʒ:H�"�%�dP�ki�lL�T	J�t������|�*�v�ԫkL���$A�l �cm��h	ia�� �m�H8:�r��禆�W-�GFvqRr�h	@ڳm�++!+,��UU�Um@H �޺���Z��lNK$�َrո�I��    �4T��
�Uz��}�T�U*�A��uU@T�R�˵]v�򴫵U���� ����R���T��;��nu�ye�ڭ�:[	�W=V�WAKF��jC�Z�/gm*�U.�s�J�Ue��5?<��L����lpp�ִ�M�@�6]a�b5���q�+��Uֺ�u�,8�kh�j���i�������*��.`��R�p�vG��Һ1������ÕZ�q�m�{r�E������:�+d���@l��i�p�K���}�u��+������w��9��t��U��W� UN�n�p �BV�����Q��z������bч�j����lu�K{Z|�����2��q4�]� ^Z���� �����oHvCuuc�i��6C@T� Ғ��4U�p���MUJ�O`zB�Y���p$I�mwE��)͖��eSg0�-�m����6�q��-�4P C���*�UUq���	ˌQ�� A�m*� �8lJ�۵�5(N��  �eɋn�lHV��p�i�'%�$ �.�ݫF�Z`  ����ynر#���h
�X��T��[��`[���v����  ��l �  i�`   �"�Q�	 	 �ƫp� 9Ci6-�n�kn p6݅�l��C��f�L�طe��B@a�2�a$�:I 		�����ič�e�  �8L�$.ض�;m���$ڶl �      ��n�`��6� l    NҰ�m�           ���m�v����ۤ�s �ER�T/n��)V��� :ٳv�Hm��    �hfۜx��l l�P $mzl鵵   �`�  6͗L�t�ٶ��I�ώ�\��m�%�m��_]����U[�@U@ �G=�J)$jRkU+̫@U:j���l۶�8�J��U�9m�U�jU[V�`�Iv��x ,6���   v�	6ؐm� ۥ��6��bJ퍌k��َ I��  l ��qa�Z�@�X���   N���`8�M���6��-�C@[v�|�h  om[         ��� ඀� � m�  �� �I!��  8   m�    Y��k��
^i�� `   m���� Hu�xH �]���n�zK�� ��͖ɪݻlm�     �    �� � �       �� p�`   �-�l  ����n� ���Rl    5����-��]���  mڶ8	e���b@��J�� M�.���m�Z�r�1�� >3����ۓ#UHt�C�eZݠ6X �vj�  ���@p�� �m���$�[KjN�-�$�OOA��	3m�)u�8H$ ���  �� @ #Zd]t�@v�l��  �q��� 6��Hm�$��m'OU��8kv�dH6�Eq�K n�-���&�9�	6݁��ݵI� l� -�А   �    � �m��;l���   h     m� h  8 M� n�mm�   h��     m��@ �  l   �`��ζ��:@    �M��;����'�-[nJ  �  ��&�kd����  -�n�` mÀ	 �` ��f�.��H�   k��M��m[[l      m     k�� �o�  pɴ�m���  �m�bM�26�    �pl��J� �X�9�nm���'Kn�pHm�Æݦ0���  [@   $ 
�uQ�+.��!7U*��I,�d����ٶ6�    ��ll�oQ'� 6٭[b��� ;���m�u�H��9�� @�M+   I��P	 I�jU� &�^�]�8�ʖ� �`��[A�`۶�`I*m�l &iE�$n��:��  [l]&�$/Y(  c[��( qlӮ k���     �VP�jmS�ҭ�U p�    � M��ht����Ě5�� �oX� �ms��n��Ƶ�����J�m6ڗ�iV�s�J�V8ԣ�h���̶M� X��$���Àm�I57b�.M��`wI��-��Y4�iA�]6]�k7#�/i��k  ��\�I8��Ѥ�ۀ&��tU��V�\�CVʳ��U���6�+�+i�-�f� ��^��٘s j�
x��*���+uV�����Wf\��\F�%�Z�AiNl	2��֛���U�3,nM�eH[\��8b� "iyS��/oeUkz�ECۂ����V��6�l����||��eU�� ��e�	&�ͥ�n�ʍڪUV�
�ݍ�֪vj�m���ܡ�V���B�*��7E�v8� �v��U����E����@��w<b�S�hw��WJ�u�)<��9�^�rp��!l6t���S݁:h�ۮ���z;EkxՔh�֋�Rם4�6�UݣST�E	��OGl�[V�U)'h'g���[���c���)Z�U�,d嗋�;>��cU.�m��B溠�����UzV�����VPC�����u%�)��NF��8��e��$���mUr@� ���U3��r��=EU�U\��ճJ�T��0�ְ6� b�z��B�r��ְ�VOd6B�75[���s�d�P�Y�p"9g��UT��j�qC�U��8A�#UT�;e��Gc�K�;l ��UT78kfC�x�Fa�_ϭ���7 $�nخl�5�ۑ��km��3]��,��s��5�GgtJ�UTF�:��p��!�gѸ�%��SJ��R�M����V��r��u��L���cm�Ȫ�VNk�a�T�N0���6��w;n� -�r<�W�	V�U�i�*Ci���V��h�m����4P:ݦ�:�^�c�J��.�U�VRLͳc��@����m� I��h��$6�+UU����T�n*Z�c��  l�MUWd����i~Ь�ힺv�e'��ꃄv�f⊠*  .� m���p{m�l[A�kt�%�`    �c���^��3hh�t�96LڹVɝ�m���H  ׬� a�m�m�]e��gM�/otrAK6���  ��M����)����n��� ��䖻k^��IҴ^�t2BM�Λ�zF�53��@����k�jV梷,p���H��Go:�6M�P���Am[V�
^-���j���5<�P8I�h����� $6�[@i!�ɵ�S�*�@V���K�-u �qn���C��v՚�bi@�T��d�6��R��w.��p.c��-��܄ձz�^8�]�l�ԙ����>�@��̃�q�|H��Ҭ�Q�m��T��DdrI6�m��;�-��+�UR��R��ѬK�%�m��`�e���[�����m l-�^4(ei���IZ� 8+jpԄ�ht�	R�p,0[bZ[R 6�Ÿ[@���͑{l-��[�Ue�j%*ѥUK�ҭ�iVr�P���r�T�����Ͱ�6��[y��1�@�@z���۩
^���l�.���Y.Um�۶��,s n�)��tu� [궢��dM��ۜ�����iU�	v�I%�-��m������J��W�ul`BΞf�p�,v[���<�Jj�{v�.�}k�
��r�j�|�7UwmTΜ!mH����6�p+���MJ��mʆ�5R�m�� ִ�,]�l���Ds{iyG0 $[%�v��`m� h�k,ik5-7��f�s��ně.�`]�FVlh���H.[�hv��WO�`�rl�P  [Cm����-����uz�� �@���VZſ��{��w�����6 ����c�`(��x�	��6� ����lO�q��LU}P������ �X �ꠧ��}8� ��]"�Շ�U�:U�YdB�Q !ebAx:���D���$@� :(9�O �;H	Ǡx(z���$�����!��!"��N� p@��H��Ҽ ��� ��|�8J`2�����(��x�h�P �·�h>O�;�PE/�I �P>W�Өz(���� A#���2�u@q�A���i;�!�� }T:
¡�B��EL`謨�T����*� ���:� :Qv��|2A0�$�ʯDC����C������(�pW����4iEF�ڤ� �`�p�'��U_�zJ�*�$��� �ʬ�ªJB(� J���	@��d��~�-U@�u�OnL�� F�  �i��l D��i���Svt�kM�G)�Bb�
�p0�i̘����ˉ��ª�3Lѝ�ۙ�c�qQў�ݣ��C��E���Ya�뗃a���c�`�6�Ѯ�[�;��۷�P�vs�籹9��Td:�nm�6�L�r���.��pc��l���u�c�{�����.�b5&�Wa�a�6���lJp�JN:�U���[[0��B��5J�,����m�  �g�q��1�Sb�v튪W���5��-�m�M)����EkcbQ��.��l!�
ڕX	P��,��lu�P�j��ɓm[8��nm�u��lm&C��k&� -�^�l���U,uUn�� 4d]B�M�j�ǐ1�j�Z�`�B�"�1J������c�� H$���E��v5��U����Ҫ�pٷcm&� 6�Y��r�ܓ��Ih�R����T"�lm��&�7l�\�ڬ*3�=�����+Ur�(k��*����Y����v��x&���up.���g8��3�ZxZN�k�-U�35ll���n������A395nBA�5����Tu��3.��׷�e���v�;�����x��&{\�]a��r� r-s�j,�������w�`c�c��!�{]F������mu�{<�d 6vBn�$!1ʫm�S��v��;��K�v��;m���,���c��H4iz��^�%(�m�T�$;&y�`�q���]^��z:K�(6u��dIi����j4Nm 梊��'cp\W4���Y��[��������u�E�e�m��5���6L��v[lJ�<AOC�����qlS=�b���7C ��n..N�']@t�z{v�oY�m�q�ݢ`�L�K�u��\��+��ncck���ձŒ�8�� d�65��Ǟ 3(�s��g���;���޽������¾�� �>�D��W��~��o{�d�^��T�Z�+ƌ�r�ڻ\�����T��97�=h�g9�>*�ݭ����H<zۍ��͝���۔nP�p�@F�n[b��3�lg{`eU�h�k�8&m0�أz:���j���1�긢�v�-f�Y6��4�mz�Ϯ�9뮶�jd�I�çV��4s6��3!m��,Fnz5͐�ӭ���W�R��jSv�0�)r�KM�q��yݑ�EL�Ó�ʛ�X�3� �M���)�/�j �y������俵 ?�]g�o�鹇sRL�j� �ޫ��wwU�ok�m�w��,�$j$��@-�P��	$���u-a�Ǎ4) '&�u�f�[l��f�[l�C�_�Ac��Rh�j�9hG5 H�jꪯ����o���ܖ��	t1����d��]l�t]cK���܎_5��%L���9�B��;�~ZoY��@-�4�:��ħ�s�ZoY���ج�b��$��%���~� ��j����@=�()�M�2M�I��@-�4U��޳@��H�%T�4�
*��X�m_(l���`k���yY��4�"�翍ոؤ� �߄�� 	����������������vl������/��f��u�I���d�g��g\ݴg��6�s6����@�sP�j�EH��.hH�Ě�rh��@7sj��3mX�m_Ca�6�̞��jh�U`��`}����8P����B(���o�ʯ��4uq�b���24�ܚ��i&9h���#���u	y2�ٓ �8�s4_U��k�oY�wYM��|X1<$X��dX�N��ܦzq�ےsڞn�r��Ū�-�u�:�΂352NE�{k�׬�;�����Z��MYqH<cH� �ͫ�7z��;�y��ݚ�o+"�翍ո��o��@���?(��g��j�;7���ƭ�7RMT����C@�ޯ@<�\��C���I	�;;n���kU�T�#r���:�4޳@��ZW��=�ckS��n/��5�Pm�AcS�\m��.���ڵ�b���v�#l�������s@-�4�ՠUz� �s@�wW$���24�ܚWj�*�^�yֹ�����Ѫ4̙1�$�@��z��>ď��M���`�5�LS$�T�*������XwuX��6n֖�7Kj���nS$(��U`��`wNwO���ߵ�JR���;�)JP��*�^�`�G6
uQ��9k�n�����9�]"���]܌$!����;kNqqd��7I�dv�2U�E�Ղ�ә`�
U�ۧ�E�W���S��++I	�IQ�k��J�Eգ뷍�6	L'�an���8�q���Yu�ǯ)��ނ���-�0�^�ٺ�.�\��Ë��`���m�7]��\mV|9�`:u�ݹ=�s��{�9��y���k���u��ܶ��c�z�;4%�mco�mز�v���i��"��^���ڙ�UJ<D �_�~|R����a�)y߳�┥�ͥD �^�m2�5*�����jR��{�vG��){����JR������)�u���)<;��#���\���sB�"D#�ǵq"~��JR�w]�qJR���]��B�x��L��7RJ���\B��A �w��<��=��߳�R�����<��/>����);w��֌�o6n���3y��ǒ����{�R����a�)y�����)C߾�ǒ��\�Z�m�9m̄%L���5B`�N�49e�c]��t��k�L����ۯ˭��f�����)JR~���C�JR�w[┥���Oʊ�^JR��=��D Q��7I���9)�
9)J^w��|��':8�o��ѵ�����m)C�߼��R�����┥'��{��JS����s4�RHQU55q"(��ҋ")�����)>��t<��/;�u�)JP���û��j7�gj����R���_����)JN�~���)y߻��JR��}ݏ%)Ozv��-kz6f���|R����{��)y߻��JR��}ݏ%)K�w�┥9�.oQ� �4�!�S$�Ļt�9����F�+�ގz3�W0�>^:��/eַ�ַ��)y߻��JR���ݏ%)N��)I��{��)�Hk�n��
M�M\B�
=���Ȃ���{�)JR}{��y)J^w��w�!-7�(n�J*�Kt:�Qd%)�u���)>���H`������R�=����R��ٴ�LM*)�5T�!B[�u�� �/>�w|R����{��)����� �@�34n��7*��r9�j,�)K�����)<���y)Jw=�u�)JO������~�wlݽhսL�)�Gb�n6��p�v8���l=��{l]���u��L�.�H����I�t�����C�JS��{�)JR}�u�y)�q�\B�
3 �m~��s6�Moz%)O�����ʬ�'{�_��){���|R����{��)�퍸�#�jS������!fl��)K�����)=���y)Jw=��� �A��h��r������"�JR�gw�)JOn��JR��]�qJ�{"�;��k�JR=ō�:�U�Rn]U� �Aٳ��JP��u���qJR�����y)Q�1�\B��۲S�UJ��[�����`1�fW��{2�������M�<��xͷV.��ru�)�WP8��}�����������)I�{ݯ%)KϾ��R��ן����츳�� �	F8I#�)JO��vJR��}���)>�w�<��<���┥���v�����[�V��y)J^}�w|R�����py)Jy��u�)JO��w�����%��j��n������A���w������\R�����py*�}��W�!�����2ʷ5E-k{��)J}��~��)=�}�JR������)>��t<��3�!����ӽ�����~O�I�$�Y`A�h\I<˸�Ѕsl�Ԓ�<�!�����gW-�񯾌�+(��vM��;�=���@�&*��H 褓bŋz��n�����ʼ�P@^� �pr�aDpQ�kvU�A,�+��dv�X���Y��m��W7���.�.Sg�ܚ�\��Fc�<�2��F-��m'&�V��l5)$���{X�e��fSmɬ�{��q�ۃ���v{k�;A����}Ez#R	:��+�����th!:\�ۜ�m�y1�%T��Ȅ!q��J�"D#=�թJR}w��y)J^w���)<��.@���d�	ǟ�����;�,�)JO���%)K���┥'��ʋ"D#`<Z�ꁩT�%U�JR}w��y)J]����)>���<��.����JR���r�V����oy���oC�JR����)I�~�a�)w߮�R��]��J�!jk�i.jiT�USUW�!{�vJR���;�)JR{w��y0�!�ڸ�!f�彙$(�ݝ�,M!&�V�eƼ;��ۚ�e�U<kD��5*`�ʑ�u5dB�}�{WR��]�t<��/��w��rT�w�"Ȅ���3qNU7AD����)JO.��D ��~2 � ��2R���|R����wk�JP����!B�a��v�U�I*j�S�)w�߷�)JO��v���/=�w|R����{��)���b㬳xh�[�{���)I���ג���~��R����t<��.���R��֪��fe4�f�"Ȅ�a�┥'�������{��JR���QD �_��q��S2K�c���lm�=����[��6rX��N�j� �\��A��l�J��K�HrU}�!,���X�)w��|R�����k�JR�]��A��X��J��UM��i��JR����)I���ג���~��)JR{��py)Jt���]6[ַ�7�[����R��w���R����w�(A:g��kj�M#`�ˡ
�k��a�$Ɨ3@B}&�b |p��:֎͋�ށ����j1B08��X1�����J@���7@<�l�!4k4����1^�'ϕ�_}4�Z4��i5�kO�$��zM�x�U���Xp�� ��N&�u�LBu��1�<^(+���rO ?(C8�ꊏP �)>�{��)w����"(�{6f��%P�rT(�!�}����)I�~�ǒ���{��J�d���~�������Y�o[ٙ�y����o|R����wc�JR���|R����k��R������J�	Bf`�%	BP����5�<r8I��<�s��"B��n����P�+�FaEvy#������yۛ;��I����<���(J!(J��30J��(H��(J�������J��(H��(J���(J��"��(J3�(J���w���(J��(J��"��(J3�(J��J��(L����~x%	BQ��BD%	BP�&��(J��J��(L���(J���pJ��(O3�(J��J��(L���(J!(@P�BW.�ϡ�ˡJrS*���B�(J��J��(L���(J!(J��30J��(O�k����%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bg�����P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'~����(J��0J��(H��(J���(J��"��(J?}����J��(H��(J���(J��"��(J3�!B/.�K��r��uT�SV�P�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	���?o��(J��J��(L���(J!(J��30J��(N���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�&w�߷�P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'ߵ��pJ��(O3�(J��J��(L���(J!(HP�B	��ք�eP�)J��PP�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'~����(J��0J��(H��(J���(J��"��(J?}����J��(H��(J���(J��"��(J3�(J�����	BP�%	�`�%	BP�	BP�%	��P�%&	���.�BP�%	BP���?o��(J��(J��30J��(J��(J3�(J������7�۲���3U���(J��0J��(J��(J3�(J��(J��3�~��<��(J��(J���(J��(J��(L���C��^�~�؃�47��� � Ѓ����@���?[A%S��'�B1��2M�Fhg5�rNWK�M�j���@S�?w����}v�޶oV���{���P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B}���\��(J��(J��(J��(L���(J��(J�Ͽt��<��(J��(J���(J��(J��(L���(J�~��	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	Bg~��~x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�%�ۿ��xf�[7[�V����%	BP�f	BP�%	BP�%	Bf`�%	BP�%	BP�&}������%	BP�%)BP�&f	BP�%	BP�%	Bf`�%	BP����pJ��(O3�(J��(J��30J��(J��(J;�����(J��(J��(L���(J��(J���(J��>����	BP�%	�`�%	BP2�%	BP�&��(J��(HP�B;��G�tU��!D�u_|���(J��(J���(J��(J��(L���(J����(J��<���(J��(J���(J��(J��(L�߿o��(J��(J��30J��(J��(J3�(J�����8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	���?o��(J��(J��30J��(J��(J3�(J���~�e���n�f��	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	Bg~��~x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'߻���(J��0J��(J��(J3�(J��(J��3�ݿo��(J��(J��30J��(J��(J3�(J��߿s�P�%	By�%	BP�%	BP�%	��P�%	BP�%	BP�����Y���ٚ�������%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP�~����(J��<���(J��(J���(J��(JC����5������J��(J��(J3�(J��(J��30J��(O߿���(J��<���(J��(J���(J��(J��(L������(J��(J��(L���(J��(J���(J��:���7���7��p�-'eؑ$W3i&���Ǝzư<tV^�3��v�����AƝ��Ԩ�;�v5G$�6"���X;���X*�ذG��f�t����j�%�\ƅ)�t#.�8j�aH��Y�v�UNئV���e�j�y�8��z,uo1m�Y�34��.1�X�i��f�9{s�A�8���9�p�^��xLɤz�>6������~��s���!cz�T��H�B����l�]�����aW��l\�m׾����b�c��v��۽�w�a<���(J!(J��30J��(H��(J�������P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'{��	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�&~������%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	��~���(J��0J��(H��(J���(J��"��(J�æ~�������5�ߞ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP����8%	BP�'��R4%	BD%	BP�&f	BP�%	�%	HR����o��(J��J��(L���(J!(J��30J��(O�k��8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP��������%	BP�	BP�%#��P�%	BD%	BP�&f	BP�%	��ڪ�T�[�sJ� P�B��0J��(H��(J���(J��"��(J?w�����%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	������(J��(J��"��(J3�(J��J��(L��[��(J��"��(J3�(J��J�2N���%)MO�qI����5U5Uq"B���<��.��s|R�����c�JP�ݫ�A�Gљ��i̊�94'����~�o�R��}��y)J]����)=���<��=��խgk[ùf�6�x�GJu�X��n.�Om1�e��Nu�kQ�����������c�JS��{�)JR{�u�?�@/%)K߿g��JR��g�ݠ�o0٣7��%)O���\�R��g{��JR���w�)JO~�ҋ"D//bи�LԪNJN���)I�����R������Jp`2O~�v<��>�{�qJR�ñ}��a�h�����f���JR���w�)JO~�v<��>�{�qJR�߳���D!a�`dU12�˪��!{7�JR�g�)I�����R�{^�� �A��C�)�S*���q�P<�7- �7L�V4.�z;u�>X�&ù�Jh���T�[�sJ>"D-y�7R���;�JR���;���)J��D �_�O���"���MMV�R����~������K߿g��JR����c�JS������P��r��s"�ANBf��"D#��5q)I���ǒC���qX�! �	�i�J�Ie��$xZR �D�H���<�s��������)JN�����JSϺwX좪�Je�Q.�j�Drd-��Q�JS��ߵ�)JO{��%(?ݽ5q"(��k���mR��iG%)N��)I�s���)y߻��JR��ݏ%)N�N�]ֵ�u��v�^�ڮ[��K�#�ݍ�g ��v۳���G��&�\T��v��l��;�JR������)>����R��}��R����q��������y)J^{��|��'{��ǒ��s��k�R����t<��9)+����,�kU��o7�)JN���%)N��?���>�~���)�~����);?t�jލ۷�z��f�<��;��qJR�۽�������'��T1�Ң���JR�3���y��7����R�������R����w�)JO��v<��;��┥'���;���~��u�'��5��]�Q�k16�f㛷Y��[6�r�']��77�p���y�ַ��)~����JR��ݏ%)N���8�)I�s���)�����DF1�$d�������ٟ�)Jw=�u�)JO{��%)K��q"(��5R'4ڥ4K�Qd%)�����)=�w�<�� FJ_���|R���~��R����9�h�k{6f��o{��)=�w�<��.����JR��ݏ%(? ��ߺn!B^\.���L�f��i��������JR�ʂ��������R�������)=�w�<��>�E� P�Ә��w{�o{�ku�4[�1p��vI�e����eIͷm��ޞKv�e�غG)x��Gl���cA�T�]��V6gy�� �4� UM�z���i���l�Tx�4*Y�4k,9����T�� Ŕ�kw<T3�3��эƺwAˣa�����9�ѓ&x%�=�nM`���!��n���mrFg�gp��4q�$�r�Q+ܶ�>ܕ�CΘ���}��{�{o�׶�\��c��/H��8��K��V��Iu�.�XȻk�8��<{'V0�]�kZ����)<���JR�g~)I�{�����)w�O�┥'��L��S�U-�9�D �X�6m#��'߿k�<��.����)JR}�{�䟀�靋��V�岪GSUU7�!,�Y�!�7|R�ʤI�����)����┥�zh�֬��uj�f�%+�G�Q0M~��o�R���ly)J|�6n!�С(9�5D �^�]-�&�eI$�R���!fnҋ!(�=�����)>�~���)f�ڸ�!f��R��:U2�PK|o8��dk�t	S�vӭ�]��#q�)�gE"1�����45*h�4��!B���q�������R���zo���%)3{�E�"�oZdʗ.�RuLsU7	JR{}��y`,��		C	 ��!	PS�2R��~7�)JO���ǒ����ٸ��&�B��ng��D�9�ֵ�JR�{��)JR{�{������k�R������<��/ 1�[#
d%MM*��L����ǒ������qJR�߳������ܪ�D ���ɮt��*����ǒ�����\R���?w?~��R���ߍ�JR�߻ݏ%)N����� ۰�n���+��uaɆ�i���\�Z�.�ͺ'rtn����S����R�����<��/��M�JR��ݏ%)Os�)C���j34Xt�Z�Y���JR�����)>����R��;��R�����<��<��ueZ�
�ڵ[����JR����JR��{�qJv��@�1ت�);���C�JR�┥~�Yt��ֵ��k[JR��{�qJR���]�������)JR}��c�JSϯ���՚�͙�����)JO��vJR��w���)I�{ݏ%)Os��\R���{V#��Χ؜v]Wg]UF�Ξ��7i'<t�����lp������r�Xkw�)J^�ޛ┥'�}ݏ%)Os��\R������R����>:j��kE�{���JR���ǒ����{�)JRy��py)J]��7�)JV�V����j�L�TʪQdB�nn��)<�u�y!����w��|R�-��QdB���X�ХU
���{���)I�{���JR���)JR}����R��PŻ��|R����uFf���V�5�y)J]��7�)J?3�����JR��߷�)JO>�%)N�Fk��FE��g�G�lhv���q��]�8ܭ�;�
N�PPqq�[�$�kCu���{�I��wc�JR�{��JR�ϻ����"�ܪ�D Q�;SD�*��5�Z�ǒ��߻���	9)I���E�"�ܪ�D ��ͥB�I(B�D,�T��	��R&�����T�'�����R�������@d�w��<��.���|R����1��S(��5R�D �	!B{�ʮ�������){��|R���J���Ȅ!��%MKr)�LMM*�)JO~��JP��c�����┥'߿��%)K�w���)I!��'�X$+J!�tE7Ȣ$Zd��1ȩ�f؅vnn�f��C���4l�D�c�	�:UӾ�^p�u�Sy�zFY��u��$��v6���6�QJ|!��kÒb�ӨRK�@��H�Bai``d��b"+J&��1� �x�#@C2El���R���-�6l��YE]X����l m��K*��m���H@�g�!���v;Yv7=F#�+VbT�$1[i��Y�fhҏWm��:�_(N�G7��b^�gƭ��`���x9��ӎ�7>܈���ۮՍ���<=К��)7\:z����Ν6t葓�)�0y$��r��q�v�4� �V۱;s�u��7�'P��nF&�M%e��9��8l���v�aޅ��j&`Wf �Zj�m�R� 6�L�k$��[qS6�.�vb�E���mY���@����$b��������fحk-�Zn ��:/J��UT�����Vr�UR�R�t���V���<�]*[ζۀ[@m�m� m�i6��-�/Gm5� ��ؖHl�I��R:f���[l�h�u�p�$�[��v^�zIU&���M���J�+�����W�� ��m5R�UVQ��d�a�&$۝��e�����@Y,D��,KdmN^��l���#tWV�s��xj�xl�k��ڭ����5�p;*�Gg\#�3�9�8����%�l�k 'I���`[zk��p��s�eUrv�m���ȓa
�8�$r�j�q��[�3�^;g�/����l�ۨ{/�cq��3�QŒ�Zl��]<�H��[�ضӻ]���ެ\�2f#�O����}�v87ɯX�֝�,]�;���[*h��^��_o����,�vذ���;�cu8qdv-y���i{<�Tu�i��	;�������غWQ�ORu���:��Y �ɆKb�csm)�4�hקn�T��!����Jn[�c��V^�i�YΏ!n��K��v��1B ��㱲�R�4{Zm��u�Bl6dwE�u�vݶ]j�,aQ+�{O7Z�Y��DB�d^9�捓�F�	�B�^̫uQ�u>:)�K���l�mgF�~����[�v�*�9�=�SBK+��	��`筞e���kY��kh&��_���SF z����G�T=�����w���~���$Ҵ�L������t����	�5۳`۞�I7TsSs��*S�>��g���%��e��#=0X͵R�!q�f�K�XI�^ ��)�n�me��7<��fu��<���{m�N{Z�[;��ф��oZ��K4�ۘ]跞�'R=���V�ՆåsŸ,Z��ٔ���+��&��ݤ/\�u�Z��֮�r�]Y4P]�W������[������Rp�,b;��ɺ�D�]))�;X�9�:�sӹ�#uBmo������T�[�c�j>"D,{ߦ�D ��l�<��.�ޛ�~	rR���`�TÇ<�[�Ҥ��UM� �A�w]���/�����~���)JO߳��%)N���s����VkE��#V��nJR�����)JRf<֢�K�B"=A����D �_{�:�T�M�*�/�������)�;����)I�s����\�����)J߻�*un��1�SSSU*>"D.{�7R�*�����C�)~�[┥'��wC�JSޝ����7e9�2.��'%W[!	\��2� ���[m;���]���!�ٸ��fދE�3{޼R�����~����߾�)JP��������g����~����):a���j-��������)w�o�i�$Eh$�*?�M�)I���4<��?g߿k�R��}�vI�����N�W���-j5�ӭ�v��)I�������s��\R��I�k�<��/���|R���|tz��B�S-�1�5D �I
N�k�R�����C�JR��v��?��3Rw�~���)�;Y��z�ޣ[6f�{���)JO>�%(ʋ9���o�R��w;����s��\T!}�-9��(D�Tۦ���P�Ԭr�{nx��3sΛv�����ږ?{���_}�íXZ��de�3[��JR��[┥'�g���)�}�����ʂ�������_��R�����V��Y�5�[�5�|R������<�¨,�^�M� �A��5D �G�4������b�>�����w5����F�k{���������)JRw����BC�M:G�E\2R����┠B�}�E�"f'Mi-Jt�T�R�����*8���?��y)J_߿�┥'{��%($? �8���Q���rt�	S4��Q�O��'�����)��s�R�u�D �_{wNd�۪mUL��n��ôㇰF6���{qӹ�ms�w��a�����N�p�[����:����)JO߳��JR�����);w��~�!B;uu\B��.�>�r*�Js3{�7�JR���� �*���wt��!B;�u\B��^�Qd.I$��^]+T�RRs%*SM���"R�����%)K��w|R�ʤI��`�R������({�v�Z�hΛ#V�Z�%+�C��5������)I��~���)�~�8�	������DL�>����<��;����$-:N�S149���D ���Z�!(�9��o�R�������R��[�q"B���N�l� ���^��q���\�;te�=Zy�p�]�)K�Ϸ�������W3j[mR�&���"�����JR���]�����{w|�%�JO���������7��3V�k3Z���)JRy�u�y��
!�K������)I����%)N��w\�]
!Bn!,[�9�mÔLӪ�3@�R��}��o�R�>��v<����������┥'�����R�闽��0ѽ�����������ly)J~�߿k�R��]��JPrP��;�\B��]�=J�St��ou�oc�JS��{�R���O�~��h}��/��f��)I���py?�?~ə�xY�+�d�&A�5��[S�ƺZ(F��܍ո|;u����s�v�XՒ�Y�ju,�q���e5�\��kOnk)U������z��ʨ#�
�MP��z\�����v$-�Тv�ڌ��)WI�͡y�<�8�;k��q��g�ő��Ûr[�nƎ���b������n%M���olni�l��L�]f�;��-���3���bX�����v�v1\���r�Ec���
�{̺��K���n�Z�����.��+�]ݛ���)JN����JR�}�s|R��������/%)Oߵ��qJRf�p�[M>R�%3R�Ȅ���┥'�����)�u���"��ʋ!r�(dB�k�$-:N��bhQW�!.�ꈲ!��;�΄���`��X���.fԶڥ4�M?��(}��~v=ޛ ��*Ô$�:��75��sB(���S�<��6�3�����=�?��Z�Z��)#K�ۉ�hE�=���㣑�[�k�6���'�^���j��{����<=�*�?Ͷ��*�Ǚ�`n���y�t��^��t�)�QN�� �ͫi$�	t��{�����`��_�P�~�??��s���7JX�uU`~�?�;绳g&�������qS��@Sc��-�~�� ��*���ٰ������b�bMg̘c ӏ@-�M��^�k�h.���Y�j��ĝ��9�*:˨�)�b��3��qbe2���둟~[��ִ���!<��=�j�<]k�z�@/Uڶ!l����O�wOs��6c����<͛�I�sYbЉ���j����`��Y1I[I)Q�(�x�zlV���R�)1~L�1H�>��o�x�vw���wf���J'+���`r�}���M�*��TU������"wu|>� ��*��t4ar�,e^�<�m�y�l�6NZA����z��ޗ��Y6i�"Ȕƅ 7&�u�hy�6��W$����1<���T�2c�9&���^�������Xn�_脗�d;�?���IHRQ.jl�w�ٛVtB���t�{�6ۚ�l�T�T�@ꊰ�I&�w�����`|�vl,I$�""%�o`�����c�����O�k��>y�6��U�癳`FOq3�-�3 =�1�M�)�]�kv=�
�z7eyNF�p'nκ��s+�D$��"�C��hi̺���~�6��U��3g�D(�����sS䤁��rF��@:�&������{�6��绳�~�I$�C��)
���UJjiՁϻ���vl��B�
g�ߦ�;~u`k�ls�e�n���"f�ÒP���t���l=���:�4q{E�,� �1�r=�ݛ�%s�����`f��-D%��?'�?(�h�\�"��%�8p�zQ�۷N�N��Y�?���}:�M���P�t��=8��9[G�22k���g ����@U/���xk���	j�\�[2
uK�����+c(�w��4�Ӱ�6qc�ܓ;9�:�t��/�c7.�t��q��ԁ�On˵AB	��hw]m�X8v��h�2\�D���R�r{&���{���}����pj{4�آ�lNr�-ηn�W`v�b�臖�:���wջcq�]��I���w�V��Vl�P�a�{���o"]�SH�d��
�u`�ھ�I�z{��(��>��ls�Հnk��wL���(&���|��;n͟�!�syՀgwU��c#lC��hi�5NáB{;�6����=��a�	DG脧���h�>Jg��F��= �z��9DC�Ξ�`y�l��5�b��Ѻ�n1crn(M��ԩ����W�/��;6R�sG���-u�.����/��ڰ=���=͞�Q�syՁ�j��Jf)�R�T5V�w]�B_F �рC�9� �H�15�B:D���L	�vL؄�DG��>>������3۵|�Cf��0\L�QMJ�U;oM�g�]Y�D$�(ID����X�~v��V�[x�S�6�����{e4l��
NwM���D�EIN�d��US�������uw?�ǝ�`�U4�tQ���G�M���#�L}�ΝF�L�.�Yڬl�<ΰ:���ubg��{����5��ܙ�ә�}����=^���͚��zCw��V�&~V۩�sCNLݴ_I���j��HnL_��M����_�b�pi�ڎ= ��������x'�$&{��N)0�q��X �w�xo�<g+��3,�=��0z���M��beBM��%e�	�׶��,N�I��GўDql"/��k�����xp&	)w���,�@��b��6{�Cv>��}��)�|��! e�*'��X�	��@: O'���N�'������^� 6�������r�������ƓR4�&7#�b�~�4
��=�z� ��\�*�˕�ْ)�
L�L�9u�@�^�@<��4�����[���c�M�$I,mÃ<�Z����m���מ�\�I�{V蝓߾=����G�68�������/W4��~�_0��`���#���T�T�f��'9z�s$��& �1���ڍ�?��M�k�*�^�~��o�wM�vo:��z��n���2�j����3���כ�`��VP�j�^�{�-QQO�AbNG�Uֽ�ҵ�Uֽ���ܠ(�U�n�˛\� cu=�K.v۱�8�ٻF]r���97;Eӷc\P�O�o���V�
�נ^v��k��s��≲"G#�h[^�yڴ
��@��,ZY�r�Q<�LhRbN-���䘀�{6�d��u}R��6I�,x�G�r����Šuv����w�QG�"mǠyzX��f�WZ�
��@�?/߿�����m�M�;i͛c<\�����Q���F�Z2 �9T�e��'l�gi�.��wgz6�-��ұ;e�7-��}[OW9uq�����oeeA��"��CY�[j�_.��q��pdYy���#�Cqs�w�n��y�F�FX{m۬�j���a��F�qi I�0v��\nقz4������0��k!�[5�6�U��Z���yr�s5�1t���ãۧ)-ks)p�T�����azU��9�[�h���p�F|֚?�m�~��-Ɉ	q�@z=�hIdߒ&)��I'�_��W��<�,Z��4�Q�@�S�X7$�9�6l�+i��$��ޫwM���)W#F�����@�X���h�k�9{����q�"rc��$��\srL@;�1�nn�=�~wڭtF�ܦ{;�kfN#�g�d�H�9-v�' �d����΍�.:��=rK��1S���<�vl~͛ �3f���<�zt��ϾM����<p�G�r��՛�� S��M�!��W}��.��@�[^�u���.fjl�͚�>{�6t%	�}�6]~z��-R<ID?�H懙�P�s�h}�6���j�Nf�Xڏ�'�77" 9#�x/���+k@�Z�sP@*�V-,,ۯ���u�NjX.����WB\
�=�����N������X�TM��bi�������1�� �ͮ��>��ps��1��i$�z.��{�f�{m�����H>�*��#jI�H'1���X�v������Qs�{�1��c�*���܀H�4���@=����ٰ1���O���`jx2�J]T�UX��6$����?�޵`�ڰ>���ߚr;&D*��Q�d���%�v�$����x��(zMnl�N|��֥���s$x����n? ;�ɠy{mX�v�D$�a�7���o"[�U)�NX��f�X��W�!$���9u��u�4ڋ	?���#9�:_��`k�l��!(I�3yU�ݽj��,�L�D�
��sNÔ$�}=�6��U`n�ڰQ�?f́��ۚ�U)�L�rʚ� �٪��
ww��<�zl{�6�MwNdR�Q)ε�z�����YwB޶Aׁ���仱�q���o�{��¤�m������O������$�v9V��蟥�ziJ[sTUUU���u��Q�!%2~}�����)��ڿВ��%''���.&51G�������ﯮ- �٠y�h��s$`���m4���3?.��N�;;���Ӻ�?G�S���M���`ֱH�Q�c����hٙ�Ws�{�6�9���"�JТ){���h	v�"]5g1kV��ud�+������:6UB;]���i�AJL��Oew35�ⴠ'BE�^��Z�j�#���:�^gjp������l�-T:/R+\ru���U�ѓ;�݃��N�(�k�)1�v%���u�9�E݅�趄8�sq`��m�ݠu�Ãct�ؗ][Qg��@E#�Ɖ��ie��5q�$�gms�����{��:}6�}oprպ��;��)&��+�m��Ƶk�������������7֯�����y��N���@;nb��@�j|�m���	U%PԹ�`c�l�興l̝��ݽVޝ�}�M��9si�,��4I�˯����hz�Z/mz��z�&�$����>�����;������(��$�����=�\����1��48�Qɠx�V���1 @�jΉw/�`V�T���m9k�6���-ڲgs6�۞�p��n�2�����}�����sx�����wM��٪l�ݯЗ䗤3���`����2G��z/z����~=)DC�ڰ=���?n��M���k"H�c�G1�w�M���?���|����@-�c�'�)���f���P�o_�����`o�5;��L��������BD<��Hn��z�P�+y?�7����ei`�tuU-v{x��Kr����g�7Gm�q�/x��q�]�^|Y����x{�a~�8��	��oד� 㚀��q�@^�*�!*S�.����w6��l��`s��7Ӛ��M��ra�54�PMM6����`c���ixQ�"&�Na
d$,0A+I
fb8�֕�!)_���3�^wz��r[f�Rt��n�����;�@}n}X�#sP�� 6̩�����4L����5�6l�}����_^����7^5�"Ȃ7��q-�Y�yC�K��7 �bĖL���:�w���q��GCK�8� �ߦ�}�M�mz}�4�F;'��6Fb�$���ͮ/�#�)����6��ls��/�����#"���h{k�5�6l�P���z�ͮ,�b��n[B�UL�USa�
}9�6۽V���r�����#��N��^�~�]�46�<l�N= ��`~���B���������������m�Ukv�K��D?��I�%1	��(�0zN���H;M�{W7maɹ��a�Hvv��GP8���J��-I%]���I^���BI}2����}�m�%��U'I̶�&��m�����ܢ!L�����ow��or�[�����m�-r���*���i��$��O�ԒW��<�fco�'�jI/����%˲�4$�i%�dN%�$��|�<I+�T�$�?m~x����m��m���2z��fn��i��^�m�n-I���J��z$����<�$�^��<�$�ް %vLJ�3Clҙ�J` "j d�Bd
�L���i�c@E�GB�0�����5ȉ�i~��F�!{�%�@BP��@hGI�.a8���*���Hp$��y�}�̵�oZ���m�� KCQ	k`�` -�l k^\�ӛ�y� �qc>K�ge8�AT���V0��D�z��`2�4�'��[t�4l�0.�Z%�'��l���g�װcv�/c3c7^�ٱ;p����ݫ�����ۅ��n��w�v�6���ێ��	�ضG-m�ӮWt������Vۜ�dw�<��=���i��0�[�ֆ7Z�G PV�U�d2TpO$�쭙g%����Ul�m���-l�&q@ i���k`m�j�<��r,���:�Y�C�-�h�Ng��=5Ut�1�
�óT�h�P �=R�i���I��9���� �`�y�6׭m������Y&� ���6�� �`�۰q�v��:S"��o0I 9m�ۦ;���Rm)��:��V���n�W��\eu����T�U*�@���pٶ���Ŵ�`T�lW.հ:�����n�6�4؅DKdm�[Z���l�ֱ�C�ܯ:"���{nYm�`Yi]��x��σp��[*յU�����3�G0�v2�6V��Q�*9j��n��*�[X�ؙ���	I�aa�G�F�kl�kn�����;q�:�
��'O8Bq�톹��.{�e�����ouE��&3����ab]�+[��i��\���>#���8tb�. ��{m�8n���`�8m�AtTa�R,��3m�ѭr8���7e\g�M���n��{n���C�*mŐ��uQӊPh#r��:�)��6�:���Ӟ)T�J�7��5��i�m�Dyj�V�`��`h�`i�ܽY\�=3�]:�M)�ɒtN�&�#7	��DM8��H�VJ��WK���ch�r���S]Js�g��e��x;jg(WB�7X<nͥ����9K�=�1¡��ɪz�ś�
mxv�� �2��dx�!�Z%�c��7)���{S�Ksm�3�_�����xv���(�|��g�S�=W���|��J��~3��{���-��W�]Έ���e�hټM>؝�g�7C7�1��q�y��;A�ڂtN��}X�K�y$^cmQԃ=08-+S��7;%�,�)j�Q�mA1��v�;�{el� �D���P�P�tGO8K�q\�����ٓs\n�EMt+�v��K�z�n:��ش:���M�	t����Nm�����GY��-�4�I�$�k	~��ߴ������+�`�c).�E��zzI.�rv�tn�v��Iy�֓Y���#	�&/I|����IWҵ�$�����%y�-I%r�IT~Y#q�#�Ē��kRI{�_3�orvӶ�O�g￡B�T�w:_��S2��d�q�I%����<I+��-I%_u~x�J��jI*�( ���89�:_|��=��'m��wz~���r�]���[�y�Ir�B,��!��&�J����$��bԒW�|�<I/y�-I%{���g��c��c��asv�&L+N�ݛ3g�u�]�����1�r��:�^�6����Iz�V�$���3�K�r��?b�e�ӻ��ͷϗH�*�T̍�i4֤����y癏����(�$����<I/_J֤�V�6�?\B	0ng���W>�����<I/_J֤����y�I^�5A���$H�$�}���Iz�V�$���3�K�r�RIy��*���"$n6�~x�Kޖ-J�o��$��������<I/x)-q�d;]e6sL(5׆5m[mW]��	sλ<�u�s�r��R�r��'��������%�9E�$��_�$���kRIW��ŗ��G1G3�K�r���f6�����Ē�g�Ԑ�����Is.�%Y	�S�-I$��g�$���kR��	B���4z������癙�w[�$����5Zq���m9'�$���n�m��������Z;m���������f���O1̊DjI.�|�<B^�Z�Iu�<�	{��5$����F��Qѣ�g�c7r�i���=��k����7k�Q�ՠ�%�5�W�cj�n�?����jI%׬�Ē���jI+z��x�W�t��<A �)ԒJ޳�KޗQ�$���<�$��*Z�K̼����ő7�x�^���I%��3�Kޒ��$�[g�$��:�ƔbbǎQ5R[o�"S;��_|�y�\;m��ww癙�o��bh���ډ�%���e	�������ff~yjX���d�#����%�9E�$�[g�$����RIu���Ē��f�'��e� N�p�C�b�m�)z��m�fSoj@�p�u�*c�u�y�Iz��5$��|�<I/y�-I	y�P�FD�1��G�%�����2����"fsj��m���������UE�4�Č�$��$�w_3�Kޒ��$�v��%���$�������͑$19���]d�-I$���<I/W]ǩ$���y�E�Q�,L�F<��$���ȩ��- �~����{������F[Vk��!4��cKs�]����L&ڕ:�����!m�V�A�ΧT�["�������W�H�"��% ͸u���=`H7f�f'+�"��m��I�muUm�C�ZM�;��֧�̇n�jq���#U���'hb��V�t�ŵv���\7�^���tǻ>i��� ��lVH&��!j3�dnӖ�	��œ��u�}���	�`L���B�r�K����i˛XXF�Q9/��,'�"������lȩ��- t�PP�w2�F�� �4�w4=}V�{m�����=YܕC$	Ĥ��[��9ɨ��]�Z9 =gU��hm�6� ���y�Jhm��<��Zz��FD)�	�M��D�*@y㖀#�PCK�fQ�u83��� =(K�f�pv7S��MnM�Y�촞�����p�-�s@�U��4;�4�ci���&��S.i|�w���%
aF(���ݭ�s6Ձ��j�BI�_j��ER&[[�V�m���js��ȩ;��ٷ-5I�9�UUXtC���X�T���Z nM@uL�d��k+����ݤ9 'c��9ɨ	��hޢ�ȦH�!�1�8�X�!���.��gl�8Ʈ���7>K�c�g0R㬢m�.�ƉĤ��Jh[f�}�s@�n��=ŕ�$Cm�19 �l�Jgf��{�Ձ����I6�rd@�"X�$�>���/[����~q�!���!d���b��R�	!�$���z!�E �?o���U��o�^w+��F�f$cD�4�]��V��ͫ�}��+ ��'M/�f�v�ܼͯ����'9�	�*@N빠y�U�,FF��Ik���*�ƹ�서6���Y���qp�*�+t���<�js��8�;�4?wa���Y1H�C�h�w4m��/t��[l�;+����L�Ɏ8����������n���l6I4H�%&h�S�_w��*��V�Q��(qȈIL����kX����3-ҙ��jt��T����?7�Jۖݞ�κ\��D��Ǟj�VQ�H�y�ϛ��Ժ3�n�6�v�d��� :8�� 95H�fmFbF4I3@���h�S@<�f�}�s@=��>p�Y5�bq7�^�7� yɨ	�*@sqR�X���Rj��N����L�~�V��ִ}빠_zS@�����R0X���wP�T����z��o� �I�g�������߿��v�h�ͼ���thc�[��:ڰx|X	x���:��6ݚ��um�ƓI�U�UC�0�8c�5��U�5f,��U.˷��a��]�l����;f(i�P��ܤ�/>��N��[۷fS��� :���z�Q�qҞrY��n�]�.㢺M��\��GX��ظ����t�{8�V76N���ݗ�Q���٭Q�Ѻ�ݽ��T��{�/�O����'/9Թ-�먬Y�v��V��=tn�^��sK7C���v�nm����H	�`�=�oް�ϖh/�����ۘ�#�nf�篪��͇���f���͵�g���@Ωj��n��S�guX{vՁ�fڰ=^�z�^��'���D��@�۶�{6Ձ��ٰ�I7��V�{�����2!ɚ�۹�z����m��۹�u� �sF$�LA�p�l����GFx3='77��蒔n����~�����ɮ3�73�-- ��f��)�{�]������i��yʯ=�w�P@���D**p��_���ok���j��'u�lK�u4M&ӡ�*��fV���j�I&����3��^�Z�SLt'A5Ef�� <�K@�j��[�| *�<Q��8F�hs�h�Ğgu|n���j��1sar����;V��sl4�fA[���v�%��W�Z8Dܷ��U��}g�v�5�@����$���7�@wH��Z ���^mM*e&IN���fV��&���V����l�<��W�(2dn��j��'uّ
�@bH�F����V�1&�df�9��0O�8�m`k���� ��!�͘�F���H������H`�a�B`�a��e�		!�03,&(f&��RHoq���7��8x��F����<�DH��
]���>;K��[z �䇤����6�F�Bnf�4FlDhT1U����$�L�@���!��|����'QHZ�!-IG�K�~��=�,ٻ?�h�w4�曙��DD'�_�; ����M�m��*���"�)6�t����� <�K@I�� 흴^*n�su��[�jq�*z{!���^<ݙsx�a�sv���o`��R�$��&�<�R�UCt)�5C�v��j�$���=��3;���Nk���y�NN���RSEnm :g�Z �I�x�;�T�����Dj&�Q9"��z��߳�{�����~	�����ż�������JɊdI����{�s��y%�=}& :VJ3&Vq˰��J���zK3��.�4���.'�d�e�v��7?���}�-�k�u���s�H<������@$��*�a5@�3K�<��o�g�wM��;���ٶ��!Cg=Z��m7I�SD�MT��z�d�?&��֬>����cX�@j)&�����z�h+k�=�4=î���i��9������I���{���LP��/���������yw���٩嵆cu�9�lJ1�Ճ��'���i�`H�=�5�h��m��W�S�i�7#����.I]gT�U'T�h���\%
� �6�ڪ�����˔�d�v�.�W'P��xh�K�=�W�s��':x�}ų�v;^��-�2n'vmspl�wav�<�hݐ����d��n�m Lu���/5^9J��Pe����N��|>�a��.wg.�eV��l�h4g�`բ<9�=$�6�izisk3!���+s�M@7�Z���ut�.�5i()"�=�4Ϫ�=���}v���eM+&)�& '&�[� ;�T���b �Px\�h�q�Xѓ#p�=����mz���Jh�o�������F�x���t�����*@z���m�aw==��8��us�c�>^X��QۃƘ1ێ���L��v�n8�����ǽ�V�V���k�>`vwU��D��ҥ:�ML�*��̭/a�  �I�p�!C�n��w�*����*����<�9W���c�R-�m��I5 wI���@;� @ܽ�S!54UM+~�� ���9����w4ظ��Q6%�= �ޚ��Z�"��Ɉ~u�.au��7dի��1�."vʔm�ݫ��*�`n[WY��;	����;l}�������R����&�=0�,/w�0����@wH� yɨ�M@{Ϫ�z���l�COpD��� {>�P��F~���:�y�Z��H��Y2E��$�=�4y�Z��s@<�f��5lb	1F�jT���v脷7�_��`|�6lhtO
I���!""���(ˍ� �8I�h�˵|�\r�1ix�6�]mͣ�՛�����& =q�@s�-W�P�L�����f���^�ⶽ�}V���s@���mH�lJ9$z�����i��߿%m�s@�_�z���l��s�L�@��S�{���ʯ��w��~�
��"� 'a)	p�r�I�JiBb��)BeP�� ����"�hrPrtX@�R�a�5��6)�fb)��8D��*�~�٠w�]�
)���H7�빠~�����۽Vٵ���D(��n��֧�����Һ1�l#k;{nӷF:P6.�����9�a!9'��3Q���
9������ ��@y͂��H�aY.�d�1�br- �z�β�����>�}��#ۃ��$� m�<�(��{Z����&�#��nٹXf�n�� =T��b �9�즁U��Pi2G3@�[^�}�ڰ36��>�m��Q�BD(DA��O<i�۩���Tҙ&����NӨ,��ʕ�q��՝-��{v�{���;�и��8ۅ�A	����z��dl�y�.��5�nUsa���vP���F�*�j�ճ@VΉ�S�Yi���)]��;uJL�L�d�tA���v�zv�^�;�9뗷@�6i	�{ql�$�%��j }�=y���a4n�M��.�B�I�u�ß	ۛ�e̐�69�"�]�W�^d�m���J�[<3��{q��.���mYp]^nx���s��nL@tj��Q��1� '&��YM�z�h����@��u �8�,�3D� :ܘ�#sP�� {۪J:�S�C(u4�興M���V��jǰ@N�R:�ta.�����ܼ����@8�T�vh�P24�y"�(�md�����;uR�f�9��<،�z�¢�=B�<���%�^��4��@�Қ[w4�Y�m��FK
q1H���n�U~����s���!m�$4D�f�u�4�l�:��@�n��;T��L��%#rM rM@9�Z� �_��M��s.�RL2dq RI�{�S@����<�vlٛVDD/v�9:d��UK}��P�1�XVT.�@��>/X2������g[�P� �`�E��1G ����9[1 ssP͂ ����)*�m��f��mx}� �j��@>�R�>YS�C`�ۏ@=����/6�6���Ν2$9�d���=����z�W�y�U;xdeK�L�X~I'��Ł��j�ǻ�`��@��#7�$Q�#���[���3�����i`}���j�$�%����!����5Rk�<��/7÷nYƣ��&@��4)7}�����@��`�}"���rfYR�L�ꉚ� ����BI$ٽ�Ł��j�37j��l햵��UEJu4�nf���� H� 9&��5}|جH�~�p�=��� �n�U���P	�	C���V(J#a#�w����?�j쩚M=�����T�;��9�@wH��`b玑d�1,i��"4�2+WB�j�<��`|�s�5gN7-�M79v��ԇT� ��ٵ���n���a�{�����O:hTʗ,���?�z����V��̀g�j�&�z��L��6���IUE���j���ٳ�M���`f�q`c��-neT��S���V�<�� ��ٵ���͵`|�OV�q��Jdn= ��h���:��*�>�uʰ��B�}� q۠ۦ�'�(__���@=1 �� �������n��4��������"�)-�,��x[�SOO�wl"���!p<�.��:o�=��7�ս|1�Ϭ,v�8�%�\����f�^��!����Ŏm_�L$�=#8r��b��|�#�F��ٳZX�s#`o��}rz1�m(�5��Md�8@́��z&���&�H� &+	2O_���&B�m�����WK,�lv�X*L��km�  -�6m�h0�yq�2�+;u�n�or�f�e'��P5
2�I���)P�&�`ذm���W`�t�\m�u��̈́H�QƮe8�N�ʔ[���;u�t �Ǳ�8��9RՎưq�WV�v��[&����V:�5�O[i�\z�w, Wm��m��h�]o=�Q�k���d��E�V54�F�蚥砚����i`Թ�6��X�-UP�\�++J��@ ��]l���^սtUj�5��x���nWf�r[+�t��Uq�"}�Ba25,�R�]�8B	3�����yӑ%�
U��P�ٵ��x2 ���Ŧ{E��Z�Fy�j�g T�f�X m�Y�cY,f	�m�hI5q�E\�쭤Z�j����%���
�U�h�6^�j]��ƭ�k����ܒ��UUR��,��]U)�J��*�U
ҵR�f�jK��&�@zv�c���횢m�j��j�WJ�d&V��ܛm\�[7l�8<����m
�J������g��OJ5ʶ��v�ر�d�^ISt˶k[# *��f�����Q� i�m�[l����8���Mǭ�l�dM�\t�F1���4�n�8Ƕ]l��=���Cq��h�3����'VS!�s3ڌ�:�Vɟ6�����M�x� ,N1ą�ݶ���[p\�vr�bB�s�6ZyR#���K�-��WJ�8�BC���9$܎Y�F"�^d�vN�b��2��乻V�X�;<f��ݮ��!Ud��h�l�m�N�4� UNRڗ�N$.��u��'g��ٻ;�N��z���� K<�l�ûl���[S�H�V��lXN�=i��p-Ǳ�Η;�� �v���ڐ�|��4v�y�KVm旝�F�۞ciKr����m`#\� �z�1��V�=��]ك[AE2�l�m�m��F�f��`{m&�Ә�e��8�y��P> 4�)���q >]�P�Uv(��{��󻻧www_Ϸ��#-���lT���g:��ڳ�Ԥ����b�Pm�BVE���U�Y��6�\�lY6��K�m,�l��qL��F]�B�eSsm�-e�m�D]BS�P
���E�i���M�t�[RIˎ봋<���q�j���{yoS��x��rm��HU�%׋n'P�[a�.�6����͒cl�<e1�[C�X�����}�{�G��P�$ѡF{8�*����k���jstz����λZ$���"^{:��(�)�u�M�ֿ�<@_��@���/�@�s��L��@�Қ��� �M@s��%�����F��ݛ����w>��j�� M������LCTR�e&���&�;��s��@wH�����M3^�m���嗻��� �EH�& �f���T�M�2A�M"���E��];F��n���κk��q͓l�*ļg�`�R&�7"�:���=Vנzϳ<A����ƻ��X��K)���+����R��?~�SP�& qR�\�i`�bbS#q��W�r���]�����Z��29"n=���z�h��@�z���4��I����7��[��r�� ������ۄ���o�l1n�=�G�RҳGp�ր6�9�.�X���πR'��L��9DQ��W�|���Vl��>a��`�e����U*�������@;�bt��䘀���#chRM�������|��C*���`>g3^w\��l�-��d��F��r-�~ǹ��1�t���V�k���𹡼&A�Aɚ��z���mz�۹�y�K򹂒()�<ngR5&�Ո��[���pX�sn�Ԝ��A��u�F&%27�{�@��j�=�����@�
�9$�&�)%��N뾈I�;zՁ�;��3۵`o��\�b�?�qh޻���^�>�P�%�7,�唒.�t�4��_�;��3۵`{�ZXBI}�Fff<������4�rH�<��2!�� }&�=&���|� :geR1�'�A@@���LAP����=�����E�o7D�/;H=v���M�t� :8���b }&�$��d��Fۄnf�{���ޯ@/�����,�ehX�dk"�M�\��5 ܊�T�vL�f7#�1)���޳@�s@�͵a�!$�OwM��ԛ�uE�V�Y�y��nEH�T��b\s}$����-!�I-qjkY��ƹ���`�b�tm�^���#]����	��B����y#��;u��U5[#��qmT;���)=��U'�����T
t]:�����Я*�]h� ��І��6�N�D�5@����`�\ۃ[��Y��W��l�[���7ce�K`QD�6��Y�b:I�tD��^�"r5�-�*�j�����^n��Î]�+��&�u�L��]l\Cg��ʍ�"�^�jz�P�5ɘ�ꦤ�O� :䘀��r*@��l٩�H�P���_}��*�^���s@����bA�G�F���<kw_��@6��*@z䘀�F�TXD(	�$4�w4z�h�k�-�M�t1Oɶ�� $qR����`��M��������w��c�% �7&��Uh-�-�.�e}j��vT8�&��]nM��NM^��׀v�؀��Ht� $qR���1㑉�L�G�[�sO3?�T�L� ����w�ʻ�]���W�{^UAFD��M

L@wM�G :�L@H�Lw�dX�Yѓp�-빠z���z�h{e4�mFI�&�LI(F���>��*@{��#���[��Oj7I��A��r������ݞݦ۪�A�l7��Wl�Xv��	�����@H�G�@H����q��
9���=�)�[�s@��@��4���k�M�r����9W��{�Xz���r�����"&�H��,�,=��ɑ�h�5&h���z�h^��-빠z�h�6$�X�Jdr4�*@z=�I �����	�Â�Y�͚9��W]���i5���Dn��
w[h�N�Hs�Zv��`��EH|� ${Lx�Q&$@�2cn�w7�H��@-�M�|@�/�L1=�$�36���؀���@H�;-�?&��d����>�@��)�}���>��M%�ٰ>�ʕ3�L$m�n����67 :��@>�����o�{~j��n�^�ŕ��w.�$�7"Q�ָx�bқ.鷶�Z݅�۽ͤ�EH�s���UW�����V��pL�Q$��T�?n���t��� %�	��W��Yz]�nf����EHt���z���
�h�cF$��<�U =�*@;�1��b�Y�,ݻ4/h����@{�T�w�b���������rG	?Ll�<������F�WLDڵ��]#�+���3�<�i���g��@���p����� ��4�HCEJ�-��#H���X,�˶ЫA�h�=�н+���A%�>�8�C���{q� ܻ\V]��{K�x�k��Y.
���ȧۅZ���m�7b؋��2X{'5<�p���q�tꥷ�Y8���"��W�Iݻ������O���:O������u�"�Ɠf!4p'���=�9�]�sP������t:�Z翿����l�nm��K���V��*��&��R��M�癳`}����vՁ�ٳ}	&�jږO9�"JH����~��<�w4^�z�����Ȧ���m�F�h슐��@u�1��_BVX	��1�,RL�9{���W�_z�hz�h綵�D�q�H�|�/,�t�4��K��[،p�b��sqv���bN<�	L�Ǡr�^��빠u빠r���/:,�&�$�ca����6��BJU	%)*��m������
����0�I��*@;�1 �9�� :ݸ[�+����m�MR�y�6�f́�m��<�w4���X�2,��I�[s�*@yȩ�"�u@*G�n!��X�K���=T��.��n:�i�9�-�,�q��sn��zx�46Z~�EH9 ;�T��nbJ
;)��@�j%�ηs@��w4Wuz�۹�z��eI!��<y�`{۶�<͛%zi�!T(�%I�CX����у+�O�RRh� \����b,,0`Ms��HKx�&8�}�1�'��̳

j3_A��ؔ�h�D�82'�.�;��_6�� >�+꧈���⫬��˕{�{Õ}���m'E�$�h���}������=����|&�)#DOMƀ�s���*@z�L@s����..�c#�(�vk�,���\�ù����>|��v���#�g�k����s���&~����߄*��Q9�f�&��� �nh.�� 9�� F�e�Q�V��e�H[��*@w8��"��]���4L�87#����{�}�h�p�^��xr���B���"�ه�|��@�*)��BM��b��H� =}& :8� �|�C�Uɳd�cfHG��4eƎƐ��v=s�@�nܳ��k�*q�z�s�E�i �EH[s������F�q�PQ����x��߱#������Z�3۶��$�6oN�-�uSe9S ��M������3mY�!$�����o�@���Zx�(	�q��*@>�R m�@u�1 �[�w�����j�׀�� ��\u�^����?ߞN_��E$�
D��Ӛ�P�;���7'�+�U�%�G$��N���g6���6��ӵ�6�2j���F�m����P�	G�H weeW-�t4S��0R�;9�)���^2N�+�6�t�8ct:�V�6����Ͳ��q�'���%*+����M��K\���z�׷RFSv)vJ71�t>��7V\lc���d�jҺl��+v(W�ӻl�b!%�U7`)��tM:U#mH��r��Ů�Q8��PY!y4�ڹw�!�$�V1���<�o�]�F�׀9ϵ���������s@��}��4`�d���@������H�*@���.^���噷��h�T�}"�:M@{_U�r�(cɌ`�,RL��ffU��ޤ���@t{n*@K9�DƜyF6�h�٠w�~<�~��;޻��H&V�S �{8�͚Wr��<v�u�ktC��G���>K���H6B7<LnM�Қ{6��P�a������'9�jI��Q.h�3۶�RP�
!G�T~H���j�/_����M��r���)�^�2d���noZ��6��oݵŁ��j�=��6��BsD��+P�K�����`?��@>�R���6��+kv�p��@z=���T�:��W�S�6 Ф��Ib�$5�\q���Kv���8������nnH���|��_h�I��I �_�4��� ��hޔ�=^��Ɩ"�����j�%	Bl���`gmq`n�ھ�ICg34����L*�L�+�wM���}�~>d�jR�L����HZ��&(���.��}s޵`o��X�CjvU��䩩��䟻o�7�Ձ�ݵ`y���{]	�&� ӆ��s@}"��& :=�����g�Y�r�n
,X��e)ܗ(qr�Pcu�h�E.�uDJ`�t��e��hU-�/�߮�rj��$T�9�����kM�h�:�`���"6{���3��X��W�	��o[�9d�iU9�3wP�� t�P�*@ɨ	N��P�Irɧ3T�9$�wuX���*���|�C�J��c�)���3��Z.((�DE$@wH� I&�;�K@I�t�c��UہtX�ݴ�vgj����Q��i�Mͻ[�N8�wND��XUyz7+��$�P�%�	$�t��=�"dȌ��M�]�@-�h�n�[l�*���
cD�ёb����ڰ3۶�脡&��t�Ӽ��oV���*�rX*nf��7;�X�vll��$�}��`���*��%���TҰ�ڰ;:������_{���^��?H8���t��i�����e,l$]#F^�x��X�:F�k��܍[��k�{g�w���-Y�;<��2O<�Ξ��UV2AO���۬�к�؂)�Kb���1L�DRW
�(l�%�(����n7��ve��y3v��:��0s�$mӈ^v.y�C�ۖj��i��tq=��[v۫q�[�Cr�Cfo<V۫'W���n���9�o�mٵ�n;Y������{���Ȏێ��n�=� ���N��s&���\���Z82��stOb��95���nZ�o���]�n�Ձ�ݵ�%0���`w#��27,�tꝀn���D$ٹ=�����`{g5�~�;4��-���{��}�Z\�1�@ɨ	g�X	����ȌrE�Uֽ��� ����v���I�� dx����9h���}�Z �P��:y��A��V�Z�ε�jn����@���pD�v���Ί�q	�	ۢ�3m ssP�K@rj��@fKz���wS3l���W�gOs�_/�P���߶l�+K �f��J!(l=��s�H��Ƀ�h���@�v� �����Z�`:����܏@����=��`}���9DBOӽ�`}�(	���D�n�u�����ń������a�t���A4Y�3�q�WZ�d�0�ge���fԝ��ݔ�ɇt���N��FF��o���� =nL@6�^���;$��W$?7�܆���P}�q����e4��cx�+�@��=��75U_�W�U��o�_I�	}(��MF�,�	�@=�@��M�ֽ����ҹ!���CQ��|����
�{��3���=��Z�]#��I����(�ٓG���Dٖ���;A�i���aÞΆX�2F�mm� =}& :=���H�a�^�*�lJd��nG�{zS@�ٶ��֖�۳|�!���'<ɔ��"��@��@�l����נ{zS@���EfLBǑ6�4��X�ݫە��B�J%BQ�|�v�ƀ}��FbxIɑ܆�y�@���O���@���h�c�i�8M6�:pj;3A1�1^�K�mDMy�.�ׄ�,� <M��dpj94k�}����N�舄�`{;���ѫ��I-��Y6��=��4�ڴ�m���ZsJ���o'��ȌOd<���@z�L@t�-������e^�w���f�=}& :H����٠^�PlHS$Ncr=�J ;�� H�=}& =N�~��U~��i�_l<����n�1 ��hx����Ù��X�Xd���Hf�.�1t���c��Mi��qJA�3�0l0ȱt�J�һ��q�TI]��#�O�^L6d��d�)�8��<���6$:�,W)���,Zh��
߾���Zս\l��t�F�ۣF   -ɶٶX`l�H\ �|6}l̛g!���)�7]�P��+R�G6�ӎ�T��JdUg�Q�76PaL�n#+��'0n�üݸ�lq�<���
l���ۮ�����'@��A��s�wP���g�1�x'��W�zv��Y,dK��3�\���W[?�����?-�&�tz����K��	��-����>��j��8`bj�i[��'Ӑ��>,H֙^	��l&��5l�l�h  �7g�� ��	vvUj�^G-���[�>�衷:\aӌ�ڦeQ�:��x��[g/[EȲKlc	YկWf�	� BٮlH��-���۰i,�� 	;!�Ky	Qm �`N�m�  5V �}M��sW	��Lm/5K���3K˲��m�b喊P�@�W���"6�)�3�yr4ʵUUR��*�U]+$��J��-Q��j�Tv]ud�sU ���2�s�Tq�k ��\mn�]�e��9��S��V��STQ6� -�K-�&S��(8��\�7������;c&�v&�:%��Y��UX�[$�P��嬛hq�-��d{Z�,���GOT����Xz��J��:�튪Fu�՞VM�x2]��b���v�{�8r�k��K�����v8n��!�sKĂz�tm1��O`���`�^//�UxZԷ�t޶�\Rj�����4�X��l�'��yڲcn�×6�i�+E�!N\�Ej�{l@��x�ы4hvN<r���]��&�vʃ�-+̝dU�U���4��ײ:���ܺmdOj���'�^���U��Re7�m�y�����Tj��z��kLPm���XW��ܢ��g�X��I%$su�s��fa���/������&�3�'=�����ݭ�<�H)�=Bmzb�d��K��]|=����e[Kj�:�,��d��N20W>�Ɋ�������ѥ|PC����/UM��D8lx�ͩ�9{����f���[)Rg�Nz�G�(Q-�X���j�u뵕�tnot8r�E*�d0����ʕ+4�7j�"i\3�U3F��K��`�.K��UmTnӍNU��"�H��ј����L���B���'�9��ٷ��^�ij����iw��:�Y��3���}�n�zO9Y��m���@�t�܇6�[3a�ojݸ��X�[a�{�����͹�)�ۀt�hO�N��.�Re5{^��/M�W&t۰r�bD����nh�f�W��ޔ�=A�%Y��dR)3@-ͫ^ń�����͵�I6]�X����$RM�~������w4޳@��a��a�##�����*@9��&���,N0i�cȤr�����f�y�@�Қ���#xɟ�&���v�eUY�۱�;u�c��N�:�;q�m�O,�J���Q�v����/ w��V�۳`u�M�z�h���i�E�Ž�y���i	e��z'�}��{��7s�X�6��;T�m���*�ͬ��@G�}h� �j��f�nVDBh�jE�{�]� ��Ձ��u�t(���]������L���"mI���4=v��v��z�h�ֵI�7�rG2`(:y)[��F��y�:�.˃�ƴ'<f۫���8GCQ�M�]�@�]�@�޻��Q03���͐F����M:)UM;7+K�	(l�޵`��`}��z��ul�r�'!�{�]� �ͫ;��!*�d�;�mq`fK{��NA7�l��q���~�����Jhw]� ��-�p��db�h[s�~���<I� 㚀������y���J�6��Hֹm�3��ȵbNu��y�b�qn�\��u�X�q�n*@9�[sS��k� ��4;����_��@����:�����QX����d�H�5�nbG�@y����Ǆp�5	$�<��h����w�+�/<T_��w^w|�ϴPe"a�&H��:���{�Y�r�^��ՠ{ԉ1Tا� ͳ:�J�*�ˍGa�0����sv9�gϕ���М�m
c�ɑ<�C@=���9^�@�{k�:�����q�M٬�aSU_����(l̝�`omq`nmX�g2����jG�yϪ�:�ig(�M���5����V&��)�mm��^� {�&�	�_Z�p�atȰ��#��{�@$sP}& {�������7i�V�r�akjc$��ൠQ\��v���k�����F�������Ɨ���mٶb��ͶJ 4�U*ժ2��Sm���c�b�l��M칗�F�Wvy'm��������h\�#kFC�����v�,Q�㭚�<��mo�3����(֓���4�����=���8��0�j�M�y��\��v���ﻻ���O3�aT���6�Jq�<������7p��\��v�ۆw,�g!�123��Ɯ��}��h��4��}�4��."I��
���۳�CggW��V��W�	6f�-L����䪧56gW�M@�_I�W9�w�`ә��Hh��4�Y�z���tB�	�Ws�9�ܦXO�*K��3U� �O���bvIh�M@N�[nQߖ�Ո�)6r�_��|}��Xԃ�ɮ{Ws�!rh+u:ka�^�t����jv9h�5 NsP�1���xL��������ؐwu�{��<Vנ^�vĞ$���f��g�j�7ٵg興oϷ������=Y�*�����&	ɠ�Y�zۘ���1 y��Y�?]��+%Tˢ�����l��B^�ޟ�=��`�f��%[kXƿ(H$5�8�e_cA�h��E��D���w<gٺ�3<�������bd�z�����4����3�$��"$�9�4ԍ t�j� <��@�j����?�4S6,1I'�[~��<��h� |�P0��!i��FH �P$e��1C����� {�Y���d���!���nZ �P�5��s�R�M����
�����sv���@���Ś��Z��T�M�<$���#��H�q��8�u�ì�7�廉6��]��iNL���L$�@/�f�}�s@����$�`v�U��a�����J���X��W�6vN�9����mX"׉,���Hnf�}v�����@����v�ܑ,x�UNjl:!(O����3����͵a�'�@��qe~��?y�U�n���hO1��"�����-빠r�נUz���p�_#�hG�4�Ő�tO��ڡS���ڱp�J�kz��q-L��h�tЦ���~�߭X��6���oY���\�����!�s4}& �- tsP�T���U]��}�!�#�h�O� ������}}V�݆���4���; �fՁ��j��Nk��B�ӝ�`c�[ȑL�HԪM�U���j���- N�P�5 ��)���n�V�p�26�#j�v���ֺ��BN]�;Y��y��#"R;0k�(�;<F�{I,��6c��-���O)V��g�s��nv2���6�h
Vb/�}���[:�S,�%<nら��Wq��e������b1�ӹy�,m�v�I�^���������W���]�����Y�7�X,�ݚ홷MR�ROB�R,h�UT�U�v裍Ӵ�Q$�>,k��мfݭ��*<�5�1cd�,Oi��9ߖ�w�� �������y�CU%�7Mʹ �M@���EH	���"Bǎc�jI�޳@�ފ���s���	��.�w�A�]�����R���sP�5 Z��!HO�q���<���=�h{�h��s@Yl�S�5��1;����`خ����9�&���<{\<Z8�v�.������&L�F�~ {k��z��{Z��t�]�^a�TK�� �fը��Q�B��I�m���@<�٠x�{kLbS�<���@���I����sP��)�6�x�X���y]�@/�� ��4o]���r,iI�d�	�Ih���sPT���-�S�C�gTn��a����Gk�'cm��nq9z����ڴ�vΠֺ��Ȼ7u 6�:8��Z q�@J��q5>[����I�����v� ��hwY�Ֆ�X�H�8��H	� 8棊�ª��QT:�=�81�;M��H@�FI�e�%�����Q�O=vhgH�ј��L��fH��	@�dy���$>w��H���X[��+�4;4kF���JB�5��f$��8)� ����z����I	��X��������:ɢ�Ȅ)Rh	$��3b��WDLk�5��	 ,#�6>�l��&�W�p�xzFy��RziM$>����۰Y�LB��1�y��Lƍ��� LTͮ�@�浶&Z�N"/=���=�h�bCf��s�>��ѐp�,!2��1���m��Bd�'�h0٥"f�5��Ȅ�eA�H ��$��&HH��A4o	��*���6 �xz��5 �R�+@���T4^�x��}���z�h�׸��7�dȘG�&����;����͵a�"v����G���Iɠ���w4zS@-�4�*�֧�X<�sec����m�N+���#����ɻPHwF���m��~bǓrh�w4zR�������z�3��9�N[	����i#� �$sP�*�l�T�)�R�T�3N�כ�`�j��H��J�̻�3i�NE#��Y�ym��<���3��ߴ�`$��\��k�~=��~2���+�/U��*@zd��w�e�g�ڰ?BK3��MK��*e��#��:��۱��<�R�g���c��v���,[ɋ��!�9���>�h{��{��/�voZ�3]6%�t�S�&����7�
"6�}V��Ձ����=�I\4)#mŠw+47 'd����1��Բe]����+j�/u������ Gvh#���D�iNf�}v�癳`n=�=�j��QD"��~��hm&�8��@�H�����뮠��6"�.���yƍC�[��%Hg�QD�4�hݟ5R����6�E���G�!���t�e��E9�h��N�8�bXӖK]<+��	mѮ�w�q �/�7]��{kK[;�ZݧN8��x��:�Nn��W�8 ]nC���|gv�(Vd��;��ȍǷH�5��TM�&S�T�U'�%�	(j�ܟ̙��]��ca��2�S�c��@1�p���v��=un�l�	ڶ����c�ؖ�؀=�@w8�;$� �9Whi)�i��yyY�{�]���Z��^���9�Q|�cx'��Ż��*@N�- yɨ���"9U%#��C�h�j�:٠^�h��hz\P.Oɑ�f�95 z9��9���K@w~�t������1z�۰X���=i��	m��Z���p���|��;����7�������@G�Z �P��e6�$jU&榬ٛW�	y/�UW�V�s��&�G3P��k�Ȅ ܚ�j�/Y�^Vh{�h{�X�jb&I�5$���GsP�5;$���~��D0i��� {�_M �z�};��>�ڰ:;v��EL�)]�h�C셆��bR�lDs�lttv�n�N��j{&7���=��'���' }����ڴ��h���ׇ�ŉH�7,�77P�L@����j ���H�&(��d�ؤ�@/�f�y߳��A�#�8*iT?י���� �_�z�jȋ�'�4) ӓ@<��8�/�����_�R�VS�5*�r�{6Ձ�DB����?��@<���.u�j�2G0R	8�ul�Է#s������Й������ŷ�ȢȡX<m,��_]�@�^�@<���;޻���b�26�dy#���\s����*@K�1 wuď��y��&��/+4o]����� ���o�ķ0/B��U���V�ń���a�D)DCJ�R�%L;4�'sT|�����`�x��xG3@���s� GsP�*@~��U�}_�n�?�8�5���'3%G.�jF�\���=�4N3��Jt9�W�9�<���\�K��~3�� �q�X����s��>ϾY�CM
I$��/+4}ݵ`k�����w�BIBM�ls7�� X�bMI�^�����k�h^VhR���%���Ĝ����@9�}h�sP$T��u�f5Y2<�$q��ՠ�@�۹�z�W�\��n`�����c�c����s//S��v����u�_V{&���#�y3ƞۓp�YՒ�Y8�rECQk�[Ce�*T��ej���3Y�b22�,*Ұ�'C����f����$�UWZ@�v�-�V]�r�#{U��9�����<絬��0��/gyݪ�����v���t;�x��k݌m�l�pN��a���=���yXۓ��d�&p�(�\�Ȉ�_Ң�xg����JN��϶�JZ���V�e�]�xK`h|U�s�|�[�h�Ll�d�4��2G�ߗ��=� :c���Z�%^�f%���������}�Lr��`�$wf�u����n!�������:\��EH��Zfn��mfe� ;��@��@{�T���4�VDX6���G"�-,�>���3f���5��˸��ʙD�/�9vvôF�ŋvS��y���d/iݸg+��H�L7U 5L�JfJ���wZ�:ۘ���- zBj[
��j�D���sJ���ټV�(�	"!%0�k�V�w��h��h�/!;�I1L��z��4�K4�]���^�^���8�1I ��js��m�@N{LJ�+��K.������ϕ :ۘ���奚{R �yrG��!m�Î_�;G�BD���uƞ+��&���\�+u��d���(�(�����_zS@<�Y�y���M��N4G1F��h�`�<�5�R m�@:��!�m4)"IǠu,�:������y$��ޫ����ǐd�#Ba1�I�u빠�f���z�R��JX�J~SI	��;�k���X{^Ձ�ݵ`$�Gw���w%�L��c٥^�n����g��sk�m��n���2�Y�\�:��w|���b q��$��#sP�&6��&�qh^Vhu� F�:d���ʚV����؃I��~�h�U�{]�@�u�����;���G�RM�uzW����ٰlkM_ғ���7����(ҎM����ծ�3sj�=�ڰ?��r�4��z�X�n�Kxܝ�+-�í������c�=�ܖ��ȖH�lx�B�$�~���= ���5 �9��?ź'�.�K�sS`��|�l37����s�>~�^���\h�?)��rh{�h{k�<^ҽ �l�;u�P�s��4
��@�{J���@<�@<�(%?7�2NE#�<^�]��!)�� n���2l�
"!(W��AW��EPU��EPU�AW��U_�T�T� ��D(E bQ@E h@ZQ@�@�TUE�"�*��"�*�Ȋ���EPU�AW�EPU��AW��U_�T�EPU��AW��U_TU_��PVI��x��@ٷ�@�����d/����� �[=;Ԋ�Q�+��>[-�{     �$(| � �>o�}m�yn״���Uw3�x=�����[yܹ��3< 3��|��������Ч���{����6�m�[����� �N���v�+s���k[��玻6��=�����{�M4�m��l�M�>��| ,��n�eү)�%�Τ�޶��s޺�wgy�J�{��Q�v���V�w��Sͪ��7U��uU�y��n�  
   R���)#�0&&M�  �#�SƤF��        ��U*T�2i��#a2bi��`�Р��H       ��I��SM�&��ď�=G�<��I��"D)E1#�� ���� �����J���~�P"�"` y����b��; Y�������h�@M�E���牠U@x��;�R
�1g��՜畷e�¦/����$�I$�I$��˻����	$�I ����Iw$�]ܡ$�I$�I$�I$�ċ��KRH�� (� `�$������I$�I$����I-����H$�I$�I$�	$�I$U��]�	$���I$�I$��I$�I$���P�I,NRN�K�I:I$�$�I$���J�N�I,H��I$RI*I)I$�$�{�;�gwF�w+���~��Z�\���ܔ<s�I%��%I$�KQI$�I$�����I$�JI+A$�I$���J�I$�I$����I$�I$��wv�3֍Z���VP������� /������@7�߀����Yկ�o�]^q(��BÅ�4���x�x8oVSa���L�����[��w�.�i'3gVw8EH�����6lì5�ҹ�卜�ÁYɲ�12�k�0{������D���� f�;Ԑ�|�Au&���[|��0;�}����D�4�1oI5��M"V�q:�x�n;�#ȯ �J$�if�n���1NԺ���ݖl��ؘ��Gr�9qE��n.���]�'�}w
�~�BE`���7�Y�(��$�`� b$2�)�J�MLc��` �HB�0��IR�� K	��
���[�L7�[�ﺭ¤�T��^p��"D:n!E����E��!�A
`PD�(�J�c4��#&�DX��aDa�r���l�&M;��1�L���$-�x�;K���,�����&�{
�e�8%0�%7$j`�3�L�2HB$�|�M���D!�[Iʖ��!L��=`�I�2#�&�%�nе�'�O�C���˒]���*�ZYV�@�
]�y7��<nm�R�HB	w�����#�x!w��9��hI���%|^j�5���R� x�Vf�,���قs2,���F��i=�J�v�we�jVV�o���fq�׺㋽����kz�[z�adKoW
����i�9��Z�h��6��D�5�j�h�|�.M��u�4s͌]R��N"k� {��!��G����8�#\\;��`b��%P�J�����Yۘ]���hM�F��T�[�B�x4�#��[���Jn1O2�%��	��nvd2�:5fD�A
iIy˾�%���������%Wi�NI�U^y��m��|Ѕ���2G�.q�֓��<}���Uw&�7Ñ�e3zRwE�sY��3�ř�/%���NM�PHF.����N�G�;"�w��]�.�x#���5�l2GUW�<�ս]�v��W���QĪҐ���}]8��O}&nu,�ʛ~x���z� ��n���3��s�������\�x'� L�A�3��[Q�u�ڡu#DmD0J3N��Q��B�9���y��ʲz)f,�9^�����8���>����|*�eۓ�q���A���[���8�vОR�����#�ɐ�FT	�;�K&˦�4�7���Lu�&wa�s���#�V;EP���i����l���L/������|������9�r�4&��A$�������_�g�d��d�_�~�P~v�Ͽ�r~�����9U�UUUUUUUUU\�j\v�l�k�nBxb��J�c���H�m��3M�n(�ڲ��,���U*v:tc�����bO���w}��a.A���[d�_?)�������ֳ���}�}��{]�r �+t���8�2��s��u#ц��Q�k�͆ݖ���ڥ���.3��55+�ۋ�\6Ę�.������h�ɎM�����Λ~7�����,�3���N��f�����vg�l5ˌ� Ş�"�y81r�!{ua��ן���k͜ܜ�f��تxH�g����]��'�X�i��UUUU[�UT��N�UUS�]��3��1��۷u����O[t!��\��m����F���eݓ9���W��j��{6�6h�P���JEj��������U].&ej�^���U t������h6 ���6��\C���O-V�yA=b��u��m�xz�UD��7\m�k�Jn݁A���s�W����vk����տ��|�R��S�iTY�= Z������x%@S����K��a��[�mU[Y�۰6%X
ڹV����¡�<Y�qӳ�k������m]�>{-ː��M�c���L��]T���5�k�)Nq�bKKs~��$Ʊ;EN/%D�a%�E����!��g�tv��7o�vʭ�W��ڪڪ�*�����j����tUR�*�UUUUV�T�UUTUJ��UUUUUTUWS�*������     �   �$�        �*������*��
�5UUW!f����U��Vꮦ�UR�X[[�6䖶��R�u5.%��n����4�� �J8�D�D�m������ڪ�����UU���檪��j���HUUUU��UUV�@)r�UUUUU[V�UTn�QQ��=[�!��a!�st�����M�����'�1O����N�-�4�{Nݎ�[��&iȤ-q+Fԍ�2-#G���,���K�>�ܶAQ�倢'c��M(�;��.�7J����SST�DDADTETTREQDY�U,EA���T�U%UDQ4S1DEfcQPLQ���PfaUϘÒeA	�eM�Uf9�2�3�(��2)0��?�UJ�R�E*�REQQUUQQQQQUQQQQQQTEDTEDT                        QUUUUUUUUUUUUULQUB1�B��C���@��@���Q͚� �I8Pq�Ⱥ��%��Z6h$�@k(����SHW�e���6f�4�ik�8:����L��A���f@���i6�2 ��810p�/u؋C*p6�Q�h�ap�����:j�4wW'%d�&)�utSoTxI�2,bKN�;�S
�;����N\mӗ�����BF�q��F�J�)�����s�p���LSZ8�&{��h��'�phJ ap���UQ�e6��\�k* ��a�u�:4��,B�o�aK��7k%UQUUUUT    �              lp    n��   ��        �    p                    l  �  l              p     ~�C��� �$�`�8����Dr'�I'wIR7wwj�P��%
�.��~a�J�	�*��!�]�!wy���2�5�!̸<�����q�2��m��u�����5 [�r�������ڝ��b�e%��t�h�O;l^݉�m����7]����~�	q��i7\@sv,�qb�m~C������W���2=Q�
�����8@u =���t��٠ٸ��vt��ݍ�#��@�7.՜N��]��λCnp����j>ѽ��,~��Ei�>��4o,�ξy�v�*��[mU-*�UJʡ A��Ȉ�*Sp��6�ۭ�9�Y�q��mLu�C��w���t*)
�Ω��Į�KR�Q�2��_b�F����m�k�C#���;E�:���fl�)��P���fD݅�)��(F�6��?�WҠ2�������ǋq,M	b���*�G#NF�ܟ��s��{��H�w�֦�7̳�L6���ç<^N�~%��݈�[`7j$��rK�b���o;;0���e�s���������<�"q��v��鴳�<�_U(<	�f%�ך�p/q�jW{�텀��640ز��2`c�˪ؘ{��/3��+[v0��Ki�kN�]��`o}9#K�1R.G��`S`�9��;2fOW1x���T�7i���g��Ԩ����HhH#2&2�<��SFbJ�����{�!�Ͳ���Q���a��f �^�{B/>\
��h��V͎�Eڢ����q�n�JH>t�ZKic;�.=��GU��1M'�3N^Fm����fߛt�e$%$�E��wI%�s�5�0 cc��`���02��kyw�$����mmbSo�"����X����E��pΫ�b��	H��<U�06����z�I�5e-hWk�)��]�2L���;�􋻇�u`;�5�@����oWX0����FK�J���y�S��J��ؗR�T�\�"4��6��fO�lj�Xݭ�:V&J; �*�:5(��C��5t��`d��kQP�-B��*hf�񛺪��9�fˉ# o��=��{���� ˾З�hVJ� n����{��段��.�����*p:�/m?Tؚ} "���Q�VhDEe�q{�ŝ�]v�jE��i��"#4���K�#������vru���uf���% �X1@�
��B��lB|z���`��W�ɐ����&p���^?��4��I�"�x�|���z�ikh���5�H�Nw���kn��W�n�r������.�ja��7�ٯ˯� ׶�Hj%š�Fkս���T��N�$\�[zW5�ևQ~������47��P˚a���
v7���ш�y�y��Ɣ}��^k�l����g��&�jO>�M�L[<ЮO���¹T�������y���0��5�\��q�j<�nh�`߻׹��vP'#����i�ህ�X�{�2a76�D9T&aX��֏��?P��z��^�xЛ%���VJe�d��"�3����iV��m�A 5n����u7�n�IQ��K�6����t��O�����\�s��@��~��+����ME|�}�Y@lO{J(��v�4� �W[ֽ�TQv�\�Pu�Ts7��y^�/�Uuv����,sً>�{�,fe�کnl0�� sP��Ra�=���/�>��mjV����NT�_�W{g�5l%�'ƵǠ���	�Q.o3KR���qjL��3߾�<�o�k�g_o땉��Z!8Z�9�������s��^�W�ʜ��0�³7ŭ-}�ޅ"�*%���S֗z��>k��p���n��/�{����㶌��3���~��FC���=_S����ǯ��X<+6u��M�r\�,p#N�M���Եs�ܟfִ���x��X�
����]��R�s�tV4�o	��־����O��"o���ov���]"�[3nw�U�9����$�+�e߭�2X:��Z��I�Z���*��R18�&��4���<�j7�N!�o�UL%�+[�����_`�x��5Cy��x�sʵ�׹^[�"ImD��Mh�is��w�]w��2!�7O�1�C�w�m^`�}�=��U9nw���� �*p�Bw��6d0f�p����ΠxvXF$Zu%J7��s�𝘾�9fz_��,H�� �A�C��uܻ
:��p����P����tW%OĖvo��Ѯ�h��ϙ�d�=�����J۹��,�P>��( p.gwD7�L/R��S1%���m�ae�!\�/_K޿7v��U���Q�5��PL���k}��/��$�����?zy#���U�}�IlD$���ݥݨ���7w���p$�ffc!ZDa x9��Ι���&ɋ	!5Ⴡ�% a3�'-�˹�����1K�e*�@ D��tb�P(�#O𐌮5���`������C����t����g��9�Y�gng�[��i)�����fWs���7Y�Tl� 5��k�pv	�v�l[1u-������+���*T��ڣZi�+h���`�<� _�^ݝ�|�������uJ�PT-T��*���N�F��غ����"��b��u��:�}	�:+���ƥ������������/�%�Ĉ2�q�0q��M)`9�*�h��H���Vq�[XZ�L�������쳎�8o������F�jw��x�{$�$�����4P%c�1i-k��mfK64�"�Rm:�T?lq�A������P�eH����;���Y�ș�F��QS��\�fj�qZF8<;��y��0ş��Y�@�Q���}_jS��d��ơ�p｜Fַ�\������E$�d�KW3�޽�Bk����i s���1�g��u�!�� �M��.�ǽ����z�s�=�{�L�4%]�<�;~T��$D�ys��z��ֺ)Ӊ������j�0`fTxe�l��bG0� |Cf�]C�^	�<��2HJ(��n����ww�IKInO{��Ue�o$Y�~�݆s-����4X���>K7���ľ����Ed���g��j��ā�1I��t�J�WP�.ͿC���|�_��kS�,�L(�>�Qf,��[���s7�_������]��|���31D�1  P�1<�f�pE]�Dy����J��$�Y$ı��%�Y�1z$�Vk�dJ�����6l��W�mD4D�LEt�[�6@55s�D3h\w�K2��y,"� ���U�T�s =�HzK]=��QGB���
�sIkǤ�D����h9��!��b�5Ȗ\y��&�$�8��!#j:�_<�`{�A���)�L�qq1�����fH����� ��~�8V��Ӥ�$�¡$��A�E���ss�yfwv�pr�sE�+�6n�j+���� �4���;����������:��@����Ud�-1�ř�bYLK.{���Q�"�c����eq9ND�V"b �y���QP��7�A�5�<�A�[�X7�E�G��բ�k��> �^WGĠ�s3���ޤ��4��R��\�Dp4On���F�7��l���暥ZWm��8����,��8�+SZF2��ô@�^3�� }#!�n�Xٱ�9Y/���=�`�(b0�w�L��2Q]���,{�߫z~�}�V�?�%�p�ᇈ��#�|���>�9�[�;+ի��G�f��OPڣ�n�KKE�F#��3#4=���h�feq>I$�"Wb�������뻱w}�2�%�J(
Z)(aO�k!��T�aY4��d�kCe�BXPP@����Z]�`�qz=�Jk��P;e�b[!�Xa`���z~��i�2�h�L��=I	���HR�p�\��������f`��~�/`lN�ٟ��������If�}� �%�
�Y�HL�K�~t95πa���C�U`隻矉餶���/��5�W�CЀ�Eh,�؇�wv�9��]u��s�zo�S�>��C1gĂX�=�	`�7�D�7c�������&�]v3���۩=!^&q�
�b�ls�����k�2��m�Mۅ�s!���|��Q��)�[��1J=A���o7�dZ�ޗ�VQ�I-3.�kT(7��(�=����|i���ff����Xk��5�E����ws�]^�--������Y-@���b<������5��c�y�澐���$|�#��4��W���;5��ԋ��l�����r�`�r�)TUM���ޜ��>QG�h<���%~3b/~$ۍ��e���\�[߁��v�"�
@fed�f��і������}�pc%֭k���k���>�=2D17q���fn<��pݰzu�tv�=�+Tꭨ�:u��{eѯ]ߘ��z~�oa�r��"����7�h�g�3���i��b/��ߪ{��YXlM�F<P���.��
��N�&`��KƕN�?7��
a��V���:��E�xA�Nf�w�<�-kA���m-(�Y���U�˾eb3���t>B��H��U���ϼ����qs�9}11%�2w�:JDD�1���}�b{�{㑗/��`{����}A;߹����S<�5����d(0�ݮȻͼY<���!��N= �M�5t\]��ŋ���~q}�L̅�{��w���ww}��#���kZѭy�q
�@��Cb8�5t��T��<ق�2e�Q'ۈ@�N��UL�%��V� k��3I���!�m��C��l�V`���˽�����qn(�<ت$��M��@�i��t���h�	i��S7�P>�+FVܹӛ���f��N���$���m�]�.���fÌHoB�myܶs�Nyv�������Z�M�]m����`�8��z�]-��[v�n)�9��v��uʞ�1l�����+5\:f�v�n�ڪ�YV�*�P   ���4�]7JlL[.�5hְH��K���۸��)V������﨨��+��u�*"�!� @�`�C����3(�$��j"���b��Z�fd��L�N?k�p�c�-�ƛp�Ç�0i�m���u�ҝ�Zpv���a��;v8!�p���v�n�P*TD���<������D$�k,��
��'��jE~��[81�����5r�D�ӓ6�W������1ج��L�2E��˕����k��t{�3hl����b�5��a��>�g�sV��KI)Ao&7�x+W�&k�D����Xkw��� j���E��3k6��6נe���蝖$R@R2��}����|F���}��[��Ƶ����������>���8O����������ȉH5�����(�^����p\�`e�����wj��al���xb%�E]W�]o�/訤�A�R<ܼZZGN���KK�a���H����ύ�f5i*�Ca.rj��N�9v�=L�QS聟LY��Onvnt$9<��1�h0��0��EJ����誓ݤ��w�����rfd�YN��ԑ���6��:-��x��:p��qW��4��Q����������.�h��5�w��q���g��+����;m8�ݾ�#]g�H��/�m����b�	o^��1C��l�}��F�6�px�����n�Yt�0"���v��b�U�w�|-~5� ք�?3���7L`��zx�ٛ�~ �mD�#������w1>��o��؜Qm�|daiOFq�ȃ��#�j@�z��{M.u�h\*�]L�ĳ����z�^ux�2+��n�Yl#>?	�/�!<F�� ��ޯܟ��H'J����@.kƺ�$�C�-9�����A�l�V	A�A��&�6l�g#m۔�
ENR��CssS����� }�7"W'=���z�E����k���g*��:�)��H�o9[u�V�k����������}uu��q����شh\8lغ�j~�.��p�-W|��\ؙ�B�_o��\6� `υ�p�Yk��H��ț�Ge���ե�� ���62�5�8�|8� J�{W�o�b}��$H�A���H�$K_�[Hӥ���d4熼�J=�[A���&Lȝ��ޢ�!k:oo��ؖ�����7=!z�R�n�W!��\��@?��C/����$������w$�DGw]ݽ��wbG�㻮������w q`�4��4�vo���*1�P(̑�cM���YC�VcA�M%���_=�?q�XF20�1ID��H�/��F�4���01֢��@��6!��$4 @�I�$a6�II���쇃�~��`�q��n�{w�20�ga�f�n�Q��{�I$t��u��N�x�$6�L�]6W�c}��4�ĩ����?�M�PO��}{8/��t��S�L�?���Uj����K��p]<�5�K���><���]�޻�3U�N��;��������vu6��.�����~T�����X��y��Q:R�a@�ZMھ�3�hJ���>{�F�L���Y��&���4�������;<�!�S���ê�'$�*�]����g6�����)7�z�uU�j��0���#�Bֵ���Ff&[������h//b�Q��}X%�鳤6ݪ��(ii#IO=�#���[N�3�om�t]o�mt��`f���m*����E��ٚ���$�c\��<����8D���2B#H�u8�p�s��ij#IìK_8�v�q�!oI�Aae
ZH��b���\z����WD6���h��Ye$($�G��>��v@�R��N$�>�o�>(H��=:f��϶��rJ#"3g������-�K�ì�#]���G���:\�c�������<��4���� �ș���!��.�O�33�lZ3���7���YX�p��z����TFl�pZ4���@�@�4��=π����0p��������!���@�~��+0�UU���շ<�D��MWC1d�S��2�viVUV��*p@���4�!�@�&,p�j�υ�8*c��U�5���M>�˭a��f:Dۇ>����%-��U+���t���T2Gs�Q�����Uh����NU��L����h��x�'��" c��{�C�����[Y�[M�-���!��`���8��B� t�ݢ@A%��<T2�q���:����~L�!��js�M��iM��8�x�C�Jϰ�~��2tUӈr8׫�i�m��X��Qu�~ 	!%�,*��,k�f�"��m�vm��ρ�!(���1Tv;ih����4@�|=>"~t	/krd��uLn�
V~���j���:��S9�Y��[�/�t�vDii���!#H�e��F4dqDk��$�`��qϐ�l7�����i���+�C<��?'~t�����~;�\"#����.���t��y�kZ֯�%�(R@#E%��&�6�� ��Mi�xH))�˼U�K�P$���yV�n�D�%v!'0;IS	�`J�'�K�I��Sإ�NPba�oǝQ�W�ȶ7�h�2[$"iв$"	�֪�������l��C�}T3�Y��*nYz��79u���a��0�Ρg�5�)��E=מ������Oi��&���Ȥ���ڟn��9�,�C�;ևh��jE�:��z�,S� �CW<$���BZZ�5R汁��<(��W4>ɹ������i
YZS%UT +��!�t�.�a�6��Ɲ��6�
�͹`��u(Ik*r�\��� �,K�Z�fg)��A�Kx��r�����a�f��h��!J��o=�3�^�%Իmx��vN7�i�"2&��.�j08U��m��D|ֈXnl����7�@��p,�.��l����b�/1f�6-�N��`;h�m<��"����E�OA3b��ضq!U�rpAE�$S���� �F4�7,m*ݴ�~5�#[�~�B��ax��O^}#�f��^W�8O��l4�g*�������џC�^�<ظS�����3�q�z�^������,nr^�qJ��^Qt��>�jf� �Zل���\1���|:S�<�a_}~����f��ޔK���7�u�rb�v�r�v�l�KY�h^��r.��x����^��8��A"�xD6�<r^͖���/�lи/�9�\O�ho>��Mm�2
i�}$��K�;U���޼��Z�Ȇ"�ǫ`��~ce��)�q8=O#Q������9ƶ(p^�%���K�����Qm"M���nN��b�n[���ϧ�N�� �݃�oVCv�vٴ�Um]K�NW^<}���o��.��nÕ��l �s�>�b�YQGZ�cy�ؽK���y�oد�K�h���њ3f��}7=%��2J�(�4�f��|��DK�|�as��>���*<���H�c>�0�`���D�<�LP�
#9�\2�����{kpv��-}I����	��`��/{�vrP@���kDNj����v[�x<K���b�����y8N���"W�sb�-=��l�8���qE,�JH3ar4�����<B-b }qg��!�����=9�9ڋ�g��y��ۆ��2��K����Ym��e	�9D ˧�pMi���U\�p���-��r$�EwTH��n0��V���W���\}U����1=5�&��7f�ts�k[c�+s��n2�Z��j����u<�`�i�l���~_��E��qa���r(�s%������
-D{����E�#�sH���׆C=��v�DV��GH��篧L[,�^	{~a~n�@In"L��ȇ��ţ��2�̨��p��yAp�yLT�u�o��%�H��6�4�%�獕��QZȺv���Վ�r����!jw~��D<wt����wu.w��ww{���4
b3�F�<6ى���:%���PY-`0`�T�(pn��¢`0���,�	FxgO��_�	�����%�1���B��֌>�Xa�����	jO�����貿Z��Ǭ�#�:۶d�Z)l�ZuÙ"�_�-Da�(�f!P�a�\3G�뺧'ʜ��v=xZ�_��k��t����|Qf����Ga <E-FΒ@<�K_?ɀ}�j �v���q���sָ��^��N���s��ot�\�}��:����ĩ���ۙ�0S���O\�m��=n��u�C1#�izB#�L�ߵ���I��m������P� �=N;�����4�#]r�l-�T��;��ࡳ�p"?@�Ᾰs3�������]���X���PI�נ��{(>(0")��Z1�~�g�zk�fC��/�n.�im���y���5Ǯ�)g���U�BJ<��T�w^q�\�.�O�x֖��G��G�� ����h-յ�,0�[�_8�%�q�:\Y���~�J���Ʃ-ߧ[��~��0�́E��-ݸ$ax�����GHc�w���5z�=���>5�Q�qq�}~�EM2�%�Zִ,[|"�	-Ñ�0�[KIg�C#������H��E��2��\�-�sK����縱~1#���,J���V�U%I	8[v�����Ó�V��S\-l��-�Lړ����v�eOP:�Amc����B�LX,�B���&�8]�Ex�c���9��~�ʴ_'�,�+�̹x5*wj�o�����0o�.y����罪���_f������Oy��D�!��Z(�g�d�︟7�b�3�	�~n 5�a̶_�Q율BŘ��9D�Z���+�.rޮ��=���k7�gSu1����R �"pN�O�q��*�#��;f�Ϋ��R����fp����7Y��h���g��;���K�������o���;��뺻���j$'HI
�e\h�dL�6.2�HB�T�/sQօ�`�	� m��3�u�Mq�II1X�׈ŵq ��8�9��!�SD��tk�y1��&��!� �D�O��?T���Cn)&�!��+�w=<y��/�sw�}w���^s���8r�%���2��<��-oV����6�́D�a 8��x��J�6s�%��&�|��R�-s��D<j�Z�E�;j�`�B�\q� �m���kJϬ@�w�;s�U*�J:��
�Uev@�����F&..�*�,m@)A��q3U�h�L���cP����@2&ԝ �R;*���m�ؼ��/O��9N�P�'jL�uT�9LN�Б܅٤.�����76M��9h���7Uu���	K��x7��9J� GAE{��w޿|���O��A��{~��}��Ϭ��-��;^j��Хă���Ǣ������s7��eຸ�����Uu|C2���/%��^$<�!ej5�֡gd��h�˿�_O`���*y�s~���z��j�K�*Z�<�g����TI(���w�
"����~�yެ{yvG̘��my��+�󇹒cx:!I	F��UQ�#��?57�����B���~Ղ��>u��N���	�#Q�_Vh�T�&d-���	wRs��rh��c*�J�{UXN=�"����0����c~��y�ēNځ��3��*U� 	��K�N�����jX�$��V�D({�v����Y� ������7Woު8n#�P���>ִ��w���:�E
6"����ַ��}.:�k�5=_��<��9�����ϼ��~�$��2�hX*
��y�#U�M�ٰ� ��#n�>$.|ٝ�[K\�m%�s���>�� *&Z8C�G��>���)8�Qۃ��/v��VG�޵ӓ6W�3�Gćh/ �:��/흞_f����x��L���m�����9=j�k�K�i�$�1;iW���;�>��S|$��M����_Ug�u��>�|���Pb��hʊԫ8��W[_3��z���m�o,NP�k�
T��=���s�7��m����K�b%�'8��0z��iY����w~�r\�������s�wG]���t�Y� ���t�@�S� �`����"�!bJ��E�:"��9(���T/�Mъ�M�3h8�0}�I�U���H�7A�u��Z @�hW(���GO���s�[`z�Ôp����^��W^�m�\�;���ڥ��B:�NQ�S�8�'߾s�x���jK�'"�d�<���غ�ƾc�l$R�	��}�#��o�h0x�)��C.��xa�5Q��}|F	����^/���1+Z�	@w�f��wV�Wc����e,�D������åH�w=t~ĳ7��3�}<�~R�Ԥ�n��~������v�"��1'�adL�鎃��kZ���e�-)d�)d��S;���w�����a���1��}��[]S�([ۊ���##߼3ӮN�,+tɑo�z,S��
w��"�3㻾�g6���󿵣����'Å�*v��Ȫ،���Y�}U����ufM,��|ش����ֻ9��Q�βXW(X�N.g�ýc՞y��3<w��,���q��.Ƴ������=S�y��Z�̣�e�ez���䍎ۗm�q�6ֶ����u�n�*�eˠA+�}螒�b��8F*�VR�a�a�>��5E
tc��RǠr��Z���۝ 8t�IS9�s������?[|蟑o�W��y�MUO��f���%��^����5*c��|��+ػ��)���Q�W�H3� ����B?	۹�d�����\S�w�b$��S1��{��9��J;�t\z����֑˪����L��"���<��N�3sy�=��;,p J�7lм�ȅޙ�Ǿ���.C�ot<�E���}���?��7�DWmTJ"���UϿ��O�y�%7��?���s*�J�jR�eXR�J ���CrR��9��#�U�L%rU!@� U���" �d�D��&EbEhE(�`A)�ih@bBA��cd��ʴS@�� ���@S@!M!P	@��+���ݩ"
��@iF���Za P�-��fFX)�{Z$*�d���IC��1�y�T�SJ U !E%f&��*J��APAUQ��DIp�r���f%�M-+�\�4p֑���(J��C@���˟���h�4�'�  S�E)9�m���?��Ϳ!�z�� ���SP�y��PGH���#&�LUN?���[�>?4m��#�T����'��u���y?��Ѐ�=zQ�֨#��E����u�O��������<�@}a�F�7��������w�'��~R(��Gg"�x'�X�b��R�a��o�P_�wf'�|w8���~�QK^���f��GA�ۺ8�*�s�{�8]�mI��.l
`��
,$��D�IQ%3�A1(Ԕ�PI$̰C,S@�C1,L�RHP@�� ��
�A1� `�`� e�DdB�*��!���R�J 
(
)
@�i
B��Rd�@b#N8�-@���	BQ-PAM0K"�HT��� Ҁ�@P̑,DTP��R�!JSII)R�\s	�*f��*��
D��@X����!��I����I �&*" � �DO)���(%
�XD���V������q��s��� ��UX��hP�w��=�Y�9ޣ֤s��Jq9���O���������G��*(Ft�{C���^�E�N�Ƀ��>w���������w�{|��.����DP7t��M'pg���
?.���9�ܾ<ϫq��EP:zAE����jG}��`,(���?�aٔ�?�_hAP�8�U����~xP��P8���?�TP��檢(���4��n�����mO��(��0������������s������{_�s�t��*�9��o��:�}�'�����6Q�!�@�|Ԣ(a�
��n_�j~�/gO��=GH������6FPw�$ƧW�=Is���s��+�����:Q_���s&I��A��u�z:y��R{�#�E0��1��7�7���������4z�]��@�T?���
({�'����k��ۄi;���v��H��d����H�
G��