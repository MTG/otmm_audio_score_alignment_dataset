BZh91AY&SYR�����_�px����������ay�     =�@Bl� ��Q � 4��@��֠)BIBB�

HD �����@�@U@H! $H(  �   �*�@	@( ���� ( � $��� )G �   A��� �4
 P ך)�������c��`� �E���Ž�  /��9=�� �&��j�� mB�&�J��L�:��j�K �LM)T�ЕYj�4�W�   ;� @   ��L����W|O'y��ye��;J�ru+��}�o��..�6���Ի\Υw Εgj�9i| &���s:�  �{j��asi嫞ܪrj���P}��b�[mɯ����K������ ��     �`�>�b�Ϸ>�{��y}��{�@�>�m\��U���O+��ޚ� 
v�K�{ۥ�� C���p���z�_x �w�j���Mqu*ϷJ�<�����A���g�T��_W��˔�� �@ P  
� �` �u�m�V���|�\ڗ���w� w�Vm�Ӗ���w-��u]�� i��Ks�;��&�Ƈux���f���� �ޕ,���W�������y�ֽͧ� {ʥ�T�f�k�nWz�/J� =��PR�  P�Q�����\��+�Om\Y{��3T����w��r}�NYs��-K�qe/p �w��s=��]^  �͞���Ou�p :d�e9湴��x��� O=R���KϷ>l�ݶ���붼             "~�SyJT� 0�  a#$�*�     �B)��T�� � 4�2`��R�mI��     0��!�)J��40##@���
B�F���6)��<���C&MF���?������S�u����ﾮ���{��@_CW�� *�@ES�� *��U�%�(�*��yV"�*���J�u  *����~mT�� ���E?� *)� O� ��� ?�
�iO�"!�"�}*��� }*/��J
}(���Ҩ��"?H*� �ЪB��
*}*��'�
'ҀH*}	���(ȏ҂� 	�B#�"�(�@��ҪJ�}
H�} }	��@� �~����C�P�S��MH}#��BJ��)@�B�@�҇�@�>���@�S��>�>��T�D��C�rS�a}�O`Oe�_�>����O�C�>��~�O��ПBНK��J�(}#��C���S���F�$NB��JP>��O�~��@�B�'p� })�=�rS�_�O�O�>�>�>��<��~�5��H�n_�O���@�P>�;�>��O�~�>�>�~��D�C���O�G�2G�E���O�>�>�~��W�������E��>�� �_��~����ҟJ�
}+���(}!I�	��҇Ї���� �}?KA�#��B}+��"J� d!� y�?Hj�A��_��#��?B}}*H��
{ {'������/Џ��	���H�K��J��ҁ�}!���_��}"} <��O�N���S�G�_$U��Q�`T�P>�>�A�UN��Yο,���k~V���9g;��E���}�����wݟFH����d@E�q��d#B
�A�B��%��		D�ڥl�tJ0#v�F�6��dR�j��v��`���`�����r�?B2�~�9���j���&�%	��5	P0�G�Д%,��p�&њ�d82j$�s,�24C������3!5A�_w���Ì`j"�>ǿO2�"�1�NC��8�58�&5��̳��q�vh!�P�غ!t%��hR(�뵕���wA�r<�'��P�&�;�N�C!��â�Rvj�< �1q��9��;5��k��'Rm5.�؍Z�h������cG0:]�@d��pǇ���[�f(�l۳9ѣ"MNw:09�4�9��I�PƊ����JP���p!�,-�m�_�`N�(��ز#&A¥�ePf���Wnc� $���x6K���P<�\��5vM��}�:#B$*p*l��jяF����,� �8d۱�����Fd�5�<٦/���w�{����y�e˂*�l�<��s��;=��(( �2Pb:\�\�r�89B��"L��Y����2qrL ��.���w��1�d�r�����9xp�T@�ʘI�<��:Q�U��m�v�		Ó0��p�Q)2Ji�����:ѹ5��8�!�ݎ�Tu�ܚ�d�Ǣub�FZ������F�4����c�8M9BTF��Mo0� ԝ����X��xw����Pd�Fh{�\��X��-�6]���7��Rq���q�����a��y��YJC���}�T�TXK�ξ����[:���BX4O��HV���s�����'���d^�����5y�y��M�DI�۾Z���z����\�*��'P�'3�(�a��=�W �gA���|�&G�ՄIޱ6�tv���y�4o	�Ύ���8�|-F�s��6C��:'�7��K�Bl(܇:�h'^o��~�j�Cp���\����0�xC@$@@Ff!��׻�ԋ,��������¥�ܴމ���X�GC�q����L����� 8d�΍�sd�oZM�Ȝ��$5���������� ��t�	C�����J��(Nf�%�f�#�ޠ������w�_9ڴe_H#SZb3XA�1v�8!�&&I�30uιLY'�V�3̃��|�ᑇ7	F59&�'p�Bu"d'y��I��R�.� @V*@�F2���΋��{��d�$��\�;�)�� �C��MBP�	BR�y��u�4��bB+�q:5m<ޱN.�ٰ�Y�xƭ$h�Dy�n,�]����D��z�I�d%�,C0w�X'!2\ya���8vo0 p��J�hY���u�{�"�T6�c���t<(]tX��X�� �!p4�LL�H���f���2Xv�qy�rd%'d�A�^`kw}����0�u.9	Ho �4owy]�7�Y���4�	A��3ս=��'Qo\���C�Q�v����Y���Rx�Z�u�CYc���C[h���o�F�79���J�$�Z4��'��E������|�z+�3��0լ=�")�a�p�8�Bu	�H��sXﳮ�$rx6��'ޣ%�Li�j"4j�D���~w흇Mk è{��4��xɒ㑎�[\r4�<�Zz1��#As.㸏q�����7f�x��)ڣ@�.T�$]��� 64�	hFf,�yd2��X��s��"�@S�`��i%ˁfA
ch�#��ݎw��v�x%��*�%5b��B�e SX-� �$ �;��`Έ��ͻ5����ɓν�ç���j�PwHy�17	��NBK���,/(��8k\��0�3��#F��:�2���ȥ��V����f��@�FW(������t� �4 �P̃��	I��Ձ�Jj,�W\׽uz�ےq2\r4{�p̓,4j�o@aIul�'^c��v^F�9x:�z:����gswu�In�a�5�A�]��;�uB[8k�Gq�I��,�ש�N�.�������N��Q��'Y�x��l��\̺��Vt�yk�P�X�'�2P�m���J�J��J����B���j�љ��ѹ�q#''=��>���7'Sdɐj�����a�N�::�g3o.ġ)%�m.Pbi6d%6��'���;��q����9�;BE	@K��$P��P���LYrBP��Q��d%P`PQ9��k���hᢽmh0sI�=2p�"BJd^�`��#C���n	A�r��4�M���N#0J��A��u
E,��H��*��X9|
��tN��%	By�%'!)�� �0��BQ-I���(v	X:u�k!:�� �B$ A$��R:3�9��@D���d�2��͘C�Y���	����jѠ�t��n��k� �1�����T�a���Y>�~�����)>2�Y��ܔ�ˇ@)��BG��i�g��֧Np��b㐔�=��!EAn��.h#Bk+�����]tvBV�I����aa��u���>c5��Iy�����5��2#'(x�6ƫ^���E84C�/��v{�Fkz��wk�:���]�P;5�C Ɍ�i�㖍zX�ѫo.=K�}Bk3Hy�g���K�j�g�X)��c�]��4��u D6ڵi�G��<3�N[39��:�N:�Fyd�}G7�����]�An��@���Th��
m��=�;�>���F��-;c5�	{|9�m�F�	�&��Ǐn�����-a���{5!�vÖ!�d'��	(��I;rq�# F�V�-e郱�� ڸh]E��r��@T�;��S����L_Xo:üL�&���&�(�L
t�5.9i5�P�3oGOf��[�C��r �!B ��M�V��]�H5KB��h�Hu P$�
�V [3Y�q��Q��Q��.98栠H�M1Q�:1>GwAAk*(� �P=���,�4z
��}�}�0�N���%�P
� �!�Ue,>6,�e�Q�Ns��,�!�蔹�kf8A�Y�]kF0��4f�V�j�P!4F�#E`��E�*$4j�eԐH;�� �$c��ػ����nZ�X!ՠ�T=�R�5 ���"�1��C+ �	.������h۬4�nu����`h�%b��.Q	�(@N��(Z��n͎z^ƶɀ�O!(�2�t��)�&A�u�	Z�^�34`����x=�ZߕɞN>�7ۚ6�i��9�@rG�y	C���d	I�f	�`�<8k���u���L�$�6�`dǒeo��1�x���v�FQ�Ѷ3��Ǝ��20��{�G��zu&&@a�q�=� 6f�� �Dr���NyzK�-��p��S���p�q�N���p����$�.����'i݈d�}�W#��Rm��Í�ָ>�Co��o������2�6q9�k15By�t�	BR�bd%	K�$337�!�:���˕݋�V��u
�E"�9xX.`Π:��,w��3���9�Ph5	BVT>K�'0����鞢������7yh$�1���:��vq|�5����,�:8�����q�=I�#�d�b4�8���!f�<�ep!0v��Z�.Y�5	�GL�I��>k4�pLД�E��#FdDUJ�`�ͦ,�[0�F���v���f���	�M�Up���vm�a���#W�1�7p�l��z�:�nb�:����sIe�'z��p�.���w`a�r�����w�Y��.y��O�^c�j(oc �p�,�0�j����x��!9�&��d�:u9�I�W4BT
"D!0̃�m��l q�V�ɗҸD0s����E!�I��rsC�O�(z��49	BX%	N�r��7�K�T��f�R4�06hh�d;K/��+"����@݃� ���p��J���BY�A��j��a�ヴ�X��C��7���uAdƺޝ�̹�=�eZt٘fLZ�4h9�К���R㐚��P���z���:�$3�Oa(Ou�r��lC�D�F�2tY`A���`����dh�W��F�4;���=��`�3���w	A�*��8NBP�'Y�Z6��ݺ���`�u:��%	hƨᘲ�p�0�:�޷�䙉�j�BS�L��;���ѻ���]y��QR`PT�I��@f!�	�`k<��Zeq7fQ
Ca��z8@d��$E(���4oM�$=�.�2هF�#F�ՀY�5�{�5�n�4Yw�FC�C"�h0�HuFN�!(�ka�#'k�p2�z�{k���Y���kSI#>f!$�&��#2r�"d���N��23�3;�N:��o�IOA�V$����Ƨ!1&	V4���/#jLNd��&���}w�ɲ�� [��!0��58�ݙ$r;F;m��f�s��������K��)6!$B؎�FX`�M��f0с=r�q��ת��˷���܉m���X�:�����c�Xg�I$�I$�t8    � ��   Ή -��8)@A�m�   H�   mK@  4W[@     H ���  ��	 p6� p9�"�G�  
P;e7i��mmö,�gnP.��xB1�v���TC�2�+I��H� ���F@
Y<[RY底j�tN�s��s�mm[$ lݶ׬u���.��T�+h�S6A0�m) 5W[m:%Z�uN����"c�!i���y��>8-A�dn�L�֝0�q���ԝ�FM��n��SlJF��:ٶ[u�ǉ$�J�0��7\5-�+s�j9XhD*�^�M��;fphmE����VWj���{p�T���j��jPp:C���U��$Od7`n���&�� �]*��:7 l���nh�U`�qǍ��ꔲ;^Kj�Uͪ�-Ө�')���&Wr�t��&���E7Zx9�rg!S]���T�c��W�U�rm%�����-�� NY�;\��tAv�u�[ql� q�]$[� UUT��һ/�"OcX�i�v���K��p�I'94�  ����� �5�6�	�ĝtZ[$�   M׵�mu���ڬ���Cm��͝�Y��   	�� ��He����(-��X*l�@�!PU��ZA��e�j����.��v�G�O�/�/��h�B�G��⚶@  -��]$�ێ$}3��ݗ��� �`� �kkFݴ��#��#�]�ئ�ٺ��۰�U��P��E���λa1���|��Ij���Ӛ6�:�6涐���*���1�� 8 �! h�t�.��-�H$sm��@,0�d������uk�A�5��wm�m �����c�A�6ذ�nR�7m��  [�涀	   Xbmqm�� �C��j�ݶ햂�Hݺm'MM l���+P�C%���b�6� ��1�g6HF���%Z����l � �v�I��m�I�  �xm6`�[���*ݷf�Ve9�D�ru��t�H<a��5�tc��O%��6�ճm���:9%�� �[n-6 �"�-��� �m�t�p��M����h K�cm��m'l  ��7���|R@mR��[U/kɤ�H�L` m����D3F�n�0H[D�"BI	$ ��Ŵj�$�$�-�p��8� ��m   �  k��m � Hf��Y�l [[li1m�� �[Ku��ڶ�-�   Ͷ �ۯ\��  �� l� ��6�m�  ᢭��kk�$ �h�m�u����=�w�m�i ĝ��	 �� j�  �I6[@8�m�d�t�zg�]o�w�;��|^�=Kv��^Z�W5��ij���[*UUU@O/����(l�iC�M����H[zpĀY�eV���AR�<Um=Tͱ����/+��6��K4�E���	�sj����i�k#U润iC�i�i�kd��$h�� ��e�R���ٳ�n�6� �l��,��A$ ����8[A���` Im�6��6���UA�mR;nUkj��dT��kj�j��U
��A ����8����ɐ[Am'5�l�&�l���    9%�ֱmI"CE�m� �2�Dz�p q����� �`� 7m���[m�m�-��� p  7m���   �z��4�v�p i�V��m� [m�ZŴ�6��m��^��m�    �m���v�H[C��` �im6�N��.6� o���mr:�ۤ���l�E��}I�ހ  m�m�Mm��0ӥk4��H[L��5U�J�F���'K�l�ԙ�l  �����$yl�d�b@H�b�6݀3��M�v��L� �M�������z�J����zu(6�m���a��[���6ٵ��H^PZ��2.Ҳ���n��(� �m��s$��՛cd���ݜpm�mt5P� �`��:`:���$����s���@Νa�����m-���h[v UUC�`��h�FDE�m:˽�������l^��l�M�mm�-�p �Im�k@#��%�[M��[dh윸Cm���B�j��0l�*ԯ-Un���-qT��,���\g2�ꪭSPN�8�i%꧞\Q�$Ud���'(�����UPq�U,
� $9�� 7l�2k�T�a:%.m"3�m6b۷f�m�kt�8	%���kh����m[dlYز�o4��.���E�P ��Sh�a	]� �gͩ t�6맙^���T�(�CF66̴m���Ucl��,��bYd8)�ź���   ,�ە��j�:��c���o���Oa����2I�ڭ�mv¶ t�m��$j��.�E�UZ����cqUy�U�i9xH-9hj�7
�RE2�T�q1�{ln�6�*J-��`�e]mJ�V��T�`	V��
�n׍U �@W=IJ���e�ķ6�a��������pY�7C�P�ڪ�W��%�k�\@V��    �i��m�(h6����UJ�J�pWl��UÒ ��n-��	8�i�>���u�� � l���8Zl4P  $l ���tE� �M��ݶ'I��`6�d�m ��[pև\.��f�ֆ۳m�89m *��i�WR����m�%���]ml��s�	�&F5�  [E���   6�@m��lӒ$Ӏ���h�)��m�m���� m��a�@� ,6Z������̮l�Nm�l$�mv� m�   l�h �8 N��i�f� 8 �u�H H�#m�m�l6�E� �kn@n� H����Un�k���[@,H��   �M�lp���UUJ����������� 5�m p6�J���.ԪpPR�(6�Au�,S��WD��$�vE�6� H�l �����l��@T��s[��v�Y�[���{Kn���yXr@��l� ,k$��v� �2�	 ];b�X��]eɵ�s���l8j@[m����N��X�KCne�Fɰ�b�vXyڥn�wm�UZ�V>>w�Ӕ�2BWs���ٶ-���m�A��׍�
e�V���]���^,��E͗M���J��Z��\Ua�Rgv�ŝ��Tz���,Mc�$�n6��<�·W\�U��p@5u�:w=*�A��ڍ:��d�`�Ͷ,kiE�� �v�!����[@8a��$sm� 	��� ���\e�/C� �l����\pm[`�I3��  m�  m&�m�*����F��6}�rcM�bI�O#08m���I=-�h4������ �mI׭H   �Ŵ ���p� 7m�p m&��� $     ��k��Xm� �I}�۶ؐ��6�������m��:�        �[Vһ+����"V���Z� -�e�%�WM��� �\�` � �m�o}���$ m��l - @��A�  שn�݋o-�� 8jZ	mm�$l   6�hx�I � m�� - m� j�`  �� -�z�  ;Z�m�� ۭ`$�l  ��h �u- ���[[v@�W�]�Q�UUU@[WB�T^��6BWb�6�Hֵ� ��e�%�  �m%���D�KU*�UUJ�դ͵��Ľ)!� @�J���葃m�h�  �,"�f`X���"��KM� -�k6�	�"YBڬsU�Kh��hmT�J��J���7j6��     XI��p	m�����& �I�m�e���m!M�0�8 u5�Cj�δm�m�\���%X��V��
�Te�^eM���mUV��M\l�khؗ���.�H�fU�#M��;/W+c�uj��S��f͛)h����X-�м���k�&
�xi�$,�`[Z��$�H�` 6�[u�n7m��6�u�� �`@ H     �$�o@h�ɶ��=�V�(�k�,3m��N�6ذ��m�-��    Hm�  ,e��t��\����I����       ݖ� ���v������ks  $  ��6�H ۰ 6�"�A��Z��*�P @�u��kh  �  lR�^vBz�ge��U�8i6�L���`�&�L !m[R ���=\ڕv��R���ˋ�l�������  6�[@86�   � K8�D�O���*�����x�(��y��D����Q�	E4TAIMa�TSUAC�A��fUCd�F�0��ʀ�#�' �*�N�FDaa�@၃���)(�����������������������������            
��@�D���(�O���,�2�B��02� ��
v��h��M���@t� t�H�P�G�C��&�<a��� �� `�@��JH=����%SH <Q�T�^����4��������cg���P:C��G�ETgC�� �"'c�L����Ǳ��D�8��	�
q�y��:!�D��� ��P�Ā]{���}�_0� �d&�)H�Q��h`�it.��G���)�"�⁈���	���2&�0#�`�'���U�@�H���*� ��|N�8�qô�⨧@�E Ëצ
��ga :{%Q��t�A���DBM�/~�0���; =C� y�M/[�= �`�������!�=!� N�YM�plHX@�	��$�)�J'��+����<OA|
@�����\{�У�E�<�T�A ���s�QUUUEDUUUUTEUUUTUUUUT                        UUU_���1W�����G����G���/���_��_��u��7�������?����J�-Q0u
�+@�R"H����J$4�+BH���w��~Z�ky��9�����c��i���ȧ2>Y�6�+�̅�%�6_wn���A:����Ig[�n��Ӵ+H	�{RuYW[.�l��^�3��ų2m8[F�H!\l٫G-�ijR��Q۝m���tlE$��]TK�s]"v�冎�ܗ08+l�;
�nm ��\G�;������`.�[�<��;mdq��g�pv������ͳҹ�G�;m�}�ҤH���u(�	�b��fL�Z���:�mU��)����A�=�vkJ���Z�vn��u�;3���"ѝ��Mc�Tm�3�mַ�t,N�֤��VI]�zs������)҇���΄��+���g���px�����_?g9���+����s��r��W�`��q��0"�9H�X�����l�4�R�<�U�UiFbZ�c]3�8��ʽj�.Q&�*cZ�mhA�,������ �s.�ǜ����i�H��(�E�V���� y�ZB5M�6Q6���W��:�I�Jn9���O[/򒀡��[[����ʵe'�0X�pif`�e[�:Xd�y5WU͜[t�ݍXh�Ή
��8�>_bH�\`+'s���ckv�Ӟ-6P�"`�f�<�ѲcQ�������`x)U��۬�5�먖��(,n��:Y��^Ҷky�k�����C6p�+h8R�ykju
�"Z#M-դ�Ԓ�ŧ@� �j�NѰ�e{?�_۷]�K	���s�3�8�K�8�4��8��zy���J�.����=�#�\^^���9'����l�k�ӡ�m���Z�
��������O���1=2�c;`T� $.�b��I-`�>�q���Hm=+-,�f�P]�Kq�岱�V��:�U�EU!5�eT&U[xޕ�� h*�����S�J�M���W��;Z�o6^������ u��n�w	�mT<m�^�:�.`.	W`t={lR�WS��{t�$ݯ6$8�o$kv���
���4����Ej�N�GvM�`�5���ڥP* 
��?7w{����	�p�,�D(� ,�'���lL�zA�P_��<D�z#�5��gg[w螕Ý�2��Sbά����[c[����+��s�5�Qͳ�Z[h��۶�����-��3�6d-�k��[��ku�Q��{95YYE�cU���fA2㡛n�2��Û&ɴ&�#{un7$vűNۓWZ��8m��zuby�;s��l���B��m�'�r��j���9�9�	�;��Wo8�!ݒ=�FV[�� ��i�&; U E
�98�E��a1s�wn�s�r�{�۶�ɱ�$��'L$ (n�P�Os�w3�VW���O}酁�ՏbA��Ȥ�,�����*�Tw7n�nM,��u`�����6��8�{2���za`w�˫˹���P�d)EI%$��酄�3lY���hQ�nزN�"kP�n%$n+��]X���`sٗVq��~�g�J�i��8�B��	��������w*����ue���\�)خwF
�*r9����`sٗVq����I<�Z��I�P�{�O^�Ñ�}B$%�	-����7yb�=�eՁ���`�Ecx��T�D�Vq�+��]X^�v32���HT�(�P�*qYԼ��V�s��̺�;X�����Ǒ*t������~�`JU�̕�;ט�'36Œpfhj���DюFYG��g��cm��kt'm"۱�W������aq���qԡ6�R+��u`s�1X����X��FB�QԒRNJ�9�Jp��# ���8��0�đp�2�8(F�=�eՁ��L,���fq��#�ؒ��
bP̨@C"��#�T��yb�9�4�$�t"�hj)!�G*��}0�9��V;酁��WV�_cb�D�:����,feՁ���f��ͱd���7� A�)�6���qx�6r�gl���#�Ս��uwO��D�٪ Cn2�(7
D6��'�������7��0��F�S2L���	 )��]X�=�]Y �,i��bA�$QȜ%�;��9���n��͐��N���0ڑ�%��v}�����*��@RA�0��
'��u�~��e^h��Q�$	9 ����n�s��c�� �UUP;��^	�A��`�\�lս��Ÿ�hw �.<����/>�NǓ�n^7==;�`�.�n�N����Y��q��ަ���"���$���m�n����33ea�uTe�5
4�R]sw`�ͱ�� ��m��N����j"Bn}�����3ls7`��(,!d���,w3`���g���ͱ�h��%%\�P5$#��^i �9`��.�J3��Xa{s���Mdj.4��n�Bŗ��h7;&ֱ:�=k�МY
ڽ�* Ҳz�h�8<��x�퍒vy��U�7/���kd�WX]C��w0W�i�}����ܺ�^N�S�]��n��v�n���;��}j��C��`�����<:P���=���K�p��N��Va6����F^�:^z�-�a����]�g�&�85�竐.��pA;�Z�i���r����볦��̮��ٌj7��k��A(�iM�-�~��E�Y-r$RE��\�fn��3v}����3�OH�mHܒ�3v����X��@/��c�	8��1$�7 �ͱ�͔/��c��Mw:ւf�',z� � �L��@�nz�3^���m�����JBS�G ����צ��ͱ�̀z�7W�����d�]7oǮ�Źۜ��6_)�g�Ð�2x���{'�]uB�.8���������s��f�/��u���oDm�Q�����z�
��A�@rE}Bk� �7v�3^��đH���)8D�9c��#����zk���tkؐaIn'	�W�;�z�w�ƻ�Ͱ����Ob
LiI#r��k�^������]i���lf���`���Jn�̊�n��ل�m��흺����ո�Zz�l	1��(Ċ@\p�{�6��l����uV��=h �Q"r���B���7)�5|udt�"k�@�����'���=�b���Ckj�EP��1����l�p��d*2��$��3]s{�c{�!��wli�S)�4�DK��\������3li�k�pnjx�[�Ї�u��>�5��v�8a��GG3�n_��v�N�`��[	lW���l9��{����z5�I����$݅��w~K#���:�ϩ�%�p�|�e	��D F��'.���H�罗Y���wls';qF$��C����X��҆s���� 0��n*�t"0-����Dd��������Y���ͱ��lpB�dDTrQ"�e]��� �x��y`�������\��^wF1�NG�7Vj�gsln��9ähoQ�(�J"����^5@
5DP�@���_���;�6�q��4�@�q�\���n��/;�cuf��Ē8��aM���,ws`�ݱ��Us;��t7� �8�md�H�wlf,�!�w4gf���D
 �	C�]їa�ʁJ���QD$Qq�mG1��F=ݩ孳���q��b�7��yѨ�d�c�q��(9�����f�k��l)D�`���#��6�m�+s�9�N�+���yvB��Ë��c�#�n����9�n���=7�-˛\�q�q�.�n��x��< �m��y�WW/@�`��fL�ܕ�G����:+v��v�e�^-�5Y5�E����7>�o�g�c�v��Q��d��&�f�6��.5Q�'������X�ki
e�=���J�w6�7vy���$�'a(�2J1�\������9�ݺ�͕��D`/da�
���9��gwo�Dn�w}���4=A��0��N93��\��\�ͱ�̀_N���mF�h5FIu�͜#¨�o�;��gwlv�A4@oLO:��cq[u� `R�-͵�Hd���t��Mo&�H�!m��p�W77ls3`��^���*��I��!1	NY�]�����
6��^��8y�5���c{�����H�n����\�ͱ�̀wE= �	�)nX���\�ݱ�̀�=Y�c��h���@Jq�37lz��}`no�cs]z���;���		��#�$޷��ۏ���vn��#�vtv�]N7����s��fH����a��{�뛛�:sCH5j4��3��~�G������j��{%m�i����E%�&B:�sWR���"~]5�U���Vfe6�w����%����;B����Å�׆���ڡ�$�����ޞ���"���@��b!��&�8Gq�L�1f�'��v4Ҥ&p<8�T5qW|-`��t�%$�:0�f�nZٓM��-I�7l*@��0ʈP4/x�0OjL"�]�:�1���S0::5�euqZ�,� ����@0����sQ�� ���� EG��P��p��(����J��A��� i.��J �0����gN�O�?{�����%)>���pz�iK߰����&�A�qH�U�"�Y�}������~p�4�'~����(??����Ͽ7u@��H���I��#�N���R���~��)JN���=JR����)@����pz��?  >�]����$2Z��޳Ւ���7h۶�us�')�r��֎6�h.��+��AFe���JR��~����Hd�����({=��=JR����8�)I秞�a~ �	�)nX��MP�3|�� 3��>|}���������R��wwޱ\ Q5C�	>z�I %8��)C߾���JS��~8qJR��}��R����k�R���ᗥ���֣y�[�9�s�ԥ���ÊR�����pz��=�=�\R������R$H)�X"`bP�<��H��<��pz��>�?Y?0aB�R9u@�(����WP$B}�߶߾��ԁ���G��d�r��~�B�q�t�q[�k�Ϸ�a��e��G��p�J^��nW�6�`;On*�����=�=�\R����O���)Jw��s�R��w�o�ԥ){�֍}�5���l�[��\R����~�|�)N���qJR�Ͼ��R���h��⟦c@�]��$~_"SBB$bXI�خ�J�����)JRw�}��Cްԧ��@�(�Y���WP&�j�����[��V�[┥'~����)O�׿g�){�߾��)A��/�}���)7�|�6��q�����ǾV�)C��}��JS�=��R����~��ԥ)��)�O���5�Z5�f�b͚�b��]���QCm�\�qZtۦ�{t�͛3r�.�m���p�݁\�l��m�����8���\�)3�N���u���[v;��	�[�ܜ/=p�k�.�T2o]�f�����P9�u;�V�����X0G����f������Un�Q;�M�ɥ�r��MR�ɑ]�E�ܻ.F�q��gei�O5�iq,��ݔq�ݷ~}���m3��o9�v�۞ѺQMyք�x5����|'&�\v��w�BBQ�$'�j����߳X�����s�R����~��ԥ)�y�ں�H�4����B"(̷wwb���<�߸qJR��}��/R��y��k�R�	��}��JS���VZ>�n5��k{����R��{��pz��;�>�\R�@d?y��pz��;�߸qJ���x�+�%j#e�$�\5@�N�Ͼ��)~����)Jy�p┥'�����)H��3�f��oZ�-��[��)~����JR����8�)C�����JS��ߵ�)JO��O��^0~u�%��[����of:�u�u���dB��l:x{n��1��|0��;�Zz����ԥ)ߞ�ÊR��������)�y��� K��?��~~pz��>_?�N\ME#-8.�T	���\�����z��:��??z��(o�ޱ\5@����X���U@��~I�LiIn]��p�������������?#%<�����&�4>����p�j�kH2�d8�IY��|N��J���pz��;�߸qJR��}��R�˙�o�R�����B"%!�w.�p�j�s}b�)JO���=JR�~{���)K����WP&�uJ�i��Iq�ZEA��	�(m�ۓ۝ʱ f�{N3��;�ɰ���j4��`Q5@����W1H�����JR��>��R��~{�)U@�^�J^�p7D�
j9b�j�*]����NJP����pz��;�߸qJR�Ͻ��/R����Y��_n޵��y���R�>���pz��;�߸qJC�e1�Hh�N��Oλ����)J^z{��)JP���feo�dFa�K�˱\ Q5C���u@��f'�����)K�=�|R���~����H���! qE���c�@�JO���=JR��g����)JP'翟���)N���R�������l6�4ӝ��!�nlsG&��F��$���gP�;�o2N�F�.�Ź������R���߷�(_|��=JR����8!JRy��}��R���(���h(�II�.�B���z�p�(�w�p�wJRy����ԥ)�y�ں�T	�����$FDR�r�=JR����8�)I����ZS��ߵ�)J�~��R���Ĩ��rHຠM
����z�p��~�߳�R�>�}���(?C�D�

)@��w�!��Z)��CX↏}���h��MP&�p�-���"c�7��R���{�qJR��Ͼ��ԥ)߾���R����~��ԥ)������7:���3���,�.�v����d5��q�Ӎ��,�'i�©����?<�b����޷�R�������R�~��)JR{��k�	ԥ)�y��┥�ԐC|JhHa�K�˱\5@�����o��'�{���iK�~�|R����{�+��4 W��֒2#�)�kg�i:�߾��J]�����w�������ܥ)�����iJN�䟌i�	�'$NX�j����}.����Ͼ��ԥ)߾�ÊR��{������I{�(ĒRrK���}��^�(��Ͼ���yJR{����R��y{��┥'�� � <_�����EBȍ������v겤t�<�<�������}���H��׎֝v�-j8U��nS��2��-��Y3/\����
V�^f�`�s�\� �ź�S�]�G7Equ�{vý9���k9wz�'6��+�r&G�lF603�����]u�z�v���k$ӶL�8i9��θ�Y��[Z��IGs�,��q�WW�R��հ9^����{�������)ۓ��=����S�[��u�ɏY0��vܻuϹ�E6�d!!5�]�F�N2&�-X��s��?'%3�s���i>�߾��)J]����4��}���(s�!�O�5��$p]P&�C۾���� (�H�^}����)K������JS�}���`4�y��}�����7�-o{��)J^}��┥(}��}��R���~��)JO���=JRn��`��lb�[��5@�^�{��JS�}���(|�߾��)M��K��Esu$�Ȍ��#����R���~��)JO���=JP7~����)C��}��JS�/~9�D�x�����g�#ɬ8������](n��HͲ^���2gv��j�Zv[���R��}��R�����)JR���|pr�R���~��)J�/�_k4\0��q����Y�v � ��|�о�� L
���A�y���Ҕ?���8=JR����8�)T3��X�(���I/|Ta��A"�z┥�}���(���R��R$�����R����ߚ┥'���B�hFDPK����T	������'�}���)O|׿g�?�߾��p�j��A>?BZ�0�$���)JO>��=JP>��~�)JP���}��R���~��(}�$�~�k�답�)u�����-���n{t���t��.Å���n�1��xsq����'��%):��{���`9��}��JS�����)<�߾��)JG{���l$"���&���H��{�+��@ ��O?>���)JO>����)J{�g�o�R�={�fe}�j2ٻ{7��[��J�}���(|�߾��!��En7o�#��S3��	��{��������ZA7Q��d��j������WH�7�ԥ)}����)Jw��p┥'x0�z3"��NH��\5@�+Vo��R�>���pz�P�{���h{sޱ\5@���"6�tC���\�\�6 �v�\��q��\��u��'ZN�m]x;Kq(�-C��#��MP$Ug��^�)N���h
��}��R��;��u@��M{4#�d�Ȋ	ww�pz��;�߸qJR��}��R�����)JR���}������W�N�ַ��[8�)I�����J��~���pC�����)N���W�ht{����R!h��U�TR��{���)C��}��JS�����?@ "HBI	���	"*B$�H$���1Š�F�a%������p� �D�0R�j4�Κ�/��T	�N|�n0�@͕�f��)JP���}��5!�����8�)I��}��JS��ߵ�)JN
�n�0�0�#idD9	$:0����n�7
k���z��2�*^��;�6��8�v�o����ԥ)���ÊR��}��qz��=�=�\��u)K��??8=�MP��_ZH�b�6܌�ຠMP2y��}��?Nb����ߛ��(~����R��{�)�b��h�+�&�P�crE%�����|�
&�?y��pz��Usz2S�Ͽ8pR�߳�WP&�nF�%e�b�2�v���Ͼ��ԛ�%;�߸qJR�����R�������\R���������"Ġ�,]݊���}b�)Iן{��JS��ߵ�)J;�ל��9��{���*��Ҵ����\��$�$!
&I`$'��`�����%�@�eM#��%怬3@Xj���ȲC�ucI�fa�e �(k@ja��H���"I
���($�@"�B�3LаԆ-@���m��d����$��j�&�x�J�6ăA,�u�[H�N��w)�]�F���O(L�A�l	QѣF$�LДD[���JT�%4�TNc�4��@�RĐ�C��aq�� ��چ9���%!<��;-��W�]C��#)f�a%�$*�LZ�:ܔKBP�%1)���K���R&�Df�/�N�n[,�Z7؝A3քp6F*'�d�LT��$��"f>۽�h�� ՊN��P@�C1$�
U2��8CDBHI��0J��K RK3!!�΄��ũu�ޓ�8�,�����z�$�߇�	�d�AD32%AhM�+B�P�QY��J�e5*i�d+�"�)o;ߓ��^ټóX�y�۬v9;���й����A������q�B5�[AF7�h+m�=�gc5�ݶ���_�����h,�<�� ^����xl�'\�M��m���l�m��n}��9��l�U��Ș�v��F�2&| �3���ڪBn���᪐U�2�+ɷ́|��w[˛n7<O�h�$12Y�3�q;�8���f�ݞ���ð�ns�r�gr�dv�[�m���/A���Y��������g("�O�up`���G���«�q�U۝β�hq�(iE�H�]t����#��KQF�J��ji���d�Jrj�I���,��{s���T!�Ð}�z�ٖ�I���'��k�l�4���Mhth�������3J�G=�PAv�q��5�Z�b�U%C���@�);!H1��W`�����;d�v_%TF��V��!O*!0p��V�v��vj�r��=��$��L��b�h�h-Б5��P�H�b�����=�2�'ě�za��nѱlt���&Ariv��du�كO=&D��WSpunB��mp�5*������΃�������v�3ݙ��P��^݁�<��Q��v���8�4�HY��y�eX8�vѪ�t��kzs����'USU/AƈD�Pd9�ZGd�K�ڔ�W�B�gD5�3��ԒѠ��/ EVW���dv�Hq��^/]Y\�:���A�e��^��uV%�]o/dL�N�-����cZ�7We���MqVf��E`�3�婪�X��%&��!L��J�nv�m���X-c��݀��/'�'l��.��l�����;B�*ѹN�P*�ej�aXj��F��sA^��L�rn���K��S�^`���t��O[�f�}�m�mQ|����휾�ԓ']=im]S�ۋ��98�m��9�T��9zb��Z����nګ�,��H�i��j 84m��ֵ��l�����
��E��A�ȁP U,~�����w��'�5��u�v)ڧ�v"	І=!�<��S�
���:?=�NHܦ�H�"r�$� �e�w6�]n��ΧK�:Zё#����Ҕ�J�{�f�#rv^fx��t/tm���X��o4[?|��\X��b�h��~+�jB:N6�{J�bƛl���$[��'�������Ѭ�qūuuI�;
8���\�Y��^�8ל�l��W�o�7.�wKɓ�����g�lʦ2��EP�<kp��c���Q�#iWP'�
eۆ�������
kv�ۋ&�BW��n^]ۯ;
Q����q�]�P	�/��&��'/m˴v�f���Uj�4=���\5@���7�┥/�����)N���R��{<G�o���A��,WP&���|�cJP�{�����R�������(��o8�کV���Q%i�� _$�@�������_y?n�y�߹���~�d=�(������*��4��# ���`=N�}��@]�S3%V��6ڒr�o�yޠ��]�g}�|(;��Ձ��o���i��A(3�5��S��h(��,��m���QO���.r����2'Rs�b��`�f� ��mՁ��o8x��jQ��RS���ߟ}�����Ѡ�	D$Ү�  w�~��,�߷��	:�|�� �>��?#�4b�K��3������|���fz�`
~�w�>�G�7EHDڕr�(��7��]���ݜ'�*�}�,�~ψ	}�PH���{�B��u��}����y�'�r���&��􉌐Dq&�7 cgc�$�rk]a[l<s�Gw�3��m*$�Q8�^����u`��y�DG ��)��н$���qe�]eVe�4�2 �Ot�S���(�ީ���lHM�MSm�$�XE�>~��A=Y�vz?�]
d%u~^��p����Ձ�W�kbJG�H�8ʪN��`z����	i�`}5�O;��FO%e�b�2�vI���t
G�Ց�j�{�)�u�l!(tE�Eđ�8�;wn���R;u�1�����:;m.�w7n��ە�J$qSD���ws�wsn��:�{�}=N� #��'z>�;Ժ*B6�r���7�>Y��.�V��ͺ�}��n�	B#
jNp=N� ����L�o/ ޴�@"���qQZ�t�TH�q�?,y��p��Ͽ7ʺ��~��׀~ ���C3�Rm��y����\����?�P1J�u�.p��,{sy�1{5;�~�|��V��uJƷQ�):����=�m�W:K��.v��cu���l�14��MSm�$iI8}��p^�v|����͖���TnD���ʺ��>T��v��h�;�7����X���l�����_󙯀$� �6�@�Rs�(}Q#�������������&z߯ ��Ƿ@�Rs�A�/f�����I�HF�������oӠuR~����� �ΑZO��W�Ӫј��h�5�v8�����q�ԉtc�������7!�7kk���$1r,�-:�3"C�^к5D8�Ye6A�]Z6c�Cm����T�q<�dF��^s�Sԣ��.h�SY�e'ks���+����#�x�H��I��@��� +ά]���ylq٣bө�{C�6�'������-�d`��ZX���m�Ի/J�Uw�|���~g-�@��&ܴ����;���hgx�e�!���y�
�5�7mnݼ�/[=��]qn09�i�ݍ��%ڐ�������������u�1/<���9H���}�N��7m!F�qY�M��� �����{c@�������P1J�u�-��͖swy�;纬c͛8mc-�6��n�������v�� �T��4;��`o���8�F�Np��܎G1<~�t���>M��q�N�n�6���g��nx7=��^�M��֣��֍c[���=�vW����t���\%s�U&�@;�� �6�@������l�#r�Wv�I9����	�j������v}pp����Oq���� $}����4��0��Oz���;�np8}��u��w�8�5���5$� ���=�7_ ;�����{� �?Lꫨ�����97W8U&�vd;�� ��{�}�np�?c�Mҥ�ۄn�#���7����{Q�ݜlnۮ"66U����3����Y�W��Rw�|�{�.�s�uRz��4���ؚqG$�,���s��DL�u�N �Kު۩�� C�vP�#q�'8Pw�=�����F�([�����<�@}�
-�4EL"��R+�~�|ā{6X����g��+$�}�	!�QFʒ5	��|$S��>���Γ��W[�܈�O��~;+��ɥ�@�A��7)� ���yv���m�������ڰN�t�mUw�4����I�߫��h�w�(����'É$GC$��ך�;�������{n`�U6�EH�+^��k��,�m�sk���U�sڄ�֐�ʑԸ:��s��L��x|���:Np?Dv9�UUB���UUW;���Ny�Vk�@�m��nI`~��y��׹���{�gse�P����� ����NCW9��宣�rv�:��7V��͍�{N�,uڬ7�i������������`�XQ��o8]Ҋ�zD�jH�#�6~J�;�U��Ot�;�>�El$I�5*W.G�$o�e���󇣜�9�����>�y���Y2���"�ª� �|��z�`����X�>Ku��H��Ԝ������`������}!�#�����r �b$�D�1ĎD�h2�L�#'F���K�ɺݓu��X�zz�#�q:�df�m�Y�uЋ��NS�n���=�������ݷkhN�P�4]��UN]�WٰM+m��頃Z�"�v���>]�C\��D�[��մ��U�M����.�d�^�5��S�@�;��9�-r�k�n�����)�L�Y8˥{���9	Xw��2wD٩dcl�S�w~���Q��]���w�΍��u=��؍l��vڷr@����΀��IE�LHt�>������ ��%�{��ۣ�5{5�]^BFkHdeEM[v��ـw�=��:�6[U��&F�dnn�m���Q)$�3��� ��k��Ż��;��`s��n�i��2G!��;=N��� �~J�=������EM~�M2��RTj8�w2X;��	6�@n�s��<�`�T�1]�;e�Nu>ѽkm)�s��c��v˷\��d����ׅ DH�I2�PNܒt�No�K$���z��i^ߠ!X*��K���)�,�w}�s�����U@W�2m�/ =��@ߒ�=�N���IDt&�� =��`��,�<�}�,���yn��Q�QDT���� 7� m�l�Aާxv{.D�֐�ʊ��\���6X}����:���<���`z������ҤIC�:�zlƟNq�;���ڀ�d�=f���}?C+��H��(��R(�rX��������@RU�G""6@����
z�N&��Ȥ���ٮ�ՙ��9��`f��8�VS�1�E%!�� r����ߒ�2%_���RmU�v�Ľ�~�}�z���c��ߒ,ZL���8YG'�u)�����T��L4�4��((>��P��)܈a�a���I��U	��(��v�7Xi4�BVj�>�^���@�@�4����B��`"k��6�.*bv��8�EY�۰�hu���w�lP�DG   =�h�ҁ�4��
�
&�`���b�8Û��M����Ç8��C�9�u�����E�߭��;)����$�e��U7[wu��[/ I��ݤ� r�*�=��YL�Su�6�37w�8���� 4iV o�^��G!u:�_����#����xnR��^p�u��m��,����݁sA9{���F�ӌ���m��~��J�~J� M����s�D�G�8�Y��
9]̖n��{�5X]���T�ʊ��!]ր}�� ��mϣ�)S����Xy�c���ӒTJI,�ۼ���V��vʡ�q�۲��ר��8�F�q�py�V�c��K	����z���I�?�q��LHɰm��.k����e��v��ъ�p/[U��ݹ����TԊ����$�\�2���>�A�<�`z��H��@��R��zu;�m��i9��� �� W��!����p(�n�8|�U��1���d�;��
ObR)BDm6�� ���V�;1*;�a����߻�
�~�>�Q�D|���չ��z"	��� ߽��i9�?D>G9b��hVQ��&8hE��L�ɈH���K�Q��3����)��+� ���.�]�`2F���7��{��o�NF��k���Yx�0���ppNL��r���%\��/�nϨ���$�׌�2Ƅn��=������)l^-���+ E�aZ#Y֞zΡ�m2���Ň�q��l/�ɹ��������v{�c������ђ�
!=�H��(c)�N��vZ�,�2��sm�����۶c��ݞ�@��SL[�]����}��x�8~�9�!Σs]�=�β�����Ў׬]3]�Occ��m͑��-Y1��s�tE9t�?��w�M��;�Np r�vy�c�Q���5"�I%�����s�;�Np-*� ߺ�.d�����jY����'5O��e��(
)}�,���s�v�QYQ�)���57s��J�~J�s*����j���e#H�Jc��Gˑ��ݖ��M���s��Ҭ�̬���l�5њ�,`�u���A�]n���ڶ�@����(M�6����uܖ�7y��9 }-
���W�u��sM�#H�9�Nc�+C��
�P��"9�?N_��~j���-����>)���E�+ 鹎�9�d�=�n�w�5X��E,ԕ22��Z�������7o�K�x@�-g���3�#�܃i�ԒX��� ��9��W�����P>W		�<�b\��Ǹ��P6_m��uiG��g��9ۺ�[ur���:%�nP2G�_ ���R;I^ o�W�u��@;�UR艙���$� ��K�w�,nn�w�5_�]ܠ6��2Sr�˒p�ݜ�Ͻ�C{	�1�RY��$ @0�C%�O�\�o��wے��h�,��:��]��ot��� ��x ߒ�����=jG>D�$��^�v�|Ҽ ߒ��7�y�)�d���U4:��㝸ՙ���8e��+�7\��������+�)a�C�:!�#-F�q�$��v ߒ��7���)��=eI�)2TT�+���l�=������`��`g�T,�ӂi�ԒZH�I���w�ϚW��W�v:Ga������9�p?U*Ǜ�� {������?D(���A����{�|�F��J9�rK ��K�w2X�n�y{5��7tj)(��S��vc��c�l<��V�Ƿb��ݫ�X��ݻ7���}��PPr�)����}�,nV�8��_򷬭Z�O��ܠg�~�$7ue���i��" ������ 7�OZ�B��RNW ;��,��Q�d�ޫ�i�G[�T��t��"��If��^O1�;��7y�*���6X]����I�MTT��Z�S��������� �ZWx�l^�JD	BUW���3ݿo�/H��ky�ўS��:���l�N��8�W�U�c8�t�N&N��%�]�(;x�xxF:֧��ۜ�<xwg�]Z�ٹ���b6Pv��u����ٚ�9��,�I*#�t㫸󓧗Z�2�S��Ss����gnq�7=�r�����~9>�qێNԧ vwa�wBͣ�Q�V]�ܕ�&n��F+%�ۤ�qm��eAHI!
8��.� _ߣs�Ş����z�Ԕ���;m�om�^��-��n�Z,�Ʊu����{�CcזּU�Suw�����>��X@}-*� ߺ����v�#���Q8�� ��f���Ñ�D�g�� }�� �{�"9ޔCTT�P��C��[����J�=������`VWw(�9L���ܻ���>��xZot�����UW����3��m$��jT$�X�ot��� |Ҽ ߒ�~j$���-���-�]����g��o���f�hۨ�"綣�.�q������n�j��;=N�#����y�D@i��n��oj1����7�ws%�J���#����9ȝ�O2��}��>��Y $�[���4"ҹ8A'�7� �MR�~���� ]��%**��i�5�U|{�n�W�]�չ��Ĩ
=ɲ�=��+�#�"�J9u{�}=N�r#���@>�w�|�ݠ74�5�ut)H���H"�ͱ�m�n�ե�%ƴ��s�z֎�g�=��W��z���}q&�"r��v71�;�{sw�+R�ͷ`ewr�j4�BS���#���s�Zot������DPW�@�R ��BI%�����E�y����"�RDL���1��9�d����'V���C$!*1�9�>���f���t��`�Y?� S{���8I4>�Q3�M�]U�KJ���U�i��>��XI�ǚħ�ː�ۉ&bU��0gW8�v���5ۂrlX �\v퍷\DlAK�wY�n��'$GL�q��͖�7y�:��ՠ���`gZT,�7�r(�r]֛��DD�"N�~���� 7��>��P�q�#���8W�]�չ����w�,nn�w�mҎ�JQ�%]��X�U�i����)�"4H�J�@?��x
�Zu�n�:;�|#Nd28�r= ������DC�����OՓ2}-*�8�Q䩱S�"Sp)I���p6�G�OnC˵�@�N��`#�ɷ	�y�m}����:��K
=������`ync��x��e���3jB9�T:m99�:�����Ҭ ߺ� i����LH{�*�"�&�(ϣqݤb�5�}�,+���������u�+6	9 ���2s+C�2������@�z�a"�8�5�'q��Z��m7"�G&}24����:�;+�� 7��"-gt��V]�IjJ�3��9�� �(���A�'����	�G���3|()�Be1*Z��y�tn'�IN�C>fq�
�Fo�xs~�������F{���;5��`/��$I	 �@2���KA$D7�h�ݎFa�ZG0ӂ��:S|�@�U;57;�3P'e%<�P;�}h���͖�v�f$Y�b%ۈ7���G�@|M����:�! �[bT���
lU9�k�ɳ4��@HJ�=xl�� �%`�6�w��(JD�9�(Ľ� u(>gH1*�O-t�Ѫ��.�� ��9�9j0�gy����X/����~w;r*JI�IB� E��)�Vdٶ �^��@V�9�r���:ji@X��
V�P�."t֫�y�v5�6��Hm�s����<��[����2/�*����T�����yմQ,���fr��e�4�[q�W[U����*��y��㮻�x�:;{���Ĉ]��u���D�b�"�yݞ���Ohb�.��;{FʩsL�ڦ�0��:� 뭞�c;ig�j��8Hۭ�e�凫�;Ǹ;uW:
.��n�p�J:u=��6�&���� VMk�8,ݝ�KR���Q�9��ZU�Ynp�����+��v��Ϫ���QN���p�nIn�ű�7n�K�s�g�4�<��ˉ�P4�,��ԸҀ8�����c%W���j��*�9�/T�UŶK,ʡ�	�µ[X�ii`
��p��Z�^�]���*��ɓ%���_;m]�;�<�$��"L���E�Aԅ�e�!��S��L�+&֛���瓪�u)��K������G6���z`�ĭ
�]�.�����gsK5*�`9���P�[=�q�n1H88��ks�<��y뷵�砋�ݝ;2ݖ�X+nXV��傕�;��;۝������t�\#��[��2� �����S���z��Q)<�lu2��'補k��J��)I�fW��2�<���ä�t]�\`B�ʛj:+m�=���C��Y�Nլ�!I��wc��]�]Q�������JۧS�gg��%�
�����:�v���f,Y�x�@Pے slIub��(�:;cN��i%R�W/2Ɠ8�5E-Hp[@ڵ��`�6h�g�^��q�ʋ��̦M�o8��m��R��8�wfPvh�
��㓐ݎ�r�pd7���.���Bd�n�G\�:��-�u��x�CdZ��VI8�Y�2֩�UUTQ)��*ʨMm��:*�Y[q����@�8ݝq@T�E�wPK���\f�"���Ϟ$����C�� t/�@lS�N!��'���o]�s���
��n�E�h"��\��"!I"�8��\c���Z��|���LcZ8����/�{<~7c�Q��A�;�;l�et�n�9�o>:��A�9fӄ���Ҏ�ڪ�1��L�p󨛬kp�uն�r�+8{s�h�;q&٭֫r��)�ݣ0n9��/��t6��
��!$99�U�mnȷOl�y8�vԙ���]�A�0\�a]���,�e���S�g���t�n��?��}֒������_k�ɋ����n��)��z.�;![�#���G'������`yg��@s��`{w7�(=�
ͺ��H�Rr;��� 7�������� Q��6�ܨ8H�>\����=����<�`yo����)e2$�R�$� �i��i9�ɓ��� >�U�A�j�fԂ��P��'8��U�/-�v�R��:�{���>��_(������釭���tm�:��7m��=�m[c�^�vW��=��ۦ X��c������~? o�\`�oc܎} �?N s�;�/|JrE
`�"��	'��K�kC�t	B�k�7��󄗹=��'�]� RG�Zx5i�JI,�/�}���j�<�1�;�,����PHH�ns�G�o�aF-�v\ﲥ��7w���7m�i��MH�$�`Ȉ'~�m��i9�;�f1��Nܜ�;e���ѽkv����auv�v����AN��\�3�&��C7��|$���� i��ݤ�܎lH)m��P��"Q�T$�X�wy�;皬,�v��%��UK6��t�NNuߚ���^g�����t���2�w�^�G����f�8��M�D�D#��������t��Xߓ�ɷ��y���.ְ[�'!"N����}�^6�@}V�p 줫 ��B�鵨+��$����cY����Ύ�8�hd�,L��|��2l�,������۠}�Np�J�~�.���RD�$$R79�}3W ��c�w�,���?��G��ڏ�j�����9 )m� o�W��9��?{۠uS�������Jr��|��6XG����uW~k߳�����\��>vV_�~k�����3�V҃�P�I`3sy�;皬	��{���?T=����r�"���,�um�N9C���YMh�b�����֍ܙ��-
����i7/���qnk���xM=� �8ܢ&*�\�T͗E�VIŹ�� U �=���O���s�w�5X���	�8�Aj���y 4��.;1ȣ�I���� ^��N	��q(�777��y����c�>���K3��m&�*		�Np���=����Kss_:��~�����A���?3Zݹ�Ø�R\�x�;v����:����[�Is/�5�/[s�tM�ӋY��,i��n=m��՛�bػ����zzŃ!u(�@@�G4m��n����X6G�lt��Qn��{�gk:�r%^:ٹ89#�H�5d�(��nMnj�9^-��L��٬�n��j�G@�glQ)E	m�m�	�Y��g�M��)6Ѝ�P�!��.�a�vg���n˳E��[�G��%���F�π/�!�p�2�� �:r���R.��<� 7��i��"9������=��,�!��'%�8I=����P	����U?N uu^��p7��&Ur��T$�X���#�6ݞ����8I<��,���Z-��N�(Pg�� k�� }�� ����7(7�
-��m��vIŹ�� Tyޫ�i�v����n&%�P]��F[n�ssq�絵�X���j��q�N�W*�ٲ;�rA�K�9I�PZ�| �e�����>�'>�s��DDH)�u�4T̷wR�r8�rY ���s���ô '9Y"u� ><�X�U^~9��m�RR���'8-�����;"G;�7sy�=�ʔ����Wu��Dp쾪�����{ߤ��Z�`mf��ڐ��' ;��g��DG�O١e?V uu^��+*�mqoC��x����\v�j7DGG ���'cs7����\e�^Ў��]j���������:������+�>��u.ąIM�NN. Nk�+�����N���yI�9ũ|���s�
@O�/�_H�n4����+ �ݖ�d��Uڪ�G�������u��uWk���We���n�NA��J�oP|{fˠ6�wy�=�5X+��<�������$�EQĤ������_{f�
<�v�fK+�F��HI�6�H(�ʩ���DX�tƆ��F9��g�[���tn�2�6B�PHH�ns�{j�<�1Հs��t���w�T��6�"�R8XY����rd>I���{t��d{���I-�{�WSUWe^��h[�� �oxs&��f;������D��T%��`1��>Jـ	%x�/��8H��%x��f�?Q�T{�w�������D��&nNp�MIԕ������	Q�&�����8n<����u�,��H:s[᳌���2Z�gq�:�%��˴3��u%x�����hJl��=r��	�������� ���p�ջ�d�[��� R���x���$��$9J9R��?s�ufk��URX�u�}�,�䶒�>		����D}=N��J�~�Dr"'������jS��iB)9�x��`{�r9��w�y��� >��`�/�c���U�@I��-9#p6�R7�����#�ʍ��Z�����7m���3�7���=��V���;<�x�:˲��vۃ-���ɶMjP�qtvj�����;]������9�Q�����]��������.�8�h�5ۖ�y���5�϶��	�P�gY�g=S����v[.�iv89�r浲o,���EO"[k�x��W;]+*auδ޻M��?~�p��
]�O;��4D
4�aI�q�px����Nڮv��9��clwWn��^ڶG*D7*'��� =��Kswy�:�5� '�$�a�ۦ��2��%� �ot*g����X�꼎r �5�-��I�n�7'8�͖ybU�z9��'z>~�������n��c����,,�v��X���_W�s6X������NSq�����9����4�� �'y�0vRU���;������k5vޮ[�s/T�`�ݻm���`x�\�գ��z��k�W���d��2���W3wxM���w�U�DDF���aF��RnR���H�� ;�o���p�dq@�)�@  T� tUV�)�vI<�l�O���s���PR��QHRrK �w\`���9�Ots'[��>J��r�Cr	�� w3e���[�p͖���s]����ۦ&D�D�G.�&���DO[��
Zu�ޫ�=hF��ZL���lFRDE4PXތq�}۔�S	uֵ�㶒݄V�n�y����V���&�ܾ�Vf��=��9�d� ����h�1}�$#q4�F�M�`qwʰ�ޫ�i�|���5�ڂ��&���.�L����w�4��?�Ȏ>sO��	�Wqwi$�JR>�\Dr   ����i	�)i���c}~�����	�L�d�8Jxu���@�|w���й2A灰-it�|��o	:�˚�fm�� ���52�10D�ݔ�MK�<|Sf7!�m C������P@Ah��i���	�]�RC&,E�������F��\�:⚚ ��F��P:h���sG��X=
T�Q,#�s�����{���P�F/ IR�
��{����C��M�l_���)E�2���ֵ֩Z����t	���(NÂbi &S
C �(��*���E*(���Ѡ�FAh�4l4h�T�H���QO����v��� �a�W�*�H
D= Ca��p ڏ��=��� <A9"����Y�vI���d���[�7q'%\����9�ȟ��ۤe�V�]U���X{05'JT�"BI��K�'X����u�A�� �i�(��	&���*B(C%S$�eB���Ou<[��wY����]�*��z���"��� 쮪��U�4���>��`A�b��
nThnA>\��{� ����Y����}A��eJ��D�D�G$�777� ���,��d���,��]Q�)>j��Ns�U��ʯ=���<�|���A��H�@eUPܠ.� �}���	'>^#�Hb���&�nK �{%�s��`nno8�w��?�P���1+�RD��4�^�7^���k��k����R�o�Z64)�ubxv���RE(�������߮X���ՙ��=��`s<E��EpNFAM�� �Ot� >��`WU�����`jN��
D���s���U�+���" ��^ �Ot� ��*����&��p=�DD�i� |��ͧ�bB�WuwNw�����*r�ր|��܎r9�y�����������U04/��3D���܊�gQ��\�s��tHE�qh�/V��Y:�0�"���i\�l��t��� U�.M����9��O�O\�vza�Uπ]���<p��&̎�w��rSr���Y� �܏�FwSWg��yq�.�&�R���u�љ����nطTQ���N��%`�i�']���-N�5��uO��7��4���W�����ڨ�?:��QgZ�Z��V�6kb�>��8w/\���}[X2��[t!J�=s�w�{���i!t�8Pl(!�Id�ٿ��uf�����1.�d�;��ꍐ�I�T"��t=N� R������������� )
)���?	�4�Q��9i� j����~��~�O�3X/�~	Ƥ2-]�� ���K$m����Q�)]U�w�J���b�#�'%�����UUU�3]��=��9���;�x���(B%F�6M[�9�5�7>3j�ˋ��x���;nݓtt��쁥*S��P�)/�b��`j�c�]W�m=�GJ$UH�&�ԅ�#�O���>����)`�*�&#�Ϣ>�#���~��/n��������$$Cr
r�� �se����=N�����veFM�Y1Uqe���~��?}�9OՀ9]U�5T3uK$�G��>�Ĥ��M79�E=N� r�� 5u^	��@[�םr��'L=��\ݰ�<��!Ən�#�ԯk������ ��]F�q�[� b� ��xm=�9��Y �y��C�HIJ�]��畲�i��� �uV�w�H�WsT��Ą�7w7�(3��v+�]|/߿z�}������׳��=��)E�w7h�)���J� ��xmo8W�2�mA�E���Ş�`�� �{���X�r#���)&�e{rs�ӳ6"u���ɍn�o`�1����m��=:J�o#Uq;||�o�'�ɩ�^����~�8i�� 1uV��: �D�I$�3w7�+u:����]W��Drf�~����s7|���*�t)��+���r ��xn����*IM�B��a�WU`���i��?A��S�"��UM(~��}���5ʏ�m~��}Z��)EZ�| ���(
����;�ٮ�՞�`{��4H�1�cM�N����0s�۰�+���Q�i��d�|��;D{ ��B$�'wn$���������u�CN�Dr�r9�����=3�
�)�#���(1{5�T��; �{/ M����DW9��q��\������=>~� ��� �][�zRu�|ۉ5�5*E)���o�A�ݖn����«�V{���yE,tTb�P���6���^ �uV jJ� � �B���|9b0�-�Q"����.��r�;y�^�n�ܜƗ���L�:Ma�9ӵ�5�e�Ӎ��ˇm��)��`y�v����T��A��n�l�M�Rl<T�`���@��L����ӷCV:L��A�u�G[|t	��T�����<hSdSj�Z�B�ֆzQ�H��T�6N��'Sfwn	��e��7N�8s��lJ��f�m&G4��1�G����ʧ�|�R&��$�č2$�;���nwK۷��u�=�'�<3Jyɝ��~�����HI>���ܾ o��u#�vޞ�aFn���
6��$E7Dn<$��� ��xm=���?Aј�K��%	$R��v����KOt��?^�mV�RH�Ys5d��\�����p�K���@r�� r����R�/g�R{C��P�);�)�u�>�UX����{�8e~8ϳ�~sOOeM�r&D-�l����ۃ��\ nzݶˠ�k��2<��;�d��%yzb�*� r�� 4]U�&�� ]N��Pn�JT�G"��o��ݗ_��s�D(�s����n�}�;����3�
K
*SJ��K7sy�'x~�#�S-:��w�}��Q�����LŕW���Drb#�-?^ s�N���	g��� 7`���Q�GWX��X@z9�p�s���w�?y�t=�,}^��T���u R$�9 �]��ܺ9�4=Y�a9����;Aˋ����Z�:��*"JUj���͖3L�p^�v��6X�э,�MĜ�$��}Ot��D@�� �uV j� g�Z���A�G���l�5g����;P��@�ց ��k��.�Y��*$�@&H�h�$�t�HJ����"'꟪�~��s�,翛�� �V��HSrKDD��u�4���
z�`<�3@�$ND�r� ;����U���LDDDC������� b��[���K�ыz9- ;�8�9�.�k�\j��H�m�.<9��l�\evø-ۮq�Z��0&��OS��ꨈ�s���� ��5|l�$����79�1{5ߺ٪�V2j��6�w܎DL���+�vC"���u`~[Y�����,�����Y�sy�:�5��w),5	O�QJ#'.��#�ͻ�i'X�܁��3�X](-�׿k�u�3ZO*&�NGNK?no8�f�Z�����,fV�����J<�Ggsd*:�}�8ګYюz�v�x�[����')�>�P�)9f�V{�jJ󜈈>M��� EòK�UݔU�d �uV jJ�᧺��eW�Pܠ+4	Q�	$S�-���0�{���`WU`�
�D� ��b�f���?r_����[�`Wu�G�@P�x��d���GʏͷQ�W���`WU`oR�6��͎�5{?���c�I7ww�s� �IR��0�)��,�32,�3�01�hߦ"kn�WR�����CF���ݤ�@�])�C��'��l��A<���b0�0dƔK�u�[S�b��R�P�П!9�Mf�ȱk�D��CKEMD�����fZ�Y����f�h(gR�Á�FAI��)��,R �(
��(�	�)����Z=��C#0�H8�R�cT%;:��;W"��# �	�Ĥ�!η��`�%d��t�0�JQ�� ��B�1d%Ƌ@p�iLL:��5�n>��ۢ�M@mT�����i���^$M[I��\�`W�r��`'\�3�Mr۲�m��W]�I�͚�tFJ
��Bkh������Z��qdm�a.s��p�>-��n��F�5V���n�Uq�Z���]r�ubֆU�}[��H������˺Hӌ2e� y<�۫n��waMg`�ܣYgZ^�vL�����Vy�V#�[v��S��*��j�R���Hc�i����6rn ��t��G�̻4q+pZ�2QW��L���&0�Ғ�hs��4�ݬk�oM�ʃٞi3=m�P5�]@x̓���ݢaݻl�y8��ې�Um��%:�O=e���ݪ6�rv, �V�m]r�B��hVU1��UtJ�]T���*�[l�2d��H��$�"pClڱBH�uʣz��Ǌ ,c3j@1������Sa��.9ݍGn��rh����e�^M�Egd쉍��S�gz5ȼ����X��E�ۚ2��T��� ] V�e<b��Ҵ+4�ca6��ru3Z���N�Xzq��g�;��4��3ӽh���e����z;+�#l�7���g,�4�ЅX�\�l�B�� Uc/g`�P���M���A���uUI���e$�+��X�6�����e)V�6.H����Y��Ci�-��TQt�����V��.{d�i���òMQ�d����nGv� �.�ޮ�j���a��ɲ�@Tc{�]�˝�nv&�n-��R�9��&	�ʻT���M��n+5k�U������h
��Y`Hx-\V��m����iM%l�$�vɺZ��9�jC��UU�ճm�$���m�!�J�+��{S��fY�3Ʃ���';�$UK���B쳠 �v]���j�7]��띶��d��'�CQ�.+]�qt�*s�\��UT T �VJ ^��t�S�a�fj��#T�/4��V��U*ԫ�E�ѝځ8�����j� ����~�{��v���*���}�ઁ��í���!�Jx!�PMt��
���T+�WÐ�1t��^&��F	p���:[/�n+�۲~o��|&�d�������D������J\]��v�cT�U������/l_ξ�}�P{Hv+�|�["f�y��{)�&�����:���Y�.m�]��� ���#�ceE�����\Y����cNOc]�v�_x{� 8#���1l���7�)�N�ٸ+@��힧�Ss��gt�g[��|s<�۴��Y��7N^������;���T7��CE��Zxݫ���eC����c��9�c�=�-jˇq�s��%���%��m�����X�J��Ki��s���
[�`AO�д?RRD������얃7sy�1n�5g����$�4�TMĜ�������y�vRu�9]U�ԥ�sI�$=PC��ⓜ'�@Ph��X��u���^1�-=�`1T�%@���՞�`�d�i��I�=�qSg�����*�a�+!�n0�h���m�ծƱ�� z^�\v��\��%F��H�n[�svX�Y������KN��}��D� �����I߽��?	@� *�pK���K"]]�wԁw2]��H���T�.
���$�;29��¦`ޥxm�8�U�Ԑ�F�IMFܖ��; ޥxm=� �N����PJ�a)	�H�q�{���O�@P��{���M���r�� �G!��\���pT�7h�<+��ѣs��<�'I�iX�y�M�k��s��=���J�j1��8�rp��s���`j�c�y����*�5*$˻�����.�ٗ*�`����M�� ݠ�SH�EI
�I`fc���=�|�I� I@{�!D���SA�"蔎�G9��C�"9Գ���n�|��Z�3B"5$RD�r�����3w^�Rw�vD�� }��D�8YS\�� ��� �N�)*��d�7k�}��LuDBH��&=u�Ƀu�q�w%Vy�<`�v�X�'cp�h��ys<�*�t�;��� 7�_��E�����8_�V�HE#%5rXU�ԯ M��@I��ҨX�"M
�]��svX����F���,�}����I+*6�RG&K��y��ԝ� �%X���.@��
`'��ϥ�OzO�4����E�"s� �fˠ9�2>q ��,��� ���ߨN�����!"u����wm�B��'a=iKv�#s�24g��N�9�
"��
nI`j��`E�fN3}���{6Xܠ3h�L�T�5˖�&�=ș��n�&�xIVz""#}@=)� ��R����߿~�
�N��9�G9>��`�n���\�%�Ur�&'�]9ɔ�� ��� 7��G"��?n�G9�����T��i��I���d��U �{ӄ�}���]Uy�o�~��B;�qF?L1;y������z��e�R��\�"U��X��#��ۛj��E��MW5<��Ev����U���#��s��]j�&�hz�G�1s��l�;V7V��tdyH����Mn�f��v{t�c�8s�C����ڨ�"��9<l���n��}�/m�IƁ���q�a��s[`�(]YY�]�H5�]k"�{K`�írNVN�9�i����� �Qύڕm@�$�܉	�9 ��3a]v�Ǵ��Gn�q�]��6�b��G�#|a������˯ ~�� M��ԝ� �{��4���I�9I�,�����u'x��`�+�:�)�5ħ"��pٛ,^��+���R��;��~� � a��j"��
nI�)�]g�C���?{ۤ#�T'x�����$r5ۖ��͖]ͷ�I� ��u�z>� J��Q1L�uW������=��3�rMz1	�or\m��\�z6'I' Q�MR�P�I�;��~� ��� S޺�D`�+�>n%��]T��"������|:
� ��Lw��{�`�X�~�p�������M(�v�s]�G=�,*����p,�v-YKZ�!qZ���n��7�e'X
Uv�`�L��̉D�RG�K���p
����3]����V�fK+}���C)4GN'C[�9�W�Z�d	�!kur�F振3��m��ā�@&R�9C��%'�f���� 7�E��u=�:��,��\��'�7��
��HU
=�zXu{ۤe'Y�Drd�\ ��E�\��]��^V�uǽx���/���"?A���� �?�: z����Y��z�]�~�d��'B2��Ld!1I,�(
��u���� ��u�Dr8oR��n�ԾZ�e@@&�� =���/�ٯ��d�9�n�e`�c'ΉM���Θ}˒��+Z��ݸ�x�ݽ]��\l�<T������w>����L ������)� oR�~�{�I� �ʉu.�I
�9���I������
D�7�`��ty#��U��1���#m(��ģ���o��Ǜ,ĺ�k���n�$�����*E
f$��	� )UDDr4�M��ˎ��z��~����}GȽS���f���2���G%�+��z��֞�Rw�~�����?/�m�|�qp &��7;�۰�7[�Bݹ�N�X9�Cץ�;���w��o���8��F�徔���`sۛ� {3e�Ş�`gh2Pch#)T�E$�:�{�I�KP� 7�^3��DU ��Z��[L�I$D���^ǲ���X�J���7� ΐ�ܗui�N�#nK�Vd�{2XQ����P�{�d���B�^i9�77��&� �M��I���� �UB���!v��ifF�mG\�^��iC�����yv��ĉjtH�f:n��J��WL�sgt�n�vv�Ѵy��n��-�P9G0D�ښ� NS(��5!��0�=S�[�Mv���\q�z�X���������Uɬ��7�ݻ!�i�L�7U>�ݭ�rVY�l����鱤1�<˂�F����\OH�w������г��Xe%T�LW����U��L�х��1�u��unv���؛9���Q�k#��3����F�a ���J$�q&����?o8�f��sX��VN�ݚ%�sI���iH!l�7{�vRu�*��V�A6�w�+����7��T��)!#�:�n� ޥx8�DLs�+��t-���p�ߢqI�r� w7e����p
���`qnc�9�(Ȥ�J�B��������*oՀ}>n�svY'�s~N�0Dʑ!$QƈdH@��ˍ��ݷ�,�tvÒiO9�.@�+�^9�F�'9�f��َ�9��`{s7� �<V�IRH�M��rU��}�9���Ε�=A�!p%J�P�@�~ �Z��{��g��u�usw�� RD����6���Q�j���޼:�{���~�>�7XI�i%��5r8�rY4*�Ϸ}�\�u'x���܎DL���0^����$r��)�9�fl�8�1�=�,nf��%���6������u�M����mԻ۶Hn8sSǝ��l�N�G]�V�����`$V�)𔐨��s�sْ���k� =�������ځr)"\��� �7y��'�ԝ�Kn���'GA;����1I,����s��� �{�]�y�����K�H" 84 Rpt� ͉�f�s4�]�ڟ��,�Wo#�� �hxkj��^a�oh�b�nWx{]2z;�W- h�ۭr�\�Rm:cccR ��3�.د}oB��H�l;Q��@\x�=���G�i�!^#����Ͼ�U���Y5�w�,��o孊C&.��@:���m� oR�����o9ăO�	R8�M��%�/.� �� ��Jw�~��8N&&�''���m���7 �[O����1���u��k�ݷ:�����o�����^����n�z����u'~���r$;>�� J�KQ�$�MȢM�`{��ܮ~H3w��N/���$f�'4��!�"�0ʢ����ٞ�� ���a��J��'�P@\�	��"���=�J�{Հ\���{	{v�w��s��~ܼ��������9��| �n��G�}\V߳�߯ �� ��edUE�!oG%��z��l��5�Dݵ\r�1��ǁ��v{7a��pT�N�DB'%��fo8�͖�� �%�F{u���(	H*&.��@n���#�$
}�V |������ i�CdD�	�5)(�ve�X�J�N�'�ғ� ��v<ߛ	�M�|$�G��K$�n��
<�5�[��y��#$JFG&j���'�@z9�D*Oՠ)���]w��_�� @�R*>�"{��HAxp 6��M��P�� �"�UR�s��o�1e7�җZyaۮ-����H[�;l4;��:���%�y�����|�[�c��0��ٺ�b������P��˜��ͦ�iz���판cn�/]��h�rʂ�Mt�F�p���y��pO�����̝s��Wd�\�{v��%�]d	��>F�k�-����(3���e{9ݻd�c�{X��ƎتݎV]��b�$&�V��v"!� ~7tkQ��3��%޷Ggvgn�;7^ݼ��9��^G�X�u�����E6�P�_9�Ll�G/@��������@ߒ��""8]R�@� W-Q	𔐄���5�s�����7��/f� ﶀ�ߥI�ȕܷ�����Ot��Dr��� �� ]���*u �"9,?�P�����2T?V�M� o�^@��r�QeD��������X�s��q�� 7� ���p��K�5�4�T�!S*{h�n�(�s�Βr�;'1e�{u�Yp��Q���iJt��v��,�̖ff��D��|�s�G���M�h�ݥ$᫿>�|���V��`�XPҝ ��0��Y��~u���u��찋��%��q��⚫��:���9t�V�Ȏs�G����vX����ai��#��~_}QȈT�� �� 7� �%���"4!>��; �ݖ���\�+�7�=�;=N��t��*b�E�y�{U�u��w��q�.��s�k���W{k�Ձo�@ `�b�&H�NEw%�Oq��R{�vz�{��羠%�׀>�/d ą��'%�w7~�>�Z�X��^ o�E�#��ޯO%�ua4L]]��7u� �7x~�C9�@d�	�~ov���|����Ϻ�*��͑�8�tԤ(�v��,
7�^ �Ot���L�ڎĺ�S3Wª2����� #��ԞhSs�����}�_�&��"�(����CH�\��t�gI�"+t͙�b�7��8���+�5Dn(GnN������uX�۷���`n�{R�l�12Q� j����r��hM� �Ot`E���&����77eX{2X��� �Ǻ����+~U$r'w9�yz�r"y�y���oۢ�[������S��S!�GB!����$d�}��\E �W�]���9���jD7JRK䗷@�w�N�~���W�}�)bLI0u��TbJ�RDmېۤ��9Ϋ8c���z{�ڜ��v7~���[��˺{i�Q1e���78 �w��^��s��V���"��MJM��s7b�z��$��Ss����ԕ|*��2����� �$�OG#�ST)����Yԏ��Kh#ޖ��v��������|��¦� n�=2��`n��%JJ�4���p�[����"<�����u/n��>��G"$Q�Ce�2ZX!Z�A4!���!�K�BӒ(d�����e�1Y8�kZ�/V6��x�	��]��zݖ�m�����Gev�˵�&�����N�;vݙ��t	���8�\����h���{&����Ͷ���1�57gm�� Z�3qm]���l��3wm�$r���F�қ��w6N��dKiڗpn^z^-���\���S�n�h�Gm[�_j�8�N���A��z�����O�VЍ�޺��DF�k-�zٳݻ]��tp�8�޴��]���W�.�8M�(j@�M� D��nK)J���_�H�n�� �8�������˼�s!)��r ԇ� Է6�ݖaA�0��Cj	B'%��Ot�n�����R0��7P[*:�N��Np�&�v�ݖޥx�p]i��g���EܗU4]T���`�wޥx�S���w@e{`�O��) I��H����V��۶��ݸ:I��{[Ǯ�:�O���|����7w�
7x�S��۬�G 7۲��F���9��M�`w=�uG询9E�}����^���+�3?*ױ*��n��q��`��DDޥx˩���a�*f��&���?��D�^�� 6��.�n�,{5��2��I�ȹr\�M��P�@���� $���EWQ�����~]��5����bl�� �k�ɹ$7�5��p�>^��O������|9�Y���`{}�����w]�Hǻ;\@{1�������6"$�JTA���u@|���J�ާ�s��p����Wr6�H9v�ݖ��K?�����>H<��d� `e� ����9��u��U{����U�FW�[6�9�D+jI���9��n��W��Cb9s��DH���t��' Ԋ8X�g�p
���`��,��٦�9^�ߐj�39�:���������p��k���76�8��ݷ�a��9�%H��H�'8�� �f��+FG9���P@��wə��ɻ���s��" ;�`���[���E����R'"��s�g�i�j�{�vZu��� �vUY�����l� UU����	8���M^����~����J	���G�?�~6I�~a��!I(�9�N/k���]N��Z08j�{ߤ%SwW0s�]vV�Za�\ֶ�i�{6ۧ���k�#�sֳ���=�W���NH�3��.�xߕ# �����G#�e�X�^�l�t���JV���36id�Ϛ{���-�%'x�$�T]�e�M�L՘�����a��s�6�K3f��-{�*H܊H�'z��X�'xz����PBKe ��)!���`{�0�9�=�;-��?������]�ݤ�IBF�$�
^�D"Q�0��I�P/�˺�����.	vx�o��w%!�p56 b���hD�'�)�0�����c$\���h�L���;�0v�k ���4l����j��� ��L�c��M "����6"�3A��+Z� 00qNtP�B�
�"�'xB8�f��m1�c)�*Ű,�A#<ݽ�K��{��Qo^ �0-��.J�ȷh�H��l�!���N��֚y��Rg�\E+Uoan����Ҩ�l�Չ��R]"�u�(��X��س��p�t� �t��g�F�b� y��F�OOXpQ�G.66-��e��4H�-'*��cY�����"a�Zi�c#��ܮh�=����ob�^�-m�&�q��vRū�gHn#b��[j�S��Zv-����e*�B��m���t���C"�����n��}9�67!q@	�l��RR��ݍpUU��Z�n��^&��d&�fjU{G���`K:��g�����ǅG�.6Ό���S!y�=���P����w���Ɔ�9qT��\Ó�:g������Ċ���ԇ1-V����Z#�Yy�ӣj��c�N��K=8�;EB�;9lF�[�E� ���v����-��B9����Fi4;,�JʎBѮ��x9�g��U�W������� Dp���l��ۄ5!����v�vP�jU �=�W�n!�%��q��pc
��3��дnw,�2����rv��6xˬM힠�)!�Ր��P��\{['G9�7n�-/=$��N�ɖ-��x(9�������^���;$�I�l���UQ֣$�H V!6|�u.���kj���/b�C�Pr�U��λ-��-��Rړ!!��.1�s2	{7na[�hg���u�g�w�ibp�hS��z2W�q��a��vqu��[���ڱƞ�B�ۆ��(��;j�2���]*�}��v@�
�����6�og=��L :[��^5Aq�	����I% ʒץ�an��թ�Z�հ u��M���+�͛��],�����J�ݍ7+�U�s�>�t����5DN�q��V�ɲO0R=n6���b�K��齮L���1�3��pWK����@�� pIm�C�N�u�,ՀF�*��uAd�
�^a�����I��BL��s�9k,�튧D��w~���w(�=�����LN �O H�4��#�&tv��B���B�}@{��-�i(���3i�)�#�Xiy�v�g�,��]�^���F-;������������YS�Ä�ʻh�߷������VW�r���`8�1tA\��ׅ�9
�k���f�%�"�a�{weݸ�Ֆ�m̵��8v(5���Ѳ�z�# �M��}�~�vn7I��<��Hձ:�M���.k���k�Į�ɮxy����է���@�&B��#���
�C��ht4�A���f�O���:�A]�;���x�n�'>}v�@:��r�������చR'�]�s�N���jI��m� $��	@R&UM�Sd��Uf�'����L�}�V 4�xI�٦� EP���~_0��$bF�%���`I��9Ȉ�I�0�w�9@�Tf��DcR��;��w�w�рj�{�s��v[u�l��M�����' ��4�?U}���ހ����Dl����@'�Iw3U�in��E�c�u��we9ۂ� ��f��.C���m!��2BB6��8w7��廮�3ٱZ{&f�{�	#r)"*Np����w��t s� �*�| ��DB�&����h�5u~��9ș3B�/�@�(JHA8�$�~�=��R^���� ��5&�n�n˝˼�9�I�0]Ot�n� 3ٲ���
P��P�D��p�9�Ot�n�u8�;�h�=ȇ	������C�&ϝո�kormn�{$�,�t8����4g)�/$�kl�|�{�x ����q�}��@+q|kZ�Dc�M�V�͗���I�0��n���F G"4j)��䊪��r����� ���O���9�T�?����QC���Y`��K�eA�6��0?r9�?4�n����dp��.d�٥��ۣؕHI�I�� ��f�G#����	;f��۠>B�^|ߝ3��U:�v^��n4 S��]W>���f�-�x>�n:����)Z� .�xz����[�`( xI�"qI\�8f�/������?%���Xg�e���
��*P���B��WS���09��ޫF�<��^a""PRNp��)o�}�ʯ���g*��w���6��(�F
�"����  |��!������ ���^�q��t�J�X{6X�`���\�8�Q15r_�6��խ��h87�:..�Q��Oc:ݞ/K{+vɤ�ώӺj"����$��4�w&o8�� �f��i%�$t]��L՘�����p�^�zp��Y�fI��@{���%RF�RD)9�u�s����DDĤ��?n�ﲱk����6�"N+ �f���8{��pk�Vr�=���"qI˼� I��j�y�u�s��������C?�S��}k�a�a]<�^ltg��Qç^ӮK��mn��m�耱Ӥ����"tI�ݤ�]�.�v۶PÄ��U�vw�ً���V���j�i��v-$>6�H������
���	��'��o$���P�z��N8���}����9����D���t�D�/SU�v�j�A���)m�Y�_b����\n�x�e��^ݤ�6j�Oh�̳�߾�wq��}��?��m���vb'�� �v���:���k��3[w<�n�L���/OG֊�ߚ�]78 �N�9̐;ԯ�� ����6GQPRN�?�V	'q;��+�5u=�DC��M�ff�T��H�=�,�̖b]~�� ���`qnS�h�7N1+JI���`j�{�u�s��"$i����fUS��l����j������=^�zto�,�̖}�W�S�T��!B$�z�����r���v��t�nnCtn�Y�n��*�G"_J�H�RD)9�=�uX{6XP{ٓ�Aܙ����Ķ�$K�6�"�o9U�����U>�U�D;Dt2�/ �?~��۬�9ɓ�<��&���$9r\������{7��w]�g�e���ŉ�u"!�Ðj�{ߤ&[u�
:��z��:ֺz�"���T���Y��=�,�̖3ټ��}�ct0z�r*R�(��h�{��7g�k:��oh��4Aiˇp'��q$�)(��Z=�-��d�u,{����e��N&K�TU�3�7w�	7x���@u���w�w�$��8��unK���pk߳�����RC�1#~$(Pb��`.�P���?�UT ���K$��<l�������'�
Np
��7f��͖�&;���Y�V�AA�R7 �S��Z2 ߒ{�)m��s��~~ru۵ũ{t�'=���q�ۅ����&5v�h�e%wm��vW��z�8��(b��˼�V�~I��mףd���76��:P��2B8X�g�rL���`�;�>�`�S���R7'8�n� ��e�W�j^͚X����U�޵#j���r; �S��F�$�`?ED.�d�<#1Frs _Q�]}���U���?=BS����98�f�=��@�� :�����rzT�PTԟ���GPn���R�u��۶�o2��fM��q�����0������K�������z߷@�� :���F�l�s5*9"�I�� ���`����a`s+3y��lϷR����!���`uZ0"""�^�����E��R'�#�ٳK���s�P���f��Vn�"ص:P���躳 �佺S���u'��oU��<��U�@l��!b5VE���uOg]�����ξ݃�N�/@'PKƍ�r���ծ�:x���^-����)�h�ۈ������3է�{7]V��kR��+̤
�b�'���K۩�s����M�����Р�p��m�t齏zGG�lA��Y3ۻN��ێ}�2u�r\�;���T#b'WsQD�;s��Iz�
�"�c������m�-
=;V�k0��z��h C�N��Ǽ�<^��t�v���p�m�n�v�r�ƽ]�vޜVti{��3��W=mǵ[������9�:���7�рoR{�S/��T�cdmSQ	G��=�W���;�4�;�n��I�Dr"8�E:��5EM��5��|�� ߒ{�uRs�w��`mfD�KtE��%1��T�w�}�7OӀw�ـjV��2����Ԓ8I�� �y��+������`s� ߒ{�lz)�7詸8E��wQc#����5�lk������c��;�Z������U!R:TFԄjE�+w����Ł�{����+<QG�?ԊE$޷��]������D�  zD��UP��w�}�p����d�����T�U}�#���pM:p�$#���n���J`�y�Z0N%�As\&쉸�������jV�Os}�y�D�U�51���#��=�y&�r5+F��Ot�9�>u.?%���+l'Igt�n`j�K��Ǒ�v��:q�.�>��6V���¿u7nM�9��0�Ot�9�>�y{R�3!$M�@N	s��]�Hř� ��'��|ݳ"#��2����]�Ԅ�
NpY���Kٷ������a��{��}��}��o}Jh��S�8�I� �نl\5Քr�*�� �����H��"*&�b�jH��c�)�'��@r�d�(��e/x�;7�h�잰�G6N��Q[rJI��%�̚"�@��He�eF�.�<L(�\������nq��(� +20��sL�H�ʙ��9D�p�N�6�5aTÖBR!��8�xz��ק0Вl{|b��-&���p�4�k�}ݪ�-޲#�fе&�����@�7�zs�g����^�U'�e�0
& ���#
B�(a��	Ȱ�V�&aU�:5S h�1A�[2N	��1�B@�Mq�n����ɀ�0�ac H������*:<��
�*>�s�� { U-���J ��������ĕ	����~�X�ټ���(�QRr<�=O���0��ۡ�t߫ 낌�߂��H��Rr�wf��U}��<��� ���`$�\�&*�5��{f��7G:r��m�$����oE����ۇW�d���@"��'�fo8,�v�O#�!�v��މ��\&쉸������;$���F�Z� ߺ��� ���W���l��a@cq�'5�# ԭ@o�^��:�S� h�9��i���ISn�wv=V{��p_{��_��}���%�r��Yh((�h����H���� С >��B�d�٢�G�IoYeDӆ�6	9����I�+V�sv�fL.$s�Z����Tƪ&F�Z��	�y�q�H<�n�Wn��9��N�m�ۙ5�A�9�NI$�III�ՙ���n�fL,�ټ������!e���[�Ü���0��{�7I�
 P���A��H�RB��$��ϦI���4�`u��.Ċ`�N	"p��U_/{7�������y��'����D�j���R"NNpY���v���d���}��	?��LP�x��~%!�B�2Mp�\W"��H\=e��.�]l6�d�Ҽ:�F���[U��5�wg'$��mیi�Xaݹ��[!(bk�&�kX��D�[��/;����u���/�����gs3���l=��wgF㩎���W>�v�@�l�_M�(�h��zW�q��l�\gl�T㭃���`-�&�����h����14n�΍������U��6�n�i�������/靳�%�����pu�Y�.:5�lu��s���h����9�u��C��g�E:R�������V3&D��g�� ��=v�z�7�i�c�O��� ������ٽ��u���Ձ�4�1d ��@Nk��� ř����_W�Y��Ձ�n�,g�`�%N��I����JN���F�Z0*~����$`)KTU(��9�}�*��d���}���3]���YC�*)S�}��㣳3Q����'�b���9ۮݢ�X��O^��:'�I$�Rr�wf�@w��\��5���Ձ��B��:p �I���U�~{�]�舏���)�Ȉ���ɍ̬W���jV��?/z'Ʉ����H���in�v}�ue��Ʌ������jA_�}�8�(�h�����jV�~�{�)I� u���4�SJ_6�wf�;��pY���6�Z{*cB%2�j%֮{>���0p������Xb�r۝��w�?mq�I!)t2	8T������]��f�Y�W_��u�bU$nI�� ���~H�ͺ�7��� �w�<`)KTU(��I��f�X]{���Ȇ��j���ƿ];b9�Y�[�~��`( jM�U�vL��h5l�7��Xz��;A��F�ƩӁH�,wټ��8�?V���d`�h�>]����vҎ�My�s�M��x1��2F��W<u��j�q����t�`�%�n0��'8/f��j� ��9�T]L�LH��q���Ձ��X�y�1{5�n���4�1ԧ�n��u[0��{��2�?V��d`v�f`O)&�'
��,�����]��n���;_S�d�A�C�D��3z��6I���~��9��'8\˔���F���ﺞ�70�ϲ���#��g�F�
}˼Y�uWP���ޙ���q�y�봥kT���[��5vр}�S��N� ��@�LR7�(�+�Gw&�{��p^�v}�uč��픩Ԩ(D�u'����������>]�`=�������m���ۮ��n�X�L,1{2o8�_kf�JS%)5u�|���5vр}ާ���w�~?N�]>�B����A����3��V����ėS��l����PY9��'Oh�D���I�ץ�xvk��9�s�F�!�-�nێ�}Lr��v��֓<�%��{S���.jq?�5�o��dVn:z��9mӹv��p���l� 狱�7%����K���x���M�I�[c�ѵ=���.sX��O0���K��Lӝ,0V�I�=�׎&��z*�u ��r���w��wU��9Y�*�B	�i�%\(�g vʹm���O]�H��l�[6GU��w��}�7pm��S��n�w���}��p^�vsv���IQ�)!�8T�}ާ� )�u�|���5vр|��1�J��D�R@Rs�b�k�;��X~�r93�V��?n��)&n��\ڐ"�;��u`s=0�����p^�v����F��Q�IJ9��ܚ`u'���X9���`�r9Ϻ
^�-���v�'Xذc�Ń��v��� v��m��n�Ͷ�#�O][X��cH�����Xɼ�s�͐��f��|̓u�I$�s��Y�;��B�v�����=�}�~p�]����W}���u Z�Zֵ5)��)��ב�|�h�>�S� G[��6�«`�I�J&��&�}��p^�vҵܭ�2��IQ甓T'
��0���@S�� �7��|�h�:�3s���9��gz��*��!Ƿv鵜�ˍp��h�D�+����s��QD��| S�� �7��|�h�>�S�
��@��qԡ6�!�����ZH�0�=�f�g��;�Q�F�Q�IIH88I�l�Nfo����:�� v��C���ϕ�{�zŒw�
i!*�������=�i��>m�`9�Y���n��NP�QT�H�8y���u`w=0�=�f�w�e"��6�o�4�.1G��+u�l!�n���Κ�#m�8�'�(&U�R��Ē��JQ�����X.�0��z��r�� >�K�܉�
�v8I�l��($ww�s��k��X�۫�i%F<��
O�)��=������D�_���u�f ���� ӎ�r��	�UUP@Y��\*������|߷�e���!C�G�W���������P�&ԑG�]�܌��F��=����CC��pm�I�k���p���n�Q���;��v85�5(O��v�[��m��[��U�߮�!���l˙;�S���u�Ȉ�>m�`�đ5�Hn%�'"�Nfo��~M����� �vю#�'��銸+�7
�9� ՟�;��i`w=0�=���p�{�K�y�a�)�*����`.�0���@S�� !.����H6"$7p���gR
�3|��yW������=߷*��7�o��`�EW?�QEE��Q���8+�޹s{� � �	(*$D2Q�iUP$TZUh�
P�A(PJD(@� �(!`�Q� �TD� �hZ�D�
Q��F�ZUF�ZR�A�bT��B�V��Z�XPiJ
Q���@hE�T)Q
��LR�P�@P� �MPH�CJ�@!2�(D���Ѕ%
�)@-!���3{4�	hT�X��P"JQ)U�DI��
E�NF@ nT� %� �JP�F�hQhZ�F��V%iQZ ��
DJD
H  ��Df E(E(T�(R��%i���Q�DhB JT (EJA�(AL��Q�T�U�HB UD��@)D)R���D��D(@R�:U���p�w��8��B(�4������������D�b�p	�������?����G�DA�����@����A�0A��r�?�����������?�?��w����Q���/����� 
�����O���_���
���U�C�O���A�?�?��⨆�������@�`������o��>�����G��SAJ����
���)(���
�#J�K*$���(J��*$ ��B�(��@�)�B��K*$�)0
D�� �*%*$�*��!$� D!HA(�)J4 Ѕ(RH��L�2(�!J�	% RJ!2�% A!J4%(R̡$���$�(H�� � @$� H�	 �@0�#H�! H��$��$�$!"J
� R�(P�D�J�$�#(H�����BA�F@�D!A�%�@��BIB�)�Be� B� %	�dB�a!	�&B��HBea!	�`�$ HB �BHFA BUXa �!H�!� �d�$`H�Bd	FQ�� `XF��aB�XTP�D�` 	BU�d I��Q�P�H�`	B	F`R�h(PhB�bQ�X$F �eIFUIDD�eFP`) �!FP�aVE �`@`Ya X�eBE�ID%	 !YF�`HXHA��`HAa���a HFQ�d�% �PQ�F X@aQ!X��!	�	F�$ �!�dXB% �	�aQ��QB�	U@�`RB�aFPP�		FHF`B �dH@��i	H@��@�&B	�%R�$%@�e`B��	U�	HFPP!TeDRP$D�	Q�	�	D F��h�I@�BaGz�oO��w��좊�Ҩ��z}]���^��zN�8�s���@_�?�5���� ����s_��(�*���� ?���~�N���
 ��!W�G�'�� _��: Uz�����;��J���
�3\_�z������:Q Uy�������@_�t�I�����o���_�(�*���΢ ��SD?������M�����0���0���<Oמ���8�.(�*�:*<����'�5� P��?���_��~�0PW����TC�Ӿ�����*����?����x����?����e5����P$��� �s2}pS� H  P_l�$ tE  P 	 ( �`�T >  � $P@�!	O�*
*P� *�P    JP
	 �*"�( ()�   `   ��
� }_m��s:����^W�{�< =�=�4q5��tt�h� 0e�`\�� _y�u�xƯ{��>/}�=9�5�����qw���n�q����|Ω� ��    A@�� �<� #@� hQ� ���:h ��� Y� �"  J     A@  @  �@@�% � =i��Y� D�b 
$4  �JP  PU  �*΀&�ʸ��W���ۢ�� {���ͮ[����si^�{�@`���E��yݞ}�_ W�����/@�������-��O.������.c�� �#'��<v����p��x��� ��QB�  
P l Q��_.��>=�y��n�� }zG�f�.6_Z}����ﶯ  �����1� u�7'M���{� �|��_y��3獧���r�<�S� S�n7B�}�O�OW��t� {�(
  
   )��Wz��j�d��q��^�������qe��ǎ����� =9��{����  ����<s����Oq�����;�y��Ҭ �w�q���x��9:rrzN   �芛d�UC#������J����d�b)��R�S��	� ���R�mEH�� Њ���j��@ 4 DHI�JSH�������/�����?�5'{�t{��{����.�������QT�tPEW�Ƞ���"�*�PUO�?��ze0�������p�@����F�i��p#I"��Q����~���\$���BC$GRK"�l`��fs�	��I~��H0����$��)����`�$H�HE$	#Sa�HC�Cf��VA"�`D�G C�����¹$HA#�kO���м�Mo$!IO������:u`�"�b�V!C[���4Ú��[���l�>�Rc+ �+(J�[?aIg�_�.q����kB�� �)?f�ȃ{`�������f�)�@���*�R�%!B$�Jd*E� d!U���`�����H���)�K�J�Z�ӣ�"kg���(�J
�?��1��r��5���aJ�(B�9�h?o�pѾ�HJa
a�IsSf1�f�j7Y�ɴ��L4�Ͳ�4}���B�dX�:s�L�B��\�Յع��|�����D�G��$B-I����}7������8rF	9k$H��DK��904²ț,D��y̎��HSZ
��HtM� h�!��TČ�숤-0�T:&&����&���0Ѱ W&ߞ���@�;�/>�2����� �:)� �>����%M!���M���fE��L��v�l��ԛ1��3.�f�L$����,��yq�D�S���kD6p����1���6�$#Sl��P��l�qd��2�eXK����٬֚)�
���FB什Ĝ֡���6?�>�0%	tco��>1ӱvp�#��;8|;6k�^�K��|lt�$(@�0 `��?e��[41�!�B!rko"�oXzr�k�h��f�F)�D*�QLF�!p����Ms��S>���2�~�kQ��z-++��8��B�;�)��a�9��?~fs	��nb@��sL,5���ILCLX��.��c#�`T�R#HW4�,+.��s\� � �����ᙐ4 [����P$0D�H�q:�I�V�J��e���{'H����L0���?-�>��
@��?g���~�2�]�Vy:d-�=��f��\O�xj�M��-�&��kW\tp�j��zJ�ŕ,���sy�j��L��d01�X��� �kX֬-)JϦ��HJ�����!H[ch��\4�AA���)�$J� ��@����0�����#$�`B�c�Ld��� ����(��B������t��-r6�k�5�BkI8D,h
U!M�x��S5錈������J�&Vx+�&�K�(�[�����\��Ȱ R� #J+�,�"V���Hu�
u4�Ā�I"k�ѿ�p,[ T04�r��b�����o�9�8Hu���,Фd��P����p��@���D��xB����(E�$�#�`SD�$�i$��!aR F�p����dr?!��D�`HW5��@λc��g�����9��g��������Y��� G̈́[ek_h�f��_��!�&�6*j%2;HT�7���r�͙M�'��unn��q�J�)�	�B�1"��5䯯�p�Z�H�TJt�0L����FK��vp�o�V;�4�M �IZ�âLA���'�\������D?���'�d�i�iM����H��C��i?�0��3Fl�@�S��|!YHS��m�ϰ��H��C��'��ġ���>;N	�l!Lӷg �ąS{fR�
b^�껹�\wsL)
B��
�=V!��l�	�5�&i"jI ���R��(�(R�L�B��6#*�kt"��㟧�(]�u���))��.h%ִ��"�$�7z#ϹMnw{;��8˔�![�جĉU��v��Mj�/ ��p�ˏ�,@�0)�� D' ���\u�nmܓm(0��R�8�$ �Mw	�|�*q�Mi5�B��i�~>�;$��B�S��2�
�D� b~6¹ h"���������Ҏ�f���}�B\�~8o�ڻ]&�!�b�"&�BK�K���H����$��6sf�]�k��
��h6��ƠF��.���6�߀�~X�����JA�� �� %�9�G6}Łq�I�
�@�q����!0#5��hB�WJf�Lt�M�g"���`�#ct���B��D8���n�,ta�%1P��@>��ٷA�n�t!q&]�w���,���q�i�+�Ն^�|'ɱ6��k|e0��\4m"A�.����oo�
f��a)�D�A�&O���>H7>浌n1b�IsR�:%�Iq]����X���7 #}��]�v���H�aYBc����±�9���\ՅP�k	���g��M!��ڲ���2���������L�i�K��k_��IY8��	g��Y��rAW��H��1$ Ձ@�	F	X1_�~���H�BZ���G�'	H�H�%ğ>љ��M����E�їZ1
c	���.��)�"V�/�).Ra�D��\���!Q 0)�����"۬��Me�L�q%XX7���w�ڵMƤn]u%3HK����!`P� �u����|p�A�0���s.K�2�	�ԅd�;��0����u��a��K�� A`H$@��5b�qjH���^�j��O(���I�OC��ɿ�GF���Iz�����>�ni4l�0�O���yg��O�����)�vq�!X�G3�ɿ��V#v����X�4�GF͟1h���K�kg�g�6�s\���Ƈas_s�a8��:+�`F	� S5�/.�`MpM
.k_�w���j�.�3��_�o>���J����aP�X��cX��H�R,!$��Xc)؄%l����+�.쐁b��Lb�1���B"˺��np7�$x��!H�	��Z4�T���'�k�3������.&�����6�D�M���P�� ��H\$��&C{~��z�ad�4L4�Ha)��a��1Ԍ��+����5K�ܿH�$d$�uI���щ BC"Dq4sd�u�9�-�gnc�\���V4!X\	��,Ke�5bI12���IK-Z[O��os_�H���	�)��[n�A	�<�x����m�eX��ת�».�� ����أ�GD��)����W@F"�"�c?�"5���1+M}�:�̤ \���q.2�Ʊ�*@���.�h!`�(D�D�%~���	�_ͤB3\�f���?O�JŠŀ�K�����!�������r�^C���Ӵ�\H D�)52G>&c.1U*�/+�{2p��F�_Tu\�d=+sӘ��z�<���*�$������P�n�
h!��p�&�6Ư>�e�4�!u�/s�Ϟ����$�tֿs���#C%�G�ݤ�js�e3x�%3[�&�p�����
�&��c9��
R�V�q�
hJ��?0����%�"�#���"0��B����wJ�)_��P�Wh����}y�����hv�.�
#S$������72�q��A
1+(a����ng���2nq�RZB��4a��2�:�bP�@�wr6��䉭Ċ��¨X�4�ЦH��(@b:�0�I��J㷥q�a>ۜF��^eJ�W��Mg��^Y�>���1"E�)�$�
�
G�-���IO�@�
��lJ$X����	!����d��	 R@`Q�P�ƻ*~RR2�F��G��F���Ŷ�K&��F��.H>�w�w]�
J�����b�`XP$�!J0J���+#.!JT�Ԕ%2=��!����Z��L)	��
1
)'�ހ����$�Ac�A��>޳t$��n�uު|�����K����r]��{����ߎ�#�{�ߗ�	l� 	  �   H   -�  m��      �  tm�$�l 8      $ [F� �   8      ���       [@@       ��� �   UAf�ݧ� P ul:�� r��l�l��gv������s5��@"��ٶ��۶�m&l�T�J�h�J�^ �vĀ �M& � X*��g����UUU�@Gn2��.#m��&ۅ&�ۧ���Ke�m�Uҭ@UJ�%u���!��mR�UR�$��.y�s�6�j�݊ 
 6FU:e��U{d��y��Z�so/2ʴg7f�M�Ht��k�[da��k%$�I���W�C`l��vU\�UZ���$��kq61ҭU +U]m,q��۳<g��Z�^k(�J�8ݸ�l�[���c�y��jؖ��nNdY���m�@t]u�d8����ѻk벽��-�^m�M�k�J��щ2ݫ��9}P�GjyV^s�.j��m���j����N�N��/��U_��)^�Djn��ny�m�nZ{'gv�㚀Z-R�Y����*�U�oy�}�[mu��H������Hk5����]�A�*���B�v�8�2�ma�F������@��D�U*������mun��fצ` �`H� m ѩݍMm�����K��k�r��yJ�`�����O+Z�񕨃��ݻp)vF��Y8N�v�ո)��ʺ$��m���� �- 6�m��  ��5�5Vݵ��  -��Z䝱mù���$� ����m  �n�����8�����\ʼ��������5G�Uٕ �����ڗnYS�%|m�Î��cA��u��l�$����i.��hm�ƹ��9a���$  p�;m�G�-��ݏ�÷m� m�88�� H�k�6�p-����/Y��[C�m�M��ۮ�� b����*��6�89��H� �� H Hlm�� ��"����F���p   �	e lH�b�]6 m���ݲړm��m�NXHH l}[:�K*A�e�C�c�������4,A6iyB���Um�[�em�mH  �m K�ŷm� "� 8ph�  �[A#mی����j�.��=) .6�g�k4��-UU�M��E(j�����vJm��J5Z��k� pm��l ���� �N�[�[6Ԡl�-Y@�^[@V�~����'��k��m�.�ݍk  �H�oM0��!���G�H12 sm����K��Z�h���D �`�-�q�q�7m�,0�l��- t�;k��ZM�v�Q��k:��J�K�}���jI/F�$�!�v�IɌ5Nԯ�K��rA�f�1[t�]�[����	�y%��������$��-��8Hpi$�������'[#GH�ض�6؜9�܇k��ۤ�` 	lt�]5�ۉ  D�G%�	��][��[� i��p۶�!�A�� ���n˯\[v�ZH6���)��� ��uRY�*����m	 6� � �mi�Z� p j��� pH�v٢�-��IBMv�r�N�@�VtVp+�6��X*���j@	n�À6�ֵ�h�I� 8�p֚M�lY!��$����&�r�ʷ6����k��`kX	#]�M�/F�� mH���L��u�u$��ٮ�q�S3�;TUW[����li/����Y/��M�s�Eז�2�Cup�
�
��UU ���ݶΠI���j�춗l8�s���T�L�9�9k�9JZ�Zm�.sVy�'k��鶸"˳lvW#ʚ.���շTS���-Z��.ʘ1�3[7b�C�B��N�`�Y�F� ��$ �vp � ��I���xz?6J�Z���v�W��a�fm���� �   y׽}���M$���ݶp�*��    ��m�l�m��AyV�*�SV�9�knm�m ����t!�V�O��Ci$C �l }m�r@� 	 ��\]6�$�\  6�6d��IR[C�I�z�{�h��Hhm�  w[&�NͰv��z� ��ͯ`  .���n�n��$6�i�i0M����K. ��{�YSo&�8���h6ʬg�ګ�����X�pqJ-�a��(J��P �Umt��l�@h�m$� I����[�����ƗK����  �l�������qJ��P*�UU@R�ޠ����  Un��ݪ]���&]�`�:�m&��6�a! �m�� � ��H�YC��֮�v��E6�.��[E�k�I@��ډ�P����\ {{��  ���l������c���]�  �Y0ʝv��m���횤ے[[l   �ʲ�E��.�UUP z�c�G#����Hr�,�Dغw9�΄3<��˽ln�Ƽ���b�B&q�.�M�-�k<��(q�+�vN�ؠx�U����m�sp*Լg)���gl9$��E��h-6q��km��       -��ge����v�I:G-� �t���aa�,�  [E��ѶĢve��ř��Q h[�J���j�
��ʵp ��@     �m& �E�[@9m��m� �s��m��h6�` 	�7m��$ 
S��m�&�KsI��8R�u� 7m���6� ������-�5u��   ��    �n���m4P  �[p�hkm��`$8� �֋h:�I0m����y�8|  �l�  �    ��$q �`-�$�km��5n�� C��J�  �l�mm��u�Y�	��e m�m�f�z鰐   6�  p��   m� [v�km�۰     ��)   ��  @$  k��  M�$  mk��v�m9�{޶�    d�hm[@6�  m�n��Z�m�['S��-�H     �� &t�6�  ��8 �����  2-�m�� ���EV�7iW �smڝD�-��lI"BN[��:@
�T=��!lё`{j�� N۷n�Rx%�v�o�\sd��'j7=��nD���W` �f�Lק6�c헫�piR\"��d��nt.E�>�v�	Vյ*�/*�ղms�-�m����6�  6ٵ���m� �e���d    	 ��f� ,�@[N�k6�����  rN�� ����P�ĺ\ 6� 84�cJ�+5J�O<�Uuki�m-�m�   m�` �   l���Ĳ���ՠm�� 8��[t�V� �` H-���z�i�]u,�P�m�jX�W*�@PUU* �`-6   y�����8��f���h���-�m�iY���@i����kl� �6mt�[N�]6�i�Z��m -��rE�B�p���햘06��� �|(��RY@e,�6�mUUT-�-�Lp���@$��e�5V�U�R�+���~Ѿ��h)^�F3f:��@/KT��5�vm��L�� $.[$-3m�'����sv�ٺ�[�� v��Yv�� Ӧ���WnZ�
�*�Ԁ�-n*L�V����P;'i�Uq�e�v`��FԤ��:l��Y�m&�R�At��ƽmm��mp'k�m��� � �jM ;����%����8�f���� ���l *����2��[+��J�P�  � �m��[�s��M�]�6̀p$v��Z� �jݱ����^�I*�6*�
��rB�2� ��$�褉e�t� ���Z��6���h�!:m�Ni68	�h�$[Amْ��*E��͛�:�,Αͤ�\�t� X` u��h[@���n�i1m  /6�m�� �m��tͺ��5M������s����H6��Ym�]�U*Җə�����FKH;W*�O5^Ӣz�ԡ]����ӡCp�̫ܴ�V޴jK-�����n���`�h��i�( l����Xlk��<   -��!���� ޻jV����H l $h�4�__x��p �` �`m 6ش���L6� "��pa�6�v�8�^��͢�   �lYi\6� 6�l �2���a��p��#RU;v�j�U��"� �FU�5����mΜI� ���i�`6�n,0  �h   5�K��6�N��]�-�T�4�5Rʺ)V���ְ�nhhi69m��6�޲���!:t��&��ES�6#�?����6�8E1s��
��j#�� )����>D�b�E�~qS���FȀU�qD���\@�P7�~7�?|�ȏQ��M8~�@ڪ�B)�|*���X���L`? i4�"3��`f|)�"(� 0�*��^
�Qz~W�>x<P�t@j��4�|q/����}�b/À'R�b�z���PN��2�@(�(hT"��
����@
Ǌ��1�4�Px�O��(T!@���@�����"?E?5�?����AUW>�uv��������4B1N��|�?��l
�p4+���O��:�^h�?�S���U����]��!���kAD��D�@C�i�%^��1Mg���(�Ӏ�M ��6EC� (�'��А�0vg��C!���$ ��
`�*��~:��DV"#)A@M�!���=U4���@���<���H�!�����������غ��־(�ņ�?DF
kk�?���G���q*�DA�Q( PX�D�R���DK4X4P+�1#Q`B ����O�p��l6Z6�m ph��������:m� �-�l%������69j@�P��V�:%jC��Ď9�h�yqp��-�D��ս�<�b RNen�N�X������\�";u�2���+��K�5v9���rB0��h���m���.L��'���8Է0QjR�eS-c��̭y��Ύ��Vv�V���V�x;+F9{tv0Q;0,F��/LV�����/I�ζV	��ompuA�������U�o`E���m�6ݣj�1ACO����+���(�$=*�@� aN��ۗ�{�mȐ�X=�*�ܷr��d!:����:c�0�Y�������>� ������E��I��[v���F)�݊ql֐t A��@7lne�vJ;rW P�j����t�K�v�D�%f`�v����������#[���z{��`5;S�Ga����c3��<U�a��ڲ���g8wn\S ��Q�;/A�#%[=���j��= v%#�����.خ�ݼ�;<��gXe^���	��ۣ��5d�:z��{v:Ÿ��vd��ĳۆ�#���U.��m������@�N}��$0�dlt�f-Cmo)�h5�3��@J�qIT��l�m�,��˵UNu��A�4h�Z��s8�T�9�����&���u�*�@-��Up8h�kz`��K�[v� �U��Z��:�G/3���Lci;\�9]ne�Ѯ�9K�j��#��Zs�ؗ*N	ra�UU����.��(p��VZڤ{+ú7,m@Ӈ����iLl��3�Q��`�"��
(�K��v���ʚ��*\��2�7Ah�[�n�N�X�I�E�[�KJ��+�ŷn	�fv���m������l9�[Ƃ��^֠��r.��v]���(-�t�q�';;���SRp�GG�Ż4m/
�m܋�mmh�U�-��ˣ$Ѻ�$�*�n8v#7P,�WXU�e{k3Y��&�$�E_����:����b��"1��6�sH�
��6(���a���AC��:[.i�r���c'a۲�:#��M>������H���[>�Unr#�Jr�
�%ӓO)�xe����\a0:W�rGD.��6�w��>³�}���b��	�d4�.p��]���s�WIƠ�c�H�X�֕�p�q����=������v����>�T�����u���v�nR:U�❤xځ���Etth���땫�f7������6���"dx�D�o��q�/<G�W�`�;l�992s�T����IC���޾ �;��^����i���C	��/�)�\ÉqHmmj,}͖fe���W��o�Ć,rC@�ˆ�W�^�7��j���i`ugq�t4���I&���Xm��5������n5"�c��hn=�w4oVfV"���2X�q�o]
�W`Z�u�^�'�A�H&Nv.��M�-���W�F��Y��(��ΰ;Mߛo���~�6� ��� m�XhSEP:˺�5V`�hˎK��*V Q��§����}� ���=2�c��fo郄N)!�r�נ[n�&��ZX�ZX�
H�A�8�r�J�fe�������������2X\|~i�\m��L��{zS@��`:�`�� z5(&��*�)z�ۗoTE��(#�[;��{<V�|�ε�#�v����do�DB�$4l����^�m����4��7�!�LRH�����`n�ڰ>��fV+h(�&�1���z��hO��]���Pj� �B'�`�Az]{g r����ۛ�&�(��=�)�^v��������X�Ma&&�^v���������4
�P¤��� �eΓ>)�n^��R6[�m5���xcO��ӎ ��̟�9$�@��@�n���M�hs�cM����T�,�e����V���v_��K˓)�1*�#d	��Ē/k
��y���=\�l���������mz�Z�#�"�	!5$��j�ĕ�~�r��ow�9�n�H=M8"`]�+E�7�w���5�m�{�̙�[,�i6���Ē��kRI^���Ē/N�n�ok����?t9���4\�>׈�k$N��G7"��t�X����D�'n�f���'j4�Wn)�..Q2�� ?���~��fv��m���Ǽ��F�̭��m��oȐR%��L#��$^���J��y�IWҵ�$�[�y�������概0�p��J��y�IWҵ�l�sw������ҭ��`*�$��R�m�"�ė߿?�ߚԒV����$^���K�-^x�^ِƚ+i<��72��o���r�|*�w~����׽y�m�~�r��m DC���CJ�-�A�Tsj��� h �&"`� ��R��(H�E�nM1S������8 I�˩2Bc�z�<�.#0
�&�%;�.���q�M�b�r�bѸ���us�(V
W�SX�ݶ��m�6e^˪w:ø�F��bJ��ɹwF�Ў�a��a����I�����l�M���Ylv��U���.$ܫiX)ZE��7��v�A��7�;�=�<vZݶ���\b�[I�l���}�w-�m�^��[V���Z��23��m��.ۋc�]�ƭ�8P��c���:���y6Gg��$Iٮ���F7!���I}>&���e��J���I%���y�Iz�L�#��b����K���<Y���m|���I%�_��<I"��ԒWޭ�<�$(��I��%_J֤����<�$�ғRIw���%[�R8�أ��kRFg��ED�A�O��9�m��MI%��W�$�}+Z�I_n'Q �K�)���x�E�I�$��j�Ē��r��o�����w�.�����s'J�����]{<�+��eޭ���� �b��v���=�fv�-����_����7����m����j\����ו���hd��CLj(��E�%_J��~���~�z@�9m�����k�7m����<I/]!�<U��O ��Ƶ$�����%WJ=HB�e��J���I7�b����GUP�J_�6�.s�l��z�J����%_J֤����<�$�V�i��ő��Y$�Ԓ]�y�I}�>��߉$�����%WJ=I%�n �C�8���t훜q��&�L�Z9r:�q�6Q�c�Aq1r//Q������IWҵ�$��|�<I*�Q�I.�Z��$�����$6(�4'Ԓ^޾g����H�f�v�o;[�����3$��o=���D�K�)���x�V���$�}����|w1!� �g��k컶�����Ē���<y��A�(�ũ$��j�Ē��֤����<�$�wqjI/(d����c�Q�"�Ē��ޤ����<�$�wqjI.�Z��$���U��m�k��M�����exu']!��n��8L9u���EWX�e���|�<I+]�Z�K���<I*�jI+���M�\��bng�$���-���#y���6�ɻ%���;�����rH��S4�1df&�LZ�J����%[��I%���y�IZ��Ԓ^S�C^D	���$��Ē��ޤ����<�$��컶��X����&�!>���/<I/]�Ĥ�b�cBq�I%���y�I}���1x�J����%[��I#�������~-�#썼�(�M�Rn��h����6�p0�\�g3+�Β��U273�J�w���e��J�kz�K�����%�`��a1�)�[}���@�@P"kZ��׳7m���y�x�V���$���5c�~_�HE�/<I*ݭ�I/om<�$�wqjI.�Z��$��'�ƛm�RD�z�K����Ē��ũ$��j�Ē��ޤ��nnbo�)# ���<I+]�Z�KΖ�<I*ݭ�I/{���$�?e��2�5�ۗ9��MՕ�������ۧ�iʋҹҷH�tT�CL{v�b� �����@f����p��q�On�cS�����8�,v݇m;�۬�9�v��]�N�h�F��^vP�e8���3�'�gh����vDۋ�9ۙ"m%���$@]�m���>����]dkAq[�&˺؍�=Y��v����۫Z�+��M���}�۞6�6�	{s����y?����[�2Cε��5Qt�l��;XX0�x�qӹMڮ?�������$�v��$��g�$���-I%�:��� X�@m���%[��I%�u�<�$��G�$��j�Ē�¤�Mb�cCq�I%�u�<�$��G����Ͼ^x�_;>kRI.��n�4�1��drx�Ut�Ԓ^t�y�IWҵ�+����y�I{��<�L �	�S7m�����r�|*�;�L����s�%_J֤��N�^�1�<"hi��.�ڹJ0j�Cv-ϡ^�8��p�c،���N�q��I$��J��z�K���y�m�k-����F�۷��ͷץ�M��jJ����[oT���/ߧ5!! MXĄT�!F�@i]��"g��,�Q�$��j�Ē�����nnbm
�䌃s<�$�K�Ԓ^t�y�IUҏRI^���Ē�ҽ�a�&1�c�#RI^��<I*�Q�I+���x�W��jI+yV�<�0s؜^x�Ut�Ԓ^�-�<�$�K�ԒW���-�� �z{9�[5�IXMi52��S�Y㋘ŧ��<���j�x�#����r�:�@Ƣ���$��}�y�I^�Q�$�KW�$�](�$��n&� �fI2�D�h�-����ٿ
*�e����[n��%��M�ߗ�ͷ�6�V�
r�U8�m���~m�;XU��5ĸ�槠-+�`��4C[I(�����f!V�KS�X�T��A�`EZ�I��Hb#b�������'���{1��؎�P�P~���ϔ5�\�������*?'�p�8���F��HZ��c	�HIEx�������8����^�vF�:�[��	�S�Ԕ�d#v�s��?ZЍH@���� ��bPW�B�@�Mt4|�`���πJ�@*�l.�g�9T� 'U�SZ�\���9R]e�jI+J�V:�����E牶,�a`gs-X�w��$�ܭ�`w|A���i��ƣQ�@�n�ﯜ����p}l�>J(Jv>S.�/�=�g�z<M���6�wX�:;nV���ה��́��bm
���x���@��Z��4��h.9��6�AH�*S�3�1ޤ�>�֖���_U�|���/�͈�bqh�_� ��X�s��78�c����1$�7
��s@�_U�^���JA��[U�"�N�������h$�v&� �fI�93@�����j��������X��{�-"��X������G&�C(m�u��7Oc�\n��,��J�vѭ��Y(���Z��4��h��J��V,_�HE$�-�Қ�w4��Z�j߿$w}4�M�n5�Y�|���\� }M��v���V�B)��9����@��Z��0���=:u:��*�R*�N����`j�r������;3]���^�8a���ۯ��(f][��3E��c�;Da^�i��c�ؒ�l���L�<��PG��]�v�q]�A�=V�zݹ����	2�،�q�#�i|?���y����۪,������Kː��=���cp]�A+:2ێՊݞl`v�K��c7�<�e�Q�Aس��is*6�wr�=�I51��h�L�E�Mrr�̧9��k�j��Duq7*����]�$7����֤5�MkF�� �]���ߛ�۟���9��ݳ� r[�rA�a�l �6'�u�|h���=��Z�j�/�'&6�BI�n�w4}}V�yڴ=�����w$M�I��h����i�����[>48��Q'H��hs�i�^���@�gƁﯪ�<�XA�,a!�H�=��������~Z��ZG#�V�"���8���[�rR3u��+�69��`�Ƴ�q�������lX�4��F���u��@����ݙ��s���;��|���:���Q5v`��rX�¸��P��~��������/�����g�*@MR��R�; ���`~�+=�%�������.~a���`}��LR$�<��hl��ﯪ����aRr0��I<m�@�e4}}V�u�h^��<��
V��Ǒ`]�9��g����nPM���k���&q�f�+���Ѥ�lNd���#R�h����@��)�u���Z	ᨁ�jE�m���4�S@�_U�yJ������H&��<�)�~�uٹh�E!�ާªb�Ǔ��h�l�=�L�pX�j8�4�S@�_U�m�ߗw��w�q�z��Hc�E���1�Is�}�W�fz�X̬,s�5=nNC�yxs�m��=��Ⱥ�;�[;%v�xz�s��%�2P����q՗.q�bj�$b�)�������,�V�?0�f�5w5���(	UV�ea~^\\R�W�2{��;��z�9�$ٽ�5�T�rJcnBJ,ݭ,����\�9�&�߾�w��@/.b�$m�G!���q$�{[��3wj���,;ĸ��n#
 ���?L& ~1�!��@��\�?~��wӾ��j D��h[f�����~<����=�ڴ�S�<�~Q�"%�;��v�K���q�z�ҙ�)���;����sY5�@�$�xs��u�M�]�@:�����;�HGT��k�^JC2{��7��>�f;�&Ϻ��G�鲩69TX��v��U���f�3r��??��8�1,��ю8�>į��w?�Z^����̿y���2�L%�%U���1��^��x���; �w*��q����nL�40���Z��՝�ue�G�y�m��\a�Z)�v�lV��V�OQ�&��xٗ��c��y�D]Q�U½P����)�c�@��\�!�/a�m��꺹��ݻn��=��e�
�1�]!n��v� ^,���U ql]26׉9�$��M�N�;�c/9�+�L�];�<iM�G>��'Nzv����p�n���*�Oww�}�������⭺��W��m��.��x�=��X�n�b��vy�<�PI����|-?͓M���w���=�ڴ����s��Z�_d�����@������9�/r>qq(���Vr{���d����xj D��h[f���,�y�ZX��v�1�x�TT�H�4=v����=��ZbWﾚ}Q��
�$j8hm� �w[�| ����=�ـyo!KU�l�k�޶���n$u���c�7\���8.��.ͭl�4$�����x����q\�h���� ����l�9�f�]�+���R��R�; �fU����I��֊#.]ih!�<��{^���������w�lޛ�F��4������i`w2�����2o��o��3��ME�qQa�y�zX��v�̫s���_��۬�R�RDG28�p�=��Z������zW�;������X��tH')�ڝ��鮽�T�yn`�ztN79�%�o/m�����E����E�?�y=��_�����~7kOs��}ٚ��֩�r��©S�䪰�w*��8��Kˊ��z�Xd��m���H�Q��"�y	1�5�'}�znIϳ�n� ��z@ D��O{�`f���S��E�ʌ�M�Uğݬ�`��`��U��<�ߍՖ��4�d�6�G�u�h���m~7kK�Ӹ���	�	��guq��d1	n�&.%�r�R�8�(���[9�����mBwѱ�H˲������ـ{i��G���^ ���4��BBrhl���=��7v�ﻕ{�6�٩�S��*J��ϻ��;��g����U���x�?t�_)S�*�nT����wj�;�ڰ;�XX>5\�i$$��C)���Z5�B45�MiB2M �?y��}�@�Մ��<a!�7&�{�Y`jY�z~���`�ʰ?|N�*F��b��GnX�)m�Fڷ\d���N�PvmkxS��������֋Z�*�����������^\�_@37�`f)�y�y8�U)UE�����3of�w_����oؑ�3�bLc��Jv��V���Y�$��7ޯW���/�kb͈!����4>^��vn֖�q�{�o7v��ֹUU��B�i�9N��ea`oٗ���{[�s�~�ܐI�b�:��H��g�lF$A6��t�C�|~���'�HM�P���H��E�!��$b$B �(��B�(B�R$f�;���y��1����f^t�<�j,# ����@`���$d��R	�Bp]B0LB�A>>g�%e٣X���0 BH!��2)#P�D�#0#��1�D�{��7����f�7�����.�B��2�,I-�S	q	"����!� ���!1!�H��~ �O��˿��gn�Q?,X�4$��]���®$�4������ݍ������ �*�i��	�G�mf��`�6� ���Zl��������ܦ�њ��	�Q�p(��xĶ,�:�Ëg������7l�ۅйD�T�j@Ql1�A�kk���vXu6hj�\�q�8�㙋�()���p��%M
I����]t;�U�E�h�m$��70;�d9���t��s��c�[�F�<�=�\=5�M\�S��SZ�v:ˌ�+���b�!��T�(�:j�]����ick:��۲=RL�0n��RX1
��z��Pc��p�T�P�z�V� 1�1���Y�r�|�'�7}�}��^�u�$�v�\FV{ܻ�<����p��<� �즴�+�4��8	F՝��A���[���X����YG����]�ɕP�:�3]��l6_��7��vʓ`����=�ϡ@6^ny�qƧ�6�;:��[��ha8i�l���p�Gkh�}�v� 5�YY�\�r9^(����ع�s����$��U-��a�������L����\նқjڨ{��s�&Zq����^��^�j:�l�XF�jr��KB+R�Fz7Ѕ��ё�����D<Q&ݰ �U0<��Y��4v�i�St�f��e���6��k���
�w� �0����ξ�Tɑ��i��!'m��i ��v�/H-��Xh�t�z�8�v��m������j�]�U�A\�vnw&ѰԫԄ��s�b�vr�:�v�m�91�s��!lp�)y�nh�n�Jζ@j��6 ������	u�Si4���	V_VL�p�7i��b]�1�+��N�m�<b�C�;쪭�Ql����:p'c�hy�e.��W��Ψ��獷Y;$��nN�vNv�,�X�@�5.�&��iU���n�.�Ez坵�K�(��;Wig�7(�]��\L6*ܣ`��A��oUD�n�-�4��1�iJu��Z��+�@��/���<m$沠m+ʓ��h�alC���L;[�ڪ��#��։�oY��5�٩�^���|i��	 x�!�#�$? S�'蟕��m:���s�ww�[9w����g����s��NSh!�دH�^;9m�)5+���zl���]$����0u�0�WZ6�э����R��7N0�`C��i�ۍ�C�\���i�1u*���n�aȲ��ְn#�Li�gOCv
yU�D�B��p��쉻8�oZ3׳a�f����e*ڸ臍�l�T��c����9�οg��Q\�um�I:���{w�����~�V��V<�J=�M۶������q�4	��c�-���9�9����7��gƀu�hs��S@��7�Ȝ�"q8hs2��&ϲf�7kK?�g8�̽/����&q3�{�5��*�nG%U�"X�%��u�]�"X�%��{~�ND��T@�Dȟ���M�"X�%�}������$~��,K����a�5un�̷Z�ND�,K�����ND�,K��~�ND�,K������bX6'��}v��bX�'�ƛ=f.\�Z.�ֵ6��bX�'���6��bX�-��m9ı,O����9ı,N����r%�bX��?N�~�v���r��혠�v$���맂�`�j5�� ,絅���;�1�9L�o�r%�bX������Kı>���Kı;�o�a���&D�,O����ӑ,K��{��)�Y)r˫3$�k[ND�,K�뾻NC�@M"���IU���P�ȟD�=�o�iȖ%�b{�ߦӑ,KĽ����" �2&D�;���Y�֜sSV��.j�9ı,Oo�m9ı,O���m9�Ľ����"X�%��u�]�"X�%�OǼj�VL�Y�ˬ��r%�`��{�M�"X�%�{�{[ND�,K�뾻ND�,�`�D���?�ӑ,K�����3	8������f�ӑ,KĽ����"X�%�'��}v��bX�'}��m9ı,O���m9�q���~����~�J�{\&G���z��n�5�n���°qF�;v�[�=�Y�����f�L)5��s.f���Kı>���Kı;�o�iȖ%�b}���a��dKľ����ӑ,K�-�e�!���qQU�w���g�ｿM� �X�%��{�M�"X�%�{�{[ND�,K�뾻ND�H
dL�bw��o��ra��L�M�"X�%������r%�bX������K��0 �cQq dL���߮ӑ,K�ｿM�"X�%��~���n��ѓ2̷5��K��F(�=�����"X�%������r%�bX�����K��A[����gq}�5�]0i�:d�*���9��t��H�b�ouٴ�Kı>�}ͧ"X�%�{�{[ND�L�g�X�Ì�@8&��Q	*�J&����1G�c�:�]�\���C��-�����j�7F���\��r%�bX�����Kı;�{�ND�,K������bX�'���m9�*dK����R浫&e�u��]f�ӑ,K�����6��X�%�{�{[ND�,K������bX�'}��m9�,K�w�\,�W4f�u3Z�r%�bX������Kı/��kiȖ-�bw�ߦӑ,K��}�m9ı,O~�&��P�@U�G%U�~8���P��z����ı,Oo�m9ı,Ow��ӑ,K���")�D����".�T�1 ł�%E����j���Vk���'$O����/�8���,�2��Dt�TTD�kiȖ%�bw�ߦӑ,K������]��,Kľ����ӑ,K��w�ͧ"X�%�~���f�hՄz]�T�X�0���	�����哝���9ڦ��2۲f̶e�[&�SiȖ%�b{;�fӑ,KĽ����"X�%��｛ND�,K���6��bX�'��ܞ��!tI�d��fӑ,KĽ�}�� ؖ%��｛ND�,K���6��bX�'���m9ı,Oߏz�9�%.Yufd���ӑ,K��w�ͧ"X�%��w~�ND�,K��{6��bX�%��m9ı,N�]=���G4h�ܖ�iȖ%�bw�ߦӑ,K��w�ͧ"X�%�{��[ND�,K�k��ND�,K�������Z���I�����7������ͧ"X�%��������%�bX������Kı;���iȖ%�bA4��N��2���5%Ԑ!��tAS�m��OJ�O$��Wn�\���C�pK�ظ�a:��͜v5bxە�5��T���/��[��%J�������Z�u��ֳ��w�l�Œ'���k��An��n̶q�uL
zP�7�0�l������;6���i��/h�fx65��\��b�����zǩ�	9S���m�vnd��b�\ʦ��8��$󥥮߾�w�x�rv�,�W`�bg���=\EW33�\�Xul��s�ܝm�[0�.G�z�nh���w�{��7�������ӑ,K����ӑ,K�﻿M��n�&�X�'���ͧ"X�q3�ۭ<�R *�j��U|_�&q8�'��}v���ș�����6��bX�'���ͧ"X�%�{��[ND7���{�M�^߬fZ�3���x�,K���6��bX�'s�}�ND�,K�w�ͧ"X�%��{�ͧ"X�%����I�2ٗ5n�����Kı;����r%�bX����m9ı,O���m9İlO���6��bX�'����-�B�2ɫ�ͧ"X�%��;�fӑ,K��_����m?D�,K�����r%�bX����m9ı,O�K�$���.��:��շ9�Ň�5����>;l}�Z譞�;l�r[��+�=F�	��?�����oq���������Kı?w���r%�bX����m9ı,O��{6��bX�'{���k4�5m.k35�ND�,K�}�M�!���Uq�Mı;��iȖ%�bw?{ٴ�Kı>�wٴ�O��{��{��7������t�)qL�m�"X�%��￳iȖ%�b~��ٴ�Kı>�wٴ�Kı?w���r%�bX��|K��4k0њ��sY��K��2%��ٴ�Kı>����Kı?w���r%�`O����|_�&q3��^�4\=MI�U*kF�5v��bX�'��}v��bX�'߽�M�"X�%����fӑ,K�w������&q3�6�a�T�R6F��'��M�n#Ơ��ת�d5�G2=��ts�zcP��{�7���{��~��6��bX�'s�}�ND�,K��w�iȖ%�b}�w�iȖ%�bt�z�$�n[��-����Kı/߽�m9�D#�2%�����iȖ%�bw����r%�bX�~��6���&q3�����<&�&��Q*���X�%�����iȖ%�b~����9�bj
Hr5��6�&D�����Kı/������bX�'��}fՒ�auff��ӑ,K�?~�}v��bX�'߽�M�"X�%��~��iȖ%��*�
�D�}���Kı?���YsT�a��sW3WiȖ%�b}����r%�bX!�~��iȖ%�b}����r%�bX��k��ND���/$��,����Ъ�(��dQԞ:玟X�+I��r��s�V�âd�Y��ŉd�5D�Tڛ�.���B����$.���d.D�,K�뾻ND�,K��w�b�%�bX�w���r%�bX��|K��4j��5�K�ͧ"X�%��u�]� �%�b~����9ı,O���m9ı,O����NA,K���Rl�k�ѪkW3WiȖ%�b~����9ı,O���m9�,K���fӑ,K����ӑ,K�������kP��{�7�����wn�'�{��iȖ%�b~��fӑ,K����ӑ,K�"����(�~��o�k6��bX�'LgorL�幫rۚ�ND�,K�~�iȖ%�b}�w�iȖ%�bw���fӑ,K���ߦӑ,K��;��Y/�}�s��y�;�\g�E�B�C[e�;=�[��=89��p��f���'ۂۂ7	�������%�b~���v��bX�'k��m9ı,O���lD�,K�~�iȖ%�b~�{���Y)fVfYu���Kı;�]��i��bX�w���r%�bX���}�ND�,K�뾻NE�,K�׏\��c�h����ֳiȖ%�b}���iȖ%�b~���m9��"~���v��bX�'��k6��bX�'���.�V�̺.��fk56��bX�'���fӑ,K����ӑ,K���w�ͧ"X�%��{�M�"X�%������N5Lњ�&f�iȖ%�b}�w�iȖ%�bw�w�]�"X�%��{�M�"X�%��?wٴ�Kı8��80~�Ÿ��|����v2/R�#��옮U���u��nWA2���׃"�h��`,�rܗH;�pu99A�e�C�ZA�Mc+;������� c'��%�ڽk�q���|���XՎ�&l� �Żu	F�ss�n�^Q��Ⱥ{ctG9:���xD#�g����}�nb��=���/����{ñF��\��8,�\���ִYu������5�|B���&�"��ks�Z�n�ts�n[�F��Yy7W)�v,1�'��������3㫵�X����ı,Ow����r%�bX�w���r%�bX���}�^D�,K�뾻Noq������������K+���}�,K���ߦӐlK����iȖ%�b}�w�iȖ%�b~���WiȖ%�bx��d��-�u�2ۚ�ND�,K�w�ͧ"X�%��u�]�"X6%���w�]�"X�%��{�M�"X�%�������an�.Xk5��r%�bX�w]��r%�bX��w~��r%�bX�w���r%�`��2'u�fӑ,K��O��p�[)fVfYsWiȖ%�b~���WiȖ%�b��w��Kı/����r%�bX�w^��r%�bX�����'�d4d:�g ��'%v9:<C�\tg�X���+�ے��R�-te�^�6`h��"X�%�{�kiȖ%�b_�ﵴ�Kı>��yı,O߻�j�9ı,O��=fh�Lˢ�h�sZ�ӑ,K����i�b;�!��5�i*):�U���H��ȟD�7��˴�Kı;����ӑ,KĿ��kiȣbX�'�{�fI8h�3FjjK�ͧ"X�%��u�]�"X�%���w�]�"X�1@ș����ӑ,K��{�ٴ�Kı=��y=�L1��MMK���r%�bX����WiȖ%�b^���ӑ,K����iȖ%�6'����ND�,K����߷/~�2�֑Z>�~oq���b^���ӑ,K����6��bX�'����ND�,K�{�j�9ı,O��!|d'2L3V]jP̸h�NU���77.�N��8����R�����{��n�L���e�ՙ�sZ�r%�bX����m9ı,O��{6��bX�'��~��
�ı/�����"X�%����_�K���决Zͧ"X�%��=�fӑ,K����ڻND�,K������bX�'����NAlK���޹�9l�]Y�LֳiȖ%�b}��ڻND�,K������c ���)�~��ٕ4+�^��Gx&D���h��
�Bl9��s`|�	�j��
����ϙC X�� ���3�}�ځ0M`�5��@��RD�jY"��STр0D"��>�D�d�
(A��cpV@5��p�q�!����}����Pȃ�A����)�'Sz�l����ƳA�KZ��D ?;��p�h��`#���(��>l�A���J���	��(�� z�N"T�D�Oٿ�ͧ"X�%���}�ND�,K��OY��\�D�f��j�9ı,N�^��r%�bX����m9ı,N���r%�bX�w���ӑ,K��g��5Jd�f��]j�9ı,O��{6��bX�����ND�,K��~��r%����=�����Kı>P����RY��c������-^�Fm�s�xn��!�Ϝٖ���G�]�룫�[�{���bY�@Ȟ����m9ı,N���˴�Kı;�{�cȖ%�b~����Kı=��y=�L1��MMK���r%�bX����.ӑ,K�ｿM�"X�%��=�fӑ,K��{����7���{�������{�e���f�9ı,N����r%�bX����m9ı,N���r%�bX����.ӑ,K�����d�L�n�f[sSiȖ%�b~�{ٴ�Kı;�{�iȖ%�bw�w�ND�,��dm��k~�ND�,K�wyBfZ[��j\ֶ��bX�'}�z�9ı,N����iȖ%�bw���ӑ,KĿ��kiȖ%�b{��!)��T�����7fT��u�{k����Қ���'ld�2P����b�+��b2�Q���%�bX��}�6��bX�'}�z�9ı,K�{��r%�bX�����Kı=�t���5�5%�&k5fӑ,K���]�"X�%�{�{[ND�,K�׽v��bX�'}�rͧ"X�%����=fj�ɚ&]]\���r%�bX������Kı;�{�iȖ%�bw��,�r%�bX�����Kı=����N5Mh�MY�m9ı,N�^��r%�bX���s&ӑ,K���]�"X�%�{�{[ND�,K��7�=��4։�����ND�,K���d�r%�bX}�����%�bX������ND�,K�׽v��bX�'�~@&�(f �"�T �D����P-P�5 `�)���w?q��ܛŞ�֑��ƽ�r ��fq�92W����M�+�����=`3J��OX���ۇJ��&��ZL��j�\��.�<��Rc�]1�y�sgg��b�T����ę�9rZ�]ßH�EK'�[Z�Z��1�G@{-�,�ká��vca�r�gx6^Ǆc=ڇ �X�l��W�m�W=y�m(�=QF��\�����O����=��1��N�];����z7^{^ն��w�-ьv�wp\g�='f�X��.��tN��X�%���^��ND�,K��{6��bX�'}�z�9ı,O~���iȖ%�b|g�_�e�,֬�s5v��bX�'���m9��"dK���v��bX�'������Kı;�{�iȖ%�b}�^����Kuar�5��ND�,K�׽v��bX�'������K�AHdL���]�"X�%���]�"X�%����f[��[�]Y�e֮ӑ,K���ߵv��bX�'}�z�9ı,O��{6��bX�'}�z�9�2�D�=�x���rrE@�U:�w���g8�ž�y�r%�bX����m9ı,N�^��r%�bX�w���ӑ,K���{=�2��#��[��{:m��Z�n#&�XN��pc�H\�g3��x�7d&+�]�"X�%��=�fӑ,K���]�"X�%��{�j�9ı,N�^��r%�bX�~���'��f��.k6��bX�'}�z�9
�j ��ƾp6�'"X�߷����Kı=���]�"X�%��=�fӑ,K���k��Mf8kD��˭m9ı,O���WiȖ%�bw���ӑ,K�����iȖ%�bw��6��bX�߽�����i��)M{�7���@ X�����A?_{ٱ$D���I�$��w���ӑ,K���־)��rd�[��j�9ı,O��{6��bX�'}�siȖ%�b}��ڻND�,K�׽v��bX�'��Cn;���쑸v���a����n��R��ٮ7���ނ �LX��jw��C�m\�m>�bX�'������Kı>�w�]�"X�%��k޻ND�,K�{�ͧ"X�%��{}m��e�eՙ�kZ�r%�bX�w���ӑ,K���]�"X�%��=�fӑ,K���m9ı,N�]=r�N�jCֵ��m9ı,N�^��r%�bX����m9�H�" �=5�q,L����Kı;�w�ͧ"X�)�]�ƵUT`�H�:t��~8��ı?g���r%�bX�����Kı>��fӑ,K���]�"X�%���.BpѪkFjkR�iȖ%�bw�ߦӑ,K���ﵛND�,K�׽v��bX�'�k޻ND��7���~��ى{��W�B�\F/<�D�ks��K�ɝ�p�[��{p�X�<��&�&�L����%�bX����Y��Kı;�{�iȖ%�b~����Kı;�o�iȖ%�bx��뙭K��53.����r%�bX�����Kı?{^��r%�bX�����	�L�bX���k6��bX�'읭�'��!(prS�/�8���.�n�ND�,K���6��`%��u�k6��bX�'}�z�9ı,O��ߡ!.���3,�Y���K�䃑=�����Kı?{^��m9ı,N�^��r%�`xC� ~����羻ND�,K�{}���ܲ���5��ND�,K���m9ı,N�^��r%�bX���z�9ı,N����r%�bX��z��l��%�RkS]u��]�>8�h8�s�Xk�їvD}����刺���٩��w���oq�������9ı,O�׽v��bX�'}��l?��DȖ%������iȖ%�bw��N�z���ڴQ���{��7����׽v���G"dK�����ND�,K����fӑ,K���]�" eL�b~��䓆�S4f��nj�9ı,Oo�m9ı,O���Y��Kı;�{�iȖ%�b~����Kı=�����I�M[��j�9İlO���Y��Kı;�{�iȖ%�b~����K��yWQ=�������{��7����������ң֒+Y��Kı;�{�iȖ%�a��o���>�bX�'����v��bX�'��}��r%�bX��T �N, D�Pi�Gd�̥��5.�fL�kH���7*�������:-�ٮnP4�5�q�g���~���V���Y�G'�ʮ�Ŷ�5�s���%t�����q>݋@]�ʽ����Nr݌a����sy#��B�j��j��P<h�Mvܑ��e,cB�6vI+��%�vx��Ȫ��곷H$��9�Ϲ�J��
��$t�'ۋv�켝u�nk[D�8�sV�7��D�a.�I�4j�a���v��^ۅ,��=�c��k�r��;�!��s�o���h�G	C����x�g8�śY�iȖ%�bw�ߦӑ,K���ﵛND�,K�׽v��bX�'��oА�VSV�I���r%�bX�����?�`�"X���k6��bX�'����v��bX�'�k޻N@lK�������e�eՙ0�kSiȖ%�b}�w�ͧ"X�%��k޻ND�,K���]�"X��2'����6��b�ow�����뗋��SO����7�,N����r%�bX���z�9ı,N����r%�`A2'�o��/����&q3�=ZוUF��"QU��ND�,K���]�"X�%��{~�ND�,K���m9ı,N�oK��q3��L�ՙcOi�$UHu(�:����z��շE�V���>Wm��kX�neh�vf�Y�٣T���[��ND�,K���6��bX�'��}��r%�bX����yı,O��{6��bX�'�C^0��e$֤�ɗ56��bX�'��}��r�#6�_��ND�=�o�iȖ%�bw;�fӑ,K�ｿM� %�bX�=�zh�]fe�SYuu�fӑ,K�ｿM�"X�%��=�fӑ,K�ｿM�"X�%��u�k6��bX�'�~��&ze�d�K����r%�b��=�fӑ,K�ｿM�"X�%��u�k6��bX�'}��m9ı,O��ߡ!.�Md3,�Y���Kı;�o�iȖ%�a����?�v�D�,K�����ND�,K���]�"X�<ow����|�����Z�ۮ�\s�]<9;7����Ct�g���n!E���u�c����̘f����Kı>�w�]�"X�%��{~�ND�,K���]�"X�%��{~�ND�,K���5�t\.�0�j�Z�ND�,K���6��X�%��=�fӑ,K�ｿM�"X�%��{�j�9 �,K���x�k!-�$֦���ND�,K�{�ͧ"X�%��{~�ND��S��I�QV�9�=���WiȖ%�bo�z_㉜L�g�w4n��J�����ͧ"X�\����M�"X�%������ӑ,K�ｿM�"X��)2'u����ND�,K����g�d5�jd˚�ND�,K��~��r%�bX�}��m9ı,O��{6��bX�'}��m9ı,N�SԞ�;T]��iֺ�p6l��q��������s��������w���ir���Z�ND�,K�׽v��bX�'����ND�,K���6��bX�'������Kı>����3�.Lչnf�ӑ,K�����i�0 ș������ӑ,K���o�WiȖ%�bw���ӑ,K�������C2ɫ�ͧ"X�%��{~�ND�,K��~��r%��S"dOk���9ı,N����m9ı,O����yl�,��&�jm9ıAlO���WiȖ%�bw���ӑ,K�����iȖ%�����>
D! @�����s`�X���ɴ�K7�������֛�抏�ߛ�d�,N�^��r%�bXD��i�Kı=�����Kı>�w�]�"X�%����n�n��L��є4�5�C��D�v��*hd;!��[��f��OԆ�f����d���֮ӑ,K�����iȖ%�bw�ߦӑ,K���ߵv�Ȗ%�bw���ӑ,K������TѣT���Y���Kı;�o�i�-�bX�w���ӑ,K���]�"X�%�����ӑ?�ʙ�/`��8�`��D$�����&%������ӑ,K���]�"X��b~����Kı;�{�iȖ!���~�������W�����{����E��=�����Kı;�����Kı;�o�iȖ%�b}��ڻND�,K�?C�&ze̔�[���j�9ı,O�׽v��bX�'}�z�9ı,O���WiȖ%�bw���ӑ,K���9�e���4�" @7�B�v�����,b��$H��@�V���!$�������A��i\�cӡ$] <���*qS�@��4���X��P��G�n���D���R��t�&��$	$UHF�P�Sa�P���� h"/�g*�ĀU`EdJ��?.�2��`�^����E7�1� ���L�H! H���N��1T7��> I4u"����v(H"���G���#`� �"�������w&�mֵrl��l �p8-�m��  [B�n�p%q��I�V��=n�@Gت��V�b*Öɫq-��A0]�*Q� �Q���)ݬ�{870�ڷN���%�\e��ۜV���h��YD���"���L,[w�(u/"�SUɪ�YY�w'>�&��v�l�6�I�cL�$�)6�������ҋ8��g/��Իn���4�������]����)�f�pK<�zCK�l�����f�efU�(�Vc�<����n�}g�X^a۷Z{n�m�����S�,�ZV����Ě�`ѭ�
����d�.5v����Ojs�0�2td:�5��F݃���:%���'n�g���7�Li�r;b�X�<p�ی5��^��íqi��.Թ�л[�#t����;e�5�����.lb��i�i�3X؋V�<WUlj;/����;]l�+��<��v,񵴻	���.�vM�����=oi嵭��S�e�l����RIj�=�ݤ�&m%^\��d�NJ�]ـ+L��lA�{pݡ��IfI��/:��$ۥ�8�GFG����V�������!���5.���V���E�y[i��vT����Y9����Wj�%p�H�m7T[vĀDҶM�Xv���Y���yP��8���/�&���I'a2r�­�5fۜ�kJ���q�ZK��Ρf�T;bx�f�n�v�=72\�[��d_B�8zP*�H��KUf��SZ]I�ZD�jG%5UK�Q5�)&�;>eC��Q]TQ�Uw"�I^وG���[��1����gDe�rl3�Kg<��Ƿ#���xx�0����_<g�3&�m��Q����R���J��m�h^oj���.��YGr��nUҜ�3Y�l����+6-�<�Gp#n}����Rq�%��Uƃ�l�>sxv�je[9«��Z��<��9ݴQ�����d`*ٍ�F6[պ.�ֲܤ֋�b������G�!����T���b!���WK�S��O��8~3_/��{����ݸ��vۗV��{9�8+��Ht���v�H�YVf���אt�ƳE�������Y��s�ە��m���)ݺ\v��Oc�رݗ^�f�E�{vf�P'j���;Ô�zs��z%��'`� 5�{mJvI�ۧh{h�\Bcs�#��<�����=5���PMm���wë��)�h����-�I��[ �6�֭�z�eq	y�e���笧n��`y�GI��6�z&��GJ��{}�DIÇ��s6ݷb�l��c��%�b~��z�9ı,O���WiȖ%�bw�����'�2%�bw��;��q3��L���c���ht�C5�M�"X�%��{�j�9ı,N�^��r%�bX���z�9ı,N�^��r'�2&D�=�x��k4�.�0�j�Z�ND�,K�����ND�,K���]�"X�%��k޻ND�,K��~��r%�bX����ƳXB��2j���WiȖ%�b~����?��2%���]�"X�%������ӑ,K���]�"X�%���)��D�����SiȖ%�bw���ӑ,K���ߵv��bX�'}�z�9ı,O���6��bX�'�'�w�C�Ѷx�¨]z���Y�ڨtz#do@ᶲv��wm�F��r3���K�۫���~'�,K���o�WiȖ%�bw���ӑ,K���o�a�"O�dK�o��w���g8����;k�B��jS֮����r%�bX�����:ӡ`c
Ѝh�|���l9����K훮����S�$��]��DرĜn8����uv���b�:�V��SĠ�ch!����ku�fVӰ;�1�y�v��7�4ih���D1�r-��b�g�Ͼ��_�}�ZX�1�gP:xUp�M��gdn�.��خ�t�b:ㆳ��Xx���ˬ˻mJе�M爎��m�����>��2��3&c�������vvc�J�Q2R USuN��2��lݛ���2���k�hb���,�0����!�WM���w8Z������*@�)P�b��;���U�u��w,���U"�I)�k�2����7]��ea`ev��/�c��,qH�r-�k�=�����u����v��P�r#�·�\;[gq<�Re�=u9�y��e�{��[��S���V��l��`a��m���k2f;�{YOW��u�wkD�J4,m �4]�~�����ٺ��+�I6gVi��ƇL�RU;���vd�vj��8��z�X�����ά�R�J���D�uT�=�$�ku�ݭ,ɘ�'9�s~jq%� G�3���"w�����ܓ����.kX��`�H��@��M�j�<�;2f;���8��5�S�i�:��.�NH3�yw4��gɩ~������sɘe�{vs?�r�Wv�B�T�*�DQ��������-�j�=�S@���R7�	0�Jv�����s�.yq%�z{�ϓy�W������1��R��Q�NS��N��fc�>̬,�9�ē}ݭ,�_��<T���67�N'Z��hݳ �W;��B���g���� �4�HX�Hh���<��=y�0nـTG�HQq�IB踈U��������;pgy��]5u�舋u�]=�}r����8p:�=]d|F�֙ζVGV�Ls�]�P�W�ֵ�̳��\Ka;#{'].Վ7�4�F��+��"9�c]��:�r�N��<t.QwB���k�-�Nf"P^8yƂ{'9�v�Z�&�uӱ#�tO(��Z$�=��(snz�Y=� iS�O6]��8�������bl]Yc���"��M�K�g5�fCXY&�3Z�A�<kt��N]�����˘���s�v�v��msÐ�$�
!�C��������=���K�I$������`�W�T�UF茕U*���r��qs�6wv��;�ZX�;�/�\\\lݘ�����(���� ﾿�y�0؉��u6�`S������)*��I%;��}�|ց�YM޲��Y.4H�
"$�����G`jK�w6��skK޲���c��G�����'ѝ��)���v3W������8M��9	t0�� �qƴz�h���=�)��3�\��fף�:�q�Ѹƥ7*I�0�l�J%�U��JT+�y�0�v�;��a~�\RͯQ�M�@)��?��zV����e4��h^ISD$�
	1�Hhg��Jfo�G`n��Xw+����>���H���I#Zu��>������wkK�Y���{���殷Q��=��Nݦ��� �� �'g��{-H����Y18�c$p�G ����=�V�v�?s��w6��>O���T�*�B���>�V���&��kc��}ͭ?s�ͭ/�9ė�R�+�'TԁT�n!�,�W��>��v}�C����J�"�.�O�� �v��9�T9�M�o �qƴ>�ߗY��@���{ְ��{���=8�cq9�J���+˜�������`w&c�9{��\'��)�8�ĴBD9�����]z���*1�!��0+n�bI����������쬎��L����Zh�R_!&�PI���=������\�l͛�������ea{�/%�<l=UR�*7DdUUQ���;�ʦ���h^�-��*HQ�N��Z椦������i`~��S���D���T>]�>/��u5T��E
�Q`w2��=��}��O�7��vw+u��8�"���qw4��ćn��3������ ��h^p$���'4abN���@왎���a�\���ZX�]Er�x��8�r-��h�����h�����q/s���C�?"z6E"�ʒ�;���`w2����nVӰ3f�?}�� uDƤbQa�������r���ܙ���.q�V�>�m��#Q�EUTX����\�K������{g���+�.y&��4ЅŊ7�5�'*J#eII�șk�5#���
�^ώb��^�����m�LcD�hɹۦ5Y2p;�a�m��k==&q�s�ݷCs��2t��7�
��7N�6��6)í�83�s�.�ir= n^:�v(R�Ch�eL���»;d�tM�no.z��xg��8�mv�z#M�ۗ���Ea��65=����8e.�:��5�jۭI4Kmֵ3Y4qꂞH�4}o26}��0�Z\�.��T�/ ����j�ٮ�z�݅��48���[���N!
������p������""!zC߬�-��|�,qDc�QH��1ߛ36��>ܭ�`}�1߹��q6|�\>�$Ƀ$���o��@���X��]��������:V(���
�S�Qz���m;�7]�����ˉs�3oK�B��NE$TJuR���j�/YM��h^�- �L�.����ݫ�}��v�#�r<�1�9R��哇1�v����x>�>���p��qx���wYM��Š{]�@��b ���RJ��v`�ل-���V�R�H#�T E��"!���@0�l��R��W��;6n�;���$���om�9������r����L�g�M�}>4~���;s�Q49�`��;f���?(�����\���ʉ�%F�E8ꝁ������9Ėfޟ��r����L�`b�hi�W��h�^���㞊�]Q��)���kg�LzۭZ���������[�D�s<ߧƁ��b�=�ՠ^�s@��.<n�d�D�	�@���o߿~H���`nn��?0����ŦС�S�4�H��-�Қ�w4���a�s��Gm����QЁ� b�����Vn4��a��,��#V�c�`q?_:T
�\C6F0�P��!�Bҩ���Ȇ&<�>L ̫J��w���^k��،���7�"A�@"@ W�&�8�Ja#�F!�7��I"k�ɩ�閖1P�p1�T�M�O��=+���^ tE8������*� ؼ?  ���t�t;��������@��b�<Y�+��O��nJV�s���{�`{6�X��������S j4b�тs4�JX��9�o�S�پ��̵`}�����PYb�n�՛uL��������n����OVy�_;P���0�q 窳�kw�� ��,[x�$��>�֦��9�F(��H��]��?g����{�������~\I�6c5Jidk�6��߾��/�)�y�N ��,�w�Sj�M����`}
�������s�=�%P�"��mÊq6rw��';ٮ�c�<Y&7�p�<�,Z������Ӹ�s�s2�t���:�TX��sc�q$�.��؋a��)�q��#������s��VJ.@u
*�UU?��o�`�ŀ{k���n� نO"�SPp��nJVs2���9�&ϻ3]��mm;���W���H�n�MH�9J���5������9ēw6Ձ��j����h��Q�J��v�O���v�͵`w3-Xo<�\\S�{�`��z�J�:q���S�>��v�9�y��9��N����X��v�j�81!T@S ���� L��1H�b!w=�����6��]�Lmt�t�8�����8��͎.v�q�{rmٻ;��u]ѥ鴎��q�}�aO���rmzۜ�Z�Y%��6y��6��9�Wr�ZC�҇v�������(L��vyݐ�m����V��x���i��{FԼ�uk���gV����ݧ���S�g=)���C<�Ζ�w�x��[�=����%1�����}��ۗ����#l�G�F��o=��{��ww�}}��9̝�X)�ݭ,�3��r����ù7]��.��/�dơ1@���;V��Yb�#�'��w$ﻯM�U_�Es'}�'�<n�d�D؜�@�O�yڴf�����v�Xm�#n�q�Tꪩ�{��9�<������j���1���-����ti�2	���׮,�Q
;������p�np0�?�������7Wg6G���X������Ӷ.n|�ڍ���)�T�v�%�9Lf�`�������M���?�`��Ŋ4��-޲ž~�ّ ��-u�w��7?w=�܇}�ۚ��ZmN�$�q1�ȥS�>�Vs�j�K��o�7]����Z���91�k(�[�s@ަ� ����|�!N��� �-|���1�LP�nf�篪�?���޿nh���=�%��������m�q֓n�ts�9e ol��n�����ܘp�Z����Y&A0NE�{l�h{�s@��Z�\��vf��Ц�#t��E�y�]�޻����@��b�\�g_4�H�l�ܦ�`n�ڰ=��p#�BR�[�s�o7� =�� t��&�brR��'�k5�ݭ�`~��j��'���Xwu�����i��"�=�X����<�ۚ���`j\K������: ��"��ֻD�Lv��l��4�!�J��5��������}o�^�$�q1�I�u��s@���篪�-}qh��q8��j7��i�+3�j���vf�vf�`~��j�ēg��ռ�T�����%+���`fN�v{����j��͵`}�]b��q$�,x��@��Šy�S@����d�"o�	t�ɫ�M~�.�-��9��m�WNЦ�#t�URRv��a`{�[����;�5���.��x��V�	�T�K�\�,Ǘ�P�:w��介��rp�,�����|�ٲ(%�:������;��̝��%�Ϡw}^,��R ���&�brR�>��;2w�?w+3�j�%���E�F5�l�}�b�=������=��- ��nG��G������������;��x�ef�`kŨ,x��������}V��\���l�&P�IB�#x�$�}��w)�d��N�un��+�͵vհ>ݎ�.-���Jc�l9$
�ؙ��.1ɻc8�W9�;N�
Qo/4J\�ض�P�h���y��X$�=�ۉ{m]g�=�4��#����[�Csc�][�#b����������DKʅ����wmìv�'P�:�]uYu�9��eh����� �ծ�X�Mnp��SWW*Ы�I�	���}�w�{ߎ�[Ƚ��E�bƞr���aӞw[l�G�N6�v�g�gfn�ݘ��1f����&5	���P=�������YM�n���\x�LI�&��Zs�@󬦁�s@�����^IHui�(��%2)N��JN����X�2՞\o�3]��3S�>k��:�Qa�s˜����/���w>��:�h�����J6�73@��U�w>��:�h[w4��ʱl���?88��Gδ��Jl�v�z�1+V�v��>�\��s;|�mF��$�x���@󬦁�s@��U��[�I27<i�1��l̈́��_D(���X�N˺��/t�p��#q�@��j��������x�5K������b�54h�SE��\���D?�\���`k����a`~��Vfc�N(��j)P$�v_{�X�Is�I.w}���w������=�L��'T萨���n�H��u�aX8��vh9�p�9kA����N]+ƞzP<�D��m�����}��۹�{Ϫ�9w\z�����Oe��TX�2����\��y�|�{�Ǡy�S@��w�7�C���~�ݻ�~��t�����Ȕ��"T�"�*���ҟ;�gM��@C����]��z��>����w�
W�mF��$�h��=β�������N�vT���(��R�w+�s�\^K���w����=��_{�X��ǘ;C�iw�j�����Hӣ	�[>2���X�H�q��d�\g%ح�m�W�ifߛ���;f���|�DBK�?�� �=�j��!Ӥ��`gr����!��T�76��?fe��.q6wwK��8J*DIE��3T�3�XY�ė�wmX�ZX|�TQc��B����U�>v�ͼX�l�܅BPȹ + d�ih��7~Ǡr����Od���n���0�� |�ؐ��M`ׇ���o�G?Wiv���b�۫��\铏�15u�b��)�[�6߿���X󸥁���˜K��n�ڰ30t�C����UUE�����S��ZX��Vw+�9�&��I�rUT��㔥������ܵ`gr��1�q=�����D�`���������������ǝ�,5{��Oo�x�:���y2`��������*�q��� o�,DCY
�b�"�����h����S�̀UVR~�d"�=%���|F��M)�ȩ�>CBD��$H	��P����9�B����+i $v��_����ր��AӴBo��� 8�����?8IjI����<�ȷZ�v�kHt����3?MY5�h�lm�n� 6�am-�8lޡm�`]UJ���B�g\�3��L�G�ڕt;08�n��-�،�H�䶕Px��6�+���h�%�thb:�� �����;s������RIĔ�;봶y�;��r[���)tK]�kl9(���(��͠bD
VL��am�� �tO�m6�%E8�pv��30���5��#Y�\�1�v�ymڜRDP����˲�#�90s�c4�pd��9 �!�����ٺ�]��d��1Ԙ�i	��c<kfX��8�{e⶞ F퍮T�5���c[v��]l>K&]{<݃�[����V�eՊ�	�Fj�H<H��/��٠�n�z�x2t�� zz�`�\cU�N��8&�qq;s�)��m���F��lܼ��9Ɉ��Ӽ���n�[܉A���7:<r�A�Sa�jݧ��p<�+m�d����@X�j��m��a1N�іj�݀2�.t����rsp��:<n	m��s�@��{3�[�U�mr���Č#K����t셮
��8.b8������i�)�6�Ȋ����7r=��utEUT�m���d%�G������	�Z�{.�Ѻ��T���C�ݶ��� b����*��mF4V�H�Q�Y`^Zڪ��&�ͱ��S�5^�`A���Ԫ�����
�]�{U�N�P��h#�I"Pm���9�d����9�lpl��\%v;E��#���!�pf�a��2�NqT�)�Z���s�yy�5*����	�(�zۜ��8�0+�T�^Ȼ��wgX���e��Ty�P��ڭvn����v΃�6i<�I�>|Fja��y�̛W4�5F��d��T�0Y�<0��.Ƈ�5ќܪt�L�=�ˀ��
G��#l=a'��\KT�:W0g������\]UT$m��SbG9f�v'Lő�@��'�\�h��x��Gl�]��d`*@��ɹ�g�
�mQ����w�)���6�* |������E��G�(W�Tb"Ĉ���g�&��8PE{�;��9'쟍;I�Ϫn�qgω�g�a+Ӗ18QFj�ח\p���Vy�u�Vm�F���3���\z��U�v:�]a�\��8�h�Ŭn�KŊ;<���e8�0r�;�H�:v��K�n9e˘2�Q��d�f�P��=MZA����c����cj0E��j���AF��9�{I@�p.�[m͞��ҫՅ摓r��D�,/Jt���|��O_^J��=�<�*wnn�����v����Ѕ#����*��оp�SN�Hv9����m������������Z�9�qq}���`n/�<y���y�c�/;V�o]�;����;�^�l��������8��>����^��W�=���ܵB�"��#������{�zX�5K;3��IM�ߕ�����mS��"��,y�R���n��n�ڰ3�XXŚ�w��9�-�QMPj��y�ܽ��e��WG7.����9�l������|��S��x�F����_�����Z�3�X{����^�`gv�UU܄�u!6]��� �<Y�
��""!yDbZ���l�5X�ns�)�T��**T�N���%+wkKw�-v�޻���^65<X�M��<�)`gfc�3;��7��m�`^ψ�|�j<���c�/;V�=�Ē���|�V�<�)`otCX.8�5lm]� �'^u�؉��8y�]���9Q��Gg1�v��x9���e�z�)����`gr��1�qK;3�ߺ�C�7�፣s4�S@��Ǡ^v�޻��E�Q|`�Y�a�kSrO_w�nI�����h�
� �!�!��!H:H��H@�� �7@t��!��,�`Z�E�*����q�Rü�8���ɻu���͵`feaa��yOW��X���R��B�0rE4z�h�M���m��/r#���I�d�,��?,laGM�l�Xƌ\uly^�d-�)��-���It��%/�n�i`c��fVI/�7smX�TR�Q�N�nQ`c�◼M��ZX���̬/�lέFk��C�*R��֖gr՞��8�����׹�X��Yb$N*�]�Mـ7� ۶`u�XNb���Q���7��"fm����SUk m�0/���l�� ���.�z��E&�p��Y;;1��[}�m?[��=Y���"��n�.݄:�s�T~^�`fea`fw-s�ݭ,
���qDc�,YI�z�S@��j����������8���g��B��	Q���R�}��`{woO���q$�=�R��������P�GJQM�J�R{�zX�5K2f;�=ɾ�|�{J�@�h%S�7(�:󸥁�.$�ku�76Ձ����m.�	@8�K'�d�I�5.��n���N7�7��ִp�cM���an�swOk�a�Ɋ��ѐ� ����ְnxK��;pq&;9��6kE�ػ�k��ع�<�f�ft����=r�n�^s������.���)����1pKuN{ۀ�FC���b˲���J�FNx�\K�������7��[��5����i��9�;t���#g��3՞Σ^sT\w���w��}�ۛh�v��ٛ����㞻u�,�+�ۅ�=���NCXq�����&��A!Ĥ#�����hz�h�Xq~a�sT�>k��Q"r9�-�]��)�r�q��V��e0ILG�6�M��/YM��)`�{�u������+mS�d"��,y�R��f��v�m�=ͽ,z�=��Tu���R�}M� �<X�l��j�Сj��K�;�v=���чՅ�.�:�
�Y�ݑ�7u,�{i4���Q�s&�AS��m�;����;�{��nM�`}�ݦ�MTt�9)Xܬ.��Ě��(����U�{���� o�x��X�c�7�p�*�q���O/$����Ձ��x�;���a���iĤ#���ՠ[�s@�e4
�\z�8��wx<q)�-޻��.qnm��{�����������G�l����q
��<Ȧd"�;]b.�����Ϝ��@���(�ۂ��۔�-�`�e4
�\z�j�-빠wp���T�d"��,y�R��\�8��R��;��Z�3�XXx�<�Q���cm9�@��Z�w4����!@ 	�g1>���?%������<4��z{b��`1ƁI�X{��9�'���X�ZX󸥁���@����<��nf�z�h^���ՠ[�s@�q��bʜ��j-/:�7_�����2ǅ�E��s���1����w�݋O.O�N٠v~m��j�vf;3�j���a`w僨�%7Cq�ꊔ������j\\�$;�J�����>��W��6~|�qR'Z�}��z�hw\z����9����a���ryO�T�~����~U�>���F�GD*��Y��u�3@�xD��Ș�ǒHhw���78�x��ـ~J��;���������76s%��"�Q:�m���s���t��0�l�l_ϻ����}��4X��cm���?���@����/YO��|���@��_B8�r6�R4�X�x��ـ9�j�����P��}���:�L���IJ�������\z�j�/�w4x���9&l&���5X�np��`}�%��~4��Q��Ġ�PR
Lz�np��`�� s��`�(i�p��vۗf��*-�T�umL���!i9�\qV�<��fiv��\urCF�v�g�r������D�ۚ]�ob��p>�S;/n_;:ӹun�	hp=p��#,t`��tnLڍ�żi��cu����pK=���w=;3l�q��s�n7|�啐��4#ˍ�^�k�:�aZ:�G�]<��5�k"v����5�O6���y��LQ�����{�����,~v��<Og��͜<�k��!�B�K��W����%��&��r<�xu�����9R��7w-Xܬ,y�S˜�?0ܛ����KD�'Q	�!�Vw+s�3�1���W�ė30t�C��pl�UUE��7T�3�1ټ\���K����Z�=����y%(�R(���Nc�/;V�z�����*�q��;� $���N-�e�˜�I{}��yＥ����������������빧��^-���ƶ�[�77�6|�vb��㳙۵78���l�����]n=�h���-�<O��r&�N]n=3���^n�0��|
*������`}����V�l�4u��Pӎ�ꓰ7&�;���ԛ���@�?�Šx�q[ƞ&�)�-��qs�S}�|�{���̙���1�u�L@xbhs4l������ɘ��2Ձ�ū�f��UE�X�b4�X�7�,�����n�p�=�ny�i������������:�5o�������-�j�;���/YM ��ncX�EܒH��S@�s@�e4=}c߿~���{��$H$����UY�s��X7l�P�{�BX�o��N����|ʟ�GR�OȖ������ /�h*� Y"Z����9�Z���#�u��$H�`	 [�nRq����;]U+@4� <٠>��!��1$!��y�w�K,K�c|%Li ,36�# ��9���X)wv�ۇ�`�Hf찰4��1�KrS��?j5��H��~Q�6�u��W� 0֖��4 �����8DQ?)���s{�.���v���ei~M�j&MNT� �����_������l�����������E!65'	T�1�,ms��9�f��,��`�}��I��]=��-�%��s9L+m)u�3� �8��N3�WH��յ�芪~7kK��Z�;�Xo9��;�}O@���6/�i�l��5!�{��hl��篬z�e4=�)�(�	��V������k)ټo�����ݵ~M���-�q5N�������!N�Ϯp_���,�n}����%\_��8.}����7p~���S��%S�N���XY���o��~7�����K�u-��51��S�9$��'`�8�)�,�ԝb�F���<�`�\�[��&�m)n�n��YM�zX�z�h\;��#� �����{�a~��sk���W���Z�&��*$���&`�B4�4zϢ�;����[��{l��iE7�&�E#�v������nڰ>̬,�N�K����ƞ'�%"���[��fB���><�?���ـ8Iz�#��J��cD�Րcf�3J��ۀ�;���yF9����vx/-i����l;����ʓ���r�cy��n�R��M&��H���8b.͸���ew`�D�S�-�p�cg&�r�֐�ce��~�TO|9Ku���mE�Ƶo��f{F�I��[
�ż뾑nӳv�
�Q�m�vZ u�,N��by'�̑/#t��D�\U���;:r#8���v��Jy�F�I�{�����ow{��Ɋ6J�II�a��j�3O���G�ڮ��9�GMۋ�d��d��������n������Ł��ܩ`}�Xy$�0�nڰ;��[��j�!�� ��l�5�f�o��,�u�&��,�N��h{n�����7mXt����짐�Q
��M&�4=�s@�s@�ӥ4m��:���cY1�I�h��X��w�?�����2��>�p��k�9���,�RΛ಺��vv����d8��n�up�e���̜;�h�6�cxv�[�`ݳ�/�Kh%��,�4u�h(i�J�(�>̬.�ńN�Qk_�N���G��QVV�|�ŀo���!�)j���Mښ�0nـw7��
!&���vwkK�e,�����d�,5y..)��|������2��=�S@�ڞ��4�&$1�u���e4�S@��)�gm�p[cz�Ї��W��;����Ep�ͳ�;;n��rh2r_�����U	�1��_�;�5���~���%����f�Šw}��n14H��hzS~���3�ZX�[��N��\R�&��#T�Uܪ,�W��;���?D�� � �'�m�9�~'���`o��X�J��24��&$�u}qh��hzS@�l���(��������"s��}V��,ܽ?�����N�v�I>�5��Wv�]�Wel�B�׍��WG�
�+�m&81������)�ccz.G��W5\����0u�N�����X!D)�TX�+�.)��'`g��������n��)��8$1��߱h_U�u�M�Jh.�)$m0R5��)��~�ع��^���s����,IH�Af�B0I��'�4�;7�@ڈ�foޗrO��_�d$i%"jE�u�M��_��x������.w"0���d�&�d��z��a#��PȸՌh��V㍜�{I%����M(,c	�	�x�ύ��ZW�hzS@�x�ƪ���I�8h]��=���:�����M�R7�e����E �k��k<�I/.I���`o��;���OƱ�y"�qhzS@�Қd���mf���-��	B�d�,�k��mn���6X��$���8���N��䦤�	��8s!�9�9�M�7mWp7S����D�Xf�[��Ų�2#k�ۋ(ukY�Y�ؕx�l�ی����o�k<n��[�=b���5�D��Hй��]���?���Ƅ��cԵo��a�E؆���V7K�ծ9)�Ͷf��'�a��6��
�S�b�l&8�ArWon�����m�w*=4,���-�ڹA�ueП�P4��|�)%�dٚ�5)�km��9�֘}�8�ls�����wc�Ƈ��;�"���J|��F7�������?�sg�3r������V��3GUMҀ�NH9I��/y��!��Z�=���Ž���$��4���G�wW� o���mN ���6�T1��9��)�{]��
�YaZ�f�����I�J*����mN ����X}l�7�{�x��lWi�u:nvǎ�X��m�BGe��]=�q��,ヅ'me\ulㄺ��N�ǝ�`w�������ٺ������4�"q���;���s�R\K�.͛_}7S�1�r_�>���
��!8�ܥ`ov��>ɘ���o^f�3vՁ�;��U#H�$R��q>�f��י���s-X}�&߼�@�߅$Jc#X�b�Z]ΰ��`]� �\��>P��L>(��nz:��ێi�
ݢ8��Z�Dd�n��tٝ�tk�}���_vbH���U>w޵`g�XXd����qגG����!�,c	�s4l��>����K�̵~K�����q�BU7�,����;���Z��I��( H� ��A`�BՁRȢ�<Q	���~��;�>4�#lY`�,ML�)C��<�K�̵`g�XX{��IqL���-�?6/�i���8�q���h�)�{_QhwW�yC�Q�}�ȓ�7lֶt94e!"��z`��3����������(�ۡ��l&�������@����*�@�s@��z�#x����)UE��N��˞K��Hy��X���>����1�hꨨ@�Q�#��>V���w4��=�����x��P�����U,<��y��X���`�8��A(K�r\���K��~�~��`yi3�ڎBd����e4k�-����w>�~9?��V[�ݙ����O�9��ܦ+[�����w)��T�8�:-\=�vQWs4L՘��N �y���/�~���gƁ~>#lY�i �d�H,����X ����8�H���M4�I��@�s@/�f�b�\o�3G`k�l�?}��B�% &���������@��^��s@���fF��$Ɖ$�;�Qh_:�5�� �xU�	%�X��#?D��$�a��]�� ��v0�C�,jв%-eDhC�Qt�0��/ڂtp#Ϲ���e�]�RA�`n�A�#�y� �Àh
@�R,�i���F�߂M���%5�C�3H����s��a���[��k�}kՐ&w����??$W:��� �"Ȃ �AM!G_w��]��>�?~�][PM��epAKi�im[xlth m��+�0U�k�n4vh4���ԱMJ�s7;�Mö�k4Y��DYg��8�&�c3WC�ac��]e��e�x5�/,�i�>\�;tV���ƛpl��ѝq.�y��V]�]u
���hi�V׮mѷ*=`��D�)� ;S��(����n�;c���;:��v�wl�]h�N��r��Տ��q�*��Ahb�,�ZmC�:zi��҄L2��d���[��mq��q��R�C��B�N�pn��[�ԯ]p� �ltE�a�x���VWT��q�a�3kM{vR�W7�psE[�Z���;s�3�e�l�ms�w�,]Z���qq�n��۬�+�+�c���P�|;���`.J�J�4�Y-՗4�g���<mxN�x�[md�֋n��Wq�e��v�i�`���n��ku�k�����eZ�q�i��7�˵J�V��m�rҬnr;;���v��]���'n�wl�`�td��@\=��|��/ �	eq<ݲD^'�GA����}�}�Iĝ[9��R[<��O\�yb��l�M�K-�J�ϝ��7%�LS1���-�\�^hԛ�Z�r�*�:B�gnq F3rt��]g@J������:�b�.�C��;GY&I�V��j�DR�Ӛ�H"�j8%�c��8[d�Z�M���G�n%��ͫk~���M�v�N,�m$;vūڍ���օ)�sg��6�Z��%�&�r�ɭk.�ĭ�S�Sml��l�*���=��۩V��q�RdUɝ9�EB��Z:ݳvL�.��ZzGr�F#8���cF0��۞R�:vw�����JF��qYm�>KRm\m�*�i25\�/U+�@^'��d��1�g�ut��kg���y��*]�����lp�@�9���WY���݃z+;����tUQ�9��F��;vY���w=S�aMjēˢ�$�4kZ�Pi�꒮�M��	Ӡ K���Ԇ��S�
�QW� .�4
��=�PR&׎�
qD:�u�4�@!�8���@�=ڈ4��h�������ên����V�[�h%�oO[tWcV��j���gG��֣�ȗ�r��*uĜr���s�߷Ѭ��=$p�ɝ��+hwn5v�G��]4�cM���ݛ�T9��2�I�}��z�62ú;쬦��tvSh��ɷ6��������ʛ8����G@ T�y�2��@4����ut���KY���Z��̒�5��fa���i��Q6o�������us�î����6:���5����e,͢:��k�3���}=��LF&ؤ����z��� ���;�Qh��8�d�$����w4��{;��1�r_����ަ�ppTRj�7)X�׋������z�6X��Vgp�N)Q�U7@�{;��1�rXfe�$��ߍ�|Fس��8�"�ZW��<�ww���V�����d���3��8���h�w���{2sF�X+����Au��6��-�xC*������DKC��s@��M���Wuz���U
���R�3�-���y�٣��b��޳��rO_��nI�{��˜�I��͖�n�QnJ�,]�Z]���w4��*�H�D	TA�T;�{36X��V��hϨ�}�X)����r=�n�oJhl�h^�@������vx}��ne2��]m���A͵���l�a�Y��϶�D71qRnR�3;XX̬E��;�y��3r��>��l��Ʊ0r%�4�.�I�^f�7+K>���6oM*H,�4�N2E�@�[��:����3���S\��!~�%�ooj�s+Q`~x`���q�D��*X{�.'������|hz\4
�W�y^q�	Ց�!��,����3r������zS@�s�Q�j���A8�MudU��n2�by.��E9{F�l����+�1G���I�K��U���)�[ҚV��$��bm5)<�K�.$ٻ����������h��H�D�$����������7�����6X�&e6�#j�ҕIʢ��\\\{�zX���������b!� PT A�`�@"��"��@O��j���w�1<q�L�@N/mǠUz��Қ�)�\��*=��Y�W-�[�0�H�7jZ����Xݸi����+�q�si獙�Su�9|� �����`kj�K��\i����'���M�ď���@3���yܖ�!�j�B`J����a`��7�7�se��������f(��Hc�$4�\�W��:���oJh[T��fBBIJ�yܖ�r���V�����6a;;�:[-�l���IY1�|_�)��DOK�=T�9��z`��rk�%�
�dڐJm^8��-�H�N�9�Nb�����ɸ����d�[mݤ��h��.�ۉi��v3���=�<�FNb1�����u7{۴�s��j�h��B������{6���甠q���$�؅��K�����H:�t�<	j���v��e9͝g,�_i33Zӫ�L����/��&}.����|]欞7UGn��:zP�[���9��9`r\�[��vΤ�T�6�����w���,��T����ǝ�a��{���%�,�Lrbr�Y�z��*�^�ץ7䏾�1<q�L�@N~�d�*�^�ץ4_U�_J(��<@�E&M���za`fN�Ը��&�|�����9�M5$N=�Jh��@:�ɠUz� ��YE���&������q���\�n9Y�"[����-�3��CFλV���a�x`��x�Y�z��*���:٦����Q�#X�ǒHh>j��J"!$�~�.^}X��� }ҚV�##��blm̚^ܖs���ɽ̭,75U�߲�SuHH�%"�C�_��h����\���^�}1��,�Lrbr���K����l��Vϭ�����,�t�n�[Wl��A�������dk!��y�mЮ�$2�:�y��f�qWu����=:�`���%�h��V��O�G��c�1�Rd�<^���)�z����\��Ҙ�5q&�jl�����9�� ��u��R%J���I��G� |hC	��"�������=�V�K�ӔTL`J����w6Xnj���2Xy���`}���N�
�4�*�Xs��ӭ�ϭ���ܘM���r��OF�M❻W�3�\y=l�GWg���sa�����L#�=Y��u�����zS@�{��^�4��q���H�#�:���$r�����&���נ_Lu�X����&)TX?���;��Vy&�}ݖnV���lq�L"���C�����a�l��V���
P�,��H�%$�c� ����[jXB�V�䒍���X���*�]�%M\�WUh�=:�`�l�6w�`�m�?w���v��M�b`���Mq�{�Wi�&,�M��h�Y��=�w���p�}��MA���?�����=^�z�.��^��<� �X� M	'3@�{����h/mz�w4-�Vb��F�qʕU,�V"���̖oM�}��˯�@��TR4���%�9���� |�,gy��Q��>F��}���"$�@�n����`��`�n�S/��ZJ�<{��{o��w��ɻ�%��x#�u���:�i��͵�Ǘ��eh�!�����t�������B:�k�iy�ӽu�k��.9p�x��0�w$;�tVn�=f�Ѯ76*�Ygm�wUK�s=��:�ܪd�护(�'6��r���V��b��6��'nD�M�t�VʨԦxC��G���H-N�g���	zxػvH�eWJ��U�f�n�CQ��w����<A��Yr]]M\��Kf�N�����5�(d�%�b�<c���b;N-l�:�ۘ�x҄&99��������h/mz�w4�M���X�8E�R���b/�6|��,��V���q%��f�#Q�N��L���X>�Հ>o��� |� ݤ�4�Zn7!C��*X{�Osw�:��,�V"�S�wvXdZpNk��� ۔����`y$�����ϻ����Z�){�Kzjh䡪�N�2�B�:�E� P;<����_}���.�e���d����1�O���4�>���a ��s�;�d�����RN4��%�9����׾~���v&�F�'w�Ձ�����V"���9Ĥ=�O��SICi�2������X};����b,���Ƹ���m�"���w���/Yp�<W��:۹�[�ُ"���S�hl�hfg���~~��j��Ӹ��00MJE�E!�J8���c�^�oD�v[�m�k�%��Ë8�r2�5�bN6�Ra�x�W�u�s@�U�^��{��1<j�LM�ND��/[��<��h��h.��W8�g��@D�M�V�3��;h��H25D$*D(DEЕ@�v�9� �O�B'�i��E��`B0�>z���$������� !�0HG����2���|P�yC��8������H	�'�HJ�� �B��sBl� �]�~?7���2B�d��1c�>���M��$D�4X�W���B��<8~\Np����ہ�t�#��͙ �F���
Č$$6� �m(C����L�Ѣe��o42������)�,	)(@`1���*���D�?b��b0�����_��?D� tK�����!,$
�)�0�i�㿴p�H$>S3�$9jB-/]�+1!�с B@����f�"�x
|�*�aT uY�s�
i�~�J�r �κ~@�!�D����S�TP��e��g�,;��Vۛ-��p��N9*����{�z�癲���Z��.?��]�׹���hjR�m�H�?>�%��s�����k�����0h(c��HT�ݖ��4s�B�h��ss��ɨֶm�۩f�۴�5	�8�cpR1��m������ˇ��=V������ �1GNf��>�@��x���=���y�s�M���ҊB� J)�%S���F {����X��� kM�T�	'#P�a�wY�{m��<R}�������jA�� B2H4��B � F�%� ��A�Z�l�"��#�u�\���*�5�����>���c_�Lm�M���=���=��p�m��x�>B������v�7Z��H�Fmx�<=�,7b�9�l�r='3��;�å6�.0��������r��;���wwmXf�I��Q��rUU;���^�I��3j���ڰ?vw�\\�:��T�	<s�I�4�~�����}V��e�@��Iā�ғ�h}��=��y`��8s�� �s���@<$���'3@�U�wYp�;ܫ�̵`jH���F�$���ҝK� ��nݶ��zj��؆���wOk��ڮM�V����ޔ���*�͹\�^��I�o7���cɭ��Fɍ�Pl������BuI�<g<k��n�hÓ�{m��&L]6�����q�]��X������c8��p(�$��/]bȮ�Zm���!�}F�"uv����a��������;r���{M�u��u�����p#�Z��d��i�
� �s���o�WV����ǉ��99�͢L]n����7�;Kj�v��W<�;:#D�ͷ�����m ���w49�Z�Q7�АHr5	&����w4��Z�\7�����|65�d�8��vՁߧq٩�ݭE����`~���O*k�0Nf�޾�@�ˆ��^�m���k٘��(��ӒH�ݴ`�ΰ�ŀv�9�5w ��}<�Nٹc����u]�P�r�J��t��ǎ��f�iv9�ªs�z��w4��Z�\4�Ȝ�1�	)�z��oy�����C���mEHss~Ͼ��}�kQ`~yܖ��������'R��^�?� m�F�|� m�Xoq�dX2(�LjE�[e�@�^�@����}V����7��HЇ �a��~z��h��l�ho�{�w����;L�0��ѩ��J�U��vQxoX��N ��Y� "�5�.HÕМ���}�ۚz���.��z�q�<���6`���}V�m��z��w6�${e{3��rI�m��z�=�� �1:���.s�Ĝ{����3]���a%б�1��Әh+��۹�w���-��^�E$����G�ffZ�<�����ݭE����,���ݾn8/dm�s(�odJe����%���dܡ��f��g3�Eh5��6�V�ms��m�y� �x��	q�d@II�H�_eZ�ے���Z�>�w�~`b�a{N�m9y���z�w4}}V�k�@�����T&6�'#q����N}��w$�s�۹(��ø�'�N �3�����ٹ'O9�ɗ)�r�����v��X�����`fw74��C|0����"n,Mb]���,�HyK>��T��c�K�ma`��q>�,14ܒ/ ��s�x���z�hz����M� X�16ۙ���u�7��s�7\���DL����H��I�����nhz��>K�ϖ�����=�դH�o	�X��� ۶�Ӽ� m�X���<�	"	�Z�\4�� m�X���q�Q!BP��w�_����݇mÙZ9����@�lh4�4�s$��e������;�%ڸ˹M�ɜ���{w��( �m��3Y]��q�;��-s2;��:��d-�6��,e�{v��n��mX����Ym����g��<h���s;N��(Mb�v���sk�� �ñ���۝��mM˟C뗚���u�8s9�͜J=9�3�ܜL9�Ζ�����w� �N�Ȝ ?}��\˭f�d�s¶K͛7�c�ڭ������N��83O��laa�DcƜ���I��|��z��hz���.����M��)#q�}�ۚ���@�ˆ����``�q��R��MZ�=��p̬E��o���`n�ڰ?}�.�u88���rH�l�h/z��w4}}V��z��,�bm����� m�X�s��m�
��~���ݵv���]n�d;oUG'FIť�2㬵���フ�hp\[��=��4�?��j����;3+����ͫ߱��Q"D�8�)���_U�~̂5�!��	 ��"Ţ�I����E�����O���rI���4m��;�w�+0��E�6� =�� m�X��� s�xӤX8��h�����h����.���lj�M&�(㫼��`��pݴ`���{��;L��������|ws���2Ì���G���e�nsp�Z6����\&�{MZ�����m�n��ŀ{�^���5�NI"�-��{l�-�s@���h��o`��1����F {[���a*!BKP�"1	��[��q[�����I���I��#ȑ�dē�ܚ��h����.��ˎ��D��q!H�&h����.���w4-YVj���� @����J/^9amԖݹ�����;es�۴��s#N���=;kH�LjE�[e�@<�٠[n�ﯪ��+�����N)&��lL��ŀn�9�vрn�b�*n$�O ��ɠ[n�ﯪ�ĭ�p�=�hP|~�\M1`���DB�����I�{^&䓟w�ܔLJ��C���vnI�ݝ��u��Rك�H�l�h��4m��=��Z�()��X�x�D�oy�Iڻe[k&��n`[���<'o=�a�'��0��69�ɶӘh��4m��<��Z�\4�ێI�bɉ'��4m�߿~l��5��Z� ��r�[:�����걬da���@�ˆ�_z��w4���+0�4����v�S�5�6X�������fx�qg)�r��N���rXy��qn�>�{��'����w$�EU�EU�AA_��AZ����("��(����H����(/�� 
� �F*�`�@��
�F
�P�� �@B
�@b�E
�@*��R
�T �DX*
�X��`�A��*� �H����2( *""�* �A �Db** �D���
����*��1��*� *
�"*`�F
���
�D�� �DH�`**`����H���� � ������H*`*��E�������E�����@`�B���H*��F�
�X��E��E��F�B"�����A ** Ƞ H�TP��������("��PEV��*�AA_�EU�U��PEW�QA_�EU�("��("����
�2�β^�(G������9�>�x�                    @<  >��*�	( U"��   H�� 
�@(�"%
 �   @   ��   #
 (� �
�c���T��Թ5���t�[�wJ���(�}�}���ׯO}�)9>��^�z���-�u� ��ͷ]���� 7P��[C�˶�-V�w��  �wUqoF�/R�+���Up  �� 
P $@%+��7g�ϧ˨Lvu�^���ﾔ�����Z�t�qgZ�� �=*ťL�/��y�JŔ� �>��ź���}w<Z�n,�� ���}k��ׯ]�����9�� ��(  $  �� 4|����� q(��@  ��PX R t� 	� ��� n`  %)@D Qi� �)D� M�    ��:  �P ` J �(+  � O=�}�wco�xz� ��8��m�Ƕ�Z���ԫ ��ۓ�=�}��]w���^� S�R�w������f�y�ǹ��� =JŔ��ז�M{{�]������ (  Œ��;�����5\�|��׷��[� }�֝�}}��ݼ��Z�{o/sV�����֮O;��;�� 	�ͥ�n���\ u�\]�t��K��y�&�׼���_m���J�k���z�7�ԯ�   4�T�%R�  E?�5R�� �<z�TJ=#L#&C=��#j���db41?�%�)J� h ���jR�D 4x���Ο����K�}�����}�.��_g�������EUWTQT��
��*�*��UAU��(�>��!i$~z�Itd�#�hb��c�Q�����i���5
�bha!�����4`�#u�j'�����g0=N1�{s@�B��@�Aa35��x�>c�������ߜ$�2l�!t�<�'$�)CC�����6ƺ7#�6s �h6�(�$B1 �><��O��<���7�a=du!��
�A�]04n<�Ј@p�	�� �td���H���*h�!'9�a��$�)N� �HJ:6��(��Wi
q�х,aL6B��$�2!�Z��].le4B�z�ńa�t���3z���z�7>ގdu9�=SA����B�*�l"I�{�B@8
:S4�Sn�C��<`ň E�!$��0`�;��8�+*AZ1�H��a')��ٱ���B6F5"�t���$�40,��DMjHK�8R��c���kD3A.o�2qٳN�l�:�J�����ѐ� ��p �A�A��i�<1�BGG��3f��!	C�#d48m���4�
h�44,�j��������#�2XJ�`@��l�Ұ
&��}����Դ��`�"�H�V@�d���v��$����p�����3!N�$n�Co�D�CB���$`D��-)SA�HH>!�P�
	��ᧂE�#�B��uY[I%1��2І�nݴ�M�;YK��i�^]�XP�����j�I1���a!H�H��tTrBH�����rGqK ���椉�����4� q 2 	P��|v{��HRg���g��T��0"Ut��C��`į�����zH��Ct
}��n0a�.�XB��3u�P*@�0��xSAD��D �]$�.��g
x"lb%WF0*i@1�L���y|xqĐBW@�b�0�Ab�XMD-Sd`S�!$t��E� T�><&���1%4`�"M�	�! 4�l�1�M<6�>�|0���AR�XD
c)� 8�%X(T 5=�����F��ћ������&p"�|�v�~᨞_�0�ˡ�c<�����Y�CHH?W�M;F�[��65`�G�n��NM�Đ�Y�@�i�"� �U��_z�&��"B"R- �x���8�>>I �F(8�&ӏ�`�(Pӎ�'|����nG�	(k�7�t�I�Mnn0X�L�]I�{���0���@#�B��@�U4�"k^�N#*B�HP�E�!B	f��V�F�q4�I_4�Q��"B!C�0��~����`���jb�}���FMc��@�
ƺk�d7#,�����A�
i�`@������0�k���C>���|L�� @O�-@�Mnp�9�<�,ss8x�y^x��`���#�ӡ�4h&�f��%�
%��BH����P�"h�R���f��]���� `B%H1D��N:�M�SXBY�7��g��i`U�6��lױ�rY�p�~ ��r&�`@<|OIa�wm�%Eٛ �!d�X�%���"F+���l�1����ؐ�����?�~�d���lp���,B� FBᰇ�<��O ��1Z2EH��!u$K�MJi��.h��'��I�2Fyt:�d�*,�AR��i��.�Ǆ�
J0�a�WL!���d�:�Cp!�R�y7�՚u�2��P�� ��SX��,k
:�w͜%�+5�f��0𚄤^a)q"ՉOH��E8��A���C�2��фə��)%,�<�����5t�G4y��!�f�t@���ys�n�.���t��E�$w�4��f�]��i�`k�0�	���%xOOtB�F��Z0H!�b6d�H�7���6R*����� %!��*����T� �U`��9��	��F���!��%4C7�wYZ<�5�]�i�01�J���(��F)"F��/��ֶ���xp��!�B���44���L�Nl.��mK�]!@`D�T�ɀ��m�'&��_Ns�I��IYYp�$ ���۱�t���9xO#�l�aH^x<%'!Q�f�O��I�����=�m�1���|8��]a<ֶi��҉�@"@'��M����=���,Gф��sP�ᰄ	u��u��9���
�	)��t�8{��ᄐw&�Cc�ǎ����5����8�9�)��i��� P�x����=��kЅN݁���aCFx�]����WC¸m6��<�5���N����͛!��ڛ�7ɬ�"|��{'�#SB#%4��7�'�EN|��5�d2�HI�)�X1�ӣXEta�
hI$4�_R0"�NF8�
�(�)'9<�����RGD!����~2@���5�&�!���8c��l���Fʐ��{[Z��0�T�yMA�6\��M��,3FK��.��f�90̼�BkWӄ9NSlt�$�7]�ͤ+5���H�#�"�d�(D�hAJ� �I�F# E�d���dp�%��n�����'0�;k��.��μ��h�eQTs�h|�UgiOC
�*�8�w�B2Oxh��Y�5��!<A��2�8�,	3s�%� l!��X� D%��+I�J�y=��]ۣ^�.�se�K�N�9���+�Dщ)�3˚9n��o��_>�&��B.�f��XEa4s/&�&�l�szB�$U*Ӂ�4etR��d9�!n����g0�ėY̖泇�S��< !Mm2�{$i��u�T�1X7Y����DGL���h9<n�P
E�r��&��5�&����*i	#]!�	<��o�Jk�>��7#���p�'����M��aCBF��	 ��d!]��:�B4�6��78x``��dL$��REdaa H�F@!"ج���H&&���>G�p�ts@� �cO�Ռ!B�g��G|���H�� 	�0�1��*���礔6"�d��oWf�U�Q�0�X%@� z�|~H���$���S7���r��lx�1����pcD"-H�B����J�7�%=�$e�J_����y� �%�bCA+�z�S'�6l!BS!u��L�	��y�����%H��	s0���Ӑ�8�z +�0�!�,��Lvs3Ƒ	�4��=�
l�
a��nIvB�L�Zatlܕ�js��M[s<������7�O�bzr�¬HBE��H!>�MX���<k<��y���|�b܇4c�7���&�5���☁�2E+!��P�f�!2再&�к/�4�A�BB�B�H����GщF\}pl �k�r�]rSQL`HB�#���p	t�'Il�܌��1)�4Ji^�n�' T;�xđ��<���������� 	h      �    �      ��       �� �`  8  � m�            ��l      $  A   ��  8 6��   8     6�nh; pl�� ��#�sam �m8%ȳ*)��pl�h 6�i���  ��    :	2�m�9�#[U[��A��r����-n��6֭�p�p8m$���l�qmi%�8��n�\-�kB�V�+r��Ҩ V��H�N�C]%�'��#������Ԫ�q�mηf�	��$pkX-�����|'J�^9lN�^�n�&����	m�KX�fR"%���Ү��*��m����J��a�Uj��e�S��=��75����A�N6�,��Pb�̆�u����SPJd��vMu��ez�����Ij��d�r����;T��:�*J��rmAүu]=�L��Z^z�����P�e�^�8:F�l�4Z�J�
ډ �6K�nݻmR�ۚ�j�t,�%lG[Ht�8Z�@-���*V`��vড়�N�nj�knI����D�	��m�KQ��B%���l�n׮��  �p��m��/�m� l��� �8  ��[R 8;m�m�pX���5���x6�Ԇ�;t�K$�u�T�u�p.� -+f�[p�8G	l;C ~���| m��ֲ��y[j���᪀��nj��]X�qS����   v� � �d�Hl�e�*�a����ɫ�T=m �
�[v��K���C]����p@���:b��ڐp$!��\#�-�۰8KZݖ��$�N6  ��2vN �&�H��ۯ^l�M!�JG��Rl��� �le�ຮ	e��m&w�����iu� $K%��d&�zA,�Q�l$-�d�v����8*y��ZWe�� ��sl���׭���/�]Tls��+vr�`�l �h,�e��n�Z���24cۋ�3]U&gb���^)�\EBEnqN�gn�A�٨l�\�����M4HĀXgX5l�@I����]�;8�N�l:�(9�5�v��A�Ā � ��⋚����[��� [���]":*U�`�ݴ��p�E��d���@[@� H�� l��I�m��qru 6�$�SI��-� m�����7v� $  8 �m  6� ����g| $m*���ko� ������8m�cm�����(�� r� m�[@   �5ۉ$�C�� �HAM�m���t�`��9m� l�j큶�l��֐ p��H�x��-�   � m��trI8h� �$ [@ 8 m�    �   [@   [��-�  ��  �c��ڶ� r�   $�   ����l� �:@�Y( 8 "� ���	6�`$��k�q�8�n �m���  $� U�hm�m�ݶ ���   T�r�*�v*��XP@*�QU���u(
jk�   p    K��kؐm�2H9"��N�m��6��L�v�U�  j�oI�䙧(���:M��N��ڪ��r��"��-�6�s�dK9nuLZ�Mٝ��2��6�[�oPv���IQ��1+�e�h
�8%`��m���kkm�    �nu���&ձ�l		  �i��l   e���ݺmvd
RC�7i��.�� wE�v�f 	jT��Hm8ר m�D��0Inv�l �H i����9�m�`�Z��ɶ����m��m   ��vRΖ���  ��*N�� �pו�b֜I �m�6*�� .^yX����
 �vm�d� R�յ[ �p�uC����M&m�"�k�6��m 	�ͳl��a���I�R�V�l� �$  �kh��3��+��IAj�H�͙6����� 8�-��[\��[@f�$6��nl � �܃m� ��ji,�$�Ȋh�k�`mY�  f޸�B� �NZ�mu0��$��v�V����/��rl�uZ�܎Z���k$6� He��&�p-� pm���`�`��ЩN�][�@R�c�fej��M�ݛvr��q�H�Y/m��m�m�	�zR�;]S�O��nGh�lM�	�J�@�j[�+���AT� �ԩٹ�V��U@Rls��T��tJ�I�mFփ���t��d�� +H�H@w�h"�UP&a�&켎��`�0�3�(�� j����͖!6Dێ8�y�s����lΙ��[���pi��K�]�����(p	$H��v���f�6�U*�mmUm�f���̝E8���U�j��K��6b�yiY��)\�LY��d-�f�$��m�7m�d������*���Ԫ��v�H��a����j��Ԗݶ˦�L��d��`�8  H�mA�[��H\�җԬ�/lt��ԯf@ �cZ�2�Nηm��p��� oP �S,䲷  	  -�l    -;b�h?}��A��p $4]� �8���6�I5�"����l�k  ��۱'m���n6�5���H86�������@�96��`A&-��k��^m �F�  ۵I���l   UP��ʵt�5A�n�ݠ�nו�  �&�5�m��!�6�o]���;��  -�m� .�$d �[d 6�Nm�]J��ʶ�j�� .�N:54�U�^Z����"G&�h�jٖ�gRL �&�Lߍ�����u�$m�[���Ѝvk��uQ���)eې�� jy4�gb���g�d�6�r��[Ut�D�U] ��]��*PG���`�IJ)s���UU<�)�B�vp�k2�U^L<��4��^��a��ڥ@jU�5���]�����I�Ӵ�e,�-��  m� M���m��M�����  	 ֖�  	 �H�m�` � �6��m��H��� ����"�6����5�������-�@� ��-   n�          ٶ H���p $  �  	M�k` m��l $r�AZ͍U�m��� h      HH�`H hm�9��Wf�m���'a	    "@H-�հ�cm�4V�	%�� �se���  �L�6�W���;l�ٷl i6��|JŴ�9ce��m h [xm�}>��   �I@ 	�kjG�|���eN��mJ�S˳�Vm�@ h�am#m���v�n� $d���E[R9�Uz�d8�lv�M٤\�H� ����s�� �4�M� 	 ��    8  �,sm� �m-�Zl Kn�Ą�oUJEʼ�����U �t�M5�gAYi�-��m*���[C����j�m��([@m�[A��mp   ��k��-���  mKtRC�׫9�H��m�8K*� N��	�E-�ӀD�۶ڶ��T�UQ�Խ��R坯Up���Q�8r+�U*ݵKpU6�g3YxVr�Ky"t׫r�v�-�������"�:۶̒�]�݉8[z@�N��u�i$�RiM�l�m�Z�J[[I�` lz ���!����@ �u\Y��@$bZh�H��0 d ݶ  ۶� H )[`�MÁ$�  ��pl m�   	-��l $�Vān��WV � Ĝ��6��:��m��ٶ H�am 6��a�ktHCm�oP$	 8�陶5l n�݀   6�   6��`  lε� #u��� kX  rKx�$�    6� Ȥ�J�m�� �6�m� �`m���    l�VK��Pj�`*��@��/5�"Z�W�W#�`⩵p9�`ɵ�`6��Ͱ ��   [[l�  ڵ��m���&9��� @�I���jX�cl �SeYW��Q���U��_-�R���Ԫ�t@9�������ڀ���WX��`
ڻm�-����  m[  ��� �qm-�Hp H  l          -�[[l[@� Zֳ2fI����*�*�~E���c
R �! ���()��8���]����t�TpP�iN����� ���Pq��Eb��EQ�o��*��?�3>��(�XT�|�� DW��*@�A>��vq�X����{h&|*
 �T�U��(������tyP4�xb>B�"�	�0�>�'�p�(>�h�-J��C�_� �)�D�W��GÂ��>�{D=D�ń �
�B2.� �A� @�RO�=�!>����x��PCS^T; Sh#�t��Q |�����mD�	��8 (pW"�>D6�t�TX�O@�|/�����pPM�� ��@OA�:ڞ |�_��]�T�AA,4�� @�G�PG⯣�Tء��F��OQD0A����|1O@G���:D4��/�s4�"�x p��|�j	D�B)�b�Ov ?��G��|�(@�FA,QH�Q@��A��M_w�k�HpH�@l�m� ����6�,���L�$$��F&���f�f�Am�������Ҵ&ݥ,�۰���)���Wn(�v%H|t��CI�t���㬄�ic7W0i���"8�J����ܲN��9���C:�;;x�v�A�I���;�1�GQk�4��fͨ8s2\������Ct�ӂΨ;a| l:t�!�����le��vK�>=Gg�������Q�	^�yB�m�ܕ(5hd�&�����@�<kMe�FwX^[sM��m��i�\����*լ)�m�=���2�^k��{i���O��6�l���`J���UW���q��\*�X���X@�p�$��h�.ΝC�V�L���6���XQ�FLu�T�3�Pd�eMiUUt+�O��n����:q�N���Z��5<�˖m%�u)��Wf��b%��=��p[�H6z�����C� U=n�U\�]���g�:��I�4���3ј��v'6�#��F}�a���N㒝�̫nE�㗞x]�^���և6˵�C���O�nn"��Ԕ�������$8m����	�5#�n�������e�f�&�*�VWd%L��-��rl����n�u�NU��j��&8����d��<��;c��6o63�ݶ�	
mX՛����a����ȸ��mn�ӻA�m�E� W�Nt&O+d�i�#;l��`.���Uڕi^��UƐ����`�U�k`��ɓq�*��0©��u��ݍ�gf��*n��gmu�;g&��%&YBM*�c�;<��#�b�E:Y�P��d�9z!�Dk���R�{n�q\=\=vI�`�f�$�z/(N�$6��GqG����m�k,PY��9n�m�YBM�ݮ.Ȭ����f� �,#bU]T�e�j�j�{`��=x��*��g��Tٞj@
V�p� �����d2M�R��� ffeɓ�J��T=EM�ҧLT���H �؜q*�~E�Aӂ>>���*|?;�{��]�L��SS��ql�i���v|�7G��9��M�M�t�ZGB�bȳ6���#�i��D��kvΐ�镊L�{v�[A�*�F��$MC+���.5W]����07u��v+���Ucq�ەn�.v��]v��s���s�i�!h��l�0�\�)���u�o$v2D�:�`ͼ��.f���XὬˣJ
m������V�T�Rjh��grrp���Ǟ<��_'�ؖ<6M���R~���4n�`�u��Wo��0'����Ws,���݁�sm_(�P�DB�Twu�h�ۚ�h�[���b�K32��07�0I1�ɱ���b�&�Mę#�4���y$�&�L'�_)&:`vl�Z�+2�n@cNf�ym���������s@�^�W�cr4)�c�	0q��yv����='�۬�֌�ks`�.,�
��sCRM�n�{����s@/�f��p�X������4�]6XO��2j!�4s���{�`�f��s@<��Ȕ��Ĥb̦��Lwf3ԗ}�:`{g�����b� �)1�"�4��hY0'vS���L��r��]!,X�V��09$t�ߪl�t����_z�������m'$Ƞ�B,��[2^}]����ܩy���/<��4Γ][=1+m��4�Ŋ93�=����w]� �z��n���-�a�qĘ�3@���ovc�GLM��ɲ��9�8��i�����<��h�a����(Q���1�O�B1�zA*��W���07�0:��JfRBW����1��#�&�t����ov���ܱ7!�A)3@����36Հgٮ�����Jb\�i~��"^펩0�ca�|��5��qѮ+���n��n�@�.(�hQ,sF~�s&I�L��ߝ0��`rH�ɲ�0;������0��hȤ� �z��n��뛚w]�Ӡ������i94$���)�[�0��`vZ�S䱸�M4
93@�������w�����;4�B�RZ9����f.}��y�|-�a�qĘ�)���� ���$���)��}�{���q�~���X�N�:חf[�vװ=:ղqֵ���ٹ�d���y�����9��
l$��� ��;��ڰ?nj��Q ����r>��_I�	8�(����GLM�遻�� ���kK�q5!�A)3@�������w�f��s@3��*k���2Ljd��vr��f09$t���N�ۭ�ݍ�a�K"�4��4�?{��y��yߺlܓ�}�f��_ � �P��#U%!T� ?T(�X�	 S@� 4F�!`� ��M)�',���!=V�j.����s�zyڝ���
��h�K˺����񮵃[��մ;M�G�s]��	�uɬ-�Ҹ)]�u�]ɻU%�V����7<)d���d0-su�c[��/��z�zN�FzJF8P[5U�78���]�6pJY�6&k�d~�����t��5-��)�j��c�J�.���Q�?V�#���q�H�;J졊������b�)8-!Ul/�;Z'&A�zcX���Z��<dy8v�����+tu���5PM''o�nh^���wu�����=�W���rF�h^e096S����'�0	����s@��K&�7Q��d����ovc�GLILM��UyY��*�$���:4��7����j���M��������VLHI�1D4�`rH�� 遻�� ����o�o�o�����p�ܳѻ���z�vn�[r7ipyz��aՊ�5��@���Y�[���\���Lݎ��f{�;�y� �V�5I�M�M�j�X����J�TIڪ$D�f�@j�G�`s��$���;�Kn�WH1^X�b̦�ٌI09$07��h�_�`�QdM�&�ؗ�}�`w��遻�� ���e�u>J�i��rh[M����{��_o�@<����atm�(�b�"��n�m�cA��]U���Š�3��:ɔ�x�L#n8�$&h������-�@��nh^�F�̒D��bR7V�f��IL�������`d�mX���Y0X��d�iɠ^�@�ߦ��)��~:�˾�[ �ߦ��q`�qbiƲFӒhYL]�l{�&�`߶�$�2<q�4^�z�����4-���R��91��F$�� ����Q��Ŷ[�tt��n��x�z��}��z�h�'�(����4��h[M���^�iб��"MED��v�s]�Jd���V�oU�gٮ�L��=K�eU9u54�%�����`r������/Y�_h��#MӚ���ՇDRQZ�z�~�v�s]��!$BP%
%*�v�Vn�+�)�n~q�$q�{�h���<���/z� �Q[1�Y#Pd&D�?�|�sٮ6��.n�y;9���\�/nm���g^B�(��#rx���ym74^�z����X'\X�q����@��}6o��1T�E Lɗﻭ�_o�@<�� �u�)"Nd���L[���f0I1�ɲ�0=��uF�9�G�w�f��Ձ�sU�	J!)��ڰ7Lf�R7R4HdM�&��s@�����uz�f��E!D*����V��cm'h�1�u�r�4lu�4m���ݢ��%7�ǭǵ����^���Z괹�#�f�q�T��f���@���o���2��X����:�8�h�y	V[Ůyf�+�%��U�9����@!vn�I�3o�v�|u	�����zx-«�i|sv�ˢR}a��=C8%�4��v��(8��؝3�d�l�o5�N��t��{�w�>"�G�WOjݗ\��&Ä�m�nz�ã�÷W\�Y��l���XӍ	��w����9wW��Y�ym��<�R��'M��fSV��ٌI096S�&ך��ds �H�����<��i�3�o+V��U���3��S�mS�-^c�#�$��ջ-�n���;��&�(��&�h[�s@���nO_ $��6GL��6[�j��uɕ�q De�,f&^��w-��xw:R����VαP7\����c�v[ ���6G^����W�0$�U��"NA,QǠ�Y������	$���	J��>ݵ`}���`};������h�qE�1�4����*:`uM��7vc�Ժ�%V�-	@�2����T�lwf07��hZJ�b��`��3@�^�`rI.���nwZ�7um����{����]�}����i�}����:�������'(�H0;:�jLXU�����3�f^_ ���l쎘J��Se�<E�U�by��(��;�w7�߿~ď{��L^��RK`v��J��j��m�[V`};�V}���k�C8�0)F8B&ouj�ȨU ��!�؄��� � 1���A!$H�
�="P �!���P� �0`F!��@�Ҁd!#���ؓ�ͩ���z׎ڐ7�L�{��!�F9���`Q^>)�d���V"��^���OOZe@�!�ߑ�A/�;�*:=J)��g����*',�w���m�?vCI$I̟��1��������I%m�}�=���ƒ�W{��~�s�%�]%�yK*�9�G1�I%��y��mW���I%�����[o��k�֭��T}��N��u&�*2�q����7@Pv�ί^�&1�� 	�v�hf::.��!�f���У_������i$�w����RJ/yմ�wjl�s�.�����Uj�� ���4�]��r��Ԁ~s2����.���֯~���-���w��������Ѽ��.�Z���?���{=�M$�*�����gz�^�y��IrHy�x�^�^�c&E!�LQ�Z�Iwvg8�R�v4�\��q%mU���D@_D��X���w�}��qjI/Y�_�G18܎LM��%]�ƒK~��|�IIq�i$��Si%�{?��f;qA�"z'6�,�a%]lgd+:�Z��=�ty��Z����<3�#�U�fX�I-��JK��I%.l�q$��Y�$�w�˞$�9��hr�Jˎ�I%.l�q$���i$���$����ǐC�M�Z�J����IK���I)$3�I).:M$��ĩ�Y ���#�Ē��f��V�O<^��z��4�^�O_�����^�%b��VM\��ݷ�kZ�zw9�m�uݗ��Z��]�u��j�]~���5�m�DO�A��v�+��&�rP�SQӽWg{�lv6l˹��m�6���s�"<��r�=u��1�P'�B��]uX�� �pt��tF|i�rj;>�q����خs9L{.�in�:�*���ۜ��ۙy;'@�k�)����^p�7��i\�n�րB����o�%!q;v�8˛-��/N�n9ݎ܍f,g�+��6�^���Z���F@���f��B�5ZH�5�<[q��e������[��^��]5=�Z������2L.��W��$��憒J\��Ē�GV�I)%L�%���2dS ��q�J�k�J)[I$��3�I)244�\�e1��'��1�#�Ē��ǩ$��,�Ē�]F������$��K�� �'�)&
Lz�I[r�<I+e�jI*��J�w���߻.xd�
B~����$��I)rK�J)[I$��g�$������İq��4��m[��ݬvLr)>�ʼv�vݡ���n�b�s٢s�uYAD(��ԒU�_�$�V�=I$�J���m%�g�I)S��V*�V�2���s������P�@@�Qˑ)�W��I/m��i$���{�[-z����1I�$����y�IZ���z������^#皶�]��7m����sK�Ga�L��J�w���m~x�U۬ԒK��<�$�v��C`�ǩ$��_�$�;u��Iu�g�$�+w�����y&7#B�&6ލ<ḹ��۶Ů-Wl�A��Ӳ�r�)n\H�I�zZ�����~;� l�3�I-R:��KnI|�IwJ�+v`�6(��)�$�[�y�Ir�q�I.v��%��f���߻.xd�b����YY��Ij�մ�[rK�k�S�|��iD�A0W7���z���|����*J׉\��AD!G1�I.v��%�#���[%L�KT����߶�C#�ё��r?<I.v�5$�ٙ��^��$���[I%�$�q$���|.Һ�4>�Ɂ�[2^}H��(���Շ'8{(���d�vz2b�+ڮ���T��Oz���Ij�մ�[rK�KnGcI%mڤ1,n7I�L��K���RIm�/�I-��$��*g9����[~�Ѧd	 ���9�RIW��?<I.v;^����������$�^�i$�z���7K\՚? ���s�}����ޝ�r�}�}�[��K $T0�hP�u3߼﷜�+L�	� �6(��)�$��r�<I/}/��_Im�z�Ēۑ��I~��k�x���-����Vz�l]2��z�ݭ����].��{h�n�Q�Y�?���w��ܷ^�2�7RK���V�Iv���KnGg��]�����%���6dcd�Q�z�K�6_9��UVf/_��ƒIz~���$��w����DW���4df4ۏ�K��ƒIoeL�KT�����͗�$�e��x�ă�$f��]��<�$�X��I.��|�Im��i$��ŘRUw�$��&I�%��ǩ$��:}~~��R��cI$���s�$W������W{��e�h����%-k#�)`ê�ٙ�ۉ�N�{p���Ӵ۠��P�:5�N q�7=+[rg�βp�T�������n5Մ��j��Z�*^6��<y��	;9p�n&[c���s��L9��8�z8�YL� ����S��n������Ӻe���hnl��ay��Q]���m�[��7�k���̦T�,�s�#BU�-���������q�|���AbP��l�:ֶ<p���6��v�|:��F ^-���_;w�r�l�閬�:�*��K�=��Ēۑ��I-쩟���P���? ��}>䛇��i�?��[�E�(��US
"��s�?ߦfv{�U�Iz�W�%���u�&�E$�H�I$���s�%�GV�Iv���KnGcI%�����4�$m52O<I.V�=I%ۛ/�I-��$��ʙ�$��IL�O�Ƅ(�=I%�_�$�;u�$�6S�8�Z�um$�~�����	|\��gg7o,kpd��R�a�����W�]d�-z��oOI�w"����~9����p�KT�����͗�$�e�y��xI0@����K��U���g�[G �A�`i}|�/�٭�m�ޯ�K���I%�]�C��qĞFE�%��ǩ$�w����f~m����I%{�>^x�^�^�c#���Ȧ�Iw�"�J^�cA���0�}U���~4i��z�1<�ɎF��@��[`{w��p�g�{r&��ԫi�֛��1���8�-���n�m�ݙ���뱌��L�BY�~xq|qˈ��O������097 ��nE�\A�[�{�W����m��������������������l�VA�#ޔ���ZWX+�tT�l�2s����j̅	+Qi	T%�{������Ł��I�p�:�;*ի�`��3g��$����܃|���=�����6�&b�=�nH0=�G��{����J�˻,I[Vx�{ݣp���-�6�M������Y<9յ'�>�>_
9%��soͷ������������W�~-S#�I�Ȥ4�m�31#��^���)�yzS@����F�r1+�`j��`w�Y&�;&0;��WX�oRL�@���M�қ�O>��ܘ�~sK D,0�Ȅ"HHH�F({
BC��@	 E���;����[�x����x���!�w��h�~Gu���z{rS@��iup�EI�;��R����.�+�A���m�u���s��n��LJd���	��� �����Ձ�5=9$�HnwZ�:7�髆ө�UUSvӹ�|�IuQ9���7;�4��4-U��m�R`��$z�e�`g۶��Q�TN�;'�����U"X���q'��8h�����sjÒ�Λ����*U���7�$s4��4U��yJh^�X�%�@�$�"E�ȥIjb�j� �D��+ �	d���X�N��F)"m
Мt��0C�I �H�!)�.���LD�lI	�1$	't8	*D�� H�I8�w1h}<���$��eF$BTt�A�Y!ĂE`�0Iz��vޞ���(�6HD�2���
i�c!��cQ���6	l�X�!�3���D��� "���"�"��$$"HH���<�!�8��1�Iń`B�e1`@���|WQ$� ��PӦm��$��(�24QJ1cF$"��t����������bJ~�$ ��dg
��˺�De��H�`a14!m�DLV�X@��A� 1��B3�"��EBA�� @� "E ĉ���I$A�$,M�9�D�!������D�ׁ�1�D=��k^�Z����!� �)BAm[M�q���%�m�mN���[QD��,��n����	�Bj%��8{b*�M���\wp{6z����������g�U��n]֋������D>]�<VY�
J�4�l��������Ç��h����(�"��%v�i�d� ���� Ca�Z��hF����j�J��W)b/v�W��;krn��v�zP6�i�֝��ς��v��خ������h�7`�E��;Z�lcg`6r�
ݧ-�J6s��lB`���j *q�>ۑ{�tKWW*�
ո:'������['i���K�U)(qT@'=��ZU�P:u��\&P�$�.��9Ty��,�v���b�%�K �y�םh�MO\���8�E0x� &�cn;Sʎ^w>ڱM���A�6�(��jT7Z45{+�T�'[/:ᔝ��l�ёٵ���*�G+ʪԫ9����+���g�Ȣ��$�.d���v��S!r�R��]�_#��웠Maϋ�8���I��ݓ$9�V�=7h1ˢu8^�݂�8�-T�,D����63�#Q����mf#���Tl^Nno �m�LXm��&�uЖRC�R�t���Ӳ&��Q���k���cv������\�tJ��-�:@�Ӎ6���IT�A*N�]�fB����Mu]+��e5�X%W�m�%*����o$H�m5��5��*�v�ZWn{��Y��Ek[l�`�;K*n: UVՁ�'U�/<R&��&�[UV�+ ���;]PH�\XP-Jϓ�~*�4'SXy]vv�i{@Fv;v����yT����m�^\tC�޼�/BD���Θv�3�c�>l�B˷&6��-���A���,�`��M����M�B�u��ٕj�ݖ1����6���m��7i]��0 �e� ��ZW�a�Oc3Ё7I9%�U��b���l������3F�k2\�C�D�Ϟ���	��z��z�tpv�!�X��񻬙�fB�3!e�M��7��E�s������\q7�l��'I��A3]!e%�cr�ӯdC�h; R�PW�'�א����m��Ud�'wp\�m! ��n��tWgs�2��F���<h�G��јA������n慺��|��7σ�bب��`8O[Y�(� &�6���g�#ԙ:�1*;a��-��1I�{Cnmw<���]1e����{����z:��Q���������m�>��f�糷-��"��{smPa5���cY�8�'���=�R�{n��^���Eu�&�5#�H��/K�(Jd��`����w6�ё�4ƛrH�9��;�w4�Y���r{z���%�C�T�+n�i2jH�s4�~���z^R�{n�ߺ�����ё��nM�z��)M�Қ{��9U�7���n�4�dѫv]r�=��c�Mӷ��t��I�WLʱ������rb���$z^R���4�Y�r���<�U"X���̳D��Y7$�Ͼٻ�V	��, �"�E4�@!���ԫ�����ڰ3r^�В�2{���DjI������h���yJh��UMȜȲ7$q���T�l��쎘z��K�{����4�6F�x)�ה���۹����z��L�ؚ����+��ɢ2�3+Ӻ���,�����ml<��a��~����x����JC�/}��\�vӹ��%侠�t���g��i<�rF�������9}~z����Ϸm_�Ttw����iԉЪ���g��3r^�|��	$L_G�����`����ͥqTږ��R��DG�W{����޵`�������`}�O��bƣrD<��@�zd �~/u� _��@��S@��F�yc�Nʰ���NӶɐ�g�|�R�m�N�����Ʌ�W�|�?2y�i�������~�wf06j�{︃�<��󬼙D�4��@/�f���~�|hu�s@/u��G����P�k#R1�&�����3smY�'n���`~�������R+������hI������1�P8��"@3�Oߕ����/}�\{O ���(�0	�1�I�5dlt�ꊶ��l;��&g�,�ΐ�v�:�w xq�w���{\��L%n��Y9F��1��VA�&�Ln�`I�J�[j�@�R�M�7%�|�N��Z��M ���<�U"X�q�"
D�[�s@/u�oY�u�)�z���d#RH��d�f�^�4޳@��S@����pqI2<i���I^c �f0=��O� ���0	�f� �D�!Ԣ�])3Hw�;骺�<f�%�I�mv�p��,��6si�N�����]b�K��Iծ��A�3��-��e�zFuܖT#u�+��K�\�T�G�n�(+�p"�fGg3�8;d� ��H�V��S�+ם�8���Kn�+��g!׻PQg�t�l��|�ĺd��6+���u�9������H��'=���8��ss���555���S&Y�&~U���{���Ɔc���Q�2�=V��#�k�;����uk�{<����{V�a�;x0Α9u�4�o �d�,��V������{p*�a5 �H��-빿~���{��06j�09���o.���4�� ��h^�@��S@��s@��Q����"��rh]��٫ �ٱ� ��It�W��O�O��M�)M�]� ��h^�@=��&�$�m���+n3v��j�����[��^���U{7f�l�����j7!1�N��4�Y�޳@��S@�{΍c#JH��r) ��w�/Ȉ��R��YHV=v����7�z_B��L��[)�MTӒF�rh�_����)�w�)��f���h��4�6dr"9&���)�N�A�n��K���e^C(˦��$R{Қي����M��S@��U�f���?�E�lݱ��q�d�Ղ������I�qun�kl�x'Q4�	�j) ��4��hyJhޔ�;:�o)�y6��@7��}	D%2ol�,�|X�k�<����ɎO�L`��hyJh��1}_meU�Z$�c ���"����$Ƀ�8hޔ��f�_s]�BP�{f��2sk��C�t�H���^�4��hyJhޔ��}�w����>��ӫ�m��3us�˷m�F�]����C�\��Pqٲ[�#�j+�"rII���~�^R���4�Y�{��+��5����I�u�`N�A�Mٌwf09��&��q5�8�4�Jh�@/�f�ה���\J�bi��4��Q=���7�������QiD$�c�����?>~S@�/{R4��,m7��'vcf��wrn�`z�������6:ѹ�vש&��q��t;��ð�����3��/^\�n��Y��z,���܃ ����`yl�D�cQHI��p�/�)��f�yz���S@�{]���	�Sr�`���?nk���ID��K�@�gƁ��.��ı�$����ɳز����`w��F��XّȈ�{T��}�M ��v�f�$��P�涩j��
n��5��J$ۂ�\Y�a�g�^ts�\�׹s��܄�-����:M���Kb��Ԓ��.�]�:
�����v?����Y�X�����d+�m&�N�f�-˛d��Ӵp-Ѱ�����[�ݗ�n��q����GO"�:���l��g�'sIմ٬�l/ ��5˲�yݍc����tH��h�9ŞK��=Yn��~�ng�va�Y�;B7�D�1����\�[����cnz�]����v�v�F�����D�D�S��) ��S@;�� ���{T���\J�bi��4�Y� �ٌwf07�d��`L�=�H�#ȱ�ܚ}�4��M�Қ��h[^�&I�L2c�3ز	��0ݘ��R^���=���,XԎ)2`�N��4wf0M���Ő`z�a�{��gV�:���=�gQnǎ9�N�cQ��00��z�8�>q���W�O3Ut��+6���&�`mvd��0$�O"�&��F�rh���˗���3���x:��0$܃ ٳ��Qٖ�U�Yy�Y���H遽܃?��F�{�_���`r��J<Q�~�2I�{��&0M���W�eOr���/<Y�D�5��y���ٟ>�? ����Қ~�,�@K�S!:����Ԛ��ݻ<���b��녮�<�en���{�3cf�#J�X�nO �u���vڰ3sm��}@g{�����hUI�ra�
H�{:�hޔ�:٠U�W�~H���D�1H⑀<rf�ٯ� ����Y�DD[V�~��&�c5�R���NAm�@p8"��!�u�!��5}6I��8�"hӨP�nɥu544A��P֒8��R�##<�G��M�<Q-����(�hc���G8�-���� ��U㜂��'��` �O"�y��@@�胈����U*!�}_���*p�*�>:뜾}�nI�O���=^�_�rI27�$s4>K��F^��vD遳c�; R��e
'$����+��u���x������<�P���\�k�u�5;���ѧ����W�[#v'cr�u��J¦K�����Q7���'#��|�4�w4��h���v+�4����x���0����-�ݑ:`y�Įő�N8�s4��h���޷L��k��f,3�.�Uڻ�`l���ݑ:`l��>[nנ[n�1���d���E�{֭�͎��%�6^���v���G���&b�v�;ݣ껟[����n�c�z֊��^D뛥��LPq�TS��~m���~�`j�������ȝ0:��_^\�L�������޲��j��=�w4=�*�ܘ6��H$��=ِ`wdN��07�"`s颎�cfG"�p��u���h~�s@�]�@�����`r�cQ�#&2d�L�>��VBK1�O�3y�`}��j���Z(ej��t�Q5�GAV�!�"@�J(��
@@M�R���� �_��5������ne��7y7o�r6��!�c��Tr��]�m���95�l<�I�o<����}� q���sõK���p��tj�uK��b�+.�mch�kr�oGi�d�6��g��2]��Ԧ�sՎ�!�����^�x��6$7��bVEx ����۟��ś��ù�Q�.�[g�N=�#M.��t�j���VQ�J��pj{����w=ޭ������z{s��t���&+��E;l(zس�#��[*t�GMV��rRE��N8�#s4_�h���=�s@����;=:�"��B<���0;� ���#obt�����܉�zݘcx���'�4{���=��Vz%�UY��M�ޮ���^�s*SRH�`�3@��s@��j�:��C�]��y�/��c_�rI27�s4v�LT�O.��N�6:`��sߧZk�\X��'�φ7=�۰>��f�糷9��ki�nm�!;a벋UvW��OL���؝06lu�����Ɂ�慨�(�29&�{z�͙dE���u	%	z�����X��7�{p*zcQ�R~x�S4�w4v�L�}IOL���{��M���X���4���s��~ �>4;��/��ׯ��}�_��BD�E�&��7��0;$N��09�"`n�)�?c��4�ôDvP�j�+�:�ܻ��i�㝺����L��-���͚�מn�/�o�����t��܋��[=lo�� �9�� �S4=빠x�K`qwe�;$N���<��U��.��R(�mXN�U����VDBJE	! � `�B*!b$��R�)D8����5�r��3��Xf �Or`�nI&$��=^�z��4vGL=�����7�Ay�X]�م�,Yyl	5d���r��O[ �Ɍ7���m��~DV�\���U���a���wTaB6q��ǯh]�m�uY]�=h�b�Ww�0`wv:`un�`�3���)�[�%�ő�N8�"s4Wu{�$��0=�Y����4�ًĠG�diI4ζh{T��%�������߷m�U&�6��̶�<�yVo���{�j�3��a�+�-νv[!�c���0��@���hU)��p���;A�:|L�*�fc\Xiu������;P�qƹK��s�vZ}�U9�4����ϗ˓Ԥ�^�J�Ͷ����0l���b�0;ݎ���<&��$�����G���s@�nh{l߿~ċ��/���Ěs�/:`w�0��96cn��6)q9�~�W��f��z�&�a���v'ၳԗ��"��yyj�/)�Ų[�|����س��=�f�Q�_"�y'x}>wѵ[X� �k��N.3{/I�e}p۶n״��4���8ڎ�$t�9�R)Y�vÅ���	
s��T��x����.��]�䄘�N7����<�8�Sg�i]ՠ��4�5�ʗmSմ��9��NYЇ���ϗZ�:xzu6_QǴ�^�@ݞP�v���h�	`�װ]gv+�)�@ַZ�V'L�L��W����b�x�v^����]���{���'aݦL��zz��ڂ��lj��-�R��8��R',����g{�7�P�g7Du��������udݎ�[%�7��hSE2�BqJe�v�^��J�BUFo��'����wВ��2�������0N)��|h.��������<^������7��#,9BIOս�`�����K��З�g�}���Ɓ�%�&&�rIr= ���;� ��̃�d��ZUŰ��t�E:�bz��< ��\�4્q]��]�=�۴j;��{��<��!e��\J��p�Y�͙��=��}����>�>�6)qHhu�ހ}1���ޤ�s�ܒy�f��ڥ7����-��IO�N5�$�{wf09أ�6d��
##��M�3�~����V�ץ�%3�������sN�Jp�̶��l�З������`�Y�Ա7�9&H'�LlpM�n]n�:ǒ��=���v������?����i�1�9�2@�L�o��@;�f�{�f��]���f5�F���,s0`�1�������y��2�g����KrLM��$���4'<���s�XDXD��T�ןf}6�����u�&�Ć���?)�:{�>�|X}��<�Q;������lǸ�8��C@��M�3��g $��;A�ϻ���OB.�T�W�%��a���A�@=�k�pp@�-�p͒�%��އ���@����ߛm�����n��;A��2�-���2�:NS��݀ff���J����O�@;�f����$qL�����v,��d�H��c �{}FV�T�����*���:"~�,s��fk�tD(A��H����"#����'ʡ�٫���}~��5L�M��-��X}��B^���?�����4��=\�.����52I�6��N��h����/w.t�z]�����ϣ�f�n\��jd���)$�9&�^�4=��h�)���}4����(�ǎ&�C���l�������;}�`����B�;uqTQj�d�UNi���{&3�|��=�0&�JS̩��u.��l��%	L�w; ��v�vՇ��u�`}��V9M����r����&��;t�����H.��`H�������� ������"4�����y�;=�G� p��^*p�LX� �	ff���
>�SJ� D
m���װ�f��,X0<��y���GG��4"1Z��T��D"E��<G"���1H$aT*�O5��@uP@�  ��ꮢ�Bc"�8�5�8�� E�f�H���U�a�$QҦ����������lG�!��U4�v�XP�R0_��֮kZ=� q� �)BAm[M�p  ��Nۂ�^��m[i �C��mXōU��%T�P=YY�^�՜�Ǔ��$�
��n�n7Xv��k�<�)ru�6� )�t�m�;i���̃u���N2.5���`�W�7L��*:m��{g`$��W���j����=l��e�5F���t��5�&���:YP��k�L^��M�a��.9�Gf��v+�<����m��'�<�n:��WX-�W�΄�ɘ�8��lv�`:!+-�<��7nʰ�Z�c��J�e��
ZP
Nؚ�� 9��R��9���մ�UMmO,��ٴ�``��[EPli�ё���mR���Pq���b���C�[Iӕ�6:씻hx�ZZ�yGm<ب
�v����Pkm'�FAֆs�8ݟ0In�t��������L� ���������n+bU� ���ڦ�T����	��A1ll���ͪ�Ê94�\�1�.
q��'�&�(�R�.6C͛�8�Re:S-rg�������aײ!���'#��6ō�������u�3LW�%.ɥ�̫�Y�܋lX��N��hg1�<��㗞���z���ԡX�ڨ)��yYY�A��]d�q"�ٞu�μi�%���Њ1��9L�<�m�[���\�q�$e(
5m%�*�둭��m��e3���r�y[U��ݩ$<+#��9b����A�u^v[���v��N�`��]�V��§U��-*�e�UeZ�@vT���UVBU:���'��������������<�,��l�Jݳ�$�ِ�s��	�Y	�dfVwm��;a�[;*��ҭJ[\�(�&�����b�a���@F{j g�xꃦR���\���Z��vyY]��
��Z�M�*�R�d���$jT6���ȪҭA�
�����,kCl�PS�����V��[�l�Ɲd�]�]�ۜ,���I�`,�p�^�v������4����w����U��p��"	�1����S��������Èx��OA^g�&�55�t����rP:fn�<n��qE���$�;���m�!��s6ֻۗ'%�y��9�Mpv�I�\D�XN�&�jB�+�L��d��Rr�H��(�l���	���:ŧjS�.ܜpn�t$��qwP�ۭ�s���8]l'0��z��\,��;o:X5]�Py��b존�tL��ܐ˴�쏮�ێq�C�*�i�v�[kL��^bƶn��d��~e����9 u΂�㩎���p7���x8v9�h2F���"D�M<Y?LB�p�/�4�������~����1�8�Ȇx�)�;2{&0	�1���h+�c_�rG"ll���4��h{U��;�)�{xkrLQ�ff%y���%���w�Θِa��@�����k8��4��<��j�ϵ�`���5�IB�Hٞ�w�z��hmcs���uݭh��l��`��E�ݴ�XF8�v��u�:欱�Xn�؛���7�c �ٌv(遻))[#M��F���7���g��~�@�`4��X�]�3iȖ%�by�oxm9ı,O���6���MT�K߿~ֹ&L��1�K336��bX�%��fӑ,K������r%�bX�{��m9ı,K���m9ı,O=��ɒ�Kf�C-����K��D�����ӑ,K��߷�m9ı,K���m9ı,K߾�m9ı,O5>��5rk��L�Zˬ6��bX�'}��6��bX�:���6�D�,K�ﻛND�,K�{{�iȖ%�b_���w%�CY��Bf�fQ����N׎��:m�v�k�%���<�<v��wYk��TP�u[��{��7���������"X�%�}��ͧ"X�%�罽���Ț�bX����M�"X�%�����㫉������{��7����߻�ND�,K��{�iȖ%�b}�wٴ�Kı/}�si�6%�b|����j�5�Y�j�3iȖ%�by߯xm9ı,O���6��c��:�Ԣ�@u�����y�6��bX�%���ͧ"X�%�߾;5���Y�5��ֳ.��r%�g��߿s��r%�bX��߿fӑ,Kľ���ӑ,K��^��r%�bX�}���j���[��{��7�������iȖ%�`�{�siȖ%�by߯xm9ı,O���6��bX�'��O�GV�/�r�N:��H�m͍�Y9�'�C	�i��Tx�[$B�<r��fӑ,Kľ���ӑ,K��^��r%�bX�{��myı,K�{��r%�bX�{�y�%�,�њ!��36��bX�'����ӑlK����iȖ%�b^���ӑ,KĹ���~!zL*!I(��(�2���4k2��"X�%�߿o��r%�bX������KʰuQ/߻�6��bX�'��p�r%�bX�k�٪jffe̹��L̛ND�,K���6��bX�%��w6��bX�'����ӑ,K1�b?��!��C��N���ӑ,K���d��53��e���u��ND�,K�߻�ND�,K��{�iȖ%�b}�wٴ�Kı/}�siȖ%�b~U?��,�u��cֳx�ku�$�6�<�����.�L�^�k���^�\��~w{痋�Ny���|�7�ı,Ov���r%�bX�{��m9ı,K�{��r%�bX�����r%�bX��};���32]e�f\��iȖ%�b}�wٴ�? ��MD�K�����r%�bX��~ͧ"X�%��~���r%�bX�����f[�S.�W5���6��bX�%��m9ı,K��m9�[��]�m9ı,O}��6��bX�'����ٙr��R��ͧ"X�%�}��ͧ"X�%�罻��r%�bX����m9İ�/�����Kı<���&K�Y5�)-�fm9ı,O;��fӑ,K����iȖ%�b^���ӑ,Kľ���ӑ,KĂ�<�DAP���h�I�GY�Y�d��q/X��f����hqE�m��F1;�����+tguY� �nt�q:NY�Z���m՝�]�&�;Iݶ����Y�Q�ۄҬA�@�%i��|;V����nn�Q�	s���C��{`��n��N�j������q���ֳt���)�N�MI�;m6�����V�Hz��݋۷n��È�K&�9l�$r������W�￝��������+<Ks�.��Bm��q��>��-۬u�m>�u��"u��ny65JL�Lɖ5�s&�Ȗ%�b}���ӑ,KĽ��ͧ"X�%�}��͇�b)�MD�,Ov���r%�w��￷��2y�fԺo����7��,K�{��r�:���%��߳iȖ%�b~���ӑ,K�����NC��7���{����_�W1UW��bX�%���6��bX�'}�o�iȖ4X�'�����H���mI�=}��][�]Kn�7��N���fӑ,K�����ND�,K���6��bX�%��w6��bX�'��N���Md�fe�2m9ı,O��y��Kİ��{�ND�,K�߻�ND�,K�|o�iȖ%�g�����[MEÅ��;7a��		Nt����l�:_WN�M��E��^��.t2K�5�ND�,K���6��bX�%��w6��bX�'~��f��)Ț�bX����m9ı,O~�n��3.S0�Y����Kı/�����6��&�"X�ύ�m9ı,O=�xm9ı,K�{��r+bX�'���d2�Lє����r%�bX���}�ND�,K�{�ND�,K���6��bX�%��w6��bX�'��w�T�fY�d����iȖ%�X�{���r%�bX������Kı/�����Kı;���6��bX�����=�ުY�.��{�7���{�K�{��r%�bX�����r%�bX���}�ND�,K�{�ND�,x�㿻�o��復�͋O?�$Χn{5�͝��]���y���-��;\V�Vv湛Ys32�fgȖ%�b_�w�m9ı,O{�ͧ"X�%�����"X�%�~��ͧ"X�%�����53WTֲ�̳WY�ND�,K��o�i�R:���'~���ӑ,|Xj&�^���m9ı,K���ͧ"~��������
�*t�`�ܴ�p���$+�~���Kı/�����K��z��ө��ND�ߟ�iȖ%�by�M��ND�,K�[ә��u�Y���\̛ND�,��{�ND�,K�߻�ND�,K��o�iȖ%��Rj'~���iȖ%�b{�mܟ�e�`fK336��bX�%��w6��bX�'���fӑ,K�����ӑ,KĿ{��ӑ,K���%�֯p�v�q��d��s�o8�����e��bö�d�tl,�u�����瀫��%�bX���}�ND�,K�{�ND�,K��{�D�,K�߻�ND�,K�O�٪Y3,�2CE�3&ӑ,K�����Ӑ� �Q5Ľ����r%�bX�����ND�,K��o�iȟ�&�j%���ۣ��\�ə���L�ND�,K��߳iȖ%�b_{�siȖ%�b{ߍ�m9ı,O���6��bX�'��N�s5s.k5�33-�fm9ı�߻�ND�,K��o�iȖ%�b}�wٴ�K��C�G�✑7���m9ı,N��sS5uMk)��5u���Kı=���6��bX��~���i�Kı/~��6��bX�%��w6��w���{�w�߯�Em���tu�i�˵��i�rhN�ݝ�O^zD��wX��S�����Y)�K�n�iȖ%�b}�wٴ�Kı/�����Kı/����S�,K�����r%�bX��ioNfj��L���\̛ND�,K��{�ND�,K�w��iȖ%�b{ߍ�m9ı,O���6���X����b{�m�?\��j9�R��ͧ"X�%���w����bX�'���fӑ,5Q;����ND�,K��߳iȖ%�by���.d��$4Ks5��K���o�iȖ%�b}�wٴ�Kı/�����K���MD�?w����bX�'����j�L�3&Xh��d�r%�bX�{��m9ı,�{��ӑ,K��]���r%�bX���}�ND�,K���_��|��Lt����Fv�;YON��L;��F���坟j�pd���wh5���/n���Ia5���k�{Wnڔ�#��{]׎Gcg3�c���3�Z��G>(�u��.Ssġ\`��չ�lu�3�(p����-*�ۍ�8ڀ��	��6x�VP#\[6��h3��=�`���(X�&:۳/i��T*�3��ɚ�\��~�!�U5�M�th�55�dnz�x.�>N�ت��v���n��X���N��]s)Cӝ�Z��U�}���"X�%���ͧ"X�%���u��Kı=���6
�%�bX�{��m9����ow���n���I3P5|�r%�bX��w[ND�,K��o�iȖ%�b}�wٴ�Kı/�����Dı>>���j��SY�3Z��ӑ,K�����r%�bX�{��m9ı,�]����yı,O������Kı<>����e�$2�[�2m9ı,O���6��bX�%���6��bX�'����ӑ,K[��o�iȖ%�bw���9���Y2�kYs2m9ı,K���m9ı,Ou߻��"X�%��~7ٴ�Kı>����r%�bX��>�%�7�L���l��m�+n�۸���N�:{�qY��f.����ws�o�>�SO�`}��D�,K�w��iȖ%�b{ߍ�m9ı,O���6�@�D�KĽ����r%�bX����2eɖ��2CD�3[ND�,K��o�i�p
���O�"4(a�8�D�KϷ�ͧ"X�%�}��ͧ"X�%��v�\/�/T¢������ ܍6
��k�"X�%�߿o��r%�bX��{��r%�bX��w[ND�,K��w�ӑ,K�������33W5���iȖ%�b_��siȖ%�b{���m9ı,O{��ND�,�{�ͧ"X�%��~!�NY���]\�̷Y���Kı=�~�bX��R?~���i�Kı;����ND�,K��{�ND�,K����cDv�M�E��%K$�5����p"G]�{i�n��l[�|�����'U����m9ı,O{��ND�,K�{�ͧ"X�%����u��Kı=�{�m9ı,O�I;ٮf�f��2�JfND�,K﻾ͧ!�!���bw_~���"X�%���~���"X�%��~;�iȖ%�bw�Rޜ��Ӭ�s5���6��bX�'����ӑ,K��]�u��K.�� u�9�TٱB	�(� �S~�Ͳ�衠҄<5�Q��bk�GO���pM� H�f���M ��@Y�(&�*�Ą tͫ����# E&�!� CD�A檾�b@�Q�٬ ���,դ���jP��%V�xR��(�Z�R�-���@q@��H�@	NO�G���T�y} ����TSh(���S�� iC�_Ƣ{~��ӑ,K����fӑ,K�����'nauc�[���r%�g� �'����m9ı,O��?p�r%�bX�}��m9ı,O��{��"X�%��w�I�rۚ&I�%��m9ı,O}���"X�%��`��~�O"X�%��}�����bX�'��{��"X�%�~>��f�]fgN��ȕ�ћ۫v�yܻ�[��s����Xp�5��n'+��N4[Vמ7|�~oq��%����fӑ,K��^���r%�bX���'"X�%�｝��K=�����ߣ�'��Rt�������K��^���r%�bX���bX�'��w�ӑ,K����iȁ�������۾�~T��V~{�7�ı,Ou��[ND�,K�{;�iȖ%�b}�wٴ�Kı>׽��oq�߽�����H�V�JV~{�2X�X����ND�,K﻾ͧ"X�%����u��K���<��P!w�>���{�.���ӑ,K���'{5��k5�HeԶfND�,K���6��bX�'����ӑ,KĽ��ͧ"X�%�｝��Kı?( |�;��חKq��-��C%�H.6Ŏ:.ڬv��7������	Y����8>w�G͢�*�=���7���'u����r%�bX���siȖ%�b{�gxm9ı,N����r%�bX������2�H�F����"X�%�{�{�NARı,O}���"X�%�߻�ͧ"X�%����u��Kı<���̘L&h�C.�6��bX�'��w�ӑ,K����fӑ,��^���r%�bX��w���Kı<������2�0�E�Ma��Kı;�wٴ�Kı>׽�bX�%���m9İE�{;�~���7���{������s��I��ӑ,KĿ{��ӑ,K���G_���m<�bX�'�~��m9ı,N���m9ı,O�|?C�8~�33�C�A����I�y��{��5�J[�n�Wd�ی�# �7hU��uۅ��Vl���ݪ;uN�4D���tt�+D�7t�q��f�v;p1�EX�bi�;�p�q��6�F�VdJ�t�{.o;���c]���D��M�H�u�v�m���[�"z��]2���&v�!�q��H8��4�X��5���ƌ�f��|�l��7m�����2\�帪�rF�����3mj��cv����0����`�.����{�ӚO�ˮ�P���Ou��Ŀ���6��bX�'����ӑ,K����fӑ,KĿ{��ӑ,K���������fd5��nk3iȖ%�b{�gxm9ı,N���m?>T�KĽ����r%�bX��~ͧ"~ 	���bt����f�\��˖ۘm9ı,O����iȖ%�b_��siȖ?����w���r%�bX�~���ӑ,K���Rޜ��Ӭ�s5���6��bX��~��ͧ"X�%�{�{�ND�,K��w�ӑ,K����fӑ,K��ߥܝ��jGZ0����ND�,K���6��bX� �����"X�%�߻�ͧ"X�%�~��ͧ"X�%��~*�1�+��7:0�s���s���h|dy8�Iv���Ht����[����fӑ,K�����Kı;�wٴ�Kı/������"j%�b_���6��bX�'����j�e�0�0̛ND�,K�w}�NB�A�i�; ���%����ND�,K��{�ND�,K�{7ٴ�Kı;�����j��ffCW&fM�"X�%�~��ͧ"X�%�{�{�ND�T,K�{7ٴ�Kı;�wٴ�K7�������P?*XpӪ�����7�Ľ��ͧ"X�%�｛��r%�bX�����r%�`#b}�{�m97���{�{������:�̐M|�~d�,K�{7ٴ�Kı;�wٴ�Kı>׽�bX�%���m9ı,O�	�)��1�i�f��.`���Lp]�������m�F�m��Ovś5r�Ԇ\��d�r%�bX�����r%�bX�k��[ND�,K���6Ȗ%�b{�f�6��bX�'�����f��d��j��ɴ�Kı>׽�bX�%���m9ı,O}��fӑ,K����fӑı,O}�]��2�A�I�.fkiȖ%�b^���ӑ,K�����m9�݃�F�n'y��m9ı,N��bX�'���9�$�3D�5%�Y�ND�,@�;���6��bX�'~��6��bX�'u�{��"X��������6��bX�'���~���rL0�Fkɴ�Kı;�wٴ�Kı;�{�m9ı,K߻��r%�bX���}�ND�,K�{�I��u��kS0��/i�=���ѼN�6��+v3���Gv�ߜ|�:�}۾%��_2�PO�ߤ�Y�ŉ����m9ı,K߻��r%�bX���}�ND�,K�w}�ND�,���������RÆ�������{��%���m9�,K�|o�iȖ%�bw��iȖ%�b^���ӑ?����bt�K����532�\�5���Kı?w��M�"X�%�߻�ͧ"X��b^���ӑ,KĽ�{�ND�,K�I:w\̹r�.d�3&ӑ,K��{�ͧ"X�%�{�{�ND�,K���m9İ"�ß�D�;����b~����ND�,K�R��2��rfk5r��r%�bX����ӑ,K�[�����Kı;���6��bX�'{���r%�b�������q+�\��b��N�}Y�����V�q�Y�1q�	���F���Y��Kı/{��ӑ,K�����r%�bX��{�a�"yQ,K�߿siȖ%�b{�q�35e�$ԖkY�ND�,K�|o�iȖ%�bw���"X�%��{�m9ı,K�{��r$�PPI����T�jM)��X��H'���͉ �'�}�&��'藾���r%�bX���}�ND�,K��ܧrjd�Lֱ�ɚ�iȖ%�bw߻ͧ"X�%�{��ͧ"X�%��~7ٴ�K�K���ND�,K߾�ֵ%�e��&�55u�ND�,K�ﻛND�,K��o�iȖ%�bw���ӑ,K��w�ND�,K|Q>�����SZ�Y���ĥ-�]ӧv͒��k�y�����%v�E��н���Lxtדv��ܴ��@�Km�K+!JK�,�([b�ܽ��z�g�[����9wOW;����E���=@l�ζk��s�w��r�-�u��n�}�&lAp�&ݏ�� ���;������.��	��r�m��)���Eg!m�p��m�ڗ ��:Nl������I���w�7"g������ӭ�O�ݛ���r�u��J; ]:�=��w�r�|t��nH�k������d����r%�bX�����Kı/}����Kı/{��ӑ,K����;�f\�u!�2]�iȖ%�bw���"X�%�{�{�ND�,K���m9ı,N��ͧ %�bX������\�nk.[�5�ӑ,KĽ��ͧ"X�%�{��6��c���j'�����Kı?~���ӑ,K��^����5#tL-���ND�,��DMD��߿fӑ,K��ޛ�6��bX�'{��m9ı,K�{��r%�bX�{�x��I��rMIf����Kı;���6��bX�'{���r%�bX������Kı/{������$-��UJ������+��7;>�\�m�L	��l�����.�Ȫ�MV�~�5�ܻ�,˓�L��iȖ%�bw��fӑ,KĽ��ͧ"X�%�{��6��bX�'~��fӑ,K��߷)��2f�c��3&ӑ,KĽ��ͧ!� 4 șĽ�y�ND�,K��o�iȖ%�bw���"X�%���v]j���fL5�����ND�,K�ﻛND�,K�|o�iȖ?��������ӑ,K�S�����B�����uO~�Ԕ6�S�5u��ND�,���O����iȖ%�b~���m9ı,K�{��r%�bX�����r%�bX��|N��3.\֡�2]�iȖ%�bw߻�iȖ%�a�`(��߿f�Ȗ%�b_�w�m9ı,N��ͧ"X�<ow��h?~�`���fN�'LF��Y�m��wF�-۱�s�����mw\.�຤|�˖��ɴ�Kı/}�siȖ%�b^��siȖ%�bw��m9ı,N���6��bX�'����ֻ�.���33iȖ%�b^��si� �bX���}�ND�,K���ͧ"X�%�{�{�ND�,K�~�ɬ�\�2MIfffӑ,K�����r%�bX����m9ǅW��F(� �U��*���,�.GH!��*�CB�P��iu����~�"^}�ٴ�Kı/~��m9ı,O5���B̹35.�3ɴ�K��@�O߿s��r%�bX��߿fӑ,KĽ�{�ND�,K�|o�iȖ%�bt�۔�k4��c��3&ӑ,KĽ��ͧ"X�%��Q �߿~ͧ�,K��ޛ�6��bX�'{��m9ı,H��p~�羔U�,Z]Ȏ��n{/�\��nc���Hێ�ݞ��p+.�K���,��r%�bX���siȖ%�bw��m9ı,N���� �Ȗ%�b^���ӑ,K��������532�\��fӑ,K�����r%�bX��wٴ�Kı/}�siȖ%�b^��ͧ"~U5����k\���\r�K�Xm9ı,O߿o��r%�bX������KD,K���m9ı,N���ND�,KޟRޜ̚ѓ33-˙�iȖ%�bw^���r%�bX���siȖ%�bw���r%�`O�C�'�*>��DD����M�"X�%��}n���ctL)�̻ND�,K���m9ı,O{��ND�,K���6��bX�'��{v��bX�'~�/εu�2e�0�Y2�om�L�����n\����X��A�Y�Kų���{�7���%��~;�iȖ%�bw��fӑ,K����n�S�,KĽ�{�ND�,K�v��Գ.Lɫ����iȖ%�bw��fӑ,K����nӑ,KĽ�{�ND�,K��o�iȨؖ%�ӿnS]̮a�k\��6��bX�'��{v��bX�%�{��r%�bX���}�ND�,K���7����{��7�������.��\�|ND�,�Q5���ٴ�Kı>���ӑ,K��{�ͧ"X�
X�{���r%�bX�|^�S5uL̆�W-����Kı=���6��bX�'{��m9ı,O����9ı,K�����Kı0�7�O��=HO|n��ɰC����Ё�dE��
���#X��� �@
� C��s��N)�*&eeQ"UJ(zf�˨D�I�C )0�����U�h� %y�yI�d�L4a�D�[��d��O}JmG��`���(�M���mp�������o�ۖ�8pջ($$[M�  ���m/Z-��HH)�M�@��$�I�U���5���-UK�l����y���A�kRctݚ��[��ڨ�n��cY���.��K��иop..m$el�ԭ�#]fzV�c�V�kfԼ��T��t��곳��(�����\33Rq567</Ev��S�]�Ϫк��ŏ:qΧ���T[�iǖ7�R���!=gP39�mz�KNr1��KU��YJϚ������r�@�m�s�ͱ�����4��k UlKW��uwn݃e��@qf�;,Yٲڶ���F�=C�3-Ip 6�t[tݵ�K++U���٥�vyx.�W���ijv
�6�UJ�Y��uc�E��f��7^�lg)݃J�� �Z�Z�wY�UJ�r�8VV�L����N��8a�R��	���!<m=bEi�-#��s�՟SX��nU�:닭�RxW]��Xظ��ef2�>��p�g�l�ݲ[ؔxz.Vo�M�[�[��L��H�]� t�m�l:�9�_�����r��n׫�;ZCc��'�Lk<�P��y2�fJ�i%���LY�b�R�U$�z�s�˴k���$[{i��Ymݬ�`B��G�0 ����U�X
q�_$�<��Wn�v� ��͌`U,��^@��Xj2����ke$t,A\i(ɻ3�P�z��n�$Z�\qƚܻ*�ԫ�*�pWݤ���HUW.�/16{q
�*�=Yb�:mW
��g�X�h Cu��$�`�ei��&,8������#)-URq12���Ynַ	ֻ&UҲԵ��WIp�g������L�[hi釦�F� �<����vX6:�tnԋ��U悖
��]j݀��B2۴�m�l��S�5-�� ��nٶ���.CbԴ耮8#��̷D6�ڭ���=�،���^�擥�n�΋/s/5X�UU@.ə��w~{�t  ���8⠡�||&ǛCIX�� QN �����#�s�U>4EEq��M���ߟ�Uvռ�0���n8:����\#C�x�m���Мh��6�笄�e�+i�:�vx�j���C��%`�L�I*��&��ϛR����1@�ɩq�x]��I$e��-��8�/j�;:�-�n��H�.��X��ieqw�6{Qn�=&��2Y�gLZ7�:�m`Z3�L^��v���e��ț���!��X�n�i�5?�{����q��DV�2 �mr�Nւ�|��v{,�9×���n�}բ޺p��v��FJ�u<�bX�'���ͧ"X�%����ݧ"X�%�{��6�`��5ı>����"X�%��㴷�e֌���n\̛ND�,K�s��ND�,K���m9ı,O{��ND�,K���6��ؖ%����Y���Z�
f�.ӑ,KĽ�{�ND�,K��o�iȖ%�bw��fӑ,K����nӑ,K��߻�2f[�Z5�T�kY�ND�,��!Q>�ӟ�ӑ,K�����M�"X�%����u��K�,K�����Kı<�{���2��ԸjMf�iȖ%�bw��fӑ,K�����iȖ%�b^��ͧ"X�%��zo�iȖ%�b~���ӷ��y��=.�O>����-��Ljc�ǧq�e��p<f�0�t;�W�s�W.��ə�i�Kı;����Kı/{��ӑ,K��7ٰ��<���%������ND�,K���묚����.�jL̻ND�,K���m9O�U�>"�q�<�bw����ND�,K��ٴ�Kı>�>��r�bX��/xk5�����j�36��bX�'��ͧ"X�%���}�ND�,K��ݧ"X�%�{��6��bX�'����Mf�2d�d�fM�"X�%���}�ND�,K��ݧ"X�%�{��6��bX6'��ͧ"X�%��O�oMs.�d���r�d�r%�bX�}�v�9ı,?"��߿f�Ȗ%�b{���iȖ%�bw��fӑ,K���݌��.���-3;c���Fm�ti��m�]�-��۴����ݜ�t,Ʌ��oN��?=���7���%�����r%�bX�w��6��bX�'{��m9ı,O�ϻv���=��r ��X!�4���S@��� �ٿ$UU�B�(HҘ�9��w>,�͛%�Q���B����"#QE4��hR���(��(��ﻝ��j|X�*��������s4=���*�U��4�S���z��{�`nק̩m�TKT�Xfb`I�IY�:`jݖͿO������\�)1���� X�#^Eꂫ��R;N��{tv�bܻ���H�V�u.f[���>,��VefϢ/��}��=�p�6F�q��L��-��V�$������H�TT���U*uJX��w��7w]���L�r|X�֬��j��$!�5*e����`oڞ�����IG�������_�����(5��@���`I#��ؘ�c �v)�5�r�U6�[�������p�#{<={p�N�.�L�r��Ie�Ѧ�q>��ݵ`nVl�����!���`r�d���)��8r�MX��7�!��������ݵ|�����*�ۤT�-:�V�{������y$�BS=�֬
���;9+��5�Cj$��dDOݪ��;��X��6	(����`w��ٲ	Ȝ ���w4�
!-ݾ? ww;~���%BK"�������O����E�=7Is9��!�6W��V���v��2=Bŏ]⎷��T��l9�gj�
�0�4!cMWK�;�ΐf�H���4�[\�nx�#q�g�T��] []d�6�鞮�.'9��v���P%���Jz�71��8yl���q�ը�mP�8��Xxv��c�5����]����%�կs�b(n��e�O{�����>���(�Cc�=��vg�����:/j�6����������5��uY��I(I��?� �٠ynJ����|h��6|�~�&,#��I&09%dL�wrwc�+2#x�0Crh[���SO�%m���}4Gu��21��$,�zX�����aЧ��|X�X,B�M��BHh�)��4�r��)����#������.*�����0z�[8�u��,nNn(n���s�MN���O��}�����*cI��U\A��eD��X��3!���nfnI9��ٸ�l@-l��U�����;�"N1��M4݁��K3�tB�2ww= ���{s�%sd��ℐ�7ob`I��T�� ���]�J�HtJ2�7w]��DB���? ��Ɓ�Қ��Ѵ��"��p�bk<S�k��n�|����'<��G%l��'?L�#x��nM �ܳ@��h�)��4Gu��27��n��ץ�!(I/(��*����`������`j�d��1T��X�,�͛ ��vR��@��"�}��4*��(��Ey�Yӹ�'�t��=\�W#�1%1L�$�C��~��Jg����˝���K2�f������y$j$���f�m��2s6�wu�} `��⪓�nq��[W	�v�g͸��xNz�۶�`�Yi���СD]����i��2���M���.���f�ynY�{s�%sd�r�Җ6�'�ڿ�DB�����`}s�w>'��ďW���^4��D@�������jcI�`j��`s�ۆ�s#�R��J��:�脡EV{����y��2~ͫ����󗷯@�{լXE	��ɒh�M'3j�7w]��um��B���(������v���0��t�{^�n�ͷ�����..Mh\��?���8�{���=�X����ӯD6���*�77]��um�s^��9;�H�D��FE#����rڰ75�`d�m_(Q	L�jٞ�%�R��Q���=���s@�e4��h�f�ޝ�͐ND��9����3+6ls5�rJ!O�˿+yt�ͭ�oR'�C@��W������V��j��
ref��TUL�n�vzikR��;l��L/JA�Gp�9�w[X�؜��v�jHÂ�btX�*�Y�LP1�H'n�p��ĭU��[v� ���vۓW76;ZLeg�q/l=�-��pӵ���˱]����� Zٗ�����V��s�JV)�l�©�!x�(	R�D�P8S���Ο��o�6�v͞�*vL�)���UWEʢ�u��B������{��o%�p�`F�"r<���g�(��)� �/a�6<��!�r�:���j!6F���G�^�h�ڰ7��^P�/�9�VٽqNo�
I�y{.�}�s@��W����?g�E��"�X91�`vwZ�2s6��Q��U��3�_ۚ�z�y��#'���uz;������Lej�^fZHq-:�V�f�В�Q=���z����r�@?P�����	s��.��}\����ݖ�W�9:�p����h�x1D�Ij$'&��RS@����9wW�޳@��.K�3#pl�nI����z�a$ 64x@",�,�M�҂?*�׳���[�go;�h��D%2g.��Sm�J��4����6wz�~�vr���x|X�֬�쒪�iTĹ���ua舄���c��<0'v:`j��`s����L�'�`�$�<��������^�^�h�z/�o_A���q���7HN�xw�xv:��'����܆���%��wvbC7C(E27����}����yϪ�/Y�y��g��y�4Fgذ��`sob`�1����07�-_(J&Cyl�*���\KN�]9�������>��c�Ok*�8��c"�`d����8�� �١+�Q���SI5�b@a��$�4IH%�!%��c���kDu�.����c$�MT2`l`7�D('��)@��*; >��|
�'���q}P@8�T� (�򄢒ͅ�=�`~�͛�,��iA���Q�$�<�˹�w�w42�fáD�ݼ���2iӧC*�9W����t�����96c��0?��}�����L ��V��H�T�ꕦzۧ��h-�����θ'k��wGJ4+���,t��>�ޛ ��������%Y�������U~Cm6 �4LPn- �ٌn�t���t������w!R2(�(5��ɠyݗs@�z�i��S?moM�}����M5l�9i�)T�mXz"!N���`}��6�s]����
uw�`j��N�I-8r�N��ؘ��}=��W�07�077���{~�WX�'���o��۞�x��n5Y���#�T�����=#�u�Yi�^�������`sv����Lm�Z���֔�!�ErM�컛�b�∊��޵`gWzl~�v�OX�q��n
c��_zS@�U��$}��{n}��\�+i�M�&�!a�	D��zl�y��ڰ7�zX�y�[�!�����Y�g�J۫�/�vk�����6�}	$� A�
*�X����Z��w~��{����]�4��=��^(���Z��VqE�m��F1!�m�F(�N�t"���;����h~1��!�*���L�I�q��ڹj�ܸ���l�'�r��iJ^8�qX���g�H�4 ޭ�Am��$����m�J.I��S�2�q�n0S��h��H��@��ՠ��][N�۷YŇc'�.[2D���\n�Wt�L��Z�� �('�XM;��'3&���[*���նݶW�n��뷏�^����{5��P��d�L�'�`���?��.�}�K�Vl�"D~�;7���qˠ��cx�ɒf�}�M�}V�_z��컚�m��9)��P���� ߳]��L���Ձٯ� �����)�9�j8�?��}��{n}��_zS@�S@󳒺҃y��Q�#�?f-�`y(��vm���_�f���-{�, �CM7�)�#;k�<]�:�=��Oon�9����gg<Ҷ���q����/�)�y�)�޳�<A����}�|�{l��<pr�қ�"~ � �DGVN�=��:`N�A��wl��.�A���L��5��ڳД%=���=�|hz��E(�G�`����=	%	Ugr�=��X���f��R���H7��$�/�)�y�)�޳@<�@;����9 ��ݞ$��ΞŸ���V�q��r�]�	xn#\�P������7����%��ͷ����`�k�ٚ�
%�C�zՀr��D9J~N`�R}�7��ؐ{o���޵`~�z_�"�>ճ=eK&��N]M6���v��K.G�JQP '�Df�@O��?s���o��@��%��L�C�8��/w ���A�N���ٌT����c�#b�s4;�4�g���_��}�֬�6Ձ���nQ4.��E: 춺��q�;���;fE��m�|���v-�[[2�j<k���< ���@��hޔ�;ޔ�<��!Ƞ�85����?nm��DD�ٯ�s_�ٯ�9�X<�F�<RI��gƁ�܃.�&�L	]����¥Ö6��^Q	Wo~�`zw�V�϶nH��*��F�h�Ff���LADP�.�߷�� �/�(�"h���1��z��%�o~_���Ł�c���̨���U&�\�:Vf5v���M�5�����۫���\��[���yy�ܕ�-_ 利0'w ���A�v[�J�6�!Y��3@����;ޔ�*���<�w4師#j((҃mX�=,�Y�g�/$�V{�j������{�m���&��'����c��c����0;�<a�+b��T��ӫ��ڰ9yGo{����nI���krJ�� �  �\?g���Ы����D�$��Cttݴ�zڹ{g@�]�q�j�Y�ۧ�%�v�s[���'sp�W��.3îĎu[=�I�x%���������5�\��十�c�j��\�[��U�vR���E$��v1Ռc���,ak��8��[�vd�r$�$��h'e�i
�=R�$�p �a�9˕�b���NҼ�2� �Bk1H![�:}����{����?��ZA���"�%��{unä��7+�Z1s��'\g�:������ rA�ǊI3��������M�z���s@���O#��q�2���?W�^��d��c�s�TC�5��JC@�^�@�:`ov:`sw ��֥B���+��`sv:`ov:`sw ��U.߯�@?�␎,�Dә�w�w4n�Se�9�09�6+�M]b����OOA!ϓn�s���h�pA��z�	��T �x.��K2[�m�?���|��-������q��LF�.�z���DPN��{��3�:K��w�w4��4=�HE2,��X!I4M���:g����3� ���Q�LI��I��f�������f�zύ ��h_�;���}��O#���rEWve�07��`vc�c�쎴��Da������m)�8j��v0z�\��/Dycry��;tv;Vr�������Fs�E+�.��:����n�L	�vx��t��ܩ}�Q,I���ڒM�֘�2Ձ���`�����3���c$��dr&��������M�T,�E���aRE�H�b����P�%�;��{��ٰ�q+�b��	�����M ��v�͵a���*���+dޡ6<k�(' ��hw]��n��t�����m)$�NO�1,Ja�Nc��8�;�+�����x{v��tA���M�AA���
I�y�w4��Қ{��=E�a�� I�a�FՁ�nڿz"�J�ή�������s@����LdprH��G3@�T�&��7c�쎘�ȱ^^�
[
���J(����`v�Z�7Ͼٹ?*��ʠu��뛛�y���k#F4�I"iI&�{��}�s@��M ��h�,�- ��b��H����O]\�m��J'��>.�GC:@�r�d��,�Dә�_m��/�S@/f���JQ���j�<��gɵ-�fQ��Svdݘ����vG���y�:�D"qHh�@�͵g(��)���Vg>,�c�6B(��1�������e4�Y�x���nD9�a�I3@���vdݘ�����߾��⚉�T��lր����"ED)���  x�_��T���+*/��@	�R�|/�
PCK!<"/�5T�������П!i����ht 2*�?x� ���G����Q�Ta ���j� ��e@e�u�F� ��T�x�^���<��k-�	�n�	��   8%��m��-��ȢB@��fh�U�9��U*��mri6��	��LPq˶�c�}6s&͉�pK=Nj��v�M�2�B݀�:��*�ۯ:��a����`ル�z��;�e�\��]h.���m�Kr��H$�@X1�ۙ�%�+�=5��s�v����e%��9���@P��Fb�f'm�nV�9�q/n۫@��[��E��6���$�F�-��GY�g�.��ۋNճ�aRi�/C�t��Ց�2��b�7�y�5��U��<flj�jK&ӕ
����c�$�ač�%�^�Y��EE�Wo�I�T
��6�mZ7UjY��lVm6�������!�6Q�~>���-\�a�%��ATU�zM-t�m�ׂcpr<��^t��l��7t�R��;s��tc�8��Y����m�?��G���=f�UH=�m��k�x�m���B���Q�\��cF��6WcgTgA�9I�x9������c��K��T��r�V���ڌ,�͌�-�#�Բoi-�^0v���WY+m�X̶�#�?�MQV$#r�u��g����vM��Q���IcIŘ�c�d�dZ��5WN�쪷Wg�f�Q۪�N'�9lUH�pDjU{<�5N֒ۻ]:��fݺ0s�:[.a͹ײ�:.������y���9��DIA�kj�RKa��'�b�m���ۡ�q@�q�౐kj�v�Zv���si"��@�Z�㇖[q�����1�{����kj�; 5V�Yd�F ���][\�&��:���Hd�	�UZ�(�.&�9�7*z"vb��b�Upa@Wlu�d�ոy���S�=m]��N0œ�#��U�F�`�0/P �Tp٣A�Pq] +�S��'`ۋ���	�JKU�T�I�����;-S��,��N���s�*��^W�ز�'��2�w]nx�t��R��WJ��� �ȥ�~{����=�{�1QCÝ:(	Q��SH��L�сC�D/�x>�mUO�P���\�ѓ%�*ٍ��f�$����X�e�l��Z�[��=�0p�]B���[i�Au�f�u����IY�ᮾ�*��e�Y�gI9j枳�8��thlg��w6�j{a��$�)�2s����%rGF�֎t;.V���=vH�ꠝÔ�
Z�����C��
���|��m��q/Q�<�8-�9�ugd�u��gv8��h���ל����z�mֳ�*�z!���Z�h�jfH�Zv�4�zd��7��V9ݝ�-�HZ�grg[�_;��������σ�Λ5C�U�ݷ���_�7f0&�t���� ��+�˙r)l*j�,s5��IL��֬��V�m��
��
��]3�Ԋ����[n���֬�v՞J!D�g>4�~��v)X� ����3@��ڰ7q�`����BSݽ�X���mKnDےYTՁ��j�����ݽk�%�C��Ձ�.�}L�m��7=��wndH��'p��'qv��c\i^un�%�,b�I�Ł��� �l`I��l��lt��w!YXefI�0�i�w6Ր��Mb�	"yD+���Z�3��X��D%
&O���
���NP��Ձ��j��͵`���w4�u<��&66Շ/B����� �{���͵`nn�h�mQ8�J#��nf�^�h�����V��Kf�"�*։�Z�I�et��/n����n�u+ۜ�^�l��l���~��slƟ�$M(��/u��77mX���菨w��Ӕ�Q#l�p鹩����W�'v�,�����ߒ�U�jLRDd�
�Н��ٹ$�߾��U�VeV�T4�ezP��"��X�!��y�rN�߭X)>�&kj���H�MXrQ�U�����w�X�����V��6U&ӔI4݁��j��%�ߗ�}��s@/[4kU��8(�|�����p�c�m���=��qo>�.Ź��������pƛR"L�RI�����޻�z٠[�s@��S�1�����UCmX���Тd;{��ݽj��n�\��R6�1H&�h�1�&�L�Iz{Θ�y��Z�veȪjnje�v�	On��`v�Z�7�~ٹ"�� ����9�*��S�}�ܓ�ϋ��l��u�\�j�dt��c�6L`I��6��m����� ����皐u��Ш��,ѫ]St���m;c7bz���n+^l��SM���1�&�L	�:�=G��i����y#�������'v����Ձ��j��O�_	�4ӪN��I����V��<�g���@>�}4���1��2,1I&hdt���6L`M��7cWY���m�l�f�}���/��O �w�X����� NF֬�Z��
2Z����Z���i&ȤK%�&�{4I�;�3�ȕb,��^�%wo���7��j�/�ŧ=��T�R\ҝ����tp�h�5 ;l�u��U�;s۰k��y�rIv��ݹ6Vܼ��M�ph�'+��8�mJ�s��HMg/m�շ`�-ͥs�.�<���
�5����W�<Rvݍ�؎��8��gI��s�mG/8Ck2Km�q��6d���Y�A�ʪ�D�Ԓ��z8#nخ���[/*$62nn�F��]r�3d���"�����73mX���E��k����D��������$���������ď��nhw��@/[48�[D��,�b�yL	�:`ÑT��v:`�uI<��$������h��X���<�/(U���Vɽ5U5�k �y���9[^�{������n�xÿF��$r5�5O�P׫oo\�f�ck��,]ۥ�L:ޙ�ө�\Nr9�<�"����/u��:۹�_m��9[^�޲�0Q9S#��f����u@��h ����~��lܓ����]�����Fd$�1��L�$�遪Il	6:`l�� ��*�.�̩i���jÒ����;��Xm��-빠y��]iA4�$S̶�06H�&�LRK`v�����������Ӗ:��M�N��nӭ'n��z<���n�qDu�)��%5`f�ڰ7��VN�ח���=��V~Ͽ�O �&1���_m��9I-�7c��0:�껵qb�1�Ӛj���ڰ73mYiz"$�@,@��
e�%AqPP��;�{�rO;��7$�����5.��(��ua�{w�+{�Ձ}�s@�mzz�p�qȦG�)����#�쎘������ �����ަf�5$\�ۋ�-ۇK�n�`51�㭜r���ӯ�a�6T>���M�z�nZ-Yvfepo�遪Il	�06I��=�D�QĖ)�m��9[^�7c��0$��ͭJ;2�j�S��[�w6Ձ��j�Q3��j���z{���j'1�dR&����w6Ձ���`�&�	@DRHBF��LP@3���rI��$�
Bc�����w4Vנn�ڰ3wmXP�di�(�Kr!��v^���l��8�Ə%��hq��<�:��-m\גP��檦�\����鯀���l	6:`l��M�����W�����$0m8�z�hm��-빠r���YnbRHɑ�I3@�vՁ��j΅;=�Vv���ܼ����F1�I��w4Vנ]͵a�����9g��̍535yLRK`I��d��lt��o�w�}�����Uvռ�0���n1�Z�����/-���n-դU�4���9z�oh���4�<�;��2;C����Ѯ�HlĪ��۞(c���mLS�K)�؃���$��S�NAM��	���:����;Gc�mk.�I�b��:�m�6G3jKY-r*�B	ǩf]��3�������\v�qq�n�r)\�#X�r��MY��X�@J��������UC7�.Y�����3S3�g��9�����1�]�Mj2�+n�3��d�c�-�n���Z�.
6�����~wͷ�۹�[�s@�mz����j'1�c�榚�3wm_�S'v��g����͵~J""�f�除�lj��2��ޞt��$��06H��wU�V���'4:j������;��4��hz�hg���"&(�ɐ*��X���D%	%���~{zՁ����ު�F��dQ<�G��,�n6���ص��[�;��I��Qǫjٰ&"{vĤhx���<�� �����ܠ����{�jֲFCq,H�f��߶oB$@�d$U��S���]�}y��ܓ�}���=��W�P�$��-��L��T��9��������遲GL���䮍A��D8�5#�<�w4��h�Jh��@���cl�bs�R&��7vՁ��6���wU��۶�m�}�������:���&�'�<��kv�n+]���E������<����+\�J��`w� ��$�{#��0*��n�F���h��@�͵`f�ڰ?mn�򈈙>Y[ҩ��.��aU4���޵`f�ڳ�N>PL��,"���ӂf�,�i`Qn$b@�>��f�%��o"��i�F�T �(MrF1��@�� �B),`ǖ�	B�XJڄ�
R
gЄMHB�$$�HH��$H|n�6�ҏ��@�)���D@�4#aH��.j�O@� �EaO��_>��P1XP�ǞHy��~/�ւW�h6�lH�ۡ	!1g'��Z	u2o	X��__>R) �.�����&ƵJ0!BB�Ő�Ab BF���
Q�=_0'���",6�$��6���~G�QTDCBQ(J'v��2s6��s��)��jjiJ�m�(��������lVס�+o�f����dxFd�t6Ձ�kvl(J6�����j�����*8FI190�&H�F4�vױ�=s��uN-�ѹ:�&^ݬ7Y�����e4��������33mX���	x�ߟ�-ە/�j����G&���j��ݵ`~�ݛ ��w���$����^��:jiÖ橫��Z�?N�zz٠wu���Ȕ����x]�08���&Ɍݎ�q�QU���
V	�=����<�(ڱdxa�����f��Q�ߗ�;{�X�wj��V�6�[�a}9��R���YgY95���u5q�\�r<O"��6�F�P���0�Ͷ��L	�:`qI-�M�n)tP�[����*�����W�^�
����V������j�
"&O����C��9�䙠z�����w]����{ĸ8�I�1��zg侽���޵`nnڰ�P��%X��U���%��8�l�1�ڎM���z�����X��� *�t��mP� �Yn�q��Q����݁���:uN����wm�>��j�Hw�����8G��g�z�;�B�@�gh�j�k���nz;!¹�&k�[5��i�U��:n�0�2�ͬ���ڵ�8;v��C��8 �ae�k�k���ň�1�k1�ځY�FP��m�"RY�9֞s�5����:pCl��K��k�r1\�X[5�G��{����q��az�W;�cH����ݛ'�v�8�6���t�8�Մ<&1�iB9���H��������mzz٠wu���Ȕ��U�
�RKă��cI�L	�h�Q�Ǒ�@y1F�z}�hfm�?��&{w�XN�U����)�u%��#
�ݎ�v:`ql���/�女��/�bR4�O'$���L-������t��Ԩ��-.�q=<̽��c���on�p�wku�@ :;P^��>|�y�.��{\��������	�1����7c��(���ɥ-5T庰�u�$��J?`"z��̛��lܓ��vnC�ֽ��JQ��l�2DҎM���7c��lvL`Pږ��N~�����z}�h�]� �A<�L��7�h.ݫ����7zՁ��j��%�.��m5 �������u�n�z`݉<@0�׍&9՝g�8M�t��3����������7c�{{�܀㑱�(���۹�^빠x�נ�f�bE���a�'(ŋ���zՁ�՛64���" P��M	d(�PY�z�ٻj����[t���r!��3@���h�٠y�^��1�152cqh���(^���_��Z�>��f�������\�.������n{/n��X|77��ݝ]rpȸ/gF+l&뀬ˏl�M�vGL	�0;�ؘ��;Z\�(G1��8F�h��h��� ��4=�s~�H-�>�%2L"���07ny0	�1����7c���m:�,!�ő���l�<����'�}�nO�j">��J2'�pA�y����y�kz�Y�\��,F	+�`s�:`~S��p۞L��@�Z�7���8(�x����u�=rl8U�u�=��I�o=�Rf9�v��­v����رbrL����_U�m��۹�y�2�	��r!��@��ؘ�1���遲GO�D����l*Zj�t��7������Vzg��s@�w�y��%)�p"�G&����$����L<���c ڇ��#���#s4m��=��Zo�f���nI��b�|D�����j眠����yn���#�n��L��Z�o�wb�5�E���9�W&-IQ�8`�x�N��
�wX2ZQ�끲�v��l㴳d�YҼ�,����eb�$�K���;\�qR�z�P�t�	t�;�ׯD	��OV9�ω$�s�Qs<��ې.�,��EM�����۟����;�Kl�x�sO�φ�i7����I��je �:?;�{���v���~E3�]s�/��J)W6����w-��&�m=��e�\�w+���,��7s(���f���~���}��z��,� �y1dn- �L`s�:`l������)#vz݃��4���Iɠ{�}��u�sO��Jg2���7�����ִ!LSTJ�Y����#���&�f096:`{�Dl��&�L�I�z���^�����X���DDB��&�2&�ʪ�ZyLBg�&��N4�O1�F^UI4ld�ܚ���\�Nr��[9+6۽�;��ڰ3wmy$���|XI��5�L��!M���ڿ�G�D
@"	uB����}�}��/�S@-�h���ґ9����e�0$��{�=�{���r�y2A��l�f�����{m�����n�ＣiՑ``���;$�&�L�07��`z�Ø4�) ��bC�O�Q2mh���,� []�r�C�c�lүb����"|{?����fp�y�vGL��d�@�����&ŋ�f��n恽���vI�M��݅'��e�M7%�Ձ�Vl�ۺ���"!b�I5�)���Z�;��Xnm�SCT�4Ԁ�Z�h^��u��دK��=EϒL�RaJ94.�L�07��0�1��t$��&;Y�&]�\�땎{=������N�c�wl]��ob$�N�~��wt���Z\�d��'�遽��vI�M���	��m�-9m���3��W�Q2���利07dt��ueڸ� efQ)�j�>��`~��Vt(S;�֬�uQ�T$M��"RM��~���I%Y�������X�=,$�d|�"5BQw�v��ʭ"��j�R��遻#��r�L`rlt�9ݭ����$i�e��f��l�W��[���]�婱��\ݖ�r�e�Uv�a`uM�>ǥ�}�������IBK�����/���F�2I1��9��o�DD��oZ�7w�X�m��S&I��y�HI�25�M߯ۚw]��빠[f�{���ps���4�hBI)������V�w]������o��'�RA�1H�&h�]�}��:��y$���$�y�7$�*�*��UPU�*�*��UPUj�����T_򪠪��UAU�@�+��$P$P�AP�BBBP��P��B�T )P��B(��EBB	P�dBD	P��EB ��P�@T"EB*0 0DX��T"EB	P��T �aP�P�P�P��`1�@T"�@T""��Q 	P� @T  �b*@T"@T"�E��	P��bDT"@T DXP�$B DX�P�1DX�B A`$EB"�bP�#E��@T"��"��T  �E���Q$B0DX�E��BQAd �"�
𪠪��UAU�*�
�UTZ����UPUª����T_𪠪��UW�*�*�Ҫ��⪂����e5��;�  �-��?���u����B�P C�    ��   $   @;�  �(�� �PPQEUA@R�P�(A@    QRH�	@(p  2�@ �� k�>��c�/���a�� ��O�&�����C�g ���=r����_NM�;��b��N��w����n�� �7� X8  R�̀4�2})�Rd&�� �Tn�d2� �K�2�p{���i�]����	���sҚ}F�A�n@p�� (  �E)�%�a�}L�}�>���l���Y4���ϥ2݁�� �^�}9]��R�:kֹh�A���� 8	:z���k�ν<����  ��(� ͨϡ�A���  � ` H 	   $ � � H �  � Ϡ } d�d@o`�p0 -` I�  =��x< �J �U{���F@/`2�{�s�N�v=A�@v�N���p 9:pN�nP/g����7�}{�p������磻}��|
H EEa��1)M4�1(��O�D�i��@�F�eJ��  L  dɈ�=U*�R       D�*�*@4h4 �  j��e��P       ��T�h2���� <��N������=r=}�R��n��c��@�B=�?��: "#�T?�UA��@EG������?�Ñc$QDX	T�'��`
�#"u��d�&��"4�iP�������\C GǀHD{(24>��b0`l'?�4���v�D*�x�a.:�N��%�sx�a��c?��Db���Q��
��E��*x�&u�anR�8d<!Ha��vc�1�F�s	�X2��f.\ǒ�M0�b��;%�hp#\ M�%���K��Oo�u��t@�
R�L�@��D�\�tI���|�s�-'%�i��Ќt�^��s{�7�z^�1��T����^]�!"uN�a���4�B��(FƤ�1$k�e�wy��w�BB^�,fB�Fq�䓬�9��&�C�
����L5"xf��.x�=����z���X��F0�AÜ�a�o��4��NR���� bB�ׄ5������0F`.Ň���z�;h�[C��!aRaBV\��_w{��� Bc
0��F�0��l)�7�Ω���&���ę����A�L�<�y,�tv#1����B>q�uF���;�h��iO<=e2\�N=����2���O:���zFob;L�E�M�íA_{�=y��:ɮKM�HP�9�]y�w�4O8D
i�u��w�1(��R�b���)�2Ve�!����u��6s״"�"0���6)�X4=Zw��Ρ6�-H�
^���32C�xbPa 1#/gP�*\�Ji��F��N���|��s�y�L"��<)� v�&�^>.m�N�f�jh��P�aNzrxxe���%Ò@�
��/�q���t�s9�y$o]�5"Ab�4JB'-�K�),9���	N���C^#ڤ	k
�9;�64�Y�D*�= u^���b�"����H���I�C�鐕���Nu#$#�
`��"B$d199B2%�X�5�q�zcQ�H�i�jI���xO�c`RR!`�"#��^3z
}DbLA��W1MN==��K��X��F$:���`� �p�1�0�S�q��ss@�<\�+����8��1:N#�xs:�=�
�N���f˚�9l��m,�S.�� �!X�2R���đ�Q�R��A�Jq�Č��s����$H!F��C���zO|G��H@�b@0_�=��9	���^ǰ���ۯ���J�N����1Ӱ!\t8u�7�s��'�ބ�ޞ�hǡ�`�0 �^	�:�4�S���ì�x����}w��kt�4�$+*�V��$"CB"�0�i�gsw@����]�7�{;�3n��:�e�c(�`�yF�m�B���G����H6�e�����@�6]1���^�	0e��RR0`���N$q��\+���z�a�U_/�����j7��tA�x����ozs��Nv0�z�-D� D,�i��~t4��tB���� ^��Q�@"�a�M ���B<î�4E�GX�U4Yq�ǈF�F���GT�Pp1"T�T�
QpC�!�7&w�=�: �H6�p��CGML,Nͅrxi�Ǡ�C H\l��B�HD�X�*8��b�J�,h�"�+b��߃��w�!�5d�pz8�Ԟ��d"GHBI!'}�g}d1�Ι1B	SX��#�1��!E�;8z��C�Oo��z�0k��;κ��Vyw�EXá@��0H���8T�!H�RL��)��j�����k�`V73���;N�{	8�	��9�K�!��4%�M8p[��7���U�˨�}�p�j��Wt$B0)�k��̝ap��<��AOD���= �"D��)J¤b��āB$	H�!B �si*@�(J2丌��.�HZB�+(K�桧 ;N�t
']����p �������"F��"�,vHV0B,Q�B"VI�����9�Y���������w���I/������G�=e��#Æ��!	z��XNL4�H��:�qMc�Tt0��W
k��*@��/NV4��Ӂ
�0����/
�.4L�M ��(�l�n�@�����	n�6���3��߮!P��B2Va�HRS� C	BP��`��\%λ7g!��޲2y����{|)�K��a�'A$�w���&a����gA뽵c6W�P40��\B���芃�J�n� E{��"U�RQ�dU0FL7{;6�|S!�%R-te뮎dC�:b%qӳ�;CS����W7z	�\��tM�#���C"@:�jp�y�n��0%1�LM�9���w��	�.��Ǟ���)
�햲L�Jl���*�0���aR]fic
�ƪhF�(HF�!��)�l17���i8i�˛��0�L7dQ�t��^@�:%��U:H�T�\'��o���FE��.i�J���o7}�%���H1�����ĀP�0��=�'~u�=<`Q#IV�!G @b���P�L"�x�7`2S	L D���H�LCF�KL��sL:
��Z��3N�~� q�1�Ț����i �Z��$)�$��i���K��!�{�:��N5W���B\�X�x� i�ID�4�*�^�u�F��4��Ilp�T00�B0�e�d�A
�
� @�$cJ�FD F'���Ӳ:Nt�	!iN���`L��*���)�6�!!��ŀ�`@=��$�(G�RV\4�8����݅�OEc �	^=��9����`gS�;��｝_p6C��5�6$ � �b@h�]W p�`�2��W |�-��� 
���).3t�֓9:oV�+/}�2������q�\ab@�aX�лC4��`,�d�xF��;�N����կ@pRpt(�a����,-�B=1n#[��a�!�U�J�`��8<�%�l�P�����5/�����J-{�A(X�������m��m��m�� @              �            �   ��� ��l �  � @��  l  l m  ��         ��                                                                         �"Y]"�e�	vI�k�v</Z�u\���-�u���Z���ܦ��"Khh�)8��+��\g;vvj6�qm��+�t�a����u`�
��:X��{����qDʬp�σ�k)�:^i`��v��iÎmN-�L~>w|i�nȵʗ�U�y[�F���ML�4�g�u�e&V��vKx�ȉy���S>p]�D���հ}��b�*��� mZD �Xؠ��P�]�X&��ӥ�r@�u���
 m�`'U��   � �s��R�U�����Skfة��j�^y�'@of��U6L�\�PR��!ö؃�Nl7i|�J�kv��`�m�U�ءU��mհ����Ā�-�*ClլWH ^�i��m�� sjۖ�l-�rE�-��8��lƹ!����H@l��e�ɀ     d�8��r�@��$z�6ȼh[N8  [@>��m�� l�q�!0J�mu���u��F��[%�k�t��m���u��  �m�	 ��Nd��Y˴�`��m�m�>�m m-�mlm���Zl $�kh��T�<��l�u���X0[@[d  �@  ���6ؓ��-���� ���8 �HH�$m�[�m$A[P��\-�6݀ n���u[��ݰ[��hGHѮ���X	V��[��f]��@Ye]#�US��W $�m�[[lh�ڴ�h   M�]l ���J�lC ְ m����   v�-���m�h;m�ۭk9�m��� H�ݻkm�N�����(TӦ�WR�P�d�OG���������խn��,r��lp.�� 	���I`m�v�ͤ�n� کV�*�Y�
�b�  �I�RF�a�m\� .�-����r
��b۲�m�k����*��U*E��$	�a�Sm���iZ��JL�Uu*�P le�lv���m�M����Z��]@u&F�mչ�N�   �T���,� 6�ioi�m�uр ��[��n���j�[�͹ຣ��˻ u-͓.*������]�����;@-�x\��X6���3L��*��A@
��uu�Qk�s��M.���K�ۇ�9S# "��SfJ $w$m�l��m :8    �` %M�^�-�l�-uR�K�l��U^���f۴��`-��[%�lۛc��8 -�$H6��6�طz��k5i#vmĲ�� �`�w.Yf�n՛��A�pM�^�m����d�$R��n��дZ8�\��>�lXe���m�qJiK��@r�T�J�R�n�/F�մ�5����U�x�յn�mr@n׭   ����( +K%��5�� �4�;m�m�  [@��NH ��mYƷ�B�㐝8�@���m� 6�G-�}d�g�@$�uPq�c �0�rU���檤&���l���0�� l �κ��n����m*�ː��s���\W[��brmsvbP�&�h[m6   &��[�ւ�$s���o���m� $[@m&�`�:Č�pp	 @m�m���rl�ZI*���  -��� $ݶT�AL��ͪ�D��6�     fu�۵m"�N ���j�n�9����n���%�f��M�  ]6�Z��a [@ ΂%���6�A���m���`�vp�kn�mf�( A�����A�'���A�i ӎ$ [N I�`�im�	ޠ:B�8t�m�m '��msu��w�^�ku6�p	 �,�h� H�j�WtK4�>�}� p��-6��$�:�Y����[\6�n�M-���Pi$�?o���z$�6��cR�4�UmR� =-T[Rܒa -�hsj�T����UT�vm�*v��s`$  4Q�ۛ\6Ͱ�mD��ۍ����v��}'�J����Y��
�UYk�@/=�ʪ��a��S�� n�ۤ�vZ <��n��K�Ͷ�� �Uӡ�Zj��� �V��e]ۇ=#���@j�zq����d*�ڇvV�T��� �T�Ur�G]`�_/�):����Ύ��877S�Β��y��n{+f�T�+۞)���R�UV)�L��DT�m�z�zK��� 8j$�k*�H ��&۰��M��J�aMɛkk�-6�H��5lt -� 5�V�&^J%U�A]������6�۝h  �����׭ �pM0$ u�s#m�@�   ��� ��� �,��m�m������`���im��p�e�o4�m��8��m�  8   H��m     H  ۰-��H /Y(   �a�`m� H �H��mm%+��$6� �m���'Kh6�mp  ���!�8 q�� 2[R 8 �mrڶ�hm�  8m$ ִ�    � -�6�E�z�o�>��Ŵ8�e�@ @��� m���8q�m�   -�   �-�l�����M�`8  H4k�ф�dvm��  �@   ��     �����8ݻp��M  -�   ��&m���a���  -�  �        �A�  ��`  k�n�H@��� �������n5n�LI   �$�m m��  9-1���I�ᤃUt�i�����th�Ѷ��t���H8
��ڭ�c�����_���� �	���]��VT'K������m  ��nt,�&��m&�M�V�p���n�e��� �cn��Dy���-�\��  ���d�g-�]�� n�	  � �^k��ٔ�媥eٕ�-��.�fm�	�� m�`  m������Z��mw:�m�m�  �ݷ �[d	6�2ԙ"���a s� �t5�K� �pI�۷d��u[I� ���m�knD����I�m�����%Y��(��
�*�*(�d�A��U��z��j�s��S$ ��8�i��gQ��D�6�m��[%-���d�� (�vհ ���A���t��lත+���Y%P‭���Խkn�W���avZ4��ζGiT�گ+%s*�tU.���ۅ����r�    6�9m��l-�	 k�i1� �8[Cl��  v�  z۶�M��9�p�Z6�  :�$Tme��  $6Z`�kX;v�i�,1����u@�;�(ζ��$���d�[Az���	 [N �j�-  $�l �d��K�8��e��_�w���w����
 ��PD����"�P����E=AS����z�� ^�H�z�aI"z��,AR�QD|p� ���8p�x����S� �Ũ�ǡ�:��9� kU�D<�OA{�=^v
��jC���{G��@<ASD����D� x j ��^�1]�EV$������
�b`C��: S��\M� )����;�H�(p�l�ǡ�����8�(�C��G�T0T;ET,T�"�S��N��|ED��A�/g �0��;Ȩ��8�Z2� .�^����x�D�QH)�a�\�(��uOTQL��L��<���GЂ�w_PA��* �ȒO��������
#Q"
�E��Z�
"5"��%AT �EU���������     ���X ��	8����l              IZ�ZRe�B�qc��v�viy���]�랬�3�n������%Gd5V%�t���݆�^�N`��]m���.]��v�I�4��l;M�7g�*��\4�6�r�J�Vꭎ��l�If���(b�(����&�'5Ol`���5Jæ�{)Y1����UU���S<T�DUNة�,Ԩ	Gd4�-��ζH�2�nӲ:�(�[���-�ȇfݱ��9ڪ��힋�M 6�����t����K��{)H�d8V�Y`
8�We.�֧5�gdL��*�l�P������'e�4UW:3Ȝ�x�L��B���\�ED�<���㣧#Vp5���5��&V]��A�W&:W��mUUJ&§bql<Qf���f�����<p���V��:=��Ĭ�s���ѵ��:�:��Gm�\��7�1<��^��K�iYgb��R[���Q�y���Na7C�"^"n5���s,n��&M�:�6'�����WUV�vM�� �]�-�#��p�Pr�P�m�
�!Q�ll��ԧ��N�ݹ�:�[{���)�ķ�a�9��u�r��U*հR� ��em�,��l��[X����dt��OLuk������8��[;�`����]�����lᢝ��$m�᝚���**r0�qI��Pˡ���q����n;l<��F�nB���N�,J8�/d1R�*�&i"6=(�+�Sf�]4�����l�칲m��e��w7v�eP�A~� �'x��z�3�t�<�@<A�ͧ��sws�6��` g^M�B�v��nm�SEgc9�)�t��!�5��k6.kK�NtW�j۵���F�MN"v{�H�㜄v;��g���^F�g>Z�݊.�[�kq�Δ6��c��n)YNɞ"��VwUnx���[�:�O7,n�B,�wn�8�w�Ix�3���	.Kdxۄq��;`W���3L)�̽1���Q��c\�_��+�L9lł�)]��G1|�~�w��C{�f�������KC놟>Czc4�ɢG�����0�8�G���M����v�X�+���Dosx��O����/<��)*6DӨu�u�[ǲ�h9�ず��9�Ч-m!=c����8@�@s�}���ϐ�F�o���ʼ#4�33xu��~��t���1HC�ӯz.��D�~����n� I)U7*qƆ��_ y�>���5�KlZ�(��@�Z=�D�9���ϐ�|Z��ZWeQĀ�G4y�4����:�ˈ�q�NN]!���c��۷\E�^tc&��j,ŵq���VQJ���p����F��t�$x`�hC
�ֹ�6��t�<���`�o�J�h�H��t��+ �.�W;��Ƈ���!w���h�is�7Ѡ���9Y��b��y�4�������1�
�k�Ϗ��r��r��s�K/j�m]2�f����I �w����!�m���ww۵���fZ���{�Mw.m���W�$l��9�׻���p����Lf�$'!6����)ZZ<�\�錏���`�1�T�o���}�O�ɗ@�°�5�D7�3^�C놾�*�Op~��nȾq�N�H���b¨)��[��n4n�mf꽮EMD�*&Sr�*�U����]iK�C��"p�w����4>�ishoF�r;���+�2�h}p���ލ��4{��%JJ��b�k\�o�@{��<��%�k3-e�$Iţ�"�;��~����w�;҈� ��%Ip����FTC L�`��@t����`�q2�5S *1P(	����T��j׻��am�܍�  q��V�Y��tm��Ü��d����,�2�w��x��87�$�8$.�Dvv�5ٝ�r���n�l�:x�r��8��[�oOX��wv�V�ⱐ�.�-��5��Ge0m�ۧj
r��K3�Vwl�d�����Xb��ɺ�"W�훦"44rLr�^����O����G�m\�^+9��f�M�-�k<�¯�č�G���p���o�@zHe�v����),Z<���C��@w|�3	�E3����m�h�k͎��0�b����� ��������G��K�!�{�X��ŀ�@{��<�\��h�v����� �6'r �\D��Y7nn��E����A$J�+2��C/�;��>C}
CO�r�3i�Ȉ�p���6B$> ��\�G��O���̻Yx��qh�H��h�i7�t�%���F���W�Qo������!���=$'!6��B�m,Z<��Ul�G�����-�]i�ݙ݋���l����2�n]���lԁth��Xr�*EZ)����tsD�{��.͡wy��+����~����h��Lˋ���q8�J�sx��� ���C�Η/�fRYk�����!��9��w!(�v�x��[#Cy�5�����m�-a6��<�q�v�5a�]�;7���q7=��Nji�e�J�ţ�DtsG��I�C��8�ZI("���9���5�47�h@
�{��$�)P�⼯Lˋ�������3Y�H�E�kdhk�f������{,ah>��ܽlz����͡w���qh�y7$��i��8{�=���v'���q�;m<q�C�Y�l�e���qy������x�+H�rM놛�Cgc5�2��fRYk���~ 
UT	�bch{��&�;�	E+����V�H���rh�\4�]���V^$�b�� <ܚ;��|�K�q���6PEb���Gu�]ϐ��*9��-����h  �Zq^���	�f����lN�:�[֤����
M¬t�ƀ��d�5p�jo=�u�Wks��L6�i�F��%���x3E���htܼmQ���g�3����6����z�tVGr�D��D���YŠ�$���.d8�cL�+�Tq��p�P�����{�]�z�u;�k�c�3��@���hq;��.��ϫ�]����m�.w���o͠<ܚ#xf���V�È�q����ɣ�p׸{��h]�b�p�Z=@y�4{��|����V M���nM놻�!��\aW��1^Z�x�{��P 73��͉w3��vi�
*M�۪���:%��n���Ό���k�4���-��*�h��N45�;�ܟP�����d����%L�����h ��$PbBQ�����u�M�C��8�ZI("��nI������m�OB\&��*Ѵq,Z=�7܆��i�&��ÖqR*�C1�45�wM�4w\5�
+�j��AT���0j*(o��Mk3 ^Ӂ�gv�M��H�d���nF���W�z%���Ww6������7x�,�rM�
(��R6���_��*�fW���\;��<�����򿐁/�	���̀f���������z�x��%c\N*u(�"Ԁ�Bp��كa£Q�Ѥ���@0"D��R!1�HB1��`F##�a�10�k�1�]1`ڬV!�	)�ΐ���\Q@�	���Nꍬ���a�<�J���jA9��Y��
>��;1( U���AU�x�� �:&y����ef�R�	G�H]�+F�m���? #ύs2Ds	Yx��Ś<��ܚ\5U\c �e�a��l3.a�q
H��ofv�=J���e撋���d�1��p��'�h}p�o�ލ=	p�K,�F�J���p�7�o�@sro���%yyw��V�È�����7���p�o���B�X3	ţ�"��G��$
]UH?�$F��������M0�7x�Z��O����ӑ���q��v��r	�'�lcj�c<������!�/%hp]��������-��9�5�����Cf�%V�!��Z4�ho�@s�h�k�[h���%u�4{�@s�h�k�r�ĵkJ�D$��I���}�o�@OBd��*ѴRX�y�5Ϯ.wr/�Y����D ���J��*�v��  9�m��&c����ӛ����K<�G@�'�����F�#\�bz"L��sq���*c&�Hv<1���G����t;�is�h��W�Ǝ�7Ϳ�����¯&똵!��q�dj�U�]L"q�b������D��ET��q��{���w��dפ��L7��>I3������b���'+�͘��A�h��F�������G��M�����"��qh�H������o����J���X��nM�������b9Y��A^-�����ܚ���QV���hӑ�����C놞�
�?��G�[��6��à�f�f�ݪ��-�M���@7N�Y�v��%u�<:}���G���$�B�܊�XH�9TH)#�^g���p�?r��З	��ʴm���Z<��·̶4Jw�����bfe�
�Xqr47͠9�4y�4��/��1V�G�D7&�.��U��mۨ��R�Gn���MÖ����v�qv��I�]�tu�1,(`C
��V-b��G��\�!���8"�r�+8��Z<\����hU]�b�#188nDD��̶5��X�� A�]T(�Ͻ��w[ŷk3-e�J�h�L���4x�u���ļ��b�)�H�7&��P�]9������T`4:�%I*!��D��n;g�؋�o[N�������#�T*T�]3k�̸���ܚ'H��e�
�Y����~(��CRO�����T*�r;3��1V�G?��M�7�( �ԑ�޾�
��\m�`���hq^A��0�'A�@��=���ן{>�ٙIţ�˯�H�{����k�\
��v&��>�>�{*����UI�ve�u�e����M�w�q�'	r�LKM��{�kuL
�����u�d��^,�I]b���&�.�|���-,ŉ]��Ib�&�,|d�w���w,�YeZ�W����\��K�5��|w}�������d&��Ãwm��&�$��.]-�ƒ�a3m�  ,]�T�ҙx�Po�u����`��պ)ں��ty���Чm����B;�3ف|Xx�ڛt��j���DmT����ܛ��0eweәS�uE�v���n�9���).�����qt�<NMK�c��)ӊ���-��vⵛ�d��,��v]��i�N''-��w.f�g����D��S^T8��/<�w��::m�W���:�\�V����nM._�I���SP�\C�Ue��$W���7�#��i�%S����8��WٙsK���3�řU�%A8�'NR��{b�֕���J�>5�[&#�^$�+4?����e֟fe�ݺed���cc�R�^����nz���gi#�:jKߧ���Ű����O���p�o���\5��w,�YeZ�W��������� ��q��2���S��r-����N�2��1V�,8�I]�~I���ܯ^akQ8�P���kJ�39�����E �]��5�E9U\3���?+��n�P�.�ߟ����ۮ�b9seNpA�K�6�ٲ���|P�����w)n�D��I?o����w8��b�]�8�c�ڕ�2�+GI24�
�]��Io�I;���\������� �ؠʭ,� ��H�U3����a���c�#�!D�o�f{x�q� ̸�wk���tJ�R��.�z@3.(�� ������V��B9'\+�s`q
`���J��=�%s�4�NM�ˁτH�8�E ;��{�\��r���n(F. ^�]�qp��2�w���5�����|3w��e� � �� �nRU?��� �\-� ̸��8 n!B�H�V8�eZA���K�*�#��~�$����M�\r���C�n�P��s��w����)@�P��H)�T�DB��Ue�&�x;����<xU�a!1p�tn�I?��$���qp��ܠ�Ƞ��#��A����.uU�H�E ;x�X�R:$t�"��He� ;z�{�\sf����5R�8�E ;x�{�\�� ��b"��B0qp�\�3��^= �$��y�D4;eQ���
���	!�\c�Ą��"-��.���d`B�``&c*BBX<ʺ�X�EsO!!<<�q$$�;0�,Hu0a��");b,F�Ы���$�XƅxQ$̛�ͥ�3|w����x��0BH$$�R`�"�X,�$`���A�@�B�	$%.�!9�]�$e�U��I$�I 6��$q$��Zێ�AÀ [@              ��t9Z�l�o���o[ �8iVGk� ��]�OU ع��9aN�n�v�t6�ܧ[+ԯ4��^��Wn4܅�7�h��ϛa"9���v�*��U��֕qv��:�ʐ=� 1E$̀�*�a梪�U�t��R��%U�B��K���F�lRgn^�R�.6CL�-.S��Z�WRl�uv�:ʧ:z�O�S���,` ��X.��<�;i\[	�+q֪��>^��p�d]�'r>8��x0�������� -$%,n����2lqj��]�WQ�����d��'F�nH���pxZ����r�eP�9%���Z�Bu��S�����s��m�ӵ��r��}��z��vQ��2'Hs7e[pi�I){-��ے(��,&�e�S���\j�=ͦ	q��.KW^���x��\[��\�I���d1)pWr͞r�p���m��hn��� �e����;���<]����n6�\6�J��&��M�k�I/8���p��J�][��+r��f���ZN$m����
�
@]�a^� �`v��`�u�m��O�e�N�I]��]�$jk�Mۢ(N����iIc���n�e쭰8j]i��Z����*q�pA����'6��v�c�f"j��q�˳ݙ��]X���0]/9�E���@^�tU,��.��r�'v �j�nv����.�x���7n1Z6ḩ���2W@I��Mj�q�l���m�V��k�M�|�6�2��*���̻��I�8������] 7l&ۛ���!�?Ǣ �(�=�� u�^���A'yy�������  u�v�9��Y\��w:ǚ�f+0�*�f�0�\���������x�Պ�v�IS$t٧�Z6!�l�ӭ�16�۶�f��㮣a �z2c���%��\�'kv痎&9�:-�����ˈ�Z}��	U�tЁu���x!^5G[ϗ1�h�6�U���m��t�᤻�-ܒZn{Rm�U7K��gԏ\��B繝V��֣��������z��.x�f\P���v��RH�I�4��B�(]����]�8�Qy�Q�9Tܨp�I=��UWm�4i&L�ʭ�z`�$�"5��8�g �~ !V�q@3��F�Dt� ���pn�w"�~p��U3��;�.����{B��>z�8��8Y��n�N?��}�#�F�G$��n�ˊ ]�����.��^��9��R��w"�� �"R��i*��$��� �Q�ښꈥH������8o3������f�P�ߓ����)�mǤ������J�q4�Wit�0	���Au�ǪJ���U$��f?��廜\ ��]�8�a�y)#����`k���b�V��f��&)�L�3�=�z����Ъ����lP�����}�$�����zJrJe�g�<��!U]�i%W8�J��>���2�����p	:o�{߿qpǤ8�%�#䁀N�w�IW2ZK"��%�&�C��K�� 	��SIf[$���KKW�<��Po�q4S�J�1���I���{�.x�@����pNE-b��/�5�w�4����[�s�$�ڟ绞:�r�)�����p��.x�y}�܊~�7�N&���N8�|w������q@޹�ꣵ�6���lQ�S��f�ˊ v��{�\^jm�NAU9*W��P���'}��I���A�Ŋ% b-A�� 1V �)���  bǝo���>�xnz9)�)�Tk��\ٛ�]���f\P��T�B����6UDQʕ(C�W�>[�9/IűW���I m�y���;�H�� ;��X^!�%5JI$\�����܊ _��;~�.�ռMϥ*�p�� �� ��qp����L)T�
`��f�o3��f= ��w���RR)���^n�pn�7"�~i&����_�����o�[@ UU�^�P阦7H�
ܜu�����-0 *hI�t2&v�&˻D]�iw��Dj݃e�%̶�0�m�*T��7;\mF���1	[��5W���F�~M듡9��f_k��n�\�s�ɑ+7c=0��zq	t*s��,裞-�S�(�9Hm����V2\f�Xm���}{���虶Ȼ{V��{�H�������3��(Y���UTa
���)��7!N.���e� .�?�}��o �Y�M�C�
�Jg �ȧ��Uf�g���f?�jd���*5��p��.��fdPۙL�@$�����3�̊ ]�max�����J8�\1� �38��� ���}�������;'lK���"rt��{c����������*pr���hn})T��� �ؠ�8�� �z@;yD�)
����Inb�UxRErz4��D���I|��.�y8�B�n>$�F�[�"KmI=�'n�W��ϩ�S��f= � ���u�?upU��M��'*S8n� /1�;w�\-� ʻ��t�DJT�%��N��݁j�M��m`��IzQ��L�%%�L\/j��p7\�y��2ސ̊{p�9*8�o�^f�s�}�Q��@3v(~� �ax�����JH�\-� �Ƞ�ID�/q�;��.���t�D��� �ؠ�8n����_%Z�� ��SP��J�. g��;w�\*�����3��SNw��k�Y��y 9��Eېݯ���tu���u�q��n���e^��"����Y���qϩ�)��2�jy�@�p�� �Y���8��� �ؠ�8n���ef��Z�%9%2��p3\�y��.ܴOUX]^ 
��kB$���,�r�A����\+6�� �� ��.�4�����D#��*�*�$�X��l��:.�����A��uM�ݞ��ct�w�m�7� �Ƞߜ�{��77x�8��(��76(w�}����HoLB�MʅA�\ �� ��qp�_}U��@76(z���:��n8�|/=��2�j��@�p֬�Ji�ϪHS��ef�/"�z���. ���.���Hڐ����  x=$ݳk����t�6蝩A3ֳF!V�wTM�<��[H2gna�D�Ü�%�/\,�Z]������L\�<rX�獴�S}�l�;]�H4��ѧ�^�ZVE#5k��n;8��vw:��%c��ln�q[�c��fۮ���\��ݦ�YK�������v0�nޯ��;�o��u.ضa�u���b�đ��/1q�i?;�� ]�_}�\�� ���9%'U\ �� ��qpǤ;�@;�*�U9H�ES|/w��^= ܊ v��6��C���(Q�"��Hw"��p?/�e�z���/47"H8p�� v��/��\�� ��}�*��}76���]��aм�c�;�ɶӽ����X���t�3b�w@3|���.x�@2�(�ާ�ݭ�����I<��xsE�~�E���Z1@4"��"���͟y�����@޹�|�Qu�n�SL�}RB�\5��e�P����7�no�.���6���93�nlP�E ���p=�J�g�tɱԍ9%'U\��@<���ޮ���@2�(���1ѷ8v���&;lh�8�����#zB3f�F��/}��rGJ�
�)T����77�\��i*�1�	'��J��4�c�R�a�(Q�"��� �Ƞ��}���UG��<L�� ��=�����f�O�'j�ps�!LhJ��&�]"z����d(<�؁�j�b�At0 �{���D!0m��5P�� t�D�V%H�M0H@��B���]d �Ȱ�MH`�H*6�Q9xA�(B�L(j!�a$� ��D #���� p}H�&��R���
"�x����؂: pN!�����c���3�"�IT�E�/=�y��/���}w���*n:� �����H^E ��6I�D|�m���Zl�.�ۦI5�,�`�=�ݗlyN�WI[o�����B�;	s���@2�(o�^\���qp�+|�iʊ���8�� ��P�� �zO*��d��F����������.�Vk� �ؠ�Ǎ8ꤥR
�� ��qpǤ/"�뷼P�3�DԕPr�\�� �Ƞ��}������ߢ�����c�1�6��l2�r̜ѷ�-;�O=u l].�]����@;y�{��/��Q���:��T��^lP�� �z@2�(�޲:�TGS��e��pǤ/"�v�(ij�$��8��� �z@2�(ob�_ox�q�j��**NGL����$���p�����$���M�H���>���*�B��
J�@*�{�������e���l  �{i��]0m�c��0Qڥ��n�SY�wn�mFVw6���3��ӂ�Z �{��[���z��<�jSm���A$6v0ǧ	V�(�����V�U7\�|m��jӠtnH족��p�uX�q��gy���\rA��C'&�n�,�n��\�����}���߿wyNs.�͆�3
S	l,̗[&���22�u������x˺� 4���O!/~vߏ����� �~ y�q�:�}R
�� ����~���z@76(m�2����	����H�k���C�_|�U�� ��qpfŭ�܄B� ��76(j�ۚpǤ��g>$��R.u�P��8����@:���UDI�b��Qɺy�Οt�oA����9�њ5;3V_��y4��H^E �^���f��p�A�pǤ��/������@2�� ����;�3�6�EI��sb�v�*}�� �z@9��#r5$�:���b�z0/�0�Z0/��q�$��U:�y4��H^E � ��T�r��)J�G�exy��3�]�Ѥ���-�]�a3���j�j��� �Ƞ���sN��k)��*AÀflP��˹� �z@;�Fs�ϩ���8���}�|����R	S��<��l������YI*	�T� �ɧ �z@2�(m� �Y������nC�^= y��_ni�36��Qj'��&��E:�m���=��ѝ��A���m2D'#�p͊�x@/�4��H0��nF���U\�� ��À^= y�q��P����ɧ �z@.�(m� ����GA$n�� �Ƞ�����%\��p����rE_J�p����@9w4�Ǥ V����[bA#����e#�=��v#qc(:�f�q=������dq�N.{�@9w0�ǧ�A��@2�y��O�8�\/'�x�e�P��<�Qt��HJj9"�!�3_��E ��(n����\m2DBTt���@;y�sN�6x�w�TnD㔝UF��b�v�a�;oH�E �$�(@@�$Qj�QN��nu�ix��-�  v�E%�1:�/A�����lf�L������ä� ����$L L�Y�uѵ#x���ݜ୍��s���Q�n��6��(��t�NdbWI;t��^Iӹ�\m�����m}������9�'=��6,��{v�ZN@e.d��kN+�����&�I铙����w�{�ہ��[����sax}��T��mȎ�ۜޥ�ث��7U���}'S�"�F����O� � �o"�ma���#��7�zO��Dʼ�K��4���ի�]�p�J�T�D�� �z(^E ����;oHf��|ԎH�����{}� ��kI-�q4�	=3y�%u7�s-�ٔ�m��/2~8m� �Ƞy ��U�R��!:i�i�'Ј��i�_�/�՗)�-���n��0��i�p���Ӓ*rk�@/2(�Ƚ�(/2x���y�ӕ��e��K� �U�B�h"O��8m�<�J������q�N��\=���p�� �Ƞێ�<T�P��:k��J�w�8�� �Ƞo�*�oզ�#d��H� �?�����p�� �߸���u�T6C���o��<w=Ǜ�s�-��mX�MfK]�o�Sd�"2C�o���@;w<p����8�����qp݊{��&����^dSj���q���Qe�!��"��'�B�Р8
(]�Ƞ���Z�Jj9"�!��U�<@3v(o�@��^g�z�W��9QF�GL����.y�����*�i��✎Wғ*QC��̯Ng�G�� ��ݚ�ӥ3f��{�����s� O~6پ�ۼ�����"�wn:T�S�
�T6��o?%���f�� �E ������C�l��I��^= �<��W��y����7��D��2C��}�I�� �Ƞ��\����!<D03�Ϧ�軻U�^+C1$�"Onyt��y�@�/�N��qS�x�K�w9��$��\�]�m��6��G]���-2�6��8��o �z@/2/$�\���P���!)�4�N.x�O/��E�E ��P^g?$�����9r��J���3v(o"�ﾪ���\5��e����S�RuU�~�/��Vo�(�� �~ ~��W�� �dt��$F�mpf� �z@;w��BN��� @� �
����!H�)0�H�=F���b��Ƕ�I���! o�I+(:jD_��� ��	��	~aQ}��l<;�.�`�D�F$I�Հ�DhE�7���FB� He�a#J�2�zހ�ł5"2#*B*��f �#�GwwO��{��~��h�� m�8E$��b�8qoS�C� [@             UL��-STuPm��ٺnt���X���-}b�,���&K���"��ni�&��赺��$h�. ��1�v�u�lZ:6"��ll6t4�gnYv���)�eb.,獲ݩY�3<A��a��kax.�\�3�4��I�2cn�N[on �r�έ���c�99Zv�������Rn�uF6���:n���Q4p�[�@��q@Ҝg���%wX ��ے j�ҘZz݋�㢰Í�B�Uq�]�]YH�E���ZQ�֍�1sA,�Tf�X�[�۝����#y��6�Y:� ��,i �-Th�{s�zX�A�qfM��xm c"�Z�l�#���UQt,=��p��*����\��qs]��Z���͖�s·��*]Y��0qr{k�Yɻ"�ȼ�6qZJ��6r��
�d q9�3!�^�ch��<���Yu��\F�R��p�KGfwWX]me{t�ڳ��1\:�����X��s+$fћc2�ρ�2Y�kex�Q'�BeסU��9�UR��*��� Ͷ�Gk�Vu�m���05uH��6�j�Wk���a%U�n �����ZRZ�h x6�iL��R��J�UUYFyYS��d�:�d�(��|�u[�"��7<E-۵�=�=�x!�Pn�L��fcu )Q�wZ�� T��6��E^YUd&Lt�f.̝�{gٝ��Ƚ
t.��u��^cq�G�;�6"��6���f! �Ucu)�jv���u��"����nB˒l���8/H���@OT����y�)Ѐ�v�@��z�=����~ߵ��-�ޱm  z6���1[��nvՌ�vٲL��%���XӪX�5uWQ��Y��U<\e��R�d��O������F6��֎x�ۛ�Μ�]'=�Ѳ4f S��H����4�[Cd�<��k &��q;= ��bev�V�إc�j�Η���Mu�h��
��ά���-���'f9籸��С����.[[��GkN������N!�4┪T�+<�]�Pߢ���w��{|E�j��F�!!�/2(o"�m�qpǤ�\YUU>�GM��/6(^g �z@;w��\l�T�S������\5��v�(W��v���	N	�$�����q@;{o3���b+`D�
��#��|�:y��gT�1�8l��������O���4�OD�����P�E �y�_�ݠ�~ �i�ە77��9�RO=����'i"�H`�I@����kI+���\�a�!s��M�u$F�mpݞ8��y�@;{k�9*'�RF��/�̊�ؠ~�������r�*�H8p݊ �]�����pǺ�~��~O��'�64=�4E�3r=���r��w��1��	��.[��~_�������pǧ�(3v([�8ӒS�S��^d��/�̊�ؠ��0��Ԓ&�8��y�B�˿1�*�e�B��$�rgI>y��ԍ�)Q�8n� ��P��8���-L�r�q�UQ�y�@?+��5��^dP�҅d���L��MŮ^98�ę�u���L���nx{rV9��Q�\�&��� �ȼ�(/=զj��ҩ#p����UFn� ��P�����A�|��M7B�!�7ފ�ȡ���7����7�� �xV*q�������f��]S���*q4�� ҰB �z
������Rn(�:��8��O� �z@/2(ob�~�$�̆!��[�ǎn08�.誻q룗d��-�mt^%�wq�qN����D܅����E ���۹� �5��#RFH�GL�����/�|�M�o�7g�^?��Z��u*GuU���s_|��Y��7b�w�*�u)Ԃ���y�� �z@/2(K���U縠�3A�M8�*�7x�@/2(ob�v�i�"����BJ�6��NI��  .�
Ӧ�S�z4�i�Pqd���@����^W���D@X���T�i��;���S�:֡���
��m��rl���ݵ�M�n��8�:��2�j�]m��GO9V�Ƚ�b�)vNZ�:�ER�a�Ӕ�M^M�[��[�6�v�.̏5���3m�[�� �N�6nn�r�����v�.��y�����<���@x�B�!`_���@;w<~�%�/�_%l7�� �-��q������r����T�i%W8�K�L;��W�6m~��Iԃ�S��o�?��_Uf4���PR�m���mSdK	 #��4�]��B\���\�}ZIw=��IQH�GL�����W���/2x�����
��mR��݁qq�7`O˽k�y�"@�/S�c\���"�K�l4���KI.T��$�@ܥx�@3�����$F�mp̟�R��>�%�M��H1� ��S�/�Q���ӊR�#p����� ��(n� �׮��qHR#$8K�[��y�@;w<p����T�'%9Q9y�@/�䲳�t��x��uuZ+�U@�CMR��7C�g�=G>��]�kJ4��t�m�d��4�3��~���pǤ�����碀v���	��&[ZIr��!Uͦ�LG+֡.U<Z���ʬ�����M�bV�Y��i-�kd�3��uO�I-���-c�:�#�:��p?|�7�P̚p����f� �5��pU���/2x��Y�� �z@;~�~X��(Tʄ 䔆U4�S`�yO�0�8����b���L�g�z�.�*[}����޶/����̞8���*���)�7b��I%T^lP̞8��?|��׵Z�J�"�.����p��y�@/�qʡԎ��,i,$E]��Us���T�Kd�!a ��HSOa���)4ܳ!�be����ڀy|�n�p�E ����3�tY��9s�u�k�E��t5��l��L�˫��*"E#RF8J�:���"�v�x���%���@;�-��H�N�64���K\�hi%QW%�S���)�=g�)�9����.��P��w�@/Z��j���H�ZK$�7��Uv�Is��K��#�]������N)
DRJ���/� 	y���]�CI*��4�L
Aw7��-�۹l  ���h�usr�g,�n�7�dм<�)v�J�P�V�e{D��Az���K���dį�wa�/X�Zӳ�[!��k�S��A�r�'gޞG��<s�����,��n�nD����neZ�g��n��\v3'nQ������%�L˹�nC7d���(|i�����[bE21R��s�6�v�c�Jq>{>�n����'�`�"�'�t��q`�ۼ��Y����$�A��@.ߵ����R�I<��4���D�mI�/�
�ϩyf�H��G"m��6�� �Ƞ��,��\�=��;�=�mBD��넗"���D�wMO�P�Us'։>f-��H�N��\3�@;w�\+6����UL�(*q�q����'��LBi�t��w��y�k��Wo绻��~~��(mtݞ8Vm@/2(�� �c�(%�PX-%���]�h���� B�PR!C�B�����/���E ��(n�������i�	TE$���P����$��2~8����"�U(Lt��qp�E ��Àef����$���Pǿ��:���H.y���?$��-{�����@;ꬂ�q	��jUI���h��p��i-d3�՝ZD�/wm۟qY�1��x��^dP��@;w4���n	���#���O}�36(�O+=PYk)��Si�Tk�fl[$�������|cP"g��N��«�$�:N�Ԉb�0"�F�z4�D����{t:H�
�l�7C�,n&`o�t�B0����F�¨�\@����'9���1||�+��](�@
�:��ET *_�4Ã�(v> �y~��'������S�:NECk����=�����~��E �����E#�(�6�Z�J��K��/3ci+�0�[��_���*0�`��E*$:m�h��÷�7�pu��@ݷVg*��IQD�N��)%p݊y�@;w4��v�k=P���U>e4�.X�J��}�\�v�������S���������E�3vx�W� �Ƞ���^)*9�Qț��z�1�h��A{�'@� ��˗\��a�T��U(��n� �Ƞ��p�ڀ~�ngi��ب�Gk8��9���>���p#���ѧJf���w}�zr8�:N��V�~�۹� ʿ� �Ƞ��S�N81ȩ�\�&���/��6�� �ؠ�~k18�(�I� ʽ��E$��*��� ���z�-M4�(�TRJ�~_%W���Uv�Io�x��I 5�i+�Mju>e4��8�{b�~I$�3�t	o�D�mI����ȕشUYWv� ��uAvI��-�X]^S�F��.�`t-��L�2&ɸ�p�8;K�`�Z�$�npʰm�òqv�gd�)�k Kh��cm���o^T�W�&H��ג�G�n��7f�e����CN�M�v�mtJre��-�ɣ�]��gWH;	��kb�gJ�%mw��κ߄�V�L��n䋅<''<��Oj[l/�B(M��r�w���>�uMc��&��/ޟ��{P̊{�@9K����T���{P̋���퉤�T�j� ��  	�y)w��l�R*Qp~��"�v�~8U�@��t��@�.&�C��� ���A��U4�W������u)�ۅJk�^dӀy$���y�����@9��(�T�M� n(6&�I�t(mb���V[[��F�i	��ƜDN0�5���2�jy�@/r/�%�̞8��y4Ӏ�q6�I*�a��4�\��R�of�*�P̊�7>n�5>�-$�D�w&t�@UP����Ir �>��4A��	ԃ���{��e^��i` ���[�bV�a�ܱ0��2�� ���\=�@;w�. tʬ�-���ǜۙ���XG|�ZVM��;8l#npq3���F0�#Q��Qt���^dP�3C���W��[�B�Q"��F��lP�� ʽ��E=��*�<��
�	�
�� ��qp�ڇR���@/r(�X�U8�(�I����i*�a����K�"9U��$���E*��W �ؠ��sN�{P/��uY[>�ӊG@�B�%�DHn��\'!���y����{?}�Q�����`{����p��P̊޽ƈ5S�:�u �ɧ=�6�� �ؠ�~K�T]+��RT��T������E�*���@;�<p�ЍF�tT�:���"�r�i���z� 3���"{�W�4C���wvI�MY�M�ʔ�Tmp�� ���g4�Y�]�P�|����[T`�L��b��fG���e�֦y��㵃�:2vG-@ۆ�Jk�^���2�jw�y/�}���@7����F�H�8U���E\�a���;Z�{�[]� I�13~��;�������0���:m��p݊˹� ʽ�J�7�v�KU2T*�Ȋk�w2x�nZ$�h"O� �5T(3B�
�Ι����u��  �7ye�C�N��to�Y-s��n��QiC'�\����֝�+���u������j,�[e���&���vѱQ��m��3�j�S�	ݛ��n8��+��A0dP��s��O��]��"�Q��Z�1�Ɋ�-�/$U֪UV�k��'ߟ��~;?���[�ǁ6����7k��'=��vv{�3iMy��ݾ�ݾ�*D�)��kި�E ��(.��Ѻ(ӎ��G\7b�v�(n��6���Gp�9dr�'UQ�����p����+T7b�]�d*J��SpU�j���=����^�P̊���k1(�eI� �ͨ�E ��P��8jj����ZknJ��+c��j���tƋO/4{����Ϯ�Ǿ�U>.&���2����7ފ�Ƞ���6�w0���7M����8��(/��_���K���O���=��4*d�US�� ��Ӏ]f�?|���ؠ���^�����U8j� 	� 	������K|�%�q����БF��Du�36(���M^lm%˷դ�"�%ں�Q�����g��Y;ml��-9�v�v�.�QG��1�H�#�):��t7�˹� ��T�"�]����9M�*>�ɧ?%�IU[�flP�� �f"��P�̵��"�IUSQ#�2L ^���|R�����_6f�����~ݚ���eI+�n�P��wsNu�P˘Sn}��}2ƒUV�It	=� w�\Idgb��@'�Z�W����)�{y�n6�O�뱭	�3v�F�\T�H�[~	>nh�K�-[h}B����%��D�ҿ�)�����2��2��Ƞ{�����U��(�
�C��K3i.r�k�""��V�W� ��#nS��5�3=���y|��z�0 _������6:p�ASp�5�32x�Y� �Ƞ{�b���%*r��
ۣ�ݗ��x|Q�Ѧ�HiN�t�:���e�Y��%ۖ�-�'�!�U[d��� ��xCS��"�W �ؠy��+6���䪌ܚSn}�u>� ��P��p��@32(�͍�m7N@���J�w�8���J��i_A ��vK�(t`n%�sZ)Àeg�w2(�� �ni�>K�VDJ�!F�������B����Ab�����'daE�F����!������D�GR�^�� "E�b�Ո�^�<��5�(;9���N�o���������[@    [\�#m�-�pHp h               �Nۣ]���4Isk��}d��Q�NÉ�����e����h���Q���B����ʃ �UZ�4�<uf��6#$'g��^�l[��\/Z�kZZ�!ȵR�ɺ�b�X+�.h蝁aU���6���x�R66N\��.��*�Y}h�F�\��Ӝ�U�I������@��HŪx�&�#�p�E�LD����o(�wh��0r��Yݲ*�ʹ�P��{y#nU��ctܣx�=�L\Ke��d�	і�i�mD�\kKJˋv��N{<�u�gEr�g�(Wx�N���(D�$L�*�b�Q�Wj� 
���c�'c2�Y՚,�z��{g^�zT�@��u�2���\�����	u�ჵ�Z��m�^�]�x��ֻ6�N������r-$E��I7^���6upz�k�W^�I=���`ums�9zK��*v2p�������!����Vq��<�ul�ݍ:�nF$�=Gf�-���w[���S�SZ�j^�؄ٕjU���-���N��2{l�[�m�*�2�H[  ��6�$:���:�U�.�J�[3f�t����66�!�T���/.��d�6�m�kA�JK\�! ʠM��l�[X-�:I������g��!h^�������c;4n����b���js�el�/,���@�g�Qv�Űg(�Act��b��Wm����e�OCۉ�%�ݴz[<�a��=�UZPKga���B�8��r����R�5l�ս�t���D_��P{R��N���J������@@�z����dG;I6�  �osL\���R�.�%�4�X��it<���B�9ڍ6�`�[O7[����r����L�A�=Kf:�mĀ�l&�G7-��t�RX�js�����L[T����u���HժR��l�iR�>�=��ٺ�z���83lS�M;VR�a�Ϯ��n��\y{']�������u�-�Bt��,/eլ�M�v��ʪ���n� �Ƞ��?/����[W�T��r��)�>n�5�3?E �ܙ�K�-|��We���^Z��Dk�fl��2�j�Ƞ{�ј��J��*J�~�V��@;���@�������zx)���eI+�wv(�E �^�p�ڀ��~]��%yC3s�{�g8�۱�Җ^���[�M�6zc��|�Np����uS�������qp��~_%��� ����NF���CI=�Mh
�WCׅۖ�>�I�ȧ侪;J����Dqp��@9���@;��.�ȍa"���#��ؠy����y}Z�� 홼��Jt���F�g��~_|��oW@��T��@/�
�g�AS�Gr��N*�k�̪��@U��\^⯬�n�z�mt�� �ͨs"�]�S�Q�'�m��K�n��76f���%�bX��]ND�,K�}�Ȗ%�by��59ı,N���'PlK��߸|ft�t����%�bX�}�ND�,K�=�Ȗ=�B��
P�� � U0"%pa�,���xu�<�tq:�bX�'���S�,K���=���i�u����%�#"}����Kı;��z8�D�,K��٩Ȗ%��Ͼ���Kı=�}�����,�ݒ���%�bX�y��'Q,Kľ}�jr%�bX���ND�,K�>�Ȗ%�b_'[��n���nMn���q��FLUk�5t�����[���n�i.���%�bX�Ͼ�ND�,K�}�Ȗ%�bu��4?N�dK���tq:�bX�'���_��4�ٗM��N�X�%���p��Kı:����bX�'}��G��%�b_>�59ı,N��{�ܻ�.k�n���%�bX���ND�,K������Kʄ2&D������bX�'�}�S�,K������̷L���K���%�by翺8�D�,K��٩Ȗ%�bw�59İ:�Ϸ������Kı:�l��].��2�7x�D�,K��٩Ȗ%�bw�59ı,N����"X�%�{�Ϸ��Kı>�i��!w$a���4�݂y:M���noZ���:�m�`3���e�^�
���Q,K���jr%�bX�y�ND�,K�ߟo��%�b_>�59ı,O|���7.�4�uı,N����"X�%�{��w��Kı/�}���bX�'~��S�?
�TȖ'����\�K�7d�q:�bX�%�߿o��%�b_>�59��*���<����bX�'~��Ȗ%�bu�g�dݹ���ܗwx�D�,K�����Kı:����bX�'^}�S�,K�ș���'Q,K��߹/�n�fl˦��'Q,K���jr%�bX~T����D�,K�翷��Kı/���ND�,K�`��<˙�һ�6m�t  7kT���vX�X(<V���V�j����`&hw[ �����{@��$�=r�W�鱹��v�K�Ayu�wPmS�1v���\m�3�݁9�R���-�ݶ�D7o`S���Z����o����Y���V�.և��v�R:�8����y1i˭��;"�$�h^�I�Jow{���i^G��,��k:��k�}n�mU՛�n�3b�X�-�(I�{ı,O�{�S�,KĽ����%�bX���f�"X�%�߾���Kı:�~��ܗL���]8�D�,K��o��%�b_~�59ı,N����"X�%��p��O�*dK��g���sf&�sw��Kı/߿f�"X�%�߾���Kı<��ND�,K�ߟo��%�b}��>�2f�i����q:�bX�'�}�S�,K��xjr%�bX����x�D�,K��٩Ȗ%�b{�=�&k4̺�Ӊ�Kı=����bX�%�=�'Q,Kľ��jr%�bX���ND�,K�w忯պ&mn{u@t��;*�H8������g��Yn�]aͻl���Lͤ�t�ı,K��߷��Kı/�}���bX�'~��@�Kı:����bX�'Xvy�7ni�w7%��'Q,Kľ}�jr��?zb��'q,M����bX�'^y�S�,KĽ�����%�bX�{�.|M݄�ٗM��N�X�%���p��Kı<����`ؖ%�>�'Q,Kľ��jr%�bX�w<�/Yvfm�f[�q:�bX�'~��S�,K������%�bX�Ͼ�ND�,K�}�Ȗ%�bu��fnK�.ݬ�q:�bX�'��ϧ��%�`�߾�ND�,K�<�Ȗ%�by��59ı,N��ލ��e�%2���q��/n��k��-9��ڱŻsHɮ���.M�����%�bX�߾�ND�,K�<�Ȗ%�by��59ı,O���'Q,K���d˛!�[�����%�bX���NEQ�,K���Ȗ%�b}��q:�bX�%��S�,K��y칒f�L˥�8�D�,K�>�Ȗ%�b{��q:�c ������ ��Ȗ%Ͼ�ND�,K���Ȗ%�by��}-�6-��]8�D�,F���~��Kı/�}���bX�'^y�S�,K��ϸjr%�bX�aߓ����n�n˛��%�bX�Ͼ�ND�,K�<�Ȗ%�bu��59ı,O��޸�D�,K�=����[u�lw-�?�[��G����Ѷ�{A�ju����ARs���wv3f]6�q;�bX�'�}�S�,K���xjr%�bX���޸�D�,K��٩Ȗ%�b{��ܽe73nS2�É�Kı=����(�`�'�y� �	=���$RD�}�lO�����y�fnK�nͬ�q:�bX�'�����%�b_~�59ı,N��"X�%��p��Kı<�l����v��sx�D�,�C"g߿f�"X�%�߾���Kı<��ND�,���S6&{�]N'Q,K����.�2����'Q,K���xjr%�bX�w�ND�,K�<糉�Kı/�}���bX�'���߯�둺�v��nЍ�8�v:�D6w8�=]���E��77��2L�i�t����%�b}����bX�'�y�g��%�b_}��Q2%�bw�59ı,O}�	pٲ��%Ӊ�Kı?{�>�N�X�%�}����Kı:����bX�'���S�,K�����3M���.��uı,K��f�"X�%�מp��Kı<����bX�'}���'Q,K���y~�7v3f]6�q:�bX�'}�S�,K��xjr%�bX���{x�D�,T[��٩Ȗ%�bw��ܽeٙ�i�n���%�bX���ND�,K���o��%�b_~�59ı,N����"X�%����������m��h  ѻXfL�8v�nJ\EeX�I��RpF��N����Чa,����YqjWi� 4��B��64ۧG<e�]�sBݼ���F���n~ہț�;��z�8��S=�!Z�-�s��{2y�pY�D^�m��@�W]��G��T;�N	l�O2�ֺ�X�nM�v=ݒ�cN�o�ǖ�m��YKs�r��ՓC�k+����^&���ĺt�ı,K�w����%�bX�߾�ND�,K�}ᨁȖ%�by��59ı,O>�<=.�]��7mݼN�X�%�}����Kı:����bX�'���S�,K������'�
eL�b~���wHi����q:�bX�'��p��Kı<����c�"D"dO<��^'Q,KĿ~����bX�'���e��i�t����%�b{����bX�'}��'Q,Kľ��jr%�bX�{�ND�,K��ω��l�nn���%�bX�y�}x�D�,K������%�bX���ND�,K��p��Kı<<��3��i-̴.vN^wfnxJ�Y�v���h)ï
�Ů�7E7LݼN�X�%�}����Kı:����bX�'���S�,K������%�bX�{��㹛2�3��Kı;����y:S�A^�K�,L��59ı,O}߽�N�X�%�}����O eL�by���eٙ�i�n���%�bX�{���"X�%��{﷉�Kı/���ND�,K�}�Ȗ%�bu�/ٻ.d�4%Ӊ�K�@,O<߾�N�X�%�}����Kı:����bX�'���S�,K��������eɻn��uı,K��f�"X�%�׾���Kı<����bX�'}���'Q,K���K~��f��eH��H�C������ݶ��nƮ{sW>�#{���w�}�wHnK7ws8�D�,K���Ȗ%�by߼59ı,N�߽�N�X�%�}����Kı=�}��0�f��K�q:�bX�'�}�S�,K������%�bX�߾�ND�,K�}��(%�bw�y�4�M�-��]8�D�,K�7���%�b_~�59�!ǂ� FH��D&�a�$ Q�%��.0�'0"],���,�J�aمq��,(�ױH4"�@!I!�$H _*s�^޻��k���H̵ �uk��s�p��P��&CXP�& y�'Aiz�=yB�1O'}�B|t�j�>�����'����T�� �x!��N�w�59ı,O����"X�%���=76f����&n�'Q,Kľ��jr%�bX�{�ND�,K���Ȗ%�'}���'Q,K���{�I�Cs6e�ng��%�bw��59ı,O;���"X�%��s���%�bX�߾�ND�,K��>�w��&a)��J]�%�2�Q�뛉��p�#Ճ�:I�+�t�)%���Z�ǻ���,O���S�,K��y��uı,K��C��dK���jr%�bX�{7ٟ�&�B��8�D�,K�?s���%�bX�߾�ND�,K�}�Ȗ%�by��59ı,O����wr]�.M۹���Kı/�}���bX�'^��S�,K��jr%�bX���=�N�X�%���N}2��!t�ww3��K��"y��F�"X�%��p��Kı;��=�N�X��h��Ȝ�߳S�,K�����0�5�\�fi��%�bX�����"X�%��~����%�bX�߾�ND�,K�}�Ȗ%�ow�?����\
�8�n¹�GW=n�&=v6��N+��<S����{}��oq��KϷ߯��%�b_~�59ı,N��"X�%��p��Kı:ÿ'���ܛ����m�uı,K��f�"X�%�׾p��Kı<����bX�'o��'Q,K����:�nf�m��uı,N����"X�%��~���Kı;�|��:�bX�%��S�,K���,��vf��r����%�bX���ND�,K�w�o��%�b_~�59ı,O{�"X�%�ߓ|ϳ$�2\Й���%�b{����uı,? 1Ͽ~�N�X�%������Kı<��ND�,K�7���A0(i"A��3�����I��  ����׮¶�X�.��6,�l�;պ�4suòƱ��g
��mɰ�����n�1��9�Ɠ���Tu�K��8xÈ�uۧ?�o�}�c��S�Ra�A��zmo��3g�µ�lbyi ���`�ER�e�m�Wn�ە�|�[�뜻9�b9�r�z���ӽ]�Z��'\�Ȧܛ����Gݞ59xӤC� ���5�����d,�ۻsoؖ%�b_�}���bX�'���S�,K���59ı,O3*�Dm�DB#/�LL6&m��'Q,K���xjr%�bX�y�ND�,K���s��Kı/�}���bX�'��ن���ܙ���%�bw��59ı,O3�}�'Q,ı/�}���bX�'�y�S�,K��<��l��Y�7$�8�D�,K��ﳉ�Kı/�}���bX�'�y�S�,K��jr%�bX�d�y>76e���3ws��Kı/�}���bX� ��ND�,K���Ȗ%�by�{�q:�bX�'����~-�vck�/!�`t� �k
]]9�&p���V���[p�r��nɻx�D�,K�}�Ȗ%�bw߼59ı,O3�}����ı>Ϲu9ı,N���z]����\��q:�bX�'�}�S��Q�P��=��ND�<�y�q:�bX�'��S�,K�F�*hY�f������V7��q:�bX�'���g��%�b}�}u9��F"}�59ı,O<��S�,K���O=���2\۷ws��K�,O���S�,K���8jr%�bX���ND�,K���s��Kı>��Ϧ\���I6���uı,O����"X�%��~���Kı<Ͻ�8�D�,K��߳��Kı)�����]�L̻��L���h�Ņ��fNľxf<ƛ�.�zg�{�/�3�7��Nn�:�bX�'�{�S�,K��=���uı,O��~��Agq2%�b~����bX�'����Y���r�4�uı,Os��g�~#�2%��?}�8�D�,K��jr%�bX�w�ND�DȖ'y'����̺[��f�q:�bX�'�����uı,O����"X�"���Q�!Ȝ����S�,K��>���uı,E�$7(9�1'.tF���D"3/F�"X�%�מp��Kı<�>�8�D�,K��߳��Kı=���Yf����.\�8�D�,K�﹩Ȗ%�b��{�q:�bX�'��g��%�b}��59ı,O�g~}!k���ល.|kӻ�)�H^��@�m[����,�l��f�K�%��s��%�bX�g߿g��%�b}���q:�bX�'�{�S�,KĽy�jr%�bX�g��d��kt͹sw8�D�,K��߳��[ı>����bX�%��3S�,K��<���uı,O��s�.�,�M�����%�bX�}�ND�,K�癩Ȗ%�by�}�q:�bX��w��6��D"!��!L�,Ħ�i��%�g�TbdL��S�,K��=���uĤK�{����%�``���zF)a M^*"&=D�>�Ȗ%�b{����.i��[�&���%�bX����N�X�%��y����%�bX�}�ND�,K���Ȗ%�b^�[�ݺ�^i5�s�[��B��ݟ��"N��YN�΋�Ȗɑ��.��陛�'q,K�����8�D�,K��Ȗ%�bwߜ59ı,O<�>�N�X�%�����Y�ܷd����%�bX�}�ND�,K���Ȗ%�by��q:�bX��ɬ��DB"�����&��2&f����%�bX�y�ND�,K��糉�K�@B9"~�~�'Q,K������bX�'�M�e�-ْ��8�D�,K�=����%�bX�g�}�N�X�%���p��K�?3"y���bX�'��{��7%��6�����%�bX��Ͼ�'Q,K��߸jr%�bX���ND�,K���Ӊ�Kı<��/���~��J`lݶ  [z��_�����l���]��(�C"9H��vG���g�-kd�F$�Y���Z`�OkX�)����mH�7<��mt�x�C��9){L�e�ne|����ȧ=\烶U-�86��H�Mr���'�t��rM:�k5�	"�`vn�k���H�[�m�;�}{�J����˼]k���{A�������ӎ*�ûh'	��Y�qq�k8�ı,K��>�Ȗ%�bwߜ59ı,O;���uı,O�Ͼ�'Q,K�����p��ܛ�4�uı,O<���!�G"dK�=�Ӊ�Kı?g��g��%�b}��59ı,O{�/�l��۹.�q:�bX�'�o�^'Q,KĽ�����%�bX�{�ND�,K���Ȗ%�btg���e�-��fm�uı,K��}�N�X�%���p��Kı;����bX̉�|����%�bX�}~�u����t�wx�D�,K�~�Ȗ%�bw߼59ı,O;�>�N�X�%�{�﷉�Kı>�~���]wc�ƶ�u�g�^�$���Μ��Zu\�\ι5�&y�yQ������{��7����59ı,O;�=�N�X�%�{�ﷃ�Kı>����bX�'�M�g����wc3N'Q,K�������	���ș�����Kı>����bX�'}��S�,K��<��K����r\���%�bX����q:�bX�'���S�,K��xjr%�bX�w�>�N�X�%����e˻��.f�:�bX�'���S�,K��xjr%�bX�w�>�N�X�%�߿}���%�bw��ϥ��ۗrf�N�X�%��p��K��<��{8�D�,K�~��'Q,K��߸jr�bX����������y�˞�ai�X֮����)j�-׋���E��m��8�D�,K�=�Ӊ�Kı;���uı,O�����`��e��A|�|��yHӨNH7�I���S�>�bX���ND�,K���Ȗ%�b}��q:�ؖ%�����Y�ܷm��'Q,K���xjr%�bX���ND���((T�D@�P�U��� ��؂�D�'�y�G��%�b_~���uı,O>��eٛ�p˗7'Q,K��ϸjr%�bX���N�X�%��g��~�'q,K�*�O���S�,K��پ��2]�.�fi��%�bX����'Q,KĽ�����%�bX���ND�,K����6%�bu���nf�.�.g�7'N�8��g<m۫�%[��ci4n-�i"��f]3nL͜N�X�%�{�﷉�Kı>����bX�'}��S�,K��9��uı,O����.]���ۻ���%�bX�{�NC�2&D�=����bX�'�{�Ӊ�Kı/~��x�D�,K���}.]	tݙ���%�b{��59ı,O;��'Q,KĽ�����%�bX�{�ND�,K���\�m�e����%�������%�bX��~�x�D�,K�~�Ȗ%��E��{P�D�}���Kı<3����vKst�6q:�bX�%���o��%�b}��59ı,O}�"X�%��9��y<��_��Yd��v3����7��ݻt�*���y`.�9��B�ޒWv�IW8�Is�v�H'������{}��nJ�:t�\s"�]�À���n�P����s��E�32i�����䪽�E �Ƞ�3N2�Q9MӇ 3۳�n�P��wsN��h�ԈPt��$��.��̞8��� �/��5J1(֬�,�W��t��o~1T�'�
�o��zP�P�D{`Ȍ�hS�7�L�@��K"B 	��!u �R!өA�{���s��U`�v�`.�I5E:�?o���H    $ ��"F� [��� m               ��m3Uju!��g�[���^͓͑��ke��U;U�� ���j�6�,����lK�T��*��'jM�����"V�C�r���8K�U8*�[�)rB�9�v�(�mW{lp�ҋT�v	��pML�S*r�)��n�r*�&�}��JVI���-Je��5\=��:9y�a��SM�,{�@nҺ�#;������1��ѵ�"�)#t�
} mɹVe�V��Bt-��7[ulk[���'
�������f�^��m��-7l�tdk�-���q�����y��3��ʭ�B�b��w6�`V�(�ʵl�����+�W֌-���;C�͛>�H�KUMԹ`��p��52@�/�g-� ��m*�v՚�L[���m���	�����S�g���Y�� �3>&�Gq��^/]�I�eAub�^�<�ZzMn�}�8�ݚ����6�j��`+P����Ac6��il4�p��I��q�mq.�t�	��J*�9v�-�<�Prqu���3���岭�Pr�Pm��-mٕ��;o+��V}�,�Xª�J�[3e���I�n��.h�"�����o+UUUʵ{ ���R��1m@UUT�!��I�J�&�Sqi�Lf��z
��(�^�1�C:i8��$�vˤ.!|�2�t�'3L����7դ�Y�v�Y�9����
=:����\�iݧ�ރj1%פ�O%�I�<nx��Y���.�- 6FU��ÚX :��Մ�rd&l�nɖ���M�f���?S�4���">���낏�X'���`m�B$� '8��t�@�����m� �nn7�-�r�G,.x'���7W`ݢ��o�������kP�VkQ��9u�$���v�oc�Ul�F@�q3�<m��lډ�1���vb�
�OZΛv糵��e�c��=��糹)ŀ6�V�9CiU0�nx�\��hm�:�<�z�lHqv6Vn���"��oW�t���2��&M�t�v�P�UKa��s���5fB4~;�1���k�:3w��lP��p?n���@/�]`EN)Ua"��4�n�������&WX���L4�%�-i$����J��k��I���J��-$���N'�8:�ԓ�n�P��wsN f����ʎ5$�ӧN5�72(���i���=�����P������.��x����nv��ouY��v����ΎQ6ʃ�>�Qp̞8��8�� �^�3N2�Q9MӇ ;����T�Ij��q���v�]����%�UG��:�
2�)�8����ws� ;���v�_%SN��FJ\��]�À���7v(���%�F8Hp̚p��8�� �^�e��AU��*�c�9q��"�m�z^��a�g6��o/d7kδt�>����3�u��?.�^��pߗ�rRr|7Q:�pǤ��_U����� .���e��I*4�P�פ�s��W�}�{Ӏn���*6ʃ�>���{��f= Ǆk�S��TNSt�����?|���<p���s� �&����kj��/ı;���	���j�5s�1�)�D(�$�I�3���˹� 2�g �����QD�8��{�Q�ɧ 7=��3���Y���%D�8s&� �ݜ1�V�IlF��M��b!�KZK �b.��Ws���sI�$ "I%
AD�w�����{���fφ��)�-� μ ��. e���i����c�P|�9 
�^�)di9#��q-��eV�� LL�D�,[�����/3��{��e� �Y�7EAӉ����|���zp���x@=Ytb)�*"�RG 2�g �zC���V���n�pf�A�D(�R7$�oHu���. e�����t�|UE��oH33���ZI��Q&�V� 
 6S�Ԯ�hm�Z�`  t湴u8��5�e��Iҩz�WL��A\����$�=N'�

wjV��>����r��6x�Qg����� �����ȝv��f���y�kt��,�W.ƍTMmY�I��<9��0p�֎:�Fq���x(�-awn;q�q���U����6-�n��_�{��{���|_m��)�Onr��\l��ƻXn��r���:.�t⒤�!*����^������u��ʱ<^В�(���7 7=��;oHu� ��qpś�L��S�nN�z@9�6�{��w3NG"�T��P�פ�������{�^��[��*S�>���p�vp���x@/mULQ)��*�"��������gvϩ�ƒ�!Րc�N5J�T�����BH�w�8q� �< �� ��j#B�ubKI>y
;B���6m�(���F�M������U7S�(�� � �g�ջ��/_�VZx�8��%I*��;~�.����w�[��][�%:QUIG ����?^����s��.�g��*:���uN��k�l�Y�Qa��4��KЄJ�g^����$I�|��rݐws��v�՛��/7�#�G*Rtܨp����qp��|��e�̄aR�9�8p��I=���rx|+�t�r��b��ӏ��x@=Yu����T$��z�5����v@9��.���t�4(�I �= �d����W���u�
��:j�E}@;f�;vevd���`^������hB�'\��m���@9��.�y�ݠ�~ Y��ۊJ�	T8o���6�5���޻ UոPȪ�����m^��Ǥ�v@9��.��_)��J���Ǥ�v@9��.K�ϒG�% )*� =�=�rI�~{��vc�):nT8m� �s8����z@<��%]ͪ�T�蠩�t1���^f@C�A�����h�еsf��4#{fߍ����� ڼ��;�H:�me�P7���P�.�y��w�u� �w8���Ө��L�9 �= ���qp��|�u>�TJ�"n���s��\j�_���x�mf3Sn)
���C�v��\j�_ �= ��ߒ��Y��H�!L��  �w��\�2]g���*�����5���v��OS$.����A����Hy���N��%Kg@q�]M8_\xݜ�z��j2��� 6�㎞W�#ع9v�
�;qT���ғe�&�v�9Mph�����;u�u��t�jv�Wo}�tk,gOG��
q��e�!�w�%����[�XV!���_�k��BEb�M�:v����l�H�8�W���;�H:�s��\u�#O�T�%��Ǥ�v@9��.�y��v�]q��)R��2�(;���6�u����<�Q��:s�U ���p��|����Wy� �nV�7����pU��z@;ۊ��qp/|����נ��!ú��]�rv7��n��AV�1�k�@��f�I�#�G`g�`s���\P��>���W���D�8�E+~�䖦
2 �H��b�6w�^����_ �='����j��ԃr6����6�u�����P��R�2*�"#��m^��Ǥ����� �F�*4���'(�>�z@;ۊ��qp��| ̭���DU ko�|����s۬�th�s<CYY�lј�9�P�7*�"�s��\j�_ �= ����A�>�E�;{�\k7_ �= ����Y@�n�"�$��m�3I>y
/`n� @��� X T�{�Bc ���)���#8p�/�i =H�G���B,�@^������L�R$� �`E��������(f�G<d�a�Ҁ�6u�d�fc;	g��.4|�K$���߂a��#B,Rh�Q� �*��lF#t'�Uˏ@tu��pp5�X�IR"ؐ$����4"����@8��z�fF·�'�׀�0�X��@�D��`��=O"�8��J�dH��� �0G�=D>���s�E��P���x�@S=y�A�'��|�t�'���I&�S�Q�D���?}���y�@9�g �f�����C��Dn&��/2(;���6�u��� s*��M�3�Q��i�3���=���e��B�j��{\�dd��:�	%F�ow�����w�ˊ�][����Ȉ���I>y
$��'}��U �����U�S��)NNz�@/.(;���������II�r��3r(�y�I'~{��O�;�@�P!!$��BA`D$��BABG�T$YHDI`�b�# X�T�B(E�� A"H#���\��l�β�\m���� ��x�y�8q� �����(ܪU �_6&�(�z�'<m��ݍ ��rMr��Yם&&ˢ�ͯ��|y�8q� �����. m��:u�b���vޓ�$��܊�f�p���y%�J��l<�'S��MÀo�(2�]g���Z}��O�P8���f��w�����놼���>�N.� ��&�u�^~hl����N�����~��z���-� ��H�y�#���vn��I�&F͜�X�6W7�wѹ-^�/'M��'$����X�1q�
q��Cu��O���ݲ7X�s����1�v�J�ݻ]-��r�rPqv6���|b̖A6,��.֎���@7�t�ŧ.��\��,l$�I��r����� ޺���l���]�n����m��w�%�I�]�۱\��4�X�ז�PC�K��;��?������C'4yɣ�̵�j�%c/1Z5Ӣ��;�M놵�o-f%�3#kG���G��?4:_a^$���i�rh�\5���h��A����2µ�h�\5���h�D$�r�K�ݹ�ۣ�%��@���2�nx�Mn���Gb�\� Vb��N�k��94{��|1���ɛ����{�q=��� �� x�t{��������p�w�r����C|�Gz�~�큖�D8�����Z;����ǌ׼���\Xm�+y�Ѯ�kx�{�M�|���tl���61u����U��tv�K�g����nRG`����i�QJ��~�z��sw����̃��k��tPE,J��rh�k��/����A����rµ�h�\5�muS��t  �B���5����.�]�E^3��k�f��&�u�[φ0sYv�I,�� >��9�ƽ����=���]����D�˝�6x���g4�tν6�u{��@�g
x�W��G��o46s@Fɘ�*�-YXRZ=�k��h�9��^L+,b�c/1Z5�k�|���k�z��Y��h�G����:��:H�F"���
7�4��q�8�]J��sG��͡��%���U�}��	� �H�);;&���	q:�dWMq�\��T���i���b��nu^W���߹�74F�Y�j�W��j9�� ����p�U@�n��Ae� �]��� ���w��C��w��g��H+�����i�hl怐Gb�Wg+
KG��͡���sC�B�C��{h��-� ��u�"�LS:��ٮ�8��7f�lDc9.�ܞb.x6e��=��í�\�uԄlE���qu*�v'Y�w�b��u�#n�w,,�������:ݳ�Q�a��vs؁k��k�*��lWB��;J�a����3������ԃFm���u�.���=����������_ ���J�
Ca*�d�g��I;����Ɲ���X�s1ȱo?���~��7��u�^���
�(��@�Z=@>nh�\4��8K�Ŋ蠊V���=�y���4��,��XB9a��y�5������<�w�1R*𡘍t��h��;�� 
�Lu���M�v����{X�(1p��u�vӊ�秵:#"m�%T����y�D��7��Zy|+�!������� V ;��r�`P=Z��Q���D +(�!I�@��ݾǜ��9׾ |��V��-XV-w>m�h���,��,V2��QȆ����;����;+0���qh�H�|�՗Z}��v�S�B��(NL�T��.z]�qYx�w\@�&&���d���e�' ��~��4>�i�hoF���ŗw�EXAbZ\4��Ѡ94H��x2���6>��s�<֋��J(�|�f��os��f ���%v�yȀ|����͡��t��āX�|����͡����"��Bc2�a�/v��
�N�i�p�h���"V豎�^�uuh�C놟6��h���,��,V2�+F������\5�'��Yd%�г�G�����|����+0�6�	%]]��b5ʦ(@4��I]{bW����%(�s�.��͡��sB>n-Y9d��������0�yݼ	�7l�4�`P�y^�l��y.��Xq��͠7>���5��0fb	^bI]�d?Q�����O�C���E%b�� RF�94>�i��7�3M��
�1aIh�i��7���M蹸M5.\	����/��b9y������L��9!!$EDe����"?��ģ������QD9����^�ݟݴ燚 ��C�H��@���AE	|� H��=AD�(�EPREJ���0�������#���6��q��W��#Η׭�@����$~�ģ�	��C�w�G����?���'����ED�!��#���(���������i�Y��}��~ğ��@ �������ȍ  ��O��D��??x{��{��w܏�.��C"W���{�E�!L��(�  ����H "��"�",B(�F�Q�"�"*",A", b��P ��Ab��  ��P�"�X�, �� ",D�,@",F(��! �F�b��A�"Ă"�"�� �DB��, ��
� ��� �H 
H*����U�AP�P��B+E�$�W�����������Z�3��������Ǒ�G����}X���@g��=M���@�>!�C�
���<�� I>��"�`~ }������X_OP�@�����'����������=?_��? >�~�@�_��_eV��G�!� �@ ��>`��Y��zh}�TA	~������F��PDv8�(?��PDka�R��Nl��hq1�k
��/��QD����|�~_���GH_��������D~c�!{x�_�T������O��A����?��E|�����>���?���x#� l�@G������?0}��u��?/Q��:A �A�tH�.{Ǐ
;���{�y����>��?�X* �����n?��%�G��A��2�H���4�n��g�_�>AHr���]��BB�'��