BZh91AY&SYР��߀px���� ����au�    ݀Pɀ�� 픶�l�Q*�CtnնY��b�[i@��%�[�!��f J� ��@P�E �"�Q ��R�*E*�*�@*��I�		JHJ��BI"���B		�    ;�  �      
w����}�W�Ol�=��[�� }�>� �6q:���C������� U��QVf�Ta�(3��YaT�J%LMR�6�R� �)[�ȥSBU14�)���         �@n��\�����wW���j盼�}yW���z���:�������ҫ�c�}�C�
���k����rw�nM*� -S��o}�R��u���W�ϷR�:�:U�U}�����qeS��@��      �ޕ7n������֜����3^��>�׭��ە����wJ���Mv�� >�=_mŽ��6\ :7WW-�Ԯw� <��]�w�m�����|/x���� �U��ԫv��7m�YE��      
 >� ���s�޴�6���ӛ�iu� 8��n�4���Zy�qjS >��Cvz��Z��纜��]� �w��.�msk����_n�=R�} �T��\�-w���nU���+�z�T     �� |����e9o\Y]9:�� f�n.�NYzӾ�}����+� }�zRǺ�\�_  �מM/˽�k��s�,[�K�=j�����w�V�� �7o}�+����}ϖ]z�>�{j�         �Rbl�*�@     ��қ*T�0 �    �z�R��Li��0`���R��J &h� LLѓ U?�2C)J���    )	T�&#Q��O
m4dфdɩ�z���'���w��������8{{}�^��QEW��7xEQU�( ��Ш���EW �T?�*(���ʱQU��S�s�QU��ͧ��`�����a?���d�P�`�`���'�'!B������{ ��v^��{	��a{*�(C��������;"v��G����	�@��C����a�=��`;!�{��`N�eC�v���vU{=��;
���G�/d��^�'g����;`C�e{ vT싒&Hd��; �E�e���/`N����{!��d^ȝ�;�� v;�C��a��N�n��w+�½��e;��v�a�'a^��C���C�&@ �^��;
����C�a{ v��G����!�^��D�e^��{vG��콀;!�A��܁�Sr��)���@�vN�v�vN�v�d; v@{C���;g����=��v^���vT�d���v��e�����v�vN�v�e�d;�����v��S��W�=�콅��❁�/!�%9���;'a�`�n���vN���v���a�e;'`�=��=�;!�^�v;"����l���}z�p�4�A�'C����q��fi6��|'n�8��p��N�MҥeD�_�g;Ĩ���d������[i��n]+��+��G���>8e�3D�{0�8�0�oF�������{�������A���.�%���!,L~Z��ZѦѻv�Vm�h5�5a�'	��K��ؾ��V�9�����Y�i�Y�4��f�y��Q�	��r�Ife1��q���;���s�j3_�Y����mׁ�����300r�Չ�D��b�>>�w0���M<�~�<�4�G�w�6f� �F���C4yo|>�<���I� 2tF�O ���|іgЊ7P�čF��k<5&��������H�is�)��S���	HQ)
�A�I��c�!�R�(�M�_'����3va�D�~|�0��v$FF%Y�%��ɫ5�tl7<u�g�h��/)/=�.��$���_SB�d�DR��@"Ns| &j抩'��W��[cD��DII��ʼS�O��h�I�w�yeΥd�\/n_��P�i}�i[1e̪�Eћ�5�b�)X���b����R�T�r ��*�(��Y9����ؾat�ѢNc�-?t��LTЁ3������}�[��#F��3����	BX8�-N&�	�*����I^f)�
Jc����'20�Q��@Z�"rp4�Ltj0� �AK��Ya�,u���`�#RN��Fi�35��-eǎn�����e������{)���'�۞o��7q�Tµ�?o��~Iʤ�*M
U	�k�0KU�F�'6pu<5�a�$'v:�3�p���s_9�������'9��vn2m�������Z�!�a�3g(.ZcF���A�>��@>1�S�&2� ��d`�����6kFiud�rq��2LL�̌�7��A�X��v0ߺ��Q���q�ӻi]Rb�bj��&��W^ش)��d}�BXB��Fh��F3L�ύ��̌��oa��-Ԛ�8��㓔��c"�)*�"P-RzV�QGǖ?��[f��'��2=�����%Y�b饗Q���0֊H`��5}�\� ���n-�Q�L4�D��R�-4!��s���<���ߛ���_���c82da������w��}4ו�\�j�9UB����5��E��<L��v]FK�sN�x�l�a�{�4���l�,X���I�$9�Fo� ��x�9�$h��4l�d�ۻ.�
K&f	I�d%PE�F�f�B�MD���BL�D�.�)2ɫ.T�!P�b���)[����SIP�>^�B�ϖ�������T�
0j�)A�5���\O8�S�*v�*_�bO�)@���Z�WQ���e���)ɱyq�&�5`�Ӻ�#(�p58�#5�Wh���N�s
�sFfF�� ����������oN�A�H�J��~��Ρ��+WV�J�Sd| 䖲!� ��A����k��43Q�2q����A�������tq��9o��}�cc��D�$S
J��t�,2�o�b�/�J�j=m4��0�$ڿ{��������7�<� ������6s�ym}�r���
R����N��q�1��,�\rg,frc3~��a�Qǉ��t�\q��2�e��s�95���5�6Q��%��Y�a�5��Qool�5�W�&FVoq����Ͼ�F�������y���ĵ��M+����V)���MeaH�DH�?,��XOڂf"VQ�T4�dT�*'Nf0���2�k0cZٛ>G7ș�i�k{�Bd%���8�"�H_�J�բ�,�,���~U���{��'��(�JW������]@�vtwj��W�ԇWm�~V!�i1Σ���`�B�P��D�WʖR�����s�����v��%�D�� ��W����;�8�AD�Gꦔ�Zr3�J�`�i7e:O�qݹ���}����a���=�;QLkQ���h�Y�ى��Y�F�#�-��N0�N���aM�2��h�f:ĝƂ4sX�Q ��Hbj�M+*D�*q\)�jf)4��!�d��D}䤚�k�u�V�(>�f�,b�Մb�S2�;h�)�R��W�tn')J��f�#V&��k����5��`���r�	���ή��Jr�|�*��pj�=JU��:��f��yU$�z��@����S���t�or��F�p.g�=��h�a���6�-�$D���hw~�j�?/������噸�W'�+*H\+WMD+1RA��!6����Kb��Q]"���r9�p��Lj����yn��_}�D�G�������H�zU�b��!"z�>'��*&���@����$Д��VЦ*jd�{�&��W��R��2�����BHV/$B�;��
���b����?Z>r.�]������Up�:�I�!�[�H���1`1�I��G����aA����Մ���&�B�ʚ>���+Y�D��LE]�:��fQ3j�Ū�I��;iN}
<��k�}T��ĥJ� P/�V�x:l�sfe.��̃>�YxZ4EQƬ�l��Č�",��2�-�5|��*q�ec`Xj´�ݴ���IZ��Ī�(��?1[���'B�ʹ�sw�qջ�����R'3w�&7�<T;�>�_K�{�J�i��iU8�ұ2�i���+�
�$DW�)U2	���=��T ^���LL�Ԛ�#�� 0�L�T��n�"JI���+*�#����R~���ԣ9ƛ(���X`��%�Jrq�Q�01	I
a�B_J��JiL�������I�k���oz*4j�V�BP�d�f���M���į#�w���;�C��=h�󴤘�@��)#	b�XDO�`j��2���v�0�##>fQA�u8I��1���%Aa���\����U�_u��4��[4y��V�1>Y�z�F�^F�4R�	4'G�c��>oP�33)َX�o���4�1�ſ���0�h!����,�a�AXn# Ĺ&��
uA;̉%� &�i��a�6����x��ێF��n�oxXs$��LA�,g���Q����՜�~s+F��@a���1�d�8�b?@>NUr\��,!�S�	KE�6DF6,�|�f�q���Y�-�CP��d�A���p��3�I�rLQ��y�c������(�b��%��`+�BP��d�%	Bj�ߚ����qߑ������5͉i�LF��j4bT�BPRn��7�CY��13xMA�9�kw(0���-�(6~��mGx�����y���L�����h�5\ɀ�IȈ0�LL��L�4�bԒ)�P��4�Of�~����[z�1"������&HS
E(�,|l(5!��0r���e�����l��<�:6��<�	�"%��
~�ۖ��ܥ�m��#�Q�*�-����V�������E4>�K��	�IA���^l'4l'<�4NX�,H<�g��#9b�2*"ID	IEi�>��+'�k78D[�0>O!�t.݈d�'�������s9����|�-����a B��B�;B�͌��Fg�<���͎pMN��yE!���M+(T��鿱b!D��g$�n�
�G�����I#*��
攧�J�z|�T,��R��
��ɫ' �0���2�池�.�����<d�c���tv;FfzTai�Ŏ`��l��*7�Z�VVL�a�a�[�EA�jp'X��P�����R�����j$�,)3�y�f�������
3̘�Z��3|Ĉ�Sr0",���0�m��f��2�e�>pv�>��эz��l�3�bj$7j�����3|l�Vy9%ç����� �a虄�A��FX�1543r��'[y5�5�Vl7��'
��H9:u&���|�VZ�<�ӲCZ���bQp��0}�-��M[��f�(5j4@W���4eNYbDe�a���|d��"')�I��d��M���y�)#�ĭ�1e���9�B�ȕB����i����ۅNW����/ؠg�4T��R�^k ����X��J���2&��$a�w���-Zf7��Q3>3����a��j�ѕ�ȉ��Q`�3$R�II,G�d��R�`��' 2�4ܻ��ø���<aݜwon�|���yǛ�M��h,�c�u�58�<�=��;s��n��^p�9����.I��h�l4I�sAf�Y�۫~ZEr��W���:����\+���������)�Ӆ,SB	T)�UJe��.�.�Oʩ�H]�#�����Z�*~�	Wn�r��~�����U�	��$�U�)�����@\�}ggN$~B
�ya��1����4r1��ko�]:�|�
��$v����P�9R)��^=�E�MTҘ O�"_�>'1�"}�ϭ+��4Qi�smZ&��τ�o�=���.�<��,�(J��)4N���Ԟ����|h��0���!�	v�40'b���M��0�#��_���ѳ{<�1�%�I���)@�nLL���d㦬C'���N��5l5P���9	N.c��'3 ј8�$%*V��W/7g5�k|�����0��P�rLMBX��A�g'8�Z�0M�`c��2Y9E��G�[��xoSM�C �q����_�U���7���W9)̯�C��1/z�5CV)�$S�r�7�2������U������0�aT�eU� ���,��"�Я��B%L)&;���,R�w+�K���6.~��,pU��>(߉�NU(eR�����$R������a�u��Y��c�S�1�bDd�I)��(�������R��P�&>p��A�R�r������o6�BQ�	A��DjtI��!���4�:H�rw���j�y6�Q�:�	c<��@a͹I���'���C����A�'�b0J|��0��s�F|>޷�Dg-� �	��<o���i�Z�b5��>A��Ձ�3Pf���ԚL�����ӽ�0�̎F�)Iy:�ZѬ����:+Fn��F�7�{mh���yx퓹ͽ+s�':��7!f��k��=�6ӭ�do^{s��{s�v�k=��a:k\���d%[�b4�a����	��Q�o����N~�M��h�$烢�l��m5L�c U@mUUF���v�N��'b޲�� -� �a� 6֢�l�m�9� 5� k[@  l     u���Zmmd]��/[Ue�h�  �kj�mH"Z7m� 	�YY��       6� *��&�c\�x`.���u�Ăڰm�m[� I���     m�a&[[kn �m�p�֊K:�  ��`6�3�=`8�l�����h׮�֛lʲ��e��@��P*��Pp5�T Hn��Y��@pm�m9m �� M��l'[Am^S>}�Mmh�ޣe�V�몪ܱ9A�{u,�-uUP�ҧ=lW!ێD������i��n
ݞ�DE�3n�  m���e�%����ڀ�V��m�m m,�$��p���զ� $ �m� ��9�k*�U|r��m �[[_vG�$�e(  m�lH9�[vݎ 6���6�� �)�  z��5��a�  lԒ`'"�^��m�gI����j�[�ٯhm�l�mD��V�-��b�]*�Rjڳ����BjVR0 �c�p�ҭa� 爪�8�y��X�$Wça����lmU7hඪ�YZU��Ry����;��K�A��2�eT❈��zR	�Z@�K��U	��@U ��T�T�%��Wl۷G���_mǎ�l�[2�p$�Q�Gk5�f�0��ZY���G�"��m�Xgic6u��Vʵu!�\�W蝱 [A�H%�M����A��؝T����H��U ��@Yۦ�R�5Ҽ��}�Ҭ��g5\�R�]]T�Sn�� j��Ά�t�miD��YT{k@��z�	mm�$ �`6��	&�[ �I��mU��,�ymIf�V�I��oHjm����Bj�b�a���g��j�#T%uV������<q�6v�Wd{X8t�%#֎�J������BJ�v�b�cql$[\5��	��Rkd��v��1L�n�����4�C��(�]N%���F��+R�1�+�k���>��r��@uy��s��P8��ḏE����	AsM|�;`GI��	$x��a�A�JK*�bS�
�
A�e��js�(nz�i�fTN�-�+sg����N��鬢:�hv�7�GmЛ���lOc
մ&��V, s�h�T���<�g���G������LM� myoZ��:�oSh�4.֩�a����@A8��,*���$����Wl��P.��N`�r�ʹ
����<vENZU�%���uz��]�65/\n7H}+F�j�Q�r�U&���qaM�!4�դZU�.���)y��� �R�&F�[\� K(�ݝ��6\���td�:}59f����v�ӏ\8 m�M#%+�$6�m �8 m&�#��ڤ�UYZl��UIX ��E�l�[A�մ�FMU�v�zN��L�nҤ� �-TU\ 8�[�-�Kͩ"�����E��u�����2��[F6Ԅ�*�k	9��%�6�m 3J��i[j�]�T�6���۶�:���t�  m� ��� �*��T
0��~%����j�i���j���vG1��6�ו;,��+KW>6�n�;j��,�[@[A��a'@ �   ���-��M��m[@m�� kV�&��"N 3�����m� 6�'$��f�C�4Y�2zT�VۦvF�r��l���M����l�u[C�4v�Ă@m$�m��`B�L�p  	��$��lŴ/Z��ݚ���;��A�n+���nf[m�m��  ��m�����,0'ej�^\�6ʶ;
�WV���6�@$M�Vk��
iM״P<T��e�Aղi6Ը�l� m���KN�h�-�sd�i��ջ�mZ� kn	wK�C 6ۋz�P-��m�6��d6���m�@t��shn��[�Hqb]'f�m�� $l m��LVН��!J΍��j��,R�l�m�B@m�Xy����޷<Ƹm��2/Y��K�c��0�Iӝ7$K�m I �� �Hn�H �  6�    l��	;E&����Ӏ�n�j�lt��Z`� �un��R�^����Q*ҭUUJ������q�U\�P�fQ���U�  �6ͥ�2ۖ���UU�x6�W��Ŕ�^�������2/�Vی�is��S�k��Q4�[:P��f���     	���-��kn�&6� �@m�m�l'�)m�VhkI ���HH�o[��
T�h 8n՛e�,��E�u�Ժf�UV�BL��U����v$ �j�G��8���V�N��m+̹NT�-�k����� �$������@`� Z�	�$���Z� Pݳ��7S�U,jxAa������,sa�5��*51��vx����(6�	���ѓ^-Ö��XI���nUU��T��4@n�U��:���M���&�	0bꪒtK6��k	��4O4��z�Q�t���j�t��;<��u�[I��  m� [Kim  n�8&�p  ���}�  UUUR�R��j� /r��UUV;m<�ҭ*��T�`���{P�yEy��hV��4���m���Cm�Z��ͪ���,���S�s@����e��n��{�}EZ��j�U�&�-�����_ }u�.ָԔ+EɳK��U8)V�C�٨ Z��P
�0r��K��Z�y�Q�k����-��6ؐ   8[A[���A9׵�uR��T����v+��0�(v]�P9�]n�0�ګi\n+WX�+/4�8��K}���ݾ�)�-M��Xt�[���n�M���mÁ��Ku׭��e�J��ه�{u�8�3S���j%�v��.�lu�^��ۘ�u�:4�E�Q�{p�UʱJjn;6 b0��=0��na��0���w���b�#9�k(�n��.+��Va1�b�I-��-�^�l�����@�N��9x�A÷m���a���+�Q�^Iuu��Ha�(�ۖ�Z�Z��4�WU +m�Iu;ʪ0�v��6 I4�M�	 ��7k�[@ Hڶ�j�U��y�Yy��j��v!�.�^iy�N�lJ+J]�����ݺ����'�����U���ʺ-ksi�v鱶Ĳ�z�-�$p��$rګR�U*�@*�m]u��i7:E!��m"��]���k��D]����v�؝����- p� �e���u���궪�g(�g���sHHe�D��۠�u��6�-�m��l86�@  u��s[v�i#N�U�  �lv�]��  m��[@$ �J�` ��  [F��m��uMYh ��+`  ��qi[����`3fPݷ`�Nض�z�dH �Nm���$Im�E�mm� ����.  �m  [UX�Q�,h�iyRAur��U��j�mYV&��n`��m � m�p6�kl�4�#�-�m@�i� ��ʖkobE(�w��[U�9�p�[jB�	�yi
v@j 6س��@ㆵ��!� h� *���
J�
� 5u+�5tٲڶcR�T�\Z6ؒ@[@�.���vn�b�6� �u�E�R�*���p�c���*4�Ү�HF�;s�TUn'8*���Z�V����I��$8$�9I�T�=n�j��
�5<��x�В��+���n�f�ɛ`�/JD�@Ĵ��)g,9٨�ȶs� h+Em<�N�ݯ/;�ʫ��X\�'d�1��V���!���KJ\�q+V�����i��q6䋊�n;.N9'n9ol 5�1@�A�ڏZ�jkph�u��yoK�Y���  ���<� ����+I�����b�Y�$ ���UV��;���G�U����x�M�T/\):ι�x�<��F���Z�Ÿh�u�e��tۧ@]%d�����j騐6�mW@�Ky/Md6���Qm�me� ��	z˭ε��M.�͆����˪�v�Y��^��p.��mf�   �b��a�}��� �յU*��s��V�t�lP�luR��L�UP�0R��R�Y��mժj��ڔ�����],R6ڀ�ܶ��m�u�.�Y���l�� �i��f��Ӟ�i*��k]�ɯ+]2�n�Y�#�ukM&X��`:^t�R�UU���56��8W�MW[r�P�'*�n�[m��m�  	 !�6U�m�:[���nm� E՚���m՛�E�ʮ����Mr�UJ��T��=]kY����-ӳ� �)�̛b]�J ��Ln�6��� �cmm�H@H-�8M� �  ,���`#�In�
m�i4�P#-u+��5]Hv��/[��6ݜ]*E�6@,����
��S��eܨ����Uv��������D�\�p��)�z(uا���S�'T�6�¹8,�Ry�ؙ�Ɉ��j�MK����i���)^Z��^�������Q�AX���c���<��<������w� ��� ��@����a� ��)((��M�A0`d�`eY99�$F�Fa���!�L�4_�{��Ax��?�mUUEUQUTUUUEUQUTUUUEUQUTUUUMU�UU�U@5UB�UUEUQUTk�����
�Q��a?�����E�q�T?B2.����L4	�����]��4!�'���t��� ��;S� �)�8x��U�JE0@<@�>��B�S�N.��8J�$�D!�U^"�����}1E>#��;�p �>�= }@Sˀ���x��}��U� z�P�D�}��F< �ͣ�C� �	#�O��4/�CK��|�� � ���V6�!�I�(�Ht��C��D1W�Sb�
 ޯ k�>�����H&��ͺ��}���S"FM+� ���J�����~�}`��D$�$П@�+��@�G�O�	�U�E>& �@*f�� � ����/����J��"|�}=�}��?T�=���E.mD1��(_ ��J'�4.*A8@�����`�����/߿~K�%��m��M��m6�m��ʼ�ʼ�ʼ�ʼ�ʼ�ʼ�ʼ�ʼ�ʼ�ʴ�i� @��� ��k���M�F��ִ~����U�����_����濂��������V�+3+5����t��*4'�ESQA(�MPPR�QTRPSHSIDAMU������4d&0%*A@QU�P�"dM-,DRʶea���	R�AHT+���LU�bҎc�����(
T���5
�(�"%J�e�Q@�KH�I@K�d�H�aF�arDK0�	�(����2G�e��N�e�*=�7�:�,��wq�޽�Gy��i�Vv�e`�Uyj���2���<�UUUL�!�܄ Un�:Y"�L�Z�Aő�)NjCH�����q�m�3jv�:�uZvf��D�O\��l)c+J�u�T�(�)O%'�+ �;qq���(Ⱥ��tk�:�*3̇A-�26wm����:Y�L�����JY�FT���Y��ضi�-�Aጛ�5��ӭ��!t�\E�k�]q
�2�5�Z]浈n57;p`��'DWxu�4�{��/e���8N�m��&��sW3�C��3��/mi�BUFq�-���p�=�x2�m���.]ؕu�	<d���Q=���\UT�O,�Ö�>_$s�k��j�� �����V�e�^tZi�n�4�ji6&w4����n7\* ��ڊ����a�5��v�%G+��+�l��$�tfn��u(	��v�O��(Ȧ��j	�۶@\7��"s,j9�Y��٧v���X+!9‪ �<,�tRհ`�R<���V`*&�줃��u�1h��NGXع�p���f�`--:L⡙7	&7Hi�����4���h���!զ�l"�ьv�(�s��`em��r�.(k��Ӵ;DK��cM��@�c��
���i��<��.�����i�����M^t����t�(G��"��XI6(���Lm��-� F�6!�]I���b��m�U[`�Ba�nt8��y�"��'`�*�ڰ�M��� ��de�A���Uhkg�R�ⶊ�ΉF���+��u�H�.Y�kf➰l"J�\�۴��Fe�Iٛj�2]�l�[.���w] =ZK�*Ӹ�92�]��0H҇;c��\�.h"]���n�W�z�(٫p	�+�Gw'ҝ�5γ+ì���u��N�V�!����N܃�$��P�c���>��c<p8[,��ҺH��T eZ�u��m�(XZ������H�(��σ�㳻Xs�:�=�&a��O�4	�� �����(�O�%�����4�AC�����~�1?Qd��-u��ک��^��e�M=��^�\P�n;s��-tb(��J��{l�y�vsʹ+�H����<��#�e�C�� $B}B�n��Xv2�'�%<�];1�Wܘ4-�i��vav-�-�=8����T+v���6����\��x�Y�1P ��̜l4��n�]�Pv&%�g �x�Ywe�5=cZ��l�Y�>�(��y�Uj�4a��<��˄�q�6{pN������좋�a���AC�Ʌ�;�����z?�-��,����˙*FЊl�71�`�d�3=0�G{酁���R�Rc�ND:m��>��7q�h{��L%�s��U\Q��%�%������:ٰ7q�`�5���Q�ӊm
:*8�u]�3� �s%��Y�`�Q�(�(��sC����n��Y:�����-��^� W@N'�U�u΀�K�Ω�#��&آm�p����u��N��c�;�L,�{"p�Q:J5���kg*���窇�*x!���.�Ș�.>���\�.%6I\!�S�ITR
���$�%�3�0�Gk��gB����V���a�����-��
�r楶X>ݫ{smX��w鞅�;k
��9UR�tH�*G`s۶��n��ǥ���mX�G�f�j��I�"�s�\�nw��6�ǖ�b,g�9e涍��J�۱Q���9cv�� �w;7��ٵ~�3u�`s�����i�T�JNK���`w��6����f�P�N�R��e�T���t��[�`f���DD/DBJH$d DLR���{�U����2�Y�r8�1D�Sq��L,�f�7�ُKgۭM5*e���9�e�}����ݺ,��f�3�=0� ����Q(�EJ�P�1�&�
g�����F�S����¢��'�����J�"�qȪI`{=0�9�L,g���%�3��܃nA�n�Jq�XA��"�L��e�w[�V�,�����(r2J��L�6X��E�}��g%2���`{5�`nc�%�:US5CKm���]��ץ�O���^��/�+��Z�9��U[�8��\��7��`f�"��W������~�M���v\t-Ѽ�AD�`^H�pr�]�g�s�7�xz�8.��n��Q`f�"���q`����FH�t�%Q�V�9
�6(���,�^��V�f�=�K@}��6�eh�	Q���B�V�{%����ͪ�<ڰ=���y{.�pLr �N9*I`�>���`	'VV��IU������$t�T�RB�;�d�'s����f��f�tJ!@��BP�D
j���@A�Y_��A�}�.{u�:0d.�U��z8�	gg��cj��3		r����^`�2��Y'��t���n�̒���%=����ӻl��d�%im�m�H�\[��{	8)i0�.�nXSm���כ�]�fyC1ם������6x�ԍ�V1:�רV�r�mk��]���W7f�L#�\� K�iƭ�iq�6��\�6�o�>:>;Dl=�K��C��n�WF�;�kl�%�2��hͲv[�X�9�)6v��*�����{u�o�n=��&7��uEP�fi�%��x=��73m{�ZFo�m}���[N�鶥�q���zse/�۷{u��-rӉt��)��~J�eoLggu�;�3��e�2��q�8�1D�:p�o�n>�k��͵�ei�BȄ�v����ۉ��Γ8�L���
�M^�
l:�³����qws�mW�]����_�{;�gۛk��ӡBID"3�z׳��4P��M7M�m,�so�P��D�fH"�֍: O<^���X�ݹ�f��Qr�ީR�ZnjGNj[v��5Ƌ'ٷf촳�͵�Ӻ�˒�%H�6.I$gf�ǳ��}����Z%��� �QRSKm�}���}����ZG�ٶ���ٕ12�4��2��I�^�=K�ݸ9J����qM��؝˸���T��M�(&���smg��V{5�Z_nk���&ZqN���4�g��K��ۏ�5�}�����m�hm9�5U%S#���K��i�)(�(ԡCܧ���ZF�̝*�Щ:MK%�����>��]����Z�s$��lr�ӊT��?_�������/o�n>�k��JեM9r�uTg��-7m������/:M�
�5����ڇfC���:T�UIN)'NK\�{+�3����q��ݵ񓺄6dr6m�o��q��Z�}��^�͞B��H���f�!�n�ټ�~��36�}��_n-.����J	��~��36�}��^�!LDA�`
J�U���P�s~m���}/l��T�:T9�kͨ�ۛ�%��q�nm�_���ڪv77�\����+�(��u�z��ӚU�^�n�ܥ{́�,Ա5T��Q��ۏ�v\oۛk�3j7ٕ�S�Z'I�N[��w\n�6��Q���\��#rRc���ԑȧ��{-x�������ۺ�fmJ�L�4�ES��fN���W�$�.�0�J�*�
���t�/}�z/N��f�ُ̜DDm�B`b.C*�����^�y��fqЃ��V�$�!��l��BM��F�r�٭��؂���
:3ڄ��g'%��hR5��ܚ1v��Gek��t��k���$�/:�3���m�]��=�(�n�r��=�k�8��pݨ��u<����"��K�ѵ픮}�ᱬ��f�7&,�Ʋ�R��4��,��3����2mG;���v����ӧG��$:�Q��]޽�����w޽�cF8��Oba58`N)|QmÌ%֐���n�Ͳ���(?S����"��@G$�������ٍ̜�f��qh9tә�M�(&����mfNl��۷n��,Z�f[�)e��ٍ̜��n>�ִ=�ۣL��53I���j�TӘ��ۏ�uƯ{v�d��-�YZMԩ�)�jS��>�����=^����e��/a��Q�r&�dK[NS۞xf��^�k��N�I��y���bM�ژ6��"e��U-�m��۶�'6c}���!D/����V��J��In[l�7k3+N�W�EP�&*�^�����͵��+Xɖ�JaS-���ۏ�u��smfei�h�e9�D�M �Ӹ�w\oۛk3+H��m���sM:���Ђ�[��f����7}�q��I~\:{m8��Q'R��* ��^e���6u�s�]�L7l�������X���w8�R�e�Y��2-�f�{w\n�6֙9��M52���R�iʳv�o�P�!{��wf���͞�w�����S*S�ԧ*�ǻ��i��P����L�[nf]UL�Uk35�s��i
fZBbH�*B-��!��س���P5K�G��~Bm�a�k`�8|�����{IIl!��D��:��|4� �i��0M4TQD�ַ��rϥ%�����5MY������*����,�T��Rg�ѕ�xW��B�q933�2����0��Aӵ9�O/���қG!����6���i�F�K�5�	ɦ	��M��/��%�,Y��z"��y*q�pG��������M���JA����Yh(H%_��C��h�_��>�*��A?rDD�)�FJ��5��8#I�����Ʉ	G��۩)1:�m�nҀ�A�5���@�nk���A�voZG���Q �>�~~o�R��;�5���F��d�Z�r�أ�B���4�'~��� h�w���);�y��pK�%�<��{)U
��N���%�]nzZ�8�F�V�7g%;�x��1 ]tL�ED-Bn�R�\�¥ӛJ!.��iK�{��JF��{�{���|������q��RB���?4�G%H����|��o�{��R��~�}��S�u�s�R�������'�C�~��>�N�L�ShNf�w�!/ޟ?4>JR���\R�);��{��R"��w�-��\'#N*�K(v��C�"��{�qJR�߿{��������	!�C�'N����9�$~ �rO��7���H�_����t��uD�iʚn�D �ٝ�����8�����>�~^���hH�{5�(�/Rђ�\�t�hZ"��U��ݎs���ܖ�5.�6�y4����k�Vݚpލ�o5��);�w�)JN�>������}�8=�%)3�}���A����)�AC����6�!���}��%(rO~��8�)I��޵"��w�!�[��*��F�ʧuwJ>"D-��W���$.����)}��w�)JN�>�����
���I�9)�J�w�!.�����JR���|R������|�B�޻�A�f�(�MЪB�z޷��R��w���(�	���]���)Jw����);߾���)�C?�c�隴������o7����9���r/m���g7g]R�r�)e i��xK���0��z�;7`12�Ȼsg:F�;l���ey"t����L�l1Z`=��M�cD�{*���JN���D���IB���&d��nn�w�p�|�=*���x"��R�	Z��rY�W���:x6��mrNM�'THNv�:s�n^�ֵ;�+r���eɆ����`V�텿����~�wW���b�g�V��s�v�j�m�@�n@��ͫ��y�]W[^�x9�i�z��Tµ۶Z��ݥ)=��_��%)Os�{�)JR{߾���)|�{�)JRw�O]]3f�j���n�T|D �[����!of���������)J����>J��I�UR��s��5L��!og���)J_;�w�)JO{���%*!nk��D ����M9r�JS�4;5�����}�y�)JR{߾��)J{���┥'����%)O���ۥ-�P�j��)�q"Bջ��JR���}��)I����|��/���� �@��duW'RL��nfDM)d.��՟V��Z,��v����l��nN��}�o��葶�c���Q��!nk��D��}��JR��{�)JRw��}��JS�{���n���Z���)JRw���#��T;�9)v��5�)JO���w�����}�n)�f)J���)����@�Էj>"D#?w��JR����>JR����\R��]ݽj>!P�H����eCm�-� �o|R���{��Z%)O}�}���%)3�{���������)=��خ�%8*��۹Q��!n���)C�{��|��������)I�{��Q��!~��I�2�RS�j������{9�-�4�M�>sr�X�O�w��I}G45����m���{ݷ����?8>JR����┥'o{��W�H�[����!vn�R�-IQ)�j]���)|�{�JRz]�{��R�����)JO��;��4����m������Kn�w�!-7�sQ�)��wۊS�C��
�a�`����,�~"&b��@���k��|�"���� �@���z�����m�P麻|D �[����!owu��JR>w��R4����a�R�v�5�B[�LcML�sq"B�����	|�w�)J=�{���)��{�┥'�U;����Z֭��K�8St�����r�1l�]d�V3��+�h��f5p�w��w�Q����j��������┥'{���)J{�^�8��JR|�{��|��>w�k��ni��m*���!vo>|/�$�L��w��┥'�˿��%)�{���$������qT�TN��C�)�{�u�)JN����� �����)I߾�}��JS��w��9tک�j�N�!(A�{�G�%)|�{�)JRw��a�R����T|��ߟs�R���O��ٛ����z6a�o|%)K�{��JR���u���)J{���)JN�����)J~�A�����-�ᖳ[ݚֆ��S�zܪ<�k=���Kg�=�j���*嫸Zcn	��KN[t��!B_��?�K�R���┥'~���|��/��]� �@�W�z�������huN��
R����pĜ��������JR����|R���s���JL���gv�Ks,d��L�sq"B���Q��K��{�)O�(@d�����C䛈�!v��+�A�yd��S�c��T��o|%)K�}���)I��{�����}�mqL���;������R���L���tM: *���sz{��~JP������┥'???8>JR�����JR��:!n�~{����'�V�2��Zx�D��(�uű��ǊS���m`G��v��N�p�8L=�4^�8�^�v;5�p�k��N��Y�:����R�9�mj�N�0����@Yv�`�sG�ϟ<�2��D�ut����}Fێ݁���M#�d&��U5+�Ջ�T�԰��c�7l��M*��l�c`�k�ڵ�e��Z�V� ���������\�!��V��5Ѭ��z���td� ÖR��ѣ�D�Ղ�׭�m�zMV}�0}��?3�q>C����}��JR���|V�������R����7*�:�5�J*�\B������J_;��R������){���금J��Vup��:.��y���)|���)߾���P�=Ͼ�\R����{����ݽm�ܢduRӖ�6�!G�BD@�w�����JS��3�R��;�{��R�V���|R������kvʩ���:*��G�B�����A�|���JS�]�w�)JO~�����v��o�~g썵!�H�
-��*�+�4�;�,��:M��[S��d�Oi�}��*W��7[�nѳ,��)JR|���J�G���B�T���"�_�!.�[RLt:N\Jniڏ��J_>����~�[��S[��h�T�w��}<D ��P�R����������wۊR��{�G�IB���۩�U54�̂'{��);��w�>JR�}�}��I߾��������|R������
�(�N��ܨ��@�,�|\B���{�x>JR�Ͻ�����>����!B���nU:uJiP�R��\B%);������s ���s���[�'��;��h|��>��}��)I��﻿ut���Q�I��r!�r@��-�BӸ��v	��=�7wy����bvSRr�ڏ���1+��� �A�s��䜇%>��}��JRw߾���0����-9RK&Zr�j�D ���y���������A�{����B���i(�S0�7{�iS(��lM��]�Q��!{5�q"B�v����N/�`1lP<T@8)䦻��g)JRv������R�������Tܲ�R:sqD@B�w��|��>}�xqJR������)�(��긄!}ٴ�i���
M�7����Ͻ�)JP��ߺ�p|��>��{�)JRw�}��5K�׍�}���ω$u�)�]+��N���ZI�&�69]/`ы�8Ӎ�{����}�)�5���y����)JP�}�]�������u�)JN���x ����}�� �A�yt��4�S�,���r��JS�w��R����{��R������)JN����x>H!�rS�a�ܧ-���MU1�ˈA�nwX�)J|���┢Rw�u���)L,�|\B��Vo4�˩���mZ��J��{ÊR�����%)O����R��!�Ő�Q��3L��H��)�%_�$��<�"�[��%�˥H���&���
Rwߺ�p|��?L������)I���8>w�O��xqJR�������ڷn�����m�Cgr�.��w��nCX[�����v�����}����s&s���R�����)JN����)J|����)>Òw_u���)J{��ˢ�53-��!/woZ��J|����)JO}����JS���Ģ!-�wL�5M�j�Q4�Q�R�=�xqJR��~���R����qJR��{�x>JR��Ӧ��7�3Vk{�df���R�)I��u���䜇%=�{��)JRw߾���� ��o��+�A����~D�cMS�,���>JR�s���(� �������?8qJR����{��)�}�sk��
�*����}���׽�������s	��H��`�2B1���!��5�S��bd`�# �&�4d9��32�T�)���;��R0��� �
��O/�_0����X�U��QI2DTESL@�"�<F53�%--٬ "���Q�b|��QN�10&a�,D�|��̲2�<PѬ��>I|4��~V9I4j��<W>�����yÛ�8�V��D�(jO����*5B�Nq��d����U�ω�fd��
"Y���7�����q���$m�9U [Km�@ڂ����&�N� �պ^��H�vR�t��ÖU�y�-�w��wԯ<�f�v��:!���M�J�Es�B��R�]cs��2�m��Ҁ�Y�$��'��j@C����'y���qT�p��6�ӵ<�O ���ɺ����Ի*¹8����5���u�������4@�tcv��s���5�u��$�u=H�Z3��n��5�@�R����*�y��H
�k��i,�̝��h��Ї9omnǊ6y1WYa^��j\ݭw;L�#�F�P�1���K���k[`�x�m��2���/���Y�`g�PYJT�6�ĪS�q���2p켂tv�� 2��DE��KZ��ͳ��`um��nGUK֓�)��:A0��	�����v���A�Ѓ��)�]�Ve�H�z�q[���&+h=���i�vt�@U*�:�7cnct��#���Ʃ"s�L�e�g��Z��Q�mT�ă*��½1��*ڞY�%X�
�9�֪��&:[)	է$A��6�H ;�̯"�lu�֮��v��l
�5-E\����+����-���p�Ƀ8vQ�\(��
�qr��n|�R쵬-ب[u�%e]��5=]�s;�Nx0r��j;Tn@�ۙ��Z��m˵����x�
ڙ
�WN��&�Yͱ��v�'3�l��ϔػ5�u�t�쪫u�$˵�'sSm�
�':�t#2�LAaV����"c��{IĠ���SUT��=\e���c"�ݧ�j2�ݴ��E�l೥6�[J�IӇD�p��ʶ�R�b��鋶��\���셧�S�l�n��8˖�����m�zu��cd�������=zF�3*��-��1���s�,n����W�oI��oNs��he�b8ū:P3�� ����2m���);v`�\�SЅƨ��p"`���YgvM��cn��|���iʦڞln:��:q��m��#ZƵ}_|�\�fl���.���x(|���tD?_��}���@���E~
�����U�>��k�u���eڥ[k�9�����:��ৗ�g|g�9���m�D8���b�v�z��q�X�Oe9d�N�׋n�WMU�gr�����\�*1>*q{s�	Ƈ��T���+��W$G]�c�\"-���F�4��FV�X��!�8�8n�*�8ь'\RV�ݴ:{\�\��J��U��'X��*��i��ط)�ז�nן;���w{��q���4����.[a4�����x#��6z�㙛K��%E9�_�_�tVx]�/e���)?o������R������)JN�Q�IG�B����q"B�Y���޳0�o36YoZ��JS�{��nWt���A�+z��D ���֣�"!{��chc�A-9tU5q!);��w�>JR�3����
a���w�pf�j���Ǳ���J��wM���D/f�,����=�֬!A�ɻ\+q�ʪ�m�����}���	D(��Z�;����=��,������]s�jE�9
x:���m�z�<t�\uۀ��"����8�����S��Sr���zՁ������?��(JC�߾� �4�[�*RuR8�$V׽�w�쇂2J��R��ሧ�`EC�W˿���r�Ͽ}��ʻ��j��B���/ȕ,i�t��K����x�5�ǘG�DSw�M���͒�T��Dڦ�`���wsg8Sw�&����D@�2�j5:��#I���RNr���� I~K��pfM,g�y��Y��m��8��`�;������b4�$���X��]GZ��N������Zd�t����&��73m��L�1���}��DDt~�ŀ}����D7R�#t���ɥ��~J i��:����6�>��>���R�քTFPȠUT�����p��<?Hzt"�U��>y�|�����=�ܝ1Ą�u2S���?���JaB�����dXӿ�'6}}ORw`n�ܧ�Ԏ5EI��?eXDD}����?f��ŀ����&bw�V�b�wlmdB�n��VOg��/]v�-n�mz3vz��������g�9n�p6E���ǭ������� |�^mp�Vl���j�dM�n�ۼ�>������'8�L�����*n�Q2�R�Ss���j���M��ۯ�ۛ�| �G�k�r�6T�SN]MX~��)�k��~;�������+��6L��P4�/�?HA迀?�����s�*Ϟ����޶Z���n� ܻ���x��گ�IRIg�=}[�Łմ��NB'����I�n��M�Q3��� p����h�F�g�E�L;[Q:D/�y����ܲF�h�K}���� �N�������Χ�N=ޚ)��j��E9o���j�(H�Q!�����׋�5<�ﾀi9/�<�E:q�TS�X����;�X~K���o8}�h��j�T�TQF�A�|�8DGR�9��y�u�qc�����u�6��dUUS�M�n�ټ���"5�dX�^��J�`~�9��}�Goow]��������^EmN^�cgU��k���ٸ�8JnX�݅� ���#�A�[ɵ�u�v��Ɏ���u�s�)�vd��nn�4qB�C J�.4�UwC�(t�϶�Eys���j�.۷h8�K���0=���L]]:�l�,����mh�P����r�-�K�/����4����W����m�e� �rSŝ'�n�Afl�Ʈ���!BV�%Y#V7TJ�*[M��R�����0=d^f۸�c�u3��8%�������}m7%���G%��Z�7����;�4��}��pǻ%H86���r��}ئ�?�L��x�<��`Iڿߗ�3�Ǳ�O�r��u�;�L�:���">��,��� R�%�R�Z
h�Ke�D${s����Z�Ks+�~BKۯ��3x�)�N�9Rs�w3mX/ߕ$�[�����gŁ���8/b�LNF�~r�T�\�%��nv"�[��:u���y�U[�/NyU;e�$�9����%�:r��ڰ71�N�T��[Ͼ��0Ƨq}���rƩ�iM1�����{5�/��B�Q�!'�V�����j��c�J&J��k~�F�MUO�I�����ٽj�(F�t��_Dp����F5HjDT�'9�B_��nՁ��ݮ��ńD�����}��aL�Lr�n����_�_ �d����w���j������~���%!���®��c�-��%��:'mv1
��eu^���������XܻU���ɥ����8s6�����ξ>g����A����D�Xz�a��@u'qb���l�:�2����s=��H�p��ʓ���j�Ͽ{��_�ҫ��+��>^��,{>�ps5GQ�䢪����"����������^��G��N������jIR��F�g �i`Du�;�;��Xu�0�C�}D���[�:JcC��'[�a�O+�j][Ƽ�.��L]=m=��/+o���{ـwS���}�u*e��6�ƩDQ����W�o��L�W�Zy����MN�U�����f*���*,5��u*e�Zy�w3mX�͑�%SuU˅�1����*e����Rw�~�g�G�}
>���I���_|��ꠈ(QDQR:�3ۯ0&wSȰNـu*e��#���y�,�vm&mw&t��'cK��#9zqkN����]t/6�u�������!���:j�������[w���}�t�y{٘��'.+�TI'**bI���Nل}@u*e�K��p��/�}�DE���ɸ5�ڥ"�o�pnϋ���G�}ԝŀ��f����uQNh��&�7ߑ���p�m����8s&��[��'M�ȝ9UU�RwE�|�����2�ש��B��P�B2"�q�UML�eL�i��l�mն��:�yk;  ��[u��3���u�t�m�4V��ASێX�;u�eq�m,��M�e�!��`9�Z��DbW��6�(f֮�c\Jk(<t�#�%�����)���^�rv�n���Ϟ��&�Y);����6�`n�iV����Ѵ��ënصvĤ�ܲLI':����:A �ˉp�9Ӷ'������{�������ChW1�v��7�mcq�-`��8+�����R�^��g��}��J)UUR��n2���}\�ɥ��ݬ�Ap�m�37dqH:m�\.眻���S/�1�� �N��]Jـ)k����T�@I5E��'����X|.�l�:�2���UrfbI����*�� ��N������S,?�/��w�߹��}��N�r�N��
AR�,>Z����>����Ł�oـw3mX_��#iboX�*�IڥT�姮K���	[��8u��WF���=��v����"�*�w\�ɥ����p���� w��O�t��6�&�"\5T�Z��f]�����4��+) ��cX����bLc(Ĝ�\X��2�1T����$2���D�"��==���녁�ܙ�\��KI~_�uf�M��U6�h�O���Z�;�����QQ
�G�gŁ������`�O§JF眨��l�:�2�m'��}}KmX��dq�*��K��t���;�4���!���I�X)s�ـv�χ��t��%��a���ݮ�.�n.��7]L��Gf�B�Mp�;��H��p\gT�TX�~��;�^��`Y4�3�׭!�"�B�Np��=o# ԩ�i<����D�'���䌁*�J)9��g�qpfM,�v��q�m�m�n��~]���RC��'��|�R\=9�Y��O 
HdvȺpڱRl���/��C��	������hvů�$�7�kf��)[I��ڞ���G��
��M1> /���>�uwϪH�P�~x � GK!���4��Ax���~y�w���|̾�����T�G�T��Y�=�X����nڰu���۱��I#*DT�i�w3y�?wٶ�����35�՘�E(JdQҧTJT����6 �V��I��î݆�3�r���h��r�1�nD�9��fڰ7��� �{5���ۻ�8�}>�0��NB���qX��0�O���`I�\�Ӧ�5*g���\�Cnݟ���3�{0�L�~����� R�'��
�3<*���W, I�Y�u'q`.�l���?�&^P
'���X�����@Rn�
�V`I�X	�`��,�����_�~�b>_S�EJ�p�����R3˶����ϵ�k%׵hɰ�ݎ ���{g�ܒ͹URQH*H�~ϯ�v�5�������W*�fn�jE �NE�,�:�,�y�d����O]� z��a)ț��D����nn��{ٶ���Ӏv�5��ٱ7M�u"t�\��G�DLk~Ȱ����I��[����6U:%&�%D���`{sm���>�5���{���;����}�0����ӵY#��j���cHt���awYP�9��=[	���oa���=����p�9����k��X%��������Mt��+pq�2YJGm�\���u�ZS��-�m�b��76�0Ѷ�����*/<w[��=G}u�q\���Z�N�E�B�Uѭ�O2��/^y�bS��:8�k�E��3�.yU�����LR���ֶu�~�����w��wW�V�:�b��m�Jf]�u�a�������vq����6���;]�3������b�|.��ʻ�_��Z���;V��zp��OJDMR��BuR�X[y�@u'q`kNـuq9��>��h����������j���m�����5��`k��`cpr�L�T��UQ`j�l�:�2�Z���(�=��X�ܨ�-��Lu̳ �T� ����xRwn{f� �k�Jl*���6�STFvmFl����ۓ����莉��#i#�,�tk�.)N47�&�7=�����V�ۿDDB���k���Y��SN����SU;����������� �%�s�������}!��~�2�OӾ�,i<�7vl�(��$�Dq�qX��zpΧ<��>�M'��5'q`$���"���.�IN��8��K�6�����dP�ygr����Mj��'"��倚O0�:�=�l�;)>X׻��~�~�e��`�n�9�y�ssq��n�q]���{sہr`�m�=m�����w֨�5 �Rq����V�6����w����p�몴葍�T#���;f������'L������E*ID��[��n�������؇��~��<����.U��?=��������5�S�mG`wsw�ک��"�O+ �!N����뜮E}Tک�-��;_���;�^������f��8 ���)J9T%NE?`�X&:�lq�^�jvb���l��Ԉ���H9"���7�7_ ��k�7y�">>�:�׋$�U�e�r�g&�y˫�`
u>_���4����l����n����:c��aL�
�!`nf<�:�2�舀���9�T�Gv4{	G�2S�D$���K��Gt��{�*��������) �%7�K�������:��U#t��#�����`�J�`6����,�N`�p
7.�-p=�IaQ�xͷ����(p�\�f�5�������|.����Xr=��� IS"�m��[�~�{����l�~�GTԎ�o�M�����*�G��|_&O{����-TŞ�����ݩ�EW&~�D�9�ﾟ����33mX����ٱ�C�*�*�o]78I�XSy��~�z�X[�TMT�Էr�dn����j��%߷�w�o�^,�m� ��V�=�}���ղ	1� �s��JX�> hݎ�l�L�фH��X��F.�r����V�/M���dй�8�ݦ�rµ�ٰ� Y{O%�2���WWuT�:<ݗm�v�U�X�a-��0\�Vx�;�Y7]v�W�"��2b��N����Q��V���52��h�S�Y�(-�D!{Vv&�XW�]�5��[�qi0%'(�.#�Su��{�}���=�{����ߏ���Cjx'�"62�t	��Z��[=��4�b�n���c��7�4�[��S��U7��ٟs�wvi`o����j��|�{$E �T#��u�e����`	'q`kM�-Qp��%�#���{��{6Ձ����ܚX��	
qTr*$P����"!jwm��;��a�">�Eo�>����ߤR�(��RH�i<�7]2�Oi���5��~�zx@��a��n�Gd��l�ڸ����[����u��5Ɖ��h��Sr)5��XО��7[�=�D����� ��8����"*B�޿k�������������Ł���`��`{��$Mr[#���*]� ��mX	���DD}3������x�\�9ӤS� )��������,7;��3w�X��.��*d���-t� M7x��,�y�n��Դ�v�\���1vtr�W�A�d�6�fZ�ۗ�R���������pw�ԉ9�3o��vd��wi<�;��`jM��7*S�H�*��z�fڰ3s7���K ������Ԏ���&ԕP�A�n� �tɹ�����?DH�_���W������7��`n�,�I�EH�q���{d�X����3۶�{sy�72'�$�!�Q�EU!`���[��m��S,�OP����إ����\k��i��dc$��mq�v�ʽ��Gn�mpv�y���B��wx��,�y�n�e�jm���uN����(��`{7us{A��������E����):JZ�S!*� I�,��xz#�D��M���}��{��hr7D� nHX�6� �M��Ԝ<����7��"?z#뤗���X}���:��S�H�*�����,Bk��@o���19u`n�;�߭N@�<��I0� ��t�ۃ�e��𾫃F5�(!��6Fz��z�{-�z�� �闓!����������H�q�����K@��`v�1����>K�>ߣ�$�	��W ���,�:�;+W,>5o�`N��=�ݒ*pG$�[�V۹�=Y���<��Z�MՀ����&aI�q@��v{7y�3�4���`v���$���`�`�`����߿����Y��Qf��<Y���dв y
�� wh�I��&(����:���o��f�ߓ�d���aRf�H%O�Ҹ@a��SM1�83ۇ�L��B@ƃ^�:pN-"I��aϰ�	��`�4)G|��*�0��s02�FE��X��o�'��}�I#�-�z�lܭUUT��� ��Tm�H5Ӛiki6�D�YVѻH;V�@[Fζs&��(��n�f��S�]n����>"M����uPY�L MU!J��QV۬�uJ��YP ێn�qm���h�Sƙ�ε'j���Hs�Nwj$W��G�gtu1�lc���0�f|�Y��vq��	��a���N�W$�㛜�tRH���jۭ�g�@Y�Wm����*e.ѡ͛;��Ztݲms���#f���=�#�Jv)���us��)Tkd��H9��*��8:���PʲTR��NC��6峈C�ְ�	R�����Z3�T����Gۮ���<�xM���+R�p��$b�lKQ��gu�n�ՋD�P�MR�u��k4� (��l��6x,��.�ۙ�]���d0��vƣjŶgU�-�9ê['W�]r�*��@��ɱ��kp�컰UN�@�\e��<�1p��˵R�L5U���h� ��UT�i�	{AZ��3D*I���ݛ^����l�\�%�2(���^ݸeVTI�Vڥ��t+p[fj�QĠ<v5����x�e�s���{Z�-,���88��QB����E�a�Q�/7�bMG�Qu��^���ք��]�n�ݺ����e���әd�4� h��hzp)�C��9�/@��6�ې�u���c	��9��u.+�b&.u�J�bH��@dv����E�I�C.�6���@f�����B�5]V�V6Ӱ� �E�킘(����v5 �����-��+�U�VU�p�nND�s�!�/�0�l��5�x��d�a)t;�Z��^�s��]�@k�4�n���-Ѻ�5oi8�C���q����۶^G `�3(6�.79�$�;ar&؉ثnӠ�
mB��Cy5�ʕ��Z�6}���V�n'<��`ͮ'��q� on�k��3�T����{���I$���Qj�5�4�<��1�(H���� ��A���l��!E?eOޠ@;D�'�QM��`���(ԑ� \R�ҟE�U�
��>���/���f�֌�曎8جv1�Y[�+u���l��\ɛ�qu���3ٝ�ir�o="FW�����d2mi�eڪ^p'0^�)W��	���S�c�1� e��dWk�`�L��p���9s�)�s��;&o/g�t#�m
����n����P<=���5��:'M��1��Ӕ���֮+#�c�{m�� C�/�wow}��S\neل|����\�;)��u��k�ӥkA��d��Q��p�}��A�Rv����������������O�#��A�{ـ{~���F5(��q��;��;��V\���`*e�����ɮTO+�G2���W�u��N�`o%��:�4�H!�MD�m�����5���,SU`}G��%6P�:��ER(�Ch�s�fl��=��,��U��{7� Z���*�D��<7M�]��Ǭ�YX)&����$�.�s�,Б�����Kv�R)�q�"HXsvX��M��5<���}�Gd7ޯBp�����-�Թ����[�����I�Pz��L|˻���<�����+ �n��_��Te{]0f���
$�`kOـu�e��}[�w�W.f�{ص�G��:�aT�� �l��3۲���eX%�#���p�V�m�:r�D�L�s;���J#�׵6�7����,.�Vlm��r�E?ԣR9�-V�U�-��XJ��y�N���s�/K�n�l��&����wuX�L�:�<�5:g�~Iq~_�Ͼ�kk���Q6Ԏr'�������5:e�-n��_��Z�6F�(�E�ӢI��٥�vw;?��<��/)S|���;,�>�s�o���N���q�B�,?/����;ݚE����R�XZ�T��u˷.T�m��ǻJ����;�٥�ow%�s�9H�`��9��m�����������|�O=n{-�YmN��
Es&�ͷM�t�8�UT� ��~� �l��;ݭDX�zX�����D���+0N����@��S�X}��|�����Q5)�R�r8X���R�X}G"V���]2�ޤÅMG**j���]�V���^��������z�r�cGO~�?�tA_Q)U9�,Wk�#u*ImF6�`g��`	�|� �j�J�`w��\.�(�88���;9ʱ�aۈ:��-��[�v�k�s��q���������rW+�E9|3f��ܖs&��{ۻ� ~_�{q슛 ��UJ� �j����:�"��M�JN�`u<�U"��T���pn�,{7y�	(������`d�eM �����fj�u7��L�mU��Gп.�&{ڵ�p���#ET��S�Xz���ΪE����~��ȏ�^���w��
Z�,M��O ��K�b���HZ^n݇l�3�:1��q���w*<.�C�pI���s�j֎�'cN���"�nG`N����X�u��m9�5��e��u^.���D\x�N�r��;N�{Z6���M�n�pn�8��k�5-�*�e�*��E��;����em���H\�̲��Rr��nf��KuǮ^�@�Yݝ����{����w�����w��b��[S\l2a��D�����ƍ�-��4b�	�v��iN��5$U�,�άH�{$v���(DDD%{��X�߂S����cYʫ�S�X���5�e�kj�����YG+�쑺�܈mD�m�����`�q͙��&��%H�Ʈs�����U5%U�
����=����ץ�ߕfo�w�}��詧)�lU"�B�5�V}F�X�����,��'~���ӹGCո��u��<F4��mص.��#��Ń�ps7U778ߏ��Hyu�$��o0N���#�}�Vױ��2��5EHX�}����=F!%S`����"�!Dx9�xX������������ϴ��nT2~mUT���O��[U`f�E����6e�Qjjby$�MI�E��"���������� �l���{�)P"rD�����5:e�}�n�� ���������Z`�cH�<b{]���˝���s�n�v�GK��R�>o!JB�e뗕���i���,�[�����T����/n�C�'N'N���3f��Q&����[�X���D��I�sި��ƪ�ԩU!`��K;UX�*���V<iI�T�Y��+�̲"�&u����A~c��Ϲ˪;�O�����*�n�ԫ�]V�)m��޴� M�,?L���`z���-����Q���~�� �>i�,���\����BI�)ؖN���uܮ�ɤ�[�\j�2��el�Pc�Q��#u*(���U$� ��[V�]X�)���7�<��"_
��)J�"�p�o�Y�U�yu`{�����KI��Z�@��U˫�����i� ��Xu��2{:�T�)Ɗ�&��v�#���pn�,��~�|����R�A`���TD)J�P��z�ػ7H�r4���I��'L�?}LDw}��5�;߳y����IJ0��R�$��n�&�>۫v��n:6�n��6�N휁�:��-r�6��F�J� �we��y�`w��ėUc٥�՛�#Q9ʶ�����8�76�O0N�jdWWﾈ��M�c�)�	$j"�9V��� ������g;�ٰ<��u��M9ș���>�� �][�t�}���W���_���RJr�D�L��u`z#�ݳ {�{0*Sv��v>���ݏ{�wq�ǽ��y�o�^�YN��G-�-�wHrg4�]+`ڂ�����c��@.u����u��Rյ��{�=�y/f�c���]��Ҭ�:Q�Kg9�tcpɷ!J5A�cv�Y�z���T����
-����,�%�w=8�1��9���BR9'���;Bd'˷\�+TY(���7b��c���u��A�zE����6����Q�^:�����s\�xZ�o[#N�i��kr�M[v�ZumC�㴜��W/a��m��Kb呉�P$Q��MVJ����Ł���pݚZ �{e���J��7J7T���"y�,��g���G�W� ��U��Ʌ���f��ܢ)R'N���7L�֪�ԩ֞`:�*�INjfGI���d;�`{u�`nno8�٥������ʷn�*U��n�`-i� ��9�֪�Z���q�!���M�L���Ҳ��GeJ۴lv{��,���Uj-�p�#�I�\���TXZy�$� ���!�ݲ���~n��l���RNp͚]��� �AP�O��DG~�/�ʳ�2��XZy��>����K�#E)R��%J�����<�}�?#rf�fl�«��Z�"8�:�8���V��,�O0N�a菏�M��.U���U(n1�i�3���#�O�� <����E��߯����2g���&��P\p:����*N�6�x.���ŷ\�/h��C��r}����E#������������;�|��$�����犪�b�9s꒦���U��C$��Z�`�2���dj0��ܸBU��pcݫ=�����C�o���y]�kU�����s��9�@R� ��P�LĨ� � Ԃ�ԉ	�P(�$��!�y��|���k.N	0L&$gɁM��c� �#?`�|�k8�����{ڂx
���@��w*���Np˞o4��s9�0�)K���CpSUE-p#$#W��]h��ј>)�Q�"�!���H�
!V��|�Q(�G����$�?���,���ެ33O��c��~�u�o����9��h6hѣF���P��~���U\v�����B�i�����=>�)���[Q$~�?��:X>ϥ���:y���$ɪ,?��{م����X�UX�0�=�i���5M��QQÜsf��ͥV�X	4� �rj����Ֆ8�3hs��#m�͗�ʸ���G,sL۵��z�Z�:.;[�����i�,�y� ӦX�0���H��H�p͚_ߗ䪍߷�p}���`����9]�<����8�9��M<�t� m*��E���6T*8�)T��8��,{��2����r�G��X�d���`H��8�.��|��~�s_���"��
	!`���UcɅ�����L�?}���9犘��&������y��H�d��M�<{q��K���]�]`8�(�(]˗R�:w:�}>,��9�76iaU[��`sy��S�n@"f��m�֝ŀ6�Xݤ_��}��RHRE2P���{��Հkm� �S,�y��Z��ɪ��̕5O*���}>�u`-T�/7�_��o�Vsu|q�*IO�\�5;�M��:Ӹ�ҫ�~�ߢ>��$I�@�UQM%E@��1�B1��w~O{��]��8�����j걃���Ju���u�vn�pl�ɨ�Z6�d#�]e7i��V��[uφ�l��a�5Ֆ�6D�sk���o]O%8L��Vcbg����9��
2;<G �ˍtA&��H�Έ�u�K`M:T��.�v�8�1��qū*v-M�mΎ
)X�fW5،F��v;Em��'�s3��<�˜&d��|)k���s<�p�4������������e�y�	l�)q�� H��x�9\������R�"Q98�Q��h]s�����fڰ����{&��/��H�����M�P�0��,�����!�t�`	7\4�4
j%��e�Vݺ��=,�}2��{0��Ł�'UȮAQ�7v�uV۹�Tg�h�n��wsm��̖+<��S�r ��,{wf`i�XLδ����"�e}��<%��\fywY�wN�Z^�	����N����^E��;����v�[n�:�[���;� �%V�i��~���^���q9UC��
���=��˫��#��)څ$(؄�����?n~�ۛj��n�r�$nErGs�g�i`ki�֝ŀF���[��U5��Ƣ$cp����$�>���=��j�3�]��ǥ�ܻy��6ښ�MV`i�X�>�%y:��e��i� ,ͤ���Q�RGJE��lv91u��k�ͣ`{xZd{=x�;�F��k�n�y�ԕʋ ת���,m<�:Ӹ�9��#Q�~����%�rp�M,�Un��wsm\�w�,Vy�Y����L�6�`i�Y���}�p�^�3�K���o���2T�U��i�X7�\������p�1O�9N��QR9�{��`|��zp��{0�Ł��q)�d"f��PK����ɧ��+����evwft�����k�H���G�Ȣ�Kw8{&�7wy�;���\�33�`o�6�R8:p��
�r�<���;� ��_Xݬ/���Q��5�T�#�H��T�8��\X�u`ov�`bm� ��2������#D�8�U{�,A��L,f��W��US�0J� %�@rBL1TJc#��pL��1h(� D�jDPҩ`�
�3��ֹ�r�>}�#�Q����(�����V3wy��w5`���I?�!(K���ખ�r�ݝ���S�6��v�βZ��n{-�6���;<(��dӝ�٭����������{��X{9���U`{ش+���b���pnm���}���y�`sw7����F-4��N��Bjwά�i@[Z� m��=R0���mJq5\�w8cͫ������V��b�3���F�J���m��X֞`m�\ %�� ��/��>>� IaN����k]ֳ{��ֵ�<�.�N��v�Z��J��=��q268��tg��L8۪�S�!���۸�;�G�h�M��mGce�tɇPU,��У���0rv���u���s!�ɓ�-s6e#��^����lv쯷��:7h��m�$'Un�A�NP��{����bٴ�,g))s3�;��j�Җ�AԊ9u�8'Y�ɞ޻P�{��mMr�ۡnPɂ�y۷m�Í�8�F����nJ�3���q�n:qJ'���E9ށ�nڰ/k�w������u��"j�	�A\������u`n�T��y�vZmX�샌�ww#q��I8{&�6�a֝�r6V�x����8Tl�t�`sww���j�=�l�Rg��`|��:���lS.����ݮ��7uՁ�橰1�� �I
F�BG�2���T< ��������;��V�m����c].��V.r��@�n��w�-�s`bm�֝Ł���)���"k���9Tg�mZ��hKW��>�-c��N��7uՀ�gUTW������r�n��.�m�?�_����X�Vڳ��d�"�Sh�Y�u�q`�u`oy�lm<���U:"CiƉDqX�� �_��m<�:Ӹ�=���#އɃ�	�^��S۲n��F�T��]�67�S8��fw<����ʳ%��7�1o���v����y�u�q`֪��[��%�R��Q��Gwsy�;�6ՁU��N�eX�� �B�����޵`��}+TW���R�UDW�W�B�����|�M���`\L�)s2T�M6��	DL�o�`v����nox��j���AI��q5�QwX�L�1�� �N��7�U�_���FKcu'R"�[��%�R�h�x��i���v�g�ݵ��r�bFb$�����-�74� ��ڰ��=�L,պ���T��"UNs�wsm_��""f�XU2,�'���&N�߿53J\QT��95`����zXϳx�}�j��yc�\��J\��4\�UF���u9y�w[��>�[(!�P�S��� = t%[~�`uVc��Sd����X�O0�wE�.�w�M�ޏ�||����-�ݍ�.Neܶz9۰�;b����m��.x��v.qV�Wm��cM��n�u�� ]�VzsT��y�=`K��R�N��7"��X�~ʰ9����fګ���r��q5�.�gv��O0����w)�����r�������)ʰ��������Հg}��\��U���6:u)9!ڪs��͵`�lVeW|��������}��H=�FA~��!3!<�����"��P��Q&�!$4CT-f�U���'�<}��줱r�ް��}�
~A����`�j~H�� h���8N}"b�h6T'Հ�ϓͨ�Q���_< �"$���a�JR�r	@9-	!�Q� N�Gߎ�5�!D�������-FIZp�ƽ�Z��
�#Fڱ0ľ����a׸�����S�1��<�V��'2'�h�iʽ�����7n�������m:N��U�f� �P�J��%�P &k�6ԨU�B� �Π%0[s*�,u�ZEl䴬���N��]����|q�*���iU�;póJ�6M�$�
�$�Y�� Ъ��7sb�b�X΂z�f������uZu2ܫ�c���[Y��l�����n��i$3^\ݰ�r�v��(�>ƲR��.#�ĂOrV�Ärc�$q̑>P���7 ��6�]w�V����Й�D��T�e˹B��7K�㉓���p�<w;� 6ۅ�]n�lF,mˏu�G��5{����s�c�l�=��rD����El�m��9fBs�j6�S@�H�07eR�TV�^�*�@�ۑ�UTl9[<�x�!1�vN]$����F�B�iV�;
�uYI='җ������x�![6�,[�Th)
*���:m!���,,N!���׆��������2�ְ]2�i]�U�}���cLFyWeڪ�N�7f��5�{��g<Ц�jƀH��ĉ�YH�Ӌ3����R���M�:�9c#H�t���u8eU%ѪU������[�g���dD�;����=wVcq�u��͎�f�g�jl�!��2��I�.��s�{t���pƵ�uQ=����s]�{f�����-ձUq����=� �J7&��۝�:,�ڐ��e�nr�P��
�A��6�nyٹL�bc[MAI�a#;����Ui$n�[Hl8±��\�$�8�i[mƊ�P�����$���;k)Z�`�`ݗ�z�15�:h�\�X�"�!vŦ��ˍ�h-��E����X^��B�:3�A��0�ů [l��ung՗�:�����@�����tX8\�d�SN��[bB�+nB�.��'',��x�15.�vl�s�`�FLl!f6��J�a����g�`����������m�Aӈp�N"�H�:�cĜS�D
3�3������m����R�	T(P�B�J��UW��+�:�Q/�M���`�~���"��J%
-V|m۪�1˦T��lM�/-ۣ1<=;����Jvc���v%�OGul�¼�����v�4v�xՍ$��f1�]�%*��P]F9,/`� OnڵE���ӡO=pl�^�x-)��s��y�LD�r�9��v��|�uC��Ms���拲��7�5ӕ�C��h��7=��Vg<l���l� �Ō�Y�g�<�ӪT5掖�\.�P4�Oǻ����{�mu�!���^[��sv�oW��sɷS��[W6	ݳ�ٖ�Ɇ�.M��D��_�@��`s��V7sy�?�֨͟Z�;��|���#��u$� ;�NlM<�;��YّlS���ȧ��)��ڈ��X#�����n�g�b"d����̭�=��_� �t���8}�j�3��b*��=�`s77�6�rV�5R�N��7"��X��"7i9�:���u�����}���?�fn���:[�\qm�e��Zڑ��/7W�lBtx�!�e]+�vɪF�G#�Wu�5q�l �����ǲ@k>��ǮR$�9Q�NU���w�tBN!/�!*I�o�Z�9O�kv ���V��ݑ����6��� ��X�u`w��66�`
Su�P1����8����Wi�*�����9Tw۶�~�����wI�ʎJR�UX����w����5{�3�.�xj�x��Q��TM����M�sa�;g�]w-t����k�XA�og5&�2,m�j����k�7 bi��n��u׾�2C�y�`{ګ~D*��H�Q�pA�7q`����y��a&�`(%�r����V�3��`.��*�J}��%���w����V�ڸ(F�6�k�]���J�&�^�����nڰ�*���X��JQuM��ʛ����ŀ.��橰:������@�P��R'�%H�����1�Yq>��zvP뭴������4��ƺ��UNs�w۶����`uW�����p�n�#��i�R"T��3��~���d�������`����5)ų�ں��,�N=�v�����p���߾�`��+��Κ�(`�q���6��{��޵h}��!D$Ҍ���BO��́���Kt9ʧS(��V`����un&N�76^��m�~�_���ֺ�{6FN3u�*y�����f-Ǟ��n�hv[�t&��=�\`�D	��g}�X�̫�����ٻj���"J�:n(�%����v&�`��� ��u~���F����5D����Q�9�w~߯�{7m@g}���{1����$h�ȜTڪs�@jn��uՁ�Թa���� ��a߿4��̈M�2ꚰ�s�=8�,M<�57q`'�(njf��5"��y`.�h��
�$A���.�j�,Jp�������pkT���������td��v�e��걛T��xl��%���M��96�k�nPb��s�7e����OZ�]n�۹�Y��5��ڷd3÷m�Lf��4
�j����� fy@:�y*WnvR2�s�-�+���v���V�6^��R7g:����{�������w��4c�D�9u������q�ĩs�θ��pUҎ�\kɺ1̔�[}�����]���������������V�����t�Tn��j"TQ������V�������G���(ʥT���I� �~�ŀ-�VgR��y�w\ԏ�1P)J�nE`�l�;������������(��⋒]��q9�16� �q`�]_&ODG�8n�q�,��\�"�5���R��E����F�<Eb�n4i ���'�8�{ـw[����,�����j̓��U���ns�w۶�AD!T(A�����\癗yجu�*���� �{�:h#G�H�Tn+@�l�z��g�]߷�pg�+V��{�9j��n�)d�p{�́���u�� [����J����q���U����p�vՀg����_�������TQ�D
uIÐ鎜�
��9��Gc%�q6v蓉4��dT�McD�U'AU$� �n�X�z�X��U����p��Ul4R�P	�,n��;�j�16� �kw$<��(���MrK��=�V3w�ya�����P�@�\����
�fd�3{S�$�QGE9V�����n��2uՁ�橸C!�\�*(�D�6���v�ٷj�3��`w��V3sy�����UTl��#t6��9�݋M������u:v�
ڲ=��n�mZ8jDۍ���H�Tn+ ��e�޿e]U#��7��ݵ`s�Ǯ8�.H;���{��W�Twwn��l,�� �{���?ƪ5Qʰ9����wZ�A��v�Y�`{��ɡ��2�TL����{;�w���`{՛6��$���d�� �l[�F�Q�7"� ޵V{�S`u�� �q`8���߼=���i�.�1pi��8�v.9:�S�Yɳ�g�̆x.�qU�uu��͕n�ʪ��7x��nS���Ǿ�>�$��ڬ�)�u�&�*��ۏ0�w�ufL���6pӮ}5T㪉�M��� �斬���r���c�7sy�36`�M��UTqXzej�Xx����`i�\����ۜ�K���I�3�6�n��w۶�����.������q��6Q2;V���s������2�ʋ6.d-�Mx�Cy�rV����u�M�{E"[�N]�����b�3�82Z��C�Q�ª��ʥINz4Y��m�gs�����um��!oL�̽���lE*�v^W<a뤬��9�e�l��s7M���J�<����#���BI`·���j鳵b���\�2�jn�϶� lh�4{�����n���/��;vI���K�S�`�0I��]nv[�[&�����Мn�q�)Tj"���3�?��g��E�n���Hn�9�7���s��R������ ^��X��U����s�*�s�UJJ� rH������T��'9�{ޮ�	��X��ʨ�)r�\��.�<ڰ9���r��nڰ�d�9�c�̊6�qB8��nU����p���`�l�=��t���*�J��UT:*�؝�a6�s����ٺMӵ۷G3k��^��J^q���M��9�;��V�3��`w��J��no8c݉�r���#D��V7���I(��j}�̧�`g�����ڿ�%�U���2�N\��%�I������� �q`�U��[�D���"��AR�X}^߷��g�Z���;���쭔Ӊ��0#��u�q`�U��橰�������������8�5�ٹ�X�6�Pp��έk1�..-�]];&�m]nt���q&��j�0:�����j���� �n��塮��)S�D��8��j�����ŀwuՀ�N������ITʰ9�����W�mYK����vC`6�����v���v�v�JY��#��d���8��&�f��1���蹲+5(豃ZQ��
�0��L�L�&M��`36Mf��J�E�9�0ѧ�>zX���K��d�"�0�p��K$�� ��Le�f�!20�K�Sv�#H،���0�^8n?<Sݴ+�d9�`a���V/��q����@�_��W�TT�B|O�:C�9�4&��/����>��� �^[OSr�TN*m'8}�j�;�l�9��@ssw�1��
H!�����,u�*����8w:Ղ;�Z���K���nGi�[<.�u�J��g���N�h���s��&�U��_����*��9U�-�sas�7�u;�9Tw�e���8�Q�Sj"��`q��=2o��,R�X�j�L���Sn*C��&�I��� ]��X��U��n�8{uZ�r�5*P
���=����VlۙFx��P�Q�(�J�A�!�Q�����=\��R�T�\��p�͎���_��o����� �{e���0q��!U���7MH4����g�u��؀�#<suۢ��v׮gl��Ȟsp��H��nU��no8 �mX3�,��*��ܭ���j�qSj�u�Zwﾈ��z��Nl�'��u��T���F�R�V�ϥ���j�G�L�y�0^�Ł�W"�$e�ubnܶ�3zՁ���{;�X\�l���yQUT���*�V=��|��Հ}�����fՀ�C!%�%PDFD��7�x.j�nJ�.��䍺�,TU�ҵ�q�V��A{f��գ��vj	��e��â9�n��w8��۱ʝ�?�.�'?��M6&�pRжO1\�G�	���WllO���'6Î�����dZ��i�Ä)zd��g�Q�[ō!K�y��I�/6EIYyqS����3h��.�t����@u�1���3L<���z�Y�4m��{ߟ�����`�ի�탶C�0.��cp�9v6�:M�ʽd�v.���s��Tn*D����9�ٿZ�g�X�fڰ>����7;���u!)ˉCm� ��Vn��5��Rw3&=�ڕU!*D���w3mX���w3mX3ڥ��2:��dR�RE�E�ﾉ��p~�ńn��;��,Ÿ�*���ASh��p�� Ů����qp4�`�ʎ9�
��%��Un���ɶ�d:ݘ�]�<��RiVwj}x-;h��Hn����m���]Xo=��}�}���Ł���N��}v�X��4��{;�^(ȅDG>�}�G���5'q`�u~��M|\{9Iڊ��F���\ٛj�=����7mX��'2�ۙR�T�f�""S~ȸ ԽVjWy=� ��W
� 5*~�7"��rX�\Xi��Rwzl�0r��P<ܺ6��.�wU;<�[d���"��\�;9^�z��nvd��DJ@�	N&���;��Zo0I�Xu��5���'��IT�8��f�/�R�7~�`����v��DL��~�_�L%�mMR'��o���Y�� �>����J�<���g~��;�y��5%6:R!�n-�/����}ϥ���֬�fo8�vՁ�{64�U\��݊K�$�n�����[sq`�Ձ����\o�������܅�#�gs<�ʺ��v�\]���G��#�kn�-�ƫ8.�Nr�{!����2.7q`Q���J���g)9�Єۙ�T�|wu���&C�ת�L	��7��{��d�~�tGC���+@��K�̵`s�f�{wmX���T�*IQ���uЈ�}>��E�^�� ��Ń�7��t�P������_=���c��TR���G��n�8�uZ��s�37mX��=4�4�(�u*[u�zg'm����Ѷ�9�}��8=s��6����nJ����M�U' �nڰw=��sٖ�{wy�7rlQ7S�T�D��TXuk���Ł���Sw w=����Wpn���rpf����}��L��\X�ά���TMQ\��qECqX�ۼ���V�ܜ�/ʽ��+@w����� A�T�RNpM�X����ܬ�7��o���@'������@F44wv���v�tlw��0�*��@[l����!�ʻ;EJ�!�>;l\�:��q�n��*�)78(�)��s;�*�)�Q�>���7fjC�5�zÎ�6�ej��Z��C�\�*�^�X2-VG�\3��+/f]����U[9���q���1e�z�M�t$�$+a�l�#T:r�z���\�7bR�ٺul�ۍ/N���ж,���k�1lt�������s'�q���f�`ۉвe�d��dw�$1��Ü�p݋�V�*B8��uH$�x���K{ٖ�����~�莾I>~��7�<z����W9Q��r�����/�}�DL�{��S��\ ��K�:u����*c����m� �w��XԮ,�ےH�"�Sj�Npfm� ��K�̵`{ۻ�7�6&��S�T���+�mU���Ł���I�X���������я��,�p�Hi�2��y�t&��8.ݦ���gJmӎ����9��n�%�����V���w�ٛj�;����g����#��qECqX�����L&�K�
�Ϸ�X �f��nڿ���T���|��8�9'8f�j�:��:�ń��`)qtW*$��MUE�wSw�n�q`u&��/ʳ�\V��G��6⋎B� I��c[y�d\n��;���}���~}���?����k$�{-Uh�]��utb�փ�4���5煁\ѹظ]t�庢xr����f��� �J�2CuE
��-ݒ)�E"��T���Q@Kj,�]Ł�ۜ��Ϧnj&9J�1���MXws�37mY�!BZ��*� DD�"`�����Q�fڰ:�ٱ�4>T���)q�9UGu��u���w������C俘��"BS)��3ٛ������߸�U߾�`s���g���#eQ#`[(�'��W��Z�wK]':XKƆ��;Y;���ڊTP�RG9�=��V�1�Vu"���i� �K��5%G$��`�yU��cj��W�O0�fڿ�*��b�(���M8��r� ��\X��u;� ��X�Q-��i��LrE`{ۛ��nڰwk���_"���3�Ձ����6�5S�UNs�{wmX7rX�e��G������4r����'�Ӑ5[���Sێ5�Φ��vr-�M��1�kWf�T�"�UV�܊���Vu��������q`w�����a5W55Su�U`	7q`֝�۸�MU�����Q�ڨ�L���no8����!5VjW4�UIU3�MH�V`۸�MU���r���o8�Vӷ
��GJ�"�X3rX:�,�O0������7��?>r��Y�Y��{��W�]��R�F�2��e�7�H<�h�Y�� 0MX���C�C�N�I�+�eI�R"㘘��lGq�5��	��h�ÊX��3E�K�:3>(#�P})Է�VAsW:�K"ZUt�1�ad9�Ġ6��܂ldbJ"A�������D�����ZL�'�k��9b亝��0�}�f�M��C	ўm���ߵ��!�6���66`0���>{`�����G�TI]��S�>��ߵ��O���>c���s�u.�2��++n;u��� 5umHU�� ��z�j���R[4Αm���pn�b�L���SmlE#��̡И�����k�Ɗ�ڶ�m�c�
HL��3U�&eP��;J�Tϭ��K��*E��/c>!j��ݺ���9���M�j�+�_���,�a-`݇��px�;u`i� ��Z�^� 6�t�!:���Fw,��ml����J]�v��xGFd�5�[�>��:�.��\�Q�wMr
�g�����s�B�u�<��s���޶�ũ�T 흶Lp`7���XH�ב������88�l�;�З	�BV2m�&KG�Αں��XtN��ZX�a�!*'e��jь�=�˗�8��M�9��� s�Sn2S�bM���n�'�&܂֮Ȳ��t;�"|��!�hU�X� Ͷ��
4,�F�ȫ�c*�0��-��v�j�H�6�v[�nڎw=<dPh�SJ�ܻm���[���$���Q�u��n~����o���Z��z�J�ZsO"��j���B�!p@��#ā�c��qL�[�OjϞ��!@��Y�+j�鸝Ԛ�rqҀ���R�r;��v4��nv(+�r��&�;cs�-W���K)/\����(q�݇���B�R���׍�6�m�d�^v$-psպU�y��6�e���tj��t�޽t�y��������m<b���搎؜vg��ڕ��A��M��*�@�jG/$D�f6�Gk�HuSnl� p��IM5M$eT#C��*ki{.�*�j��9�T��#ٸ��5FxַY����gm��h�UZ�ڶ�3��u��*��.�����]���{lv���7=�!Ӷ*�ɀ�r�;��+-ָ(�7Q'��؍�Q�S�n��+n�Z��k�ѧ;�7f��JZK-60.��u�g�dϭWS�5���ō���K��g)�{0&�&mE����RN���ۃr�E�j��!i�2�lϲk��s��p#	�a,������È�� @��hT~s�?:�b 8�����簩�b��c�8�p��l��i-��5 �nD�Zx\V�R;��s��TcO!KQ����nz;�.�ɋ��V]�NB��lai|ͩ�m�=�i�Blvtp ��.���inP�یF�i���Ԧ�g����9�����ک��p��ã��)�a�Y!
� tnl7lF��̘�= �AL�v6�M��+2`�q��w���mw�pVXˬ�l˶6�g�΄���q8;!�݄���&��k2Uҷ����-��u����,Ud�2*e4���(��%�;��� �͵��:�%���c��>Ͼ�5$R����O9$� O޸�MU��&vS|�5}�s�j��N��MЅ�Tn+ �nU��Թa{�^`���1�uUQɞG-�9J\nT���v�ټ���V�v�`o�6,�R��$�3M�r5�JX�����*����J��nrV�s�inpuۛ*�d(u��S$R�����ٻj�9��`w��U�έ�a��R� �{�ȯ}��� �D6)�E�r��ʰ:��l�O3��DL�oܛ��ADȜt�H�w~�`w�2����pf��塰��m��8��Մ֞`����D}3��V`�9Ȧ���E1ԕ`w�f�{6i`��b��U��p��L����j�J��OCa��u*�\���]�a�ι5۴��v�Zi��:)��F��EM�Ns�{vi`��`$��}�Hj��`^�#�ɣ��E�̶� �{]��
"ɻ]�`����}�̙���Т&BK?w��i���i�v�����lv�}���p��Q�P����j�=����wjkeә�i��54W*l�'�vg[���֪ə��eX��	��:�(	� ����$=�DD�y�`	q��;�`|�%��ٮ͗��ɽ�D�q�R�s�Mp�m�i5ː.����f4AէF.���M� f�V�� �� ��q`b�a��$d���8��Ձ�no7��mX3rX��n�<�7T��r��� ��ŀbj�Υ���p��~qStS��|�%�~�߾�w�v��f�aD/��J��g����͊���(�*7�s7%��<ʰ;��� �nڰ3��m7J�T�y��N��O�8�����-Y
q�4n��ޒ]�M��!n�JR�rp�{�`ws7�ٺ�{�Zܖ��9U$�:�r�US`u��=2B~�ŀuyՁ��ʰ9�mm�C�R�q�pf� ��VzgW�|��0�>E���)R�X=�,��U�;��� =��X�-F��Cr8��\�U���;�<˙#[w޵V��߻�w�R�.W]�w2�\[m��j0ck�Jۮ�H\��"8�Z��]
�ǋ��^�v.=����k1u�7n4�ѻ��,���^眤�m�$wK�30l9�1��ێ4�y.ȇl�H�L����$p%,��W���@�wsg�7f�Zy���w��A$��99��BV�q����m9qu�Siz3���5=�ծ��s���^-��A�1#���(1�ن���ww{����a�[��8g��=�O	至n���3u۳SFnݯ\�;uͰ�;.(�N����~� ��ڰ/���p��}�� F������8�v����C�ά����O3�2G�=�TB�N��h��8���}|1��t��� ��ڰ';���Gҙ,�%'n����=۽��gwZ��%2�����3�:d���1�RJ�;��0m�XkSV@n�)�3����U88驶���c�&�]`�[�F��l�䮶����px@��i5nR�v��~6ߟ���Xt��;�w�M������&�F�hr�E6Հ}���*�D)��S`f�� ������Rs�\���Õu�j�s`wZy��e?z��;�l��2~h�����G`u{�y�jn��15Q`vu.X[��ESU?8��)�pf���������v�u���� ~��'��ET�qZ��� 9�J�^��=�:;.�c@^z�g8&`�U"�	�t�"*��`w7-X�fr��I���~�Ł���TQq%�/�Erg��o�ZO0M�X�Z�=ט�H�*�mԍ�R;���\��{×U  �~F� ݯfZ�=Y�v���֢:$�PH�0.'[y�Su����^���n�}p�J*�H�E`ss-X�f;wۛ��ݵ`w������q�������F)��ts�Í������
G$�&��jm��j�N'$n(�S�\��j��� ��Ǣ>���$:�L�Q�i)
1�"#��;�o�~���߾�`{�>,Nnՠ<���\��2�D�fg���D��X��`wx��֡>�A����T�锣D��V~�����U��w�ʾ~{{�<�>��R@���)��+��lU˶��`�n�q�j�s`i;�57q7!��Łމ�)߮��ŚdB��VW���u֨9�Q@5��×�x��ی�V�jV����Xi<�SwkWgR��ͭ#n��#�	� �nڰG5����r���=L�nkܮr��$�	����mX�f;G����� ��ڰ9�Z
�$����Nqp��vu�����Xz>����_�E��C� cQ������pn���j���ڰ1ZQ�(�EQ�@���v*�\���F`�6�s#�=&�{Y��-�,+�.���1�vˑ�^R����2󺳪zVS��ڋ����g�O&�kf��M�;t;0/6슊�k�݀ym[E+ˌ����ct-/�k;��ܬ�S�]-\�kF]���t�<�$̬�]-AEF�bz���)Ֆ���N��n&�Nv������O���J~���d��N*�`
����nU`X�q��ے��X9��fm�ʦ�ە#%F����U'�߳�VSW����r��M� �Q\����)Ҕ�UVU�nE`eg��������V{���)��c�1�\Ud��e����Ӹ�3]"����ĊP�rJ�$�����pf��م���c�9����UF1��$���.,��u�,Υ�;���.;���8F�Y�=��q�[P��jQN�k�:죶��+ l�Fod�i�]�V�m��3���=�`{�n���Vw�Al�$m��M98���u�~���Z�5	4O;ﾹ�7�Ձ��`b�șUU���ƣC�����{7mXsr+���`o�kڑ��N~qStMV`���:���;:�,?}����p��"HFʥ)�qX��VgR��i���� ���9*I�&'B�M�m p̩�y $�g�۵V��M�p��)J�rSRȚ�V�J:n� �f�;�<�57q`bp�,�ު\�UEG$��r;�Q�i{��ݸZ�ܵ`,��;��Ke6J�R�u'8��,M�Y_�?�a��&BfByU�����@��B�Xad#H� A �B�NCl�df_�g�2
-��ߘkgNY�,ݧN/���"�0�{QE(��~���>��3�2�j���ɤ���ci�D%%%4�3(�@���]�x0�E/�|G��i�~��s�DL�DD2ACG0��ǈ��͒&L��9�Ȓ"""B�Jm�&	fE��Z(�J��[� "\2Y� ���e&π�'��D���}τLT�}��>�,h���RZSR�j	�ϛ���/�d�(d�)K8J�h�HO�J<�0��2O��Ҽ<�L�	� 0$8CA���_S�eN���JJB��h


T܁�������灂dᓙAFl���T��MJ�4��I�(� ����۷;�����;��R����E���)�AM4���2ii
&��IJY	����u2FI�u��p4��[�8J�B�ȹ4Do��@�/�A���ڇ��:��!X��D��� �'ADdD]}}�>��C���7�s#J��m��FئmX
�Y����ݮ�;�O0=�}��dXZ���
���*�˜1�Ղ;��� ��ڴWkrX��^O :���"��R�Rr\:ݶv	�-a;l�ݣk�s�{]aa�b���~q��Tq���ݮp�ݵ`�����.P,ǻV���ꑒ�N~qU:��f��� ��X�Jn �I�zd�����(���"%TqZ �}����eZ��7�ۻj��פs���ճ�uʪ��s`u�y�kn����-qDr&�fgX��P+%@RL�̈jE�S{�u�d�fDD��A�w~o�|���Z$QP9%IR8�U�;��y�=��� s���]�f;�-����#m�po����+�s�<��x�w\ŧJ���x��6�Q�TT4R��@���V�j�Υ�G�d���f��{�1\���t)�m� �{��JD%2,�����g�s�{7mX�Z
�T������ �M���20M�\ bn�Z���&v7I��6���������� �;��=��6gw'-��m9P��m�pf��{vX��y�`w����}
!L$��f��u2��U0���Yn�e�+r�)��r��7J�Oj��e�;\d7C;�>B�;�)x�bt��r6I��^�L\�&WO3�79Ď�L�9v�"m�cթ�m;�R���<WJ<m�gR���Q:�x���}���n�Թ�t��m��JڅMR������J�W=DZ^��s�Y�c[�n{;��60�4�lm�a��K�CSļ�%�O��eL���Np�Ze�)����͗<U؛��n��'\nu⭍RG�U:t�D��^ ���`w�2�u]��rU��V��n�q�|lwWA®�UX�77 w��a��� �ݗ��*Tg���N&�)�GRJ��j��;:�\Xku`wx��ӗ\㪨�a ��Npf���`v����ۼ\sO]F��T�(�+�u�d�S����`[��>���w���q�u�nMD:0l�:l��q<Xhvtml���r�'Bэ����qR���*� �M����. 17,�(Yi�"2~m��U#�;�n�B�	!!C{�w�p�W�{��W��c�7ۻ*'��"m��p{u�X&���Թ`w��`i�9QU©�R��8��ݖ��*��}���ݵ`�f�Z��r7WW@�q�8\nl �u��5�q`�Ձ��G~����v�Pn���	��}�m��rv�V�R{l�)�RI�봎[���⊒�m�3����	?߳ ����9���Ħ�ƶ�:j�&0�Bu'8 ��ڴ�ݖ��*����ndM����q�!6ڰ�����6��H�!�Q
?'�c�/��>��Ձ���["�#m�T�<��.76rb{�<���� ś��Ty��"���j�ʎ;����=�� ^u`wx��A�֜�MV#��p�Y��bm9����I"n��㒛+�����6��%���\�7� ��ŀf�VgR�i<��i�F:N�"F�{r+������o8f���z騹Q��C%�UV�����o0���MՁ�ɍ�@��:n�����w���Õ^}�w��}ZG 8���V������D�C��3vՀf�Q`vR\�;֞`������~�7N����"�M9��Ukt���C�:��9�sɮ���	��,�%;sW~6�wޫ������羈���q`u8�}*�u$�)G)˜1�Ձ��w�wZ�����J�Jj�395��i�s�4p&�l����{0��Xku`/fL,����G#O�&��s��o�� �����T��;�'� �|�U���EUUV���ٓ���owM����(�FrJ&����UnT���s�Gl;��̳���D��,�����ٕ��b�֗b����TI��z���>�tY-n=�������v���Jf���M��.ݵƧc�i-���2U:��I�ٲiz�Y�g;2=h(+�m�k��$���de�Fa^+��W5[�ݦr�x5v�`�n����1���d�۳=n&۲����!���q��ƿ�;�ǻ��<��7�!M��z6�g�F\�m5v;�̇S�q�A�\�x��VG������q�4A�?���n��f�ڰ{v+��X7p)��!`w�o0�����,�%6CR��S�"�UD!�s�b��V�;��`weX���n�Z���*�F�	��u��f{).Ys޴� m;�3��6R��qJ9N\�ջ��ｻ���j������K��R8��Z�u�۵��0j�{hN�m[t���3�x욲�:�(���T�����~� ��h�v��[�`vwslm̸���5�f��<���x��$D��8��U`F.j�:�<� i��8J*!�H�Q���ܖ|�*�U��o8�݊��i�cd�ʖU+C.�*�0�����,5��+���9T
qӒJ�{ۛ��޵`��w;3^�ytl�9S L��-K��\"W'��,".ݛ�tt��扺�h)���IR"*� �D�D��{wmX:�e��0�;�n�-̋Tq�S�Br+ �}�|7f���}����j��Dl�(�G%)G)˜;��癗�}�|�4".Q�ST�����?L6!o���}&w;ىƪ���	Թ�XA��y�&�ŀf�V�H���T8�ꟜN����uK3vՀw����a`ws7�|�*^>7��:T�S#�3Ł9z���@ɪP�'Gg�uɐ/<T�rX�MBQ��"F��s� �"��y�jn��z��2䊳�pr��j� ��u����, 1<��^c�GD�r:rIVw3y�ou� �;]����6>��r��D�R����V��K�y�a�F0�#�F�
�����E���I��J��KT;�,��l�����,m���UTUv�V��<�gu;���u����Es��)ZK��Nt����ܒ�u9��築'�n�́ש�`۸�G��H�:�7Zq̙iĺBu$�6�������'���Հw�l�3�0�>���$s�i�6��f �w �ʲfWU"��Zy�쭞j��j���(r���"!)�g�V�L�;����L�3���er�.jZ)͹m�g>,����`ֿ-�s�������Us�**�������P$_���9���Q��E2F%�" :� VE�D�$A�E1@Au�S4�@@
*2Ȉ���Ġ������U!�TH��R��
��E�	D�������R�
��E�T��@!�C�?����o�  �R(��������|�D���0?�(�{��(��O� �"?�QF?�O��o�����S��Z�?����_����)��������QG��?�����z�������������������uQEW��~�P JDT���߷�������@��y���_�P�S�TQU��������_�����?����l�Q�������y�}�3�₇�+_���'�������QHQ$�TD�E	Q�Q)Q A�RA��� "TIQ!�R �UD�YQ$IQ!!D�Q&D`�THTIBIUaD�HTIJHaD�TJTIaD�%D�aD��RTHRI IQ%HU!D�TH@HEIQ%@!D�H �@��$D�&TIP �Q)Q!�RQ%!D� JBQ$%@��X	��		P��$%U�� !%DHQIP��Q��X��		BBF ��		Q��$ 	Xd  $$%dFT��	 ��B@A$% ��	BBP���!!!	RB d$��	BBB�����&$BRBA % ��IHd)��$&B$$� d$RBT��`QHH$ HB!�)�(@��iBd 	D 	d%!		Ad ��� $!� d $	IBR�� ��BIhB$)��BY�%`(F�Z �P)!�"B@��!�$VP�H!	@��`	�� aXBF@�$	@�HBQHB R@�A$	BA��0ABA$�d	R��!%	B@��!$	aHXBXB	!�JP�d$	$	B�b �B$!@T��m���ߏ�TZPP�g�ю�3�O���_���/UE_�?�5�?��מ'��?�?��Ƹ�5���Us�߀�
 A��o������G�P���E_�y��X����A��s��,<����~�h�����0���]�(�3�����#���χ߁�TQU�3��?�������g�> �d��?_� ���~8*(����p�����⠡�?�����M�����������g?�����_��݇��c�/��QEWg��+Z�iП����b�!D����|�'���/_�TQU�a���PP�f�|>��(�����?����á�������d�Md$ɘ &�f�A@��̟\���@� P��   4  �x��$@U*�TI
 
 �^r�MH@����JBU�D��� JE�������J��R@�������P(�I�       � *�� ��f{���;�����9h�9� 8r��͔�ғ��{;׎�� :q�fΘ\�\  Mqo���������}(�{�{�����y�F>�Pa׮.�z�y�w�����3�aU� � �  P@� m�y��> =,� i��(�6PR�>�S�JR��@�,��
bi�8�J
0 ��
)�` �Ll�  ��i��f�R��t��)J1 �vR�7���r�R����)OM���J)M��4� �     .3@)LF��y�WU�wo�O]����{km��l�x�^n^{����\ ����}q���[�|  �<�ռ������Ҍo��u������\�U�x >����v���:�{���r��� �   
 � � ��L��5��rz]��)�E�����v8�L�� _n���N��ü {�ro�ԯx }<�Z��g=�י�z�#�׼ z�'�+si��]��� �z�  
 �@�z,gGNY�� ��x��� ��vuK�㽵޻�}���}� y�O��O!� �s�Cǻů*��΃'��{�����W����A�ww��]r\`�{^y���    ��*{iJ�  ���D�*� "x�T�H�  '�T�6RT4  ���j�*� ԥ4� h�OQ>�����������y�>��~ϵ����@_����U� �*��U�dPW�"�*�AO��'�_� ��P��SZ4R) �, �C�),!<���ʒ��l=��d����$�1�V5"1�]˾g���hB�(A#
�c� ��JR�,(Z�41��Z���73���}��!\"�D��F��F�o[�K�vC�u�Q��Xo5�48�5�0�ca�(�@���<�q�P܉�]I��51�bQ!d�1��%!&d��<�����	���Ja�R�B!cJ�����ů����qv�/n�!p	L=a%�%!LHԈ�cd�B��@�mhCXD���C�т�$}	V�ė5��!#�c$1��V0�"VB�7hI�B@(���E �K�q�icaBf�B��l���F�A�i#XŉXHSR�:aL%0bM씓[ 2�p�%�@����cF�r��PƘC3{.m�3�dbFR�\��-�N�BJXE$�X�A$
@a����y*�}�7��T�B$�������@w�ϗ�O�-o�!Bh�G��<�O`�D�2b�`�X�D���B��I�µ�M��be%)��s+�$��F���䋏�B�R��M$(F�X ����X#.|���_U��Z[_y��.h��/�e�
0&1 B�������}�7~��6��>y�da"YFن�e�a�f{=���U�Q	S#5�X�ZyuYr��:��V	I�r�k��>ڵ\4Ɠ�E)���A�Q*��_}��4�K�ҀI�|�X�f�vx�9$B�p��C뤆��T�D�d�R�8�0���Nh�!I3[e���g����;��b���4'	��4��B���!�Z�G�|��ZG�LBG.�J�0b���0��={v�T��\fs�yl̺�
���ϼʰ @��R5��#%���o�(�`��$F�0�.�h!S`B���)�d�k0�.��%3q�:��0�]]�e�n�d�r1�ÃȔ`e�1�d�-tx˚F4�]��B�d� i#X�hax{���,��3Y�u#_Sz�4±�aV!#@�V��n�X�]!(F�#�����J�BK�
`B�I(dCx�]�m3�I����HF}�F�i�$h0 �*B��
�S�Ƥ.�%�rL4F3PH�!ψT�%Ð,H�X@"D K�nk.�ܺ�V$BLYHo�k5�7 ȡ�5�F�,649�Y�P$7"����WFS��WS5�'1�B%�`\9�ƾ�$�
a�LL�� I`�M�H$	FW\�~� @�2��Gt%�D��!r2\\Hj�#M|C�&ͤlH�8F�F�B�b�<�	VbX�	H�F�R��A		 � �$$��T��<�T�R��5�D�ALL�ZB��D ��+B4�R1)aK�ki�f�FUĈ4=l.h��	���D��MXĎa�㠐`ԔaI]0�!�Ԭ.O�a��P9+Ϲ�_aL�ЗP�BOwY�u���p�0�p!S!dC4%�\4�X�y6�$,Sψ�&y8Ğ,)�=їC�0J���8l<>�H�"��U<cL�.a!�S��F��%P�C�O�������&@!�:07�̍�H҅k)o	�L*H,����	Iq-34{�zIHF;��$�e�Xa$��l�V潡�A���4��7�@�!	#<���L�|���B�hF�$d�e�e�2a��G�ov2ZS�c"{BE�͒�h�����y�������@�6�K`B! 0F����5���
U�|#01�(@�0����S(��I$dH���s���HK�['&NT��&�T���d�C�Oa��4��bmEpp�@�BbZ��/���\!๬Z��کhM4$!��ͮoy�_�IɎ��>��;u���q�8�r����#�h��1K� ��8l�w��wd�L`хm˸��"x���{��uƆ�n��p�m�sۗ{L�/n9�'a����2�۞{x���88��x�@b�wKfBf�[�����Z��}�6��F�^!h�b�e�-
cb�E�F�ںFL�R�v��ۆ�m��4mF�Dmw���7��!$��)�0�od{��'V��z4JcQ��v���0�i�[ɩ��C����w��<���*�:�k���RbRH�%$d��V"�abĒ)X!m2I�]�f�q��������O�H�#$ F"B1�r0��6����a.j��7d(H���!"HH2�X�S����r$d �6��.J�r�$M�.��	�:�,N$ED�F�u��Z�h������ͽ��Ki��Y�Y�*X�����G<�oC�@a��H�,!�0a�+&7��F���$Ns�S����PJbJ&�с�
ư����𙁠 �X�d�P��j��6��+$B��e�(II�)�B�F@(�Y�r��������D�+��B_c��0��Gv�k�N���^��:���D��k�k�|��m}�#iMk�u�bJ'�o����/�y�c�j]��Sɛݤ��LtB���!hƔ�fwJkb��q!�|�/�Br�@'�$�a� ZZO�sFN/��1�F��f�p�e֓9��������R8�,[���4(@����Onh7en|���b�CQ�!˄.9�/	���b�@���s\��-��$�E6��ʦ$Z�g�l14D��sQ K��XT���]�#�����!r4��aH\IrHRc�GR�N���pfF�h�H�	�$1�f�P�r��s�B�F�
�����)�(�$s߼/6��r�D�}�_$�b1�!Ĉ}O�����jy
aF����e�!3鿖w[�`i��Z��]���I%1!CaH�SU�E���x���b�}�ԾHO�|�sUicJU�)X�!I<�@��15�FH��0"�Y�M�@BU�M&$��r'������ދk��ߵ<%9���pؑ���GX2N� �䄺 ����=�!}��[�L߿|����#�!!	�B�8o1�B1#x���ˊ��y<JDG�L��"Hd ��6{w��B5���9&K�F�
ۘ��V�Xgs4M��iur�73,C�ˋK5py.��N�XիF7�0�,-9�X�|���t�����a���ra�1F���%i�0��T5���Q(�$Nj�J�9�m|;�9R��C]��ԚK�49P�$	_9yy�z�����@K���1��i"R!P�MI	���~��x����x��:7���`fE�1���J�@;S��p�ĺ�g�t�Q��.S�4�ܻ�a��1��*@22IX�`�!�	3en��)�0HDHb�#�t���-��w{�:�K䚸����r�^A��L� Ѐ�p#LacH�F����I~M���G<k���v
�"$`E�@K$� ���ֆF0"�,%!F!"��,`ĉ	���H�2!�FX@�$�\E"�Fb��O���ŉ`X����2\<�D���fr�s>�,��ĩ�	������ ���@��F�Y0�RhͲJ�b��i�"Qk���H� ���=<<<eq�
�5�Y"YhF	�0F`�	4�0�����1�	�G���<<�Bhy�HB���1!�jFJ!sj1Rc++-���a�'ؘ�$U�YŅRQ!"XH�1��`@���jH- 4bؔB%1���)���*(%�B��Q�h���$!4�	�����̈́��I�t��@+a��j�Di�˛9�y�Ld#W��@��<��RF�F" �)HHH4���������!�������Z��`� B�b%�[-��Ẑ���Q��
d(��L0���(D�$ 3KV�cؐ(�1�*xؓ�شӢ\$e1�"�H5��h�e4�(J��&��I.2���.�]���0��f-a	���w�r腁aa��7���ĒQ Ѐ2dH�5bBF#B$5 ��Ĩ(	ˮ�G��Kn-�BKT;��kl�ۭ� 6�� atۤ��j��k����+�H˵l�"��	۳��y���Ns�c����U�1�l�V�l��SרH���H/@U)�M$�)U���N�N׵���rI���5�m#��p�z��=r��I Vڷ��ѭ&��b�� 	�OC.� [��r�R�FڀG -r<�r���Â,C�e�]:���Ԝm]P��]�@���$���`p��o�[e�א�$r�$�%�1mュ]�!��{2�n�[Y*��R��-g���Ա�9��J+gh��,	e��k�g�j�A�C��eY8���-�S�v��a�t��Q�� 6��6��Z�j�E�6�M�H�bޢiT�e2*�V�R�M�檺U R�Y-�N,��讐�	��2 *���Ut�[t�]�n��[x �rۚ( 	6� $ m�l�6�&[@:4Q%�u�����`�H� $�K H Im�d��	� �Z���o��8*ڕj�d�'S�`pu�6�,�n�[@7m�o �6��Ln�4��fٶ�Z8 �d� �5m��N�tm� m� ѶͶT�H  � $�m� m �  l���� m���  �v@jU�N�j�V����>m�l�a��Zllm��Y0]m^`�!�6�m�h�mIvă�l� ���m�0M�^�V� [I6�6�6ؒCmͱ!��.�Uc����j[@�`6�� l�H���YYT9Θ �+UUJ�UR�̨�̶���6�" $[@ ��8�rA���uT�0����8  4RCm�l�Ko m� ���  �`հI���l �s�{2��)2�U�o3e�KБ����,`�����ь�T*�M��6�&��m��Ͷ:ڽ�͘� 	 �Z��mZ� 	Z0u��� [@�۲�̺��7.�WmWK皷69ۛٕ3u���u�1���)D��3�bGUUe��rp�pEq��]/��m�m���r�Fn�&��m:���{^�r^�2h3mR[5m<,67T�2�+�T��y�b����<�}����Wh �p�ZUlֺFe]�lB�˷&�j..�۶��wWi� �6�` �v� 	� 	d��  �  
��V��;��E�F����R�Y��UR��U$6�@[uV�[ĩ�
��C�UO*Ӯ6�˭kom�i����W��Blv+f��j�m�
@[PL�]ʵV0�j�� v�X�1�,�Տj�UOl�h�en��ۢ��7l֦ �c��G�o8p���촵�$=!�e�bJP�>�Sm&j� ���T�W*Ŷ�  -/^��[8�ڙ�i�a!��I����Ԝ�D��ɭ�[A�m��ݞ^��".�e@j�k�� �T�]*U�[[T��I��Z�!��q�6�ٶm��m���$���ʷTd�VvZ�U��enUV�r�UT��� ��6ٶ�����sibB(�8j�Yٍ�%��@�
   �l�d���H�ݐւ5�6,�%�V��g�	�̤��m������eZ�`KDU��VԺ��.�^ntT���[8����i��gy��ݞpl����;B��h���U�1�Pq�Rtr�7Q/U!t�q�'K]K�(�B��G����r{l%l�n��Iz��
��Z�\ձ����h�z�k���r��@�$	� ?o�m[hڳ]rDL$٥�F�	�]�T�Z���P1�n�A5Th��e��	T	Yy�V��j�V��)d�p�ͶhR��w�}� ,��I	����g`6��mm˻���Ed�)���3����m��Leʁx)`BV���� i���l$6���l� )v睡̭˗i�(
�WUJ�*��i9���,�Ub�ݮ��T����EV0T���J �h�+v˻3�[���Fݳ������m$�i^P�kN�^��>]��m�A!�	�bA����U�g@l�\�M[<X�*� �V��+V´U/-[�� c=vu�#B�о�-�oh5U�ʴ��J�@��Cen��G�V��%ތ� k6]t�)R8��� ��t��uv��n@�Y`-� H���J �S�mn  -��� I��m$     ���������[v�SI����m��kX�ʭT�)-*�Q*�T�J�ɉ]VҦf�!��Mn$��n����'mUZU�6�U�*�[��vں�������F��jU��
�] p��﯐���Q� ���#	"^[�	9�mLȮm����dyz��걊�A �m,-�܂�� *ꠥ�ح�c���c#���v�vK�m�wÛ�?na��(���(]�hm��aV7$�MףB��{h/*��#�URZ'&U���{la�`sq�T:*���*��r�:�f���hԯ-[m;��PE	��j��YvVq5USh{l�\�hM��]�t���y���u��U�W���X��旴���ۢ��%��'i` 6� -��sn��9X֮�*@�#���@��N�-�  6ͤ��v[��>p�6ֺ��K� 6�E� �@m� �#m��*��(
Kl�R��Ua�� ��OK)��mN�h��[�m��H 8 �ȵ��֝m�d��[KV�mH � �{{t�i���M�s��m��
nR"�Ulm@m:��P�Cm�l�Z�|�P�s�lF�Xc�a�m*��Tqm���ωe�}kb�L���hk�\
�Z��)��B�ݍɮ������Y�pB������l�{TcZ� 
]�Z��W�jV�T{c�Y:Ytu���T�lj�ݰ	�]��l�d� ,K��j�*��A�u���f岖I8�U@�gJR����er�6ӱ�,0��]v�s0]S�{GnI"b�
nI��cc�ճ��0t���UWKvPs�=qL�9���r��Pv�UX�15�m�*�.UXO�９����3uˬ.�-�W����pT��o]l�ʶ�UmS���*��3��R��@*mV���3�9M%/J���u��Yp��� 	+�d%���m�v���!���V��;`U4�U䳵����\$-�N�\h9�ks��m]P>˯M�m�,�J��8��v�t�T����ߚ�p�-6�V�F�n�4V��*�A��6���^�^��]q�� *�ճ�2�Rl�Baj�A��Z� ��`� 
��U�-��ԫU��\#�Ni �h[[e�l�`[��Hm��4��'3�Zմ@m�m���mWS�˷++ی�    i�v��M���
Te'l's�& �  6� [C�E����� h� ����vm��f*L��2�ܐm���5���ذ�/|�t���nē��.µ��J�UU{�-�T���!m 8��"��\ �k^�AK��ʀ�7(d�f�M���GU*���    ��khm�m[�m��|H{I�l��Ză���}��-��i��@m,�Y�7mۀԉ6݀[@�M�a7J�&�� �� �۶ZLѹ�'��"j���c��:I�9��]�8v��
�m��66Y�Zi��RWE@�z8�U�"����9�r�ۯ�iV7Z@��m�Q�S��d��g��GKAaE�[x4t$r"���I�gm��ր	�m*�[['������y�Uy���y]���l��H�  [c���� U+��U�R��Hږ�-��6��	oX�v�m�I�jt�&�,�	��d2�ف�j�"QV�v)�&�`     ��     ��cyK���ڲK��D0h�2ȖQi� �  ��!����� m AD���R��b���$�θ��UJ�ʴ49i	Bj��B�]*ʵ�i畼�3P �d�ګ�br��t�9R6�6��7h�lN5�[R�D���m�	6�[h��T�2� ���h�Vہ��$��8$A�u��3�X��X�%�]�E�<*�R�ӱ�j��;��ym�V���7�jS1��\�/Hlڶ H6���t��'EK@��]*�������8���gE Ʒ��P� ��8y��յU�@mղ�ܮ�4jUvU���
�F�ƽM�		:�ր8,�8��[u�mI�C�!K�I�(���^������+jk���,����6�-�2��[v� �E�����PكI-�!�d��m�$06���mf�r�Erñۢ�$-� m�MM��ݤ�e6ږ��m��[  �����ۖ�8��d`�-��[�hm�۠��$8 u� p<��⪕Uj�8a�!�p��kX6�f�*� h]6���Z886�L�f[��\$�����m�����aN�H9��ͭΑ�e��a鵮3�����J���I�zÛh� si��dŲ��&��gl���!Le�'�j�Rݔ��Tk��P@�+{v�x
�5k��n�ɇKҒI�6����� p��	-��Z�Z֤��ˣZ����*���HlTj�`꨿�R/� �h`�Ƞ3��T�W�.�����=��@� �lGy���4��.*�����4t����� x?#��68�HёU�F@�*	���"|��`Ca=6.�_���j0M���؈ ���(�U<=E_W��^ ����G�<~P�O 8��F�x�"mV���D6�;}/W� �M"���h� ����!���8��:UpH��>v���>���,>QO���DJ�hUL�	q@�P�H��R���G}�����0؀�0^h�Qg��F�������(B-�	�(�f��EQ"�HD��+�� �� �&>�o��|)���&�"�H( $4b���x�������D�C�_���ુ��l�&� �ł��>�G`#��H�^)1,I(������Y C+���F� �Ac| Ū�x�a=U�"/H���X��-A x q����
��=Gh�B+�ȡ�$3pS6
���] ��1D�J����kZ˓2�Ŏ�$a�$V8;rN�;[B�m��P0��[B�9�u�4eJ^m���mluv&�[OM���3����$����d�&��J1�;AEc��:vW�w��A��:�a�U��v�%�e%JKT�N;4��K��Ը�`��) �QĶgD�m�8�*��:���m*��@��-��l ��:Uݙ�3��`�gDE����,λr^E��mk�9��[mgm�GH��f��Q�6%�j�U�J��Uu����we�N:�ƥ�b���i�=Q����:���n�I�bLun��k ��QM�lCq�����9SH.��mєu\� ���M�5�Ί���u�L훘xv�'L�<*]��G^��; ���9�b<��T���D	b�G�L�Mfs�YrUK��c�H�Vk��M��3^@kbj�'nY�]й�6K<d��l����x�ٞ(�����G9f��s��hR$������Q/J����ѻKMv��g�L�N�v�M�qK�ZL�w$j\�;-H�,�nŸu��u���,m�#a�u���A*T��`�\��퍲�J�۶��m�V�#o]6zH�N; E0/F�s&��^��4❠#��ru��c��l���e���닮o6ڷ��3�X"�q��gn�����pE�h�"/l����B���5W����A�M�r�2��v2�0@*��*HUj��T��h9QL�4�ڵ.Q�v8�6m�m.{G���MU)-x��/2��2��{t���5��zԦ��v^g6��v(�z�F��v����(�*�S�M{ m[^�m�I���V�]i��D$.�C]rS�H�K{q
�"�/Gg16M��k"�gV˲=���^�P�������
��8I/�)�!�Y-pPf���O��Q��R����)����5�5�y�S����_F=���]���v22s�\���Q�'Ax��"���_W�S@�����D��'�Dv��|!�  |#������m0�ݫ�u(�Sschwa�'ds��J�9�Xݬ�J�[���=�-d�t� ���An3�WF���M�\s�*�g���/ �#��)L=5!e��#�Q�!랽dN�η��U��k�ۃf�:D�v&e.�G9s��l��"��$�.2��9qN
wf�5���d�����rK�Z�m/�9�c��<Z��[9Ѓ����x�}��v�� ro ���2<�����g�l��x�y7.P���{v���Mǐ:�4��@7��� =����[���bd"pRM˭{�#��~�@:��4��@��uHL�&,���MǠ}�X��l���˭z��'q9�Q�H�$Z�hu�@��^����hu�&,�C$���l�<�נ}�,Z��n��b��{��7`�����.Z��̸.;K<���`-���a�7e�rt��5�ޠ8,nA6��W��}�,Z�hu�@���@�$k����{�}�`m�!$I0h*%�cͤ�]���i��4�s�@|�k�=�PN�'2c�LnF�.��[f��ֽ�ek@;�R�8œcQH���@��^�޲��yu�@3��U�Lqɠyku�~�n� ��u�ۼ�([��<����S5Ӹ�ͤ���/Ohlnms;���'3i���wl%��r݇NR&��_��Z�Z���@��^������D�"pi���ֽ �l�<�נ}�X��$������8�l��4�{�@|���ś���K.�EH#L7���sWrOo����g�9�� 8,nA4��<�נ}�X�.��[f�|up���H����u�-˭z�٠yu�@��醲�����Q'k�r9+�Z�����9SE��o[l�Y�U�3ێuc8i�u�1�$�-˭z�٠yu�@���h�ζW-��G]�@�{u噊&M��X�_\��n�j=�n�QT�j�K-�>w�@o���G�I�W�����@���,nqDډ����w8�[� ���(��I��$3f�|w���r�����84�@��^�u�h]k�;�V�z�����mܘ�q&�D���]k�ۅ��\��'�^�0h���ۛe�����,�d$mI�u�h]k�;�V�bK6Ï����Wd�J�F����t�Z������^�u�h���L0���7#�;�V�/uz~���H��~��~����'c�1c&'&��p:"!DN־� }�x��u�~�,Z�e��Y$M��@:�t���֛o|�^��||��m�,Ŵfb���4���v��	mJ��;��Ƈ��q�^��nwn{(F�i��;F�=t�c��������uq���4Աu*�::lX��z�#lޅ��o�6y��j֞�x0syw]s���ŰEp]����i�K'E�m�vg����5��	dP���9��:ƹd�I)`q�r-�������f�\�[��΀)U�p�\�;����A�T�l�9��X�gës�h���i��C"�N��˲���'��ènM�I%߿I�$��/�I.]w��]m�|�J��Acp�M���jI/���K�]ǩ$�[g�$�^�MI%��N�s�&�dRcNH��$�u�z�m����m���t�o|�^��m�ֺ��N�UIdn�4����,�$�뽶�]����K�b����q�I%����J�9i#��m����m��w]�{m�>wJi���{۽�߳U]�Q�&���e��[���Q�7�:+���`�B�X��n.�g�v
z�w=)�-W� �;�z�����)��o��o�,K�m�{���K֚'�cncŌ��$�}�Ir�홿<�dx��0 �2@�! � g
����s\嶷���6��;�׽�33��B��u�`�H�J71�I%~�>�$���jI.��}�Ir��$��yu$����"N[�����I�z�6��=��m�OCI/^��H�d���mD�sRIw���K�]F��^�g�$��k��?��po��+<����u��ub�a֭�n�Ů�:�j3ۘ�1
7x��#����Q�$��Y��$/Z�����M����u���UnF;Y��K׬���sRB�]��$�s��RI,�����q��'�$�^�MM��w]7��bWma�s��OM����n��V��^I��#k���&������K��ũ$�����K�ɩ$��Չڤ�DԬp��{m�rwI�������m���t�o|�om���@�u�r8Y̑u����v��$�/�\�����Z�6�;0��
BԨq� �����|�Iz�5$�޻O�I.�w��^
����l5�� ���_~���T>��{m�����m����������_Z<n`�M6�nI�$�߷���$w]ɩ6��s�{m���m�m��u;.YUp��}�Iw]�ԒK��>�$���jW\����H�����s��/�a����U�m6�}�����)9�[��|�u�{m�s��i��\��9�X�F�uu�+ �瓨uzyѧ��n]R�B@RS����ڹ,���0���� %�dԒ^��}�Iw]�ԒK޶}�I[�9VI��#k���&������f6տ�CRI.�ߧ�$�^�MI%��5;�����Wm7���;��m���n��Iz�5$��v�|�E��Z�"�����$��l��K�ɩ$�����$����7������r}�I%�dԒ^��}�Iw]�ԒK޶s���B�@H@���B"�~}��qW#�u��䠢��:sغ�0l��^Z�c���e�q�'M���In��Ee79knF�㞑4�ҷ\uh��z,�=;9��=�4���e�NḢ���4>�N���&c�,�=n��暜F�M�m���8���� &.�yb��r@D�c�U�{EwmR����x���ٮӖ��5�j� ܩA]��ңƹi{��Z6nyi'��!*�;���7��w?b[ԃBqm������ܮ�,i��)ps��E�5� �b0F{n5�\=�U)�س�j&�I%{����K��^���I/[&����.���b��y��$�u�I%��_�$�^�MI%�]���c��u�*EU�m6��}���$���jI/z�>�$���jI%�v<w�dq�N1cn?�I$�l��K޻O�I.��K�ֿ�I+pd�YBKm�m���om��3���m���zom����m���QˑP�J����N;]ms��v�֞��ny �was�t�]ۖ9�1��71���$��$�u�I%�����m��{o�bX�#o���om�y��	ar��m�>�f��bX��  2 �
�M)�Į��v�6������|�u��m����ԑT�to+�om����m��]��$�u�I%��_�$���XLM�Lq�DܓRI{�i��%�wCRIy����$���RIy�\Q�Ĥǋ��>�$���jI/?Z��$���jM���om�垁�G��ʂ��\9�	�si{���/^ىt����жš{oʘ�^���@�m@�$�>����I%�d�m���om��wZ6�{����U�'#�)%��m��{n��b�7�{^7�۷��jI/?Z����cm~��'�	�#�!%���9�x��o��o���@%�U/�bB	E"0` ČX�A��L�H�HY��Sb�"`��V0wpI
E�X�qW�B�`A�HH@ ��0�h�=g�f��_p҅ZI(d�kX@�ac
X2�ҖFA�KJ��tҏ��B!!!	D$��EH�	 �5��=9t��w5
�����h`e���ժi	1�!v��F$#t��+�FC�!(G#I$&	�x:7ǫt��=�jC�%"�=����Fs�0����
��(HU����4pG�;:����PAM���U_Q��ө�������T�H#�f�﹜���k[������֬���Y%-���s��i�����om����m�f$����{m�������N������M���t�o�ݭ���u��m�)����?v�G\u�e9l�(<V��;�u���n%o�:{[e��stݷ+���zY�?��o���m�ϻݭ���u��bY�	}ku����,��&'&	�1��Ǡw�Ŝ�d�w��ϫ s�u�|�B�:Z��MՂ��t�T�������=/]aСDL�����b�6}�������u5R]ف�
)��Հ�� �7�$Ѩ"�}��D�����ƀ~��O��#�q�q�{��?/�(K�Q��^���zwf��ދ�:n���d��6r�Һ��nxzw����a�ւ۶��U�GN��~{�]�|�r�iO4��~~�� ~�f�z��N������ncŎ!�I��4/Z�
������;݊�2B,cI8h^��{��=�)�_t��x��[cy12	4��*�W�{�S@��M�ֽ ������&8ʕsWX���v���;�X�=�7$��=�@��ZO�u��Yp����vb艛�c���)]�6'�$wa��q��=w	�p'G[6LD擮�V��i���a";�5��>�e��l��g�m���,3U�\��Vl�XbDݙu�l��ܛ��c{;zԑ�-��+I��l&���g&�$���@b©5�t� �n�\'k��vݺ��)�m�T���Fp����4�;7k�Kq�`HìQ8R9)!{�������D�6Qn��,�����,�Yes�o�9U$茶�H����Q�ĞFy��~���@���@��^��YM���A	��ӑ�C@���@/��޲��Jh����x��xۏ@/��޲��Jh^���)^I��#k��$z�e4�)�yzנr�^���:�'1���$��ץ4/Z�W��=�)�{�e{��m{^4�<H\�'b�2��hӸ�5�kY��n�u�c�H,ナ(�q�$�yz��6^��=�l�DG����u�Lo&$���Ǡr�^������@�Қ��{� �U?B"I�n&�e������m�tL��u`����\Q�ĞG�7��hzS@���@���޲��,�4��Cr%!�yzנu}V��[��u�M٘���l*�I$���tR�-���'�\��f%��{	�3uH�^^n�f�s�k�5WE*����}8���m��Q�>{�@yyu�L�����E�h�׋9D%#�|`��e�䒉�����'1���#��_�~4/}�nh7�d ���R�����V~��� �Qe:��X8ƒp��������@����y�X�D�y� h��f�jmL�ҙ����5ֹ�>_D$���/�u�`�?����~?�����b�acs3�v��P䕺���Fw�S]���z.���wx~:� ra���^�����Jh/[\�BQ�S��7h��n��ک
�sV�{lϔB��BQ���}X}]���x��P�$�M�+�Z-�d����0��]k�:(�3�݋ |� ��jiū��*��UUu��
%���u�,^�01B��	'�J` ��N�3�w7$����q֌�kU()\���kŀr�}���=;�X;;נ?fff'���
�*v�4Җ�X������\���+ �n��{Z�F{:�}��<���Ncǎ!�)3�~����>^��]��g�;����\��DS3V`���|�%�IU�}���ذ�S$0��mLN(7��@���p{^,>J|�Uw�_��������"I��������˻��@���z|�`}
>Q]�wӀ6�{�5J���f��.���m�В[[�_�}]Ӏ{���)D&�	%@�AIֵ5},<
��;����(-"���dL�@�*<ې����`�nٜx�Q	���$����:�:nʽ�]�iSr��Z�bt�nΜ`գd��j�gZB1Y��.���$-I��\�[u�l��k����;�1�Tţl�7�v��L�x�l�۶�eP3�RA��$�$gVY��s�Mˢ�[$U�u�vٕg���}|u�v㟟w��x;o�G�8R��"�z�jE�WWm�����c��_G/e	��6�H����GF��k�F���ce��`�\���]	/�����k���ԕWe*���5ֹ΅2n�ŀ>w��|�g%	L��9���U!wR�������`�هD$�S>�������h�"'^D�<x���4?�!D|�Q
��|`/� �M�BK1>s����QI�IlmXX0���|�`
#����n�ŀ?Ss�{�����	K;6��\9��5g���G	קi����ئN��ˀ��~���[�}��p�eT\���9���=�x��nz!/�]������8�&L�<dqh�]���`b$) �
�6�*lJP�EΫ��W�%�,�V�pK}Z���ױb��r�l�\����\� ���?O��>��QU�W}8}�-�x�Xh�а�r���=�?�=Հs�Ӏ{��`rJ"'��� 7ds]����]��� {Z� �/�!C}����������@������4˞�amIv�h2Qm�qj�Cr�{/�jJ��F�,w�1`��Z�j�-�U��9�i`������D$��u�8됺�W5j�*-UY7k {M�|�>�I*�e��`uwӀ{��gB�	L��,��*(��&�7��߿=�i�ə�*���`�� r"� ���"����ٹ'����rI�Ns�FGS��&Wl�ybI'��y�q�,�n�:B�V�V 1wu�J�����Ң�� ����:%�ϫ����@��ZY�X�Q�d�dIc��#����<���m�n��r��z�ns�c1_����dz�O��Hm�Ng�~_��|�k��sД~��}� ��]A����(��&�� �>n��B�;��p�ذ�W��?�:����x��xۏ@�����׋�"#�U���Հl���SG/^Z�c��ŉ��ր��{��r��ٹ!� �(E`�`|DJ{�K��{��Mgi��3!E��&�`[u�|�G�
6��W���� �����ɊR�]�.些6�k��Bc-�=�)s�&��e�[��6�9#���0s�VG$K�hm��]���+�s�{��tDD~���Հ�M�諸��\�� �k��%
d�}� ��Հ~�7YТ%2]��T�VUrE���� ��9%	Dϧ{� ����@���R���������fb�BQ���V�����\�|�K�C���٠[�Y�a�Ģ$1���z����!}w���`[u�(N=d��_11 c#���i�`�ִ�}��C_�G�C�x&��Y
)��!�d���q ��@�'��5�#@�dBHF�$@�@��! 1!		1�D�Fzq�
F�ZD��HĄf�b��H	�b	r@�
+E�,�d�mee%e!HR B0�d�D��2B	(�FF	�2 FHFI"$	 0"��A"� ��d�H��� �$I�&Cɠ��B Ń �TMx2����`!p`8xj�%����b1�dc!�J�0b�R1b�,�1S�,�J�(A�#HA#,a�B�
��8��)���%�Ĺ�>�M��I�PFXV�%
1e��m�X��v��v��h��r�)q5��X\���)�me���Q��X�������R�֗�.Ú��Sƒ܀��l�8��9�\<�t��]��ۥfL�6[�h�qrL)����X�6�WfT�m�g(��������G��:$,�2�X�� N�dCU�m��8�ڔ�cJ!t������;*��kk�1t8bX8�yۃ�v�q-���=<2�۶�絷c���n�_��c�yZ ��ԫR�5X���:$��,�mӄ�,طF���Z�Ŝ�p�p�3ĩ3�BT����N]t�Ú��2���LI����Il���s=��"���ų�EJ���]K����o^�om� ĝ���3����=q���;�Ah�$m �J�vb�m���m�RKə_#�� sK�ѫC���C=�=���b�3���'l:ݐ55]+N�4l�1A��Nr�VUSsk+� !�Qi闝�Cb�L�������Em'Vn��Ŷ��6��7[1�zx^!��'g/+�n{Q��zp�!omq�T�U������ h�v]<�-K��Ux�ݚ$�Y]�ck�Ey-k]��ę�c��㞱xP�C�yᇲc_g`�b�jݵju�l�6λ���@:�<`ڨ�Ƶ��d�2m^x�[��K�T���-��ͫ�iJ��k���3�������[9Y�Ė�o���.�'ِ�/Ru�BZ��
&iUM�Nn��*һ V��7#��86)6�匆@1��뵶���&��s:݄#���3k��t�"��c�=�:ڬ���4 wmג��SW�P��a�db�­�ڱ��n�:AS������S^��uʲ�R'ɓ���H
�֝��.��F�)���S�	�mG\n���LjŶk�{G���1v�Wk{k�h�]������7�u�Q��Y������Ub���홝����F�u�K���Lu�GkU��ؠ;;��8�#lY�n����n��������q_D^���'����"����U�Ҫz ��|��|�Q���,��k0ԗ.h����v���=\9�v@P���P�b�u]�S{S������>�%�7\>4��_�?o���P %s�LL�����e��vݫ�ʉ�9A57W.2i�g;�`b��0��:�3�Nk���풲m�c�����o[�S�j8�s����l]X����S*5�V�=u�;j�`��I]m�ȓ��Y'Zm5;-�:).ɬ�@@��7�M�˚�&��Ip+]"цp�:�h��	���t�؋�%:�:�;]#��5S�ʬ�9QI,���~���- �뮈�!���� �.�H]ԅ�����Y��*�����e��`]�@��aXӘ��&7&h[^�9|���B��Aș�~��6��bX�'�w��"X�%��~!����k-.�2ٙ�ͧ"X�-��{��ӑ,K��u�ݧ"X�%��w�ӑ,K,N�{��r%�bX��}�w3%�YK��a��ͧ"X�%��뽻ND�,KO}��6��bX�'s��m9ı,O3��6��bX�'}�v�{��'uGGt��A�ػB)�`{1�x�Qq8��Xn5��?{����m]�Y���Kı=����r%�bX�����r%�bX�g��l? 0O"dK���]�v��bX�'���������e��j捧"X�%����ͧ!U� ��:*-o�*�dND�5�s���Kı;����r%�bX���xm9�C"dK�ݧ�*n��HDKf�l��L��\���m9ı,N�~�m9��,O}��6��bX�'s�w6��bX�%�}�s��f���F���r%�bX�����r%�bX�}��m9ı,N�{��r%�`~D�D�]���r%�bX���~yj�-� ٬[1313�w}�ND�,K�w�ͧ"X�%��}�siȖ%�bw;��ӑ,K�w�:�xn�� J&�
���.��D��w5���:�-��ٛú{.�6���㑹�2h�&f�ӑ,K��w�ͧ"X�%��}�siȖ%�bw;����@�&D�,O{��ӑ,K���x���Ht�i�����{��7����siȢ�bX��۴�Kı<����r%�bX�����r �X�%�}�{��2��d4d5sY��Kı;�}۴�Kı<����r%�C�q
�� ��bw;�fӑ,K��>����Kı/ӿwF[35&��I�.kiȖ%��(��=��~�ND�,K�~���r%�bX���w6��bX#bw�wI���{��=%�E\�K,A���n�H�r��ٴ�Kı;߻ͧ"X�%��w�ӑ,K���;f��r�����
�9�[�QhW�lJ� gun�Ѓ̞ۛeL_w��������n����"X�%��{��ӑ,K��~�6��bX�'���G�,K��w��l��L��O�}'��r�Ii�ͧ"X�%����m9�,K�~��"X�%���{�ND�,K����bؒf&bf.�k�-Q�t [n��,K��߻�iȖ%�bw;�siȖ-�by�����Kı;߻ͫf&bf&b���椕F�J;V��,K?*�"~���ͧ"X�%��}��m9ı,N���iȖ%���#"agbq�"w���l��L��_~�kS�6��FI,�r%�bX�g��m9ı,?) �����O"X�%�����iȖ%�bw;�siȖ%�b{�);���,�fh7[�Rɧg��e{
*B�
���k�zݖ�9�ԺĐ�jj�*t��U�5�f&b�,N�~�m9ı,O}��6��bX�'s�w6 r%�bX�g��m9�����Ow�F��ڂJ�ų�bX���xm9lK��w��ӑ,K��=�siȖ%�bw���iȩbX�'���w,�ԅ�k2\�W4m9ı,N�~�m9ı,O3��6��`��bw���iȖ%�b{���[1313=�E�F�j�h���fӑ,KlO3��6��bX�'{��v��bX�'���ND�, ,N�w�X�bf&bf'ýs�U9c$��35�ND�,K��ݻND�,K�C���i�Kı?g��ͧ"X�%��{�siȖ%�b@"�v�������d�b�Pf烱P����k˗�S<��KqԪtXnh���d��=v�n�� 9a�t�u%��5�%���k�K�E�WD��E\N�λ��[���ة͡�ȝ���ۃ�E3-��=�cX�oآ�jx�+]����zt��am9���p�ڹyh��4V�Fѩbn&ی�'YD��Պ�wt��4ݡ��nKx�0D�<ѸA��n�w��{���ޯ�s�5"Z���qlM�<][�5�1�Q)<���q�Ӱ������WO-Q���Ӯ׬[1313}��[ND�,K�߻�ND�,K�������Cșı?~���iȖ%�f.w�5?:9U�
���k�L��N's��m9�ș��>���r%�bX��k���Kı<����r*ؔ��_{��O:Kci�F�%�ų1X�'���ͧ"X�%����ͧ"Xؖ'���ND�,K�뽻ND�&bf'�ӳ�(�S��AWl�-��KV��>�siȖ%�by����Kı=�۴�K�A,O3߽5�f&bf&b|;�Ur�K*d���ND�,K�~��"X�%�删~���i�Kı=ϻ�6��bX�'���ͧ"X�%���M̷2K���m[
�\�3����Yf8�k�h:��u$���n�|�q��X�dе���j�Aȫ�i<�bX�'�����r%�bX�g�w6��bX�'��{�ND�,K�~�ֱl��L��\�u�)Uh���5v��bX�'���ͧ!�Z r%�b}�w���Kı=����Kı=�۴�O�șħ��g솋��35f��m9ı,N�_�]�"X�%��w�ӑ,�,O{���9ı,O3߻�ND�,Jb�@��ժ0��+���L��ȂdO~���"X�%���~�v��bX�'���ͧ"X�b}����r%�����΁��I*�!T�v�bىı,O;���9ı,O3߻�ND�,K����ӑ,K��߻�iȔ��L�����[,Ei��-v����-�F�Ln��'y�s�3��m�-JX:��u�o��~���Յ�����f&bf&b�s��Ñ,K��>����Kı<�����%�bX�w���r%�bX����;b�;]v�bى�����;�M' 6%�by����Kı>����r%�bX�g�w6��6%�b^Ͻ�d�ʙ%r�bى������}�iȖ%�b}�wٴ�K*;H, Ҁ:^m 2&D�=����Kı=Ͼ�m9ı,O}�w��3Z%�k2\�W4m9ıB����iȖ%�by����r%�bX��{��r%�b؞{�xm9ı,O{���HJ��[#r�ų131}9�Mb�Kı=�����Kı<����r%�bX�}��m9ı,Oȟ������:�z����+/kAmg�76وl��\t�a�o=�<φY�p�#l��Y��%�bX�g�߳iȖ%�by����Kı>�����bX�'���k�L��L���y�TalSY��r%�bX�{�xm9�,K�{�ͧ"X�%��{�siȖ%�bo[��_�_"(�D)!7�e}6UZ-�35.�m9ı,N���ӑ,K��=����K �,O{��v��bX�'���ND�,K��o�jf���ɬ��5���K�lO3߻�ND�,K�뽻ND�,K�~��"X�+��������fӑ,K���N�X��N[��٬[131X��]��r%�bX�{�xm9ı,O���6��bX�'���ͧ"X�!����������g�B�)���'��\	�5]��s�ъ��[9��S�zw�o���9��9�Q,��W�_��������bؖ%�b}�wٴ�Kı<�~�lQ�Kı=�۴�Kı=��v2Z�-��*�Zų131w�׍'"�bX�'���ͧ"X�%��u�ݧ"X�%��w�ӑ? �Ȑ��]��E��%��F�5�f&abX�����ND�,K�뽻ND���@��=���m9ı,N���M�"X�%��}or.k�՘fkY��K�@,Os��m9ı,O=��6��bX�'�w}�ND�,K���k�L��L���y�TN��Z�m9ı,O=��6��bX�(��w}�ND�,K����ӑ,K��;��ӑ,K��sϤ���{�R��v��v�Bc��a�݇h8��d���m����-Tg����ekU�uRxz3����&���=[���:�;pC��}�h��"��V7�vՂ�r��z[1W=VJ��&ub�6y����������۪[��6[�P}�ENnA�9�m�Sa^��������ή�^u��u\]x鍘z�gͨ�-��lcA���x덨5o��-�-�{���(M��8�%�=tzP���rh����GZut:��M��}��8�j�QXIGj�-����b}�w�m9ı,O3߻�ND�,K��{�ND�,K�~��"��������SҒ�ڲ�۲�X�%�bX�g�w6��!bX�'���6��bX�'���ND�,K﻾ͧ"��,K���~�rh����]k6��bX�'�����r%�bX�{�xm9��,O���m9ı,O�;�[1313����"Z�eL���ͧ"X�"���w�ӑ,K����fӑ,K��=����K��!S"w_�~ͧ"X�%������Y-C��Ir�bى������kư�KıO3߻�ND�,K��{�ND�,K�~��"X�%����ߢ���Ծ���z�jn�f��%gi��Xק�;g�.{:S��3ӷ7kf�S��ӑ,K��=����Kı>�۴�Kı<����"��bX�'���6��bX�'�}���h��.f�a��fӑ,K����nӐ�~"���lX� �#�FaF2�~b(G�<@Jr(.
�vH�H!"�			�|USO�2%�bs����r%�bX���}�ND�,K����ӑAD�,K�!���іj�&Xa��]�"X�%��w�ӑ,K����fӑ,"��\��=ϻ�6��bX�'k��ӑ,K�������R���լ[1313y�zm9ı,O3߻�ND�,K���ݧ"X�(�by����Kı>�V�����Օ�ݖ�ų130�=����Kı���nӑ,K��߻�iȖ%�by����K�7�������\Zg�<k�E[2�<�oA�ލ��{�cn[����.���,��9S��AWl�-�����������N%�by����Kı=����~ �2%�b{�w�m9ı,K�oi��KUnB���f&bf&b���֓�,K�����ӑ,K��=����Kı=Ͼ�m9��"d��]����Z�-��ʵ�f&bq,O{���"X�%��{�siȖ0�dHET���lH�ZF!a������al0�� ѥG1Ҝ6:��;B0*�h�*B���FRR4�H1�BP��B��)a���BBB)�(̉�`�,�1�Q�!0�đ`�K@$5T��rJ�
�JRH2�B0�a��P����C|���ں��i��X�AOw"IHH�5Y
#���^/������p]D~<D=A���>Ч�E>�]}�.�F�'��|A=BD�>�|�m9ı,O��xm9ıL��wMz�
�h��v�bى��%��{�siȖ%�b{�}��r%�bX�{�xm9ı,O>�xm9ı,O���{��sX[��L�k6��bX�'���ͧ"X�%������Kı<����Kı<�~�m9�7�����ߛ�j���kk��Z향�S���Pv��pI1��k8�������~����]d�&�Y��Kı<����r%�bX�}���r%�bX�g�w6�By"X�'���ͧ"X�%��Ӱ5?5d�D���լ[1313���m9ı,O3߻�ND�,K����ӑ,K��߻�iȖ%�byߏ�[4��BV����7���{����siȖ%�b{�w���K��ș߻��ӑ,K��~��KĦ'����p��W��k�L�����{�ND�,K�~��"X�%�����"X�S�D�_o���S131?q����J�[��f�lKı<����r%�bX�}���r%�bX�g�w6��bX�'���6��bX�'� k��/��VY�j��s>�X�qv����g9���i��N��M.vN.k���٦�j�8B�V�|bf&bf/{��ND�,K����ӑ,K����nǑ,K��߻�iȖ%�b{��^`�B�UKdnլ[1313�߻�ND�,K�뽻ND�,K�~��"X�%����� 6%�b{ڟ_��v��u5%�X�bf&bf.w]��r%�bX�{�xm9�,K��ND�,K����ӑ,K���=�5j���1D[f�l��L��A�=���6��bX�'{���"X�%��{�siȖ%�b{��siȖ%�����椖0��Qڵ�f&bq,O��xm9ı,?)�}�ٴ�%�bX�g�߳iȖ%�by����S131k./˫�?u�\�)*���L�ě�m��!�@��h#`�{:ed+�Wd��Oc���m�!܍��uՄ��VDmU���ۓ��Ucs[c^�h���7,IF�ds���.�V���S�eu�Mp]�k��ԛ�I���[����6���v�獁���v(�1H�ֺ4�+	Y�lp����hC5�״�rj��R��a�n/^qBR�b�,x����A�R��+�,�^WN'T�u�����;���x���p�~��.�~l��$�V����7���'����6��bX�'��{�ND�,K�~��"X�%�����"X�%1?���F���+\��٬[131X�����9�,K�~��"X�%�����"X�%��{�siȭ�f&b}{�P�J�����L��X�{�xm9ı,O~�xm9���� r&D�>���r%�bX�w_�=bى������_O4�v��
�6��bX�'�w�6��bX�'���ͧ"X�%����nӑ,K A�>�}��[1313'��R�BZR�Z6��bX�'���ͧ"X�%� �]��r%�bX�{�xm9ı,O��xm9ı,Jy�'׺֮��F��mt�F3��6q���	�ݍ���q:(]X�=n-��ԗ�u�&���w�{��"X��]��r%�bX�{�xm9ı,O��xlD�,K����ӑ,K��Н�i�0����a��]�"X�%��w�Ӑ�tM E"� ~Ja��pS���bX��y��ӑ,K��;��m9ı,O{���9ı,O~��w335��Z���5��Kı=����Kı<�~�m9�Rı=�]��r%�bX�{�y��Kı;����L�d��u��fh�r%�d"؞{��7��]ӊ(A��p�P�\B|�ٴ�Kı/���ܦ\�0�j�\�m9ı,O���v��bX�'���m9ı,O���6��bX�'��{�ND�,K�߻�HfOƦS���e{�mf���8&Ҽ�����7e:����q��|���XDH��J����L�ı;���m9ı,O���6��bX�'��{�S�,K�����iȖ%������Nڇ%���]bى�����~�fӑ,K��=�siȖ%�b}�}۴�Kı=���i�!bY���=ؼ:Җ2�k�L��X�g��m9ı,O���v��c�
E0S@�RD�=����r%�bX�w���r%�bX�}���h��YsZ�0�5�ND�,K���ݧ"X�%��w�ӑ,K���o�iȖ%��'��{�ND�,K���}�4a����a5�fӑ,K��߻�iȖ%�b��~�fӑ,K��=�siȖ%�b}�����Kı>��췸.�p�X\[�h.��7F˥�:;�Y7 U�r����=�v�;[��U��+a���Kı>����r%�bX�g��m9ı,O��w6�">DȖ%�o�,���$)!I��aK�WUvM��d�5v��bX�'��{�NDP�,K���ͧ"X�%����"X�%����nӑ,Kħ���r�sV\5�.���r%�bX��~�m9ı,O}�xm9�ı>�]��r%�bX���m9ı,K�}���.a�0�3W5�ND�,Q�=����Kı>�]��r%�bX���m9İ:	��`�j'ٯ��ND�,��\�k�͖�;,��r�bى���'�뽻ND�,K<�{��r%�bX��_v�9ı,O}�xm9�f&b������\��UVT��We����c*sx��=t�v�j�d���*b���}���j�`�#�W�[1313'=�\�bX�'��ݻND�,K�~���Ry"X�'~���iȖ%�b}�i~b��G-j%�X�bf&bf.{_v�9�Tș������Kı;��~�ND�,K���ͧ"~��1C1~��k�R�i�Wk�-��K������Kı>�]��r%�bX�g��m9ı,O{��v��LL��_s�Ӟ�I*��+r�bيı@�>�]��r%�bX�g��m9ı,O{��v��bX��d��}吿��$)!}܌+⬚�&���%�]�"X�%��{��ӑ,K�������<�bX�'�w��"X�%����nӑ,K�ҿ�(���܇w�os����^vkt�u�<�GxѬc3�����̤�j83I�8��>�y�a�V�n�\�kn��6�y���ָ���ӆu��e���vW��lt��{u�v�v8lxn@��ó�N�^T�Fl��aگd�nM�v�v�ں鸽����B��Z��uݢ��W��h�jՒ�VۅWS��ͥn���]�t����x�]4�B����(�����yd��5�Z����4�ըGv=�*1u��W�q�Ş`-��U�]��w�L�Z�G
��VE]�X�bf&bb~���]�"X�%��w�ӑ,K���w�iȖ%�by�����Kı/a��Vd���a�.f�k6��bX�'���NEVı,O��{v��bX�'��{�ND�,K���ͧ �b�����u�l���db�U�[13���w�iȖ%�by�����Kı=���r%�bX���xm9�31r{�y�����2Gl�X�bbX��'��{�ND�,K���ݧ"X�%��w�ӑ,K����}��/�)!I
HM�/���*J���kZͧ"X�%��u�nӑ,K��߻�iȖ%�b}�۴�KĳӞ��-��������5<�V�F� �V隁�ѵy:4n���c�[@�����j�::wg+��̫H�MZ�j�4ȫ���N%�b{����Kı>�]��r%�bX�g��l?(Eșı>����ND�,K߻���ff�a5���sFӑ,K���w�i�iT_���&�ı=ϻ��r%�bX�w_v�9ı,O}��6����bX���h�%�t-��X�bf&bf/���m9ı,Os�w6��c�dL�����iȖ%�bw�~�v��bS15���F��NWc�W,�-�������ͧ"X�%��w�ӑ,K���w�iȖ%��'��{�ND�,K��t\�0Ѭ3E���fӑ,K��߻�iȖ%�a�#߷���yı,Os�߳iȖ%�b{�}۴�Kı>��r幙�tɬ�e��d���a�T�4�q�n�]��kuv����M�]}��Ӧ�l���db�U�[1313}�{v��bX�'��{�ND�,K���ݧ"X�%��w�ӑ,K��{�y�*n�UnGl�X�bf&bf/3��6��X�%��u�nӑ,K��߻�iȖ%�b}�۴�Kı\���Gi-Z�l�-��������ݻND�,K�~��"X�W��
��Ө�z��A'�9�~��9ı,O����ND�,K���V��,"dU���f&bf&a�w�ӑ,K���w�iȖ%�by�����K��3"}�}�v��bX�b�|֜��Ub-�V�Zų11,O��{v��bX�'��{�ND�,K���ͧ"X�%��w�ӑ,K=��~�~��~�%.$���J��$��է���ɣ/#� �+1�`�:��Ũ�5&k0�5v��bX�'��{�ND�,K����ӑ,K��߻�iȖ%�by��۴�Kı)���ܦ\՗5MfCWZͧ"X�%��}�si�%�bX���xm9ı,O>�{v��bX�'��{�ND�eL�b^����Y�H����+�k�L��L����ֱlKı<�]��r%��F!�2'���ٴ�Kı>���m9ı,O0e�[��U�[13&b��w�iȖ%�by�����Kı=Ͼ�m9İ*:���G��b���]��"X�%�{��l��-�tj��f�WiȖ%�by�����Kİ������ͧ�,K������Kı<�w{v��bX�'{��>߫	4��-�7a�׵b�a�l����+�Z=���o<�d٢-9+<�������r%�bX����v��bX�'���ND�,K��w�j"X�%��{��ӑ,K����o�֌.��afZ�m9ı,O}��6���%�by����9ı,O3��6��bX�'���ͧ"~ ��,O��7s�IS�l��U�[1313?~5��.D�,K���ͧ"X�%�����iȖ%�b{����Kı=��7�-�ЖHJk�L��L���4��bX�'�k�ݧ"X�%��w�ӑ,K����r%�bX��}{��r��ՐU�5�f&bf&b�o}v��bX�'���ND�,K��o�iȖ%�by�����Kı<\��06
y =\h�tC�k
9 |!E,dM h�\��+�[�
��1m������BJx�� {��J6"]4O`��	l+aH��Aa��M��p!!fdS�f��9�
�0�Bj���b�z�6���%
�	uٸ�ّ�A�enݮTI`����J�lU�OkЯ�!S�Z����[8۶]�g�;F�2�t�  �:u��tYۥ&�ˡ�!�O;Ju�󚓳!�=��[NP@ȣ��嚮NִN@�G�U@Q��KhI�H��SID�TδvL9q3�*�5ʸ���+��]�rat��3�.Θ�nR�ܮµ�J:D�H57f;]���^�j%�mv��;�$�͍D�p$*ݮ�NV,]U�  ]w���n���2�;>��'mpusAc�b�N�P���H��^�>0$�ۘ,��/���qg)������ҫ��	j�n6�ht塺kף"x�:�l�\���*wg:�˳�5�Q��V�8#m�v�n�cRv�����A�B���2�Y"�0vw3���}Q흴<vӹ��Bk�:��Ix�:��A��L�(G��4��Q+�m���3���I��v,ʪ�l��q��86Bђ����f�Gk���w��"��aq�\7�p�fݘ�G�v �R��.�c97v���l��M���j��2�'��ѻمS�J�C�
�-�ݵ΍u�S���[��;�ӝl����؏/R��3m��1���u� �=Y���;Y�����9ؘٞށ�-�f�;J��S��v莝��T��4��T0���ܠ�]�]N���3у�\C ���Gg���A]��*��&�	Iz�+l�\Ӵ�q�8]�X2@����ʵKj�v9�9�[�2����'m��%��xKw>ҡ��9CvX�� �Y��d�ԍd\8������2l ���J�*�h���U�eU�i���kl�Zݑ�F��ƶC�q��Q==�^z�k��/dhm&2��t�7���E�͋g>�e�n��PJ̾V�]�F���EU6�a^��;�sk�s�]u��99a��ɇ�n�I�εv��&��i��^v �}����$>� >�M�#����C�H"���h� 
�=��w���U�zvg� 
�J�]jt�48�5;�V��DB�^�4N��$�N�T�5�gC��܏gF} �r6�uCX�ںX.�V������Z�`�k;���kv^�n|��`�7g<)�5�q�zԗO�[L�%�=n�k��Qv�[]vX�� M�b��Ѷۮ�.��;'gBVF�zz��Q�K�,�Z��	A8�$���,�,F,�$��}��	
��Λ\�t{	q��{H����{b���S�zw��w�ﭭ���E���f�Ȗ%�b{����Kı<�f�6��bX�'��{�Ȅ|��,K��fӑ,K��;�?fY���)2��h�r%�bX�w�}�ND�,K���ͧ"X�%��}�siȖ%�b{����Oȃ��,O����*eV9)Mbى�����>��6��bX�'���ͧ"X�%��w�ӑ,K��g���r%�bX�r��#�r��E�k�L��L����ݧ"X�%��w�ӑ,K��g���r%�bX�g��m9ı,Ox��Z�t���Wk�-���������ND�,K��o�iȖ%�by�����Kı>���r%�bY��������G\�)��
�Q�b�9�by�t��'N�Z��b���h'a�_|;���[�WYsR捧"X�%��Ϸٴ�Kı<�{��r%�bX�w_v�?
*3șı>���m9ı,O�t����mn���SX�bf&bf/�=��<�� �@n%�b}�Μ���$)!H��~_������cN!7dR=��{�柿�/ߋ?�~���u�0o&7�dqh�]�ӥ4���?+�_�@����H� &�0k$s4N��>W��:��@�u��-x�,\%\�# �AN�6�@��z�anwS�a��4v�hn�ur�,��J��[-����;4��8�^/���A��_�ϭ}E��3J�	�E]����|�(����Xq��@m��������Q:XLqYl�_b�6مD$Х�E�H��ۯ@��Z��D��ۘ�i���9Op�g�V����D�����qd�	"Pcln-��z�'�� �� ٶ���0�\��ˉ�K�q�AGisV��kt�K��i��.��}��f���3�2�K?m���W�w���-U�z����:��7��qH�����#����@������g:��Ͻ���NWq��Z����2��N �� �ڂ��0��H��9���s@���$��~ٹ=)E8����FBD F!"x@�l4�h��)�+�`:Hf+� ׂ>讖fcŋ�O�=�ƀ��j�+�n+@r�f���Z{��iҚ׮���?�߅n���\E,苐Mri�;st�G����ػ-vcu�84 &/��6��\�����G"����iҚ׮���Z��D��ۘ�i�9��JgД}����ŀw��N�׋ ��*�$�@�����s@��Z~�Ēo�ﴴ��|hg����jjT�Z��s�o���{l��P����ր;ֽ�ʉRR�B��=��(\����>ŀ7Z� ��ѝY�t�&FH�E�4(�"n�he�*�Q�
��Kin�ӳ�۲�#�y�#���Ʊ�m����#s��E� ��t��:ҐM&ͅ�['4�+�T�4�i���s�UrN��[H��U�^�C�b�h�fܮ[v��m��˭��
�ۋM�p!lf�4ՌJ�MR�3���@��;f���slS��=����ďbܻ`��8�������wxI,��1b��ٷ����Kb!lWK�7n�Ys2Oh��R����zis�qsC�ە8Y�[*�^��7�wK@w��~Q�(I/Ps�`ϐ|�]�­B/��4�n�U��{��r���~Y�����J�$��nUe�@~���=�x��D�Mڰ?y�X�
[T�j19bğ�s�Z���4����*�^���ȝx�s"Q8'����$��ߗ�:y�`��0�r }�T)(����p�F�H{&c��uz�mN�"�9��� Ӯ9lYbٜ�SV`��,��X���J#�.wƀx���i8� ��	��*�^�)�)�E�E�Gh�*Q�s�y7l�?y�3�D|��?~_��cpȚ�G�[����M�YM���sVŊO��J����G�*�}߾0_� ����-���Ԩ�*��%�����B]\���� ��f ~<#_H�n,�]�Z��8'�ڜnНb���u[9Г��ݝ���X+e�7Ko��s�{��`=�r��޾0�S���Dհi�e�@}�;��ؖ6y{��{�OƁk��bG�����8V�v����v���1g�#QH	"1�Xx6@��hWj�`��������I���f�}�M:(IɍLop��b�~�Ɓ�󿖁�kŁ�Jys�0�%��L��5jl�Dݘ����_~_�����?=�hϑ�6_����ɬ����i>$ӱ��9\sqO���� m���.�vY��s(���f��;|h�����/Oٶ�����~���Ġ�����M�ҚW��;�w7�G~u��X�2?�$4w���*�^��u��.^��=�ՉH�Q���h~���Հn�ŀ4�ـ�yTD��(���DTM�_o���{��}Mh�.n�SJn�{^,�
%��}߾<_��W��;+G	*���!6��k�t��Y;it��&6�:�ɚLsj���F��z3q�M�p�F�Rf�r�������U��|�����?[�G�P�#&51�i�@��S@��Z��s@�zSؐg���N19�Hh�;�h�]���M�YM ��"aLnD�h�u�Ɓ�?Y��>��������{�>�~�l�*�7HڶU�{l�;��������׋ �X��'#��Е	���h�ZV4��.��eq�̋��y��0!��m���gqh��d�noD�Y��Zy�q3�5�V�`6��&�ӳm�p������r�3�;Uͭ��^;=�ƹ����>M0݈��q�0�lZ��p6��%�8�m�����M�\Ʒm�H!�g;�u�r��`�dY�5���AM.�'hI�䷒��cac��V[�l����{�����(�$��nI���MY�3\�kE=�#Z�r��m)<V9�Cy.��n`f�M1c�@s!#�nE�:�M����]�ٟ ����h��bR�!nd�� r��|�M�ذ]O� ��lϖ$_�c��cDQ��$zu���\���>���*�^����;2&�8D�q)3@�_U�}�)�Uz�ى��ր�z�g�Kkj��G)�7�)�Uz��빠\���\0E�#��G�����f7��ͥؽ"2���z݌������~���>�g�����<����XN���� ����IE\u�4>�t�Չb�BB0dd eTM�������W~�{����9�L�ڞ�%[�X��m[*�^��7�oM�o��-����=�[.,�d$�K0�v���8���>P�|�������H49F�F�Z��興�}�~�;� ��l�=椷V���JUA�Y�����k�h���F�%m�ɗ��K�G^xc��z��=�ޮM��?�n�ŀ4�ـ~�|�~��Ӏ{i�?�nc�J7�4��7�����ŀwS��=�x���tɲ��U�uH���������^��U$�BƐ�!P�TH`>0$	! <G������.�(0�!3�4 j Ԩ� 7&q����K�7�>=~�6@��12B�d~"�#�2�؋F-��ҥa�@���Gc���Ɛ`@�A"b�����@��a,,$�� �V2Э+)		,M�G_(n͑�a20����! 6�T�D�!FR!B�+b� D�E�#\!v*�B�>�:�)�D� ��`@!	��J�)0��5P}"'��Qx�A��H1(� �8�'���4�!�
����Q�4�A��>ٹ'���4�q��僲��C�h?f,��}�wӀ7�b�{l�?y�X�Մ���"h�-��M���w���߷4_U�wgD�V#�#�-L��h�IR�`�,c��de�d���۾��	4�%�V�UJI#Vڶ��|h�n�k�{���:�qBbDɐ����0�o&N�}8��XN����Xԍ4�ڙ��Uz��׋ iֹ�?y�X�)7j��u4�v٠>����]�������b�8)d>T@�B0�!�4��t�L��_f���j��4���n%&h+��n�k�h�]�����7�Q�Q��D��jʥ�غ�svۋ�ޭ�͘k�z9뫆�@c�X�Adb��6��w�ۚ���=��� ��]Zi8�O�j� �k��׋ iֹ�?y�Y�2ſ�L��B&�"�;����}V�����-}V��5lI�	2je]ݬ���[��=�ذ�\�rIc�;����y
�2��rc�������s�{���:�8I,�|�=� �X��dhP����>�0�Z�2]h��j�&g��{G��(;j��Cm�8�'���鰵�V�];q��,�6�[Hc�8g�&nњm,&���k��C�m7$c����[ezN�X���-i3ud�4TM�4qȼ0�5�v��H۰�6��]��I�f�z�C�uhPm��+�[�٭"��zh앳���JWog�X�m�0���N��:�P�H�ȋ�܌��w��x��ǻ��	��Z{s�P#���	',6e�tt�pQ�]���{:���cR4Ӑjdrf�yڴyڴ�k��Q�Cw� ����R�*�^(��@���@�_U�{��h^�@��udnAB%�I������ŇB�Jg��V���tɱ�(4�'����n�U��{��r��@>3�V�N1Lq��Nf�U��{�4��Z޷s@�{�T+�E���)�ۮk��m�taר�JvX�����71�g�ݖ܉�����Z� ���tG��0:��"�*�X8ڶS@qrw�I���3�
!�h�,���q�wwZZ���>�����{b�B��24��r-�[��z�V��t��˓�z�{�9h9VZ�Ř�z�� �w��i��?y�X���J�t����נ>�����.��y�w�ۚVנwvS��6�d1�a�q�.��[���dԝ���ĸ�4�li6��D���' ��Ĝ4�ڴ���*�����}�d���Jbxۋ@��M�k�;�S@��^�|��q�4@X����ڴݶajD		B�IKu-��� ��ꁃp#�dqh�)�WR�`��`r���8�uu����]��S*��`ԷXD(�������h�w4��-#j9$IH�c��5�\@F�%�n�m�5��V�3�Q�Z�V�g��I�iL�7������Wj�;��h�k�=H�N@M���h]�@�빠Zկ@��M����K�*�)��թ����}� n����
g��� 绫 ��*�ʻ���v(�JL�-jנ}l�����;3<�$v�@��T!�
i_#�ۚ�P#�,�A1�16ӏ@����I�wW�}� n���>Q�Fu����D��& �jD�>j��ۧ�n�]��fO<мkaݶ�Ì.�p������wm�u-��/��0;�@np�n'����қ��v�e�Y�/��".�꟨SB�53%S`}�_}8�,N���>�@��aq2b�Qƣ�9�����n���8�{�{� �w�e��F�&�r����4Gmܓ�}��䘎� A` �"F.����:��m�D6ݔB���>�d-�� �@�\����5�t3��[T\�;x��f��I�����6�,j%K��-F�����V+]��6��r��ǅ�+����������6:���FM�)1�b:t�;.�2[=A��xN��i,a�(1��lS�P��vf�2r��(�l ��i%��5�:ڮ-�)��6Ļ�����8�;������\�Y[�\3�AVQ�i����k���;7E�v�¡�o!��	�����w�y�1-�
�>�~��֭z��h]�@��ՒI�#xȔ��kV��m��n�ݶg�EQ��Y��WWd�Ҙ�iǠw��?Ɓ�����-o�� �����NP"%���bX����� �����n���0=�� 90�$I��zwJh�k�>�S@�mzעK*��R�N9�З95�VU�g�=�wE���7�"�vN��ޚ5�Q�r�Ycm�e6��4��M���wY�|�0��1F�#R'�@o��5�X�ř�,��d�_�����h�k�>�H<n@J)�Uf�۬ ��x}	)�⻧ �u�uK�&8�ۘ6G���+o�~�?ߖ����+k�;�dN�rHһ��&���np�߾���:~���s���bI%�ވ~����Z�m�Gj6n4k��0���n�h�tq�J����i�1I��m�����=���h�W��f�h�� ��u���L��Uـl�u�%27O� �}X��N:����D��Ǡw>�I>�/�f��>���Z!�f�(�
��S~̿��ﺰx��tU2�mWk�~ı'��z�z����@�}V�����0��G�U����`�˾Ͼ��]��Ժ��x�N���j!�Hy"NL�Ŷ�ԇm8�nNZ�6�F�E҅q�:<��V��+p�Sp�9[^�����v��� �u�w.:.��7Uh�.����9�Q
d���8�����Y�ɭ����"Y$m�G��?;�h[)���/����@���@��&6�7�)�����?7l��� ݭs�p�DRP[xP�k�u�]�'����r���1�!�Umzs��ڴ���/�#m�cy��q��q4��Қ�����3���%Y�81[v[d�.�l���8��q���Z��Z׷��~�������յ��:��v-�v��e4
��@�}V�����0��G���@��M�k���Q2�>��Wt��m�svR��
��SUf(Jz������:np9D��8�;��wEک&�E���Z� i�s�~nـ9z� ��2Da��x���Xč�X�A� F$�1H���� �! �M*q���B,�������`B�B�F�*! eXEH�$D�}�$c1�!P%�����!D�D�h��xCA��l���#0�='�z��+���F#$�9(Č>7�"��2꣛.ѣ�
2a�B�T6.z�a�+>$xz/1!�4�S�/�8�5����J������	�H��H�qD$H!:�Ie�K���c���Ը�����+I�4��/A[ ���O,�t9�6��l�pi��L��U�6��.�nv2���X��9�l �˘%EF6ջ�,`Rj P�b�^��a�*�5f��[M���0���$�\6���&R�t�p�VҜ�8���u;n�j獸���GL;��x����VH'Rk���*�%W�I���rq�.�aܡ�G%�sq²���Wh��M�iv�Ͳ��P�iV�W:�ջS�њ�ֱE�9�-�6]vHL�A����#mrQ�Fی��gM�V2�f�9zU�K�˜@s�en��Tv�.ԧ�5�H�Xuiv���g��q���G7\Aū��S	V�+<�J���2�9�+���zW �Z�9�d NvQ�c3q��i�Y�m�U�9\m>�ʹ��P�u9�]�d��HD�M4��$p�͛-�YAr�#�*�ĳ���U���s(	gvL����[�1ӂ��v�n�fz�lˎ$��v��8���k�nƵ��	уm��y]�pH;��vk��Z6ٺ�x�ZvL�K�Q�����9`v�-��U�#��6��Ż�%�Oi�ũ�'��=sBd��i��K����3�J0�@�����_konMg�4bޙGHmq�vѳ�;Dg��o�,m��W*�`��i�G&��ɤ#�ëF��nR�1��x1	��X �̣� #y�p)-]+l�L�U ��,C���K,�4�ʻs���0�-��F��W 5+9���]�Wk[j���P+�tr@�띸��6Nr;�Z�."1D�Ŝ�dV��s�,ٴ�3�UH	,�5���U@ JZ�*f����u��[�l�b�)�1a�NHeǪ��n7����XXx�{[vl�sm�]�vzz�C�u�,y�{g��'N#��N�M��dr�9�2*�؎CV�܇V0Jk���ۚNm�q�99&u�<�ѷZX��浗�kZ�3S&������>G�����a�;��Q��� �)�	�<6
8/����D"&|'��u̺�5gY���r����&�H�J��E��qű�6�D|幰��S���t�'v�+z0�p�e����F�vŶ�����]g�#=��U<�&�;������v��ּ;�9����`R�D��ۉ׈y�����\������Tƴ��cv�	�[��4:t��1t>���M	ك��'����]m�Fŵ�5�Bܒ�kګ�.�yf�U#���'�+��Ki�e�ӥOB���N]שz��\v��r2�uJ��m�^�� �ݳ r��DD~�n�N�����Ɯ��jcxۋ@��M���Ϫ�.W�h�guJ$�d�,��U����h+����8�y2<q�#����ح���?g�-�e4
�W�{<�i1Z.fe]]� ӭs�t(^��?�ϫ ݭs�t(�嫲T�5=E+�WH���h��O6�
n�+��N��/�wAҫ��6D&LQ���Ⱦ߿OƁU����=	%�C�S��<���5e)�������}�f���ҫ1�E;'v���Z��h�-���`�$zs���Z��h^�@�q�c���F�qh+����*����Zף��1�1��T��� �ݳ �]�_�n�N �v� ��-i2q<CDƈ���ʣ��gmsD��7O[���K�Q��v��c�%�brVנw>�@�_U�>A�ߧ�@)��`�LoCq8���h+����*�^����T������v���oMX<C�^"�_��ܓ�3���=ìjTZY(�A%4X�I��kƀ���@�}V�|YM�}a�����ۆ�˺���Z�e4���>�u��AD9bQ�c���q��5؝;������1�.�ru�+��raG0L�=��Z��h[)�r�^���;��2(��/S:$�Ow_��X�k��e\�6�7�)��Hh[)�r�^�����@�O��a��(��Q��,N��6u��7k\�Gl�m(PG�b�,Yy�zh�v�D��2Uv=��Z��h[)�r�^��c�7~6үl��G�X�cb��j��m��t����������s��v�[�5�`��_����@��M�Z���h��P��$#pQ�7�e4Z�`��p��g�DL�t�˚��Ԁ�Sp�*��=��Z~�K�?OƁ�ߧ�@�3����(�
G�w>s�=� �ݳ�D)t�� ����A�9dQŠ^,�����.����h�g֪�"���N���v��5�s�qF��.�T�4-�;�[/B]>��6ӬR	��+F�K��\>d,�뗒�B
{JV�f܁S�e��n"8wY��Ơ�[g����8uuݡD��ѪLi*�*P8[�>޷5�����.=���R�������#�m����q'�Ϙ��m���6�K%�n֠s�7�0d�nv[����V=N�$�[��KC,%a����9���X�n6�R�	�v�=�=sp�{q�uб���ncXҘ�$����?.����hŔ����I�(�br.����hŔ�>�S����N�ER�Uj�殰���Ŕ�>�S@��^���NdI���Z�e4���9wW�w>�@>����a ����hWl�7k\���p��0��"O��6�un��58#C�]B���qAV�pd��N�^�����JU��-lIp��
�����hŔ�>�S@�#;����Q)e������$���R � `#@C@��=��x�;�)�r�@�p���v�
�@w㷦��{zh�,l���h��hw'�drcJbp���h�Y�w>�@��)�a��(��NA�X���z��s������h�5�I$�Fۑ(˝1:6�vآ콡͹��:��q*>��̼a�;��I`�LL�Nɠw>�@��)�}l��{����kHs &�1��8hx����h�Y�wt��w�
#"�<�}l��<�ߵ��B� �"�`�)O��,bɘ�'���@o�oM�Nv���N@M���h�Y�wt���S@��M��q�Ȃ70xۓ@��M�,�������h{:���F#����@�n��	���'ɪF����[��f�6�9�(��ni�V������h�Y�wt���wN���kS���>�S}����)�}�� n=�D�bs#��9 ���;�S@��)�}l��{�-�1����#�@��M�,���{zh3�ˋ3�vww@o���5n\N1�,��@��)�}l��z��wJh�u#"H�$`���ư�㮍�&mƫ�L�#ͭ� XqV��λF�F:L�jdx�@��M ���wJhx�������M96�n��h�)�}Ŕ�>�S@�]�u�����NM��4{,������[4���jc�#O����e��>�S@=�f��Қ�9:�71�"b�$������[4s�������@}�fw�f��Ȫ����<�����v��A�+��X4f�v�N��5��l�;V�\��k�u9m��^ڹ�������Ղ�ܢY�%��ֳ�	ѤW)����b��re���ը�=a��;�x9���m֛\�7m�ON�9<�Ό�+������ԋ��9zLsOS���hުc5˙u덞�T�m�-��½ɽ[qu�))j,�33x��Ѣ&5K-e��.����
��תss��uo17���=�8�p�5���G��r����7vـ{��>I~��u����-�bqA8'&��Қ��S@��M ����س1bl�9�1�h�,!V8h��~4���z٠wt��{܊��a0s �n��h�l�;�S@���hs�#�4�ډ�h�l�?[w����~4���;9����'�ǒ ��cq�=OQ���8^��E�]v���ǜiL;��v��rm-�Ɯ�s��YM�e4׬�;�>�	���<"�-�,���X��P��T6�	'�jx��@�}V����H�#����Ʋcy	!�{����z٠w>�@��oM��:v�[�Ud��M�b����|`�;f��f ~<6�`�LN('��;�S@�Ŕ�?7l�y��:!$���$�Ue�)�9�]'.���nW��:�S��]�s���$f8�b�!��m����=����>�S@=�f��Қ�r*I�Ȣ���h[)�yzנwt����)�}Ϭ�$7 �m�@=�n��9zhjbW3����+�tI�B�߭OxD�"!���c!�I ��A�A�� �"2E���&���K� ��K��Y!#�h�JF�@�"BB@�d�@�. �$�V0�_ k�@�	hF�*BË�c��<�����C[v�@�"iD��� ��|�@>|��pdv*�G�>U֐�(x��D�Kc�~�� �m� �:��*ǋ#srh�)�}��h[)���@� ������0���>�e4���z٠wt��k�W�n͙��ٺ6�j�k���V=��8�&����X9ga�ѣf�-ӓ�^�[�>�S@���@��M�S@��RƢN19����h^����ċl�h���h[)����ǃy18���@��M�YM�e4�٠{�[�C0Q�d���V���k�$����Ҋu #�'C|#M��v�\��Ny����h��QBG�n-�e4����|�~4u���Y�9<�nH�c������9��O��7�]������tv��N�/�;��frF�4��@��M�c�@��M �b��<�0��Ɔ�wJgBJd��]8��� ���B�P���,�H�9a!�u��}lf���G�׀6�wd-��We�R�U+����ϻ���u��l�=�:�
��[�8��F��@9�x��0k�s��w�
� CW0�)|��O�3Z�)uK@j9(53��
���K�6q�G�u�E��]g�[2
�7 :� ��������i��5�\[<�S-(��L���y8.��2�2�KŹ!��k�֠�l��-s�Qǵؽ�N�ե�&C��'v���[>՟��ﳺ��E{y^�-YF�nQ�5�T{8�9g��z,�r�jk����۱xV`�i��V��%ř���G�Z�z�kOo�˙�'v�G��s;�G�᦬� b��m���/��@x7��	��<u���e�@>����*�=�߿!d�0S�H�{��h�٠z���4�T&LY$JD�	ȴ�l��f�����Ɓ�����t�!#C��&�uWx�/�^ ۾0k�k@>�� ����d�D�4G$�;vـ}�:�����^��?2�����ptpT�1���V��[�Ѷ�mѨ�e�\��v�ӶX�y�v�ݘ�۹�ͻ�z��	~�n�Ɓց?E!�Lo$�- ��ypBJ&+�
ДU�[��7]�{��h{�%q�H�PrM ��ݶa�)�}}s����7Ah�V��������B�D*�����- ��4�Y�y�$I�0q�d��݆�}m�׬�;�S@m}�DHu
�ڪ)S���6�U65؜�;id�N��-uQ>���v��{�/�:㜂q8�7!��~�4�Y�wt���a�{�+H�N@$27&�s�y�26�_vY��w�芠�OE+VM�+U%�������s���'�!�`T�k��$;���|�9֫��[d�Gi��c���f {�� 5�wm��Er��#ɍ�C@>�� ��h�l�=��(��B�;��Yr]���Nx#i���jõ�8���;�[m�g;��1a�D�N1IjI��M��4u� ��4���7��VU���l΄�ɯ��p��x׬�ؑ˿?�� ��	���@��~�@>�� ��h�)�w5�	�5*�WlN[^��{޺ ��9��nMa�
i�"=#@��1f�����{���8�8'e�׬�/t���Š��װߟO0�su���Ա$n�h�Z�{�,�ڢ�v�㓮v��W��ƞ�9&�{�4u�- ��h^�@�Ƴ�ț��Pl �4u�- ��h^�@�Қ��+#�m,�4������ 5�9BIL�w���톁W��bQ'�8��h]w�=�f�o,���w^ �w*�"����%�@s��4����^�`�׀���
(��BV
Dw��dDN����9�=�lՋp;1�5nz���M(;gs��iɬT��mϝӉu���m6ܗB�U��rPhz�+���@E<�Y��X۱m�63Vņ�m�֫\��cf
���	��-=\����c�یb����uv�K�|�R�����\���UAx*B��;���r�IIpe�,�bwg'l������+�Ʃ|@t�$Kv9MI.��#�sd���x����y��9��pW8&�R�Eb�j�:Xy��fѧ3�Ӱ=d�?�>�����!��Z��U�Y�����0���z���H~�~4Z���1c���r ���BS �����{[�0nې�"M9&�G&�u�4�)�{��h��@;�ο�&1%�drM�Jh�v}l��f�}�gW�9"�a!�{��h��@;����;�V�9�y'�%*:��mƝnzg�Z�ZX��k�(o`N��V3��B6"by#���f�w[4�)�}�,Z^�-�D�b���۠s����Ė�I*�I*vv���s���r�S#�)�R�U+WVdNɠ~�~4���_[4��@����&@o&1��8h�+Z ������'��0�/��-J�q�q��� ��h[f�{�4}����,����WXF��`���������;r�GWV�4 �\��۞����8��m�5��> ��~�wJh��m���P|5��U@vJ���4� �t��f�u�h�k��Qța�}�X��~�������d��E�d,!��˘�Zgu���ܽ4�૝�r�lD��I"���@;��wJh~������aK����Y2F��@7[��"!��~���8��x������R�H��e�)� ��f�y{A��A�s�йw��-������\�t�Ârh�)�}�,Z��hu�@��97���@��X��n�u��7vٜ�Q
dݩ}%R��"<�h�~�4�٠wt���YZ�=$i� 4�(���� {���v�p:!Y���,X�O^�t�{�P������h��� ��hu�@��i��$���L��kP�1���&7b�]�I[/^��n�WI%/B鴈������ ~n�[w�G�t�pZdO�bs#Ɣ��$�@>��������-w��>�,Z�uh��,���@:�4��hu�- ��4AŹ2cp#��rhϪ�>��- ��4��@���$I����E"�>�v��h[f�=�=��I�_�����
����@�<�4��m &	 704`�	pQx�S@qn�4:�P�.h܉dr!�#9�mL�@�'b��(R�7"F$�"�a	 #	�0��$ B�'�9��"��|M�a�myȠI�rC�!*���$O%mx�F1Xd	 a��*C/��� �!	u����N"�<�E�9�H<~}$;(F2��3�e"�,"��B0�f�R�y�Ӆ��b9y�����9��'GŊ�n�1�kp�t�c���l��۬� i�����Ӧt��͍���>˥�ݛX����e��jWm�� �HaBP9A,p�؁)&8����A�PR��洫+͵��m4�gZc�2mu!���P"PP��j#�Իr��D��ض��%�"��ݺ$�8�A���6��
�l8��	2�m� Ԑ<�n��Iʻ\��wm��f�t�W]����۪�ivZYWq�5 ʵJ��pF�\aѷ��.��I˦y�<�9���EZ&3p�шĂ�Z�����va�P.1��D�P:����Br�����3\�1ZK��������	���k!Р�̝nC�Þ���X�J��`NX�6@zӄ���9EK��mrt�����Wdv��ŵs�:�%G[p�G+W<E�ss�&st�-��]��Y�R�㨥M1kb셪SmL8��UZ�X���(�j��)��N�n�L獺�̠�Ͳ=kug����]�-��]nc���kv�m��\���ش��L�,�6j΄M�z�I.œh,/L^:�8�@:��WaۨA�����`"�: j��zXe�'�A4�v\�1o5�[��6(�0��YN4��0�U��b���5��EtqY8����ʍ�9;��ў�+s˘/&�qn�ƘC6�enT
����u�S��hn��Q���n{4��� ���D(&U�R@h
/$A�"8� øض�zr�Se�j���8�j0*����Glpr��6Ů��:��9o4�ٸ�hκI�Ԛ\8�66W�ؾ����F�(8j�%�H멞��V���r���3[��V�ؒ�ztT�f�xd����o��ڹk��#/V.�����)�ϻٮ�,;� v���s��E9m����:�������t���1�j�u �2��%�w�,1�^�eݮ&�Z�=�n����9���{����{��(�F'��S�����]���UT�/!���"l���k��2�Lѩ��W<t��9���qAf��c�y^-�/M.2VҜ��{Y�xM:��_�d�1[�耘��r,ή�Z���)�q��[Aa5߻���˴y����X�wh�"[�����e<�m6Z�����/!�1�\��C\���
+έը8�5o7;�U���z��i��	����8ۮe�}<��\������.��n�\�uq}]�[�S5f�k1{i������V	^�y�wK)C�F6N����\sR!���5<�����@:�4��hu���Xc�&���Y�@:�4��hu�- ��y�	L��S�
n���� u��@�YZ���@:�4����d�#M�#�@���h��@:�4Ϫ�>�2'[��LN)#X ������������S�{�������	أM�&�P�D��.��8G\���-܏b
����l�c2hks#�I4�٠^}V��YZ��f��V��������o�����Ua$FE�H��>eO�h�~��l�������$�@i��H�w��- ��4�٠w>�@��ꅎa1�q��@?6� 7[�v��B�>�ι�<��4Ӑk#rh[f��ֽ�Š�f��8�v	<AL~�.��p�j{l[�g8��C�lM��=ڸ�wi�Y'��Q�6��9zנ}��4�]�H�� z�O�]�R�ꪐ]��`���9$�"&Cy�����w�^X�&��W= �V��-�� 7�^ kn��GO�2�D,Q	f����߿l4�x���,���9&�u�h�k�;��4׬�9����ܚ/Z��{����M �l�>�L1+	�4T��1t���\ue���u�#j����3��Lm�"�$���
1��@�[���f�u�hzנw��c�I�ヌ�h�@;��^��������!#M9�&�G&�w[4
�k�=�+Z{��>]�������Z���QսՀn��N>�ߵ�=DBAFEQ�)��D��,K�oz���u�b�9����@��X��Y����Z����x�w\ܥn�rk@V�v�v�ظ�c��7��@� N/,���:9p�9:�I�^�4�٠U�^����h�_s���[V�Ic����n���ӽՀ{z�� <���6��U�A8'&��ֽ�Yb��fbG~���[���<�]c�2��bX7����h�Y�����z��\KȦE�<�h�Y������h����3339ө&�նAf��>��z6�[��kd۷iT%F���H��2��Gcj��;!��k�<\�ba�X�]�6|,��v���ulΰۉ�P�
-�ۂ�HE�Ĳ��e���nQ��82:R�b�s͛�ע�.�v�ⶒ�7�[ӉQ�,�{e	�۰��Q(=���0�p����N�B�
a-�6�Rw\����y��&��_����www=wە�`Y�
jg��6�6=9�#[y�ΐ�mH�i�;7\a#Q9
9���7&�[���9zנ}�,Z��h�/�'V�U5w�l��ϡB�=�}s��^ kn�BJd�B�Ҭ�QWuT��� ��~k@/u��٠U�^���vA��&'�� ��h[f����D%���pP���sws*��j5$����Z����^�4�`��E&�ũ57�M��i�^���6�,��uz;tW��T�!�M���pnO�����}�X��Y�m����y'���K��>�,��IBN=	D�Vۼ �7x�7X��\I�$�pq��@/u�ջ��J&zw��>���ݚv\�ɑ(�G&�u�hzנ}�X��Y�}�8��70xӓ@�ֽ�/og\� ���u��?mJ4��_����71����r��Y�x�,�D��H���sۉ��OnX�\��{ji�c�Yb��f�w[?|���ߞ��TI��ndŌ��$�h�@;��^��z��{�T���d�6�Ww��� ���BȈ����By�1\X����z ����aýV�L�� ��@�ֽ�Yb��f�D(�o�����
Ue��7EJ*���e�@/u��٠U�^���!�v�N�����m헛��	����Am�G�u�G���H�a�7V������ {��[w�9�u�(Q�Cϯ�Z�_���70j,Qɠ����!L�;�X���p��?ml̎.a Q�Xۓ@�ֽ�Yb��f�w[4�1�Y&'��m�H�z�D(���u� s}x���5DBV�4b�h�C�x�����nI�~��>��1c&&I$Z{���f�W�z޲Š�$[�q�y	:n��GJg��v��s��)�:d_C��4CkӦ)"�##���hu�@�ֽ�Yb��f����7�q`𚵀9�u�~�s�u���,��H��_� "(��n=��~�@/u�u��^����ncnb�	H�׬�;���9zס��,s��z �;=B�5d���d�@n�� �[�_����� y��Q
.ffqqA��Vȫ����n:#r��kgce��HV�gm�+<V�q�:�4����lwGG<�s7v�B�74�Q����guk`��덻5�������Uum�
G<T�\�2�=�Һ86����';<Q����r"�k�8`y��3� y�R��p��m��jR+Y�ukbE�dI[pǶ�W\�Y�-ŻM�JS�A3�{���������o��i�]qp6^�,C�q��7Kd�+���,vŶ�9�7f��=�a���Wh�ۓ<��^����h�Y�w[��w�}VI��8�xd�G�}�,Z��h��h�k�>��sfLL�H�׬�;���9zנ}�,Z�3�R"�##��$��&��,��V���� y� ��J`�LMǃ�9���Z޲Š�f��s@���0�AG24<Qe�sQ�O3İnms;�+�oi�__9�_�C�LR&�PR/��d ���@�t����@���q'0Rc�	�M�'=��n����t�Yg��ͭ�Nu������a��=B�5d�5F��:����{�U�}� �����$_�0�(�$ܙ�{�U�~��� ?kw�СN��� z/�Yl1����G����4�h�w4s���	�Bc�ړ�)#ز�<5��<����^5ݲnoX�^;c�X܌�<Lɉ�9 ����������� �_� ���J%FLq�5$�=��h���>�]��w���݋,s�bd�0Nf�����u�i���pT�BH��`
�n<M� B�l �U��WlDĂHH0��%4�`ETB!@M���L��A��I�H��>~���$��Rh�����d��krA�
t*�
�>0�0�P�H�C@�H1 HH0##�$F	��� HHB, ��%��J�"B+�k�fj	F,ށ���d$u��4���G��~���j��<X|�E��K�  ��B0!��#!D��F�@��=�1M�$X�R$H1�LN*݂�T�dQ�4����(�(|���iUO���;<P�Q6��x
 v��)�|�O��6����S�ޥ�_krN{��4ݍs���U;\r:;^��?��n� ���n�09DD)޷Ӏv���)���BG�r޶h��=_U�{�vu�(���f
@�M�6��mB���gusm���m%���n{sl��X����ME�94wJh���=�yg%�>��<�̩�E7V�nL�=Ϫ�>�]��}���n���H�_�!c����-�l4�l�:۹�z��@���v1��2bd�C@;�������Z���P�^�$R����$�D(F� 4���u�� ���v��S'���S@B��n�]b�XK�@n�� �s�~�yf o���K_~���ڠ��	�
Fh�kngœ�ݢ�v����Ё����Ó�u�<u7e�1�&�~z�N����n�#�}ذz5�VӵT�q���zw����	%2{� o��Z� �ۚjf������4�l�:۹�z��@���h{�����X��C�(��ߖ�O� ����n���,W�L
9��&h���>�� �7x�x�_�(H���:�T�+HD�����lw�-Å�0��N�6�6Ta�غn�'v���l)UnK��֞�!�̀W$�֍��T��1��V�x���yS@sH66.6�n��qp�m�=i�Z��xi1Q����ez�s\K����
��$ʲ�*HnJ\	��ݠ5�Rs\p̿��lf0=����W;[`�<�o[���-U�ʢ�;aeK�_$�fe��r�&b�m�fgP��sRೝg��.����H]lE��㱮�m�����+��qh�߶޶h��h���>�N�72b�LL��hz٠wW� �s�~�yf}	B�!s雙.��ҍI4~��=_U�}�v�[4݋:�`�LLq�h��hz݆�}�������u�b�&)M�)����h�l�;���=Ϫ�*��bE�q���BzԷ=x��<�zΫ�+�9,E;t;�)���e��7$�H�X�#�� ���u����Z޷a��Π�0�F��޵�'�����< �J+�񼙙�.�{��4�h/v$_�0�(�&ܙ�w>�@���4�l�;���;�3��F$i��8��n�@=�f��n���^���"u�9�2bd�C@=�f��n���^����i������wƄ��$�m	�*����v9ιѳ�u�<(4��;�ه�jr�9'���4/Z��n�@=�f�{�u������@���@���4޶hu�@��ıJ�v��u�f�����n��3�!:�R�3F!��(&x�b��}�]��}49��Sr�emHH�nC@=�f�w[4/Z��n�@3ֻ$���G&�w[4P�mk����,��n�M����:�A��3�[qրw'��m֛�-Iq�q{9{M<�mq���o�{��>�� ��� �h��up����3������h޶hu�@��W�{܈�pNdǌ��#���l�����^��[��a�ԢD���mF���٠y{��9��oSr��V*PG�Q	|�Y��Z9�y12D��@��W�~��� ��� 5�x$��␚��p ��d�C���� /,�r&�֍ٳ�qt���m�X3uŉ�?����0��� ���$�Hl���:���JL�ı�G�r���ջ�=>�X�o,΄�$�Awu.�W0&B<Qɠ���@��W�u����� /���Z����A�'k_V ��(��n�[w�?"��0��f4��;��4�[4[w�z}��	I$�!	$BP������]����}9��K)�anր�nF8 UA!�,��ph�Q���l���)�z�t�$��d��s%�2Ubzuٱ�;$���0�띫�*�n�"�M�g+m.ɗ�0�n6: �t�u�f�pi�"�sN�q�s�+�l]��jM�b�^��ByV�'���ꓮ�8�m]}�Y�$�d���=���<�U��n��⶗.��I7(7�߽���>�w�ￊ��5<f�b��;V:5r�͎ú����c=H2����wntdf�tǌ��Q�|׿M �l�<����u��)kQ&�,r�ԓ@:�4/uzz�f�}�f�w,]E0o&&8���<���u� ��� �h�Y`<s&((Ƣ�=�[���l��f���@��Ĝ�k$x7!�z٠����u�~�yf�J#U&.�8������L��n-;d7r�Ļs�1���C��������܎j�EX+P����[n�;�z���� ���Έ�����5�k���S�[�>s�ZĽ��fU�y������BQ�!x����x���/�gW�H��q�z݆�}�f�w[4/uz�ȉ��Lxɍ�C@>��@;������[��aKZ�8ŎdmƤ��l�<���z݆�}�f�z�E����g�l|=L��=Om"Nn�����]�l��u��'9�nۡ��^�s���m˯�}�v����l�=j�`U*���#��4��uM o����l�<��������c���0��� �n�I&��"6%%��"%%�RQ��N�V�7�`m��2L29���I4�٠y{��>�� ��� �����Ěnb�����py�� ?6� 7[��{��Ï��'�Q�WP�Puظ�+�#ŷOZ�G�h�m���]v�vZ{9�u�!#_�&���ߵ���hu�@�}V��r"u�9�8��f�}m��l�<���=�u��R֢N1d��RM �h]��z݆�}�� �9u������C�D�7Հ{{�� ������RI(�,�A�4*�b��k���Ns�]��V���u�f����[� �n�N��(K��с�B��RU-���<��p��2��k�#5E�h�v����k���)y���> ���hu�@��@��X�/W�&,�C$���l��S&�}X���p��x�V�8���c�Q�4.���e�@>�f�w[4���&?�5���z�S��� ��x����n�{f�;`�UE
�V�^�>�{t�f%���l���8���I(�����
��DPW���
� U�(��Q@_��*��ATG��
� �D`�@
�B*�B�*� �D����*P*@B
�Q �E@ �D*
��� ��
�`�B
�`�F
�H**�E�� �A*
�D��`�@**�P *F
�P`�AE��P��@ �@Db�ED��H*����
�X
�"�H*`�E*U�����,*`�F
�`�@ �D
�P���*��X*U`*Q`�DA��
�
�H* �E�� ��EQ`�DT*TD�� `*PH*��"�EH
�
�X* *`�F �H*�"�*���E��* *����D �A �AT��E `�D@��UR
�A
� �D*
�*�
�F
���D*V"�* *�� *
�T��@H*R�`�A�X��`�DR�
�
�b�A�`*
� ��@"*b��
�H
�V"�`�@
� *�"�B�("* 	�@^��*��U�(�A@^�
��E U�(��@_� ���PW�E U|E U�b��L����v8C�� � ���fO� ��|�AAJcJ PQP 
'l��R m� ��h�    �y�
�UR�@B��BD
������BP(� �"�D��%QU)P�*H
� �   � �P      =�K'}�m��'���wm^��(��m�����-{j��{{ǝK� ����o���޼ μ��y<�. }i 6�^�n`eW��EW-z�W��:�����r˖�mT�5h ��@   � yUY�֩�fr�&��= =�U�E_{��%e�m�]U���B��;_my;� q��UY��� ov�wۯ�W�7I�s�ҫ�J, >��mm��e����u�U�j�x�P   @� ��j۾w� &�)f ��P Lt���Y�L@��(��ҔEh�()e�(�  (,Ɣ�14���:\��,�iJ]۔�JK0=t ,�(/v�@
Y�)E,���  ��  �   �!�e(4�,�W��Y^���_mp���K��{������͔���R� MK������������^�<��M� �O[��R��zu�����+���Oz}N-�[��_{�R���| �  �(   �����w}��<��������z�n@���ڕ�۷�O,�zy:z� iY���>��_  k�O����v׼�>�L���^���n��iz�=��x �-���_+͗-{�w������׀  ���IR�  E?�e3U)P  Ǫ�J��14�F=��@J@  OЕ6ҥ)   "(&)Ri�bq���?��/��q�Y�9������s��(*����"���TU?�"���H�
��PUb*
*���gǒ01�)�_~�~!��!Me��n���V��<[�v]���VXӕ�8��� �w��#��R���u�A4���:�E�8�Л��%3���������&�Yx�F����n$1�K��SX��E��0a�)0�)�o�h�C�+�0$�B�3���p�
���
Ǆt�y��1�0HV�$/>��>̢�R�����7h @ #�R$Iw�v�u�>��S@��ff)���������8�.�¤h�&4�s�\n�a��8+��B�b>}�>W������Q*s�$�b��%0f01�7JbT�$%cq1���!F$I8u���2f4E�9U�@f��1ܒ�p\��c�$�0$.F+CI�H�! ��6�Bo	���C�C��&�K�ή��vGN� � ���D.5�cn�̈l�)��Y>�ג�w�}ɬs�}�H�t���5�`�bƸ��,aK���~-3pF86 `�A��N8h����$#�Q�"�����
���ؤ�`Im0baH��@#���$	#�X�$ @da>� �T~ʜQ-�������Պ�*����� F�A�� � ��#1%�e.3#$��t����)�,`�6�H�$.!q����H�`�b3t�d]@��_
N�+Q|e1
�p�2�W��:lG��T�y�p�"�b��bϹ̉�9�e�R�)A=o�2 ;�A$u�bL�ã�A�2HƸs����54Bc80h��'�Βa3���e����<a�|Ԗ^B"�8���L)eξ`�M�&3�����.s"BϠ�����m�	s��Hآ��V%T��q5�IS��P��ɧ㜉T��I㌸�$!~�faH��0�˙Ld�B�HrE����BJl���$!��3�o�n\�8,%Lv���қη���� E��`�K��C{ɣy��c|D#BE�$z`���0L���yw�0�b�0��u�\���4�"G��M�2�f>�A��h�
�F�,	
b4�
a`��
R8���e�$bU��+"Jj���/٦3���&@�B 	���a�W۟-�������lqW��ds�#��}>��E��@a�)�HI����YpD���	��-a	 Vh钦�@�B��E�$�CdqO�Q_�3-J����K�3%�>� WY!VBD�d$d�D]ƈLgP�.L�B�"���H�)�T�Li�Ϧ�Ӆs��ȒO��_�7�ۚ|}�<޶|!��H�ad�%VB,HVa`^bf����i�����."�!]1�Ĳ`Y��x�@�`D����!LR\>ޘ�D��j��B ęւ\fc_trp�0H�,k�XA�>qY�8��!Yu��ޯ�MA�IM_f~RDN�i �y�
3k$��H��@��.	�������7�G	�]����AZ̼?=��(��t];�\BB� �G
^4�d�[U
)iRM���R���	 ��yK��Jc,1�NW��k�f`��~_��G����a�� ��(�a%	YXP�Q�� B�$.3Ɍ��S!L9�%b�b2+
�Xp�l���!)�2�D�ƴk2I�]Yy�O.f��D��0�{W$H��BR�2��&�tsx�$5H�X���8�2$1D!���r�Y0B��(bBF4$tf�sy�A�@�b��$cF0�����i�7#̆���0e�$f\i�5\H���CϏ�J[��$�R1�~��3z�f>w�8��
$(H1$I$F8�C�7�ؼ�9��@�|��oL5&��M��^nm#�c>�L&CS��/��yk,'�;tdCVq!�6��8�B�j�1i6}+݌j�*B�PbH�BA�RW�q�w������
B��&3���0*�ڟ*ŉu/�&�CS�:'q*MA<Wb� ��s�m���/#���qzך�������U��3>����c���nS%!Hd� ��&5F�C��1`�i��Js� ��	Ć)�U�C[91� `��ϡ���$ `1�0�a�2�p��f�9NS0a��,��`�dh��r胬kI
%0�Būʑ1��7��.tˊS��4& M	�8����C�2���Y~���~ka�@H0"��A��X���a 5p�+"AiRRK�H�� B��$������
a�Q�	pHA�&��Ez��O�q����hn�a3��x���4��%pF�
�`Ę�i
2@ Bp��o��@�A�+�+��1�G&A[ؗgo!�K��+C�i8��$#VHXЌI0��FH�%0JƸSe�$
��n3b"`�$JF�cX�,	��`���X�ս�0�
0J�.s!)�G.H�)�a��ֵ���م�3Չd�b08�X. H�,(A��T��p��K�c��ˁ8�#�x2&>3�'s��jA?"ը��T��>T\0T�$$��a�p�K��
���B���BRq���/�Po?#*2v�����)�q.I���?�H�������w��3��9��p�$�Jc$k�%9#@bA`�e�vk�jCP6G��q�XYL�J@��0�,��X0"6,� C#����"�#�D"�b�a�!"HF!#(F!",�W;���
� @�aB$�!B�R��6��}�j�l�ou���L��1,ަ��~yu�u�ȭ��߽�Bc����ś�.������I8�O�l��o5�����]ƿ$��FCY����ġcHR��w#���ԅF$(��`��.�hS�0��P�CR��IX5�
��`%���0�P��c_'��l�0�$pF�)�&�1�����0|BBĉ��
�F�bU$m:�u ��)�z@)� �B��K���F���X�0��D"acLB$
�
��ˈ��!!���F�!�B� U�H�j BrB�8��k�e��\�*Ć �H !\�:��{a_�1��|C��D�̼��&~���>����K ��E�Ą1c� K:`b� ȋ#Rl�d�6bj�j�$��h#�d@�dq�a�b:1p����,�������0`A�e!!H���RV$5F�	���\�O��mt��Ǖ}��WW��%v�%���T�i���%.(YY��1$�+&�	m�.\q� C�58p�8�CiK�_��*'�NVeeee�e*H�$ D T�IV�d�,,�$+0!,�$1�!1jC�HF1�� ��W�bHq78��H��	dk9�L0����q������� F$# ��4 |Ơ��C�QFX����r@�2C&�2��C&�ox��	�o���{!�I���h��+�?@�C�\b��qB��X�¸2�|^�)H1.ك+�F�Z� ̹�Cl�m!D�	M���!"1"0�i	!��cdB"�����@!��0��!L!
$(ĩBJ1���B��ĻH�q� ���Ld�5�eLHW��V0 `���I,`�a!�,"ĂP���R24!^n+��	͚%Ld�"E�)�T�C) ��IL!
CW�����s�s
a�0��#a\�%�M�2ƘaB,k$)���.xO��r�g�0"E�D�+	�B�A�8�q��F��^�HHƘ̲1�
��Ł8b�
FHP�	F�nP�cXS0*�)z��I����(0�'�B��+Ro��FE�a�0�LGF�;餔�*Čn>aq��P�tK"`Πc:��ވ\��i��!I��H�	H@�R1"@�,�aHP�HH��a�22BВ����������!e�!@�B$d�d��q+0�$� (�A ��I!#��b|BN
�[�u>��W��Ԇp�n��:����8'6H\�C�j*8��>7΁�R����'��ܙ�}��9��E�s�|4�D�eHXV$�. \�IpJ�$�ۙ0M`�2�h�$$$R��GhK�|kP��"\�93Cx����b �?r�o�%���H65 FF0���f2�c��JGȋ�&ТB1�#?+����D��pJB���_�  �6   6�$[% ���)r����{k�հ:�:�{=��g�m������I*�N�s��ζ�%�n7f|�Z��V�xвP*�T�.e�XV�.�ӶȋUUF���J� ���'&๬�h��5��f��6����g������Z�d^שc�Y�ej�(�[J�����j�hr� ��Ur�pR�6�3m��!i�7m��$4]�뮶�'I 	��˗mk��U�!ԵJ�K�G
����r��+�6�tU�qj&6ۮ�ej�|�*ѫm�7i�6Ne�`6� ~�g��>�}N�e&Wey^y�ʁ*�Ѩ.Ie��6Ͱ  m���h6� �!6���` 5�Li�6�4T�)�- �	- �e�M�L�  ��ڶ��� Z���nm�� 8N�"N:,�m�d$�b��n�T�\�'Ke�RYV�@ Z�v�e*��o�o���^����W��E$ �H 6� [@��  f�i;m��ۭ� ���Z  lm�  n�텷;�7ZnB@�n����:���I.�Y��sm���4�mm�m�f8��:P��� 7mnmm	e���V3UJK>c�[6����v�H���@6ٶ�헨 m�� ���6m1�ml��6٭`.�V�#]g�Ͷ�m�@m6c�[��C�g��d
��  �8 6�s㏲ D�޴�   �ș:�	@T�:-���nZ�
�h^�3m�m H B��Mm-�׭�k ��($�@�#�^v��(��v�/�[x� �Z��Ά]�n.[���6W8�8�͈���^H�R��,�lpWAg��X�����4�z�	��8Ί�]N3֠�L��t�<�V֥�Q2D���pU�uГ�z�$�؝���pGU@C���0�m�9���p-����@UU*ڶ�V(�C8kj�N�j��]�k� �t��9mַ5��  n�����zж�����m&�0 IrP$m ����m����� H E�[_ -�D��H�`�&[q�l ���6�-�m�  m�"�6� lm�  m�mU�T�PPT
5�2t��`m���:   �f	t^��L�`�$�i4��6݀ M�V:��۪[Wc7.mm+FC��mMU����o���ܛ���!��Ί���YZV�k��r��{j74��s��'���:���GAU[�βsr���Ի�Y�2��m�����8�4�r8ۮM�ҷn�f	�HG%]�ۺ��Y�i�F�ry�Nb���ݶ�2��/`^h*�A�,��~�}�ӡ"jU:��Tr�U.���ko@u[r[r�E�y��@�9ݚ��9k�������m��m� Y��݀
δt��۱�-SR��4�uJKu�T�Ԥ�*�*1��K�s��:�	�k��@��R��2[�ŷZ����ă�l�@l
�/Tr9�^0;c�`32��T�*íL�5U*�[��jhR�W��@ RJ[v�J�m� ��h� �im�j� 6�  m�!�,�B۠ v�~�p-	 �i6� 8�`;H䃵�ª�v�+)n��UC��d� ��u� �`[K�Ai��1��٪�i�m*����ꫫ�k���q�4�2sfe��8��i�����9�6��Z��kr�E ��q⤋HԅҲ��wm��B����U��//kUU��R������y�mYH���F�T����:ٟ%�����VV����{'T�1ζ��3T�6� HX�`[R��ddN*��:6��NR�U��ز���U	3+T蝰p2X�U�ׯ�[~����>v��U�+i�W�;y��cm�U���X 6�ڶ]6�m{iʻ �[g�M3��Uv�� -*N�ji���  '����� ޶�6��;m��lUUU*�e� Ca`�U�U�
Xv�R�TP �u�&x 7џ*e�f�`Hl�N��m�m� 5��� � [AB�n�V���U����J�� �R�e��i�d�ڛvi鄀Z�P��Z�{dTTm� �Mf� �u�z� ж�k`$ 8� �bCm���ڶ�U.������l$�h m[ -��f��`	 jٴ�l�  ��    [���zj�l�۶M��-�3��Z��j���j�Ȁ |>�}l����\F�� 	i�kX ��b��S�niV�	�IW�eZꪜi���eq�m�84�l�A��:��U�ޖ\&FH��vێ8�tͳ��k�e���HUm@*���fnI+m��t䒃��tӦ��v�m�6�	Kh���
��:�~�D�l��u�[[ -�4�h)!F�� �����i���=cf��	q��S����@h�Y�h�Nb��֩�+��Uu;���l[*�;+V�@bu��NM�s���m�ų�^{p3I�n*ળ��e]W��0`�C�8f��	F������5��}�qeұ&ݷM�Y5�!�Q��F,���B�y�A���qu�É@�����q����,����W1Rm���WZ5��$��n[�m��M�E6/��K��u��t��l�  -��Mp�5�I��D�C��rA�-ɤܧT���. n����o�  [d  ���Ce��m��ڛl�.�kn��WH8��l��l��<hԀ��+{i�Ѯy�F�{���ݲCC�M�Y���A���%��UE�\M��S��v_�[��bౕr�vF���vV
��+ɥ�c�X6����U��d6��T�-)icg��b�ݪ�N��)l��U}s�|� �}�W� ��.��MC�u��%�j퐗��wi[Hqm�kzܥ#��r��UT<�48�M��rIx$-��ۄ���s��q"KhR�֮m� ����Y^�[NU)[k��IÅ��kT@)�N��۵T��U�K��X�۷m+%�A=r��J�e�*�gjVv%�P6mS*�m��7�j���X����à6�Z������ �� ��X��H��XN��-��:M��&�(���[��d U�x @,�-�tw22d��V�媠1��9���o*ʶ�-��Y���p�oZ@� 45I���U�m��t�M�D�L"�[Gsn��M#Z��$k0öY
W.ڦV��\�v� [M�`K	�a���
��%q2[A]�kiye]��+��v�1��fU��l�l���Ŵ�lDZ$�  h�
RZ�����W � �eMI�Ύ$7}	�n�L��]�
��Շ� �˗t����o%��Y	!#nu�Yl�cb,R<4%mDܡ����j�ҫX�]�"�k�a�� m-���GB�UUN*�R��!`�p:�:Zs��Z����;mn�R��TyU�V�����6�m��:�\�6Y-�oU�Kc��Ŵ��	1J�cm��n��,U�A���8�UivZ�T�Pg�����p$m&ĝ:�m�  #��l   mn����^�F�n"�[ma��ٹ����4���`D��l����/$Bt�n��������KStu� Aw��4�ɴl�g�z+[\�6]��,u�J�]�`L�&�\.Nj����b�n��8su�ۭ�I1&M��Z� �+Nͤ'F�r�uP�J얃�[�m�`hp�e� $�+m�Ŵ�����Hݵ����Im@m�  5�4��u�bDI��lUJ� �+j@�!�EV���[��a�
��UU����T���v�(�����v�H�]m�p�z��Ä�oQ6u�Q([\���<��;v�m��c��j�)j��J{ �V�PT)�mctKs�6��j�yi�j��w0	#Y7<kәy}���q�I�h	:F��lU�,=�Bvxv6vM�+Ү�9��xW�{kiv6٪�6H�e<���i�[j�( ��U����l9��Ͷ[I�:��Hp 	�V�j�l�VʰYLԭU[�!��*�~�?�@��U����;� ��     	9"۶�p   l�l�ꚛ�� 5�e�pm�l��v���l+� H ��Ñ`m�d�N���Xg��K(�U�k%�6Z     ��p��M�`[Z�[V� [Im��I�l��m+�`s�j�[@�`m� [԰�k�	 -� �]�V�6�ְR��` �j@vݙ��t��+�U����(r��UmJ�*�P�T����P]S��� ��[*΀����m$�j9����Yy�-��zBF�޺@$M�����  ��jå��A�����m��t8���zzl�d�Z-���:�m�o^�m�-� Zlm�	$�[d���7B��	$	�����  � m�o-� ��׮��m�Hp  _��>� �l	 䎰��(6�&۶�[@�f�ld-� m�`�,�$���  $ְ���δH�d�e�s���#m�q��������������bd ����U ?�C�� _�Q$$AȎQ|�T���|�.p��*�̀!�"myU>
�+�Uu��@ &�C�Q4�J��M��ڛ�Hq\=P����*mr2��zp�&��H6E�8� �6�L(�кR#
v-r��� SH"Q�@C�UaB|��/�q�qM�M|�^��*�P:
&����
V"��0X@L�
���	�2�P1�P
@:"B0bA���~A�)׏�42���tU�	������2�?$W���������!G`��8�D����&�P��2��"�M�H	�:8�B	Bb�@t�Cj~E ��Pt0�Qʩ�/�$"0H� �� �|��#X�_��<� ��I�^�=��Q��FDML('Qj�^���`2)2�P8C�qP� |&�W@ĎB�(p?A �I�P8	���TW��$غL!�aT`,��	��)"0vb) �0�Њ�p�A��I$uG�S�q
"dA�� �*�
�2 S�h��戠��G"B�b�E�,�Q"���&�8@�"(�

$ 1J - 
�_wowx��w�?6��I�W/P�7	!����1˵�iN��Z덻��0�:]�+��cVz�^v�lBw8l�Eiv�n�Jw`�56�m��y��;�I���]���h��Y;�#� T�nqh�2l��ֻ<�-[p�hГv�ID,��X�م��N*e�(�]G;-MI��m�Ĕ��nb�
���U<Gm���&�i�]�|b`t�Հ;c��l�kt�Wh4�eB ,�FAK<��X$I�ɷB�m�Hŵ�YG���]"8vUss�f�q���l�v��^"Sh��u��v��t�����%���Ιx��2p��7@9rtg���Y�^krK�S@J�����[1`�G�[�P��e�=�Fn�#��=�a#pu������˻X3C����֐�1��;T��mU������2�d ��q3�,��@*ӻF�q�mV�͐�2mZ ���6y
2�:&Y�V��Yiʀ�T(���n�1�m0%ٺS�W4�h�(�܃�s>�Mw����sd�O#\m�n�r�8�=[����m��q0h�N�20
c��\����M;�<.7S��Ί1��g�=Z/pWd�K�$r�g5��m���A�]<���L��Z6%Mm�6�P{er�m�&�u�Xם�U��i9���kvъ�����!X��:�p�'9�@�����\l&��P�z���0M+9v��U�[�]������չ�8��͈�`�g�.];Z6E&���m�²��kQE���J����$��v�kp�Ý�b2�uλ%n������h̀�6�3�� ��[5n�"��q�s��\D�6�cq��6B�cԾ�n��Ÿ;i�sU�G��n� ���*��� j�Y%��ܸ��Ŗ��:��VV��dā����4��(WlԪM���s΅���|d���/X�ْ7n��q�>�n�u����':* (tM�ڷ�lBFk�X��m���w>�s�{���O
#��
�t y��&���ʝ@�@�;�:D��������ox���iLZ�]�qs�a1�m�L�.im)�ƶ�;x�vni�Z¶p��b�dv��c��l���n4vѱ;E��u���p����8Ҫ�0vĀlRɌ]c��4�3m��ݰX���g��u�h&$Hl�	��v��p�OD�n�6�ZCcf��xچ���<5���l��u�ci���m��':C����6�q1#���u�׾���S۷Ɏ1ۑʧ	�rs�y�p���+�EWl��y�9j�ϳ73���t��޴�ܿ��Xl�ŀw��$��M���)eX��������d���)�����1+`�&�GL�:`v�u�l�{k�i�*h�W-�?ow�GL��l�D�ݩe
^eڴ��K06H�۝-�wH����.s�O�ע�*�X䊸�
��b�T��<��a'V�d��-�d���vz�&�Ӳ���b��e�~{7� ;�ۀ~��,��ŀD�)5��2Z���s�V��̉U+���*!B�$%.�U�3���x��]s�u��o+m�(*J����{����XlDL�����o �]����-Tⲱ,��L�:`{�����S�wߖ�k��z�7C���`�:� ;�� ��x�6�`�P�u\��A^[X�]��g�ѵ��h�1I��xŷ�^M'&mír�����;[����Oߓ���d����l���_+R;PJ���q`n�,�gu�{�sˉ&��k~D��mAK��&�����RM�������1"�b�(�$�B"Ei{���{���Q`A�,�*ۖ$���Ζ�;�LwGL�:`m�_�+
Ɋ���������ŀw��x���#�����S�HIۛU-��H��h�i�֭ՠ
����z���"��M�(*J�����q`n�,�gu�{�p�hl��U�R��`m�͙8���{��}޼X7��I�����,� ���x���6)�7����,��XU������"`{�:`l��	��*���\��~�����쯖)�
�v�����0="� �0%ʏ��]uG��"��-ړ����tv���S�_Qn:s���#���=�줕v㊫_��ŀ|ݳ ;���"!} ��X}�X~��[r�j�?n�0�D���遲GL�����d�aH�L՘޷x{׋J&{���nߌ��SyX�-��d��.$�^����,��޷x'�K���j�V)lnU�}���۷L �wn���;�RL���%T�ww����'b%�My��<Ŭõ�

�N��-��-�<m!ʴ����n7G��������]<��;Qdf:�ڀ8�CEء�ý��� Y���խ���`1*T�P���ۋ�a:�iۛF�C��Lm�-���@c��P����a�y�t�OF�^�[�n��!��{�����T:���Q�z��2h���+���c8����g?m��W-~=Ǿ���{V�N�<����zS+�نkj�n�qpM�<��L�]}�������,��o��� ;�L$t�ސ���&�����L��ŀwwq`7l�?ok�+�Gj�[n��q`vGLH��7�Luu��Q�k-%B�7ukb"IO^�� ����w�w��Xۡ`A�,�*�+���zD���遽#�꫕�.I��I�v��HᶢV�g��j�X�ۊ��,:�X��:l��ܱu����׻x{׋ �[Ű��	} swo ��)�U��KUv[�w��Y�.x{BH���E�!!��!.a0{��1�%�>ѩ$�ۀ���>joij��V)lnU�l�� ��0�10;�:`v���{`�#hw���q$�w޸��D�����#�������"���0�107z:`v��{dL��o���s�	�ݪ��-;&6W�	���I��Ӻ�c���V�yf<��v���w��l���D�7���w��U�$v;jN�V߷q`�D�7������Һ�>Y��5swk >�w��sxD, ��3s��E�}� ��ذ���Ԥ�X*ee�� ޒ�w��l���D���T��M�@��e��ﻸ�쎘�D�;���+��f+�����L����5�n8�j&�5c���s�ŋ���Q������R+I%b�Xܫ �۸��"`�b`n�t���W�y2����)eX��۞I�����;��,�n��q6w��º�>W��p�����GL�0l���ֲZ��+1b��V��GL�0l�RN(�
��#v�*�}־w ���z�+�ڛC�U�w��X�)�wo��ټ��ŀ>S(�\�*�6W��غ��зu�t�^P.��S:	̈́�����>7;:wK=b��m��?&�]�GLt��u��ϰɊ��$��tL�0=�5����:��49S����VUm�$���� ��0�`z�uGV�X���V�����n w�v�}�� �޺�sccq�;�YS �Ș�tLގ��0=��%)E`���U�0 `���~��G`-N����`9Ї	��<���ӸiMgmnv�r��F����ZD��[��SnH�J8�f�8x���f����5��S��lD�	��=���>���ڷd�008��m�c�6u�Irk\s��sa�3ֵ�B:6w]�u���ΆNv�ܚs�R���M9�Y{Vզ��RĜ�� �ˈ�k�°����m�S��-̜�_�{���u�}��e�q��N�V��]<vZG���6�V�ݎw�KB{�kq�1-�~���0=�0���ٮ�I�"�����n��?}��l�������+1Z��]�ib������`z�����>�B�G�VKc��V }�ۀMΕl�:`M���[\���>YX�$���*�::`M��t�p�F����,D�H�-�yS����n�ur�n��q&�Ռ�-�<����8��-��%ҹ�ີ8_^,� u�ߔ(���=پO �{h?)VGX��r�$���(!�(�0  ���!(���d�u��I���˩'{�ŀo��͍����)eX�wSnt�`wtt�����h����� 0X�nt�`oH�7���ݸ��l|��ETce�<������� �"`MΕlvL��> {�؋,���ܸ�q�x�\K��]s`���qh�h������X���W}���z:`$L	�ҭ��GL	�Բ����X��ڰ��sˉs�����)����:�f�Jdr��lQ�WA)e� �f�<�����\�bW�E��g��K��HEH�-�>���C���Cj�@�b���2bP�i��1������R��̒�x|16�.�c��ܬ��É��Ʀp�`\��mӲ�{/��#*P;Пe�!��0�pg!���1�n�h7�$n�DF	#!G�:A�$�_��FIa���D���`�BbTd9,Hɐ�۹�*�$x����+�����m��&�D��LB�d��0�9M"k@+�C��aD4&ÃcPP��J�:�T�;M(�����(=JP%	"!.%�K�ŀ6� ;ƧPT8ꪵ/�<��ŀo��X���.s�\~��'�|��7�5U��V%�b�ގ�t��7:U�6I� �~�I<�@�9`�R��Pj�,�'K�Pۣ��gnl�J�V+��6���2	(��.�| ����֧ �o�P�0��������ޭe"||��Y-1���]*�뻾�:�����{�ww�4?˜K�F������5	U6�*�6�������zz�뻻����.�~����U�RWU�6����}���~�۷��5m�}�:]�ۇ!"E�<�V�V\)�o��5m��8k��!�,���W�Ͷ�����}�}���6���������l�����V(����1��S<�!m�v����.X��.�Sy�\�X�'9e����cm�ݽ��;������oOW�ww}#C����J%C���R�YS�����q6�~��_�6���W��#o�_x�6��{p~��T��R�ICm�wߗ�ޒ3}�Wm����x|�{�f6����7�H��,������ߕ��oݾ��~m���6�߻����ѷ��R'�ƨP%���ݘǹ���ݶ�D���ܟ���o����{��8���gV�k�<�V$���R��IO����Z#u�A2���9'�l��(����n�lO{h�٭ ���4���#��N�U�a�&6x�H���K��j����e�b+=��&ݸ��oG7)bNmغ%��C��Zt�X�[�8�vyι۞�I���q����ݶnt&���d5�ɒ�9U��:r���;Yw7N�H,�u6�46�N:M7�ؚ�㓝z馢�^���22�-T��m�\I#��IO�1���ꨎ�el��n<�s�!�s��ԯ�\�=c���I�F�UT�YS����?����1�߻�����Ѷn����I���?ߛoڊ�^RWU�6�,�3�F��{������b��#o�w�����w���0m�n�D�V�c��W��䑽�e1�߶��_}}��#�$�}���m�'䧫�9b��L�RF��|��ͷ�z�<��o����Ϳ��;��Lm��w��U�-E�vT�~m������m���z���m���cm������F�}ry؄�t�v�,�&��&GJ��-s"�%��s��-�:���6��)$j�c�R�IQ���M������}�&v*��{��(�\�L����T��=�rH�D��(�_�6��w��O��8����?���g>�]����l����{�7��Dy+�����dLLJ��*f�̙����)��UU:��33/��-K������1��}��|)#�����������\F7䤛�����m����ߗ$�z�����Ȋ��%u[Sh��Q�\�7��~7�m���3�7�[}�������tO�?���ÿ����q���ݮ��.� ;E�]'k`�Hsq�-Q���)ȅ$u''R�\�#�[,U�Wm]�m��������o�]��6��n#�.s�������#zO�OW`r�G,��oݻ��~���}q�o��~_�1���ny.)#m}�G��9hWK�ʟ�ͷ��`cm����~��\�� �J�^AZ�)�'|^r�syέ���׭��νrF��:�-��1��%'���~ݶ���9ն���v����\{���ն�w�rz����m���q�ߔ���o�[o{�jM[m������8y#�?+�`�Ӥu��=z�m!%NR�4�&�a�N�Yx5B^HE[�*��K��E���>5ATH����������}��6�߻����$���F�}����{q�Z�RGU[&s�w�m�;�I�����@ֵo�{����m���έ���m��
�����I-��6�,�1���}�~��m��o�I8���{<��ͷ�{01��{�x���b�r�j���两�����H����n�m����5o�� �����*�.s��ڿ~m�Ѓ�S���Q[l��۾�]�{��xO{���[m�;�ݶǻ�礍�$��S�{�&8�UH�,m�H:��:�E�mĝ��^�E��1V��v��!��r��)jd��������3-�c�;�ݶ����;�-�{���ݶ��Y�F�RZږ�ef6��������z��'w�y33?w���<���v�$ͅUޞ�9=����Rʿ~m��}.7m����o�_�!�kZ��Vj�o���7����G��
��,����{߽n�m��}�5m��s�7�o�_�g�c8�o�a��ㄎ*�m��~m�ws߬ն�ʉ�{��Ü��{��έ���m����K$�Ķ�]p���A�6b��r�� �hN���.�#�������o	�%��q�څڧmv�.�(�6�Geu�=R�mn�s��1��m�C�"R��Ň��	C�	ex�tm�4Z��l��.z�>���i���|����z�u�;I;fv[Hc�:�-�Y�m�X0�YD�c��z�H������B5С9�s�I���u:�3,�5��������Xt�a�J�q���M�n�[u�g�?u�g�.�]�x�=�w���W�I%�ڛE$��m��������������o�{<߸�%Ͼ�������F@M���c��W�Ͷ=�K��ž��w�m��Y�m���ٽ�UBH�H٩OG`*J+e�m���7������Vj�*��;�ݶ���ն�������Z-㔯����q$��K������[m��~ٽ�c���3�n�@���������νg�*��Ե�+2�o��l���7ﱝ�e�=�[��on�)�����}"��Ed�RK9*e^�=m�6&�\X-t(��Q
.�ּ�=ޟ�E�D�C���}�m��z�m��nk�6�^�)�/�9'���~��}��G�|j�d��um��w]�{�p��F�Y��!�"�⠤U%C��//�cV�~���7�m���s�"����ﰟZ�Q�Q6��~m��{F5m��s�7���s�}��s�m���?������My�X��KT�߅q�s�����w�έ�����v� ��~Sm�u7�[,U�Wm_�6�g������(�Iy��������b���������m�t:�Ѐ�T%�U"S���E���`#sq�-ʶtv��Z����w���Gb
J+e��m�����wq`޼[��wo s�Um(��,���.p>�Y��S&�������y�..6��O(�dp���eX��hԒs��u?PBe51 �Q  ��F�Tf�w�[�'~��~�\rl��6�yK*���9Ŝ9�	*��o ��fp6�`j��Q;׿,�i�3 AT8���[�5B�	ww~_�{� ;�� �7Ut�X��ygeH�׮����v]���O�h�P��P��N�ȼ���	��q�TNB��~��� |�ŀ}w�%��o��5l5�BGc����-X��Ŗ�B��o ��fp��Y�'u��	�r�b�r�j������o��U��b�<�ذ�Q#J�M�*�wWx;�͙��ŀ>u����%+� ®�\%D�@R��)TppT�i�����u$����E]�e�M]��m��<�8�{��}�\~ۭ����P�����B���k�ե1q.��Z�9�,�8,X.��d�m���Ӧ(�I*p��Wj���ŀ�v���oߘw��X��\s�EC��լ ��ؙ7�{3�w^��:�f���O�@>W�T8������^,<�Um=ŀ^��)�ws*JT�L�]���Q���� ��b����(Q�^~��8eNϪ���WJ�.h���>u��<�	V�z����8I�{��St��\|HGb8�� ��°"� ܑ��q��8@�j,�"_�ms�.a�)���`�MsA�G*���E���Z��5R7|ւH\C�ف���g�}��	��Ɍ��/���a0����w�h��������L��ai����H��`A�@�21�`Loa���i�
K��&$)H�S�xmi)B����� A�	��BD����$b1XA��a�F����ٸ���Yd�fHP�X%��H�Bf��� `�R�F�Єa aA�RXSB��c�l�A��B5~ ��}�}F��)"�#!,����Ĩ.'�$���p\\Nv��o�~���MF�aom� �,�
�*S'/:� �Ol;�p��Sn&��cnT�=��,��w9j���X��[��*�uQa�ΡY�+�bLe6�;rU�Z���-`�q�pKz�P�Xruu�/K����-��N�iР�f�G�r�]4�V22e����932Ҫ@��UZp�t�K���	ɳZƙ��ѹjNj�h$��������)���$�ͩ
�+]��V�eZ
`�$��&iw&��VW�^���j9�m�F�N� �JAjL�rI��ҕμ�v4z���V!�E�5�M�nڃûv�rݑ�K�����5�\�v\�5�t��z��ž��T�1+EU��A�����n0�JNkk��v_C�<D���<ң\���>� Dgf�U���p�C�bS��u )Hh�+t��e��{O-Z�R��n�!��J�N�=����N����U�r� +ҩ9����*�R�`�XU�O[��c�u ��\0v��2T�Q��]!J�yۇ9�=�nK�g[HL�.8ܘ��^��`:)�N8X�����Iú�r��6W�$Q�de���>����nj7(����h���R�T;釞�6�ь\���	�b�������Μlӑf��#�:��C�s����p��S�-��'#��d.ж�M����7���i\��fҌ=��S�l���8٠�kp�b��z���<�,�vR�)�"1zb��n6;m���nF$(��8v�(�q��=h.�f��YI��ۣ;`dy���Y�Pμ�N�#��N�-��m��$����T�J��/\�TP�Sۓ68ƛ�������E�K4�1�Zy@��I�n�J�69�u�v��]��k�-�v-�L� Q5�u�p�D�Cm:6af���ˌ�F6�*L��nUHW� �l��6�XZ#WG�z[d���Zv�q���`���CeeYy���ڷd݈�7i[��Ȓ\G��? w�ʿC���Z���=�<Q��V�6��`� ��>�3p2f۞���UZt�:�Ҏ��D��ր�ظ)^��g����,�k�⌏Y���խ�\�Վ�961����[�͐����[�<h�7�C����#�-���;��q����,�3ן%��ڮ��k��`��g��[ey#^��1�Np�YڂzW�іyꎤ��H�qp���^��"Ѷ:'INI��� 8e��B�R{ߏw��w��z��_��4�n6R��6.�.u4�76.3���Z���-�:wܽ����D�2��X�v��o���7�g ����_Ho^���jU�7H,��]����~D%UG5�,x� w�۟ɰ޿)�q�Z-㖷�}��X�^,=
!(�*�w}x���8 �t{	%dp���eX��������>;s8�"y��,{�sS[uJ'�yK*���p%����f��7w �׋ ����r��Y*�Uۧ's�4���sSc\�'��7�b��u]�w(/s�"ڰ����U;o�=�_7�|�ŀ>u��%J!r���^�W������M����}��X��$��@�p��3��jI9�z���o?���)yG��RJ�W[�n��ŀ�w���Z��g �ŀ}�N�OaK-U�WmX�{�z�����m���D/%^{�,V����v ���[�o�u���_{s��=��, ��ۀ}��q;Gk����S<g�9�w;UW]�=%�u�jb6p�A{F��=��[��q�Z-㖷���� �׋ ;޻�$�
���w� ^���UrT�qWuwv`�x�TDB��}{x�ofp�m��"��M���L��E"hw��� ���m���|�QP�(c<����'��jI��c.jQ1s�M]]�z��%��3�w�~0μX-Q�Sݫ��d����Ȫm������o9ĵ�/������o >��"���K)F��lj��[��iȼ�:�kn��DmuŪw���28���b������ŀ}w�>;s:�} �ޘu�t
�
Yj�r�j��v縓g��1`���~�Ş�5v�S�؁Y�%�^���nهڢ�ow 7�x��R�E]�e�MYs��P�z)��x�=��, �[�G��B !��Q�!)������x� �Χ�UZ.�K����� |o��������p�n����l������+<V�#��Vn+�{��ϙ�N�4�m���]���U�H��4;�;W��p�}��y}Ϡz{ذ�<�W��*�-� }��9�%T?m��<��X�7y�$���Q����H�#e�<��� ߷qa�7���=�|���T�7\V*�q�L$��}�� 7���7����8���}��!�RKUc��V w�w�yD&��(����;��{�RD�� �  1i��qܘm�vX�\�j�۬�#4����"��T�<wn���R��$��ٸj�jkg�:�5ڍq�+�]kL�ƞ���zE��D��M�[�v�0`��k3��% �+mc8�8^��%wo.�JMd9�иԲ�������)�n[��^��랤A�fV�W=�q��r��7M��0��[�[gstX�V�X�����S�sú9��� �Zh'���wwt�����Ņ��ʯ^W`�n3㛪��7a4k��ܽΕg���ԦGb�j�o@����|�l����"9@k�^ 3|�Q��˸��' ��ٞ��{�� >�� �M��P�d7fv��	��l�� �}|`~ݸyqqo$�����o���drk�HD!�G)��I%2��x��' ��aBQ;��0�<�+�@r�p����z��߼p?_� �z� �ҥ��8mغ���姱;�n:��<0r���J�e�Z��a�u��{��}X�'���.쟀���>;f w�ޤ�&��=��O ���zZ���ES��S |v̕Ș��\J<�Jh7}���~S�q�fy(��BJ�~�&�G����\�W5V`�x�u��bL�v��=�_~#f�6;'kV�p<�8���8woL��06���o :?#�	�Z-㲧�}�t�?%��t��;$-�/C�2Z2���6�qgGh�&�JӍ&��4�V���c��:��V�.$�K�u��Km?���}w�>�dꈏ��� ��6�X��꣔���s˜\l��x���L�Y�!%2s�f�Ђb�j�� �[��}�avD%�6P�Ж%�"!�v���X��׀s��lo�rH�A���{��O���{��, ��n�9����o�~��]��vU�Sv`���5$����u�N��� �K��ޞ�:�U�J�jЎ ]�#gD���d�������]�n][��J����-U�W-_�7}�of��7l�}!��ŀ>�L�U�7H�ʻ�����檊������ŀ�]�z��G�
QW`Ywwd����0&��wH��B�t�&uSt���m�����ߖ n�����z>IBQ؏$�����|����Қ�
-R-*`�&}R,��6tt�|o����zm��]�qv�P+��8dBt�;�䈤�l<#x���5	{0��/��/��S�,	����x����n�����޸{�$���rH�BK�S�q��͈��M��, }{x�n�?���R��o�Z���EDvU�y�ذ����)�u�N�����6���X�rՁ}�$��n����S�}޼X�x��*e�N����Uuw�>�d��8���{�� >�w�yB�*�gf�]�V+�Eϡڕ�̬X��ta:%@q�\�N�֠ˎ�^��xn.8�<iǿϾ������mԙ��`�<��,�V��Zǈ6Sqc��S�u���m�^9�@@G!�P���\-�cN��4��N�-�u�ݮemF�ˬ^�SXg�\�.��'C�̎gm� k6�ێ�g ��!��׃��J����D[-��6ˮ�9��{I[�[����/��8�qKmF��H�)�:th���v�4ܒל:�j�z�s�����шȩ���,����x��`����ݾ�?0��xxZ����7J���n� ��,��T{��n��pw��l����z��`�yGj��޸�6N�S=oq`��X8�e�)��V�Wx�u��8[�X�x�<�G�EV�z��}U1Ub��aD�V� ��ŀl(��������k�����*�U�����lRڛ��{x��n����~�g���9Keٷ�����~|���]��GQ�|���`~ݸ�wS�Iq/�;��,ڵX��JGj�p��RIϻ�� ���2&�Dì@<*`Ȇ�p �a)"$�0&�ȩ !2�@(�da (Ф���@�R���(�#0	 � �i�"�\�~����~ŀ>;fj��%26�%=��V�pl���}��XyBQ���U������hqSa� ����������`M��m�����������:ҩj����>;f�DDK�����' ��q`���Cj+vp�NWS�")Uz��n�!t�f�6:F�R�Qv�=g���޾ٶ\�4���(�? o}�ogu<����?0�}|`ﯚ�'�ƨPr���V����lP`�'���������y\���U�]�$��8�� ��,1�HB��B$@�R��X��2q�=��*l��q��[R:e��! FF%	h����Y�H\.~��
b:����Pފ��2$��P� iM"��eގh*i |��b�~>��4�T����8���>7�@!A�@&]��Wb"S�;v��)��-EZ*TW $ �NT؈���N�߿\��y<~�nm��T�nT벬$��{�������O ���X��b#�R;Uc��V w���65��?�{� |v���9qD����c�q�:i�=[mwSg�@��v��p�[[%���(��7R���V���I�>}x��l�^�X���;�y�j�
.�n��� ��߷n����͝k��XK�*��\ݬ{�� ;��(^U^��)����`��C�"l���Qڰ=�����5��8^,���"���`��b�>��@q�p�}��X�`x����$ڽګ�Wvu��
n��������<Σ�`sV�P�V�(�EYY�-Wq�JR�B������ŀ|ݳ ;��R�A�z� ޻���r�Qr�[V�v��v��}��Y���n��'�J�U��� wo �k�NJ������w�Զ��)(���.$�������;��,��0�n�s�"�j�
��.�N�׋ �D$���x�����֧ �%��d���DX݌yv�;0ͬ�h1 ����Hڶd�@��N�gl���]�{e�3�{S�}���u�uƥ���N�[(F��rZ�����L���ڕ��gU�3>k�\P<鬝nj�f�����\;�)�cF5:;s�=z��;6z綴�>�Vk�qٍ�A��yb�M��%-�����ܤ%�<O��x�F�I�)ڂ�'g��������=�c}�z��΄���8����b��,=h�{�� .��+����*��a,Ct�Z�v����, ��&��V����J3����y�Mœv��n�a$Ҫ7kqN�{� ߷qg�8�g}7�W_�P�8��z� ��Ň�B��$�U^~�, ���p�[Mq�KZ�TV�*x��ŀ>7� ;��a%	N�z� ޻���p���ʡmX��� �K�q�}��l�'�}��X��{G	!m'mZ����G	z��D��v�R��u�vN��.�Èm� ����\r���{�\��' ����$����XaS>K� ���ۀogu<���*�x����0��
�$� _��ŀs}�X�7x ��-+�5v\�v� ��ŀ>7�I(S#���پO ���+�Y��T�J�X���f���^���T�8Q?>���"j�0N�U��v���V����lP`n�j��]�Ȫ�׆�7qgt��.Iㅬ�s�3\�Slu�A��{����]|AT8忀=��x^,��5B�@}ݼ��n�y�D�n7*���ŀo�t���p{�W=Ģ䇻���W	jm�UEݬy�� w��/B"*"T�BK�+w������.����W�^R�C �0�:a�﾿��~Xt#~K� ���ۀ�u^����|�w s�w�6&��Q]ڮ��;g�Nr���&��[mS�uě]@�\p�'ی���ip��^��erS�H}��`6�`9�~�^������W�u������K-� ������a��� 6�^�7� o��N�L���Y5k 9�� [/���wq`﯌�۱W�PU9n���z� �ŀ>;feB�	.��S�� �z�#�jWQ�ܪ�ow��	i�������j���C�߼�%��-��m�fΞ�5��7d^K�utz7N�4f�F�q=�}+��J��ݯ�������޵~Q�u�,�����VD9Gj���s�ˊP{w����,�Y�<��7B�|����]�����|� ��ŀ|���v���z�i�B:UGj�����wx��ޘ�7xQ�QU��+��{�tU�7j��\ݬ��0B�}ݿ�5�W�q���>U(Pu59��q���l�Nr� �yJ�UthL�Qv��9|��F!7vM��ƛ��l�d/hy5v�-�z��)UU���A&�mc������}o��kjU��K3�����0J�T�j�E�ۖ0n��Wkg���c�4:{Ͳ���y���gk+���Z�rv#^d�	
��4������v�b���u��s��9����8��$��: �6dT��)����(5�cP��یB��1rc��f';�8p��%�w3u�Gn������v���<��*Ȣp�N������ ozR`l��6(07b�J��/�RD��� >���Jd�ŀov������zC۞p�Y�A��U�;��ؠ�;dLwJLlY��#�FݥE�`y$��{���pz�x�DDz"���X�B�=E7jn��R����#�� ������E׶4�r6�k�r&�*nH��v�c�|s���3�uG&7x�<��p+u,���]ڻ������s����Q	/$�K�u�N /o��,�U�T�pM\�9�fRJ�%�/�K0�v���� �wq��ě:����n��j��V`ݽ0�M�J!B��� �v��7Bul�q�N���"��pop0��f����� ���U���TD%� ��p0����{��,�Ӻ��푵�q�A޻#�s�+�h^�(xI��k��1��be�L�Җ?�<�jaY�A���}ݾ0	�:`{s��'t`�݋3"�,U�v��$��0=����0`~��L ��sU�;Uj8��`��۩'9��MO��$Ȃ��!��$���o� �^��>�S#I�H)%I^+`v�`��������v� /n��Q�ꩺ^P�?o(0?�����od�loF	}Wu�0�6��ѻ\�u�QӝNE�c��F�9�mQ���9k���~{�пp��Xvn�b<����Ζ���`���t'Q&ȇ�Mڰ�N��$��g��oGL�Ҽ����h��� ������f��B����,�?������8rZ�0,*��\��^i�s�q`r��	��!Q�I��.>%�{p���m�mu�eR7iU�ـ}μX�K�	.����u��,�t����%��TFH�P1���g��r=b��ؤ���@-�f�<;�����'�#0J��Y���0=�%�=���t��8�0���X�`������ZҶ�A��U��gt_������-�q$�a�=O�F����x8U�w�|`s����v�g �wLX�,j�Yh��YXf!������-��Ł�q>�s���I��:�uSے[� 遻�oGL�qxq||D�+H�TL:p��JF2�:#�)b� k���	�|#� �HSy�4�ư�9&2��h�)���%�Dɐ#�92@%�1�3������#��l�AN/�w2���bɑ9>5v�}����g9�qK���"^��'
��p�᫗��� �̧<�qAIla��
a�l��AG�y�C����P��H�r���J�`�Э[90gJl �v�	i��[����۳m\[���]�D66�����[D����d�]X��q�m&�;66r .�����;j�yv躣���y�ٌ9ɛ���r#��,��˳h֣�[i�%ڳ����N�ScFll����^
Z�]��[T	��\ֽl��<�چ�ao/��5�s��۞���CМ��h���&�mv�d�����ф*�uF�� � �2K��1v��N��;qI)uJ�:���`�/m����N\��+���b�LW=��<z��݈z�ҳc�ti�v�gvi�0J:�h'�F2���J�r����	���$�j��HV�ج�FW��gm��vM(Y��ej���� ��!@m҉ō�����$������·��[8iƨ��s���M�mɆ�F����7������A{7g���sn��p�m�m��S5��<��N�]��(�ČI�*�m�������[��.�'�F1��W=�"�)9�lu&R�=�*�۪!���)��z�s�m+'e�MeЕF�g&�]�n�He煤[>�l�X��g1z��;�/-4�uhC;��U�
���u�ի.���\��%�7S��d&�#t�%Ր:���;�e�d�m�N�.Wa�m���X����f�2��IV4�ݫ��������:^,l���-)�&�(�nݐ�
�� �ʙ�o":�V0u�ĤFs��)��g Y�dٞ������.�5i2=h�yqF0oc:Ɍ�C�m�6T�\�,�1n%*�M��e]<U.^�3��t�@
��*�q�elϘ#��(7%V���ӘH��1α��n���8	�C*����T�meʹ�=`�x�!��p-'BIs%�8���F��
�L�+�z��iP��S���C��uO� �R� �8A�*|"��'\o��ĲS0���+��vn�)1��m�Ћ�]�	gv���¦���u.��Ӏ5��B<���w0�̶^l���Fn�Ƹ�r�9�Guuy��V^3%�N�7#l�>����p��Yq��id�h6N,vn�&����'u�9����J�:�ne�e��s�]9B��V�I4p��W<����.%��	,�*�Y`\[�h�`�U��V�}đĕ��`c!��v���3���C���m9+u����W܏Y{�w��eƫ���*�I_@��,�� ��x��B������ ���FJ��J�,���(0=�0=����n���/����g��GmR7iRI����ܒ��L�P`oz��j����$�`y��g����,��T�~X�N�.˴\�*Yx���t�������H}�ߎ��?}�^]t)��5�����\�@�Q�K,睎�g-V;,�9ߞ����~�:��V�l�&�_���}μX9MϢK�~a�}� wZ������j�1��&��tk$@��m�U��k�Ƿu$��w�f�q,K��=�M&�X�%��Lޖ�8��1ar�&�q,K��3�]&�X�%��=�I��*�bs����q,K�����&�X�%����`��ea���1���Kı9����n%�bX��}��Kı>罳I��%�#bs����q,K������͌13�bY�q��Mı,K�Ͻt��bX�
����i7ı,Nw>��n%�bX��}��Mı,K��4z�9�)��u��yn��Tѹ;�8�tl�L�6R�vl�,�O<j�J�B�������,K�{�4��bX�';�zi7ı,Ow�����1ı;���y���g8�ž�fN(HZ�Q�K�I��%�bs�צ�p��1��~�4��bX�'}�߮�q,K�����&���bX�9�g�L�g$�&33���&�X�%��{�f�q,K��s�]&�X�`oM�z�@ٸ�D�}��Mı,K��4��bX�'=���S&Ks2ˉ�I��%�';�z�7ı,O��l�n%�bX����K����Nw�����g8�������,D�Z�����ı,O��l�n%�bX���޺Mı,K�x��&�X�%���޺��q3��L�k�ݍy��B�D�%��^��.w[��R����e����.��hz^т���!nri7ı,Nw���n%�bX�sǶi7ı,Nw>��&�X�%��w�4��bX�'����7��d3&.1���Kı>�6i7lK��s�]&�X�%��;�Mı,K�Ͻt��bX�'����ݙc��Y&q2i7ı,Nw>��n%�bX�s�٤�K ��s�]&�X�%��=�I��%�g�՞��e��ݣ�W�_�&q3�H����Ɠq,K������n%�bX�{��4��bXp�P>�g��3�(�L"�:�O�kܺMı,K��!u���L��.ri7ı,N�>��n%�bX�{��4��bX�'=�z�7ı,O��l�n%�bX��ӧ���[�9ű�Rط2tZ���j��.+�K�Z��V��SyĒ��aaj+D��ל_�&qX�'����&�X�%���޺Mı,K��i7ı,Nw>��n%�bX��N���c2[��ٌ�Mı,K�Ͻt���bX�'9�l�n%�bX��}��Kı>�g�i78���&q>��yK�:ꖩ%�8�D�,K��i7ı,Nw>��n%�ؖ'����&�X�%���޺Mı,Kǳ<[��2�K�K����n%�bX��}��Kı>�g�i7ı,Nw>��n%�b����w�4��bX�'���s.0��2f��t��bX�'���&�X�%���޺Mı,K�w�4��bX�%�}��7ı,H/� �(!�����hD�&Ɖ�.XI'dH��ٓV`n�]L�[�y�&�mg;D걞�m��9��ZY�\ӧjw `���C�y�Y0Y�6�E�P�ƞ�q��F"ڜ�u*�A�3�r�]\�݈.,����z�+�͛��v�]��Fuju����yL'Wz�z���\{ZB����[=�ayu
.�Ά�uPZ�%1���y��08� �=L����u��{�]����>���D��[���p��6��i���`!�Gp��ʽ��:�:#=��ѯc9!�fn.M'"X�%��~����bX�'��i7ı,K����~@ �?D�K���~�4��bX�+�a?�%��1�H��/�8���/��l�n%�bX������Kı>�}vi7ı,Nw�ޓq?q&qo��d��q�j�FI-Y���g�b^����7ı,O��]�Mı�ű9�{)�$�}��F��I���j�R����X(@���.k7吷ı,Nw�ޓq,K��;�Mı,K��t��bX�'���Sɒ�̶���n%�bX�ｽ&�X�%��s�٤�Kı/{�gI��%�b}��l�n%�bX�9&e�����̜[]����\�Z��t�ra�h�^��J��s����73��Z�f����,K��}�Mı,K���4��bX�'=��Cq,K����78���&qyz�g��tw��g�,K��}�M&���@HR3��� 0���eD �bb%����f�q,K��s�]&�X�%��{�M���1�LD�9���q��ᕎs	1q���Kı9���I��%�bs����q,K�����&�X�%���^�Mı,K�{؛�8�,�I&%��ɤ�K��1D��~�t��bX�'=��4��bX�'{�zi7ı,O��]�Mı,K�����Z�c��J����&q3���Mı,K���4��bX�'���&�X�%��g޺Mı,K��U��)���=�.��t�$�j�i��:�'%�<��q���ǧќ��ɗɴ�%�bX���~�Mı,K�w�f�q,K���]�X�%��;�Mı,K�3,���g�3rc8�f�q,K����٤�?��&"X���߮�q,K��}�f�q,K��}�M&�~AHb&"X����~S�d�3-��4��bX�'g���Kı>�}�I��>�IO�-�U��01���D��A� �g"r'���&�q,K����]�Mı,K���s�,�srg91�g7I��%�X�s�٤�Kı;�k�I��%�b}����n%�`~��O��NB��$)!I��j�UՓd�,.[s�I��%�bs�צ�q,K�>�}vi7ı,Nw>��n%�bX��}�I��%�b}��l��L�6^ڬ�^l����ޚ8Li�h��s�5]�۪�-�˧���ޭ���{��oq����I��%�bs����q,K������X�%���^�Mı,K��7nq��Ysqri7ı,Nw>��n%�bX�{�٤�Kı;�k�I��%�bw��٤��&q3��wH��Dݥ�W�_�&%�b}��f�q,K��}�M&�X�%��w�f�q,K���]&�S��L�﵋'<�Ij�FKmY���q,��}�M&�X�%��w�f�q,K���]&�X�xe�J�U "�@�/��&�8���.�ў�,Ej�������bX�'}�]�Mı,KȌ^����I�Kı9�߶i7ı,N���8�L�g8�@[���Y��v8�"��F�uњN��G1���my���É����KE��2V�k��}��oq������}��Kı>�}�I��%�bw�צ�q,K����٤�KıM=�Y
�U�I-y���g8�����4��bX�'{�zi7ı,N�ޛ4��bX�'=�z�7�b�"�����������؝T����q3��b{ߵ�i7ı,Osޛ4��bX�'=�z�7ı,Os�٤�K�L��}�����-G)�_�&q3���{�f�q,K���]&�X�%��w�4��bX�������Mı,K��_���#��K,�&M&�X�%��g޺Mı,K�+���Ɠ�%�b{ߵ�i7ı,O{��4��bX�'���Y�~�,��d�2e��k�:��.ol�!B���rtXƻ�/\l�ZC��:x�u�9�.�n��
�x�M���ɍ�50��lx3p�u�/ D-�K�^1�EExq.G��wX�kP�;f��8�<�F���ݭ�c6��"9ь/iK8��琛Ǝ����(ʄG;�O6���e�rK����zې[��v��Z�!S���W������v���ݴ���3��K�kP�M@T�u��!�ӳv�u��5nKN�.-R,�iX���;�oq��Ns߶i7ı,N����n%�bX��}viwı,N{>��n%�b3���,��!%��m�g㉜L�;�k�I�~�&"X��{�٤�Kı;�?�]&�X�%��w�4��b���.�ў睱��-�����g�b{��٤�Kı9���I��%�b{���&�X�%���^�Mı,K���1����nf[qri7ı,N{>��n%�bX��}�I��%�bw����q,K����I��)�L��_��`�n��Z���ı,Os�٤�Kı;���I��%�b{��٤�Kı;���I���g8����D�DL
�]RKi�d���'VH����q��Vإň#�ڻ�n-p�)Tu�:�%Y���g8�ž���-ı,K���&�X�%��g޺Mı,K��i7ı,O��Ob���s�!.3t��bX�'��]�M��	��22(�H��	 &�4L��f%��gۺMı,K�w�4��bX�'}�z�7�*b%�����v���XYsqri7ı,O~���I��%�b{���&�X
�!����g޺Mı,K���_�&q3��_n�<�rYj�-$�3t��bX�'��l�n%�bX��}��Kı=����n%�`~��b'�k߮�q,K���X�?\S93I�9�ri7ı,N�=��n%�bX~c���_�'�,K������n%�bX��}�I��%�b~1�[����q��!#v��p;cv���5SCb���e�uI5R-��9*��;b+D��.st�D�,K��~�4��bX�'}�z�7ı,Os�٠�(O�b%�b{�~�Mı,K؝��~q..rK32ۋ�I��%�bw����pVı,Os�٤�Kı;���I��%�b{��٤�Lb�"X��}=ssf	3�rf��1��&�X�%��w�4��bX�'}���7ƋkK'D�(�P4AT�Ċ���Sg<l�E&�ϝ��B�c0�f&	 L�Dp�!2a	Z��h�lO�!\��ĉ2#��0CI��m2�\l
�D�¬P�8@\d�`0cA�%�V\ �M
�LPO�����	��}O���?T�:@�q:��L_�2�ѫ����L�� �{4+l��گ1��Q±�*��3"�P���|
�ϓ)�އf�D= �; �AH� �D�N{f�q,K��s�]&�S��L����9=-du�:�%Y���,��C=���4��bX�'�ǿl�n%�bX��}��Kı=��f�q,K��}��\�5��L���f�q,K����f�q,K�9���I��%�b{���&�X�%��{^����g8����H�\RXӕTG;j�N��K���k�̵���b*S�.�O&q3nq�兗%�M&�X�%��g޺Mı,K��i7ı,N����n%�bX���l�n%�bX��L�V8岨�Ik�/�8���/{�٤�?D�K߿k��n%�bX����I��%�bw����q,K�_{��P�q�j�Gm�g㉜L�;�k�I��%�b{�}�I��%�bw����q,K����Mı,S8�]T~^%�D�$����q3��,Ox�i7ı,N�>��n%�bX��}�I��%��FE � 3�
C��Z&��O~��Mı,K�I���\\�fe��M&�X�%��g��Mı,K��i7ı,N��٤�Kı=�٤�Kı?<�KOߜfK�Azz�n�g�y���wg�+U�Va�n��\�l�s��5l�RQs�������x�,O߽�f�q,K��}�Mı,K�;�Mı,K�Ͻt��g8���1�z+T��:�%Y���q,K���4��bX�'�w�4��bX�'=�z�7ı,O{�٤�Fq3��]�a��(�ÕT*�3����X�'�w�4��bX�'=�z�7ı,O{�٤�Kı;�k�I��%�b{ݾ7nq�兗%�M&�X�%��g޺Mı,K��i7ı,N����n%�`~O\���߾Y���g8�������rKeP%��9�Mı,K��i7ı,N����n%�bX���l�n%�bX��}��Kı8 ez�J�� �JUrDG
 H� �{�qCa��Y�d�S҉�&�a�R��-��9'5 �Ź��n�3��8��]��0s�p�����&]WvP��*��Kb@1��'o^�������)�n��
b��r�1�;me]ac6ƞ�GE*�3����m]���w�=���tlp�F����`�������v�ӷbNư�Q䗧cq[c��M�v��l�	��l򻎮]�"t�U���\��I\�F��E��$,![��x. l�\��8�-���1v]�`�K��v{V�I����U�-8���&q{��3��%�b{�}�I��%�bs����q,K����Mı,K�e��[QdM�ے����g8���-��7ı,N{=��n%�bX��}�I��%�bw�צ�q,K��$�s,�s&)�%�M&�X�%��g��Mı,K��i7��$1=���4��bX�'�ǿl�n%�bX����Z����K^q~8�����=��f�q,K��=�M&�X�%����&�X�%��g޺Mı,Fqym����K�T����q3��,N����n%�bX���l�n%�bX��}��Kı=��f�q,K8��և^�A�r��'Q-㜶3%֖�n�Cs�iE��,�x�f����<I:I��{z��n34��bX�'�w�4��bX�'=�z�7ı,O{�٠�Ϣb%�b{ߵ�i7ı,O߽�8�,�Xb\�4��bX�'=�z�7��,�5Z�@���,�<����&"X�k�l�n%�bX����Kı=�٤�Kı;��R�$�U��k�/�8���/{}�I��%�bw�צ�q,K����f�q,K���]&�X�%��Q�<�qګQ�eY���g?�I�O{��M&�X�%���~�Mı,K��}t��bX�'��l�n%�g8�о��Nڋ"
ے����g�b{�{��Kİ��G����I�Kı?w߶i7ı,N����l�g8������X�q��"u�-َ1�:"��h[��ͱ��C�X�U�HW\nԚ��%�Br�+�/�8���.�q,K��;�Mı,K���4��bX�'�g��Mı,K����`N�k�)%y���g8�ž�~4��bX�'{�zi7ı,N��}t��bX�'=�z�7ı,OϘ��V�k�Zg㉜L�g���Kı=�=��n%��7	�85Q;��wI��%�bs�׌��q3��L��}��u�|*`W)��Kı=�=��n%�bX��{��Kı=���I��%���������Kı?w߱7nq�兗&q���Kı9���I��%�a���|i>�bX�'��_��q,K����I��%�b}�=���3��wFLz��ɣ!�����vq�O���%��`K��u�'�#��f�9Znv.&�ǻ���ŉ����I��%�bw�צ�q,K����A����bX��}��K�L��Q�3߅$��(�v���q3�ı;�k�I��%�b{�{��Kı9���I��%�b{���&�	��&qwC�$s�RZ�ԭ�Jg�ı,O�3��I��%�bs�ﮓq,��;�Mı,K���4��bX�'�''��0��Hfaɜf�7ı,N{=��n%�bX��}�I��%�bw���&�X�'��F �#+ ��b�a �� �+���(gE0L�(<& � }Șɝ��Mı,Kg��B����UqI%y���g8���w��n%�bX�w���&�X�%��ﮓq,K���]&�X�%8��\J/k~O��eR���I�j1ε'���ldfņ�ܠ�yH��LL�FrR��1��>�bX�'��_��q,K����I��%�bs����]ı,K�﷤�Kı9�����ea��	3q���Kı=�=��n%�bX��}��Kı>罽&�X�%���^�MĂ�F� �'{�P�T��iM\, P��}8��"o��)�$��'y�zi7ı,Nu]��/�8���-��~R�d��R���n%�bX�s�ޓq,K��=�M&�X�%��ﮓq,KMLD��]&�X�%��I�O7x�ř��fs�&�X�%��{^�Mı,K�3�]&�X�%��g��Mı,K�{��n%�bX��X,RB(@�"D�Ç7;�S6fe����u�� ��Z�Rm�Ҽ�h�u��ҍ��s��J���6�ͫ�3zy��u.�A�x,a�;\v�ݱ9������\]�;��c<M)����l0�s�f��֑�t�х��;	lkn��&Gi��kH��K�������!�M��yBkr��n;L�)=�OFMp-n�u�!�GX-����r�ÎҷR�D�FN9t5ė�9�b���7QS�r;@v���v�ڞ+��p.�=Y\�j^�����{�!�I9�X�ԭ�JgN&q3��[�>��n%�bX��{��Kı>罳I��%�bw�צ�q,K��-kQ䬖!R�Umy���g8���g��Mı,K�{�4��bX�'y�zi7ı,Np�}t���"b&&ql���K�eU�$��㉜N%�����I��%�bw�צ�q,K����I��%�b}�k�I��#8����~�*�R�:�����q3���X&"w����Kı;�>�t��bX�'���4��bX�'���i7ı,O������V���7�Mı,K�3�]&�X�%��w^�Mı,K�{�4��bX�'y�zk����&q3��Uy�W]�jU��N!g9��׷Z�5�M,� Yn�������;��겼��q3��L��<i7ı,O��l�n%�bX����Kı9�=��n%�bX��u��+VJ�P%N�L��q3��L����M&��N
�C;�b%����M&�X�%��ﮓq,K�绯M&�X�%��d�'��L���ų8��n%�bX�罳I��%�bs�{��K�1;���4��bX�'7�?���q3��L��B�I9�,U�+e�ri7ı,Np�}t��bX�'=�zi7ı,O��zi7ı,N��٤�Kı>��t���̖d�st��bX�'=�zi7ı,O��zi7ı,N����n%�bX����7ı,O���=&���da����1����f��A�9�0��Gb���s�i��R"3�&�yjߏw�%�bX���~�Mı,K���4��bX�'8g��Mı,K��4�8���&qym���j�F�M�L��Kı;�k�I��%�bs�{��Kı9���I��%�b}�k�I��%�b}����沰�̈́͸��n%�bX����7ı,Nw���n%����ΰB��a��.. ���(�X������&�X�%���k��n%�bX��Ը�c�d�\��n�q,K?�;�o��n%�bX����4��bX�'���4��bX�'8g��Mı,K��I�kU�ژJ�r����g8���}�Mı,K��^�Mı,K�3�]&�X�%���^�Mı,K��I<*9�v�FEY�#����k;KWѫ�x}vL�e��5�v������ٜ��n%�bX�w���n%�bX����7ı,Nw����%�bX���~Y���g8��ޗ�s�X�j˜fi7ı,Np�}t����s1,N���4��bX�'}��4��bX�'���4���\T�K����~JIb(�eVל_�&q3��[�g�[�bX�'���i7ı,O��zi7ı,Np�}t��bX�';��g�*2ʫ�Ki�_�&q3��_w���7ı,O��zi7ı,Np�}t��bXw�$
eb0��AȂ@Ð��(2�'�~��J�q3��L������e���SvU���%�b}�k�I��%�bs�{��Kı9���I��%�b}�{fq~8���&q}���zF�W$N@�ě\]͐�S��Fvі�3���Vzz�f�ó��Z;+��(V �S8�L�g8��w�I��%�bs�צ�q,K�����&�X�%��{^�Mı,K���9���U��㉜L�g}���Kı>罳I��%�bw�צ�q,K����I��%�bw��<�j8KP�\�q~8���&q}�{f�q,K���צ�q,C1�3��I��%�bw����K�g��/Ē�TN2ڳ����&!P�������Mı,K�3��I��%�bs�צ�q,K��D�~��㉜L�g��$���*څc����bX�'8g��Mı,K��4��bX�'���i7ı,O��zi7ı,L����˥�z�@�H�S$H$D�iT�0���`b2a����$A#FF@���5���1"�c0��$H��,.�:C&�(AI2�p$qv��\JR�k<�3,��#$��$ �0}�SY''M�t.��� �)"H	�C8�J���"-dH%�LۓD:s(e�%	���dE��$@�!�Uk		#@$�I�b�!��"ý$��|3�!����+��9̴�,a-L��H� !$XD�#1#bHŁ0�^�;�.,�h�~2�� ��s!5�aD$�L�)P�D����(/)�Fn8���	܈t�b�6��@.����E��$���3�	�����AM��;����<9%�[�c���(s԰c,bXV���I؂u�UbօI�`��+�ō�m�R�\9Y.�m]5�%�D�:"v�۠�[j�*kd
��)5l�s�L�dL�V��.��5%�����b���L�� �VV��A
Sj��r�l������˄�\�J�rW��.�e��JgbI�vW+� �m�����J�U"����Z���ڇ8Pڪ��5�v�a��v��gG�x�%�e-[��5�@����ۅ�A���6{!%Hc���"&�lc�v�r�]���ݵ��v[�`�+� ͖��f��)����:m�$h���vStRoi�y�v�&W�[.�"s��B��t�t�[![
n�v�(�^�ڷkv^jδ�6��Ɛ��]A�6��۷a�,��)��A�Ӊ�룘�O]d�Ҍ�m��W�[Q�+NR���`]%t5T�b޺
�8�XP��Ȳ<n*�nx�H�m�f͛S�p�sj��NYw&�%:$����;Mh9L�:�t��<���+������c<Z2������%����Р.��g\uWn���瓔��{����+���� �kk�U���i��j��c��A5<+��ڱ��D8v3n��.�һu���jR׋��$h�8��ڞ�䑆�0[F���qK��S��ܚh�h�%�q�Ҁђ������秙���9Ɓx�i2�ݳZ��=t.Y\�%h%'Y��X��z��&�V]����V��c=����s[<����C�s�MC�(̤�h�k�LO8�iݕ Y��6/���`	;H����'>ɢ���m����ҡ=]CuvȮ�m�p�)	�#���Ȫ�T�-S$mڴƄ�Im؀��n^*�7d��0��-@V�X��*Z�Cfz
�[���[��0�m�f�ι-��l��Om:�V�i
��jU���6g�E�Wv��1n"s�).d�379�©�ȁ��>��(?"�~]=@CH�>Wj ��z��X%0��)A�|��_� �SC�m�yfsn3d&s�S��T�58-�Z�@�]�&"\��]�'N��b�2�s�l�imI�U���ؔ���ݗR{;[������JEkJ�:�^%]�]@�s;1�[�Z��s��t�d��Y6q��*Ll���&�ktt�rlb`�Z�����']�F{[<��f@XLpuH�z×�ObfMu���g7em�%� ���p�\]I��3sq1��/#�uÌ��okf�5�t�ngk\=��q>�C�e�:�%�:*�U���N&q8�'��zi7ı,O��l�n%�bX�w���~	�LD�,N�Ͽ]'㉜L�g�����j�����gı,K�{�4��bX�'���4��bX�'8g��Mı,K��5���g8����9=iTem:���&�X�%��{^�Mı,K�3�]&�X�Xb&"w���i7ı,Nw��Mı,K������p�a�q�fi7ı,Np�}t��bX�'=�zi7ı,O��l�n%�`bb'y��i7ı,Ns�j\b1ǲI.L�7I��%�bs�צ�q,K���~��}ı,Ow��M&�X�%��ﮓq,K��*�;=|Y{��`�\]m�8�����ix���\����d���mCsv�nS��q�q��X�%�����I��%�bw�צ�q,K����A�},K����I��%�bs������1����LY�fi7ı,N����nA�::*8���'�g��I��%�b{��zi7ı,O��l�n%�bS��=�G9�,U�J7e3����&q19�=��n%�bX��u��Kı>罳I��%�bw�צ�q,K�_mO@�!-��/*����q3��#9���I��%�bs���&�X�%��{^�Mı,K�3�]&�X�q3���/R�5FYUqIm3����'�����&�X�%��H����i>�bX�'zg߮�q,K�绯M&�8���'�-i��W���; X��\V�g���
Wi���qጽ��iq��x�n7
a�ڜ
�u7eY���g8�Ž�x��bX�'8g��Mı,K��}t��bX�'���i7ı,O���vp����S���w�|��n��;��0��Q�p�ڀLuY^I>�9۩&��{5;�&%��\�ήs��﯌����]�T�G%�0�SuW8�B��ߖǷ� ���p�;� ��ƃy�;]Q5,v��uA�6���7���&�t�;n�Ȣ��������YPx�;s��9ӫZ����e�/���IayS=Z��}���gK`ogK`M���nY*�C���Y^�gu��.6{��X��� ߔ��VҺ�+vU\RJ��7���(0&�t��t����&�S�[N�$� �ݺ`�ש'��;u �:0�9TW@�;���v�(��',��)�x�t�ގ����ud�ɈAY��rGN���M�[\��e:�m�v�;�̽�h�T���*��(UG!Ò�c����;� ����(0&�t�ur�Y�Yy�XZ�Y��z:`v��Ζ��gu�l��cA�<�����;V��� |U�8l�v���{� �
e*��,YJX��Ζ�ٝ-�7�,=���c<����������z:`v��Ζ�ꯪW�v���ڽv�b�U�ƅMm�λv�!��<�ق��0�t�vŧXݳ���[��q�Xe걺�ݶ��������ЉQƝq��!��uR:B�K�v��L�Um����n��1n��嶒:a�x��(�<��X�r�[�pn���s�[Hu��)�hݦ�y�;]��#���:�fX�ә�#�I�u띠D�	������Y�gGmڶՅ,����{��<��v�7����6�tŭC΍�ag����nL�`��mkc������t<�������k:[ft�]��&�S�[N�$� ��t�7�:� 㮹�:�g�L�ݳjɺ���1x|���Փ��6d������(07���-@1�ex�7^����(0&�t�uu�YwYy�XZ�X��&�t��	��-��7^�{�Ӫҫh��eP�Tt�d����퓰֙zL6���v:�n�p�v������;W�7}|`�׀}�u��w��is�e���Ge0'~1��|*iC! ��(�@���Ū<~  �ɩ���ޑ��(0=�d���ىQH��us�q�\��x��IL���oT�<��TJ�eU�$���w�k:[{$�����"J�(EժY����k:[{$���ŀ���[��U6D�[��k�l�۫tsVz�(7�Cq:�]^�lΞ�����%o]�����^#�M�P`od�������� ߦ�c���c��`vIl	���ފ	��	��%���K*cuZ���L����C��J`��P��N$*�-�0�w� ��X�S2:�jX��A�6�A���-�7��[�Ee����)�o˷L�ۺ���ފT�+2��Yxe��V[SZj۴a����
7=v..a^�chKA �N�T�JIb/*v�ݛ� ߺ��ފV��t�^U�+����fbV�����]��RձA���(�z�}���"�I%X�t�=[�%�7z:`l���Y��]���^!�����%�;z:a���D( ��V�����U�
KX�[{$�oGL���^Ɍ���m��iʜ��,�F2�mM۵���~�䳛\�%�v:�S��g�����쥉_�07��ײ%���Xt���;�m����Z��9L�v�z�D�����A��eL�̅,J��!]�C�:,`ogK`N��ۦ�����I,�Z� ���������&����v�R���J������&ݝ׀w��>Gk�-m�	��i��	�X]bg e�h$	&����.�v����j67����┴�P`�촜g��%쾍Vʜ��.��6��l7n����:��+r�3�4�h�_R�z+k�dkC�<5�H����ޑ�q�/hl;K�g��K���=mE=x�@�e��4d�p�\&Vr�f� �jr�B�l�lt�c��y[`����u%D�����;2�p��e��w��#\��a`vz@�!��64(��Ub5�3u[#+i�d����� ���n�gu�s��{}|`o�����Ɵ,��`od����A�����������,G-��-�\�=�ouA���LL�j��3�Yk2Ē�tP`oE��$���Y��UMK���� �כ3�����`Jl┗:���v�÷f��g�gps#��[�t�:���0r� c�����i��������R�ݒ[�(06Eޒ���Z*-�L��וu.s��ĸ������ ܽ��jI��=��}�s�\�I6wb�=`�+���rZ��{�(3�w{"L��l��w�+j:؝VIV�{�� ��޷ �gu���,��{(��q��G)�z�D�����t���UUoRK����]�4�Nhu�Ю#ţcU]��iTQ�$ݥ�n9�g��gm���i%�$����:`zE�dI����l|�[*��Ymx{�� ��`����;���7N�%[��f*�jX�X�ۦ��^b��T3�lŦ&S�#a�+���T8
�+Gi!X"Č�!|*1�g�l�`�"FJ��0l��74���&+(`H�!��d��;&�u�!'@���$�0_�<D�pm��(��VBC�@ٲ	M��t
gTD&�@";:	�Dڅ��Nl^/(�0t���S����� Tx�5
D$��]�K�����>�� �
]�I���[T��L��v���׀w�t�?n�0�Ƨ��$�j�ڭ�ݝ-���A��+`z�!�_�$�Gi%cAs�{'azÑ�yh��l0��-�le����".���t���A��+�U�	2~��km�Ҷ����l�`�n��q���z�vo���� ��[�ݜn4�X|����0'gK`wEء�~XpP��B������v���05%0ДJ�H��$�!F�<��P�a���u$���_R�9]�B�e����,��8��g��}�_W�ogu��ݑ�-��K.;&v��஻�m!nŮ���R��笸�m���,�"f@��&����w����`NΖ���t�3켅,J�f(��0�M�g�L�������?n�3ɳ����܄�T+S-������a�<ݽ0뽙�9�R�jD�u�\NK^��� ��t�>��o �gu���ޫk+N^7U�U�zE��[�:[�GL���PFAj�+B�m��J$A*�����g���sn-snm:��ʳ�(�b��6�#��l <j޷��M�f�ې�F�m���u/n{4�ix�&�d��ݎ���;j7q�z�i:Fv8���;2�o�;s�0��G�징γmZ5�p��hC188|����g�V�;X����.h�B�f�y]������6:��T��Ev�Эխ�����W�2���>�w绽�����s�d�t[��-i�BMq���0t�4]Uٷp�v�#�I��]_�
E�8	s���Ζ������ ��7��o ���0�t�oGLH����`n�*,����QJ��׀w��,��� ��v���׀}����2�H�-���<��0ݽ��;����ŀs�.�I�Z�|��L�m���w^����(0'�}mP�2�0ˡVm=��fl���g;[m3����R��w챎S��H�O��r��b��^����;�w�v�JD} ���8])�Ju+���WV���p�r!.BQȈ\Q�[w� ��ݷ �gu���ޫk+N^7~K0="�^ȓ�:[��� ���K8�,����}�p�?[����(0;z��|V%�%i$��Ζ��tt���-�/dW >���lQ$V��E
�6�a���Ƅ�v9��.��mx�[��k�-դz��긬U�$������$�_tI�ݝ� ��je�)*�vڰ�7^y%
d췷xt�p>�Y�2uv�1N/Z�|��^����{;���a�J�B�M�xϴjI�c޺�n�u��Aʪ��-��{�|����f��>�wl�>�[��e��b�X��7�:`zd���΋���K��{�kNOA	�c�UP�����
j��ї��{a�MuإƇ:ͳq�	�l��
��U��=�}��ـw�����ŀ~ݦ�eO�
r�RJ��7n�bdn�� ����5D��j͢#�-����vo�߻���7^߶�x�M��9]�)T���5(�׿,�[��w���)�Dc"�Hq>�\HI,��<�`]P��#*�I%LL���El��lw�� 5w�ie���qW�I/)-�U�`����'V�u��۵�틷�����|�Bĩ]���+`M�+`wgK`v�t���u��M`��r��b��^�Ζ�����[�(����0ʹV5IS��e� ���X훯qq&���� ݛ�wf���aZ�T����%�;rd�vt���䟽L��?X�Br4+I+�:�ٷ �M������>t���aD)Q
�	 �F�J
DP�"D��J��*��JB6�ל<���4�B���j�*���p�p���;���q�;p����F�=K��nh(7��%���V�ۜ��b"�K���Vܫ��$1.S1��S+��ݻ�tɷ2��N36�۶�i�ۧ(�9����X�M#�i6-�Y�� �nBB����=yf��keg��d써����[���Y��d�����zZ�PH��ݳW���Asη�F��6.I���l2���^5�U/<�Y��*���KR),�@���s�w�x��7>Q���l��u[U�I,��am���wy.q6}��<{�� �gu���ꄅr��*IS�$�NP`wgK`t�避�sEe���[��n���������$���W���Ā�����;���:tt���-��:[ ���?��@�ZM����g�	驈5pq�!l3��ٜ��ۘ
��Y��[�f�UbI[�GLL��9A�ݝ-���oamei��T��`�n��{��.�
���)���7k\�}x�R�}�Q�����X*I^���}��l�0=�%�=:�˺>+�*�bC{:[gGLvIl?}Us�?��k�ξI%�4�%������>�78x�;]s�j��$�N^�)��۔����#���g[-{�d�Za�<�����en����W9`n�uUߌ3��`v��t�W�6EHmd�sEe���[��}:P?}>��?ww��u��MO�9h	�� ���n��w�ѩ�[a4�\}�k�@~n���T��(RU\��k�>�0=�%�:�La����~�L�w�k+M�:�,� �ٺ�s�ql�<L������]�r�#1R�,���6��I^���(�t���HV{V��ơ�C���=+��X�i�Ь$� ��v`vwm�;���$���L2��Ī�����Ζ�����$������6wu��_$�ڢ��l� ��ذ�Il	{&06gK`zQ�b��b��UHKmX~�� ����>��x<��\縸�����z1G<+-U�B�V���cft��%�:�~�_�֛��rm�R\�)`�C����F���+ZS���5^�Yѷ]�nk����8�pw��Ss����8�u�~<�G��IUr�m� �{t�;rK`zd��ٝ-��%�ŉ`���֫����A���-���L�v��n��hV
�W�~ݺ`���ܠ��d����;��>+�*ʴ���Ζ����$��]��|m)���ޥM��VCP�¶��>V��"A�ѝ�&��3	�"sd
}� �����O�h��"4ۧ^�cBմ���Ƃ!Q9�}�v�6��ѸPu�����#i�C[�QqvF`����$`ȱb�	11�&L\�T���Y<$�b�b�U~R�!"�>5��f �0�ȠI�lP4���'��mșp� $R D��H@��ZJ��,V+(�D	�y}�.}�k��8�}?Zڤ���T=�Җ�nm��m����cp���+=�o�I����˞ݭ�B˸T�sŁ|V�l�R�8�	��WSV�K��!��F6��	u^�Bֵk) 狵Z�Z�`��@�wh��^�L�$s��C�C��*�[��HZhy �VP�(KʰY�LQ��2�]�%�A{+XCyQ1Y��m�o(�]�ŃFr�v�q���c�m|=�d�A��l�W'��E(Y�J�[T��m�h��mOi�>ܵ����m�A���eue���7TI�x���'�Kݱv�I�i���`c,d^���pQ;�l���Ķ�F�fM�3'&���ƧT��gE	.���أ��pS�li��ݡ�f5���	n�4��[)ٮ�Zۄ��Ȩ �G�w���'���:�=[!p!P�n w<&��ĵ�Y���V��ζ��X�fCX��l�ɶ�Pc�\��S�D��V��0&@���-�"4*�m@�N�t��;ӝd4���h��ƧW��n6+[M�X�`܆�^�+���&ʷ�����;DX����aUCPp�Fج�+��`a���l�J�ۚ�ݫ��sM�ۇm���{3�\㇁�)wk{;�e\�����ϳ�m��(��J��8�dɾ�#6g�|貆ݭ���@��ݝ�@����VA���6���b�4��vY���6R���By�pQ�{Yݙӝ�]�v�[�>p5t�=N�.�H:�)G]c���۬�m�Fzܩvn�1c����p-7J��h���]�p.:���$e���3XƦ�^m��E���iP����yʄ�\kE�.6��;�q,&6<[��蝡���><v��9+���'��.��Wu�q����;�5P�UO�8��Ɩ|�����4��t<�:���ܨm�'���pi��"k�v��m]wX~>~{����jlA�$��΅CHlMJ�?"�?rr�m4�t��ֱ�n����3�#����¨��XpQ�1 �6��GO�?  �}�����j�t����~�8y1�rV�.��V2<��4�-�m/hh�N)�km���i�xa";l)��B����;��v�ܱ;]m�:�&�Е���o&���u'3�#�08�8C����m��]9]���-���	��t�2\��1OGj�g�kۀ��C��Ԩclu�מT������š��(�9�]�l��+��4�5��Ԏ7ij�vP���;��Ӳ��ũ�^���w������[��k��Mn B���M���~K���#�2\�v:�����&#��s���m�?����vIlؠ��Ζ���R��K1b��Ib���A���-��ۦs��wOeT��[R�k�7��ၽ�-�����0*Y�`V$e�07���6r�ݒ[�m� ���{�J�Uʭ���� �	q����n���\�|r�R�$��ōs)��=u�5�:^�i�;�"��s0�Ժ;�ͪ�vIlܒ����9A���q�u��Ь$� ��u縓_#�L"�"�R*��� hĝ�}�����>�79�DL�U@!RUE����:d�l�����-��7^��i��I-�D:������ ����v��Jz���c��J��eR�L�M׀~{�0�w^���}ػ��AUȬn��{v&��C��lٵ�vm�%f�f^�l[���Tg9�%���n׀~ٺ��7^����q~a�=�wӞg-�>IE,� ��6"P�Mn������6!q$��E�Fy*�W*���n�I�c���8Q�|X@�G���>��}�� ��z�B�\�$���;�K`tΖ��9A���Ș�C��X*I^ݝ׀}ݺ`��0�7^߸u�,�ʢ�A�Nv��y�JE������e��:���a
��sC�%�VY^�v�w{t�>��xvw^���l|��j�*vʰ�����-�Ӕ�A��K(Z�%�YT��S ��u���0��0�n����d��[R�k��Q����0��0>J!C%�A���A9��"��ݺ�?}!�
��$�KL{�L�mс;$��(0=S.��H����#0Q�r��૏Q��㫍V4mN�SnR�m�%Q:��J����`}ۦ��� �gu�ݺ`�׮Yd+RK�%�ݘ�79�D�ݧ��k�� �� ��f�݈q�+I+�>{ݘ�a�DL���k���:�/&�"��,��,`N�ؠ���[o{� ��u폑�ڨZ���~ۦ �M� q�� ���!$��ͫ�7]�zݣ��:�g>�.S�4v�÷a�3���B�;�����\m'J��V[(��R6�h�%Vm��I��B,�Ν$��K�ށ��g�����x6u��GN&��[p���5ʕ[�[[�nبAz8�D���ջK���2���7f�
\����l�#l�������)M`�d��>s���V�%�o^ݙ�j,�FN9t}���w��{��r_K�Χ�)պ)�M��Þ����W�����<I�]������������7o�2�MìX��3�?��9A�:(0;b�}��d��[R�k�>��3�I&�=�X�ޘ79�2;:Q�U��3�����Lؠ���[g(`�^��"��+��ʰ��L{������S�w�7[;5wuH�Y���Yi�%�6r��GL�n�����m
���I����-ݝɦbh��Y�Yf�sM�[����\���XR3�6r�t���A���� ���KR,v��n��Ī��'%�$��P`N�ԭ�5e��Ki�w�`ٺ��I��o���� ߖ��q�ij�$0'd����tP`l�	���H+e��+v���ŀ{�Ik���;�z`�����*g,	�ZK�'h��)��ںR��d�����-��e�::���W�R���Z���{�L���7:�/��ŀf�ԋ��_*�_$����K`wtt��ۦ��׮YdErJ�%�� ��۩'9�����T��#�s�w��}����8����hV
�W�w���]� �o=�ݜu��d8rZ��W*�;ݺ`�w��׀w��Xݏ�����`T1�iN���x�R[�9��i��լxQ��z��Y{Xmo��-P,R[L����>ٺ����B����� z�������whSuuk ��5D)�������>oq`ޅ��$��[��^��q`���GL	�%�=W��*UbjJ6�XI�}�0��ŀof��A��!�H.F��.�{�RI�poC�����嶘ۻ� ��׀w�����0��ZqCX������!��Rz�޸x�9�/6ٻ��RNqK����v���[�J�%�U�of��;��X�n�ۻ� ��O]#hV
�+`wH�:(06H�;$������k�;#||��b,�`�_ۻ��I�l����ŀoz;��GIj�b��� ��� }�� �z�`yDBS��� ���'%qKP��j�7�u��0'E���^e}�����H�n��\�Gq�h$	3�4x-Iˌ;s�:�r�t����nɛlvO=*�$�!��[����N�n�\�t�v7��v{���^�R'�f˶-���' FC�99��=][�V.����z�l[�1qG�f����M�v��-�'|���=�F�*ɵt:�DÊܲ�NѫX�8]]rv.$�S[��͵�:q��26k��������#��MN�+����u�adGl�^y;[:��ڢv1l�%�nMwV�q��L�~������:(0=$t���[�m˲�V!U�b.�0'E����K`w��X�uR,�^W/-�`�wvIl�A��λ��,�`�Č�T���[����P`{wq`����Ѳ6�`�%x{��`N����rK`eO����f.y��k����ӵ�	%��.�a�n���`���EF�uH�-vF��-��Y*��h��w:`{������P��1e�-�\c7RM��ѭ�������Φ��7������K���m�|��C��X�S�g������;:[�w�t7*	 ��*ܭ����� }���>m��Ԕ)������/%)SRQ�*�7���ۻ� ߦ��;��, սڤ�$��6rV�n�Ӳ:��\���u���[��6^�u۝�}O]��b�W�嘭��#��Iln��ӭ��W$�R�9V�Ζ����ײc�GL	ܮ�tl��Xr�^��q`n�>����ӄ���$X0`ňH0"E�R�H"K
LJJĤ	�D��+�zٕ�N|���[�P�0`$H`� 0�&s�d$:�Nf�]�����1"F1�d�&�P���SID6���A:��d�a�$��)��9�tںUw!MBP��90��/x��0!	�VL��Hm	H�� ��7����A����PS !�'D��H����~6U(;W�Op�a4���C��D�I�~�?(S,$�7�[j@�$U8	��r�"� �T%X1D� �I$"��$����CbBڻE߸h�i��U�#�PO��i>4C  ��_���#L�u�&͂Q���E��^=U0A�� Ђ�:��{�RN}���I���;#||��L�������z`ｋ �����Iq>��� ����%-�
�fZX�ݑ�vt��P`Kٳ ���5�J����'B*�����&軵��Z�ƌ�׵�v-��nc��⌴�j,��{;� ��`�ݞ\�\�ý��`���$��-U�[���A�/d�쎘����vw��*|��v��}�}��,{�ŀ}��0��=�Wd�+���0q�X�^,�v�P�3	J%�����i1�(Ҵ
���P�E0T�)��������v`{����
않ZG*�'tt�݊	{&07dt���W�]���Ѳ�m��ŕ�:�%�*�je�-�Dk�g@��PܡˬX�2�h�d;qz�v���� s�� �Ű�}!��,���;#lB��L���5��3�q%'{�� ����f �����UX���Te���0'tt���n�~��wY$��P�e�`{�Ju��`�z`x�`�x�7%�L�V��V�vՀ}��`�ݘ~�tjI�s�5$ڦăXxJ�<�����-�^������Ifƃ�@���5 �g�W R�]Vu�[�V���n�euwP旚�m��w`Gg�tC��v��뱷Nb�ԚqͶ膷l���u�Hj�bl�8�.w1�6������$����[�m�܉=/��������t�O�\Bm2���>@umw:X�6u�n�P����ڳ��������2�Ó@�c���Q�%�J������]�:�w��{�N|�Is�,SZ[��u�#�%���&շk"PGe5��u���وH`z����l���:`l� �uR�Y*
��r��n��7�x�>�0<n��
&N�ڝ���wD���G*�=��X�ۦ��ـw��Xڻc��6FН�� �{t`K�1��#����̲�+��ZC^Ɍt���:`ov�w�6�h%��(����-u[����F�xw����w6��m�����v��t�y���K<�ߝ0'tt�����f���d��mM��*�7���T>�`�O
���Lg��jI��z`��� �u�jd�V�nWmX�(0%���H�;��[�u�ʥj���$0%����wF���L �uR�Y*
��r��o �׋ �� s�� �Q+{��1)s���W��'͡���r�j�iz̎IyÇ�Gm��;TWE�����?I��g(0%����q�6�9��(�X�ۦ��ـw��X��� ߵn;#gQc����;��`}
)	�� ����5�t
�p_��{F������>��m���KP�j;f߷q`�06r�^Ɍ	�>�,�1	eL��ݬ������O����`ww���j�$Q�P�I*��
���ڔl�ݛs�J嵶ź�9Q��Ŕ��ZJ�ܠ���c�#���� �u�=J��$�KL_۱���wGL�P`�.#물T
�}w��0'tt�����f��j�)+�7*�7��Z�}�g�RN߻�jNQ�T,,/��9�)�{�~�lp�"r1	�Q�L�P`K�1���wGL����y_�KG��*�b��ȯ(S���s��;-#�d�bZ�[�z�G�W��O�Z.�������[ŀ>���P����� ��G�_#㖡4�v��wq`�x�s�����Q
&M�r#pr���;mX�}� ���0n��۸���v�G9l�V�vՀn�^Ɍl���:`u՗*���e�06�L`{dt�ݑ��}�3٩&�Q� F�0��.5Z�u�Ҽ3�������(��ؒ	Yv)�=��;wt��6)`���vz�8�ʬM�Qѐ�[=�-���q�NW�=��lkl�:���crY+d��Yp���m0<϶NuΈ�m���-�]i�mO;�e�^g����K��)\��uŷ/��)�[��=0����<�����,�l�"YDfQ�-��%a�p=,ҏ���������~{���Q��Ƚ�gFמ��;���N�v�9�:}5��ѳY]���q��l���ݴ7��w~t�ݑ�w�{&06DI�Y	+�7*�>�w�ݺ`{&0=�:`N9e��y�j�ISw�{&0=�:`N�遽Ұ�&�՜E%���ـ}��,{�ŀ}��`�u=��>9jMWl�;dt����g(0%���}��N�����w8Ӛ�����Ύ�җl��#�*iz=o7Ro��|]�.�7g�1jx6.�� ��`�m��7^�	/�8�q`��}X���X�r�j�>�n��%!)DtsZdeJ�2�5L"�C��%����'}��ԓ����??���]`��%���ـ{�t������}+">�����}��0=$t�������l�>ݦ�e��IX���L{�ŀ{�A�/d����a����� �(�nV�v�����u�U�m�5��ke����'!!#�����Հ~�n����P`N��{�3U��K>i!�/�����:`{��~��m����P�j�f���`N�ѩ�ψ šQP( D �"D � �"�m�y�}0�b5c��[aib�:`v�\�N���e����[��V߻t�5�v��^,��X�$��tUT��An
�\\���TL�n,�8z�S6��N�&ݤ� ���ePU��2Z~���H����%\�ˬ�AJ�رc���I0;yA��7^��6�,V�%b���X��nt��%�=::`I֯2�2���_!b�nt��%�=::axA�"FXpF��*����*��WP�Ͻ�RM��51bj��׀u���?ow�o�W\��-�P��UU�ɧg�] �v���C�rs����>:[)y���F[$V����M��g�>����ŀw��~_�k��0��j�������u��5$�S#�=������ŀwu�s��nW-X~�׀$LN��$t�48��a/,*�n���
v�v�k�Xm��?vw^��SԈI(*ܼ�Y�~�w;	%������ �;��<�(��_�"(*��_�DPUj"���_�����AU� ����,
�*"*T��DH
�R���E`�@H
�Q��EH
�@"*P *
�Q��A�
�EX
�P *"��
�H�� *��@��F"� *��F�
�0��B� *��@B�R�P��@E��D",H
�`*�2�b*Q��D@�"�B�"�� *b����"**��Q_�PU�"���EW�_�EW�(*��AU���
��PU�"���A_�_�1AY&SY)9��HY�pP��3'� ao� Ϻ�:�#-6���   ��@�@ �` 5� )�a���5�e $  ��O���h	(   h  h   ��� P�
 @2��h��C@    
�'      �
   �������á�9�z\}z<;>�s ���{� ���f�`}�{��=�d��
h���ڟG�� Z���A���^v�a��A�}��r��  � �@�   �������{�@w`�7����]n>=]�(q�� ��;���p+�ςV�E�=�{���ٞO���=�@d� �}➷6�>��w�{�>�p u�ր�  ��t���;� |]��u���6��y��O�6S�=�������f�O����|A�����t����}�}�}�O;>����p������0:d  �� �    �8�@��>���<�z�s�/�/�6�z �� ;�� <�)�{� �2��)�Kw��
z^gJ zi{۞�Q��:S���W��g���{��җ;�
u�Ҟ��)N���ց��)��tzt��zz<�Jz)u�  w   @ �76��h砥�sѦ���P g��}� ���\n�.�C� hR�1}
��>  #�}���[��(�ww �a�}�p=;�c�zd��������>���"~�Jm�JT @��R�'�U  fU%3j�F  ��M�*Pd ѡ����(e)P  ԩ2�����������������}>�_|?aϿ�DW�֯�]�"�� *�����tDV�"��������8�f���)�m��2�����.�O�w��uxV��WZ(K��eC30�IbU�4 0"ĥ����'31�WS0��*@�	
�+*J�Ć0�+
�1������B�L�s��2�O�´�o�)��O6+/�����.d�i
BI�`BH0�ĄFW!L'Ґ�!1%!X��b��$b�!XVP�a�`q<= ��|��! �����l�)$*Bb�RB{�3Z	p�ީ�'6B�)+$�!,%�$8K! K\��cbK�]��Y	)d.��0�Vv��M3S��M�-�ӑ��S{�#�.��W�x�\u��)%��Ř�J�Mp��>[��s�#���8�$ԼB����f�|ݹ���"�R �#MƄ/��棣#5�:6���HF�T9�~��؛bae$0� �� bM�c��Wэ�M�.j\<���0���zܸl)
F��J��%��r��J�v�H7� )y�No M�p�����RT�&�ju8��OM:|-�����
iu5��7��75�IH@��TcB�0!\\� �(\&f�{�N��]1&k{�M���Diֆ�3GՖ�N./���Ž�U>MZ��طYvj�ֱ!BHI(A$H�!�d
A�(E�$��0�]$p�a�B���!Β]�Y
r�Y�.�rK�\�<�H�.8�;8�X�ù���%������+
C95�w�J�i�&D���*0Rn|��٥
zz0�:�\2�S	�$��2\�BKs�Bs[�3{8O5/6�v�����w0�!45tE8/
IS'g;��Is����#Q��5�7��..�K�.����R�Y�#  B�3YL�lѩM�p:Hu�&夗&.�.i��߄����F��NT0b�e��.2�K��²��+.�Y�S.l�4@�3�7^xS"20��I0a4B䒲���nBLH�%f9�.8,��X�Q�,�IcAf]S3sz&��><p�V�H[9���9ɬ�.z��!�J���HD����2�H������`F1���e�b��B3$ą��7��N �$��X1(�B�K��-���{�_}_Lώ���}]���i��Z�o��\�4����J�q�cH0%��X%%��a_��d*`L��эXLaq!XЉ��sA.ie�zAӳ�}�s�4K桉�����_X���2�$��m ]�h6*f�Hv������.0��*�.ͳy�6F������D�&$�Lae��I,V5�	4�<H�F!OhP�T�!BRH�ǁ�D$�00���!H@ ����8�T!v�K���~y��:!qcL!r%$aa$�@�
iĤhdlK!�$� ��0�A���������K��x8q�0#bT�U�B6a��p����޶I�!�M��O	Yv��^x���!c��B��H�IHP�"�7DjE8�d
� �B8&���ķ$4���1�r}���P3kʲ2�#,�B����ɩ���Qa
f��#FM��D0HU$��B#X���M��h���᱔�5Yn$��j�e0��¤�kM>�1."�����x�e�{��Us�WpK�5�W�
s�H���P|;�.yVJrڐ�����;t�2��d�aC���8M���pѲ�B2��a�HP����>����KM:^0�� ��)	
F��R�F� J��B��cƄlK$�g�y���.m�jSz��,��.%�p.`g!V0|{����(B�@�)J|���2c���T�$-i��I��iZ�;���Re�˦���6p���	tB�B� SX���YRc�0%��[�������<%����7�bc2�[������4����o���钢];Z�	gȷ�HE��h%߇�gZ��>�4B�SS	P Y �]:.�������1�B!�q,�ԦOf�k��sd��`A#1��X���iojYe��.��Ԅd	��M9�ILfg&�g��\�a�S	���*@�00O �r!�!
�)
z*c�\XW��n�����/8ā',�/	s���1H��� Ƃ�1I��9�y������K�N����� ��1���R54���)1#���LbG�0Ӭ�K��x����1����K��4�u�e̎$��\���=�:0�%����;7{��C�>����BQ�4l#q%P�0&2臾��#�����D�bE�"0�1`�%ֽ�����ϼ�Ρ 2�bؑ r��g���kid� pD+���@!
�$ �A��\`\�B��X�~��A���ಲ�H�9�}���Y�0��Cz�p�ʟ��f�1���$�����f��HX#ra!�!XP�H��1�6lލr���^y(K.2�nsis[	*�F�,X$HE�F�,�3170�1�)�x��Dֈ����r�)��Ze�F�L4n7�cLHP�q�L]��u�>n���2�{!f2�-�S�ĕ%��K���fUf&��U������Y��
�T'���[����I��%��vh�۲�D0��1&��D�4�0I�`�i��C��S�A6n�RX��>f��w&/�f�ԛ�%�d�C/�[��s���2�_fm�&�r����H�S��$b�E
�d��y�n\�:G���,�H2I ��aMI��y����>�6z{3F&0�̳
P�V�c)����c��
D�+	���d2�$�h80&��3MB@�ub�[N�D��*���S[�a&�P������R�,�	4���o��)�>�g����u�ӹYeԼ�BB���x@�+
B�2�*ċ�0��u�G���D�����M�M�7�i��e=�A���(���.�sPœc� ũ
4˭{
��
&1l�d	<a�&�a�A��,$�e��ef��z�\w�Q	4�1�,(4s�����۾Ϸ\[Mۦ�Ms�t�ՌRBV GA��B�p��)MBA������N���.�+>N�xw|%��^2�ٲ�Ƅ����qվt{��"#`D��!�i��		I$ (� `��*��$�.�Jc.H]fg�]|0�bD�L���4��p��c<�z�G�Qr2-��S�K�%.�9�����F���%܌2�m95_ߋ���Ms�~y�<���8G�2n<���w���Ev�.��M����O���5��q�E��L4o��E�$!!�%%�t�����ɖMt�� @�,���#e6F��]�SAZ��)����
�����u���r�~s#����q;468w�����m��.�a���	K;���f�J�:h!*e��#Nf��ZAh�"dH&�B�M�o�d.�4(�w
p/.a&3!��.R[�����0�+1 @�-,�jpٞ�Z���+��.����&�Ҍ��p��b,F����f��RR[��B�ZJ�����Z�u�\��;��%cYX��cF�o��h�'H��i,�CK��?g~g�:���f�$�Ѓ	y�p�>M�<O�S�0�4`Y4`0H2�!v4iB�.Cb��0�$)�� cB)��2�R@��J�d��O8,I�"�$"�ĉT�z�!�T���-$$�šC&2�y�a7�S#B#H$�����Y��bϤ�0�JaѦ�\
{e��7��d���&�s~��%�=�W����L��|�8=CB���$�' 
�{8rT	y�.�v����K�!-�
FH�_����|¸�
��H���Bİ(@�+"
HD�M$REX�"A �!���=�Bfg���oe�!� 4��(țP R1 5c �cB&�����g�9ᤞ���Ab����I
�f+�����ks�_$X0=$�uL=7����̆\��T 0X4�k���@li�, ���B$GC�f����D�hp�$�(�)
�!���Y	4^���D�	�7����$b��BR� ~�	!�� ��\�@�j��	BP#H� NkV{�6OHI0d#���3�߾�j $IX��4��@�D$N>���p6\�ٚX�܄
��@"0"D�!�㙒P���"J�"0�����HD�i�Ō���(Jʕ���4�!�F����їq��!�)�t/�n3�=�.K��%[��q�_o�\wq�?}c��{��Y@�$Y��6xr�k�q�M6�^I�����ZB�HH,54
���ԅ��=�AA�a@�/wΌ�ׯwY:�׼�����*��UUU_�w��UBl��UUUUUUZ��UQ���*��U]4�Vʠ�UF��U�[j����SU�[v�*��U',��*ʴ�5T,UuUUm�碆������ڲ�xy�G0V�
`.�V������ڪ���V�;t��ʵ�T�N�;s�U*�P�UC��G@*l�Y-�6�][5�DVŪe%ڪ^Z��������U:( *��j�����Wn�*������UV6�M�炠�{�}����ٮU��a2��UPV ���UC#t���UP�U^�
��  ҆�]uT+S���v�`7�胐��2�(`SR�l������hCe�vH �T���*�ҭS���쵷*��U
��V6M�����`%e��)MMU_}�@�8>�Q�M��sj������W`*�`8�Z��������e%8

�uUu*�J����*�Jʠ@R���;,R���Wl��-�*mb�jeZ��tZ3˵j�&��U�
����������
�u.� ��R����h*V������5��SIW��N"�
�r$�~w��n�QY�ڕlFƎ[��i��7cB"\ftl���@*@)�&��R���K�����o.�p�fS8X
�%P(�������[�{��[����$�vj(�ٕ���-�ڪ��U �q��iUƶkj�u��#DUT��U*�[*��T8�j����mTᣚ�]Ms�۴ �VԱl��Bz몪�%�-�m�����v*�-�D���ܒ�U!=8��y0�Ͱm]cR誥C���d.j���j��������UU�UV�u�UUJ�UUUUUUmUU�RC���Z��@j����U���j����e`v�4��遗b�
��%y��m�������W�Z�b��f�������ej�ȡ�R��Tjkj���ZWf�ꀺ��UPR�UUVԫQ�QH�v�*�UuUV�U*��2����x���V�7][UUU�ec���JPVX�	����@Z����)YYV�����}��-PU�T���V�Q,�ԫUJ�r��UUUUUUJ���X���@UV�@U�N�qL�z�`6��
����US�*�U����V�����*�YZ�����Wj�����
�����r�`ܬ�ʎZڨ*j8 ��%v�cVҮ�0n���G�{�n�.�j���*Z��UT�J�R�4 PUUUt�e�;5uUJ�*� ��U�UX�� �����r�UmJ��T��*�[U�̠l�gK�T���,�;TJU�T*ں�Y�^��.ͥ�e���'j��[T���UTQQ��t�Q������+}��ꂈ�j�����6��v�UK���؍!Q���WO;/�ћ�u��YP9�V)�v��cJF��2���MZ��Ђ^n��]��m7�d�@�[&]�r�wmsVԂ���`�������솹�&��Y�qr�Ub� ,��dAX���Z�m[���U�t�c]�0U�Q����l�UUUJ�0R�������P��ɷ@5U@E�\��u��%J�R��@AK:���y�ܣ��N����c
N�h��������+m�WZ���3\ RշUU�ȷJK���+���h͛h��F�Z��:�����u����Q��3G�xc�S�U\�R����Gn����S����)nT)�Z�m��sШ�k+U���8�%d�r-��ܗ�z��nV����8���Ak���Ǫ:�4���d0�t���6�Nv���b��k�Wtt@ )����k������q�K�LU@sn�.�/=6 *��Y	�VX B����rj��r��9��Y��;m���]�j��cRS��b����c�^����5*R�$HJ���l� �Ҭ �A��UtQUP[uUQ�
��j�Hj���U������	�⮲K&�eΒܲ��Sj��b� Щ��m��m[����]Uc9���)P��v�` eZ������R����°;;nZ�A�L�����u���T��U:�g��C��n��_	ڒ�T��iZ�u@+��FYh���F\]��l$-USj�@�q��j�V�V��Ml��@U �U<�mUUJ�umU\�����UUUU!IAUU[@�5UWN�j��V�eiW����A"�ڪ�������O<���+#���q���94²�n	�]q���*�RZ��Ӭ1Q�ɶ����PU]Un\�R�J״��b��{zl��pmJ�T�UUUK�U�Pq�Ev@j�����y�,�,�`I���<�UR�UUt���V ,U����]��6�*��ԭjv���;UUUUUJ����� �R�)5%·Zt5UTQ��v������d �(���
�ٌ��UVճ���RUV�c��=-�Wj5\ی�;Ȱ���ԩ�����]�β�ˤ̼I�I�b�-�
Mȇ���[U�Y��z5uC @�*����U.��U��UA�)2���uT�{p��2GUuT]K�<�JɌ�8�6�fiP.��-�%��Zt�;Sj� s����n�1�q�`VM�^���4��#�J��Xec]5Tqm)vV���
2@�<�PR���K��<g��)��s5K� �T� ���qn��³hZ�֮��V��mXT4
)�S���,j��խ{ �ݰ&�z�p۬#Qӂ'��k(Qp@)r����Un�m�N]�݀ҘH�F�������i�tU�xA��u�Ԋ�n7fدQ���皣rp��Ol�<��릗V [F�T���4�Q^��Ūl��GnO!@#�5�^;:㱰ն�ؒ�I�lr�=��T@U�P���q/�iV���e�� �}8��02v��T]qη&���8Z���
���)�v7�z���P�B^y���U�K-� ��3�K`o��V��c\��H�nSlR�5UWUl��۠���6@8������:)UW�܍U +����ݷv�6'�;P<uml"����$
�����/>�f+=��W(�j�U*k��V����V�1Uڇq�"�5�V!܁��`��y�Wa��*e3���eF�j���M��V�Uj�����Ujڠ*�j�/]UT,"d*���l[WU@T�&�UT	��]�WUuV�UmRдي�[t׮I6���ۃ�4�n�t�X��cm��b�� uUT�tQ���T�mUUT�]J�������k���{l����iV�8��[B���^�D]mU*ԫUsg�i�I��M�i�muQ�9�(jfvy��`88��=e�
�
�������U��UV*,��UUUUc!(R�������A������eb�Y��UUUUUUUT � �X*�j�K#]ppWT]���PcV�UU@UUUUUU\m�Z�j�Ub�Ml�Uʂ��Um�>�
�����Uu���V�R�Q�s�Glu&�� UUU++SUZ���r�n�UUm�GC�%Z��e�Z�P*۪�n�@H��U@.�Hm� ]�UUT��k`퍫�u���j�C�5+8�j�l:��Nꪪ����mN+�9��ccf��5`dS�	���e嫶�@�R�EUUUJ�S���P3H���t��ٸ�jtJ�UAKUUUU�)V����
�ꪪ������vv2UJ�T�����Un������Sc�*�j�T
���Z����U��T�j��WUU�UL=���=MR���e-J���6��U[xlB�\�$We��ݡ�{�0�P*�q�ݧ��讨
��f��l��Q*���宩���=+#x�y@��l��c� uU�Z��)yzR^����v����V���������b�ej�*����E���	����P�mN��]B�yhV�)@�V{ev�Z����Q�mCl: b
����F�y�5UY2�L��j�����^ �n���B�1�J� #��=L�f���3Gg���H
�+��r�̸)RYk`�WD��,S��qU��ێ�c�`��g�{;3�华��C&ోj�����a�����8تU����+j]�j
�Z��(�P�)j��n0���VܦO[pU$!U$ZYj��{U.� *ک�Xڀ�U����2N۟Jɮ��(*��.ؗ5F �3w�@ᱬ��ڍP!�-ST�U�*�.Hxeݫ��.�b����Վ�6��ꀭ��lc���Rܬ���kg�;����A�!V��6>��~��F�g[uFG�m�j�����r��o����������B�m%����1��:-�U�T� N��z3J�u�%8����4�N��[�ﴜD�WUPQl�mV�j�
yU�WT��[m�z�U�X
X +j��`j�Mvj�[��
���j��<�UUr�\몪�U����^���x�Y	��
�j�/�Q����������Z����nZRY.�%�����%�����d&�V�SUUVҭJK[U*�Ps��U�n0UUUU*�u�u��*�UUUPjke'��mOR��\�*�l�j-�rI��[uʪqtE���I,pUU[@�N�Z�j4F+����[UUUPurүT��UQEW���R��WUT�J�Y ۲� UUUX�
����U��h .���P�Vݑm�����+�#�����m5T��2�d�{E]UUPNVV��:� 
��ڪ����Yv@j�v�S��ɴ�̤�J�$�UUS�nʲ�UUJ���*�uX��k�����������:m5ƕ�V�:����*� Q�e%.�m�e6�_𓻺N���h)�#�p
�� g�A����V���^
� R"�/�@O}vGQ0�n+� b���� ��l]��h)�ǂ�H1����p�b��Q��@">�����`@X{�T�` >�'�8)�Ϟ�"��!瀆�}�X�%(A �B)�T�l�����x��a�OD(!���U����Q!�	�/؊x(z��Ex�@MpDC`(��� ЈiT6z�#� !�8T��@7_QCbG�~���E�Q�� iP� b@@����0��B A��D<�M<���Dp}D�|�lP0R )�#$I0A�%Q�#����W�� �Q|��9�-!jZ��Q��t!A� p 6�P��H�F �!F� <���<P��$ �Ux���@U|Q��z�Ȃ�P"���QJ�]:Y'u��|<�Uz��&��m���c*��m<����`��J�Î|�Y#=	��2ĩ;t�nk+�!=��W��vMڠN�)
U�Q��p]������i+��2��=��༼�%lDcr�U�Vs���v	�i.���l'�X���s�s�"0�YQ����z딤a5���k��t�S���C�>7M[ ��M��v0��Z,�pm2���0��UBL;[' $�)T��]֝g�Wam;$��[��&8k�ULn�b�6jvr�q۞
������4q���N�YʛA�n�r�2d4T�����sA�s��3�v�T��ќ���qpY9bq����rBb}.;j�{q�:p�%��p��Y���aμ�`LaSI��A.i�9'�����j��UYmE�b-��Ka[�5�����+s��@����h4X䠝�˧����:�lq�M�e6�eX8��T�����*ju4��ڶ���M3�+H`�vٕ�c�6�C�N�;�q�,�5�u6�n�f%	i#4���H�\L���u�z����&����wci�4�g�	���r��%�c�s�1��&�m��\aI�g�l�m���\��2c+��#�=�'kVp�$�6d�N��# ϴe��vL�0��lm�Uю��,�R��OF`eU�&������Ip��b�Ns�n�0f-���:��C�v����s�l��vQ���]�y�W*�����Qd��n�M�6�8��'n���v^����Y�Ô�l���� ���e���i�WEV;8@ۓZ��67�F��q�ՊQ�mX؝1g��eN,�PP�q�,�K�GO�av�RI�
.ˁ����ۋ�p�!b܏b���ۢˎ�������T/@Sc�]��d��x����HFEc���e�A�E&�^8��j'���U�P@k4d��]�\���N���q�HE�b�[�5��u�4j�Et�z*�6)�N�~Ew���!�'���N�:$���Mi����3*ff L��*�t1��s%ɯ(��O�W.�s%bCb�@�6d,D}���'#@�,&�J�\1�T���Z�d1B�j��)���fR-�&@��:w'4n��gal�X}�]��@j��),ll�:iKY�(�Β�l�������Nl���N��*���3�@&�2�[W^�Ib�������wN��k<��K�4��\[)1 61l6����"��.2�_!�q�����a���Kс�����|��������V�W|o �u8`Se�m�X���n�*�TӴ��7m�� �/ �\� 7�<��p�;"q��e���h7xݹ odxz^ŀuM��l6���)S|N®� ������ �/ ���`����{�!�6)s[���b�;��Z�PΛ��:��1������� l��av��T��:���>��X���Y �[�˶�v���~�����UO�� �+Q��(eU������}˹$��~��w��/ �wj�(�����x�8`�G�����`�=x��ic)S��v�ݻf odx��p�:����+��3�����+
v�WH��m���`Se�w\0{#�=ʪZIw���������B2:�d9�S]�ۚ�rv$��[��cw9���j����H�{7C���m���׀}�p�� �e`�8�ue[)+��w�w��`�G�w�p�:���${����e�N�m��o���ԗ��r�D
�E� �����Ϲ��{��X�s 6Yv��m��/ �/ �ob�� >�mD�*-4�;k �/ �ob�� �d��H',j�WJ�6��0e�*��Y\`�f�g�����%j�w	���s��APYF���[�bM��Is� 7�<�����x양F1�EۻM[Xٱ��H���+ �}��7ob�%waWe`�.�6���yX��x{�\JK�X��x��V���ڵn�l��`�%��ذ�c���Q�*�R@#j�=�����9�N;N���J�n���Xٱ��w��^�6*�eݺuoA�Y�G+GnMm���\����:ה8xY7U�w[82��l��EV���<z߶�^��/ܪ���;�<���ܼ��X��w�����^��ŀ� >�l:��-4؝��w�"�7��a��y����`.�TER�,��)�����f\���}���/+ �nE�w��
�R�V��v�������L���%Ȱ榖�#ZbᬜL��J1
��Yy�Bk�L�Y��ͺ��!��J5T�J6V;a�:(�ƽ�)s��F�&!��f��\�[�2D�.�vyD,�G�ŷiM˨��hJ��m��;0���r�.�%��5��;:2�#�(�\+s�f^Iv{ej�P��Rr�)�<$��;�tX4���R��:��4JP�S��}�o�S(��=-�3�6�������CR�1K
P+lF�]q5�XW1c�H"
��ee�f�jE������X{r,K�`{#�$�ʴ�7lN�M�V����/?U$I~�����;]�� ��ӫ)1
��xݹ vlx{ke��%��9C�U�v�e[m�r��q-���7mO^��^�ob�;�����0t6�x{�e`�%�m�Xٱ����<�I�;M�mu�m\�mHa�*�A����\v9b�ұ��E-2+͚�\πy{��G ���ʮr��A���V�%W�N�E
ۻ�x��;\9Ü�!\���F�R��3=�[�y��� �܋ �uT� ة�.��wl�͏ �ٌ�5vK�&�:l)r�;c��]����[����5o�x��X���	!2�m�����[l�:�%���`{#�;ۑ����	ܗ�j*Z�-�4���������+��2a������fX�,�%�;= n��ذ������ �엀}�r�uWt�6ݕm������w�܋ ��ŀw�(UyE �L�w�^V�܋UU�`{#�>��Z-��wwC�m]۬��&�`fǀvl���UN����X�p�͏ ��onE��mҴJ/��ue�'@Ӵ]�v�� 	�l�@̌f ��;Tɳ�.��!Ce�;I�N�ٱ���{r,w\0	�aK��퍂.�6��%Ǟ�s�o�X��� ;6<HL���ul:�ڷm��%�G �dxQ$x�v�,����x�p��G�v�p�\�.���/ �Z������h�vـ� �UUm{���5o�x�Ȱ�k�G#b��-�=�.z�����m�]�G���y�Ҹ����-
�ten�\�6��;R8`]��ۑ`{#�>[�T��&Z��[h����^z�=/�X��<��ݽ��S�0�݈wm`nE�� �r���X��!E�HI�V������R\x{r,K�`�/�i����H���X�Ȱ��krO�x+A���mbIJNy<|��\�T��5��T��m�ғ����o�p}�!v��+z�f�U
7�BIi��F$S`���P:���x�pge*z��i�{=��{l�gp�sZ�Pe��9���:ݮu�-�ȟ���q�g���s��;r�:�A�4m f�]���y��sl��!z��g��g�[*q�S�(��)��-Y��Q����`ڹ��&W-AF�p����X�R�L�
�8���J: ��V�5�L%�%р�\�ȑ�Y������+M���߼�ˑ`{#�;��X�r�N��mj��6\� ;�݉� �I/ �Z����tբ��f n�xv' �H�	#��%
�)� �:�o �� >�<dp�ݏ �M���	0�V��V�0�#�$������6�k��d�����U$�-8��)������֫>Q��V�٥��Q����ГM�dp�ݏ �����KIpm��z������� ��a-ܒ{�k~� % �T�N}\�&|��G�wnE�}�QR��n��W|-��uj���G�v\� 7v<d&U�j�X݊���m�)%�ۑ`�ǀv��X�r�|�]&��U�o �܋ 7v<�� }$x�[�G��/	�tժ�WLi-�!4�J�(��5Щ�k�l8�uX�c�A������N���m��$�xa0���	�"�7d�V1�C���t]�o �#�z��ă����~���˿kKZ��h��!*��Z�������>�>��xGӄ>�4�V�Ot��+�a��l��`2L�8>1�Bh��P��t��Pخ�gb��`ŉ�-#"M�z�d#E&��!��3�ŉ�!��`ŋ� ��g|uf���En�.�ox���� Y����j��V�ܬ�$oU���e#�'��&k��M��$�O� ��\ s�N*���T�� ���Uj�AR'�*. l��*��Lٱ���� �wj�)�I����7nE�ݏ ����*���~���T=�CeҤ���� ��xT��/ ��X���y�YT��َ6B[/W;�6Ӯ��&�>�ӻAe3�n݇CVUƛ� qE~[7�~x�Ixˑ`�ǀl�ʺMZ�vU�vݵ�I��X�����,�	��eZ�11�v��6\� 7v<��� >�<ek�:g-_�e&�X�����, �H�.�J�T��̮d�g�7҅Xƕ�v��;[0�U^���/�X��:�:������v4�Y�����Q�n��d�Lu��Ts\kT�+��"�"���m��;?y�����[%�v��YN�L������;�� 7v<�� }$x�-�⡻��:Wn����F���#�;�� �������U��_m�F���#�;�"�ݏ �	�J��ى���@>y�@��=����$�ﻭ�<�}���(&�� �:w;��(�֖�6ǪS=En��&uƒ3��#�}����z��k��N�+Tk��*.���q-���Z2�Zց��.kq46�J`%�C�^��P!	��sq�9����g��:�>�wB[f��zu��%����P��m�kw
�o]D0�̩�]��6���S�d������2k�՛��Ɇ�DxW(q+k����KfpV+��#�d����6�jݞ���scvmb�ܺ����3�3�d蒈�5�p�ŭ�W���߼�wc�;[0����I&>&Rm��ݏ �"��ǀv\� ��B�tP�eպݷ�wmIx�#�;.E��<�$��B)�.�!�i��͏ �����R^���,��M�i��vG�qI�?�����G���v�uZ���EΕL֫0�3kД���mvL�ڧ���(<v����.����Z�x�����9\��{��6���xF��B�9�-�m��&L�ʫ��1��"�ݏ=_˳�����Ӷ�Wv�v� o�ߞ�{ n�x�'�$�2˫wi�����{ n�x�w���o��C�RC-��V����ǀ{�=2�� ��E�/ ��{��:v�t�E�]�t;4�u��؃��GR��6az#���$�agc ]��U~���^�x���^��r���$��5o�-�,B�4����<�Ǿ��Ii�y`�� �ke窩"lw�YE�+v�ڴ��=��� n�xmUWܪ�����tX�]�k/{��O}�u�!�؎*�J���4�X���R8`�G��S��X}�.Y�ā���x�r,�?U_��ϠO_�� ;�˶��k]����R�K(H��Iㄈ��`y8ݺ5��B�]z�lm�9=�ݒ��Zj���N���cg@=?~xۑ`f���9_ ��?��?S�iӵl�6��&܋?r�U_��U\�	�ߞ��~� ������W'��C�RE7Ʃ�ݻ����	,�xz�T�'��/{׀vIIb
j�0v��)���	=�E$�s��/������d��h"����� ݑ�I/ ;$x�R^���+��=�,�[�9�T6�Z�es4�HR��~��3��5��Nې^�a��
d9,s�1�E�[/߿^ vH���� ݑ��D��h�#�e�m��f]�Z����m�{� �d��l)r�wJ�j��m�dw odxz���/)�^ o��6*�Tҡ��]۶� ���	��`fǁ��=2����~t4�n�ݴ�m��E�/ �\�~��ߟ@������'�}��$�,��9''!NI>����C/en�g`�'5@j�٤7Cf3��3i��;���l�S��C-��܋��9G������^�Kd��>���#0��d]�)6���.�gk�k�C��.:Ty	])am�����}_�)xj�l��h\�!l��;�U�8B ٔ7];ѵ�y���:�fa29���sX���#<�J<�(Z.Wi解i�}�	��ۡ�c������Tw0Ό�6��F.�=n����]b��ʰ"ʷ��yv	ݻ��|���^ od�_ �����z���1����m�-l��U$}�yzz��c�s�U\Hվ��IP픶m����o�L=\�W*�7���'�O^���,��+�ڷm�+�W9UU�g�� '�~x{��m�iih3���o��$-�e	M� ���W9[=���	���7w�/@���Y�i�j0�M���c0��Ь�̩[�%��B� �m��zv�l�_�Iڥ|-���k� 7�<��_�>P?{�@�����Dm�3�V����>�[�Ac�
i^���_������;5��ܪH�xO���uwn���m�V�׀����Uw�Z���~��I����Wi�ZI����� ��=xٱ�z����� zJy!:�9Ge��ɶߎ�=x���� odx�{I!��N��(�\�{<��qÈN!ώ���#����e���l#u��7Uv�[8��=y����`�{��K��/���f����:�!m� �7^�i~Zմ��ל ��_�� }���{Z֤����Y\-cN�^���^p;K�wl�!��R($�*�Q$!+W�	�U}>=�?^p ���l Ϻ�hQ�X*Fɠ��y%�-Of�� �y���f��ZI)'s޼�s��A�KJ���K��̼���kJe�Y� �g�8���l �w�Т-i��-[	�Wr�Ķ�!���Un���o.M�#S>��"���5�� .����nL�� ��y��3q�ik� w=�� {�_'Uz#���KM��̼�JH{)�ǰ �{ל ;۔ߔ�f ��W�S�Ky�e=�� w2���[O{��� g�~��;��7XV�uWl���I;��� ��Sv�o�����nTM@R�� p��Z�HZ��]χ����4�j�v��{��`�%�/�=���@?z��6 w2�LY�mM8��ղ�Y8j�:�F����x���P;&�A���&����$*B�
@%�i������8���6 w2�}���`���Dz��\RM�� ����ZII �{ל �g�� �����֖�$;�{څ��(�e��̀s޼�I�&��奭+i���� ~�?mM�w���f��#*������t�{������l 3��y��3jl�Z���[{�߯8��_�ݭ)��6�i6 w�y��_�~���> ���� t�ڛ 7��O���> �n#���H�"$b�r������	f�O>h�R��IIQ�ya���i% ��_�I.�-!J���-dȚ	�B�[+CZ�%j(�e���� H�!�&���[l!2� L"ȁ�Rh�a�b#,`0��d�"db��"� ��F�#jB�sL�H���S��!�1�0% V���H�RRV����$$�0HklP�Y$�!!R�1ddY�����c�	<	 B��)xT�"AȲF�32�ƄX0�D @�����7F"I�B!0 0HCj/���=�N ST���XB BFZ��T���C	���YIMl٬��nȺ)I[�y4 �r��ځ��)�
K-)�Ie�HHKiR
��(�6QK�$3�"�m�#�r<��D��$�`H�d##$HD�d�a��0h��#��"��� p5jD!@6��D�Uly��)	j.�@�"1��C(�!95��f��Z�Tn�Fq��j2Q�&�ì�g���r��n1{s��P��UPtO�ƠɃ�_b��z{q��#h	�v�æ%�6����$&���V�6]�e	P�h(zˋL6<`�F.���7$�h�ӍuP���㈢^�U2n^��e�
�mb�ʆ�2n�M��۶�T�MUDoϤ>��5��v�Vm{�U� I�:�b�LWdiUUV�����z�;=+@�UkN����NeR4�sEJ��b1;N�жR"j�(�J�� n�&�����x�Mm),JFz��J4���I���4CB+3w5ƔܐD�К��I^'�( �d4W���h7d��&xls���x�sl��v�)Wc��p�[��k$10�j(05A�n�;mmO��x>~K�TK3�dWi�n�js�8v�Nχ������z�3ʭ�UmJ�5�p�J��r����ZWe�6��m�@3;Z�)��U����7fq���jLT�h8ofe��� 6�\8��:����m�R����%3%�-�/�-5�/[��ܺ�$�a�24�I�j�ڶ�5�w `�pڹ�f��8֣�a��-����5��Gim�v��ʩ8:��H ��;p���SNP�;G�[2�ʩ��];���SN�
�<)�̀0�ʁ:��K�H��5V�Q19�ا4X$Wn������kI�Ja�V�o��������ئn��tWRO,��Ss���R����R���m��q3!4�(H�Fx��%�#�Χv�.����A�@�F2 m��!k��t�َ<�nu�=k1]��q�S�K&ôit�Q�a;Wl�&�q·�|�	�[4r�`�[;M�0V��=�����jGdZ��/l�b�%ݗ�6ַ�@��:�AĪ���R��cm��VU���\��c����F�q���
�+�d���ؕv����(��fJ�`Ҋ� ������9A�J�m��'I:H����;��tZ������x�<�(� �TD��[�f��#����.qB�[���#��!/��t$�e��j4峈g��Ӄ��wRf�Ǒ׳�
����:��L\���-�k��CI�X�i��R{Di�BQ���8_1�0]���ÞXj2Uт.Z�V�Ƴ	j�s�!2�a1�=R�l{m�I=��A4g��u��J���@5[�LB1��Sђ��:�j2Ś�I'�NrNN���`������K�����n�3���U�+=���v)�Q�eiue�-�(ڱDT����9�`�w/8�3jl ;��� ذq:0.���;+6 ���?�I����	)����%!nIow/��h2��p��� w;��<����/�� �g�8 w�$-�b�%�4�� ;��� gaq̀s�y���.���#��
�i�o8���6 ��� gp� �r���u�JSL�I��k],U�R�sX�&H�lf[p�k.z�7$u8+��̀s�y���.��ܾKI}��mM����J5\"��Ym��n{���]�D��	�O( "�;���v�6 gr�Z�꽶�iJ�tq�I\� g}�� ga�S`�;�� ��ڛ �Pe�FՊh��m��v�6 }3�9��ͩ�=�-)&w޼��/tc`����;j6 }3�9��ͩ� �w/8��mM���!R�Iil,p�����*���[�K�$�
�[T�f���kcTm�
�[~��{j� 3��� gaq��Z���/� ���^p ���i��)`��݀w�y�i%�$=��s`��ל }����-i%$�<#��
�i�o8�r��-����k���Qb��DG{ޯ������^p ���
K%	m�J́�ZZK�I$������ x����;ܼ��kI+�~e =�~�2��Q�h��p�t� Ť�}ܿ|�r�� ��y�� A��X:R]���ύ
[�m䶳����h�me�J�&�1W�MYݷz����l��� �sל �r�6 �r�k�g����� �Y�T��p:��o�JH����<M�}ܼ疤��x{�@�F��H�� {��� t���{ZRCٞ�����6 w�٬���*�9m� ����ZW���������ך�]�����G������~���?!���@ȭ+vXl 3��� ~_����y�� ���^p���� vw"�\T�[$��#ӡg']R��#\�6٣�ΌƅK+�
�X�=��;�m��[�آ�i�o� ?c�w`�f^p�����\�ٞ���zm���b����>̼�RC'��� ��� c����${�ߢ�B(�4巜 ��n=�}ܼ��I��� {�� w*ͷz��`F�mS`zI��8 {��� ��y���S`��A
Q
�$��m����S`�=�����|��>�^pkZ�c[��TP�I-pV�ʢ�Eb�,�l�Hݹ�n�g:��i��ܹ�ф��f���{b�����Ɣ�_lڥ����0/%����SGeV�S��=����:��L�ę<�n��]Mn�+�h0�L�Fŋc9����2����]��ےv�96���S+S��Rps��6|;���\uΙ���4���б�ڠ�S*]G&�����/��Pק��$��{��S-(gv6r� ��-1*e�k������۱i�T�Ѩ��z�E%-� ���� >��v ���5��� ��~�`��k��E#����p�w� ��/8 gi�l 3����$�T�2頻��E��nǀ�G��<�{��J�c�S��|-���Ji�< ��� ��Ł�N[�z���}��k
�tS/@'dx��\���ߗ@?{ߞ N�<���K�m�m�k,h�DE�b⍢p��u.s����BUj(Uբ������λ��k�m��<�nǀ��ܮs���x�׽E�2��v��J��	����竜�ap�� =���7ob���N��-��͌�f�ʂ�[o�����<=T��<��y�eDc@�P��Wm7��R^�y�\��	�����M�|�(����4�m���`ݏ 7�[�	��\��:;%�j�d !r�(�SLB���l���M�J�6a����n;(�Mu�i�m��='� od���?W�&���7a�R��ժj�]1;o 6l���U�~��<��~X7c�$vG��Z@�:)��V����x�`���8/���W+9U꯰��� ;��xؓ���ݮ'V����/l��<�{�o�A���m��,^��9#IL ����S|�� ��� ����i�.cupf��o��mi�`���N�fnJ��-��D�M��۶gqPݶ�{x;#�7ob�>@zO<���X�
�C�][i� ���I��, ��x�(��c�z�i�J��v���=/�X7c��[�	��鴀�wN���*�ԗ���	=�x;#����W9\����d�w��S�J��V���t�� ݒ� N���X7c�?r�t��p���	���#��<�H���[��ձ�onj�P\�'�'l��3�R�e�F�������7�e`ݏ�\��'�o ��O��N���յ����Y�r�ă�y��^x;#����W*��{����S|W`�n������Q���W+��y�y��	�RV���[��n�x�+��R�� =���7nE�v<vT���P��+t� N��r����� ��x� ��!'	�~�O��JfcV66&t�������a�8S�S��ܚ���k��:��Nk��;;,�Ў�3���� ۍ�1�z�i�3�/^��I�I�����v�ƌ\�cT��7&D����1[�Jж���W%8+3׊%���G���A㨂�a��I�d6L#n�Z�l@i��Ջ�a�c�\s�lg��\�� �،iu���*��P�%�t�������~�'V��**ۄWSG�3	J��uѿYx��g���,�m�5�Z9�L;�tOw��:Z���n��ߖ n�x�"~�W9����է���tRv�m`�Ǟ��q �{��}�<���$n׼��uj��WLN��o�o >�<?UURSc�O<�딐Ɲ�[��un�x�W��M�� n�x�t����}�>[}��_R�X+f7x�\0W*������x�y��|?6yt�1�"�]b�Ld1�N7A��=��P����Re�U�c�Z7�v	+k 7v< �a�_�\���$�y`��
��o���m�I�O��O�@*��T> �X����k�,��T.�b��2�� 0$H�d�@<G`�0R�@Ch⛥�TU�'�+Y����m���wc�Ur��U${}^�����t�I�������"��� ̝�krI�O�ܓ�d����j�'I�i��7nE�� wa����rK�{ﻠ~��ya�E���P������r��K��O�:��^��6�U@t��7J��	ݢ�c]�s����b�4{�mqu�bTˈ�����I�b��wJ���}�'�|���ove~���s��=�~x���Zj�unڵct���)%��X���{�|�t����ﺾ��*���\��O����rI����<���B���DM�t���6 BV]!�i��":BA ���<�]h�I�%hS@&�9�r�1PĦ�$�!V�KƑH�7T#�H�V�i�JR�@��ZJJ�:�l��հG�ћ&7��µh�Y7���,�р'2��tp��&�� )�V�J���������T��J#�ڀ!�W�>���E�z��]Jvʥt4�I6�=ʪJI����)%���X�%
�J��HN��j��x��v��_�wny`�ǀw�q$�-�=��\4ng`˧`�Vx5���n_k�s�I&���"d�٫�������e���� ���xݽ� 7v?ܪ��v��=��,�?"�)�I�m�n���X������=Ĉ�{��S�Nհ���<�t������U��~������;���x;�*���x�%!<���<��r�ʻ�c�;�r�n��e��m7�j�/ �s��������Q����W*l羸�j�����nr	
l��4��A�g�
���H>�	f��G1�иo�l�ߖ l��wT~�W�"�������WWM;,M� ٱ��Tx����{z�Ă{ޡ[B*���n�x6/<T�xz������	��Nʔ��*(|1�V���9�/�׀wo�X�c��Q�vͨ+G`�U���<���Nro|��z�y~xT�x�r���T�EX]z��
�U+踸�\���&�֎H�a"F%�X�j^��	L��M��(��T�C�.�qq�z�>w�l}��c�Fn�^N�����v���Mn� �Ҩ�ֱ����n.���M�\L8�RbŻF�n��@z�MZ��RZ����I�r�X���z��\�y��=�B�ORrtL�v�Q֎��\0Q�)?:I:HHN�law���z�����rs�x���d��c���ÿ́�u�8�CO�ww+{m��ౣv�����x��<�l���݈A�1�N�wCm��Q���5zz��?�c�s���G���hcuht����v��=xݎ+��\�Ur���~x�ߗ�M�'U�M�!��&� �܋ 6lx4��=\�r�J_�� 쎽M�U��N��k 6lx����U)����=x�{�Q����;!3�lT�Q�ٵ�t�f�%��Fj#�r%�k0�%l�aѼϷj�o 7�ǀun��>ۑ{��+��>@v{� ��{��R��6S�E��un����@���U*$?�> ��*���g�n������=��~��}/aV���6��m`m�X�v<=ʪ�URQj�xv� l�EK)�
�d�����ZII����:g��}�ф�9\���� ݞF�m;���4��5ulxݽ� �ob������|��͌��b-m�P��O��kHl�Ӵd��c�����ǡ�~�{�پ�֫�ݍ�I����,� }ݏ�k\̆zm���E�Q��Q8�	L� >�ǀoon^�ob�s����u�m򮮛�V	&� wg������D�>TN�y��gyw$���n��+9n�Rt;v����x{{�c����w�x���X�*�:c������X�U]�<� �����ٓm��E�h�-����Qb�z變��B8����A��u�f�,����O��wV;m�Xݽ� >� ��ܞ�ָ7����３^�X��D�L ��<�s�ĉ�/׀n���>�̬vA �j�R����{{r��{�9UIw}� ��<zk�t�iһuhv�v������s� ��e`���9K���/�c�6iI�g�4�J�V�����=U����?��T��>��Xt��#�7We�CM[���N�
��m���H�X���y�Ju����w��ut�ڰI�> ��<iwe�v�/��}=����y��L�T[��m�K�^{�*��~��	�߲���yꤏo��X��t�t�t&� ����;5� >�ǀm.�xT��%N�m[,wm�X�R�O}Xݞx�엁��W.L���z���Rav;�t+k >� �\�rU��s� 콋 �+��A�E�`D�j���/����X���bq�P7;26�bmIoUŒ	���mn]���
)�KU�ap-����P�3:#��=:��\�<�j��u�����[O�4Ny6�q��f�̙��5�rp�z�N3���]&� o�ۃS�ȃ��cgk��Óf����֖�����ҏ.� ^Xۢ.�˺����D���x�[ј]XV[a2�-A��ӿgFt��t��>J?�0�.]Z��F��QĦk9�x1Wn�BNf0��F����'$z��v������5m���~���ŀvG ���5ʺV�:Wn��.��v�,�s�H�\�����ݗ��9�i羒���b�ށ��N�}������p�>��U�ʺ��j�v�r��Iw���&��w\7'��!�s���rI��˟�Rf�eE�m�{{�v�,���x���������h۶�Of_��{c���q�:��d<
�x�2��o���׏�(!:cb��@�~���8`������9�}������������&n��u��ܓ�>��u}P_y�ɞ��nIͽ���{{��*����,.��t;f wg��v7��U%ݹ�n���7�(Tb�&ںT����r�J\�o ����;�p��UR]��He�N�*%v[v����6�������w�x���6T�����ˬ��$��\c-v��pl�L���4�2uP&_�K�+�-�j�1W|�>���x]���/ ��V�)]�J����y�RG��7�uI��o�6��7�b��9cQZݶ۹'�ﻭnI��f�H�?UR�D� ���A��g�o]��O~�� �*R0|T:Bt��m�~��~���$����x�J\�o ��J��Ui�M4�ۼ���ݞ�o �we��vK�wL�m�]�޶�����n��tc�鸡*���,�sa2ܯ��;� �,�w�t;g���n��x�v^����B�16�ҥwM6�[#y���r���~����`۱��\��i�:�E]�����{{��s�f�ߞ�?~o �
N6Rj�*�J�M����)�y`d��$������ ����ky�7��U�3�vV� }���ʪ�\�Us�����^���>��v��癎����ԣ2[�G�ZD��E�΅B�-K6\�#\�t�Qr&�n��.�M�oc��/ �����9��|��x��R2�H�ĝ2ح��|���ܮr�������E��ܮW*�:�R�'tՊ��v�ۼ��� >�Ǉ��U%�s����� �J �U�WN��� >�ǀM����v^�T����x)V�m�J��4��"ݍ�-�xݽ� >ݏ ���9��W���L)$�R5 T�l4�֐5��dI$ |� ⤁@}U�d'�5��kɽ�С�Wf����4rI�i`q�4)��֒Ɛ��5�1@�$�� ��l�!�	  ��5ϼ��k	�u�s �!�D�j��i�	m�&V�X찹B�,!�Fu=�ZBP��Xw`�LH^���b�m�yv����$:RY@T�C�R)ևt��Ts	��Zܘ³�� ��2�e�s]�+v<f��8���."\O�1�)f�a]��ȎjJ�],t�۶%"�h@1F2��&�=��J�Q+�Xؘѵ���b���@��ّP�X�n�*`��X��q̴�i�]0ei��Q�,e5���9P�7+J�K[mp���NL���l]hrt�yy� ����mk�Z�@�7K��n3�uװ%�j��uR rQ��ɰ�9��ᖈ��X� � ��<j�8�m��@֠PWYV�U�Sc9�8@
q��Y{:R�1k4!I�^H� ���K��mf���t�0Sm.¼f�ᬥ��y�k��[u��I؜X�]v�Ȳڕۡ�ʷ@m��D�AN�&x�g�z{4�ӎ���pӔ54m�\4�����]> �@��@'��^���)=�͍���	��<g&�#p���yO;]z�7m�ι�Lu�Ɍe�t�c�˞Բ\˺�JnRG.�$ꭧ�6�n����N*��Х�����um� P�ikl�.iiuk���R�:�Yɉm���*��vZ��.#k���b��:���+r�!l
���Y��1��H�#��I��6���yn&��<�(��UI�kW+����Uݲ���5T��m�W!$��
�����T@S�[RQ �R墨�8ڀS:Ej�d��G]���"��-e�V�s�lJ�v���=.����<ɒ����c��D��m�ۛ��oX�w��S��ýl�n��u�u��l��ӆ�r�!�<��G#c�P�u�B�2��D�,���1]X臓(�y:�˞v��d4�F{v�и� Y�:�Ze�ꮷdsgd�Z,�-�U�R&ƫc�m�x���O�Q��:�P�	&I�)��S`G�t��Z�\n��&jp �*)��]�����x"	�=O 4�0 +E�D�j�"�%��߶�b�B���sьv
�q���0i�dq�î5מKkS:�\��*��u�bA��-��V�J�;����y��ף��It�k�����xڇ3�6�v�\h�0)���n�1*$Cx�T<�%М�lO;�m
��m��p=8�㣗k&7%Ƿa'J'!VP\��[n�-��Lv�}WI�i�I��=�0��v��/XT+칈�0~��O�O�.;�^\���	�Mɱsl�<)�`�*WZ�M�e���aG���8�P�dU}/{׀}�ذ���s��+�;a�O~o ���'������]X����ŀnǀEݍ�-�y�������<��+)���W`+�`�ߞ6�;�>[���0�jբU -�v�x[���/ ��� 7v<vT�e�C��i6� �I/ ��� 7v<m�w�M���n���X�M�o�m�6����w���vP0p�5#^������dkjۚj����ݎ�� ���	��g�Z��ǽ����M���T��ـ�<�NU�p���xT���0�@�XSwi�E]�]��	�����^�c� vlx�U�[��:|���n�]���{ vlx��� ����gN®�Ֆ��m�Xٱ��#�Wd��a�&sjƉ�G6ģ��ٌ<k�[G��@γq�J�5Qc.I
/.�[��͏ �r;�5vK�|���� o�Wv�qV�1�m�nGy�s���׀vy��͏ ݕ8���P��ح��j엀}�����Vv���xRF���`Ʃ]ۦ�w�}�� ;6<-��Wd� �m K*�݉��� ;6<-����+ ��� �tiQ��Z��2�S�xL��mF�Lт��Ȗ���i'u�w;�=����U��*mS��tU���o �v7�od��>�ȿ� 7�� �����UiӦ]��o �ɕ��I��� o���o �o���bW���u�}ۑ`fǀE��7�e`�u*��QcT�m`fǀEݍ��2�;�����t&���aJ��P�i�4)�9$��nH�	�DߨG��}�w��rI�ߌ�g�S\Li[xۑ���+ �c� vlzϧ��m�[��i3���aa�s��;0r�v�d�ƥ���;5}��gyN���M����{+ �0�c�&܋ �o`1&�J��6��68g�����=/�X�L� �hYWN����;f vlx�ذ�r���mm������ٍ�n��%$R[p�e��2�	ۑ`z��ķ�� �����7M����m���+ ��� ;6<.����9U*+�Ԯ�5���N�cP��(�q6���MH�ӳ�����(惒�`M)��gmȽx,l����ô#Vǌ�05�3�i�ni��m� ����7c���Ф��#�e`�$���1�p��L��<�6��R�#lQ1� 3�nְ���U�ܰm2���pun}W!�ԁ�;tuų�Z��t����N]�F�N5*��·�����Hu�{�HF�����Fcj
�-3.�њ)��)(3<�k��l7,�.Į�T.&Y�������͏ ��/�W��+�퇧��X�οU�L���e��k ;6<.�{&V;{~�+�r�v�z�Z?U*�O��+o ���׀od��yĤ�0͏ ����|T_-]��s�[�>�O?ٱ�l��}���>6�]�M�u�M������<��x�L� �O���i��`��⭆�3ZJh62$u��٣�E�f`�;������0�c�&܋ �ɕꯐzy��}���PRE%�m���6ikZ~D���(/9>�\ٹ'�{���'�ܻ������/�(�R�Q�m[l��e`I2��c�7ve`��;��'�i�m���s���{�����7ve`�2��J�X�T�;,�f vlx�̬{&V�kn���G(��tJk^p7�n�47N���)��ɛI��f��Ț�9:�h-�wfV��+ �G ���	�y��1`�U���<�ﳒrIi�y�����7u�=Uʤ����L)�wV;v� ��`fǄ���W��
� ����S��@|y�w=� ����	%QR�L�7uj�l�͏ ݽ� �ɕ��R��<`��!n����dD����m��ֳ���{|�`fǀv��Q2�N�v�]��Z@]�r]���#�-!t���b�^=�%P��J�D[i)��~���o;�ٱ����K��툥�O��-�m��n�	�� ;6<mȰ�[�KH{꼦�T�m�W��吏6�X�L�lp��ڻ��R��*�Ҷ�=\�R�~��&��Xߵ�܂n�U�6�Y��krO��������i���{&V���?UUW�g�.�O���	ۑ`l���vʜ�
u<�vh^l\�a��d��n:�0Z�Ӵ�jeг$���ۍ�t?~|0�c�'nE�|�o�����+�R�t6��]� �v^;r,vL����h{�6'���"G-�m�ny`�e`�� �v^:k�n�7M5I��k���}X��������� �)�춝�����X�p�=�s���������7�e`H/��F�JO��Z�5n��Ctaԩ�lګy�kB7O=����E���y^#��`����ڛF.c�,�j��V�st�Qtq1�:�g[Gb���9�݁�P�P�݊��;���,��q=��2�t�X6��%v����s�%ۜ����3�Y���+�f*�]��-שj)��i��]����^�����f+R�+5p�*����xs����[�d���-�nģ�W3#`ݜN ԇa�=J�Ue:��*���r76�I�vO�>���f�`�2��p��ڻ��8�&ZV��{~����V7�� vlx�H��()�i���L�v8`fǀM�� յ!I6!���t���'d��͏ �r,Ԧ��V��TW�B��eZ�`fǀM�� �ɕ�Nɕ��ۨ�S���Z�k=�%�X1Pe�WK��e�ݷ&�k ��5�ج�qۡa�K�n�K������+ �ٕ��4�*ݤR�y\�o@���;:s�䓐9�Np��s%W�U�W����}�X��x�س����zK�Y��P鲳�{��{:ٱ����I{ny`}�鮥.2��wt*�n��c�>]�x�L��奤�����m�{�li:��	^����?UM������e`fǀw~��Z5�����u�\����ne�D�Q396�0L�0�̯���\G^<��^i����@���+ ��2��c�s����:�z��{�%n�*t;'n���ٱ�.�{&V򒨨�4�*�]� ;6<�ݗ���U�!��r��R�-ϖ4��.��Q"{��"�@�!MMO��C�4��4;AC�P����F�i��xy�*��Q�>(&���[�p������H���1�0!5j5	G
l��y�,
D��`��<D�0�D4��E؀���{\�Ns������ܬ����
�wI�ݴU�+m�z�T�{=x�{+ ����4�*ݻ�`�R��V���+ �����ob�;6�!��Z�cF�鍐�.�����	lU���q��z��;IY7s���yf� ��2��c�>��X�L���R�2�����6� ;6<��ŀod��>�̬ �M�dEP�ګeZV��ob�7�e`wfV vlx�TG/ ��V��{&V�vea$��~����@���DX��V����͛m�|�	P���YV�>ݙXٱ�m�X�L��Uʒo���s��%U�\:��0�;aX���)��0%C`.l\�*��P�6\L�ۯ�7�� �ob�7�e`n̬���I�h��V��>�ذ�X۳+ ;6<n�)6�N��]݊���2��fV vlx˻/ ����J�էt��u�}�2��c�:���=���� ݎ�J��+�i]]
۬ �dx{{ݓ+ ��~ٹ'��UNh�"��"0!ES `�$ "���)$B@ amH�R"�֢�!#�.��5&d�5�]j�Q�������$ły���Ӄ�ٽ%�t[�sG�E�jz]�!.��v��&�] �Z���tr�u']���1m�s*������0<k=l����� ibbTr�/.�`m����+!�X㱡�v���mclOc�f�vz�%�3�9+�s¢��tm��������(朗���6UZ�(n;uS�56m)�I���Ќ+iT�ѷ`�%�y��=�-lp�h	)�fj"��Y5Zj�e4�}eȰ�X�ٕ�=�M�y�(�|t�իk �ɕ�}ݙXݑ�v�,v�
J� ��v��`wfV wdx˻/ �ɕ�|��#ʻ�j��Xݑ�m�XvL�� �$��l�v�*����&V��ŀ��̻m�|�2k�ڪr7,`A4r��5k��1�ۮ4u��:C�Τ�5EvJ㚺T��U�ح�ݓ+ �ob���֗�;��m��1�wD*�9,Tvչ'<�~�Ϙ�"�ϑ|NrO���܇V�xvL���R�6�J��WWBM� ����{ݓ+ ���`k������Z�m�~Z�>��m�=��� ����Q��|t�իk �ɕ�}ݙXݑ�v�,��+慚�c�ڸj0 T�~g�>8>��sh�p)������5#I:�+nŵ�j�n��=����ob�;�e`)*��6�ݔ�6� ;�<��ŀwd��>�̬�D��Ӻi:E�+m�v�,�&V�8r�mwfV vlx�NR�n�Sc�Wwv���&V�ve`vG���ʥ�s� �!�|E�m$��-��>�p�=ʮR��?�ݹ�wd��>�5`�7m��l��<A��ѹl�-����(��«`0Sr�kq�f˦��:���=�ݱ`�2�����(pJ�-��M&�ݎvL��� ����Q�(�|t��ݳ �ɕ�}ݙX)#g�����$dt�(N�mQv� �܋ 6lxv�X��UQ��,�^�(n���������ݪH��6<�s���z{+ �܋ �U��9U%:��e�]�]<�q�ۢ���9����X�p��@������Pu.M+^m�r����w@ٳ+ �܋�+��=<�lOԩ[�[������6e`ۑ`͏�;�7�׵��y�C�hqF�2E[}��, ��>]ݼ}�+ ��Wg
즭 ���6<�d�f̬r���,a���r���Lm��d�f̬�r, ٱ�\�QU�$�Hs��c���)36*�8�J��juS#�7���ͅЋp8m�0�H]p�k���m�3vJ;ID�H���3�I��l�(�o=fӶp"Yŧ5�^�ye�9wD����n;�Ѷr���&����d,�{�in&����h�lV-����ӌ�>��	1R���!6��Ijk��L�]q=�Dh��79�q�p�t��F1l�Q
��]���F�^�s `z�V-U�a��	r�(\V@�4��6�f��;��LvÃ�:�M��==��wc� l���Ȱ�,���N��;j��Xv8`͏ �܋ ٳ+=č^�1[-��i �f OO<�r,f̬�0ʐJ�i�I�*��;o�9�s��˞�ߖ�����wnE�6<t�*�ڧn�t�]؛�f̬�r, ٱ�[%�I�.����b�M;
��mP�gU�`�77:.��dȚVX��5y^����ջ�E�_���6<�d�f̬w]JV2���һ+k 6ly++��Ƚ�� 鱗��Ȱ��N	R�ut	����;�"�6l���%����� ݕVb���i�6��2��p��ݹ|�X5U�R	�V�vfm����~}z�~X͙X��r�T��+ާm X�u.B��k���&��vI].��挛�.��T!)m��v�"�N �)���g�ݹ�fVݹ�R	Q�R�M>]�'m�ۑg�H����6_��fǀN��_�ؓ�J��m`6lܓ�s���H/��Vr��9ʥSܧUŝ�<����;���V�c��U�۬s���9ű�� '��ݹ�fV��R��[wt+]� 6lx��_==��wc����i�~�$��4���<�Z��n�lX8���H�4�6n)���x�ڹź-��wnE�lٕ�wc���@OO<OW�@��LI��lٕ���\�H��� '��ݹ }���tݫ-��۬�0fǇ�R[/�X��V�6���V[��Av� ٱ�[%�6e`e.Q\r���s��b,!#!�!�tw�睛�y��	Q�*+eZ�N��;�"�6l��;�"���%ԧW�C���ՖL��]V����)�^�[w\�.@�筢��
'Mf+u|v�bv*Wv�k ٳ+ �܋ 6l~��l�y`!K��e7l���`ۑ`͏ �܋ ٳ+ ��R��[J�,v� ٱ�ۑa�������6y��;[)2"��o�*�m�z�\�[��	���0fǀnʔ��E*6��k ٳ+ �� �dxv�X*��Usj�ҁc!!	F�2.�5�i}�����xI5��h�4 Ce�(4�!�H"�1�>#~�S� '!e��>VH0B1 h~�hBJʁᬡ�mc@��"�E�zqSየ!=���LtxQ�,͛�f�
(X�&�!�n)��B���H�Dx�� DN]1<7���@	�	.0�����y>�}���sا7�A�Du�OEa9��HD�E�$���_-�۰�d4EHBA��NUvi�>��OO(/� ��v��(�BB0�#0�<�BF4���!!$�o�:�vctE�钎n��Ŗ�k �,6ЖG������l��7Pښ�R�W̠�����L��<r�x�Y���5�{hΤ)V�W�knں����JT�L��Uz��(�,������aexS�x�2<���I|�M�qeEY�v�ni�;���.�eC������HrT6��5�aR�x��u
�Aj0�9٩f����3 ��T���.6J�����FXY���%���͗01��X�[�騐��^v-���ݍY̡r9�-�q�WR
��]Q�!�W7Vn��5��c�}kd���4a��p�e�W����u</�]��f�1R.�Dv^T%p֜&MGA�4К�ŀ��6�������gMls�y��p=�6pv鈉`.K�ØǞ�ĵ=n� Rq-���yع{&{rj�d+6�����`#=���v��3�;,�\��p�ۍ�쭢p�Z3�eIu�O7E;yf�(��xP. ��z���e	q���mn��![�6:�u�����;E&���x���#���sr`-t;��N빫t�ٷHr8뷀�j�6�k���G����G\�1�v'dΡ4�^� ���9�/#����,�p���;85����	�q�z�՘��i	��jy�����.�̅hvl�ֽ��t����C���-8��v��� ��Q����be��ų�l힗��e�ZaN�!<�EgX�Z%��{v�E��D{e�f�����6��4��;Y�S���g�UÕ���Y�&�T�lY�l��v�c@�i'iୣ����Rt�fly���\�����l��g!�Lb�9�3��rsX�Q��3n^.LY'l[ a\�z��񱆅�T:�7\�E��WƦ-a�f�����T�h�7"+���m�e� 	P:��qZx�zB>�f`���vͬD�r9��U��)���f��;iJ�ݚ��R@�����.��]��
b:�֓Bp=G�DLx<4J�z�p���
��*!�#����ә���]�g63��N�Ҽ��ucj�v嶠�KY�xjV筘`x���\��ɞV� )��E6�ːv������8I`ٍ�e�4A�WU)�QHD	[d��^7vҝ@1v鵪��F�m��������+P�qF�{;:�W�I]��h%�=��O<n̨m��z#<�m�ln�1�����]�[b��퓁@�X�Xi��&��q�/H<̭k��Ny�M������[�W��	Y�-^H��ԙu��إv*�6g�>~��`�G�wnE�s�����X��G���n�ā�0�#�;�"�7ve`ۑ`ڐJ�bJ�V�NـwnE�n����\��_�����:k�t�StӤ���7x�fVݹ���d�mi2��&�+e��m�ݹꪮ�g���=��7�2��䴒]�?6.U	#�!A��M5��*�˄+H+H�6�.۬��,�u����y�m�t��J���?V�x�fW��7����o��^CM�4UZ��������ٕ�}�� �k��*R1�q>61�n��̬�0��`[%�ڶ�	SbN�lv��`��w��ul��}�2��j�e*V��Ă�{��?y|w���;�� >�R�n�.6��4�s����2`�e�
�7`i8yw\�;�u@8���!���Ƅ�-[Wl�;�"��� ��w\0	�\��j��ӥJ�-֯�,K���nӑ,K����iȖ%�b}����r%�bX�����q�HzC��c^�E+-nJ��kWiȖ%�b{�wٴ�Kı>���m9�ߡ!� �l�'�9�۴�Kı<�]��r%�bX�}��eD�T��p�{���%?�$��D�{��iȖ%�b}�~�v��bX�'��{v��bX�%���[ND�,K�Λ���Hc���e֦ӑ,K���w�iȖ%�by�w�iȖ%�b_~�u��Kı>���m9ı)���;��`�5�����P�k�q;Ht��IM	�uK1!�]	�{<�WR�j�9ı,O;���9ı,O~��6��bX�'�}�ͧ"X�%z]�������}������ֳ5�]�"X�%����fӐ��"dK���M�"X�%��u���r%�bX�w]��r%�bX����
\�f��L�M�"X�%���o�iȖ%�b{��۴�K��"dOk���Kı>����ND�,K�>촜Ԧ��ә����ND�,Kߵ�ݧ"X�%��u�ݧ"X�%����nӑ,K���z�b������iǤ=!�K�y�(�+�I �ގD�,K���ݧ"X�%����nӑ,K��߷ٴ�Kı>ϻ�ڸ�=!�{�^A82�IcՉ�*�M����P�u��qZJ�h��ܶ�jE��3�1k��O�%9)�NO޾�v��bX�'���ͧ"X�%�~���ӑ,K��;�siȖ%�bw�y5Zr�T���ޗ��=,�o�iȖ%�b_��u��Kı<����r%�bX�����r'�ʙ���g㔚a&ju˭M�"X�%�{�ߵ��Kı<����r%���Dȟ~���iȖ%�bw����r%�bX�}ӥ�$�M:5��u�m9ı,O3�w6��bX�'��{v��bX�'���ͧ"X��RdL�~�ӑ,Mzk����z�0���G)�O���,K��}�ND�,K�~�fӑ,Kľ���iȖ%�by�����K^���'���}���f� (�!6�{V�aR��l��N"5�e�e:���YkkpK.����)\�#7m՛{<��V:
7���6���z�m��k|9�mh��^[��@b��jB�N�X-�a�z尋U��L�8\�6e0e����'���:�� �6!�ӎl�(۩J;������x��+j��ˮ�+E�R"�eq�\���N���{i�Å*�c��\],m�u��k�w��N1�7Y��ku�aJ�+��Ӹ�x$���=�bX�'{�}�ND�,K��{��"X�%��{��ӑ,K��{~{������^��`�B����jm9ı,K���bX�'��{�ND�,K߻�ͧ"X�%��o�iȟ�eL�b~�w�5���kD�.Yu��r%�bX��߿fӑ,K����iȖ%�b{����r%�bX����m9ı,N����k)ssY��n��ND�,K߻�ͧ"X�%��o�iȖ%�b{�w���Kı<�{��r%�bX�}�ΔѪ��4fI.f�ӑ,K��߷ٴ�Kı=ϻ��r%�bX�g��m9ı,O~��6��bX�'�@?���]Mn�]s��t�:).�dgex��PY�u絹�s��Y���؎���4�6[�,K��;��m9ı,O3��6��bX�'�w}�ND�,K�~�fӏHzC��g��p�M���+-���Kı<�{��rF"A�������� �&׏�=�by�۴�Kı>����r%�bX�߻�m9ı,O=��vR�V�Md��j�Y��Kı=�]��r%�bX����6��c�"_������bX�'���ٴ�Kı/��'rS5n��%�]�"X�%��o�iȖ%�b_~�u��Kı<�{��r%�bX�����9ı,N���S��X[�ә����ND�,K��{��"X�%��{��ӑ,K���w�iȖ%�b{����r%�bX������0��v��'a݄^`B睮�,�e�"0�.��-�����4T�F�C+�O���4K���ͧ"X�%����nӑ,K��߷ٴ�Kı/�w��r%�^����3^�E��]V�Y�.=!�,O~��6��bX�'���ͧ"X�%��}��ӑ,K��;�siȖ%zC��ͯ+4䢲��ZoK�HzDK�~�fӑ,K��>�siȖ0��d���W�B��
z����=���fӑ,K������r%�bX���Ӕ�!�Yn�r�SiȖ%�b}�{ͧ"X�%��{��ӑ,K����nӑ,K��߷ٴ�Kı>��[�d����&f���bX�'��{�ND�,Kߵ�ݧ"X�%��o�iȖ%�b{���ӑ,K���]�fS:Β��G]�$��2�~}��l�k�Va�dI���N��2��:�L�^�+��|���bX�'�k���Kı=���m9ı,O}���r%�bX�g��m9ı,K�z��]I�6�sWiȖ%�b{����r�$��wI�$�y}�shH���>�I���bX��1>X�A-#��W�.=!�Hz]���iȖ%�by�����Kı<�]��r%�bX����6��bX�'}�~B���$���q�HzC��w�ͧ"X�%���nӑ,K��߷ٴ�K��>3q.��K9)�NO��ߚ�+�U�j��|9(�%���nӑ,K��߷ٴ�Kı=�_v�9ı,O3��6��g%9)��y�}b���M��l�SKc�ǔ��v�V���iJ�Ja�#��E���AƳZ�[�]�"X�%��o�iȖ%�b{���r%�bX�g��m9ı,O=�{v��bX�'}���jɖ�ɚ���SiȖ%�by����r%�bX�g��m9ı,O=�ݻND�,K�~�fӑ,K���o4e�4����f�iȖ%�by�����Kı<�_v�9ı,O}�}�ND�,K����ӑ,K������]M��55���m9ı,O=�ݻND�,K�~�fӑ,Kľ{�u��Kı<�{��r%�bX�Ϻ�֍Iud����Kı=���m9ı,K�w[ND�,K���ͧ"X�%��o�iȖ%�bx�߯n�۔0��[i�.8��؞Q��erZ]�ŀ��f�i瞶�p)�5�v�L�y��tmƆ�2Z8�V���H�s \��&�J<�5�]Apd�j�����a�
S	Y����%��W��!_<�ɭ�L���6D֫Tp �O���'c�ڲ�dA2�!�e�D��b���:��d!b֔�b���;H�B�75�8��U�M���:wK�� 恆�ے�5��,l[v۲�l�v�����l��٭B���&n�l0�oΟ��^���/�w����bX�'�߻�ND�,K�~�f��'�2%�bw����r%�oMz{��y��R� ��t�zk�ı<�{��r%�bX�{��m9ı,O}�}�ND�,K����ӑ?#��zk������j�*6�A�O:|�bX�'�~���Kı=���m9����>�]�v��bX�'����z\zC�������*��,VZ�M�"X�%���o�iȖ%�b{���r%�bX�g~�m9ı,O=�{w�Ǥ=!�K�y�Ȩ�;RV�-{ND�,K�u�nӑ,K����}��m<�bX�'�k���Kı=�7�.=!�Hz]�ͯ!I-"e#��U�Z<����,F���4:qgq��Q31�Y��+��O�%9)�NO��{�ND�,K�u�ݧ"X�%���o�iȖ%�b{�۴�Kı>���E�EK)lޗ��=/}��6���<P�{|:�U^>��%��w�&ӑ,K��;�siȖ%�by�}��r'�*dK���O��SE�-�3SiȖ%�b{����r%�bX���m9ı,O3ﻛND�,K�{�ͧ"X�%����)9A�2V�e{��������ޗ"X�%��}�siȖ%�by�wٴ�Kı<���m9ı,N���J5p�6�Ο/Mzk�^�������bX�'��}�ND�,KϾ�fӑ,K��=����Kı?�z|��Q�[\k����5�;Rlk\$��x�v�v�㢦u���3�x�ٮ�Y��%�bX����ӑ,K���ٴ�Kı=�_v�9ı,O3߽7�Ǥ=!�K��^V�%	b$m�jm9ı,O=�}�ND�,K���ͧ"X�%��{�siȖ%�b}���.=!�Hz^��.EGDD�j��M�"X�%��w��ӑ,K��=����K��C��:RI$GDJ@��[@\�; �v�"ČOIWa.���)�"48c"�5[56�&�0䐕�h$Ԇ*a	���l�d�1&�.�D�������v!݉��
� O�Q`�@<L(��TD�{�z}q=Ϸ��r%�bX�{��m�JrS�������� �b5��Ñ,K��>����Kı>�~�m9ı,O>�}�ND�,K���ͫ�HzC��ex�'*��Rٽ�bX�'���ݧ"X�%���o�iȖ%�by�����Kı<Ͼ�m\zC���Ջ[�m ���R�a-��]�
��5Z�^�1�c��R�!��X�u�RJoK�HzC��ٛ�ގD�,K�߻��"X�%��}�sa�I�L�bX��]�v��bX�'���	g��e�#q\���rS����{�u��? ș��;�ٴ�Kı;����9ı,O>�}�ND�,P���=���U���z\zC������ӑ,K���}۴�Kı<���m9ı,O3�w6��bX��}�C�"(Ӗ������q�Hib}���r%�bX�{��6��bX�'�߻�ND�,ia. �bSŠ��M�%��m9ħ%9=���b�H�0]s{���%�by����r%�bX�g~�m9ı,O3߻�ND�,K�u�nӑ,A�H�蟛��)-����&P�T��V����.7ȶ�Μ�0�,W<�6�m5�P�ֵ6��bX�'�߻�ND�,K����ӑ,K���}۴�Kı<���m9ı,N��[�9J! ����rS���������O���r&D�;����9ı,O{���ND�,K�߻��"~\��,N�G���f��sWw���NJrS����ND�,KϾ�fӑ,
0ș�����r%�bX��{�6��bX��3�I�4"5X)%7�Ǥ=!�<���m9ı,O3�w6��bX�'���ͧ"X�%�����iȖ%�NO|�С�%B��\���rS���'�߻�ND�,K����ӑ,K��=����Kı<���m9ı�ڵ�.%��K�<k�v����Oh�]�7d�9�e��snL�Ϡ
S��ߑ��+S��pr�� ]���E����99G5s�k��&���
;*l�;YH9�%nf�7f{vݶ]]e����XK�`P+l�JR�٪��28wb�mL�6]��	�(��	vy�!��,�Pir2)r��$�@\�t���!WQ���kb�Fv+�������w��1�sr�ᕳk
��Rt��{x�ə�le���%��ƈ��f�ʴ �	����Mzk��}����bX�'���ͧ"X�%���o�iȖ%�by�����Kı;���1m�j
)Bٽ.=!�HzY;��ND�,KϾ�fӑ,K��;�siȖ%�by����r%�bX�w�;�tQ[Z�Q�ޗ��=/����r%�bX�g~�m9ı,O3߻�ND�,K�u�nӑ,K���8���&�����rS���$����_��6��bX�'��fӑ,K���}۴�Kı<���m9ı,N��l8i��Zk&��kY��Kı<�~�m9ı,O��ݻND�,K�~�fӑ,K��;�siȖ%�b_��o��;;.s^:k���a�%��*˥�+xlv��:�-e�O������5�U��fӑ,K���}۴�Kı<���m9ı,O3�w6�E	�L�bX��{�6��bX�%���?d-�k!�i���ND�,KϾ�fӐ�ډ���Ȝ�b}�ﹴ�Kı<Ͼ�m9ı,O~�ݻND�,K9=��B�Ď��Ѹ�N�|9)�NK��{�ND�,K����ӑ,2&D�����Kı=�w�m9įHz_yf��(���
e�z\zCҳ�
@Ȟ���ND�,K���ӑ,K���ٴ�Kı<ϻ��q�HzC��,~�V���E([7��,K���ٴ�Kı<���m9ı,O3��6��bX�'���ͫ�HzC��}�\�ʪ
5l��S�����,�$����ݝ�f3��<��H�qH�M��qc�w���NJrS���;ٴ�Kı<�۴�Kı<�~�m9ı,O��}�ND�,KΝ�|`�E�j���rS�������ݧ!�#�2%��w��iȖ%�bw����Kı<���m9��eL�bw����4Ki�,��f����Kı=���m9ı,O��}�ND��������E�C��y���M�"X�%������9ı,O�'����`+�;��JrS���}��6��bX�'���ͧ"X�%��u�ݧ"X�%��{�siȖ%�b_��N�%�k!�l�5v��bX�'���ͧ"X�%��u�nӑ,K��=����Kı>�_v�9ı,O�:C߽��ܱ%��l�qv�&�7J� �t�ܶN�n�Q�),(�lAa�n�lXd֍k%�jq<�bX�'�����r%�bX�g�w6��bX�'�k�ݧ"X�%���o�iȖ%�by����ꚺ�ɔ˗W5v��bX�'���ͧ!�V9"X����9ı,O{���ND�,K�뽻ND��TȖ'��0�5�bڻ��JrS������z��bX�'�}�ͧ"X�%��u�ݧ"X�%��{�siȖ%�b_~�wZ�3�,сWw���NJrc������r%�bX�����iȖ%�by�}��r%�`m��
�����&��}���������N��k�G.�ӑ,K���nӑ,K��=����Kı>Ͼ�m9ı,O=�~���rS��������0m�.�i\c�n.����p}�n#�e.�>1p� ��W��5q,ԋ
Q�˘eo�O�%9)�NOs��ͧ"X�%��}�siȖ%�by����r%�bX�w]��r%�bX�x�zZ
B���\��|9)�NJr}����r%�bX�w���r%�bX��~�m9ı,O�߻�ND�,K���*&�-��O�%9)�NO���6��bX�'s��6��c�*�"dO{���ND�,K�u��iȖ%��fx�Z+���d�ս.=!�,N��m9ı,O����9ı,N��w6��bX�dN����iȖtצ�?=�|�9�+v�	�O���bX�w_v�9ı,?"G���ٴ�%�bX����6��bX�'s��6��bX�'��b�EI'8rNBIhY駳0Ä�V�uާWE;
^�y�c��-e#={\�R��ZR�t������s��c	B�SH�f�\&;A�l��8>Ѵ�Ϙ�1&ܜ�z஠��kA,-629ք&�G��	p�dŵ ��`'Wl��I=��1M�Qr@�Ic\ N�僐Ħ$���U����T~Ka�77EH{746�e�N�m��N�ܹ������T���c���t뼞M��Ԫ�%����ۓ�����me�fNؠ�yx;{Qs���J��z3M�UX�-����NJrS������D�,K���ND�,K��{��'�2%�bw����9ı,K����2LU�`U���rS������=��Kı;�����Kı>��ͧ"X�%�����ӑ,K����g�� T��'Ò���'���6��bX�'sﳺ�r%�bX�Ͼ�m9ı,O}�xm9ı,O�yxk��ۣD�Y,ޗ��=.��wZ�r%�bX��_v�9ı,O=�xm9ı,N�w6��bX�3���H0ֹUW��JrS���u�nӑ,K����iȖ%�bw=����Kı;���iȖ%�NO��K�f���h��W���yscq�o]���ihlTib0�7j�*�d��v�l�5v��bX�'��}�ND�,K���ͧ"X�%�����6��bX��zw=7�Ǥ=!�K��#|���׬��k56��bX�'s߻�NB!��DӸ��bk�^�iȖ%�by�}��r%�bX����m9�S"[�����a0��v��y���MzX��v��ӑ,K��{�siȖ%�b{߷ٴ�Kı;�����Kħ'�}���33��UQ�y>��%�����ӑ,K���o�iȖ%�bw=�siȖ%��	�?~���ӑ,e9)�|���ɓ�P
���Jp�,O���6��bX�'s߻�ND�,K���6��bX�'}�ݻND���'�99$�{���$�8X�CH��#I(܅ND��v1�v��M����gE`�1 e>r}9)�NJro;�6��bX�'~�s�ND�,K���݇�`�'�w�M�$�͖�M��ֳbH$���}�M��K�����iȖ%�by�{�iȖ%�bw=����Kı>�S�l�Z�h�.���3[ND�,K���ݧ"X�%�����"X�|��%E���л<��N�}�6��bX�'����6��^����$�Z
W"�%7�Ǥ4�,O>�xm9ı,N��m9ı,N�����r%�`~����ٶ|�5�Mz~}���������,K��{��ӑ,K���1��}���yı,O���ͧ"X�%���fӑ,K����gu&�Rk�8��vC��^�p<��ķln�W`���.YA��]4ô��t�zk�T�;���iȖ%�bw>����Kı<����r%�bX��{��r%�oMz>�ϿF8�1���O���,K���ͧ"X�%���fӑ,K��{��ӑ,K��}�u��"~$7B�צ����D����r�t�Kı=���M�"X�%����ͧ"X�%�����[ND�,K���ͳ��NJrS�ϑCcZXĀ���Kı;�����Kı;�}�kiȖ%�bw>����K��mX� ��������;�ٴ�Kı?{��I�R��9wy>��%9=�y�kiȖ%�bw>����Kı<����r%�bX��{��r%�bX�}=���(�2d�m�:�ǢP�l-�Om���e��A�4ca�V�ֵ��r%�bX��_v�9ı,O3�w6��bX�'s��6�y"X�'����fӑ,K�������f�jᚶ�sWiȖ%�by�����Kı/}�u��Kı;�}�fӑ,K�����iȖ%�by�ݹp��]M\��ɭk6��bX�%��bX�'{����r%�bX��_v�9ı,K�~�bX�'}����kXa�j�p�f���Kı;�}�fӑ,K�����iȖ%�b_;�u��Kı/{�u��Kı<�N���Y\ŮW��JrS�������'Òı,K���bX�%�{�m9ı,N���Kı>8<y�~@{DŇ��!Pш�=���H�1aS�N=ѹ�_b+���t>���c �} HR�BH+$$����M�����O>IS�� �P�U�)$��)�@�Bi-$�&��� :B�M�iO��c�����椄!�pYH��	�!@�K��*�q02���(idv@�\�0F�},]	c�� d��y����!DXB����	@!aD@� @DG��v)�}�v�����=�̐FB�$P�Q,���7��L,�B��ͮ0��f�<�g[����@t�l�g���L��&H�ʦ́I�m��v�5�E��B5�^��L����.��-��!�b]��E+��J�nDDdѻJ�*��cT��˘"P���݋n��3��(cY�b63�Ĺ�6~�D��Јb��xt�\��fM��,R�).ʵd�k��c<��nu��J��!�u7=���'�6��yj��Lm����:���)V֠�[s���JdZBj�)X
�m�p���v��'2d�5��m-t�p�ݜ#u�a�3�	�ΉA؝N�Ćm�[�%�e�=흵���j"���T����(�t���s�s����d0�蒨�::��׳9ᝀtChCygj�lU��lԻ�8���Z2K�v��U�u��Gj�X������4q� ����gte^
sU]N�P���=�)T���[TK�@-��)������(����cez�n��j: 2�m�&�`�ã;![7g�OR�yͱ]��t�ڵr�Y���6"�h1�d�7��'�OE�S��oV�8=Rm��՜��t	=\�nH��PE�T���9�T���x&�^[l#H�@�e��)2�^wD�PRK%qk��g��6�'x�b[���M��S5K�K��q�f����N���xj�����S�8��W�.�f�F
�*#��q�U��Ur&�E���K��Ј��I2u�����@ĺ��-n5�v��]A��c�>l�#�$�F�˶)�ɹM烛2\���`x�xE���;�pt�t��l�n��v�U�v��],�v9j�f�pٌ-�aѽ7{)��2l6͝�ъ=9��\&�9��́���V������ ʤuV�[���
	WU%\�cc���%U��c�Vw[��3�a�Sl-2�l�ݾ���y	�T����+���%I�Ȏ�ڀsJ�*l�ekr\/w{��;�N�	j���Lbp؊z����<�����y˚�b�#5���$r[�TZ3m�hZs��kb��n��`6�Q�Ⱥ��lH���1��[T�k���Ơ�;b��#��3\�1��$�1*ۋ��<�j8nQ�h7`ca_\nnΒ뗭���l��kǡ�=��V傥!1\8��+2�MH�Es���db��uv�6�@k]B�Sf1
�+b��k6t�ZK����<�fTj;
}��t��2�M�uD���q�)(�r���qWp��$�^��7S4�w��n{���{��ı/���m9ı,K����r%�bX�ϻ�kiȖ%�bw��nӑ,������.V�rA���۽.="%�b^���iȖ%�b}�w��ND�,K�k��ND�,K���[ND�*dK��~��XR�՚��ֵ��Kı;���e�r%�bX��]��r%�bX�����r%�bX������=!�d���5+j�8R�5�]�"X�%�{��[ND�,K��{�ND�,K���bX�'{���������S�jG]+浴�Kı<ϻ��r%�bX~c��~����,K�����j�9ı,K����r%�bX�zh�w.��\�є�0�-̬��bRY��m���ٴI�OG0�=J٭B�D�E��
��O���5�b^���ӑ,K����uv��bX�%�{�m9ı,O3��6��bX��{��5um�)#"��z\zC���w}��rT@9D2	 *@��Qv�'"X�]�u��Kı<�~�m9ı,K���m9:{���^���=�L�+21nT�r%�bX�����ӑ,K��;��ӑ,KĽ���iȖ%�bw��u7�Ǥ=!�H�=<P���Ti�ݧ"X�%�|�{��"X�%�{���ӑ,K��u��6��bX��3�����"X�%�����5&�1�e�am�kiȖ%�b^���iȖ%�bw��u�ND�,K�ﻭ�"X�%�|��w�Ǥ=!�K�ͯ!I(Z����j��B�L3:��#��&�K���1�i�Y��#a�4E�����NJrX��w�]�"X�%�߾�fӑ,K��>�sa�'�2%�b_�~���"X�rS������ �v�����|9,K���o�i�~ c�2%��w���r%�bX��߿kiȖ%�bw�ﺻND���S"X�����3WZ��d���r%�bX��~ͧ"X�%�{�{��"X��!Ԇ�b%�� �ḞD��w�WiȖ%�by����r%�bX�w���e.��f�]d�k6��bX�%�{�m9ı,N���WiȖ%�bw��fӑ,K��>�siȖ%�bw߻�i֮��&a���ӑ,K����w6��bX�����~�O"X�%��~��6��bX�%���bX�'~�y��	�&4��л^�s�*7nƀ�4��{ ��F�d^���p躐MbG( 1nD����r���~��^�� $��\�x��N�8_t�J��:���I&V%�� ��X{RV0v�ā�(J���<H�XRK�>RK�7eDe�����q{��j�I���7$���rE@����	-T��kZҷy�v�����5+t`Zi��k �Ix�Ix$� �?�	��y|S���\lA:=�N�uly���뗴�uGX�2�U��{�;s��@�����/ $��c�`\� �H�U�ZCT��I��� I#�W+�����z��|�K�'vaO�����,����lq�K�a�W9\K�{׀����.��V���Ir,�$� �G�Ik 7�����E4�	[X�Ix$� �r;�$��s�UG
�UJ���y�6sX3���C7�ْ��N���Xؗ� ��.�Y�\��Ό���ݭ��ȶ��1��s:�t��jX��*�%!�Wf� �r��B�l�[���y#�g����pvmƞ��D	�/"/GG&Z���9�wO��H�\�m�:��R/�O� �}k=�8�H]�fm��\��:#'b��x{9���%6�k�
aX�m��O:wBt���rl�����$Q�X]ۘ�d$F�hx��6�����dB�1X���B�aBV�{�xۑ�%Ȱ��x�Ki4�R`�m�x[#y�#޿y`S޼ �G���q")^�**���%i���w�y{޼�^ I#�&��"ݪ��e�R%n���x$� �8�������xg�Z�������E�7x$� �8�������V�MX����DlŎ�l����(r���e"����wT,�3,˃"��G��E���r�<���$��$� �G�}�L�MUݢ�*�[�����ʮJ��+��\��I$q� �ˊӻG�`
���G�H��W���w�y{޼���ae]���aI+o $��\�����I�*R�v�H4:�o ��w�j�^ }$x�G��g��4��˜��K�1fI��J�;U��<Q�u�fWa�pT��E�hFY^]���w�j�^ }$x$� ��w�v�]�,�c\HJ���G�$x�ưRK�>�Vb���n��M� �G�Ik	UϹ\��%H�AHXT_H5�9�}/ >ݏ �م>;T��]�M�H�XRK��G��K������t������lv��"�^ }�< �#�$���(E�;iӡ05v�Ƨ�Wj#W� �0�9�9�2�LgB-�l���3a�Yu�t�x��#�"�7�r���A��z�ڞ�aL��ƭ��x$�=T��=��/{׀l� ݕ)e;J���c��m�l��I/ >� l��[[*�4a9E]��Ns����}��< �#��9Ts�W9++�UV��� >ݪ�j�M;o�m`�#��<Vɕ�j�^ IH��WW��[(#3��ɮicN-�-�G�q1ed�,x�3v�Dl6Ճ�SWI[��;w�H�		2����j�^;�
|v��7ae�5m�e`I/ �$� �G�}%L�MQv˶���)%�I/�G��<��{+ $�r�����`	��	$x$� �$����UR��޼��ZTSWo��m`�<kve`I/ �I/ �yFϡw_eڻ%�<���1ն��'��c]���(��K5J+y�.z��i�5�)6G�b-k+E��L��)H��������NW��M��i��c1p!�����.�Gm M`����u�mw��<���Z=���d��[u�3mi��pA=�����;$��vN�?k{l}�-�l��Ų���B�h��&aXn�')r�5i��������86�'9�#9��w����2C�+��Y�q�a���ٹ�����.�;�r��:��cp���V&���
���߿e`I/ �I/ $��ml�J��@�i����`I/ �I/ $���̬-ڨ�	�[|HJ��-��I�l��"�^�ak�Yb��v�w�H��fV����X��)�,�ui�e�5m��̬)%�mȰI 뻵(^�OG�w#�2��v�R��#��b��|�����@ئ�&���lM��d�|R&˻���l����6��U�]X�M����7�-$��j�UϾ�s��'^��̬eȰ	���M!%MՉ�j�����2��"�>�"�7eJYL�H��n��6�fV��X��Xʤ����b�!
T�wP��IV�}32m�̒, �#�6�fV;�];�r��c0�O�����ܻ=<n0V��͈���Q�2� b6��T��e+����m�&a���H��ٕ�l�$�k�Yie�J�k 6H��fV��X�r,wf�2�]5V����6�fV�����<=��O���@@��n�<��� 0�P$���h0�u)i�"%"RY��ES�o ;p{� (�`pM"dd�V� �  ��@Bڣ��6H���CǄ� ��B��?|�d0�!D<��fD2Hi��<W�H��+��>;C�KĿ*��$*��y����jd���O��[ E)8mU"-ϼ�!Ĝ�"}���t�<�J�$�D$�A�@!AR$La	"l�����Hy
;`��	�+B/���Y���J(<@�*�� �=TЧ�"�W�C`bT�(
zm�0����U\ ��u��{�ܒy��krN{���e��ĝ:����$��܋ $��z�\��'���#�>+�`	��>�"�	$x����"�n����/K�4��l�m�M�5f���tm̦����,�#��4��,�V0x�$���H���� �I~�9\��u{޼OW�e!�L��m�x��ŀE$��$��Ix�6R�V��-4�'m`�K�:�����ۑ`ͪ�j����)!+w�uM���<k�e`z��W(�)*��tHCJ�B����P��|�nI�;�+��љ34�m� vH��ɕ�j�/ �/ ��yo��B�0�2�ͱfJ\s��=�]kv9{Z��Ձ�.\�EarF&l�f��t���mvL�V�xT�~��{�m����EH�J8Z�j�o��z����5zz�}�<jl��7u9e�t4�˷J���T�xݑ�[&Vݹ:l��HJ�n�L��Xݑ�[�+ �܋ �I/ ݕ)c,TP�:m�kve`ۑ`)%�vG�]W9_UU\�+�z�gMg�h@�����'�[Y�:��:n^��#f.ãS&�е�=#���:��ܮ����۬�YU�2�jZ]ڸPL�����h����e.�ֶO���9N�Ti8(Ň7�ŹnB9��a.Ȧ��u33`�[q=������pŶ`;P�ݙ3�m��`2�$Or�^�օ�k=�Sv�w\<�p�v�c��0�AE�I�N��$�ww�/�?]�Ƨb(w6Jv`U��i.Y�/}�%����.I�힠P�fnO5U�V8�۵��j�@;���|����#�7��V vmT�T�[E�I���v^ wdx��o �܋?�I��Z��Z�N�˶�m� l�� od��wnE�j���'d�N�L��cV+�� ��o ݹ��� ;$x۵2�n�ݧm1ݻx�Ȱ]�xݑ�s�]���f��6�v�J�J:(6���ږŶ�(���1�$�f*6�b
�mMեn��[�-�xݑ����[%�"��Ң�n�+gn��#��*���9��mJl.ղ^ջ/ ݕ)c,TS�40j�x�$xV�xV� ���	�H*Un�j�];v��xV�x��xݑ��(����%V0c%n�[���#�7�L��d���s�JU�ށRZ��+��0�+]V���)5Min	c�Y*Zv^Gm/Oe�[��6{� ��2����[��	�1S�,aJƬWI6���Vղ^� ����je]&�:-��M���v�X[��^+�rU�*�R��QG_}����䜻� ��r�gZ���V� ���]ۏ ���M���wI�+l8�w�wc�=U�{/��;�������o�ڱ
��T�-�2���&`�pй��gU  ���ƀ+.�.�6X�����V��5wn<���������l�T���Wt�nݷ�wnE�|����#���x��j��j��0@����/ ;�< �췀wnE�}�U�.��uwm!�xݑ��(��Ȱ>��S+�1��A~�7�nI�~�tљu(E��WI[x��<��v^ wv<�Lt��
�[�e��v�Ԉ"��i�q.e�f���t�K=��3�əi��N�m]�x�r,V� ��x�qK�>�NU��*���+k ջ/ ;���R���Y�W9U�H���VU�;��É[� �<����>ۑ`����R�;4�R`��m�m�w�ul��j���� �d��V�h��i���:�K�5we�wc��#�U�Wj�9�:�L��D��qʜR��H���;2��K�&��%�׶�M����v�"�9�*�Rk�i,b��n�Rakem�#�t��/#TC9Ζ	����$�V������Îq�7;�f^?����;�#9�M=�:֌@\�v��y�On6�ƃg���a�T��]���X1�AN-��/ v{.�n��l��qcq�m�v[1'�H83Y[�ݎQ����t��:wM��I�N����4��aZ��#�\Y��u� j=�n�5�B����b�M{�;R�Ʃ��p��� ���{xT�x{%Z��.��J��i�������:���5n��>�b��X���T�Лx�ˏ �/ ջ/ 7�<��2�n���Wv��6^�v^ odx��w�vD�����P+w�j���� ���xT�x�םyQv�i�tթ�tj�%M,�֙���R�Z0��h8ř�-���Pf9�X89nw�?{��?}��xT�~�*�Aճ׀I��1Їi�am�o�N̛�F�MI��$) ��RRE	b�0q*��d\��!Aڋ��ﹹ'�_��� �d��V�i*��i�w�uM��}�ذ{#�5ulxݪ�*c�J��m�X�����xT�x�J�WF]��B�v�m`�G�j������ذ��Y�6�v�;& mvM�pH)Yq��K�o(��8ci�p�
uWD�>5\�/km�ۑ��6^��� 7�<��2��Ӷ��n��ۼ�l�v�, ٱ�ۗ/ ��vS���n�[��fǅ�y���U�+��ʭ�Q�6��;�5I/ ���ug���8�������x���w&�}�'�u�
I+rYn�}�/ �6^�ݗ�6<��r�Kv�~�����ew)OgM�Q����4�,����@�ft��EH��Y��� �V�i���=x�{ odx�� wj���[T�(BV� ��ŀ���q`Se��*Ձ�hjЮݦ�X����q��l����g1�j�ݤ]�����:��f�}��P�oHT
���̘��;�L�C�i۶�m`Se������`�����6>Z�c�Z�H�(LcLB�Sɷq��e��I��)8���Եn(�m�6�z6�n�e�, �����;�:���'t��)1�vwm`�G��9�q#v���^��� ݔJƅ@�N�0�M����xT�x�{ odx�H$�|���x�9Ko�׀v\��� �on^ wj����;Vʴ%n���,z��Ϡl�۩'/�{��~�������"���U�`DV� *��U��
��_� �������DW��_�����U��
�DW�� *��U��
��D@U�"��� *� *��1AY&SY=��o
�ـhP��3'� an��@P)TIGѠt  t*�LI4�@P (�=�d  ���h(��   P   (@      �@�    h �h`4 4� �� �   �  �  (�@ 3��]�)�#@G��zi��4y��,�.�z�{�����P{�|��G�  7y��v�)K��.�;a�w��w}� _x:;o�������}���o}���  � >� ����ͨ*�{��{��}�����o@�xh�k�v {�@w }ǣ���#��� ����u:����\�=�{��`>a������_Cw���;�p{��0p �� P� �r�
�u�<ڃ��H=�0� )ǡ�7}��oOC���������|�=��w�x��v��*!\��@�`}�G������z;��|ػ���� x>��    ��)�/ �������r=i��.Ϡgc���Y�Ǡ��g�r}�p={��} �}N��w�{����C�lxl���;�k�  �  �
 
1���s��`�{�ڇ���K�:M�}�==)M���)����K��R���h mQB�R��f����  4��K;��J8�6S�4��P ͔���tѦv h
�[ ���h:9�ҍ4{��J)�g@ �2SmJJ�1 �تR����   4�j�S'�( �Oh�m)J�@  �Ѫ�%* �"B�*R��0x�R�����?�׿�Z����n� &\�-e˝_פ�����"
���"
��QE_�"
���**�QU?������������� SI,c I�hI���H���Bl����.'6jP�ILP� �;���I~HW�F$�X0�4X�I"U��2�T��Ia.%�q/���.�	��P�+*B�Y�#$*|�
�J�!
B�kJJȑ,�L2�GJŉmo��6I6l®<�G	4!d`P��p��5c@��Jf�=�:$0`���������v���.e�$i�.0�X�,��P.$��u�.��5 �~髐5$�	��dj������3���x�#�Jt
��hB�
�a$b�c
���1��"JJ��(���#k
������̘˄��Ja.�B�H�R$�)�[����k%�Vp�����RJu!H��B�.Z4�u��Cpc1ck	��2%Ιu.��/|_wy��^!3�w0��\�Ye����7�nɌ�+
ă��l��O����x��1�{٣��=H��]?���HB"p! �L�����`Յ��B�}���$���f�E�"� D# 	�@�n#��e�������Lv�@a7�����i���IR�4�F�3�T#�"i	 Ȅ��\�C3�0����:s��B�%�6�s��@*�0�`D��1"E�!�agi����Io��~�R%IR_�26D$�VC�0&���C3u4��{�3�35?f~�},�Ёԍ�T���[�1�W �cRX�/I�5Oҟ3�	La��J:�˞'/ZǠ��z�u�g����X4�D#4 �уR\ֲl���B��!\�pL�)�c�#py
h���m��d-0e���[��52��V�#F%MD(!��\+L�ˠ�p�$bB���
f�Ez�L	w�oi���O��S�i����@�3�p˪�oI9��|@���)O�Zi�J��Z���.B��8�$I#�R�8$
�.VZ��`$�I��4̦���bn-q%SL��׽�����B$CF�j7N�k{5�&�Ԋ`%k5��s\�N$��	FC�R3x�"B����� CVfR晚�ޱ����H��q,!�B�A.9tM�$LcI�:�@���}���!`Q��!R1"�k�d	Fl�!ll$�a���2�d>�q�Y4O�-%��
D�!�Y#R\4�� �U�P��B�b���B!B��$���#�HHp��c@�\!Lee	C%�\fY���B�������j�2�6��&/cI�����
E��J�
�J��
��[�2���@���m!�?: ]Ĥ#*¿$hF��D�)����6V\40�Bk4�s�7��.�yF0 ��0#eeHĕ��B�q�$%c��HYf&��
����|���z��'�TJ����JKt<O0v�it&����8��RBc�k!e�,l*q?���{�^,�$  IaKa:XHW|̉5
M�ےI)��a���П������k���h$�I�}1������!�C�$��d,�#�$�+d,�BL����(a�t� ໥Ć�݊�\�,&:\�7B�9�5�p�"�
�$J²�#$)Vy���;�^��$%����������M��]�d��C��B��RM30�p��0�o�7��gѦD�_|Ml��w��Uv]M�mozb{Ė�K��BK���¤�+
·G�$%7�xK����/B�N!s�t�@�K!����X@|��Oø$3ĺx�xJ�Ǜ�4.��%Ļ�s�h� ����I�����`D�a)��Jd)�����ϒ�3�����"u�=�B\�Bc`���̅��oMĺBF8h�7��?�n��Np�+��� G[f�۲��!� @��F�,m��i����"���b��7����#XQ�B�2D���`j A�~�#!L�42����B$ ��"T��h�$$	s���͓Xh�X �3rt��"�w*k&`J�|B�(K�.$��`Ȅ�!�`X`Ԥ�&GP$Ӕ3)�X,L�^.:�XK!a%:�):�f��5q��+·		�Y��\����VL��2��Z�s�.�!F��
1i�?@�� �2I �U q�WIƌ
� N~!q ��6���]A �j���$$H�aw�!��#d�!H�4�D�1�2����W\��V$"E�`�R0�f�	����1!9f��Hjfn\
V! ��4�h����op��3{�zwL%Ƅ)qṪk��d @ 	�@�88�:�Oĩ$�@/Ĺ��C �Hߝ���O�
Y���%q�>�i��LcЕ#L��D�B���A"F� ���@! ��"�1��	p�D���w>?�FX��p��	Cy�|~a�E�~���$$��cM�af��D��ǋK��t���z+Įᰔ��\P�i��S%�	�ɜ��Ls3@` ~�\��r�d����ߌ���.P�		%��BW��0ֿ��|���oXP�~���I���-J�m�g�܁��"՗d�5�A��62�#
����f�����ƥ �x�ZƐ)���?4�����L)b��% M���Ґ�����CY�jrw��[0�IV Mv3mHi�F'�C�A!���-H������D�bB�bJ��):�E�����&0��!�f��]������!~i�yB1�!��I�j	�D�D��Q�G�k)r���߫#����!i�����'��&�-X`	�S�@hI
B�B���H���ċ�,i#�� A�.���G$���+!h@��
��!p�W P�IB��al����II��HP �:�%��B��|�{�������}ܭ�j��CϺ���4V[��~u����}��3�2�)�ap���
*K�$�$
AjaFaRR���*i��C��N�k\rM@�R^��.Yem�Y#��S! @� ��	0�HA�`X�dI@�,�ȵ�I	a!�	�6;���Ƅ�?�5� Ln@�,��o$<7��	d8�0�B�fA�K�/C�%���<�d(Q�d#��i�����YͿ�a�=�o�5����|~���S�4IR,�Vђj~��~�.h�¦B������'d#w��@���+��)�\��Q�%����f�H˟���2����	p�=�
g�sy:�"IaHi��c0���@�F�@�
i�u��HR4���|KBbX�aaHW���&���?<��~aB1�܅0�!XP��%e�96�A� �b����|l�$�����6�e �1�`Hh�B)�s�����K�ٸ~E��_�pq�nU$B1d��r,�e �������X��5�DJa� D:��`!LM�8v�m��,��_s��(��R��ߞ�ܗ�&7�,�)e�pi����q�̆y�`��I���]�u�e�[7HDb4�����i�1jF�����~�\r�܃$'3[��������B%�SL*@�D+���BF�h!qHۦ�5
V�Z	X�ݻe	XB��.~d8ē�a��Z�[!2J��B�"B��B�*@�
A�+)F���wQw���.�}9���z�+��uÈ���&"S4l���&.�*I�}�}�s7��2f�acea�'�+	oRo?I9��$���Sg��χۤ�	a^%:���I� Bl��Ա�!#�B$"�%�c$$1+?2Je�\�iF�m�,a��a#Q��(`H�5J�.aP�Hȅ#D�*�@+�Ĉ@#�e�Ӛ�FB!�l�,jB6u�s����������O�3]�t���d�]����pv���$�	����%�BB��+
��D�
�k2)�# FƄb@�3�0Ϭ�7�q�5��%������I$B��$wRt�J�D$����!ݸ���\����{�г����
kp܃`$�&��4!Rqt���a��%1%�%#��RE)����"�b@`��*�I������aS����%7)-@�4��j�7�	��m!Y"��h8�c@���Q�X0-�*��`$��I
P��$i��%���]в�7Ϫ�������ڪ��&���ڥUU�`ڪ��UUUV������*�V�4�*�J�J� m�6嶭� *ꀪ�����UU��������ک���U���U�WiUQ���j�ee��v���Wd �'0@R�L��WUU�X�cu��tM��Z�n	�y�N6�� �lmJ�Ҭ�V�@5]�h��Ho4���{�h	�mO@���UUx���Gn0�JKJ�v�@�U��[i��;ED�t*�+�\��n�]�ٮݫ$Pq�eV(����Rb��WU����]N�G���_	�g:Z��U�
p =/&�LW@W�إ[j���+j�ꪭ�����61R�Uu�UmI�dnU��B�5�k���UR�[WR�A�-R��UUmV�]M�ڦյB�eP*��+=��V��[�HMvԠvpp�VյV�]Qu��`�J��[c�*E"�{�+Rll*��3�m�Gn�;\�囩�S	�F�k����)UV�UT�����h*�r�Ӳ���j|9����h�ڢ�#���L�
�����UUR��V��MWV��W!��BW������VV�V�v26�;gf���V�����Z�P h瘽(R
�R�i5ȼ��VBeU]R�Ő���!i&r��UUPJ�UUUU+�*�*�r�����zӵ��֬�
��J��x�ʵ!J�{J�G�H��ܵUJ�U[UT���
�p�n�un�m��5�F��k�x�j����U��n)j��v:@������j�j��Bj��ګ]!UUT�U]R��
��lCePUTUX��X�k���[���(8f����һK+U*W���������B������-*�"��ڪUU�	�
�[T뮖�ꦫ4�UT�UTT[UmU*�UUT�Ej�W�SrSkm��������(v�jh)�����v]W5TU��y�-���T�L���v��lR���
�
�G[P(���uR��	iPA��^�j
��-�����T9`*Uö���cSv�C���P��uJ��ԫ�\�'��uT��U*1uWU8xx�j���k�Y]���]UR�N�Y�%�fu�*��K�Uur�.�+mX�1m`-R�6�ޞ���UUJ�V��UU�UW:�f����W����`�V��v�Nܒ��T�+v��V�2 5P�_tq��Ь�[\�UUPU[@[tڽR��7�̭��j� �o�W��U9��ն�z�UV"��i�ҬU4jZ��rpT�Um�l�I;��+�Ҽ���%�΁:��Z�W��U�(��	�P�$�E�MM��Jj-�^Eez6�n���UW��}��G���0�k�r��6�x��U�Hm��T9��SR�US�ݽ�ӫ3u���	��AP�k��̭J�Լ��z�Z'�� q�.�[�pҲ�UT�J�@z�
�mUTO+uV�!5UV1�K�J�u:���mt��0b�A��
Rej���`%+R<�����Rjń�����m��SUUT �Uߕu��P�5C�5��1Բ�vr��*�ڪWj�5%�l�n1l;�ڪ�V��5UN2�0R�H\�T��*���^]����m;'?*ԫV�4�J�jj�yZ��k��iU�\�5\��ty��+U�UQF���]\�ye[�@R�Yj�b4�U�UP[2��v���R�ptq�V��q-v�+;-J����vun*��j�jꫪ�
���b�UVv�m�
C3U<�ZG5Z��
�ڪ�-*��+�偪�j�� �su�z�B��U�1<���m��K.�]mT��-Ut��@F���*�G+*�յR�UR6������U����j�Lj�*�^q�����̇<�n�4�?.�;���vۓ��{#H
��Ƕ.�;�݌mU��^���tUUB^e��()j���V��v�t��Uu�	�����dtª�A���siZ�fa�Z�6�d�l�Ꝫ����j�⪧�U�UJ��J����������
�UO+UUUUUUUUUUUU�kY��V�	y����\D���@Ҭ���&��J�p�(U@n�	��Z)yd%VA�R�^$�����.���#;M֑n�n
�N&�ʻ6��]�A�*ͨ
�*��nR�HEٺ�YV���J2�1��*�]UUUmUUPV�l�Ue�
�j��Kb@�n��Si^� zü���m�^Y����UPUU�UT����m![u�`*�[� ��ٽ��Uk�'m�pp��R��GK�쳢�Cm�Rkes[b��	��[<�ꪩvvs����C�V��/XrNP#۰ܙ3Mܴ��Z��-T�WYZ=��s�Ur����3
���48;F��]b�mt�vDN�J"���h���ɦ��8W��n���kYd��q�*�us"�s���-�cf�eR ���k����E�
�CaU��m̀(�4��䶞�]��j�V�`�\X&p[�[R�b��U���ت�^^�W+�� �-UK��Rlr���n�k�
��F��[i-�8���Ǟ4�=UJ�T�t��P�ەMp�SvM��PR��p�mp 5uS��[{j6
������Z�<ls  mR�UUu/-e���T��U����㞨�m�X :mP���`  �	�f�/UZ����H!UU[Z�U�^���mq*�!0q�6����ej�ڪ����}\��>�UVԜCB�mQD���yI25!6�UU��]ѳ$�R�b+��L*2�;0[UU+*�^R���UU����UU��UUAUv@��j�8�ڣ��UT�v.�j���������ꪪ����v�d� ��[l.�⪎
������T���m�jO���r�@U[J�l�皣`�m	�U*��nڠ�jy�T�[�᪷Tѐj�U��%����v�[3�[U�����  j�ڠ*��7P�ʮ�*��%H4<Ϟx�u���|���`:U��3mR��U�ۇ��8��ٗf������j��5J��1],P9@���c��S���ڪSITV�d�#nZ�ڕ٩IjU�Wm2�"����_z-R��uUPuTUU+��W@T6�m<�� �UU���v]γˤJ���mLY��*���)KN)U���V�R��4�H��ߓ�}UWR�uUT�˶3��卩yhmUUUV,RR�]�UR���� TUUY\ۂ����tp\���wa�
��&�.�M���i^j�jXM�n����P R�,�h�Yvj˰�+�� �v���e�]���P᮪U�8)e[��j�rN�F�UJ�U�-D�J�*���("�%tNԫl���u��r��\���0�U���V���[�ۗ�`���UUX�5\=Thv{5�T͇���ViUh)j�b�D6j]b�����X�i�:<	��.3fZicY$;�T�V�f��.�i^v�3�.pAQIe^W�k5W������V�T
�5Zt�iݍ���8�j��*���W���h����V]�Ep�s�*�ܫC��e"kq�*�@���ݸu�lq���v�f�x&�6C#��s�lz"ێ��Z�VUo*��=��S�vC6 ;`է:{i�kV�[��*ʷUUUR�+.�r;u��rm��ͳf<۠9�*��PV�%Z��
��u��Wh�6KrғNsPU�KVm<��
�+UW]mEWU*�!'��<��ZNw����*����ͭ��|�|�PR�UUUR��&F��)[pqŖ2*�R�ec���܋�^�Xt�`T�F^�Z�K05!�x��cZ��yY��n��Un�Z�-T�;mUFpo-gDYP�gc"Q+ ��E�v�k*��\O�Z������Z��T�c�j�*����YZU��v��0�L���R�T���Q������
U�����u��eD�V�
2:F���6�.W[MVԮi�Xj��u�T��h�	�FQ����X��U��mU˳t�U@�`��[+U+Z�ݕJՙ��y٪�ܻNQ�Aژ�X+��!5W:�U]	Ī����v�U,UU�e�ʪ����UUUUUUVҮ�UUU*�ն�v����ꀫh
���LUUT��UUU��� ^;�A8�����T9%-���A�BͲ���S���j�j��j�*�UU+}���UUUU@ZGe�m�PJ��; �UUUUKm�J�Sj���*��ꪪU�
ګj�I��U�*�\1Kr���j�UC��v�J�*�����Y���WR�;-U�UT�ʲ�y�*��d���ۖ'�[q���� k��f\bj��ʵUUU6���U�U]JK\���2���UUUUUUUUZ�������U�(8��Bj��
�-V�UUUUUTU@�4�����UUmUUT�U[<�U[UUU[UT��UU6��p&������ں�(RZ�V��ڕi]��	Iz���jڪ��*W����~���EUt�U]6��yy�����keZ���<S�J����D��MUT��-ۥ��eknPZ�  ��[e�媪�
���.�5Sm��^���`���A�����z��ka��\�N��f�J�PV�M��U�R�Q��W�y@٠'����Z�U�V�$�eꪪ����YVW��2�[Sj�M�UU*ܨ�h媪����Z���vZ��પ�������U��������������������*�V�����U��������*��j���ت�	>_��������������묣]@UXī)/UUUmPUuUUuӣ���Z��<5��b��f��33Zֵ�����*�M���v@��?�@?�����$D�E�uȿ��mj�?Q�t�E���V��j?�h�}�TEW@`,H�u�8p� �U1  !� ��0��q�buA�q)��?�*"��Ά
t?�AN~� s�? �p�#������(|DSb�!E"�dA���~PK�T>�5cڪ@C���G�ʪPT�|	�S��v�1<D���"���s� UWG�A���4�	߅A���tQ�JU� ����G���>�3���|�Q�	 �# 
�F
!��= 0"�hO���ߔ�@C�PD8 ]�0H`�P�S���U^�/ >衎İKZ��k�@���4����V������! ���~ ��AW� a���4AQW���Pv(�ʫE��X%dV�Z�V�*���m��9�R�������[n2����&"�v�v����f�Eg��!NZ��M2!�g5gm�4�n˺�2�;s.W�"��
�u�L���Q�˻I��=�j��#q���\���l�-+��V�S[6�;͐�r �Qם\��0B��ZkN�nۍk�Y�#�GD �J{4��S<s�N[i!ӳm�!$�Ob�p���ƃ��Ft�Li�ؕ�Kvɘj�fɹ$6�k5I�J���1�sJ%�}����M��]�<n��˟X�����%ns��s!�9Cv����q�{l֎3�ܮ�;"�i��.��UP7$v�����=clp��l��Pu�a.޸5m���&Y�U�@��,�5�� u:�v���!12胅صR���f�ڲ�Ҭ�+�VC�Z����[�A&(�a�G6�� Gcb���,�:l����Js7�׫m�h�G%4�� �A4"�p޴�ܥ�]�{h��0�3ƴ=��	
�M��nM;��*�/<]:�"�e��/Vh�@u#-�K�37h����tq� �v2v�4����M��ŕ�K�X��4��d1�5�@���p�퐦U��M�胬�n�����%��UAJ��%!'l��is����|���,���.s�.^�[ABa3&�K^�c�⅏Kl'a���q��n��΁�SN�v�d]q�9:����[!�����$
�esn7d����:(�v'��ƴ���w���>9����eZ�h�@�;^K�=I8#�X�lknej4�@i"q"\�8�O8q\�N�lj�l�vF�:�G6�����nƠ�d�U�F�R����VA�IrQ���,bt��A�tQmѫt�۫�����+UUI;���\�F���J+(p�#q�p�&�����D�������n��L<M�%�6�j�K�ѥl��4ԫUUU@)*Nd)��{�9��N���j�� ����O�~�hUA����~����=�����*%V(�K	�ڞ��'=��sU���]l�4E�9����ٴ�9�N[�L�ю��Vfdr7@CP�ڳ1Ih��P��.�0&�y,N�:%�v0�`�׮����m�[���^@��ʎS�ӣ��@.G��V]�"��J˳�ǚM9k��O ���S�\Ց)7n�	Z�a�yYV�.x��J6�������$#|{�[���=��&y��Ƚ����Br5P�F�D�I�bX��������� �	"}Ͼ�n	 ����`ODȖ%�����r%�bS�ϳ����]pMH�\t��N�����w�i�x�DȖ�}�Mı,K�ﹴ�Kı:g��D�K�)���g�ػK��D��t�t�K������Kı;���ӑ,K��wYq,K���w�iȖ%:Rw٥�~�u�J�[�秇Jt�X����iȖ%�btϻ����%�bw��۴�Kİo~�i7ıC��ζ*�L��J�������O�k��7ı,N��{v��bX����&�X�%�߻�m9ı)����>��/�:�[0.q����eb ���t�j-ٚRv��ԴT�Qˣc�fk!�4�P�ՉȖ%�b{���ӑ,K��w���Kı;���ӑ,K��f��q,Kļ'IӤ�B�V�p�ޗ��5����m��|P3A����M��J�*��↌E�)���w�,K���m9ı,O�N�R&�X�%����nӑ,K���.�!�����)�Y��n%�bX��w��r%�bX����"n%�bX��]��r%�bX7��4��bX�'�;;�a�]j��F����"X�%���wV&�X�%�ߵ�ݧ"X�%����I��%�NU͑�+�g*�U��ʙc�˻Xh�kV&�X�%�ߵ�ݧ"X�%����I��%�b^���iȖ%�bt�]Չ��%�byAG�|__k3W��Q��9��c[xc<n��1e��,��b�(Ƒ����c�Q-ٶ�%����ŉbX>���7ı,K߻�m9ı,N�k��7ı,N����9N��N�a����qv��j�<8�,K���[ND�,K�k�����%�bw�w�iȖ%�`�ϻt����ٝl�%�+%�2��K�,K���]��n%�bX��]��r%��N(A�UJ�$B! H�(b�����gݺMı,K���[ND�,e'{��g�]��<:S�8�;��۴�KİgݺMı,K���[ND�,K��wWI��%���b��nHR
�c�����4�gݺMı,K���[ND�,K��wWI��%�bw�w�iȖ%�)��߻dQb�c,�Z����a*��/�rG\=x��l����M�7;-�˶��h�k3WI��%�b^���iȖ%�bv}���7ı,N����9ı,��n�q,K���g{5��ZY����m9ı,Nϵ�]&��9"X��^��r%�bX?g}t��bX�%��w[ND�,K�N��K���%ՙLֵt��bX�'k��ND�,K�}ۤ�K��/��kiȖ%�bzw^��n%�bX����	٪�W�K��OGJt�JN��}�O,KĽ���iȖ%�bv}���7İ?|��! ,�������w}�ND�,K����K�$'��M6�������uIx;��	r�W��Rwt���;�Aה�䦮L���=�v�|�sI.'D��-��Rڶ�-۶��\w�N�/ 'v?$��߳޻m����m��A�.�$��	�K�	ݏ &�����r�Wai+��ۼ ���l� ٮ;�&�/ �tQJWv����M7��W*���=�OG�x�%��ǀw�	
T�L��:v��6k��	�K�	ݏ &�����U���y�PdSp��Er�GG-m�
��$^y��,gHЅ\��<j�!m
��=������u��$��:�d�ͳ�<���x�9+�C.B�1�x�gۭ�)o%��sg�t�\<�������W;c�1��8zٶ���.���"��	�բa�/W�՞���sȶ��=��!SX̦ZL�"C�5�C9n�������+�1�Hm�ҳZ�T�1�Ζ=S͎�a��t�\�y�q�6��� ��r�K���9k;��a&��g��M�ظN�Q�}�޼ ���l� �[/ ��Z���i7hT閝��ǟ�����x�O^5Ix�u%�LHt�M��:�^5Ix;��sB��-��v�7��s��_��^���	ݏ &��	�*Jʻ�aM��&� ��� ���l� �[/ �s��qz�v t豃���;�Ơ��wbB����Ƃ썞kn^Ͷ.)�7\�ܜ"�j�b���l��	�<ul�qkZK�~��m�u�O)$�mZ��k[�N���iç��@A��Ȗ� X�gڟ���ܓ��޻�N����Wf��{�*M�]X��{T��T��� M��mk��Mݠn����{��_��� =�� &�x��x��j��t�S�Zw���I���=x��նZ�qΓ�k�'�5e�lpDT]cc(�v
�(ط2��nsY��ɰ��|7c�;ղ�	�%�ݑ�sB���h�ݻm���x�����l� �h���Z�)�M�5Ix�dx]R)"l� �V��;W*J)]�CC(n��x�dx6G�w�e�T��v�(�Wj�\j�]�x6G�w�e�T��vG�dM�'�Z��D�Hհ�v=��6ݥԧ:���rod�۪�E��ϛ>���ƭ�uO^5Ix�dx6G�}*;*&ؐS���'x�%��U]�w�x��<�[/=�]��uAm��L�� ;���	�<�[/ ����.Ҩ�I]>$��dxz�^5Ix�J���9�b� ���'t7V�E�v��;ղ�s��G�_��y�� l"��mZui_wlSu�Ԗm��C-�R��B���y�m����ۊc��������T��vG�dxz�^ڹRR�Z@��:v��ݑ�v���7T��T��v�-��)q�ut;m��ޭ��MR^ }��\'%�e'wV&�7�w�e��K��#�&���>��n�.�5|I;�'T��vG�M��ܓ����rN"P��Ak�ӯI/}�;�y�p̐���*@��v�����]Y]Fx�̮X�V�g�m!��� (�B�l���`�1U��ZC\��k�_��Ck��o5�`̪m��!mj�;,X�bS��,֚3LM�.{��=�V�����┻fn�I���:�u���E��t��u[@d0���B��-���iYyVɈ��tL�4�V�XY4�r;8��R��U�g�ižr&p�
j�� �J%i�U�j͵�X� M;S���9�0r��8:���-;����&���;ղ�	�%�]Iv�BҢ���4�o ��+ �V��'T��vG�m��[����E�4� �V��'T���;���==�����,�66S���j�����	�e`��xj�IJ����)�t���#�&ɕ�w�e�T��w�,bP:h�M�.�!�+Qu�6�4nY]N�.L�H	Rn����$K�]�ccQCT��v��&���;ղ�	�%����W+�w�x��{����;�h��$��g{w��:!DB EX~�S�zgWe��ǀMٕ�}��n�SI�q4� �R^ w�<n̬�R^/�f�Fv�N��� �dx�e`�Ȱ	#��ԗiB�*�-17�I�+ ��"�$� �v<�ʾ��+nƬtYBtR�	����7��V�yf�4���v.%�w`^��t1�l��-����� �8`{��l��>�!�e�lE6S���Mp�W*�UWa�<�{���>��ܭhQ���D$�F�j�W���s�m������8mҡ`�>"l�����a�w��"B$&��F����!�,�O�\k1F(X��Bl�:��&�R������Bb;Wn�{
 �.	�������qM�M�sJh��!��!��2��N����X
~�!�I�~�1��1����@'��6"���B��
8�~~6?( ������.ͪ��W����� �9�{�b �`�`�`���o�b �`�`�`����f\̐��E$�k[y{���A�A�A�A�����A�A�A�A���M�<������ �{��lA�lll|��?��u4j���sF�A��������A���o��}`n�<}=��~����V�;Eoڿo�}8r
���*%�8�3.#�:a����M�*n���x�x���1o;;�߿��0���͙_��÷���={vK,�պv*��`{�����V��y`��}rZJm��m�o �+ ��"��]Ƚ����m�m\Bumզ�-2۬W9W�~��/z�~��u�)��!��f���nI�Q�eݍ;E>7i��n�/ �{�`�e`۩��tiUٶ��V��c���%��i��t[ď;R�h�<�a�kf\m.㲚,Ht�v�[w��ǀvI��}}�`�K�;͓�Iӫ�i��L��/ �����c�'.�l*�1�RE�X�R^��+ ;ݏ �I��wj;(I]��wgM`�2�����̬�� ��f�b�ƭӱU�n��������;{�,w\0����T���Q�uvb�n��;x�w�]�垳58�R<�=PjC�(gS��y�7��D�"W�$hk�',,m]v
�	aur.тA�RZjR���:l��]�_�&�5���.�hYQLK53KV#w\V0��7��j�<䱜�7]�*
�K�w��c�ݝhe��Y��Ch:kK�l���'��A�i��&���򵗉�'E���۶v��4��gZ��Q�쎱����:�-�)��b�N]��c;��-�<&�Al運��!��������,�� �v<_kj�!��Zl����`uIxۮ��x۳+ ��V�˻wH��i7xۮ��x۳+ ��K�>���DP�"���f w�����>���\0�d�TZ
(n�]M�n̬�;�޿��� w� w���n��Z)f�67l<�a���v�0�����f��@܊3;-+!0������-:���� �u� ;ݏ�+��+���g<�~m��M�w@Ӽ�����"���L�ul�^�j*Ԧ!6+��I�;��l�X��xw\0�v�('i���CM�l�X���� �v<_kj��(n�l����`_dXw\0�������ޫ���wm*�v7�+� `�`ݣ�!���X0R�-�V��\2�2̻��t�|v�w�'��+ &�x���\�U}a�^��W��x��:E;I&� &���˰������;�2��Wf�O{���V+m�I����$���n��T�[b�B?�r����+ =�y�ˮ�9j����L��:���L� ���z�{�xw��כ���� �&V���O?�'��N�/ �\��E~m7tSNSX�4���P-�˄����KjZ՜F����a��:y�y�|G\1��vO`߿8ݑ��K�9U\��<�`�x��4ίn�V����~�N�����&���ߖ=��0wc�Ur�Uvz��]ߙM�Z|�B�������p��\��$�x��xТ��˺i�+|m&������O< ���>��>m=�y���;W��X�Г�m$�0wc�� �� ���+��s������Q�K����$�b��;�=s����g���ϫh��B�,�-�='���6��ڳ]m��O~��vG�wc���='�4.�y�'H�(Kv�y�e��>矌 ��xݑ��;����N�v+�$���� M���U�~H��������>��ED�N�e.ZL��ߤ�����	��g�����/��;t���[�� wdx��?/����	���$���$� 9N}��\�5�����9Ւ⛵�����ыn�wJOb	�1��y^�3�p���yx#�X��EY��\m"����6N-X��λB�M+*��b��c����}�Qa�8}��uf�ZY���i�o>q��R��&l���rBb|qַ-k�b�3m�UN棶�p�X�x�� ��J	.�x*�[N�b	�ga�c�ٕ;4�)�ԝ>B����&J6M&�L�l�l��͜ϕ{�}.������0�(ff06y�v'�ݫM����p�	�?�Ϭ���=(��YV�j����M�ݓ+=ʪ�	=�=�v)/=�W9Wf����v�uI��u�{� ;�<=UʮU��{׀l����I1�.�f5W��;��t�6����������vL�r��˹'�9u��Ū�j�N�7�}��z��g��|$��� !Zm��v��i*J��X������笃�%��K�.�12ƺ��&���J��8�X��V�5�<�`�ǀ���������:/F�+d�tjh�����}�o���"tUhdh�˾I�{� �/z��p�r��ܯY~i7b||�V�=�}���W9��)�����<_kj�)�6	�j�x��x�?�#��]����Deߩh��ƒn��p�=r{�����;��I����N�BW�bi�rƌ*Ƴ��Y�ms�PY�єҬ�3)a�=.Xe]+�n�4�n� �y�vG�}�0��\�{�[m�/{�RA�duF����~�r��*�?E���߿e`w�w�$4.�k�L���(Kv��s޻�~��ٹ���*���?�(�$
�(<�ߧ�=���>~����}�{����wm��~�;�^�g� ��xݑ�z�Uʫ��z���z�Z��;�\���v<��s�{=����^ݎ�6�����Җ؄+&1�N�%���vL�؄Wfn�T�[���Ӻ{Ϩ�r��:	��=�v)/ ��Ur��I�z�6y+UE�)	n�|ɘo�Hs�� $�xݑ竗g���Z�V[�6S���g���v<?~�H��������o�|�'*R�%�m�Zfz�I>ｭ�;�;۹)�@�EB^4?(�;����>7$�{�����Yf�+m�vG�~���+���߯�O~���>��v��� u`�RV�n����U)��s3����E@�����{Thn�>mϡ�Ubwi��xvL� ������	�ߞ��vW�ұSTӤ$� �ɕ��r��$�x��xz���Ur���ב~�m��vR�� 7}���9w����6{�X���(ݦ�*|j��o�Us������ �~�xvL��ĒA���m���O%eL�e!-�o�R^�g��|�<��#�.�Uf�^�vDa�@��XF2!B0Y:�j-�b0�r a��Ì`D� �#1� �D!X1d"B$ �`�#b@$H��,��͑0D�R�0&��u�# FH�	�&b`E�#"� �0�3c���`A��$B��V$��1C��	����-% XA�-%��Q��il!��a1C
FXF$�A0m @���%��$��
F2���a1#$`B!�B�H��!�,��Rj�(��%*D�l(����\�[-������5�g��@������"�3o�ҧ4ld(sP���)�%��H��5��5lG� O�|t��$��$!�F�$b�����*R�V-�Ja,+$����I������c@��->���I, YbH��<.p�MH�X����� �,��փ�AI4A�D �&�F @�gߞ��Z�P�UT.f��ʬ�Y������SAC1]���NU&I�е&�Z僐7;"5�K��u8fR[�98ь�,m2��+�gӳlB���=��J��t]��ȫ=5C��-�ƺ�U��N�,a 6�U��v��+��s�����<��YIB��#V�¦юwE=8���(�C�v,m>)m�1���.kIS�X�U�.�*ک.��iqK,��������窺�4q(ghڵ���
ܮ�Ĝ��ڄ���VxuvM�gv�Ý�.oZj�.˓���z��,!a�625���݅&)l�΍a{A��	���%��$P!�P����W��[cY��Y�m;s�Dj]+]�*uǐ�g~�y���l��*�f�Z�DL���#���d-�q��^M�2���ḫӓ�h
PW��
�`���! N���c2gɖ��]&�;6a�N����6飡��ժ�KvMƸ�*�g�q�j%8�Q�f��X������ܜ�uil�d��Sh�5#*4f�U���+9��hr�x%�U�� �=C|�� }<�
\m�ȡvB�.l�Q�ULT��U�E=�-��^����R�(T���R�56��Z�j�V��4�<r�iF�� i�M�L�� �`�Y`����;�΅ⱋ���]�ccV-�0kh�d0��92 
���]�[n����.��㜣N�+��i鶼�(�{tZ^{��K���Ç`�0����HY�'dXd'm@��&�Hsk���YW�[:�#O4Ps��ѻ�@$������s�����l�%nQz8R�m���#����� n��g.�r�n�������pE�!Bj
�<L�e�UU��rP-�)[jM��uĨ��#i4j��e�»*�U8��Y��im��(.��ky-��*ܦ1�H�kf�f +/>jڬ�ڳ����u=��%a��gNZ�����ʵ!!�͏������l�1�kY�
4��.�����T����s��] 
��P��׏�ݵYb��h۴��e9z+��:�+B���r���4�T*83����Goj���:��������&��⭖�=��^��v�흖�,�c;��x�����x�'�s��8\�fY��Nrױ�f�6
��W
j�mMPR�Ž���X��ly�R!]`-��ƨ.��T�.�:j��M���Hd��T��kj���t��y�?ĖRr�nkrms�.���XƝ�uaН�\�^L�#��keQu��
Fl��߿{+ ;� wdxf�`��<0`�ܩKd����~̻�%�kZ@=�o��wd��>���vZ��10B�� wdxf�a�UUW䧿~��Oߞ����Z-�b��M�z��<`=� ����#�>�4|Q��T6�'m�vL�׻�?�6{� �c��[��خ�]&ʲڴ\k%MJT6��X���qm��Ge��jy�r��i���M� w�< ����8~KIpo��mm�����c�����ܒ~�������	 �"H ��vL� �dyꪫ�װ.��U�Wo���k �G� ��2�{#�����h����6��+n���+ 7�< ����\��L�v��z�ae�N�6�n�{#�����፾}���o��T��H�����L��e��7anm;��[WM���`Vƛ��ɽ�"�"�1S�+m�ݞxf�`wfW�U~�s�Oߞ�\?P~�Ҿ:\m�����s���ݞ���y��ܻ�������c���G%����s�7$��w���X+�jg���$�����o�>���&c����wN��R{������0%z��-�����YK�$�]��۴� }�L	�}ِ���V w��
q��7v����X����B�g����c���kXV�y��ݏRo�,�M$�v�o�;�~0��+ ;��_X��{h��i*����Ӥ�0��+=Wa7�xog�ۛ�~�<�yHAT��KV�o;�]�wc��w���wg���rJV$�X�![o�?-sߖ/��,����?�,P;]��ߵ�'[�w��c�:�6�o �͋ �W������� >�ǀIwR�;\�/�c�+)�m��]��48zxK,���nֶd�(!ɻ*V��N�n�_ݞ���ǀwc��7��zm���+�UTsD�m�w�z�;�� �Ｐ��+=˳��)y+N��|nݦ��<���,=wݞ����K��CM+|-[i��� ��2�������	�7�+���Cj���X�ٕ�Ur�}��vy��ȰWʾUU�*���r�ko�� ���C(���.���Ќ��A�Tv#c��Gs;K[�g�n��%�`�i�ݭ��ÎGr1 dÛ�T�"��[n��fey^m���:���Y�fb+.�e!fU�[�(::�J0��ĝ�[$vyNH���Z��q����g;Y�s�Cu���}�����63X��`�Ж���[��Nha
��ڭ�M���EPP4�Y����[��z�{T�B�̖{��t����1�P ���̆朼=���wT�w��o� }ݏ ��E������e`��I�Ac`�m� ��z�ͽ��ݞ���c��r�����;
m�l���9��3h�{RC��^p ��Y��׽L�H�Q��9�=�N��� �sל >��ljO�}�� zxUG'���E�-F�ﻗ� �S�޳�Ӿ�� ;�q� 9:>���04�G����f�GS�G��k:�ǋ�Y�Y�,� ��ۦ�㕫���߾ ;3�l ��2s�vf��� ;��� =2�z9Q-�d-�̀�fNsz��/-�fzsh� fg�8 };�o�KZ��`���-���*��s���`߻��?I��� 3��9����8�!R��-F���^p �w,�߮a� }ٛF��sy� �v�%����Y��\Ü ��6���ܼ��TL���5��n��;hٍ�6[�`ă���@sŚP���2̥�']V�-� 3��9��.3`�w/8 };�l ��wcS,rK+�nYNp�ˌ��JH}���ٞ�`~�Ü�)!邪9<�)P�4IY� ���� N��Z��\\���>�� �Om ;�k�X�*��ui	o8���Y�;s�8�fm gr�;[29Gj��v�f��{�8�fm ��� N� ?//g���,"t���4�2YH)nR���Jr]x�u�F �e�i�*ƌ���*2��;��F�32�ͩ�r@=���T�t�h�d�[$��`��y������sp���7���?k?~�p��v���p~ڛ 3.a�ԓ�/�� �{ל �]�����5`J�������8ܗ�� gs/8]{֖���|��9�uM��{c^��¨�;m9��.3`�̼��f�����8�Ik-^��U�l˱y^l+�քT%v�1א��H�CA��+l�^[�N��zk����KwV| ���� >36����<����d�f��kX�m���Ky��ͩ�ii-I�}� ̗�� gs/9�-kZRC�+g��v�m[KT��� ��6��������y����]0���$Te�8����N�ߙ� ��ל ��mM���s�)��#�%J�$� ��� <�Z���qN ���ݗݶ�h$�Py��l�r�f��D��J���3��Vp��]vΈ��Q��cX�@�C��k��7����8�e`��+�b�[0�	D�r�.2;X��b۝@$��,�m�p�I<�g9u�~����,�-�m�KH,�	�2�4!��	ص�d��`�ƶ]·T7gɨ$涣�Άr��EG�7!ઃ"i�k.�nC4d���;�`ز���1��ͼ�b�Y��#v�es�Wq��C0�k�U�h
G�����͂��--��rHJ v�-����jl ���� }ٛG��� ����jc�mI]�j��M��0�=�-I�f����8��ڛ�I��=�Ե�h7�Ӝ �K�l 33/8~ִ��3�S`�}� ��U��EF��$��ZҒ{��� :g���˘s�~ZK������� =���E�R�ꃒ�p㹵6 y$����|ܗ�� ff^pE�&��E����rv[�1�c�S+2]�X�Ol8����Ӟ��[CU�2�,��m-��l ̽Ü ��6��gr�KI%�����=�VU����� >�ͣIAz���dBI���i���ڡB!�B��!�e�$D0��!�b�	�S�D A\ E�DUy���߻m����9m�_~ڛ 3.a�{I-kZRC�yVz(��*R�$�� {��� >;�Sa�Zִ��kZKZ֭��_ߎp=/�l �gs��AZ���ݖ�ͩ�2��ݗ�<��������y����n r�Ձ*� 3.a� y%����~g ���8 ��� q��1��[x�E�_i,���t�d��3y�fbe�Q���S�t�ޑ�.�6a1UO��=/���3'8 ����%�}h��� ��U��$ti��J̀��9�ܸ�����rfѿ�~�Z���Z�?D��.���s�߯�v߾�{y˶0�0>Ů��������!�@��&� �ԡVK
�vQȌZ�0$��Ɨ1����&�3k����Hibn��Bh��Q:�q��d���ƴ���������9�� )�LLd��Bp	���hI�$]�pRB1$�"*�'�[�UO� Ѭb��UM�>~ �O��:]*�?�~P|	�{�gv]�h{��� d�L�e�ڭ�+��I��x� 3��F��̼��\w`|�o!B��$Td�8ܙ�l �ҟ{޿| ���� �op� v����n�zs��T[�r�5η$!��as-4B�\V��e,&�����/�ɜ�L��;�y�͏ �[/�s���=�{����߲���]�`��k 6lx��xŲ�������9��Y�+C��X�޼b�x~��IO����=��`�U2���V��5��s׀H���	6<�_T�`v]:BR�I���� �R^�yzy|߽��d�m�KZZK�b�'�P�J���IL����hLY��(ʸK���J����9�W|��<ohl#�y5�}���_6ے,E��U���޼�暦7M���+M`��`-��oT��lx�m�bBv��J�5�}#����=Wf��m�y`�7���ӪM6�0=UW5�׀'��� �c��&̫��.�S��n������������7ߟ� ީ/ ��v�����߶�XV X�W���F��%���	�V`��J�ڈ�\b ^u��+�ˁVC�l�[�#�[�J��Svp��!��	(�U���E 0*�Z��[���v$���Ž����dL۔�0�۬� ��s*ͦۻ����|��s�#"���y]�Q
�b���k�Al6r�	hkGq������ڎWH*�(��S.����{����s��7��b�����Wt�8��k��L=�2��G����%��q���Y���>K���i�[o�	����>��oT��ݏ �T���X��m��k �c�{��]��޼ �<��dY��W.��t��E���)Sf�����Ǉ��U~�+��R�{��7ߟ� �-]JBM
�bn������`lp��W9\���z��Qs�k��v�i���r�ʮWg���M�� wv< ޟw�"��L�ܩ]*�t��1j2̃sI�T ��Aк��t��5�ԂɎ�y��X�0�`wc�+��s��÷��l�q��ui�&�m��\��M��D`0 ��M*� �~��9ʮn��O����,��*˱S����ݏ ��"���W9\����n�z���H/
u|e���{��9�K}�����w�F���}���o�����$�+	d�m�lp�;�%�wc�;}�`�VZ�Gօ��4p��vwfs���ٹ䭢��箨��H"��ӧJ�xgKj��D�|��� ;ݏ �͋�U_Xw|�`�+֮��i��bn�����ذ�0���ʫ��T\�i7E�[�����_{ٹ'?w]�������KK���=ɿm��޻m�ˢy��(
�J�5�}�� �R^ wv<Ur�{�XvQt��,�Rm�ـn�/ �9W�y�߽�}�� �e;�p�����g2�`8��.�E����(�72
���#���o#�4l�ˊ>�ݏ ����U}a"�� �o�׸�.�:�0����z����l^��wc�;g6�BI�bM���8`j���*�ݞxܞX۷M[T��e�*bl��/��׀�� ��Ł��q� �Em��J�;.�bn����r�I���?ڤ� >|'ϫ���fa0e��Q���=�XC6!A����Fn�wa.�:x��>]�$�ے,��uIx��x�H��HT��]:k ���?~�H�~�x=�� �͋=UvweN�"�uM��f5{׀ݏ ��E�}�� �����v*uhi����� ��y`lp��U_����`�����v1�Sm��Ȱ���v{=9$��k�rI�ﻭ� v- �@ 	�@��b*>���?���e<�i�M�;v�v�_ �:ͥg���Č��F;j��%[[���vV�V/C]u��[7Z�E,c� @�b඗����=R�ScӶ��d��F���6��cCV�D�=�l��Ő�6Gm;�4�mi�߿��k�r���za-pn0��7a�JT��A��n-��v��앛50�U��R��-��b�U�ZU��$��:y'3��'l����>���klv:6�(�$ڱ �6&hS=��a�a�J�;��Z��)��$�5 �y�0�8`wc�;}�`wn� ڡڷJ�Sf���*��d��6�y`lp�Ur��j+�/X�����0d��>���8`�`D�U��˴����}���I��k�rN~�]����U�ߞ�ޣ�e�-SG��i��c��u� ;ݏ ��e�컁fZ�[C��#i�9�
�A��$�`�����/Gc̆�����I��y|��lȪ�z�� �v<�/�~�UW+�6~��}����H�F\9< ����ǧtJ��+es�U*����<�v8`�g�����悔�Q�tmV�m��3��c����z�vy�j�6ⴕ��B�ۼ�ʮU�}�0Ꞽ �v<s�����;%�G��պWJ��0��^���ݞ�S׀}��{�i>}k�̺R���ɢ��k��1�k��+&l�ny�!u�$�_X��Z�0��w����>��x�\0��m�#fd
�K��%{m���7����wT���p�UU�=(�e:T����H�� ��w�e������@�6X�G�������;��n�t�Z/�l�m�ف��{�<`c�}�%�~�UU�}� �mO`RH����]&��w��~��z���e`�`^�%�:N���Zfz�ZXM,�99���/�#����}�=)�`n\�W��:��v�
քcs}�����xݓ+ �V��>��x�����$�H�I� ��2�����ĉsߖ�{��E����4A�M1'X�v,��ܮq-��������w��dvݾ6S�um���r����z��O]�9���ܛ�|�Z��䟿cgre�%�A�M���0�o���$�U����@���ڶ^4�.��\�h�GQ�����h�����K�8\C�m�D �eT�V�h�,q�&�f���>�<w\0�\=��9��þ^�����ߒ��M�M�Ӭw\3�\���;#�v缰�fV~�r��vo6��)Z廻T����?ײ,?s�\���e`#�w���b����)�I��}S�Xw���7u��*�}�=x��]�զ�.�m`wfV��^�s���'{�u�'˂B-9�?3�{��:8��!&�T��)�C��S�R�Xiح5�(b��\6"�64���1]�T� ������Ns��PP�u��@� 2���� V	��#�5C�I��n�7������Ͳ�ج�7T�l����i6q�3;�ar�t�c�!�8�;.��dN�t�Y�U�=�����b��nJ5�Q�L<�x�4jzRb�l��B����c��]�"�p��%�snsU�	�l��g���u�Vt]R��(N�u�,j���,��T�\�;94�f��lŞ�B'��;���Ġ\K��u�.ؘ:�z�u�Є#B��%Sj��-��J-
&#�ݡV�:��<qYэ�x��;h��6��`\;�9� �#^�Sn̹���)����;sۚ0�g���Lr�V�Dcd6�OZ99ѰG��;k���قUa�]�<�n1vTXݍ�6a	�� �=�r��ۖuvqe�dll@�gY�O�AZ-��fX�&�l��]:h�H3���x����H�ƆS�UJKUU�Z��(N���sR�^���R�)��x��WaXH��dx	�:��ۛ#8��zi6}=:ӦAx�<������q׭s��l/����i�Z�N�m�N��*Z�7N�,Z]liu˲���-UV%�я6\��>c:vưhc���K��B�Y��,���#r��q�QZ*݊�dr��,�l*��[�=�ŭ�&��;pk���@n�̀'f��b_Y��ZA볡�vF7Rݚ4G4mu���-�-�7i�4�|�f�K(��Fy3eЍ����΋b]�Xw'e� Ę�C��P�c�� ����c�#eL���]/j�1��fv8�d�pDΩ�=M6�3��g�ۂP�G	j�T�k2���b�/W;.�nm8�[S��fpc1�f5I�4칚�
��=��q�Y%���`V�(�.�V�P���L��B�{C�Sb��sӢ�8�tg�:򩑪��^XƩx+f��3S��YW���ve!����C��
m]u�9ѭ�G+]Y�D�m��jڌ@HUUUUR��J�@\�T��j9�f�".�B�(�	Z C��� ��'��~Q����:@��+�I��:w��;�j	JomƋ5�EnH�Z���!q�$=t���B�e��<үNvZ���dZA�1�d1�
�:�H���%cr��<8��r;�����b�����M��uy���s������ʖQ녅���q��Vܠ���q�*��E�l�x0ul��5`θR6���P�n�m��Z)�ۀ�\��u͜�E[��J�z.�|0yj������}��ף�W�)����̯�C���18��ب�����^[�$��{_U�3�wt��:�=#�}ղ���~�s�?�{�����'�}��O�9Dy�*`ul�nlX�ٕ�l���Ur�R���~��;��2Sm���m��d��6k�ޭ��M�,t���;)��w�}6e`5� ޭ��l[/ �v�e�VQI����u�l�{�Ų��̬�|�+��t�S;٘csЗ�Ԙ�N*�I�q#�^+� �] 7?ԻWP��dR�d��߲{���>�_���U}a<�� �o��Z��Jm�ܝ�x��.ִ���s+ �-��w�e��p=r˿S��"�i������e���x�8`t��Bi���Su�v-��}ղ��p�>�̬u,��iۻ-�m��[/ �R^�ve`u��>O��C�<J�o3�X�g*c�,��!�t�ܮ:ܮwY��Nz��͆n�՛
�;*�Zw�K��ve`k��\�ú�� �P�wn�vSM�n̬�.�z?b��\س���J-����gm4� ����[/T�j������+ 7���]*bUmSI��l�o�,�+ �[/ �v���V��l\T�;�7�K�>�2�Ų���xޕ��
���6���rne�J;yu�i�\�y�p�1��ͭ���]�-�M�2�ۼ�+ �[/ ޭ��oT��}Җ�m+m��E�i�ٮ�j��^�� �l���g��)y�m��bm��=x�dX{��*�q-���X����>��HղժI�V�� ض^�ٕ�l���-�@$$��b��vn@�HK��5 
f�W=�S�����k�����m�����UnƫU�w�}6e`5� ޭ��l[/ 3�`Z�$�9X�KZ���iH��Q]�	�/]K3	t�%.�� (��o![hye;6Ӵ��'��N�/ ض^�ز�y�"�1�����w�MR^~���RG�/~�{���6-��Nn��J����NӼf�`M�+r�������޼yr�Qw(Ln�����}6�Vض^:��W*�UW5�׀wJP�-�Li��Ӭ�l�~���I������׻7$��>R$QC䳧I���q-\�A�3�[	�=���e��v�E�p��9"N$]�@wa� �q��L��B��XT+��i݌��<V�r�t���6Π�+/AI՞Fxp���{h��)�����3��p[��Ѽ �+�]x���r��1nز+���
m���%q���p����E��`X5Dvw;�r�N��rf�v+u��ƍ �]�\g�͎�:��J|�:t�ӧwG�=��Ѓb�ѕ�'�sl�c�8ō���&��.Nv�B]��j�BZ�X�:m�-	�h/z��Ȱ�ne~���s�U���� ؃���j������x�dX۷2��p�>�0���kIH�{��Ң8ݭV
�%�a�����;5�	�]���c�>ݢ�݅ZGH�L=ʪ����;��^�R^��YX��Ֆ���U�NӼ�Ix���_�vO,� ���	߼�������6q�x��Y������\d�����s��p<4+��z�yuش6ϛ~�/z��ne`�����x����b���t��o�}ͭ�ֵ�Ť�k�~@�9�>޻��9�w�rO�g{s����;�(xI�M�-�Ӭ �O<�^����e`��V(ݶՃ廴���UU�9��%Ｐ��������)c*ګ���i��6,�"���"��Bo�e�a�7[L�N�
�{��E���cuq��m��ԐunG����h1��������6<E����}�L�hX��)%��m���˿kZִ���޼ޏ���2��\�*�=��]ڲ��U�;M��f�`]s�^8�Kmb�p��P������nI9�<rTq-���i���/ �K�X���=Uʹ�=x��U��4�cB�� �e̬��<�� �� ��+T�irƭ'`2�Q\��f��T��y.3�pFi�34�vaQt�h��v��ƮӬ ����e�sb�>�V��mX�v�V��&��Ix�ذ�E��6<z��)c(�wo�N��Ȱ�E���"����I ��bL�>�,� ٱ�)/��9�r�Q�������{m���Y�!	ʑ%��m�������������}$YXf>M��at�UX�9����6����]�h�nQ���PZ)LD+t��&%lI���o �Ix��}$YX&ǀNJ���;L;N�	5� �K�X&ǀI��]��V�X�)�7i��z���lxz��yO^�)��7�0�C��4+���� $��	��$[/ܮr��_���H�b�m7v��&�"�x�~���}~��7$������),���Z.����3��Ɣ�����N�Ab�i1� b:+�i,ۥ؝�K���C��,t#��n��\���8;;Kн���
�\bU'�<X���&Uݶ���M�lԃ� �hm-�lu��Cg+�FKlnm1��w4�
%�&��	�����i&%��-
�B;�f�@�9P�����Pf�fcB.��їabB��ۙc�"d�We�Y�դ�kZ��q��BY�P�͡*�kĶ-�2� ���(1,n����!��H��b[�3D�M^\߀n��.e`������ҵMQHab�&`vE�����o��d������{��{Ɏ�h%J�`Ӭ ��<uIxf�`vE��J����Z6 ���x��Ų��"���9w7�x�����5b`��I�ۛ�dYX����� ��u�k�E_�xb-V;J��aT��X�9�L�;^w[v����Z����$�#TJ�bT�o�l��e`� �0�ذ� �ۤ�v5i:��w[��?��M
|�@�����w�z��"��'iV�6�w`�n�m�{"�%͋Us���Ｒ�ޞx�Q����-��ZM`�ŀ}�s+ $��=�W*�W�� ��Wj����E���.e`��O?�����$[/ ���,�\��L^��[HϱV��f��[��4ٹ�W�Pf�3��wF�
4�)��j�@�}���Ix�e��Us���X��껤�'H-��o ���U\��<�� ��+ 7�<jA��Ӥ�>&$̒w���rN}�ݛ�
�"�����D�?%�`&/ۉ*ؔ4�R��X�J���2Z��Q�O�P�
��P�)2����e��LM��Hk}7�ᣥ���s0#@�Y,@��"�D��`b����$�dDC��͟�TҎ��9���!��JTu��<�����U�-��"�v��~�?s�}��v���~xŲ�	��7�0�n��$��j�:�	6<�<��=�=x�.e`{elv��ˍn��V<�����X�p����S�����ƳDe�]�Pz�e|�����	��;��W��=��H����i�.�v�k �l��-� $���"�7tr�V���L��Wi�ݖ�lxܑ`��;6��gN����u���IxnlXO�|B �	Яȿ'�2�k �^�u,�c)�*���x�%���`��X�c�6�n�ۦf���}���f9Yo&l6���7%�F��M���M4�lgk�Pc�*�@}���`��X�c�6)/ �T�{D��'hI5��� 6lx�%�sb��]�A����+Wv$�� OO<nH���`�#�7����66���դ��6� ض^ we��~���z��&�����)$k �6, �eǀ�<nH��/¦Q@�� j�QGLE
X�T`�Aa� �
�� !j�F���P VQ`X�T �@"� �e���d�5&k3�	�LN����s�SkV9vDtW#�[I���ki6���� ��!��
\��2�D���f�F�\Xyer�ζ6�ɶ���8fF͵�B �3k�jg���1�<�T<�m^1�@�k�Ɍ+�0��4�;p�=��[��jv=��x,.	���e�B��v�e�4��bȻc)+5��4.b�ͦԛ@�V�Oztq���`���,\Hf�����lj��td��hZF�%���R+r�a�2*�S.�Qi��>�q�� ے/}a�=��o��]�uV�Ҷ�vG�m�7fVݍK�6���	H)��U�;M�{"�$ٕ��ʫ�<ׯ =��vT��"Ҧ�t�n�k �fV���lxܑ`*�6�)m��ZM7Xv5/ 6lx�Ȱ�2�	p���'v�X��U����P�Y� �uл�+/n���5�/�y�\��ae6�}���o�dX͙^��}a'���i��66j٦��kZܓ���7�6�`� ����}�ﲰHׯ 7�<uQ��M�h�|-�M�n̬����v{}�K������MU�L��ui���W�ؽx=<��"��~��Հo��:�i�I� I����I�+ �ƥ�^����:t�iS�l�t���"��v�hz�����B1D1��V��]��-��@���6)/ �fVݍK���<��=c�Z�ӫN�-��$ٕ�wcR�M� ��%R�ҥ-5e"�i��7cR�M�UO���Ȱ	�2���&��t�]�5m;��߽<�	s�X�2��Լ{Hڸ�m��v�j�6���`�\����W�I�x7c�=]眻7��m�=v]ͤ��Y�ZΕ���#�ګ�1p%f�f,�~K�J�˲�Pz�����~���wc�x7c�6�E�K޴b�؜��
�Z����L7�h���.{� �fV�h�(Wui�&��5�lxodX{��߽=��l^�,U�R�*vʴ	�i�od[�w�wf䟾�������B",�
��بsW5�nI�?Y�U�wi���	6e`�\��{��zy���`�U\�9QB+E�v6�|�&x�>�({e�s��n��$�Qe`N��Y5"�ME#-FIe����~��m�v<��/��9Ϭ=��i�V�&��+��m[X&ǀm� ��+ ��2o5�ߖ���~�k� H�&�I+o��ߖ���[z���<uQ���Bj����n��X� vl�o�I#=}�m�ޱ�ɫ"��+�uK� &�x�%��e`���C��o��[��ځ��X[��h�mθI�2��&n.�U:�p��Z-��yl�R�kDnՐ���WL$�QX�M�hqh���/O���/:�U��e�ԍ�ն�j�r�n�9���P�!��쒤e*]{d��5r:Ռu����HJLF�cmB�.�/l3 �ۄ1brN�N1�ji\�E�n
Շe���ɷMz���Tk�?w�ߖ���m��0��e�S5���t��4ÔlVq���ۍu�d�׮��N��C޶�e+e�&�zy��K�6l��7Q"�%_ap����T�u�v)/ �fV����+?W�H��~����4�m��{�V��ŀ}�b�o�3���S]Q2=FYe�m�IW+�����X���b���̬�5ܴ6��:VYm���&Vے,{�+ �D� ݌�H�E�v���;W�����.�e �mf�"��HX����n鎭4!����N�u�v� ����7T��	�2��
V�����ݤ��'d��T�7Q"�;�2�ܑ`��+t����U�;V�`��`�X~���{� �Oe`�WV�
�-:�l�����+ ��ٳ+ �D� �}�V%bo�ջn�ܑ`ݙX�$X�L��\��{��|���6��2�5� ����M�F&ˆb��(l��w����k��m�U���擾��{�V؉��+ ���T����Q�E��u�n�E�ܻ;�{+ ����ݙXzk�hv��H��S5��s����?^�����SdT�Ȇ0>��� s��Z�͛�~�'�����>K��ꋇ��g��'wt��^��6{+ �D� �l��;�6���N���ݤ��7�2�UW�{ߗ@�����v� ;�r�D5v��J��%�ةe:�m.ݴhlO(E�T���i����nƭҫ|e�;V�`��`M�Xb���W>��{+ �J����Ӫv�hM`l�Y���s�vo��x��u,U�X�Z\t����;��n����+�Wr#�X}�e`9,r�V�ڦ��-��7ve`��d���vnM�GpL�Ȅ*,#0H	��{�߽w$��y���-���u,�&Vؤ�wskm��c���MRA���R=^��N)z��F1���w���t������I�O.��-�5�}$��;��n����#�X�@��U�۱�7m:�;��n���7Q"�>�e`�d��V>ݦ� �ٕ�n�E�꫾���������V�:Ak�,v&���r��r3�X�������{������A0�(FY6��fmm���<wfV��ŀ]e�\\��9T� :7�CL��R1�f�E��#F2ڲi6MCu�Q����D?A���p:�qF(@Ȅ L��b���$V��4���1��HL� �p��l@�wI�\����BĬ�8G�F���B#@�b�&(ri $H�?����h�B��\�J ��iH)6���(j���&���#��������|����M/H�����0i�HGR�����;$���T�H�Hww3�C�R�}���TUX�TSJ��Q�ܴ%=+���Zl���`}(su�tR��:`�v��Þ�@s�p��ű;xͩ�8�0�݂�F&hZ6ik�i�2�H���](g��7.�A�ق[v�/`.�l�1g7l,���5�, R����6JPf��A�`h3T������m@3�9��(9�3��C��c<�N#�F\ssH���RP�C��lL�mD�݀3��j�kr3���P�G ��ۥ�fc�6ٸ�Ӄ�m��a+�2�Qvp;�#N�<�OF��q���	��d֧9a(�3�8��f��g�h��֛�zJ��Ѷ��c[��-�bc.GV�V�VE̬d��hh�\��D�N��5����sƻ,�lڍƎ�૥U+CB�w��7 �V�V�Lv�U�UA9�ƨ���\y���J�D�)Wu̙ �n��!�	ư���D����c�3s���]�3�QÎ���h�N:�p�:A\����D����ĘɌ4n{��ԻCm�Wm''�cۅ��e4!�ܙB�M�ӣ��i�2i�h�1���c�4=Y�v`÷@ƣ;
�3�%�s]�k����b��4� �5�AU*�]�
x��B�����H!�f;�������O(;Ȏt��Q�Z�֨Z�έ�����#8U���ˁnLQ� ���Nmj�L��f����J�*�i�9�a���������1��q(Fe9j�x�`.�ӱ��4�.vR:���,�:�u/:FH�u��49��A����Xt��լ�J:ղt�������J����꒛Q�%�t�TY[��cf���1[��ݲ��7 
�HG!Fg��w[=f��۪�inR�]���Z�����Yn`�Y�Vy2+�v��Dڬ�ZU甝��G��\	�[�na�ʴRk5��Ӹ�CeB�@SUUUUUP
�*��S���E�f���WZ�Z��qw�b~v�ЉQ�hAX	Q���8%C(O���Xo���lo0m6�5,ٳmB�^c�Ws�'e�r�%�g<Ѵh�4��ݝ�t�}��p2���*�,ژ�KP���;h���=�9�$���g���*�Lu�5�kD���hw��X6nE��LJsh+�3,fn�.�.�mY�N���I��Q[DLn�h)��#��30!+��0�W���R��VR�KR��85�йN,�WV��֣M���6�_^�K�Ͱ]��C���c����.�Ub�mnz$/"���.Ղ��B��
k�y��V}�lx�̬uK���r��Xw��V��߂��i��n���7T���L� �#�;�A���+�V[M7X�$X�L�=U˳}�<I��5��[�"�lM`z������ �{� �ٕ�n�E�oQ�j+�I�v����`d� �r����D{� ��+ �r��W�<ƛum7|�L�l�ma��@�8��pX6[�9�O%�",�uy���ZuN�����o�='���H���^����{� ��yZlZ����7Q"ϫ
���e`͏ ��mm��u�����m�ff� vH�ݙX�$X��.U��||t��`d� �ٕ�n�E�}$��6rX唭��t��m�wfV�����v{�X�#�	�ۍ�y�O�i�灴iZ��v��Sc:��ikf��2��%Уkݫ+%
�ѓB��=�#�X�&V vH��̬�5����hE�&��L� ��ݙX�$X��j�-&�o�ݴ� ;$x�̬��
��S�U&�,wfV�Tj�R�wc���I����\�I� ���>�e`d� ۚEi�]���bn��H�	�2��G�Mٕ�wM�^]�&��wM����`��q��:�� � }E�[�Pf]��t�*�eYi�+E�&���X�#�7ve`��`���E�B��6� ;$y�$���$G���L�g%��:i:\c���ٕ�n�E�}�e`d� ����Q�N�i�� �D� �d���jUs�U}$黻��}}O �����b��]Z�>�2�d� ����7T��	{I�}�xC2�mR�,�Ų�{���!Q�#e,2��Q7� ����&tE�[�B� 6H�ݙX�$X�&V�U�Z�
���Zi&��ٕ�n�E�}�e`d�=Wd�B�m�WE�0�զ� ���>�2��9\�7���$���o��VF�K���G,�~>��Ű���ݙX��\����
"�ܻVS��m� vH�ݙX�$�m�[m�w�IknA,�9�82;MC\qa㭄�[���nc9�ܰ�r���-�8=F&0=�E]feT���1DYĽ[[�H�qȼlf9�OW\�m��X�͉�cr%S�*��r\(J�0mc�P�g��_)cp�q<W3�ۓ��y��.��v�Q�F.�M�ZK����Q�Nm2��ӳnP-�L�@���:N�{��̹����y�[��a�J�
W����)e8�����%c54ҏjg�5:\b��@���u,vL� ���A���`S��i��7Q"�>�e`vG�wvegꪻ&�����,����{�Xݑ�wc�;��`���Whv���u�� n�xu,�&V�U�Z���i��x����H���Xݑ��W9U<{«_[�e��X��v��$ҁ�UG�:�3H�&tg����j�9��͖�j��E��M��{� �I��� n�x�J�_-;)њ�5��s����X��� W������+�ʥ�� 7�<���[J�R-!�ӻn��#�͏]�G��	��V!R�*�V˶�卦��c�;��`�2��#�>��
�D�㫱�i���;&V wdx7c�%�v�]�Y�Z��+�;O�ʖN\g�n�C����u�/�욗Q����S;�>�����d� &�x�$X�+lR�Um���[�� ;$x7c�7Q"�'d��;��KT�;-��I6�nǹ'�d�sr� Vh*,���E$_�C�P*���=���N{���;{����	��Ai�uK� �fV l��͏ �����*ӱН���fV l��fǀn��x�zS�}h�2����Mi#��v�Hn�:P�%�4n��m�]�ٜ�,f��&��� ���fǀn��`�2�	Ҷ�*Ֆ��W�;m�fǟUٺ��{&V wu0>� ����㰱Ri��R%�od��͏ ;6<�5���UmPӶ�=\�_}�}X�O< ���;9��U8�_� ޢ��-�n����j۬ �lx����n,{&V��M=���XАu�yM3�	vHz|��f�6af�����̻�VQ��l1t�=s�W���>��� �fV }$x��dt�he]�M��n,M�X���M� �����Wi�Ln���X�2��������6Qr����۬ �lx7c�7V�X�XҶ�*Ֆ��W�v�X7c�;�.,vL�o�, �UI�̟Ī�p���rÝu�.8Ex�q�0̓-���CgA���"�,��X�kl�����L%6��ľ��]���:J[���d6��X`Ŝ)�6w�N�;Ctpv�kY�5��SgVVا*p��"�-]t���3����������SB�
 ��!��\�%�WXA���ܛm�j�� �;L��s@�ZV�Nf�q��b� ��0��㤓����9�߈��1\�ùW��üs���ܚ!��g��2g%�[)�%�2'ln�6�]̲�f��7���od��6�"�����x|Gg���`�b-�m`�2��Ȱnǀw�\Y�W+�g�,^��RX��m�/}�lxz�ŀI�+ ���KJ�N��n�M`�ީq`l��6�"�6�K#�hC(�i��R��===�|��� l����DI�ҷe��e4�V�7j�-��ġ��oAzw�3�f���ɦqIdf��sGt[�m`6e`}�`�ީq`��v�Zn�t�wm����7�)�1"D?tl@�}��<z���7�eg��T%��Rb����v�X��xz�ŀod��6�"�',+�ȓ\t��I��=W��~X�{+ �� ;6<�k��IS�hE��{&V�� vlxz�ŀ{�[=�v/	 �2�&�n�����ei�)pp�v���V÷U�����C<��biq��ݷ_/}��ީq`6e`uV�t��Ӳ���L��ީq`6e`ղ����j��Qb.�x�R��6lٹL���~�H�h���r/�B$B$FM�f2$�J��#g��&��:ܣ� "h�GHw�m�J�� m�iH�)� @���� �@܈p��c��4��ڪU�@.��O���G��&���!���
�x7�}����<em59j��e1����'d��7T��v<�R%�l���UiS�ӻn��%�ݏ �T����fmm��f&nn)\,���׳�]a^wl�l�Yp��b���OoLQ�s���Ǝ�J����i:\V�w����w�\X�_�U���?�a[9��Ac��xz�Ş�]���X�?&ǀ}vA�I'v���ݵ�I�+ �ɕ�6<�R��7���m2����۬\�{��	��w�\X\�=�TT�"�}>z*?_f�7$�p�uL��I�EZe�u�6<�R��6lŶ�~���m�0&)d*U�v^vɩ�h8�b��/.���%k��^Mv��ݸ�:� �2�v��;�.,{&V��+ ;6<em58�T�)�Н�k �ɕ��&���I�n�y���<(�=j��aN�N��7�~0nǇ��W�� ���XҶ�*�մ���n�0nǀw�\X�X�8`���TM�:���i��R��$ٕ�od��	6<꬯��Q�*��$�ӻ�=���ML�E����"␳�#M�j�M��F�a�r4ȍ������VI�����l�һ;g�Ƙ,�=6v:�xywm���l@te3U/9�����`b)D��؁��tn�-#�`�7a�-��:3��۔�Y�3����!�vʘP[k���0���X-�{�bֽ]Bf�pP͍�F�:��5��zk��V��rspWnW l��T�%N�o���싏��iv'��h�:���Hh����<�[�-�7]����%v.�MEvhD�v�f�+ �ɕ�6<�R��7����Bi��۬{&V l���K� ٳ+ ������ �4U�Wm� l���K� ٳ+ �ɕ�m��ڱQi�X��x�ʽ����=��V��7c�6V�J�&�ct'n��'d��7�� &�xz�ŀl�ڲ�%V���C��WL��&�^A�n'�0c��d.� �0�b�\��m�Zj�T�wm���7c�>ꋹ�U�O}�lܓ݇n���Vk3F:�i�7cϪ�U�r��������n��X�8`����M�;6��>�,vL�?Urﾏ� zO<�;G��U��;-�m�k�J~�߾[m���� &�xuj� �Em��ջ���m��� ���ժ,{'���I��썮u�rD.h��W;i�i��C�`+L6̶\Li����>�rzzz�kV&��n����y�ժ,�+ �k��4.'n�Qi�X��xuj�?r��Wgg���w�z����r����g���a�R&Ak��?y<�s��n��N"�>?~��o[�s���l��]J�I5Bӻn�	ղ�nǀv-Q`�e`��w8'Wl���+n�nǀ~��9�V������V:�^������Ik��O�U�.fe��;�� ���9y�-�B��B`"�PÝ��򯎐�5���M�����,M�X��x&ǀw�w.��e��X��M`l���s���;��`�<���?�����Z�V�&�4�`�~0�c�;{�<{&V�Uo%��T����w����RS��<_��<{&V���W9�Wٯ엀K���wJ�SZo ����L��^ wv<�l��-q:t;�`���*#���K����)��e�@�e����zx���ui���1���v{�X�l� ��xo�#�6Qu*�$�����;ղ�����܏ ��+ ��������0nǀv�r<?s�_�/߽�+ ���J����5�­�m��ۑ�l��;�p��w�O<t��ut�-�j�'I7�Nɕ�{���R~������v����j��s��
@V��D��w<e�2~���b�=`�\���F�Dr�kV������,Eu�;��w#;g�3l	u"�]�	k�u(�m:8j�&{�Y�`sr��+r��;Ɲ�+�4�L�v6켪;!�n�R����J�3i!�:dtmqJ����2�3��_��lkr��� uF�,{pH�@�6�E���-���������9�km��0,k�����>t�:O{о~)ݺn�u�Z��a�H��G�Z;O��KзI=Bވ��3�m�	hIl�"���v<�ۑ��e`�S����E�Pݍ� &�xo�#�'d��;ղ��ڻ#)ݪi�E�-7�v�r<o�ޭ��M� ����,�E!0b�� }�ޭ��nǁ�W�o�x�.�V�&�`�M�_v, �lxo����~����}tمe��a|6�T��k�M��
��fQ��t5��U�17&^.2f��6:k��y�}�� >ݏ����Xj���¶Sac��xo���k����U�s��܏ ��ŀnǟ�f����e��X�զ��y�_v, �v<�W�`���Q;Wm2��ݶ��� }�ޫذ=W}�� ��^���E�P�$���c�;�{ }���b�=ʪ�T��R�_[��2tsR��6-�iQ��Ҹ�k �����)/&��lR��m��7��h搭._`}���`۱�_v.��v&���
,�;8���X��`e��X�̻m��3&��~򘠼�#�5e����>�wٹ$�~� "8�T`�7Ϫ�r�f�ŀ}�K�;Z0�5e�N������c�;�r,�[/�~�(�,j����6��X��ޫ�`�U��Wc������nǀm֟'�j!r��G]�6�q����tBc>І�ݺ���.tҎY*.�b�i��V�Xڶ^��ŀnǀw��X�+j��4��>*e�xov,�ʻ��MW�,�݋?UUU]��׸�7t�m7I���y�j$X׻�݋ ے�#�|T۲�vZo�r�������v�b��\��r�ꪮr�\�T䪬�W��{�,p��i�Ę'ck >ݏ ��b��c�;�r,��I���hц��/*���#mf,�%�$a�-ر�!�If��2����7�v��`۱���ʯ�@o�����eڻh�W�Bm`۱����ŀv�b�>���n�'lv:m7�oU�X׻��ܞX�<��)B+v�i��)�m��݋ ��ŀnǀoUȰ���ˍ���>*wm��� }��W"�9~���$C �mP�BH1،�(?��~��� �"��"F,��z-4@FBD����	���F�DGF�qC��$Y�D�<@[H �0C`@)B�T�(�!"$!$��$`�#��d��U�R�BH?�~(i5'�BX��_��0� `��a��<v Qq	8DLT��B���`B1�I��
��.���a�H�N��V�F0���`BHI!1��l��^C�-� �"H��B!!��"E�Ɨ����XF�'�3�H�=V�fXIi#��ӌ1�)Sj !Ċ k����[�ֵ�kUUXk�2ْ����%K[qE*��^-2���+��W�"�"�f�ݳ�5C�L�*rKWK���F1+!kbU<�q���i�֎6�8�ppIj=B(���jmtQ+q�	��<�cc�1�7�b$
������ņSYVӰ1�3��uc=�y&���F7lh��ɷj]d�<ںf'8��ø��B9]����������*G(�Z���Q-�m��T��c��v�Dv��q���J�ۅ�ݬp�R�qu�K�Z6#g���r!�^m�m�e�YiݬT�3�i(Xsт�<���K�s��/U1i�a^X�C�ɕW�uiK���Eóg��*�ӆ�S.���5�h�\O;ex}nz�;P��k=Nݎ�Z�v69Wsdq�
uԜTE8n��ˀ�mR� ~Ͼ��c�2��� ??o����A#ѝ�.��J��Ѵ�C�d�k@_|E��o��ܖ����;gs��_mNtL$c�<�Iŝu�U�**Q�� ]�#U��	�v�d��b�� 4k3ϭ�l���m,��IӦN�f��`�i\F ���S0t�nQRlƂ�h�i�{r::eA�FG*�`���:��lM��ޅɘ7\mb6��dˠ���%6�m��K�$���R�N��Kf]�Bv�d��f�D�'MF��5�Χ���	MK	:����	��Q���T�p����sa��V\����FA�s�Z��SX��hF�-
Jآ�=[zC/j��I��s\�a�>�Ӱ�H��G�c3ˋ�'&*M�g�\"�j�(����G/R���]v��j�Kl�\�SF%)(}}��SPݑa�&s���e����޹xQ���yj�Э�	4MX�83h����2�.�&�\�up��0g��=�NY#7��������l��US$m*�R3e�����d֌���� �գ�����]tQ�S2�M����jM�Ɋ�`C���5TOUUUUUT�J�mհ �=��tYi��!��"�N� |*��!�� yء���>C��W��?`��7>�-���5$������o�����˞�Q�	�eґ����;� ]n;[պ�L����5��a�x�	�9x���[Fœ�HF���m�ѻkT�'�Wm��`W@�;hӚ�k���8�v��7�*�2]lm� acX�]��!6�A�3��]g��ܼ�z�,��<r��p��t-ݚ��v͑i��X63YN�tvke�&D�T���kIh֒��Js��Z9H�A��{$&��w0�<;���֤�.`�4�?���'���]`�߀?|������`^�Xov,nJ,���mv��xډ��ŀv�b��c��Z֐>�aO 4J=I[�%�m�fy`^�X��x�^ŀIKiY�ۡ�j�N��v, �v<z�b�>ղ��InREۢ�S㡶����Ur���_ا� ��b�>�j?��-����Ÿ�m�==\�b�'c���v�Em��{lѭ��I��R$��ˀoU�Xڶ^��b��c�>�TǖJ��G��Ͷ���7u��/=-z"dU� �����������^ŀ}ev�\������_v, �v<�W�`j�xuT��+�[��$���c�;�{ }���g�/��7v1�l����;�{ޭ��}{�`ݑ�m�d�$���d��-MI`j�;dmm�6�0j�U 4f�	����7 ��k �V��>��X�d~��7U�M���1A�8�+�r�$��|;ܛ�l�����'~��f䟿}���Am��zߩR`��O������꽙��Bl��"C����^�g��/��\���M��r,�݋ ��ŀvG�}�Jm�t7B)�m����Ry|��<z�E�wc.��*\c.պT5 ��0[���A,J�W�0vͷT�u��F�y�9DR�Z4R�Ͷ�>�O�\zC�"X��}�m9ı,O����iȖ%�b}�w�iȖ%�bw�,���fi�њֳiȖ%�b_�����Kı;����ND�,K�뾻ND�,K��}�ND�,K��Io��uM�B]Yu�m9ı,N���fӑ,K������Kı>��ٴ�Kı/��m9ı,O�;f�cl˧S5&��k6��bY�(@ȝ�}��ND�,K��fӑ,KĿ�ﵴ�K����D�AT���C�T���?}ۿfӑ,K�����������gy��ҝ)ҝ>��ٴ�Kı/��m9ı,N���fӑ,K���wٴ�Kı�>���߁�p\��Q#�YX��h�M��`]�ū����˺y�bz���gc=y�ֵ��"X�%�}�kiȖ%�b{���m9ı,O��}�ND�,K��{[ND�,K��x�5d�5&��m9ı,OwW�ͧ!��G"dK����iȖ%�bw;���r%�b��}��.=!�Hz_u�}�[X*R�5�\�m9ı,O���6��bX�'���ͧ"X���/������bX�'{����r%�bX�d>/���5���F[�fӑ,K���wٴ�Kı/����r%�bX�}��fӑ,K����iȖ%�b}��]� �g��.󧣥:S�:_~|�,K���^�6��bX�'���6��bX�'���ͧ"X�%�Dm4�����߬�X�)�u��d9�mƝv����ȕ4�}���rݝ��������
�.�"z��ذ��(�/n:�F
�D�^|��춽a����{v�+0Lq�$nh�%����[�4:N�Z����
�Tk9��:��q�����h���@�.|�8���k��ƚW����]�Z�U��5�ŽW`������ΒHt�N��F̆up0-��WL��$�m�n;7�6�m�� ۭ��b�Z�v0���4f�	ue�k��Kı?{W�ٴ�Kı>ϻ��r%�bX����6��bX�%�����"X�%�ߎ�~��K���	f���=!�w�<oK�,K���wٴ�Kı/��m9ı,O���iȟ�TȖ'��C[6���v�7Ξ���N���~���ND�,K����ӑ,K���N�6��bX�'�k��ND�,K������)��w�=)ҝ)������r%�bX�����iȖ%�b}�wٴ�K��RdN���ͧ"X�%�>v�����HЦA��OGJt�Jt��O{6��bX�'��}�ND�,K��}�ND�,K����ӑ,K�u����Ԓ7lV+,L�����#r\<�ZSD쫸��,07��rQ`��d3Z��m9ı,O���m9ı,O���m9ı,K������bX�'��{ٴ�Kı?d>/���.��ӣ%֮ӑ,K��;�fӐاTzc���b^���ӑ,K���O{6��bX�'��}v��bX�'��߂�32�Ξ���N��}���ӑ,K���O{6��c�2&D�{�ٴ�Kı;���m9ı)����-��k�.���OGJt�'��{ٴ�Kı>ϻ��r%�bX�g��m9ı,K��{[ND�,�N�~O���4��XV�����N�%����ӑ,K��>�iȖ%�b_�{��r%�bX�����iȖ 􇥞�n��Pe�n��+��\�o2�\�gc`6�u��r���I�۫���7gK���CRf�����Kı>ϻ��r%�bX�������bX�'�=��O�2%�bw����r%�bX�=?�����a-�N5��r%�bX�������bX�'�=��r%�bX�}���9ı,O���6��bX�'�v�=��e�������k����ı,O����9ǼcM�֭� �H�10�yz�GH�D�v'b~�s�6��bX�%�}�m����N����O�~"ƶVlL���,K����ӑ,K��>�iȖ%�b^��kiȖ%��L��w?~��������#��9\.��֮ӑ,K��;�fӑ,KĽ���ӑ,K���O{6��bX�'��qoK�HzC���k<�0+�_.ap�2쎳�wL�5e��p�nkvNG�V+^�1��Mn�C3+����N��D����ӑ,K���O{6��bX�'�{�6ʬ�"X�'s��ͧ"Yҝ)�������)������ı,O����i�ș�����6��bX�'s��ͧ"X�%�~���ӇJt�Jt��}�o؆�)���y�"X�%���{�ӑ,K��;�fӑ,Ŀ}�kiȖ%�b~����N��N�G�'����͹g�Ȗ%���{�ٴ�Kı/{��m9ı,O����iȖ%�� ?|? �z��6��bX�'��}� KC����oK�HzC���絴�Kı?wS�ͧ"X�%���{�ӑ,K����iȖ%�b{'��P���r���/^��Ha�b�x��G2��i��:�x�.�]q~o=��擀m���ı,O�����r%�bX���p�r%�bX����m9ı,K߾�|���N��N����������,�fӑ,K�����ӑ,K���wٴ�Kı/~����Kı?}��fӑ,K������K�f����֍�"X�%��>�iȖ%�b_�����Kı?}��fӑ,K�����ӑ,K����Oh�fY�BkFf��ND�,K����ӑ,K������ND�,K��ND�,�VdN��ͧ"X�%��j���SD�j�5��"X�%���O{6��bX�'�w�6��bX�'��}�ND�,K����ӑ,KĨp5����rju��\�7
�(�z{A���G����U��� f��gcB�S�Z9c&�4u�kPۭ*X�f
Tf�=� l!��M����W؎���L��1�]r�p�Nx��3x��:�A�A,�h�NK��i*\���:�.6Jq�I�����j�����=.h��;��gs����k����}/)tO�^�t��.՗��z��	��!�����:K$�$=���=�Nq����J�]����0�SQ.,԰���!Υ��"�j1���8�XV����ı,O��ND�,K����r%�bX�������"X�'����ͳ�ҝ)ҝ?����8���Y�r%�bX�w��ӑ,KĿ�����Kı?wS�ͧ"X�%������t�Jt�O�I��ɋ�F3E_8�Kı/��m9ı,O����iȖ%�b}�}�iȖ%�b}�}ͳ�ҝ)ҝ=���oܮ��A��OQ,K������ND�,K���6��bX�'�{��r%�bX��}�m8t�Jt�O�����ut�lJ��:r%�bX�w���Kı>�}ͧ"X�%�w��ӑ,K���O{6��bX�$C����]R��	�][�˅�����jv���fiUa2�k���*�3 jan�J�i�����t���秀�	9���đ	��q=ı>����Kı?wG�ѕ�5�LѬ�m9ı,K���[NC���A � �@��
=D��>P
��O�,N���siȖ%�bw�{�ӑ,K����ӑ��N���}������T�Ԫ��Ж%�b~�ND�,K����"X�%��u�]�"X�%�}�kiȖ%�b}���C�Vf�uf��ND�,K����"X�%��u�]�"X�%�}�kiȖ%��3"}����?+нн>|��g��c%�ՙ֍�"X�%�~�}��"X�%�~ｭ�"X�%�����m9ı,O��p�r%�bX�}��j��.h��L���,��g�Z���c��N,0&��Fa�	�aB��3SiZB��Kc�W�OgJt�Jt�����ӑ,K���z�6��bX�'��p�r%�bX���ٴ�Kı>�]��*�@Jܶ�K�HzC��ٯ_fӑ,K��}�ND�,K���6��bX�%�}�m9ı,O�C���� ݵ�ek����N��N���iȖ%�bw;�fӑ,h���(�O����]��2H��~�`�� �R��H�!��8
q	"#��$CX-T����bQ�A�B��>*� ���+���B0�"�@�"���ċ�Cb!T7��v���� �Dڏ� �j0�&�	��
M��l��?O����' 7T@��(�RD�#��A4���~��p��W�W)D���$A�1�GB0 ��(P?$>G�y��Bt��x�j~��'L���a$���� ��(p>�U�J���w�L|!��tS�eh	�A�"'f?�@���UD����>=�_o��r%�bX��M�q�HzC��m�~~�V�V��ND�,� X����iȖ%�b_����m9ı,O����iȖ%����"~6��bX�'���_��l��fWy��ҝ)ҝ/￿>'"X�%�����m9ı,Ow���Kı>��ٴ�Kı;��\zB6��6�I+��Z����9įg�G�쯚�ǭ	sl6��V��V�D5�r%�bX����fӑ,K��}�ND�,K��}����dKĿ����ӑ,K��OrHa5afh�VkY��Kı>���iȖ%�b}��iȖ%�b^���ӑ,K���O{6��bX�'zk���fL�4�њ֍�"X�%��w�ͧ"X�%�}�{[ND�,K�u=��r%�bX���iȖ%�b|vMw���f�nj��&���r%�bX������Kı?wS�ͧ"X�%����6��bXȎ� �Ea,Q��'�P"�T���k����t�Jt�O��R~�4����OG%�bw>�����bX�'��p�r%�bX�g{��r%�bX�������N��N�7}���V��&�r�d-)�g��.��jwFt�"únw3I�3=ų��ڛ����K�HzC�����ޗ"X�%��w�ͧ"X�%�}�{[ND�,K������Kı=�����BV�����q�HzC����ގC�U�DȖ%�������bX�'����[ND�,K���m9ı,O����ˉ�6�]�OGJt�Jq~����"X�%������r%�bX���iȖ%�b}��iȖ%�gO_�]�Duh�+G/�=)ҟ���v�kiȖ%�b{���6��bX�'���6��bX�%������bS�:|�>��~	�ғ0MU󧣥8�,N����Kı>��ٴ�Kı/�����Kı;�_{[ND�,KbC�﷫s2�VkY�֤�^Jq���3��a�@r���c2�J�L+z�䝛��]��c�J�/�2L��lɱ�430��CS����n�f��I��U��%�8�j������z� �c��vEn��p2] 6����2��A�8�U����EDx�ɸ�rf���/����;=\ry��J�<E�J��m2�ҭP��];W��I�-֜�h<
��]��]f��Vk���-�8�Cv:z9�*�ZU�lp�������7�#6���L<�̬���ҝ(�'����iȖ%�b_��kiȖ%�bw>�����bX�'{�p�r%�N���}>�?M�*��Ƃ�Ξ���bX��{��r%�bX�ϯ���"X�%����6��bX�'���6���"��zC��L���9l�\-����"X�'����[ND�,K���m9��HdL�����iȖ%�b_�kj�����7�1�Б��[v��bX�'��p�r%�bX�g{��r%�bX������Kı;�_{^t�t�Jt�O؟,?�u�h�)��Kı>��ٴ�Kı/��kiȖ%�bw>�����bX�'��qoK�HzC����x�Q�FY��'8w$v"�,��Q�Fg)�5�D�Ź�p*c)�klRkuB9�]�OGJt�Jt�ｭ�"X�%������r%�bX���iȖ%�b}��iȖ%�c=�Mv�����n_:z:S�:S�����Ӑ�~��<�����?D�5��ӑ,K��{�ͧ"X�%�}�{[ND�,Krx�[l3D�˭kiȖ%�b{���"X�%��w�ͧ"X�%�}�{[ND�,K������Kı>�Ŕ�f�I�3ZѴ�Kı/�ﵴ�Kı;���iȖ%�bw>�����bX�'}�p�r%�bX����L˗��d�kZͧ"X�%�����ND�,K������Kı;�{�ӑ,K��;�fӑ,K��{��[���h����u����;-��(2���Zgڵ��Q&5ݦ��f�(�s�t�t�X�'����[ND�,K���m9ı,O���m9ı,N���r%:S�:{�����K��WΞ��%�b{���"X�%��w�ͧ"X�%�����ND�,K������P�=,�tM�a+TՖ��q�,K��}�ND�,K��{6��c(B�4"�`+�'�'��b����9������Kı?����"X�%�ߴO[L�2�h�Y�3Z�ND�,K��{6��bX�'��ﵴ�Kı=�{�ӑ,K���wٴ�Kı?{^2�x�5��Yun�Y��Kı>ϻ��ӑ,K��?���ߍ��%�b}�{��9ı,K����r%�bX����ff�#_U���s׶q��v(e�h0u��q�B�+�I������,�Ũ��L��,K���{�ӑ,K���w�iȖ%�b^���ӑ,K��>�{[N)ҝ)������K3�Y�OQ,K���w�iȖ%�b^���ӑ,K��>�{[ND�,K���N=!�HzF,o=\��:UTQ���Ȗ%�b^���ӑ,K��>�{[ND�,K���ND�,K�u�]��t�Jt�O���v���n_:zı,O���kiȖ%�b~���iȖ%�b~����r%�`|�'"!���9�ﵴ�Kı;����I[���VR۽.=!�Hz_{���Kı?}���9ı,K����r%�bX�g׾�ӑ,K���OT���nA��1׮��JlWgbݙpY��! M;X��m1�ܛfy��G�Kı>��v��bX�%�{�m9ı,O���kiȖ%�b~���iȖ%�b~���6��k5fkWiȖ%�b^���ӑ,K��>�����bX�'���m9ı,O�k��ND�@G*dK�k�˙�jkWE֡n�����"X�%��������bX�'���m9ı,O�k��ND�,K������bX�'�;Orfj��f�.���"X�%���ND�,K���ӑ,Kľ�}��"X�%��}{�m9ı,N�k���R�5�˩�֍�"X�%���w�iȖ%�b_w��ӑ,K��>�����bX�'���m9ı,M���d���ߪ�����Z�&�GF����
v�.3���N#�$٠�T�)�[��Esb���_S�ܸ��,v�6���]��J�J�W<m��C��ŝS��r�á���rm�����2�e"[*I`��[��a�D�e����Q(�ew9��N6��7cqYTp�2�<���e6��۷t�1�x-��ʰ=��ƛlK��U����t�󻘊@R?e��V�2���-�,t�ic�Z44.� �4��}��֭zJ�3�Þ����M]jL2]j�?�X�%�~￵��Kı>ϯ}��"X�%���ND�,K���ӑ,K����z�5�7/�=)ҝ)���~�|���bX�'���m9ı,O�k��ND�,K������bX�'���=��\����Y�f���Kı=���iȖ%�b~���Kı/��kiȖ%�b}�w=��"X�%�����-�.��SL֍�"X�%����ӑ,Kľ�}��"X�%��}�����bX�'���m9ı,O�/�U��]�ZoK�HzC����]�r%�bX�g��kiȖ%�b{�{�ӑ,K���w�iȖ%�b�{�z��;Ti�b��p^�d0��^jb�RZgL�jF:��x��ݸ��j�݈���'�%�bw;���ӑ,K�����"X�%���ߦ��T'�ı/�����"X�%���z�nj��f�.���"X�%���NB�?�_C!("Q�;�� '�݀�y�K���M�"X�%�}�kiȖ%�b}�^�^t�t�Jt�O�#��f�L�2�iȖ%�b~����r%�bX��ﵴ�Kı>ϯ}��"X�%���ND�,K�w~$��d�]d�%֮ӑ,Kľ�}��"X�%��}{�m9ı,O}�p�r%�bX���xޗ��=.�������Z�.���bX�'��ﵴ�Kı=���iȖ%�b~�]��r%�bX��ﵴ�Kı/�OR��el30�Ma�e,�tݍ��,bx5x"]ò۪6��&�D	smΤm\�ɂ9����ҝ)ҝ?|}��Kı?}���9ı,K����r%�bX�g׾�ӑ,K��tY	�%pQVJoK�HzC���k��ND�,K������bX�'��ﵴ�Kı=����Kı>�Q���u-�ޗ��=+����r%�bX�g׾�ӑ,pP����DH _ �v~��'?k��ND�,K��]���N��������i��kU�"X�%��}�����bX�'�׽v��bX�'�뾻ND�,K�����=!�Hz^�x�� ��j]T�m�r%�bX��^��r%�bX���}v��bX�%�{�m9ı,O���kiȖ%�b ����3,���ԥ�Yj.H�4nr��R���H�ZT��yt�b.�,�̸�3	��٭�&�}t�t�Jt�>��v��bX�%�{�m9ı,O��絴�Kı=����K��cy�'!$Td��i�.=!�E�}��[ND�,K����m9ı,O}�z�9ı,O��}v��bYҝ>v����"�/dn_:z:S�:X�g��kiȖ%�b{�{�iȖ%�b~���Kı/��kiȖ%�N��O�R~�����1Wy��ҝ)������]�"X�%��u��v��bX�%�{�m9İ(zB�>�j%7�~ͧ"X�%��>�p�bl��%�󧣥:S�:{���v��bX�'��siȖ%�b|g��m9ı,O}�z�9ı,O�=�߯穜��u��w)��]&�W*6i�bY����0�#�Mׄ�넎�W���x��X�%���siȖ%�b|g��m9ı,O}�z�9ı,O�k�7�Ǥ=!�K쾌g�Pl��J��ӑ,K��ϻ��r�G"dK�����ND�,K�����9ı,Ow��ӑ,K�����̶��G3N��k6��bX�'�׽v��bX�'��]�"X�%�����r%�bX��}�ND�,K�!�I�0�XjL�˭]�"X�02'�����r%�bX����6��bX�'�}�fӑ,K�����ӑ,K����ߤə���4a��WiȖ%�b{��6��bX��5�fĐI����M�$����A$O�TU�� ����TU�� ��QE_�D�TU�� ����(���A�B@C�����
���**�TU����AQW�QE_�D�TU�`AQW��E_�D"
�������)����Ā����8,����������04�>�>� g���mi۝��s{�( (��QBAOz X�S6>�WhC�� Z�\�p݂��iJ��CJ`-ЈQ�g^���R�ȅ�B��ՇM�Ή d8V؂[4R�@�-6�ܮP(��u�agBT��╭m�WZ֔�f���BQ@���5��`r(���ͳkl�eڤ*�Bu�J�*Uy H
F�%J� 4     ��*D%R@444  @ Sm�H�@    �Ѫ��)�       $��	�#Bb<����R��))F��44bi&���t�(�;Q ��$		�B7C준����?����X��UPTM�  ơ.Q AU&kҙ�;o �ɷ�W��o�K�V�0�d�6Υ�},�����JHĦ�B��w��od8	�(��HA��BK6Uc	��>`�J��	!#CX��;G�u�,�f�ƶd�_6J�/[7�fe�+Y� BR@�@�,�x�́%�ՙ���!%�K8�t,Ř�a�/��I|gY;��!�bY�tz���r�d����5:XZ`B����dܾj5)���&m�j��AX����	�"���@�G.�w;tģ�=#-$`@"!��(�0�{p;{��Xq!I!a)-�*KLx��5`�1� ��(�B�xJaA�,`��XDB�!D)��J�am�PJf�:�BR@�����`H٪9/4h�a*�!t�Y�8�^%$��t.���,��]�Y�wCb%��<|
y��u*&MH��,e�_n�
XC@,����A+XeZ�wa	
�E���_�XJcD�(��Ä)�B��4��S-��DHFzF�Q%�	a(!	 ����	fL,�ė(�FH2"$dqy�4�9sd�yx�t'!�c
$c HT��ݲ��G:U7�Ĳ��HH��1����Axj����wd@*H�DjIL�PFj���i�j�Ғ��[����x����d)�]��1z�!x���2oG����  h&��)ԑ��J���:qЉ:tH0�л�k�Y�[8�C�!	,:��o����Ų3y4�g�J�/R��.%�]Ļ�Д�q.�q��,�1�BB6y'ߓ�1f	C(�L("@�r�NaA����Y������(B�KI`wc�*2�A$J� K	#�l�����\H�q�HbK��d�z��5y2����%h�Vd�i*B�*�H �A( �
	Li�
%�
k��=��U*'\��V�d�H=�y�֑���ˡf8�#"r��1�Ec4[�,IwQ��'�4�>���z�~'�qa/b�JK4�I$I��1!e!R�R�,��N1,ޡ���e��L��6��غBX>u-�d���e�q!3	���B\8�1�4PNM��!e`�!A)#BY�X�8T��V�|Q���*��8D�P.):��",`j�UB��͎��u��(��#��JYe�o���a8.̤w�o^�& 	�g�b�.�T,c���Al)��,H`n	Eq�u ��<�4l�2"瀵"�*�h��<_E�I��U�E���V&!��-g��5�
j��bн��^�l�M��)��ud-W���r�gCp�d��)���$Ѣ�����*�[QzCQ�HK�v�^��x73������س��t��}��=�{oFp
)��gU}��+-O�-kr8R��âS*G��Q��@�,�1�$���    
�������)����l�5���Ub��@-v�.�ڹ�&���bC�ki`�@!��ڻa�ٔ2@@͇��p(f���@!@L�AUTҺ�Qh�e(.�*�UUBZYs�*�2�Ȁ*�B�b�� Cg7i�SaJ�%�;;iuʱR�VD!�P&�lg&-� l؀�A�V�P5Vb���[u��5v��6�H.�[�Z������l3�\�B�!���
�J���i��6��E��(�iKKM�jh6�h�@�֋�9�du�e��@m�U��[��u;j�9a�miqя0�1XQԔ��4�6ypn3�6L85��m�@�C40^Q��k�������X�UC!�kU[UA�m2���ͳ��nZ5�R`UPԆ[ UP ��l��e]����������*��B���a���Ɩ�*��-�eUv�@UX���ղ�:႐������C��V��ݵ∮[��7Nꔙ�bL9ڑV��5���m�܋H:��j��c2�!u �g`�ª� �2����֍�*�lPvR��m���f���l�����m�m� ڣU��U[lV�b�+�m��UUx��#�ʻgc,��*������ ��m� �ڪ������k6�QE��C 5�Z̪� 1h`�UX���*��j3a���cS<��M���T3�U\f5�B׀.�[c�.��i�[p�(���f������P 5���L51����ٶ뚲�kmA�:��݀0;&.�m���]��UUU��6P,T]UUPvu�cK,�[�*���P/�f�,E2G�mP��i46���PR&��l������	�he��K�g��.^�J�C���fPh�!)�,�׺]�u��:�c[n\1L���3�nuPdkM�m� !WKm�q�Z�k,m�*�
 ��Q;U��6�sk���mC;"�j��UUUU��	�KF������������eUUUvJ�mUUUU]�j�+��1��zz��l,��"��,�����+�TA[
�UU6D-�l�eل�\����u���:ڴ��-2
Wlk*�0�m�6��8⃳�mÅ�*�ȭ�K�U �UUP���6�h�� -����k����l��-G
�@�HP��t�f�����]Iu4�[��Z$6�+�W��Ǩ�GU���6��
Etr*ml�ڃ�uM���[��sF�p���q5�@�b�Ȫڶ�� ��li����ڨ�ܠAUx���UUUUU]�ڀ 
�������;]�Vၜ��F���UH-��R���]V��3L��X����UUUU ��Z����Y�� ��P7M�� 6/"LQ��&�3	~ڙ�����{:�lA鈸� H�!�a@k����:"zD�J-|�7����G�`���]�z�_�@������Pl#��� �A��pI��Vz�����g ��6B�{,IB@�����	��MVE��K��oǁ�NЈ��G��S��<i ��!(p!�Wj<t�`�x	���p$:8^::3�m6����\)6�6��lx�,^�'�4��Xr`@�c�!}KW���B���3pa��0�h�_�p�fҘ�ghT2ED��**��4\�f���HW��~�7�|��%E��9��+��ͱ�M�A��9H��9(��6rJe5�f P	��Z��FRU�T�0f�2�6j�T��6�ML�
�3�UT.Ur��HE�QLnŚYvus6A�j�:[`�E[a�dL(*M���%I��qC7Z���ƈ(;��.��:�UM@s뛨s���n2,4r���V�#�k�DE@k��Ř�W
�[���ԉP�5�5�������\�4̹`�]�V+C�]��q��#�$hW5Wg�mmM����Amx(�~�;���8w�^�])8&��%j�BV]e�-�Ы�k�\)�-hhKJ�r�&�jh�mqE�m�X�*��L1�j@��U�I쓳��w�Y�m&�&և�I������׼��f4�z���yBut�<r���v���O�K���D]+����F�h���n}�w A����]w�%�V?Z�����k�9��~ �f�B����*�e��L+�z��>�Ǿ����ۢ@��@�fO*�{Y�����߿~�ڻe�0V��02��wQ�A*�7�'9Z�*�7˽�)`��������)""o$���6�]|-�@6i�8�Q�"� |��M�w�K���{uy�A�A�}���H<�9�A�A�A�kګ� �R!���b��'9�� � �A�A֩y�>rM���ڋ�):�]t"�q�-��ip0ZUu�j43��[�]5a��Zl��-�*�::f����e6qeq��\j�du�;�t���w��gG�������b�5�A����sWh<� ��q[3��� |�CޤDD�u�%�yh<�:�<� �t�ﵳ�&a�xe���]�Yp�/2�4�؃�R{A�,D�A���� �����\H� �jt8![�D�lb��������R���H?f�*��Q���sg��� � �R{�'<����/�vh;l\�F\�̹�h<� ��q{3�ٚA�iq�{��ʿ^Z"���!�� =�A��Y�ܻ� � �T������fR9H9�A����Nw�vߣ�t�LU.T��I��ZA�iQ�{�f�*��~H!����9H9��s3H=�7������2��y�A�R"��}���"8ssٚA�iq�{�NV�$əu��%Y�+�e^^R"�9H;� �=�]�{u�A�iq�^�fR9H9�A�A�A���V�{�A�A�T7�A�V�YWh<�:�<� �t���	��I4��|=*`2UH�:�\�[���b+��Ka�[�j)�3&���������j�ڗX`.{9�Z�}t��Iľ]��5��V�6Fa^�N|�7������e�]�󔃚�D�]��Ofi���~`>�<� ��}yyH=�9y�A���}���>wo�_�Me� ��r�^d�x��͵�d����+;o�}��r�f]͎���9��'�Nd��y?O��k�p@3�
�`�~|�ϲy廏M��n����z��=CJI�d.d��/�e�/��W�� �Z2 A�b0�	"$!#$","��,��t���q��G?{�'ȏq������(ً񧅔����:
�K';�o�/�7��N��-�Q�� N�A$ߚrs���ͽ��2]�%�6��J*���"�{B*�t"�l���j�ت�!T�R*���� ?����^�U�hZ�U�Uw{3�~h֨��p;�g�Q̵{�9��~r�A�k�ϟ7'�����OMl�9�:�f^B�v�y�'Mn�ͷ�6�n��@��u�f��v�o�m�M曒��w?��6 Y���.�V3(�B�\�.+��3D�T!�P̦.-Y`9F[Vm��eE���˳a��|�Ɖ-]J"C��ˉﾪ`�����ueUMDw��fx]���e�ک��O��n�+(vE���/�3����j�%�wd��;w ��ٰ�h��Ovc%߾�������`\X�Ȫ�����v��w2O�[��f�t��f2���f�pN��6��{f�u���\M�ݐ���I݂��j>��\�̓���v�~y������spAMtX�l+�GtM�`\N�� ]�0H����k n�jǧ�t6�XIt>�s}�/����� ���ri�Ô�bTJj!��&[�}�]�_�6�X����=��o��|AGv� �ﱿD��7`���;��� A0���3L9Rs2�9`�B������h�MLm��R���qPB;0�]+-���2��+�]Ug���M�>K���i��2͊�Y�ޯ���~�e����^��d�� �-��2荪�{�{Ͼ�^mU�7�v '��(��	��`��Q�r�ʀ��)6�Ç-��H� v�����dE��ӧ��5w�����w�ڇ{��݆;��7rHn��G{!�͠'v��ʵ%-�K.ba�R� ��Uw2���"���%��:���෭F�����T��7�pI��d .�����$�<���~�n�n�������{[v��ݽ�������ݻ���e�y�A i�	g2;����ge�D?��iXL����n�����9�����Oh{�tIwﱽ��|{�{EMO�u_X˰�_7�YU�~A�Y@"*��%1�$!!Q����t�H����e@/)�
�%B��L(���ċ)�5'�6\�I�Q��	��#�#�I0#"���@!4Jd!	 %��dHBD�!B,!!MZ��'��0!_��<A����vU ������p�Z�3���E+
	0-�Qquv��F浻8�lJdjT9�:�L�eTv�X���lA�2���\#�0��]��4��
[l� Ȫ���{�� 
�mpl��6{zW�q���T�bb��[V6��c
U �c�]��W2��2��tʶ�8�]s%�� +�vHf�9�]�)��F�6�`�f����Ձ��`��� ��0��nPlj�bV&���U�Ճj���6�ؗMM���mh�3ʆ���)Eج�A�qrj� ��\j�b� '�O��''8N|��6�F�k��U�kVB�������� �;���V�&I(d�!�Z��1�mh�p��M��!��R�
�XRhV�h���e%�|<�8�v�$���{��܌�(WR�ŘS.]��UN��^~Q'����}N^e= m��ͥ�*�7�cf]�,Q��&\ÈQ2ډr�&\Ko"s<n}��s���7j�D��y��wk�m����d����w�/�t�V˳EL7���?>[߁q�|�(��Mm� ��}���} 2 @�I ��S����9�ud��s��w������ˌ1�+������ߕP�z|�z�n�߽�/[ݮ�~r�-�� �d���Tv<���E��r�R%�2�Q1��r�*�����̨�Ns%�U	���VUC���v�@	 @��>�ov��V�y��nǋ�hD"�Z�#շj�e�.M�Z�h	\@�L�������ƕ-���j�aT��g0��QTW���#�>��د)Fcѷ}9X��VeT����9���:��	Hٲ�k��h)���<����߉��d�Z�y��ڪ�z�^7�[s���׽�����|�s�Bh0
��*�Ǖ]7؜�x�ݻ��[y,F�����q�
�>����:��eeV�W�kMFm��
��}�z}��>�[�W=N^e?��x,�Qcv�� �DP :��{������+2�-t/�ˆ�dKr"bb"�s.�؝�7>��s����"�>^ov�#H�ȼQ u��E}��y�Un܀���@�;1-���/�w�m!�k�	��X�EL�K��6 R:8��j�H�՘��@
Į#t�@)ԢK���٦��=�?ߺ�i���,�Q��u�g�sS��̪������h����s�����g���J��6�i�-��M���$]�Z�y�������!R0H 1b%�PlB �
&�������r���0 I��l����w�=�Y��wI$��ݸ���P�"d&҇:@3R�9����~�7�9���g�.�}�a�P'��G�8�6廬PUBA[lHЅ6k����T�D$�,�R�M��%)� �P��tN�����O/7d���å��ov���	��&6��~rU�Ag�;�ϟ?�<O����X�[��A�����Afچw`R�n�����b��!��[�G��:�UI݁��@ H�t}�2��D��R�[������*�6��@�q��A�(����ڠWt��72��\����c��n��{#��>"3�>�2�"�#�Ș㪢M��!�j0�h� [5��e%ul�m�0*LFdi�0�''9�&g|��e�D��na̸�86t�����w~φ��^���wA݌$*�N7'P��Lw@�g�M�zTC��f
�6���� \C2�z�(��2(T�ى$R�^ϗ�Y���99$�{�9���y�f�#�H'HxEL��֨�}��n����%r8��,�P�a ��b<�wd�f������{~��;;P#1��z=S�,ϟ4H�_h����UQ����^M�;�)> 
�^B�֨���yCv,��N9l���@�|�yL\堡Ȗ�ĵe�r�n�����C�.�g�#�]��gj�������M�'�2����43`�r5C�����8e��ʕ�-Gs�t���fAw�=��r�!�oA̋Y_NL�u
�;�-�+�Ѐ��́��A^R�s |n��>ѹ�
i)��i��5)��hK��gZ�֘Bl�r�#��h"sT
`[�&��X]�lfZ�I]�{t�^w��gP�maV��c�������w��rqx���^	{�c��]@�m���p<@!n��u�$� ��r�#�m�7p���m��J9B\D���j��e��UA�������fh��Sh<(������ �mC;�)B��=�fhxtC�1�sӲ��:����D�A˕!��v���q����Ǻ}���<��Vdx+GP̊]dG��F� �$��#���_�s-��!wv#��|��=�#��#=3�8M�2"��e�s�6�(gv#�]��g�L�_}�F��A���ܹ8��[�1�G���.�j�A4�+P������~�����oݿ�i�,9tYi ��+t5Cv����[8������� ���7C�dF���Q�@�q2K�S3CQ�7`��g��8z,"t*&��B�b�KJ��aO!$�je���cYW	v��rJK�k �˵�0�k.!6�5bj��&v��@TV�-�����ʒ��Z�(U��.�9Թ�c����A�v-j0�ˮ.�q(*P���"�ر�l9�&\$3ՐA1��t8λ$m6��X�
8skDpj�]2 <Tu&\
#Sc�q�`#r��Z�������Q�Ll
!���U��a.Hd&��m5��e��	lH�Z����Q���J0l���6.U,:l;M\P&����Ô��U�D[mm u�Q*��b�a�1���6��4e�u�]T�<"}?x�/�#��pSo<�i�_�Ы�\+��H��L�m&��\l�k4З\ƈ�
�䕮�q��;��攳k`%��W��S^ގ@%qv��hK�'�ng�	���4;������U�'.�
GP��7b=��H�6��	d˛���Áh�uJ�S���0���ۡ����<�ݿ�h�G�$ dj>Bv,X�_s�349C��p>�l��́h���sCv�>^yg�従^��e���"�.d
G4�̂�v7CW��t������A�@���k��wA����AfTC9�4�C25�&9�)BQ�e!�>^ygϛ�y�|�|Vq��@�gpt��݃U ����e����a�cۘ��h[u�>>�g������i�׾���4�D�12��gu2���[t7c�!{��<�ݨ�s R��~߇L�F�݁Ă� 5���:��Rw`b4~�/|����Q-�����䥋�.�LE��b�6x�4xfXkJ�ݦ�) �(��ĩ4U��O��s����ٷL�k�0S�����O����r�l��r����q��q @��|�#k�y��TL��m�݁��1�n���>�{g�gδ���)�gز�uc�Ѩ��s������h�H�m��1(N�ˏ�K���<�p{�Z3�����=�s y\��_KgvdC3s����u��̡(VՉI�{>Shn�!�/ӓ-�_Upw`b>�>��n����Q��:��]���
G��/��S3C��7`��a\G��D��Z��K��T�.�������.hn�����a��l�@�q�3v#�����D��@�ӳ-�C�rwt���~~�y���I��v3�*�n�����>K2�́H�q�?o�L�F��2��[ru��@�9�G�f�t����@<<7�LM�LL���]���`[-�L�B5!���&3�5�����B�7E\�"�IF�^3L	>��iӷL&�ɱ�%f����t
G���7b=���m�7p.�ne��:����c���k j�Kv�݁H�pf���[q�r�ә����f��hn���*�-�8�$2H�l0T��1|:�hn�uQ�*Þ�l�@�q^Iy�;���m�7p'���mt��<�������s3ĉ�?/d��k j6�<�mĳ��p����B�|�8�FB�`��Yi����d��/��/_Iz"B頯��
������������҆����t�X�HE����34=�q�9�%_�m������<��~��<�
b2�7K�X��hn�uV �!x*z%����.��؍��j6���]72��Áı�D_��{O�S�^h���v��7� ���mĺb? ӽIgv��]���Xۡ���n���g��B���<���W�е�S�^c�Ѩ��=TCƔ��I�N�_ �D�6���6�X!c��Q�!3V�S`H(�TˊsF�,m�`ae�Y[.]v-�W;����\M�il�M�Q�W����>|ߥ���_�2[:�T��ϗ�]�5���G�ݧ2��G���b��t5���h�~�_d4���a���Ɏ!Ng�1�ɚ�R@�SQ�.ßD�s RB�3 �`���j6���]1r��*��@�g�Ljj�$Dʑ0�s.T�r�f�����=q�᳙#�fA���45��Ǳ��9��MÁh���sCv������ژ-��a0�]�r���;y��A2��n��hn����錖Π��F痮]�5�57��ݹ���=�-B��>�ȉ��R�D���nd�2��#hoA��.-y̜B�������݂�GP�z%����4�Iy�;����n�a2�+�=���M�Zɋ.�P�B�W-��B�Kl�W-ٙ6��
��I6��nn�M���[V�{��ƻ1Fe&�(��L�r��*��@�nuz��݃YQ�{#)�g2��]����4<M��m�;�%����)�́h��Du���9�L̂4(�'gϛ��/<��D�e��A@��u	�3�2y��!�����l�Ps Z7:���݃YQ�?I99����ܢ����n,6w`Z:��xf�D��Z�n�AN�=Yt�� :H�"����Q�|�\\��A$o����q
��y�s Z�y���?k��i\�\RnΩHt5Cv�}1r���8���V5��K���#hW�eL6s Z8�gL�=V�rE��������1�$�I�Kp�!Ng�j>��4;�����a���s Z8���ͺ�Cv��V���*��@�VJ������Xx�,ă��J�gk���`q�20#B:-Y�4���	$T�Il!�$���j�BI		!	!SƷ�G��H
F���� �^�3�D��p�	��Fl��627d\�����+��Z�`	�ɠ��\l�bLM 1��]6b�����aEU��+(��� �*���2m��6H�*�&M4��庨mn�#�u4�n�ܔ���WX;[�(QX�b�([E.�-�ɦcd�j�im�řW"C�ℤ\Zi@X\�[�F��ն� �nq�1s�#�UV���u��nq0!F�Vk��T�W
j6Z7
ֳb��
����.Hd�f�E.�-m�V���l�@-��Q6��\�S16��'$�B�ô0ݥ�#����^�N�F �L�t1ٷ�ErUWK)�]efJ�Qpq(�5�,"0��\�r�K�[��%��vv4l���(b�9�4����wy�ף�(�`�ð�T��k r��1��r��G���b��t5�������Z���բ�f��P5C� {fl2)؊钳D����O/>Y����6�j��hwA݁��n\B�́H���ˡ�FЭ��-���^t�����gch)�j�z1�#U�/��!H�@�u�뙡��U�	i�45���>�<���ǨZ1T;ͺ�C��Hw���-	p"I��E2;���{����{=�������t\�w`R:�#�i��r�4-(�{�=�ߦ]=���v�w����E��̬t��ˁ��a�D�̀��){����n����j�S�C�h�@� �~^�{>^>i��l�<��UUs֑�`l�P�j]C=�3Vk�`M0�8`ZJX,vR��JU���eV!��$��W�;J��bmJ�HfQy�杧P�{�FZt1X
C����9��R;�);�����!��L��s�;y��s��ۿ��v��\� �"[nƢ��d�.�;�K�R&� �t�{�9^�y��������l�@�q
G�Z�SChb5P&� �Sd4����]�����&��;y���c�f�#.#Hm�='2A#A�� 1�����r5�=�̡��1���8�!����щ]s�V1&
C:�R�*�g���{y�;�:�����)/-EE���@��̏�-�A9Ղ�f�#.#�?O��u�n�W0��ps�`4q
F*�O7C�1�[3���)��N��t1p1+Cr[l����v����}kB#�R���@[jP,��ۃL��Tp�h\�l�7���\4�+KeV�f�2Y\�:{�P�_�����M����$�>�p=Q��0u
G2-!��왡�ˁ��aϢdi -���h�P���b4����~��f9eR\;mq���!��j:��n�G'�z!��F��^rܶw`R��|��1�#U�Z�2q
G2#��=��ta�9�Fy>^�/;g�#+�'2#�R1T#y�����
K�ء1\�Y#N�S��i>f���ɄJ$�R@�\?������x���B��v��	��:�<)C`�u�/{��ry
G2#S��]E�F��k�ë(�m"��t���ih�{��!Hj7q���Q��0u
Gv#�c�f�#. ���c%T��t��v��~�����2���J��t1C��Oz�8��#�׉(c��CQwQ�+�z�����)k-ME���@� {ڔ8�
aC�!.�h�)�����.�L �0�Q���lHcs%h �]aU�ʭ�V%H�*�9��[���3pmv&��)����\�T@:�����铙��)���F��j�Sއ.!���ϟ4������i��˒b����Cw��@��g�}���� �C�{Z��C����s�j��G�Ǯf�#.#Hz�B~��JA6"��W���z��N�|��Fn�W�����!������˃�45Q�bb�.~_\����![�[9�<I�:��Sk���(b"�D$���$HP�SChb5P<��`�� �Gv���3C��:Õ���#�#�a ��zY���t5�5�<����i��t��Q?���?����\�<�#�����ˡ��V@�m��l�@�>�#��WZ��C�w�W'�]��[�Q��4N���:#�ػ�
���a�P��m��f�q��݁��Yvs #a��]�@���ֱe3j�r^��Bb��@��k>O��������O�9� �Bы��t1C��O���8�#�����dˡ��@�i�(�����fQy�v���O/?Oط��5�@�hj5�<�r��)�`Z>�깡��B���+铻��) 7�У&b"�ܹ�fS��N��o#Hr�)
~S��8�#���Ho=�.�Gc�U�"��4�G�_�eKgv#�|GĜ���oj��Q>^y�~��?�d4���vs�3�s R>v=s41|B�j6�%{EJ�d���u
F�?����iC����@#Fd�y1�l��d
F'�����P�P�)V��g����v���{��@�q
G��QChb5P9��9��R9�)v:�hb2�b4�87B'���6�m%��H��lm`�)���+�B�BAD��@��#P������X�",8����.���3�w�6K���k��e�@�\Un��A�٨dCl	@%v�&���l�!��6�c���6I���4Ҫ1]��t�,Ɏ5�K�����:�i�r��
���8���VPѵ�q@e��`��ݝ�Z] !Q��@n,r �S5��\�����b�m��( I]�R��U5M�	c3�r�63Z�ڡ�2�-����Q�lʄ�%@,���\4%��B��7U06���P%��0jݮ�q�U�S��� �\�؊LVlm�Z�[��F� 2��˖e`"V�re�e�\��T`���F��%� +�����z��ߊ���r�.�35ba�6���	���,j���eM�l�ն.�S4JCMuf�Ttr��_wv���4�|��l-mn�5�S�>��!H�7���mF�?�Lz[:�#�����e��j�b4��wr�{���'f�o����f��&e�˼����r:��߫.�H(@E�#ʹ��{�9gNn�G#yF#Hu�+�Nd
G�j�����iF��������BR&��"��j<��n;Ͼ��h��
�{���� Or��fS�ѸpĀ>@8��z���]��ȴ1�q}`��d
F9Z��;i[]Fܠ½����v���t�́H��P|���!��@��~���	�n=��`g�h2<���{>^w�{y�>�o�.̠L��a�r�9�-B��ֲ����B��w�1y̜B�ջћ�n��.'P�̹���Q����>A3��j�"�Z,�aCnL,���ͻ ��4Wa@v��-m�dH�nf��J8V��6A� ����9�b�0Vh�۱���T
}�r������{&]F��HWC�K����=p|=�q�/=��t9{�~ �a�,���s'�s R3Czۡ��x�$	�%C���9�)j��~^n��Hb5P)��˃�uA݁h��Y
�6�PɈ%nr*����{�����3��Ѹ���nsr�r9>W-(����(�E�8�nd�fT1���;}Ca>��H!02�H������Nw����}v۝�z^<�㺦_�*���GI���a�瞦��]�\ͲSX�D���f����\�+1����o(OtNd窨?/7��N{�tJ���2ӄ�q�Գ"��m�]M�&W+�6̮�)1�����m��5&V�h�8kr�tΉːr-�߿W}��|n��}�/�t������s���Ј�N�� Ćt�j�*��{�q��`�{��GkwV�<��yY��}�>/����ћ,�6�"�ļ��Å](���z��h&H 3� �CG 		�6n��6A^i.���ʹ$�;��A�y�@�mN�d��P���EPF1�
�H?G�"���>SM63�(D�8/4>�Æ�7��#�D6�G>oa��_Xz'vq��zT*����\F*��?Ns�;�}�?;�ǽS.۶�^edx �	�D�00A�	uFͶ�r���!��LL�'*aÙi�Vc�5�w�5��'��8�=�8���f:�<��!�G!��Fku��@c[A������+�0ڦ���)5�)����;TV=[�/�r{$�9�w��g���k(Θ	�L9ne�z��%�V?��yj2l�^�g���c�9���o��}QL��]��fۜĩﯪ�}��w��&��A��4���{�r�o;�%�V?Nn�ߦ���J��ق������~�_��Vc�7���`τ��AP;��|�}�bF���o��r�ږ\K��K�Ģ>��W}��|_{��Cy���R�Ssr >'I$�'�ݐ���{w޻k]h�T\¾cǔ'WNc��j��yX۝�z_�#kv������?f��m�П�.Iu�u�(�.��@,X��j��lp�f�k�7#�3e6آ��\�P�27L����$��;��"G2���U\�~����WJnm����r�1�M�ͼ�<�s���?~w���k�v.
��B(�cnw��y�����` �{���r�]���D���í]L\�{4�P�0�D	��`���T����|���<}�>ߧ��Y �P�"mz^�m�z=/c��?��(��������>�ϯ藙x�u����o���ψ{�4 hV�7�6�G��ܩ C����!2��<r���w�eUN�=/cs�T˹v�k藙x�d��) �_��I$��$�@�����'	;��$L=+�u[�?�,u UD��������H��H�(Q	0aE�#
,b�3��%˾�C�7) ���j����8g��W�s*�~�����Ʈ�G���Q���oSFr���� ��5��?tuI����~�U��e;����8R���94߫��e��~<)|���oNS�2]*�G�w�K�����������X��K�O�=�W�Z񈖋HKQ!$T�$*T�%)$**B��Q�(�(+DV� �m����B˾w�2?v��=  �܌�[{��5M��Rg���fd�q��_�|�u�;�Y�`9*{f���8yG�˲_+��~QhY�8r��.�~Y'χ	�\��RI$���t�����^~���<��ʧk�9���}�Jp��ګZN�����FjI��=m�_[��L�7{c ��AY��yp�`��[�|%KL&1o/�I$�]�D�n�I$~�'��������	��n�$�n���o��OPx=q���i$�@�I�;�������F<s{��4�#C���;9��R�����yi����i~=:I$�拌:+>��{w��~*���	��dڨPģ����萶�9�A��/-s��Ʌ�鍤��*_:��/|�?�.�p� pʾ�