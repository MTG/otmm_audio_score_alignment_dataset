BZh91AY&SY���K�y_�pp���� ����a|_  �
� �  
U  P  @

 P�      Q@ 
 �xP��P��* �*@
�UD$TJ 
 R��)��P��!U%B��I@J��R�(
UJ�     h (@   �� �������7�}uw���Pw�����v:7�o���>��	8��ǳ�Щ	���{ڴ'��0C���73GZӉ��i�У���kVǼ tw�S���T绽QMy�v[s�MP��z  � �Z� ���J����r�M��znX�� *�U��-\�t���n��z Q�I,�8k�n�z ��F���c�8 t�ꜷ�G��{i��mk��'����;���0�����®�U�       � �z��c��{i��᜜�� )�U=�91�W�Η��g�y����d�;�� t �<Aݽ�r�=�OzQ���s����e�q��Lq;���s��fN��y+�EP��      �� t�>f�a�ZI��:, =.t.[�!ݏy�+6�� ��!��i9�@U��2���X�����e�̜�+��a�>� w ��1e���9�L�� � ��  �   nn��>�'ݒ�z{����}��R���)b�r�c�n��Α����e\�p@"��T��L�� W�ޡ�o����{�9��Op �p=��y�{����.*�       i�6ҩT�P�a1 щ��0�%0�5%J�      �=UJ�20���4214d�4=��(d�4�     "���E6�R�@�  ��  �A�T�2�M5=CS� 4�CM8���_��Z�g�������u��k��DU~_�
"��TTUO�AU� ���/�����y`������?�DU^�ÚU�3��������6���'�?ͯfF����9�"���֒I�GS�Q�����C:h�V��7!� ���n���y�/ā����2M�̢�o�Л�j�$ˊ����#x]9�CLwף(�,ͯ�p�*)DSۻ��}�F�ĳ>Ƽ�&ԤCG^���B��;��=ζy�L�~����&���X��J,� ���\�E�����^�¯��X����/8�(��2b��B5�� ~!�DF}$�י��^��̈���9�o{���I�[�SN�Z�X�^a�5鲬_4�Kwf�Fp��f��&�}�lW����x�L�F ^�%3bȎ��U�$k�	�:�>��֮�O��3F�i�4����E�D$��s�|"�� _|�ú}܋ ڠ�D���<Y�gEt�ܤGRF��%{���+�o�yj}{��NǼ��ō�D�����W����0���y�,f�yK�theC�iP��������O5���ܖh5�5C��L^����
�|�t�XL���p��).){�2o3��Y˳�����/z��.Ovu^	{o~{;���|-J-DX������jf�.�	Z�$��B|l�_VB�dd�	�O���$c@�M<��Ϸ�_2b	;�y�k�Æ�V�%W��h�a��+��$4cJ��D��8�}�vsB\�*�H��t�ǃ#<�f;g�D]*�r��kA{��\��D�A:�,d@�����C3��Kw;���1�P�!���0O���I��&�f�V����-����.���h���t�@S�s7P���|^;w��R�K��59��i0m��V`��%	a�7�xw��<::7:w��;ӫQڙ.���}�9{=�F���rrc�~���KI��{k����|G���K�K�X�QD����e爷�/�z�Z6n)N!�]߱��^��f��5-Ꜭ#�5MWԖ7�?�rl�K�N�S�w��r��y�Z�v��߷s�X����s!yb<����"�(,h�cɌ�=�A�1�[�1�2��\�6������ϛ$�	s#xCnG�A����m��C�s��SY�/k�Yu��7����Ni����4���%MK���Ȣ4Aϗ6�C��VCP��P#mFഗAB�o2eͫ8�ֆ]���MՅ9�NB��v���Ið��{�u���-�+UY��m�Υ>��Ċ����Z�M5My2��CP�p*
��G;�G�?]���w.hȃ���0HŘ"��}7��w7#~��H5�Pvjp֚�$��L`�� ��ց�p|�u���w
�  i�N�ˉܬ�v8�I����cb�2���8�(�'1Eq2�	�k&3���h����7|�^����N���j^SV�2��K5�պ�U��c;���d�i��¬N�������<m\�cꦂw��v2�܅�,��Y'0D�XɈ��>�q�����r�K���v�>N�Z9�g%[���^���z;/F�:���K����~�ٻ����>ש�u$����,���x<�<��ɉ�C@�.C�>kbF/�8f���d��_t%�ݻ�=��}��}�㷗I���B"	R47���9n㎚��W��pC��q9E3���^�-��y�:�w��qgn���>��|�3)og(|�Sʈ��C���&TV;�q��� 4ch�j��D$tTU<�:0�oxpOuj�/�ED>9�h�˘���s*,sDLDL�ē�:���sXADH<�4�I��B�XVTO�8dC�M�l2)�kD	`�8��SX�	}��g�!�C*`�N��Q'm]\��9�X��gS�q$��\����j3��4y�������Q*|�㹻���kٞG�k��5HDI!ޜFʶ��w�T�3�X��o�Y��n�5�gT�Tǎ \�l�y%��#w�tI��݁%F�z�Z�2�q������������X�Yy�_�ތ�ZD(|n�E�8�'��:Ƹ9'2���
	�
�D�eX��S%k�p���\ӁAZ��r����C�歯�j<�ۭ��%�����4>O����Ө��ȶ'[�^�NsݼǥN�8�NQ������3�O����|�J�aE�7�=TXܷ��غ���8sI�O�N&"�G���ӈz��k�8$U�N���u2��:�:�!M�z�ub���38q����	�� ��8)w�˧5B�Q�}�,�G>	�(��F=}�E3y�1}�c�컧7�>�
�@Dw�b����>@�p!�=��+JT��D4�<��<;��&w"lI|H���j*����ۿ:7ߦ�+E�PA FSLHX��Lp2a�VuY��Ν�w�druk�ߜ�����\�E��:&��o���v�ι�����)�����sЩ��`�-���;��×�{t�d��G�D�N���Cڧܤ_{����U�}㷛�f�&6�X�_Oo��v�la�Q��/�����k��/�1b�IB��Hs�E)q7�@���E�%�+߄��z�:s�ߩ����5<�y���=q�^�A3@���M��Z|qc�
���\��PT9���&Lx��!�Jy�H�Сx++9�άfL�;�&�J��1���M��~&��_m�%�}��{u
�^wy~�>H��]���%،��T��Z�&���Q�V�'Y	�>8�(&��C�ϐ̻y>]ϜB㢰�.-��n�~1��ݜ�����|47i��������A]�j�c"�7��x�wf��[�V���n��.�76��Β�S�7�s�����C�|��J���8wRs�I-,�{����N��u���K3���)iZ`1=�����?	g>*�e�L�"3��;y��]9��ط��.�A�4��CI�A3!D�c�G����o}=a��ٞo�}��GWa�s�b[M[{���D)����1*�o'54�ugWF�Hn$�'&荚��M	d�N8|�K�C��!�'E��ix��3�o�+�q��
dC�l���'yx�=���j�>Ak�74�T�RrZ>ʳI�8��m[��CLh`�ŋ�y�4����u���I��8#�|���t����L�v���{�oxd�w�̺ϪΊ%ԙ�,�Xf�=0��Ա�ѳQM:p��鍼��0DMf.�yt�qf5��,�=0�<�a���~C�;��*a�8;>>w^h�%�fy2C	�?+ZIX��1{]��s�)��78��(2�p#'l{!�c�}�TFE������h�ǔG�sp�W�uq�����t��+NӛÈ�Zz7����o{N5����X�w*���p#Y�İQ]����X�(�ӈ�6�f'%�������r>
�q�Q�o<'��.�t��e~d��VΘ%��s岱)H��>��|{}Ǔx
��c���ܔ�l��z|�4�����w*��e|_,��?�ANi�~���_^��UV'�/�yUg�\E�:�V�L��cF�Z'��pHRclC`;P�J�T�k%HY2��Y��[�R9Y��q�dQL�G�,�	�☤ǃ�* "!�<��ŉCw�{�n��Ld�־��Q�w{�-5Z(�^�Щ�f����A��=]YGR�GM��.�I9�T,�-�P�v��1�a�LL�	(��1L޵�20̈�D�is3���h�:t$	�`h0%� 0�(Ųn�p��h�&�%aE;ӌ�]����F滘���z��2g�_=�D�p2�	�1�'Gԫ�o|��j�$s������xc��ɋ5Z\>+	p�f��������͹tHL�T(nT̙ŀ��ʡ�A%�0LE/����@CC2E�:�-���[w�;7qk�N N�ϖ�̝�D���MLX�"�M��D��aa��F�ki�R:���w�yϴw�~Y�l�q�'��C��x{�\�CPO��;���Nr+.�4-��ē�t���|����W��L.��#.�c�;ȞL����H�i�-%����T�9^����_Q�ND�6�/�xn.N�����[����{:滯^�v�מES�3���߭ع��C��ٞY'�������o8���R�Dw���ٗ��w�S�8ܡ)WT�N�d�k�pQLS��(�;�[��s��7�Y�Vq�\N��9à��qc@3�wA=,")��ȇ�1>�8���{��5�|ĕ����C�.��No�{� �=;�|F�$čL�h�0B%�߅���">��K��c�'*���s��'p�0H�#� �a�fq�&!�F�P�Zjb��'�!�3��t\�#�\�[�;������<f�G�K1�����%�����C@�3���8�R�G�t=���YLK4�"(|'r�D�ED	�� �xp�tx��>����bi�X4B�ST��C���/3�
SC��İ��Јє�|�eRi�/���hh�<j�'�⒧��5�PZ^ZX�״`���������YA!�b"�k���$,sP���#�!«]Q��D�SDsdM2�څ���C�'�X��_/�$W4������b�"&)\�5:Ҝz�|�"�}��]�ϸ�ge}�zeF	`7��u<�'*G%�8���i(�.)w>仉�q������F	%���;�RިX/xUӢ{�5����&��t�����S���Īǵ�c|���ݧ#�\����Ï>�'�1����ϑ�x��[�{��Ga�%_�Z�T߾���x�R�^k:>o�(�/K����9w��Q�BIwEa΢x��cy��f���k4_kA�1�tmc#(#! R�j�V	��x�XsR�,�=Z�fv\�yw���h��yE_y�ӟۿw�H��!��$��v�9Ѡ%�p֠0�4Z���Oq
�WV�99���οNg��+S|5�y��{�Μ������{��QN-9����S���Ӽ��[���;��u{d�v������}i�/��9�5��v�C��ȕ��Ō�N�-T�N��p�<yT�>��Qj2Tq�"q��c�!��&2�<�2b� k�ǥ������i`�k4�P��;�p��2���m�������X�߼��;�o8�7V8P����fu�2*�����ɛ��*~���vxY
60*���xJ#./�D���B9�)�'��>{���u=�Z�Y�h����v�>o�s���в�U��\�g��u��yz���W�Q�j'7����~9�N!wu��q���k����LR������0Hk#L�;�"�Ym��^�3Z!(J���x.�H�R���ۉ�s�'z�*zE�w��Y���ҏ;͊��c��syR����]���oo_ŝ�4D�c^l�Bu���J��y���(����g=�I�$�/�%�9.Fy�����S��b���}���;;Óy�'5�zH�N)��F�����K�s�L��V
$>�k�s�aψ-ŷT�iiw���O����!�F�"�)L�h\�~A�P��b����¬�1�
���ܪe>�A@Q���+���7�_{ھ�}��𜺈��D\��	���]���;��=�>@�P���a!t�ӈ��3��$c���5;���u�>ސn"N����jщ�w��so��D��O�Ḙ���N�m�h�,[�1Я��
���Y�깧�ɑ9<->h(�ܜĭ_|�B��4���(߫-i�^<Q�T�g�;�<���ӛ��{�@�P�8 ΀�  5�@���m���m�` 
P` [E)�h�l   6��   ր   ��      �T  ;e��b\˶����*L����Z�� WT�9���]RkFyZ� ��h���U���g)@Pڴ���ķ�tꛥ� 5��s۰�lԫd��cW��bh0���-�u�ۣ�ڕ��1{e����Y$dyj���(�8�0��T�CvG,6؃v��;l^۰�yl�UUJˤK�.G�ב����H�q"�m��3�ƥyM�Q�Av�m��#y�e5�U��<�m!ɤ|˓&�]�@S4죗kq���j@���v�V�s���6N��=�5��i�rB�Y���鐘5�\ܔ�P<>֊I���3�ƐX*�R��Ò�E��ڴ�ɀh��m۶==�tÉ�mW<��HԱ�0�z����Z��f�`���N��V9��/���l!�۵��C��b�K�Vm�:Ci��fT���S�Sa�'m��`ؤ�6.�]0��e�+�W�zU��H��]���tT�L�(�&-�J��E�L\@4��T譮��lS��"���Z�n��=E�V\��3U/-mU���ݶ
8�v;�G��mmÄ�ඬ�:�2h�S��Fkq!�@J�K{���,���K�H�vjX��g�n 8�ν5ܯ6���KC�ʗ&��,�f 8�m���[��5c��9�9�ƍ��#[����m�����J���V([��iS.�^x8�86��_ 5JL����Ç�X+�ܩ���A���!c3��,��U������ҍT�5�M�����*����*r��n����)Cm�:su�lUj����]���΢�V�mrM�.,%����tۮKFC8[A:R��ݶli�P0C�A�\�>N�����鵴����[�E\��En���V1j1�`)Nu�*1�ڤ	]c���9B���v}Rtر���ʆǾY��I���i�t��f��i�i�\#�.s��'L���G��K��,�ܻZ⤧7V���-���X�)���/+��2��UJ�R�Æ�ۖӶےK�]"GD���"ܑz�^�$g���k�m��f��`�pm������n�����Wi����}���)�%|���j������||Q�pҭ]@u�L`wZ�VU�_*�tUE�H��66��K#v�VԄ�nC�y+j�N�#2*Cm�-����p�I�m� rBp�^�mi��%mUL�۪v�@�6�
�����S�<с��Q�vի\��G������ݮ�a����:�k���eq�5Ok���~{9�dW�pݪA��Q����D���+��OhAܕ�plq�s�r��������z��#ْ��Eֶ�s�.��b;J��=��5��n��$N�Sk�t�s�,��	D�{���P�(e92i���dI��	�Y�S��)�B:�t��v���A��q	��^� ���Q�,�6��٪�U��ԇ�Z�r��<�5#��j�~GΒsᶥɇ��'a��)+��3��lآ,&��{[��&-��e-@r�UU@t���P�m�f�uD�� W���3#�j��^�q��\��줗-UTQUʻ�[�B�mSX�fm�i� p6�,�ݱͣu��4�k���z�[v�` -���Y�]�8�m���t�� �>w�}u����]VC(� 6� r�nV�
��K^T�G�A�Ӷ�TQ��Z� $�kOB�[J�����n�a�H��E-�m�B��
4�8�T��D�g���\T���������z=�\T6.�'[;R�u̮-�n5t���Q�J���l]@��c`.�D�ur�v�9N����]՞.�t��<�t�o:.�;p�k�a��O5�!u��ݞM�e�k�Q���8�Lc$��%[����y��:1�Hf�:�^��Βl���4�#�'j	�k��tr���I�+��:�6�P/�ɛ��7H��*��%ʛV�p����B��.&�zی��O�h������|�һ������l3�D]�tt��������v꜌g�Ƽ����6�lM�;�:6��{]�n<mX{m�i�cy����j��!NT�\��bj^\nӛGi���A{��UV�6�`��q���u��5�>��
x��j�K�d̮��U�xaSr�7��5T��d��q���lv���̮��w{nЛj�Ek�Zn��8%�V� �����Z���.
����[@u�]R�Uk�[@ÉwkD�`�6��j���vJ#�{�qK����n4�X������*�7۴�m�[P�hj�]����;=c=f�i�ST�!�61T�8����ݐ���8�ۅW[]n�*� ���l�Yæ����ݍNϚ�v���n��^���[�~��6q��X��m��+�@�����WV�q�ۮ��m��,{M��k[��u�j��TP⪫n� ��@oUJv�am�W�P[U!9`A	:��6��`�;m��pN�Hm���f���VԮ͵]-���u�ll�I�K�(�t��nH����Kh��^�������lr��Nʨ#����ً���KT��UT<ˌ2�UUJ�P<�(n�tUJ'i쵸�PV�!M�7jW��,rA��a4�J�t��5t�U��(ڷ1gi�'Aִ��ͷU]��i�l68�ORԃc�#���l��@ !6�3Hn*rX�m9�2nW�ݝ�d��V�T�H���<�gbT�	�IxǺ�ؑllIZ�V�B�J�,�ZJ��y�zGv�,$sr6�Z�n׫�fl�E�S�j����fi.�ܫ�iv�T�W1�vhp�Z��p\�.��'�7^�!Ŵ�8I{[%K�<L�U�a5+��O�l]\�C&�m��V��D����9�l�m�K.�M�mdH��V-�.�[�+`�n���p*���=D�գ��zw+e��k��G+� �۲�m�e�7n=�R@%��jNu����@+�W:�N���P-��[�f68ݷl�i_g��UU�Nˢܭ�2��f�ۃ��$6���.]�T� ��ܒɑ^l�����f�2��gm�����u�U�j����x�w(՜Uu7n���P�8xl��l$$�Y�(�n�[�ݻX�t���	m6u�>|>$�� l��]+U�k��I2�� ҭTUQ�A`Giu�jZ�V��&N �H�
��ҭu�k��j�hr�~�~> v����R�+e�
��p��rG-��z5���iG�0���ɮ�gc������$vN3WU��:5[�g�*��*����
�UDs�l p�8��Y�.S&�V*��UHc����8�۞YY#Z�n�[Pp]Kp[�T��m&��e�ce�ں�{n�j�ZU�.an�sI���l$��iV���*�j32x�:�����XĄF,�f�kmm5�Z�{b*��؃�M��U@OW��[��鵲�rN�t�ʹ� �@a�pqtcl��Xێj�UH᫫ջd�� 5�0���@ BU��VW�uCn�Tly�����j�����kׯ<�%]�+r��<]9;�yxUq��@<��sR�v�}O�.�����y��V�*�v��m�)(.�1��x<u�F�Y	ܽv�\�]�8h%��U�������N³������@� �h�v�GbKY��`�K�[!�YG�n�8%�˱U�er�Cq���C��\�[���\��Ė@#S���UHM���S�����@@@`K��U�D,J����UUWJJ6.;K'E^�^r�=���We������M������j��B��sy`iV��vG��6��;>��d��Ӷ�ms$p�L�t%"So:�Ӌ-����9��"�9�����0� GHT�Yִ^��pm��z���'yDĀ��j��.��eX`���v��{ H��l2a�䭭�4��?n/�l�U����!�d��=
�ڂ�I3���T+.�.�7i�gDjv_����Vqv:��=��(|���i8jT�2-pi��;k m[O+�܏��9 ��b�����ݢ�/�6��.0��']+l�%�`�[ؘ
Rek��wH<�+��8V�	�Ԫ�g��V2*���JpA�U�U[vݪ8 -�Լ�Q�ѪU�e�hk]��hd;D��U, m]��
Wf���!�vۤ쵷l���m'@�nض��Q�e��V����Ԩ�E �m���6��t��tĊP �b^y����m#=,�ܦ���n�Zͤ�$d8PiM��l�¿��k�
��*����KWm	�m�RAes�f�$���j��PM�j�;e̵W)�������L�yv����8ŕ���ںU�U]#lGY�[m�`r+��U��`  �ru�Z�-�kj��6��ª��RYB e���mPp�5�]u�j	:M�v�FFV�ٚ��Pݶغ�#v�OXщ�tVyrm�[gcF�,�uU����l�֭�m�C�[S�l�UV[D��#(�i͛3p8�pC7Z��@ZńMJ���n��Q��n�Ip2�+� �*�U)@u�bAz��k�dHz�@VR��UV��$��m%�Bn�--�%�mP'�f�*��K��Wj�P�y�����۫���Wt�[Amz��� ����06��	�q�yg��Q�J��̰�j{J�j���Ӳ�@�T��5pmn����5@�K��� ��M�l�UI���}�㴫�ّQ��OuWPJ�کٶ{lKj5݆��AΦ�j���B٩`��\�q`ۆ���N�2�f��<�u���U_�o�Ъ"������:�������'��!���Ђ?/j���� 	�JB@u�B��P@4(�{�!�� t=�H!�g�**x��!��T�WåC�Ǿ�N�6�=� m �>$�Cᝀ&��� ɈfH�`�'��(@@$ hC}+� ä%%S�TqSf��$ �ȑ�� ����BAءڏc�,��>;���W��@H$=SBd�>_U`=pN��@�'J�]=��EH����x�>#�<S�T8A�8*��hA��VIPSj�$|���E]+�B���=@��S�P�C��Wb���="���J a�;	Cх�3�|AЏ�x��(�(���4 Q�
���6�=�M"��`	ҏ�@�+����@OA_OTE�h$!a��FX�Z0G R ������/���U(�$
�H�"z��O_��ΑXBN�"�d�bZj�
P
U��(&�R�`$$H�"R%)��bPh����)V"
eү`��$G��Y @~P<Uu#B!PI�(�)�L�P�"�b@��P0E����F@%�C��ġ�1�JP�j���0�<F�{W�O�$B �>�aIQDTHC0Z>u���P�X#�~Pp �D>N�J"� ��X��О� `8�� �$�t���ȈH�՟�"��k����=�ϯ�G��@�"�X	Y��Hh$$І�&������s4�
b�(RB�t1-�H� �a`����{�W������}�<�\��l����M��h�S�M�݃�{5�4um�3�G>:�z碍�V�@�]�VOc<m]�K��]�\�'�������[m��C,����X��4�QcvvΦ��ܻzˌLV�jva�jv��4��n�}��l�Y�:�l C6�tk���'`�s�7]�h<�&ݰ��n��rvj��j�ѕYkƘ���Ԙ�lnN.�=e��˹;u�.A�^�nQP,t�0Z�f�Τ�s��9%�pٱ[oEͪ��z�;i�'	�,6�m\�+NG�f%3���cpWy�z�Z����T�/F�4X8�9��m�y1L�]�� ҇ 6�T�mX�jݴY�K6�g�SN�m�)5�1�r�A�e�<������Y��62�s��쬱�kՕ��bS�+Ƨ�DX�Y�8��v�ɤ�J��.���b$��s�%'NNwNq��]��6m�D�8�r�=k��
Gv�{\���u� �l�I��<��=*��x��@� ���$�֫%�����c��Ob4a�c�1١���n�ԝ-�����$hrx�z����1����e;v�ⷬj
��spb�V���!�8ݻ	�ϵ�<�bۤ�vhG;Q�����A�z�˱�[�r\�p�i����s�����l�����l2��2�*����7 ��礘�+�;Y����h'�@�H�i��6#Nʹ����"0�v:�q��l�UVq;&��94�C��	Ђ�zX�;g��g���kѹr�S��j��@p<���7&ڽ;r���N�=�n3�ZhI�Y�:�o�ï=�GbĽ�LlcPp�$N:�a�����H��v�k�f�\qcp
�{)�[sj{�n��Ҝ�9�4!��v�]�p�\㵙�P\鷎��R��-�m9(mN�K���X^зt�h7�x�[�F�h�\�1ݙ@ɰ��#��w[�Lu(Qa�����k;�l��;ˁ���U���;V�XU�'���Z�ΰil�q$>;�w��}�{��=� z����_"mU\�#��4|)#�!�+��0ǘ0�K�7]��l�1�q����Ɨ�u�"���{c��'���,�N�!�ĸ�n.W8N�������ջ�vn7l�;��؎��`�Ͷ���ɟ��q���U�6U��zMm��p�N�t*�k�۳�ػn�Iv�a���`�0nR���n���7𣖎^ʢX8:�9���2��P��̝���C1�����D�q�RI�["jen���pf�8�E"�Pk""dII��s�s��aw'�\��A�$��S#�8娫��y�Iw�H���_�U�'G ��ݷE:m؝����}��+ ���o�ܰ��rn�_��m��}��+ ���o�ܰ��x˒�R�V��RT�V۬����_r�{��}���9{�lI��j��V�~���s�>�ݕ�}���<�^9��Wwi�tzVs���r����8��r�k�khݝ��0�ؓ�v��]���,���{��}���>�|`��,|��%m&�ب�庒�~���C��2`�Y�e��W�D�p�>��X�w< ��+�gR�cwv�n����~��s�7�vV {���se۫�(M� ߯�d�ԐwH�{�V�^�!�wA��;-��V�ڴ��{����+�g�������(M�32����҆�N6�=��zA	�K7m'+��y$j�JY%Hm
�cY(��[m�K�{����s� ߯ܰ��x�J�K�7e�B��m��>�|`���w<~�ed����"��BcB�1�l�>��n��~����&I�ȬB̰��P�����,	��e`w>0��w4�n�t�ڵwl�{����+ ���o�|`�]��bj۱Ҧ��~�e`w>0K���jI}��u$���zS(� ���l팓�F��Z����/�����]>9�"�����hV�n��M��s� ߼��{����+ >�P�������(M� ߽�Y+�U~H;�x�镀}���=�j��-�n�jڶ�`���}����$�|ݳ�|�����Ut�	7cm��{���������ř�"^��.�6|?Z�h��61�X�όz�� =��}߽���W}�A�**��72(��1���R!�vm���������͒��ѫXu�@&M�ـo_r�{��}ωZ���X��v�n�lv��v� �������>��X�{���Wu���;��t��o ߹�}�ܰ����� ;�x]�Wh.�
Ս��M��P�|���>. }���;�^}�%���W'-z��~���粒`�>0z��_���*��Vڤ�:�\ۭzY:9��vqM�gL��u�l �����|���ƌ�V�E�:2����D��㰤:��� �v�6�ںY�͍����ؼt�s1��Μm8�-L�5T��1�q�w	<�ήM�ЋqۛnVuA;8Y�m�6n9�R7v�R)9� [�������������$q�%^Su�ފX�M�v��Ku��3�L*~^���_c۾�ϱG.p�,���='������"�U��lHn��R��&����V���[�j�u�#��X�ό�_r�>��+ �YG�um��BM���X�s�?�~H�\� ����>��������?JQ@E��U�/���}ݕ�}��X�s� ���s����U�3VpD$��o��y�9�}����oX�s��ݻ��V���� ��8{/��xp
G�x��+Q����J�RjYVZ����Ulv4W^\lz�NK�BN;=���v��{���3�xp����B�����
�+��Wi����f޾咫�7�o>�&dA��&4e*�Ab����",v�p�p��Í%(=�,��wV�[�E%m�ގ{��s� �_r�=�SJ��c��Wv�	U�����=��}�ܰ����7������m�i�l�>���ό��X�ό﯋ꫪ��H�z������+mjIzq�^d鶄L/UU�ӳ���Q��v�A�J�X�Qd�R]���y�{��o���9r䯄��~��Jـ}�����ό�όz�/���ݫhbj�ـ{����/��"!TW�/�����W^~Nն�&�ـo���>��X�y�{���
��ζڻiU��0�>0��� �s� ߹���D��y�I1G$Ǖ�eU��A�s;��b,b�����u\%n+�������nd������r�;���7�|`�|`����+c�6�V����J��/Ix��}��,�u�K�]��`۱�ـyzK�;���>��{���g� �)Tk,+�jK�z�jK�������u�����I�ਐ��|�]֭rI���.�l�>��� ���N��\� ���}�y.n�t���mu�������uT�nUz��)�
�*.��7�>���ZJ���0�}����o�ܰ�>0��r�7�=I�C��ݱ�j��}� ���`}~�{���
��e�-ջ.�Ub���_r�>��� �s� ߯�`�]��j�)�TRV��>��� ����_r�;��`�P$ub����j�ـfe��;�fO ��À}�g �����<_�ʂv�9)$�*�r�SZ�f�ᩐhxҌn��Llkp�-�i�/=�@Q�/Fx�c��&��z��j�qv���Ƈln3vM��ݽ�ci�S�ܺ�v6�\�cp`N��˗�LS�~����ٺW�;Ȑ�dؗ�.up�&K��6Y2)y2���2f�����㜃���<�i��w�W=n�v �8�ttM�T���!\R��"��IZ�陘�p8�|V���%q%�6Qю<�;���0fݸ��:��O���[��Wm&:ln�0}r,���_�`���>��*��Lh��Վـws� ��� �s� ߯�`���I���.�l�>�ό�ό�y�w��wY��;M���V[Wv��όﯹ~�w�+����_%�_6��J��w��y��i���=���;�޻v��6�M�9y�s���&ط��n�.�R����fN�+o<�ٗ%�'/G9k��{3��-,�36�����-�}�`����յ�n[�{���f`�@1	Н*c�A��~l��ߴ�������^��QR�k�U�����^��=��>淪o�!z���c��n�]��{����}<�����z��IJ�4깹���������K338�>̨q��]����F�!�<N��s��ݢr�����;\lI�|]������s`����Z[���Wwwe|}����+|�]}v�`պ��j���fgBPx�u|_}�i�$.��(r����,�d��x�u�fs��8��q�A�3CQ��,����H���C˖�H��1GH��}��퇹�k)h��<=&!(��+ZLz�

:{������Ҙ4&��Ϧ�g��+봖$�`�$���cf8�8%��h!�I��_��l��B��p�z:#��735��a����m�lN����TY���79�mw�
�>=���/��R#����=�������K�38�p�ө �`�'��3�����r��z�鹁�H����0�D$��X�JA0��2��q$5CSIAI:������u-2Z�Ӭ6zQ���g]vE�q�d�e��d���Ě��: ����O��'1�Gp	�V � l��D~+��ׇ���������"��P1��H������b����� ��z��QD�4�����D)���ͩJR}��scܥ)1�QR����T�UWuȄ<��=�R�g9�mJR�����)A�P�!'M�r!BǠ��n�Օ7z#z����r����s[R����6=�R�g�s[R����s��)O9��Bps-��v��!��2�T�{n�n�\{`���{=��D�����]Ӫfã��SmJR������)J{�}�mJR��o��A��!z^�r!B_6"S�JUeBu�m�L���>~�鹂Y�9�9��R��>�5�)JNs�sc���>��d?IH*Ғ�c�n`�aC�s���)Jy�s�ڔ�I�s���A�9���!&��ɕv �Ѯ��o����R�3�s[R���9�l{��=Ͼ涥	!���	�tb�� �"T�!=:C�f	�C����cܥ)�~�͙����E]]]�!BM����B�	lJ�X��Q��Ģ;�ˈQ��]��/��۴�=0�nw�ι�7�Y9�X�#��kv�{\����h1}�V*�{��u��)J{�}�mJR������)Jy�9��JRs�s��)K˜֭2~���+"rٹ�Y�F~��ߴ�,���s{R���>�6=�R���s[����I���J���7wL�ĥ<�9��JRs�s�� �>Ͼ涥)C�}�l{��9�Ù�뮺�5u���u�ԡR������)J}�}�mJR������)J��s{R��缄��7*��u�m�L���<���jR�~%����l|��=�����)I�}�l{��>=8���&������i1*�䌱�E�84�a��x�+p:�&�S��Jc3�����ջb狢G;v���{U^|p�םqPR.��q���F+Yy�u����b�ٺ�ܲqgD�M����ݟd�l0���jd1X��vdI�j޽c��9,���H6�����ȡv����yCq[Z�َ
�Y��ѭ�v��d�	���@N�]U�
3��v+�����Cfa��n�`�:�H��m䊬J�"S&!��V*�eN��"o�[��ۥA��H*2B�9gs�������L�����9�R���>�6=�R�g�s[Q,�,?~����-EmB˳m�3�0�<�:�iJNs��ǹJS���kl �@���tJ!}�)tꬫ���%]M՜��P��A^��GH�	�{��O��d?����r������jR�a�������U��9t�,�,����kjR�<���ǹJSϹ�-�A	�o�:D �G�uU$�쩺�r��uֶ�)CϾ�6=�P�EI����ڔ�'�~���R��>��ڔ�X~]=���H� 񽶩F�l�����'�Í;��;%8�j汆�0�s[s�{O��Q��k�oZ����R���u�jR�����ǹJS��9�����J����g`�a�����e��VWd�s����6=���!�a�\ڍ)��9��JP��y͏r����\��� ��JO9ȳ���uu�NgSuuw|Q�!Bs��Ȅ<�����+��g9�mJR��y�l{���ޞMC���U)
Ie��$$g��6=�R�g�涥)I�y�l{����m�"D ��P�L�Ys%+���[��)J}���ڔ�>�9��R��9�5�)J}�scܥ)�C=��n�ǿkxL1�uk]�����e�!�g�[-k�� M�9�?;��?-��m�1��jR������r�����ͩJP��s�C�JS����ԥ)??��2��UU��Y%+&��>"D,�{<I R��s���)J}��ڔ�'>�9�8�ĳ~��q'?X��'k��%(y�9͏r����9��O[䨨,�JFS�a��#1	��ւӎb6�@Ӂ`�J�NǴi;�{�ǹJS���[R����߄�S�W%�6K��qf	|��5�)JN}�scܥ)��3jR (x�⎑"fK媵u5j�T�\��Zڔ�'>�9��R�<��rڔ�>����)J{���mJR��Ͼ ��orw���wd(Gg�s�h؇�ڸ�t:&�n���^��q[��FmQ�]g]u��R���~��R����s��)O}��͠��'=�9��R���}IJ]�(,%]�Uw<�A�C��t?)*�)����ڔ�'�~��cܥ)��3j�R����kW:3:���4u�[���{�)O}��ͩJRs�s��V���s��)JN}�u�{��=�D�:�utV]W\�@�O|�)Os�s[R�����\��J}�zLJ)����,�8 �`v�� s7���)JN}�k�-%��B'.�Ř%�}�{��)J9�9�!�R��9�5�)H���"D-�����Q7ET����������h즻v@5�O\p��K9�Vv힉N'V�f "Z�iͩ�m+*N׹�Y!kݽt�A����!BO|D;��=�\�mJR��~�Y��:�#4k�fk���)O��9�iJN}�scܥ)�5�fԥ)9�9�!��߽g��#rR2Y]v���N}�scܥ)�5�fԧ�J�I���^�:D �M���!B]��s5e��fu�k�u�[�(S�k�fԥ)9�v�"D,�7<�@�jQ$-{�ŜY�Y��?&���LJ��Id�s�)9�9�!�R���@s�~ͩJR~��߶=�R��_s6�)IäT�����9Ό�F������Qu���io4<H��Ʈe�գa��/g��]-�	l�nk�M�V�X��6䇰O����:�6���i�X;n������}�k�;�2�l�ñ8a�˽��d��D睻7iqaղ᯻��X��6U)kk�<��ܯh�w ���pz��3������� u���"vӍ�74>]���vO^�ٲ]S�������s;n`���bUH���>0?�%||v�`㭮8���q�U�bn�[���<��]q<��u��������\���֎z�_��ܥ)�����R�����6=�R���<���A	�v�"D,�R:wJ�֭f��:ֳ]fԥ)9�9͏r4��>�[R�����\��JSϾ��"!.�9�%՗wv*&��:D ����u�)JN}�u�{�)O>��6�"Bx�⎑"�d����U�Z��3]u�)�H䟹��_��R�����jR�����ǹJR���ԠR3���(��#��cr�8����lڔ�'>�9��R����u�)@��b��"�s"

��YTR�
�� �ۭ�x�nو��Ʉ�p[��lO`Y"��8�Q�-��s����߿i���/>��mJR��}ιܥ)�����	f	a�yߨ�,E���=�R��}ζ��O�(i�P!�'��zM���&�h!1.�ҡ�� z9)I���_Cܥ)���ͩJRs�s��iO=�,�g::�:�tZ�]u�)JN}�:�=�R�}�6mJF�����)J^}�:ڔ�B~�s.�͂���v]�8(��">��ͩJRs�s��)KϾ�[R��O1�t�A�qH��+����	���յ)JN{�scܥ)y���jR����u�{��<�_s6�)I��3��u ��m[�Ŵ�/vS�5�ϛVc/n���gj���؍{d!�Ж���is�:D P�	�{|�A����GH�Jy���ڔ�'>�9��R�����C�(岕��-��,�,?{���ŘR�}�s6�)IϹ�l{��/~��m�,�#=�~�7'��%c�uŘR�}�s6�)IϹ�l{���aQ�	��BJ� v����9�[R�����!���?~�dK��&R�e���0K0����ǹJR���ԥ)9�9�!�R�<�\�mJR������u�ֺ�2j��j�:D �G��!B�<�n�)O���ͩJRs�s��)O��_�]���h{a�f�X�z�nY��\��@��$��	حV6��3,�5��ΰ���Z�]u�)JN}�:�=�R�{�s6�)I�y�m �R�����jV`�������)QY��wQ�Y�Y=M�Z(��!-ǻ�"D#5�[R���s�CܨR�g�\�:�u�Yk]ekZ�k�ڔ�'=����)J^�wȄ�	@�D��ފ:D �O+u�`�`��y�ߥJWmrơ�L�R�K�}ζ�)I�~�\��JS�u�fԡ5�H �. K�\%?('B���~���=�R���$�j���ڹW35wȄ!?c�'�J�	Ϻ��6�)I��~���R�����jR��{�5D���Z�" ����ۑ����x�u��y���k�W[8�K��3%�7&��D��n��g`��{�\��)IϾ�6=�R����lX��A���*:D �M��:��.�뮺κ�jR����9��@@�/y�:ڔ�'�����ܥ)���ͨ�Y�Xw��/O�ZYX۶��g`�a{Ϲ�ԥ)<��}��P)O��6mJR��y�l{��=�g:n��+�u�]k���/�d@�>�����)N}���ԥ);���ǹJ�	Nk��B����ڙV��UU�uַ��{��>��rڔ��D�7w�>"D#5��!B^�V9Q�!R��<>������ f��T�i���F���e&Y��5����Z�LQ�z��E�@��p�Et����A	�1�=�dk�i�A���v�6�Q�^`k]y�����f�h�[�3�M�6�f��ЇPE���â1�aCR���\q���Q}���<.������v�D�z�F�}�J`���LX"v�<�Xၜ��vq7��VU��eefFf8X���p�ZH�z0�&k�T�'OR֎�L�������Op{�rn�����^!��d�2�5� ��+������Q�����J
o�n�Y��CUh�&;�g[�+fCUv�Q��*� òe5�NF:	�{��������(ŵK�b(
ԜAk��$�/������J� 	�"H٬b2�Y���-�ѦcڙLLl��d�a�X,�9�3t�k��
���X1�$�f�u=Ŷ�Q�Y�x�x��7ŀ�T
�T볲�b���esn;2c2�����<��#XWu<�Mػ]��� u&�����wzȋ��1d�/>�m�F&�wP9��&:Nu��[X<���i�gf�ח�r3��wX�*�ݥ����vڂ�9��ڝ�����(1E�v�g�lݱ�HM�h^[lܾB���<���m�F*�!��vF��SQ���d�D�!���li���''1W={n�p�n8вq�1Ŷ�Y-�l����험�!&�;;p]�'"�i�`�v5л-�۲#���ܻvf���ۆn�S��ڕjf���(��9������]�R�hA׆��m���vd��z�'�n���ѭ.v�=�Zi{kB�յz�)�;l坡��r��IvU�i� ��z����IY�kCkL��,E�E��D>K�C�f�lYݠ�C�l5��i1[cY㞟jl����,���ϋ�|l�r\˝c�6�\t���]=m�V�o,�M��0�=�0{n�:1�^N�������D�{v���^�Yn( �G���L���gd��ۢ����%tK.n6]��:厬	Ŷe�n��o,�vڼ��,�`xYm���m�[���Z�;6��*8�e�h10g'j��.��`�v�МIHp
�b�4��8+ ��uܨl�X�N{p;/6NLl�;V=k�w���p��bg<�[d�5,C�|����ӤU^N/$lr;S!��n.3]�q��J(���H15k�Z$.4�t�����k�lϞby�Q�;��O/:��㳭����m�]�7f �����˵&��u'QS4�3�u���zZz��Yx'.�"�dW[v
�n8ŉ3�J�7jU��_�ʷ���Ӎ]��^NN��@P{�p�n�lm�;bvV�<�t��ݣ4���K������_��Hȧ��(�G������!؈�"b�(����h@��@>����0�ɻ=19gv�ٞ�ҋ�g�lX޶�moFq�dy:T4^ٝT"���n�(��m���ڻ+�&�x�un-�[%�uW�
�@��nq���`8�������\���`-��#�ڭs�Bs�ݔ�a�i� ���	����Gbո3!�LBr.��(c�h�kdd��?}���QK��l�z{9�X7;���F:5mD����03�¿������#/gf�mp�_k�qv՞z��ؽq�y�.v�,�����_q��6������D �Au��GH�α�")I�k�`��R�{ιmJR�����Ru�\��D��8���O~z�I���s����)N}���ԥq��" "���st��	�Y�)JO~�_s�JS�u�fԧ�	!�y�߿l{��>��~ͩJP���U�v+��%�/���BQ���jR����scܥ)�5�3jR4�̬r��B��uC.�-Q7wsuVmJR����l{��9���R��{2�ʎ�"{-��A�f�;�+n���ݓh�89�I�]=�z��&��G�'v^&:�U�|��m���Ӡ4���{��A�u�y�7�t�[5(K�Hk���c�)�As6�]\��\�}�o�~��1�L�42�8�A 3D)b����r�\���@��9��㝝�	V�����h�,{��?P}/��'��h�"\e����.�յ����&�u�x�|gCbb�ݞ��U�˶�n��˷���XUS�8h�`�M�=:`R����-]Ю����wl�팘�u�<]�/KA[����v��ny_����^Z��Ʈ��[X�L��޸�?c}Ԓ�DB_�Og��Ҫ���ʙ��p��nx�@<���<����ΉB���ɻ��E���M�����:�<>Y򈪈P���!)o��:��<���UwArww7wކ����	f����y�@�Ss��
���{�r*R��ڕm�ݵ�w��UUU{�|`�tK��qi\aeU��%e:�)XS�a�=���n�Z��uӭi��VH18�H�q��S� ����*tc�N�a�w�E�N�n��X� <o���H��v����Gwj��'I7J�����,t��}W�����l�n���ot�� �3�D@g���6�������خj�b�xP��{�Ӡ<w��\���}���	,
~q#"���Wm����HUE*ظ��S3w�=�����B׻��m?�N�!�t�ʫ(WV�՗t��4 UW+m��DL��Ѣ�J����y,-��rJY�L0�m�)Vbm�ucm���`���}/��7�DB�@g���;�[��] �]�\��zα�4�
!Hk���8��z(J >�dʥ.�s%�]ܶ�t�������$��}=�(�*��;���~�U��t�t��XUD�2u����՗SwV]U]Y�c}���!(������Ӡg���.�A0��("0Xs��1�l�W-U�MJ�R����t�Q	x������A���G��s�1ձ�D>miv�����r�����4SW	��%7Z�] 7^�я{6��b��VZ�vQ��\�.���;kb�ks���u�t�Om��9�A��ηZ�4�h�NB�k&�#Վ�n�R��@���=<�{1�h;t��`-t�ćK^��nO]���1X{3.n'����'��{���na�⛈DcP�D����eCM�[].s�����iRB��(\��"�?fciT��i:vӰUe�π�����=�!�w�����@�*SW`M��Tլ{�C@�t��'�M�>��g����aj��?:bwI+y���镀Ot}�:�<��hD�ʫ��6ۻ�`~�{���}=�!�W��8`�P���/·Wnݶ�@�_E�?P�a-Ƿ��<w� ~������m���ɺ�c::��2�^^ƃ'm<��<�)�e��mȷ+Y��{��@�}v�1�Mݵ�Ot�hz�X�I�U�{��`�.�T�?ëv�op�>�ȱ�DG�DJ�@���@̬s���Ԣ!D���M����WSwV]M�\����@���"c�:ަ�g�&�X�n݂���+���.�x��s����}��1�
�n��ۼwL���_E�OI7@�wK�_�OOߪ
9q7���mGR�R��nӮ�9:j[����]sW5�?{����vD��q7Jfj�à}��x�o���uȈ��N��=%%�m�l�m����?6��(J��u����sĢP�(\�Z�7m�{�|������.��t�B@#�A�	YVTHHD �C�N�QV��[�`w���q+4�t;j�n�?DB�C��΁�V9�}�	B���K�'�]�t*t�v���4��. %	D<m�}9��m�b!K��������X�L����Aqō��n��P�;�$���ع��eI�ݬK,`��B*n�΁����Nc� �2����˱�ݻV]��>^�|Q	 c�:ެs��}J$<����]�5uJ�j�n=��V5�U����7@�wK��K�E����J�a�U~�_u�X�I�˺^**v�
��tuϺ�����y�MGMYM��m%m`�&�/t�_��t�X�lB����h�R�&����; ��0<�4��k��cm�{��q�G�vY���0څ�[kQ�Ҳ�%�ԗ�߿��u�������${���=�ɩ%�b�t;jӷx��kJ�߃�_E�w{z��u�I$BQ!�����%؄U[�I7��{�,��7J���t�d�k@��K��0�ci�k����7@�{��'M��_E�w���Q�vݶЩ�ot��^ ~���N�]�������߹�u`v�@D!����xߩ�i-G
����J�W���2E��]J!�G �ҍY�8�ħ4rg�z�v��Okgs��'oe��V��L+�I�6�:z6�Xp�`���D�Bvϵ,�]��4�ɷ)�O��.ʖ�5ϯl���1�F9�b+���xu΁��	
��͏@����g�l�1x�z������]���)�=r�.v�Bn��d�:����S�ET��5���f=J�?�����œkg���Z�tv�p]jt��6�L�̇!�������{]������T�]p{���}��x}�}J@�}�������p;�I[��>�6qB�3����Q�� ���Ԓ�1��ѳj��m�]��Y�7�zә/���Ot�h�p�7���#hhh�����W�>�=�!�w��TB!%����f֕S3����������|g@��p�o� ��<�H\����5E0t�Е�WuC:����<�]G:y�N�]��G���V6���e�cV�.���{���_E�Ot��zG���W�'�d4	ŤK��n���v���s߹��>�7����'?!������'���F��&
lSHa�Z��V�D ��׾��7��i�=��<��I ����.���EU��y����Λ	$��%fS���w� �9���UuWSt������΁�����z������awh���J�a�}��< J""!�7΀}�w���=�?4,�L�UTS$"ʅJ$�:�&�^��U�,��OG�3���nv	��������{}�{U����� ��{������$�������7����6�_�m�m���:��۞�����o����(�Rc���Nթ �]\��]p�{��>�g3v��11U�
nJ��2m�
4mНL>��f�4ƅF�����ʷ��2�B��C@����%뾘�$���'�
L0����vY�w�`{Yc����)��=����0{IѨɒ�\�4��͘��h(�(/�3�V���Do����>
b�D�Q'�=�������SC�.�Z|!����B�=�����K$BB�"X!��$3-�ib���.	!c8ؑ1N���:��	�50P�eT[�)��ɇ�K����T���]���E ��iA⡴�����=���N*:����VGh�
��+ҫa�A}N�M=���#���}�S��C��q���m&�1h�U~����'�M�>]��	�r-�!T�V7e�e��{��BQ��p��}��<�9utwZ5�����ϸ�6�Iݮ�c:��y5�i�����s)iߞ�����!� ZC毝��� �����l���u$�Hn=���{E$ګ����uwu��۞��-���@s��
{Wb���wI+�ŠN�{��6���II����7�N��dۻE�ԗ\���Y�IB������?Ssʹ���.�$	 �X$�w8`ux:ț�Ӱ��j��z� (�Q���:�[8�7ށ�������IUsx�)#�����Y�
G����ܾ]I']u�ڤ8fa�n��+�WW3uw<q�4�<�p�o�D(����<�����)U�����@�峀?c}���<��Q{�J���КMYm��I�z��(Hy���<�p���PZI�$*���_�UWz�,wL����zI��E,DbV˶Ӻn�� y���	@��{��77w���� 樄�B��('EHUw3v"��*)X�u�t*Ƶ���(<�pZ��w]K��ۋ78��E϶��h�T�E���/a\+�6${����(��Z�uP`�+�]�}����fywXû�� �ۄ����{�N]�]��w���cs�c���{x�V����O�A���B�{T���6 s=���N�cD'
z3�ep�Ϋn|F3Ʀέ1�[�V���&�m��as����	��
ݏs��trû�뭺�[��"�^�+]�����+����
KrD���n��.��K���ƚ�N�t	��	:d4��񰴓n�J۬N�t���O\� ��C@�镕_��qGY�M�J��շ�z�� ����!A	)3^�pǻށ�q]Х[���;i;��	�� ~���"�V9�x��XU�[��{���镀����3@�_E�OI��'ZR�h�Jݫ���6.G�W�ƺ�7����o���*�3..7\�Yx��;�КM��`�M�;��`��"#�?e��g��h.fj�L��Z�]�W=������b��a����g��;�����o���.���u���M�����&�+�t��X�|g@~�gD!�7ހ�X��t
�˸�wv�M����Np`N�7@�_?U��8�>�/N�0��ݶ��0	�t	��	�{�5%߾O�~�[jWD��۵�!ƞڐ�:�<���4r!1hUn?�_�k�e���ۻv�h��`:d4�8eP:M�=#V��[���lN�X�>�@�s�>�7@�_E��~{ܡ`�D�]M�v�=珋�?����B����# �"��҆��\����Z��M%Q���Lv���X�7ށ��s��۞��%�����C�Հ�+t�&�ot��XU���\�@�镀w�M����t��%N��mn�x\��t�m��i��gWngl��s��$����ny\�.5!7��g�m������? �1�p�o�D%�>��\ ��MK���vKGl��ė}��n`$��߿s@�wK�>�r-�K�����v��]��c}�Nc��P���۞��{��������RUI���m��K0�3��u�>ym�@�1�p:�J}	(�1�7@�F�TV��AN�cI��=9ȴQ���g �}�Nc���LӴ's���^^2��h��rk&k��c�n�;U� ��طJPT�*�s00,�a�*Q�7|��>̶p��zӘ�R���{�:f�3+n�)e��Uvp6�{��P�D����{�Ӡ}�l�B�Q ���S6Ijf�L��*����� �!�w�� ��n�}�)��bM�M5V�������&C@��� ��n��0�՛��f΢h�ٻ�3uv�f�:��g ���߾ӏk�f7�t8< �&�t��!��?���rȝ��h��q֝ym�̝���}��mѮns��˝�n�J��k
�v��V�)�8�nyn.^�Ƭ(���\܌8㴛�vkp�W��gl�m�j���SuIj��"kmGJ�9��M#z�a�l�z=��\v8:L[��ru��uj�;���xv����K2�u�y�G ��.�K�p��.}A�{n��6��V�ì�i)�ϱ;SȲ����V9��߯?���k�##�W1�G,c��-	IwQ±���cUF
e�V��8�nO�4�CT�hE�m+�`'n���K�;��h{�0��Ү�ݱ
���{�|�����&C@���zI7Jtj�K�o�M�;w�wI��>�8`�M�>^�x�]0t�X�M6�����g �m��}>n��DDD��4��.fV�ȩe��M]�ͷ���^�&C@��� ����(�Ϯv��/�r��حîx�[u�)����ˮ��m��X���R�MQ�F�b��]7\1�3�{�l�P�d3ww� �k�şЮ�䬭�5%�~��>s3.!�GaB\�3��ߞ>���� >��خ&�v�$�f-���I�~��}9�\������*T�wT�T���5Vp5BDNn���zsv�c�硱1��� lY�:J��Q57E��z���l$�{����zp6�z<f'�{��ɺ�8�G�]�8�͉�,q��=snWk�H��Q������o�j�[��9��s��$���/ ދ�`��)'I��1h�8ePI7@�zK�$�!�U�������Jf��� �o���u¢��|(J��G��K" �|玁�;Ӏ}�haw4\�ժ�4����؉��Y�\ww�t{-���z��Ĳ��i[�I2U{��I$���ߦ��>���Tn	Ĥv�[��L��n��F��k�3<p��D�ܭ˘p��s�w��:���4�;wI&���I&�/I{���i���U.�Q5uvMU���{�)P��ӛ��7wy�@���͉��k�B�]ҵ3Wwww}��ݮ �|gH��{-���z��(�E\LT��suu���P6��=�|\+��9�u��!v$�$$J���>�)�zA�z�����R�s�R���������5BR������׷�o��y���S$�W�5���;{W��؎'��x<ۋ��!K�]��
Z*���ʺ-��+Wn�	$��y���nR���=�|\��C��suSt)�5Wހ|��6
"CwovzǼ\��{�DL��݉Rl��UU\��������>.I!��z�������i��wI'��@�s������;�DBv��&�TwJ�n��X�M��G�Iι���7W��0s�bC�LP�p�-$똁���::��w�N�L^g����
H�}�{�|y�3��0:�D;l"]�"0���x�M�x.�3��,��\&w�����0�ҝY�0�A��w�γa��̿d>qO3��C��0�䘫@mbah$V F�R��݁3Y��`A	�wѸ�(���>i�+V��@p��{
D�=��LA�r���L��+^UZp���#@+ �+���̘eG����RYKm�n�s*�V�R�`(
�����������K�l�vt��a�tWW(p�ŝ��:���t=���˸�Fm���h�܁�ѭ��b�w6υԀ�)�Ty����ĸ�g���$ڱh�����"�۲x��6��Z@�gg<�.-��J��3u�ʏF��s�^�x9�;)�8g���E6�2	e��m��v�͉ �c�ay9�=1�`3q�%����e��iE��� u۫/���.˓se��N��\�jA����܇5&��sl��K�����;l�]Ϣ�^=�rBl����c{;�v871.�#2�	��[1۫�}�ݲ�I�N��,\!�j�ftu�N\�D�:e:@�Au��ѭ ���la�m�v���Ή��'Y��ǣV�>�D��{G�E�]�D�&�ѬʆN3d��B��.щx�ۗ0"t;f�r�sn��v�P�ϐx��w7j�cl�D�q�;vΨ�n6�gM�ds)5�m�� �����bݠ-u�v�a6-Ȓ��qEЅ�-���<�,;8�sX-�5�2�vu��jY'������=�s�s͌/%�H+R�۞�*�t�C��8��+)�a��pe�e7n1-]+s��8�X�9d��A����a�83ɮz'oN�ғ��;�XN6�#ۨ;i3���v�ւ�Z8R��;7^.x��nK8);4b���lk�#�땝���,��pa�{e���I��,Ph6���0����i�*��I�:���ܾ[M5�1�5"�-��w;�����d{[<�l�Qz�
�wX�[V��Fu����m]e�8�V��0��2ut:�]s���l���d� 1��i�,�l�v6�n�����q=yݯc���ָm���(��6玩�mgJ�*;m�w�:�z2�K��؂�ʇX���ݤ!�+e8��]U�ol��g�ř�[+	z��q�殀+�M�N��m��[�/\��a^ޛ�(`BX��E�$ ���
S�]z���kl�㲉[VW]j�;��ww���*�_:@8 �<G��ʯ���N��@��U_�z@� y�3�Ɵ̓���-l�r�"�S���a��F�:�m�1g�'/a�U��u�e��q�:u��طA;�*\����s�V���D�N�(B�.3.�G�G�jWh-�s������K�6I�l:�<жc�����;6aԗ�5�,��`u��VF�Y��#���--�m�OO��W[!۞9!��s
hC�L���d�\��.ܷ+�uV�F�w0L̜��1J�hn`a��z�����=2Uvݲku�����A��圽��w6X��lm�I�m��@:tx��==���"7�7w�ށ��%�U�Šlm�H�Z{�V��n�}�!���Tis$M*���9=�e`�&�ޑ�H�Z�I*ꌫ-��+Wn�(��7@>���!�}�2��Љ[vS��n�+Wv�����n�t�7�\3�@�ǧ�P'bi�$�D�DnY*���i5�p�4e��Crcn�sRy�.6�G�\�]p�|g@�1�p�o��D}!�ok��:��Rm�s57jfn�à}�l��
�aDG�$)�.��@=�w�>�d4T������t�6�]� ��7@>� �t�hw8`��Qv�e�M�wm�}����>�p�;�&��0�)M��BM�M���!�w�� �t��N� �"wT��:;Fƌݻ{�Y|�4������7^�0@�ch�8����O���������g �{z��z�Gd>x��@r&�?�RX��Z�%�}���� �����N��h�p�=ޑ+M���usJ������;��gӽ�$""c1p�`S��u�\�W�zM��E(.�N�i�T;����!�3�l��1����׵�c���S�6˱�I[�4�8`���t�~��h:"��I,��Cn��ug�s<c�X� ��(�3=���}]����.c�ʮϤ��vƓ�hwO��>^���ݐ�=�p�>�D�QWt�n�����u�ɓ���:c�8~�}�l��(�iЛ�ۼ}��h�8`W�~|�%�����ӿ�WV�����9��p����}/p>�I*����a���d�eRb�B�+M kIi �¢��:@�T�X�A�ֈ�B~���+��~߻�.����U�R�۱�'vـo���)���vC@�s��D����'i$��sמ���\�F�ܥ�'i=�u�;�u�~{�+�ĭ7I�i6���o4��x�vC@�s���7@>���"0t۵r�j��s3��P�M׼\;
&~m�zν� }�8��5j�ˢ�I.��@��V��7J�_�"�/ ߻��wJ�C��H��.���b~�{�@�׵�;����	B���p�3)�UJ�\���SU}�|�p���>����jK��߹Ĕ�xw�{�n�*��[.�1pL�F�
붫��B{l����F�8�1-������8+{�JM�U��'W\�`�;�:�oI�s���J`N������N��0�!,�M���u��-�k\���.�mt����3�ٓ6�m�ʂV/ ����1{J�����"�3�;8z;t��Ƀ���9}k�B��9ѣ����.N��8Kut�=Z��Y.AO���e��;)h����.�����q�r���g�7/D�=�wXvٍX�:�)�LI��`
�N����!�<���;���b����5��]_���]&���@��+ ߽�ty��������2M&fS�`�v�;�Xޓ�tzG�߿%����c��}��R����
��� P��s�7��-wL�~�Q�t�7n���o �y�Z���t��7����xOWP�*��ZJĢ�;��ۨ���Q�8{-�m�l�Cuo�ݟ̳��!�ݍ6��<Z��+ ���t�H��UP�r-�Guu�N���m.���^}���T	M��!�J����{���{6Q!�i:�.�Inڵot�����9��t��>�t�R�@Q��i m�ۼ�_��9��t��>�t���/ ��W���t���Š{�2����zG�oyȴ�Ȕ~�N�*�F����<Gn���hm��k��{��s����I!S���i	��X�t� ��UV��镀{ޕj��MP]�Wwހ}��5(�>y{��1���g�����)-%���Sj��EM]���vz�P�_D(B����8���Bi	N�F�$����
b���HC�Z�Q�	(]��{ހ?f� >o(&�Sn��chM�ŠW���镀}�t� ����ϛ��ݺ������U�\�7X��M�*���#�7�r-�镂]������'eD%L�T�7�غ
�.�4�=�.���n	� ���X�q��v=V�ս�>^�����@��eeU~�{��Pt�i%C�����9@���p��}�O��D% {�AJ��R�V�W��@��e`{�7@�zK�7�r-�%�R�Cwm!;�u�	{���>�7\�e�=�����%ID�0A82�9��$��_ M�s�pwJ�5l�l.�M
�{�|�%��߫~��{�V��M�=�0�I1��ƶ{<�u0�[�{Eky΀+F�ms����-�y�T�	"�N$:��,�dnY�.{��h�L�{�6�Uhޑ��u���v�M��
�f-�镀o{���n�s���aB�#[�RR���RIM�J۬ӧ��ޑ��r-�镀}�:5J��T�v������H�s���{bJ!O�=��n�l�j�n�Qwe���筹�$�=��1�z��|�x�!B�bb�	HA# M��K+	
�C,A@Eʜ�c���*�\����f��VJ�75v笇k���ܸq�ۓg�ɏ=���7;ZQ����ɫ���m�[u�kHv�-�w�ܧe���S��M0��7b;N5��ےݵ�tϙ׬UO�Df�yB���a�����V�r#k\q;��n�����f��ش!��u���8vM��+�%P=���p;uٌ��5�F�g�����Q۰Go�ԓq�"�T����gs�`��N�ː�t������A<���5�J�k>��tm���� ص��k��uˇ��m�\�����	����w��t���P<�Z")v]Kݴ��۬��ON�� �r�g�fc��>������me�����)%�<�ZwL��}�_j�6]�v]Z�w�l�h�2���n���$� ��-�bM�ڵi�Šwt��;���Ix�9�=R,����j�L����m۳��ͣz�uԗ�����v�Cxz�GE��Y��{�@�f+�R-�j��;���Ix��@�镀}^'\T*n�o��k��������zaH�D�.�~ =��o���s����l�^��>�b!L��(ڸ��(�����}����>.#��>���� �3GM~@�Ӥ�s��t��=�t���끱���g�b�ڢ��j���I����=����lB���f�t���z����j[�7@D�+�����T���*�]�e+^���km[��NEir�m�A>�-Z�d�MQ3rU]�>ӛ��:�x�{���!vA���z%�;sV��T��R����<�-��+ ��t��� ��-�����Z��1h�L���M���A��ّV1c$e��fb�'AR����tk��Ps����۲	MN6FObj'@v�2�4	�H��n*&��u�}�jGq�t�M�ch�Ë��Α-�G�{:��dtP��gFf���5�7Xa�8e�JzX#��Bȝ{���2��1�����)$9$Th�(�X��h �:0�E��ahz�L��1C0 B�޶��&h��"j��h��Ձ�����6���6k�B�xř�Dfs!�jN��0:�*'��Hiǵc���i�Ƞ׺��L�������ޕޢ�����e6�!�	�*����OE�	� z��/¿(�(�hB!%���k�{��bmL���DȪ�j���"_��z��� ��㞀{�<k�߮QV[mZ��ˤ�g�E�� ��t��K
�r��܁Χ�ɇd��i�ű�b:��8!�SP�ۍ���N�&����Ϣ�wG�w���H�C��.:�t�t����wG��I�?�@��׀l��T�v]KZ�HM�o ��t�Ix�9�{�<�.;�خĚ.�{�|�K�6yȻ�������'Sy��J+z
>�)(�Q&����/IN�ʺU5uwV���6yȴ����t���^������?O���9��2X����vvڍ��&��ػ<h:��<I��YPn9�{�����Z�x�|�<��M�>]%��r-�AWR�TU�V�]��{��ށ��u�;���w͈IL��k��Qt�\]��M_z�wk�w�m� ���{�7@�Y)n�Wt$�ݕw\J'�o7g����{z���v�hڠ��Y7(�-L�y��f;�����}-���>3�?BQ�� I�
�!H�MN a�iK)��u���b��՟�[`��;k�br�mZ�kqV��F�N=���kPE���dpA��9�l�ב��0��vv"�����Ld����3J���q��@�2��i�xBM=k�9�N�����$�m����3v�˛ۥ���.�@����Wp+�6�'�U��4o9.����S`�cYr<��<�vss�n�g��v ��tp�&�W]��pV���̒e!#R`���n��7%I��*Q�hz�Lɽ��ss=ɶ�ۋ�QX������7[��0�N�6�o�o���Ix���$��{|�V�+n�ՓTT�����Ix�� ����t����wR�V�6�U�ۼd솀wtxjQ-���N�� 3��#j�]�7%ڵi<�@;�<��7@�I/ �;!�z�'Wd��mյv��|�K�6N�h���7���
��Y�����iݗ��ϝ��t�s��9ֻU۷����hò������2��������~������P��x��YA��l�5A$�ݗW\���$��RS0�`b��ዅ�&=����(��>?_ �x��>�n���T�Ze�t�t�{��{�<��)yO���>���Ɓ����]$�����P����=/v�~��tَ���*��6�-]�����)%��L��wtx��M�9Q+�:g�ݥj�0Px�{<[bQ��ށv��A��X��ʼ�z��R���lP��[ed�Y�.w߷��Iwtx��M�>]%�}^�H�VЮ�իj� �tx��M�>]%�=2~�C�QX�۫i�x{�7j�>�5��T�F���\�|� �tx���d��[���ݥot�7\�ό���5D%/1��YFʙ�E�@�K�SW|�ό�	(����c��w�{
p�*��.�cv��.ݺ�3��],dz����&��]����њ�)�����I���V� �#�=�t� �G�o�d4	^������;M$�m���n�I#�7�2w�ID��k�*�Uu56�d�Uw}�������۾�{z�)��E�c��mRI��o�d4I�w���~	L@�)S!i}�?I�./H���P��j=
>/����?��Wnһ�;�w�h�� �ُ� �����5DBI<{������wW:���w�y�&�5�B�}-���p�E���󜽒WQ5�m��������<}�!�$x�T�.�����ս��<~�d4�� �����%�Tj��gU�U)���c� �eX����ٮ�_xR�Z�]�ҷ�hI��M��<~��h���m�6�x��7@:H���!�$xUU`��ɘ30���m	zOÒ��j1V�apۇGZs�s���aܾg�h[sa��U�9E��ȗ�{n1���kH�:�r96isĢe���gsuv^u��g5tk.����Ө�n����"�K��L��%�i��ۚ�l���&y�OF�ղm�ݭ���7GX�ìp=�d�յ�)ڱ�\��!��fbT�K��`��r� �GS������C�YJ��U�w3�oe"ʨ�M&˝&9�$n8�<��3����$�s�������3��۴�[)�+��T�ߴzG�o�� �#�7���Ri"�F+-�j���~��hI��M��_6!D�g�$t�jꉪ�.��àwo�w��ޛ
d{�|�c��ꉩsS$���77W|P�S���� ���o�솀I#�=�F*�c�IX����t����!�$x��ė�����v"��2�i2�X�+�z^;���r�%kHt�/c�BYଅ�����t�QI4�]��}�3��	$x��7@$�����J:�I;�v4��$�[�E]���������9���ϻ!�O(��t���v����7�� m�ᰒS?y�i����?a5-�v���m�t���vC@�t��������t��Eԫai�j���~��h.����n�{�<��٭R&`ҁMȪIUE�6��Qu�:�:Nn�sɽ����*��������#�6,ݵy��r����7���H��ݐ�%qj�YqZ�ۤ��x�� ߽���^���I��j�f�\����w�;������@-H��3
#e���^(@���^�I��x�໔�iէw��ID��}Ӡd��p��}����	_x�(��R)�]&ս�@����o�׿|��|�{8΁��2�Q5u4��λ��=Ih7nu�5���z���XY�cxy��[.�+WM�Cwi&�������H�}��h^��	=\����WD�%�����ẅ́�d�c�'7k�w珽�
&O=Ss3S�WSE]�ʒ����Ɓ��/ ߧM�zG����	]:Ct�؝����~�7j����u�3�Й�!~Q�3=�{�q%�����$VZ7e� ߧM�zG�{�vC@����N��s�C�������z��v.�q�;=��a5v������"��c5�9�e�+{�� ��솁��/ ߧM�9z���jl�rI7j����Y����9�\�6��y��މhv�R��2ӷ����/ ��M���Gw���;���Z�,����Cwi&�����M�����m�Cb�f�p�2kj�WN�M��@=��s�h^�[��y�w�]���j )�|O	/\�~V$�b �E��$S�KL��HP$�@�E/SBѤ�2N�,�2���h�)i�
)�`�������p&�rĜ�2q1T�h��+ɨ����g��bn�Op�f�ib����x�]6)7P�ah03,7b��R��	<��Mc�)b,����hK�DeV��`,�U{�gmFU9��f�T�a�����̰�����:"`!�`���"�z75�J	�"AN\ǘ�C�!��o������5؛�Y� �&)�:�p	u�Є�IXV�Y
m��dy�o���bf��:D;��ab*�2{#��QID��jGz:��ؽ݋_@t�W�:	q#Z	�f��A��)���e�1��QF�"�h�4G���h����Ε|=����UV��0H۠�&I��С�{ӭh����]�.�5��׃�n�$�/`�=�`P�>vN�[m��k![���W�$�m���iZ.�z��zvsɇ�`3�[l������r�Q��;:T�u�pA�G!�V{�u`�A��D�r���fӸ�vvq�Ƶ�{ng��T�����1�cx���l��b��-9��k&9����Q;���utj:�t��$�+���;�qafple}�'���ˎ��W�5��;�p=���숶t/�ը�n������YscQX��m������=�{6N<8δ�-t
��;]6�2��7<�K��-[`z'w���G������X7�;lP-�9�)�E;c}�U�s>oip�h&����л��nנ8�q7-����f��mc9N�p��\Hs��5�k!Ի=����]��k�ؗ�z6X����L��Y����E���3��p+��ڷe��Ȗ�3YK�utuYk�j���8�8^M,�c�vӐv��.�n�]��l�s��v`���9�K��u$1�� ��(�QUݥ֝u��%�%��nB�N�6�/6�^pʶ۔��)5�b�֋ q",�"3b���Pz9��pRi�f㮖*J��K��y�,�]�6��u�F����]%2O�����ݗ� J�s�7��Uv��]YV��[�'�����pgfv�Q�W5���n�a����L$:��ݲ݌uQwb�d������������/cWT���Ƹ旣����I�VxٶR6����\X��iy�I�DQ�֮��;j���@��8�4�<�� -G��v�]M�����^MΓmvg��^u��X�8N�a.6���M��U��n�[�&��j���a���w<x�WEd�GkOhdm��z�nB�N�A��<���)��6p�*m����2 Fwbw2�G �ي�=�#]E=�7]�u�62�����S�M�ek�=l��c�{a
x�[�n�R�6�t�!�����َKm��.��/]m#vu�H�Q�k��Cjκ�p�h�;�m�f�QB�H�a����7���O�:z� أ���Ҭ�"�#"2$�b��BOh�U�| � ֳyY�n��׉Ƒ�f�ywT�\R�S�b6�N�n��w�/���^)'H�X�$�;gv#6��a�9s�-v��G��׃��\��%Ѭ�쎓F���ck���y�ͣg�M����������^�u۠�ѳ���v�"^�a6�;�<kp=�\"p�j�1����Gf�m�����Y�l԰M�o&�H,���x��{I=�L�j�L�p�&}�������P��ڎ��TV�H2��ͳ�`�vwj��m.=bnո�ݷ.^�)�ܵ'�p�>�@����}�&��#�OpF�7E��wcY��/Ixޒn�{�<��"�%q��ԷWtRv�v��zI��H�w9���/ ��ъ�6;N��tս�zG�{�ȴ/Ix�$��֎�6���$��SWw�=�m�@؅X������y���1�3[j�R���J�f�7�g�q�PӶ��tj6-��Iص�6v�]�wC�:/UMX2�o/������I����]���vz�T�M-�R]�7Q��ַW�s�ￄ ��QN�^�>x{�E�y{��P�p����6�Cm���#�=�r-��/ ��M�=ғIGv��;mڤ6��s�h^�xޒn�}� z{�4	Ӣ��]Qs�rz���lB�f����u��9�*�Ո�TV��۶�Ӄ�.��qq>ݵu�to��[�����}��kYn��J��V� ��M��#�=�|f��2q�pf�L�Z����t�m�}����=.E�}�M��}^�uD���i!&�[o �t�h��t�7丵BP�};^�{�����D�Rt%sAeM��xt5$��m��?�����G�{�2#�KW-��O�k ��M��G�{��Z��=Is����$��r8�B�Q	^�ܜ<�8Q��x��v{mӉH�E�����Z�|�6MO]�m�:��m�w�<��"�>��`zI��)4�jݷV�iR��{�m�uDB�S'��� �n�z��|P���Zt6�۱��Z��,�F��a%2<{|���<�t:�AAM����I7@;������~q;W�z/��wﹺ����p�5uV��tս��G�{�d4��X�$�zD%YEQI;��n�V��My�u�aWV�n��pr��u�;t�8�V�q�3��]��C�t]��{�d4��X�$�ՠ� ��"R��c)X1�����,�n�w�<��"�ꪪ��;SS�r+���n&��y���=���9����=���M4]���{��G�{��Zގ�������;��B/���M�Ҥ���{��Z��g �;��c����G��;��n���g����m�w��q��i͵�S��e�w9���
 <�(<�ա�s��ӹ���P��"�]��N�nW�s�p�&yc�wh�⢧�`*m��MC���Ѭ�(�ۃ�l\:���ǫ�wۀ��9�)���u���v8 8������q�]��nj�(r]�³�c����ތ��e���2E7���9*�rEn;�2�%���9ʂ��{k=N�u[�ݹ��i�8�ݍ�F�=�l�n�Z�5jd�*ҥ%%��Ԯ� ���>�&����w9�߽
vKuaW�۲ն`t�t��^�ό�{-��S#�c�j�.lV]��{�yt����!�}�p�>�&�WZ�m�I���Eۼ��E�}�p�>�&�/t�{ԉJ�S�5v���>�8`N�t��^��E�jJ""u�)H����m6D�Yf�i��y��M�s���n�-��耠��H���*f����{ww���:���~A����?�����m]�m����kz�(F�V�O�Gi�K��Ym�@̬s�>x�zy���Wv�66�*�x{��@���a���^���۠yt�� ��#m6��5��@���`zI���/ ��"�:�D�(��
��m��I���/ ��"�>�8`wDQU�(N�0��
˭�q�)�m�v)9�v�P�vS5�]�q�B�*챠�2�M���{�|����r-�s���7@��.��:M$5n˷xw��@���}$��O_E�O�"R��cJ�5M[z�h���^s��}ݟ
��Dv�8@*e��$�
DG{��g�wv�g��]ML��wvX����$�/IxwL��:�,��T���ի@�m�����d4	��`I�tT��R�U�G1�$��l�(�N�:�q�����=��B=Ie�n���ZJ�!ҵ��L��:�,��7@��^ O�Etm]ۻuwm:i����H��0�%��>0��wb��W�鍡[m`wM�"���w��Z��1fb���mUU����k7k�<w�=�c�_
��(��|�@�Oq��-$[��n��r-u�X���@s��c�)¨��U�ʹ �6���v�R��[�<�Þ�E�6�{s���䝣<�n3�t�b,N�o^-u�X�t�ϛ���7��= {3�5;W%�SR��k �N��E�/ ���h���;�"�q�i�v�Cm��^���u�X�I��)4(���m�R������{�:�{<���9�ޢ�6��7j�WM^a�N�� ��}�����>3�5���2��OdV&�ܛuc��Բi��7D᳠{-��
7��O��j���&)�m�����8Gc�۵��C�͚���]�Fw������k{x��x�M��ְ�v��qԷPc� ��r��M-l;(��S��/��pgd�j �ö�3��YҞ!UR�k�U�D�];X�z��%��g��{>�sΜú��5�-�i�=QK+��������ڠ��1��#w+�Մ�V��k�9�p��&�ϟ��oK8�=8�s��G<mj0�;o�����;�������"/�5����l����Л�Wm�=r,��"�V9�<���(��=&��JU]]��� ~w�=�c�	)�k{ށ��� �z�)]Jc�����'_E�}�&��"�=�r- 蒊�X���Z��m`zI��Ȱ{��@�}�yD�����v]]Г���gf��ݰ�{z[�W8ss�pha��Ln�;�^�5���5t݉i���Ȱ{��@�}����{ғB��t��n�;�w�{��s���Q!X �B�ʤ��0��(�����3tg���ϛ�jJ�n�ڹ&�]�VӦ���?���}�M�'�E�{��=Ɍ�T:�$,��j�灱
%����7+vx�[s�V9�b�)�2ݕn�;@��=r,Ӝ�@�}ޒn�޹�����e�J�trSۻ=.í���ikslb���>�8e୒�mgI��-+B�vݶ���E�N�� �I7@����*Ԧ:,N髷��:�,�n�=r,��"��(�厝�ժO�v�����E�/]����i�5����	F ��2B�41)���?:���E�aQ��wW���)ԮHDD�d$�JA-2��W8�[l�y���HG
(�.�
�E����F� �4tI�G���L;ІIA40���Da�Ѡ������pDDa��l�`�I��X��,���I0\8�tFd�Xf�طl�����̎ef�^�
&���*	B`�&i�-F��i�fTPVY��y�u�2l�i�gOZĳ�#c�QT@T�FFDQnw�:��3$p�2�&�������J֘G��B�4�3rLܒF�kTE�j:6��n�A��v�B�kD��H�Ʊ#�gn]��fZ0�sڠ`�
�*��z�_C�S��aS�dN�_DO�%U$@�]�SJs?z���=�������'j݉!���/Ix��E�N�� ��M�=�N�Q&ۺ-�j�ݻ�=�r-u�Xޒn���ޝ
+x6�Ϙܘ宵�`'n{h��{q���ɮ7�'s��r~|}��� �Xi�}|=�yX�y�}�|�lB�n�g�b�s&� ���I����m���)�g7k�cw�=�c��,�aH�����P������E�N�� ����|�t�⡗b�M��X���I�Ӡk���>��z%
�	DS
)B�$�ae]*[�ֿ~����%u�LtU����{��:�,�n�=r,��!�}���괝*J��vEM��l�x��n�q!֜�j�����8.��4+Wl-ӻ����k ����O\� �t�h���'�ȵq��U�������ny��1��]=��~���� 0m{�ō��ܵ	�++�����t��xj��)�f���nV��OQ�v��m�۷C��@�}����E�/ ��d4TԢ+�*M6�m��}�&�zK�=�u���]t$0q%��X"H9���k��53���F�K�t=fI3ֻ	v���nf�e��˃��D�F�N�GN�c�������lB�f��V�\�\��e����ݶ.\t`2�n:t{[m���A���;	�n�9�b��7��y,���p�n����HR��O+���ծ��	V�����x��u�U�u]�"q�l��Hnqe�u�6�1�����G�[�F�u�X��{����l� ��dJ��ҌhV[J�HVl����<F��iٜ���n�En:ܵ��s:�.�:�n� �c�:��<�m��|�t�+�V�i��wL��:�,�n�=r,OT��t1�V��������I��ȰwL�@�\�9.˪�53jj�x�DD����r�g�{1��c� ��M:��Hn�&�{�O\� ���'_E�}$��t:aG�]�cT����М{Lv��ʚ#�z���wZ;u��v���O7m�'OI�mQv�v���!�N�� �F��"���< ��=�-U�*����owus�}��@���!=-�����"wt�h�v����,n�۶�	�&�zK�'��h���=��j�
��WE\���z�B���ݮ���:��<�7ށ��2��2�R.�m���'��h���'t��O\� �D�:����]�e�9���)s�l؍�A�⣐N�8���XΣz��M�T�,j�V�p�'_E�N�7@��^=&C@�H����j�iЪ�<���I%
dܭ����i�V9椢ɾcU5�%Y!$��z�n� ���t� ��8$ %p��NC�Q�=گ�<ws{�=殤����UUsr�j�x��w{�@��Ӏft��Ir, ��� t��e����0��g �c}��s�>��΁��߿��ܣ�����nq���n��Mƶ�z�������>�*�����i�1vU�h'���I/ ���hG��B��V���fj���뚡B�2y��woN�c}��:S5�,�R��˻����tݳ�}���I/ ����GMS(��j�{������i�<��z��p>�YJ���Ҹ���a�A�w�s��v��Q+hlv�V�5l�>�t���t���$��(���-'����ReE�T"4�!jCe/n��y-M�k]��A�t���ˢ�_�X��ot���t���$�I�t�S�KcUv�wWwn���Z�� �:n����@�[��lw��@�[87��6"IL�����og�y0�]ԷH��tU�l�:N��Ir,�s��P�wy� ��T�Z��7Ws3Wހ�7<b{�{?��� ����g�	BP�!�*nj�B����)�;[Q��*G�۳�7:C@ӎ�ܽs��rr��s�<Im۱�6���(�<��&�b�y�����]��[�7e����-S�Zvݛ�$�qk�9�"�/m�9�v��:���ч���Z-���BiE.�,Y8�Y�;����bn��zø^,�d�˧rn�����mO���tv1n�f�x�۰����OL�m�d��)D/W��Ͻ� wݻ�Dƞ�b��q�7a��F� �ێ݁���'b��a�R-�V��bM���e��k�$��h�g �x���(P��ݭ���Ѷ�R�Eʹ��|��۶sbd�׽�������-��%%-X���+N��`zM�$�'>�@�8`�%��ĭ�m��$�'>�@�8`zM�>�L���1]��Z�k ����$��I��"�??�~���n�0���cYƥwN;ywl�;d��A�^���:�F�s���|m���j��f-H�N���E$�z>�@�@�]�˴"�tU�l�'zMޭ��؅�z�p��6��P�ɾ1�m"UZ�%M��U_z��� ~o��$��I�/.��e$+T:����?;�=�l�<�z
�n�p�Ѷ�b�R+����zn���}�[u���=TBP���\n�K�9wF�F�y���n֧����zV��D�n��x$uա{%����n��7M� o/��A�e�ߛ������l@�m�˹0;���@�0	=&�t�\.�ۤ�����Xyx�6�<�I� @�%	D�HC@�$BH�PJ
EH U@�J�JG"��u��7X����!jm]ۺm؞f-H�I�7@��/�D(�Jw_�@x�T�lԒUݡT����}�齮�������q%����#��;]I��rH�hiFd�
�������m&랰��>^۫�؞��=v�;b]ի{�r{��Z�8`�����u��V%v�;N�n��E�|ݳ�{�o�'1�5(��5�N�m\â�M�ּZ����oN��r{��-�Ғ��lhwt$�f����d�:��^9�lBK�K鈈R�"!8���so�p��E;��Kbj��˺^����p�6N��yWTPt��l.� �tRi:�^����gt2)���=`�@����t��݊D��	7xw�E�}#��t�ꪪ�R^ }��M���];��b�>�� ��M�9wK�=��-���\M��j�0}$��t�ޏ��>�� ���UԫN��*n�]��9wK�>�}����7@��]r�nЋT;N�n��E�}#�ﱾ���\���\���H��%V�5�ã;tbɚ���졊g	(/]�X�h0�Y��fi�&�[s�F�p*H� ��gfj�4�����yz�������E1�QWM��m���WgY����89E]:��"-P�9��6�
j��Y:�PMMS�c:�#�$	�����9J$Ƙ��,�ة�06e�����"�.d�A�=j��P��:dN�Z�/�9��{�ѫ,]'
��H��9VdQ���:"�%",�`gi@d� ��=T=��T��1	cD�GPw��0³2"�
���/STGV:L�0��o��@��a��rW
&��5�{{�^�a��u*=QJn*�33؞�x8�ǀ�&��	�'q��c�gQU i����Hn�.����}�2-K'�?���s����uR�=��}��cD쵠�*��U�����;^�-`�]PF��bF�q�;�>6�+!����p!/��ݞ��d���7=v݉�]�'���$ ݀��T�v��8l`��;Q�,�p$��r�\� ����4�m��V���&s���&��� ν��t.ۦhnf{b��v�E|�ɶc���*�z��&�!���.s�\������W+"휎�9༽(l�.�0&65�4�W���@��C�nB0f���VeNm<;�`��<��%�eI�CP�F2�Q!�"Bx�h����ѝ���b~���/n61�2��+�`sͺ��j����lks��v�&d���3�Қ�#H6�sq��c��c* ��N��f���#��A��7N���'�2=��z36h��ޮ�z�.6�,o]���i2�r�7���pE��z�x0�� Z�LX�;��w5��k����Eu�`6�Ѥr��m���s�-��=�������UNR�c�r�X:&�lQ3u�a1�kov.�4X��yk��Y�C�Lv;.Ɯ⎹��y0�+�m��n�NI�4�i��(��OH��N�ɪ���5���]��x��z�r��[����Uf�(��`��2O�R��u���� �����i�t�)���ghBwc�j��l'b��,�\��ii�	Ƈ\����sm�c��vg���zis)��kd7o�r�lqc�mR	��d���C!vܺ�}����$=n�:mb ,�:gh֛A����.m�at��n�3�v�����:.�O��y�+Y�`3ۍ��p��7j�p6�;��93ׇ��m���/1,�9�G��lnݎ5\�\i������6y���댮7+�7�v����<q��='1�<Y��%�<ژ4	
xXD���1��;x�jj��u�`���)�7�صeݛ���Km�K�ӫ�;�=����ȑ�u�6v<�%wU]����r��FSrFvɲ�y�}l|g���m�l�1�x�Z���3�\�#�Zۖ��N�������������Da�@� �4(v�|@���1@ͫ��K޿��������;TK[[�	Q;pIF��i,���N�iT�E�.�7c=mΧ��j6&�mY��L�f0ے
�m���ګ��vq�Qpkj�KpN֢wq��l�6��2n����}D�ێ
����Wx�b��,]��[��l9�L�B뜉���x���qm�n֜�㎍���Ό��"ʂOnM�qr�۷g^4��2�n��$=��_i;�yL���f���AT�[bc��!
V�oQ���Oz�f�^,�q)�<�oj�Fܛ�I�e��?��0}�n�˺^���/JJZ���CBtճ ��&����y�9�7l�舙>��Um��-6��"����E�}#��M�>�L���e�e�n��E�}#�亂�r��:[����N��y���p�=�I�.�xޏ��:t, �P��@�G�)�N�,ON�Wrq�턷�}��8�|7>y�W�����F�tRV٠w�������z>�@�GW�qWR�5cM�+��.�{����ɓv��!M��(�H����g�=�g ���{��&G&��n�
Ҥ�;��=��-�0}�n�˺^;ԉJ:iկ�Sc����6O�y� �=����\I$�ټ{='5L�U+��tLڹ�8��7@��/ ���Z�8`������NW��Ξ�0gs�+E��g]�����t=�cj�{�/}7�8�O����	_��o��u�;�x�|ݳT$�!�o{�=��?��V�%�M�5%Ͽ_~|��0l����3��zNc�j��֚���Z��WUE�9��ݽ8����"I- �A�)��z�s��T������Ww�V��V�� ��&����z>�@�GW�qa*�ꕓ%�)�����\a$�F=��~۷� �ُ���ZT�t�����;��5�G<��͸��2:�[�K"�u��0#gj����6ӫV�۱[�}E�}#�ﻦ�wG�N�T�p�;�֩��׋@�G�t�������IK��cT$�'M6`��� ����E�}#��ԹZ������SwUwކ�-����{=��ۮ����1��i()pΥDv#�����<��&:EݕWe%I&�����p�7����$�{߿$%���%m�Kr�E|��p����.�ܵ�l�bdae�1GS)5�Kv�RR&�Ӽ�Z�8`�M�� �s��JZ�O�V��VـoI7�DD$��6��7og�|ݳ�5�1��wc�j��wG�}��-?������>m�zتg*]��5!sl����}���t� ���w"�+�lVRT��kŠ}#�ٍ����|ݷ=�DB��vߥ��t	uP���2��F��9�6T��"�ݙ�r��2�m�S�v���D�볔 �޴.���1[m��s X����W�M�n8&�:�ns@�9�Mƻ�%�v�ڷ7nQ��'n�����r�.��Sp�T��W X�������.m�4/Mc)�6;h뮹�2\�L���7�@r<;^��C����V���J�kő'*nT�*��W�< y�0˲$�ږ:&��rA�����p �J�����r]=p�\�]��c@�q]��t���<��7@;�<��@�G�EK�������j���ݎ��
�=�{��=�zp�o��J&Ol�5UuswA*fn�{v�g�|ݳ ��7@;�< � �$:l��iR��9=��3�@31�aB��n�vz���ڭ�q3WT�SWg ���@;�<��@�G}ĕWE+0���<oSƻcc+�\wmqɭ�w���h�`9:�0�n;���JX�̸o�Ͷ���� ��>�� ��7@���r.
�(ڶ�%����_~|�fd����OI����O"����j�
��x��p�:zM����RD����9���(�ht��jН4ـt�M�� ���hH�zu*�j�j�L�����������>�� �{�n�:L �]�զ��!݆V.�-��72��Mqq˳�@\����E�m��m����wn���$��:y� �����>�3�a)���������W3J�tnޜ��}�f;����=�ZK���V��Vـ{���w��w�E��K�]��2p�@2Qq
:w��pg����ɗ%�դ
ڴ��wtxH�os��wI����E�"��t�-;l���H�os� ��&�wG�mN��AUp�ë�aW6�����6��z�)���8����,6���WJ�]	��cI��@�G�:n�wtx�>0N�\��ZC�v4ـw�M�� �G��όޔp���v��$ƭ�wtx�>0�|`��t��R���Wv�������S��3�|ݳ�}���u��,'��4	!&�J#�#�}�� �2��ʻ&��3�)0��t���$�� �Oy�H�q�5`�u�<B�dMG)�.ބ�u�L��/=<�����D�����^�nU�`Ӧ�wG�I���όz�uډ'nبVՍ��� �ώ��Àcm��'�*F��-T�ۥv��#��ό������]J�]��cH{���co� ��|��Q;����KwRZ�S%�Lݢ������l潾����e��?G��%���R,��.˹Mqbn�C%*�YjD�q� ����軮{v�+m��í���i@�(��nU��mf;6���c
�^���o�Lc:����H�6�Y�E"B��gN 4c%rŸ���eݍ��&��{\��0w�|��ʆ�Z�C�����i%�^�t�\���^י�ǃ SOv��Z$6ܻ�,��p]=�i��\�&�9�5?��Θ�o$8�n���=�z�kFN0<77A��nM�&)n����ػA�b�&*��ۻ-�$�������<{����Ӻn��Qk��[m&�
�V�;ό�s� ��7@=:<IzR:���c��z8`=&��G�Oy�{�.�%��V��J� �:n�ztx���~]��?��ʹ]ۺj����{��>����w�M�2��I*�=�OEnl��М`9O\�����<���n����r��m�`�ѵ���k�m=|0>����ݘ��<��WR����Z�WY�]��\��_GH��!A�����@�� m��2�v�N�C��lM����۠yI/ �ό�ό������aB,���@�m� ����Á�q���҂���J۴�`*wv� �ό�,o���w�%�\ �,�ME��C�n];��r����m��rv�Y���^8kc�iVO�+j��x��p�>�o�%�[���g �tU.����[f��I��#�>���=�|`x�Q��t�%mX��zH�9ξ�>or��w�u�u ���T�����fa�|��Q@P4#��*P
�&5�oӰ���<.��_��N��[�#�����A����u�o�ڬi:���Dl����}4a�A�
Gf���5�����R���қ ���-���PT�f1Q��) ��țB�v�cqi^�n���ʾ͛�h�� �<� {{�l��
;՘�T�*�1��j:��en�Y�gkWK������L�TU��I��k������M���	'�}�P�G�}c%�ف�]}�FZ.�Hͽ�a�D���ު�${�tIAYkE]�m���/�����MM�ŉ��H3Iؽzv����N�0�N����*�j�x��F���= 1B||�-<��"��s�L@�!�G3�TLo���^���8��{��.���E��:}D�_U1E>b��"O˂x�Ggoj/Gi(���E��eH�)B�"�4!�H l~��0�I��)4\lu���tջ�����^���C�(���ݾ��H�����Iڶ4�ntp�=�M�Iӟ����/�v�����ګ�by��Px�gGp�2��=Z6�K�lT�ƭ�&�+-[i6`�M�6�y�ᰗd3��<ѓ4V�J��X[{��<ӟ�όѷ��%2{V�Ң�䛰%M�]���{���=��< �DW~�E���Ӽf��8`��n�t��~���c_��c`��6�h��"qLٽ��M�i��R=�;5�A��g}��v������m]]�`����I��ٗ� �J=�Ɂh��w.G�Ӯ1��;�ԢhX�gs��nܴ����؎�
�2�
o���o�������峀{2�Ԓ]��c��j*G�ur\M).캻���g5D(Jd������I�A�ԫ);��ӵ�h#��{��I�ǧ��W*h���n��J'1���wo�y�g �e��1<XL�L�T�X�{�$xtp�=���>��IL33���f{����̄�V壗��=k�c"rd��`,N��v���z��!��v^ݚ��l@�������N���u�n���
B�y�7Sr�2fM����p�rX�����'�#٘۲�W.^SY��5��nN|u���Ҷ˅{	t�8��W8�.�D[<���GF7Q�wO�|����n�n��p��ݘ�^��"�b鶜���
w�8�l�Ӭk������a�e��|V�JT������g���1qv�,��Z8^�K���Y{Jp�Dܶ�IJ�IQ�-�K��_-I}�8ٟ���Hwo�{"�&��UwM+I<��p�7�&�I�t��S'�NKT�݄�uhD���>y�� ����L����;�ZWJP�
l��m�zH���V�s� ����}ãi�젵nӶ��t��=�|`ޓt�G�oz?U���b:�h�[V�A�G-I��P��k���u�IFB
��)R5aY-�ė���0�I��#�;�X��cWY��Y����uw���}����$��B������|�c��f^꒠��m
�Ћ-���#�=�X����wM�>���$+t;`:Uv��=�X����wM�N� 7� ��wm+I<��0�1��x�{����DD/���Oo�=i]��������W���nsn������y�����i	F��B8�R�$�tB��ԗ�����:<�镀{���'t�"6�V�۵wot�G�}�X�ό~W�HR�%ܧc�?Z�����=��l�^��_[��>0��MhP���]��'w]�s����:�ԫj��ok@���:n�t����V w/]��cC��bvp���@Ԣ^����=���^�����?WI�Dd@՞�(cv+=��n[h۰��.-����\�e����y����vE��� ���}�+ �y�oޓt�w�t;i�]���L�����zM�� }<�v�I۵i'��t�~�M����e`]\��W�Гv�� ߽�t+�}ηW��͛�A�" �)JP�E���""�(�S���*�@o߼��usϸIUNI��V������ ǎ���=�����;��{�6Vҭ��W7qRq��ә5�;rl�Q��s�l5������q<L:2���en���ƙI۽�?����Àw����G���\=�)����h�v�V�k@�s��wM���t����U��$%֣I�VZM�� ��w� ǎ�lB��=�����>Z�&i�\�Z�(���Ca%2�������=�|`�M�>��!�ح�:Uv��=�L�����t��:=Iw���O�6��
K$�+�qԌ�	���nu[=�%�d׶h�9skeݭ���!��Sgf8n�r:ra�-�G"�v�{b�R\��ԧWn�xr�wmT�%|[�+I����c]��]8�J'�<��.�����v�lJFuGc-�78���6-�p�F��v�;rb0� v� �َg���.�Kl�O[4#D�̹�7�c��g��z���&�U��^QNe��!ɇ/8�1�E��0�ֻmg�KL��ݏ\�v
��+�}r��D2 _w���������:n�t����V��ɫE�ݺ(�l�7��t�G�o�2�w��v��I;��[v[ot�G�o�2�w��:n���A:���1;����V��� ߧM����WR����t��U���:s� ��z������~(���4�ws�c#�^�3��L'��uzc����;jؗ3��\;v������.N�6��}�{ހc�|�c���^��d�;����*�*j��x�Q0�
!U~!���&!����$HlL@S��f\מl�\��0��M�:��[�l�n��U�o ��X�ό~�7@;�x�-RPjГNդ�V��0�t� ���L���ɫB�C�j�[l�7��t�G�o�2�������5	��\�<I�J��5l`�[�c��e������Tk���йBpN���� ���L�����N��},�CTƁ�M����V�s� ߤ���<�Ȯ�p*�wc�*�������6��J�G� Q
T$,	S�H �R�����^��6n��.K�Lhv�Z��l�7�&�t� ��X�ό�)Ewq��ƚ�,���t� ��X�ό~�n���?~����4�"�$"�Ip�R���uk���v�8��kp��<�^tn�8��f�VIv�J�[z�?������&�t� =:+HT�$�ݤ�V��0�I��#�>��V��C�_;O�v�[f�I7@;�x�t����;�wW��:6�N��t� ��X�ό脿:�J�WH(��	j��LA2�A
����>��{�<�C���Yr�6��=�L�����t���_m����_�;�۸�ʭ�˒$絮���v ���u��h���`ۖ�[=x����ET�Y*��_��� ���z����L� ��_4�К��M�ـo�&�t� �镀}���=:�Wwq;�j��{��<�镀}���7ޓt���Ymҷm�ҫV��~�˽?��H�o��n�wH�Ӣ���j��.�fo��y�g �Q�n�U�ߵ�]���7V����XR ����U��O�炨?��oz��*��� u��T%(Ds�mi��?�"(Q�/��'���?��~���W�:�/����������W������?O���9� �*��_�������U_��$Ab�W��K�#�����"P�(��������_��_������:�O������y�?��w�������B�9
$B 2�J��J����(��)��(�)
2�J(�B�0�
%
%
�H�I ���B�@ʉ#
$��%*$
L(�B�2�I �
$$�������
$��*$�
$�"ʉ(����
$�
$�J�)*$�*$�"K ��D��J�(�*$B�0�L��*$�L�(@B�(���J,�����(�,(������������) ��ʉ
 J� 	*$�(� B� �B�J
A
$B����
$J�,(�̄�D�@B@@HH�	"�����(����, HB�$��!
�BB@)!�!
#") ,� !+! �J�H$$2@I!!)!,�$�!!"�@����!(��$���*)"H@���H�2�	(�! H�HJ0��!) J���$� B2	! 2+ H#! !
�HJ 0��	��@*�J�@�H@�!2��J���*$$*�!***HB�$��+ @
�@�HH�B��$�!)! @��*B+ 2�	 L����� +J!		 H��B"�*2�B�B��(A AB@K R)0 D!0������B�@B� B�J)��B���R�2HH���H$�(2"�H������� 0�H@2 @����� J���0�(@�! B2,! @��J��Bȥ*��J3� ĢJB2J3�" )# � J�*J�$�����������*����_㗗�G_����~U������G]?����������_��g�"��G�����g�ق�*�����ߢ5�?�DUu�h��PEU��k�?��3;��^9��Z::DUo����?����DU��G�?����q��u��*����*����:5G��=f~3�����������?�=�[DUw�xY����y�~�("������{ο�ΑX��?������?�������)�¶����hl�8( ���0��  }5u�*�C�Ȃ ڛf�
���{��  Lc��5k !�E�[�}g����A�P�� �6��wp��Zt: :�:
�
 �@u�t v  �  h ��� �����   � tor͠h4��(���]>�}��#�È{�s ��cG�yC���4����]����{�9�#�M�[Q͋�@�\�Nv�ww�}��|��]���j��U=�����:P+������Ý�{�<����  /
z�[��J�'m�w��G���uk{@/,����R�R�`���f�)JYe(
]�t��R�c�=n�e)E1 z ́�  )K�r�
;2�)���w�,�Ks�(]w(�
t�n=���ҔR�4�;:J]۔�Q�w(  4���L � ��u������^P-�J_{�v>��{�p���5��=͠Z��z�a�ӻ�����u��,Ͻ���t�@0�����xy�ڼn�{������<Nv��[xmAf#������@�=� *�h �|�^������@��a���󾳦��m}�w����m��;>�zx�"��À b�w��xz��	=w������|�__O�M/P{��͏����s �  �Q��Wv  ���ׯN���k6������`�s �WM7����M�!�{��}����.��ޱ��P�������}���b݃�1�1����}�=��n�xۓK���6�a��     �I�mJR�  D�*�*�ͪ�  	S�ʪ�h��0�L�@�����کT� �?ѪT�R�H���jR�� �x����?��Y��������χ��_}��TU�.���E] "����
����*���TU���p=dI�|�0�3{5
�#[��/����BHM���K_N��s���l̵��W\V�(�V��Z�N��
(:^!�S��y�o=28�+�����,�O=��ߣI�X�����'�r_��]���,�,<%�<I��#=��1�O5�NlNm��8�$H�#��`ˮn�����<0�r������g4yu4x���Mıfh�߷۹�v}��w��)P���
)�������k��'�.�%�~�)��^A
f����d����jFF�y��zB��z��2��B�ap��}Y�EP^^�����(�S�qv�]�p�_[3[�]�����o�CG�HO0Ԯ���U��[�gk/os��Lo(>�U\�Ū�w*���w���K��V�ǥg7�n��!�eԺ�&�XqԓC3$��֘R0�Ɔ5��)�P�$l��0�
�#P���-tVm�B���	��!�B`a� X%(&;aq�1�IH5�`V��o���!��
BC�a��Ґ�a�D� �"�Cc��F)��Y�8�m��@�����$I�b\&���7ᰱ��@l�revAb$��0����p�����K��4xЏ�A
c����1߱+���$�ߚ��.Zj%���Gz�MKg�����n>9�w�nr Y�1����l=�u�[�e�79��F�ay��T���:޸'�st"h��)v�s���QO.������_Z�)�.yY�g�S9�w��o$�sVs*�wC�ʷkMBt��vs�k/�G/�r��%����s<�t��὇��z�ϩ����_qa�'ߕ[�����T�\�-���SS D�-
��c8w_k�Ugi=)Z�|�֕<ў<�}�9�!�n�_zD�|�([�|a���R�rxV�{���P���Fy����r�����h��R�eޫ���ܤ3L�:����dGF�������S���I�}ݻ���#��)Y��~��J��Ϲ.���6_{��8����Z@-��تͮ�O�Q�a�{9[�Y��Y�E+�<YR�k3���Xj�JJ%����f���5Nv�[� R�]�EY��TR��y�`��!R�� 2$bF���S�(d@�xD����W	F�0�߼=�L�L0�N�^>|O�6�OO��\޹O=��=ֱ(*�eP��3��4Uv���uo��w
��s~�[Gr�}]�ԕ����ޛH��u�,�j���.�ۺ�E�W7�;ٵP�6ǝ�M�ej�7����9��B-;�=�����q��ݱ�{.��/Б�H\>8s��h�֥/&�l ��s�s	�o~y��f��F���"@�C+�Bk�,�f�!<�&g�.k\�hdY���a�.bJ^�C�9N�����&���e�(�(���wY���x���+yXw�wܥ�O/CE'���+"\���nm�2�\ ���=̾�s�y�ׅ)�뜓�<!��31������l/57�h[�ӕy߳wh����gy���Y��P���36�-m���n���W�}�י��70�;��+�
��Ŕ�ھ��q���E_3;���v���>��)^o:��~�����ǷƫK}�Wo�);#���֤��R]��_l�([#$
Ɖ�֧9䛗��p)��ƴ0!L����x��S	[�[�<�9�g��
z���`)|/�뇺��oW�0��
Mޜ�4h%5�#�$�ۜ�'�����0��%��e��w|�^j2P�+(A��H���ː5I�����%P�Adc�Hf��FdK����9�&�?���=7�O��L³�M}�oyÏ����pW�G;��_o�9wTR����>H�'���B����pڵʙ�pN�t�Uv��F5�}t�.���U�W���e���+p�]��/�Ue!�r���o|�?\IL�\HC�Kq��ni1>���!'e�&���Kٴv�}�����P|�����[��}(��*9F+����딫��N���xO7^r���d��.k�
���B(��h�n�?��w�b����A�]��Q��1!r�(S���L!BX��J J�
a
��B�
&$,*BXZĘ�$����bR���i���tu���H����=
�g���=ל�K捗�6��i���¦s~h�B��/9�'�y"L��p���Un���1�kxL�$��谷�W6�ο����N�/��ev�(�ܭ�U��<���"�5��/��g�/7��2̿�����Z���C�̮v��溯,kl��.om�0��g�9�9��r��K�@��fkl�Fs|����f�-�.�q,ļag�.�4a.�y��sB�
j���(\�0��+30V�K����|�怉 ��+��7}��K�/��!�5��a��ф�熝:�����k=����<+~��8�>�L�%��/!0\�cAl�yo��t���x{8{p��~��8��^xM�m1�,���Fw�䜼q��=ӄ��fn�ᙯ^L&��6Nm��{a��ύd�Cf�7h���bI�aOP�O�K/=e>����T�I�a�|=�����}���9fm��w�|�ʝ�s�s�.�*����u��,��h������V�`�^��+�>6��ӝ�S(�x_�Aw���H��^o3�����=�d0�.i{�8��.$��J�B	���˒�3��H���y͞湔�5�1������㥿|&�KdϒSWRa�'6߽�8��rH����.o�	9��B�/���o�D�e�Jx3F�u�g��Ю��X2�1&&��e�.�˞�ɫ�M{��π=֞�ݮ
r�]�W��뻺I��V�g��wt����e<��W*����g����kw���>@�ns�{����hߺ<��fOu�~��n�R������f��
�%0fh&��a$e"XR�
bb������0��ņ,
(¸�acV�*�$hD�
�
ˉ(D�-4���0�d�@��H!Gg���`i���M���"�h�-�����Z��,7�����7I�0�����Y�8f�6W���4U���xxH�M��B��R�"@(�"@#
�+(��Z�2�/����w�}��]���ss!����S���]�|�5]Q�n󊷆P@4+�/��wv��9�^&w�q4���=���̇ۓNyf޾k���[~�dg&���Ɵ�������rFj�s�/�?�7ܖHW�w�����j��_<�st�sҐf��h��aIJ9���zl%�l��.����/��#79�>b@����=�w��c��!���%ɓ܁�<���gѐ�4I��e���n#=��˲��B�^I����%Ԝ��MK�+-��-�	ak�����������~������g�y�|xY�ۈC��i�����^z���QӐ�d�>!��U�xV����V�*�iX/��n�gh�|�aK��M�}y�m�\�n��侒�HF��<��@�H{�z70��(U��ʟؾYήl�t���ma�p�c�[�s�L�y����s5̇��[4a6�߫��/a:J��$�2[��8y�	p�z����6���rϨ�]ޔd�÷Wy7Nv�*�*s��hK6�1�~�_y]�G����_j�N�U��!q�9Ϳ����U��76���_W�M��;Y[;�:�!R�����)�d�H��σ.�>r��s�}Er��i�N�8�NUo�+�]<��J|��eoA*�,�o��[|����_ic����v>�rr�P)�;�WiveM�櫤�)U�s:SN���_]Q���\U��)X����ˮ��]�}��+hǙ�]���vkl�6�dB�.h���}����g�&������[!Q�"�"Leۭ]B��G<��<�3\�a1"D��(J��+
a)���۟nK�m��� �nlQ�{�H��$av@�<n���o~����L���K�]l���܄�1)9��i]Gsw~�c�E����'+����n^���r��[Fu��|�B��uQX#e.]w���(]�+��/�\;�In����R�{��k��j����r�U]z����U������y��6ڹ���v��5)&��%��u��)K��WI*B��#�
!nڐ��߷�dlXᠮЅ�w=�9����F��~I�����+G��x��.�˞I<O'!ss��n��礦D�zp��]�2뚜�q�!
HǞ����R��F8��P�0aH�eʐ�.I��.�1��y�j�M��x�X���XS/�i���7�+���\|�)P����`s�w��9�s�j]i�	q�h�Ĕ�a4Ynjf�$���8l�e�e�ЗЁ5�O=��d���f�%0"B\(���Wܪ;]ۮ�>[׫3��J��e��al���')}�R����3��s�=���f��\��g]��+e���<�5��/�y�l�g��5u�.��s���j]i�4�F�a
��&�sL��YL'4K�.�+8Ng��������i�8�>,�[�(�m�"�E��Q�7A�7!�7>ܞϓ�s��J���)��Ӷl�4�B�F��`E(�<yp�B��aH�%G!#RǑ`�)�������~I�=pH�p�I�˳�"� �aP���|��z���<�%3W||7�D��<]�!!��i�����^{t�Cp���^�%�$��B�&���.]o�|�\�r�[�B��䞱.�bJ�Зi_/����-�RR�R>�O_}�K�	V/�n_�w1�g�����!��w��`{+i-�\���q��R$ą�%��o>�r�v���oٝu�*��}�Iv%˷����Ѭ�7���0�<��8�ƍ�|.�ݪ�������5o+�V��C8{��2�0e&aX{�j�����7�P�3{��5�3[�Ix˜6L��PvC��0/�D���Y�N����x�|��
���)�w>�+2�-0�P��ĕ��H\%r5 5,ġ�%ř��O$�ox�\�]3�����Z!q�+&32�ᄡ-e�����5�ݛ0��ۢnF����
���`XB�צ���}!��߹�&ؒ�b��
LU|:�y]_g+7~@����_m]m���F������:\�����\����7�ub]�e��$kR�=�.nBM�ZB�e�. FS.�ɚ�dHY�#�=��Ep�HQ��A�M7�!���9��lѲ$�O8�b��E�2��s�W���H���Q�|Ѹf��o�����ɹ��Ӈ�l,#)��<|8i��i�s��<%�G�cr!V G4F0�Ӱ���	P�"ͺ#P�\5�f�;�s'�<����>�p�Z*YQ���}
��U�73����u'�I���o�։�oL���<$�!\�IsIdhJ0���a� ���"�%H1 E�ԅD �:B\H]�t��ep�4�8oF�N$�{��*�����
���*����*�*�����j�*������L��6h˶M����9�a��I]���cG=ql�ђ��O*�M9��;F�s���b�HgTf}�#z^<��W���t���ʰ�V��$�:7�Nϻr�&ԵY{3*�mt�l�'m;�W6��S��Cۊh�W�,n^����Ԭ�n���}M��k�Bx�*��9�y�u2h�6�Z���Wl���ѵm(�q�5��"�1R�ښ�-�(�k����(j�l�
�U��GXwD��UZ�X\���k��Z��,�l+�;n��Lm���y�[k�N%x9U+�*�Tm*kq���������;:F�]�#ܵmpN���Cn�
���rl��_a����8��+��4q��G�ms�6�zyZ���p-@ձ$�W��b�jݪ�f�T��������}}]Jg���x*�5IaN��T��g��ɂ�vڞ��R�4�S;8��jꀢ��9��twn"8�&������<Ol��T��c5b�r�#M����$�W��z��(�tq��I�sH�5-UV��ID]BV� �Km�S�4U[q�e-X�q;,�UVS3E1��<UQ�േahwn�O�6����N�E��j��쵶�eӷ�Nވ�mWT��U/��m�a)MV$�PWm�R[,����e�E���`CB<��e��w;>:���*dS�u�\=/T �;�F�������׳�-�jk����YJ3m٫���~v!�y�\�e�:�pB�b�k��N�Sp! Ѥ*{�R��2��l�Tu��:��'mױn8^jY�\tpꭁ�fr�j�G*�&f5��E�Z�#�=�'.��FgFW�����vv2�&4���ף[<V[�n�z��t*�1��F7.!qv�M<��]U���{v�Y��ij��^��.H��,%?����g�z�T
�mV���֗cS�G�Y�UP]e��3$X���U+�Άҙ@�)�px �y�ۗ$H�.R�������UUV�דs�Pe����0�;��n����<ĝ����"8��ѧZ�>�ޤ�x6b����]�ҽ���a2�8���>y���1��.��0JI�6�`1U�j��{%6ꀍc 3�k��q��ԗ$1�U����i�9�D�=pVy��8���&j��k�4�ض(��S�����R�,i�\��8yS�f�+v��f�A�UƼ��=l��;a����ݴp}��9D��Y���j�e�*J�ҹ]�.1*��+%�tZ!�n�8lR�Z�<�qNg<��v��HU�
�����5uTy���+U�l�j��U[Uc�&�Q�;�V�ؖzi�SpBu͍�W����i*ؔ��l��7k�#tWA�U�m��mʇ@#T��#H�qFƪc��5�)hh�3]`��N0׌.���F�v��^٨Զ�P�NUX�-8{qP+ʭmU+߯��y_��.������̅-UT�N
Қ�]�r�APNL��U�81��yJ�_����BރƮ��.�
�/����r��
�j����gA\je]b�y�釳��p���w2��R�TR+ؓv⫺m�:F$x���>�ͧ\[kUUWU[�Ğv�ޝ��-�jh��@sj�����*�]nա�hW�V���'U�Rl*�mUǊ	��#T�!qU��@����ml%��@6����Tb��v��Ms�X��×�랛�v�N;k�8��P�q�����V�B �@ы)��rͺ�p�1�٧v�%f���T���:��{a�ֳ۳��C�����Dض!�����SL�ì�^2X�^�;tOt3Ϥ��E�B�B(��,-�jvӮ����)��k�|�S��@U[J�tjT䙸�5���U�քF��rMP�4��Mq��LU��o\�CksŷNP��M�
D��`�me���
�0[UQej���8#:�W*�U�P�תm��	�R�e�4�[Q�nҰl R��pUUch�P�R[�[UUJ�����<j�,�P���mTm*�U@=�cWO*��%y����a!@�K��QF�-6���I�g��W*�P��*UX����`�88^��������v�u����*�W�B[.��+MB��`b�j��l�J�q��䶊��g���L�]�:^.f�v�5�p+*�WUJ�W]%vD�J�$�=��� \]_U|`�u����^_U�<�Q̨�U���ͅ`yZ�ꯪ����f�R�UUUpV쭗����f���W�lp��S�&E�[�� +�P�UUlpUc
�UUR�C���mϊ�㸀���*��(Hw-����U��uN궪-����U%�T�@�1=���w/]�����c�=���<R`���� D���j�UU($��`Aڭ�����In�SUԤ�*�Uv�W�����l;1.�J�U\xU� �
UU� 86b�5/h���8x�u���Ɂj��ڠ�*�	��V��jR�N��Y�s-pg���cl�\�蠳�U�ʴ耪"k��;m	*���"�e�T(ejų��K*��Qj�T���ڪU[:��^Z�`*�U����^ڰmh��[�U]!5uUUme��UU�UUUUcqU�]U�l���UUN��X e���g�6��"����f��vj�Z����=P ��8m�+�2����+�
ꪪ�[j�*�@.[h�\�<a�EmWUUUl�����BU{+3�m��VW��$U�X�ڀ�5]U�U.!����mA��VU�@UUUUZ,[T��u]E�i�j��"�QjUUVm���T[*ۍ�ԅAT�U�U�����\�UUU�UT��`j���{7$���cyF��,Y�Xո��JR��n�������e���!X������x�uO ��UJ���Yv���*�� )W�
�ڪ�	VVN�����y���UO[��ѳRDҫj���Wf����
���W4�]�t��;r�UT�V�QT�Bj����*��j���UUUUUX���`�5UUUqM��v٪�����@A�R�Z���A��VʠR�2�V��UT�R�UUT����PUU]UUUR���C� ����j��Z��衺�5R�U�(�Y*�S�mJ�c�����>��r�c5T�vn�=��  �jU�:��䋓�K 9���U[���J�J�UUl��E�h�9��U���Ucs�Vm�2	�J7<N�k]���/���U���]���U�L�.��t���.��R�>�9�a�[�0{	j�.%���;k�h���J`e����T��j@���
^Z�����%�U_UUuT��U'�J�Skj���*�-�����UUݐ 6'P�fV)j��j���
���tTkL�:����ݸ^��J�V��˔�U��J�P��UV6HA{m[]Y��?����
��pNñMմ@K[�Z�;�Cd�9���u���V�$UUVQ�.�M�`:yZ�T�������tI������Ӷ�*�-���30�c=K��N:c�v�]W2���OFܱ��o@�.ʸ���k������LX������y���\i�lC��@���F�)v��0d�2���5$�V+W���_b6�,T6����Հ䗎���6�UEۧ�5*�*ҮK8��}+�mUUmUV�[��5V�X���$������|��� �L�6eq��\az�Œז����(�wsn1�[�P�.��U]@4��;,������qR��j�ݫ��Q�kVR�A�V����eY���ڣ��j��g�R�T�U���|}�ۍ�R��H5e��+������\�4�=����֠2��!`BlN��ȫ�m5UCb��x���8��ε$p�@v�FyZڪP�gEv� �V��
�TgY�`zj5��/R}��|ܥQU�R�Z���^We�%Q΃�� 4cMciTb.�)6J�i��4UN����Ms��Ί��YܨZ�;Y{g����`EUC%��.|u�s���jr��T��k��P�ګ��V���)�S�Nwn�'뎦�j�j���8
���[�����z��T�9j���Z��Sw�Y�Xxf�iI��������Z�9�X���۪�j�ۗ�P̹.g!��t���m����ӓW�1t��nv@��V���oN�A���Ɏ(V���R�a��mU�g�׀�ax�vn;>$Z1�s)ia�5nDG�=�W�Ft����I�W���=�I�����2g/km�K��떐ݭy�)�zg��m�m��gͺNC�I�%Ӑ�k�N^�q��P�E4X�y�٪������Ewk�R���ې��*\�	OKc@�$����X*�y�G����H�cz4l�q�K�]��v�ŵ�ʴ�xɴ���ݑ�@]�;Q��ͣ�b�u�T�AnnX݆��[ڒ۴{��i5:�öZ����Ћ1ҪoZ^܊��;��-���� ��@��8�z���V�W�v�Um���]��l[72 Um�^6k�����/�[J��[��UB*櫶�p#��!*�]��TU�h�[m��}��yZ��������U�[H�ڨ�䝐��R�RYVꪪ������������H���y�8�cC�js5mP5TUUR��1UPR��+�*[���6��tu[R�WUU]�*�UmUWU�٪��U����*N�UwqUT T�.�R9�꺕j�
��
���J���[6��N�,�����궀�S�]:쏭���gp�M��4\� ���k.��d��+�S�M�UUUUUUK��UUU�m@���.u��d�‧�Ѫ:�N�O!4I�j����8 U?����?p����E���
�m?���b`��
F�
��;�,H A�Q4`���������lpA|0Th�S��'�&�6��)�(H���B�H)��;���5O�� �t�m4 1"A�mD � � |��48
p'Ʋ "�O�W�@�~T�g�D�WA0�R,)���m��b$"�*pؿ �/ô�bOV��O�} `�@M�8? �S��_E�Ȣ|A@Ҩ)SEH/h+����T"xx�`�4<"���a���ZLЮ�=@��*@�� ���B(
x���g��TW�x*/��𫈇,�IHB@�c"�� ��$	$	! E��V@�I �$�	 BI$$��P���5E� <QP�8��a"��[KJ�I"D�E�H"Ȓ����X�B0I BUUҫ�G� � 	G�S�C����>�d	#%�����J�a@ځ� z� �b��<Ws�]"�U���UU
�P\Z�M��|@4�� *���`�B�P!(C���0�F@�V�s�Yos~N�Վ�&�6����r�<��;��hp���W��Q�
[nk��x�ۥ����#r3��ٹ8��ZpMpI��1�u�c Г��ez��6v�2;�)��V���¡�u�Z��K�H��;����1�j�+m�2����e��m�����-�e8��.à�M��vɊz��5c�1�r۔y�GvyM��<t��M���+���.��Q��w�^�G.���ӭjc��aS�ѹ�nv�-˗p=c������<Α;�F�^��1�gDQmnˇr0n����+��i��!q���g5��m]����S�5[��m�3�h���z��-�V�wZ��	Q0B�LgBj��Y."Q����Z�-a
\��[�E�47m�N�1�V�"��x����-�A��Am���87b�TO=����3�'l^m��������Ƙ�LxX�Lho��H�5�틨T�iZ8j��:���)�N�v(������v�:sL�][Z��]9����)-<�fi<6�:ykGF��a���e�z�
�3�ut4�mD��(T��)�l�E��01Z��P!���ʈ�Y��]��{f�=��1�ٍ"����`(bň��k]��`�B�
 U4�f8�-mUJD��q���H	�톬Oq��>�R�n��t5u.D�WB�8��]�cv[6a�aƻ�cu�)��:�^\���`Bd�C��%2Ll:僁��g��p�6�Pmb���]-���]p�1�⃩x�;v���rgl�qq�n����oӻW�\s�ج�z;a޺�n�E;Y[�����Nx�^̜ݠ=k���p�۱�\��'`���I��کL`F���(�<A�J��n"y4���$�x��ͥ��yR,�.��g��W[��ͩ�����w/v֣i�gL����3�l�VçH�Bu����`k#�[����j��]v�{[F��3g�	g�ċk�����Ê�E��51���V(�f�]��II���	��E���G�<�C�~<4��Ǐ|x���een�wmp�.ʻl�I���b ɮ3@Z�ySA� ͖��%]����JrM�I�<��.��ہ��m��@Y�Wcc8窥���c�t���.x	%�k��5�W��M�$�d�E�u�8m�f�����Y�WN�7a�S Tw����Oc��i�"M�3�s���V,�]�g6Dʉ{q��7n��qu�ک��C$�r]jLК^��&�fϾr��s�Od��9�l"�s�7l#ö���W���a��_�J�]���M�f͙X��`n�u��W������=B60wM���8�K�}�G�~�T���L��P�Z�i&�ZlV� ��w�un��9$��8�K�'n����ݶ�ZM��:�e��e`[%�\��WbbW+��ݫh�w�rI��ql��I{�[��T�J���I�����k5�XM� F�A��u����5�\�s��-ci�e�Xh\�<|��g��������ջ/ ��+ ��R�!�q��;;�{��]�9� �CIJI	$�"%�ڀ���/ ����8�%���J�*'L�e۶� ����&����uo�x���`���V��N���$ٕ�qvK�;#�`]�x�e$hc�t��n�.�xdq���/ �fVꯪy�W����Ī鰤��f1�k)���S��A��{6��6�3-�\*k���CE7Wm�������:���	6e`]�������n�+N�XWd�M�XWd��8�{꯹���%f��(��o{�|�[<�}�ny��"x����������1�����/ �ҡХ:*���I��:�%��ư��x�2�v���P�����ݻ�;#�`]��	6e`]��z��rT:�O���c.�4��+��N{\*D�Þm��ur���b�:�u���}���^&̬��^�k ݽ����N˴��&� �fV{���Hվ������]��f�
�鍖�cnـuvK�6^�x{���o�x�?������E�)����u�$���ٹ'�{�����H�X,R����g��nI�Y��֍k-Nݺv�n���x�`]������������9	P5�kn�4Z�Yu������@&�gڲ;����eݚ��bVЭ�;�Wd�e�w視�V�׀v�C�{����m�Wd�e�w�uvK�'u� �j)�(MЬB�˻w�l�����xy/H�`�޼f�)7B��������U}Ko}��=#�uvK�;/c�v����5i��n�	��uvK�;/c��l��S��|#�Ϸ��c�s��pvr��u�5֗��1���66++��gw(g^ț��y �эM�./7��m ����YI��t,�	jzJq����e���=�gx{t�e..��7�ɐˢwnxt�G"Ď%�۫��-�F.b4�`;���,��2�kef�� 6:q6���x�O,`�8:��§N�G�����	{m����3ݴs��㮘Y{fQ���o!��䳒I<��
�ҥ5bg�����n����|e��́]�!�W�E�F-L��������{��]�Se�u� ݉:�����[eۼ��;���W��=x�~0����{���v�P�\ŵ]�=��^7\0]����� �ԀvR����7eۼ/I�0�޼��;�:���9�����U��V�Wd���;�:���&�꯾��y�	�]1[ySk�.��M�#��WQ2�/�����5���H�p�ݚ�3۾���xWd�n�{����߿n��o�e@bg*����~��D���
X0���˚�r��d���U�0�4j8`:�I@e�i��������"���v^�x��C���I��n�	��`]����� ������X��2:��~���������7�<� �엀M�� �Ě �6�*n��]��;5ư��x�ظ���pߥ�n�Ys5kq������c�Qv�v.�.E��9���8��z���A�9.�����{�~�v���xf��ɩ �D���݊��ob�:�%���XWd��F�ĉm|[��m[0��xf�����X$"D BO^I̼�8`���ۥN�m���ٮ5�uvK�&���/ پ��K+��6�������|��:�%���X�F*��l)�wfZk���2c�y.�M��	��Æ^��j�F���sM�F�B�p��Ӏ{}���q���^ l�P�����M��f��/=�W�����}��&�݉4A4���m�n��q���^7\0��xV�Ѕ�v�Wj��uvK�&���/$�>�lSB#w�}�j�IϾ�I�w�݊��u� �W�W�{�_ �G���Xjh�V�� ��ys��rk''*�;m��k�m�$�Z�*�CCZ\ĎqG7' �����uư��X�p�9�)�m+�e��m���ٮ5�w�"�&�����>���FV�5��+x����	��uvK�;/c�v䦊����էv%m`u� �엀v^�xWd� ٤��I���N�m� �엀v^�xWd�n�`����⨪ѱ��g�$�h�D깺�M�=��դ�6�m�lZ��Ճn9:mq�g$�������`HH8۠\By,�݌/6��'Xvnsҧ+gv���x��9Y��Z]9c1��q�uڊ{k����m��&|�A9��lEr�\ggZf-�K�w[��������\���C�[F��LRY��q�j�Z��謲.J�eefaw����'$�xc�[�᭳�[���xt����vEOS`�տ>�}���8D���"���v��Yg�������^7\0��x�HЉ]��j��uvK�&���/ ���95*):EKk�	���&���/ ���:�%��6���Smvճ �엀vk�gK�r+ĒSw!�$�v2�V��ڷI�;�W�$�7#\�Iu\��$���s�%�fU�I.t�r�2�*�v��#w1*��q��u	(G.v���:���nz�7F�fGk�T�����M���w��-����3��(̶�߷�^r�d�e:E�tR��l�I%7r�k h 	o�]ٛ���u�u���|�w��ߏ�2���V*���KV̫Ē]�c�q$����I)���m�O��*�-ٛ�������%�/IM܇8�Z�ʼI$��DJ��V��I�|�Ij��I)���KT�W�$�7#\�Iz����	x>ߦݧ�\\m����1�K�.�7�g��x���6��6*b�K���]L���g�q$�GĒ]���q$�\��$�6��ĕ�>v�E�V�q$�G�W�wio�y�q$��y^$���s�}Uwkgi瑻1�r��� ���O} ���\ݼi����}�p�8�e��>�i'�r���]).�	�����px8mS���ř�y0�#	���Xf@5�f�F�Y�5*.��K	'��%���(�ᤀ�9�m�qcb},�.@�=-]�w������������nG���_B���3['��y�g���x�$.��绛	3��G|"<��'���t�������M��$�4:�0�'$^�֦��̫�.N������	-)8h�5�	�V��BG\I�%�2���-�TĘ��H�Ê<�!�S{��foDɬ	u9�k.Y��s�g�V����i?Ngh�/[�K�|�Y�6Mm+���&��y�!u����u,�h���&�wĤ�I���x�zlW���A<O<�T[�a	ĉ	$bE�� ��uE )n	����D�U_V�gNq$�lʼI%�L�ӥV�V��˻m�q$�\��$���s�%�~�o �䓛~���=����룘K��
�x�Jn�9Ēճ*�$�f�k�@?���� ����c��f��'
\kl6�m�<(�p�e�5k�*���LԦ��C�1�mfr��@?��o �~�5�$�Tp�}��r�%��I/]���h�i�� ?}�ϓ�@?���S���KT�W���IH�(�[C��N�\�IK�z�IN�C�I-Re^$�ٹ�IH�	�F|۱�i[�ĒS�b�KT�W�$�nF�ĕ�m=P�� 0XYU�0F@"�t�p J+5��nn�o~a�꡻,V�\�Ij�*�$������$��y^$���Ē���&����\@I;=K�(�n4	�q��I^3s���+<l3��	n�ca2�2��� ���5�$���^$��{8�Z�ʼI%٧��F3a��ʻ�@?m��x }��q$�lʼI%��w�$��:E�Nڢ�Z.��ĒS���KV̫Ē[�|�Iv7ĒJMR��ջm��Ijٕx�Kc��I.��X�Jwr�IK�R�4'e6�����I-�c�q$��o�<�I{fx�KV̫�m�a��g̢A����o����f�C�c�;h�2�GRM�44Tُ�
�V-V�{���lm�w'2��m]6K�r�����U��]s���ll��I�zF[���f���v2x�{FD�l�/e7m'a��˳�b��N
+'�}������z
٠UM�=�P\<']�ݲK����4�	��	��|����)�m��x��0W��2�^e�.]/��W�Fkd��g5sE�q�ql��<�f�2���v�n�N�q��==e+�E�������� }��<Jwr�Ij�*�$�Ǳ�8�JD�N�&�۱ۻ�ibI)��s�%�L�Ē[�|�Iln%�$��o�b�T�,���I-Re^$���;�Kcq,I%;�q$��X��];hM�lj�^$�ٹ�Ke�,I%;�q$�I�x }����%mu�\m�=����bI/�UU�{g<w�%��x�Kf�k�@�k�i�m�n�:�#C=���&,9�DM��m�t��N��j��SV]�	[$��܇8�Z�e^$�پ|��Ns�����< ;����j2M�ֵ9�m����߈��%T�s[&k\�Iv[�ĒS���=_U}�ݯm{�E4�!�����~��.��x�Jwr�Ijٕx�In�m���1��S�@?���� ����_}Z�e^$���;�IMH�&�ݧn�m^$��܇8�Z�e^$���;���}� ;9$���[�,2R1�X;�.1��9�؛�[��<�Gk�۵��e�7��+�1qY��\������� �|�Iu\��$���9Ē��Yy�.:�X�3x ~������|o Jwr�Ijٕx�Jn�ʺj�	���]���%�r+ĒS������Uʩ�dŭ�I,a����JH$�$qnA$�}��Q�/fU�I)�#�q$�k��2�6YwI�W�/���x�J)�Ē[���{�ߗ�����n�j&�-e��9Ēճ*�$��}9�Ԓۿz�߿y�����99���͌b7Pݯ3�.��sG<dleP+���8�r8䍑���rA��y|/���jn�������Ox�]��I%7r��m%�U�I%���J�Ɗ9O} ����m��3�8�QOe^$��܍s�����(u�)�S+�;x w�����＞P���8�K�9�m �h�M�˶��wfVٮ5�snE��������##ALDx>��7$�ߥ�؉��������n��	�2��̬�}�c��v��0t���&5Eu���=�鳛����l���]#�k�f��
����[��߿^߾�XwfVٮ5�wve:C����$m`veg�#d�V���`۝���n�Q��c�����y8f����/�X��V" ��RN���&��\k �^7fV��9$��|�_-�����(��4Qʰ?R��z��UW������@�O{?������x������Xl"�ŏ<%5��ެ-���4ȹ���tW�V{��m16�Yq#meE@,Md3���&0���]���-��1�s��nR��8zs���R�5��A��QȈ�܆��$�9ى`����h�+l���# �/;<�Qė��s��ʮ�=n4��;�׍�z�ɹT�<et�;���J�.wh4��w[*�	��Xs���VQ]�9$���%_.4�aK��z�&�\	p8�a�@Di�>Rs��K�.bN_?�Ú��)�����;�����8�I�8}����S޾WvQ(�/Y�h���d~3�I�~k ����^�~���/����բ�fnZ� ���L�\�{׀M����������"\5j�l��y����z�������0�`z�w�<���S�;-:i7I����� �l��w����Ix�"'���IRM��[4��v�M5Ȯ:��PS0���f�ֈ��T^�د/)&�m�Eӫn�$~0Mq��Ix�p�"��T�Wtդ�Z�Z��y���W~>�)�T�"H�I`z�FLF	B�,�!$4�-F�57�/fNw7�ܓϾ׌wfVz�H�
SŶ�ؕZ�v������M�=II=��o��X:�D�+���[n�ۼ-����Xw\k�K��z��%3�ݢ��j�V�wfV��L�\��������w���;t㥭���m��Б�������5�ؓ��ć0���|��C�Htն;�\v?5�ql��wob�}�'��	�z�4St]nիm��d��ԑ���{+ �uƳ�RF�{)�N�N��V������ٳsG��hTEd(�PB����r�y����{~�� ��۲Վ\��-�~��.��V���x�x�����^��I�wMX��[���;�=�ݹ�_ ���wve`v���v�Łܷ\������J�D{;M)���Ɗ�����nyv@[K�
�m�����ۑ`ݙ^�� �y� {R����wCB�v���&܋=U�F�����x����A�D��Q��Sj�۶�$�V�{������U]���������gk�d��UGfp?y����;�:��x��*�+kﾧWWW�ԘiP
|��;��}��svM:ƁSV��m�Ų^���W���g�ˠO{�V�{�*Lb�V�os�[aW�X��M6	��y����	�����4+�I'�|�c�W5*g{m�۽<�ݎ%�w�����T�� =�I4��s��x�u���y�Z{�w���^6�Y磌�*���+���m�ـw�<� ��/}��R^��,������wd4ek��U���'�G>�~��?w?~��y���nO�~U3��������G�n��+wj��6�,��W�W��������@��ߝ�RK��z5����@���p�rԡ�t��o�3�YĜ1��"FF F$"�$`Ȱb@��J�k�E!+�H�F�c#6!ȅ"j��I����"9IY� �������Ը���p-I��|�����Ot����Ҭ�N\�כI���!�B1B$�����|֎p!8�nP�p ����#)*A�`A�%�ܫ=�C������0vI�aKe!�1�q�#	O[���.h#���H����Fb���҃!Ĥ(��c�8�0/��f�0����
d��y$bI�{�q�0sE�VKI[X�Ki	5/$a�$a$� {�fy�<sG9v��l�vCf�6
k�T3y/�d�#@���I $�D��3��Pէ��!�1D���H"�0�����D�$�0��$d�BH��$B`�9�l[�)#$I";���C/Ĵ���HD��kZ=٠��Ֆ��6Yi�I��	��<��V;d���Uφ�-k�l����9خ��[u�xq�I�4c:��qD[�ܷ�x�&{QF�x�S<:�pf6�i�EV��&�1,+a��cv�:�EE�g��!͎�B�v�'0�ur&ͽw��%Z�v��	X3��=�J�E�\]�l�oe�O3oN]�衄Zn��Ƿkn�æ�gk(����g���v���^�����e}��ѓ��C:�n��s�7�|�����-������]���%�z͋�_<5���|av���G���sEg�r6�P]��NX��v9�#"J�)<��,tv��&���k���-Wn+�	:�s����zLu�<e9q׷''U�TOnL!ٙ<�D��nژ��uw-�L�L��cu&
*��8���qF�v�v�q��ۄ�c�c[@lh46؋nH��fM�n��&MA�pų7'(�a�8��Ӓ�.��kE�!���e��M����`�.`8KL�t2�kp�C�[g���k1O "&��t�q
�Dpb�"��Փ
�K�ƀ��Q���4l�gs��Uf�#WOE�r��^��9�< u��d]�t=��.Iݗ6!,0�d��Y�T�J ��;�0f�
=����f���/h�.m;S�=�#���&�i���c���S�	J���Hg�Ɏ�W,�t�4�� X�Z���
eI�Lm�-��녢V
Y[�&�[�03�����2aƖ ��ql�3�j�ݸ�����|�Ƌ�_3�� ���CY��u��� N��=�(/��spf�KG ��=�:��I�n���'b�広iVi1P�GԎ4�1��#�=�
n�|�������8�$=��	��cլ� ���)�4��$�sf��&Q��a�5��C1e[0��7r�v箉Z�O�W��2v�s�nҴ���Bm���͸6è��4������k�[0UG� ��PV�Oa-'MV�.�q��l�QVR㰀��ٶ@��dM��zڃ�7I[P)
힪V��R��[8<w�{���z�E��UTO��EN|+�
�*-=QP�T��kfHz�qy�3C�ֵ�a��n�{�;;��T��;M���ח��Od.���^`��r��*�:�N�Q�=t�����֧l�xp��pvx0�r�,��I�"�׶�xL�5�nH����:J�"�FYP����H���+�<t���흧4���k�gּtgs�ɜ����]��#�Sm鎣�)����k	r�Ԛ���?��6r�����!͋��I�5�.(�\OYxP�:=nG4f-M��v�y$�`�9Yb:�]��?~��`����$�U}�q��,my{ڤ�M�4ـv^�y���#W���=.y`��=��W�ǽx�7i
����^�� �{ϫ�W�U߽��0	���X$�M�����ݻ���UR��� ���ٮ5�ﾩ۽���{ߎ�EA�c6U�[~��꯷�<� ��z�	��vGg�X�2���ƴ�X�T��%�6)DY���@d(7S)���rO!�	�CiJ��e�p�~kԏ�o������Gԏ����o�a�@��2%�bw���m=���/!y>�ó��YQ�p�<�Ȗ%�b{��si�u4.���E�P�����Tم��
6"�0	�T4�H��bo�ٴ�Kı>����r%�bX����Wiȟ�
�L�b_ݷ��ڷ5�d%�f\�fӑ,K������r%�bX�}���9�ı=���ӑ,K����nӑ,Kľ|O�$�;���r��ӑ,KK��ݧ"X�%��~�uv��bX�'��{v��bX��dO��?M�"X�r��K���Zj.uf�W'���B�,O{�����KİE���nӑ,K���o�iȖ%�b}��۴�Ky�^O�קOfE�̫6v��rny7)�I��H�:	��솆{K�p������ݍy�%x�);aS�Oo!y�^O�{۴�Kı=����r%�bX�}���?
A<��,K�뿵�ND�,K�߿p�:�3M�jjˬ��r%�bX����m9ı,O��{v��bX�'�k��6��bX�'�k��NI9�!y�^C���K�l�v��bX�'�k��ND�,K����6��cP�( `�2%����ͧ"X�%�߾�fӑ,KĿO��t�f���kS3[ND�,���A2'߷��ͧ"X�%��o��r%�bX����m9İ",O~�t����������T��X�ꟑ�cĉ�}��E��u��v%�bX����iȖ%�b{�}�fӑ,K���}%�lk�%��+��p�����[�5D�M����xc���I$|@�<�k.k2fjm9ı,N���6��bX�'�w��r%�bX��_wY� �Kı=�۴�Kı/���]ZjۗY��ND�,K��m9ı,O{����r%�bX��{��r%�bX��_v�9ı,O�'f�SQXh�S>r{y�^B�~��]�r%�bX����m9� �,N���v��bX�'�w��r%�bX�vw��M9f�j�3Y�fӑ,K? �Pȟk��fӑ,K���w��r%�bX����iȖ%���Qd��x�	����fӑ,K�����nx9�S;�Oo!y�^N���iȖ%�a�*�w�]��,K�����Y��Kı=ϻ��r%�g!y;;����@.b�^)��,+���r��ޅ0!��|cԣ[\R�����������$�e��B�����r%�bX�����9ı,O;����r%�bX���w6 "X�%�ߵ�ݧ"X�%�~�߉ٌiI��O9=���/!y?���6��䀋�2%��w��iȖ%�b~�~�ND�,Kϵ�ݧ �X��/'���uج��ZQ]�'���,K����ӑ,K����nӑ, ���w�iȖ%�by�}�fӓ����/'��/�r������OjX��ߵ�nӑ,K���w�iȖ%�b{�}�fӑ,K K����ӑ,Kľ|O�L��B�[�Y��ND�,Kϵ�ݧ"X�%��`������i�Kı>���m9ı,N���v��bX�'�>o.Xt��)ejk����R[b��iG4���mf�]�{�O�lO�������r�%.8θ�og��v(��cb�
�nRO]ٗÚ�n��ռ�a֥�ηk2�in��c )U�s��F�1h%���$wK�g�=�,���%v6-FP����5�6��H��ֆ�� x{q^�w��w���1��6�+���<�h���dc�N��{��k��dڰ�W�
Y5r:Q7��`$�^1kQ�}����;���9�RV�hg%f�W'���B�,N�����r%�bX���w6��bX�'~�ݻ9ı,O>�{v��/!y��o{�%y�)\e�T�ږ%�b{�}��r%�bX��_v�9ı,O>�{v��bX�'��}��r�$/!y����֤u��楪�p�Kı;��۴�Kı<�]��r%���by߷�]�"X�%��}�w���B����t�ã6�lf��m9İ�<�]��r%�bX����WiȖ%�b{�}��r%�b-�ߵ�nӑ,KĿOo��.�֥֦kWiȖ%�b{�w�]�"X�%��H�}���m<�bX�'{�߮ӑ,K���w�iȖ%�b_=��0��^+p%�3�ϟ���n*v[�q��WR�r/<�@խ�1��� ����s-S-kWi�Kı>���m9ı,O��{v��bX�'�k���Kı<��:�r{y�^B�~ݠ|w"�f��V�Y��Kı>�]��r�EpWQ,K�k��ND�,K�{���9ı,OsﻛND��W"dKy��{�?�Q6ɲ�r{y�^B's��ٴ�Kı<���ӑ,P,K��{�ND�,K�w}�ND�-�/'��{{�laJ3
��9=����<���ӑ,K��;��ӑ,K�����"X�%��w�ͧ�����/'ݿwzJ�鉗+���r%�bX�g{��r%�bX�����Kı>�����Kı<����B��������Z�L�R��MeZvģn5e69�nyzc'���{b�5Ugf��I�@_#4�+���������,N����r%�bX�g{��r%�bX�w��Wj�Ȗ%�b}��siȖr���t�ãͳ��ȳ�Oo!xX�'���6��
X�%��~�uv��bX�'���6��bX�'~�xm9d�s��/!y���vcmCF9��Kı<���ӑ,K��;��ӑ,q4�@��(�*H�:WB��b"w���ӑ,K��;�siȖ%�by�B�w-�4I�]kV�f�v��bX"-��w�ͧ"X�%�߻�ND�,K��{�ND�,PV��o��ND�,K����u�e� ��Oo!y�^N����r%�bX"'���6��bX�'��}��r%�bX�g{��r%�b���>�� ���4���9^���M+��WD[��j�^Yb��]��k۫XV묚��h�r%�bX�g{��r%�bX�w��WiȖ%�b}��s` r%�bX�����Kı<���y2f5��*������������u<���ı,O����9ı,N����r%�bX�g{��r'�"D���w�{�ޒ��jgev<�����bw��~�ND�,K�}�ND�U�,O���m9ı,O{�����Ky�^O����3
��j����B%���߾��"X�%��w�ͧ"X�%��~�uv��bX�@iH�ɵS"w����9ı,K����p��ak�3�Oo!y�^O�{��r%�bX����WiȖ%�b}�w�iȖ%�bw��iȖ%�b~�=�C���K3�4�x��'7
���g���9��9�f�]r%I�����o��'�����3Y��%�bX�~��j�9ı,O����9ı,N��xl�Kı>�����Kı=ϡ~��sV�dA�y���/!y��^������,K�}�ND�,K��{�ND�,K�����9�r&D���z�#�]�h����B�������iȖ%�b}��siȖ*ؖ'��}��r%�bX�g{��r%�c�~���������0��Oo!y
 X�w]��r%�bX��_wY��Kı>�����Kı;����K9�^O�����k���nV�y���"X�'����m9ı, ���m9ı,N��xm9ı,O����9ı,LGD ��w��tja&���]�vG��:;J�]J�vubcq�����h����[����n�����}T���Gn��]�8�Ga�-=�Y��o#L�n�!�mK\�u�/p��)�y�Y�1�=�.s���E�I>Wm/Qv��V(UM]\��ю3շ@�I��{J�F���%iJWM����0x�&��a��z�8s�R����7�k	����S�w���2�?�]������hh�P]�����ۥn-vG�B��[���u��r�u��w���y��vr�9=���/!y=�{�6��bX�'{���r%�bX�w]��+Ȗ%�by�w�ͧ"X�!y?�w��#4�D�y���/!y,N����QlK����nӑ,K���u�ND�,K��{�ND��^C���p�n�m�Vy���/%�b}�w�iȖ%�by�w�ͧ"X��%��w�ͧ"X�%�߻�NF����>����m�a0��r{xX� !by߷�]�"X�%��w�ͧ"X�%�߻�ND�,��EA2'u����r%�bX��a~33.�6D����B����n���Oo!ı ^����r%�bX�g{��r%�bX�w��WiȖ%�b_>�˜":ɹ�<<�tID��7m��
t$Eg�]��We���k\�����z&��6��bX�'~�xm9ı,O{���9ı,O;����ND�,K���ͧ"X�%�}��RԚ̳Vk&�k4m9ı,O{���9��o���Ph䛥�V�)�T��CF �*���jVB��&f��Wl=`!�"X�&s�����Kı<��~ͧ"X�%�߻�N@DRı��{�~8~��2���O��O%<,O;�����Kı>ϻ��r%��"�Dȟ���6��bX�'ߵ���r%�bX�vw��tkR��f]kWiȖ%�b}�w���Kı;����Kı=�۴�K�@�=���ӑ,K����f��hպ�jɫ�fӑ,K���o�iȖ%�b�u�ݧ"X�%��u�u�ND�,K��{�ND�,K�k��]�F+ô�i�iݏnp�`���|�R���;;F�%�F��<������kT�5�5�kSiȖ%�b}�w�iȖ%�b{�}�fӑ,K��;���@9ı,N���6��bX�%�{�w-�0�.��h��]�"X�%��~�uv��bX�'���6��bX�'~�}�ND�,K�뽻ND� Ar&D��״���q��"S�Oo!y�D�~��6��bX�'~�}�ND��|HGĳwYI�rJfa!�lHzP�RPO�2Qb�$b�0�I��vI&�R,6Z��x�F�+R���7�}C̡��,��aaf��d̶an$�,�
:A�Z�Gjf���P&���o� 1���0a$�&s�b��H#��2RY5�kX��M��!�c�!%�2��I0H�`A�l�Wf���1�"E3zCa��
�X�j6RRBD�м<K=�9B��,�	�{���BD��t�1ٰ��u�\I���>� 24ll#!W~w6ncl�331̵� ѺĤL�3��0�Hy��h@�A�8 ��/G�>D�������_�� /��t ���A*z����(2%���>�ND�,K�~�uv��bX�%��g��+)����r{y�^s�r��}�ͧ"X�%��u�ݧ"X�%��~�uv��bX�'���6��bX�!��Ғ��;1��'���B����w]��r%�bX�����WiȖ%�b}��siȖ%�bw�w�iȖ%�/'v����(��h˭�#3k���rq�h�7n��%�b��(%˴�f��<�I8�g:gr������B������Χ�Ȗ%�b}��siȖ%�bw�w�a�D(�DȖ%������9�/!y;���oa�1�vv<���,K��{�ND�,K�k��ND�,K�뽻ND�,K�����9��y�^O���HͬctKQw��ı,K�k��ND�,K�뽻ND���"dOw�v��bX�'s��ٴ�Kı/��l�YsP�2ɚ�kWiȖ%��X�w]��r%�bX����WiȖ%�b}��siȖ%�S�H@BDYb�y�'~�:y���/!y�v��t0e�TE�m]�"X�%��~�uv��bX�"	�w�ͧ"X�%�ߵ�nӑ,K����nӑ,K���}���?CY��ds�=���n��}l6�+��0��fڷBa�G3�I�r�u �1`�`r�rT�,K�����r%�bX��_v�9ı,O����9ı,O{����'�����/!��_��F�e�.m9ı,N���v��bX�'��{v��bX�'��}��r%�bX�g{��r 6%�b{�Ĥ6u�e�\�us3WiȖ%�b}�w�iȖ%�b{߷�]�"X ؖ'���6��bX�'��ݻND�,K�Iٹܚ��Mf��Z�ֵv��bY���D����]�"X�%����ٴ�Kı=�۴�Kı=�۴�Kı;��s�5�:������Oo!y�^N��O9=�,K��ES�����<�bX�'�����9ı,O��}˴�Kı?�O��_Ǉ�f���j�œ�񒭡������-ͼVT�ƚ�t��'��Ȕ7�q�m�T�X޷I�.<Nt\��ȗ�ۍ�6(o���
�/}�H�4�4�n�v��cp�595��	S�l��n�@�8�q��`����m���r@��Ac�:c��N��2�d6��/<t��{Q�@�ъL�z�f���k�4Xa�)#�Mn^�H��0��'�u@�a.�|��6AJ��FiCK�v��3�ͻp�n@��l����>ysc6]	�Rf�v��bX�'��.ӑ,K��u�ݧ"X�%���o�v��bX�'{���9ı,K�{�2�\�&��fk3WiȖ%�bw��nӐı,O��}˴�Kı;�w�iȖ%�b{�w�i�X�%�{;�vܷZԙu���33WiȖ%�b}���]�"X�%��뽻ND�Fı=�۴�Kı;�w�iȖ%�b_!;ޙ�e�,�kY.�Yv��bX�'s��m9ı,O{���9ı,N�]��r%�`%���o�v��bX�%��g��h�ͅҫ�������������'"X�%���۴�Kı>���.ӑ,K��w�ͧ"X�%�߉����_EД�&�����0Peɮ9Ƥ��[.À\�Q�z�4�:���HD�Z��r%�bX��۴�Kı>���ݧ"X�%��뽻P�Kı=�۴�Kı<��M��ˬ��h��jkZ�ND�,KϾ�uv����<�T�D"�����ı?~��ӑ,K���w��r%�bX��۴�Kı;��s�4a����Y�˙��"X�%��u�ݧ"X�%��u�ݧ"X�bX�g{��r%�bX�}�s�ND�,K���˨je��
e�f�v��bY �'��t��H'׽�lI�9�f�pI ;���'�����/!����Y��γ5v��bX�'���6��bX�'���ͧ"X�%��u�ݧ"X�%�ߞ����^B�����������t�*rAm�l��Qel�f�sa��x�qpq��,���9Ns�1�P�j���y=<��S�b~�Nm9ı,O����9ı,N��xm�,K��;��ӑ,K9�~����`5�E��|�����b}�w�iȖ%�bw��iȖ%�b}��siȖ%�bw߻9����^C��Tss \�O9=���bX�����r%�bX�g{��r%��QlO�/�%���w��ND�,K�u���Kı=��RΙ0�e�ˬ˭ND�,K���6��bX�'���˴�Kı;�w�iȖ%�'��}�ND���Jy=�;x~ƨ���]Ws��y,K���}�v��bX�(w��nӑ,K���o�iȖ%�bw;��Ӈ��Jy)������*���r�j��:���⇐.��.���6h$�@kD3�[irs��TD���Oo!y�^N��M�"X�%��~�fӑ,K��}�����&D�,N����iȖ%�b{���Ma�f��aL���]�"X�%���fӑFı,N���m9ı,O}�{.ӑ,K����nӑ,K��۽�*L���.2��Oo!y�b}�w���Kı=�]�ND��,O{���9ı,O=��6��b�����z�M�6��`gy���/K�u�˴�Kı=�۴�Kı<����r%�`z�@�'M"�����6��bX�%쓽�a��dֵf�j]�"X�%��u�ݧ"X�%����}�ND�,K���ͧ"X�%���e�r%�bX�}&���������L9ב�g�E���U�pi�ӡ�T^U&R�ǒy����g*���]]�"X�%���fӑ,K��>�siȖ%�b{��v�	�L�bX�~���iȖ%�b}�IHo?s	�.M���r%�bX�g��m9ȁ2&D�>�_�K��Kı>��߮ӑ,K����iȟ�H��2%<�t?ׇ��Kb�����S�O%�����]�"X�%��u�ݧ"X�%���fӑ,K��>�siȖ%�/'�����9�U����B�����nӑ,K����iȖ%�b}�w���K��r'�o��v����/!y?�����GK1m�y��Kı<����r%�bX~V=�~ͧ�,K���~�.ӑ,K����nӑ,K�� ��A ؀X@Jj+"� v��	C���!��3e0\��#JxT�q�n��VQ� ùnK�ࣛ+r�[V8�o@��jŲ�yw������;nWz��+)�c��[���r�oF8�v���u��'l�v�/k�P�l̳���Ɓ�&v��Nu�6 ��n;&���9�Ȳq�w\-�&N���v��p�޲C::��S�Ь-!5�.�L E�O*�G�&�`�ˏ�#�s���4|��a�b˽K��%��cn5�9:�!$󗍭��n)a�t�ߤ�n<��VkMr�<��,K��?w�m9ı,O}�{.ӑ,K����nӑ,K����i��/!y�}}�n���C;��bX�'�뽗i�+bX�'~�{v��bX�'��}�ND�,K��{����I�^B�wK��nw��J��v��bX�'~�{v��bX�'��}�ND�,K��{�ND�,K�^��r{y�^B�߂��Gf����֮ӑ,KlO=�xm9ı,N���m9ı,O}�{.ӑ,K� �"~��~�ND�,K�Km���b3G�<����������ͧ"X�%��u�e�r%�bX��]��r%�bX�����r%�bX���|tFm,[�������#!*O�9B�l�H0�gl���g���������:�Z��k6��bX�'}�ݗiȖ%�bw�w�iȖ%�bw�ٰ���E�&D�,O��߳iȖ%�bt����F��(:�O9=���/!y;�ޛNCA(8��"X�'~�}�ND�,K��{�ND�,K���˴園�������\Ir!����<�Ȗ%�bw�w�iȖ%�bw>�siȖ?�!�2'�뿥�r%�bX����ǜ��B�����{�MT���\�3WiȖ%������ͧ"X�%�ߵ�e�r%�bX��]��r%�b!bw�w�iȖ%�b}�>���E�55d֥��m9ı,N���.ӑ,K������i�Kı?w_�]�"X�%��w�ͧ"X�%�|���)���g�Z�3�温�p�wm�rU����e�b1�$���p�R]G4ne�r%�bX�w���r%�bX��]��r%�bX�g{��r%�bX�}��O9=���/!y��;N�[�L.�Y���Kı=�۴�D,K��>�siȖ%�b}���ND�,K��}�N@ı,O}���y�e�a�5�Z�֮ӑ,K��>�siȖ%�b}���ND��?��@��	����) �"! �(ű�D�G�P6H���~���Kı?~�߮ӑ,�/!y;�_��qL�[�O9=��K�k�˴�Kı<���m9ı,N����9ı,O=�{v����/!y>������f�A�ZyÑ,K���}۴�KıQ���nӑ,K���w�iȖ%�b{�}�y���/!y�~�}�FQ�\A��z�����I:�1�7i#u@�[]�pb���f<��*��u��*�)��'�����>�]��r%�bX�{���9ı,O{��.ӑ,K��=����K�������)�̡r�<�����,O=��6���X��L�b{�]�.ӑ,K��>���r%�bX�}��6��B������;ҰڴuC7��bX�'}�ݗiȖ%�b{�}��r%��*&Dȟ����ND�,K�����Kı=��}ٔոk,�j�\ԻND�,[����ӑ,K���o�iȖ%�by�wٴ�K�� �����;�}�|�������;�ԻP����ND�,K�}�ͧ"X�%��H�>��?M��,K�����]�"X�%��}�siȖ%�b}�ߦ^���gh��0wl�v���!HawX��R챻�ښ�^Yb
59j��պ$p���Oo!y,K�뽻ND�,K���˴�Kı>����E�Kı;����r0���/'K����f�Z����Kı;��N@�,K��{�ND�,K�}�ͧ"X�%��{�ͧ"~Qr�D�:~���	�5���un�kZ�iȖ%�bw��~�ND�,K�}�ͧ"X�%��{�ͧ"X�%��u�e�r%�bX�w��Զf\�j��a����r%�bX����m9ı,O���m9ı,N���.ӑ,KlO����9ı,K�{ҙ35L���u�fj�9ı,O���m9ı,N���.ӑ,K����nӑ,K����nӑ,K��u�k�S�Mq�ۤ�2R&�����c[u(f�l�C{v<H��$`E�$!	�3�D�!	�˔a$3
�P�Ʉ��@1�&P�փ�bI�D�xR�,�BI��<y�g_<��}�-��-�%Uc�jBl�BB.����@!$�`A�HF#"�H1b������I3)k�Z��,��1H�ZrՒ,�ٰ�B����r�$����p-k�V�VV`Bws)�m�s���.��cA+�D��+r�X�C�cn����L/<al��-��,�(La�%ك�$���`ݻ-؞�����3:��.�{�V��-�l�%s@�$ˈ�%,���T جA���4��1�U�mw>7^gT��uXᇗs�L
8v�//	&GΪݽ����Z��+�<��u��v�����l#��*��6n���өu��GjKu�m��f3;�sc��[\���j� �j�.�E�fc�"�;�<<���2n|���a�b��`7J@eI��D�t��A#�5�J6�F�3WC���Wck� �\X��O4�o'��ek�F��3j�V�f��a68����S�����&{0pM�Ӗ�G'h�p��؅���4�U�v^�浒����-�ێ�ZNy2<9���!��ޢpuǻ]�&G�N�Y�!<����fL;<�js+��Rp�n���Lb1���n��L�Z0��<pp�Jbۓ��l�q��mq������v0F7k��
@ԶZ:���D��ښ���ViӍ��pT��rn��ev�V�ˀ��ۑۜ�q��'���q�q�v����3���{8uu�j��j�(d���,�
�\is(e)Tjʙ3�oY�gM��W9��\��bH�j��¬fj	0��
����ź4�k����X\�@m�hv\*Y3v�+�J�dշ:8���Wmȯdݓ$[k�VѤ��n�� s�XV+��a�I�pŚ���Ÿ�º:uKf�lɌ�$h\vz�eE�]#s�v�9��[�(�6�gv8�ˠ�jv�Γ�ӎ([���E�.KQ�]�т�Mog��l�8��^|�u�z:�šj��,X�]bѠx-a�@;��]�#Џ��<s[����[V�^��խ�fTϓ�,r����r����#��.�l��%��b@��V��0��F��()S�X� Bj6z;d�����ۓ�Cb���ɜ�A�[��j�^�X]e�ً�2+�A��azA�.�k�F�Q
���>P�4*x
l � p��W�P`� �LS�P�<�vbmm�b�0����ьК��8�2탗I�5�bH����K�ݡc�g����]�6W�#�r]�Dt��r�#;m/m��ӱf�Ye�gc�;f'H	��D�=���O�����6B�5��P���s36��G��Vސ����*I�i�m��Iy�g1�0fF�v^zڙ�R�,�r9�Zۭ�)�y}n�� �Μ۝�"]�������]�K�p�ѽ��S����ݐ��v�!'7X.��^$9ܱ�y%������>���[\�9=�bX�'�k��iȖ%�b}�w�iȖ%�bw�w�a�b��2%�bw�������^B����;�vX�q+���E�r%�bX�w]��r%�bX��]��r%�bX�w���r%�bX��]�v����dL�b_g֟��Yp�R�ֳ%֮ӑ,K���~�v��bX�'���6��bX�'~�z]�"X�%��u�ݧ"X�%���[HN��y&��uu���r%�`�'���6��bX�'~�z]�"X�%��u�ݧ"X��ߵ�ݧ"X�%��I���mX5��S�Oo!y�^N����9ı,O{���9ı,N����9ı,O��{v��bX�'��%���3Gn2˹���ѥ��.�qr�G���,�ܶ�f����E
�&����:b�9ı,N���m9ı,N����9ı,N����?�&D�,O�����r%�bX����ά�\�Y���f�v��bX�'~�ݻNCMuM Cq,K;���9ı,N����ND�,K��{v��bX�%��MLٜ�
�|��������^��r%�bX��]�v��`%���{�ND�,K�}�ͧ"X�%�zztJ5�k�y���/!y���z]�"X�%���{�ND�,K���ͧ"X�-��뽻ND�,Kܝ;���9*f�r{y�^B�z��^}\@���<pz��oo`���e��1�T�9��d�1�tZV�\��]��2@j�;i��wY)��a)�xf�`\� ���~��v�������IQG�,X�|Zvճ ��Y�ﾯ�=�<,����ob��$n�<�h�E��m� �Ix*u�}'�hAa����:��Ϯ�y���N��ɠ謨6�T���M��~���ߖ%Ȱ?/k��y�拥I��e��w�M�� �^��� ������v\�,�Cv;�X;j�V�q���4��mWX�$!�'h�;+gֹ����춒M���	.E�M���"�_������R�4ڦ顱ݵ�M���}I^�� ��y`\� �R2�����CVŀE$�mȰ�%�_��K� pԢQ�n���N�6��}_R�~��=���6����z���B��cV Y###���ԒB$�	��hX�%�dt$���VE� ��XHQ54[#��:[$�B)+h�%���F18��� ��^����~����L�.�e�k4�%Ȱ	��XRK�"�/ ��,��Mx��!⌸�0����ʳi\[�a�Y�7B\L�nbW���:�[�jKm`o`����E�^%Ȱ�"ʺ���)�v6ŀE$��RG��� ���X��,�9M%tտ�6_�7x[%�\�}Iz_�K ���x�%*�.�ݻ�I[N��\� ���"�^��^��^ z�K�0���鱱ݵ�rk�`I/ �d��>�>��I��#����e�5	����,jr�-����X̛ܺC�딞�;�d��L1L�dJY�v�,0�11��p�a;[��Gdo!�;�u� k"7�1!E��\�Pm6�5����,;�{'oC�zɶ��s����j璞]�A���j�)yy@e퐸����d
�:s;u�&��s/lR����f����Gs��f�Y-�m"q�Ӏ�9�c[�n�B�]�����燐���T^1�h屸ѧZ��޻d��ٕc�b٢� ���1s�cJ7e��-?���v��^�� �d�K�{靖;��� t�D��˿U��cM�-�����rk�`I/?y<����l~���a��S�(�Uw ��~�x&���$���r,��S.�.��"��z�N�KX�~��&܋ �IxԄʺ,���)�wi�X�"�=U����<��^;�Z�'woW02�˦X��g%��.�ӑM��%x����D](����	�7U�j��v\� �Ix�\�靖=��� w��.M\E�s�o{��K��y>ʮU]�z���X�#��U���Z��j�li�;w�zy���Ir, ��I/ ₒ�v:[��v���_��~�ߖ O߿<)%���X�V�cj�����m`�ﾯ_�����,K�`CQ ��㭌�Yq�����.@h0;����^4/��=-�f�1+,0�:��U���vٮ%�Ir/Uq=�<v���S�V���wi��6k�g���z�����"�^~��5ǝ]Z�&�՗e���_��l��P��EU#�>�$B�D#FI�(�Fj�ZE����!"FFI$D�b4X�+�>ʬ���y?z�M~K �SIZ����-���������z�	��X�s�z�������]�Z���<��.E�~�諾&y.%�,lp�$׾�X�c�Ց��Yn��e6�r�]̎[�(8�6?ic1�,X�،e\5j.-��=#�X��X����︃��y`P^�����m�n�ŀM�%Ȱ	��Y���W�a��/~M�Yt��m`�~���,f����=8��,�{]��қ*��w�y`�����ꪩUT}�P�@ �	dW�� Gҕ�N^�DL�[
���-�`5İ�W����t������w��yh�˜�5���,P�L�m!C���  ���*y��m��y��X�\0d� ��}\A=��=��CUt�i��� 7dx&�`��X�\3�W߾����]"��&�
�v����f����V�x�[j�:��M1�v��Է�<�6?���?}U��.�g�����(/��ݓ�}��N��<��&����y$��u�nI����rO��B�@`!�F)�"АU�"�EdT��E��V^��f���Z"�6ShS���f����8z�Xn][��7u�4Z�nշ��S'd�Q�"�c�h��H�zw��ݺM����wf�&f�)I��X�Š-f{����˶ h�q�k�۟b�ob�<�����s�]��4B�b�p]F��n�l#a;����q�rLbY^��2ة�K�ֺ�P�Δ�.MLR!����1|T),�]Cf���9Ü�5�e���a�M����r�w�7��%�1v��qe&��>F�X�X�9���5��~��|��k��fW靖&���7|�J�u��"��b��ɮ����z{+ �s� �\3��I�D�}vSE];���0z{+ ��ŀI{;�Q����6���Wv� ��� ��,w\0=Kޞ�`�����O��E��'nE�N���&���'ob�6�R~JLX9&�GD�0e��)�yC��u
.u��ݣ&K��؅�<��>��7=����I6��{+ ��+ ��� $�����J41;v���0	6ed�U|<LT�6�t&L�o˹$�w[�s�9���-=������I����� I���� �fV B�lvݗn�i�6�M� ����#�XQN���H�[o �����zg�%�,)���'���p�m,Z]��`ؕ���[z�W	�ַXw1�vv�Uɗ�����Ε�wC�pz?��X����=-��^�-���oY���n�-��v�,Mp�9#�&�`G��v�uh��X�ȰH�~�uC���eH�R�&�e�U���9���ӛ�"�#.���sCP'�6�%,��&�. $��w1�-��39�	fS�)9Vs0��)��.�������b�5@�V�J2-)e!iJZXolR���˘�f��Q�x9S ����w�81�w�ZJF�*l�#IU�	h��r�͋�2��5��&�b���Iʌ��&�Lt�r@�$�$BF��}�讦xj��KC-*��"���u�!lˡLGC
sI��D����H�/�&"4�D� �*��Q���+���T�������0�Ȱ���_]��+��ݳ�_R～0	��`��`5� 94�%:`���m�� ٮ��X�p�9#� rRZ�+q8��a�����������+�����!�q��-��bA�b)suXKWB�'�\����0���R;b�)���6�M�?W�W����ޏ��{��*iEi�J��m��8`5� ݽ� 6lx{F�jP�t��T1�f�\0�ط$����܁� ���
�[�y}�zpi�N�F9���cfp�ذfǀr\� ٳ+ �|�[��n�&��x��ݔ��\�{b�����R��j�'v0�;�n��;U�x7f� '���r,f̬v�, �v]�Eһt�t];�`�"�6l��7ob�$���_|��B��l�MSl���Oe`��`͏ ���i,n�Hm$�n�=�Ԥs� ;=�r\�ԶL�*/y6�۠�I�m`6G�r\� �����rO�iAO`
"B#������,��E4�Ad$ �YP0����cPVAG>o.Xh˔%%�˩	&[��1�(��	�����0Ťq�d-L#Lb����n�^�Y��K��6`���%���pu�)��,�ۡ�쎍o	�13���hGriX�6��e��X�CH�݅��ː}��\�	hR3��]p��2纹�ݨ��r
����8���\����ޥZ������L�lK4��1"�4�Q����.�ul�khc����{òN�����ɯDcfڲ��gc.K1*D�<Wm���U&`$�m`6I��C�Yf��ذ�`�e�������x�B��J�H��wm`5� ջ/ 7�<��X�a]:V�N���V� ٱ����X�~0	�Ɨ�+�H�M� l��K�`5� ջ/ ;�R�E���T��5m��"�$�V� ٱ���uSF�ՃO6Ҵqb������� ݂��76ޝ�o]"1��sY��wn�Sl���\0[����������;����j���*M�텶� ��f�p�Z�)"F�P�L�,@ ��O~澛�y�}���e`+T���iU�N�6� �0K�`$��5n��7�$�ʻ���[l���W˾~��7��V�v^�0�4��h,��2���;$��=_K���y��95� �t(tݵ�u�����M��[a����p<	�ǖ;G�-�]4���EZ*8�lt��+u�oob�5l��r^ŀvI��M�1����Њn����{�&V��� 9]��i�ݺt����9�{�ܓ߾�f傲�T'�g�^ }����蝍�Ŏ��o ݓ+ ��ŀ�<R���:�g��K*�d.Y�>�}��?O<��~��>�\��7d��=�����_��ݶ��g�P���h��P&��˹{N�v�������[�F��f�sp���������`d��5we�� s�N؛�6�f�{$�X��,Hឤ��/[V�]��[.�������X��r^ŀ�H�S�m*wN˱[�{{�ɕ�r\���L0�ܲ,#,$������Z�)���R��l���$,���!�����ٸ�����n���M�X;0Kذ�fV��� ��}�W�V���V��;�#��=b8}����9غ�S����ɳ�4ن0��05{m�������̬Wv^��/ �%:j�'V��e�X{�+ ջ/ �/ 佋7�"���v%t��05we�]��;��'ve`4R+i��I;am��6^�{�ٕ�j���7�$�VU�4؋��x��X�fV;{��/ ʿ����ȵ+Ug���155��Vb�`*;sŋh,���7J�<Ժ��v�����=��
\v슚��;Es�u��.����ayn�c�q�P��-���ۋ`tid��F� ��8�Vh���ѩ�c��nur�1Ph10&@����%B��;�/mmsO��-�zf�ю�3�,p�=�eq��.=���/��"��n]��l��Ck��k<�y-	�Mf�Ŷ�OJ9Vۮv�޴���vKr����&���R)b����tιo�}�{��;��N��/ �����Ҧ�����V� ���v8`ݙX6L�_:j�6�J�l�5we��� �ٕ�N� r���j�v�t� �w�꯾���g���e`��w�"�94d��`�lwM�V���+ ����;{ oiV������ݤu��v�޸�u(�N��k�:�6���h�1VU|j�S!r��~zp�L�v�X{&V i��[M6�\�ȹ8}�y9���I�O'd)~�n7fV7\0�D����ڶ�m�� ���Xz����=��s�h˖���m�[����X�p�&���'c� mJ��P$���n�	��w�� ��{&V���vB9��J��R�u�e��Ƶ�o.Gۣq`m��d]:���ꭢ�P�0�ذ	��rI��M� �wg�դݺ��Hw�N��L�n�`�KđɭTb�l��Ӷ6��L�w\0���}E����(D�# ��F�3N�Dڬ���f���vnI�=�)6��6ZCav�`z��I3��� �ݓ+ ��).���t�+�7l�;#��r,f̬w\0�Ӡi��hP�K�X>����LQ딶�͠�V��ڋ��p�ZV[l�m�%Ȱ	�2��p�'u� ��	���&G\�f���y9�O<e�$~0O8`�"�}��$��ί��%B�n�	���9.E�rk����' ���!0�h��,j� ����nɕ���U}E�E |B��$��b�>��|�M�'<���![j�WV�&�ɮvL�{��#�&��Rv�WV��V�t�A�S���v0Z"�У�B�W�J�Ś�̙�UM���m�;cl��{+ �� n�����`���M����av�`�p��<��,f̬*Ԥ�C����Wl�l���{��+ ����J��	ݷljۼ��X�X�`we��2�4��l���v�;�+ ��v�,��X��R7�\����k��]_'�8DԤ�^Iu������*B !!0*�+)Fā$�Fz�ڨ�@���)��ނ3�2"f�>��i�%�(�L8�Ja(f���!(�G�!�:}W�T�WB�����s/g;ަ��������8Nk�s3�˩sDۗ�pٮsD��2^sLyT+��ֆ���>��#�	�����
B�!20���׆d!@�v@�0��"��	$�d �y!d��������qxd��)�21M��F6�RC�I.��,�j��1����dda��1CDL^0!1$�N�Ȳs��������n7f�	�a��CFJe7�sd�L0-8$a�a&��g��N��=��yg9'*������ve���2�F����L��J�^F�3j{����H@�A�.�hP���$!�ؐjJJ���H�	F$ �#, ��h��	�ɽ��A��a9��a�0!��s����|��-y�o�%e�$B��w��?1vU�eҽj�L��+����`��Y��R.ډ�fQZ�l���RaHܛ�5	X�B����O;s�q�^V��f��w]���n����ap@]�:��M��a������!vi༂����0\���.�����v�*c�tt�t���cÞ;,v����ٳ����:����f:�R�6���p]�gG�p�,gWj�Rd��=Y�vZ9�����p�v��pr8M�W^5Φ�:NdvwY�0=��ñ�V+�1��X��;�:���g�8�����qL�j}�� i�'��qmڶ�%�sWcY"Kcs�ٝ���m�ݳ�#o#Fϛ@r�-�k���j���B��l�R�cpcʳg!�����vͧ�틂N���ic\�[\�(�شY��q���d9uӗ��9M��I{{l�KetZ�d���6m�x�GȒ�J��*�jr	���X@��Jy�n,�Ÿ0����\*ꀙp�.}�Wn�v�Uz+wGC�c��vS�L���ʷN�.wd�ADµtl�d�P�y� ��U]��y��Î���(.0��m�!=k��m����.#fH�[bpA	;���Uf��YƲ� ��Qf,�s���b�d8.�zr��%$R���ht-H`�e��K�+kĤQ�"wV���K�j�4&]g-MV�ړ�؅�����Y݌9vi�1;��99�-A˥�j\�I��ɇ�;aɜ��;v�\�p��D�׍�	֜�X�x��*5Q�ݬӞޗJ�c���.�}GX僂�֝ՎK�$a�T�=n�1i{H�n��qq�Xo0�k��^8}���-�u��Ĝ�5��ٴ��[���J656���SY88͵���u��
�p�)!4^`*X5cY	�T&��fP-�����3�@4�u�B��8��\��n��&��ͻ."�ѱN_a�a���n�@9k;�uA��"՚D��-^t�x3p��&�բ��2w0�vl�kSB�-Fش{�h��5f]f�N]Y���K��S��(�<M��?+����@Z('�)��@�0`A
QЧ���h⋉���}y�L�s�8�6���	�Z�׷$;�7)���9Ʊq��Ȕ�Ր���k�\&�I�-h Ȭ��4D\��wY�;R�Uu�#�i':�&�qk�v��{)m��8��.����j��Xy��)��⹲C�f!�]��wBm'[b����q�c��|��#�"�Q�-�����=3uݻ#�[=��Lp�^P�J1��I'$$�9k�b�����zB�M���v�S^����x7��`꣨�h�%E��U�ZQ��p�ק �b�9.E���� ��e`�{(��j�ݗJ�ـM���X�e`���S� VʵWV�v��8`$��7��j�^����:t;n��f�L�{��#�T�ŀsK�t��6���u�ou� �W�Oy����&V����Cv5��l�\:�ױ���@q��6�n��>�Z�])�̧alͿ@{� 佋 �+��G� �i:��[u��\��f��>���Q|�����əX7\0	�"�9�4b��,V�ղ���$�+ ��H�r\� 6�#���m�hV�V�R�܆$p�9.E�I&V�&V�Wm��T6�H�r\� �L�w\0	K�Ww(�ݪvYKB�狣d-����*�k�r��8ݮ��ci�b g�n��![�]]Z�X$p�6I��n뇫ﾮ �����5^av�`���`$��7u� 7�<�8`zi��E�5��8�|���}��;���D#" ��Q��Q���=��XTj��C�wj�vƛX����)���;���ٳ+ ݽ� �MJ�V	e	�@��x%Ȱ�e`��`fǀj[-ݺ�}[�շV�O\:�M�]n�e�Z��n�����v*0m�|!�W�Y�nnGf���y0�ذ{���"�	]�:m4��ĕ���7ob�}_U}�A6y���� �ٕ��H݊aAi��h�E��wc�'nE�����{+ �����I�§V�+o ��6L��}�{�ܜ8�ot($��}��=�٩p-[��c�m� �ɕ�M�� 7v<v8`�)d���V'WB�zS��r�&�\�o��D�Pղ�!�C[�1��.ڳ1%q���?w��{�\v8`�2�Tj���vR%v�v� ��y��=���;��w\3�W~��i��+�t:�@ěx��ɮ��X���m1K�v;M[j���]�x��x����s� 6�t�c�&�X�0���{����`��?�_J��}_���[�f(�k��̇jt�`�M��:2s��@�Ϟ�)p��ru�XeG5P��1�D�ي2�/]����d�$�62YP�Rh/�i���g�^�&��kjD�+��m�O5�x� vq��w�RYm\e��D����gbY��;Y ���U�Ɨ��Bw�����m.%���f�[ul
�r���c�-���s͸8t�b�72����sE��m�dr]I��S9��HƵ6K��w���� �zpMp�'ob�wT�$����:�J�w\3R;�2�	�p��c�9��pm]�SmX�l�9�2�	�p�ݏ ���]Iwn�t�m��n�	�p�ݏ ���L�U��t��줮�nـݏ ���fV6�,�W�������$;u��W^-j΅lX�5����pa�������%�:D���T��0����,�fV;{>� 6�<��Z�,m�95�r��߻��I&�<<<��a"�������*��X�v^ N��	�ذ�"���:HjՊ�`we�7c�'ob�9�2�	ئ�C-�-Ҵ���c�'u� �ٕ�N�ŀ��-��Ӧ�]��N܋ �ٕ�M���}�^ }>�\m�Tn,ř�\]u�s��<nP}`�v��/2�ts5.�zڒ�cMX�6ـrI��M� ��x}�Ӏ{�{�p዗ll��M� ��x�p�96e`�M������v�����	�Ⴏ:` (�!�)BB���C�{���w�k�'<��I��eҤ1&�ɮ&̬{����hk�J�2�ݰ�Z�`�X��C�uwe���`V���t�+�$Yl0��S,��^s+�: ܭ�93q[hl��:�r7�/k�����XWv^�{�ɕ�wjL[Ƶ3*��o�ws�i�wDvL���s�~C�5I��x6�,��+ ���ݗ�se2�V�j����m���+ ���ݗ��T�����)W���,�]Ijݖ��v��V�`�p�:���KذM�X�^�.��R��M�I��К��U���:Xp(g��NîLl�!����I��Rn؝��g��{ɳ+�U�q۞Xt�P�۲�4�!�6�KذM�X��, ��x45�\e킶7m`�2���X���Kذ�����ت��V���7��`���KذvL��R`�Bl��V���{�{��+ ��iZE�*ZV]�� �eje(1���V3\�����.1��cOM=j� �Ǳ���!��[��w7�NJ3���I�	�m��c\��>�*9�m��Y����-�hG�v�pg����㵠S[�d��<A$e�,;�x��BӰ�Wnj�{M>z�'�w3�"�ы��dC�B	:y��׶�Z!�[��9=C��M)��8�їR����缓����2�"6�7hCTϠ�\IEI�^hx)�pJ\eY�":E[*ltEۼ��y`�e`�������W���;������e���2��p�:���r\�=�~�*]t]�r�ߺ�8�Ix{���`{�XTn�N�:���n؝� �^ɮ�X�\0i�j2�cEJ��ɮ͙X�\0Se��[H�Z�+6�!���iq� �Tq����K�B�k�ٙ����2�:�r5N�~�&��T�x%�X46g¥N�4\�����=��}7���@�A �M��PY'�Ͼ��oob�;6eg�����`촄؋t�l�"���9/b�96e`���`}v�M�t��x���|��w�~0�p�5we�]�\)����e��Mp�7ob�5we��"���C�ПM�"��m`�V���v�5��6�,��v��nݱHvi.y�1��&�;�E�g ����/ �ɮTn��'Lj���k �ݗ�r\� ��v�,�4@�X�Bi&� �$p����>��R6���>����!�<%4���t`D"@�E0� F�I���Y�i݁9RQ�B���dp���0!BȗD$�0�r�vkSZ�,X��t�ڤ6���I!J&%�!���$$Yhn�!m$!�y
O#��835n��s��`�! ��O8I0&ap ��!	 @�V�����[*%ZA��*�"@! D��&��&A��V�+��P,0n�C�8am#
JXXTA6n�XM�Bii!�]�ڭń1���4�
H�B�HM!b�!##1�	�Wbf.�@>��\�[B%.@ (��i4 |��|Tp���ߨ��C�@���4��Tߞg�]�<�{�nI�$��X+��1��l�9#���V��\0��L��v�V�]�l�7��jݗ�r^ŀrGdj5z��p�Z7��q�f����������R���s�(����uF�yv�H�ElV���,�8z��� �� �O�lV:�H�.����g���#���Is� 7v<���7e5V���[k ���X����"�;ތ��2ܮ���{�Ӏ{��ܓ�g�]ɧ�*�2X)T
F  �VN�M&�o>�~0T{�F�+5I��;f wv<��\�����v�EAux��k +�_e�獹�z-�&�=���؋d���M�mj5��I�3(�5�LZ� ���͎�`wc�9��h�Ӱ�:�m&��3���${c�'� �=9��'��};�r`զR+v�f�� wv<=_}I{c�vy��;+fR����'j�6`wc�'u� ��w\0�[�*�V�.��'u� ��n�`wc� ���(�A3�o�fMCP֡�%њ;.ɗ���DP�غ���(!��&�-(��Xu�kf9m��k8N6��`�õ�Qr�����l�6�Ζ�5�p��uk�n���v^^S/l������}���9��nuB�.s��W��q��^�Bظ��QgLne�9'�8�<qWcŇ�<�0hv�w'ZJ�F��YSqSr�(ލ�j��R��ĺ���;CV�%�������be�/,\n��m�e�x2�Z�$�ۗu�g��{!�y_�2nlݥ�k�vՍ��h��`��jݗ�r\� ���n��-�0�p�5we��"�95� �7Twe۫��tյ�j���9.E�rk����+R�S�n�E�����˾s� ��`�p�5n��9��h�Ӻ:�cv��0�`�e���`i.�t�M�mS��i�nθ��ԅ��lGM�]ӻkQ�P{p���eۦ&���f���v^�{����;<�`*{)|�v�պnnI��߳~��@��K��Ϲw$�Ϝ0�`wbK�*�V���x%�X68`�p�:�e�[>�:c�mX�-��諭����M��ջ/ 佋 ���m	��6�-�0�`]�x%�X;0	��Xnŵ.���PF�fC�u�nM��=wm�v�s<R9k��h�[T�e�Q�GV���/ �����\0�>�{M����������I<��Nl~0��yﾯ���������N���f��� ��� D�	B2��0�@�a�$"�`����n����x�e�Wl��_}Jl��=x&�`��wkfR���S�n�M�ջ/ �68`�e���;H/�V[�K�r�����koZOe�H�7p�����F���Db��IpE��l��޽8��z`�e�]�x��)�c�6[�e��Mp�UW�|���-����������u���i��s|��������K�`��Dj؝��Ս�m�����^�^�_��M��rH���-`�0L�6Ut��^���s�{l�WWcut����"�95� ջ/ �ݗ�jIlN��
Wn�u����C�:!x�4Z����E;���5�E���⋦i:WV�0Mp�5n��5we��"�7���)��m[�ݻVـjݗ�ݏ �ɮv��|��CJ��� ��x%Ȱ��UUIw���"�׀�(E;47e���r\� �c��v^����-��M�x��n�N�����X;0}_K�����r\� �U_K����p嘎T�&�6��{n�Q%�W^��K��&F�ƞή{��뷛>W�6��)R�(gcf������)׎D��9�W'�<�-ʀ<�P��s��^�`�jK]Q^3d4X��V��u/7��YMf�(��ͤ��G&�ݶF�դ�L]��r�V��h�N�I�����)�7q��W��+�na���n�B�@6$v�d�°����Y9�g'ne<�fڋ��~}��g��f-�(d.�7;2u݉�:���LV`Ջ2�����
{m���� w��r/�}����Aݿy`�)�!��*����~��I���L�~��&�ŀoJԇW�ƾ�wI�x�Ȱv�X�ذ���t6�4O��m�J�k �nE�E�/ ;ݏ �{����5m�v�[���0	ۑ`{��ob�9���K>:ֹ��L	-غQ������b��� �����J�fj��u&���4Cv� w�6�,���Ȱ���C�M$�,`��m�Y+k�U:��;r,��/=�U}�F�����de�-�����;��o ����"���7`�;m5t�m�;f;�v^v^���wfx�""��N۵e�Mۤ�v^v^��6�,�U_w\B��;�3�Ȯ[Oin���nb7fh4\b5èӇ�d�äIm4p�ƳG&������ �ob�&�������ΆҦ��n��Rwi��9�с����8���"엀N������ݧm]�`o~��r��ٹ��F(0�@�D ����UUV}MZܗ�w��vh��J�eۤ[k ����"엀s��꯫�^�y`�z�!�c.�%v�n��%�����\�������{ї
�L�4֋u4F��������'K�:3d9��T��f��Q��]�p�&�x;{6�,��� ��^�S��M;�v�[V%m`ob�9�ذ�%���Y꯾��H��W�M4��M5ui��wny`vK�9�ذ	��`ߴT剃�u`�ڶ�?�{����'��ݻ�}�{�ܟ�
D�������˹'�I�X[�]I��N۶�w\0	/b�9�ذ��p�Ie�]ҳV�FW8q*��g�m��r�I�H��T����٬�:�x[�5��$��Kذv�,)���}�߫�<��x��@�����V6�ջ/ �l��0	/b�͔�M[�+t��]��"�/ ��=��{�<�Rz�m�U��:��n�vۼ�0	��`[���%�e:���N�J�jĭ�m�XWv^d���h��)S�R�0A��Ն�C��f���:Q�/�B�b@�M'>��M�$X�0 �,T$$R!`P�B#HH2�rd`�+	#MV�.�f�e!Iv���3{�	B[JJF-e��Zm5	����)ˎ���h5�4Vb�j
f��D��` @��aF$�̥��el�{�$c �	H�B$�$H1�FHB�� Hn�y�7�I���)l������||���s�<��߯��ׄ�&�3�!bĄ0��
H@�D�`AH�P�R1�d! d�I!!�J�$���݅�km���A��5���m�֡�R�@`@��3	eIF�	i�cHHߴ3{�w�B��Fkr��� ��aZ$ H@5��L�����R �;	H@bB�0��!��`HB1�BH9K&���T����$H�$bɢVYXP�$H�aBo�GpW8o�2k������|��^���Vޖ�Ě��۴��9��H�������s�4�Ѻnڋ&6� /#�������rRә힋�5�s��ۇ����q��3���7=B�c�Wv�tqcO�vsZg'[�t��V�6��6��c���S$ e��Q�e] e��Obn��<�'k�0�d�
W��V������O�^��wR�ǆwS� ������\m���#ثcl��K�riϭɓ�n$zS����]
`4�r�ph���%���[+���%;lk=e��T\����
�!gW)]Srm�7
mL��ԁ#MCH��7m��]�5��^\�M�kl�l�DXb4l��ۀ�&i��R��q������8򼶍!�3�0�M�b��p�,mvL�
�{�^mJ���y@�X[ �F���Cb1��h:TŘ����j}�`S����
T����?}����c�#|�ퟴ
#�2q��{b�Vvg��[��Z,U)�Lǎ��s͡��9��i�KB*5n�4l�]=�;Y�=��s�v�+MWb���H��Q3m3&9�m:�9㮺�(����1vp�B��bG�)�Om�Q;���0RЙpV^�a�.���Za�ԅ+)q;i�ۘ˵D��g���@@-a�����Xr͟ �L`Rn@�!��nJP���`ݹ�ؠ��Pލ�-�أj�g�rQF��3TU��ܝ�a����zr�f�ѩ�R]�gØ�ktg��\#�Ģ��u�mO�V�b����%�%�d�(��d:��x�;c�E�,=�^ֳc���U��`�x�]Mc�k`ۧ>[ql�+Ϣ�}��v����l��j�vݺV��#jr+a��sɮ}p��>>���jóXuIy�FX�0����W�70���R�[;E%�n�(N�7!�.<a{u�D���L�ոM�b�m:x�Ƴӵ�a�3��6�/U���kl&���AK�����ϓ�Vּ�S�y�\��svcah�#<��L���ԙ��: :M&����(�DTڏȃ_��W�x+���!��ɒ۬����6+t���y��|N��S�l�S�F���Ǻ�$�n�D�k�P�&�5�Z��Z�T  :� ��]^��׎,�'ugU�z�v�ל\�l�0;���v�����Id����b��:�wc,�6`�s��&,����䷒�!����=;�.�M�9��C�6=`���Z�13�ܓ�ĝ[<W羾x�WK���\ʅg9rm����An&,-B�M�sH��VQ���l�'��{�'������;�Zm@<�O׀E�/ �c�6�,�Z!�ct:WV���d����ذ���UUW���́�L_���E�Rwi��6~�m�XWv^d�{[/(�7V�m]�`ob�:�e�vK��˳�� ��{�Bܤ���·�{~���v���͎�ذKZ�*V�lE'M�}��N:q�����[�,k$��rs�F�kv.2̷��i���4�;�v�����^�m�XV��r�M���M�z��9���o��?�5 <Cb�Th�?�3�k�ܓ���srO��}���^��γdL�k�Sf�m��=�Zun��"엀sc��R�������[rz�-�� ���}_|�&x�;*	�����`�	��"엀snE�M��v^�+B�K��m���+P���	I����V��t��J���h(U����7�#s)O�9�"�&�ջ/�UUWyo�x�;�NytU�[�� ��=9��'�y%RF�=x��׀sc�z�H��{*�J�)�i۫�ـj�׀E�/	��Uz�(� H*2����У�/������ /��Lv4]]ۼ-�x68`�"�:�e�SbM鱂n���lp�=U/}����v^ŀ��j�M:��E+�l1�.�D�nUN5�����[�o,�lat:盿|��l�Λ51�O�;~��p߾��;/b�9�� �i����ww`�� wv<��,�r,Wd�zh�Q�YhmЮ�m���`ۑaꤢ�z�d��9��4�w_0�m�k�UR�~��"�z����g�'�pA����s�.�|{~�n�h�Ӵ�m��"엀~['� �׀qI��;�{xۊ�)���M�%���A%/E��ӎ���!l��xequ����ks�[v� 7v<-�x���%�l�ñ�հv]��E�/?}U�URGW���<�޼ ����$��V�v���Cjۼ�{׀E�/�}U��'��'� ���m�wm2���d�-���e�l��ujZA}v����݃�x����^�=|�{׀E�/ ������&�� �J31�)tq)�C�T�۰�����a5nҼ/g��-/v� ��n۰���n�ͩ�@�
�+ S3[tC�V���8�v�`{f1Cl�w�L�ķE��[H�V84?���wԩ=�q#j�8e��Bq��l�[b�5l%���"fR�
ns/Evǳ�@&1�������|���]cmZ�0�Wl0L_���Qe2De��,&eə�e�t�楖�=>���3]���phc��'6dr�y�w<>��X�52����`+巧}��9�"�"엀ݏ 暄�B����[�v� ���}��}��?)�����<-�y����Hݨ�e"�v�ݻ����}���ǀE�/ ��{*e�J��݉���w�ݏ �v^�0=_U}K׾��O{��[���ݗm�we��� ��/ 7w� ���y]���M�@@�pr�����K;t�z�����C�l��`d�ٺ
�+h��w�;<�`we�[�����	 ���vշlAv� ��/����~�F��x]�x�x�KH/��u`���ۼ��/ ��/���R]����׀oMN�F�+��4;w�Eݗ�s�� ��/ ����9��4��Q0�wi��9��{���׳�| �<����	4���v ��Y�'f��7f��Ng��r7��;6�s��[�-�/����-��e8o�*����we����?�֒E�v[[v�����we��� �����H��۲�$����'/�}��ڕ%T�J1�Ĉ��� pPM��F N���DZ���M�۶��$�w\� 7v</k�X����un�m[V�n�	�r� ���	�ذ)%��/K��iLWT�����:��pq�	q\Prj�>l9C���󖻈�"�j%�Kbݫ� }��x}��qI/ ��(�;�S�R�0��cv5m�u�=IRz�-���{���P�
��>��v�f�6^d���ǀM�{QC)]�����m�����z�ޫ�	�� ��'�@F Aa#,�D���y��绀}��в��.�l�n� 7�7\0.�x]�� ��}��0!��P)g`��K^j����v9S0���]�	'SqQ5�z��.��'u� �^��ݏ 96 �j��ڴ۶`��X[�� ����'c�{睊#����:�I�vݴ����g����w\0v�,V��I�I�Z�j�����/ ������_UR���^���%�AwC4Л�w\0v�X]�W�uwe����A�����-W�V�`
�,bů0Vh�x۷�qrQ':��Y=��k[j�۵�`w��)�A�#�y7N�F����(�nҜ񳃌z�Ų�L���ېm��܍�/���=�w����8LPe3��`q�iC���Yk]v�Tp�Ѩ)O65*7�z�qҺ�"���.<m�pPY*�x��P�v��ܘ��Gl��K8�^b6qՀ��v=!Ui�w�''%����|-=�B:T�zm�vxc:-�V����������ㆳ��a�R�P�G����o�~<��we^�ݗ�N��֨e!ZN��+v'm`we^��/ �����Z�/�;�[)]۫�:�%���w�"�&�`wv���Ֆ�t����� �nE�M�(�:�%��H-�T;E��0��,n�F��/ ���ԧ�t��D�74m�L'�Z1�f����pA���m��/b�&e�V`�����PAO�o~ݡ�����ooF9}Հuy-"WI�Zf�[u�&䜾}�o�"�A6����U��*��$�%�X����R�VZV�	��$���� ��R�8�%��m;������N�l�9�ذ�ʼ��/ �\0��C)%n�Z�k �l��8���	5� �ob�m*��wv�M��H]���UF��	k帻���SVz4<�������m�WZX�6V�n�}���vk���ŀE6U�rl�E��wWv� �\0v�,)�� ����	�P.�t�(v�m�`��X��~3s�&} \0�\�u��5��'�ȵjV@'!�`�@#�� H23~)��C29~�FM@���a	�)�Ч ��t:`�)��q>�_�}�:�!.�S����$����)+.�3�p����Ú9r�H���������������|�
�%��̺�z�ٓn���*i"��wH����Mu���d�r}%���)�ӽ����73�0d#"�!�d�cJK	tI��S��zз���c�'�᯶�2�d@�BB! �BU$	��Z�6K����5���[��-H�H�BB$����0��>!��3�	w�����v�`]����O"Jy�����Y.��|���d�8G�"yo�nk�d4��
d���BM1�"0���BA���g��7	yL ��k�<�0��M�@��! � �H$@�	#f����#�����OZUFI�Ĉ�O
&L ��h3'��b��"'���h@4/Z /��׊(�R�L~4�늦 ������0"C��U�^�D �z��Ͼ��9���nI��G�۴�n�m&�k �vU�]��	����ﾥ��JJ���������8�%��� �ob�"ݕ���}��i��siw	��P7�oM��.
T+[��{<�u�]�#��!���^5:ɜ�	��'c���ŀE�*���qV�׀wBS�H�^��'cl�;�ذ�e^��/ ���#v����E��vi�m��?Q�qvK�$���{����}��������Xp.�x��`��X�Ԫ�����ꔏ}"`:��4`��Gj������ '���_�ճl��� �ob�$�(�8�%���^�{�Z��2V�B�txd�X�1H��L�e��!e�iMM�\�lu�n�&f��wny`k�`]�~�����=�~2�߻u˜ʡQO-�~��/��>��#�g� ����9�ذZ-Q+�t�J�-$�рqwe��� �ob�&�`���"&�J�ʷhM�;0v�,m쥀qwe��m;�����?���`�`#�`]�x�p�*�����ң�(����h�c%0�;��E��Z�U��{rY���^��p!���q�rtkXݴ[�C��=�s��[�J� �0[f���r�[;sٓ:�q#�'#�vwl�;��sq����#>�r�����6 nn��	���� Ψ���Mq��u<�]&�O{_��l|w��9�AA��S����g=��N�.��۪��Hi�W=�S\��։���*sM)����0ԒVܸ0ݴ�vv�`9���t��ì4�Q#��M���jMZe8~7�_v^&�`��X�/�N�Biէm�Ų^%�Xv�,��;��I}<��m۵`���s� ��ŀvl�`[%���$1�-�-ݶ����͘��d�n���w�JλTp�.�����&ղ^6�,v�X�BR�*�\�<7Z�[m��k��2�ea���1��u=ca뎰:ȵ[�T�x�ذ�Ȱ͘�v�;�`�jJ�9������&�~��I E"��~)����ow ������hm;�����?���X��X�q��l�v�,{���*m��ʴ�;k �{�Se���`ۑ`�8]'V*LMm�xT�x��X��X�������$�n��!��X0�tʶ㞠pgMr��*m��f:�m��qoi��񅨻U��ۥN����� ����;�ذ��Xd� ��B�@�[v��;�ذ��Xd�v�,�Q��ՙ˶m��w�����p�~Y$W��H1Bx��DP6��A�=ϻw$����rOo��g�4�Z�V;JӶ���/ ��� �ob�6k�`kS�DM:V]X��7x��X���sˀOG�.�xk��Ҙ93@
5�R%ĸ��-�]T��۲'�Ǧݗ��Ma�^���^ cx׉���:�����Xd�v�,��LE$�un��WNۼf����/ ��/ �ob�;4p�N�$�v�v�w�qvK�"���;�ذ��X���������v^���]�=��}��:p�"� $`�BE$ D#�"8�I��I9m��-��߻)Z�u��w�uvK�6k�`]�������}�;�1��ia�����؅�E3r;�\��O��nx۲��Cr4�D:v�ݱ7|z?5�uvK�"���}��A�}��"�*x�ڲ��m���^v^��/ ٮ5������mD����T���;Bn�-����^�\k �엀sCi�$��R)���n���x��� �엀Eݗ�w��Y�M�Z��wN����;�:�%�we�]��	�j�����|@�V�)~��$�vfKnY�	4Xm�(˥b�Yv��q�ܰ����/i��8{-b����8Hp���i;%����ts���l>@̾���֕�`�S��[!�:wny�D���.����!��Q��S�)\�����	!�nM7;�&v:���Nr�l��X�7n1vzȒ��������b��%�l�R�5��]�5�B!4w+5-շL����S�Es�.�n�f�5�f��М�ח��t47��td�9Q�ld�fQi�xBF�ɨ�fiS8�W�����;~�^��/ 콎�wah�պV�'L.��n��:�%������/ $6P�6�4ݍ2ۼ��^�{���o�x��,��uq&��'m��[���;�8�%�ob�:����R}i;(�i��ۼ��^6�,��/ 콎���QK#�>."�4��x���Ұ�*`���'�;���[�,�F6��0��u*�߷ݼ��/ 콎�.�x46�J�V:n�Z�]�<�{�o���Ȑ�I$FHն$�B� �$�8��w׀M�� �u(����m
�m�ٳ�qvK�&�ŀ{}���}߇���ʂgl� ��e�ob�5vK�;6c0[�h��t���0�w�M�� ��/ 콏po~�����gf�]������hs! 49�%�VZq�9r�ҖZCl�4#�bc0�66&���6�[�^�{�Se�ob�7H�F���'m��7xe�w�uM��M�� ��/ ��"��buj�۱ZM��:���&���UAW_}K���ճ/ ����4��n�6�n�	5� ��/ ��Se��m&$��O��u�j엀v\�����	$��?}_}��ﭢ�	���1`,���Ct#OAޫkS���c�)���a.;nU�E��a۾�_�� �/ �L�Wd���z3A�8�˸��ws�������E����#�V�)��+���n�	�e`�%��#��l� ��B�ƛ�cV�`���g�k7$��߳rji�����\m�B���+�Ia#1�Z�
�"�T(�d�I�{�y8���wQs�Q��W`�#��l�I2�]�x���iz6�cVV�48���_`ű��W:���wYmq	f;��z���w�qM��I&V��/�A�\�k|���Yw�Nմ;w�M�+=U��l����;�8���9��T:J����NӷX����;�8���96eao�����h��U3\��{�ý~���׀rl��5vK�9�8N��I�-�v��:����������@7��I=�<�Y�'�QW��E_��
��� EZ��*��QW� *���@Uʊ(��AP��T �B�T �B"0T" EP�	B��T  AP�B U��P����P��T"�AP�)B �U��T"�P��B(�T"�B(T"�+B �B*�P�$B T"�U�B(�P��T � �P��P�)B,�$�� !B"B
�B"	P�+B(��T"B*�T �P��T"�B T ,#B"�T"�B �T"�B
0
0T"�T ��T *1*	B(�T"�)B(�B(� �P��1T  BB�B	P��B B",B��0T"��T  �T"
�P��P���AP�,B�T ,EB(AP��T �B+B DT �T �	BB)P��P��T"0T"0�,EB#B
@T B ��AP��EB(AP�	B
�T $EB �P���B �B�T",BT P�� AP�0+P�+P�B"$�� 1 �T"��T �@T �B	B@T ��T$AP�P�B���*��TU� 
��PEZ��*� U����@E_� �*��QW��*�����������e5�� �-� �s2}pS� �!O���!�`e��@'S� i��Z4޹�Ӷ��v��E����А"� ����@=ښ hӦ��U���tY����+�GIfº� 
(h����  j�t�T���:.��K���    <�T�h*�
�M]�=;��N���r7��� ���k�x����a��`t�`��W�����8 �y�;�p��j;�� v��'-�hS��CE���Q{�j>Z9������{�  u����#[�s`5v���<�ֶ�<z��}����f�uO����� �;ZٜG�� �gR��� �;-1n��υC>À���B��۽�Vͥ�O�y�:��}�wZ<wضws�7����Xqz�C�y ��N����4�� Sx���>�u�=�{��O�M��:t����6�(��y�zS�u�GA���>l= ��ON�g�(>���()k�JiA@q4 �t s@�f�����h��(���`@14�{�=O)�y��)M���=����=g��� 4�u�
QB� �@����� bz:zSop=�����͸>���a��}�;��=ҥ;ۻ�\Ϡg�pT>����<��Y�O����]a�����{ϣS�s���}�;��< : ������Ć�d:U��V2��3��@������ͼ� ����4�{��|��;'�>�8�ր� d�����kx����C��ɹ�o��o��x;w�1 ��<��� OЕ6�*R�  D�*�5M�  Lʔ�m�J� �5O�j��jU(2 h��OF�)�T���C�
l�P� a)�'�����X�����������{���;��  ��5��p W@ �� ���*����  �� U9�_�O�����Hi6;tJ��\!];4No[����0�������� 񁤉� ��4o[9���0���l��s�~捳�Ͳ�����XF%"V1��%X��$f�/�����.j\m�fK�2�2ZKXa36&`|�Ώ��yYC2����}�~3}�nh�7�����ѵ�O��D�w��%ڐ�4��6����Nk>�l��߂]}��������K
~eay�L۽����h��Ѓ��5��^h/4�	�͜�����7��JY<�����4��Ƀ�����s>7�Sw���IBP�d�ٔ��MM�&���/P�x������*a��i�fs3�6���߸�M�^B(�E����1���M����7���~��֏�,�庌�����0������p��p�	���7���o?k��#�i����P�T��9)F����(�L~'���|h������r��l%���l��o4������������~0�s?~��oT������n�>����0�37�O���l�8kgߋ��BSg��# ٛi-�B4��e̞F��!4���Bi�/�z�R�_w0����.�0�sd!������0S�g�]�O�0�1��d{��>�_��L�s������;�p��7�Aw���>�����K��R]�᭒�ČMa
���c��K��9��������a-�>�w��]���		G��	)�o�?<��~Mguy�󤸐:f�|JF�����4��)�����/Q��(��m�^�.�s��Mw�?��1	�}z�j�����������&$$�%c,޾�����̿Ͼe��m�Pc\������qs������߻rr[��
w9����_���5{x^N�&/�}��~B���ၝX`,k&��z��~:�~>�>�C[���s����_�CZܼ�)���\����,{!�d"e��.j��O�w�/���c)�ѣt�͚�L�a�\1���u��r�?n=���_�_��>�\S{��'�G���}�xo߻���̚�`����������gqwq'�-�
no���Nn}��|N�FL�g\���0In����'�7���j�<�f%u��]0���_M�0��s�f��?fG����(~7���o���9�[X(@��O֝27�ӱ�SV��?<�}܁%:s[�3>�h�X%�U���_��̘��>�f���9�,x/�7�FE��}�����sa���%�a.~'�޷��>揉������9�Q?Ӛ�?j��?g7�_�/�0�GI�cO[��;���P�B�pu���.a/g�������t~7����İ����)��1�Y"�������c�Z���>G��!>!HZ��Đ0��{Rm���7����3b��
m%S��J7?�:V�*0i���a�.)�@���Mr��z	%9�ӽ�7���Tϯ?h��د�t����}�/�Ƈ��]X%�~�z~_�a���pNf���9������k+>�Ro��^ssd�K���.��c����RJ�O��y��Ԗy����'�}�7�p�kW_����7�P����Maаi����S7��}h���F��S��)�I�ȟ�ُ�.k�.ka
Ʊ ����Ǹ!}?C��L�i����	�����}�M~e�a5)f�~��Nf�Oٮ_ۺ��y�7�����.g��������E3�y5��%�ILHP� �H!
�a�j��@*a�|�y�>�?~Hfo��c�M����o������S�����n�~
�8�ILo���w���m�.�9�k��Ͼ3z�޳�8}��N%њ�0>sf$��f���7��>��Kϡ?���Yxɟ$���$�h���t�"�sF�W!`�H�2�$�2�t�2a�7]�0���w��=,�;�=/,���~�_���Ϙ�����B��?Sr�������Y�6CZ#:�s���&w쟧y�o���n~�����������5��!��w���[�M��>���a���v]��w�����כ���7�o�'������rd��������s��+�w3���&cq
k6������{�6K�����s�lHC�\�o������)���RHT�R4��
a
��YF�Jc
�+�B�0 �F�F�
��
0�d�(��i�(F
c
bK����k5~ݟ@!�,H0j�%0�$!%�5d^;!������{��~9I��a�S)�h����'�ϿrÁ����t��22R��@�
`F���|of���D.rI%e	���39��JrY��%%>�x~�oEL8����2��to����M��(dI�%XD������_ۂ�����_���~��?���K��i!aLe�i`�F���Ãf��G�����|����h�o=4.�%XY��t$ФI�]M$,HB�)!( J�hL3|77�5g7?M�l����)��ߎ�~S�������d�����w��;�3	! ��b������Hib�'fl"P#Cl�K��3{$�!]$5!I"H� 0�h�R��B8:`���1��4�ۦ1։�f���~x
��e9���4ۤ�P�Z���gS�����Mm7����x}��A�B�:�S���>'�8���M��?~��71`HCD)��Bef���q���FQ�hvm�a���1~�b����oM��I�,;���z%�0��Лѿ��o��Ϛ���orhK��n� ]���	a,�����a���.�w�����	��eK��k{7�nF��]��>HC�33���A��ƺ������P��9�f3[>3�nu~a�_w���`�?w��O߷����\�ni���湜fN_�����:��f��o�]koّ���>(�Ѵ��1�:HA��>Ĺx�޺%|ar���4��3����懚w��xw�'��wcq<�`{�Ŀ�d,�_o3��I��o7>���>�[�>�	�+�Z�����?�}W�~>���v<ŏ3��������,��\6�X�c�v9�?j<�7Ze�l�$���&���XK�玄�:石��k>�'��}�:�ל��ļ�����|�q����&���o��-��gw�~������p�(}��a�I��ߤɟ�~�ן�P����?�ss5������_�s�|��L1�MǞJy�<�ز��2Lg�\�d��܉��׆=|�͹L	�(J�͕��~������`�˿_��~W��g�8/�l��?_�~]�k3���-ݗ���n7>��f�߿~��k/;H/!�D�Y�f�f��͘\���g	�CD99s�na���>�|�����s�}�:��i�s�N���e�A�l��9��9���\ѽ}���3�WWFw�5��������dY~�}������[�>��X�ﳻ־���W7�n)��,�M�_#g�3go~�mX��''�}����	��;7�Lg5��}��)��3���L���Yۑw^'��'�;�ٹ�fL���;�3���엽�����I�'gwﷷ��eϮL1>��^����_O߰~�^��}Ø泧��rh�s�̹���8��B�!H]���Y߾�_Ƭ���q��
�����\�O�R��[�?�曃0a4~e��@4o���[��ֹ���l6o������0��]���s��ϟ���zt�8̌0��W�D��i�����ȝ6MS��=!�����e�x�;%�1���%��8b�>����٧z$��ߡ������~��ZX�����}8a�����Ջ�%���`���P~ϿN�p��p0�Kg��~��S�A��O�Vs^�~�I��s/>}ϸe�a�o[��]�߹���.g��K߿NŲM�f3f~ϲ���q�2�YI�c;��|О������?��䔙�ɼG��{�i���Ƶ/JR�5�g����˄ß7�|%ĿJC�{v�sq��t�%��q�p����$�4%"XĬX6IxM~?@ֻ�S��}f��$&]B�l"BF0�d���v��/w�O�=��=qA�bn�eH�-e�~�&k�Hq(bFeU�²I�e��X�$VZJؐ%eI�s���n��!�a�u?��s�w?}�����H�L����'�ٮC�?w[	8�H|5�p�2�㤹�U�!\!Lar���&K�١�>ZK�w���ߏ�xgMpɿ��d�;��g׫��z~��.���~���������d�a˼e�c�3�6̈́�a-���g���%��t�9��O@�N������q��~q������7����5V@!���6H۽6���SL�,�;9
_��;�A��e�n[�2�:),��K��
�*���)���S$a�6N9�,sY�737͒p���5?^�����ɗ��9˫�NI3/�7���~wf<)?������<ӴO��C7�ϊ�n����dIw����[	��e�Y�5��/�9�����O�f~�K��g�>�w�.p7�9��$xF	Ȳ�P��$$a$)�B|6N\�G� �E��FVP���ɺf���aK�z�o	R���0�sh�u�9���ˋ�阱������B����ޔ![��
n�����~�e���o�G��f�K�I��SB�Af��<��Zj�9/�q��m*������M��.i�7�-�		R!d�^NU�&�B4%�)/>Ĥ��6�dH /�W1�*h`�BXGC���/C>�%��B�D�%�4�����<Y�p�;�a$����V1椩c�v�ap�)�W���q�{F����;�]֦�ߟ������>M��A�eÇ����AC$#��2����.7�nl�� S�K����8D�Ł
��d��9�S[�Hr2~�}�}K�c	G@�33g�D���L4]��ߎN�h��������n��<R759��ǐŸ&)��}���o~��d���z�g��˛����wX��}_N���j]�n������϶��,٘&?��޵ǻ��Fk�ňĖ4ɯ�?�k��l��;ƚ��j6�!� 5��P0#r޷��r��k������'�ه��i3w_q8���c�Nl��~3|�_n����l?s�:!��0$�$d{��f�������ˆ�������ￋ���jc����a
c����	"�"@�� �$*$D"�1)���$[ �� �@���,"B@jb�(@#��1 �
�0 ŌH¡�K�V��A���
P�4CBƌ�o���~����~������f���}ӛ?��Jjo����ϹϡWN�������N���'������nw�d�n͙w7�|O������r�.h����A�`C�~�������\�g�w�MsVa6��..`WA.i�#�R��`�LjB�!HI���}���_Ĺ)�4l���~�6<t��f�~�������9�Ró㡭|2+���5���Ƒ5,J�̙ד���op���v�����F���Ĭa���/�^$e�t���At@*K���0a4~)�M��L��]���,H�z�m�}�/`��l>y�s_��-�?s��o��$���}�����UUUUUUUUUX�����������T�UU�UUUJ�UUUT�UUPq7e";Z1�j�ťCn��O+Uj��k�[ ��[�P!��5T�:R�5UP�1���U��ʿ����vҒ�UR�kE;$��ԶNXȵ@]*ʵ@+�;j��A�Z�p�`�	5���5U[r���AUUHYu
P�Ms=�B���z��͞Y8ѵ&�M�:�vʷ+&^�ڪ�V�sA��  �&f���*�Hsc(n�,N)G�$�p�v��8��Ժ���喨ڣN�宍u��j�y��kEn���Z�������+��u��4�́T���k/��6�@���ob;䗳�gV�)]�-�f��9�z÷��yk��hD!� F�R�A�/`��t��`�����؊���e�:`F%���.�=��#�6Ѣ�%���WU[/=�0t
�a��o�h��n�p��6Mڶ*#���@<�+N4�@N|�:2�c� q�h]�,��U*�顰6��K��V.�( �UUb��v���Q��YPΜ�� �o��f_0���������f��(�=j�we����۫ԯ�;:���R�0-R��$��%�U��ۆ؟d[r�z�G�]&��pʹF���K�R����l)x����v9�v1�N���jQ�˫��an�f�"J�U�rl�
��c��U� )㍧��*X%�i��u��ݡ̶���v�0�ِ{�I`�� m��X9,�ra/��	�<�F�*X���&�w����f�WX��Oh���3�5&�\�J�l�p�w]pm��g6ֈ��nA�	�͠y^a��[���X����(7]B��-��"=�`�[�Ph�Dpݱ�T�u��C�N��2�f"�+�w]�(^���kpm�qY�\y�i����ȲXЛ�]�uZ-C`+\Ԙ)����목�{m#�FAL�8^�,\Ů��S��&`�\]����چ��Ix-�VӶ�pVح��V���qE��q��T���H��TJ��b �UD\�,��vgER��a�\UUAE����5$nN$�ݼ��Y��U�W�I-b�Bdh]�KK�ےX�P�[�ɂ�]�XJm&��h�8 ��R�!2�&L�v���Z�aF��uAb�u�(#���9���t*lc�q0�p�����DUFmŖ�ƃ�r����@5+SZ� Z�4ٲ�ǳ�I����S����+�����\"�u��T�=�%��S�B ��b!��ҭ�unչ�xBɰ\jz{,�V��hwC��U�\1�v��N,���H�$bZ�еOul�q��O;5UP9Q.gD�Auu���;v��P ����N$��[�̪]R���)cmz�m�f8H�Hʫld�,�2�D�\�hEa�
n6�ޓO�Ҫ���m�p�6�ڂ�q�ǳ'�]mŽ<��u6q�M�ҬK�Q�e����┝hP�b���A���.i�
�[*�Q�lPRR���mlMǴAӕ)������h��pqR���`2�d��=��/WTKZ��n�p��u� �[��s:�+m�O{�[T�%Ms��U �%�Q�n3W�J8�ˡV3Գ!���fU�A�4c��U��0���i	GSv ]ƒ�-����屰M5�̥4�Z���4c�n�nȇn5"���n)fM��u'˳���t���t90b-�`��by)y�.�K�ɀWnkz�,�r۰�B�ڹ^N˘Ň�� ��(1�m�m\;l�E]����:��wl�2�Q�4�m]� ���J��E�\���d=�ۜ��q��m�L8�A4��
�]�m@Nd�.�Y8}�,�2�]�:m��0	J[E�6�-ˈWDi{,ճ�8���x�Z)WgGm��@@m/i3 �՗4L"��c������s�vu��C��y�Kw��T!���W��^@��P1F��n%[[)H�<\\���f�IAn#q�Hx�ڥ\��q�SVʀ�I�+�Z��h�-b�;m��i����'�޶��R�F�v�,���>w;�|���L<�Z7SUWm��ue�Gj��@uQm9��ma�@��ڨ�iea���n�jR��n�V��es�Ռ[UT��7N��UJv� ��bj�`��L�Zn��A�YACM�CK\k:�"�\��Z�g�:��.���D�"qj�I%�:���-�	������œ7��ԸSh�Y�����Ma6��F��s��7`��r[E��5]���
JR��Mi�%QU�6͂⯒��5�q��J��<�A�9�TF �Ʒ�����tEUC�s�3U��J:"G�vK��j������kqڨ޷
���Uv6�Ξ��X��@��c�%�v2�c�x�Fx��V���{P*��\	�LWMR`����N�Ų�øo���D]�t<J�-P�;�J�k�m� *���Z5=.�$���Z5�T�횔�h6��i��]K��\˺��[Vu&��8�U��U�
�]TY(Χ��Ul+eGX�UA��URx�v��UTUS��UU[UUTUU�UUA6�p*���3�GaY�D�R�UJ�1ɶ�;uT��WmUF��ī�.�䶪��jU۫�m��$�Sfwl�-�*�iIm���#UUm� �lU�UP���ʪ�Ut);Bꪠ�7.86�P6�����V��&YZ����Sj�e�*���&UM�D�uUUUU*������UUUUUV���!�n{�0�Pn�uWUUV5-UJ�TSjU���렢Z������5pqUu]U�`�B�2��-�����y�n�a�mUZ�j�\b�6+��J����j�v�n۫��UWh
���XFڥy� �UՔq�3�L0��[lT{ن֠
�+r��[cPŵV����K��R�U jdx�N��nݗM@�d�`����j���Vj���UU@ST3�U��� 686���[���ƪ��Nf��)�@ a���j)�滎8�wI.�W-u�'�8�Xm�!]��`�<���"�e��bCmpM���S-M�����Z�C\��[P���s�t��ڃ5�m5vP�5�0ht���9Wv����͔'��P�*��tkpeƛ&n�F6�P�j���]X��H�و��m��ڬ��P���٠��ICh@#+�>�����OcP<�86kqγ�i3ѥ��V��<午5^ZJ�eU��8��kEF��s�[*	T#���%P-���)�����/,cQ\WS� v�k�d-;ju��+X9�5�p `�n�TݞĦp�-On��uAԫp@���r��L�K^3�� �cn�ڒ����Њ� Ъ�*����
�`�힠��wfb.|��U�\���
�	�RN]���Ks��zqM�jL�]���ƉL��UU�mP㣥�s*�5]���d��9��	�h\�v�OTuÞ"v���b�������j��R���UUT۪�V8*��`��z��ym����j�@�Q�yj�j��mȈ�W��A^]�x7�˶@
�N�Z�e=��z�f���@��]���V�@5mU6^$�h����8*�(�UVغ��
8Ș'�q{TSs���oK���3bh �m�JM�n�������O)��o�շV�A��]�U��:�
�
[I���r��c9H,P��R�Z��k�n\�UUV6���L ���;8l3�h�e��j���P#;l�UVҹ;u�L=�vY!�*�
����P�V�]s|o4
_2ܻe��P�B���j��� (�k�-��f�9 ����6B�ࣂ��燭���v��ڕ�v&���UuUJKUS�U-�Uǭ�<Q� j��T&��	�������Gl����(�ڪ�j�
�U�\���UT��hᠨ(*��U*���1�ڕv�������R�JT�mUb�*�T�ch�^ˆ�T��a}�^�T ��" 
�4ͯ���ʴUP�ӕ�ۜ\,T*��$�IlT [kt�
�h�M� UF���V+�=�UV��rӓl���J��A��UUF�����j���5<UUUUU�*�UV1U���PN�
��W/-\�@e�R�C��0��om�
���IdiV���UT@*� ���*��<�>�P%5�Z�UUb����ݍv�j�d���d�Z�RR�����Z��������Z��������j���VU�V�YZ��8���UU����������Z�j�����b���U�m\��M���UT說�
�۔�yڊ�lWU[]TQ�J��,'�V�]UUUUUUU��d�p��٫a��WlͰZ ��j����h3s�m!�Kk�����;SӲ���UJ�J�UUUPUJ�R��ڪ�*���U�+j� 
ڭ���UH $ ]��K b㓬;� W(]r�mR�UT+;؞�@��Ի5T�Kuq*p� O 6�*յ��Q�ԫUmT�UUV�]UUUUUUUQ������1N����dCԾ�B�UU@UUUUU@/+�l�TmUѠ$r�*�\U8+����b�������ܢ$�s/-��a�n���je|�_;�z�[l�dUV�Z�(ѵ��v��\��Pf�DOBdC���v�J*�J$��Ih����Ԫ�Z��sU]�J��һ�j����tʪ�&�:�4&y���9Ÿf�kp��s�*ݐ�6��A���������������X��]�H�)Zͥ!��
�RY�[h*%�ĵ�`��.�	��Vť��9�m��뤍m��v̅��Uv ,ԭ(��Pba�hF�V6兄j��c[VD�c�6[[c�h���  �TF��
�lT
�a�W��� �,P	
.�Tt�AY"H1? ���
С "��p@x Q�%W�D���?DM�b����l҈q�T�j�B �N�P��]�8�"�/@��AH��8� S�`
�mA� ڃ�M��B��_�^�� ����T���*'¢|.
�^�1Ft1O��@��"�����R
*T��.݃���v��� Lb	��:(�؃��C}~
�(~z0� Sz�"�ؑ��J��Sj�A�P�pt�l@�<t�u80�@��L �lO��CVO�S�HE���D$T"D#�U���XT��2
� "� ȄH�T��?����$�X-PʚDv���S������DKY$�F0���#"Ā`Đ$�"��D�j/���'�P�
��"|���I# H�H�!�@�a"�	 Zj��h��@R!������v[#llB�HBB��V	-dB�J���@$U�))[IK%A�@��!�"h�#X# �*��)$@�	�w��*��
mX �����p�p W��+�ъ�kX$(JU)cR%ZR0a,c�D$M��T�qXg�[u�kY��N�ҳ��ݗVMkjn�:��M�+i`��p���u�Ms5�:{�F�Q��f U��X�݅�SHI�l�h$%(;<M(p��[ZU���^%�����H#�N���,+��C���E�,��7X��RFW9ez�-��8Oc`�1�L˂�Ie�-��j�M�t���<Qb
���(� 痑��c��c�*�Vd�ġ%�!X�1������{�š�n��>SO@m�]q>�P�Q��%���y����[ �9;c�Eg�/n]�Lczw�S;l�C:ւ�s�A7K�E�m��� �5�Wbf�`�JEYkQ7�x�𠵘��.�1�{W%	���i+��w�`vx��5�I�p�U\�'E����ٕ��ey���gF7b��.�B���6�#3V����-2�܄l��
�b�1Ս�f��X�BV���y���nܽ\�8ל.G��M/��ӫo;�qb9Nۖ6���'i���܍��P�DlA��.ш�nx�W[�'Rg*�v밳)�t*\ve�{p�i�`;h�������6$�M54����Dvw5.����T@��b�P��aκ1A�-)1nSh;�F�-�Nہc��ǋu���f�>��b�;X��s��tW��-p��N�4�8�,�l��w1�v�E��=�=yܑ5ݍ���n9�����x�}<3`fgT �K��Mh�5 씅��4ڝ��ss@YCa���mٺcn�qt�6#AC�i�Nǋ��7=���1��/K�î5it����f�De�X��`tZ4���� �goKg:e�UW��8�-�d��[�;X����MWUU�����[TeB��椠�dPR��t0��݁��.��^&iz���%0:;e����Edjё0>�� (���y�.Ul&'X�6�f�v��i��iN�r;�N���rE��b�ɻ5��P�1�F�%�f��F�A�PCˈ�Q⫱O "�G�	�H��A���8�q1F*6I���b�z�W�gv�"\��WA6T�xP��a	�f���׫RU�VڢM��+��S�k`,ʯ��'�����9c���=-�h��<���;d��&�7cvrr/�b�Ǳ���Z���G�ɺN{s�l�Z׋2&:q�%�#bK�.��0!�­�дp7�;q��=�xT���7r��@s��p�N���Kz�f�SK5:t����&�ww�-�ْe̲��c��.ܠ��C��;>�;s�L�1���i���N�f�޾� �_z����s�]�����
D��Dܚ��h�V�k�Zm�@ꫥ���pĞG �l��k�Zm�@��-��î�X��A��R��h���h�l��~�Ų8��(�'"�m���h�M�ڴ^�|♰Ԭ�8�n��!Y
�B�&�XR��a��l�BvKP4Xe�p5ڈ:����?xZ�S@��� �٠}�@��a�Cp�H-�)�f`����&T�F9J���H�3��s>�s��n�z~�h�E�}������F�Dk"�*��@-�i�����-�~��>Uto��E�9&��@-�h�E�Z�ZW��~��+�H�1&�mɠZ��k�h^נ�4g3/r���%[�Ra������`�8��#iq��t��2�V�c��&6F��U�l����oyh^נ�4]��:�\:�ŋM���*��@-�h�E�Z�[�s9���-��CP2Ljk7$�����;��e�����"@c	F A�Ũ���\��v����}mx7��� F��94]ʴl��U������� ɍF࢙�k�h[^�[l�-v|wm�{�M6h�dЬ.�「�[u<�::�τ��q�W-x�6Ė祇���L�@����f�k�V�k�h�Y��<��Ʊ4�zm�}��31#�~�-�~��*�� ��q
����H�&��-w*�-v�=��K����{ޚU],n"8�I�s"�-v��k�m��y�9�C��A:�w�f���9V}�H2(8��ŠUmzm�@�ܫ@�ڴ��#"q<���)'����zn��uB�l5R�Rh@�Ɣ���Mh��^f�T*��1��S�� ���Z�U�Z�_ٜ������;�y���l�&I�Z�U�[e4]�@-�h}P$�^L&8��jdZ�S@�ڴ�${���=����;���<�Œ6ډ����9���=���4]ʴl���U�o,Q�BH�&'�[l�-w*�-v��j�g1w��	���S4��I�����HW[���B�l���Ws��sfKM yH�ġk��{hz�e�Q������-�ūU�m���s2�H���5B4l8���sY�X��F�4E&!͍)������{C��åG�H�B����65��y1-�v�Ą��1�Wa�Kv%�
�����z8k�n@���q�F4M?w5F�f��K54�0���f"����Вt�5� ��[6%�*Jإ��h$�j��kn4>1������YHhf�r1�*���m�s�@��h�V��mzUY����pĞG2-��o�s9�H����
��=�r��>��,dPq7��k�hVנZ�U�v�V�m��HL�0s�NE�����*��=�~�-��h�V����މ��H)�k�V��e4]�@궽ٜ�fwo�
a"�$�����Q뢌]s��;E��cR��0V��P�A�$�Ly��2/�_zx�-v�������~A�?g���|�Ǜ�D�q���շ���\�ぁ�!�R�+AsB2�J�	Jq,���"]-n��Ӊ$��RI�#�GB/�Kw�^��疁�e4ʬ�yb�b�8<LN-���]ʴ�)�Z�Z�����sQ��=��g9�ޞ�-��Ɓk�hVנuU��H��b�$�9�v�M�ڴ�k�-w*�>�:��x�&!L�C��nJ֩�g��,Ȱ�&�*���eN���[�Gj�!�Z�ZU����h�S@��[s���F'"�:��}���?g��}��@�ڴ�Օ=c���G�Z�U�v�]������&|��w3]��Wֽ�E܋c�H�E�v�M�j�:��@�ܫ@��׏��&����-v����]ʴ�)�uv�#Cq�cF72)��sX�ۣ6kKX��!S�瓷WF��d�͛
��78��18��k�-w*�;l��k�h_��J�E1qcq���-w*�fs/�<h�����mzUY���DbO#����Z�ՠu[^�k�V�Q�l@�ȣPnG�k�hVנZ�U�f}�s�m� �s���w�vK����F��(E�u[^���3=��������k�h��Y���0A$jF��)��1m�r~�>��rl��]#pY�[�Opm&�	$����yh�ՠZ�ZU��}RX��E�8�P�L�@�v��j�:��@�ܫ@��׏6B$�	'"�-v����]ʴ�j�?*��剸�&'��mz��Zk�h�V�e����'�ō�#�@�ܫ@�v��j�:��@�qp�s?,����<Q%PC%ʌ�v.q����]W�A�[��+��1biT4*ؕ*u��T�i�[Xn�V�S�Sr��b%@7�\v��\64�$5�	���/`�]v�@Z�iR���j�=�\����mF�-�."�x���_,iŷ^�� 4�%�0���:���9��v�����i��m͐�`݁T�[�y{s�;/e�XkuŌ�"|���N$��WNܦB�Jgc���x�[d�1�<S2����!4�U�v�v�v��)�8�"�|��Z�ZU����h�v�	���7#�@�ڴ�k�-w*�;]�@���H�8���ȴ�k�-w*�;]�@�ڴ�t��؛D$�R=�r��ڴ]�@궽�K]ɋ��DE2-�ڴ]�@궽�s�o����Z�0�e�16q�%��LTS2E%��h ����3�6�53�U�u�G $�@�ڴ�k�-w*��g9'S�߹�ûo��}��0��:�S&䓽�u����,
Ā�
�#N*&�wy��rN����I��{w _���ĜS7#�M�r��j�-v� �٠uU��E��$�9�h�V�k�h���r��ς�mb��7#�@�ڴ�f�k�V�k�h�32凟�#�p�g�0"�,,�Q̀IL9y���>��i�݂l�ˁ�0���-�?��M�r��j�-v��*z<D�s��-w*�fs������?yh���fq#��K{rb��"���?yh�V���9�9�0H~-����ĥ�bO��!ͼ^:��3�4F������WG8���Fś_�ٙ��0F��F�T�x���������0���h@�ٟ|�kA�������ߋ���c��KD��;����@kO.	�8]�~9�5\�fN�%l�ow\ഄ6o��-?:~n:5�;Ye�ԁ	x���?:�ʩ���\����i�0�u���3'�0�DvN������I�HZHI[f�!  �8��Z#���d�}�Y�p�0�����f7/�O���8F��F_���HLq�0�e��ksl�o0�;��,	� ��`�0�����*R0f���9�L151��{ě%l��7�$�f��g9���&`H���~!���lU8.�S��QP�EDM�C�� ,j<�b���$F�Q��)M#C`��C��
?�M��u�'�g�n����3fH6CpH�]�@-�h��h{3��^����}�ј��q�bqh���r��j�-v� ����A��<����xEM*qΚ�Y��b��X1� �!��+����N<r��&�k�V�k�h�W�����{�@��/���"r,I�s"�-v��j�m���[��Ċ��{��4�H�F�qh����[l�-w*�-v����&4A)�P�@-�h�E�Z�Z=�{�9�p�(D�$��(0!�(��$���s9��vyh��Q��l!��4]��?g�33�����������y�:�`�m	Z�9��7 ��׈Ɠ[�G:bǁ�����%��7\z�uR@�_|�_j�m���Z����̐l�dpȴ]�@-�h��h�V�~�Gc1H(��@-�h��h�V�k�h���+r1q26ܚ��Z�ՠZ�Zm�@�;b�92G%29�h�M��Oy~ ���Z�v�I�
@ւ4cbS!	::�O��4e�,t�r#$Ht��l;uf�IO%�p���z�c��D���0�d��Ԁ�ή��	�uj�� ;D�����R����j.jK����KŴ��f�ԈS�T0����C�֋+�2Pٚ����ǳw�	e��1�ze*e��ݛK�Yx1Jq6�u妺� �#sh]vxݚ��.�IZ�;%�`�b&���6�)��M$�}:��OK�oc�[��e&au
P˪�w6�D4BZؤ����\���m�>��mV�!�/#q8P=��- �٠Z�U�[e4{pOd&<�S�<�@-�h�V�m��-v����f8)AI�I4]�@��h�V�[l�>��.]ɋ�$��MH�]�@�ڴ�f�k�h�kǛ1�5�& �Z�ՠs����{������k�h��#��MH��$�4˝݂���B�u���;�k�f83l`�t2sN��Q��@-�h�V�k�{9���? ����ݬxx��94]�~�s99�s;���{)�Z�V�[l�g33�ye�Q�������@�]�@-�h[)�w�a�idq����w�ՠ�4���-��{h'�)��)�P�@-�h[)�[e4�ڴ/'RI���X0�����k]m�sq�ҐC�(T#�4f�8,ppE����D�H�I���Ɓk�h�h���b��ɒbq�4l���H���@=�zh[)�~����L��8h�h��>��r���!�"�BRR��������
F#bBVY��f t �߳{צ�z���c��nD�����%�{�@�<h�Ms��Z��<<����$�M�e4ff{������@-�h��g/r�����)t��0��e���j�����5�馅��TD��c�K���:�.O�o�ߟ׻o��ՠ�=������Z�Շ��K#�8�N�v���g�s9�l?�����|����m��s3��;o�OX�����r- ���}�jz��39��{����7`��~��h��k2�|�uԛ��� �9�/� zo�7`F���,V���2�P
;��=�s���}!]�h���8�������<� sޟ�$��k��K���з�ِM�+�������'
�^ź�<�ٚ�qf	?I)�����0챍�o��p߿RI+m��$��k��ͤ��o�ߒIv�M�5fk���7`��|�����"�s��� ����� {��m�6�sߦ��E��r�_< ��� �����ɶ�nsn���<(S�}�[��X�)q�I%m�~��]N��$����~������t�%�#i0�һ&o� {��m��ԓ��s��� }�k[����}���!�@�a	����=a���^�sV:ݸ��[X�eSC0@.ծ8�̛�мB�ף����2Mn`�@�l,⚒vo����5;θ�̇9㷫q�Ls��͂.��ׂ�>���s��Q.�k�7I�"�.�n�����n��.�%��q�$�D�=uYJ����9�F�Vɞ�<s��Mֳn*�њ�rj�nu�@�C�:�#P��j��k�YӺ~�����V-63T؂��Ĥ��	�5 �@֚��d�=�%U�%�	VmY�L1��I^�OߒI.�&����?~I.�~۰�g�x�tsl5��r�x �&����?~I.�kz�I[l��$��l:{�:f����`�}��� =��ޤ�V�?~I$�l��K�����p���o��'RM��v �8�� {����m�s�_< ���m��s\d5��݀�}���o���s���$�ݭ�I/�.��&<�8�3 �l�@,���j�TshX�إڸ��SG���9�K��Wk�5ʹ���q{ >����x��}�<���< ���H&�Ĝq�4I+n�����~��9��$��ZA�)��c�$a#$���!IT�`�Hr���U_.��˜���m�����$��\�g8�J���=�D��#q8~��U?y=I$��~����b��{ 9�w����6ݠh	X&�bz��s��߽�OߒHW�sRI[v��$rI:�g�7`�O��5�Ya�\˲��=��� ~�O�u?~����7���}�Ϟ {����H����jv�e�k�.�vy����a��l�1�Gi6����v�[��������W����_< �;[ԒJ����g�4�WޓD�ﯛ���6��x�������e��~|� 9��� }���|�I�>>8Mز�S!��v� 9ϸ�� {��ݺG�U�Db(��D#���Px
�;�?�����T�n�7�!}{��"m��I$��%�fq�}�5$��w���%��oD���{���� S���pf��+�ov��$��9d����I{����K�ɨ�~�}��n�f��j�r%��l� W<t���^Ă��v��-I�ޝ!�WOF�TF��� }�9�`����� �l��g?6������$������iDH�\.݀�{�������� �.���$�ݭ�9��V��y$35��35�r�mｭn�o{��9����ª�o߶� ?~��� =��a�;e��7!r�`ru'Sns�9|��ͻ ��u�[ t����G�"E|�<䓩����� {Ϲ�������U�x��}�`�ԟ��H���Ͼ�?~^������ ��(�dњTuݠ��h�d�U���/<v����6lv�zI%}�C�eX�n0a�m��}?~I$�l��J��=��s>���~�}�����j�n�r��x ����*�o���s����{3v�o{�u�x�u:�`8NnD6`#C9�� s�w�����rI:�ls�q�� ��^�w��>���F������u���맏�� ����< ~�{�RO�u'K����y�7?M�n6�J���M� }��>x�N���RH����ߞ^r�~���ݶ��ō�(0�*���~aq|�)�+�ؔ��)�Lp�M�B��� h����̄!	YK����?T�&S��]$������q�
�&� M2�@��X0��ct~��C���)�G �I0`Bm U�V5ZYl�ZB4I!2U������	�Pa ��$���u߁��1)(����B�(Bˁ�L�8^�D��*�������̒N$!	YC�e�!.��R&�_�S	sZ.'�00�X�KK
M�fe�u����.MU�	�ǔ�p��13����9h��"�����ֳ0�F@�JM\��M�s�6}�r���e��RR�K�2ɻ��T�]I6�kZL��e���	�)�"B|�M���	oR��y����m�l�;ʳ���V��q�v�%�� 48d(ti�q�u <�X���6��,pRq�]��b+�J��z��t:vg[Żs����q�����z��3w�c��+��Xᓋ`N0e -���!;vpg����Ƙ��\�91�A���em*m�d\1o0nz��qAivn2jQD5v�0D��!*Ky�������h���ʑ�93iin�4���ҔR
��౴.��&;qf��6��,��@fP�8ӵ#�ef�l� F[�(��*ds��Mχeؤ�Up��[e�Q�r��-���Z��2nN�ɥ��%熣P'�]n��X�v4&�rmvˣ���x�Q�76.�;d���1	���C Ű.R45m�X�\#Þ9�l�㮕�xx�/�C�	:��eN1;��۴��̖�VqvЋ[i!\�M�o7>����yc^!%�{���JIR�Ƥ�S7K(�4�7����m��tT���b�0%2,VZ�u���p��-������]�6SrD���]Z�%�j�mE�s�n�:D���2��s�t��[s��q\s�U��
^ݫ�:��T��6�F��M�9�cu̅�8��b
JrV(4��k6���^zg=�	;v��r��w�� vl�)�.+�𭏊�MCpj���F�/Fl����gaUy��β��5%P���iiYk[��%X�$-�0��X�9���Й��U2ڱ`�d�v%Uun�,��z��;�َ��71���A#Elaq��h�uWU�)h`��CM��Ӷ�9��f,�&��f�X�!*��vʺ��m٣q�lڀT�U嵍� ����Dj�"�cz��D��UV�ڕ�2.����V����%��R`�j����B] �����H���Y��U�SԵ*�`�j����k��+ts�n3p�Ӈ�B�6�ܗ�;�:��%�#,jZ�&.���m�;�n��98yw��ct���f��ӫM��
�K�kqcʴ�
�-�t[J����w���'�����(��_�|���q z��~U��>Γ���:O���\�E�4�p2ghz`�g׌���B���hOhD��hPR��3v�;ɉwv{ ����.��ۦ�a��u�^8��4pNt���ih� �m��Xi{r���\&�����S�2�)��=�A��R��"
B�b�b�g!��]k"ks��^-�dqّ۞�Z�!��e��.�5ݠ���U�㺱o.�Gٸ�B�IJ�Svfr���I?wt���ai���SR݊%��GO����cM���	��K�.Ѷ"L�I:�;'a��Zj�m��� }����Ͽ^r�~������m���s���x�tlem�9�ʽ�|����~�Iӓ�~��`��?=�P��}��'S��{�sjC%�j��)�m�m� }��>x~���N��ӟ�/`S�矏<(z{�&��F5[��ɻ�u:�s�q�� ���RI[ݧ��/s��u�y=I%�U��Ƹ�tk�U�� ��I�S�����I*�����V����_btea���[�05��t����.��u���� �KfT˅�ZY���t�����Xf�e�[}��Ӝ�߳;���m�����/��ڴ~���9��5#��-�������
	k"��IB���d�[i"!
���������$��&����O߽��q����ޢ3b�긢�� �>����/a���6��|�~~��;��ȕ�"�D�I��s�ĭ����Y�@��V��9��I�?~�������w��������[�M��g;��/�����٠\=��l�F�:c�K֬���a�f���X�km�^���9#��6�:wO{�]�0�7aI0����٠����fg$�k~��wm��?bn̮��-5�4�پ��3}�_;�}]�}���$v���Q<X���4�znI�s��ϊp�'�@�v�~��'�_M �X��#Pq�)rhg9��
�{��rN����ܒw�w[��������^"d"�7"��>]�^s3��ퟀ;�zh�S@3���CfF�I-��:���k�"\<٤h��ˡB:��Jdx��N�;���=5CA�8�+��_M �m����g39�U����dK��7�7�@>�}�fs=�<hW�zol�s����Y���Q(����=��f${��@-����mOF�q!c��hfg?����g����{�h{l��@?EaH�0H0 tS��t�$����������MaP��-8���h��s�39�~����?-�mz�v'"S'"S!&!�H��z �H���.a��OQ�H�VT��o�N|��&�cPx�9#r~ �ޚk�Z�����s? /���_,^�)��"PjG�k�[���s���9��= �����w���9��$�K�Fq�#�@������i�g3��o�4.�=�ލ��X�NDĤz�fs�o��[�M��^�������y�\�"^��,k$n �M �m��s���fs�_?�������l�&g9Ü̿Rı?�AnZ�6xz���!*����-؎�gb{rW�qW�A������]�٣�ҝ�[�H�kqv��f嚛Z+uX4����Ok�R�5�k2��!Ʌ4S	IBQ`����c`um�`�]�n�i	a6h�
��f�)c!�t�@�`�17U�,p�kiQbb�1�aT������^��nFZR���U�XJ��ٌ:��6˜����O�ӻ>��k�^,yQ؆���XA����X�Fˈ�6�i� Pg���ɻ�.nlq��HrN�����w�ՠ�����~@w���;�y=i�8��I����ڴ��4�l�*��ﳙ�Hﯚf�H��� ��Z��M ��4�33�w�@���@��Fݮ��a�S/v�u$y�=�_;�|�k��fq+����)���R8��;_j�?��g9���g��������߭�Q�:��k Bf\	���%�w9^*��f�%�)a�ڶ�"{9��i��D�nH��W���v�4�[=��~A|��uZ6����M]:�-�f������-N�.I�{�ܓ�g�w$�{�sʋ���?�ydK�ȱ��8�94���h�է�9��U���_{�@���t�'D�$��s3�����}���g9�K�ޚ����<mLs���>Vנ�� �m�k�hw���8�*ڂ�c�v��zg��Ui�h�q�5ڳ����tv�{�Oo&,�J18� _{�@;�f�k�{9��������;�6?"!�$RM �m���{��]�>���rI���߅D�N�b��4�ȔXԎ94��Ɓ�4`�H��D "��D�,�Wj	�
�;�{[�}}���R#	�$�o���9������}�v١�fs���{|h^�O�,�c��1)�w�����f.�z~���|�k�?�3���d��ݺ��/��zյ-!k�e%����Ib�hN`wG6NKH��rtU����zh[)�|�k��fg? -����\1s�LYĤDRM�e7ٜ�Ď��= �ޚ�m������3������z&�FLE )�= �m�{9�Ď�zh�������G$��ƞI"��{��ĭ���v��@��M�T���oٹ'��3'�n�ŉ�#�I�v٠}l����@;�f���s9��-��	��Ć���F��&��.v���d�-�����Qen�$��źA����9>�O�@��ՠ���s��ޚzy/L�&�xㆁ�]�}��$��@;}�}l��fs3�ٜ�ʯ�4��Y �'"`�Z�M ���=�Ļ�Ok����Ϋ��ȱ���(���31+}�wޞ4��h{l�>�r�1d�994���=��識� [�M �m��s7��T�L��F/\8�:1,ڌHTk5ne[h�u*���bfF�6�&��+7BP��&�JjR��#��5̛�&���C��f�&�9���ʼıI�T,ш�Q�F���](�<泎r�#S���-���l�5Ů(�G+%��������}�,t�X���Ӄ*��ngsN8G�ӳ�0S�BӴ0�n�QZ��)I@�2���\锚�A	wko�����x���;�MX�j�Ȗ���S�\<\�{�1e*7#K�˶���I(z��# ,�@R����w�� ���g9��wޞ4���h܀ǉ�HI�w���33�zh����V�oT�ơ1c��$��l�>�SOg9��U���[�M �X�H6�LpƤ�ɡ�s3�����:�����h���g�g9�￿��z��1�#�4�mz���b��;}�~�~��}ǜ�Vc\�+[c����1���m&�E�x�-t1̈= 	ź��Y&JNDĤ _{�h{�4ݲ��9��? �{�z�U�ͬn���M�O�����:Pa8�HF�X!�qTvc����@��L�AH�`mM�El�h"��`�s��<������M�>��@>�l�s���Ď����&,�<�Hֵ�'��^��r������*�d��4����>�n=mb�b�Hh��������g3���/��Ɓ���y�R	�d�)�}�٠{��s9����������ٗ��	�IyH�C��n8n�l�Vn
M���L�2�'.���z��t�r;֐�f�B���m��?v�h���g�s9��0/��4��<��i�D�H�@��)�~Vנw�h{�7�33�9��l=��/� &8�Dy#����������&,A0�Q%�H�x��#�F���U��2%�222��ß�O�R����)!��,.�9�?��i�}1�k�HD���y�T5�1���$!D�$`ˈ�v�I��զ�9��@��$�G�q�ȅ)�#�3�a[��E��B�c*��(��HB#&�����&���ɭ$3�sq!�˭�?��l�i[)F�e����)��������C��ѻWI��&�H;*�q��K��d�i��%+H30��tCzہ�D�,�W%�� �!!!)``��b�M2m�(�J[g��K 1`���Rf�`��"�"�&�H�63sf�l(Q�HE�� HĄt!nR|"4D؀�� TD��J*l�O��|��
täM@"&�
#����!چ ��\�޿w[�{�k�rN_��s��(�'"bR=s9�Ļo��[}4�v���:�Vcx���I&�w��@�s�Ϭ���>^�����n��~_�p[��K(�Yl�C>���@H1-�Z�a����p��Q4tv�O�N������œ�H��?�~��?+k�>]�����$�����'{�]K���ɨ�Y��Š~Vנw�h{�4�v��s��z���ԑlm�"��m����i�����9�7�?��u=����!1q��ɡ�s��J��|����r�����QE�$�����[�v����$y�rI�~]���3��?{��m���٠s���y�	0��,Ny�\=h��D�@٦3�I��>u	�4��?I$���wR�̍v���_���@>�l������? >���:�~R9#	9������4��h+k�s38��Qd�1��x��)$�}���Ofs1.�{�@-���;��͘dĜ#@ܚ����s�}����h��- �{f�w���(&���b�C@��V����W=�k��{���ܓ��7$�iڒ��� �5`�Z�F�L�gVe�*;ol�Q7df���/>Ų����u	�˓�2��	��(ц!�m�g2/fJ�8����n8,�����v�&����gl�q�o6=e�u'��y�m��ZH�wǮ,wTp��+(\���-����2L�V0�H�iZɣ(��f�%��L��6�l�f�	�eɕ�� Nxw�t��졉n�3�t����I:��($s��dň�k۰��chݱn����n�<�nu���������(
�w�m��~�&�w������ڴz�cC�����R'&�w���fq#�zx�;��- �{f�9�H/�����<�N8��>�����Z���?���g�������>]EJ�1��9!�}]�@;�٠�C��8���Ɓ�h��GȘ)�w��@�f+}�����@��V���U蜍D�bn6��eHCjV��]K_���<`���Yfa,��Z6e�\r&<pM�H������?[)�}]�������@���l�"�vL�krNw����(�"@0����]�>���ܒ}�{��}���y\\YHhWj�;��i��bE���>��������M	�$Zg�8���zh��@�����ڲcMx �b�4'3@;�f���M��Z{۹�~κ�\~^u�6�u ��,-$x`�b�68�:��JY���;{�!�WF�"��zx�>�ՠuw�������ޚk^k�,2c��rC@��V���נ�@�l��9�$u\���#$�"`�Zm���٣��s��9�D��@�$!	1«U\�s��3g}�Ɓ�;�}z,�I��RI�h{l�?[)�}]�Cٜ�V�M�˂�f��"#��Mɠ~�S@�ffw��_�-����4��Sd�`4���eh�RSP74i��h��s���6G�qGVZ����4N�т��}]�@;�٠���s�9���;��?��{���<P�	7&2H����s31 �ޚ���}]�@��&4�"ưJI#NM �m��e4�s9�K�~��o��v�㭱�8�8�C��3����Ɓ�?yh{�4Μ�00�y��pm�4��h�,Y1�(�9!�}]�@�s��Wo��}�~�S�m��~�c�����F�V2�5FȚ�"��7u��b�ka�ن��T���;-C���"`�_���= �m��e?�$���y�ûo��8v�5��PUhݶo���fs;���h���hu����I��N��>���{3GTp@�;���huڴ��V�}�f����i5QG�&
E��s��{�@�w�@>�C�9�g�9��o���/����,�BMɌ�-�ՠs3��ޟ���yi'ﳽ��lz�b$H�l��E1	�"��y�(>=u��V�� ��h$Hk.,u0=���p.��۳�q�t7	D�l�6x�� i���aH.��3+F�f�)E���.���	�kY!������.�.���]�N8U���/.��za����]\��D��!�48�y���6��B�m�7��t��o��@�Gk��3/4�*�;�A���-��*��O�n��Ԓ��[e%�ɢ�Z��z���9<.H"��a�*��&%�HP��^�̓�a)�[{TK�m5����t}}�@�n�.�&F����M�]�@��ՠ|�����m����D�M�]�}��H��|���o��Ď��4z%�&8��$4���@�w��{l�?v�h.���p�N8�'�����o��[�M�l�����9���g8���-�y/��5	�F��hݶh�e4��Z�}�@�F[1��I���M2�����h�<�\ۧ7�e�t�]3>�IOO�ٚ:�0�-�_O�v������3���s3�����-�(�I���Ȟ�}�j��b��4���ϳ���'>�u�'>�����v�6�F�A	''$����hm�O����yh{�z��w#Q࣒bn-�s����4�����mz�s���= �k���7!��94�v��9��s����U�zm�@��>)��\��1q
t����K��j�WE�2=i���-�6;�뮪����#E#��_������{^�[l�?uڴ�zݑ�I��9����{^���Ă�ޚ���@궽�39��K��j�G#��zh��ZL��bŌ�	�� E�FF	��E�AI ���.� ���{٠^��h�w+b�Lym�NM���1}g��
��=�ՠ��ﻉD��b�)��mz����l�_�/��~�h{� �ƖG��,�3Z��#Y`2�-6�4�gq�#he�r�dɵ�I�xP'���]���|��[���@��j�:�k�-b�R���%�� |�����I�?ӺN�/�=����@꽯@/�x�o�`Ȝ�I�u^נu^ק�9�ٙ������������ժ�r$�8�n8�=��g3��_=�_= ����fa�,��A�k_w7$�}��k3Q]���vw�|�~}���'�wN���������U{^��{v2A䄀,5��U�yyչʖ�'����0m)��4��p����N&�0x�$n9�[�4_j�*������9�����r��M=&,��q��@����s���H����/_= �o�39Ď��Di�=�a&)qh{�z��i�����E��4y�-�����ȢƄ�B9�k�Z���_j��g3�����;G�g�Q���cn-�mz��l���{��w��n�]�kIX@�#%�Kl��>%Y��JGk�F�-�"́��"���D����$֡	I`K��d!�JR,J�o�.с���trB2�9�W��@�'[-4meu�lʻY	@%挰�7��	D!$�������4�����@�:Cl	$���pBp_$S��$��H�3��'GH3�fc��E����.r��{4nl�Lt�9��P�Vo���C����en��tX|͸-y�8tU<m��Հ��Xr��l��*�ǆ�:RW��v:W��1չm�ۢJ�xL�x�G6��
�6%�X�R-�2��4la�Q�oF��l�Z�w)�`"q:��D�����YD^��3�ډ�az�Q�����.M����'<sw�Yt�����Ζ��p���|Gg��U�bv�7�-Ǵę.���Ѡ����/Q�V��CVP)oYV9[��ф���<�r�v/\gX���R�Ζ6�
L�[FF��X�mH�݀�U� _g��=�4%�l;&-5��Y��LRb�"قf�d�����s{@�hZv��uq�t���U�TeP��K�0�#
B�E[qѢzפ܁mps�6�=W���8|m��6�r�]�6�R�xW%���#�-�:�k��z���n;8� e�n=��M��cF����ZV٫��;$��m\
�7R��e��cbͳ�ԜmcEv�I�7C:5T�m��!��5�$,:b֠j�݅c�',�L���\S��X@yT��Dh@k�<z^<�h[f1�ɚ傥UZ��P��s���,1�-lrnN�s�*u��r���&<��2
v`�ˬtWi�Ŏ�t��n���	I��)&Mœ{m�퇜�pcb����Ҁl٨�c��'�孪�D��'nD�}���<���B8H��Ӽ�nT�[�5t�S���n���2����3�����2����C�����<<n�v4N��Mu���(��3d�E�p��b�j��i���/!�[-Uv�v�\�ms��/M���m��V��e'Z�3P��Z���ѝ��3�
s��Ɛ�O,���%3yuU[�kx�Hm/6��rMUU�@R��26���Pc(b�uZ�*9�1ˊm�t�d�5�i�ZJXN �%�>7k����'.at::����V��ē3��m%v5&u;m+$��.����ٝ�A�ڬ�	ד(��{/Wc>f��tJmb�zwt�N�,��& �> 4��N���Sb�8���QCb�
@
'�"�h��N(�G쓹5�@Q.e"�h�P�k����]0I��E�,*4�����
��s��u���uɲ���z��@���Wn{n�r��<@s�{�qդP����']�q�n<��N�
�)�|��I���� f�!,��J]�b�h6�l�<:��q�{:1<=b�q���g� �E"v�yXѢq;+$�m��i�q��mR[v�͍�F��?����'�On��.Em���{q�����mP�afXkhK����B���i�����/�]+\
/�z�yh]��V�����fs>a����;����(�q�#�@��@�v���Zk�o�33����ʯ��NI"���9�8�/���}]�@�v������J��Ɓ䑸�z�s8���-���@궽s��~���r�^M�"�`7I8��ڴ�k�;_j�;]�@��ۓ�b�6�fV&����+��(���1{'c��E[rp3mm�ӧii|���H,�征���zk�Zk�g3���/���;o���U�K��&Wxϻ���;�$�@L"!���������{;�'׶��;1:F�Q�$�'"�;]�@�}�Og3���@�w�@����6�m��qŠv�ՠuvנv�ն�Ix�v��n^D֨�*��>�w��%�bX��k��ND�,K�k��ND�,K���6��bX�u>��*\�v8�Y�f����*�udԪ(�Ԗ���ҝF��F���̓MW�֭���r%�bX�����Kı>����Kı;��a�?DȖ%�����m9ı,Ow�����lԵ��Jt�Jt��������DX�L�b{?���ND�,K�����r%�bX������,K�N�ffre&��5�ۭ]�"X�%���}�ND�,K���6��c��D ��� %b��Ac�Q9^׹v��bX�'}���9ı,O�e����!��Wy�ӥ:S�J's��m9ı,N�]��r%�bX�����K��&D�����ND�,f�?��>S.�h��/Mzj�'}���9ı,D��]�"X�%���}�ND�,K����ND��/S߹��JgZ6c8&�#-���Ԛ����+fd&��b�VٗA��cB��m�#�0��ԥ�j�9ı,O����9ı,N���r%�bX�Ͻ�ڇ"X�%��k޻ND�,K�z�2{X�p
�t�zk�^���~�=���,K����ND�,K�׽v��bX�'���6��bX�'���Y��Fū���Jt�Jt��~���Ȗ%�bw���ӑ,Vı>�wٴ�Kı;�{�iȖ%�b~�^��
��{
l'�|�5����d/O����v��bX�'s��ٴ�Kı;�{�iȖ%�����$�)l�X�(I"�*@�!@�hEd�tJe�ed�2{H����H "�@��>z lF��;�����r%�bY��� ~����}O/P�B��g���r%�bX�����Kı;�{ٴ�Kı;�{�iȖ%�oS���Ĥb�*���B�i����04)u&�K
jh��`kݣ���	���=nI�L֬��Y��Kı;�{�iȖ%�bw>��iȖ%�bw���ӑ,K��=�fӑ,K�����][��֮ӑ,K��}�fӐı,N�^��r%�bX�{]��r%�bX�����Kı?w��ÓU�Jk�M�y�ӥ:S�:}���|�Ȗ%�b}�w�iȖ ؖ'}���9ı,N���m9ı,O�۹1����;�yz���^��~��Kı;�w�iȖ%�bw>��iȖ%���k��ND�,K�{}� ��S�>^��צ�?�^��9ı,N���m9ı,N�]��r%�bX�g���r%�bX�{�wN��<߶�����mXK��ec, aVdĹ��A��$�77l�t�C�-	��tڍ�vDac,a�P�����Ѻ�i�,;j,Bк�ƀua���us����X--���9ܕ��i"�l;�M���kk6���i�:�d�l����2#ڠ�#f��h���X�fX�d;Ws>�]�+�9�h"�&����һ[�vcf���z�Whd���I%�����|=����t�uh�B�;i�u����D�Hm+�
�������,��E���f���Kı=���ND�,K��}v��bX�'���6ʐP�"X�'�����Kı>�ٙ�hg����=:S�:S�����Ξ�,K��=�fӑ,K���]�"X�%�߽�m9�U�9"X���o���ѡ��\�Ξ�)ҝ)���{�6��bX�'}���9Ƌ�����pI��}�RA$O��׹��0�0�3I�$�>��k��ND�,K�{��r%�bX��wٴ�Kı>�wٴ�Kı>��%�o�5��SY��ND�,K�{��r%�bX's��m9ı,O���m9ı,�_K���1�s�]����s8$%j�R:�Yl$�!�E���>N_.݆��P.
/ne�:��b쒹�Jt�Jt�����9ı,O���m9ı,N�]�؜�bX�'~����Kı>�n��v�4XCd����^�z��s���0 O�>(��T6؜�b{z�.ӑ,K��{�ͧ"X�%��k��ND���2%��_���0�-k�D�O���5�O��߷��,K��w�ͧ"X�%��k޻ND�,K����ND�,K����⼹h*�t�zk�_�gB������ND�,K�����ND�,K����ND�,K�׽v��bX�'����m�hg������ҝ)ҝ>�~�ND�,K����ND�,K�׽v��bX�'s��m9ı,N�v���fm.�R�f�uւ� �m���,<]���[��f����n�I��(,	��v].�Z�'�%�b{_��iȖ%�bw��ӑ,K��w�͡Ȗ%�c����3��G1�s;r�6��a0$��\��r%�bX�����?�1ș���fӑ,K��{�6��bX�'��z�9��L�bw�)-�[ը;�>^��צ�?~=���ı,N���r%�O�xOɒH$!�4-�!R0LI"a1[$�$�FB1�l$FB#$!-I �E:�>��O�k���r%�bX��_޻ND�Jt�O����K�]Inwl�Ξ�,K�;��iȖ%�b{���ӑ,K���]�"X��ȟ����{���^��ק�����P1���ND�,K�׽v��bX�	�k��ND�,K��{6��bX�'}���9ı,Oǽ��Ɯ�.]j��!V�mq�U0F&j��j��-��%ΚRm��vk��0#u��:zt�Jt�O��}v��bX�'��{6��bX�'}���ND�,K��}v��bX�'���f�aH���|��ҝ)ҝ=�{ٴ�Kı;�w�iȖ%�b{��ӑ,K���]� 6%�c?�ϰ��Thg������ҝ)ҝ;�w�iȖ%�b{��ӑ,K���]�"X�%����ͧ"X�%����~��-���gB�|��ҝ)�Q=�w�iȖ%�bw��ӑ,K��}�fӑ,KB�,B�E�DK"�bC�0 ��r&���[ND�,K�N�ffre&�5�E-֮ӑ,K���]�"X�%��k��ٴ�ı,K��kiȖ%�b}�w�iȖ%�btϻ�+<6��7G�5ō��V��Dm]浯h�����4DiQ��P�3����9ı,N���m9ı,K�w��r%�bX�{]�ڜ�bX�'}���9ı,O��0���հ�5�f��ND�,K������bX�'��}v��bX�'}���9ı,N���{����K!z��?����߲���6��ֶ��bX�'����Kı;�{�iȖ%�bw>��iȖ%�c��ޛ��s�G1ϟ���m1"˚֮ӑ,K�;�{�iȖ%�b{>��iȖ%�b^���ӑ,K� &D����v��bX�'�_��̹�CY�����K��Kı=�{ٴ�Kİ�H�����i�%�bX��׿�ӑ,K���K��Kı<=��E FE�DB�b$P�A�A����G�	��'-�4�������u��Ц�Pف�Sv �[��ڠ��gb�+�%�@�����5�#��Έ�Ao6[l	k�%E5cRcQ(#Q�z���iʸ��v!�1�
�y��^dពAC,�=�����<��d=my��;X}f�6�Q4��ٵ��2H�i�%2�h#ʹ*�� ���C��G��`7�+9���V�MxE:
������FhK�n�u�8պ��p:�XGk���;\�w@3tjU�V���(�ާר^��b}���ͧ"X�%��뾻ND�,K��|]�"X�%����ͧ"X�t�O�>�_��X����r�:zt�X�'����9�9"X��׿���Kı?���ٴ�Kı;��}=:S�:S�ϳ���ޚ�����nӑ,K���iȖ%�b{>��iȖ%�bw=�fӑ,K���ﯝ=:S�:S�ϳ��:��p.�3iȖ%�bw>��iȖ%�b{;�fӑ,K����ӑ,K��w����Kı?w����kP��֜�k6��bX�'���m9ı,O����9ı,Og��ͧ"X�%�������#��b9��Obn(%#p��)eȐzm6X��1� ����1v�tq�:pq��Ja�r,��O���5�O����Kı=�w�6��bX�'s�{6��bX�'���m9ı,O�ߠ}�0�k�+����Mzk��}�L�r*b)��Ci�q�"X��~�m9ı,O���6��bX�'����9�2�D�;�k���@�؉A���>^��צ�?�ߏt�Kı=��iȖ%�b{��ӑ,K��}�L�r%�bX����̺���n���m9ı,Og{��r%�bX����Kı=�w�6��bX�2'�����ND�,K���]�冃 ������צ�5�����iȖ%�a�(��L�~�bX�'�w��6��bX�'���m9ķ��?Iӿ���}����,�\m��it'l]mʈ��M^"����J�1�b�a�����}��t�Jt�K����>t�Kı=�{ٴ�Kı=��a�)?DȖ%���]�"X�%�������#PF���ӥ:S�:~���iȖ%�b{��ӑ,K��u�]�"X�%�}�}5��Kı?~��m)�"�,��.�Jt�Jt��w�iȖ%�b{;�fӑ,h��^��/�p����ΆƝX`'� ��$�?J�d1]!���mC���̸�L��9�&-���t�7&�CB]��B�0̆��ݹL�RVVR[	�ޤ�ˤ��#۞�I�J/2 #$)�d!B#��d�eNB	��u�&� K�Ŀg�2k+M4#�D���+B��%	ti%�i%e%T�
�Bp3�������i���� @�.�vq7M�Rf6ĉ
$B�HI&�LHzn�a1%�t��.�L$�U�u�w�,#t; ����))Cx�"[���ZZ�SN,���c��$��./�M--JR*@ @��,#p&c[IR%%!Cm6�5�,B$�	#��+,���ak,wt2rB)�U&��)e%e��ܐ�'�]R�1q�I�X7�$�i`�^�����M�c�fp�����l4o�5��H		e2�@�$�N+�@v
|�У ��d"͠�
>Px�����O�������� ����]
A�D����m9ı,Og{��r%�bX��w�f_f�u��k!u��ND�,���?��fӑ,KĿ����ӑ,K��}�fӑ,K��u�]�"X�%��=����l�����Jt�Jt��}�>qȖ%�b{>��iȖ%�b{��ӑ,K��u�]�"X�%���w��ɶ��z჌4=�8��7�En��� �3�-�LA��b��n���ZkiȖ%�b{>��iȖ%�b{��ӑ,K��u�]�"X�%�}��=:S�:S�����c�-�ִ��m9ı,Ow]��r�r&D�?��]�"X�%����[ND�,K����ND�,K�����˚5�fk	u�]�"X�%��뾻ND�,K���ӑ,K��}�fӑ,K����ӑ,K���o�3�2�D��Ym��m9ı,Og�=�ND�,K����ND�,K�k��ND�,��F,!�su��ֽ��r%�bX��z�f�=a�MMպ5�ND�,K��{6��bX�'��}v��bX�'���m9ı,Og�=�ND�,K�s���֦�$�I�X���^���p]�u҆����8�Y-3j]�x�
1�yi�{�D�,K�����r%�bX���ٴ�Kı=�t�m9ı,Og��m��)ҝ)��ϾM6��J��W7�9ı,Og{��r%�bX�Ϻ{6��bX�'��{6��bX�'��}w����wHn��O���� �iZ�kZ�m9ı,O����r%�bX�Ͻ��r%�bX��]��r%�bX���ٴ�Kı<g�s���Ӭ4ff���m9ĳ�D����iȖ%�bw^��ND�,K���6��bX�ȟ����r%�bX�g�'�f�fh��M���Y��Kı=����Kı=��iȖ%�b{>���r%�bX�Ͻ��r%�bX�&)���t(Hш���2H� ȨO�#�.$���:�YB�Q#�������������\f��݇J<��Ck�jxn"�s�\����؄m� ��r�]�b��;u3������nӆǑ,�݂Z<�ni���0��Pp�;\%�wQm���3��m�.�J�j��QE7W!����q�y8��p���!�ΐ�%`�i��;1
��dS��q�λ"r��+�&�Cm�]M�b��q�y�3�Y����Ŏ�3t�d�46����e�9͠)q@��lR��%��4I�X�Q���:1͗!1��<���֯�ؖ%�bw>�iȖ%�b{>���r%�bX���ٰ�	�&D�,O����iȖ%�bwޔ��9��ԆkVIsY��Kı=�t�m9ı,Og}��r%�bX��]��r%�bX���ٴ�O�ʙ��[,�����5�_t�zk�^���}����bX�'��}v��c����?���ͧ"X�%����[ND�,K�~�{�*ژɸ��t��N��)��k��ND�,K���6��bX�%��=��"X�%����ͧ"X�%����M���]˒����ӥ:S�8�w�ͧ"X�%�}�OkiȖ%�b{>��iȖ%�b{�w�iȖ%�gK��h+�0��Ě�Z��;=$�.��Cu8q玪dv�s�v����F8��]kZͧ"X�%�}�OkiȖ%�b{>��iȖ%�b{�w�a����2%�bg���ND�,K������e֡�љ�Z�Z�r%�bX�Ͻ��r��"�|�
��$-�V"�b@��$fQJ̔���
4|~8�O�,N{\��9ı,Og��m9ı,K�{^t��N��N�������Qz֕vӑ,K����ӑ,K��w�ͧ"X�%�}�OkiȖ%�b{;�fӑ,K��}l�r�sF�����]�"X�
@ȟ����m9ı,K����r%�bX���ٴ�Kı=����Kı>�eg����!�Ւ\�m9ı,K�{[ND�,K��k��ٴ�ı,O����iȖ%�b{;�fӑ,K��={�D���KH2��V$�e�r1�M6+�T�\v8�v�1�7Fe��[)JB��n��OD�,K����ND�,K�k��ND�,K���6��bX�%��=��"X�%����[�[��51�5�ND�,K�k��ND�,K���6��bX�%��=��"X�%����ͧ�Jt�Jt���M���]˒���ӑ,K��w�ͧ"X�%�����iȖ<qP�@HtQ�q7���6��bX�'��}v��bX�'����2��S
�����^�z��s{���r%�bX�Ͻ��r%�bX��]��r%�`ȟ����m9ı,g�~�:�-����>^��צ��｛ND�,K�V?�߿���Kı?���ٴ�Kı=�t�m9Ρz��s��SC3`T����w7\['|qO#�8ͪƝ�n%ێ{Hנ�r��#V��9�,֛ueֳ��%�bX��׿�ӑ,K��w�ͧ"X�%�����iȖ%�b{;�fӑ,K��}l�r�sN��5%�j�9ı,Og}��r%�bX�Ϻ{6��bX�'���m9ı,O}���9�TȖ'}�a?����!��d���r%�bX���ٴ�Kı=���iȖ%�b{�w�iȖ%�b{;�fӑ,K���m�<���E�Gy�ӥ:S�:~�~ͧ"X�%���]�"X�%��｛ND�,/���?�[YZKJB�IlI�T��m%����I%)��P�h�	V���m������r%�bX�����rR��3S&jc.k6��bX�'�ﹴ�Kı=��iȖ%�b{>���r%�bX�Ͻ��r%�bX�����0�W����]�Cۣc';���s�q��<��]��K��y�x�c��6x����bX�'�����Kı=�t�m9ı,Og��m9ı,O}�si�ҝ)ҝ?���c󨸲�v��:z%�bX��t����bX�'s�{6��bX�'�ﹴ�Kı=�w�iȐ_�0I��������%��&�pI����͉ �'~��M�$O����Kı/�禮��bX�'�ӿ���iE�Wy�ӥ:S�:~����ND�,K��}v��bX�%����ӑ,K��}�fӑ,K�������n�V��}O/P�B����8m9ı,K�魧"X�%��｛ND�,K�ﹴ�Kı6u�[�|M��k��ip冢�����&�JA��i�eZ�{�1�k������� ѳ�Ll�K�ǂ��7Z���� î7g[��7fHC��Э�dR��� -��Q!�Q�I��Vs-(��j�b�m�� �ً�>��X�K[�s(d�4��'���Pk��M�a�"
��]B��n�bU�v54JM�8�r�^g8�-�<`Y��F^!��׺t�	Wyn��k F[��%%���%˨&l%R�&U�@,�CmF]ff4[
J���KvD�7���,Kľ�}5��Kı=���iȖ%�b{��ӑ,K��w�ͳӥ:S�:|�>�_-���3[��9ı,Og}��r%�bX����Kı/�����Kı/����>^��н5���~'�t�V�i�ͧ"X�%���{��9ı,K����r%��2&D����5��Kı?����y�ӥ:S�:}��4��T�b*%�j�9ĳ�H?�����"X�%����kiȖ%�b{;�fӑ,K��w�ͧ"X�%��=}�=���s��5��kiȖ%�b_}��r%�bX���ٴ�Kı=�w�iȖ%�b_w��ӑ,K���{=e�L^��\<�\ӹ�p�2sɺ�75ۍ���x��p2�i���D�Xm�SV>��bX�{^��r%�bX���ٴ�Kı/{�kiȖ%�b_}��p�N��N�~7��fm�Qx��o�=�bX�'���m9 t@~WA�q,K�~���"X�%�}��r%�bX���z�9ı,O}=o��%�0�5ff��ND�,K������bX�%���"X�)��>�����r%�bX���fӑ,K��ݶz��	`�daU�Jt�Jt��~��"X�%�����ӑ,K��w�ͧ"X�%�{��[ND�,K�S���i\��|��ҝ)ҝ?�?�v��bX�'���m9ı,N����Kı/���m9ı,O��}��M�5յ�F�i%��)H��Y�!���K�M �^�6��2Y�x�5v��bX�'���m9ı,N����Kı/���m9ı,O�׽v��bX�'s��,��Թ�L֮�fk6��bX�'{�p�r%�bX��{ƶ��bX�'�k޻ND�,K���6��bX�'���d���4Iu2���ND�,K��x�ӑ,K���{�iȖ0>~#0$`�1�L?�]2F$a	#�)H��B�QѰ'��D�L�~�ͧ"X�%����iȖ%�bx�N��
��"�}���MwId/O�����ӑ,K���{�6��bX�'{�p�r%�bX�Ͻ�6��bX�'�����a�^+m[�ON��N���;�fӑ,K��{�ND�,K���fӑ,K���{�iȖ%�bs�Þ03s@��;Z�q��\��������9�[jɭi�^�j,Ê�y�ՙ��m9ı,O��p�r%�bX�Ͻ�6��bX�'��޻ND�,K���6��bX�'��{��0�Ӛ��\֍�"X�%����3i�G"dK�����r%�bX���fӑ,K�����"(�S"X�����Y����a�/Mzk�^�O���ӑ,K��w�ͧ"X�b}���ӑ,Kľ��5��Kı>�t�U�3Gu��t��N��N��Ͼͧ"X�%����ND�,K����ӑ,K\$v���2���@�!O
��cȞ��ٴ�az����ύ�"bU����Kı=���ӑ,Kľ��5��Kı=�{ٴ�Kı=��iå:S�:O��'�Թ͎a6H��Z�`sfaQ�TYl��j7j�m�71�H���%�h(5�l�:zt�Jt�K�����D�,K����ND�,K���6��bX�'��p�r%�bX�3ӹ/�˘%1c�/Mzk�^�O����Ȗ%�b{;�fӑ,K��{�ND�,K��x�ӑı,N��~�3h�^*w�=:S�:S����iȖ%�b{���"X�%�}��kiȖ%�b{>��iȖ%�b{��}�\��L�c�2�Y��Kı=���ӑ,Kľ��5��Kı=�{ٴ�K����6��bX�'�~��X3�e�t��N��N��{ƶ��bX�'��{6��bX�'���m9ı,O��p�r%�bX�=��a|`J�Nl���.̈́/p&P�Ҧ��~�*lJ6h���ԡ�y�	�	p�`�I�h�v�f��S���4��A��55�@�%��dN~�&�U�$c�G�12�rd?/,9��l�T��6!X @�+��yu�2��1��	�)���Dk(J˻q��3�"�q��&B3sH�(�u��p%�B�$�c3��;s}ڜ#�\"�\�IX"D���H��Q��\C��`� �����C�%� 4�f�y��Y9�?I�s�d:��"CF���a�:r�˚g3��p�Rz{Y��a�/>��ߞx���06���l�P�ޒM���F��L�Y��Zk� ?�w#D��a �_�	wĸi	I��pC	���_�0��.B4̙H��ÈF,s�@��	ՁX��y�4���M��Č�8|B⒘˅����\����E�e��5�	p�4@g@�<�($H$&���l���F<������?;}��8��� ���\�C���
[�պgG8�Z�4���n��\�=��j[�U	�����*E�3I�h�4�0F���@rn5�6�K�Vkbb0��\�A�-����Dq��i����P�q6��0ld^�ɝ������6��2������h����U��O&svr���a��=�Np'Z��[��D{�PI�.�M���0�r��SDŢi�k;h�9���pj种n���\�v�\m�@l��q�y�ڹ�2P�8�Ps�7DV�Bj��ڼ"8��
2:v�V�<v��I����=�r:-�4r-:j�,.ᘋ	��Teȍ-�r�a�u]
�poZ��6�6:}H@mp5���:Q�l��M�=\�u-[���R�-��A��&�\l�;��j���� �y���9ܖ�-��̒�۞�0�	XsᘼNN��m�%|���p<�2���)��p�l���m�rR �Bչ�݇���M��ݞv�kk�Xu�!�֮Դ�v
�n��=�X��3s&NH�5I�	�UR-��s�E'��j�9�`��-*��>l鍩f����|�:��E��h��< n�5&W����쾦:����[ ڝ͓=s�9h���֍o<�ĬǱ	��Nn�y�t���=�`[�;
��q]����-�E���IB�0��Ke*���2�25u��B�K'��:#{)�RV��Hn"��B���"�/��=s�F�۰<AgK�r�u�Vs�I�GXy��s���j��-/�{u
ɘ����XF�X����ͮv譮F��9���βA
�r����WjM�Zm��xlp�U�jޛ#ul�(;	��rM]U[UJP*���dZ��[
�`G��6wgZ��*��e��l�-Av:��on������=���ST�J��K��T�ջpf����m�s��p� F���C5��F���lU��ڍ��!Y��7P��v��U^�i�y�2=ӧ�����FD��~پ�����N���@A��"B�Z�DҀu('���>U���>�cWv3�h��l�m�h�@�q�:�t��j�B��it�J�:Q�mL�Kj��OG9��E��l���mL*@{qu-�C�ݶ��(���9[u� ��b@t�ض��X{a�Z����_`�8�8�e��p�t�)]���66��v �9���H�
B�5�9D��G�M�7Q�1��hM�g[�˒����$�N�C�\.�0e�j�ٛ/#��M�30JL)եMt�*�a���b�;kj�(�}��Kı;��iȖ%�b{;�fӑ,K������1?DȖ%�}��{�yz���^����*7%snk6��bX�'���m9ı,Ow���Kı/���m9ı,Og��m9�,K��nzꚹK�Z֍fk6��bX�'��p�r%�bX��{ƶ��bX�'��{6��bX�'���m9ı,O��}�ڥ4h�S.ffh�r%�bX��{ƶ��bX�'s�{6��bX�'���m9İlO��p�r%�bX�3ӹ'�\ִ\ɗkZ5��Kı;�{ٴ�Kİ�Q������~�bX�'����iȖ%�b_}��r%�bX�������*�0�n{Tmk�NดS<�n���l��3�Mnl��Ld���Z��b��~�bX�'�����Kı>�}�iȖ%�b_}��
��2%�b}?�����צ�5���m��(��	3Z�ND�,K�w�6��PT���6&�X���m9ı,Og{��r%�bX����Kı>�l'J�W8�;�yz���^��}�[ND�,K����ND�,K��}v��bX�'��m9ı,O���|�� �i�nc�ON��N���>��iȖ%�b{��ӑ,K�����"X�%�}��kiȖ%�b|����OiԬ��s���ҝ)ҝ=�w�iȖ%�a���{���ı,K����[ND�,K����ND�-�����K��fd��e:���f�F�h�b��]F�H�a{��OB�kX]f�ӑ,K�����"X�%�}��kiȖ%�bw;�f����dK�����v��bX�'��o�_�R�Ԓ�e�˚6��bX�%���"X�%��｛ND�,K��}v��bX�'��p�r�bX�3ӸO�f
b*��>^��צ�>�ϿOqȖ%�b{��ӑ,hR$E��@�	�6dND����ӑ,KĿ���r%�bX��vn��E"�P����ҝ)��Ӊ1������y��${�ۚ���4
����,��0|�jG�^��h�ܚ_Z�
����ֶ����x"$�!y�]��t�����Fd��I����kauԜtN<1a1�8ӓ4�nM��^�W{^�����>�D
r���q$�M��^�g9��$y[�w�ۚ~�&��{S͘�))�>4��/_j�>���{8���@���@�ϭ
�8(�5$���@�����i4����D؂���w$�{or�V���Q��s4��M��������s�>�o������Z�������41`�bӛ��]�x;Z�d�t��6��KW&ƞH�4����ڴ��� �v�@�"��P��8(Ǡ^�ՠ��@/��4����ďS�G�c1��Z}}4�ܳ@꽯@�>ՠw�X�����ڎbRM �w,�:�k�/ϵh{��J��h�@��6IĔ�4�����Z��4�ܳ@��}Iu��Hlrn�C��B{������Y��2^�6�'\<���M��<]�u�Lvݶ��s;9�>3l����vp�<ogv"�	I�����9���N��^�R��8�WL��m\����6ڸ{)�,pQt����D�Q=�N�n��o;p:�y-]��܃���K�Ck�ѷYfSCE�.�f�KKRWB$���mXh瑏lK[6컫��;��4�ծ�ٲ\�(��6�FR,�j1�������M�
��CX-�pIHdI�|M��u�- ��~�Y�u^נw��*�"��&H���٠��hW����o�G�­�% �q�NI$�v��U�z��Z��4���r)cO$p�U�z��Zol��i4�t��1BC$�G�z�V�[�4��M���g339}/�JL�ԛc���҃�^ ��^8�×;s�h,buf
7�`	���fk	�ZF��ym���{ �v�@��������ŕ=x�)��W���>��Id�t$;�Ab�$T�ccC��99�*��@�����٠}ވJQ&H�R@��^�z�V��G���v�����^	)��>$��/_j��l��i4�����в��F��c�ۋ@;{f�_�I�u^נ^�ՠ���$F%�&@���b�g	n��E�͔`�8Csł�V�&&��q�)ۓrI&�_�I�u^נ^�ՠ��@����q�I��&��{^�z�V�v����G�_�īs�,���z]�zolٳI�l�F�
�~��f��s�|�e�Wֽ�T���L��R= ��h}ܯ@��^�Wݯ@��X��RX�E0nM����}k�*����l�>E�ɆGQ1�`�T���6����P��fŅ�F�J9��*%�(2��LR��}k�*����l�*��z���h%Yd|IǠU�׷��_v�@?w�{8�߻,�,q��1LQǠ��@����}k�*�k�? �V$��ĜrI�U�h�
���w��}��˜33����BN٠\TYr�8�H8G��}k�*����l�>�����Uo15P��5�Fl[q��Q�Ŵ�h�gv��S紳@Oh�� � ��D��E�[x{�7v���٠}_]��g? ���S�)�f7� Y"M����h}ܯ@��^�Wݯ@��X��RȆE0RM����}k�*����l�>�D%0���$�����
���}����4�ܳ@����A(�Ȟ8�ӏ@��נ[f�_��h]���s/,��5F�*B񴢙r ��=ԝcpn��+p���ʹt ��J8icj!n��UI��K1d���	�0b}xw�Rf�F���lK�c,��F]�8��/]��	ɩ<MX��2���Og� k���zݖ�0P1a���8P��c��v�l����Љ^l�>΅.N�'O@,�m�6�Mm6������_�wd��_Z@c�S�I�N�4���a���8�u��<�;�V&a6����Cj�f��th�-6X0[o�� �\�@�������<���>^K�z�i90NF����4���
�����7���1 �Ys��#�H�M���@���Of$w��@=�g��~RU̒(�L��
�����4�r���^�zT���o& �8��:�k���4���{�ۻo��{�h�b�*132�C��{j����Y�^��;9ӻ6��=�9d������1���r��mz]�zWmz{�	L*h2d��iL�@�{����mR+ ��R#`�;�����s1��z��^�_�Y��$}o��7n<#�'q�V��]����������u1d�nLSq�{39���= �nzh+k�*����J�`�b�'�8��ܳ@�[^�Wݯ@��@�fb����0vˆq�q=��v�2���d�nzس�ԍ0�v��vHi��D�b1䟀����
��zWmz~�Y�v��*�HHd�
��}������ܳ@�[^�z�1���Dԏ@��@/��4X��3���㿀v��rK�a.i)7{e*J�K Ja&2�0���)�Sx�S{�c�I��ECS� 0��2'+��.�#l�$RBt���e��HXB2k]�[ Q�d @��`�\�I���`�C��~��K �@���������v%�`�YHE������K���Y% 䙄!y��O7A� H�)-���B&�����d�%��Hn�҄�(P�Cd�	��L3r$TÇ�˥O�>-�+��&%֡�4m8���'P? 	����4 : �#�x�"�B����"�~DN�	��U��x ~�ou�7$����䟿}H���&��n= �w,�>VנU�k�:�k�>�D
b��Ɏ	�ۙ4���W��]����4��?gf��3(��Gt�J�fX4�fXCY��C�1QE=�������N=�������ܞ���g�^������?7�$r"dN- ��7��bA�_d�*���-}�@��U��LNL��4�ܚWmz��h�٠*ŝˑ��Г��ɠuvנZ�V�}m�����<X��$ EEmm�4����?�ܚ��K�d���@r=�ڴff.�ޟ�=��Wmzϭٌ�#����d{m	4?�� ɥ<�l��f�Z��9�R�V+u!]E_�;�zh��4���_j�>��+�A"6�H	ɠ�����f$y_y��Z{l�fs��H�1f	ƛ�4+�=�ڴ�9�����M ���h�^<Z$��	&6��*��@/m�onM�����`�oH&�2az{l�{MnI��{��v���䟀�H�����RD�D��7{Hfr;��V��:��b�T��'���PY�q��K=�	K�1cec�sk viS�BXk��:�:�m��.ߟJT��KSK��4��KX�P�2���lw�u+@K�5�Z`��\�òԌu�&�/Z9�<���Z�-e�4��H�Z\���4�oܶ76�C��h 69/lvz�ܫ��Z������Ѵ��2<�)ǐ�����N�;���M���&�B�� �M��l�[Bh!4Rʲ��\���c�t�
�(�D70LI����ɠU�^�U�z�r�]���Г��ɠU�^�U�z�onM�RU̐s� �9�k�Z��� ��&���^���D��i�0	!��������f�{��4���{)�}�V�qA"4�RD��{rh]���S@>������0�����z�ۑKt<k�	�س�	���m@\�+��sL�f=�}=����S@>��s������h��=J���V;;�>���<�;�|��������L�6٠[rh]��}��:�,�M�2G ��4�ܚ{��W�z�g��*�W#�Cs�nMs��b^��M���@�YM ��hâ�Q�	<�L�]���)�[f�^�����w�y6JƉ�R	H���ZT״��rԝc��zB�8*�	9ܺ��9�g�C.���_��[f�^���:�k�?S����02(�4�l�g9��f$��4
������fg9��X#�qA##$nF��[�Wmz{)�0��0�HB0!BA����HBI$!$�$$�#�F�~ 8)�Z�fo^��N{���}���{�Bb$J9�C��sw�z���@>�� ��ɠ~��x�$�RN6��/�S@>�� ��ɠuvנ|�ۛ1Csf��,�� G�Y����[���My���enI���B$u�X�.����h�nM������Ȫ�\�$�	�ܚonM�338�U������uv׾��3a���BNLzW��U{^���^�U�Ǡ[��+� �@r=s���rI���ܓ��t�ɴ��H�FEL7(�H!��,��k(BEJ��h�ؒ#�	T��o7�ܓ���k�I.h����= �m�{ۓ@�[^�Wֽ�����X��Ă6�T�D�),��ϡ[�8����CY�mfV�j�H�1�I���4���}k��٠w�K+M�8�X��4���}k��٠��4״x�$ �#�F��*�נv٧�3�ď[�U����݌��ě�&G�v٠��4�mz�33�}�|�/%�#�0n`�iɠ��4s��w��I=}�f����$�=U"N$���H�?~���,�k�̴�LX+k�u�u�U�W�kM�ƀoj��=m4[?!MBz[��%Y�]����%N���l-ԩ�C��d��Y�*VϤ��c���{.�@�2���ZFK1�[�b�cD����Ƚa�&݀�ϟ.�'�ǳ&�H�9�J����7Բ�R6].1+�m���Q��2��]̆R�6R��
:�Dar0.	f��L��ww�:��{\�mV4�J+��9�Z��1�t��a˶�B<њ8�����i�"y�:����U�z�m����9����M�]
��8�%�z_Z���9�o�4��&���@�N�^<m�X!�= ��� ��ɠ|�k�*�נ}��,��#&<�F�{ۓ@�vנU{^�}m���X)Zo	�&(�G2h]��^נ[f�[ۓ@;����A�0�8����<�����c,:���t��h�[*L,k"��Đ<����ǠU{^�}m�onM����,,$OnL�I�}m���s0�g������@��������9�H�^K�(9�p��4޾ɠuvנU{^�}m�r���ऊ O"�&���^�U�z��h{���%�_d�=����$�ɉD9�U�z��h��4���s9�g_�����Ls�I-[��|k�C���a�m@k�*��vH��2\49ǎH��Dԏ�}�M ��&���_s�
�Tﺱ,��<h��2F�߻����zU�z��hw�
*�D�&(�72h]��W�7 '� �V i��N(�����rh��W�D�����G��{^�^�4��&�����^w�z{�0X?C#�ے$z{l�=��}}��W�zU�z�*�@/YT��=��nV����R�݅�`�����7]
H
�z�_0��4
�k�:�k��f�\�:�)D	�$ɠU�^��{^�^�4��&����$^.���IǓi9�W���^�4��&�Wmz��
^,m�A�!�Z{l�ߺkrN߻�ܞPl`hC�A1�ߧ����bY�Ƞѓ�BI���4
�k�;_j��f��"��û[�4�f �F�TĢK��!6��f��:�+X����{W��|�U�^���V�^�=���~@__d�>��6bI����I���V�}m��ۓ@��@��y#�ێa�@>�� ��ɠuvנv�ՠ~EU%a�$��N�4��&���^���V�}m�r����"��I�@��@�}�@�[^�v��$�l�����,h��B2���!��X���	e�0��I)qO�洙���e%#il�����kK�5��3ZK���i- �f�O>�7��	��k\+�M!(�$i a`�� `���!B�DgR+hBE�	��6FB���%�	`A�.�B$ ,�C\>,�%�%���kjs���,G���1]�6h)�\vFCI��ַ���i���P��uٔ!>��[%ӎ�`�۶n�%-����Kv�=�M��g01����BT�	ă��5s����H�o�9&���X_Ŗ���k�7��H5�4��erg��7�C�����u��{��_���3fnh?]��P0�ſ$M~�BB0#4 e~�iG��L�0��.�b��+�4~
Za��4��@�E����xj;+h��l�k���akdG��.\�)K����lS=����| );��⧳���6,K6]i�f�
�e���ջ�܏#\�Km����:�CZII�Ur,#Sm
�մ�ؒ%Ҙm�#�ե���P3��x�s	`jm�xe��srW%4Ԗk��Qٗ��٤n��౻�s���exQz��R�j��Zٸ�N��n�]�J.�c,��I�!I��Ţ	usPe^��%���Q��Wq�B��R���nܹmeڋ��z�џ)'c���1����x�9{7[���$�Yج�����q�lUr�wFjЉl�b<�[b2����p+��#caPe��)������Smq�g>V�j�-j�
��R�n��*��A�J�80S�/�I�l]Mn��ˣNhh�vD8M6��t�Hø��r+s����tcm��C�g�,�f�p��)p�����F�6�RZ��d��a��[�6�&�*��zw$�ִv��9έ����Ƿq��9ā�eD�>��7��l*�6���l��e�s<�K,'��]#�;Kn
���ݤ��⪕��vy�6�GL�k)�����(5�i-��X��C3��
�ͮ&9�k.J�s�ر�|8,6�ӗ8Q���6����!��}tM��z%��-��H3Ћv���eū��ǝ*��W�R(Ƌ����\!�"Ӷ���Y��p3���ۈ�r��Gk���c<ч����:lh���m�.��X���4I��aa]�070�K1l(Lk���#��ή��l>�U�Ӱ1��[B��[{f�.a�!I鱷2(q� g2�6��;N���ݖ,v�$al��%#�5��j�zQÝƌ�]U]J���V˱m=��b��i��nյWl�97h�D���@wI�N�L�;:̈́�2L��q�"h��JT�#�.��U����t�י(CX�KVW���ԃJ�xͅ�g2�qk+�tC6��:�x��3A�Vٚ�� O(�|
�b)Ez �SC���]E�:(�EM���+�srk�1X��e4x��x�<�ܲb�VV[�N땩}��n{��!����yE�˃��0
6[u�\�݁l݉����k d:������m��c�ĳ}K��+��V%�
"�R���2�-LZ�X�#0��R�R����Zb�P� ���2�
�d�B7� t�m�m/c������w��T,	�����q:k�v9Q鼧Ō�3~��t��σ��at�w��e
LK7�h�=Yr8�c��Ħ1�KVM��bZ\��2��w�>￯�u[^�v���:��@�ޡKŎH�c��ZU��onM��������s��X�{`����dQ����&���^���V���@��KC	�pqdnd�>]����h.����&����͘�����2I���M��^�[i4�mz�ڝ.����aJȚ����Ȯ,r����ݶ���l]>��ާ�b�Lh.���ܚ˶���h�P�� p#�9q���4Ϲ�p���F0�@�O
TxjM�o�@�ݞ4�m{��f$�,�dmH��'	�u{�z���:�k�m&�q!v�A�LQ��Z���:�k�m&����b識��P����� I��� ��hWj�/�ՠw:�`(��"b"�(+��y��z�E�ڲH�&9w��F��bF�d�R8���h+k�/���g9��W�z� Q���q�s$���}��s��G����U���^ܳ}��G��y�Q�䃒h�{�rO���n'��	HH� �*%jt_���6{[�N��M��S����M�bjE�uvנ��4�l�/�ՠ~ŗ:�hS"�9q��nMً����=�OU������LǌRL��#9.6^Ncx."s��N�s�����`e�q�ɣ�5R&�<�L��l�/�S@궽 ��ɠ\G�V�F�Ǔb�M��ZU���nM �h�P��csd䄎-�����&�v�4�h��ˤ����2(�z�g��ɠ���/�ՠ�9�p��V���nIϻl�Ft�5�A��72hm�@�;V��mz{ۓ@��eq�Q��!#iH�v�����]aU�h�@.��]]-���idDĒnH9&�~v������&�v�4��0`�#x��&6�ZU�����$y[�z}�M���ز�Qbm%2,�7�U�Ǡ��=��g3����*����z���CN5&= �h^נu[^�[ۓ@�_���b�RI�U{^��mzonM �hg9�م���aA�e�TK�[���;.��ZM5p��<���l{>6�d�z�M��4�.�td]+���1F�=,�#���M������q�e�C��aKu��#}�[n���Fž-��;7&lt�����;����).5�ͥ5d�*Z���h�)A�h�6�)��q��W�B b��˸P�4���]lȎ�� �֎��X��gt�I=$�%���OP��uu� ċ,��j�
����;D<��BZ!^.������R�ZMט5#�|����{rhm�@����ubYt�<FLD�D��{ro����$���<�|��k�s31#��S��(�N<M̚}�M����k�{rh�n<Z��iH�$�*��@궽 ��&��33�_{�@�`����I�$zU����4�٠U{^��>�ˏ��$r�E\1�����:;�Z[�uPє&�l���r�X�DH�4L��nD�zm���f�U�zU��tJ6�4�Rd��f�s3����ʬ�@���@-�ɠ^/�[�yRG�U{^��mz{33=��������
^&�#�N85#�:��@-�ɠv�V�U�z~����0���zonMٙ̾��������oۻo����8J�H;��ҥC�&�iF��2v\3iG��Y����@D��[4ED�x��4�j�*��@궿s3? =��޾ǚ4dD�&91��U�zU����4�j�>�T�����o$����:��@-�ɦ�9аR�B��@*@�Y���@Q`+�k����I���Z�W:����$�mǠ���;]�@���fq_Oyh^+��ԃ#�)2hVנZ�V���ZonM �ާpjH7q������֖����;�Ҽ��Y�np�@�cO��l0��yRG�Z�V���ZonM���׸��RBG��p�@�v��fbA�_d�*���_j�-�ŉl�fD�"�@;{rhVנv�ՠv�V���@)���QD�xۙ4=��s�U��z�Zk�hw�1A�V @�b�>����I-��@��G�4dD�&I0r=�YM�ڴ�r����fs�{�L�tj$�κ���=ZB/����e�l�,�0=����ghOY�Òۧ�*�R/�_?yh��U���h�s��<L��ND�Z��f��mzz�Zk�o���ď+S��P#0�$�*����ڴ
��@>�,�;��r�� �(�rG�w�ՠUmz����fs���}j�s$���	ZVנ^ܚ]�srO�g{w$�mxI>�H�HB龇�O,�������mF�]�'�g�hi�\L�QФ)5����K���b[�:��]v��6(,v2���n��s�g	�K�(P�C�=��۵r��0є:����32]u�v�\�� i���Z�<J���
\���l��	fT�"��j���x�^�
�f��.�
b������ޢ�z2`����sq�=�
����V�l�r�]�$�t��'w{����n�h��Ćl%���`��a�]5anFRcbY���-�����
�F̂L�����@�ڴ�e4
��@��@)���F�xۙ4]�@��S@����ۓ@��G���Ȍo$�ԋ@��S@-�h׷&�k�hS�^G�5$ƣ��[l��nM�j�;���?"�u�DLj<�G&�}{rh�V�߬��[l�_���R9���5��<y"�xxg�08��v��9t�ҵ����ȴN5���0�d����vt��� ~��ɠ}��%r��,nMj�I���|A>Q^��D`�л~�]��k�o�q#�P����$�N8E!���4��ǠZ�Z~������d#fA&H7&���]�@��SC��%�{�@��3�ǒ6�cs�k�h_Z��f�}{rh���C�A�1I!6R������m�3@�{q�qX�ӺhMl������Y�Ȧ
E��٠�4�ۓ@�ڴ�ى�Ն<RN5$�m���ɠv�V�w�f�~�G\"r(�1'nM ����>�w�s� �4�x�b����y�XT��ɉI����8́�ö�w�˛7���g�Rr��Y/Y�N�wis�N{,�p��&�ָ\�o��4�?2�c���5,���n��w��5&������f ��jh�~��BF�	��O��:��@�0�J~Ҳ�T�FE�6
~ 4���Î䑙�p�4����� �M��)`B�t�X*:�B���HJt!��"��B��\��!!�JO5��J�	eVIL	}�/{�5��o9������w��IK�1��a����]�`f�j�Q��;8'�H.��$�Y"Be��n����?�4|ID�.��b�"	>:K��:����&���$�{p����?@��&~8*�;4&�ń�W�?�)Y�H@T$����D��+7,4�&�b�x!D��W��~���h�Q>6� BQ!c$T� $	2��D�dQ>D���'��!��~�������4
���xLN1@	&M�ڴ�[4�١�s��b]��M�:����"��$ZWֽ �h׷&���Z�}�I�O#Ȱ�FE�n�L�q3%�aR� 0�m3Wr(���d�R窑�1�8��٠^ܚk�{3������@��ą�!2	2A�4�ۓ@�ڴ�[4�f�/jF{�#�#s&��?yh~�h�� ����?[S�hDDC��Z߭�m�@>��4&<�9��P���N"KX��2V�@������y��rN�}��K;�kx��rM �٠^ܚ�ՠu}k�=������F �C�	��Ëuq�dF&�L�ZۥہLe�W�����v���<�$�M����b�-v���_���~@{���<�~��Dq�	�Nb�-v��s��H����{ޚ����:��K�Z�YM�"�:���������-v����R(��NI��h{8���=��b�-v������-�ِ!$�@�}��]�@�}�@���	�fs2�k��+)�&Xb�Ghج�&%�R�]H\#,C(^�&�]�B���w�;ovҁ���Z�Vh]��5�K@������0]���
f�\�n�0�Z�q(U��`DaX�pUء]�K	������w���ۍ�/@4z��V:��+���6:=1CM7&���8փù惢ں\�57n�ż�F��:�a���\�3,�^�I�N��믯��+q
�dFY�Jˣ�9	S+�[��V����el�n&7=9����=������V�U������ڞkĔDC���Zk�ZVנv��Z�տ��H�`�="ňo$�ԋ@�����ۋ@�ڴ�ڴʇlXӒ7�$�#q����k�h��h[^��W���#���N	�Z�ՠv�ՠUmz����lu��i��Qŉa��E0LK7�`���0��MP�ұ�u&����.�/�A�ܒ/�{��h[^�k�ŠZ�Z��
^(�r#'$�ȴ
���uP��� � $���"l��oeܓ����Ik�Z��,OHF̀�	$z���k�h�ՠUmz�U�#�ɓJ8�Nb�-v��ڴ
��@��-���jH���n'��h�ՠUmz��h�V����fg��n(]GZ"��= ȍ��-6�6m`�6�k�m�'u6<��m1ۅb�R/�y{�z��h�V�k�Z�C�6�nI�7�k�Z�ՠZ�V�U���z�mFH���)�Z�Z��h�����9��a�4BRP�lT����)��s7�-��hF|%ܭ	�M���-}�@-�h�E�Z�Z�����H��0r- �٠{��=�~�~��-}�@�w��q��0յ,�)�<�c�G@f���9�r�Z#m=ыqM\WBˢ�b!����}���k�h�ՠ�4��F^L��Q��Z�ՠZ�V�[l�-v�@�{[��J6���E�Z�V�[l�-v�@�ڴ�]I�Xd@�dȓ�@-�h�E�^�{w'�P#!$	dT�A�R�R0$BD��Q?�g2fr]r��B�Q��(!'"nM�h�]�@��� �٠{$��>����14֩i�e0��zk�9�ш|&��x��cn�n��&,H�O"�_�����
�k�m��33�y���*3�W<Й�A�܎-����f�k�Z�վ�s3>�
{IH��1��{���-v�@�ڴ
�k�-��!�Ԅrh�E�Z�ZW������� LOrF��k�h^נ�4]��?s3g)�8���ғ�B%��}�RϫEv{$���ak^K����mk���0ζ�Or�Ⱥ'�ŵ��wW�.��z���v��;m�j�B�6Xr ���՚@H��e%M�^8���larkL�K�wPLe�X�\�+�1�>ȯ����m���ۛ��F]g��YU��)W��WV+A�³��3)-,AL�.6�Y�N�і�p�b6�b��6f��I�w�$�!:I9oψ�L��p�b�,�^�F�v�5���w#e��hƬ!����
.[ID�m4�X9@��|��f�k�Z�ՠ}Z�"�"��	�N= �٠Z��k�h^נ��p���(bC�7&�k�Z�ՠU{^�[l�;���ڎG�E�y��-v�����f�k�ZQ��T�̊����*��@-�h�E�Z�Z�g2���:��0ь�l���֋��3Şı��u�D����bC(�T1\v�8���Z~����M�h�]�@�����yk���W�>��~�ν�&��� �Y|`�E�5�����
�k�m��T	)�GjAh�V�U�zm�@��-��lf���x�D�r-����f�k�Z�ՠ}Z�"�"��	�N= �٠Z��k�h^���R}�;.�^�"�u���w6j`ɋ��mX1��ggB�9�%P�����Dܚ��h�V�U�zm�@�+�cq�&GȤ�k�h^נ�4]��:�\r�2(21�&�U�zm�O���p�g;���,�frs9,r�@��h�w���C&H��zm�@��-�)�U{^����5(����	$�-v�@��h^נ�4�fg�|�3&���1�st�+a`��f�۔/��a��îR�G4F�Gh�um��"�����@��� �٠Z����V�$(�F��W������-�)�}ֺ'��Ȱ�H�'�[l�;]��-��U�z��@+Bqć"nM��-���ܓ�߻����}�j�P ���BUq7�G0d�h��y��ǜ��n�M��v7����m��:�k�m�k�^ O���}�1��!(��
Q)�%=�e�9[��e���j�����qgO�C�c��qHhW������/s��? ��<h�=�b�r%���܏@-�o��f$_?xZ���@꽯@���c�Q�@��	$�-v�@��h^נ�4��)�0H���9�ޞ��=�|��f�k�Z�U^=Rm�#X9�k�Z��{���'��&��}�}w$�  U�  ���  *��� *� U�� W�@ _�  *��� ����"*� *X
� ��A`�D
����EH��V� *�b�DB�`*B�"����"* *��D��D��D��E��@��D"*`* * *"*���Ă*
��D�"���"�b�� *`�� ��"��� W�� W�@ _  *� U�  ��� ��@ 
��  *��  ��� ��� _� 
���(+$�k;nJ,�Bۛ0
 ?��d��0�
} � ��rB@ �j�S�]v� ��Vt���逬�e	 
���%%��� �͘ � R�@ PV�� h��S@�4
� �ZR��  h4 j�� h��    ��2�@�h(P+�zr��N� �1��t�>�h�o70�9��e��-j�x >�ht�c�D���`�������[�f���#����{�p{�|�8=  �Q@(��5� x��kv�|4|�������ku��������Z�}�m��Q��}��y�ץ�wTzݫP-��#m{���g
�w��Ϡ �������� ��z3���1�{�'�wx��f�^v�z×G�}������@�CB�$m�P! �n3���wo�9>�������M�p��4�������a�:w����I�g�oaϣ� 8w��zn��>������ǡ����:$�C�`������8�� �E #���h �)�#�>�}��k4 /L���T�μ �tPl�K0h�R��h��);��΂��)�w)@��R�����-�JR�,��{wE(͔)ye)@Y�Cc� }�r����n��;�JP  #|���MR�`��[�#6�Ҕ��(�� ��_��tS���]5�`3n�#y�����p���p @þ���7|� �z�ݻ�\��=���w{���g�۫U��f��� y �2o{��'�4�ڔ�Pd21��U)Jz�� � fT���R   j{EiJ����d�a��U$�R�@DHCR�� ��=D������m_�u���d��}�����PU~j��TU�*(*��TU�eQW�(*��O�����%�2���i�Ȓ�g�����w7r�/��%5��$���0��o5�畓���C�_������L��%�u4����.�e1IB]%7����0ޒM�=��&�<)�.2���"ی�-u�W�˙y��ٵj�୵F"�ڢ�xQ����{�e0cLk0�kD�hc.�hd�f��>��Gd��Khfda��$�u����>t;�A~��|��!p׉-HҦ2J`XR���B���6����F�>���g��0�N5��jG.�7��(�:7��7���>xp�����s��6B#'6B��H��frG6y���&K.�|�=-�K�˳��d�lǉ��d����7�g�����B�����g<xg7�CA�Ic�u��ą�M%���i&����B����6h�rM2�P�t�6Fަ��A�+`\2�	K�e��S���
�"bE�d
š$B�(H�`E� ��$0 H	��$c�Vı�	���ѷ��K�d�5�y����jRo��BnKY�Ko����y�����7���!L���\�!
��������{�<,d�{����G3	���]�g�!+3\�yx�5_c�W�G_j���5����_o�;u�x\=�wZ�y2ѹYad1���"kO���*�wO@����kXK��j��/�r_u�|:���~|9���V��ِ�	}/�$7�&L�e���5Ǆwͅך�f�xK��7�����n�3�3�����ě0��˾rGZ��'���մֈ�o;�-���~��MM�6y6���T�$5	�i�
$X�$�$��.0i��J`A�
{�U�N��]QK~>��tX�ON��]ߓ����󭣃����W������g��J�!C,��5$�Gs�����-���CĖg�4��)����i�$"�a!/�p�y�2{��t�p��K鳇�T���C�xa����6�����Io���r�|�X�Wv:�'�}/�sV��Yw���g��8�x2��{�h�/�����Ȅ����"BFkF�[���v�u������*�ҷ�w���(*�ϋ.���쳟pE�>5��|U�(�V�;�"��D���Q��%�f�s+~{WUE+�W����u�-to��AWn�>���f�>WUΔ�nk|���/ܜi�,J��U�ԐhbhC�`�w�P���ѽ�7�o��<��[(p�rM�DX��{4l�7�
�hߔ�4�ܼy��s[�|4M����K���xyɧxn�y8z��5��]��=ۭ�,�SF�ɣY6����d�F�ߚ�@�=4x�5�h��Ѵ���O�����[L�+��M�{E:��\�z���w��t]�p�ۭx�^p�p�)��-r&��ϦOg��8!.bԑ\4�+!�)
aBL&7�������T�H��p�.��S�q����ɜ֦CA!�#$�!����0���%��7��8���#'�5l�W5�eKɉ+(᭒�䫲hݖM$��!XYIN9�$-��]�u	]�͛љ/��R��I�8��	�d"Nq�f܁rh�w,o�|�5��¤g������_q��y�Y��z{��f�=��o�L!u�z�xX>���f�s�w�X��1���)��&)�8K�\�M��21"V-d`�Yto�ɩ���4j!`X[�Ȕ����Y�0����(at{õ��)���pT:�>ǝ�����@����~�W߅]�u��}k��J���=꯰��y��+�[�;��*�޾����i0��A.&��o��=B�y7�a�v�}�ݩ�4��i4T��ed%���Ï��[e�oˉ3Q!H�.h�ih�#�J Jc
�3|���I�S9��4s�5���s<�O�ޕG۟v��/k�OjU�Ws>��|Mf�߾8���Ѕax�$�!�O%:�c;ߵ݊���^�"аO.��׵��9�zlӲ1.�,	�A�G$ѱ��4�V
A(
�0����ĀF$])Db0���p�H����0*,H� 1H����"@�h�Bdh�
6p�������������!K�7�'�����6���?��D����u1��\m�@����W'6�O|�	����0�5�فh�W��Eߝ*��R��)���N���t�>�|�[X��YnK\w������xY��P�l���3[7�=�6q�as��}��SoOM�6�����z��ث��Q[���uE.PUӧY��n@ы'�C�5�g���>��=�!�ܾG+��!7�J_�B�"��%�C���]���F�;�;���C��#�/+��|�m��IaR���1�+��`�%G2BXL���o3-��"����\���,�
�5[����S�s|��$5�^j<��2��k[%לn_��L���5����	/�SL,�%�8��og3�g�n��n<�t�1`�o>C2�u<�%����s������mM�ɦ^NK��[OA
¤"���|3g�9�{�E!�+��糜�U�=a���4K�	R �;]H��;���������k�|nk�y$���� iӢ@��0��!�6aI�����fg��OI8���A0�F(�!�6x���z���%14���L*���$=��&��g��B���K���1x�Ơ@��!\
�Fl��oA<�yxq�y�2�	#cBE��[ͯ6_\��r�|�y��)3��<�'�0������ɜ��?���%��כ��!��f�k�4�fp$�(KB3��y�S4�%�����э\R4���P�	%HP� V5�$P�R%���uI]��_~�[Ⲇح���y�K�y/�.aR����[�;�ka,ˤ�'�^r�Æq�O1��i�&�ZQ ���K�P��;�!ӻeg~��_+Wͤ��.�u5�)Uw����j[�h������
�}Yw[��ô|���[���:����sk���J����˦oo���W�[+_A�_,���	Mf�}צ{�����,i�L�Wp�,0�Ro���&����¤�!e���~ ��MH$<�c�!}B\D�a4n�p�g9���9�>y�8{�o9e�ѿtC~����9�����^x��@��HSVo�Rff�w��;%5�s������.Ƥ Da�H�2��rŅ�K�04��@��%�P�jSS6K�߼.�rlܤ��W7~gVЫ���h����Z���[�M��3Æ��tp4xx�+��T�i!I CIo��d��\��6��Qs�r�;�N�Dk�l�8�>of��N�b����P���|B��q���nn]��_5��l���fm���}�L�kgf����}�zf��\�[!5t�83[�zIRT�%V���ė��z3k��s���O	3^�א<�&g���-����<�x�$���Bo�4,�S)(ċ��@���5LAa%��H#R,]!s[%eIYR�b��V4 ċH�T����T4m�%x1�x�A��Y�=®͑��%�S�@�I��!9�|�y��g�"`T8�\tR�7	��$�"\IdI�m sM"o9��d�f��y�4I�>�!sI}����t��^4����]i)��'�y&�� ����Л7����7q�'̡Q��P�ۡ���
��/�/�|�q�K3�Y�Y�%%x��̆@��_��a�4����|&od��7㴎(P-��o33��~��ZFH�L�h�JbB�X�4�����7�{�t�v�NB�=�%L\����{�HRL"D�!X%0%1�#HP�c@�"CT�!F!����I�0��\e��T��)
��%�B��e�H�Hqw���$��#\e���%�L��}<��)o7����B�^W�߳�����AVo��ݧ�UBV����������h2��ks��t�щ��5��x3��4O���'`��k(�`�{37'j�0�ʗ��	r��x��k��}��<�L�'ԉ_��kk�!���h����F��H$!LMoZߞ�Wy��HΔ2�fQ��z��Y[�u�.ozٳA^>�$7�����P�K��ns����.���.2�$�B�f�	RbԅŀB`B$ Ā@ɚѳ�y���ٙ�w�%)t낶�|�w[02�+�ef[yv�n��J�ϝ>���#�vȷ׌�ߩ����G��X%Vt�!�$�D��
|p�H6,��Ņ��H h�4B56�ԧ�� .�g5�����<fM�ÌO{|<	`p�gO�6nsZB2�u����9�K	*�&�Cf�l�����#)�����q�V��JHF��*K�5�l.ki
��!q%1#sH��m6h��&��=��r\�t�e���B@�!I(����$�$�����̥�xH���=}��{X[�����(�}�7���C����0$t�o&m<v�)���p�5�p�W�Z�[��]���Y�wU<�w^B��YG�<��f��qV}B:;���>�d�M�Dϯ"ON�䜎��¿d/3�_�,�av��?�����I`��\�Ky}�|��a���r����u�!�6���u�������9���Y�i�{�9�!�@��ˌ�	e�</!���wt�.H&�ܲ3��hӒg�f��Y�7�w�v��d���렐5y��s�	�	B���o0
�N���}�U�ˮh�-�5��_Igqv��v��Z��fЪ���/�y����<9�K��Sz��+��g��'7	o3F��7�9��ɞ��
�Õ~�_.��gχi�}e>M���cO}㉰$MyM��"a�D#�B�w�y����e�'�����3مnT��iQ��Wc��v���tW�;*ئ�����k�ڳ(EU}W��.c$.�g٭���
`���&�,`H�tݶ?����������Ws�Uw���նm���{=�l��E����gg�k�����Ѻ/*It�Uep�xsh�AB�<��9�~��y���5�L�'.���xz�v�P��t�}����*����B���v�3����?���������Ec������eg)�}D��'�+��U��)<U��V��,�}/�>��j(��qW��ܺTW���ϣ���
6��h�/�J�۲�<��9�eI�"WO��Q���#B\6q�%g��)�r��sp$��^g���I�<0��%w��1�r$�H�ϵ���
yw�3���Γ��|�C����*�����UUUUUT�U*�UR�UUuR���8�\\�:wl�ZX�y�����e�����F�=��ڝ�
��ҥ0Xnw+�͞ݒ9�ͱ�YZ�t*����x�S��X�v횅����3֎���^��2۬TX��P�%���J�d6�E.�Ue&��}� ��	�T��]���v�
	��ElT9�uAe��v�T�J�LjwF]p�KU�upr�z����� �.iDX�˘P��b�]$��A�gb0���,���۲//>KWhB�Z���m�AT�K��*F�T�d��c�p�(�-j3��CEY`B%��n�Fж�����o�)W*ݲ��9n�ֱ��J6�;�8�����s�UNu�V^�*
�]P�<�僳seh
�]�P��^.,��j�hƦ�÷�{>���R�Jz��
��<N���ۢ�z�t;�ҭ]�r�{j�5d�[Brӱ���N�gl��y9ݰ����ur��PUT��Tq�rfv86����ÛT�
�fw �K�)\�\
�v�-WJ�j54@F���jv[j��`#a��×��Unַ�+ʹ��RN�ƶگ�K�����#e��)J��P�\.��e�� 9�Xni�
T^���V�z'��	��V�{Y�u��5�����eW-n��.��D���FQ��jg=cGr쫂�X4ڶ�[@hj��B8�@ٷs�{E�˸햨ɭ���Fѓ��m�\趮TiΕ�i�`��VТ<�p�U)�.�UM��A�'��)F����=�L��]�T���gOi ٶ�+������UA����t���Wvto]t� 5˲��P�%�UV�@e� �TA6�^١*���;*�*յ�K�׍UE�s���!J�����f�I�vEԢ��Ip-Pb�ʶ Ӗ���檥���'K芻J˺�eԶ5�U\2��mmr,T0���F�w�p��g�j
��a�����b���s*l-���r��爚��W��2��UT�ŴQ�UKɄ�O,m�]J�u�����n�bpl��]4m��5�ʀ�T@0a]3�{�k�T�y;@� h���,i�d���W@UUU�������Y@����A�����۴�PC�6x\9%VX�4�LD��T���[�3£��dO	:B�T��j��V��z�*ɵ[;��E�B�$�����*����7-��ptpÉ<�+W�K��ԅT�vP6����ܽRqKR]/PT�˱(���a:(�e�d�V�ON&�yN����M��*�Ɩ������6a(�;X"8f����`4���Gq���>�-��ML8j����"	Yc���*c�.ۉ�v�{4�Tvյ���ڥY䠪�(8��*�r����+U�*��OɭZ*�rԻ���̪������UUC+�&��v���*���`Rм�=l����S.͌O$UmV�v��c��ʡ��b���6��
�1V6���TX���*��h�M�v�����T���UU[U/-JcT\J�h�9�W�۩�쪪����UUUV*����鶭�gC�-r�Pj�*�R�uϺSl�UP�1*�]���-�e��UVV����j��� ��	V�����
5T m�·��JڋUW*�uUUR��U�UV��9�Z���wl`Uw�	d��55QJC Z�A2�Ŗ۫p��d�L�V;.vCa�ꪪ�]������j��
��.��������_����U��j�
���Y]���xV�UUWUTU]J��TU[U]T��W*�U�]Tb�!���8�z����������%n	���^ 9�����@�v֯0E@��T�
��Uav�AA��Xƥ5^�&���YY�ت�a�J�3*����,UUAWl�	m��Z�X�5�����
�T�O/J��
�~m�������-��U�n����V'�j�U'iZ�Y�U�	�X�'��4�61x��MP!N����Z�.W*.���U<�W���0t�q����j�Z�APPUULWUv9!m����c�ꥄ�V����^٪��@�@��n��U�Yʬ�	�����6�Ü�H�䢍LZ��
�@n�SU���2��gtV�&kX�����USfܪ�5:kE���L.l�v�g�Jp۵@���gn��7 5ut9[��s����j���8ĵV�q���-K�x)v��[E� ��h9����8�]�s���ǜ0e��^UF=[\�l �����u�����8ʵUUv۶�T�mQF�'(�0s�㡺�کy�&\�vܦ]!P�䣫`ㄍZK�9��\U��	����,9`�sM�Uv�˰hlJb����@EJ�BP��:o���n�����N�\c��d���ΰ��l�����qS4
n-��cF���T�(6�v�Pح� *�j��E)*��5�b79V�`P"��9B-YW)H���]HUn���`���ji䙧� �)P�;M6 ,��[��J]�:�w�ge�XA�Ѹ��{1�qU�I�KPo9익��<�.���3�˰�q��{I	�TP��5�f㭪� �cOj�<��-�MG�*�Z�v��|s�(������<�_��y��Յ^�6�`�%�L�@UWQm��;UTEmEF�`%9����Z4#�G�C]J$[����X�%� F��A ږ�V��+kt��;������Bv�	V�I���ҭ�`y��1�^ڊ(,�U�ׁ�����*�@�/��e�0��[*��[��0�`�m�*��Ԗ�îH�A�L�ʤ��w����uR��a���{n� ���j��V`�ݒ�Y��mm]�ڦ�mļ�ű��(��ֲ9ET%Y`�K�U�<������z�n�"^����n0�xˍ�0m�\ڪ݂����rY�mQ��!�5�Cv�����rE�)O8�v�kXk6T���q%|�=�:Vv�s<���v�1&��b�[*��j�8�`p��h�j� X����@&��#n��c�Zgg���TQ�%��3�٨5��+�o3�,�PUuQ�$�m�{�mUUU�H+�����^r�e��A�7X�g�����IUv�j�����Z��]��������
i�9���UڃP�Y^8 *mSh
���^��^8fUV�@UUU^�in��H�uQîԩ�ղ��8�yU٭ST l�.�*��J�1UP:��u�I;��3F�Uv�`C�*� k��5TQ[U)-��UT=���Wn�D�t�9\2�P��H���+�kR(�[�U��uJ�,��y�*��L�K�YU�9s�m�嶪��k�Uv��qK]X+e�UT���M�藦E�t@X�ǁR����w�z�{�m����-u�*���9Ł .w�m]�U��5<����=��J����k#r�@C�^�D���.����];b;�$�D�Sq��g�;\�(���w#�Ԭ�o3ت���ҵUP�������`9�汊��b�ȴ�4�qd9���x��V�
��W@v����"C�)[��� 4&p���JQ�]??<ż�=%����z(ꨠ��r]�v�A�:qO��i����)��S&7H�{PH^��LVۘ8W�t�{�g��2�X�k�V�!Z����UUT�nƩ�Dv��� VLN�UGN�Ւպ�C�z��ccj�6#d�rHM��j�@j������U������ꪪ���hrԬ�qT�UUUR���e#%UUm�����R�h)V�r�\��H���2��*�TP�UU[U*�l�ʻUHM[UWi��]K���TP��dUUT��UUU<�M[hҀ*�������UUTj��U�؜��j*��Vjv݊��U[U���LmUV�W*�_>��U�غ���ꪥP*��������V�� �j���
����j��P�|���L\�`�[+r�UK��yWfꪪ��
��T�J@�X�*����U٪�#�UUUT�R�8��J�UU �,�#%�UUi��@Y�Ҧ�gA�v�8C*�Ub�*������Z���V��m����]�����ګ���VP����%Z�������UUUUUUX��m
�V@��+)�nJ��j�8�p��U[mUV�WUUM�eڭ��h
��jU���j�ʰJ���d�Җ��f�
�T�y���~1Z��.�) 8�uWR�UUJ��U[uU:*�������j�*���۠,b]�%�<���\n�U�r���������V����lԫU�tuU'E�5TpU!5��g�2��6m6�t����YF��% ~-�/�U�R�5UUUUUU]UU]WI� WmU�����.��UAUU�ʨ*]�JUZ�R�U*�UUm'QJ��m([L���3�D��AUuJt����WT���Um�tQmV�	Y��f �(�+UW[*��mT�(Z��jڨ�A� h�tUn�H�fZ��d���a*�[#+�Ӱ����4�	���{۔�=���z�j��n��U�����hƇMmMh��1����
���u\�wUUV�vGAU]Qx�5W]N�jj-�`
U�#)��`���8�wl�T�];
�×j�M��[<�{%�Ӎ���8�붍W4��6cЂR�+;�����>�T�f����s�肣���)<B[��ђn��m	p�p��ɷ�����Sy7���]�]m	���wR�JαT]:��,�v�ul���PlUY���4�*��a�)6e�Z�ݸ�R˱g����QΪQҲ�湤'j�Z�����W+*�Y�]v͒g$�?ꂊ
�"��N#Ex!T?� ����������@�� �⩷� �"b��AP��P�!A_�/�R��:P8;G�ځ�\Q�*h�h�iUj� �""�/�+�F� �^E���{U�0"� � '�U������ x�	_���=@8#�'�������O@��]!���M��<�<E����9�p���D����Q�O�� lWM |E6�ȚG�O�򇢈�~T"�j��������O��B�D��(�z0��z���� �1=�q�H���@~S8��F>���z������	 �@�!BEB!"@���Q�H'����!D �T� �,��V�4 �mE�c���H@Z/���� z�ȏ�"z�$4�2$!0b�`�*�H@! BB
H$#		 H�	!@�d#E�_V�="���O	�C�a�a��-R-[@(�0"2BB���,HȌ�"��U�H��"A(��"�� ���� ~�~P�<��0]��
d���@��$ 2a!�4b��! x$"�b��Oh%@O�A���| 	� h�D4�#@�W�� �� ������!�)U�Z�
�1�D��2"L��֤�[�a���	q��40�f4e�f*�e�S���V�� �0��m��+0Y3��<N�d�:�l7J��7"t]d����F�v��rV�F7h�'Xf�;�nn�D���q��-1+k3) z�L�2+KeK6��G�K�m���B&��N՚R�cu(�%)�72�F�K�!.�J&�r�:nם��1c\'�&���m���T�R�lt��:Cf)4#0f<�0=TrE�CZ��yq
�����0�6nI���'//��w�o9��٥�0]�@L�[+
�ٴ*�Ӯ�]�����H��H.������P�aa�4�m-u�ҕUd�Ų���^v�'])f�C	�8� �*��Y�FSp�hz�p5��@f���-<f㚥�r�r`�u�tmVU�8dqEWnb���v��M�v��.r<\�㌄d�����6�����aʻv��honM)��4l*�������EA�\l��[�ڍH)%�$���q:��odX�GB�R�ܜNll4����|=t1����|tS�2r�W f��f��B�����oa㍣�K�l�3�,3M	���q9ۜ9c�]��N9<�vy����=p�vMݭ(�
��p�-�/�k�$;�[Č�i���⃭��p�kg@22v��T���.�Vd�5���L����-�,qK��\)���ӵ�d�Kvxp�8A�¼�Xۑx��ݒ,��
絰�iō��R*R��a�6g�Waz��i��h�G;o<HJ����Z�peT�k]
S"�M�zrmK�%[�<��	�O	k$/h�l�#����!���2����U��)K��k��:���b�&��%u�)�M�%ju�������<�m����\k�,�4�z���*ַ��3�ge0]��.���<��cv+'�L��U�9:�-�(���lʱrC�B�Hݮ(Ȳ�3G\%�m��7���Yu3Yt\�.hU���mR �P4P���|��B (�X�˓߼�nm�p��,��;���ێe�f�:+Q���Y]��s�+%P��pF�HL�8�h�u�eu㴄+&7v�pnibn�80l��rNڻmn 즁A� �Ż�b�.P�S�F�!��v-�94�#Yo:n.��5�a79�s�V���,�]qGl�\e�In a�l��Q��˔�y�U�T�mGZ�ޡ%,�d�lȀ`6FH�R	�$cq����#hNIAbqF����t��8`-��;���nW9�|�v{+ 7�y�[���ZM�Wd� ݑ��Xdp�7b%,����'V�5wn�vG�w�e`�� �엀M�d�ĭ��v���w�e`�� �엀�<{ �b�m+ui�m�XeȰ���vG�od��=U���n"X�Ԫ�P-brJ就�5R#c
Hʨ	D���Y�e�0ٻD���s��N�_��׀�<�+ � l�8���C��]Z�� 7dy��@�!����Z,��ҔX�Z�HBA��H#F,�#�(|'ʈ{��{�f�y�}vV� �i[�%i�mմ��7�e`.E���KW�� '��E�j�餕�����6\� �ݗ�H��X"Q�NӶ���;k �/ $���2�	.E�{����9�	P"KZv�X�L��a��K�VL�W"m�q�hitD5	�(�h�J�Q����������X�"�:���&Ě�>+��T;N�x�L�K�`Se��<�s�H����-+j۱75�kF��w�rO/����S��� !��
�Wj��d���2����n��5bBv��:�e���ɕ�M� l�8�T��vS��V����ɕ�M�ջ/ �B!8]1���lz����:�-�c�}��� l��Xb^�h-��쨌p�Zf
�e~���e`nE�un��	�<.�V)m$��'n���6�Y��T��O^ z{� �ɕ�R�N;I��Ӷ����l�s�IM���K���%������t��n�l� ����O�Ͼ��>���E 16�)�UWj��^��>��ʸQN�iP�6��7�e`nE�uM��dx�e�'�佗h/gu]ezzcS��0gcl:Қ��F)�q8�bdೆI��]�M��6^ vH��L��rqP����V���0��x�#�>ݙX�ȰdR�l���vS�V��������7nE�|�e��H�N�H��v�x�W*��'��K���ݗ��e�u-���&���`��{�ۓ���y����������ҕcQ�e�:�#
��݀�-��BMͻt��ݳ�J��^^q�v��p�����K�z	/�bSL�h�i@����A�vݠi	75y�\q��g8�ч��j�Mѕ��N=��i�$�tl�oE�;x�7T�q�d��^�#������x���@��v��@E�GnQX7���ey��^�iАm�#���S\6�&��aՃ�ۇ.���t�wx��C;F+;9ttbv��K��V18\��.�F�ak]��Yyzsa�zqX�+N��/O^ wdx�L��r,vBїB|Ht]&�[� ����*��"o���l���6^;�W
)��*�����+ ����:����G�w�),-&�vU�m����{'�0��� >���+ �^�*I�&�wB���l� �dx�L���+ �+�U���)��o�-b �[ǎ�+�g���qà'd8�my�-�L�"�e6�����x۳+ ����*�_ ;'� O/�i�Z`�s��>}������N����z�wt�4�9H@��%%$*憍��R$`\�e�z���؀����͛�Ny<���v]\;���I[�-��;�2������ݙX���bm+�j�0=\�*��吏 M���ٕ�vk����e]'V�t*N�[x����2��p�͏ ��o�Ꚋ�.� i�.*�W��qe;2;���]<�J�����=SĮv���M�m�ݙXf�`�c�� �vRYV���ݺ���u�vk� }6< ����̬�Uv��݉������{#«�ÕUA�9Uʕ��js��3���>��EVҲ�l�%V�x���ݙXf�`�c��.X��Al-�n�{&Vٮٱ��G�oc��;i�EN)�C\�F�@4�9����6�/�p�
��%]��MX\�+<����ݏ 7�<�+ ;(�v&�|V�� ;�{��) ��<o���vk�{�{ţ,�I:'v�� ��<{�+ �� �lx�we_%2Ӵ�;o ����6k� }��krq|�"$"HH�+��Q�o>x씒�Tݷwn��v�`5� �9ʥ�O?�'���ٕ�nܢ���ڧ�t�c@�t��v�@�N5nk[Xɂ^.B�G�q�!��-�rx���fǀ}�2���`ȣ*�V]4�*���	6<�ٕ�I{ }� IP�bj��ݤ�Yv��ٕ�I{ }6< �c�"캔�HWV�%mU�u�I{ }6< �c�>ݙX �%N�د��m`۱������$�� uU?�:ww��Y���t�3D��d��;\��ݴ���Ok�k�7nx�rK�mڍ�'4sZ����s�Ԇ��ѵ��������3��£�փ�ێ���j��v�k`2�rE���&ط����J�M��b�6�D1P��������}3�m5Z%��+H����˭������:p����8x؅�m��˻6F��Ӫms�pЌ��a�t��N�M�޷�,�N��*�e�+gZ��JK���z�e1���� ��Ql�j8+�c*��շ�vy�ݙX��`�c�'c�*�V��T����7�2�	/b��ǀlx{���[�ݺv�ݷX��`�c�	6<{�+ ��aV�ݰn�C�����ǀlx�L�KذMQ�m]��v�ӻo $���X��`f�������9�E���[tl�H2���F�j�[=��&��e0��[VQ�&�˶��X��`f����\��}���߾���m�j۳�Y�^şo
�s���������< ���ٕ�ĥ&�&�|M�m`۱������$�� ���Yi&��:�Iݫo $���fV%�X��x�N�_%2ӵJ���{�+ �{ }6< �H�UUUw��5��8�v��2f�L���̛g���j5�5dʗn{;��<�Ol���A*b����$��M� 'dx۳+ �d­U��݊��ݵ�nǞ�r�o��	��X�س��8�{޻�e]��c����<{�+��QG
�$!�*f�f��Iȗ��ulH@$	E�d$a	D�	2Y!)�w�,��2��<JA�"��ԭ�E�ǻe������|!���(8�!� f L0`�῍�]��@b0ؚ֗3\MQ��1�s`��p�bB�Hh������.��ÈNT[�r�B1��WWWa��8��8.$��'���MRf��.��N�g6�5�%2�� ���˨h���&bodV�Y6��s8K�.�W���f��"G�0��1�J���a���<����B�!�8���fa2�bܾ��n���/4l����"H[B���T<C�� "� ���H�Z �r�d�"�"���Q/� $H)�y�}�ܓ��~��$�Z�ME�I��[x�fV6�,�6^��T���x����n���M+�lm�6�,�/ >�<��6������]������vڛ�-h�ּ�2q��4�ѳz�3���fӉƐlUbn�k �n���� ����9���d�m�}��PE!,�l�H��L�v�,�v^z����o��W�2�ݔ�;�m���V�{ջ/ >�<��Ie�j۶���v۬v�,�l� �H�2�UUJ���Y�� !��%W$�*�~�� ��
*��P�;������I/ ����7oF�[�Ҷ���C���z����x�����N�F����� 'OCƦ�WY{F��L�l����̬v�,�6^ IP�*���;wn��o ����7ob�>Se�� ���U�㫫M+�t�u�M�� �I/ 'dx�̬ �K"���vSi[X�Ix;#�;�2�	��`�ZJ���:J�V�� N���̬m�X�l�kg�*%``�̕Ąp�-�̿u�K����[7N���21��q�\1cr�v�u�%�=>��<���+q�齲����Ԁ�+*�!H=���`�j4�1�;mՄ@Hu-���6SV��R4d�Vۨ�2�
k���BzS�\"��G�WC�3��y�ѷL�H'X�H�� La�HM���A�Q��4q��-)�1������!��P^��[�;�x!�o6�5�3.�'��E��.�L�*�N�\�/�VtՕF���3p�3k4d�n YRZ�ƙ�����a�&�˗�����&��/ 'dx{����v�Z�v�ݷX�p�>Qlx;#�'ve`l�U�,n�b��jـ|���vG�N���&� I.S�V0E��i��lxݙX��|����(�Tݤ'n����Mٕ�~�s����x��/y���x���\N��+% (�"l�%��9S��ǂ�a���!��k��eͳ`�ۺm��$��� $���W*�U���V {�V���M��M۶`-R<�W+9ʭ�UUW՘μ�&V&�g���${}�IVX5j��Rj�m��<�͙X��|�H�	ؓT\�M�U�v�o �ٕ�I��T� �6^�d��VYm+V�-;n���|�H�Se��2�W3��'�����U���+�M��i,���Vjғ �mX�nb��ٻE�ggWT\�|T^��5M��vl��6k� l�*�|�i�Qtڴ��5M��Mٕ�l��� $�Eʫa`�t��xݙX�p��*�S�s�\V�0�*	\a!#��*�*���Uer�x�R< ����]�%]:Ui�v�n���|���͏����`��u�؛.�M�n��T� �)���ｕ�vI�����~�}���0����b�8����d�v/u�@�#�;x�p��7m5�M_�҇|�	áRj�m������Xd�^�W�:�{� ��My'e	�)Rv6��ɕ�������߲�Q~��d�=ʤ��I$�!��e�շX����}-l�=�RD���l�V�d���T�m!��;u����x��x�̬uQ�pj�Dx�h菝����_���vӫ�i�� wdx�\�l���=��ke縑����?!{���Ő�p%��1������[@�u�;�݂�@vh�J�N�y����J��p�+o@����=Il���������|�T�z�zG�U
X9,Rڶߑ߻��[<�_���q����O;�vo�� ��.�`;��)?�c̯��=x�l����9ڪ�]���+ ���+�����n�2�"�ͷ� �{�|�?��e`=�=���\U\�����~���hO��e]'cm�z�w}� ��UWyS߿xy$�����O}��nH� �B 
 	�w����-�0��y�d03ɲ�ڶ,���*콌Wgmf:;��Ԩݩ�oT����U�H���8�އdE���LT��]=�%DC��mѥ1�Gl��r�JM[�p5��z��P=�mk�7`1{x5�C+
�f�c�K���i�Ĩl�4
�jۘ� W�c������co
�n%�������i`5G\�%�� ��8М�cíD�L���/iiy$���nD@�P$MX�-s$�%�n�����T��r���-n�WSG뻕�2Te2��VX�u �'���jz� ��?r�A������w}�\,�M��i*���ݵ=y�_��G����7��e`�eg��$z�e7˶�Z��զ� $��;�+r�-����w֧� 7kB�	��t
�����������'�߲������q)=�E=v]z�ҫe�ۻu�vI��{����Oy�M�[m�<څ%�бQH�GP��f�TT�.��vm�]ŀn���d��,����27'��v���vG�}6e`�� ��J��tZuj�E�� 7dy�o��bA0	J��'ૣHQ@�ů*�ܪ�UUU����ۯ����xȔʴ:C�L�N�m�vL��8`v�����d��S-ݵe��Xdp�>��$x�fV���@+�e����l�>�[/ �r�������X��wv��i(Ʒt�a�hI��lsϬ.�2�d��t��U�qc=��h9uyz�qu�]Wx����7fV�8`KR^ n֑ڢ�ڥm��m�ve`G�jK�	$x����)4˫�t�u�I����s�}����0B�Q U\���Uu\l�#�;$���U԰h.ݎ��v��jK�	$xݙX�� ٲ�*ʺj�Z��i��	$xݙX�� �Z�����CEZ�h�i[M01�a��n1�^Y�o�����Y�XR�Rge5`ecI�E�&���$��ԗ�H��%$%F2�ݻ��m��$�e�/ $��d��>� We6�WiU�ـvZ��I�R^��V�y��	6��|V�j�m�������<ӽٹ'�}���� ��!�Q�i/r��|m����E��*�,�d��?s���߿}����,)%�ܫ*�YA���$�qK�P��"�K6K�3Vnl:��Dձ�k´��M畆��d�ѪM��{������ʯ�{��V Hz��C��un�ӻf��z��RG����$���	#�z��I{�b2��Z�V�4m`^�� �ɕ���T���� �.y`"S-SE[�L�N��x���s�9ʿO߻X�ߟ� �^Ł�%�{� ���T�^q;�wWv۬H�~�9\�\��=�t��ߞ�ɳrM3��]���	e)���II`�Q%%H4��\���cD��$�HXF���"��$j�0"A������Ct�i�FH�k���<�Շ]���yø��D8:Y��&����$.2��Rd�	s\deĐCW\q=�4:[�3����B\%sF�LpK�'3@�q� v/��s���jBՎ�*�@���F�̞�B2�$cK	"I!�

Ƅ����#���ٽ!��2I			!�FB\����[f���9�L�a�+�[)kD�B��p ȬH0 F1��G��ʦ�fB��U m RB�XB1a�b��%bR%�b�	V�$JI	00D�#�� B��hi����&���
{�Ź���8��m���`8��\S�0�L5�e/���.�]9��e%|�'l�=�	OF�}��c4�}1��4J��R��e35!5���j������|���U`[��_��{i�Ի+ۋ`q�����X�I�N��s����A��\�=������9�#���vy��'�N��n��r�'\iZ���j��f* ���S���n�LY87Dl�9O����v��)���:fʅjg,�Z,��BH��m6<O-�!�����c+��`+g�9-� ��f��@l�\�����FZ ץ�)�h�`N��VP�ۍs��7��5�780�;E�qh�aSv�+5�gll[���J�tUb����K�@�������5�p3\��Ɏr-#��Z�Smzs�յc7l�R8�T:��E��v(���#�˷R��j�*����B�J��K01#\�ƣSR�V�%j�6���-;��xS삩�7.�˻WQ�J���ﾵ����є#X��ЊU�qm��z�qōB���C�uô+vk��mr�R�����$��;�d�8�B���w����ݑ��e짱u��Ncbj�s��e�Mz��ٖ5�\�v%����G6.6v�a2]���Ȯ�q�=���C��3�xz�v�筺(��[`�k�֤�Od����7K�"gE�Y�}��+��z<�C��٬�`g:X7Z�<��#s٢��<l@���1AUu�h�ЊH�b��ƅ8�V	��;v.�s�l�c�\�O[�˛F�Dp�Om1����tz��&�+�c]���ԥP�`��� ����Q)6I�@�\%�)cZҮ\1�Y��V�g.��f��
uۮ|vش��ܯ�a���(�Ԧf݋h�W������P��͛k�pv��d�*�K�¤��96�������m���G+8����ʳj ��Y�6`N�ͪN�Z��l�NM�%���G6�%��������s/ ���<����!y���Ը�ǌ9����Y��$��{����{V�${tɊ���x�����@�y	��`S��8{vt�
r�Y�6�h������qH"Ey+��ٜ6�]�K��d�5�b�'��Ut �P�!� � �|~���(�������J��5�̷jpX�<%�iʈ,n�esvƽOm������{.�"buq�:2�&�gvu�W,�-�#N��*�m�sp�<�Q�c���5љ����d�2�r荽c2�6���v{5[ue�c��cBہ�h �}lw���7v�m�t�f�wX�3�'l`(� ���@�b���a������<Z]�ŭ�:�1Ԏs�ò36��-��֦h�T� \����	|��1�j.�@�u,����F���jE:��X�ԉ�JA�n{`��t�#�-��)�heo�|_�, �G�}�ez�_ ���`�Z�1�iݪI�[k $�窩#g���{�~0��Y�$T=I�M��tZ����V$p���U����y�ߍ���߿_�\}����*�VE,M��Uq~���ՀH_��I��ž��� ��y�`��t���Xt��UU/{�����	$��&�%��\<3p!���	�Z��E-n�h�*��K���XF��������x,ބtta�u3w���<�L�I2�r��r��	�_�^�ߒ����-ڦ]'v��L���D� � ��Q$>��O���f�{��ٹ'����_ʹ�߿~%-�v�f]a��kF䟿~�� �ڒ��+�����^jI���$��mg�#VW	Bʹ�=�%3�{�l-�����[l��kv���GZ����Nr�?OC�ⰱ���hl 3��� ��H���x {=�.p���� ߿m3�e���!k��&TxŹ;cF�f΋[��%�v�������7�y�iKlWEݷޤ��{)�I)�}_|�[忕W��m������m���'�Y4ak�Z�e�� ��qs�KII�/��$�����$��)��U]�Ka��$�J�C���pޥ�6 �e��\U��@zޯ{�7m��~�r�g��G~���V���[�'t��I:+�~�9m���l��m��~��[~z(k��m���g��$����!m� {Ti$���Uʣvv�Ԓ����$�_l��f&��EG`�j��%�J
�nM����l�[���y�* hb�Q�pl{:O<��[iw���E������� 3���;�}��}� ɞ�`����#VW	:J���~I%$���8 d�Y���x��-jH�Z6ⰱ�m��X�Iv{��I-��%��U���� {��b�):���(Ig8�%�$����n���qs��n[�o�PĄ��"��pG�
��������~�9� ���uDW�B�m��{�\���ױ�~ ��^p ;ܷ`'X���8;����ۮX��e�5Ϙ܅��m��Ŗ�i]����w��u|<����Zj����}�/���I}�?�I$�c~�*���Kd����$o�CnH訬btnZ w2���Du�[{���������[o��k�w�4������UEE��y� �y�I%������W*��A��$�}�?�H>3ǻ,A%�J�݁�-jL�����% ��ĒK�#�䗪�˻���$�}<|P����˺(i�����bV�¯�{���{���k[����Ü���I���cL����e��e�����*�0�%�+a����N��
m�M �i����W7[��.�n4۴�Ӷ�Զ�$�	�O�Nղ����nA��i�6��[�MV�

۱xY���y�Â\��rl�Q�m���3+0ˈ3�uV�ց�@�Fo'n�P"���W���n�m�"�� ]�t ��S���ZTf�X�e�0Ͷ�V���'�wGxy�J+3	�3e���]qr��!��7p9��i���8|m�ٮ'��0{�b�cuс(�� ~������Y�����+���JA��$��^�]!�D��8Ky��ܳ�I3=�� f;�`�̼��$��x�~UJ���-RY*� 33�\�z�l{kZRC�{ל �ڛ �☢,NKhە6��^�r�3�#I.��|�][2�{II���s���ܑ�*	ѹ(� ��� ~ZI/�K/�|�����\�z�l{ ��'%�J��6Nl@�g��������LcG�]&�s5H��t��=�-uF"�e�|�=�6 �v}_|�[���Us봒����%�ޤm�,%�JK*� ;��8kKK�i|z���9uɮ���m���뜶�/�l���'�tV߿����ĻRm����{���Ē_\���{�˻�=�x�JI�9��܅V���@���`ykRu�޿�I-S�W�$�^���/Ur�C=�6 ���TV �EY� |w6�In���Kts�$��%��IvȌ]��H��ċ*�L�(�k&���ގc����쬸�
�Q~�w_{z�(0����Ux f\�� w��ǰ�3'�ֵ������ f?)��br[P��i� w���i$�����9���������{Z�֤��zF�U
�BtnZ >���8 ��m]���KZH @�x�� S�9����� �v�6 g�8>HZ1�Y��/r�\�Z��SĒR9���%4n%��_��I[����s�~����rJE,�Uv w��s�KKZ�=�����z��$�ٔ�$���&��G�6�e�����A�M��,:���m/`Jכ�H�չ�LI+�DV��Q���c�����/�HݙO�+�U��JG<��$�q�WS����������y�kZZ�h��OIH��$�Ѹ�~�W?r��������+�ZKy��~ڻ >����-)'���� }��� �#r��▩B�v��'sy�{٭v��m����[x�����־�纮��y�P��mBr���$���,I$���$��e<I%�{/ϖ�����7���oM��Wm� J�SD�jƕbpR�QID�`����_�t���O
�c�N��Y� w߿^p���q$�u�^�Uw�����K�䗂�.KA�e����ͫ�kZR@�\�ϒK��`bI/�d��U���U�����-����un۶�	���M$���\�]S޼ ��x�\�)]6��i7m`z�\^���`^�� 7dx��X�i��Uo�U�&� �I/ �9�)=��\��&�e`�r�Q[Y�9����������PP*B̖hnaq((��s�
F�Z�0�ѹ�24X��Ui���.��E���ʐ�f^ָ�5�V��B��YWϲXz5Yu��@)AU�Sd�h���YT�YC` ��	m���n�
7h��Ե�ջ��<�.Xj̅�v�D�p�.Z4�g��]7�
p�e�\nl-���u)�����YQ�d����8�X�{�=�#��/���j-���6�@������F.��R�ٵ���l�2��}�<�z�0iv�]�
��}�� ݽ� �I��s�S޽��=�<J7k�Z�,�m��;���*�={+ ���vG��ăa�=ai��n��Ӷ`�V��/��*�6{� �� �`\���:T4n�=�W8�s޼ ������U���{;��rO�~��M��殭�-ԷN����9�ql�!=��}�"�o��8�RX�"j�RT�-RX/[��ןld!���\�ć5�.���9�E���v� ;��l��>����r�� ݹ�w����m1��U��m��>ٳ�C�HT=��$=�����`��R*�X�J�Z	$���q�uA�Jm�P� 'ܞy�~��}�� n�y�s�\�7���e'HT�\�L��y��rO<�~���? �\�=�~x���X%B;�$�����l�;�ذwc�;�L�Ur���g���޻�Wv�Sb�n�����ǀz���*�t�������w��`w�ͨRXۥ�(�WGXW9tf8q�d5�mvn�"d#��Σ���'Cމฬ��ut*i������}�"�;�ؽT�Ipm�3�m��d���T�*��ܷX�r,��� ;�ޒeg��~KKZR?��?M�nJ@�
�i��d��$��~����e�l+!)HE�-���$�<$KhO��&�RHC]x�#��1d��1�呑RO�+6F��#�A.3Z�P��-eVP�R�+�aBB�1*�mD:~�|&� p��͙�MpтMBH���َ����5�t#6H<�Ѳ�.SĈD�C.�B�S+%A��&���B �A�	 ��'7�;@����x�8�iy�
$ѳa�d'1nF!8l8`8���N��l�PN�&���H0�b��X�h����H B,�B�(E+H�(�H���Hcx��)a6]��1�����-�m$H�%!H�l#=���Q=_��C�ѿ=W�4 �p���N(:���uG�b'�;�s�U�o	ܬv��%@�m��[N���X�9\�Kd��7I��$���ŀ}#�E6�;+�m��+ �W+���޿�ݹ���d�7h�a��N�erH��f�-�q��bYQ*Mq���m8��t���2�n�h�n�n�������X����+�� >d�}?~ٹ$���O�5M�pцe�x{{ n�xzI��|����r��^��/U�Tخ��v�X$���y>�f��P�"9��߿f�}��w$�zd�#��)j���ݷ�ZGz��-�uOz���,	U�q�*�w�|��n�պI*t�h��>[%��s���s���� �M�Xꪯh�z�M�mˈ�㤒��-ƞ7��a�f�ٙ�KԆ��t����w�?��vZL�,L��l�~X����&W��UU�����x�m�ح�c��wc�;�L��0	���+�Ď���MSc.�$Z�v���V�z�����~0I�}��5N��Ӥ+v+u����_����~��~��� 7v<�I��E*RQ4�$�ӫ�JـM��r��+�Us����?~��>��~��%�����Z��٬�˴*	���A�֌HP��L���k̠	P�#tX�)�.3�c�rV�Y9Ȯ�Sc\]#r�8lM@`�v�TtF�˃G�&{`��ض�d6Dns�݋=�8熓v�:��\`��وC�^&(��v �:ƥ�z�^9K��÷�]\�WG*e��]��s�@�m�c�C�6E-���&G[ۊ�&^�X��%|mǊ�-=����I�;��|c��u6Ӷ�!�d�v��Z�{fv��&JW�v�ۯΒq�$=-ݺJ�T��x����BL��7fV nԹWV��m[.�M6��&V{��:��x�{+ ;�z�H�d�c�T ��d�m�����;6ea����r���~x���+ ��Lht]�h�	����fV wv<�$���UR��z�Sǀ�ݫ��`�� ��x�ʮ�����{׀M�+d��LJ�H'B#M�
��,R��lιr�xn	K��5Hl
���)�z�Vr�c�]�o �$��>[%�ve{���'�����l���Ӥ;v]��>RK�(��@#1+����@�߿}������&V�JU�I+e��[�n̬ ݑ��W�{+�{ޛm�̘:�R�)Y\�m����]�z�����woF�T�6}X�^�Uզ�l�]
�����+ �f̬ ݑ��F�i���TV�nm(B�j�듞^��\�e��J��e�ӡ�����Ri`й� �ﯧ�vl�������;{+ ��^ƚ.ݗV�4ճ �ٕ��<�$��;#�{��$j�<�t�Vӱ�lܒ}�{��9��훕 t�1�E�1$FB�dTaC��#���D~��y�o_�����	�9LM&��t*��m��$��;#��&V���JOy����[��l&�����r,��r��������;��X[ݹv�ut�1���[���0�bG^�tCG.���[�"����T���u� KFJm��fmm��#�;��_���\�r�a?_�� ����C��t[�v14�� n����r��������� �+ ;�.Uն�L�wISV��$��;#��s��K}�e`�����:-t�h���B���rO{��ܒ{��kraED��'�߸nI�~�Y��h�	����L���W*������Vݎ� ���V�t�j��u[uC V�֐�Lܒ��p�k�u�&��[`8	���G�
�-6+i��ۯ�6{� �2��ȿr������=��V��V�+.�m��fV{�U_�\�U��߯ �߿e`�?W+����*������wl��"����I2�wc�;�̬ ��Gbc��M�J�m`z��qw��ՀO<�l���9UT��g�W�~Bt�ҷwv��M�����\���I<�uٹ'=�_M�8�� �!A"��`���4'�ؠ�e��WD�,RR���44�+��I���B��UJp�xέ��R���Gq�^�)ے��v��X1�f��)��Y�ә8���ֆ���e�aҺ!�e(����`��Ű��Wh�ގ8���n΋Zla�e3�SEP�nӞ�ƛ7.�B�Dn�n���t��E�e8�s�+��Tk�B����챬Ļf���I�5kV4HaMr�$:t�ӻ��ߞt�B�]����0��K���]�q̆��4��]3�Z9jD�$�|�� �s.��T�o�wO~��>�� �c� n�x�.�	4�Eҡ��u�}#�{��)#��� I<��fV{�UI�$���N���&��`��� ����+ �\� >�F�4�bm;6�r����� ������?�E�)���?M�?};�z��欗%�v���2���x�\0���>���txQ��X�V�W���e�*cF��3عMi>���	�Ro��҇�cl��C�ĭ�@�_�� �k� wv?�q��I�{lܒ~�~?k-��m�Z�nff����}7� bTv��I�<���>ۑg�����t�V��;�n�I� 6O<��ea���e�� ���.Uն�L�wISM��ʪ��/}Xg����r����޻���t�Z�X�8`�U��}3��O<��� ;"Q�-��ʙ.���)�a;J�`%ZkM��<Ci�-F���nm~���?!��:�˂�l��?����N�8`�j�);t�7n�� 7v<�UURFȟ����}5�=\�U${I�wI��J�˴�dO��W�0�� � �� �""	#��H�b�� �PQE=��}R���1���x{�]�����-����K��zx�������E*T�ӷI	�v����>��`�UU)'��l���>�"�>�$'P�i��V�O�ӵc6��f)hc<���F�ڛ"�IR���'I/��F4��h���&���$��;��`H�}.E�ڗ*��];�����6egꪪ�ܪ�r��ߟ� �����ݏ 7e�@Um@_۬�0����9�s�H�y�	�}��$UX�a]%{o�-$�}=�M�'�}�nI�߶nM"��EU2�\}�!��WI7E�v���X������?Ur�\���ݮ���?�����}�,�x�ktQV�C��Σ�)`�Y�Y4�oi�n�k��ep��B�@�v���wM�X�8`K�{��Ur���� ݏ�X�
���c�`Hឮr��Ď���O<�lſ�I$Ǘ��v�A�[Sm��~��7ob��s�\�Ka=��w��,�KV��]۷Cwn��p�;�̬�r,r��r�|��+�꺶�i�N�&�� �2��Ȱ���}�_M�=\қY!@`�!! y
L V0�$ B k��$a�{�#���H��8P�a�;�)irh~aqa�Fy]��ВHK$��2��U$��	�U�]��[	n]�	n�q��hJ�$��цL~�ld���F),,�%��15���[��JB̥.�' ey��IKd�%���4���4��c��-�-�YL�G���Z*��i#% Y��!!�Hib�cFkC��!$!$'�C��$��ߕU�}�U%f���k����u ���nY�wj#r6왖5�F�Y���c�#m{X���y8ރd'y��¹�Qɸ=uϓ%+��x��r!��9�N�Ӽv��DsR0�vGu������a
K�Ա�5B5�4n�p���M�C����m����y�ƛ$�:h�-�Қm;q�K��s��{1s���;M��B�R��k����l n=�oik&��y!.�����]�k��YX�hiZef����&��T0R�F˸қ����-t��-m�Gf'nt��m]-*:��9dLmdA C�P����p60��ͩ�KAB,ݖm���U�{&�S�P�&�e�ge�Z�i�&tUu\�Wl�*�v6Sd���ns�"�݋�ݐm��:@�
�cZu\!�!��s�)-�C�9:76&:M+��� �Jں�MkchMˈ-��SK(��f�i���g���i�6�m<JuiF;Ykf�5��a
�keGB��Vf��rR4�nݐt��bh�hrݴ�<�a�C;E2 �퉳ˇj�ey��S(�:�'A��v�6��F�F��&��
�NN=�)�����-ٕ#�IX�.���g;m᲎Sqd�7u��R�s�0ӝu����18�ӂ#�u�r��h�˧�9��:^��u��-(���lV�[]B���vc퓪���	r��RY��]od��B��jT�X�^\#t��a.�-��nᒁ.�,����V�� зA�Tfy��Љ�0�U�\wQUT�E;�7L�����#P֤���m)[=6���s;;pna�@��R�L��{��lQ[-`�,6)m*�����9@�c��q=d��%B���@R�l۞�s����c����8��v�-0l�(��R� ̝��&i6fw�LkI�1�)����h�R�v�kzN��ɷ��L�B�s��ݶ�MaMK�.�z�6��ix��g=�����4Ղ�kt�?�Hwt��
�S����%"��G�4�Fm��@��C���~qSB�z{	m˓����\H��rI�z9�u;
���J\xc�s׌tk�����8����̋v��7Ft7)�6+��yp��]a<�.����z�^�O>�c�T��V�v�B�CKL����@��$�6����؋q�mм�Te�"j@rTX�����J6����T���[b&��
�,��t��-�¹��ۍn�:��հ��Ƈ=���X��;�C�OR>�h�AinF�J��uH D5,d�(Ԫ@c���`��$p.�vB����s�c�V�t�n��<�����p�+����{+ ��$�b���]��6`)%��2��+ �G��r�W9UWa��U��P�1�v2�w�{����wM�X�8`)%�I1�U�j���[�Ur���V�y��>RK��9�qI=�`#��ڱP��v!�n��Ȱ��x�̬tٕ�}�J�nĩ2Չ�+���62�3��(z]�@Z�#s+FR0f�K��o�Ҫ�ee,7Wb�nұ[]W�~�wfV�l����}~��5{�e���eܹ�ՙ����=�߶o�|�$ ��Ux[3�X}~��>[%�v�ʺm�i��M6� �6e`K�a�U%�~��$�� we�(T�W���u�}#��܋ ��Us��'��}<�_-؝]$��l�>ۑ`
���I>��$'���p�;�Z�ҐHP��U`�m�a���pz:�m�X ��.�r��h�
��.o�}��� �6e`H��UW�;<�`����,���;���fV~�9I������n�ş�ʤ�#��c�t$]4!�n����}�"�/�o�s�#FH/�P���5���I��L�)[J6�Ywm��V���[��	/�X�&V�r,�"�P��Z-7v!�X�p�=\�J�������ջ/ ����iݧ@�L*�u�����TQU"hP��/m�]�k���j��F`�]��m�i�j�ղe`�"�:�e����I�� &���
�J�XS\��;#�{��H�'� �����eg��G}<�]6�ۥI+�ƛ0^��v8a����S���7�~0�*� t�۱����r�I��v���y���nOq��D����a
�$\�  ��&�ic$EB4ˈ���Y���6�3Ѩj��%) !Kk
D��0ҳ������jVФ$�@��h�ȝ��~���w�뺚(��i4˺)���ݙXdp�>[����E���7t��ʳ��j�n��Cq���պ�Ѩ:Yc�0h��dJo{��VEQ��Z���|���ݗ�n܋ �M�X�m)CV˻I���v��6^z�T�%�� �'��ˑ`R(�J���1���v�X�l��ܪ����,��׀ڗ*�v���wi�m`i�+ ��/ܮR��� &���*m'������X��,v�X�k�I6�"�!<�O�E�˚̺!�����B�C�#4V�S��ٮ��['(X��J3��ŽgO.��TϬ�f�Įlmo9Ð�2����c�Ӛ��zgr��d���4��svu2,v6XѣP�s
�׬��ٛB�g�J&�f�V�R��cqBXX��HU�#�����7n�ev�B�lq�+@��*h��K�v�r9�;e�4�Is�����{���y>2����F�9�Rs\OF.��
�u��wl���I�����&�O[H�RJ�1�k@���n܋ �Mp�UU��������}���@鱻v0�k ݹ���vG�{~�W'�v�����萚:����[�}=dp�s�ulLۑ`[�T+.į��V0�9T�&C �y`�� �Kذ	,�)CM��e�0��x�UR{<|as� �܋ 7kr���N��I	j*�,�j �.nRz��vI�^2^����p� �h����v8`i{ݹ���^�� ��������V�����^�{�3׈�D��CC��7�ܓ���]�������r����w_�Um4���m�/~�x��Xv8`B�,�"2��J�C��m`~�\��3ߖ=��0�{�0�C�Ln�m`�"�=��|9���?};��}ɉ����T�q4�[���]��V[P�E�9!�4� f�06�V�1��v�2���/b�;#�;{���	/�X������į���[Xeȳ�9ďm�,K���/b�UU�t����_�5s��sno��o��O}Ͼ�� ~�J����10�h��@�$*�l�HBHS�4
�5���n�w=���#*���i�+m`~�U)�����vG�\���, �^/Ԛm��Rwi��`B�,�Uo��>�s� ݎ�P�)�n���uw �Q;$�H��;Su�EII�4-�Q�Y�r:�������l��)���;#�;0���W>A�.y`���lJ�;�馛0	��n���� ��U$��2���R��� ����^ŀvGv8`BLT�wn�&];l��s�|9�o��`�k�0_@��bA���H|0I��#��E$[��즊`���8`��{}�>O?j^ŀ5߻�ZJ���Zt*�+am!A�O7r���P�Ƹ�,�Z�Sm��:���lJڻf���p�;R�/r���?��1ҫl���V�v8`��Xdp�'c�~�U~�*�'���4�mҤ��Wl�'���`�"�'c��&V T�q�*��(\j���=\[��,��� ݓ+�+��R�<`��E]:t!�n��'nE�z��UW���k�Oǟ� � r�\���,� UH0���#����q$��~��=�i^kfB�@�+[`ˮ��n��1�G'k������]�ϋu�T���^ˤSܔ{t�ȥ���Aa-a-�ct!61�����-c�� Fۥgqlۄ�H!^7#�w4-�7�0�4���v[J-��^[k1c��g��g����;pC%���\gn�j^��R�8]J�n�::`�+{1BTێ�g�ݭ;��[Fl
�)T�)�wt��O'�|/��[uy��6����g�����b�7s�:.E�`2{l�v�v˙��ΐ�E��n�+ �5� ��s������P�J�ݪ;�Xa���ʪH�_��m�� ݓ+?W)#�~�RE�lN�av�}�� ���O{����K7����c��M���Ȱ�2��\0?r���� ��_�ҫn�SO��v��&V�k��0	ۑ`*�¯J�ռvJ1�E����F��*�%F��g�h�e�E���0<���t�չg�7�~0��N܋ ݓ+ *l�[e&R�[f�r,��8UU����|��tNy5�y۹'}��7�����G}<����ӡ�;������ݓ+�UIo��`�����,���;n�t[k ݓ+ �6e`�"��\��W�g�� ��~��+�v��M7Xa�+ ���Us}�������&V�w�Y�b��o��Z��Yp4���7dք-%��f���__k�Ro�&�̠H-�7c0��@����0	ۑ`�eW*�A�'��z�^:����m�f;r,�\H����7��V�0�.1"�����k ݟlܓϧ�l��v�LID)k�	�OI�X���x]�xR,���R�#dT�I�_f�p�aR��Rd��B��eP�0eͷ	�K�+�&����t�p��j�S=!Wԇ#]Ba"D�����t�C}�M�xV�M�K�y�>fX�XB�sA�JMLˀ��މCF^!M��l��5u���"k�-������ F�BH���|��5���3iH�0�QL���	�Ў��I!�X���$r�:bk���pYI[�0\-�IO��%F�²�$�)�ʸDf��-Ob��L��5��-�.ac�H�$��K)*C!6��@��%��iK iD j��%X�g�q= �Db� ����(H F�`�E@0:��Q@��;}G���p۴�'���9R���*��O���X݀Ji���.��շX����\�{�k ��?�;r,vL� ��r����e*E۬�8`�k���I�e`�̭��3
�+d�r����,�	e�.ѻ]�ɽ�8y�'o0L�C�-�\�v�aJN��ـN܋ ݓ+ �6ez����� ����YJ��X�:-��nɕ��\�$o��}~��'nE��#��{+��Be4�`�{+ �;r,vL�v�����݌�۬R�?y`����&Vk��Es�"��^
!�J�	�g�xnBm���m���-�m�v�X�Xa�+ ���]��K+�&��͢�4��m�Q�Ƨ49�Z�t�ӭʁ���-��yw�ٔ��Cf����� �6e`�"�'nE���nګ�i&���;�Y�H�y��=��,vL����$������T��X���;r,?r�II�e`�{+ �lW����]���M��\^��,O{+ �M�X��UN3���Z�_��V�,l��7d��;SfV߾��rO|Ͼ��z
� ��C!!F "���E$���bX�"���1�7�]��g6�#.5k&�C��W��b�����h��X�5�=P��s�KGkhT��+�]ЋV�Y�֙+�!簩�2�İ�,3kH���q��;cp��"N��,�])����@�YZh�׫nр�
���kM�AHm�kO��Ȕ��Fb�K���M�v0ml@8�0)(8u2�Me����yĺ/�R�\�̺��w}��I�$;��|�놃Z]��{DYY��mH�����=�������'8�[?��z��l
M������?e`�� �܋��$�����r�M�]��:u�vG{r/UW�$����Oe`-mJi؛c��m� �܋ ݓ+s�Io��}�� ���1>;��	JK�Xa�+ ��Ȱ�*S�i�h�$��0�fV�r,v�X�p�>쩔6[��&I�$��Z�^@w1՗w�m�-3�a
���rl����l �R�]��;.E�N܋ ݎ�9ʪ�����;��x_ӥB):vݵ�N���W{�r�� ���X,$�'ʞ���}0�I��v\� ��R����E��t6�v8`�̬;T��"�'c��Cf&	Ym�+�N��[�{��7��,v8`�� �l���I��hC�`�"�=�UU{}�>O?a�+ ��(	cbE	;,���/k� F�_�!s�n&��kU�[�r�UqՒլf�*�n�US������8`�̬lp�:�VD�*m;t�� �2�#�ٕ�N�v8`d�N���E��j�a�+rO��_M�@4	B>�k_{�}6�p�
�QTt� ��H�u�M��p�&���-�=�`��%t�P�WN�l�'c��s�\����7��V�0�֠�.ջ�E�V�;�ͣ�c��*1�0{th�'=�ٻ�mR��Ђ�E����`�� �$��;#�� �0�eګ�v�ؚ�nـve`�� �0�ឮRGT���;t+�4Sn����lp�7c��I���E���*���v�0	�� ݎa&���Q� �V�j�"��$�!al����-��-%���{|�y7$���ga5�SZ�֭]Z�`�� �$��;#�68`�t�������ڰFǵ@e���H�h�Yf%fa�K �)9b�n�Ǌz��J�v�Wl���e`�ذ	�� �c� Wb��][����$+u�un��&� �dxa&VNs��*�����(��զ��� ;�l����:���	�JpJ�m[J�Xݑ���XV�xJk�`��e*ʶ�V��ve`[%�nE��|�\�UK�����:���JW���<th�S:�����eCY���|p�G��ݕ`Q�bxM�u�;���J]�� �7n��"�t-��ݜBٴqo+�ӻ����q��N�J���kvzె��cX�4Œ�D���4Ʀbz"�5�y'ml699�N�u�uC�^F�@Q��N��a��m�^ICJ)	��Sqf�R�B�GKfԳ��I:_4+����VĤ2���:h71����Y�pD$��m-�&�gmR�[V軴4Sn��6�Xݑ���X�څ�-6�զݶ�	�"�� �$��;�"�UwZ_}�OAl�j�i�o�{����Xv�Xۑ`쨆�n�%i;J���=U��/|{ݬ�~��&܋ ;�< ���l(���n��Ȱ	�� ;�<��+ �Z�0%rTºQ5m�BISapG({v):�[w;g�e!���T����u�cqt�m`c� wdxa&Vղ^6�N	��[I�`vG�s�]��9�s��Wy_|c'r��r,lp�>�ȭU��n�ؚ�m���+ �܋W+��.�<�`���mȭU�[����L��;�"�&� ����L� �mB�t�E%j�n�X������;�"�=ʮ�S�b7ڎ�x{:ڍ��r&1�\���sF�6���:s,k���c��瑷��y��L��r,H���Ce�uh��Tշ�vE2��Ȱ	#� wdy|H+�E(���(�����X�d�H�s�UAEU�x\��q�a �Ip@(�@:Qׅ��}�'� �0�e��IRt��w��UR���0g��ȦVղ^%���v�[I�`vG�vD�ul��I0ˀ%u8�T�}�v<�r�k����΄pa�85�����[{�lvU��uwbj���ȦVղ^$p�� �n)e[un�]հ�5n��ȳ��W�Wg��� '�� �eg���H'���`��V��n�{�~0�#�;"�Xv�X�ivTE1մ�Uujـ����;}��ܑ5!	���"b�đ�#!$(ZL=T]
T�����HM�U*�'nĭ4�5m��L��d�H����R�VڲT`<��'���:�N6Ȑ,̰�	`!��V�i��m4諶���j�J�`[%�G ���ȦV6 s�J�����$�ݑ��L��r,J')Zj���m�ݑ��L��r,H�}]����1իV��꥾=� �~��&�r���<���e[un�]հ��`ۑ`c� wdxa0Uur�|:���̹�&�Q��ɼ�="B!#2��	J�,k(JBBF, -)V�� HHS(U�R}Y`B��~`R�!�.fP������X�"�
sR�j�����6�p%ō1!p���(Jc.2�Ͱ�ĺ������4�v��޷��paX��3^k��.˄�%R��&=l���$�i���wIy<]z��{���o�5�2�&1����6���cm ߾y�����It6��-)�q��[���M\������@�IRQe�H�V4�aH��hP�a�B�5��I�ri�{�	4a�g�7w�bD�����-o��`@!$�EB?2�$���C<<��`\a	"1���ʤ�H�Jh-b���f�<u#!$d��� !"!		�K6`�1փ_X�8p�g�M�9�ނ]��hM�J(c�RP���ͧ�#<Cs���.�JM��k+,"CA).�ٔv���r\3鬗Â���-�"��ѫ�\e�\�� \5���K��(��8��|�>~�����6�Ac����pM=���B�v9���ґ�hF�C$�4R���\�Bd����\`6�ΰ�d��t�Kv�B$���Upr�ۅ���:��{6a�y�gq�1��L��ёS[�%�8�l�Q�4n��4���НF[0�%�(��s��v2m�ԁڔb�姴�I�6���!6�m�N��u�}�A����v��/���+�_'؟]��XA.ԔJ�G6�n� ���
n@�.��m]S�#��Di�����
�e-�m�8x`�[�rW6l#�0n�Ͳu4���nt5��Z� vmAQIO\"]��N0��n�e��y�q�6�`���U�)���lp�$^�g� �&*bs��HM=N��vyq�jW���w;"s��7TX1#���[�� PmK��P[�q.�e�V��t�tq��9nhu2s�:��1]2�J���]
 ٘���ř�a����</`�U�k&X�Zxݭ�ɰ��>ZIb����`µv��Ǻ"�[N&'#$��J(�[JRx����W\tB�o1�M�v�A�+�����B�q6��`W��K��ѴH�!I���*�]0�˹u)���m�q�j� Y`3j!vY�p�Ż2!�]�p��w9#XKDv܄e �v�:˼��F�,�7%�n�Rx�;=��-��M�T6��:�E��kk�3a�˭�<��c��ݠ �7L�)j�ևq�ca��X��,�klq�S�<jKPz�>������$=:*l��"����=�Bjy�M��r�^8:�TBq���艺�5R�,ݩ#�ۇ�95�W+$���n9��.g.�s�Ib�h�g'e���袇AKj@U���P(��Imќ�9��;�Y�����f칵�� �5�ܚ��W@I�R��ەuO�`��[Xݶu��
��ܧ�d8��3fu��pp�6x;v��m'P��lt',�S���y����:6n���.�ֆ�t"K�)���j1ƛg~�������ۻ�CHT� ��M����W���?
TBH*��Q��x pOP�� ߿���ιn�O-��B�ƥ�!.���2�b3F�jE��u�ё�z[�7�,bϋͧm���wa��͚�A�t�a&�D)-1�T�Hm[�`Msi,p]\p���mn���[Mn�dz�y�B44��:5ka�J�cn�؄��3M��*ֶؕ�n��!]6p7m؀��"�ŷn�P�0���^��J��f��3LjR�.���N�I'nfO#����Kl�Ų�YtS�NG�lɩz�\�;�Unn"���Z����䔥��7u� ;�<������6_���x�Hc�i�ˤ��ݑ��p�;�"�&� ��U*�'n�V�5m��p�;�"�&� ����R��:����0���	�� ;�<��I�`���V�Ш�wi��&� ����L���d�m��N'�����B�MH�n�S���pwi��^a�#����L�n�M�
��FA��[I�`vG�ve`[%�c��v�WK�ZL�m���l؀@�"�֥���nI�����#�>ۊYcl�j�;u�ul��M�ݑ���X��X�ݕiݦ��XJl�`͏ �$��;�"�>R t���v��+f wdx��ǽ�|���68`*�άjXE*��#qKQM���Ԕ��8l�m棞R:R�X�F��g����&h�5m���Xv�X������x[�{Ԫ�t�
�bB�Xv�X����I��M�&Yj��Qt��68`vG���PUr����T� 7���훒s���'ޓ���5n��eT�=�=�t����z��ı,O�O߸m9ı,O~�{v��bX��?w�?M�"X�%�������W3-��5�kiȖ%�b{����r%�bX�����9ı,N���m9ı,K���bX�'���u���,all���H�e�WGKb�Dc0��F�-�3hM�CQS[Q��,K���w�iȖ%�bw��iȖ%�b_~�u��Kı=��xo�å:S�:_ޟ�\9I�uW-�r%�bX��]��r��DȖ%���kiȖ%�b}�~��iȖ%�b{��۴�Kı<��a�h�3.�j�56��bX�%���[ND�,K����ӑ,!��>�~�ND�,K�o��r%�bX�ߺS�h��L�Y�SW5��"X�%��g{�iȖ%�b{��۴�Kı;��۴�K����@+�"�Ȟy�w[ND�,K�{ggI�h�$)�l��iȖ%�b{��۴�Kı;��۴�Kı/�w��r%�bX��w�<���N��N���m��\���-�+Oi��C['<d�MY5]`�lK2ǀHr�5��]+�PѦ[�O�Jt�Jt���iȖ%�b_~�u��Kı=;���r%�bX����m9ı,O�'^�ۗWLԚ.kWiȖ%�b_~�u��Kı=;���r%�bX����m9ı,O��{v�����,OO�O�0�&���L��ֶ��bX�'��߸m9ı,Os��m9ı,O��{v��bX�%���[ND�,K���S9즃3Ο��N���뽻ND�,K��ݧ"X�%�~���ӑ,K�2'ߧ��ND���N���=�C8Ȧ�֫����҉bX��]��r%�bX���m9ı,O{;�ND�,K�뽻ND�Jt�Oӻ��8�e����R�!s�Sp�:�l�6#p[��Wk�l�ݔ���b��,�A��Ѧ&�`�(4U]��ZE�Mr�a8�qq֨%k��d�j[�:�j�U#�� �m�D9�%����qd&l���fi�'�m�.E[y�ssQm�
\��=W#S��2\@�kֲ'dB8�rZ�7�@Ԍ&v*��W��V�6!�̼��=q���[�������sm�}�#ywZ�݈�H1ȓM�D���W:�X�ۥ�ez��1����\�1��j��ı,K����m9ı,O{;�ND�,K�뽻ND�,K�k��ND�,K��K�3E�D�h���kiȖ%�b{����r%�bX�����9ı,N����9ı,K���bX�%=��L3F�!MKe�ND�,Kߵ�ݧ"X�%�ߵ�ݧ"X�%�}���ӑ,K������Kı;�i;�ܷN�,�j�֮ӑ,K����nӑ,Kľ���iȖ%�b{����r%�bX�����9ı,N�N�幒�ᩚ�R�ӑ,KĿ}��iȖ%�bxw���r%�bX��{��r%�bX�{��6��bX�'�>��a��#X�679p�r,�Z8җH�k��0�h�1��bs��/�fؤ;U~x�%�bX�����ӑ,K��>�siȖ%�b}����r%�bX�߻�o�å:S�:~����A��fӑ,K��>�si�iS�4
AV$�:���GOb{�׽��iȖ%�by����r%�bX�O{�y��ҝ)ҝ/�O��uȦ���]kY��Kı>���m9ı,O~�{v��c��DȞ����ӑ,K��;��m9ı,O3���&���2�殍f�6��bX�'�k��ND�,Kÿw�ӑ,K��>�siȖ%�b}����r%�bX�ߺ^�tf�]Y�][��ND�,Kÿw�ӑ,K���w�iȖ%�b}����Kı=�]��r%�bX�{Ӽ&�3F����sv=fC�����On\ón4b��7&ks.H�Vi�c �%��y���ı,O~�{v��bX�'���ND�,Kߵ�ݧ"X�%��߻�iȔ�N����l�|���4i�����ı,O���6��bX�'�k��ND�,Kÿw�ӑ,K��;��ӑ��N����=���n��J�Ο,K���w�iȖ%�bxw���r%�A�����@�:*0��"yY�߳iȖ%�b~����r%�bX���	�E�j[���Z�ND�,Kÿw�ND�,K��{�ND�,K�~��"X�%����nӑ,K�����TX�k�\���ҝ)ҝ>�����Kı>����r%�bX�}���9ı,O��m9ı,O{�_aO�Z@��YoX���&�]��%'9�vWEn(�-Ōi֋�ݰ���i՞'���Z�'�,K������Kı>�]��r%�bX�v}�m9ı,Os��m9ı,O3��;�m3S-��]�Ѵ�Kı>����r�$��߻��A=�w�hH��������ҝ)�����l1�0s
;'�>D�,Kÿw�ND�,K�뽻ND�,K�~��"X�%����fӑ,Kħ�/��34h��ԥ���"X�%��u�ݧ"X�%���w�ӑ,K����iȖ%���Ρ�Dћ�ӑ,K���p��a��M�5���Kı>����r%�bX�}��m9ı,O��ND�,K�뽻ND�,K�u{f[ۗ5��ʶE0ZU, \����ggm#�n6�GD�&��#=��r�c@�f��d��å8�,O���6��bX�'�~��"X�%��u�݇�Ry"X�'~��O�Jt�Jt�?z��eV��t�Kı<;�xm9ı,O{���9ı,O���6��bX�'�w}�gå:S�:~����Q��� ��x��bX�'��{v��bX�'���ND�,K﻾ͧ"X�%��{�Ο��N��}���V�hٝEsiȖ%�b{�{�iȖ%�b{�wٴ�Kı=��xm9ı,Os������N��N���맩��[��f��"X�%����fӑ,K��ӽ��Kı=ϻ��r%�bX�����r%�bX�/MBK~̙�VjR]�c��m���'c���0�ԫG	��(�LMI�=d��ݴ�\�\"����*����q��v�3M�wHI�d�.���cs�nN���F�Bn=�qW2s�9��Cu�a.
�IŇ-s�pb^5΃�#����]�#�um�<V�+\����k0���au��C���&0錚��7K�ڰ��c���v��~]:]��%��2	���u�NLg^o\	���蓮ڒڗAc���b-�H�FU����?�}:S�:S�����yӑ,K��>�siȖ%�b}�{�a�Ry"X�'����iȖ%�bS�׷�&�	!ufh�r%�bX����m9ı,O���6��bX�'�w}�ND�,K�{;�iȟ���,Ow�×n��I4j�ֳiȖ%�bw���6��bX�'�w}�ND���2&D�����"X�%��w���r%�N����{Ǘٍ+R��'�>)҉b{�wٴ�Kı=���6��bX�'��{�ND�,K�{�ͧ"X��N�����>R�]���Ο��D�=���6��bX�'��{�ND�,K�{�ͧ"X�%����fӑ,Jt�O��-��a*�F;iN��3i1�4��&�ܹ�[qv*��^���n�k�2jMY�jm9ı,Os��6��bX�'}�}�ND�,Kߵ�ݧ"X�%��g���r%�bX��ϻ��.�֦���kZͧ"X�%��~�fӐ�)a�^)T<�Ȗ'��{v��bX�'����ӑ,K��>�siȟ�2�D�=�߮�u�F��c��å:S�:~�����å�bX�v}�ND�,K���ͧ"X�%��~�fӑ,Kľ�ӥ�Z�em��<���N��c������yӑ,K��;��m9ı,N���6��bX�'�w}�ND�,K�v�{$�4i�5-�4m9ı,Os��6��bX�'}�}�ND�,Kߵ�ݧ"X�%��g���r%�bX��h釵c�ٛ���\;\]���ԄZX�TH��m-�	A�����������)��BS��D�,K���ͧ"X�%����nӑ,K����m9ı,O~�{w��ҝ)ҝ=�x��h5*	ry�"X�%����nӑ,K����m9ı,O~�{v��bX�'}�}�ND�,K�ӽye����jᆮ�v��bX�'��o�iȖ%�b{��۴�K�����+�$���Kמ.�'R�� f�C�H���	!"�5�U�$�Bu�wyސ�ŬHU��t���	uL5�$ef���x�Na#�s<ֲ���.�\M��t�a��9$!�e�Ȗ�cH1e��ۮ�B�Xs���R�A!���0p B��pnBF	B0��,(T��(B1��!!AwCq�<۪j��ٶ$	�<g�f`K	����"oP�d.l&��D�S4�o-� Z��J%�L�*K1�0(Bb"/��(&�|T�H�M����U�� `��x/N�ȟo[��9ı,N�_v�9ı�����{�4��F��t�t�K���w�iȖ%�bw�w�iȖ%�b{��۴�Kı=���6��bS�:~��������������N�%�ߵ�ݧ"X�%����nӑ,K���wٴ�Kı=ϻ��r%����HE*tTө�����;�����3g�'�@92Nӎ�93b5�F��F��eپt�t�Jt�O��}�t�t�,Kӽ�fӑ,K��>�sa�'�2%�bw����9ı,K�鱙�fsLۛ�O�Jt�Jt�=�}�NC���,O���fӑ,K��u���r%�bX�����9ı)�Ͼ�o�i�!�%�SΟ��N,Os��6��bX�'~�{v��bX�'�k��ND�,K���iȖ%�by߻p�e��fM�u��r%�bX�����r%�bX�����9ı,O�>�fӑ,KH~A��� �XXS�N�;�N�_�fӑ)ҝ)����R�6�R�9��å�bX�����9ı,? G��y�m<�bX�'��߳iȖ%�bw;�sΟ��N�����-��V���Eu`��1/b0�;up�Y(PM����,�뮬fy���Y�V���ҝ)ҝ?z~���9ı,Os��6��bX�'s�w6��bX�'�k��ND�,K�u�슚jK��5<���N��N�w�}�NC�1ș�����6��bX�'����iȖ%�b}���6���ʙ:S���}�����j��s����N�K�~���r%�bX�����9���"dN�����Kı>����N)ҝ)��{���e�FҮcWyӑ,K���w�iȖ%�b}���6��bX�'��{�ND�,K�߻�gå:S�:_����nb�3�a��'"X�%��g���r%�bX��{��r%�bX����r%�bX�}���9ı,M��_
�`�H��# ?�����~�j�f��ۡ�գ�O(��ۆ��P�݃�n�r���6���4�K���]�����]���yϞ^մ��X��9�6���"���{�7���*6��kq=�V��eŀ�f:"U�e��u!T�.��0t�����)�t�P��9M��W"���b�lem�9k��FӰ�m�	`1�k�۠�(�j��J���SCU�cn��wI�ߺ__>	���d�������z�wQ��&ul�e�Q��%z�$�j�@	bZU<��ҝ)���g~�fӑ,K��u�nӑ,K���w�iȖ%�b}���6��bX������K�B�c@�Wy��ҝ)ŉ���ݧ"X�%����nӑ,K�����m9ı,Os��m9ĳ�:{�{)��q��1\�:|:S����w�iȖ%�b}���6��bX�'���6��bX�'{��v��bS�:O��O�Y�V�f��Ο��g�D��;�w��ӑ,K��;��m9ı,N�_v�9ı,O���6�:S�:S�߯��T��t�ͅO:r%�bX��{��r%�bX����r%�bX�}��m9ı,O�>�f���N��N�{����eb�iL��&����DL��kP��bu�	ӛ���"F��Xх��å:S�:{��۴�Kı>����r%�bX�v}�͇�I�L�bX�g�߳iȖ%�c>���o�XE�\�[�O�Jt�J'�w}�NB
A�� �u��n%��O�ٴ�Kı>�]��r%�bX����r%�bX�ߺ^乣Z��4Gd�å:S�:~��秝>,K�����iȖ%�bw���iȖ%�b}�wٴ�Kı)�oפ.Ԅ3P��Z�ND�,���������r%�bX��k��ӑ,K����iȖ%�b}���6��bX�'�}ۅ���9��F����r%�bX����r%�bX�{���9ı,O�>�fӑ,K��;�siȖ%�b\�; �]U�r5U���PX��z�0h��k�����x�ݱ�q��Ơ�k��Kı>�]��r%�bX�v}�ͧ"X�%��w����șı?~�]�"X�%���[˗
]d֮�M]j�9ı,O�>�fӐ���G"dK��fӑ,K���]�v��bX�'�k��ND� �L�b}������遛
�t�t�Jt�O��fӑ,K��u�nӑ,o�"�IBBbF���'Qj&�g����9ı,O?N���r%�N�������.��T����å:Y�H�����r%�bX��_�]�"X�%��g���r%�bX��_v�9N��N���v�,0���Yvo�>	bX�'�뽻ND�,K�Ϸٴ�Kı=���r%�bX����r%�bX���Gl�?CWY3)tf�s�v'�����=Yy˲9�����Ĝug��B�g�1A�c��ߝ?���N�������iȖ%�b{�}۴�Kı;�}۴�Kı>�]��r%�bX�����a@�I�*�t�t�Jt�O���ݧ!�Q�DȖ'�����Kı;��~�ND�,K�o�iȟ�2�D�=�\��I�nM�sY��Kı;�]�v��bX�'�뽻ND�,K�o�iȖ%�b{�����Jt�Jt��{}��6�am�W7Ο�%����=��~�ND�,K����ӑ,K��>����K���� ��)KIJ-�b��J�0��.I*!�`0SJoȗ<�o�>)ҝ)����m����VhջND�,K���ND�,Kߵ�nӑ,K�����iȖ%�b}�w��O�Jt�Jt�������fq3 ����-3iJ�e&��ly������V��eHan�5��k��9�:)ҝ)������Kı>���r%�bX�{��m9ı,O��xm9ı,N�o�z�Ҳ�2վt�t�Jt�O޿v�9ı,O���6��bX�'���6��bX�'��ݻND�,K���V�m�.�+��O�Jt�Jt�����r%�bX�����K�C"dO�k��ӑ,K���]�v��bYҝ/��e�˘��Qk�y��ҝ,K���6��bX�'��ݻND�,K��ݻND�,�̉߷���r%�bX���;���Z�uL�捧"X�%��u�nӑ,K��߷��i�Kı;��~�ND�,K���ND�,K��� �,��Ą!�"E���?~$��,3�
M�t3�l�� ja�e�E�Yc"���)��6�2�dxc�ږVj��ͬ�i��&��A��Xqj��u��3tn�&({ �}���ɛ�y�a�` zT�=�n��.�3p�y.M�����hG$-!��nFY�{u�6�5vc���IT��Hb(}�]��E�cs��1q/��ݫ`h������՗RN��'vofib�f��c�:˃��[Y��,Z��v�b$�)!�E�j`pg��h�f����bX�'��~�]�"X�%����nӑ,K���w�����&D�,O�k���>)ҝ)��g����`����nӑ,K���w�i�~F9"X��w��"X�%���w��r%�bX����r%�bX����ys$�Y�Yu�V�WiȖ%�bw�w�ӑ,K�����iȖ%�bw���iȖ%�b}�۴�Kı/���;�[�L��4L�h�r%�bX��_v�9ı,N�~�m9ı,O>�{v��bX�'���6��bX�'����uu3E�L5�.�v��bX�'�߻�ND�,Kϵ�ݧ"X�%��~��"X�%���,�|r��G)�ЈFW�M6U�$����Ќ�4�:���J&	]�n�۝UFX��4�X��t�t�Jt�}�۴�Kı>����Kı=���r%�bX�g~�m9ı,��{-�]��(�ss|���N��b}߻�i�D6<�Q5���w�ND�,K����ӑ,K���w�iȟ���,Jw�{���I2]a���iȖ%�b}�����Kı>����r%�bX�{���9ı,N����r%�bX�}�l�y�曖j�Yu��"X�%����ͧ"X�%����nӑ,K��~��"X��dO�w��ND�,K�O���.I�f�i�Z�j�9ı,O��{v��bX�'{�xm9ı,O{�y��Kı;�����Kı?!�}�)��-ˢ�ʳ��PR��J@�x����ps�э�6��M*�46%�=	�(��~��ou�b~���6��bX�'����r%�bX�����q6	"}�{��A'߾맹����.g��N�������ؖ%�����ӑ,K����iȖ%�bw��iȖ%�bw'~��*Q�,�����ҝ)ҝ=߿{��Ȗ%�b}�wٴ�K���D)� a������&ӑ,K��=����Kı<��s:\�SZ�f�kY��r%�bX�{��m9ı,N���m9ı,Os�w6��bX� &D����m9ı,K��I���1�r��å:S�:{��=<��Kİ�����i�Kı?g{�6��bX�'��}�ND�,Kߺw���QQ��GI*hq��o#6�iV	sem�(5VLV��7,tq\��l�O&5���Kı=����r%�bX�����r%�bX�{��m9ı,N���m9ı,O�흖p��K��f�\�m9ı,N�~�m9ı,O���6��bX�'{��6��bX�'�߻�ND���S"X��~����2kV�5��fӑ,K��߷�m9ı,N���m9ı,Os�w6��bX�'s�w6��bX�'��v�fL5��jۣV�WiȖ%�bw�o�iȖ%�b{�����Kı;�����K����HDO}z(~D�y���p�N��N��������
]�i�<�Ȗ%�b{�����Kı;�����Kı<�]��r%�bX�����q�HzC��b�lrq �Q�U;[�X�X��7(4)-PoM��sc���p���*Q�,q��:|:S�:S������,K���w�iȖ%�bw�o�a�y"X�'��]�"X�%�������ҙeV���ҝ)ҝ>����r%�bX�����r%�bX��_v�9ı,N����9ı,K�����8�C.\�t�t�Jt�����r%�bX��_v�9ı,N����9ı,O>��6��bX�2Ͼ��K����Ԫy��ҝ)҉����iȖ%�bw>�siȖ%�b}�wٴ�Kı;�wٴ�Kı>��vӅ�H\,�5r�iȖ%�bw>�siȖ%�by�wٴ�Kı;�wٴ�Kı=Ͼ�m9ı,OP���&"p�W�1#�	$�dBYIHЉB,H��A$�E	!$%@�$�X�C�9ơR�3���1 �p���%�p�� �"@��a�09�7��L�"�s��G;y�<XF�d4�8��W2�`����IHQ @�-a)E���(�cFb0� ������H]�����ՁA���%�BF!��5©D���Ĥ"A�`Č6����!�k���B0 ���	�Y-!����؊[��.�Wc�D��y���c��f���%A�N$!	8�fk��u-�K	K-�@���>~���V[��`5ame����إcOa������C��!J���Xl��IF F�\k_�Y�=3U���Z���a/>�u%'=�j�@v�9G��������{v�lp�Ͳ��㧋a��X5�PlRR�2]eҕ@����c�Q������cm��@wn5���]h�Z$�H�<���.2�X�rp)Ί���2�m��q�p*k43��8S��`:��륌1�[܃3�㧓�ؠw ��.R��Ptm�rWhǎG�煪{5��?F�mXK����T�q+1�A&wv�%շA��p�mdϮ��6��9�1�ɮt�v�h\�I@���l3���1+X�یO(�ڊ[�Щb%���:�k�r��ѶF�^m�: hA����ճ[�����mδib�g��ή�I8AZ��&p�g�kBGTp��qR��Yj�]������2I8�� GZ�xyݹ7F����WC����`�-tPr{iZB�V�BĹ\�E��n�[`�ک�$q��g<��VU���#���هX%,��`����D�\œg����ei�dqU�	R�rn�7H�Y�gdMٵ����-.�{dx#q�����[�*{Wk�5�J�MR�¤�@�u4]k��k��k�y��Q.����r��4%�WX��P������g�Q7ϲ�J�%�3�nP�F6�uT���[�(�n
[��,����]o]�����xؚ6a�9P�'�����Jq'��������v%��2	�N�2`�[6P����F�%GB��nUbk����[��l�+��VՏ`�B["�UE6��v�ۀ����6�PRҏe];y��x���D<��}A�������l�;���yP�iUmKHm���L��������7K����i�[I�_twʠ+@�aP�cun��	˘�FɑBٓu�C�Pܡ���a,���+j�D�Q��R(1ǋ�܀�47�H󾳇e�qӹ,B��܅����/K�1
Y�q��j�p�55����rasZ�Ux �|b�TO�� ��x�|"1�<B`�zE`/�� m�i������>�ѥKۖj���m�M��=��ʷ:�0M�
E�uٗ;B!�۵ìp����M�!�9K������f�I��l�˓c�n�p��S���S�z�/�P1}�mt�X�K֚��.��$9�ͯNԭ�6&��ݞH���=q�,��+*��0h��I�n�v�SM4�-S@j.��#3Q`c&%i.KV���m��n�u%�I�v�vŢ�� !�8�gn�]\��۵�#�`.�T����]�S���bX�'����iȖ%�bw��iȖ%�b{�}��r%�bX�ϻ��r%:S�:}�{K�U�.m�'�>,K����fӑ,K��>����Kı;��۴�Kı<�]��r'�I�5鎔�~�������-2�ӑ,K��;�ٴ�Kı;��۴�Kı<�]��r%�bX�����å:S�:_����ୱ�*jl�ӑ,K����nӑ,K���w�iȖ%�bw��iȖ%�b{�w�Ο��N�����m���B�]fӑ,K���w�iȖ%�bw��iȖ%�b{�w���Kı;��siȖ%�b}�vwY�4]]f
[`�*YX��q3�X̎:ۮ�dkz����-SaF�Pʵo�>)ҝ)������r%�bX����m9ı,O���m9ı,O~�{v��bX�%>�}�ir4�Z�Z��>)ҝ)����si�h�H�	� �/Wo"n%����6��bX�'�뽻ND�,K��}�ND�.TȖ'�����p�j\��&�]k6��bX�'s��fӑ,K���w�iȖ%�b{��iȖ%�b{�w���Kı>�����B�զ�\֮ӑ,K���w�iȖ%�b{��iȖ%�b{�w���K���L������Kı=>��^f�YjҰj�:|:S�:S��}��Ο�,K���ͧ"X�%����fӑ,K���w�iȖ%�b}���ݳVF�1����;]��V6���E=�8��jQv���(���RiH�S+}ӑ,K��>�siȖ%�b}��۴�Kı=����~�DȖ%�����6��bX�%����ՓYa�kff�iȖ%�b}��۴�? �1ș�����m9ı,O�~���Kı=ϻ��r%�bX�g�˝�5�j�%�֌ֵv��bX�'�w}�ND�,K��}�ND��8��	�%Z���"�(����ZU�CE���g~ͧ"X�%���}��9ı,K�{;.d�L.�Y&kZֳSiȖ%�bw��iȖ%�b{�w���Kı;��۴�Kı=����r%�bX���v��3Z�)n�Yu���Kı=ϻ��r%�bX~?��߮�Ȗ%�b}���6��bX�'~��6��bX�'~�:d��3!s4�f�%ͽ\8�bN	%�[����\sS۱1����s�)8���ߙ,K����nӑ,K����iȖ%�bw��iȖ%�b{�w����N��N����z[,[c����ŉbX����m9�r&D�?w��M�"X�%��w���r%�bX�����|:S�:S���=���F4�k�Ο�r��G7���O^�0�8`�.�X�n��4Zm��\[rz�	<�`lp��)W��}ʪ���ML� }SK�;V��wI	��7c����8`[���J�YY�]����W42�[�vmc���$����
��kD���X�Knt�O ��8`�� �ݗ�l��J���;l-�nـl���9U�H�'� ��y`lp�
آR�]��MZfջ/ ��Xz�ʮW���zy��7b���t�T����l��}�� �0��x�\��X�SiS�m��>��vG�v^�d����\+�E�Z!A�۵t�y����]@��%����Dŀ����6
<;`���n��wkp/%��Zj�f��t�IW�d����O,���%�qm�qj!m�V�������
�Kd�F�6⹧�i�:�6�l�c<�:�O	�7���dȊ�V��׳H�m�&'e8c����n1ê��vs������Jp�"�LẌ�)�����i:H�0�p����ǉQh�[/;T����*�O���.��Θ�M�:i�:��V�V�.��ܸ����d��P�	�U-��O^{��$E=��;<�`�ឪ�-g��}��s�
U������l�Xv8`[���tWP�h�B���k �d��;�� ��/��I#�}�m���^ ��,�����wc��$��r,vL�{tmǸt���j�=��k;X�g["�i�V�.RMpS���6� �孓��o�uI/ �܋ ݓ+ ݎ�R��T1�]��V���8c�+�Hݓ+ �c��$��V�TTU���:wm�vL�dp���%�{׀I�� ����*�'Cm��0�����wd���]ܫb���4Zm�V�x��H���=��ǀ����ĵ8���L7K�
���]uv��gB%�N��I����s
��LH�w�ul��nɕ�wc��ĸ7����o�d�jȨ���-�a�&V�0�%�[%�d*]�ؐ�N��u�vG�Ixv���#$��B@���(@_R� �*���}��sϾٹ$6()E��we���l�V�x�L��8`�D*ˡ�[��MZ�x����L��8`[��Ϻ��G(�-j�Ԓ2)%�6������3�!4m��[��:5e���#c]�l�Xdp�;��{� ���mo�+H�8]�'Cm��0��X�p�>�2��˻�lV5N�C��fݽ� ݎ�&V68`��S�wh�N�hV�X�Uqz{<`}��ܓ߾��r*�$�I��^s���>XW`]�T�Ӳ�vʻl�>�2��� ��ŀl�UjKf��i����ۊ8��[�a큠�ǂ���ɺ�Ck��W%�%"e�
� �0��X��}�e`lPR�V�wt�fݽ� �r,�+ �3�\�G����,-���v�=~��>�2��� �ݗ�n�w/����:wm��L�dp�:����s�JOg�k}��LWm	��u�vG�v^�0�L����~��ұ�Q[-HFbCk=v½Ἆ;7c��WOlQa��-�s`�Lqu���������H��c�v�^v���I
�x��k �a�g�֍�c�'d��Z����]��G�[��7:�ni��Ԑ^s�ほ(TWR��8�6�y��Lc��雟]Nyū9	]��B�@;�t��vS�Z^Q�u�@�I-���FbҺ0�LiHTJ]?>���$��y�L%�l��xr��(=�=u-n�y��n�/����R�.i�����&٠j���7c��ɕ�vG ڛ�v"�:-����� �d��;#�ջ/ $�J��m�I�m`l�X��un��"�/ >�Q���c���n�	�� �ݗ�E�^�ɕ�ؠ�An�tS���fջ/ �$��+ ݎ����m=f���Vƭi�k����� ������M�jrL����KFW�@�MZ�} ��l����7�運{��wkST�r�e�v�o �����s�������9ɿ���䜾{���z��T����Wt��+���n�O?�l�mȰ�X�L�ct��ӫ�E�ـuM��M��ɕ�����Dzy[���m�� �d��+ ���v^���ʌvGm-
҉�%��9b�]����Y;:b�����%�%K�o:�l=1X��x�&V�0��xT����鱴]�l�&�`�� �/ ;$x�L� ��t)E[���6`Se�d��kj�QE<�
`F0! a`B��$Y~�i��(NJJ���]��D�p���.K_�_��GS���]kG7��&b�R-9��_�1&���O��~%�m|����b��j0�I�$����'��!��@���)�fz�)� ��"�l�� H!5r�TŒEFMN�J�c }n1�n��n4d���Yᬆ.1��0��"���7�W\\!	�/��F���fT|�_~Ѭ�c�`C�ZY��2B Aդ=�,
a���0����	��i��P�|h��o^��t���Hr�%�ݬ���՞y�*�����:&�JBo���D�`���h"�T� c���E�q*�Qz�@�2 H��HB1� H�
����$`�I2`*B A �@�D�C=⁰ N	�5̬�\0�-!`'V[Rjջ��q)�y�}�dp��9\������6W�^J�e�j��x�L�v8`Se�d� >컥jYi�s4h�c�z96vݒ�e6a5�՚����C��X�	#UVIFUKj�o�ˏ �/ ;$~�W9�	��V�{ح�i4�ӫ��l�:����<{&V�8g�ď#��j��H�an�[w����7�e`#���/ ;(R��t�I�Wn��;�2�	#����rf׀!@<5�	K�dR�ۋ$,$:rBN�H��N�;���'w>�_ ?}7����L�۬H�uvK�	$x{&V���ً�T���;DG#��M9`m�&���`:tI�Ok&r��t�̽��OJ�]�&πվ���<��+�\��zy��$�z̥`��T���x6G��Ur�7}�g����^6��ueҦ5M]�o �d��;�� �엀���j�MZhN�m���ų�� վ��vG�w�e`I�lt�wN�������^ wdx{&V�0����}�A"����]�s��WY�3q���n�ڲv5`����9%�ɹ4��	l���ۤ�]�g�j�#��v֪ӎV�)��k��vR�?J���$�("��1j��$oi�ou
ú��}��T�;��ټ#K��X�HלZ�-Xd�=xizx�=�A�ӧh�l��%��j�M�b�K�Xë+���Ixmb�a3F�%��x� ���K38\m<�Jt�\���!��g�O-ĳ@X+������G�=�Q\cF��߀?l���L��0��x%*�N���;v��ɕ�I0��x$� >�\C�����e�6� �8`]��I�d��
��P-�j���[f�ݗ�H��L�dp�7e)X��ue�&��� l���X�p�:���;�"IS\�ƀ��&�[���E.r���A���t�#N�X0�T��ns�M�
���L��0��xݑ���W�򑺍�g�}��<�ӧ;��:�L�uD��nk��$���[�{��+ �J�v�t�wN������l� ����Xv8`jUڷB.�4�[w����+ ���l� ��HwWm46�۶��Xv8`Se�vG�z����o���-M�2�a1�m5�KNL]Mk���ufĳW
�5ӊ���mi�]���un���<�+ +�K�X[�j���ـun���<�+ �0	������.��t��n�d� �d���UΔ��(��R���$�$ RC�
�Ep�w���'/�w7$��g�31�j��x�&Vݓ+ �ݗ���l�wW��v�C��u�wd��=�UUm���}�<�+ �r����Z����������rnם�����$�Y[�t%v��#��RU�oV� ��l�X�X�6��-Ћ�4��d� �d��7d��:�e���e[��I���;M��+ ݓ+ �ݗ��< �B�4��@�ݻ�.�`�� ݹ���f�׌!D��	XDB�($IF@x(�|s���l��x=WV��bl�&܋ �^6L�v8`�Uz�Vyݶ<�����jN9��ӳ �M8��]�[SN���&�Ql̬#4e˥\�����o �&V�&W�ʯ�z_��J/Ǭ�WM�N��w�M�+ �ɕ�M���;�7䖴�~�$Sh�������6{�Xۑ`[%��e`IS-�,M:�.����r,�d��L��&V I��Yn�]:I���d� �+ �ɕ�n܋ ��w�w��?��q��4��-��#i8�Q��B��E��	Pl�,�7#�-�Sd�5
�@i� ���ڃ��9��AN��Z$̯V�ݴ��ejd`�%Hd(�5��M�㎷m�Ik���a35&�ʹ���]SGh͍b�6#�ix�F�QrP�IX���+Kh�A�\]kp�u�Ƶ��I�\Q�u�t;ܭ\���xL�+���`KYc&_�ἴ�(!�!�LCVy���\�%˪��T1�Mg�(]��5cK5����h�'i�s\ ��ņ
֊Ū��߾�<��2���dx$)\�4]ڷj��X�2���dx�2��%)];������68`�6L�l�X�JQ�t�E�WI�M�6G�M�+ �&V6�Xv����t�*wi��	�e`�2�	�"�� �\���J��ꓯjV)ԥ	���Ì�r˅�,����&i��F�B�@R�iQ��m\m�=|`nE���&V�eLL��Wi��Jeֵ7$����M�H�F�#@�$$�h�� W��y���V�0M�+IЋ����[X�#�;$��7c��r, ݥ[R���M:M����L�v8`�"�� IGbhT6ն��u�l��Ȱd� �+ �]%.r�V��t��uF�f��%'s$m��0!�����æ���tҵe&�v�X�G�vI��l��D�YWM[�t��m`��&V68`�"�7j&)b�Eӱ�[o �&V68a9O�ʜ�s��U��>��y M����*�m��t�0�۬lp�&܋ &��	�e`l�����ګeЩ�ـM� M��d��;#���qMS��ݯ[��`�aKl��cJ��.�gu�5�g%̡�OCƢ�#c=y��|'��	�e`�� �r, ���U�t�N�n��o �&V�0	�"�� I�Шlv�n���M� n��	�e`v%)@ƕ��I6`z����� I��rO>�훒��Y�K��JX��V�j���i,J4M���`؉Ye�v	:�I�v� n���2���n܋ >�J�E�2����y)n|<4�/�T�6̇[���%���H�V�)��vB[v��36���n܋��9ϐ=�w��J���
�Cm��;��=�URD��, ��<�L��&*b�uv�jĄ�f�r, ����2��p�	5JV���>[������ �ɕ�wc���/ $��J��6�۶��L�{��7���@��&��$���*��ATU�Ƞ�*��TU�
���PUʂ����QW�("���D�@	@�ADG�E_��*���ATUꂨ�TE^

���PU҂���E_�*��QW�PU|PU�b��L��ݫ�v� � �'����`����|~  0*�(��`II$ 
�I(�[hI5� 2��O�    � UU   P      %(	UTAJ�
 ��F    � �    f�ZCY�u�$�4�æA��$��B��5݁��mn�&FA���N	9�r2waӰ � �    
��v���F��9w`w88·#Gvt2<<�������< ��t����� ;�2ތ�:2��Ω�< pzfaw8���wU�s4.�     =㛀�n:;�����{=�����.�
�C-�Z��A��=��� ����� �N��{�� �f��=�=�92�X�C�{�t�� w�@    3 �Y��w���^�s�Sf���95L�p
�y�=�h#��/y��806��O6rL������dz=�w0=� �     c0�l�����aށ�4y�6� � �4݀ ك��G�L빺;��@@C@wX�p
`z,��d�MWs�� �ɠ��n�S�:�]�  y      ���OJS��UU �A�� L�  4�QR��      ��U$�&�4� ё��2 تTL��M d� � ���1JU���0&&FA�# ���jIL��&&I�A��S��S��}����~��L<�5ﾆ���ϹDA�T?X(�j*��}� ��!�o�'��Z���z���?��������@`T^ _�$��ED�B"���H�1��1��r��/���ƛ�wn��vgv5�� :	 T�Q�Ib��EEU �6$�H,�#MŐ�6$�Hz��g9 
'@���eN�J 
$��wd  ! ;�U�{�@N�{ �S�@{D�@N�U� @; ;�U; �� � C� N� �\@B��� =��`� /`�ت�  v	؀=�	ت=�؀b ���=� v*�؀v  v )؀���v 
v 'b�`تb b�*����Ħ��PZ��|�G�'��p~�����-/��a�jx��>�x6����R�E���R�,uxf`��s}�5T�E&�v�*�SV�#q� IIR�q�֌/D�8@�TL00-ѥ�Y5@d�w� ѫ���{��8EV��l�]�ɯJ��f���(�YL*5��Y!$�eV���)A
"�	���Q���D��i*�X�[*�U���0������HA*�ю���8�l��Bw� xc Ă�^�p!9���1#+�d�e�h`@������ZMQ��  �@Y�6$v�����{�p��D�D������D�2/F!�N	��)��6��)�*��H�h�	�y�X���xҽ�*�8�H�+3 e]]��(6ư�vz嚞!;�n��!$	0JN�QVR�̷׷�NFdkul,�WmK	W
�[*�Y��,-��A���2�5�_<ԗ[4����<7e��!KBͰ�Lh�^����e��1%FJ��1�Aߒ���Vm!W�L!�,
L!x��b@�0�LK�7P��݂Jy�o8՜h:����R�xm'�vU��H�d�T���twA��#j���"�*�hY��T4�3��X/4M-HQV �\�0$Lг"�2�a�j��n�ǷoD �X9m�����/�p2��\X5fjo*�j�0p�`T	V1K�@҂��
h���۪t��E�(�h"�N���l0��������(V�s���V�$��%�e�$�7*�^���t�x	7����QHF�B�aEB���F4��4D((PŔ��!F��V����H%!b�&�IE�wʯK�����[��Y\�
�
I�ݜ�ny�T«�#4qkƦ(h���&� BE���E\�����p��!Acc.�d!��
X�m�E�V��Ġ�T���j�׆����y�J���̧@�P��	�`� L�s.p�5��a�3h`3�(�b)A�(�$�Vm�\�x�yZ�Y����V`3OV��e83T̺�YV4*��92��̳82���1C6v����TAc�ڨ�Oj���L��
��rjI����r��F��XC�(H*֦����%�eA�DJtj��4J�E[P��D���7�����IT2�PJ(�\%��d(b5(%$	R2�`��RA�!�Qa*�[��aH£B�IV����@��,��]�a5��z6B�����mQ8 L"�ج�:R����ZbH�]͉�@�h2��JT��n�
�R�J�����ލ$62�UY�����QH�%a�tl�n�����+xB��*y�X�˘��(�+ӎ��ѧ�Ͷo��rJ��O���8@�)��#x���%0CV��rP��EKx�f�Xd�;:�ʩ�$hZ �8�(lqѳp8p�
t��"0��A�h� [� b����-���J��P# �����ֱ��g᥽hS�N$�M�����I����b�%�����!a��A �c1���Y�&0� `6�
@"���;6a
<B�(�XM������Uӆ����Z0�`�Xa:s[�s��x2����4m߇����%�CF��с�&GP�$7Y5�ӿ9A�o��J�4�����!W�%^��M��W���٠%2�¬�U���k��
%p9Q!�<vB�d��BF�aLGxH�������56B�Kn�5��M���H֬�M%Q(�	�^� �P�Ad���$B�5.�o5^�A��������I��@2 RW��`�P�;6� ;,^��E>&"I$�Fb��7*�$N�@3eLl���Z��)��
D����"�Ղ� �p�F��5\8fh�ٔˬ�e�mhq@� �M
��]�g`�o�H�䉔D�ɺ*����%Ѵ۷z�J�
��R�S
x(Av��	S�����d�QpNA�cWP�%D��D(�9�<*a�������Q�`I�7i6sj���3d��*��Z(IWN�h��e^E�-:jN8 �!*v��@;W9HNV�Ƞ.�]�d	ln�Ŭm��`EI�UtL�!Z�T�eL`I��K���C�lI�p#	��8Q�>�T(��,"�VW8�$�ܦm���:1]\UOi�=No,@�hK��}5|Ψ�NU�����l�%;��V���	�ȑ�\o�4^he���+3BJGe�nFF�dF�1BA�:E�HFB��`QT$�=�@�m9�pɕ�&�����	+e]��3ӀB�dcA+�i(㫯}6j�M	� �)�v���݃Gp��B���4QN�k�FB�e��uz줧�}�!Ke�J�ap|�e��4!K
��no)�:"{N٫��6o����u`3T��gi란6�ڜg�; RΝ�f��`�%.u��j��2�����5(aE�!�Oe�
l�	惹��!9UE�9�t����L��8��b�v�kVN�ѡ�T1�,%e�D����Q��W�z�7�r��'fm�(A�#���&o��H��	5���jSc�	�HM���UP&����W��;�v�@<���ĭB�F��a�`���HsU��/���m��e]ߵ����ЩǤ$bAAX��o�	a��c&�N����� ;�vVX3Ӄ�͚3�q��@ALͷ{$`�
,�6��w��8Z�0N��˓L��q�8g"��Hٸ��X�'#&�^[�(���X$�ʺXM%6k"�Te�fP�.�x2��E8��{�WU#E����K�1u�b��f$�� `��e>��Z�\�^Vk�<9d��n�U8q�$�@�����ƠTB��djQL���Vʰ�#]�h�(%y�s���	��p^F�"��)"CL�E� ��4��aVƂ�,h�E[
m�D$)����xVer�=4z�(2*.)	Ы����B�35S7%�9,��!K�`m�y��`�k�YH��ၑ�]�Q��%7$i,	EU���$*�_����*��
��;�:p9Zp������82����L��
l��X;m��0f�f���ŦP�LQ
.�Y
J��Z�h��Y{%^\��Y �K��I��4�`���
�:}��	g$	BYB��HW�p5I�m�5B"��P2gBU �	����j�Ag0����-әGC�]���A%V��$#!��IVI IEf6�B��7f4e�B�((�faP$@�ā@A����ʐ��1�dX@�B�P,�H�%!,aD#+���Li�ZJ��	4�"� *4�	1bF���`�`�0�F�%)����M�E�p���!c�w�e�0�RQ*�eU�0��h͗�Fxc
�04�]�HA�
m�M�����|=$�%
��2�TVV�A2�����01r D�.��D�Q� ��6�a[�*��lʛ<8@�Y�$5�6+�̮N&nA�,�$�e`ۭȁ"	M�X%�*AĨ4��J$"����1BL V
E�K�x!L!,Ġ�8hㆊXU^k7�a| ��眔o��z\�v����x6"�v룃g�c�����Z��G:��}��K�n�;��Q����lV�av�{Q��F�Įyzۂ�`N�Ѱ�{���Wg������n��jݰ�:�#�?���*��?������l6�Á�t�T>��.�F'���}��q|?��&j����   0 � �� �@ n�   [d���m�                                             �@                                                                            ��                                                                             t                                         	���7&cwd���f��w\9α���������w0�dgvh���b�`V�j�UwD��p[���J�m���s��B0��n�����`�W"�%5��Uv���y�v��uʠw�㯓��\\!9i2��B���"�Y9�)����y�PcB�	!�˲mݫc&�իc1;��nZ{C�b���8�;��	�<����y]�;�9��%��DB�O[Y�`�ـ�wTuSmKęص�B\�^��ﯵT�<��S�D&��[n60j���+ְ���A��V˃�P0�-tԐ�]��n�Ui�ԮV$�#c*֪�q[B���[�UG;��u-���t\J���u�l�]�J�	t`;c�eZ��v���{vخ�L�kv����7n�j�M\��u*��z�om���K��v5�D�*�5�-¼i��5@M��S6^em��6�� �m �9���jK;p;d&��nGe;3ETv�u��EU�qTf�Ut��_@uT�*��ۻ�m�� [#P͝gmpK�(��>U�m�`d�5�HA�%� 6������٤�[kmr�66���nW`��R���K�56�0� �� �ۺ���՜�j;K�V�:e]�
��[T������pHk�m 1cW$��JkA��Q筺P�����h5#�Ez��n� �g���pTL선�d���.T�\����"���(>��	��ӱT�9en�ā�*�uUGK}����۶-]�'��� �cS)һ�+.�k��8��.�NsҨ]x�T�>�kV)Z�
*�.j^Zƕ�_UA�E����;6:9ቝp�*H��;sf2#�����+֊e�d��^��wf�pcu�*��/�c��pUVSp��lݶZ�"z��UUH���������'j^B[d���ۛ*�ag��Z4]5�K��2���U�ݫI/���b]t����5�%��-Q�6��T�;ME�t�����.Ze2�e��1N�M�\�u&YU@y�������)%��m�t�x۳�V݇���jݱ؝l�`ɫÙei9<�4�bH���«�j*�IK�ӌ+j�[��;;8}TR�������nʱ������㚫�cJv�Kլs�����
��&�L���by�Y^d)�5UUU��qFuۮB7.�@x�)�l0��X�`;��T��F��z+NBU���۪T�
�ҍ�m�q��`�ۥ�5�\��9��ؽUyIj��i�ۅ����Wb��P�Y��Ȫfӵbݜ��W�����yБ���|�Z­V�q[u�R�3�1s�X���K���O�K�8��Pg:�٣�eJ�
4n��� cg�v˷� �	U*ڴ[1;wZ]���nsWhUwnz;"�Z��*�Aع6�M�������|/��p˹�ӎK���6VT+�-��)��g�sʞ%��NGg�jonv�,k�������8�v�U�@*�5UԮ��sj:e��[�t�WR��^Y���ܪ�uR����3Xԏ��s��gcv����ŉ؄����p�Y���k�n��ѴuЫ�Aa 힊9H:
��ݸ��;�9x�ǱU�GnN�b����EP���`��R���̹^C�F(�"����j��tmq�����vҧV�N��;q�ѽ\�0�d"i� ��7] ���Q���d�)�u�u���h޼��K�3��d��g�;��;E�7=����ۣ��:ҫ��K�S!�ݥ|T� �6�b;ep�mױhj5f4t��m�=]�d*�nsf�ψ�!ك��z��v6c;�o��m=[��,���Upy�3�/J��`���[d6�phj���v�m9;k����e��"l��V���݂U��,���[����?�T	Fgvz����}���j��7F�6Jƭ\�6�j�� E̍�$&��b��>@]v�9�������UUY�D�SѨ�А�̑.�nɴ lU�@J�R�n��]�F���K]Rl�*��TUm[T���'g$�l�m��	d�W6Z�u��d�-����� ݒB���[,Փ&ɹ]��W)m�V�K��iۖ	�T�TQA�� ��#�� 7v��U�C�
��}������Q5b뱉�>�ځ�An5;�m.Ŕ�*��� 8�j�`�Q�Sj���	�U�WRQ�o��������̂ĭ���V�ڨ8R%������� bf��e�յ�����0T,�mbL���+-UT�lT*� �&�M� -�@l�F�YnɷkX+��+ln�M�\�ma�en���%Uh &�����v� � 	�ETj����٠*����6bde cwA�i� 7v
Rl��wq��n� ��ё��r���u��UGj�f
Z���t)�N�tԳ�ZwjU�Ӄ*�n���� �	���\ڥX
�c���^C��r�Z��ѱ&9% [kw@ 1%UU+� jj���m@]r��q�6��5;Gj�m7t���L�q��[URŒ��m�� �����vv�ǋn8�p��UmVڕkf�^�U��qţ4�U�@#�d�M��Wk���X*���(k�l�X.a�U�H�MTO<���@F��GS�.̫ �8�r�[����Md2:�^�"��6�n�q�������<��^3�������*��R$u�6ە�
�y��\a��(vZ,�=c&�3v*���� 6x٨b�U.��ä��c,�O@U�����m ���%���.��UG�P���J<$n:�r��l�S��������s�7\�6d�3PSiyf�1P ��x��$�Y6c���"���UJ�����7Vv*�5�pU�UT05��+][[W]U)���b �g�*�cq�Q���R�u��q��h�+�v��U�[�n���:$6����ꗭRD��v�Z���ey��^�k��m�y%���մ `$-�U�� &˻���- ĀIm�n���  $	4�ʡ!m� �6M[�p�Ą� [�@�	  mʐ7t	��c�%���ڶ�0�� Z����Q����U,UŇ9�{N��7]���@uhIm�����UT�T+-T�5l1��u���l�]UnP-�&*����Q�V^9]��Z^ek�uԼc���MT�Mi�uQS�qE3��J�@J���������ue;z�T�R���>��I7�A��+��t�z4���V�I��K��3�4T��:���D���J~�
��?�Pt7�(ό�!���C�y														@@@@@@@@@@@@  �$������6>�adA���	# I�0 h�B �`�) On������~?8����
�®0��*�
�®0��*�
�®0��*�
�®0��*�
�®0��*�
�®0��*�
�®0�Çv1��Ç���lc
�®0��*��;����ϻ����x�PhS�~�P���G<L$  -����JN#௰DҶ�� 6��X��R (�8x��/�R����-P⦗� &�7�C�� ���b���
��B��b�
8��p"���J =����8����z;T@ ��A^"�X � �"�+�_�v�v�O|� �| ]�D���6�LO|@�`�j���}T[.�@u�x"!�P��"����P��6�J�h�S�LE�@Y hȬ4����(G��OE�U�
�4 ��0K ��� �"0"���J	@,x���P�G�b:A^>�����rE���HF$�x��0/<���E�N�� H�jE`�!	$�+����)���x'�ԨT�$Y�
`J��L"TiF�����$aK!P��PS* K��X� �<p�8�X!J!ꂘ���O �(��C��A�D-0��@DA�1��ht�>�UUU˻������������u�K�b��H��P���H-! �5RF����  A�D��k�=�wn7/�9��c��+/)h�(�B^Y��Q�Dٻ*����t-�/#h        �              m�              �       cy,ͱw&˼�nv�l���Xy��^)��۷a�uc,^�6�v��[7��6=���8�Ʋ��l�&�n�[u.p=aՇn���n���vdܦ�ݛ�ԍ��*��<�v�[��w+�su��L�qÕR��8�J�Rwod�s� ykk���<��$.��ٜ�ۦx���Ί�<�9!�!�C=�:�3t=�- l�=e���.�P�ug�8��-�Y�Sø�na&:�}��lw����N5k�G\Z��h���cm���:�m�Bu����a��\�*�[��9���ZZ�d^�d�1mۚ��bzz%㚻��틴�cnp��'��!k
��e��Z촦��{e�Oeh\;���������[��6�@d�d|��v�G\��x�뛬�N��d�ݯf�E����W�;rPh�溶r�qY�*��,A�mkcy��!�1:{/N��Ȼ�(	4ܝl0�(vT���^��v�,�;��+��l`�,��b��Ƴ<u%��nu0�:U�CE�S��O`{�R��6�V�ï;�3�\n��Cӧ�A���qչݵ-��n��oc�WGm���[=p���̓�oC����0��\�-���+��%�v!��nvr�<�CVuV��{u�pFP����6܄
)��`�;T��%�X�`G"hU������ƺ�;un����M���6���Njy��g7v6m��eM��`*G>��>� ���#�#�z���'��D-E�S����`?���<��;� ��  ��  ��nꮩuu&z�;��cd.�3i��1�PK]y�m�;��W.6�1����--v����ˆ�L�� �MN��Ɏۭm���`�\��\f.үS]�F�r��5��-����r���;n4k�+4Ֆ�^�8 ��U�wwweʕ�\��'���{��8BAH�32�+��uLV��8���C�P"�f���̹)9,�rˊ����j/��g�S�����-��)�j��0��e����﹍�ZJPa�Ԥ���co5�_qU���I�[����C���_s��D���,E����m�ك'�v�`����tm��tceN��( ��S�J�lKo9�w�٬u���<ԆĤ�W�9�,���$I�YCb'�/xj�1�����/-��9NAFS`Wo1�����y��@<9�u��a2�j��o8��b��+����̹)9,��i�_sx�}��^k�@0��m��m���*�6v���\�؛�����O$=;\�68����"�Ȗ�f��k��}�fj�ZR�,������co5�_sx��3�Á-�3-��C��8��hl �D�@1������4��R��ĩe�i�_sx�}��^뎾��HlJA����@=�q׺⯹�����m���j����`�5�dۊÊ����5T�݋�:a�s(�M�]���늾�.� ��t�i$�L���=���6F���(E�ky�e�I�e&i�_pqVqG�@5��=��77�����iK2�����=�<��&Ń�`�Au��s�ߤ��S%�Ԥ���U��7����x3�b�^F�(�.�q��eh৵D���/0�-$�&ĝA����՘8��cb9"��Ǐg))NJr��qW��Ó�
��:�X���y���X�I�9��{��;;�Vg8��Be�,#)��D@��c���_���@<9��I$�d��u��*�x�}��G�SIKm��l       .�l�i��c\Ԋ����q��f�X�`yx���lPj,̶���L*�E��0g�������)�`�vBxЭ��ڭ�ܻ��a�cY�ӹ�,v�6�AN�^4�`3�6������9`���
��v�֮ŵ�9�H��r}��ݻ��t f�ԋ���n֒.��jŝi���7��X9h&e�H�BM��^w1W����^k���ȶJd���R�^o1���w�e�8��1��AiJd�ܥ)�]���k���*�#;X�CD�L�fe�����/=�*�G�Nhc��))NJr���U�?�P+��z�k�" ����m�UwW�՚����V�ӷ8�q�s���������Ԇ��LI����{�W�_�"��q|5t�˔XDJl�k�p �dA�IM4�� �		�4�#	#%2����Wg��f>�z35�Ei��e&%2�j�{�qY��ޠ�����rRrZ���qP ���c3����{48��%��fZ��<���+ٮ.��h's[m��`�.%�c����E���[���c1n�!��7iJ�fԤ���b�5�gsz��Ѥ��a��ɗC;��"�sz�w���FP�y�򲪳s�p���P�P}U�9��b�u�_i\�lL�����@;�b�u�gs�њ�&T��)6=^��_w8��}g]�s:��< wef�VlV'6zy��6�l('B����	�#���IFE-JN.[MX�w���e�+:y1��̹)9r-4�ә���7�
��+�5��χ	D��,�T/9 �u�����nj�ZR�%�wWx��9�3\��9 R��ੀ l����D��a��ɗB�o8����xм�_����m��m��3*d�:3Gm��nh��lClS$G\��G��������Vo1W�
��+�\u��Ȅɒ�2�/9W��vk�����4Ba������m�Xpp�)&%�m5C{y�f�x��ùg�e�Iː�M���m�/;��:��` tG��}         չYy�!&����t�n$Wmm�.�Y�ٍvK��pk�w]m�Mm���r�k�E�򹺫��ۣ���n\B^���<�Շvˢ��-���.��k]��Ibݻv:)w`a|,�����K���l�S��,ʲ �sνvۖ�u��Ng�9��� n��ݧw`�ѝ=��:?��N�����t��ή���l�߮�^�����nj�ZR�.[FS��ޡ&����@vѤ�`���dˡ���Vo?�f�/=�x�N�BRa��̷��6�W��vk��ҹ�)K%Jn�f�^�ۮ+7�7�+[m��{����F]y�PLgZ1@z��t<Z0@7��zw.m�2����qY��x�o	ǆ�r�b[��T7���L@�L�.� � ����|�v *�X��f\��D)i��{��@^^����wxph��ʔ�ˡ٨
��3�\Vo&75j-4�%�h�`f�����y��@z"0@��� [s(ٹw6�n7+/1۞��[�cp�1x�%�R���,1&[&U��y�f���}�_L��
L4ә����m��������{��!2R�J��o .�^}��ז�m�  ��~�ܙ��ܦ$A�BJ(�z�:!+V(T�������N��&A1�l >���MӺ~M��a�y��sP���XML-�(V�w��0���L5e����쫕a(�#��x�������ҵ&��x���`j�� :9=�
��1����d �C��� �(�w00Hs�tRo-�z��/�ǻ<ם1����m
��u�UE���L5E�Q����*�"M��L� B9xJ�!�,0�ehѪ�,e�r?����~x� �|�"��6v PV�!0��!��W�A ���IG��hF���Jb		�9�3�}�Eh�r*Yr�M�y��5�f�1� ��G�%K	�  �M�߻�/{Ŋ�@;���%Ͷ�m�ܣP��F��t�+
������%�{\�Tr���L0��1[�	��C=�㻼<%6�	��B�P{�}�ި��?��\��-6�S7�1{�胛�+q}z4�,12�2�����s�� ?  ��<�,O������ ��ח�9=䟂&mɖ\Vo��ޠ3}�*���ϗ� ]��v�͚�Lif���ra�;1q'[�������NOŦU"%�I�g7���U�����8��B6��)�/=�U�y��@V4�R�l���y�⳹��@;�c/'���h�-&�*���X�z��Z�wxph��p[���{������qY�c�Q"#>�$'39�}�fϽP        �����/���Ύ�@�W'�n�]�[صN�R=vz�vq�w`ǇN�{M6'�W��$�|r�َ,ٶ�7>����ص���x�v��$����%Ol��7hnrt����qn,k���V]U)�OF��P�p��K膠@�@���m��m��-XY,��=��Mk��]�2T�ݝu�^�:+t*��Kfe��y�b�5������=�8*KL�L������U��/=�<{��@��N\�n+7�Vj�����}�r!2Rh�M׎~�D����g�qY�8��Be6ģ)��� ��Qy�2u�κ�� ���˛Y��s��sqX�d�k�����Wv͒0��XŁzϟ=�λ�Э�= G�/���?	r�)p��i�_���|<�(�Q����7ߘo~y�A����j��)P�y �5�9�������)$�b[3.>7�y���~�=��������Xbe��tg������@uf��@�}Ͷ�m���2�8�[���Gp�C����@;^�=���{���������5�w�㳴�D&T�� ��}��͡���u�`�r)�%L���{{�s����F�[iJe>���� E!H�B+TR�`@H>� Ru^�������!�L6�M�C3�qW��n��f��>�JR�K�ӊ��}� �f��q�": G���������89�mι�#�WoPé����Uc�
)1A�BS�&e`߾_��c35� �/7�^�6IK%�.dKټ��D@��y�o|�ޤ:@#>�KS2�2[��Cw�d�����rټǎ��E�&[ �o����5����8@�E!���tP�!Э�o���}���%4�$��@m�w��9�؀s���0��[�"�.�n�ɨ�=�k-�i�ٻ�.KRi�%L�����^늿k��xpv�Ĥ�l�ڡy�� y�b����32|%ʔ�!K�ӊ��+5՚�_hq��85$�d�N��!�U�b﵏DD�sܸ4���.K3,^��9^��|�k�,>�ۡ��?_]3���         H%ݬn]Yf��t�����\b u�d����{IE�4�L��v�J�;<v�`�zslxֽq���W�r���i��'\��P�n�s�X��N�n�����77c���;v������q��O<U���cC֠��9�/Y�9����2�W���ݑwq�Z�%W��8���i�9tg[H\j	������+�}�B���X�'B	l�(L�}�V��5����x�����i$��}�� ��9>�ȫ�8��B6����~�@��c3��^y�D@�������I�R�j�g���yޡ}�
�k��몪���D�v�Жy��N �Qs�C�`�8]Z��T剩R�D)r�d����+�`:���q��B	�&Lʡ}�~�4�A ���"R�f�D�)�U*��Č�D��ֶ�}��s� �j��JC9s2��w���c�7�����f�%�2���˨�{�Qy�1W��< �y�9��P(K���*��~D|#7����כQY�u 5c�����wtJ��s�<��j�]d߿{M3R�Ji��v3yD���{3_� "��qz7��l��S`W���GI����x� �ӣ�a�RrJ��oy8���}��F ��`z���@ �EU�>�!�>������+�Hh��!&�OOD4~S��~�c� W�뎾��h [r&L�B� ]�H�7�^{�f��m�ÒR2Y�%M��ט�O[&�7l�wR\�6-߿ww�>��4b ._��;7�U�B�P�������-��Cټ� �E�y��@W�_ ��(%��L�qy�xo���"'>�1���#��=-��ْn����o�=û�}�����@�H�� �*y���=�yܪ�fa�˪��_�������\f��*��d^|� $՚Y�8]��F��B����7���V�￟{���p��@�\ʔ��{�{���!��  H�{�v���eJrYM�ۊ���""�@{7���  ����h �r3.�f��k��f�������]�IYYUX�:*�|���;��[��r|@�"@ު~�x��2��3,��7�}}F�ޛ����X�0������J�� ��;��'9�o�s$��!#��f�T(->@��DXIHF��+_M8�5�.�AfƊcK*��!����Ȑ��*��
 �B@�P�B0 D��HI4�e�l*�fc�����Q�ID	���47D���*�U����|��d���5[��!	F��l�%j�M�p!�D�Q(�$!(HS)�J/)��	��0K�v����oP���,j5��:
( �HńA0��I�{�Z�M,�   �� p!
T�L�b�%mŶ����   �@                                           m�&]]A$����y��H0>�ۧ�v�-v��&x�/^ݷj��ŋ����M�K�s�v�ڗ�7xh����1��!� �=�6P�am�k]�(�ú�Й{�&֪��8ث�=4���UQ���W\�Ф��i_F^Ç�y��El�7ݺ�X�l�DwJ���K�WmF;f��M\�źB�rzrE�dr�t\6��ܛq�u�t�v��
�XL&7�W�ʹ�C<h���{1 �-Qt<��S��n�kt�r�ٵ� �K��uh��;sI���v̅���=�yc�%�z�[��x�۶L!{�$����o���p�wG��bܢ��e�'�l[����^��.:xWN���2lu�����D�;�\�a4�N��Ө���rp7eT�M�u��g�����ݎ�|��Dpٴ��l�A�ir����ɐ�Ȳ�P�.�8x㘵V^��E��B��+2�7!�˒Էj6���SM���W+;l�̵��㐛6$�ۙ&v�����Kp� �E�8��켈N�ݐ�q��]ő�%������M�q���tg,x��A�&ƌ�i�F�5rn�"ݍ�^�f��Lr�C�]����8�⌾�Q��6�j����h����d����{D@�;����s��I��!���J��2H���Qf�k�c^�v��_���h)�?H�W�@�i)>�8J�߂�}EZ�E��  ?@D�����EzSm��m�       w���ζ��kW\�(���3ё�u�"�%��>����o;rv�;^��<�v��r�͈�Q�O�'g�c$�km�}v��nڹ<g^t�\nP�'��Cv9�Z�Ĭۀ�4�nG�2n�Gcy���N;c�s�ݛv�ZS�e�o.U�VK¬�W%��MA�fg2��]��ٻS$�3q�n�u�OE�e��.�,s�c�$� �njJ!-�ḑ{ߌU�՛�"��yǳ�}-��ە):���"{�{7��y�~�"��$�����ϧ��^hc��� K7�K؃#E�c�!�Paʡ 'N��oz����^(舃��csg���r�m6�y�ǀ�X��=y����m�qvl�l��FM��&�.��1ۥ�Z��pN^�߿{������&܄��c��`u�1�ٽ_ �$������^�� �-̰>��� t-
�"0)$�Ū(*4JAv4�N�U�q�;���I��>w�IiL�Ė�e�߽��ǀ����/ӪudKd332�"�����ޡ�� g�돷��,��e��_j� ����y���J��m�[�vX����s�u�r=`�:���n������}�L4�آ=��3���s��"� c=�����(0�4ҡ��� FH��:7ڀ��C؈�ww��rSE�-����;�7���Ѥ ؃ۤ������qY�E�&Z��>�����b��cG@ 	��Ώ������ne{�h�[�B��s��~��&b�nY�WvJ[x�7&,���Sò���ȕ�]�w�tIiL�L�s2�g��*�X��=2D��}C=<��&P-�\̧y�興7ڀ�o1~�}�p��e�-�-7C=��� �9����2 A�Y
\�fYwY���������[��>�� #�
��_T>
?J/~�a���߈h�r�5C3�|"#�3{��Y����|�o���֥�mc�gucVx��t�����
�5!�A�.\�m��~�{�y� DP��8���)�&eгG�� �>���y�^|� D��JJR�$�2������c� �o����{;�-)�ɔ��ˡ�"{�Qy�b�ꎈ��y���D�Ne�Ţ�w��T9�t<��k�<��!���<6O�@        ]VT�MՃ=��l��q�Ov3���J�7t����Ere]sGk,%>�i���%sX�{r�E{Z�]i��	�]�dC]����=Y1�<�f9��]����|��tv�5����z��j/Ы]��Wtf�s�[��[���Y]�x�y��g>s3/9�wۺ 	�M�����ej��{<7On�A�����%.���������lM=�{�o5���~� "�G�_�Be0�JS`_�����M�y��C@ zt�qT�a�I�3����| A��{y�^x�\��n\�m�����^sED��"��Q��"Jp�hP���D ��~�X9�z���b���m�ۭ�ś��L묖{x�ծ��ȵ��1�ڭ����u�m�[$�2��p�b�5�7��DCs���xx�)�
S�.���/��
 t�=�>�>�5��4y�Նk�g��W<�yL�L�Բ�̷�y��Q� �y�>�q�{9��R̶�t< Fo�{�W�X� y�q|;�	��d%)�={�V��_k������m��rC��+���)�`:碘�����8�M8�������ۡ���j�{�⯵��C�@�={����%2[�2�qY����@ No�gy�_�����Jp�J���n���j+F! � H�
#�b,/� g}��n��v��iL�2�ʊA�w���qW�c�D^s=�ĹH�R��t/��< @���
���y>u���� �l�#V����\�ĖӺy�X .�yy)8��FR�`�L5,��m�W�b�Q���@(_��g���nT�-�i����F�y���q���>�����fYa�R���{�nm A�ߝ�@no�Hr���i5C��w�/7�U��  �>��D3����&\�r��o��� =y�u�z��F���6�m��,G/nM��nu�Ĵ��s�1�<۵��.�{���N�2�o|���b��~ M���I�]T�
9�@{{Ϣ����*��"@�@	���r���M)LPAo�@�D��93�ͨ�>ߜ0�舷��@)nSI��!/_Қ���p�*�ʠ5^bI�KCnF���c��"2���U w�,Ȉ��2s3��g�����        D�40�������v<�ݞ-�/<Gh� u��D�>r�X�퍏lk��v-+�h���˰Cl��0�v�������svl�n�0Y�3��m��Q:Kmr���ڻ���9��O8��F��qv*�Ѱ�����s�Y�wb���-�߿���4�� ?_�Y�e=]=jIO/8�G��n��N��]?y�$�R����8`U��;�c�HSy�$���*K	̴�rN{�Uq�z�X�8`o��o�CDL9�D���^�;�pˎs�m�v�z�*"e��S4׵�a�kٵD��< ��ɒ}�~�*L�e�-)�$�G��I� E���$��3']�ē~�Ϗ<�f��r��+Υruy8�ǫj]:W�\嶅Kׁ�]�߰���j�={,
�8�s���x�ݜ��	I�I�3-�$�y?���  ��aU�KmrQ	+@�(�j�[�l����y�9�RN|�����t@� L���}%�r�NCM�D��0�;��?�Dz��~�UN��2I��iKL��t́�ޠ�9��D��o�&� M��d����S-�KI�D���Q'� ���*$�s����X�w����@�ۚ�KI��<�];���
�[�5���׽��y>���<]i} ��+��ԃm��DG")v�*��͊�șp� ��s7:ၗ��ڢI��O�#���FKfe2eKjRM����$�oU;���I$���m��I&�t0~` �A��HM�7�RJ�Y��놪�sl�!�	RRe2�%������6�b�
�9W� ��9�!Un$��T�#
 ��A��M1tH��&� y�x��%oxxI5�C^�R�0,�ai
#
(�@B��CƸ��qB��s5`h����&m�%It�ʌޫdc��,��*��`Q
j%H�����> Q���tL�E��D��qC瀡��^�t#^(�Q�C�Q����8��":��ϒ������y�53*\	KBqA��⿳{@��_�07��Y7)\�i1����%���w.�����t�_>��]I=���� ỬbA#���c�[�\�=��-��Hn�~�3�zN��[���I��	;��d��m~� �"1w�L���*�d�b%&�P^8`v�u@�L2��"&I���)i�%�CtŒw��ONo����s�O��'��BL'r��A��s�z��}����2O�6����B@@5���$��
�I�-2�}2s��$� ޠRm�P}����Ż��m�ۆ�]��vj�^#)[cm��jx�,&8z�ϻ����hL������q(�fU z�w��R�0/o(jfSp"Z��yT�d�+�����c��H��JY2�Li�2�ײ��ۆg9�Ko0+�yށ���ܗ-�M�D��{�������h���
���7�D�ۊo0>�""�7�Ig�����D^ff~fs�L�~�>L��ɷ���         ٶ��.�6mf�Wq��%䠻<v!p�ؘ��i��S��Kr�ٹG&�4����:�U��rۣ]�q٭��gQ��Ş��ݎ�Yl*р��N%j�5VX�h���`i��j7�N׷V5v���9�v�íN��G M��=���w�����UU[!҇���-�t��(2�7���c��ߺ���t�.�iKNY-&��'���¨�o92Mn�p4~��	��m�o��sfO^�`gs*(��V�	{�BY	1%�f[tI��������@O�ͪ ��X�p5(�$ƒqA��n�(nmP���8��`^�P�̦�̉��P�ʠ69ٳ@w��|�*(�e6�m��.2P�
�ƭ��=����i���<*�hP�e��}�ߋ�`U���i������_ٵ@|������eJe�>���a�� ���bCd���K��z�{>g�$�y��$9��[_ �q�\m�R�[b�;��d��ڣ� @#��2N{�d�x>����K�У������I��L�X�B��ݺ�]�M��p�*[t��f���p����Wv��;�]���n���Z�����-��-�:6���<�b�ߵ���4q.�%3�=�ᘗ�!�R{qWb:��l� ��)�e)i9����P^���T��`Uۇ�	��9m��i��bN(��ޠ=�,�Ȉ\�D|DA���]���5�F��=�a�OznR�	��c��: �ر��p��m��G���V�l6��ؓnh�8`o#ٕ�wە@͖E�'uUUn��Dv:7\�y��9�t��n���A�F�/�I������fU v�| �Nw�d��>���l�)� ����*�8�{6X��E��b9	��Q, �e��tI9�L�Y�3�3#�ܨ�;��t���ؤ5
\�Jf�@�����2M�6����G]_&�6�Թ�A�
b��d>0>�{<����v��y�'o� ���<�X�A�6,k��6�݉�Ց�[���~�J�vsbN��ͪ ��*����DRn8a���R�-�cP�7@˗���{�d���3�9��W� dBG���~��m�6怿���n��u@��$�,Г1%2e�(�@��
�e�P�e����O�;�>����P�����4r�0;�̒}��?�#�A����9���g>g9��d�ݓ�        *��=s�m3���Nuu���&��4�^:���{��m�sۂմp	�������Ǘ�z����!���8����$�n���v�cU�V�m�B�i3cڈ5��aY�e�^!W[��v[���k����l�Xƽ��w�ׯ~����O����� Y�ֱ-�r��:Bv6غی�] �#�����z���\��Զ����_�e ������R�0����;���y�[�m�Poe�9Ď��6����!LPjŮ��@=�����p�G����ʙa#bN(7�����T�y2M�1�'�@~��I���L�Ķ�I��v���^�d�`{q����mkm��m�!J&	>(v�����]���vݩ�Xcv�N����7�j��?����|C$�gu
$߷��z �;�$�.�I��	32�b�9�0�`z" �s�T^���@o�,�]	�7ll��˖��f�jA�͖~G"�}z�y������M�6�n��s>ϥ�W��n8aq�y�2�b��H�h����IY�2O�@��(�~ޯ��I����'ϒ�� �6f���Z��t�s�+/U�=v�V���6ݕ+~��_\��]k�F�{����u@��_�0=�wfT�	q�A{�U�s��f�ݷ�yȈ������cIL: ����k�a��4��Ȭ� �(D�LHB@$ �*�*ާ\03�ʠ>Y�lJ[nf���ȅ>�����I�f�M�$�,Г0�h��I���$� Fv��$�y9'^|bI�9���� cU"湱�'2�-�pZ�*��v5aq�����{w�n�Y:i��{�T��f�ܷ:��P��̚������oy1�����!#���_��U�y�R����%3A9�0�7��=�� 	N�޻$��ɒj�t�S-0LhSܔ���8�Ϫ����{�I=�{�ԟI��� �)P�����yfT���'����?���d��0�7���6-O��m���uv�I<[��7Y7�)�]V���8�x�np��&a��%.�R�l�*�����{�3��G)��[���ĥ�&�h�~�s���'=�TI9ޔ� �9�z&\KKۊ>��;nꏹ�${>�r�&������M&��P��Po%�Go0�G8��P�ܼ���L��-��ٱ,�8`wm���J���������$�I$�6�m��I'C��O�B0#
%6B�1�P6FF��p�J�4��Ѫ!%.f�7upۺ��T�϶l�uT`j!I���*đ�(�Ejh�!IC�M��#$$�@!$dAc+�q		!��FB� d��7�$�6>x�h��R�3-	!�e $��a���D�����Yn�                                               U7=��Tp!;����U��Wme���b1�#M[�p朄�:R��b,��ZRa2Ӂ��n��f}��IN�:�qA�Bm�Ol����<<>Ԩ��#0q���#�
u<��K@�:�썋Gua��7�������j�G\����%��k�#q�t�-��6����F�7����Yvu�w���ϒۍ�Ճ9Ӯ����9��a�q�u�z�6�4v��IX3;�-�*@l�݆ ��LA�����Zp%:=�A��Blc;P��m�<97қ����e{#�θ��$܄Z��ڌ+Gg�P
c�]����k�-��ٷ)�(3�[n�;m[l=I�y틶��z��Bc
���v�Bv$�˅��� nP0��m���p�q*.��m�m�r6¨3Y,9+q���9�,��0��C؞�����j����mɱ��Q�^Pv��kZ�{nÛ�4mOgeOFIzL�<3��Y��Gf$��j�v�<i��dpC�͠ԯ�-�5��T�0sl�vd�[F�U�ܮ'8�BX�]Ғg�Y��ЩU��	�j��F_��֫Z�xw\�n,hz��Q�Ǘ�����+�{e�N�c�5�\��= �th.��Vꤺ5�GW���b�e�힙�Ƨ=,]/�Q�6WlX6��8����Y��l�ݸ�`�ng��#���8~����I
#�(UT�(�*E`
�����'��O�}� >��#��8*�<v�-�P
����D>��w��I����ٻ״         |�t�;ޯ'3(�0 s�����Zv���g�-�.]]7��N��z����f��m���-���.-�n��$Y&�Od/O�ϓ��z;a_�݉ �쉎�BQ�6�`��#;�Q	��k�ٻ����y�Z��%=�Fe2R-&RD < ʁ�ݶ�wq��D�e�b�SX֍Bv�f�9][��q���qӨ�5.���ksj$^[�}�_���o9�H�KۻM�2܂�4���c��B�2�ٳ�����,@H���m��*[3,]�;�}TI9�,
�0;��ܛ�.%)��bJ]�!/f��yQT���*#�����t�1�)lIÙ�R�k��2N���]I'~}�'/���e�g:]t�l$nrf�hөtE�\6'?�w��2\��j0�t�p����H�l���p���'{���ĦT��@'LY$f���,N0��T�{����j����I9�8��yМJ�̶�5+ߥ����q/}���P�[$�L�'!*f��c�n�0;ܺ��B^͖s2�R��jRhS�06#���@=�jIמ1$�~|�@#)�[����Dx�h�ͱ�\ۧ�$q�u��t���.�m����_|��`Uۏ���d/�p��Ӳl�S28cBn�;�K�9�s����]E����곑	���\1�nR�9�=��$���=ח�S�1S�~7���sZ����r�N��E�!��Be�(��N��{2�1/f��A������9s)�Թ�ċ�ګH�8�6hn�`w-�$����w6浻p��m�6�sd��݆ tJ�㇊�Sb�k,[U:�N����������Վ."�wە@e��!�N9	Q3@v���ďf8`wە@��RK�tڔ��8��q@{1��e����`w����I9%�)�'��G���#ٲ���eCȁ�1.D.r��P�$�a�Q�R���]�?� 6~τ]֊$�/��RE�XIˬH=����[�i�p��*���}�@f���Z��Xɹ�E��ˍ��sv8zz����7��L2�-��m+78�y�I��&��TA&������#��E�!��Jn; ^��m6]�� f�,
�p���L����MK�ޠ�ݪ �l���,��d���3�?wu9r�$�-Jm���\jGrp�A�c�}�T�����ა�3@v�j^�p��*��7�L��~�$@��{%��m��     UUUh��:	�;B�i:�b����݃7G<Z,gW=�k��,g��̦�F:�����G��p��b�U�>";7g�%��.�Ύۡ�L.p]���*ܗ9��,k�Φ,v��ri���fv*��݋j���Rڀ,VO�{�{������@3l�ËNn���6�{m\tO\[]�̈́�]�wsMS�����X����2� ;O�>�����ϱ�$��	6$‿o�D�/y2N���7��� ��9��>	)�hc�t{��/�c=K�LHﲨ{���L�JRa�Y7���ܨ�/׵A�`{�vJl8��I6�i{#07���C�{6X���o�UU[`i=U<ܐru�;��Wt�x�m�a���d/�%7"bj\�u#s~� �l�/�fR{�d�wu9r�$�-�tI7�^����}S�`zX�nw��oU'O��F�7�«� BG���R�KD�AQ&�~�p���uA�{6X��9C�9(>��}�a�G�v��ϥ��ǥyo!$��SbN(�p�W�5��с�[�^�ζ�m��"^�@
痶kq�\>�N촑��\K�
��.���-D$� {6X�)�W)}�T���$�-�-!2�n�7�俄	�����Poe�#�n<�8d���I�2M^��$���G�B,
#�I� I)(�b�I!�6������/$�^��FI'<����q)�Җ�8�{�� ��+����^�*���R�˄9�m��G��`TGo*(n8`Wv��۝m�U�\h��S`�}Oc����Z4 ��+ع��%!��2T�@v��ݷ�:W; {5K�@�Sf1X���%��U e�;�p�!#�o!9�,ؓ�׻T~�`W���o��m�vJ�˂\�J_�/rX�pɺ�|�.��`�		ȥ
���ҤP߀��s\�rNy���2e��$iQ&��d�������Y'7�MQ�w��I<��x &MeśU�4g���=]��`Nq��)B#st��^��W}��~�wX;�ʣ�ׯc�=��{,�Br��ТM纨�oy2Mf��7��������MJI�*[ ^�>��p������nU~��&���P��3A��mCَݺ���Ȅ��K�@�I���`�P�|`o�����/~��k��2I����@B ,D"���!J���1 |�K&�em         6n�i�;,\��T�u���n�;.�5f٬;u[������q n8ۤ�l=�z�&�&���TdQcsH��pA�x}kN�\�ň9tv�S��1�t�]�=�9=�+�h�BQ����v���E���rTý��Bo�fg�s��L̹��� ���VL׆C�^����1Q��Ǔ(t�	��D�#p-�+���;}TI7��&�X�m�w͆I��.G���.\%.�;{0��BGo0=��]۪������A���%�@{5��nݺ��KԌ����1��-Ê�\0=�\� v�XlB��C �٬�嶜71@wە@��_<bI߾1$�;�������ˬ�M�./V!}�����.�I���?~���B�i��u��|`{��]˪Yy[	4�V8U��Ԓ��tka��x����o.��\U ��� {6_�H�̠rK��d	����}�Tg!#����	v��p����S7*e�bE��P�e�Wn}͈��{i{��6$S)�NZ����z��9��/�* ����w����|�m��pp�(�L��+W�=��T��aV���7rZ�+@�������7@s�n��[�Dw�BW�Mj�Md&�-��=�8`w�u@̉`Uۆ^�C�-�.S��K�����n�9�<#�_�����I|�i$�I%_� i����J~��I	au'aE4Q)�UQ���hb�ż��d%2UĐ!a���3%�Q$ BH)��6$��-$�#,2@�!!�)��RB����%
�!��-�^.A�;h�#!(�y
�HP*Y	�*6��X���0�@�n����0#(���VJ�MJ�~
B0&�vGZ�8�
���VB�IUL�U�ʎ�7���P�	VJ�beH�$%	%F�D���e)#$aK
HRŢHR�$"F�P�BJQ`J,!L�iutJ��2�>g��!����Y,��4VU�*�d�3EՖG���}��{Fj�v0XN��*�P!&)P$�pR�p���!AQ�(��B��Qe�Xh�ѫ���8���`�<q�0q��:��p��P�+��!��z ���ޣb p���/����DpG������<����^��mJS.9�m�?G#�_�İ;��߭���TI���fZ0�	��*$����n}�T��`�]��m���U�U�];Ÿ+-�.�����]ў�*V"�����N(5^�C�̪Kٲ�#ӎ���Bq*(q@wە_Dr8�{6X�p��ۆ]�rTH�SR���R����\�]E.�g�����0�1�K��\'4o0*���˪q���P�P֯^�I<�=��AC�nf%6��`���� {2X~1����fy��@��2�c*nX�Ka�)�;��5�g�:P�:��[���m�������D�*����02�鹅2��̶�����[�e�$wە_DG75�	5|p����=��Wn>���T/f����0ہ1�L�+�j�eW���a�!{\h���(��8�\$������f��80;�a��Cj��Z��� # �u�
%@��U���V!��Rzm        ��%�5/M:�g��N��̷u!m��۔l��3�Rw�<�����v��]�.#�^u��@�5G��n/;"�ӷ;�vàL�l9����F��DZF��t]rn8�(�'\���-��nI�ql�u�)���[�s�s��%�@���uκ����X����U�z�z(�x盄W\�tb#p�m������v��}�DR���jإ�S-����T�0;�]Ps$h:�r[!C�)ĩ�P��
��Q���ȷe�ۜ{ƱTˀi���_��� ��H���8`j�Zhr�Bs2�Τ���`v�{�Qԓ��}�'�����7x�5�9&�n�]�V�]<`�qvyQnb��^�x~�~.rS��3R��W܎G:�%},�n�ѐ�%3)$����Dd	B��b F6$�F
$e(� $bh@����TI9��&�i`{.脚8�\$��^�w�ݖT��=�Q@{g$ȒfF��B�A�#�f��h���Sw쨠+�]P�D6ɗ-L��K�50>�!�v;����I'�ԓ�|�o�2��7u/S�����)�)���%���&%.��Y�xc�;��0+�u@˖/Z`��9M�71AK��� {�,
^����W�LIʖ�Nf[w���>K����X�A,���3�d�Z�<ޤ/��������33@u^&]�`Wr�;�,���ȓp�Kʠ;���-_Dr"�}��}4U�`_f�~`#-l���K-��i���tx�H�:�lH��q�kp�8�\$�z�j�;�,
^�����ܗL�4&�t��v��m0+-���^�{�Ez~��-�#���9����A���� ��:�s*�C�.IJZ�;��]�� �d�<-����%\�SCA�%�(��(�%P1�UL(IEQ
��rm�S �l�!���CM��B����R��np`Tm�s��DB�2r��C=�Cd�nt����3]�vz纬\k��.h�&�8Nf[} ��`R�c�G~ʊ�ܪČ��{r��2ff��N��Uۆ��[��e�q#3
%D�T�0���4���w=,
��e�&h�\$���+z���;��[nٸ�R�����R�Rn�i�pƕ�n���ܪG#�ؒ�x�        ]�)��F���u�:=+5V��.�M�:�U��&p�`�������/kv��f����5���h�mr�k���1k��[Y��yd��ږݜ�q-���z�Nv9p�eΈl=��٪'F����ئ��끛��κ:� 8lݬ�mdI��!�Y��[�Sb�8�X�lc ���m��Z��;��}�d��\0=�ʠ�L0:��p����R�P�q���̪ ����0
��b��(i�������5{vh�8`Vۆ����jR|���ˠ�#��B^ݖs0+m���"�o�濠NR!�	��i�p�K�n��T�w�ڒy��<�o&lG5���\#V᝽s���g�r�0�F�	��̦Jq@w1���� �d�+��컢�0�\$�o;�� � d6L�&I��&�Xd�ɹ�R)S�8Je�$�%�뻨�;�����Řb"[S*\L�3@w1�}�QAK��� {t��uv�U���K��n(�8`Wn�R��#~�$���>o� �,�fi��:mOj��m�gz r���&E?���L�!˙r����� �d�*���ӆۙ���J����r�{����
�p��r�#/ {����$Nf���]�g�4�O�����$X�	�JI(�@`� 
ww�mQ$�jd���\4М���#鿾�0.�j���,�8`{n�0L$�	8�=�ʠ�N��8`wq������m��Wd�\��u�v뙙:�s�<k��z�u�
��[��LhS�;�,
�p��˨�+�u@b�1�%L�I�4s?�Ȅ��0�9��~9��� 3s�|��e8�m�|����H��,܌��
��b�؆��ޠ��ڠn����A�m�"U��D\���d��8R�>$�\� �d�*��5.�8`/{Vw�v.��m��p�C�KI�ў��mXA��g9!��+�s��.�u��~�~??�
�p��r�H���̨�d���q@w1���� �d�*���wD	�&6$�J�v���e���H;��ݜ��"�,I�
]�	{�s0+m��{��@�[��&$BM��Kts0+�����jP�Jd�����"	�^�����I$�I%www~�
 ĀB#��bā�!!"�$$ �`������]@���A�Ã	���T�$0�;�A�aa�L��"��1̗����h��"@��*aM������%%@c#6�ͺԪ�H�"�$ 0%j�����!�K�ߎ>�o�'�<������P�bJ�q` �%���! �/�e\��J���dJ�p�w�f�*�w��m�߾L���Ud�͡��!�)eiIkF�P]B�Y�n�!6��3�q�D�������BB�Q|]Ne'�9tn�_W[ $`�!���kZ֢V׉ ���J3��!"@*PD8@��t
HT�H�`PB�PB�UJ��UD��Q JeJ8D�H� H0��q�P(؞7����}�+搞�c�                                                �l��C���-r[�0��������8��UŞq���á�G��qyw���f��c�#q�j犎�Q�����q��ި�`��yܨ8^^ƶn�gP�l��=EC��؉���������Sr�ls��ZwB��d.��g��^:�Ӹb�J��\!��1�.nq[��C��v�t�1������v�'�����ͦ�m�>��0n�tl�Hָz۱9�'<�m����l�݇u���=Wk���N��{�lr�t���������㳹8�ݓ�.40f}�=Q������wa.�wZy <�-�xe��gm��>���\�ܫ��6�EP�	��{1��^�t�:5D��ӭ���5��ܖ��8��b�"s�8ݞ��k��9��.�ۊY��K�Xz��2E�m�ڑ]ղ"����؃0��k�G��ջ<khE%�f�ݬue7N-4�$�,�f1�`���p�����h�Lj��l�s���\p�)�i<:�wm�g^z1g.�,������ۥ��è�v�6��m�(�n���N��#���I�0\��x��E&Z�Wmu"c��c��t�щ���b�nS[X�u�\�pY:'u[qp��8�mK�ɍT�O��|�@[����tv=v� ��IԽ��/,�[6��l�J��^� �mشl�z�J'=�ݢ><T:Σ�W �z
�R*�@$PW����W`�`�Y�;�\�;{�         '�5�Z�)n:�3T�|ݰ�k�3�qq���m��oS˴ۣQ�Fyd>���8�X��g�K��zĚ��t��5u+���-�]�ny���BZ���d��4��q8t3�m�s�=�؋[qv��V�ݙ�䋂y4Q�b���{�����{ݘ�ꪪ��]�B#�̚vj:��;m���h��,(`���ո��&m�$�k���6��d缿�72s�X���H�@�s}�U w2X]�
F[�_��8S2�%5.] w2}H۟R�p��rꀿ[�Ȅ���}ٟn����n�������$�[r6�n�K��ၱٽ��I߾L�ku2O� ��sm�ۣ�6ؼS���n���4L�����{"V��vP�FĜt�ڠ�K*���uw�d����Q��S-12�}2N}�� ��sc��`�e�E��0=�ʠ6a�����4��s%���W��Pw%���\��L-�m�@��v����+�,�#��f�T����׻T���h�#ٲ����u��� ��m�*n.����S�9���[q��N���z2픺Ͷ�V��$��$�|���ʏ��r)��2���JdS3@��|�s0;�ʠ�K��K	��I�IQ&��w3r�v�͈ E��@�<AZ�׾�N�M��ɪ��� L8��'r9ř�ݬH/\���K��TP���JNe�˗	K��K ��`V[����Pxֶ�UV��5l�TZb�힍H0n9ذu�k(�n�n������b`Uۍ���o:�uy2M��:hڕ)�Gfs͇���G��T%},�C�^���e�!�s��T��e�E���L}�~���L�|�Թt��`R�L
�a�7@�_nQ's_ҙ��M՘�v���� w2X�7� �6,.�jݗp���u5��hq�!��ۮʔ&���Jp�D��Ts0;�.�����ue���	��6$���ePs%�K��Gw*+��vu')�˗	K�}���v����]P��15�r�-9�:���2M�mQ>����{3��@]EMZ	&JJZ�;��]�� �d�)z� �d��M��         2��˕61�e��(�7��	FY۝���Vw�.1��Cر������5�ϳ�P�sև��}������_V��8L�,kOnq�Ywf3ap[�M@����s��Ŝ�r�q�Y��j�k�vc���7b[gޫ�� ��,�&3P��,�up]���#R ݱ�\	(v�Xҵ��O~vח�@̖(��d[�_��Ȕ��%9�����:�
]ܮ0;�ʯ�H���e(r�)�@yf���
��PY�wu	8%�',s*��c�v�����Ii�컢�C�q@wٕA�%��`u^&_|bI��fs��̞u����$
��-����2V�qs�k�n9���I+1��m��s]�x��|>��r��[t�1��W�2�e�I\�{Z�6� H�� �H1���i_�y��$;�]Ps%��ے�bT����Z����2����e�%嚘l�?B̍�ƛ�P��T�d���ͦj]�07/*\�fS�2���%�K֞�.wr���}�� ���m�����+�h.�]T��Zڬ�mu���Tp�m uX��34U�`U�p�����Yr�H��|NB\4)c�TJ^�p�#�̪ ��XټU�BF}�x&	���'���jI7﷙Vl�dHHā�BDd�B 8�T������Y/���79ϕIBr�̹hR�F�:���0+�u�A{;&�i���fe9�<�S���.�����yܶ�m��D�cZ�^��Z.sj���*��5���1����
Z�;��i}�T���AܜI�v���52�Թ���^�U�A�R+��=�"Ofe&����E�ӢI���4�����{.*��	�ڄܦ�t�ĲMn��7}�D��`��d�3=�	�6�K�@w1���� �d�)z�ԏ�9�2~m��mË�:���z�8�v�GnA��Kixq�z�-�[Ȧ$KI���I���59�>� �h��\0/���JC�3)�B�A�g�l����e �*�պl&�R�r���L�s* �*�=�,�ֆL�c�KU�|���ڠ�x����*��_̷5.b�H�ݪ ��)]�m���s��cЂq�        �t���5.l��eؠ9W]vw2�\]�L3S`у�c�_l��7����B��`+v�7g��M��e읐�H\N!�ׅ:�o7m�2tjn9W<����1�%����avm�U������$t3�[,��ύ&tpNL+c���g7:�z� n��g[�ۋ2[�:���\�^B6���j�rf���*Ͷ�V���O~�,
V�X���9��ʠ2��2QI�fh������TP��V$ݝ��ȉG�}�Br��
XԪ�\0;ۺ�!#۲�H��L�pL&a��({� �d�)]���p��Gf��ʖ��NZíH/vXR��&o\2x�{�Tu!m��6�m�%,n�b�� 5����A��sl��u�uƫH�$���10*=nܺޠ/vZH;e�]�U�*fV��\��d؀�HAI ��B8���I';��U�� �ܭ�RKpR�(>W�}� ��)z�U�ၝ��N̧�MK�A�s���o論嚘��`W~��/��(���34U�f�w2a��nUN��RO��=��}�\ٻ�]�c�p�8�f8����'N��q9.�<'�o������E�fUbAﴖU�~H[�|�$�$ˊ�ܪ �d�)z����d�\9Rۙ�	7@̖/Zpq�����ͤ�I$�I$�0	'̃ {k�
�n3aT,��4^Z$H3ZL��i�����{.�$#LѰ�F�<��U��Tb�Cd`BD!9�H2f��)�2���	,�k*�B�e��3L�R�AT��5`B$��Ʀ�*y! 8��� ��j&b��
%gT*4J2PB�QƊB�
��lK�CWYc.!K��q=z���T��==R�``&�'"�����A��&!g����uS�yu@b�2��m�Nh�Y,
�p��e� w2X{֚��p�8��T�w{�B�ڠ{%�K֘qw4۪��bU�V�=��nc;��5��Ƕ��a���$�z�S`�)�d��z���s�L�s�?�""�w�p�J�ܯ�J��-K�G����9�嚘�0+�]W�y�J6���Q��vᘗ}�T��aK�n�9&[�d�T%��ۺԒ���4�MH,~QI�TFHU0=
N|ך�jI���	���%�2���*��{vh�Ēu��$�}�΀I�	%���սz�Vݵ�B��Ծ)@��a�h�$\lW�m��~�|�Vb`wq��m��0�ClC�i5D�����7��$�{��ɹK>�"d���R���2��'>���۸�29�ɟ}/R-N�^���ԉ���s�����n�H:����eC�i��Lr��2��w%�%�x��p���s���9Ørs��         �����Ι�n6�k�9�>�;��6Xui�9e�\��;�v�::<;��XG��[۴{\��]u�9�v�vcyܦ��Ia�v�q�r�r.�ی����u�x���&��Y���v}r�Oݧ�l�S;���T��aɒ�v�eƸ��ڨ�s��f�gN� �2��u75N��L=�^&<�V��TbYy�:m���^�/����
�`���� w2Xwu	�2��̱̪��>��eP�e�J=i��|��IrL��;�ʠԽ�,�K�10;��[7T��)��n�󐗾�`ue�`Vۆw�T,�Bbm9�4VZ`}�ʊ�yT�����Ϛ� L�Y�Ԩ�V�\��V<<���1I53	&ԅ!�)����M�&�6����s���-0����LjĴ(����V�   ����+�,[�����y5�$�O���,�s1�Yi��ۆs�T��	�ڒX������Sۮ$}�u@�1�
��NeG"�5+�{��~�� w2X�������m��	zz�\j1�����]�3@vΫu�x�+~����ql�e�@�ͪGs%���&�r��K�\O�6�(2șn�'=�_��伯�jp������"9ș>Y��ClI69�怵��v���  �dBHH0d��	$`H�>&�} ��f��sZ�O;��$�n�!���n[D�@����2Of�Pw%�˳�L�r��H��9�1@f�F��ݖb]^����{�u��UŌ/�s�v���S��۵�76��N��{\�B\�R&[n] wrX�<��wq�).�L�/�	�l�X����O�G�30>�ٽ���r#�H�ǂrK�8RƥP�\0;~���K��8�n�'	���qA��7�@��D��|���C�A�GӲ4�FYq1`�H2I#D��~���&�~�C&[�	cIK���H��L���p����n6�m���K�M�,�%]{VJ�0lؕ9:�.��c��:Z��m�Yi�]�:��uAܼtܼMBd8sL�s4}��#�nk�<�S �V��11�s.b�״�Tc��z~"%-�{�s;�0�=�.z�8�4ܺ �׎����#��>�9^�7�D^?���6L��e ��K$��Fo�Y'>�UM���c�@|�79Ϲ��s��r�         .ب I�v�u���A����U��k�C��ˋE��G���<qqf6G�O-�̷����-�U��n4r͋�R�n�,+i��0m�l<���:mnM��_[��]c�ۆ!�ϵ���XL�E�:�3YW����̋��f\�|��G] �95�N�m��Q��R�c-8���V��"A,s+ �c�_���^?��s�<�S/@'�$�$ˊ�yU�Ȏ~DL���:�|��p���qpɖ�RRƒ�Z�{s]�S�n�.��N`�M�婙����X�p�������t���9�
%��mQ�z�÷2^gj�=�x��<������ q68D���0٣k�lg��Z@g��2���s\�"cL�n;ԋܪ���:�����eEwi�*dq"i�t�o:�� � \wrg�Y'oXd�go]��H���0���%��:럵T�c�~�� wo������Ԫ<���{Q� �ͪ �ٮ��s����&^<�N&I.I����x���� �ۆ�G;qu:�m���/Om1�����k`mY�:��f.�Hq�78z�-.�P���{s]���(�.����{!{��������32�bA� Wm���Tݼu�i�2�&(�*Zԓ�w�k�y�H���VVL��-{������&%�&\��ͪ�$j�����z�}�B��C�i�$J��ĉ���v���N�;�bO�����$�?>� �w���/a��c����,\N���,�r��Eml�Y͊�����q0;�p���� ��:/2�'��%�Jޠ��P�켪 �渠:����Č�y ��I.I�q@^�� w3�A帘�8`V���d�&�A�{w]K�q0'�ʊ}�rH�%������p��\ԓ�{Yv�$Rۙm��^[���c�w�T߾��Iߞ=���\܉��m\���L�j*W�ָvsn�Dg�b:z�Эm�?���۷� �f?��G:��q0f�jACc&\��=��@�c�:����{��*e�E.S�@��@ue�{n�]P�x&&X1�D��-0;�q� ��U {w]��P��[IƥP�8�A켪 �鮀��I G��333i$�I$�I/DH"$Y$c$$�!$I�.���#�>�t�%/�h$�__D���"�@�,�� $F,a A���@!�)R�Ł�FE�DKaB¥F �!�H��IHD�$�	x�$ �����	�j$$�S��%��`��P,��.� �i�1�J#D+u&�#�$L��K�Ѥ!�
5(��c�&�h�B�SCURWr�P�ǚ��z�	Mnd�Q$�IL���Ϡ޷A$������T%E&4$b�����b��VVf���' �P�#R�I�9E���x3��޸��Q��BJ�(�#QK��R$ �Mh����"͜�Zw6f�ʲU��!&�,p֩��v�����K�D,��*�/t��n����?Sw�����i@                                                k&�n��KRm�WN�N�f㵤;j���I�6^3�en:7�;��I�eD�g�.o�w_ �`��-{�����!�Vأ�ܖu����z�8U�am���<�[Aq��/.�cC����0���OGm�8:�h�sӺŸy�����j:w���y�zV���t�㓵��n�I�)Qs����iL=ro<���_p�6.���n��/kvI{]�\[�c��d���P
�:;P�G9r�f޺y]2�;j|�������/mg����q���gXv�u�Y©����Oh�ͬ\׭���]�qK��c{=<��ڤ���s��́�e���nq���6�`8��%�@��n����^�R��v�sWLn���i��`^���xvz8�km �wc+v�m�=��p��I���LЪ���4\c�}vՔ��7
��[���0&�'F��cv]�n�u�/l�������ӆ2�K��Ae��pS���q�u�xk���j;Y��Qg����8D�[N��OA�2�Yņ�n%���沥�U�wO4�)��ؚ��Ʒ��w#uw';spr�k�
��nk:��Qu�����C�V��hkk��&���B7N��-�Q`��=�Zʽjt�
���N݋	l��a��D����^�ڃ�7M�t��n�ם����Ēc�]�P�F��3,� ����M A]A�C�0��"�+�C8���Ѕ��I������       <�oy{��t�bٖ�i��9����Է;lj3o���|Yunq�X�@�C��\���^7��6z�zx+st�n�jΆڣ{=c�)�u�+<�.�,.G���4:�;e.5�Ob]&�8�uJ�z�;Xr*�j5ǵڣ��ܕ��3����~{�ۻ�������"��z�N�M7GX;s�8:5rr��Ja��R�P	�É��.>o�z���à<�S��=���jY2��ĥ� {w]Ֆ��`w=u_��${bwF�6H�[����-gɁ�c�}��u��D{sS�sK�R�+�p���� ws��L�e�Ȥa�r�����bd���O���} veĚ��\LD4�ui�w�MS�ڱ5���=0��E��)�m����w�u{2h{0;�]Q�e��a26"�V^a���W�����|�6+�b |7N�СD�W�TO�s�y��L���'�`K���3>p��^W���%_��@y^����'�IrL��;��@�ǽA�z����r!]�FR�r5����"a�)t�]�N����ޠ�9���m���h&Hp$�u�tB7/f��׋k���]p"]{N�f-%u����?�h;�p������G:������9�d&�L�'w�?�@� L���Iϳ]�Ny�BG܈��鬄�)NH&pܓϝ��I&�����/����^N�P�p��Zj�L��Mˠ��;���]��\�/;@z��8&G"%����p`lw�Q@wo*�;�z�I�g��@,�3u0�̚ܧF���u��q=.�r�.Q28��	8&G�'%�c�_���6��@z�F���'�IrL����� {s]$��pa��ʆ�rL॥!0ؔ�!{s]r:r�G!	�3�Q*D���15�TJ�~޺�f�`I�����NQ��R��&�TJ� \O=�ɉ���TNy���Q*%D��=ޓq*%@���BiG`�����q*%D���{;�e�(�.��i7�TJ�yݘ��Q*%D߾{�&�TJ�Q9�{�&�TJ�Q9�{��n%D���zWoy��UV�g����ۚB�nc/l�۝��Z���z��1���ʅ��MĨ��s�{�'�����y�wzMĨ��s����J�Q*&��MD�����+U�K��Y/+2�I���TNw��I�|�K�Q<�>LMD���s����J��L�z��`I&o}d�JE�R�/4��Q*%D�ى���K�q7�tbj%G��q<���I���TO>w����Q*%D��ʬ,�ʅd���iȕ�TO7�8��Q*%A߾{�&�TJ�Q9�{�&�TJ�Q9����L	0$����L��(��LT�Q*%A�}����Q*%D�{��7�TJ��3�Q*%D���15�TJ�O���>��W�*_�����        ْ��Oӫ���ۛ�m�JC�;&��h�k=�������75Bv�rk�g��۴k�8���Eg�選��mLZ0v�zȤ�Z��pnmv3W���v�@�
m�N�0�-��2<���]�wl(��fx;v.]S#�2�g��P@+ra_���@�
����fffff9�d��M��N8˻�f�&f�ȑsB
��z���n
����TJ��ߝޓq*%D���;15�TJ��{�Q*%D����I���TN��ΙyyW*�2�34��Q*%D��x��Щ�q*'�wF&�j�.%D��{�&�TJ�Q<��w��O��%Ĩ����fY����]]��n%A���~h��J�Q*&����7�TJ�ϝ��;�Q*%D�ى�5�TJ���˹W1��Ѵȕ�TNw��I���TNw�ޓq7t��s����J�P>"��{�15�Q�&oO֤��)�r�u�	0$��>w��n%A���gf&�TJ�Q9�tbj%D��}���7�T������5֝�vru�a���n�x.1`�U�%�{NL�	H�s(9m:�f����&�TJ�Q7�tbj%D��}�{�&�TJ�Q9�{�&�TJ�Q=�����K�d����J�Q*'<�MC A
r&D���=7��J�Q*'����n%D���gf&�TJ�Q=��zIXf��˼4��Q*%D�}����Q*%D�}����Q���dL��gɉ���TNy���Q*%D�����.eaU3%Vf�q*%D����w��J�Q*'<��MD���o����J�P.\M��y��J�Q*'K�gL�������I���TNy����Q*%C�<��MĨ��s�ޓq*$�`g���0$��L��m��nN7N���*:.9.z�[����k:h�lZ�<��G��.��i7�Iq.�wF&�TJ�Q9��I���TNw�ރ�9�TJ���bj%D����n��E�RVa��J�Q*'>{��7�TJ�����n%D���gf&�TJ�Q9�tb(��L	076}jII���-�P,����s�����Q*%D�vbjGf,
Д� ������<��Ou�MD���{�=ޓq*%D����!�.�%K����n%D���gf&��J�Q9�tbj%D��}���7�T�.'�;�MĨ��|��|�X]�VY2V\��%D���wF&�TJ�Q7��I���TNw��I���Ty����Q*%Dٟ� &���5�7��2DEhڵ�]u<m<\*�YR���!s2\��I���Tw��I���TNw��I���U�s�vbn%D��|�F&�TJ�Q9����.eaU32���&�TJ�Q9�{�&��#q.%D���15�TJ��;�Q*%D�����n%D����gnt�ˬ�feUU�q*%D���;!����TM����Q*%D�|�zMĨ��s��zMĨ��Q��;EՒ�auw�I����`\O=��Q*%D���ޓ�R\J�Q<���I���p ��3�)"t@��"k|���J�Q*%yڝ���Fd*�&�TJ�Q9�{�&�T����}�4��Q*%D���bj%D��|�F9��l�l�l�w�_�kv퉳p�ӳ	�r;te�a�Rp�\�DA�m�b�}��d���s�����Q*%D�ى���TNs���Q*%D�|�zMĨ��{��&\��*�++3I���TNy����Q*%D�=щ���TM��w��J�Q*;��I���T2ќ�r>߫�9&F����\���r�By����Q*%Dߧ��I���TN|�w��J�Q*'<��MD���{�\	�aJh��@�L	0$��w�����TNw�ޓpj%D���;15�T�.'�w}�MĨ��{��@9p�ؓu���G!�+�w���r%D����u�bn%D������J�Q*&�y����Q*%D�4" �$�_J���?@�       ���c[�ɛa�]�N6��f5��*�k��.��k1�a��qn���[�<���Hg%����;�to4\ݶ^�A��r�n�oF,�3�z��'F��x��h�7Fu�xNFx.1�YyR��ohg-�"
&!{Y����2�>g9��{� o��D��&nX������٠pft8X��k�g��-߯w�{��2TO��f&�TJ�Q9�u����TM��wZM����s�����Q*%�%����FU��auw�I���TO<�5�TJ��|�zMĨ��s�����Q*%D�ى�������ֲe����A$Nw��j	"���u�$D�;�PI�=�A$O7�v����̕�YW����H';��BH$��;�MA$��0I�5�=��AsZ�e�jQe�t  ��pj	 �繂H$����&��	����d�̓�33�����&�eݮ�������`���en؇�\=Iŉ�ǻ�<��<�w�0N��J���q5 vs�L��*T�
��@$@&����{�Ԃ"uT<P炫J��'y�В)"y���A9�p�$D��==$˓0��2Uf�pI�o��	 �&���j) ��`����o8DD	�<%4ҙm�˼В&�TJ�{��$�s��H$���{��$��?;c��w�$D����|�*�Y�WWy��A<�&	 �&���ME$}��hI�7��PI3����� I���&���a���p�s�d
	..��L�F�L�����γ�&s$�w���j) ���u�$D�;���E�Á�� ��}'�RLK�r���RA<�wZA$M���A9�p�$D�|�Q7��_��J�^.��4$�H��{��$�s��H���333�$�I$�I+�8� �dUv?*<�!��g
�,sI���A�<U�n ����yF�L0�U4A��e�(�#©C{8�AQ�a@m�S8Y		'/[�©j,�"� l�Ja L������P�M�g�M��J2<S)T�<��XTU\*��*���	�@��C{�WxHI&U�5��D �u{ �z�	�/ZG:������b���5������U�Vf�6������	��!S��%����}���f�IFS�0�q9�sF�l�!�'3,D���s`�:�A�P=��C��d&�@���B ���,�J��P]��
OC@@=Dz��KHZ���46���� $_@^*���)� ��
��8BD�y鉨$�s��$�H���N�¬̺+%e�7�O<�$�H���q5�M��u�$C�EeD�>bj	"�vw:IXf��˼4$�H���pu�P���BH$��w���H&��$�H:���uUUwb�p]�x1l�D���uN�bHq�7\�0�.L�T3%Vi7�Nw��BH$��w�� �	�{��"�D��zbj	 �
�gK���2��BH$��|�&��	�{�	"�&�縚�D�uP��	����? �RKe$�I�$�{��0I�5��j	 ���В	"o��&��	9�O=�fU�%�a�$D�}�&��	�}�ZA$M���@��&�ߙ	nB�TP6;���$D�W�;UwxVUe^^�pI���ZA$M���RA9�p�$D�|�PI���ϟ�~�	�fk$���Le==-��T�)�!���s�-�b�d�%bZ�;�ϳ6s�'3�~kPI�=��I_<��!7�N|�u�$D��|��Yyp�����A<�b�Q֨J����MA$ϞwZA$M��q5�ON{��V��/,��	 �&��q5�M��В	"o�鉨$�o��H r=���D���:�t�@G#ۛU	"�&���j	 ��`�	"k�{��$�t�}��yy��ʪ��	 �&���j	"����	"k�{��$�o�{�	 �%���>{�ʫ�ڼ��    ~�t   7��ͨ&n�n.��fNl�$��Y�%���M����ɠ.���n'��\m�#��l�Fnq��Uڍ{c;�M\�Q�>s���{Cf�mi��K]�n=����幮4��arp�)4dN#3��%E[hGytr)�l����s3?9�9��s3-u� �ٷj�!��WL#)���̀/=�H����W&ڰ��{�XI`�	"k�=��RA7��u�$RD�;�MA$oڞ{
̪3&K��BH$���ى�$�o�}ք�I��q5�Nr{�	�%P�'���T�U��L��yzM�<J�+�~kBH$��w���H'9�$�H:��j	 �����BJa��r������
�H'9�$�H���j	"\M��w�$D߳ޝ+2U�E䬽&��	���I^��&��	���$� ���D@$@�S˛m��`�(�7�O^�i��c���n�fA(�k�}�?s�dg,lI�9�{��$�o�=�ք�I|�q5�O9�$�H��V*�%Vi7�Nw������"X�P�Dm8
y�7�wPI�	9�0I�5���ME$�{ǂM6̦�e:		�y�p(��7�p�$D�|�PI�|�ZA$N�gr��!W����n	"��`�	���q5�M��u�$D�;�MA$oڞ{
̪����0В)"o��PI߾{�	 �&���j	 ��`�	"| C����ffffe�Q�;^m�x��������)�BB�c��9��+)a���r	 �|��ZA$M���uBr���I]��MA$S�y�L����2]��fhI�7��PI�=��I]��A$}��hI�=�ޝ+
�¨�����@|�`�	"k�=����|`�!��A�D�x��
��A3��kA�A$N߾p(����h���)1B"����MA$~y�$�H���H&��	 �';秤���
��U�I�$�s��ZA$>#<��pI���I_<�PI��}�ffUW�1Ϯ��u�X�#���[���1��
-״�l�W�UW�A$M���A7�L0I�5�=�A�g �	���ք�I����6��2��DD�0�D�5��j) ���BH$��w���H$ߵ<�f]�*�	 �&��q5�M��К�D�;�MA$7Xb"06�}'��%�e9MT�	PO;�kBH$��w���H��$�p�!$B0�dB0�#���5��q5�M���R)�Ri�t  ��p(�$����I]��MA$}��hrd�d���fs<����� b�sb�Ww`��ag��kl<Y9zc�.uuӂ�ͅ�{�;��	�0�$D׾{��$�o��A�A$Ny��&��%D��I�uxL�˗xhI�7���j	 ���u�$D�;��7�O<�'�TD�;���`�ĉl̺��""}�U@�A$NxwX��H'9�$�H���j	 �+�}*�33%^eU^hI�7��PI�=��I]��MA$}��hI�;��w.�¨�%]�pI���I^��&��	���$�H��{��$�za=V��"@�H�H'�da*�Iy��        e�h�3[��8P ur"玝۹by`���a�W\+i��'��K٢�� [z;i�/W�d.W�}����bCJ:�<
E��{q�3s���%wdf�	�dI��Pf�'�t�/n�6Yn��fǎ�sY�-،۞N�N,�1��x�tU�+�T�^�33333Ye�ѝ)rC�\��y����j����`��ܦ��Ӵ�̫�<A$O|��&��	�}�ZA$M��q5�Ns�0I�<ߕڞ�]��%�^^�q5���{�	 �'<︚�NP���H$����&��	�7�ZI$�r�N[� � ���D$�s��H$"k�{��$�w���	 �'�{Ӧ\���R�Qw��A<��0I�5��j	 ��=�ZA	�y�8DD�|JS�h��	"o���j	 ���MhI�I�;�M�$|�A$O�G;��ffeV�z�xw53�w[s��N�+<s�u��%�sY��ؤ�aU�*�i�$�|��5�$D�;�MA$|�=�A$M���j	 ���Rm�2T��Yt  ��p(��a��l P0a2�
S�6 ���H$����MA7T%|��hO�J�$O�|�>e�fE�*�4��H'����I^��&��	��{�	$��w�����$����VF�%�b�D`_�� ��oN��I}�wPIpg=��I m��OL��)��d@$@�w��Sq*%s���L�PM��0I�7ߞ��L�I�Ͽ=�� 3sXkx]�z�M\�V���k���Ԓ�=�N*�*]e�o�ݷ{�M���A=���	"k�{��$"�z�@$@&oxx4RM2���� U	�p�	 �&�{�MA$�{�$�H��{�����Γ.��W�UxhI�9�15�O=��hIOb������PI�a�����	�d̶f]@�$�{��ZA$M���A=��0�H�L
��D@$@��E&�s)19y�$D�;�MA$_�|��$�H���q5�O���hI�:���o� 	�&蛱f4kY�Ma��.9zn������h�[��FcWfWy�NA$�{�	#�Z��g���H'�y�$�H��{��@$@7�W"&Kr�b�D`_����H'���hI�7��PI�k@$@&���iJ	��r�ȂA;�{�	 �&���j	 ��`��^�cs|�
RR�)9nS@7�y��,3��=��QUP	A(C�J�.��7p�T��.��D�(-�/8��G�D�̔%3-P������u߾����n�p�j�R㵶�\z�$�s���P�m���qh���v�w}��?Lm��C3P����a�J��ˡ��~��y�0r�0�X�;��M&�SfZqW�����:�\u���HlJA�����8&�y�X�qW�qX'4�Ô�)�+��� {{��7�:�� �o�cO�2I!$�H�J�(���T�����b���a�'��*���5��4SĀ��$=��@�|3	wK,VU% �U��(O�@aPTp*��QT9		0�
G����Ab�@$T� P���Ŋ 1`�`"� � ܔ�h�B@ �RSp� ���&@bA$@��[E�B	b�S�PE� R������:�"b�@""<�� c'���5Z?Ċ���}��� Q{!?���מ��T?�'���*	��A?#���p�"�a��4��*���%���P+��� �PO����"` ~��!����I$�          ��            $�I$�H2�I$�T`��oHzqPH}����b��?�<T�[�l�=����|���?������C����A�,}� �����P'�!�'ѯ�O���k����B��r�����q�?��f�>�h?�C��2B2D�BFI	$�_� " �?�_�����6B�`�=���bg�O�h�����Z��f���y@C���'�C�?l��B!�o����'�3���U%n�� �EREP	D# D �DE	 	$ FDB0P�dBD�VE$@	BDT�AY �%P*SDY 	VE�I	@�@$@�	 $�Ea!a@$ �I�PXAU�EAA$E$E�EdD!�e)D@�	dFa$c$?y��2BB###� 2!#"A� �B$RB)$$Y@�PC�� W��1�N�C�``~�6%�!���?G�P@z�6�����d?3���}�� �o���x?y�\��k��?�����~���"���*X���� ��?bc�vC�?�����>?��������O�?��l�������@DA�?#���~��?��'�~��4C���~�`A?R����dO�@DA�y�	����ZO�`��4J�����v��~����~4"" ������,�%!��t|*� Җ:��O�F���UP��YH	A ?Ƞ8)�G��!���M����xp�����)�����?���?��"��ϰ|A���������|���-�����?)���'�0��J����O� " ��)�#����H��@DA��*�A����|K���O������&���4�!�$���|�'�_�@?G��_]��}���%6�S�"������	#���m��W�CG�t��� ?��ؾ&�>��&��"'��c�?# D�������a��P�����D��������6h���k�p�F?���?b��â���]��BA/�M�