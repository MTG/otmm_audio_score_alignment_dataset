BZh91AY&SYs��� �߀Px�����?���P�����6x-�7;��$H��h��Si1��2Fj�	i�      I��5 Ѡ=!�  M�SҏSM6��4�  � E4� �S      �E�h�$��X�[Ud����
D�)��l�C�2E
L��t�6wa�Q��L��{Hi�Yv��8�
����m�RHO��9!(MU,��UQ�LHS �زH��m��N1V�gB�]� ��!4���w�>yj�&�`�DC걘m�!�gy��.6�[�k���T"�BT�r�W�.�����q���(��/5�F�.iP�gTA��1"ce�l���N��AM�@�Α����y���Dcv��B˭Fåk��)B[+.YRɹ�a���{4��W�w���3�z��ȄP䃛�{Z��\̍<��?.Ji8SZ�9���˜@�m���f�F/�ľɽB$$ @ԣ4����"b�9p�>����ezb�/H���f��	�Qb�1��eܾ��^�d��)S	6��X�7D�ȗ�vz�$��,��fs+��l�@�ӻa�nr��qBA'�I$��FI6E�X/�*C�sXع5ր�ɕ�Y���Q&�jd�bItRҐ�E���u�ܘ2�ר͛f� N���|�z�	羭~Ym��S/��3]��l��4?>�K�^�G�>�R����4d&�����Ƿ�|֎h�"XS�1ϭqw�k��q$�@jd�3.�?ďr��T�!��?��!a���`gП�HS{
�0�f$;'�X�QrAv.�B��X�g�t�g~j�,7�S<����VĠ^��˾�[���UP!0�	V0�@�+��E�S慠��F!�ⳌHU@C�K��SƊ��)��&&�ǆ�.���;�հ*5XE�(l���cR�وJ�Q��y�f�y������r�V�)�l�<P%{88�}p먅��>�8���� ��|Q�6]�#?	iزHJ˦ �[.��	%�W1Q1e��7�� �4�o�h0V[�Ւ��P`�	����L%&l�0.b��۳L�!e��Q��$�V�KRv�g�׉�w�( �.wkvn6���À�GY^�,`;���B��_̋П5�qY@�H�$f	1�C�,s���ɿ�d�eʦP��MW�$)�����"2v3ɦ4Ma8	O�E�r*On켬"ͭZYRG��"��+�l�Q�*ډ�7(K�_�y�dT��A������;�����.�p� ��d