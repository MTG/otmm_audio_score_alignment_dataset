BZh91AY&SY�M��«_�pp��b� ����af_ �
  $   J@ 	 �  � 
  �   O�I( _�(�� (  DTI
@R�@)U ��*�I)@ ���D@(��UB�AT� Pp   �
  A@�14 s�N�:�Mzn-.�R� Jd�w��\�W�'J���2����z�  )N tN� uv�.3��Z:[W��k���D�Y`)LN�P�j���:� �@    M�^յr����؜�]����Y���=K���z�q��f��t�r�T gU{sn���� �嗯]��� ,���֗.,�n����U� ;�,�UX�u[��-ǹK� 8�  �  �` '��qnR��M�t���H�� �/MŻVrݫ.n����v� t�Rťs����6���ͯm���ܽm�wM.m_Zr�vrw���z���w�k�;�x�WN]ڭ� �� �  *�d 篙��t�T������m�p *Y:�\Z�w/&�mŕ,>�ޖ���[��| r�j���OWj� ;r�-�e�ڼ�<��NN�m��=Ը�����yj��g//V�    @� 4>}Jͼ���M�\M]o��^[� ޒ�k�.Mz�o6�z��iq���=.-ҷ7K� oo�ί}�����{Ҝڥb�mqi|����\ ����o-���q�w��yK��      ��56ҪR��h&h� G�jg�0��eR��ɠb ���M ���R�@�4   4 "{J����     ��$�R�P� �`   A
B�LMM�B'��G���P��O�??��/����������}{���* ����n�PWh�"�@PW�� ����TUo�9b
����������O�(�����/����'��0jK3(�!+r0���(KO�-k�?�8w���G�k��7%U53�{����a4��R@P�bJS��-2R��0����%��(&u.��5ZC 0��BRm2;�����M����7&��������!(JV�"�Ñ���\uaR[�h��:��ٓ��A��A&�����GTr�䡊�C_g�eT;>r�
L�%.F�d4'P�:֐�%��%�F�w�Ǯ�GZ���#75���k����IF����n0��'F�����X�5�5k�ߛ9��%߹�k���%�,�8� �ѫ-����Yî]�qvc+�\VK�T� q�9����R�'2�-㋑�sX��o=P������kS�zjsA�H�7:XdE[��i����f�٭�5������v�!5�%��D�� 0�p9.9�s9��2�n���F۝ws]��}�;��vcc���5EA�f.�tI�Nf���w'S��t���uͶf�4Fjq��ֱ��Bְ��Ա��;w���3{�$��$�F�zy	��P�&��\:�Z��N���#V��z�!��5&Fd%`����#&�3#NÛ�@p���'q�{������㠇�Hk:�);$����1�sdkf�1,�ѷA����(����#�͛�k��7�V��`Js��cs����tTmh*�0;�a��f�F��E��V&[��2p����d�����ή����at9���c2Ӡ��2C2g,C#$R�()��&S$�����(4�dDcF�i*7Y�r��~/'�9���vopa��`i��Y�9Ru&{&du�tZΎZ��;�E�t�ox���X�9!j�t�y���f���:�F�w��xC���8X�w&',�M2�8�	����J�g$ĩ4����d����փn�A����wl-m�8��έ]�:��V���3y͛��r6q��`e$f�ր���V>����kINFF����Č��G#�\����c#���t�7q�vnM�����ՈdGa� �޲{���4�:��)#4�����N��s�u�6p/ ��WE�;�w���5f��Մh.�@fkT���:3���Y�7�)éq�pu�p�##*��7�jd�J ���;�!���+Y�Z��"l�"��Gzz��6o�泇\F�yf�	#��� �a&�BV0��r�:w���r��{��Z0���0<�j05͞]>�xjֳ�����"۫8�[�e;��v\��.t�vG])EJ���]n�_��ev��R�ma�D�=�:`�Nf	�0��J��|w�/�u��O�u��ԫ�)9,,q�����_R�{�U*��S���v���g2η�;:<Å�^�.����7ˆhј��"�NL�4g3�wY���5q�f�((舌��5ܚ�A��.�F�Z���8OO��o�z5�8�t�8� d-1�Ն���è8���yם��1Ffh&cX`�b��l�,%��8�5h"r2	�J�I���f�3z���`S���Dd8&A��j�C��N��0�����j�4ƣ4T�E�J�lWw�G�:�+뎜T�T���]�A���kN�7�'%�#2��cb�]�"��!98kg]��l1�P�4A���$����Q�`�UR��`X8���^vf��#���dw�u�Qu���h�ܒ�����gy��8z,(8@U�ce�͚z�Gu"�i��;��;������ov0��t�5̀�\rq# ݢ7j5g�&����4 8u�]�%'M�`�Hs7��.i�E�Hփ�ގ�	b�Q�T'r�C��ӊ��eU#�X�]�ç#P�N�8`_�]�Mй��h2524&&h0r���u<�1d'�u�)8����i�1��	X���5� ۨJ��&�,���l�kA��	BS���d`��=�5��3~����[I�;u	BPHA'@A2ywu�zN�o�ѷXh�V:�uk[z�]��� 
R�����q�)M��ث�ڞ��:ӽ�'F����.\6q��M&͎Od`�:�z�sU��Xr��,u!��M`hr�#M���7�kC9'w��9!�!���,�Ɂ�Ɏ�Bw����:�s�Q�iq���y�d'S��po��h�d��A��r��S8�:�q�C��h���V�o���jqѳz�Fm��ۤ�()�'Ǩ�.dx��g9��g� ԝ�l�K#��%	`�b�;�3���5ӝh*�H��-FJ���(=�O	ˣ �cE,e@T��ȓ	�j����aCN�0a�0`�����	��Wd�<��i���8�)N3�@xe��ձ�12A�,��I�κ�w�4A��8�t3�׏q�����%�-�'5�0j�e��F��:0�7�լ��N�C3b���u�53m��2�a�#2�20сޜX�Pd`A��da�6�YVN>��vd�19bh�z�4Ns�:�]�]��z�}����Zr2��M��`XDdƲ0���t�`�'I�/X6	C�:71޶lk#&�c�1MLs3Hnqr��4���f&�����j0*�+��ľ����8�ڑ�TOſ)e[>t��/���{�TU<Ԯ�RZ�K��5�	ֱ��nt��f�Q��r�8�C��ޘ8fV΋z�}��߭p���k�)�I�Sܣ��)�WG.�O�N:����U��㯪�*+G-�5�sg3��t\�3<�F��4�>f42ă,�b��j'!� 24�i�u��A�#A�ђd1���1�I�I����у��֬�oe�З^��}���p�=F�-n�2Lc�c��Lc,Xܼ�o�r32Sّk5�v���u�84�IK���c<�n�a�4s'#
���뷁�f��zl�љQ�"Dʢ(H�sy�:d	ّ��eY֜��h�6�w�Ӛ6��lģ#{5�9��<�oU'(���9T99�I���.׺W�\���gN��2��04����#��	֞��5��N�g�6��%	By	�`�3��}g���Y�6s������S�NBX��A��Xh*�0A!8SM$R8@`��k��0��Jħ���j8jM�:�Θ���6r�N��8tѫdo0�[3�� �#5���.hrr7L�:#�����
4k�����Y&S���Վ�P�˧�f��j	BQ+���3��5�-��z:�9��[�����A���Fl0w	m12�А%�̡�8�δ�NA���	40�4f�;.���!(�#(��90�85���d��X4�R��h*�	q|��}H�:J}��(�u��F�r8�D�P`l�Ȥ�'s���Ç{��^w�����=5bEn0�2��C-�F@e�8=XJ�"��I�Ō�)�p�̘���%۽�4�����e�5j-BX	F�`�%:!)v���D��'��L�BQ�1@a����!;�N��Q���ܙ�h�G��Ӱ�:'y�J7Dhի{Kre>��	@o��f��Z�uk�k^�۸�::�g}A�cQ�:�	BV�ޥ�-''Q���l�x���s��=��XL��HD�8Ҏ��a�R�bYj4��r2Lc/XrF`��Xi(�3A���-A�h�9�(rC:��FN��	Bn��){7��0����BR�<�LYib섬%�3�{�b2[��z1*�dEhՆ�C��\l�kfs'��c�hц���2�l#F��h���f����ӣF8F�e����g�� �K=���BX��6up���xa%����@e�t:�'���F;ML�kQ���h ֧p�f�ǾrL�����p�ê<v��f.��:\� ��[������&���;�a��w�5�G|y�~����=TS�N�R���՗D��������8�U�r	�L����K㷉��軻{v퐮��>��os���'N�4r�ZMjN�	Z���F�]�pA�qpE*pn��ή�*��PR�	=�sF��UV�L���Fv������V����1�5dfTG
JO�S,N�E*�}A��Q҃�I�n�()�\R���$:T�_kn�q�֣g6�ӣD��N�F��z�A�O!7��Z\������S�)BQ��](W�u|��(�N2�!��JNDd �u9.)��h�#,&s30-o�:�͞O���2MDn�1�J�e&���9�C�����f�#����4Y:ͻ�:-!�e:�!+L���w	BW5��ӿ3�[���(ܹ	���A���D��y� 2�4j�n��ѳvum���hլ2��,:-0�X�70��გtNF��C��9�����P7	HfXÐ{Ue�nLL�� ����G'�7����u���]NI$�IYv�	�� $  �  -�(��E� pm�I   n��f�u���HR���$��Iΐ�m���Yr)|�R��a�n��(��j!v㝕YV�gʇ��w��t�-�jڐ�f�8�M\��ϦW毭���������� �+�6���� H��\�QB�Y2���!i��4��� m��M����!�n86�6mm�K(����Q�Jꣂ^���nP�ۭܶ��� %��r��F�UW<���UTp �ͷ2�A\��m\t,ƞ
����ꪥmY<Up
�K�j�ꗖ�j僉V�@h�
�V_�����u����Hm��[Vԅ�UTWUl*��.&Z�Tb���v�z����l{e�a� �i H!�I�ɯ]�f݂@�  ��@�am ��kl�����}�-�����m� pH����@ 	eY�`m�`k6��R�UK�UP
�/*n�� �`?d�m�� ְ �D� r��b�6� ��Y�� �.��4�7h��� �e&I�V�e[B�I���� ;  m��`�6��`ㄎm��l�� �i"�m��8a�MͶ�4P 8�f��5�3���H �XXa�� ���`l�S`��m m�`�m��t��)@-���#&9o^�`��-�b���` δ�ݱm-����a����  �C����W�It�3mŴ���]U��M�P ��[$��cl�*�`�UK� ?[W<�2*�J���V�����NT
���D�On���Rts�[Ү���$�a��E6h ىv��6ۂ@l  6֒M�2v)#m��> �m�rdv�q'n�eY�����k&k37j�#!� :��R��H� ٶ  ^��ZKbIdk�l䈸:\1'�ݺ1�h���T��R�]9Wu\� Ȗ�i�mA�V v�a	;�Y)�n�v]BBd�s��r��-��� $��[u�t��[xm��ꪬ$-�TY�]ŞL&�Uպ��o0H�Nk���m� [A�kjݭ��k�ЯT�Vi�B�ڵ�
ZU�X+���]P#@�[N�Bu[T���U����*�UU ,kDk�lѶ�`V�+)�BU�j���e��0
����*�,EL�۬�L�4ےH�ޒY@p�m���M��iѻl�ӭ�A���(�i{Mŷ�8l� e�Y����_^������f@��i��Ŵͤ�����oˠ)!�;[E$7P-��ղ��` 5��Ŵ��6�u( "��v�B��g]+�j�����e��� 6�m�    �l'M���u��m�m�!&�t����i2I� -�b�ņ lֳE�&� �!#m"�+�@]Ҁ�s��eP*��A��I�[ͪ�K7�	 -��m� X`��[�%�bc��dup j�P  �fض�h�I�f� �\$	  6��u�I���p='K\F�h�r��ck� H ��Jjj����5m*�n��m�	����e��W6 6�k��!y{c��0��@�R�u��1Zx�w[�,N��v�7��#n�w:�j�&��	�q��Y�h�N�cr��@5k��U],�ׄ�d
���#���>E��U �v�*��o�d�>�<���
X����=�Mm H H �qHN0�UQ�/UT���rH� 
�[F@�i�w���@r�UU �s��T�Ү�`��� I&̋h�MuM��M!�$6ضJI��kn���c�iyp6݊�\�8�&�h�� )M���g�'�5�v�m� c���` �[��l [JW�h��
[h��	6�ݶ����j٭o�� .��  ��h��g� �-�$p�m��he6m��2)f�'7�o�m[s�d� HH����Qm�k@ A��ְd ���l*���கh�(=J�-�� m�m�l�d���/]fX����$��	~�n���/JU�U������ 2�8�<���
@x  ΋{:���rGM�p�g#��t�_R�����u*�M�@�-6��gYx{\��ϛ������8�L�ݥ�.�mr��I+��L����A{t�Uj��'@ �jP-�U��%����|�6 kob@I�ꮒA�tq��$��$$:��]j�m�Y-�hڳli[uV�$Ŵ�P8�`靀�:�-i2�6�M��Z���ҰZE� �M&-�/F�i�m�V
�J�p
�J�0  ��@��-�k���� t�ź�ۛfZ��[@����gK:Mz�;m��$ְm��ճ��n��v�K���jm��{cTn��y�d�g���n�jvZ��Q� [m�� l  ��[x�(�r�J�u��ԫUJ��l���n���U�ӛ�E���[T�� �����z��d�*T�UUU<�P
��ؒI5�b�E�@�N$��\��p;,�R���e���)V���Z����k]�9�mU�LbE7^��nӦ�y6� m� �ݶ�m���X�Uު�m�` �6�`�m��-���n� >��b��H[R���f۰�ݻe� �[[k�l m����l8��cv�kk�o��>$l�� T 	�j�VUU���m�)$�0`鶨��l���v ]6 �Ckj�H *��H�!0U���m�$m�lH�jC�-��wf��nm����� "Z�`n���-�p�޴8&��  ۯ6��0��J  ���a�m��n��nٶ[E�$ � �` @�6�e۶Ѷ� �6�A��@HVٷ]�;�`�^g��HàX ���)n��F�Ye�@��PH[@[@ �$pX�T�@*�UV^L��� � !���� m���A���� 	 ⪩vZ��G*�AØV�NݦY[�*�UU�\�*�n�9j��/0 �l 8�`A�$h�m��H�� � �b@	  $� $l h 6��D��r@�9$�6�d�p,�S+U@UH\��-�Vԋiyqt�ms� 8���f����H,]�@v�V� WT��Һv��J��GjA
U�6����Z7Y���L�0#s�[h    ��N5�-��   6ؑӠ�l 8-�&�rޡ���  h�`H HH�����E��[+������p�  '@ X` $ )V���Ѯ�MPt�������m�հf�Hm��mڐ6�#-��$�Z�5�J,v�� )^��eeMt�m�cH�
�
�*^Z	-�-��'=�-Iv�:� $���4��l -��A�� �� $ ���i�im&�� kV�	Žm�M��n���h��� � 	  �j�eZU�+���A�� �-� � 6�6ض�-�   6Ͱh6ۛvi5�l� �i��鲔 KX�#��"�R�R�&ݴΜ��Uf(��7PUTHu� t� 88m��֛lH����z��I�,��m�Ҕ-�6i-�h  [n�Yp [N  ��(�<���ڨ���e�U4S�h�G5ؖ�m�䍶��q� *��H�UU�P=��a#�4��9�:\�I8m��vQ�W*�mU�)@v�-���&͵y��z�6ٶm���۶�L�	-�a�  �l�m6������Z$�v�IwT�RC� @۴�    kY���Hp  m��m� �f��h ��A�� �n�Hl� ڶ  �`p   m� ��Ŵ �� �mm� �A�nݲ����Z��$m   � �@h v��m  ���k��  ���jt���M��
َ����[U\�ɦ���lA�3m��E�P	l���hM'`�k�{n� �@A��m��-�  HA��I����UFD�Tm��kX� ֆ�UJ��z��m\ʻCm��� �f�ie     ٙ�U�P�MUJ���R� ���Z�-8U��c�@��mUU, m�6�H���]WA'pmT�~�mHZl	 I��(���HXkk�m�퀶�&�   ��m���m�nؑ"ėi3�[u��l �m8 ��HH#���m�:�mp4P�$m6蹀��m,��ier�U�@WP
�����]��i�ְ-�o�봛�-�J���	հ�d��Z���+3i�I��%�  � ��'Yլ�0�y��7����������
��s�����?���_�>z�������"����������!^��	Tz�4*��_؂
8��x�U[�B�x u������	:?��l���X/�@��P�H���)vS�=*��;P��׀(ly�z�� �F�z�T"Vd�&U�:*�x2��"#ત��;@�x�����U� '����N��
@��t�h:<B@ P�x�j��BK�@U�}@N	ؾ� �8'�
/G�A��
q@x������"b(��vih@���"�/���<������}�Te�Te��"���S�����������h���Q�=�AWa�}$�"����v"QU�h�Ą$2b�8ؘ#�+$�M$�	 0H��)PRH��5%%a!4Q��.1�b`�D� ���؈mp{š�����A�T6s�B'H*���	��ED�� Ę�����4�'G� U_�?�ݿ������?�Z�����\P�G��@�Rbba��������zw��W~�ߥ�sn�Xש�;;e�x�ڧ��.^�S�s�*�ص�[V��/	���=Ȏ�]i�O5xYa���z:��\�����Μ�Mr�!�̶L��e��v	Y�v�΅y�@�ql<pإ����I�AZѰ�Rs����=�yvZ��m<�W9�����V65m�F��z	�%��=��-8V�dur]w"��_wZ�����lv�V��$��6A��Y:R��j�����ҝ�]�Y��,�"(�UW�\baCƣ��YFW��c�j�:1�ӎܜy6G3�@pl[Z��t�h
�)T���d&�s%@L&̌V�ʵ�<I �Fڹn�ђ�z�Α��:a�ܧgی��֧ &^+����ûn���c�Z����&�l�ѮR�Ip�&���I&�b�qe"����3�"YU�=*�&��Y�ђ���Pⶬ��¶�����E�b0��ʨ-u��h�ZA�M@���U�Aة�g��:J�G�&v�[Y�Bq�] �cJ\�*Γ�U�U� sI��0T譎���Z��4�miun�`1�<��۫iyN�8̔�����xz�v�+utt��mu)U=m0�>����l+
�qs!*��z�M�� ��lT���(L<k��4'
U-�#���n��KV��!�@Ym�����,�Sd=�nt0��jK�zɅ�@J��\�ƅC��#�)Rē˧7(�5�����lR��jl�8�3�-���'E���J�#�[A2n9j�6�%n�;n�mm�Gk5�E�F�ZH���t��mIL��s��G[0�*�5�����u��G3�u�<�4��d��%6��Td�s���aT&Si�yjX3%�)��Ve�M�V�9��e�rJ6�ޤ��Ҩ��Ѱ��٩�����`�K����ڣhD:[d��Gd,`�\WPQZ�%ʄ��n1=�)�h�f�]����I8���[���ո��n�Z���^�'+�	�%VRKy�����#��U�h �<=@�C΀_d|�f��M��Bk�y�(�fȷh���l]��u�kfD��Qm�һT�z��q�!��Xms���\�;t�DdPKۋ���:�v:�qP�p����/�%М���۞��;\\�td_$�X�i��%�K�uY���Q���E������`8+=�ql�م��7^�WC0#���k�1�{l�tQ��䉗�{$��M�#)�0K�s#*����7��w}�w���g'�wsܼ/�|g�����G�
pd�(7N�lj��[n*���9��{�8~~�<��vW�X�)H҅��� ^�x���O�V�V� ��n�IEJi��,�����c�>�L,>�K�x��K�V��T��� S�U�{�� �^ �5�7M`��!�#����0���,�����c�;_B��eȕ)YۓB���:t�Y�FK�t�4gv��8wg�d�@�"�
�C�$����,�����c�>�L,�ƛ���#j�r(���Ʌ����>Us���y���l��3�d�>���̐�B!Q � �ܫ �+F /r�ܭB�b�r�q����a{��s��o'x'l�qG�듬ҡ��`���(P���g��`}�X��;�d�����&q���I)'*3�����v9�b�y��9�<n�C��y��	ȃ���E)T�������0�1}�v�Ʌ�g��`{�� [��#N/�V�V� ^�x�Z1̞eH:"��H�StG��٥�g��eUU}\&T�@��=߷*��y�r���G�1EB�ʒHX��,��������0���m�x㑥J;����ܭ*�8�Z0�+�o���o�;���Z�L!��W�Ѥ}���F����Vz
�h���{��n���Z1��Wv`����h�\� �+F��e�Q���6�$�+�d�� M;�9;fʹN�ЉDT\M�L�Uv`.W�{��2�'8f�,��*X袢��SHJI`}�r�=מ�*��w��� �N�B��d�;����T��i���?)�=�р�^�V� �{�\�EFu�Oh�Gj�xs�m�u�v.��Mv�Y��L`\;��V���Q��⏶��h�\� �+FʹN���QAP�r����K�d���?b�>�L.�<�䓤��#j�RTrK�Z0U�pq��'l�Ӽ�*���HD((ܐ�=�ج�� �{%���a`z�2�8��q��9.� �+F �SN�Nـ%\� ���)w�3 �*\�M��*J�^;y�J8+m� ���H"ʛi��T,��%�L�vm�Gh�3(��Ё��:�<*�,�q��=N6
��
�BR�mȓۉ�t��� �k��l.7m���H��'d�������\𘋲Z�ܲ\��Qr��vyNm��ظύ�[vr�/���3���}k/Pv�T�Ṇ�4���5�>�؂��R�^-�)7]������x��F�pY�L��/3���O\}<�����^��,Ņ:W�s�$V���ČQP��������0�3�X{&�{ʖ:(��*���X{-�"&F�9�9;f %����?R�aR���1����a`�����0�>ƒ�,r�StԊ��'��ӼܭU�p�N���
�*I!`�����0�3b�>�L,�s�����bRT$\S�Lf���p��t�P;%úg-jK��nG�Eɲ�I҉��Q��ٳK3��d��33%��,��d��
%o{�W���nzz4P��&�5��`��`}�^�[�pq18ʫ�����`\� �+F �Z,�aK�R���M��Xo+�In�x'l��S�{�� =��*)J�4����Ʌ�������0��d�1W�c�'Q	
)r"���c����{U7+1�4��8��m�㭘�/���EHӅ�������0��d�>�L,�I�6�����V� K���h��U�w}RpVG:T�E`��`}�Yڮr��R1d�`}瘬^𓧎6�(5e����h��U�{�)��K�YK��	$"JHX���u%8 �+�=�рwD
b����1�WB�x���{��^:�<�h�� 57/V��t
#�q18��#�;�<�`	r�ܭ�ʰ�J)T�q7t]LMUw8 �+�=�р)\� �R�`W��c�����4����Ʌ��r��IN %��9)��$��EHӅ��=����1Xg�Xs��!�	y���ʻ;�W�(��(E7C��y�+k�[���{6i`b�c�>����̧I8H:���s\�3��̝�y�N��!&��5�v�(8�d��G:T�E`��`}�X��������Btc��JN˼ܭ�ʰr�`\� �J��d��$��1g��{&���Ʌ���ˁ�	�m�7.� �+F �r�ܭ�ʰwEX�TJQJ�&��,Y�v�W*�{Y`9x�}�����U�Rm:������,�cb0�N#h)��n(ی��n�<y�7p�d|�2�2����f���`7)��wX��]��m�5`�v��tf,�f��>�H|��n�mѸM�ݹ9kl;��qA����<����Bt�(���7�욜!s)�!�C[�^�]gd%�aӵl��u�;Pj�Hv�n����Yyj�c�	8��AT)*�>���W*t꾪�t !Z;r)�:����Q�[�]���r6�w[
�Q^��幎�۷S�� )�m���f �r��IN �r����`�L�.���>Z�d{�)�%�#ܩd$��!UM�$UAWy�J~Ir��*G33�u�q#��(��R�r.fg���cÞ��˯W���y�RN����@jH;��r�}��Y�J~Ĺd{�T������T��f�(����78�v������Cf�5F��ILMSt�$��$������,����]}�xs�Ͻ� ��i�6ܺ������(xT�%4�@�f���B�R���`%%&�E��Q)M
l�T���z��k������~y�X�TJQJ�&�$\��e��Ǉ=ｗ_yf.g�ب�E#Ji$����������,����]{
�aMQB"*QR4��w�d{�)���T��C��L.�-�����EM�e�vB�[Y;7���#��"��£jP�lrNױn�^g���cß{�e׽ďP�GIJ�HG}�ί���z��u}�DB�[mL��mQ'"r]{5��w�e����WNW+��ĂK<��!��zS�df���b$)� ����������HdD]tlt�,Oz�� �L��ftA4�JX&$������0" J ��	5��n�%'�Ę$w���RC�!#DT�BE��c!A��DF�������]��oiqp�h�Pnq��D��y�t�@��&D�
^�+i��@PD��0��ֱi"(�4TAT4%P��BP��ZKX�Xf��-!h"hr
Cb[$����9R8����ڝ�*z���!H�� owZ�;a^�h4D@0��x
B�;]�JZ8Tt��~0@v+�*v"#��{Щ�o�H���>���b!� mU��@%7����)H�ws6�9�r�Kig6BI�R�w�@
O{�=�Cԥ)�o�R��}�pz��=�\R���o�b ���Jܷ\��Ps��ٷ�)TE:��~��)Jy���┥'�����R���F��9fZϷ�zS;n.ͷ>tϬ�s�v������\t��v���������5�] �[�{��������R������)JR{�y��Qz��<���qJR���F���f�33{��)Jy����-)I�y�hz��<���qJR���~��$JҞ��h�.dl��Y��R�����ߴ=JR�{����*Ru�����!B�>3�"B��J�e��[���R������┥'_y���)O=�\R��D��(���
�	���)I����=JR���>3�k7fkv��o�R�������ܥ	ت /�~��_��~��^��ݩ�{��8��p�~�d��%��c� d���M��N��xe�U��W8K��w�}��P>e��o5�淾�JS�~���)=�<��R�����8�4�'_y�����qm,��I$I qI�(9�V}�{���B��߾��):��~��)Jy���⟘  �JO������̳[ֳ[ՙ�o��(N���ߺ┥'����EA�<���qJR�ߗ�]s�9A�Va�V��)E)D4ۗĤ�����R������)JR{�y���)Q|���)JO�>��F���f�33{��)Jy���┥��>�=����JS߿~����'����JSϾ�a͛���o{� �������rd�P�����OMe�f����am,c�q�,U�gF��D�N��.zs̎v��;�r6��S�=X^yC��QG��c�Td�Ү��գ��kE=qէ�,Gj2Mi�� �O7 Y�h�r�����l�/M���1FtiW&N�E)?����d�vm�T����i�c1�kѝڝźÞЛr��j�i��㻻�w���i�8��]���B�V�ێM��t�y���M���gV��47q����벝w/m��u۩┥'�g�~��)Jy���┥B��}IY�!{؄!ZƁɪ>ֳe��[���R������ R��o���Ȅc�� �A>�c�ΕUA�ViMijqҎ�FI$/��R�����R���k߳�S�
29B~�{J,�A��i؄!6䜒~���-��{�k{��)H���~�)J,�}��Y�!c�3�"!+~���)Jx��z��[�����խky�)JO{�=�Cԥ������qJR�}���,�A��9�B��6É���.|:�a���*��N�V�;&#ΐi���3���{����6+p4���[懩JS߽���):��~��)J{���8��)I�y�hz��>���GR�R�CNH����(9]�f�s�t�O$T6��!�DZS�S��B��K�J,�A��9�BԢT rR�������0���6k337�R��ߵ��┥'���~��CH�@�䧿k߳�R�����pz��=�>�5�Y����[�)B�ҽ��r�Ȅc�� �A
���!)}�^��R������5���k6Yֳ|�0z��=�^��R���~��R���k߳�R��{���J}����_��Y^A�Ms;I�U�g��=m�Z�v��uQ�����\��fF��w���q���[ћӣz��oy�)JN����R��7=�A��ՎR�
,�A��s�)JO�+��}�h���ְ�[��v����JS����8�!JRy����)O~��g�):��~��-)�K9�IH܊��r�����U��R�����)Og�u��rA�㳴�R����R���kﳊR�W=[�؁HRN(��n��Nr������� ���B��ި�!B{Og�P�'���~��R���_gַhٛ�I���s�؄![x��Ȅ
#c�)JR{����)O~׿g�)�����oÿ����{۪
��+v��;sŌ�ǖ��z��;V�J(�����;tF�V�7�r��ߵ��qJR��|׿`�)J{����4�'_}���)O~��aE����[�)JR{�����!��~��)JRw��߸=JR�u�{
!+M��T�uS�H��y�s�JS߽���):��~��#L,t��!B^�V9QdB��G3�~�oFoN������R���߽��ԥ)����┥'���~��R���0>L  6�k��┥'^��Y�3�޵���o{���z��=�_}�R��^�V9QdB���A����G(9��Y�5 ��p$��J�IT�Q�+��)�v�
���:�'p{d^:{?w����$�$��ȯ���(9^�<�\��Pr7�v!BV�}J�"����Ps�̭�؄�@n29��UΜ�R�{�~��PL�����߸=JR�}��)JR{�����T@�+1�4pu)E�$W�Ps����TY�!}���BQ�B���*.R���w��)JO{�����#y���5�R��������)I��߰z��<�^��R������R���G�Lh�;#Z�kw�)=��{�R���߳�R��}��pz��;���qJR�`=����ۛ7�浭l�Þ��tՂG� ��ڵ��O���e�ݻu����1�;)y�y7�H9����Cr��^۔���>�L��l�6܊����Y��6��z&|Z�a�:7C�n�4��Bk^�0h�\�.7�M;�s��3kmð9焸�yywKM������([�tݐ��P���X������Fn,�6���`�zBw���L�2�[m��ޣV����TO���]�|3�k��z@xݢ�m|����9�m�[Iغ0���rl����#�ͅo��m�(w�]�˛��R��k���)JN��߸=JR������)I�k߰z��<��>-MAG�Q����r����w76�9�;���qJR����~��)Jy����s������-Q�D�r9uΜ�������)I�y��hz��<���qJR�����R�����ϝjַ��fV�Z��)JO;Ͻ�Cԥ)���R��w��pz��;���qJR���f�
T�8㈊ܷ\��Ps��ɥ�)K�{��JS�~���)<�75�:s����P4�SJ)H�J�6���r���.��P�e�zu����^sr;}ѫV8:���M7!|�9A��ۛuΊR������)I�y��iz��<�^��R���_~�Z"7�Xl��5�R��~�������IReR0PPؠ�ǂd�&�Ϻ�Cԥ)ߺ��┥'������=�=>��r���k5��R����{���JS�u���(O;��=JR���/���(9]�IڥZڔ"�r��Cԥ y��8�)I�~}��JS�~�������~��)Jx�Ѩq(��2Tr+�(9�W��ۧ�JT�߷��)JO;Ͻ�Cԥ)���┥'�����[7ox���77Lvۘ�=�&2�Ӑ��<�3�v�r<�ݨ������ԟx�Rv��j��~���	� �߹�┥'�g�hz��<�^��AF�����ԥ)﮾2��*�G&B�Uñ"B���ҋ�B�)����qJR��?}��ԥ)߿o���9A\�}���'R��"+r�s�������)JRy�����C����M)�~��R��������Zr��G%)M9"�r�������ԥ)߿o�R��w�{���JS�u���)JN���쵢#{Ն���[��)Jw���┥'������R���{�qJR�����R���^{��	�/<��1�����OX�#���eX�\��5�r���nzݹ�ض�+���)JO;Ͻ�Cԥ)���┥'�����)N��\R����32��J��(E6��ۮt�(9��<�uU����������)O>����)<�75�:s��y-�P�Q��d��W��'�����)N��\R����)�QdB��s؄!{�9$Җs���[��{��=JR������)Iߞk�z��<�^����d$����8~�� ���$�w�y�\�)O��u���-kf�eh���R����5��=JP�g߾��R��y��TY�!}���!B^OHUºr����7����ח=�]�O t����}R��?g�8z�31����~���{Ǟ���)JR}�}��R���}�qJ�A	��ܨ�!B�)�T�K���9S:�k{��)I��}�����;�_}�R����5��=JR�{���JR}߯�f�F��Vʷ�o�ԥ)ߺ��┥'�y����V���w��)JO���=JR�|�}�,�#Zֵ�┿��������)O~����)JO���=JR>{����)\��RF6�V����.�W:s��{�g�(�A��~��)J{�����)I��k�z��?��yؐ����$q4�+�����5����kd���Lo��E	Z��Zu���X��J6��%�w���$9ګ�WR�
C�
����;矷kY�֍k[ѭj.0e�v۹;v�+����2�0hluҡ9��l��Ҙ����7d��1oQ����r}��Ş ��Y݇���v���B���k\t��ѡp�e6�5�0��Rդ32�.�;�.NԩC�/d���/��ʸ�ʛ�����ݥY�fαnv�T���K{�G(��M�Fݢ]��Ó��9Vm:6We���`Y�]�
�{gaIN�y4��8c�ŶĵA�xs��/9͙-�C�[�#�/s��0�b˻��V
�O\1m�`�^-+����*�F��Mڝ��� �6�@UQQ˫kEy5,:����*볘��WL�U��A��@	0v��YN��m۰/����Yy��r<8:�'��\�m�vA�`�Y\��97-�q��/;����1 j�4Oe��=6��V���3�3��a�F�.Q��!�JR�6W���I�g���ky��)N@�<ڍ�3��G/��s�&jpt��l	�Sg��É���[l!���{l=F�7n�|aj��*�1 lR�f꫏n��	��&�`ٕ�'�;��T<lMuƖvvUU�*��%N^����Y㴓Ҝ�RmW,�gl�;���A�U
QԪ˭nm�'O��}���@�x���c*Y�e^U0H����4`�{K�Zl�Y���)A��Aʲ���u���J��A ��e�[�l6��l�7�~�����&��]r�6wWn���WF�5��ū�Wn�e�A���͌7�fI��A�ܻ���9�;��I�Ȭ�7��ti�j�*�<��۬h:��f�4h��.S� U��:���nn�G��y��2��U��ct���ZE�+�2��`e尣t)�,�5 �����Q���5�r�V�I��i���$8���r��hԯ�����t���9�eޤ۩�n�N�@Y^���P���g�Uv�MF5&��{B�Ur�d�2��A�X���]��������*����f�{�v�����?��lt�S�p��E�=p¢��d���k]f���h��޵nH7Q<�9�ۢԹ��3��l�Nv3\X���y�J���M!�St�3��ԑ]M��u[�(���3kf�1�
�Z. �!��������Xz�L\�0ζ	��RA��"N�6���`ܚ��)۴nI{]	��gV���``ճ�D����[j'��F��s��ڨ�J���Fv���>G�{�����8D)��r]�	͏&6x{9���뎸�l�;�5�v�<+�;��\|j	狮�>��o{���׽QdB��|gbD ���nTY	Jy��8�)I�g����������٭�ԥ)�o�r9)I��kvTY�!c���B����TY�����؇M�p@�n�Ps������=JR�{���)JR}�}��R���l���r����f�J��Bq����Cԥ)���┥'�����*!{؄!?K�J,�A��RD4JR8�i���+s۷\��PD/c�;�!'�x�E�"����(9�W�{�St4�&H�r*l�Sp;Z�e��vF�=r�v(��7U��"=:T�A(	��NU�f���k��nu+�כ�`8i�Z�J싈SU��ʾ�_{����T�P+��h@�G�U�*y8�ov�d������&T�EQ[y��r�� k����X繯���hH�t�J�� k����`��Z�;��p�ө'G�F���9;�=�4�7�s_@�=�`n{w��h[KSHt�R(���O��۝̹)��Pv��g�/7e���S�q�):lnS�Cp�7�ۯ�{)���n�$��ǼӠ�qJ�.I5sUste^V�ʛ��7�'l�7�s_RFm~��(��6�q�`~y�v���IJ^I@�s+����Ss�/��*���9��r�6DD����7+7j��Ss�j}��db�
Z*QI��`|��v�y���{w�ٳK��#)hґ�"U8AqnE�s��K1zuˎ,a���˱n�<F=�mҨ�`�l}���=�uX�n��{6i`o��_@�`���H�t�2"'s�>��@�����@�M��=�:4�ҢpNN�f�,��u��M� ���%����⬘*��8tC�y��=����7v��Q��"V��*���E_*�ſ���o��S�Ȅ�nM�e^V�ʛ� �ﾏ�sy�rv��~�}1��1q
���$r���I��[e:���3�vw�L��Wj�C>Ǯ��w{����䈁ԥ#���qX�n��{6i`|��	+�M�@���UT�)S<���tNّ�DD�M:�9Ss�fy��D@db�9@�]�q
j��t:��@�M��.��@���kT�[�M�ۻ}��uX��{�=�4�>����=K�Б(��q%ɮO@�y��6BX��X��ڰ=���ʴ�C*��s�R�f!���o�o3z��ժ�J1��Q��=2�v-<��#�EV֤�<�z�YL�P-�&�%����v�h7�m��筠%U�7�iN��=c5q�ַ/�:�c`Ws�:�5�논nv����{xsu�3�q:�0`�v5����E�2�4���<�sm+Y�u�\�T�Ь��ԕ��(sr+�p���]:�H�*H�fLm[&�N
��Txɛ÷-v���{�{����m�s˻�8����=qF���gy���v�,��i�%�W/�\�/�|o��GJ��9/�{��Ł��n���{�s��=����+l�鱹N
�Uf�M:�9Ss�%����0=��S�*!8��S�-�c�Vg7�'l�<�Z'rȘ�����������.otNـ>��h��;�Sn�Ҥ�	@H�z�f��DD(��:��n�@y����d/��t�l�6*;c�pCsJݺҜ'6�/9f���i��{=V���w|vݎ��v骚� }M:�9Ss�5��h�� �
��U��H���v�-�wvD*P��n�{8΁󧎯R��LKQ���H�t�2(9����w�f��:Mր&���E%@˛&�\��lB���tm=ڰx��Ԕ��݁�i�Ҫ*������p�:Mր&���{�&����7�U��֮|��4dv�^{t]h�7]�vy�0�C����3㊴������՜2�s��|�<|��n�y�u$~�L�i�Ձ�����R�R4���`g�w��r��P�G��tm7�`��(�
��]*JR�@H�znM,��k�꫃��H)�`	I	IA�Ƞl��^����^������v8�5S\:	B�γX<|��7v�"!D=}Ӡ}���i�����m������`���!y7�jـy�N��^M�u!�#յ�]�^����Iom��[�@�k%=��
B����24ݣ.�cO=0tU���otճ �G�}��`�0EDiI��@�ɥ��Y�����}���)�RkӚ��QU!�prB�����[��9UF}����4��׮�$�m�)��}#%㮁�cw`c�3�v!B�!D$�IDZIR������YK�K��7u3UsWX�otճ �v��
w5������*�B�t��H�R7	Elɽ�李!4)�֗oޮC�N�5��E��w}�[��T�A((q�����`g�f���s_a�w`4�"t�����k�@�v���)i��m�g�>��5K
���WȪ�M��`9׵�=�n�W(3ri`{�3W@�cKi�Dt�U�s7u����	�f�Zs����ݬ�ti#�Dj9��@�ɧ@����6�:|ۻ�$�`�r��UU<�X�keI@)NqNVi��H&#8�d���6�.��J�.�+�����u�;��p�֧��.(ɱal�����b\�T�oL�q�G�aX�}Q��ʤW8S�����Z��TF+R���;Y(���P������x6�F�l�\F��LZ��/V�p��gzԛ��o4�1�l�U�m0�.{E�	J6�6��	u�p%��ꎻ�����<v����n8;��N�; $�ۍ���!K���p�������_p�crD��JrB��ߧ�ˠb��`gۻ��W:nM,75��)��n)$���%��P|ۿ�DB��A��?l�˿��\H���uԧ�'"rt�ݻq��<���1��@~�
mֺT�A(	�@�ɥ��l͛ Ǐ�S���X�I�J;DMT՘�i΀��X>otճ ܯf�IEI�($�U|#$��OVk�{F9g�-��̉58�G#a]�:st�QS���	�x4��	�f ����z��[Z%:��I`f��n!B�q&<�:�8��<|��`:4�Ң5�rw�f����ɺ���,���@��m'M��J�)�ـ.v��i��7�jـ�k��m'qHK�] �͖���@M[0�m΀BBp3��e]Ը���ۓ��������Q��]<r�N�N���n�aN���%:�⑤�NN����w�&�����@N��Jb���LM�]7{�&�����@N�����L��I��v8�5S\:��gU^�����ΌO��L��2��0R�1�M��WgiBg���]d�HPR&��o
FN�p(b �<�6�a��H�TjGJ=&�$���6�2Z�AA��%�1������2L�IJ$$�P���h�@�������T���ٶ
���0�D�#� ��� :A�� ��Q�&v����<T<��P��LE���T;Ђ8 ����&����X�P��ڭd�E7C��� ���{�.v��[s�(��F��GN��"�X���@���,�&���H���Xme�ߥH�m�>���ni7�Fׅ�y3�D�����y7Q�})XJ,�Ң5�8����,���@9�y�� �7�L�Qwe�݄�V]ݘ���@9�x�ot��/�� �f�l���q7�\��<|����b"!	D�7�t�����Ou��R�R4���aUU�w۽�^����W�{�>��E�FED��͖�f�iֺT���5�@�l� >���J٠Ӽ>otL	T��H��b���{mu�3�6�1yغSS������v�1������v��n՘ic4�w�'���h�� �8�TEL9.ɒ*��p�i� �7��l�K�|
R�aw3uw2\�� �7��l��u�:-�vk��I*#Qȩ9;�*��l�u�:O7X�7�pˇQ$$�
���,��j�痷]��y��=��tJ�!D$��`�7���8�D�%s�'tlq�#��Ӑ���4�GHl�n����Wf8g�Gk�&���<�W��p#�tg�T���O��î ,V�@*y����[�OK�U�`�*�vzC�']u�W��..�g�<�Tpu��,ܺ�%��uZ$�x:������^Î��38fen����vZ���n�ά�psg��Z��n�-��CW��������>���Hth.Y��]�{�ו#�+�uGRSt��2�g����%+_�����~�vα�@o��6���Q)ԧ�&�q����@�^j�7}3W@���`na�N�ҥQ��&���:�=�s���yOg�o���bb5�P��J)RN+s�5t��V���X�[��T�L�Ȫ�r�'@=�� ����I� �Zs�5�~��3����2��Qv�i��b͸�v�uƽ�4N5:�8#��`=h�jx�x������{�{�9��NtO'Xk��I*#QȩI;�>��Wu|� ��I���]_}���uW��k�7���@��R���!$�P�n+���@��u�?4�@�Rs��)�Dbq7��k����T~�����@3�Ob���]>Ju)�#Iĥ� �7������@=���#����7��x{<:�h��q�y/cu��k�z�<����vR�H��S˧�������tj1	������`o�f��}��u@?&�@�_9��A0g�LL�� �Zs�zy:���@�Rs� ��b_�꒐H���ݮ�}��`n{w��:r��D� �b�eB``B@�)&X�)� )ƻ�^����}��gU|h֣I(��ujI`n{w��<Հ>v��|{��c����.���bf�tu'8C�I΀{���߾몺>��!�Z�y�?0�<.���I���wAd=�KS�g�/a�+�-��N�u���V8U��yZs��� ~M���{�9����)��n)r�@>�l�Up�7vެs�(W!���l�7eW(i)J)�NK~�����U�9ʣ}�5t�f�su��*�F!75{�D}{�9�+Ntܝ�zb>�>�9�۰<�ˤ�v8�*f�=��@��=�� ����I� ����~[�\�6�O9`!0��{&gZ��W]n�Y�u+I&͸9mѻ���k�>��Ti:������u�?&�@���F�~N�́�B�4��r�.R9��9]����1'���@�|{6z��@��C9*��ȩ);�>ך��L��3�5X�n��n�R��R8��T�m�a�)�}{6�{=��݆�P�S���`~���M��$q8+��/f�V�����{=�9�l
p�DQ	G��M��g%<llO-'[gq�tR�m7Xt�ϛA�^Σb�ޮ�l�>N��b�:dq�������Z���8{;q˯X��q��e�u��WNbԯ:t�z퍮���[��W�s�p�Q`�Q���A�5P�l靶qg��Wm�6������ai7����6����mp����%�8���������Όݔ^�j����`9붣����w��n��������6��n�=�ۙm�.�|�ݍ�.6��ګ��{ �n�����qtT�U������<�9�+Nt<�����u���bi������@S�� �����̺��`Ϯ&`����i΀����7���V�P�X�nH��INv�t^ͬ����'8Jӝ�
`®K�������p���t��+Nt=�,���M��c���T���u�Gc5���9��>Ns����*����r���:#QȒ��幮��d�] �f��$��z��է��9\�s�J����t����,��"TD%;��t�s{�>[��|��4��F4�)	�;6��΀��5)�N����{�:��Ҕ���(�cJ8�?s��+�'�v�m=�����XjJL<���3U�)P�5���z��U���T��oO�yOg�g���J"3Jt��	�O�:x�n3������7;�틠t�)�]�=�]���v;^�;m���3@]I� �7��'8jI�tC���.�.¯p�Rs� �����V�6��A��[KP�#�Q�$���3ͻ�>u�zl.�(��%	Q����:���6���6(����IN]��P�D�^�=�����X��==���@�)ѕ��q��6����lNt�Rs�5���i��}	���q�\xu�k��q�K�:8���q˴᜷H̓ts��Ur�w���9����0}�́��s�y��>���DDD+���o��?k�_�R������(�7=���%*Rzu�t��ٰ3Վ{�(�7w��T*�F!1�ށ��;}�5Y�"!$BIH��@כ�`5��] �U��%BN+
�홫�g�j�7<��П,��� �!J��A�07��H#�u�������R�V�$Dj��;v�y��*��-����{i����9�>�q�&yT*��m�ķnz��a��{pj3�M����c�.;��di���	m<�����������Γ���@]I���suN�dn*��k�W��#�l�ˠn=���7{�ԑ��F�%F�1Rm���;�@]I� ���Γ�Jj6��L���%�]<�U��f�z��U��ɚ�ۓj�DB�E#R�p���t����:�Np�������h���f�I� ��:^�!��"&��i��n�!%���兜��$d.�<W��t�ljPT&r�w��>6��a�5��g�ZP��p$u�Ta��q�H�H����rx�-�q0SC��h��Zd��̭���7PHKP� )����4�$3U��v�y��0��H��`twoi�ǣ!)��r�)�Bi!�����H��h
(Sp�O}�U|=<�:�!�\X%Y�����w�4kK�)�$"
��f����n�߮��_����� �����8*���ٛh���	���-�+c�{T�y[�-�-kaÂ��7P��i�t������ru��'SNj5������"gDŻ	y��,�g���.�5/N[e��֧L-�U=�X�$C!��6��Q[E<� '<�lR�f�$�p�,;f����%���ʻ.9$���\��i4*ͺtg9a@�ڸ�R�Q��D�8[��2����6\�K�*�b� \��t8<�l�u��6�.�cWnù؅��b@�� v�:�0ƥ�Y`�ܓ�۞�@��.l�Y�s��;C�a�Kl�C��!J*R���S]u�o4@v�l���V�,�
��g�gr=��ն�%�V.dA���\����7-'��'=��:�Ar[�b:�駜E��50�Si:�FcHX�nR��7=���QP�*V�ٴ�[Y�WC���S���0Ar�����!-	A��pغ:`(5cm�nh�L��8�{h���@i�C���`u�*������Z��5U�VUz�
H�E��C7S��ۤ+@�s��pP���z�ЗK:9���66 ]E-��v�9w&3k\���wf2Q�Oc쪚�b�
�&�j[�� ��Ԇ���$ �q���[[�wT�f��s@U(*�s��-�������)�<�R��8B�T��,��cV���	��t���V���\�����ՠͬ[e�<XZT�H���.h&� �-�x�v�ۓb-:�*�@ �t�,@R�n.�G1�[gWk'6۲��)��[&�<���������ϝ��	�U�[���[s`���n�;>³��vx��������]HI�e��\M�v���Y[�D��iV��g@0MU �U�R��s���X$کT��g��5�uN���UH%&�vFv�<��*�A�ķV[q0)�3��F�#u>�epO,��t��n:���WA��3�t��F�wYm#��8���^���O	��[7��Vk5�fe��s��*�����D��xv���k� �"����@��E4�ҵϧ�3��q�� Gm�f���<�i�����v�G���1�
�l�p�v1�;OSM��'nB�l�:!�9�t�Y�c;��b�+*m���8TC^�l��5�Y�gsF��.�� �,C�N,-�nz��A����I֙z�eq����%����K���έ��1��,�S��X�	�n�>j��h�6��N8Ӹ�ڲ�nǶrn�n㌚�W���{���ޭ����\�G8$-�\*U;�]��1����su���ur�v9�Ƭ�)NV��U�Bm9�廮��d�]<�U��f�z�sR�AB��Jj�8��β��V9��n����I)�7P�/��ۑ%
�����n=���7{�>[���e��6�kkZnt�:%��� ����Ӭ�X�u'8k��b��D��T);�>[���Ē�n����z�� �U)AN��[�����iv�øu��¡x�RƸ;gX�qڵ��N�hY�m����3Վz��I%􇶞�@r���`�d�IN��皯���Um�M��i� �,f���O�As3q77tT��� ���Γ��X����`n��ҝ
�Q�Lnw�\=�p6���Np���s.� ����������X��'8�ozy�>���M��EQT����;��]��p�l	=�n\�NmS��#��YS��"JI۵�=�5X�n��g��7�3W@����i�Ө�H�X�ot�����::Np���6(��L��B��<�U��ɚ�TGJQ��t�=�n�b��.r��2:q�"�>ܙ��{^j�3���C�*�nOߕ��o�R	8��ē�4t���{�.�� m,f�GG��~x�n�E ��WW!������{}����Gsr)ұumGJ��3���$S��rl�ݻ=M�@o3��<����4�S�Tj1	�����W���)#u��`f������s.�"Nȸ�W&k���c�α�MP�"&w���z���X�B�knQ*%9۵�<������nz�4��QP����w.��kKi�M@��GDm������� mZs�9�� ^����tM����a�s�������^!�շ�B�3uۭ�yq�-����D���c��_��� mZs�9�� o��8�KjB9$���qȬܙ�����I�n�K�IDL�v�t�zN<aО(�q���k�j��7}�ށ��U���5t͋JN���⑍(���w7~�V�����s��?8�l�H�ʞQ$�U˰V9��!n����������v�yB�B�	G�]8��k��"m��9K6�`'��M)-]p!��m�t[uB��YM7��.�}zNU�B�y���,�M�¡�h�ar�r�Ð�y��YZ�/l����b4���&��8�P���=u6��]���Wm
tv�Kp;�ɽta��PH���W+)��d�!��ya�<���D��WWEfqE]r�!�Unђ�1rgV�5���6}o�6�!i(F������vwd�f�MN�ؠ��J�:�c�ITI�
R�����w왫�9�� ~I��T���$��]U�Qd]���N�盬���T��t�]�Uč�im?ɨӨ荷�������z8���c�����@���Mӡ:m݁�~�`nzf�ܮs���~Y��?{���@ͧX��#�H��Ȝ���Nt�n���<�`���~m�"V����ǭ�˛cpI�}]q������/	a{��ml?`be�}|~���� ~i���� �Zs�rw,���qH�E#�7���Y^��hK��<�c���uݙ7L�S�$����J� k�9�=<�`�;�>�Ne�J;S(&�]S�:�t���`�=�:y:�59$uS�'P�*Nݮ����6��s�����y{5����@�U��Z�:j�q����k���7.�t�
rq^ƻ�]Ru:�;O�.B�JS��Ө�4�}~���^ͬ6������p8��T\�u\�s����u�1��,����(J�7���ށ��֯�$NG##d����β��|�t�I����J9Ou��O�Ձ�wh��	8���6�΁���i���� �X��ܲ&J
���(���6��<�`	���<�����VQ���j&ө)1��s�m�::��:��y;9��o=���P���Ix+�*�.*fj��t�N��{����v�!̺@�Gc�e�+�ck�">���[�6��<�`�̚ڥ���
�$����`f�oz��]���zt�ik4jt�0�Ur�7��O��@�󬰴�"0P����o]����hأ�Q27N��7]R{����ݮ����ߟ��L�1�RY
)�A s��]�]�ۧ���0p ���Ƌ�m�E�4�uuWu�&���:y��i�����wh���Q��r�y{u��=�:y:�i�hN�1EM����\�� �Ot�N��{����Ś*t%R�I�'z�c�ߟ@{��X�7]Q��׿XN6gj	��n� M�f���� ��v���@�I/�D!(��O�(|�<v1�y��W��1C�;����z�n���V� >ŬnC�՞���i����z"q��&`	�F}7nʆ��Һ�BZ�ʵ@&y;X%Q�u�����a-��^�طZ���=r�kmptF�T;]�l���@v�Hu�5��y�U���Hv1�`S0���#p�'�4O�Ne�xkk��q���&z���Ħ�T7[\�Wʨ�-���GaJ��Y�=&r�҃��q��p����[=n
wSg
lۃ�e���ڥ��I�:��vm=�:y��k�8�$�eM��T\T]MU� �Ot�n���h����x6�$t�&G"�$�@���`	���:y��iT)qwsR9$nG`f�^��ۮ�����/n���jA�$�wg@��� M��O7Xmc4�%�c�'2���1<�Ztg:w;V�6]"a�#Upv�q���n���z�l1Nt]� �Ot�n���h<�`�X��S�F�SI6��@����}�Ur���)I� �OtB�̺��`Ϯ&`&���h<�`	��@���`{u$-�-N&�Ta'l�^�Xi��:y��O�8�$�eO��qR�MW+�?f;�6!(YY�V��t�=>n�1�J��T�T��<�o\,�X�c��w��:�X�C�c3��Nr�M#M��:U#�%$�@���7��Ӡy{u����@ͧF�#NG##e�U�`��4�N��=�=<�`}�6��	���wg@��k�7�}����~@N��_�
V�x�=c���h�"IFY&���c'n����Ũ��������Y�Jd�D��<ӝ�nh�]�����xi�L��O�Å���ٜ�JBI&	 �d`	BHe��" ���f.��OOR �: <6�/��h	���Y��A�����wߚ�]{��?]A���t��@n))H��f��|�����h<�`�
T9��n�b�fI������<f�w7x䷽w"�t2D�F�)���
�
Qs��<	@K�gC�ޗ�.���t�v��q8 v���v��&`&�������{�t�u��B6�ַD*0��t�ݼ�Ot�np���q$�eM��E�E�Uw�>I��M� ��3@=��`m{��i#�Q2I����7=����y�t;�&�$�D;H�TC��;�3ߺ��r�� ܒFF��X�m��:y��$�@�� ��B�EE\��-q��Y�����f\��s�\x��5ƹn�-;ry�Q�%|�)J.�$R@n�vt/7X�������4��*,��q9H��`o�7�8^�vw6�`z|�w�$���ֶ�"yRU32M��
W�Հ?'��"����Ot�+R�@
��RT
G`oٷ�@��u���j������rI6�T��$��.��p�:y��$�@��� ߳oN��P�Tr�^��8�ڨ�a�{)u����ŨJӝ,n���n�	 ^��G!�l�����R��c#�n�S��:��v�3m��q�ʜk��6��̛�C�Ș�h�j9	�z2��jN�c��a`ԗ1��2����K�4\rKل�*�f��r���ɲֹ��B��q���i�[P۱�P���u7��ۚ�ft�:�d�Ӡ�vk�\'\�=[n���}ߟ{��}|��<���n��c�qs�u��W	�mù�����5��s�q�{��J"��57R��v~�ozO7X�x�����p8wR]M�uw�O7X�x�����f��(7uJ��#��F�v����=>n�lB�����m�������imHH��7Q��·�?~v���t�np���+uT��]Wrk�������K3��`o��N����`wk4�n�T�F��r"��nqHk;�ӱ�<'7h��V��v��ήdwݧ��B�b����V��zt���$�@�̒�	��.&`�������[J���*T!(������@�i��M� �I#���4\TYAw�hsw�>I��M� ��3@6�Ec4jn�86���f��e~�8�x� �n��H�e�HE�T\������ɽ� �n��oz*��Mҡꑺ���t@|���ɇ�Wl)u�����]�aJX�n���]����e������j�p��ƀw7x��^�vＶ��R(��Jmݝ �n��{�t�u�jm�h	��EYM�R�JI`{ٛށ���eUr��)0? @$��B)�����k�����x�i��
��HRw@��� �6�4���;�{�y@�5���Jj�H�}����{۲���7��ۮ��Q�޷*'R�SMã����i�n��н�������k��8�:M��4"6�F�S�TpRv��n��i�����o��¡�\�UeU]��=�:y��7��hs�`{Ǒ�i#AQ26E$�@���7�{����=�s`�.�����������7��hsw�w$�A����@M{��ֹU�~fЩ�%"��&�΀{۲���7��ۮ��oN�啩�T��$�&��3����'׎^>�1�srNS�b�ڎ	�ڣ�
h%8ڕ$�����<����v����,����ДH�$�w�O7X�oc@;���'��#�
"�š�$T�PMO �7vՀ}�V�ܷ@����C��]���Ⱥ������ �I������3@6�%X͑R�ԧܖ����^n�����=���X�\IDD�$�ʮ.Q��TU��ED�
��'Sh]p�Լ��ʎ �+e \#���#��j�3�{=���^۷<4��<�����j��y��F��;�g/�V6 z�QĽ4�ŚN���m����-��u��p���"�j;<��i�N:Q�ӝ�\M���yZ��m���X^�����@�H�M@����!0��7'!��A�N=��Ǯ�:�7L{-ې+�zn6sAg��w{�6{{��l�g�+�b����&�ۇ����oD�f3uۭ�
�p�F{Z�
��5��f��ݽ:�n������U+eJm�#�ӑ9���3@;���'�O7Y���&A{�H�Q(��n��g������vj�3����>���`c3���!�\���L��jQ��`d��t����=��`g�RZ�ӠU�$���˛�Sx� �n�I=�?DD}�{�x�W �KiǇͶM���==�g��.G&i��t��[��v�^�;b��<�~�ƀw7x$��<�`Ƥ���m�"S�ty�|��p��G"!(�9����st����L�M%X�tF�S�������/n�6&~{���̭��yzF�s� �4O*n��t�n�M�4�np�G�GӋ3{�=�m�T��9$nG`w7q�u78$��<�`����vg`H.&Y�<C�nܹ�nĎ�<�Hfn.^����,*��}Ө�-�~�~������{�t�u�jo�&+uH��N1�H�ff��y{u���Ӡ{�uX���T�D�I$����u�/�,q
#� ���	
6S���`�1���	J9�87��@��݁� s.�+�\T�M�`	�nt���m��ۮ��IYKS#T���{vtOww��������8�jY�]7[�u�����k����1��<)ۂ;q{�Ū�i�sp�h�:�\]QS���������`	�nt���$
\h*&(ԎN�/n��Ϲ��Sf��?ut[�������f�\�ڒ9%�]� �x�JN��{�z[u����-�R(����tY�����Kn�������s`}�8�JD�Jq�P�q���ށ���`f��]f��F$���$�8ӧPq�1p����˺��{<PSú�E* �N���ڊ���i$���-�vn����u�&������	�Ϯ&`'����!D=����9ǵ�1����^7`wƤ��oS��5Q��@�{���ۻ6�;;�]��t��"űJIT�*)������u���e����wy�=��ѧ9R�D���@r۬7m΀�78m�п��R���T%�
B�(� ~���c��V�:QCx=iM�����}+�I�& d�(@�b�01mݐ�x>�:���=�ZG��I�C����(C �� R D�&��Sh�&���T�(�h"&�f"��("��R �"P( �"�4SC�2�3����P�Еx��Ћ���� ��!��.�=�0�7�<,	
KF��Ѝ2jM�DR��4��*���'V�h�����F�A1�a!�&�M��š)@RT8�G�\T���ZA(��T�$�b;�H
d��a��SՓK���^o3YY��{�����
�X ��7k���#�`�.1���D�������n�Xݶ�Ǥ����m�I6��Trta�9"j�l��"�Z]�l�eZ���]�C^��۩
c�I,�Sۢ�p0�G&t䗱��#K*��#S�U;�3l���䫮[y�6s�e�;'6�B�. �L�h�Waj�g%�)n	��(�۶�J�l�۲���[#ki�j��l��rk�cmRft5�2���*��A�mv)ִqv���j���
���xegH�˗�^��� ��u�<��If9��p筋=/ls�V�U,�k\���vV�B��͝'7[Ҝ��D4��"N$��ݙ�dK$Hq�Yy�y2�M��콱q�c�J�����u�io[K«��zʴ931`�cڭ��X�7i�tl�'Q,��Q��m�iJ$]�Kk�:�t��6��e�����h
x�C[��+�c'Wn1�,ڵ��]�@36�cl�m���uR�I�i��Ɩ��NB�vy�2����&7b�b���N���P7�g��-B8�櫀���'�d�c��s3�f�@.���z@��2]��9�ݣ�r+/�g�q
kkC.zUv��J���s�6��m���kP�d�ab���.�룞�Ԫ�)�*��V[إ³�W��N�mf}H5*�N�L��,@*��!C�e��*ZV�)^g:]ڞg��"rl-V����RA,nԅ( 5��'uPZ�W�;J�%s*�U�m	۴�Vv��g���r�-�!6�:&,�2�؀��Y�cX6���N��J�:��x�G	75��L�ײ�{n^ph�6��J��e��C6����X㳭I-���msS�-UR�c�3m�7i�ٖ�`��� ��'j�t�PgL�t��H!Q��un�"���R�g.ó`�n'f�L�J��/�RɞBye�Ca��Z�{<�[���"��D�UU˭�xA�q�����
�-@QI��5۩櫮��eW8�k��l 8b�v�`p�U��T_&A]��K� tTO{������sc��Fu���n�����y�6���V伾.�ܡt�S�"�n��S��\�L�ˎD�%�����4l�c��<s����g��+Ea��ő�G'n�f�1�K���T�H��udvn��VB����ѝ��v^u�c����`�j9� Y淛:X���:`��[��n��-��ʷg����Wc;5SB�!<��l��א�mm��4��N�﻽���O��"F՘��As�w���E���WZ�z�e�f� ��ܦ�M͵$r6H܏�����7^�3ww�������`�_��ꈑG�5wk@n��6��[u�jo�&+�K�Jq�PܑX���@ջ��ԔB����Kv�g�gމu#)�333�]��]��n����S�'���]@����7u�jo�7M��'���`�Ԑ��zx�=jw#��\.���X!1��f�&w�M��Dnݴ.Hzv��/�����t��fc��n�$��>{���6�ȭ��JIT�*)�����+��s�D%
*�<n��Ϭ���y{�Ѥ�D���ށ�w]��ݽ:��V�3{�7�(���qȤl����f��'8$��9i� �ӨKjR���bQ�:��V�3{�5nk�;���@�zlZD:Q��)�5�=���t�'u���\���!S��=�xظ�+�\$�K�Jq�P�qX���@rӬSx��Np��]Hʀ����������� �O�7I��Y���PfbZ�"�(`)��f�,���Ib!(�DB����;���`o��#i=l��5R5;gC�*��w�g�{۰�uЄ��c�,����"II*�%D�>�f��j��`wٷ�@�y���ͣ]:t�����y9�{uOh�$�z�d�����(���.0��8���{�ul%H�TLQ�I/�j��`{�x��NpsOt�H�,*���˩9ʮr����^�D(��M�{=7��j��|��;�ImDH��d�Q�4�9�9�{�9i� ��3@Lɭ()�9Cq�`{}�ށ�s]��{Ϯ��eVUzECi��ϳ�o��]-N�D�D$����5���f��'8>Otr��PE��YE�5��;b�x����fF:^��un���ݎK��Ȑ����#��) R;�隺t��ܞ����`�9���T�R�×�̀�7=�Q
"d~Ƿ`l������f��m��؈���RTR,{���n�}i΀�78��h�F��ҍI$�@ջ����f����U��{7�}�Z\�ABDD����ӝ�78�'��'XG+�V��[�JE	N���H�C3sy{ci�;e�8:P��Ӻ�i��k���irʶ�G9YŎ�v�`a�d���Ӏk�z9�$��g�s-M�L4�9�7]'jG %�4�v1�R[v��9ذ�sFN�f�\��;kL��R�c�͞�5A�C8�6���vzT�����nM��k�d���3�-YN�����lw��(9�k"%δcqɝnѨ�p���u��|&���w4\��r��7a9�s�<g�q��:����6M���\�N�m�}�o2x��~�{��ғ�_Zs�g���R��c�7$V}����f��隺��U�+�f_�~i�8�M�W�K� �֜�T��ܷ��k�l\������f���I� ���$���9��拊��������78�'� �w�?�3W@3���!T�1GDC�!)Jۋ�����݊5�W��ęj��.p�3%O]�s�DpIT��V����36X��j�_ ����?i��G�F��ҍI$�fc�i(�
!U���l:nz�ٽ����Q7�������߽3W@��s�aD��݀6����h��E��Y�x]M�N��M� ���$����j�����T�)�BrE`?r{�	'x�Zs�y�s�?Bd�=��J3\e��ӋF�wn9���<-і-�V��v��⽵exɼOH��F�m�����9�<���=�<�*F�[��)*RI`o�3W@�^�������3#��T\T]L\U�;6Λ����we.P�BI-"V�!��������W_d���Q�����	*����߽�� �w�>�Ntͻ�K�e�̐X]����$���ӝ �n��۽�.{[aZۂ�#��j��f��	����r��'��(m��'�ˋk=H�r(F��rX���@>��`f�w� �͖}���d�8vK��@<ۼ�O0$� �֌w*�
n���7(�I,g�{���`&�3@<ۼ�"UC��
����.�v�S-��@z�t��|�dDL۽�eb�k�E�K���$��e��6� o�� I;����QW2��$u8܁q�5��f���� �Y��a��8�&��pљz���}�[m�6� o�� I;�K���
DpIT�I,�n������̽:���p�2�"�F�jI'z �w�6�3@<ۼ�ot����"�h�7%��r�~����@=������@N��`�e�V^VT�f����{�	'xic:���aU�攴n��QJ�Gt�Onkh�����3�	�Z����rv������q���,n�Ak����"�;�F�N�Ea�4m��%�e�Sq�knt6�-���S��a7ۢ�x^mu�����]����#;��E�h���t��9ˊ��;]��Y�I�M���G�n��=d��堻&V�z �(��n�<�Ue�V�:�X�rv�)��n�(9�������wwo�.�(���y��7����׎,}���6����x]q�d�X����M+m�'A)�nQ�x����w������u��G��w��!�S�������I� �,f�y�x|��铘�F�;H�*�<�9�7q�K ��Κ�(���{v ��t��#��R�*b��4ͻ���@N��f� ��EelD��U*J$����oz �w�&�3@��� ��0I�q36�3�$g5� l!=[�.2v닺V[1��ݣ�Q��L��Q"�b�I$�@�x� M,f��m� �7��VDӒ�R(F�6�3s/N��s�\���s����(��Gd�m�@�f;�3+��(�K`��7;�]廮�߼��	Rs�>�Nt��+鸫���n�� ~��@J���Zs�z[u`ex�c��t�� �w�f<�`o��s`}-���7v��������Fc��H�m��6M�x��myظ��k��q9+��
��DI���M(�]�d��@��� ~��@J����#��T]����^�N��m� ��'8�隺���%I*6�ԔG��{���=:�*D+�D��G�C�� ��Ap;HtM"�h2!��CHP֙2
K{��\z��oK��d؝�kb���"�)����h��,0�`���C,D>fk�4m�h ZZְe��$M�8���)a����5�83UPD
I����cè�x>�@Hi |҃�(��J���DH�J�wߪ�]��)$�C���#�� iD�Z	�P��SB�C�:Ї���
��l�N�U;P�U4x���`|QW��E D�L�/��{ߟgU{�}�7LF����&(ԩ�@�<�`?u�:��X�'���w7v]�Yu%�Us�?u�:��X�'���Vm{hT*��A#�:PeG�ݹ�n����ѥ37/MQ��t"��Y+r�𪋩�̝�Ӭ���u'?����ɿ�@���Z��P���)x�'��Np��@��� \}�֪N�R�4�Iށ�y��߽3W@��9��c��2bc�;P � ��g��OB�$�N�:�lmn�@{�b���h�D=z���3�y��e��;��������p�<����@J��7�zt�d�3`��U*�Ɖݹ��nvy�	ی�����=��,�3Ru��nEv�	�E8J�Tmө*)�����ǚ��e��>׺�¼�QATLQ��\�2��u%2k��,mn�@<w�I�6�JQ�G��V�Ϳ�@��s�RQ3�׷`7Og�}�I|&j��𪌊��4Kn���	Rj���^�sVڡa������*Np�c4Kn�	�lC[X�El�T���l��W�����1W+��ECm����u��m�J��f���)���;k�=��÷N�=T9�ö|��i�;���5ۚ�s� f��9[x�.ƺw�[��tT�p�jҫס�ָ��Z�q�6F]��]7d�[�;]Y�C�W����rµf��ڇ�z�,,cL�6Z����$�[�{[s${F{tn��yѹ�ص���w����𝱾j�v�91p�����p���{=�-pA�
�J�/(]�K�R8x�lrDs��v�g�7��XKn�~n�Ն*Z�Qi��M(�V�e��=-����@J��|)�Aú���������@��� O��*Np�^��Q���T��n�"�;�W�_�{@n�����=-��8%H�PUi��zc�V���-�v�{�3Z�z��CCn�j����ms�u����I�`n�a���7e�/�N�0;�$p�m�`n�/N����`f�{�%I��PGeM^�^Q�SY����뽈��)B�������r޻w�zt�[j�4�c�9$v|��
Ru�7��z[u�oD5R�M)���Ds���J%�{]wt�>��t����*]@��H.*�.��c4Kn��=��� ���OJu)�)N�Bq7$��	O��ٮ�#�	z��>ګpZ�{�K��x�u�L�I\���ۮ�߱݁���b"�7so��=H?"��*IQ�NI���۽P�S#����>�`}-���D(�7L�������NG;�5n�vﳟ]_��P� �1!XdHJ� B�P}4b��R��v�w�}�P�FI5��u�7��z[u�7�'X�hԖ�c�w,n��wg@�n�7}�ށ�3]���:�`��=ln�{����.��؃1��/8��ܛ<F�e)��C&�]s��P�J��(rH��f��bI� �,f��m���K��$����G9˰2swRP��7q�Kӻ���;��<���씅�S'9��������릥	L��۰���/�)V���F�!���>[���f����uИ�B�T(�J1�?����V�J��NI������5�n����w]���f���L�8��gW�,�[��W��a&Ǫ���n��%8wg��(������N9;�1fk�>���t��37{�>ܨk��$���TM�� �X��۬���
Ru�w�R[Q�uܱ��iݝ廮���ݛ
!%2彮����X��&�����
������
Ru�6�3�|�u��4��Sb!9T);�2st��w��zwv�o�IBi		a�X�%`�%����I0A�do{��i�;�-�n�Ӭ�ܽHn{l�g4.:�[l�����;�r:7��V��z��P�[���|�u��VB�l�P�ʒ歚�h�ݧ��iAܻ���n�2l�)k�އag��q@ki.��F�y�X)� �؜n�=sn�n�kI��B��[�hV�)�)���=��R��k/Pv�����$cYU��q58�7�+.�r��9ʪ�UV�X�УP"TNF6��j�ۮ��bNy��\�ີ����s�E��� IH\U2s��~��,�Qջ�`n���
#�-�t^d�V�٢��b��4Kn��{�)I���zw�UTԃQ[�*8�e(E$vm=��� m�f�y�x�
LF���&(ӎN�Y����Ӡ|�u���ށ��"z�l�:j8�Gu�6�3@<ۼ���
Ru�t�~w�;�2�Qy��s�>�;�IͰ��pvțjM���w�	����l������^�*k0��� �Ot):�k�nf�(m	�c�G$�����W���lP	QF�3.Nc�����,��wa$��>����U!E9n���������Ӡ��`n�ozո���-4)�I���3@7xm=�}�����)�&Q#�"�b��4�w�6��Vf�wr���T����1�N�IT�ˣKtr���;��E�3A��E��q&jc��l�I@DS��)@rI�?~����6st�u�} y���D����O+��4㓽 �� ��^���7w7��ʃtld��QƢrX����]����]�*�b�"�@�fF(!�ٴTv,[��몯~�����j�':�X�]4�΁�w]���bDD������zX���&��(�(RH����@�ʥ����7u�K'��@�m�SɮW��G�-ˣk;��m>�g׉.2��Px�j˞R#�P�E9n��� ���wr٠)�� m����&@MHE�L]]� �Oc@S�� �Ot�� ��$R��#e�I�������{�'xm=�� ��K�����*n��{�'xmc4?} :dW0�L�1�	�V��`�5�Z��\������������u����@Ż�������x�'IV�!�I%m�[s�{&�x���:�H�E�]�N8�e6�)$�MGjG`f�^� ���@����D(�@�����;$�	���yҩv������݅
d{�n�5�偛�zt��e
�EB�r�$��M�� �w�&�3@s���"��%(�#M�rw��%�6X���@s�� �Ot80� 2jB.*bn�΁��Y`9�u�f^�۰oy�ؐSCTP��P��n�zP��s��\d��}�X�{��B4�ް5�nı�efb� PUf`ZG[0޺K�YX%$JP���C^������v��Y�MNР�$1&RB��R�0Q4���I�
	�)�
ݙ�A�p�=5�L4�&��D�t��9�2J��	0�̃$�#��ɥh��\��՚&	I:��dF��;:@8�P�o��N&fU�td�w�Ns4�;�i�����3�4AM0�nM��!۾�#�w`j)(

-�*i�E3��ia$�;`ͨ��i*��!J(��:�wZ5����d��S�	b5�N[�d^����;����W]��r'dz�v׆�� �Q���=F+nj��e���En����B܁�4	�5�`m(m��l�k��is����6��E��o`ԙV�R�Ca	V �u�kzKv�D�F��0��Ɯ�� W*�-�-���J��Un���e�&��.J�NUúM���Ɛ�k���.���
pnN��vݷL�-�V9n=���@S���7��m��\�вD�!�gP(-<���Assjdή��W\Z��ڥE�ͱ��v@�1F��S��mW�쏞Ii��Z�ᴴ6ʴ�����ۭZgc]:t$�+:e3:�\<�l�sfr��a��Q�\�:[���'�t<]����ӱ�q��`�!�y3�����Zumu�N�	���/c��r�*��In���\���0�����m8������c�t�V���!�1�L��n���n/B0�H��8��QK6���vyS�,�>�
͹	J �����Yv�^r���N��ēU�s9�N7�1��@�D��n.�/B�)�7�3�[s�î�x�(U��/�Cӱ&�Mr烉�M%C����% �)�+�:&u�5.-cjcR0�n]�����'��V��Mt�2!,d$�U����-⇕D��Z�tcJ{���N�EF�0㴚��B�vM���q��*�kO��m U-��6��삈�V1¼Ȫ�;Us�8�\k;mp��R�PZ:�I1��r3h����d�t���12-�'p>4��n'�\흆��d�o����g�ܬ��:����g�la)��\�9�ԭ��z�j��V�vEZ�j�����Bf�P@:�]������ӡ�kZj���m)/�Of� �.K�v�;|w��~�D/Xs��ö��`��+��U�x%�J��`��[���mցT��aڜ��3�	��uu��4�*}>_��l��ζ�\g�mJ��Y��3� ��!�B���@Vq>A_��=��`�hM� �Wz�N��:���E�kz�hݚ�ַ��}�}m�������+�f����tc���Z�)�t��y�N��5p�tT�;[r6�Ɠׇs�8]v����s�=yz�l%�BƦ���cG�Ѯ۵ƕz���)�d�t�b�65*8�r��ڷ(̵��)L<=�s��K�@Vݮ�<exک�[m��nA�q&n7 �f�ބ�'CZ�:���G5]���=Z�c����ww=��e�2K��9{v�n�;�ъ���fR�����8�{mrcR�4�(��JN,����`f�oz��,��Ӡ}H5R�$��j]� �Ot�� M�f�y'x�<)%*#N9;��6X����y'xm=�9���QWqQ2M��uw�&�3@<��6���w�w�i'�);.X�[�:�f�5����	�����q.`*j�����]&竳���<X�o<[�,�l���˳��"n *(Q�Q#rt��w�I� �X� �N���*\��N�n��њ��꫿}�|��4���a�ȓ�$�	PM)�0Q	�$B[	(�g+��X��:o�=����;5 ��f�y\�@�ן� �N��{�I���I(���+�W/���Q>oy�7u��ُ�Jwuޖ���¶g��.X]U� �Ot�;�k�I���Vl'n�luM�H�49Fx۲��;r��N�u���1ںݣ�6v�͵����iq�ހ}����ܺ���r��r�ff�z�j7F�I)�B�29,ֲ0{��	&�@<���2w~��5��_;ΕK������:f7v}	F��%�J9�t�_W@�{+�T�QWE\uWxBK���9�x]l���,i����n��� �7x����[0w+�5&�@#�>?oln_�s`�"�����=s�.f�`�`r��z�lYm���#n�5� �[0w+�5&�@7xxS$L8�GpE���^�'x����vX��X���()�n� ^M�>n��ـ�^ ���������vX��X{�ΆD$���$���W��y`}�q:5�IN�q�$�3=4���X�{����8�QQVX]\���r��'a�f�c^�7�X�]��+�]r��|gNW��';.X�[N����`w3w� �n�3�K�ye�)�EC�r�ʮs�^cw{	L���:y�:��s�{����j4�7'z�ݖ�[0w+�7�{�{�� 2�d���&�� ��� ]������偕��R�b6QQ���l��l�/����|��q�{��%�2��#�~��l����5��ٝCu��;s�]m����{���,���+[V�t�ڇot콅�=�-�����Ϝ�vh�Ӝc[�s����ݞ��;\��J���38�s�ݣƺkkv:g��1���d#��%��	�@w]�9�,b�j"�����rtz8���;�X����slX�%���9طEY��ڶ@�s�Z��Z����rN��z�sք���=�;��s��Iv�rJv��#��8;$��{t�介���Iceۑn�%�5*J
r!�0�?;���%l�ܯ _&uw�HӍ��}�/�����`����?w��������b�:hQ�ܒ�M�� Sܫ �K���� �8�RS��r�𪋩��@r��y'� �vX̚X���(�uSr����I�>N�Jـ)�*�99�co���-�қ���[�i�6v��b��c�I�
EK�q���W$�h.��@��� �;�9+f �ܫ �I��Z��K��brKٓK��9�r���`�{����(�&Q#�#�+��},>�]�1ݚ�d�{΀��Ł�1ySX(�H� &�;�������[0U�p�c�uw�u57W� �;�9+f��N�����.b@��i1Tm(�q��b�^�l���4���I:�#ۙ��*��ܦjqD�GrKٓK�����7� �f���W9\H����?�Gۗ,n��]�~��p���� 䭘G��G��r��R�+���z�͖U��;1D4|>�u־�}\�����ʽ[��H�5D��� �f�������
��7~�=��v���U?\L�5wx�l�5W)�7�����`z�s\�H2�)�rJ(�q�m��W�
��,�4��)�����Z��p�qpE���^�y�s�os{�����K��T�	H$S�����ިQ2�|�4��잁�/��-pT"F�Nw���`w2i`g�ج�۽��t���T���s��j���ϱ�@�{]�jJ!jJA�T
H!D��R�$�D@$	(��{΁��j�T��v𪋻��4<�`����� ՓKِt��M��I�"+�SED>p���;&�V�2��v� ��+$\5v���h��&殰�ot�w�jV�O����X=h%EQ$Ƥ�@7ٲ�ԭ��r�{���˨ ��'늚&�� ԭ��r�{�� }�,� R���l��U)���5{5��7v �����(�����>tjUK&y�dU�)��t��݁�%;�y`|�4�?{+�Z����N"U#n"��:lt��j���V��ٻW�u���tE��U�h�E�1�)����m�e��4��T�5�8�=�n��ܦ�ۗ�:�-<\$X�4��ظǛz�׷Y��rn�5����m�q�2�%�,'Hl�unx�h��ٲjn�uP\;���SR��y�n��l��CzzᆀnMU�R.9�5���bΓ�)����l���t~�����>{c��m�3H�8$��i��%��Hl$��Td8�0����D:j��dTB7B$i���o�t��:O���BP��3ٻv��3T����#q7$�;�4�1}�v}���}�,mec�'e��t�r΀������>N�jـty,�8�D9M�V}���}�,�M,?W�f�?���P�TD1������[0>�X�7��~��?>0�b�[�sj�Όc�Q�9tIZ��8���:���w9�P;>ݡ��%Ww�y���}Հ{�f /r�s )V��e�Nv΁�ٮ�9WʧE��݀}���/3���DB�>tjU-�H�%$�>���� �f���K��`g3MTh���4�s� ~�΁y�g@���]S��߬wh���qȚ�9RK��K�Ur�Z������ |��z:���U]�U���r<m�
��Vx�Üun:���pv���N�JT��\�Zn�G.΁�ٮ�ϳ��>l%!��N�����SRLC�ܡD�3����P�6X�4�1}�v����tJ����s� ~�΀�8Ο��o $���&%�֬�(j��5��;`b���L@CD��,5�����5���cF�$� ��&�ڎT!J\T�L�cP�E�0���"�@A&��u�]H����erp�.oFLm��[(AѨS`Bhɠ��hw�e%�hd��=::�
��$�Q�)0�B�4dA�1&���ꥶ�E8`C���$�)���ӷ ���p�	�_Il�n����)�0W�X0s�%I�[٫����$���XfjL�#FF(Pe�Y��Kf�L�
>���%=�v�hN���|_}����z���~�\��>����č|(��rSLNI`nd�����]>�wa��	L�=�@���~�"�.*��'X\���� �ɥ�}�'��Q�%(���d�RuZ�OrI��ץ-���S=Eg����q�"��	�A')"��N;3ٽ��6X�4�U�皬���!~pT"F��w@'xjـ/W)���@���N�r&��
I,ܚX��+.Ot�w�{���N��o,ɪ���Ζ�c���f;��|�u%����P���c@2A�3���|X�[j��(�#���`gٟ���� �y�r���a�\r:u�4ꧥ��w'<jv�u�7k�rf,)Ҡٸ��SQS�	I���m��z��΁���������1��`<NT΀7��MWw�&�F �ܫ �� |��pK �PE�L\�{�N�I���� �Y�H��95�5R��L�+����ow� �{΁��u`g�جW�F�8*�$����� �Y�r��ot�w�������/$\�:��e-��@��;;;���c\[��c�yҜcf��M"�B�P��,��+qil�2���7&��@�M�勾���]�m]M^����r�!�z���7v�f� r�3��/VCOE��K���f�\���%l`m�m7ilx�Ѵ#�M��SWa���ۚݶ��]�1�Ν��3�G:�����Py�Be�;�3r˰��mv�F�.c^��V ��Y2�k���^y���aJȸú�lh���l�ò���	�xO9�Xu�t����=���
/���,���Ru��v\-+n]t��V$���� k���">���s��iA�H9C��`o����}�,�˫��`o��u���R�m�'z �;�k# S�U�rM�$��R�Ji��,�M,_{�����}�,�n'�RU�F����LoN�޵���عk]V*
�Եf���Ok�<1pu\T��^�9�� K�� �n�w�K<шaY)6�8%WX\����鈐t���� S��`g3CCEq�I;��l�9���/W)�;�{��&��SwuS�����ͬ�ur��ot��?r�����'_�'��iX�r��?m?ӀrM�>N����=�Q�
ce�	��:`�m\����m�$w>�� ��v�\�UB�E�T�k����.1��&�~� |��	���/W)�5�"bMR����jN�}�,�˫>~�`{3w���+�Hbh�R�d�9΀�ή��W�z)K��"�%	|��\���P��۷`�y�^A#�!�qS5{f����y7� �;�=��X�KTVBA6�8	�`wɽ���˭��r�X��~y��Ƅ:�˻#�Dvr=�vu�rE5\uu�'vM�#͵�����tU��m���˭��r�y7� ���)krF�Ț�X�M,����f������	Pʻ��2f2�js�'8�ot�w�r�f���"�ڔ�V}����6X�7�����L!��2UŕS`&�E7޼�9W|{g֫fo6�S5TW9v ��:�wK�c���g��@+���Ji"�r�PaR�q�B��[��׮����ƺ��q]E�M],�q")J�4�ܖ��K<����v��sw�ubٚ
A�$�!s���`5I��7� ����f�S2�a��!�I�N+�����vY���q-ܟ�q������GB�9\��jQ;���Ϛt�{'�^{]�,���nH�rH4�3�X��O@��w`��T%м�$��������o�j4�Ѣ� �9�!�ˣ<���J�-��u��7�l�@�4��v�T�¦�ܮ����vv�H>����D����bԨ a��gnȢ���n|6ۡ���c:�ݍ֛V��5��g)IHan�8�;n��$xwSmmLqńq0;��u�1lPVڰ���\�U<=z n]�t��j���ݛnۮ�
�Nݩ �F�<�nJ��������������n���+�ۜs߭�¥In��x��gm��i�8�����Sk�^��Oq��w<������&br³��p\�����ϲi`z��r�r l�r�G��M�>n��`�����`�������vX�&�y��߳w� �`�[JU)�&�;�ـ.�S�o�{���3���W�˒.���4�9�7ɽ��e������o2P���P�q��tԥ;t��{lI4��v��]�b�HÂ6E�vɢBIڤ�'@�7���}�,g��y������GB��몯����?$0��,��턢!*
y�:t�z�5݁��TU1j�@��'%������?b�;�ot�w�tt8��̳&brʜ�@j��y7� ���;�ـtrYp96Jm�Ln+�f�z�ݖ��3�g��=T(Q�hJ6��	U[�%]�7�.E�uU�����]��-pM�%���g�:�:R���)���|�7��<�ـ/W)�7�{��C�$�����&�� ���O�V��� |��3O��pZҩEH�a�5{5ٜ��8�ي!(�)%	@y�=��zph�1����;�f�z��x*jp>�X��"MՓ�Www� �;�9SS�/W)�=ɽ�o���~��`�)�BBF.�˴spͼը��P%�;/��W/�N�9U��3 T����f�ڬ������������J����Y�Lef\��9�=ɽ���ʚ��%��eRr�q7���w� �n�����~�`wr�H�JR4�Clrw�������tu�zz��ЭJ��P��_D� ������u�W���jb��(�M17%��{���?b�>�7v ��:6��og���T�8KϯW����x0j�q<�Mu&���sZNT�[�9IP�1�:\iT��~v�����`{�{����58�R)(�D�ܒUE�\������ �MN ��+���QAP�r��w���`4���8���N��*]]��L]]�sWxNр.�S�.M�>ݖ��K9�v��hTI�tY��
�c| �� �՞�����3)�"J"��� ������S�8*�����7 UW��(���0QD	 TV\о7��BIDDD��?��?��'��_����O���W�~�ο_�������������?���	%��o��_��ͯ��*��?��* ��vO��D��1���?�?���Q�b!$�"",���?�?�?r/�o?������G����������ϟ�7�U2FIXQ%A!�P�RDaD�!D��TH�UTHTaD�X!�A�   �Q!AHaD�� �Q!�HQ$�THQ aD�d�D�Q�T eD��QRHE%D�IQ P �A��AQ$�R@�P�aD�"E%D�H�eD��RIHQ$�BTHPeD�YQ) �� �D�HQ%D��A �AeD�PaD�P �A�H �Q(P"TI%D�%D�D�Q�%��XITd $$P $  $Y$)�X��B��
�
Y	RB	ATY	BE  B ��	$"d$$%H��		��`X
@�)Y����H@d$d!�$��	�!��	�"Bd`!!�!BBPaVYB%"P�"P"�$!YB@!	 ���(AG��PP�P�BXV��`��!�a!@�F �`�d�A �RQE�FTI%U�Q%YQ D�RIAP� A�AL�3g��/�_����PU����'���}�v^����^������9�����u��O���ο��\�ʀ*�y���?�y����TC��@U_�� U_�a�Ј
��?�����9�W��z;����f���<?����뗟����ﳵ@Vo���o���*����ّ��g����_���@W���z�
������z7E���̳�;?���������������9�x�����x�:ٱ����z�=����=�����c�u�/�o��t������?����?�G������
�2�ʗ����������9�>�����3f�  �4-��ݨ  ��  h	  �   �a� ��IJ��@��B��Z��41�"� ��($@R����P��D�TR�P�@ �J8   �@t�� ������=��w�Q�{��� }��g�dك�����m}7�*����sj� �������WZ�>�� z2�Ҵ{�׭v�ON{���=}�>���Uف_wp=�{W��� �� �Z�Mw��J��P�s`N�� �#JS���o��t�Jnw( b i�͝ 6P X
+��:Q͔��e(  g` �a�Cu��Ss�� ��(PMgM(Y�Mp���)M.`=������}470:P  O@
 
A���zYp)M.c�A����N��0�z�B������@�n��|@6a�d2��Q�m�����Gw�<��)�>��^P��k69���x�  ��� C�ݔ4iA�N�S�{�!�=�w0 ��q�{����=�����=� �t��F}�_g��A�����N@c�k����w�yS݁��4 �@  ���n[��K�2y�\�>�v��}��󡝴��������W��}e����> ����J>��.z�@݇�כN��y����lϠnãs&�    ��)��)P  "x�T�Q�  '�T�I�=R @��TLR�@j~�R�R�  �!M�)"� �<S�N��?��?����?�5'{�t{��{��zw�@QW@* �������*
���**�EU?�������܆�`��	�X��]	`�,$
��X�$sg��Ჵ �$�S�;`��Q�R4Յ	d��s�Nf�3�6�����zg�'o;�����^��ۡ4�M�^�{���^]��{	��d�d�4J2, �dk%�4B�#��IYB֛�LaZ�	��.�e-8S�@��/	��)^5�B:�sF�:"F+�6�`M�3L�J[������L%Xhe�%�B�C�^���cˡ�<Yji^FY,)%%	A��J�è-�sM�1HG]��R�D�r5��
$*@��L1�	p�İ�!XR���D7
®;c^�Z$�1�n�a�[a�0w|�\v����} �B�(�z�˪?�wT{���P��,�������ne�b�u��s��Jo��3y���̥>�eL��~����նf�y�4�%���Y$9n��$�e�6LIIp���[i�a�-0-�`m8h�������(B!a��/��@!�$"|@!����dF@�d��$$B!HR!��ce$6q�V0�`ԑ�A �s�+�%1�@i¦���`FB¤B��D�R�@��±&��1��[̙���������1��4����X�~���N0��d"SP��V$S#L��1ˌ�h����p��e~
�?$�O�
����M�����XY>�ϘK���f�:�H4#RM�>������7�����V�P�� 0!B�
C��Sp��P*`cF) ��ā HBMd�9~�X�� �d��bA"Dh�B@�$��O�d���	�D�X.���H�y��w�%�f��4���cF64�)@İ�"4�0�:���I�\�!R5�HX0�0����$����3>���@��.I �N D �[$(A�Xх��8�FJq���(:Q��旅�Pނ��s0,jHP�%ò扎��ɼe��]������Yav}�i�\5
��.�%q��Ja.1�GN?;���a�k4ˁ(]N�6ꑔ{��?C��A�ɴ�	x�>�~����x}��"C��4�ӚN+"@��aZW
g��Ц??��f͇���#A�@�esF�Ԓ@��!+�cG	P�H�`ō1$���@�:2rv�ȱ ��H�\����)��r�f���w��)4�²d�WgY	׼e�	$����xM�9���$vm!R0����Xc
��6�B�.��y5�����I���D)��Jf���&Ws��
\8Y�w�w�(aA��y�J?�=aq���|.���?}���W_������c���g��&B��������1Ќ�$䅘�h	�F]��&�xn�&����$���z*ݝ�f��JŐ(;IsA.7|پo�!�ԡ/a�࿷?����0�B#V�F+Tb2M<�w�0c���5@�p$t|Mn���gCP��r�[fkc��/�?c�*D���(EJ�1�"E�bġ���2D� �B�(c*Ș�K �ŋ#Ǣi�����������f%��UHh�8`��}���0��ɭd6�R�4v�Ld
��$)��@��D4H�HH���J�c1��a��B!b��RB44ī��A����!�"E,�!�B�Ł�َ�L/P�ơp�����
�*BH,#	!B,c$�t"HL$�h�H�`�HH�`1��
�H��CDc�
P�©8� ��SO�]E���i!%��I��H��bH�E��8�L�o��S����ײ|�YH�K�Ͻ��xD�"K֒,���,*%0b�d���M&4��0�6�$�!�0I5��M���&�@#$l+�� �`CV1�e�A���(E�vn]Wk��

��$"�HE
6���g	~�]��%��I��C����6b�	,l
a���w�sz4�W�T1*�M�08A�@�A.S�]Ml'�~��>p0��Z�H$B78�Xo�\$���*c2�	B!3�T��Z�� -X�H%�65�h&L!H���HB8��A��0��4H� ��E�	!�d1b0���EMI!�HB1JA��)(D
���"M#cJ@�	���¤SP!	�aT� $�`a�S+*@"���"b)(P�MT��2�
d��(J�$n���+�h��1���I
P��\j�0��(@�����˭�l٢u���wZ�X����\7��$�	p#H�	IB5aL�s�淳�C�aґ2VE�!L#YBUN��0Ѳ��n���N�)��߲����q����;o�@.���󗄖��5c5��6��B�D�`ȄB4B0�jm��%�YE P�D��X H@�����G�S>/���$��)����)K�j���a��e5�g�K�{n�!��P�@�ˎ�kP�q�˝����xw�M�~��))�K-���'ا����;�}a4$i��LǄ��9w�?rW��o��hO�h��A$#�+��k���2�MI`JJ|+��  ��..F�a&�J�?d����hD�$+3ʒ�q���I���lw����$���"�� �2	"2B,�!���2`B��f�� I�B�j��#�vw���P"T G�_����P�� �y�l���:F	 ��I��L��7�wKú���o��q�h&���K���3f�����!y>e$eXR��aB��H�����ٌ���J(����$	w9#$8Hh�������>隇��@�bь?�(bcS>��A����r�~:oL� GC� �6,
J�G�A�3M���,c�jIDa���S!���M�O��)7���/���h�``F���bA���	�\5Bg�Y��HCD��$�`"bB@�n��˗�pa�1��I�i�Y� �0!`�%ft��!O,�
��3Od�&dd+$�J0�� �B�KƬ�*İ�
`�`A�a�H,$�A�� �bf���p�bF�� D�Q��
`� �����؛!�)�Bep�RT��@�#aY,0�nLۺK{�lM���HB�"�$�F |&�cV5��cW!BFbM1���)1
��~��#HL���%0�!0!e	YIL��#$`ȓV�\%`L�0�HGP�HB�#]˄i*B$��!H�0� I!aXX�$bI#IMBʐ��ʖ�#
���°��,���IH����2���G���kV.K/$l��-�Cp����a��/4�!��ui/i#���n�B\���
���ib�Ұ#����5���f��f�q�Ð��L	@�T�W$�GL.k�.kz�o_�����2, IB2H!�V?G��Y��o��Ft�np�����J���i,���(K��ZKIi-%�s��T�YRYp�"F�!HT���H�
 P����$tV`F)Ad��d��R�IvK�[
�)I�r���E���S%��!Ba�"�	�XXV5���$G -"0"�q&��!�k�[�� H�h�����1Hք��V1>�R#@�F�b(�g�4��J�p�D!$dP��B$�!��*Al
��X�F$#L5���`n��5��3i���7��6�H��$"Lb�vh�Д���5�c��Dia�HV01MI#s������9�R���	�ga����UUm
�@ � ݰ ۶� ,&�֡Zy���U����jN�[��mؓnu�$�[U���l��dj�V���ʱ�VI ?Y!�B@h�݃�ԩ0 zzFj\�@AL��m@UP$�Ut��ې���锉F� �@䆍l�U�!�� r��oHV�m� �a�Knd싔�b2 pR��t�m�i�@�А7m�n�  6�@[Bޡ�
Pn�F�v�v�	R�*�իvږS3}U�݌U*ҩ�v[܃s�$�K6ڐZ)Ij��4$��,�6�1Gkz����[��ml�lqt�U[��e��
�W�Ŵ	�`:Km�d��^�  ��@�5Uu)*�[J�ԣ��g�[Fݤ��͔� ԫ��\��ʪ�mV��Hu�B�m���,%��Y�[d�Ͷ imp6�!i���Cm�ٶ� 9����m�����F�6�  �`�� ^�:ɥ� mm��m�` 9m:@�ζ˝�f�� ��{v���UU �m��Ƀi�2�$H�pB� -�q6굒 D���o.��m��m%� ��im	��۸H-�m����� 5�m�C��]�K�^�N����7��-����,��eK��n  �`lѶ��#m�h���Km����U*� u�UPʵ@A�*��{f��ɩV��)�kŹB�A��UUT��; �  6Z4^���j�bmu����NU�U핗�������b�Mq#I'n  ���+"��6�W]�5�bBW�h��,�U@���f�í����$����@�Ë	�i��o�ԫ�vqsUR�EqkJ�m�j��d��r��MI ;j�:��lY�g��b]���S�
����*��ڞKU@ -���햁&Om����� �� m�  6��}R��+r����Ҫ���nf�lכ�  �յ6�Z��`	e  6�^��cm����lkXF�cu�3����F�
�ʪd2/M��p6�&�nk6�Uk�� I��R�	6.��k&�6�M#���J��cS*� mUSʁm '[4�7m�m��	 �`�g ���I���6� [[l*�m�u��u����� �c�~��j����M�jQ��)�c�q%�@����md�$5UV��)��e㭜2�ҭ�p=��5n�UUʀ�U�p�����j�͵�,�`�[T��ugl�,U(�W\#��4��Z׵�`�vԥ�5�ݢ��\e�-A�[@ ֛i�D�WM����Pv�[l���]6�����UC�r�[u*�-G8�UݩT��Tk<V�/�����6[E�[MJ�K��	@mN��-`�  i.8�D��o ��94�m6�z�Z�I��ĕ��^������uF�e8���;���u�ݞj��:ʐ���$���p��_Mw��n�bj�IV
�Q��M1X|1��n�͔�M��۶�ո6��' 5v�m�E��8��H ��m��N׶ �l;�ﾫt�9.�H)ؕڨ4̇���ޔ�k]�2�yۥ[���H {P-�Up���h-̫@m���    ��[��ڤ�Hcj�I��� ��&�r�p�M�U���lm�H �ml�c��y���pL千�����Pkp;8`kC+�����,�`�]�6�o,��K�vR�K�M����=�iV�
.�U�M�@�r��2���p�ٽj�uIz.�n8x�����	l m�H�m�Mm��  3s���v�/6�U��,��� p6�m� i��am[�� �� '@�    M��6�BCm�sU֭�8h 
�ʵ���$�UUPqR��Ul��Uթ
����:�l�
�y��q^U�6,r���ح])���-�K�5��f	�oR��L�6��m!'KU,$��u�q���'�?+K�Y�ʶX{s��
v�Z�u(�f�'Bp@BR]�u��d<�]SU@gV�R�J�^ŵr45�ڤ����6���m�#vȚVض���n�L ����kZD�� ���v��&�l�A���k~��K@$H6ۀI�V�t��-� ��	 m��,$m���m�A���l pvkp�m���$ �i6�Im��L�j��
K�yґ-�I�$6ҩ9����6�=���[̵�`stP:G+j��V�^Z��x�v㥩���(DT�J�nܗK�HN�;J���8 Ѳ��e]:�[UN�Ѕ� ���b.��p��Mc���Bm�o��ˁm�9 � � -�Vč�m��U`���۰9 �Ί��V^ZBj!�V�m�kh-�m��$H� [P�k[��lH  H � ����n$$$]6ݶH�� 	i�M�$��l�C�em�m�� [@H�p-5�m�#j��L�  ����B�y[<�u�]=��\����t�5�;��������UZ\CuUI�$��&�m�#e��f�j�.�N�ձm�	uߴ>!�ݭ������������-�a*���_�x�5���QQ�tc;H�]V�A��ж���� $�M��*�a�#�������I��� 		 l �  m��;vJ]��� h  H� �fӧ`-�ɷ6�*���UYP)Ij���ڶ ����d�  H�6Ā:�;0�qr�sK^���U�ڹV�jAԶ��c��q��Au�x�Ft@��k�R���r����j+0]Riq�U�mۭ[.ì�Шэ�Pl0-�ߝ�'����3��M!mp����6�-�v p �I�H�q6��$sj�I,�����C�� 	 6ؑm�`	ŵ���;gG6[j�Z�>^�}�Ơ8����rM��zZ���bD�R�Y�4���mI�mז0.�s�1m���hm��	�ӭV�Z�5�Ƽ�-&�DWs���kv�ct݆�S�Z��i˱UV0�ԫ��V ��"ѱ��6`jk��J6�$�}hj��#�� �MդͶs�&�L�6�:a�fͯ3�m�n��v�W���^���mvjE���.�姘�$v��nx���6�+e��5vT�B �;
�����Ul@WJ]�-�Z�PW��*��KR���id��}�$-�O sh8�h
��.��5UW<�!;v	P+j�eUeZ4�vҠ�M6����p�-UT����W$����mv� l�N��6�oU���		ڨq*�nV����7a��
](;Ub� �m��?�Ϣ�fհ`����l �2M�g��`	V�A �`�ֶ�  ���M� �^��  [R��n��4�hl�$ ��Hn��屮����	6m�  8�`m[F�۸�m��  H��y������m�´�UU�eP�Um"^g 'K҄�v�13۶왌�UU�BC��j�Db���c���_Y�I��袥嶪X.�#�@	 lm%�gd�#"Y:�l�<p$�0hv�1:  I�� ��'M�K�[m� ��շ�m��h 	,���Ҭ�����&)����RD���Zq���b� �!6����ն�U�k���w�5���8N&����&����RF�Z��c������p�im�8��ְ6�e�wWL/�׵�n�n�l;Nn�$CumT��!q�q-z�tkC���h�FEUz��H˵R�lK�i5�� n��5[ɖ�@k�\$�kh  �Zl�kp�zOT�m�uC�	�y`6�	���t� �� m#m��nIk�@j�t��T�k�ܠp֋�g  -��5�[dֶ���	0+j�d��kz�I-�t���^�� ��M����;�sJ�u=�A霉����&�[��$`-���9&��lP�����	���T	����޸  �mk��m��m��ΰ�im�[%8�I���@�lH���I��Hm
���`*��:���*�-��I��S�U@�   	i ���j�s��R��M5/-P*�n��]���mv՞KE*�qt ��-�[D�:@�m�e�r΀  m  �@h     -�k�h�n�3Z��i6�8r�� 6C �2ڶ��M�i6f��X�F3����"m�n
��Cm�p6�i��ؐ-���l'd`�m����ܛV��6�ŷ���-m� ��[��i),6�ݶ !�͛lր ,2��9j��v���](�$n�:I  ���`m[� �f٭���m������۬2p7<�D
U���o�
���m�� �@��$�m#m�ʐ�>X�ت�ZU�;M�e�ܐ-�m��[�b@m�e�� ���-�tm� 8�t��m��.Jm��-�z3� �)R�\���WUp��-���l������h?��,` -��n ��@ � m�ہ������{�T�h�@v�'����  �?
A4<�J�@�8��[��"/��|/�EC�(��z H G�ôz��C@��BB
� ���;O�E�0"DS��%ҭ`��� dN���Ϫ� �6?�?
�b��:l !ċ b����S������TTt��D�D@?*��j �S���= ���Wf���|)��t��C�P�DL�����)��i���:>��N*��WZ>Q �mN�4�~T�A��v�&ѡ'�p�&�^�Th���"D`"�"�"��4 :�8h4�ȔU0��V*�����`�H���u�D�T8�(��3�Дڊu��8�?��G��#��^��#��!E�!�Q� A �E/�����C�����"��b�ҏ�S�=At���U� v)�bAb�X#��#�HHE$���RҔD�B	X�RF� ��:���DU�$"�VI$"E��P�TPҜ����k Ev/������&!�(�Wg	�*�h39�pQW��U%�b��@��{Y��Pn�6e"��-���"^� ���G�PdrR� �ci��) /<x�T�T��+bd6l*v����@$�ơvY�ym�#;:y����ւ�� Vu�R�݀+c966��F^N��A�ݷ
Aɻ'PF,Q��^Wc.;��@�ѹf�Jge����WG�SKͼ��L�6[
sh�ז2Ԧts�̪���]�m�V�nE�0��K��++[\I�V�"he����I�MZF��3u]��-9���b�`m�f۞ԫlYn۳a�I��:XuS�۱���� �{cWq7�i��L^��ST�Q������B���(�@Im�*d8�B9�Z�qG�=����喖̒����v�i���AHh��`;g3T�@�m��2���J��dG�'��u,Sv^��\�c����F+v4l{X�aͥE؇]zm$�&󘱊mz���(M��h�'@��˛v�Vbj�j�P��'4����\:��l�<Y)��)]�#x�8eWhw\��ۨ�A2���smI[�`�66�$b��Ӷ�Ȕ�r<a���/uӌ+Yr�ԪUC��b5W9H ֹ�f��]����c6eb{Z��'��;{aw���ʲ��O;=J:v:ؕ �\*#ɥ���ZG8k��Ph��V���c������A��)�[�n�+4p���8�<���-N��\jÑSܴ�[V�;ͻv.	b6�:��;�2�.�G.�o6X-��%xh�gs��&���"b'C�,�N�Ẑ��f�v�kdR�mۦ��6��s�+͕f��#�nA�m$H�[�]B×<�Y:��]���^90\ݶ�sj�t���:І�JcTn�ѷ\����vx,�h��Z�7V7^�\�=s�-E; ��5Y���즌�� �jLh�Dp�8s�I۫�Ȝl�ЛR��0�8�5۲ �u�������i���X;��4P�I%�U�UK�����`�Q]��:|���G��]�*h�Q��v �p�4#BN}�K�;�K5�1���Fj��M�X��q:-�����q��l���^�֏n�����ś^��3��	Qcn�hi9N���L��]�L�rl��%���,��b���/)m��gv�x0l�A�J�YE6������ڶ'��4G-z���,r$�ٙq\�s9�)��m��A4I��bP�)����&�#E:ͬ��,�֩������I�fS�����[ "�< ��(@V������@���ud�`[��ξ��_ 7������E:`��jݬuȳ�H�d��uwc�;[���ݪ��J�v���o ;$�����X���-�n�];��� ����x�`E�s�;�n�5m�ݫj�]��]���"�>��X�#�<熔�M�\ژ&�m��
'��-��G.6�\s=��j�
��Z�iG#v���
ݤ���E�}%İ�K�5wc�;�]�E+v�X�ӵ�}%ķ�<CH'`	�ܙ�{[�v��rO���C�%�����n�ݥ��^����X�\K ���m�贛��� �ݏ=�UW$~��;�_���s�o���	���
t�ݦ�x�`Iq, ��]������+�*�;/;�<2މ��1��l�b֋`A����
��-�;X��f�vJ��`Iq, ��]���"�7���n*m���b�K ;$�Wv<uȰ���z�7O{)SV�ڷb�Wwx[<��"ü�U_��+{��*�.*����kv�I?~�u����5N�իI��7\� �K�`d��jݏ ��tJ�ڠ��ӵ�w�\0�K�5wc�7\�V���/������Rf �_K�m��R.���]]�e��,��!yi����s���]��%��c�7\� �=� ����7E�c��� �ly�URD��X�� vIx!Ŵ��ݦ�x�`�a�RF��z��=������h����g7�lŀ�^��+��_9�s����r�ʪ�&dXݭ��pTڠ.��v��K�"���X��X��XY���f�hku�f��m��rg+�U��n�-juU�7<��62T����#�7\� ������� �y���]+��jդ���E�H�7��^v<����T�Zv�	���K��\�^[<�	����-�[��+cwv�=Io���<�y��E�l{-�qWb���+n������E�l{/7$����rLS$P`��';i��O{��Y�
9����9.pf��ϗ�+^��N#f�V4�렬�gx+�d�4��7��'Xf̡5���+.����/"	�b�.�����z�=gE��a����{1�ڞ�\W�%�n��"XUc��L
ځ�u���fۗ�m0-��Em�85�e�������U��ĄېgzZ�v��s^4�Zl��%�%��J� W�a0�}����Ni�NI t���d��ɇ�s�$yț�z<���Y�4`�s���Ek`c���4����� �{�}�q� ��[�����JVZV+�j�v�`v\k
�K�5nǀn����E� Ҡ.��J� �%��c�&��eư��)S��V���ww�����x����eưl��kL%��]��+V���Mr,�ˍ`�/ ջ7@�rrI��{=&3M��RZ6k��������pV��5��r�\vwn{�(�!�[�AiU�k�;��� �%�[��\� �������XZ�J�$����~��C����Ck.<G�`wf3 ���Q��Zjӻ��v<k�`wf3 &�xޜZ�HaN��nӷ�ꪪ��=�w}�f vIx����t8�n�t�]�n��vc0l��z�������X�m�um�BH���c��ֵ�<͍��+E�+i��3��p�k�s-]*Hn�k����i�f vIxV�x�`wf3 �b�:vR��n��ջ��:�c�&��vc0l��|���B�ݫN�+�;x�"�>��f͟R�T�UWj��>���uM� ��q4R�j�ҫN��vc0RG�unǀlr,�C�"vӥahV�+�`��  ��X�ٌ������[�]�,R�sA�y�um2#4qЇ9Y8�=^U���>��Yr�Чn��[��� ��1��#�:�������ݦ�;x�"�W;���/{� �ݏ ��ӧ��JӺv�`wf3 �$xV�x�"�;�6�_n�tҶ��#�'�����>�w�rDM~�lDҡ�Y�s�����t���fJUl�\-��v<�ʩ����wg���#���3�����K����l���m'n4��9�\�7�H�\�U��$Ů��e�X�#�>��f�dxu�Xخ*h��j�Zv����j�ջ��Xv��C�N���Z��ـj�ջ��X�ٌ�>���Ln��N���[���E�}ݘ�V����-d�SL�l�k �r,��9�Wv{�|���rO�gݻ�*�*2 ��>�˰���us�Z�X��Ȓ�+�a���'Gr����V�u��K�cpϵi�Ԅ�����]6���q�6{[��c�����B�"��8i�ݶ��C!R,f�Z�u��!�ke,X(ƶ��E a��*D�/K
�؆���x�umI')e4�l�+�G{-������EX�UK!,�pfMF���kN�흭�� �n.Ԩ�m�:T��9�)�9���R^��5�����g%��8,�#���s�ѶlFzq�-�vX���ͮ��[��ߠy��� ղ<��,�Ȱ�6�.��ͥ���� �}�z ?y�����$����>�$��:���N�2�[�x�K�{�$��px�K����|���{^������t�+s��I-R��$����>�$�K�Ē]�ؾ��q��Qĺ��W��=��}�Ij��$���}�Ij��$��s��N�5�)즐9"6�k���z�o�fr]Q� phV�n˷L��`���.Iwob���.�U�i.�����`p����j�p�v�@��o9�h�P�Q",
�Er� ;T���vf���>�I-R��$�YҖӜbL�l�k�KT�<K����%�Ȟ$���N� �ۮe��rVt�j� }�||�Z���I.��_|�Z���I.����"�"餕�}�Ij��!n��g�%�\$��d�>�$����^�ٴ��)�֭�DV�ͻ��4m�Ē5�WW N��Ğ�KW���8mn��v?�Il����%��#I}�||�Z{��@~����Һ++s�� �s�$��>�I-R��%�7�'��vs�qSﱾ�����]Hm�����$�-���vf�� ���O�Q{O��r���Y��UPԆo��>����HE�$���b��1�@�? m�]�ĉ��<�c^p��;41����v|D6���
&���r00`2$"�!Q�P8�+A��b&��q��$����C��n CR�C�A3B�,axrH�2	��MĐ���E��X:e����B,�r��TtH"���P���8 Mp Hq�!t�J���`��@B�����'� @0~!�G����	���&��U~>�
=1?Њ�5�������7����-�ʐ��e�k�I{�U�q�<<I%���$��1������'&�Ͽ��ﲇ�c� ¬��d� ���Ӿ�>���'��w�������.Iw�7B}t��P�Yv+�v�Е ���-/��gXl\6ݳ>6��?���'&׫���������}�zI%���}�Ij���*�U]�IO_�/�H?��4g�l��SJ�� �y���USmE���$�˞_|�Z���j��U^��������\�2��������K�{�/U6�~�x�Kvy�_|�B����\��W�>_=�ߎ� ��sv�~��Ü����,@� $-b(��" ��T6��~���7m��=;.]kSFkRfL��^r��{�{ٜ����PE�=�ku$��_�$�ݽ3K�[V��.m[;�=��v��R�Nrv����4Ǯ
a��\�Ÿ��;_S���k�]IM��I~���}�Ik�Ē]�ؽ�Wz�Q�yz <�]��͆�C)���`>�k=�Us���\��䒍���I.�c����9���O8���1�e�Gm���{=�w�%��Ŀs��*��ݞW�$�~�'@���<���-�;���;�{ٛ�����p�-��v�"���^�w�������Ԭi��۠�����$�Ur��s�{��u$�����޴�_{�� �9g=�^�Z�i�D���*��tc��;��Ä�0,��r�;^��A��nw7�m�bfL����.��s��Om�),�
~}|Xq�X����GS��,[���]c���7���Υ���ӵ���"�JI"��9�$[�淞Z�g��V������ga	���47d!2]"LC��m�)J.ո}Pl��)2�2#��a[9��N��:�,�gSA��{2|�[te�{���6z������{0���5���w�q��Xb��3�Ϟ ?o�� ���Ӿ�<_}_��@����� ���H���,�k�� ~�y��*���@�o~�}�z��N��P���F��h핣+�=� {�� �o=�}��s�ܓm������￞� ������]P���^�8��O[�������5�$�������W�~۠�e��?L�kt2�v{����t rs����޾���� ���n�߷���<���J_Xt��Ñzc�&t霚�����5���M��lB���>�y�]Q��-�;l��2y��I%6]�I.��[�_�\�n�K���g@����X6��.�� {�oH�D�ցV��9�K���������� ~|�׾����I9�m������ph�cl�}�g��=<�׫t�>CZ����9�m���kv�~>^��Zm��;l��I�'���ВZ������^��*����|�A=���\K�1���@��={���A�ߝ��߳�`�ok��'���}�����lX�nm��%��*r�e��,��d+��a��-ҵ"��{�|�~�����Ϟ S���t ~���=�����f[~����[o��n���a3Yk�u)�w`�o~�}�I'>=�W�Ik���HSc��r���[(�B~��5�L�=����� �<�ﳹ�'��+�6�y��o�K�}�ݠ~�}�{���=�eYnQ�j�ܒE�{��}�S�~w@���s�`}�9�z�� 7�ߡaWa\��!M��$�U]�=o�=��`�E�~��y7�,� �sJAY\�n1��XZ��XZMq�X�\hڲs�Rڔ�;��._�9�n��wn�t���x͸`�E�s�=�{z�'��2i�f�5ʻ�lۆ~�~������/����췞�+���y�,ZY���
����o@��ذ�*�.�=o ��� �m����][���C�k�T��y`�z��nM���+A0>�9���r�Ώq�V�v��������r�=3��yzy��ǀZ�je8��-���x�%C��m�;N�c$����[<-�����9�����up���e2��m���`M� �6?r�U������T�y��7Aln�ـE6<�ʪ�s���U��/���	���o ٷ���*��Qe
z��E�jӷ�O9�v9-��s��%=/����J֥&�I�m�V]��X��[������`M��rI�ɽ��נy�?��d���&k�v�n�?O?���� �r[�W9������]T���X�h����W:�\�k�V	Q��u�K�S:��L^���k�vC�̕�C�Mɖ9�9z�Ĥ8���N˸��q�;hM���J@:���lW[���bף�b��S�hɕ6N��uJEɮ��9N	��{]%֬����R��ҩlvۅ�m��;�^0��!pT�Q��u�S;`]���I��2M:	����Z՗�T~P`�';�΋Ҽ�$[�Z�F�6�E݉���[�{"FC+y���\���CF	�d�u���-][v����N�� �r[�'^ŀ}6�NZWi۴��N���'^ŀv9-��b�"����N����,E���v9-��b�"�:�,t��GE�N��[-]���S��`)���b�;���V�h�I&�-��v��ǀN�� �r[�'^ŀ}J�5q�b���T�k��G���y7!��x{qu����R�Rw糭�̤1:������,��o �{��/O<�����.�V]��M�?w;�f�6 }eF)[�K6�&�O,���=w$��}��w���ߔ'%��g�Q���tL�*���締E6<=�Ur�����o��o !�pq����voC�I'9����w@���� �r[��9��9�q{ny`�W��V�\��j������=���9$����k�XSc�7�r;E�ګ���|��`)m�A�.݌�n!,�r�ih�f�746��y��99��y���6	G-��9$����o�=�y`M��r���W�=�y`?y�N��ҶZ���N��?s�9��g��ߞ�z�c��z����Kmy]	5Am�m��<�<�	ݸ`�>����s���\���vݿ߭���� ���R���ƭ;x����o��o ���e�{绠}���6��
��vV��Kx�ذ�ǀN�� ޲�m��b2�%Dj�7%�;0`�S���5iF1�Iu�#���7e0v.��ӻ��s� �lx�ؽ������7���Lwe!��n����s�g��~x��~��N�y#����wui�;m;Wo �� �r[��+����� ��{��>�8�%m'j�����-����k����Usk�*���v��R�����rN���OR,� �����痠{9�I�?���@���� �r[�B���݁mU�t�v��=�[�����$4����E\�]�Ϥ�8�O��էm;_���E����W>A�~��5j৩5J�.�jӷ�E�w�\��UUj�?߭����`M�?s��ש�U�;uwL�n����[�'\�r�����<���<�y(ɏ(�#�2��rs�O�&��?~X��ߞ�xc��b�WLn+��ٽ���7@��I?�����_�N�g���rN����H%4 }�LN�W���0��9�0SaT�H�b�oO�]sp1K�bqO�,D0�,�wG݄��蕅 P��6�~]��B+�L��B?�q�Xb�������$`L�G�Pm!\�f�j�JU�%�eŢ�!Q��H���J��9�6�6�m�V���(I��t�F,8� ض"�Lc)t:����tN��m��KK���;n�
����~�� �h~���}j����nь\����h:�L�FZ|g$��
�Г��v�Y�Z�������Q��Bh��\����5���W��̩ڃ8;͋�؈�Y ��(&L2Ҡ[+Yk-@��>�nzy��,�Gh1���m����6�O t=;`4���뜦ֈ^Zn!44[u��Dv�+�f�x.x|��լI��'�Y�r�9؛��/�m\��=��!s�IT<d��èT� �m�K�F�l� �C �ז�� T�I�.�u�اka�-�ә�В�)�2���'"q(p�5Ca��+��#k��lH����lRm���|��1��Br��R9.M�]�H糔��gFA4`L�p�����Lp=i�Gn2�qr!�������v릢 �n8(h���:`�H��X�]��y��~_�8�	����ڷJ/-r��;vӛfui�B:��W��g�ÌUU\�!++eq�(m��H�6��1�Aq�ENlu�1F��q��&'��I�K�=�	Wb����YL�h����L�a��Ie^��4;x�!��"ؕ,:���M)�EF��5jc,�,ditgK�%Wa��O	b�+ƭ +�u���5�WJN�$���%��G0�Fmw;�u�M��v��'3@�(��[WR�/9��[`;2�֒��v��$S���=�����1qrZA����׭6B�hYvh���:. ��3� +�UJ\�.�֫���|���5�9Ui�*�Xӧn�^��=g��lU
��x�aͰ�0�<gd
z�@���kEع��|F��!�bd���mr��=[�0
fW�]���&���cEhL�!4�n�/E1���:7U���u���6�ʫ9ܜ�����9�4���*AT;� �~8 =D��(��w\��$o�lk���®��t��B5�0�JXC0e*a�D���ē]V���D���[p0�m�6��B�yt�z��]֕�d�]�d���o#�=+5U&�01r���iZ�54��G�1; I����k� �<�Hb��[O6�E1�2��-8����N�ݜ�գ�h�g'������$����g�A,��&;=��v��߷Kg�a������:u�vn�r�;�E(�n���bo��'����]١���U�x�<��%�uȿ|���� ���!k�͂Se�����NI-=��X����y��6P�z�WE+E�����{_���Ǉ�����x������m:���j۶ݬs�K��� �� �r[��r�����j�ħ�ݍZv��c�=U\�o�޷���,)���IBt:�������,!�MX�&�3jM43��G�]%�2Ư����7��sp�+�|>K������ND�,K�k޻ND�,K���6��2%�b{^����rS������YN���.�W6��bX�'�׽v��O���*��\#0(�B"�GE6"r%�����ND�,K��}v��bX�'�׽��r#bX�'���h̆�K�R̺5����Kı=��iȖ%�b{��ӑ,ı=�{ٛND�,K�k޻ND�,K������sEҪ��듻�^B����~z��Kı>���fӑ,K�����ӑ,K��{�ͧ"X�%��;��ik�Hb�]�O�%9)�NO޾��"X�%���]�"X�%���}�ND�,K��{6��bX�'�����ht�
�a4��2��X�N��6��� �;\��ecJ�ά�l:��%@c��f��ND�,K�׽v��bX�'���m9ı,Og}���2%�bw�_��ͧ"X�%����t���ՙ���f�3WiȖ%�b{=�fӐlK��w�ͧ"X�%����k6��bX�'��z�9ı,O����	&���W5�ND�,K�׽v��bX�'�׽��r%�C��`Ț���޻ND�,K���6��bX�'㺽����չ��"X�""w���ͧ"X�%���]�"X�%���}�ND�,�K�������Og��3�·-�*��@��N���7�N����z%�bX��ͧ"X�%������r%�bX����Ǻv�)��4eH�R��m��`jU���4�<�u�s�Vm;��6#`��7fj�9ı,Og���r%�bX��ͧ"X�%������<�bX�'��z�9ı,O���3٢]j�nff���ND�,K������,K�׽���Kı=�{�iȖ%�b{=�fӐRı,N�������Y�P�f���Kı=�{ٛND�,K�׽v��b�%����]�"X�%�����r%�bX��&��ɢRMˬ��fӑ,KlOw^��r%�bX�{^��r%�bX��ͧ"X�����T+ � �ȵcE�j�號�����JrS���y���K��`�gl��|9,K�����ӑ,K��(����6��X�%����ٛND�,K�׽v��bX�'�޳ŒNh��Ye�� #u�:��� �.x���ͬ�F�؟IiW��7�f�2�f��fk5v��bX�'��z�9ı,N���3iȖ%�b{�����,K�����ӑ,K9)��x�=�(#h�-s{���%����6��bX�'��z�9ı,O��z�9ı,Ow^��r+9NJrS��璝�����fU���Kı=�{�iȖ%�b{;�fӑ,,K�׽v��bX�'�k���'Ò���'����b6ctv��r%�b���｛ND�,K�׽v��bX�'�k��m9İ[��圯�R9H�#��Le���o3Y�ͧ"X�%���޻ND�,K�!������~�bX�'����v��bX�'���m9ı,Lx��$��*2�R���}l�\�5���g��Az�;]D�&�ڠ*gi�����$���Jy�ik/Z�$�8:��Jƶ��`������G���� ����`����,��� ��@cf���q�6ֶ��{��&�P6���C�t݅)2e���39���i��Yj���tr�iNw&Ց�uhw0�^6[�q�a'�-���v�%/l�#�qq��Bl���?y'c��P��q�Mwex���35ú�j�2��u��K����_8�U����:�ه�{y�^B�~����r%�bX����Kı=���a�șı=�o�iȖ%�g'� �{�����wy>��%���޻ND�,K��{6��bX�'��z�9ı,O��}��r%�c��>����Yp�s�'w����b{;�fӑ,K��w�ͧ"X6%���ﵛND�,K��{6��bY�NO��=��)���w���NJ%��｛ND�,K�k���r%�bX���ٴ�Kı=���iȖ%9)��x�=�Dɰ�Wgw���NK����6��bX���G�^��ͧ�%�bg���iȖ%�b{���ӻ�^B���g�ξ]��������T���FQ�A�A��չ9���i���[V�Ok�/
�3\+��O�%9)�NO�����r%�bX���ٴ�Kı=�{�cȖ%�b{�wٛND�,K���2�--�ҹ���rS�����yﹴ�7�țR�h
w"X����Kı>�^�fӑ,K��w�ͧ"��2&D�=�o�).k&�ֵr�˫�fӑ,K������ӑ,K����6��bؖ'���m9ı,Og}��r%�bX��]���5�%�Fd5sWiȖ%���(������m9ı,O����m9ı,Og���r%�`؞��ٴ�Kı?|Mz[�.B�I�Yuu�3iȖ%�b{;�fӑ,K����]�"X�%��｛ND�,K��xͧ"X�%���І?|C�n;$�bFs�ë����������-�q�/S[�}_?Q�M)���r%�bX��{ٴ�Kı=���iȖ%�b{=��9ı,Ow^��r%�bX�~��L�K&�˭f�iȖ%�b{;�fӐ� `"X�����fӑ,K������ӑ,K��{�ͧ ��bX����ƥ�0�ˣ&���fӑ,K��{�3iȖ%�b{���ӑ,qD�D�"1U@�&ՊlW�2'���m9ı,O���m9ı���y�y�Z�h��Y����%K�׽v��bX�'���m9ı,Ow���r%�`�؞�{�m99�^B�|�~�A�8�a�q�'q,K��{�ͧ"X�%�{;�fӑ,K��w�3iȖ%�b{���ӑ,K���^���u��m��n��;qu�i��;#�<�q6�6uW�uM9���(�C9@S=�~���/!S�=���ND�,K��xͧ"X�%���޻�,K��w�ͧ"X��'��/��2cd�9���rS�ı=����r"�bX����Kı=���iȖ%�b{;�fӑ?�`��2%��I��n!u$Ѭ��Z3iȖ%�b{_��iȖ%�b{;�fӑ,E�,Og}��r%�bX����m9ı,N������.a&�Z̹�ͧ"X�b{;�fӑ,K��w�ͧ"X�%���fӑ,K�"	��D�
��:���޻ND�,K�f���3&�˭f�iȖ%�b{;�fӑ,K��w�3iȖ%�b{;�fӑ,K��w�ͧ"X�%��>���0�����vr����)7n7���n5
��@F��g����r�{]��3
���}9,K�����Kı=�{�iȖ%�b{;�f��Kı=���i��NJrS�����UGW*��O�,K��w�ͧ ��bX���ٴ�Kı=���iȖ%�b{;���QlK��z{�.I5r�R�WE�k6��bX�'��z�9ı,Og}��r%��bX����m9ı,Og}��r%�bX��{��.k4\ֲ幖kZ�ND�,AK��{6��bX�'���ND�,K��{6��bX�'��z�9ı,N�����E�5���fӑ,K��w�3iȖ%�b�{;�fӑ,K��u�]�"X�%��｛ND�,K���)��-`!�|Y}'2e�֍�VW&��
�u���n�Ƣ�X,���^κ-ɸ�\�[�M�ml���nmb!�Nݥe9y�ў=&�ݴ�D�,uE�q�+uyd4�6��K�\����(�E9ͩ�� 9nS�v�&��)b���.F7h�h6#t�"s��1f��׮�i�v�1\�կ9ӣ�;`���ۺ/�~~qѫw4�Z� S�9���;v�:�Хt��(���5a�/Fwc��2iX��*r�F\�ܜ�wT��]I��3V�Fm9ı,O�����Kı=�{�iȖ%�b{;�f�^D�,K��xͧ"X�%�z��UO�[�q�'w����/'��:N@ı,Og��������,K�=��fӑ,K�������r'�eF���{���.F�	�=rwy�D�?����6��bX�'���ND�Rı=�{�iȖ%�b{=�fӑ,�%9>�;�I�ɰ�Wgw���D����ͧ"X�%���޻ND�,K���6��bX�2'�����O�%9)�NO���N��iETur��ND�,K�׽v��bX�)��}�ND�,K��{6��bX�'���ND�,K�a�o0=�f�e�0�sӌX7�cX���x����W�:�s���5�HI!�� �)��W;��JrS����|�6��bX�'���m9ı,Og��6��bX�'���m9ı,K���0�����j�����%9)��׾�NCܝU6���7��{�3iȖ%�b~ϻ��r%�bX��wٴ�[ı;��|J��3Q�2f�m9ı,Kߺ{[ND�,K���6��c��ș����m9ı,O����7���%9)���>�����4u���"X�%���޻ND�,K�{�ͧ"X�%����]�"X�!b_{�M�'w����/!���T>0-�kWiȖ%�b{=�fӑ,K����ӑ,Kľ�|kiȖ%�bw�{�iȖ%�b~�;%;K=&]]j�K;��R�`B��^<'a�R�-,&���,),ڨ���8��eu����|9)�NJp���ӑ,Kľ�|kiȖ%�bw>��cȖ%�b{=�fӑ,K�O���ؗY��)���'Ò����wƶ��bX�'��}v��bX�'���m9ı,O�׽v��bX�r{<��f���uUX����NJrX�w]��r%�bX��wٴ�K�����Z��:�(@*
h�x��!�"�0���a1Xc��R���$� \� ��H�qi��&�� @�3��A��Tik�4�VS����� �@18�%��r��'�o�� �"��b�#y"u�P�A~�i�?K׊�|(4���P~~x��!��|*��(��� �P���t��Q���?D��~��r%�bX��{ƶ��bX�'s��h̒j�֦CWR]j�9İ���6��bX�'��~�ND�,K��x�ӑ,K���w�iȖ%�b_���D֮�&�k&\˭kY��Kı?w���r%�bX����"X�%���ߦӑ,K��w�ͧ"X�%���x�k.����8�s]��غԙ�Aɍ;Y�}Z�#S�:W�m��8�B5�h��֎:�Ȗ%��2&w���ӑ,K������r%�bX���ٰ� ���,K�k���9ı,N������a��Vk,�֮���bX�'��}v��bX�'s��m9ı,O�׽v��bX�%��}u��,K��!ӹs3�j��MjY�jm9ı,O���m9ı,Ow^��r%��(T2&D����kiȖ%�b{��iȖ%�by�Vw��ɖL5��W5�ND�,Q�׽v��bX�%���kiȖ%�b{�ߦӑ,K�D AF؞�w��r%�bX�>�ߍL�&�CFL��j�9ı,K�魧"X�%�~���iȖ%�b{;�fӑ,K��{�M�"X�%�ߵd$��}O�^\N�-5Ӹ#��`�z꒮ �(������ٽ���#;ҝ��(�kF���bX�'���m9ı,Og{��r%�bX��}�h r%�bX��{ƶ��bX�'s��h̆�3F����sSiȖ%�b{;�fӑ,K��u�]�"X�%�}���ӑ,K���ߦӑ,KĿ���Z��f�U]�O�%9)�NO|}�����bX�%���[ND��,Ow���r%�bX��wٴ�Kı?{^�.C-�d��ɒ�WiȖ%���}���ӑ,K��}�M�"X�%���}�ND�,K�׽v��bX�'�&���`�@��6G��JrS������6��bX� }��iȖ%�b{��ӑ,Kľ��5��Kı0A�C�H�{��gٚ�d�asYk�Q�p1�4�ngb�����W�78�*SVN�d�;��/4�������u�n2DÝAt3OYCPL�y٘u����ݡK� �(���gBY��GL�Sev���6�S�s���I������.�
�l��ô��v���vmTa$m�	Ŝ_E63�����D1ka�j2[d繮Y4���iYl#JZLԹ���	�e� ?
��ɻ��I�f�ImЗaź.2�򌌢Gn-�vs'�&��r,�'K����m�4��T�'�%9)�b}����r%�bX����Kı/���r%�bX�����r%�b��y���Q)k6z������Ow���r%�bX���m9ı,O}��m9ı,Og���r%�bX�>�ߍeɪ�f�5��ND�,K���"X�%���{�ӑ,�!�2'�{�6��bX�'{�]�"X�rS���=��(�-Wd{���X�'��ND�,K���6��bX�'��}�ND�,K����ӑ)�NJr_}�{X�&�L5֬�'Òı,Og{��r%�bX�g��m9ı,K����ӑ,K�����i�������o���h�j�Q�9�E��K ��43I��㒜�tGfOaUmLWZf������rS�������oxr%�bX��w٭�"X�%���~�ND�,K���6��bX�'~���Zk�֎:�������<�ߝ��(@> ��@v��wı=�o��Kı=��iȖ%�b{��ӑ,K���׽&Yf���[�fkiȖ%�b{�o�iȖ%�b{;�fӑ,~R"{Z�ӑ,K����ͧ"X�%��!ӹs3�j��Mj�j�9Ĳ��{�&��	���]� �'w��pI�?w]��r%�bX�>���5i��j���fӑ,K���w�iȖ%�b{���ӑ,K���w�iȖ%�b{;�fӑ,K��P����	O�WZP��a���:��f�GL~�l|X�Z�l��C��4��{H���4]����O�%9)���?���ͧ"X�%�ߵ�]�"X�%���}�ND�,K���]�"X�%�㤝=�j���4]d�u��Kı;����Kı=��iȖ%�b~����Kı>�}��rbY�NO7���R��5aV����NJ%���}�ND�,K���]�"X�q�8I$HQE��"�0	�ィAx?�dK���[ND�,K��~�ND�,K��}�Y��ukh�
��|9)�NJr}����O�X�%�}�}5��Kı;����K�,Og{��r%�bX��S�d���3%˙���Kı/�禮��bX�)�w�6��bX�'���m9ı,O{]��r%�bX�� 9��@��>z	ѭ��e�bQ�Ѝ��	��@����\��,�J�1&���nͣ�Z:�����NJrS���{�w�"X�%���}�ND�,K��}v�Ȗ%�b_���[ND�,K�:z����-���rwy�^B�z��iȀ%�b{��ӑ,KĿ{��l?�'�ı?����iȖ%����xF{��P�n���'Ò��K��}v��bX��s����m?D�,K����ӑ,K��w�ͧ'%9)�NO����p\&F&���O�X� %�}�z�iȖ%�bw���iȖ%�b{=�fӑ,K��0A�D��w�iȖ%�b|}!�r[5Mj��u�]j�iȖ%�bw�w�iȖ%�`��=�fӑ,K���w�iȖ%�b_w޺�r%�bX�����IQc,�,lf�v���������Ś�=]]��l��;&˥�y�s�6��b��g����r%�bX��wٴ�Kı?{]��r%�bX��﮶��L�b[�����N�!y�^O?��{�p;\�ff�.��ND�,K���]�!�*EAșĽ����m9ı,Ow���ND�,K���6���L��,O{��iXd�rwy�^B�����m9ı,N���m9ı,Og���r%�bX�����9ı,O�A��\r����y>�����P5�����Kı=���ͧ"X�%����ӑ,K� V	�3����ӑ,K������������55��ND�,K��}�ND�,K����]��%�b_{��[ND�,K�k��ND�,K���@
��O�Iy$��ΞZ�	�,�f�F�:`Nz�?#,�n6�+w�Ɋg�4� 8�ָ;Dj�f�qt8k���9]����q3�;��!]؍�ٲ��È�;>��� ��:�vU��g����]F����-�k��j��̉���#��m��3y��=�֧�z�]�:�^�r�x]7�ɛ�YWe�RXa���E�콬�Ԡ-�[>����� T!�o%�w�3Yd��f`�p�f|v'90e�Z��f�|v���[�Wd��pTßy;���/!y>��rwı,K�wƶ��bX�'~�}v��bX�'s��m9ı,O�C]�-&T��oy>��%9/���{ÑKı;����Kı=��iȖ%�b~����Kı<vC^�iW-*�G��JrS���~|��9ı,Og���r%�bX�����9ı,K�{�[ND�,K��������aV����NJrS���ͧ"X�%����ӑ,Kľ�u��K��	�=�s�m9ı,O?����M2eڛ=rwy�^B���w�iȖ%�b_��f���bX�'~��6��bX�'���m9ı,�>�Ko>��ղ���ͰE��Ýɠ8қ'<,r] �Y.a�[��c�i���f�5s5v��bX�%���kiȖ%�bw���iȖ%�bw=�f��AI�&D�,O�����Kı;�k�fYHk4K%�k5u��Kı;����8:�<l�Ȗ's��m9ı,N�]��r%�bX��﮶��bX�'�wr��Ĺ���55��ND�,K��}�ND�,K���M�"X�%�{�z�iȖ%�bw�w�iȅ�/!y<��O�1ڷa�\��B%�Ȩ�ȟo��iȖ%�b_{���iȖ%�bw�w�iȖ%���Ȟ����iȖ%�b}�k�Ʋ[�ja�.���ND�,K����ӑ,K�������~�bX�'�{�6��bX�'�k��ND�,K�A��̧2��<;w�.<]m��y�;x!.*�[���������m���x�����W����bX�'~�}v��bX�'���m9ı,O��}v��bX�%��魧'%9)�NO<|X��e­�'Ȗ%�b{=�fӑ,K���w�iȖ%�b^����r%�bX��]��wy�^B�y��=�7`]˵6z�Ȗ%�b~����Kı/{��m9��8 D B Hv�T�bn'��]�"X�%����iȖ����y���1����rwy��@ș�zkiȖ%�b{����r%�bX����m9ı,O��}v��bX�'��w��	K��,�I���ӑ,K����ӑ,K����iȖ%�b~����Kı,���+㔎R9H�Ip�um;C�$k:]���4JW[���37 <=�c���ڳ�x�{-���{u�Էh
Ds{���%9,O���6��bX�'�k��ND�,K���ka����L�bX���v��/!y��ךC-[�0�N�%�bX�����9,KĿw���r%�bX��]��r%�bX����m8rMy1�NO���3^R�j����Kı/}����"X�%�ߵ�]�"X�(�0"dO���ٴ�Kı>�׿�ӑ,K�����dֳ&���̺�ӑ,K�;����Kı?g���r%�bX�����9İ?#:T-�����t�E��D��ﵴ�Kı>��HED�XU���rS�������iȖ%�a�(D>�߿���Kı/}����"X�%�ߵ�]�"X����=��k~h\ꅙ��Ͱ#
��X�rn+lF��뉶9���>-�Ss<+t:e�W.�5�u��r%�bX����m9ı,K��{[ND�,K�k��^D�,K�{�ͧ"X�%��ڞ<a5�Y��ə�sSiȖ%�b^����rbX�'~��6��bX�'��}�ND�,K���]�"#�2%���뼗�B�����rS������{�u9ı,O���6��`ؖ'�k��ND�,K���kiȖ%�b~:ww\z�]�)��O�%9)�$��������ND�,K��{��9ı,K�{}��"X�-���ߦӑ,K��c�޺�d�3V̺���r%�bX�����9ı,K��{[ND�,K�{�M�"X�%��=�fӑ,K�����sg�Ч�pj����]_!B H���?�!�gĮ�����`BB$��I��4~��P`@����D$ $�	$!"�X@�����C�lbh@ߘ��qT�6�0J���@H�C����À~@����ʕ$�	U�6~#(<Rr0��~,���/�1�R���C(@����B�">"�"@���c���ϵ����4-�r
Lu;�:�T '[����ml#R�m�l���:�:����Jϖ
�K�R����D`'��m-���F��]�ŵҫgn\����Rk5�"�Z궕�S{d��C����WkVk0�{K�2�֡�N�ma�g�³6*��0IA�2;/5t=�N���]5=��q�n�vZ¶L��PA0�uvəq�!Z%%E�Ue��b�j��C�VU��tjHI�ڹL��"묦ڮژ(�Dl�}��pt�u�e���X}��i��4��	��$�Ɨt�s�8Ȫ�;%VU���lHǳc��9��N9Ϯ��j�i���#ل楸��Z亞�ԎJ���anZ�m�xFl�]gd�l�l���m6ЭAD��c��	��S��V������6u�Ӑ�)m�;[vt�urޚ�rmq���kZ�v"�tᬳ�ml�Ӧ�B���AcS,�
�H���0�cSąUҤHph)p���8v�m\=$S��9��� Z���(��P�Î�� �U�����f�ՆGV���&�F��[8�zT%YX�%el+,MH�pE���g�\e���b��`53���lB]�ў� �b�ET�r�i�Fe���R�+a��N�d�.�ƶ�m3��5sv�N�E�䘼h�	�r5��9��Qv.��q{Al���&���qXE������cp�0�+�:�=hȵ��i�t�Ճ�[�bm ���dv/P	c�H&t����[»D���5��Ϋv M3K[f��Ʈ
�т�<Q�d���#�g;r���A��SC	s��6�Iq��,Z�^���RRVX&x;�rv@�b�i���5�j�a0�%Z;Kv����^m@n�F%%�x)J���X36m.�A�Ԓ�۝К�R�Z#fW�mO3�/&���'Vc�t�N\�\�@y�\73���qA��Urڠe�7�I:�����po�@=�q�����>`���@�~�$�y��Ǔ�?_iI�q�M�K�!������p=��.b fn|�%lZ9����t���3z�ڨ6��������@��Z�a�X6�kL�z��Pr�w.�%��;Zd֍m�c�6�J8�6UP�i^�-��d�X �W68�q���,YXE`�2���C]A�.8vv^&^��j'��/c"\��.�ڽ�����m���t����<�W윒{%��']^Ά�{�3��X,jm*��2i�Y�F54���G��i�Ue]�:L�$íi��n���O�,Kľ����r%�bX����m9ı,O���6��bX�'��~�ND�,K�d4{�]kFM��W0ֶ��bX�'~��6��bX�'��}�ND�,K���M�"X�%�}��m9�ʙ���_�HE�p�N�|9)�NJr~����ND�,K���ND�,K�����r%�bX�����r%�bX�}�w��EGkkr�wy>��%9>���m9ı,K�ݾ�ӑ,K����ӑ,K����iȖ%�b~�G�72�4uz�������>����r%�bX*ǽ�?���Kı>�{�6��bX�'ｿM�"X�r��t��>�ٛ��qf����g��:^�Q��v̗g�j;a�^�u���7jId�eֶ��bX�'���6��bX�'��}�ND�,K�}�M��?DȖ%�{�_�m9ı,O��˟�֛@R�y>��%9>�<�w��6̂� �n&�X����6��bX�%����ӑ,K���w�iȖ%�^O|��߲D��
�s�'w����"~����r%�bX�������bX�'�w~�ND�,K���6��bX�'�����5���WZ�ND�,K���kiȖ%�b}�w��Kı=��iȖ%�b~����K���׽m5V��t��;W�n��E��e� &�W�N�U8����X�M�ڎ%8��h�F�o"� �ν��C�b!ڮv�2)Aj5m��<��y�ϮE�v+���~0�y�;vSwcm+v˻x�r,�U$��v_�)��F����_-�[��� M��ܓ��f懪r��i���ջ��&�*-���W�n�� �lx�Ȱ=ʪ���x�kjZj�tZ��(.��"��r, �e^���jH�H�J�v�I;��)m�h����v��I�[(XB\��c�%�UgJ#���Iv�-;x�v< �e^��� �lx���U���I���H^z��H�� ����>[��O�[xݭE�կ@�����"��r���T�x��+�;ݺ.ʵt]�-]��������:���	'u�>�S�$D�!�����?N�~:���.Jf5�����>RG�l�wnSc�&����1�2X�,��`ݶ�K:$��yz�"S�$8���.W��7X/5�ᖷ�l�wnSc��9K����7�V�!�Qn�\@ӻ�7vឮW<�<����UIu{�x�O^��m��픛��(.��"��< �e��p�;ӎ��!��&Zv�=T���< ��� �ۆ���A\�)S�I4���/ �ۆ��䜽�srJ��H�v���e�C�"��띍���n�6�`g�5��<���n�w<���]q�y"�j�3lrXk%��>#��3�!���$�6�9�
�n��S��e���*�(�˼�s)m<��9�GcE��KE!a����v=�&�n�ζb�$ek��j'(l��]F����tR{VE�d2��<�n2��ö�iq1vM8��x�ZP���=��P���Ke�<��.����=�2�40�m�u��ze�k6�l-��4Z��@�����<�c�>RG�l��ۡ˲�0�VZ�IـE6<�$x&��7v��s�Z~����LƍUw@�}�� $�x}�%��`E6<zŴğ���j�7{��w���s��/O<����;"����]���)#�>RG�Ix_��@E��jK��d�D�Gi�9���a��2qS�jS"�J͛%��̥��qS�y|�̀|�� &�x��0�㥱�E7i2ӷ�|��/���W�9/ �v�E�<�Gkǯ�b�J��v���� �ۆ��)#�%lJ����i����w�n�� �H�����^����vU��]�j�'f���9]r[�	6^��������ׅu Y��,6�����l��(�d؜mv�pv��̞�����;V�L�����u{�x$��n�� �H�	�k�v��݅��j���/ �ۆ����{� ��o�c�E��q���7v�E���9WEU7��b*�
h������w}xk���c�teݘ�y���{� &�wnt�t�R lӷ�|�� ������e`vG�M�)�t*�v�RT�BtN���N���}�go��M7�������2�bR�*Vm���=x�e`wf��({}���=�{lf�֭KU�z�eeW ��<)#�	�/=Ď��]��݉�Jݷu�yo���� &�I2��]]�����m]ݼs����< ���I2�r�TUs�r�sy��)r�������[��� N��\�\������@���<)#�>��-ZN�4�&���:P�g�<,�s(���r���y1&�&�	�&���и����7v�Eݏ �I�_ =���[R�I� m�]�v`nǀ|�� 'd�wn��&�N��j���4��^�� N�wn]���R�Y�M�
��x�^�z�	%��69�����9ʄ�����<���8��-KU��۷ܞ�y|W��$�yUU
�h4"Db�p���fC���l�2(]��ҙˈy��]k�K"Y�j0u-)�[����÷=W#��5��ݬ%��lJӸ�׭������E�v���4��m��E�h��1���<��	2duv]���d1P�c����n�n��;y�l�
�sm1�;4�������:��!���WS�	���p�]���'�mv��O�+��K(�X5�rrr~䐝�^��M���1��;D��֞$���u랞����d�V�-�1�ubm�iRWi;>�Ȱ����/ �ۆ�Ȳ��[WJ�[����|�� 7d�wnc�`��r����v[��� n�x��0�"�>RG�}����IQn�\@ӻ�$�+ �r,)#����;]����te$�� �=� �\0{��	$��6%R���uhA�ɕ�ys͗8�g1�܉`j����5\�o#�E�Ut��T���n�#�`���$�+ �9!R�Y�M�
�	;0we�.��W9T�$��;� �\3ԑ+bUt�6��tڻ�wx��e`G"�$r, ��x��.�m۶���N���X�Ȱwe��p�6He]���Е��X�ȰUs�l����`G�`����}[�v�Ҭj�Ͱ*,��\�eҁ�4r] �!�i|Z���qk�m�Zp컳�	�׀n�� �=� ��X{�[#h+wB�n� �n��X�b����6�R�P����(.��>�b�"��_��r����e��Zlʆ����
kl8D�:)F��*�A D����ى�:]Q�5QLA��k@\]gЄ! �!#?"F�����M�ڦwa̩��� R��b�(�v('E?�uDD8�߀<�����g�}��?~�]0�U:[T���n���we�m� �=� �.U�T�@�i�����$ۆ�{���@�V4ݻn�t*����c�2���m�'���{���i��/e�X!���3��i�wv��ޗ� �=� �lx�����ue�.۱+����ȳ�<�<�I��$ۆ6C)۲�
��cN���we�m� �9:ͧ�˻V��;���/rN��vnI��{w!a?E(dX @]#������s﮲w2��n�\@���l��>��E6< ��܌�!y/+�n�$�	��C�ES�{�t8.x����6��{ls�'UZI������w��`M� 7�/ �fV�)Wv6��6	[Wf��{��	6e`G�g����^�U�I��I�o $��M�X�Ȱ��������vX�wj��z{+ �9#ذ=U��~��^ o����.�jݍ]�wX�Ȱ	ŀ�/ �fVک�R�s���UR��$y��6ņ�\�ј��2����T�*Nl�/fS5��	�i��e�g�c�rN�WY6�onK���1��Sڐ�MVCݴ�4kN���!����{T�ms���Y (R=&I��-��t��� �1W:Y\�.�At�_O��	�W@4]�'lU�7s�2j��K�˵��&vu��v�/l�I�v�u�	u0�Q"䓓��9�s���<'E8�K��T��H]��H�dv�Ҁ���b[s
��r�u޻'ftZ(�+v4�|��, ��x�2�W�;��,��O�,/�v���wo 7v^&̬�.Sc�Ur�6Oy[?6�T[�;wx�����}%���9ʤ�����g� ��KMT���te��W�S����~���`���$ٕ�}�U�Lh��� ��X�r�UU��\����������}%� ��S����Q�����b[��\�A����n��:6�Ɔ�T�N&�@��B�f�we�l��>����A���J�*feڣ.��z�~󳽒rY䆀J^�?������'���7$?~���>_<�3Dlb��V՝�0�"���H�z�z{+ �!���i'`Z�e�f��we�l���.��� ��S�h�[�llN�����?W�=�|}��E6<��¾�U�`4��
-��4!�c�ۯ]Wl�vx˫RX�����7c��W�I�+ ���H�, �v^�ږ��We�]���.d�`{���2��J��m���+j�ܓ�s���O߾��1H �" @A��/�w�7$����܇�%YLI�+nݬ ��/ ݓ+ ��p��9K}~��%H�_=M�N����� ݓ+ �vg���?y`�ٺ����=���.رT���֛��y�y�����^�mKrK�$Zb+-ݴ����i+��� ��p�;� >���7d��;�,�n��텦����;%� ;ݗ�nɕ�}�p�'Y��+e[�ln�������2����\0��iN:T[�wx�[�s���ܓ�s�����?��_�6# �4�?OٿkrN����M�]�����Ȱ��vL���D�O�BM:m���MP�m��q)I�- �YV4+����`ʼ�!*�k�S���v|��� >���7dʺ��wfV���Bj�V
ݻX�v^�&V�ve`�E��{�ʦ�I�!���$�����V۷�@>}�Ǡy玾V0j��U�g@��2��p�����2��)�˱զ�����\0��x�7$���f䟸�
n�����˿]p�Ul�+g8ٽZ�9���&��É���ڝXMn�n�&.,��P��&��{tݜ�T]�;k&����;!��0f���^�fV�F��-�ݤm���֠��x��y�`�b�-��� �����$��r<I����^mnîi��g���݅�x.�^'Og�:v��g�v��v�<�	�	�F\�+�T�3B+���9����.���J�ۊ�H����hGv��Ug�x��&�q̜��n<��B�1@�,�;]-����=vL��ɕ�v9��)Ң��E .���2���+ �r, ����y�I-?{=n�c����t�=��v9 }ݗ�nɕ�}�U�1�4	X��Ur����� 6O^�&V�ˆ�A�J�j�V%mݘ��x�X�.d�`�UW'�k�Kg�-pB �Zf�U�+�X�J�"�ݎ�6����I�V�b��tu�m]�w'���}��vK� n��&4:tcVڶ�� �K��2�W.��Gd�`{���2��(�v;�۱2�n��Ȱwe��W����;�_�u�Rƕ�t��t����/ ݓ+ �K�򫜮-�q`��j2�*-�$R�� ݓ+ �e� �r, ��xʥ�T�6TMq����j��a���;u�v*d�է'E�jiY�e�c-�Xl3�}%� � ��~����V�R�{�m4�V+� � ��x�X�.ܒ��&��bV��`I�ﻭ�>��ٹA8���/�"�iP�D&&	s���?{������]m�jؚmT���e`l�`�E�ݗ�n��Զ�E���u�}%� ������׀nɕ�N�9��*Le��Bm�t��8���4w��g��j�bc���'���b��93�-p���>�������=vL��.�6��+���-��ݘ���ܪ�x�6{������;%�=UIe���$�)ww�I�e`l�`���/ �i�]Yi�S���ˆ��X��x��pݓ+ ���H�6`��v`�E�ݗ�nɕ�}��l�{�'Y�hX�F��Q���k����p
��76�wj=��.��\�v�	���l�� ݓ+ �e� �r,��<k�v�[�$��߾�wm��_��Ȱݸ`��:u*�am�i�`Ip�;�W+�JI~0	=��I�R�MջWn��0�"�7v�nɕ�ꪥ�{<`�J��v5N�ln��`�p�7d��>��rO����IXDa F@0M��d#��c��cHI	,##!FB���0�P� B$	"BBH���!F2���#� �H�B22��,-�$#�݀! �!2�S�F����$�B	!!?qCi��`^uG��jHut!�D�F��@�O�Ȑ��m��#��$᳦η��)��$�`8&���*&+�!���E�H�X$?#�$�!ɤx�6��A B1HN���������@"D@ 0`��E�I�"EH,J���#  0Y0��|�!� ��S-��|����t�$M��%[�B$�CBk�6h�0b�B;�t��F��E :ҧ`�����NHb,!c#�$d�� ��l�b,~��	�"HD 0a"�b��#�$B� �+!�#�a�0�!�$!$# � BI$dd$����%$��$��%%�	KJ $xK	C�0���R�!H�2c!��1�0# ���D�`B0d$#��$!H@���bA�`F ��V
�E������!��;/����XJJ��˷�z�3Wiۣ 3�@i챭�V�[� �-UJ���-�3�Bv[*ȫc\�ٱa���ٻ:6щ})�+k:6.qE�b��;�T��kV��S�V�e�{cv�9̦�v@gk�۝�h�_Z8ֺUᶮ��/S�C�:5a�o^��^���Iӎ��SN�u;�<N.���)�ᣞ���k��:����R9�U�"j�]����*��k�4���Zve�t۶S�S�M���n�cQ��	�2��M�Ma��b|��pGHq[I�ƛ�2�n�q����@^�eM���ZH�>�ɻ��d�f�Rv���Ʈjum��"]�����g������D+A�ηh������F���@p���q6��ƒt�t�] {@�M��]�c"q����0�cq�����%-Z� �4p�h�Ssa��9��m$i�:���"��u���q�i����T��ۘ�d���떔��9PK���]
��
�Xf�d�.-�l�e
����*r��\-�*��H����V�[
�vD���Y��[�5�V9]�{X)^��n��:����v0�U�c����4Ҳ�Óve"X�l<�� ��ۖl��&�CJp*M�����u��Lչbc)�RE��r��z]�ZVݛ�F�H��r����E�$��"�jL�&FwnX�z��2��*}0�y��ڵj8�ȮMw@Ύv�w�����.,�j�6T�ԡOF����|��.bv%u���r�5����t�9�3�:B�S�ݰ�5����P]�k�[4�qj3S��37=d46ջ[�Zu���le��klb�ӁZ,Xδ���3�ٗ��.�z�$k&�[Զ���U0(������K�%'U��QY��K�� H�M��`:�%����4�A���i�Z�(�j���G�p�m ��R�m�"&T�ڡL�tY�-Q�;Y��{f٩6�5(( ����6 ~ ���'4��A�D�/u0A6 e!��+�_�)�C��8����c7�&�&V1�<�eڈ��.�l����gGb�U��sv�WLl�AX�Ÿ�æ�S���v�Z��^(2t�n)C�vt�;���),$��B��su�am��!{�ѱ)��0�s�0N68*�K���u�T7b��mY\[#���i��-"ۈ�$.d.��&f.uwZ.��N�Gnts�&�cH��/huc��;t:urh�6V�Nq^v�ڦ��L@M;iS$:C h�k<k�;7f���bM�M�f���)E�0�̬��Ȱ��0�X㫲�;
a`[��>��v9��vL��R�%6�@�%b�0�"�7vᇪ��)=�����>��Je���ջX��0�2���`er�eȰԊ�J1]�˦��wf�&V�����7��X��0V��+��H�ۡ7eÍ����з �e.�OWg�:�م�˳�6�3C ��2:wm����vK���s�\���I�e`�{(�mÚթ\��>�s�ӓ��%�`l��>�p�'Y��]��e��$�`�p�7d��>��v9��R �`�E�0�2���`�E�n�� ݈��]���0�-�`Ip�9��g��d��Xv�IR��t]SM9��Ҥ��m��J����=�*gi�
���m��V+� �r,��vL���A�VpN��b�n��ۆ�&V�ˆ��Xպ���6�쫦աݘ�X�\0ڮs��U����A�w5۹'��0vP*p���m[N��\�.�g�|��wv�nɕ�vi2�Whn�&��-�0�"�;�p�7d��>��w���AV�X$�m�[,	j�0!c�(ۜ��Y�v��A.�ŭ��Z��6:.�m:I��7v�nɕ�}%� �r,��Ri*-�.�ݘ�Y��9ʮU$w޿��� �ۆ�cU.�Wt5E�n� �K���X{����`{�Xܥ	M�&�+ـv9��vL��r�UQA�;t
��yɹ'�;�D2e`�V���7v�nɕ�}��v9V�'��y�}q���������;K������{[6,�{1���6}�R�I�TںN��	=���Ȱ��0�aJ�R�&�[v���>�p��UUč����_�vL��b�T��+�vX�ـv9��vL��.�6J퉢�7Bv�ݸ`�e`Ip�;%� ��l��H-ة�-ـnɕ�}��vK��� �wiJ	b�n��,N��!ڂ;��������k�bì�u.�vp���4�c.�K����FB��5��ZgN��Ў:J�N!҅eI�%�8��9��6�F�'����cY2������V�VTN3�m�:c��t�Gmrv�F彶VYt��Ϭ縢�����v�{hKn0�OhWe���㮸,]v�k���k��H�d3ma%84x��j)�c�c
��zR��6�I��:3ۡ�bՇ�])��{m�����T5E�n��;=~0�p�;�p�7d��>�*�6���+� ���v\0�\3�RG|q��c�
v+J��6K�nˆ���\0�u[b�N�!�j�;� ݗ�.c�`�p�"��*mF�i�iݘ�\0�"�7v�nˆ��a ��;����E��{Y$�&cy�ȳ�H�V���3v-ź�)K��]+��+�>|��n�� ݗI��}}:��磅�l8q�.o@�ۆ>s�G+��ʮUT�D�p�6K���X۶�8��T��[� ݗ�=��[�_�d��h�妮�j�Wf��d�`�p�6K��)T���Hl�]��p�7v�l��.�j���f5ٔ�
���K2�46 c�����bǍ+6vR���o� M�b
�m��E�l��n�"�;�ԭ�Q�wm��t���l�uȰ�E�M{�)S%��HVݻ�0�����I�s���� �+"��-*�`����n����`$YJ�,Wat�+v���{5�X�&V:�X�H[��%V���N�5�X�&V:�Xu�V�=g��-\��X�I�a�3vD�Q�)�h뭚�.� �fNѺ�^�Q8���¤�wk �d��'\� ��� ��,vR�Rn6��j�Wu�N�JH�Vױ`��Xr�ou��!�J��`kذ	�b�>ݙX�`8�j��ح[��M{�ɕ�N�+����b�7j$�b�M
�t���}�e`�E�w^ŀM{�A��";N�m����x���vs@PnFZ������k�H��=k7<L��2��I[un�	�"�;�b�&��ܮW�;=�{�YJ���v"իWk  ��,�+ �r,c%8�WI�l�7Bv�	�b�>�2�	�"�;�b�;�أ) �b�E�����9�]��V�~��>ױ`^ŀn�V���i�-RJ�	�"�ſ���ܓ����IϾ���>�U�c�̬��
���XW$˅;Bk`��sb����|��k\V�i#Q�.G��kk�j�@������{hۏ]<f{B�6�;�f��"���n��L�c@AӴ �a��w�(����/�K��v��Xv��6`ao3E�\�,��c9��9�� �ɬW
�N���C�8�t����W�R���[��5V�����9gVނ|��[8���@NΡwgokc�Rb
�;K�����#�tW���v���+z���7^ŀ}�2�s� �x��-$�ح[��n�� �ve`G"�>ױg���G�y%c��S2�7k ���'\�s��]�y`�y`H�2�$��V�� �r,��,kذ�L�d�)Rb��n�5j���;�b�&�� �d��'\� ����ʵf��Y�*����	<�X��m�suvM7�du.۞WeS]��r��Н�kذ�fV:�X��,�-�Sv.+�v��fV3�#�!�u�/��n��>�ܓ�fŀn�V�r�j�%wX�Ȱ��X�ذ�fVڥSc�am�wk �^ŀM{����'\� ��UhI�;�v�	�b�>ݙX�`kذs��l�Rt�����.'Ls��v9y�)����Wk�[�씉�����x�7Aqݷ�{+ �r,�{5�XR:L�6!�[��u�N���� ��,�ٕ�I#�T��ݷi��Z�X��,kذuڧUg*r��
�+��\���4
T����]�^��P4+����I����d�����!�-(HS;��r�wP��$9�X���R�H�XX1 �+@h�!���y��d�w"}��&w@���l���8��ȥ �M��X!�x�1�M����Ǩ�ELUM�π�@@?
u8���`��8��h� ��P����\J�r��;�X��Y��J�WM�l�7Bv�G<��fV:�X��,�-���Qn��bV������'\� �^ŀI.�.�T)];/�ۄ�8<V(N#�{nqy�ݎT��3�Ҹ ��fܶˮ�Q��՝�7�^����$�z�����J��6����Eݬ�{z�=�_���e`9�snr�L�N�jݬIp�'d��$r,kذډ+��v첮���v`{��UR���V�?y`^Ł��
@V��(Z�P:`�s��9����>S]!S%[��I[wX�E�M{$�`�e`�	:�K��B�V#����K�����D���+(+JW�rK�(��M78�b�k ��,Ip�'d��$r,��C�Zi�l�7IݼIp�U$zOe`���dy�q#g���Ш�b�ZH�f�=��H�Xz���^[�<�}}:��J�|�`a��3�y�`vG�l�n̬�["Cam�wk ��<Ip�&���69 >W
�ʎ+*ӧV])����˘8][���^غ��f�2�<nyBi�Ė��\wj��%�T��S3�V�Wi=�֡P8��`��2b��{k�#%�.�O���%��5t*����i�T%tb�8 ;$�6��aG���û�`De]s�fU��� ��f[cD��N��Ӻ��=qrɃX8F�ڔq���G]a{BB8}s��v+��׹'$�]I�E�:��B�&"1��ld�!>Tݝ�m6��tsّ�C6R�f�̱m!N�v�ށ�K�Mٕ�lr,.��	�W.�v�ꮬ��v`ve`� ��<d�`k����i+eZwX�"�"�ǀl�w|��~��٥Ô�SU�oC��_w��Oz�`�2��E�wZ��-�l�7IݼIp�>�2��E�j�ǀ|��$*�X��T6��l+OcTq�n�Q���.IdmH\���LI�J�S�rn��T�J��0�̬c�`���%� �e+C���w@�T[wX����$P"�IW��&�[����ɕ�}T�H��[awk ��ǀl��ɕ�lr,aǲ��6p�b�Wo��r�O{<`�{+ �Ȱ��x�D��t�*�V][�0�̬G"�5wc�$����C��𞛥���6n5�ͱ��J��3�v�d�5'gWf�-��+�m1ix�)6�M��b���~��5wc�6K����{+ �/e���]��j�`��竜�'�~0�{+ ��Yꪪ��u�����6�.�{���9߻�s�y	I#~@!V�dP-N��F "����E�� ��dE4Qn�H��[�˾���	��,Wv<M�X�R���ݡ�����	ŀj�ǀI�+ ��e`J�E1�ݗH�c)��6.3RW4��P����nz�{�t��`Q�un�MM�Eݬ��&̬�ɕ�H�,aǳ��&�R�]���I�+=UU\H;����XWv<�������Je�L1�� ���^�#ذ�Ur�ճ� ��e`�(6����-
ۻ�;ŀuwc�>�2�'�&�*_��krN~���I���ƭZ�XWv<�+ >엀n�� ���2��T�$�m4��nԫĻ�A��E���z m��+���b���m�t��[����ɕ�vK�;�b�:�����)�*-ؑV�j���xcذ��x�L��J�M��t�M;��&�� ��Ǉ���)/o����z��U$mR���ۢ���ݏ �fV }�/ܪ��\��'�9�+T7��]�M�X������'���ܓ���srO����
 ((P���J�j�U
�%��%˭d���c@7\u�S+:����1���M��r:��i���]t1�rr�4�����첷7lV�½h�Ɨ�7b��.�hDڡ(뎙
tE�[9ݵ�Kb�VU�c��Ge��8����� �-���X��! ]�ק�ڻb�tʶ��K�ӹ�:��mQ���rޓy2nU�����l"{'k�0�Ǎ���ŋh�I�b�#���"9&�̷�ֳ5��������!���sص,/��#����c��m
dV;%-У�]��cs> y���=�S�=s��5l��+�\���V�=@鴼4�at��w�l{{�Uč[<�	�� ��^J�U$.�E&&˲�SV�]���&̬ ��^#ذ�Im6��;���'v��2���xǱ`]���F0T[�"�*N���xǱ`]���2um����/�&�Ĳ����.�pm(�������n^�v���vc�"Kj�n� ��,���fV�d��;T�dcM�M��Eݬ��}ZW� [�� Vȉ�_}͛�w��f�w>����;��+T�TR�]���OOe`vL�cذ��xڀ��
�[c�um�`vL�cذ��x�s��z��`o���K�l]+�`ŀuwc�6l��>�X������X�
9�-�K�-�����7ּf�ݜEr�u�\`wT�u�t���;SR�$��y�6e`vL���68_��H��L~b.Ɲ���wo �]X��V��� ��ǀvK`�%E� �C�7$���f��}۹�� � �P ��������7$�~���9�JV���'t
��5�XWv=�?������}�pܓ৽��r�6�]��:����W*��������XǱ`����C�n�Pҡ�3F�j��n���L�,��D��"�M&���Ҝc�N�v���fV�d��6=� ��ǀM�B�`�U�]ZwXݓ+ ��,���fVz������y6���X�� �s� ��ǀj��.Rbn�]��Wm]�	J9q�M� �W(��堨5�� �@A��T:'�g�7�1�R.Ɲ���wo ��<�\0	�b�5l� ��Jr��P!6�Q��L�U�as �a[F9���h[������*f�V`�rZA�����.�b�5l���s� ����;+ԭ��XX�]��b�W9T���<��.j�II���v�[#�6=� �cذ	]({8�l�N�v����Xd�`=� ղ<v�%h�����j��ـvK���X���6�o1=@(� 4: �I�"I�II#!�Br� � ��� @� H� �M�C`"�+�	=�oA@c+�π�

f������$�����ām�\��e����k�kD&�&ߒ	�$����AP�.F	��:%9^@Y��9��G`}��� N
`��	S@ ��^"h�D��_�C��+�1�F��9���'ȿSQ J�E?~��%@H�$Ua	$��!��Y*�D H�	�B�h���U�Lߗ���~m>�JJ �uYV^U��Xm=��HHs;]�˻ +��d��V�U�<�0���mk��z3-B;/Z�3�W�
�X-���t���-p��,�*�r��v��e��ub�N�Q�h�Hԩo^i��gd�UR�0p�A6�ۂ3�׈8`�Qp����<tꤸ6Z��rr���`���bG���m�*��ʅ����u-���kf�@�i��2`Z-[@�^5��PH�k�e���k��sQ{�Uo] �L��r�@�8Ш[�1��ɸcP��be�q�Ti�xӶ��`u��`��Dc~��L��ܒ��Q>�����\ĝɵ`ЩA�m�ʪ [�:{[�c<zeUj�Xۊv�x�,��u'52r��m�.�g��a�v���Yv�5�d��>��L��]��Arv��^�h�<���r�8�jTul�6rKE<�b����YҶUkƨ*�*����LÜ畣�x���W=���(�\E��[,@�i��vq�c�F� p���{0X:�m+�;��%����0$���P/a�l^Sj�@��6�PY����wc�[:7g��pusTR$�m����(�Ҋ Uم[���n�!;.}8#gNq�Ŷb��]�����<��GNè��QG�񎅴4,�kr;3���i�3���SJ�4��d�$�9M����=��Fm��0�����H(�4���,�t�gp�s���V��i�"�^2�K��L$m7Y^�d  1�λn���NnC��,�VG:���f�ڤ�6�N�r]���Qf6;3ǧt�vأmnWl����(ǲ4��MM��
�g6x8U�[����%��[�-y85�Fm�$( t�N~>��e.b鋍�H��%�y؈�:Ͱ�us���K]K˶��;5#%�1�뫦��]�n�ɛ��f=(��J�K�Ks�x��@\�/,q�<�C6�]T�n$)0`�9ZU*62����qΰq	3"�*��k]����'��d�䜉>O ��ʿ"�� �����;H/�?�|�|�'i�>Mn�D���U& ��B�&����T �;X��*�W]����KJ�nT��r�-�i�׷N2r���ѳd� ��TT�skj$���W+4�Gn-3�\m!�cp�m����,�ړ��h1XTf�6g4bPt�y�z?{��&�	���k�s=�tq��������:��Q��CiSL�Z�����V�Će�0x.�9NNn�ev�/bSn^r��'l֪�mZ�����d���AcUe&5�f�Cj�p�:�X���m� �{�e��ӻ�uj��j�;.d�`^ŀoe�j"��Ӷ[N��6�vK��U�%<����-�JJ��"�@ݘd�`=� ղ<M�`mJV�]�;���Z�0	ŀj�&�0�p�	�R�[��4�T�`*��ͷ�0�\=�r5�mt�w!�g�j���Ў l-�.�`�G�I��\0	ŀJ�O\�RuE;ڻx�p�>E~(%@�)T�Dq"�D��3,׷�M�=�;�'�������'���kEYa��@�﯌cذ[#�6m� �s�o�
�?6�L- ݟ��W8��y`Oy�6��s�K}��{b�P���wv��]�v��"�6m� �c�z��9��rd͎��ԕ�V�4-:B�ǎ��:���Ѫ�s'����R�9ٶ����ӻx�`�``�b��������/2�E�*Ҧݘd��$z9�E=�Nˆy#��J�O�an���i�`�y`�G���s��\�q���vI��mR����������dxvL��L��X���cg
v+�v��X\�W9�%��r,V��	]e)�y��b�ر�M�Y���n\W'��.�3�[l�(��vbN�3��s��K-�vD�u�vI��w\� �r,�&V obSLah��.�`�2��00��P����mէnݘ����e`�``��oe�%�WcWm[N���e`�``�E���UR�Q�W[n��̏ ���J݊�iYwu�vI��o\� ղ<�L���@��ٺ�'�&�6�9�m�$��ہ�6�nJ�<A�f�.��+�%�����o<�V���Xd��J�bI����X����s�H���{����r,�8=�Ll�N�v���ۆ&�Kq.��,����;[Q\�e�e��N���M������ױ`�R�SiA�0�U��X�nRG�o^ŀI��>�9���j�@!A:M�3�5�"l��\�9�l�p9\�f&�l*T�P��\:
:�ۖq�<ܨ[qr��j]���k\M��{�X�p�om���Mm��L�rc6bE�ck���[��Ld�tC��Ǆ-D��SWl���ڄ�!Sp�<�'h69#!ԍo]<��l��AH�m�K�\�aj��������#Ьv��&v汞�]�;�L�MY�;%�Ke������gD�,�YhP��SY�j�l� ��a2�GQ����ӣ�_aA��2�Zk��m��rt��������`mİ��0	ݱ�4��5vձ����{~�q#ޗ��_�/}���rp/�|o����B �[~��%�w��E$xz�X�R���n�Ĭ�;K �m� �H��ذ=U�R��y,U*��t�l-:ـE$x��X�q,��g��iHn�#)�ܻY�%���ݧ`]����̌�u��v���m�o��آ���<�	6�X�nRG�v�yjo��Xk����?>[�$�%T׷)#�5wc�"��P��A�L-���>�p�"�<?Uq(�y���%�M�ei��c*�۷f�����mİ��0	ݱ�ի����v�]��r����y/����"�<��ѵP�t��H_9^'c����6�^���)�x.!�cN����LI�e��ږUe�m�.�����@���0RG�ݗ��W9\H�R�	�v��J�-�X}/��H�{�����J�bN�v`������w[�&Ȩ@�BG��;��5�M�� �ZU�*�k��MZ�x��X�\k �m��9�s�?{� ڞV��;V�tZ��wk �ˍ`M�`�� ޽� ��Ҡ��t��AiqY��i-��i��Ŗ;Y�=���W��v�Ҙ�P���'V���{zT��ױ`�q�lS(CI���U��n�T�窪�\����y`}~k �m� ��L�RwVݺV�ӻx��X�\k �m� �$xdWSE+��H��wk�\S}�k ����rO�{�ܜ�B��r�
d?��S������I����¬J�-�X۷T��kذ���Ң)�X���.&��M��NKbVԈi���.ts�e�T:N�09j��i�4&�ӡݘ�#�5wc�7��X�n�9i�6��wcVݼWv<l���ۆdy��I���j_r�����=}��|�n]�����H褆҂Le��ݥ�}6�E����������}��{���\K�ͬj�'@��<ܪSg��==~K �m� �+�<�5U�3_���_d��e�l�g�ny5�P��m���z�M�%�ۭm%Vʼ��������Ÿ��k�N$"�Y�ݝy�H	B8�8�{]����1���Ǝ�R�k���@YNǣN�3c�uv�AA�\��܏kB�ؗ4J�P�����QuH3�pn`56�ۑ-�M��78zu�,5�.4i �����HXQJ�Ae�
lJ�Ymf�VPU6MU>Nr�I��G�NϚ�}��t���;c�k��l���	p�sl��_��70��ڬl�ߠ���z�ۉ`n�?�ʪ����X���Ԇ��wj�i��;��>ݸ`^ŀݗ�vj�F�һ
�+,N��>�p�&�� �ݏ �ۉ`���ēam�n��	�b�5wc�>�q, �l�n�V�&pwi����j�ǀ}6�X��x���R����1Gyȸ>�g@#;�ݻH�'\m��ŀ�Oj�%-�ϴ&a����������f�o պ���� ��:(*��!n1����|�u�{g�s�)�w� '}��'v�Y��9\��^����2���+�=�y���߼z�ۉ`۲�	�i�U�����ln������&�İ���=T���y�Ɓ�������ߞoC�o�s�]~��O<z�, ��H��˩g�<�F.y��v��V J6	��`X�U`�b���m+�fء�K�z��ǀuwc�7�b��;���8�O&�M���wo ��ǀo^ŀ}ݸ����-5)��C�M�v��>�ܓ���m��]��D�I�M1lI���$�HO�����h�!.&�0�Ag�t#;�O���������'$!�0G �$�f:@"5Ln�b�b����#�(P��i�	�ͻ&'��"��!�8��# "���Uw(b�1E ��a0�~���Y��v�]�(��a q�/GB�;So�hw��T� O�]��uV��T�<TB�~?��/�^�<�_{�7����l�E�A��@�����@��c��K��9\�R��uH褆5�0��ݥ�|�c��K�7�b�;ݘ��-��n���=;oX�+v�]oC�k�i�8�֖ݽQ3l76t�ZN��Uj�wo ;6^���و�9_ ����&������le�w�ݗ�w�1�lx��xdWIJ
T��R-!;��>��F� w�/ 7�/ ��[#��vbVX�р|�ǀuwc��	�ׁ����� ��|b�0
	(� ��'q{��o�	���c [p�v��ݏ >�/ ��1���s���>�gR
�3F�����Z\pu%�(�h����f%�U�����	q�6����׀}�1��|�T�x��ޕ.T45WUz�߼�;�;'� �'� ov^�uQI5R�L,M۴`�e�f�����;�|��O�y�GV�X�U^����/^�� =�׀n�X;����`�妝�-��v�we�����x˲<���%9�+V��I��:�89�zn^|�Ab�ӻt[����p������Z���V�=`\6�v�)T�lu��&��5��F��v�K kg2��F��T�\�F����t�+7e�y}�3��~/����'e�r��P#T\n�h^ь��#�8v�H̰Mķ[����j�����I-�C 7�+��v���M�'������Z�U-����TH��O����>vj)Ih�:7LE=v��qm� �׮��-=���`�n�v^CL���,��F�e~瞿�����=��?�s� ;'� �
������+*Ӵ���xWdx���ۉu�䜐/�'��� Yn۫o����ױ`ݸ� }6^ޔ�2R)>�6[��I��ۉ`�/ ��ǀv�R�v�CW`����İM��uwc�$ۆ7lN�_�C؄ۗ��;��2�X�\��j�������$�F��DLj7YA-��`�/ ��ǀI���İ����i����r�����ߜ��	����� ��q, �e��c8�v�WN�v��#�>��K &������T��R-*��}ݸ� I��{���#�=ʞ��Q�wJ�Ĭ�;K�I�����$ٕ�}%İ)��U��ա4�J�@Aa�a�������$5��Ƒ"�e�u9,0��	�-&���z��2��\K $�xzq�ڔ�O��Nһ�M�X�\K $�x��y��W)!B�[V�خ�N�N� �9�	>�<�t1������;�~�����	�	5AH.�����;UT�{/ >ݗ�E����>�?y�M6�b�j�+�>�߼���z��ݗ�n��>]�J+j˾+.8�&���$�c	�q2V8"-��j�	�s'� T�E33.�Ь������7@��1�7e�]��Ȯ� h�wj�iP���ٌ�	6^�ݏ �lx�j�EN�wEҥnһf I����xSc�>ݘ��U�T�����nӻ������+rmG@U  K���έ��kr��^�R��7m��"���\�s���ޞ�����9�it�N�܊㍸ri֚3/ bZ�e���ʣE�����;�f�9��ٸ����c�o $�xWv<.���E�2�][Wwm�ݗ�uwc�"� �\��#�e�Lwv������<)���K�����=x챑[wCj�
��N����� �~�x6K�5wc�;"���ڠ��ӵ�}�F�l��j�ǀM���I�6��Q�8 �$�2ޟv��۶�;\�;�Kv����0��Ռu��x灭m�u���yz�Yv�P��&n�p7j��m��\m6��d5'oAe]��AM�u$�2ʓ�"Ή��ۭ�&`���8��uuW� �Z�2�1`2�l��u�t�V�4�x�P���mѸ���(`�
C@P�e����n�E�A��!�s)\�Y�
m鸍Wڦ��M��f��?��Ϲ	�9?N����-�ɭz�'�&᪴���%��(�
\�f͸��ϥ#��M�]�8�i} ���x��x�"�>ױ��8��[优!�-&�;��5l��&������/ ;ӉmN&��7m��&������/ ��ǀv�WI�]��V��n�����d��M{��Xf���UT��ݵwm�d��M{��Xױ��'�'���-6�hL�*F벩����;Al�u<t�ru�;2v�F��v����Z��w��5Ȱ	�cx6K�'v�8�t��t+c��`��n���D_��DTM�OG�7����^ŀvEpH)�[���V��k�� M��	�b�&����I��v�V�7m��/ ��,k�`^�����A�1�-&�;��&�� ��Xױ� �%���r���R���H��O*��9ps�g���Ywg����e�̈ܠ�&����S�v�n����~Xױ� �%�^ŀv�V�p]��V��n�5�o &�xױ`\� ���J	1�ӻjݷ�d�G�d�O�TRg���ܓ��{3rO�}{�&髫j����=� ��Xױ� �%��i�2˶��
ۻ�0	�E�N����/ ��ǀ*�\�t��z.L�BmCm+�`�[�E����v�R5��5�)�M�5��n|L{X�ӵ��y� �%�]��	�E�n��#E��E+v���l��uwc�&�����R�IA���v���]��	�E��.��� �%�zq-�I�)ӻM�v�<�/޻�~�wٛ�N���rok�D "	��:" ��7�f�;۬'���c���˷k �^���K�:�c�7\� ��r�z�q{�v����ҧ@����OK)�mY�)�<qR�F�A���#2�Ќ�l�i1ӻj����޼��,k�`u�o �u]JJۦ�E��ww�uwc�&�����d��u�9NӶ;��I��7\� �^���K�:���خ	P>+v�X�ӵ���s���޼����X�B��հ�)[�ݷ��^}���y$���RM���fnI� ����T� EE_��EEZ�**����� "���E_�E@Q?���P��T T#BAP�	BAP�T!BBT T"�T"$�B
0T  �P�B(�*0T �B*T �T"T �@ dBAP�T$BT#B$�B �T" �P�(DT"T  AP��B,B$U�T"0T �B��*T"#B(0T"�BAP�AP�T �T!B0T!B0T!BT$BT!B00T �P�0�AP��B
B"�B
)B�B ���P�$B)B@T$Q0T @T"AP�P��P��B$���T"��T  �P��B#B!T �E�P��T �BEBT#P�@T!@EPH� ?�*
��������**�*
��PTU�**�����@"��� ����**������"���QW���e5����F��� �s2}p��    (  @=@  (   $ @�    8HJH�BIJ��RE
(T(��(�RTH)I� QH��� J��)"�U$�IHH*(      � P   
�
}ﴜ����{��,��y��� �����n,��&^���W8��y��}��K�g�� 5y`��� �w�V-�Srö�3l����@z8�rǻ�8�� �  �  �b �@�9����79��� �//����nMqj]�6���0t�ĦO��ӗ�k��d� 9�Ӗ���ɯ/W�T�}���n� <��{۪�t���ht����x �  �    @ <��U�@�b    P�   "  ��� �     D h��� b  f =����pP@ 6` �pt�    �   t  B� @ Z΀ �'K��}�^O z�L���k���u���ۖ� >��|��Y\Y� �y=/g}��[� ;����C�ϯ���ޓnmJ�<��ާӓ�=������^�y4�� ��

   ��*�a �Ԭ\s��z�m/[�=7� ���2j�n;]�nN�׼^WW }>���W�伴� 6���z���s�� nԸ�)�_{�x�W�y�\��} ���)w����9�f�:�\{Ϋ�8i�
��R�@ 4 ��������J�  �=U*Tc@ d"{J��QT @����R�  �!M�) �5>D�=�����_���M�ggs���{���TUz�������APU?�QTU������qEQV(
���O���W.���L?١���[���w��)�!�?F���0��FH�"��G0�y��B����	F2d� f�%c@�%�#$��Ji"D��dHFP�d���U�	��?�)��P#t!
A"@*0+�E�$�!BD!���""�0�)
�H�>�/jh��ޤ��h"k�)�q`�S�$�R&g�	4с�m3�{Ɲ�z	!��F�`�d�� ,���5�7IFBE�$H�� 0�05!�I����Ѩ�m!'��A�J$���) ��Y�9"q~a�ZB,F�"��
1KȺ�O�dJA��Hb�`ŋ�@��!R4	"0��`F�����	 V���R�Wєc�O۶s	M��)�"Fp�C!�f~�L�P�� ,��C���K�ʒH@�� ��(P�r!
���0�.,(��P�eL%2S4ˋ(J�T�!ICD+�
��Y��� �q�B6�\����8�,kJ`JB�����(�\�2R6N�,�9AJB��2\c �H�#��1!�����@��i�,R�jD�� ����s�����m���+k�.�3y��]��oA��m���g%�s9��7sf���(RIX�?]�{���+գ؉�[	��&�8M�d!�c3���틇�acH��\%q����\%ąLtB�Je��~��S��p-�L���߿sw�N1�$l������ka��2�`@��F8b}���7G���2H��
������*A5yk�*��阸 ! ��*��B�L�.0jd(��#�j°� �$� ��j&	.%�74�u��HI3a$	#�k��d�rnoT�f��J���v�b�$	 ���oȥ�A�A�db膖3$!0ن�Ÿɺ�bŹ��HD؝s	
`ȑ,�V��`�a�Ċ$11�D.h��.j}����X��o��R$�BRBH�!�@�#S2BX�$)�C`AaC$�1�YG�M���6�cH�5%�!`�1�k D#a��5%
��	$Z�O�xF2�s�~�$'v2V*C�(@�����"Q���R! �(@�c�R5X�Ք��5�`�"��D�\�\1�e2-�A4�H�	M¶��%7�ԒNJB$���#�,XH)(�S�$��dԁ� `@cő��F,Ԓ���w$�uS(�%z�z��e��!���b��˛!B�2KD�d,�����d��fn�
���,�-��0	 WN	�8����NoY��C�H�Wf��'
]�֙v����~��?�Fơ�!#
W�5!n��bLR��3[�9%���?bD�dX�M�
a�	S0Ӳ�&����q�{���"?"�6�odw<[v�����oZ_��)�H���7��C�s[�\v?$>M�+�Z��
��HƦa��?hՔ�5�9�B\�!��T��XQ!��I(�1`�FA�I������(�����xYS�HB�@(-(���H0�BB$$)ԧ�� LIB0���@ѢP 04ġ������ �
E�	SU'�$�!T�#�i VH���D�`�4\%a\��dC�g�@���Wph�$�j�$�lKvr515y�g�3CY��`�JILR1 kd4��^� f}�zx�Ku\ ��*J�*�@��) �H~c@� �R6)@��i�G5+���cS	 �pL"d�fd�
MֶI��2�,�
��#$
��!!�j0�@4S'\`ȱ�I$H�dF?HB�@�H�XȰٮ<���8��s���q��>���3A>��0�u���.�&�0�5#@"�2�$�Gd�@��c��JK����%��kQ��X�ԑ�6l�3�+
1!"�(Ku��&I�!M���GXh#d�"=~��忔��xH"����9��X~�o5��fq)"P�#���	�4���0�v�e[�i�
�Ejї4JKto�.}�.f�R4�4�h�����s�.��޿��IHB%�b�4!H>X�� �������XFB�A�@�CXo�;�?s��s����o� a�}?Iޛ!���,)"�) �1`�� R!de�VH��P�4��`8~)>YN7����$ct|�h���W�3?k��Zh�k��!ċI�(BD����b��< XA� �?r�IL�\
��GŀY�P!c%4d�xZ1��BM~1%d�G$؛y+ Ct�!���#��`|R!��	A��A��HE�!$Z�SP�0���D�B��~7��ˣF�F<�#p�!C��	�?�_��9?l8~LF%4���P&�mtЁ�dn	 ��(b���B�~�0�S|5ME�Z�i%�S���\[��sL�&��M��"F��2\csInh!�Hj�9�!�$��1r������{{��v}���\5.	LW!FT�P��n;�L
J��Ey���"f�31"�Nf�)���Ty�]����)��	KX]~�ϥ����q�s�;ĩu�kS��������d�RĔ�Mv��M[B�Fa��I��p �BD HF
c ��i�����Ĺ���sz���¸hD��a�6�s�k�wt��p�0"�".2�tǀE܋Є`@��b���Č� @� � ��$�H�$BB	$,(JF��B��a�X�#CQ�
ܔ�%�VH@�A��!F4�	H�1��!%	BR1���2�R�X05�m$�\u��B�i6*�h6�aq�ۮ����;^��o���n/� ��f���Pῴ�����lKarBa�������R	D��9��;�6���J2�ĩH! �&�~0�!��:!�#X"�RHK3z����D
 p�$�R���R��A^���U��>p����!LB����0'T�_�0���f��~���bF:��P�,�q��\�u�Q�,*I$i	)�K��@��0�G �4m��sZ�!�a��\��.�&�Ӡ˅�+�!
0`�+b����?�߶�z������p�nL�[$#���� �HI"�
�Z� �,aa�������c��!jV�-���ގ����ނkJc*Mk�A�f�bcBD�B�*Jd(���Y�jK���%�����������F���7*�1�)1�a7��y���ѩ	���/�3Wo�Mb3%r�#!FHB24��T�eϘ�#Rc"�4�h%�n�l�1,6�o��y�5�3�Nf$���B�
��H QaHP��b�H�"���B�����%0Б�h�� i�D��# �ЉV�K�~fa3���s�)(B�!��f����%"�JF���ap���6bR�A.�\0`Ĕ�B�� �10ې�
LX��� �"�`h�8���3��O�(�ƆB�HFi6&�ɩ�%3�����3�ɼѳP�I ���n0�0�m��$��	sP�,D�� @�#B"�pHXK�jfNT����IiUȰ�P�WJhd�LFA��TĈHF�sT�݅�������[���'@�9�B�$�
I,�$I����,-���6�p�}����F��F5�FP�J����;1�RD5ňlA�HƑ`B���ݟ�  m� � ~��o� m�m�����  mA��TUP UcSѹ�us�R�+@�4�-M�LO*A=V�URrC1E��g�j������t;�����5�O�'��&�S���UJ�Sʉ�%��Ӗ����*��5V�ћ�ݷm�N�Wl [@)���m�'Y@a� 	v� ̌�����NI&�U@�pF��>�%�Ub���]����\�+U1# m���� -����M����`I$6�5���8X[�[m����n��[b�mf�m��d��'���4\ �M� l�
�U,7��N�j��m�i7I���H��㎐5�6��i�٬�8  |�mRl�40���0�]UJ��KX�u�Y{m $m�bFa�;E@m� *���V�V�J�R �4kp mmm�m���J��I��T��qd�V��9���j�W�	��U�P[[l[I��l5��z�5�ˆ�d��h�PXt��s`ٓ�6j�A��l�O+!6ؙ7J�+���� �^��˶`9��*Z����� msm��[[lM��$�[C��� �5���۶�e�  ��X�Ш��wgJ��� "SH��ҋK��������#� B�wRR2�*�UUV�R� ��ʪ�z=;S5���zI5���V^��$�d���$��r�UR�˳ʠUR��N-L�K� M�e�P $�G�����c�  fCm���N۶�e[��O���倥XM[� �  �õ��V��ϴ�J�J��6�X�;"�yI#m� 	8�۰���W �UZ�jycb,ҭ*pI��n^����!�6�m@m��:�ÁJצ�pl��P j�y�)�Pt�H   HT�YL�m��k����TUĆ�����*]��UR�Rt��1b��` *�L����,�UUPA�:[[lڻ`[��O*��V��A��U��Å��n��6��   հ�C�m��R�UU���k�e6j��YNkH%�]��l-�F�&���^���ۭ�[V 6^�Mn�M����M�UQ�E[@R�5���h$l�Å��.�lm�ie�N�ȐۢI�G����n�m:l]$�m�$�m���'B�-��YeeUGu4 n�Tٶm��ݳ�� Nmm��	 2+�+i6�m�Z�t� [��W���
�S�͖�StSI�[@�lm9۵���   -��d�O��V��jB@t�  mmrޢq �1��VQ����b�  �[�� mIm*���R��`5����C�3]uU@u�2�kntSϗ(ri�������
3�(�h�-�ۥ�`��).;J�����p����� sh�X	�]�a^���s�Yge���q�t�=�C<�im씶�)�.	����*��e�Z��U��U.�-R�c��>[@۶C]d:��j�TԶ�&Î�Z����(i�(�]UU��$r�l�]m��}:}�jjm l ia�� ��mٶ�޲^�a�m6���6�M���Zf�6�[Mjiĳ�[u~7�|m��ӧ\l	v��m� kn�9m�l 
]���h5p�֩���� �l E��-�5��v����Z�bx��PmUAf� #ZZ�J�ն���Kh��l�"i��R�ɕ��jUV��	��W��Ê]� HA����cm�� �n� ڶm[	�^���k�'�W[�R���4.� $.��8 m������W�qK��� *�P!���J��5�R5���H[@-�f�
�પBA����d�	$l�Y5���cm��j�8:I,�YZ󛔈,Zڥ@eZm@rq��]*�R�9c� j�� m&ŽBC����������&eTL-F�`�	 u�`H��m@��ɳ�-mwO2l����ٷm� �Sk�qJ�u���
���5U��c5Uɜ��l�f��X[xݰH��z�m��  l��Н�vm��H���
�K��  �����Z�+ �T�W*��spp�`]6� � m�HD�U���l��uJ�W[[�t�ۦ�f� 	�kXHM�m��ٵFڥz�\� �ETK]9���N&�%%@j   Fc5��k��p6�-�  m��z�c 	 � �0n�:�RUUA�m�   'ޝ8�����IӪL��4�$z����N.�-�v�I���]��������� �4�ΒY��$l6� p @� h�[mk5�Iz���N �� �m���6ٽ%����hmIm�ƽ���8p��t�� 9�l�-��u뵬�۰5J[B�m� �kh [E�-�m�ݰ d�� ű-m�HH@�`f��^�w ܨUU+�0*�UJɀr��6�m��6�6���`m��%�m"K�  H 6�j�m*�K]US�^lm�"%��a�VkY`�0$� ���V�v�V�nN��ɹev��H�qlr6�j�C���z�٘��m�[������Ԃmsm��8再���8�Y�rC�i�m��l�/`I �H�e �hڞ`�W��iW�m�гh6�$m����m�ݶ�M� 5�`m%��n����ٓΗMo-�H�˳�5��m)-�����ڶ4�����`C�4��`  ���B�m�UU�[T��m�F� �m��mmh�tu���m��)Wf��e[b������UHMe4��m<��]��0 2˶�"Am���`�v�m�� ��mS��ݲNm�m�@]x�a"j�RZX-�Vڀ2':�,v�ilٳ��[��$�p�� m���� m��(: 	 ���|�D���k@�� m�m�[V�	 �`�` $� ےC��GY9R�l��N�ֶ�,i�l�@�8 l��@ݰ�`��H��m�F���8�ρ"@�Um@R� *��N�<�%��7 �5��ջ@
�VԬʽ���U��6ĉ -�X��"N9m5�"L  	�ʎ[RUS���l� I~�E���(��݀ZU�Z�d&U�k��m6��. m�o[M�,3Բs�Z � �`�[\m��շ 0n�4�[@�4T���0*�U�hN���b���uA:�)V�@Z4�I&��]���-�<n�v����-҆�L�U/-��Ɗ��si4����}�U�5��[��vêAUʻP �;����Uv�d��6Y.6ۤ$	  �ܚ�D�!m�6��Tr�­U�A�@ts=�o�>[��f¶��|Œ��hn���d�V���WW6��t� k��$�Y%^����c�*�Cf�`�glm�� l 9��l$��   `�R�Z�"��.�N8�m.� J� �
���VV�y۞Wv�Vilն�  ���ڮ��ܫykt�G3ê��b��;I7�6�e�I(n�ó��8ْy��6$6i	�-�Z�,.ۮ^kb�M�H��6�FLE� �$�m�7m7�.�Yy��3�Nj���U@j��%^�{$`���I��K�m�Z� $!�UJ���Se�q���ڥ]�j�Z�U殨78�M��pp-�%�v��\	�l�UTvE���kg��|ij���N������3� �VL�N�N8Z����4�%櫇�m�<�j�Y#�v٢��bt�ښY9��/^���y��Ck�@Un�l*��UUU!5�t6�vM�sm�� l�@�mq��L�]H[@��&  ӥ���쾹N]R��W+Ӳ�Pp+�u�몰���� 6�m�	��� ��m��jD���@���N�]6-���rE��Q��Sm�e�
kw6��k���[u�q� �`M����f�6-��`[tIDڷlZd�k\�^��!����ꕣr�*�a4N Я
�9�k�۩i[�
�y��gM=����:�莼���l m�@vҪ�*�UU�jUm�	��gn���G 8M�m��,�cn��[  >�m��ݛ��U��ڣT� *�t^I9��m rF�M�5��  ����6 I��a���Y��BM��rv�[��.����&���r��~�|�n��+c  9&�����-����8��RKo-�[2���� k� �����`�l��M�h�[B�nH�v$H�i  L���#Z��m�$��Hm�c��m�-�4�-�m� �m��6À�� 	k�� 	n��v�d҅���`!&�-��71q���ڱvn������`�` ��5����lm���d5��  m� [x�aEMa�6�p6�	���ܷ�^u�I�Z���)�6�`�n� �{���wyR�8��*�����4���)�ث�?�A� P�\ZR	A 18&�^ �B�4 ��0���P/��� �b�1#�W� |.�~�1��o���H��N$���ʫ�v��E[�IO�
~=^튚.~O�'���"�@�@�رb~_�>Q��m�� ��8�PE��a�G�� ���?|��:
���`���lb	?D!�0�����1@����TR��m^�a�D >1H�i�����6���TS�&
���Q"�X+H�#�`z�C�LPA��`!���G�b
�8�]�`���T?@O�Ј
 C�- ����� W�)�z`��)�Ch�A�LC *!(�_�`�f��pEqC�p��O�� 6�?���M�D��@m�X5�P"2 �#�H	 %�~�1Ax'Q�$�$�T>D�+�q v~+�a�>Ңh 	"��E�4�Dv� 0��Ӣ0B��"�D��M��QTU��A*$B)��b)�'���ֵ�ffkW"��:V�"B�]��^R����lvq�'G@2�מY�LmtW]Ӳ/3�Sʀ]��.�^��;c�f�)�`B����/<9��G j�Z���*�1��eч*Ava�����;=xɷ�Gu:#���^�mG��D�9/.�C3���m�ݸ��9�r��p �c*vz���&B���+�B�Z�g�%ع�!�����6�2��x�ez؉�y�nu[�ePOA� �!��mJ�=f�K&vҠlS#k�KF���.NZ{;AJ�IQ���d�i�	��b齸fv�f�A�װ�\���ׇ!����α����:=��"$FrA*�a�$1tS6���M��T��Ju��<�]�L!��i+!���9ն!�]�2 5m��U�m�b��)�g�΁��w�B;N�$R��N;`5�Id7<Ǡ���h��1�@�l�C�V8ݐ���&<�ά�K山������vM�Í�����n:����@*l1m
oi���e��4v�q+
#�*1JKTji���R.��sL���m��8�5LXs͝նE&
�:I���+s�z�.xa�َێNې��S	�gn���ط-�d��
@Z����PAg&�,k��=����[:��k��x�[2K����ܮ�V��)r2(���+&�ɱ�Me�%"����R��@e�
{;�!G1��]H�3�f� ݂�;��NB\H�"���6�`�Ճ8�u`�)D0<:����V9�az6�N3��È!���]�v������\��N�і�b�\X��Y�]��l�Kk��V�)sZ���K�]N���+�c�S ���KU�F�b�*ԫ��kO'&�{F�Q]�qӻ<i����R�O����<s=����C�����g,�*�����&�`�Z�d���$�\�>�i4�u.۲�w!m��X=]R�p<�d���dt���
	*\�F�n9i툓<[*Z��=��wz����+����^ ���	��i�M/�S�T�� S�����~ Ҍ	NəL2K�d��f��nۈ۩5�	��p*B�\>\����m�� Ǵ`�!��w)��(�嵜�]�������&f�bSm���K��W�[t�v!�	фy���;q7f�I/\���D���h�� �H��3�<ɮ,�n�#�3����ݞ�Z��z�8:�&���r�pr���ViҲ�3���8��rZS4椹&jL���^�D���}���x}�aU;vs�S�ÞN1�;C�N8˓ʇ�IX�<I�_ǐ9yf��9� �{q����׀#yL�u������:�v �2�+������q*xӇ�B94�]� �`��X��9�)����ˣj������ |� ��n,���\
F�x�6����@�-�@���@9m�|���uA��D��Z�����z�ũ64��;v8�J��{��M@�6/#��"c��rzG{٠7�� �v >]�r:&�n�WY��d�ַ$������b`DN�9J�Q���� �n���x�Ih��oy2)#�[f�_��m�\�zWV���cĤ� ~n�(S#��� �o��J%^��@8a��ouH���M���}�@W`����}���y�3� �jzvt���E�`e��� �7�G3�]v��zFދM}��?�� +����W`h�on���ڭ6�r r� .�:�vW9^�ď���;j$�	�nM ����$�����ڈt`�X@D�R��(P���� ?7x�l�UX%�xLQ94"�4
����٠�f���81�\�H�ɋ#��r r� .�:�\�rW[~�=�@��76����r�y<�81���s�� 	�GjUa��}*u`�۞�*~�r� .�:�\�=̨m
�rxƜI��h�٠q٠^r�h-�@>�b���*�h��I&�6� {���������K�8y#�@����[f�'w�ܝEЈ:��M��w��T�5��k	�9��l��v�+��� ��y�~�����Y��p&w��91)�nx���R,A=�l<�E0���amD�!1���y���W`s* r� �򗕙����6�o7`b� {�P�� �٠s8�m
(�Ɉ�@����m�BS'ou�]�x���NĢL1��#���<J����w�@�-�@����-ajȜ1	8�)$��`Ԯ��T ��`�~����e��Ө�dQ�<й��=sǗP,ov��6[�6ð�*�л���"�[�u[�jX������]����՝ۿǾ��>�FK�)�әrunC	�v���Kh�Gb$]�'�n��>�q^y�gc=h�)@���`�ػ'+�k�x<�� l�:mK^nz)WWCs��P�8����p�h��֡`�����ݜ����u����������u��ǝl�w5�Mv�WN�x9�b��"zv�6��k�)4���n�j졍P]M�߀?.��X������{��8y#���/9w5��P6���u��ۼ��9�YyYto��ͨ���y��+�^]�����bmD�$C��C���׀]�x�x�[w�~��������6�sv u+�y� 9]��w�tB�M��IJZ���J˕՞���m�9s�,;5��\7�M�i�5 ���1��mH&�X�brz���q�x�]�Hwu��R�ɛ��T�wv���c^PDF�BKTj��D+DDG���x�y��5�ŝ(�-Y��Iı�
G����R� ^e@:���5�Ywf:Y����rIB�k�� �}� �m� [�4 8\Cʞ4��#�@���Z� ��J���ʳ��;���f]�|n�q�v��UH�^sͱi�ٶ��s]��ϩ9^N�u�����~.@�`R� ^e@>��*ܼj$�"F�zo,�e�h��hVנ{��by�`�c� ��@��u�'���79@j8��{�W��Y�s���m��R,x��@�PVT 着��~\Ŗ	D�cɒG3@�s@9yf�r�4^]��������91nu��9��y�V��v��9�8� ����4�g7kl�(��$�XƔ�4+���٠r��h��h��X�E�#�&�z���e@9YP���u��Ve7���~����<ʀr���h-�@�܏�co�y�9���`�np[w��,QH�Q
?
�q
"��k���>�/a������j�s7k ��s�t%/�����`m��>�Bx��rLL�8� �D��һW`���ֲ�v
�9�ck�q����k�A�����pi�L#nE��{4�n��n���@����MX&�X�'&��-܀r���[����wf]:��Vhn�m@9YP�r r� �n����\�q,cJI���W`��+* x��.��®�D\�U� kn��(Jw~_�}݋ �m�Q	(��L��ʛ�D�ő�v^
pN"�^�sks�K�]˷] 9�΀h�=�v 
��/��p���Έ䬯n��pnnt햶�v��Rn�h��J���m�MG:l�Nr!���
!9��c!q�::P�-(�BMt��{h$M�� �nlI]<�e��^�t�۝	�4�9�ל��$gF��5p��ezx=���[<�	�3ZneԄ�S�� 7�-��8�.�`�l�n�p���0i��qt�Ӳ��G5G=�'&��m�f��o�w��+*֮@W`v4�Y�YtmV����� �W +�[w4x�tm����y�4Z� 9]�r�����S��Mڻ6�����܀��9YPVf��mz8��V�<Iɠr����Z� 9]�z�+�N��ۅLOb�뮦�g
-p`0[m�%���灰��34��[ҧVŇnm�n�5�� �m� kn�K���X��X���4�XƔ�4+k��fa��*�/U�X
�R��Z��ߝ�>�T�̨��]�n]��YF�fn@�vܲ��e@>Vנs+1�<I���h�P<ʀz���]�}��;�Y�YtmV�y� �̨�k�y� �-��;�ngV�׉&���"B��@�<W汶CK�i��Ԍ�,r�\�Խ:�N�N��q%����I���������9n��˹�{xeb{&$LjxD��@�7� ��,�^,�u�՟�D$��k�&���H��������>�;�s�B^��]1�/댄��!|#�C�I�1�fĪ��mr1���)�)����V �����i���1"I)1�L�kP��"@�#�A�`��C���)HB�#	$�����ѫ)�ü�N9!Eq]��t������~A��}��5����T�_� ��S@�d>.�ċ$"�����V�X1HZ���p��l2�R	IR)-�V�+�D	K,�H�"P$��*aN~�.�5M�!q�a!�D!�$��kRE`�"0b�!%�`�H&��|�h��_��_�| 	�����?&!����k��T �:��!�DH"�\T���(Oj^�`�ذɎ�S��&�U��լP�)|������7����y��+��s@���%ر�8�1�$X��XDD(�}ߗ�>ŀ{u�h��&��V4G��O�nvm���Nƫ��z֞����`̽�f^߾�w{����>z4�"F7#������s@����
!/�y�`H�z�\M)��,��X�x��S&�ذ<����x�_$������ �nUM*�ZVV���,��8tD)�>�Xs�X��(u5Ss2���W3v�9DD)�Ӏy�b�'{��ܚ?��!����Q,B�P�"`������s���1u9H��M�wUW8�/>���y(I%�D}��^�}� �ݛ5=��n��ښy�u��C�<&�� ����P���N^z��j���w��xS�����Suv� ��ŀy�ŀ7M�D%�@��f�s(����0�E&h^\Y�"��]Ӏ>}� m�Y�/�DB�:�/D�I�i��)&h�?ߖ�o��9$��=�ذ�ذ�It��K��M]�B���L�}xwv,^�X
�_t�H�z�H�UUd]�]� �x��/�B��＼�W�OТ#􇻻�R2B�mUUXR�v-k�v.����e�:�î��=V�u�r �k]q�\��&�+P��B[/:���2��LlD[�&�J�(�Z�U9ڻj�;8�tc�d��'w������ET�Ѣ���73p��Vҭ!��v�Y����w]<�/';����pr�\�����!���	[���j��s�Ҧ��6�ӫe{j���j�3!�:��/Q����Y���d-�0ݹRt����w\�Eь�RmT�aױ1y�Vۿ��|�m���v����͍�� �78��.����ذ�N�ZmD�6�2%&h�V�<ď����;��`��g%&�㨪��IJ�໪���݋ m�XQ�IUwwشߟ��@�泘�0N��NL��P������L�wذ���$�����8���3�
6�$rf�y˹�}
/�%�����>��ŀ6�,��o']������\�m��R����Sl[=c��AI�:�ؗ�'�cw�w�ۏ}����VMEL���uwN ޼Xm��D|�Dy������˫�dND� ��@���7PS�0@�����D(�x���Xk�Xt��оJ%
����M"��.�����}� o^,&!B��	%
���� �}� ����e�)4��ѹ<�#}�����{Ӏ7�%�'����6E�'T�M�ʪ��\����� �	(�}�~��s@��s@��[�E�����"�۷u��R`�J��6��*��M#�T��ڇ���w���m�<jxHۋ�;����w4���
K�uwN�&�W)�5�]Mܪ&���;��gВ������]Ӏ7�rJS!���Z���B�.��`ϱ`�s�%�/
!R��`š�:tT�=��nh�����8+&A��'"��
'��� �}� m�X�)�}�4�ꫫI'"FNE���9(�����fN}��ff[����&~�r��~��x��� [�%kG��O �L*�\l�/fx�ⶫs;w���}�i��}���L�|�K��߽�}I%yv�J�j�f}�I��jI.vg|�x�2s=�$�זg�}
��~���~��>��o&fe��/���r�����0�'V� ���z��$�y\Ի�����=�$�ov�K�_+o�CƧ�����%�ƻ/TԒ^��Ü��߻�M�b|������B���7�~�ל��_R{&a37&��cĤSRI[o��%�1���z�K����Ԓ�sRI}C�����bQcH�Qv�۞�rh�m�J��B&c:�rg�qJ�0���1o�(�ىD��#�>�$�ov�J�j�Ԓ�s�ffz�J���=�$��.�@���'$5$�,�{���<��""��'���&fg��/ߦfe��3�fff6�\
�����#'"�Ԓ'�U������~�?/�!B������2fI�/}I%r��p�9$ԗ|�<L����s��=�l����}��[��|�~��5$�{�q��E�<k	��{�I^+ə��Gл���������]������{�I?3<��jB�
�5X� BB9!��q&�0aE�h��I��t?��}y>w8'�����\N �oN&���Ѣ�X��v�H�i'����	wE���f�o6���9�g���%Q�	����l�IY&旳�.,n �zQ1����Z�̚�a�����v��q���v�>B�f�Ohn[J�Yv��9驡���⇧]t��cv���[�7��G�0�V�LˆB�53�ff>���x���5��vs8�39b��ذ��t�;��o�9��)8
�� ?������I%ydԒ\���|��H���Ԓ_\��6ߠ��O	q{�I%yd޶ҽ��=�$��욒K�r�}YC�o�r5"ǂ�MI%{{�{�I%ydԻ�n�^�}I$�{&��_y�Te��I�I3�RK�3��b��I�$��w��ԒJ�ɩ.�������F/-K�)�dĜ�RIr�U�%��잤����=�$���jI/Y�`	*b���"`�����nu�n��VRv:D�
�Ό]yI���~���||o��$�H�	Ⱦ�$��욒K����ԒJ����=m%{/W���Yԣ1���f��ֵ��m��w�9�C����ޅ\Q��TxS�_�n��;&���w��RI+�&���i[�~v5��k��Rf��B�뚒K�r�}]�<��ػz椅{{�o�%�3�U���D��㚒�y�fcw�z��$���7m��������\�}�ݶ��==�~�5<$mž��W�MI���fe�����$.޹�$�g*�Ԓ�¤L%eQ�'�뎛{:װr��nh0�v�\7w��jT�o�w{���Q�{{M�_陙�D$����ޙ�'�U����s� ���m���kv�o̝�g��R���s=�$�y\�߳�̒%�ӿ�����w�K�����獴�e�u��H'&[��n�o}����/~�kv���UQ?�n����{�I�9�$���Q�$�H��{�I
�$���群��+��K�]�����T�1��nI$�jI/���{�I
�$���{�I
���w���q\.%ݻ=ю��6����.�6��)s���Z���8�Q��G���bng����+��K�]�����+��K�r����\C8%[PK�Kn9�$���{�����5$�-��%�v��$��2���<jxL���RH\�sRI}�_s�RK��ORI{˴�Ԓ��*ǉ�ԋ
G5$����=�$�N���o>��9�o���%:���+��?�o_�u�m��I�ŝ��[�0ӑ��Ԓ�;SԒ]��3��z}�Iu>�=I%�9}�}I*�0��[�x����"�����Z���Jѯ �m��u��i]��POŊA8��ORI{˴�Ԓ�ڞ�����群�N��$��Ü
���0�9}I*����g�x�s27-��%����$���O}I."��p�#��I/���{��y�6��z�����z{�I��jI.>y�V4�JfH&�{�K�g����w��I/�w������椒���群���U���D�m��$���O}I.��y�v��RIr�����_'j{m�G�	��8P�������}��BE,V`j$B#%8 PL	$	������a�����ZӥbB(kX����ĉ2-F�G#��4Pهø
��w7��Ԅ�YX�F�����ᆳ��kZ�fd�;e��ў��#v���uXu`;;`!���]麍dv�hT.��XʬU gk�DWin ����;�ɵp�6�Ђ˳&]��.<	Lq*��M#�1�c%-�ګ�d�YF��{;$��2<���<VWJ���"t�U���*X��d��uv�L� ey��\l��l����������~���mK[��J�Ƒ5��h$�n�@�l��P4m/�uV�3O;A +<@nX�������=�6��'0)���t�
���D��g4ǍUJ*Ma+�\��v8,TZ1Ru�C.T��| 'n������ų�:��mP 6n��@�A:�U�jR#+��r�;-�N�%��7�[�Wdd�k�ۑ��̻kj�B��n�f:[t+��+:�VN&w(���U��K�Nﾬ`3 H�řIGe��F���3��Z���WE����&P��9P���bZ=xQ��)�c��3[z�!�aj�/:^C�'O\]r�*Q��c],dڔ����� ��'�q�6�f&�k�hEq�u�e�eY��C��-���Fڥ�xcSY@R�-�8w2���[r��'Se',�)���ö�v).S�	�6֧u�b:K]m�y�up6y�����
'�9e�����Q���ȵ����@Jr���Lŝ��&�
�S]����gP�j6��)gOC]B��Y�
X	ݛK�R"I�l*�q��S��5nks�On��%��Y�E��V��)�||���8�YT�m�c׷&��ݜ@��{<�9ۧY9-�л��������H!�v��=��^����țRcb�#�)�gtc�Wm�����WF�Ī��ۦ�c��P�d�uUٯVӗ�6�c�3�|>K��-`2f��n��-R�Rqv%��Rl8�Nf56��݅8�����X��P+Ƶ����'
��<�[t�E���2�� ΍�uS��W$�T�V���3A�\c�@���b"����	��P>Q�|�T�h��%�h��]gn�6L7���m�K�R[lv�m��i�N�;�=�TZ�ZF4�J�����ݴ�#oQ�����6����Hu���n��fv���;�����cs]s��3Qp�ͳ+���Om��㋥�M�.�<Qtvg�y���a����N��s\+%	�fy���u����0�n��SY���]/LGM�p��S��W�T��Z��R����}�o����)����@�pvֆ�k.�H\\�,uݸ�?���G�+��˅m�r^�KkRH\�\Ԓ_s���Ԓ�;S�g����ޞ��]E[Ky��c�H椒�����Ȅ�_]ܹ���ə���>?~��'u��q��Y�{��ĢOy�g����SԒ^��=�w�m�޹�$�o}�}I$��_��pdm8މw<��v�{��sRIr������y�>I޽ ᅠ��5$�br-���@�fy�e���.��@�|�@�^q!�*hY鍻v:�:�=rn��c����+���e���j�$�癙�3R�cĵ6��$r?@��ŀ~��`�\��>J!z�����>���SJ�L�Wd�Z�?Kn��8D$�Z2H
T�R
�-
�� ;C�*g&���ܓ��}���������εLZPK�K��z�}8��:L�}� ;{� ��M�����O	qhw1.r�h�����^�q^�ՠ^Ջ�~&�r5"�M���^,��{��������7���U��{Bi�%.]�����k�M�ڃ�U�Й�34�A�ݾݷ׏�HPUe]ݯ����5ֹ�{]��w�nh;Կ?)�ܚ���9 �P�������qB�k�jH#"��Z�^���sK�B��T.�W����;k�p73t)S.j��.����IB����� 5����\�yt*�}VO@�D��3V�d�m@�٠?��o����2���1��~n;>�=���{`��f����v����ֆ7�]A��R[�7n���}񏐰s�M9=�ޭ ��Y�r��w=@}��h^�����Y1��#n- ��Y�ċ��� ����9_*ޤ^Ջ�~&�#R,b�M��s@=�٧|�+�z��}x��\S�&�i
���Z���U��������{]�TB����@�*VER�����s�� �~?%���!$�LQǠr�U�r���u����X�����UT����9i'N���]�lV�w�j���j'�erk&e���w�{���7G½�R�n������5�ŀ���J!G���tt�1b�M8xF��@�������IB����׀w��N {��9DB��p7�I���j�`���u�p��$s��@����=眉*�X�"X�j�����pu������S>��h^�������O	qh�r��J|�����]k�DE�&!��`Ad��P���� B~?O��3��3U���!R
�fV7�Tq���q�]����:���0���v�FW�[���0[n��u)���-Ţ�n�4��]�� �" �;sAc�c3��j䃰��]����F�m�z�`ݝ �Tm�	���&�l�c���Ŏ��-��q�x#u��Z�\�=�;jKc�96�6���l�T�-#�c�1ڧAWU٧��(��P��]�*���wp��s���'�.��j���ݹF��3=���^�)����r��4V7ˇ�z�1I'�{��� ��f���Vh�r� �×�[m�<��s4߭�s� ���@<���S�n~�����K�sv��@>�s�+* }�Y����(ڒȰN�����7��`�k���8�7�&���jj�.j�� �o��I/�k��w~����+��>�F*%@�d���sr�չf���M�d��q�)]j���T%�]�����L��0"M���^�����ܳ�z���w4��$�5��D�4���lɔ$�B@�"�yЫ�����X���}	%���S򚪀��O$�C@-��}m�ӹ���;٠[��@�����o7#R,�7$��lD �.~��, ��׀n�fB��}���>�(�y�f�{��@�u ���<��_�r��2�K�2��ˀ�A�{g��8��0g'<��2�nx��A�R���1�$G'�[��@=�w�y���~�=�׀\���U��B,&��{]��(��}� 5����ٝ	L��j�]4�j�.��� ��ŀ���DID"!
�aP�Ab�d@�!�ݗ� y�^ z��2SH.f��(�Jg��x}|`���9%��}���.��!�#X�rh��:J'u��{� ~�w�kU�T�}j:5�5nǻmm=�bɼH�m���)�]#�T����;�*��K�5��o��w�y�� ?y���H7�� �����܍H�Dܓ@�۹��<�ă�w^ �_�k��">P�U$9�Q�ȣl1��&h/��@�,����9�٠s���z�%^ �M�	ɡ�B��8��׀y�� �"`�D���[�����uu$���$��}�4�x����u�0�K��$OM@{�����������f�99��V�b�g��n+f�q����E1�D�'�r|����~�w�n�g(�����6D6"P�s$�� ��f�<ċ{:h9{4����<ď�X�.�@cjF�4���� =�w�B�3�݋ =�׀~�2�����F��C�g��9{4��s@=�٠}_*�9x��<��ԹWsUwx��X%	O����O� =�w�DBJ,�i1�;��*e�T�/Y�/@g��G��	���:[ ;6$��@W���@=�7m۸�6A�V ��9�v��=�h����=q;4��6��� �pj�<�=�2x*���{S���9�[Vw��B�t�;U���V]�����G���|s�e��kb��V�u�h���9&rF��9z,�cM�p:+"
���v)(�k�ZX�Z��m7;F��u��fڻ�������;g�|�8d�]�۝�CЃ��g�u�q�k���3@7B��#'�L��"��������:�8�k��Q�A�v, �&�z������%U��Z�:"&Cu��"!B�!��`���BS&�\�R�.�5w8����x���=�׀s��hR�cS��xF��C��+��� =�׀yֹ��#�UM�׀t��|�2W���ـ���	o[���^��YM�R�c����<�d|�q�l��9y�m��姥�ŗ���B�!�F�6�kNO@�]������>�� {{� �tuUX*Uj�����{]�@�c����$��~���� ?� �s��G�W*�D�nF�Y"nI�^vt�~�i�1.uޭ �/f��<��2�ĢO#��~�w�yֹ�{]�|���� ��]x�4���ɠ}_*�:������4߭��8�1y"ǃDɁ�����Z���yj��"���ם��I���~��cV���8��NE�9{4}e4߭����Z:tQ��xю�f���@�� �� ����W����f���	�8a�4���}_ݻ�0��!��T�@EO�b�+H2pN)��v�� � l�JÇ��E;�HTM�6�`��	�H�ϔ6 7�!�-+E��>@��O�/�H���ѽ�<U�n�����}Ω�*�iБ1�BI��imB��m���M ��b8� ~ ���D�~O���� �:P�W�8 Q�b���hT∦"�ځ@���\��ܓ���@���T�6�kNM�v?� ;��w�H��`u#�fd����qh�r���ޞ�}��hWʴ��&�+!4��@x��w`��ZLC����]���=����A�����o��rO�r5"�rOC�.�������ε�(_/P�׀9#��>V�nf�Zf�i >���sp��`�Rx�g�Z�_�#�܈HnM�w�@>����(�����`�����L�T���"r-��x�9{4�Κ���[������]}۹';;R�ʞ4c��i�4}e4��g���{=�w�@>��h\�����f&�um.��z�]�s��N��͑��x�{+@�y���aB�0Eũ©L��\�]��=�׀yֹ�{]�I~�{����`ꚫ7"Pi94��Z�ܳ@��S@=�ٽ�3>�|�i���x�24�Z����a�
&Oou���8z&��3K��ʫ�����#�IWw߾0���}]�@>��h��q��1(������l�;�s��^�s��@�� ȅ
����ҧ��ڠ�,*�]�.0�F�e�"j@n[�{������ۜ�]m���n�.~v.V���huv�Ԑ�N�r�\�Yڨ��lx�[V$�uB@�6�n��nyK����l��wg���:"7K���v�1{m�K���Z�k�;u�+���8M�tc��H���`�=.,�^�m��->�^U���3t)J�^W`�鬎�0��v<^9�k3� J*���I�V7Y0�f�m��؈񍜑h�U��U�#v������8�?�wܼؖ�A�	��;���- ��Y�s�S@=�٠|���M⩥#Fj�p��y�27�� {{� ��9bG:D�xَ���-���l���:�ՠ���8�/��F�)</7H��`�[��; �u �xVۀ��J'&��v���/g�r�t�~�h\�)K����(�77mho�Ms��:��s��|�A��DcM4�#9��9@귯@��@˰�H=t�^QyR�ouL�s5��w��x`&@ iG�"}_��u������?H�:$q
4�p�8h�٠^YM*�+�>�S@2��
�dL�	ɡ�_:�}�@=�ƀw�� lv��{�e��@�r�Ԁ�hr�h���2�reX�`u��4�m�}jSrb�&�.;Ü�]��RS-\�sV��"c�<$�G���4�l�>����z�#��ѼJO$�����@�r�u'��?�X��I�1�x�rh��4
�˛���	#60���"х ��U�1|s��k�`��@��UC[�X��d���gu��� ���r��8��r�x'��)9����e4�y��;�������!D-!%��(�I�n?��m;OT-���U��sc��<�펭�j&��t&r�e �u��ŗ��wV`�w�{]� s����"=@��~4?yދ��DƜHHnM�YL�J"d�o� �����ou�@�ƞtiHЅ�U�W�w3��{�?BIL�?����00rZ�:SB� ����J"w�8����7]� \£{����','_�٘[��Uv`�w�tDC}�~�����4�*����Y`��2D��e�i�-��]��ĭ:5w^����J��{���w�u���nE4���ogM���e?y��;��hΝ]M-c�1�$r��9�/�P�P������^�v��}��9}��H�X���UZ������� .�=Τ���Y^,M��&jfk57%?�� ֿ����������BI|�T������E��"cnHnM���\�x��`�w�l(�HVD$(%-���￦?}�B�e��@�<��+0m8��\�l�A6��Z�Q���2\i�d�X�u��s�[r�6�ᇪ�Wi�.ޛ�26�mكpB�X^uۧu�	���`)�uc������ű�m�01�6��ny�5j�Z��[ �YZM��E�t��n��޹���!��]:���a�8�[n��z�L�"4��L�kM؁{KO�q�S��z�+u���{��{����}*��ЗNL�q��gu����N�ܼj'�es�&I��]�wgm��G��Q�"p��;��r�h�٠}�)�|��'�*`Ӈ�����e4����@�r {�ߺ����ݪ4�� ���Ԁ7����h���n`�D��\�ޚU�zܲ�Ļ��h:gz�jf�[��@�r�u ��u��=Yp�*G�2s �$bMݶk:^�`�Yvc`�[3�T�=SA����{/\��c���@��M �[4r�w3<�����b�6D΢O�&nf�VU]Y�$���[��"� �D�P���� �� ��@
k��r��˼��ԕWx�`u���3��� v�M�08�Ӧ1H��ӆ�s<�<�7ߖ��� ?7x�%��0�����Ӈ����ܲ�|�w���}|`u��<�(JQ�D�����t�Q�ѥ�x:����Y��I��I�A0��K�"b�O�ő�i��	�h�٠}˩ {�Ps� z��B�̣3hk"NM�YM����{��r�t�>W��|ă��i�!�Lq�h���䟾�7*�D���u ����`�ـn�:&�T�M�ܪ�Sv�9$���S�|`~� ��fϭ��|��`%x894��X$��q��ذ�l�=/]Rv^�ҏ<ӆ���G���=&pl�x6B��d�8��|-���[���"���*�����o��$�!G��}Zk�4�xI�p�9����?yGw��9�����3�Jd=���iU.�����j�`��z^�á(IG�
����`�� z�:�SVE̕v`tBS�ϫ ��� �7�RIbEʴD"�
`�PBNIBJ�k�iܡ�ܔ��EJ����<ݳ �$���(���^���h+��q���q/"YA"j蹽�K<sjm��D�lm��N���<�M�֜y�\г+6������YPs� ����z������՝bx7��)9�H�k�gB��g�V���|�,�BH����Or8h]�z�v�>�S/{�`���l˨����2��/w �R�YP�R�����z��m������N>�������0DT^Bȴň�����9�D�",Ix�T�0!q�$�k0�`'���A! (��"|��'��	|@��M�	�4I�x��%�^�t	�k�~H�8ȉ��,$������� ���%��X���p�<(���G @f~PHA�`b�Pn���@�L!S(s��@�i!�A�������>��խ]h]��� �"5<y�UuTs@-Uܫ>]����]V�1ѶB�h�1�
�mcX)�*���u˝Z�a)�c��&��G"L��ۺ���w:�����4Npc���k�wm[)���K,��pE-v]Gj�g=�;��0T
�kkzB�C���級M�Ǵ\ҨR<\I��y�ь�A�'J����=*:���gsF�m�ִtB%����g�f��@5mp�����g�el覚J:�
�Ҋ�Ķ��k�1s͓����u�,��w))���RKp�UN�PeѻV@��T����e��u�-X�g�!�l��"	��x���zg�q��ue:!Qmʝ�5cmTN��=��!r�5��zJ)��d\G 6p�35,�rJ�NA5�&Ήh5�n�nM��6ig`�۲ͧ�� jat\A�se�b�n�-�*��07iz�ۚ\�6EY�`F�lZ�x��Q�uˍ��AL ��e���b�a؍�)�r�)&��Ҿ��l�#(t��\m��k���\0l3��Ue6w$@�] �X��������%�VM���0�-�Tc7X�.���ˢ7 �8����J0a�o5+-���T�\����j�6��U[F�;u�(OR�͑��g�#�r[vL���R�6�g�Ueb�T���m�xwml"K ��!��ق��^�V�Ơ�[�탈+�T�6X3��F�7U]����{(؀:�3�<od�R���.�,�e-'[K�M�k�]d��0�m�ѱ6�	vlCc�>�8+�sԼ�m�9`�˭����k;>��0;�;�^0���㎝8��HP=v��<dX
�TCKTcܲѵ��GNp 6��@$���ӓ�h�,�<�b�j��Nب�g3�%���c-*/-�lu�mԵO79n���;m	�,=���Ce�ܹ��.��˄��]�۝(m<�d�,��Y�Y��m���X������z]�qR �F�3WSq�� lz
uU`h�ؐPC�~��� Fi�?�A> >P�+�����co����^��n�{P�Z���h81�17a�4pV���1H�p1׫9济{q��xƼV�[Il��m�x��'7G!@$�O&����ss2���](�'Q-�^,
����f[
ssq�n5Mt��͔�Z���@�'&�֨�^��UΣ;�r�7�i��.�勀�UX����x���
��bݖV�#�Xs;�{�������w|���m�sPO5��wH��O �Q�Ee��,>�zY:�[U�;~�����<𹷴����:h+���l�g�/;�� �i�η�8y���@��f�o���(����\�����n`�8�z��~4}n��YM�y^�����ۀ��c&8�4;�+�ߖ �_��P�{���Q4���nn�U����n�f�%
#k�W�7���7���=�@TR�"T�<��N{'nzƔ��;=mͭg��=�"5J�y�37�$��<2H��]�z��`��}	/�����z���USwX��e��ԥ�}�����h�gM�y^�x�\m�U��t*��0�x��lâ&vy�`�}4��<I�YSc��dnf��YMӺ� �v�IO�w��$��-�g��3Qճ5���Kı>Ͻ��r%�bX����6��bX�'�w�6��bX�'{��m9ı,N��rIt�ݳd7�k#��:��7@��-�����ŗ�����ŭш�e�'1O��D�,K�{~�ND�,K��ND�,K���6�"X�%��>��j�B�����X�]U�$�V��WWf'"X�%�����"X�%���~�ND�,K�}�fӑ,K���ߦӑKı?t��K���WZ�k&�Fӑ,K��}�M�"X�%��>��iȖ<�C�CG"r&���m9ı,O{���Kı??Mt�ڒ�[��CZ�jm9ı�}�fӑ,K���ߦӑ,K�����ӑ,K�FdOs�m9ı,Jy���Mk-̳4eֵ�ND�,K���6��bX�'�w�6��bX�'}��m9ı,O����ND�,K����vۿP�Oc5�v�z^2t��8��x�]é�vΈgr�H!mvclOϳI��56��bX�'�w�6��bX�'}��m9ı,O����ND�,K���6��bX�'�'ol���33Q�5sFӑ,K�ｿM�!� 1ș��;���ND�,K�����ND�,K��ND�,K�!<���fL�u35���Kı?g��m9ı,N����r%�� �2&D�}��iȖ%�b{���iȖ%�bw����M�H��T�������$)>HJ�]�߾6��bX�'{��ND�,K����iȖ%��?�? a�_@-C��d��X�ډ�s���r%�bX��Y�+��D�������_�RB���{�ND�,K���ٴ�Kı?g��m9ı,O���m9ı,O�?~�?n��kثF|8�d��uf�&!�L76y�v�)�k��@[�����Qβk4m9ı,O���fӑ,K���{ٴ�Kı?{���r%�`L������Kı>��O�In��f���5�ND�,K�}�fӐ�Ac�2%������ӑ,���;�p�r%�bX�����iȖ%�bS�ݷ�I��ne�u�fӑ,K���o�iȖ%�b}�}�iȖ%�b~�w=v��bX�'���ͧ"X�%����ل���˭[�56��bY�
�ȝ￿ND�,K�{s��9ı,O����ND�,K�{�M�"X�%��N�ܘ[g������6��bX�'�v��iȖ%�a�1�]��ͧ�%�b}�o�m9ı,O��m9ı,H/�璘2�%�Z��%ջm����爐�+��񸤩zs��S��M��&v��Ҕ�Ay�	n�\71���\#�xx-�h�5f�'���.:
�kZ��v9�=���N:���4T��/	�hz�B,k�p].v�,�2D���2�+��\��B�g,��n�pl=�t(I��үV9�;B�%�C+K(lκgh1�:���W�����l�]�{/\O=�[cz7�F�/�k�o�GE��i햡d��u�M��sQՖ�S�Ȗ%�b~���ӑ,K�����iȖ%�b}�}�iȖ%�b}�n�6��bX�'~��=e՘L�)�3[ND�,K�w~�ND�,K��ND�,K�w��Kı?}�siȟ�eL�bw<��։f�&��kSiȖ%�bw����Kı>��~�ND��ű?}�i7���6��H���L�%�fe�34��H���ݻ��r%�bX�������S"X�'����ӑ,K��}��iȖ%�b~��'�-�˄�C.�jm9ı,O�{��r%�bX����m9ı,O��m9ı,O��ߦӑ,KĽ��H�ԅ��[�&���Z}�u#��Kn�K=v��j��9�.ސ��Y��sE��m9ı,N���m9ı,O���6��bX�'�Oo�iȖ%�b}���ND�,K�$�a.e��u�a5sSiȖ%�b~���:·0V��D�K;�M�"X�%��w�ͧ"X�%�߻�M�"��{���w���o���o��̖%�bw���ٴ�Kı>��ٴ�Kı>����r%�bX����m9ı,O��I�)=��5�W5�ND�,�`dN���ͧ"X�%����iȖ%�b~���Kı>�W�ͧ"X�%���n���&f���]k6��bX�'�w~�ND�,K
#���6��bX�'�j�ٴ�Kı6���_�RB����������r*��=���r&�F��:�ø�d��*�wn9���|�νH���nu��������bX���7�M�"X�%��ھ�m9ı,O���m9ı,O���6��bX�'��L�\�.��Lѫ��ND�,K�}��r%�bX�g{��r%�bX�}��l?�'�ı>����ӑ,K��;��'���Yp��e�Zͧ"X�%��w�ͧ"X�%���ߦӑ,zhT�@��9��� �>��Ow�M�"X�%��u��ND�,K�{�}��Y���F����r%�bX�}��m9ı,O���6��bX�'{��]�"X�%��w�ͧ"X�%��ڒ{0�2�d�հ�����Kı?w���r%�bX�w��]�"X�%��w�ͧ"X�%���ߦӑ,K����ٓ.L��NN6:䃸1]�u�:9�]��yͮ2��G-}����z�%��������ow���y��Kı>��ٴ�Kı?{���r%�bX����m9ı,O���딷�s5�u��ND�,K��}�NC���,O���m9ı,O���6��bX�'����iȖ%�bw�.��.��fje3WZͧ"X�%���ߦӑ,K���o�iȖ%�b}�w��ND�,K��}�ND�,K�>��\�a,�4dѭf�6��bX�'��~�ND�,Kﻼ��r%�bX�g{��r%�`i�$d@���w���m9ı,O���f2p���3F�jm9ı,O����iȖ%�a�1����~�bX�'����ӑ,K���o�iȖ%�bw;	m��~�b���Bqs��cO+�����L��ԘA�� �kw5ά�f܊��9ı,O���m9ı,O���6��bX�'��~�ND�,Kﻼ��r%�bX���_f�f3&�]kY��Kı?w���r%�bX����m9ı,O���ӑ,K��;�fӑ,Kľ$�p�����V�����Kı?w���r%�bX�w��]�"X�%��w�ͧ"X�%���ߦӑ,K��'{s2��\��������r%�g�2'}�g��r%�bX��{�6��bX�'�w~�ND�,�"� ]D��߿�ӑ,K���Y�)o�\�G.]f�ӑ,K��;�fӑ,K�����iȖ%�b~���Kı>�w��ND�,Kh�ȉ�����%�L���a��P���ޟE�M�g4��8�=��絮��w<�����EFm�9��	(keF]��r\�.�3�&��Σ�y�/9)�x�k���u��K8�r��ڴe��Sn�rH �c��]��;��&Нl�8)�p1���L�J�x��Ѫ͹�m)iL��:��8{I����Al9\X�����1P����ۮ���Osԗ�1�ы`�	�&5"Aís]8�l:����]�vz�;=�OL�9ִ�34L�j�Y�v%�bX��w��Kı?w���r%�bX�w�~�ND�,K��}�ND�,K�>����K0��k5���Kı?{���r���,N���iȖ%�b{=���r%�bX����m9ı,O�}완��.��L��kWiȖ%�b}�n�6��bX�'���m9ı,O���6��bX�'��z�9ı,O��x���L�桗.jm9ı,Og���r%�bX����m9ı,O{^��r%�bX�}ۿM�"X�%�>��x%ƛ 5${�zy���#����Ȗ%�b{���ӑ,K�����m9ı,Og���r%�bX��ۼ|��ؤ�`+��1�I�j���cN��!Ո��xv!3/E/���mO ��ln܍6��bX�'��z�9ı,O��ߦӑ,K��{�ͧ"X�%���ߦӑ,KĿ};�.e��0�&����r%�bX�w�~�NC�,�	'_���~��K�{�siȖ%�b{���iȖ%�b{���ӑ,K���Vu�[칚�\�Z�ND�,K��{6��bX�'�w~�ND�,K�׽v��bX�'��ߦӑ,K��ަ�u�	��e3WZͧ"X�%���ߦӑ,K����]�"X�%��{w��Kı=���iȖ%�b_���_]If�5a�f�6��bX�'��z�9ı,?��޼��O�,K�������r%�bX����m9�7�������w���dn)И]�ۂ�v��ˢ���D��%�ۇ������cp�{�77r�˫���xTB���t��B�ı,O����ͧ"X�%���ߦ��'�ı?����v��bX�'��?�-����C3.jm9ı,Og���r%�bX����m9ı,O{^���L�bX�����ӑ,K��η��S-�a��tL�ֳiȖ%�b~�w��Kı=�{�iȖ4]�� �`�}!�>��!#r��FHB�	"$ �b�$���`F����KO�İ��ڏ� ��dя�o����T14�M�<^p�$cH�I+'h`��&l0��U���
	�(���6��#�$M�@�I	�B1F0I"4JC��&� 8�XA$a6B� G�B�aE �HF$�QM�-��H&�O�iT�� Q@�C��G�U��@���R'��șϮ��ND�,K��}�ND�,K����˙�\�Ke�M�"X�����?�ӑ,K��}w�6��bX�'s��m9ı,O���6��bX�%��ze�0�k.�ֲ�SiȖ%�b}���m9ı,N�{��r%�bX����m9ı,O���6��bX�%?|I-�����uf�.�t�9��x�9��I��I��)$�e�����<>iu�35�n�6��bX�'s��m9ı,O���6��bX�'��z�9ı,O�ۿM�"X�%��M��.��fh�L�ֳiȖ%�b~�w��?��DȖ'�����ND�,K�����r%�bX���ٴ�Kı/���/���ѩ�֦ӑ,K���o�iȖ%�b}���m9ı,N�{��r%�bX����m9ı,N�x��̜.��L�5��ND�,K����iȖ%�bw;�fӑ,K�����iȖ%���`  Gʴ*�5T!��~U�4<��{��ND�,K���d���Yp��fe�M�"X�%���}�ND�,K���M�"X�%���ߦӑ,K������r%�bX����ne�.�d��B1�1Ǟ'�O��gc�ד8�б�6�V���"9	yT�:��w�{��7����ߦӑ,K���o�iȖ%�b}���m9ı,N�{��r%�bX��{	�=�Y��˚�ND�,K���M�"X�%��{w��Kı;��iȖ%�b~�w��O���,K���-�a���5]fkSiȖ%�bw޻��ND�,K���6��bX�'�w~�ND�,K���M��G�L�bX��v_9K��fj:�n�6��bX�%�����Kı?{���r%�bX�}��m9İ?������B�B�����}+�LڤUZ*U���ӑ,K�����iȖ%�b}����Kı>��~�ND�,K�����"X�%���	��6Lp��8�~��WL��E��vѷw[�7t��p�4���rT^�9r�k�i�θA�
ݓ&��&yn���Q�Νr�Ӷ%�vw�Fi�-�8n^*w/A����nˠ���۬���d���u�]m�硝�<��51[�0�v[�8#F�[\�rd���G�kg�v{Jz��֨���M�x�Ѳ����7K��ٚDQK N�=rpw�{��{�w��o��<zl㶄ы���u�M����`;��.�v%Y/��:{E��,��;lO��v%�bX�{���r%�bX�}ۿM�"X�%�~���ӑ,K�����iȖ%�b{���32p���3D�jm9ı,O��ߦӑ,KĿ}�kiȖ%�b~�w��Kı>����r%�bX����,�.��3S.\��r%�bX���m9ı,O���6��c��� w����O�,K��w�6��bX�'s���2�ff\�D5��m9ĳ�`dOw����Kı;���M�"X�%���]�m9ı,K������bX�%���e�h��԰���6��bX�'�{~�ND�,K���^M��%�b^���[ND�,K���ND�,K���ݻc~���E���&Y�䍴�h�:(���Xz؞��X��nK�P\�s�/X��f�6��bX�'����iȖ%�b_�����Kı?{���g�ı;���M�"X�%��G�ͥ��35\�Z�ND�,K�����!� =� u ӷq9���~��Kı;�o�iȖ%�b~�n�6��bX�'}=7'�n�&f����ֶ��bX�'�{�6��bX�'�{~�ND�,K�{w��Kı/�{��r%�bX��>��h�34jC2捧"X�$���s�m9ı,O����Kı/�{��r%�bX���p�r%�bX�;;�3�p���3D�jm9ı,Oݚ��ӑ,K��c�������X�%���p�r%�bX�}��m9ı,O��I0�K���,���"yѓ�x:sƹ�cF{X*Dj�+v�[��tbG�e�{���ou�b_�����Kı;�{�ӑ,K���o�iȖ%�b{�^��r%�bX��7���u��r]I5��m9ı,N����Kı>����r%�bX��׽v��bX�%��{[ND�,K�C�������jXI5�ND�,K���]�"X�%���w�iȖ;D�"A�@�1D�@R �P_���K�w��r%�bX���p�r%�bX����ar��\�SR˙���Kı=ٮ��9ı,K����r%�bX�����Kı?{^��r%�bX���܅��������j�9ı,K����r%�bX$}������Kı>�׿�ӑ,K��f���Kı>���-�f\ k��-��C��&'��4e�i���
�r�M/+Q�v��gkc\�[�u������X�%���p�r%�bX�����9ı,Ovk��ND�,K���[ND�,K������2k5�	��6��bX�'�k��ND�,Kݚ�ӑ,KĽ���ӑ,K�����"X�%������.rK��S55����Kı=ٮ��9ı,K߻�m9ı,N��p�r%�bX�����9ı,Oϧ�,�.��3P̗5v��bX�%������bX�'~��m9ı,O��}v��bXZ��)."��(`b�� P?r&d����Kı?������n�3.K��ֶ��bX�'~����Kı?{]��r%�bX���}v��bX�%������bX�'����ff9m�dݴ�s��x���8�k�J��箹���L�ݺۮ�j�YUd����)!I
H\�ύ�"X�%���w�iȖ%�b_��kiȖ%�bw�{�ND�,K���3���jjR\��r%�bX����6��bX�%������bX�'~����Kı?{]��r$� �H_$� ���*h��X(@����H�~�t��H��?{]��r%�bX�c�2����$.gd�I%�EU�)���m9ı,N��siȖ%�bw�o�iȖ%�b{����r%�bX��w��r%�bX��><{.�MMf�!33[ND�,K�{~�ND�,Kݝߦӑ,KĿ{��ӑ,K����6��bX�&�H&��#�F(0�@'ݳ��}u3VY�S��Z Es$ÇDc�N�Ռ�M%��u׷éWg������x�}���CL�`���v1�\7p�܇R.����i6�/Up��Ƅ���d��v:���mk��\�]�V3�H�-$��T'k�uʶ�B��R�`غ�"㰺N�_BSx�Gkk$D�#j�9R�v�b)��]�d�:E\�#4�%�9�rM ׿���{���v_�]�G�S��qk�ի�k*sՋ��y�v���U�ׄ��N�E�5$9�S�G��1g�'z���bX�%������bX�'~��m9ı,N���m9ı,Oϧ�,�.��3P̗5v��bX�%������bX�'~��m9ı,N���m9ı,Ovk��ND� ʙG��Q�?,��ؠ�7����!,Ow���ӑ,K���ߦӑ,K����6��bX�%������bX�'��ff\��SY�c5�ND�,� dOw���iȖ%�bw�^���r%�bX��w��r%�bX����m9ı,K����L�_\���%�M�"X�%����fm9ı,K���m9ı,O�{�6��bX�'~��6��bX�'����m̤�s���L�4>�u�z7M�m�ø6�+��e|t��P�yn��a���\���3Y��'�%�b^�{�[ND�,K����"X�%�߽�M�"X�%���߭�r%�bX��wvOYf�&f����ֶ��bX�'��NCJ��Ԉ��Ȝ�bo�o�iȖ%�b}�w��9ı,K���m9ı,O�>:{5�K��֤&fh�r%�bX�����r%�bX�g��ͧ"X�$2&D�������bX�'�����Kı=�w�fs�]]j���֦ӑ,K��>��m9ı,K���m9ı,O�{�6��bXD�=�o�iȖ%�b_ǥ�g�Yu�	�Iff�m9ı,K���m9ı,O�{�6��bX�'~��6��bX�'��}���Kħ����*�,1���1��I��/m�*F8�H2��l�E��շ/H0��`�m�![��I��k��%�bX�w���ӑ,K���ߦӑ,K����6�L�bX�����ӑ,KĽ����˘SSY�aeֵ��Kı;����Kı>���ͧ"X�%�~�}��"X�%�}�kiȖ%�b^��˅��j�����Kı>���ͧ"X�%�~�}��"X���ʞ�0U���(D��'�?�����bX�'��o�m9ı,O}���)o�fj:��k3iȖ%��2&w����r%�bX���kiȖ%�bw�o�iȖ%�b{�ﵛND�,K�N���,ф��2����ӑ,KĿ�����Kİ�c��s�m?D�,K�����iȖ%�HS�������$.i������݌An��wci��u׬;�!����k]ۗ�ѦI�����TbN�g}��Ou��=�'~��6��bX�'���Y��Kı/�ﵴ�Kı?}�p�r%�bX��;�˅��WZ�k.����Kı=�w�ͧ!�R�"X�����ӑ,K�����6��bX�'~��6�����aQ
HS��~R}`M�H�EUU�m9ı,K��kiȖ%�b~����Kı;����Kı=�w�ͧ"X�%�����2�332]�f���Kı?}�p�r%�bX�����r%�bX���fӑ,Kf��D���w�kiȖ%�b^��ٙsWZ�K�Ѵ�Kı;����Kı=�w�ͧ"X�%�~�}��"X�%���{�ӑ,K��-��m���f^��[nlpb�<k<�K�n�k�P���z)y���`xxG�N�Go��̖%�b{�ﵛND�,K���[ND�,K����"X�%�߽�M�"X�%��^�e=�e�GW5��m9ı,����ki�%�bX�w���ӑ,K���ߦӑ,K��u�k6��bX�'~�ܞ�٣	��e535��"X�%���{�ӑ,K���ߦӑ,�@�Dȟ�׿��ND�,K�����r%�bX�d}�=�֥��kR34m9ı,N���m9ı,Ow]��iȖ%�b_��kiȖ%����"}����ӑ,K������r��Ir�T�eֵ6��bX��$������~�bX�%������Kı?}�p�r%�bX�����r%�bX�S��R$�Oߍ��O�"�bFX�c�$Xq������]��.�$ S�Hq��T���@`�!<C�G��,�D,V�
��J$�A�"}��k��Æ��� !7�:�;�� گ�6���B� ũ,$ЈA�_�۶h����T��a�T8l�>٤~�ŐH�"D���2"@��$�dc@��?�H4�Ǧ�ҿ�b�*B$RB	 F2F ����"@^�B��9��H Ȱ갰���|}���㯹���~4E�1a0`A�X`� X��Ц,$`@�A�E��ą��2X�g_��v��IU]W;�r�yY�x��vh��86W8�8����DѨ-.fa�C��d����qkx9[��#�*�����$	�j�H-Z7mq�6���ZI���\�Ŝh���D�=��ss��e�{e]��L9wX;��-���16ZT-w0s��6vz��X--�t��˕��'�h�i���8t��������U�v)�l�]Nn0��.(x��fU�N`�[l[gkQ�Tp[pj��lms�n8\���j�V	�V�N�M�a�۬�x�9���mB�]�](c;n�����.97Bh�b��_8�$D����V%u���n�C+"�:��j��9�}R�HJ�����mʥ��X�tA��6�b��D;���Q^��¤��+v�Ǖ�9��8ٞ���u::��h��:��y�[{`�-����l�����nMlړ/��<',lwR��뒰��vM �����v.�T���%�Y����/K�ꓢV�R�YH[o.�e%���;)AEU��k�v�
�ՔL�e��9FZ�kP��mp�d�jx)����	z�n�����p�Jg�vb:ݼC<�L� ,��F��7+M�����v�W��m��lk�5:�!��3�0���D�L�q�H!O(l�\��
I���9,�gX@�T!̾���w"���J�i��.��B�`�n����5F0�ؤ(��Sk�Wo!��m!��8xI{]�lu�F�&�[O8zm�	�L͑P��l��� �S0H�@E�}=�Q:wi̜(ON�yr�	�#Ag�It宵d˘#��۫XD�����Y����B�O��L��UY���k�d-��ym�v��f)K�	+�ܼ�I���Ζ��1Au@��܎��-�s��Β��Lh�W�d� q�i�-Ѷ1�lmj���]6�:��Z���˜ݑ���Җ{"aܪ:4-��fӸ��*n�m����[m)�Y:v��$v�����ߛ���H��m�@�=^���*|��b��U������O��8��?	7�w���:�ag�a[n�s!���p�����V+���ʦ�@�����#j��Qt\�3n�P5v^�狱s�n����=��:��]s׶|Y������1�s�%�7N�<�
�s��l���lI8vy���.8W7�A���Ee��u��k��-�-�!��jAx+�Z�n]�X��n�&���6�<�$�Te;.��D��e�`SM�CT�	�WZ��!�ф%�˸]�[6L�8�-��y��4�l��AR��=��N�.ݨ��a�]�i��~d�,K��{[ND�,K����"X�%�߽�M�"X�%����m9ı,N�Ň}	�W����ֶ��bX�'��ND�,K�{~�ND�,K��}��r%�bX��w��r%�bX��{3-3��֭��h�r%�bX�����r%�bX���fӑ,�XdL�{���m9ı,O����iȖ%�b^��d�fY�YMCT���ND�,K��}��r%�bX��w��r%�bX����m9İ0dN��z�9ı,O}���/�anj:��ֳiȖ%�b_��kiȖ%�b~����Kı;����Kı=�w�ͧ"X�%�z}m/i��q�&�\�&uf8��m�<u��@ݞ��<Ez\M]����\F��ݓ��������ŉ��{�ӑ,K�����ӑ,K��u�k6?DȖ%�{���m9!I
HRBtG�U����]\���Y�%�bw�{�i�~{�EB�D�K=�~�m9ı,K߻�m9ı,O�{�6��bX�'�;=�䙜��֩�˚��r%�bX���fӑ,KĿ{��ӑ,K�����iȖ%�bw�{�iȖ%�b_ǥ�g��\&�L��k6��bX�%������bX�'��ND�,K�k޻ND�,K��}��r%�bX�σ��՗Rf�!��kiȖ%�b~����Kİ�1I_w���i�Kı?������r%�bX��w��r%�c��?>�|��ey`�gάkVv��:�՝c���G�YP����h㓍*��*��֍�"X�%�ߵ�]�"X�%����m9ı,K���l?��ı>����"X�%�Oz��L�o���u��ND�,K��}��r%�bX��w��r%�bX����m9ı,N��z�9ı,O}���/�anj:��ֳiȖ%�b_��kiȖ%�b~����K���]�ș�~��r%�bX����Y��Kg~��ڤMZ*U�WxBIN�����ޭ��Ǡ^Y�|�/Y"MG3l�w6��[�=��@<��.����C��ddc�(3m���\I��^M����]��=SG�[���m�R,q�"�/,z���[��s�j�*��"���LnG�]w��")��݋ {]Ӏ=�wXϳ9�Ȉ�o�dnM߭��9�h��= ��� ��+cX��<��7���k]� y�Q(���E�� u~�8nI9����ɝ�.�6�sn �s� <�����j���XPXe�F<�y�X�9��xsv�f�Ñ�j�Rl췜���Yڣx���8�z���[��s�j�/,z��.	Lx70jɠ{�x��(Q2=���9�� ��x��-$��d�G3@��ՠ^>X��; ��* �Å�f@�r�7/7n �v9 <�ye@;ط ~b�\�Q�I�m����4~�s@��ՠ^>X�Wʼ
����EN���p�+r..��V��\㫣�]��8팲]g�Il��q�
dn�b����M�;7(�և\Pv���.�m��;�� F�cѶ��7n��K%��Z�U%0H�/B)%h]b�T�P���O���ikQ׳l�0�ےd���$���y�J��]	�l<�TYj�����yv����=��c����i���=\�!��;�.8���:�;�\�=k���ƍ�U���}m�DG�x�7'�{��s@��ՠ^>X���4���yLjD�Brf��Ÿ��� ���>�ʟ�~�����x��ȗ�b�-��Ǡ^Y�{���>v��ל�5DĜ<����着}� �b���r���%1�����rh}n�ϝ�@�|u�זh�.^�1��
n��s�«[&��{Y�m��.�P��(��^2@RH&G0����ޭ�m:�=w��7{�`ɝD�U`Y���YsZ��w��;��*�&"�HP�B�^�_�3]��^,}M� �B�\�Q�I�m����4��s��^�t���V���M\�aT�6��������[�=��@<�ی��S�^!93@��ՠ=��@<��YPY���ӭ���ۧ7i��6�(էOfj���ћՅ�V�v�,�.Ftn&>�~_���<��YP�-��]uY���w�~���܀y�����[�<|u���E�)��d�@��tܓ�����C��PO�C�aDA�?��V o�^�mJi���'��h�ͨ{�gc��; ��w4��L�Dj�@�|n@<��YP�-�W%Y�p�X�������j]F��g��㋞���[;��K��l�c.5��Qg��v�,�{�gc��~�ˑ
<ja��4��s~Ďq�x���~�o1�l1��8��NL�}���gc�ܻ ��T ���h6;���7�x�c�>\����,BQ��m��?I�m
��Jf������ ����YPv-�����JР�b���ի�'瓑�ܛk
.�Wo�V��	��(嶣�&�b�ݪb���݋ ��s�=��_DB�!�{נ}Fgs���L�2a#��}�j�=��@=|� ��T�)��3 Y�z��� {;������qڴ��*�X	D�&6��C�x��3�����X����m:�6}�.D(4��M��ӹ�r��pt� =�� D$���K��D�[��;q���.0g%���<y�q�]��I`��\�B�v�in;u)[��-ڍIp��Иu;�+Q�a�+��� tՅC����KɚLV�z�.�M�o�]VC��JC��Ƶ�v�̶{I��]&�<��A���l��69[[�lcjڙ��p�\YMں0�fM�jy���Õ!�l�)%�d��̝�\�d՗Y��MY�� �3{�CX�;�ݫ��bt)�����l��ݮ�aMP�7^M$��ٍ�χ[�������~�}8��u����(_�7{�`<r:�<lsX�&��/z�-��[��}�j����g
�k�bND㫬 ��x��,9(Jg]wNΝuh����)��d$�@��w4��gc��v�SM^�����ѻ�P8� {;�˰y���˄M`�Uc2
ĦE^��7�uE�1+�u�ɹ������5Pb��r��m�e�n^n���r w.�=� ���J�Q&I����r٭%�����(U�[�ŀ~���k�@�����50�$��[��yŸ��� �]�|��g��*�6�
�3v�qn �v9 ;�`����qc68�d�n-���@���YP8� �+�U{�~-W���aۚ;C���<���np����/6Nme|qn�0�yn����Á����m��������qn �s� �u�6]�ǃs�E$�=��hWj�/,z�[4s�.(�I��L$��<��ֻ�-W���D�DB�Z5L���w�!��|`dֹ��$&��d�|bA�0��Hߕ��(A�B"c�Mi �懀n3.u��#'$�����N��9��D�i!8��"@COA��)��0b� �EM�:e8��h�h�L�"`p~����?pB1�M� ��(�
���E��o�q�I#$A�SN��4��B����q?90�pcdb9��k�&�B�����(��� �䀨~P]�4������ޠmE:����!�D$� �SH�V�~LD�������$�ݻ�ԏ�L���r-��̀˰������컶�t�2Lm9�[�4~�s@���rɠTJ����L1��`�`;�6c��C=��uT\iN^���pǭ��(4�9$�=�����Z\哹�{٠s����gLQę�nL�<�΅2t��x �u���, {�T��(b���@���h9l�=��hWj�*3�sƨ����IWw�ДDL���݋ ��s��$�� ^����krN~�Y�m�F��Y	$�=�������^�v޹�r٠^g0#Q$B&�b�#�ܛT�7��46䃭Z$9q��K���X�o��:��28Ʉ�g�r��h��-�����_(�xނ#P#NE�Y7]�Тd5�^�݋ ��s�?EL����1�rhܶh�w4x�+�V��[٠q}��B�O(��݀>YPv-��� �v�Ǐ��܉5���}�j�=S�� =���k\��"17S.�xG"�i-c���`�u͘���f��ƪ|nS�`�c	� (Nc&ʔ���U�D�Z�p�C�㫓P��4+�crO��ixNx�-�z�w%�{5 ��p���1��}g~�넸�֕�,��=N�;`���e��*t�4�:�M��vɻ=c-�/G���N���9k�W��n��̌�L�6�Q���;cf#�&(���{��u�����v4]=��Mm�`+�n�����+�g�W�=]�/E/2�]&G�&��.?�o�����]�}���=ط ���}��&$��Y#�@>�@���hqڴqs����Ԓǂs�I�}���=ط >�s`�v݇�Qȓ#��$qh~�<�\��Zȷ�@>�@����=��'��"5;�ۀ}gs�ܻ ��R�Ÿ1g��S&QǊ �)�Cj-����C��3Ɉ�b�=0(�t�!v�o <j�m`fn�r���H��������������F6
a�I4y�MТ�P�(�.� ��}��h��Y�r٠{�q���f7"N�374�{�n����r���M���ر�%"�17�s<�|�{4����䦁�mz�υ��x���B94�٠{�JhVנz�r�癞z��q%��i��K2")5�B�a�u7>�Z���ZZӲ�4�s�9�N3-H�x'0k!$��Κ�����@9m����e��28ɒ)e�Y�2zF���u��m��<�1#��N�'��"5
H��[׹$��� ���*, 7قD�9, ~ �o���nnI�｛�s�J�,A2Lx7�q+��h[:hVנ{���@=�R�m4^�[�� ����u��������=_T��L�B
I24c#:՝�d��[����Nx}(�I>ͣ��v3<b���374�u��������>��8�̩����D�M��qs��(��S ���7|`-�Έ�=&���top�,�Ǡ���=�%4�y�x����@��z>�Ԓ#	�V]��rS�� ������.!�؅䒄�e�w�7D4��]��utZ��� *����`��>{RϹ1b*�C	��ǎA�449�e�&��y4F��:�-���4q�ZW�8���hm�n����`��>{R *�߼i+���2LcNM �٠|�� U�������n���1���$�h�Jh��;��y�%��h{����7�� R%6ㆀ*��=��]��~���lx&��#̍�ɠz��f��]�{=�� m����I	
�"��!(E|(UB�@� �h@�*{V�$d�˞�gk��ǱfUd��j������ѻn���g�ۏ\s�ݺ�
ú���';5�
Bh���K��'h&3�;3��O&쎿ˈ6�|��*Yn�E�jj�g�N�C���6pح���C�s�M����2���SpV��c7q����v�e�AnB��Ft�G���d)�`:������4ÕŎ�+��ڥy��&L�f���A�"k�h���l@�p:z���XѶ�`G5��l�g�:����r\��]�u�|�^ދ~m������Ĕ{^q����%�=&����$�ǂs�I�{�%7��y�C���I�� n񨄔��Rk��!d����mz���h-�@��Jh╋7�Y�$z�{����>�j@:�����Z�� PLx�$z�l�/ܔ�8��@�3���3��4<��#�8�^�;��O����D��Y�]�n4v�F��7q΁��F�K�$�h�JhVנ{Z�z�l�/��`���pMcoY��'׽�o�00 $bB(�D�E��T�D@8����_������/ܔ�ٙ�g�;[M�0]R<��N=�z��٠_�)�q[^��/�.x�I�ȔN= �h�JhVס�w'V�h�c�I��d$�@�rS@ⶽ��+�m���h�]M����WE\�ظ��.܀VP�2�D�lt�EĦ͇������u�(�C#�1�!�w�z��^�r�=�PZ�;��ӬX�F�AI2�� �wl��R֮@>�a�W��&�6��@9m���ҰU�H�EH�H� ��A� �  l?�B���{7��{4�e�
	��L2I&���f�۬脽N__��
"e�u�E����5kq�@ⶽ�g���z{����M�}@K��,u��`�HNm�]��
��<�7P=�m������鍺dAs؊{�F~������r� ��HZ� ���}�Zf�<�D��[f��䦁�mz���o|�H�:�D��<�5��M��� j����`+�ޱ(��n!�c�������z���h;��riE7�XRZ��BQ�(I��^s���D�UXF�AI�����l�=���8��@��9O�MƠ�Lc������ FW���%��Cû[T���q�:��	���@9m��������<��ʫ٠tΆu�Pm��$� ��ٝ29���=._^ kn�
�qଏ��5���q[^�����l�=����Tk'�U#̙yy� ������� j��G��1b�4��R'&�r�4o-��n�ӳ��WF�$�4�	H�`��]���p����`���`��@ H&���(be+����4��PD@�t�?�?8�|.~փv�B���5��BD�I�C�Qtҩ��l�D�UR�,H���q!���h�A \B�k��pO�J���|;O�C�	ǈLI���4�h!�}�ֵ�kD��L�Ʋ^��[�-���J�l۴=�mɱ��6kA3D�I+�Yڴ�q�kNݱ'b�MS�J�ڇ^-�E���$���l�-��i�ø�\A�Q�UG2�9�1��̺���N�x��0v&PwZy]�q:����m��n�uQ�	���E�=l�i:up��%6Ɍ��ak�j�	�-q��ՙ��g�c�l��`Un�x-��m�6��GNcmO7Wv�u�x�`�#Y���Yz�e�:ti�v�d�B�����^�5P�)K+�R��Lyl�).Q]���"�]��[��/l1��K��9��1�[:9���c+��N�#Oje �Q��d\�l��"���g<��n�s��	�]�n�Hrl�ೞjyC�y�tQ�:� O��uU)��t�&�3�]�n<f��8^�U׭�*R��m�-!s�Խ�e-���u=B m8*s�ɮłi$�wTU�Ԭ��=���FxL�;�X,+lVz��[H[5x4$�����[��l�Ͷ�Rɪ�jUV[�� �l�����/����W��j8��L��S�,v�-��0�o�����K%h��z��۶�= m�s�Z�;x���ÐM [�T�ꐧ�Vj����:�T&X��Rl�Ѣ�YI r,����F�h���kh7k\���3����64;`�ukv*�[�s6�S"���=�$7*%��6��t	�����AJ�g�BRB�#g"[vݰ�<0ȅ���WYU.ŉ��!��Y���m˞�M� /X�l�Z����3�nc9�]���>�۴�0�O! Q\������֭�I��a��]4���ñ&��YËPT��l�#揾����9&��e�lt�ks��hӭ�b`�:]ۓA/F��j�jqۖR�5M�k٬u���-��l.�"2-�g�`�Z&װ�1-�Oc	g�n�*,�y'!ش)��" '��T�Ѻ=v�J���R�n��X��� �*����ɫm�-�f�Z���?)]�@?�
�A�>��tS@�&����B ~M��E����_�O��g3T�8�vb���
ո�nc����d.�v�۱��ȝ��{!�mq�d�H>�dA�ӌn����]�K\\�НU۶�m��.�vɺ�����͐�u�nz�C�x��u�d��6��qW���Z�����Z��ӗMl�����<�u��(s��ld��k k!;\^�Cacq^�5�+�m��=o�p_h�V�W�Oc��ͳ�ə��K�v�����}����s����>�b�g�`�3ctE����Q9��p�%�j1D�!%1������p{:hVנz��f�r�4�L2��2Lʽ��֮@>��v r� ��H�)ZC���$z���h+��Ԁu����YmX��y�՗{� 9]�|���\�}|�f�{����Pm��$�@��R֮@>��v r� =��~*��P�[��ntbz^S�����(Gf��)PW�..�8�I����;	>KhY��o�����������>{R y���/*�n��j��rN_����P8
E�J�@�@��Z��M��H��b��H�G|�Y��ܓ�ݝ4���s�ď��,�cNE"rh���=���>Vנz��f���e$�ڤUZ*U�w��ID)�<� ����?Nλ���[���vN�n!�c�������4r����M�-Ka��86�<�a�v����7�5�����mqמ�sݎu��$Pb�k��盀��)#�=\\�@�-��=������Xqw�z>f!w��8LB�݀w,��j@=j����`�EQ�!A1c�s4o%4����B�DE�˜����`,ƚ�ƦA1�4����.Y�s��h�Jh*�ǂ
�di�2���~���W*�ڐZ� �X:�Ń�M��x�g\`z��q��/X�Y_[e�Y9��s��t�{ov�vܲ�=� �������_��0ILx70k�����M�W __; �YPޱ(B�3l�v��ot�z������;�T�4np�X�F�AI����I�����9ߵٹ#��Fp}��נs��+��"p����9n�� �r }�; �	m�[:ʼO��&��7Ńp\�ס�S g�7/KPs�Γu��Ͷ������� ����9�rʀu���d~%2	���|��{�fbA�/f�o{��{y)��`��fF�wX�Mw�n���>�|`��8�υ�b��Ӈ�894r����M��Z���h�2�S���ͨ���<�����`�*T<�	��Q"��!���߸ ���];���.3Mˇ$/^�v��mv�=U��n�nQu�Q�=���>Ԙ6��[�R�i�ݻ��b;��I���q.�Z;���`�鸮Ʈ��!Q�v�]$��re9d7]n�O�X�-nRu�-��Tΐ�h�n8\�Y������u�9q���6^����[�����z��Q7̧��[<nzg<�+���fh���W;����»���u��}�;〧�N-��>׳ڧ9/Mz���$<Y�/�o�g}%ݞ)���u�xf��������u�X���ZV,xނ#P!�@���{���ċ{ذ���:ns�"d�Ф�Ru�7�`�#�-�w4��4��h���@���2�(7�9&h��`t���5�(����� s��@�^F�7$�/�@��r���� ���������Lx������ ���Yq�W�K<Z�.y��z)}Ls��c��247���z9n�{yf��v��g��1eli�ȤNMu�X�Q�*���]k�����fY�Jc���^&�h���:np艟:�Հ7݋ ��N�����˭6��77 qn�Ü�w,����8V,x�`��G"�9�� �	$���� {�^�M��{�p����vQ�A&��C�Ps�f����q.��,��v�2V;9�a�Vء������e@�v��__;?�(J&OGWP�䛩�*�.��`���qn���� �Ap/6�kj	��hWj�=\\�E�d�<1{�R���b&�%��gb��׀k�<M�%dY����W,�9m���]�}��� �Ij�⨙�#ov�v�ʀ<��u __; �V#^!e1%�E�$iL�V�������qm�q��V�vZ�s�۪�v�&3��� �����Z���w�����֨��q�ǉ�&��v��J�2z\����X���Z:<{0Dj#�h�.Y�s��h��hWj�=ϝX��a�D�1	K�u�X��Λ�Q�� \ �By.DSC?���}�g�x����\���R������<��-�>��vܲ��R����Y�ʕ�v;�:��ń�מa,!Z�O&�ɂz�}�jv[x.�疯�yŸ����;�T }��o�x6`��fF���=Ur���s@��W�}]�y�#8.�u��"�f���@�9 �p��v �̳Dǉ51�&�h}����h�λ��J!(���,�zYԊ�����H��>�ՠw<ϟU��{�� ~�xY�(IG�&GS21Uښ	n�'���]H�uI�c������[�c0h
��d�ݤ\YX������X��^�Rmτ����q�0g�k���Q�v�j����U��.ۊ.��.B�Ge �(�]u��z&��\�k��K}�&�6���Q��<3�L�^K��`�IΗ:ygS�W:ӴR6x�

�áE�R����nW��9�gt<����qO�T��$��u&]YI���v;;vޭ�ũ67J�[[v8��ض��T�ŵ
pF'�LH��G"�uq~�4r�� ~�Ȅ�_�7��p-w*��:�/s4ڲ�w`�* |�8� ���f����xc�I$� ����[�q��9YP��o������fn�����s�y� /ܳ@>�P`ق�G��@=��r���v�-�6�Ǫ�]�w�c���e��������kjv�nv�/D�<�%ͬ��z��H��L���~~~U�u�ݐ���	޾�y�v����ܺ��f��'w�����
���W� ~s׀ko}
""d�eu�D!1�I�^��h��4[w4�Y�{r���ɉ��Z��w�k׋ �x	K�}8���UI�)����f�� ׯС(�������h��4�pU�<y�∤�ɍ�ݓ�vر�c�.[n��]/f4u
��$�!X�
	�8�L�yf�
"&_S��wO_B���b�6x;�Ӈ�5i�M�� ��f��˹��� ��F�l�W#̍E���x�x��{R�N!@�D*Q�N��C@�E(s�b��*��t�z�!K"1(~T#	c�Cq8�Cd�^ 5�~5�8����Nb(oF�` ���iL���@��RWSύG��F�"������������(�P�B1 }��	N�j�s�@60Ǡ�R	9��4�~ %G����bl�'�'P��_�������� 'A�ء ��<��@~�w�}��;��V��#��ŕ��$q�4^]� o]��\�}	%>�]�1�D�y������ ��f��˹�g˙|lē�����rF�=�919��r�D�q�b1f��Q�#�f'�mDB(��+�Z��f��ǋ�(� w>�ܸ�&�e�KU6^f� �m�<ʀ��9�n�q��,1H�'�E&��˹����� ��f��Rı�ywwk �x��=�@�t��5	G� ���"0H���J�_��X·�ULՑSsu54��v�sp�`�* /; �Ϩ
��A�S2)�Ɇb�Ǜt���2ם�e:J���c�]�ڜ)ؚM�3F ~n]������пH>�Ӏy#(��Y�ƞc�7&��˹�H;�٠^�ՠڬ�/,t@�1�D�y��Py�9��>��`�*�#�U�6�!	�RM��瘯e�z����`�* /; ��p���E�Yznf� �m�<ʀ��5ֹ�<�*D%	�����9��s��D� �j&�+[��]�,�搵���k���_7nR�ӧk�˧mnl�V)}����N0�m9Z�%��'��w(�q��'ˡ��l����1�Q.utm���n��2X��n�v�����N��+Bl�-��t[��a�YE�(�s�q(p����ڋ��s.�CZy��������v�D��K<�N��*���︽�ی��вv����M��9�&� �S��c��'��v��qP�g�Zbh��"p�%����s@-���?��?HWt�*�L����7wv��s��-� ���y癘����[I�Ƣ�4�I&���� �n�s* /; =^�.�ī�y�c�= ��f�~���yf�Wܯ@���,U��cr5&���Py�~� �n�;�e^��m��_]��ްJp۳�A�]�c�����;6��G5َ�F�qsɯ����?� o���\v ��P��mX�j"!�I�q^W��g�y��e�߷F�rl�e@�`4��I�&5(����f�~���yf�_�f��s�cE�$rd�(��s* /; s��`���w��X��D�cɄ�L����~����˹�w�{@3�1���n�]��r�k�6�g��Փ�t�� �gÉ��rݶ�#bp�(�M<RI�y�� ��f�y˹�|��@>*\bi
��7w`�; {�PZ� .ʯ�y��f,U��c�7&�y˹�?^�����^*{K�*��Cg��׀t��� ��w"%M�U%ĕ��P>��-\��`�� {���\�
4ڈ��x(����@�$������b�?Kn�4��-N�˸α�7A;�8���-�4]���g2���;]E+���˪��%�C_m�-]��ʀ}j� |� k�n�����92b�h�������l�*�ɠs��w�0Ǔ	$� v >]�}j���T�B���⃂i�M �[4U�M	߾��ɰ7�j�+Q
�A"�������{�ܒ~���.ZOM�I������w�|�(P���� ww^ ?7x(Qk�O���(���`�m�����8wӮ���GE��	�j2��H0�lǑ<i�9����� ��`���+�q
l�/+,��hfm@�v >]�}b� {���.W�F�Q�RM �;��?)m��D�7ذ���L����D��l.nj��K�B�WwV��s@����l�.sE�$oM���r �2������^��$T����!�,���c������ط-vĺ��"�x���z�.�-qV�UM`q��-��ٞGJ��7��Z��KNi�EIoI:��:0���<[l�t�;y,�%5��:��9�3�d.�m�D�dÀ�	��;]Hz��gv���m��&�,)I�;l�`�ٮd-9N�F5<p����R�~>���G�\<.:c�TTV�^G`x���\��4MY��o�(R(�{�8�������A�녣q�(��؝�����M��iw/54��<�ۛ�a۞�Uv��~�������b�Xř���޶'L�@;��h�v �2�����Y�am�埶��݀6+��� m\��4
��ǅxۇ�B94/��#�e@W ��b� ���2��ڭͨj� |� lW`���o<���ubI��X��8Ѹ�8�n;rt8�*�������烈5/N�ӯףi�� ~��M��4�]��k�=�J�ǳLq�NM�;g{�oc��A�1U�`ThB(P���?u�� ���Հ�� kY����JF�1�h�]��k���b� ��9EcE�Eem��P�� ���6+��ʀUB���⃂i�����h������� �!B�\��fhU���b,�܅5ջu�pmV�yŎ���pd�����O=���	���I���~�����s* ڹ s��,k����?m鹻 }̨�� }��E�h��i�XL�	��m� ?k���(�$�D�I}׀w/w4s���Lx�rh��`b� }̨���)��mmf�{{� ���e@W`���>��.D�u!ū���Wji�F�q���71n��%^Yyy��<9�$#p��I=����[f�_�f��[f���ǋ,�Ǔ	7v�+���v�+��ʕ��U[��	��I4��4X����ns* r� <P�f]���Y�ܽ��X���T �v��GpbA �H� ��	� �b���9��?Y'g�0��35]���� 9]��`b� �;�������7~�={�ծ�H]���^.wڜ��Wd��m����t\��ۑ�h�G���կ��� ��dm�(_�;ow4���:F�x�6����z�Q��h����l�=����ͬ͢ܣoo7`b� {�P��~�h�3�E��5	��@{�P�� �v�+��w)e����a$�4�٠%~�z�w��'߿}�rO�QTU��QTU��U�TUsE_�U�(�*����*��
��� ��@��A��@ ��+S�ʊ���⊢��E_�EQV�*��E_��*���(�*��QTU������"����U
*���b��L��h�P�� � ���fO� ����  �UUU* �D��@AA �-��UIP�
H(T�EU)@)@ ��D!U)D��*T���P($P�)T ( R��
�     �    
a5 i��Z�6��uﻩ{}�oe[���Je��:�Y֝�tzy�p �طF��:� y�.y�=�8 z���ܳ�k������^Z�� }}7�����{��n�{�����<�   ��U � �|�sg�i�Uڳ�Jrn0`G�gbk�ӛ���j�x k��z�qo�z�k� ��}����x��[}���m��3�&�5{�}�}<��� 7)�}����uz�ů���e� 7� P      ��_ks��I�{}t���y={K�C�Jd��\�盫ŕ������|�m��M۾��{�^ ��iv�[���>�}Ʈ[�wmy��ӾΗ�׾�_q�@�W�]sW���u���W� � � 
 P(  W })^���+�wԥ唥��R�` JR�YE)LM(R�YT���(�B��(�)@�Ҁ )K,�(�ݹJR���r��14R���
Su��biJP� 6R���Ί
14����R�3e)J �
(�QE
�� ��R���$�ҊR�)����>����r�ruKz�}5�wS���J����Ը��{{��� }����}��iV@=<��[�+����Yw��帲��� ����]�s�qg}�������^ ��I<*UA���hb'���T�A�F�"x�T�!�0�&�"{J��5T�F�"����z�)H  A1J������'����9������1'g{��{�}�� ^�s�( ��AO�( ������ X�����䅉bC�̸ͅ��	�#i�cP�Bҙ�B�CX����&����>�q	-���d��#XS,*`a!I ȄŌ1�\�R�9����&�_I��!����CWw����{�)>����#��c���e��W#!����&���]$j*�d�B���]6Nv��!�᜚t�$p� �)�2% �R0Ô��^ ��#�%0�B�RF\2W�k:.xn����qr�Ƥ�a4(F�I0�,@�!Z�BEBDc@�Ќ�D!a~X	CaHD�b8�63��n~ųK��\��HH2AjF1I��9M����:���Bi���eY�b�,\�č���n���hJF��Ůd�c�c����I�B�����HWLyj8ԠB����)�m����(D�H@>�0���w����	,"��B`�F4$3��B�>x��
�j� �.	fna�P��B�r��Θ�9M�
7y%�AdhEd`V�H&A�0�i��ecSD TÓd�B�.�#L��\9Q�х\1��VI�#���`�H�!��X�ddb%RA#2�h�BF8�Q�"�4�D$ #$n��K��B5�!��]�+�Y���G��0��!$����) ��B �G	
`��K ��H
6kFH$f���S0
���FH��B�d�H�1�Σ4�%p̭��1�W�Y"�J��c���>:!�Xh� �L.!]n��K��'�MG����zY�ŏ�b�9���j@�\\����Sn	P̣!lJ���f�%&��2\a�!D$�@6����5��J�p�1�&I�hFc�H������C��$,*�T6�F�jƨbH��J$�����$��	�1RA(�� ��c�D���ő���d�$X�H$#�jF����*��i��B$"�*H�ґ�S�%�h##Ce��E��h��!J��&5��0`�6�d�L!`C�8pkz������܄	!�Rz�.	p��� �`�/	�/�T���&�G�=�eǋR�1H�@���k[#��Ɔ!?��Bq�*m}�W؄Ԧ��lR��J`KL6\��hL"WD�q=i3Kl���M|�2cD�!��q�,�24�ɔަ��U&I���R��7�Z[� ��"U�@!��1���D�Q���"��R��G� ��a$��!nV��pe�0U1���~*�_�j���r�dBQ��j�Y��J`f��E�����je7*�6�R�v�50Ǒ!���By�'Rb�u�!�S��>>�s����bȑ�C#\���z��ͭ�x�E!�U�H�1�	�
	S@ġ�c\/5�rh�d.ȴ����b'��ΒpG���}�St�Dζp�W�AU�Ĕ�p��nH��അ4��󚳋���okY���*�eܦ��Qk�i�JfY�Y Q|'50�~1�%�Z�|G�O��Ԕn\'�V�T' B3�!5�ZƇR��|a��0��P���If��!H���U:$���`Ő��Fƌ�����Y�b,cXP XBj�8aHV!��H�y��Ȳ4�c1�I�$�M����L�cC]|k,,!��D�F���((F�*Q"D��ȑ�/�������l~�0廤�5�D(A�2�Y4�Ə�v|=��D[s��j�����._�e-H��)X�(B�)�x#	�֔�+$3Af��o�f��HQ$$��������g�k  ��0b�iIs��x�	L9�.4�%YS A�Ms#HM� Ӻ�#�zBx&-LB&(��i�A��46�����5�TZBzZFK�*���@ݯX�-��_���z����$YF�
|����m|)���u�B�K��8H��%+#K�hX2M7ΉRc��&�"���&����Tw_]�DƘg e���;����H1c�-���)dIqČJK��1
jB$!"C�+��b�ă#$
��Sk��dhF��!Ld ����,�b,�4�t��tA��!h=�K�Pj}�O��^!8�1&���D(
�FG-B$L8rlUċ�,B$(A��ġ�� ��e0c��\gX�Cy�+)��@�Yxp���U�$�����b����&�c10�B�t�jc0�%(2B3�p�c�CR�	��
��+�#A�Q#ZLc"F�(��H�\����$��"$R��$�,������6b`މJ,б, ����.cM�Ɉ��#!!����+��p��1y�i�X`!\!
�"��$�_�d�3�FO��.Mh�jA��h���π��HSF�8a��a!aB�aBR4�>bS�ń,i.3p�'�ß�Yj#�ɡ-�Q1�5� ��$�D"�"�.1!��F�2I.L�9#Fm���j۟���K�Ɋ$���vΡ��E���_��4l�z!��L��Mɲpo>�D�eI0n$8�BKW��_��&)t}�YlI���42I)��L��c����)��p�ˀ�F)"0 e�BL~//k�3���D
a1�1N�LI��0*S8�1��pXm0S1����F�*�K�,��J�b4�~5�1<`�iKsHMߴ����~���!�L��CB�i�Ld_۹̼�oY�u��9��.Cd)���po�!�@�R�+a!R�����S�ƀ�\&B���Ð"���b`�\Ȱ�:�H?|;o ���LH0
��R9tl�$.)q�\`9��B8��Ϗ�W]D!��֮=�L�e��Rւ�UBH0���ɔ����##!bE0�
��5�!P�#�$3�W��f���|��iX5jGxv�j��+	�$1���U�p�c�, "�,"�E�"�h�"`q�� �b1A�q`X0aL�� �~�Y>0?q1��+�R�0a F���6%$�"T"�!�b�:B@�g�+�e�i�.��L}эV4�
�5���ϱ��t�n�XR,ay��@k�fE�	������{C�>_��Ia���Z0�`F:d��F�X�jAb�$
&3 ��4e�p�,�aFIB�(@�\�5����~7�y��$0`��"T�"A���>`č1#��!
abU�P˔�F	cG���]����/�n��������q��ad�h`�\2d�3�$C&R3�$2aD�^$$э$$��qa��N`�B��ͅGh.�)�tY�f�0)�p�����S,u4��Mꄧ	BT��#X��
߆ᑲdɣa�3+�W0�َ~�C���C��iR���C�&��	#�۟9�Bz�5r�?�����M�K{е��#��ƒ���`J$n-i��9����l�H�萡�b2@��'p��#	7%Lii}WT��Ҵ̆N�F��- 00 � � B*t:H1j���cC
bH$r�hE"������BI[X�l�������H�X� R��+��`c2����0ˍϱ2t�d"A ��]4��"э`ф-B�(�b8,V�[�h��9U}r��1��w>e�ݦ�p��!�E#� D�@���$c	"V`��|ҝ�ݬI���
`�׮y���        �   ����  [@H �    	m����-�֮؛\�x m&À       �  �m��J�a!WJK*�������� 	�kVK: l��ڶ��M*�<��u�KӈM%�n�0֤]��K�*hV�Bj�gl�� m����XÖVV�	���,�� ��T�I����azY#�v��� )V_����@eH���g�H��vI����W!khnۭ��۴�q����MU][���f�	 � ���h��� �`D�-[Pd��3�8[u�u�l -�-u�E�q FNqUHE�1�A�A o\�� m��-���Hl6�a��	�ֻ MRS��`bN�v�e�JZ�� H�m�۶mb.�%h�m�4��m!.�  6�i�Ŧ�Xq�i[�����r�l�    �n�d�k�*��P�
ej�������  $p6�  �j��a��W�U!!@-�k���_�2/�J�����Y����&E�[I��$h @��쵶�lI�����N]��� ��l �l kVf    ۶���];` ���,0$h ��m� ��&�,�����PE@!5 �m����h ۶ ��H�$   m�m *]�j�
���/&f�X��t����[/ ��u�`���[@�m� @    6��e��   �K�m�k���ZyZ��C��jeW��ポ�y�ح.�k��Xä��Z��m�+fѓ�m���:��`[At� [Dk�m���j���W��eZ�)j�j�yP�Žl��إ�o  �հ6ےslݧU�/K"N�8�K�͵\�Հ �t�X�f��5R�vҵ�ۜ���2�4�-�m� kn춛f��� 9�[�����M���^:���հ�� m�H��������
���m� n�O+|���I��'=;wS;V�Q�n�v�"�KHMU\^m�t�`v�Z�m�lM;v$u�\
�u��;n�j�`IuI%��u]$�E���O�D��9_n��	If��H9-�U��8Jvm�[D����C�ۤ�o� �����2]lY�&H�k�T�$H-�� ���T	ĬUW��V�a�Wl-�i;L�`�]���cv�>��� m �[dr�Ie^����>�c�X:��I��i�[Z�8�l�^���-c��l�����q�&�;�Z��ۥXZ�E���� �E������6��s�����)�H�v����ҸkoT� 	ep   �d��I$�]�9�6^M[lm&� 8� [���  h'm��N�6������"8�mm ��I6Mn��4{^����[I�`��jAm�d�r�UP��r�[/V�S��]a�ܛp8�@� 8Hp�l�}�I~�Z�U��
��#��	Zԫʥ.��e�����5�vU�`�W�6�h6�d�H  �e�g,v�%�i%�6��WCnzۛ������cd�b�'�9k�K����H����iz5��` 8 [Km�N��m �&�ִݮ��p  ��m�h�i��ඤ�km�m&շU�`���)q��׵��4�  �/S`�8��lm���Ŵ$i�Z�k[ �a�� �ۅ���m�@ �5�ɐ6�m�     ��m��m �`䁶ܶ�׫	,Q�T�8�WHi'j�2��[IeӯFm�H��1c]n {N۴Y8��x�����+��IY��F����^�K֚7}�s|���-�]2�;r��Y��9֒  �����5]o-�][,��ѺP �v ٶ  ^��9 [UP1J��V�d[�i��j�hmHq  *��cP�ڇ�SdͶ� m� Im���@$��d���z���6�Ӵ�3!� $ ^��bY,�N�s���ԫ#�gk8����� ��r���=�$�(vq�8ڞ\� �M�i�e���fZl���� [��e�p P�4�	$ � m�Z�i4��	'H����R��ҭt�,Y7ij��U^��:��wl�vs*�a��%��<�l,��	��T�lL����rE�m�v� Ɗ��:@�)o�5�����	l�W(� q:�P:B��v������x6���V�= ��� m�-��	�]M��������8���FʽUK�U��'hh���	մ�����ve皫�l�p�].��l� 6�kjI%�L
j���� -��t��,��:m��K#n�m����m�  � -��׳���U;B��UZ�����@�t���lm[� ��  ]3i0#m�%�� ���3�gj���3�Ze�b�j�_���a�)�k3�m����-���H�VX��TkX�d��N[�ޣ�M+)C�e    ��m�����k[]���r��f��R��J:زSm�ᴛ8�#Eh>��� m� ���m� � -�  Hm�m�F�n�  �`�m��cZ�]+[cD��p$7Z��*�  p��kX���   mS6�M���8�d�� 
�ׅ���fճ�f�3�5�cMK�n�Z	cI-�j�6]7k�� ��� Κ�j��[�\� lHU����Si�t�����h�D��y���d��ʴ�� aE�����J�@J�S` [tU:N�h6V�D( �õUUH �6�@�`&;Hd�mo\:C�q!"�f����S��;�4m��2f�k4�:�0w��.=U�����s�^�Phlu�[RM���T��Z]������j��95�&���` l�m �@���Í�X����$��� XI��gm���hJ�6�Ɖe�ͶҎԫ^"v^�]�4GE�7$��첃�i�(H$�m.�ݻI���n�<�S���P m�m�"ڐ[%[Sm͍��mU��<m���H �`�  8ڶQ��@R�
�uk���Hmj`]4V�^��P��u� k�� [@ �jm�:R��Yն[�J R[-��l�\$�d���`6��Bڷ�	e�����^� ^`�v#
5@l�T���i5�[@  6ͧLm��q���l����n\��;EH��i��@xΩ:m�-�[��`��O��� oM/<�R�UW<Q ԏf 
W�b���ԼT�싯('it-���iy'V����l	۵l��BCm� -�[Eᗧ`�"fl#=UWP[��:F�֦�-�� -6 m�   ��m��n��� ��ȺN��.�V���n��jjݨ�eeh��]*��$8      m�m��m�e�Z��­�3ɮ�u�:t�i$�� �6��}�����1����0��z�l��Mn -�� -����6�i�m�v�@ 	��k��W��[ 򪽵][mV�  [\Zfر'�`�� 	5� -ؕN<UUT+F+g@[������V���� �
l�Jl�e��S�Ԁ�D�&22u�����lD��9��B���u+���	�
�iv9 m��]���ඃ�Ѷ� �La���`ֶ�	m����X��eKm��5��$6��hl  ��N��?m�� t�6�h/Z h�im�۶�q+R���3��S��(,3ԩ�jZlհ �@�lۤ��� 	l�@  m�;tP�fΒ_FT�S@�o�� m���(!ri.�K�Ā>_��-�������kR`�2�h�   � ��F�.9I�ms�:l�e���T
�U�� �� ���mۜ����j�$!oP 8�6��`�7I.�f�Nͻk"m�D�"ŋ���0  �p U�K:�am���`m��	$HڥYgf� �$$-� qŴl�mH�ic$�ܬm�v�8�Z�"BM�-���e��`p-��  m�m��gYWVR^j���Q���ڰ�	ۛa�l#m��-�m�H艶m� AKU:)V�c���J��i�$��3$�!2m�K�-��� $6�_T�6m� �[��c�L!����,�R��V�s�FDm��MGNY�I� c����ZU����V
2;.�^m���+�����,6���b@ m��[�m�,���   J+e��.Z����m��6�8d�Y0 �v��K!��4� �mD��kM�v�'I̋�m���׉����kE7��fI��n�i2�  E�ὶ�\ [@-�	 6܎�׮��xm��Hd�?�g� ����� +�-l��啤;avٕUj��m����ۇ ݶ�����)�b&�@؉��!���4��P!4Q� &�]�j�b*t�B����T����p�H�pZ�PuF�u����S�� 'ʃ �D�?
'@~4+�8�@"�HjP"Z����)(���(`����DJ� d���� ��4�qPr�����FPS�(˄:B ��(�zpD6�L� ���S�ت<A DwHE�+� Tx�Q��Q��A`H���p@��̠�P 1�F|����x8*�C��P�/3ÈO��x�H����@�� ��0�5)�z"��_�t
�s���@z�p��@����A�?_� dGa�������4*@��	H,*�����AL�<�  ���}�O�'A®��v���D��@��4h2(F�E�@>TW��C�*lWy�D�@舝 p���#��2�"�H�X�A�"�D8'���@؂m��TC�B�lj�T�Q_�\�U@�b�	� tTҋ�g�T{�BZ��O�hAH�aj��hAH����Q��һUC,,A$�FW�����;9���A^�"� q�@�*�8Ap�2�X����@�@(��t�������U�_Q������Y�{��V�� Xgm�m�r���ϭ
��*Ѹl�����-���k 4�/%�t8�<r��.��.�v��l,m�U@W����Έ	[H����4v�������p T8�Y��R��v#��ۉz��r�vE4�� ��	���9���:�;NG&�1R(��Ap!��ݨ��R222�+,�q�qÊ���V�i�]U�wI��2n����ۣm[ KG�:*��=<c�1�p[:;v-͒�k�śBin�U5��:�.֭�
��ʀq�Eml[��RZ��%���h�u�s�i��tP���V��Nݽ6�S�m{k���/Sm@���R�ʴ��XL�1K܆�v�����!�ƅ�4���m��έ��eAj�*����Lҭ���UP;���lz�t�+��ا�m]s�:y��������Ed�G4��� �r9�3��g��b�&V0^�	=�:��P+$Jl��\�n�2������� � 7����w	��\a��6��Ce���]�*�`n�i�6�EX%	���`G5��%�]��^�9��V�p��hL�m�^eU@j�@��Y��t�:(V����Sp�F��uU�S�o;l�y��M�P�[J��)-l`䶎�5���Kű��X'�Ŝ=�(="]�+l�^x�� r撌qŶ��a-sO]�g�I7n�\��[@^�ەt�x�CM�\m��=W/T�;2FJ���>�tD��i�6�=��JO=�@�̍��ztTեc�5�U �P��U�	��n���*�jژ���u>;AV��!�qn���^^��� �Rƶ�=��AU�����\�e.��N�1C<�iY8�F��5PK�;���[���U� �7Ue��%�P�:�J/��e�͍���Wļěm��/7v��n�<�'A�Wh�¶�:k"��(I�J�nrgf�Aq՚�0]�F�ei�x3�KUu�甘���1�cT�9�dʞ@��] �ʯ�;�*Q��U��P����A3��pʌT�AT;�Y�k\]vb��tK<s����L�5$���K�:lZt���(�Kev�����@�am���ۘiI�^/Cv�"%l��;K�q��l-�l���^�����ݝږ�p�3s����5<X�#�7f�q�M�g/��{n=h�v^�p��G%���pb�n��8�Y�q�Cɘ���r�����MYt�8k8����C��w��L�Dʎ�&���1	�e�,8�n����d�"�Ȝ�;�(ûs�6Av����gۭB6�����/{���_�%<��D�qₓ4Wjߒ���;�)�r۹��\ ���AUw(u�@n�bj�@\\Θ��	��X�94��h��h�ա���4���0�F�wubj�@��u�_��'��pa���t�R5@1ިG<Ȳ�$z2�&�׫W�wѵ�q�-�ή{�䚸����ݠ7]����0Y\�jH(�ԋ@;�f���δ[h`%����D�&���@�{w4Wj�*�B�Xㄪ����� 1�����u�vԵ(�6������r۹����Lu�(�� �D�}� 3zf�l�țn$�PRf��]�@�m��9�����h�;�F��A�9��~�8��M�N�ڭ�κ�81p�uY�ƻ1��0q6�LL]��>*���ڄn�n؀��ՠ\\��5r#k�L�9�j�P��i�@n��t��r���Yd(B�V��{�-��8�?��B� B�@B�Pֻ��F���3٩
�b��G��"����V��۹�w�S@�s@����Ȇ���%M\�7[P��v�6� 1ֹ@U�$��"�G�<�b�Y�(kX���� �Q�,�Z��OYl�Ѱ�H[2D���f����\|޾�P��Z��ڄ;jŤAII�I�������2oS�@=�P��v���m�\�Eq$҄��9_j�;�w4�~�ؕ留��ƀ[]p�,���q��l@c�b�ވ��DLG�.� �L
�����RM�����Bdm`�!ɚye4WڴW���s�Z��Mv:�Q5S`��ӵc��O<�l���Z�4���7B��Е��۞
��do��>�w�@�}�@�-��_0��zh�	�GT,Q��i����mBq�9��8�Y\�jH(�Ӌ@���h��ٙ�uv���ZNТ��8�G3sW:=/yp���Ԁ�Z��6�@�mX��#i)#M�p�8���u�Pcj�؀Q#`��#ފ��g�i�>i��H�(۵�J�$C���7SKc�������*vtu坞y;��t�Wps<<٤V��J^8��K�'�<=��wN��z��+V�8�Fu�z�G�ӻ=3t���Xֶß�rH�%4�����R�Hv�ػ7�^�G��gO4���cv݋\�G����XG9�\�mxx۪�z��9�8�JL�1F룠˩�-sT�D�]�����z�����{��������KZ��q�(狨��r����ٴ���q�ӹ޻<���(�z(ۉ&�rG�>�Zܷs@�,����נ�d�X�F�_��ZܭB�#޾:���\�Kg���X7�rf��YM���@�}�@���h��b��6@rG{ވ���ԀާҀ�P��v� �g_��#ǂfI#�9_j�>廚ye4.v����gs��R)�0�H��m��յ��30N�C0�#���nӮ9�F��'�E�Q!��s����v�Nk���}!�O� G;���&�,�7\�@o�/mu<Of'�k1}�z*���j[���o�箤���Ѩ��m%��I�}�@�}�@���h��>�JU�<�6পn��Pt{�;��P���؀�j�m�~�ıȰ_��Zܷa���\|ξ�:�(�6'\T��t��v�1��pEɚ#%��'E�<nz��-�ݨ�)�.�Jv^3]��q�9���\�>�� 7[^������8h\�{���-���w�S@-X���G��"�G�>�9۩&���jo�G� F�Q�=��}4�>Vנ\B���QF�_��(�� 7]����C�� C9��(Т��!8h��;]�@�Wj�;l����lClmLX�nz�ї�qZ�+��*��kƛ��ԉ�<����(D��sa$4�j�9�ڴ�)�w�S@��)VD�(ۉ'7Uw(�M��{�#��| 5ӫ@-��?%�Ȱ_�nE�v�M��h�ՠw:�Z�ޟ�W$Dm`�'$4[w4�j�;�v���fW�Pt W�Q]�y��'{ۿ�)�<Q�n8h�ՠ{���,���_zx�9m��>�S#���K.Hx�3ۭ��N�>�\Zf�ڲ���� V�e�v.��	�X���(<0��-��j�;l���e4�j���"���Q���Zm��9l����Zs�ՠNgr�4(��#HN-�@k����ܠ5�b�nbQr�J9�����;]�@�uڴ�)�r۹�^Ԕ)ȣn$��ȴ��r��D{Ϲq����@:�ddA� ���^ىs�[��r��Hr�
�v�_�n~���h�����<�<b�Q�;z��P���'���+4�oM<;�I	�n+�p�ZA������F�-���-;�:�Pw�5g��t�8齹f�f���x�\���8,c۫������-����odj��8L�52�r����i��\l�xm�½k���b秓-k/ �v�n9�p�a�Ex�q�g9̛�
�Z�]��1���/�tB�m�&���X�hQsOjqt��6���nǍ�M������X/�7"��4[)�v�V���h:��+�X�7$4[)�v�V���h�S@�,�LSx�d�p�;]�@�uڴ�)�r�M ��h��#x&a$Zs�ՠv�M��h�ՠs��H��_�qh�S@��� �����\��ؚwU;��/5q��޻*��4�e��7Vh�C	s����Y��I��i[}��?n؀�M�!�sޏ{�����-�"6��cl$����[�߸�?g�E�a�0�V!���h���ϝ��/l����M���Yȣn$��ȴev���h��;]�@;ޫ)�/�E��cr-�� 1ֹ@k����ܠN��wS"6��nHh�ՠv�V���h�/ՙضw���R�Hԕ(��m�f/,\u#���]�+ruۣ[�U�� 4��b�l��R/��~��;�v���h�ՠ׍\do�"$���ܠv�:nPt�_t����F$�!{����r
/�ȴ�O;�v�p�Q*w�$`�T�#EthR��b3(�00p:L)E�6�U�7!!&[� Eep�+�b��D#r¬�B�C"L		���)2,�)�e�jA���`߰8	�)�A��p%D��k;`�����z%n2�)	R����4��"S�1�B;�1��d08N�y���8�A�7�2!H�FG
�`�;B!æ�H��,�BE�0�0%XL��۬���WFdX�L�jm@&�]� ԗ!	D���`������E�r�n����Ϟ ��d��G���>� zG!�`�C@.�_@�D�訉��
pڨAP�pAO�U_c��.��ǽu �w�QF�#��'~������9�޽�rs�A�I{3����7�y����6�H�@o��z���%���? ���� �S�us6]w]+�`�����t;�vzzn�K�;B����]���7�w{�ݾ���蕀Ih�`����l@n�gG�=�Wt�-���~K���ȴ�)����o�����@�Wj�f${nb�k!26��nHh�x�;]�O%�����}��@��&)�<Q��rG~W�޺�p�=�';��jL����
�AZ����?����~��Oܿ�,'�J�`��k��'8��/b��}��﯍��� ��n��2�6�sW��n���3�u���3��wn�t]����A	wm��}��?k�nAE�� ���?����k�{?g�;�w�@3�hxQ�D��jBj��.�{�#���S�@o��5���Y�C���z+#n�	�h�����mvw�G�,ŉ�w����oM͇/�*쒷#�Z��Y��'���P�� v���%��J}�q��֚`�������,X��}�����������6�6��Z�+x)9wW`�inV��ơz��hF �+����>�d�``\�n%�y�M�a�箅�u��iNv)8��=mAtm)�l��2tғs�K�������ȱaY��mu#��`�HS���z�n/i0��n=�k�n����Ѽ<F��狪�3���β�������.�����[u�N았N���kc6�U�SZ�p�[���3���76Kq� �JSe�ޣ.#���ջ�\��g#+t2�6�J��	闧������������k�9yf�����������H>�P�{ݿ�)�5�	�4�j�${<��q�������l;����Y���k�]���|�&�䗔�����Oy����Q�I-�W�Z�|��i���[� ����l8�l�֥���hs����%����_�{<��u[^���%8���%��\��m\)//]��$�a��v���;�l;����n%�H�6��FH�_|��\�����9<��/�=��=���|�qWd��rנ8�Nq���%�~�~Y���|"k�럷�I>�;�';����?��IHw���.U�'0VZ�_��9��=u,��9�޽��޽���,j�Y$QI-��ř�������^���7Ǡ�bK��{4;��T⍑�����@�v���?{=/��W��h�7Ǡ=�-�g~L�6�q��M�-�cuԈ�Eĭ�r88n�v7Gd6�\n�M�fb��(�k-��n�����=��rh���Աg�9�޽�Y�oʶz��8��_�q������M��9נ9�޽��o�]�I6�|�AѨ��#I���;�v�V��/߿/�0��
�(� c��㧂�Q5��ǹu$��}�I>������6�v���$��޽��ν�mz���^�|h�IO,��Q�u75w(�Z���C�\|޾�xhf$�w��#v�2ƣ�e�#�.�Sq��v+p2V�N���9��bz݇�c��t%��	����#qpO�@�,���g������zh�)Ɵlj�Y$QGm4�ܼ5��X�C���8���@o��5Ԓ�M��oES��Y+c��M ���c�r���z"e�_���9�E�e�m�MVf'��]�RN���ԓ��{5'R
�R���Δh�� �����2����m����Q���%p�Ƌn����mq���@f;w(gwSm>t�	��cg�e5xfny�FMT�普���7�\���6���{��>���58�i	àO��;l���Yb�K>a�����z5��#n�����/,Ėy,X��9���}=�7���Vf$��{���U�l���u�M�����Nq���bŊN��ƀ�|h�w���,hxZ�I$�;{נ9�^�|���b�,Ē���z˽(�X�*�ȢnZ����@y{���x�9����9Ǡfg7�����l�5����Bg���T�6���1�[7���[�����]v�s����F-�z�3ר�5��m<�]n�76����iI�"M��`9m��N���;��Q��ڗ��V1����v�U��3vvJ� Ĺ�ob�+m��9j�{4��2M��6�k���#v��S��E:˵R���4��Wd�]�Ę����w���*�K��q���q.2=A� @��n�n��������j8۬�릻�x��]�g{[����iH��ϻ�g��uɴ�Ą�O9e�@�v�fg�-�ƀ{�xч�H�3"JH�s����=!�Oy���ƀ�9xk���Tl���"��-���@�{)�����w���@�
���(�q�����5�=�z����+�u'���h��,ZD��q�8�v�M�yu��>��@n� ��]4�%��N���G<V�H�4S�9�mCn�ێ�o)m�}X��L�R�
CG�m��}r��M�wm�H>��@6�O:�RƇ�%�@o��z�f�f4��p��f��d@�ʂ"i !��*��C�57�٩'=�z��-����L���Bdi�x�� w�]7(�L�����wJq̤���#"I�4=��b����;�^נ7��=qff'�s]4��(�w,`��%$Z9e�@�g���/����<h�S@�q���'�b���"s����S:��m�WNY�:M2�&;�ٻ\ݼ�����8�f�4����E����ﯼ�v�J[�~���">�z�P0t�ꅒ��k�נ?~��ג�bJC���;÷ƀ�'8�Չ���F����۱�J�z���7����fby��@�LQi��T?���~�u!���^Ԕ�	�M�mE$4=��Ѯ��Pmk�/�p��w��P0��~�h�ՠ{9e���OxvS@��ܸ<X�x�D2��ݼ"]\wb��e��4��g���s\-�N,�{���65�%����NE���h�1�m���H>��@k�.&��.譹#��󗆽䔇xv�������s|z�bl;����n5[r�@sg/M�Nq����^Y&�;�;�_�cH�wҍLM`If~W��Z�㾺�s��I�HA덄���|&%Vfu$���1~׍w����3��J7-,����7Ǡ<�K<�������zk�h����5�Ŋ�ms�[���qZ�+�!W'W/]u��:�u�ϫ!�6����۱�J����Zp�b]7=��Hc�Ҁ��3gV�H�r:�@o��]Y��9�ޔ:}(m�]�{�����E�M�V4؀������no�GVb��;��h��4�z~v5�"6�<iȴ<�X��3�u�=�{�Z��%�Y�N�^����S����$v��s�Z�1b�$�ÿx�}=�>��.��s����h�3�0�bI�
]��8���7�api�>���1��MCn�� h$�Eb�VD��N�6�4|�~z��B2E�hK�!)�0��D�>�a���f�%�P&���f2e��\�� ���j8��5��o��� /[e�IӡP�U�Ag�:]��
�Z�֥�f]�QW+���gDf�i���{0��I�f�K�xSm� b��=���
�v��@l�L��T��;�`g�$�q-���6�Cf;[�Nm�ݝ"Z����14�$H��t���Z��P\ ��ghF�]��-R�J�9	�ayӵ��Zn[�BD��.v�Qv׶�^S0�X�Z�����X^��ࠔ#ٺ��

bnѺ�Vض���&�ϲ��5���E��
��j�C�[�՛.�O`���ڗ(�=��n��`.��J��Pgr�������T�Gf!O�ql`����=��p����N{h�;�#��Yb-�� �Q�',�0J�,B�T��a�f�,+f�km�a.��xq��..�Gɵs��X�0®���q�p�<AѰ6ڗ(�t5�[M`ۭՙ�͸ъ�n�V� �Qۢ���֢n���f�D8���@+�;@�e`�f�
{W�j�4R9�l2�g��v�u�=f��p� �յUU��m)�]�G 1��ۯ�-V�լ�����U�����a\��*NB��1�-�s5R���t���3���v���$&��=���(�a۱mmS�ɻm4\[��6 ez�'�2����
;#\g��ֲb�ZTp�q���i�˔�:�n����b-l1����c�b�[�V��B�$�ȍē�;d�gZ��2��{lZjXÎ۴�$������>�,�7��M� ��$���[�JN�D��@��v�<q�l&��voa�k&��vs��aF�z�iuMUX�i��lTb���G'"��J�N�M�a��ٔ�����(h�j�v�C�l9KgUQ��^�JV�V�E�������rc�^Z9�r�H���Wc!��O�ۋ��6]�v�@]���k�Wdj FC��s]A� �A��oSea�NYa�P�&iZ��$nDք�����q�+�A�&�4a �ЉƟ@q�*�:�:��piQ^"`�'�QW 3�K��5��P��!�ۯN���
T���FA������!=��]�2�
�*�d�k����z�����<Z��غ^v���v�*=�v
�8�[E�"\��a}Y1�8�smV5 㧆��#�q2�<�m��v-�盥�'F����`��s�����Ӝ�C����$��ȵ��Xu��	�^�$��v�[������
A����E�
�#2�F�����{����q��w��u��s�&���{u�6�3�.,�8�J�u���i�v.��k�c�pv���;��8�� 5�r��k\�D} ��B��l�'BH�u�Am4�9ǯ�y)�w�@w������w����9ؙ����s$x�"�9]��;m��߳��x�/���mX��#i(�cȪ�z#����@=���M���ӎ_RIz�%��O#m��j(�}�Iw��-I%���?f_o��Ē�s�Ԓ]������0�M�&���تu�ˆ�u�:��e4��.��f�2��p��;��r�����c�bF �K�W��_|�\�Z�K|�>^ř�Ė�[}�o��m��ޙ=cV��"�9k�����x=\Qf��f$�R ��A"���B @`03T��p<���_}��Iv�<֤�흫｟��m+�&)�FD4ԂԒW��g�$�zIRԽ��6�����s�ԒJ�֒����fD�s>�%���7|�������K�r�[~�췾ﶾ���l�'�H�u�A$KRIv�տ$��gn��$������%ގQjI%�w�&���1#��n�� 04cva�ԉv�p����������F�������$�l�KRIv�������^�3<�Z��|�����枊�6��Lo#q-I%���}��fcmZ��4�o��������x޽�X���w���2c��j$�$���%�RIv�ս�=P�� E_
'��>�yn������ose���&�Q��  �s�~������[�m�w�ٽ���ř�e�\������vƭe��)��$��Q$�����r���K؝�z�K��O�I+��+����c�1�����=��o,\u"�D-,lq[���ַ�	��{����hU;BB�VI���o}�~_|�|I���$�۴�����4���KRI/U�D��m�V�m�)7�5Ԓ�#|�u��o����m���>_}ՙ�G��g �͵�g�oRI[����%z�KS�X���{�����s�sM����⅒��K$v�|��f)�k]oM�������[��q�[<$F�uV�T�* ig��y�DO���sg�6ߧ<֢�,��RRJ=6���s��ͷ�Y�g���I���{�x��ڽr�RIZ.$�"��@��,n;8��B|�g�U��8��v�ul���[����{��@}����H����0~p�?���\5�m�v�}�Y�������/�m�vt�H�)bi�
Id�m������^X�b��v_M���{��ͷ�&�&��bII{������F�R�O�m��^�M��s��}��%�)'T��m��w]>���9x*��!l+$�����̓}�/�m��9�4�o{�}�o��N���m��>��'p�+nJ������#�m�$�Y��߼om�������s�/�m���"��F*�{ώ��ZH�sش��jqw��۳|��\��v�V���&NbiP���@"��wW2���q�)�H�.�tq�$���.��\<h\�m��yg'\�)qw1�����uʮV�F:�c��ײ�mҖ����4������ρ�nt��>��mʫC����>֜��NU����>v@mcn��+�w-;����kK8j7.pg8��1�8A��.�K���2k������v�7-�犷5� f�nv�M���S)����|���Fw����������$��Z�K�߳�'9^�g�Ԓ_z.y��NB6ԇ�$��Z�K�߳�J��jI.��>��j�u���,�vJ���zm����/�m�'�ZԒ]��}�I^�E�$�ږ��<���M�9�|���K�kRI[����%z��������tz~ �$!G,zm���\>����{�����~���}�I\}��I%�w)���$ll�cyk�"�4v�ӛ�N2��h��quGU������{�8:/�F�DF�7�I�I.�7I%m�g�$�q�ZԒVݧ�$����@l��Gh��o��>_}�̏4jffs�.�Sw����޸}�mF��$�I}��m�w²IW�6���zm��s\>��I���m����/�m�M�1��Hݎ�]��䔝�~��ͷ���m��s�/�m�K׫^���߻A����M��R|�]�n�J�~ϾI.㲵�$��O�I.:��P��;:���`��;me����N*�M��@�7�q�藥;u�G@iLKr�]�@���K��ũ$��O�I.�7I%��iH�H�Q&�9�|�]e�-����[[���|�}�����|�9������G�M�b�NE�$��O�I.���5lFP�,X"T� �X� ~��s��6ov��N�ٺ�������5k,�K->��ԧ;�|�6��{ߗ�6�������,Rw����6��������6D170ԒV��}�I{[�u��m���]>����]#M������w�mA� 9b��5P��t�.y�ͳҥ�y7��ƎN��ݷn��I�{Nàm��K���Z�J۴���l�?��b�F�{������:X�'Q#v:�*;k�m�s����Y���F�m�����o�9y^��g�3[[�h3�#�%��#�����}tm��s�/�}X�%$�;z]6��{��|�{|�OU�Y�Ihi�ԳI�����6������9�vov݂��
�D
.��ԳRI/��m��´��#����3�K���RI[v�|�]����w4������4�S6���������z�]��d�9\��5�;q�7Z�}v;��w�	=DP��4[�{�ƀ��sK@[n�g�� �=}4ܫ��k$DmeTUU\�5�P�#�2v�(@99�����嘗�$�{�N�HY
�I.���#�h��G�y��@>|� s�dd2X�J��Y���;P���5�P�xڄ�6����v:�ev��������o��|w�hԓ���Ƥ�Edb���v�����e��<ñP;�����v���t�G���/l/:v�-!b.QOWT�[s���9_j\�玵�WT{���8y�t�$%Χli8�������F�8��*s���;VWb�n��7�4|OJ�>sr�uJ��Y�ӿ�~�x^6�\��{q���qI�2�,ؔ�r8�7)Qq�e�L�+���n(W�K�i��@��q�zC��������õ�jfD��+������[��w���5�OKaZ���n��� ��)������O����� ��F�6�&h��o�~�ĎmN��bX��=��=��Z�X�l�9��Y�j$��I�;��Z��Zfc{�;��;��K@o{|z��'%i�1ur��<���7_(@<mB���%7ůy��]y=cV��ԊI+��Z�DGow���]Ҁ{Z����v���.�s�q��p�=tф9{[�<�R���t�n�'j�o\�e��8ZP��"����=�Cu�޾Bw%�+$�h�)�=q`�&ME:EB��*~@���c���y�-��斺�cg_NF9:���B
��y9נ?~�4�{^ıI�{�Z|S�z�\7�<�Q9%�B��f���@dN7H;��z'���W��� ��F�rL�/-��=����������3P�n�i������rt�t�9⵪L���l�6��fێ��s�ݮ}8��w{ܶ>��z� ����|��]�ֹ@n�Q��D}!����-��^E���,X�7$�/_j@nkP�xڄ�7v�~�{�T�ӓ�5k,�H����w�Z���-]4˹��Rw�f8��t\�H���Pp?Pv hEҡ��C2\0� ���1"@�$ ��[cT�C{R�sOV��F�ɗ"?e�15�G� �M<U�	�"��A�b@�кH|E 7l��%P�D$J�Ga�? ��P¦,iU�|�hk�d�6?U%��,3X�`������0��P��Ԩ�A��|5>:�a�A~�"�l��@����S`�S�:�hDz�p� 	Tؠ�DL�����r�t)P�;��s9ԓ��}u$����Lf�B�[p�U��,X�w�����t�h�n�Z���q�&D6�8�����}��_(@=mB����Ee��'S�UFT�	�5uJI3�bMr�e:\Lx��V���}�����fҍD3$rN������s@��s��Ŀ@��n��^;�<�Q9%�B����B�j8���7+��$Uڱx�#hQȓrI�����u��-��,K�fI��y������Yȣn$���4=�?g�_}�4W�]I9�;�Rd8�"+*�;�w��;ʮjȰ17�F��h�{�_}ϹBg�@~�E=ߝ��2g��G�����;��뉊k[��ڱ/`o<�V
ޮֿ�������?I�iN^j�� �ߔ ������{���߼���<O�6FɈcnf�{n恳�ݠ�r��֡w����*!;���J���t79ǣ��31+�����]:Л�6�j!��m�y{1bS�׼�y�ihow����h,�h��1���"�;ε�G�9���9���nP��bIfē���:Ӎ�7��+J�h�%�I,����S���aT��4\u&��.��:{S�zkf�-).���v���b.��xv��G�ͣVz��-%��s��t9�B���Lh�l��S#����x�;lݱ�IU��=F.9���u�º�Q��w9���9-��Xv�hks�s�k�x� �um�ĢfRqc6'VĜ�s���h����M��F?������f1��ĸ�.s�v������W+�����'7jGR��u������Y�AB�D��L����4�[&��;V��v�h�%*ȞEq$UUU����w�=2=��@o>P�ǻ�]ēf�ޭZ&���i�Kn���z��o�Z?�3��9������ �ί�ƲD(�or-����9{)�ur�4=�^�yh=Lx��lQ�QUW{l@w�V�W�=��@c۹�r���~qL��$�ɍӪ,\IW�������i�r7g�և<��=���n���t�ܦ��Z����<hT�	�`�Q��d�I�w����"":D\�  �ELQ����l@l�wh�4�T��ȴ�$Zy۹�r�S@��h�h�]�r$ܒf�عe,�n��ZX�j���͌���q$6ۆ���d�;�j�;����7xh,��݅�o�
U,�����uqW�q�g�9Xc�Qo;fl=����w<���#Ǒ�#rO��~��;������W-�@/3�󱬑
3mȴ�j�؀�����ܯ�2�ǉ�b�Q��Ĝ���Ɓ��d�L]cXXT��Qڠ�t"%}���{�RNs�ѩ$�Q����L��!�ur�4�ڴ�sCػ�4*V�߰m(�EwWv�ܦ���z����| 6r�4	L�U�f641LrO��>݋�\2�������ܝd���[�ׯd��Օ�Gi�$��>�n���M���������- �U~�mDӑ&仄=�.�{ޙ����f��IB�<�6�Hm����h�ܣ��DL�P��w�5�U�C�+�Ym��KO�����;�RM���jLx
�so��s�$�ˏ',j�;"�Z��o�Z��,Y��||]��@�j�>��Uڍ��i�b{4�'Y�xGn5�5�ic+r]����H��o�,KԹ�I�;LMʾ������wh��?���}!��B Bw%�+Q�h����fb�$�R��;�-��^�ybĒ��������fI$����@�;w4�e4�vɠ÷��8cnI"K����D���| 6s]��1{̜����xl,���U�e� >�l@l滴ek�f��W�(�
��t������8�7��E�:��
���U�z���gon��9;N��`�jP�d���M�����x�o3n��X��y�"��y�-׊�҃6�u��S)���]��^֝�X��
ĸ��X�mkcj^��L�\ƹ���}��aw<X9�x�Bʆ���B��R2Y�E-���*�tހ�R]�$��Ԗ�h6��9�b�2�*���U w���{�����s�b&�(C��7�q�qm^K�Ұ�C���X�m�i.5�����j����V9[~m�s����Z���B�v�kh��@�QX���m��M���g�2C�ﴴ���@m��-�s1��ï'lj�:�UUw(��c� 6s]�2�z �|Ȝ�N���bnU��ǽ�]4��t�Ӝzfbļ��;��@�����2,jC@��l�8�Z9۹�s�S@���
W�IX!-��w'��VdS��-I��f�m:p�$IRzK!mz�~}�����Q��$��Z�����v�h�r���ė���w��g�G��E.3����7RO��tkH�@:�������Kn��M�艐�.��NdN7&h留�vɠs�ՠs����IJ�'�F�I��8h=�bKاo;�t9=�?~�4�I{'9�hw�Z��	�+�Ym��Sr����k��7z�@9�wh��w���}��K�I��=h�r��x붪�g-�`��W����>�?�p=���:�\努����|�����v�̦� [Տw��LF$�h��bE�}v�ݮ�@fkP�"&C�YQEw������*���8�Z�~3���F�
�J�@p�(TR��4})�Uӭ	�	�E̒Iw����G��������؃����h)�O��8cNH�Šs��������9��h�nP9$˗%͞�7cv'8�vڸf������k�]qr��q��4�;E�;����;JJ7"Mw�޾9���Z��G�����_$��D�Fډ1�8h\�}�=��꡺��P���l_�2k|+��NX���m���^���|����X�ؤ�=|hvw�h�y9cV��	�נ�{�{�����@~��$�<�H#��"�U�9������/�I��= s�2)'�v:���h�r��X�Y���?�N��廚3��]hk��r<� ˷���
�� ���G����Ǝ�i��O�g���<j(F�s����}�@�-��|����yR�&�	���I@fV�_��꡿ߔ 5���6��/Ж68u9��QG-�2�����h�e4�Ļ]�zz}W]�mFԃMG&h~\�Ɓ���9�ڴ<��}��@w�mӥq[$tq�9M�Z���P��@}�؀~��/���1��T�UМ��e�V6 ���A�`�\�h����Q���^�6��:I�G%!h~G��7��i,'�H�a� 8F�"0('�I��0��"A ��!(C+�Z�dR{��>�쨟:z$b@�3�29�4�sa_�" 1�HF� %4^�IP��/694pg/ƪ�).^�
B �dc��}$j9\Kx�#�
a��[��'-��kvȐl �m�d����T�`Sv�2���6-��,���a@��d�v��t��b�iT
yvB�9�jT�;� c��<˛m��,�Oc�
5*˳0WZ��U[��7V�n�箩Bg-}��q�h.�Q=�P$��.54<"u��[pm@�5T��-Ւ-f�l�JaUa�6��tL�xX��n��c���
�duXс��]Y�h�Kx����4� �.)\�Ժ�r��=�g��m�չ�l�J�I��[��r0��K�V����Τ T�t�c�=+Ӑ����|aR'(��lX��y�j� @s�s����׵,����0+�)�U&��Vȼ���q�&J�.GV���n��4b��]m=t��5 �q�+�$uք6J������H��pn�`}�&@����\:a��
�Գ���<�:up, �X�p�Pu2�E�@���P6�9<@1n.ж�q��B����Gd��=6�l�e���2#�y9�V:��,��ewk�	ے���Z�b�ZW����U�2콊���գ��Ŏ	w�]��z7&Z�ܝH
��U�H-TT n�a)[<n�(�sp������v��`�Dbm$�fH���=��݇t�Э��,j�풑ukx*m�Ѯѭ��9�9'��x2C1%�5	��#��WklZd%�q��*�m�����۰��t�F��d�n��p2Cb-�ݽO�pmŶw(���l���tutIE�a�(5EW*�UH9���ۄ�3uy<�ghKd���Oe3��%�1e���2�Î�7ln�W�1Yh����S�ɇ�U�펪�hM�I��U4���avĴ�R��m�`�$:uT�:��Q�iѵ�r�E�CƖ@zѲ�Q��/5�vx7��ŕ�d3�q ���kʋk��x���B����mG6�e���6Ќ�a�x���HLsgF��h�Ӭ9��l����=������d�nl��m�D@Η*�8�M`rB=E:�0��8	@ٴ�p�DH �:�+D���N*��A�̕��?���:��ƹU��X�ݪخ�Z�*ʘX�9�c��T ����*�`�s����;J^�=.�"V��NH����0�:㍩��Ki�<�l��@�u��nݞN�2�k%�-��l�Ξ����\k�	݈8��vq�K7�GIu��F�'H��3�5rr���mY�j�<bKh�
Uw$m;n�u˴�P���y���3V��3^�k5?����{���~��d�6Rƚ������b�%]9��S��i�-���+(��2���b��(	�+�Swu\mwJ1���?G興���I��������H�����9�@f�b6�� 2u�_������dRO'h�u17*�﯍�s|�@qvנs��h����	5#�w���U 6_u 3P��ӯ��+Bo��#�#z��ĒIo}���9�ޚ���&����{��v�]����������I�õ�6En���-��7�;8�����G�>��vN�Yu�7���l@fֺ����{�=�H�U��R5��v�M�̂}^�B��V?��R'���ڄ�RP�O$m�&�7�}��V�GD��r����pX4T]A$T��Rޗ]�H���l@f�kz�J�;��1�M��r���즁ξ��+k�>�~eUL���vK#�-��s�㞖!2o}�t(t��xx9���6�)��I��;�)�fֺ�Kn�ޏ�7{� ;i�Wz��㬄�����&��16m�{�w4v�ht�Bn�lP�b$������}�{�R�� ���&��Y��ξ���"�F)�E�8�% 3P��v�mk�A��D�>�@��AQ� �Qɚ;e4u���qvנs��h���I�Bx�'k��'"�x�j�SU��ۛf�=vog��9�۞}XD
:�K�m����?��~����1��l@f�
��&�ebdv�4�rk�6o}�;zh��o@>�W�cY"#�5zcj�؎�G��t����� >_�w��LF$�h{?.�o���c�}y��Rs���HDpb�b�`-L�s����{��}5�t��#�h��4u���qvנ}m��9�)�\�J�dM���b��[s��Ƹq[fi�jW�2�.<i�sX�	���sС�I�8�k�>��h��;]���X\��1��m�٠>�9���fcg9��Gؓ|����:��= ���$�NcN)& 7]����@d���mB�̺p�+d��8G)�������M���@|�P��v��q5
$����"nn���ۤ{���G�7��y9�4��9�	`%��mk�q��x�lU�굥�φ�T�W)�����g.���u������v�B�6�,Ńjݍ�h�W<!��㫭�^�݁���m����ڜ�Xծ���:_C�96�!�8�
��u�7��
�N���B\:�{:��=u��+m��¡D9kh
�z������-ƺ�M6N^�.�u^�v�%]��`町���nN�a�[�Ͻ��=�{|G�vx�d���G��p��x2�q��j��.�����y&ekz�]Y<�k$B���#�9m��;�)�v�[�8��@//獻�AF�nf���t�R%�H�jD{�'k����G��8h��o@ⶽ9��\�d���À�pm$4`6���+vPn��l@k��1�ar�&69$�9"�>��h��;]���hK�6�<0N6�Enްs���Dta���i�]0�� ��k�\]d\ڌR	������+�o@�]�@���h�%
D�m�������'���cZT����js�֮��w�s@�l��#���<�3$��B�)vR]wJ�mB5��l��J�7F�D(�������}�@���4.Z=�v� ���w��O�L��5�8�H�nPcj;Ln�3#���%���Lf,#��b4��]M��m��;tیe�k��N|^��kg7V 2q���ܠ>�� 3]���Zw�QF1H��uڷؑ���Z|��??��5�ٷ����*���\������Z��xh�%��$bV �"�*)A��W8& �1��D*#�?�o�[�@�}�@>���mFӌ���������g_�ͦ��D����RP����&ƚp�8��R�G��t��_�l@8�"����k��7^t�7o6'�\[g���e�k�n����x�䁻�L<��n��F"*���ܠ3����G�:�� �<�7ᬑ
1�q��r�h��8��=�v��~��{���AH(��������Nk)�M��v�����D��8h\�z:�Z�o��R:a!�@�q�;�M�V�����Q�R8=�v��z3yq���@d�e mӸ�*S�a�۱�I�.˶0V��w`fk7Z�k'N�iX�=u��a�׵˒�X������ 3]����@}�l@�d�3Q��q�hs��;G�}��h��g���"r6�D��g_��6؀�v�ٶ�kp��d�<�QE$��.v����>���A�ı$�7Γ@�{2�F��袠��c� :#٭q�:�+RM���jI"��(x�)SD��3Ʒ��Պ4JԬej��$�k����"E�۝��BWd^Gd+p����>ME�%�G�g�w��6�Փa-{\�����b֭ۄ�vS!v�'ggA��ӢHkbi7';L)��M�I!&��1=F]�n�8E竹;b�$���Ғƹ���l� �l�=�lk�����J�+Jiy�֓�i:�!�nF6���:���l���f$���K�~��dv[ET�Iru����m6r͕D��ӣ���N�|��bAF�!)��M����9�j�9�)�^:?����M�ㆁ��r�DG�Mu�(޾�؀�Lu$�0m%cR9�@�]�@�,����M����8��/�cc�H�E�&�_}| 2q��ٶ� �����q���4��M������M�YM�ēʆ��҃,cc\�9Up������]-������&1B9k"M���@��n=�m����m��eER�"�
��sss��ԓs=��+�2C�SBD\E������l���L����#�0�c�����}��h\�z�즀^_����1	H >Ͷ 2sYH�nP�؀yL��_�c��8�qs�z�v�y|�_�l@w�t��}�\ܖL;]�nO[q���9̛���t�b3��Id�z��lm�B�1��	�/����9�� 3]���#�u�h�ꠘ�\\�I#�)��[��s�S@9��{���Z��J&�bq�ܒf���b ��Z3ޏ�}�<DؔF�����i�&�$@��H�1X�bP�WHi$��� $B�$0Bq���D�*�!��Z>����$a"g;�dc$�@�HP��"M�bJ��~
$���Hc�)f���!5G(�M���&�*H��B��0f�T�q���ɾ&L������H�*B!�`�q*qS��eP�W��0��BBHF*M��P4�"���� 0R�'��
e1�0*�*!�@��� �<�~��(J	��D�#�b���֮���{�P/
�H����'��8h{�g��� 5�t�3P��v�n��V]`�$�9!4uڴs�s@�l��s���/nF�����5�8b���r��y�TK�H�8{`.��^�#`�`} lS�rd�M!�Šs��h��s��:�Z���+)bI9�;m��������@}��@k�Ey_�c����4��ɠ}��hܶhs�����70M
(�s&��m� }����b��(���DA$
Rv�A�@Cb�}�>&�W:�,��"��8�r٠}�l@���f��h\����@��v;pN4�;v��S6ڑr��tM��[�N�E����Œ9�������@���f��ݠsnb���YccI�@��n=�vS@>�9t߷xk�$�7�t"�X��n�7W��w� ��ٶ�Nk�@��k$"i$4�[4���Nk�Aމ�k��ި��ɻ&8�rhs���=e����@���Τ�0pQ�\X`V���Պw����~������RX-���Ӄa�J�	حuFĞ��p��<�d	e]��yz�y�������5&�:�kۡ5��;� �2�7Ͱ���Yݰ��4�E:mD��,�c;Q/kɛ�h�똶�f��t8�lFk95ղm�t�Dݔ�e��53�r;%�=Zs��mc�T{<�gsm�e`�LI�9��f�\����5`��Ca+nx�{�^�=��J�5>�#B�U�V�Fb�4�ˣ�c0:�;�����������O�n|^�q?���}����;)��ٙ���4���L��!�`���f�cv��6؀ݭwK��{��z*|�ג��[#��� �=�>���G�33}��l��w�@7�!���,n+m��������ݝ���v� ����T)���'��%)�9��Y�=��g��\��������l��Wz�Ҋ8�5)#'�Y:6x���S9��S����/Jm������;=[l�	�I`���h9l�9�)�1|�o|�4���#R������M���Zr�� �P��@��}3�����������f���۰D�8�Mɠ}��h\�&�����@�{t�8)��Z�̪ub'5���6؀3��Nk\ /��452&����I�}��h�ӻ���Nk)�"�fu�k�c=��'�8ٕ�õ�6If��b��m٭2A���LɑF�p���Z��b'5��{��| tL��Ɠ�$��즁����s���[7��#��Y���'��$�ԓ���Ƥ������
)��Qh�T") P"���}��:�s�S@�{A��24'�%�I��Ś�w��f���� n7^��0��<��r٠��9۾>��7�}��h\?2��6��m����n���n]��&䊳�]�P�I�5�&�oL���O6��b��>��ƀs��hs���-�k�?���O��;�=sh�m��n�f��u�Ʋ&���q��>�e4
�����M ��M ��`��L�r74UՈ9��f�z��g�
#"�>Z��!��U@��𨒋$�v�F�6w�:G\��˻�۶� ޹��7(9��X����T�&HH"�E�u��������睒T(����Z�VI�ҧCʒMY�s��7(9��ݱoh�=���D�H�S@�]�@������sk=U}>�&�h���]�z:�@��S@�]�@//�݂&A��7���M o\�6����_R�����\�\��ㆀ[ڦ�λV�W;^���٩ �����, �,������CP�NT�1 :�F'�Y�Tm���N7f���;	*/F��v]y2'I��t�ڀm�oUO��<����m��=��]`INP�Fl��N4���nv��lY; ��ݭ�Z��8��L�jy��`�`�Ɛt������0=�6���]�t�Mў���6�8؂�%��do�pb��'ZΤ�5�kq{�<���{���n-?�>n����Z�:z�u1[4�#Ge�1�_f����_���,)���ȧ ���@���@�l��[ڦ���@Ys&D9m8�Z\�z;g s���ۼ5噉%��}�1Ѣ4�i49����h�j�f~Ĺ�<hV���*Ȝ���<m�'sY������o�ǽ�h�n��/(����O"#�M�vS@s���m� =�6���G��=s���lu���m�lx2�q�\�j��z�6���]�O�7ix�V�lt�Ԁ�6؀�@}�l@���eT�X�\�@}�w��Y�X�ĪQ�o���| �@k�Ez_�d�q�@/{T�>�e4��ߒ��@�l�uS�8�6�H��M�M�x�}呂���ً1�n����@YL�i�F�4�j�?������y�;�>���@y�u��q8�;��iݻ�51X��g�vk�W'R�+;�� �ֻ^L]9��,�B�8�m����4��M�vS@�}�@��c��m�������hs��k�Z�}�@�讨���O"#�M|�{5$�q��M�D�@w��+C�&Pr�0>�� ��]O|��������d�jTYQ݈u�Pmk������b |��v�i5$Z�}�@�V��|-�4�ڴ���8f)1̟�s��;Ő�}��V��\��/X0Q�M�b�g��3��'���c"�h{j��즁��W��9]��8��&�F��
7.m��~�DD���J>���޺�cg��T5ܪ2;k���hvs��ֹ@�͠>ݶ kpI6T��&4ƤZ�}�@;�T�>�e4/�ĳ�s�w���[��9d��䌒j� n�6��v؀�Z��ֹ@|��'x
<at�L�u����}���==�����7�ڛ9�]�j��8�-�ݩ�эwWsh�m�u�Pmk���� �;_�ı�#x��䆁��}/��r���hw���i�;S ��&��@���hyj�{���K��������F�?��@;���n��A���Je�H�1��Y#�F�S@����;]�Bo��n���w�:�!�,`SH�d2N�6u41`�,X��A"��2H�/��b�@� 	�K�h�0�P�Ѐ�b�R��%HԀBH	3ԉ`�*�D�V�p�(D��F|�A�B �b�	RU�T��m4H�IDB8�P�BLK� \,��9�e� ���p� �{��>�q��!�0�#I�?���SS1B!r��F�+a�"���lh=IX�`�P�(��Hc���h�##�dH�,#"1 ��As״�+�!0��K��a#��!���a$o>�����3�0��
<M�Θ,H�D H)
E�7�����aE�1�1#D�ȐX����Y���O�Z$� L��ŉ�����nϭ��im��PqUU��B�7R������ͣl��kqV��IekcqU֡d{V��vە�	�Eɔ%VW�u����%[�.nְ�H�{�����",f���4���Y��{K��ãR�U�r�!u*U�6�q��:�6�.ȥ[Kp	�e�X�S��l�Y҄#n�E �R�U�*�r�Sٮq�#⮐�|vޱm۶T�6 "�d��ֵ��gyyv�e�N�jnU&�0Θ����©Op'nU�=���r�0��';��p��<<���X�՛n`3��Ʊv�f7��:��>b�gBD������t�UP6��b���㍠6oc�q���@�����o=�������54ڧN�c�y���EH��6�ɵ5��m.2�t�l�UP�m�ɞ����[���A�-r�uq�v�� %^g�f�GJ�+7ST�A�#�Ym4��{��%��x.sa�d�x�$ܔvǛ�f��n8s����s�i�b�mcn�8�&"m	�]�n��Ź�E䜛�].kh;$��5�h֑�	2�	)����f=-]��d���ёi	�ei1D���kQ���΋d֚V�v����7�&4�E�rr�Id֢��"�q8�l]�5I}��v����{um����RҌ]�צ,��9�7��aU�q�y{n���ڵ��'�m꣨kj�[�X�4��s����݁�^g��b捓#��rup6t���Z�<v�A5d���\�u[A�,�^%� ��^u���Fƶ�s���v$$5Ҷ�im��
���D\�e���-�7���<��˔Cut[�����
Q�QA�R;���Se^�5�-��{����cE �����T�#�����nGͰ����u)-n��:��� I�v�K����n�veIC.�"pJ��k��=����#ˮ���k���Yf����{5�M�ЍףM3T��M�ؒT��H@צ{'^ܴF�͒�t�&~QёD��UL�� u*#�F%C���@�A"��D�6������ qA��
���Nn��*��S�0bE�Y��y��P�u��:�*�:wVi���7h�F(ܥj��BO\J���n׊I{eֶ�R�/]�d �[\s���d�͸fq�w�A�`^��\ӧ�{&��q�)�Ͷ���Վ(8�[<y�	on��z�ú�q�9�]m�F���v��6�\�vE���>JrW-�9�=S[V4���9�t5NV��ffm�V���=�������˓8��V��n������8��֧���vI�&O���#ɂ��cCREp���@}��P�s}�(7�����$Ph�)�%"�>��Z�ڦ��{)�v�ՠrԣ�mdM�!8�u��۶�~�G�_S�@c�Ҁ��]Q3	1��qȦ��{)�v�ՠ}�ڴý�M �;_�ı�#y1PU݈/] :"1����t���S@�g2缾q�mI$2d0Qō9������]6r͖��4{Oq�]5����ѹ���rL���;������}��K�}�f��gE;�B�*�v� =nmG�D���Q�wm�/] >��[����?4y�I,��r)�q�� �H��� x�������44�#C�Vנ}�ڴ�-���n����
�#IH�mk�����;��1�� �[�:Q(���"�3�D�L��Se�K�e%���n�]�u�����:�}�>~{2��&�	���{�@����*��3���h�x�3"���C�$���bηH��� {��2��$R�Ț���@u�����ٓ�~�0dʷ������I7��S�����y��s�N�;j#�٬_�K? �1�׿]&�X�%�t��:Mı,K��^�Mı,,Oc���/�L��L��ފ&w,��UB���7ı,K��t��bX�'��4��bX�'���Mı,K��u��&bf&b�����FA0l�GU����E9�S�;
Eݺ�"m�<v��@^:�y%�u��ldh�Em�/�L��V'��4��bX�'���Mı,K�羺��&"X�%�����7�f&b߼����FG-,d���񉘬K�ｍ&��H�&"X��}��7ı,K�����n%�bX�w���/�ę������zt��;a#n�Mı,K�羺Mı,K����&�X�%��{�M&�X�%��w���񉘙���ӯQ�%���I1��&�X�%�}��Γq,K���צ�q,K��;�cI��%��P
z����6+�L��}t��bY���ލt��E��6�b���&b�,O��zi7ı,Oc��4��bX�'��}t��bX�%�O{:Mı�{��������T<�NZ;\���u��![l�h�ա��)ּ�k�;�F1O�2+���k�&bf&b��{5��ı>�{��Kı/�{�І�X�%��{�M&�X�%�}��c�Dꣶ�;e��񉘙���r�X���LD�/��gI��%�bs����Kı=����nX�%��^�&w,��UB�^�|bf&bf'��t��bX�'��4��c������߱��Kı9����n%�bX���@]b��8�vȭ��񉘙��}���I��%�b{����Kı>�{��K���1�����n%������C^ʣ	-$d����bX��}�i7ı,?���I�Kı/��gI��%�b}���I��%�bi���J'�_ә��.�\/���]3���:��uF��&ݍ�$����WE���q�Su��{CW��5o[�T�u	�@Ö�.�֦�a�q�I��sQe@��T.�/7]��c՛lE>��3���m����t�wN/V7n�����u|�`�c�8���6]�;�V�Iyz�`zLj��Ge�=��������O[C�x�{l�;��T+�^�Zۿ�	����&6��c�J�.6ݵ9��+mH�k������o8�8��3�[�6�,��LS��~oq�������]&�X�%�}��Γq,K���צ��Kı=����n%�bY��:�BY$j�	#��b���L��_t����Kı>�u��Kı=����n%�bX�w=��n'�b�&&b��5��A�(�%�۬_��ı9�k��n%�bX��ﳤ�K�,O����7ı,K�O{:Mĳ13��ّ��Q\l���X�11,K��t��bX�'��}t��bX�%����&�X�!b}���I����L����I'q�GmD��u���bX�w=��n%�bX���t��bX�'��4��bX�%�{��7�L��^X�b��Z�� ���Hw7=ؤ�9��!�ky՘��ì�n�Gg٢��,��UB�_ؿ���������7ı,O��zi7ı,K����~b},K�Ͽ]&�X�%����My�:��i�"���&bf'��^�M�{ G�C�Þ����Ȗ%�7��7ı,N�>��n%�bX���t��bX�'�d���ZH�,��|bf&bf'�s�X�11,K�羺Mı�$LD�K��gI��%�bs����Kı/�=��pqW�X�1313�^u�7ı,K�{:Mı,K��^�Mı,K��t��bX�'}=u��I�BH�X�1313���gI��%�b����I��%�b^s�Γq,K���ﮓq,K��3??.C&aK:h�m�:C�S���T��˧8�(r�6ƻ�k��8�Rv�z�pg9�n%�bX�w���n%�bX��ﳤ�Kı>�{��Kı����&bf&b{[�b�mJ��f	��3I��%�b^w�Γpı>�{��Kı/�=��7ı��9���񉘙���tR9�*��$�sq��7ı,O����7ı,K�O{:Mı�e��"�"+��
�E0$��Ӣ�
>9������n%�bX����:Mı,��\��gr�X�T+���&bb�����bX�'��4��bX�%�{��7ı,O����7ĳ1ogt��u��ӭ�.�|bf&%��{�M&�X�%�y��:Mı,K�羺Mı,K�����bY���tEO�E���2�G��4��/5n]��̋L.f���$�[�tVNv��}]v;�\���FK)�_�L��L������&abX�w=��n%�bX�t����Kı>�u��Kı)�{%��6 ���u��131~��^�|!"%�H���e5�O���i	�>�9qh��13:u��\�H�rK�f�7ı,Nt﷤�Kı>�u��Kı/�����Kı>��^�|bf&bf-�]#��(܎�8Γq,K?�b�'=���Mı,K�߿gI��%�b}���I��%��3�q����o:Mı,K��cjTW"%��/�L��L��s�Γq,K���ﮓq,Kļ��gI��%�b}���I��%�bwѷ�/�O6��t������F�l��·�Z�f��N�:��;7��r��.�Wg6�9�n%�bX�w=��n%�bX��;��7ı,O��z�? O�b%13�}�_�����~�L�Y,2bf�7I��%�b^tﳤ�Kı>�}��Kı/�����Kı9���I��%�b{��!�\�n%.s�fg:Mı,K�g޺Mı,K��{:Mı,K��}t��bX�%�{=�&�X�%��=⒞rb���+%z�񉘙�I	C�=��Kı;����n%�bX����t��bX�'�Ͻt��bX�%>�`��:��Wv۬_�����{���n%�bX����t��bX�'�Ͻt��bX�%���t��bX�'�@�@�������ɜ����2�=�������� ո�휼���ڎy���졻 n�i�66�l��Ξٶ�J�S�@��Xh��b�lL�!��6+�r�Y�a*�v/F����-��Y����m-'p=;�7nmip�Z�=k����GF�S�HTm�%(y��f�9"<=;JԶu�^C]�Ci۳���h �:���z[�'�5z9��K׮���{��w���Q�e�ܜ��rv�������E�u�Ғvt�c���y�\�t4�������oq���}�O��n%�bX�s>��n%�bX��{�� �蘉bX��}��7������=�m�(��[�_X�%��3�]&�X�%�~罝&�X�%��g��Mı,K�Γs�,Y(bf'��z(�Ԫ�#",�n�q,Kļ����n%�bX��{��K�@�LD�����7ı�|���/�L��L��w��uQ�Gq�1�q��7ı,Ns=��n%�bX����t��bX�'�Ͻt��bX�%���t��bX�'�ϡ��9�&qa�79�Mı,K�Γq,K��y�~�t�D�,K���gI��%�bs�ﮓq,K���B�rf��Wuы�"n���N�\u,�i\�=="F�2�=u�v��v�ݞ�8�������K������Kı/9�gI��%�bs�ﮓq,Kļ�g���Jbf&b���r��KI��b���X�%�=��7�@�$aZQ�5(x�(��q,Lw>��7ı,K�v{:Mı,K�sݚ�񉘙�����H냘:��9�n%�bX��{��Kı/=���7ı,O��{Mı,K�����&bf&b�ӯ]j�l�+�H�1���K�1����7ı,Nc���&�X�%�~罝&�X�%��3�]&�X�%��zW�ͦnq�fYq&3�9�n%�bX�c��4��bX�%�;��7ı,O����7ı,K�<{:Mı,K������;6���Z�^�8��-q���S
�g\<�i��&�L��vmp�&n�L�*^�X�%�{�~Γq,K���ﮓq,KĿsǳ��Kı>�=�i_������ut�uQ�Ge	G-�n%�bX��{��Kı/����7ı,K�{��n%�bX��ﳬ_�����{�L�YB����bX�%��=�&�X�%�y�{:Mı�s?HE�|s	���L�g�� đ�� D�1�M���c j�"H�p$F�3Ȥ��\XR�$"1� s�Rƴ�0։	�� �7� �8u5�U'~neFC�3S,���4�D`R�Cf6`L$*�V�t0�5!��c!B���
�t{DЄAxb��
X&�'�2�a�����d��@ڨpP2�x�9@�S��U� t]��@4�%"���AN�B��Q
-y� �蚉q｝&�X�%��g޺M���������c���v�U��񉘬K�����n%�bX��ﳤ�Kı;���I��%�b_����n%�f&b����FZH��k�&b�,K�w��n%�bX��{��Kı/����7ı,O��{MıL��^J/w��XR 䤔A`�[�b)^Χi�b�%н����F���ccsS���/�&bf&b�/|���,KĿsǳ��Kı=���A��LD�,K���t��bX�'==u櫖��F�X�1313���Γp��D�K�s��I��%�b^�߳��Kı=���I��%�L[�����c�c�-V��&bf+��}t��bX�%�;��7ı,Os=��n%�bX��x�t��bX�b{[�b"mJ�r2c��b���L� @�Lw���&�X�%������7ı,K�<{:Mı,5#*H0h@V���@��cﮓq)�����]褝TuQ�BV���ı,Os=��n%�bX��t�t��bX�'����7ı,K�;��7�L��O��Ie����n��$v�b��ޕ]S�3��^�wF�G=n�c��3��\�1U
�z�񉘙�����v��,K��3�]&�X�%�y��:Mı,K��}t��bX�'q��Xy�����m��b���L��]��^�n�8���%�}�:Mı,K�s��I��%�b_��gI���W1�O~�^ʣ	mr���&bf&a{�~Γq,K��3�]&�X�Ea���y�߳��Kı?w>�t��b315�}>��70u;-��񉘬K��}t��bX�%���t��bX�'����7ı,K�w��n%��L�����r�#VH�$���&abX��{��n%�bX~#��߮��%�b^�߳��Kı=���I��%�by�2	3�w�n.,�2g�$�Β�y^�-SF����@$A��g۲��bՎ�l��ݹ��ѣs\Ӏ�j�9�n]�γǶ��v�������-C���n:�X4��wH�@�)s轷G&ԩ+ǆ_�?㾱�kA�a##Vgt��`�W�=�5�ZB�ez��21:��!��v�)ۣ�a�j�՛�:Tdv���5[-���t�0��ۆĸ�RM1�l��.eZUNh��d�!�c6'�-�����nl�k;!h/ݶ��s��:����"%��L��L���y�ı,K��t��bX�'����7ı,K�=��7ı,K�{�dcR�܌�;^�|bf&bf'�|��-ı,K��}t��bX�%���t��bX�'����7ı,K�ކ1;Dꣲ���u��131ww�z�q,KĿs�Γq,K��3�]&�X�%�~�}�&�X�%��s�`gr�X��׬_���وJ�����n%�bX���~�Mı,K���:Mı,K��}t��bX�'�����"*����u��131ww��Mı,K���:Mı,K��}t��bX�%���t��bX�%=��.\�l�ۃ�Ϸf�>��{m�+f�S�fSMۛq�׏=�z�^�6j��q,KĿs�Γq,K��3�]&�X�%�~�}��D�K����=b���L��O~��FX��R�9Γq,K��3�]&�,H�SdE�E��M;���%�~�t��bX�'9�z�7ı,K�;��_������=u��F�����7ı,K�;��7ı,Os=��n%���������7ı,O�ϼ���131w�辱���!.s�&�X�~@�����~�Mı,K���&�X�%��g��Mı,K���:Mı,K���)�������n%�bX��w��n%�bX��{��Kı/�ﳤ�Kı=���I��%�bp��o�-�s�G]nE�Gsxݮ��t$j9�cSvQ�G����Aۋr���O\�}��oq��K��}t��bX�%���t��bX�'����7ı,K�;��7ĳ1~��gr�X��׬_���X��w��n�8���'��߮�q,Kļ�gI��%�b{�ﮓq^Y�dx����:v1y�����d�&�q,K������n%�bX��w��n%��q��*`���H���L�A���L�?�t��bX�'}��4��bX�'��O9#	mr6ݯX�13<��)�w�Xn%�bX���~�Mı,K�w�4��bX�'��{Mı,K����2���`;m�/�L��L��^��ı,K�w�4��bX�'��z�7ı,K�;��7ı,N���1�&Y��!�q�s�q�&�˙����Z���㭙�2�+�nɶu�t4�Ң��I��%�b}��f�q,K��;�M&�X�%�~｝&�X�%��g�z�񉘙���ө�_X�lr��[2i7ı,Ow>��n��"b%�y�~Γq,K�����t��bX�'��i7�&*b%�}�~���3m���st��bX�%��:Mı,K�Ͻt��c�b&"s���I��%�b~�~�Mı,K����_e���TU�n�|bf&y`�1{����q,K��}�f�q,K��s�]&�X��!�	���Ȇr pO�����t��bX�'9�C�B�k�&bf&b��w�_��%���޺Mı,K��{:Mı,K���4��bX�'�R��3rkq���m��n5�eNz��N 
R2��qmۘ;�ձϞ�.�N��vq"���~���bX���߮�q,KĿs�Γq,K����M&�X�%��w�4��LL��_�š��Q����׬_��%�~罝&�X�%��{^�Mı,K��i7ı,O{>��n%�������}#,mLn��n�|bbX�'��zi7ı,Ns�٤�K�EHb&"{��Mı,K�gX�13136u��\�H�n) �Mı,K��i7ı,N��4��bX�%���t��bX�f"��}�X�1313�y?�-�Q��1�d�n%�bX��}�i7ı,?G����}ı,N����I��%�bs���&�X�%��� QI��(��?@p���vo�y�A^�tj�� �qۙ��z���N��n�`�]:�P̳4z��ps��+z��b6	�KsZm��8��lx��ZuƟ�˲[���c�ꔽ,�Y��]e;N�F�9��<E��#��A�d�u dnp�/Wm���ۜm�	F�z��=hw���bd����l�!;��S�n��zCn��㟾�\����z�n�$I��w�ϻ��w{?|��*y�sV�s֎����N����Ψy��fۨ��k���>�C/�e`ՖY�\1313￻u��0�,?�=�����%�bw���A�},K�����n%�bX���~�G�Q�Q�n�|bf&bf-����?(�LD�;�~٤�Kı=�~��&�X�%�~｝&�|b�"Y���Sr�X��SX�1313;�l�n%�bX��}�i7ı,K�}��7ı,N{���n%�bX��;3�D�C��d��b���L��]�}�i7ı,K�}��7ı,N{���n%�bX��}�I��%�bw��w:�	mn�٬_�������{:Mı,K���4��bX�';�l�n%�bX�w=��n%�bX���o���#�*ƅd���
�1W�Iv�u�
ې�-�'�����Œs�ŗ�t��bX�'��4��bX�';�l�n%�bX�w=��n%�bY���{u��131o�^��r�#U�1�K��&�X�%����4��B��� !�(�]8���&{�oI��%�b^w�Γq,K���צ�|b�ŋx���������"���c9�M&�X�%��{����bX�%���t��bX�'��4��bX�';�l�n%�bX��ﱇ�c&,����t��bX�%���t��bX�'=�zi7ı,Nw�٤�K���1w���b���L��]S�1��J�����s��Kı9�k�I��%�bs���&�X�%�����n%�bX�����n%�bX��Q?{�q"n��'Z՞�2�
�	r���2�q#�enwGg٣�s�̺�������u�bX���l�n%�bX�ｽ&�X�%�~｝Ѓ`�'=�e5�b��ه`��IV� X����5�,K��{:Mı,K���4��bX�';�l�n%�bX���k��Kh�v�u��131?��n�q,K�罯M&�X��:�T�jD� �*�q5�sf�q,K��=�cI񉘙�����}#�'Y�Xn%�bX�����Kı>�}�I��%�bw����K���&��]b���L��]��5\�HՎ9qn34��bX�';�l�n%�bX~c����i>�bX�%��:Mı����릱|bf&bf.���Q���-�k�����
���*z�Fէ8�-#�C�gN�[��G�Z^�lei��w�{�K��;�cI��%�b_��gI��%�bs�צ�q,K�����&�313�9�0��J�lj�,�/�V%�b_��gI��%�bs�צ�q,K�����&�X�%��3�]&�y%(bf.����T�D�r[�[�bX�';�~�Mı,K���4��bX�'��}t��bX�%���t������}��V'd(B�Mb�Kı>�}�I��%�b}���I��%�b_��gI��%��`�uT���h��> �l��/�~��/�L��L���9��C�C�,�d�n%�bX�s=��n%�bX�����n%�bX�s���n%�bX�s�٤�Kı>�&K����b�si n��l��]&z���4ș��Iuvcۨ.�s����ʣ	ml�׬_������߽�&�X�%��;�M&�X�%��w�4�},K�Ͽ]&�X�)����1��Ȝdc��b���LK�w^�M��$q,N�߶i7ı,Nw>�t��bX�'1�{M�f&bf-���Z�[$j���Mb��ı,Ns�٤�Kı9����n%�bX��=�i7ı,Nw���n)���������"��G$�ʵ��,K��;�cI��%�bw����Kı9�k�I��%�bs���&�&bf&b|�;&1�Tm�We���%�bw����Kı9�{f�q,K���Mı,K�ｍ&�X�%��}I������>
)���)�Q�tXQ�G�>`��N�  Si�T�_�ᓏ�LD��C��X���ݠ��n�H!�)����$7�L#�pG���L��@�E؃��q�F+�I �g���w9�M,��5��j$��`��	����HA	��%px��HM���g.TM*@�ٺ��>C��c�Gju0�&X��N�cB������ E��c�~[��T4�nBU[!4eҋ�y�g~@�Hz��6�ΒE�*��UVV�#���U����b} v̬˴2��>��꭪ΉTٸ�dR[m�@	U�CR�v�:��@Sō9��C��8��
m�H��-JF3�qK%ȰsK�e�ΛY]4�u�dgj2�5:��C�VtRf�$����]��;��0��6�m�hIe��Ɩ�=ڮ�;�+bp�m�e+����u��tq�2�n�f�+�@�~G��u{�����q��)E�~zu��&ۍ��v�A�<�V݉����I��Kr]�6ݺ��kl/I�ԦʚF�����
�&��8!ļ�>ϒ6���X%u�I��T��Ӵf�ݳ��M�I�'��)9W�Y �@��LӍ�-L�8%235�2��`�N�/�����L�M��<���5&�t�
ntZlʻJ:�A֐�m7m[P8�)��I�#.� c/V�<+X��皪�)U��:Oko��zY�!��R����u):�#3@\yL��`�7�֮�)Z�m�0�H�S=+4P[C[v�8�T��U�����h5v:���+�G7M�ق��U�
Z`�b�f�<.L*֭��l%ݷE�%�`$=,�FjS� �@��0�I�.��GI���2mֱ�Fw"�v�Q�>�%ӑzCe�ua�nH�m��x�]f{]D���u8M���f�T<�m`���G��1�[�ٱ�vd�^�����an���c��	�<૵��Ӓ�m&m�Y�d�
��n��3a ���\9�R���e�Ӣ�5U@rmj0ý�w���lLP�[];>�^�]����k	��v�n��R��P^�9��S�v��! <�I,�OS�vtO���澉�mht��
=HN�c
���E�^[P�����F۴˲����t#�H��M�B�kaf�N�5#���w�j�U�.���o��m�b�R�%�ų���-r�恐����Y�jg5F%s�e��l�ܢ���*By�m ��D�1��\�dʆ��T~Ax�@4�]t��n	��32\��c�wf�я6R�:��ef�v$�̣�4�C��q�]�^�IAY	��i���H�J�=:춡��1W��Z��.#�;-&�A���-l��ZqX]����;>[����ӷhN�G8���;�-.8��F���au�~��}����˚�sP��6���Ss�؞���b��դX���kf���-+��%�Ǵ�ı-��̟�+�J;M�v��`�a�CT�ƗX�r/\�:廵ڃ��#��R5NKg�/��������kı,K��i7ı,Nc��4��bX�'q�{Mı,K�ϽL�"��[j�/�L��Lž�-a��%�bs����Kı;�{��n%�bX����O�1S,Oc���!ѡ�I*�/�L��L���~Ɠq,K��9�cI��?�b&"w߿l�n%�bX����4��bX��ު���Q���7Kl�/�L��N'q�{Mı,K���i7ı,Ow�٤�Kı>�{��KĦ'�|>���dq9,�/�L��V'��i7ı,?G����I�Kı9����n%�bX��=�i7ĳ1o�}���G ��jF�d
֩� �^��n�V�ܛ]Mu��]	����;8�1�[��Mı,K��i7ı,O����7ı,Oc��4��bX�'��i7ı,O�{��ng3�q�����4��bX�'��}t��P
e�?���L���j T+UxF��\~���'�~���n%�bX���l�n%�bX��}�J���13�{�21�J�li�k�n%�bX���~Ɠq,K��;�Mı,K��i7ı,Ns>��/�L��L��;�}T����rK4��bY� ������Mı,K�}�f�q,K��3�]&�X��X�!�ם��/�L��Lž�y���%vSX�1313w�����ı9���I��%�b{ﱤ�Kı>���Kı8s���3L2�1y��ݹ�N"[\Ze�ҹz�*\���stoX-�[iݛ	���w�{�K��3�]&�X�%��s�Ɠq,K���צ���O�b%�b~�mk�&bf&b�C^�(����Mı,K��}�&���"b%�����I��%�b~�l�n%�bY�{���/�^Q�&b{�A��vFD�b��9Ɠq,K��~٤�Kı=��f�q,j���@`�j�D�N�?z�7ı,Oc��4��LL��]�F�|Y-�5c�2Z����bX��}�I��%�bs����q,K��9�cI��%�bs���&�313�����dV�+��V�|abX�'9�z�7ı,8��{�cI��%�bs���&�X�%��w�-b���L��]\��>����ʅ�6�;l{^����Oj�O&���J�n·R�"&5,m�Y%z�񉘙���7�cI��%�bs���&�X�%��w�4��bX�'9�z�7ı,O�Lq�R�F�i�,�/�L��LŽ��4��bX�'��l�n%�bX��}��Kı=�w��n%�b_��m�xF���I��}��s�ՠU�נs�S@�^fk�s�ܠ�@f;b�LA��b"5 p�`� %
�C`h�w}�4w/�I�8��v��v��j��P}�4ꋻ�&��tv��qp�.��{).��#�7)vW��OX�OђE
F��Li�zܲ�׷s@�j�:���ʒ�kjF�U��S@}�����ě7�νǻ�}�)�s9jL�7�$�i�92���k�t�o_�| n�hB�HYqhrנ}�)�^�S@�j�.+Oɫ�b��x�7% 3� �m��nPq�@?DG��  ��8�|Og9�ə���<Hu�aΪ���G]u+��&����S�/��Y�:�L�:�H���lT��L�mT[�I�h���m����t��nII�͞
�N���W]��k��c�V�'���=f�w:�q!��Y��4�vY.�I,�d�:nsm�Rqau�kF2��1{=6��<�.�XԔ�l��`� ]c:�p�܆�ih�sy�R[U,x�f���K�%�l-십�n�7U��牞�M=�k��z�b�� ۟��4@d����e7(8� 3P��c�D+h�KM��������{�f����K@s{�5�ēg:��uFGmn�j�ӽԀ�mB���ܠ��B�Q�O��n=�[��^�p��M��;�����{4w��D�Zk"M<nL�/{)�s��hrנs��h�aq]�i FG�b#�d7cWK����El��uΕ4tu�p%�q��Z^H���8�4qڴ�Z�r����;l�@:w�C�ƒF�Z�7K"=���Fly![J�؀�v��]_�W$DmcOr=��s@Ƕ�tDDD��wJ��R�ֽrVD�4@d�f���M�v������s@�x�0�Mare7(�{��{��7{� 1� Cg���C`�_���'[l���&:N��e3�F�MRn�ӷ=c�]Ǟ�z�s�%X�����1�{l@fSr�ޏzPs�/F�<#I�n=���4^�h�h\���%LZ�k"M693@�즁�;V�7��3>?~_f=f�Tb�{��RO���ԓ|��6&�4�M7���;V���^��[�����]���Ѕ�4�������1�{l@fSr��\�\�$l��&�mfO��2ce�������K��`��n0+�G��=��4�#�UwH�� 1��M�} �{��}���4@d�f���M�~���2n�t��u 3P��c�D	�#nC@��@��@�-��9{)���e�q�� ��qh{��߳���{4���h���ά��31)�J C 41z� ���ﮤ���	�F�21<�@�-��>���9�j�:���ʱ)ZCnE���8�^wN�:'r�:�b�1�뱞�Ժ��7gv��L�#md��&h^�h�h\��廚�-bؠ�F���U�؀̦�����ڄ�m��l8s�tQ���6Ƭ��Ǿ�h���� 3+\�2l�j\]�uRQ3Wt��mB5�ݶ �FbX��;٠9�wYYc,e	]�hm�@w��� ��Rq��	*4Q�A�@�A�Ov� &Xי�M�S�Q�\1��G)vh� ��ٌu�v�ݩ��ۆ��%!�ʳ��FwT���kl�7/[�����ø�l�N`�U9��[rb�\q΍�zYW��z65������6�b;jʻM`�y�H).�oF�f�nӳH]�[1��=�8�q�xݵ֭lܜ��a޸z[��-5�@��AΩ�嶷^+�cW'fY��_׻����/���0?�ru�wV��^d���/"n+i�n��gn<qQf"XFә�=�g�������/ffb_0�{�- w����TdwvM��݈�n�kj�P���M ��pB�Q�n4�N=�۹�cmB7m���H��f(�E�SQ6493@�۹�s���:���=�r��f��{�[��q����bgu��mB�mBCm;�K�s�;�������1Н"�7�3�y1�铝�v<��&1́����m�̀�uBwn,�/D���Ը���1��g8ԓ|�tk����> ���P�׶�N�K��G�26�z�.�����@ow(@f�����۹�uZ�"��5�m9�;��ηH��;ޝ�� wD�1�ꌎ�:�v�o|���ĳ�w�/�����9��h\K�������x�m�����9y��܆��K�y�̳Ib�(57!�8��n��n���S��
���_xK�H�n8ʒ����ݶ 6u�@}��@}ӵ��A<�'�q��9��h]�q��|�kl�t ��X	F$ �r ����$���*�ˀ�2
��#��'ݦ�#�����묗�*����F](� (q"ň@�B$A�hP�e Vi��Gyk&�I�Į1&�J�#	�P�0��^(���@� D��!ʹ�`}�3�;����4Z��Ã/ȇ�pU#� �P6dD �\	�p�ҁ�S��0x�8=!�N��CN�����Mf-��NkK�0�;�- s��U�Y#K�����^��m��9�w4;����M��ǎ>�UdMH��������ݶ 6u�@c��K�z�\Z9՞�R�S˘�I����ewa�n*��.��r�t��n�cX�@��ڄn�:�w��� �Mb<�$���h�e4����n��n�[���Ɔ���E ����������m�Mw(59"���z����9m�Л���ԝA�d �W�B� (DH,Db�0�P E3831�����o����~�[j=2�$�WEIWp��ڄٶ�ηH�^��}z4���ڄ��,��Y�\g����b(�^θm#�C�gN�L�q�(���q�π�l�uvנ}���|����4��"Ȅ,�k��Wk�ވ��d�|�ϹB��b�:'{15���&<�����{n��;)�U�^��ۿ��4@d�b����<���k�u�@}�� :�OY��Ě�&���vS@�[�٭B�j��x�=�A���{n�??7�$���F��2�-��Nuԝ]�z�h݄��m�Ƙ��Au��J��`�hwMѲ6�z2_4�/;Hĵ���t]1;�9�v�D�m;��FI��]�V�/j���[�������� m��$���u�8[��Vr*�;����N��:��)(��d!Գ����ː�{o:��,�,�jMev��<�B�*�Fj������bj����W�D_�G��4�!�^�k�Zh�P�2�b.-��{WJ\󶃱�c�\�� ��$<�/��?���;w4�w?�������4���B�Qc�b���f���@}�l@9�t�"=2r�$��JF�q̌��{����;)�U�נ}����;ZZ8����*��f�w] >�jP�;�����A�Hhw��s�s@��s@����/1��X�o�W��nc�hBp�ۂ.�++���͐�m��nK�\8�Jf&�Bdo7�7��;w4��@}��Pw] 5�^�*�.��13��ԓ��thR	 ���`�c����IJ��H�Z��ٯK��5�Cs4��V�U�z����-���q`����ԐQcr-��H�Z�z� >��(���/E�H��%#�[��������>o�@u,X�;_gQCdc�P�N^C�R���u�]k�&��D���/V�X�JF��rg�{�ۚ�}�@������h�i"O"m��՗W�����H�Z�z�-�H{c�B��X7"�*��@���@Ob��4��&�@�*�4�?~�4jI��~��;���	��X�$�z����-֡�ֹ@��^�뒠������@c֡���;}? =��۹�w9L����y1�@���?3��*:�[�r5��]�s��]���s�wzf�����ֹ@���֡�n�[���Ɔ����hyl�>�j��@}��Pn�K*nb����M���/n���Z�[4�ڒ�&��%$�$4^��I>�;۩$���u&�
+樟j��Q��*!�U����{4;�%��ym�6���ڴ�{ވ�o�������ޏG�"��8����z!8��l��s�=v��*���K�<�:��w7j3T��c�'c���e��� >��w���(����Bdo7�G���M�۹�r�V���׾�ٙ����!�(���X��ܡ���w�ޙ�o� �_o��c��MƊ�*�u,���ޔ ����؀ǭB��󊑩 �CR- �-�����9{w4&��v�I�����0�S������6��k�#�GRi�n�"ײ���}?s:�Z�q��B��(�z-�.n�W��D��M��d�[�9.�����NCM�����N`o)���j��QRb�;Pc7g"70c��t��%�l���<b��#�[a�7dz�n�^�V�s%.�=�{ZumŹ�����(W�
��vθ�s�1�B��U�
�(٥��/
w~�����{�׻�ĳ�߿IU�@�Ӷ��q�*� �tC'��Xb6��^�L���N+���<K��Q��;��nh��hu�� �m�ݵ-��HФ�m%&h��@}��P�v��v���n��DM��()3@�v� �m�{e4[w4�c�ĲB,ȴu�@n�b�mB7(��5/!27���&���M�[��r�V�?~�.��ı.͝�9dT�QF�zJӜ�H������dS!A$�u�[[�+3ٙ�"a(��>���4Wj�s�h��*���Px&aN�}�w�^M����I\ QM�)�3@\� ����*@@�"��ﳩ'�w?�����Ѡ>��Y\hjH(�ԋ@9�٠w�S@�s@�v� Ϲ�EG���b��M���-��+�h{l�>�j��6����-��:nP�v��v��z"";H!�k��{h͢x����q u����Y�H��dpǐj<q�	-��X�Ŋ����wJ �n��؀�ڄ ۧVA,K"�`܋@;�f���M����ڴ��?&�Bdo7�NM$�;��I>�{�S�pb0 B"f%嘒Z����@�{t�s��ʋ����@�s@�v� �m�����9Z3��Y�D�	��>��Z�ݠ>�j�P���G�1�2ʡ�9G��s��۝p����m㗘�浧��l�]��GJ]ǭ�z�s�%X�%���>�@}�� 1���ֹ@dK*Xܙǎ94�۹�#����ՠ�@����F���m���jmk�9��v��u�@}�f�D�qₓ4��V�w����5&0�� QX�@�bP��E ���������=���q,p��r- �m�����9m��>����,ŵ�޿��v���$���wJ6�k��3�\�]P귳n�_Pnż��	��X�9>��s@�s@���{?|��ޚｿ�&���I�m�]�>� �u�>�jDL�����d��&��Nf��w�����-���/�I*n�z&[�}| 1������EG�,q�7�rh��'��vnI��2I���u$��Ƞ���
���@W�� *�PU�J�
��T U�PU�J* ���F �E��b,Q#P��b�cE�P�E�E�DX�cE�AcE�QDXE`AaQ DDE �E _� ���@W
�T Uv* *��PU�J�
��T Uʠ��� _�PU�PU���
�2���G�@)Y��@���9�>��|      �0%  �   #T  h�}h;��$��T	 R�  �   IP�
$J�*R�%@"�R�( �@  �    L ��  (@�)JS�J:s��E=<l�(�f�W�x��zR������NO\���/}�@��J�}���6��  ��u�rz�������m}�Z������_[���n ��,[�W�Z���,�.N��
 AE V �M�R�r3�ͮ����]�ۅW��}+�n���[�}i�w���U� ����9�� �r�Kn-h� ��+'vz�Y�x�uk��7� ��K�9o�ί�{�}s��W�rj^� ��U@    c� 4����X�W6�']yw�ʦ} z^����Yoy�{�w�K�Ͻ���{���}|��i� ��gK��uK� �sk׮�.w��OK���ҽp��ԦOvS�\��}5qev�   � P  ��w�X�J��^��ͮ���yʸ ʕ�z��>����n^��iS��m7���� ӗ�ow^m髀��J;�NO�^�OS��m=7� �=K�{e{������}���J�� � 
  
�@�_mso���Ϸ�My�|���Ү� �S�JR��s����%�s�JP�&�R�J�JR��JR�i@ tӉ��)����� ���M�)�J\�t��q4�
14�(��N�SҜ@t��(�K�
P��)* OHI�T�  �RmM��* �O��*~�i��2=��)�*@  S�	S�*R�  "(&)I �)�P��{�����������Km��r��FVVu~��U�Y�dPQW ���pPQW�H����b �*�8�!!��1��$! ��b�X�V�H�!dHI����#R"I����E`�쐡�8H\8���b@"Ą�F��$$R�B+dx��4J�� #\��� ���*0(��@��"�V!&2�����"D#V	 $H֤��`E�dD��b`�`�H@	"P0�Xl4˛��L����e�%e$��Ѱ�+L�!1A����!$����
��� @�H�O�\4�R��z:H�q��&�"��BC�#coM���r�Xa>�E!����XLM�2�Y��̆���˃$`2�
`�t�x�%�K�$�YfB�u�h�*� E�L �(d����$��t}��	%���J�@�J1H1*�0��!�#"E�0e$�C$@����R$�9T��X�YIk��N�l���bћvP�V!"E�n�1��D�h`2A(R���4cI"a�Vb����5. �/�`�!P$$�	�
b�@��ÓA��I���l P0F`�B� �^����
��#`]�d+�Iq��Ɍ^^3��C�U�$Cc)�㗔6Ĉ�$9�>�.1�D5��%a��Ca�ԏ�5�kX9�Ð�X��� �XT�._��#K��e�)�S�A"U01�n]�i����H�!���11`��",J��z	w���!{�sr�0�f�ٜ�$H� ,D��h`B	A�%��#���$Մ�4� �H2!$ a!LDha�E�!
1��� a�XYq�ٓY�7�s���8���l���.V!cB0 B-	�e:L����0`&0¸�1)��cH0`�(H�\���ɸ�cu�THBa DL0�� 2�̘6�	6���Ԧ �  U�\ĶgB�`c:�c9�\��|�}�Hd����u:���]��_.��\.j�8-O���qLT]��r��MW����aIBLԁ�P.
K�l��6J��.�K��8�5�3��F'!T�Zf54cy	��2�3�rw� F+�5B\A B���9���asa�p��Fk:�J��d����3r�Š/T" �!H5�c�"S��k�٠$b j�:�n#�D�!I!$ A"�,.� �2��.>:�8�2,y�P0j�
b0�	d�55+�PL����O�.t>*G8FMX�\M+	l�>J�JSWb�\  i٢dgxٌ�7Hk��`���̟�!����9�'3b�b��/�|h�5�v�	���$x�̒,`I�	C�6��$$"Da$�0�IC3�0&S	���:B%5	+���h0`�@�CL��,�2���Bk��e1�����O�HM9u�i�����
�bP���b�-#	R`��%�f	npE�L$J$)�`�(�0&1�6�a2i�m���pdXWX`S�bT��0��Å��f���°$� �(X���}1�X��`>)~�pF�HA�İ��2�&)HI4���C��$--!p�`�)�0���B�$\�,d�`H��a�[,B��Y1�bx)�ZSۙ�����q�!Wny��HU`H�!R����ݒO����J��HՉ.�����d>I�ݕ2Hfċ�cE�Ջ �@�b�@�pi���#.3	hJR*J�	q*BnXH�ΒD"�D�	@!�/�Ba���Fȩ�|bS�ٳI����GHo\.&��T>4һv�s�@�Cc ��cR����+�B$#���0@����Ù!d S�\!���"I�kL�ы\2�~�q�9���N`U0�*v-�6p�A
�s8%R	L�1�Y��glhB8H�ԁP0�X'J�
$dv1���� �+���+�y܄������7�XS�)p4�5�K$fLS1�\hƲ$a`$ܒ@���	�$�  !RFᗈ�D�!X����B$$��
�ZȲ&�F%01>b�Fp��c�pB% ���`��@i�"R#D�V,�D�
1 8�r5�@"��U�#� :H,#p("hbF4�q.%�L1��0&��[�Q�.	##!!%{���$B@$B#��F!0l���94rI+,`D�i
$Є���	#�	h���Ƥ�'icd�H	\9���\*r\R�0H	BH�I	 |���s���O���T�Dhu!�7�Cq!���Q"!��D7�o�,����H��F0X$�*D��ŀ�B�)�0 P��8aR�0˂A�	$9CR��$Q\��ӟ�hU�bb�<�+��6\%�	p[s)�s.�}tT�&.SsW�U���a"B+!�@�Ԍ$d���g��a ���.�nVIYHa���F4�[rb�n����e���� �	���c���fI�f��}�iP.�ݥ`� �	�+����{�L�#d"�J�� �bňI8�S�2pe1���C:7ψ`�#2�� � � �AB0N!(Jl�1��!X�e6F�#���rXi%0�*J���R4��Ѓt�>7uu�� �k����Y8��%L@m Q"K�%8"�`����A���&3�����˧g4��);a5��l̺��Mˮa�2��$��!H���,�-�#򒐿|L�>ɒH��mC2F;0���2�hƬ��2m�0� ��B�H�D:�d�'؄7��`a#��10�X�aG��\��B����{�a�	3��l����
�5�����v8��RS.P�$�`�d���~�S�FeHP�R!����*Fg���%%��d4aXu�YS�У���q�cI��)���-.H���er�AX�s��%t"QN�YI�s��6i>��R���m��%.E\�Qu��d%!hF,�b���5��㤒HFB?ZBBB���#ӷP�SC��1
B�"����H:&#��4j;H`�17�{3���U1$�"�B��@k�ʐ�,H�HEc� B!���Ꮷ�H@! �"�2X��"��9\GfМ�$L������I�!@�B�.�%�у8�r̘�	$�bd�bL,*�>T�rU@��C	��!��P�jF��� �A��X�p�X�g[�B���g3��$cāC4
��0�����^���we�^��>Ǳ짱�A�!M孉�S!$!�j��0��*�>��~����������j1(}^gY��nϋ	x	L`C+l�F�&2�3���9~�~2B�!�`A*+)�\]l�6c$H�V2bޓ�B!
�����2�HH = T�X�GA�K�B�R
\����4P@B4�׺���7��I��NN�s�4#���X�2��M���Si�
�
�F�����0dHM%�!}�7�T�m�ڭl ��8    � �   e�[@im8�?^��2�����ݰ	�l��	V�1�棱�uյ*�E��,]�T��/��rڝe[%sZ��0�쫳[! A�@�P)^ܶ�-+`f��H�i�:�m��i4��m�&��VăȔ��m����h,5�U���  �j�l�-���H�7-�5��� �l l��부r����+2�T��
�V�&��+��@U[6� �lհ,���k�8��5�`5V�/R�I�8�G ��U+.�l�UPj�;��x���m�T�(u�4����U�X���)��ZMV� �nh[��sm;�[@m� 6Z��%����
�YL�  [KoHu��������v ��Ŵwn:a�
�6��ض�$8-�Z�싱J��`+�|�v>mb���̴����.�e�ۋ���o0hQj�Vr�3�J�*�0ų[d`B@5�L
P�m%�v���`-������ mٶ �� m���8%�v�6�B� /S��������ذS�H%����	�zX+teeUT�%emlU]M�cm� �u�-��	6� -MF�[׮������lM�뫮 �l�X�m�:�m�� 8	 ��k��H���T�kY��.� Ԙ    �`p�&G-�[@ �a4�n��ku�K#�� n�N�� �ݶ�p5�R� �i����k����mm�	 m�m@+/5UU�G��[M��m�l   -�V��j�
U��zU�Kz@ m�ڳb 9#�i�`Eˉ�gj�VU^e�]�.��@$o�{���m� $ �E$  6�a������e���2�p�U;`H�@ �n� қsY�����$ m-�@[A��i$� ��ڶ �m���6�m   6����  ����6Ƴi���^�ݵ��rl�����@ �[� ��    m�l$   m�p�>v�m$�m�  �l9���%( �	�� -�,��M��0m[]ye�m�mXր��Ji�ԕ�  p���V ��m&m�	��K��	������v]� ��Zz��	7Y��mU !�F°t�M��C����-F"��n�9̳G�
U�`�v�� ��n�`��ź���m�MT�  l��l m%M�$�[V.�M��$�`�-*Ԅ�(��!m9:^����($�` �E�����[E��V���'�કiY�5,:�m� v�ֲCm�[Al�հs�ZXmjL��	�\[Kh8$6�-�qm8  m�m��a���l �  [Ki�ְ   !��[&�� �m� �q�lm�4Q���k���I� �`6�n�` ��%p�v��]��qm  �l�����l6�m�m�m�lH[p  Ѷ�� �i ���Ͷp $��p$��&�m�  mڶ�m��V�,�մ  |߀ �z��-�X`�nm��٨  +�&��E[Z��J��`m���ܐc����� �jͰ���6ط���  H� ڐ�@ �۵� l�9i�zl��C[@-�!�):P��6���J�KQ[��kt����P M� %Z�⪯J�w��%W� [@�Zmm�v[���Xb��km�T��5m� .��[;
�dZU
Ukcf��m=k�B� ź�%��c]vU�N�;����y��wl7i$� i�6�����R��h8$��5�$m���� ����"@ ��]�]XH���l��$[B���`,Iv�ܷZm Gl��a}����θr�լ��أ�ֳ;tb ��<�J�/��U��kn��,���W[J�ɜrڒ�$9���CZ,0 �!�l�am$� ��6�p��@��݀l��  ����    �[[-   �m�p����	��m�ۇ  $[Kh�Ͷm� *ҭmr���] �+�@�@�m[~-�m � �H@H���0psm�lm���  m�l h�`  �`   ��e�ɤ�I@����٪�j�m� �ɶ�� 	  r�X�� m�#m� �Ԁ5ه[d  HI��[@��5�l$�K{T���;�~����@����m�`��̓`[xp�n�Ta\͒�Z�����K�n4�+�n��9R��Z��-�����x�e�Z��B�087Kl�G��F��YerKU����̯-U/"�;COZtUU+�UW[NB9��E�@J��V�Z�V����A�[�h3��j)6e����j�o`2��m%v��[�[���e����rj��<��G���]ձ������jI��w$�[C��n��U�sf0ңq]@*ԫU�Tvٹ��������IoP��km� ����	 ��H7e��H >]+o� ��6���O5UU:��ϊ���km� H�� (    �yUQ���ڪ������H �GHlOmt�������� H���*�yٌ�T�ʬR�]���Uj�[v�`ⱐ٧@�4u*��Y|+L�,��z��5�-�v� %�t�d��6�m�P��V��S�9Y�e�m�m  ��+��$[A��d�hٶ6����iyQ���n��l��@  �� m�Y[l-��:@)ն�UF���V˂@   8 �K����h	�ie͖t�,[� @GT+���UJ�����m�K���   �Rtmm�'N��֛��!mI����vZ�� q�8ju�u*��+����F�6X)��-�<�5ufd��F�;��@R�iV�4J�mm[Z�� ��N��ײ^$�d�0-�ņ���ٴ�Mv�[mĀ Y�MU��� �e ��sCf�mj5`��:�:06�6�$,�ےF�  [v������6S�^�$��~�Q@7'6��W4香�n�غl<�� ��[s�m���:��m��=��[��8H 	i�����݌`�Ҭ�+�xh
U�Y��'a�L�nH�PWP,m���m�CY��$���	�.�a��]��n��R��{Im[h,���Ujj��p��-��;t�kon-׮m�"K�pqt�P6u���f���m;3l�I�e��z�m�m���'Yn���Sm��E������<DC�2��XU���V�@�Wn��kٵ@Qg�����U5����ܝ�ҐJ�W4�UU[A@ 6�SmzԞ�K�չV�R�*��BS�N��3��v�m�8��&�iv�k�wq��ہ�n�pٖ�5Snض��,    [z$�[�εn�� �m��m��fvF 8]��z��p�i�h�8�8�M�6�mm�%�H mVi+j�L�����@XbM�,.�eJ��q*��F۵*��N���l �Nlp  �H��F�Z�]��� pVڪBke@j�6�p�*A'-�n$$q��[7\� ��� r�6�m�m��p[Ԑ�~�}6��$86� �o&����Wae�@l��	,$���� m�[v � 'm�[# 8�An7K�#�9��\1�H"Yv��h��M�[m�j���
��J�J��zZ�V��l  ����-�#'�v�m&��;F�po�m�� ��-�B�ȩ�� �4���[x-�$I�m$4]� ]:N� $� ��-�HE�`8Hև[3�_�o���������]/X�$I�m�h�H�p6팕2�"I����R�K��l�)/��h�h$��k2�ԥ��UZ���J^�B���fI	p ���BG-�y��j�70������ڒXf�X[s���v�l[@�YN��@�fMt�14��$��m�[K�(
W���m[��.�$&�tm�im��v�� �H86�JU�j1��ݶl�6�j��ШqsØ��]JM�\�/Y2� �-��-�mp�f�nٳl 	:Y@-��  �8-�ſIe�[~�ض����-i��bI�Kh   6��l ���� 6�t��	  �6� �� � � pm�9m�!m9%�ݲ�iK��kyI%$�e�l ���	 ll �6�v�m�� 75�jݮ��f�iu��\	��U���-��m�Ҷ����{�{���R.S��]��O���O��� GȃG)��C�%��,�D�U��@�04�4�`�@R�.� %%U��H�0���&�C���
E �Uп*)��ʜQں�����M/>CP$�E� *B 5H�Q��|�� ���3�
��"EPc����=��| P��E�8u��T�N�TTА"�D>U��U ��P�  )� ڦ:�L�.TpⰟ#� �Dx�����.��0f�
�� &V*B0b�W�~C#�"�8 :C�h� ��DH�������z���E�˕�$$����UH��p(�)�Aҹbac�,zra0��O��@�;'M��O�
g�Dz�Z#F�'  ��L�!���Z��sQ�;x�D@�hL���"=��� �R�� ���X(AE�H��T1r�;v"�7�	FB!"Ed@��B	���uW�S�l�.��~B��iB@�`2 H�@~W�T�beJb8�i��	�'^�"pN
�`@ ͕
A�E2��
��^*���g�T��((����� ��@H.�.����I���[Am�Il��n�K�4�%H�'Nz�Sn�+���A�Dec<.^��T��;�[�n&1�SG�p�⧜�π�s!�շi۶�b�M��:�)�:��Bqɑc���-eI�l7K*�,�a<��@�k��A�b3�n�YJ����V��c�� 灭�vW�.�#$�X{l�����sv���J�cY����VVN��u2��K�*��Rk:�&�����N�ʭ�T���V��0ざ����V���Nv���0�H^쭮ݰ��l��ra'I��:��j�N��E�^�����V�zh����J��v&�U;���p���f���8!�r��4J��6�m��R�V9�������2��fـ��i�g���W`��:����/f����\�,�q�i铯J�7j�g/6��y�ͺ��N���T�z�̻��u��U!
\6�<6��We�lЫj�3e�,]����ѧ��H;L�{=)�Z�I�Ib��9&�f�f����Z�;hr>{(o)1��%������e��#�+�u4�PT��o-T�Aev8��[A��Z���2BE�ٶ%��ii	ꖩHs�,��V���J��*DX���	�.Uy�J�]X���T�UeXH�b��@�^���$r�Z�U�\S�d��؝@e)[!hQ"�操���G�P#v�.�x%��2�lxؤ ^���[{(�u�4���:cv� Z��`y���.�����88��F��8׎S;m�,�)ձݍZ��)]6�FA�,�0j5�-��5R����ev��ݶ����+[�P]�:%�]�0�=v�:����F�'QƅU �Cb	�]i���Um��jY�v5ӗ;�L��
�B���&˴Gr���N��ͻ\&�c�1�1�"�H�//j^mԇgt�*\K x�+(�i�ج�a��W���W4Y@=�;f��X&iZ�)Ƹ@SF�c8���^. R#�@���e@2�~N�:Q
/�M�E>ڬCp"�����M��0 Qh����q�!�b��̪��k�͒�c�C�q����,t�;�Z;s)8�`A�R��-�Fkm9�b��q)��yN����]�ܸB�.U�;a��l%�*	b�vT��� �j��ٹ@�6��Lvm0��m8���Г�;m9z������	�u�eӹ�9�{���]�&�p�9̝m��A7Ik�Pn�,�%{�;���Qr؁��sV�Y�b�&�Ǘ����������p����H4����t�&��5���A$O��2��H&��1����D�K�������bX�'���Б�%��R��ɟ&|���s��n%�bX�b���j%�bX��;�&�X�%��&{2��bX�+����n�⥲�%�۟/�ɟ&|��b���j%�bX��;�&�X�%��&{2��bX�%���t��bX�+�Y�ƣP*��5d�|��3�ϓ}�w��Kİ~��fSQ,Kļ��Γq,K��3�ښ�bX�+�������u�V˟/�ɟ&|����=�MD�,K��w:Mı,K��;jj%�bX��;�&�X�%��?u;�Ο%k�=vڸ��jT܏3Sq�j����V5�i�v)�kEٹ���LY�̦�X�%�y�;�&�X�%��g�5ı,M��ޓq,K�ê��VBd&Bd.ໜE'4蚑���c9�n%�bX��q�SP�!��dp!�.n4	��Q�G�5��󿮓q,K����&�X�%��~�U��	��	�>1�¥�'RTn3�SQ,K��s��&�X�%���=�MD��C1���t��bX�Bܩ��Y	��	��8�Ʉ̒��bg�9�Mı,K��{0����"b%�{��:Mı,K��=jj%�`yFb'��}t��bX�%�;�Б����7KI���ϓ>L�>�q7ı,N�8��%�bo��n�q,K��,�fQ,K�������Ы�W�F�y��Z.v'g
.��l�J�vcZk�|i��u�ΓS����1��>�bX�'��z��Kı7��I��%�bw�g�	��%�b^}ܫ��!2!w)�U-KR���q�SQ,K��s��&�X�%��Y��&�X�%�y�;�&�X�%����p����I	���{3<��"���P�3���Kı=�3��Kı/>�s��K� �T�Ej$H�bb'y�v��Kı>�yۤ�	��	����iIR�i�$K&����%�b^}��I��%�bw��mMD�,K��{�&�X�%��Y��+�>L�3�w�9]%�V�۟�bX�'y�v��Kı;�w��n%�bX��3ل�Kı/y��^��7���{���;_y
��d7g��U���r��4�,aʒո�������ۘ0�8��_�ܵ��&|��g�gwf&�X�%��Y��&�X�%�{��:Mı,K��;jj%�bX��I�i$",X�,ϗ��ϓ>L�oYva5!D�K���t��bX�'��z��Kı;�w��n%�bX����a#-��v+I���ϓ>L���{�&�X�%��g�5�ʐ�LD�;�cI��%�b{�g�	��#>L�o7"7k"���%�۟/�ɟ%��g�5ı,N��4��bX�'g�a5İ:(>H-؉O&Gq7�k��n%�bX�{&��q��1��`�|��{��7���{�&�X�%���=�MD�,K���t��bX�'y�v��Kı/V���wmQB)T�5S��n4�v.�n��0q�뷷V�
�>���]��kX�s�&�X�%���=�MD�,K�s*�p��L���N=I.0כ�`g|�C�����0{�p��x���{�t�;���+NQ�GUV}9����ɳa&�1V���Xy��G\A,/�r[0<�O}}�zJ��1/d� �6J9ʲ�Y#��{�t����5�v`�s٩'��ۨ�V%9��B㰴�qu��a8���lˡ����1��J�m��ӫ5�O7+�oi�XC/=6�^g�Q�ƌ��]�v�@n{&D��g�wYۗ��=����-� ^T��wA�|�Ƨ��%��M�ނ�(�Vg�#�rע&��z���챕�΍����jbz��k]u��npf�n���^p���\���u���v�fpՐzS��5λY�$�ff�B#EH�s�R��6c8%7g��赫s0��E�N6�r�N���V�L�)~������v+M ��؀��-�2�dTr�2ȩd�Ie��ɺ��6s}|`�W� s�ۀsc;�5�U�q���s ���A ksy%�7\���#���B��^��`���7�u��u�掦�B�ee��R�I1�nq'$�[�������;����P�=����(���m�e嶖䁃&����d��U���F���45T:��<͛2s���V�q��{� ����u���RYf�7^�ű$A�o\�iA"R#�94�K �{�`q��7�Ca��5&+BBI^��|`���?>�f�7^ p�~�H�I`�;��I7��V�3f�̜�`s�U����� �T�X���pϽـn�׀~�U� 7wnׯ�����)Zc��]s�8c���b�r�bq/7^�m�=�&/�����@��8Ֆ�vn��z����pϽـs����GQkn�|̴u�$���8��{Ҩ�P�YX�Q����n o��u*�b �q�@���l���7��x��kj����U�K�b �� ��q�@��	ζ]q��;-�?n�0t�� ;���n��7gv�'	H�N �����|���J�æAUv:7g+Ef�*W\/a��A*C�AKv���{� ;���n��?wn��M�Y#%�MTӰ�ܫ�M�wv��kK�Su���"�EK%�K-� 9���2�Z �� 5��r�끕�e���f :�A �rK@��M��H�ʋ����:�l�?w^���T�mТ,�ީ�����\�wf��r��:������6�m�Ijb�"r��\9���]-����`�K�r��5Ξ���9���1�$��d�$�w��j����U�G-�8�v`��L�Su�;ݸ���Q��P%� :�A �q�@��nI�(ޭ	!�����i�w�w^ w�ۀ~{�0۷L ໢�H�Kcb+W2�nb�_}���΁��x@7\rԓ"�$UG��u#1�vf�9�-�;T�5r̚��]`݁.��uY�ko*m��i��u�M����l�-g��'5���`�ٙ��$e�[�۠� @c\i$��e��	������؛`��X0&���@մs�z5��q���xRM��=�ֳ�طl]�0޶��6��c
bS(��Y��#��W]sh�T�C�t�lJ7�<��]��I�Z1�����[�ߊ�� ��U����!�b��d���,;C��3ĸ��m������s��n��ӷ����TA��d�Ie��|��v�w�w^ w�ۀ~�hkmW��և�fq�2�Z m�@v�@s�z�Z�S�N�r�:N����p�wf�v�ozU�++,+�s2��@$�|r��$�����QT�qV�� ��ـk㖀n�%�&ȩ7�8圲�����p���҈�H9I��*B卮==WjՌ_��-u��Y~(�0���S���2גP��ڰF��s-�d1�\�8�ԓ�1��P	�<I��Y-@/0
p>�w|ލI'{ݸ�w^��ߦ��"[��&ȩ l���@7\r�c���R�b�9*�ۻp���S����,�{C[j��-hq�fb>9h�Zl��d����s��>����uZ�@��Q����pN{\GB2�]�a���x��"�p뮲�/�}J���&ȩےq�{Ҩ�P�YY`��� �n��$�>{�6���S�w�%	Bl�g�z�����Z�r� ��ogu�� ��tH�`I�E$��8#�da+3j��t%! t�f��� ��D���I�Cꩨ$��̩���
!ϱ���l"��L3!�z�i�k�F������E؁�j,2���GN��b�$cEmH�2 7�X�
oHcS ���)	4�b0!q(G�(`H�H��r��� ��hC��])@~��ڭP�D�&4$h�:r.����knn%��A�� �F�P��P�°�����L`@m�� �s�k�F!��8��l�O�p�܂�"	�'���S�|(�D>�9@��B�A^�ӢC T^�� �(8�)�U�z<�6gݺw��١pA�A�A�A�'g�\�3��fI��8Ѓ� � ؠ�>�{�pA�A�A�A�:k�B��`�`�`��w�4 �66����t �6
P�	C%��	�ET
j]UM;w�4 �666(��w�4 �6��"�w6l���wkge�N�������&��z�	2T��/��PV�G��}�\�.����{�w|���m��q[������`�r��{��Д$���U��=�Jrz�J���S,Ұw�W�	Bl��k�>�U���w-_��B�3Py���QT�-T�M���9ު����~��ǻ�oN���[�8VWLsN�TBf+����ڰw�V�? Պ@:��)�D��P(Q	w��y������US*H%M}ܵ`uy$�	D%Y�������|N�w���HڲYSV)�MQz���003����'��`�A��~�����uک(�XIW�o���0����/�0�wذ��y�XX'B�-@v��/U}��$3�\���/ߩ/�R���5$pV��� ��_>�Z�a(��>�ڰ>}͛E�rG,	���D�E��
""�7��>�ڰ1�ܛ��	<�/K �vSS�%**f�L�niX3�V�	/Vo��7t�}ܵ`
>M'�=��Oa���3v��Z��W�+(��q�_�zᵞ�ٺ��67R�I�ӱ:�*�ۚ;=qݘiե�{V�7.@��,� c��%���X�d�Г74��*������j�㗣;3���岽���sc������v���|LrRѶ3f
�[jE���]"���[�tS����WsX��J�hQ�N!���3d��nK��.AN*U]�c}?B�����e�S�;�wON�EN��Qb��ls
�.��۵���M���G��$s3 ���@6̂k��U]�7�ـoO?He��8WQ-�{������b�{}p|���g�J�<�b��T��M�6Հs;�g�/L���p{��0��
����j�ʰ=w�����q �2=���v���=c	a`�
� ����?�����x珀�o�X3�V�J1��UKuN��O��K���$�s$ۏ;�/n�,�D�t��ёwRKO侐.C	#��uH�����w-X3�_�<�}!כ�ǽ#�	mm
���?s��/��>I �]�Z'�O���׳�'�=�jI���/�
<�$�C�����%**f�L�sJ�;��Xw&Ȉ���o3
� �wذ.v�k�W����Im��_����w���ԓs�5'��� ���!��*p*��[0��a`j�w7��nmXw&��(]Sͳ�5�ڎQ�T[P�A�+R��9�5���K�=X�,C��6��_/�b��CVVR�S�*���o�X3�V��؄�q�zN�<�DnѾt��hsCTɚ\ �sj�	B�ϟsf��I�v>�Z�/��&�wJ����N�l� ����}��{u6�iZD��`��w��/��9��ѩ'o=�h��$�
�U�#�`y$��K�Z\�޹�����9� T����5T�!�4�}ܵ`lB}�mp>��u�����#����j��:�V춎vgg
:v�I��fY3Dj�9���s"je�T�X�`�\ ����?>wf�u��w}� ��U�ڍR�\q�Kn��3�6�����`|���g�����SQU]D�`����qR=v��q�縀��u!UXUH�dV�|�������M߹�jN#� ��w�U�������.�����eEVQ�5Y%H�� =�s�����u�Hއٷ���D�L�a"n����f������My;Z�ț��\�m�������ڗ3�m�� ;{Nq�qW��� @�S�\�P*t�\���N�ߢ"��S's}j�;��8��M�Ca�ln��5T��,��j�9�r��^���{��wW���bjm�T�X�`敆��w6��sf��˵���B�B��o�V�z���-QN�˖�]UX�s�W�k��tsʐu�@_�&���n��+��@+�T4l�a���8�RZNx�φ���m[Q��h���s�6z��i ם�dg�6N�s�VR �c�rdx%�g�ơ���H�V�8vM[AUn@E)��җ#���=�m��y}�3v�§��	ι2�f,	�����t�ss4���#nz�uŨ����r6����,nN�m���)��|��S�u�������h(A��f�1��Kne�2tvmK�fH�i�n2�:!���P]���
�~�cGd2V�MJ�Kg����� ���, ������>���z�«�r�� ;�*^���=��=�v�i�_6n�OUB������ �w���8�}w��x@k�T���Q��*X;�[,�����`��b�?s�� ��v`Q��$��U�#�`�EH느z��s�q���#�7�ۈ��n5�Ω*q��r�t][)έ=�u�m���&٨;x�w�� 6�� ;z��� �ʵ6ªY,R0r���ٜK~����>���ێ����TT�'o�|@M��@w\T��U�<�.�uJ��mYl�8����-�a��o��b�:��������SR�uف絛]yx@k�T��nq����x縀��~���+*vF��� ���,�J#�Dv�ޟ�����w�Z�8�q�a��l4zn�-��]-�c&��x��t�j&佳��{��>n�]l�Xlti�\��ٰ8��M��ze��IB��w}� �����K~t
�����DB�P�d��֬��Ձ��d��l47���8R1WT�Y�n��,$���M�T��)
���Z�\�<�M��sf�:|2G,	����Ұԡ?���`|��6�ɰ���t���D)�
�d�H�ʰ�������@�_� ;�*@;���ۯV��8����b���<����b^n�w���!����5|�N�8 ��s�m�� w ;�*@v�N ;:7�#�5(WQ-�{׸�����b�8��L��vg�g����^QYYaep��R\�od�?]�� $��X{ݪ�Q��Z������z`>�́�ze�B��d���!T*P�\%����v��+��H��&���)�M���rl$�/f���w7֬ϛ� �&�,ER�4�n'�e���|#[�Qxf�Uq���ȳuKdz�/a��~�;Q�RG
F*�c�����X;�� ���=����� i�^�`KkhL��@k�R�}_]�o�� s���EK�$�w��l�eT�X�*�8��L �&#�UWnCʐ{ʐ�eݩj�r7M�����J"!yD%3��U����Xw2Շ�G�S��zl��%�s4�h)�5UV�閬DB�^�7��|�}�ʰ-Z���؅�!'�sZ�t�y��Dic!<AtČa�A�b,bX�a��x%tH��B}�3Q���	��'*`�6"��*�`��a3�h�oT��';t���Q�W@g,���/� !�t��	1ØD>��3ޓ��8����:���v�-�msgc%�Zv�O�J����6���NU���֫��D��QS���:t����+�����$8;k��v�us��F4݊�8�r�{gZ)�j^�]V6u6��.j�Z� 4&�������r���L9���:s;0C;�ИS#�2�&v��M�ꪭ�e۔���JK�� ��e^�U6U�]AvE!�N�Z�a�cM0�$�ܡn�t�#q93;UU��P�]�j��Jl,&�"�-ku ����`K�!t��jmns݋�UgYpC]W�b�Aq������+i��km�ū��g�l������f�j��i$���\���r�7UE� 	Ulb�w�b����t�Z���������:M]�;[�Af�D��"������6�p;FF�K�l�KsϑS0n�G4�X��c��ֺA[#X�5�"X8�(Y�٤tZ�7�eغ^�A�y!�����(cUT�eu���'�9�`� nl�g��k�:X�v�RX�g`���K��h��\�BV���q�3������\��vm��
�7a�H�Rr�/m�6���@P�QPTi�/&�����DO*��A�ŘU�+��n�l��R�s;��u��xùK�FC��]ɞ����;v�v�fe���;\��	oJ�H҆f\aG���[v�2C1�N�I҆�8��<��m�6k�2�l�@�E��r-�#���ֻ 5��֨^�"wSU/;p��Z���G}l��7lFj��˼y��+��*��f.j�[s��l5l�V����%1UiKt(���6�];J�����.��v��ԥ�"���j���v��gh�j�dѱ`2����ނ�#DqJv���{m���f���K��m*�gl&�0v�&��
�ͣ����=j���n�ڛ��˳p���m��� Ft��i��p�m�5��a���m�!��RˌX[%l�S�5���r�7i!T j��g9�3�cm�R��U6��)|��<?-ن�ry8'�E�7b�PJ�/D_�=��w}���������0"B9��[���M�ɋ��'6�A����U�c����:Huż���!Żeu�ݘ�WX��R��x�cF�l˲]��8�&�6��cj�x�-��C��A�S���{�V�g��T����,��>y��퐝��X9�̵UH��K]��`��drPJ�^���Ӝ�ڑ+�C�۝��	9^m�+#���R�q��V�.�.�}�U�&C�&u775�.n%�[���d�̽�L����.Rz�]�T�e�`�佷?;����Ȫ���YEi*����N���[�>�j�ݓuҠ�N�*��&iX�{��QЦC�����ְ����|�=�O�#�N�vW�c�l��
��G�&{���rw��:��ؤ�*F*��`y$��� �smX�{��aBy=͛ 頷dr�MT���*��ܵ`lB�����>���]0�u��l��*#�&ö)4����`��7�u�]Jݺ�l��������}�Y�&̬��K �_�����:��M�ϰ�=�D/�;���w}j�f)�31-Ͷg��r���@!�ʥT�P(�R"5�T1�I;>P��j_Y�ºX����9�����d�y��j\�	��T�T��=j��w-Y�����1�6l�S܎ETVV:�+IV�O��~X�o������O���� uR��8��p�2�x�=�N9�t�~T��{� ��5�1��Q�5+�� ݬ�E����r�;�"J盋�K�k;^�r��t��x��Z޹�츩���}�l7�|�[<z)$����6If�m�H� ��@;�8��������刚�m��+��Z�;���.��E��(x ����jI���F��u�l�t����$�iXz��
w/|�y������S��*3v���B�n��k�8��@��k����{�N��9�dz���Ij�
���5�:;QiRV��z�:Q�z�����]p���&�+	B�Wm�{��X����;��~�/�5�}0uM�r*���Xa�/�H�/]��z�����Y����
�H�VU�of����#�m�����T��*����^H���v'��`}�6Ձ��Z��@�� ����E� XX�r:~C��7��IØ;�1�5D�UH�3S`s�2Ձ��sx�vo�����9�{�杲�k�-Y�sq�G$خו�RF\�I�a��>g�u˲������\��D�6��J���� �'q�w'bIq���mX��)�i�����$�iX�{��/B�
&My����֬gr��BJ!�3v��ʠ�F�TӰ1�6l��-Y�
�sq`��<�5ks���ʋlv�P�?��x��6Ձߧ1�lD<��́ީ��ETVVP��9V�{��$��r����}6>ǖ��)�C����B
9��Ƀ��.L��Lf@B�OLF��iݨ�M���ll�	ҶM�T�gv�Q��=;��u�ty��n���/C9�ֹgf�I(�Iz�gCڔ��Q���D;k�lq�����YS4#4,�/f{h���µ���}�Y�ƈ�N.;�a�)��]�{n9�.S��v6�ӝ��]2ny�!4�Y�F���6~s+#���vݎqU���"��V�rs]9'��Ϟ�{���x�_I�ۄ"DM�t��*�v��c"2/9��'a�Q�tOm<p� ���3*-	H�VU�;�� ��v`����9��,����(���hz���c��x�]��/z'#�#�l�����X������f���}p�զ�F"[�Va̤c��x��bv\ŀ��f�ꥲ�9V�N��?"#ӹ��������ܵ`u>�y8涹��e��:����[�;k��E��a�b]�Q��y[�#R*�u�Y_��ݗ ;U��|���y���⬌���l�9�{�;?4$�!BY	w{�~�Z�>�����ߢ"|���7�ȬVVTK)� �ذ�r���\���_� %��p�/8r�Z�$��}�I�n���}0s^��������{�^���*�����8�ݗ ;$T�{�- ��o��M\�7i.������Gn�M���Nċ��y��[s��+j�Ӿ]��¯Y7S�/��O��R�EH�r��l%�� ��^$R1�GҹV�wqg��Q
<�M��;^����yj�6f9M���Ke�r�{7� ��va�ҤR1�|t�W����_hԓ��jC���cj5B�n��k����w� �u���j�a(O;Y�����ͺ�qVGX[e�`�ŀ{�����~{7� ��v`�S[g͞~��Z��7U�l6�P��9+���ô�=X�m�Lu4�z�lrR*�*%��U�{}� �'u�w'С(��^ڰ5��RU��%U*�f��ߧ��b!D&�}͛�׶�gr��%��&O{O]H:��������M��ǖ�ԒP�ۻj��m�uv-؜��V���0<���ۯx��vՁ����b)BH�HP�M��>��D>�5���$�=��1���G̤ٗd��y%��8+��>ǜ\�m�DFa�mL�f[�UJ&S@t���u�vgg
.{\d��]�ֹ��ٮ�덯�{�!㏗7Z��8n������>���<�Sm���<�؈_}-���E�����mKTH�6ʚ|�m�̵7��e���x���{�t[m��Y���BK�U��?&W�$mS7? ������\m���E���S3����6޽�Sm��\W�\t��ʉe#�~���������R�m�ku󍷏2��m�}�8����Ov
��nR����m���ߛo�/����6����.q��v���۵	  GA�4>�Nc�B�g9Ű��~�/�e6���p�mnɳ<T\�`A'Y����If
�R��&�8��̜�W)�yڙ���0ts�c�GBs�� �.Q\,���`�N��.ںG���<�&88�vmҘ6+��׶{=%�uz�9�`�C�g;t��N���·�e"��7:n�V ��n��hl*�m��ʲ�b-t����K-vww�����_Y
Q�ś�ܶ[2\lѲ�۵Vxm��oO']l��$�no��w��3)¨:�_��m���Sm�:���m������Dre�����6ަ�_7#�	��lr�����7�����RK{���re��y󍷯6�ޥ2��]��"��-(RU��m����m��Vc��DD��͵6�o{��s��>��i�V��X�#��m�}�R{��?ߛom���y�L��~��IUg��v�o7~w��mE�L}} ���~ ����/�m�ݭ�m����|�m�'Sp ����tj��3�x�.�5��8��7m��Q�^��z2F�5��m����6��+)�m����K亮�}�cm�����JE]e#���~��w�繺�)��w!<����
}���w��m�y�Sm���.sTBS2��o��87)Q�-x�oݾ����������Q�EU{w�\�m��z����t�ԄaT��������o{���m����(Jg{{��m�Y(�ne�A1N�c�Sm���.q��D$��{O����������Z�m�����������j74�C�� �Cv�9
n,VxW�]Z������X�*�E#ZR�K�m�ki�m���8�}}�S�%
#������ﯠ~~~κ��9J������|�m��-M����8���ee;��B����6כjZ��tK��SO�m�_~э[m�9ݛ���P:�D&
��a��C�I�2U@0�W��X-XHH��2���20&�a��rf���D�%)`SC� �`�XB#�1��;-ؘ�F�0��ξ��j%bu�����`@XO��HD����7��¢Yʣ��<b$�]	�t�4(l�t��`5��(�D�d?*P�a�ĉ�����P�Ԋ A�W�%@~U*qt�T_?!�_
/���3�n���o��~m�]����⬎�HKT���$����˜m�ݭ�m��+1����1�����qVU`냵~��o�YN�m�r�_�6�<�Sm��38���|����[-��CDtLU߬�Gd�Y؅�+ �6��Ҹ&��/l���u���E�R(�m�_��~����ͷ���1���g�B^�	w��y��;m�����r:e)��|�m��-M������m�����ef>sbL���+[�rPLS�l�ɍ[m�{�ݶ߻����Ȋ�F*���zy��׾�6�m�.�d�r���B�sK�m�P����Ӷ�{;�<�m��1�oPTЄ9��~7�m��\Oj�R[$v׍��m��6ߒ�哛�<m�����6��+)�m�-�f4��ۻq���d:�t��ݎzYb^��q�uϷQ�^{��+�|���!���[o^���m�����6��+)ꈈ��o���������郑�YN��������8�o쬧m���������Z�����ʇ�~~ �Ѯ.!�w��ݭ�m�����ǰ�BS3�6��m���.q��Y��!�nh�*Snj�����DB���>q���M���{�\�m�������wG�X��/������}}�Sm�����Wz�o=^�m��������(W	�8�7�OF0��Q.�h���cb ��'=���Y����ڴ��W�9P�6ݻU���t_�����`���3�)ٓ��#��;���WX�[�v��kb٘L��x������r^�n�˔�L�[�y�4���9"8��	�xm��;x#Bp�nܝr���%	ڞ=�\�/��Ͷ�v��c&�Z,)��'u=dv
�l,���C\�NԖ����@]
9���3n3I��&.1���O�;?0M�U�dUs�:��B��Z�u��;^�����D�2���E���� ��~��w��ͻ^6������m��qLm��}��dN0&�����m����aDL�{=ݞq���ڛm���qs��B��<� ��UB���$˪�m��{�<�m��-M��z"*�۾��m�����v�6ԵE:*G$u�?~m���)���������|۵�o�O^�������ߦGdu:BZ��m�{�\�m���>6��������1�=�k���Z�U�����(�6ܑ9v9eI��^�*�p�Z�������uH0�eN����ߛl��.6������m�wr��۾ŀs����T��EM�n���w��>W"���
��H"$�Ȅ�^��ݿ�X��Հs3+ �zn+e�:�f��q`���&�{޸�����4�8P�[ʻ/�H;WU��b޻����V�{�H8���>�U��v��s��T��qR��U}U�%��~�5�e�c�b�5��\ch��7�a��F�v��ۢ�ó̐�qLnJy�U���縀m�H�~큾���2�˵�t����{�ŀ~��, ��� ��v`�٣��YN���$�y��M��Φ�ҔE�TaQL��d&�
8�p��Io���{��;��,��wH�uVUC�y��R ��� qR^�{��o���EVG)Q6�_;� �,��.�͵`�ʰJK�%6���tv^�9ΰ�:���.v�="�8�.��7��k;^�B�F�������{��grՀw��򄗔/�5��l����u$��69�`s;��TBl#��-�q��H����������V߳*��g����}��V=�b�:��'���v�	l��|�O2�]��͵`s3-Xq%
aZ�D$��|�ٝ�� �ڶ6�T��Hݖ�T����Wվ��] ���|r�λT��$���P�[c+n�2��\���]�2S4lХ�5q�����w�޺�~a\U���	j�=�b��v�����þ�b�5uM���ʪ%�9V w�ʽQ
#ВQ&���Z�9����z!D%2n�ñRu-��Js3U`{���@nȩ�"��& 6HZN��Mԉ�L�S���(I)���V}�Z��̫B^Q	D�����n�Ø�B}]M�*�?n�, �7n���ԓ���lV�a )�p�Dr�0&W5�F5!���0�������v.Ӊ��0�7UJ�(V�	d��� $�s���<�ig�W&�Ո^j� �yb��	'�.zKG]��d@,H�n9��:�qW���Nc�������;e����u#�nሹvͻ)&���ًvr�m.�1�.�m��� :-�u��8��m����i2nܠGb�Ö�(�p��'7��ɛ����>U�ou�Ƴq���gY�k]N�::��aNە�qp���S�1ۇneg]V��
U6*�L�J	�D�����b�9h� ;$T���|U��mK��$�MU���q��(�S&g�j���V�ٕ{�f�R�mKTN�s�]�2��ʐ�*@�b�9h�F�4�VGS��Ձ���� ;�ڰ;��;(���wx�]�4ni�YU	]�U����;��x9�� �����v=Bdj��KS���gm�j�-�c"2/��؜	�y�{h]��M����>k��"�'$���|�sw�wqyB�0;�ڰ;���Q%Su"t5Uu$���F����B�uA;�ꯛ9����b�9k�]����	�mʰ{�ŀ����7�7� �}�X��wT�'Ĵ�4�*�؈Q��wj�ܜ�`}�e�P��w� �����IlP��p��R�wx��vՀ}�eX�"y��;{�ۮل���i˜�vפu�)�u*"nӈtݻ]߯��ru��Bc�m�~�� �1�����9!du:H�X�wy6�pl�<��ŞM��^NYUeU�\��;�ڰ3��vuE��8HH���:�D��}��o���I>�1;(KsD�R���Xj�	y)����~��6EHvL@k�e��y¯���@nȩ����] o������[��~���������/E����F�v;eqKL�n���<V֏�m|�	�mʸ��b�sv����
q�{�j���T�$�5E4�*iX�fU�^Jd�������>̵���:��g��R�%���7�����VlDB�DL�=�V��U����F�j������|�{�~X��b�$���:� �C%jR��|��B�|��;���X�T�t�U3J�3�ʰ=	B��
s=��l�n��?'��C5�mR:���[ZS���7i�� J��E�m��R����5���UTv;e��n���׀s��������{}���nR(�rKp��j��^�2f{֬��U�}�e_�P��^�j���:IV��ذ��U���;�ڰ33mX��3$����a����`��X��B�>�������I���i�� 7d�n*@nȩ M����eU
m*Bf�"IQa0!�H$Te�	ď	�z�Z�H���3�f�NHt`IIHB����i5�f�`Ǥ�����1H�$E��C`D! "k��pd9ě�.��t@SRJ�b+(4Z]4@�'��ő2���Lg#�t�
��@�G�2т#��� �H3�͈L�!0Um�p�Y�� � $� ���UmU\vT�p�6E�v�M��av�@yra	Ơs4��e"�st�bxy��T\z����ۭ�V��]�c�YÑgn�a����1�睹5���q��3�lkEr��T[e��0��Y�W�˨���h�8�i�lTg���9��"@�$X`�A�v��Mz��f�s�]6����D�LB�(�"�-m�ډj�g,�AsM�۶�:�ޝ+��Dd6j�cS%�;t�N����L�f�j�M��W�C�gu������/OL����)�5ǄkLp�=�`�YR�5&F��0����W���O�cS���;;m�R�H��ٮ@���.��@M��bۃ�W�1�Ҁ�t�Π�;Jk�9��P˘��](
K\v�t]��u�#d��w"�aNMڠ7
���+n�2b�TJP�Yv��[ ��Z��=^g�K����՝�t�Tc��<�T�J�E+�e�Ɔ�vD���t�e1�����RZv��D�QEM�u�T6{l܀�5�մ����k�.����홎©M9\�ܝ��Mi#2x�N�b��On&�!�f�em-�\)ơ�fr��Y�v���
��:�
ώ:���g�^!��nk;E0@��]����jݬ�++$�Ҍ원!)���m�[qm>I��
�7hjT����j����d��#ev��c�Ix�u��[a�����u���=M�� �/r�)�qNa�%��7�=��t���<c�cl�C,�;v�l�ٲiM,[3�ckm���0�4�f��[eT��tq�N�:��l3������F��-���n���Q�U�,������\�O��O;G;m���*�6�N�7U,u�Ů9-�
Ipnn4�̭�eV�ָgk�\s΂)��q�8�x�n^gvY��gjݦ9��E�TDᶛaV��؞�V�R�g���j�Y�)Ԣnv�Gd�L�2�-�o���8�"=z��@Qx�*@6��ڊ<z�P>��7��G�"!q��TԢj���T��6ͳP6�޽����%�K�Q�҇\6��];�<�m��عιZ�1��mH$紐V�`�2�ɱm8ST	3��z�p�:t�6]]h����cv	�ڜ�e_\p:3�Ӷ�zC�W�\ѧhv�g7k��5`g��mds{�mګ<�/���q��;^�ӺI�������c
���Z��r0�F�Z��EPٹ�o�3�L\8���.1�"�e�cXg�\��������\�x�����o�{>h�U��ؙ-��{�ŀs���>̯B��@������^�ԵAT�G<���)�"�6L@�b7/�B��;�����uI�I�*�f��w߿b ݓ���"��fJ�s2*�,nYn�ɾ�޸�}� �7q`y}�|��po�2}S��H���-X�rՁ�
;��. }��`}�X8u��K-nPN���R+l���^�v�����My:�#��v©
�K��F)V�)J����.��ڰ�2��+�a��j��"^h����`�4���W0�
-$�$��B��߹ʰ;�ZX��, ��9�J�T�� �$���#�Wm�ʐ~� 7x�,ڬ���n�����<`ｋ 9�ہ��ɾ�޸�j�mF�Z��9� 7dT���m�����@n̂���4�\R�i��+ct�gͷ��n2�Ld����F�k��Q���L�F����2�였7d���~�U��$��ŀ//�����]c���[���(��;ݭ,�vՀs�ʿDBl�ݜ�T�nR(�rKp�o���ł_.�DDE&���B��g.��fU��.�Bt���6�P�}���w��`}�VI$�ݽ,���L�PL����}�eXJ!����;ݭ,sw wN��l���%�J���u�b�Y���V!Pݮ2 �͊x�]W��6ƮT~!iZj�ۀ���9ͺ`��/%����� �f�=lmKlA-��� �W���p���HO߱ nɈ�[Q��$	i�s����ݸyB��3=�3=^,��1d˪T�j)j�U���o��� w���9��0�PY%	�ds�(���D�XV.\DC�w�8�i�x����?����H튺�Ur� �7q��� ;�*@�\�8g>��w"<k��9qզ�!��)���\CJܗ�uUG�d<�µ�m����@nȩݑR ݓ�Aaft�����-_���3=�V|�$�3=�;ݭ,���K��	�Pg2��*@�b?}v߳��yR �YՎ[�$�TӇ3J�ДC}��X�< 7dT��U[~�i ��fr�9�R�j�����,(������� ��ʰ&#�,JF+�((sS=5�[��j��#RpF*㎨��v��ח!��۞��e&LRA�Ֆ;bi�|vF^Q6s˳�Y,p��J�w��STn�]0��"�[m�v���R�b�Sl��m�K��U��)�1�&��qXM۩8�:���F�O3�Ac��<�����ۮu���e��� r����V�v�@�[�7B8�nN���b��~�g��}�?41q���lv7s�]pBq�V�n�W
)ؗ�7k�uϵ��)\�XڍP��9 KMw�ŀnȩ nɞ����7���ne��r�*����V�n��sv���0�k�(�(J&O-^��jeS�:TT�2��{� 7fA��nL�vEHvu(��Q�C�}�O��� ����ݑR q�@7*qQ��s+>����`�q������v�==�א�;��-�*�ZI$#�?����LR�)٫K�lv����秖vY�v6�۱7dCY����t~� 㘀�y�U�v�zg� ��y���%U��*��v�R�U	eQ�ʲ��ea`s��W���"d�������ӕ؂[-�7}���vEH�1 �ʜ��]`f^p�s�����������*@9��t�?>��v�Ua*)h�������nmp�+K������n5�67C��H��Rk���i/+*��Y��k��W���f佷=ۚȲ�F+�����؀�y�!���k�� 6{9�UJ��T���n�w�L�7-Xs�W��L��/M��
��n�[���{���jI�����E�Z5 $Qv�S���;��I�s=��sBkߣ�'�V� ?sv�w�ps�L=�� �F��n"���/3�bu�<� �Ɉ7���}�q#���;��!d�N �T��n�.��=���V�vy�F��fs1��A wd�ݰ'�� �ڽQ���$	i�w{t�였s� ��匘s��2���0��vL@9�א@8�LWCj�$�*�,�K-��_7�ݫ�����v����	����%�ɼ��5��A�Q�T�[�s��`�	%�}����zՀw;�`}���g%�x3���Wqvz�����H��V����s��n�Zi��Q�RkH�s�Z�"� ���s< ���u�������ŀ���9��0����6��E�����]��R ����� 㖀�ȩ�ц3*���J	���B�(���};�`s��V�ICy��`fe-�b�Z�*�@��vw^��\��~�N��Τ��;�RL��cB��{�}���}�w��D߂sM�VZ����e$��ś�i���Q���p"Kvʴp�+�/2��k���������X6�s+U�=�ĬZCI-+�N���ۤ�nص�`�\!W��2��Q���V�����=��˴C�<�2�0䌓pώ4]yy9JݻP�u� ��6��j����+۱j�ʜ\��K#���U9��UMF�9C�enR�������>�� ݾ�����lZ{'���*�IHv�.A��F3%R��2l�m�z���Du�ɢ�0�/�� �*@9��U�����o��������lU�Y[�U���_�f�m�6s]��fZ�DBl��C�%Q(�In��b�;�����, ��n��&!J�c�$� 㖀�"� 㘃�W��=�@?-����
�++�7����ݸn*@9�-ݗ��,�y���$*WS�:"��c�$���Gf�1�6-��6�5�c�!A6;%\�r�&�4�3K�����T�s�Z �& ��Y�y��f3�Lg8�u$�9���`E���	�J��UR�{h��@9��vI2��b�Z�*�Fܫ �M���v���f�}pw}� ����5e�5 �e�	�b q�@MqR�U\�OZWV��l�"��V�`w�p/���\6s]�g�ʰ6v�vP"dt�����uA�uu=�c�����J�瞺'���+#R�eAB�u��$����b�;��v�w+R�\`f�Ձ�ճh����:[^ݝ׀����v��ݘ5Wl�8P�XY^���Τ���s�����>��1`$ �R$X~���!�mH�HFB�0��6;XP	��f!0�bbO�Q�0$��HO���&-���	0S���e(!a� B)A
�$PadF c��� �o��#H�$�P���2����q�c�a滰�,X�@"R�p"��%�#�	�0��$�I�z��1�BP�yن���(B���>:nt^�:D��BO�0�B�ؠd�:���G�����D8�/�QE�(��ސh�����I;�s^ ~Z�kdn"�ӱ�p=��$��� s؀s�Z l��|�`�m���n ~�v���x��ۀ���5=C}�㊪��Z��;�-�f�'t5�6�5+GNdDM�����w5n�Z�*�Jݷ ������� ��n ~�v��\�F��&���u�^���'�� k���r��G�l��R�����ۦ ~�v���x��ۀo;G������o0@K�8�s�Z �� گ��������}TJp�� �q!
�F �D�Ni]k���'��l�T�J�n��ـwgu��p�n��wf������*u��V�|�2p�=�=�I��U76B�hM殇��+��mu����� {��w{t��ݸvw^ ~\z5�7	V]]�̤� �;�b�9hu���_6kѣȞ��KlL��`;=�8�똀q�^T��+8�e�I%nہ�{�x�������I����;����+PvYH<̴�s<� 8�qB"����2 �D{���~�^�㣙��7`flT.�OmuΧJ����u-�نʋ����뎭���� zz��t�b�� V���m��mtvD��u˗!�5Xђx;gm��R����y������ۮ3��agaX�y6x��9�'��pv�q�nV6�
�v�a�=��7&��m֔yZv��ˮʅqY��C�� RAr�l����Q���c���ٹV�������w���������'b�]')�m��q�nxn
�@J�t\�t��,�N�;�|�|�-=�ns)�����;�b�9�a�yR�l<�(�N*ꭻL ����;���}ܵ`w;X^�K�L��/J�H��t�AS3U`o�|�}ܵg�!(�o7+� s��sz�6J�	����j򄧹��X�ϻ�`w'���,�c��%�*i��+�����(����};�`s�� ��#�2������E68h:ܳ�R
.{^9��y�u�g���~���a�J�Yb� ~�v���;�w-yD(�0������-�R�V�ʤ��m�;���|�>"IBa��P��������s�Ϧ��v��c��PvYR��ܑRǐG���n{ܞ��Dɒ[j��\�U���۞0���ݞ�����X��5�hn��N�6��& ?}S�=}�yRǐ@o���f$����@e�V+2v(��n�X�(-�^N�GdH�N�u��-����l�9��s�Z�"��!����� ;��evB��������ŀw{t�s�p�����è�đ��iSM�4�ܭ,ﻕcQ�)�
�"�" ��y�o�RM���ԇ_D֧�J�Yb� s�ۀwgq��2Շ���������]J�UL�T�V�vw^�\��~}�� s�ۀn�bln���O���f����x�.V�-�H��x��m�]�mL>9z��7/A�dMH;k�?sw��� 9���;���]ѻ�Kej���\� �y�� 㖀�ȩ{类��\�&�#��]U�i������x�n��;��`�[1�E*�жKp8�;�*@8�;��W�:=_e���hyr��wﳬ�I�xϳ����>9Y�9���ȩ �� �1ݝ׀y}�O}��,�K-M�nGeꨎ����LJ�kgGJ���q�v���"#�*�$���0����;� ���X_D֧�J�Yb� n��8�&�� ��.��������MH�p�P7�|��P9�^��wn��>��Ee�5 � ��� �&���A)�2]��(�jYV�ۦ o;� �v�jI߹��)�yi���iU&��_%;��[k�`��BR6V*[Lp8Z��ݷ���O\1�t[�N�u�8t��l��y)k�H)A��;g�AkqK��u��4;NOE�F�zt����`�8�&��22>c#+0g&��f�įl�D�4T�n�{H:�����t�\��N$���u�X��.��y�YV0ʷ��+�8絕�q��ju�-n95��a�ж�܍��L�ط>I<��"��!QN}b���N�k.9[��5�<���gڭ��Ur^��	��.��˻�:�L@72	�*@l���ճ(�t�V:�n��� ��ɐ@\�ﾻ�g�3.�(O���� �wذwn�{��w}p﯌ �4����P�r�$������<��d\T��Қ���PK,AIi����9ݺ`��,�;��/�Kg���;j��cv���;<���Y�Xz�T��b^�ݯn�>�C�Aʬv+���$�����o;�������v�ȟ\�"��ȩ�Is��'~�tj�� �n �Wj��QR �L@w^A)�0��-MV:�Rʰ�����v���;�ŀ{��X�5�J�*�9V Ms� &��W�느Iǔ�8B�d� ���X� �;��yݸ��w=k%j0Eu�<������屨��9jE;������6��ngכ�����
�+$�p���,�����v���� 8�;��DGiX9��Ru�Hk���qRk��}Z��h�ʰyݸ�n���S����R
�
Z2��W{�3��o���I>�2w�����%-��>w���w}� �;��yݸ�'�5H��&�	2�\T��*��� �=�� �F����rT�E������S�c�ʪ/m<�tq��"���nK�s�I��Y�U�2�� 	�b��}]��K 裏�Ԥu8����X����_(l�����m��w-^���fn�N��
�t-����b�7��X$��wذ��\{�l�X�	�n�@MqR��5�@��Gʾ��Uwn{� 5o�$��Шr9V���Hk��5�H�Ng.�9o-tU��W.��e�*^��L�.��=�G��+\;<ɸ늠33�@��m���느\U��k�T�~�^�s*�Z�*�R�p�����w}� ���, �wn6obz甊�"j@�)�<��qR?W���vy�b\���)6Wk
�K���;��>�U�ϻ��5$��7��ܝzƦ�j�V^V_/�Hk��5�H���Ԓ��p �N��X��HDo�cp��x��Ap��@`�D �t|�Ѽ��$ᣋ�1�%��F,F��=S��#����� d"!&�`p�a
U�J��  A�=:0��"�#E.��:�\�c# ���~ ):��Kze2� �ГYb����H20�D� ������kd$ �O��!�D�8P�K(H��/ h�5��2�J1Gbv����ڟ!��J�7��dC�I�g%�9�sB��f��I��'Ce;um�9��@\�@1�]8��� �p��Ku%��bF���� ;*�xy���)�:��g��c�k��P�3uz-D�i{j�����whDzi�yh+2����K)7k
JA�ׇ����6aAHZ���xVl�.ݧvٮ��b���u;� .��Lʹ����/*��wh
V
K-���Uy���)*�eZ��d�f2e]��wX�WfU��V�K�f�á��I��-�X�v����=�msn�j�z����69T3�eBȅ�ֳvV�q�-�H� x j���\���%��Ӷu�9��u�tS@J�vGj��y�ʠ5R��C�y

�E[Z�Si�spR]�Vlˬ+�H�y9�.���Ʊ[�:�qW8��;p/��q�*մ�(��\�<c$�G]]�NA�K�]X]g�l��t�Z�'��┖�L�4Ub%	4p'LcS�P++8� q"��U-��
��78�r�ўq�ڴ�:�@ՂNv�8j�:x��<�-�pu���2L��XT��!$S)Y�h�OEn��Y�㍙C5��U\� �vD���mS�Got�ns�d��XV�)��J[��Qf�N�Р++<U2��ĵ*�@�;s�x,�
ӎ{9��1Y��iT�U�b7"9vZ�v��-"�L[z�>3�1^Z��%8��Y�u��1�Y�M��r ���<a½l�s!�X�3�{cd\�ܝ>��$�d'9^��۷l���UV�8Ԩ:�Q�ݹ6{)�z�ڱ��>��	�6C/[URV]h��@��.� �"���S�"��Cǥ�'�����6v��	ékGX&�B^:.+#.�t�nL%915KtAE���ڽ��x��V�I�l!ԯ,�q=i�ٸYj�)m�������2I�����CR���c	���z�୶��J���w{ۨ��E2�p��6U��u����0P>Gb�|�iTn�	�6.�7�;�-�O\���;[E��i���a�q�1��
��t�5u�e�t��h��Bpj=���Jl��u�1�m=�91R�:��ts���l��Н���83�g+y�,ҩ���b�������6Ѷm��4D[�������Dn}��/M�N�i1z�idZ���zs�#m�6Fm���;v��R��t�9:�����KY^�M�gE�@������/��6�$p�qü��9�f�����U�^�.�z4Om.�N6�T$���]%�-6#qRk���z�`y�b��^�J�$(_��v�y�ŀ~�w o;� ���, �4�I�P�r�u�Hk��}U�޹�H9�H���������ܫ 7�ۀ~�w�������︰���%��k,�����느\T� Ms�������?8�qm�;'���*�z�;W ��1�%��5�dٮ۬�toa�q7��s+�y�*@w\T�&��������N��]�
�,Nʰ�qR�U}S��}�`c��� &������BTE]C�� �wn���H	�*@w\T�rU�ya���^g9��5�H느~�����ze����nՀo;����] ��u�Hn�]�p9��~�}�:�9l���lH�3���K����6-��X�5�G��$�-
�#�p￱`�1�qW��퇜� �u�=��Y\��U�w̤5�@w\T��qR�;��������%��k,�IKm�9��F���;�R�2�9E6q���ۋ ;�� ;���Pv; �$Ұ�%���>�V�߻�a���,�|��ҹXX셕`��ŀ\�[���*@m�ɟ��<r���U���:���55�F4 =+���vЮ�$R�|�y�	�A�E]E�����@u�����v�d���+�
B���l����Ş_/�g=�ŀ}����w*�	Bl�ֶn���J
�j��)��T��qR?UU�� 6O%�F��I BШn�f���Xs�w:�o��I��8��?�x߿r`��z��)e�(�X�wn��n9�[����r�9��eڈ�|X��kl۱;��(��c��
�t��X�V�S�k���k���r������>� ;q� :�U꯾��`G=���mT�Ӧ�LҰ8�7�Q�fm� ��Ձ��-^��z���|�L�J��T�Gl�;�b��p��7��b�8���wlz�%	QuJ��w*��{��<�M��%�Ow}�=�����!j�P�Kp����?ow���-X~�U��Qdth��5Oh�F������4!ue�k��l�=��c�PE�p�;v�b��"�Wd�v��-cV�7�-�X�������v������[�)�ugPn*�m+��4�h�k�;#u�jMg%�]`ㅶe吉�u�A�p�z#��n���=���b�F�ڝ� �`�]=s�p��8�[m�ꀛmTH���h�4[�V�_~����s4���Z��V����3�t��*i���/]���K��Ԓ�d!B�D۵h���ŀu�� Ms?�Wݰ�<� :<O�9��̣(�r����qR �� :�T��wqg��l:.�3��&[+AG*�9�@7"�~���T�~�� 6<�rZ�T�ʤ�����ŀo;��n�,/�o��\ ����qA��J�9����� 	�b� ?��$�����zX��:�N��L|��hm��,m7�@	�y���K�R���кef�]�3�y̮���*@\�r*�_v��}� ����hJ����U���̂�|�:Ms{�]�I;�;�R��XwV�+
B��l����>�Z�У�3���X�ޫ3ɜ��B���,� ��q`��X�ݸ{�� ?!oV��J��#�`$T�&Ɉ�T���H�|��T��8|�����*�r�㘛/<N����r�β�k
��Rt�r��1 ܊����EH�+\��*��%-� �wq`��,��� 7�ۀ8�v�(7]`H��MI;�;�RO���Ԥ��T`�W� �DB�\�s�~�ڰ1}ܒ�ԕ*�T�'eX7w o;� �wq`��,vu�m�BTE],�`�ȩ5�H�*@M%�|�s8�vs v{UZv�59g�&����xz��r$u��4zL��H馇k�����̊�\T��"�5�@HC&f���YV����ɳ��P���9��@1�]q��G*�?7 	�b� #qR e:vLtȧ5��+��7�ݫ3vՁ���������f��9��\�����9�s1 ܊����EHl���kbi���7���+
ʆ�a�ĉ9n!�����m���ja���n�5�����9����H�*@d�}_}]���b�<�}��ʡS��,� ��� 	�b� #qRN>rYu��9YyFs�Hl��nEH�T�����?wv��F��[p=���UUr{ݤ��� 	�bBm����YV����9���y�p�w��Iwj�H�u[Uu4k]l�5q:XF4�s�)�e'E���y��x�����Ÿ�5=]u�A�lO+u-�����ASIm�.�����p.h����s�W'�7J9u@l<󩕛��(�Hq���<.c�(�3���:هTlq�X��{c�J��������n��o%�XuӺ��@6�S�b����N.�l��s�;�0�0�X���V�nFa��ﻻ�Iv~��yS*��ݣ���zӗ���
��I�V;.m�j�w\j�	�dq�9QP�r���`�v��e�(�K�73mXͧLL�s>���1 ܊����f����j��b��U$�����,;ܵf�I��֖�ݫ �|���⃱�)��{�ŀsv��ۀw���]��#��S*u֥�`$T�&Ɉ�T���H�L�D��M�7=�v�;Q��˅[i�Z�7k��X��K�:�[[7g��-�6	�b� #qRd��rs����-Q������ō}�_�A>�
F�M��PƧy��ԓ��tjI;���%�ɳ�<_[Ia
� ���<��EHl��nEH�Tu9ˍ�G*����� =�z���,{�ŀ:f�_�d�2�U�d�r*@F�� =_}_WӞ7��ߛZch�ҝ.�2a�<cI�3���G�4K�m��ۮ}��ó��k���r����{ʐ���EHl��k����n�`�RJ��w����ۀ~��,W{���Tʬv)eX;�ŀ�ۆ-I*��#C���l@Đ� U��&�]ʟ p��}�M��������ra��jPڡPL�c �ԩ,�C|��U��D�!��h(}���4^@���d4�RԖP�at�jPή �h!dW{a4b}0����T2�����$��2D9�IG��WIS	�{u�N��!�� ��@��ͷ�o	Eh���z�T��S�^*��p{�A>E6:��^�b��4�h�-EO�":Q���ŀ~�w�;&�������y��&Ɉ� #qR[��{�<u�!j�Ul����� ��q`�w o7n͚�q���1� ��'�����������^�^h;@�K���j[*��~"*��}� �{��>̯G}����-ų,��T�2敁�{��b"��Xf�;�ŀ:f�_�l�rU��ۀuȩ5�Hn*@=�S���̬�*iL�UV�ٻ�`nfڰ>�r֤����� h�ȠD0��_y4�9�ٗ ��;6�݄�RW9̤n*@z��'�] ����"��f��	mU\�Z([dr��f���ʪ/ms�n4�[����Ƭ�l��]ju\�Y˼39����6L@uȩw�͚�Z�+abn� 7���D6wsmX��VW�X^��gsuL°�-Q������b�7������ޮ���o�p�֮�T���g2�ȩ �fA G& 68� ~F�Z�"!hT9$� ���0\����r*@]��UG.���]ݶ��t]Yg���+��[7h�x2���9�\�n���-��9ڠ)c�DG\�dP2#Ր1ŷ��@�����2�
��o�|7n�g�.sCT�	�r �Z�����i��zQ�2V�4I�[z��8����Z=Ǚ�c�6�qh.݉��vؘ����t��N�N:P�i��s=g���T��`3�nD��m����Ўn�ig����{����N����=��]��̸�//j�:�qr������6�vy6��F�j������ߞ��� &ȩ :�1����k��$�����,y�� :��p{ݸ�=sY�d�djIV6EH�Ɉ71��H	NN^�mP������ޮ�� =���ov���X_6jmZ�+am�s1 G& �b9 [& 7b;�4�;���?�� ��9s���y�/]�H=qm+Ó�>��Zt���S��c���EH�s=]�==�@s|Ӿ���~"��p��,i|��m"(�
T�{�&7��I7{� ;�ۀ��V��ZI- Q�@Ɉ��Wd�� ==�H�C��clV��#R[��_&������@G"� �d���2�*�Yd��� ��n��ŀ\ݸ�ݸ�# }��N�B?��rѶ�S�I�j5�.v��i�ٺ�r�]ۣx���*�6㥶���X��ۀ���0;���<�}�]t����;V u}�W�l7wj�;��`ffZ�P�f��/&�	Q���-�{޸��w:���d��� /�}�oF����pwuI��R��V�n�M��bޞT�;[& 	�v]����e�vۀn�q`��ۀ�� 9���?s�E����G'��4b���[�땶�ͫ�k����zذv�m�kjvuԒ!hQ�%_�8��\ �ݸ�wn��� ?�m��[kL�ՀffU�D(l;�ڰ7wmX>3*��{�b�N�Ye�Q�p����ܵfϺnՀn�Ձܖa�9$)M&ܺ&j�6=��+ ���Xgs:� �J0rSF�Mj���ƞRحcU��U��n� �L@�b9 ;��9�(/�����rpQGj�p���9nH x��Մ۴��V�R)+�S�%DV��	n owq nɈ�T�;���뒹�e�X�Q��v� �7n��ŀ�n� ��n��i���(_����y�j�9�Vj�
f�mX{�V�iծH�!hQ��X�����v�9�p<��{���[b�֙���������g@��� �&)'B�p�4T������"�H�A�5X��=�kS2ɋ�'3D��;%��t�e��^(��y	����]u���{/07vm��v�Vո��{#��ٞW:95$�u=h�1!���<km���s�V��j.�yRp��V�s<�J�&��<Wb��w, ;^'��8VɎy����<c�ݻP���z��Q��vsm(�&$-�u��mvU����~{���p]�[��朋!�ʚ�\�Y+���o�ww����S<<nz�L�N�N�k
.�`g�f�:��'dn�S��W+���+f���~~~��0{{����n��P���ͫ6Y����Sn:In��ŞK�aΞ��n��9�p[��,v�k��3�H�I�71 nɈ	�*@~|z�u[l%���� �6bl��t�rW8��Æer�+2���7d�� �& ����E�7juKm������;BIXڬ�	���v4�s���7���ۘ#���5�|r�y����T�;���#s�ۀF�Z䍡X��j��7ntڊ �:�	���"}އb��6I��T�}_W���iY�clVZ&G	n {}����7����ۀs����N�Ye�RK�vL@G"��$��������� U*c�$� �n���7m�g{�`}�V��1N&�cͩ��O"v+�]Ń�5�n6��%rM4���=t\�t��T��j��[�Zƫ),��:{� #s�+�&V�ۇ.p�/(�fp���@��޷�	�*@�v������!j�Uk��9�p��w�5:�E DA�� �@XE@"@ ��B�d���
#s>��s�$�;��I�����X�B�E����X���;ܫ��C}��X#LZ�e�*�����+�����{����v���, ���XȤ�Ps�>J(8n��e��P�T�׳�oL���˧:�K&��e�h�� ��� �7n��ŀ�n�����-V�Ye�RKpvL@G"��$�����]�ў���
�Lp����{ ~�p{�p�ݸ�kز�mV���9��@�L@ɈvLA�_W-D��H�)A`\��Z��W��V���=V*�v�L���7d�r*@�L@M>Ͽ�$���r��k1���g�4��7j�;W:�j艜��2Z�dMלVb ݓȩ wI3�}������:h�b�H��(� ����/�_}v�{�� �1 : ��.!X��j��7n o{� 9�ۀo7q`�-Z�lY/��;V ks였�"�t�Rd��9�Z�e�IIm�sv���X��5$��;�I  lNq(FX��鄉��D�>i��
X�V"v��0��(�Łv�V� Έ$��p��"�6�XS����! �S�F��mҏ��N�«�pT �&G샤4 ��I�`Q�Ї>]�U�c�sr_�ȠD)�*Ʊ�"9z�];��"�u�>@!'G�p�B�\�7��J�fj���UUR���vb����7Fp� k��l���퇵���\,.8���V�i0����m�h�ղ���[v���$�<���Jv��ޥT�C�1q�nǞѰ�'1�X�R YeK@�s����࡙u�v%�Z�Pm h:R2����!M�	cbv�L�&��-˓�om�������-��lM�7�,�+#�*��rF�YPe�sM��5�*,�:,�NG'Z(v`�0Pb�)�[pk1wKI6Ќ8�Z�R��-�#��x�8ݫ]�`�]��3:��l��b�0�8J	�S�,�2�``I3i6��*�w/XE�(6FSSmW�h�4J����wm�R�K����I�Z�P����U��b7#6��� ʻ�JUk�H=u�V�9�C<���*��.z<�m;��;(XīΆ�UL��aݧ��"�P������]@\u�7F��ȠZ�l4�7J�v�&aX�H2;��y4���yZ5!K7!�q2�J�[>ЀD�C��+��'B�r�9��:���1�?1�|��^̋�PR�	��&�胗���Fn��/��ƴk��&�[�� ���ѧq�(O)UWH	�I��O6ҲI�z�s<��q��;�ܠQ���+��6�U�J9ntT��9�"#r����5Tq�9��2��1�hr��,*j�$1zr�,�/+U�a.��p�[v[`�'`v;q	 c\K�P�A!vٸ5/n��8�t����u��WYC��gm{[:�A��۠��"�{j`<m�kP=\r��CT���cUf��\�"R٥��0���6��:鷘��[']D�;<�n�U<�Z��ka�	�l�8����L�ʧiD��V�ܡ�fZ�wd��*�.;p�
G:(W���%��*�I=���&��q��j���;��CtP�TY҆���nQ�̺�b=FY�pV1��:��6�4�%P��*�>h
 ,4b�1���vJ���@
�Y��#���ߖ��\(8tU��@�<���- � �G��vH&��*�DZ���G`�q�g8&Z6���LݫG]q7*@=pe���:��ב6�J���8{3��1���
�v��C�[M�m�Ka�n�4ky L��]�k���7h�Dj{{m��LD٢�J82k��rg=u��c����W\��!S���(�UV Vߛ���z�Y�\�䰯���h�Y8�"�r��A�:�2l� k5���n�F����n��������{Ӡ���\�<v8z�]��H����C��^k��k�����/X-��
�Lp��������, ��n��ـj�vE��b�����H�EH71-��� :��oU������r� ��n s��g�������nڰ9��3e0�J�.������& &ȩ�$T�#{p�:3f8�V_����y�� �*@��vL@l$���r���+��َ#����Ћ�UX�SX8r�Քm�s�ܐ���$�!X��j�?p��@ɈvL@G"��*T�38g�LLLg:�N�Δr�R4�D"4Se(�G`)Ka(�il(��=�*�߻���u�_�;�{�j�Z�,��[��z�ȩ w]�@Ɉ����8\��%5V�7x���ڰ�eXlDB���ڰ73e��uT��D�Bu9H��b �L@rb9 ���LX鑵��l�K��"r�V�s��'3���tk�e�ӵzMʒ��ʲ���y�91 uɈ�U�`k��@s}�&�!l��m��ݹ���77mX�ǵ`�ʽI�: ݷ.AS*	Rꪬy�6Ϻ�Ȅ�H�^�℡s�6���ܫ �3��"�+�� �ν��ݸ��� ��ـk�k-���ߚ��� �& 6��}\s�:�{�@�s�hf����#e!��Pl����=Z�\ܨsy�N[�k�n����ó��]]F�[<�@rb[��뼂 �L@l����@�T�
In��� �λ��gs*�9�ʰ?!nf�\�t�c�na�g8�n%�bX�s�^�Mı,K���t��bX�%���t��bX�B��ٸ\!2!2�+A�*t�J�˪.L��(J��>�z�,Kļ����n%�bX��}�i7İ6��%�8�T��>��\!2!2۫g�0�tMH�*���I��%�b_��gI��%�b{����q,K������n%�bX�wv�L��L����L��-Ln�Dv�]�L��*�eIȼ��l�ԣ��;i��pmy�ݵB;tk�������{��7��Ͻt��bX�'��צ�q,Kľ���&�X�%�~｝&�X�%�x�5l���*�Z���;��!2�v��I�~@8���%�����7ı,K�~��&�X�%��g޺M�d&Bd-���
�A4鈇N��\!X�%�}�{:Mı,K��{:M�dz��$/z��p�Bd&Bd.��p�&|��g�}���%��k,�JIn&�X�%�~｝&�X�%��g޺Mı,K�v��I��%�b_{����	��	����ږI!Ji1�D�gI��%�b{����q,K������n%�bX������Kı/�����Kı?)� �-������o{�������y+���[���IIF���&��1��@^Ƌ^{B��<�Ԯ�XM�6.iB�ݪ�=p������+��N��F��Ęִ�;��a]^Kr��M�lt���;e�`N����3Ix��˂��fU���O�u�9ݦ�w��VnL�b�� ����n��;�pܚi{=���:$�1;M+\�h�yى�=�b�a��Q�w#p�51����ӻO�o�����I9:5hܱCɂ�"��\�՝1�^vb�q��r�*t�4U6�n�������L��_g�����%�b_{�Γq,KĿw�Γq,K����]&�X�%��&}%�*t�J�˪.L��L��wj�r�8���%�~Γq,K���?�]&�X�%��;u��O�	���d,����0�tM)j�S����!2�߿gI��%�b{����q,K������n%�bX������K�L�����r
�PJ�UUp�Bd&Ab{����q,K������n%�bX������K�����Ls߿gI�!2!=G�/K��B�%��S�[�bX�'��צ�q,Kľ���&�X�%�~｝&�X�%��g޺W��ϓ>L�w�y�#M:���$
�o��F뇤�a�^��,s&n.i㭼��k�g��AR�&�0���&Bd&B{����Kı/�����Kı=���I��%�b}��zi7ı,N���h��U���)%���|��gɟ'�����:�#�C��Q5�����&�X�%��;u��Kı/��gI�!2!wi����RS&�rQSUpn%�bX��}��Kı>�n�4��c�D!���~���7ı,S���p�Bd&Bd-]͖�4�h�m��fs��&�X�%��;u��Kı/��gI��%�b_��gI��%�H[���L��L��J��*�J�1��n.s4��bX�%����7ı,?*�����}ı,O߳��I��%�b}��zi7ı,N{4�1LI���q�w[u�V�T9s��B��N5�u���#i;-&Ϫ�k ś�������"X�%���t��bX�'����7��	���;����
HL��O��U���.��p�~�K�T�T:Tꪭ7ı,O߳��I��%�b}��zi7ı,K�w��n%�bX���ٸ\!2!2�i�e�̢�r�M��7ı,O�ۯM&�X�%�}��:Mı�GQB�È��7�]���Kı=���I��%�H[=�,�i� eE��	��
ľ�}�&�X�%�~｝&�X�%��g��Mı,�LD�}7�i7�L��[�{�D�*�Tʚ��&��N%�b_��gI��%�b{�ﮓq,K��;5��Kı/��gI���3�ϖ����T�V"
'��-1a�ŪSD�T�5=1�7AB0�;7n��D�Z��4�r虪�\!2!2�f��Ȗ%�bs����n%�bX������O�b%�b^{���7ı,O�~ĮU:�*��2���p�Bd&Bd.���n�c���b_߿~Γq,Kļ����n%�bX��}��KĲ�ײު�ʧLt��*���!2�}��:Mı,K��{:Mı,K��}t��bX�'9ٯM&�X�#!wul��ӢjF�T���\!2=��Ls߿gI��%�b~��߮�q,K������n%�`~ �Q�0<���Z�j��F"a�D$�D�����n%�bX��y��K�T�T:TꪮL��L�����7ı,O�ۯM&�X�%�}��:Mı,K��{:Mı,K������v�9+�7|���6��m�j��0k�:���K�BVw#��M��mA����k"vq�s��r%�bX�����4��bX�%����7ı,K����7ı)v�]��	��	��{�4(���L���f�q,Kľ�}�&�X�%�~���&�X�%��g��Mı,K����I���qS,O~��d1s�8*�SS3D�U��	��	��}�U��	�bX��{��Kı>�n�4��bX�%����7ı,Nw7�ٷ�L�M�tL�\.�	��v�]��
ı,O�ۯM&�X�%�}��:Mı,�"�Ls����n%�bX����+�N���0�EUS�\!2!2��צ�q,K�������'�,Kļ���t��bX�'����7ı,J��C�$D9B��Ƿ���Z^n��&�v�r�b[�Zn:B[�Tػv���ҭ�g/��'��)l�sp2��6�&�`�/n�N�HJYK�Q����l�cdC����`�b�.�
ؖ�pipE0C=,�qݛ�\u���ً%E�����c6o7bu�\�{-��i��79h�瑓��ɺ�E(�puV�D,ql�#N듐l͊�R�U�Kr�	j�����{����}|~���t�rQ��S%��J���jn9[�C�=X�ۧ�ا1!ua�]JV��~�qı/���&�X�%�����7ı,O{=���D�K��u��\!2!2{���sMT��R泤�Kı>���&�X�%��g��Mı,K����I��%�b_{����!2!oC^�I()��t���&�X�%��g��Mı,K����I��%�b_{�Γq,K�����L��L��qks3(U$�SC��Mı,K����I��%�b_{�Γq,K�������bX�"~����.�	��Ӈ�̢R&�[T��Mı,K���t��bX�'�����Kı=�w��n%�bX�w�:�L��L�B]�<��eʥUU��a�x�5�m�v'q5�;k�͚Z٘��y��Eq�]=F�[5}w�n�m��?=즠�	�㝺D$�MD�FBd'��W�&Bd&B�Sǥ9�
X͖b��:Mı,K�Ͻt��L o�Ө��bk}�=t��bX�%�;��7ı,K����7�!2�{�+�N��)4R����.�
ı9�k��q,Kľ���&�X�%�~���&�X�%��g޺MıL��[ܶK5UU2��-�Ӹ\!1,K����&�X�%�~���&�X�%��g޺Mı,��N{���܄�L��Y�/O(m�:&�j��U7�X�%�~���&�X�%��@B?�k���%�bX�����I��%�b�wvnL��L��5���ꓥ5UD�O�_[�����ݢ��`ĵ<��z��t����H�Ѯ�tU}{���7���'�����7ı,O��c�I��%�b{����"Ϣb%�b^~��:MıL��OP���fIB�%��S�\!1,K����I��%�b{����Kı/�����Kı=���I����L���CYD�MT��uE��
ı,K�{��n%�bX��{��n%���O�#��!��O�
_� ��04(̩ԙ���0"?D�Q��>���a�&80W;R�I�Q�p}�a�U��U�3�fT'ˊ�RS�~ڮ��Mpv�9R
���|0A�G&���r���j��q�P�E���%1I� o�΁
|�"
4;vՋ��@�d��	6Qr ��J��� ~\�F?�)�t*\(�:�z ����]� �CǢv'9���7ı,Nw�^�Mı,K��8;T��Yd����~>L�3�ϓ���7ı,O{>��n%�bX�w�^�Mı,�1�~��&�X�#!f���nZ��4�K�f��p��L�����]&�X�%��{u��Kı/��gI��%�b_��gI��%��{�������zy��dݮ;ua#q�K��#uk����1���;g��z��i��&fq��&�X�%��{u��Kı/��gI��%�b_��gA�g�0Bd&B���w�&Bd&B�m�Y�T\���ŷ�Mı,K����&�X�%�~���&�X�%��g޺Mı,K����I���qS,N��?c�6�R5N�T�.�	�������Kı=���I��%�b}��zi7ı,K�{��n%�bX��=��e�S*)���&Bd&Bݭ�i��%�b}��zi7ı,K�{��n%�`i]/�<B`�,H$a �(�vE,
D�]A/���wx�n%�bX�����̒�RT�uSp�Bd&Bd/���Kı/��gI��%�b}�{��n%�bX�ǽ�i7ı,O������Mqs8��q��6y�%����"�^;^���9-�g9������{�Hm�8���}ı,K�����n%�bX�c��4��bX�'��{Mı,K��z\.�	��77���ʪeMN1��g:Mı,K�{�Ɠp�$q,O����4��bX�'=��I��%�b{���&�X�%�����6☓*i��D�U��	��	��wvnL�ı>�n�4��bX�'��l�n%�bX��{��n%�bX�=�b�nq����uU7�&Bg�!)!wu�����%�b~���4��bX�%���t��bX�'���Mı,K�j�nUM1Җ��p�Bd&Bd-��+Mı,K��{:Mı,K��}�&�X�%��{u��Kı+�RDB P�n<S��J���u3J���'S��p�-�̡sn�N�q�r�I�jtݞ��s��K�и ����/l��DlN��ؒ�eU38ݞ3�c��[�u���%-��U�P¡e�vF$��6ػ+u��dS\Z,!ĺ`�������{\�c�y�[S���r���94���ͳ;�b�x]u١����	��f��-��d���7n��-Ӷ�pkVI�]{���{���G�ҩ#N$❇U��ۖ�W�� �M[5����uӯl��7@�R4�I�]��&Bd&B���7�,K��=�cI��%�b}��zh?��O�b%�b~���4��bX�'�<��ː�TS�T�M��	��	��ﱤ�Kı>�n�4��bX�'��l�n%�bX�c��4���QRBd-S�<L�(U!%IC���� �,N{�_��q,K����Mı,K�{�Ɠq,K����]&�Y	��g���������uE��
ı,O{�٤�Kı>ǽ�i7ı,O{>��n%�bX�w�^�M�3�ϓ>[����v����r��~ı,O��{Mı,K�Ͻt��bX�'��צ�q,K����M��	��T���c�mɭK%44�ƺ�6c���.�qXk<N%��׍��D���3I�B��-T�M��	��	��ku�.	bX�'��צ�q,K����Mı,K�{�Ɠq,K����.8�h�c
TUU;��!2!}��K�p�����Q,O����n%�bX�ǻ�i7ı,Oc��4��b��g�ݫdG���ec�6�3���1,K���i7ı,O��{Mı,K����&�X�%��{u��JBd&B�o(m�:&��T�4�N%�b}�{��n%�bX�ǻ�i7ı,O�ۯM&�X�%��w�4���L��^]�<��e�S*)�*j��� �,K�?{�4��bX�'��צ�q,K����Mı,K�{�Ɠr!2!y(Q���7U*f�7*S�C�Ή�2�SB/�1`��z�
�e�u��:�W��$�B�!aGl����gɟ&|��]~�Mı,K��i7ı,O��{Mı,K��}�&�X�%��t��T��� U.��\!2!2��l�n%�bX�c��4��bX�'����7ı,O�ۯM&�|�����{�Ժ�R����2��+��!2�{�Ɠq,K����]&�X�v��>�"�
%GeEx�@CIP>D�M~�u��K�2g���p��L��]�fmK$��5e��q��I��%�b{�ﮓq,K������n%�bX��}�I��%!2ӻ�p�Bd&Bd-]͖��S��ۙnfs��&�X�%��{u��Kİ�(1�����'�,K��?~��&�X�%��g��Mı,K����ر�d-o&��N���D��s��'�]-�N��:���/m�G/70=1�R�4��bX�'���Mı,K�{�Ɠq,K����]&�X�%��{u���	��	��E��%��DҖ��u�i7ı,O��{Mı,K��}t��bX�'��צ�q,K��=�7�&Bd&B�Q���rʊt���4��bX�'����7ı,O�ۯM&�X�%��{�Ɠq,K��ݛ��!2!b��3-�T��%7��&�X�%��{u��Kı=�w��n%�bX�c��4��bX jEv�
��-��)�l@,
 7٘��7���K����CYR�SSLT���p�ı,Oc��4��bX��A�3���i>�bX�'�����Kı>�n�4��bX�'���g�9�l�΄�n��`L���A]�n�zS����ۧoi!���q�]=jg�j������oq����4��bX�'��}t��bX�'��צ��>���%�}�~Γq,JBd,�g�S$����j�jnL�bX�{=��n%�bX�w�^�Mı,K���t��bX�'����&�~R�I	���ޑO(�ESn�說w�,K��u�i7ı,K�w��n%��b&"s�~Ɠq,K������	��	����e��*��RKw�Mı,����L{���&�X�%��~��Mı,K�g��Mı,S!}��K��!2!f�w�KsN�����3�&�X�%��=�cI��%�b}���I��%�b}��zi7ı,K�w��n%�bX�|H��{ۻ���v�@Y���E:�]��B��::������� t͓Ff�	�v]���sҕ�e뛵�̈�g3�m��+��IͮԠO��]�k������Y76������[t��K���,��
��H�붶����&�>������v.�3�v��`ϭ=����=(�e:kA���	5���ڭȝ�Ό=���ۆ�8����,5����������Y1gͦf1e�y�p��I����ʓ�s���59�F�=7f�����4L�
e*"��yHL��L����n%�bX�w�^�Mı,K���t��bX�'����&�X�%���̒�RT��S�\!2!2w��n%�bX��ﳤ�Kı>ǽ�i7ı,O����7ı,Oc�CYR�SSL�*���!2!<�}�&�X�%��=�cI��%�b}���I��%�bw����n%�bX����dv�U-�),���~>L�3�ϗ����&�X�%����]&�X�%��vk�I��%�b^�Γq,K�wk=�$jV��Ւ��~>L�3����ﮓq,K��;5��Kı/y�gI��%�b}�{��n%�b]��w������z��mUF�F�M��(s��tC�=p��^�g�\�*uDZ�ٳ0�3���Kı;��zi7ı,K�w��n%�bX�c��4��bX�'��}t��bX�'�'t\x�Ƀ8͙Ę��Mı,K���t��P\�ˈ�A��F$0"Q��~
6��'�,Mc���I��%�b{����Kı;Η���	��	��E��%��Dԍ:��t��bX�'����&�X�%����]&�X�%��vk�I��%�b\�m\.�	��zގZ�L�C�g9�4��bX�'��}t��bX�'yٯM&�X�%�{��:Mı,K��ٸ\!2!2��4��P�BJ�6�7I��%�bw����n%�bX��ﳤ�Kı>ǽ�i7ı,O����7ı,Oʡ������ɜRH��skn��B�S$Kح�e�y���=m������pkh�`9�۬��^��{��%�}�~Γq,K������Kı>�{��Kı;��zi7�&|���o�'�8�l�Ie�����bX�'����&�X�%����]&�X�%��vk�I��%�b^�Γs�ϓ>L�wk7�8�
�m��%���ı,O����7ı,N�^�Mı��:�T�����;׳��Kı9�{��n%�bX�w}��]-m��VZ����3�ϓ��צ�q,KĽ�}�&�X�%��=�cI��%�b}���I��%�H[��NuIR�i�"%�E��	��
Ľ�}�&�X�%��=�cI��%�b}���I��%�bw����n%�b�СFz��-�}U3M��Zi5B�HuG��ȏ2�R�;B=v�`�I��wц�R4ꉚ�B���L��]�{�p�B�,K�g��Mı,K��צ�q,KĽ�}�&�X�%��Ok�.i���2Lg9Ɠq,K���ﮓq,K��;5��Kı/y�gI��%�b}�{��n%�bX�1��LcP�BJ���w�&Bd&B��z\.	bX�%�;��7ı,O��{Mı,K�g��Mı,K�����$�MU6*$�.L��$%$)��gI��%�bs�~Ɠq,K���ﮓq,K��G@�T`� [Z�ByDZ� !�J��W"�3���i7�&|���{ߓ��H�l�Ie�����,K�{�Ɠq,K�������bX�'yٯM&�X�%�{��:M�d&Bd/B���h&�ʦ�SȉD��j���u�8�:�;k��F�wi��W��ٻv��3H��u����w�����ow�����7ı,N�^�Mı,K���t��D�K��?~��&�X�%����3�tU1�(�����!2 �;5��Kı/��gI��%�b}�{��n%�bX�ｽ&�~�LHL����%J��R��M�&Bq,K�߿gI��%�b}�{��n%�bX�ｽ&�X�%��vk�I��%!2�Y�T�4蚑�TL�\.�	�BRB�{ޛ��!2!{}�\.��bw����n%�bX������K!2!oMn��jS�*
D�T�.��b{�����bX��5�}7�hI�?{�즠�	���A$O�((������ ����AEZ

*��PQW������

*��E�
�1 ��b(@��T*����* ���Qb(V"�?�Q �" (#��PQW������AEZ

*�����U�@�����((���AE_�

*�

*���d�Mf��.�l9f�A@��̟\��� z      m��t�  �   � � @ ��TR�(   �BB��*JDEU
�� P�H�QJR���T( *
J�(RK    h@E ��{�,��ZW�WY޷_/��h�h�����g@zs�
S=�@�� �@�s�[�4 (X ( ( (   � P    ��    uLM+�N&��4����0���R������U1Qӝ�]4 �
 "�� �(b N�Jb�LM��p bt�p �|��{�.�;�e���{^������}�yμ ��N�y�@O}�k��׶��z�����:^{��z�Zr�7�{�{ϖ�Lvz[� }�UP *� ��
=��-�y��9�^�^cNox�����k�k����y��[�� �q����{yn� ��n�{������ w��nwy�o7W��OS�כҞ��
<���Z�k�/���/^�{�m� �� ��(  ��P�=�&�����{����m�7�� z�Nw}{�y5�7{�w��w�w_j{�K�{O'�׳��x ]�ݭ��:�\ ʖn�7��s۫͞�wy�u��� ���)�|�qg//=��ܛ�x x  @    }��O>�˝�F���ٽ�������� ;<��oM{}��_w/6����Ԯ����-ɥY�� ��v�n�g���@�����Z]��嫽ܧ�x�}�� 9K'+�:��gO����ڼ S��T�%JT � O�FԤ��!����O��'�F�h�=��I�JPa2 OД�)*��db40�!&Ҕ�Q 1)�'@��?��?�?�����d%=�	��g����n�qTW���/��EQ]������AE�*�����+�����A���!'�H0ӱ$1�0�A�I�C�.C�8�朳g��?��g�sf���NM%a�XX��#Z��`�X،Jc��cm����s8�����,�퍿<5�SlK16da�����!�X#0B0�4�dP���y�8�Oߒ��[����"�o7�gf���x~�8y�`��¬�����q*"0���pI �`i�0Z��()��4��9�{ �0#&�`�\d0��y������cg�f��l3Dc`�!�Xry��:6�d0ԆK��N�d�,��f�LAYh�kc�:�&���=Ԕ�@C������8�8$�I!),��>����q�d��<��qC[K5��z˙�GS����8F6��DP����p�ћ��~t�\�$I�<z��o�����'5���5�ZVd�0
XIԹ�`CQ8i�֠�4��zl'J~aqM.�1�����/]F���`���$	�pI	&��Gk��f���=������$�H�#æ�YQ�Y�߽�s5�=�8���a�Xke9La������e3��g�L��yf~���������ͦ5>,dc,$����;H��Q��.��5DjtC��s���6[�qٯ��oѹx�.���(,����1��	��O/�a��h�'J��
d���tF���³[<��3I�|�t���g5�wN�6;�&�!S�n�z��Ω��+�,�H�g1j�޷����푽l���_�9-RRh�4>����n�F�c��F�a!��zp�F�A8�
b�!rL��I`"t��BIBb%$I��#E514d��n��8i�BAD�AT��H�5i������ke����
��<���`�B	�Iqȁ�1Ӊ�
q�#��p04�P��o͟��8�d����Y�7��EXZ�ֈC�0��"?6l7E�=(8Tlxk��~����H?����&�1��f�3N�sHF��F�䆝Ǐ��Xe�6�h�,��	&2�N�8�_~�Tr냥mP�
���AT���7{�{�����߮����n��¼߇���#�>~�^~�ן�	#0�	��m�r����X$I7k�����h�F�Af��Z�kaa�6Fe�ccX{��Y�s\�����<���³$���ER|wS�c�������s�ʔQK�J�F�ه�s[�٣Lf�0d����IkPzPY��4y�,f��a�8�h�pd8p �'Bl3Q�s	d"H#�C)�~Fkz�>G�?+K�]~_��Y�P�@H(����ف�w���u$�Ri��He�V	�#�e��݆�݆�u���a���ȍ��LƑ�R3F�=��l��5ݼ~ߚ�Xy��W����F��O�ߎ��׋�z�!��q�w�=�{����5���N~ۆ���`a�s�����i�k�7�Y��h���,ȱ�8�L9�� }�>�w�).>p��W2�>��>�C���Q���#4hsK4�i�'1ѷ�bu�^��{��Q\H�$8�RVG��f��6Ea��1�l�F�M)�A5fxzq�#��hƵ���7�'��%���'�fi�A8��h��QI��v�v�HrX�`2b��l�h�Y�4������g��#I)�h �C`�4bI,f����m9�~�$�����4�`�E��I&3�(�����Fk�~��K$a����5�獮8����k���yo�6f�~?	��?%�����F�0	ǌ��l�hbߟ��xkFs�gd�DAF�mS��%h�N�04Rf�`�����z�c� �e1g ����1I"4bI�9��pBL�#��!��JmLL�c�u"	P�H`��fl�k��Fko"���3���'E2&	%�!�(� C��������ޏњ6�h	gdΜ$��<c�F��гM��
d1�O^'�)$�aꔪ����ok���q�09V�U�U,���&N�F!��� �a���ԓ2�e�~0 ��`F.�eJ	<'�[Ca���6m# �F�VkLb���1d�Na����z}�D(d�(?Kx�i5�����ȱY����-q�c��I2L��!!)�9��_����Բy&,$�#�%��}sZ/4��#4k�5�J��Z����6��k�~����٠������X[�Z3Y�[�]C�َL� AQ �%�4��Dc������q��'1��?n#�4xzr�Ky���69�0��rp���D�ct7:��pc4n�j��2ĸs��� ���F�%��޳��B��捌8D����2�6b��6a�?{�kX@�˅2��C+�*�����q�k��h���'�$"��D�M�Ei�ٯ�oÆ7�Df�[x��[�[�%�HG��&� ���8��IFSn��`j 0��v�:6Qi�i�[l��v$$B6BhŔ�0���C�:���R�+f��k6NZǖ���!c�'ax�{����3�5��I�"d�)>������pCKHa���2"�Ĕ�����4;M�O�Ȣ;R)�M���tI��R_:⋂b8%j�D|�Z�+w"�ͽS~����_�!	a�ĒU���ɂIa�p5�"�I���,�IŐ�t�$L��KF��'^=��h+����?��2�H�-l�Q��g}9�y�����o��{s��p)�p$$$�`5D_�+:i��A��g�LN�OBՆ��1����=4k���?g���!���)���.рa<@� �0D	&)�g ����2�.���i0q'�R�ɿ�~��O�I�t'\BM ��d��~��た���z�����-l#F�p'b
��d���W�<���"I�A��L�Z9�{~�����{��g6��	�6F:0chy\ҹf�3f�LBp`�;����>(h�י�F�O0�%�-�6X�u���K���k��#�a����������88�%8�ReD5�~y�ޘ�g0B4�Z��[/��C�Y��8~�y��,��H�Kl��ѐ�BI���}�����;�l�M��4�h�,c�I�#4v�h�J,Ӱy�<��%(I &//�h��g27�/5��7���9�o�9��A��i�Ȣ$a`FF�h�������<M���BH2q$2�����"b"w&Y���_�ɹ�_ܴ�Yv!�j}�y�¤�ڿ�?(���Ml-�l��|40F��bX�����D��4 ` ��L��t���'��S�b�厨�|�^�7�32�ؚu��=�oι�Z���}c�oTFi�&�J����h�ҌX�!�`I>�����Sǘ��6�1�����FZ��̽�h,4���S�q,]M
F����oC��O;��d�4����:7�����h�ĝ:�t����hT�,@j�ÍC�S b،�'d�h��iiv�jٚ��(�e��!��QDg��f�����8G���L��7�k5��mҖ$`@������������݉�����e�0Ŋi���X/מy����4�mݎ�wF�14=3�w��`l���  : �$ [@8  It�     m� ������e��[ɺ�m�R�|%�Y:ISUU��/*���e�T���[�m���Y��k�㭠  ��R�J�]U:.�ꍖ�[[M����C!���U@��b�Pu=H0W]U ��UR�ʵY�^
�G-��]PP6X��D����wn�5dQ�ڪ�u��js�U���In.�em*��p  H(�v�kk�mF�(�R�Wj�K>�����m�{I�8����  $
�	yݙ�#VԫOٶ�h[@�D�۶6�m��vPA�V��U� �@� �Ûm�9wKn�׋n�!b� -��-�@8  *t    �$�mK*Gm��m�-� F�ڴ�� :�ВY�d�l �д݀ m��� ��m��n�Hz�R�   �  �2m�[�mZI6�ۀ�V�A�݋h 	�5l6�m�E�� �`  ۶�� �H m�������m� -�m$�mmٶ�p :6�E  ��[&�k��� n�L��n�@�t����%yԝ�#�f�2M��Y[ �[p ���m-�� l�m�!��qx�m]�  ��@�   n��u�ݹ���np�a���lH @ ;m��*��]�j��`����m�� � Z�-�m�	 o$4V $ 6ݧDY�֗�j:��t[�m,��p�HT�F򑙪�%a�-������ 4� �[���y�l�  �� p����Q������P�� QUO1Ď��t/U�V�^���j�U����p-� ۉ��6[m����O8�9$� X�����am.��oP	uȎ���b�m ky����Y^g��j^8�̪� �N��@��k�b�yd�W���.�e��*�,;�c��R�R��l ��l�ᶒ���p�a�l��F� ��I�[`�)u�6�m� ��` �>4�퍶�\m�a.�[@��l ����M��,ݪ�p  UR��J��㊅YVtUUJ��Bj��b�ܻ -����$� u�a! �m�e��jU�yU����&Z�E��-��n� �E青�ěk{6 6�m��khm����h`� l���ާ@6ٶ�  �o��  :�  [@�c��m�ǎ�q*�Q�k���%���m�Hm�������  �`���O8��l 7m����v9��5U):�OW'�»�\��\KJ�T{kj���� *�*����*�۫T)f��W��,n��gP��SdI����6ٶ uT���Q�n�UV���dS&��.�[q�� m���!�l�n��U�8)yG�̠5JK����iV��<�K<p*���kn�[/D��� �3R� e
��'���*�9�V�VӜ'RI��v� �����㖹&v�-����d 86�����6��l�j�@E�RY^�2�yn
ݪU�nݜ�K5R�,���YF�"�q�%y��ֶ�n[d8p� 䆶FH( 	ӤH5��oݹt��c\ ҩ��d����,dz�h ��Am��B� ��fV��YP� 浀 6�?B���V�K;��$�@�M�$���!m$I��Ͷ�im6�`6�m�n͚�Y� �  8.ݍ&�[��U�h�;+�z���v�e�)��l$Z{gd��ݞö֟Y,��l�|爉gn����B�j�   �>  
���&0�j��.�`�h��6*��۝�5,S  h�r��l  �m�kͶ� 8���m H    q=zIF�C�nL����0[x� 6�ZZͶ_��> m��m������$� $�[[I���� H �K)��^�m�  �k��抷Y��#m�� m����շ���[X-�i��-�@K(H � -�f�H`    6�fհ   �ޒ�X�V��ZE��� qPm� 6�  �$$�c�Am�[@�E�ږ��^��-���6ٶm��n *����m���T�|��KL��BD��m�  �`�-�m"�m�6�6�ޥ����m�    � �-�	8-��X�-��7r��� p�z.u�6�y�w&�:	<�ڪ��96���U���UU� m�:ĺ�qͻm��k�z� m�  ��t:�J�%�[RHH-�s��R\І
�j���i,��=9�y�Ek�$�8ut���6��jP-�m�    � 	t�
�BMɲ�U@T�첼�UR�.�-����M�@r@ %UNZ�I�-ڵ)�I�:˥��^��!m [G� �� 7�ŷ�h��g[�ܖ6���`ְ	M�m��[ldh�Mgb­�r#V�:lH� 
2-V�UZ���f�n�l  R�d -��  m� 8m���۫�i�ۀU*�'KP �WU��IƟT珞�� �l H�[Rh�٪M��&J�6�UUNR�6���m"C�)M�i�wg�U]gn$�� �`���lV����e������e�n�J�j�
Sk[�-��6�j.�]� ��-��I� H  �,�[m�M� ���� -�lp��Ŵp �m��imfR��f�Ҵ��m�6�"Kh ma�;j�I ��&�!BY�`Ry�<�� �'d�-U�)Z��
��i05��'iʒ�T�,B[��2����ݬ���l�ñ�g�y�ݨ�tl�9�H�彭���[�j
�WU8�Y�,�����6��~����=u� 6��	�5�2��*f8'����p;�R�ʿ����WJ��R�/-T �j���w�|��e%�y0[ J[Kĵj��X�lU*�*�@U]\��ʎ��El����9��<6�m� :��[+^��$�ՠ  ��ն�^b�m��]�
�e���$�r�)d	�t�oSm�Sl $��6�IƷ���ٶ�$ H9e�$�#m��p m��,VԧL�E4����*��U�Wt[O*��V^�r�U@��h$m�m�C �x  �۶ͫN� ]W$���j$���bVt,Sm�bۮk��mK��-���  <���	-����jP�l��ͱ  �en��Ir�צ�� :���(8�*�WEU++�Ơ��S^锖��z�]]���kAJ�tÛ�/��j�t�9���s�mI"GK(y�(����3K�vV�g6� $ �i$�{at��m���޶� ��Tb���|�\�Z��W��XR����  ��u,���	6�4���߾�&۳Y��8�lνh   �40-�����6�̒� ��lŵ,���L [u�07ԭ&�|m� v�$�h����$�7l h H6��i�t�\]6  m�  ���e�(m�` m{&�Ti�`U�\i\��n�� ��i.�ڲ�f�`U���ᦶ���ʫ+T@���6��@n2��7`�����P%��Xڗo]@�]�Xv 't��m��W]llOI�L �  �di!�K{v�����`oYZ��cm&m�m�Ammy&��m&m����   �e�-�[Cm�js�S�h�im���p�v�� ��mR�UQ�r��$�mJ�' 6۝��c�Ad H�[rD�l 
������$��[\mHMUu�]*f��V$���cm�$��G��V��j��� <-���.�[פ[[m�$	6��`�`����  m��; -��{ni�d׭H8�� ` |���6�N$!kI�m���c�ր$� ��I�mfa�lH-�ڶ  	  U�ݷW<�Fڗ��T p���I��K5Z��t۝%�C;3K�p��堮P/Sm���-�p���6:�l��[@l m� imm�r@��V�+��6)V;S
�  H[M�m:lm���o[d%�H��� 9�퇥շ2k���S\��z����!#��@���I�k�� m� tN9m� �ݒ�$p n��S��H#�����&��Y�v��ب2:Z���<��\Sv:�RYؠ��Z�'h����5Ӏ�(ͩ6�
�Uo E:A� 7�!;uJ�u�9Am�[E����˶ۓ��88	6�ɛ[D����U�����Wf����U]�heA��Lj�H�z���;;n�S}w��k{޷���EN��]�$Q�0�Ч��������b�8|(��j���H؛`Y$�:�D���U��`z�.�]�L@�����'���)#,����S����@ׂ�
⿽	P������z�3����*���S�@(`��[ډ��'C�B����T�W�©��$������F�Ӡ�{�T ��t��`�\�QaX���">�
���^���hD=z�����'�^g}��Q�
�@��^2���qҀ� �Gg�wӣ���=UB�L��\|vh���	� ��}�OS�E�h�PC�:` �	B}Q3i�4�^ �1A8 ~� �� 4	~\��+��ҪN����o�/���W��Dh�Y?�����L�C����/A���lb��1I0L�$�!�)�
`��  hWb%�(oh�*��^��
t Q�h��A�H%BRb��
)����% �
P��_�y 0B>	R���I_��U�)� Á�h����I�CΈDWX���P@: ;@�A�1CJ�x���D��� ��.�H��$^?��� ��U�G�(03�a��~]�}����������5�+ҵ�q��1��ךI!&�ډ6͠1@H8�+v GJg�ҵ�iӻ�l��&�Le�1����q lJ���+�-<��J&Ń0����WkS���mgq��pfM����L`���!*�@�޻��e�W�R*�0�]�͉%�&���s�ca�`* :ݴ�+yW���F��:�MiٷC�$<�fܷ� gJ*Z�4��)N�kl6����\�n�a��(:r+{P�egh��^vi�a��.l�����}Ϋ�f:ɰ��U� �(�[@.�wZ�UX�����$��N�p���ڇ��Ajc�cH�a���V�2��V�&V��4\,dy�yK�猣�"m��l�۝ф@CA�HO/��M"���i�=�f�3�6�:4lR�Ѯx'���Q.��� �*�nL3�H����vۂ�6��r: ^�PE�\��,�\ɮ���V��Xm��Um#R�q�V�t2I0���UA"��������h�Ҵ�Y�A�W��Ŷ�7Mmm�mUUJ��
�˔\��V��������Բn^�$�i��:��(�\>�J!胝�����.�Q��Lu�.LL�תt�q�H9��;r�[oZ�u�ti��p�XΒ't�r��q�r��ј��`g n@�ls�I��X���i8nK�H^�*��n�J���k��ĥhGb�wf�vJ9�y���R�(��k\pY��Y�P<g����C�f������L�b'� א���;!Σ��b�����9�j�	�l�Ol]����m�[B��]04��v)�`����sWR����K�'A�-)�����J�����C���K �-V�-v(8�ACk�e݀��n(�v��@5]���`_0m0*�F��津���p��)h˫��,KX�ڳ��ݹ�m����^����vK���em��9뗖�"���'@��ޭj3[ulѻva��邁iA�_�?"U�� �Oj�ࡱڪJ z� �x
E4���X6#����ۡ��k���+��D�jl���:07:`-��j�cT�%h[�cb�˅����*W���GS���"n9�1ձ��fٌ��	s�ƧK�P�n�-!�3l�k�����Fv5t�DՍ�
r�.�����1�pR���R��f[���[�]; s��&v��`J���ۣhWLi�;Mԗ����P(�pG�^X�5��ff��YY��{<�3ۗ�8v�>�'aNM��8;<�g�����c����0����uު��/O[ ����Ҕ�D�g�ҹg�j���ǚ�[���f�`nة:1NH����ؘ��`sfA��l��f&�c�N8�[���f�-�vq���S�MTc8�l�05vK`wob`uM���r^b�.�H��=mO�JnU�Nt�6�ɫu�ٱk�p���٢N���{o2�s�}Wd�v�&T�ll�0'e��1')�NH���W+���;UK��'c���Ql����fM,]�v�i��8�S�I��e�`uM���̃?|�[�[e�&R�h����	�`}�4�1wu�ǚ�=\�?o��{|��j1ʉ^Y�'��o�l��L���ِ�?e{oԨl����Rn6"Ri���]V���@�b�P�����t��d:��X{983�řy|e�&T�ll�05vG`op6Țm�pj�8�:�5�ِ`j������ݽ�v*�B�Q��>͚X�����Us�r�W*$�1!��/{�s9W����*+��=��G$�RHX����Ș��09� ���F+����˫��`wob`v^���̃Wd�m���?f?;N�]���Nd��k�#T�z',�r�9í\��qn�:��͵�aK/�l�6d�%�;��XK���Jr��T'��l��T�����sɁ�6[ ݕ�Ye�F�Q��Y�}ݫ��q��.qqq��ͫ�٥��Ր�Ȝ#L�G%J�;��0:��`sfA���T����/�}�P<P]@~ֿs\�ｯ�D�hc�U)��չ���6i`b��;�5X�/g��F�I9J���&�x�#���8�V��:8��vE�ܼnj�N!5Q����u`b�� ��{�O�B�R��>��┥/�V�ڕ$QIS���A�.��*��JR~�=�%)O��{�)JRy�{�r�r����ѶME)�)�NHR����py)J~���qJ~��?wﶼ��;�����)Iޝ��[��5������x<�����_w�qJR��~�k�JS����R����{��JS�?{�6[5�[�[�5�qJR��{ݯ%(����qJR���~��)�;�u�)JL@�!/`���=ۻ������ ��j�{g�vv��1�iA��c��.yfKn�v\��Se�H��9��Ӷ�'�9�m�m��A�f��ȕ�ۢ#��`�v2�ɚ܏*C�v��_�cD�g,6⻅sϠ+��X�j�u�z�3���&�'Vmnd�7&�|sX�mZX;��]Hc�W\&���ld�z�15JWJ�f)�\�fѼ�f���{���dG�� q����w�ςnv�q%��l�+���]����]���{X�aݘ�ҡv��-�"����oW��s��R��Ͼ���)?{������u���)<����R���2:��	�H�W� �q}��k���d����g�)?wﶼ��:�u�9A�Pr�sA�&��B�8�JR���{�R�����k�JS�{��R����{��JS�u�kF������f�Y������~�k�JS���k�R����{��JS���s�R��w����7�oYkf��[^JR����\R����{�JR���{�R�����k�JS��}�њ���F���K��+�2�/fzu��"@-�-l�;ZMqrQե6a�[hd�7S�O�������s�`�R����┥'����/%)Os�}�)JR}����n��l��[�췭��R����������G� Ъ}��5)I�{���)�w��R���������i��J%9N	�(�W�Ps���vs�)J~�{�qJR��s���R����r����֛Q�Q������_�$'u�����)I��~��)��w��)JO;��y)J~�]��5�3{�[7����qJR��s���R��'��ﳊR�����%)O��{�)o{�������ICg���W�J�����|�H���zul�{v��33۔�m�B9�Y�۷���y)J~�]�qJR����^JR����\R������<��=�惦��(���W�Ps�ϷvW.>$2S���k�R���w�JR�~�}��)K�,;��oZ޲����c�JS���u�)JO}�{��W�"2$��M ��J�Q�Jg��n)JP�����R���K��v���Z���f���R�����������n)JP���c�JS���u�)�,ņJ!R��2��%F�g8��^~�}��)C�{ݏ%)O3����)=�=�%)N��3]�l�u�t�+��)s֫t��V�|hѹ�;[N��Ɯv��R��S�q��(9�
�ۻ+�s�)�~��┥'����)��wۜ�9A\��kM�ӔD�?6��s㜢S�{ߵ�?�rR������JS�����(|�{��)�k��f����ճ{��[��)=�=�%)O?{��R����ǒ������R�����c�ԃ"�*��9_w'n)JRy��k�JS���u�(LUX�Uҁ�Q7�'���Y�Ps���A�T�Uě���I�{ݯ%(�g����┥'{��������n)JR{ﺵf�a���B����-,��F��gr�s��q���;vz*��n�^�t�:�ʙ�3��{�"�g�{�)JR{�{�JR�~�}��)I�{ݯ%)O}��ȷkz޳5����o{��)=�=�%)O?{��R����ג������R���۱�q�dC��*��9_w&��P)I�{ݯ%)O3����)=�=�%)OL��l�f�f�f����n┥'��v���<���\R������<��|���qJR��zwY�fl��y�����8�JR�����)JQ�3��~��R���w��)JO;��y)Ji
�w�s���߀\aQ�I��
@�ۖ���#�� =��حǉiSF��ӎuI��3�^#Zu۴��W���Z93ZV�r�|e8А'F2�܂�3�km�:�a9��%@+�u�hWŜe�e�*q�b�s�zzD:��v��佛�F$�kK����v��l	�yv��ݤ���y���g�#AO;�ĺ�3�5�i�۲��a^�xC.�v/'�������{��w������G6�nG��}?�l�q�1E;�8�F�
�����m��3=��=p������[�T�)?���`�R������)JO;��y)Jy��)I�}�9m��R�8��s��}ܚ_9@�'��v���<���\R������<��=�}�a�5��y��Z�kw�)<�{��)�~��┥'����)��wۊR��{�ûٕ�o7kf��[^JR�g�{�)JR{�{�JR�~�}��)I�{ݯ%)O}���"q�' �$w�Ps��Ś��s�Jy���┥'��v���<���\T�/��X���"�7�����+K�=�U�ƮVѻs��g��݈N��B6p��g��yk{ݖ��JR�~�}��)I�{ݯ%)O3����D�%);���<��:g��͖l�kvkyk[��)JRy��kȁ: By�Ĩ� |������qJR������R����/�A� ���YSqTDu!����R�����qJR��s���R������)JO;��y)Jxt����Vo{7f��oz޸�)I��py)Jy���┥'��v���<���\R����"M��9
P�*��9_w&��)I�{ݯ%)O3����)=����qy/�.�UQ)�Q�#�U��,�	V����[.�d��0o=S֣��ma�����e�V�Z�┥'��k�JS���u�)JO}�{��JS����)|���w�+z�n�͛޶���<���\�rR������JS�����)<�{��
Jw�/�V�J�:��ERJ�q8��1��9�O?{��R��{P�G�Ŏg9�k�	��Î�M���A�'���i3��i؆�í�A"�,đZ�`�$�����)�D"HH�J� �H`���~��}S|�j��ާ�Nu�����[����.����
@4�6ɠ��1!#�*~3�O`��@�c�;���C5��� iM�g?�z��&����O� uE:"���x$�����.HC�?'G��l�(����ĀЮ/�+�{Ͼ��R�ǻ�|�q�XRt�R�F��#%LJW�	����R��}��JR�g�{�)B�f������JR����J�GQ��B���,�ȹb����{ߵ�)O3�(J���}���(J��(J��"��(J3�(J��J��(O���^x%	BP�$BP�%	Bf`�%	BP�	BP�%M���. \[��J��TnNNF�X�t=&*���sHN-plwPZ6Aˤ���Z\�q]7DGR
J��. ��<���(J!(J��30J��(H��(J���{���J��(H��(J���(J��"��(J3�(J���}���(J��(J��"��(J3�(J��J��(O���^x%	BQ�H�	�%	BP����(J!(J��30J��(O������(J��(J��"��(J3�(J��J. \Y��ߣtQ*H8�rT�ߗ
��(H��(J���(J��"��(J3�(J���}���(J��)hJ��J��(L���(J!(J��?{�}y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	��}ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�^��y��%	BP�	BP�%�.��P�%	BD%	BP�&f
��..懮7UT6��Q+xpJ��(O3�(J��J��(L���(J!(J��=�����J��(H��(J���(J��"��(J3�hJ�����(J��<���(J!(J��30J��(H��(J���{���J��(H��(J���(J��"��(J3�(J���}���(J��(J��"��(J3�(J��@\@��q����j��7"��T��J��(H��(J���(J��"��(J3�(J�����(J��<���(J!(J��30J��(H��(J���{���J��(H��(J���(J��"��(J3�(J���}���(J��(J��"��(J3�(JU㲜a0�W��mW��%	BP�%	��y�y��%	BP�%	BP�&f	BP�%	BP�%	Bf`���q��/��5�@ITRJ��(J��<���(J��(J���(J��(J��(O���k��(J��(J��30J��(J��(J3�%P�O���>@�@����뀃@�B{��A�4=����kz֝˲%r쓀dg��F�����`̽s�ķm��Zw���7ݯ����nk����P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B}���8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	������(J��(J��30J��(J��(J3�(J�����(J(O3�(J��(J��30J��(J��(J����y��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BB��V���R��7RFJ��. \T%	�`�%	BP�%	BP�&f	BP�%	BP�%	B{�y��P�%	BP�
P�%	��P�%	BP�%	BP��%	BP�'�}�8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	�^����J��(J��(J3�(J��(J��30J��(O���g�(J��0J��(?�\��(J��`�%	BP�%	BP�'�n�q"*Q�d�P��q�����(J��30J��(J��(J3�(J�������(J��0J��(J��(J3�(J��(J��?k߾מ	BP�%	BP�%	Bf`�%�%	BP�%	Bf`�%	BP�}���	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	B{�y��P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B}�|}���[-淸���	BP�%	�`�%	BP�%	BP�&f
#BP�%	BP�%	B~׿}�<��(J��(J���(J��(J��(L���(J����(J��<���(J��(J���(J��(J��(O}�>��J��(J��(J3�(J��(J�hL���(J�����(J��(J��(J��(L���(J��(J�����7��Vo{ݚݖ�����(J��(J��30J��(J��(J3�(J���}�pJ��(O3�(J��(J��30J��(J���Ur��=��^x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'����8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	�^��y��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP�?�
���{���a�	��e�tx$��-���8+�`-i�k�9���ڒ�nx�b�9G����q�}�w���P<�5n���lc�j�lu����.ewku�c���H��&�c���a��<qڛ$$���`��6���������fUAJև�w"^MӒgj�!<��e[8t�-��YY�ˮ�9'-�[��;B�!t5�1-=S<-"]]\Y������ww�{�{���k$Ve��]МŮ�5�S��c,c�DD�;�k�mGc��;�����*��[�kV��8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP������P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'�}�	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'�{ߵ�P�%*�	�%	BP��%	BP�$BP�%	Bf`�%	BP�}��ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�w�V����[5k5��x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B}��p��%	BP�f	H%	BD%	BP�&f	BP�%	�%	HR���~מ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP�}��ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	������(J��J��)���(J!(J��30J��(H�ߋ�����ٽ�Z��(J��<���(J!(J��30J��(H��(J���{���J��(a�JO�Ͼ���~5)�~���)JO����%)O}����J�:��ERJ�q9�I�[�u�%)O��\R���{ݏ%)O3��_8��A��̎5!n���y)Jy���┥ʿ��lJR���k�R���w�<��?~��ѭ�N��z\1-�/2]��瑕J	�78*͇8t���=�����b�s�ƙ��R��}��JR�g�{�)JRw���"?�~��=�����)I����"��u(RT\��A�/Ͻʴ�K�������:���yϰy)J~�w��)JN����O�G�J���7Tԩ �$����/y��<��<���)����c�@�+q���+��l�6�6�eGo[��| $'�Ϯ)JR}��ly)J{�^�8�	� �}�}�q8��4�#M�)�)�B���$�{ݏ%(�{���qJR���y)Jy�wۊR�������}�l3��i2����fݥ���ΑTgj�v6{Qq�'rs�w^O�w{�s���{���]��JS����┥'{��%)O;��p>A%�JO���%)N�����2��L��9�]ǘ�,_ �)����R����<��]����ż\��q}�JOeF�#M���޷��JS�����)=�{�䇂�����h�%@��8t��}�S���jS�u��┥'�Ͼ��)����-�6kvkyk[��)K�'~��%)N����R�������R��R_�w�\R9�Y�V�q�TQ��)*.Y� �k���(�{�}����﻿�)JR{��c�JS�����hۘ:�L�����˩9kY��=�K��z��v���z������y)?���������}��)I���O�/%)N����R����k��3Z֭a��սo�����}���R�����c�JS����┥'{��.YżIp\g8���
���t�(��R������R���w��)� 2O�Ͼ��)�u߳�R����ڬ����IU,�j\\ջ��)JO�Ͼ��)���z��|HT���T@�G�=�PsRs��ly)J}߫�U����Y�٭�ַ�qJR���{��J��{Ϯ)JRw���R��;��R����>�d�z����5*���fDi�: ���v�Zz�ѻ[�M��p�.xD?��w�}���Q��6:����8��[�<_8��T�����R��;���.JRw���JR���~�e�F�n�o,����R������?�_�ԧ�����)JR}����<��=�^�8��b���|}�޳6kf�5�F���%)O���k�R���;�H����}��R��������qw�՗�p�(r�J�qR��d�}�}��JS��~�)JRw��ǒ���������qJx�����#uUE4���F�g8��]�^�8�)G��c������)J{����┥'{��%)L�ӹ�kE���)(��(��˷Z,S�j�f�S�v�PW��'ۂ�B4�/"k�Lk=�N�+g�����"�șet���;9GF���Y�m�r����Z7i��c�9��K�m�ax!]�6�e9,�œ�u��t��yVڶs�-ev��Z:��]*�
Mh�M�]�-�v�>�Ӗd83�(�c�2�딺{�3l�gi��z�hѴ�� L6�g��3R@Lc6�Vo4Eq��tt�/Y{	/I5�y#�]�dY������ݾ�}�ˇ[	����)JO��ly)Jy��u�)JN�;�O�/%)N�]�8�)K��lCnB��U,�s���ʴ��=��R���?��y)J}����)JRw�ȹg�.3�[�`R*dR�e95�)JO�Ͼ��)����)�$����R���}���)I�m��j��7RD�F�g8��k�v����JO����%)O3�)I�s����A�/���8R�A�c�G|�qR{��c�JS��{�)JR{��py)J{��qJR����2����VoS��S��zSjg<����u�D��ѻ[9ź��]��F�JS�q��W,�(9��n�r�JO{��%)O}�}�K����v.Y� �ubۍ�5*H9G%_8�JO{��#C�K �p�qS�8+E��	i�m�W����o��)<����R��;��}��'�O����kZ��ktoV��JR��w��)JN����C�����w�qJR���y)J�v�p*��1�d�uP�q9�&qn��ǒ�����k�R���w�<����va|�q9߱6�"m9H��Py)Jy���┥���}����}����)I���JR���y�5��:���qX$�YnlGi��+�\[Q!�:b�B�RՕ6��ͷ�m��&�ɑ��)>�>�������n)JRw����/%)O��~��)?}���TMT�h�Q��\��A�.�م���?�WJRly)J{��k�R���w�<��Aa�O�{߬�lѳ[�[�7�n┥'�}�ǒ����{�)Nޜ�6;DGl���jM}�}��JS��\R���Ք�dUn�
J��s�7��p\_V��R���>�������n)B|���݋�s�9ŝX��t*�*A����)JN�;�JP=���┥'�}�ǒ����{�)JP�w���J<U�z�+֦�m�tv����7���p��۷n�3=�L��E���Ls�JS����);��c�JS����);��py)Jy�{ZՆ��k2ޫ5��R���{ݏ#���O��~��)>�>�����}�n)J����CY"r�I*���q~}��R���;�H|�������� ��݋�s�9���b�2Jr��kz┿�A�w���JR����┥'��v<���z#���C�>*�}𸪏����|�\R���tt�G)S����!���s��w2i|JR��������c�R��>����);��py)Jw���f�ѷQ��o��r�k��5�i�\�Ӻ�Z7)gn�J��$�\������"�A�eT�~�s�8�w`�R��=�u�)JN�;�O��R���ɥ�9�[�V�q�TQ��)+c�JS���� �I�JN��}��JS��\R�����ǒ|�䧾���tQ*H9GR��A� ��{�r�)O����R������ǒ����r����eek�&�ӌ�QH��	��'~���R�����c�JS�����?�O��I����%A�.�-�R��&�2QN�� �q~�{���������\R������C�JS����)$:h5ւ�ǁ��gi?n�	��8l 0�:q��K���Ǟ A�i�p"YK�����:,��[<6���`stz��Nk=��n�&����W8Vy��gB���6'� s�I��w��#����RUeb�O|���v̄2���!�4�loP��
��L���h7f�q43���� ����F�Ӱ���h)%����1�+
��q$�瞆�@&�P�p� (�_��ٽټ���a 29ͥIu������Ce 
2;8����x�<];�zSv`-���'
��{Pl��aW�U��;c[#���[�Z*�� ����s���{#�UUR��f{P�Pq�;F��-�۱�Sat�r�8�r�.�Y٭ W����`���@�㭹�
햮�^�u\V���FQ�xߗ���N�ͦ�2���vU����M���V�^�g\�X2�BUBUfӢRZ�7���_�@�&̻GRl2�v�i�bQ����URJ�,�J��lj�LI�fT
�ƚ�n��{(NWn�����D�:�9:�iŵ�q�I��lB��q�n��6gN5uFZ��6zm����ܙ��4ۛ�L�Z<qt��*b�n�WiL��Q�/�ɞF�&�y�@��pMUT<�Ob��*�ʦJ�6	Z���j�+R<N��U�3�\�;STݪC��@v�D�z]�l�v��R�0}�����#����^[F�@�i3�L�
[{7m�v	ٽU�I�u�Y�	֞��,�  ��S�we�1�f�q� ��ܬ�`9����Jγ�aX��0u��S�6�Wl���o��m�Y�02��q�{0v^DV�v���5�C��>~���{v\<ݍ&^l\�k�9]�'�7a��K�vie��z���n@��E0�z��kP��)ew%�c8p���m ۖ9i'm��4:�������z&6�A8=r�8�ɑ��C�ӳl�9���t9{yֱ붱��ֺ{l�k�lq����kr��ghՉњ�k$�h5�Ƕ�����l8nVsа*�U+��=S�q��p�v����ӫCn��̼:v���S4�֫d�M���nƧk�Yaͪʼ���1@mƀ�����T�Q��:��>Z���sgM�����t��lZYl�N����ÝzY�6q5�N��CPmV.�shU�g���ΓG8ӆn:T�v�F7a�\센��{mF�[-��G𦟏�U�����������|�(^�g|��/A(�#��b��~7��q[ �6�cJ9��wd�hwf����U��'Yؘ��!���v�=]�{Z�����V�2���sX�q�n��f�����HQ��k@q�[p=$�(x��]�\�l79���zb�{P��5싳O�mѭ��5
9���\Z�k>ic����.���=Y�d�,'kaE�8��sP��g#�i):�Rf��0�4���ͳ[ݭj�Y��*���?�My��8~��s k��$��ka�)k3�2=v�Z�3��{����﫱�cof��kk�)������)=��t<��?{�xp>AIrR��w�%+�Y���	Ԋ���TS�W� �qt���?�@�CR����R������%)O3��\S��R���Zʉ����J��J\��A�.�m��)I���k��R2S�w��)J�鹴�g8��_���8��EPuU$8�/�I�~�k�JS�}��┥'��C�J�%�{���#��VS�E�G�w/��s�9����qJR��F{}ߴ>JR��~��)JO{�v���.��c5wVoY�f�7#�j^�;�sN�G$.��a�x���n^����{��wsw�}
��,������ݾ��JR���xqJR���ݏ��	����)Os���\R�������Y�V��ޣf���y)J{���#�S	K`B��P-�� K��e��#�И�9)I��}��)����)JOn��/s��8�(�r�יj�r�(�R+R������%)O3�?�d����JR��~��)J^��0�i�2E$����I!q}Y�W�"R����C�JS�����>�Vnl�,�s�3�!:�Rr9UCu+�R���=�%(�g���)JRw����)�{��R�����x��u��Kl�eWQ,�<�j��7U.���]������������:�����aj�[�������8�)I�}�ג����{������JO����JS���|8��EPuU$W� �qw;�^G�!������);�w�JR���xqO��]iJOo��g���ke����9�/���s��?�qJR����䄇��x��16#���Js����)>��my)J~�t�7�֭�[�f�e���J_��R}��`�R��￸qJR���ݯ%($>�s���9\����M�i�T�$U\�{��P}���)J~���)JOuf���9[�A�t89M�"q�S�`��X ��w6����ф��7�Q�c����{��G��R�m�d��H�s�9�Y���%)O;��R���=�'���JR��~��)J_~���{,3[2���z�ג����y�>rR��g~��)���R�����k�>rS��}Ȍ�����7�Y��JR��g~��)��{ÊS��w����)��}�)JRy���]͚7�xf����ox<������~8�)I����^JR�w���?"��!
<��R�H����π��̓[����R���~���٣f�f�����┥'���^JPO�}��┥'~����JS�}�)���{����K20W��H�t=&*Ѣp�uhA��c���]$/&�_�����>q���y�޿�9��JR�������)I�s���R���{Á���)I߻���r�����z�m���Dn;�(9�$���py���.!�O�����)>���k�JS��{�)��Rzt��:uAETb���r�q8�3m_8��A��Ef�s�$��wj�ͬ�`~��p)II�JNP�H�5.qs����V�wj��Wq�j�8������wul���*$RJ���3*��^���9���>w}j��w-X��_9�?�w *�73aV�ٞ3Yh�x��n�l��b���]�v�+��@9����J��b��t�'	ɹ�mѶcJ0:l1=����Y\F���F�5K��Nҽf��{(�<6C��Knm�5�i9]c�vo�q�[��7.��7	���6���K��M��@���sg�Ҕ�O'��f�f�s�Z(Pmhm�b"n�M�y��j��	U=E�'��sn�[ֵ�֫X��%�a`����Q�B�f�/\�Ic�����6w�ĒU-�'Q�ܕ*�uR���ၻ��f�^��������;���ʺ��fR������f�L)#�3ri~�$v��h�%:��G$�zy��Il�%=3�I�L)[O(dUn�y��k�y���U���K��Z���s+�Z��JT�r�yl��`UI=���ΘRK`~����Z͚ĳ���t'1k��P�yy�s�}9�fw��Tڎ�g{s��E�����8�Θ6:`qI/�A=3���|�h�(Ĝ�`f��]�w�!�/^i�(8W����U���*���W丒M�����QQ"�UE`u{޶��3�RO:`OO:`n��'Q�ܕ*�uR�<�������͵`w;��7�/Wg��;��z*R�T��2�fݎ�6:`qI-���K�4�L��"r�u�P���$V�rl���:8�6��B�l��P�8���x��̦͎�RK`l܃wc���,FU�bW����u�:���\��?�To�x�7w֬�r��l�W��N��
A����fmՖ��%w��'���_s�p�_g�|��l�&����*Tr���}Vnm���ʰ�9�*�o�r��)FIJ8�D��X��yŵ���ܞ,�۫�*��~ֽ�SMn06.kٷXx�]\�@u6Wk��a5]���pζ�IIT���)�T�H����3ri`w�{�/�1�mX��!:��*J�:�Vs��q$ٝ٥��sj���r���I{�\�;��z*N(Ӫ�'$,�O^w*��Iq7׹�`f�����{��DT���*�a�I$���ڰ:�6��f99Ӝ_$������Ny��}r��O��j�f�X���*���K�L��`Ñ_ٕ`.s����:Q:mP��J��А��27�壪���8==X:�-j-������{���pr1H$���o�OŁ�٥�����q$��0ܬ�`}�6�:�P₊T���d��qq$�1�v���v�م�s��9Tw){�J2�)Q�R�`k�z��w�����������وk$Ct�R��J��.q�L���L������l�&R���INJM�G`}��XĖ�oO�c��W}׽�U��!lHU�G���~v߯~����@��5ʐ<�MeW[dK��
З<MR]�ӎ2�nq��d�.#���k�{���ݷi׬]T��{q�1Mpg��1�l��5�������iy�TFA�/.����s���� ��<���3Yu4ʛZ9lf�dgj���S��3L�N��syRvi��ݎ�v�L	�[aZT�p[3h���ʍ�r��L��*�4?�Js:�<Y�lC����4�\��Dq�筺�jlX�T�:o�Jݖ�.*R�Ӫ�'$?������l	��{� �L���/ObhR��'#p�3�4�s�ďk�+��K>Ʌ�.%ě>z����*(�J�j]��mo���vag�8��f�wf�z�e�UA�C�mʎ�R�}ܽ,��,�����.*�����^��N��PQUHX�L,�Yݽ?�Y���;0�=�'���rUIN;D�䒻�\��K^pN��qv��nϷ;=�C�,�墜�"R�q���������`nWq�gf���ݚX�����R�%)%HX��;��j]J.$ĒGY�p�@�� 4H�����9��!�?O�饁�]�^�l�F�	ָ�T�JM�G`f���ϲag�8��9U�[<X��;�aFD�S�$䔜���٥��Y4�7k��.'�����{�1�JD*2J�06V�����2yp	�� �3���V�qU1G)@� ������n�y��%���r[�dB�����z~��~�k���W�ի�:������va`g�0�9���Ĺľ��-�,��댩�� ۗ���r	ِ`l��0&���U��q���یt�6ET���٥��Owۖ�E���t.ض��G�)�'{��4���/� 8��?3F�6�Ɛ�Ȍ�mSI��	��@'� �@�S�����CO��4��3c�?��BГ�<��a��G�S�ʡ�F`�^���N�W4R�X����=�i $1G�T��CI����#���Q�m�z�	���D�E��Ϣ�z ����m@4 qzH��O���z��ͪ�^�9U\z��36x�>�ؔ��L��C�P�Թ��<�/Kr�]��va`g�0��b��ET�)"�m�LUW�W�����g��܃6���?w���:a��qX$�z�<�غ�>B���R�l�)�D�RՕ6��ww��n�\q:��)7U�o�x�3�X�ه����\����;��G��(�:�̥��vd+r	��06nB����l�=͎��%"%T,ՓK;]�g��s�����l�`{=<X�.��E�_�Z���y%���`f���ϲaa�qp\HI�م�ެYq�MG$Q�Tvs�y�s{���3VM,�w����pzJr:�����*���m�$vz���&�s=�p��nۇt��
��K�!�WQ��U6ET��{=<X�م������s��ܚXv���R(F��ㅁ�Y4�7j�;��X�L/y�ē`���͑�UNR�N�`nVk�;��Y�I.&��4�7ճŁ�
)�R�q:I��<�������`{=<X�م����>�"��iGI9%'!`ovi`{�#ߎ��ʾ��r�{��r��M�1�T�!Hq@��0�,��Fg6�:+��5�۞���g���Yc�I�Vk�f8�i�f�rM�7���c&���:�i��څ�^�Ō����1�+z��7i�6IOhX�V��	-�٪yzf)����n�FQ�i�m�͉V9hÍͭ1Y{���0��0h��B�m�ۧiͣf�1�i7!�#*��Ζ��]���H�f��s�.�h9z�k85�Ĺ���r�9>��_S���9NQP.Z�ͨ��NWN�>6�ӆ-�،�Y'��������B�GQS���|r���`n<�`l܃vdR�ԱW��^_�N�����w�s�I�7&��f�qvaz�\l�Z��n������ܚX�L,��9�qs�[�Ł��>��V���m"B�7!`ovi`f�M,ǚ�=U�[�q׽����b��+r}��O.=3�vM,�A���:q�@ډ�NSB�<�Ud�gvv\�uku������l�E��<�vǪ�Sj:m��Vw&���W9�i-����KXzS~R�q:I��s33?w�v���0�_�T}Dy�5�>��%�y�4�^��I)w����T���qМ>�$��ZI,�9����w=v�Io���$�iH�Z"R�Td����7?iv�{U�Um������ɉZI/���"S�q�*ll�RK�s�m$�f�s�%72$�If�z}�IW9�R���>iF�)A�F�R��N����g\CyC����m�=��Jr$��� �B�7Ԓ[�����ܙi$�h��$���v�Ioql�)Z��$*Sr|�[�jV�K7��K[�n�Iwr����:ۉFGF���ZI,�/O�I-o5�Js��ժ�Uq�����.
��_��w�^y��}'���J��B��BNSj:m|�R�e�I%7\9Ē��i$��ÜI,tl(��JI���M��$��^�|�^�F��I{�~9Ē�{.�I-��߆+�[�-�;*�i�y�Us��Y�����8�cq�OQJ�d��76H0����$��ȓI%&��I%6fW.�[�z~��}Ov�8�J5Q�UF�ܚ8s���%��ƒK�?�Ir�I|�b%9Q'���RI/o���]���/�]ߥ��IOA��Kn�GMTD�N%�ZKܮ7�߼}�I{^������}���33�=M�� �UG�rZI-ȶ��&�i)��I)��M$�����s�z�Iz{1�����������s�WHcE/j�a�u��+��>���urnX�Y��';���	�hF��Ԃ�$��K���$���i$���?��Sor���m���>l��!)�RJ"�����䗼�����rH�w������������?/߼��\\RG��A	לT�����[m��_�ߛo;R	����s�$�٘Ē쐾Y��\	�@uߛz��.V�޷m�������m�;�,=��%����,��:c�ˬUx��x0;$0͘��̃���nU�(z��V du�*$>+�#^��Vj�z�f��آ�]�6�-�s��K$Rz��+͹�XKÛP�]w��c��+�y��0s�OU����76�R����P�{k�6H�zP�6vi8�,�5�6"p  �x�hy}.2�ڽb&829t���>����u��K�a���&��x�{&��)We��Doe"c]Nݖ���ܒ��<����i�vy����vRb^���3ㇰ	.s8�Ē�,�TӸJ�"n�:�)a�u�)�Il��Zv���@�a.��g�����H��МU'͗e� ��`w�07� ��t��R�bJ�b30W�ʩ,���K��I*�s�Ł���V�͗�r��#<�לBi��!Q�B������t�;6c{2vTq)N827I�W9�Y�x��=�,��qqs˜�n{�� [�M�SQ�����`��`gvi`gvi`wwK�Wq�[�6S`�R7MT)6Hk��f��	�5��sV�l�X��';+���������QI�`�Dn�ܟ���������3^���{},��U�
��Uu7Y�ܫ���npP0!R%V@i�M���s-ｸr�����Vwf�k����TT�$Nwk]0	�1��)=��<0;�ڻR�EEE?�-]���߳ޖf�,�f�q>���kVlm�Q�A�m+�`ñn����;&0?��?,GEs%��K���3�\hN�vS����u�t�L۝�mGc�?�q|}�1�e[,�ÀzL���0	�1��2�V�JS����jB���W�H7���������az�`�57͑9U*S���E`��`w�YI}�s��!�shLp�6	� �"[���ʼ�����.�#5�@�nU!�%��$�w߼Xݞ,�kn�{�,�tvʎR���	��7rW��W�\ ����ݙ3�<��U�V'��l�mP�Y�kb��v� ۈm�5�Iɓ;�ﯾ���]Q�:��;��Հgْ��ra�s�K�̚X�b�{C�����͖�����$�ff�,̚Xf,�z���kVlm�Q�A�m����٥������?���yzՀ{=�`~x��FJ�*�$%!a��Os/K��Z��2X`k���r�:"�"+�{�v�^�V\n���5*�9;�Z�<��Kˋ�W�ޟ���`g{0�1�J�P��Ai�ظ�f�a65:�\B5 �������Jrs�{u�.k��q,�<Ӯ�`��� ���}_W�A���#tBu���*�ܒ���0�s��K�����`n�ū ϳ%��qq&����r�
p�'۳Ł�����8�����>ݚX/�.:NPH�U#�Xy����7�������=�q�v�X����#�9S�U�W_ {=�`rL�n�$N���U_|�ypx~Dp�j�C[��: � ���X%a��Rp304-	5$�y���Ҙ�C�B��U2���$8I`�1��9���d�� �#^ĐH03' ������O$�\�o�$	d%�֬M��ٰ�� ! �gj��.��2&���A:��q���
P�J*j�����X���4�"`p� [��$`��f$L�L�KA0S��x���K�,��0@���n��z����oZ5�3u��l	�kJĊ��%�e����MF;;'K��ɮ�g%��%j�6��tʵРڳ+�5u�O�V;!v�͢ثӴ�2r��f@�AK`�F4m' M�ѻ55��N\+�9��ֆf��mFۀ/Ke�k{f�%m�	u-T��%�m�`� �V�HA��K�sHN�Y��ݢ������j^��0��aӴOW*GeJZ�O\�/`:�v5L��W0�3�@ER�T�zSMm��W���ó>+�52ctG8m���!+ �IeZU��[*sS�K�L�u�L5tdF��+;۱�\Km�k�Z��Ķ�L���6�-���N�Ҵ��2�!�q�ز�uۦtF�lGK��zʞ�$������KQ4� ٫���U)um��P.ܼ����Nk��϶5UU<l�Ñ�m�WejvV�
���	���*���l�F���1]2;���V�nij�	���u%d34��m�9
� ,[@ġ5��H��'N�2Ŗ�.�kW@��+�Xv#s���U�m$�ig^ͰD���b�v^Z�Z
�N�W�l��F�ۓvv,S$ꗕ����;fʓ�U��fv�l�coG4���,J�guvPٝ����6R��2��+;wa;eʽ�*�O�et���f��*jq[d��#�G�m1]5g;I����hKI�X1lhj�W�E-TZ[�r����;����*��9�%Ð`9d�vR3��r�;k'Ij̸ɑ����K葫��Rv�w`k�;q��x��,\HoiƜ�23�:�[et��M{���#=��2� *U8�[�Vd�^�:����M�'�zܞK��
��`��(m���l�ۜu�CWc3Glt�wnr�ؠؚ�nnql��l��P�t"t�v�:A� �Ca��5��B� ջu�v���t�pd&�U'x���q�
����(q�\F��n6�[H�;<cV��s�Rk���v��"�ٚ�fo�pt�E�&�1tQqqEeS�T�����p?>�/�UN�&�@�J~:q�zOw���w�׷��H�e­�9�N<8z�ɍA�Q�C��n�-+]���d�8{uӻ �8�ώw<�&{*Y�Dnn�l�Q����K㧱v�8�R����<�Y2�ηy����d ��r����ɇ�e�UGS��!��hY��qgB^��M,]F:��و�v��6zCm��wm¹�p�b.#LL�#W*ݶ5���&O�{���;���{����������Ύw3<��e��ZD�F�\��q�綱����������q*H'I���O�M,��u�Iys���K�^���J����w ��"t�'d���?�U~��J�����R�U)J��r��;V;&09&A�7r��K�K.�%�T���.7�ݖ۳K;م��7u�V4n�N��B�R�09&A�������#��'���NɌ�H�h���H(�B�plq�c%�n'T�I%��GI��8p�.xG�wo�����*�R�~s&�fc�`�d�8���{�K�������5QH�,����
z
�W����7����7�;�<X�4�;ה��F9Lr��v� owe��d��&�2i`n�VZ�܍�h�H:��RX%�q�v��72i`ff;VM�we��kl��m"BSr�M,o���|�����٥�������JQ$R�;Q�b<�X
['U��{v�l����g�)���n�%(�S��33� ϳ%��d����ݞ,n�6�H�UI(���8�vL�������3�d������q��R�Xn�,�f.�䁂"�7���Õ_�w����� �8�Ԕ7R����7w]� ϳ%���q��zX]ݵ'($Q��G!`w3��{����f��M,;���lGSjJP6�,9�����k���%�q�U3n�����>��O�F**)�5un���zX�&w��~a���X֬�ۦ�����rK�d��ĒKܪ=�<X�yڰ��/͝ǩ�DGm"BSr�g�7uZ�RK�G�},��Ł��Yq���H�#�NB��$�w_�`��`~̘]y�������fd�Tv���0P�tɊA���_���~,���\{(��%7�`ܘ����$N���]]ܬub��gqX,�m��W�:9�	]���y��x�v��%�+ø�wnX�M�{_m�_� ��܃d�� ���va�R�D䅁��������Հowe��2a`gWr�8���F�)���D�NɌI�`M܃��WO*:u�j�_���9ē~�zXݚX��,?���+՛t��un��>̘X\�����m� ϳ%�i&���ώ�C
����JK��u��Ƴ6	�p���L�L�k��x��P����Չ�t�U��ܝR7b�SV�qqr�Y�����������ghsp���KV�g`����Ų���ز��w<(��q�gH�X�|ǡ�ȇ���&ܘK�����N��#�g��s����1�ݐ9�sWD[�dˋ��{Sb)ˢ�[s�����8�yq�J���8F�UTDm�!��;^�x:ƺ4�nѰ��m�n^����jr�Dq��$%7!�nl�`f ���W�;�On�~M�t�d"�����_���>ݚX��/W��P/o�|�U)�T��{7���J�K�p�6H�05����bJ�]�z��Rf�������"t�7����n��RP¤�)V�$��Oyr�����0���lm���Kl��4�z��#�E�q��N�{[t�	C"���"�9A"�TR9;��X}ܖew�����l�`nV�?*r����?���k�ۛ,��?'�-q'�}�%�&7r	�'O��������:h�H9�RX�o����a`gsՀ}������q���qX{�6?Oy:`�cKؘݩq&�:N2Fԅ�����/g�>�{�`nd����6�O��ӎ:�zrI��b�{5�(U#[ήg;����`��ўNt��4܃*'�~ ����Wq���=��;��Ձ�׭
�e�9T����s�l�ɥ��3mX}�/R\�*�����:!NTrTvW��o��_��;×�?�
��&(⒀H?�@�G��Rd@�6 y��������U��{�r��}��qR�F�)���s�V�ݖ���Os/K<zʒ�QQR7m[� {}�`}�d���<0;����F�CVҍ�R��N�7Q�U9��b�Bnqbڰ��x�6���R�g�)���N�U��	^_ �y0&�A���0"���=OdDq��$#q�`nd���ꎘvK`r^��RF�^x��U��Z��]����/:`�c��&�f���+"r7Q8܊�W9������k5���,)w��Ë��q%��U����`j:�QM�`��	I,�]�`.q.s��8�����f��� ����Z� NF(�(r�6ڋ��]�K��l웭��g���N5��g%k�n�R8�̚X�[u`j���9\_�}����͵N*R(�E#��;���]����0&�A����g����ԈNT�I�nԺ�����`}�5X�4�;�����[�MQ*H)��,?�K�qqW}{�`{vx�>�^Z��K�=��Ձ�v����GL$%T���f���������zX�����b���?���r��:9��f��l�8V�ٶ]�X4k����q�t
�Z��cb�AD�u�כ���1�s�K��z����tm��f\�<)mŁ��[%�p�#�/3S�Dj�����8v��ݍL��=ël�t�g���ͫ�ͳg���O)فɎ�@�F��ـ���PLe�W[��7��J��7S�$�b�H�j+<�2�ˣF�:����N~��٭�f��2q1֢�<��);�r-�a��׳/3�7�-f;�有7)ӑ�5Rw�n�{�,�]��_�nd��sS|����Q����V�fK�8�l�k5��4�>�^Z�s����tB��AUU!�%��\�`I#�wTt��Il�W	I�H�)V��Ձ�ŷV��,5%����`unm��r�E����Q� �L`r^���GL��\$�%%؜���M�F�Kg�n$���u�t�.��g��h����,��v�:��߿c��&�:`wumՁ�[�MQ*H)�rXk�V��3 I�`���}A�ߓ��v/:`I��*;F]e��]��`I#�wTt�$�����V�I�M�%�Mʰ;����$���0��{��)�V�R__�)P�7"pr+ �̖�l���ݵ`w۫��W9��u��M���nD�u�3�r���S�s�Mgiܶ���,v����R���(��`��	I>�~�7wn��w-jIs�wvX�ҝ�'@���^,����GL�� �&09�2�6�)J0��d��`wۮUw��|�^� ��3�"6k�J����	�C�C@ҁ������Y���8'�;�:p�F����z���b�t��0.�B����3)1c&�-��Ä"kb�b�ƏCa���h�8SFA(�o��7�v� �C&�@�s@8 ���(:�2�x�;@��D?�렚O� u_��Q�ꯂ�P����=Oી'.u�Vsv��ŋ��������r���K��}�`}����e��˫��v$��S�)�rXk�V�=�W �O:`d��.@*�̴Cn�YwN�&s���L���qH(�һ��1St�Du$M��n8�svX�c�6L�������W�%w��H�)�*I`}ӹj����nn�����`�ͦ�#��q))AIV6L`r\��M��c�К!:�AUU!ʒ��훮�77e������x=%�����GW���X[�5u%*JdqH�77n��� �&09.D��Sؼ��^�QX��p�X�M�6N�8K٭�7���n!���$<�\}�_X�����L��m�<{�6L`r\��6GLZ�EyQ����E�_�77e��l�ku�����ז���%��ַv6�) �Wyl��l����-��������6�#�"l$#q�a�{}���c�V�fK^�w׾v�W�7QD�4��i�Vpͺ�?,��>�~�r�}�xr�{�O��j@�N�
��l D4�"ҙ�����[/WK���h��<Y�э	�r�{Zu�[7;8�bZy[��q�crX+wl9�!�h!�`.z� �l�6v����^{-h6D'Y���[W��Un��IX�j�͜�R;˕�sL�kԝмv��N���ą�+�qƃ���l�#u�j�kl�a�u��Y����2��[�2㞻U9u6е�t�Z�B�>��^�w�������=�lް 4 ��Ng�u�0
�6{]:붸3����y9�=�T?%j\�T����F�1Ȱ���%Ș�:��q�y� ��(��'7DnK�{���ݺ�;�e� �3%�<��^��H�"�TrTv�j���r՞\�gwvXmn�w-G�"S�T��5q{��o�L~���"`n�遫V��3�*�I�t\����,俗}~���z����V�wo��u8�L�t�R�&+٤L����y�ۣ�n8�rZ�[kp�	FVf0J���"`n���6:�9ė?0;�����[t�JH�BUMo9W���9�@�~LRdA�%��̼�������>׺�̭�����7*��0�1�K��y0$��0
���G)��RA�IV�ݖ��U���Z��>��XCpB{"���F]�09.D��UR{ܮ��t�;$���:6��TjAGJԔ�hpFbC��K�v�Y���Q�Ӈsk��挗Mŵ^U�e�b`n���6:`�g����Ձ�smG�EE����0�1��6[vGO�IE�d�UG$���-~ �{����Vq.r��qB%��{�yÕy��Z�>k3#n�$�:�n������v���V���V˜�}��`b�[t��8�D�r8��۫��������,��囩��ȔII'6ˆ;Q�ø�ڎsvz,=q��n_m�w�۔��v���$�N�JF�����u`��`}�5X��V]��n�r�n
H4�e0�1�#������t��ꎟ�$Ҋ^��p#tF�;�V쎙��E�L}�cvDZu���*��.�vGL��vI�8��\{�<)�q)�!b�3��../��:��ۖ����J�����ꎘ�[�{8}sɁ�#���۴��J)*#�D�8�9�Άr���ZM��H���\[�N����M�U�	�h������{vGL�#�Un�I5D�D�I4�>ך�͎��GL�L|����,Uj�vZ�k ��t���+ 9����������r'Q��Mʰ30۫�lKؘ�:`����+����0�љL[%�9/b`vH���ʓ�_	JI{һ�<�U�@�8�����0\�v�j�r�#2%�Vݨ�u��C�l@��p��`�7���S���3�筓���.�<�[���:��^�aF�=����U�Rde1����IϪ�ܑ�b&���P�<ۨͷc�Ti��)�2�d� �F3��x:o9������qq\\�N��Y�sk���Z,�(̊�Ғ�\�?��7�a�~�潦��Ѭe�MЭ�� ��a�.�C�{;L�exw��RJt��M��;:�U��ݺ�;����ś����CW)��)��Ș�:`wuGL[%�7� ��D�͵NPE �*rB��V����f�$�{�K��K�x�	QTp��Ԗ������z��f�ٓ��WVUn�I5DqF�HM�`f̃�d��V�lU.֯�2�h�p��W�M�����x1n�����7m�/L���<݊�aZ�G �{<0;������ �١�n'"��NB��wU��/���r��:���cS%�;�"`vH�W{%'Q:Q�)!CQJ�1f�3������4�;��j����By"��F�W�^[v�L�0;������i+���qJI�`wwn��bt�ղ[vd^��b.�E�$[b���s͊��ɪ�7;q�nE�h�#u%p�ԕ�J�Iʉ�_��+��lِ`vH�W;��/*�^,��̷\)�[vd�:`vH��9���j���"7���K��xr�J����� _P�	�C D8&hv�~O�}~��X]�vv��Hn&�!�d���:`j�-��r&���q9(5nU��ݺ�=�Y�z|溜3v���^S��i�jT�=�\�g6��Of�U(�ʰ�r�z��bm�h��r�II�N�n
HPI*�;����م���Z��û�j��Gu	�RSuH�RX�L/��8ٙ�j���ڰ�2^��l�u�6�TQ��`fnڰ>��Vy$�;����٥���|�R�%HSMʰ;��V�ݗW��}�Z�H�qA>P��s�ʊ���H#��qO�M����zX͚07dt�����F�U�ie�b��/O�o�A	U�.��#)�l�z��JY�ܦ|�ēTJr��9>7�Ł��u`}��^��wvX�n�eT*:l�2���0;�:`�c�2��l��ۍ�GP��9N�+��i�vI������{<0$��0
�vR��ҍ�I
	%XwvX͚X���7�q/$�Y����ƌ��q�m]їy���07dt����vI����8������
H�)彧M_��:�8�k}$X�v'���=?'?��z��G��}HS��G�����ČĐ?�E��P�N������/#�]�����@����A��4K��s���L�؂~4�������G8JNݪ��]����ހ�D�'�ˇ���k��%-��0��c/%cur���	g�I�	)�5����
��^��ۧ����������n �����ģ�y���mSí�W<�
2�j�R0�.��/n:��^�n|5�Z�� ;X{K���Ͳ�X�����tmr�O��84�2���S�j��>����"�Pƪ�K�V��5aְ��Y&�PRg��A�<�
���*4+ԙmQ7 TJ��̼�V�.���u�g���@l�ˎ����X۱�y"�&a�5����Z:���+j��L�l��ET����J;��5-ɞ�/L�f�ms˞R��D�q+v;�@Ku��Z��k*�85���Dڟ#�`3ZWY��^���LӥI���̹۝7e�]MmdvV`��t�5������/"���9��2m�n�5n���.��ά������gq����.z�"�a�eM�!a�Ys{t� M�i"ػ�/��L�S����K� �9`h��И6j���$ӕR
,��K���Tv��Gh��SJmt@�l,��U�,H�3J�0L�MUR�ݸ�d`'U�箲�[��u��;C)�q�u�=. t���δ���Uv���"wW+�ѐ[k0:ѷ�vĹ��͐�J'=!�jٹfځ���Ƿ(������B^�RtQlR��S������ۆ�L�.�rtX��#
7r^�*V��t����i�tP=�ka�	�c���������l�`�H8PTl�MczNȻM��Yv�81L� f�m�qT��]v�A�9��YP�s���M"�p�Ԏ��S��䮩�]�u���6ܬ΁85��'�5c�aݢ�S��Z�f��ܔ3%:Ѽ�Աf�
��9AU�f,�&�v�Ǵ��m �,Gj�m�M�d5m.ɭ�0�ۋ=m�=;+=��V��	;vR�h�mYF��h
ڕ�Wl(ۄkN����L&5�su�/5m��̫h��g�V�:�b�������b�dxu�th��>�_uՎ�����t<���z�z�
��6x۫ob��S��>��j�M���@���4����=������ �W�P?�Muk��+��s���IP�6�ؔj6�)):�'�����r�ѻ[�y���u��ɝL��2M6U�*���`��.��ݥN�i�=v=�oBi#�d؝j�ٝY�����f�M�Ut�4�d�� r�6��N
mV���g��`�9�Ŷ�++븮�U���2�E��&Ѻ��=v��<gJ�tg!ٞ�H�*���3up01//^:�:K���w��{���?>�;Ol�bKr]�]^�UpAf�Z�]&�Gn�n7=oh΢'��jm��N\:d���0�3��}\A��ၺ�o��($#�nB������fK�����;0�I$�/��i�����誮���zXw&..7�ɥ���]X>�ԓTJr��9,��0;7 ������RS}�`M��i��1HH����y���n�XwvX͚X������%8څn6u�:����Q=x�Q�ף^I;7g;���N�����$�l�(5]}��Հgwe��{����`�si��ҍ�I
	%0���}�s�?���l�A�I��۫�RA��E/H����7%����vl�vGL{&0;إ��8
"E�,��,��Հgwe�󏹷����o��($#���,쎘�����{8�g�ٳ��7����[W��l�t	���jvmc3թ-`����u��=���>Ci��u�U�����Xw&�w'�\K��w7mX>���4ER��Ԗ�Ƀ �ٌ쎘�L���h��E�*:i�H��;����������6�4�� �I̽��*���s�w�Cn$�l�(5"nKܪY�{��l�;��v�I��l��sUR����+�(32��L`wnD�;6c�6���n=MF�M�7#t�A��&6�t㙚˝ntsm��϶*�B����r�F�qU�;Buq�7N7D�O��~��l�;��_�ʯ����3<��W	"�N&ٳ�H��:`}�`wnD�U}I�6�qR��������nڰ��,�8���V��l�>�9CC�H��Ӷ�}�`s�"`�1�����@8����w����}��ff��o{̱��09ۑ0͘��v:`�1��׺6H҉7*S�A�����ʩ]�Ft9���^���4٤v�;,d������vl�{�� �ɞ��������`{t=q&�d�A�rX�m��6��`}��v�w%��9�Uk7ҩGIʨ9 �r+ �������vy$���X�� �̢��N%%8�T��1��ܖ�w-Xo8�^�J�sޖw��۸IPNJ�:��>�1��v{��	��09ۑ09_U{꯺�I�*���U��7�`����%�KcN���K8�Ru���lN�r囅��}�_��6�N���t*�����&��{�5^�h��lu�uh��5:�m�����c��i`����3Q��ˆ��6�{˭�^���ÈMw&�R�X�C�ueݷeI�sA���X�:�M��dN����bQa�*���+�O:��LN�ءtĽ�v�!��.����@<�ҝ3!c�;5�C�g:�j�kq[k�6�-�dp�6y츷Ln+\�ER:�,�m� �ْ���f?��~`wse�i��)�����+���o��v�L�f0;ݎ��A�}<����������������K?�9��f���7=�`wv�#�A�HF���vl�{�� �Ɍ=�}��缘�\I�آ ԉ�,�6��3�����uXw6X����?kk͹�$�h�؜�f��7e.Ľt�\���z�Ѽ�Z�	�*�U(�9R'*"���wvX�Șf���W�A�<�@��~���7�[5�����?k��qUr<@�}��u���07�:`�1�͊ZI�#��)bqXw6X�m՟��W�q*�sޖr��`f.�9	E8�1]�0;ݎ��L`s�"`�1�i��@�����wu��,��w'�� �o�����Xsvp�N�$�c��v���&G�ƝӴ�s��.����7s�1d���'MQ*H�rXu� ����ͺ���;��iƠ�$#����?}IO:`}�`qI-����n68�5��36��3�����G�2���5�#
��q$.s��^�Ձ�wmX��r6���T�NEa�7�ݖ�wj��3n��۫ �2��S�INStH�8�����遻�� �Ɍ	�L�ߖnzF�zy�pI���Ż�Ȑ�<�rN���H�sk�q��ā����S%�_ �O:`n�t�7�c�Il	+6�JB1�F8$�X��W���=�|�v���S�$�;��4ӑTy���-�����Se�;6:`ov5`ϻ��DU#ddn���\O��ں���p�^���9_�	b!}��˫���j"B9$vw#��c��GL)��[P�0��	%$�K��T�������]r��ӱ��m���M�E6��X]ě��"A'+�7'�07�:`qM����� �O:`o���*jR�N(�IVw&��s]���-X��j��`f!��P�R�H0:�=lM��ݎ���09�Jm�$��Ԩ�T�q..?�7�3�Θ��08��`IR4R�+,��.�yL��L��Se�96:rO߻��w�t���h�%H�Gm�%����9�%��Ƌ&�93����Qc�%pp<�n�������g֭�.
#�.��͚�6M�0tW<p��1qv8�ɵ×��˳ˎ�m�˗̷W0:Nz5lu�q���f�l�a�{7\2癇`蔼]�MYP�
��f�|��qm�^ �@�b�.+l���sme�F(����&չ?���{���ww����|}^|�8���U*�͟6j+�%�����= [\+/'4imt�2��V�JvR���݀{�?����X��k��I$�����Հsپ��)#d`T����r�ٱ�{��{����H��H��XSd��$��͵`w��5%�U��Ł���;�06�M�I�A'*���t���A��6[�c�U���ۅ(�IVw&�������������X׺F4�*NS������h�@u$�>�qh���s�N;A��z���a�NB!��HX-�vۛu`gsn��M,�V���GR���7��}�q y�ʦ`�w�IM�3mX�4�?<�U�$ٺ�m����F�ӕ`no���M,�]{�Vۛj�0�1�l�G#��uv������`uzz��07�0
��i�JT�""$�V�s]����X�۫:�U���s�[X�xpC�Ӑuv��*���P��l2s�Gb�Om��9���L�
�_�®�%Jr�D��I_�o�Xݎ��ؘSe�9�+�B�0łW����t������-�ɻu`j��7 �q!�DRU��y���;�u�f�q��jJ\ <?b�/<V���w�%�����/1�6m����7��x����#�9���ω(��b�����qf8�~Q6��Y�iI��!�'�� `��N��;�~`L��Q�x�*N�l����P��d�	�p&�aS (����~��S �0Y �L \����W@H�x@����Ez��6��E4��ӺxH!�����$*!�(��W`�
'T4��Lם߼,�6��+3(Oe8I"Q�N9��6[�c��c�R�z��^���GR���7����X�۫{�`~yܫ�O�ű:P�r�pr=ft�]�;rj���s�9G���]'1�vp�HD�9MJ���+�77�V.���Կ0�smX�ݎ�%EPu�)M� �g������:�=l�y�{�ՀWw�ڌ�$DD)����`}6:g�Sg�0"��`wBF����ҢBI$�q������͵`u�ܫ	ăz� ?Z�J������W����uM�5�u�߻���f���~vۛu`}܃��m��NF�˥v]�L�@�bs�Vf�E�r��;u�[�#���I�Sr	��E%X������ͺ�3��VY�B{)�I�J�$����_�K�G}��`no�Xw]��;�^i+����q&�;���{��<�[=l�O[J���aK*�V]�j�~Sg�L�z�Se�96:`E�1Z�*�)^/��ۮ�[��'��w�Θݎ������G9�U��ܾrV��Sg�$���QP�9WO�p�	o^҆�C��jQ��r�\�Q�iݫTvQU�j":Tn�\nU�LK1��ϩ��#�e�s�v���]vʮ�HD�a�%^�1]��jy�v�ۭY�ۉ;SK]��6�E���ŲX�2�-����	������ў3)ͱA�?ߏ�۾3���3��]�:�ϰ�M��t���5�4޶]�^y}��{��I	hū�ݕz~-��AѪ���+t�.wl�<w�f{r����Ph�e�~����09�05we�;��iƣ)T��H��6���3n�]�v�3]���ۉ6�m�QT��7c����&�LU����N$7*%%X~�Z�|��=lM��ݎ�n�
�U�,�J�2�fe�8�e�96:`N�遫������ډ�F�M@Q�GSAjλR]��v�p�Y����;�۔I�7i˗�]�96:`N�遫�/�}�RmX�v�
���P�E`gٖ������	�TK��[�Ws��W&�L�&+Te�Y���mc�����v[?}�R[��Lo��Wf�j��$�����Xo�fՁ�͵`gwn�]�v�b�h�5J�$�F����;#���l�e�'I7.n̖ۅ�u�9����^)��doJb����2\s�PZ�v99�������n�쎘RK`E�/�q���zxT܂iĆ�8ܫ�w]����[�Vf�>̵z��`��C��T�7U"��J�5�mX�e�;ĵ!.s�U,%����9��}ʰ1{���Z�W	�1��M�a諭����)����0:����v[JʹA�Q�E�G*����X[���e�7dt��4P�S�3FRY��ڲ�+�vny��c�b�z�q�u)x�u��=G$MQ*JR/��K����y��5�7dt���� �lR���31#�W���v[�_|�'�����0:����I6}��m��9C		$����L	�3Ԗ�{�������%v�uQ�ԧU��s�{��X{�V>���O���D�@�A��]�˫Uwu
�r�N$7nU�ջ���v[vGL	�0'nK˼���-/'NAe������B�h�\��a����llD���Ҏ\5���w�O��l�쎘�:`vH�$R�w�2��/��`n��;#�d���5��m�:�j(��9V�GL�3�}��yI�`I�:`E�1SD�)���ܵ���{�`}��V\�{����{�[t�$���+̦[���Or���t�����C���?!?y[l������o3z�=��k�v]ٗ�
�k��}|��6�f��
bS62��z[�N�I�k�O�Aڑ�]�f��e�.�:�cn�x�
V닕[z�������z{7#�t�t+N����kM�c���q�B�K���9�9	�ru��Of�[m��l�<����f����R�]�jy���P�H;3$a�՞[�t�q��u�]߾�w����L�!�l,��+�:���K�wlGk�h��N��.�<�i�X�`�fs�	$��{��`gٖ���k�_�k�����]�����`��0'dt��W�}�L)=l͎�WdB�NRiĆ�ʰ3��V��vw6�����Xfe	��MIN����e�;6:`N�遽��H���)�SrH�q��۫{�u`gwn�Y��Ҷ1-�'N)Q�Q1B�2vkby������U��Xޚ��:͞{.-��u�Q85%X�۫;�u`j������d�j��+2�b�m�u�'�}ß�$T�4�Ȑ ��w<���]��ʻ�����\Ȭ�/$���$DD��`yn���ۦ쎘�09�����e��ffe�;6:`N�遽��U}U�/\���<J�$��V��)�;#��GL�e�;6:`{꯫�%z��d�@���xh-'n[���s�UϮ�E���q�2�ۗ��1��1�Է~�ߟ�y�-�l͎���l��
��̥$�MIN���]� �;�Vwv���7n��Zҷ���䑦�;��ʻ�����z��(B	���6xB+���w�*�w��*�p�du�Q85%X�۫�ݺ�1��V�.$�s7�5�v:h�E"r?Uۻ?�nڰ<��6�6��͵`ovi`}[������q�H��W�Ȯ�k�6J�}qn����E�P.�Ȑ	��#���`E�-����;r&6mՁ�m�G�A!$�;��u`N��͑�-�o�U$I��I+1U��+�`{}�Ll��n�`w3n�U��N!��7$nU��n�ʻ���r������E��#�
�6�y���ÕG��Y��[��.�ʼe0"ݖ���t�����ݺ�7+"t�ډ�iʍ�T�%(�̃Q�e�<P�.�v��L�S8��Nw �7��8����f�X�۫�ݺ�s��s�[�v���8�1��pjJ�'dt���}�RGg���'����遏���Q���WnZ�ٻj����;�0'dt�+��IZ3�F#y���v[���vGL쎘`f�Dp�&�I#�;��V�v�U����*�{�uʿ� /G�8*Y�
l�}]�E��[P��N�nk��bk\X�_�P��Y��'�{� O���/@���F���2�D���.z��?����E_t���2I	D��lGBmC`h6	�����E�����!

�� %6XD��&�K��;$����x�s��@;���J�� 8~�<��5�$h��4�4�a��y�����V����=�s���D�L���u�Gl��6åW�m��������%�����/����	��*nKj�`����+��R�F͵@[U���ev$�g�8��UJI�m�vU�S�Uq���l��ܘ���-�n����nÞYrZ%Ѵ]*�Q����e~���]�И�f�+v�,Z-��V��J	<oh�ۮrF��ҩ���^ѧ�\��b�l:�(�N(I-]jBUy�X���-VØ4ۣ Z��Kp[���a�ӧ7|�O�2�ԫ*dHհ��J���s�֩������b�&�����g ��k%.��]���Fn�R9�ީ�y���Z:��"�n��z��g&�gdͷnNg�l-.͌j�+*�흻m��öʽ��n��s�N�0���v�벵UU�������r��T�y��N�4j�p6xi^e'�I�B�&��J����RZ�ɫ��'t������k!D���M�25Uu����G#�X�k�iӳ�Pz���m�nN6Z����ȍ�tW)� �P9��{o��S���l�"��Aɼ�]E7hrE��2�6�G�?���0sJ V�6��%V�-���&��`kj��z���3��k��r	����8i˟V<��AN����C��dۓmG�X�����{f\C/d����Γ�I�� �,�S���v�;�ն�8�ud;#&��l>M���e�(Q�,i���ɺ����w=�&˞m�h�cJ��!�j����]�e�O)��f�v�[����z��U��=�U�L��|�(���֮���"9��і"]
��eΎ5�Ί�:��%\�]��Y�a�@A��d闄�E��l�*�]����m��l�1.Nun�U;c>��A�U��	��Ki���bU����� �(���i�U��t9���лhҴj�ԎR�T�m�	��]\�q)���p��������DO t�'u� ��|q@��@�;P �Pv*B	�C�����h����]����%��el踚��Ɖ\�	zt�%�k9.����۞��h.�׶��:y&I26qu�-��pqFm�����8�o��|;D��-\�Q.X�7\=��u��M��s`8Ův]���9t�ո3۬��9D����.������m��ᵞ;���I�7+]]r���]����,���tR8��l'��w��s}%�p̗��6�p�S�\��g�䛗s<���/m��3=�MN�&ĆEMTr���Ձ�ݺ�5fk�;��V���N*MɗyL쎘n�`vlt�����_}��fbȉ$
�EJ9��3j�������/o��7�t��)i;řu*B8�M�`��`own���Ձ�3]����du�Q86�7����0"ݖ�콉�vK�\3���q%�dPk�Jn�����Wg�l���-�(��:���uw4J"�9�YWk�7=�VRK`v^���GL�5KJѕ���yo3[�ʻ��u��W�O���4��p�x� Ρ�������t�����#v��w�,Vfffe�7�<�H遽��)%�&�G�]���Uj�Yx�H�߳-X�2�7��I'ݙ��ֻ���x�^*Wy�fS{#�RK`v^���ݺ�1n��=�JA��7�(�7Ruu#πV��Y���m���=Zs�v�]�3�̫�Y���GL�ؘH���9���wvՁ�״۸IJ)%T*S�Xew�\�f��;�j��̵z��ٽն�ꔢ���!UQ����/w�9z!�	t�F�w���^�ؘvLV��2���[-��}�L	$t�콉�$��vj�����Sq���X���s���3_�7wn���Հ}Z�[�8�t�i�=fm�s�0�[���J}�΃����D���<݊���0��nU��y���ݺ�3���H�7B<J�T�b�U�����GO�}�L	'�0;/b`qWt'q4�܉IVwv���ͺ�;�5Xn�ՀVfP�J���S���/����xr�~�~�U�{��¯�ဉ�*��������ʼ��u��	������Vu��ݺ�3��VfmՀwr�&���g���<���#�h�y��-n�p�on�P�g�GRG#���`}��Vwv���ͺ�;�5X.����������M��?��}U�$I<遾����� ��V��)R(�����۫��U��\M�������ܶ�U	)��U�Y��콉��#��GLݎ�t#�J�!Z�j�Yx��:a{���ʽ����_��{���W��Q�|\\�j��ڕ
$�N��t�rb���jv��&+!:li�f����c�n�����sQ@[�Z���`��ژk:�xV[��T��`,n6.n^	5ҷJgOPg���h�C��q/LX�/�u<m]j��`�V0k
�G;�F=�z�ô�b�FѤ6��[g~�uȝ�ug��F3$浰��m�m����6��K���[i��,��� �?�w��s��}���W3�>Rz\ZKV*�ɫuu����I�8���u�[�#���͵�a�w��e@9���wc�e�LIX�z��!�(�$T��X�r��.qs���Y���wmX���qq��ݦ��F�(�phrU��{�`}��VnmՁ��u`nVm�J:�j8���&$��6:`n�t��U}_|��y0>}ݎ�"����YWk�����c��ؘ�:`n�

�;ř@��ݩl�%�& ���l�5�\Xwn�U����!{sh��j4�%9Q(����w}u`l����#�͎��E,.�U�u����^�^�9���'��,�|���GLݎ�t#ċ�B���`��09$t���韾������y�|����Wp7�8��܉IVwv������{�GL�v�3(Y�eQ"����{���]ٚ���ڰ3��Vݧ��\m�9��8�k�6��K�-��y�9Ƴq�F�+N�6��ƥ(�phrU��y���wn��������V�͵��)ʎHIQ��:`odt�����{��b���*Q�~�T����V{ܵe$�k�C0	�d_@pO9��|�����+��Zm)NQdI�Vf�L�ؘ� �����ѱ�,.ʻ��e%�L�ؘ� ���遙�u`}�7�l��Ĝh�I�]<��xF�yٮ�X���7o��Y��'9٠E��j�Yx�� ���遻�����]��4�i�I�p�3��V��L�ؘ� �+whS2�y�+3*�e07v:`v^�����Vٺ�l��JI��%X~�W9Ovf��٥��ܵaՋ�Ӈ.	�KB�����y�ʿt���ލ��oX�0̼LI�`ow �����{��r����>q)IJJ��p���6;7<��lslP������t���=MBv�����x^3�z{?ݎ���0>ݚXwqkI�S�E�fm���&$�07���ﾪ��7Bz�I��u8�%%X��+�٥��ɥ���u`op6�M�M�UV$�07��`n�t��UUK�������q4�܉8XܚX���~���k�g*��nU�K��Бw���?�{
��Uul<R�X,��L���\r�A�E��)Au�6���ٹ��Ac�n�lP�d�+[j�;�%.�x�k��nq; �V����j�&�Nk�3��9�=1�mV�%e�2[���Vۣp;�6]9f�බ�N��2��]Q��!�Hzc�5�����.<ֺ�Bhn:-�m�m̥@p���sN{q�����<����*a����i~��2T� ]��#��ym�Svh�SYe���5���<k��Z�ܗMث��	\�V������09&C�W�WM����SV�8Ԥ���9*��^j�>ݚXܚX��V�l��:�RBe�`rL�{���LKؘ_fGMTT���P�g�����`ffڰ?ew���۷��-�6��E G,Ĳ�`n�t�佉��2��
�����D�J�I��JP6D�Ψ�c��-j�P�B�M�{����]�v[Ys���%%|�� �Ʌ���P��u`f�měn�n&�����viu�S��+����>��u��09/b~��:�4=ƜM8�7"N��fmՁ���`}�4�
���B�6���I�07v:`r^����6?�MZ �JR�F���y���+������ �3�wc���j����:�2l����\d���U�^�7���9u�<�MB����FFI ���vi`gri`ff�{���՞�MQ)ʺ�x�^��fx`n�t�佉��٥�V��j!ʉE#����uʼ��r�$�� �)fXG@1��� ��qS�^	Ȉ�9�'8��Ё�n�G��)����k��*���.)�O�QB�^'��2�x�&���m0tӰؖ���.��-G�ͧ��<Ox��������y�4�� -k9��C�@�[����m��C ����xp^ `(:PG�銨࠺u�X_�W�|PI ����h��v�f����U�+��s����UY������hͱR�mS��))*��^j�>ݚXܘXy%��3+{����UUQ�Pr�09&A��܃wc�%�Lm���֩8vhѱ4����܌n��[�j׀��]����,���]�#�@ف�܃wc�%�^����T���(RF�RS�$,�۫�y����0�;�f�$�3uk��T��$�we�S������rݎ�ݭ�F��Q��H8�>ݚX����^��xr��d��#����a����^}�U韾�͖�l���/��Ƹ��ၻ��-�lK�X���9�v�6�8霡�p�Ȃ��x{6^z\^���.�'\��ፎvb�*n�I�7bX�K/$�[���"�{vi`w�ͱ�
�j��D܊����^��g�[�������{��[7�q����j���`w��V�f�fmՁ�3]���oq4�܉8Xz���^�?	'�0"ݖ�� �6��P�����RHX��V��v��{�����ܫ_�"�1�����o�c�(Ƹ͉3�8yZe���[��bF��t�E�9�Zug6���vI&�ͤ��)w\�.�W;��i��zv��8�U*�Bۮ���;��vr�*�;\�5�׮���cvp=U.0.�.a�g��\;^#�ٞ�1z�X��v�ݓ��Fwmu�.���-�x��0�g�Y9��z"�.s�=-\xI��3�4,��m��DF=���w{���</�H�/G8�ŎeZL��D�2�t:���ۜ�,#�9��C��QQ)D�6ڒ�]��`~��;>ɇ�ĒK��m���n�u*22IN;�y��������ڰ1��W�..6|�n�"*���?U�����07�0"ݖ�佉�V�-i4Jr�QD��`gsn�Y����{�K��6�J�N��L�[����09� ���t��'c�t���l8c��\n�l���p��NB�۷陞ܦ�ڴ"��N���%�Ll�07�0:�e�8�07�8�qRnD�VٳKʪ�Õ�Q�A��uD�-��ʼ�}�W��U�V�P�J��Ԕ�Rw5���-��{wr��j�/���6ڒ�ך���7&�w6����m�5J���D���ob`l܃{�� ٳ���ꥻ���[u�qk`ȸ[j��b��,C������R9�zN�8ӏ����]��l���~����{�� ٳ��0
�b֓D�*%R+;�u`����^j�3^j�;�3lT���q��u^���y�{���;�8 ����C�A�6�D�*��V{���7�q&�MS�U333��06^����t�6l�ʳxӉ�&�M�`f��`z�ʯ��r�6{��0�l�r�+ʺ��Ţ8�BEA��7]�{G����w�ΎP�X�b�:I(RF�J�E`gsn�{���09/b`l�N����RW����`ݘ�����&�۫���8�Sdd�Fܖ����&ݎ��f09K�(������<Ƹ}sɁ7c��ٌ:�	ь��Q0H�e�@��� ?"<\�+���+ ����%9Q(���X�0?UVܞ�6����܉�ﾪ_��?��H�<�Vڇ��r��������e^t[m�zfg�9�جp�z�̮�O[{r&6�^�ꪪ���Ձ���ěm5NT�Vu��r&f�L��O�_$uV�=���ӊ�p��`w_���6��Ur��%�Y���ku�����"nT�JR�T����I=�`l�����r&�V���JI��$���U����uy���^��xr��lQ���o{��{{�ߝ�m���:qY�嫟Y9���ls�O�:��6�\���)�fV��n�/c\<� �9͡p�OEgNڍ(�̅@S�W���n�zLP�E�۱�e8G��ŹU�{=#q�����u��kv*��U	;W\R㛓���n�S��Jg^�M���L;���j��\�p�cNx���Skv9�Q����BӦ�9�������\s������������z��])=��ܔ��ʫ��<�X��n�m{u�ϡ�n's�ev�U��\�8��������>Ǻ��۫��U��Y�)D�Q����忀�yX�0;��08���*lRҴe^V%�Ėb`n�t�������{����&46��#nU��y���ݖ��܉����;�%wv�Uኲ�/�{�r&7c�v�U����Vn���&Ԏ�.6�q���RV%%oK��2�,�Yv�y��A�NV��0��n/��yX�۫��U����`��
��J8Ө�Tr+;�Ó���*a��+)2$HZ?l��� 1!��/,ֹ�r�~׿g*��w��7�Z�QbN8�G%Xǚ���&6�L��L�Q���UٖffR���佉�͹{���{���4P%J�Ŀ	�_�~�1we�;��09/b`~���RU�r���'�#u,s�l���[9�"Ů;�b&��9t���M\� ���#@Q�m������;��09/b`snD��	�]M"rD���<�`}�5Xc�V.�{��D�i�p��8�>ך��=�{��AE0�+�m{��u�;�5Xך��N*t�F�>Ǳ05we�;��09/b`�(Us)(8�%J�E`b�k�;�5Xk�V��U����f��S�\ljF�(In,(M�Z伳kΚ��۔4��НjӸ���8��SC���q�k�+�y���6i`b�k�;�͸A�R�JNGJ8�Kؘِ`j��`wob`m-�)D��_�寀��x�1w5�ǚ��� ��Z�iJr�Q(�a�Wsj��Vk�?ew�K�.#��c"��
�!�Pğv~���vƝ"��9#�%Xv�&%�Ll�05we�?}_Ul��:��t{4��9�]<��os�u�Fr9�q��\Ø�rs��B*��:�c�������̃Wv_�����<�okΚ����8��f��Y�vr�]���r�x���}���bn)�++30`E��������-�͙�kU����*GN8���V�l�6d��`IP��/.�����Ҏ+�{��Ww�x�����~�9W�"*���U��AE�AEqU��TW�DEQ_� ������������"�"�2�Ƞ **(�� �Ƞ0�Ƞ H�� �* ��Ƞ�"�0��� �B���(,� �
"?�AE�E�DU�U�TW�DU�Ȉ�+�""���DEQ_�E�DU�qTW���+���
�2�ͧ?8)������9�>��     >�               �   Ъ�D�P�� �
*R�
� B �P�IAD)D���AJ�   �PA@ �US    @�( ���0� �z}.-�o�y�֮,��|��+� 秭�y�}���7=j�u���ҽ����Vo}g��^ y�0=>w���� �����`  "  ]��>}T��g��o�����7T�ܚG �x      3 �>�n�e{��ٽ��z��qj�� )� D f ���P D�S�ܠ`���h�z  Of �F ��s ����� :b:���OGG�  f���H�S�;�
  
 P 
�V��)OF S�N�9O@��OA�fP � �7ϔ����u���.nN�_=@$�����������7}�w��o�nW�Ͼ >�[�{�/�y{���������o��%��V�ҖM}z�{.ӓ�[��  � �f I��^��������}�W��Z}� wS���Z��k֮}�Ks��� U�*�z:rk�oy��[�s����{ʧ/.�����_|�ޕ�Y]\�S���ϯ_O}���������N�� >��P  ��{髽ϟe}�pK�{�����Js��ɯ�O������Ү� ��qh�O_ ��+�}�VpM��r}t��q����W���y^���
���-���c��}��糥^ ��*oi*�  ����<��R�  '�URM�E  '�T�JT @�����J� 4ha!JSH�����~?��������w�Ώ{��� *�5?� *� 
��� U�@ W�UUX�������H��f�����!�����A� J[��ߞ3=*��!p�-���ɇ���RK�t@�h�hj0H�$I���h�O4s	K)b1��Z���ɚ��0��A�*�@��F�,�3�zM��\�9�a�i)���Q� 5�#FE�H��}##}XL�V�J�H8� ��J�+J���8�(K$K��Z`��BR����k�{'��E�zrf����6!])�@�Bc4�aF1"�$ E$`ą50�S0HV��z���":0��!�F�~Cy����\�S���������=��3��=`đ H1�BRf����\������eф)��T��@�"��
���)K�HB��m�&x�\v\X�cD� �
Fup�f�X� ƌH0��,�d#s�{�3��y�4�ȱ� @`@�T#� E�������R5���� �lJ,
�H�����!p�)��x������2k�ɠ�=�cp=A�H2&���$Fr�F��,��c��!	!2M�#��� �B����u�y-���ss�+���q �@�H�1�.Bp�� ���}� P"R��e�B#YI@�$``I#$X2�ӄ����(F$*�'�E�I#���%��k5JD!$H��pc5��Vh���i
±���R�@�H���H����9fݳ$��x$8�b@`A��C�,`1�F,c�.�
�WBc#2���4��HP�
P����!P���e�A߁$x�f���74�l�.��S��C�]��o꫋�ձ� N%S�������!��v�©�!\4l#avK(B�+ ń� �2�9�<�HC���J�Ő�#�"y<!n������
͋6�� ad�0MI��w�w�!��p����7�x������#p�rHĚ"P���!s�p��bj'�!RH��� Á 1)� ��`�d#"	C	q�0�DRJ� I������@0r%��IH�&i!�A؁�h�=�L'���	�5�pѽ��xC�)��B$��aR,2�C	�����9/�r$�a.2��K�cR�p!L!sC
9����u	5�Y	�z]�gLM1"�,F0#$H�F�f��5%HX0	HHD�RFF�,�	3N�d�ѻk�mIv#@����=�_5�jJa
����(b�bd
$ @��5�B{�.oG_yZ���B�B�ń-$0�(8��g�!
f���h�F'�%�r@�Q�@ �2���@�C��SZ������c.a�kJ`ˑ!)�nHL�h�B�tJ���!�,)-&B�$�H�1�"IB!F4�ѕ���HZ�+$�ake����2��Y�.�a��B����0�L�}	xB5��!B�x{�����3<����֤���+
Ɛ�nB�Hby���{	�H�n���n,����#cB
H���.kg��k<ibz83Ӈ�xD)���0�H�#L6�Ƭ*��D��bP��6�J�:p����f�y��ĵ"�$RaVP��<������y/8^p���{9�!�5��zݐ�@ �B�D��2=��9p%��I��YVP�֔�%R����(L0$I��Y6aahB� � ņ����!fd�-�]�.�ם9p�Z�����ư�������h�ԁ"�����l&� �$=%����xŤc��熎� l|8h�a�3�Q�F>� �l��BW0�ћ�.kx��73l���!#$! Da$H�F�0�e�!�<7��M�tz{CQ*ĉ��t���k��h*a��@��0< 0�� �)8A�R���)��F$�4��!�Y	z�8޵����:���dP����i��/Q�m<={
a���< ��4l&�R$�D!�|��G��I�
���$�F$ 1#���a7�{��y��]A�0x$�X&�Y"D E"�	�b��XrB0� �H�"H�d�cBXFf"���`B:"Q�  V"K��%��
GP#
���h0b`bGBW�$:h��F�iu���4�a.��ozk�XFJ@��	$��!�,<5�I��B�,hE�@��2�2q�RGF�F@�A���a��HG�4l� RbQ��%RB%����4K8b�2	�8�%)!$�Zf��35I��6��K��6b��	
0�+0Y�dF� F�!!$�d�	 ���y ��Z��@��!� A�E��C��H(��  ��� �b��
D�Ԍ�D����c	 �$0�K)�ro57��@޷�4��a��1�
D����]����8�/$��
`@�D$ۊ@�"�I ���$"Ń�s�pg3f�i%�D�5��+FSfof��+�5�a,� F��I0I,�h�@� �W��e��B��k�7,R�	\X\H�c	�����$.�2��4�&�3��;�2I��
�����́�F�0�lk#�S���0i$mŅ�!<���}�K���% �$$!g����ݚ���谺���*Z�1!�
�8%�	�E�l��$�eH��IaF����7�$���SZHC4�Bd<��d_9�כ)g<�3Dl
y��5��e�d֍G!�癡��^{,�[m������M��Ύ��|d���mX�$�XX��aT��a���y.i�"�%qHҦO|��!\� ��)$�!#�$b�E�"���#F�UӁ�
0�i�%H˹��:��#���!#��
G	v�!���v0c�$��FH�N�J�G"A6l�$�A�w�)�@�.6d�;�m�kz&��,�{�"թ�,��Y��<�h��=˯s9��7 ]<=X�@#%�l.:$6���!YR4"IV4�!Fc,�6/&��#Odٹ�ݝ�;�F��<z�������RRQ��9M�B2� GL�Fl)Oo�Q#$��i�2�3Б`�<h���Fxi7���,��}�pH�$�!WX��,��M���j0^�
�#Ej�F�ĉ��$*`d�C^�|��RV�!R$B��@(F0* @�\� \!�iH��'�4^y��I�5�]N�l�/�2_3[.�0�#;���P�"F�a$A ĊI"ł�J�H�ƒ21H�( �I,�FI!�E���B�	#"B��F,a#@񅄒�E���!�$,J�)"FbH2,"�BB�A�K
K#{�������| � ��6�       ���   �    �          ?�>                                                                             ��                                                                             �>    �lـ�޹dlm���q��	 /i+l4R���R��3��4�$	���Sj�-�Eq,��,�6Cvձ���Mv�	)@ �[Ku�m-� 2VͶX�9�v�e9�Y]�Zꭨ
�$�� -k��Ӧ�[���9ݩ[ �*ʧ9k�9��m���V��)��]�s"=�*�V�.ʹ�U%���M�k�Hkd;j٭ko .����ۭ��)�-���cU��� mu�� �|�5V�T�p&𰶻m��Lf��sd�9��[h��6�	 6�V�5��m���Hb�iv�O�Q��v�YP j�U3T�U]R�t��� #n�ޘ
�Vd
�%*�=m�R�Kr�e�1��j۠-�"��m,b�m�,�Fݛl6��$:�v �[T�6���T�T�  R�P�/H�n����Ja�ύ&���n�-�� � 6ؐ [m����I� @�M��$]W.�k�B�vZ3��Mzӆ���f�$ $�ӆp�c�� 6�M�
Ytj�]�YV��V�Z�Z�jyZ�vU^4k�V� .��AK��8l5*�PVؗq$Z2<�P����QΊ�ܓ��6��� 	�vm����A�k��W.���轖�z	mm�M�]cZ8  Pq!5B������N{
 p�b��j��HUR�@6Z$ m��Kӹh
�*�VRY27uK�-��`�n��w[%���)!�L�@b6��8&װ-�z�Նm��/Q�H�lm[m�rI$�u��(��m�sm�hsnYͤ��*�]@=n��RS��&��U�.n(�	 ���V� �Hm�m�X-v [m����l �;m�� m�$q��I[ ���;�m�\��m� �l���/0   0kV��ֵ����6ܵ�Ts�\-��2ղ�k{l\�m [m�v� ���f� ��Z��a�n�k��r���m�h�`0 ���a�lpCZ�k5���f�Dv� J[@ a{i��ݳ^дm&� �$ ]3h�sS�� �e��n[j��y�������)�V��p6�S��E�T����v
�$M-  m���J� @FcU����[i+j��Y`��3	�V�It�m���D�6��Hk�MoP�\ N�&��Kk��VڞZ�]��� �(A!o-��H�Ʋ���HNl��-�8۴��k&[�DZi3m�ݶK+e��Z
Z�k�)��j]�m��@ぶ͎P �~|�g��ɭ�(Y����[|l�]q�[RrE�d���MwY�m  $�^�lH勩zMs�鍤݀6ݔ�U�pX�mPUskӒ��c�v�^��m-&G�z�6��g��k��7R�6Z���Hv���]iYW-mV�Vm �nn�z� ү��}�TjnV�V���]�l��%4�Xbz����m�H� ��0�2ԫ��V����-j�1sEp[B��^` 6퀐	�����[\�o�6� �ػxҭ�qm$� h6ٶ�i��vĲ� 6��m���ݶ�`� l�:N��P%��	��i�v��N�J  m��p �����m��o4 �UJ@f�jc"�X����U&`���U�Tʴ띖�r�\�igq\�S����{i\F��Cu�S�@z4��`$ 9 �m�`mm۱�m��H-�6�$�� &�	�`	 8m��cm�6�m���m��-.�-�� m�m�|$>	  m�p$ k5�m��ZkT � t��ԫ]UVԬ�*�U*��U: m�`  v� ��ml  8�����)!��  �`m�� d �f�l-�8�-�Cv�e������&ݱz�A �]fvNCX8X%UU+�'m�.�� �� �	�a��  �ɬ� �� �^����hm� � Hm  �  �  [I �"B۵ӏ+m<�U:(㊥Z��iM��	 ʜ�+J� 9�i
���  6�  m��n	&�H-�j���?��85��m    ��q��M�֠0�*�F���R��/l[m��6�m��  ��e�Ue]�b�vWDm"��bMn���im j�m���"˚`7eP*��X$&��U[�k�%URP [M�6mm�.�Hm6�[m�h �TQ(8܊��uIu�.��4�>�['�|�߀m�m��,�m��mKY�z�[@�6��M��&�vٴ����	2&հ�B3h ۃ��e�K��ɩ̷'tGK�d���/��<�L[%	$p-�����$ q�l��:��*u��UUU*���P�	I����{d�e��Z�,��9Z���J�P�wl������ ���lt�,[G;Z�Z���u�=jWf��6
�Z��q(�V����8�ַ�(~�k檪�CҒ��s�� �h��]>� R UJ�]U���@U�.%H�`�  �� [�� �  U���n�j�i啨
5�.ٛm20[@ H ���nDF�m�[A �`�>m��m�+r�9@�FZ�����    $���4K��l6Ͳ���f�6�  u��)�Ď�\��Cm��T���k���Zp�j5 �U�U�@n�7l��@�m�Бz���f�m�6 -�8t�p  fٷR鹁���-��H  � j@ pH �j�����nʪ�p�UR���V��w�>���m�� 6� �]nH�d[)l:��M���mm����孷b�m�@K�-ɪ�����m"�ԫZ��jYWa��E���/Zm[�Hp   ��` +����Z��jtK�T8-��,[Y:�6ݓa��F��l��Ut�Fհ��M&�n�k� �qc'Ǡ�+c�-��u�W��.B�â�\B�ۧ@�4�L9ct����Z�g+��@�Xqm 	[v��M�f���i7�h��i#�$n�X[Am,^�ԷkX� ��]*(v�-��kn�l��m� �  $6��qoli{J��@����� ��(_�|�� �m�)�v��M�%�����l�Լ]6$� m[6ط$�r� 2:@� � ���l]��m[j����[@�J�m���m�-�%,j-l�ki  �( �]��&�n�I���v �		  	�\:tl���I6X"K��Jkn  �Iԣi6p�az�m�m��@[@v�Rō",���[U]+�n�]�s��UR��K�&N�S*�0櫓#Uz;mW;7RHb�#[�c[W��qzٷ\ml�UUeb4��j��@�� )[lv��c;3�#�vŰ�m�Z� ��]�\8�s�UJ�˯T��nf�}�?(�rp���� ��YZհ �[U�*�
�R%��d�����	հ,1m l�@�аoi���>I�O��i"��m��� H�mz�m�-��kvۣ��� �M�.{�=�Z�e@|��[Ŧ֭���3���-�%��m�� �� [���-�YD�� [C�8  ���� -�lp $v�wj���: ��Zm�H-��`���m�[d�nۃ���6�~lm�� �	 �8-��0<	�A��[m��vr���v� -��9b�m� �`��%t�-�� m��H �m� �J ��u+�ڬJ��mUAMl�I؝d��i���n2m�n �`H  �8 �8 �٧�l�6۶�]� i��-���izj%u���UR��㟾 
������tݒ"�+�P�i$�@@�5�ʳ�W�:�Z�h 6� N���]�dmq4WuT���I��W��l��+b�����ٶ�W;�>���{��T��Wi:���P"�!�
:�(�j pb
�J��"`�x��!�T	BET��x�u�P���(y�`�4"'��_UOT��$����A|Wщ�ٳC�Ш��t���SJd=Ҡz����q�
��S@U8/= }zz� �<�j#*z'�xvz��A�ߐ��A�$X
c��")@آ.S`zDuJ PE������oQ�@`D=D�=v����GB�b�i�x���� �@|U<:*`	��D��v� ��QPGa�T�L_Eਮ�"	�Eg:�AE�;�TІ�SJ
��_I�����	 $E!8�:�\��}T:
TF �N��`���UO4��O^��@�����y�H����Ћ螊=D���h��6!�<}A���A�<X�^����)�����mi�!���zo���y BCJo��Z��!�4O����> �'���� �`/�� ��Q��&A� 
0@�*%J�@��KU,EO��ffkZ��i�����              l              ���&v�筱�٣
�MrFy;f�ٞ����η;]C����j��)����	�n�ܵiN̹j�^ɒ��j�;�����l5#Z淍h�"�r�	*���jn8�ss�қ	���嘍��\���j�ݥ(�nB�1(]r�m�;��mU]�MÝ�k[�7aŋLo�An;9�R7#l��m9FU@�l�p���� ��`�30t�J�Y�nm�n6�+mr�c;]B�V���lltB�N'�8�R =GGC��\Vl�..��,�ڛ�{gnS(u���mЛ�a��RvI���{N�::8lJ��R��V��횕�.x�"�HFH�	-*��f䊶;<R�j��X�!�vu��,t�x����-��Ύݦ��X���x�%`*�$dN�s�7[;.Y���`դ�F���^����6��	�` ���(�e��nګX�}�i��Qm=JknS`IJfwl�v�SlK�fa��Mс"n�r��c�GFm\�b�G�٢�8e�,i;a=7�����mܙwn����T���fx��kqul�+�U;��c�wlX��̤����ce7Ő��⸖�*�^��s�8Sh'��î�#�#sγ
��bJ�9 .ܵm��.��=u�ʁe� �ۥ&;I<�T�K�P�.4D�;�w�Jͽ�b+�^yig*tl�r�d	�J�c�C=Aj�l�Kn1e ��&����ey]R�8j�Y���{^L7nY�[�-5u�9�l��ca#�1��]�$u�슙�gX�kv��*p+vA�M�;,�Ίh���#e��u�(9*v�Z�����ۻinx-�� �\뗲���5�nF����I��85��7�^�PV���d5u��֨MkV�d���-�ȏO߇`����?�qC��+��!�'AW�"x�OGJ�Q��wZ��շY�ր l  U�ȝ4���N�	�:.@���q׌��N��f�� tt�+�]��=V���J&mQ�o@����Q 9��:��a(ɂ�$�&�4rg]l ͇=�@�c�0j���$7ћ��t<��܄��oE��lP�b��p�Z�����l��o\�����.���O�r'�'�Й�o{���w{����t�y�y����K��.0˗caȻ
�&�ȡ�q���M�`�3�M��<�j������6wv��$���0���ҞG$"�	�4�)�Umzם4�f��yr�2D�4��巬Y�0mL	b�N�j��q����#����4�)�Umz��Z�q19�6�m��,T`\���K;F��?�������ڱ�͐[v�_n����͵n)魕.:3�(ܜ�=]I]��X.�tI/����巬Y�0mL�͵f�&A����k՞y��8W��] (dAqьp@j� 4T=A���'|�97$����^��?.���c�4�F��@%�� ����*0.[z�6��s�L�<�F��4�)�U[�JD��\`wuM��]]�sv�ԓX���m� �v��S	��_�~�@:�k��T�:��s*����ؔ��{p��#\����瞛D�F��p�o�M �Κ�hzS@�;1��j'�CQ�4�:0���Q�I*`}"��B�LNx�M�@?[f�ץ4컞g�<Ą"�Q�1#Z�D<�<̐�����@�ݑ;�$���tI&�Q�I*`�р}m�s�ڳH�Ả� ��4Y�0���,T`�-I$�-�0�<)��ԚŮ3n^5�z�-Ղ�mͰ뗜ֆ��o���h�>���Q�I*`NL�nw�By0y��@?[f��$_���o�@:�~��
y��Lx'$�5� 7u����Gθ�����TW�#K#IA�hwY��s�rI���܏ʟ#Ċ�	�0U�G >޷�ܓ����2Y�!�ܚם4��hzS@;�� ���I$�a�11ŉ���N��"D�����+�5�H�_#Nީ���XG�(�p�z��Jh���	/��\`o+��Awvj亵Ԙ�F�m� �v�ISs��t	"����mzo:a�!(�}xs�0��f[��J���s7WX
!L�:� }x���� �3�:��a1���n�^�0�۬ ״��J�(�����������ն�      /Tّ\�e.����� �TUm�i���ŭ��y�b�<s��B�C��v��㵷a��m����y�����#H�4sp��k5��s���A�ի.��n_(J`9���]vc�mu����W��*ҺGj��B���q�[IӐ yÙ�M��q� ��ݻRm��m�:��_���M��Ƙ�ߝ�������{��|�:k���9*Ėq�^YX��6Dܱ�n:�WA�;S0�
yi�0x�rP>��Ɓ��נy�@=�٠uh�\"��,�%����z�%�� ݵ0%���r��s#OƇ�8��:h��4�)�z�����CP�&)Q��0<�)����;� �~n�^�4�܍�a����&�}v���z�,�� �*`{��'��I$,K��TY&����S�J��,�j�\ c��F����^��5�mOGB�ܡ?$�o���X �i���|�!/��|`t&g�&�**j՗5w�v���"!H�!~�9$HH�H�!!�l2F$$X$H! AdAH�1#��:EY*<��W!�^�u����IFf$�~yxbO&Q�h���.�F��0'h�>���HX��������IOog�>� }Κ���V������"Ib��*`{������_&ڨ��@rn�����^�*z�nR�-��J]�K��V��������֡��&qw�0'h�&ʘj� �ʘ�TUB8��A!Hh{�h�)��Y�^�M�vF�0�@R
n�j� ;f ~z�V����DD%�fy����{��;��ݞ���ȒH`[SȨ�$�0.�F^�J�ǌīNM�Jh{�hj� �ʘ��ԒI . ];X�OTrj�^���\��t�˶G�d�X��c��1L�F��Ƀ�D��Y�_l��~�f�{�4��zHH��L:�����ДDL����n����߼�/�g�FA��%�8h�_&�Q�M�0.�F�����s���ܚ�����/�SI§���EDr�޷$�gu��2�8��A!Hh{�hy��w���߯�@�ҚGu�I0MA"H�i�$!�L��[.�yݎ0^-�:�XMv��s͹�#��(�rh�)��Y�^�M �z���m��	�L�I��0,��l��v�074�W�0csӓ@�Қ�����h��hq���<1'�����M�0.�F��0,����e� �(I��$��)�}�g������wN }�� _�!%BJj��t����ޝ���;�7�      X����,u͓q�n{g�E�l�筶�9� ƨ�m��=�";mh�L���z�n6���OH�vӹ��Y�x�m����W��)��+�@�=�P�#��j1��[E�/_/ոIW&b#vG�b�Y%]Heզv��mE�IH�L�b��.ؓi�0��*.�;��l�py�[�n���^�s�Z�����=;������[��4�2\��$4�i+�;d�
�'�pp���4n�]����82dI,Q��_��/;V�{�f�z�h�u1$����hj>����� �*`YU�����5X�#��C$�@=�@�e4�[4�ՠ~�����
D�K�I�eT`KS�یd��5�m�a	�L�I ����Jh�S�T`nm�I$�pIf!u`+�;�V�ڸ&�ڵ��j�vsm�m��].�Y��R@J8�Q��Ɯ���{���l�(_��u�Kb�u4�&�N����O=���D�D�� ��iH��0u��� �ڗ�D�(I��$���h�h�S@=�@�:����X�� �Z�EF�T��UC�1$����hj7&�{�4��4���l�-,,�I&	)ԍRu�tn�����[;�W��˸ 'u��6���`m�0�H�NLHR�u���h�h�S@�ݑ����	ĔYޤ��U����*0���~�f$Z�m�<#$O"�C@=�}4��78p}	ȅ2��Bbw�xlw:
O�D���A4��UHp�ۏ�@�2:t��"c$ D�23)	P��G|G@�=�@H,HÀ0��8΢E>Ho�_���j��Cg"���"c	@@oD� ��*k��m�Sk���l�-�����`mxJ�3ͼ�ni��@��(�*P�X��RF	��6���FS�� 8"¡T�9��l���� M��|c�z* ��	�J�ħ��Pb�D����|��ܓ�{���Asu��71�94>��<���� k}x��0<��DEV��x�p�t���LҴTU՘���(�������`YY���K�����:5cc!��Ju&�d:�F��]������GO�w{���ں�>Rk����n0�n��l�IB^P�>�{׀w�}'�Z��˔\���� �[�興Jd�� ��x��3�yDB�C�4L�׋���J����;��, �[�:$�S<������>�wR:������j��`t%
"g_u�����޷%?|Ob+ �Sʺ`��"��Ą��!*����>|��ʦn��&�j� {Z� ����ޯ����`�rI����$�Z�f�a��ޫjN9э;q$��,�ݝ6�+�s]���ͩ������{I�K;ėz�����m|`-^���ߖ�~���S1�bnM�n,���x:}8��y�=T9����6�I��������^}V�{���n���W\�aI�ƔrhrS��N k���,I)�}׀u\�����J9�{���3�	%��|� }�^ �����B��ӽ��zw���}�����M�   �!� K����]B(�e(۶�m�͓��8	������1�W)�P��d���5�y9R��9��[�0�Ɯz:��i����m�][A���q&�y�ݰ�Nkk��:�N#YY����m.���m4���`m`muT4h��c7�2jv�v��݊ˢ�O��+�v{<��>�=���]e�������ލ�~ {�>|������:Ķmq˳�uJ�O!'/=��d�*�69�\�}��{I�m�Ě���u����z٠~{l脔B� k��鹞�������&�j� }��r���d����� �z�o��bG��o�iF��D��rO> �`�`�`�}��kb �`(X � ����b �`�`�`�}��kb �`�`�`�ﺿfg�f��ˆ�k56 �66 �7���� �666=��p؃� � � � �{��؃� � ؈� ��w�؃� � � � ��}%�3X�d�j3Z؃� � � � ����b �`�`�b�� ߿~�� �`�`�`����lA�lllo���lA�l�g{��w������o�R�s��un�n�P�-gI�t��C��ȉc�gV-������fI-�D�Yu�6 �6667���� �666>}��6 �6667������666=��p؃� � � � ������u5L�Z&�Y�lA�lll|���lA�G�S��6h����A�A�����A����{��<������}��<��僐A� � ��Y��d�f��5e�ֵ6 �6667�~���<����}��6 �6667���� �666>}��6 �666?w��,˗>�k���f���A�A�Q�A����A����߾��A���ϻ���A��,}��p؃� � � � ����߲Mj�Y���.e�y�~�[y A�����A�A�A�A��}�b �`�`�`��{��<�������w�~������+�Ɂ�D�mq�ۈ
��Xvu���n9X�3�����{���������֤��5nkZ؃�lll}���M�<�������y�߸mU�A�A�A�A��ﵱ�A�A�A�A�������h�a��hֳS��A�A�A�A�߿p؃�"`�`�`��{��<������}��<�����wM�<�X � � ��}%�3X�d��sY���A�A�A�A����A����߾��A��<�F�AP*@���D<�A� ��7�؃� � � � ����b �`�`�`�{�t�fd��4L�]f��<����X �;��؃� � � � ��w�؃� � � � �����A�A�[�߸lA�lll}���ˢ�j�f�L3.�Z؃� � � � ��w�؃� � � �"��{���A������y�~�[y����??�ڪ���t]<���e���à*AD�=��53Ƭ�6��F���{�Q����uV\�䚫�2B�A�_���X�[�����!�;� ��!53U]uuL��ݘ��zP�	B��z��_���frI)��鹞�������SU5k >}׀~{lÔ%3���ۚ���ڍ��r'$��<�^�w�[�0�^,В���PBKR�Q��ռ>k�>�$�r�3>�4f����s��`l��s�_}π6�Ɂ�����w���������wf����ӫ4KE��N뭌�sp)u��jئ��w��c���FR�����s@?u�@�zS����:���s瑶O&5� ���z#�%F��� ��Ӏo��7��<Ď��_j��s��rh�o��s��B^��UϽ� 7���=狲�5�XD&䆇�b�/�@�� ~���P�o����됚���]]E5sWs�o��`�����s�4y�Z���u&�I$�I    աS�ч��}қY҆�<Xp^.�Ƶ"���{rh�tl熂8�qWt�/;vd�s��eݝE����)�h�TՒ3��v^\@m���7h㙌U���;L���w<��۲��k?L�tpg��&�v���q[�q�Y�L�b��W���Y��mZks����h��ٶ��ܽD�a��酌;��]3�U^,q8Y�oe��G�X��٥7;iҬ�4�����S�[�����_o���i���i��o���?^��=��}���~Az���u���R4��I����?����}]��9��`�n�%
&O�z���VR.iZ��0t�p�^,9(�2|�� ���k��sWQ7AD݅M��y(IyD*���`��x��P�]�� lMu"�y0q��h�hg�]��W~Z{�s@�λ$�`�<�Lo$&2a�q��t`�n��g]^9��]Fkc2����\_�����"I?��|h����������uyY�Q�DܒnI����H�����j�+��S�Y��n, }�x����ď��i6��?������� �jg�3}W�����t��/A,I���m9��u��{����Zx�_�f����R4��I�4ו�{��_>0.Kz���RI%�gs!T䵱瓒&]�Hݝ��N$�޽]:8���tv�F�W����m=q6�m��t���X�n�!~����oW"zj�&mM�T���kŞP�B�U�޼}�� {M�tDL�bk�UA3J�wEլ ��x��'RP�C�)E��B����~��r���ۚ�q]S�����&��b��"~�`�p�^,Q�"g��M��ϔmƒ &䆁yڴQ
C�ߗ�}׀~{l�ԷvM$i�$"YZ���[�����k����<'1��v]������}��D~��L��U���ŀ[���g(P�~����Z�|�_0�H�MA6�� ��y脽�*�}�� �zp�^,�^${nD��8ԍ'!�M߬��;i���P����`��x���S�-UҒ�]�5fB���� z� ~�w�)꿔`�� ��H!T#�"�KХ���?W��5wښ&칺� ߵ��=��%[����_��즀{�ݒI �!��GoȢpW*����=�F��V&�RlzZF?{�}|v��+�L$ds? {o�@�zS@��)��~Az���}�/��)(�'�rM��frQ2|��=}� ?n��Jd�X�|��nܐ�=�|h�]�>�"��h�gƁ��$�۱��uuv`z!B�Es�|�{�x��D(���V�~�y����L�����Ԣnj� ~�w�z<���x����l�$�R$�`�FS�@����æĚ]+"!	�\�I$ Hʦ)�`����b@�
JD`0��*`iMRt�z�c�!Fj��x���R2�.�IUȑ�A�n��GI!��1N�= qB�< �p �3#5�����bz��0"B1$�v��ā���`C	�8r�<��$4�H����S�, L	HL�<2��9�5t.�IHk�h�	��2;D��z�o��c���j�                                 ]Ӕ�f�h^�'G�v�嫌j���Z�� %1�[���=����f��V5�C��y��J���s�.U��\/9���#4��-��蝬VZ�A��1�����b��(�̈́��&���:�v�K��,)s�y�F�B.��(���Wn亶�u��x,h��_m��1�v{�rJ��f�x�Z nA� ���ҵuV�w>J�[`ͷQ�v%��p���Ҽ��FyU�ȵ�눸�m���bZ��ck��-�<4���:�uϐ��=m�l��s�??|[�N0�=L�rx�<�T�N;��l�H��F�8)��!-M¼��]5+���u�e8�Hm�ZUەg>ě��+���B�U��8+���%ۭv��K�n�v��er��8h1��4'Ó�K�3��@��z�f�Sv��mA�h�V�6T�6�M��g��*�+J�mژ�sd�#a&��P�e�*��(�\ֶ�̌�-k�8��\�n�2��yֳݳ��MQ��쥖ɘ�b��w�uXB����rUC]�V�g���9�<�S�IS�����݋��q�m0[�-*�9mh�v�)Pvs�JKUt�kF�em�N�[1�g��)l(��t�S°�93�0U��;t��۵��R�8RY�'<���{\��'O�%m��xܦ�'�B�&V�.Ԇ�q���]H[�K����j�n�� %Tj�복(����*�lj�`Й܆5�ض��s[��V�%z �az�+��/Q�+Ȼ��&(��P�W/l��
�*B�#��,��2��SV�(�˧��)��`ɶ���c���Y�� ��}��7�<���Rˑ۱Eϐur���������ԧ8G��V�U�]S9i+�s.�>��
� �T�k�яQ��|*+�	�D<EJ�=z(�C�������      ,J���Yz��z����m4qֻk�RP��Y �fR)�+gY:��܎���m�g�At�.�U�띖y �v���v�:9�ghݦ�OQا<s[cv����V㜫��S��.\k��9g�'A�w�m��r�����\��(�m�*p�0&�UEԛ�ݝ+�v����V�xm!V^�Eac^�{�{�����w��U�KM���n�( #]�N���x0�V닇��n�����̔�Z
��9��`�m���BQ�@�����ꮨ-UҒ�]�5f�vٟ�	Dz�Ts�b������3�(�:y��x)��AƜ4��� ��f�fy�{���ύ ��xF�$�a#W{3m�`o����EF�/�� ��}�H1G1<C�h�Jh��e|`ISgrT�Iq�g{��Dql�W8Z�ؘ�븹N#,�.^��ˣ���2(8ۃA7$4�Қ{�V ~�w�	DG���w\�T�nj�Z��s5��ܓ�=��݇QN�*��F�ک\�
Z��>��x�0۶��%Ty����$��M`�s4���h�Ji�%��@�~��/vD�1Ƥi9��hr�?s�0��0�^,B�%U�޽�_ͯ�&91�B'�t�����_}π6�&�*0>�{RI$�i\�.`-�����u.�09����y��b��0q}�n�SZ`�&)p��ذ����g�Q�C�� m�<��y0������o�${���ύ�빠�V)�b�bx�ֵ�';�7$��s҂/ � "%QU?kŀ6� �iN�*��M���]ف�S�y� ��, ��������@>�菛ȢqH�	7�����g�U��/�T`}��c�j֪����^�+�UlX.y�L���ưZ��2���â�$�Bq%կ�7׀~t���m�	(� ��s�?��"�drFӐ�I&����<�DL�7|`�ŀ�]�DD)��i/��c�$#qh�>4|���O���>���h���"mMd�MY��QСEww�X�޼�����C��#W�] ��O�'��߿� ���#l�L$q9������%��z~]{Ӏn�ŀ?�>���b���r�!��IN��[kI���9�+Y'.�������x��n%]��>��������tB� n���ϖFF�1dۑh�v���D/(UGw{ 7޼��:!)���7�D��m7�m�s@����D�K�XdL������Kİ}Ͼ�Mı,K�N��ܷY�4]\��Y�iȖ%� )"g{��q,K���}��r%�bX>g{t��bX �2'{߼6��bX�������"RHy�y���#��e�S�,K����Dhw�]'�,K���p�r%�bX��s����%�bCh��1"�t��sV�k5�kZ     s�i+FٽǇ)c^s�ֺ㮱�IT�V@R��'�v0�@���C<[]qՏN���9Ӧ
�Oi�c�F��� ������"K����Z������ɓ���l��c���U\K��Gm�n8���h� #�zX�zc��@ޙ�lܵ�뵫��u���cls��m����>�>�ۖ��::�.�o��{�{�}�wz>~o�9'�]M�� ���m��i��s��m�cc�Sؐlc��:�Z�����)��5�Y�5�Y��'�,K��>�t��bX�'���ND�,K��wT?��Po�5ı=��߮ӑ,K��g�\�B]&�.K�]&�X�%����ӑ,Kľ���Mı,K��{v��bX����&�|(�TȖ%�{I�Y�L�h��j捧"X�%�{��U7ı,Nw]��r%��C"dsﮓq,K��{��"X�%�g�/ut�jd��35���bY� @Ȟ}���ND�,K����Kı=����r%�`|�L���}���bX�'{����ɬ�Mԗ35���Kİ|���7ı,?�
��߽6�ı,K��~�Mı,K��{v��bX�����*���4�����C�*a��.li��]�����S�u�͎�?�w{�F�z#5uu,�335t�D�,K���iȖ%�b_}�q,K��u�݇��"dK��>��7ı,O��]�~�Y�Z�W),�h�r%�bX��s���q^"�� @a��ȞD�<޾��9ı,�~�Mı,K�}��"&�5������2k5�f\֦��kU7ı,Ok���Kİ|���7��Dȝ�~��Kı/{�j��X�%����2��3553,�Mfj�9ĳ�~��=���I��%�b}�߸m9ı,K��T�K��}u�o�ӑ,K��ωr���5�r]j�7ı,O}��6��bX�%���n%�bX��۴�Kİ|���7ı,O}�~� ꗫ��3�i,ӥ�sti��k�-�Iv㶝�0e�mJ��r\v�%�#�M\�h�r%�bX��s����%�bs��nӑ,K��;۠�r&D�,N��p�r%�bX�{�~��f�,��35���bX�';���9��+���`�?~�Mı,K���iȖ%�b_}���|9S"X����k5s50�����]�"X�%��}��n%�bX���xm9�(�K@У��,��D�K��ک��%�b{�-�?b<�y��-���E��0M�f��q,K>��;����Kı/{�j��X�%��뽻ND�,��F�t�,!I
HRB�:rfzK�.ɻ��k4m9ı,K��T�Kİ������<�bX����I��%�b{���Kı?0��>ֵ�����mQ.��v��َ�L�7g-;��g%��B㛑�䫡��̣Z	����bX�'�k�ӑ,K��;ۤ�Kı=����~	�L�bX��ϵ^�{��7����ߟ�w�me4�c��bX����&����,N��p�r%�bX��ϵSq,K��u�ݧ"~O�kQ,O�~%˗�%�rf���WI��%�b}�߸m9ı,K��T�K�a�2'�k�ӑ,K��>��7ı,Kﾔ���2I�W5�6��bY�"g{�j��X�%������Kİ|���7ı4X�S}U>A2&w�zm9ı,K;�~��f�,��Y����Mı,K��{v��bX����&�X�%����ӑ,Kľ���Mı,K��~�Zֵ�h�2h̤�W1�`V\=]g�����5���՚�77f�S)������|t��㭅h�=��Kİ{��]&�X�%����ӑ,Kľ�������,Kϵ��}��oq���������%�
fj�7ı,O}��6��� G"dK����n%�bX�Ͼ�[ND�,K��n�q?��&�X��?]�Y�ɚ.�RY�Ѵ�Kı/�g�T�Kı/;��iȖ?(�ș����Kı;���iȖ%�`��㹙�kA4{���{������ș��}��"X�%��}��n%�bX���xm9ı,K��T�Kħ���ZYI���4��|�ǘ�1b��w�I��%�a���xm<�bX�%�s�T�Kı/;��iȖ%�bh��bAvw�w&�      	�N:;)�d���sj���k{k��\oOF�I��FX���ۦ�n�5��RiC��-���^)k#��8#.M�ѯa��gns-�c�G-�ݰ{v�As��9y�n��d���tT���k��G��V8�҅�̙ؖ��]u�����l��$�Wv�6:��A����Y��3�W�n����O�w{���_πG-��n��g�6�lI���GN��6CV��I]m�a�����؄�v##p����q���ǝ���ӑ,Kľ���Mı,K���&D�,sﮓq,KĽ�JO��̒e�D��f��"X�%�}�;����șľ}���*dK��~�t��bX�'{߸m9��Os�������/�M��Z=�D�,K���kiȖ%�`����n%��dL����ND�,K����n%�bX����v��\�e�ԖfkZ�r%�g���>�ﮓq,K��{��"X�%�}�;���bX��
]D׿�~�ӑ,K������ɫ���SYm̹��Mı,K�}��"X�%��	�s�T�Kı/�}����bX����&�X�%����<�j�w7k��u���9�8����v)�(K��^�Z5ź��\�Bv4ݴ�Kı/��uSq,Kļ�{��"X�%��w�A�)9"X�#}�d/�)!I
E�꺅7WWU5v\�f�Sq,Kľw��Ӑ�Z����A�4 ��$X��#�a�y����D�K����n%�bX�}��ӑ,Kľ���M����w����ߟ�w�me4������,K����Kı=����r%���MD�K���U7ı,K�߿kiȖ%�btΓ2�v�L�����n%�bX����m9ı,K��T�Kı/��u��K��du��I��%�b^��'�]\$ˆ���56��bX�%���n%�bX|�s߾�[O"X�%��}��n%�HRB�x̅��$)!I
S5����*K�\�j��ntkFN�R��Rhi�q�Vzֹ�3i�q���}�Eⳉ�x�G����%�b_~��m9ı,3��Mı,K�{�͇��șı/{�j����1b<��+>YMƅ�ܓS�,K��;ۤ�Kı=����r%�bX��s����%�b_;��iȟ���Q,O߿n�\����e5��˙���Kı>���M�"X�%�}�;���c �;B��tŻ(��D�P箅"���#�P4���'~	���k}
#Ȥ 0��xE\F�z��!�`a G�聂���u@	4#�&�! 0 Am�I�1H c�4#W��,q	$Z	4�X�Mz�Si�q@<�A�n�6������h�h9*�BL@t�Rp��U���')P0�EXZ(�A6��<QC�ꢴ�"ޝE�y�
z�1T�EBB)�JmQ�Z���Q�^ �(xyQ.���r%�bX=��t��bX�'|����MfL�ur�˚�ND�,�D��>�Mı,K���kiȖ%�`����n%�bX����m9ı����9�̣Z	�����oq���[ND�,K�����9ı,N���6��bX�%���n%�g��w�������Uӳ�6���%)(Z��K��(����bq��5��{F�F��u!�M���-�[�ּObX�%�����7ı,O}��6��bX�%���~��&�X�%��ߵ��Kı?g�\�3�-�2拒�WI��%�b{�wٴ�Kı/��uSq,K��;��ӑ,K��;ۤ�O���,K����e�Kp�5r�ӑ,KĽ�}���bX�'���6��c���Q5����n%�bX�}��ӑ,K7�����x��n2���{��7�"{���6��bX����I��%�b{�wٴ�K�8#2&{�wU7<�y���^�YVGq�Cӑ��%�bX>g{t��bX�G���M��,KĽ�}���bX�'���6��bX�'�G���z��ѩ�V�fMjf�v�<ݧO<�;=J�y[mb9+u��A�.ˣ���}��z!������oq��������ӑ,Kľ���Mı,K��{��y"X�%������bX�'�Ϯ��5�����e�M�"X�%�}�;���bX�'���6��bX�%�w��n%�bX����m9�*dx���ޗ��L�5��=�oq���X���}�ND�,K�;�i7��dL�����ӑ,KĽ�}���bY�#����S&7&�b�=�?b<�~?-D�����n%�bX�}��ӑ,Kľ���Mı,K��{�ND7���{���?��+I^ﷸ�bX����m9ı,>V9��کȖ%�b}�}��r%�bX�y��I�{��Y���=�}���cI�      ��i*^�S�v�c1�{X=��utw�8��>�8���98e(���0����x]H8�lpс^S����cÓ(���]�]oX1Nv_Yګu����\�.j�^��6J1��`mq�6�2�y��]D��J"���N�$[&t	݂B��ݒ@��f�n�[�
tqƸlvr�Qz8�KU�7,#8��ݺ�o�$���vE.��ۊ�/L��a��jы�
�3u&ǩnX���w}���x�e�D�˚�O"X�%�~��n%�bX��]��r%�bX�y��I��%�bw��iȖ%�bY�K�]kRˬ�p�3Z���%�bw�w�i�| șĳ߾֓q,K���o��Kı/��uSq>A��,N����5��f��P�s5���Kı,�ﵤ�Kı;�wٴ�K���������n%�bX�����o7���{������C�g��+W�ı,K��}�ND�,K��wU7ı,N����9İ>fD�{��a
HRB����8.�ժ���l����Kı/��uSq,K��X�����yı,K=��i7Ĳ���fB�B����ͱ���ݩ&�:;Tq�cHa�Sմ+rR�����pq׫s!�.5�W���̣Z	�����o'}�{v��bX�%�w��n%�bX�����|,�&D�,K��ک��y���^�}���Iqo����%�g����Q��5gG|���r'bX���6��bX�%��~�Mı,K�뽻ND�,K�5r��-4e֦�R�ZMı,K��}�ND�,K��wU7��Dȟw_}v��bX��}�&�X�%�{�'p��I�W.jm9Ĳ���ߢj	 �w>��I�y︚�H�D��s��Kı,������jYu�.fkU7ı,N����9ı,=����bX�'}�xm9ı,K��T�Kı?����UWI�U��e�x��
��]��I�'�	��\k�"kS�����釙1n����=�bX�~��&�X�%��{�ND�,K��wT>���,K���ӑ,K�����j�段���f�ZMı,K���6��bX�%���n%�bX��]��r%�bX>{��7�*dK����>5����e�Y�iȖ%�b_{�j��X�%��5�ݧ"X�� �!��S�B]+� �o�X��g�}�&�X�%���}�iȖ%��{�?:_�BjQ�q-ﷸ��%��5�ݧ"X�%�g��ZMı,K���ND�,�D�{�j��X�!I	��]b�Wj�Ww5W9�
H,K�=�bX�~�~��yı,K�s�T�Kı;�۴�x��{��??ʪ�ٸ��&�#�nz�%5r��@A���6�ym�Ź�ي��BY�.�5���kZMı,K���ND�,K��wU7ı,N����>�DȖ%�g��ZMı,K�ޔ�aup�.&�k4m9ı,K��T�>#�2%������Kı,��kI��%�bw�{�iȖ%�bY�x���X��<#G���7���{�?˽�ND�,K�=�c��"dO�߸m9ı,K�s�T�Kı�靖dq<px��Mȷ��y���2{ߵ��Kı>�~��Kı/��uSq,KHQ�x��L���iȖ%�by���0���]RI����Mı,K���ND�,K��ϵS�,K���}��r%�b�Q��WRB���3pwwwwjKB�͚,�YצX��Ҧ��u�۫3�����rQ��Z����ﶞ�������{��,K�s�T�Kı;�۴�Kİ|��4�șı>�~����oq�߿��)=R��R���%�bX��]��r	�����~��I��%�b~���6��bX�%����	z.�Y
H]ݞ�����VJ�����r%�bX=���&�X�%��}��"X�%�|�;���bX�'}���?b<�y��9Ѵ�0DƤ#r�h�n%�g��D��߽6��bX�%���U7ı,N����9�@��.�G�~��s�2&eL������x��G��������)�w�Os�{��Nr�D̩���}u��&eL��G߾��*dLʙ��xkiș�2&eOG�F@B;|�Hf�qB{ӯޫ��}      b]v��&v��\t�%�1;H��$�)#v�J��b݆	L�{�:wգ ���F����n7l���ur)ظ����V=���#r���Շ5�V�F@wK3Q�l�95ؕε����[=�V1�\8���]�ʗeo[V��K��t�YXy�7O��^�%�5�b6}�4A�\�v��7���8X��;��������w���ꪺM	s\7Q; !��RU
�m�Sq�y5u�� ��I˩����w���>��A��<#G���=��)�w��߿��92�Ḍ�{�I�Tș�2%����ӑ3*dLʙ��T�*dLʙ��Ӛ5��f�Ԗ�kW[ND̩�3(����s��#�k���L�~��m92�D̩�}��S���3*dK�ۭ�"|(��&�fT��Nj����]RI���֍'9S"fTȗ�������S"fT�}��9S"fTȗ�w�[ND̩�3(����s�2&eL��{wr.�f���e�Y�[ND̩����T�{�j�9S"fTȗ�}��ӑ3*dL�>w�4��L��C��&��������S"fT�񻟌ˬ5�f\ц���T�*dLʙ����iș�2&e;�Nr�D̩�/�������S"fT�}��9S"fTȗ;�wZֵ�IĮ�cI�Kw���8�FZܚw]�:���D���7f��t����r}��Z�ũ]]q<��S"fQ��i9ʙ2�D����r&eL��S=�;����ڛ��S"^��뭧"fTș�>��s?BY�.�5��sF����3*dK�᭧!�В,$<T�Qu�+�S"fT�w��Nr�D̩�/���[ND̩�3(����s�>]T֪dL?8���.��C7_{��ܧ��婝�}���L��S"_5��m92��Hj&�G߾��*dLʙ��p���or��{��;����.5p�����L��$D�w��[ND̩�3(���4��L��S"_}�m92�@����M��~�Nr�D̩�?~���f�������j�iș�2&e;�Nr�D̩�/�������S"fT�}��9S"fTȗ�w�[ND̩�3/����} �̝��ae�����sm:	���d��x��JrN�\���籙z%�v���ִi9ʙ2�D����r&eL��S=�;���L��S"_5��m92�Ḍ�{�I�Tș�2'}��!��gN�n��7�Os��{���*��L��S"_5��m92�Ḍ�{�I�Tș�2%����ӑ3*dL��������OT�sԴ{�����r�2%�]��ӑ3*dL�>w�4��L���R�@��b��v�QZ��~��5��Lʙ2�}�wU9ʙ2�Dﻷy��њѩf������r&eL��G�������3*dK�᭧"fTș�3�s���Tș�>����﮶���S"fT�r���-���7^����;ܧ����᭧"fTș�3�s���Tș�2%�]��ӑ3*dL�>w�4��L�������??�Un�u�`w���գLc=�n�o-�1��6�XM�it�p�5sY�[ND̩�3*g��uS���3*dK�ۭ�"fTș�|�xi9ʙ2�D����r&eL��S'��~EⓉ��F�w��{��S��q�ۭ�"fTș�;=�Nr�D̩�/�������S"fT����Nr�Ư��s�߿�w��釙1�E*o����2�D̩���19ʙ2�D���5��L��D֪g�ϵS���3*dJ��9�g��my��^gZ~��Q�E�-ֵ����3*dK�{�[ND̩�3*g}��9S"fTȗ;�s[ND̩�<WM�i���
#7jvs|19ʙ2�D�{7y$ְ�jd�K-���r&eL��S;�wU9ʙ2�C�U�k����y2�D̩���19ʙ2�D���5��Lʙ2�_���g��,���Ĝꭳ2�.㜴�1�Fs&�	8��z���I��z�Z��Tș�2%����ӑ3*dLʝ���'9S"fTȗ�������S"fT����Nr�D̩�;���e;4fjjY��\�f����S"fT���19�|?����L�~��m92�D̩���ک�Tș�2%�;��ӑ?��b[ܧ����/��FJ��7>����93*dK���[ND̩�3*g}��9S#���SQ.{�٭�"fTș�>���'9S"fTș��S�	��&\4M\�h�ӑ3*dLʙ�s���Tș�2%�;��ӑ3*dLʝ���'9S"fP�Rj&w�xkiș�2&eL�|_ؼRq7���s��{���󹭧"fTș�;=�Nr�D̩�/�������S"fT����Nr�D̩�1uHT�0M�) f��N��ѭ. @b�A��B�@���S��`F��UqN<5�w��s{L0 ��Bl��[�c�}yW��vt�h�0!"x�
D i�N	
���^O|�"sH9�0<�a������C/2�!&.!��s��k33Zր8�l�j�                                 T�6��Ҁ��kW�7bvqkg��J�h8�l�z2<8�n�!�q�zA�,��aq���6ݱ�v4j������z,�Xƪ�1�.��^e�ᬀ�ul\���	��Nsr�;b�*���=]��I��`ܷk9�IΗ$-:�&��\ܰ-���SbN�<l���@{7Zq�t7�X�-�]͢�Y�F�yemS�u�U��:&���2��U����n^8�yU��ݷ���n\����$�t�s]��D�^;K����B;5�+�݇ACLO/:��� �5��k�����]Wv�	8p��VTr��+�[![U/6n��W��!�V�mJ�Yl�ĩ]N���̥�����=/;V�j�ín�&�Q����m�Jځ�*�0PM��nԶ3�&�.5������ �B�BX0K� T��vm2��+ʭ[Uu�ػ,��J��q��v�1̱�9V������a%`�\�9�qTqK��k�n��dc$��]�Jj��$����u���V�q��d�Q3�L[M��g-k�5�p�C���ۓ8���&yvz�i��������a�!8NݭmQ�������Ҭ�QtTZ*���0��[6Z�U��B��d�I%W1�6��d唧��#`2A)�{N�YB�j7�j��U;[��1!bI�jt���ǖ��5<�,����f�! R�ݵ@Y{k�(�<�����˴㭘zp���)6�kj�n�'lӜ�R��4��i��gG6 Wm��l�Yp���.l��K`�nr
,�
�2e������Oc>��T�n�jZ͡�����+�]�5�K��((��꒰��,�I(I�����.'B�[���*�����G���+T囂���W��r�M��*% C�׊�A�'U��O ��S��T��$�`�E���W���w?w�`     j���	.�rt��h���;�i���6Kqss!�\��1��i�z�tW )T.�WW�7�{�7nJ�OD��e���h��U�(2�&rnZs���cU��u����yJ��sѵ�!R) $����.c�Q4
��NI�^˻[���	WbS���ŌWo�F�Y��2ɓ4kN���D�L��Wo�����~ u�:����t�gt]������]�i��9�5e�r�0qN�?����_S2c��o����=��)��߿����*dLʙ��xkiș�2&eL��P�(��T/���Lʙ�~�}��or��{��~���K�-���V�bs�2&eL�}��5��Lʙ2�w��s�2&eL�s��5��Lʙ2�g���T��Wx��L����w���j]X����w�{��;ܧ�����S���3*dK�w���"fTș�;=�Nr�D̩�/�������S7�Ow������O4�ץh�?������)Q3^��kiș�2&eO�~��Tș�2%���[ND�,�fHUκ���$)!ss9U+�UVY%�j�k[ND�,K�����Kİ���}���yı,K�s�T�Kı/<�u��Kİ|��Zֵ��Kk��=Kl�s�ç�ri�M�g�u�ls���n��8m�n�����*���-/Cs��o%�b_}���r%�bX���uSq,Kļ����)<��,K�߶bn%�bX�gzS��d�.&�k5��"X�%�{�wU7b�`"�"��DȖ%��}��"X�%���혛�bX�%��{��"X�{��7���x��n�����D�/<�u��Kı;=��Mı��Dȗ�{����bX�%����n%�b<�y��_�8�#b�Q�$�3��(�~RD�w���bX�%�����"X�%�{�wU7İ?ș�}}��oq���������#��U�q,Kľy�u��Kİ��}��U9ı,K�}��"X�%��^*��)!I
HRӝ�wwwj�F��'[��#�M�,��i#�N��D=���Ѯ-��h�ZmK`�_{���oq���^���Mı,K���[ND�,K��������Q,K��~�ӑ,K���~��?�Ry�.�+G���7��b^y��i�~c�2%����17ı,K��[ND�,K���n%�#�G�{���Rc� ��Mɾg��G��`����n%�bX��=�c� ��UI"^���Mı,K��{��"X�%��t����k-ֲ�k5��4��bX�%��{��"X�%�{�wU7ı,K�;�m9İ>Y�~��4��bX�'�ޔ��5�$ˆ����kiȖ%�b^���Mı,K���[ND�,K��f�q,Kľy�u��Kı)��u�kZ�dת�m��幌6E�GUhk:9!�]|p&NGb��.\Qx��n����X�%�y�{��"X�%��{�I��%�b_<���r%�bX���uSq,�Y�����}�4nŗ��p�����İ{�vi7��DȖ%�����"X�%�~�}���bX�%������ߩ�w�����ߍ/D1�kF�q,Kľ�ߵ��Kı/}���X��C"dK�}��"X�$�9�+��)!I
H_n�,.n�����e�Y�m9ĳ� dL����n%�bX��~�[ND�,K��f�q,K���F(�"��
�5�"�Q�z�F�tD|C�E�""ȗ��5��Kı=���r�)u�Z=�oq����?���m9ı,�ݚMı,K����ӑ,KĽ�;���bX�'������'KȒ�t��VS�=vmkM�� 18Ѩn3�5�2"�ֹ����ֶ��bX�}��&�X�%��y�siȖ%�b^���Mı,K�������{��7��9U�ݧ��n%�bX���6���,r&D�/�ϵSq,Kľ}ߵ��Kİ{�vi7ı,N�});���L����k6��bX�%��T�Kı/;�u��Kİ{�vi7ı,Os�{�ND�,K�����u�)u�.\��T�Kτ dL�����"X�%��~٤�Kı=�=�m9ı,K�s����%�bw��浓Xf�m���k.��m9ı,�ݚMı,K��^���yı,K�s�T�Kı/;�u��Kı8�|FzK'��݀     �aS��u�r֭,�ekS5iљ^����Rܕ�*��5�ہ�{v���t�ov�A����.`�/]�F�m�]�NTt���c��Sf/n7�a��ݷ�;h������]�*K�����,lC\;�����ԮC�[��&�y��M�Oml٢ɽ�<��szWa���G;��f�K�4���՗0x ���T�9 �m���ȗt�Z7n�Dӥ������v�ֱ�H��&����\�֍'"X�%���ͧ"X�%��T�>���_Ae��K��a���u�M�0����W�6T��Gv?��ҏ����ۓ@=���=�w4�x��W ;�f�ލ%�6<f'��z��l|`l��M�0�T���m�a�JȜ� ��Y��@?{�h޻���vF� �tM���J/L墹��5��Z4�stm���b��Ra�8���٠��4o]� ��Y��V)��$M=krI�=�D<@L���������� 7��9(�2w5�wEҫ����,]��&��� �eLm��}���DV�(�QdI6�s4>Ľ��`{ɀ}���_H,��u	w�a�.��&ژ�*`m��~���>���O��I1	��E�qF���2�m"�qv����ɀ/]A�x�h8[������ۓ��~�����{��{l�/r����� ��NI�w7�:!L����{�����9BS#���?	���FH�h�~��i�A�SbX�b��&�H�p8v�����ذ?j�:SsH*jЯ:�� �j`l��%���0��b�)1�RA4ӓ@?{�h���*`mLfV�I..�8fb[vn�s�Y�������.��t)m��4�-�GQ�2I9ܙi�4�w4�ʘ�S �eL	b���X��qfgzuuq���q�m�0����+��$Z5�|��"qLHX��@/}��{��=�w4�ޯ@��u�iG�F�q~]�R`l���W�ٲ����(I�Jb!!D���vn��2�VISw5wx�^,��k�� �����f���$�c�%�Q�ۛ]��FZ�wC  �e{��=u�:�f�%�i���G"s4�ޯ@;�f�w�g���w�����<Dx���#qǠmLl���W���?~�{��%<RcX��i�&�^�M��s@?^�@;�f�oe�$rcM����(��~�|�{�x�7x�Q3�M�b>o"��D�n'3@?wY�z^�_����>z�`��(H^�׽��|��[p   �  %�
�I�ȵ�nza9��ipk롞x�cZ���u��4��6���{'^���7k۩J�'j�Ł���Ů����8�؁��ݣ.n�NZi!s�n�۶��6X�W(�8�q�Ny�����\����@�W��%��jQͥe���k(=Z�N���<]��x�uh�$X%s]�����}���w{�o{�4��?���TLGX�:��\M7b4��ޱ$��v�wN�4�JÌ��=P�ن`���Y*`ISl�������;���Ɣx�m̞Fܚ�����DD��݋ �y�`�w�IL����W�:��ı$���� �J��� ��f�����0r4�ؤ������ ?n���J{{�,�yJ>x�x9�E�@/u��h�w4�٠~�[�$�dh���LN��eW)u�J*7[f���lus��ִN]OO�x��<RcX��8��~ ��h�w4�٠����#"y ۓ"������,�_�$�IA��Va"� � ���p]�o�.���[�O��M ��4�[ȢqE�$����� =�xr��M���;{�`�Pu��D�bBQ�4�Y��f �oD)��� mS�U3t��f��uUw�6� �v�~_�� {��I?��������rN-u�7^���;H�:s)6�ӗ���n��E�l��3_�w���W���"�I'�_��� �h��J~�>������Wu4]Q6��7eO���`z�&��L��0"���4�NM ��h�m������ f:��*@�S4\T��� ��  \��]�x�7�&��-W��f��b�9�1��ݚlF"ɣi) �Ç�8@	"E�q0�"DB$P��dI|qKDB1]��о�4H5�p Hā&ͯ����04���6�M��pS��G�tQ�#�Q�l:*o�@h�4���������f, �ۼ �ܻ���*����\�]��B��B��w� ���`{�h�@�{.�ȞH4�ȣ�Ԙm|`eL�S �ʘ��>�{�������X[}�MڲNm����[C�nHI�k�6��r�̽�t�u.|e�`J��U����|`^��I�7HJ9&�^�7�bA�>��� o�� �U��L�*�������&�ژ���7eL�S��m�9E ���w4�=�$�����Xx�mD�A)@,�T�(���5��7�D�f�긹��&F�JL��S �T�>����0=��� G-GV;v�km��t��t�N���[����qlQ����+��{K�F��� ��� �mL��0�S �ܱO#��)"N(���f�}�s@=����f��y�G�\�dq'���2.�w�0==���*`J��j`u�V�(�QdI1�ɚ�f�^�x����DB���� �)����Wcq����h�@?{l�/��h�=�$�/�x	O�!8�L3(f"f���5�ֵ�h     8�nd�d��t�f���N�N����=�ob����{+�v�`�/&닳�˵�-'q�9���9�f催F��z���lm�����K���6����b�:,kG;@�������-c�����-���ٺ��K�w%β!��zCqt9+qk�j������<n�>�9�M��X�.͓��������w���UU�d�9��ev�m`��1��j'9�b�ն6<�vճŹ��J<m&ərh[f�}�s@=��������h؛�# Ȥ��v���*`J�6^�&^en�	���F�&h��h�O��J&\���;{�`N�J)�EMU�S75w�С%<�^ �_V �o ~�f�~�X���mD�Q�4^�l~���==����0%LتI*��*[]]F�]�%;L��Ʈt�+��� �Ӝ�c��99���dk����, ��� =�}��:�������N(�$���� �z;y�y�E"0��(�Z AU�DMbUJ- �_JjN9f�~�@�۹�~��'Sc�n5�f.�����ژm|`���;�%�n#�ۓC��/{女��>0�S �T��,�{Nw�]�bF$�m|`{�9̒�|�|��m���d�BA�drc��&ns����'Du1unz��n.��X���w
ω���F�&h���{����?�!~���ŀ9�R�Er���ԩ���`J��j`]��nʟ�s�`o�/��G1�G"�I���M�n�JR��!D�>�]��w�~z�]����q�4>�1}�}�4��4�Y���h����N(�$���� }���<�B�o����x�x�����$� 4D��(A&�0y�c�"���$v^^2kT=�0��h�����}���w3�ԗ���`m��d��}�4}ƺ�iA���L��4����No�`����w�n��U1Z��GE��`Y+� ݕ3ه������@�qV��ԉ27���������?(�IyL(�	�P�*?u���:_)D���UUjT�M]����=?ou���X��� �J:�������n{�!ڽ�ڝj�'3.6����n�WN�Z�rQNe��pٚ_ l���_��ϰOy07�>�&F92(�rh��h��� �n���y�Q���W����U3*j���s�^ n�X~ݼw}� ���'Sc�n4��rM ��4����]���M��cibO�\]�R`m��d��vT�.ڙ%6��2��vL�ֵ�     �S�������A�$:Vr�[	�u�;���9X^��[�O3�t>wi�N�0M��|��ǣv������Ivdr78:8v�ccSC��f�2�����ܘX�����u���C�n�f�4���ek]��4&���H�Vl��:܉�·��j�ng����L�؊Nu	��J�n����K�|�[v��'KȖ�n��XΚmM��[���/�V3�5�8���qtK�:,HĔvW��*`�f�~�٠r��u�)�BG��}���������g�(^UG���R+ʁUU�S55w�~����h޻�����9����vU���z#�Uk�� ��b���x}�4ײ쌍�#�q�4�]� ݕ0���ژ�ޜY�$�U��xշ7ZM��t��"�t��l�YѸg��c�"��)�C�mW6	/� �*`m��vW�����M�A�Ą��h���7ĳ3'� �mL�_쩁����qw���RX��ޤ�>�S�_�s0��0w�M��M�$dI$�/u���S �j`m��2�/{{���B�%՝\`��v��>�S�w4�<�/����I!�I�rbr`�n��X��s\N����Z�j�M���,U۵Ø�s$ӓ����@?^�@��s@;޳@:���Y�"8��@>�S�_쩀]�q��s��2<s"�#�ɠ^빠U�^����> ^�7PыǻEP��NZ��Y�_Gk�(�QdI1˛���=\���{� �x�x��}����S(���h�)�}��� ���������RS9�\B��[@�\]�7N .7%�y���r�sQt�lʘJ���e� ���v����U]�eݗwx�x��(Q2t����� o]�%29�=U�ڛ.lK�:���z���[��S�_�����s(�@/�ՠ��X(J�dBR鿫 ?1�~W1�G�R- ���/u��*�^�_U�@�ڞ�$�#�S'�n6^�.\���u�8땎Y�^cu��ts%,�"�9��i�&�{��U����ZoY�_Gk�(�n<i6�ĸ��e� ��� �T��W�z>��m�ą�8���Z^�ÔDB����ϫ ��[MT�ҫ���m]T��D)��׀s}� r��������I��Y$�BIe|`\���sfQ�[*`g'B*Y����h�@��@�y�b���Y		B�_
����\�Jټ(�S�]��|}v �:P"�Lc�}�x��`C� �Y��4$WHAe�E��JEc<|`yᾰbČ`��Z��oG+SD�9$x��0B���h���)�� @u���~~v��'~O��߆���i��                                 k��*p��C�<�*�u��fa��`���r&���)�6��p�f�4��W;����;n
N�'(f�����F��wbl�dN��1]����gf�JJ�l�z&L�<�<\L�x���V����۪q��.YW���R��u���N�L5r璹�����aG�@���6��"6�֧v:��H�����p�\6絻j��ݥ�^` ���hm��{vkK�Gky)_/���q]���\<ai�lѮ8 *�&�M��gw7 F.���'Z��Y�Q��\r�۲�ۑ�Aר���kl�vuf�狴涃uG��0�����N��QM��h���h����SvV�{S���.(l@/*t�K��{g�TU��g���h8�gf�	�3T�C��4�HR�U\�*b��ɴj향�h��zң�Ү�UU�IQJ�-*ǃnKv�����8eZ���	ڞaV�d�4�b�P7Fta�t�	<��Y�eL���u�.�qO:��p�zyN��:z0��T �\CM��:�)u�wl[�ڶ�8����6�u�OZ�q��8��R��l��n�Z3.�5���86�U5��I]�=�mG:bݜ�+/6�(sH:n4����t���l2u�pV��-��u�ii���t���q�ѝ�L��5V&�x��L@VW1�� �X���1�dP�:eU�B�\�L�g��n42�R���u�:�4aC]3::��'I��Ч��>K�z�Of�q��]js�O\�v�����̔��X�����(�R�Y��I5�d[jB5��',6��!�2�ܽx����t s��52s`�6���3`��Bq7^���Ԩ�2[]�3�ƌ�t�!ل�G�4����L6�c��������'QOP4�|�h���Oc�����:b>�������{}�;���u�����L      9�/�V�^���L1������ێq���b�9m���M�ֲ��F�O�����]��k�g�Ʊ�u����+�������6�a��9Bw9ov��.v^��a���]��9:5��:�ҦY�9�Kd!�&nuA���;���C�P)$��n.�����b9��;Sl�$�ŭ:��x]�J�����=��z�|�q:V����\h����NKa��{9c���9嶓�#3Wϲ��$ds4U��zuZoY�G�o�`-�W*UV�M���sKq�]�0,��rK�);��yC�l�h�٠^빧�y�
g����N��?7)���t���T�M�4�w4
���*��h�٠_Gk�(�iA�ۑI�]��D(K�N����x�x�Q�#h����z�3N�;-�zg4����%γ��˷�c]��zR��^Tn"��W~�{�S �T��%�w;�(��9"��Z}�o�����1\\�IB,c�����s�}󴛦&H̍A�4��hwW�U��h�٠r��u�F(E	�䗬�K��vW�Ɇq�6�,Q��W�U�}�f/������rK��{֒I..��C�#��t��mq.f�/4�i�&�ė�n��&�G��di��<�!�- ��4��X��]	B�!ӣ��>��.o#�2!��6��/�w4
���*���l�/��ƔN54�p�f�v��srN�'�����T������4�w4}k�u&�1E1!b�<�Sգ�������`w]`�>w�� �b�qh�f�}빠Uz��N�@�{[�I&@�Х��1�I�#�1շ���d�s.SM���Zi�"M��3$D�rM��s@��� ��\�D~�;�^ ��WT�l������ؑ�������_z�h�.�m�X��=�N� ��=��`-�`�ښ�V�yC�$Z}�h޻�]��8"x��(��G�3�no�'�|��ئG�dCymɠ_z�hwW�U��h�٠r��$�L�	M͑--�F�eZ��i�h��E��m<�r@;�����Ok�p̄2O ���������~�9��8 �n���k�X�KEt�*�Usjd�7WX��s�ȅ	L�ou���������1"�:�����9"��:��{�ɁvW��/X4��7LR(��BI4�]����~5��B��QU�w� ��Uz���"d��f�o]��N�@-�4�]��3ř�}�MbI�$�I$�I     ��D3$�#=�q9�u��8���Լ7v��-��*板��`~����m��F���r���g�\�qqW7M��q�`�qN�0��l]��J�Ƹ��d4JW�'M�[85��P�Ui����mn�=48;v�mm�l�������fHx�5������c����ۛ�[�G>0��Ƙ�f�豧�LL,b����S磌]��]Ԁ;�yy��j�]WO�Y���q`�+0���sv�vn{#V�M\խ���p����x��������Z~|�1�q$h�h�����`u���k��(��S'��>͊dx�D7��ܚ�~��/u�����q~Z�}��/��ƔN54�ޡ%���0.i.0������~��w�'��qLHY��U��`�����`u��<�6�ˮ����;��[���uؓ�8
�x��Y�k�]��J��7�^f�'��E��?�m�����Xz�r��
>�<�8��6��r(�#�I4�]�~<�0B�"�[���L����4��� ���9\U��#"�����7� ?�\��Q�G��x_��4]�q��qq9���.0���+��_�w;��q�#�pQ��_m���{������s@?z������I0M�Br%�$�ڻ!��7<�
�a�-���Y�Š��P�l��E2<s"��nM��w4�w4�����@��֢#q����Ը��W��ف�/��z{Ɂ�������ۘ�bBDrh�WU���[�����Q%h�6�fg�x�߷4��M�:�4�$��1qw�Ռ?��==���|��,�0�:�����1H�$Cbrh�빠J�ے� �j`n�ԒHH�],��ٶ�s�X�Asȗ��Ӻ�0��p��m�^��ٽTT9N�$�~� }�.0���+�d��^b�;�� ��&�~�u[�$��^빠r�� ��Z~.�ő�<�%"���`]��Y*`r\`[9x�..�C�ymɠ^빠�� ��V���0�<��q�4õƔn74��X���w-�v���W�I?��}�7T�htȗ�����.)�y(3c<�GMp����z�5l[���0+sN�#�@/�ՠ�f�{���g���4�u��%	"rE26�ZoY�^빠��}V��lM�c�N`�,H]I�d���S ��� ���+��_�b�P���h}���|��{��.ʘJ����8K�O8N94��Z}�4�]� ������3�kP��I$�I$�   ���2��v���HL&�	2�	���7U�ɞ���+��賍K��N �\����c���:ڍ�܍۫W�t�3t	Nu�6��Q(�$���"<���6-�d��dm���������,�S�l�'v�����#�=�Sl���Io[��vgD^%�0iqő����g|a~:9�V�C�G3ٳ�����������N��])�����k#g�n�1m^T�C�	�l���mw�ڢ8��D�Z�_��}빠޳���<�����h}s�ؤ9"j<�7$`]��]�0�.0���~��{���F�Q�I�	&h�~�}]V�f$}��}������N��s�3�u&w%�vT��+� �,�;�|�4��"rE26�Z}�4s���s�K��.���m�$��$hnɭ`ޝ�
��tR�zRu{lq��m@�c8DC"��m�$fF��NM��s@/�f�_WU�޳@�qV���]M]Mk&�F䝾{��X;T=4��9J���@����9{�qG��7z}]V�_z���s@�ޯ@=�4�VcH�byJE������0=/�6^��.0-��i8�9"j<�7$�/�w4
������ ����}�}��I!�)�2`�[S�u���D
��k��v$�L�;^�qX�H����F�Q�I�	&~�����h���/�w4ޏ�:�M�n4������K�쩁vW�͗��;�Q�q2H�m8���h��70�ꤑ"� ׄ����!w�КUł�� +�t�! zwÊo��NP"BD�%<dF�!I$	HD!HŀHäu�� "�J {=qH&k��v����0"�"���	XYIYH����8x�^� TC��BF�T�h ��hc �RD D��P�%��O=�έ@#�C�l�|p�4� p^�W�U=PN�(h4�A�5��}��'����I睉�Ll����I�^빠U�W��j��Y�r��u�F)�n.�0.l�`r�`eL��0=�����o�	$���+̹k�'�{N�֞ݪ���(������Z劻vn'���.�uw�L��vT��+�����sOf$��'�ĤZ}�7�P����ӯ� Ӯp�5�tG�8ڋ#M�4�]��z� ���@/�f�}�F�Q�I�	&htOV�� �Ӏ�w����$B���F�O<<Ϳ���:��u����FsWXܗ�z�|�|�,��$���S�Ys�Ŧ�4��\4Imt%e�-#�F4� ��l�A�#Z���'N- ����Y�U�@/���;�vx�#"#�@/�f�(�S'N�V v�����9)��.����P�rM��|����>ď��h�~���î(��ӀD�I�]�q�Y*`eL�m9����DȢR- ��h�����`�u�R�B�$�R!$(�����;޽=����~��      Gnr�i����kW���w�UC��yӶ����f�gi������[�w.�p\.(��Ñ���u��)$tgO�(�i'`�n�ɂ��U2e_.l������l�с�����r�kf�d��F��(��#�^:�@����F���݈�^{u:��Es��Ѕ)ړ�xruCV�(Gb�S>�06�����%UU��������؂k�2����s���nd�Vݢ�8hݙ�gs�Դ{�|`mL�K��f�}�F�Q�jL��@/����f�}빠w��N��q�ޙ�a�&w%�d��vW�}�h�5�D#����iš�瘗��`z_>0��w%�ڳ;�bd�d��nM��s@/�� ���@/u���d�L��!(��ư[sk�.0qz������a�ڌ[����ZxF(AB'� ��4��� ���K�k�X�B+��"��57w���9�
���D�7� {�3@/�� ����Y�b�"dQ)�Y*`]��]�0�.06���##�"�ŌMɡ���߳@>ﾚ}]V�^�4��pj7��P�q�]�0�.0%L��0&O�g�XL�1�Y�,�	�e��#G �����y��ƻ�-��<Nn����c�K��K��S쯌�oX�k�&�I$��Ӌ@/u��y�y⓵�,�{� Ӯs�Jd{�3Uw`��� �}� s�u�'H� �R  Dd`D�!3��I%0�y8���-K�u�6Y6\�լ��z����_N =�x�����0둍�ӘFԏ@/���B�:� kŀ9���:k�����!̤�4��W%�9Z�k1emNss3����Ջe����5pq1��ĳ�[���+����w%���.I9Rcrh޻��$|����_N =�y�(Jd�+�����j<bmBI�˾���uZ}��bG��4����vz>�cq8�ORI�С(S=��p�����X���<�<�'yl�@�ƺ�h�8�N6���}%L��0���]�q�o���:F�ěF�.n�i���H:&b���6F�,�hd�^�o `�d��NƋ�z�쯌�0�.0�T��qV�1�
8�h�z� ���@?{�h޻���îF6Np\P�.��>�S=��3=/�,��=E9���Ĝ&E�h�z� �׋ ���0:"!L����6vZ�$dx�QI�Mɠ_z�h{�~? v����k��KH�&�$�
;��u��޽�޽��
��      �8�w�{X��7U\q��3�aS�����Yi3�͒\g���؊|�tk��!�u��ݣ����F��k�$�:�c1���3[`+�ht=YEBvN-�։jzס㭓d��n���f��y����ј'N�N���Y����k�`5(��@�5��n:۔�y��]��x�[���tf��e��>�{��| ;�����E�Y�Yvy�ήӶ��ӻ\��q� �5��p�{\��l��16�$��_���4��� ��Y�3��>���s�q����x��$4�K��0.����b�o;��:�����iŠ��4�]���)���h�Ct��F<���ɠ]����Fw%��ʘ-;���"q��?{Қ}]V�~���/�w4���I	�)��5me�M&�G��&l�62.�ơ�v`[+�����4���4��� ��Y�_z�h��M ���<E��$�2)n�w$����|04�>,`m��5ݚ����_WU�g��˕ϲH��Ȧ%Ιޤ����튌�K��h����n517p�?{Қ ��s���x�DOk�0�����'��B������f�}�M��)�}���>U�$�O1c"I������]v��:V2m]��I��J�r��C�$Ꝯݩ��D�dq8�q~ ���@�����ޔ����� ��M���FF6�o`�j� ��� �eL	������"rC@��Jh�uZz��1E �F)�֧�ݚ��=]�qLx�NbO	!�r\`l��v*0�9�+��'�V�#�bN"�H���f���g�}�~?�Y���h]vI$ƛ�	��W:w\���%�HL�a�l�e�Y���8�Uƹn��T�.��'�����튌�K��0.����.�wy�;�B�lT`r\`l��}�M��3<ċ����n'��B��L���ʘb�튌	�����D�d����~���/�)�9��ܟ(kH �@�^^}ۿ��{�&�19�(�ɠ_zS@��J0�.0�T��*�I!#�w�����ջ'<������\D�ղ��n��h0�@�i�LjL����)���8��w�!D/����6Z�M�1�1)��������H=���>�>4����{L�"�Kp�JL`l��v*0>ب�.����;.G�5&A7&�}�M��)���h�z��;����j<i%��*0�.0�T���z])��4��A�Z'6QX�PڱR�J��x��4$��� ��:Q0#��Q�hiA��b@"Ł�7��U��	 �d�B�S8�)�dR,�)$��� C@z�F �"�B?(�Bx�H���>$B+'�`��KsR�R%P$VP�$V0�A���&��Z�D�<�Jmӫ�JJ�*��$&��0�$H�m�� �}QB�0~"Q~@ࡾz{f9�`IJwIvaSlP8ŀ��"D���ȠGňD`a @���%A���k33Z֍kZ�MR@��                     ��           C��P������͙�\�f.�;�����N��;�cQ�6�"n*���e4�Ηnwc#	E����!98[�*�lS��v�Z�4%Gb���ʫjU���z����T7�/Sw�^q��[�ݻ6�lJ�k���6^�Y�6`wQ��p�4ֳq6wd�<�7L1��<���9��N�ggtH�E\��S�:M�P�\�i&Y���4�6��g-v���ac��Z�[t�SK�#�ۮc+m�J�N{�4�6k,�ιmH:G^�mtд�[	n�u�y��8-]�)6���v��/J��y�:�i�]���}&�5S�9`- =n2��kg�R��'��ͦC�	�&�j��2�ԫ<�"nwe.��窠��;�6gƝAГS�DJ�	a��-�veb�U\�)lF�.����.����cur��fV�#�����-$��s��+��uJ��5Uئy�:,ͮ�'(Xs���>F8�V�B6���H{-�sK�.QL�`�;��v����+qc;W[,p�C��;.��m<q�R�gc��i	g�D�������55�Kj�q�&ј�;V��9\
�WONa��c8�.D�e�m��%x�ش�c�B'/ �k�vZ2e�`tnm�բ6R:Ѷ;��0U�ˤ��bó�u�����&Ɛ�u��Wu�h�3��t��*�ܸ�Ѥ:eX-E�����j��T-���Y{J�K�-��Iד�q��=:y��=gŹZ�m��k6�m�/}��O��X��F:{$�y�und��삼�pڍ�i�n��'����9�/ P1U�j����p*�vƫB쁬PhO;{����ۄΰ�J��Eǋ\pslݠ+�nK��(���<my�j.������# �z�����t0O�Q`��ϕGb'��E}�����WK��=����|�w��ߟ˾�`     !�h��^:�t3�&�ݦn96u	�nٞl� 6Vy�\#�h�r`����oD��Xv�GL2�!�6��u�a���q���`��'@����F�v�V��uґ�)�m��k����'[���Ãnz�h��جf��)�cv5���[�n�G�Z�T�2���l�9���U�yOGn�]� �����8�Gf���%ik~�w�w��/���7^��s�z�On{sW3H�a������ZĘ�/��6�n��V)l_�uu�����ʘb�풚{�덢E#d����~����l�?}�� N���D(�����W�7"J"A�4�ύ��)��g�r�- ���@�ULT�cP�y�	�Q�]�q�}eL�Q���a�ǌi�JAHh�uZ����Q�6*0s%I$�pHY��`�C���+�z5����J��ӷH���ItM�\�3O&%�8L�%"�׬�/�)�w�)���hz�#���֍K��nI�=�f��|i 0 !K�h��pD����.[Fmߌ �N�p��y�;J��Q��x�J�@�gƀ_WU��Y�_zS@����[q��OĈGf ?�\�����09B���ߖ{~�ґH�2D�iŠ��ب��W�w%��mI$�YӮ]�f3�Y]7g�Tlڌ>a�v8ؽ��9��{A�6҆7"J"A�4�Jh�ŀ��<�~�;�^ 约���l�h���0���Q
&C�_N w>�����
!B�6Z�M�TTթ�������p���J��t�(Z�!DF(K˾0�x��-��#�+p�JE��4�ՠ[n�^V��G\�L���&	�4���+����s�8 �w�?�[�t��Ď��CM��v����9(�Y�ڀ��3�+���t�%�y ���m��̷����w;�8�q�c@��@/+V�[l�/;V�[l�?{�뉥"��d��Ӌ@-�h��@-�h�j�=�,iS�% ��j�ou�$﷽����v�$"�n`���E�o��zܓ��r���&5&E�@-�h�j�m��j�?W[�I$ �%�I��y���5�ܶ������U�W����:�\1Wn��1�1(�rh�j�m��Қm�@=�9���BppQ�' n�!L�s�0���~�s�r��"S#rF�ɂrM��M �٧���h�}��/��\�G�$�7 �٠���f�yڴ��q��lƁG&�^V� m���s��xG(�]P�ӽ�t�{����$�      �n�$v��M�\��-��(I�k����8��k��e�A�˺ݝcad�����Jvc�f��弖Z���o������Ŷuk]c�c5s�	���lG[6��G`� F��Bfs�-�h�0cp=s�щz�0Y�kQ�u\Tt�8��K��j�t#F[���p�=���sϤ�vl��=3]�P��ٷ���{��{��B| �.v��۝�ї��b�Yb5m��c:�-���� �7R)# �iŠ���h��@-�h�j�=���LnD8�D��hi��BJ!L�wu�9� m��^f$U��i�a1�A2(�Z��}4�h���h�a�\J`���F�@/+V�[l�/;V���}��M ��O��,N
5"�mL;n0mL̷̭$���t�/JY����sX�
Z◬�������̺+�KDW=���Y�q�[j`e��-�0.����F�ƒQ��[l�<���3��U��4�ՠw��7�6�hrh�j�m�}�g��%�|���h����5	"ddm8�������f[��&�1�Ģ$�@��Zm�@/+V�[l�=V�$�dq	FH��D�@[sk��U5�{r=v�+���j�Z55A��ơȣqh[^�^V� �٠^v���0�L71���L̷����������T�X�jE��4���b�V*:+U�CJ���@/.�@�W\pS#r(�ǂ����s��x �[��3��x���}&5�$�nE��4�h���h^,�I'��"va�'h��i6KZ%b�]�g�l��E��g��bi4ڃq��lƆ��h�j�ۼ�x�"~�;�� �QO��6I#�m8��f�^�h�� ��Z��6��H% ��j�m�yZ��f�k��nU6Y4\�U�DBS=�׀�p�w��'WЂ. ��%
N~�8�BA6����swWxf[��S�ی�Sm��@u^����I��X�W3t7aX��pӂ�5�5�e�:zwX東��lI"�m��j�*��򼩠r��8)��$łrM�}V�[l�_�>�s� 绫9%2>��:�*ڄYJ7"�*��^T�9[^�޾�@�>n��㑳rG�~���e�X�Z��e�u�j)�CP�&G7$P�9[^���~_�s�Հ~���WD+��W���5Www`     �I��^�������{r�����c:�ѹ:�bq��h�w#G�:R���ѹ��n�>�\Aض6,t]se���+�e
ݵ�a��8	���v�st�%����Ns��N�^yn��$u]$E\�C�;s�$iGF�uFz`�v��3�S��VA�Ǡz�.2]V�;���2ɝ�"k��v�	�U�>�Vs���O�Uv�c[.��c���k�ڮ�vk<�s�I�׳D���ۭ�8�+P�$L��)�}���h��@�/e����H9����uU���,�-F��9[^��^T�m�z����3����70����^T�m�z���k��Qc��,A�jm�@�_U�Umz�yS@-�
y�LX'$�;��h[^��^T�m����I$�?���������&��:�NڣV:�{v�aMms8��	�ْ����o���7�|hw8�����|�n'�QRUU�� ~{L�

!T(�
m�޾�@����<�ď{*��CP�&GFۆ�}��M�}V�U���Κ��T�@���z���n���f%
"g����]Uu�1�A��7�U��f/~����}��������I	�)�8J��z�+k%��ˮ�nS=��z��f������10na#�= �y�@-�h{�h[^�u2���`�"Q�0mLYS巬Y�0m�7"$��NI�z��k��{B%Q%��4V�����9!5���h�U5�D�A�!	xM9�"�M�:C`E�눎b!�j�hxI#�_tYST"E3����2IK����D�`ȱcI$��v������*QL!���2#Q�B8�)�p���:��H��<���t��$XC��f�EG �ͤ�Z�`(8�x.�
/���4C�v��ǂ���(D܈���_���Y9޽4�f�ժ��8�"ȒDNM���� |� m���DL�}z���7�D�hm��u�M ���%�0.[z�4ܝ�$���3���i�x�k����"K���+=mv$�]�7����4�s�$��E�6��4^����� wOt�ں��uv�6��@-�h[^�Z�Zm�~ď��[��Lj�)$�>]�X ܷ8 �w��x��#\
b`��Gzj�h�� �ٹ"��.�Dp�Q"�Y0���OM�V ~�2UuЉE+)\��Zm�@:�4
��@:�V������?_w��\�fćhӭ;��`:I`��UY�ІWk�9�%�נV�A24�܊)1�����女U��Uj����h�>pjdI"'&�U��Uj�m��٠w����r'�CnH���h�� �l�*����GqBH�$Yn�L�w^ >}x��`��`�#u�rj&�c�h^�@��X�i� �w�%�$!(""���������O�zۀ      �b[2M3��8�Q�� 79"N:۷k���ݼ�#�g��W1`ٹo;uF���9K�:�v�Fͱ�A�j�Ƽ���;�7X�lFL]f�"틱��pm6 v��mq]�I��e*xN^�Wk	��hq�.7>�[c��m/�ڸ(�ZndJ�ck9��s�t@���u���i�h��H����{��w��w���5��8TՒ7�����7=.����[�cc]�V�V6l��V}�g��d���=ΰ^�0������4U�����70���u�M m��z� r۬��o	����X<�Ȕn��}4�Y��4�:h�����Lx'$���m��K;Fm��/p��pq�E�$���Vנy�@-�h^�@=;��I2�L���o�It�7g����Zp⳶8��u��&���,7�4�hi�&�u�M �٠z� �٠w��*��$Lp�"mɹ$�{�o��v�*���&k]��-�4�t�/vF����M�Τ���m��[;Fm��y����1�F�A�&�[l�y�@-�h�f��vu�S�,�� �v��S �T���������@t�H���&�/n���1��3YǗF]�⦡gs�m�KH�;�slp���]�> ����%�0-��KΚmUG���ǂrM ��h۹�y�@-�hZ.WƤK#I94m����y���<H�<H���W
A�+�([������׀n���mS*�j9��� �Κm�@:��m�@�s�UBH���"m�@+n����}�;�� 5�3 �>���F��Ӧ��j��u�d���g�g����ٍʹ��n�<����iI�I0	eL�S �v��SsK���cPDy	$�m�@:�[l��f��vu�S�EԘ��`ژ��m��{L�c�`,O �%��[l���nI;��[�E�GpF1� M.v`�����U�G$"�	�4YS ���%�� �����j@�����Hi�]+�;kfQ��Q������5x�
�ih5�l�A��� m��{L�۾�IB_�ϯ ����q8�OĆ��h^t�m�׬�m�{���jD�W"���0�� 5�:Q2ww^ _���/vF�<�B'���x���0{�LY�0mL	;����#�I$�m�ם4��nI=���D���FAC]3���`     *����[�ܑ��q[Ies��u��Z�M��B�gW��%�pÀ�ֹ���|�����ͼ k��d���j;�]����gvc��`�쩆
+�aG�X1[rE�mv��E9��S�`���cu]��F�����{5��N�;��;]$v�V���m7km=m86����rΥ����2o�~�w��������	:Pt��s]r/C����.�V�m�=��g��v:�\1Wn��9�3_Ͷ����@-�h^�@����gSby�(�4�f�u�4
��@:�[UQ�drB)1���@:��Vנy�@-�h^+�@���$D��*�� �Κm�@:��p�ٍ��Q?rJ�{L�ۼ ׮�-��<�~~o߷�UW�S2��v�����X%)w-�c���� 	��l�t��92Za�q7SUg����z� n�?H���>�"c�$��rM ��k@� �H�4��*�E�:P#�NI>��u�$��t�m�s�ڳcpQ<�rF�oX��`ژ���8!u�)�s#QǠy�@-�h^�@����gS��"Q��S �T��m� �v�~�����?�Ut�:v/RY��!�
�t@X�lc��l#���d�tFC��"K�V�1������4
��@:�[l�:�\���Di"'&�U��^t�m�׬�;��[n7sQ2UU�� k�f 6���#�%EQ$  k����krO��w6�9EP�#���i�h�� ��h[^�u�M�dN�	$��X$� �T��m� �v����I�;���o�w�<[+Nm%l��]v�S�ˣwi�܏]���3]���ͩ*T��cpQ<�rO�|���y�@-�h^�@��.�(��9�������4�Y�Umz�3����ĞBdJ7 �٠z��k�����Jy�E&<�h�w�9m� k�f�TD(I���X�S	X� �,��d"�����2s�� �)r갻��4��@����:h�� ����I�=������?�����擴Y�R;1ֻ%c��7BMϲ.��K]�6x���\ˍ��Hm���m�@�ҟfg��|���{J�>j���4�4��:S#�|`=�X�i�Х[�?���	H5$��ύ�k����4�͵f�ࢥwWv`tD%	OWwV >u� 6��zS@��.�)�ә�= ���(Q]����gwk �$�W�� "���UAW�  "� ʪ���U_�  ���A�A � `�P1�E d dDPE b
DP
!@� b(��(�P
�E b(�T��@�E `���H"��PE�  ���UT� �� U� "������UAW�� ��� *��UAW���
�Ҫ��⪠����e5���A�`%� �s2}p��    6��  �    
Ъ�}�|       ����*�J�J��
U%% P  �   PJ QB*�Q@R�      c(|��MRž&�νw�s���Nr�sb�su�&���'�wǀ>��R�����c�zyeW[��O� ��O��=�����_O�     >2�A��=�<�&�e��,�����
  �  c�7Y�T�m��q���;uL�,����qh.�}�qj�n\�����Q�y�^�x ,���^�](��
��7;וqo��͗M�ut� ����7*�\�˛t�����x   �(( �1@;�V\a��Y��j>O�ײ�8N�h(�@�v`QO�; �� f �� 	�  �   �0 � D @  V    �    ��  �` � {0  ;2�@ � S��>ϲ���^l���ԧ�U�}>W޷�i^Mp >��ez�y����
�Ҝ���O'�m�﻽l���y�[�����S�����z�nl+�  �  P �$4��Ln��m����rysqp�8����n}���x�|����g��m|x
U�Jr}�q�p _O-�os﷗���9�������δ�ӽ�Ou�ǅ �Id���ϭ�w+�q5� i�
��R�@ 4 ��jf�T��4 "x�T�j  '�U%=�(�@ ����%JT @DHjJH� h�O�?�����Z`����m�����{���w�U�n_�P]DES��P_��*������DDU8�����������#<�E�K�L3$,!�@��Y%Y�I"J\`¤B�� @�.s�<s��s����I<&$��n�)��n}LU���[y^]�g���(�u�������1��e���o;#��`Đ, ������
}���Ɓ�2H��!�4��a�3�H�)����I�♐�I��O1�aX����U����㷹Q�)A�15�3���/��=,~���y<+��Ͻ�4%�y�f�a����1�L��0��c-0�RL�RIBV^w˾nO4���
9>��o�B2L��R_O�H߁��@��Z�0(`B�/��;Չ�L�4� �\��4cT 1 �b5�SST0�QB�op�_9���HS=e��\�YsM�4�\4#R!R\�.o5!La\ԅy
a�)���@�hK���lk�i�
a�	sy�sSSS<T���F�T�$!F)h�G�FV%B2H�P� A�ђ%
 ��Hфj�\��]��$	¤v6aD���9��n�3	��J���XS.�6�4�B��L�\aBZ�ឌ/��|�`�A��z����͒��/��ٿp8O3���p��$�+����*O]!�$j�D
9��\)$���P���B,�_��$���<a���ߺ0��X@��Ȑ:�=�B�,�I,-u<5 ���"D�xK����������v������X������ς\���Xsﳑ!�>�2�7���0Ӂ)�Xn��] �5�l#�e�ӛÇy��s�0�D �<;���X�@�H���E󹰻{�Uj����b=��)+��0��B�14\	��5xz�4��{<a�� �i�ͯ�	��%5UU���Fb���m�E!"P��-�	�Ze�*��r�QEo®�	q>�=�]Ð�\�������o��	�C6\	y�򞙃 D��b@��H@`F!B@��0��}�M�Ys��]�� �@�Z0�b�YK���M	����B����_d��J���+(Fp#bD����[��i��{�;��hRS�L;�f�HCHP�FVXؐC@�$�/��sy�=�w�ac�y�J��qЍ�W_Pꨥ/G_S� B-*QH�s�3lߏ��s�^p���!��5aX@�b�CQ����S=7�}�^��t�7d!q`P��@�B4H	�"�"�1 �"T�ЍIsy�.�y-�u����#���߼<7�48�F�4�F�1h8��'�		�F�B*HZV�R�n���0�4P��t�30���,�'���4������ 1$
$B,� �,B#����J�4Ӟz.�$�}*�0R#`	�� �X�bRR���J�+����q�P���c� ��-L$X$#Q c A�ĂD�b(��0>M�!\%Y��^��{���! �0`�q��H�Q!B��D`j: 415xF�)��������⑤K�c�c�+���4%�
Ƙh�J��̦��@�[���ir^{�����0�rn2��'7��=SB�qH��)_�JF�m��<��M!	o�x{�c�3M9<��y��U����=�i��W�n��/-��t�/L#�hE��h�n�����3�i�i�}�=%���Fʰna�����5�F�H�%
D�E�=l���y���#10��e�@�%p �XW���h@�*F�=�����^�_#I7ФqaV]氦I�����o�.o��!-����ϩ�H�"D�xh�&��0�G�e�b,b�21�+Ba���}����w�i�B0!�
�)��,��fsc�Ӈ�!�Y�2�C, ŁHЍH�H��Č��wR�g��_�܅�5!q�\I�CsHsxÚ�%p�RO3Ͼ���c��L~���"@`��t�F,�y�z�!ML[�D��Z�H����"a  kǌ*x)�ϴ���4��_4�����߳7��\CK��;�38y\A�XP�D��$IL�fa�j@���H��MVA�.���O�|�9d='�4����^Ji�W�YO�Y�).�.� J$�`��D��	�ϻI{��C~��;nY9�Bx��rDə�t۾��}�J�l J�F��{�����9(�4���cI!�qӞ�i�"j��|5���y�}$C1"c,��R��-�t�ZȄ`!�@b8�`	���y!��H�H�1�BV$"�E�BBBb��HXubƇ�k�
B �E�$A�R�`@(a����X��O	���M���y!��۬���ύ=>�ט��2�h��B� � � ġ�%�:vLg�P������ ������|�l���[=ԇCۜ�s��'������+/��� �Č�D��)
Ĉ|BBa	
��s ��������"e)g�#�>sxM"WJ�I#RR� T��>R!Hz�S?9D�\	)�b�H���B\ԍ	x˼L�������Jkٍ�eRŗm�+�K�|}���(��������5��3��L�csǐ'7��(JK��x����%�eٱ��)�w�,焥�rr���V�7p����&o���.�Ի�a[�������k-��yXp����v�m��<��7o���'���
��[�^i��w�{u<۵X�/��	��9O)��㻡æ���}�-}ɾ�2y�B�K�L4!��niye�8���p�8x�+�=燋<��.���K�e����i��tk��~����ՔS��-�=�Kw�?nn71{WZmB��_ʦa�m�x�h:�����k���~e���'�s��3��3�ߏ��%�!o3=|�B���É�����S6�"S7�\�$瑃+2��xO9���q��Ia-"F6f�-�HdI��KB0�Kd��;p̙��m�7�<[�{c>˼{�2f�Ny�7T]��!��ЍK�.7���fX�����й�G9�6_:Ne��e��,�%����HfaϜ�;ӏ���������!Y"B,H�\��|�s�t$��	�=��|x��}a�,��Љ	�(B�7��H��g=�~�V�[¼��{���?|}u������3=�����<����$���p0��Ȅ)��1$!k����m�9�筐���D����W�d�X�	qٚ�|�I��>�\�Y�a���w�3vxO'u�����W|�w�'���@�J��}�����                       h                                                    m��                  ?�>              l                                         �@�H                         m�  -�     �          ���                   l                              �@                         �`      �|                                                                             >�                                   X�:I�������Zm����*���{��\��zݪ�k(�JU���S6v:�ٍ<ĭJ��R�����lfZ��Ð�yV��-�GG�)s �"n���D�.�ˤl�I��|�$��ےA�U�L�f�/:�^ѱ���e`�{F�!]cmZrs��@����c�=���b�*���k�3�[�M����LdZ�x[�!8�:��Np��ծE1�����T5��z�nЭ��Q&��I�Q���p8�c��m-j����ƸyU��t�:((8 r׮�,��l�@  	 iͮ��eZSi�VV�nڞ���`�� ��m��v0 m� H[@ݶ�h�%�-�m��m��b@���  H�km������ʪ����	��     �6�  5��ٶ������ ���x��z�+rD�ť�W��j����lj����	�͹׸]�l]a�`,�`27m�u
���yUZ�c�mN�Mf�$m�`��,��Im��sm��   $	����  ��ki,��j@:t�ւ�2�h�5VQWf���m��n� 5�m��  n���IqUR��U*ԇ
������Mm�6�� V�#���n���UZT�q�|�Y����Wd�i{-�l�K�=��(i�q�k�痚k��P�'ee3���۫�` @�f�v�'iI�[U��j�P  �~�| 6��ku�D����k6H�:I&��	 J^m&-�.�86Νc-���z�T�	��:�@ w�|    v�����5K��%���sU�֊$nӦ�-�o ��m%j�mh s�)�ڇ'�F�j���d��k7m��lXmk2�f��mv���y`�p�9�n¼�9B
Zܓ�V���AUs����;@�=��ݜoy��v�*��Tg��`�YV�����ܪ���2���<t��i�=v�����"�Y6��Q��`Rܮ�iU@J����;Q/m��,�Ѭ�C5��4�'C��am�m���mm� � �`�[� @v���������ms� �m��-���H6�ۤ]np���
��UU�� d���T  �Y
v�� 6݋���j� �Z���VKm������ꍶt�����	�kt�� U[m�V�q$�m�{%�H5�,x��ݭ�I[	��%�pN>/|�erU!J�6ܚV�UQ�gcq�sMe��[6��o�lN��6lNn�a]&�]�eeK-HM]Z�n�؝Q�U�ei�wM&���Ŭ5�I,��OM��i�Ŵ�J��PPJPur�no;$�8Ͳ(���6H��l��h<��@I�m�nٶ� YD� �  >�N�}�� �m���R�WK�N��lsd��IL鳝6�i0 ��`6�m�f��\� ��`��V����j�p  �` n^�vݶ�d�l�:ې��m�   h��t�`��$  H��6Ӭ́mK�i�@���m�XA�#̫�
�UR� ��m�m,��kR ���lN��mҶ6���@-�J6Z      [@7p [}%� p m� e��� �� m�    H  p�� �`    	l�`-�-���ۀ��  ��l 	     l    	��`�s  [[ֵ�lݺŒM�m���  ZM�c���m���Ym�O���l h���kq��� �M)k8�F�6֬�$%q39�Z����mT���W-.��8���n�   �` @ml�tU���[W$$�&�L���gI-�h  ��9!��$6ZH�	�,�Xm�e���@$m�  &�&ٷ    �  ��  -��:md��oͶ��� '@�    ����    @  �`�`   8 l   �� �  p 	�  m�      ����   ���6ٶ�kn p^��R�,����];9�[y�[A $�V]�i8 m�[-��M��� ڶI,�e��m���m	-�Z�6vy�e�e����C�r�U�  ����hN�I�pll ��G����̍d�-͝�D� �  a1�m%l[du�kk�-�[@   ��(��  [d  �� [@�  6ݤN� �  a�    �~�>�� ��� 	h[v�7־[D��/ϛ/��cS�d���e� )z݆�M����@T�Q��[J������^����p ���  -+i ���n�����z��` ��m������$6�'@�Q� ���Y%���lN�[�J�0���5,��B@m ��6�mHݵuUP
;�ڬqg=�P6�n0��Umm+�l�Sʨƪ�r�K��tU�*���P8	F��w<��Ͱ�n�0�-�F�k�7D]F!I9,��m��Z�7T�p��Mn��9��2�NiϢ�4�-�v�r�֪�Wp�U��U�㰣@�m��lq�  m���Y�U�����aPv��U�Xm��[` G6�D���zk�6��͖v���ӎzMGIz� 6����|Ζ�z�l $ z8�n !��` �Z�䅴  ��O�|nհ���  � 8ȶ�=�,��p��� �]-�Yl� i�]6l�u��� �;v�SZ�4��-��d��9��٠<yݝw;p m:I4�Zv�ol�A����P����
�$  :�[�f�"��M��-��b�$H @�Asm�ۀH֘[�����j<�G'Pfu�;l6����J�'C֛K,�Be�N�S���9Kh�>
km����t�t����¶Λlm�DQ��${Ur��*U�V����n\粬��P���v�Ǎ�N6h6Cnnݝ%�n�n�:�n�6OM��ىIV��󷆕m����6,�ՁoPm�H��ml 8ݲs���ݤܵ:��o � ��  -�l�\s*��l9e�j4f&�loԀ$��m�( $.�E$��fj�j��G5<�/0�	6�mjKpAĒ��
�������u:M�-v͕� �ʹ�N�,�Mܳ��~O�� �j��ݐB��մ��Pp	[v�5�Jv ��"ڱ#$�[%��$��+[%�!�� 4��=0�Qt�*�q�.��~���m͢�ʸ%� p gI�am     �m��ݻF�  M�l�tm���`����8����`H    m$�,帶CAl��4[��P]s��C2��]V��5�� $J�]�λ�Mu�F3��3`	zT�U�K^���÷bi���	���F����������0�!�5�<�<Z��@1k1��9�n��[���A���]r��	h�B�5�����c�Z�� ������.¤ZXvh릂�����ܹ�rI7f��(�����#@�#T��S� "���$"D �|j/�<O�X������A�@ u ���5T�	��AB�P>A��1 �����!�O�b�C�x�8Rq� �t�Bx(��B!�&��R ���
��T��⨇�� "q��x�F��x®��Bh�U"9��R�r
��֢�zj�8����TD� *�@����V�S�h��z
����T z�_P<@�	��~C�v"�*'R"� �.�����#@���h<qT:����H�R��%*�aD#X4`H��Y+2��1G��:OD=�L �"�O @�0z"�dN�C��C}�_���*��p���)D�-b�D��5���Ţ����PX���w����{�~�  � �          N�  �� m  @   v��   �h ��         .�    � �`              �      �!on�$7]g$����xN*8˃�d�t����W����4sʤ�^��.�]��n��3Z�Pw 1�����n���U�Gfv����l�D��)�v��4#ی/'�ח3�v6�Ls�� ʗ[-4�1�cs#V^9Dj�9����a����O8pkx�z-�.zι��C�����3���H�f�MVӪge�=�l�e���c[d�Į(�N�_<s�pql��&��uc]�����hT�A&��v�. ���p݈vx����Y�Ѫz��u�b���8����Σ������ӈHZ����md9��Oom�g�a�ɭ����*�v�r�%J�6�bUj�)y�۲�����n�go]��m�
!�"�ٖx��	��G9��D������4ö�ls�Yà�}���UU:ʽ��!��Z�в �]&�ڇ*d�I�[UUK��-��T2��6�Kl���g#�&A�]��<��lT5�P� ;N���V�'`&�b�,$ZT6��[MN����c�玻XOn9=���k:����[r�I�������!Om�̅FΕ���M�:>�E��θ7]pl���'C��Xmi�;(WE6u�Ӆ�n[(�����n��E<Ġ�xH�a3�{:��[��cf�.��[[��{X���m�WD�<pM��X9�==9ۙ1�r��x���P�Z-�J�,��'[���nl%�C��U^�sq1 ti���Yv�I=<��j�i�!n�Ը6�@�8`��U-$����%�
�8�Δ����8Պ�Gr\��.˗	�v�����V!�R��|

sP<E��^
����ꏨ�>x���{��~~�	  R���h5�a��m��  m�  m��6�u��ڶ�=����lẃ�-�U�W�9��'/��/Fn�0Y�N2�-���Y4����q�PYfs���J�C��F���f����JN�s��Pk��e��Srq�mm�g��5[�EͬĂ�m�<����]9`"9�s���ơu�jۻ-�L�&L�ߑX��,��d&��c+��=�r��ɶ0"�nQ]��8;�8PQw#T��P��C��ŀf�_ٷVs�V.Grd��tۅ8&�`�1�����r&���]>XXJp��ے��7���ܬ��U~K7�� �w����c9�D��U��r&�����0=�0=���ʉy��ĳ/��� ��ގ��ܬ~�_����H�0I9$�)�i���D\5�<�k����,��j��]�톕3u��7NT�I�|��K�޺�7r�>͜X���J�J:�m3�?���UT�	-�0=��`����`k�Q*Q�6(�%X�"`n�A�l�oGL#d*��$B�Ɣ���6q`����7���ܬ\���%
�)�9*�6t����mȘގ�����)���l�	9�U˹1#\��bz#��m�Qu��Z6�ʹS��[�m<��w��7��Lۑ0=�0�1���ڮ��tH*�U������o]`u�p�׋:�����2������������Z�y%"�B�D"B�y$��޼X��8��y @ܢ(�m7*��{���7���ܬ�z��Ŧ��TjR����������r&�����0:m�}%��1U�4��
�ӺW�of��6]m�8����q�v�ہ���6��8�ˌFfS��LoGL��`{z:`|��)�9"J�R+�޺�U~���,��Ձ����ˑܙ$�T���VM]��m��kŇD%/k�l��Հi�z�IT�%'M$�,=�xrI����I=����*����]q`j�mWSn*$	)*��}w����0=�0%I�bʽ�j�s�W?��o�[���s�Jľ��׶��rPa���Pλ:�^6�G�Rc�m�~�b�<�ـ{��}�A�wN���d$�:�F�qX�yX��V��V�����Mo��Ӕ�A��R+7��mȘۑ06_D��4:�(�(�D��=��~]��Vk���������u`|��)ʑ9"J�R&��L��07dt��*������~�  �` �Z�v�`8��}�    /L���M/1���˦��s@����	�ێ5�u�[�2d͹c���-�ݸ���kA�ɓ���ku;�v�q�Y�4(p�@l�U�ќ��-���zz8�J[� ��-t��]u%��cF�t��Йui6��oZok:�[�V\X�fe�[љ掬�kf�S��w��>���M~+F�:� 9Ĕ�YӃN�q���X��l�A[�����@3���S�R-�?yX��V��Vc�V���8�9):i&�3;���"`ñgd�#��U�N����	,�`v܉��#���03;�����B��B�Q�`ftt���쎘�"`z���$T�q�ܫ;g��u`n>�`{��`$�!v�gM��)$�����fB��]j�,�ܾ��[�@<��w��[��g�XےTi�p#rR���]X��X��]
?Ho;� �4r��*n���X���݇�U(HP��P�y%
ԋ���b�?s�0�ot(����x�?4�4�4�V�z����Ł����L�:+32�,U�M]�P���`��X����ו`jރ��d�I�I'�7r�=[�����,�{�)� 5U�z[���ێ�l!v���Σ��v�e-��c��d��q�:��
�o���L�06vA��#���YB��aFe���Lގ�; ��������XV��T)"����X{l�?y�X$�D�	%�E޷�p����IQ�)ȓQҎ��遽�107z:`l�Q��)b�Q�$�`f����;g��u`n�Ei���D8Inw"F��ڦ0O9Œ�:P�ܕ�1�Ѯ�i�9�6Jb��ۑX��Vv�,�������X�ɒJAT�rSgd�07�&&�GL�]�:�Jr�7M$�,��7gE`n�遳�#WU�R�����HK2�ݓvGL��`}_U}z� u1�~��rI�^�%,�3�������=��`
o<���ذݝ��8�q�  RI)��������ㅢ�q����m�۱V෵��Rq���|a����&�m���OguՁ����3;��Zk}%F�)�t�����遽�10=�:`l�������t�7 �P�7gE`}��Vs�Vf�Ձ�3��?$�1P�mȘ�06_D�ݑ�{�b`r��L�R�t��;gguՁ��w8��, Z�@�7aawwwvm� [Mk���  p    od���>u���ӤW���-'&�`ntk��U.z�ۑh9��'����kF�iKH�N�ٹ:�v�t�+��I���k�iKN��9-v(�e��MZ��@�'n���e�.ё��f|��l��lg�]�u9���\w/��k�줻I�[��v�2pi� 6���2��̙���1����6�ۦCQ���kۮrqŴ���1�O����؝@`�P���7����/l��vߟ�07�&&쎘; ��5uX�I�TT���7gE`fw]X�8�3;�����B�}�F��+6d; �ݑ�{�b`z�r ((�m�;gf�Ձ������X���J�%n:JE`ott��옘�L`l����-w��g��j��226�Fw���h�Gj����t׎3�8�#%���M���uM��=�n� ?kw�yֹ�!%�C[���N~I�b��ۑXz�%��N|+"���B(>�ٟ��גO{������X�ɒ9�ӧIBs/�`ott��옘�L`E"O��(�*St����7gE`ot�3��>F-�#�I9QR2�)���106���`l����#�m�m���u��5U��4.� W�%4�Uc��X� �Gu�ݫXMsi�^����ky̵w���oI���06H遽�1X\=�	$t���$�s�VguՁ������~�H��7�*4���Ӥ�V�u`f��꺻6�`4
	3k��!|GЉ��|HD8p�|>7�� >��0`G�}1� 7:K�ˣؐNq	�z%����xp��NvS�P��7q� �	>���#��m@��h�O
BV�)BH�C������@,���O���!B9l��0�"�,�B2��]�<O���1��$��|E��\��'���>� #TJ��z��DI ��Â��= ,?�����B�� }�{����y�w+Y���鶓�d�$�7gE��w�z}��:Q����� rw�
���c&܊�3;���߫^���n��V�Ί�+�z%"���$�)�Tãs�$��l�u�n�� �nrV:7a�`�����KE�d�~t��RP���{���o�����^����>���������-] ����orQ2=w�8��x,�w��_��QS��$�(�q���� ���Q3��� �}� ���P�O��H�rEa��_��������� ������ P�_B��,�I"~@X"��
����}��'��~�K']�)�������}_���D(O����O��� �Y��	'$�����9�$�EH'd�F���eI��N����l\=U��~�w%F�m'��H��{�V�m���7|�I~���Հl�]r�c���ܕ`nl�߿~��f�����Հ{��g�䒪�Y%]���"�j��p_�^���áL��b���V�F�r)N�N*r���Rׯ� ��ŀo���)����:{�k��D��JG`fw]X߿v��/�7}��j��2��r�	RI$�I$ ��m� ��l�    �
�:4���a���t�܃�H�S,�z���#�q�ێ'�'����t'4P%��Um�� sp���78r�#�u�A[UGh:�maݩ�(B�s�����铙3�Q%8����b�^ͥ�K�8��+��dz��㳭X�7�6u۷%:۫Į����;\�vm����Q�&�ͻ�m�v�f���l�� �cb�c���HM�t��U?8�����1	]9%)ERV��ﯮp�n�O��~��}� ݇6�H~���M���Ӌo;;z�����_�#+�� H��m�.������od���Ʈo��I��i�$���޺��K����O,�v"�_Sq��n1��ݬ}��p�����l���=��a��}����8�*�c�ƻ��nzN�;��p�hCFjX�θN���R���4N�nE`ft��ś���޺�76tV.Grd�S�ӊ�p�1f�s�A��=�Az��%���'������3�$��:x��J�*�+�K2�'�L�ɉ�������i�TRS�PE%X��vd���6tt����P�ڹU�-]�`����l�0;y�DDB录�w6�&f�����]IT����u�\�K�mԯl�W�fA�å��ᶙ��D��Fې�[�vv�Ձ��p�7:q`b����JF��H��0;z<� �ս-������lm��NIV������ř�q �j�DZ�F1F��� � A�
���y�{]���]X[�S��H)�Dۑ`�a�;:��w_�m��qɒH:8��7o;��Ł����7vq`{�/��FD�H���U�94�zw/6�ӓ���:�[K$f�TGF��T��7l����w��A�����N>D����w���A�666=�y�pA�666?g���|�����>�2Y/�n�B����A�A�A�A����|�������� �`�`�`��}���� � � � ���?N>A������L���wr�n����lllw��8 �����>A����߹�pA�666=������A�A�A�A��oY%�lݳww33vpA�666?g���|������s����lll{�y�o �`�`��Db�A!�s����;���pA�6667���g��\�wr�7w8 �~���� � � � �����>A�����?N>A���������A�A�A�A������I��b�#k���h�^�Ҧ����]m�9�������v���Wm�ܳɞg:wwg��A�A�A�A������� � � � ������ � � � ��w�pA�666>���ӂ�A�A�A�A�������n��n��ݼ|����{�~�|������g �`�`�`�����8 �������A�A�A�A��Y��&�e�6���l���lll~Ͽ~�>A����߹�pA�6 �A� �~���|�����߹�8 ������\�w3q�$�78 �~���� � � � ����|����{�~�|������ �{���|�����;,���i3HL��8 �������A�A�A�C� ���~��pA�666=��g �`�`�`�����8 ����F~��� ���km�k� ���    �νd��h�h+q�N6Ϩ,Og�R����|�:�2�Sn
�3�v���IrYГ�ĳL����n[e�����> ;Gn�-�j�b�TblQ��:WR�[X5�j�R묬-���fP-%�,�[ygsG[��]&�A�.��t�2�x�:�ٞ�q/Z+��k�Vg����w������??��j���To�m�
�V6��j�onn7b\�Rs��S�N��c���sYnn���666=����pA�666?g߿g �`�`�`�����8�������A�A�A�A��oY%�l7M������� � � � ��~��|������s����lll{����>A����{�ӂ�E�A�A�A����g��\�wm�n�pA�666?���ӂ�A�A�A�A�{��x �[��?N>A����������llQZ��~��N����H|���������\�w_���u�ДB���0O��u!#N�nE`v������U�^���=��,ݝ��r�dm��$8��٤�^ku[�X����[T8R��s�q=��{���T���q��:�6�������� ��w=�G�n����]*��ꬨ�A3wX ���j��^�B�1 ��h�
Ҁ�`�QH6�t �}�ό�͊�����ŝ��_�#���=IH�(��I`wt�Vn�,�%�}�`�zX��J�M3��E�+S����V ?7x���s�j���%DB�R�&�,Y��/o�>����;vq`nNQ�I$�F��w��-�	˰�g�Z��V�i�{v�7q��UZ����)�
�FӢH� ������_���C�=�<X�����}M�M����.�� �זgB������ r�����_�$mw�S��28��D���?w��rI����MC�(
������BJ5|�������vY�l�MsD���Ԋ�p��׾�o�,ݝ�����Ł�Ǔ�`�D�)��� �����ι�7|`�7Y������
.v�����nN�t�c5�k8��O4Gh��un͜0c��o���ӵs��*J%1�>����;vq`b��Т����ݢT�J��E����� �m��!(�6w�����ݷs�	L����(W%������6w������/�DDUwu�s�}� �K�`�mL���iwX
Q3��xn�� {��>JyDFBQ
�LBMD(����~���w�ʪ�UU�e�ww�n���"���ǀr��v,�v�j�q�) I$D�8��s۞obu��d�u�Ŵ���8�;\7g���V쫅H��N�nE��,X�`|�rJ���� �d�.��+�Wd�Y�z|�g�B��Q���`����3�%29㦺h&�R\����ӽՀn�9(�S<��n�yX ͦ3�2�jQEG#������%]�������=�np>��СDU|�����D�
��K������ {���J�""y�����^��,�0�s}
��Cp�F`Ed��c�F{�i7�R�J^�Cꄐ�KO��f�30Z��>�6>��p���BRt�漻�w��:��_  h m�         @      [@��@    �p   m�[@�            �\    	                        Yέm��^��y�UNԱ�o�eN�/nW��1�@�Ge�V8ެ��sٷV{v��n�:�k� kmƸ�B�[үA��`�����6v6Ij�� ��8ː�em�r�pep���*ʻ�&���I)����F�0[�s:����=�kPv�TV�:�4��㮫ɛM�%���X.�@M���0���u�L v�Oc+�m��uM�y�9\Y�]�7+غ�����҇��|���b�m��gaVK{bU��Z4��z%�ݮd3��K���0��3��=��M���t�m�<��0,q��6����nʲ�Y�)	��sɂ���A&�n:&�`5"�JlZ�r��NM�8��<�UPpڀ��r�V�yUj�P��Uj����UJ��Yf[;�Lgfcl�O��+@�U�@���iJ3���V���m��vX$ [�}���:�S���@P�UiV��c)p
���\�X�Y�N7;�����J���(^��m�`XHA���R��:�UU[���Ş�L���z�fm'<��e�v�>"�r&
����t/g	�1���B.�j�Pt�3�ԭ�Q����t;8x�m�]d�#�ngY`��W��9ݶ�ݛ�2�j�����k��>��qۅ�p�|G�gw|�H�"�s��Og�ob��͎���Jz�Ƃt�Cm�|p��ƥ��nY�g2���6Y���ZȐ	Q�E��;��
�e3����v5�1�kz呣;�Z�[�^`*XT���	UU�-�=��@B�(t����J�n�ڢn�N���u�l�a�ܛ��Q����^"�B.� 
�|"��z���(	�S�}�͓www@6� �ְݤ�  $    mbnd뷶qwI��f�O	��WG��p��O�C����xs����%lI��u�g�����;T
`���]�l,�
�"�$��<G:�+l��e'<$�^�[����E��J�;p�m�p�m�h,\9�7ۗV����Z�\τ�K��L��7�J[NgO\�e�a�l�n�<T�@9䜞y�RI$�Ӗr�����G�uٺ����� �K��q<�'�Lg�����O�`�Tr��U��߫� ��wm��I/��x��߂����F�E"��霒Jdm�\���z|�gDD)�d���n66ӌd$�X�=�۳�9%
gg{� ;{� ���.iW53h�����IB�o8�6w������ꪥ���Z�y27?6*�Q� ����9(IOou��}s�=�f~w���\�Q���띜qm2+��u�]KV�0�'Q��X�����m��V�9@���o�,ݝ�۳���(_D%�r����|���4�hEM��I>����r�j��@"DR�}��hU��������=;�X ���BJ"d�7jd����"�I��87|`�7XtDB�������R�7kH�T&��ۉ�T%;��8N�V�Sjp>�DD*���ŀ���
jRC�u�����脣u�L���0z��R_�\�M�v�n��̻����'=b!�-���6L3��q�Q��)���>n�?9eL�h��Lw���;vq`f>�ꪪ��������)C�mJ$�n�3�%&�wN v�^�k�3�B��ɾ�dnB�BAGu���;;�~HID$�r�J�o�������/׬�4�0͒����?�*�g�� o����0<�%��UϪ����z���%2I,݈�w�J'���u>� ~n��z�赶Cf���*u��AE��C��\W\�dǝڱM˅�6nm��D<撖L�smv�7w3�n��<�\��wТ��C������_�=����5?6�M�X��s�BS!��x�}3�=�ftUU~H<j�~
jR��S�������s8r�IL�w����/m5UuE*��76]��З�	*�߾��>���9$��og$�A=?��ê���������'����ɷI��2�6ʪ����0�DD|�?��ǀ>}x��J�+��H�1	�'�"D�'\g͟ҹ�G�v���<�0;u�$��������Y��dnB�������;;����s=	/���9���X*�V5f ?7yТdz�pn��<�ٝ
&OHkTQ+��HEwx�}3�=�f	L�;� ;{� ��D�
�N�b�I���J'��0�|`gt��R���Vuq�$	���⪻0=�`���_�����2I�������8�|l m� ��p�8    �z!s�j)�wfA���(]F���Q�Bq1c]r`�-��5�ݢN�ZE�����뭍���t�6vݮWf��v�T���a9�Zy��6�e%���l�H���7&���{B:��ۭ��6��6&��l���\������x^�vrԖ;s��g\����w����w���ӡ�`���$��a:�y��zRA;t����u:[vrh���ϙ>/͹.ԑ:q�@��������X�8�3�q`b+5�76�(�RG`nl�0'vA��t�[%��$J����`ܦԢA��=�<X�����yo��ޞJ��v��܄""�GJv��`<���ۙ��J{�q�r����))(���M�`r��`��	!D}����>��0O��g���'A�6٪��em�{X-y^`SV�c�:�t����X�V�:lO���|��cヨ�!U]��5����`�7\�!~A���3�t�R��L���X�ٞ��.��EQSϫ ��Հn��}
�|���Bd$�u2U�Wf ���p/]a�D�n�� �w� 3��*�SU3wSJ��p>��������V���N ��0=	G$�EO[��5��M�J�r�R�r;wg5`wnA���&S���!339�JTF�[Z瞑�ktgrgm�J�3�����ڦ�����yn����%ڰ�~m�������\�$����N�{�27?I�E�.�w��_�$zw����N �m��!L�x鮚�LݡU*�����{� ��u8b"D1�`H��!�S������b��>F-�!u	�	E������%-����0K�X�P��{� ��Ғq�I�Ձ۳�UGB�Ko�W��o� ��u8��t��nv�./OR��f놹y�U�-�L�_bÖv�v8I��u�X�;�������� ������yBP�Hsw� x���Ҕ��i��v,�w��_��F��N�����%脒����ڃtӔ��I��z5`v���
&vy�`;�X�kX]�SV���vMU��rP�y�� ��Հ9�u�L,NJ:!E�v���:M|QuWE�Y�����t�[%�;�%��Xˎ]�"D� ��)(�<I��r��Ŵ`�2�k��Nv�ZH�]�#�����;��pBp*:pq`˿��������(_�7����e�$�E�\U�Swu�n��3�D%2sw��O� w��9�����>{�IK$���v�ٵWF�u�`u�p�
S=;�Xo��v���FTi8'!a������s�����7u�ݶ`=.��aTU4��� ~n�J!&�~����z^��-$�ע�/wZ@ �m���.��  $    I{i74�T���M�/ѯ��:l*N�i8N��4��C��Ѫ^��5�t˅���a��1�6Iٜ9`f���]�G]X�Zm]n���e��d).,a�
�:H�f�(�l��]�r,8-�.y�%im�Z%�!ƬX.��]�:Z[=��MD��l�����w��x�*��i��iGN�6��{v}
A�N�<;{q������������~r�9sq����vQ�=�f�z�BK��ޖV���ԂjQ ��X�8�(���g�V v�^��q`#�QuSpU�YvM՘�� o]�СD�wy]X�O�9>l��E'Nuu�В���׀6�q`���D}�;���ds�)>T\��X�7wX�ŀrQ�q��}X�7X�G��������`�.v�w��� ��	.��f��x�j<���,��uQ�K�x1��Ӕ̗wu^����=/]`|�"~��}����z$%IJ�A�'!`bﻜ�@à#"�SZB�5Q� ��P?��f��g ���U�=�ft(�6z���WU37U4����{� ݭuX}	|�U_w_Ł������Vk�mF鶥(�RG`nֺ���0:�8�������K����\�-WU�=�f�!F�w��yo��׼݁�r�dm����enfN22K.�v�B�2<�k դ������{��|�gKyn�j�M�0l������7k]W$�~����y'��M�?9Nn;�o;u�:��f�z�>�_$�*��}E�*�B��������a�U�&2T�:t��F}��>��-@B�B0� D�HI`1C  ���@������&b��A��}�#**Ȃ���� ��� �G�1�=\��I�$>T5C���>(�(²�� Lg> �
��)R��-�ܰ�C�H��Lۘ��6RRf�Ü\�������l��({�}�"��z'}ؐ�.�
��'�� ���t=:
x	���/����q�!Ǌ���Q"��q�B�Q�s��K��{m�2�E$�$n��K���`j�y�v��7^�vmi:$%IJ�:j	�X�����ϫ�����`�w�X�t�s��rr�j�Ű��M�����J���n�n�MZ����~l�QZG����}W��~�}U�7�BJ>�_��v"����Q�6�F�$���{�Xz�`����w�
dki��4Ԣ)D�8݁�w��]����{�,��n��v��M�c�T��:'y������U�J~��(� �X�b�H���{��'˵'Ҥj~r��,Y��~���o�=��;g�ޥ;�)�!:W�����nN�t�e�B�GH�`�a�#���$I��ߣ	ʶQ��E)#�=����X��:?H�׀z5�%Hy!8*IH݁۽u`gl��;;������U$wW�!*JTq�PM��7��9�u�BS-����X�.o��Sm)tㅇ������}����o;Y�����B9%�����=^������vݿ�����~�?��i  m� i�a���l    6�l����ǰ�v��x̂n'�����c�f�[]��v;jN�n.��0���6����9���ͷ�w�����l�T�<�R;;1Ŷ�mkp5��2�5�p]T��Y����i������I���XgB�k]\��8��쫮�k��$�h,9���x<��GVxᨑ+����'���Y-�;$*9��7�ulu��v��v�lN6�9��z�Y3��:���au2"�J#����V.�vݽ,׼݁��ᒛ���T$��]�Y�L�s����Xz�d�	r���~��'$u &�<��v��oJg��,g�V�C�E	Ю��B���v��`�ŀz^������`g��I<�u#������V�_���;ϼ�׼݁�0�q� �J9g+�q?���s���n�t�ptX7$�X,�;�v�2�sA����X[�6߿��N����u_$�H>}� 8�ꮓ%�2eݛ����w�wy©�(�	.�����X��,�v��,�ͤ ��c$�X�y��z�Ͻ��7����=���2��R$MH�ISh����(��ߕ��� �mX8�Էf�v��ᒛ���T$���78��X���`���?�˭��E�0��q\��-�L�d�5�ۛ�H�ۣ[S�.�ctDU���a�ܕ���`M�����pmk���gB����+o1��q��9�����:vA��r&��?�|��I���/�U]"�����;��{���1
DW�U���+������tHJ�iʦ�W�07nD�$���i�'GL�\��Ƥ#��Vݽ,�ȓN���"`{K]1x]X j��f�<<r7dvԜ�����J�a�5���\�8�!Q�M�DN�C$�����0$�遻r&Ӧ06��R3奉fR�K1&N���"`:c3g%`b7xd����	$�3�0����뾙�5�ŀkw4�[�nF�@#��woK3g%`wo]Xg����Ł��2��Ԏ�(C���&�07fA�I��~��[d6j�z44.�B)�R�n^���m\�j����\mX�ͦ5�x1�l�� o^,�m� ޻�P�����z�����!J�
	�Vv�/�Jd>��}S�k׋:""�v�o���HE$N��X{�,ݜ��GLۑ05�r�������$�n�j��޺�3r��%��Kk_z�%'$�)B��{z���B[��?�>�۶�p�x�I~;������;����D� 6� �ְ�I&�8 �    ;5�G&Ʈcv�Y�ۥj�<�x�6�ы���<m�r-������W`֍���^Nl���iz�v���:^P'\m�RR�G�Lm�]1l�� �U��@�Pl��7������Πs�i�%���ڼ�[�1�VM�ɣ��ogG���I�3f�]�I����7[�jj�w��=�������8ˢ�|�0��x�x����8�l��c�l7.�nqY�-��E�AI+@�����zX�9��z���|�G(�:��8��f07�%��07nD���,��rF8P��X�9�{z���}�����%��K?oJ�/1��47#�^�X�M� k�x�N��S�o���~�B�ܫ1�+ ����i�ӣ���b2�WV	&�B�]'@�u�jn%�e	ٺ�Ǣ8ps:[ �����Ȉ�')�JF�E"���`{v�N�^.���!�]Ӏl�]r���)]L�E���ݷS��J.�{�V����woK�)#k_z�# �jmL���ϱ`�a�(S's��7�y���%7)�QPpRJ������ }�}x�۩��S����WK�r���)�i��7�������7����X�wE% $����u��뜼AMb�n��;�cP�<C��ݮtؒ6"�ʒA�����X�06_D�:t�����)��e��2��GL��0�1���-Xդ�~�B�ܫo; ׮��#�B�BrW}�yS�v�ʰÛ�br�����vݽ,��i�'GLS��5�r���.�]��/3ݒ�N���K`���pgt �RI?H5#D�J��<��vv��.�4D�S�v�.�#{t�8��N�k3�,�L	::`j�-�I�?}��<Ձ��xd��1� क`b�u������p^��Q2>���r���Ӏ���;��`n���G{�,��+�b�"�ߤ���D��>R�Ω��׀yֹ�Ԣ҅	�쪻w�,��(BВ'Q������z�O��׀n���u���`����)�{P�U'+��ev��ʡ����]���uͅ�G&,���OJ\�`j�-�I�ݒ� ��0	�7���� �G"���~H���8 ����7Y򈄦M�k�UR���F!�I,�j�7����;��ooK+�"FA���9���`b��`����ou��Q�ᒛ��(��)%��;��ooK3g%rI�~��I�� }�*��(���@Vئ`��D��D�!@�PH! H @H�H��"I���B�CQ���(R�HR��A� ��B̡HFIJ�Y� O�+,X6ZJ�R���a�i�'�P秿}}zOow�>�w{�ӷ����  ���                -�  $ �  	    n�m�            	��    [@                       1<[�p��l�gix��u.��ۍ�.�u��l0l�)�`���s��3gj�K���A�YL��l`���.��	����W.�*�6��eٞ�f�0���r�7��v;x0���+G �e6�b��T
i��^^��������F�u�h�u�ǶL#�m���I�z���)L�R�X 
�we��Z��mel\�;	�n��e,�=�����;�5�\i�w��;R��:ۃi^b�����hr���q���;v���c�^h�ƽD��9^�s1���l\�[��ų<;����r�/(n`d��!^�* �u+%�)%ΉU���)Z��t�+�� �Nɹh�mi����*�[��n$kn��l� ��
��Z���@��Vqۊ�e��e�
�`+��qU.X5v�; ��1�Z,@F�N�(M����%A���v�j�t ��J�U[�.
j,v�C�/�S�2vI�[Hy-֓&0@2�
A�j���E*@&�S:�sp��Gh�<��qdu��M�{��S�e�<��ٍ��M����8�'��ݫY���ûk��P;D[F24݌��VF��t��i��[[%R�'�87H&�����ʇ�܋R�0/I����S=D{g���#��Cj��*.[�����q��Gb�;����M���@�3�{A�Nܜ[�=���V������{N˖���v+�l��Z�q��R�ܽ�RR��E7=O���*�Os�Ɍ���.U����*��;����M-�s���A���Q��P��E�N�����}�OE��x���w��4����� m��l /i� ��p    �鵵,��IU�:p�<���x����u�E�6�.%��V��Ǎ]�W�Է*�a{���c���4�8u�D��I�\	ũP�Jg1-�*;���C��_����9�"��%�gV���ء+"\�A���k�yㇶ��n�N�c��Me��@�J�r���Y�K,��q��'A�6٪5�Ɗ��zx^�hq\��q����T�k��s&5ک8�r2R�QӀ�����`fl�^��(_�6w��I��f	虻*���`n�D��1��d�'LΈ��2z5ڙ���.�ԓWs8��cV�lN����07�����N?9%��;��woK3g*V�IwoO�I#���18�)�7JH�I$�t�y$�H��K�$��?g��Z�A� ~�����i�����f�;Y�:T��WC���\Rr����5�8l�q���5I�1RI��%�'*V�IooO�I,O�?~����I.�z}�Ius��H��2TR��R��K{z}��USmb}��I%ٽ>�$���J�Ic;xdc��(��3=��r+i$��3�I.��t�I%ݽ>�$��'q���E�)������=��Iu�K��I):g��Z�D�$��ŬE%ߒ�QP��}�Ik��I��]:g��Z�Em$���=䒕�?J.v�ss�3�g��4gd�%��fϔ��)g��U�m/��75���WI��]:g��Z�Em$���?}��}U����<| ?���c�gؙ���X�rwꪯ�M��{�>�$��^��[���H�s|Q	�(7JH���]:g��]}�	��_]���=��r+��X��}M��#$�|�Z�.I��]:c�Ij���K�L��K��:�#�2TR���[���K譤�]:g��]}�	���D�,�.�q��W؎�c���[ �ìB� n��V���d5s�6t�77k7b���Kn�i$��3�I.���I):g��[ϓ�S�J6�@��I%ݽ>�$��I$���Imܗm$����"����4�MI>�$��\+I$����/W�޷�7i$�{�>�$���BAȎT��
�^��_�6�����%���ڶ��~��嶾ʪ5�L��B���Pa
�:���n��^[m���B/C�9>�$����$��ޟ|�Z�.��[���KXt��(<�E$D�F΋SGT�Y�.��Z:�;;۬w��էcKm�/gO� �����K^�´�K{z}�K�\����Z�~��I3�E�U~~ ~��� Ӧ{�%��V�I.�3�I%��r��`�d��(+I$����$�'ܝ��[���K^�´�X����� 򅙞�Ij���K�L��K��A4�K{z}�Io>N�FB(�7NN'i$�N��$�꯫��/$�S����Ijߟ�}m�{ޝ���{���Ā .���km�k� � @    j �"8��P��s�p�b�6*�-��,��1�;���N^8�;�ţvz��{�)�fK3V��ٖ�	�[WJ�[,Zc�3%��gs�nn�U@6�:J����-��ᩕ�C1��:��9-l��p=�#���:4�m͝�5�n�]����]��7jJq��S�v�\d�ͮ{^M�1˃�:�Cr`7D����z{tS�+�Q��A5BjI��]�p�$�ߩ�>�O<��3*dOs{ۜO"fTș�3��v'�Tș�2'���['M�n��]ݗ��Lʙ2�}����ʙ2�D�7����&eL��S>�wby�L��S"}���<����ؙ�>�����c�������{��S��q���&eL��S>�wby�L�+��>�{59ı,�s�G�,KĿ_�r�,̳359ı;�=��r'�Tș�2'�o;/��Mڙ2�w��jy�L��S"_���O"fT��S���?_����4�w���w�2�D���e�y2�D̩���ڞyS"fTȗ��n�<��S"fT�~��O<��3*dO~����͚d�����M�Q�]����<���<mp���j!�lW`�K�n�,��3.�L��x�D̩�3*{�3���Tș�2%�{ۼO"fTș�=߻��*dLʙ﷝���LʙOw�~�s�unn�l�����r�ȗ��n�<��ڛ2���w"y�L��S"w{��x�D̩�3*{�3���T� �Mڙ�����˻$�4�7m��x�D̩�3*}����*dLʙ�����<��X�C"fT��gmO<��3*dK���x�D̩�3*����]�X��fw����;ܧ��bw������Lʙ2���~�<�D̩�/����y2�D̩���ȞyS"fTȞ��	l�����-��v^'�3*dLʞ����2'�7q6�>�߮�<��S"fT�{�r'�Tș�2'��/e�y2�D̩ݒ��f��I%�����;��}�:���t�l��+7:ܖcAy穌�Ā�7v$f*{�L��S"_���O"fTș�=߻��*dLʙ�����<��S"fT��gmO<��3*dKݝ��\�۷7r䛻w��Lʙ2���w"y�?�c�7jdN�����y2�D̩�y����ڛ2�D�o��x�D̩��;��߯�)g�kQ#N�~~�{���>������Lʙ2��s;jy�L�ʈ��FHV~Z�CO}��K��˼O"fTș�;������;ܧ�����~?x�쳮��ּO"fTș�=���S�*dLʙ����'�3*dLʞ��܉�2&eJ!n�����U0��U0��L���f��ٗv��ʙ2�D��{w��Lʙ2���w"y�L��S"}�9;/ș�2&eO~�v��ʙ2�Dû��
.q��������;v筦L������l�o7̜^�u�$�\�
�N��[�nm�'�3*dLʞ�{��*dLʙ���x�D̩�3*}�3���Tș�2%�{ۼO"fTș�=�/�20��Y���w"y�L�r�D����O"fTș�>���S�*dLʙ����'�3*dLʞ�{��*dLʙ�~�-��\ݺe��͗��Lʙ2��s;jy�L��S"_w����&eL��S��w"y�L��S"}�9;/ș�2&eN��e,�\Зr��ڞyS"fTȗ��n�<��S"fT�{�ȞyS"fTȟ}�N���&eL��B@H*��a	A�>��}ߟ����=��m�~���CH�[w��Lʙ2����D�ʙ2�C���'�x��̩�3*w��֧�Tș�2%�{ۼO"fTș�=�o��7,�SYHh�s۩�(B�{"=��I|��^ɘ'�([��K<�Z�*w��*dLʙﷇe�y2�D̩���ڞyS"fTȗ��n�<��S"fT�{�ȞyS"fTș��3���&f��n��l�O"fTș�;jr%�bX�{���yı,Os�܉Ȗ%�b{�xvq<�bX�'rw;2nm!��.l˛br%�bX�����yı,Os�܉Ȗ%�b{�xvq<�bX�'�ov��Kı>���snf��3M�vۛx�D�,�"}��nD�Kı>��Ӊ�Kı>�{�'"X��S� ]���~�x�D�,K�-�����74�i6�m��Kı=�N��<�bX�'�ov��Kı=�{���%�bX���n'"X�%����F(1T�D߰�@ l �kXom�  $  UUT���,���n�ÍG������^^`�m[��Ɩ�[�m�D �L[��6涤;v����6�չ���m�ۘ�8�-�:ٌtDd����
�� K�%˚�O3���sʋMפ�+oHA���br77$�K���kfu�ڍ�7C�X����WE�mH�ι�\()�C;w��D�[m�*�v�Z՗�ui7/ p�@�U�K�y��]e�����m(�r�y�����7���{�~��Ȗ%�by�����Kı=���ND�,K�t����Kı;��l�Yt�K�swlND�,K�w��O"X�%�����r%�bX���ݼO"X�%���ݱ9ı,O:v�\�ݗ6e�7v�<�bX�'�;ۉȖ%�b{�v�<�bX�'�ov��Kı<�{���%�bX6��3.�0�ٛv��Ȝ��DȖ'�i�׉�Kı;��֧"X�%����'�,K��;�Ȝ�bX�%�����ܙsl�n�M���%�bX�}��S�,K����oȖ%�b{���ND�,K�w����K=���v�?~�8�U���ãl��0OK���8C�3rq��vz.�6[�ˢ+��t�CsH\ٗv��Kı=�{���%�bX��{��,K������yı,O���Ȗ%�bw;��͹�\�ܻ�nm�yı,Os�܉�z(��Bg3�S�"y��w���%�bX�}��S�,K�������Kı=�[��L�&i�i7.�D�Kı<�N��<�bX�'�nv��Kı=�~��yı,Os�܉Ȗ%�bx�%�v���ܙ-�v�<�bX�'�nv��Kı=�~��yı,Os�܉Ȗ%�by�v�<�bX�'~�N�%ۗa.��͵9ı,O=߻x�D�,K�~܉�Kı=�N��O"X�%��۝�9ı,OʧO��~��n�U�z�I�=��DH�N鶞x�&1��l:���%9rt�p�ȺA^���bX�'����ND�,K�t����Kı>�s���y"X�'�o^'�,K�����̴ۅܙ�m�܉Ȗ%�by�v�<�bX�'�ov��Kı<�~��yı,Os�܉Ȗ%�b_O{�,�ɗ6�6�Jf�'�,K����ڜ�bX�'��ݼO"X�	���Hy�+�a�i�8�S�����t32d�(0	��*�o
R �����a�2�s$�`��0H,J1�bbS(K(KX+b9¡BGA�
8������(� j'2[�0+Q_ra.yi���h�2]F�GD��4<"��b�CDz�QA)�SŘ���N��=�r'"X�%���}���%�bX����ɹ�&搹�.�Ȗ%�by�����%�bX��{��,K���>��yı,O���Ȗ%�bw;�n���w.��6ۛx�D�,K��w"r%�bX�{�ݼO"X�%��۝�9ı,O=߻x�D�,K췽۹6٥�F�����h�r��$���',I��75�zS��b5���g0�g{�oq��K�t�oȖ%�b{��mND�,K�w��'�,K��;�Ȝ�bX�'�{��d�˗wl�nl���%�bX�}��S���1ș�������%�bX�g�ۑ9ı,O=���'�,K���	�#w.f�]˛�jr%�bX���v�<�bX�'��w"r%�bX�{���O"X�%���ݱ9ı,O~;y�C.n�6m�7v�<�bX�'���D�Kı<�N��<�bX�'�nv��K��y@_�`UT͉�o;x�D�,K�߳�e��.�]�n��ND�,K�t����Kı>�s��"X�%���oȖ%�b{���ND�,K��oߟ`��1Uu�BRk�-���I�vv6ќ��q��r�k�	�.ݗ4�MƧe�tnJf�'�,K����ڜ�bX�'��ݼO"X�%��w��9ı,O=���'�,K��N�fM�,��K7e���"X�%���oȖ%�b{���ND�,K�t����Kı>�s��"~Dr�D�?g�����neܻ��nm�yı,O���"r%�bX�{�ݼO"X�%���ݱ9ı,O=߻x~��2%�b}�����n��Ͷ�3sr'"X�%���w��yı,O~��Ȗ%�by�����%�bX���܉Ȗ%�bx�-�N�̻�fKpͼO"X�%���ݱ9ı,O=߻x�D�,K��w"r%�bX�{��8�D�,K��l(0b\�:�P��7�l� 6���i�a{N� �    u���؜���X�I����^z�|V��8����Tێ1��>�ڱJr�%��n�z0�Yĕ4�Z6�k���M�P��� �^;�6KٓƩ��r��fU��"'m\"*�R�Gj}��ú�v�g+�۞�Y9�Җl��7.y�0c]ywFڍ#/Z�Z�uq��w�;�}J�%�qzz���-�@�Ϙ0���l���Qq��MF֬&a�s6�\��ؖ%�b}�����Kı=��r'"X�%���Ӂ�P��Ȗ%����9ı,O�~��e�˙�m�&��'�,K��;�Ȝ�bX�'��{N'�,K����؜�bX�'��ݼO"X�%�a���2�]�s.ͷwr'"X�%���Ӊ�Kı>�{�'"X�E!�2'�o^'�,K��?~܉Ȗ%��dL���~,��37&�w%ݧȖ%�bw��lND�,K�w��'�,K��;�Ȝ�bX�'��ݧȖ%�bw's�&�m�&M�nm�Ȗ%�by�����%�bX~�����O"X�%�����q<�bX�'�ov��Kı<���w&�4�I�\]�6�χ��ӌ��>�!�([r���a9�ƻU'b��Q��0|�~oq���=ϻ��,K����vq<�bX�'�ov����"dK�������%�bX�d-��a��4Ͷ�r��ND�,K�w����>+��B��R,������C��n ����K��v��Kı>�~��yı,O~��Ȗ%�bx�-�N�L��f�s6�O"X�%���ݱ9ı,O=߻x�D�,K߷�br%�bX�{�v�O"X�%���'p�ܹ�w37v��K��"{�;��<�bX�'���br%�bX�{�v�O"X�%���ݱ9ı,O>;y�L�s.\�m�7v�<�bX�'�ov��Kı<�{�q<�bX�'�ov��Kı=�~��yı,O�'y�sg�b�.:���q!��sɡ�r&��ӭ��n��1 ҍ��ܡض��-�"X�%���Ӊ�Kı=�{�'"X�%���oȖ%�b{��lND�,K�{��f�I��4۹.�8�D�,K߷�br%�bX���v�<�bX�'�ov��Kı<�{�q<�bX�'r}��74�ni2n�slND�,K�w��'�,K����؜�c���1�M��=�{�8�D�,K߷�br%�bX���۷s72�]7\�nm�yı,O~��Ȗ%�by����yı,O~��Ȗ%�b{�����%�bX��-���]�wl�M�ͱ9ı,O=���O"X�%����~�Ȗ%�b}����yı,O~��Ȗ%�c߽�__�; �:�6+m�θ�/�ѹ8\�L����WY��4ek��ci�H�e��Oؖ%�b}���'"X�%���oȖ%�b{��lND�,K�w�Ӊ�Kı;݄�I�su�s3wlND�,K�w��'�,K����؜�bX�'��ݧȖ%�b{��lND�,Kώ�v%�0����7v�<�bX�'�ov��Kı<�~�8�D�,K߷�br%�bX�{�v�<�bX����7w,�$ݙ�nn�Ȗ%�H'��ݧȖ%�b}��lND�,K�w��'�,K���#H��(��,��AB�"5J̉{�l�Ȗ%�b_O{�,ۤ��4˹.m8�D�,Kﻜ�Ȗ%�by�����%�bX��{�'"X�%���i��%�bX�������E��j��t�n��.��`V�[d�iRi]��N���`�6tޖ��v'�,K�������%�bX��{�'"X�%���i��y"X�'�w9�,K��{�ݻw3rK�5ݶ��'�,K���ݱ9ı,O=���O"X�%����D�Kı=�~��y+h�'���L�2d&e��$�y�w���	"y��;�;�w��'�,K����؜�bX�'�{�R��33rٲ�ݧȖ%�b{�s�9ı,O}߻x�D�,K߷�br%�bX�{��8�D�,K�w�m�ܹ�Yv�flND�,K�w��'�,K����؜�bX�'��{N'�,K����!���2%�c�N��ӿ����~�p (�A����Ӷ� �    T�_&��N��g' ޲��g]��΂��i����ngcN�9����M��nj�wV�2�m��n�s�`�7YV�g���mc�,[3��qT�@tYf���ʲ�j&�ª��vAy̯@f��uϵm�-�Xk���΋�5�x�ch ���rp��j���.������d�cI�PyΊI����]����ƶl�ݦ�螜�l�i�s�r��v:�n]�woؖ%�bw���'"X�%���Ӊ�Kı=�{�'"X�%���oȖ%�`����wr�rMٛv�n؜�bX�'��{N'�,K����؜�bX�'��ݼO"X�%���ݱ9ı,K��s��t�7&�w%ݧȖ%�b{��lND�,K�w��'�,K����dND�,K�w�Ӊ�Kı;���ɹ��C7f\��,K?"�������%�bX�w�6D�Kı<�~�8�D�,K߷�br%�bX����nə�L�5Ͷ��'�,K����dND�,K�w�Ӊ�Kı=�{�'"X�%���oȖ%�bt�s�\�S����;^]��s�p='N�`V��k`���L�;v��Vd�����,K������yı,O~��Ȗ%�by�����%�bX���l�Ȗ%�bx�%,��L��6[���yı,O~���` � v&ı=�����Kı=����,K����i��%�bX���l.˛�K�3wlND�,K�w��'�,K����dND�,K�w��Ȗ%�b{��lND�,Kߎ�v%�7v]�rMݼO"X�%����Ȝ�bX�'��{N'�,K����؜�bX�'��ݼO"X�%�g�gM��K�nL۷7vD�Kı<�{�q<�bX�'�ov��Kı=�~��yı,O~��Ȗ%�b~�����.6�l9�sv�ܰ(SZG���3�����1�����a�w%ݧ��Kı;���'"X�%���oȖ%�b{�����L�bX����S��Kı?d�~�76ͷ4��并'"X�%���oȖ'�*dO�o�9ı,O~�ߩ��%�bX�}���,K��w����m�&������%�bX��{�'"X�%���Ӊ�K=�� Ƥ@	#?�7]<xybo7�؜�bX�'��^'�,K��!/K�Ziwe�M�ͱ9ĳ�2'�s��q<�bX�'{����Kı=�~��yı,O{���,K���zZY;�n��m��q<�bX�'�ov��Kı<�~��yı,O{���,K������yĳ�ow�c��u���W=���u���u�̶��f����\�Ggn��c.� n42l�nn�Ȗ%�by�����%�bX��{�'"X�%���i��%�bX�}���,K��㷝��sMݗvܓwoȖ%�b{��dNC�"R"�"dK߷����%�bX�����,K�������O��2{��?M��t��=Y�j���{��2X����N'�,K����؜�bX�'��{x�D�,K���"r%�bX�d=�t�n����f���q<�bX�'�ov��Kı<�{���%�bX�����,K`¢W�Kȟ}�;N'�,K��O��&�ٶ��ܷ6��Kı<�{���%�bX�����,K������yı,O���Ȗ%�bS�~�۱s�5F�۵Vv9ۓh�&��Ͷ�yڤ3�pY8v����GM�n`�yı,O{�l�Ȗ%�b{���q<�bX�'�ov��Kı<�{���%�bX��%�{KM.�I�wdND�,K�w�Ӊ�Kı>�{�'"X�%���s���Kı=�y�'"X�%������w2�n�m���yı,O���Ȗ%�by����yı,O{�l�Ȗ%�by���8�D�,K�w�m����e�swlND�,�	Ͼ�gȖ%�b{��dND�,KϾ�a��%�bX�}���,K���;y�L���ffMٗvq<�bX�'��6D�Kı<��vO"X�%���ݱ9ı,O>���O"X�%��ω���O�O���9�4 ��A7Q�O�9��@O8��B��)��*������e���|��M&�BBB�^h�)V��b���]�a��<Q�j��Ȣz�0	aXB
���N)���B!$H$����HyWSz_��	�\����1�X�|M/��{������  -�m          x      �    �  ��   ݰ�`$            �    �                       S�Q�6���`痗�,Y [!�=O;�ci�kD�Ʉw%K�/ec��(������ )v�s�i
ڪ�컴nΦ�R죝�hV�
٭t�-ɰnۇ�}uk/m���;f��#F�lnp9�<�Am��W ��{74X�cj�s��0�q��ur��wa�=�aK�(�M�]!4�-�q�^պY80Aٺ�nu�h�Oj��<]+�(q���Z�4n�wk�3����ؠ�n�]��ɹ�vml����T��]`y�l��pk�̅u��6Γ�$��5,�דSq���v�NX1��v���<iP˴��6����Ԫ��+,��;�m�FZUH��B��4����<�v��'�����@����[@ �]n�Y� �@Us�N��4Z퉑��,�j�y�pD��T�Q�Z��f1��&T���F�ړ#)<�mUU*��72U� � eA@���9�vPXq��@��@��:�R��E���<�c7:��08���Ix�U@*��'EUR��˞nb�XT0γ��v����F�\7���.�۞�h���=��{t����>f���N�ѱ���ҼrNw8ĴN�1;�3u�Y���ۗ��h�c���[v�mSƙ3�VjB��^8�c�<�m@/3�W�\����`ӷ�Mc���؛i���]h�pq@��U	�q��N�WCPUvSG9�7��:�t3��q)��f�c��X{)�ls&�� W����/����&ŉ�U���q�����e3�+���b�a�<�ummゝ�5dj�]�@�PC�?!�׽�uC�� Ph�C��U���w�����w�����@ l &�ۚ��`8��     %ŵ�ݶ!�"�iӭ���]�ݺ���Yc���m�⓵u�w]V���b�g�z�WG���Y��؋Kd�[9�^]��� �8���j�	ƙ��vbp��c�g�`Z^��d�oC��5Շ`�b��g1]\k���/d�-��v�{I��I\���w�E�4��`����磦��]��XBԯ@�'Zk��v�v.]F����ɛv��ȝ�bX�'{�;'�,K����؜�bX�'�}���{"X�'߷�؜�bX�'r~�śt�7&�7%͇Ȗ%�b}��lND�,KϾ�gȖ%�b{��؜�bX�'�oݧȖ%�bw'�ٓsl�sHnn[�br%�bX�}�;8�D�,K��v��Kı<�~�8�D�,Kﷻbr%�bX����nn���w6�6�f�'�,K����Ȝ�bX�'�oݧȖ%�b}��lND�,KϾ�gȖ%�b{����.�.�I�wdND�,KϷ�Ӊ�Kİ�(1�y�lO"X�%��{�Ӊ�Kı=�y�'"X�~�~�Uw�/z(Ȕ �$��r�Ɨte:M��yc.��eE9��ma�u2��������7-��Oؖ%�bw��lND�,KϾ�gȖ%�b{��d��&D�,O{��N'�,K�����m�I.k�幻�'"X�%���s���: ���blK�w�"r%�bX���v�O"X�%���ݱ9ı,O>����e���ndܙwgȖ%�bw�ݱ9ı,O>߻N'�,K��w�br%�bX�}�;8�D�,K�gs���ن�ͻ�wr'"X�%����i��%�bX���lND�,KϾ�gȖ%�bw;�Ȝ�bX�'�{�,ۤ��4��.l8�D�,K���Ȗ%�a�����{ı,N�{��,K����q<��{��7�����R�j��z�v�g��W������b ����3�2�悺�gnn�v�sr���,K������%�bX���r'"X�%���s��~ '�2%�b~�����Kı??����l��b[|�~oq������v��Kı<��vO"X�%���v��Kı<��vq<�bX�'�zN���˴�3v��Kı<��vO"X�%���v��K!��> Hr'"}�s���%�bX��{��,K���zZӹ�w7M�ۛ'�,K?"	"~���br%�bX����8�D�,K���D�Kı<�~�8�D�,K޻ܴ��\�%�swlND�,KϾ�gȖ%�bw;�Ȝ�bX�'�oݧȖ%�bw�ݱ9ı,O���w&�4��	3Í�k�k�����8�[�f�u:�Y�+d��(ܫ�%o����,K���D�Kı<�~�8�D�,K���Ȗ%�by����y7���w���_�%��:�*w���bX�'�oݧ�~T�L�b~�����Kı=�y�q<�bX�'s�܉Ȗ%�b}����ͺK��I��3i��%�bX���lND�,KϾ�gȖ%�bw;�Ȝ�bX�'�oݧȖ%�b{���͹��L��2�؜�bX�'�}��'�,K��;۩Ȗ%�by���q<�bXB"�ȝ�;�'"X�%���{Mͺfl��,ͻ����Kİ{����Kı<�~�8�D�,K���Ȗ%�by����yı,N����k��j�z�L�1�h�r�F�n�7[��g�lv+�֘�m&��Yg�����bX�'�}�É�Kı;��؜�bX�'�}��'�,K��w�S�,K���zZӹ�w7M�[�'�,K��w�br%�bX�w�vq<�bX�s����bX�'���É�Kı=��Kl&��%�swlND�,K�{��'�,K��w�S�,K��߹�q<�bX�'{���,K��v�L�.iw2nɛ���Kİ{����Kı=��vO"X�%���v��Kı<����yı,�Λ�d�&�ݺ[�u9ı,O}߻N'�,K��w�br%�bX�{�vq<�bX�s����{��Y����??$H m� [Mk��l�     
�m�.�3�u��M�L����&�*��rX�v,��#=�N�u�QŰ$�����;�N��'���4�[��u�R��p�6L��B'ʴE�N����U�u��7��	�m1Ͷw�E�x婶���㞎��γϻ=[����GS����~|�����qK.Ig��}&�婺�(<Hڂ7��]��s��<	ճi��&Nz�ƻb��&�m��j�.nM&i��N'�,K���m�Ȗ%�by�y���%�bX=���r%�bX���v�O"X�%��O��v���!��nm�Ȗ%�by�y���%�bX=���r%�bX���v�O"X�%���v��O�ʙ��~��Y���n3���{��7������Ȗ%�b{���q<�c�$2&D��v��Kı<����yı,OrK�;	�n�������S�,K������yȄr&D�?~��br%�bX�����Ȗ%�`�;۩Ȗ%�bx��-i�˻���.fӉ�Kı;��؜�bX�'����O"I
HR(t���z���9D$����n.v�.�ũM��r�Tnzє���Y0��
]�G�暎�xP�7M=��Q��{�~�"`n�B���0=,`T�Uj���
�0Λ�~�~D(����	B��6ne�`�s�~�N,�#�Tj�R)IH�͕���&�d�"`j+e�F,�^Y�^U����0=� ���3eq`|��$T㔩£�N+���L�ʃz�&��^�\m�U�=q�C�9����7 ���^s��)�S�=]C^�����γ-d���L�ʃz�&�d�yQ�F�t�����`f��`}�8�>�ܬ�c�J�sjG%$���{k\������Bp���؅	BB����+�u�`�+jeLȝ]�»������-��w����}��r�T7(���H���+w����}�d��2,�ˤ!eT�Y��5�bÝ��i�j6�<:�:���ƽg����Dr�P:��JJE`fo_���&��lK�05��#P�,ʵ�wxS��'�H6K�=.D����h�t�S�R�
�4�V,�v�Ș���u�LS�����eD�B��s�Vf�*��{��?"8�9��{��{d��vv�7s7	1^��S��&��lI�`~���~�\�U�]3��:�>~X�ø\�d��$�6-��g�6�'��q��T�W�x	.~L-���!�U}��A���Xߟ4*A^r?�m9"�>Y��� ���0;��`z�Y �QH葑�H���f�*��{���gs�>X�}Q���Ԅ�R��d)��}�d���05��")Cq�
Rn`n��g�,[�;=����޿�k�	RI$�I$�I �h6� �v�8 �    6޸m�˶݇\q��M�k�$�E��\5y�S���9'X�c�{o���ɾ�ڮڦ�pH�<o�cKv���&[�8��umgA-�;�еC�^����l�P�$�-��n���.���&�7,�a�/<tݧ����ݍ'*����7�k�X+2�Mm܊|��3f�n��˓K$�Uã[�u���n�H�j�a�DP���v�i��!�Ȫ8�q`��v����#�G����y��WUp����v�Ӌ3z�X�yX,�v �GH�$n:�VoG���&��lK�0=�ܤ��Y���RK3�u�L-���"�37�����zЩs��i����-��r&�G���& �^$������մgN��/J41�b�,'E�u�wZn����E�&���h�M����Lޏ�u�L-��Z�r�)����v�v�I�w�5 � 1`�� �H��/��9;����s�V"��R �!�JO3�u�L-���"`n�B�Fw&G)B*�4�V�߿RǾ�3��Vf�*��{�����7!*)�e�e�=.D���0;��`yos�=�ӽ�Jb�F2S(�R	��!�����.k v�F=:�[����̳����$n:�>w�x�7^�>Y����߱�%H9���EI'P�7^����-��2�ʃ����R#�6��X,�v�Ӌ%]VUN+) � t�l�q�B�������BH-�J��k�H!j��4��$�7�"�U"��b�`E`A B)���B1C�Y����S�@�J�#�F0�E"q�!Ã p��#��ݞ�	�����������e�N�gѧ� �/����  Ɛ���(������xF�S��y�@�q>�@ ��c��!=u@|��T���<8�6B��^m�f�M��76�P����D�R;��Ł����7^�>Y���#�Tj&�r)J8X�*��[%�=&A��-I�/q�Uv)su�%��mv�q"����;,�`�V5��u7�<�l\/[���[%�=&A���P`y!"iȔ��I�`|��ߩ#=�����^,׼�]���nT���8��lI�`n�T��0<�K`j�\�$�$n:�,͕Ł���$�_{��4�H%��zGf�;8~��AG6��H�$���V�d���07{* �,� 	A��[�J�����ufm����V��M(�ݺN�#d�s��'�1��V�aF��m�����=&A���P`w_D��H�YFe�)�.˛��?7lϢ""d�v����>Y��ߪ���Z�?Tj&�r)W���e~��0<�K`zL�Yϩ���8)I���������-��r&�eA��l�b�yAyEe�x�[%�=.D���0;���H���;�7���Ā .���ki�b�� � @    D[x;>W^���=,Sp�ê�(>�YG��+[=�ԝ�cҶN��І�����$<����s.�q�m�6:����bW�4�� �Kk۶�[D5���N#��b��y��`�/U�&�.Ja��8WV���(趹�m��;f��q,�:i2�{���wݏ���Ypu��(��v���k���F��z;f�y��[z\�L���gIH�
G�}��Vf����{���gs�1u*���J�,�ʃ��&��lK�0=��B�W6��H�$���V�;���>�`fl�,��օH��Dm9"`yl����w�����U�������R'J)�G`g���͕Ł�������`fwDGLNUP�Ȇ磪�mN^p&Y�x��I�
��K�Sd��Tj&�r�MH�͕Ł��� �>n�$��!���6E�\���]ݻ��s��}~���^z�N�Ӓ���`n�TF�a�fyEe���[%�=&A���P`r��`j��	�Su%1�)��lၻ�P`rޖ���-��6"%��n6�������\X�y�,�vݳ�9��dH� �JtJ�c>�	wFS���w�m�2�¸�wkh��2��1�b1�#j�N�`j��`|���v�,͕Ł��zЩT*&�r;��u�	D��w���g��9(�<��<P�Tj"9�G`g�x�36q�����0""0����"�	!w�D$~�s���l���ӈ�����)�S���������O����-��2El�H̰Y��Ŕ��`r��ﾯ��e�=&A���� ���mJb�JqF�G	���g���<��cն1qrDt��t�:T��"b#)���+�`yl�����d�y��yA��Ғ�"����ٜ�S&�0-�`���r�IL��|�$��Q�N�O�޶��lI�`{�$�R˼̻U35fK���N�V��f����"z���X�S�%HQMX�j���-����`n�t��-�+{."�Im��<�In�gjV�[��	���l'��+E�@�΄�I[��%��I�`zvA���������l.G>��JL��,��Vo;�����q`b+9�"F
F������u�~�7Xt$�}���7_b�>Fw&�J����N;�����ـ{��`t$�K���<�l���-����v�Ӌ߫w��|.�;���?Ue~��mt	$�I$�6� i�a�I� �`�    
9K�hݷ3��<m0&/�7#�&���2�;�h��pV��Stv���M���0rrb׋uӺ�7�-�[t�]����o�����F���[��n'�<p�/׮A��m��_Wvn	N+�V@!�N�n�7a����aC)�x��Bƞ���y�#�K���ws��h�:�&��e�891��^��(�Fj�<�v�]"Jtv��5�%Q��t8`��V�;���䒅�C������B'����(��� ��u��L����]Ӏ{�|Xo�e%H��Q6��,�v�Ș��`r���H�Y���*7Q����+3g��v�~_<�v�Ϫ5R�:r�R��X��`r����-��r&��1,/�b��R#Q��t'SώpG�
86l��cn6�q��q��C��n"vYӋ��ͷ��-��[��L��0<���W{��қ����$�_{��KO�|D��:���� ��u�B���wM�SSj�))�!H����3g��v�;���0�I@nq�D�`fl����u�~�7X�(J}ݜ`����Py��lbI��ջ���gs�>�X�8�:���"��$�9C+��=kCv:�΋-��)���d{g�j;E�hT�8RM�$v�;���t��������p��N��IR&����� ��8`E�[�d��D}P�)�S�ӎf�,[���ߕB�PWJ����!,�$AB��Q
�e�� �u�zE���Q����)7
�ߨս���gs�?�}���}T�z�X���r%NЮ��������9B���g��wŁ�w�����E% $�)�	*M�.y�m���FU�g;ub���sk��Dq�((��)�)��G`}�8�36q`j��`|����9���䠉�����Il-��&A���䌭~c"2&ڤ���˻���d�����d��J�B�b���32�z��K`zL�w�?}_:�%�G��%$�}��X/�o���݉^,Yy�����d���<����Ӕr:B�H�(nIHt9ܹ�l[0�M�Wc<v6�wv�Y�g���:�2��Y�����&0<�K�>����_ �~�5�~�t9"�R�p���~��[�;u�����Ł�3��7*&�*�P���;��������� �����%F�8�1�L��Ș��`�c�d� �G	@RrPF�36q`��΅3����7k�p��\�j&�%y��	@��x`��5�j(o	��:�q �`F	7�M�0�
�k`|��{���N"�>T<���'8��@���7@��Ɩ(|@����" ��
*B�`�5"�6#��bf�B���%e`??zB���/�i,��	�>"��>{��L_��Ty�U[�q�&B�BB%�����FUV������,�<>��#��ZX4��x)پ������w�����=���` m �          '@      �  � 8  ��   ݰ�`�}��     m�     �l    h                     |  �g�d�#�[�I���;sֱ�,h,9|q���и�C�ݕ������Z�*�Ú�F=h�sգ��l�K�L����+lv*S%C�'[���T�]�Y䉞Mہ�����Y�@�u�Yy,�T+81v��#���8X���q��9�V�q��O;��U���e��.5���!@��j��..F�7g;3��;iz�`y�C�ni��J>S�vJ�3����DNm��3��5&��+�6�pV뀉�|c|�e��l�g77I`3�\�2���k�k��ik)�y�M Ɓ3���������#��sq�D���6�=kl/c���V�e��ua�UV�U�u��Վ&qT��)���a&���m�%�Z��h� 

G�Āͨ
�|��gi��K[�(��T/(�� �UN�.�m���[F�[�yګj`Hr��UP��qc#[J�f�j%YV���qB�A��v�R�D�l�	��/�m���tqF��'0�	�b�a�h�KB@e�#���*K����j%�l��r�r��:ޖ'�wF�T��M�7�/W C��N![k��.7�܎:������gu�+��V�j�NF5nQ��ɍۗ��N��U�[`�	�:�-
o<\%�:���e.v��HVT
���	k�=XP�
��yŎz��S�\�|*Y���dy!�R�fj����f�'N�:���Rɜ��F,� O&v;^���&O�ݼW�s�4�W��Pj�5WO0;�ՠqSR��0�;N���q�9Nns����^��˺	Jw	w4�F�n|��?q@OW����'����>���
J ��w{��_��܉  m� i�a{N�  8    m�5Z�\��9к-���k�sX�"�`���evN6
1�K�ݹE螗�=����v������v3n��I&:@6�:m��,.MIK�d׶H$�i�kJ�\����mk�����?,X8�le��#\�&4ZC����YWhKa�N��.��8f�x���7s�G�UR����ͷv�[sww{]<�����s�9������k��uaM�;�Y�I�&2q*hbI�����,��lۑ07{ ��|vRT�
�
.�.�1��[vd��`�c��S�jB���qG#�3:q`f�A�nɌ-���r��P��+-],���`�c�d���X��}J(�rER��`����gs�7:q`f����5N�8�%-������e�9x�����.�Y;Z������1�\�j��3�~m�߿m��2��09wK`j��e������,ɷw9$���t�D��$J�T��(���%~:�~0�������_��5�t)�("�&~���<�K`zL���el�y�*RD�>�w����u�~nفД�y���2�yYF]�fe�<�K`zL�{�]�����q@(�O��N*�ݸ����m�۞y����4M�ی�z)$Ԗ���n�� �ݳ �� ���(��bK���V �����$�-]M%,͜_���9oy���vݳ�YϩE)ӑ�Ҕ7Vo;���áG%�Q"%�"#��ο��g�`|��$Mȓ%*�1H��w;��0�%3��,��Ҟ����RRr�)�H��X��V��v�{���cމH�1	�#)�9?n��-��>���j�V�ǃ&���Ե�"%���8X��V��v�{���Ӌ����tsj@H��`j�-���[�d�0=��� 0�˻řl.��&A����Ww;��S�jTJ��DR;[�`�x��n�2"GBDB_%�%J3w�V��|���4j�mM����<�K`zvA��,��&�; �Wb��X�K�5ik���8�Y�e�L���.�Sq�I!u��`rޖ���-����GL#;�r&�*�1����;���#=�Ł�޺�5f�1Wo)#r�c�dN;��Ł��ug���`b�y��]�$�)RJ��7���u`rޖ���-��}Զ!]��f��2����<�K`z_D�����I?^�w{�??>��  m���t�p      d���������.lU��u�e�zs �Zex?��k���uEtq�kf��q�uKAx���L���7�����c[Xêa�A�ö��R�jۋ<���T[�����-b�V����bȞ�&�S�UeNg��+2mv��A�϶�%�^��f�iZM�Z#}D�����_<��f�2�3wvt�Z��[��Ji⫃Lk���כ�72���z��GIR R�ۍ��yw��;9�+7g��v�ڧ ԥ��7u�yֹ��J&Mn�����?N�Y�""dr���u6���Wsjf�po?S��<�K`t�Q[.RŌ�F���,]����;{g�(S�����˪���ԫ��/-���[��07� ��:[ ��߰Qs�5^.�CZ����15��{qF�&c] ӌ���[׮t��3���3�%��W�����d�KuT�H�5.�)N8�GA��������_�%t(�f7ެg{� �Z� ��u$ӣ�ܡ҉	��՝���ku��
&w����b�?ljeH�_wyw����-���&�GL[9�Wj�R�Q�����{��䒍�ߗ��u`����u������5U�u1��ê�������<v�I�ƫKc�K���i�K��]E�G��09l����-���&��\�`�j4�5%X���-�vs�Vn�Ձ�3��n�$ISq�GrO/��rI�s��O�@"�`$H
DH@���E��rI������ռ�����T����{���޺�5v������y/xd������������t���l缬�tQ�"  rI)���}v՝ќ�r��m�,��6Ñ�+��:���O�Tہ(�
J�5v�>[��缽��A�޺�3�r�*@y*#n'��[��?\����)���@%H�nH(�v��Vf�Ձ�������`j�k��ԡ0�t��ÔBQ�������?O��i
"@�_��2!$ ��ʨN���7�^I?X~��Ŋ0r5R�%X�y�,�v��Vf�ՀWwt �RI)��$Ƽ�CI�0x����::'s�Ws�ۧ������*D�7$v�;��������u`j��`j�w'r����v��8���
?H9�Հzw������F%#Un+w�u`j����-���&�l�Yu���\����6^��?O��]k�J"�Է{�U�����R��tH�N;�Ss�r���}?��}� �z� Պ�����zo����@ l�M��5�2p�l    l���t��c�M���6�m���I��V��k��u��E�m�[�"����������F���c�p;a�hCj[.̧kk5+˱Eƫ/m]J��)�%3�&֩c��{���lH�=	�^�,��,��n�Iwn���ݟ4����qn|skSqp�n��lٶ��$n�������߮}�ߪWi-�W�1�ֽ�%�Ō�ܶ�/	�zv �x�k,ɣI�\�k�*7$JH��~�Vf�Ձ��������V.�%F�	��%"�3::`r�-����LEl�K���Ҕ9*������r�7��37�����#t�2R��$���.D��}w��)���$W�nS�� �I�`o=�`fo]X��Xc�V�ƭ�"D� �5)!�vP�N�r��h��:J�sN�S-�S	����Un/���P���z@>ך�A�Cn�Q$�PD�9$���o>D������zUT���/&������t��|vRT��w�Fe������D��}�����L�yN����(��X�yXf�Ձ�����=�`b�k��ԡ0��t����7�����/��}�`g=����ݿo��x�*���-F�$��]�w��1���v�d�^��n �IZX�Lۑ0=��06_E������Ձ��x�n�)Sq�"�>Ǽ���/�`n�t������$Wr�����I�`}�yXf�՟?�A��'�ا���P�� 1�бD��;��`/}�2�O��:�.h�8Z{�BHŝ	�NT��o<�y�����%�}�n�A<|0�-�t�Q�ξ@�,Y!����,�2ܦYL2�L��̹z|U$�3a�5`�0�I`��L�+�e�!	,���� ��ރ4�> I�f� �GQqU:�B��^|)�S�>E:�'�(�����!���9�����+ �K�eI rn+�޺�7����Z��IB��}8�7�R�")�D%%X��Xc�Vs�Vٽu`uwG�E)�I�"q�"��*�T t���V��Ʀ�nvYy��,뵯#�RSq�#j8���+9�+����_��t�O������������}�����Lm�L[�t�������R+3z���}�r&���	r�%��Z�Sh���o���?z��_�7���d/�@�T���T:�;�w�䓶}��8�R�)Rq�"�>Ǽ�缬��+q�+�Y�+�Q��J@I)ĕg5���]�hD[�l:�)�Gf���tݸ.k�	'r�����JE���V������J#􇶟N 73�**�B��r���pޭs��DD%2=���=��Vs�V#!��Ԏ��$�����}e�Lm�Lw�e%Hc��Q�`}��X�yX�yX��XWr� Ɯ��qD�������Lۑ0=�"`e}�Q����ϤH m� [Mk�I�  p    kJ�B"q�s� k�R6�t@��[F���H����6��~bA\��ͫ�N�" �z�2�Q�c�B�n�N��+*��v�"i˲l �m�30N5��,�		:G���N&�Iɱ��`����#5�\�3Y��N�x��tV��<�b:�,D� �Wj�ca���ǻ�ߝ��}#������՝f髚�Ņ�n��8�sWc=����:�s��J�
U�K�J��)&�����}���r����KQ���Q(9�)BqX��X�Z� <���ծs�(�2zM�,��'?
��)�����3����=�`n>�`j�w&F�'IS�Ĕ��6t���&mȘ��r]*�$�ST�m�`}�yX��Xc�V��,�{�)�	'$�	GQgo���ێ��n8c)���ϙӅ�69�L��Ȉ������;_����+ �ޖ������6R_��6���<�>���� ��AjJ�Mk��M���� �ˋ}(9Pj8�RE���,Ǽ��ܬ�Wꤳ_��]�zJ�F�**`�1��}��LmȘΘ��`s�Q*RH���V��V����goK1�+�U_�NW裍2Q��W�i$�9���ڧF2��qd�v�77#:`6�]�n���ᐣ�m�~�ߓ ����0;nD���Y�yI�L��'�goK1�+q�+�}��7Rޤ5M���nK2�����W�P�b_�D(_�nWt�ݾ��3���G%9CI7��r&��LgL`n�D��|vR_*9�*$mG��>�`����{���}���o8� )$����T�8!��0`���4rrs��n�p�8�jnl1��%$V��,Ǽ��ܬ��+��IQ��5%D�I,���"`{o�`:c�З)D�I"lR�qX��Xc�V��,͜X#;���JTIƔ���>n��]��k�Ј" BB$y�T�@<z����|��}~��2G):I�N!8�;zX�yX��X,�v��Uet�D�R��䒝;ٯn���-L=8�z�r����1�*��Բ�JJӔ��i�����V��V�;�����,A�3ȎJyE���0;nD���-�l���y�Pg�gt����l&�e���'��߭�l����"`z�r ���(���aꪪ����,��V��V�7���Mo��ԡS�`�cw�ۑ0<�K`:c ���{���/�� ���`{N� �    nyј�	��sh��J�øP��z:��)�mp����z%A�[v��7T�;+m��M��v��wi\'8��u�� �Y��KU�GP�H�Z��+�sG8��M�iZUBI�y<U�V|Ӂ�)�)�Nv�{]F��b4�I�
c�Ř���|�.9��Br^�B������wsh�F�<�T؞���<�^�RqK���,%�C;p���q�+%�95���RH�Cp�=�|��w; �ޖf�,?�3}�j�j��JE`b�߭�l���0;nD��#��2�'I�S�I*�3������q�+�Է�Hc�"���nK7�ۑ0=�:`:cPl,�Y�K*�I^ۑ0=�:`:K3g�;�FB �$�ą��]��~|��J[uWc��W��uoJ��v��k��0�O�JqQ#j8�7޺���`fl���}����}�7(��&�r��{߻��2'����ɿIŁ�����w]X���J�JIYw`�1���mȘ�0�2����J��&��,�ܬl��Θ�����
̵Yv��E奘��0�1��}��>m�������\�W�n!�ls���0#Wn�����9��u��j������&�N%$��7��`f=�`n>�`}��V���¨)	��i��36A��r&�GLgL`j�e�3)eZI]�`v܉���7���T(Qd�w�~�k�����bQ-U�/.�^&�GLgL`n�D����� �J�EI9V��,��8�����ŀt(J��r]5��5R�Ц��hul��vxF�x�eI����la�b�Օ���]+�W��������vGLgL`yr�%JIb�N+q�+3���3��������3��TӔ�4�Vl��Θ�ݹ��L�:+29I�nक`����}���}גo�HO��r�@`�ן�-�¨)R~n�m�,Μ0;nD�ݙ��03��bRb�04m��U΍%d�v�GN�]\�q�u��j�,��]�.��0��vs�q8�6���܉��#���07fA���줾T)��X�e�`n��l�ِ`n>�`}Z>��*%J4��`:cw��mȘ�05q�s2���*��U$��B���ߖ ��� �;��;zX#_R�R�Dآ$�`v܉���=^ �/ ���0?���W��TW��U��U��
��"�*�򊀪��
���Ѐ*��"(�0��� �"(� �U?�
������*��U��
��*���*��@�
���*�򊀪��*���
�Ȩ
���(+$�k"#¦ *�k0
 ?��d��-��    ���     
   "P   �    h|  8�@U 
(��!�J((���*���Q��B R��RETTDUT   5*     �e�]��\[׮o.����{�rӶ�x �iq���g��V}���o�ϩ|�= �2��:^��  O,_Z���>���Kۖ�K�w���s�[�yG� �|�  =� ���/s p<      Y`[�ɽ����������z�>�sC������ ;xN� \Y:s�\� 1L����zkq�vܱ'�� <��\n�����5����y�����*�@@ � Ϫ��ݵ�Z�f�z���_p
t�M�۞���w��J����� pN��jp �'/���>����ݯ�[����n{r�� w+�������ׯ[͔� |<���  @, �>��o����{ox�m�y�u>�� yח�|�F�&����H� ���Y��S;  ����@�� � �N�i���� QJD
P" w � � ���� Ġ   pʪP P � 
�0 )JD:w  )�� w u�( D���o-=���{}����� �)Y=�� ���v^�/�� ��'�ӓ]o���K��ͽY}��<��3��O&�7��ͽ�׀ D�F���J� h?�SoUR�h&F@<z��mULL D�*������S�	G�RT���C�ԕ&J4�"������������2OO{^��{���
�j�슠*�QDEO�*��������AQS�����iHD�"	2����!?��H�s��D����h�kl���!,�3y�ST�bB �6|Mw��uJ��2�k�>��0�{�������a� .�ćIs[�^�B2�پI���F���nc5��4J�U�8塚����(���ZQ��'y���kF\�~����-�ɬ�7��l�.�t���B� @�Ά��i�o3{|1���޴M�8���}���FMrP��׈RP�6��(B$B���)���#��r�K��댽&�s!R�n]p��2�4%�J�Y��p�4|��f��H�@w� �JbB�3>�	}�<j�,jA�A�f�A��������e��a2�9uɮ]��v�!f��HF�a	>�ɁϏ�8�! �ho$Za���h�K��;�k�
�*�G�81h�$+�U#A�1�1cCP�>4R4��5H�S/׿h#X���"R]�'S�1!D*@��!�J�`�%	fl��>���)	�<4��.:z�٨��@�n��6@�F��W�L���!IM0��) jg�4�^�Ir�#B��������%�:�l��,�O��{7�Д��Ϗ��6���/��t���c3���\@�Ye�h@�{n�{A�g�1��6|L��-�!,�!!,���/N�&���a��H0Mp��0#�B$��h$�R7c.asC�����Y%�u���}�kn��
a���ނ���Ϥ�Z��JF$�A��h���=�峾b߽����[��cd���\�׍�iK�q"	Hhe��"R�$ajfr�۷3\�1ì6Nk~��˚͚x�X�"�:i�d{����]ow�եgС�~~�E���y�y1�����*�Wwg���ق�/~��Dd���^ߵ/��K�o�Ls���s��x'33L%�s�����+�c�"��%X4R���7!Y�ap�����z1������6}�sz�}��Ai��i
b�`1�#p���s[H�B�A���D��$R���;ɢC�CY5���l�#��u��m!ZVXE$!��, ��R0#@�A�HĀ�R&JjLѦQ�vo{$%��!0�!�@��w��R[�޹�h���0a3|�o�{f;#[B�)�40��(bJH(D��e�@�`P�A���5X�	6��X�H"h1 ���)!#H�h�2h���D�!L�D`�2HD�ĆFq��1ۮFJ0"D����g	pw��\��;��u�
0���
G��y�2���o�9욄#bB$�(��P��	��h�+�atI�d�!���V���5~��A GdB.��!��5�Y��~�3�t||�n���L��7��f��c������f�Ba(JB���,+F,��oW~e��ȒH�$c�h�]xsy�]$al��2�xg{�Ȓ0��fk%�����a@�]�)��5��5���2I��Gy�qq"�	��<m�C�37Np��=�R1�����pH4���%�B#�B�, �"T`�D(*H�I�
A�	#$B�BD��+
1B,�h@�B�Q\
�S21�H"b`ƣ)"H���$JQ��9�4�XF
I�R"D ) �"�V1�`U��lH%�I �*04�n0!C�Q���/�Rj�H��H����I�FR�wE��%ch�4�d���Ia2�l,�4�����5L$��RkR��)2��,$
䤄L�RBXi�6&�!(Q�i��kR\���k���)Im�Ɇ7�&'�k�^���ۚ�&<0�!)�a5{w� :�36������lI�Ww�I�%	�``iaVb�@�9�$�04ofr�5�����v��
B2��HhHD�3Z>�F# �`F$�cï��Dng��a�xp��&BE��+�$���~H���\�vh�� Ire�y�o����}�}S��n@*˼14~0`�0��rs\��v��h%�D)������S���\��̝��5Ӽ�}��
-��	�����P�T����\5��h�i�sl��+�4l�04�*�@����Cq�0 S$x�{��%o3�}
���w���o_mԸ�s�k�r$�*N�%C!X��P���! ��dH��E����9�܄��9�8�9u7�k6m�5���H��a�lJA�p\D5y~��HX3+c	bF�
$�BB2$cK2\���"+�C�	�bH��֠F%�{�L�X�B- �swz�y�K�����&�7�p�͵ ��R$$�$j�B�����jv����8�1��B��ǂ��k�0���`�:ky�����Źfo`'4{���2'2)�#c�5�K���,՚�)����4q�տF$Yۜ���1����km�\��e��m�`�7͓4�8�ܑɃ,�6GF���q��wM����D���ւ^�	ӗ �JE3�$��H�)�������r빥"Y �,��B�`@ $Xѐ�R�q��Cr�)fh�wRnRs3Z ��%�q�F*XH�� b@1/���3�@��\�CXB�F���5�-�II]a+���h��� Hfa����	�� �X��BY�Z������:ǎp�f��MD�I.@�!���!�^� �FtR�%&$k
���V7�����7��4Jb[##!a�[��캛��9.�A�f�$���K�4�Ɩ+H$HH�kB�5.����9��p�G�ă���I:HH҆F���ٹsA~��ŉ�ULD�Ͻw;��w�9�W}�p�w閦����tro�~B������I(������	.�߼N;���g�3�4B�����'2��;��D̜�
�"@����c��5��d�ֻ�gy�ܦ͸y�3��u�$�4鸑#2�����kۦM]��u�欷{IM��f��%7VMB�<HIqS�A�a`���5%$Dݷ����w��y9�<��bحa�M�~0�����$ �Lf ���a.�1��S&4�9��q!�%K�0028i�3p����z8r H�-aB��75ÿl�ׂOfB$��![%d�#iIK��C4L�Jj����%a\%3S�v�3�&�m
��5��3�w��,�a�H��Y�2ˌJ�F8�D%�)p�	rSeaiIZ�Id%)!H�˒�K�Z4�$ F0%�i�R�h�WHR�4kD.��J�$���D)�Be,i	���iC5��85	4̒�-!i�Camr%4��3E��S;�&��C�D8s�
Cw�d�0,�!0�Z0�(`¹ "V A"��a�h�H�feΐ���h�2��X�!�!u���S
SH�j��%��
IR5
HFH�V@�V! ��"ZM��+�%�i��@H�R@��Ԉ�(l�#WVi"F� X�IW�,5����"hb��E(P�@�AĈ¡$Z)4I
A�Jl��00%0��p\�!p�j��1+)d�2KjB����\)	$$-L\�)��"B�fC5q4D����1���JbH�+��
VD��ef���� E"�l%�5y�B���y��O���<a�r٫�3�k���K�q�]�!E��l�Z�Λ�`C`JD�Ȕ����sz,Ϲ��>��!5��/9��9��vs����Ń
�7g�!��K��B��̀ ��                                    ��m       |�     8          �^�         �  ��m�            l�        �     �[@�  Il��n�o�^:$tȬ�k8�Ե�N�T	Kh:�bd�`� 59J�!pRm�u*��u�5�ePٶp7 �m˔r�m5�6����5�JKJO,G]l)�pV���I[;m�m�s�-�A�6hx��(  ��۷m�llp m�$�����-��(   6ٶ��`�h6رv����ݶ ۰�m���8���I����6:��R՚��M)r]���aQڭ7a   $L�*�H�e�Uڪ�˃�:L��/u�m@    m�  Xe�Kh6�l�    �mH$����$"@m� F�8����    ��m� �m���4�`��m�-�����7i/` [m�ׯPkz��.� j@ ��.�0	 u�w5�c��;YM�TT���Hj�p � �   m�l� @ۮ$�ai�Ā��V�.��ڕV���p-�  �m�$�v�   ��� �  $  �	     � 	  $     	 �m�hsv�m�pm��l �khG>��VU���ڀ��ʐ$p $�V�6�6ؐ    � ki�]�[x m   ��R�Ym��m��  =��m�V� 	 v�k�!  ��     ��pl [Gh 6�-���    ɰ��-��eejT7a�
ZN6�h � m� [@   H      HkX  	]�`ݫn-���bwE����u ��UUR�/6���\�+]kl  �`-� $��ݬԑ��`     @ �  �8� p�� hs� -�� 	 8l�$�ݳ�f��Ы���U�UU��Z���FԤ�P����F��  $m���zٷ#z�d��l�jف��������D� m� � � ���|> Hm%�M�e�I&�Y0H�  �p�dNL�n݀8�$6�Ue��`���i���ve�a�L���i�qr�ȪL�N�9�<�h@'�,�[u�UV�q����ds[� 鳑݇l�}�K�ݵ�J�u���Mg���e��Rȷ��L4vg]� uӀRJ86�͸�	�\�$���j�7$2�ݛe�m�$6]�[���`p�� ���Ysm��P�S.�[��gï��>���+j�9e]���WfmK#gf�Mn�  lڷcm�@%�f�sl9������h@�q[��i^j���d�I�FH$km� �H$mE�m�Gn���U�_e> �C�eۗe���ӫit%� h���Yx�nC&�\ݶ[d�٤��f݇N]J���/M)r�T�=:^�jٰ���:��e-�JW4���#���d�$.Mz�%�lH  8bm���@ �kv^(	��vs�P�Ӹ���0�:ڐ)��m�u��4����m�I� �Hm�H %eh�8��k���g���j[u^Js�*��NK���q�-�kn�D����M��`mK��f(��g��u9��cKad��rڲ�W�1�N��Ҳ�ac��026�m�Ė�3;vTK�Ts�J~.��J5���n��q,�Y�6��nHs�ڌ��3�v���H�	-�pp�ۭ�/N�L�J�u�i���xa�Q
���iZ�s�%�>����N��o[�q�����Ն� m�լ�TA�ذ�6+�^UvޅH�Kҳ��IWn�^��m�:)�
���ñ�3,�s�h� ��g�jYW@]]F�dK�	��܎� ��Ғr�I�i4]�\h���m�m��kY�0m�h�5���Y�NKX�m$B��mVjd �q� m��i� �H\MJ����~ñ��yVU����Kj�mp��79�ؖ�%$�յ�k�k��v��   �p�5�  �v�[Cm��@ݶ-6ִ�f�kvؽo���I�p�Ekb��
������  $��-6p-^�`��]uuUW<�F�� vKp j�  ��죝�� �`[I���m��` [S�Iy���5�h  pp�#vD�n	^j���! �V�UT  � -��h�mll@t�țe[C�۰�f��i$���&m�5�M�     ڶ$��n� j�Uyp����Ӎ���$5�ui6�[hm�6��K(ƄƒL8�ٶ lnk5Q�vٶ���  N��^�22D�K�]��%�M��ia'i��S]���$9j�{SI���  ��3������T.uq���7,8�sm-ն�k�c��Ym�
��ʪ��x � ��Zk9�r���Ke��==8��V�M%����M�Ge8�t�ۚj�pi}�R��܂�d�q�vZ�*���y`�$���4�N�k���;a[sP�v�M�5�]� )��U��4}����� �;f����2vt�u�(̒6^ٖrݻU��W+�}n>�N��iz�%�V� r��3�'^�V$KV�[{nY.,k��ܛl�I��.�9�S�L����v�犐��V�uu˚YUW(�����y���_H6�d�"6���9ZU�9�;4Y�j��*qH� *��Hm6�֤��m �6Z�����
WX�lh�6r$b��aĵS��nŲ 
d�U���M���pv�p-֩svSf��S�^k��dk%�h:Ɂa�m&�$N,�h$p �ZlÛkm˶���޷���r�e�Kƛ �Ij�U�	��V���ͶHl�'@mn�f���]��l��� ��$��E8���[@��Ky�f� ��ݻ]	�/8�uv�¤�>獘�X�d�lf�J��:v[��h�dr��2�7����_+�pBB��L�oc��0+O�7k��֟i���B��s����ne���6  �v�kI�H8   �6�  � h�m� �gI��cI���6��/J	-��ӡ�۫6��I�]$kh[@8 �[D�R��W[TH�km��h:�,5�m� 8 ��1m�cF��m�m�� m%����*�jm�fs
�L�HB@[�G>>O�>5�   m����I�p5�Ca���U������6C -�e��۞b���ԾZ�
u]�Ӣ�e@f�����iY��G=
�9�*�n��ݘ�ڶ�t,�������� �4���[Ru��� ��
���[j��mU]JJ��O+!2���u���q�l�I��	T���&��)YZ�U�v�h��#�S#�  	8l �J���e����V�c[W�R�R�cp��ګ�LK�U�q@T��Wf���J�ݺ��g"�w`��@$� ���ٶ  m��|�Mn��H �m84[hjv��R��l  �\�4��`8��m~9>��}@U�ʵUf��үZW�W�놪U�*�A��������j�* [M���H��$�m����˓Hݽ��"�U+1�p�bA6�n��ltS���ݨ.�0×�ɭ0����V�    6�m��ڒ� �:[:� ;ml�w6�v�9i[�u�.� O-�\@-ܼ����$�k���i�iV���kUë�X���ek��T�$��P ��I��W��m�u��Z,4N�:سK�t���G ~�|�gMg�� ���L��R�u[l�8��ԫU9�̢�Rmܜܹv*�j%����N�2�R�Wmn��Uw(UU�W��P�H9tΊ
v`8�h�^�Knֳ�F��n-Q���6���v�ci&M���  �����V��o�����mv�ہ�צ�H n1!�T��l�@TV�� �I��۶�8 *� �   � mK%�pm����E�ׅ�n��m  ��հp#���ݬ��q[U¶R�j�Z�ܨ��h9� g�U�5V�#�l�m�$-���H�ķ*�3rЧe���`�J�"sʷ\�.� �bF  ?>.���6ذ���2Ν[ki�tdū�h�MŞh��i ^��J��6     �m����i�zI����(b"���E�D� �G�qE@BT�D`A��E��쟢F@��W����S`��`V�R�@>T(�gTJ ��:��P0`�+���h/�}]"� ;[ ����*;��s ���"B uP^���^+�/��� H�`���N���~A�*tD|@X�@*���h�� 1N(|�?(��<0B��@F�D6#�E:(DEȠA |N�!�a�H�����ǔ�*h�EE��@S��	'D�P"#���<W�mDN�>T,v��Qk���D��U#��L]��`)�������O�<G�!$J���2��V����e"�IH�#E���6�@##$X���@�dYt�(&�4 H0@d�> *M"(p��'�O*� ����8����U@Uڏ���@"D�@�*� A�a �E,PJX�c(D�����ff��kZֵ�     �P�m Y@ �f�l  l  �8��{D�wc�]��>��n����&�C�v��&�\�]t�A�$��ɶ��RAr��v{i�muU�'\��N쪗AZs�@�Pl���Z�*��Ց��\GQ�T`L�n�$(�1�j�u���YR m�Tʚ�9�\�.���@ݺ��4YG+2��)*���V��24�ZL�lI���rP� �z�jA�^R���W���W��V��u��6�i�(�kV� I�%��Xk�j�l��z���N�]�\;Pl\���-+����ηQgH��1���ֱCFD8�]q&.B���1�ێ���΃E��̻���f�B�vh$wQi�Ԝݝ����񷋠�ͳv��(m�w�;Nr��#��I�E����-#����7k�=�m�6�>CYW��ö��75����ę����i��rOUp�r�	m��6�k��rN'�{�
@ ��jum���ZKi7l�;���X%Im�mn�,��`���\�����r��Ʒ�eQ�T6���m=��=mJ�N3�����8-[�T�u"u�e�]����l�[OC�[[���k{qݺ . ��v��ܦسhzy��]������Fܤe�����ѵIN�\�.9�dX�FRݖ��(fz��T���l���3Z�ugv
�@덊�,s�;롤��h8w��R���;<ٍ�˴ K��kM�yy�1�cO!�m��"\�	�n�C/6�0m�I���R$f}yb1cOq4��x�nm�@R&4O3����D�P�GmƤgEe��l�sk�-��)Y]�q�i+m�O��sU�:Ȫ��s)3[����4��.1�l�rD���4C�����yw6�Iurm����-�;lsz���1����j��6��r������c9�ɜ[�-��j�s$��[rW2퀤�&�׽��~�O�Qt�P��:�?8'�����T�0T=3� �M&�ȷz�;t��!9_#�H!��c9��n�,�����F�-%�.A�6킖���Py�n���&Ѱ�k��L�<-��l�]ks�ܜo��0�B�<t�<�v�O�}�����$�ەp�v����V3ېć 	�h犦��3������6z[^2أ�ي�(��ڧ�p���K�9���P��u� ۰p�J<��2[,�%�̒YnZ]��r�ώܻd���㱸�<Om ��&4	H��u�s@�s����ͯ���L���ܓ/����26ڒf���Z�s@��Z�[��{m�7�A�c�Š^�� b��P�n��Ҝ6�J$s4�ՠ{z�h��@����>]E�����ȴo]�ط ^rT�[�~�����ο��w�Auެ[.4bѵj��(��ƶ�{�zgxs�-��U�nj�F�;_������� {��ʀwtQ��o&8LhR-���ۙ�x��89��ED�"7��M�9��;�w4�ՠ}�șcX�?q	�iV���ށ���i9ʻ�$�Gss@(u&1��&�P�-��s@{��ʀ=�pW�L*���3ko37wj �-�rT yv��ց*�U_���bTV]��	����^��S��gY˙���f�=:����sM�M��ebF	V+�$��������yڴ��hD�$ȱG3@]�|��ط U�S����W`�y Ir�,���Z�&ր��w�:��D�@H�"C��fIo��� ��h��u��5$6�ͨ���rT |� �Y�wF�Q�F�d�ƅ"�-��h˰�� {���?7y�㔖�v��y=�OW�;v���{G�����\�v���间��\�1bn�m������+* �-��T @����v����^%�~m�o�\�W.��K�$��nh�٠}�;Fbd�NdM������@o�����*��h�mh��LQ�o�$��@��@>���]���0=^gy�y�)j�=ϻ!ZK$1&E�$rh�٠^빠w;V���@��y_*��"FF�œ��0�5��rZ�z��ͯ>N]�z7�@\�D���"�ĜҒz�nh�)�v�ZS��UW��"�\-��e�Ȧ4�h�)�r�d�m�@����/���m��	�L�*���+��� �YP����ժ�*�Yk/Z�˾���I��w��h[d�
��f85�#� �YP� m]��v�o�����,��uN��Az�s��C��d�UgV�m�4Q�r�ݡV�^m\ٷS\�f�k�eC��[p\bC8��U��<�(�u�ќngM�&q�V8�':�]�.�Sl�d>;mt�v�Yg;���4�vztg<n",�����tGH��X�c+�lc[v&)�6�)q��E�����V�݌��'f��L���`�{��ﶋ�v\������Jv�Gn�����0j��mH��P麧����uhn��������߻�j��+��*�w0�̺̬H�*ŉV��m�����;&ց�n�s�ZK$17�b	$����,�rʀu�� =ɉY{�	��M�&�~�s@�s@�m�@>���Quq�F�D�ә�w,�Z�����ʀ~�_�~�ݟ�o�g{����S���T؋0��

��Z�p�O=�t�T��z��6$����͵�?��J������s@��D�(�)��B�9&�}m���|�O�2����>>E�'w�4���s@�m�@(�Fc�PK*�6�v�,�j���hW�l¯��bIV��9Uq��h�h�k@����}O�J�˦��6�qɚV�4��@�۹�^�s@;�0EH�4�1�H��b�^p��;'s�*���vE��n#K�wHv^e�YFn���`+* �ʀUm�@;�tb��H6	�I�_�* �ʀu�� ]�u]7�{���h�&6�h���9[d�fy��y癍��4���^˲8�������wj֮� yv �e@/[��{�dN���4bq
4�yv �e@YP�w`z��㊃��hxiƮ�=�pqƧ���97<F�]���I�K$�d�-�nQ�I����* ڻ�����\��X�Ve%�bIV�����s�d�"Z�@����}�ץ^e�ebY�^$�h�� ]�|���*�ݦV�#@�D��h�f��s@�����U�v����=�nI9���aip����1%�|���'9�|_�~�@/u��Xa�M��#1DFɒ�٣#N �<��s��$�������#������ ��7�21����h[d��f��s@�k�$qF�	��%���w`���e@,��X'So#18�rM ��h�e@,�j��rn�Yz]�]��n�>VT�ʀ6�� {��=ϝ�1d���G#�L�/��h��ַ$���krN{�ٹ&���(�h T���# W�g5�j�U��V����!�J��ZwQ�v������QvԐ��;ΐi��ed��(R<ю:5�8�cv;l���u�v�@\���Kyj��g����lqڽI�\��lz�ػvP>������O]�[��	���9R�H�끪uU�\m�84G5��w1s���q��1����:������Jݞ��u�A�H�{�!��m�:��^�2Q��_.⇬WY8�!y�n݆�Txʸ�Ś�Q���'r'$���~�&�^�4m�������!Z�`�D�$�`�; �YP�2��� ;��I��rh�w4���U�M ���b�Υq�9#&�@;�ʀ6�� ��`+*�VԣrF@l�Ĥ��Um�@/[4m���)�{j��mb`�ak6AL�^.�ι�{a�R�V8y�k����ER!2Y8'o#18�rM �l�/��h�3��}`�H��@;%,�1[p˚�ַ$�}�蔇c���Oi߈~]� ����)�]n��i����� yԀu�� ]�>Y��e�16��N7��M yv �e@u uh�ᙹtfVݔn�� yv ���R��ɠ~����1�k$I7���DBE9��n����^�R�q�)��/My���h���#=(^�/��(h�3@��ih�@�T�RnA4�D���z�h[m- ��Zm3g.�]jV%k-Z��T����?\�- ��Zv�W��-���!6�����B8l��K݉�aR5e�!�&M,B�&�*`�*h�T�A�aKh���f�[0%hԧ�`�K(�"�"Dv2ZFt��"ggBT�,KQ���b��1"EF}�{E%���X��|	фHK����BJxrqٓ�����zt�{�%�����iS��>A"f������d�⑘a
@���HCn��!��fą�.�m�#;WaI�A
N��M�#<���N���	�#w�dc��X�1�!	��q�:M�Dp�M�����>T'�Ͻ�8yQ�������@:$hQ�>@D��O��k�ܓｯ�p>�tm�c�'�NI���~��C@}i���*�d�- �vJXH��I�N)&�m��/YM�m�@/[4��E�7Ɏ(A�8�a�'&�%��5�G����8�8��L��`���:�nX�FI�Gp�/YM�m�@/V�>��(h��y���b���,�h[m- }mh����l��S/e���Ihr-���>����&�vrꁹ��$�+� yԀ}k���?~�_�E]/3ř�����Gl�@���B��"���Zf�ڜ���s> �E�wψ��ȦA��$�F6��Ş9ջ�x�n�'��m_�m�q�6~�p�=i��H�	�	G@�u��@/[4�)�^����n���~$�i�4��{R � ���Z�V�1]�V^+Ih��>8��}m�4��@��!�L�)��p�u Z�������kE�y���bį�[xց+�UqȾF��>�w�>r�9]���I$����G6���t��i�7k͎u���@7+�� ��KMU�ya4��ܸ,������5}󫃕N���ŀ܈/;7.�6ɐ9n��zG��s��D�ݸ8�u��D�K��v۷>'k<�S�]�p�X&��g�KqfHn�Y:��(�)�;A �a�,ZݶN��4�� �yٵ��e��ԍw]������y�v��_�{���}�����]Zݘ8�N�+�M\�n;FGeN��2����Yh`���po"F98���@��4�ՠz�vhg.�i�	�69&�oJ@Ÿָ� yv�g7��^LB�n�j�=V�4��@��4_s��(�S���@������s� {���132�˼V^bĖ�>��Ssa��ߖ��٠}�,2��HLJC�5�5�͞;�Í��#m�Ͱ[�xy�u���FnZ���P�'�A�h���yڴSxԮr����(h�\��iX�Z�����@Ź����UVa�\�`ڐzSffbG���ؓcP�F�r(���?� � ^Ԁ=�p�Id�Ȍ"FG�^��wJh��@�[^�˒ꈜ�(�`�Iwj@Ÿ֮@u ߪ�~���?)�w�M�-�Wt���+����yS���\�s�镴
S���q<V�X���$��m���4����μ�^,U��Qx%e��䙠>�M��4�ՠ}ϱ�6�1���\˚��=���'�}�M�U�A�1DmAj�b��V)��_<�2���۲������R9ēƠ�4��/YM�mz�)�_���)#S#n6�^u Z� yԀwv��ݷ_�������-�65n;F�NN�����-ўɧXv�p�:����^3�Zf���nI��L�;ަh�3@�i��J)ፑ##�/YM��4�S@�[^�˅Ց9�QD��wj@u Z� yԀz��6�#h��n�)�z��@�e6O"E���H,�y��nf}���V��rB)�	���W :��Ԁ+� ��{������9x?b{k&��io���{w�'g�y�ۗ���s�� �#azs�d&ӏ�?����wt��m��=Vנ�s�d&6�P�-��7��<�$��f��7{��}1芼V$b�y�3�6�4��撪��L���~4q^���<y�nI!�{m����@�z��9�U\�a�~n����.�k,���n�	UU_ʒ}������m�ڮUW쾴�I*HH[ymp�M�tQkk�yC�������2%A񮝁^�[E��f��Ȁ�;j;f�\It:�����m�;L���/f�M<�u�m8��z�Y�v�{!m�5�P�\t�N���-�Sn+��l��l^^m��a2i�:.w����a:�b�Z`Eӓ<�4d�nocmy ��6K��6԰c�ˌ6�x���m�+�yy΅��̝͘qQ�C�����]���[kk�v�
�g=9
$m�a��qͯ;"��7�Ʊƹ`��{��~t��(�`�9�����-�����+�XI�^�ں�I�Ҳ�e�
��h�͜�]��I��%��S6W+�$U��q7"�d��E���=�n��U���[P�#����Zxg�sd�˚��35�y� �����b �`�`�`��߷�6 �666?����A��@�A�{��؃� � � � �ޗ��k!��I5�]L֦�A����{��A���@@����6 �666=�~��y����b �`�w{���wx�o���ݗ;�/M�;I�W�Ѷ�����v���$�c�a�E������ﭭ�j&�jf�\�ff��A�����o�؃� � � � ����6 �666?�����lll}�o�؃� � � � ����e�fjj�5�֦�A��������Db?���#� �
�����¬h�E� � 
uڪr<���s}�y���6 �666?����@�A�A�A����ִIs.��Z֍�<�����k���A�A�A�A�����A� ,l{��M�<����~��b �`�`�`����_ڗZr���\֮�A��@�A����b �`�`�`��߷�lA�lll{���y�����؃� � � � �a��߳WSM��f�VfjlA�lll{��M�<�����A����{�����y{��6 �666?g�O�̟��m�U����2ꞞQ#��=v*׷g:�'q��*�5�=��eئ�k><�����W����{�����y{��6*�����~���A�A�A�A���L�.a��,��.�֍�<�����k���Q,ll}�o�؃� � � � �����y�����E�A�A�A��/��ѓ52�k���M�<��������y����b �b�,*� �Z(Q +�*� �Ҩ�;�����6 �666?{�b �`�`�aʮN�Ax*V%I,Y���Us�U�,{��M�<����~��b �`�`�`��߷�lA�ll �A����b �`�`�`��?~�2�55sY��kSb �`�`�`��߿p؃� � � � ��~���A�A�A�A����b �`�`�`��߷�lA�lllo�[��d���f��&�fC�H�1u��m�mqݟR ;{nܗV�G�Di~��{����n�kZ�%̺�ִlA�lll{_�]�<��������y����`���������=}=���֜�����x���S6s��r��"���I��7��ʪ�U]���T��йy�$�hE��֞���W��\�g����E�@���4�ĒX �K-^#Br��\�$��	2K�i��*��(���aj-���X H��Eqϔ^����}�7$���\�s0�e�\՗F%Zx���r��W9^����{�Ɓm��L�qY�48�D����ۧ�K�`.��v�[�5ɭ�^��-�S7~�ww����a�e]�%$P�i�m�J��U}a$P�?t�
E�X�$�fb4�f�W+��.�"��$P�i�9\�*�v~�r^fYYYHV�bđ�I4�f��\��]�4	"���[���K(/2�Y�b�	Uʪ��&�@�(h�3C��9U�s��r����4K�~E��Z�u��i#@m�h�9�UW�U�s��x������hHS��=�)�`�%�H�Y�q*�b�no)sұ��=h�"-2'�S�H$�MG@Z B�Ča��>���V
���Hw��qt��Պ��֠sRMj	e���(H���	�=;�?7��       '@  �� ���!��	   �`��H[ԇ7Mӯa�iX�ΗK��d�Hm��7lcm���k��JKK^����jM�;`��X�J��y�@uuPY��R�6��]dp�j*V���0��R�Gj�p� ջUU� ����`$�,iڶ�X*��l۵V�5��$�����,�نUV��^���V�2�����Y.]�d~>��_��(�
�W��mtN�k��D��tf��v�n�Ю�%R��s����j�g���� y!��[���y����Em�Mz���Mv����7=�b#��&Ln��ףt-Ύ^Gl8{GH{6vi�[[6�l�'��b�nqs��0v_a.mh@u��&�u.�R��v۔ޓBu8�u*��.��w-� 7��ė��y�u"/"J�s�غwg���^q�x�K�ص��z��'k�n�ي�:��O/vgq3[\�	��Z�е3�=eT^N������Sjv�x��n6�v!q)��R��t��5 .ֶ��,���.�:�US��* 'Y+�W`�(���[�W՞G/k�F���N7����n�H�ٶ=��q��.�7fR]ū��0����7�0���<pݻljs��3v��4*���n�c{y.��)[J�!�p��Nٌ����>ˈ	����ݫg8:Թ�.�u�Nz=p|��゠�)�j�j���]�:v�&0��[�!�a�������s�����6�OD�jnq����� ����5�ӞtvxO=�a�U�sv�܂��=�7`�'X��Ʀ�\�*=�l��0um��mgmE��ОԎ&]��WS�0��}�|�X��N,�[P�V1{V�{a.��y�����cv��'Ig:)����i�3�4kd�ɮ�q�I���ԸsA�zAխ�m���] +U����\�<���X�n���\i�P0V�{��-�]�ݣ��RB:7w��*u_υ� �P���yAJ�∝��Ay�;�kZִBY]mp⮙:ꝪNݤ� anw!��%N�9�pM�i���ŋf�vq�6[:������F`�ljpt��4��VW���Giv��w�.�¨�un�����)�*����npH���cXC!<�c.��5L�v:ͅ�{)��[�Ϯ�f��r=���#�M�f2�4��q�!��^�3�"�u����볦�b�ێT���l�՗,�"��*\�'39�3	�U/�����wg���n]�[쉸��=�X�#�3s3�7��cpCl$Hp��?������NW+�X94}y�I`�!e��u�����Wdy%�E��l�+�vu�^K��Xb0�+J��K�:�f���.��mh�}�,0-U,�,W�9\�6qC@�okBs���ԗ�~���R�*Ib��h�3@������ↁ��4�e�є[��)b��%��m��ܻ�x��ݛ�^v۷e��<dP�)�Umn��fYYYHKZI#��k@}i�[L�s��W9���Ɓ�<V���&�h�9��)�Ǟy�a��{�(T �dT#	(��U���W*W9_|94ơ�u�����ve�R�\1R��ʴ��94�f����rM�H��:�?W^*�E��b@ZF����&�@�M�����W9����Hyz�ĒX*+W��ok@�U$�|�C@m�i����K����b�an]��k���4�;\���.y���ۦY�8�/��p�a�W�5j�tbU�E���6�=U�UUW�{���x���0�ZF��L�U�U�$P�$�k@m�l�+��?WrB��.Ҥ�,�F�$P�okO��
�r��*�UUII��6I�����
jkY���kSr "g��~���z��f��\�W+$� >�񚓒<0n$I3@�|@.g�_�X� ���@9YP�q2���F9������`�������4���M���Wd
#�}�����}�+y.�y�����C@m�hm�Ns����C@�tu�,E��b@ZF��L��r��rM�H��u�͜�.�O%N$�X!!R�x�I6��f��˹"��'���>�y�D��L���f/�l4	"���L��W.�|*���S����\�W+���u��~�,ˢ�f�H�i���\�^����{���k�}����o~X���@���.����ps]=`OltlԏL�󃡹��9��s�V����Y����(h����*���(h�䙕�̫�$�F���7������Oyx�Zf����*nbJ�V^,�ıqC@�i�N]�4"��v�ݷWx�b�u��i#Br�ɰ�#�[LЕq͆�*ì�R�Yw�ii�L�=\�{�x������h}�i$�Y��H��8�Ggh�#;D��sGD@,��͌C�7�/ ,;��%�Ղ�j�:r�"�C����t��G�������T�Jmq�1�׶��Z�p�q
x)��M�	g�<��i%�s;!�l�{qu�M��6P�ŻlW*�r��ձ��1�(wH[o�o����܇'��iS��X�P	��;�鸋I��虪A%��ڍs�A��w~��}.~�R�\t�Q�-1�3���L!�d3�{i�o���Ɏ�}��&��U�I%� HU�,D����h�3@�i����qC@�j�&^e,2����ni yԀr�@u 
�l�]�e��f]�0�ZF�$P�Zf��rE8��?�Ռ�/���f#BU�6�C@}i��S@�9��7�Ő�FG$4Zf��U\窪�=���{�^4֙�}���mӬ��.��Lv:�4�^@�5�г\��95�؍����������G},ŷ&,�Ib>8��6�4֙+�����H���ɗw��*WYYV�4�f�r��r�9U\HJ(hE��o�(�?6O]h�jYn[��S`zyx�i�Nr����ↁ$P�;�>bBJ��T�X��UUW$�h����*����l4��"���y��@��h�M�)�[e4��q�)��	1�D���q��C]̫��m����.�:��z5e��{��?k�T�2�\�Z-#�$�m3@m�J����H��N�Qs�Z�2��]�h�͕\��$P�$�m3eW9v~��fVg2���ZI#@�)7$���MʈXF"FE"!F�$�ڡ�rUUs��C@�������I,�Į�X�	��UU�6�C@m�hNr�\��l4���˼\�VU�����NW*�U$�W�I4�f���͍�
Ȅ�HR(��y��A.����q^p95ڮӷX�ur�;������BTZF���ր�L�Zd�W*�_XI4reʳ�$�*V$�@m�l�9�UU�P�$��{[�W9�s�\�`�K�f���Fbб�������W+�rI��I4���*̲�f�HМ�W.I��$�k@m�h*��r�s���+�"��qp"&7�8���m���S@��h�M�Ϻ,���iH�(�X<�9���ȣ�QA�*�|:3�4����Y�z?��[��2��1e��W�=�/m3@m�Ns�XI&ց���nbIe^%t��h�͜�U�$P�$�k@m���9\�+ܮUf��<���!]eeZH�=�/m�i+�\��M�H��v�v�,��\3,HHМ�r���$��s@��h�M��\C�E$nR�jҭ���	��I6$P��߿;�{����߿� H��hsx��\��%BZe�P�A������A�Fݕ`��N�s�%�%md��%�nnz�1͸��v얷c�r�u��^��;\�g���^2�����ƻ q�k˰�.�)��z��\qڠ�s������V��M������sY:�=f�5]�������i�g���"Wd�o������L�Ԇ����߽�������'��\V��������w�c�=�M�7�(��2@�[��d������Ӟ�ю҈�x�i��{S�_XI42�T��\���H�i�9˲96������mh���mp/b����v��6�ր�{Z{���(hE�uu�Ywv�Y�-%��'+�$�V�$P�i��9^��{����;%xͼIfQ�x��$�h��r�����M��������V�b�K/3�7m�F嶞�I^·]����w��>��`.�U�8��cǊHh�M�)�6���s�	"����ȃ�\3-Z�.�7$���M�"5��PS�"X�! A��H"����"HČ`�$ D�B,"	 $�E������Lр,�F0����B$��E���D�b@��a��$@��H@	��T���M~���;�h�͕ʫ���Eyyk1^$*��W��$�k@m�i�Us���g���@���h��q����Z�v]�6�4�f��LЕ�\�}Z!o ����YYhč���Ns�M��I&ր�L�~�n��8Z�J[r#��)��f8�x�,]i�m�wf��=cM'+�iZ۠��3+/�G�I4���i���>��(h�9WW�ZJa�I$4�f�m��-��m3}UU�s��\=��k��Y|Ē�=�/�L�kkj��T.v��QN��8�6Ȭ"��W�3M�� ����0�M� �=��Մ)`��H���CI�c{�W�i��D B$6©!�q$_�C��|]0���l"�"w a�gH�UT�hbJ�"X��ĪjiSD
�k�;HCJ�a7�A��M`�,i�
���֛�D�`�"Y2"���A"���@#�%�FH:;�ؠw�!�| pUO |��@'A�� &*�x�<��T�^�7���"��~m]���Z��ʴ��9q͆�.I� ���Z��ذ�I��l�!)����|�C@}i��wC/.��ے$�ە*`{d`�;;[��g:�k�A�5�N7��	��<���m�?m���>��r����&h��.e�b��G�@��h���U���f�Z.t�a�5!�>���o4�vG"�$����t�j����ZF��d�4	nL���7'�:T IBD�{[�ܓ�ϽWW�]ݪ%��K4}o4	Q͇�G4}o4s�r\.��h0KJm��I>��]�ݯ��T}�{vJ�8�>�����r<0N%��?@�OƁz�h���WZ���ؔ�Ȣ�<St�<�@��|� yԀu^Ull�7"#��*������.��P�;_���W�-!R��X�Br�73@�(h�L���@�]̭7�c�1�,IǠ[e4߻6.I��������I%IU�u]X�[u�uٳƊ�㡁Ί��x���N� @hU�Mͫ��Z�Bc��Bہϕ�Rp8;��e��7i��R�س��r�v���� z�E����u2ֺ\�v�Nt]�u�k�vd;�=[qPW2��P&�,v�;��=�1k-=gm����ܲ��/b8MZ�%���~�hӳ�;��l�����Z�1�;��Ͼ���v�|�� 9�z�y�Z�6��&�z�xǮ$8��꥝�S7����Df�Pr����k�*�@��h��A�4�4m��˲[�4	"����6r��nU��e�R��V�#@�����f����ↁ�d��}ތ՘�,�3"X�#�;�S@�e4k�h~��_��4��3���eZH�Zf�+���&��%�3@�z��>����{qTWl�k���]����s"����������&0�&!�I�'��pJC@����[���d�s���qC@t��$Iȉ�$4
�׻���<ϳ3 1QaUP�~9���_����~���Z.�"�L~F8%�H��L�Zf���Uw�d��Knf�w���Ve������s��*��`��2K�߻�W+�����<.K
�+"�!�{l��WuzwJh�)��,Af64�$Xc��o6�:^\�Y�qLZy�۰���r�\I~���q�1���I�n��[���)�_�d�9_X~�C@��b��Y@f+��b�wj@:��R �s�����g���1R,���4	ء�|���]q�r��ʤ�ۙ�>��t��q��4k�
���;�Е�\��h��"�J��Vb�2�+�7���ڐΤ�9����|��m��v,Fk��/9�^8���u�)jnND��]��x����ZgNF���π��S4��h<��Uz�`z罚!~�Y�,(-eڻH�Zf��λ����}`��4	�.J�Z��m�!�{_U�Uֽ��M���*�,cŗ	$g�8�
�נw�R ���y���×2�wr��Wu�K4��f�����?Lr�
�נwU�ǋē*i�o���M7")�&6�^��못u��n �;76&��nb�ӹAǈ$��/YM������y�es�֡�:��2V^b���1i�:�g9ʮsه�{٠G���o���`�z���J��]�2�+�=s����M���=���9}�V&�1F��X��@�S@�e4oJhg�^���h��ʖeҼ�Yv��4֙�{��s�{��������}UO�b�h�IO{{ֵ�kZm���9��9��$�v��6�Y3`�s�v���3�H�:���:eum�r�j��ա��[����q��Ɍk��N��-l�0��v���'r�Pz�@9�6��.�Si���Tj�ӁNu��v�M��Tn��	{��3T��7>�!e�x۶�V��l���"v�sӶw#�x����o���h81�vcݮ\�kt��"뗀���{���ێ��e�:�]=�u ���y6�z7Kv��Hb.�@񃡹ｉ���B(�6҂��/���hwW�w�)�_���U��chYp�ƼY����6s��Z��;4�u����#��zԒ<��28��~4Τ�9�}�@>�����p��U�I�W;6�^��y���9�ds���\�V^%wFe^"�#@��n �.@;ݩ yԀ{��`�t��+��n�� �.p:)ʻs�N�<)�1=��go w��p$������]���W�\��@��h�3�U�z�`w�=z����LQ���$��;���yy�V�3�3@���@w��e]�eȩf]
Yv��4ↁ�λ��ʪ������h��_-
��^ah��_蜽[�4��f���l4	2QWXe]Jŗ�x�@w��@�q��>8��|����at��t]��ݵ%��Y't�WD0�m,��vt�v���1C�%�G�9 l�~�z�ƀ� ��H|� ���������J�1$h�3g.�Ѩhܙ�w��;U]Ɯ$�pjC@���䞿{ٹ��"�'�h�"@�s��d_qC@�]1Ӭ��]�+31$hz�c�4֡�>�������:�ҌQ���&��;��$�a��P���@��tS���X�cm&M�:�fw�۶�ݺ�������uۣ��=U����-j�f�]�����(@>{R ڹ �v���_��on������|����W3\��@r/�)�w;�,m$\$q�#p�*�y�~�S4�9�UVg����=��>�7��bX�3u�Ś�U}oa�G�'>�z�J$ Gi�p����nIr����Ȇ���z�h���>�K�	nL�?w��o��0���8���䃣�T�[ȩ�7lv�9^ynj%6ۮz��,b��$�<q�@���@��zu2W9U_XG&ց�fH%Ib��Vff%z���9\��Z���Z��[���$Z�?F�(��Ĥz�P�[����U��^�-ɚ�.�	�&0iD�4��h���}o4'-��4	�.J�Z��̼���j���\�w�R �ʄ�\�D���A����k � ��R*�|t#�
��P�Hde�v��*(kx&���b�,�Q �ס��lU�Y�#��-� Iޝ������N�����       ^�  [@ 7m� � �����jL�ӰT�p�\1椹cc��ȍl��H��"E����-�9�Hچg�})+�m:���<����A�EeP�����l�/  �%�_m�In}@�#mp!�)Ͳfj�Tnm�j�Wl�:��u�sLƋ�
�r��m�.�/n��ՠ5�&��ui��������y{l���'h��*�YA�۬����X)sMUV�t�J��G)&��]��X*P�<� by�|��o�ݎ�lCN�8ح��y�s.���%kְ��p���A�M�����u
)Ͷ�MM�g8`�Y	�/N���t�Em�i��n����ݍ8���/����e���&�l� '%�K����ݢ�&Kz��[#��{v�2�s�v���z|���Q���Og�+&ӵ��n{Z��RvnI.U�g�4r;�9�xy��Xz�Jk;��0�b���S.�*K����r.�&�7Li�&���������RѹK9�f�U��;�y���Ipn�Tް������1/>�!��������<\�L�.U2��`���76�p�u��m�pZKfz�-����167��ۈ�{t<���I:��$�z��]l��]rgms��B�HW��N�hȚ3g���r����㎪��:7N�n��.볳=h��\v5����8;p�<��tٮ�GUñ4�KFsm�;:��^;m�fBw%@���k	>v�#���0����9�5�<�����\��US�n]�])�(܈'G���v�X4K�]��0�ܮ��.J�<ͩ �
p��6�p�ht����^�<p��`��[�[��	����y���H9�tT�ƌ#�����3c��LnML����%^۶�r�@Z�<�!�֩��v.4�1/m��#�����qG�U��\���\�@�-�yF�O~@�*�����#���� l���
�/�)�v��kZֵ���Z�D�utbk�9rF�ZL,X�m��mm��K�h'��Wmv���yH�7��0:�9�v���n�́�azI.ʛ��gSɒ�u��
v�ml%�϶ݓm�y�P��sr���d�0��Q��].�v���Y`yٍ�#rgm��5�<����]�-��!�d6�@R��<gZ�l�=����Z�6�����Ξx+��.��{��u���Â؋`N��6^'�u7S<�ru�ƞ�ld4 �sOG�q���r��BX�)f!��䙠w�S4���\�9��W��/eK�m�Ŕ�/u�q��Jh���=�)�Uֽ������v��=YbH��ĬH�==��Қ]k�;��;�[�51D�,�%Z��{ۓ4��f�����}�>�ԙ#�'�$4]k�;ݩ �<ʀz���ve�f: �G���>�sE�}#�ω�s�۔Wu�1f�9��I��Q��by��~�z�Ɓ�ʀ|�*֮@�v����]������9\�w��;'�Z�?=��M��h�P�%�ly��|�*֮@;ݩ �e@,�\"�3#�4Vנw�)�u�kB_��ՠ~쫗��-
��WXZY�w�S4	�$���jm��������ۡ0����N�0i��"�IGonWsQ��=a���N�1]�捪��u���|���v�y����W��qx�.,?/��Ɣ�$��{_U�ٞeUU��ɚ�P�?6���gi�W+-L��'6�ZW��wt�����s@��V�W�Τ�LO ��X�,ЕUm����Z����� ��1����(��������_���ܓ4��� ���t^a@\�5�	�ّz=r�v�@fm��.z(���^�r)�4��D��	��=�ՠ;m���2s����mhd��2��B��
K�;m�����P�$�k@��Mߎ�j�r0I���G�wu3@m��%U]��%�䙠��)���TU�%`�F����I>��I��{7 P��(~S'�����h��߽K1,0U��@��n ڹ ��H��[t%��N�2Z�4S��i赗�g��Ú9�&{]0���]X��]��ec���� ��H���-�:�]��ejA��G��Қ��i��%�����?+����.�k	�Q)� �YP�r�ڐ�n9<P�$�ly��{l��˭zwJh���-w���R&d�|� ��H�*�p����߻} ������7_I6vͷ�C�Ĝ2XV6N��l�U��n1��;��t(�K�#k��F��8�riT[nx$�!��,��p�t��[m�s���.3��uђ{'W-m�e�p{[]��.��`�a��!�ɼ�Ú���v;v5��WZ�k	4�:�wN�׋��j+"��Z�m4 ���a�@5��s%�U�L;�Rw6t⣶O��8���uلC`j�n�׮͌阶����Wm�v���g�����7$����)�^�s@��V�WZ���Ma��$� ,��-���wj@:���N����$���Z]kӼ�.�H�w4��ho�i5�u�� v�� �YP�WeM��y�ĤzwJh���=��hu�@;�V�$�~<n%01�s��r�����f�;��:{k���n�M�JzU���(���z����s@��z}Қ��vO"�#D�h�ʝUYEf|� �v��?�UWꫲL�U�eݒ�i^�*�%�3@�v�� �u x�I{Y��Qx+�,Y�*�\���m�4�6��T�9u�@�^YpQ�0ŎLY$���e@>]H_.@;�R �]��(�*��ɧk��{OJ�68�v�g�-j�y�z��΄t��5r�Lӡ��$�u |� ��H�� �wU�V�"��b�8h�׿���<�H��Ɓ߿~��=�S@�3�m��y�-ֳrO��^��w���ȧ�+ (Xҫ�����$�ۓ4���U��� q�Ĥ4����ڴ]k������']��rЭ]�Y�R�U�|�d�� ݩ ye@�.��ڽ��s�v˳�D��X̏N�qT���=�-]k)�R��6%E"fE"�*�r�ڐ�T��{�ۗ���"�G��қq!u���ڴ
�נ^ypQ�ı'�$4Օ m� ��{R�a�S�j"D�$��Uz��������@��@���|}���sZ��VZ�Wwif���9UUR=��G?nh^�@揄��I6
b$2���ƌ�հ�2�E��:3���]�k�$�i�7� ӂX��@��4��h^�@��z~\�Ʊ��`�Q�Hh
��群�v�5$�}k�Ԓ���r�_�B&��c�s=�$��Y�$��_����t5$��}�}BV��,lKXE"dRLz�I^�{�I[f�$�[�{�IUn�Ԓ^�
�T��&E�O}I+l�5$��}�}I*��{m���{\��1 ����+Fw���?~�8��k�
���^Ъ��Lu��T�Z�NI�L����؜pQd�Y�j�,ȷQ�FwF���^�u�i�nF3�h�uՕݝ�θκ�tמ�Nm�l촆�W��Nq����Fu��)���m��x�aλ�:h��g�=��h�b��ۭ��z;��.�i;&��+m!�q���[W�q�dܩj^;c�сt��݈���H�����y�&]y�\뛷�G�d�Ǣ��Zؤy0P���5�I����o��%U��RI+��}I+l�5$�c;,iDH��9���U[�����I~��O}I/߿M�RI^���Ԓ�r���F(�$���$��l�Ԓ���RI^���Ԓ��ǩ$��s�7� ӂHRO}I+l�5$��}�}I*��z�I^�{�I�vcX�c0q(Ĥ�RI^���Ԓ��ǩ$��g����n�K�a�߄�\���8hcuЛs�t��E�����n�v��/.��,�&zŢ1�͆��%U��RI+��}I+l�5$��}�}I+]����DȤ��$��l��0�`��O� ������v�}�����U[��$��«�19!��^H��Ԓ���RI^���Ԓ��ǩ$��g���ܡpp�%���$�RI^���Ԓ��ǩ$��g����n�K��ˍ��%���g���V�=I%�2����뻹"�6���[�����s�������-�[k=��cFXѝ����V�ёyLK�W�����.D���ݪڮ��?�I/�����RJ�7I%z�s�����~�������_�/L��_��%m�����o��%U��RI+��}I"��m�1��Q�I����o�����l���_#�B�!q*��$H1M��	s���Ad�1"p� E��!R1`��0��""���eaq�pCA$�BF�T ��0"X�e2�H��j@� �BP������&�`�ܬ�)
��	 ��6�1dM�di�f�g�!�h*o�`!��$�Yh@�	���l�)�������@�E�w	����+�
��ѭI���AbH!aFHT�4�%IP�#H- �Y+*�A�a&f\,�<��t �U�P_#������SB��(;�����-��{[&�_�k� �B��9���������Z�I~��O}I.�n�J��群��ቌKPE"c�LZ�I^�{�Iu�pԒW��=�$����$��Ae���K�s�V�,��!q���o(ӫ�b��p<�Z��AQLNH`��9=�$�ٸjI+�����]]�Z�I^�{�I�.�<q��L5$��}�}�癍�?ۋRI/����%���RIv0�v\mL�,�s=�$����$��l�Ԓ�f�$�[�{�I}��.%&�6�<I�Z�I^�{�Iu�pԒW��=�%s��|	b,`B"������1jI+�+So#�b�����RK������o��%��ũ$��g���ή����Xɱ��U��M�rgm ����s��X����=]��r-p8��2N
a�$�[�{�IuwqjI%z��%�����J����XƜ��[�s@[Z}{Z�{[9U����]f]�خ�Z�f%Z�@o�k@}ok@����uL�129��H��-�T� ^e@�`�hњ�W�f����@YP�T yvI=ｳrJ�
� UX��C�w=�{�<{ǽ�~_ʪ�^��U���s�n�@� \�0��mN�7h6w�ܙ#'An�u�;7j�5��"G(�^lm�:�p;�c���x�76_��u�V��A�V�o]�%A�.ԕ�̬���9�͈��D���t�.�n��v���GGm S�Խu�:��ۚN�n[��zH$�#���5���u�I�6���$�f���십XiG;Z���w����q��:J
q`�۔h����֙N�Wg��yG��bv@:)tI��"�.��*��׵�������W9_XG����l�P��6�4'3@/[ ̨�* �ʀw���ۺ�X��-%�7׵�>�����ͭ �~�הv`�1��SMɠ^���* <� ��>�sK1E��<���-빠�� ���>��h|�׉�� (�$�F���I�d8���9���r]�1��vعQ���q˅p�F�� �h�f���s�>��ͭ�r�7Z/Wx+��-{�{[$D,*t ��(*Db�@�4(12B%PD�R	@��罳rO��lܒ{�Y�wc�pP$X�8�I&�z��y� ]���;��������n�9khNr��r9�hr- o�h���>��*&��s���Z����ɵ�7׵�~�u�����h��t�Ɨg��%-��ϗ��ݏ��۶0��	�:73 �M��춃6������* �ʀ.�<��;F��f���y��+* �ʀ�4޳@�r�Ɉ�($��Ȝ�	�}훒O�����Dw���5���h֫��$�"nܙ�˰y��� ^e@>y�7^����X��7ִUs�O��?~��4�٠w5ɇ��L��
���Ǝ,�5zt����v��r�ֳ]�a4�u���h8�9&���s@���w[4޳@���ʰ�d��G2 �ʀ˰y��� �q�X�LnD�S���� ���>��h���/�s�L$��D�7`�+* �ʁ���U~�KurdE�W�8a@�Ȥ�Y��g�}��~����������Ɠ���* �ʀ.��`��������Nr�eS�e��½\ƣ!�v����-t<�kα�*�Xz���IR������ ]���YP丘�JD�&�3@/[4޳@�n�o]���;�Ȟ&'���� ��w�k@��J��v���ո5�$I�^�s@���^�h�f�ً�h�d��G3@��P�� ��� ���(�����ߟ@ ����׻n7V�VI���R�,���+�m�؛s&6�\0�񖀅��1�5�^y5v��E�zrp,V��d�\��nٻ<�)Ѳa.ݻuŘ{.Ζ�#ڻn��mtsǊ����y��k���
�^U�-rC����2WQ�kxY�����+��8\��wm��6�	@=K���b:�x�1�Y�ti�����\��t�j��ܬ����]'EK��Lp�X��&ud��q��7V	�mLY&'#i��	���l�y��* �ʀw���t��3M�/w`��Ty� ]�}xR�&0j'1�ܚ�w4
�* <� ��>;q��u�iwxe�+�Z����\�}Z ܋@�Z��� ���Ƅ�RL�(�� �]��+* �ʀU���]X���umڌ&��Y��[�l�Z����څOm����g�����MÆ�9��l����<���* w.�;�ne�H�48�9&���s}�;33+�s@;��oY�vb���E2A`�h��h���J�$qh�mhg+I���jcBs4]k�y�����T�Y�f]��fi�W{� ��yYP�T���m�����N�w~��ҵ��7"S��s�K�^�u��nȵdt�F4��2](�fFD�4���?_߷4z�hu�@-�4�F�~,��I�8'3@���|� ��<����eeݩ$�&
93@��zoY����:D�}�؊�8H ��U۹�}�]���'2cr R$ȖhJ�r��qhɵ�7׵�;�y�wq��y$Xؓ��h���-빠Uֽ ���/r¶�c�Li���h�iA��'3�ɤx�0����]�\0��O$d������[�s@��zoY�^�s@�8�F��rF���^*������U�H��#�k@o�sfg�r/�MDҘ7�)�~�� �ʀ/2�������ỉ7&�z�hz�hu�ri��V�(� U<׵�huQ�<Y!�Ɯ��׮��.@y�Τ�.�nQ�xj�j�s<��v��8q$�����X��4�Z�Q�E��D��H�0�ɚ]k�y�Τ�e@>幷�[Y��U��ỹ 9�`:�y� o���SRp���8�I&�z�h�* �.@y�U]yn�p�.��{�@9�T�\���M��\mĤ���<I��*�^�s��u �*�����*������D�Ch�
*�hj#� }.�48��h0�6�4M7F�T3I,RД���"W4�%ĀݯP���P;��~���H�ߐ`����w�1ꕋ ��3a�R ���$h�j����-��"1��~$�:`)��p�)Ԏ��`�A�0a�.��I�r, H�f��.�
C���       -�� �  �M�  �  �  �8��a1�{��������p
��N�<��jJ�8*0کh��� �vu���r0ErZt�i���P, <��@Q�P �Y�Z���2@N�<sp��� �����"��
5��mVʵGH�u�s��L�sg�lK)��|c@P�����sK�%^�ͣ,��#3:6��
�U��n^lOF�[N+Y��� �۪�(-�WI<`<��{.�P��1��` ��R�9�+3c�Z��y'ŞK8ӻv��o-�%�y���k�;mK��{^��&��u�S�Q��.1ї'cCdf"v�ar(�QhJ�u�l�C��ab�h�k+��Azs�a6÷�7=4 ��N%�js�wY�cq��Z�<�R��W�z5͓CÍ��Q���v�=������=�"�<7\�Y��^��-d��)�vX�W���ҹ�lgg�OWB��rncI4���]�Qs-�%�Ӥ&0�ޝ�v.Ň6��مU*n'k�tj:S]2���Nڰx��kpb5bTƺ�M�m�b�q/�V�v�;w/jMk�&��+ty��Y�"�(�y�3/�{m;ν�]G�<�6:3g] ���q����R�Ů]5RD�J�[�d�ɳk��=����@���9G��h�47�����0]�f���qF!y�ʊ7:�7Tn�M�*����X;qٸ:��l��2�uN�9����wm)���<�ؗ����t�ڦ��j�8<=�T<=�Sۢ�;j��gk�I	$��Zl[9طY��Rt��k��Vԩ��xu#��"t�\���`�:�)���Vl�	JۮG��s��!��;;�9�E�hݽ��V��&-�3�Ȧ��a�#h��z-ۡ�|��+�m���5��RntƳN�&*�=[/F���dH{F��ke����v�1<J7HD��+�u�������{���b�:�T_��6@AdD�)� #�Cb��z������mp�b��TQ���sg�EC�ә6��9�\і-�Z�T�[�S�0;(�6'���Ч9zL�F�b=�z Ѻ뎎��,"��G�Q�!ۺ`"���h�U�֮\㲻��n9w6���q�!�p��يUj�M�!cq��;lٷm,U��`YC�ݯ/c]s&l�Û�{������xx\�gm�[R����P���;��{������֬eذV�By�M`��[y0�".�xyч�/4�rD����JF�Wig��k@}i�_^ԯ�%�3@�E�sƣi�4�S@��s@��z׬�/�G\�d�I��/t�s̨|� 9�`,��TI�$��E0�ɚ]k�y��* �ʀ}�sov��wB�V^	,��k@��+������6�}o4	U��ru]K�����be����ޖr�#�h�=;�lo\��[�.6聹�X�N��#cq!�'�~��nh�w4
����}`~�-�\�+R�aywt,F�}��lN�� �fO\��rI�u��w4��X7&)"��9�|� >W`,�w2�~����m(4��%#�{��/[��{�w4
�נ}x�Ԕ�j69$� ��� o� ���=�8��Qm�cKt�s�6����n��٣]��ً�'vt�����g��uh�l*��׵�;�y�w�J�U}a�Z����I)"�4(�������h���=�jؤɎH	H�$�@=�@�n���Ǉ��g��Ƃu^)��3�ٹ'o}�ܓ�����K00��vbIhJ�r��9>��ss@��z�u�f+U�FF6�F����T�\�w; ye@?��\�̔t��Oja�Yў��;nͻV�wb����ld�2$ϗ��Q��/6��� ����*�s*���Rn�N	bN= �������U��Z�Z�����W��2����̽݀<���� o� ���/��T�d�Ii�9�����z��f����܇��DӲ����H�6Ej!�3@��� ���<���� ��].ѹG$�9��⃪ۂ5�6�I���瑦�����k��^D�]Js���]�$���} ,��e@��<�4��̢��6�wwH�* ��P�r~�M�k��Ɏ4�,�C@�uڀ6�ݩ ^ԀuZv9���$BlhNf�U����4zSC�g��_�����M��r	��IǠ?�L�'*9>����������*�Uڕn���d N���Ny9n5���
U��rs�wF���NR�v�%֬�)��,nv���h@�;b��S$�Ӵm{G�V}��%��V��$��-��g��:©�3�R���Sm���d����X�Epvs�N����a��6[DJ��s��:mi�F�sP6��ʝx�j��ʻܶ��Wc�vrl��RvȺ�1�~ww���۾P>�vl�ED�.t�r�&pln*��q�k�<�^���s��^'l�Ѫ�ݷ�������2����ڐ�w|���tۻ3��j ��P�r �� /k}�Ur���rTFV`$%��a��h��d�j@YP�ʀ|��n�<�A%$L�=�Қ�w4o]������ �J$ĜJI!�^YP�e@����g��Y���'"X�%���_fO�B�R�іf��D���H�:W�zP���;��dv��\��9ƛ����q��oq��������ND�,K�}���Kı>����r%�bX���ʛ�bX�'ü�cq�"I�!9��zy���#̮�ى�a 2t �� *A|"	�4�/"r%����M�"X�%��{6D�Kı9�������{��7����eV��8f&�X�%��~ߦӑ,K����"n%�bX�����Kı=�տ3O1b<�y�^5ّ�FQ��5���Kı=�fț�bX�'=��m9ı,Oe��q,K���o�iȖ%�b{>��4֦��2f�f���bX�'=��m9ı,Oe��q,K���o�iȖ%�b{�͑7ı,K���&I3Y,�Y�C��M�.x�T���\o�.Ę댈Wl�Z��Y�ڳ,*5�{���oq���~'����bX�'��~�ND�,K��l���%�bs�{�ӑ,K��fl��II$���y���#��~�ND�,K��l���%�bs�{�ӑ,K��_{17ı,O{랐p�DƜJI!�g���1b<�nl���%�bs�{�ӑ,`^��W��"� v�D��,L���bn%�bX����6��bX�-������k3	Iu�&�X�%����m9ı,Oe��q,K��~ߦӑ,K����"n%�bX���ə��kYnl���"X�%���bn%�bX�w���r%�bX���dMı,K����r%�b�~�<#�~[G���a۶x:�L��&���x�m����1ghq0�_��ﾻ��YUnL�����Kı?{��iȖ%�b{�͑7ı,N���ӑ,K�ej���<�y���[��2(�`%.k2kZ�ND�,K��l��@?(��$��߿i7�O������H���i7�Kľ�[sƚkSV��u34D�Kı;�{�ND�,K�}���Kı;�o�iȖ%�b{����i�#�G��3޷֞F�R%rjr%�g����ى��%�b}����ND�,K��l���%��@����ND�,K��ގ��VवK��{��7�������ʹ�Kı=�fț�bX�'{�p�r%�bX���f&�X�%�{�~��o�n�s`�q��7=u͋6�6�D�@S[�8F�O9�_�G�w�͠��Y���Kı?~��"n%�bX���iȖ%�b{/���Rr&D�,O����iȖ%�b�R��[2�֮ai.�D�Kı;�{�ӑ,K��_{17ı,N����r%�bX���dM��L��,O����L�Lֵmі˚6��bX�'쿿f&�X�%��}�M�"X�%��{6D�Kı;��iȖ%�b}���2�2�h����5���bX�'���6��bX�'���q,K��}�ND�,K�}���Kı=�]�F���L�.�k2kZ�ND�,K��l���%�bw���"X�%���bn%�bX����Kı:���kZֵ��¶�U��0.$�*`�V�:ȳ�8��m��ŗ�i��]���dꇳ�G^�Y�䧪�6����q�M8���z۱��s�`��y�3o�O��ݻ��K!�>su�v����F�@Z����m�꺞6���2�.�X�n@Y�48��nc9bM�8�&��n��:ջY�2هm�r]��N9�u��2�V�-�3kn-�і��_�F�(fMܶ��R�r8$I�P�i�ۀݖ:z[/,Y����m�fJ����V�\Yn����,K����"X�%���bn%�bX������L�bX��~͓����oq�ߟ����vՐ�E��9ı,Oe��q,K��}�M�"X�%��{6D�Kı;�{�����7���{������-�T���%�bw�ߦӑ,K����"n%�bX���iȖ%�b{/���i�#�G��3�=QEi'�p��Kı=�fț�bX�'{�p�r%�bX���f&�X�%���~�ND�,K�OfK2��k5��]h���%�bw���"X�%���bn%�bX����Kı=�f��b<�y��/r�%�!&!�[rc����f�^6���X��,����suc]�i���kV�d��Ѵ�Kı=���Mı,K���6��bX�'���q,K��}�ND�,K�칖�&f���KsY���%�bw�ߦӐ�&�VVE�BU:��lMı3�͑7ı,N���m9ı,Oe��q,K��|�̊%�l��zy���#̷ٲ&�X�%����6��bX�'��ى��%�bw�ߦӑ,Kľ�Ks�4֦����fh���%��D��ߺm9ı,O�~�Mı,K���6��bX�'���q,K<�y���$G�HIMɛ�zy���'�{�q,K��}�M�"X�%��{6D�Kı;�{�ӑ,K=��~�{���,q��On�F�ݹd�y���4r��1��u��$�L�9�Sv��uLu:�֩.�n�����Kı>���M�"X�%��{6D�Kı;�{�ӑ,K��_{17ı,N���f]]]e�fj\ֳSiȖ%�b{�͑7ı,N����Kı=3޸��bX�'{��m9ı,��/�ٚɬֵ�R]h���%�bw���"X�%�����K����ab��5"�I�n��2�J@��
�i�m	
R���J0Hĩ�J�7��8�&�ݤ���9�[h���B$��;�FBB�:uKbB�D��H�*��J�!��k+D!s���$$3T���K 3%BVQ�*B��$���+���5aX�$e���Be�FSJ� <�  ڠ� C�  4|����:�U��E�/v&D�wM�"X�%���͑7�q������䭚�k8+��7��bX���f&�X�%���~�ND�,K��l���%�bw���"]�7������EX̓�����,K�׽v��bX�'���q,K��}�ND�,K�}���Jy���[V�PBy�m�2(��3l<��Y�1�گZ�l�+h#n�&��`B,�]Y2ٚˬ�5���Kı=�fț�bX�'{�p�r%�bX���f�r&D�,O����iȖ%�b_����cu5um̗S3DMı,K���m9�r&D�?e��17ı,O����iȖ%�b{�͑7ı,O��������&��7����#�G�Z���Kı;�{�iȖ%�b{�͑7ı,N����Kı;��f�^���_w��oq�{w;���}���9ı,O߿fț�bX�'{�p�r%�`b��DA4 ~"!ȗW����Kı=���f]]]arLԹ��]�"X�%��{6D�Kİ�G�s��v%�bX�������bX�'{�z�9ı,O{ԛְ��B;[���%ǰY�=�N��M��6g�<G�s�![�[3F��:{�Ou�bX����Kı=���Mı,K�׽v��bX�'���q�#�G���Φ��$������%�b{/�����#�2%������9ı,O߿fț�bX�'{��m9�*TȖ'��3��e�Y�.je-�f&�X�%��߷�m9ı,O{ٲ&�X�%���~�ND�,K�}���Kı=ٯ{E��Y5�3Z�S5�M�"X�%��{6D�Kı;�o�iȖ%�b{/����bX�'{��m9ı,K�}s��f�][s%���q,K��}�ND�,K�j�����bX�'�~���Kı=�fț�bX�&�;7��� 	o-�Ȓ�פ�.i^	�:�4�Yx�B��,vճ�M��0i.����n�E�m��H�i/�nw����)�Y�!���M���-هu�;�O;w2�nŜ�fTad�.�ƈ�=�mtW���Ԙq����\��v��mϟb���}��Z���zM���ܜ�&�J�B��m�k+�[x@��ܝ,�0�EC�R޼�Zݐ=�w������9���u��K��۳ۚrp�sՈi'n!��i��w8{hn��h�8�]����=�{��b{/�ى��%�bw�ߦӑ,K����"n%�bX���iȖ%���������Aj�����o'{��m9ı,Oz�Ҧ�X�%����6��bX�'��ى��%�#̿rڈ�j,L��|�O1b<,Oz�Ҧ�X�%����6��bX�'��ى��%�bw�ߦӑ,K7{����ԅG\v�ﷸ��{�N����Kı=���Mı,K���6��bX�'�u�Sq,Kgc�]Q�9"I��JL�3��G���}���Kı;߽�iȖ%�b{�^�7ı,Nw���KǍ������X˰�#qSk7kk��ў�9�t<�e�X�[�����f�13��KsY���%�bw�{�ӑ,K����*n%�bX�����gbdK�������Kı?}5��-�N��l��{���oq���~~�=�B
y^b&�j%����ND�,K�}���Kı=߽�iȖ%��1S9;���8$ؠ�����1'���m9ı,Oe��q,K��~��"X�%��]zT�K��}���#�$ �R	ɛ�zy���b{/����bX�'���m9ı,Oz�Ҧ�X�%����ND�,x�����ϩm�N��_w��oq�X�����Kı=�J��bX�'���m9ı,Oe��q,K7�����?;[�y��-F��E!ܮ'���u����X�� �A����@�<sΥ�f�m9ı,Oz�Ҧ�X�%����ND�,K�}���Kı=߽�iȖ%�`��e����[�j�)5�J��bX�'���m9�r&D�?e��17ı,O�{�,�r%�bX��ץM���S"X�3�=�����+��7���{���O���}�ı,Ow�rͧ"X��	�P�$#!	 �@�C�P2'"g�ʛ�bX�'>��ND�,K���������8)}�oq����{��"~���ٴ�Kı?~��*n%�bX�����Kı=���Mı.�������؉V%�}��oq�X�'�u�Sq,K��~��"X�%���bn%�bX���6��g���{�����Ǿ�0㱢�Zl�nq���Y��]�v����rOn:3vY���;�52�K�u�Sq,K��~��"X�%���bn%�bX���6��bX�'�u�Sq,K���\֮kRMkZ�L�h�r%�bX���f&���DȖ'�~�ND�,K��Ҧ�X�%����ND�.TȖ'�/���e��Aj�����oq�߿���Y��Kı=�J��c�"~�߸m9ı,O�~�Mı,K�����,p�Ѿ�7���~�v�"~�w�T�Kı?}��6��bX�'��ى��%��@�֨`�� �����x��"X�%����3Z�u�SE&��Sq,K���{�ӑ,K��_{17ı,Ow��6��bX�'���q,K��?������؍a7����.��lݣliL3����g����[��|hȅ>9�a���֎'bX�%��/�ى��%�b{�7��Kı=�fț�bX�'{�p�r%�bX�L��MfutL�MR�k17ı,N�ޜ6��bX�'���q,K��}�ND�,K�Zߙ���1b<����F�M��S0��Ѵ�Kı=�fț�bX�';�p�r%��C"dO�~�Mı,K�~�6��bX�%�>��1�52�K���&�X�%����6��bX�'��ى��%�bw����K���ȟ��8D�Kı;���kZ�a�I5�k5��Ѵ�Kı=��f&�X�%��#�߿N�Nı,K��fț�bX�';�p�r%�bX�|��ݷ������Ŗ�'ln��U�m���--�i	�*cύ�􋾩z�q%�m;��)kVK��L) ����t�c���D���m0g���N�(5���ލ��3�� ���(�7	����y��c����2�Kێ�D�B�˶�5�i��D2��#����6��v{:�n�lgj����rt\v(�,]�;`˧���9&�x��{��?c���<��F��ձٝ��5�����Q���@n��;�06j:�6sK]�N��_wbX�%�Ͽ~�6��bX�'��l���%�bs���򈓱2%�b~��ى��%�b{>��f\�����K�f���"X�%�｛"n�c�2%�߿~��Kı?e����Kı;�zp�r�bX?e���̗Z�0���q,K��}�ND�,K�~�bn%�bX�������bX�'��l���%�b|a��OY�sZ�sF�[�ND�,K�~�bn%�bX�������bX�'��l���%�bs���"X�%����zk0˫�fjj��Y���%�b{>�=��"X�%�｛"n%�bX���iȖ%�b{/��Mı,K��C�٭qR�ZV!y&��r�Cv�rzk��=���r�Ւ�Uq$+�����ı,O}��q,K��}�ND�,K�~�bn%�bX�Ͼ�kiȖ%�b_C��L�4L�˙.�戛�bX�'{�p�r�X�L�bz}��n%�bX�����ӑ,K���͑7�eL�b|}��5�Tֵ�ff�m9ı,O�߷���%�b{>�=��"X�%�｛"n%�bX���iȖ%�b}����k$�ְ�Z��f�7ı,Og�g���Kı=��dMı,K���m9İ?*"~���Mı,K�j����5m�MK&���ӑ,K���͑7ı,N����Kı=>��7ı,Og��kiȖ%�`�߳'��.�0���w-�ػ���{c��9���p5ʘ��p@�i:#4駞8+��q,K�����"X�%�������%�b{>�{[!�$O{�:�H'J�쾳%�j���.�lI�>�}SQ=ı=��{[ND�,K��l���%�b}��iȖ%�bq�t��QL�XI����1b<˞�{[ND�,K��l���<�ED�O��p�r%�bX���\O����{����t~~�,�K��Ȗ%�b{�͑7ı,N����Kı=3޸��bX�D��{?kiȖ%�b_�������[r˩��&�X�%����6��bX�������r%�bX������r%�bX���dMı,K���e�˚Բ�	�V��NN��5lg�E|��x�	!�5�x9��������{���oq�X���\Mı,K����m9ı,O{ٲ&�X�%����6��bY�7���?���Ob��/���7��b{>�=��"X�%�｛"n%�bX���iȖ%�b{/��M���ט�1e��"YPA#�|�Oı?{�l���%�bw���"X�%��{17ı,Og�g���Kİoe��k2k5�0���q,K��}�ND�,K�~�bn%�bX�Ͼ�kiȖ%��z�DQ?{�t���%�b~0�>�ڹ�f��sF�[�ND�,K�~�bn%�bX�Ͼ�kiȖ%�b{�fț�bX�'{�p�r%�bX7�����L��ޝ�������;��F{m��s��k9�$)l�^H�-�������oq�����m9ı,O}��q,K��}�ʓ�2%�b~��ى��<oq�ߟ����2�bX��7��bX��ٲ&�X�%��}�ND�,K�>���Kı=��=��"X�%�}	��n9�3Vܲ�fh���%�bw�{�ӑ,K��_����bX�'��g���Kı=��dMı,K�}��4kReֵs.kFӑ,K��_����bX�'��g���Kı=��dMı,K���m9=���ow�~~{�=�L�﷋ı=�}��ӑ,K���͑7ı,N����Kı=��f&�X�%����I�:5ذS@J�P��"$H
����4�^�>��i��f`�¬�)�i?;� �F������
�9�m)
+N%��H�8�H�H�Cc4�t	���]�)�&�}�D�@���t �
���� ���*B��	0�",�X��I60�E4��B ��|޼�&�&
i}�~r)����%)h�!���),�������֐�!����#!˘�F9�n S+��@�!9�t�iǫBvRV\v��u�y�]�\0;�"�6����2D:��i|:%�]���"|ˉ߾�`|���.��X�]rh�X1X�Sd�ixt%%��:dy���q Q�1� \0���0q�0kl���1	��9)X�5e�7)
1E��l�°F$�� ���Qb�ĉ$XДHѣY 1�!3N/OOw���{������       �P  ��,� m�H  �  
�kn��3�\:��5o9��.���Y7aӎ� �F��^�2ŵN(�H���R��́ܠ7A���U����#�5]�L*]��[*��UZ�,�e��mt�����Y�+c�v
`)5:�٠+`'D�0�UP�{-N��p��)[I&m&��5�*-�˺u<����W�M�n ���i�.M��J���(FZۃ�a�JػhFZ�vwj��.MROn�gv�_���8��s�M��\v*�G#fE�8���XAC��͌� ՋvwG%�m�ћJ&&�{���ݍ����mʜu��&s0��\�B�pQɻ]B�(���^����u��i؁k=��ʱV�9�d�sm1�m;�f�IS�I[zU��ç@���x�[�1�o;��Sl�*N}�ph3�����#qz�ay�-vV��χQv�^�P�I�lh1���66�^Uz�N��{,�ڮV^]��U��äb�,���sMJ�)N��ez�N�)��i	j�c�������ɧi�U�d^��,�v���"n��"�۝��[]v�Wn4��(ݶ�e؃�C���v!)lxp�,�q�N=�4�M�eH�`�͞ɫ�KFu�����mˎq�[.5��g�7i���p�7�T1�2*�b^�m6�	%���fOpz%%͐���8���F8�l.Z�c���.ۗ[��lq����m7*컁Ⱥ��|���]28z��6�l��a���ҽr�FCe�� m�D
Y�AƷD]Wv��h�BH�j �'Q�:�Ύ�K�������|+�
t�͹��(t�`^���Cճ���:���p�E�.�2m��emm�Z�fىs�Q��!�%D�p"�H�V�ό��q�z���<k+k/T;&��,[Q�dL�+����>��[%E.���V#/�#���ڤ΍�oYM��P���n����hfh�4ŗΝ�Է\h��5�?�PQ0A~� �B#�C�|���"�L�u���j�^�.�n��]tp�*�JG\�&;\��S�.��0�L�;߯��2�ӌZ�nf�HLWW<�{k��]��7]��ђ�'�k��.v�h�d6��j�9J�cU�RN�k763��Urq����F��n�W� 5�ⴈq���]g�5��nGC�� ��`ڽv^tƌٓ��[����&�.t�D덊�6���!��w�wx�ccl��eё)�r7
qqh�#mا��Du�p/�n�����Ғ:�̀�KS_{�w���x�=��l���%�bw���"X�%��{17ı,Og�g���Kİom>/��d�kXaIu�&�X�%����6��bX�'�����Kı=�}��ӑ,K���͑7�ʎ����~~���M(�@������x�,O�}�17ı,Og�g���Kı=��dMı,K���m9�q����ҿ���e�pR����%�b{>�=��"X�%��{z�7ı,N����Kı=���&��oq�������!XX����̖%�b{�ޤMı,K���m9ı,Og�����%�b{>�=��7���{��?7�C�ݓ�eP�̋͛�C�ܰpu���ېz���nF�d��7j���Fjۖ]L֤Mı,K���m9ı,Og�����%�b{>�=��"X�%��{z�7ı,N���3
hѣ.�����ND�,K��k"nȌ�1`%TgP��n&�X��}��ӑ,K�ｽH��bX�'{�p�r'�2�D7���}�Y�sA����{��7���=����"X�%���ޤMı,K���m9ı,N�^Չ��%��3����C�K#q�	��zy���b}���q,K��}�ND�,K������%���������"X�%�����k2k5�0���q,K��}�ND�,K������%�b{>�=��"X�%���ޤMı�#̿r���L"#m�" v��v؎�e�p��ke�Ͷs_N�I�K�kZ˙�-�Ѵ�Kı;�J��bX�'����iȖ%�b}���� NDȖ%��߿p�r%�bX���3�m�S����4��#�G�{��m9�1ș���oR&�X�%��߿p�r%�bX��ץM���TȖ'�5/��0��Kr�3S.jm9ı,O{��"n%�bX���iȖ?� ���Dx��M�����Sq,K��}w�m9ı,K�'��̆jLշ,���H��bX�'{�p�r%�bX����&�X�%�����r%�bX���ԉ��%�b|}���JhѬ�Z˙��ND�,K�>���Kİ�Y��6��bX�'���D�Kı>��iȖ%�b_|8�<~nm&�3ۑ��$u�/�k��/=������=�.,�kuZ6iJJ\Mı,K�O���Kı=�oR&�X�%��}�ND�,K�=뉸�%�bs�}O�5fe��f��SiȖ%�b{�ޤMı,K���6��bX�'�{�q,K�����m9ı,^��=�u���֌)njD�Kı>��iȖ%�bzg�q7ı,O}>ߦӑ,K�����4��#�G��>�� �9�֍�"X�%�����Kı=��~�ND�,K���"n%�`QuUK���6��bX�'��fz�0s�����y���#̼v�|9ı,O{�ԉ��%�b}�{�ӑ,K���z�n%�bX�{�y���p����pq���4aaLt�n�H�s�,�Y!6�H�нr�8�Im��ND�,K���"n%�bX�w���Kı=3޸��bX�'��o����b<�y��0�f8$�ԉ��%�b}�{�Ӑ��ș��3�뉸�%�b~���M�"X�%�[v����1b<��Ʊdd�ԍffkFӑ,K���z�n%�bX��}�M�"X�D!�2'�߷�q,K��߿p�r%�bX���jj��j��u��\Mı,K�O���Kı=�oR&�X�%��}�ND�,K�=뉸�%�b}�_��Y����h�SY���Kı=�oR&�X�%��}�ND�,K�=뉸�%�b{���6��bX�'ȳ�޵� -���^Z��I��GRX갂n��t>4�Qږ�2�ܚ���ӒY@GV�v5�m�˝6޳�+x��g5����"����op(#�y��Ƽ�{v�`�l�[�V�'$v���@mG�Ƌc����Du,%�+	2�W�	�]�Ԛ�̸��W���0�Y�D0��Q�Iw[�H��YL,ȷM����d��.�m��U�oT�ְƶ��[M�d��C���Yb�6�G�6Kttϔ�苶�uҚXjv;�����K���p�r%�bX���\Mı,K�O���Kı=�oR&�]�7����?�����ֆrw����X�%�����?�9"X��=��iȖ%�b~��z�7ı,O��p�r'�ʙ��{2���&h��Y���Z���bX�'�Oo��r%�bX����q,K�����"X�%�����Kı>��3���5���Y���Kı=�oR&�X�%��}�ND�,K�=뉸�%��I�?z{��ӑ,KĿ���j�!��5m�.��R&�X�%��}�ND�,K�=뉸�%�b{���6��bX�'���D�Kı9��ҙ����N17��%�gkg�9��p���;Գ�m˭lѹ��4«]�����K���z�n%�bX��}�M�"X�%��{z�7ı,O��p�r%��{���o���+G3�a����,K�O���8�DG"dK���"n%�bX���p�r%�bX�����<�y���{е(�2���Ab7��ʻq;�;���'9���x���g�@���R6F�r<��r-���ط x�Hط �_]���I�^e�U�>�w�Nr�7{��_��@��w4���ǒA�H��)\kc�fu.N��qj{C�r=���m��k3�i��j&�9��I�`�Z�R��m��7�+�XG�^�Wc�e��Y�k�N6�����ߖ����h��@��S@(u#�I�B8���srO}��ܨ�b2����E��9JhW�hpt�a1��m�&h��@��S@��Z�<�]߿{����lRD�R19�Š^�)�>Ÿ���g7 }�\��ͭ��I]k:�׺���'%�m�F뜮�v�聹��.KZ�]e��6�m��?������:�W+���n�4�j�0X+ň.�J�ߛ���r��Z��@�;V�ع+d�b��M�6�b��Hط ��T���w������tZW�*���r�w��'�g��rN��ٹ8�I�T�'�g�ff�{�ՠZ�<���S$�i�'ط ��T�[�=ש ���{���X��ۗ\�"�:9�-س��5�Fҝ��k�W=�{ltf��5�;\�&-f��YP�n �^��[�{��CɎ)�rf�y�Z�R��ڴ��sbG��7$m'%��m�?����>Ÿ���g7 �Xe��d$�8�4�h|�ր��w�*�ʮU��a�9�.#3Ȝy1`�Z�[��^v��)M�=�{�rN8�@� �D��t������@8յÉ��99�İn{]���6���'�P�Mz|
�]XĦ�=<�9p��nݎ���+����Ź5ۓ���Wݺ7-�,�Qm�w���"��i�/��w��"'�zV�i�-�+�<T:ݫ��v�cvlnmlu�% 1zl�zSFv3���R�<y�r���6�T����a�\�v;<o���}�]�~�.p6v���v�	T������{�����s����d�q���I��V��l <$���v��H?���;�-�
| ��j�-
\v\�Hط ��T��������ȰR-�)M�h}n�yڴ��tĦ,I�(]��n�,�����Ԁ>]\��1ēB�qh}n�y�Z�R��ڴ���C��"���ݨ����Ԁ>Ÿ���=�-s��&8`�юb�k�M�]Hވm�q��/�f�j:��QP�(9����2޾�{�2�?�h��"LDM�bN�ڷ��*;@^�@����ܓ�Ͻw$��]S@��\m�@��&,�@��w4Ϫ�;�Jh�j�;%]�2)�&5&h�U�wr��/�ՠ{���.]�7$�7&E�qhܢ@b��,����>�]�v��v����}�\S����l�m�U糸v�ͣ���#գK3p��`m�����7 ��* �sp�H �����D�M
Š{�����hܮ�~v�����8����_��]�>��훜4u�L�Wg��ȟ���z�'�!�p��Q���,:!:;&��erU��*���; 9��1!�a�⩰x�x������B� ���ا"�Ĉ�-����Q��0*ϣ��GK��U6.�|�6�@v�@���D�����ЃH`(X��H2 WF�[�|0؎�p�>��LV�H�$��U��$V} M.D���U����O"Ux���@6���6DG��<��8�)��ٯ�_]�;ｳr�U�9䍤�N'����h����7��ꪮr��N^���Yv�Y[�nU���@b��YP���^�)�r�͔�a1'�O�E1��oV�N,�`̜�-��n��ͥ���GLX9����h�U�wr���9\���%���̋1Y�+FZU {9�w^��-�>�ʀwe�X܌�ܙ	Šwr��/�ՠ{z�h�U�_�;1��1�N6�.�H�[�|�* �sp7�W�~��@8"U���}{�nI;$�����1ēB�qh}n�y�Z�Ws@�;V���ߙ���$N$�*اr����uǎy%1�O	v��l���M�<���A1�dpi93�?W-�+��?��ʪ�+��M��r�^$f$�.�⴯@}����W*��/@�d��s��s�ʻ'b�X��U���bW�P����{�* �sp�� �l�mHPE�}�����h�Jh�j�;$��2717ww�P���=ש }�pye@����߿�@6�C]3���3��z��L��ټqWQ����.�Q��곴� ^{mph��gF�FW�OS����t1�⇱Ƴr^��:���n]���v1���ű�˶܎�Nj(�{�/���Gs��۶�殻;��7>3%;�'�v�9omc�[ 7������Er��\�;bs�����m�)؞LWcKr��	��ԝ����1�����w������l�[)65
�;������n�������4��C��H"=J�-�]'�ߔ�4�h}n�Wuz}c�#x�ŉ��pI�@�;V����hwW�^�)���� �����2	4(G�����Wuz�Ws@�;V��wJ���G��4
����e@b��YP�nm�陻�e��ṹ {�� }�pye@/>�@>���R�4�1�H�yX��κ�q�iݳX���0�
���"4�Q�f��5"E&h�j�>�����ܮ�{z�na�D�,�@����@�H�H� xP><�Lm�Z[^�~v��_%�Ʀ(���Rf�y�Z[^�~v��n���QD�1��E2!H��rT�[�{�* �sp��Ħ,MƓ��f�~v����/>�@���4�y��W�1�b��� ��:S��e1��z97=8���h֭�t��HLmD�hP�/@��~��/>�@���h�j�=ϝ�1�1���ڀ=����� }�p�����b��i��R-�W��_�޻���E���!�"�w�f�|��-�|��C�1F�$s4��>�ʀ=���rT ��l��Ҳ����1+�?~ok@�F���m���/�ՠ^�:�7g�!�"�ɶ㔭����csۨ���L��tv��,t]�`�Ȉ��4Ϫ�/u{��ڴ~�s@�k���51@��МP��Pط ��* �s��z�ȱ)�j1�G3@�;V����hwW�^��4��I����m%͸�YP���=�J����������EA���~��|{>�2Y49��E�f�Wuz�s@�;V�����W+�%���.]f��,a�%�v7L��k��ݹ�����5!\���T�$������G����4�h~ojr�������u)Y����X��m@b��P���/9*~�s�����Kb˥��(į@��6����=�J�>ŸU���L�2H������z����Z������F�m��@��� {�<ʀ=�p�W����t����Ӻ��ޝ?w��q#�[���t��[��rƺG3egq+�C�����wA�G\��W��ج�-�z�u�2:p��W��<�9��a_n��mg��@�u0�8�Vv�>��Lq�S���mt����'c����2���S��k����[*.[��D����f��[ ���x�'P�@t�xr=���Բ툷.�ݳ�%l��Җ9I.I\�'d�v�W�
 ��v��t��&G.��R����Es���=M�.���Ѡ7F���,�y$X�����Ͽ���빠^v�ޯs@(Ř҉�&�Znm�>y� {��J�=�pq}h��G"�93@��Z�^�yڴ~�s@��ZI2G"��ma�� {�� {�ye@����e�O"X(D���/;V���T�[�ws��uѮ��Y����h�vv{&��BO��"͍�A\���;r]8)5���Ʋ7���Z�[��^v�����/;V�ؾU�0rG5�5-֍�=�{��A69��s�|}�fց9z�׵�w����m��@�����h^���j�/ܣ�"œ����[�y�T�[�{��P��85m���/u��/;V����4�ՠ}�*,li�0m�]7	q)����t/��g'Y ��f�f-��Cr�Y$�Ls$n6�f�yڴ�W��^v��]�޵lN��1�Vm���9* �-��T�[�_�k,y"H�h��@�}훝U�QS�kZ�~�w$��~͛�U�.6�Y���r-߭��/;V�{���/;V�ؾ���0�E$��ڀ=�p��P�n��T��w����>_�jη�jL�:D�8�kvE��z�'����[u��st�Y� ���p�Ф^����s@��Z�[��^v���<�,Y1���LQ��/5��YP�n �9*  {�k�M��Z�[��^v�����/;V��/��Ȥn6�$��hܮ�yڴ$���y�q,���,U!-
)�W��a�~�vh���'7�A�c�Šwr���n��T�[�w��+6�3�[�͝���.��u�zSq+�뜮���Őni2(�ơ��&A(D�L�/;T�,�ط ��e@re5���,ŕ�F%zߛ��U�Iznfցyڴ��m�9��) A)3@��p�rT�[�{�*�ۖ��%����,��Br��UVۙ�h�"�>����ڴ�Q�bɏĜB��*�?<n����O��	2߿w4ܓ�"�
��P�T_�"�
�U@U��UW�QT_�T_���A���P""$E `" DP ��T�DP���@, `�E `@�E b�T����E b DP
$ `�E `"1��DP ��P#���P�EP�@U�*�*�UW�*������"�
����*��*���H���EPz��*��b��L��n�x��Q� � ���fO� ��_ �@�J 	�bT  �  U@    	Px    �CAD
��U P %J� P  �@( Q(�  P �
QA@% �B��D�  P�j��R� l��JPX��J ��SF�� :q�.�)��X��-�W1˛}�� ������ü�x �X���̝�x�w7�V�|��;nZ�=��Mʋ;w�<�j�w�
 ��4  �pPT 
P ���B��r�ڗ�e����]���:��]���ӟa��ˢv�� ���n����X� ޾�罪�����*���U�=�{�{��x��xݵ� ;gϫ۽{�K/vF�j���:�|�
@*�P ��Ǿ�c�9�Í���e|-�!� �'ҝɯ�����N������s���8����|��m���u�� U�1o���0龌S���0L>��glns��M��o�o����P �( fG���v�}�;�n.�}�{{a��
w=��{����k��^��s� �z��j��>�|�����3� �=���x��ϼ�c�����v����}��p�n8���	 
((� �@���vk����ϻ���aﳞ�|���)]����4�h(�R�y� Δ�14�)c)� ���LM�9�3�)KM,f�SN��Nvt 9��� bh�i���"�Ll   =L��)J&�1O�I�6�J�4���z�Q���20D�*��QJ@  O�2T�ҩJ@  �h�IJ$�`❥K������s����g��N���kٹ��lޯ�IU]����
�TTQS�H���� ����"�
�QEO��	���c`P��7�l�C�ٴ��������J��tj7F}�MsXr�I?��+�� P�#
Mk���ݤ���O�>:�	r�7�1 ����f7Y�ؐ"����@����5�!"�ѳ�n�bZs�(�6�K,Y�\K�-��h���̼����w%�1�tbr|�hL�.1�ٓ~��n��%�L�s�!Bn��~aHXSLc�lH2�&�\>�}��_�|k�R��ĝ
�M��Z�؁AH$XD�A�F���Ԯ.����R 4����������7��ѯ���Q!�UӂB�u��﷮��&���7�1� ��5��)���t4G�Æͥ�m�39�8<>޼fp��7���2��{̮�m��G{��ċ�F5)
�t��\p��p��i!t�M��u�$�8wp޽:]��׷7�Nn].o5�0��2�,%��-�7�t�2X�ºe����+�X� �hN�,q4+��H��S_R��L�1֓{�к���H4��]��i��o|ֽ�v�;�a�\fE(�
�H�Eh1���js��w�����!��Z�w�R�].���p��ȡ İ�i��X0ԌX�-dԁ�R:J1 �1(h�i��Mjk$��7���*0XB�iČ
��رBFZ1���5����B)�4䮤�H�E!u'.��P�r�(KHj�ri��4i��)V�) B�h��i/	&f^�o�Rn�&Mk����Dm!!`գ&�H%M?' �M�Ζ�g0�!Ma�	~�}ی}�]7Z�]���J݃wV���5j(�.ZōB�1
'B�+�-�_�Y�X�>A���!I�Լ/�&�77�t/TT{_wRgݳ5xk�[�%�_�Y�� 9�SwD;̚v�b�[�Һ	uk��ɏ��χwл(c����?LGw�5����Ò�"@"�IgP��Fl���S�~�ǲ]eaXX�`���wDjh�5vJa�Ϥ&��@�����ޛ'й}y�x3������	]A�����t�@���JSF���}b6�%���i���ń"E�e��I��>�GP�:�9������u"0�c�]c.�n�#H�LH�E���L.;�1�6��&��Ҵ�E"��+�S��B��$'��j�� i��;u����{��Y�]B[�s�ץ"�,H|1�m�}��:��0�3����#%�rSI�i�Jġ�`�B`JHD�KIl���.��	$��o��s��9�q�l,�E���Λ��D��f}q�>Wa�m�I�ﾲ
$�x�E�w�(B�[�69�|u�����w�|��)	�,�-�@V5i�׉��H��x}�d5w��D���1}ϻ�Q ���[׿�����N�f�7tp��h\X�B
@M�+!�F	 �A�h:�l�������ks3S|�Ja���H6�X�{�K��|4����*$��P�0*(A* F�����2B0�~���Jo��
0��#R4	��#A�4���:��#�@�1��jX���o{6˚��Jo|هSX�!�^�|٣�&$���e��1ػϽ�!.�P�M�&�ϳ�p�͆������{IN��.�,m:t����$R,X,b�b@�!R׆�\6x���y�0�W�XP��$(���]i�l�6o��ΞBC(�>�L��D"���bEb�R�*K���BNe:�B���S���P�y�-�,��P��8�E�W_!�gO)�!6�e��0���(�H�4�`���>�����'y�ow�)��!��"Hg��~��F�	�HEH�"�H�"@b�t��=ϧ~�;/]e5�ۥ!�	C�v*����$A�@� ��#�c5���!���'��ӒbR�~��}��l`�`щ*@B%Q�^�
�(@(K�]��Ɯ!]�0�f�������%�>�p>�ßHB4)��9���o\��)	X�"HI�����K���n� ����oze��$M��7�}�!�k9���tB�&�$\8B�h��$c�*i�42�0ܓZ�O�'�1:�g7�o{ۜ:�|P�$#[�!1��*A�B5ad��!n�h�{�SL4|B�]X��(ʑ!F@"D�T�`�S�6˼�P䋓XP���C�(��;�ɮ��;�F`�� Q",7�c2c$�@]��h��VQ�H�Z�MeT�R-O����ox'�RBd'Z��$�1b@`tC!!$����l���$X�p��*Ab�Hă��8�LV�>Az2D
�aMK��3[�
��`fa��=�IIO�`�+
0a+���d����$��.J��Of(]���`�e���BV�k{��T�z���ɮ}����"q��D�V0 �aFY'oL;�SFr�.��~����Ā��]��bi͛6���!s5���o�Ѱ�9d!	"��!0$ H�e$``HS��XSY�$Ku�$'{��4V�p�EaZ�5"J�$3]��$�#��5:Yl��
1�2�\�7��fK5 �Q�߹�c#��Xք
$H�����vj�ϫ��n�W8��Ӝ�˾������I�ˬXД%1"��1M�X�"��)��U$X�M)���X+��`�FTҁ�B*D��"�IQV��D\ȇ�^"�H��[E��w����?�./��H��{˯�Es��n��h�9��L�)`ń	,�HHicaZ��ۉ�@�5�hH)�HH0B)(Q!(D�) @�H�21(Q"5hH0"Ԉt$�AB*� �F	�F�Q"�H�$B,b�H�b�H�j��F�R ��H$$F��	�t�l֢�e֋
�-R���P5�X$J$P����11��D#M	���l$R#�P�
,D�B��Lk� ��������:(b���IGY	��.�a+	R��RjC����.�Y!��F$)�� L�-���!
j�E�%�!� R���! �!	w�}�H&(Fta�}�t#~i��B@��}�zYIe�9����%�%��k}�w�e�meXMa�]f�n��t������K��>����v0�1a��f��,~J�_��n(�5$`�f�8t��!���c��]8�9ϰ�|�����B�3T���7Revp��L�;3'>J?atIlfk����]!"�r<��}k����e�1<��f8���>��X"�i䱒B2��Z0i
B�~:iQn�/:� ]aąj��.�E�H�CD7���Ѡ�XP�6q�@�"F$
�R���adw���J�HD���o���w�;��ϝ'۬.�V��-Z�]h�-XV�����M�(�ԍ��l                                                                 hz                                                                    �           �@                                                                  � rv�u�zpi���M���u���uk�7��&8
0z0ħ��Wm<ݺ .���['�Z��w�e�2�p�.���V�T�Y"�ŀ�� �[\�XԵmSk�Kр6���U�Yj��Y�KHG&g�U;bk�O�Z�����j\����<Mш�OHJ�kfr��'E*�.N���+X�@cb6�N�M9hܙ	��z]�\��]t��ƕn�gc3�T@d]���{4쪖@̇!D��*��&����v��Ir��I�[^H�� :�6�`�` lIam��Z�&��;m���ﭶH��&���v&�[]7`�o��3�Hf�dS�2�R�J:��YV�a  6�Xv�4��g[��:հ��Z�%�  H���^�}���m        6j� �8�n2	��6��$�o$$%���]T��UQ�U*�CWeQ�]mr@�6���'Ym6�&�H���}u��pl훐A��M�������AK�M	UU�eԹ@�<�^m�b���6yZP �ڀ���I��M�i�𥤀/��r:%UJ�T�՗�FU��#�h0#+��Uh-�Y�Zmm �5gm6�Y��(�U��/I�e��cm�� �i�vضZ�������(�r7HGm�H���-�v�	�i
�J�R۵R���Z�mlL�[qm-�  ���5�m� ��M�n�Cv։#�MoB]m[@e� pnBI%��qv��m  p Zl      ���%v��  @h��i��mHl@��f� �5*�YD��:v�X�cŻ�m�0oP �[�p  H m��`F����` Hp�u�P ��ж�il^� -�٤�K$����n�ݰ/]UJ�t������@(
�UUU �/1�n2�.��Z��U8m��#��ҫ̣�l���\� ��ref��ګh
U��vV\�h�ڀ	�U�D�w�w� ���e�R�`��^hF�Mn m���-�lq��ǒo�6����7,�A�r]f�Uo����M#e�������m�	q��lUX��� A�C���]��n��kX$B�ic��Y\� ��*�T�6��v�;e��e�v�   �m�lٻ6��ӅFq퓨몭��jn�.y�<���+0 �� [%4�a�l-�@�$�$	 	 	$J[A��  <�s���� � �`l    ��    ��@�`�   -��Ā� V��i�v۶�55 �ҭV����v�m�lm6�  ��  �m��   [@ pԍ��v��$���   h[Pְ�am   -� ���    		6� -�   kZ� 	[@�-� �˦�k��i0� ��m$G'#�u��jU�B����� 6�ڶںkn  �ݳ`�\݀  �d$   8ݶ�  ��?�8\�o�pm�,0�j�M�AVH�h��iJ N���.�s\��{g):���Q��#���PWk���m*`�8��H�$	ӂ���kY4��ye^ڪ���]J�����l�7kl�h� �۳���Z�/P mn�����k��:�+r��54$��i1�mR&�k%� �m�@ m� ,9���'` 
�a�����ݫd+[ K��� � �� ��     ��� 	   �]��/-��5��'@�d�m   	Mڶu���� stIv�� m�@ �i���UUU`%YUV������m��  �` �  �   �   ��  �  ��9��͗���v��i�\i� h@��6�  �����vH ֲF�L-�xm�� ����@     ��   6�L�m�I�l��`4�Eg��x����  	    Z���GZG  [Rdkit�v,�ۺj�T�XQ�ό|Z�R��_��|Saw�@ $f�6�����(�*����NZ���ήц������F��㷉S����l6�r��6ۧ/%� kY��e�MNζ�$8����g]w�6� ������/.P�v��cb�̈́��Il��,��Gk� [׵���8[I  6�D����=��[6[i���ʛ��l����Ă@ֶ�� rN&�dٜ ��WH   [@   $m�L [V�j��oו�c��-���u��m�M��I�  n�T�p�� l[�� p  8  m���        �    �oC�i��-�[m� @�� �   v�h �`�m�  m�sm&� 9%��ڥY�8�es�T6�6q�8H첀m��MWt����K�� �m��q#m� �n�  �   ���āއ�8     H  8    �	     �� p�        �    ���m��-��    @-�$ z�m�H � =��� 8ڶq�Ѷ�N�m%��oP���rm��ۄ���i0�m� !�V�T�t�6�|��n�D�$�-]Y�m�$��b@� � H6��m���ݒ p �  �`  �� -�  ���m��     	 �m  �m � 2m�$�m  �� ��  9�p�hiͶ�8�6�{��V���i�*�]U���:K��ipm�lɶӧ  	��|���4��
��MJ�����W�KvV��am8��m����� � �`�n��l:��v *�������Hj�N���YV-�6��m�F�m\���u�m5 �5��`^(�t�n�^5�� �m�]6jE��i6�m!� u�A�ccekHܜ Wh��Cj��&p9,��"��f�K{�$Hpm&�H  ��I��A��M���k�`6� $O` ӫv�*�ۜ\��k����Ӥ� ��ְ[]u\&��� N� ڶ�k�ר 6�),J�VUV���� g��5��͞����W�M�۲f�Ȑ�m��Z��|���SgR�a�=�X�c[\��T�VƦ���"�pU��YV � �J�j�{THMD��@���.$9�ZY|�kv�.�3�J�����(�'Al�d;���ۮ�)�32Pp� H��<-�#p/W6��p��B��TIi�m�$:�m	��f�$Ύ6��J�bDGK��q��.a� jm�I�-�Ͱ��Y�$�x���/�Y.�m�GI&�^t�6�X�g�Y�C���;�tU�K�S�R�=)�(��Xn��<�:*^�'OF7K���F�XQ5\�V���ګh�L9j4q�5�*�M�7M�t���N����,�y;Upl�Ah�4źij�� �黥m��m�$�T6i��H��ih	(�S�V��G�5o;�JE�N�wY	-�@ ��m�se�� .�t۱F^§��UZ���멉�@�e$���jmx&N�m�uʧ��gkK;s����m��{���m&��V���   /�ڇ]�S
�f� z�U�lQ��.��l[@ ,��oZݛ-Y{h0کvK�:B���PlO�B�CJ�C1F[m��SJ����  ������H �,�z�ݺJ�$�  �t��I�D� &�  ���  -��  � @[Cm�  �[�Ā ��К��n����T�lh���@:ۺm!�2ff��T� ���(�8�UT�A���' ?� �$E� l��x��O�Q�� PR��*�����] �h���C@h^�TW��D:� N����~U�Q����JT��P&*��_����� �S���@� ")�����u^�� >����T|���_ �Q��k��By5�`�cC��T�;E ���j��'Q�Bh*����v�	�J��*�����~D]��j| h؎�C¨ �@<h]
A1X��PM�Z�`�M��% � �C�B��|���DD�U����<��+Î�z�' _��*�� �$"	M��WP�<
?*'@~@��H���8*1��6��iH�XB���P�!�I�A�� ���DU�U��U@���� �WjDbC���
�<(A ���  D���,��y<�<���_��           ��      8      m� l           ���Cg8�p�c��p���z/;U�\�͑۴�Vg2[�lvXщ1�7-�i�v��ƺ闙!�=�� �O��/6��π�ˤF]UUUʁ�O%�h<豴�n��>t�K-nx�[�N/IĂNF	ɖnۜe��B\V�v;vH�3���%��3�3@m���ۍ�K(�g�$m��D�vGFk��N�����m�`� N0E�$E�EU월:֞����/]�ݧ�b(�Hu��-Q�N���Ǎ��L��b���E`MSZ�� u���%Q6g&eU�m���6�ԍ��[d�M�n�#��hUd�6Ba�f�j�j�<�=���9{k�Y�1�P:���N4��h\�\��m��n���U.��
.ck%����c����`�4��m`%ڀ��*�UU<�mG-\�:{e�r��̡qA5T���%ZU��km��69oF܊U>g�5�7F7]B��֬��l[���k�vْy�����=�
WD�m�)M���0ݪ�4��x�`���l�u���kj�Nێvԑc%�r!W��dk��@��Kp@�MJ��H�mm���YL��l��2�p� w(5�h&�;gq�49)0n��n�\PKWW4���H9��s��S��O$�:�Qܛt����C��eњ� K��l�n�� 7̷i�����â�X�v�x�\���f�Ә���؋9CD\�S����5��:�g ٴ�f��� �|���[����V%��vP+�+�t��q���s�FW�/;��iCX�v@�� �� � �[�e��t�:η70!Q�u��
qX0�+#<� �^ �5x�ahضѺ�ۤ%�O���o+� �*?'�TꮐH���*? �y'�C�C�؂�@�|�����������6��۶� 1���e��N��=�K���O+��U��۩�^�4�s��M�����$�M]l���ݧ`����x�U�J�왐�T�ר�+v�7	e8^�nyż�ѳ�g4�h[B���<m�(�v��kz��y8���ؤ��wE�:k;N�3�\��㋗]��`��mr�.CZ��̗Y,�گU��^����UP\eC��q�9^{r�=�g�c>������7b�c�bn��+�)#IAR��ű$D�ױ2	 ���m=ıV*�w%,)YJ�VRݝw��-�(��5��ӑ,KĿw^ʛ�bX�%�{��r%�bX?w���KĲ�ۻ��_��e+)p��F�h�r�r�5��7ı,K��ٴ�Kİ~﷉��%�bs���"X�%����XR������v����2Gr]���r%�bX?{���Kı9�{�ӑ,KĽ7ı,K��ٴ�Kİ{'�Y솮:�2�&fbn%�bX����iȖ%�b^�^ʛ�bX�%���m9ı,�씰�e+)YK�i$���z6����m;�{F^�q���ug���1(nt�e5�{{7]��c�֣C�b�N���~{���oq��K�k�T�Kı/~�iȖ%�`��oq,K���ND�,K>�����l���|��{��7�߻��r}b?+����ND�}϶bn%�bX��}�iȖ%�b^�^ʛ�bX�'���e��f�2f���ND�,K�{f&�X�%��w�6��bX�%�u쩸�%�b^��fӑ,K���=��Y�f[u����a���%�bs���!���j%�}�~ʛ�bX�%�}�6��bX��$1W}�+)YJ�^ٮ�sZp�Y�&k3�"X�%�{�{*n%�bX��wٴ�Kİ~�zbn%�bX��}�iȖ%�b~E����uV����1�ׁ���X�Ŷ�v맬����$��z�
J�j�3��̩Ȗ%�b_w߳iȖ%�`�����Kı9���ӑ,KĽ�.���e+)s�����h��r6���ND�,K�g�&�X�%��{�6��bX�%�u쩸�%�b^��L��Kʓ�L�b�w~�g���r)n����bX�'߽��ӑ,KĽ7ƀ<"� D"$ "�V� B��K��iȖ%�`�����Kı;��ۢ����2kE�a��Kı/{�eMı,K���6��bX���LMı,K��m9ı,K�}u�u�sR��Mj\̩��%�b^��fӑ,K���鉸�%�bs���"X�%���{.���e+)of�I$���"0C%F�m��k�{i.R�Y�=�c�(��ln�[�[g47:P�W���{��7��g�&�X�%��{�6��bX�%�u쩸�%�b^��ͧ"X�%����Kq��n]�G!)aJ�VR�9�{�Ӑ��GQ5ľ��eMı,K����ND�,K�g�&�YJ�VRݝw���#�0�8���+�bX��ײ��X�%�{��6��c�U!������bn%�bX�~����ߛ�oq���7������rqUSq,KĽ�}�ND�,K�g�&�X�%��{�6��bX(�!"*;x!��Ȝ�5�T�KĲ�9�5���;��rI��)YJ�,�����bX�'=�p�r%�bX��ײ��X�%�{��6��bX�y߿A�a�j�g-u����w<q<�=9�Y��%���"�m8�!	��y�.�f�bn%�bX����iȖ%�b^�^ʛ�bX�%�{��~A�D�K����17ı,N��z�����Y�d֋��iȖ%�b^�^ʛ�bX�%�{��r%�bX?{=17ı,N{���Kı/��׭֦d��$��s2��X�%�{��6��bX���LMı��D�O�~��iȖ%�b_{_���X�%��w�Y�r�\s5f�3iȖ%������17ı,O�~��iȖ%�b^�^ʛ�bX�%�{��r%�bX���5]����BR���e/�w�r%�bX��ײ��X�%�{��6��bX���LMı,K����  mm  d����t���l���V�ףM��ƇI����76X5��J�Wj��Y��8��j�ɍ���W Q\$�h�72k�����?��`+$��[y�kn�=������7<a@ݗ��ˌ�M:IR��ܲ�ݹ�t��r��[�{�g�ا9�k��J�5�䈍�:*n���5���K��q$�YFc��nB
�Q�C�k��`�|bC�B�s�ӂg��b�>}Qd�S2۵���n�����{��Ľ��eMı,K���m9ı,�����bX�'=�p�r%�b��ߧߒ�ڒI��Q�����ŉ{��6���GQ5����17ı,O�~��iȖ%�b^�^ʛ�bYJ�\�l��N4HH9NI2��+(�,�����bX�'=�p�r%�bX��ײ��X�%�{��6��b�n��G��ؽOKi�������D����ND�,K����7ı,K��ٴ�Kİ~�zbn%���e.>��v�m��չR��bX�%�u쩸�%�b^��ͧ"X�%����q,K���ND�+)YKʪ�U{s�$�I�K�r��.��b�kF��d������r9�c�\�OkQ�@��\침�~oq����}���m9ı,�����bX�'=�p�~Pg�5ı/���Sq,K�^�7�X��ʑ��K╔��b������ :����D�B
0`��k���߹�ND�,K���T�Kı/{�f�╔��e-klv�X�\%9c���%�bX����iȖ%�b^�^ʛ�bX�%�{��r%�bX?{=17)YJ�VRݝw���Kj0�8���,K? �D׽��Sq,Kľ��fӑ,K���鉸�%�bs�ߖR��e+)YK�or6�D���j�3*n%�bX���iȖ%�`�����Kı9�{�ӑ,KĽ��t��e+)YK���$�H[q�qZx��&N�GAԦ�a�k�9�<�گG,��WBm��BK�=�'[/������2 {ָ���=ƫ��Z�?������d ��p���{�����UM��c7qky =�\ �{�ʪTW%���4�9��Xݽ��n�%��t�� ����t�}����ݘ�wS���ʑ�� ����l��Z�wW �m{����y�n��Wb5�2su=['Gj��Y�5����/V¼�u�-z��������zG���GE��M4��S`�N�ޑ��ǀ{����d��Ǻ��oSԙ�� ;���] [f@z� ��vf�׺ō���t�}m� 9�ف���*��\�IVgs6`h���Rݩ��8`n�,�J�U�������=�� /um��lM�ڬ^��\#�ۙ8z�� ��2� !�qu��%�ܸ�pP��Ȱ�ݘ����t�}m� :����O%��t�� ����t�}m� =�\�:�g��'���n�WH�ِ޵��V\���Ğ��{��d�l��Z�wW ���E��M4��S`�N�ޑ�������w���ܓ���nI�V-'y�>��@  mm  d�#�<�rE-V���+v�8�+\�Aɸ�E�y��4�����đ�+�+���k���%���b%Bwn�iC�ӗ��Xk܋m;d ��'!�S���979�l�,����0[*��A(��d6;��v��s"�����<�e��.9iZy����v�nb�mL1d�������-�����|�? ���Y����wMBn�:��!�a����]Nx7V���iZx�����}8�] [f@z� ��vf��LX�n�WH�٘�H�wc�=���T�]6��Ǭ�}m� =�\ ����t�z�͵IF�M��Ui��zG��ޮ��� UVջ�^$��=5� ;���] [f@z� ��߿%�QBR���x���a��)�;]nMە�mV�1��-uu��\���.a8�&�l� �wq`9�?*T���ݜ���䯐˫i���ـ~�ed���BT�j"$u@_���7�f�'�x�0	��4�un�&��� �k��\ޮ��� ^V=��z���m����=�� ��2 {ָ�Ȼ�D�����m�=�� ��2 {ָ���<�R�n�I$�������ln7Z5�:	�qu�p�BI��6
�p��%�Z�tګi����� ��x����p�={fڤ�J��e���`�#�ݏ ����I���U]���]i�r�������9�L8�v�9}�n1M��f�*��k��4��8��y�����U�C�$F,&G\S�W���L�9��v���:'{��D#Bҭ(��BSB��ݔ�f���":��i��7���\��ba�$�tM:X��eFRT�)�beX$R%�^34GI,qO]��X͖�\Hx�l�cIFP�IF,�
U���Iu�R @�!��6RQ�H��$e@R�H"0P�VbP�RZ�i(J�(�(� ���D��\�X)�Y&�ՖS\!	9t�`�H�I���:A��>�]��~\6 ����X�b.ҥUI*�%�9�ŀ���7����(��)-�[�ʕ_{�|���� s���UR�J���~��_���7p�q��i��0�����N�{�{��>������j�ո�����plIp��y��+�ԒY�&ʓG��{U�M�m��< ݑ���]��{��_cI5Ct��بm� �������ό ��y�f쳖1[�Z�6ۀw~�2���޵���5]�jcZ�����^@>ݚ`9�0��������_%ԒK�����Y-!r�7�-U�� ��x��'/�n�e`�]0?n�4�&�fT��9��ٷZ�e��F��S�����rsry��;@r�£xlث��?�߮�[2��d ��p�뚍��Ԟ6�pM��l��ِ޵�ݏ �R�Q+eմ?���X{��W�����I��H�\i�ۤ��m�y =�\ ����� [f@>��{���S��pm���`�]���{�ŀ���9IWvl�  ��  6���Y�My��z�nB'��
���k��`�c�Meh[���m����������-)bU6�8�A�l��;��&���SVw[�C0l�r��p��qjݓׂ�Umv��dݱI��-��k.�Y��_����C�]�؞\�f\�ov��g�	n��vX�lF�M�11�ٞ.����w����u5���A�����J��e:�#[�.t6y���ɯ[F`p��k%��@�U_ͷ��e`��X�H�wc�=����4�]6��cN��L��.�w�����I��WfܲZB�ջ1*��`w�� wupzِ�� UV�+��-0-���rNx�vV�I���{�� �ԭ^}m]�nҢ�x�&V�U{��W����7g���Ni{]kSӔ�&�m[:�N��N�\���_���'g]L��.o8�_��we`�#�ݏ���Xn�e`��~�9$W-�RG s��*��5J����7� �}�Xۻ�?$���K�i&�m�hT6� I9���X}��]����w����1[�;�CxUU{�߫ ����zG��J��M��;��7�ƥ��i��`�L�������Bs�=�2�Ԓ��Oz6����m��Iv�-�vuiK����%Uݭ�Kwb�QqD7DS�R�̳-��In�A�nE��ߦ w���9���}a��ذ�T�߯����$,�H6��	%����ꫳw�+ ��e`�#�RI]���'n�;����r��;�{�9���sb��Z�E �E0ґE�"S���7$��O߳rO_[n�j�����%W���X���t��;������X��M6ڸ��H��sv`I%{��|{�b�>��,���I"�BK�+r<:Ll���ۂ�`i��Bv�����[Wb҃�m�ݐʪ7s#r5��#$����� ����?l�]U�~�7{��,�V�cdN�D$�9��?*��Sg}��, ���`zwfz�*�;��[��ԷM��X�vV {�<:���$'<���`���[[n)r�ڶ�ꪻ�}���`��,���IP���L""Q|/T��s���ܒ~����U���l�lM� �6<�w��~��� s�� �����zI$�]�N\W;�I�X.�uɄ�)q�h.{:1�G�7=�ۛ֞�%Wp���Q�#�8��ذ�0ޑ�߬	%��:���V˫j(2� ��4��/ԛ�ߦ {ǿLޓ+=vlQ^4�I�HN�6�0�ݘޝه�U�&�~ŀwߧ� �m�i6��i�m+��껐���{�vi��R_�ow��n��� ����D$�9�� �J��w߾�pw���ݘ �U+)%���$�I  ��-� P�����!���̜�]�.�)Q�����v�xJsg����۶�.����3��G=Rq��W�0�������w>n�&1���f	�N�M���Ԓx��Dh;������YY22��?��Ϛ� Gm�r�v�J��W����g����l�b^)�k-����v��\�t�;���w�{��vY������Թ�i���o4��G5�\�
�N͋����yo-ƥ�#$#�@��?�lx�l}�߬7{����Z�}iӷ�V�I��H�밐�������<���7��g����
�� 6��I��W��ߧ>0w���إ�Q�ˑ��`�J�=�߸����`9�0=T�RW{��`�������Y%�X�٦�%W����		� ����%�T�n�ҡ'I]�Z��J$�^-!�Z��D!��0Tk�7Zv?����3_i����p'�|���= �6<ޓ+����a�ό�/���Q��w-�I& w�vg�U�Z���(����b4�b+��:�<��z>0ޑ�U}Wf쾴���ؓ�[T1��n�e`�8a�}vn�< ���h��-���7hM��X��vq��� 7M���{�V��KV������T$� ��x\�������|�6�m��n�[f�4��h{a��+�\r��=���tQ�rn�C����-�.H+prO��J��ߧ�w{���?��X�� �D�v��m;��&�n��ߩ&����`��� ;ӻ3ʕ]��������B]�ŀs}<`9�0�I~IRT(�Z�WT�@
��� }�����7$����6u��܎\�Ki��CԒ����x!9���X_UU�vq�{��4�j\n!�wd�`zwfꪮ���~ӟ�H�^�m��n�n�'[��X�'���������H�d�gX���u��<���/-�R5-یw!$���Ź';��ܒ}����NZ������f�A������W_�fan�)�fjf�؃� � � � ����6 �*�����~͈<�������f�A��������E�A�A�A�Y뫫��L�殉�d؃� � � � ����؃� � � � �z{�lA�lA�D  j:������A�A�A�A����M�<�����^��l��"��nI����IU��Q�A����؃� � � � ����lA�lll~����y�D��B%t�� ~���A���;�y�d��k��3.feə��A�A�A�A�o�؃� � � ء� �A �s�lA�6667���͈<������f�A����%Z��F�rO�RF�˖�b����'1'C����iFY�wF��=ca�������޵�j�&.[32lA�666=�����A������f�A����޿�j�� � � � ����lA�lll{�=���k.e�tk332lA�lllo{��lA��z�͈<����{���A��������DlllW=��r�r��$�%_
������f�A�������b �b(� � ����6 �6667���6 �666=��p��3Z��.h�����A�A����������A�A�A�A￷�6 �6667���6 �66
��A_�O�ٱ�A�A�A�A��ں�ٙ��dɬ���d؃� � � � ����6 �666(�@׽���~������~�͈<����{���A����_1�@
��c��R?~�0�o4�q��y�Zt5у"da,�麘�.��:��d$	(Fl���YT0!U) �?k #��("�2B0���̬&�a �G��L0�#'	��Ҭ���0����d�$�L�SE�%I�)ZJ�Mp���E��F��]�H0��y�Ν�|����                    �     �l            �@����cì<���pv9K��trF��9�`͒Ŧ�ɇgTe�̦�*5��)絸9m��!�Ɔ�w�
��u���8Ɩy��^���jnCR�����Voey���8�p��ݛkq<��\/GI؜�n�:�m�s�b�)�$Y����[� �nٝ���V��R�AEu�A������FPB�����ڎx�j��cs
v�TV�=�8=��c�͌ob�K�Ӭ�6�;���u�ҡC]1�ئ�w��a.��'�X�-<�KV��l��M$� :ej�V��dk1�,�T�ml�Հ#�$�k5r��T�LYM8��4���mTUI Q��FӇ9;x;Mp��9���c����s�^�x�岰�
�@#` �c��X��j�YYT�H5���qĆL$��R�UT�O�{SԨ�@30f%Z���ʾX)��'
���3D�]�Z�z�� �k:�q�Rmۥ���\'g��݉`�����YN�͇���b�p��e%U�m��̴�]A�h��3m�l)@[V�U��n� �];���<���{10��.�g��Vδ٪��M�! ZR�5Q��5W[e�U3f$�n��籭s�=�B��49�ѽv����/5T��<�ά��9V��Yљ^�6眖��ݻ;L��L�Ĭ 񹆪�T@��;e��R�Z9Ӽi��.�ْ�nWM*[/������ۭ�=�z��ML�M;e��a�k��m�泭Xݻs�hL��E@��V���:�7>�uÓ���䶘�5����S���tm�0���!���LA�������vW�Ttn�[:�V ,׬fuۧ�E#V��wqe��ضѺ�ۤ%�Y谌N��{���������8������ yz��=W�:��@�(	�D��߾�  ��  ����k�����3�C���Yr=ۙ!E�DbgO�2�qWI��$�1x�2��Y(����e��v��j�N��-=�k]��Fzb�$@;;��1����mv���J�d�h0�N�V�V��PjiWT�Lc��)����6�Wn:�յۗ������Stk��r�tcWi�e{�;�����������UU��f(/Lq���ۗ��=Y.��吲���O.��Z���{�)��
�9�	�f���6667����b �`�`�`�}��ٱ�A�A�A�A�o�ڀr666?{��M�<����X�*����y�P� ���1RU�lllo�=�6 �#�*�PA�l}���M�<����o�lA�lllo{��lA�@�ɾR��rG!d�%_
��%V6=����y����A� �A�A���ٱ�A�A�A�A����؃� � � � �����~֮I�0�rٙ�b �`�`X ����6 �6667���6 �4����Bs��_U^�g��V؝��qE$��sv`UT��M��������mզ����D�#ݒ�<l`���ŀm�y#68#�tS�7������4�T���]���Bs�=���>��?R���%U���� �����H�r�ƈ90sf��v��%V�(� �T�I � ��O��ό �9���UUU]�����]�-9##��������T��$;��ό��6�M1��Cp��J��� n���9͚`~���U*����� =��[���.I��� ﾪ�w���l�� {�<�����yjs��'��7Onݤ��Rn��q�+*ڭ�g'Z�Q�\����u;�Ό�5V�r9>���s�4�sv~T�R��0=���`�~_��̅�VGd��7c�w�}�]��s�	:���pΪ����\�����i	Ӧ�w���	'{�����|:E?(�s������u���ƒj��鶮��o���~UUT�o�����~0����R�IRow������#DM�$�0ڴ`J��覆fC��s��q��������ʵ�R]���ۭ��l����p=/�R`���c��{����G��3k�M��cL����zG���꯫���>0_Y֐�4�Hn�	3 =�uW�a'_<w���NA}Ce4؄�m��|�z8a�]Ȼ� 7{�<�bl��i�˓�/�w�ߌ��^ s�فU�"0 !���E�����nI�O�����w.X��H`�ݼ�U%}��|'_<����l��m���c�ڶsf���q;�y�\��tu`$��5�xs��\��=��j�V؝��'N�M���� 7eǀ~�p�+�����t�ƒj��HL5'��ꫀ}�� ��T ����ʭٍ�7Z5=��n���uIxu]��� I�� ����n��v��f\���vs��q�z�@>Unn׺ǌm<� =�ـ*��}~���x�;׻xU)]�|}��   -�:@  �uۖrt%�m��6�f�Ԩ%ܩ8��q���j�%fe�dٱj8�g�\���֏0�2�S�r@>�U��j�uG'n�lEr��w%��w[g�-0X��J3A�b��U��㱇s�M�*�xzt ju�A.�ԁ�vp�^m��̱�V�K�[��i��]n�[Q�֜S�X�Gw����w�伵MJ���q�j�r�ֻ/�jzGh8�-�����3A4�(�F�]5��M������� �RZ�����u5�X�{��kM�>�t�wm� {�\ Ys�Uј�M��ݶ��up���z�@=W���v�:t�n�?ʫ��� $��~�p���}׀{��4�T7#�D;����of�UK������;����������t�m��$��]F Kv��k$��Q�]nl�խq[�l]u�$u���fe�o�K��ƈ�O��}<`�������`I�� ����۫�%�I�w�4̪ԩO*����& {޿L�l�?RI~J�;��m7�7	RG�0wߦ w�{0�U]�0�Oݽ�6���p�&�Ԓo�����?{�L*���}0�]µm���M1�o ���n��up����cm��{��l��+`I�{u��q<�K�+{i�4�5��sm|c����?*E�0��A]ˊ�I!�=����ǀ���������%|�셵M9!��vg�R�J�a�~�� �����٦z�%vs�~�ۍ���qɀ��L�l�UJ��(��U+H�)G�?|��~�>��O{ޘ9��o!#�-��ܘUJ��{8�$�� {�}UU�]��� ��ߋ�"2F�p�{�L�UUI_{�� n��0��L�Io��KX��Ƶt��3���ѧZ�Q��8���=��cK�{$�����X��6G�:l��I�� w�{0��Oԕ%U��琉 �_���+�G �r`{��<�U*Wg;�� ����vg�T�*��M��^��܎�$j�P���;��� �vi�W�}��f��u��%� �heݴ��6ف�UU���� n�x�.<��J��*�K��� ޻5�������m����uU�>�t�wvi�~�K���m8��K��!l��2���:��)�tl^5���ƭ���\A٭����q�2B�\rp����6i�n�/�����X���/�,cT66��h���>��3�T�Wf��� ;����of~J�K�I6wÿ��7.�#Q�G��^ s�ه�*UI]�u��=���?\�Z��J�1�N���u}U�}_]��x'_<�����P��E���=l�X���Up$�R���<|��� 9���IQ��Ϡ  m �� #�5��vM{%��؈��Na����tKU�k�s��"E���i	�3Oa��P�k���檮�ˠ� ��<)9�[�;UK�t����Hl:m��3�S�\���Ӈl�g��6݅���whb��"dy�u5$�x��9A�x'F^;Iݩ��gmZ��+���ۇK�Ό�۝�`Í��1�m��_�_*��^�F.�g��F�;����:�Ocs΃f��Ʈ{m[�?��w����"RZ��ڊ����?z�o 9���%I%������=z{�n2q��I�{��J��Wa���%���~�� �}<`�g[���A�(�nK�s�0��ه�R��w������>���mƈ��,��������N�x����?%IW�T����n��[�.4HH��T5m��0�����_��� >|�~��~��~���,��:�E����\����P��n�N�]��bw��d���7t�cL�7T���ǀ���J���}<`�Y�v;�m�K�!�xI>����|�TdH�����X@�XBH��H@'N��KS���!��V�}�_&�~�0���y%Uv����1&4؄�M��|�ގ}T��U*M������~���m��{����p�] �j��W�R����� �����]ȤnH`�� ���vs�'_<����~������KSa7X�km��p���w\!<D�.���v^?�����|S��Ht�Rm��7g< ݗ��ê�W���0{o�q�1�H\r`{�� ��4�;ݚ`9ݙ�U~J�l�����\h��n�Dw&��?��znh��!	P��H� ��Ґ I4�t�"�,"��/�hC�e4Q]��h���&�$��<C�1d6�!��VU`P�	RV%�"��$e�%�t��wJmhi@�%!0vm�VT% �-%Ii��HR)J����GaB3G�	���:�+��D�1�2�H!�%�J� F$#�"
B�F� �
Ŋ,
Ɖ�ƀ�jK�Ab0�J���
��B���D)*�,�i(���Rj���Ж�fL���&ʵ8���h������<U���+�}��@�8���U'�UIK�Us���L ���`tz��Ę]&�Li�UUrvq��� wU\�WHʢ�F���3Sׂ�`���_U\�|�����0�������.u���h�[׵��}ƪ�s[X$fi��c�rlM����O����D�&�ܟ n��0��L�٧�I/ˌ�~�����w��$$�0�] �� {�\ �1#�p�he�t��[l�$�� {����&�{���w��`׮�;���;$�0:��vs�	:���0?U%�U$R}����v�#n4F1�,��o 7eǀuW����Iό ��?d��wy�}�� .+y�9+X�3�J��큻cZ�fy*���]�% ��ݨ�?*�Dd�w#�8w��`��0�������|�Ar��m6]&�Li��p�{c��q��3���_Y֩.-�e+���3 7g< ݗ_}w���"� �r�	J�V�e$ě�ꪫ�:���|`�K��W /�V�^jz��[ci��G��G��7g< ݗ����߿���   m�h  &����Бm�;y�ع4c���ݳB�[]k�{b�F[�ԍ�P�b�����z$L�v�n$kH]��W�k9Y�>��PK[����$��m�4��s:��ջ��sֻaLfKK��&��v�JG�YrL��r�5�ƣX�
�'����s��s'\��n��;]���#]�ˊ;�7���o?R�U�W�s��m_�z����&�]�[��u��t����19�tg�tu�M�#�;���_��W$������/���{c��q��0Eƚv��v:I7x�ly���I�� ��� �R^w�]��}�$�p�Yqɀ��L�l��I*��&������L����DRKc�#��ގ�����:���������+�K���#�޽��<�}{���	:���0���m��L�:�1��N�ܩ�=Y��8�r{1����CN������;�r��m���߷���ގ_}U��E�x:�Uiy]��A7���ofb�U�T,K*���I�^��K�}<`��^ s�� /�V�^jz�z�M�>�t�n�/�����7g< ���.��(�]ȝ�.�!���UI'�g��� s�\�UUssL�~w��r��<��� ����Up�] �~�d������3k{BpG��K�0�uΪ�� �ع�#��S�������>J�N��[M� ������ �R_�$����L����c��IlpDi�ޮ��@{���W?fg�g��Z�ۻ���&4�E�x���nkpD��~E_¿}#����|`�Y-RUt�M�I� {� nˏ ����_\���u���M�RLI� ݗ�}����.��zG�:��}#iRM�G<Lry93���Huz�)�;6�ڛ�C1��Fz9;�Й�&'5j+�m����`�K�zG�U~�$��u��4�'m'bv�m����w���|�z8`�+��v��v:I7x�H�v\xu]��� �w^�m�i&�hCc��m��������� ��T����k�{ܪ��{��l��Cv��G�}��w����n�ۦ�bI��4�;�����F�"����dl���3۞���2CqT�9Q�G�{������og�K���������^���;r��ݙ�UT��7}~�{�� �^�窫��u���6؄�m��|�z�@;�� =�\ ��Z�y���$$�0=�����{����sv`~��N�x^��I�v�S�퉶`���UU_{�O�=�L�٦�UP,�M��S@ﳙ����  -�-�  -�?���i0�(I���`M��*��g�r�T������X`oW3=;7'�lj�8c�tAd�%��l�.'/We2-M�zS�c ]���i���7nN�N�6u��4[*����U@j����ͱ{B�{]F�Gnx�g���Ʀ�����Clkkm�7k�\f��)벢WBۊ�n�%��)/,��$�I"y��j��j�ڪrj��^*NyӺz�o��6x7Ⱥ�ɴ\�Fa�J����6������yW ������ו�V���FƄ&ۀ��WH���H���$��X�����e[xw���y^� =�\ ��pq��,M�����cL���Ӗ n�< �����$���{���`��~��_�rEm��� {ָo*��t�y^���>���S%SR�7l�<��V'&�,��"Zf�oS6�!ּF��/ﴐ�6!��&[o�t�x�0\ؿ�������L ��?[���9q�HIr`��0�J�Ki$�������� �n<��볯N��t��T�1��`}9`�#����;���7y�z+;o\�.[$Nܑ�~�����z`�_<ގ�UU��� �K�j�T6'nݖ[m��q����g���� ����$���$�I%�M�1�0�`���<�J<WYC.��9e��wh�����vIyo!#DR(��ܟ�zx�9{�`���yW �����m�M�T�cL�=sbΪ��%�� ;���>ݚg�Uvr�g����9"��;r<ow� 7{{0��(UIm���UIfw���%����-Km�1��+v���������=���=sb�6�b�ބ�bt��m	�7m��p�;�����V��o*��cm��In&��&NN1Gy7�FN�^�<��q�;Ǯ~|�ƞ���?R��a�de�P��o��<�u�o*�Z� ��rۭ6���v� �����K����_�w������+���޶ı&� n��`n�0���7��ߞ���<���y��Qۂ#�0=T���x�;~�<�����E
�i%]���f�L���Ա���iSm�3 �͋ ���ԕz{ߟ ?~���۳L��ci�C��7ZzBxY�����;��.'�7������/����s���3�\��ꑧ���݋ $ۏ �#�U}�����u���p�A6Kq��ofz�U]��������svg�J�Wa����N�vЛcv��ό�6,?�ﾻ7{� wK�K� �h�I��f�z� ��p�U�=�� ��r��V���Zm� ��x&�x��znI��}��8�b�#�"���������� C��9|��M�������+��;QĀ �AF��D1��a
Z#�eN} �"�B,VA�����lV	�
�&(��F�B�E��m��6�a��!�B��T����P��B����I$�H                        6�               -�[]l�c�#8^ъf5�Nv�*��rz�ۛڻB�q��nz�#Ӌ��o\��n�b ���T�Ӹ�J!ˋ�n;P+g{6�UUT94��L���s���������N��fx^X��p��8
۫����YJw`�09��ijB��)�F;2�`kn e$Tk�E͜���2��5�,r����ݽ���q��>�X�9�cW]�YW1\E��XG4*ؽ㮻c���w9��a˭�ζ��z�XM6%�ݖI�l�mfL��j�TԪ�-Sm��m�m��zXjL2�j�P��jj��lU��UO+�R����9�R���`�m��%�j��PIt���v�6��:ۧY���<�	�YmVܺ��/]3�G!s�1*��[�瘟*�@��Vʲ��廕k��v�!̅f��p�`��bҒU�=F*������PM�e���I�l��X�ing�G4��y$��z���s�������+����5U酳�	mv���
�,���p]uu�nm���Ґ+��	V��������d&�j�C��6\�ʺN�]s����n�&�������b[�����Am�m���uf��ԝP�<�#�l�q���/=�mAKKS�;���*����KՌ[]x�s�fA;$r��`���۶M2��d�m�	[;d��p�-�W��6M`ط4-Ϻ��r��:�:%4+�q/��@�X��,��6�綶��hڛ�|b6OZ�v�<nvd��)�k����b��;��=��Q�v�c9+:�\�M˶��C�՝�`�;]r���7`y�ݕܝ����Яl7�E�
��ݹ�E+JA��W�a1�3��n;l즩k��n�@v��n�QO��`������ ��~��S���^�Z���bEZ.;��ٙ�������� ���   �vb�����@�u����ºE���i��fa�*xxz�z�K��չ2%��۰�S6��-)DD�OA6l��5K�Vs��ʽ��O���%ɪ���մ݂��R�Vֹ̛i�-�Hm��@���kjv[e�Sf�;���n��]�Yͱ��uļ�תc,/M�K!�3Xk5�_*�V(��9�֍k33Y�5���1�׃��5(Nv�6�m]sa�fĝ�Gd2*,�x�D����߿�O���p�=sb����`n�<N���Mbx�=Z����t�y^� =�^ n��g�%UJ������˒�܍�#f�Ӗ {�< �n<ގʢ�A[����ޭo`�k���WH���.�m�X�fn�[p�U�=�� �v {ֿd��7ߠ۝�+���-� �Gp���¥�g�e�ͫzw7&8�zą�3rLHM��o ���� {�>�����/��]�\Ս�V�X�0\�yuZ*R����f n���9͚`�+��ch�c�趚�zG�j��WH���+���Zi�$�p�U�=�� �v {ָuUlz��o��ޮ�+�`�k���s�����2�t���6�vBW<Yxeg�5��7b'Xs�n��ف�)�5��ͷ������H�M��ꪯ����=}gZ���-��G� s��<�RWa�m�`���=sb��Eli��RLrL ����9͚a
_RKR�*����k�z�j5�5���6��p�6�ŀ����︜��:��v4؆�m��ذޑ��ǀ{�� �64�&�դ!�XM���m�NY-�ь�g�:�I/b ��cn���(�MD�=:�������߷Ͷ����t�r�v��c���zkN�wv�x!��}Uvn�� �Ӗ {�<v\��[T�7N�j�&�z�@9^� =�\ ���\�ݩ�˴�Lm	3����.��w��I�N�7'�~�Fd'�`IC�� b��[!X�X�`FF@ DHI0�����ݛ�r�g�4y�b�Ҧ����zG��GH+�`���m��[�`��7s\�v[m]�#�J�l�X4�
��b�шb�M6���fn�[p�U�=�� �, ��x�BZ�4Zh&����G���_w,?}Wf�s���R���^=OP� �� =�\ ���=�� �UO[i��I<y�[��Z����WH+n�>��z��OMi�	� --psf�ow^ s�� �_uQI#w�   ��-�  ]I�5ݬn�˧[+���.we�X&�4�Nz�]����mFR�a�#�\k3��r����J��1�Bn�t*+���M�-�ցh�FvU�l���F�v��K�E]�]��$��T[�\���<�:5.) Ü�^'^�YUǘ�R68�4���]&ޕ���m�YtsFMt�1�)[r�����UU��Ě�7=��n��šm������%{g�]���;j�ջ8�ٺ&?$�>}}���m��Z����ʭۏ[i6�	!&`rE�� HH��p����_Y,T��-]4դ� oNx!#��}w�06� =�jV��$�В`���=�p�6� =�\ ��V�^��1-z�6��t�r�� ��p�� �m{����=S�&\��\[s��O\Ge�aMi��r<]^����*�ZMp�j�������_�� $$x�0�+�&յi��'nG����$�UQ.�V�����ގܑg���]��}�[j��m��V6� w� ����$X�n���׎\i�"��Mr`yU}U���q�K��� $$x�nZR�mݶ�chI��ذޑ����{�� }�m���u9<1���ܩ�=qqm�0�x�Cvh6&��5�$4njoE�Տ^�o`�k���WH���.׭�m6ٚ��x&�y�}��Uvn�� ��� =�\ �ԫV���[Ե�M�=��7$�����Tە5�����}� ~��\�U�^����SHm��lX�H�M��;ﾫ��� �\��M�j�'wn��� {�< �Upz�@<�]�|�km��x�[���]��t�97*�붧k����㧘O3�����Z��h{$�~��^�?}] W��z� ��ѽ��u��Spz�@<�]��� [ʸ�*�n=m�޽c�7Y �v {ָo*��t�|�*75W�LE4զ� {�< �n<ގJ��A\I!UI)������9-7m�RLM� ��������?/�, ��xݘҤ�v��e�e+�c�|�ݴ�t"N��̶�ycG=���r�5j{�5�K^����] �]��� Zup
�V�z�oM!�@9^� =�\ ����t�uڮ4�Vն��t�&�ޑ��ǀ{�����ו�S{��Z�4Ҷ��	� ����6,�����x�|���I;n�(bo �������sv`�ݘI%N���@�*"ET1_�~�  ��  ��M��Ʃ���A���ԕn8[<��ue[��f��t�;L�&�r�-k���V�cL=X��Z�
;u��x��=�.T..Q+Ih��V��լ�Ī�b��]@�k�@&<C;5:�؍�/@��ۜ���'g�w$v�9ct�@3x�:�^Kosk��.5���<�&v\�EH�!n[5v�Uj����]�eVѴ�ztY�x�,��k�l[�x��Skc;i���!n*���L�8
���z� -:��] )fڰ��T��MZm`�#�	��WH+�`T]�[Z����bm�N��WH+�`�k�z�j��Vn�KZcpz�@9^� =�\ ���e���Bo�!�@9^� =�\ ����t�I����@���dt�sv�*'C�KVBDh����&���E����l���2�R�0'M������Cc�=��mλ ���׸3V�Z�M����b|[ u]��s&w��ܓ���[ �6<v\X���vݤP����H+n��W --pUU�q6�Z��7��d��`׫��<}��Y���:iS�V�X�lx��_U���c� ے,�������%2S4�5l��=;�k��+���Ş!u��ֺ^��`y��%T�Rݱ�i���s�7��m�}���9����j�WI5v����}��V݀^� ZZ�Yi�n�X��5!�@9[v }z�\�_ݟ�$�F4P7�6�1�����0HXX��*j�<Db���7F@��ډjQ�5��*�O�QѤѡ�YE ��J�]@��B���h_��P�
�hiƂ&ڒ4A �t��F*A� �@%E�	���4��V6�Q�B0��Z!E���M(:E:� W�yU��ǁ'R�������v`sf�u٭���N�:N�M���ǀ<}��V݀}yX�7����M������H+n�z� �����]�f�f�X�*sJQ�ˎ]X�[S�)2�'\�&s=�
Uݭ7 �����`�k����^�{d�ݸ�R;���מ��Wa�����x�0\�m!AӴ�c׫[��Z����WH]�@���z�[i���ۀ��9�L��o�U���B}�iVg8�}	jմ��4$���=�� �] �k����m�x��Æ	��ڂ:�	pO\�N���p�'?����{.�M��[2DJ'�����޵�N��WM�$��v���浸�^6���IwXȒIZZ���G�ww����*��m�}���X!����l�$������KʺlI%��}�I.�IwUw�5�u&������IyWM�$����$��������~~ ~�O�ROTgY�$�^���]�2$�V�_�$����[���7zh �*Q��R	R�(� 1��`�Q%�g�s}��   [@u�  �k��]��Y��ܛ^)5@�Kyy�-H�"\u�2�tޔ�6;;oqHc
�l�5��4U!;�&��\*�̧��7U˙啐IC����,��gvyƻb��b6��V�v�m!��%ɻ<�'C��:�+A逐<�:�{ٙn�vn3��SGV��nzu�/X\���-��2����w|o���ͤ�@I��;�'=1��F��O;��݂�gu�;���2.mt,z%h�� :�ȒIZu|�^U�fg۩+����� ?�����Z�:�վ ߻�����Iu}W�$�$����"Jp�Y���� �o�� ~��e��}�$���3����q9��ww$��%��1�[6$�����I%�c"I%i���IyWM�$��v���浸�^6�k�K��$��������\�?�������� �~�e�h�(F6��s���N%�����^��EWR��5�1��l�$����Kʺn]���%��}�+��;�ww'_/�MS���6�!$�뻾^�j��$�J�n��!l^�����9��T���D�J����%��V�������m�u�Iuv��I%�c"I%ik�� �o�� ��7ۥc�+G�$�g���dI$�~?~|�^U�bI.������ O�ڤZ�:�վ ���KʺlI%��}�I.�I~|}� m��Z�cv"im��8��c�ce����E�\���Q�U&��r��k|�^U�bI.�S�IwXȒIZZ��$��hֽn<c�lI%��}�I.�I+K_�$��tؒK��U��mf�ZI���}�I.�-��z{��^�O��������I^�O�I/Z�V�ưC�4�m�$�����IyWM�$��O�I%�c� �ߧ����*VU�j�? ?��.������w�=뻻��̻�������~�j�����m��t�v;T�+�*�n��n����z�pۛ:�4�3KQ�6��lI%�e>�$�[I+ů�K��$/mG-�ܯ4�f1jm�|�K���$�����%�؈�K�ϻ�� >���dZ�:�U� ��k����DI%��}�I.�2$�_z�֧��ך�����$�Wb"I.�ߧ9m����n�� ����GIa-Q�T��`ԀFTF�i �\��[�����֧�LZ�h��x�'�$�[)��$���www!#����c�f]��UW�s��$��b�m�9�ѭ���[���z���Web�4݃ukt�[�;]r�������I+K_�$�Wb"I.�S�K���z;�D�[� }����? ?k�$�Wj��]ld���������4՚�[�,�ݑ$���"$���R$��tdI$�R���%�Ȼ�5�O[��m���$���_|�K���$����K��$����M��F��f�����$��ȒIZZ��$��Iu��|����>���   �   �65�r̡ԯjY��Ed�R{5&'��ֱ�Cat6�l��ӧ=.����%le�mz���]g�[��5���Gf�Ru���Й��q�ػ=a�+�Ã�k�bx� �VsI�6�a�s9�z��z�:�W-�g�9g�8�������ڟ�ǘz��b�Ut��Y��̌�kr��������)�)���n�:[�$�v����L�sF�i^�*�wX�Z�5S"�Mu9��$�V�_�$�Wb ��] u� �UT֧��kĞ����l�Z� �[2 ZZ�t�5���lcא���d ���=��Xu����r��n�0=IR�������x�L�����?H��{�a�F4�o x���f@?n̬�&V�UU�'6�m�V��WYw4X�S�����DM��',�Qu[��]��L�+i�5CB�ƒ����l���?oY�u� x����ݘ޷��{��z�@>�"���<l��� ;�f����>������RJ�j� �ɕ��G�U���d|`�d���z��6��@�k�{�� �s���l�yUS�O��z�6��f@=�� �[2 w�\�R�{��6��Wq�n��(
l���Q�,p�@mf�G�<-׫P4���|�o�������-�^w?� �ɕ��G�{d��6(�4�C�6�f�+ ;Ů�d�ΐ�zW�^�X(�K��, �ـs����"I-&@�*��]9�f}7$�훁�;z�4F;���AɁ���+���d���ِ�Z���ݘ޴�{��׺�@=�� �[2 w�\�l����m��{�4�$�vcvםѺ�ѵŻ^���"&�x;J�qz*��r�Lm�3w�@=�̀�� �[2��H�E�ך��m�m����vg�URJ���ذ��;��<�UWa���}n�]�Wn�,m�;��w:@=�̀�� �Q�O����אw:@=�̀��d�FB$*U	X� 2��
��*I��w� ޽w������d�l��-pu� �g�O�ߟ} :�h6���`^w3k2�u���G2 4�W��u����,�fz�cэ$���-pu� �t�{d��?{n,Bj��Ӷ�����������L� ��-,dp�%����{4�9��Xz�J�Nx���,�HJ4Sn��I� �f@���=�́�����Y˭6$��6��`���l�7$�{���}�}�rMTqMA�x�&�Z������b�����"��H�E�L"���'�$�: ����Bh!I�h��#(��	�t�ܤ�M��Ҿ4qH��D�����(!Ī�ʭ�Wo�Q����A4�P%juP��s��l��h��ԑf�!�)�06�� �0y�рҍ��u��Ԅ�͟�=�                   �     �               �rs��h\�������B�\X0��u� �6��	�%��u�k��6�����\m�ztU$l�Vysn�vsv�6l4�ԸH�sfk4ȸ �tIe�̺��l�ey�8� 
�<$dhi��R�7^�$%��6^�������&;	=NO`D��X������)!<��Z���kT�A�������z�\��e�M�
tYA݋ϗke��	xt ݲ�/pn�l�m���l��q���묕S�6�,�N�T���-%lR�Dt;m%�I�m�lH�V	&#Z��+��UT���	V�*�
� *�����H�9&
S���� �H܅F�g�UQ���e݁���:�K��V��N�lX:��gm�p�6�1*�h:���i`yj�`%e`ཹ�S\	"Z�z]��Ұ6�
��Z���Pu 0촒٩'�EUC��prσ�fUY	�q�h��f�h�܌��=�.�X�>7Z��]u��Y�ħe�M�d���ppF٪s����Jd�k��l �-��$�:A��U��ِ'��6䜻�Nwl�k3;Y��4�e@%��Uu@TJ��r������[��j���'����q2��m�Rқew+�KP�ڴ9��䲤t��G2�)�,1�ZH��I��Ֆvz2[�l�im�Z�gI����eh�ɱ�v��T���v��I����>��R�	�:q�v���8�\�ِ�m��z3���<vw*�q��}��,is�l�#)m�lN�QM������a����n-Vj9yќ.����Rrv<\2�V�9d4v�K`@
��ٹZ���h&t�l^B�c���{X'���&�4�i%8�Uv�A��.��Y����"��S�۾��
�p�U�	ر�"�T߄A��E
p���@  m�[@  Y-�%t��\�1�M�D���Y��N�����i�v�����O5e3���U��K�Jurֳ��5m���e�K�D����E�΄�5$6�;tW<�N�ۃ�^��}xk�@�;7h�PQJ�NS�UU�M
���1�ʽ\Z#��:��Rk��hM�	t�4��R��L�Tb�c��nZ)}IR˙��܅�s�u�={�:-�<N#,]�Y�7���i���Q"����k�m����+ ���{�2�����4���w�<f�'� w:@=� x��ޓ+ ص\i&�bH*n�0{fV o������ݕ�zG��F��mSTRC�M� o�� ��3 w:@=� {�٦���Z{��6�ޓ+ ��&q���X�{�0*I{w=$�I"vڸԷw��c���ƴc
2���c]������kc[b�����pz�z���y������d ����_Xs��,��567��$J6��nI����� N�(�3$ﹼܓ�{� � U*׃׏[x���@�� ��̀{�̀{�f@ʣUO��kZM�޶d��d��2 }ָ���k��OLO^@=�2���g~���� ��2��� 6r8k#���ݹ���8�IN�@Ɋ��7�3�iׇ]��$�gu�ў�n��;+ ?l� ��2��������X��9��C����n����޶d��d��2��]�k����m�nL�n��9��,3�UuT��R����J��ss w{� �v���F��r�$nE��T�%|��� �wذ��x�I��z�I	GHI�;T�u ��̀���� ��� �Z�*P�S .�lյ�(4��LM`��ٺ����qֺ��B������+ ���}�f@>�f@=� �;ۊ�ۊ�[�nL�n��UR�vs}�X�� ��x�$�Hi]�m1=y ��� ��̀���� ص\i&�bHv*m�X��+ =��7$�������_@��o=��ܓޯJ�[��Y�1���@wW ��̀}�̀{�f@>��m�m��o5Zs�a}�׭%�뫬�6tCi�,�^6��27q�8�r��ڗ$�>��,�� ��̀�����Ǹ=i�����ɕ�Uvn�������b�9{gX��D��܋ �;�����>�� u� ]t�ջ��oz����>�� � ~]��� ?U��'�R׉5�&��[2��2�u� >�\����[m��  [@[@  U�����ՌM�1��5.v΃h�
�0Y���ۖ�0�@V+ua�;VF��&�UYy���َ�[�]��gp�mЯ+��/6V�>�C��� �o%lk���t'`���q��S��k�bS�p8�[J�.����.�f8��F�͒��5�0��֕ͳhwni�;u�.�dA�.ιgM��w�o} [w!�erةݝ���H����u�ͷ'?���1�Ie�2B[�㻸��\qp���wq`�k�}�f@:�6����{��n6����2 }ָ޶d�Γ�ff]��h�i;���;��� ��x�[2��H��d�r�4׸<m��n�Z��[2��H��d ��p�UnƓCѦ���o �t�s��X�wf�7q`J��}=��nL�N�rA.�V��\��nzv���vz.k��h�n��{&���s]��6��ݝ���G�~��]_�6G��9	]�6ڗ$RGr, ���%*T$�M� ��)����ٹ'���ܓ��� ��5T�jZ�&����>�� �\0꯮�ge`��z"A�&�=LO^@>�t�{�f@���}�2��E���J݉�f�l�����}�f@>�t�U�w7[׮�X�ci�=���F=Y��,lW��ݺ��2*����Z���ߟ��o�}�f@>�t�{�f@>�+�M{�ǭ���4ۀ}�f@>� �Y����Z�݌{��cLm��7$���f������$G�.>x����=r���&:E��I��{���up�l���dˮ��k�coX���@���}�f@>� �Y���m�j5����Z��Y�{/b,t��.3@e��4r�P�c��"M�x�-x�Z���zِ�����d ������k��jhm1=y ��̝��� �������im"�m	+t�:�=�2���x޶d��2��J�koǭcK\� >�v`_7^�{��5*UUT�>�s�s��x�"�A�mK�`/[������d ���˭m��-�7iO),Κ�d*�C؂�z��j�b9۞��^���]��r��7�O۳+ ��e`���ﾯ�Xz��`}~�8��L�*[NH�s�� >�v`/[�����]7צ�4���M� �������d��2 _)b��%v�]�N�7��U�{�V�;*�u� >�떚�k546��m���2�u� >���� ���/y:y����>�  �H  �ܓ�w<'u���/�9�S%ں_f��xM�l�\���K��k�<�Av�٪Jm�lDKT��w.Ş8�E% Y�v�%����^��:�V<�Ѻ�s���%���c�����7J�m�۱��H<����c�d�ѷZ�ɱκ.xӆmqc���g��	�<�	=t���q���z����{ǽ�x�?%��Sj����mh1����N��a�ݤ��W��0Z��D�"�m	+t�:�t��۱�����I*�Û�ŀsތ�v�"-G-jo ���>�� wY�{�����Wg;��q�(�$�j\� �}�X��d��2 }�\�U[��py�����y ��̀{�̀wW ��� 򪥸�h��k���zِ���^�`wY��um��ll���]���l�D��U;6�DbyZ�.�C��.�d=���M�6����� �z݀}�f@=� �Q�S��u��u��3rN_��oV$�H�P���w����;�{f䓝�p=*AZϓ��j���?l�X��d �up�l�]�umf��ٻ���u��U�^��Հ����e`���ֽm6ǂz��n�����zL��ɕ�{�2���T��m����sE�"y���ɒ�����S&�Z2un�$�����7Bg�(��~��� wY�{���up�Un�=i-ǚ�l�{ ��̀{�f@���>�n���m����n��`��ٹ$�{�ܧQ�d&{a��VT�DHF��5�-�XV�G���Í.��@"ęd�"Ce��e�i��q��"��BH%ѭ#��ԬbWn�,!	M�t�\ �d�u��H�< � x`m����<���:1@�.����� _ yЂ#Tx*����ܓ�w� \��V��M�6�y >� z�p���zِ��Sũ6$ִ���k�}�f@;�� >� �&4�&�-��Ҳ�B�������0H�-�cg5�9p�7^�qi���>|�G�f�M7�I�X�X�v?������	u��k�Iڴ�j�;N��2�����s���~ݙX�.7m��������up�� ��̀w[2��]�k�5�owq��R���ޘ7}� �wq`EJ�%T��K����f�����]�Q9r+����2�l��up�� ;��.k���մ�gE�qele�뵩��瘂
��^�kګ,�����^��Y �d ����k�}�f@9yѮ!�.I	.�X�{�=UWa�{� ����nɕ�U_}v/�W����wv�wi� ��x�ٕ�]�ݕ����	j�R���j�M��fV�l��up�� ���K[3Zլթ�� �̀wW =mp�����/y�����>��}   h���8י�^�qs)��]M��c{�uK�rn^�w�3ڻjq�3F97d.�s���HgUu��uca�iǶ�����mt��!.B�Ù�T8����ړ�����]u�V�7PzEzsM��F�jW0dt����.MÌ��V/U���s�{�C���&k6)��l�6.nHC��g��r�)@lZ���c�y���0� 뱠����R��t�i���ք�BG=f���Q��'g�z��ko(���[\��2�&V��qbT6'M��;m����u� �d ���֪�f4؞�6�ěp���u� ���n��9{f�Mꌹ����R��� z���l���d��w��i���M� ����� wY��f@;��w7[�V��6��>z���K��uV6Y�4�y�I��n�[���x�&�Ou���=m� ��̀u�/%IU}`sw� �x��x�,�$q���rNw�ٿ*?"� �w��{훒Onǀ$x߈��lCCB��<�w[2 }�\ ���>� �ƈզ�E�mP6�`uUߤ�����2�ِ����Op{���Ѧ� �k�}�f@:�2 }�\����WU\���+$������児�^ܛ �K��n����n���T؛y ��̀w[2 }�\�ِ^�븭�r1G�,���<�*�I� �ݕ�~ݙX߬���$���r, ��ـwwqa�{j�-���KԒW�g٘��� o/lw�������x�U]��x�vV�L����iV�S���o^�n�[2�ِ�����wX�m������$v��H���2W-Q)�NȮ��Fʛ�����׮�Y�:`k:���Kw���� ��x�G�~�2�zSDz���i=�m��� u��>�2��eg��f�X�J�ڷV�Hv��	�� ��ea�}Ws���d�~�r��v�lv6�-�XU~�߫ �����'��rp@�w����^�&ǢoLM���l�����̀}�̀_oW��M�����r�+��ml���S��vڬok���s��Sv6H�i��E��v`�ِ�ِ�̀ʣUO��I��� ��� �l����iV�S��OF��k��u� ��ê��9��s�6斢��!�Hli��L� ��x�G��_�w��7z�9�M�-ݵ@�u�ݏ ��{��9��,��� �$�I-VN����   mm  d��U�M�:�m��V=d�@��U�Ac:�y�����|�k0T�����k���S��;��`i\�\�F5I-ͬ���A�R��"Q�j�+=%հ��v���t�qs����j�Zر���Hպ��wk`W�6��<��g�������d�ݩ*�E���zlv'B�7T=y&&�Y��ݳ�umV+���=��y�uo}R��4�Yu��ƽ���ѹK�u���&���j�b�@�N�^a"��d�' 7�ـ}��Xww�I/����s�=����v��զۢ�x�+:����ݕ�'< �#�}WbW��x���צky���u�d �up���[2�ȺVص�Z3[5��� u��u� �f@�Q���RlI�ikpzِ�ِzِ���=���m��[��#�*7kj�zin�G�}��q�.O�\_ ����� �۹R;���ܑ|7�ŀ}�� {��wY�Wun�����q`n�3VR��RT�V`ws� ��̀}�f@>���Sm0z��<oY >� ^��wY��� �ܓU��kSCպ4ۀ�\��3 ٳ+���I� �K�KlZm�� ��̀u�2 }�\ ���U�Oz6������!m�G.�Þ<�\�e�@��z8㛁�m�����d�̍4Rn�N�:vV ~ݏ ٳ+�~���M���њ٭� ��X�t�� z̀�F��-���\�r`��,��q`*U_A+���CY�s�7$�w���;�OxkS�oS�^�{� wY��f@�c����t�K�/��Ȧ��l+�`��,ԕ*����� o�� ���X/���nIi������䫷�T'^��ݫGG�6	���g\n�P\�Uԕ�I�66��up���>� ^t�}�Wf���֦��ti� ;�\��2��H�us�ffbGw��n�&G�[o��=o��:@�c��ǀz樭�4��E&�[u�}��`;ݘ�wf��UJ�*ԕgu�,��5��m�# ��� _up�ِ�t�^�[m�`vi[����!�j<p�ڰZ�K[r�L��W�uX�5��5��˘�����d��'�ë����s�;Q�;V�M	�i��۳+:�폌 ���{c�6��M*��];o �� >� _up���ޯJ�6��{��������W ��̀_s��r�7^�&�4֛�M�}��>� �� >� aޤT���M������q>~�Xl���4��:��������Hř+����l���{6tC��@H��X�RkN�2!�l! �b�����(�B���N[	�PN�������؇>��'������攎�]?4�bQ��C��@F&�4���b�
*.L� 0*��
`��M: 4�L D���@�����`H:%�2��B�5XG2)�"HJ�:~y��[:��߷��w���                                         �M�^��v^K���8尘ys�s�`�n�\;YŔJ�ks�у�l%�[���W'5��n��N�����X��KY�GP�T���M�sn� n���E��MC$�&��+����{�^Km��d�\�l9�ւr�v���h��a1a�ܔ���	�U@u7]D�Ж�^)u�MFV
�w��Bn��beej���l�ٝ���:��՘x=��v�����g��m�U.�k���B�JS�q���吰
��=��R�r$UVJ�C�ڨ��YT�R���5R�T㧦��B���hK�kD�� �U���ԝ�k�ڪ��v�U�2&� �WJ�8�'��­���UHZ%�!����Ҷ�n��ה\!VԄl�v�mm���jW��;m�Qfm����U�`G^�l�sZ�[������@9Bz�*��kj!�:$�a��e�*ph��u�9ͥ���l3x�-X79܋��s��I�L	�n����)ר뗃�	6շ<�Яv�\����v�s�7Q��eM��I�G#��8�b܇�Z���+h< ��I �I:^�@i��&ʝd+1!�d��$��`U�A���j��P�W���U[e7c-���%��Kq�'1�6�4)�i���
Z\Q�ڥLֈɳ�]���þ:��8o]��ղ�6+v2�vޣyF������n�-tl�lcs�q��TݗN9t�v��O��kln�p��{:5��k<v���;uj�����Pt�;��9#�n��v(u����%A�N{,�uuۓ��]�V
��g�
P��x���i4�q�M����|�n/v�R[:r]��T�/I��+�୓��aݲ�e(J���g]�c�.���!<lv�t�l��\l��5u�k-�I��a%X��S�S@�ኇ�O��iQ���$^��|�)��~�sy��fff`  ����  �Ѧ�%�j/6n�GJvˬc�V�E�wD����f�v�u��82a)NT�⮸�2�l���!"T'vڝ�]N{]9z�D����al�ݕ啻������0��j;\O�;v.ڿ��c�[*�f3�)36�lu��R� F�"4�������/%�s�����fq%�i�N�qf�svb.8�q6�Z-�$�U%UJI�I�Y��21�[D>����U1v�7X�<��u�s��:DZ�j�}���d�ِ�����{n��i���M�i�=&V ~ݏ &�x��������<�9qH�8�H���p�f@>� [f@ʣUC�5��5���;�̀}�f@>���۱�� �^|�M4�`����ِ����f@*����u<�l�l�;jݷiWAc��v�:�� �p�V���[��sؑgt�Tc����� ���;�̀}�f@>�zV�G��W �X�{�;J�U+�Z�B�V0B"�b4D������s�۞ŀ{��Xۻ�<�+����f���֦��n4ۀ[L�}�f@>�̀wW ��U�M5�E�����:�'~���+ ?nǁ�w�s�6�.Vؚhi�t�u�OI��� ^��u� �km��boQY�2�<�ݓ��]]r��[��h�k��/ �S5�4lڸ�3��d���ϯd&���?l�]U������ �r��I,lr�ɀo{���T�]��{����nǝU_]�+�V�>M	��q`�{��Ň�xI!I$ �U$�*�If���=��,��-뷯L{������� ���^�2�[2��ҽM��I����[����fgr� u� [f@<��v4YةZ�v�ece��w���l��s����3sZE�^!"=&��ِ�ِ[f@wW ��U�M5�D�o��>�f@=m� =�\ ��=y:�q涄�ѷ����ِ����\�do�DD�V�1;u�ݏ 7d��9��f��� !�ALM��9�� ;ʣn����7Mikp�� ��̀z�2 }�\�����`q:�.M�ۭ��{t���\�l��.q�v���&�sMuy�u�˝���ϳ �̀wW �d��mպ�i��K�`��Y�UUv����� ��2�yEq�m5CTҫlM� ~ݏ 7dxw���]�N��7�������{����Z-ƛp�� ��̀z�2 }�\�UV�i4ּ�޷���wY�[f@���ָ ��R��T�
����I$�I$�@�@  a��y���z��Mm���d�^�4�&&y�XuH�=���0<̗e�k�8S����<������ݡ��s���ݖ�F�����tFv��8���sY����p=�:�l�m3i�&����L�[���f����+��:����ю�q`�]��"�vH�9m�5�rݧ�a���;��Y��rT}IU*�U:B����$�I!n1^R]�ݮ�u�69��m;z=��]+a��^��Km��r[$�䋠o�ۋ >�W ��2�u� �ȺVޭxތֆ�@����"��d��� ��2y*�I]���g�. ��1˷&���@>� [f@���we��S�^��^�{� wY��� �����*��w}��6���;r;�i��K� [f@���wu� ��̀}���ƌ�^�Jݍ�ig6v�y�4\��ڄ�z��y�ǔ�.D���SS7F��I��wW ��2�u� ��2��W����vH2ڗ$�;��,uT�\If��vd�ِ���z��f4�4e˚��f��bX�v�eMı,K���m9��CQ5����7ı,K�{�m9ı,M{Z��e�j�kS3��bn%�bX����iȖ%�b^�^ʛ�bX�%�{��r%�bX?{�17ı,N�z��5na���YffND�,K���T�Kİ�
G^��ٴ�%�bX=��f&�X�%����ND�,K���i�u#�n-lsϫ�H:9�Ը�ӗ]��+����l�ոV�F��'hͣ6���%�b^��ͧ"X�%����q,K�����"X�%�{�{-,)z��e+)n�xv��q�v���,K����17ı,O��p�r%�bX��ײ��X�%�{�{6��VR������� �q8"H�n%�bX�{���Kı/{�eMı��DB 	"@�PJ$b*j�iWq7���m9ı,{�17ı,O���}���z^������{��7����T�Kı/{�fӑ,K���ى��%��	������ӑ,K��m��q�rƤmK�],)YJ�V%�}��r%�bX?w�17ı,O��p�r%�bX��ײ��X�%�����ϵ]Ur/6N�e�c�i	�&�ڛ3nL���oW F볷Vr�t[Ok&k4K�ͧ"X�%����q,K�����"X�%�{�{(~ ����%�}����r%�bX>�����e��q�qBH�,)YJ�VR��������&�X���쩸�%�b_~��6��bX����Mı,K�}g���R��e5�k0�r%�bX��ײ��X�%��w�6��bX����Mı,K��m9ı,K�}f������X�nK��+)Y�$$�[��ӑ,K����17ı,N����K��� T#
i � ND��k�Sq,K���ޚ��u�˫��jf��r%�bX?{�17ı,N����Kı/{�eMı,K���m9ı,ON�y������u�PnWv�gC�\p6Z�SF��\:��T����=^}.���$$��6��^���7����߸m9ı,K���Sq,K���ND�,K�{f&�X�R��y5;��Gp#R�n9R��e%�{�{*n%�bX����iȖ%�`��l��Kı;�{�ӑ,K)YK�o^7q�XӉ��$�K
VQbX���iȖ%�`��l��Kı>���iȖ%�b^�^ʛ�bYJ�_som����B8��YK╔X����Mı,K���m9ı,K���Sq,K����߿~̥�J�VR�V�͵�.�'q�qBH�7ı,O{���Kı/{�eMı,K���m9ı,�혛�bX�%B ��g�������� 6��  p�T�����նҝ�.�1���#ʛN�n�ȝNl�u�V�4��.ѮNL�Z������?��|�g|�l;m��$��8*��bd�����*��,U�ʶۮjOj�n�n�]+�8���5L��UV��*��r�;���6�&�޲����]vdml	 �5��f�X!`C���g���V�n��{�����/�����C7P�����dXyRy�՞s���t��.�oi��v8��hJt�s������{��7�����Sq,K��}�m9ı,����MD�,N����ӑ,KĿ��c��Y D�rK��+)YJ�]�ͧ"X�%����q,K�����"X�%�{�{*n%�bX������r����s)|R����U��R�ı,K�{�6��bX�%�u쩸�%�bw��6��bX�'��K�շ�vE%E)aJ�VR��7w唹ı,K���Sq,K���m9ı,�혛�bX�'~���Y��Ke��YK╔��e+�^˥�,K����m9ı,�혛�bX�'��p�r%�bX�	��2���%
�1�ׁ���X�8�k��l7f%5h5�n�()=�<���UD�I���7�Nw�`�! ���&�z%�b^�^ʛ�bX�'>��o�.h��+�2��+)YJ�\�ŉ�|"�D6�Q�Mı;���Kı/{�eMı,K������/*N�2���~m����8ᩙ�&�X�%��߿p�r%�bX��ײ��X�%����6��bX���R���e+)u�ͷ�;��',��iȖ%�b^�^ʛ�bX�'{�p�r%�bX?{�17İ?)K������+)YJ�W�Y�����fK��7ı,N����Kİ~��bn%�bX�{���Kĥ+�^˥�+)YJ�]�ݒI$�vӗ�*7k���=��ez�vx��g��"O����u�;nW%䬔�Cw������n{���Mı,K�{�6��bX�%�u쩸�%�bw���"X�%����		;�6��]{�oq�������ND�,K���T�Kı/{�fӑ,K���ى��%�b}ɩ��r;����e/�VR����{�eMı,K���m9Ɓ��BZ,�D�����۱7�8�O$C�UwC�ye���.�*l�6K⚺���L�k@�]F�����<�u<�4�$MMh3 E`U�����A�5MR0���I�g�5YYR6 FT�a`Wb�3��9Ą@@�(�Z"���,�jF�kQ��
`b(� r4骸���bk��|�tCT(��߷g�)  �
 Q(!��y���J� � z�D�] �4��D�L���f&�X�%����6��bX�'ӷ�޵��p�5�K�ffT�Kı/{�fӑ,K���ى��%�b}�{�ӑ,K�j&��~ʛ�bX�'�����K�$$�]�2��+)YJ�_{�17ı,O��p�r%�bX����Sq,Kľ���ND�,Kﯦݰd:�\�9n�)S��Ws�K�b�w�
��.��75��P���s+�v%�8jfa���%�b{���"X�%�~7ı,K�{ٰ���蚔��b��JXR�������5�I#rk5��ffND�,K��{*n%�bX����iȖ%�`��l��Kı=�{�ӑ,Kľ��{53SY��̳2\̩��%�b{���"X�%����q,K����ND�,K���T�Kı;����㫙5s5��fa��Kİ~��bn%�bX���iȖ%�b^�^ʛ�bX���4�B���� i�@��( �q?{��m9ı,O>��r��(Ɯ�nE)aJ�VR��=�p�r%�bX��ײ��X�%����ND�,K�{f&�X�%��>�����p��k��\pDΝ�,��<�vѪ��j���
<��������a��Kı/{�eMı,K�{�6��bX������D�Ke-���)|R������o�����0ɭ32��X�%����6���U:���~ى��%�bw���iȖ%�b^�^ʛ�bX�'�v��\R�F�	#NܙK╔��b�n┷ı,O��p�r%�bX��ײ��X�%�{���ND�,K�^ִ]��m��$�R���!&R��6��bX�%���*n%�bX��{ٴ�Kİ~��bn%�bX���u�r]��pW�R��e+)YJ�ײ��X�%�y�{6��bX����Mı,K���6��bX�&*:�ϟk�   [@[@  Sm�j��8�����0�i�M�Đ�L��\�j
)�Z%G�NK�]�p������e��v�풞�l�Uz�utt�;v]�Z�r�mę�A&���3�;�6W��@c<NJ4\�@ut��m[J�h��*��p�NqΜ��msd��cB�5�p��˳������j�ݹ�\dkL��p-e�c��ww���-�	n�ؒ�jMY�T��������q0i�<�u*����3��'3Z�s2��,KĽ��ٴ�Kİ~��bn%�bX��}�iȖ%�b^��XR������[�w�K�����fm9ı,�혛�bX�'{�p�r%�bX��ײ��X�%�y�ٔ�)~T�)YK��-ܷq�2ڒ���q,K�����ӑ,KĽ7ı,K�{ٴ�Kİ~��)aJ�VR��9:�c������0�r%�bX��ײ��X�%�y�{6��bX����Mı,K������+)YJ�\;{�����(6�feMı,K��m9ı,�혛�bX�'��m9ı,K޽�K
VR�����ݒH����n(�WY�%�ctKfs�`[v�S5m�K�ˇ'k���i�"�ӵj��{�7���{�����Mı,K���6��bX�%�u쩸�%�b^w�ͧ"X�%���Q������|��{��7����6���� E�Atn&�X�٭�Mı,K���6��bX�*��)K
VR������۽��-���6��bX�%�u쩸�%�b^w�ͧ"X�%����q,K�����"X�%�}o��nk3WY��ɭK��7ı,K��ٴ�Kİ~��bn%�bX�w���KıW޽�K
VR�������1�(���p�338�D�,K��l��Kı>�}�iȖ%�b^�^ʛ�bX�*��ٔ�)YJ�VR�J�g��i�$rO<���6�ݺG�V:��hӫb ��G\ݮg�+a��G.�H=^�������,N���ND�,K���T�Kı/~��iȖ%�`��l��K�VR�N���Gp#�4D�)|R��ı/{�eMı,K��{6��bX����Mı,K�w�6���UJ�]%�F�j�Ƞ�$��aJ�,K��{6��bX����Mı��p4��@��]"R�=����"X�%���쩸�%�J\�om���K#�4ۓ)|R���������bX�'��m9ı,K���Sq,Kļ｛ND�,K�ߩ���#\�Ϋ�w��7���'��m9ı,K���Sq,Kļ�}�ND�,K�{f&�X�%�u����UZV�+v����n����f��wN������{#��u�B39�(]Y�ӑ,KĽ7ı,K��ٴ�Kİ~��bn%�bX��}�iȖ%�b_[�[���ֵ��]K��7ı,K��ٴ�Kİ~��bn%�bX��}�iȖ%�b^�^ʛ�bX�'�=�M^9up���F]fm9ı,�혛�bX�';�p�r%�bX��ײ��X�%�s�2��+)YJ�Z���[�dN��5�17ı,N}�p�r%�bX��ײ��X�%�y�}�ND�,Q�"��F	 *��"�pt��}��Mı,Kﳺ��\��Gdh��R��e+)YJ�ײ��Kı/>�iȖ%�`��l��Kı9�}�iȖ%�b =�?�����Z�K��l�u�i:d":J1���.p�c���y洍-<\5�^���9ı,K�}�6��bX����Mı,K�w�6��bX�%�^˥�+)YJ�\�om���wrF����r%�bX?{�17ı,N{���Kı/{�eMı,K���6���A]T�Kڿ�t~�\���5��S3Mı,K����iȖ%�b^�^ʛ�bX�%�{��r%�bX?{�17ı,O��;uu�f���d�.��"X�%�{�{*n%�bX���iȖ%�`�����Kı9�{�ӑ,Kľ�{^��fj�Z��.��ʛ�bX�%�{��r%�bX?{=17ı,N{���Kı/{�eMı,K��O!چ�����}�   -�:@  s��,��BɌ��m�Qa��b�z!�M&4���'�D��ɨ=�]�b�h��`�8�1-T�)�m���;;3]����؉u�\�@r�E��)��iƬ9M�7tA�s�eIf�/��Yxz#�ۍݙ�	�+��ف�ݛ�ܽqO=z]r���N7;-W]��1j�$"���<qKpW%�)~UU�J���w���|������z���l�X��r[\���jA�� 
Ew�Q[��f,lw�,q8�.I�^)YJ�V*��~%,)YJı9�{�ӑ,KĽ7ı,K��ٴ�Kı=�����j��Y)�5�17ı,N{���Kı/{�eMı,K���m9ı,�����bX�'����j�j�f��fa��Kı/{�eMı,K���m9ı,�����bX�'=�p�r%�bX�N�o5�f���d�kT���7ı,K߻��r%�bX?{=17ı,N{���Kı/{�eMı,K�}u�d�&ja����fm9ı,�����bX�'=�p�r%�bX��ײ��X�%�{�}�ND�,K�U��{�fffe�['!.�m���k��k����cɜ]���@ �x.���z�4��k���ı,O�{��"X�%�{�{*n%�bX��wٴ�Kİ~�zbn*�VR��_l�z�#�չR��ı,K���Sp�Y�hԐaO�PP�~k���b^~��m9ı,g���Kı9���ӑ,C{��>���ղ�a�G����bX��wٴ�Kİ~�zbn%�bX��}�iȖ%�b^�^ʛ�bX�'�=�M^m�I��h�36��bX���LMı,K���m9ı,K���Sq,KĽ�}�ND�,�e-}5��b��Zdr���bX����iȖ%�b^�^ʛ�bX�%�{��r%�bX?{=17ı�<�>}� :��
�)+v0��-�:y����-�y�ɛu[������Jf^�ՙ�f�0�r%�bX��ײ��X�%�{��6��bX���LMı,K���m9ı,O�o��ֳD��3.�is3*n%�bX���iȖ%�`�����Kı9�{�ӑ,KĽ7ı,O���ֹ�䙩�r6��e/�VR�����IK
VR�,N{���Kz@@?"C"dK��쩸�%�b_w߳iȖ%�`���~���.��6��7���{����ND�,K���T�Kı/~�iȖ%�`�����Kı:���D�Vd�/w�w���oq��{�eMı,K���6��bX���LMı,K��m9ı,O����w����伴�J�[����X�*[���֎�j�l�����qjR�F�d�d��f���3*r%�bX�����r%�bX?{=17ı,N{���Kı/{�eMı,K�d��kd�Y&�ᩚ��r%�bX?{=17ı,N{���Kı/{�eMı,K���6��bX�'���L��C2۬���fLMı,K��m9ı,K���Sq,KĽ��ͧ"X�)X��4���e+)YK{:��q��3Vf����iȖ%�b^�^ʛ�bX�%���m9ı,�����bX�ދiV@E#�D�T�! �=�|��r%�bX��~�ۍ[��W$�K
VR���{�}�ND�,K�{x��bX�'=�p�r%�bX��ײ��X�%���w��߿�ڮ���Н6�;g��[D�6���6y��cmq���ځ�¢-b�t���ܓ�\)YJ�V*ｒ���bX��}�iȖ%�b^�^ʛ�bX�%���m9ı,��˚��S0ˆL���Kı9���Ӑ��MD�/���Sq,Kľ�fӑ,K����&�X�%��v��]_]a��2kE�a��Kı/�ײ��X�%�{�}�ND�,K��x��bX�'=�p�r%�bX������2\�Z�&j�̩��%����w߳iȖ%�`�߷���%�bs���"X�%�~7ı,O}��ɬ5��d�ˆ��ͧ"X�%��}�Mı,Ky�{�ĐI��D�$�O����$D�U_���
��U_���PU�*���������
��T�_��H�@�DP*T��E `	@�DPT��E `�@�P(�T��@E bDP 0T����P AP
EX�(
�PU��*���誂��*��AU^����"�
����*��*���誂��"�
�ꊨ*���*��b��L��kFov� � ���fO� ��� } Ԁ�  u�(  �  *�U��C@(k@   :��RU!*"�AJ��R�	 �	P*��IUU$�UJ��T�TP )!T�`   `      &��S��νg�oO'�����}� p�����9΅wt)W3B�� �n���@   �gTvPn( ê�@n��P�4��
� 3��΀S�S�!� 4 
   U  '@  0        �          �1�rQ�tX�h[��.`�n�p�
uK>����r� Zs2��Z 5K=�٫��V�܅�W������웞�}c��q;�����Ox��  H  
 3`�����Yr��m�o��g��� �{)�77t�����g���@����x�� 0���{��g¾x ﶗ�k�l�m�ty����xyTbԋuǾ�K͊综����      *Llϯ��X�S�v�������9�p�w{5��}��|�导��n,�� (���r�{v׌�� �^OJ�;���� ���9-�w���o%睎���
�׃�˶��}y�}��q��| �@
 P  l Qϑ���W�u�ǋ��ɪ_pG��l�ݩ\�wݧ�^�����P ���i��� ��g�6�z� �{��f�o�e�t����w�*�y+�n��{y�d��<����W� i�
m�IJ� ��M#ʥ*   "x�T�f�OI�FA���U)&$�h �)����R�  �
BM�)� �S�O������?���o�'�	5	K���GX�{=��� �*�079� �*�QEO�(
�� �*����" �����jI�㦘��Fk�D�q�F��a�lt�f�9�Ml��CIi��lݯ�޷����<-�,��lPBp�a��=��D���p'�.Z���~��wF�1�盓�"�02	1�tbHi$"�"37�j���G�.?l,�� �%���[9�s���h��&���$%5�C\&z �X�3^���~���TP�L�>`��@C:�n-p5�!�0}�� 3[8Y���o��oDf�O�?���-�M͋q/�Nu���_XF2CN20��٧�x~��2�~�� ��V�;)�G���f���)�f��e�s�w�yg��<,�Ґ�8����3K9��E��,Ѹ�F��b�����akNi-6ŧ���y��,.����p�#($��b ��Ԍ �~�����,��hJA*o.�`�گ|���0\�M%w
1���qch�0��l)P�U�dM�J/ʾ��;�b����l����a?e羪��n1���Z�li3(4p�~�e�ٟ�n2)�C �IĀ��`1"���!�*"	�"q�̮s������dm�
g	H���#2+�񃆢��J�ٳ?s�<-odE�4�l4j#ٯ9k\�ɢ����-	�Ijip��4da��,3Ph5�y�o����I8��`i!�H�eXh�Y9�F�������y�ՄˌL�����%���ߜ6^��yh�@��g�ƒ7���o��PT[3+R�N�f	�HcN������=7l����7�^�әj���1��1�Ń4f�&����4o~g�瑫���O���1��l�-�4󗊧�~{�ǹ��m��$���b��F��Y�y�s��N�c`N��x߶��O�~������	��&# cԱY��f��_��vîl�m��DIA� ���DL�Y;����XXVLV{�����f��f��"�o�`AoE̲�Y�ms�����2��A%���Km����}���Y:3aÇ��a�&$���� �	��#	�OH�Ijq�=��bD<W�����iÏv���A����D�'(	��3"J!���Q���k�p�f�Y��-���m� ���Ǚ�< ���L���%�/����D�y&@�Ok�/���~�ǲv�S���
/�yc21�v��	Z��@{�dz����1�)ɽO�md!��m�4o�����s��?��{�g�秅�<߷��^��M�0h3�10`ˌd-I�k{��{�Fzm�[�w�+��~�*e���9�ߧ��~���9�"��@��0)RJ��(r0�����zcQ�㪵Qz�o�3����71�p#ǐ�Q}_�f�֩���v�d�&�a���yfe�	�Ut��ĉ��`M���\6Nj�3��(�f!��0�xt4��}�mN�&	����#(4f�I�9Ç�#o<7�za�L:p�aX�cf�x��OX�`�8L�f���X~
`�E:,�V�~w���O��D����i��3F3�~H�F����!��a�؇x>X��� �5��s[�<|x~6g��ˆ�͙������$�В0`A��#$É7���ɬ�рó�OϾ�f�hII'R|8�7��e�hc4c�dc�06��z�f��@A�=X!�:޿a��^xc���z��p��06��َf(w�7��{x٭�]SJHdHF���I^&�Lb���Y�/߄�v`��L�n�f͓��ɍ�bl�,�'��)!*���)M��ٿ�*O+DJT�@�+ޅ��9��HH��'�t�55�z�]�f$������MS�k�Rd�!�1�'!��o�jv`�0����\�m㕯9��q6q6�lcɄ���Bc�r�0��g3�?kI�sykl1�O�|6���Jmg��/����k���vC��3S[���V���=f��Y����9�͘,�'���r=�fDA�di��y����9�X�����j�G��N`X��+[��1Ix��y�2ty�i5p՚�`U�5yA�z<�[4$NFd��f��E5G%���#fZշ|6��#~yo��:��[��(��G�0�ߘ�f�p��k�֭��fk��tA>p�|$1�ᣇ,�g7�� ��=���٥ �I�a�7�<��i�82��8��M�y��gǞ�8U�6q������<%A��gx�8ꍇ���~K5�y���85��p���BC���S��ѯs����3[`�[��23���-0I2k�j�����o��/����9h���#�PH@a8x�.��2�Q�{�����,ӷ���G�%oN���w�.ٌf!�����/�����&�}���5y���S_�3Fk<���I�N�.�A5O�	!w~�w���ٛ�a��Ԃ�)��v����I�P-�D��&� Y9~ý�sF�߼���#ݧ��֬���"%
Sk))=~^̂j�K+0�&�wq���)8N"�X�	�(�ua�䵣�a��O&!���7���1�I��wsΛ�Nc�a��kg8~�%����Čt4�[�xI���Ág�hߜ��qto_����3I��4m�f�g���V�tA�/kz1�ٮ��e��FU���e^(���zX�4��� � $���ޞzxp�2�lxDO�Fk|���l�7h�6���Y�q��a�ɞ�g��ı��3F�����ĜP�b	sF�5�6l-g������o�1�`A,&:a�(6d`ch�lSg�6�h��#�G�4�*�T]As��iϲ�
R?'�Y�w�N�O��}]�yq��I��=������p(���3�/g%!�I&5`�0Ն��q���H�=�%;�̓�=�G���>���y�oa�l�o8lLIL��D�l%	*5{�|p��8Ꝅ�q��K�Fkgo��4�o��Y9xTb�HH�$B��&�4�9��
���Mf���E�6�4Z�f�٧\<�k���b$�ń�%���02pƦ&�V�md��?*s[=��?g�h6��O�Ə8���ќ�[�3����̌����	�p͛�Ƴq9��<4C0f�D3	,e�a�I���=���������߿p�}�7}�7v.6f�yk~�6Fh�9������oÚ�g��A$�+	K$�,�A!"@K3����0��/�����5��N��<�zډ^V�Ͻ����_��i\
U$)I��A�!��:\�FI���d�DD�D��IA$�A�d�0I&ή�Z�Gq�a��+/^�䙽�kә�d��`D��!ČZ0*0-y۞���P�Er;��p�	(0���lc'��	#IG5:�2��8y�D��Ț�*q'@F!��ٮ\�3��3�0��"�b����	�_B.���f'��E;9�	`�{D��x�y���_k�1\3eyg8~<=N%2��?�!(I\0,��,5�x����l�T���Z����Ե;X� Ba��5k]��$���\�xc��Ǿ��}���D��
8H`�ʛN%��x`�1���1��İ#KN�4Fk���f�F��5w����ݎ����������q��d�cRa�|�?7���7�f�
HE_ؑ*���s���Ц��}q��0K&�$��=�����=�鞻0�G��5��mD3FA�2K$F�	�U�_���#|�Z�&�s^o]l��bf0A��#�H&H�(4p��*�vkq�f���3�p%�r�0�Ç3Čp�Nhc-��p$�Č4�i�Dp���z��Ӹ04�Șr� 1Â�H�bA$2�PxC�� ����7B�8)�����$��\�WC)!:gpߟ�2�ȓ�N�6H å!"HHI�  �Ğ8B�H`���4~�ͱ�0WIb$��R$0�CŃW����� �      ��  p     � m�               ��                                       �  8��     �           �l  -�  mg�v��u��ўvk��鶻Z�8�i��m�K&������[s�h��[E�^����l6݀  �M/SE �`�ö�m���m-�t�nĀl  m���Vk�		 �m�  �ӥ��Ѷ̝"�s���l�8.���[$��` ��H,��@Cv��m� 6�Ӭ�ƌ�f؇h����X���mm�|a$�F��v���-�5�o��g&�B�ړف�^�U��nZ�W���6�;|a�U�d�9�
�����m\�9"�Y]����M� 84P�nٴ�DV�)onY�Ue��d�k�v�*it6��� c\qr�[���}�}Q�F�ɥٶ�k�U�W�)��A�h3�-�fٵ�    2ib;&`kd�ˌ���[k鲡p:�j�ZVۀHl-���m۰m��6ݐd�$-����,[��*[U�l �lV�J��l��J8��^��of䷨�mUPVy�s�*�T����h��6�6��ڪ�; 6U���6�t2��m}���t�{Z���<n�Dd��@!��n�m�6ʹ�� �`  ��p�  �}�ό�m�ͭ�i�[-�n  ��d[L�� q�kn   �� �`��m%:k�n�lR�ʵ�����PU*�b�Uy�꣍�j�yW�cP���.�l�q@.�\$K(I�m��$� ���;M5�pm[qWUR��&g��$kix+V��m�Y-�  �U\�/-��-�T��D�T8梏6U�Y�!����Z��
�R@��I��lk7] 7l�$��:�H�Hݷuu���N�I��zI�]4�@r�Vqm�ijLt�l�   ඖ��[�'�z�m��oPwf��ܼ��֕`:�j�8[C˥�gj�6�v�*Ъ�L��wcr�mUT��   l�v�mE�6�6�9'"�*6[�� �&���i�N��&�3 :E.��BFM�b� ��j���K]6U��5�r��@8 [d i6  ��Z�Ua��L�ey�k.m�(+��L�U��� H9J��g7j�:�ke���c瓾!��mH�-����me���T�@�ܸBg��d����Xp:A�J�04��eݵ�[)�+�m�P]P��^{(�Mhp[�$��-�l��6� qd��H � ���mm [@moVY�p [Ym��� ���� Vղ�8�5J���RǤ  շ6�N��Izm%�\�U� lip�Um]�!*d�ei� �` �ޖY 6�  m5]��w[�r�! pn��0[B@ l �-� H  ����m�,�  �xr��@�[�[u�6���nհH �[p���5ﹾ����vI%�@ ��  u�V�:�( �[���� h#�1 v���aml��7�g�.cj-�l�T]sb�     m �-�   $"ޫm��o`�`-�   �l[Zmx-��Ժm�i; E�ښ鎓�-0R��޲6���R�R�$5@U�[GԷ�R�S�;\��H�5�J�l5@[T�m��86� �  ��h p  h[dm�[I�   p   	      �u�  	      ll�� 5�[���Z4�WT�R��KĀԥUV�T�V�Kʹ� f�`�hh ���  H  l  [@m�r@ 8l�$i�ŴA����0      �#]�`ZץCe��v�$� �J6� �  o�����h���     n�d�ya��ۀm���zv�ٱ�Q�O\e��nTTC�b�`���:T
�t�7Q�%,V�
����l�km�m�'G&� m��h���m���r�]��&��6�[H]6 9f��I�´p8�[[UP%Im��J�3M�D$��� �Ŵ h�/[\��"@pi���iR�t�$�n���+�夑+�6[@��� �����BK�@����6,<������5WUA ��6��x�D�'@mU[l�m��x
�h
_9l ~��v�|�M��Q  �4�v�� k�$�m�m���[R[���9,�ڶ�6��:J���W$�9z�� ۶�i���nضK:-��)W�U�'�a�\��v�X֚:��������~�����H�UPvt�m�� H�`�2��ͻbD�M�m��6���7n���Xq��@����3�զ�[\6���6�@m�Bڷ[�m�Iz�l��l����۶E �Iw4Y4u-���S��a�Yj�� ���]{I�[�:�.i�u%H ��Ua�� z�-��	 ��h      ��[@ �ᶳ2@ [@=	Z�nm��ym��L� � 8m��\ ���e� A��2�]lTpR��= 9S���vi�:YE8�!�	�m�E�p��kj��n�e[B��� ��J�R��]S��[C��m��n�  BM�m�N� �z��&��Kd��P`ְ  m�bʡ5[�Q���lb�nCa�Uu8q �R�IWk��gf�B�ݪ�h%��I��8[Gަ�  ��kn[Mo0�i!mm�k�����h�S:��٥��lN�t�v�fZ �9$u�-ܷP ��=� I:m�7O������U@\��η
�U������-b���չ�L`܋h$ٲ���« QTT*�;A9�5�Tk�	@�ց�Ƒg'iV��޼�����Zꪱ��ml��u\[BNuҴ���(�V^����@*��5@�`m������l�/1TT�iV��"KؽRu��Z݀$m;��ڠ�'FR��&��M�t�p�Ӷ� H(6��֮���Wgj����4}A�;K,� ��f��]��j�l��mͭ�Km l�  ���K#m�o*v�@EjD�}nҭ@'D������۶�#�[|	�M��	   &�ۛn֛a *�3�� ]3m.�h
UU�nZ�S���m��[@ �cj'������b���uToU�[H�`6���u@]U*�t*[-U�m&�� �E؛�Z���e���,]U*� ���������*��@*�iZ]��%�H���t��Ut�^`+�ĵ�]�h�;l��յ��8��,��v����>Vv�em�kӷX�Lp��&I�*�J�n�P��d:k�5.5�t�V���:V��u(�j�vm��m�+,jj�8e@���l�d�H�[��0m��{c��mpΝYwm�m�6�ո �5�ۮ�X%Z���.��6��  �:�N6Y+z��)e]�5mT��V܏.�.�}��V���v=�ҭUc�pJ�1�YXrʛ�ݥ�ڕ�v����Q��l�+9P���P�lވɻm4����I�v��Dt�\�wSek��K�]�I'GU�� �t��������6K9e�����;k���	�'~}�n���Pz�Z%h�6�%�%g�2[)(��Y*�?���l�iL�l�'�u��䏋7|���:ꯁ�ږϑ���>V��C����N��Wb�OF-�:��y%�kd`�4�e�m&1b��ӈuΠ�T��ԭf�wZ�Ė���ڶ��Amk+'�[@Zl۵�mӉ���a�v��U��B��딬'4����e�m� -�Yr-��cq�	%�mp]�lI¶m�F�z�33'[@}�π[\[Y6� ������n�pm���w�l��^����X��8�u�lH8   m�s�۶�հ�  o������6�olݲ�   8  [x^����n�  �l���l�q� $nY��l �������U@m�M�$��[=�+P �ݰ�   %K6vm��u�yn�m�P-<n�n�c�g��Vl 5Ul�R�������m�hHEڶ[M��e���[�8!��^�N$��ڶ�K�Z��ـ�]hIKƵ���7����5��y�V�b:n�����C�Ҥ�(b�Y�/N][V۫v���az� m�/ 6��b\  6��$uUv� �shiv�{B�ʦ���T\�]�e;b��bD�[�À �`ݠ*��؞nlS��E,��-.ѓ$�Q��@�MV�[ٙ�foZ�͙e����T@qT6���A0�d���aO�/�t����B��A� �
qD?�"?������~dx/�'����\A� @�:��@��:D���x�!/Qʁ�v>��� �L/�������P6����je6�wOOȡ�C���F�(���Q�z��*����� C��l�({p� $��_�#��6�/���@���z��J� �QS�Qz�ߡ�E !�HQ���A���z��=(�a���*����8"�1� �Gb$:Wh1CgB||W�m�����ء� A�����!��!1���0��P��v�G��?*>*"�N�SG����hT<4��@���
�� ��D"��x��m#�B�$�'�K��AG��u��.��N���%9�0�]����`uN�% %X 	�CB@^� �>���1�v��-��!�J*o���(
���B}$Ĕ �A4��J�Bʚ%K0�d$�{��~�m�� �� �  6�       	 �%�����.�p]
�K��B��N�)*��r��
���^�W�<���	5��2)�=2�<�Tz.�z��hPZ�G�^l�d��aQ֓�@�t�����/[�r�7[�\��]�k��D�vq��X���r�D�d
���UK�k�s�uP���A��Q��K��ڂL\��m؁�z��rX��j�Q�h͵�-F3��ܙ�wY�l<ܚ�tV��V�.�@��
ٵ���S���t���ls,��+A��m��i�-Jt��=6�ڝ5غ]��J��6�J�,�Ƥ.�MJ��8��p0(
���*�����0M��j� Um$Y�\fg�rfQ��8� t�"62� ����u��9h�U��X��W�"+�壃��M��a�m��*��5�
�/�)yk(��UWe��볮�ss�2�cj����7�i�кZWg�.���Mu���X�!L�'�]�5���3ӥhʖ�9��in�l�2)+8�h���9�4/<�&��� ��v�rOl��jh�=H�+uF�Bxu��:���t�Fz�Q�n���ӘYmnq��U�l=v.�����cmy�y��-�.�yS64����%��st���8`x�}�^G��zR�kr�]�r�W`$ʞI�ìbtURu*�+���d:we�t۲�j֬KU8�iKg#n���v��np�S�Fm����`��9y��O�6��v7��^nnܙ�Jzq����
@"�r��B�����u����H�!&��`�{��n6��ƶ7	���rvvC��;m؃��=(�M��n9��hq6���l��1��(���6�΃iV�N�;���䪹m@������a��c��*�y5��q88�F���]�n���װ�l\�]J�-�e�K��u�ٝ>k��q����[Ֆl�Y��
��>Q?��G����:��Ci�����=�~ ���w��{����~��l�
�UQ[����������Vx6և��8���^s�z�Ӥ8GWm�]�E䫡���7[ǆ� ����Y�N�l�:�n\n :�s)��<��JY���ιq�J�]��6n��i��/g���Z��K�<�)�q�pj�]{8��`4�#��"۝��u;�}]���wQTf{sZ_
��lu��m�Mz�p`�V~���s�{�}w�)�78Å�����
x�v�c��.���#��/=��¸;q����ܕhd�#�%�y�[�2\l�7���qh�S@;�f�{n���Z�`���6M��S1� ���Yn�@��V�et�"�O�rB@��+�h�S@;�f���KH�/�L1��M� ��0u���� ��(����_�{�]L���̓*r�ٔ[I&��n_h��vjeA'n��G�a�	�m�6���~��ƀw������ڴ
��[�8�Ǔ��� �m���}�O�B��b#�$��b�>��8��?#;��ł�����/m��=rՠY�� �נO��س� crL�9]�@�}�@;�f��v�|��|�U�UX�H)���ֹ��� ~o�M�Т���T�\'M<Q�ŷ���gf!N3��u�2n����[�N�Ϟ����넿�1�]�؊?X�߯ ~o�M� ��������ҹ! rM����ڴ��8����IDL����=2u\ą�U^�U�����]�^�9(z�*��2ʘ��	�"`�I!��������ԓ��L�#���yz\�	-z}n�@��V�Q�+v'x�|7#��٠s��h�ՠqrנqr�PMD��$!�2��\67#�m���=;��G�]�Ǯ�gv4f�#&8���!}ܚ9n���Z-z��4ø]�	�""��k ��:�2l�u`_u`��X��%x9#y	�1'��s��Z�a�(S>�ذ�� �yK��*��G�*���?w�s@�v���H$���N�s���U���+���������9]�@�������G��##��c�������IVȸ�M�'�˨9����D�flp�[W�KH�,œ�L�9]�@���������v�s@�tu%��O��28�ZW��)nh����-ZG.u�J<2|6���٠~�n枈Jgz�� ����>�j�4�L�\I1tU]�tDD�_|�������6u��^���M�ۓ4Wj�9D/V���r�� ���`�!����� 	���%��E�d�ժ5�qq�s�Z/�����A�'!�:�ؙ�a��_}ط-lvs�66os��7����k&MR2Q�L��*�p���8��{хl��Yᔙ���5���Z��^smʢc��q�۪���}Z�9�"p�m�55�U0��ch�q�=r�ֈ�3�i�'n�M��7U�b+q�N個���޺>��/Cfx�y:i�^���y�ͼ-���콬���7�&~o�&9#y	�1'�:����������9]�@��%U����a����W�z�v�h�ՠ~\�zWh��+���������9]�@����E-��LK�\k�\|]����'z�� ����6u��>��Z��+$�|�a��"�?.v��[��kŀy�s�r��z���Dբ��p���#�%rvzsu)̋��Q�0���q^�!붷]+�g�]������/��{^,Λ��P��N�V�O���%\I1j���{^,�'
$%�Y%%�4��1]�z�Z��^���^�#Ը{d�i�`���`��8��� ��� �����+��n�.������	)�ou`_y��n���Z�`�_����a����W�z9۹�r�V��rנug2��lm�$��7�lE6���a���S5���@]qqA�v�p�쓫vY���\
R���{��)���s�R��_��%)Os��\R������@:�JU�����!B��")I�����R��=�u�)JO߽�ג��Oֽ���{-��F����R��_��%)Os��\R� ؘ��
O߽�ג���׽�)JR{GM���U��YUWJ0�A�u�Ȅ���{ݯ%)O��{�R������y)Jy���sF��[21٭kz┥'���k�JS�u���)<�w�Q"ηY�!-�h�seZ.��'�u���M�L�qP��FƧ�5���0
�d��R&ӌ"G'�i��}��ժR��_��%)Os��\R����w�B�ޡ[���j������@�'���C��d2S�߾��)=��my)J~���
f)C諾���-�kZ�V��z%)O����qJR���{��)���s�R��_��%"!l�&��T�,�I�U�dB���{��)���s�R��_��%(6<Q�� �[)P��R9�����ʻ��!B��!)J?�B^����JS�߾��B���F"�G�h�������M�v���[��v]��2�[:�X��$7��m�5�V�����[u���y���)<�w�JR��)I�����R���u�D �AA5�T�f�ZE�Ut�)Os��\R������y)J~��┥'���C�JS̏O{�7�Zّ��k[��)?~��^JR����8�)I�����R��=�u�)JN�h�˹����&��#�Λ��T�'���C�JS�����)<���y)Jzw�7�F��kN�Tfoy�)JO/}���{��┥'���%)O�׽�)JR~S� ?B��t����M� �-�д�m��i�<T�&�zzBcx��v�]`��gO\Լa�f�j��^�ݭ�-nMk3��]��c��}��_.V���%Pu���d��Sg{f�M[�5(�������9�h*\mf)�=csG�uK�����6�O�4vk�nݓP�V�a�7m�����ٝ��$���יλ> +���i��������ۻ�ww����sțf��k��V7�>+9�x��Q��v�ݳmv��Z��pg�����2���:g����m��3���\R����{��)�����*!/��J0�A�|ɪT:,�I����)JRy���R���{�┥'���C�JS����R�����FWu�h�f���)�����)JO/}�������)<���y)Jw�k���w�ۭ�o[�o8�)I����R��?w�┥'��ݯ%)��Z�"D ��jڪsE]!ZEU�%)Os�{�)JRy���R��s�"B��t���۹�� k�E5��Y�z���"��Q���]\�F�tsѮ��z1��\���v�JO=��^JR����8�)I�������;���qJR��ݏ�{���kz���������?w]�p��8 ki'��CJRys��y)Jw?{�qJR��}�ג���}3y����Z7�s7�┥'���C�JS����R��{�v���?w^�8��
7�/�f%UUWJ>")����)JO=��^JR���{�R"B��t��g̚�@S��$�-oz┥'��ݯ%)O��{�R������y)J{���┥'����u�`2��F���]�b�A7k�;P:Ѹx�%��򸖻z�6��n+k�)����┥'���C�JSg[��A�ۮ�0�A��[34�շ[�޷��qJR���{��)�{��R��{�v���?w]�qO�L�)>��u�}��oDl-�ַ��)���k�R��{�v����HC��8�E���&�!XM���ۼHň�#5��ټHI!����4�ͦ�$F8L)�g���7m_��$�V �<$t	1h2`t��������nY魆�w�3�OXKl k���Xa�h�x���0,h�/5���d�l �0Գf�c���LE�a���U��J�L�#BF��A-���J�y��M�L@W<�0��Ў��H!����M�������ġ�~�*Q��#�a�k�`$��	���{G���@l�`b���l5�T%�Ja�"a�a*��)����a�<��	����G�ꁰ��_TJ
>��~�16� ��'�K��a����qJR����C�JS̏O{�ݙ��e�lֵ�qJ_���{�ג���kﳊR��^��%(?�������)JR}}ٽ�kZޭ�eo5��%)O��{�R����w�h|��;���qJR��}�ג��������ݓ\�*Us���-�,p���e�����s6�1��e�ݎ|\3�t�Q9��qJR���{��)�{��R��{�v?���R�������R�?v'���0)UUP`Qut��!Br��_�%)?w�my)J{���8�)I��Q�B�������E�I2����T�'��ݯ%)O��{�R��$�w�hy)Jw;��┥'�3�+���q��ג��B{���8�)I��~��R��=�u�(I���4*���2M���ג���Ѯ��ٛu���{���)I����R����M?}���~��h�{�Q�_�f�����Y]����ڠG��6�����G���S���Kߞ��sm�ڷNzC�JS�߾��);���R������\������JR���w�ky���e�lֵ�qJR���ݯ#�C%=���)JO�Ͼ��)�{��.���A	���˪��.fB��0��=���)JN����,d�q�VD �A���!B��M�
�3��s[��� �>�>����s�}�)JRw�{���K��}��({�g����Z�Zֵ\��ox>JR������)G�/��?�}���)Jw����R�����py)JuT=��޲�k`6��e-�0��i4Y��������l�<��e�kn$��"�l�*�],ˬ���g/[�a��B��Y��������(ٺnzaJ8:+	'F�۵[��\OmNۖ@:��O�y&l���spƝr�]
�Y6���v[���m�
��s�ͷ'd�ۍ�I���"��!�;��N��8�Ś�#ƬGA�^ӑ�(��������׻��w�|�u��qu�x�Q�%�����6�\�/g�v������\l�?�&����}�q�?��m�u'��my)J~��┥'g{��y)Jw;��┥'�3�+���V�7��%)O��{���JO�Ͼ��)���k�R�����y)Jw��ff�ڛ��usw9�!'�nT`�)�{��S�`��￶���;�]�r!BM���5St�h�]ܧ��������);���R���{�┥'g{��JS񗧽���e��e5�o\R����k�J�	����qJR��s�y)J{������ow���=�4p�cf�mTe�!��8���zv3ɺwWntv����A�9��%+���fV�[��R���w��)JN����$d�s�}�?�]�R}��ג�����o�E�����Nf��R�����py}@]@�|���}ϵ�)JO���^JR����8��"��TBȟ߿��n�Cjn�G�%)������)JRw�{���d��kﳊR��{�}��JR���a��ֺnՔf��qJ_��$��}��)����┥'}����+/u߾��)?�a�X_ox冣z�ג�����)JQ�?w>��JS�߾��);�{��)�"���_l���+�9�v^�4n�V�dd۳��åtL�S��zq,������wP�����1G���R�������)�{��R�������y)J{���qJR��O�.�j���]R�h�]ܨ��A��ubK�I �����}��)�����)JO����|"�䧦];�oz�-�326kZ޸�)I���ג�������~`s1q]H	(
�$ 'H!WW���.�w�}�JR��}�)JT'��ܫ���.fB���0�A�	!'�oﳊR����}��JS�����>,����%)N�t�����ޝ�9��qJR��s�����]��qJR����%)O��{�R��_�(��t�uZ-J��MT�M�
�)b0$�O���Y��5�ۧz睤�;��?l_?��سV-k[������渥)I��ג������˒����}��H�C*B����d��dB��_v����1Jw�_���)JN�g��%)Os��\S�C1JOǹ��s����o[��R���}�qJR��s���¬d�s�}�)JRw�}��)�ѯs3Z���5���y����D�$����JR������)I��ג��_�J*��"C�;N/Ș��|�8�)I�];�뚙�E�+���Q�B����D �(�'������kﳊR�����%)O�=׿f��o5�7�3z�9�����,n8�.���իY��=qm�������1^U���ݒH+UUu�!w~�q��?w]�qJR��s���o%)S��Y�!.�wL�u3SWAr��ג�������JP���ly)Jw;��┥'���^I�Jt��}�e�ٽ;�s7�┥�}�ǒ����{�)O�ˀjO�����R����~��A�G�%�_�aE���Wv��J�!>����┥'{��^JR����8�	�(	��������JR����ȵ��7oY�f��qJR��{ݯ%(�@�L{����┥'��������{�)JRx���b+����~~n�'i�  ���T��[LM�Ψ�v2b��2h�v6‽:���sm֞��٫�5lQ���%�a����m�dL����X���.�s�6���[�����%W^:;؈�A��7 �F�a�'7 >�.��������p�X�g��z��[rp.�;r��.S�8�rz�=�m����Zp%t[�8��:E۲�1�ه$`T�c���~����߾������r���sT9�3�^�.�3�d�'G]=�z��:n�/=
N��\����o�AŌ�o��{_%)O����qJR��s���)�{����'{��^JR��S���r*�usw9�!/9׃��d2S�߾��);��my)Λ��\�)����U�53t�E[��[��)���k�R����v���2R����)JR{�w�JR���=��6ff�e�lֵ�qJ_�����ג����}�)JR~�{�JP|�,��~�\R�����ٚ�6kZޫyV�{��R��w���(�EI����>JR������)I�����}��a��S�@��N<H��*m=vRs§L�[�zN�؍�m�9��H��w{��5�ݭٽ;ʫ7���)I��߰y)J{���┥'��ݏ���){�ב"(��K�XQu2�UW*>��;���q=��h�i]H��!\Sb������R���϶���/�����)I���py'���ۿYaZ��v�#5��R���ﶼ��/��w�)���=�;�%)N�~�\R����fa�٬��Q��z�ג�����}�)JR{�w�JR��	�Y)�u�a�!v����ݫ�U�+Uww�R���������]��qJR����ג�������)I��N��*��Gbk;���S�f6�Y�D�z0����6m��=v�q�o�����m���>JR������)I���k�JR���|�\������<��?t�}�ٙ�ݖQ�Z���)JOw�^ĞJ^�߷�)JO~����JS����"L� ��]�ԩ�UWAr���a	J^�߷�)JO��{����0�l��t�����B?�d�ٿ��qJR�������=;�������"�o|R�� �=�;�%)N�}�)JR{����R�����!B�_R��WU+�k[��R��{��┥��}�������|R������<��=�����r�w1�ٻ����<]e�-ۨ:-�c�����M����{������ّ���┥'}�_C�JR��{�)JR~�{�O�A���;���┥'�K32�kY��q��z���)~�� �D	�JO~����JS����)JR{���<��!�O��w3>��l�[٭�{┥'�g~��)�����D� ԟw�_��R������)JRt�Ǻ�w��ދe��[��|*����┥'}��%)K�{��J��jO@̀�����5�}�y���JTԟ���S3vI �Lՙ�!-�{^JP¨ ������)JN�g��<��=����)JO#��V��kq:^ł�+]j�6f�<a"�vH�]sp)�� ]�Έ��ލՄ��Vv��{�JR�����)JR~�{�JR�����|�.JRw߾��R���O��j���v�+3{�)JR~�{�Gȉ!�����┥'}��%)O��\�B�
��@�XK�_�@��"j�x>JR�}���R����v���Qc%=�_}�R������<��/o{e��u՛25��┿���`jO�����)��g�)?w=�%(?��A����?�)JR{���>����n0�o[��R���w��)J?�?�L{��`���>����)=���y)B)�I�gO}X�$���F�7�j�{�˚�mv��3�4L��#�H`I"�h�i~R��$0� `1���g ?z�ņ�>0A4�&Bcor��[�&�z��	��WQM��~��ZI#y��z5�]˙`��D�њ�n�+��n{wu��ݚ���)��)�6�����%�&�4	�L�C2 :�w���La���^���m���8��BFB$w�Q86as5������lEz�S[F0כ�Zֽ���m���            � ��im*���i6u�(�4`���#���]u�F���aӬ���s];�ζ<S3؀Ç�D��z�`�������u����6�����%s��>�?��S��g��n����a��ݠͬ�g��E�ٌ�E��^BU�JC-���.�����Sdy���ت�i"q�wl�i�Sܖ@9:8�Q�� M�V!M[�(&��=MWKcd�����!(�L�9iE��OOI͝�.��>X8�+Vi'	c�����_�w]�/ږA�:Z��;/n��K����]��|u ��87�*�j��s�U�P]l.˳օ�Ju܊e1MUR��u�*��p��8�68�z�S8b���`.�;�\:JZ�j��lb�y��Sė ��;t�Jͨ��U��qs���+//VW��V���ݾ���G���>}l��/�Wm�-�(!�n%��ÞQ���smŒ_�/�wm�}l�C�8U�!��dy��L�n\冪����6tV�R�v#n��΢.pR�l�r�\�����D2�Wd6f	��]G�7gW-�e�<�R��n��s��Yz5�;<5W,pg9�lnV����G�9���YU[���Y������]�m�yt��ӷ��.'���ճ�68Gp���T{�
�L�$��u��i�6�Nf�c��U�����DMm0v��\�N�y�;n:�/Di6�uTcv�Ν�&�󱕇��e�qn1��o8�l�'9��]w؈���&.�ұ��q��
�֍5���S�C���s[]���Tmꗀڸy��^5�Ds��pb(pk�N ֑'��v��$\'7	��vM�ٞb��6�vi�S��I��-�@�SeC�4r�c�	��U@�� ���8�������Iيĺ�V��g�gc8�zѽ�M�S��jY�`�93��P��Ғ�4`CY�<�^6n�cf�f�n�V��z��O�ȇ}���������������q�������Pz*�h�`�No�|�\ 	���	{gT������fـȘnL�d`���;L�p�=4�֊M�z|�tMù���l����hX��T�,c�`�Ų�΢S���z��V4�^�7h8�X;X,�����wg�WBmۂ�V�qg]���T�zьnm�g�6ݜ��3��qA�@����a7� �4f�ܧ�-�� �\������JőuU�왷�Ȭѭ���2p�^ �y�5����+�ۉ۵�d�v�M� ����)��]�qͮv}v�5���n��>��swn�7��JR������R�����)=���~/%)O~�\R����N��n�he�Z�"D-�lė�(A��t�R��my)Jw�����)?w��y'�C����w�j�fovYF��n┥'}��%)O��xqJ~$�����)����)JRw���֌٭k6[0���ג��'�}���)=��ly	�&f	BP�%	�%	BP������(J��"��(J3�(J��J��Z3�(J��}ǂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	��k�֭������<��(J!(J��30J��(H��(J���(J��=��p��%	BP�f	BP�%	�%	BP��%	BP�$BR P�%	��ϯ<��(J!(J��30J��(H��(J���(J��;��q��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	B{��xy��%	BP�	BP�%	��P�%	BD%	BP�&f	B�
(^�]K��SJh���n����Mv�N`Ӣ�A����s�#p�<vI:��x���}lo�7�e�F�5����%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bw]��y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�~���(J��0J��(H��(J���(J��"��(J߾����(J?�Y��J��(Mf	BP�%	�%	BP��%	BP�'����(J��<���(J!(J��30J��(H��(J�ϯ���h�_άّ����P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'}��<��(J��)�)��c�D�F�a�1�0�	D�4%	BD%	BP�'3�(J��J��(O���<��(J!(J��30J��(H��(J���(J��?}߸pJ��(O3�(J��J��(L���(J!(J��;�����J��(H��(J�30J��(H��(J���(J��?{k3��f}��j7����%	BP�f	BP�%	�%	BP��%	BP�$BP�%	B{��xy��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�����(J��0J��(H��(��30J��(H��(J������(J��"��(J3�(J��J��(L���(J���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'�����o{-������g�	BP�%	�%	BP��%	BP�$J4%	BP��%	BP�'�w���(J��(J��"��(J3�(J��J��(N�}�<��(J!(J��30J��(H��(J���(J��;���8%	BP�'��P�%	BD%	BP�&f	BP�򒉐�	BP�%	����Ǟ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP��t�5���f6ջy����(J��(J��"��(J3�(J��J��(N�}�<��(J!(J��30J��(H��(J���((J��o���%	BP�f	BP�%	�%	BP��%	BP�$BP�%	B{��xy��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�����(J��0J��(H��(J���(J��"��(Jߏ��o5���owjW=m5�)��Ű�9��Zt��=�J�L��ɮ����|n��z��m�+?���(J��J��(L���(J!(J��30J��(N����	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'�}���	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP��߸pJ���T2�`�%	BP�	BP�%	��P�%	BD%	BP�'����^x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B}��kFpֵ�-�[��o�(J��0J��(H��(J���(J��"��(J߾����(J��J@J��30J��(H��(J���(J��=��p��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bw]��y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�~���(J��0J��(Ab��(J3�(J��J��(N�t�^f�n�ݼ"�{��P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'�w���(J��(J��"��(J3�(J��J��(N�}�<��(J!(J��30J�U���ت	�R��(J��(Mf	BP�%	��}ÂP�%	By�%	BP�%	BP�%	��P�%	BP�%	BP����<��(J��(J���(J��(J��(L���(J����[�#5�a�ֵ��J��(O3�(J��(J��31�2��(J��(J�����<��(J��(J���(J��(J��(L���(J��p��%	BP�f	BP�%	BP�%	Bf`�%	BP�%	BP�'�}���	BP�%	BP�%	Bf`�%	BP�%	BP�B"&B�w�<�R�F=�ϵ�����kFFk{���w�y ��	BP����x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'�w�pJ��(O3�(J��(J��30J��(J��(J���k��(J��(J��30J��(J��(J3�(J���~���8I�%��箉�"7%�ݹ�|�lu8��%��NK}��{�;��<����z��	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	B{��xy��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP��߹�(J��<���(J��(J���(J��(J��(N�}�<��(�(J��(L���(J��(J���(J��;��p��%	BP�f	BP�%	BP�%	Bf`�%	BP�%	BP�'�����o{7���o[��y��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP��߹�(J��<�iH��w��(JN���BP������)�%'������ff̈́n�ki�J�߾��)=��vN@|������8%	I���i�J̏V��f�AR���P�G@����p���=��pJ��}�Ӑ�?��
_�((����k�R�����k[��խ���y�nJR����┥� c�￶?�)O����qJR������R������'qJ�M��֭�i���<s���m�cqD�a*Dx����������lkG�����픤�����)�{��R����'��)��}ÊR�>���kvdfkQ�ֵ��%)Os��\�rR������)��}ÊR����v<��"���]͔R5wY�!'�}��)���)O��{�~��R��w��)JO?Y��Vwq�0�oz�<��?w���)JO;�v<��=�{�qJR�����R���׹���v�5���{��)JRy�{���	=���8�)I�s�`�R����D �A
�ȅ5�ݕSWwwwwww���j��R�[K�3sZ*�N��(�r6�'�^nѺ#�<�Y̶����mc��u����Ge�Pv�sk�!s���DI����K�v����᳹���������w{&�bw	"M�ӷ�V$�����ީ��»���U�V�F�m�sϭۍ���ֲ�8�n5\u�:�,��[��:��h�����-�k5i�VY������{���������Y]�����j/�v��ٻzuN��=e"�z.�c�g�����E�����JS��߳�R���;�JR����┥'}�v<��<�����ՙ��e3Z�qJR���{���$2S߾���)>��ly)J{��┥'��K����kf��o3[��)���)JRw��c��2S���g�)>�}�%)OS�/
Ua%�(A7v�!BO[���=�})I�s���)�{�R�����s����֧ff���)�~��┥����������R�o���"D ���Q�B��k]\��x�k�j�Щ��u8��7R��̝sX���77	�ѷMv��=�=}�wo�lg��g�JR����`�R�����);�{��P���;���qJR��ٙ���V�7޷%)O;�xp@��N�)>��ly)Jw;ߵ�)JN��vI�!���?��_ff���f[�F���g�)?�����R��?{�qJ~TR$��k�y)Q��D �A	���w(�hVV�<��� ����┥'��_C�JS���)B|��I�~�c�JS�G�~�n,��,�F���R�����<��<���)JN���y)Qg��"D ���NlUE�%]�s5-��zub��b�<a���۬�-��tK3����WK��w{ͻ���ЫX�ж�~o{�����~��)JN���y)J{���p>DB\����k�y)Jt��>�[��ȋ7��R����Ǒ��"����o�┥'����%)O;�xqO� �R���}�[�e��ٙ��y)Jw���R���=�-�fJ��CI� �"��P���s@�� �QV�*$���Д(J^�q�{�b�<����!B��}�� �鹚�ꩰB�e�\�7l�:D%Ͼ����7�ـ}�����d���$	H�İob�[Cּ&.������f�WZ��5�Q��ܠ5uƤ�uuV|���6}���~Q���ذ��:�U�hE�^��u��$�G�|`�ذ=y��%�%��r.]�j�IV��T��� ���ͼXr�P���������C�dI�)�����s�߳@ﯷJ�=���C②Qқ� �|��g �{ؽ�	d"0�I3@��t���k���,�D{B�g��M����6ض�����RsOrL�ҧ$�:G�_:�:6zȟٙ�'���0�bNN��=����o%Hv�f -�z�GIuuS )���ֹΈP�d�wb�;{� ��u��BQ�DBUC��nf�E��l�Ysw8��� ��ÔD%2徬�_�V��;�\]�+������)��� ۾0�ـ|�ŀ8�FӹE\�eU��l�9DD%ϳ���������g��v��iI$�I,�l��T�:�"���ѷ#̜Z4��ih�ʯmk�ے8V�-E6��<��Dn�P�����3��j�����t�e��J�.�QtVa�:��d�rtܩ;A���fw'<���X�pź�&7l��&$�^�N9��wV�sM���KT�;sV[����{�jٵI{u:t��&¯J��H���=�yCk�����-;��l�muM�\�u<ᱍ���9s;��7���Ӌpp\ܟ���y�w�|U�eU�$)���;��ͼX�^tB�H6���;-U�UwSd�MU�ͼY��L���������Xھ[��H��b��n&��`���s�ـl���B��^�t���X ��4�H�&F���g�b��=���@����DD%�""���� O�?��~�j�MU���� �/ww��7�f��נg׃����1� ��da�]l$`[��t]���[��v���l�r��hAC�b���mh��4�w@�K���}81S���\U�+����w����O�`���ـ�%�����Y��"���`��tH:!����<�KW�{��r����r�;��΄�)��Z]����"����}X�l��B��D*����,�~���gs�<�X�!<nG�^�M�������B�t�V�p��Ud�W%̢�j� ��� 脡{�}�]�w��hs�5\j&I �BS%3�=��e�N��u��D�v#q��o��<�@���{޸��x�MB	a��g ����@�{)�w��yB��C�݋ ��	�U`
i+Uuw�n� ~�s�|�ŀ?k�����/�0�C���Ɯ4������9pڏ�0��8txU$+�mt�C�,K��#F�z�� �x�M(Y$J�P`]�l60����h�?�2CF�[0cc,I'HQaNa��23�x�c�\4m�K!,�HPžZ�t.��m��"Im�1��ûHi~6�� ��.9'�9�4��A蘉�@�)࿕�:,�꨾���m�I� �	� �T��T8<~��<��h��4ת$�"���ǐ�E��I)�w|��}X�k���� �Uԓvb�8|drI�\�z����|��yh����T�84�$���c;:{[l�u,��m�F�-��O<��c�OH�%ajs.�U�hWuW_ 徬�����/�D/�������r��j	c����x�Z�n�W{^���׾�>H��c���&�pwv,��?/ЕWK�Հ~u����q]lq�%�
I�ϒ���W}�~�U���s�!! �4�w�s@���Ÿ�f�����~Iv�t��� =�x�(��5Ժ��N�}P-��ָ!����
�t�s^@�ӱ�[��Kv����K�|'1�{~�~u���6�`�w�/�w��so��b�&B'��۹���@��f �M�t(�;�Nfj��Ю�����o� �V�ÒJg��� �>ŀ5'��W�EU�]�rQ��N�]Ӏ|����� �V˫�2�Ԓ
�U�`���
�>�|��h\�z���b��y��$�I$�l��Xv���㶍[7L��Ѓj��wy8�;CYV�,p4�Cآg��~~�?v`ϙ��;���`틷).n{v�����Ǝ�Q�<lI���<�p��\q�+wJnsv�xy�"Lٴ�b�n��f��ː]��$U:��j΂�Aٜث6�����\��m�ح���Y4eZB����BZ<�AZΧ�;so]ɬ6��w�������������-�����!Z��6ÀS��!�7:�쫴n8#z�Dw���ݯ�D�q�b�)�;�����٠us���ՠw-�u���2#�4�΅	L�u�`��8�^,��G��%��=��37�����z�p��Q��DUo��� ?w~� _'.�Mc���7�x�Z�۹���C�g�f*�|�z��x�~� &B'��׋ �
'���:���l�=��7��.����F{$�<�;=�7]�\^^��e#Orƙ��ӗE哋n��̫��u���u�?;g$�%����GqW�s�``�nM���Vk�q �G%�E�?
��|���=�ذ��="ճ5*e��AR�����0�x��Q	D�����x�;�(]S"M8�Xd#����DB��}�o� �m��Q	K��h�q{[md"0�93@/m��t�,��l�����.�Ył���irJV{��[o������Nѵ�ɉܷO��Ӹ�'�DD(��	����m,����?w��0�ـ|�����@��x ��|�Ǚ�����4�j�?[w4��h�e7�g�f$s�D�ē�AD$����ŀu�D*I}jbID%��k��� ��t�E[34�թ.������� ��������K=}�4b;��E�� �ɠus]`�o�~�� =�x�9�%�穞Ҿ[m\]l�� �<=,H��Ը��c�Ŧ靊�ܚ�ny&x(66疟�����=x����u�`��ڦD�qİ�ӆ����o�ă����Wo��{�M�n+��6��0�;������u�B����� ��.�T�KK"n����>�X7|`=x�>S ���r�uR�� �� {������������h9۳q��8��s�O�J�Dj�s8}��%F��5�h��z�����Ь.K*�π�u�������!,�����c�/I2b�28�� ~n�Q
&F��sw��ot%��G�W�s�`r94l�Y4�w�}k�<�NE[�	�"AR��������, ~�x�/�?K��z��ڦDƤk��׋ �
'����}X��0J:	>SB� �w�7�Z�o{�]��Z�3��-u����H�q8�`V�s�v�&,�����'�!����5��ynv݈�mќ3�`��v��v��؝l��j�[r\]Idj��@�m��k�Ӹ�n��i��=�c��,�,���ts�nn笝��%
{RC�6�����X��'X��̚�eG��)���v�)��î�bh������4<68��0s���ޞ�ﺎ��v�skŭs[WV�;Ok��-�G�7a�p��1<WE��#���=ź�#L�F'&~ ￿������/���}.�@����׉	���n���_V~����k�X ���$̫��y4�	Š{�x�/-���٠^�ՠr�D��۰�D�ʺ��Oow� ;{� {Z��!(_�+�wߌ��WL��V��HWwWk /�z��@�:h��4"E�X�P��b����[[T�=q�l�\b�ѳ�b��J�I{���X��,���$c/�9���� ~o�
_�@~�^�Q�����yc�$z�e6f�=T#J�@�]�;Õ]��(/;f��L�{TȘԍcۆ��}� ��?DD����n��56��*��*D)��X�W�����߯ {��ߔW�߼�����윙&��<o����#��}.�@/�z��s������#��'Á��4�3:t=�G]�sh�r��no	y�t�n��{���-��:F!�?�g��s@/-�y�4ת$�&��B$�ㆁy۹�Q2�׀�^ �m��'p���]ڵ%\wuv��������B#�T��������{�*M�r|L#�ɡ�/[�z��@��s@/-��:�P��hA��I�Y4�w�}k�*���Gʙ����	]T#8��S� |��컟n�<ݺ�V�5`w[1t(Ty�[}�߿կ@/�zR\�/����[�w0i����Xހ_J�~��z\�;����}�V��?��hD�ߔ�~��~��m�~S'ou�k���ʙ�"�����n=�y�4���M
h?z�^w;�k�y�sy��m܄�
8h�l�=�}�b�}��.�=���x>��H��Tb����	����V8.��M�z����YLt�#5�h��Qɓ��$�h�@��u�=�g�} v���T��隸-#�ɠU�׾ϱ#����M ��o�g���F{/�$m�A���n������%2v�^��� ���dM��<��h}�\�4������נ^�S@�[���"L�Xa�m���@��dt��^��6�5��zz��#�	��;���:@���<2�
~�ꄉ�o��l����9ǖ�bq��	�	��H�b�I���9��
���@�:��\T�*�=}����ெ#��f�=ȜD�%T<�P�S�"A����m� m� 8m�           p -�����X�3& ���!k`xͷ�{)�
u�h�c	��Ű�m��7�w���X��uǲ��R�;���]�J��s�����m�����ٺ�(�B�e�٫�I=�v���0VX͘B�v� ۬)�����m�]����d�V�ݺul�nƝ�l�[T��]�N�1՞�n�)�n#m��=���F�K�l굼�N��5�a�t=�6����ӤyHN��iָaR�.��I���n屷��M=/8���΀5���������D��e�,g��WZ�bwH���tJL���� )YZ��M�UUpV(�fYZQ�/TU,F�cF%�UHA��	��vS��{,�5�oa-����y�-�Y��ո���%�m� H�wf�xޒ��jP�+,�:AeeZ��@U�lj�9�N��;(�g�rc��ܱp�'m��[�Eu� �8�]�T���9AW���*+���9�3�b��2+7�e35Kj{*;\�l�	ŭ9u�nSj�8)c���z�����hG&�[I� ��k�Rv�]a^�]W�,�4���1�6�3��a�y��YM�U�Aɹ*{�0�;u�*�YQ�6��&R8�Ġ.�u��5���v����������q��҈Si{<P����h�$��ŗ]���7lj�0R�Ӭ�_5Z�#=-;jy�0�Bi���nQy9�lʎPY㛴�.�.q�m��ݩ��w2k�vsBv9;.{['!�8R��Y�ڱ5��5�A�KI8K��8�\�n;CvAdE��P�&w;����x��:�<f�/l����^ѷX_I�� ��i+d��I1ɗ.��'d��[�N��v������f9Wf��ʵ�A�-m`�6�e�۶v���`*��-��vZ��02����v��KK5�<nhӜ���Mڙ����zMs�8��A�������q�w��";��C��zF�=�bDG��4�
~�+�S������w�w��k5� �If��.z�v@��Um]�����ukf8�->Y�p4��;�-n�E�#Y�t����s�d$7-��yM�V��ga�X�j� ����Bc��u�tV������٠��Xa�W>3�CnR蜛��M�7p<�ze޲�䀑�I9ɶ�dt�:�)5XM�q+�i#�l4{htu.�iT9��!�6^��;RAԟ������{����V�|�qqRr&���{ksf9p��=�7IW<m6�{z�gu˽�gp��v��wѦf1)���=�Xݶ`N�_�G���M �yb��y��ƌBrh���>�n��]��]�$�Dɼ��e�섉
8hW�zy�4.����>���$��1���W�yIs@���T�4	y�S+@����8�{^�������V���v�����b	�,JD�s���b�VwB���v�Ӏ�H�6�s`���%��y"��hA�����V��s���v�fg�]�z��j��3$����V�.s�q}+�<���w�*�;���ȓ!�8��;f���s@�U�w�j�;98<���<K��m�����t�;�h��@;ʸ�|�p�G�1�dt�;�h�@��k�/nSf6�"�G i�v��M/�F��ZsӲk�ص7a�`T���7K�H�H��I�~�h�w�z}��D%	} s}x1S����
.�E�Wu���rJ�6u�`7�~\���ĺ�XHa00n7&���u�u���ВJfw]t,���}�Tgr�Ȳ'��<rG�u��ֹ��w��	)�7Հ=<a�S"��I���ɠ~��Zy�4�.h��@9=Ux��k�1����Q�bgX��>�M���l�ٍ�q�q�۔>pk<<N<r&�a�ԋ��}4˽�@/�zfJ�98<���y����z[���2�� �Ӏ��:!J�*��i�G�8�ݾ��ՠҽ�K��M$��ci
�Ww�В�;}8����u��C�w��biM��3*����82X�fF�W����7ʽ�kԓvLb���qh�l�?.v� ����J��'*|3bi��Zs�$c���Ӻٸ�^�m�F,[X�GK�&����t%�	&�$�?.�� ���ՠ����gk�dO#Bx���΅2y������>��X�
�1qcia���o@��V�_Z��.h��ܷ��`�c5ÀԋC�{���/]���٠~��hV����.I�#����{O� ���}�Ӏ��1	G��'`��� :/^��mSe�I�	���tr�tjݜD�ـ�͑m�m:��9Rں`��:�c��"�]׮v��D.N^�q&�j��pf�2���ܑ��Sg�����G�ձY��[���'7 =�t��{yy�{wX��Pi�v��� Tv@�5�����c��ts�{����n<e�h�!�۷vI�n}1cd�Xo��k��r�N�v錶K�Z���V;��e{��h�+�[�浆�8n<M6dȌ���٠~��h��@��V��Is0W�cI>��>u�p�]���8 ���)�񎤛���'�&��@=�zh��Z~������Z;�K��6a�M��D�\����>u�p�]���v�G�FHI�^v������_�=��w��hYWX�n	H����qQ�].�

���E�p	y����ۋ������ �'"L_F��?Wڴ�h��<��;_^��ʢ��.P���p�]䨁��D°{O��ֹ�>u�s��*��.E���2䛒1)����_�� ~�s�|�\��w�NS�Z�
¢I���
y���=��- ����*�;bi/��/ƒ�m��%Zl�@��V�nJ�N���N$�p����ǀ�Q�X�z�tv�qy���nӲ�,d��x��f���0��5���	�h�@��V�T���]��U\���Z�:"!DJ=�|�y��@-�q��""p�L�컹��s�|�áD.Q!BQ��d��׀{���h���k�Lő����ՠ�4���f/z{�@�_b��H�G�Q� �נOd�@�-ZnJ��?o~����u���d����-�h6�r�z��C��l�b�;j^g�\]��~>ǧ{��i�=_���k�h��Zol�e\�*B|����h�@��V�[+�'�U�v��_�^1�%��ZnJ��נOd�@�%Z�y������,k@/�z�J�3��*P�`� �\�����^�h�C	���ɠw��h笾_�����f�˝Q���R<$LŶ�rN��;Q�Pd-��c��Y�WL��X��Ȓ�,2BH��ڴ��� ��h��ZzP�fFc�6�X�cZnJ��נOd�@�%Z3�Z9�dx5"��f��>��ֹ�>u�p�Qo���"m,J����<�NΟN���S=�׀�,�~1bO!��
E�^�ՠ~����� ݭs�djP�������=��;��������k�6[�n�r�0x�&3l��T��{[۝o%XԨ�w$���z��t��+��t���\�몁���C;;K�ûj �H)U�۬l\��	��X��v�F������S2r�8��gt���'u�^�yO>vM.�n�i6N�tI��:mdX�W�v���oS�/;�^{i�������%�w[Y�u���\�-w�����ǽ��ww�}���6n�[�/`y��`Y	�x:$C>�gkG	�KE�6��ʐ/�n��K����-Z}k�$�V�fJ�	��+m�0M� ���d�@�%ZnZ�	~�L�p|c@p�y��d�@�%ZnZ��נN"r\���K�Gk@�%ZnZ��נI��N�.��7�b8��cZnZ��נI��̕h�ٗ ��cy"p��	2@9���f2[˞8�]���U���qS�`��v�qT�u�bƴ�נI��̕h�*��E�֯$���*�����s�S �*?5w��s�y�^�9Qyl�eX��<M����"�/_j�;rU�ֽ{%ZlM,ϖ,�c1%��ZnJ��נOd�@�%Z�y������,k@/�z�Q����O� �ֹ�9%�6/��Ps�En%5kc37zC���-�l�]\�d�c�����Z6ݖ[��{O� {Z� �ֹ�������@����D(�x$d��h��s��S'��N v�^��s�n�4<���ы#N-�}�@/-�s�2��~nb*c�y��&�h �?'��CA�f��6b�~�'��K�J�Vr�٠3HJ��diV	t�p�@�U��1p�PH!,L@�!;6b�$Q����	�e"!����$��(�p9k����&��`F�*�ִ�Zth���h�D��p3ب�6�`A�MAOC׊tN�'���+��*gAE�I\%	��{8����Z�*r���WPEM��~_�B���~��w��ֹ�>u�p�Qo���6�%WW ��N�(���O�{����w�~�>�270b �6,y�y��ۭI�^m͵��	��N��t�Ggc��O<��g�M�̕h�*��_��PY���=lI�`ס4�)"�?Wڷ�ϲd;{� {O� {Z�?BJdq;$���� CIǠ�4�}�@�}�@�����h�a2��7&�����NΟN�����B(}� _�J�e����zw���o3�#����2U�uIs@/�z�ՠ~�fU51�H��NF����ۋAy�c����哳�%�y�q�����:w�M���F�_���@/-��ՠ^�ՠs-�V-q�,��������I)�ΟNΟN����!BS'4�}�j�H��Ī���7��N �����}-�`ou���mK%UQb))���ֹ�>��8 ���%�>�1����{�&у��B%�H���� ?7x�Z� {Z� ���*"*t��!M HT�`�� L,#�gAu���Z�o{�����VصI��U�#��Z'f70�K	ur8K����n�{�Y��zQ�KZ9��ܼz#�by��,c�J���pb���E�-��.���-�q�{d��gp��d�ps��5�����֖!ݻx�Ϲ��cθ�xM�\�Brub�5����k<�=���.����*6���	��ƧO�n�<���8�=@��f�j�׽����ɏ����֡�����VՔ-�f7H/H:�������ݣ5���wu��A'3���;�M�_j�ֹ��K�:}8�R:�U��m���̕hd�@��V�_Z��g���͞�\��q��FL�E�y���mk�?B�;{� �Ӏn����2)��,�8�?�>\��h��M�_j�/_j�9��!y��H����9Dy���t�p�u����躭��������'��[hWt�n|z�gq'n�Ín�=����1�w_�t�p��p�u��_H�׀�Q/�R���RS7s�=�s���""�dd�Ȁ� �30DV���}4�}�@��I�`��,RE�~]�zyl��|�+�Z��Z�q��5&a�i8�?��	L��^�O� {Z������*Eo��DDܚ�ՠ^�ՠuIs@/�z��\��H\N�ːn������)�[��uN,m�J=��9��1AǍ#&I"�/_j�?.�� ����*�$�@����q�5�uIs@/�zfJ�2U�s-�V-�n<� ����٠~��%%�Q*�ֹ�>��X�Z��٣HX���O��-̕hRW��� �eB�x��&bR-�k��"#��W��׀}��p����E۞Y݊��p�Xq&�����]v�������s�7<�)�5�ց�%� �W�vd�@�%Z�y��5&a�i8��٠~��Z�*�:���K�D̫�����7�vd�@�%ZT�4�^�8�r*�	��|m��[���K�W�������A���.(��\Ul#0	G����s9��L<����LiŠ~]���w�{k\�k\�	BR�������e�`.:4/^I��̒Ex(vv���w���s��f�<&�G!�����M��V�fJ��nhH�٣HX���O����2U�uKs@/�{؏�*�p��fJIL�`s�Ӏ}>�`�=���hF���4�mhR���^�钭̕h��#��4��A�#��f�ξՠ=�s�};����J��5^�2�� I,�s���n�%õӠݳ�pὢ�-���ArOnH�c�֚㗖��p��N�S9M�����s��XLz(
�	+θ|�s�F`]�[zƗ���n޺7n��'��Mƌaeیe��j�cۑ8���6��۵��x*H�u�c]q���}��E�q�Uz:��]rN.G���Y����~{���찋�V�=&�����Ψ�[7M�=�P�-�h7]B�u�׶y'�dB�0�``�Mɠs��h�*�k�%��$�����ܗ1���|m�ޤ���-I%ܒ�z�E��RI~��_�{j�3������'31�Ԓ^�gz�E��RIv9Wz�U�V�$�2�W�d�B�|9��/}�>�1~��z�K��˽I+��Z�K�%��$��?�^���o8�1�$����z�W#��$�rK��I:=I%���w����\���r�[%ä�<��`A5H���a����an�,7\�^\�^أ��I/�_�Z�K�e��$����r��$��I��� �X��jI/���ߙ�>���_�c�ԒV;Wz�W#��$�~|B:���3�I���I��RIw��~������jI.?_?ߒI\h]����1��ǩ$����I+��Z�K�e��%y�J:=I%9��.6��ǘ �cmw�%r;�RIw,�ޤ�c�Ԓ]��_�$��3���7�����JS�Ӣš؀P^xΛ��خ�J鬬��5^wny\U�땓� �?���������r��$�GqjI/r^+��6�k�>>1��RH���I)�*�RJ�w���Ys�I+h����%������ff^���陗[n�&b.%�g�,� >7�o���E�4Ϛַ���$~���$��*R�q�����]�K���}��.��I%��y���E�ԒR9Wz�W#K�ŗ�f$���Z�K�ڻԒ,tz�JG*�RJ�w���꿲�pHdc�h���!tō=v�qw8���L��#�ۣ�cCJ7v�8mw�$X��$��Uޤ���-K���ߒJ�x.��}2``�Mȵ$�y;W��Ͼ�1�����$�=/���$�e�}���J�;��̉㑈2BH�~I/+?�$�\��I%c�jHS�Uޤ��r�l�$ČY1�Ԓ_��_�$�{���ff{�~�<�34���E,P�H�!2�B1l�$�)BJ���<�u933:�R��Ws7sǟbmw�$X��$��w�%r;�RI~w����I\�.7��o�'����}wط�ƌ�^�ݢ�;��Ͳ�t��)[`xv��y�$�}��8N$����_�$�}��I%ܲ�z�E��RI/r��M��l\mw�%r;�RIw,�ޤ�c�ԒS�Uޤ����>1e��.,o������/e&��g���6������jI.���u;Nf����/e&���'j��$��jK��'����%�O}O�L��MI%�N��
�����X��0
Z��Dl$�!�"Bv�G���%�ڹ��9�)�p��1���a��<oC�9;G�q����k׺����8~t�3��P�G��R燆��͆��S3�1���&�Ĉ���ܜ��w�N	�H:�(+�`�%�lܮ!��I1�Ї��:@��ݫ�	����3�8�t3�'��@z- _��6���� C�)����ٙ� �^��          `$ �,��Z�Ay��wb��ٶ�܋�9BS���`N0J��m�����;�C��tm�N6�%2;�i�u�j�/;�]�g.�`�1�wL��Z͠�4�48�«���+i �d���[&�R���\��Z8��EP N�Ƚ�SWm�Om�]Xr���V��q�"g��6�h�m���tk
�;6�]R�^������D�\��R{Y��t:�r�4�d�����Z.��������d�I타�F�üŨ�^���`f�oC�Y��hE{J��Jg͚m5�a0	b`�]���0e���YP{* K�ddȡ5˖jy�B�@-�Z�t.ʥB����:�e�^�$�h��Rcs�᎖6H����W�&P��-�:��+��å`.�P�*�Bh	V�rct�U�t�j��.��-Yv���<�N��^����I���w"�y'�ᗏe.�˹ګ�8���`��/�%�˻��مK�ݳ,�<��� x��m�`�rU�;�Kڀ��s�է��[��l�Ӓؖ���@�zѰJ���"մ�����2�e{t�a��Gpy&�E�\�Tґ��VF��;9xUZ�����́���p!��ٺ�����sv½�O;����aLG'J-F�c�ܐ;���#'��{���hV��e9+���v��=����.s�.�NG9�skh���W��畽>{[�t�v���=�p�v�+C�٪�gl�˷L�F�ȕ͡b0��ݷR�br��\�Vpv��ԝ)�;v�Sd������z�b\�։6�Թ�n�b�Oo0عt��Z���p=���6Iyg��G�($t���kG�^l�f2�ml[�;�`�e{b������7X駶l�NՅ�n�$�әd��/	e1�&�!7`���/�]U�qe�����u��{��>��{��@�4�E*���ԃ:��Q�x�Q^�O�OEC�Jz[�ޭk7��H��K�zI�e�+@Vy#J誩�y�%k�ӑ��L�m�hc-�U�[v������V�;t�'��]��]<时we�1֝.� [g�g��ۖ7F�����N,�z:9�D�0]�<$l,�g	y���r^��\�6��ڮP�s�I�������=�Y�山��.z�;%e&ݞ��o�6$+����w{W��h���O\��YѮ��6z7)�BB7�]y5,t�[��	��̉㑈2BH�W��������ߐZk�L���ľ\|�ǚU�4\�hd�@�ֽ�ۊ��"R,����Wڴ�k�:"e��V�����"}J�L���M��n_�@����m��%Z�T)[cx6�G6��nh�$�]�_�O� ݭs�rMm��D\8ڵ�[�<a�����NYIe]��%ky�����Lk#�dn��8i����u`u�pݱ�/��u`'d��u�MZB��n� �s�
ABP�"n�� s�� �[u�5����?��6�5�IV������Wڴї,�dOD��p�@����m��%Z��hg]L���d��z�mz���;�|�m�����^����r4<�M)���5��9r\iv��}��۵��l����fg��[�x�)9�dǠr�ՠw������}!����9���R�S3A���k�[Y�hz��:���z�@?eGky2D2D!�h\��^g{�r��I�����Q��5���9l*�:�Rc�j�i,NG���dDD�����}8����%.�����S�m9�dR=�����*�:�k�?+k�;����n8�m'2̖�,��D�;q'Yw;[�=Zx���r[�XO�r �L�9�h�aV���^��[^���Zh˖G2'�� �*˜g[��
�==�X�wN�$eZ�p⊴�&��|����:���v�@�2�/K��/���Kk��1�ے�Hʴ�.`y
�+�	E�7�`ژO���X��X�@����"���u[s@�_j�9�}�dn`�Ĥ1,�
�$�u��6�,�XG�IS���	�_G�M����E>nd󍤸��Z^�4�nh�*�$��@�T�ό��6�BX�@��ے�Hʴ�.o����Ѷ�b�4�z<��h\�z�mz�<+��"R-wls�l�]`Kn�9)�[��vzG2$���p�@��k�?+k�;rU�IV�~�99.�1cm��ue��j����(W~�x4n6�ڱp�;&el� 8̮�M��v-쵕���ml�2v�ꐒt�ԑ5��"�mr�l���`��SX٩�Q�.�۸��Bs'G���n͔ilZ6櫒0ct�f;,�ǆvt��8Wk��km�\�^r�6���y�*�Q�G<[��Lnl���W����!�q�me��\�S?��������9��K�+�q��<Lyvz�p��լY�Ӓ�6���r��]P�K���$z��~��h�aV���ȗ����<k��c��%X��� ����>��g�D����_�jI0�I��{��ZW;^��[^���ՠ���2c���%���@����m��%Z��hJ�x��#�HIǠ��@�_j�;�c�gu��(��/�����f�MkC�^հ��([��7�4��yĘ��6�RX�ĕ���6�b�I?�?yh�aV���נ~Vנ\�íԉ�&{���{ﻻ��6"� tTS��K�IOw� ��u`:npe7ȣL	�����?�����-�-�xbꤘ��|����:���v�@�2�/K��/m�31����1�ے�Hʴ�v�� ���ȞI�7���鵷vn�E�Oq��:r�7ly��l���#�[���ZMBh�	��l<��v��ۚnJ����`��fq���k@���v��ܕhFU�E*Y�A���m$���v��ܝ�XuP��pD!��C���qqL����w�ʽϿ��*���"fV�1�16�ܕhFU�E�נ~Vנ\�·V)�&IqhFU�E�s@��ے��^~T�&��d���e���#l�A��Ms����c��i��(g]3tNv�j1�hz\�:���v�@�2���$To�cG���6�@���$z�FU�yz&Q��lL�x��p�y�vd�@�2�/K�U�4�N�;�RX�@���mg�N�y��u��� Q�Ҋ���Z��/���7�$��hd�@��ۖ�Hʴ��B�c��I��;]�z�u8�.���;����l*�"��*�oH -}��V��;rՠIW�}Π,���~Q��&�>Y	�@�_j�9{
���x�Z�<+ub�`a$JE�z�U�ҽ{-ZnJ�C��0q�Y0$"���^�M���@��V��V��Ò*7ı������Oe�@��V��V�I+�?]�߽�ӿ+�� m%���	�S���U�9��,�;/V�,�/�ٸ�N1����C#t�9^nu�����K�Ý�j��}�^*�;nF�j|۞��{u���.�8�%���-�^q��˳��^�����Zl�Y����^�A�4�v�ջGN���;8�����[�^�m�>﯅7�mvKجmS��|�ַ����S�3[:v�p��������w�����r��+-�h�`�v����8��L��m^�g�ܔ<�������q��Mj5ګ��7J$���=��~��ls����BJ>��~��=�x��RL3A`�_��:p��7�������J&C��ܙi�,DdZ�}4�v��ڴw��@��&�Mߠ�HnM�-Z�J�Hʴ�^�>^B:݉��A���/�@�{
��^�ٖ�X]O�cX�8���4�'l#]�V��fv�����ظm��u*bػA�I����5����865�h��h���]�@�v��e��<��2A��r�������RTHX��B�P���6��Ô��wN����Q��3�z)�s�/�2I4_O�h��h�� �/
��LX��!MU�����[�� �ye4{Q���ɩ&��R/�w�� {���`��������U����N�W9�=��ŉ��XD�gJA�[����K:t�8ӣ�m���h��/�@��*�*�I��4��$���;�)�^>ՠr�h��@�/!+fcgˌmc4��8���N�/�ʴ� S?W�0�<b̅�h�Pq�����l?kc;U�NdP���Z:�xp��#.��\��2���؞tI�� &Ȑ��fZ�%,3d�ŉ#��0ӎcc����0AC�L��6�f3LL��aa�h̩:B�T�z����s`(��? �������PW�C�,���:"�/�:TC8 ��}��W�}�m�n�S L$"qh��Z}+�'���}������l�0�f1� �����@��V��ܔ�?w*�n��Q��XGGpe�	�ぴ:����<������H�v��f�����M����h��M ��Η$Ƞ�s���䒙7��0����l��O��&����R/�w�'� ��ye4�ڴ�bT�&(&�B�Lp��
g����t����
�*Q�}�ՠUʓh����i$'&�=���-Z�eZd�@���,�l�vl��vɢ;f�i��u��k� ��^ϖ)K��M�h���VZ�:Ա���78��� �<�_�=����"� L$"qh��[���� �����8�79�%2k(��w`<�2A�- ����V���_���-������ђI�ve�@��V��V�Y+�B�L��1a�H��j�9�­ ����[��J�}�֝���n� ��oL퍭[������l/*�i�vf�����̓���=���]v:�A�ip�&��]��T
�Kz���P�(��nEnK�=���֜;9ɝq��έ]�\Y�ۢE����<������|���=n���=q�ktu���P,��ܕ���q�KZ9��;>�p��6�s��8����N���ww���{�^W��Bظl�g�>{��lnY�eݹV��S`�&��ign�ٍ��lɩ��L
E�=�����@;�f�x�V���J��PM8����ҽ ����*�=g4
�Rm4��$����٠^;V��8�J�	��r�cl���{o�p毌 {��|��8�ń�	�Z/rS@/{f�w���ڴ�em����B�[i�\�m��z�9�JLM踼�ܽ��J��L�H��$Hh�l������䒄���Μe�=sH��	���� 7��\l/%�B��ڴ	k*��^�z�m�,x��	6��h��h��@'�� ����x�f�`)&�~������k������\���c�ŋHC�� �����@��V���h8�f5���d�s ���H�,��M5ʩ��\�Ӽ���Yz��ݵ�0O Ř�x$���zW�_d�@팳���7׀8��N��*��!auwx�79�'����o� 7u�t��i]r��V�e�\� �<��!$>�P��L/�����]Ӡ~���r@@� �CCؗ�����h�ՠ~��M��J��<|/���uz\�/�ՠwӎ�y�4��˓F!���919���qr�l�^n�ٙ5嚷Y��i���,t77@`�z��Z�w%4�hO�� �B��x��ebU�|���?D�{_^�o� �}���L��R���Ӊ!4��h�{^��.+|�[-�_jQ��>lI	ɁЧ��V�o� �v�8!(�1>w^�>^B.V�m�\����K�deZ�+�:���{�L���m��lq����랮���PL֜IM��b:m>#�x7"�} A����*��W�uIs@����v�^\m��`�l�5����K�T�4�ʴ�s�*�qf>���:���>��Xr�����gN {_^ {K¶��<h	��:�.h��h��x���V��]��^+���w_����?DB�������Հ}>�X�8��R��yt�ʩ������,���A�Fޤ�ι���[�6��\�h��y*�I.�b,�l�9H���n<IvM�Gn��]�G,Yxq��7X&�%�*ʩGX<��p-�G�,�1cLU��X���L���rb�:^�dͬ�J�N��,�mɶ8���ב�Cƪ^�9v��k4f��sqʉ��{N7]�nn�˺�V�Mr;g���v�j��\�IQקw��w8��l�4�/7=n�O�p$K�3�՞�q���:u�8�|�֎Iz$��<���� ;�Y�~]�zӺ��D(QHy�|`t�fP\�U\SBrh�{^��H��@�<h�+�'��E�ٍ���X�y�uIs@�t��^��%�����k������d㦀wҽ�K�W������l� ٌk@;�^���s@����wѕhKʙ���:���b��Kŝ���rgŲ<%ry�u���S��7�{t⇲����O�o���.h^�4�ʴ�K��^��t���"n� �w]g��"��"%�f�p�w�};����ϐ��Z�Y3Fi�ᷝ~�����W�uIs@��k�e�J�b�&���@�����u���]`~�S����=��fA�c�0K�c��K�W���2���k�=���<�c�0rd�&�D�	��q��<kgno]��k��[#͈-���f�/!���&����M��V���2������V��<+�a>�	 �z��L^���K�T�4�/.6��0`�ƴ�.hR\��*` ��:w{���r����� �砫Yı?�|����:���uMu�}�c��
g������v��M]�(S7s�};��Q��ç�7�~]�z��N�2'�B$����OD�۸��ɵrOM������'�<8�ܽ���=�Vfsx1������vJ��.h�{^�s.+[&8&�I��@;%zfJ��.h��o���H���$an|В�@��@�����ʴ�W�O���[bm�.3wXӺ� �v�8Ӻ�$���Eo�����{��>�	 �z���hd�@��V��%����#CZ[q:���4�Æ4��q�ӭVn���i59�er\��tնm��jͣ�ۮ�������#�7gN ѝ�z7�5>�d�h��V�#��=ֳ��:�����s���؀y�uz\�;#*�:�.hR\�/mo��ߵ��`G�[-��nhR\�:�.h�x��>cX��I�ց��s@����s@쌫j����& �c��^��6+��JN rTt�������Zz���	��od	ABD�@����܃���20�|ce�x�x��&~�Q7�H,�R_&	�IZ� lI�>�M.�P���M@��ӎ�]��E p��X��ۤ�!v��@���CR���D���7c���x����a�!RX%��>�P���"����W�N0�<9��#�f��� ��ӻ��{�N�{���-�w� v�p �          `$ �%�!l�Z�Ws��u�RY�ܫvL���j�P0���3�:8�κn(�i%��B,���.˒­��ƞwd�%��Uش��d�ܒ�Y�A�YX�� 8�Ǝ�q�'6�W���0n��e�Z۷Ku�D�N)�#Q���n��*�Qv-�]���٩�V���˵�x.��,�덂x+dn7c�Ku¦g��*�择RY�-�Ke�*���,f�Hq�D<mf�3� ۔�h:���o��-mM�F"�1&��q��閔�Uⵇ0�k��e.ܛK.��*���p�[����eڻ*l�T9�Xݠ%�<$47b��}�_8�UU 9Un�@Z#Y�I\	 �x籔���gZ�
��ey��ݖMV�� 
P�n5`�^�wg&�Q�.0ʶ��[ͨ
�ɉ�R�1�v���mmF̙_[5d��jZ�]�R���M������1�؄x�9M:��ƜJ�6�.Ǻc�d�X�g.àl6pZ�3\��n����[����8��0�AC�D���1˷X�&��Q�e���p��ә`��i�Lp(���۷:$��e]��`���b�RCF{s�I�:a�Y\�rrq�=/N8�.��kK.)=�;����qX�]v�q�.�9R�۬�:1�H�vI�4_f��9���i�}d��U�D� ��8�t��Wnq�eS��{9���a�����������` q�[O9M�3��m��݁7c�����e	����7��M�.M���7WGxz��l�b8ݹ�1��;�un-ĝ;�۾7���3�E��@vp�Q�k�F;;w7ͯ���+��Ъ�ޱ��P@G2��Y���n�*����	vZ�����완���2�j����:UZ��ܥr�.޼�y��7,nhJ��[<-J7It�nы�pX�m�{ykz�5��oG��@�G����/��hD�8����
!��ڡ�����l��@�T_w�ߧ���\ 	t[��*cj�jܻX��q�Mm�.�v'z�9ڑ�;N�yIyN{H�kf�!�����Rl[�2�ԯ\0��=nΉ G</��]�یݠa�I�g1�+���nC��9��]	#���� ��s�v͞��q���vL�cg���Gnsb,p��#�z��D�>�����a���v^uk�t��ٌ���[i/[	�t
+�;������ˇ'V���9����� �8b��S����<��Z���
�L����٠uz\�;#*�:�.h��"�؛gˌ�������V���u�};���D��i]r���@]�wu�y�:p���Q>���N������l15��6c�:�.hR\�:���vFU�Ds�*�8�'�/�1��T�4�.h��hR\�m�w���kc���)'��tgnzd֊͵�F�xYcq�x���Z�v�����7���٠vFU�uIs@��{h�ߤ��O& ������d���A� �4�H�*��NK�����o�k�l�Հ};���I%2�OOeY745�'�Z���@���%��2��_h�0��>�Kq�{��o���o�����Z�\v����#�r$�>\f&�hR\�;#*�:���~]�zoK�`�o'Ѝ�F1�p	ײ�͎�N�5���G�����ɖ{�-��� �1��;#*�:���uIs���}�~A�o����y��X@	���u�
"��o� ��Հ}�c[�*3�/F�&�����@��j�=�������4�,� �%�J����6{�`�huJ��1�� ���K�deZT�4�.hZ./�[7����o:�g�^{-y�uIs@���s��Ě|��f�t���C�\�u��N�a5\�V��˒��-Y螯`�m��4�.hR\�;#*�:�D/�ݑ}K��?.���ϳ=��-���@���@�ˈEVF�!� ԑ��j�;#*�*��}���>������k@�2��.h���d(�IA	(<���s�� ��<�9���2A�-����ڴ�j�/{
��ʣ�Ȓ��L�3�ӑ0玖趰2qv��է&��\�7s�1�j|�H��j�/�@��*�*�k�t�V��1�!�Us�?Ss��!L�ݝ8K}X�7:����E��x�pIH��a�9�u��
g��� ������J�U����&ȴ
����j�/�@��*�*�f<iX}K����b�o�p����� s�� �DBG�w{�w���Y� �X��t�G^\Z��ѠݲJB�lgN�Ȋ�v��t�.�څ����J�
�<q,�y��f$ˍ�r�S��F�uk��t	 � $N�f�u�g�J9[&��Btm��iN�t�;�۷���Y6��f=��J��V�/n��m�ќ�q\�;���ێ�.%#;��lF��l�}[��ҫr���9��vzI5�M���Z�Ҵ�������{����Y��j�[.��ɢe'L�;�ǳ��틃���	�x'9��=F24�>��ڀ=����,��@�K��Z������3r'�{�U�U�u�?Ss�?Ss��!(�����H8E�y[�^;V�x�Z��hG)i�b��y�_es�?Ss�=��tBQ
'��� �{7�Hڑ���/�@��*�*�k�/,���.Y�6��dJ\6M?��X����zM����V��Sv�V��K��gl�� ��b�i�y�$�\�އ��*�k�/���}�� �.s3�x��J����]d������`ծp��-�Q7�VD������`ծp�P�S<��8N��bu[�n8bɆ9&h��h��Z\����h8v`݋	���9��ֲp��V�W�s�ŀ=�s�u�cu9������(����=p����͵����>���g�c]#i�͸lm�@���e��̕hd��f$u�$���cn=����,�V�fJ-�[��^3���WrPT���ֹ�ֲp��	B� ��1ƀJ n�{+�/m��-��?ۍ7�7�����8�7X��`~Q��N y��O&<�i����*�@��s@�}�@�}��.q����4�	��^�͠�ڸ]qI���=s��I�x�X�cU۱7pM���dI,�@��s@�}s�=�d��N�V �\���ʫ�R�R����k��N��' <�� ���3�f	��I�c�8�]���^�lt�=2U�v��1��U��.��
ϟu����=�����|�"]04�PC�C���x-�<yRD�S�_F7&�oe4�ڴ]���f���eɍ#�:%�Q��n�g�����[�<sѺ��q��o;Mg�2a��rFԈ`�p�/_j�-v�@/-���h�������4�_�����٠[n�z�V�~�.��0�i�����f�e��̕hd��*�f1+�Ȓ@���h��h��h(IB�3��x�r)��WWhB��X��8.v���;{� z�,�������g��?>����j #��X��n�bW����춛mgT�|tv��w].�c���[�%���÷2�]�q{6�9����b�j�P�rWOlp�qĠ��ꩌT�N��������Z��f!�m�����j�Ms�.�Y��:C��8��q�[':���,2�6���;�m��d��n���g�[Xf�����j�6$,� dl�6�u8����wwu��W��,ɜ��]��Bn�uv�g#՞�u��	%1��^�Y֋�a�a�k�ݺH�Z���h�@��s@�}�@�\�8G�HI����w��*�,�E�y����c����-�hd�@�*��^�s�·�H��93@�}�@�{Zyl�/-��-���Ѧc�q
E�z����������s��Su��R<�& �|d&�k�|�S���s�y���,z;d�==��b�ѵ�Y�33�������06y�X���T�V+�%wx�x�DD*��!G�"*"!)V��<��� ?;7�/˨�4{#� �crf���U�ֽ�]�y�>+�I�d�8�^�V�^[4�w4=���_-���N�c�EZ ����ow��9���>{t� �}�����V���TV��cv-��ѭ=�̅��u�]$��p7 �i�[������x���p��9侐;{� 5����#�H���&h��h�c�@���^,�B鯰�TTdI7s��� ��6�BT�)T��(�ƕ�N�5����������SG��(��� m�:QĿqh�R:Sb�!�?2�Nl$fx�L�چ(~G��=M#�h(%�\G�Yp1" �"���&A�d�$"L�K�SA:m)��"�FH���H"]�����0Ąc`�?�BVbS�c#��h���w�p_˾�a� �َ�@��0�:bP�X��3����2���]0�h|4&:O�0H	,�5��$7s)cK�o���$�>N�oal�_�IS�!����XEP�S���C�@/U~��)�G�B�y���D�j&*罻�x�V�s��W�N6ۋ�B�������8	D(��z��.�M���@�rM���Z/c�@/-��p���H�CQB��x
q��1���Oa���=���1�%�x����7)���ە�����:� �ۧ8 ���ID%�k�0ZY�~�'�f$N-��ՠ���s@�}�@�w+N�c�D� �����42U�YV��e��I��/��@��s@�}��w����+��vmPdt|B�*h��������U�o���i�i���o��*�/�Uh��@��s@3�*v9�<�$xbS�����1�6��t��v��y��;l��ô\��ܽ�?ߜ��1��!H��ؼ��٠^[���f}����h.
�L��N&����w�
J��݋ �O� ~ت�*�l��r@�rM���̕hѪ��נO��r�+ǉ
Ъ��$���������� ����.p��;O��2H�Z�d���� ~o ����P�!@���ӽ�~��}߉����|M���J�Y���U�pr �����ޕ�#�:�1t�i�b�	M��x䄸����mO�"�۰�uZ�YC�-b%+��yX8���ƨ&���u����Ͱ�;Wd����	�����Ո�uۃSK��ێ4m��S�WoUډ�gm��\kg�'��9�:��T(u�.,v&�H�&h	�R#�sy�7l��-�{ߞ�{��}�ԭ���l�H�r&��h��`ssV�s.lv�S����v1����'sn$j(���M���������ݱyhFx/��&����nM�������U��}�$v����QȞ c�4��-�U��@~o ޡ�꼪�EE�3w?��ztzנ_[��=rU����8�lp�6�Z�[4��������U�ugzY����Y �NcPje��X�l��t�r�U���F��z"���+��lI�@�co@��y�z�@�5V�w���.#J�a�m�@�~�9�6�,�@�]"n���j�	-z�t�/<G�ex��Ïƴ#Uh��@����J��gr��E� H�Qhyl�/��h�*�,�U�y�%�ĳ��xf7�_K��=rU�Y�@'���{��~���/��Ą�V������[TN��:��?�����w�9��͢'"x��L����h��� �-��x�����*�QQiL���v��� �����4\�hg*l�'UEX������w�?7��3�Q	Bj(�
R�^+�}8�s�l���`ҹ! rM�������U��@�ˈ�R�G�d�$�`u�p�ד��������>���^� �z�+�\�pۈ�/[v]��Z���7�H�u����n3f��wn�mhF��	-z����-Z���q�q�� H�Qh{l�/-�h�j�/�UhG'	q��نcz����-Z�j� �נs���QG"h��L�9]�@����*����+�<�j�!�(b!���ʽ�����͍c��_��l^Z���z~���M��mr�]E*��.��t�#j�)���Mʩ��m�$�-Ӧn4cv��ǂr8�(�0M��}�^[��=rՠ_F��"�X���c�co@��y�z�@��U�Z��Q
"dq;"��黤�hWwk ޮ������L��^�� ׍�&��>�0��hyz�^Zo�4����ڴ�gr��8�ǓA�- �n��x�:np��I(V{���{����v�z�t���&� .��v>�ѵqYGS�ѩL�f1.�,+lG"f���nM9��b��$�=5t1�:�X�;>H�7"�GWmR%�P9b t����mA1�Gm�]�w��!�8A��S�ǰ��7Q��v��c��:W�ƽ\�:�/���ZG�;�c�V���lq�פ�-��j�XK��R��v�ܻ5�B)������;$�t����~�����޻��}�>r�-XI�=��۵:r&[\�H\F���s�T��nky��Χ$��6�����=����ڴ�­ �נz��m&�6�8`��떭�2� �נ[.�@�Qp���ֱ���N/�{�Z��4{w4Wj���Z�I�m�$��Ik�-�y�z�@�2�)E�>W!ā�4{w4Wj�-�,��w�~�Iw{�h�VUv�nɭٍ�L�96�Z�<a�y ��dݟ.[�\�Fs-v��%�0Ɇ9&~�~��-�*�	-z��4��e���Ïo9W{���'��zD�EP�]�Ў�3�G C��������� �￷4Wj�9Y�+�c��y0$1�h���w��Z�c*�?#;�kp��_67&�on���Z��h��м.�o1��ªn��Z� ols�����}�h�zg��MǉD�2bp@��Ͼ͐_o��v�����Sm͢�l����s�>����JAL�π����8�n����<�Z���[ F�8`�dZ�[4e�h�*�-��@��X���e̩����׋ ��D/��(��FD)�ι�����6'�)s.j�$-�o��Z�+Uh���w��в��3�mhV��	���`t���D(K�7TOZ���;ev�Зgp6��Wa9F��vz�z��-nWc��t�̯=vԑ�m����@����ڴ�Z�gp�r`�>B���4m��9]�@��U��@�K��"RI$I`�s4Znp�ـ�� ��Xz���9�*�mH)���?BIO���� o���{Õ�	 PH H #�*8���iT�3���r��,���lib�`�c4K^�e���-��`�D&�����tT�]�z^8�lK[H�q0h�V���� p񞣇[�C�q8&��Jd ���?��nh�ՠ^�M �m�1q�U8�L1���<�Ι9���^ ��X�в��3�mhWM �נ^۹�r�V���.W�x�`ISv`rIBS-�^ϻ�M� ��h��Ϊ��|��crh��h�m��7L�{v��	D$�"?�%W��@U��A@U�W��_��(
��(
���"
�� �,� ��$� �"�2Ƞ$* �( �($� ȉ
�0�H��( �� �* Ȁ$� ¨$� �
2("#
�0�( 2��肀������H
��
�(
�
���_��_�P*������_�
���(+$�k%V��`�M0
 ?��d��-��    �  t}��     @    ��  � ��TQ �H  ��@ P�H@UP"� ��T� ���P ��E0      UA@3 4�A�}�|��{��{���ޭ�}�{�{�j�}z��iK}��-�O�x�zR���y<� ��N77u��> >�}I���ʼ�rk�Ӗ���%]�[���p�Z�0h�<QT  �  �6({�Yo!�{�� =� 0L  �ww��ܯ y� :8� �����  �   4v �,  �� �  Pa!l�(  � @ (  �� P �  6 4@�0  ( &� L  f �  ��<i�Ծ�����6���6< W}�<�}�}*� �l�'��O'^���om�����Ξ�=�����{��v�m�׵x�>��
 P  1� ������)�`��|�y�]y�w�w_6S���|���}�qy���x�;ݧ�˼Z�� s��;��Ÿg.���{�� U��Wmɟm��n�w�y�|  |� � * $� P��Yo|��z���s�oVϼG}nm]��v��Ͼ���\�>��O�*�n��x�� �x�������<C:���`����ל7���T�����}��{��Ƕ\��{ϳ�j� =AT��T���CS�Q�7�R�h&F@<z�TeJz�  =��I�R�L 1?�%�)R� �""I��)�@4�z��������}����'o{���w{��^�r���*�*"����*��PU��EAV
�(��Ї�����t��0?���#E���%q40 Wt5� T��/�&o.gLeĻ�s���Ϥ��Η�L�B�.��hB�!C �s�RP��RYQ%	#	�X�5$�Ec�$	�q6�E"��P`������S�XG� jd! �,AF���B�8�Ak�	�Ť���$Z� ��J0("1h�
%��s��I����H)��H�cV������39�'�����%@�I�b6A�$bŅ|D�#\H�"A��RB+�%X�A�`U#BB5aH5�X��`�"aT�%e�!
�J@���c0!VdL�9�ܝ���O9��(H����K��O�#u��R�S%3ؒ��[�/����Ƹ���jD`R �#\M`U�!
��" �,Y����g��G�@*�$,�f���!���9ĒW��.s��k�y�3p��.��6I\x>7����|�@�8YLaI!3�(`�i��=�y�n���鯾������}��U�)�lFi�o-x1�s����#s���"�S4ׇ405HSa�.�e0Ӈх4p�\	L��Ja�)������.ċ<)��������o8��y��<9�&�x��$�s�n�)����4�'�q4񦆍�<��s�6���p�n;�g?L5����>�����|�}}���5��%�'7��k)��
���@�#xB��
���Fo<e������U:����8,
k��I	���bǌB,�a�LO^��\bB%L9��&����P�����<�:_Y�39���|��r^i����#<�ݸ2���ɜ��g��X�o/5����GaL �xB��Kw�z~��T�zI��J�%.�1���	-�+$-el��@�d ��)�J��([��u�Q�"�au!skecv��Jk�5���'�8~9$a]8g����)7k��<ٍ��HE�20����<|`HD.�M���~ӿ������s�yo��OIr�K���N��BRBHBDb�����?t���9!'!L�d��y������h{��3�?SK?d7�|�.��!����oH9(B�߈���B�o6�6f#L%2A�e����(����?0�4�������뿎������_߸��.��_^B��3�0�{��K� �N2�ɚO��<��~�j��Wo?�8�{�ɬ�c��+
��������ld����!�*jJ��A�2�!��@�.�H�0`J��*��pyq�f�!��2%bX�����6`BV-�F�{ǝ��&�/�#	'��������?,�����e�9�/�a�%�m�v�v�;u�g�:�:��{�<Zc�ư���Q�g$��տ��
d,��{���Q�Oӟ��CR �bVFF!e"��H��X4 P��� �IHR)HX[K3���Os�����0�\3YL42Ŧs\�ݻk{����� H0�$F1 A�Ð�,�Ir&Ӎ��9��a\!���ێI�i��5��!a�F��o%�w|L��k�.k�H�:�~.�3O˞}ه˾��sκ��Y��Oza�r�}���c�rfC��؞���~��4��2�HF�E�
yga��r�\��������$"� 4Lt.sy��_8g������r�0#	��˄����7u�t�!-	t̑�2Sg����d��3���\5�����o��~�fL�=�5��X�T�8�7	=�����^�V_	��Q�ԀXW9����m���ס�Wȱ����!sx��x��g�������a��L#\
FB��PІ�	X����#\G&��$�`K��B��|�)/�˄(gV_Y%p#D�1`$t�$�w�������ǁ���K7�p�|m3�4�$
�r�3�����oX\0#9�HHE� H@�$8$
6��0b�=���(�(T���d��w��З�柉s���2��arq��*c��	�m�I$��d	BF�4�4(@`	qB�m�a	�!q���Ie�%6�y���l)�s��6�[_!rB3���y�ӆ;aNr�S�Y�!�3���S3�%,,ajJy�/�l�d�$��4�H��H<EJA�р�b��`�T�"Pp�C(R6�1�P0+$�V,�Ab0	�@`5�@�DI���A`P$��
�Q!X�V E`�`U H�"A� (	!��(R!Z��h� 0����Z��a[n	Q�bF���X[�ā0�hD�0�`�	R�����la��J8�j�#97���p?k)��F�I�Jd5��\�FRcd#lÍ���J��Y0�$. qHU�N\���p*�(RJ�R�e�d� �$Y	#c%�5�����7�NN]�����az�\fs�}��NT%��@��%��_3}��.m,��o���J���i�lp3<��n���i���q�XH0�#H��{����8�`JbK �2xy��0�����sw?g���Ě�d���!sR\�s�a$,<�~<�s��˲Iԃa+o(�±)$�*C���g/�y�	�����M_eH�ԉ$7������̙�t�O<�=�36~݌[�5�7��?Ƀs�3<y�<��
d�	��xx��10�HZ�i
0�H��(B�*1Z��D� �H�RV$!i��`@��e!�P���<�6y�&�$J$` "�F�$�5���
Paw����"РA���R!P�L(ьB�ĉ�X6$�4*d�	#Y D�d	p�HS<e2��P�����S'90��C�ͼ`B�M"c �B�
@�!! �%�,` XP�D�S06B�I0w��Ƹ���$(�* D�JF�j,a�
��h��(�Ɛ*�#�T�<�e�?XD�����bG���fw���%1�y��cU��BHԅ%��
a.�?��,�O
�Hx��(I��B@���7�sO9�ن@��BT �hKS aX�2����顾�)��F4XD�@,R�@�V������]�,�L5v���� P$H$���}3/�����A�K<�c$i)4ӄ����q����<93��8'�20HHA��B�,0�@%�)���C�d�?O��������&FlI;�ө?+�
�P����`ąe�aYny�8D���t�<�������A�H�ȁ� "`Ċ@xt!���7�I�~$�s4���Ld�c	F�V"?g3�V��\7��������k|�~aB�#_=�
F���������+�!"�i���Ӛgwb3_�3Ý˽�g��_��$#乼�R�� �"~X5$�� 1��Y��]��}�<�##��%�+��%�Y�ӒD ǈ� ��,���B&d��F�j�k"F��E��p<?���A����Kl�$@�$Q @� ��~�+l���ݷ����                                     ���                               [@     �>                ��6�  m  &�                                                                   ��    �	���]V�^�9�]T9,�[[*��R����-����݉�pl��[@ [d㭭� $&� hm�m��t�m��Hm�r�  H�d ��H�� �"�m  �&�m���֏��  m�u���m�ۭ�k    �����r���� �����m�^Pn�mċkm�[@6ض�m�l�m6m��ih���E�6Zm-� �ޠ6�`9VStV�����#Key��Z����8#  -6���&�i3m�i��[U*��q� Sj� ��( [Z( [t]�f�L'C�-��݉I{(��ڮ���V�8�>ڕ�PK6��&�i؝$pl�Z�J(R��2�-uUTJ�@m������jͭ��'[l�T�ee��v	h�@����К�!�h�&�J��O+S��
K�m�
e����2b�s*�W���w[�btP� �2�kd	Trѩ��(��9��ӹ]v����@t3�t�L���j��^&:Wr���` ��]NtMu�kn�Ԑ$  �� �ݪl�2�)�A�m�m�m�����z��i�l	&�-�6  H8 �4Sk���6�kc$v��Ma�lt��� @#���+�Vҡ��ʭ-���*��mU+�4ۯ!"�['\��kX A�� u�n%-� #]���e���8m�v��g���m� pY�l[M�6�jQU��[+U�u*�Cm�� �����k������  -��]6[I �  8qm 8��  m�_�>l -���AJ���a��  -����  � 6� ��b��N�VW�e]��UT$)j�U�ڪ
H-�6nsT��dm�ඍ��vŴ �ˢհ� U�UWT��c���U�9j
��:���   �/6��    :@m$  	    -���	E�@ m ��8��F  ��   ���� �Ŵ�      �b�pm� ղ@�� d���l$�U���@�6׺����  �-��I�m��6�$i���$  �I H�l	��6����3l��핊��6u/+*U@  ��%�  �b� ��� ��  Hm��  ��`p�  �  �` � �k� 6�m&6�  -�$� � 8 N��m�  �ԙ"۶ɥɶ�km�	 m��u�ɍ�`  
Pm  �6�8$   �� � ��:�l��1US���L��m����0�  �-�'�i ְ  p 	� @ �6�v���g#�P��.�;UT��� Ү�WT�   p p   �m[��״�Jľ�`�DS�W�8� k�[N�� e��ڤ -�Y;^�9[���O�zմ��&���=�f�s��Md{��md�hIn�e5��t�̯S`6���x�-�)-U���le6�d��R����Ϟ�|���;����%M�yڻn��-ȸM�Cm�^y�@MO�z	]���6�rˎ�8���QT���F$	$XC��4r�*Wf��h��6�m�r�,�r�Hm�^҄�l�(6ٵknp���j�[m ����g&�+o6�f΢Mmv������6�#�gC���u�n����4�m�����$l� ^�^g[|�͋��`u�Ph�97AkZvѨ�g8�yV��-����t2����#�Pڨ#��kkh�r��mP].�v�pmW�˕
�4�!�E�lҵU
2ML��i�ZmT�T�\�ٴ�L�#6�mi+�D�uٳүV�v�(�U8⪺��t�T�veV���m���-�m9 m��@9u��U�G�c�GdҲ�q�m��   K/�
�i��R�,vp��G�sR�ʀ�]UTU[F�s�Go��}.6����i��-PE�&����k�s�)keYV����;�~~�jX��eT�-lګ:�ؚ^g��HH#<�UmF5	�89 m��an��Q��^��x6� ���@X�Q��m�H��-�\ U7�Mc�l.�D��p^�u�kR�l6ۍ�m��s̫�J�c�j�e�vj�d��ԯ7:9GTf���gD��A���ƛ�c� ���Tn�Mԩ�xe�a^�v�ڮ� F9ج�*N�F������ҧIp<m��@r� �l  ��   �(i1l��5�Z��%�;UA ��$lM��4����^H L�@ 6�  l�  h [vۇ�V7Nx��L�����}�T$� l� m�� i�Ͷ  �m�����p$8    ��   س�	  � �m��    m�}����� :�ɭ�h��D֙��]��iUyovj�   � m��ׯ0 �  ;m�hm&��$�[@���  �8A�n�ۭ��`  	h  m����mm�sڳ#u����m �v�ܒ��%����� �`l  [KhkX&�ۀ$ h ���&��T++N�k�)� ���$lm[@ �%�v!���lf���g�
�V�-�3 ��:k�,�z��8�6�x%�Fi���XŴ�M{O]Z1�U�
�m�U*ۇ��n��I��`   $
�K!�A��u$�*��}�bmp� �@�	wX�f�th�N�-*�)<�W@R��UG�E�6�m�v��6�դ [@^�H�vհ  ZNٺYx	��c`�M� [I��8��r7�VS&�)�"���3�\mN�WJ�{��*^�e[�[r�p��X���.9Ln���0���,=��OF�<2s�8=-T�U� �v��0-��-��t�Fض�ٶ�  m�6�ݸ���֛���l�Ӷ躣��k�� H����I6�N�Q�l�lv�Fk&�%�Pݶk%�8mytX��fɦ�[`����  �ݷ[\n�$���U@R��Q�)���,�lm5U*�U{����#�m�MS��rS�[�F�h
���uUl�uo��|Yr�v[˭���K�IA ��Q%� m���i!���`���Y���i�h
S7�yL�UYV���7�iX��bI�Y*��n���r&ñ՜�5� ��]5�	  ��t���Pڧ&f�)iUV�)j����m�v�]��0-�u�5A��nGg½5�j�5�jw:Z�M�k�5�<M�ǋl�-��nI}#d�x��L��[q��3{�ͣv[V�Ϭ���`w�{o/;:�n���n�udc��V��6횶�AP��c�Vݛ��t���[hU�M�)rƅjVY�4"�[Sm5� [��h�i&���RI&� pD�6�Ͷ ��I3}�>@�[u� [@   ���� �e �m��K3m�Im�i�`p�J   I��h�8 Xm�`/Y/k�m  �5l8-����6��i��Ĭ -��ɡ��j[{H�I���l$����D�"�:(���׈-�r�1�ӵ��p8�EGkv��W+2�PR�s�j-�+U*��l6�&&��kZM}X*ٵJ�U]��L��� ���Δ���+m���s�$6�*2��  	�8v�G��D�d�[l�\� �m�L���m'I~�*�vB�.gf~~�>�*T 5��{3�F�Q��jV`盌�B�J���کVցۉZ۔�j�C���l�sj�t״�7$�-�6�Z6ꀠ_O*�샖���׭��m����m�v�` ÑbN���Ɖ(��lm�í��Z����bU�}[*Ia3iz�M�P��Z 6� �� q�m  ���[sj�'=$�ɹ�ʓ\�:���HZi�AmÛl    �m[@H �u���l  ������ݵ��IZt�vM��w�UDQS�`'?�_Z���@�D���ʟ���  � `0$`�����x~T�_�R\�N*>(G��
��*�Ȁ 9�D<@��C�~Wp ��OU��� j'���A���A�
��B��N�O�:t@��R@������tP�(sU'��`��O�:��OS�h0�(h+�uD|�Q? w��` '��"@�<u~@}RT��uD�C� ��?0�)�����TU8����T_��Q�qE_D�gQ��q�=ڢ~PqD�#����/A���DEdEzu'`� $a"0c��`�T�U<CׯPҏ�`��E��(P� O���q*�:��� �^��z����vB,P�x�čV�%F%!"�b�d�Qd��F~��EQ|P�F�"��Q�?	 @��4Q� ��Q�US�� �
�!T
�S������*�Q�U�ER��HB�T�E��%D��"%U*a@�E������       m�      �`  �m             m�$r��d�/7���%U)��7��=��b���2d�,�S\�16v`B@P:��>gkUt�s�v�� ��h8h���@��:@r��"�'C4�ɮ�YsZ��E���g�<NB��tV8�*bOE�6[S�v��"%�b|;ujCkVt�dJ�������r�9�yv�<9.�*8�@q̯s�[]�:�{m�g)��HZ8�
m�["��pV��5Oe+��&ٸ�	庶��Q$� 5J�jm�{d�l�����g�$�bsJSm����T�J�j��+�Χtq�Ɩ��R����R���4�+ׂeZ�jڕ�j��W)��P<wmnN<U
v�u�X��FRy�!z��Rk!4��ݷQ�u��v�$M�ĝ{�6�kwcGpgru���IE{<V��m�M�
�#�.ٙx�;�������.�d�dk��L�=	����Nz�Y\�m�>�t�6�h5�)��1Lr�������w��kl5������w �U¯P$S�$�e +���������*E����A�ٶmۭ�&����j���A �R�RNMf�I�S[�� �����+P#R�C�H
�wmV�7[��W�2��s�^۶������ �9��Y���cFٍ��1��X��V���kix
��9Ʉ���콼�I�]�v��(�f�@n^oom��\������h�H�됶vI4����!k�h�sL<����h�MΤ�m����e�m��wA1 uK^� ��;�]Ǯ�(xj�@j���U�I�8�k)P�����c�et��I��i�✰ݎ�s$����y���V��ی�1��"J�A6���$�Jݙ{B�k���:���n�8�^g6�lpܰ�llPN$ʫcmŌu/]e{��w�����@�������
3�}P}E�<\z�������w�w������l&�� SW�u��v8��l\:jܶ�����Ì�c��c�Ļ6Z����K���6��wY�m�]A yp���Tj�\�����}ZxG�˖�ނ�U�wl9|ݶl��Z�L���v ���{WcB��q[���v��n�+���5���u���8:�^�&����r�qGn��6��D�CA�;�ْܒَ��nW����av6�v���yvQ�g�ß�8�n�;`���R��[S �L���?��>П���n}�BNL294��f�,T`OJ�K*`ze��D�ڎIa���sX����� �T��l��L�����_��v����W�YS�/0%��M��R������c �T��m��	b�y�\J��W<�ڽ��y����70�n�. ͎'��l��;u\�����]���&��d�Y�$�&Lx��"�I���>z^��$�� �T��gCK�p�8Öqݛ��{{�s��@�Ҁ��V*&�Q ���8rI;��I'����7$2�HXa��[�sK^0?=�R��#�o �9�kZ���C��]��0	eL˕0&�y�z���,c&$��c!�@/4����<����~{�JUU���HJu��2�Z�zrg�Gc\�ы�0u�N�f��t�J��*f咸�������`ʘuˬL���O͹�91$�z�w4�Y�^w*�9u�~���A�W�Ex(�	e� ��x�|%ꤒ@�$/�V!F!"U]ݾ��䓿��������IE$�@�ܫ@�׌mx�=mL����v�a���bL	-x��׌���-�f���R�$Odi4�D��H�$�NH��'8Ȳ���rY�6�[����כ���7WrX��׌���-�SKw4q��\���f�{m�*���	"��7'.��p�'��@��,�"rh[�hzSO�2�ܓ� 8���&���۽��7ٺ�&�Q�-������߷?'�/��iK�hv[�k'���91!�0%�� �T�%�SX��>���It�X���8hQ8�Wn�=NҞ���	����}`'�G[�ЎvnWP����/5 8���Ox?k>T�X9'f�Յ�	Lx��"�I�nY�K��K*`}��m���!���w������o��]�9� �SxZ���f� ��w���pD��?� 8���Ox?k85��[]�h,�r\��K*`ܩ�,T`Ik���2[�I$�I$�HI��  	}���6���µ�ɘk�!�7X�[y�������3��K^^�}��S����p��	�;^����ۂ�Х����; �F�r9�z�oM	.�m'&$tQ h�9n������h밳�ݻ5v�]�e��˷����\]�]�1��Ź�����HB�3ȱ��í��3p��VtG#iuU��xO����;%[f�ӛiS Q�[v^)����t��,���sbsq�\n!y(������*0$�� ���;ܴ�F��Ȅ�I�u�N����ܜ��7�?6����G`�wr�$�ӹ	mx�%�0nY�u�M �˱���m	�Д��q��	"��y�Y�6�.���b��"c��ɠܳ@�Қm��?=�%$�%�����l�t�;	���f�Y����+c���q���v�իA�zwJ[�ټ�W�m���_��m��?=�T���$Sxlv�,ՠ�w���p�˚J��uIZ��	�B9��_$�}��}����<��誮��ŕ�Y�����_��-�SX���׌	2�^����-i��n�D���"��8��@��� ��h�����j<Z�&�Q�m���mʾ�������-YE��s�����4�l������:�Janڧ�'�=Q��y[�%���`[k�,��[r��S@2��uD�xGDBs4�Y�ܩ�,T`[k��vJ�Vw	���rL[�0%���̹��+v�h[f��tAF�2/ß�y&�,T`Ik�,��zܩ�6CJ�r7��!�%����f�ץ4m�D��c�4�Rfԓ��Nb{.<�S����d��m�K�j;g!=��1�������3@:���f�,T`Ik��Q�;�vo%����x�i�EWc�a�9'. ��ފ�ݟ|jb�Q�H�1)�h�>4��`ʘ�*`zR�5�����f�܆��`ʘ�*a߳33�?�~���<��e�F6�G�q�D^j�?=�"�"���a�y�˃�����qf`n� ds)��+���u�q��=[&�q�v�`�cq�tdt�9�$�-�SX���׌YS�AasE�#�����bL	b��^0	eL˕0&̛�3V#�F���0,�� �T�,�SX��[����O�S�G3@:��z�L	b��^0$ʍ�ܳ�y,7��� ��L	b��^0	e�I<�V F0P�@`��;������?� �M�  ʚ����@�%^7[�'N2�-�hF�k5�N��Ӵda;;N��"���E�s�=SN	$�"�[����F���ݸF���.s�m�]=z[��m��tTNNM��N��	��n楁a�-PM=���3Nj�l9<�I)RQ�C�h��a�ĺ�3,Z|v�?�>����Q	�׆���srQ۵h�׍_��6�5g�Ɣ�*0��u�z���rf����s &5Ւn-Z��5b^�E�0-�� �T�-�S��%�?6�Aɉ�@���u�0fT��*0���ܐ�˻E�r�,��[2��Q�l�4{r�c$#N
G&�[�f�=U��zʘ�4\b0��{�&�T`[+��*`̳@�BH	8i'���S�'y���f��vKi�K����sJ�S����-��ݱ�'�[�s@=�f�[�g����X8���WQ�e��soup���F�%h��B;�w8wx�Q�l�eF��\����0fT��*0-�� �T��ܴ��"Q(8� S$�:���oW�YS �eLL�������#R�ӹex�%�0fT��*0>����(}$LrCȠ�md��i�E+�e힍�nܵ͞�x������d�%�<#��!�� _��@-�@�Қ�w4{r�c##N
G&�u�{�U���p9ˀ<����<��D�n#6�1n�=���ˏ�S������R���| Q!0�U��$�F!#$"�7��`k!S��E JEy��g����S���C��5�B��~a��R�z^{BH,�Z��𔿀=�"zi��4���~͡ ��\�dI�t|�p����`���#� N�I����_9�I"@f�� �|��M�����蝀B�A?y�
=�O���1"�"��G��H����W��27:��Ċ@ %l�ʒ*`�<N~{� �OR�)�:��U8� �� ����ш�Ej���z��b��-AT��{�o$��zwy$�vrT����8hz�h^��<���J�V��pV1\YFї���K���2��Q�-T�9^�A�O�Bra"��!I�\���ps����4�c�Vy�յ�nm�p2�A�'���u�M������X}�4s����"DPQ�BS$�<���v96 ��m=�*��������me�/u]��p��<����]�E7�q�8�v�3t�F��^^�y�J��q��"��y�Y���� $HT�U䊪�����NI?{�}s�̙76�͗w7y$�R��'�����?���������k�{��II���F�-��5�CNʽ>�[�ͷ7I�F��n&Q{u�Ϊ�Ç4�,ܚL��s0��I����y�g y��T��"��;i��,XcpN$�u�����~�dSx?k:U��cŔmz������ɀKr��Q�-T`I���$�Ō�NM ��^��-��׬�=�-51H�)Y -[����ʩI:�9� �O~�~_I���o��� �.�  [������읓Z��6-��Y�bq����J ]����mƂ6W],v�%���u��ʍ�n���D�,(�n�]g��.W�vl�rs�ru�f\f{�N���^9ܳku��+��\ԝH;cX�|g�����ɍ:�M�����]��a�ے8��s�Nᚸ��k��mOe��������z���svh4���#�  n�$<��s3t��rdˣl:�v���-��C��c����#�צ�r,2O�L��s �Ć��w��@:����^���U1H7�q��f���-ʘ�F�Q��Ǉ<��dq1�H���,�;�(���0YS��t6担�n�wv$����	j� ��0	nT����:�ncq'�u����4��4��h���$�'9+��Yӽ�1�zh�Y�se�4T��q'�9�ۉ?͘�?��51��!�޳@:ܻ�{��}UK��ɰ�<��a��]�j�ɳ.n�I=�N�=~��>�P�7&À��À??=�I%v{�@�6$	Ɨ�L�@����@��hwY�ܳ@����ܘ��1ɋqh��'C�#sx���JUs�%���c�xGC�n{��>_}�M�{$����>�I%~�j�w�9��L^��l��״�%�v9s	P<�b���gk��dFI��sp�[o8��rz����x�� ��J_���~^Xˊ��Q��ڼŻ�7��J���$�\�8����Uvz���K��f��ݾI����UKP�%B�H$R �� B�H�E"�T�B
�H��'��g�E7�����<�<X�Q����ӂ$�̒g I��n�"UW'��_��|��n`��(��n]�"U&��I6��p*��a6f]�j�e.�������5��.�ك�����q7W�ݎ���PlҾ���>Ͼ����=m��R���o���W�U�����k/6�7�流�Va/�� ����y�w�*Uv�&)��6��N_}��nY�ؕUۙ%�M��z��f ���4/ws�RI]��̒�޳��R'P"�x���� �  >'_�%��߳�N�3��]̺KL��1n��w�JRN������@�������$�<l�&�Ȓ�	��e��rE�q9�fhz���֛��U��sw���>��n$Ф^����?�������`�I|���,�h7V����m�}U����}��>��޳�Wd�i0�Ֆfj-a�{�� �Sx<n��U}T�d����%����~���v���n�K�[�U��_ ��p��$�T�'�/���S�W�U�����,���<޳�����M�}��'�/�������I?��{��~�?~  $�F  	5�We���5I���Ʋ�&U����G�L�)ۡv���vc�戛����e6݀�+�6�������`��鷧>��m�i�m����5�T�qP@֐��v��`Ꭳ�� eSY{uѬ�Y�{u�e����7�"����P�b�.��T;k�\��͉�I���t�7kzmJ���H�곩װ�\Lw��`⤍78[ي;	�ð�HnΝ2Ν:ӛm������\NУ�V�����>�5��͡�7
�_��ܳ@����~�I6�̲�F�ޙ�{����ޕUv9�_ ��p��%J������Q��5?4�M���@�e4���U۸�p�M�?_�;a��hY�f+����r�*��'�|p_����{�*�UUUɮ_%c,�(�Ն����;~y�D�*�V�S�����h�
����BR$�REً�(�kvŬ)N��ץ�$�#�����{���v:�X�Ɔ�"�? /�g�@��Z��ET�_���{�Dve�y��6K��$��{�Ψ�D
(T z@0&3ą�Z�P3���*PX���(r��oӒ�����U%v~�"��j�sV��/v�	&Àv��UWd�M�'��� �UfIam1�h}��q��	"��7�˂U+�O��H�L1\H���4/ws�i��UW�/����O�@��z���O$j%-�TlHntk��m��Ҩ���vv�t��{ASo�Sv^n]�\���w�'�w����.���J����Sx_�.ջhY�f+���y�g}�*U�}O��'�/��oϗEIU��cŔmj�ww5p��m=�h���UE"���	*
b
3��x�����{��s@���i�0x�/ss�URUv�Sx	��y�˂*��s#��{�Dve����f�z�x��p*�rO����p�Ox���Y+�.���s�@�H�(�������iT�.u+�G�6��ww�����}�n�wQ����� ��� y��U$��}~��~_3$�0�6�����Δ�J��o#��6�tJ�+�E�a��F�ޙ�{�� �Sx��q�I%�U*Y����}O���_�<[W���V^�^-��UU������$�����<N����	H����-R�`t@��<��y$��;b[����b��\�|���T����~�}����@�����psi,���d�6�\q�B�M���@�tP=+W,�ؕ*�\u��mj�ww5.9� �f���$����r�OI�f����b�v�78���IR�vH�.G9pߞtJ�U��)�i�ff�u��o#����q*�*��/�@>�y��&"9�G1"I�|��Y���ˀ���g 6ټ*T��UUg�O�. ��`�v�ss//p���;~y�}I$�ꤒY��|o�>��p���&��p�c	9�8H7	\@�EP�!U�TJE$��+M���c !p�P�CSR#��C�@���,�=��q�Y��bz�C�7�)��,,PsW�-�>C��t�U{矽�  �!�          p    8 m�              �+]/-��&��*�Z�`X�t�����l��ڶ!vm�U���fgy�C�8mk���pYƔ�r����N�S��n*Ǔ<�F�݆YM���Wk#sk���P�k;?=��c�7�l1Ⱥέz�j�<8	1,�Sq�PC���ޣ;�֠�5�T���ĝ�$�]T�7ceU���h؝muS�v��i^73[V6p�Rl<l!6�)��]c<�\� ҭS�ꪤy��k�j��	�T�jm�1�^�w���ncҡ0�	�t�<M)��`*��J˞�v�N�:y�%+:�jk���4+�.��uKδJ=P�Q�ݮ�����q����8�ɣ�5:.�"j�\gO5&����ݓ���=��8�' ��=wDl*����/|����Ck6��\\קۃ���Ѹ�6)�aT4-Z������t�+�%R��-�#\l��C��\܅w; F�]�3<Je�=�a�z���99�ck�{��j|�*����6�-�-@aĤ��,��gkŗ�-� U�� ��z]��$�@���0�[v�IӰ�3e�5�ԭҢ��\�B�7���9ZUU*�)Cu��� �wQ���Վ�rKӠv�v�T�l�%�V�ڷ<a�u�u&��)�Vⱡ�Dh�q��u���s]g��U�T�V �m��1����P1m�����6[�� fi˳�1K�:�)V4�q��i�/mb���	ǲ��6+�*[�% ��=`赚��:��n6�Pћ1z���@j�������Gi��@s̮��
qF����DV��$f$;�z���Ѥ�5Q�@�uR�Sq��+�*/+�}�o�z�Gio�:$�TN�N2͚6n����:;][�ݺv@�g[nx�^�tU�>��yQ�<b���V��T��U z�������.t(�y�󛻻�������n��  	t�v��l	�SX�ƹ�:�@K���.-r���&�D����)��8�U�m)k*V��N(Ƭq�v0�s�l��ȓ�F�G�p���p맷fznCݫ���ی���m�+�s�����P,��v�e���7\�l���],�Zۧ��ڶ��D9�\�L�Μ��$n�4v�����R-��#l�{6F�*�{���{����m��$\)0W0�����V��v2v�mx�ví��7rrZ-��W7���Ʊ��xna$Y$ ^��������)R��	rL�?/2���ޅe��o �|��%U_UUf}>��}}�pm�ҒWg�ȗ(զ���1^�G9p�y�ԗ�f}���}�ܸ�յ�mj�ww5pD�d�8I�o�I\�.�4�fj���F�7oss�l�*������������(5&	��9 �Ʋ��Sa�b��cxÁ�r�l;��ěV������I���HO ����o]���ϒ�����|o��W�U���w4�n��'{��suR~B��A#BAa-P`@]*�'�Ĺ=�<�~|�R�	�w+wo1��y{����pm��I]��.G��X��CH��[����)]���#���k8>�I%�,�~��@���PK�S�S@���)F��K�g ?y���f^���I�%�KN��ю�ZvmΛ`�v\]q�Hb�U��s������'��G"Nn���7���<��;ߪ��J�`}����X}j�YF�Y���Ӏv��R�����G9p��tT��OI�f��s	��G�}o�h����Y����UR��RW�^À�����f��^f�k47v��ꤾ�I*Y���ˀ�M���<�򊪩UfI�?y��}�������|@/�߳3?Wm~ [~S@�����Y"c��Qٶ�h�b��y콓\tmۖ��\L��<���tݟ������D/i�I�o�����8����m�Q*�����8	&�$n��i�n�p���D��b������Â�A�A�A�A���ӂ�A�A�A�A�>������ɽ��7%�\�˛w��A�A�A�A������lll~���pA�6(�����g �`�`�`�~��]���lll}�d�|�7iݳ�� �`�b�L����N>A����?�����A�A�A�A�w��A�66
��UX$b�MU����r?��~8 ��M�Կ�3I�&������lll~Ͼ�8 �?�"�����?��`�`�`�������� � � � ��y����lll{����˻mɖc�[�R����bo<�1m��nG9��$m��C����٦�:9
��{��������߾��� � � � ���xpA�666?}�}8(����>A����O��L��r�l��ɹ�x ����>D� ��������|�����g �`�`�`�~��]���Tlll{�������374�3t���lll~���pA�666?g�}�|�������}w��A�A�A�A������lllo��߰�ɔ��r�nK�8 � [���>A����߾��� � � � ���xpA�66"6?}�}8 ��4�L>	����3ws��A�A�A�A�w��A�666(D�������lll�������lll~Ͼ�8 �=g{�۽��������� �	��  ��}���N���n2�v�ڰ��/-�cW�dE^.b���UV�� #M����^��d�gtU�co)�#Z���&�ñ�kO7�nm�]�Ӻ{s fݜ�v4�b#Wgq�]R�U�<�[28R̽��x�dy���6�\Ƃ���!��v��{v�M�2E
=����3����1���P�)r�aգ�������5�W��L��u���9v�c�l�1�Eˮӳ]x��{u�~�ퟱ�7%�k�Ysn�A�666?����|�����w�N>A�����ﳈ��A�A�A�A�w��A�666>�}>f����م�ӂ�A�A�A�A�����ȏ��A��?�����A�A�A�A��]���lll~��8 ��6}K��L�d��ݜ|�������g �`�`�`�~��]���lll~��8 ���>�|����~>���.f�]����>A��F��߾��� � � � ���xpA�666?}�}8 � ���ﳂ�A�A�A�A��'�fi�����f����K��I9pR��U%�����_�}� ��� ~��1Ͳ,U��Z�ݦ�\�X2Q���m˄ײMι㞦���巙�o�(K���K�.�2��_�����p���I*���>�h��_<jcX)MF'�k�I���UJI*�	'��=�_ �����" ��?��>)��M7n�n�p�}{�7��*UWq��.I����.�ۻ����ox%*��M���Àv����]�����BQ2E�I�)�{�4
��@/uS@�ڴ
�T�ԉ&19�I�l�wb�(���'`�u���I�-�Y���Ć����,[��01��!�/����h�w)$��#{�4��7������� ~��_R��}�}��I�V׿g�ى�����ۄ_�	"��%���b╕�%Ki!	PR�Z@�Ab�`jj��2&D�>���yı,K�~۵9ı,O?�B�kf�neͼO"X�|��2'Ӽ�br%�bX�}��O"X�%�{��ڜ�bX!2'�s�Ȗ%�b_����]2���t�v�r%�bX��{���%�bX|�s߾۵<�bX�'�o�^'�,K�����r%�bX�����8���Њbl���k��nN�6퇘���6$�:Č�̎v�nwG!��a�~�bX�%���ND�,K����<�bX����C��L�bX�}��O"X�%�ߤ܇�6˶�.��ݩȖ%�bw��g�|�r&D�>�ߦ'"X�%���}���%�bX���ݩȟ�����lK��_�i�Hnm�]͜O"X�%��>��Ȗ%�bw��Ȗ?(���/�}�jr%�bX�}�>�O"X�%��d�/M�XL����ىȖ%�(�2'�}���Kı/�}�jr%�bX��y���%�`P ��e(9�����e+)8���/7I��m�8�D�,K��۵9ı,N����yı,N�{��,K��{�'�,K��s��n��E����q���rgX.1{��Dg�^��[�'l�n��w{}�r�*�=[TG��,K�������yı,N�{��,K��{����2%�b_��n��Kı?zw�᭛�]�e��8�D�,K�����>�DȖ'�}��Ȗ%�b_��n��Kı;���O�U�Cq6%����p˦R]ܷ.仦'"X�%��������%�bX���ݩȖ?2&D����yı,O�~�Ȗ%�bw��)p�&�70�34�yĳ�DϾ�n��Kı>��}8�D�,K�����Kı;��É�Kı?znC�6˶�.�.fݩȖ%�bw��gȖ%�a��~���%�bX�}��O"X�%�{��ڜ�bX�{�;�ߟ���� �	5�  K�a��}��dӻ�`��Vvm8���l��n;Y 1�ֺZ����.�z^�& ���w��^��笝ҧg��14�^P\d��c��9��.$-��+�\��'$P>��;,ɻ��R�ZH��앙��[f� 6�2{<��۞�c�ua��X�W$�XѧK��*K��R:ilgir򝢆���=���n�T*�b����ѳv]�E�qQ`1�E.�>}�.5��8�g�ݚD����̷����ı,O�����,K��{�'�,KĽ�v���2%�e)'C���e+)Aa-\[�X�������,K��{�'��#�2%�~��S�,K�����yı,N�{��?�ʙ���ܟd�ܙs6M6nm�8�D�,K���v�"X�%�����O"X�ș�߸br%�bX�}��O"X�%��p�e�m�wn�7v�ND�,�`dO��ϧȖ%�b};�ND�,K��|8�D�,�_�.�����S�,K������[.�6�fl�yı,N�{��,K��#��}��~�bX�%���ND�,K��;8�Oq����~�o�8�+-�
�e�ݎۣ���m��<����|��ʧ3K�H�ճ1�t�K�l˹.��Kı>��8�D�,K��۵9ı,N�����"X�'ӿp��Kı>�gm.}!&�70�34�yı,K��n��?�~^�hϒ�`��Y	 �Q�B$�"��0� ��F B*��F0�"� A`����x�	�Fd"F DBE�c�Y$���:�2��5�<��,M����O"X�%�����'"X�%����O"|�TȖ'�7!~�m�k�v3n��Kı>��}8�D�,K�����K�?���؟����O"X�%�����ND�,K�~����v���p��8�D�,K�����Kı;��É�Kı/{���Ȗ%��$ȟ}��N'�,K��>���mfif��i�Ȗ%�bw��Ȗ%�a�s�븞D�,K��Ӊ�Kı;=��ND�,K����n���.��WF���ue�ص��Ӱ2u�x^�hRl���=��u��$�[g�1]���%�bX��븜�bX�'{�vq<�bX�'g�ف���&D�,O���'�,K��O�ᙹm�wn�76�'"X�%�����O"X�%����br%�bX��{���%�bX������O�C�q6%��O��/��]�m�,����%�bX�������bX�'{��q<�c �
 � �_y��N/�0���$"0��Hb�B�<��0�v��x�B���54	�	٢l98x'�!�p��q08�<?,p-8���hx��K"d$��6"�"�E���
@�)!�A�L�%`.�0b~pN3���5��N �D�cH�!e�xD�VH�$g�t1��(���*h�/�� @C|���(�=N���B��� � x��TA��S~P�Dȗ�g�q9ı,O���N'�,KĽ��i��m%۶eܗ6br%�g�"}��~8�D�,K��}w�,K��{��'�,K���{19ı,N�g�ܳ��l���3N'�,KĽ�v�'"X�%����ϧ�Kı>�ߦ'"X�%����O"X�%����9��%�w.��\�#��ʹ�3m��zQ!\��q�㴁�i{A[W�u��`q[���~����%���s���%�bX����'"X�%����埢dKĿ}�]��Kı=�d�|�7i͗	����Kı;=�ND�,K��|8�D�,K��۸��bX�'{�vq<�bX�'a���7[I3L����'"X�%����O"X�%�{���NEYPXR��Կ�VR�����,��,K���yܗ�s3d�&��Ӊ�Kı/{ݻS�,K��{��'�,K����19İ:#�dF+"^��O"X�%��s�fn[rn���ݻS�,K��{��'�,K����19ı,N����yı,K��n��KǍ���������Wk�ջTg;�t���jcvㆮ�u
�6��Y�Y-�Ω:��.�6�Y����ı,O�~�Ȗ%�bw��Ȗ%�b^��v�"X�%�����O"X�%�{�vf[�e%۶eܗt��Kı;��É�Kı/{ݻS�,K��{��'�,K����19ı,Or~��w!�M˛��3N'�,KĽ�v�ND�,K��;8�D�,K�����Kı;��É�Kı?{f��-�m2]�]ͻS�,K>H�����%�bX�N���,K��{�'�,KĽ�v�ND�,K�~����v����76q<�bX�'g��Ȗ%�a�G�����ı,K��mڜ�bX�'{�vq<�bX�'{w� �!� 4ڀ 
�H-���*68Ć�@�bW7k��Wv(=���8@{��hʑ�RW-r�Usl;�iP�W�9�_+�LM"��TѺ-��ʏ��cJ����pd�D��\QD�����Rq��tٮ��k84n��O*�k�e#a#�5�0p�ͧ<�፹FG�̝�Ϟ';��W�VL��n�����خ�P��-���w���n���	�����6z��6'�63d3AW2�/�G�����^�=,�;@���X�%���}���%�bX���ݩȖ%�bw��gȖ%�bv{���bX�'�;��i�.l�d�ۺq<�bX�%�{�jr%�bX��y���%�bX����'"X�%����O"��2%�ޟg$�ܶ�wI\ٻ�jr%�bX�}�>�O"X�%����br%�����blO����'�,KĿ���v�"X�%�����_l��ۙff�'�,K���{19ı,N����yı,K��n��K��&D���q<�bX�%��l̷4�K�l˹.l��Kı;��É�Kİ���}�jyı,O���N'�,K���{19ı,N�{'wl�p$A\��څ��콌��:���:����Q���u{Xz��$k��Ȗ%�b^��v�"X�%�����O"X�%����`|<��,K��É�Kı=�϶[v�d����v�"X�%�����O!@�ՀV"�Eh|�G"y��}��ND�,K��}���%�bX���ݩȖ%�b~��vu��aݸM��yı,N�w��,K��{�'�,~Ea�2%���ND�,K���'�,K��2v���,�4ɻ��19Ĳ�(2$�m. T�&�ڤ
�R���¤	4��Q
P}��+)YJ�N)��L�wI�Mͻ�Ȗ%�b^��v�"X�%����q<�bX�'g�ىȖ%�bw��Ȗ%�b�s�Y+��h�]<�tA[U�K��=cxÁ�r�l;��	���E��{���o�/Vƛj��ݻS�Kı?�����yı,N�w��,K��{��$�"X�%���ND�,K��~��r]�m�fn�<�bX�'g�ىȖ%�bw��Ȗ%�b^��v�"X�%����q<��TȖ%����4�K�l˹.l��Kı>��8�D�,K��۵9ǀB"H�`)�11��������7���yı,Ogw�Ȗ%�bzg�����e�.n\�8�D�,K��۵9ı,N����yı,N�w��,K�fD���q<�bX�'��d�m�v�e���ͻS�,K��{��'�,K��#��>��D�,K��É�Kı/{ݻS�,K�����2D��A�$g����WK%N$�j��8��r��k��q����<GEzg'Naw6q<�bX�'g�ىȖ%�bw��Ȗ%�b^��v���<��,K��Ӊ�Kı>�O�~7Yd��M��ىȖ%�bw���1șĿ}�ݩȖ%�b}���q<�bX�'g�ىȖ%�b{Ӽ��-˺L2nm�8�D�,K��۵9ı,N����yı,N�w��,K��{�'�,K��ӹ�3�,��Wvn�ڜ�bX�'{�vq<�bX�'g�ىȖ%�bw��Ȗ%����"s�wn��Kı?zw���\��n\�fl�yı,N�w��,K�����~8��X�%�~��S�,K��{��'�,K����m���`��ڶ�!���D�]��F:6��P<-L(��Kc�nO���wʭ��۶eܗ6byı,O���'�,KĽ�v�ND�,K��;8�,�"X�'ӻ���Kı;��{>�n�\˸iw4�yı,K��n��>TC��bX������O"X�%��>��Ȗ%�bw��ȟ����=��?8����8���{���{��'���?�Ȗ%�bv{����bX�'{��q<�bX�%�{�jr%�bX����zˮ�n�]͜O"X�|�2'Ӽ�br%�bX�}��O"X�%�{��ڜ�bX��b~��O"X�%���Կ��,�tɹ��19ı,N����yı,?�F9��mڞD�,K��Ӊ�Kı;=��ND�,K�������C��R"$�{��������$mp  6�N֩��QM�;���t4�ɢ5ͱ�٣m�� g.��qm(�p�j2�^T�cr��8����psX��k��,M��w*q8���y�vƗ��U���z`�!�{�8[����䣇vW��{��LLL�/g����?^�ս>�pW:9�؜.�H�>*�-��7�kc�:Gi�uh���9�3�b(��ny�-ٗvۓ.���E��N75��<�l�4%cM�gV;vz�o����Y��s7d�&�����ı,K���S�,K��{��'�,K����19ı,N����yı,O};��p�%��%wf�ݩȖ%�bw��g�|1ș��w���bX�'�}��Ȗ%�b^��v�"|�TȖ'�N�I|5�sK�2�͜O"X�%����19ı,N����yı,Os��ڜ�bX�'{�vq<�b�oq���8�n���������ş+"}��~8�D�,K��ۻS�,K��{��'�,K� �E��}����Kı>��O��ɲ�2�]�8�D�,K��wv�"X�%�����O"X�%���xbr%�bX��{���%�bX=�{m�ܶe�-��k���d���1��c��\tu�NG�v�cc��k������*�s��Z�w�{��,O���N'�,K����19ı,N���� ��}��,K����ڜ�bX�'s���̺�ݗ����Kı;=�NC��&!�,K;��q<�bX�'����ND�,K��;8�D�Qr�D�>�O�~7[I�L����'"X�%���}���%�bX��{��9��!�2'�}ϧȖ%�b};�ND�,K޽��m���i�wn���%�g� 2'w�v�"X�%���s���%�bX����'"X���]��������%�bX�|g&\6�[�es6����Kı;���Kİ�T�ӿxbyı,O���'�,K��;�ݩȖ%�b_߻!��ɻ��a�fۡ�{S����F$��<�ײM뎞����
��@	Nq���fiv�Y����ı,O�~�Ȗ%�bw��Ȗ%�b{�����Kı;���Kı/}�v�ݛ��v̻��bX�'{��q<��1ș��}����Kı>��}8�D�,K�����O���,N�����$�K�w.�O"X�%����ݩȖ%�bw��gȖ?�{@H�H+�p}�HX�D�y�ND�,K��}���%�bX��.��336�d��ff���K��H�����%�bX�N���,K��{�'�,K��;�ݩȖ%�b~��e�m�d36\.��'�,K����19ı,>T��}���%�bX�Ͼ�ڜ�bX�'{�vq<�bX�'s����W[m�[uϳv\�Ⱥ�;.��
M��^��m_���u������m��*yı,O���'�,K��w��S�,K��{��'�,K����9ı,Oz���c�e�0ɻ�t�yı,N�{��9�O�J�M�bs�q<�bX�'��
��bX�'{��q<���2%��O��.I2���3n��ND�,K��Ӊ�Kı?v��ND�����؟����O"X�%����ۻS�,K����Y|5�3K�2�͜O"X�|�"{��§"X�%���}���%�bX���wjr%�`{��V,�\�-v%���Kı/}�v�ݛ���.]�wJ��bX�'{��q<�bX��?������?D�,K����Ӊ�Kı?v��ND�,K����]�˻��a���)k\#l�Ds{M��筰�0�'7=0�2���ۓe.e�4��q<�bX�'s��ڜ�bX�'{�vq<�bX�'�����&D�,O���'�,K���qq�eXqZ�Q��{��7��;���>c�2%����9ı,O���'�,K��w��S�?�C*dK���_�.�!se��l�yı,O~�p�Ȗ%�bw��Ȗ?��2&D�>�wjr%�bX�}�>�O"X�%���aܛ��˦M���ND�,K�{�'�,K��w��S�,K�����K���߯�9ı,N������w2n��8�D�,K����'"X�%�����O"X�%����*r%�bX��{���%�bX�_<A�� X����T�� �:	D�$!�8$'���]�	������'��w��,`p'>�q)�,XX�	a8v�DT��!(A"R��RBD#	�B-"�@�@��}���             �   ��              9ųY]l�X�ݥ�0�9@"����UMt�yH,�@��6��8���֝�ka�y�Φ�W�EYE8��pl���Aga�����MԹ�Q�j��H+)�gk��C�N��[�1��G��f��M�oSU[W��%�����j{\�X�x.y��`��mqvvjU��ca"`h����O+P *��uW@[j���^���<ݍ��h�r�ʀ�,&ѱ��6��*pl�U�[v�	����Q�y��m�= B�S�
SQ�N� U+���z�:�Oэ:�DI�m���b� �]qG5!=P�t�9�Qj���4�h�@v��A��]Z��c]���,�WKa�w�=��7^J��)��5zi2Z69UT,R�'1kl���h۲k�9坃�F�k�]\�]q�Os@�H"���o:v��A��������V^�	�*wn��Ԓ�%qY�����D�@L{o	����@�g;)ι�9��v��i��%D$:���5��K�c�`
�ڮ�Z� ����$��C��SVT�n@q#m�K͵�$�iV�62�+;�
�&�g&cpҋU�)*�+��a�է�����8�g�ս�tN�`Cp>�j��F�y2s���5��;lc��j�#y���[�/\�\/m�����h	sl8�y1�\�q�mk� �����;6�E	+�=bx�n�Z.���^�۰6w9������t�Ѽ��%0㴻9E)�e�pUc��#v��`r�z읞y[��ק�iH��vN���л5J�qt��<l���E�nf�P�q��E�F���8�Lv�2@m�{6!���������Ae���itnS]=�nͰ*�i�2f�Da���S��-��u�-�j����� -�<�̲\$�ʡ�D�����@�4#�z�>�#�� ��CDJE=;ǀ��G�A�v{�@ h&�� *����Y�uۇJ��(^���x�qq����$�����\p�S�9�[�E��=��n'�Guv�X��S�|Ak�VI���-�M�0$�6�����y�uu���D\��s��k��ŗ�X��.j�82뭕�Ki���-�v^A��g!��sq��b�[���2W]FҚ;%�M�s2雳i����� /�;�jf�<��l �`�n�aq�l��{��VG��Қ���q7W�w�}�G��Js6���~�bX�'��Ӊ�Kı?v��ND�,K��|8���؛ı?��?�q9ı,Oz}���L�.�2˛x�D�,K�oxT�Kı;��É�Kı;����r%�bX������O��M�ؖ%�����7$��v�[�T�Kı?����8�D�,K��ww�,K��w��O"X�%��oxT�Kı=����mɶ˓7.f�O"X�|02'w�v�"X�%����׉�Kı;��
��bXL���}��yı�{��#��ZW�6��{���{��'{���yı,N�{§"X�%����O"X�%��w��S�,K=�{�����;�-J��k�R^�L�Z�k!�!�Sv�<�7h3k����v�l�[�x�D�,K���Ȗ%�bw��Ȗ%�b{�����TY�L�bX�}�}x�D�,K����n�I��&�niS�,K��{�'��#W���G�2%����ݩȖ%�b~�~��<�bX�'gw��,K���y{f;f]���wN'�,K�������Kı;��oȖ?$2&D�}�LND�,K��Ï~����{���?}�~���务9ı,N�{���%�bX����ND�,K��|8�D�,�D�~�wjr%�bX��;�o��34�p�.m�yı,N��f'"X�%��~��O�,K��>�wjr%�bX������Kı/��m.6f�3[�0��YA#d;6=�v���vys�+�H�3���]u;�R�����{��7�����yı,O����ND�,K����?��o�6%�bO�����bX�'�;~��˗m�fn\�8�D�,K�w;��� �r&D�>�~��<�bX�'���br%�bX��{���'�2%�ޗoƗ7w..lٛ����bX�'�o�^'�,K����br%���=S��,ND���O"X�%���ww�,K������ˮ�\�r˻x�D�,�@��>�s�Ȗ%�bw���yı,O����'"X��ȝ��}x�D�,K����7[I��&��ىȖ%�b{��É�Kİ�U���}���Kı;����yı,N��f'"X�%���훳sl����e7Lb��#հQ�-��6T�n���0��Ykuv�m�1�2�d�ۺq<�bX�'��ww�,K�����'�,K����`|�<��,K�}��Ȗ%�w�����쮎�Q>Xj}�oq���X��{����؛�����19ı,O�����yı,O����'"X�%�秽o�5̹�m�,����Kı;;����bX�'}�|8�D��?��bw?��w�,K���~��O"X�%�{�[t�7$����]ݘ��bY��2'�����Kı=ϳ��ND�,K�ｼO"X�NG�蘰(@�T@�(�.�N��;19ı,O����w,ݲ���L�Ӊ�Kı?gs����bX�'�ｼO"X�%������Kı=���q<�bX�'����ݘLu�fZ�� ��:�v���piL���=��|F��j�!�=�_��2�K�0ow�,K����׉�Kı;;����bX�'���'�,K������r%�bX�����뤗6ܒ��'�,K����br$r&D�;�~��yı,Os��w�,K����oȖ%�bv;N���&i�w6��ND�,K���'�,K������r%��C"dN����<�bX�'���br%�bX���/nXm�w2n��8�D�,K�w;��Ȗ%�b{�����Kı;;����bXȝ��~8�D�,Kޟg%̻I����3nn�'"X�%��}�gȖ%�a�*����byı,N�߼8�D�,K�w;��Ȗ%�bAz{��@ ���  6���f�M%Iga:k�n�IV�ut䍔7\F✾��&^�������;K�*vү 0�+�b���緵�;������ҫ�&�^U��s�f���0���:�Y��;�X��T�7n)���������	�;6ܗ3ÜC��Z�\�;��O�5���C��n(獬t��Lq;�1���CS~��w������%v��uڣq�G0�>���^�q�jKr-T����6��jn/�*���o׻��bX�'�﹉Ȗ%�bw�{���%�bX���������lK����N'�,KĿ�]4��.仹�sq9ı,N��|8�D�,K�w;��Ȗ%�bw�y���%�bX���19�Tʙ���g�Lܳv��n�̹�Ȗ%�b{�g۸��bX�'}�{x�D��ű;;ڛ���xqI�?~,���d�K�ndM�I�@�'��~�O"X�%����T�Kı;����yı,O����ND�,K��{/K.�I���.m�yı,N���9ı,> ������%�bX���n�ND�,K�Ϋg��G�G�G��WH�!!b�u��Vm658�m=�]�C�B�*���]�f딙�eܛ�S�,K����É�Kı?g{��9ı,N����>��dK����*r%�bX�|���M0�7&�O"X�%��;����5���T�["X������Kı;��ʜ�bX�'w�O"*�ø�����r\˴�n��s6���r%�bX��o���yı,N��eND�,K���O"X�%��;����Kı<��rn�334ݺR����%�g� ���؟����S�,K�����É�Kı?gs�S�,K����'�,Kľ����Mܓs-���ݕ9ı,N���q<�bX�'��w*r%�bX��{���%�bX��w��"X�%��,��E���L	�;l997f�k�����ɱ�e���G+��͢��;Sf\Ӊ�Kı?g{��,K����'�,K��۽�9ı,O��|8�D�,K�K�����ۆ˛6fnD�Kı=�{���ȠG"dK����Ȗ%�b{��xq<�bX�'��w"r%�bX��ǲ���t�%ݼO"X�%��{*r%�bX����q<�c�CȒ(��C�E �����,N�>܉Ȗ%�b~��}x�D�,K�d��3u�L�2�M͕9ı,O��|8�D�,K�w��9ı,O}���<�bX ȝ��ҧ"X�%���ܿd�i�nɦn���%�bX���܉Ȗ%�b{�����Kı=��eND�,K���O"X�%����~ښ�(���7nג�!fv��L��n7�8�*�xz��quh���J,w6��ND�,K��{x�D�,/���-x��m��-�Z���bZ�sw��%���^0&�y�gZ���+&H�P��9��w4Vנ^v�������pN%H�i��9[^��v������?�1���"���sÒOޞ�qLr8�A8A��k�hg������������z��F�Nb"W ��Mĳ��cumzK�M��g�7#���\�r7�	�SS�R!�R-�]�������k�h��YY'�sK�R���`M��׭���X�ɏx���L�=W��=��`OZ�%��k7�V�ݩj�˖���[�	�^0$����ٟ�c���n}�3dSr)�	Šw���=��p�����w�U*T�UJ�{���{����� @i�  ]/5�f_Y6$m��G�gX�����W97��7��w�����ɮzF���:��U*��M�IӲtݸ��\G�Ò0�u��mCB��r����݋2b3\�V��zT�g*�D�X�`)��ưk�����8�$�u�C�tL��A��"d�p�.ݫ���Z�]��DcNd�=xl�"E=����wo{����Tp:�ܼ�61diy�;%���m�P"4g�Dik�v�]=�-f{v�.弳�-���e��[�	�w4�y��ؠ��m���������2K����y��=��Vn��b7�����[�	-x��W�+k�9vp�$����iH��w4	%x���y�}��{8����n��;�q�c�^0=��`_u��������$ƔɊHdJ ��� ���・D-�X�vvV��Hݹ�ڇ�'\�78\$����ηXZ��n��e�4�,R(�G�@�v����$P� ?���p䓾�w4U��.Z���܄�bĜZ����`{l�����i(� H�DQ&���n��^���Z���y��</�'�����?[���I*od�����?7˃~{������8�8u�͵�7*��Glx[�X��a��zⱧf�lLa�u�:����}��0�'9�|�����۹�^�s�?x��s8~L���kB�v�/v�~o�|�����z��?cw�{�Zxn��3Ve�����p���ԕe$������_P�$H�Hj�ኦ.!��0��k��g|��~
@�Hd���$df�ʒ��P��P�	e��Qd!aY.����]
C@���:	<a��"FQ�Y�N$ӀÄ�D�C�
A�)�,����-Юd�f$��$�
Jqh0D?]#3�L$5&��H��7?pH~D�V�7ȑ! �����]�z��Q�螥���;���/����W� ��1w��?yy$��{ÒN�{v�ZՋ/KXn��>_,{��8���Z{n�z����ti�X2I&���np����O��rr�?[�� �x2� ���d#H��q��`��xy�׌:����9�w}�߾�q�R.�,�Ƥ^{�4��hz�Z�j���!0mD�jL�/[���1]���_I|��|���xƱ&ț��3@��j�/;V��w4��h�@�j5ȓ��E�{]��O߽�I=����=R$`���`��J8&Os�^I=����ۿ�~Դ�Ե��J�%�{���ڴW�R�$Ci�A�23���7d�Y.s�p��:�����^���ۜ���^v<0sQ�L�;���<�ڴk�h��s@��Į5��(<dd�4=u���w�~��ˀ���ҩRJ��Rp�ȆI$��M8�����=����n��ՠy�k1l"nA��R_���.�o����	J�6K�K���EQ4��4�w4=v������ϗ�I�!%�z��%������m� 	 �\  �m�n���$Ӗ��풕�4��\��ƱXKusk��įfU����Wz�7 k��獭�b�諦�f�sOQ���h3�m[�!�[�͘���r�Km�i�	�ێ��3ՕA���.��f��B闞�^n\���vpuۣ��a���㜬'�WQ������%��B��U2Nu�F�N�w���j~*MT���+\#v�d!���v�c=Mq	m&'c�)���Ľ�.�����?��w�~x���y�/����-���j'�'�@��V��J�%�{���d6���?j�2�v�߼�p�|���]��I|���{q���O�1�������]�@��V��w4��J�Y֣���K{���[�zW�	-���*$jLj<Hjd�18�}!t�k�Uun��y�����䎈�����sY������v��z�h��}��g�=���@���3�$��(�"�=��xqd!�JH �i����1*
0L�5��g�ٚ��N�X�n�		N9�$Cj'���;���<�ڴk�h��s@�G�"dI�&�i�Д�U��_�_���.�o��q���O"N
)��v�����������ՠw�C6HFȇEד��v9�P��k����>ض�ۙ�Mv�n�f�7&��0J~��H���@�޻�u����V��v�ی啒~9��$��%�{���[�I^0%�bW�Ɣ22I���Z�ڴ ��tQ����I;�{Ð;��i<��r~q4��=�ՠ{�^0$�������B�\�R���o���>\I7'����/���ՠu�b�c��X䟌i$(ų���rthq�n�f.��w�ɹ��4Yf�s:՜�kLmD�ds<߾��<�j�=�ՠ{m��;=yq�,p��mG3@�v���Z����������Ra��D�	��"�;���@�۹�w[��w;V����	L���iH�m��y�\����W�$��J%�r����P"�f'C<�f���y񓴯�'����C@�빠w;V��v���g))4�M5n���a�Ÿ1�m��z�+��z��%��m��vfR^hV����Ɣ�&x��v��e4���y��I��ۋ@�x����p��.���UE�5 d`��� ���@�ޙ ��ܴ9��@;���Bcj'I�@�W�	:�`_u�������RX�8�bRf���Z�ڴm�`Y+�����������I$�I�kX  .�,<�q&Cny��)"8f�](Wmm�M%�='�<�]�GZ�^&Nr���f�3�Sr�KJ>����9�!N�2�l�\���)ũ�N��;8���uj�<��;��i6
�e+j�؞1n�2<n�Vn���\�+gZє�`�9�k�ۦL���b����r�˝[^\ݵ���@g��3s�:+�)�����������[�a
�5����Q�ص�]s[��C<�nS�����CtH鄂Q��A88�^��ՠ{l��{����Z.�J���a�H��5��UJ�'[��_�f�?��ba?�$r����w;V�}v��e4X+��cJ�W�T���/���/��޳�~��{�[�'�܄��M���hڨ��W�	:�`{�]�v���I��cv˂]P|�uF�c���T0[�6	�I�խ�+gc+J_���������`I����� ���`��3fne���O}��9�*�����μ�>�.�=j�g�.^[��Q��Ƥ��ڴ+�i�g��Ɓm�s@��&	F�y��h^�X�Q�$�u���2n�ƬF�Y�jZ���u�$��n�<�ՠ}��������#�H��K��؜�ѳ�E��:�D�������m�m�'!&�)�A&)�x����v���Z��Z_�
�y�x�L�=:�`}z�`zu���W�	��O"1�	?8�qhWj�=�jӿfV%(�J��n��Q�J�bBFl�ˀ�y%���˵�m�f��ͽ��o�UU+��/�m�\�e�@�V�wF70��88��Z��`zu��������u�oP�j���W`�����pY�Mٞ�vƳA�^r+��z<��
��s$�n'J9+��������ӭ���`}2,��Q<�yr-��[��Ď�ۜ����R�����34Enj�5-`K�����W�N�X^�X��I��~I�D�Zw]��v��y��o$�G��,D�
ĔQX�:(D�{�;y$������ٗ.�vp�䱁�������[�%��;��A�0M�S�$�	$M���	�;^���An�u���BM��=R��{�k����T`Y+��ڴ{-if�(��#��R-��F��`}:�`_u��$%3��j�4��7t���p���J��{$Z[>4���ư�%26�ԙ���{%��%���gUq���4�/��j'�O#�E�_]���]l�5[o}��ym���w9m��T??=w�}�j0�"�pP����)!O�����|0���D�Nwx�7�Iׁ����&��&��6�b�Hċ44O�p<�Z��<��a�&i8L1�I�p�VI$Q��OY ��}$��������p'O@����=�ā2'���$-�C�?ozL�? �B�o;����                 d��              $�N��=-�U��v��('b-q�	�B�R #��ᵽsl��Ꝕ	Ű�(\t誫E;���4�g�N�i�d��٫�j,�+硕{����	����\[��-�2��Y�<qm��T������b�:�s-�r���{,kY䍬����s�!����veixf��E�U�Tll��n����m@���:2Z�I]���r�Kn{Z��ڦ�VE��4�$�-[%� V�� pI�Q�S��r�h���J�@����`�V��H� �m+(l����t])(X�-H*܀�#��j��b�	궎wVR��8A���[2�Tnc+��yv��66w[�D$ň���F�4ZM�H��Xç�kn�`��T`6��;X3��z�X9�8��d
v�k\�ΰ����ۅ�.���f힊+M������6�Jx��*$�ڑ��ƗY�^:���m��<W9tK3F��2�6����������6Hnqd©�ۘB\8��U����[��[T۳���� @��F�n	 Qn�[d�uj�B�U �p����5�J*vq=�Svi˓���U��e�8(�ٲ��ݪ�(��v���v'EV�鬠Vs�D���(v���+�]�J���8]����Bj�l㤺@��������n�����<�����J����mu�ݶCu��kq��=�%@
��K���k@]�����\�^yΎ6#�&�
ڃ��z�n�wnÉ�Lv5�n���V�ì�T=�تU�����Q��q1$����`����ѐ����q�O.-[Fv�X6�M&捓���gH�N�,��v���<�K\�.ʥ�[l�;	q�Ll�x��ZS���J��RNP�)�
������j(�S���P4�P{Ǫ�&~@?"��_�w��wwt $�P  '^B] c[HjT܀F�N�4&c@W{#e�T�`<8�8��%������4�Ź�J��AΛ�OKѫe�& r�b�ە3�K�c��R�sk���]�3q��ʬQˎ���:9k(�!3��^�k.�5�n��\��7U�ף׮���m�)�B^�C�&\{u�=x�v	����g��w�����T���As,�غ	�[�n���ϧ��8z3r=��
��We�:�5��������������}[m�;�ϕ��o���_<��㝉��O�	1H��jI+�|�<I%���$��Z��$�ٸjI+]c�&�ǌ�rg�$��lz�J�-^x�����jI/����Ē���xL�G'�nG�$����%���RI^��y�I.vǩ$�쵥�B(��#��H��$�ٸjI/�ffe��s�RIW���I/,�y�A�������m�W ^��uz�[�0�iy�;%�-���Dh�K�꒸�h���VQ�Y�l��$��y��I.vǩ$���ʪ��.�ɼ������^\��^�6�wO<���w����URݷ7m^x�]l�5$�w_3�K��1X%����=I%喯<I.�n�K����$���5$�>�H��!���&)�$�[��K����$s�MI%喯<I.L�p��`�J@Ԓ]�|�<I/�ff+>�OI{����%�������,������vz ��S�q�wX	�-������Hݹ�ڇË��c�H�&y�I�SRIye��K���~����V߼�<I+C�'�H���m�5$��Z��$���Ԓ]�|�<I#��jI/{-ig��72H���[�Iu�I�m���|<�ο��@��A�mW�=I%���$Z]Na�pq�I������?cv߽�<I%_�G�$����%���RIv{0���11Lq	I�x�K���I/,�y�Iu�pԒ]�|�<I%_T�I,��nDB!�s+/-��F�z�7/]=��^$�<t�Z���7�qG$z�K�-^x�]l�5$�w_3�Is�=I%ϳ�/��a����m��m����*f[���<������Z���W�$�6rC�O�	0R%&�K����$������W�$�[7I%���V8�n,x��&y�I.vǩ+|����-���xN[|�Q�����[���x�]�wZO"$����ۑ�I+�y�Iu�pԒW���x�K���J����'~�	�cD���m��[ч ,��xy��Luz狴tw�����ԇV�n�ӍȽ�$��M�RI^��y�I.vǩ$����$Z]Na���l�a�$�u�<�$�;cԒW�j�Ē�f�ʹ��`��`�,jb�JL�ĒU��z�K�-^x�]l�5$�w_3�K�ǅbZ��(�Dܑ�I/,�y�Iu�pԒ]�|�<I}�?7g�G�$��R>�L�����^x�]l�5$�w_3�Is�=����~�����o�����  k� �Jv�oIf�bg"����J���.���94bGc���[J:#[nz
'�����@1�G3vn�n8v�E���7&5��A��Qv���&�ίV�s�q�RY��U��H)�.ݢ�;���VWd�:�C����<sRr&ztmt�����u�N��ˠ�]9�O[��q{%��u�	՝��(�]�p��{��{5�qP��ak��f��}ulv����s��lq�glg���={s�]B�3v�����)0�$��}|�<I%���$��Z��$�ٸjI.�
��Ēk&21ɞx�K���I/,�y�Iu�pԒ]�|������wr������ �*��
��	{����%���RIwu�<�$�;cԒ^�Z��!nd���ȼ�$�ٸj[�J�OZ�^�Xҳ�y~�ݫV��c�+�=j`}:]`z˹�}�3����I$��M�(8�u6Xz�.�Ż����%Ң[F�e3[]�K����,��ﾚ�����s@��h�v�k�b�M�4=�{y� �Z��A��U���3���$�����{������.h� ���xԵ��+��>\JI]��o ��_��z�ƍAv%����0>��`֦�K�Yw4q�aX���LdMI���4	�X��`}ex���D�{tC���Ƭ-�����6�u��Ⴡ�#�/f�9��t�+�kC.��I��ߟ��=ex����OZ�e���Wrė��-`z����� ��0'���:������S�L�<�w9$���w��ؓ��['� �� �T�*\���c��zGˀk�xƷU���բ0Ա�zZ��.�=-x�����<��,�	�)�7$�;��X��`}ex�=-LYCH]�4R�s���ٶ�ȑm�-���bhx�ۙ뇭�Wk(E2A5�(�S���Xԋ@����>��`���K�l&�բ���R]�Y^?f�Ky=���� ��XsɌ��3@/[�.�=-x�����[s{D�\�䷻�`Ot����x����d 
(������wӽ�Nl۹�j\.�䵁�Z���� ��L	�h�(5&4�F���$��	l�g)�b��m����?������p=%FgZ��zc�Ě�<߯ۚ���}W��;��s@��E�50Ƣ!��4�m�	�X��`}ex��ΚTv�GvjՋ{�LzT�����+���4U�J���s9&�˾�y�����=j`Ҧ�v��`n�a�n�������OJ����w�O��_���  -��V  �ג���^56��[y#��ܚ���t���<ⵐ�w {�Am6dUW��Z�vNtݷ$7$���J��]ug�ԡ;��uBPP�r�s]<�y��X6���-��z�uE�"�\��j8�	e6xɍ<��b�h�M&��e��_T�v��LI�5��ŝv[Y�ѫȇS��M�S�mvr�-��Iow� _@�(97g,ݛ�f���@yn��]͞	:yS#Nb<�`cY@�2��B��0�E�b�CY1�5&hﾚ��{�~~|��T��?G9p�ۊ�Wj]ܗ䷻�`IS�W���{l߿~�ď�}�K6F�9PjH�����I^0	�S �ژ����~[��!f��cI^0	�S ��4o]��
Ȇ��D��=j`[S�W�	%x���ʳ��V�q�ʹV��&�lvK���`��p�����&�F+�GP\�i�]KS���W�	%x�'�L	�&�%�]�[�d����}�(qD��	H3��b��$�����m{�fbG,�_(��%����0-�����}mL?>\���-����Z��3upJ�J��M��M�??>\��ˀ���j�gj]��[��0����+����~ox	J�{ӥޙ{��ի4/r���d�m�櫩7^��XJ�I:�`ѰLjٛ�iB(�s��5$�����wu���٠[f�֗�O�<c�ĎKJ�OZ�������x|*��0Ƣ %&h{l��g�� �x��((0�D�1**b�Dj�d�0������$���wA�t��B2���Ā@"JJ"���1�N�]�0%�sr��@�byS��!0��F2� p�8����-����%�ZJ�=׌|<��v������9��?'�)����?���~Pz/�k㟿f}��~_�����K���o~Ļ�L�������^0	�Slɻn��n��_��LY^0,�� �T�/�L�Z-.KR����@��ɳ��\$���V�k��B�ҵr��H(� �%&
AI���� �ةW�����	�qZ��Y����*`֦��`^빠we�s"��	�Dۓ@/����J�OZ��on�j��@�	ojI��+���`֦	0�QO��N*,@��}��I���~���!ɚw]��ߕﾞ {��M��s@���$�0�$;cb��3��<a�1�ݸ�l�ye䲙q=�gqt(%"L�cQ�4��h�٠z��$��K���r��.Ļ�w�?�{ҕ*����\nr�~oz%J��vӹ�/kv�v�7w��s��y��U��&����~���l۽�R�R�KJ�OZ�����빠[��ǑY1��L����/�LY^0,�����3��̾����{������~~�� 	$�  m��v�Cp2ۡ :6B��F��Y�֎�j, �v6���K�� p."�����m<���Wx����#�ܖ�u��mr�;_���|��b�6k:���L�D�ts۶w6wFG�����g��ӴK*ۃk'B�֢غ�C�7T���K�6W^e��]j�Cɣ�tzã0:�{/cS�E����߿{����-vnf��;�-�ح���3�v����n�t�Eр�1�n��)���M�= �ﾚ�����s@;�f��u*4q�<�#$MI4l�J�OZ������su�-���NKJ�OZ���@����/��+s5"M9�ؕ�����o������p����'�G�7$�/�ՠ{z�h��h{l�<�Ԕ��2%��s�=������7�2m�(�E��k�й��ޭtI���n�Գ{R���J�O[������a=�_�M�恪��Q{�{��~�����I%�����f�׮�n2�WDd�F93@%�0�SY^0,��L��o,Z�rĿ%�y&}j`K+���h^�@�;-i��##C�h��d���}j`@�[+0�:��O7't3Nș��m�Z'e�]���;jn������5�̱�d����_Z���`_�N��X�QA4�h{l߳?~�H>���z9ˀ~���U����fi�yF����� ��x�ϗ%St���ImURV�y'r��7���z�{ZeѻW���)R��s�p�ˀ<���_Z�rC7��`�Ku,`Y+�,��_Z�������n���"��������)�����Ip6i�mZ�I�nz���'ۣd�9��m���ɀ_Z���d�eW7�d��b��D���~�H�_�4��s@:�����H�|�$�QE!9$������^0	eL����hj�2���a���7WUq����﷒I����D��, ��X-	��ř�޾f�xtJ����(&��=j`֦��J�_JT�Y݁����V�K�]m�u̽cΆs����C��tb�u�:��WiP�id�����+���`֦ٓo��;	~�I0=ex��W�z��/�LnHS�`�冥��0��p�{Ī���=&�Iˀ�H�	d�F93@:�4�86�pD�[n.�4�3Vn��Xi������T��� ۜ�ͽ�?*ULHBB��R7ۻ�� $�P  %�Y�4��ڜ��K�q��+Sv�\Ɠ�w7��zl��\5�]��6��V7n� �km�H��YwTn=�\�ɍ��^�`]qw���4u\�\�sˮB��P�Y@�l�	�9y��=�JlK<�d)�v��7���\��l��x�=����n����s�7��1��>����[!���]r��w'D$;\[����{�����I���C#���.�E���e��8:�xy�L�z�G��o�����ݺ��"��O�m����~�����~{�%IX~�&p�^���1ɂjL�;��oߒ��4W�|�����	X��c�GӘ�=eL�[�	�^0$��L�\��
4�G#�M��Z{n��W��T��2m�5~A�	g�0'��I^0YS��I^�
�Գt�n��]uì��vx탎6Րݸ�F�8�m۞��]f{]��Xl��W��T��������	s��� �Ldc�4��m�=���fA)���S@�z�oߒ:�����q`��-����`OUF���Y�{���q&�j9"`ܚ{e4�ϗ ~~{�)$����"+��_����{y�^0YS ��h��>���~K��H�BN��&���B��C�+�v�Nnz6ٲFt�f�D��sq���s< ��@/�f���K� ���v>�`�y�D� �Ӑ�(0/�x�/�L	�&��q�8ū�ܓȨ����/����T@A�Gl��w�I���he�xL9��N���_Z����dT`[�7B�b�Z�a�f�����"��r����8�]���TH,�"��CR�A7`F����k����h��:���:�n���幸\�_�i�&�K�"��W��l�=�3\I�$�<iŠ^�g �y�����?�y�D����q��90M8h�ۚ}�hW�h�S@�yΨ9j0��3@�������k8:�)K)�J��J�ˀ�d���л�Ż�����^�XEF�����$��%��e��[�Ֆ"�f�,�巤�w�]ۤ�!$%�;X�]XNI�N�'��Z�m�������ˀ��$�_���KR@�s �4�]� ��4���w4�� �2 �&21Ɍ���>����`OJ�����O�!I4���w4	�^0�S�-|�R�I-�7��,��zW�����l����S��B4� @���5��$�
��lV�0R��`��D�+��<�ߗ���(�	J$�ӟhx9�S>���>� �0���!X4�O_���|8����|GHO-	�$�7�n��?&����j�j	��p`��n������@�������a7ȑ�?z�1r�Z~���s�JD"@s�-_3�d)@���P��?k�ݡN`���P�  �
A
���,B�JE!�����R�6��T$~��fs���a����IC��d3$�p��W`�� ���"�	 "ZX��!V��Į(T)�	=�:)�� T����~             @     �               I�k.�Vۀ��&��R[!�K�K�R��Kd�ֻEsM8��$��]�T�����6��]�֪�p���t�p`[	bv���S��CkM�.�SK4��Y��,�\[n��@ڱ�:��3)C��� ���Z����s�\vy�����?.��x�,�d��nwAT���0j�M�f8�X�ӻh�Q�<ls+��m�g-��a)�8^v��v�Şl�m�ְ�6� �H��p�]mX�	U-(�0�h-�%ԥ��s�^΍R��m ��D�����\Vl5�U���n�v���ϞE�R��vwf��w�%�ڥnY`��jT զ��y�l�ԩǧ\����&l��ӫ��k���zw/�b����vvU	�ٺ� V؎�n�)븵k��v�Onٸ5c`���Gl���sss�vxM1�q�smaN%�u��p�;�l�lF+���8nʹ�A��gAҙ6�ZZ����X��� mnuh�|�\D���Ƭ��mj�^]��u��{knf�6�3�ɰHW��r�R�>��ٮ����n��w.�� Ԩڻ[{ :M���oY0Y�����XM��FJڥn7R�r�,��Σ��kp�c^���S��]�-�a;'Vۚ���|QV�Zr�*v^��Gϴ.�nerX�.����4i��8�8�A�x�.9�yuq�Ʈ*�Q�K��u�շ7XVy-p��e�jV�v�q�^��b�1�MFe�Y�wL�R�X�9�O��l��qqI3�"��@}�۾1����;tgx:.�Qm-�K���lT�ɶ�b�D��4�DۓHQ�p0��Bs���64뇬"2��2z͵@�D�]{��|�R�,�M�78,v]�ۛI�[m����6Mh�ٹu��V�����g6͑T�ڃv�$�0T���}Q�~D x��"|
$Q��}Dz)]A��`j)������������  ]��5�NۨpJmnѳZ��зߗ����3:7gQu=)+�tkk�Y{nV΢�m�I�d�yꮘ!G<���Q�u�ї\�.:Rx��[�p��p�X�z%%�f�ne�0On�Yǡ���*�g)�u�
�]e���/[�C��͡9{H���ҡy�ě��Oo�GF�y�b���h�%�ߞ����]�T�Z�Il`ڲY64�d��ۚ�-/���x��I[3��N3"��&	�3�>��4�l�<W��/u��;�Wa�@��"m�`֦�e���`OJ����~��[���	�%���4߯�@���zW��������\b;-_�y&��`OJ�_Z�m��rҝ�o,5-KҼ`֭����]��aQ!&LR
6�<k�V}9r���vR����4� E,��u�"AdALdc�4�l�<���,��zW�L��ܳ�[��+.��I���o1<
�O�`Pbx�R�]t��쏧.F�p����T���}���ٻ������F�.�W����/�L	�����gv��v���^0�S ��0��q����L�W�7/p6�3W ?Φ}*`Y+���u
�;v�PL�̀gv���F�l-����:���l�k
�S��l��4�}�������~���?�|�I*_����7���74���37x�>])U�<�. ��x��ޔ��얤!��h ��^��y�\ �7�J��
��UU,���r�	=9p�=v5�KW�Ղ��e��w���^0/�x����sq9	��)&�_z���Ҽ`Z��Wu�a�����cv\
L�@枨5�c��r�rSd�.��bc08�(�#�"I"�ܚ�w4�^0-L�T���\׼�ū;�,;�,`_J�Yj`Ҧ�J��
��0��"m���Y�Ҧ�K��^0=3�զ����[������U+��7���/���q{H�K,���
�����w�=��
d�9�qh��h�]� �����Z���� M��2-�@��ɓ���d����p1�ш�JKJ��۫Gn,A����jZ���� ��0>���/���:�9"��,PɌ�rg ?�{�U*Wg�_=�_��|�참��NBc )&��}V�}m�RUv��. ���?y6
�M���$��7��/��`OJ�Y*`}_U�uθ�8̎BE&R-�빠�������Z������$� �M+  �3p��$�mͯb�!�/7N��n�l��aڈ<E*��rX���Lm@X-���L�[��" 4Cs�(���[r�r<�뇇.�njm$�m�%��z^��e뵍d��,m�ʫ$����v�Ӣ��jw��~��mN���p�Y��gh����:�������=vz��5��Y�MS7a�6dۻ����#�d��n��$͸%X�!�X�<e����)ܼ�]O)�H��iQ�Ge��s$�
�������@�@��V�����<�gX��bxdnFܚ��[���>���@�~���f��-eK�J2X�Ǎr�����`OJ�Y*`}z]`]�J,A����o-`OJ�Y*`<����\��|�vE�KW�,�q�c �T�������u�=.��ڔ����jL_�LQ�x3n���pz�-Ut�E��[P���aHY�I0>�.�/��`OJ�^�4{-[㈒H��@��S?~��ffY[�d����u�.K�S���$R`�"�;޻�{���ʪ���/���/�=�C�E�r�o��0%L�K��XҼ`}�γp�xdnFܚ��Z߾�~<��s@/����IID�<�=f�X������$�n��N��u�q�XG���2H���Lq!b�4��/t��߼�p���T��?Lr�	jB�07���Ҽ`֦ץ���:�9"��Ɍ�rf�_m��y����("��V�V��30W�S@�������q��&1��^�XEF��~�������:��-�q�I!#�@�Қ�������u�[B��wrZe�p�״���dl"g3���sm�F��fI����8꺼�A���'�������ox�w����oa��.JJ�Janf�_m��bG�;��>�|h�]��Ԙ��n6ܚץ��Q�=+�}j`I�ݪ�Vm�j�V,�����R���8�9p���R�J�B��iR�ԑ���	jB#/V��E��i�{��. �����Z{e4^�JH�c�h��q��@٬�)�`����èp؊s�j�g�nz@�<cH��D&21ɚ��4�K�	������*.o,������0>�.�'��zW�׬߿$uϾ�[�rH��@���`OJ�zʘ^�X�o�|/��Ia����������u��UU*�~� n�rU��r�Q�������U%�k����p��ˀkl�`�$��|�������� 4�� It�ɡ�֍�%F�
��]4�S<�um]��u���|8�Ga2��pV�&2��fq+�-+d3�'��s+�'0e�<[IK˴뱗p�E������S�f�`ڝ�v6�Q�������[���d�en6^͎M�k{X��N^�uu��n���O�v@.0u�SZ�vInE���yc��s�;v5��%�ٛ�����y���.e�	nY���Ū+����I��:��7WA=H��c���� �Lk#Ja�I�|��@�l�zW��T��:sW�7p坝���=UҼ`��ץ���p�ya�o!�=+��*`y_U�w�S@�䋏�@Bc#9,`��ץ��T`OJ����#�294+���0'�x�=eL�$�%˹��Y�s�u*�Ͱ��5���;��D&RzdJ�~_;�����HGC�����|���9 �zk��o����!%����I=��xs�H��d���x��Z{e7�V�%�4�{�c ���0>�.�'��zW��ge��F���$�@�@�l���|�"��G7�mc.+�3n�W�;;ykz�0'�x�=eL�K�m�����+���q���x��E�.{;m�ٵ��q.�v�[����%�.���R�CzW��T�������3>о�Ń�"��MXn�����ץ��T`OJ��7�#��$�B'&��}V���M<y����ߟ� �A��Hg	TL �b�!�@��YRHԖ���ˉ �H�|�x4 �o �?c�8(r2"�ҫ��lO;�~b���OD���!jY��TL`�k��&-xE�C���!�#��������X�c<��$_^����'�[��V[���+
 � �v �T6�cP�5�A
��(�h!�U'���〡��Ee��~!��Bqp�M��<fu==� 4�D��C�D?<E���x�D�B0X)B}j��‬̟�g�����}�S�-�׉rKL��s;��t8�9p��URU��|��Y�mnf���Fe��������u�=U޷w���Y�X�p�ôf� $���[JI9�4v�ӫf`�o;�Ю� �����y�|�=dUUJ����[�����4����I&��}V�ު�	�^0YSL�m���;V���=UҼ`��ץ��M��r�R�CzW��}��I�s��I��M���C����
B�{�NI>�d��,�Ldc�4�Y�y_U�u�M�빠}����H,�$m�Hqծ�\��^�>E���j6�N�����,��ۘ�n1�&G��NO ��~Z^��=�ϔUJ����H
�n�n�n鹆f���gJ���v?9ˀsx+�{-�k'����1�h�W�YS���z�0	7/Tgv�획����)R��sx��ߪ�zW�	3�mXh�u��$�L�K�	����� ��0?O���N���~� $J  �I,���`����Iy�;��&�&��uv.yl)�1��x�������H^M�z ^�n�2�
u������3�JsV7.�v�Ѽ^�2ܫva�J)tGmN��t':��ڕ��I�2ٶ���h��i��.^7e�s�p��sW�'���	�1�է=�JkՙȇI�t���'e��.�1�q<����rsR�{���x�n���h�-�8��J�6��Mۣ-�b��V�q���DV�p�z��p�0,�_�zW��T������	�� ��Xj!�=+�,����;�<���U%Wc�w/,[hZj�q�c ���0>�.�%��	�^0;�¡���294+��Q�=+�,��閆kĻxG$���KX�F�����J}��?���%t%H孝���ͅ���[�=�nk������z��>'76���N�-�%�����<`ʘ^�X�M �X�������Dۙ�z͹�|E�`��`w= Yw+��Q�=+���/,�n��݋�I0>�.�'��zW��T��"Ϳ���`�wo-`KҼ`ʘ^�Xa6�$ �Xj!�=+�,����u�=Uo�{������5f�-Р�sգ\�k�\�g�gsI�[,�:r�t�J�n�mւtvF/ܸԳ�	������Q�}.�ݖ4��Bc ӓ@���@�*0/�x�%�0=2��x�ݺf����������ˉIWEB�C��� ��e��o$�~ϻy!�揅�w/ܒÖ�Ҽ`��������yb� �LD�o35p��J{\���À��h΅�1G1A�r&$�i$s1����n���k���2L=�[ħ7M��)��Z�I�}��X����� �T���i�qo�,��Z��*0/�x�%�0/�]`M����3�a�\������.�%��q���Y���G3@:������O{��rJ�����H20`(��;�w�$��XVӈM�����Z^��/�w4�Y�}����(5&	�DӮ��l���v�T���`�i�)Oj�@�V�9�&HF��,JE��>4�. ���_����jJ��k36�ua��0/�x�%�0,�u�,Tr�*Uvڹ�����5yy���ɁgK�	b��W�L闖�����bŷ������W=�_ ��pҼ`ʘdY��Ӗ�����	b��W�YS������{���}��ޞ���w�  ��mp  -�o!n�3���am���S�]s���k4'SsU�
�^�0�y�2!�k��/}r���%���2쭻U.�DzQye��9zֆ���"ԠO�A�6�f�X)�n(�5�&6x��y��-d�r�+�<�	��V�Ӑd�-�',&�;g��f0�0:��km�i�p�5���)+�kGm�n��C�#�>s��ͳvY��[���=�.����.s6�5��]��'*RZU���@���#��}��s@:ʘ�.�%��s���sqn����0	eL�X�F���`�Bn@x�4��<���:�F�����[��ąڎIa�jZ��*0'�x�%�0>�.�=2���_�y~Z�n������ ��x�w�y�Y�}UU&���xe�/U�m�X���2�Kv�npŧ����^͸��N:m�D�iS��
���o����0>�.�%��	�^0=8�ui���ۓ����'��{y� z:�� ���$��IU/�I~�k8������9vr�DC`�6�Z{e4�������u�6hbB��Xj!�=+�,����u�,T�:�9$�,�d����z����X�����m�u�p�5�]�����l�������6(�:��:IQ���'��1�$���NM���X����� �T���C^����tԵ�,T`OJ�K*`}z]`ze���v�`���rҼ`O{�w��O��T4t����:��@�e4�su�6�
"anc �T������*0'�x���PՆ��-GbԒL�T��*0/�w4�Y�}�ߧ�$��"F���qYl�Z�"ɸRܛ������qs7l�2k��Y�2$��0s�nO �Y�_z�h��}*`M�
���;���`_J�K*`Ҧ�Q�nq�ǑY?8�&h^�@/��h�F��eF�9i��a���L�eL	b��W���~���D�E% �@$` g��L	2�5�Q�,45bL	b� �y��?=����������M�ekI9��+�|��s���vxܢ��ɮ��ٛR���ӏV�jI,d�H?9ˀ<�������X8� ��{���Z�����~{ҩ%Wg�|���{�s@����R(<Z�I�}fT��*0'�x�%�0=�,u�h��Y��x%U%V��p_�YS �̩�7$(g,X!fj/M�8~���l�q���i'�o��O�EAW��EAW�"����"��Q_�DT�PU��PU��UU��"@@�@�PDPE `APE c@��@1�E a@�P0E a@T�E `�@R*
����*�*��"���"��Q_EAW�_��"��� �����*
��*��"���"�����
�2��G���������9�>��� @  
        (�     � 
  xE
� �(�@��
 ���T%U%D@�J�ET ��*� �(
�A\    �$  �(��2�c��w5�u�N{S��v�0 (�}�������yL��p ��K��rz� g&�' ���t����q��6u�ܯn�7t�� ��8�q�0�z����:<�P 
 H(�b hy�>�>���p��x�S��z��Cm�}���   �  �w����z ���G��]׀ ]^g�^�OJ`�;�N]�U��׽���:\wJw��@�͹�飏s�qqז�j�� ��
 ��@�
� }w�>���^��u*�gu�����{ϠP{��\��[sc�ӛ��14�����S��  ��)@ 1 �0hT:R�bhL@ D Y��G��pz � bh�@@  w( )@ 
HS 	� ���4b ��� q)������@��I�a��7�3qy���g^ n-Oz�<�� Ξ�7{ܮ�wo.�OEۛ:מ�U ���r}����/ ��K� w�  � 
 H |��w�O}�>��:�ru�>��W�;R�w>^�O]��/+�xѣ|朻�� ��ޛ�x�t� Ow�..�����{5���������9}.,�gx����l� =!Sx�*��db41�P�yJR�  D��QD4��фOb�P�) O�%O=J�� ��	��	� ��t������������՞�{^��{?Ъ�+��_�*���UAS��UQ_�
����*���T>�����W�Y��l����,���0�!R!$R�\S���34� p܆��Q�@"2�g�g*���u˄�]�ՙ��t�Q�.���z�U�5s�U�/���Qx�3���%��o������p>HXR�HHLup�u�K��V\¹zl֠K.\�5����*c b��O���(Ek�<F��޳Y{�2S]i�kZ�2j�
+
R�l�p%cm�$i�Y�%�@H��ic��)P�T�^�`� R4H��k
)$��� H�$�j)c�u�o�aZ��
����HT Mo�sG��]$��B�=���N�@���_�

1�X�dA$,I$f2�і-Ԑ%���l,��k7~�w���Q
j��!!!�0��5��M!+0�!H@�)a)������B����=����SGXB�.:�q#	 ��\t�$��<D�D(|��ݺ�$!�������BT�HT!@�)D�� � �e>m�F´��T�
�@�%VLiK
s���g	&��F�#&B!p�(@�˞�p��G�D��G�āġ�X��8���ԁF�I�,$K�#�:<�p�����6 Ќ�� ��!IY��	�M�@"  ="Q���HP"�:B��3[�w��}�
1*�X��=.�I�s�s�>������!z�	%��a�g7�BU�R*@j���S�X24�h�\�R�'�~�5�(�]���$!E�j���3�&�B|��(*�PȔQ"�4C_=~���B�J!�B) 5�$1�fB����k}���}�ݳy�sQ!&�߉���5��7����2|@(l�ĉ�&�HM�}�T�ɑ}���I|D��B�aB-�X��HXT���6���jC!KY++��$(a��x��)$�$.:�G�A(f���Ħ{� 9�y��sf�.ok9���s4֌$Hk+	�,�zO}v�0���p�#Y �.i�D�b}���S	1`%,���D�
�	 H�$�B	�(��`D�0`�H�#$LM�K�kkRe����>��1Q>	 �`@`?�E"1���,�� �B2! ����J��aL$	[J@(¹�f�@�x�<oz)sN��� Q�p�ف�b1R
��VF�bB��E�.V!V��q���$�!�LaInB��t&�P�!k�����y׹��6;Z���L(Wa��#�`F���WS��t"�сy D����<rM���dO�KjF���Ŭ��E��²2�,ag]����0��ZɸÆ2���Pk��]r���e$���¹���3|��ٿs�m�,ln!r��@���#@�aP#CE�7����/���S
�����,#	��JFN�xV����c�|����`H�%)�`�#`Q!V�E�� �XL4x��RR�H��G��Y������K��5+)B�Lmș��57��)�%�\3[���<8����4�P�в�f���.�����!�K�H��%��LtK�7{$
��$�H1�ĤH^,̚�F�:8�T��͆���'�01+ T���P ���Lli@���5�.�0��w�&�gHOk�sC�"XD#�s7C����4c� F��B+�2�.�]�n�SM�#I�}�s�ɫ��B��,�
H��!+		�z�4��s�XсBb�#$nB4"@�Q�����0�-�5�p�a��a��"@�Ff�IwϞf��_�ώ9��`¹3gę��a5�����s0��p�s9��0�f�S1�l+k E�Ւ5�H�`μBsQ��SD��H��I ���X5$$�0瘲 �@B�a4��)iՀ�"�}	 �+! +� �KJ��(ZF),F�,hc$��0��tst�wy�p��X��S!Q�M++�%�! � ���zI D*���B:xh���F�m�\澽3I���!m#	(V��� �$$��h프�	BB$�c0)�,d!]T�P vj9Ӓ��Ҩ�����aD�#1���)׵S暎��O����\�l�'٭s�X_��^�����F�X�~�r$D⦛o�	�ڢ��N�dK!4�FXT�1��.���<M�U�KT����~�c��ȕ+g҄(B�����X]�!�4�c�6 �		"�!����h�3�p�C�H\"���(�ʱ$l#$BX��$"�GGC�ybA�Ú)�|{C.V�`E��HS�=҄k����8�c� I#��l S,J�:8;415�+�� L4m�<p�4���A�H�,��� ClX!��n��!�RBD�$ �U���X�����sP��4F�� Q�F��f������,�]s�4Bfv���V�~����<��`���$jD�J9	ЍL��¸jI�4wz����rI�6C|�6ky9��C�,3L!�m�$��K���O������������3G�4C�w|�h���p$cB$2[����,b���<�y��*�1bL0���$������#H���&��!4�ģ"MҒa,1@I �0,F�2���
XF24�	�ЌĤ��T"k�%#B`FjHY���S�"`�İ�H�F-J�}�!l��JJl�:� J`l۴ޛ `���L�°+
���\rE�Y	 N/��9�8�#bz�(H���D�(E KI�$G�B,J�1k$���FE4�(k����J�,JE����h4$
0+�M�Z�F:����cBH+W�	$p��\)$4���-�r2�EI$Ⴧ�$)�8��V_�&��f%sLi�
`D� ��$)��CS{w���~�q��B%P�P�I@�)�@#����a�$�$$bV��iU�HԋX�
�	+i@���.K�~7ɐ���v�����DbH@�@��u$����n�L�,.���(f��)6tk�v�|��<��;���@�!���i�E%p5���!��V�)#ْ ��I"X�%XW�BF$�H�#
9M̜scs]k�N��R�`1Iԃ_�Ċ`�R0��)�Ǧ�	�B,�^�z�)�.�	H| B̆�Ʉ����.B�kDִjo���X&���v�(��6c����3p�D��Ja.��1�,!���8s59x|��>�O���y�Jg�����59$h��h�`3��>��� �a�-r�$��<)��/�{_e���&27���XK��&�q�4G!����,f�����jF��1�HWT���\>�����ę���k���9�HVY##	#m>��~��	��}�2>��:zQ�$,��P)1L1�Y,*�k"�?~��o9.�B�g��\VQ�pԹ�35�p�W4L�Row�$20#D�-��Q��Hh=X��K��g{~��:0���� WP�aXW����7L�Ͻ֖>�n���%,�Mj���F D�"2V��"L)�`R��#�)5~ټ��Bi��6A�1 ��Ȑ�$*@�@�-��	hH��1�� ۚI���$��m�d*ƾe0���֒E�5��	��a��"�	�	����:��ڤ&�D��UP      �  �    � �n 	 	 �P   $� ����  �6���cZ��N��4��)�8z�� �`�`�oIKu��Rkz�V9km-��A��Z�m����a��X۩:�tN�.-�u�w;\�ۓge}�;��h��V�j�.��3���6��h��U��
P6�i2� $X��7m�[5�.�)��91I-*�����ݸ�,��Ѷ� ��ڶ  �}��m�  q�N��    l A�	Z����DێT�V��)@��:A&�M�L�d]��%L��n���-����e�-����Z�m1���R��)��	=-UN��8�;0)KV�6ؐ -�l	 �&ٶ�qz�'@-����[�h��� � �`�ݱ��b�uUR�-�[@ձ6� 6�  ��}��   ���h�l�"H�m$�쑭�����UUJ�J�Q�K�h
U�F%Z�j�Um �m�ն�m�m�m� u�l�u�m��m�H��� ݷ����m��m#'TҰ�Jٶ@� p��,�@UrUK�q�� Y�X��$IJC%l��kր��   [_ǀ�ɵ�8m�	 8�b�nڻ6Ā p ��Ͷ �l�H �m��lkX $tu�RI4�'D���m&ݶ��� p h�Y�]-�5��j�]�p-���:q3?i����Ξ�ˢ� �P:_��wL[�ٰ7"F^V�v6"t�k4�3E�� y�m6טH�S%�J�(��7+*���UU@[Bu�:[BA���m����_\wֻ@-4���lUm���� 
���p��X� 6�M�9� �v��m'^�ۂN����K�֪������HFob[��VvxB҂�J�UV�v�Z�5;랩�[ j���ɲQ;5@T�@˪�Mȵ+T$H��n����Ź٨3�ڥ�č�rp�E]Y+lUAD�Xj����n�i5vc��1��6T]<�6��e)\u�t�� ��»m��-j�^e^��'9'EJ� � �b	��ջk]�94����o)�@��Cd
��Q�yg���D}ol�a�B]#F΀�0l��-�ɚ��U��vx:����`+�@e��`��䀋h�`A�M�[@ -&�E-5�� �@   $ n��0[@$ mH$�[p�Z�t�M��
YeN� �H�P�:�ݶ���� m&�m�ѥW�A(�U@���  ���ͷa�0�l34� ��F��L  [@	��mm��!���7�U��q�]g�����a�mm�%� Hm�m:�-m�m�   8	 ��l��  ���,�p�d�v�u��;$   q���~�@4V��$   �@H��l6�m�m��  �   $ ��-�<��ҭT�R�/[� I�m�ͤ؛] ��Md���` ��dH[m;`m�	8()i�T��U��Uک��-��n�[i�l  �� m���Vؐ[Ko[@ ��m�� 	  m�ɪ��)V�ݦ�ۤҰ�5�m��M�mmm�	 h5���Z�N�[w2��9�� $M����	Y�jZ�v��@�^b�:����V���Kh*��PJK6����u˫�f��*����~����ͫ�����-��h��m-�^ۄ�R�R�<%�j���H#�N\ ��H�$ ��1+]wm�:褒 t���������X[H�oH�`<6ٷ,J���<mU*�q��]��m*UU[C�U��l�M�Ul�`�/ s�6�Ai�
U���e��{GS�1z1�^g&�kh
�VU��6ϕ�L���84u �v���T��!*���U� �ݖ� ��R�]<����7h.I�mHI����-���V�*�A�*����}�ݖ�`-� m����)x\C�J�6�zَ��UE�嚨rp4�!n֨�m��+�m��-��g&ǡ���c���-%���P   �`��l� �i6�Y*jp���+Z�행�j�`��]�yy꧴U@�4.���-�ʜ�cj�rn�!��`�/YG6�v�k��O��vΊ��۶�@V�Ɔ
��  (lvն��@5U/(Tۍ�+g�K*m��k]��tm� �    ���  �
��TgCr��iV�� (   �� ���FHp�x�v���� �lp  H  [GHlm�٫i��l�m�s	(�\ ΀�� [A���p   u�F�6]9vH�ލl���h�M� 3�gm�����N m�����  �R�M72@  �t�2�[v���` hl��G[��@J�m��#���m��5�(8g@8<�۶,kN�	 =���hj��v�f��۝z]6Zu�v�9�,ƶՆU�
��:ts�T;�\�f��%�-�jg���
2�5@P�r̹R$[K�b����U���'I��ş�7�p $H�'8   �6�  �ؒ���8��:a{fk���*�i��M/3m�  BAɵ����[nղ�]�6�ܶ�D�!��lUR�ʪX��2ǎ`
�ꪪ��M��:�8着$��I[ 
Sv�͝ֆ��J���UT��$$ ��#F�J��1l cs�e��U��$�m��m�q� l ]Wr@6ڪj^���7keT#/���|xN��e�m��e�A&�ljV�sm���ns����[Gᓝt��l�l��/TU2���]���` %�li.� 5��$��mڳi1m�m��Zl   �a��Y2�$�[S�i-m�g-�Im�n��v���NӢ;I�i-��]m� ���U@UW]H�"�	�d���M����]T5�ÌC����R� ���ҥ�z����8 ��k&��-����� �s�ݬ���  �:v��rX9�-'h�����h�פ�Y&�]WY-Ŵ ��e��k�ZL �[@6�@    k�H�۶��E[x��&� �igQmBFm[@ p���lH pm
�UOe'�eB@�b������-�A��m� mN�T���R�ڝ������r���� ��z��l[S���ګkl��@   t�73["��@V��{+��N�n��� Im�wP9�%��m ����6Z�m $6�`6�  H-�U��$m&�$����@|�_��� HHh6�nl�-�   ���u���ٶmJ���O�6����S#ʭ!*�n��݊��Wf���``+�^%�"�n�{&��		5IYm�ݻn�i�I�� �D��kXm[o��� �`kX�R[wUk3m�pUvQ���gl*ʷmU�\��4�mB�2��jVT
�UZ��
�h�0�kHm��-�qU���UUY�p@˔V�#���fճ�/k�J�]!*�p
�[UK�	i��/[�w_���t5)$X2s 6�n��lX����M�  6�m���88	V���VU��*��5B��q�m;d�WZ��e�h$"Ͷl$��ӶY��ZĀ��m���$`m��	n� l [h���Jؑm�m �l����`88[@   �k���d�+n3U�V�c&��ebҀ@�d�؜�v 6ؐ  ���@��@ �vҥ�s�H,�6�	Vs=@W[mJ[@Դ��!��R$�m� ��ٷ[%�i�������˶6e�� �,*�.j�kJ��*Ү�F�\i���4ۤ�� 8 � I��e�l�UU�ʭ۵T�(�7�o���e�v j�N�� 88��հm:m�t�I�  pu�H�n���з۶��$u� m� �e�[�ͶjƳKgfsEh-�2�Lz�=yV{Eu� P��qV0�` [dm��B��<�*�V��|lc���V�$�i[m��Kh��1��	յt�z�-�n ݲ�  -��'D���` �` �խ�m$m�`'A�� �R�m�Amm�ؒ�dE�&q��� @p�f�����m�j�N�� Y�$87m�,b@[Kl㘓�	a&���H�I�ʪ��. Rΐ�2][U^�J��۶�$h��m�ٶ��l�p��m�9��Z֐   ݻLdk�������[@ p8S\�L<�mWKs���`+�lE�-�m�%��{���¤6*���J&�F(<P(��B������;H�H��M��6��>@P6���'C 4���6	��ЯP P���R��*	�DN��||�Dx/�G��@�	�t ��<Gx��1`c)0�1@�(`��`B $�K�uQ����p<��S�M�yE:'PC� �+�c�@`xI|����(�C���!�h�@FE8*�W�Gbu@6�t*�p�A��Z��<��<N
��@�ǣ�`|���QS��M�#E ���UOPM(yi*��F��A@��G��V#�#��Eп
���`)�
�+G@�r"u�mV��£����� ����G��uZ������"z*����B)�!�(,
��="���`����@��C�."��	���GUx�H(5D�>A`$P"� �b%MU�C�=DN�v�R*@`ki�E�����P�������BP� �#TzXU����"�d�/w�)���!�@�6�
�EF@A"�O��P��V� `8�u1D]@1��D�A �t��@��������������@��1DƫD���Q(HZ�@�E����E��`1ZA(A�ƴ�`�@5�?k@p�6�m�mpH����1�Iݶ��R�=f�����r%v�ۦA�����6�-�mo0j��*��[;C��nv�6�m6��*��w�m���9�VBn�����mA�*blݷh����1ecR�t����m�։�T����٭¯���[�η]f�)6��8�E�\�s���ήcY���8R��v�t�qvV��Bs��b�۷4m�ˌ�q�Z�F�X�[k%���x���6���ӥU��ed)J�>z68�N�x ���w��K7@t`�gJӳ9iWm�tQ�vQ��k��b-J�e��i��c��Pَ���L��"mmWU]nQ�R��'d��v$ջ�@@[��$ض����ҙ�pj��9sHn�v������5�m��l��R���DlІz�o,�@���n�d��˷J�%���a9#[a`yÂ�buX�o&x�m�nI�Y,��p�hح��q�E�H Xg�]6�չ�������6�/��t��%�ې�r�a�l���l�7(��m=�w3�5�x�ۮ*�)��QnMd�br�GN�dU�]�0Q4ԏO=	�쌐���` ��:�����3���Kʭj��9���ʠ�^tX�6ڝ/���t�YY%M�8�tUzK]�����Uېö�l3�,�"j��9�۴"�Z�u5�X��uOl͡�F����7�/oe��Z3����-l����ꦐ�@�t�zڝ���6}6�[���X���Kn|R�q[D���\��aqv)��k�b�/��Ku�z�Hԛ�h������R][�Ԑ픡�m�i��Wbt�*k+�FI&gt�h5{i��i��"VE�d��R˶�X��/=Rj�βu ���ń©��$��,u�:ֶƨ%tfڑZcBV��v�3"��k�0�<8�M;m6-v@��D{T�*=�r�SV�^P�(�T0*���ʨxGJhP�N�;P҅O(�A<��A �Eb4����)ڔ��ԅ�N��Wmt�݆:M����)���M�pt���y�����M�.�m��V�2��!����dl��ڰ�\/m�,��-�Y,\����D;/Sl���U�uѮ�J+��ϫ���s����]U!���t��}�ΰu�m�a�Cs�A����L�����Ap=r�؉�R�Jnӎ��	��qY&f���I�&��e�6
�PڅP8#^s����e�2ffaf\�����.x{v۝�]�
c� y��1f?�x��Y_j�;���|���~AU�����$5��(〆��-v���g�$q�ՠUmz�ՠ[����D�O��h��V�U����V�k�h�Ux�[P��djE�Umz�ՠZ�Z��r˫@;��pM�`D����������v��`k�ٰ9DDB]��n������C[�rh��*�tC�9���k��'��Yk�1ؒR�u
�v�����8��@K�b����5QLR5L�Nf���'5��#��"
�H-U�G��5< sd[�=�ڴ]�@�s��F��y�y�h	rL@q㖀�$�8�|}�V�)�S�uS`~��w�Bl��`}���9B}=�6˺�%�$�&〆��?[)�~��ZW{f�����J!C�|�e9M��n�R����:�NwZ�8׻:$�顮Ӹ�O1=sgI�H�bI����r��uw����V���M��l�4�b���@;nb��$� 8��^�꯭}��	�F"$�N=��-������]�� 1��C^s�s��?.����iVL��jD�Cq 9&�ǎZ�sx�9�S��bȇ�9�_j�:����}�@�l���eˤ�'�0I�M��2Y�6q��yLk�xR�룗x�·��C*�N�nj���3f�������h��V�g�I)�2'�@����M�����w���wf�����IL��@�v��_j����U�y���h�gn=�8ē��sv�x��1ǎZ}��:��8�� x/I�k^��IϽ��2]����H��k�?u���ڴ�}�@���1�'��d���Bx9�j����.�^����WJ��i�Zz�.'n�t���@q㖀s$�9~���aW��z��y�&
24�Cqh�%�8��@;�b��uUUvs��'�ő�Z��M����]��h��Z��i�b�	�28	������ �OZ̒�s`�8pX�;��/���#�9�ڴ]�@��)�~�ՠ|vچ�I��������J����$4�*zw�`�V����*�UyϞoi��i����sY�,L��O	G�p a�s���}��4[6������S�܈EZ�6HC��Y�B��ף�(�']a�q�d4i$���C�k��٪��3,�c[pR`��n�On�q�u�x��Sr6[J\��OD���-�����B�͵������{_#�N��)���`����cO��ێ�t=LL���p��bR�����8-��6����92z�s`���-׎Ze��6E�<Q8�ݲ����9��-����}�@�-l޶����s3D&9h�r�=��l4���6(�Ȓ��H�=�.�|�z���M�ڴ�ĕd�`�#M�7�oe4ݲ���h��vBP�̮���8�)��$t&��'U�]p�]�{��D������d�75g�.�q�őr����Z�V�ξ����ûk�����ҙ�nf������:�><~��D�!*�C�a%�/јNO���+��mi}
!����T8j�5T���v���?v�h�ՠrٍ�J���h��a�!C��������7g5���Z��WșǍ������-#� ;�W{Ww��C��on�I���b.ٹOqv	\W e�
����+�˓�R Ϥ��������9h	2K@rc��9%J/2�rZ��QSUN�ϧ5�B������w�@�ڴ��+�|�Fԉ����'���ܓ����!~$Ra�R&fnǵh��Z�hjr}�Y����/j�-v�����j�;ô�5�i1}���@�ڴ�ڴ]�@�}�@��jX�a���<]kv:����)��l��l�����7�'����H@�$��$Z��Z��/j�/]�@�lƖ%ALRGqh�S}�bG����^>ՠ\��ǲ&F1�M�@�}�@�v������h�kcX޶����@�v������h�:�1�.E[��~��O��Ĺ��2��HG$Z��Z�=}�?�yh�ՠ~�-�<�&FblDl�m���Wxw���������AMQŵ;���%$M�M��_O�h�ՠ^�ՠ^���&A,bȇ���h䖀��s`��(/2�Ѵ�� ��@�v������h�ՠ�B�Ȑ�!��z�V�{e4�j�/]�@�tIaA�RLp1G�{e4�v{����Z���O�2 �(D
QP-���~����,�U�e�v�U*Jᕎ�3�WX)y5֞'��r�r��ӝŊ����/W�=�#�L�۹ɭ�:��]�c��Rn:B��� m��������t��_�w}���]�}����l��]W`��`��D�S'��%�9����c��	8.�i�]v
�[t[.㝛GX�@���Rc��(O�����]f�d5s2\�sZ��Wjg6^�X�*�kl\�x�0]�.�Ls��س���s�d�;�ʣ�(ީ�����C�9�[~�c���$�x�#�z�`�7���C�D��/]�@�}�@����h�ܸ$�YS$qŠG�Z9�@N䖀��1 ����'�#mțx��@�l��x�Z�z�ϱT�V��v��&A,bȇ���;�Z��x�8������m�}�'��u��5��'Am�	=��4����ˮv"g��9ޤ���� 'rK@q͇꯾��XzI�@3�B{<d ����*��x#�R��A �Q�T�H �Y"#b����y�W�mU}In�@N͂����1(9�I�D��?v�h�S@��k�*��@�[����#�m�#� ;m�@K�b�l�c���!�'$�8��������l��[�4}�Ξ����id#cx����N�d�0�ʎ�㤖�r%�\s����i��&��Ȓ��?�yz���e4�٠qw���fT�L`�jDܩsS`~ͭ/�CaݽV=ޛ�������/o�S� �H�4�q�@;����'5يW���ED�(T����a9�����ع��.�"�P�o4��b�0�5�([J��y�aa7����I�(	�l*�_�ƢE���y ��"C@�VR�RʉJ�I��g 8B�2}�d�.��lu�ÜvD�����t�xD�^!�.��D�ǉ �D4T8� ׎�+��aSȝ�+��7�k{��� C���(p
B$�D�H0}D�Aѽ#�Ѡ�M�y1�'P�S���Џ�A~J����:�ōT��	
t��|y"� ��)�U�Ī )�HP���IGo:ܛ�k��٠7#vRjH��������wzl}�6�����%�S>�z��M6��¡b�n=���}����޾�{^���n�	�mF4�I��:�c:�so*q�n�ul�k��Pw�������Y��lؤ��dN?�r�x�{f������g�^�z�{�쉑�x6���~M��zl}�6����铷ޙ���Hy��4
���u^ק�������@?w�\CDmdIL��&á(����`}�\XnmX\b��
*��؁�mC�PO��~���?w�?��\�P�ʗ56������%	(�����5�zl����łmʢ[�z��np�7����u��6ܜ��5���`1�v4�\��$򈈈�wanj���*\�������`|�6l���$�?0�z��3���)5DU:sU`|�6o����Os�>ޮ,�j���B��&�a��ANjf���BY��?�oN�Гff�Xz����aF�7��#�C٘��y�f�X�6l9Bew;Wr�]UL�$��\Ӱ�ͫ�B�B��z~6}�`f�k����)�!:4��U΋ե�bM�����^�����-���@ȶ�-��
�R��΃��ֺ�����[k���swX1�ݨ����;}�뛻��v��{��øt�4s�wE�f|C�yv��]�f��˷@8KK�	�@�v5�n&R�(��(��^���8�f�Qmv�v�&��ն[�s�N����B�̞�k��H\M;r�%��<�S�܆e�r�X\��W%�����{&�����G<>��{jݷi��޶{qD��䒁������u�����f�X��ɒʙj�S"rG�~�o��H�w�@;��u^׾ϒ/��̟4F��i����y��f՟�(򈉞~�M��>�?}�Nv����Ir�T�;I%	����C|�ޛ��a�	BOz����w m��ԑT��U��sf��/����/���s�h��%`b`%�-���3�f9���n��֌�`����)[��P�Zm6��PS�����=��͜�`}�^Q舄����������)�2����9��!%�!	@�DR �W�`��D9�3�~Ձ���?};��	%�$�N]�򺪙*I%L��`��1�l��(���f7οyh��h�UhC�ӄHx���Ô(Og����'�����:Iw��@9�}�CDmdIL������`tF�o?���`c�ٰ<��[���񿻛K���#��@���W��n9'�=�nM����du�X.H��a��μ�A�D36��g�Z �\���z�aמ��<��Q��[�TSS�.T����3z��6omq`}�����w͜��	9�Ō�D��/��~�is7>���E  ���"@�TP�C @���X��?(Z�V��V���v�wU�/�6��lJCCع��-��- �;f��W�|h�$���7���-�r�z�{;�Z�UUU��FV��1ƓM���)�	s���ƻ�év������i�'�k�v���V�t�<��| n{P=���/�ܰ���@w�y�cn(���h���bG:���ޝ�`}�W�!&�3�%2YS-Sn�34�ͮ,��vr�	&ϻz��|���+'��sN5!�숄��y�ݽVnV��!"R0��DJ5��~R��??}�o�{�4Z���A,����#qh#���UT�^8s| �-��������ӑr'@�%Q4�9�������y��݂�< �Y�Ɍ��պ��{�__{;�ָ��������� ^� �9~��`w��@3�%�g� D�7��vS}�Ӽ��ޫ �ͫ�	zd͕ķ��50oR�Z���?��H�}�^��@�h��H��<m8���Հo۵`g�ZXr����_y�����7$�6�)MUU�o۵`z{��x�=�M�~�ڰ1B�D$!(������Z܆4����ȱ�$m�zڀ�m�=Zۆ�Y�Q���5
]��].�n���\����)��:5�����Y������W8�Xdnܨk���3lu4�����m�@-���ۨ6����	��r�a�g�:�+[��FNrK'NS�U�dn�>����]Ӻ��/F��s7m=���7�_|[T�L�O�d:�xČ�-T-&�]{���q�q秝�o��nv��ܙcu�z��:�v�&�W�"���k��y�&����u���_\����������/��̟<J1�M273@���}�$��`��`n�ھP��3YNz����\�M�M�woU�nf՜�P�v�s@���#��3���$�)&��C�G�P��ޫ��Z�5��6�(IC}��`sm6�L�5.j���V%
������`��a�_��c󷃇�P���=N��i�[q��v�i�8X�\�O1)��\}�w{��,|l���23K��lw6�s6�!(_�woZ�9o"YUU%I$����ﵳ��jT��|$CF��R�E�uF
ELG��v��C�s��=}��U�^�������F��$?��h�}4{w4�%�������ߞ!�6�$�&���v��`s���ڰ��f�X�H�'��sL���*�k�<������h��ht�O��4�X�P��\k�������=��Y"][�3w66b��H���C�P�US$�R����z����~ �ޫw6ס/�5�����A,�QI�5SN��7v��!��zՁ����7sj�"a�6�aˁ�sUSU`wolܓ���nT�9b� ���@��?�>�g���nI?�}4�Φ�TL��Ԇ������b 淋 vI�=U_\qx@J�+��FF1��@?^٠{��1_{ӀG<� �I�GW�+j��3+6�ci�;=\��7;���+������p�(�t��~���0�^$��ۍ$<�$��/��gٶ�y�=	(������3;�S%�2�6�:���3��W�^P�L��ޛ �w��>�ھP��{i%D��I���K�,{�6�f՞J#Тg_��=}?�����Dd���"��gى�oU�Ϸ��߲���P�6!j�*i�4��+�C�@�P��o8�4�����E1f8��h^��J=�߼|�=�`�mX�����;r�<k�n3��H���2����G��ZX�Y��������}�h�����s| $�- N�����Xz��b�V˖�0�Hi�e����P���9�t��V��D$٫5�ʪ�*I%杀voU�fn՝�>KݳƁ�?yh�kē���I�*���JD�w�V��Ł����(Iz$�Ϸ�V���S%�2�6�9���7�,(IG�Q}~���ޫ ���ܓF��t�a߉)��X�c�>å��ҝ�\!� ��e{[��8�P�P߅��A ��U���J`�K���zs�C��iT�Z�����@��b�;�>��?���[�mpM���]+�l����v���{%���l)Q8�Nz ���m.94��l�A[UHh���{m=���p���ݲITFڀ�k��Rb�2���r6�k`����)P���:ՖY$7Q�*�n�Gm;��Ue۷`�Vi�5J���h�l�NK�kN�n�D��v�EA�������\��e���r�|���v�n�1A��d�ѵ�[k��R#�4�֎�fn.0ҽU��S�n�G��n����^����cp��Y
�]Om/FNJ��&N{g�j) GIu���Y�c:�6�P��%�Z:%�n�t[�L��C�Ҭ��m=�cC-��Nݥ(�87N��X�zI�㝎�nw���3����#i-[�۫6���Ƴ����\�Yjd��gk[#���R���1��+6��=c��o,��F��(���VuyUiQ�(��]���{
w���`��1pd�K1�\��u݄+�[m��[l�&��i g��)�D��Kcy� l�@pJ'��ݣ�/*�!$9wf�o��tM�<�,h�`�2�zvN�ixґ]��z��\i3	��iVy'eJ
��.8�m�Y��t�lƄN���us��
��	$�i�@n�Ib�ۍ��u��I#]$�ͥ���5��ʸ�9����#%��Y�2������Y�ʍ;j�7@[�����N�h0=�ڂ�A�铳V��A�wm����s�Ujx�Fe�n�7SH<�MNh�}&sm5��
��7Pc�f��Vu����x�f:,d���qg���ce�n�v3�#�KjjT��v#C3�e�yy��:	��^f���zq%(ZI]���3L$���,�=���n��״ESrm7b�b[�����l�q��j�mڞ/�|����;Oh����k=XQ#YZ˚ c���}����P���J��ݵ��3a���\�!gC�OV�/' K!5MB'_S��{�����:'���] @EM�v��T�������p<#|(|�U���Qp�ɩ=�Ժ�m�M�n��M��.̼8�p�t��DKTO��e~�#ñ��fڱ��3�N����^r��;m4�;���3n���0�xz�����ud,��r��S���i�c��Af�� 5��]�����͉�&�GEȬ����7:TB��J�Zl�A����iR�Z6jI�k��\���݇�;<�n��U5ٔ��w{����{�Wߨ��'c�a�q/b'WX):7Zp���s��Z��%�ljj��O���I�=d�⍧14�R�?- ����=�~A���@�o����FH�%H:�`�m_��L�w�V��Ł��V�1"���C�LY�$d�h��7��Vt7�=��;7��Ƶ�a�A�uD����I>����������V�!7��V<4���6N^m 92K@z�﾿9���ڀ�qw�o����_���^[D���0V㮘C�qv'�m�:��Z��GzQ�Uo���7o}���$�K��;7��33j�߳myDy%�����=��M���sR�&*��䓽ﵽ/تؠ�"�i�qU�*!BK��gv}j�ޝ�`�m_��2�z%e��j��9�������]�O}����M �ޚ�f:��Q�擗5.���P��f�Xf�XyB�P����X��-�TST̒�/v�#����U��o �yR�$Z��`�Ǜ�IG�d�$�����;�*�^9���&�j�N�'����}vɞ��ҥ-5_�7{��߳mXl�DDz} {{�`s^byxL��r��߳m_$�ft�; ����37j�	/(�2v�Kk�%�l�sJ��O��$�����������D����nI��`j�@Ol��T�%杇��B���o�V��U���ڰ��
!N����<q��m!�#�@9޸�������W s=�@�j�����d�\����Ԇ�����y�[�n�$�j�]�wW�1(K������a��]�� �<�ْZ }�}�}_r��{P��ײ|�LNbi����v��ٟ$��`��`}����&���e["�lx�H��ޚ���=��m���Os�67u�*�	J�Ժ���(�D�wz�w�j�����?B��B�B�X*$�EbR( �A
���@@�1Z�V��?"'�k��u�'i�a,�^S*�����77mX����y�����33j�Ź���)��-Ԓ��u��4o,��"v��Sul�k��Pw���/��/�i��,Hs?�?yh-�@33k����Vw gYSU%I-��v��W�%2��=�����پă���I��q��1�&�v�M���=�q_y���4��"*�h����O{����{rj �vh�W'�D� �b�f��vנz���_�3w���ݵ`\$BP	A�B�X�
4h@k����Pv��5��q,˰��ʶ���'=�u+�EU��7E�4�<��⛝իuM;�k`�`�Að��ckpc���J�)�m����:�%Z=Tk\n��c�4����Fѐ�l�]�����cJg=#,ڱ�ѡ(��\�2t2Gc��O6m��Ź�v���-��e��8�t�o�[q�;��u�Fz���.�mѴVw��C�5�Ɇ\�dz+�6a�im7���ܓ�:��MʣN�߂t�_=�b,��G]����K	?պ��ڏ�m����z�����v��ۈ�_�gOs�5n�Liʺ��+*���@ɨ�T���- r�7�bEY�`�#��D�&���V�;��P�3���7{����7-�XK�4�9�V�y���;��3v�:C�����@�YUT��mʖ��9�߿kb �`�`�b��UH(������ �߿��lA�lll{�_�]�<�����n�w���v�x��+ �D���d�u�8ܛ��iz����wup�1v�o�����sY�3Vۖ�k[y�~���<��������<����k��E9�߿kb �`�`�`�~�?~p�Y�2h�R浭�<��������<���N(�Db �T���`������A�A�A�A����؃� � � � �{��lA�?�"*�����2�r��Թr]f��<��������v �6667��~��A�E,lo���� �666>���6 �666?���K���Z�ɆIu���A�A�� ���� �6667���[y{��y �����؃� � � � ���fL�4@�)3Z��A����߿kb �`�`�`��~��b �`�`�`������A�lllo~���<����O��~�ܒL0�R�8T��1��Ș�0 :��2=����+K�xn�]�w!5f�4fkZ؃� � � � �߿p؃� � � � ���~�y�߿kj	� � � � �{��lA�lll{^����e�K��\�y����b"?�� � �lo������A�A�A�A��kb �`�`�`��~��b �X � � ���B��ֵ�5�ۄ�5v �6667��~��A����߿kb �b�(� %
���� ��>��A��~��A�A�A�A��~�v �6667���&\ֳ.k2ֳܰZ؃� � �
7���[y{��y����b �`�`(X ����[y���)�j̚-ѫ��kb �`�`�`��~��b �`�`�`�w��~�y�߿kb �`�`�`�}�ߵ��A�A�A�E�I{|~h�4�K��P*�$��H2��U��n;E��M�Y V�봓c<�5�)[^$s�K�Z�����A�A�A�A������A�������؃� � � � �{��mNA��������A������IsK]k3&%֮�A�������؃�������~��A��������A��ok���a/�B�:;��ںBR��j��;��37mYС&��wuXѰ=�Tۗ4��U�$���~Vt�; �wj���+I}	tDU�wU��OL�\���� M��9]�@9m���,��V�>��E2S(&����6.{W;�ָ�+��,�=�#vV谷���{��I$��x$��������4��\�?0Ξ�`�҉sU$�9nX����37j�(�ٻ�j�Ξ�`n�_�BIyB��]��Բ�%&���X�����gDDCfwuX�uX<�aԹ&�r朹�aДCή�`�����r*@F��H��w0R- �h��[�O�[�nhl�+J$_��<6�n��H%7F^�@z4(����ݵ���U���%s�\�i�sv�OB�h�c���s������6+����^���q[[�m7N�zR����Mm�c��*���<]�We�̠+癴���+��Z��,�n�Q�ց����W[9�^��'����8>�����#m]��b�2ز]eLj��]۞��\��Ӷ�K�N:���{����;���G������Í �\4�˂2x����/
Bg]g�&2�A/K���Nﯽ�Wd�K&j���>ݵ`}���%���_M �y/	x0�iƤ�yn��&����
%����U�n�U��N6�+�ā73@�v� ��f$[�M����;�
]#���O'4�:o;z�����vՇ�Q��y��zA9��f��,UUU`��`t-��������ͫВY�{�=��뭀���穄���!q�.��u�6�et��f.ɣ��θ(�@G�*@q㖀;��r���n�tK�#���.iX�s]ꈉ�[�ň$�~�IcbO�� �"B"YT�k���ZH$X�����"I D�,R1H�$�L�l���P��Q1��.��`��3��W�	6nw �lCT̒�S���ٛVz#�!)��zՁ�=�`c36�,�ǎ5$����@�-��?u�J!$�v�X���r7��&f���@>ȩ���6z� �=��٠~��\�1,XB(A���w�:�㥓eKL���dn]���J�y�����2�� �bx�&�~��-��� ��g�/$�_Ho��Vy�YSU%HK�,��@;rb �P�*@u㖿}��J!L��zBI��f��,
�� ����'���na�HH�� �{�ԋ�Jl"����CB!�H|�m�4�f��N��\;	.ka�tQ^�X��0(�ȐHQ `���D�	
+��T3`�,�0�� �D7�4��=RO&ç�@t#z�F�+	�A��0RA
-
�����!"LA�z(|�# �����v����d&8��i�� �z��'b� ��b!½D"8� !��y>q^�E6)�����D�D`!��@>Dv�A?
��g;w$�}�ٹ$�z�9�II���j�Ô$�ww�`oOs�:�k��f�k�W#1(Ҙ(��Ұ3gu��Il�t� ��<�X�}�nh���m�����1��
<w=�����e�bBe�Y�6��p���;����^�����R��BO�����>��]	z>��y���@�6����Jswd���R���ܘ��tKĨd��$�-��z�ZyB���t�wuX���R�$���73@�ڴ����١3���D�T���{�����ۚ�i��Ǎ	Šuvנ�4[w4]�@�g�ĵa�`� 7��l�U�z�myO]�ĉ������@��(����vsH�M$�=�zh��h�V���^�~�r�bQ�����h��@I�Zۓ�jL�\�*�F��F��k�h]��{l�9m��/;P&�D��F�0R-|�O{���;$T���- ۘU�RY�����z��4��h�e4.����}��1�j����m�������j ���ݦ�,Z�ŏ	�iW����=N5GYx��y���o�g�=���EhiC�S�9.n�Mna'��:٠�-*����g��3�R�.X�<�=)���g�%�Rmp���zZ�.{p�躭�㝬�-�k$n8��<4곱u��է]��K�Vb�62�:(]��lː�c��Ǐ�Q�@�����e��I�ѩ�`����<�����+`�!��zX�[�8��v94�䍎I�?s���?r�h]��9�4�׍�V2cO���,�ۓ:�;&�;D���ݒ�J��4X�vl�ٵg�Q�t�[g� �{X1������$����1 �Ih?�W2{؀;�^Ģk&$�H�����fe��_����@�s@�]v4&E�L11F�,���N6���>=�ӯ�|Ӭ�/scSU��<i���,Q�0Q��?�Z��qvנ}����~a�{����`�U��Y���ܓ��{7��`����ġT$�!D-�B��O��X?o���l����o�hF�3�#��٠|�vl�7��Ł�{��ǆ�5,������}��f;=� ���|��P�7�nՁ�;*e.�JR�e��� �- �Ɉ�M@v䘀�WU�$� ��6$�&AH�Ys����r���l�C���*��e�]{������i���nE�
�����hV����? �����4�bpiH��M@v䘀��- �ɋ�U��v�&%Y1'2F�h^�����V��Ґ.j@�X��%�!(P�B���:����`nΎ�>h��������h]��������t���ʰb��[Xnn�ۓ��?{�����f8�	IB_�BQ�"�5N��ԴR��X�2k�Ų��봜�0��Ѥ�C��B���ۡ�H�b�dȜ�����l�D/%�>������xӌ#��q[^��W|�
�������=�{s@�ﱼ�1�x�Ԏ=����������*@v䘀��T�f��<�ڑh]����hVס���>���!'j��X1����h��슐�& ;}�ܘ��~���{�]ZܹK�(r@z7%=g�w'<m�izj��rk���9���k�p��끺��_����`|�ݛnϡ%��gu��~�|�SӒh\���"�S'>������XۻW��"d��0jf-1Su-��l}�M����V�l�8����m6��b���T�zI~�BK�
+7��`��X?�f�н	)��zl~9��g�PMK���@�j�UW�<s��%�{����6�!ȩDHAH+<~���ݮ�Y(݌ lW��Mbԝ{CKo*�p�H�
�l8q=���7b�g*E�v�pFꖮ���)���*�M�h���t6ʅ�m�Z�˵�`vY�<��d�g��j����נ�:��١Jڃ��lj-�OZx��o�o��å,]$���`č��nfq�컞v�5��.˦��J\��sk���NAi6�$�V����w{ۿ�����<��r��宗J4�����ۧ�L	ԁ��r��(�������/w�c#ə���/���nL@s�*@�j��Q��xG�cƔ��]���H�}�� ��qs���䃶���'�@n� :��H�M@v�� ;nL@�-C�n�Z��Қ��a�
��oM���ٰ�IDG�)�w�V�|5����0Q�I&���נq[^��8� �Ɉ�����V�yZk����(�՟�wk_=�����]�����o󻻲-�7���cbr>W����?^�V��_�Dy(I}!�{�`ow�L���ELѣ5�f��}�zq��D�9&{~�f́�wf�"M��ֆ��
�jjhsJ�7�����l��I(M���{�ۚ\��ec���!�I4=�yB�������M��fڰ�IyB����V��zK�t)�*[���1�����ߗ���5��6��?���P{����O��%���&wd��OQSl�΂y��l������"����sʐd����1 �Ɉ��pM�Y1'0q��vپ�1 �o���}�^v�o�H�~�M`�j`�IuUVٽV�7f˅�0��HHh��D~J�;�Z��wU��wT��b�R�IUV	'���`}�֬�٠�l�;��ocx9�}!1�1����{x���L@v�����g��j���#kYٹ3����s�1�2=�r����tu��ro��d���ݮ ?Oj }sP�a�������r�K��rܦɩ����6�С�s���޵`nm_�D6f.IsN��6�Hꪬs��ۛjΏ%
Y��4���@?w���n&�FUXt$�ݽ�Xv�X}�V�J�B)"���1iȕz���k_krI����%��M�u4��ͫ�DyB���W���X�����T����F�4�L`k9^s�]����-���^�I6$���.�؛S��I4�hyl�/;w=�}��}}4_{,o��d�)&�g۵}�M��֬;z�~ͫ�Q���ѼN|fHF9&���nh76��BI��z�s���O9��6��I���4�hyl��|���٠����1��x��M ��� �&�'\T�;�>�9T��[�ؑ�$�6���B,�7���`���7Dӧ�ȍ��+������"�0X�X��
T��E� ��t���$���ՂT���c�,	 $g�.�D�e�ЛZ�˔�$b��	N�!���<oc�TH�І�0-� hkt@#�!�� F, �!���&�FI����rqipf��OJ�e����b�gwOt������p� �kzɶj��Ժgd�"m����pܧ@�7h������r�:np^�^�	�誫h#��E�;=���[���[>��8`� p�]*�QI���l��b�#H���T���XA�T�[Q��2.�ݮv�,u�V˷n«.ae�P�nP�t��h�[Y���C�D��
�"�m�q�V�kl��m�u���k�69j�]l�M졮Hd�5��{GNU��F�q9�b;tѮ�3��e5P�"�q�яm���g��N��j�[�h�Jv֡���I�� sU�Dn���U�NMgP��6�!%�/@*Re�4�y��845T* ��S�p�t�9��v��aE��#�W��hrD�mش���T��ù�D�zSI'$��]mX{[:��2�tb k<c�B,���hH���nU����E裳f��ٜ�@���`��΅�
��-�+pv�ul�^v�ϸ�d�[X�����i��6d��*P�El]tl
<�{.�பy-��c�Zn�ڗ����� ���+�F�r���u�����S��R.����m������{y^�V��`�4�8��l�b39Y�ͩ2&��r! S����� :�uɱ<���#\n��`����j�ŜtcO5<ͅnV,sV���r��8��9�>�IV�"�f�7n�d ����;;@@�;���d��X�[��KX���)P�4ڷe�v7rd�-v�F���������[Q���on�Y�=�K��݃�����+�%Ѕ���ltnnLvG�_)�C���ui�j��&.�7C�4�����X���[\0]iT�&�nZ9:sLʯ�st���*:��ˇ���TXj�pq]�ԝ�:Pνjj7%�]��=,^�Z�\���UVIʻc�s�փ0DNה�U�,��͉���\�1��6��45���97vvV�c���q� ���ƶk����p�hN|�!�� i��
#��R(�� `�PzT�v�J�}�:*����`�o˻z��`.rF��iN��أ��NR}����M(a�X�.yٻi:�pT����N�n���k��+eax%Ω��r��ק��]��Wjɒw�%��/M�oU豘,�ݍqt��E�E�=ӗ��S��]����qq ��f2&�OZL�bG�D�0�����ࣞ����TW1�
-��å.���
R�UK1B�'����Sr�������0\��9�۱�[͹�Y`c��7V�'D���f����,x�$�ݾ���j�3skС//�oz�;�!#q��i4`��v�hol�����7�3����0P1'1�� 	��@뚀sP�� 92	��S��I4?��o��__M�;)���@��ǋ�Q�)��w����/ ���ι������\���ưY�L���v�7g��vϮY�=<�ͪjZ�&WK�n���Ga�u�H�5 s�o��ﾮXK��h�6`��� �IHhm�fg~(�S��������@v�& 9� "�DϫM'�8�����l���ٽj�7����F��\Ӣ�J��wP�j�qR rMA뾹�@[|����i0rM�;w4}�����\��$�nf��³+��n�W\��p��I�-��%��6�].��L�LOsNf�v�4�3j�37k�yB�C7�j��Od�Jq�0JH�@?s�o�g���_y���� �wj��&��]LŦ*j�F��w���fڱÂ�R��!(��h9l�;��[2<N`Ȳ1ʫ�O����;���ٵa���uX�6`�K��Q	9��l��sPrj�qRvQr�W�^�V���\uu�O������*ZedFy��X�J�x�o>�dbx��M ��٠uvנ��4�٠w�U���`�R:��n��G���7�j�7��X:�r���^�]��f� u�@��g�2f�����zl�dj�&F��M�䯽����:���?��ąt��LΧ��~��<��e�
6�	Irh�vjܓ느�j�W^�׷y��5��!�sg�����q�`Dwq*̺�仝QU=�X���O�7GK��[o������qR rM@뚀�d1f�Fl
�MR����ٶ��I���?%�H�o��W��^>��&����w�H�5 s�jܓ느s���c#ćrh{���U�zl�fڰ�o{���s]6榊��*GUU`c�ٰ<�!(��{����W$�����_��,PH���x��k/rݎu�ny�Kƴ��=���ez}��;���K��#f���y���	�lv�Rs��<�I�*�P�W�y�T�tĴ����ԹJn����j�*d���]S�gI��I�=lZ��qt!lҙ��]�Ӳ�p)q���X���$�ޕ�W\;Yڥɥ���Og���n*e�V9�z��\!m��^���[��O�{��w}[q߯�8TW�ێ^\l�5���r�x��W\pTt��,�:�3�V�@ǎ4�i4`9@�����f�~�6�%�}�6<�T-�I�L��`c�ٿ(���ޫ_wM������H矒o�,#m��H��v�hn�Y���J�ǻ�`~�S R軼���ےj��� �I��sP�k�����M�;w4�& u�@I�	m�*��Kۥ:��j� >S�v��9��vŶu�,O.�ۉuc`�JH&��� ��٠�����C7�j���NH��T�Sd��n�u�]���|���>�b����,7v�Д$���܏5�54T��X^�� ��ߵν� rM@뚀��a$��T�,�j���B����ߒ ��� s� ��P㕡yw�"dmbjL��f�~�]4�٠~�6Ձ�B[�ɒ9����	�t��Y�[����֜&��?��|�%�%�k������Rqn`���' ;|����������{���l5ҭ�MMU���,{�7�	(I��޵`��`����z&N���r�S�@P�����7�f䓾����_ဃ#ȨȌ�-`� �^�~�{�3�'o{�7$����4��)���+�zh3g��͇�?�{�9�̦.b���Hq�&�~�]4��Y|���nh����s�� C� l�m�j���;�����޸�KK�i2��vR�Uv�wL3�H7*GU4X�s]���_�����%�y��[ND�,K���J��bX�'{�Y2a�d��[��j�9ı,O�}�p�C�k���b^�����Kı?g�k��bX�';���9�ʙ��{��Ir��̥˭��bX�%�����"X�%��﵄Mı,K���6��bX�'��S
�L��L��X�Ϊ��ff��ֳZֶ��bY���?kߵ�Mı,K�k߮ӑ,K���bn%�b�أ"'� MD�k��ӑ,K��i�7c��ZԸ[��&�X�%��뾻ND�,K�O�����'�,KĽ���[ND�,K��k��bX�'��Ofs4d�f�S^�h0���L�u��{P�ͧ��0�:t/.��Obs<Xn�[��������oq�ߓ�ى��%�b^w��ӑ,K��w���r&D�,O���6��bX����L����&j��S
�L��N%�{�m9ı,N罬"n%�bX��}�iȖ%�bv{�17�?�Y
�L���L�/&)�&SSUSUp���%��?���Mı,K��m9ı,N�{f&�X�%�y��[ND�&Bb���njUT�r��Q
�L��/BiQ;���~!2!2��T���%�b^w��ӑ,K�E�I�o�����L��_n��\��eֲ�,�ZѴ�Kı/o��Mı	���N+;�WL��L���T��X�%����6��bX�'L�m "|ĨȠDB�u����1v��t3Et��l]��!�nC,=͠�Z�la�&�u�s$�*HMV�ӌ�rm��� �CN�� ���	,�;j�F�n���t���Ԏ7��Bhn�U%P����][��M/i{df�oFtW�s��m�O�v�Y(1Gn^�N4�/s��ôEm�, �]��]-ʈ�R2/n�g��S[ �\�Rm�l&��j �A.M�C7.��,ɬ��P��c%=���]��m"t��.�6s��/l�u���;UO������D��ߵ��Kı;������%�bs����>��,K���U7Ļ�ow��~�l�U�MW�����bX�������%�b^w��ӑ,K��{=�7ı,K����r'찤��Z.��U�)�UC�榇
�LKĿ{ߵ��Kı;��eMı,K�����bX�%�=*n%�bX�{��̺�4I52k�sZ�r%�bX�׾�&�X�%�y��[ND�,K����7İ?ȟ{߾6��&Bd&B�S�d��PK�SS5S�X�%�y��[ND�,K����7ı,Nw���Kı/�}�Mı,K��w}Bf�%�K�jj�f�ѽP�}a��Ɛ��HQ;'(;ҍή��v��!�!�ɘS5�f���%�bX��ߵ�Mı,K���m9ı,N�{f&�X�%�~�}��"X�%�������֦�e�R]k��bX�';�p�r�BF.�P�SO�1�'"X����q,KĿwߵ��Kı;������%�b}��	�2s2�Yn[�Ѵ�Kı;=혛�bX�%������c�!�2'���aq,K��߿p�r%�bX���F�.Mn�fSZ�h��Kı/�ﵴ�Kı;������%�bs�ߦӑ,K���'���񉸖%�ow��_��s�F�5{�[�oq�X��{XD�Kİ�B?{�?M��,K����f&�X�%��u�]�"R!2$h�����*��@������	�Nw\��[Z���Kn�p`:�k#�p�v��uώ�U�*eUP幩���!2!o����9ı,ON�f&�X�%��u�]�"X�%�}��J��bX�'��r]iD�*B������L��Zf���Kı>���Kı/���C� 3�2%�b}���6��bX�B�S�a+�PT麥0���L�����ӑ,Kľ�g�Mı����
Ք�%�ɹV����Ć$MN��q��,(@��ɜ!�j�&9��v`SA���&�[O }>�	ޤ0�:��V!$!Hс�4�b#X�#PB�`@1L�$5Y�4܌B�x�b�H�V�>~���`�e%fk h֋�]���qXG��X�L���" RZ�u�b�����`�T�P��0:�D�`��GN�"=@b �/W倦 ��D�M{{�m9ı,N��f&�X�%�}��L��p�fk5v��bY�D����*n%�bX�����ND�,KӾى��%�b}�w�iȖ%�E�n��*�r�ꦇ
�L��N'~׽v��bX��?��p��Kı;�^�v��bX�'s��7�7�������۟��� �E���I`�:�p�/jz���e�������5O`])M�Y-�]�"X�%���l��Kı>����Kı/���Sq,K�����ӑ,Kľ���rh�tk2��֌Mı,K�k��NC�șĿ�f~�7ı,Ow_�]�"X�%���l��Kı;�z\�d�m��-�\ֵv��bX�%��=*n%�bX����Kı==�LMı,K�뾻ND�,K��}&��f��r��jT�Kı9�{�iȖ%�bz{^���bX�'��}v��bX)��C�ءT
�� 1
 ��9��f���	��>�s�]iD�*Bu���Kı==혛�bX�'��}v��bX�%��=*n%�bX��f�����L��\��})��,%J�$a�UI!!X�5�ɠ�xΔ��죗�&[\;=m�i&������{��2}�{��r%�bX�������%�bs��ӑ,K����17ı,K�z`xɓY-�����r%�bX�������%�bs��ӑ,K����bn%�bX����OȆUI	���QUJ�Fܦ�U(�d&Bq,O����ND�,K��ى��%�bs��ӑ,K��=�a�G�2%�b}�~��2s2�Yn�Z�r%�bX��_�*n%�bX����Kı=������%�b^w��ӑ,K��w�tܚ2�̦�u�q,K��u�]�"X�%��{��&�X�%�y��[ND�,K�����Kı=��Pъmd�4��hW����v�9���u�Z�F�O;q"��39MhF�A�9����oi���(�\��dvځʼ�]��;8�x�=v�8��m�f�U,�t
�4h[��ĽJq'tl�U��!��O^2�cTH�HIK�n�]��������ŝ(M:wV�aC����k��^��C��^�m9`�ғ���&ҝ����_b��{������h�\gj�n�P!��tnr9OD�6�E�Y03N봃���Vg9�5v��߽�7�ı>�{XD�Kı9��iȖ%�b^�{X�r&D�,O��~�NE2!2a�J�EL�P幩�²ı9�w�iȖ%�b_^�X��bX�';���9ı,K��zT܄�L��_nk��S&�IR�&i�/�,Kľ���7ı,Nw]��r%���Dɉ?{3��Ȗ%�H_mo;����L��ZJx%h*
��Mk5�Mı,�2'�߿]�"X�%�{3����%�bs��ӑ,Kľ���7ı,O���<jd�Kp��k5v��bX�%�s=*n%��L\G�{��|Bd&Bd'�z����%��뾻ND�,K��HY�˪a�uAg``m��O;�Ͱ�=-�I�Ϙ{O1;9����WS�x�S����,K��}v��bX�%������%�bs����>��,K����!Y	��	��;�6�O�.�[���S�r%�bX����&�O�mA ���1v��^��W蜉bg��ݧ"X�%��﵄Mı,K��}v��bX�'s�Ӧ�і��e&��kq,K��u�]�"X�%�}��J��bX�';���9ı,K��kq,K����s=r�٭���kWiȖ%��D��3��?J��bX�'�׿]�"X�%�}{�bn%�bX����KĤ-CЕl�����sSC�d&Bd'��}v��bX�%�﵉��%�bs��ӑ,Kľ�g�Mı,C{�_��~w�,��xq�W��h��ٻ+���6Z�]��c���N�r\���6�Γ$���r%�bX�׾�&�X�%��뾻ND�,K����7ı,Ng{��r%�bX��^�a0􆤖kF���&�X�%��뾻ND�,K��k��bX�'3��m9ı,K��kq,K��;�CƦj�.f�WiȖ%�bw=�aq,K��w�ͧ"X����j%������%�b}�w�iȖ%�`�#�g�kZ��2ᄺ�7ı,Ng{��r%�bX����Mı,K��}v��bX��=�ߵ�Mı,K���%����Z�p�˭fӑ,K����17ı,?~����>�bX�'���aq,K��w�ͧ"X���7���|!�A�u�qcΆ��k��-/��.��u�6�]���r�z�E�F�)�f�q7ı,Nw]��r%�bX��{XD�Kı9��iȖ%�bvg�q7ı,O{�.g�R�5�[���j�9ı,N罬"n%�bX����Kı;3����bX�';���9ı,OC���n�Y�֥���7ı,Nw]��r%�bX���\Mı,K��}v��bX�'s��7ı,Ot�r�E�I52k�3WiȖ%�bvg�q7ı,Nw]��r%�bX��{XD�K���P>S��� TSA���"Q`�[�������9!2!2�+�P��sNa\Kı9���ND�,K��k��bX�';���9ı,N���&�L��L��	or���*jJ�P*�k.Ůvtg�W�eKL�O$!��=,If�Cuڙ���0��5��%�bX��ߵ�Mı,K��}v��bX�'f{��$�L�bX�{߹��Kız�~5�jk�K�aq,K��u�]�"X�%�ٞ���Kı9���ND�,K��k�����H���ҁ�72�f�X����r��	���pI�N罬"n%�bX����Kı;�oN���2�̦�����Kı9���ND�,K��k��bX�';���9ı,N��s
�L��L��Y�������ә�m9ı,N罬"n%�bX����Kı;3޸��bX�';�siȖ%�bo����T��*r$6��y������*�a���^�%�8���#��JJ��s"����]����j�5˶C��Y��2�Li����tsd��.m�ܩ`�v4�����P�:���͜�Kr9�L�=[�[8�fZx�7&W�����| r�qV�k����
Y�u�u�hɊ���q4�K2jΔۢu�ۊ��yݹ�3Xl�*Jd ��vۧ����m)�����|t�N�Jݍ�0";�Tf�9/sn(��[{[p�poK1�=����7����k޻ND�,K�=뉸�%�bs��ӑ,K��{��&�X�%���}���sL52]L�3WiȖ%�bvg�q7ı,Ng��m9ı,N罬"n%�bX��]��r'쩄&B�S�a)� ɧU48VBd+��;�ٴ�Kı>��XD�K2&D�����Kı;�Ҧ�X�%��u�c�S&�[�5u��r%�g� dN�ߵ�Mı,K��߮ӑ,K���^�7ı,Ng��m9ı,_u�5�jk�K�aq,K����ӑ,K���^�7ı,Kϻ�m9ı,O���7ı,OȈ~����d�k���nʸ��7c4R�s��=;u�K�c�yTu�K��������׻����ŉ�]~�7ı,Kϻ�m9ı,O���7ı,N}���9ı,N��Ӭ��2�ֵ�k5*n%�bX��w��r�ڨ�"�@`(�B �P�bT|5�ND�9�ް���%�b}�w�iȖ%�H_c�+!2!2ef�sS,�C�ֲ�Z�r%�bX�g}�"n%�bX��]��r%��dL��]~�7ı,K�}�[ND�,K��u�E��f�T���7ı,N}���9ı,N���&�X�%�y�}��"X�E��}�"n%�bX�t�r拚a�������Kı>��\Mı,K���[ND�,K��m���%�bs�w�iȖ%�b~ �������ͭ!z�� �b� >S��:e��`�8�;���'��1��-��#u�3Z���Ȗ%�b_����r%�bX��lMı,K�k����ı[��p���L��Y��#�R�J����kiȖ%�b}�f؛�bX�'>�}v��bX�'{u�Sq,Kļ���ӑ,K��wY�5�Z�i��i���%�bs�w�iȖ%�bw�^�7�j�ފ�ך��3jC�D`��0��@�;�.k���Kı?{�m���%�bw�{n̷Z�p�ۭ]�"X�~D`dOz�����%�b_����r%�bX�{ٶ&�X�%�ϵ�]�"]�7�������.B����}���bX�ϻ��r%�bX~H�_�k��bX�'�׿]�"X�%���zT�Kı>���K��R]��Y��e�3q���=i�g���҂��m���ǟ@�M�Z%���ֳiȖ%�b}������%�bs�w�iȖ%�bw�^�7ı,Ng��m9ı,N��׍Yk��f����7ı,N}���9�,r&D�=�Ҧ�X�%��w߳iȖ%�b}�������ʙ��~�˚.i��Mc���ND�,K޺�*n%�bX�ϻ��r%�bX�g��"n%�bX��]��r%�bX�L�Sa)� ɧU48VBd&Bd/��}�ND�,K����Mı,K�k��ND�,
l'p�F�(�"�XBF @��"e �A%4��D�߽*n%�bX����|jdіf�k6��bX�'��k��bX�'>�}v��bX�'{u�Sq,K��}�fӑ,K��=�����NWx2���A�s�zp=�Im�	iA���vR�Upu�,���3�7ı,N}���9ı,O�{�q,K��}�f��'�2%�b{=�(�d&Bd&B�����U6�1��]�"X�%��+;5����Kı>���m9ı,N�}�"n%�bX��]��r'��L�bw��蚺���tkZ��֮&�X�%��w߳iȖ%�bw;�aq,��2%�����"X�%�ٞ�q7ı,N����˩��։3W.��ND�,�02'u���&�X�%�~�kiȖ%�b}3����bX�L������r%�bX�����j�a��f����7ı,K߻�m9ı,O�w�q,K���]�"X�%��w��&�X�%��� 8|g7�
�Q�:� �|.ӂ�@����7�t���Q4��:aݎ�lB�lD�w��H�#�"�j=80$R�#��<*?q�"�6M1P�� ���X�Q|.E48	����
G�x��9��P����.�t�`顀�c��Ґ
�	!|����? Sz��l0�JGb�t���!� w���}� �N��"�ڮ���	���A�M��+u��-��c�N	��dRu.��٨�j�MK�,�`$�Ab������v��v�p�5�����'bf��"jgEX�[v�$���:�48�w��r-�5!A�×m��9Y��W"
��U�6eq����=�m������O�y�򝸮�#���
U�tmNl��ciMѳ�C��ł�cs��l�&#J=9���CQ4���fɸ�;u��U�`'�n�;�n�R��v;�ےAe:�׵em��)KY(`e�l�(sUl�� b��c���,'Hd\�r���/[����#,$U�v���m]\2et�Xs�TlE,I�ʮ#�4
9c�p�N�]�eń�݄q��n��z��[j�k��.��Έ�v�:���X(I��s+'3l	jL&qьpZA2�WS�]���TM�	��Sni;81���4j�l���a��3�|\�5]�և6�UИv�[����e[vSF]����2��J[-F��Х�લ���
^�-�tuZx��R�DS��F�|��k[�jNѽ���v�El�j��6W���C	l���y؛� �]�!��̮�4U�m���3A*�q�m�ؕn�_n�]��o;-/g���[C�#58�,��A��5gc�M�	�]��l\nNݭ��'X찜Ɠ�Kg,�ղ�G�v��[uU��d ;`��-�1���9uR��B�N�5N�焋g�:!��e#���ݭ�V�����r���|T����dc]"��E݃FKTqV8.��4��6�1eۗ[3��F�dFl�Nm�:��ِި�M��n�A�l�ԁ��$���ڬ����I�W#����N�e%#Z8�Q�'i��"]n��[i9��3�њ[Sdű�;�l#,�h�\j8l�Ywn�z�[m�g'���M!�lrn5��R�Ú�U�asv��������iA�xT�	��N�� �(tt�#�E��AT�DJ*?z(��A�U���1��t~~�6�^=�TuV��x��I%�M�Lu���ΊL뛳�<�ap�
�t��u��m�k��;X���;L��gF#�^8�g2�t�"��8[��+1��������O7*gPr*�`˧�X�&���ڳ@��e��]S&��ַ-j�8��z�7K�BN;&ʗfx!�&�3�M�b�tg��D몥�z&G��}%kv�`v���:q���ϻ����9�i4��^���9.;r<�u��{P��k��i.Ν��y ��t7��t��~����%�ٝ���Kı9�wٴ�Kı>��X@�T�F�Q,K���_�L��L���6�$<
�eUVkWq,K��}�fӑ,K��;�aq,Kļ���ӑ,K��g�q7�)�2%�����j��K����r%�bX��~�7ı,Kϻ�m9���Dȝ��鉸�%�b}����r%�bX�C���kWF��rL��aq,Kļ���ӑ,K��w^���bX�'3��6��bXE?���߿k��bX�'���a��]k-���k[ND�,K��zbn%�bX��]���}ı,N�k��bX�%������bX������~o���\א��������[�eN�,�GK�����E�N��������*���UUJ�sD����L��Y;ޛ��%�bX�g}�"n%�bX��w��y���L���
�L��L����%��5�0����oq�������7�|�L���K�׹v��bX�'gu鉸�%�bs>�iȟ�TȖ/���h�ֵsT��k��bX�%�����"X�%���17ı,Ng��m9ı,O���7ı,O�w�9�Mf�][5����ӑ,K��w^���bX�'3��6��bX�'��k��bX�&��ޫ����L��XO�	O��5�kZ���Kı9�wٴ�Kİ�40�w���'�,KĿwߵ��Kı>�צ&�X�%��_����{���É�$�j�FѽP�}vۋ��Y7F�G��;�����>�}�s�����k>Nı,K���XD�Kı/>ﵴ�Kı>�צ��DȖ%��w߳iȖ%�bt��W��tj�$ɬ�7ı,Kϻ�m9ı,O�u鉸�%�bs>�iȖ%�b}��������2%���~��g2٭[p��kFӑ,K����LMı,K��}�ND���ڈR�o�tv�O�s>�����%�b{���"�oq������
�U<�g���X�*�"}���m9ı,N�k��bX�'>�m9ı,O�kI�d&Bd&B�2�ItKM� �su��r%�bX����D�Kı9�}�iȖ%�b}=�LMı,K��}�ND�,K�ޒ�!Lɺ�̜:^�cCȧ�t��Xr�zY�%�9Ѧ�]rOjOI8v�]kZ��e˚�q,K�����"X�%����17ı,Ng��m9ı,K��Z"n%�bX�t�s4k4��٬r�Fӑ,K��{^�����L�b}����r%�bX����7ı,N}�p�r%�bX�IO���T*����VBd&Bd/��}�ND�,K��ֈ��c��Dȗ������bX�'g�~���bX�'s޹=,�C4asW5�ND�,K��ֈ��bX�'>�m9ı,O��鉸�%���'����w�{6��bX�'{HXk=��\-�k5�&�X�%�ϻ�ND�,K��zbn%�bX�ϻ��r%�bX����D�Kı/;,�ِ��v4@8Ei�n),��p�^��&Jn˽&��X��!��l�!��U�{�[�ou�b}=�LMı,K��}�ND�,K��ֈ��bX�'>�m9Ǎ�7���?.`�!uS�6}�oq�X�'3��6���9"X����7ı,O���6��bX�'�����WD�RBd,ݾ�]өmR	�.�n"X�%�}���q,K�����"X�%����*n%�bX�ϻ��r%�bX�}�%u�j橗.kDMı,K�w�6��bX�'޺����%�bs>�iȖ%��Y�3���"��	��Vw�UM@��T�Tm9ı,O�u�Sq,K��}�fӑ,KĽﵢ&�X�%�ϻ�ND�,K`H+���'�t������]sh���펇���=F:����#��PN.��ӻ�UXy{��3��3��U,�5Ӯ�#��;��6�G]�l!��y�vc���q!b�ս]\�i��$l��ڝZŝ�dX��qkK�hU�Od���o�����Q���vz��Nז�ri��G��yڣ�VC�]��cJu�M�U���qJ��#Ai�M�����6���˱� �-�M��cd��[�	��Az�W���)W-�� ��7[cTՏw�{��7���g}�6��bX�%�}�7ı,Kϻ�m9ı,O�u�Sq,K��z{/���f�H[����r%�bX����D�Kı/>ﵴ�Kı>�ץMı,K��}�ND�L��!f��z�R�X�����ı,K�}�[ND�,K�]zT�Kı9�wٴ�Kı/{�h���%�b^w��̚�Y�[p�kZ6��bX�'޺����%�uS���ͧ�Tș�2&g}�����2&eO��6���{��S��r�~[����-<i�bn&eL��S���ͧ�Tș�2&g}�����2&eO��6�}S"fTȝ��K����2&eO£�}d�5_�Ξݥ��o=y��N�pmڍ�"ݬ��]�WI����	���ځ����2�D���h�M�̩�3*s���i��2&eL�ٚ���Ț�L��S��߮��dLʙ����+�kW5L�sZ5Sq3*dLʟ}�|m>���iJP"�
؊��G����=3_K����2&eN}�z�>��D̩�3=�h�M�̩�3*}Ӿ���5�aul�9u�i��2&eL�������S"fT�����d֪j&g��Ѫ���S"fT��������r��{�5��2c�u�)����fTș�9�����2�D����U72�D̩ϻ�Tș�2'�k��n&eL��S=�e��S!��!nMf���dLʙ3�֍T�Lʙ2�>�6�}S"fTȞ��K����2&eN}���>��D̩�3��v7ݭs��b���cv�w;��v��Kv��TuϘ{O1)=Ƴۍ�Y�vl3I���2&eN}�|m>��D̩�=3^�q3*dLʜ���m>��D̩�s=�3I���2%ʙ��ոf�l֭�[5�O���3*dOj�y172�D̩Ϸ�]�>��3*d�{�n&eL��S�w�O���3*dL��[h+��Zx���}��{��S����i��2&eL���a�M�̭C�� дS�P��]
�P�@`�-Q)؝�O~��O���3*dO�?l����S"fT����՚�]f]I&�s5��}�L��S ��fi72�D̩ϻ�Tș�2'r�fbn&eL��S���ͧ�Tș�2-s�4Lu�j�.e���Lʙ2�>�6�}S"fTȝ��q3*dLʜ���m>��D̩�o}�4���S"f�������Ӯ��5����kWHF=�s��v�͖�95��m��N�v[��i�lA�˭O���3*dN��ˉ���2&eNk��6�}S"fT�7�ٚM�̩�3*s���i��2&eL���g��2˫I.kY�h����S"fT��i�ԨG"dK��Q,K����� X6%���ʚ����MD̪����Ƥ��.i�M���
HS.����4���L����r�{��˻m��v�ߒK��b2;�1&܎cԗ�����~��-����˻m�ϻ��-�l@c"	S�D5���ݶ������"D�'�L��$�]�Z�K��k��$��kǩ$�s��~��\�)�h	��<�^ƇΆ�r����7;!:�3�Y6Y�]���smz�r��W ����_���l���}��z!/���t��m���m/�d �7#��$��+ũ$������I.YbԒ_�-�$�q|�Ƀ�I�jG�RIs�����\�ŢI~|����]]��RK���l�s Q"<b�z���������@vc����H.V�Т2a�̎C@��k�9_}��'�w�7$��צ�N�1�B+�}}/�[����K�����uڳQ��cv�����pm��WU44=]-��=[V�M��H��˹�Ḱ�*����`�$����X�F�'V|@���6<]m��;Q��x�3����s����F�dy��|�u���	.�N�q���7��>��aɠ.�C�n����L�^� 6yڷn�ˋ��#<��ɬ�d�tNɒGg�`���{��pQ
 ���Sv�.����Md԰��`�`	��شqҖ���Md�zX���<������i������9�����$���wM��P��z�R��R�oP느�%�9}�뗫�T�a��Dʚ�ʦܰuT���v����Т!�syՁ��j���4)�UDLnG�)��rנ�j�9۹�r�V��v�Cik $M���r����\�=�@r�& %� �v����u���M!���9�Pw�V��t��⊳Ϸ��u��P�-1}������R�$�/�b }r��N`�M�$�V�a��F��=뺁�1H�1�A6��?.�����7$���9۹�qr�P�IDd��$�@r�& �/Q�类۞T����@�!��i�.i�M�D%�S;���O~T��f��였�p*ʙ4lLdjE4s�s@��)�~\��ۚ���DwwD��2��*t�D�x�p����x9���t<�Ϯ2]gc�yTu�T��O�������ȑ"I�RL�����?.Z���M �;f��w���1�
8 9}�c���sP��/}���}���d �7#���M �;f���N��;iD��nυ5�$���h�G0���h�|s����Y�'��!$1>/7�
|b�B��@1R��]&� ؃f�H�g*b&�d�	��+lF�!�J+*`����X��*Zj����ݚ1ME&h¦��02ѩ|��� Õ�����K+kҸe!!5͒d�?
҄(J��A�
B�(2��
c0E>"��q�?mQ�`mG�=A�!��� >`y"'��64 >U�.*W�{�צ䜾���:S���A/��8��S@�o�4�-���^���%�_)�v�3d#�q�3ݤ�ɨ_d�����qR���~ov�u;�/^���x��k��k/'X�	�;�GK˧pq�1����;7u�똀r�θ��U~����?ޟƀ_���1�O4�q�oj�u�HG�@r�� 8�ʙ4�i�l�H���v�h��Z{�K������7�3>ă��|�9$I4H�?(P�O��`c����V�MZ��������7$ﳿ����S)MUJ)�;盳`r�脧��u�	�ߵɎZ���)f֘nV�x�Sc�-��h��=i�e�w�?�	��;SU۞�S�SP�Q�� __)��@�_j�8�k�;�)nH%��'7U4��>�ڿ��_�d�Oy��ޛ ��S�>�1#���!��BcQ�@w�=hۓ�����\�o�tТ2a��NE����|���M�;w4�����h���Ƴo7�^�9� 91�@r�� ��U�� ,=���g$���uk��ĕӷ��w'<{]#�Bu�9i��LY�و�ݎ���V�Zx��bqy٭��!4;	��+�D�+t$5�B�v��Fy퇙	���t���"�Zx�5�&�s;Y��ͧ^
G�B��Z9P�����7Z1���b�zsmC�ֵigp�5g�.\�.FUn�W��eJ��h%�x.v��n��{�_��� �NW{z�O3$��;��=�pE�<�H3an�Vs]61܃Ƙ&�Ԋt�]��}�@������M ����x�H�$Ѕ��Lr�����/P���w���L����@������M��k�?Wڴt���-Ɣ)MT�B����u`|�zl�9��������� ��H�X܎)�~\�z&9h_\� 㗨�ʵ�f�TZϯZ�q��]��+����{P��k��k]��e�q�B9�Ȅ�MǠ~��h�ٳ`���DD(��>��V>�<e�WT����w$�����Ck�`�}߫~@jr� 䊐����� �x���@;{T�?s�s@�_j�?.v��^	ev������9� 91�@r�� �@q�'�bD�&�JI���V��s��w5Ձ���]�0s�|:R�J���Lv�.6]��jN�,�F�����]��W���H�b�)�HȤZo��v���q͂��9Ff��@�ݽʩ���W�
>ޮ,�w����ٿ}��{$�I���4_OI�g}w:T~b�P `�+���XJU�/AM��-����'?_)�s��[&G0#��ϗ=/� �Ob q��� ;q�@��)19���נ��h�e4�����]Y䏆5�c�M�$Yg+�h�}�\����띝Փp�9Aޔg0E��Qō8��/���9����}�@��k�/,�,n�Ȝ�nE4�͵|�g�;����t�nk��>���x�$H�h�I3@���?.Z��ؑ}|���?yh�ki�(�����E��v������Z���B��V�W�9���Y���ږ��osw�^�92K@rc��v��x�$�d�2I�k#�ō�	�(�ڷ>����ݍɰk��ֹm�&:��Ճ�C������z����1 8������ɒd�1C#qh��ZW{^�v���~�ՠq^㠆%��Nj���3f�3s]Y�����s�Z8�SH�#�q8���D{6Lr�{�x��@w��2�3Вn7"�9e4g�������;{��nI;�����G�E�D"�@;�j�RMj]�0�BK�P�H���Rd$�@�
�ݧP���WI��K����ݫL�<�c�,hʄ�����k�,`yF��(ε�M�9a{gK'e]���JneB�cg��R;��nڪ3�4��4�MU�A�Z5ӑ�s�x�l/0�����6+bq�c��a��NE��[F�K�ө�+f�YʣEJN8rV�k�u��5Ɨ��Kϻ��{ާd��� �����Ol<�IЦ��Sl���c\�G��@K�h��{���Q';����Q�~A޿yh��k��Jbr2G����$�6˺���vn֗�%�{����J ��9�v�@��1 �� �1 � �mm�n�ۋ��8�Zm��8�k�ܶh�n&�L�&(��r-��h\��m�@��@�ꦧ���{���I�]D�m�k��[jyHAz�S� �(��QĜ���1I�8h\��m�@��@���SHf�������'}�k[��H?&}���Z9e4.Z�ى��c�H8���@�_���)�qrנ��@?w�|�9$C`��@������vls6�:��]��3���"	LNL�C@��@/{f��;V�ye4fw�a�����y���6��^{�nr�gu<{V��k ׷d��`�i采���D)r?���@��@���? ��P��v�_I"qcm94[w�>=b��1 F�e\���d�2<c�h�S@��Ng�,� 1Q�����
D� !(���DDѷ�V�������h�X�Ĝ4.Z���h};�á>ξ,|3��+���&����mX�����Ł��vtھ��Z�h�&�I$�Jd3֗y�v8�KtGQg���y�e�ŗ�sQVm�qG&��;V�ye4.Z���h����� �MN-��h\���l�9�j�}�o��DqJbrd�-�����٠s�ՠ^;V�y��6ŸҀ%"�G���@�����{���䁃��S`�S�q�=�,��	}$#�iɠqrנ^;V���^�^���jK%Ȟ<�7(u��n/U�`�{v�=�ݳV!93���ٸ�ge���W\A�yJ~�~~����ۛV��\�~`}��`c�S��h�X���Z�v� ������ڴʈ�1����9475�였��- w�j9�ee�I�rh\���ՠ�@/{f�~�j�<r,R4�8�ܒ�{&���o�b�}_V�pK�����%-��}�ys� �	���C\��!�~���Bb�u�6�C��g �0BQ��H:���)�#  �i򣋧�6�o�8�1��P:|�$�vp�����	�i|?��!��!`���&��B�!S*~<��:D� �rk���ð�;��O;�Q6
$ 0b0�@`A���1U�� n)����m1D5	e��@���"��> uZ){ňd�*�v~O�b�[�����h��bBk��81B!@����B�ۡwUUUTUG@D�M� �$���:�v7n���4P��ox�*T
�\��̧�rP���5*�)���V�9Ls�������,�s�k��Q�n��\�ܙ����b���f 黵�qZG�!��qdX�e��htWCbU���
�Y������7Ex�<�eq���]=�)�ۘNG�o��^�W��m�9��T�f� v�8\)Q��J��8��&�p�s�2\�1 ����Bn��,��⭧jN��	j=m�����f�m2�4jUI�v�%��y9m;e�[c�u)�G[n�6�cv9ŕ��d�tS���?[���m�v�X�Z��x��玬��/Wk�ۙ�U�Nv9G';:UE9*A�����N�n�nmY��9^��6�6��Ճ��ˌ	�̛��	ae͹�&�E6h.� �-���ڝUҜl��;mUW f��n�m�anm�8�Lڦۧk�.��<�Np��r��.���ӭSr��%�ڕ�R[�����n����pj�j�ٝk�ZqJ���,��K�c��d��)gI��:Z�!�tV�f�66�m�&�s�1�m�.�����n�"W��s��Ѵ���f!۲�e�@���Zj<9H�EU@ka�]k{a��Aj����yCus1li�p%^K,iX��J�$-k�Q��)��r��;��sv�M�֭�N*�j�ڋ&M����ER=��o����������H�+@u�n���R��Z��r:�ќcG-P�Ch�1vB�ԙ��떝�Y��Ź�������R;WH�����ܿm���d��ݚT
��E-uz;rk���P�z�a6-�u6PlF=2�@\pD�S�g�R�=�����ik����U���涎krcT�xL���v��a����+�ҕ�C��`�cZ͹���
�Fݳ�Iy�i�j�'�������k�I{v�<t�	*��{0l�D�'���DD��/𢏐Q�`��
�yW��]��iLP6 �U�y���_;G��`�q��Y������0�ec�9Ҧ��u��;���as�#���E�7i؜�*�im�z9w��Ut���&����jdӻki�C��kv{���q�,(��9N#�ԓ!���D�u͛�E6q	�;����5j���JPM��,N�KE���9dx��	H�I�j��v�0i���UP���O7���]��=�p �{Vݍ���C�gfw;����c�]��e�
��F�5ৱ��`F�Q��o�����nj��1ɒZv��3.�f(RF��������ڴ��o��gؑqg�����<m�&���؀��-&Ih75;%^Z�&L�Lxڑ��ՠZ�Z{�4
��@���A��1I���	2K@��	rL@N䖀��]~w|
>���N���t힠	ָؘ�,�By7Y��bV�6�1���x�l��	rL@N䖀�$�m�eK"r'�B94
��W�|��}��1�~��$I�2<��PM��vt� �ͫ�P�Ca���$f)O	Ǡs��Z�ՠ�l���hs����MǎH�9BP��]��;w��33jÓ��`s�}�m-�2`���- ������ڴ�ڴ˖�
H�2bf��@A��Д�n1͇<[�z��;,ik�z�*=!9�"2HG6ӓ@;�٠^;]��gu�DBK��z���2��R�2�R�ʚ�~��|�l����n�X�f��J39>)e��'N���`}���s6���J�KRQp����6}=��3�f-%Ԧ��/wm F�9m�@N䖀��- p��dM��l�rh�{^��Ϣ(K���׽�`��`fl=�r�x��NS�퇶m�*�s��س��睌�Y��UnU��y(��[�A�~�~~�ʴ�����hVנ�kBȔ�MǎH������hVנw�ՠ�v���ɂRdn= ���nI�	ܒ�c��up+kl�!x�NM*��=�~��^ٲLE|cI]�D7�]ﵹ'{�.�&O�J!���@�v� ��{�4�Z�[Cbf�$J}>�X�ݯ=dM�t�l��^δ��@��],O.��֞-���#nG���@?w�h\���{^�t��ܢQ�ōH����U}��d��b�'� v9��g]�b`�!�W-z��ק�I�;z��ޫ��4L�5-:�o*��w�� �5 q���\���"SI7�G��l�ٛV��ٰ?<͛�DbJ J$�ݻ��ߣ���k�Q�G�.�Z���� 8�
co8�P�������d���4a{I�a�Q���ks�7m�l[p\��M��[MRi���׮ ۓAö˵n��I��ՙ�v�ϱ.�'Y�&�%r�b)4̇5����1{WZ6��0jm�����TId6q��V�q�[m]��&�R��k�.ƨi{'k\!s���BRڔs��O��{���wn�w�}q�:ܗn\Yq�ss�����-��O.�_��iAn��6�]��5��<Nc`�ww�����;}s�%�vM@;*I�$#�iɠqs�����yh;�M ���#��[$�>�Vnn�<�޴ ۚ�#sP$���ۗ�%�X�1��w��@/sj�?f�XtBP�>��v�����(�bƤNM ������ڴ���\1<x�F6�Ʊ��M��T�9�=vrv�w]��nj�Aޔ��t��ax�i���8��-����@��4˽�j7�F��)$�?.�bt���O�� �sPrj�d�{jbȔ�NG �z��4�{f�����8���÷أ0�����@nj�d�-���ɠT��dFI���rh\�����I�����75�V����D�k׭c#�-���z�+�O��]1�]���뗱3p�W^ ��
~�~���f�>�ڰٛ\�~a�;��(��6}��|�Ĵ��#nG������W-z��נ�b�Q(�bƔ��ܒs���$����� AG|:"F.�$u#8F�}��o���v�����O#�#4��@v䘀�1 7&���W}�۠yv�D�y"I���˽�@��@?w�hVנ��wlO&D��=� �j|�P�rm��W���q��k����wmLY��I���@��@?w�hV�����8���t����c"�U3S`�m_$ُ��������k�.,��2#$�q�crhV�@r㘀v�� ��9�*����l:n�(n�l:J���`k������O��Aŵ�d)�HB1��O��o�;��s���Y���.]e�� �1 q��ܓ�� =�;��㿸�r8d���esmj_g�^�nݣ�6u�q����9�1�.�m����� vOj�$�-��nL@
g]�y	�NM���˽�@��@?w�hw�M<�$���w�� �1 q��ܓV��Ȕ�NG �zWmz��ڰ>{�6	(�O����x	�H��U3S`�6�P�'���<���;{�f�~~	�
ຽ�gu�����Y��g���66vn�W+<����+k(����
 ��#vm�Y���8�;\8���N�Xtj���mK����U��l<\�3�tr�v�����q��O2��E%�y�x캬Ɇ8�tu�y�N�u�u۴�lr��$�ͨ��t�t'N��qgK/F���a�tg���]uT��Ĝ�<d�u���N�1�&�����|	���܆�������W�9:�{	c+�G������:]�۱�6%�]�������f���\����m/���_\��&9`u�j�x̵�>Q(��R=��k�:�k������K�LJbq7#�;nL@nj�$�-�������S�cJG��徚W��~]�z��U�y�����l�`H�rh�& 9m�@�j �sPW#��g�n�	�\���=k�w�,�SZJf��I0�8rN�t�x���۶��y�h�y�v�� ;RL,Yu4ۚ��D�M���k���Il|�$�BI�Q��ofU����?<͛�&ð��(��%"RE���@��@����Wڴ��Й�cM�Ӛ�w�1�nb��@nj���L�(�Cƛ���{^���}�? r�M�����F��i�CU�-���n{8�'<;�ζvR��c/J��$�������M ��٠|�vyB���=ޛ �`6�� ��˼�� q��ܓ�� ;1Š��.��&�iɠurנ~��s��0�I\�J� ���>��"=\�|���� !;��v�	Q�$		�)hx��aY0A�R	;�\,	� ��!�H���h~G��P4.�	�y�K�M��I�!Dw5��<�X�BR � �$mD�,"1
1D��V�*V�`	wQfC�6�y"�6�D��qx�G�~��']���YN��-�"
��.�H�"���a�H	�44tW$�<��t�`P��w��g���6�LC\5� ��I��8��h�>.y
q@= P�t
x8���^*iЇA|��"�҂r �Q���J���hG�` �꘸�� �Y�������;���hW�HDdc�$�D�z��נ}����fՇ%	=���H˗I�'$�	#�9_j���W-z��נs3�f<1��bY>#h1�r��z�n�8�� 5y�+EՊ5�[eq �n���v�3j������f�D(�����-غ��ș�cM�ӓ@w�1�nb����U��Y�ɑD�	H�+|�Wڴ�{f���^�~���LY�LjG`}����f�(��^wM��Q��'�J��LA[��hG�����zl�`6�� �
\�4��d��Ɉ[s��8��+.�Xhg��dì]l������v;C������7i�%���;��Wl�25���~�6l�3f��g5�DD~`}��`|����%I5M�N��M���l�(�	&���- 徚W-z)n6�)�(������r���w�1�nb ���b�,�R%$Z��.[�U�y��{^���V�qpK��dFIYy��y��w�1�nb������*�D$$ҞӃ�M�j����-l�)�v�i��/%u��m��8������.���b��ѧ`��LVbzv�f�����q��}<�|���qWk��6�θr�y���:҇A�4k��⻁pr�'�4%�0��tXw6����K<I����M�:�D��휳�קu��6"�m;���sq�5���+l��r�v�l�\�=cR�[�k1w��b�E��}�jkZ�a3&Y��5��Ėv�v;<��T��]�A���K�14�ܙ�"!����q����W�v�3k�/�5�t�����Jt�5Y�Y�����- q��}���_%�}��l��!S����}�ڀw�1�nb��.Q�ۙ��G�4��:�k�?.����� ��٠~���H�'�����{1َZ �sP�& ;�W{Ww,�#ڷně���c�����w`���� e�
��F5i��As��~�~�����L@rۘ�%u�/0����7UN�?fm]��!@�!('E|�� 6��M���7$�����9_j�..	u�L��1��iɠ;였�1َZ �sP�s,Ȍ�nG�~]�z+�Z���`c�vl$���Ca)Ӥ�sNf�8�OZ �sP�& 9m�@z�������;<�~�GӢ㋭nc��H��v�+#�W-�pn�ť�[�x��8z�����; vOj�d�-���r���X�$�8��rh\���{^���k�ٛW��J���6��M:�`~y�6��(I\BKR��M��G �N���nI�s߮�9j��Ԧ8�r7�r=�ڴ�{f�k�Z�ՠ�\�&�Y�7UN�?fmX��uo?�}����ʴ��a`��ɉ�X�`,���{��x��JMs�����QTY�{5���m�&�k�Z�V�k�Z����:�N̈Ƒ��$Z�V�&9h��@I�Z �(.̫�ں�ͻ��@I�Z �sPc����V��p@�.S�dL�- �{f��g}w$�s޻��	Ce)t5��C��
�w�g�]�;�=$���$��mɠZ�V���}�ܳ�_�����6�����k�S�6��BI���:�s"�s��س��� �Y��U�F�M�� ��Q$�N9�9]��-}�@?w�{�y�-���1j�����6����75&9h<�ת���H.w��M
4�	H��hm��-��g$��g�����_D�e*t�R�fe�U�(Q	C��`}���ٵh;�4s�����F1dC���<��d��:���%�;+����?1d�n��i�n'�UԆwjlZ��V¢���UU������6V7)�u^&Nci�+�Ŵ��@kv��Ke\WZ!ѯn9�BZ���7u7�ё��2v���/���grir����}��k���6�[*9�,fW^p0�GC�i�S��no:2NI�`��
���z��5�y�c��Ƕ�\�rz ̗Y��0ɩsO�A6/��Ep_]�{�������p뵵]mְN��Yr�%�z�/gD�b\c��������b�m���&,��m�����Z����j�?d���`�l��!S����f女k�h��Z�ՠw�����LQ�ۓ@�ڴ�v��j�w�h�
���Q$�N9���ՠZ�Z����j�9ΪЅ�"6�F�Z�ՠ�l�-v��N�9BP���G�75LȦS�S�����ۘ|b�˔��������9�b]��n��id�(������k�h��Z�ՠ\��Ҭ�XF�m�&���޻�:���R"?��)�W���l 7�����'����@9�٠s�U��DcH�q7�ǒZ\�[���$��NX4��ФZVנ�l�-v��]�@?$�����G�njL��y%�%�1����[� nYDw+��M"c�r��}dݒ�nj�Aޔ������q3eZ�m����ǒZ\�[���C)뉨�'�@��j�*�� �{f�k�h�UhB��K#N-�{ٹ$����<:*��򈅤�
H���vl�; Y�Q3#�DC�'�s��@�ڴ�v��k�.p�iVL��m�����@q䖀�$���?}U��rװ��@�q�ֱ�U����;��9�ƴ�]1�]�:a�/bf45���=��f{ր�$���$�-:S�L_b`�ZV׹�g��l�-v��]�@?$�����G�njL��߫뾼��䘀���U8�Gӓ@�ڴ�v�$�����>��BB�X��b`
 ��S�Q�����@�<{��bI��r-�]�@�$���$�-��n�z���I`�l�]%����D��W��Z:��a��N�Ԅ��!i\t�~�������`:���%�8�K@�J�fa{AL�t��>�ھJM�����{��U��8v5[S&(��m���,�-޽�\�;&�8ܱ^n�1H�2U9�v�(O3o��wM�~�@�ڴ�;L4i1}��qh[^���r����� �>uh�*����*����
��������UU��UTW�UQ_��UQ_�T?�Q��E b �T� DP �@��E ` T�+@*�� b@@@� `�E `�E `!P*�E `��DB* �UU����+�����UTV����UQ_�UE�UU�qUTW�UQ_�UEЪ�+�+���e5�Isp	��� �s2}p�� }  �    
     h          ��T��P�Q J�T�D@ 
 �T�@" J�U%(�U$�R�  ���*� ��*�X    2� � �@ Pah�yK�ž�t�k����z������S�ס�g���}7�> |����l�y�x  �^[ٽ���p �+;N˾���ew�*�o&��� Ω˻ͻ[�ז��^��px |�� (�  PZ
w��q�'��S������w��<ʖ[֏����8�� _{�  �p�  ��-}<��  o]�ҽna�` ��[׮�]/m9ht��y� ��}�}�N^��ɪ�nMS� |��   P�@@����6�iq�Z��r��m�{�(m������{�O'^f�����������ӓݗ�wK� o]���nOR�{�Z{��\�^�z.;�^m�ެ�� �'&�p��u�xN^��� {�     E ��30V[���s�9;�p �,g�^�Mzӓ׀8� h�Z'G���)�14h �1�4H�/@� ��
�GM" �M�  1AJD

D ��
D   Z      0�i���=�) �PQ�i� �AHJ����E��p �{�VN���  ޻�s���[�  ��ݔ�;��W���T����X�l�&�׼Ν�ޕ^ ��*m誕  �'���@ 4 ���R�F   ��T�iE"b B)����R��  ))F��i���S������������������������ |?�P p EO��� � *��  �@T�?�������)�L@�L0!W!T�cV@����!�F�h����SO�	��ƲN��D`8,��hK��y��ɾ!�ϷYo�o����2�M0&a�4X�aV�MB�
@��5���\�I˯7]�@����ɴ�f�283�|4�,J(�4�G8�K���|i���5������6>�a�2����B\��AM���'��ٹ7d���ǽ��>%���70��u�fB�
@����
��f��כ�!Y3[�{�� �;^}�S$H�1"��������IB�w:~L�Xٝar,H!�X2H��U�G	o�!M:aFS[aB1�t2��)�V$�0�(A�!���i�"R\���>1��.�,���6SW�#�pC���#F#X#(@!�H�@�P�D"`�L&|q]�D���)Bq#X�� a���s[&�[�a��������׺�0bC�!
�p�C�	��d(��BiA�����VK"2,#J���}��ㄅ��h��dH����L��,J^������������g�I�>~���|(�w�ú���X�X�D��3Zeь�)>��gn���ߡ�,����|��D �bD"Yv�I���Ǝ�k8�$�`B^���n5�/7�@$7��u�7��R����$�3_o4����caRd�č1!p��d.��*K��-(F�t6�KRtԎ����g�>aIqٺh���n��:��%��,*ŊV$�ۨCpdH�#@�PL�b4�F A�bԉb@�L	X�0�t@f騁���7OY~9���`E""�aH0����fE2#as	�o��ѩM`t&�����ه8ˬ�IM�۲S6i�0!VA�������é���bҌd����J�A ��#��@bHm��Cӛ��Zt"P���B2)CH��İ)B8b|���Ս`�H$0��Sa�A�kP���|�t.F��kZ�t$��k4�BKa,&�@�H�H���cJ��	5@�˛��I�.�r淽�>8��˾$a�8K���
�a�ayL�$�nD�&���|r�E���d���z)�����L�U�@��ݶ{Y��$왪ph�œF��oL8Ӧ�O��='FO��,F,�BF$BK����0`�2c,�@�$�dHD� �Yl�!`��1	J��"�+0`Ă��	0��Y��!$�7�HY3Z�}�/~�N.�;�i's[5���B��t!M�tN���s|��A��榓`�sP���kH�� c��a��������I�We�N����	2�d	&2���ۍ�fl�S�z0"B��$+(A�J;M) H��u�=��������0�@��)�l�%�]���	��O*VQw�T����l�B�-�m7�لfkZ��
�hHH���`R�B���wjv.c�SLN���#G!L!LaI��LbBHOX)��4qHX�k{!!]��Z^�ԀP�@l�/ba�oℭd �e��5-��	p�K�M�g+�� 5�nLd9,�$�����&w����dZ�$M����Qp
b@��Q�@�n:X�XLA�iu$B�huC9�, i*b�j�,)�@(b�H:;yxL���G5�Xe.�k n\��S�vl2���V P j�/FS)e���n��L����{�WF�hA����"5�DH����oW�)ܤ琅}��s!�a��V�s4���p��s5��R���.1`D"R\����ğI��{M�$}����`j7o�MkQ�m��A H$��L8M{3݃�T��cR!A�\*>���c�_���Q����X��VB���D�C3��i�j�
4ω�Ca�L6��$3)BN�A�u��4}����X�!p�@��4,`�?,XG�ȓ
�)�H:�A� ��rvϐ뽐���s�!B0t��F��
(�Ó�)v�[6l��r���ӧ�*���غ��VH��@��@�P�%�>"H� ��ҁRF�X`�+4�B��HƥpbHS$�J2��X܄4�#+�¡��ae�����3�a`͚�E��(D#�H�������h�3yB�,�sr\����ޓ�.���!L4���_&p��Wa��!	<�X��CL�1}���I��Ѕ*�X%�%���K�.Ɇ������g8~��n�FH|�1�\��d3��.c.M�g#)�5%�p�n���	r����X��\��C��*��HёXP�S��\53���ӝ�3�]�BK�:H�0�{;Á�|��oǶ����&�SH�"$�"ԈL V!P�B0�"Ga(��`DbBF h#  0H$�T��c�rϜރg�$6���H�`H@�X��!�Ąb腈A�FB�`EQ�Q�� 5p�TĒ+D���$tӿK�H�8�����3&M0�$Ԅi���
`c�����5�S�J�����"\#�
L�W4�$&�:�I!C{��������)#8SAl���L��D�0�,!��dd+B`����]�ϵ��\~4ţ~����%i=9ߪ�#�������(��tA6uץ3�+N�$��Ӷ߾�Z&�Û�٢�}���	4l�2-`�hS�y��/��CL@��W�3{��gٽ]&�a��H!�h���0����)��+HA�b� HA��+$dn�jV0�FF�YX1���� ِ�
B�	u�u�IB�����wi.HP�v���`B��O��a������M�<��FF�3Z���d�!R6,3.�r���73.��SڟNA��|�r��t�#;BŬH���m.���t�H��E���d��I�@�Uew{��i������hn�|>D�D����36N�h�ݓ�cti|M�*¤LYs�����a3[�W_$��}H�$����0�����a��p��x�%�d�M�3�7tc	HP!,Rjj5���6@�rd�Gf�P$!���-֎zt4�-0���X�s{��i6��%��H�H���S>�}Ii���B�HZ.$I�BT��0�i��H�(bRD\0ki(d��*�L$j�lR��8D�J�$Ha�ָ��n&��B �	D��Iŋ$��:�B�,�ѪB�%�DɅcc#R�d)�; M1/M�~���k��U!H�38˚#%1�!]�!q԰h@�D��x�W�!p���>zF?$d"@�e�2#��֧ȕ`�41�@���@�}� A�	#DdXC�%0���5��^T��D�f���&#�$�8�L#�#I��K�Hi���oM��������ac(���}���l!��=2A4� U�hIiN�P�2���H�i,+]���>P��@(-Ϧk������p�	\āS1��0 Q�"H	��h+p��ɛ�=`$!����6$(@���	z�cR(FQ�G�S��:����V�#��A�
JH�,`IF����!6[2R���Lo��"����6���M�bT�ѺV�q�L0��GJ= I �5�B@"x�"-HJ����]�w/.HAd��Ϗk}f���c��9�Y����d	��)c7��f��u'zY�%����ﷶC��$�|:J�K�a�ޥ�e����"ԉV!H��N\��	J�		$�#8���D�XXa��ffsZֵ�kZ��   6�m�   [@  �     $ � l[@    $ H   �h  ��     ��      h  �*�܌�J��r��J�e���c�ةYX6*�Y&��WJ�q-q[d8(-S�«v��q���-���08t��l�5m�:lOB�� +v�jڔ�Uj���G�`ZY�� �,�Vl� p���eڨ��j���J�[@m�	��<����ky�0I����5L��UT�P��p��V��J��p����������w|��5 ���`+n��{Y�)�
��؛��l5��ҭ�/;���)؂@ Bje��J�����)[M��[�9�6����=�[[Y'F[h��s�6� ��[�b�f�[���l  n����iV�T������UT��[@ hJ-��l�ͺM�m������ �v�޻c���  l3���z��ږ�Ί�v�[p  8��%�4N��+��Sv�6#Vc���P�+/J���U2/A��_V�9�m�8R���nX�Z��c.۱u,
-��%p�4��#D�H8  ^mvm:t��m��n�[xHm +�]�j��;C���UR���Թf�����8Z{Et�Ct�]R��&J�����τ�r�UpRqq�-U��W���Ʃ8�UX5 �u9ٝ>|�x���xM�V�j�:��l�3�@v�q�x&�u�*qdn��
Uu�,I=��vkn j�]��� m�N_I]QtL�$M�y�v�*d;eɯ[����� l]Xp��R�f6�j��$-���^U� �_*�Z��Zڌ*
��K-TV7l�y�ڥX,�s��n�B| �ꪪ��,�� �*�R�E�!���I�d��'��V]�6�86c�-uR�ж���l�'G[K��k4�Y�F!#�<�\7Q�2q�6y'�vkU�(2�mJ��!�}m��l]Um*��ݴ������V�����H�[$�^�H ���,���͏���|�u��!ڻvXV���Iz�� 6�D�!:
kw��k�}�m��6�@�m� ej�� |�����i|���%�-�8��y�Wj��<+�4��s��UTpK[   ��	#@��� H[j$�� �ףq�Ͷ+�[@l �̸* �mm�z���v�� �Y��n�r��	 	   �`Ն�H��	 2��[�
�[��ڶ	n�-6��.�݀Hݭ�  ��p��Y!m��k�6�  6���m�u�$8�  6ٶ�il�gm�ޠm � [�� 9ŷ����� 6�-� IJ�^�r�]���5l�mI���R��3;,0�����d$ 8��2��i��[A�L�l 6� i6͖�ۚ\9�l6� �-�kX	�Y4�4T�-h�5k1�  p [@ �` �`m��� 8�`k��%�-���it�Sb�ZWeV������zv6� lf�u��$���ŵ"��l ��m�� m&�$$ � ������ ����ϸ���W,]PJ�P����hJUU��I`�.Z��7i5ۜs�>o=l'ȭ�n����֙ސ��;��<G\����Y��ۢ[S�!� m����u/;�T�J��Q�M�m�6� l�kzO]�̣⊕n�[LqK�U�+���H  �`�޴S���6��K�0��T*gi�նƴ��2� ��(��m��R� ��]�e�-t�(�[\$�t���cl�3v��!m����MiL�+]�L���q�ڗk��ɭ���	/Z ��m�BH���eێuړ� �:[6������m �u��� �v�ڴ54�ѻ[��ko �����`ڷ��-��6jͰ$��{]� �hN�����@iV�ã^�U::�8۞(
��`b�	�Z��Ϛ��|� �CT��fֲM� �d���m��нjiRv�m -�ӫ�mp�Y��,2K�j���m� 7n��ے[���-�'Z)E� <$ۢ�v�n�R�{L�m�&J�p"!u�N�L�Pn� � mm�g���l$�'�E�.Ѯ�m��>]jG  l[B�m H$��6�!�M�W[��m�#�  ��l�[c�� j�` 6[��/�]~�m���`�a:v���l-6�l�Ͷ@���¶�$�k��i�D� m�����{��$ 6ݐ������6�$   �U\�m�Ry����@��r������J�J��� �n�-���` n� �vؠj��2+ķAUV� 7m��)����lmUI�el�*�` �l u�z� pm�j������� kX-�Ͷ6�@   ٶUU@T���Ue eP$�����f	�d�UU@�T���32�u�8�� m��l�{l�2�U*��VZҭ)*��b�J�UTW�k�۵��H	 )[fͱ7K�A���� �����~|�m�Z�UIv'��9¦�R͖��p �i�m�%��`]U�@eZ����X�j�[5m6��m��( ��� l�cj�H�X $Cm�J�rdj�V�6Fxѱ�!� ���p�[T�F�
����
	�5O:����gI,�$�)% :��b�n��9 �c� h�n���k�L%��6��m�i6m��y�]7e%�,���A�a��y���n�^�(i6ΪM�8*��*�l����2Ɲr]��� ��;�9 �D��9c�.�k,�q:{&��@���WAJ��� *���!�Tzt[\.�&�!�d��q��H;�mv� &�k�R���%�t��N���mյ�-�-�l��`*:���Pp@���À��tx�uu��1 u���bM�v�m�h���GUWTD�`�`ڐM�m����i���)��FC�l���mډT�h�3l��&Gh붖u���8'��t�m�a@ IrRYx�e�ŶCU�p�����5��*��������U�N��3�S�*Kժf�U��k���h��� �Q�*x��hh;S�;U�*�5m�l @�$�]6k�jclm� �A���A�[BBݝAWJ �� ��0 ,�o  ,1�̉ 8Hn��ж�����h '@� �� z� �`$�kQ+�f� ��p$	��a��$ �Wm�	   �� V.n�m���ăm�-7n���� �m�ۀ m�� �a����@�am�GP �l�Zlp�F�   ���  kn[M�`�T�cf��e���ZRZ��H�l� p�[@-����h�� �ɥ�Z 2� I��h#���n���uf�m �m�5�UmZke[�������m�m �{� ��m��$�����`��Kh햓k�ݰ p�cZl�K�h
��] �WmTm*��rJժ�#؅�R����iέ� �o�[ S��ֳ�eucUI�.l����vR��86���B��ک@Y�v�M����`�����$ ����Ϊ�,�� �8	&ݝ��� )[f�I�کV<l�on��YO6� �ko $�b�:ԮSf�����M�6ٰ�F-�����    � k2�wViR lq�5���e����i�[_>�����WmSU�K �T�6A��8*���	t�y�>�	x���z@�������w[#U@K�@[Kj@m�m�N�nĖ�$$��8�`��  @   �}#j�m!%���`  n���m�a��mt� 9olH���)B�����,� 8e�M��Y6�ޭ�M� �m��Ci�'4Y��/6vZ!�m��z�V	Æ�UH��2�v�u�*���P���m�Rm�,ײ�� �E��h�����mrBM�I��%�I�l 	:@8��M��`BK1�7F���   �w��  �`  ݛg-�i H  �ݶ�� lq�մeo/���?+�U�O+R��s��r�T���]�P��������:q4����P!K+W�*�ؕ��T�U@Uu�T����^��  ۵�zkC��  �O6�[�m�۶� 86�}6^����n�}}��n�)J�m��=-�����A�6ہ&� �@mt����U��h�m�Vѫj��Zћ\�����W]2�)�;ح�VN�[����I��m  `� �6ͱ���6�`  @$[@6��0;n�ӕ�m�[\Hs�c�l84t9l�l�:E��!q�j���n�'8!:-�ܪ���b,zmk33��6����~H�x.�"�_�U`��|+�J�B	"���VE�O�@R��hS��Ph���Pt����~BhCH!���Љ�t���.�������(��!�C��8!��"�S��\�c`""ȡ*�8��p⋀ ��	�ꁥx'��@
|��(� ���B��@ڢy.(��;��;M)N������`*@E� 4��� �A}� ����yDv'8*Q`,@�И�TN*p@��ｊ� �*��"�ʞT8!�h^	�� �h�Ab� �>��ހtO�V#�-�@q>Ҧ�Ҙ�|����!E4�|pU6�����^ �F�hT�6�E��D�:�ᨸ��6)��6�T!����P�|� z	06�tE>5h�� H� @վ� *D !�>v ���	�����8�u�yPк���'ʃxJU0ӏ��")�AЬ�� ��P���#� 8��X�@!  DA�M b �*(u �!��Hy��5X�bԢ�B�hH'�u W��:���@��8`	� �(� ��(��(�T���|kh�A�r�O�?
�U8�� O��v�� 
��_�`�Z㈩��ʁ2�*�H b0�X�I HD $ Q�T>�{z��Z�V���m�$���h1��H�I&�����Y�6�u�*��[ũS'N7j�9��Senݼ/4��H�Iَ�s���$��^U�8��Gbq�����b�����`����+֦�l����n�Llr#]-�����ݞ�����C�FA1����i;��f����=N�ِ��Jgnٸm�񺇵�#Ӱt��OO�����٭pQiby.��<��{F�ڸ�2�i�)�ۭ=CӬ����\��`����lT��T#$�x:
Q5Rc4V�\�h�18�
���c�=�9��m.���QzQ�Y,��DL��+l�vũrMm��Z�XI_L��<��<S�7!GQ�m�j�÷.�톧psg���G0�.,��-h����3�B=���rp�`۰���w+�eͳ
�� ¼u�fd��ܜ��n�:�,9��d�-�W"�d�vt�i�x��ܔ�.��s��d'�!�XF3sV����o���3tv�k����I���.6�y�]dF���M:�ei\�ܴ�[1�j�n�U��p�i$�-$����N]`v�J�@�n��9�H�a ����z'	�6уɲ�Y=!�qk��b��E�k�ۅ[gn����3�5D��gV�uKyk�k�6��ݙ��I��ԫ����t�m�	k\]����4�yv6<Y7"Q�� n��������J��e�ݣ�'k�m�;��,P�K���P�
���^y
���8z�f�!����0�ʪ4�Xn��tg�;@Y�;7�T��h7�g���p���l��`�u�J>�N$�MR����&�ۚ�R���#���2�!g�X��q�e�ӥvܰ6֪Cv,��vz���gN�;s��s:=%�^�]�vVU��i��W"p�<p[z�����
��;�����LlW<�$�	n6�3z��;d�Z��u�Q�F`!J�V��k3Y5u�ֵ�q��T�LW� 	�*��N��D\Q��	�� �	� ��z��V����]>Pb��d�ߧ�S9��^��\�n��j�]�k�䎝0�\��d\��vˢ�NdY�u��a�k�l=j��i��3s�x�y��v�c2�EƑ�v�f"��]�&j��!���[`�N]��m;�`�;�TX�]X�= rzࣱuF�L<&�V�8���v4u"n�Eu،���lE���M��ssǳ��s^�&���ʇ7',xό;j�����i�hF��W.I$̛���a�+ɐ999;"r��
c<���E9�8���zݸ9hmށ޽g��XI<����h�Q��CR-�ڷ��B��/{w4*Z��-���H�"�7v�ȩ���Ih	ܒ����	��`�4����ڳ@�v���s@��,��&G�{����.��%��R7#o�wq��w��p;LC�D�դ\լ�ۚ��lv�y�Y�.4:�{v��^Xk9�+7p�ݺ�<�� ܊�����Y��u;�G�$�6�Z-�o���ybq!tD�0t�C�t �!@|���s�7$糵f�x�Z��ea̍ƒ�f����H�9w�����H�]�Q��x�0Rf�޻Vo�=��-���4<�}�٠w��{ �i4Lw��t��$�d��ȩ �It��{��w�}�~���GKls����\����8���T��#8��G�=�v��S����7+o������r*@7�] #v���S�<[0�<&�3@��s ���X�78ͼY�(�2j��"ɑ�<&()3@���4�jә�@�
) �}���[۹��q���F9��4	ܒ��*@F�y%��ˎG�&<#mŠr۹�^��h�f�x�Z���U��HPq(�q��������iM��+��N�3�6$�6Fx��"�g ����4�ڳ@�v������cd#Ƣo%�H�K���˳�=�@?{ʐ��@�;u��j4��ے,�/�@���Q:�����X ��UR|.��4���@vH����H�URE$E pD��M x��k��.����0��4L�swi9h�K��Ih�|�~_���g�KÛ�)9����kGf���)��Y��S,#:�gy�V��m4m^��h�K��Ih�{��}a�o��w=�OÐm@�#�f�x�d��ܘ�o�K��>`�e9�L�0m���[��U�ק�>�+]���~��8�u�����!�V�6""'i���ݕ�?���>m��9�v6B'�6�cN=�v��5B�^��ۻ� s�:�w2T)XBw������,�6z�ug2k&��YqHk�9J^keC.�D��6�ۖ����b���/3,�;H��8J�n^�ڭΖfM`�������Gu�9^��g��8���$��ya�V���E�Ce��>��=�E��ZXy�����=��sٙ��]���R<=v���T.�Z�.�$"��˪��omp���1].��xN�Ͻ�}�v��S|�!��=t�bќd�n,�#<��������ֺ�m<jD3�NX�\I�[v�{��h� %�1 �It��jJ���d�E���p�x��"��o��k��h��h�Z�1�fD	�rL�/�@�]�4�j�9]�@�Y�!L��1Aȴ=�}�{�4W�-����h�܎�rq�br,�/]�@�즁z��Sr�J!-��A��$���*jbS��� >^:���3�pC���%��Mq�L4�9�L�0m��;�<h�ՠw�՞���? �~��8�֗�4�6'�ɬ���'����<���?���(��X"j &T�"E0�`@���~D�=�_�[����V���S}�G{�ll�D�D�3h��@G��H�K@}�-Ɉ��֛�Q����qf��>�^��H�o�x�qˤIf]��H��rE�~���=���/��/]���ڴ�s�b��H���	�m:��F���\lr�o����q�5�F��L&�����v��/�@�즁r��B,�#�b�q`�����$�M�ݬ��L�np�nGV71�%�F'"��k�9{�M�S���Cýۚ�nI��M��w�K��#�&LJG�r�S@����ڳ@������.F�Ƅ�di�@����ڳ@���^�h�t(ޤ��mŏ#�3�y��g͓]�c���9�V�H�"tq�Xmu[�I�8��ڳ@���^�h[^�y�u�5�I���"��k�ffL��z`;�X���f��2��2���27��Y�@����ڳ@�����xƞ�L&I3@r۬�M����вQJ�"�T(<��o�x�N��A�L&(ӏ@�v��=���f-�ݯ�7�� r۬�-CWJl��6�����v9�ȫ;�^��e7a�[7n���cqcs"X�br,�*����s@���Wj����R�q��ɖ�*�y�Y�!L�;�X��e`vנ~GWk#N6bx��f�Wmh̒�-Ɉ�T��na�m�(�&LiǠr�Vhvנw��h�ՠw�cHj�F��i�E�]n�I&�/�k���>tܬ�
>��H0XP��8In��E4d֧��}c��c^�e�L2#oAb�V�t�s�Yr�`���"�Ǌr�&�nWV�%K;(m�uW!��Է��g�yꭶ�-kzB���.[
s�C���K˶�a"=`m�ك��v9�+m�������K�9� t��Vݘakvf�v�R�>�ɺ�X�sǫ�����v�ݏa&��}L��nՃKk;c�z�glW����w^�����ٮ��i�M\��;��{ysq�t�(b�B�vYH�FA��Y���@��� #�-ْ] %�1 �*<bOZ�&$��U�^���Y�U�^��۹�\�Z��dR1F�qْ] %�1 ܊�䖀�nGV71�%�F'"������q/�bW(nl) 뮯enmf�n֫D����o�Fמ���ŀ?�j�N��bm����b�jA#����.�;a�d�x��v��N&/n���gH�U�f᛻�_\�r*@N���+>�����s���ɑ'�%��q�N��ٿ����|B">���;3�h	$T���1 �=˫��1�4�s4�ڴ[w4
������ ��P�s�"1���j�����T���-�
�X]�j<&)��L�*�k�;�w4�ڴ�x���b�:L�L�*j��Z�G��E��7"�vF�Y�Y;g��/a ��;u��ݸ��N2) ��N?�[�nh��h��hs��-��71��Gs��r�~�� <�z�z������*����nL�>R-���4�ڴ銚>&O�7|~�<~�����(Jl8�.�L#�a�F�F0��%H�{謹W�ț��Є�8t�Md�hD�`��@dU�	�(P�����HEX�=�,h`�G�!�jłl
� D��aF`T"�`#
Q��8΁�|��!�6)�p��oP�B����N��6�%SFT$)"F%̢�����(h�VwX0��gBV	��H��ѭ��0Ć5��$X�|��A��M`f�V�Tѭp 	��H��r��Č���d�~P<''����<��ΐ$c�h��S}$�	���a(tb�F$3��(��$�@#
)%�逸�Ap-1{�4�H$j@�=6�����E��!�S� dA~��Y�H!�QdU"�D"�,H,*tU�:������UN�,P�%�	$�g��X�=���Kt]MF�Oc����fg�ݗ�@����*�ΰ:(���w� ��˪-\�Qd���M]`�x���^ݯ�{wq`{���ϗ3��y�6��G�'%��	[�'�����"���s�'$���v������_�|�� �i��������hv���B��w� w-�*f�	��Sb���\���& �R[s�Ur�w�y�z�a0�7$� �����۹�qw����h.v�"��L����J[���K{XͼX�� ��5�� 
:/y��k���@��܌��(,r273@��k�:����������V ���j��UT���v��Gl�ݎckM����sk����R����Z׵7�s$�&8�2|!8�w��h;l�;�w=�U�z�W�4�f,��376��M@7"�m���1f̞��\ҵs4��T�uWWx(�{߾��w'����� �{P�n���Y�m9�{^��۹��l�����f�w�|��� �C$��m��::+���݋ �}�X��;�|�G�Y��w<Ekzm�Z|�d�OE����ك�`h,a�'j`�Cfe�D�`+k�E�v{cn8�nv�2�K���񴐄V�ف{2'6��6f�C�nHr�{3WF��=���>��ˆ÷Su��n{1�����[��U���O�̧�S�� \l��R�N���F�P�[d�r�s]&�Y�1�.N6��8�˩������]��ݺ�o������]�n����L�6��'87�����ƃu�Ϳ����<��];]��6�}?j� ;m�����z���8� x�rM��s|��o���zx�ݶh;r2��qAc�������d�#�ʫ��������.��Ƥ�O�)��e4�m�m��{^��]W#N6bx�37t@95��{��s���`���U��!��#�F$@�f �e}�h[�`�����ʜ)����=��|o���<�ê����=�ŀ}>n�7l�Ir���/����i��&dc�i���8�mg��DRDB��4�F|~̽0�{x�x��(K���ޒ�j�HYJlWu������@rj6�� �L@7�懭F	�q�C�v��@���4.��=����@���zdX�(������R����`�:������������p;]Pp�s��J�@���H.�䳕;8��Ƈ@�n���\����n�Ad��9��=��h;l���A��,�yr/T�����J��j��v�Έ�S!�x��X���5DDbGQ}�'1<q�� �����{�74(D`�BK�h����1�j�����F"Q
$jDX������$��K�ߧ��`ݽ0�7�4�ZOK#qɡ��_{߳@���;l����ϒ����ޖ5���� �V�����
9$��~���׀v۹�g��s�|����L��X�Ô::���g-q�k�Oa+gX�J�H��n^�:�\?7y󚆓� �C$q�O�@9�f���-�I~������mEMa7E�R���� >�w��9B�7��`w���)���1#��y�crB x�rM��,��u����e�ޘ�x��5����P�9�ϳ��}�{��~��O��krqb D�d �C�{���N��tܓǉ����u�Z�I5u�y�f�
|�o�wq`]���g�2���B��7ń�ѻDs�B��k{m���|��r"���Rfĝ�o����nlrCƣrC���?ɠv۹�qv�����O;�lO&D��,L��]�m���EP�{� ��� >�w�/��!p�k(�F9��������0�2y�� �w |ל�MZ
2�J����`�:���*A�}�.��=���OE<I��y��5D=����{��y�f �
��w{������)3��%ٌ�<@��k�8��uUSv������c����%�i����7 O�WP<�c;:0�{q�Y�k������������5b[��8H���Sڱ�Wk��@��e��:]O��$�9��'bu6)z��g�sb�g�Z���83���[��Oi��r�h��њ컃�C�.qS
sn�E��,���+rbG�����������8�p�lk�x'J�]@�k�y����]���1�3,e�q���6[tr��7u�="�mɈ&� uɨ	]�k+�(dP�9�mzm����4�w7��9���^�Ԓc���WX{���7xj�>��X���.H���5�f����g�6����ذ����(�������v'�"I�,q���;m��=���g]���/��� �m����l�GP��Lv ��n3���2�Q�k�s�ۡ�q������}�ن�5��5�c�hi��U�����&����ó�T��Vz�&��6+���>��,Q�p���^��0�G�M��EQ�(�R(i�R�9�j׫��o�u�<��rb�.��^��k	�E)���X�x�7���WU����}��[B�2,nHDOwP9 ;nL@u���=�@z���y�dL�`������������{� ���`J_zڹS3uWr�͌�iS�����]&1����W�n=���o,�=ų�Lp0Bq���s@9�f����{��:���#����Cʛ����y�ΈK�U��X������gىｱ<�D<�Ŏ5��~��rO�}���D�)�,�- �#YT��h��н����͛�U���s�cX�F�Lr1�h{33�=���ŀ~u�8>��0���M@�!ۏ@�m��=�g���_��<h\�z��Q�\o$B�u���	n� b��)ƕ0ݰd��[�W����;v1��}�H�׌ORl&qɟ����>nـ��{	D/�����kЉ5$"�#qh�S}��f$�o ow���9�%2}�w
�TU��J������=��a�
*���8�0��iժ���VD���D%-��XΞ��v��|�%B6�3���+����CNy�P���krO�d��M��]ئ�swV�ޯ9�9B�P�$����@��PH��d��WyFee�]��g�n�ulv��$b�Ĳp:Ӡ�-5��s4O}�Mٱ<�l�Ŏ!��}��@>nj�{��ó'� �/�.�4˫���$����}��}��ۚ+�Z-��gٙ�����` �mU� ��,���p�P�L�v�����=�'J����E����X��ۛӀ>�� ?{��9(K�I%[��,{��d���܅)WUs�|ݳ �.��Q^�����X�W����"(�H}�:BX�1�/ғ@'�p��A�M���3D;t��ŉ���>`�O��$���^M�H�}L��D�	L8�� ��wA�M���ϸeaU�^L���@4PN{^��Mg��H�%��@� ��
D�GL�	sK�j\4B'>bD!}�~�h��=���S�4G�H�#C������'N��0]!4Vd�%F���hbP�0u��mֵ"ۭ`�6�nZ�l ���t֣n��A�y�;g�ɰ��-�rI�1s���B�����M�<�m�Z7;pkCF�r�䎜su��u[zv-��	x��M�ٺV 'm�*�UK�5�Z�wn�Xs�*�s0[_�%۷��^��=��K�����a��n6�v1\uHz��Б�ݻ��V�:���CW4�<���X3��=�٫�^y���}��p�֦�v�6�;���m;�K(�pYynte��phՔ��X�-k�=-U������Z_��ƃ�3kFI�d4\�Wd��Pg���B\��j"�U4��u/a�eT�u�I��MS��t3��݁;;U�t��� ;��Z:� �v�`�l�U�"j��C��pss<��Z6ͥݝ���FQ�6�8���l,���;.�Z�B�6c�Rp��Oω�����.�(��\�A�ct�t�jgEj�1�*�a���J.�9��h:��U�\�9�2i����鴙��,��䏛�K$�[UE]Y�yĺƴz��݋sl�@��^$�Z� ����N9$�����Ä������eU�]��э��UtjYT������mݭ�糓�l9���q�;%�C��
��Xdy-���hM�$ײ��l�	I&�!r�mZ.�ڍ���u/Xo �ԧnՎs���\j�j�96ۦtA��]�Ң�5��7`�@T��:GF�b��{Dt+)A!u.bV�Ύ�V����z�ܼt������O-�
�E%��'cP4�b�jݢ$��"�� �q��O>�v��F�D��� �z2�pi0�Q���U63Vbx��l^ؽXV�ކ^�������k�Ԓv����`3�Vԇ�^����ܽ��-��;���P..ոÝ/c�u�ԫS�Ҏ��\��qi�|o�S:˶nMi�Z���gc�G���8G�3��Ν��pSzv��}��Kv68{+�$�2�b�:�35�[��k0�eM�\� ��N��Gc����$@���'��"'�~|�gAC�O 
�`���{왚�f��Z���۲3ٵ��5*��V��z�V�JHȽ��nu���mU��k��I�[��c:�iA j^�#'���c���2�/7=<N���笝�m��;L�VF�]��Z����3�gb�Yx71!;bI5��Iܱ֘bN-ЇZˠ��ׯ��A֭�GڥLnX�������iS���F����wʬ
��Q������(�{',�5�֮̳5ke��ՓV�u�q��J;b�V�A�2���=kf�ח�{���|��+�ڲ�Uݪ���ϯ �o���:�ٟ�_zx�=��	�&8`���x���D.JQ���7������gؑ�v��"nI�)�R9�+�X��aܔU���7��`��˚V�M�X��7���W��Z�}4���}�|�e��/������S�$��h��=\�rO{��̞�fI6�~�7�����d��=]xw/�����7��Z�ݖY0�{c������)��ڹ$����{�����M�(K�B_P���7x]T)U�H�Z�������ﵼ���A_|:�I$dP�@ 1OhS�	�����p[��=��gDrQF�V!\�U���Jf����8��xl$�[���o�����Rc����Z�L����7�� =�;��$��w-���D��c��	ɠ[n��ϕ�������~�� ��n�6�^ָd5��3�s���;\�6�ۆ�sn4�[m�	�b�9�ٺ���'&I�9��9��-{xt�������wv,�{"y2$��brh�V��H=��n����w��Uw�*�]��6��]����{z��ŃO�PB �9�s����nI��{�����U%����B���9%�DDB��� k��np>[	%Z��|g�1=I0��$9&hy� ��DD7m��6u�`�� ����#�M١..��X;F�Uܥ�Ş^����gq��v뫵7~�w������-(g���n��������b"�}�x+/�I�s$Ksqh�l�}�ٓ&��, �n� �79��L�4V�͓wv�\
n����X �n�Ԣgv�V�z�M �β䉸I�9��9��.����^�]Ӏ�w��4(P� ��:��;����7$��oV����W2�U�Uw�7M����������X �n��r���YU3Jtۣ�azy�:wXN������p8��X{]���Ѹ��rcX�72I�����-�s@/-��? ����
���6���I(���or��T�� ����پH��y�5 �lrL�����s�̚����� ��^[Ńr6��(���^����z�M�)���K�������n&9�%�9�Us��w�rP��w~��}׀7^�ܓnD4�8�	R�����Rh�n��q��؞	�Y��3'��%�%Q�V㡩U!f��"3�LR�:� �e��N�Cm��v�V$Kz:�S�-kMS��S��غ'sҙމ��Ҩ�k��Y���:�3�bbjLo0����Czl`�#��imnOV\F-�܋F��f��ά�1�\�<��KsLDQ����%�v�ϖ6�>�:�����y`�)���{������S�2��k)�[����;v6�uY���	�R����V�s��1J3(˪���VSuw�}�|`�������%J;���X��\M�S	���f�fg������}��[e7��_{by2$�ıc����7kvp�<XjS;�z`�v�w�R�&5�̒d�9�����}�4ݽ0���jJwovp;��UIh.���DM��v�����s�����/{w4gmz�Rd�<�LM��=���>)�9��;��j��<���s�U���=26bf�D���? {���:�]`�x�%�C۷��Bw.�*��Z�an�k[�v��������S�*�]�ذnޘ �n�(�U�=��D�1�c�6�z�����r�M5B�
d�n� �����ST�j���X"n���I%>׿� o�o =�w��:!DEv�|����]̪��)�]��� ��Prj7 ;$T�w̫��,@���,�H0&eLn���vy;r�A{G�� z ۳����o��]t0)UtU]��ݬ���o�P�������}�d���I2F��@��Ŝ�QTn�b�}׀}-�͈J��y��`F����[�nh����H	@�"�k�j��g�g6�s�@�o�4ڲ�ba�(ɫ��X�"&w۷�zwv��<X	%�	*���`��t�UU���Jf����X��k{�~��X �n�����~o������5jN.tt����H�8z�B��ՙ��@��G�Q�sC��]]UU��5�ŀ{����w��:��=����&��ģ�4��Y�BS!�ݼӻ���!)%��[yO�"��A� � �����5�fkZ��f�4lA�lllo������A�A�A�A�~��6 �6���{��<��������<��������̚5ndԥ3Y35��<����`�����lA�lll{߸lA�lll}�߸lA�ll9�� ��_�:x�v=��~��A���߽���֌����\ֳb �`�`�`�����b �`�`�`��~��b �`�`�`�w��lA�lll{��~͈<�����IDo-韮������wv�T�
�*�GE�E��V��6Q��&�,�q�5����{_'�,�&�˫,%֍�?A�������y���kb �`�`�`�����l9���y~�Oِ̓���̗5u�y���kb"�X � � �?~��y���y{��yO�  .A �`������k,���kV�-��kb �`�`�`�����͈<�����{��<���X � �߿p؃� � � � ����[y�����tf�5����f�A��Ql{߸lA�lll}�߸lA�lllo�����<����s��ٱ�A�A�A�A��k���.�Z3R��kZ6 �666>���6 �666��~��[y��߳b �`�`�`��߿p؃� � � � �mg�fe����Pc�����M��^r=y��m��bI���Vb�=f��b��-��y�5a'2����Hg�������Y6oK�o=(��Rxm����9��q������ll4�mG`	�;c�jٗvn6�	��p	�å��;�H�1b�㡎y�W��u�� `��������Og�x��Y�]g��؎����k�5p�Y'�.�0�ה�?����g6�i�RM�i�pװ��[c	�#o��#��g��&m.�߾����b��Ⳛ�p�ۚ�}����؃� � � � �?{�lA�lll}���@9~��M�<�����~��\4M\��.Md��lA�lll}���6 �"�X � � ����6��~�A������M�<����������<�����߿r�Zє��Z�Z˚�lA�lll}���y~��M�<���67߿~��A�����߳b �`�`�`����?Y�f�5�]Yf��yT�A��o�؃� � � � �~��[yg�~͈<�����0PL����]�<�������_�a8��K�ֳSb �`�`�`�}���lA�llP�I	D$�^�B��Hn���]�������o�~��lkլ�N��emW,NC����M�t���+��vp����D��nn��u�`ל�~�tDD~�=��v���"b��2Gn=��]�M�J:pjB�i2�)�,f�b�"�ޅtj��q$CH�5�����N�~�U�{�>�"�p~O�QɎ	bMK��0�;Ò��%�V�oV������kwm�")������sc����Ur�����[y�	���&F)&��{^�����ޗ���x�{f���1�8��"�ҥv���19��)Z�� �ny{t=n6���R?}�}�a7u,�cX��Hӑ��wӀy�ـ��DB�С(��g�� ������0#B�FH��;{)����~u�7^s�	.J��{�uP����&蚻�� ;�� ��:£!$F�4p!\�H2p�#�.�`��y�!�@��01`Q�����+(hFY2P"�2Z��ȫR$D"D��H���Ԍћ�15���� �hlڟ9���P iC���B= �LE�PO�H!��;m�9��	� (�I�X2bF!C
�_���bR,�m��������3�!�e.�T�H�|�����.`��@�� $�I��D���0�(�P�⩎�8�P.�OCK� ��b��A�*��(���|��� T xtW��4�S�hπ^������ܓ�ߧ���܏rI&%�C�g����@{�=h� H�:�6�SMdqF��9l����>��? 7�xtD˝{X�[�h�f��T��qcV��yyt=�����"�s��q�F��S���d��z5���!7�_Y�@;�� ��:�	.�P>�� =�Uʮ��")����@꽯@岚oe7ى��lO"�8'#JI�9׵�|ݳ����������wR�&5�̑�9��w����7$�ｭ��`�`�1=��@/-m<J1�oe4��o�u�`7l�:'ۻ$�M�*��m]�5��>Ltz����;\`^��E�By�X���5�ٍ�8��r7 {���@꽯@岞��/��{�ۊ	�$��I�u^נr�M�ڴ��h��q86�8�q�ۏ@�2K@ɨrL@:�/!��LpK����f|�����zhVנr�M ��ڹjH��diȴ�5��-�6�r�����~|�	gj���sNmew\�a,t����Y��܎�n	�u�|���r]�n�3�v{]�m�m%&jb۳p(zp9�e%�yu�i��6��x�NzX���
����`�7.�X�/V*�k��5[p�[Aums���q���t!ۮ��r�80����)���:5��3���ؘ��ncV���^��j�(��[�� �i�=�ݻ,�Ȃv;V�7��{�>c'/�{*�8�s��]��^��':�Q�m�ab�����tcW!W�m�}��~`岚k�h{l�/;�f5�̑����S@�v� �m�U���M�G�F!C@�v� ���9(Q�U[=�X�07)ҡ��NE"��٠u[^��e4=���=���ܒD��E&��1�q����Og�h�5 돽������cY�����v]dU�wXƻ�9Sn�ֶ���z�n)s�������%���r��'��@\���j91�,Bnk�k��fxF*�(��T�~{�?s��䇭��9l��~�n��b�r, ��� �n��
!L�v������v�O"FI���$��{3��������f��UW*�ۓP�n��cX��H�9��e4�j��٠���쾹��F��3C,����z���n�k݁\��S��&l_����7&�6�%�I��������Kn�Q�A�0�+iUMaKQ��R- ��U�����;]�}�ff|��T/n(&�r���L�����f����H�D��+��>�u C�(������I=�ޚ��Rcjc�Ȝcq����<��?;�ԡD����>�+f���2c�X��4���}������:��=��h3����m7�&')��\�nzCIF����^���*i.��p;�����](�d$�Y2)$�/;f��mz~�tB�K������4�L�
�q�$�8��}�G�g���?���������%����H�G���{)�v�V�ؑ�_M�{�@��ih���D�"Hh|���������m��x�Z�L]�ٽ��;�S�d�ܷDi9�@?[f�������l�v�V�xc��1��&)�CJs4�єȹ��W3�d�w>8��6�uv��� _9�܉�	�'$�}�M�즁��_�gߐ��4V{ؤmLq#�rh�����U��8�� �n�\�Q�EmWMMիUdʒj��7��p�&�$�o`�+�3%f�Vn�%�"NE�������;��h{>�_Oyh��lO&%�!�rhkw�t(P�6�O�=���ͻ�!B|���) Ne���
��.�!�������~�%�2��WV6�FX庣�;��mw�{���vrMn%�lH�v��֑ҺCsL��c�%�'b�@�#vݙ㢭n��qnV�I�m�>�*&��p�M��Wj�k���*��A�kK<��v'/v�WGm���D����pQg�n�zA�������ӊ��1>��#q�hm�����'��k;��r����&��F��9�.��6l��a�Y݌}=��w���|�n�þ5���;�RF�4p�p�.M�k�n��ܓ�k��?��z/���&'1ǒD9'����Ɓ��Z��4�k�*�ih��Q���m79��I*��w^��Հ{޶f���g�1��NE"�{ޚU���e4�j�-�J�8&�Na�j��6����w��M�$�!r��w^�Mܖ��Wwd�Uu�{�`�s$���P�j ��3M��::3�#k6����Lngt5gA6D+��k�-�?}�����n��q���l��g ?6� <۾J.I/�7v����+�����ʥs5w8��yj F����S��~�'��krO��M�ڷ�}�$w;}�9�Fd��(�]�׷�{޶a�%2��� }���?�s*���5j����Uw��	%[���z�� ?6�T(S/^��ޗ5J #ģK$4�ڴ����{�����;��h�9��Ri�H�H�/l�r�]�Њ����l[��j��<�m�<5��1�Y1��NE"��{�@w�o`�s������4��"RI�u^׾�>�-�Ɓ|~����f|���{#�2F�G ۑ��� �9�"8�$yD�R�DHq�P�B���+s��6~{X��S��1�X��4?�>�W��h=�M����(J[y� y�l�d�wj�)\�]� ~m��	ֽ��6�L�����u|Y�bO�84!,��X6����UAa�6˹�Pys��@�A�g���ۏ��`Q�"$�8��}}4���k�Z��4�ıٍ!�Q�ɠw��g%	tDEQ�[Ӏ���?;��ijb�<J4�C@�}�@?[o�QToo^�����N�XL��#IȤZ�3��U��w��в�00�"7j�l>��Sf�{�]�;���ٚ�Y��Ԛ	����=/ΰI.������7�zp��hJ[�4HH�&�$o�V.mW)>��r����-��t����v��Tm]7k$�dr����S@�s@���fg�{�z����9��&�y��;�(���oN��Հ~�g$�H9|��9&$"Q��;]��;-�áD��oL��,��<��S7B��"��:��@��)�v۹��ϳl�Z�bX�1�Nd�$x��@��� 䊐x��1 ��ʪ��lj5�9�����|񆎝B�G	�F1������%T�1���=�WG�&�))H��~���l��>1#U8�z'u�7K$�!�S}�P���~6^}���b����$ ���E<
�$�[*��7@K�zxq"@�K,��������#�:�) �4ocf�K��/��CA���ߤ�[u��`sZΐ�sZ�mm [\[:X�ݳ[۴p�>���嚺���p�&tO4��U��"D��@��2�>�ۗˢ��$tt4�t�CZ��T�v�!`՛Nv����m�*��E�uf�,4l�śd��78uڶ`]�6���F,�G�2�5;nN{Z�z� % "g��{v{e�T����-�z�v@8���gQk��\���7O\Ð�7]Y���nv�l�r�3r�mk��O]T�[�:���y��VyX�8u.}$� ��4�y�	����v�!���5'sn�%���Z��;<���G&�[����=�R`�����dewk=Vw]������ѱ��sYx{i���i+����A�`l���@V��u�F����8s�L.H�h�kZ���_]N;y��P�L�q�]�9uL�v�pr.��rB��\t$I��t�-miX�Ɠ6�e;jx�n�#�p�w��J:�4-HU�+v��{e�t��=������b��Kv�b�	�*Nܝ����pR;��V_M�6�mA�N���{�����G�lMoŕ����]`P�B�t���Rʅ<�ͪ�x9vB_eNwd��v�8x8�8y��!�u�SizŃmN�QT&��Ȇf���*�d�m:#b�,bv�ݤ�.����^��M��i��w���<O�أD@ `#&.����U�qdMD�k_*w:ʶi�ۀY�( .mAJ��E�j���� so>�
�l;W��Z��KO$�) Z�fT��T�dͷ��2:��pq�\*�ɂ�4aSz۞��v�KsL���i{i��ރ\V�剺�r���v&��HGF�\@2ѥ�D����n�v�[\�F����8�.�oi�;hݩ.�Νq娤ZU�Y�S=��'Gj�ŷ;s�K��@=�[�5��@S$g�����d&��66㌎��z6:V��� .����5���kZ���jC.�.��
(48���(W�*`�H*l^�=����*�"hE>^6q B�����@��p��I�Ѷ��vù�ô�莟#֒Y�uA�6�cl�Ξ58��֭�6d�n9M� 5nN-����}���K��ܗ�{g�`냓���v�`˪֩��9x��6춵��¹v�6Rc��u����Gl)rqʮ���px[c$�HgTd^v���+���V�,����YMԑٔ�9PxM�Tї2���ɭdeּ
����9��2	�g��sێmf8]�t�lv�k�=�������z����w���B���fT�vh7���^s�z[uДrK�o_�J�USXT��.�j������pKn��v�ͼY�
rJ��ٙ�Ud�Ywh��UW8�wV��S@�s@�_j�?u��s	�F�7j���TO�sL��,�W��j�u�y��?7�8�<pK����n�׎Zܓ9�@ve;��]�Λ��%�
��m�a%㭸�߆�!�"��>����D|)�ܐC�b@�%�|��hrL@|���\��'��HRyn�Ժ�ֵ֬d�j�I��{7~P;��ȧj��9����rN���f�u���,n�bs$y#��z��D�*G���n�� %��� �%�^��<m$�����f��o���mz�f|�}�4�,���Ѭq
!�7i�똀�r�3��|_���#o�}��}���׮����$����ayv�P�t�j���YV����'�&�bĩ���=-��??[06�t%
:!|������?��I��F�71���?_[3�"!L�wq`|��Kn��&M���s8%�m�@���4�v��!ҐB¯�z�rf�9^��e4�k.H"I��L�Z���ow� ����?7l��Q�+�{�h-��&%�"8�N=�I�ܪ＼|��� ��Bfo�g�S�.x�[���Nvf�B0G	��K�Ҳgj����r9�n����|�� ㊐����>����@��l���� D��;{w7�|������ŀ~��3�B��S���J��nQWwv�O������ʫݷ���nh�U��F��,Iǡ��%��� �]�y����Q�P�W���*H$c�O��0��� A#�� @dB1�V��4<��v���& �����$�<�'�~@��s����w�N��F�kZ˭�Ҳ�6�G�@8����;w4�e�Y���0Nc��$�I����M�������E��y��#\{)�����3sY��Y��|�����T��vS@9�˓"NH�cȔs4�v��
dz��~�z`^��<��T�H�pQěq������M?�����*���/;�f5�̒d��4?�^�ր��T����A��==� �{1��Q�r-��s@��k�;{훒s����[�>V"I%�y$�{<�g��-�܃��ge�I43�T���Y2,���rd��y6�=s�*Jj��v����l;#N.\��9S���]=s�Q��jA	w"�u���Uf̝����>�2"n��I��lE躩%�X(9���Oq�����:��8V�g����:m �$)�f��s�u[n��.B��Ύ���iNFx}q,�֡��ȧ���_�9�庥��Վ�Ko8�r��4^��u�<ݸ&�]we�$p��I��PkB�$�(]�z��,����D$����Xv��bqE���ı'��۹�~�h�����:��I%G���WE�Ю�Y����s?~��*C�.ݹz�*@7F�/0� //C��s�V�R���@����?qڴ��˒$��s7V���:�6""�����vp�����Lz�i��ǋ#mC$$�V���Q���X�؄c��n˂6���y�^�ntZenf�� >�IhU����w���w�Ѭ���I2G�I��;뽯��V����K��k s�:�<��g$�:P>Ӫ��B���˰�7m�����똀q�H�v����kB�$�4?�3!.��oz���X啕�<��`�+���ۍ<Kq������v{���ۚ;^�ߕʒ.G���dy��eFݎ���<)�5��8׶0��l>6P-�z�qI1�Hds �s4�v���s@��k�ߐ__nh���N"db.�6�8�~��9ʻ��@OO*@}�j�}�}�Aܾg�D��	"Q��;{�ٹ'}�l܂$��荒�M�h�R $"�4H؀��U|��}�s�s����h� ;Mŷ�ٶV{�V�n qR�䖀q�H=��f.��=���o�X��&H�1�rK@~������@8�p�����l�r]�.��x�>���X���֭(�ܴɄ���ۧ�N8�T����@8�}aמ��'�����X�X9$��qs��>�#�����ՠv�վH�|�n&�Rcn4���n '�� >�Ih1�@vۘ���Z���I�C�f���ՠv���I�����蜔�T����ګ�g��'�L��L���4k%���@9�Z�r�����'��H�$�~~~+��T��*��Ʃ�ܒ,]S�W��	d�k�'Ijt��NlaՖ�e�q'"�8�k�;m��9�j�;]�@�vƩ���y�@�s@��@�v� �m����;1�nd�$u��H��@9�Z �I�$T�>�ê��
�I��*J��][��8��ͼX	)n�� طjb�	�W$ܕw7s��w�j����n���'}��ܓ��P���,���BI�d�ՙ&���50�\��K`{C2��ݭWM�5۫d�����5;@���Ғrȵ��n�������7`:m*�Ӗ^�'N9���Wve�ܭ��G��67me����x�Z%�Y{�����p7@u�ܨ	-�v4���]�Bқ��A��ggm��L^v[Ԥ�&��Z�\V��u�3�-���+�Xj�b��!y7���{�ww~p�A�C|�}r��Xf��&�Kl���Q{&(�q[ό�9Pώ8}<n��ٸqjrȚII'@��s@�_j�;]��g�=�M���rbY$2IiI�z�VrJd{[��n��m��P�O��521	'�|����@�s@�_j����$��!�Iȴ�&��R�r�z�s��Z����"#��$�on�޾ՠv�ՠ��@?pK(��G`�������:;[e���v�@�Àqq=������Z��i�ds$xԙ�]��;_j��٠v��h9ڛDń(�,FkWrN�;�6�F(�=z#�\����KP�*@7�Z�vFW���z%�"4��E���4���?�J�|��|�ݸ]�ŒD7"bD�h8� �9h1�A��������@z�ީ��j�]�����X�^s�t(J�������� ԡN�I�fԪDN��m%n�l.�c��1��Z�ť�Ӌ�GU7�(b�fj�u=�������{�{�����q�H��@�2Y�'#BCȓ�h�l�}�$__nh����~A|ܾ�x���LprM@8��Ɉ�W9���.�r���|r�F`M��B1�(���
��F�$X�ȑ�
�[ @�mC!�#��9�4^1� )
��G�>��14�~u��QOr�F�U�}����,��R#_��@	�,fp��a�HD�O�/6�RD��D^.�^]�І kpJ@�R�<V�9�	äJA��v�4S>�(|@�X�@�`BN�����r�P�c��޹H��z�U�,`H�`��18���D�S§�1~����~��
t8(��8*�j�QH�����������;1�9�L�cRf���!V��z�� >~w�y���s�m�x�X�9"�;_j�=U\�'��'�� >y%�>��,���ܗ��]���ˢM.�q�N��q��$���u�An��9� �GͶ��~}�`q�H�I~�r�����@7(�*8�r&$I&��n��}����Z����s���>H���Ԙ�c���ͤf{րs���qR�C�tj5dbR-f|������[�w������>�	0 ���ꘚ��kwrI��d�K��Yvem�n� �sP8���- �:��e_� m�HDЄ�J��j�^1\�q���w ;�<�� z ۳�w�p��F����8䓀{��ۚ�V���V�s��@�{�f4�1I�LjL�?u�9��S#�{8���?<Y����i�ژ���ő��|s��J&^�ŀ|�vp|&�b�	�W%��]���t)�7��={� ��np5G/�~��-����iq��LH�M q�@~��;7޿����@nj�G��N0<�SL(%BU(�ҍ{�{�|㭾��;F�1ڇ�j3:�����WE�����Q�����X�eMϢ#=��m]tm�\'[N��|[U��4n����6,�sc`8n�h�㪍o\��u���t�P����nwf*Ƿm׳żU��숓�A&��q����%Y9Q�mk��q�Z�k���#���ku�=��6ݸ�ܱ�ͼ���(`�e5tf�l��UxDMbo����V&v����=��sf�Iwٹ���$�cp�³��5�ɤ��!����t�'� �9h���UU��==���fMA�L�B$�@�}�@;{f�v������ă�|�d�r4$<�9' �� ��9%3)(u�k�i���X�QI��I4<����*���ڴ��h�cX�Ʊ��EwrU]����RK�{7���׀��@��v�I�$�c���'X�v�h��Ɯh�U�^ú�������i��B��D���=��� ����?��>������@�3�k��KDi9�rI���o�:M� �� ș�[@���Ǆ ����u�'o�����h�ҼD�8�7"`��@�P�& �- v9�dp��bN8�6(ܚ����U��z����r��䯽�s��g�Pq#���2K@~�U�Oo�����1��{�ퟻX�Q�hGE>ήuҺN-��o��Hr������Y�w���3��ls�w������$��� �-��ȅ���8�@;m�U�zk�hol���zƱ�cX��&K�*��:��:np�+K�	%"JC�g�} �l��٠�J�S�4Ab�܏C�b������������3���8��r)�v���P�����:��:np+�=��=[��/����&m���L�u��>�^�ay�nm�X������5�d�#�n�����$�- �IhG5 콣Rc���rh�վ��H�{���o <ۼ艓�U,�*l����%��� ��g �9(������Z�-u�$�Hyr- ���ͻ��9���/���)P���]Pȇ��<2���"����Sa�U����w$������(̄�0�I&�v�4�>�����ݜ o����>kM�?Z)ML�\�d�RQ�ӻ/<���� ���{t��v�#d�9���&5���d@�������;]�@󾈅�@z���{3S7�jK%M���s�#���Pc���r�Qvn���lԒMT�`�ր:�h�]�:�����ͭ�7`��@;m���h�ա�>�K޾�G���ƚR
1F��$�- �IhG5 9&�*��W9]�����������H�g�ݜ#���� ��]�Xԭv�h��Lї�^s��Y���k�9����y�-�.�[/u�÷�pV��N���^M̥��>֤��5��sl�㛖wn΍����	�p����adn8�0�t�����Bz��O�e����eb	=n��h]��"�Ay����Έ҅�ny�ݜ;=L�M)��vE]/nYs&6%xl��w{ܚ��m���,k����k7c���W�,t�x� ������؍q�+�}��.O���κ�ƒ����� H����ԭ\�'$BCȓ�hyl��٠r�ՠv�վ���H�v�߰Q5�na$�M ���+�Zff%|^�����U;U*��WU%U�QДS�ޜz�� =�w�~w���M)�ȇ�X�NE�v�ՠ�@;{f���V����g}�P��0Q3v6k<��э���tnP�װ$�����.���4f��o5�NE"������٠r�ՠv�ՠ�EDL����h.�� <��_BP�D�F�Q�f�����-�������dq)Q�swP���-�ʻ���@�ڀ���L���KWD�Sw8
!rQ[ٽ8�� ��>u�8�n�����-L��f�� ���`�!V����ޜμ� �
<�٢�T�MUJ��Nru�7g�-���F#v����K�z�vݷe�{0�<I�"Md�G$�����9_j�;_j�:�k�?^Ʊٍcrdmɠr�տ��ؑ|W}���@;�RiO�D<�łr-����v��f�M� 6�� `1 ��J��1 `b��C��UUu�}���� �S��1xhnWsW8���^ݬ z���y���V�^T��dq�RG����jIrP�7��7�zpO��薞��m��`�c[ Y�u7�r���ca�[r��!]V�r���f9h�r��&z�\�÷=�@u�\~��&F&�N-�}���"���@���9_j�}���{=潒&�&$L�9�W}�~]����ىw��h��h�v;"Md�G#�@��nnI�g}w$���]ɳ��,��%*�`��PJX�b`b�S0��C "�T�$ �V4��� �����'���?Lk��#bN=�}�@�_j�:���˶���,"�Y1A���wCux�m��x��A��]M�B��aܴɄ�T&��dMX�NE�s��h\�z��u��~��i���b��&h�]���h�1�g�v罈�9h�r��}�|�����ۍH��=��؀�c����s�v�OZ[���9��ȚR��=}����;]��;_j���Ͼ\w�z.�	cq�#��ʹ^9h�5��1 �9h&"S�����%6�^0�æ�BP�0b�湆��8�e��$�4)���#3�j�=�FH@I�&�Z�I�� P ŋ��m@�����`|n�2���BJm~�'Nؒ�6�BS�F��R^���?N#	 &|��@�H��
hJ�8!��	�blP�=A�"&��K��0V�[4�$S,��H�"�"c �#s�>Ut� B�f�0a	;�"�|`rj��G�>>���U�����?:����q�7y�ϟ�>�U���UUUԂA p�`kX��7cu˺����ru��Z�T- u�����X�e�h!vL���`�ٱ���[��K:n�]�u �ʼ�P��g"j�a�7R�:x���+��P��А4Y��9��cA��n�p�lk�Dv]��l[Q4.+v{xf�"Hlg*WS��8����r��/7 �^{Blcd6��Ů��q�a�{vrZ�ᗪڞ�;;�m�086J�:s�n9�Z�!��溕z��'�uA��]���zq�n8��Ņ^���d��M�
�B�1��,a����Kq ��D&���Xzp��b�N�-1�5;$�[UW�d%L�jv�T�����؇hS<�R�[��=#�]�����q�,c �F�/hbv���Ɇ䘎&�7�������u�$&�gE�74crk�ǮmQ&؎VɎp��%yN���KF�v-v�f��.�2�n-�t�^���r۝�]Q��H�Z�H������*��q�}*�k�vp+�� Z5m�-i\�a,��{2ܻm;<�-ST����@W�-�Mq�6ѳ�v47;��@V<��C��d�&VT+��z1͇�0@���^��*����G�ny��Q."�C�u9C#���h�v]�s�ݣ[��*Ԏ��aV�L�鴏\�qf5�H�	����vm�`��ڥ� 0���c��Q���;���#�6�D#� �˻!��=p�e�c�*Jdٲ�ճR�v^��8l�L[b�F-N$)���S0�m���o%k�rΈ"�ӷ$�mqv����s�q� �Sv��&�4K8� [A�昽V��娝�^zg1�]`�h����s'F֤3M]�d	�U�S�,q�#�v�z�X��u���gYD���Ğ�t/-!*��%��(�5�秱,jcv�lx-�s��'��x8��vx�0.���ݙ�¶�r�ù,�e8�WCmC ���ݴ�(����4y��5�^����(xwA����#@�P�A0�/���p��a:��õٺbStup��i�7"hˤP��D]�k���Wi���'Dgv�TZ�zYts��lk�nBL�.1�x�9#�n����V}�3���KD���8��:9k��Ҧa�s��g��)�[e㑇[v�`���z8M�rt�:u �<.Թ|s�v��7���)),/Z}�@hx�u�9TMi�=���5�3-��Z��\�PSq�ffd�aP^ָ������ݞ���X�l���6z�]��[��{t��ЗH�5�4}�o}�x��u�yל�D.P�_P=���._G���md�I�@;m�k�Zk�hol�fgؑ��7����I2F�$�/���;]�O������r�1O�D���Zk�h����w�.J7m���ء=d�1��@-��g٘������Ɓ��Z���B��m�Dc�F�����G7`QVθIfZ��Ɖ˹y۞O�jl9%��2��EYWwEԓWw��u�7l�<��J?H�� �׵3u16�1F(ܚ-��ϳ�}��;]�@;�f�v�7�>� ��W�,r5211����@;�f�v�4[)����nH���'"��٠����h{�W��Z3ޏ�$�iYUh���� �n�P�۹�����{l������М��<`u�v�����s�=b��p8��Տl������s�cX��&H�䟀�<h�ՠ~]�J����ۺMq*�l�13V �-��1 9&�{������bL�Fcr'���y�m�N���&�qB b83#���k�Z��R��Ƣ��9E��(�J�{�xn��<��ԣ�W��� �;z�n�MT�a75w�6�2K@}rL@I���ɋ�9��mjε`��ǋ5у������{�S��c��Ǳ����K�j��kvp�۬ �n��n����{#M�,�r-���}����4l�v�V�$s=���J&��%nn� ��� �� �-��1��5��i�̑��4���k�p�۬��I~^QQ�%~�s�� =���#b�b�'�����4��h�e4gz��ۊ8�����|��[R�Y���]7C�o	�>\�n��-���2a��8h�l�v٠w������4w�K��E#�h�=��&�ܮU�{րs�� v9�ԣ����Q7V�j�	���]wN���P�d��� �ݼ "]9&��S##qh{�������v١��^�yh0��F�� Y2F�4���
"|�o����y�0	��������������@���=:��b�o�{�͸~u�P�cU�.��K5uYxnچ�ZzGZ��niF�,F۲&.vݭ�V�j�sy�O�gr�O
lٸ�|�Dyx�zޕNGG&��*�S�Mn; {n\�J)���\�k2�5�m�/�k�pΰ>�)gL�c�.x�n[ �lf5��sǇ�H%�����9"u%�b	Ԭ�Cw;�����:ףn�tpb�jІ;L��j��B�ڶ��<�#�˲�<E&lY���`4�ݫ-~m���ڀo$�\�>���@v{r�=��$�̍��4�ڴv�h-�@9�f��gؐ__$ҟ,��%��ȴ=�c���c���#�z��!�{d�3$p�^٠�@��C˷��@����i1��p�M�@rj���s`�;$��s���󾟯�k�(NK�:��랚�%�
1�(�J%v�YaY׎��U�HM������_��v�h-�����zh���R69�����v�l�Z��E��0_i���Y����v� ��n\�NF�*WuWf |ۼ ����Un�t�����9���D�A���rh;n��-�6�M@|���d2�'26�$�;�j�9�)��� �m���T�1�RF�&'�`�Ó��+��C�L ��;���m<�;c=��"��pH����Z;e4�٠�@�]�@�L��=�2a��8h,��:��r*@u͂�们�(H�	$�v٠w��h�L��d� �|A��9�,��~��@8�dndR|8
,�@7"�\� �5 uɨ<u	�I���I�;e4�٠�@�m��8��Ђ��$;9���9�<�rzv�����AO"���ņ���;�����ǒ7!������4������2�5`�1�naR= ���yt%T7��=�0�z�������5�Ʊ��1�9&�{���'�K�׽v��bX�%ｭD�Kı/}�kiȖ%�b^�ڙ�VI��K������bY��V��~�����r%�bX�����q,KĽ����"X�ǈH�Dh�*E> Cב,��bn%�bX��=��jܚ&����]�"X�%�{�kQ7ı,K�{��r%�bX����Mı,K�׽v��bX�'�z��FgQ��0`��^���]n���xt�.�uZy�\6݃ﻼ��|7;)�Si6��Ȗ%�b_~��[ND�,K��ى��%�bw������DȖ%�/v셄)!I
HR�^���Z����.�k[ND�,K��ى��%�bw���ӑ,KĽ�����bX�%��m9�*dK��/��[��K����֌Mı,Kߵ���r%�bX����q,KĽ����"X�%���l��Kĺ�����ə�[%0չ�]�>��3*dK���U72�D̩������Tș�2'���172�@��Mj��s����2�D~%B��Z�f��|��=��-L��m>��D̩�=5�ى���2&eN�~��}�L��S"\�������2&eN��0M���̺ɭK������RH{N����	�t:������t�Q�jv���{L�B$�����[�v��0���X=w0��\u����s�8S5]���CE�V���;``��w2���U�M��^wm��h8,F�zWp�]{�vK��^%�֓���y��m���㧃��RZ�ii����/f�@y�a�q��W3Yu������*�Y�ɜ�Q�Y��\�H��d�x�j�n����{t�6��ݞ�����;���L���~Os2�D�5�vbn&eL��S�߽v�}S"fTȗ=�f����~����
�aV�u�/��TB��TB�����-:�˒��Y����2&eN�~��}�L��S"\�������2&eL��m>��D̩�=5�ى���&������i���r4Ʉf7"qo��/��cu2%�ߵ�����2&eL��m>��G���{����_۳q3*dLʟ�;�!}�¢T¢T��ASTU�ue�Y��M�̩�3*g}�ki��2&eL��n�M�̩�3*w�����dLʙ罬�M�̩�3*wS���o���b����Os��{�������fTș��A�V������Oz�D̩�.k5Sq3*dLʙ�{��}�L��=��wu����b�]rێ�:��O<=���<	N��Lrg����^�xf�md�5,�֬��Lʙ2�}�z�>��D̩�.{��T�Lʙ2�w����}S"fTȞ�����Lʙ2�{�>�zr�ls�4|�����=���k5Sp�d O�!z���@jP�M���
���Lʙ�s��}�L��S"zk۳q3*dLʝ���������L���]�k
��4ǻ��)�w�Os����[O���3*dOM{vbn&eL��S�߽v�}S"fTȗ=�f�n&eL���/�k��!$��~�q}���� j'�ܳq3*dLʞ��߮��dLʙ罬�M�̩�3*g}�ki��2&eL�}�jܶh�k%��k5f&�fTș�;���i��2&eL�s��j��fTș�3������2�D�׷f&�fTș�?w����|C�؍d�����ю�G�Սr���2b���lu;�H��Z�{�?*dLʙ����T�Lʙ2�}�|m>��D̩�=5�ى���2&eNݵo��/��ck�g���Cƛ$���[sY����S"fT��Tș�2'���172�D̩�o޻O���3*dK���U72�D̩�Ow�ռV��m�W|�����=��}K�T�Lʙ2�}�z�>��F!��#5����'��[���
�Z��+)-��J�D!)�j��	$�B@ċhk��$d�.1�h8ち��	�y��:uIa+�:f�d�pHt7I�d�P�8<cQ�$C`a�H��Ү�A���$F$d!��07����K��B$a �!��� 0�����%�R�B���ͤ6�J��6�*��D`�xR)J�#	�1�'y]HB��]��=�m��ވ�UR���c:�=R��ʃ�DWƈ�?EN	�(�MĹﵚ����2&eN����s�=�{��y�x~��]c#���ٕ2&eN�~��}�L��S"f{�֪n&eL��S���6�}S"fTȞ��i��}����ck�ͮ㐑�<�f�v�}S"fTș�������S"fT��Tș�2'�u츛��S"fT��]��Tș�2'��d�s/3D�ӝ��C�\�8���F�ۉ�0t�:n۶츳/���(�e�j�w�&eL��S߿~��}�L��S"zk^�q3*dLʝ���� ����fTș��kZ����2&eO���a��!����5�W4m>��D̩�=5�[����2&eN�~��}�L��S"f{�֪n&eL��S���6�}S"fTș�z5��X۞�����{��S�����i��2&eL���kZ����2&eN����}�L��S"zk^�q?H��}��-3��o�� �1��~��X�u��;�ߵ�7ı,O~���ӑ,K�﮽*n%�`e�QE,i���|�Ϣg����r%�oq�����g�sD��w���ŉbw���"X�%��#���ND�,Kߵ���r%�bX��{Yq,K��g�K}�X\��F�������ș�gLR�7�r��T����������]Bf�ԺѴ�Kı;�J��bX�'}�z�9ı,N罬���%�bw���"X�%��;��f��u��Բ�5*n%�bX�����?���,Og��ț�bX�'�~��iȖ%�bw�^�7��eL�ow��_��5���+G�w�{��7�����Yq,K���ND���"dO~��*n%�bX���߮ӑ,K=��>���Y�f������,N����Kı;=�LMı,K�׽v��bX�'s��D�Kı=�n��d3Z��f�j捧"X�%��]zT�Kİ��~���i�Kı=��l���%�bw���"X�%���;����i���V�4� "CRz���2a0��&J�i�m�r���{r`�'E�f��U�q�F�ZHp���ڸ-pU�HL	�[v�'��ɒ�NgPR��l�����G��o��o�>����^��;U��;q�����{#�¶N�A��ݙò��,�n��nF���r��-��Oc��sՓ0���HS�\Ͱ�y9��7"�Y�"U��7lc��m7{�{���mYu���5�mWo&����:�2x�'mfєT�vlmP!�g�Ɔ5���%�b}�^�v��bX�'}��q,K���ND�,K�����Kı;�x���)����3Z����Kı;�fț�bX�'}�p�r%�bX��צ&�X�%��k޻ND�,K���a��u�5�˓Vf�D�Kı;�{�ӑ,K����17ı,N�^��r%�bX���dMı,K�=�kV�ɭe�&jMK�ND�,�A��=?o���Kı=�_�]�"X�%��{6D�Kı;�{�ӑ,K����V\��tjY��LMı,K��}v��bX�'}��q,K���ND�,K������%�bS��̾�qȝ������y-�Z���;,�H�9��-I���2#��֧tsī=���7��bw�͑7ı,N����Kı;�J�r&D�,O~׿]�7���{��?~���\.�g����%�bX��}�i�j�h(D1 ��j%��]zT�Kı;�{�iȖ%�bw�͑7ı,Ow�y�e�Z�0�h��ND�,K������%�bw��ӑ, 0ș߿fț�bX�'�{��"X�{������z�m�%c��{��2X�����Kı;�fț�bX�'}�p�r%�bX��ץMı,K���o���jfc�5���r%�bX���dMı,K���6��bX�'}�����%�b}�o�iȖ%�����>̩^kF���0�u�(��:(�v�EEn�4�jl��P��f]Y��q,K�����"X�%��k=jn%�bX�w���~}"X�'�~͑7ı,N���kV�3Z�T��5.�m9ı,N�^Չ�~H�L�bw����9ı,O~��"n%�bX�����O��2%���<?�a$.���������ow�����r%�bX���dMı����#�:A�b����D�'��6��bX�'�kڱ7ı,K̕�Ik"ɊF�[�~>�}��gـdO~��"n%�bX����6��bX�'}�j��Kı>����K�q���Ϩk�t��j������,N��p�r%�bX����q,K����ӑ,K�｛"n%�g�����>���w��a��ra����݌ݒ޹�m����y��uԈ��VՏf�/)s��a�ѫ�8�D�,Kߵ�V&�X�%����]�"X�%��{6D�Kı;���iȖ%�b{����f����d0�kV&�X�%����]�!��DȖ'�~͑7ı,Ow��ND�,K�׵bn'�r�D�=�~l��Y����2e�]�"X�%��߳dMı,K�{�6��c�"{��j��Kı;�^�v��bX�%����$]6R�5���{��7��w����"X�%�����q,K����ӑ,KC�]� @N8e4)v�y��l���%������##$X8Rf����b>,N�^Չ��%�b}�w�iȖ%�bw�͑7ı,N��p�r%�c��w���&v�����nus:�M|�������sd�8�0�Y����S9q!�R�sV&�X�%����]�"X�%��{6D�Kı;���iȖ%�bw���Mı,K��_ֳ2����ff�ӑ,K�｛"n%�bX�����Kı;�{V&�X�%����]�"X�%�}�e�Z��CY��n�Z�q,K�����"X�%��kڱ7�� �ș����iȖ%�b{���q,K��޻�3/������iȖ%�bw���Mı,K�k��ND�,K��l���%��dOw�"X�%����jܶi�5�V�ֵbn%�bX�{]��r%�bX~�����,K��~��Kı;�{V&�X�%����Dn`y0�D�ل��WZ�3i���z͘콴�(�{CA�U�n��eq�Yق��cV���Ǚ1\�ut�ɍل7�g��vX�6��VH�Yͮ�8��:ݜ�We�nv@ל�����Jg�;Y6����n9z�Q���x{=v9�˻��N��n���Bj�.�+/R�F�;!�HC˓T�vrK=���/m:Ƹ�T�ޑ&7���㛳/+�r������w{���&��a��9�R��D�麫�$j�.sOF�z�N�P[�˚,�jfc�2�ӱ,K�����"n%�bX�~��}ı,O~��X�	șı;�^�v��bX��O��s�.�	s�������ŉ߽�NC�!��,O~��X��bX�'k߮ӑ,K�｛"n%�bX���}��њ5u��I�u�iȖ%�b^���Mı,K�k��ND�,K��l���%�bw�{�ӑ�{��7�����cX�5��7�ı>����Kı;�fț�bX�'~��m9ı,K�{Z�����������T��V>{���bX�'{u�Sq,K�����"X�%�~���&�X�%����]�#���n���m���Şա6Л��'��\�0g\^:M�n]�<��)3b�n�aN���Y��n���Sq,K�����"X�%��z{V&�X�%����]�"X�%���zT�Kı9�����j�kF�h�r%�bX�g��bn���U5Q,O{��ӑ,K����*n%�bX�����Oɕ3{����~�������F�|��{�K��~�ӑ,K��n�*n%�bX���iȖ%�b}��Չ��%�b{ޅl��ff��ɬ�ӑ,K��n�*n%�bX���iȖ%�b}��Չ��%��P���~�iȆ��oq���^Q"��리{�o%�b{���"X�%��z{V&�X�%�����r%�bX��ץMǍ�7������������ygRXr=U�A�L��a�ή�,+:���&�Z�����fjMK�O�X�%���?j��Kı=�{�ND�,K����� �$����M�$��\�j˅�[�R�fj�$D���q=ı;ۯJ��bX�'��p�r%�bX�g��bn%�bX��׳�5���5MWZ�m9ı,N��Ҧ�X�%����6��c�:AY O����H7��"�"�'�9�Oj��Kı=�w�iȖ%��}���1��-`�������ŉ���6��bX�'���X��bX�'��z�9İ?+2'�w�T�Kı;�]���C5s5�W4m9ı,O��ڱ7ı,?${�]��,K����J��bX�'��s�{���oq���~�S?2i��=t�c�d��3��Z���5�;�g����r`�i��B7&mz���{��7���׽v��bX�'{u�Sq,K��}�ND�,K����Mı,K��+e�34em�u���Kı;ۯJ��bX�'��p�r%�bX�{G�bn%�bX�g���r'�Aʙ���O��s�.��jǻ���bX����6��bX�'���X��bX�'��{6��bX�'{u�Sq,K��N�ښ����P�Rj]h�r%�bX�{G�bn%�bX�g���r%�bX��ץMı,�9�pX�t"���3�?o�ND�,K?^�b�B��������d�=�fӑ,K��n�*n%�bX���iȖ%�b}�Չ��%�w�����l�۠$H�@YDna�9�<㮸��[5�()�A�	;,F�S
]D�G\Z��fӑ,K��n�*n%�bX���ٴ�Kı>��j����DȖ%�����m9ı,K�߲�֭ˎ�5��k3R��X�%��｛ND�,K�h��Mı,K����ND�,K������%�b}�����j�kVkZ�ND�,K����Mı,K���6��bX�'{u�Sq,K��{�M�"X�%���ڷ-ՙ.f��L5��X��bX�'~�}v��bX�'{u�Sq,K�绿M�"X�%��z{V&�X�%������L�[r�j�9ı,N��Ҧ�X�%��k��ND�,K����Mı,K�k��ND�,K�Q8ڠC������ s��T��~�@#aQ�4hf�$<���� �9Cs�z��Zĳ�D^!�t�\H�`�7�3@�΀�$�1]!�DX�"�	=U�'�Oډ����U�k M0�J��	��@��D���gF>W۠9�z@��ϟDq�P�tDӈiw�b�(�6'�(`��ʒή!��3� �4��J�7�R�D��M���,h�0=�����o{�����@U���UT	$8� �`pn�ݝ̨�3aC\��w2-�Y-�pU��m��Kiv=�丞9D�#�GnM�A��[nl]��n���Q��Ŋ�Z�	��bv^V���y ��eWm���i��-��H�{m�Y��ʅ�-5ɧ>غSv#=�n;s�r<�[��]��l��f3X�w6x�Nv�B�`%m�m�Cr�О�h1����N�TG��c����K�sWa{e���U�����Qۓ�kd.��<�Ԭ�ؖNfjU�V5u�l��C��%�X���JK�c���ꈱ`h�;h:��t�Ӎ���ڬn4J�je?˪8>C���+k[ۥq��U�n�;��bWu]zZ�!���FRN�n�.�	�0��ʥ�Pp�m�.#�:��Nv�q�;Wv��bgmk��3iu���͕7L��5>C^d�/�Z6�ɮw[v�&-�;���S6����s����ҭ'Fȃ�\�qÞ���N�K��[^�l�|�^�~8���A�TX��e�۞�T��ۛ'f1�l���;4N�.M49] �/b��b�K+us�[�Pwu��@��m'�{;�vq�*Tգ�3�fu����N}�F��k]�hڙ9�v��b���D�`0�RńC�[�k�ˎN1ת�4���a�Wiݑ�t��v��ֶ,�gȋ�:�mʷ2K���Z�j�m4e�j���%�*�x&2q;5�&��B��V�%��IfƐ�]��y
�Ŷ2L�X�@��r�,kE/ĸ�ɎLp�����.�?|*��s�O7��qdW�Fh��sӻNs����^�:i�.{\& MP��`��N�쭔�m�	�n�f�S��O4�&�Y~�>���n��u����ŷ��E͍�]/7e'����J�K�r��Vz��+��8h�6UL%�+�Uv+\"�M�󕭱��I��۬s���'���b՝��i�mm1��ܺ�{��pz�҄H�)�U ?` T�>�D��VxXނ�C�6�ʁ�<�x }���n[�d���SV���J��D�j�A,��iu���sl.��r�t�>�p6�ל�����ӷ]����G�����~���@퇎ݛ.+n74�&P`�u=��e��f�ș��v�c����y|�cv�m��&�x�[���uz�u�JۡvLӥ��XM5t�L�G�ᡠb�Ǜ]��յeF��k���v���v뵥�k).�.a)�5�d�Z�&*��9����|��4�L4�[k�x�v	86b4�-=���ag�۰i)�9�ա�kZ�?D�,K����iȖ%�b}��Չ��%�bw�w�iȖ%�bw�^�7ı,Od�|f�Yn��Rf��6��bX�'���X��bX�'3��m9ı,N��Ҧ�X�%���~�ND�2�D�/��\�����d�5,�f�Mı,K���fӑ,K��n�*n%��Dȟ{��6��bI
H^�6䅄)!I
H^lɧE��^�[��W5��r%�bX��ץMı,K���6��bX�'���X��bX�'3��m9ı,K��)�jܸ�3Y-ֳ5*n%�bX��w��Kİ��Ǻ�?j��Kı>�{�m9ı,N��Ҧ�X�%�Ν�����<�<����͓C�e�c�{]���G�O1�i ���S(�,����Nk|�Ȗ%�b_O{Yq,K��w�ͧ"X�%��]zT�Kı9���~����oq��/�8�pԻ-�17ı,Ng{��rp ~k��� bUJ�zP^
��bj%���[�7ı,N���6��bX�'����7� �S"X���Y/���[d�k6��bX�'��_�Mı,K���6��bX�'����7ı,Ng{��r!����}��\�K�BUX�|�,K?�����iȖ%�b~���dMı,K���6��bX�D�����>�}���V[�s�7J�I��Kı=������%�bs;�fӑ,K����*n%�bX��w��Kı=��!��Ժ��sY�nJ���`��G%��9�8˄N��k��y�=��eѬ�tj[�dMı,K���6��bX�'�u�Sq,K��{�M��g�2%�b~���dMı,x��Ͽ��'�PUp��������ŉ�]zT�?�r&D�>���m9ı,O�~�����%�bs;�fӓ���wr{��7�����K������7ı,O����ND�,K�{�ț�c����5Ps��@�b�H�:��PK��o�m9ı,N���*n%�bX����f{2���0�k%֦ӑ,K����&�X�%���}�ND�,K޺����%�bs�ߦӑ,K��/��[8f�i�������d�w�ͧ"X�%��?�]��9ı,O����ND�,K�{�ț�bY�7���~Ｎ���9n6./6�����v�8u�ݮ�+��e��@;c��S���ϝi���f��O�X�%�����Sq,K��{�M�"X�%�}=�dMı,K���6��bX�%��ٓ&k.�jMd�5�kR��X�%���~�NC��L�b_���dMı,K���fӑ,K����*n%�bX�����9��3P�Rf��6��bX�%����7ı,Ng{��r%��ș��Ҧ�X�%�����iȖ%�b_�3٫35�]��3Yq,K?���>׽�6��bX�'�߳dMı,K���6��bX1\�T�)ҩA��sq=���"n%�bX��l���Z�Z�	���fӑ,K����"n%�bX!��~�O�X�%��ߵ�7ı,Ng{��r%�bX��v�_e��d��5fMf��Ɂೢ�k�m��0t�:[��HC/�����hˎ�5��kZ�q,K��{�M�"X�%��=�dMı,K���6��bX�'�}���X�%�Ͻ�������Nk|�7���{�����k"n���,O����ND�,K���eMı,K���6���Q��w�~ߤ�F�k������bX�g��6��bX�'�}���X� �ș�{�ӑ,K�����ț�bX�'{�VK���[d�k6��bX�'�}���X�%���~�ND�,K�{�ț�bX�'3��m����oq��߯��d���]Sp��bX�';��m9ı,?�?�~���Ȗ%�b}����r%�bX���dMı,K�!P��M__0���ㄦ�u�Oj�9�sͷh��y�k�lp�	�yH�;Wm5�86xK��\�[�1�������N(
Ef;k��v���ꍇ^l��sqeK/�GAv�-�v��;9DL���9�*�7il��<v�k'.��&�,�IE��m����nM�^�XzP�Sc�.;h���&�SNs���c�V�s��e��]k�(��e�9-sspm����u�S*�G\p�4v���y4��Nۑ6v{WM�ԙI��Ȗ%�b~���dMı,K���6��bX�'���q,K��{�M�"X�%�|{��Y����Զ�ț�bX�'3��m9�?º���'���l���%�bw���M�"X�%��=�dM��Qʙ����g.]kR�Z��5�5��r%�bX��~͑7ı,Nw���r%�bX����D�Kı9��iȖ%�b_�즲hˎ�5��kZ�q,K��{�M�"X�%��=�dMı,K���6��bX�U�������q,K�￷�̿�)�p��Y3Z�ND�,K�g�q7ı,Ng{��r%�bX���ʛ�bX�';��m9ı,K�6;};�6����]X�z�v4�0��Wf�gxƝ�Y��e�,�����vס�X&�q7ı,Ng{��r%�bX���ʛ�bX�';��m9ı,Oe����Kı;�K!%�Mf���f��ND�,K޾�Sq����wq,M���6��bX�'��뉸�%�bs;�fӑ,Kľ��vs%յ�曏w��7���{���ߦӑ,K��Y�\Mı�@!�2'��~ͧ"X�%�������X�%���w<f��&f���5u���K��D��?~���bX�'��~ͧ"X�%��]zT�Kı9�wٴ�K=���}�f�����w��"X�'3��6��bX���~��*r%�bX�g}�6��bX�'��}�7���{��;���S�ȝ��y�]��l��v�S�\�)�z5����eg^�0�	�*�Oi~{���oq���}�_q�q,K��}�fӑ,K��Y�\��_�j%�bw=��6���*dK>���:��1��ǻ���oq��g}�6��bX�'��z�n%�bX�ϻ��r%�bX��ץMı,K�{yL��Ըau�ֳY��Kı=�{�q,K��}�fӑ,O��ԧ���$�Wl�8��
�|8��(x!螉�n��7ı,N���r%��{������.^�N�ճZ���{��'	Q}������$)!n��0�Kı=�wٴ�Kı=0��&�X�%���,���5.�f6�sWiȖ%�b{�^�7ı,Og{��r%�bX4�}�Mı,K�k޻Noq�������_��έ���]�+qSv��HYuu���-P�8C�4�jm������*�m]�!j��Ʌ��$)!Ii���Ȗ%�`ӽ�i7ı,O}�z�?��L�bX��u�T�Kı?{S��s�A7�7{�~>�}���Q�q,K�����ӑ,K����*n%�bX���ٴ�Kı/�a}�֦�S�����q7ı,N����r%�bX��ץMı�a�2'���fӑ,K��0���n%�bX�����kY.��)�ՙ��ND�,�X��Ҧ�X�%����ٴ�Kı=0��&�X��	Ң~v3H:�3N�-K �eC�!��dO���M�"X�%�}��㮸t�[��oq���~1�\��U�w3*K@8����������d�Ň�m�gN��v3vN��C����>rrg���a�X�z$�z������ze{րq�͂�r��%q�dm��$Zoe4۰@;�b[$�ꪻ#�aA~U����I��z�nhW��p�h���S8���c�C@⽯ s��=�`l$�DN��0m���PJqǠU�ՠz�������K�����|BK���w4��痵ڰ�0�Ny+ds���t�6��ud�,�=����)D�'��w:vuE����>Q���s�d�L#�������△"��ڕf���/[�m)���+���Iy��]m(�dSs�շ�R'n��{BnnЧW9=��zyul�6CD�6v�`��q��Z��JM�;�cY���fdq�t�-ۮ��36�e�SZ��Y~G�Cʎ��K��n\�1��ų�v����igx�k����'�H�{v��^*����\�?ͷ�� #�n9��Ϭ=p���=b[#��Ǆm8h�S}�V��T�����ՠ��˓��$�p@vۘ���-��-� ;٭c�cy���#�*�j�?uڴ�j���|����=�D��k#l�3tݴ�$�y%�;m�@Kd������o�jH�i��'��`�%�s���7Ks���5�)����k��-B�cp��!&�_��@?.s�@8w��}��w��jd�A1����ٽ�W�F@�_�O� ��O]�z�:�Z�o��#�����2&���@򧼴�v��ڴ��h�qY$RG�䉱�-����ڴ��h{3��Oyh�	Odb�<X����z�Z�[4
�Z�Wڴ��PY�bDxȤj0#	��g��Y�;�x���"�\�b�n�aqհg�!'��w���������ڴrƱ��j	��$�@���@��-� ;m�@|���Y����ڼ��v�<��͂qҮV�2�Bw'S�:b�D�x"{�(��p�oC�Sh�(�!	�
јgT$!�0�(�A���Н!�w�����e���e;���K�S��U�$Ta���417)�{��;{��������u�A4�cEbt�>
� F1��Ɓ���5>�ɍɸO��p|r1$��8}�,�����'��ӡ�r6hƀp��� |�G#�������w����<�� #��u^�ĸ�Q��~�|?+-�=C{(�*y��CB�ЂUO�"��%"��]�}�p
��P�0��"	P꡷b��v(p���x�V�\����]/��{q!{Q��m�N-��sL��� ��s��)��������jd�0��s4.��[$��$�r*@|̓l6��ݵ��N����{4�A��a92�p%�]f�쬰�덬6�׋�,�3�m���~� ��np��lB���Hz[��[�k�D�x�H�"�?uڴ�w4.������ؑ��%=��䘲ay�����@�j[$�f9h�V,�'�Q	8�4��ht�l��g}w'�	�XAh������mH��BP��Ұ �F�X0� iGH�}���h��c�bdǊH7&�S$�f9h�� >ɨW}�e�o&�S�Lv-��+<�9m��Ohv��[���rv��\��҉r֣��{8�`�n�!DG��n���A�����6�I��{e7ٟ}
d�o �f��:��Jd5��7� L&9$4�ޚ]-Z+�Z��9�u�1
d�<N��A�r���� ��ր�l�M@-�d�H����"�9�ڴ�)�}>�φ� ԱC�R�D�E!T����o�n��Fֵ�5u����I=qbR	m��-��pX���s��-��م�����Ɵ*\�������7����r�p��o^�u��1n�:��3r�*u ����n|뵤̫v����{m�*{<n��^-�3�6�c�]{y��xwv�=C]j������=;d�m-���X���!��ɵ�u���K��D��'R[q�k74�����/w�|{�;����~�s��(Ӄn8�`��0"@���Eۗ���0��r�93�8���ʘ�����q�����h]�z]-_��+���s�b�dĞ"8��n{^�WKV���ՠ^�M���X��Ğ<R8�z�/����ՠ^YM���@�֗pyF�1���AŠ~�h�`��1-�Z�ՅY1-�ц6��/,����נUӵh��Z��Q�\L��"�jHbm�Ѷ:#���sg<���F�n�nVܔ��veaۖ#$	��$����נ^��Z�V�ye4[
��2I'1���/p�é���,��Wʍ9��}��@y�| ;m�@��������Š~�h�S@;�f�z�h�BR�jI&<�Fۋ@�� �&�#�r���?r�m��=�F���~ ����z�h��h�S@���gݹC��O	��Nrs۬���b��n����!gs=v�%h�tT�m�r4�x�I�����r�ՠ^YM �-���5��o����V�ye4��h�;V�ċۈ1�18�k�Š^YM	;����j��@>���(�x�p�U
=�}K�ηg ����ڐ&��[4ם�@�}�@���.XW�)�H�L�h�9h��?l����� }�P��m�}�������������ʘ�]]�^�`���a룲�r�xf�y�S��f9h	ٰ@�j<�- ���#RI�&���/,��w����j�9_j�q\YrbO��bR7 �&�;2��f9hٰ@w�qcj�����nM��j�9_jН���ܝ��$1XH@d$$X�^ �� ��G����nI�e���M�6Ɏ-����������o ���R����*��.������Qr��e��g1ѷ#q�qp�1\�;���O����a�8�{�nhyl�8�ڽ���Z{�&܉�(����@�j�-َZ�]��ٙ��G}�������G�`9&�����:��G�Wq�ʐ~��	Rb��2D�����9_j�;�w4��hT�ZxK�F��L#o6��*@�j�-َZ��#x�E@��:K�����-l-��Ø����\0OO�қf��Mn0dk�M��qgB�U���tc����ׂl�Z.u�����N��n�b���Ɨ�� �,k=ض3mu	�3�6�\�:�,�Ն�d;Oc�5����m������Bj5k��i�n0��c���f�1Ju����=��˸G�;-�٬3�mj�
�j�x����cv���hm�I�2j�.��"'�b��2e̿`)�����O`�Y0<v{]�xؘ�F�ݷae��YAq�\.�d
��v��s��;2��f9h� ;ٹu�q5<x�rh�;V���V��[���@�֗pyF��q�c�@��- �"� �&�;2���+(\�N(��@�-���٠r��Z+�Zyja���)��a$�욀��r���>r*@+�^�ߛ�?p~��ً���4:�:��7*�s����[�pk¹���][r��i�:uS�ї�� �T��;1�@|�U��9�}`^��@.{ؽ�$K���-���y�b-j�8�b�F����H�{P�9h�%����&9�m��ݷs@;�f��ӵh��h9�,�1'�n4��L��؀��@vc���ȩ ۋ.�/s.x���@��ڴWڴݷs@;�f����b�AaVxn��G���k����0�E�t6یiݵ����9'7F����A��j!���|���hyl�/])�Uۏ%g�(��qŠG"� �&�#�P@vc����1�6a0xL$�f�w���̦���� ��,>G��9�ܓ����9r�� ��E�4�2��r�ȩ |�� �J̗��E�G��}�@��s@?v٠?;L�:!DB����UQSR�.K�9�nK�ٍ�Sی=Nz�`ڛaӍ��ν�bխ��I�Ls�q~����ݶh�e4u�� �z�"�Ѹ�NI1 |���*�m!׎Z9 �{F�ǎ5��M�}�J�������+�j4��dի05O���^�, ����BHC�7�
�/�PA�sy�������N|$G�-��h�x���W���$���隚�����v˷@W3�����,\�;��+p�<�h7X�kɄ�L	#��_z #�A׎_��Xz{| ����6�dp�	���7ٙ���h����l��#���ד�qAc��!�̞�d� >s`�o!:;�F���6�Z��1w��\�y >�Ih��^ss7D�C@������;<{ˀU�(>�7$� _�� _�
 ��T _�� W�T Z� *��� *���/�DR"�0A��E"("�0X* �� �H� �H� ���QR�D��U����Q�(@ �@��B"�1P` D O�( 
�� � *�P j� ��@ U��@W�A _� � *��  ��� �� ���(+$�k"�e@��+0
 ?��d��.�P @�(       � P       .�	B%
��UPQT*� �@%BIR��  %AEP�!"QB  * (�)E )AE
�    ,   ��  ��  " H @ $A�  �@� �J ����� )��xp��n�| ;���J�ܛZX�gP�ކ9>��׋E�w�:�� (�*�۾ܯw�ןn��w��xxP 	 ���� Sw��e}��7w�Nx-��w�o� +�|�\���\�z�Ͼ���o}����I��   �    ��\�R�����|[��O�ޟ-g��rs�������}����k�{w����ޭ�Ž5x >�  �     4=/���mT��ꜚ�۽�s�/� nJ���-�Ͼ���0;�>�>�K�޽O����� ��7C��Ƕ����>�K����}����{ǻ�� ��'{=o�!��ޞ���W���  U 
 �,[高uӓN����\�/p>�7o��y=Ϸ+��t�� �C���@�0 �}��� �@0��!��Y�� ;� t�>���=}���ӓ�׀ ��   �T � ޥ2wj\Y%�+�'ץ�>��ǥ�n&��sە�<J  �

l� ^`      !�P��)EA@�  N��:b PD� �A@N�� 4�M�%R�  5?PLԕI�d�@<z�T@�M h�Ob�P�J� h�BT�ԩJ@  ��Ԕ�@�)�\O�������޹���Jb""�N��OW�p@\?� pU EO� � � U��*�����!?��D�����2�?۞sd���q�cB)� !V,2@�H!B�(�S�=�"z�f.�pj��x{��̈́cBB22�%>���V��X�`��X$T�b�M9*a�XƐ 00�1�o;��pHB+B��1�	�y�L�O}>��Hjt=�S�%B X�D_Pa�u,�`�"bLu#aR$�H7߆�p<�C��p24��h@� U��"�`C
���"�Qb^�|�!R�e#F#c�`�W<�2A�N�HR�xi)R�*i�.f̡ff��,�$�,JĠ��3�+$�Ȅi�/���s9��g�@�4����k8䎐1"@ �#��!NL���(F��ë���YbPcC!H)��%�#��C׌+�݈!W{�EYɻ�ej��#��"g�LY���H$)$d ���� x0!��CRPaaC�A��64�R6S"��4c�%�� RO!kB%0�.S�k4mX0�cD�aI!HU�$a@�ɤщ$ֻ,U(��J��3�NpKpt8�IH@��\��H�1�������s�:/�|��>ISG��.HK�sd�8�ԅ��b�	y�l��}��p��!$#{7<�5��:s��! \u!CH􎩍)�*D,�BE,+P�D(S�&�W*k��-j�}����L���!!����<��c�2�ÛI���������):�Wjza찁��dd����	�@��-#Ж|�rI2ذ�dM<!cB1�`��a��qԦ2�4���ao<���I�w�=9�B�r�!LvS%:�#��<>p����i�HF��x��M���<M��sL����蛜�C�čGa$ ����\&����Ą�	� F$*Hdi��K�����VZB��B�L�ad�< ��=�s��J�.B�$�/���Z�X	���+��hD�
�*�+$�E�,H���t���M�y�!���7��#b���Y ��@�!D��%��CF�)�z���4S�Ac�5"�!!��')m���H�sT�,HY-&Jli����2R
N�П1&�xf�3OBH0Y\��)KϮ��v�����W4����H�a��k��z]w#��T��JP�0��䙜����ϼ��>+��a0��$b{>���y�;sy_!<=)L}d�XV]��/�$*B�,��ϻ>��=�p��$�"0X,��B$� 5"Q0cbX���B4	B,���ܑ5�������'=�fL���t�L���	��,�)�
K���|e3���� ��G�4!	w�9�4�>c$j�(īD�jHe�B
d�&�h�?Jf������3�㌎���H�!xG���#��m�V�%B!�(I�)�$��e�<��&�����xC1��+����dL�ġ/�45��A�$�M)0�0�ϺvW<��HN>�5=!�BY!0���aO�����*B��RI�n�w}���F����#z��p��:�|<�iY�0	\ܼ�zĉ�+"{�"H���0��Yg%����E� 0�cB�F�$�J��`�U W�0bЁ�),X2)�$T�	 ����I�%�$�Y�8NM�}ߺ�愜��N$a�1���$�d �1("�\H1Ă�%S!e"�Ӟ�5����jH-z{�	C^!
K�fr���D������r@��x����9sxo&�+��;�g�0�� ���	R���\e#�@�ՖddG5�!D�H�_g�zz���'�����2����Z���B����bJe!����
B F�HQ�X�
H���$H@��3�����XF����!��zx��d�S�0<a@�e�ϼ��!�~=����{�OyO8�{��S��ąq� �b�@�E�H��R�GWb��3{u!v#��*&Vn���	$XŁ	 5XR%���r�oy_�g��$//�!顰��O�\��!R� ��,R-Y'�d=��k�6p%�ӈ�$!��;
a���B��D!
&T���	#Fep��p;>�X�<�$���	$-5�� �i�IC��t���!S!!X.����="X�s��¥��-�0�iY!B�1�(dŰ�a�����/y���s�+� �8 ��6NF'��=����01� XB2�	3|9%���p%�d�I�	7��r�g�jD��@�#���IJnd��w]��MkW9��⤄����R	4�D�}�syd�:�*f����O\� "X�p�}�й�I�K��ƌ�D�`�;����ɛ ֘I,nH�,@�$J) xz,����������qH�0�H�R@*��8�m���}�)�����a!�&hĂƄ���E��jd�H�H�b� ��@$�B�X��M#If����Ibȉ���J�*8�z}B\�ba�s8S��H�&B�HB	"@�@"$Y �hx� ��*ʹ�Ƅ.����4c\e��M�9�)�&�:@�Õˣ�B&����b8�[�3��� �S��Ǒ�z�p�9�q�&��@bA���a6e��\|'I@�!!���43N!*B8����d$@�2���I��0��1-Zd�X45y�$+(B�X�!���
�Ir6C�3QЅ$%��XF�)o��P���cX�����t	>��ǳ�90�N�^�w0�K�KI
��d�H�!fhhu�� B0�ӆ4��ϳ��n��a���rb�H�$��P��H�"��=+�$.t�ݍϰك+�w)���<�\�#	��6a���,��<�	8x2�< d�"F�i.4�N9���gt�"IB`��3aq�0��q�ԥ��p�,\H�xX$"�f�d9���	�	!��,! @�I�/S��k�A��R�	��B�6�taH�#
�
C�����ᮇ#P�R��]�Lw<�$�D�)(|��"����$6E�Hȇ��	��$X�9$ �@��!@�Ĥ�\$� 1� 0�B1$$`Ő�a�!1LhA� D�
Ċh�,��bD�����iP�B%�P��VEb�IAcXB�}HB	�l�'�'����H6HD��I0580R1a/�H�T�pP�HG�1$>>-yK	CbFe$)!�����3H�>�B$�<���ea��
]�"Ã�φ����g�){�l�<�E) �4��}�ﲘjB�w�2�K�.L,��eХ�>y����R!i�*�B�T����C����=KS$�ƌ�� ńd9$,.�Q�7�w>�-!t�.�1O���,Є	)X1�!`B#X�"� �)�A$F�$I#E!iB�V�c����hD��"\	$� �G"Zз�H�;H|xb��D$B�R)�sHVQ�,;
�VRZI���F������%��FI1���Y�̮\)HH����vx���H5�UI	F��м���,����%R"�FYUk��!R����}ʿw�C     ��      ְo�}��     $  �     �h[F�   � �Hr��ʰ[��7eIu�UW{Ft/���p;<���n�s�
���$K)���b�"ʵmm lg� �Xvs7Vtf�㋐�p��;(�@J�U]�6:jU
P*�U��@�5*��JKte8�Z�]�,�6�v� p�m	 �a���c:��$��n�:3�넝� hZ�vʂUG6�!���M�� Zl;jͻ$�5�m  [@�L[m�6�[I-��@ `��U�@U+����.�)v�tt��U�RZ�U�R ���;T!��m��  p  �l ��`�����g���
�t�8�v�H�n�mm��-�Y��8�`	6�H5�m�l�~�Y�-���l )dqGQ�r1�����t�[c]I&�v�a�kl ��m��` �8p�Ţ�hXa��� mYoFflʫ�u UP���t���ڪW�A�VڪUr�[���N��$@AK�WJ�J�J�R�6�K��ۓJŉX H6�.ٳi0�RT
����J)UV��@*ܫJ�J�-� -�ӌ�*�05��sn�1������km�E�8jڛ�ӃTM]l�,��'�*�2u�4YOZi�PHަ�݋4�BM�J�U+��7�hi��I{`X����5���4�8�Wf�m��D�i*m[�K�l^��m^�u��D}\��Y2]�KK��ͶͶln��$ nƻ�	N��� ��L���2�f�   &�68[V.� 6奴֛l:�
�V�-T���UVۗk�m� $ d�+amm��c��
�a��&�d��u����`<��%#��4���*�O7lc*��52�.�����Шp��)�K[]G u��H���m�T�&땝n*�q�O�r&wNwkr��^� ��⪪5J�
er��
Y�ͶH8��ơ�.�W��@D�6���/o����%;v��8{>z�O�Um�:�X�j���m�Ơ @	����\�n$�� 2-�YԻ)���y���]�u�l]6�� $�g}����P`�Y����� Ĝ�J�� e�m��#]m�N�=9d��t�h�p� ᪰	  	 6Ͱ m������ �  V�)��v6��m��XY�Iڨ��k@p�jͰ�j������[B@��< H���kh"��߾�����I $  H��j
��p^�qpe������1=���D���d��[F� H6Ͱ   h� $ [)��b�Iv��Ij%���Uy.}J9X6wl�hA�����Je���� ����m���h��m���  ��6�[@-�m����lm���m�m���Z��f`q��kp$��� ۴['@m&�Vêꜯ�n���T��
�ʼ�@<�h�	V�sm� �i.�8 N(1[L�5HM������n� y�K���-����kH�WM�hp�5�����,]�V��`X�E��e��BkeV�uU6�e%��iWm����Vm�dj�уE�l�2޿��|6��3E�jKz�^Z�El�@�eUq�vU�*��,��r^U�v�m]l����(N$��K���X�Zw>4'N�De�W�>U�d�2-�6[h,2Ĝ�dS��Z�6R�eV��[l$�-���ɘ  ��M��Kd���k�m�.�,�j���h �m $[V� H$�$� m�Im�/5���l[@     �c�!��� �e�uPJ�F���^Z�  �m��G �Cm���pm�m��    ! p �u��	4U�Pp �    ���k�Ě.��u�m�m�  $9m[@�h�l$c t�@Í�   �.���6�o��� q�� h�$� � [@H�� ΐ�%l    �a���$H-68�%m�`��l   -���Y�Ͷ�����  �-�  @ [�Z��֭��[@  ���f�IGk�9m�l��d�� pm� �$�����h�E���*�Y���5K-�uU�&��U���).�k��� �uj��(/;-Ut�T 6��͉�ZBA&�mVnM׍��a��h	H�E� j�۷` .�Qm4�f�m�`9�M�m� ѭ�YV�
����
XՀm�gE �-��v� m�MoN���m[ �ݬI�����r�z�,��P�ݣC��/G/Z)/R�ݎ�^s]0U,�t�ruU@[*s�l�ʹ��pA�mRl ^�� �[@Ѷ�M!$�YյV�.���~��H����F�%�Ij�������d�q�c��n��CK$�˒Fہ ��;k����k=�,�v� ��ڦ��6�اY x�+tnӷDlԯU\<Ql���v=m�Ⱥ!d�p$4CYZ̀ miN�[n�6���� �k5��mr� �bC�/Z		*�B���\�5U�Q�(�6�d[J���@bU���.$��5�n h��d�H� ��n՛`	6�m[:�p�Zm�(pN�@�q�}��KT�S��L5�i�@U�4P۶)�7k��r�a�^s�m�ڭ�P��_.̯��5 ��wb��z����=AvʵV�7e�	����l�[	��b5)�Kp�V�V^��m�l\�r�+/;s2� R=��Su�� qÌ��K;9B��y�%�mzY�z�j��V�x�M���Ā/�}��]r�It���,��l� m�lm�%T�U�	��5J�UE�ӕ!��U�Xl6ݖ�D�$ݵ�Y{hh�U�`� m  m� 	m��'h��H�H���H���  ���6�m��}M� I�r� 9�˶�Fݱ�o��6�Hm��m��v��p$�dm���L��� ��� K��6Ͱ -� ��p�K+I�n�m ���`��� ��2Hڥ\-�E� ��m�[V�5�8��t���m�!���R�M�  ��Ag@[y�i4 ��n�I"� h���F�[[��d"�/5K�j��K��؛f�\���5&u�4�T�x͐�]����h��u�6K��9�巍8l�Lt�j�nÅª��uV�I��e��_�-�@��]7`lְ ;Z�  ۪ۻNkps�6ۍ�n'L�����%/6I��Am �l����j�a ݶ ݲ՛Z	-��	jL$�� hp�� �� փm���		6� �}o����;7Ij��� m�.�ϗ���"�s��J�e��U����g\ԓ����o m[[A�u�Sl����h�[����[����[@ 7�ͶЪ(�ZU^xUj��IE�l6�.m��M��[�mH�n�-�[�� ����Z Z��H����{J�N��}�ܒ٥����.Ą�[@9�� m�j�ݭ�e�� [Vi(a����l+m��m�r�e*���مj��Xiv底�T�uJ���ӥ,丶�m�����v�U���۪j����;�6b�s����f�T	y�{\��8U{i��V���y�:[����� ��v����m� �	�V� Ӯ1�j�{R�w"c���p kh�H ڶ�� k7[R���P` ����Un�v��(�u��oPk�n׃u�p �kkU`HH��m�e�6�%�JD�Nʪ���ppV�L�A�� R��.��ۛ`p ������M�2Z���  ,]�ʬ�Ͷ ,�^� #�	�. ��o��� 8  -��kY�uI�!%�m�i�հ �[q H�h m���[�n  rY@΃i6-��̭��P���V�j�  �e���9��h�����[mt�Y�� +m�V�4��`��m�� :K����`h �����9���@ -�v턈`kn�ۃ�s�6�,���K��OT�UU���!c������[i@�\��KE���F�[�g�� 0�j]�_|���iYq��;)�7n�m�hlp 4P$mm�m�l-6l hd6Z ְ[\'E�煆��$$�A��̷ �Ij�UC�n�'FF�  ��À�\-��N��6��  ע6ݭ�%�IC����-��{;a*�m�Ė+mu+�Ph�HXf�` ���J{i��l�f[�I�����n������b*�'�
� ��Q0�E?�0�C�z�(�D��#��%G<*#�\ �
�%T5��D���G�=D�
�:�+P�*�� D�a�S>P�T�ʿj��	���R"�E��"�", ��1u����a"�)"SH��<U)�	"!���� �D�a�Zz|�Q*z �p =(�� X�<Qx.�>>���| �`s�x��]T�D��"	�V(z|||��E:�����V��PC�t �S�<=� �(#��ʚ����	߅��� 8(|>��*b����|'�$"������T>�y����� ��-�5�b�W��_SD,O���9}Q~^>�U 1B ����D:@>S�H��Q �@b@FA�!�u��Ra����:�pOJ8�	�$�K�
�����:� $"$Tt���� |�u�O� dDx��D����5@C���@c��­����\�j������`xD�H"'� ��/tGUyĐ�8��t`"�Aj
��
x�ꯪx(`z x�z�" *�@����� �hAq(�@�(Z%�
�Q�P�`@� �H`�\�b�(�,�j��!�F�F0��s�7ws$���ݓf� ���v��m�z��赪�,p-n���D\� ���s���x���B&�2S�h����.�I/T����E�ڠ�e�h�x	�@@k�����/\p��AKn�U6���,�II�@ݮWg��5���<Q��Y
�A۳�h�^��Ғ#�Ў�yt9�,<�m;'��mh��!Uuҧv悸8�*��Z� ;(=�z�����n]�a!c���U�M�ѬOH��'�<XC��Ҋ�m)�<v���P����RN�H��K( ��Z����W�[5�Y� �uCav���0��⮖eY	-ʪ�+�b����Ŏ�A59'�ZB�u��s8y�{e���TSŭU��k ����N�P{%q�g����I��ZBR�g��#�Z���e9�Zj��rRtn{9v �M����!��t���ܓ�n60�J���hr�2e�JV��k���lO�SaN䘺�׬�/Il�:E��[V��˃1��v8��X^`H.�#�sl�ý;:Fu�i��ewg�nݛ��s0���븎�z۞�H�n��,���:���9�ܽdx�d�Ix��t��Wm�75��u��ۦ�ˮ|a��J�>4���3g�5 QB���e{v�h!��<J�u���Xv�X[;��k�e��j�ҭQ�+ny�!�u�H5T���ɋ�]�˄�ɻ+��2���n�ԺR#p+Q�X	,Hv�p�+Y�+nxn
-��4n�8�B�����jدd��F�1f�˶���(�D7Aѱq��ϓq�n�<�ijm�W&I�s�]]DN9݃N6����֤p�Ny�=���m����[��S��9�<t�u���ɐ̡�tN�tY�v'���N"W)!A�ܸ�ve���iP�14yةm
�-�]��Z�x,َZ�v�%.o-�'e6�˷J�+]�Rsu֍�j��BS=�aÖ�hJ���gi����{����qO�SuS���A�z	������<k�aEz'�'�)��O�Q`p@�`��,�}ݷs�톒�7n�d��u�v��!�p�� �n�mҖOF��K[���� v�䫃ULV�R�mv�B]���.�/e�:m�Bk[�[Z�2i}Gb[s�2��ms���A653���{]�N�lhnW��hs�s�˻<X+r�N��r�VNL��!qŜN��؝N0��Rt�Wg�u�V�ƹ's��Arg��/m��ksvf)� ��@O2�q�^y��y��� )�q�L�C������v{/d�L���G9��9����H$������$�y�}4?�R~��,K����'�,KĽ�_�-�ݷ.��ɛ��,KĿw���AU��bX>�����bX�'���q<�bX�'�w8D�Kı/O��Ι�s,ۚL���O"X�%���٩Ȗ%�b}߻�Ȗ%�b{�s�ND�,K�߻�O"X�%�}/{M�K�iw4���59ı,O��|�yı,O~�p�Ȗ%�b{�w���%�`|�̃�of�"X�%��{�J[��sL���yı,O~�p�Ȗ%�b{�w���%�bX>�����bX�'�w�q<�bX�'�Uwf�t�k��Y얧m<焺n�LڎK�����n�oI��OU����&�y�@�ow�{��ı>����O"X�%���٩Ȗ%�b{�{�Ȗ%�b{�s�ND�,K�v����5�im��37x�D�,K߷�S���H����	�'j�>D�%�}����%�bX���p�Ȗ%�b_��w��Kĳ�?��t�Ek����oq�_��w��Kı=���'"X��Dȗ���x�D�,K���Ȗ%�b{�>��d��30�˹���%�bX�������șĽ�����%�bX?g]ND�,K�߻�O"X�%�g��Km��[��K��ND�,K���x�D�,K���S�,KĿw��'�,K������bX�'� �w���&�L��0�e�4=*�[ѓ]5M	��7��<� !sۅS��T]lm��͹w&e���=�bX����S�,KĿw��'�,K������bX�%����<�bX�%�����IvM.f�swn�"X�%�~�{�O"X�%����9ı,K�{��yı,~��ND��TȖ'{�~�in��75���'�,K�����ND�,K���x�D��*֒�R U*c@
�P���"l�����bX�%����<�bX�'O��9�2C\�ɶ���,KĿw��'�,K������Kı/��w��Kı=���'"X�%��~��ۚ�4�swm��'�,K������Kı/��w��Kı=���'"X�%�~�{�O"X�{���{{`�w�[]sr�^q��<�!+آ��Qv�.砳�J�\1N �r��Ls8�nm�٩Ȗ%�b_���Ȗ%�b{�s�ND�,K���x�D�,K߷�S�,K��};|�7Hfau�sw��Kı=���'!��DȖ%��߷��Kİ~�����bX�%����<�bX�%��l�n�B�76]3sH��bX�%����<�bX��of�"X�"^���x�D�,K���9ı,O����\�rY�)�����O"X�%���٩Ȗ%�b_���Ȗ%�b{�s�ND�,���O�@}�zi�9؝����<�bX�%>�~�72K�i�I���S�,KĿw��'�,K������bX�%����<�bX��of�"X�%��z�v퍹#�\�6�/G]7N^k���7����v�&��T"�t�"����m�u˻�O"X�%����9ı,K�{��yı,s����&D�,K�߿oȖ%�b~;o�s.c�ɹv��"r%�bX������%�bX>�ݺ��bX�%����<�bX�'�w8D�DBı,N��/sfm݄�Kw7&��Ȗ%�`���jr%�bX������%��"}���'"X�%�{����yı,[�����3��׻��7����n�{���~�'�,K�����ND�,K���x�D�,K߷�S�,K������n����.��Ȗ%�b{�s�ND�,K�s��~�'�,K����jr%�bX������%�bX���w2v���I�#��<�3��v�����T
ԫf��$���p�S�ۭ�e��L���S�<�9ܼۚ��e��ݰT�Fyڥy�;B�v��6K; �BQ��UY"-ó�4d�Xz�\����Y��$�\]�aƹI����8mm�A;��hu��
�Y�ljr[����ݪ�Cf����69�p�������Wd㧪W�Űp�v�:��;��]�w�7�r�6�B=�s��+v+[�����ݪ|NS�5�9M��(�����ݓ�%�b_�~��<�bX��of�"X�%�~�{�O"X�%����9ı,O���m��v]�0�����'�,K������T��L�b^���x�D�,K���9ı,K�{��yı,K��N�.IvM2�33vjr%�bX������%�bX�����,KĿw��'�,K������Kı=������7!6��.��<�bY�H�����bX�%��߷��Kİ}�{59ı,K�{��yı,N�[�s.c�͹6��"r%�bX������%�bX>�����bX�%����<�bX�'�w8D�Kı?��θ~�Y��l^;g6�u[�W���/4we"<ގ�.�g�-���1[��K5��~����{���wMND�,K���x�D�,K߻� ~Dg�2%�b^���x�D�,x��������3��׻��7������x�C��8�`D2* �F���4#�ObX��3�ND�,K��{�O"X�%���٩ȟ�2�D�?}'g��I�C3����O"X�%��g��bX�%����<�bX��of�"X�%�~�{�O"�oq�����d
w���{��,K?
@ș�߿oȖ%�`���59ı,K�{��yı,O~�p�Ȗ%�b|w��m�۳r��s33wx�D�,K߷�S�,K��G;����{ı,O�����Kı/��w��Kı>;'g.dn�I�&R�Y|=��Ζ8rLӋ;����q������/ʓȘ(`ې�f�b>�}��m�SȖ%�b{��lND�,K���x�D�,K߷�S�,K��>�����7!6�ww��Kı=�{�'!�9"X���~�'�,K����jr%�bX������%�bX�$�;�˰��ܛmͱ9ı,K�{��yı,~��ND��qj%0��E8|6'�/;��Ȗ%�b{��lND�,K����lͻ��im�˻���%�bX>�����bX�%����<�bX�'�ov��Kı/��w��Kıo�ܷrl��wf��n�ND�,K���x�D�,K߷�br%�bX������%�bX>�����bX�'�}�2y�i͹�Phܦۋ�a�{FT���t����}�yO)��׎�Qy��ڻr�^�������{�K���9ı,K�{��yı,~��ND�,K���x�D�.��~��B��zbr0{���{�K���x�C��DȖ���S�,KĽ����<�bX�'��w*r'�ܞ�{����o����b�e���߬�%�b~����,KĿw��'�,K��}�ʜ�bX�%����<�bX�%=���nIvM3rL�ݚ��bX�%����<�bX�'�nv��Kı/��w��K�✋皇~B7�9��jr%�bX�����kn��wL����%�bX����S�,K��1����x�ı,K�����bX�%����<�bX�/ݲt�l���[�;\�rf�L�f]	cj�WV�rFolU䌝l��xa�ﷸ�bX������%�bX��w�'"X�%�~�{�O"X�%���;�9ı,O{�3��6��a��7.��Ȕ�$)!3^*���(�BS/�� ���hm�@���bRAc�R�nf�kn�s�,[u`k�j��kaŰ�m�
94��hm�@�����f�s��iH���Gi7 ����>�� >�]k� QB,Da�"Q=�e��l�6�ݶwO][on��n�P^�\���)l�]T�ޤ�[���s׳#�4̓j�8Kp.vh9�]������%Q�-��v��m:7[�����ul7���/&�50��JV�\�.��]�u�g\�C(�c��;+����۶�Ntt�DnQ%���<VjP����`+��ں��&N�$�m���3�mT�s@��,�����9�&І�\����B)���.yr�6�4��NqnË�xv���(�iJ�sK9�v�@������`��G 񼍶��/�4�٠v�ՠ�� ���YcSi���f���Z�l�;m����5��Fa�ԓ@�v� �h��hm�@���c���q��15���5�j�5�V���k�M���6�>�IȤ�@�s@;m�m�Z�l�.s,�F$dj������ZZ��jex n�nT�����/[�UԴq���n�m�������� 5�~�
?Hsw�ڜ�Vd���]n�ӒN�ݝ��E�R� � @�D�.�BD�H"D 2(!���!����w��y$��og$���h-�����II6E����������­��v%P���6ےh��h��h�hm�@:r�cL	�L�-��V ���#� ��Xg\X\�;�������E�2Ǉ���6�\�`�w�eݮ�X�l�����I$^�,t�y�w4�jR��Q�mՀ�uŁ��V&�O��䍲- �h��h�Ł�(���ç?B�;iʩ��b.�Q3SU`y��X۵gT�-�Zz�(b���2'R�SHb���"����|+o���.3{x��R p'����N<H|S�O>| b�`b�{���/#"{��g�eq@�xa�x!�Dy��aL���U���ɚ(z�X
�L�|c)	.`9��:E�ޏ��@��t�}AQ�z8�? t` � x�C���Ƣ��:
��OU¢��E�W/?NC�@/��r�7bQŎ4�#�Ww8��}��`�gN kn�=	yE{��8�r��U�SrQT���ݬ��s�rR���ΟN��X��wߑ��o�����tX�2]qGo+.�V��*Ȗ�[K�n�������ہ��zb�K��;���k\�����}A��=8�����m�񬍶���[�H��ŀv��8���Jd�t��	��Sh����wb���8tBS#���=]��;��>I��a$Ĝ���Ϣ��8 �����p%8��L*�	CT0�Q�g��ɇ�˫����WWT\��� ��^��IG����w��X�6��qtǸ47�2DC&7#���9����q�����s��-��h����wwo�p�t`�`��8����-����¯fff~@_{�@�}�J8�Ɣ�8ܻ�[x��!L��gN >��k��{��{˿?�ޕ�2��/7]�����~����u�k\��� ͹�8���'2y���%}�M��-[x�:'����wd�UU͒��誚���k��/Dw���y��N k�hs��C$xF)dX.wA��<��d�Q�5��Z�\:� ���!�[�0�L�:��ctm�6�:M�� ���m�PRh���h牃d�l9v�5+�N��@�ȑ�����:�S��[k �/��ƳIʹ$e�f��u<sc�iN����N�A͍^�^nrM5)�q���u%���8-e�\�s��$���[���T����{���{��t,���%�v� �w-�1`�m��[�Ҥ�l>v�Q���¶���Ѿ�WecS���{���s@���@������z��s�%��'����93@SNs������ �O� m�YВS's���O���<�@������8!B�*�{�ŀyח� V�R삕�f˫����P��Ӈ�)�{�ŀv�.�(�
z���ڗ�SujU]L��U�]���� �^J�yz~�������h� :��O|�t��������I �s���V�z��9g<7�{TI����Y�޸�Q�o�E&p����h[^ ����(�D(_P{��, O���5VN��\�d�6�I���9��`E"��(������_����8>�X��s���������uUW6J������uw� m�XBQ�=�˧ ����7kX)�	��Sh������������@���.v��;tDĞLfLIɚ�;�h�V���^�m����eǝ�LńȰ�0d	hs�Sة�P�㌛8���n�n���T��c���>�3y#O"����qrנ[n��;�hϳ��e^S L�%�8ԓ��M���Vd���5�V��s*9�iI�9 �h��i��U�ŀ	$B�3�I�g9��Ι�eX�^,�ve�UL�U*�&����_.� }�xvSCد��٠�_!'&F6�9�W8���9B������`�Np�����������cjs�����]/4q��\U)��K��3��K�¹�jn�w���V"T�]SWw��ޜ[x�Κs�gߐ���;�O7�0P�ja�Z��g�%航<��Ӏ�z���s�D%24�aE��V�E���]��˧ 5�xrP�L�Ӏ�� >_��'���(�E����+�zh��h����=P��:�*�pw{���gٕ�9�h���jC��Ȥ��ֹ�:"%�u���t�������?�ۿ9��L���)t���i��z
�����]�.��H���I�g����M�8Ғ)�������^;�hm��g���h�:ߜlQ�o�Qɠ?��9��U��^���m�4�GCa���rd�7�̘7�h��M�k�<�^�T{���u���5��uUQAb�F6ܓC��_- ���^;�h������F
L ��@n�BK�y������ {Z� 6 ��-�k��۬,6wf�$��Jۊ��#\	�u�7lۦ�M�nAz�e�T��^��Χ��Lo�9��r�ˡxʩ�(�F�͟;��92k�hv��cgY��]�Ƴ[X�b�J\ٶ�;F���v����5��n���W�{�l���jv��/\�y1FB8�&m�Y�I�4ܦ���[�6HvJ <@øA�d��]�6�!d&r�ۡ޺x�H��܎�g#[GW�gbڗ�2n���ލ�6����<l�7[=�-θ�ݪㆻ�m���'8 �w�=�s�_�;��`��t�<�&�ș�@-�o���g���@���Xݶ��I)��>�U7b�7sU75UWxmwN �x��J&y��`{ޚm�W�b�Rš�����!��+���X����ۼIB�����yh���q�&mϔRf�wm� �
"S������o�T]�P�G��f<M����.��������Kq(� dײ�l�������/�dZ芕Uj���? ww^ ��� m�]	Fg��{����A)�f6ܓBw��o>T}0:@�0�f0=�5��9�zn�a`f��,����ȃ7��x��H��a�Z��nh��Zyy%T{�����N ��jK�iZ�v�MU��Om������ֹ��\���4�
zGO�Q�S"��]������݋ SNp�?K�q�.�ö�Í��Z����¥�3��a�oG](\gܕ����甭�9��~���tB�_z�wb��ӟB_��^�f_F���Ɣ��7��۹�ؑ�g��[}4�ڷ�/q��8�L1����M+�>^� ��V|�i$$���"5���DF�R��ݮ���>�{ /��f��\�Ԫ��*��B�m������x�9O�=�Zm��$�(5>�m�&�z�g ��w~_���:pw]�'����kf-j�|���)��6+\����]�v�pmm"$1�n���}6��"�tKr�wb��Ӝ ��}�C�>�ݳ�ȇ�!8����^;�o�}���	Uwz�uw� ��Ŝ�L��2ΑǓ��Gȴ��^�է��������W���@�_k�ԆLR$�m:����o� ��b��ӜD(ė�����D|<�������'�}�.�2�f�EU���ŀtDGm��� ���/_j�/{q�ۄ�q�D��f�$�j�#N��Ҏ�sn�7��}�f�P�:�[AP.Yf��S�ԙ�u�<�����_�����g���ԙMcr �E����Q2s�Ӏ}ϱ`�i�rS'-��$�(5>�m�&�����áD�mr���� �]�R]YrT�,����Eo��,μ�8�k�D(�DW�;Ӏy��ErR����j��� �����J�s�_�{��8篇$�>y�m�|����}Xޱ<����d�}x�>.o��nψ!f����@5O1^���g��,q��<|�����h�2��� EX�<�"���W�`�C��1ð�� ����އ�;���Ӻt����M����*�uU��6���wD��XB��ݞ�F��<L���9�\;���˴s�D�D���7oi��t�� �KK4.��;0-uCӶ8��cJ`���p+�Ps�^Y�v�<0`;:�0ˁ�ոۜ�S�
��!Fq����v�۫�D�,�Ξ�lhwg�j����mj� sU�]��c8ځV]�<�sۨ-�b/3�6���e�&c&����q����N.�سg�������̢�ek�U[�Y^����T�V�u':cGˣ||��S�rԫꭺ��g ��uC���F�hFB��8����ԪdV�����ė[8�ѵ�K&��趻L�t��7륄k,�p��ĳ��'7%Mg�Ţ��;n ˹ל&95��"9��E��6Re�i��۾>�B��#5l��9�
2nn��U�i���D�cD@��8����,�5+r�d^�u��\b���k���V�#��I����+,����
�Ȟ�GFQ���E��Yre��Ci:�گ@�B�]t�tVzM�l�p�!]n=���^ۖ�h+7h3�=x;vЙi�֤�ʦ�.݅�:��:�HM^�]k�iv�h�N�d32��kOn�=6Ő�n�đ�;j�^c\*ia0����һ/��<��ʷ�NjB�72`�Z����PlJVv� ���Z�;`wg��vxN��u_|��݋۵���$Г7V�^��s1]���4���.Z�#9xD��ĸ��ӵ7���glL�D�ܑ=��3��s� G@��'aZ;nwMGT��K sn^$�!ͧ�v��e��h:]sW�G>� �X��\��t�ܪX���8f*C���0��! wT&������T�C`T�+-;lX�sr����B�����K�S�(������d�I���R��^�v�q��]�lp)ׁ5�t؍6�k�ٻVqvI�ۥ�2���� �za�~}Zu�|C�=����@������0_Q�>EM\ ��M�3��v�>ԝ�d�nϷ�Jz�,8�c)�N��WP���x��ѫ�8����z��a��gDݺ���;�pq��&�ѹ��JQ-����M"n%:�ukusV��)���m�O=Tl=��Zm�{1��x�g'&�0�mڭ��X콊Řl�i��_�o�ºe�Z�]n�d�yC��* �ЯnݲQ*H��wL-ِ�7&s-�
��)��nS��kL�#���p0��u7����e��KqE��m�5fzJ=�\�������tUZ� ��^ ��f���ߤ;i��:�6�2b�'i�4��o�#����=�}�@;�پĊ���G�8Ґ�	�h������Z{/o��{g���j�7�<۟6��.z_b���w���?^�� ��I5&H6�9%&-���^���z�s@�}��؂�$����4��,&_/<��ȇP�A��F�O)&�c���(j�A��cm�4��h�n����_�%��Ͻx:�yJ��]+UV�&�̒y߻Ú�H�� V�EH8�DDGf��N k�~o ��uK"&Hd��G$������h廚�۹�~\Fv�#��dƤjLX���׀=�ŀ~z�`z!/%O��Šw����jC)��nM��s@�3��]}/�,s]Xl�&��T&�a���ãrͅ�������]�*F,nYݏ`�vգ���䞸�B���[o���,�kS����^���~���7�<۟6������}�ى�׀=�� ����z(�>�L��թ�DULʈ�Q`~���L���Z>���"?�}�=��I>�;���y������ے�w%�wy'�������x�7��Xε��k�P�EW>��b�I��XI3@�;2~�Ͼ�j: ����v��r��M(�`7t�^6���)�roP��ƛe�w1��G,�<���f-���D�Dc��?�;�V����v���v<�j�ݘ��SQ��ALRE&- �;f�/o�4z�s@�_n-�$qv�R1H7�rh_b�?=x����� z��'͕t�J����n�UkТ=[��� �g���I>���$�Qb��H�D�D��"R�� �4b,h$�#@1@�@��"��bb4�=W@?4C��~��<��'�����s,�&L������~u�N�^UϽ��ŀ~���\U�L����n9�"d>#��5s�8��fR�ZIPF�s��g�\�������̢*�5J0��U��ݫ�]�����;�쉦%>��mI4�Y�P�O��,�>S����L��u�ئd��L�9����������@�}����ZYQ2c�c�䵁���)��� 7���}�`u�OE#�򂘣�d� �;f��������X��Xu�V�*夹��.J�,B�S�d�ɳwLsd�a�m�ʍU�1K��x;@��v��R��6��'F����m��k�{o���<jݷ:�g�XE6�ny�����^��1�[X�&Dvy�������8�D�;��ɞ����ڞ�,;a�7[z���1��Ň8z:���ub�ɩ�T��i�ǃ]���a.�5'[�M��E=m�����g���Kr����Q(��w�܆��o��r����Ksw��)����8�3Y�􎦐\oU�kgD7i΍�$��~�>�DԆ<R⍧'������?^���Z�*!._��� }��+T��f캵3V��^,�(�2o>X����7��o�bGz�'�l�6�6���|�`����{݋ ��b�>�l��#��ĉ�<�����o��{�nh��X
"w�/� o��n��h���U5Swx���DyDDo��/�~�,Z�v��vŁ��$qG�ҟ/�q)0�.vnQ�g�t�6;[�3�ㄬC����xY���H�,#��9�����74s]y$���W�#\�/AJ���SF�{ߺp�H
H�T�������?}'߾�y$����������2}ܷ��ۻ��n䛻�Z�6{�X��,:!(S?7ذ������&�1�n6���ٞ���k{�,���ֱ`yyB����`���U)USTER"iX�v�zի�����nՁ��f#�=�WeL�s�R�R�Ӟ�3P�Rل�G8��\��R����sq=Q���cncjL���ٹ�~[����]
?H|�b�7���UT�j�j��w]g%#��X��,��77�bE�����bS鍬nG�;���9$��ÓU��� 􂟐������:����˒2@�r	v�:O���o>X�Ӻ��R���h��k<���#2)&h����t(�����v��~�x��GʓjW-��i��w%�-��Ϊ,VF����=�2v-��v�^wm�����窻sw�C!�M���,�_s��v��Z�3ί	�ym�1��ye7�}��$|�b�7�,X��u�J!/$�U����V�]�7e]�j���ŀ|��X{>��K��=����;�ˉ�l�c��U7k�$�y������~o=*'}5S��}�ӒO�3��wf�̨���J����s`n7j��뵀=ֱ`P���% �݈US.�6n�R�z�C	���.���;�N�/.�Sw��Ӻ�H�PJ}1���������?w�s@����fg�V����� I�	��� ���gDL�ϖ,�o� ��z"<���]z�W�ڵ%�Z����?w�,��ÔB��^�}� �?I��#��c�$�3C��ً��= ������h����~����ym��fjlq��=�s�ߺ���Z�:����ǟ�R�䈉5&D�7�!lXb���t����xnF.����]p����y��tJh,�h�ۧ��K��z��3�j�k��=gl�T�7�����K�m�����-� �L9�������Bׁ-��Lu����n�1'A:�<��hGu5��9�e�E�FŹe��<�.�7��d��un���FD.m!��ݘ�'���ɸ_{���z�ߣ�9��q��p�ɞH��B�C&��]�,M�m��gC��/~������7;q�&�y�j�ǭZ�;�|��`��X��J6��6�6����77�b��o��	(���~���,�-��$�m��d�3@������i��|�-���_f���d�H���c��9B���`7ذ����%�B���V����.�*��E՘�}��~S���xq �`�`�`��w����A�A�A�A�߹�pA�666?�����a.�=��z��^�,Y	{Y�Z-��2&]�g�kq�����΅N���E�h��]��~�x�~�<8 �s���|����~��ӂ��A�A�A�A������ � � � �����n�ݻ����N>A�����g"9���0���Z�iO�����:�
�1@��h)���p�@!E!H` �b �`!Rb� 1��
y��?��`��yϧ �`�`�`������ �`�`�`����xpA� ��������wa�f��l���>A����߹�pA�666>���8 ����A �������� � � � ���g �`�`�`�z}��pҙ�.nn���>A������� �`�`�`����~�|��������>A��A�A����8 ��~�6�̳rd��3.��� � � � ��㟧 �`�`�b ��{�8 ����ӂ�A�A�A�A������ � � � �����na�':��=��]<�Nz0�l��Wi���^�d�I��{��}�O��Z	n��f�>A�����g �`�`�`�����pA�666>���8 E=�A��������� � � � ������776[��2fn� �`�`�`�����pA�666>���8 ������� � � � �������?�X"�A �`�����6M�7vL��I����A�A�A�A����8 ������� ؃�^j� �"~%F���P.�!0v�Y����(
~Wj	y*�E�$�zq�;�>�Bj�i�=�Ug�����|�@3J� ��0��		��i����$`Af��a���(#")�)��}������b�����L��A��� ��.0 k�T�(b�)R0�F�x�Aq��G4�P�: �,���_�u@�1>�{����QtW/��q�_�}������ �`�`�`��������lll}�m�~-�K�i�]ۺpA�66*!`����~�|������g �`�`�`������� � � � ��xpA�666>�6������n�7v鷂�A�A�A�A�>�����lllP��?N>A���߻�Â�A�O� 	�A� ������ � � � �{����̓�3$���L�ە1�\��꼖�G�F�{s���r7C����_��nnc0�33s��A�A��"��A��������lll~���Â�A�A�A�A���~� ?��>� �`�`��~���|�����?w)�����.����lll}�xpA�666=���ׂ�A�A�A�A�;���� � � � ���~�|�-���{��I�w32nL���e�8 �Q$BR��t�K}XzG���z�`�����mrL�iH�ĞE��\u�`���?n�X~�$�DDQZ����I#lħ���z��9/����->����<��Ut�]=��=���rj��8S�%f����n��i1��S�c{��<$��Ȳ7�{ذ:���w]w�޾0��yZ�2!�dȤ��U��z��נ^YM�{w7��T�<�'�H�E�}-�`ݳ����X��Ӏ~u��ԆH8��M���)�~�n���U�~]�zs��Q�Ŏ19$�K0ۯ����/O�l�z�nف8�Dd�;��l����K$�t���=C���ԯ� �[����n���춵�uu;q��}���-7#= ����:Y�\�l��[k2q�{m�\��7)dha�ɝ�TQ��s��k� �7j�k;����ۮ�ǱQ�㿞}��\�$�a�唸	W���0H*��qFKur$��^�N�"s>��q�����4]��N)�F'PO:�S��������z{��=�ݹuۛI�m��GlRƝ)ֺ㭒4���}:Է��v���[��^�>��l�����&�u�{���{^�ye4�����Z�rL�iH�I�@�;��������}� s�]gD��^?H�f%>��7#�=�O���i��%	z!Uzyw� ���`|��	�.�&h��h�;��X5k� ��.q{���̘�Ȇ�E$��湰<��F7���W���Ձ�5Q����q�s�md15�q=�0q<Ɲ�k�'�n��ڮgHh�Zfz��l�3����V�L�;��{�\�`=?M��uxmHc��pM�&�ye6c�a��ABN: ��T<����ÒO�����ݶh���y1c�NG�Hh�^,έu�$�IL�ou��|`�\�Fۉ�6��rf�sٙ�}���yPo�V��@��Ĺ���ޏO�\�bCI��$z�����h�n�Ws������4�@A����۷�f@�y3�F�X��6+�t�_�{����$�
3�Lci�?��x�9��X�Z뒈I~�>}׀s}8�jW�L#���[��u\�z�[4��o�Ͼ�H���LJa1�8�$��;���O}�w��#�J�H�ENA!*��OTA������pv�s@���&���q�D���s�� ׶��ŁД������xdf8�<�RM����������v�;�9$����$�
�X`� #B D`�d��;m�<Z�s�v6���2�2��l,cygq���u��䞸�p����~�׋ 5�w�~��\�H>w� �.�n&�۟1ɚ۝�|�οyh������X�g������S57a4�� ��k��>y���g_{ >��s�c�&ىO�1�ȴ=�+�,��V�k�$���اq`=�!*	�H����k�`y(~O��9�|���h��\�&)�<���x�'�^ٝ���|]������=h
�N�M��x�R��Ja>p��E&~ ���~��Zoe4����?^��&���sH$�� ��79䒏%G{�� �{ kZ�<���7��|Qt+��j�����=������j�5�u`w%��;��7�f乻�eݜ��A�"?����� y����������~�t�yz�6�McmO��� ��٠}�}�g;����x�35ڰ���R��s��h.�\ 3�	��Y�l����c.k�q�����Q_��.�q/)m��R��U�e�w=[��{\+@��a�q0^�i-��Ε�^�vt$�s<qm�]��94ͱJ��6ŰP�S#���;=�ZN���n[��Ѻ�up�;��Y�r������ {3H�ޤ�͘n�#�&�����X06�P�:w]�alu�p���:2�Dkk6�P�Ѳ"�%�T)�ٷr�����y�r��	��swe�Sfj�Tqɼ3]74E��Y�]��\�
���"m�I䒁�g����9۹���4��V	C�Lcp�;{)��Ȫ�b���^��lΉ��/�J�)R���&��7_�X����X��h�J�Ħ�"��)3Cؗj}x�݋ V���DB�%M��,�(�!���)9�c�@�-��/lX��XŮ�XKs
)R�Q1SǬ����C�nku-�NW{x��)wmv��=m����M�-�#�ȄG3��Z9� ?����I}A��ŀl��*���Lܗ77K���O}��9B'���q�[��M�����[��"�x=��3j|�&h���@�,���}�|����ۚں�n91!�܂O.��	N�gm>��Ł��	7�s��@���/��}1�I�@�}�`}Ż�utڟ���t��\�����8�5����Zfj��f!F�щ�Y:��r�&�fS�F�Ns.c8a�\�	������ x�Ձ�ݫ���i\���|��I�y��}����݋ �Ӏ}�x��"d���J�]V�U��Wx�v,��W� ��P��$s�N�}j�:����q��V����fK�X��$�_�x��b�g;f��ع�{�hG����0q��""��35ڰ>\�Z�]7޵`w3@���%��=7H��<r��G9��<[�Z�jY$=[�s�j�gr8�K���|��]؝wLW$���?}Vq�Vq�?.vu�s@/����Hi<nby$��YL䗡U��`��`���<�(��Iz5ßLcp�;�O9۹���"�i�� ���}�w%TR��(SE��J7_��V��`w2�y�P
�F,THA�0qI�Ei�D�C�(�}E�l��Ɓ��+���H�8ܙ�Y����.k��������j����o��k�b{u�8��Ŝ�=BK��ɹ;q�l]�ñ���u�T	�׆#5X�L�;��`fk�������/y/�ɑ��IC@��)������P�{ 4�׀~��3��>�]\���`��AHh���s9l���ϳ�}<h留�г"x�1<j|ɪV.qDj�z��W�1�,>�9�߳@/���(�O#��=�-�`u�e���Ձ��\��M�K�����# �Ed;�,�-����y��� ��� ���V1aL0�E8a+�	 �"��`8�#!��Zt�`���>��HH��ac������A���$��u�Ё$>�|DXO#��M:s�o�����Q�	Db�&9{�Ç��)!"� ��c��bB���:��+�B*@ �@H�>%%��$&��%-���$��g�Q8�VP�t��XBE��'�q��Q{M��m��b�b�b����6{l�����۹�h{EG�^aէ��	�ӳöÞ�m��PHt*q$h��j��ݥf�(
@�ϝe���W,�n�C�7	jG�*���t�n���0E'�����O&@��ۭ����d����X���\j����n��YĹ�/7Z#l�	�j{u5clDR�!YB	�C�=�iݎ�6�!��5bՒ|�u*�.R	�m�ӹ��<���T�!d�$ UO�
�u�I��� (
RZ�MR�&B�&��4�я`�.�P��H
�WW;.9���mE]ںM�������h!�t3l���3���g�A4�LjVH�+nX�'����Mg8ik]V�9�+T-�<&��ۆE��.q��8���T�T�
4s6*��C��Vj��Z�%@8MU\���+N���E�2�YE�z���򬲇�դN��%z�U!5ՉG���ls��|X��S�����5li�c!;<�˻$3�ۙv4�n�j�Q�dvd�W�R�<ð���Gw'lK.�ے	݉<v��h�dԼq,���R�R�KvR�q�j�{f�3���l����f,����v�k��g�E��A���ѱ�v��f[��f5�m/+���#F�dF������շe]�8�ع���;f�kPt����A]�Jkg�#u;*�Od�N:�L�]�d)c�ͳY��vx����n���V嗕W�`�RUGc���% V�ظӵ@M���.�R���,��Ղg=��P�(��u�����.���=n��*N.1#[[�ub��l�u�*0󧔜�1��ڕ�As�PU�UK6�i�V�ַ:Ҳ�3v�w&X&q��EUm'e�S��*ܔ�3:ka7'MPpH���N'��@ М���V���vq��L �e	.C!�6�t�m�v��;���5N��gR�M%@���4yZ�M��\b5�R�<5Gދ҈t�`��(u?/���b���Q���(I~��ncQ�m]�����a�'{#�i3�ŕ�W��4��������S]���pa��5f��X�nҗ>��ǫ/v$�s	<�,�lh^[�.�c[�=��;<�[Y5���g���G	$�9$�b��	Sj�+4��[0â��M[&tF����P�
l����΍���Z8W^�ܹ��Y�]�Y-���;On��q����<s����٤�?�Hf(�Fc�B��2dm�F���jɁ���ѳ���8������֖ƣ�s�bRg@�}<h�n�gV���/�5�ذO�EIT#ʕA1B&��35ڰ25k��ݫ���^J*�.O/)�W"���UuWk q����7j��e���Ձ��bMcy>N(Ŏ=gع�{�h��4s�sCً����8��22q������t���������h�U�2<��	lC��I�3/�z"�ڋ=������V�ڥ���?s/N��j��*����j������}Ĺ�.��}<h��2	�"��&hpn�S\]�:�*���5�Ձ��Ձ�v�h��Q�6��NM �7V6�X��Xh�X��!Ԩ��c���r۹�s���Ζ��-��?Z(مǑds4f�V�5��t�zՁ��V��8�/isp^8�<��@�-Q\'�vls˸����o
��M��.�4�2�}�߿�w�~��X��/B����`�3�ZLo'��S$�?r�����Go���w�ۚ��4�Ԩ���8�#�`f�j���j�8��s�\k8�ɮ�w�s@?e�����)$���fk�`�Ձ�nՇ�k�����S �9��9�rf�s���-��9�w4s�s@�*.n<#f5P�2=��m�a%ŝճf�kݦ{Fw�xv�wc��m$���0mc� ��h�[4v��������������לn?�>��crX�ڰ35ڰ���;������x�K��CY������v٧���~����X�T�MLڸ�������`y)�}׀ou�6�`	TF�C� ����U�����?=OJ�G���?{ȺLM�y>s$�I4�-�=�X��X�u`u�Dr93*fܛk�p��.�z�61�D��3����'Nܫ'm��C�)�-8'J9����`fk�`�Ձ�nՁ��52�BjH���4X��_ˉ%�?��3�
!L���`���7�d�jK�Z	S4���`�Ձ�nՁ�i�f�Zʫe������&��;�~���Ɓ�v�hyl�9�\�?�9\�����Ǵ��K�����W@���'��{9$��>�� F!�wwݿ��P7^�*��t�: �N�S��e�b�/n˶�]k�u	�����V��[(ń�V�b�'9¦sI.P��Nĥ�ݏ]���ݺ�m(���{l�tQm(��9����j���MwX�і��j���k���76�B�i��;�x|�y��;<�nB8���qy-��6�6c�1ڶL#�%�{A5����n	�rY�i*CfL̛��4�\g�g����s>N����w�f�1y��Mۃ�X����Z�Y�C����l��m���� �n���|��H?�_s/�S'ɸ�8ܙ��@?r٠r�S@�;w7�3�=��M��̒	�,_�U��i�w���t�q��;����D�14w+K�]� �nh�[4��Ǒ��b�ɂp�35ڰ=}��o�V=v����g�vɺ{���z&�e�yi ӟ����|/3ܓ��MmR�]x����9��m������u`c�e���Հ3\��SJff7asww�I���	膋�G6K�f��x�~n���_ʡ�yW���9���ۓ@�ޟƁ�v�hyl�����tJ�'�Ԫ�aPMQa���8���{����`�Ձ�i�d�n\Jd�7��4��h˽���;���>��X����U.����5PLM�s�-��Mq9k���'���ã^=N�s�	1m׶ЈM��̒	�? w���9{)�s��hyl�?WEFFd���m�$�>{l�I(��7{�`����n�IyU���]R�AV����j��{I'����焂	�1��"��$^��#���wG��7=L�=��T�A*��v�<�gw��w���v�D(���� 8;�n�Z*��Wb�����������w޵`�������&���qL�<��6swI�!/&η*ț%nv���2OER�7�*-U��t�1�V���1��1����ɉ��4��o~�>ă��h9l�?r�h\Gr�L���iJ��� ��V��X�L�����K��fO��1�&�s���,��{�{���!�U���9ϻ�h���̙���4ܲ��7}���V��XX���0TI�W/<'ct�e���vx�^��qu���ō��B�f&8�<���a�' �-��[4��h��*��)�	��9�NM �-��[4r�h9l�g�������r��h{�M����[4��h�T�7����nMb�}�4����s�͓� I s>����ޙJ\��J��b��0�w{���v�I���I: Q`$Eu?�ȝ�����[�޵4q�V��n#nwvx�'E-����l�Q*��X�c[=F�Y��9���nf8�v��kXT����������z�Rۈح3:�ʯBD�nծ"�lI��:{:���5g��^�^�أ�q!dN܆[�M��fDaZ$��U�^:[���+z�ڌ��!�ݩ�i�:�-���cS����J���2ӧ��E�U�|.{�X�c�qO/�gv��`�ckl�]��nsawG�1]�=��H]��M'=-v�����t� �n��⡠i�'�'�4��o�>H�}<h{�M �;f���Q1��28I0nI�w2�3� ��V��X�r��o&0s܉8h9l�s�h9l�?r�h^Ԕ�G��Y��&�fk� �n��v�1��1�"����i}�G"Λ�Һ�a��!ɻ,:�G,E�/l�[n�.og�ɱEsvU���� n��`w�`dcs`���͖����fk�L�����{�D��b�s�9ũ$�$��U�.6���u`�f���TI���ɉ������ ��V��X��X����UnF��nM �;f�s���,����]�4{�/cHM�>�8I�� �(_og�7{� >�]���WKR]�y�ϳ1��	p�=:�8�S�a�UŸ܎����Z�$�����]4i�d6���� �n�3]}����X��<���a�'�����H;����脢?H}�|`;�L�M�-��D��Xf������;┗���I@�1jId�+cxPD=a9�C`F6uO�XRYH��̟�������Ŭi�V �\3�H�PN ��3�M1�`&��{ŏ���	�O� �:6�u")�"@!n&:}�	��x% bʥ���asTC�aN	��������18}�~�/���w�[�����LR.��9�]�u��;�Հ46�iM"feT*����F�V�^,1��:�h봎9ßLcm�4�(�;�����N }�w�6��(A5��� ^=�mso�PJ�х�-�Z�W�7�p�%�69��bfLL�G3@9�f��:��3�.�=~�`n�C^�)T
9Ǒ�4��� �-�{�M �-��9��4�����ۋ@;�zh�e4.Z��ڴܲ���ɑ�H���m����@�]�d�z�
�p0S"1�Ĭ(�p=W��;���I�����4�2a�N-z��Z�[4���;��6�����'�O�O$�ٜ9�l��j$=[�r�K�����F�v���x��bM"bj��~�,1��7v�`�� ��T�����Ȝ�@9�f���S@9�f���V����bE�����'��nM�<h9l��.+|�w���/��]Q*hG*V����0;��U��ߦ�3�.r1��`n�W=�L���kF��?.�������Հf7VIg�.RHIpP���oϫZ��n��v	;q&�$�M�7$D��-�05+�E=
�8[K��{]s$f�k����ā��(8�&�^-�n�'l��״�޶���mkk�O�eC��j�\��d{t�a�]���C��}u�t�`��#K;��+�t�Ύ��N5��ɮ*W4�;,c��lp��^���]��>��.2���������X�\�2i�,ި'Ç3Ip˻	-I���;����nF�����y=�ڻ�;Qm§�f�Z�Cmd�D�JG@�w�@���� �-���נr�7��� ��M�������[4˽�@��=��J��}^T��Z��E�]�v����n���Ģ!s�n׽�� ��20�c��94=�}�c���M����X�L�21��k�5*i3(��T�T���X/��'�w� ��=��k�;]u���Q���$���#c�30	l�vsu�l󼀄��q���)}1�6��?w���[4˵ע!D~��w���u]4��]+SD]n�I'����hb� ���"D�z+���6���rI����rI�{)�w�.�JdF7#X�7&��v׀|�ه(�3�� ����f媙k'�'N=�ϳ��]�v��@7��СO��� ��WIB�*ɫ)T�n�,q��;����`~����o~��Cjܻ���f�{T��;F�n�7gvK�J���MpJ���yuĴD�`�Ձ����Ǵ�.�ku��=��x�h�c��94˶����;�M����A���ȁ��uʩ���7μX�L�x�/��B3>}�H�-zz�Z{`�"��O�1�8h{1v��U�y�W�����-�����7�����^��:����|`�\�N��
�� ^����ە�s\h3��u��l����m���������/�\i�t,���z�����;_j�:�k�?s�+�!��|�q�#�9{)��"��-���@꽯@���3$��r��8�7xr��]Ӏo;� r�4�7��Ɋ70R- �-�mz/���<X�}�k�`*Ī	��b�
�P(��>����7V�{�����)��rh��-�\��`�Ձ�9�����ڎ��n���qe�u���Q��Xu�L����klm�2T���l��݁���|`m78�7~Q�Ce�V �ApQ�I�М4uڴ�Z��nl{L��q}�*�ޘ��b'��&J���l�lPܭ,���`n4�D�Ɉ�F�q�]�����9�j��ث��v���!��}�n=���:�ZW-z��4�6B�OvM�M�&ۅ͛M�ƫi�ӳ6+�8�l��ي��-�-�n�p�]v���c��V�`��8��t�s�B��NWZ��\u��g\ōH�Aaл�f\��-�\n���]�ج��ʌ�#T�3c8�s��3�)���%Σ464c,�{X���E�A��m���������NGX�9�6��*@��T��Q.��[E�QKx��[G����G����a5�6�8�t��Tؖla�ɜ�:��m����]u�t�����;羁�Y�͑�p�|��Z���h���?+]Ǌ<�&LQ���h\��ol�9{)�v�տ�$��c�G&71�����r�SOf%|r��@9kb�����b�C�}��S��� �Wzp��x�]�]�;����'͂p�;_j�ݶhol�9��h���f}s�����m@�B'���.�t���L�9zA�ݸ;=a�c\�b�W'F�jHbnyq~ ����v���즁��V��4��
d�Ilsy$�w��8+T�A�"0K�\�.BU4m�2�{:��;�Ձ��Ɛ�Y>q85$�9��h��i��#�ޚ}}4�W�$�D�N&]]����� ��^ k�x�P��\���Z�<Q��2b���@?v��z����e��uŁ�%�:?Q�tQ=��=���9�Y�㚔1*�ϯ�ݾR{�wr)�V�+���1k��~�����ـk�s���׀�U+����ϢRI�v�SĎ_O}}4���4���I���8i'�w{9$�w��'ƨ'��Q����X�S��%�o$����4r�u$����CC�g�}�������v�S@��)�[ؕȅ2|����94�����?���@;{f��Q,�z��ܘ/��1��q���.X|�i�ح�[����vܲܤ��.A[y>�85$�;{)�~�������}4*y�L�#dr-�m�<���|��[��6~n��O���<����b��' ﯦ�s��O���_O��ܸ��8�1��4�Xn��61��;��a|J���s�`x,D��FdRAl"�3�S�ӷV�٘�4���5ʈ���61��;��`�Հf�����|o�s�ui�g[���"P�[h�غ��\�"T������+7-�u�����L�z��3u׻ �}�<ף�JH!���$Z�fg˾���/w^��u�k��<�&Nn�y\�j�nF�Ȝ�}�M����ڴ��h�خ6�I��D�Q�4?�U��z�� ���I*���x��R�H̐pc��#�;]�@⽯@;m��}}�s�N�8D�*���^��#�J�#���+�a�<�#!<�C��N�2`ʷ`"D#%���������b��S� ;�� �%}�:�2���D����}���z���
��� ʾ�jd ЃF��<����O���4��WN�`��8���XMR�JY}>wg ex��4]W� <@ yG�� =M F����$!�Y�ńJ���.�y&���q_K�==-������nE�c��eo@UvͶ���c��t���;Z��n�J�a��1�ΛeA֤�:Һ���m�V²�$8��ȓ<�f�b�UVn����dж�=��r��g�NFT�"��Ԅ�s����
��9Vy�\�A���! �6��p�khG6c��N��8U��ۙڶs�e:��!Q��Ú��m�B�d :G']lp�g�vV�!K����Ү�c���9nx�=Z�n�Ӟ n�F�-�8�8R@� �SW��W�����6�h�WNh;n�jUXv gI��zE�U^���ݹ�-�]qm/S2��U@*1U���P�X�xW�L�yؒMā�[��]��->GR WMw#���={<ׁ-9k]�ˎ����L���,Bn5[N3(ڶ���]6l�2����%F$�%@�� 4�n�eh�qn�t6�	ڠ�YZ��!h���[�]�n,0��'X�	���E��Jl�}=�Z�i�51f�h$pa��*�FGv�T�H �Z�vB�Ֆ����ǲu�6\\��ނ=I��m�t��\�َ��9������a�^ul]%�t78����n��8v�gq��[�g������@��;��s^-��YX��Ѷ��Y�MÜ��,�5\Q� $���hyKڶ�
�< <���5Ʉ�"|ו@��ؙ,���&���n��[�x�ݰb����N[�Z�̚t�V��qb�l�sgf[Jvl�kl�[X���kNn���]�n�&�;�lm�Tź��8x�w]Wv��Jqv�	,���z��[�H�9����óa�6X#X��9Lk�Nwd�����]�S4!���g�]��	˪�;F���\-B���-F�`vj��)N��j�T��V�'m�2���k�v]���<u!n��8��
�6�d+`Z�v[��]Z� f
]ۘ2s����f��R �#�N��l�
�6��o�*�^"�A8����T=QC�����t+!SӝQ0��S�S:|��w=v.(�u��؀�
u	ȑ=bU=�W��2[�-=���b�6N�]�9�ǜ� M�P��S�b0�fe[��l�=�0��ˣӋvK�q�\$����*g�l�j����v���v��pv�]f��U��3���x�s/.w5z�A93�����͒.#;\�u�͹��7L��O�=�
'����:�Kf�� q�W���=B�} b�ۄ�sh��'stba{qˢ�ck��nY�g�cyΚ�y>l���$�_������٠uq��BK��{Ӏ˗�]"��U��I
I�������ڴ�پ�{ͥ�`�x��)$�/����j��f�s���los����qI�λV�v�4��h?���g��}�_e��) ��G��hkw�yBS��� ��� �i��9sx��ή���\���xۀ`�{v��o㊩L�y��%n�nN ]��{|tb��T�b�� }�^������/����9l^��i<�H���M�ڷ�������qw�v]ŀn�V��_܈2�S�3$18cn-���@;m�;n���Z�����O�&(܂r- ���:�`w]`t�_t��5���8��jbB�h]��ٙ�a������wN ?����o�<"�X��������ŹP���ܺ��W�����91u�S^q@�#�Q�^LX6�9����?�������M ���}�nh�4�9��Rd������M �h��hW���G�������r}}4mڲS\��8�r9�,�Y6n�`^�%rbS'���xӓC�3���]��� �V��	yUw�׀k�ϕSm'��q
E�u^נ[e4��h�V��W�6%1!L!�A�;i3��6�0��C^:{[����49�v�ߟ����(�n?�{ޞ4�٠[e?� ���@-�ő��6L���r�]�DD��݋ sϫ ��f ~�p�#�X�51(��{n��mz-���f�~�*ү&,#O�5T���ln�`�Նs�o��@x����}�y��'�����vn�wM�����e4��h{l�:�kݷ����˳�=��!x���Ty�ڱ�ˉ��n�	���<gp\뢱-�[i��Q`�Հn�V��67L����JdF9"orh{l��*�����ƀv�7�#��^ƛm<�H'(���9�Հ|ݳL��^ �v,��ז$̐py#�9l��v����sC�*�|���i��Bdn� 5����� �V�wM�f�|g����9�y�ch {ls�՗����k���h��P���>�n�ey����.�z�&@u�#i� j���.|���'X�Ghc�D�4�HYKILؖ��{6&�k,�4٪��vq̒�����YYJۣ&��1R �q�FWS��#�2Dm��`�ɶ^�GNQa]�'�:�	_e7\�,m�6�uX�q��2]F8WPV������z�������}���tE�·Ji�:qK$���,溑3�F�f�����ں�MV��޵`l=s`c���5� �r�V�i�&������ڴ��h����ى퍿G�������?yhol�;�w4�����6����rE���@�m��:�k�9]�@��;���H�I�&��۹�u^נr�V�v��I?*�~�^����m��c�d�nݶL�Tb��:^�g�$��o3ࡆ&��Pz�A8�&~���@�v� �m�ϳ?�0����4����2A�Ġ��@�����qi�@"��H��PbY�.%�����;�j��t�6[� �{qƞO�&F�d�- �m�{m�tκ�z�� ���]\��JbQ94��hW���ՠ��@?g+iW�m<s�ӆ��{^���Z��4��h��ck�L@�Ms�g7d��jЅ�j�&77]��;�On�v0�J6�s$���4�n=�ڴ��h��:�k�;�(�s���rE���@�����������Gr�S"1���-��U�����] �/�(z�p*?�U�A"��C߾�y�rI;�{��{�u\cO��q5&h*�|�
�����h��h���L�py$����u`cnՁ��́Ս^�����N��޶�sp�xmts���4����m�`�X�q�t�ҝ�s�G� �$׮���`l=s`8z��75CSU�qc��Ģrh�S{�l=|�^�z�u�� �w���bI��ϓ�e��y�l��z��m�Vsb���$���������y����9���$�@>
$�/�*����I;�(�s7�7�v������������®�	�䆲'��҇��3ư��TQ�c���˸���A�àM6�dQ"f�R
<�D�''�;�{s@꽯@������h��16���7&hW��]��ol�9m���H8t�=fL�"�$zW�z׮�mڰ63\�q�52��%r��I$z���������Cث���\/����1��D��9m��63\���^���qp�\9� 1U=��\��4ͻ�K-�p�z�i�9D������kt�=`;���y�3����7H`�o;]NZ�w�"8�&���[k���\�٭�]/���:!��`�1K��H8��]�s��Aӯ$\g<4;-�0�n�M�V+:�9����n�+�ˎ�(.�Itl=R���-���O=��a=d��[m����)2%��tm�z�B7n�C��ڡ����w{���������{��5�=���E�t����j�Y���
5��Iq�[\�����e��OT����}s8��ZWmz��?ϳ3? �����7�&I1I>m��ZƷ6��X۵`nθ�%ĔA��71p��q�w�z-��{>��
�����W2(�)cq���h�ՠuvנuvנs���&�y>�R&���ڴW{��_u`6�`�w04Q MIg<v�Ǉ:�a�Eu�l���cH�F�%��۝'+�tKQ��3&G�A����^���^��n���Z������}�$�����{��ńj���@�ۻ���ZWm{䃽��	0�,s��z}�nh�ՠuvנuvנ�������ϣ�f���ZWmzWmz-�����L�b�|�QH�������[w4Wj�9���#�@�B<a$`�N����]�4�L�\Bn���\�L������e��7���^��n���ZWmzWY[�@&9"Ln=����ڴ������q�q$�o'�
Dܙ�r�V���^�'�tϳ>ޟI0@0#H� ��@�[c�"��jÔ��D%$�" ¡��i�ʐc-m�`���j���@����Wz��>z�,.\ȯ�/u�"B��'�0%F�!`K*�EAGy�=L=4M{�e(�Ɩ���B�.U���)���O�$$& �:'��@�~ q�|'��芁�M�Q ��E���PP��4Ow��y��y߻ß��/�Lɑ�dPiŠU}��@�s@�]�@?r�q��6O��$�G��@�s@�]�@��M��߿��MQ�tQ=��=�x�i�<�5��Pҧ���O�JOrN�u���mst<N�t�(�����}j�͖������s��zhp;O8)��x���3@�]�}�EW�z��M����z�j��x����R- �m��l�9m��;�j�g��bD�n��̉�c�"r~�3?(IBJ����&fg{����fe�y&L�؜ ��`�?{��g�[o���N\%��,I�5$�-���䒶]F������J�&���z,Y�U��7�\�9���q�:٠�̀^-���!:ϝ	���2GFƆ�%��d��H��?~BV���$��m��$���jI.[g��$p�O6%�E�I�RI.�����ϳ�m�_y�I%�{߳���wqo�i.w������)29$��$���椒��~��۾s�ԒJ�z~��B�gnD�FA�jbQ�椒��~��]�QjI%��?~I!v�5$��μ�7�x��s?~I.�(�$���o�9Ē��Ԓ\���ߒI��x��F)B�!�zZ����u^v���cu��9�M� �۬��!l q� ��Bp��n����}����撕%��^vLc"�^�^v�:!E�nǮ���4��d�n2i��i�g��AV㴳�f0���Z:u$� ��;-���n��M���]�r�:T� Z�5�8h�(�#�#,�vb�j�u�TzH�8/'@q���9�Y�Wlx��W{�}�{�|=����1��M���Q�IW�<��O]LF�$.�q���0$�M<U�k����o��I���$�m���$�k�Z�K��ѧ2$7�7'��$+k��K�����IZ���]����]o5<c�%�8椒��~��V�E�$�{l��$�msRI.qUq,Hy>pR&��ߒ_�f}�?zo��$�����$�msRIr��?~I#�kǱ�d��,Q�jI%��?~I![\Ԓ\���ߒJ�(�$�������س�)��'8u�Lba{5�ogd����\Ę����ۗ^��N�[l��sym����ym��oe��~m$�����$+Q�⌃��Ģq��DF6���թ.�j����9j.""#ol��$�msRI.���1�Lq���$�wqjI%��?~I![\Ԓ\������j�넑b�cq9�R^�w����$��y�I%���?~I+]�Z�K�;4�D��8Hܟ�$���jI.^����I+e�RI.����q����sԻӴpp>;OT�؜���pk�!ca�G�D�]��v��Cض���f�$�}}�?~I%l�ԒK��~��I[dԒK���X'��"rL��$��-��}��I^����=��jI.^���������fġ�#��`��RI+�z~��G{���~:"�'�� � o��tB��s<��ym�����[m�{�v�˓���RG$��䗚���Ԓ]����� �Y��@��QrG�8��jbB�X�ڰmՀn7V�XM������=�z���[���,�M�t��l�Y團��M�Ra1=5\9�7�J��ﾫ �n�mڰ1�`f�!�Ib��jI����ċ}��޾��9]�}�G;}�9�!�N]]��b�׋��ޮ���נ~���j`�IƤ�}�޾���}��Ղ�1pU�$���}����]��<�8)19&�z�Zol�/m��{f��V�F%>H�.�g�&7j�g��`�<9�K�8��n��������afF��fL���$��{f�{n�[�4Wj�*�]Dk'͓裌�M��s@-�+�h��@��q\�b����Ēs4�٠r�V�[�4��� �:�;"��<s���9]�@-�{e4=�{��@���HE�<B�r- ��h�M�q��ذ�78�_(ԢT��!B
�[ Q�dx�w��u�u�s�×i�o'N�d��ظsŭ���ـ�[k7o��z>\q����Zغ��ZC��ܨU�&�J�P�!=��f���X�ΩN%L�%�j�!�[7v,a��^��"u�v�牋�j�sa8�q8ivnm�&����E�6�4��'Wa�$wmXM��mpdq���Ȝv�X�%ɸˋg���wb�ӱ�I�y������-�=9��d��.=���J���)t.����ք��]�|lh��n%1�7 x�!�����=��}�~z���_��׀}�ꥩ��I$K�[۹�ċ��- �����e6��}����	���H��4�j�{f��e4{w4��6$̙!0!�@-�m��-���;]�@��uo'͓"�2I4�)�[۹�v�V�[�4�6��o���KvN��z�t�)]�C�;58��lk<��:��ݬc3��V������=����ڴ�٠v�M �:�;"��<s�I�k�o����.�q.�&�����z�X�jb,rbo��@-�z�Z���+�h�۩FLn �8B94�np����w��3����}T�0P"�4���on�r�4�w�n�s�rP���&�v &����#M�My���ю��x����[����5�=��%�y>pR'$����4�٠w������2s�*lI�2B`L#��7vh�݋w]� ��X3e�F�cdȣ��M�v������_� D`�@U"�|�I.Gz�Z��<u`�Ձ��CUT��1��(��-���[f�[�4=�b�{�@=�}19"��7>�ԙ�6� ��������x����z���2ۓ<�ى�&-٬�\����%n�'�On^\ �;O	f������Ձ�-ŀ޻V���;�����'G&�޻V�on�r�4�پ��H�K��S�@�����Z��nh-�@/{f�޻V����	`�O����4�٠��I>�;��?Q<'����r���9$�r��bL���94�٠w�ՠ[۹�������0x㑡O<�g7����U�mG�^n��u�Xuέo
���6L�H���;�j�-���[g��������Wh��LQ�s���\��ŝ2�׀ϯ ݦ� -]��,Lcs�I��l�{f�޻V�on��v��ԑ,#�)U`�����v������5D8� ܚ��S@��NI'�}��w�wy$�\!WH�<�Q0D(8�c	$�CP3�WSĂ�xG����#<���X��<����
<A������>O�OA5B
>�|�`H�F(��yN
z��I멤`��YqO!� <C�>	��b���<|��{6�q><��O1@xxpH�T�|��Ys����(�p�$R@&l���Q>C�D<>����@�iw���dBW��b$D �, �0�E=W���G�6�lqÀ�k�]G�όhxx�<�X�����!��z���u���2%[��i�1[ 0)��WR�!�*ڒ쭰(��<6��ڰ�U�tl7c"�7�"�؀�:�h��͈��sհ��v(st�@lr��n���%�k9l[:�`�9y�)��ל����N	�g=�G_��~��B�co]i"�$�^T��'
�� �n�-ä���q���n.�6�u�Dr=��S��MF�×������(���kl��
�QVQ��Z��@�J{n�*�P	(��8�x�2�]�J�6��:*2S�\2l:�j�AJ��:��9Ѻ�s�"ml���&":V`��u����khi5�kTv�N9s��l�n�j��;۶!�����Ö]����U����s�Լt��MUR�\�!@T���H�U�ee	�yvg�W(��N�U;�O��Vv�&�Q���N$�4Q"��Iyf�`L�N��<j����U!�j��K�N4��6FQ��jP4t��Y�X�%�\h0�i��5��d	�s�D�� �x�<de�/5�>��@��i�^�5q�uYt�&�ո,���nk����cN�Y�!˃���J����7\j����t�u���B�Y�˺ܜ0v���P�!��=�^e.�H㰭��&�ۡ�rrhݸÌ�ң�V�.3�N�����T���3t:I�ސ�L�wc�q��8�d�j!&[���	��f��v�
(ͷM�
D�
v��]�f��װ4�ph�{Al��ۣ��4��I͞�b�s�&T�Ij���z�]5����v��S��M�׭l�[<���{T��m۴��R.�V�E;3�5GOs���9e�����������Jt:�]�L��t��Z��R�iUٰu\L�m�X��Y��)���>���.Yle:�6L����Ӫe٤�W�Ĺ%�-�,���Zٶf\�[	&�Y0�,/1J�P>T<<����A����O�>>�E 4/��@P�~:�3d���4���ݮ6�m�����e��i��=2A�R�B�Y�l�Ns�yI��L��z6�b��0 �:��Ȏ�U5��m���۱to[�#Mgul�lձƻ'M�.ɦ�C�\�j�L2-'j�m�B����n4�Hl	��j�@h\���õ��cJÑ�ppv�a�0��We���Y����|齧X���u�n%�� �F����o����G�dg���V&�>;��u;%�+��9���89;t�zD
S8��ض��b(��@o�ՀwuՀwuՁ��f�x�ZİO'�
L�ɚ���@;�����2�;���J kޏJ���T�!G&�r�M�{)��3中��[�~W�����dQ��$�?w������;���;�����!��QNcSnC@����.[����h��M����A�Ls&(�@���Mu�ڛ��tH��d��]��yN��gU�f�����7>�r= ��٠~]�z��S@����r�z��G�x�RM ����jV���&+ ���F)Ij�Q��}�����9�s�}�����D8��<pcrh�x����;���1�Vsa�+�DPE$iBHh{>�����r�M���.[�4�O7�`�O��4����VCnl��,u����;�6us�k� '^J2ʭ&�Ë�0h��շ���[�3ezEۮ�;\M}�����l��,��y.$� c~�c\�8�l�p����M���bG-��r�M��k�|�Wh��L#��j(������j�;���s�%Isc�H\8�s�Mgdǻٰ:�x��](���1�Ϡ㙠��4˽�@���h�۹�s���d�<#�(ڒh�ú�ĹĖ�2��t� ��x�ߟ;�L�ev6��.���(���Ĵ훈�n���]͆��1�6�6�f���2�ݖ��;����ḿ�ܘ��@���(I�v��$��@�����즁y�[İO'�
Li9��VCnl��,�n,co5��&BG��94=�����9l�}���O_���{�o$��:�8�O�&ELrG�~�e4��h��V��mz�t��70QL���q��.m.�	��W�9�ȉcr��vƼn���I1G���ې�;�)�~��Zmz��S@/WlR5��Үn�~�s�����e�V�;� �jՠ~�k؜$�26��@��@��2�.qr#_�Ł�_��׮���b#���q��e4v�h��Zmz;k1kĠLRF�I!�s��`uθ�2s`nm2��.(�.�������z�p��"}��)1:��S�G�S��{ly�e�!��eY�s��	���8�Q�vᩫL������ӷQp��<ܓnXh����tG�ĵ��7fcZ���.a牎x��p��ꑉvݤɌ��a�+�1<�{�F.���z�����v��盵��r7��5�n�5���g:�2ur��@+���3)p6f�QՊ�Ʌ����yx��1����ggζ[X^m���u��Fz۴lD�m����z�i�V�ͷ���j�8��@�;)�w�S@����@���qhV׿��x�-��~��o�Ď���q��6L�I��=��Xs�,����5U1G��ě��;�)�~��h]��{��>�^��z��Lj��8���uŁ��́���5�,;�'��n#���Y��rn���ۭd�U�+Z�\��Q��WM��� �F�6��,�L�:�\X��C��ӏ@�;)����9~��Gd�h�ՠqvנr���
�$id�;e4���=�b]W�z�4�+x�	���țn��V���^��vS@�]�@����@���(�Zmzy�M�v��}�@��;^ ��0Ơ�X��$I�M�\�����μ��ڸ�gu����h�nf�4�ƣ�܏@�;)�s�ՠ~��h]���3>�H���I1G���䒋\��`wg\X��ݦXgl��7�n}�-�_j�?.���"xA>rP�@�R_@�� H���#
�x�x�)qJ�]���,n�`wu�37L��NE�~]����M�즇���/��o��S��ӏ@��2���e�ݝq`v5��23T�������c��Z�6�.��[<B���G�����춼�x�*GQ�A>�f�2��θ�;���.�cu������4	��Aț��վ��+�=��;�M����a0�)��;��ݦX�L�;��,�u��4�`��܏C�b��@�ӒO��w9'���1"B2$iZD�"��a$�h��>�o�g$���%�&(�s�r9�즗�}��.}�Ȝ�bX�'��{�O"X�%�߷�S�,K��/w������3�i�K�8`�ss�k��/S�t���Q#�g�rb�w75��M�l�-�߿w�{��7������"r%�bX�g��q<�bX�'g�ىȖ%�b{����yı.�~�?+��"��9i�ﷸ��{��g��q<�bX�'g�ىȖ%�b{����yı,N��܉ȟ�S"X����dܷ6���nl2��Ȗ%�b~����,K������%�bX�ϻ��,K��>�s��Kı>�vS���&�wr�wvbr%�bX���;8�D�,K��w"r%�bX�g��q<�bX�DfD�;���,K�����fd�k�3v�nl�yı,N��܉Ȗ%�a�X����8�ı,K������bX�'�}��'�,KĨU�
~м��������M�g�����)��k��e]e%��ܼ#kWmVM���Ǫ������7#m#���VJb����7l�fϜ�ݝ gm�_��N�s��T�Gbv8�n"[���K��΀�k�Խ�n�����nn^a�vHוyr��QH'&p�b��qnL�:�[98�nn�ٵ��a�(y@��!�D7�bsYt���.d�nM�W���'{�ۻ-Қuv�<�S�i��K�����8�w'd6��8��5�V�O<�Y^�v��;VY����,K��;�8�D�,K����,K������%�bX�ϻ��,K��=�;3nk�m��fn�Ȗ%�bv}�br%�bX���;8�D�,K��w"r%�bX�g��q<�b�ow�����a�+,���{��"X���;8�D�,K��w"r%�bX�g��q<�bX�'g��'"X�%��w�Ṧfɓ&f������Kı;�wr'"X�%��}��Ȗ%�`��y�Ȗ%��L��{����%�g�������r��]^�-;����d�<ϻ��yı,~�59ı,O~���O"X�%��}�Ȝ�bX���9{��0#�LQ��s�K�p�t�$.���ݺ;�\��M�]]eg�4�,͆\��I�}����O=�~�D$=�bv%�by�w���%�bX�N��7	�6���ws7S�,K��������(;����'�,O3��"r%�bX�gw8�D�,K���S�?���,O�~����.��ٹ��8�D�,K���Ȝ�bX�'��{�O"X�%��}۩Ȗ%�b{����yı,��9�2CM�M7Isr'"X�%��}��Ȗ%�`��v�r%�bX���;8�D�,�2'��ۑ9ı,Os���s\�l�3d���'�,K��>���Kİ������=�bX�'��ۑ9ı,Os��8�D�,K�o��K��l��\6��X.�^�vwnZ��&ή�:�b^nYs�&�+����ı=���8�D�,K����9ı,O3߻��T��Ȗ%��w���Kı>�����2�2fk�7vq<�bX�'��w"r%�bX�g�w8�D�,K���S�,K��߹���%�bX�w����&]7]ܙ���,K��=����%�bX>�ݺ��cA���ю�.!.逇R%D �b�R1�����O ���
0ayϗE��$��=}<|�� E�t�VHđ BED��Ü �� ��q�dI+!0_�f�7�MU�$H�Bl`O� �N(���TQ��R�AJ@��x���$$}�z�� �4C�b�F�ЊA`@�3�!�>��*A<h�w�^ECH��$�@�T(I*s�Vq���{�᧩������H�7�&`�	��@�>G"!шU���0|�2@FU��� b'Qb��Z�QC��}L��(��* z��E1:��f|��)~�؞~�ϧ�Ug�2%�`����S�,K��?~���m��m͆\��yĳ�@�?o]ND�,K߻�Ӊ�Kİ}ϻu9İ? �"{�w�q<�bX�~0��nɶni�w7n�"X�%��wÉ�Kİ{��jr%�bX�g�w8�D�,K��n�"X�%���>�~~s�V����i�<���4s����`�0��l��0<�۱���a�՞���8�D�,K�of�"X�%��{�s��Kİ{�v�~Py"X�'�w��Ȗ%�`���3�,��6�n��٩Ȗ%�by����yı,�ݺ��bX�'���'�,K���٩Ȗ%�by��;.��,�%�i�w8�D�,K��n�"X�%��wÉ�Kİ{��jr%�bX�g�w8�D�,K�ώ�si�eݗ776�r%�bX�{�|8�D�,K�of��*dK��>���yİ=Ѐ���"���D�>+U������bX�'��ߩ3�.ɓ&f�.n�Ȗ%�`�����Kı<�~�q<�bX�s��ND�,K����Ȗ%�b~����S��j�k��.z���E`zB�Z����eM��ەݔ"Ӳ����V�ߨ�%�b{�w�q<�bX�s��ND�,K�������&D�,O���br%�bX�g~��m��ٛ����%�bX=ϻu9���ș��>���yı,O���br%�bX��~��<��*dK���0�&l�f�wsv�r%�bX�����O"X�%�߷�br%�bX��~��<�bX�s��ND�,K����-����7n��Ȗ%����?w����Kı/�w��<�bX�s��ND�,K����Ȗ%�`��᜹I7a��7-ͱ9ı,K�wx�D�,K��n�"X�%��{�s��Kı;��lND�,K�,������.�V�ˬ�v��%�\��n��-��C�h#UE ��ځy$�8�2��� �9x,\�g�t)���U�Ѹy�tv�۴�۳��-���w8�Ja]=�H���I���Ѷ�8��b/�������}�B�oM�G7] #�aa	f�u��ˮ��:�M�3[����y���%q� ��GX�0l�1[]�6ە�3)�M�?�}D ��8y#���L^y�:wfwa��R����������ݠz�Э�o&���qW������X�������Kı<���q<�bX�'~���șı/�w��<�g���{������ܕ�f/w��D�,O=��O"X�%�߷�br%�bX��~��<�bX�s��ND�*	�2%���ߩ��3dɓ3M����yı,O���br%�bX��~��<�bX�s��ND�,K����'�,K����L3��e�q�ͻ�br%�bX�ϻ��yı,�ݺ��bX�%�ﻼO"X�%�߷�c�}���#�붴dc�o����Kİ{�v�r%�bX�߾��<�bX�'~��Ȗ%�b_>�w��Kı=>���&]�n�n\�������$&�8rL�k8����q������dft��͓l�ݗwwn�"X�%�}���Ȗ%�bw��؜�bX�%���x�D�,K��n�"X�%��w��[%�]ٹ����O"X�%�߷�brQ��~���>>��%�y��Ȗ%�`������bX�'����'�,K����9r�n�i�72�؜�bX�%���<�bX�s��ND�,K����Ȗ%�bw��؜�bX�'��s�6�f��6����yı,�ݺ��bX�'����'�,K���ݱ9ı,K�{��y�q������K~w�I�nqX�bO"X�%���gȖ%�bw��ڜ�bX�%���<�bX�s��ND�,K�
}��L=�v�a��m�q��]���f�lH���`��O)÷^܍��VS.��&L�f�777<ObX�%�����ND�,K���x�D�,K��n�"X�%��}�s��Kı>�?6\}]>�&w��oq������x�D�,K��n�"X�%��}�s��Kı;��mND�ʙ�w�~~&5�i46p������oq���n�"X�%��}�s��K�_9^D�S��GC]=��O���Ȝ�bX�%���oȖ%�`����{6Ѧ�U���7���{������<�bX�'~�6D�Kı/��w��Kİ{�v�r%�bX��~�B�.�˺I����%�bX�����,K��#����x�ı,K�w���Kı>Ͼ�q<�bX�/~�{n��Q���q�%��U��k8d0���Uں��$b��%&^a6��:U�ND�,K���x�D�,K��n�"X�%��}�s��Kı;�y�'"X�%�|���6�)st˛���%�bX=ϻu9ı,O�ﻜO"X�%�߻͑9ı,K�{��߭�7���{�3���jg��V)���,K��>����%�bX�����,Kľw��'�,K��}۩Ȗ%�bw�S��7Hf\3]����yı,N��l�Ȗ%�b_;��Ȗ%�`�>���K��F'�@�C�7�D��
�t\�O��}�'�,K����	�o77.��˻7vD�Kı/��w��Kİ�V����Kı;����yı,N��l�Ȗ%�bu�{|����a�b1���y8zrT�z�2�9�v�x%I��Լ�Ɉ�i ma��߭�7���w��u9ı,O�ﻜO"X�%�߻͐?șı/��~�'�,K���c���ٶ�5�k^ﷸ��{���>����%�bX�����,Kľw��'�,K���٩ȟ�2�D�=���m-��������'�,K������,Kľw��'�,2&A���59ı,N�{�8�D�,K�w��!��K�36D�K��(�2&{����yı,���S�,K��>����%�bX�����,Kľ{�ٛsY���6����yı,�����bX�'����'�,K����Ȝ�bX�%���<�bX�'N����3HM�f�Y3�3,۪:�4V{�v";w��!�󂝃�նu��*Z(!_�t�ƕ�%�U8��//]��Ǯ
<�.��nDE^��0�A�c����ݸv������{r��svl��W*[�y (
�NOZ�Srڣ���ɫ�B��,[L`#��Ɓ턷aKGu�mɭY�uk	�tABu��\B�W74s&���>A�h�p�=����i�Z���7lH6��Q�ex�/�֤�(Xܳ��s��*�g��))���{��X�'�gȖ%�bw��dND�,K���x�D�,K�of�"X�?�C"~��~���C2�����Ȗ%�b~��l�Ȗ%�b_;��Ȗ%�`�����Kı>Ͼ�q<�b]�7��~'ᔙ�����ﷸ��ľw��'�,K���٩Ȗ%�b}�}��yı,N��l�Ȗ%��{�����f4�6�������D�{��jr%�bX�g�w8�D�,K�w�"r%�bX������%�g؏��T��p"#�R9	�i�#�BX�g�w8�D�,K�w�"r%�bX������%�bX=�{59ı�{���{�?����Y|<^C nm�qp'�e�2�`��"s�{��m
�N֚���f˛$���=�bX�'���Ȝ�bX�%���<�bX�~���O"dK��w����Kİw�˖Cvn�ffl�Ȗ%�b_;���@@늞�p,<h���
��E��dM�`���59ı,O��߳��Kı;�y�'"X�%��{��͹��J[�s3wx�D�,K�of�"X�%��}�s��Kı;�y�'"X�%��w��'�,K��w��Ls;��׻��7���{�Ͼ�q<�bX�'�nv��Kı<�����%�bX>�����bX�'ݓ�;ᛄ30�����Ȗ%�b{��mND�,K��{�O"X�%���٩Ȗ%�b}�}��yı,Os��[��y��=+�V��mt�ۧژ�Ö��F�*��٥�)�sWE��Ȗ%�by��s��Kİ}�{59ı,O�ﻜO"X�%��۝w��oq���~?�����i m����%�bX>�����bX�'����'�,K����ڜ�bX�%�{��yı,OI�i��.ɶni7wsf�"X�%���{�O"X�%��۝�9����+���`@C��=�y����%�bX>�MND�,K�w��[.��74�7s��Kı/�gv�"X�%�{��x�D�,K߷�S�,K��w��'�,K������݆ۦ���ڜ�bX�%�~��<�bX��of�"X�%�����'�,Kľ��ڜ�bX�'����L.g���1�$ͺ�d��Ơ�b��Ƽ�j�v���n�9���4͹��J[��sw��%�bX?wMND�,K�߻�O"X�%�}�;�9ı,K�~��<�bX���N�L:sP�Z�}����oq���~_x�PX�L�b_��ڜ�bX�%��wx�D�,K߷�S�,K������f��.�.nn�<�bX�%�����Kı/�����%�@V �����Kı/�����%�g�����O��b�蜴{���{�� dL����'�,K����jr%�bX�����yİ(!�C
�JD ?�Qh"T�y���ND�,K����,�L��f�ٗ7w��Kİ}�{59ı,O�����%�bX7߻���bX�%����<�bX�'�{��Iwsl�#�/c2�p�Y7=��bݞ������F�X�X��uۇJ�՝0��}=�{��b}���'�,K������Kı/��w��ؙİ~�����bX�'�~�il���3v�n�Ȗ%�`�~�jr�#�2%�{����yı,����"X�%��{�8�D�,K�����݆�ɹ�wsS�,KĿw��Ȗ%�`���jr%�bX�w����%�bX7߻���bX�'���;3nk0�%��77x�D�,��@�?w���"X�%�����Ȗ%�`�~�jr%�bX������%�oq����8�Baҕ5�w��ou�b}���'�,K����w�h�	"w�jr	"�{�MA$O� U��D U��" *��" *�W��@_�A �" *�Р�!��*@b(��V"�1�(� �Q��UH* � � �D"(
�1`� �"�0R
�0"�1�	?� �A � U�" *�W�W� �
��� *�� �� ����
�� *��� ��� ����
�2������R�����9�>���   @                 �5l ����BR�"�	ARA@� ���*�J� U(���AD�����$��PA U�    h  @   0Z
2�}�o^U��޳�]�{�ͩ��} +���o�S��V\ڞ{}��� ���( �     P��L�X �@� '@� 
 : "@ (` @    � $@� �Ġ �
D  �J A�4A� (E44�h�� =�U�p�.Z� �嫎��@  @y@  �M�/�wO68�*�i]�T�W�r嶺�s�3ɪ�nMK� |�  T  ������^�֎1���''��w���ol���Zrz^�N������R�n�=��� 5޷/�[Ү�}ꕋr�9o��&����C��(��}��>����O������7�W���      �@�O��eշ'_^���O'����9��sg����׽�x�{9:x�G�ާ�㷭�}�s� ��;���n����}>�7*w=�W� rb0@{�7`q�}5��ק�o|�� �      (
a4 ��NO��/�{����z^��ojn �={g&�Y�_^w����x��=���|�����o{|  ���<�ǝ����-�}>��]y���y�/''W�����nZ�6���ܝ�y���_ ��*{iJ�  �)�����J�  �=U*Tc@ d"{J�RUA���hb*�Jg�R�  �!JSH����߿�����������N�s��u�J���B���UU�*�
��UU�eUTW�  
�UUN'���(�FG�5��#0�H���0��2�#33��%�SxQ� �!$F4���sS�h�k� ���F)�
�d�e� \ѲL0�{�6��@�(1�4�$!I�M��,m�k��L��yO!w��ST# #�F&YK<C��6c�J�Xka���n�!L��$*@�`�(�(b�0�6I�Ѩ�Ȥt�"�5����G`�@`�����$ă�i	! �0�p�c����$�b@� �d����\,�i	�CP��/.h�hA�a	
0 �s7.R̬�F���#�,�)�F�22�0�nf=y_)HbB�n>B�"h����%u
,!5�2���Ip���.2��@��)�#$!@� R�)B�X�+
\YBF	q�nHWS1%1aV4�ۨm�ad�!���$ChD"�"�#�����y.j�2WH0�L	��ޒ7���̄��KrQ�50� @�@c$`��a`Ii��4Cx>lv$ Q��1-2\8"$R��!��Ɇ���eޮ���o���l)�L)�5�4�Z���|�$��\�ۘM�V@R�zV�h�B��ԗ�g�U�$�q���F{�O�a�I-y�>oNjZ�oz�RHH�t��H�=���¤1�h��l��w[/����q#R�H�5���OR,$�I"�
a��.��B>xkØ�r�zkzvba"F� A�d��Y� ��ƶ��A"D�i��sZ�������iMɰ��.��ƚ��]�w���0*a�{��Z����^�f��5�ÜԐ�;��c�~sW�\������#f����;��s�a���HK�HԐ�"d�1b��B�XCp�Ӣ�25g�k]��D�.k�:�M�zf�RZJX�#�(��O�3��tS2"xG�$�HNy��\Mn�kyn��ߗ�o�y:�=`m�+ۧ6^oz;�bƒkK.�p�<	��fC^j��(�d	!K �ޡ��o~r{��G���$B�
�`�*D�F! Z��AH(@`B! bD )�{}ߐ$��욦�\��6�	�H��D�BB)�dd�l�l��*�ƬX��h�d˹���B@�!�pIxJH�R1`��X�R:sRn�F�4�ٸ��;��%����G����āM��l��<�
bƉxA���jdH0$cB��K��s̅�6ka5���"f���8I!��j������n��� Y1��$�Y01�6z˓Wd�˝}y"G�$O&�g�S�!sS��5тP�%�\��7H]���%�5Bm��N^�i�����{|�.h%���-�"4�g�x14h�JB� !"Y"P#
$R�LSLf�L�k��7��.d���C��� LMK���B%X�7�cHԍ"HV�%%4xp7^�̉^�q�n\0�E����sV�v�ox�e��7�y�ysa=Ѱa��5�-�F�yM�f��j!� S!N�noZ	�$
F�H� ���L�{ר��Z�`5cP�HV]��B���H1�6��	 �~u�O)��;�B�5�
�@($l��%	a;t��oiw�W���rC��D��E�!W-0�g��C��%�ȅ d�!2hֲY�����s2ђ��Յrj_9&��ndp`R5 �B$h��F�o}Pߓ��Vh��B1���K��q/�{��4�HE�)��#�g�R	ԈЂ��3�פ�Y���5�a,�)�����{��}���0"R]��fk���v�A�A�A�Y�	�� �� l�I	�H��Z�a>-+F$Cy�r��7�<�5���a���{a0*���l$
&#
�@��(`h��@�Y�$"������0���Jq��M�lS��0�!��4�ۿxn�5<�N]p�!�)��j5B���ƌ�B��dhL�.�i�%dad�0�aM0�,)$�+0;����F�hA�*�+Ō�Cl׻�KRJB��F�\H1�xx��t���^A�(�����xc�$K�p�0�0%�IR7���0��Z����.kG=Iu��5`]Mfy�k�Ք6� u|0`� P!S�Ġ�Š��I �@D+"A��4�����M��x�p�j�P��V� �� ��,=�-tx��9禃3^���6F�H�b<$R	�H_e�kO�d$$Y#C$R�����xp���p�%�kf��)ŖP�r���9+
��8�Y뱺�	f�fe3��y������Lp��La̩+,�a-���gx��H5hS|<����68g��$)��#B5��HY�+�.ˆk�Жg�-͐'��k��q�|�}<��HK�`a��FGRB�B@�0�k� S�>뤥Z18��yJd.1�Y`V-i��#GF�C��7����'�o�]k�l)h�D�Æ˭llM<A������1a��!@�!Tc"���d�"@c���"�@�1H
��A`�jD�A�
H�$�g-$`�$X��{�i��,JH�J�
c��1��#�Q�3�!Lr�eÎ�M�R�#�I��)�MJ*��q��i`�BB�!!,�:Gi�k0�CP�(����\t;"Icrf�ۘ�ӗ7�u�o6j�u2��a(�4���FH�&H�HH��ᤒ\ѳ��HD�I	���Q!n��K0�[`q���j�(1B$K!$k �L��d�q�.���m"PO=��Z�!Q���]�N�������ѾxY����L%�2�_vxn����u�FHS#S�,6<NH=u!A!�cA�,"D��D��P)�jH�Y!Ie��1�#HML�<�@��jŤv
"z��6��0 Y},
�5�cX�a�aHX�4�tB��.�Й�OH2BVXq`@�HQ�H����ޙ�]oV3�q%Yc͑���p&v�s��䏧��d��H���	b��ʹա͞�C�&1����Z5��Ɖ�$�!=�,����=�j0�͞q�x��g5�!��/=4���������g�5�f�)���CE�-aZzā"�,l(@�,a4r\u�+M95�{'����!\��CW0�� H��E�r����׳�c�5���bA�����3�F>�	
Ǉ!�xor^Irh����6�/5����p�~�7B�>;�
�#q'}�}�q�q�H��@�0�/J�V󇤹����j��nH^뎭-4cY�$c��L)���$!����Jf@�R1�2��F2�Ĭ"�R�ZҐ�$�A.Mj�S!�db@�V4���]C2I%��;��c�Rg���n��-f������,�}��7����O]�Qn�:���k=���d�i	I!urI�2�p�H�WC[BP�5C1�u�r���0�.�me��˭�Y��幭y��{��A�U�g�!�iX"즦{���M:��3sw9�:.o�.��Ŋn�8+�_�h=*_���w�A>��oc�����~��}}ݾn���o��8���.i.L�����~�{�B�k��±��k���S���@�%b$]�K�|�!N�XG�<�Fp��'c@�G��(B�%7�wА���\��r�+L�@�b��͹�X��@�4JDć���0�I0ŅL=	q%�4zk\�'���a��L!�!���4]�L)��Hs��z��s=�{

�����)��/���F��3~��L;��p�&k|7����a�hB�!
S'!��Ӊ$$JF��Y5�A�`����1),$\�Ӑ�0ٮ>Da	�B� � �E4a�'�I y��*�!!�A��D�M���́�.H�f�1����������:�����XfK �
�I$�G��  -�ݰ  8����   �[l  @ �` `�UUյ9yn�v�R���� ִ�\1�C��5�k�k9zS��w�m'` 6�[}f[�;m��    �oj�Fq&�ڑ����7M�ʓ`(i���5�  ����Y�ڶ�!�H ����j�6�K$�^�-�UKjvZ]d�%�H�ŵm-�m�6�`���
-�����8�vM%�l\�S��Hl�M��ҁ�6�� �  I��E�^r��[Yh�.���"��P   �`�k�k��lT
�55̔YU�Ua���i�E�c���-5�kXڐI&ٺM�-���nit�i!;9�km���g 9@��V�lJ�m[mvհqr�\-�(Vg�wl<5v66h N��J'��������i�ܑ�[�Y���ŗ��[dZl ��
��Y���6�ئ���l �`[A�ck�V�{6��J�O;-&̜����i��H �Ω6��v>H���ۀm�$85�� �d��p8'	�.��y�fV�[g�vX
%t���gT�K+��ڨPm� 5k4���_�I���z��KV�GKג2�
jA�g���jU�MU;˰��e2�6��_�]|�J�hk�Xa�����H B�W�Ґ ���j�Y^�\Us��KKmU*>ת�`���+�糌m;5+�k��Լ�ª��+��� H�H$�n�M���U	�eyڪ��eZ���*ʁcMU[T�*�U�
\��ҭUr��]K����U���y���9�U]V�� ʠ�$ W�|�߶�t��,���}�m $ku�� p�tݵnY8R�벛 �&�m�e�Üm sm��k�����D��sE�l4+eA��ڨ)@u����m�n����!�5���kn�BL���K�TfYʻ��uت� .H��ysGY�F���:6ݸ�Wn�� N����,�[R�����!��˲�=c4�3J �kimdk[�8�g��`%X *���	�4$gI��m���0  [@-� -��@!��l(ҷ<�m����*^h�pm�T�UX�&׃m�m���ũ��鵜�͛���@ �׶��h�6�H�lX��Z�Ͷ  ���@@��dW\9�������S���Ā�H�mgi-��!  � �  8   � 6� ��i�;ѵ����jL  ��(6�3��%  ml� (l  -�-�m��>p ���@�*���m# m���Z@H�6�[@ h�` 	���i��  ��!5 9hહ�j٪�"�< 8�d��S�Vs�T�
���@oR���v�꣌���+m;+��s�C�;@
۵
U�2�nSH��KM�+�$����   �hXI��e�K��5ғ�]�w�`)8�j�Ike؉����8��c&��C�
�WIM��T�MU:.�. ��s�����;
�2����������6��pz0� ޠ8�ԗ[�-���l�Y�ksLn��J:��8ѝ�ـ��`�e^�bZ�Cf�ڷ����r�㍖�$���N�צ�Yŷ06]����\�2,	L�Ff		���V��+n�r���Ttd޺̹"�U�+m�<��q�mS��]@*�u�̀]&ɒ]9�Nu���ot��Y�`[VXI�l8	:�\��G&�d�X�U�W�k��"V��a��[� :ƽG6�v�v�*��zRZRL�6��6st*�UU\�e�v���a�����a��quT�PT}/�o��6�6�]��  6��tF������Ò �a&<$������[��< ;e�X�K���U�c��e]�������i   	��;5 �-�U[m �r�f��J���m��d  ���::�T �甭�� j��bճ��^UweP}<��E\Լ���{eqĈ4�K�||}US�y�H})|V��l�'��J��`A`�l�IX �  ��Y/�m�m��檁6+R��YFkR`�      ㄀ � �  	 �t�    m$l�   �������l��6�^�$yh]6���v�٠5�++UJ�Qa��@m��    	 [G� X` UU`�5*��@c=�v����P Ԅ�KR�m�]ͤ� �6�����-�����lI �H�YA��a����    [V��i6����]�mm��ɭ ���Yڅ��8�&ԍ�oV@%�Hl��H<�.�-���
����p �UP
�D��zݶZ�g m�:*��R��v������sm�    miW��$�3m3 �Uq����F��o	  �8m���Ie::C k�N^L���.L[:�>�}�}��庶�j�r�T�pq�`
��Z�1�o84k�����v[v��ٻlQ�.�,�V�kl�$ְm ����ayk�VVwk�A��m�[֓cv�  �vJ�^����( �Sl��ʼ�7��X+f�p!������Qzi8Hj�M�Ie<ym)V��UZ�	��Wv���!{E\��5���+g7|/}�,�:�����j�x ����ҭQ�*����U�Z�U,쫻,j�����ŻU��b��d���,Ѥ�l��̖к���-��u��[d�� �&�3��Q��kl�   k�[R�
��e\�,T�*�	v��<��]UUG+4Ѝ�.�V�%vҊ�:N  m��v�#b�g�`�JԬ��Ѹ5r�-@UUu��b�$2�U]R�l�PpZ�ͤg H�u�6� �`Յ���꽡�f6�$-��ܕpmUP
�	v���@��*�5UU*5��mR���� ծ���}3��H��m���]K�)EU*���.�rgi�Wf�yeF���[�Y�mm��@�J'��8�m�Q�n;e�uYћ���BV��^�B�� :�eD�okd�  i�e(-�8����m� q �m �-��H*�1��J\KR�ʰU*�qUԖX��h�
ܫA�­!��T��@m ��W�\��a:]�+mQ����P뮶޳��6Ӧ� ���K�  $H�eK��.�ꪹ�KV�pq��㪮�vF�Vsh73[7gFE6VTVd%u���W �e�mZ�#j볡�)da�h��j�Iӂ�Z���m����*���Uy�ҵ*�/J�m�l  pp$i6�WV �@ m�4�1I[l��8p  H[Cj�� �nEӶS��ʺ�n�T`A� Ѷ��6�j�� s�@�z�@շ�P,�K m�հm�m��඀ m&��m ����	�,6R�Z �ɴ���M�@m��hjq��>J�V�ꀤ��7eڪU�mt�g�`	cda���H[[lg�Z�6�L��ٲI n�X�y�i�������Z]K���`/G0 �e�Xl�kWQ��HM�h.���2�]V�	jع��nSv�`hm�i6l�   ��`6�`p6� Zl�&��ԁ���ZĲ��[@��u��VP\vݜ)�{u5d�hr�x��]l5@���m�J�t�n�Z�]SʅE�,-76�R�K���i@�q�ҧ�1 ��k��m��D���gH�&N`rti���8m�2  ���K&[]m ѻ:��tH7*�m��eu�r��xܠ]9�[������t����F���m��8���J��
���\�7[�[�zm���ؠ
�Wi����n�6��n�P[M����}'�o�K);k���ݶ�d��״�Ü���f�E��-�M�	��m��[BKn� Hm��5��m� �l�/P�b�H -�He����`�0p�� ����%����U�n�N�^�;@P����H	�A��we���mӶ�`� �H  d�  X`-�m�l��M"-��hղ�h$���>-� mU��Y�f��jћM���:'n	����-5�r츺�Z�cQ�f)v�X�f
����,���6���C�PQ-U%��V��� ,]�E -�t��0  ���HH˳6��}��ie$8���l$ @�`pp  M/jl6ؐ m�l.�On6�-�lp8� Zl[A���`:�m���'  	�kn�6���-��&�c�Z��6���ʪ�+UU*�R��a�`m���ᶑ��"�����h    m@ma�*������[U[�ms#�ț-��b�*�yeZ.�h;m�Bb�$��UUT0SWC�~A<@Ѐx�TS��Q�+���SO�H�F.�"� �o�DOb��҈����`�D��	F��k�*�$����]�"!��@�A��*ixiҧU�GOC�T�"���^"�@�xD<�"�d 0Av�J<E�pH�*J}Jz!CN�A��(�(z�Q ��AC�}V����UQ�� �@^�xz
�B"�P����۠}B�bTu���J�*�/A�����
<�R:���*��uQ4�XT8���|��_`	
�4�@h�C�z=@ؤ�HJ�9����``�8z�2�V$! �T��|N"�WJ&�A���P
m`�TX��P�80K�u�툏�������G@
A��=OQ�`x�Pt����X�S�T�:�^$�ذDH� b�#<C��S��)B��HRE���;�0����i1����,B2_��$ �R����Q 1�>�������N�"�:@*��� iP<B#���)݊���_�HA$�*ư$��J��Aiʧ��H��)�(��(u�Wa���^#� �
���Z"�A�@�/��  lR"ࡠ���lU4�*��QT ��������uGh�x�pi``�C�)V�
&L	�5ƠRV�QOf��w�[u��3Z5��[[UT���J� �����%.Il��^׆�d��c]�%��:�qm�Z�r11�&�^K�ף��V�v��P%��2�N2����vx�q$�L�k)�@��\*���%��͸���'�PDn���ˋ��n��s�R{9����%�����Y�ݡ.pu;3�5��"���,�6+A�Gk���6k9��d��'�Tvy9^Kتނ�F���5)�!�vh
�tnUM��{VSv;K�L�n��*�<��ت�M���%*��[B�t��`*PK4ԪJ�U�܆ ��Q�yt6c��*��t\�$
A�L�tn��b���bX�C��7�Yi.�ϳ�g�əWy�e��ku���V�npU��2����gJ����t�u���9NU��@�:m��,��學�b!��cm櫤�=F1'����K�J�t�)m ���M�B���c# C��$�R��*��l��.lv�^H��8j�CQ=�.ʳʎP:(m��0 ���arf���Xv�:*�c�wKۍ7 �:�n�qݜ��\��A��$�֚�,����L��/nd�t'OI�5�n�E�ó��kg�4����̡�;%��v���k#���S.7=3Ƣ������%r��q����P�wYb��<�m�Kg�PqL��9)��c�n+vr뫈�mӮ�#&*L�]��נ��뛧�z�5M!s�@�;Tq����-��ũ�����;C�V����1�f�x4��=�e��0Nq`��Z��V�J[Wf�z`��C�t��Fd�pc1n=v��.�.�8)�w'�[�κ�;�6tO]��Ujl�>��9:֋؂[����v��+O�%y^����-v����`�����j�;d؁��� ��{��ϋ]�>�����#��W�h�UX-ڱ��R��%^�Z��Bf��*�U+%�9�kR�Z��I���)�#�$c�A����H+����W\�U�OW�@�"����اAN���US��D4#k ����L܅���3Y����ɜ�1{mg�]h-"q3�WKmζ�K/��a���uqu�	ծ�y�a�G=W���Qџn��Mn'b�q���w\��<�ݗSQ�����I��lu=��ogL�RQͣ���`�[.TI��m��7imqӴVK�{FR�6B��m�tݣ��WGF`�Ux"���֘{/�x�0���&ac�-֬��U��G�9���nYI%��˄�̄�̛����
0;l�r��,b��1�5�?C���@��� �s���߳��4b���Ǎ'"X&����)��U�7�P�@wd����W#�Ȉ�lNf�s���vS@��@����/i��G��m���=�`���-�qRU�]�vh�ci�����!�s�ՠ~��X��X�m� �J"9���l��Q.��.��g�zSD	C�E��8�����q<��Y9ZQ�ͷ��ʐ��@{�� NsPn]���M����.�`}���KyD!oJ�@�aM!��%��)�<EP��D)I4�"L�����׋@�*�(�xDd��8���M�{^�K����*���9iq�Պ8,����?K�YД)��� �_V����9����4�����;w0�k���ـ~u�pJ$�U���Ź��^����P&.�f�J��7X�1�t:ٌ�:��#%���֝�;�H ��%���@zc���8���D�r)�G�}��hWڴ�׋ ����P�S!�˦�����0�]jnI��߮�����Q=��ID��	TD��k��� �Ү%F��ick$q�s�s@����vS@��s@�itJ50m�$��� $�-�6	T�m�H	\����������l��95�='�+j��r-�v�gsBn�����Oh�>V�m�6	T�m�H	1�@G�2T�Y*�JUwV`�ŝ
�~��=����e4�uw�<iGE]��7u��׋��}�|`�x�:��+28̘�k�h�������0<�����(BS)L_�>��k�k�lܓ���٩��WY�3ov��6��`����T��۹�r��V(���A�ԃ�!���T��ؗ�B*w!n�!�:����P��*��9���9�_��a�zx���%�7X��Hh�b�� H�9���U]�̈J50m�$���h��h廚{�~KݳƁ�_nh�Xe�"2?͸����{��`���<������cU*n��u%"��`�l�:��ߗ�;_b�7���*"DT(��A`�T{l������[����w���us�*3����ys[s������r�SĐ�9z.����ʲ���nH��:�׃�(n/XtunM�n���l.y�5�Qѵg[���P�N�'������Z�t�v6˞WܤT����M���r�֧�w]�WV����)��;D'q��vM+\��s7��mʬvhwV�홅�h;Qr=J����8���{��ݝ��?6'u7K�0�-r'L�b��ȝfDd����қ<�;h8��\RHi��[������� qRs� :��K��5�mcNf�y۹���1"��s@�l�w��h�n�B(�3ov��6�T����*@Ns C��s5S7U4���Uk�DB�ל`{�`��`z�`�je�yy�e�e�{���T��qV ����D%O�r�����4UZzi��}Y;tG`�b�c��qջm�b̏�|�ԉ6�ؤ��L�v�s@���h�l�	/�_b�9�B�I���Uf�hܓ���7��F�U��`)���R�.���q��G��`ϱ`��g(��ɼ���4�#C�I3@�l�w����n�����>���V5Dq`�F�ДK�ߖ����ŀ?m� �+2H�LQ��s4���ٜ�����4�s@/3���Q5�N:n�&{I� Iю��Vqj땻{gi���cң�"B(�R,I��>����v�*@NqR ��K�˽̼��4UZ��ٝ�G��p�ذ�n�g*W
�Cd��
C@�j������%
T�!DlB�Ǚ� ���h�K�7��6��-�s@�qRs� c����Q�V�ٙ��HG '=��9h	��h����hNd��Idɉ�+�l`��mV۩8���Tl�����Ũs�mh�ۖe���q�H��qR����.�ⱨ�#�ڒf��j�qR��T�}�]�`�~·u���k��/��4��M��s@���hr�d�r)$�h�gf����ܓ��{w&(n�Q�U
A��1���nI=��t��2�&Wf�^,�B�;��>}� ���@���=�l��ȜM�~�D�"H�-�3��bZ�j/\zm%m�:�'�ݧ\ ��2�7Y������T��=��hv�lM�j5	���s}�\�<���m9ı,N�~�Sq,K���iȖ%�b{�i�]ɫc����&�X�%��=�fӑ,K���]���bX�'<�}�ND�,K��6D�Kı9��a�!��Mf���ND�,K��vbn%�bX����m9ı,N���q,K���iȖ%�b�o�wV�-��R\5�����%�bs�wٴ�Kİ�?w���,K������Kı;=�f&�X�%��ث�J%A 1HP�2�fk0���5�aѭ�;:qh�J�.N�]"U��v�rok&��'*Bv�a�IL=3����2�Q��O�.��N���wE�qv��͒�F������ 5X܍hy�����9�&�=v�
����z�O[U���k�ky����qg��g
\`_\�I�GW]ri3]@>7N9:��V�]3ֆ�N�rx���ЂN���������]�4�9\��^\�:̚�.���$�H�I��t����Kb�ِ0v���9Ս�55�֮�4j�e֧��Kı?}�6D�Kı9���r%�bX���q,K���iȖ%�b{=���h��E�����oq������ͧ"X�%���17ı,Ny��6��bX�'s��"n%�bX���gN۬�Y�	0�5���Kı;=�f&�X�%��=�fӑ,K��{�dMı,K�{�ͧ"X�%�O;oI��r���fR]jbn%�bX����m9ı,N��D�Kı9���r%�`uVdK=�f&�X�%��{�9��\�����֦ӑ,K��{�dMı,K�G�{Ϧ�Ȗ%�b{��Ҧ�X�%��5�nӑ,C{��?߇!����f��5��/(�I�u�'�tT��k��ٽ+������`�c����D�Kı9���r%�bX�v벦�X�%��5�n��y"X�'s�k"n%�bX�w�r��іa�����Kı<��eM���)��E�Q����R
$@��Ub lS�Hؚ�b{�{��r%�bX��{����%�bs�wٴ�Kİo��;�u��f���Y�ԩ��%�bs�{۴�Kı=�{����%�bs�wٴ�Kı<��eMı,K�'���kY�M�����r%�bX���D�Kı9���r%�bX�v벦�X�%��5�nӑ,K���n�5�5u���WZ��5�7ı,Ny��6��bX�'��쩸�%�b{���r%�bX���D�Kı>O�{�G9?z7$�P�ZJ�m���pkD�C-uũ�rݢ��y�砐�{g�kq<�bX�'�]}*n%�bX����6��bX�'��u�7ı,Nw��m9ı,Jy�ܚ�2噫�̶]jT�Kı=���m9��DȖ's�k"n%�bX�}��6��bX*L���J���*dK������.]Kr�	sZ��r%�bX�������%�by���r%�C@Tā�=ސv�Cl�R��N��� �JJh"�*�H�$) ^
y�xI��"�q BR��T�2IK�M���S�h ��{��cYI�4����q!%�H�h���Ms'C��!�B��!0 ȉ m��6>�Ge)K.�y�R�Q�p�C ޥ!M�޶Ѹ������H:0/6v�������T��*q�I��<GI�(2�� ��`fB�F�*� <�h�<<H�x�JK�;�����\d�21�`�#5����᭜�dM�!�Bn�@4�'=��qD�Q�C�N��*���W�-b�A�&�<@�X��x-<A�z"� <0��'�L,MD��_J��bX�'{���ND�,K���I,�j�k��f�&�X�|�"{�y��r%�bX��u����%�bs�w�iȖ%��u���Yq,K��߿\0�5u)�,�33SiȖ%�byۮʛ�bX�1�����yı,N�~�D�Kı<���m9ı,O�w�}��Ys&Ir��4d]F��ݞ�۲g]�<�-��ܡ���n��J��؈�Ad+8�M�w�{��7�������ӑ,K��=�&�X�%���a�_bj%�bw���Sq,K��$�~��ֳR�5e��j�9ı,Os��"n%�bX�y��6��bX�'��쩸�%�bs�w�iȟ��MD���o��>��Y�S���}����bw�o��r%�bX�v벦�X� C"dOs���ND�,K�ߵ�7ı,J{=�;n��f\$�ۚ��r%�g� @Ȟ�w����%�b{�w��r%�bX���D�K��x	�J�@�DX�	B���Q?"��wٴ�Kı/ݿ�K���1��{��7�������~ND�,K
��¨���� �	�k�ؒ	"s��MA$y���am^��X�x����6l������+�cp2UÇ�r��w��>�7мf'�4��Kı;��Yq,K����iȖ%�by����r&D�,Os���ND�,K�}L��o5m5�ff�Yq,K����i�|�ș�����n%�bX����6��bX�'��u�7�~Mbj%���߮r��іa�����Kİ=��r�"X�%��}�ٴ�K�2&D�w�dMı,K��M�"X�%�}���[��n�	������'$%D-�Ȗ%�bw;��&�X�%���fӑ,K��߯ܩ��%�by�vq�Wud�W$��]d/�)!I
H[Z��Kİ�!���~���{ı,N���Sq,K��;��ӑ,K����w���Ren�vv�v��q3�RB����[ȃꅪ5NSn�s�\�ji�w��~s����e�0�����^���h�9�^�2����,cD�\�;B��v�8�ճgmٍ�ᣝ\
���ֽ�]fآ+�6�Z�6���j�ݩ*D�mQ�3h��a#����WgPM�\[.�@U���sh^�m��4�Bp���Y]�Jhgv_w{�����{�ݻ��}�޹�K�ݢ�EXz����a��\�3f]�z��ͣ�5n�~�>�~Fr�S	�kfk"v%�bX����ӑ,K��]�7ı,O3��l>I�L�bX�������%�bS������u�p�nkSiȖ%�byۮʛ��G"dK���iȖ%�bw;��&�X�%���fӑ>S*dK�����y\2���ǻ��7���{����fӑ,K��=�&�X� ? �5Q>���M�"X�%���_�Mı,K���sW0�5mˬ&k3Y��KτD���&�X�%�����ӑ,K��]�7İ>@BdOu��fӑ,K���S)%�z���33Y����%�b{�wٴ�Kİ��~Qk�ן�O"X�%�����m9ı,Os��"n%�bX����!����< 78�#J����j�s�V��S�*�+�;gqBv�����������tX�<�jq<�bX�'�]}*n%�bX�g{��r%�bX���@�+�D�D�K�����6��bX�%��g�[���S$�ՙ��7ı,O3��m9�)�1���\��,N���D�Kı;߷��r%�bX�v벦�~D?"��5��'��/�Z��ѫ.kY��r%�bX�gߵ�7ı,O}��6��c��R���>����q,K��>���r%�bX������tMg�OK;����o�wy��;߹��r%�bX>����q,K��;��ӑ,K����ț�bX�%;�>>�Yn�.am�jm9ı,;��&�X�%��w�ͧ"X�%��{�dMı,K�{�ͧ"X�%��;~���jf�˗D�j��n���7� :����"����ۀF���c;O(�^W�)����oq�����_��,K��{�dMı,K�{�͇�'�2%�`����7ı,O¨����y��Y����5���yı,O��k"n��L�bw�o��Kİ~��t��bX�'���6���)�2%���S+-�Դ�9���dMı,K��M�"X�%����I��5�:AF#hT�"F"��D���8� '�DȞ�_{v��bX�'���ț�bX�'���9]Jh�0����r%�gʐ2���I��%�by���9ı,N��D�K��BdO}�>�ND�,K��Ϧ���Z�%ֲ\��n%�bX����m9ı,?�+�~�D�%�bX����M�"X�%����I��%�b~��g/֖��sUdI�3T��m���4ڹ�KjE��T��v?����}��2�Ll����%�bX����ț�bX�'=�}�ND�,K��n��Ișı<�s����$)!I	�Ӗ]Z����]�E�k"n%�bX����m9�~P��j%��>�t��bX�'�}��iȖ%�bw=�&�|��2%�O'ӧ��-�fL��֦ӑ,K��;��n%�bX����m9��PdL��w�dMı,K��M�"X�%�w���t9YSi�����o�{ܰ2'��>�ND�,K���ț�bX�'=�}�ND�,�"���� �t���Ga���P֠�|��7ı,N�߬�afjۗXK3Z�ND�,K��u�7ı,>>w��m<�bX��߮�q,K���iȖ%�b~A~,�\�g� ��Nxc�g�U�^Mp��\7j�L��p�Y�����'��w&�G�X:|�3����ı,O~��ӑ,K��{ۤ�Kı9���|$�&D�,O��k"n%�bX�{��95.�2�2�jm9ı,�{t����uQ,O{��M�"X�%��?~�D�Kı;���H���K�����n��]k%֮�q,K������Kı;��&�X�E�%5Q?w��6��bX�'響\Mı,K��vtɬ�d���ɚ��r%�bX���Yq,K����ӑ,K�����n%�`~?%�O����iȖ%�bv~�?t�J�j�K;����oq�ߟ����"X�%����7����%�bX����M�"X�%���u�7ı,O�W���d�h���je�%h��J�ʵ����W���e�ޤ��M�l7H<���88�DL�^�Sn�/Nk�-��:��g�L/<�	S\l�sAXX�E��y����܎�n���rcHk�t�Xs����0�jL�3�����#����n��5�m�Mϣ��n'qpX�F3�q�g�}����H���0g���N�[0j�
��n*͕� ��ߝ��w���}���!9y��WZkpr�jp��.��K�!s�!m�kD>��4����}�%�fL�\�'�,K��g�&�X�%��=�fӑ,K��w�� NDȖ%�����ӑ,Kħ�_�C��)�v�}�oq�������}����ʱș��>�Yq,K�����iȖ%�bvg{q7�Dʙ��߾������n]K3Z�ND�,K���dMı,K�{�ND��A!�2'�;���Kı>���m9ı,N�vee�ɫc����D�K���D��~�߽6��bX�']~�7ı,N���6��bX�L��w�dMı,K����MJk�5�֍�"X�%��n�*n%�bX|�~�y��yı,N�~�D�Kı;�{�iȖ%�bxOn6:';�s�	T�]ٻVW������=Oa+�6|ձ퐞?}��{�������[��S�,K�����iȖ%�b{��Yq,K�����<��,K߮��7ı,K���|�Z�Mm2�SiȖ%�b{��Yp�h�(sP
%�����CI�2!�6i! �@3 4����|Q,Ns�8m9ı,O�w뉸�%�bw�wٴ�{���r{��7���O�V�k�O����bX�'���ND�,K�;ۉ��?���Q5�~���Kı?g��ț�bX�%{�����u��
ff��"X�|�����\Mı,K�~��iȖ%�bw;�dMı,�	�>�~��r%�bX���~5���e�&RkZ���bX�'|��6��bX���_���YȖ%�b~���6��bX�'fw�q,K�罷�� 8r݉��P��z���N�5fn��K��v�:2>��{���B���l֧Ȗ%�`~T�����'"X�%����ӑ,K�����~r&D�,O=�M�"X�%��g�+-�MXk��f�&�X�%����Ӑ�?�����'響\Mı,K�����Kı;��&�|�L�bx{��95.��0��Ѵ�Kı>�߮&�X�%��;�ͧ"X�^��!�0@
U��Dly�#�|,MD�������%�b~���6���oq����?$���Fw��bY����s��Kı>������%�by���K��BdO�����Kı/�ӳ�&�Y��2�L֦ӑ,K��{�dMı,K�c���i�Kı>�߮&�X�%��;�ͧ"X�%�{��R�WY��[`�v�m�z�Ӷ�:�6�T�Y��ݗ=����ϰ������g�_���f����X�%����ӑ,K���{q7ı,Ny��l>Fy"X�'�ߵ�7ı,J������u��,̹�iȖ%�bvg�����ʀ�Q5�����m9ı,O���dMı,K�=��"|��TȖ%=�ߍfe�3YnI���\Mı,K�~��iȖ%�bw=�&�X�A?-5Q;߿p�r%�bX��}��n%�bX�y=���.][s4ankSiȖ%�)"}������%�b{�~��Kı;3��Mı,�S��O�Hi�t�����ȁ���?M�"X�%����2���Ն����k"n%�bX�y�xm9ı,?*���鿿\O"X�%��o��r%�bX��{����!������y�L&�.bڕ���v��x�b��ԜP��&�.�\^ �[����ڗSf3Z8�D�,K���n%�bX����r%�bX��{���	9"X�'���ND�,K�/K���e��Yu�.j�n%�bX����r"�r&D�>������%�b{�~��Kı;3��M��2�D�/�ӳ�&�Y��2�L֦ӑ,K��;��&�X�%����ӑ,~XdL��Ͼ���bX�'��������7���{�7����h�{T�Yɸ�%�����5����ӑ,K��3�뉸�%�bs��iȖ%��?
-�O���Yq,Kį�ߏ��[��0�fe�ND�,K�;ۉ��%�a��
����6�ı,K�~�����%�by���Kı"t���D �.�u�݉H�4dԗAqѤ�
o8�y�S��Xp��x��tMi�c0<ݜ����|��O$���]D�4�.��A�� a�pC���<�1a__�9$�lS�	c��6�=��� �K\w�Ca�!�o2�pv����?[(�������/cm�Y"��~��UKQ]�)��b�6w7:��U���e�E+�J��Z�D�e�4�N�83��b�vˬc�0��9��]#�Ń��
�0敪�����j�ō��
70����3���]����j�������ݢ�	gVq�;i��ȐF�-h8ٶq��(,�a�ngVVg���N�	هur���y\0�J�7Rsk����q��ͻK�ڻn(8�h
�jӝ�S���Yr<����J�r�����9`�3vy톪�X$�c;mQԫ])6�\�҅-R�3�ӜZ�a�g��q���(yՏ]�,;� �l��`�3��6S�:踉��#����O�+��ƇI׌�cz�����M�R�ʦ�6�q�m&�Z�Hu�:�AvB��sr�ی��U�Y� �GR���^gn�0�q�Y�s<ZH��WGjɺ�� �Y`Z���D��+hI`�ej*�8�Ӗ��U@�"R�SZ�ۍp�W8��]���t��$[2��x���XW#�u̲TJ�:mp6+���m�9Χ�v�ŮQ�S���*�V,=5�k-8+<��5c���"Z���!OY8]����^t��4cs���Ͷ��,�:�͍,�M=���wF\Fܫp�UOk���y�!�`~���hy��3�a汃{fu����S��������{Kd)r�E�N��M,ntSk,$�i�$D���d�Xr��]��`���*��^3�s��ظҳ���9v���X[j��r�g6�h��ٍq�mi94(0��V���v���.z���j������q��#,�n����uy7/b�5]N��V6��3n����q�&x���M��ͺocoG�Qp�z�"ٝ�4�c��%�v���&�����9*��Iu��p��1b#D��	�������ۍY�1� ���ӍpC����;T�[erMq�]��'&&;m��U��"�^p��O�^*G��;Q�&�O(�>U������Eꇩ�T�Qj�	� z����CJ����jB�w3.��MY��#lg�(ĥ<���n��T�O���Iv�N�&�y��*�f�Z�{3�wk�v1v�׎�R�j�և�����%��6
 -烂�a��j[���[:+���l;r;˹�W"vd�^ׇt�$��:��0G���3�5���N獞9�p��<��nt�t�.��gP�<P���v�JF"=.�]HX�:��cVy���ULC�e��3��4M2Mfjk5��n�nv�t��J�؀���x���L�<&�;����0]��l��w�{��7��������ND�,K���"n%�bX�y�xl>T�DȖ%��Ͼ���bX�'���g5s˩�.�-�jm9ı,�{t���D��uQ,N���6��bX�'響\Mı,K�w}�ND�L��,O�>�Yn�j�X�L�j�7ı,O}��6��bX�'fw�q,�Jj&�{���6��bX�����7ı,Ny��0�Ժ�h�0��Ѵ�Kϐ��>��뉸�%�by���m9ı,�{t��bX�!n���_�RB����멺�.���4e֮&�X�%��;�ͧ"X�%���n�q,K���{۴�Kı;3��Mı,K��;s0�Ʉũw7S!�v�-�N�ܻk��KKb�\�q���%�9ίپ9��S��;5������oq���I��%�by���r%�bX���n�g"dK��߷��r%�w������|�%��9����7�ı<�^��9 �h4 ��.�Ot��"��iD�M��@xȖ%�ٛ��n%�bX����m9ı,罺Mı,K���v�d��f,��j�9ı,N���q,K���fӑ,K��{ۤ�Kı<�^��9ı,Jy�zj�[�j۩2�Y����%��D�߹��r%�bX?g~�Mı,K�5�nӑ,K���'鿿\Mı,K�~��sY�e��f�K5�M�"X�%����I��%�a�G�w߮�Ȗ%�b}3�\Mı,K�w}�ND�,��n��~~=a�sF+��]=�#r��a�uP�j��Ճ+��y�1��;���:��9�3Z�ND�,K�u߮ӑ,K�����n%�bX����~@��ؚ�bX?����Kı=���9f�Ʉ˚�ND�,K�;ۉ�|1ș��߷��r%�bX?g�]&�X�%����iȟ"�L�buߎ?d��N������oq���~��iȖ%�`�;ۤ�K���)�L]* �*����;�s��Kı>���q,K�纳ٝ5�kZ�E��35��K�����?����n%�bX���v��bX�'fw�q,K!�Ȟ{��M�&���~~���z(�T]�۽�{����&��/TP#ٝ���%�bX�{���r%�bX=���7ı,O{�c��sY4�Yf�q����c�ZYk�:��Eg��#���w}��ﰩ'f,��j�<�bX�'�>��n%�bX���ӑ,K��w�A�9"X�'��]�"X�%�O~��W2�3V�I���\Mı,K�w��r(G"dK���I��%�b{���r%�bX���n&�|�TȖ'�v��sY�2�[4R�f���bX��߮�q,K���{۴�K��DȟL��q,K��߾�ӑ,K��gfV[����9�3Z�Mı,�������>�v��bX�'�~���bX�'<�y��K���"��T�.D
$L(�H Ҩ-@�ZJj�:��������ˤ�Kı>���9	�F��a�5��r%�bX���n&�X�%���׿s��i�Kİg߮�q,K��{��ӑ,K���]d�5��a�v���6�s�����v4���^ˠ�e,��F�~��}$��p܌>���X�%��u߮ӑ,K��{�dMı,K��{�ND�,K�;ۉ����ow��7�9�S\��>�7��bX���Yp���&�X��߿fӑ,K��3�뉸�%�by���������;�ow����q]2�E�bn%�bX�g~�6��bX�'fw�q,K���wٴ�Kı;��&�X�%�^�};.f]e3�]\�m9ĳ���>��뉸�%�b{����Kı;��&�X��2'���fӑ,Kħ�[�n�n��MkWq,K���wٴ�Kİ� G�}��'"X�%��w�iȖ%�bvg{q7ı,C"(AJT�Q*@)�N�d��w�Cq֜�8
�q��Cڴ+7c����ه\��#��{5����ֳl����rc]nj���U]��gD��,cnv���^����+��Zm�XrU�B�N���	�g��۞Y�$�	���1quͫ8����=jru�Z��(ܻ9xl����6��1�����_�����E��nmY1�=���넻g��Rd�_ CC�f���亚��K��l�m�7Z�sfx��WL�ζ� d���������7ҽ���8*��w�{�K����k"n%�bX��{��r%�bX�����+��"n%�bw��m9ı,O��L��y�i�s35�ț�bX�'3��6���X�L�b}3�&�X�%��{��ӑ,K��7tB��T¢�����K��.�A�LֳiȖ%�b}3�&�X�%���iȖ?2&D�>�Yq,K��;�ٴ�Kı=��K�e�[5��K�2�Wq,K>X���M�"X�%�~��j&�X�%����ͧ"X��2'�_}q7ı,O���d֮�٣2�f�6��bX�%�{�D�Kİ��� ������{ı,O�?~���bX�'���ͧ"X�%�����ۯXn�X�B��f��v.�*4�7X�fWs]Y��<��zK;��������M]j���D�Kı<���m9ı,N��n&�X�%���a� �"dK��>�Yq,KĽ���&�˗V���u���r%�bX�v벦��EH@v  lP��/"X��w��r%�bX��}�D�Kı9�����O���CX���{��v��\�[!�w��oq���o��r%�bX���D�K�R"y����r%�bX������Kı=��ܳ���Lնh��֦ӑ,K>���ț�bX�'�߾ͧ"X�%�ܽ�bn%�`|�̉�{Ϧӑ,K���S+-�Դ�9���dMı,K��{�ND�,K�{���Kı<���m9ı,N�{����%�bq�]�K.gr3���ؙ]Qѹڃs�V��3�34ٹ�ȗ'nˣ_f��7	�Z&I�e֯Ȗ%�b}��q,K���wٴ�Kı;��Ȅ�L�bX�w_}~�7���{���w�� 4ӊ٧q,K���{۴�??�J�&�X����dMı,Kߵ���r%�bRۧ3\���D)!u3��.��dљi5�]�"X�%��w�dMı,K�뽻ND�Ñ��!B(A����Sj�\,L��u�Z��bX�'~�~�ND�,K���k�Y����}�����ݻ����}��iȖ%�b}�g֦�X�%����iȖ%��_ȷQ?o��ț�bX�%�v~�f��e�S0�m�j�9ı,N����%�a�	{��v�D�,K���ț�bX�'=�{v��bX�'��}�Mf���33.�����z��cF�����U�*�ۀF����O;
.��q0{���oq����/�۴�Kı;��Yq,K���n���"dK���_J��bX�'}��/5s$3Vܺ0�Z��r%�bX��{���|�"dK���ӑ,K���_J��bX�'���ݧ"~Q���K�����nl��9���dMı,Kߵ���r%�bX��벦�X�C"dO{��v��bX����腄)!I
H[�u4�~E�(�d�k6��bY����n��7ı,O{��v��bX�'s��"n%�`UC�	�T�. GH��j'���fӑ,K��N�]][f�Z�u�s5*n%�bX�{�{v��bX�'s��"n%�bX��{��r%�bX��벦�X�%��P��}�f[I�˖�J,�j4��7������.��J���佴$d�=�{��|�0�r�j��bX�%��>�����%�bs=�siȖ%�bwۮ�+9"X�'��~�ND�,K�ߦ��h��f��֫��dMı,K��{�NC�9"X�v��Sq,K�����iȖ%�bw=�&�~_�&�5ĿN�߮�)'/K?{���oq���ߥ�a7ı,O=׽�ND���Dȟg~�D�Kı<���m9ı,Jy'�\��5�n��[�J��bY�!*!k�Ӑ���$�>��?N�X�e4����6�I���-�[XDDB�>��7|`��8B�W_���?�q�J^��� ;����L�,��;8���;��]F0�ێ#,�qe�Sյ@��Lf�[��q�dt�s�wuu�<�#��?��s��v�l�-Ù�>��u-�m����iʯU�vf��1�Ub,��Q)���J3k��]�d��6��kcZn-qj�q�.1���`�z����M�'WE��⨽�ɷY����z�1����k2f�f�շ5A��sS���/4P����˳l��sͻ7E=���#V;p����\����'�G��>Q��m�k� {���Z���@����Oi�$���9�{�M�ffbG]>�∄������=/���dd���H�F)"rC@�w�@/-�~���.+�=��]+VG$1��Ł�3��x��V �m�B���S����?���Ds	�"�d�@�v׀t.o8��}8�`B��]O�Bp��]MG8�;3����v��B*�pv�i�}���1;	mbRN^2C?�9�� �ֹ�����!�}ՀB�[^�$��JC@�_j����� $`F0		 �Q�ć�xW�Hg�H��L0 �*K!C�L�Æ4Wjh�? �G������&�yw��@���1"ڼ���c�!�j��� ��� �:�a�%�P�����h�e_���J�N)��^��m���x�B���0��iR�]���wXݶ`�DN���w�Ɓ��@�p���b�pS`J��N����s�n�C�����S<e����������lj4��b�'$8}��^[f�u��(�$�����}=�����	��$q94�)�U�^�{�M z���%�
���ӒU�suWJ��bf��>�����
T�ҁ%(Q7�`@#�J�)
$�R+ ��D�/��9����Ħ��D�D��pm1Ӷ��A���4Mh�}�<9��ÁM��
(a�]�t
H�(8b��j�C~x� �6 H��xm(��@IQX%��B�4K�v0"�*4 $E�E���$	��c�P�w��8���f����X�B$��Qӯh6�b@������dȕ�D4�pPҞ����.8�q����)�:���}@P�ĝS�P�W����E��A<�#�t/BQ�*P��!)�����0E��	��X�!��z����n��{ޚ��*�� �p�u���aR�n� m��9B���?��Շ�!b^�x�/jYM���1���F�RF��ݬ��n��#�æ���n�����w�����I	̘�$�w�ƁU��v��D|���}��}Ҿ�L�b����'��U�����m���)wQJ��������"���w�؃� � � � ߾��lA�lA��A�o�؃� � � � ���߮�A���7{���wx��~q�$��v*�<���!`�{����<����}���y>��]�<����+)"EFX��
>���y�������e�A�����n�w�������6 �666(��k��A���ϻ���A������6 �666?�Ϻ|��Z�\�%�.	���=�-1������ ��ڱr�gi,�����{���D���o������s`�`�`���~�v �666>}��6 �666=�~� �lll{�w�؃� � � � ߡ�oή����̳,�j�A�lll|���lA�lll{���b �`�`�`��{���A���ϵ��b"�`�`�`�Od�;�~��k.I���Sb �`�`�`����y���6 �6*���k��A���ϻ���A������ܷ���l��D�f��<���� 9��?M�<��������؃� � � � ��w�؃� � � � �����A�����>��3����B�jlA�lll|�_}v �666(~F����� �`�`�`���~��A�A�A�A���b �`�`�`��� !����'��Ifk2�3&�k5���CC;���涵����ݭ���吠��(��j���N��57 ����.i�trk�Հՠ�9��v���mtwd2p�҆�:�����F�6�\r(�x���rʹ.x�ΐ^kT��i��PEYy:�,:Y'��oN�v0L<���[vz�I����b�>ɰ�-l�c�g<P\�R����um��w����G`uT�8Z�as�e���5u5.n�5�1���1%ֱ�KcX��]�un1�-�w:ˆ�ɭ$�2�Wb �`�`�`�����lA�lll{���b �`�`�`��{���A���ϵ��b �`�`�`��'�/�˩&��3Z��M�<����{߸lA�Dlll{�w�؃� � � � �����A�lll|���lA�Tlllo��C�˩r噭k5ff��<����}���y>��]�<��?�Tb!�A� �����y����<��������L֦��Z�Y�R�jlA�lll|�_}v �666>}��6 �666=�~��A�A�U�A���b �`�`�`��v���Y��u5�5f�Wb �`�`�`�����b �`�`�`�w����A�����M�<�����k�-���>A�_�f50����(�2'w'kW�ɫH8z��f��������v��(LQ�)����즁�v�~������4j�M-�8��0���'�{����/D	lP���K�(�?=ެ���X��2����R�N˽�@��SOf~P���}� z���)R�]�IJ���ˡ%�s�,7ذ�ڰ���~���Z��=qz5 �Li��7 ;��;$�t� ?�]>ߢ��#��ܷM��q�~ۗ��d�ݸ�tY랼`�[�s�s��{����}��,"f�䪵�w/�`����r�I~��}��__=�s"�G���8h�ՠ{�ـ=׋ ���:IL�+��\���՗r�Sus�n��=׋P�@��+F��j%�F��c����O�K�}�rnI�s�]���q�ڮ(��R�n��;f�w]`tB���� �s�53�J��&�Z.���;fСz����_�׋ ���(B��'(=f�r�6k��ӌ�����Ξ۪�y��#sv���Y�]	<�������=-��=�l�?n�_��@���?�6<y��x�#�9�)����}� �����!�o� r�jz�l.n�E"IŠ}������b\V������w��[PM49#�nf��[��v�t�t��o�(<�!R���,�v��s#�G�ȱ)�ڴ~[��?�����^��1�4\U�YħSe����Ue�ք-,�3��K8�.a��H��}�}�dmGk���m��O�{���$�~���ՀzV�EUuU]�ML�w8�׋:_DEQ���`=�V�M�|��J���jg��2'2a�����?���נr�V��z�`��T�g,����M\՘%�U���`����?n�XB_B���|`��Oi�&@i�$�@�v���Q����}|`�u�J��)�6�aD'�D�4RD6�=���?6�..-�7)u�;i��eЃ���Lʴ��3y7m]H���Y�OYĉ/��D�s�c1eM��^p)A�:;E^�^L�&:`^�Q;M�-��#CUcS0F���ld\8ݫm��v���\pZ��ɸ�^|N�nծ���l={nK�8,�;!z���]����kd�f�=�YC��Q3��W'��y��렁������{�{����G��r�A�\d�Oư�C���i5-��8ۅ.���b���%�U��a�ݷ����s`���1�$� ��W0�6�rG�������1#��=�~��>�n����=��Ndq��I% ��� :d���qR��@���q�	r=~���{�@����f�DGТm�}X�gHUW�Y��xu{�h7 #�����j��x���4�`ڑ�RD��m[���+�6A��O<<�'`A���C���w����js�����@�w�������	z�{�ŀ|���J&r˚����\�ܓ��{��i_AО���O' ��ŀn�fr���t}4�`�-XTҢ�� ޮ��?n�X|���[��@��@�9�R(D�y"�C������� �;��>��!*g�-ȫ?���&�NH�������G����oWt��^, Q
�w'@ݯ8�+KCtnl.cp��RP��՛-v��OI#���w���~Ḧ^*x-<\���$����͂ �˿��Ɯ$XLQ��Wj�g�ߒ9o�4}<h.������ŝ*ߓr742]��o�`�هЗ�^�"&	(G�t;�&��o7${]Ӏn뙩�&h�T�Z�]U���(J����l�}X�78O��� {�<k�8�18�4�{^����;��/����;�)�}����&��c�C�؝*7�w=A�!f`vX��Q�g�"\P�;Y=�3$�Zx�L2x%"����@���h���U�zmK�(D��EQrM\���3�%�QTw}�,�{���տ߳�EGVQy�M�����0��`��Xr_(�T����{���/;S�Nb���9$�h{3?b�ٹ'�g�]�9�uٹ �ڋ�QaP�XAV$V$��2�PI8K�D/��� M�Û�����Qj��� �� �G�"7����;���˽�@����7 �'2�h2]m�ڎ�[r�S���n!���]dȱ26�4���v�h��8�����~�W��__$��&AbNc�9u�3��&�}X�wV�]�>JbE���D���p�:���9-���Jϟ_}|`{.��,E�ER������Հy��n�����٘����j^�B%$�6D�n <�� �� :ۘ��b�DĒ@��z��t��b����0��h#�q2t��`��"> b"1#�Ќ& })#�(FD���Q�� O$ R�Ϊm��HBm�A������|�	�R$Č���$#+��(C�8F�l"�g�\P#f�e���"��j��]$�=hP*`�b;�5�j�_(FR1�!!i�
al�1d@�!�8�����;�jR]�ŶCm��t�v��q��45N�ũ�7a�����];��^q�۱�37���I��D��R;�b�+���gM��YE�s�Rr�K��\�#���c�R�������A�!��ײ\K�6{]nՌ�j�nXTn6�j�͕�E��4A�s\��v�R=tT�v��.��r鉒�W�*��q��g� ��5e�3���<�\��N�u�U��l��lp��nvo^�JL��5�!�A�5��`s)�n[h6,`6 �D�̵T���]����;I6�TKC�L��6������q�<���t�H�N�m���pؗx�Uݙ�I��R�s�;2��ڻv�e*U�dZ�:�;OOCjUÝ@�V���n:�bҦ|��Hy,[�q�����:��j�!*u
�2�4�$����C�L��r���D�n��h��һ�y���K�.��V�-U;��'@R�t��J7Ztݛkf���VU����5N�cX�&c��G*^���`�Up��[�5�me`'d0��n�r2i+j�9[Dd��K��zM�9��o.]muj�h�s�o�Y�\���3�s�[V�[�%�Z瓊�������pi�օ�Vn���8�k �]<,�]X7;�,�+�X�%�m���*��rJ�'1�ln��m��y��{j_v^�΄^ÉNn
6_mj%t��9��u�p��	2�;GS���Z��i�$(mI��㎽J֪���pu�	�\Xm(�0b�:�i��D�X8Aeȫ���fQ]�M˷�{2���-u	5��ʹ���+O�	��tX��[�(�Pq1�����"�/d�tԘ����C�nWZJ�z6ɵ�I�;X.�[����c	����n����l�)bkT��o9eYiD��[W���)�uv�ݧA��i@�%��ʩ�.l�0I�u�*]m����a��*����KT5��k5�I�)u�B�Dh�G�����T�x�V�S�<"��z�D�������h�����x��Qv)������{���!
5�V�����lť�qb��;u�՛�����n�m�{Ocb����K�\��z�@�;]@�6+�8��{0�R�WN�t��͊�g3�R���*�82�\�fv,q�Qu�=�㎷k���]:1��T.���n��9���H�n������/M�KX(�n'�Onˣz5Z�3�
�&�����N��6Q�F1v�w��������w������ٴ�n�fl�"m��f������t.+��97��{��o��;���$dr���נur������߳3�;���h����'28�qȒ�N��u�l���?k�`u�s�J">����z�~�R8ӄ�	�9������6��:ۘ��K2����`ҊG���\��|��ס�߱W�y���4�I�X����C@�Z��O��%�߱�6�0���`8s[���8���dv�.,�̼�	n�wN�8̏u���瓀���n-5s�����7X�vϡ(K��>Z}|�ǚcA2`���\��}���*qI���;����}������נ�U"NI�dI8����k�9(S;-�`w����:V�D�I�����V���נurס�ߗ/�Ɓ��k �ȣȋ%$Z{^������?����r��m����~w|0���U��ynNB�+���L�U����q��i�<��8G�L��E����gɺ�?k�`u�~����Q�{�� \}!�Q?U�T�R��Wu�~�lϡ(��7���-�`���?��bG�|�KD�s�h��7$���spN�@*11`��=ʴ���-�Ė���(7P�i��ή��?:np>��;�8�>��KR�H.�mjs�}���y��l��7Dԁ6;�ig�ع���\n����Cu�vܺ����o��vx�N=�<b��Uv]J�6߿����ݲ�k�|�����:�,��YmH�r-��M�ڴu��@�v��3?~H�����EsI9�wN�d��EW}_}8�� �/(���	�-���e���-�y�uٹ9��"z�l �E��M��z�/��۹$;>A[����pZk�h��;]�@�_r� ��� ��ib��͇�e�����[C�u�Ms-Z��ۧAfxv�s3c�4�K���'"�_Ok�h��U�v�V��k��k��ئʫ0t���!/�EP��}8y(IL���Ӏy��7�j�,HZ�U ���6|������D��0-�`��cP�I&�%�=�\~�����gu��D��u`M�Ϊ�sUJj�W8���"!F��W����ܓ�3���h
>�#�}�����2�\N��ӲNA���y"^��v�M��jb���b�jj�ˉb)x{A���z�WX6R5=�����Z�e�b��;�:���O -�s�E{iy]�#��ٛVRzn���^�\j�b����f���:$��\��VL�&T��q�ljض�ͫ�:E�	æL�M]��u��U�g���Oe,����)��!s2\��$���jMkR��sr��Qxp�ڛi�G�S]^��B˱5v���;Kfv�6cE-ΰ�2����`r�� ����z���_B����`w�{?�$�8H��9�����q�8��`�7Y�(�(���U?X�`�(�O@��-��i��K��@:�ҽ��DLBM~I����h�v�~���hvIhs�]���$�87���@������s��Z�S@��?<N	4d$��cX��ՎäZz�5!�ln�{q��ո���iN:ܛZ�U ���5ֲpަ� ��}�_= ���/��"RI�dm�-�3���Sŀh�6�9'u�vn�u� ����$�K꣤�\}U*榒r(Š{�;^�z��h�h�k�d�m��nCC�3?~��v����k� ����?7l���LNHӄq��n=�}ʴqڴ��`�7XD(�ӸʅWeЀ��um���㫳��;-��z�vtv�kVx�i�cI�&Ɯm0x�X�����@�,����^��̵�ܭ1h!�	]�
���v��ID%2l�u`:��@��}���j��$��L��6I���rO/�{����J� 	$��Ƞ�J9��}�ܓ�}�����<�	��#�@��Z�z���v���v���_L�̫�d��6�G�s�ՠs�S@��@��Z���u�D�P��jcn��7}�l������sk=Z60m-ٹ�9Ս��)�4�rF��留�����k�9�j�;�׬�72(ۍ������1J���ۭ����-�6�_r�i����q�\�^��;V��YM��� Ϻ���i9`�9u�����`���1U�z����"B�� �
io�����;�J��'%#�n-��������:����9�j�8������8���rж3�9ϘBn��Z��i��uv"��崢P0i�i�C�8h\��\�^��;V��YM���<�	��77}Rb�$�t� �- r�X�H)$�㍬��Wj�9�)�w��h\�^��qe+j	����"���w{8��Ӏz|��I~��==�^��Q�Ndq�M9�r�}Rb�$�t� ;�uT�U0D�`T���d�H���63�ɨvP��u[���*]��t�"pLW8/O7'[q�k��une�����]���.���N���v�Qx�S����x%x����`l�`m6�A��	�6�ӎ�����nɃT�=�L��ӤeD;y'��#��H�^Ln��g���|�4���sI֍&k����C�۝�:!Ӵ틥�;k������8*��եyg��֬��̉V;��ۖQKeVL��g��\��˛�:�2,	�5m�ʓ�%�;����b ��d�Ɠ���z8�[�٘���x�:��=��k�-�Zb�C���<�@wM����_T����-�ޔ0�ƙ$1�#����^��̵��h��9mM��1�&L�w�h��1�Z�l㖀��3�.���4��b��@�]Om���J����v��[��6�ò&���Wg�˭�@zd���x�:���Ŕ��&�NE0n-����^��HF+'X�i v��_K�{�����k�>�ՠw��FA9���yyy� �-��& =2K@wM� ϻ�X��MĚȓ�-��k�>�ՠs�S@�_j�/R�6�NF�4����v�߿fw��k�Z2נ{��\=W�yB<�ژ��8-J�=$'&�#�Wh���˓���p�{:���DZpBR<���O�@�_j�8������y��@��a�2HcXJ� ݭs�%2l���]���!��Ɓ�?yǏ!�a2`�JE�qs-z����qt oD%�[,���0�0! �"H��D0��H���a�Pr�M`26�x8�&��p@
������,B%p�A 鯞�bi���Ɣ�;WjD$HR$7���j$R� og�`�4����$��;����`�`C�P����bPvI�)�����;�4���9) B�L�Ƴ
B$5[eҡȜ�D��HY-&���6�),���0h1,���6Gڂ>+�aP��A��@:�t4�]�}x'� ��F���P�0�C�� �qH�DA�v��k� �r;�Wd�ݢ�]T����!O��� ��v�� �k�8�,*��$��l�@���D7o��:�� ���?6\���M���45�ӱ�k�'b%�f��4Y���\4��Pw-m�+�VPZ�m��Z� s��`�7<�G�n���ёƛ�5�'$Z\�^��v����z�V���H��<��m9x4����?yh���;�ڴ
�����V����"��Cٟ�z��ܓ���w$���srp�DR��1@���g��@��W�Z����N4�!�A8h�9h	}Rb�$�o`�vKyw3q��K��iV��v�M��:�[�%=��n0�k�"\P��]~����3�[���aB��~�_�b�$�o`�o�$E�d��L8����v���ߒ=l� n�N �ɺϒ��CvQ��Sd̍Ȝ�h�x�;�ڴ��K˹�=�~��;���c�m��nC@�^�����Λ��_(U���� ���i��YrE�U�W�}]�@om��k�!Z��
$%�+�������	�S���x��ͪ��q�i��q���N�^Nݒ�6:�d���xu�b�Mq=��܁[gm��FDn�v�^�	����x��\K=t$�3̺�����.Ǹ	�Ma=���RI׮��Rr�:�/+�NJ��d�Ό�e�5���ڜ�qrM�䋒��;wD��T���
��D7D�z�ͫ&�N-���u&j椰5�2���T����k�6�99ne�盬��\���ζz�Y,��:�ۀF՟τ��wo�*�J�F�.� �wN ��0��?$�/�;Ǟ�m�4�ji��A�N-��h��p>c���9BK�IU=��a�2HcPN����
�J���31���s�0N��Պ�L�Z&�f�p9/�$��V�W�N ��4��� ��ĲAI&$m�=�� ��Q	}�~����N ��u�����~���iice�tM�.N�56�i��:X�B�&9t�d����%,Z*ɻ���f�Z� s�:�"�!�?yh��j1�L�$��nC@�_jߠ��A!آs5L��@���#2r���ܓ߳�]�[�M ϻ�X��MĚȓ�-�1���s�%
&{��7O� �Ir��NF�6G����~����-޷��Z��I)��:���$ɪ���A8�{)�fe��|�|y�Wj�9n$�n�,Lr`�As1U����FK�:�f�z�ە.3"n�s��&(�i��j	�@�_j�*�+�>���(�!��_L�X*�3qh�U3wh	}	�L��=��r�类���/F�AI&D��y��@���Z�"!	""�(�7k\�wGX�9UmA6�Ԏ`�Z���޻�@��-�R���Z3���ds"�84���;�ڴ��>���y��@���;�˙���X�71��d�8�1�b�م�ONc�qj�]���;��i�?�r�7��7k"NH�˾<���h�S@�_j����Sm'#Ll� ���Q2w;� n�N ��u�n�+M,ԛ�,Pd�@���z�V�ļ���@矼��zPdjH����Dx�%�& =2KA着U��0Y�?E0��<��(p�y��nI�~���2���.��"�*�+�?�����z�z�W�o�����~���.^���X��ew���$���s�W�e��HL�׶C�c�p�ٮh�.��_}8{l�7k\�?Ht���w�ͨ&ؚ���@����k�Ϙ� ������v5�\�S���M�y��h\��ޭ�������iȆ�$�@���@��V�oe4<���@3�^G�lNH�������h�S@�_j�N�;;��+�!A��{7L��d����YM��	Δ�ۡ��މg.֮�j�N��-�s�G������97SW,8資6ڷ9o]��ɇB�W���pE�r���[sQ�=���q�qθm���AO�c���f�17m.�I��at�NX^�[s�%�{q�7�zbS�:�K�m����	����vlT�Ak�n�ݝ�M7�����n��F�����ww;ݦ�㬉rn�-�qͬ�3�C.ӹmUm��2���qtg�n,���,ԛ�,P�!8����w��hr��Wj���F�5$L�5�@7�Z_Bb�$��`��3�L��
�3qh�U3w8��>���@�s@�_j�;��z�GrL��w5��(���o��Ӏo�}� ݭs�j���3�V�dM�Dr`�Z��X�k�e����s�|�"���]��t�l���+=�^�.�U�v�8��-ٹ�������_�WL���p
�����i^���@�s@3�匎4�I�#�G�uZW���~�D�R"���.�y�}�܇�����נx��7�8�`��� ��np6�a�IL�����Z��4�RL��	�C�1w��٠l���6[`j����m����J�uwSe����Z�=>�X�Du���xu�Ӏy�� �BP���"��J�j���&t����/9y\���j�R���\N�q����,���%?L��?���<��$�I :��@6��˭ͼ�ݡȘ�����${�x�:�|�
�J��ֱAH�!�0n-��l����� �^yTL]43�X�cD[*.��0�R=�-?(O��>z|���/s�p���N'Uk�J"'k_VӼu`�M� �{��uw)R$��dR9�Wi^���!kϾ���}� ��]`��p�u��Sh��-�,綮��эyY����c��Ob�Z����h^Fa�3.��?z����`�k�P�Ht�:���4�RX�X�"Bqh۹�߿g�H����<��=�;V� ���dr5�P�f����U�W��~K�~��=�ذk�N1*f��6wX�c�����5�Ł�$�ڨJ(Q$�� � �"0]C�'s�|�_b��rL#N�qڴT���1 �1 G�9��w�n:���ٯ��q��y�0�ݦR�prZ�E�1�c�V�ݟ7X�H�()F4���/��4O����:�G�mwN�>�&j�Z�84�s4��g��?���<���Zm���� �Us�qH���H�z��V�����Q
e�v,g_V g8��[Ĝq0hq�=�;V��^,��u��DK��V��j��&eU��"Bqh۹�qs��v��y��ܓGsPvT��6�]�B	x�$i�-�����F��$4�b��0��� �xW�:5�a���`$`_S��Ri�}Kd�|4��}(C�
�'`��!��|c��������=����P|3�1	A�Bl�X��O4]�b������@�iCh��
���<"B%x�{��� �y����P�k��C��6�#�yxav���F�����&�Z	]!��0X�`���n�����w��]WT�4ԫW3�(MW�`Mpjiӹ�	ͅ.̵�t���:���@)]v��OCdu����ie�I�;���2��� �j�X��g���s n����Q�b��2�}�r#�jv�����J�S��:1�sڅ���L��][	vٺ�эF�22d��	]�:M8$�Ojb�+������`I����
;��W�N�F�-��z�:f۵�ح˞}1����JMl9��cu�`N�^uԷR��)�g�ܻ5���UP
��w��;R�q3�
�ڦ��))�r��Sj`��G];��.٥yl��;--������K��tL6ì�2�W'���K5qn��ƌ���Ƣ˔����'�v�m�E��+nݔ�Zd�c5�¶/����e�{f��r��.jz�Lu�J���S�͝���7,�狷]�u"���M��UUI�  �̬*ԙ�ι�WDL����m�����h<i=��cm'Q�᪀�C�3�9X�-6ƻU(`6m�iփ�79��y�:n.zSB�$β�md9a.�y�Z�h������rt,Dl�J�<ݩ��e�μ��t&�X����E
�ݻu1ed�{7�����Ղm�&q��mV:�bZ]8���"0�uk��ûj�zNA�d��˼�/i���!F����]�HP�
ŭȑu�t�Ў�R�3�h��U���,N.�vM��*۠:����B�\c������C*f���Ơ��Q�Z��g+fќ��mL4v��� e(mJ�V�e�"�3b�lI�+�fw��瓳�D���ɌSeic�꫏cb5;�6��܎��B�;�;��<[=��鴼��Y��y��rl=/N��a���m˹�kT��k9��Q�	�\!�l!�[�]\�[�q]�5b���4���`1�vI�-<�GEm�;r�;r9�q2���^4+@Q&v�mlg[v��{��h�t�<������(��b����E*�04� x��N���߅�v��]�fDNT��`g6-ۛ]CW�s&݂Z��C�2�ms�u��yem�f�i�6��G��f�8ۂ5��V�c�V[^	��X=��]�n��T�ƨ�8��B�,	���Wb�z�r��QP�%"5�[e$�ː�ט�]Xw5`ɹ��v%�y�=q���-{�2͜�M���N���jG��$�Ѫ��nmv����N�m�9�t���t>9�c�s�pխsOV�Ű-�S��BA#��G�s4��z�c�����DG��}�ذ�L�� �%?L	#�/iw4��Z���;^�=�#ڔm�0r&�&h���@H�_9�	Њ�8u�D�d��n-������@�cŁP��DW��V�����7u56T����l�]`DBJqߗ�=<��[)�{?f{,K�#�Ō��6�v����q���d��l�tg���CW\���������nh�$II�,$�>����s@�^נy�gС~�s�� l��z�UusAJh��`���(��J ��W;^��K��[��1h�8��q���@t��sB*@z㘀:[D�F�i�!�us������� :M��wR�uw�m�wu�kcŀtD(�W>��ou�l��~�B��!�i8@pGPsءw sq"%F����h�[��6�p�&��X��nf��@岚W;_�~�����
v�6�����piǠ}� ��ȩ�b���]�\R4���4�v���sO�,��Jr����sJ�Ve�y��v�S@3�.��BD��,	$Z����J_qߖ�}Հy�fD)�o� <t=�y��q0hif���@�x��T���e�\4��̭ݸ��J�v{v���2:���x�ܓۀش�!�δm��YX�J��q��S@�_j�;iw4�mz�� dr5n��Z�9B���� ����=l���Բ��%?LiH��]��Ɉ�`��Z�d���j�273@�vנr�M�}�C窕��B'w����O'��̳UI"X�N=��h��Zm.���@�����Ӂ?28x7#t5��<`7mc).(.-����J���ng�b����'!�urנv��hW���S@3�.��BD��,$�=Z׋9)�g�V ��ϛ�艐��K�i������W�����M=��*��=�/�4mi���N4�������q��L@9N*A��y��=��B8ӊC@��@r�T��bǰ@}U�;`]Bjf��*m))mbͤ �55���hJ��m;�����pV�l��v6���Ӿ��4�]�]�Ν���F�׹�n{Fܜ]5�=ł��tAj��y�u�zmPM�;�7��8v�ݎ��:]�YВrΌk�Z�,���-�kj��ݔx����rj�aYȻ����f)[��cȑ�Noe\��L���=:0=H1)���z����w�}}n1����%�\��+r�h��:�V�We��mnD��7ke뭃1)�`�G�}�ۚ�zoe4�Z��Ԋj�&�ĲI���^�0�7X��|�S'/��/�<QǠ_Y�@��@�����������I�R4�ś��I�)�H�� {�qur$��a$q��۹�q^��5� ��u�rQ�r�
��V�n��s�꛱�C�'-��m���M�<���CD>��c���m'O�1�����k�f���~�|��wwT�����͗WU7WX��g�B�B�$ �U�� LA#��d�ړS� :㘀*IwF7r�ƜRW-znv�i�ؗW������X+���V�����5�j�q�@8�}& =m�����R`�Y$�������W-znv�h��TF<H�
8��񼘙�Ik���C��-�0��X�R�9y&v`�=�Q*���q����;_j�;s�s@꽯@�s���)jbr�� � �1 �� 8xA�H��E��G�v�n��{^�>��6�!�Q�A^1 Q0�/���:wz���u35uS�eVf��s=��sWn�{kM,�bq�#����;{)�;�b�qR�s�U՚^eC9���K�H�\��v�+e��lC7��ܺ�2>=r����O�,��m�??ߏ�� �1 �� �JEm�w�mZ��)�K�v;����ީ�H�w�%M�&
%�L�:���� �9�)�H	l��2��ݻ�.����`�w������1^��srOO}ԅ�܊6���4�ڴ����:�k�;{)�w�ܹ��M5�x�%�L���rAkN�/s4r�Ξ���9��5�s�s����E"JI�-�;w4�����h��h8ZI����nb�s�� �9���rbif��(GQǠw�S@꽯@������� �jX�W#��ڗfD%.��`ʟN����o����&��+�����V��6^��7���6^��=��QP�	.����ѭ<��ʷ0�l�Ӝ�se���묃m�ρ�WL�
�%�U�nȑ]�ٶ�j\c�N��Hڟ����1�(���Լg�J-��.���ф�9�����m	�`N���]I��@m��$�z���f�h�7Zvi}t�C�뾾�
�fZ-bHg�d�+dvb��O$�}w%��Bn���͓=E����&��3$ն�Xj�DV�����綺�/�婲fyJ��%���"��s.�����w΄0���s�)�&Z��D�ʛ��O��`��`/]/� ��-ʞ=@6�?5z��X��X�� �z�9$���2��"��"os4
�|�Vv�=���Uz���ۚp�)$R$������<$��� H� �v� ��VĜm<��@꽯 �����^����:5� ~գ�*h�7`+;��]l��Y�<^Z��e��э��,OƝbD:1�L���o����R�s0s㘀*IwYu2��ueT�Z�6^��P��(�2�BȠb�hG����>�nH绫 �7�>��7��Θ&��������~��� H� �9���,J8ێLI=~�٘����/}��������@�yKŃn#�/sq �EHq�@t��@;�=߲����i7�m�D�ȌQY���n�/j�Wt��3��;��.y�XM��tK�D���π���@�gk�:�k�;{w4,��uI�)$XH�zk;1 �9�T�w�	D�.�s/(�0�w㘀q�HT}N��
B�++�ćpx M�d!�F$��(�צ��MM����Bn	���@Bn���0���{{�1����jA���f�C�@�p�� q����6$�=�P���"wo��k++),�
B�����w�j���/��n�ёJG}#0���-��R��J�l	B���%����6�#m���!FBB1��B@�D�D�A��8M��4���K$B�ZJB��X�
i"@�|�5��7�!��4�ҧ�(z���
�Q}�E<�Si�*(A�T=��(�YIC�ȈS��� �Ѯ���2s3���P�$�z����{^���נu^נokd#��pn73@w��9�q�@8�着M��ys��å��-J����Ӎ��أR=k����7�\N�q������t�]~�� �z� ׯBK�}X-H��M�&
bH��W��/��4
�|��v���7�ܳ�/sq ㊐㘀s1 �k�舉��eW+��W6UD�Z��
���>��� �z��%��i+P���!(����`<hu��M�����.��tk��Buϫ��b�6ok�9Ι1�ن8��?I"���;j�7=ו��ۜ8�=��j��d�!���g/(�0�w㘀q�Hq�@:�נrړĳSX�j$��@��ŝ
"��V �;� �z�9%	L�{�͐�F�IƜNf�W���۝�a�2�V ��,�[S7 �.�wS� �1 ㊐㘀��H��q7�)�dp�:�k�:���6^��5��`RJ�
���H�f�`�Z�0�fM]E�*s�˴��m؝oƺ��NzӳtWX���94��r�!sG)Rs�;m;�C�3�՜k�������le*���j�:���dn3Co�}|Q��ɢ��-��UȆ��c]ł��vtrٝ�)�2�I.hyG��n��x�؃�^��3ʹ\F��GE�gMԴ�#��Zl�a��Yܮ��c���eyL�m�Ƚ;��w��콷}�`�:������>Ϸ&�p�ݦS���nZ/i�cr�f��e���W��1�(���������;)�u^נ|�8u܊90Po�nf��{Z�{�� qR�)�M�������G�v�e4��������� ��\i'O�1�hd$���Հ>}� �z� ֶـy��B�m��P�$�zon��{^��=��s���ύ3J(�7C��k[Y8�1��\k7ZuX��`2.[��y�r���M8��8������;)�l�uВQ�>ŀo	Ň
f�������m�)"")DE(Rl�u�v��hW��w�R��nI���Gf����^,:�sϫ }݋ �ykrLX6�1�(���+�{��*���;m��:�k�8�8.܎90Py��m �1 䊐㘀rEH7����ߘ.׶��"�lt=�����\a��2�W�[L��B9�]��z9'%�56�����5�� �z� ��.P�H9���ؗ�I������hW��(Jd}݋ sϫ ��,�7��jE��y�"I���{s@꽯M�y���� B�*��00	(pEdD%1=w�ӯ� n��������8��~��~�z���U���$�oo���%�e����ci)Ԓ]��g�$�o��I%���}�I
�������~�9=��̦xA닍�:온P��^���#B��gl�n"Cm����Z�I��3�I/7|ޤ��{~ϾI!^�5$�ݷ���:��䘰m�cPQ��$�;��}��h^��RIr��f��U�����iq�xW�r��s>�$���5$�ݷ�����m����$�m����%m�ІG1Hԍ��H������_{��[oٝ�3v�|����-���m�@�S
�KL]�9ۭ�m�|���m'O�i��䒭���$��߳�H��MI%�m�>�$��F~ZAC����7<{]m=��y�p֩��\�;p6�����ܨ&,��������~3�H��MI%�m�>�$�}��I%���@�6�IƜNg�$�_j��K���}�IV�[Ԓ\�o���%�e����ci)Ԓ_v߳�J��ޥ�;���H^�sRI}ދ/�dq7$�L�ɟ|�U���$�;��}�I
���/~�����ϾI*��odō7�H�q�I%�}�r�~U.}߳\���~��9m���������b���a� ~�$H��]�l\=��kV�hz�jE���Z�&knlC�-�3��t(N�-��gaѮ���B�QC�m���;t�d���z}���\�I�V�^�.y�.����[RP���A��J���S�cA����v(��7$3<%�����*���.�k�o\��Ҟ<<�V����g��5�{-r3ʬvz�sm��0�b��k<G ����v��!h�=��������峛k�D�a����L��Q²��ڍ:K�T��g�WL�Ň�V�ffI���ə��y�y{�3=T���D|�K��������nb��Y$��I%�m�>�$��kz�K���>�$��\����Ie�.%[I�����s>�$��kz�K���>�$��\Ԓ_v߳�H�R�Z&��J$���I.w����-sRI}�~ϾI.��މ%���|��q�q9�|�Ir�5$�ݷ����}��I.w�����Y�bRcK",.uL����v�+ts�K�e����Q�b�9xb2~a)� �ҎI�$��g�$�S�ORIs��g�$�\�MI%�z,�%��ܓ	2(���%��S����ϰ��~����٢K{o���$��RIrݧ�y������4�̎DӉ�I+}��I.[&����O�I.�ڞ����軍7`�C�ә��$��P^�M���~���}�@���nC��M�ڊI͂Lr�ȩ H�?}�Ww����99nt�]���Zҳ�c�Zd"�r<w]�C3�+ό�v�pJ���>�w�@��s@-�>A�� /�%F�7P�F�4w� 9����h�ՠ}Ϊh)IƤi�Z��� ��0j"��B"��U�H�PhEN<*��p�x�1jI71U$�� ��0�\�[Ł�DL�>���5"8��a&DG�ڴBQ��/�ϯ z��&�(�$������K\	ٸ�U����5��У՜<�"FG�Ƞ�x�F�mŠ^ک H�#���:�rV��� ��h�@��������H���nC���j)$�}׀7Z� z�,��� �5L��q��xA�4�������m����˵T��u{��������3�J$��@�m��>Vנ���}�@�s:�&�yP�1ɆGdNi|t���4��Du#�77-sBݻq�bGǮ`WX(�H���|��@9m�z�W�3?} �v,xM
f��.������@7�Z� =rL@y�
������7kB�u �9h�T���1 r�4ܫ+��4�̍�ۋ@�mT���1 t�P㖀렄�n�m��ә�|�k�[f��>ՠ{�{�rNM��j6�ؼ8�;��B�TR�C���8kZ��"�#�{C�M�A8��8$UK"��4tG���a� 	�#O(B�G�w�@��|t�29���O����|��'s6	Л�]l�޴�BmO< �c��.�G�|�m0B�"��� �sKf����$�0p�.��� 4��/�tuLT����cO"&mP����0���}����~��.34�� H��@�L��$�B"H�p���rMz*b��3P��g��OkH$H f���#]G_}�e�g[Np]��n�5�;	ٳ5Yi6XĝN��m7=q��v��ɭ/�!��r�l몤8X��iWsD��nkA���@�t���YBu�M����9�ۂű��([l�"���g��她�{�q[DD��c��X�P��;×T�;I�]s�{V�����{ u+F�bJ�c�����u6:�����ˮ8i���`hZ{{r�j[�vκ70��V�_�~l��5s�ʵ\y[Ag�= �,�mi.��ڕ4�eۮ��v2UUlK�'h�
��;sU]���j�2�@{(�f�+l�'�I�n�NW盵�i��v�P�6�q�sJ���1����h�k[�t�i���>�˰�d8{]���>�,��=R�殶���b�1Q'qA�p�j��]X���Q��y���N.�n�Me䕉{� 1�Z�:��.;N:w`n"0�՝�9�`s�f�x$ 6����HMeMs���_lo��	۪궵]$�eu��.���nӝ�d᪀�i�6�
S�
:�m�X�r�n�.��{ 1�kj������e�u-l��C�	����MGm�v{'���m�-�%.�\��tG���Q�֢�Wld� �aC��g[��Vd7�V���#
\P��>�bS�]�y�����	!ʓ�Eʕi�Ga��-�m��g	9Y�'�\8m�q��Lj�v�l[ )v|JN��l��מlN}�;	�w=���ڔ�K+�Ҕx�CŒ+�vRu�ظ؞�zS4��6� f��#�ye�7^����Xa۳�`7E��L���f�(ͥ��2�d6�'��g3>�}�5ƫ=�Sؼ;�&-Ռ��Y|A2u��m�\uՓ��al��̗T�O
�\<�6�\V�m��6&�W[h�A�g ܖ�kv�k�uSV��+�iSVE�a��1�!���q�]�o]5�-i�$��'kdu���r�Z����z�Z�ۥ����{��X�;�ѩtMK	�ۗ1 ���}���E|(��U?*
G'����uD�^�� 1ؐM'��6
)�<}E⨐��;����f5E�V킳+u��L-���W^�~�|r��dF�#i�K�vqn�8�Ʊ-�W�S��g͍2r�ˆ�D7��̀�ݔӻ[���q\��d�U���ȼq���R:�;��l��m;��p�&�ۘ��Y58�Z�+���v$x�Y�Jc��s4=�s�]��Q��貭� �CtK���sj�A�\�tCu� nd*����������}�;����'9��궨�v]�N@�����Ϋ���]�kf���'����R��� =�~�v9h�T�����:][�V�q��xF��8�V���M��u���}
!L���S+��U]L�w35W8�|`���
!)����7]��>�kf�8$�jF�����^�t�P���R�N�(�2?��z�l�=�w��[�nhrנs�9���hN(�nA�28�/C�+��2N�әt[����7l���[����aja'褟�g���s@��� �h�Օ�hx�F�mŠw��k��!="#�x({����@F���*P��J�G�ӝ�����=��9���M�Or���*�**j���߱ t�P���R�;څ^hH���(�z���.�ޚz�۹�|�k�U���cNF�G��r*@z�L@t�-��_'�l�K*nC��{'dZ�z�QVK�#\�լ��O��Ѓ�e\�Z�Zp��`����M�%���}8-�f�8$��iI�˖��g�RoWt���p��g(��xL��]]]]`��8�Z��'�TKQ؇�9�}���;~�^��N��aM�0�"R-�}�@nEH_I�t� 'S���,2�ks6�3m��������7�@s��h�t#�&<I'1�����7\��c�ɪ"^�-��ˌK��rua;k��"��~i��>\���ՠs��h�s�S)�̒6��n=����L���p��`��� xd��i�������9�ڴ�����^���Z��Wx�c�,m%�%�w�zw��:np7""	I�(�s�
� y�Z��i�I�ȓ��|�k�:d�����T�K�&L¯7���Z�tasu7���`"lŚ���8vo2� d�d_�k#�qǠq[^���A ܊��& <�QF��f�Ѻ����=�l�P���v,��� ��^�y�J�46L��7��s@�:�a�B����[�0JKj8䍴/�9�˶��;V���S@�;w4g:�S�#mA�(�zݒZ�� ;�T���1磌�T}�������?w�Ρ&����9���F:e!�=�]s�3�*�%�
����ʎjL[h�ɭ�ycۡ�ѱv&v���ۜnPqRt�U͛*m��}Q�\�qP�8���ѹ��^��;�;8��=j��k�����P%��&����y��X�X��.�V^�щ�fJ��N�JY��:�����_o��,�tm���WN��WHƪ���������{�����ۛ;9��C�M�1u��#۫��0qב�J�ƛs�3�v�c��� �Q������׳��9�����^���@3�J�ox�ici
C@�;ug�L���X��� ��9$��9��i�I�ȓ��q_y�qڴo`��qR�)�m���ۛ���ަ� �� �����
�S����H#���I�'���S@�;w4�mz�v����1�m0ō��_��[�ݓ�p�v�o=���2�zY�1�+vnͺ�3x�r49ȜI8�����>]��qڴ.���Ӯ�Q�ĿTլ��u�Q�(��T�N�ݯ@�;w4g:�S�#mA�(�z��X�u�(�2�v, }�x �WQ[m�#O��Ǡu[^��۹������;R�Ějci\����,��u�g�� �m� r�V���O"Hq��$�&)���B�С�u���Ͷ1���S��3,��0�f�ݤ 䚀�bܓȩ~��S#�8霨��WQu55w�l�u`䘀nEH�5�:��76���.ՓwX�n���Xz�BB"TDB�(T60�&��M��dD$�]��=/]`��]eԅM\K"q$��;�)������=�3����-x�H��1��� �PrL@;�b��@J�2��v��4���Ŋ1�x���,9z�fӱ�21��]κK�K��u*YK}���7� �m���	D~�w^ -�l�m��i��Bs4�k�g���x��zh��hv��7��kW����� 9&�:H� �I���٤N&���&'~���1+�zh�ذ��`\��D"t�9�y����rO>����V�e˚���HrL@>qR rM@~���q��g���А�λm��u�kg�24(/fv��$;u��ӫ����~��� $��EH�MW#C�dN$�z9۹����[��u[^�1#��xO�"oƚř��'�ߵ�Rܓn*@Gڷ!��RH�PRM�v�hV׀~��X	D%/�� ���UUSWu4�D�V���`�}�~ }�xI�=���8D5	J��}�y�y�ˬ�J�]@�HX<�;�X3s�W,���ݬ�`�O7/��\���g�����M���k3�^���k۱@9���v��ݣ%n3m��w�%�Wv��e�@έ�s��V������S���y��C-�=M���/��
��X��3���.�fnə9/G��a�Bgs�%l6��Ud{	e�_�͛��.x)�� ���&yu.C2\.�r���y.����\�T�˒}�K�p��g���&<M��J'�{빠���v�|��{�@�l�'I��w��� rM@y�� �I�7 )�A_����e�����HrL@}��� �h�\z�AǊ6I�n� �1�qR rM@{�T�=��F�I�8�q�s�s@�vנ}����}�@Yy���(b�&8����6���1���%�K��3nu˚VI0��!R&�Li�ә�mp��T�����@>��iY�F�nY���ܓ�{ݛ�AB@⸈: ��G����kŀ~�n��)�[��sm��i��$�h��hs�s@�vנ}��� �u+�1�l�X�Q8�s���& =�*A���I�'��"q8I�s4�mz�s��g�u[�}����]w�I�,X��*��'b��&�v��ݮp�qL�;/K�{Y��E��a?E���@����{^����r�K��Vϧ�d�����ҽ��ݤ[s� =nL@{�T�/3��&��ȜI8��۹�|����v��x�pGO=��!��d,S�L�_o@t�C����iD4��/�pZ9�t��Ł���`�S~� �A���*lb@��h��0}��ȐaH��� ��� �z;4�ht�f
�d�S�R��I���	+�N�^"�c��ݖ0��fT��#��W4RR���$Jch��H;�#X�M#�lF�� �뇰ޡ�Hb6I�}!4�ﱂ]-�}�!�0�SĂ�l� ��C���=B�\E�hb"�Q� ��
u v��E�S���W��ADp�t"@��"`�*�m� �<Dd�׋�!~���Հ7S2��.��jf��`rS�}Հ{_b�=;��:/˝��4[�na#��iD��>㊐m�@{�T���1)ϴ�n���s��\�Zd-hX�li��V�=�[xh��8�y�Ң2�g`��M�X�kŀ~�n�B���!�}� ���Lx�!6�N=�v�h.���۹�qw��w��H�M'"P�����1�qR���s��;��X�߷>����@{�T��nb�{ݛ���PH����*j����Q!+��/<��3`g�_��b��NL�I�{^��T���1�qR��]�/0�ܯ\3%-r'f�M]3]���"�c"��6y�lv�q�O	V:~�?��ϻ���� ��x��Q�6[����\uwR�W53SV�ӭ�r�	(�=��`V��s�s@��[�̊96�Nbs��m�@NqR���]�Q[m�#O�3Cٙ�����=�����^�y۹�Υr�4<q5��{y�����Ɉ	�*@u�1I:���>��e����]kV���]�>S;|&VI�]�ԩnm�7�>8���5�����Ғ���d�B�'-ݫ�.�<W&�q�nջ=����RsT1��'[ǥ�jQ�-	y���·rf�m���i���n��u��s	����K4�ݼ(���c�y�E�@��}�7h�΃�ΞŌ-@]K]X�!������	�&�m��͸w8���v����$T��]��䶗&f�5��f��60s����u�b1Z�f'��V�n�d|[fER����G2����y����{_������}V��Ј��7q���`��X��X���9%	)����z�AǊ'&(����=�s@�vנ^v�h��F�I�8�{�	�*@zܘ���[s�igJ�#YI�3@�vנ^v�h]�z�n�w9�2�Mc9�d�����$Ӑ$�9�IY��r�a�l魫>G<֖'�9��A��q�s��{^��;w4�mz�²��N6�SSrO/��7�=B+�J�J¨E��] �ȁ�No�lܓ���f�}��hw�\������҉Ǡ}� =q�@�5 �����h�p��G3@�^נs�h\�z�kŀ|��(����r+�������}xϵ����`���"#�_�n���L6�ȝR=t<V�gK�'<�ol�h�����]{d8�!sY�%�諀�s��� =q�@�5�B+D$�ȜI8��۹�|�k�>�e4�v���?$Z�Y
�#YJ��`����ل��"	P��P�H���G J)��s��'���f��i���HG!ҎG�}��h\�z����>W���
��M8�x0��� ����>��}�~�ϫ ��h�L����2c0�H�$�Ls$N��=���5�툍��]�����<&�:������f]������9�s� �@�����R$(ԍB9������|� =�*@8b��>�ܼ�@{�� ����H\s4ڮ=H�Ǌ6I�G���@��{�rN^��ܚ}XEXr��I,��+����;����yggo�ʈ9ȜI8��۹�g�ٜ~����@��k�>����T�?Ѳ4(�h�v�����vD��g�"^�3<��K���mX�Y�#YI�3@�^נ}��h\�~ϐs�ۚ�� �"�B�3w�@;�1�qR�������ؑŝ<�6�N6�R]�z��H\s�@��T̬�2��UT��]`tDB�>�ߖ�]Ӏ~��h\��w���JD���G3@��-�{_I�s���UG�����T����̖�@���õc�F.y�.��{N�n�]8����lPp1*2\��=�����z�)�-�3rC�N��=���VrɭמM��[�
v��2![�����W�ǰF����VS�v�F	nm�]R�ԔLXY.7<����ënF���v⊬t��y��o���w����Z��	 ��W6@�<W��E��b2jR�S3���	�U�>����1���g��.kI�sqLݎ�Q���d�����f�n-q��[F������7� t���8�ݎZ9r�"q⍒dQ�@>�@����8�V��;)�TR���,��NM��v9hs� t��o.�Y$k"�6�s4q���vS@>�@�����v� �ȣ��i�"�=�`�=�j��v9h��ﾯ��߻��yw$�'Xu�o�k�`�ۑ�iH�c�,�'���	�ʷ9t����w�x��ڀ�8�ݎ_���9�� ��+��cq���7&��;w7~6�wf��4'w�1\ &	H!�U6���OV#� ]ϟ�@���� ������ւ���/w/Mͤv9hs� t���v�h�a���" �4F��>�e4�&�=�*@wc���\�Eѹ�[w��[{� t���8�ݎZ����s�@��l`����$3��f�>�;���u؞�-��ܡ�en�ԇR��g%'�wE�^��~�*@wc���=� �[4������dDM&���}�@�=� �I�s����36��.�*���� ��`�7x(DBP(�x�AE�
������y��-}���i����`���t���8�ݎZ�����Z�Ln4����>�n��>ՠ}��0��� �(��;��<)��I$�+����Og�n;Y�fG��u�Zi�z�*�9�r3�I�(D�Ƥj����-�vS@�����8�#�*,�l�>�73m�{���g^I�s����/j��E�qdI��˖��v�hfg�}�@����."�X�(��Q4���������7i�����	�	�c1�D�PO¨�
��]�ٹ'{�Y���d5une������sP��� ����~{�����v.�v�aa�շd��8z�\�͙w5릌v�G9�u�B9.s12�o3wo���@z�L@{�U�����:y���q��`���>\��B��Ok�X�>���ـޙ�2Ƙ�ick#q�s�s@�j�>�e4�-z��I�"A)�H�#��脒S�o� ��� �>n��׋ o��-xDd���s���r_y�$��hԓ��=��;�UUE������  쪪��UTW�  
��  U�Ҫ�+��QO� ��`� � �"�0@��V�F"�1
�1 � �"�0"� �"�1"(�(��  *�T@?�UU��  ��@ _�UQZ����  �  ��� _�  *�� W�  
��  ��  ����e5�E��<#�� �s2}p��{     
                �	A@��  ���UUER����$
TT�A(H ����( ��`   ��  ��
 ���ʾ�s�y�3�{MU2��o� t���ﷺ�N{yy4����}� ^��-��/��v��sya+������}i\F�g,��g���u��k���r��}��x  @@(2` }�r�,���0|�rzW��BA������iw��_Z��[�x�� gT�bh"��t�*�j���U7 	a�(�      0 4   P P 1   �t8�U)� uJ�&�TťJ��t�*�T��8 (AA@ �`	t���*�ҩW-"���*�� .�s4�U��*���R��Ԫ�p(��q|�۾�����[�>����/��
����s��g��5���|�N�6�� <��w�|��o�^�<����ʫ��  � ( c` >��9�;�[��_O�ϕ}���..��+͞���ӭǹ�|�};�..s[�{π ���k�Ŝ���s��sr���n}����]���\>�w��ʸ�}j�mUW�UW��  P��c`
+����u^.��r�w���O}� =�zru�]�s�]��wK�]}�>��<
�����W7O�������{���m���Jn��5������W��}��[�+��)}�yz\�s־��W�x�(� 4�2��)JR �O����JR�  O��'�T   D�*�"T � S�BS=J���F#CRԔ� ��?��?�������n����K����t�����v�TU�f���EPAWh��*�� ��ePAW�AXTEO������M�n0��	0���t���42\s5f�/�oV��eA�0a���Bb�&,���28ԕ���j0,tx/4�ci���|q]<��3|h�gBA���F��u���Đ� "��1������� a��B+����?9?�ߗ�z��i�H�+B0��u�Ѹ�;�/�Ǎ�{��4Mp�+��0�`j�0�0�Lʙ#a�	�1Ć#1%r���c%�İ,1!���#0$��4��d�5��u�3V9��q�ջ.���9�0�f4Q��F�#[7��#1�C)��	)1\� )�b@�)��d��`et٦RuF�!:��IH@J�L�$�C������xF�~*14ˊV`�`#�4o�a���7$�H@	A����|��	�>��L�G|�7��y�=�y�0�6'g5���k�s�~㇆>�,0�ٟa���1��l>KԘc ���DX�D�����==�a�n Ø끽��"*b	r�V%E	R{*��]'�J�y�����8x$F�,Jouar�~o��C����$�x�QsZ�Ӏy`�"B��>�N����IU1==�O���14l�Q����Hp2��K&�Y���Y�,ћ]x[~:�&:������0c9�����J=��IRT�C@�H	�B�@����Xp��5��x��^P @L���1��=w������D�%&sZ-�~�ϴ����%���F�a�$�ӛ5a�Fy�^a���X�H@F����{nּt�d�{��DT��&�.�1�fZ�	�KnL$ǁ�:���R.@a�3����ֳ�9�Fo�8F3�)�M2���X�A��������y���5�<ނ�F��fSb���Ff>�>�ֶ�O���|pH0R��##N�I��ͤ�h*D�!�I	!'@=���O���F1I1D��͂NI�2�S��N#9a�s��L7����}���C*Y�Ӵ4�� :@@�����-�\��_yG{҆�v�])��/�3W����p
$�㰓�������(��CQ�1��5�Ϻנt%�IL%D�2@�@��2RJ�d`\d�IBL'K�V��`i'�I$!!��#8)A��Bc�r�f#��I8�1`D�#$�8���I�  ��`����8��Ӱ�F�'g�����b�y��.H��5�'�f�SS�l-mHۛ��\��[�溢/ޞv�F8����q�d0La��G-�����,;�݌`N=C@��@2�m֦7��$2=t,�`���IM�$jׇ(�LL4��)t�p�(�=��E�0�Z��' � d ���}����f��E�}���l���5��4[�ke�����D��$�Pc�a���2��
jS`i��<��x�Q�!�Y�������	0a�3�����ˆ��TRk^�a�Fv	�S�l��t�a&aB�94D!
Q#�QL����4���M0��ə���1�L�,�u0��a��Y��MMil��_	V�{4Z �1�cD�5�3S�a�ysXVU��A�$�XSh�=;h6Dj ԙe2B�WhJ�5B�	
�cW��B�>��"��ʬ,t榦�cE�bY�9���S8���9;�r���N�3��Ju�4d��h�Z��מA�� �g���>t	nt|oF1�T�	6kO#��_pݳ�g�DP}��f��`1�4AP�D�8L������G<��ޜ��M�'48�0:����~@�HX��V�p�y�x��V��A9�L��R��3y����}�Y�e���:,t�A�O��TAch�F-�A�;$���5�$�Ѽ9�RPRDG�$�,L�4ɀ��a���N$�	H$*v��y�-�����񁅫���>����}���| ��A��ie�&  �q���9�5�fYf���L��KVVZ���E���k1��F6dB2sd.: O��M��\���M4�bG��#���ll� �0#��Ibd���X	d�a�Yf�Xa�p�$��d� ����L�h��p!��5bY��������Ń8ScX�,e�$6:l,-2� ��f��i,�:��4�$a�%3Af��ba1M�k5j4ku�3|U�0��|�t䞇g���h$�a�Jd�@�2b˔H����%A4@�D$��0����p*cA	�C�2�6�k����
�Q%$��I���.$�:�	0㲍��`�Z>��6U�a�k��>Ȉ��C��*B�E�c��ǹ��9o�i��rRYX1i(,��,��m�ךvb����Ↄi:Wa�\��l���p熯lK!���#��ٜ~����4�$��b�I8̬��,�8N�:�aZ��sF����20�	hő�(�$���MI���qe`�Pi`p�
Z% �aĜH�d��� �׉�!�N�-���o�=ߤ��1��F�l��9j�$,�K�A�=��r�5�������H�"J,�\���f�l�^;����>��z>����a8�b�&L,�3�.���M��[5����) �@F��% �p�������o|u>61�FX�A�Ä�*JL��g/4}���5��Kl'N:��:pO�C�V��i0�֋� Ѡ=�3���<�4l�p0�
'@�$% H	q1	 ��Pʱ�"'��p�K�:Y�4�ER6:��]3�40�$�8I��8��h
$�d���34��q� p8ĒP���q�0BLYqBV$60c0��$�̒�bBI���H$��T�$�32��rSt) JI$ld�p���1��:���#"-k	��cX�pth�o��o�|}�m��lл�X���;Yy�{��=޷�����e�2� qF�������4����F�99U�y�k�[5�k=H���p�����ϛ��z���,B`� �w����{���� -�H           �`                    $  [@ 	    ��                         6�p                       ���                             ��       �6�J�}�J�¥C��2�a�V��    /]nh��k�8 v�HI��[Kjn�L  ��@ �l씫5ٶ��	ѴS[�^Ͷ�*@������ E   GP���f�Xmm��n�9 �,$��m�j�1�EN��^9f1q�62��5:  ��6��m��:%�R�����|n_Q�6�ޣ :@    	6�' 5[��m�/i�m� [Uch��I.۷8[�L�l8&����Ͷ �.� :���%@j����U+��� 	�4P m�l H�b�� -������z�$�v�K�m���� յ�m�  h��m�@.�5M��ۛk�4��@-�q��&�$��l��M�  �j�:$�caM�  �m�4�m�հ�඄�"]�2�H �2ɦm!�f٪�����²���]$�5��6Z kn�bA�[UX  �,���R�l�Э�:岭ҭ+��)���^���� 8C`*�)Z��
q� Ň�8�H���a瞍��X����l�l�(���� V3��S���p  ��l6��7m�-� H-��C[�M	���[A�.��tQmְ \�Ym�ٶ���0���%��-���� ��i�� -�mڶlIm�~��-�h�F�l:�[{m�Hm�M����M��`i��Ju��m� ڶ�M#�n�H �I& I � ���[@ �K�U���s�,����mpI $ݮMMv�[�� v��v�o-�p
P ߶},�}#(�^Y�5Vp	^�VfٹH�]�	Ĳ�m7u�-�p  <�h����Bm������Ω� �E����$V��L&*�r��T�ۀ�T@m�kY������gK�	�^m���/n��gn�#[U/-*�Vԫ*�l�jm��]ηa 7i�����:_��-��Զ�^���m&���6���n� ��rC� �[�UU�u�Y0�@n1*Ͷ��հ������5T���z(R�9� �ͷ� ,1��$��E�   ��m[H��@��x�6�-��i�H0���uQ����hm��N� %sJ�h���X�[j���m��m�-�y��Ѧ���m��6۵�   m���V(e@@�@V���ዖt�m��`m��jֲ�R�P���z��U�j�m�ݶ �Ͷ�N�U[T�[�YZ���í�6�68��t\7�}��J�7>h�j�"��%���k q��ml��svٶ��E��Zq��\Ib�����uq�0L
�n��۶���е'�ͺn��ٯ(�cS� �5%�Y���mm�   �5�2Cm��>�)Mk�*��[m�怺�M��[v��p 86�  [I�]c�lȑ�Jm�E[tIF�%��e� I��f�q�k 6݀��8�$��  6� -6��P�Iz�7%m��}�R�̻=UUme��$�ܳ��l6�` [@ �`m� ��� ,0H�`��jCm�qm   H    H��� -����l�$�p6�p�H*M�֦��D�IS[�� h6� l � ��  �J �m� ���hm����j�U ��      �-�  �  � �$ �	   ��6�&��-� m��� �`���s^m��϶�}����\��v�R�*���}� LҒʃ����6Z���6�6�m��� ��Ie  �   ���  h[@,3i$ض� Ś�l�m���yv��e�d��V��R�[������m<f�5��zݶ �(�)�k�Vl
PKF�۶���Cj�ְ l�l�YͤZ��7i� oP 0%�횗���[
�q�n^X�!!m  m�h 8  -������C��U���ՁCm��+m�� 6�ׂۗ�k��uҁj�s[ �T�K����I+�I�U��l��4<���Š�6؅�s�Ē�$*�|�S(�qO��]��Pm:I-�[s �	 @ �km� �"޻��mI`�V�8���	̽v.�! M��uV�̼������Z��9V�V�
�Z�j�U5���%l�Ӗ��5�ɋd�6�C����z�I�m���M���k%�%�	 �kd��ӵ�Ͷ� �l8M4���l:�0-� �U[�`��������� ��M�J�@����תLk�-6	 ��-�mm];i 8[B��h -�l�6�* �A� M��u�VIݳUҠ=A��qR:Wc��	Y^R]����M��M��@Im$ �Ԗݖ� H�[v��Y�n�f` �M��i6��V�H��� �   ۴�� #]��J�KJR���J�mT�` mm��`!��!m-�?����m�86�F�H   �������We��6�b����VUU��6�U�| 4 -�h��mm$ [@  ���մ$ �� 6�m�@  H ����[���m�� h mж��e��` [d�  ��� "F˭��i�  "J佋[mm�m �b䭶 6�H�of�6�$��L�   �Y%���L���` �� m�[m�j�t   �^3mQal��v�uV�h`��n�
 ��KQR����t�XbZܴS`�i�v��t�v3.ʹڪ8A��W*�6���!�
N���++_��I�5U� u�-�-��-�յv�K^���Դa�tt�N�� h��  �v 8���m�p�)@ �d�iMsa� �r�6ض�� � 6��ܻi�Uv� ������-�-�ٶ����� N�m�I�^` �5UJ��U+�4��<�����3mT�		 ��v>�}'�HI m���lp���[z�[A۲�4PͶp[��Cm�l�����|-)L�UW5
�� #�Av� 	l�b�@��[�� �l�X���v���Z�Z��-"E�h�8Ŵ������Ӣ$e�m��m�C\�  HL��ܫV�@j����'$	-�Z���l .ݘ�m���l[[m�[@H!�i1,���@ ����Z޸�    �`!oW-�5�Kj:��y���$kpmR�m-�M}n�c��   h� $
V�;��;S]@R���6�h�6�6ٯV-����u�@ @�  ��8  m e�	z��e��4�P5�5� �[@ 6٢�   � �F�H�n��-�m#f�e`+i�R�5]N/Z Cm�6��    ����g  m� �vͱ�6�H�� m[[y"��Z	6���pT��(m��kh����� }o�|�� @�! m�V��-��[VӜ $I�� HI,��l]���`^�j�m�` m�  �l$v� �@�A͖��lR��JKztP�&� �l  N�6��
 kX�����@s��5��p�i٪�&�]�UU[g��6�) s��*�����Q�i,� 6����[MmY2�B@6���P'6ŵ�ͻ` f�Y �m(6� ��u�l�հ�n ��	V�r�˳UP �K� [@ 6�ɻ[4�qm����l  �>$6Z=#m��+�  M� Z޺U�4PH6�Imm����C-����[m�"�/  �D��Amv�.� 5���mC6m�[��   8  ��em�@� ���M�-�� ��]5��.�ض�8`�-�@ Ia�Z摶   ������Cn� +����UUJ���}��{��T⠺P� ���@'�)"�D��@�1��4�$��?��.?iĀڧ���>�&~W�_UT}c���{���O�!��WBl����E)�h|qS�Q�*�[ńځ� 'GA� p��@8��C���@��"��W��'�*�� �� ����T�������'��}���q@"��>h4��q@���4p�%P��臨o�
t����)��Q=C�О '�Qx������T��"l�h�O�$ I|Q�l�)�& qDIXt��/� <_c�G��A� )�;�|]���x�������@�(�m������<G�C�6��uD=AG�v���o1� W�~P��qS�Q��= b�!A�C��:���E�:SB( �G@� v���ڨ� �M'�*�G��?�+ A!��f%�pQ�e\%	ݽ����@ p   M��j�f�    '    m�    � $4�j�m�^�s�J���˞gj�q�e�{X�Y
ym�e-��X�PQ.!'�{��=#��s���h�������ҘBtM՚keaT뜆*��lc��aK<�9y۶묩��pOlb��v��\a�S��m�4�mWGD��CəQ�=��&xL�W`�q�γ�km�+�v!vN��8�ʲ�=��;d����g�4�hvp��ѝ�:�I�t�\=�зHm;�
.�&ό�r��	�v�\��;�<��m�#��Z@_�m�*�:71vղ���$6�P�����������F�c3���̖���βH�m���\�a[m�ʯ���
ٵ�c�;[Q���)�@u<�(
�MR��P��� ��F���H[׭�^`W:�r1&��uu���%H��P����m�5�<Ƀl�܂T��f��]���B�R�!����2�a��O�.1˻hˤn���HɹR �v�-�;NnR,�%d��N���7��%t�+������� @:�[e�C�˴�.3���cN�,�z�nZ6v^l���0-Ғ��ڥ��溁�,����l��` Wj]�>Z��V��M�ppT���[����4E-�kYa��[&����G�Tŵ�ls�%�r�Pb�F�X#)[�Lצ��:#�m��rnqhVwc.;ۚ.�D{!*m�nRWgv`�Ypf��D�N)xn
�SZ��rN� ��'
�\�� �;\�-�5ִ�J��)���x�(�Z[H�ѓg��bA�e���q�6@@���W�$l:�9y�H낪2;\��i�Za��Ip7`@
���n�wj�i5=�U�gMҙ6��r�+ ,J������v�l�_.ܖ�:6 kiM:�]��[U�v�+�-�۝E����ʛ�M*��!��/�@��>|� ���"����`C$����ֵ���`�6�k��W9V�T�ȪM�&�W!��`mÓ�a��wV�a4kk�W�!2�>�� �jH��/J�9��KS�K$�)�EnQ;.�@�m��:�$����c�m�yrܼ�ȝ(�9z��A]qHؤ�p;\�7j;���cs�-e_=b�\K�Xc�#C�.�V���޴V��8�6ۜ�6�u�{����� ��p�Qjә�Z�F�,ֵ��n��y징wa��<�~I�1�!4��ǟ%����;��s5�3�N0
��Q]]�#���Wj��f�{_UW�F遺����f�}���I�x�q��9l	�07y�q�L��f�`�e�ƛ���0Ć�π����� �����UV{���3�߲���ږ�˺�0	�[ ��l	�05f�����{��������C�����Zll٭�u��ڍ1lV��x�+y����,�� �46�r|�_M��s@��r� ��h_ԭ�1�"R'��{Ú�&�]<U8��}���U��ޚ��9�����Q�f��6��-�vl�ݎ�A"w��48�j> gs'5RI]�w6p��.�W�ص�n�Y���)0R)&�}{f�{۹�us�^�gs' ڪI/3snզ���j(����ݕ���9��Noj�%&8���Chn-��G��Y#��=o�4�w+��f�}{f�v�li��<sHi��l�q�L��f�`M������#֑����<o"hrdz���@>���/O�IکJ�����y���e�>�^Q㱍A���qɠ^٠^��h\�W���쿩[�lc�"�8��/{w4�w+��f�}{f�gyڒ̏�4���,�7;s�#Fت�Z�U�U>+��$9�LS$M�	� E1d�f����zyl��l�/{w4�Z��T�48�j> gs'5U�wsg ����\�W�i��9&"E&
E$�:���{���R���-| �n� ~X�t$��IG�^��hW�^�gs'�T�
���U.g$���c�m��<sI�9���z��h\���n�ZU^<S�<�<��oVͫ7a5rU��x�ɴ�	�:�,\�G;��ı�yC�#�������^���8��_�={�_ ո����Q�ۗ˶���ݎ���� �%�����_ԭ�؇�E ��@��s@��,|6�$������l���[n�v�"���3@��r� ����廚�-Cƪac�Ǒ�ݖ�;6[d���ډ�����{�mh ����ޠ2v��Tr���2��J�䋦ƍ���t����u�[I�˝ՙ6q�R)���]���.6�ۘZ�&�@}F9I��r�l��v�A5�QO0qSv��Y���Cu��e�������3v��n��D�`x�#%TZu�!�#c�3�Ͼ���ዄ�������8f�xc��!�u��c�tS\��eY���_}������sf�F8a�3�v�w.z�;T�9&r�d�5yC�KQP��ܓ�"�t��M䎘�ډ�M�l�*�wb�	����廚~�\�W���@>��@=z�Nx�l��v��&�ٲ�$t��[|����-��Q�>�T�]�f� wsg �[��us�^�\�q��� �<i��͖��#��ڜ`v[�W��??���;���]Yrӷhƭ�8ⲍ��̜��B��UVܷ�,��ݷ>��P��U����w��z�叀�d�I/�v�h�ɶ�&H�DI�W;��� P" zou�s��W��' ��8������w��.&�_�z�f�`L�遫6�\�YS�b$R`��Mfg���{g�05f�� ���jB����pk$�h���W;���l��l�;ZJ��ibi�naCQB\���C���x�S��
αm��]�\o���(��9��9�Wny��l��l�/;w4��ti���&�&G���|�û�8�o ��� ?a��ݐj4��nN ~�d��g��z�>Ȳ��!�=Wͭ��:y�T^[4���oF���E"qɠ^v�h�jq�L�l�e�76.s����-G�05f�� ���f�`^v�hu�U�Pn2f<	i��9���qQM��Evv+1N���h�@sغs��%�<ǃ�#��٠^٠^v�h\�W�s�eRI��I��94�e�}_|��t��e{�f�`�t$Ȟ�5�I4��������h׶h�:�Nx�5��q~/ص�;� �����*�*��ff~��y�իRMD�7�4��#�	�-���������t�՛S�����x��q��]<5�80�h�wg�-u��ٹi�4ޱ�$���vy��g=(�]� ��l	�05f�� ���e�Jލ�����&�y۹�us�^�^v� �����M����"&Wt�՛S�f�`�-�3c�ʔ1V��1�����h׶h���W;��\�YTrc#RbRI&�}{f��v���
�s�@/>��R�(@�C0$2CFw-ߦW.o���� ��R;Vۗx�vzn�MlIDK������ns�y��
�)�ݗ�nf���&�y��zڵHB�^Q�cnA�jpc�k����6"�u�h�[qr���)����QQĭ��t;	ܹ2�+.�k�\��]q�����բ�v�y�6�U-
�W=5ڴ�tY�\������ܖ���aɨ� ������w�u�.��܅�6͵f�]��]:�y���Vj�9��:\8��{s�$$n�dׁ�@��t�՛S�f�`�-�w�ʞ�d���6	��
�s�@/;f�}{f�y۹�^�ڒj$����92q�L�l�e�&lt�՛S���5\#C��m6�����n���>R��]�}��~YXck����r�/�l	�05f�� ���f��m����>^����w#@�sG:w�]W*ݫ�gnx�k �y��$�uiBW���E��wLY�8�&l�ٲ�}���.��Aӽ���q48�| ��';� z�H� 0΀�B��q�P �*�U����\�W;��\�YTrc#RbRK�`�-�3c��ڜ`6[ �\�� G���I&�y۹�us�^�^v� ��� ���/�Y"x�5�йu�"�^�)M�ٲ�6:{o������`���3շ�����j�l��GP��3�v�l����i�$�Љrf�`�-�3c�,ڜ����!��6�RM �������;}����*���l��:���e��n��-ܓ�o�x�o�X�~]���$`4�N�QX���k�x�j�I���L���f2"L^Z�`�2.���y�'5j��S*+��1k�O%َӯ��O% ��H�Q���b$��Ï��^xb��先�
�l�����d�ы��iB-mC��90@���%9�L�>�꧃�:"�EA�S >$B~ 6��>�:*/�(%T�PG���o���W���|���[n��	,�C�j����� o�g ?w2p>��ʓ�7����t��h�C�G��p���_��f�p_|�����Ck
إ�V[5t�6��[�[e砮�7UF_V�$����c��f�#5G&24���I����y۫�z��W�}�8իG� F�n�+���M���"-��0	���;6�o� ���O�p�� �F�s>��?��7$�~��K=<遾�t����Z�0o"bNL�Cٙ���4z�sB��w�+U�1�DCP*$�U$�T�R_���]| �����K����p����_W�T��-��o7?��}޸�έm~QI����cs#�(�a�U�vi��RY�C2v|�2K����w����F����E#�����x�:�ܯ@?w2j�T�Xwsx�{6�w��Ie��9!�=}��ͪ��vp�o �}0�Ծ��Z��;��#E���Q���*�g�O�wsx�}w����~ů����U��R	I$��\��٠w�ۚW;��yl���	<m�;�H�s���>���������N�����/km�&<m�$��I$���J�뜬g����{�⁺t�1�q�]�  ���;hSvz���`{XA�gXSR�/3-u�����H�R���]��n[E<��
dXȠ��k�9-h���]q�s�����Q�- I/�Z���ƭ�!�a���3�7���VY)�-*��g�[ř'1�*73\+�du��+1�q9W-Y�{������v�{��|?d;+����Q+q���ݕ��Hݶ�n�܃z.�m7A�*2]��~�߯����9N�m��>��|���N�=w?� ﯷ4V��MD��yrdlrK~�#=<遾�t�՛S���$����L#kRM����9{x���|�UM�毟 7>�p�+�_�ԗ#���m*J�W�g4�~ů���8I$�����p��w�n�E`9NHp_|��J����v~����s���9���[lI���G&A�T�YL 붞֊�ӻ\�٨X9n5��=��w��n8���O�S<��wޚ׷W �}�Z�%��/ص�ux�m�"f��ݙ��{�*�w�=E�� �0���㗜��6�V� ~�d�ʒ_Sa�����	<i2"I&h_=����$����vp��. w��4�-;�7��%z�~ ;���;��.�_o���c��Q,x�D�N8= ����7ۛ�~����=}��R����D�#���3��lXs1�:�<(�j���i9�n����������n�w$�����;}�>��{IR_��vp�R�Y�||ڿ�����r�_���5��J�]�~� ;���;��.n~�����i�M�D ���@��ƹU���i �+ �B ! (��=��}Õ}���\��1:w��.&�U*�w�n�������iU*�~� W��)$�H��I4^��ٟ�:�|���@>�@��,Xآ]l�a�8�v��9:��i���un��)1ķ��X+�Q�?f%�4zx�dD�L���>��| ��ɵT�~����p����\ Ӑ��8����h��T��IRM��� Ϸ�.���RUJ�ٸ�6��M6���q���ݜ���ᴩUU߯ٯ�e�u����9.CQ�Mܓ�������\����=}�|ʩ?'��!����CO�����o�{��5���8\�[��v��|i,~��;���;��.�*V��ۻJ�MD�sI	�N�c�%�с��k�F�]�����<����wSmjM)�s�r>����~�d��g��_�_ ��4˽j�E��䏀��9���3����e����Z������A�Ϭ��1�'�Iwl�01f�3��E��o�l�r���4�$�4.v���� ~�d�mU|�����ٯ��p����8�������W��}������;�������{���O����m� 6�tv�.�6�I��Ӓ����:�?�����2�u��}7N�jA˼f���L'=+Y[]��Q�M�[,�L�cn��P����J�WOD��3�h�k�M�=4�Y皰�ȥt�+���z�uV�hnp�3��]'�.I���[f����R��7EӑE��u%ҭa�9��m�.S��{.�n�%�K2L�n���N��Kv]����^�� n�93s��q^��gN����ܻ=D��;����L�s�ȚI� �����۹�qs���{u��U޽#�����.I�;��.mU���k�~�| ����I%v{kCY�ݎ�.FG ��5��s�����ݜۛ��=��ݜ��X9V�|	Z�*I�����vp糋��*��_��_ ��4˽j�E��䏀��8�URI{s/�z�������o�����y�^�#v[3��ZG4��#�v��E��K�mj������w{=N�j�H�s�|}}��qs��\������`w۳�Z�ziݲY$��U�{�uΠ��"���]!�ҪQ*�Z��]����| �f���qsiRWa�f�����Ӹ�q�o>���s'�U߷7��z���{����<O"i'$z��.v�h������5+����x�Q��i�n۷-��c���l�:[�q�w6[ ���qں�0&ٺ3�ն�0��݆�}k�R�U5�-�J��n��>���"�Xb���Uy��������̟U~����4���F��� sԏ@��}�]�}�8�7��v��|�J���4˽vF�Dr �g �{8�1UW�AOD$W!_P?��}�?k�w� ?.��nH�%�6�rI�ڪW�����ٯ�{�0�j�w�n� yj��H�I�I3@��k�=�+�� �}�r��h�%SŊ��4��2�6�mNK]P�붟m\�I�:ض���W���x�O���?��X�q�����z�-�����U~���5��y�v얚����� ?w2s�U|��lϷ�.������>mRT���5;oI,i�n�$���.����WʕRoo>����Ӏw>[ۧ�B�\����ٺ�]Ͽ~�*����+k�!����V�+Ē_��U���ˀw7�m��n�@Lw#���>�RK�I�>�t�~��9_j�>��x
�s1�m�)�M�{uH�֓$9���b��1�c^z[�އu���G���rG��4^�����g�U�y�	\�g�rc#N��I?��qsRJ��k;����w2sUR����ס�M�%�I ������>J�]����=��\ ���Y�t��q����US�o����� ���>K�O&oπ}���vKM[R�v㏀��8�K�U�������r����\�F��2@�KG��7ɁⓃl�MpL J[e�@���[@�&��i�`4�&��!`v��(oN�YHX�ݙ�A�f͖�BI�8oA6kdf��6<���������N����m  �   Ko�(     t          ��	4��ʠ--٠¨L/�[luHMF��fXw=��l�7EӚ��T.8�((�5�l��;q��'���*�ݢ�!���G���e�?v�;�Y�"�e�u�FK%3/Y����C�lm���5��c7��wE�c���Ӑ�Y���p�����Wh��[nI\g��'+!��Y�v%�ӈ��
g�C��cldH�+㳻,�C}��<��s\�q��^��� m9�P �ة@U5"p�t"�ԅ�����k8�b�����z㖎A.���n�"#Iň��6� @����F�	�	�$�ڱr��v�\r(���m3H��u����l�؋N]�4�V�[]����
��@D��p:*\����M�]���[@)�G�6�u�+�+6�4)!c"�.�4��q[R�5*�甙t���T�R��k��������p�]��Tj�a�s*.�b$��P��x�%dLh-�m�N�=��um
���c�c��Z�b�n5j�mR	���s�ukc��cm���ݐO\r�!�l�B�^�۶�Ǫ�Β��8�[m��� \j:�	�'"�j$�F�m$�.���A��d�˱5mKVԇ+�J�E;����E��+mVvN�'eݪ�E\ۧ��.��Ѕ,�����SA��m�v�ڙw
qF*`����4Wg5��v�N���.7n3����spç$��Q���9�
WiT�e-�Dk#Eo��o�e���uJ���K$P�@Pu�oUn�K���V��o���r��[T��8:�#
��PP�ca�	��Y^���9�^�Ƹx�J��C`�H�m���r��4�5.��_}�'����*;A�g�Pې{�M�:����g�e`b�r�UR���m�W8�r�_/%��Kd6,�K�ȗ����9��Ms_{��������������^���Ȣqp�P���G��	� :�w�D6�v{���������2�p8  -�v[�[;�MK&���S� ����+�NF����\�h�7����m�5�ڑq���v/OZ�v�<F;k���>6�*մ����Hpq�:`��7�.�q%��)v�ڕ趮��z��u;��
J�Mh���5{k����h�G4�k�U᭗Қ���䌹ش �
���8��`���&�{���������k�l�Nv��\Xh�m�W=��-u���8j�z8s���X����Fy�A�_ݶ/{��g�N0͖��P'c�t�rI-��=}�>$�/�>�����{�h^׾H�o�m�L c���Z��y//_=��=�L��xG���'"��fb\���6�5�_}���U{�6���fے&In���p��>��%�ٯ���h׶h������a����sf�X��g��.����ԕ.��\����k�����&o�zG�'P�?����@��/���>_*�����ߟ ?�ߥ��t�,�q����o�\T�~T�J��:U*����߃7������=}�>mU*Wf�6��i�j[-[���͜/=���U%w����7^m��؝���4Էv���j����k�~�|����ڤ��w6pj�m�t�rI-��=}�>��������8o;^��j��JLk��q��z�)��*ݫ�K�����v��l�ܳ���o��M�� �1��U�y�׶hW�����䫬6�~|��`˿���q49#��l�~�Ď�_=��=����ff$�Y�$���N`�W������j�R�j��KiR����k���h/��Ly4��q�f%�T�f���}����NV�J�c~�p����pm`��nO���X�������}���we�6H�<s\xx]�ڶ�k=��[tɎXn���WP�7m�v�������{������\]c�8����hW��������
��= �O{"n���M7��{��-��*������)[Z���RI�@>�l�:�k���4+��s�m#Si��lRM��_}�r�����W�߻�W���@ XIE�$�@L�
^J�$�<�͜/���^���q49#��{' �J�y�k��͜�����RX7�5���c�9�9�u���\�r��Wn��{i��nj��b��&���9��hW����W-z�{f�s.QЙ2<i8%���e�5d�`ݖ��6q�&�^G,m`��nO�������4+���������&9�!���}�-��l� ��lY'k$�W�!1�Țn94+�����O�����W�}���2�� �`-ww{�>�����\@ �[n^�dY�2vj:�*�HfѴ�/Y9�(�O�F�k�K���J����!c$Tu˻��;tNe�wk��g��J�I�YV%6Q+l��fP\���N��ĥڞtV��e%vK�Xn�.�	<�Y"f��ΓG$�i�9��3d�]֛�>�}.��.F`6[ͻl��mӲ��8��粖m�����4�ﻻ����������O�y�#J7'$Q�&(�E.��S�˴ĝ�vet�^M�D�^|vnIn> {7' ��1���B�RIrÊ����M�jm0�9��ɠud�`�-��l� ��l�C��xG���rG��l�8�k��l�:�k��
ʤ�"p��h��0��Ւq���O[ ��x�QF�ۅ�#����8�R��ٟ> _{�hW���R��caK�����ۡd��7jT��܃z.���획'��_�������8��.I<׿�π�-��l�﫨���5zy$r՗Zټ�Z��o\��﻾p@v"�����%�T�8K������=}�|�*��$�{>�K�K��Rݦ㓀e��> wd�z�����}�0����}��M�V�ێ>�URI�o�N��|��{'RI_���f�|����j!��˶���7e�1M�`�-�~w��~*��W';�]�F�t��.l�F�X{H�΁r7-Ʊ�Wk���q�������<���}4+����=��3�w�z���yI&2E&	�I4�{>��U6߾�o>����Nm%�s�1�&L�N	B8��ޚ��{�[N(�<A@�D���_w}4+�= �^����9�N)$�>I%z�ߟ =���z���UI]�7f������2,M�H�����K�����=y�|���?c��n��b��5��j����槂�f���M�ncD䫩hvy�NY��z{��%�5M��_}U���`{J�m��:�6�q���'6�]�{���͜מ�ϕ*I/��37�o��ۻa�l�' ��~| ｓ���������>T��cm�#ǃr=I+�fl�{���ٓ�iURWKk=|�;���Ld�L��hSgvK`j�8�3v[���p��������%۪1�뵅G��F��s	Ր��c�%�<R�]K������]t���@=�}8�=��w��z�Xe�u��q����8��.I? o�g>J���<��~�|�����_U*��k��wn�"q;Vݑ��3�_ ���ڤ��_}�����ۑG"ɏD�)Z�J��5�),=��p�AT��r������py)Jw�ۺ�5�̴赭k7�qJR����C�J�9�����)>�����JS�����)������~���E ��Xu��(�nrh��k��Ě)�`ɲ	�'i�x�ݥV񳧪�v8�jN)�+��D��qư�s��c�\^�[�,�ݦӡ�2<�l� �BM�\����6��[�-�a���D���H��e��5R��:�ɮ��3�k��������m�TK���h�J�����ɱY���쁡6����нr���w��t���f鱂u�;vx�Z]pf�u��[��v⻧���w��{�}���  �vnr;��)J]����)JR{���<��>���p?.JRw���<��=�����m�Nܓ�H*�R���j�/�)�������C����g��+�R
�f��U �AU�Ǚ�$��\�f�����JS�����)>�>�$?�������┥'����JSH����(ӻr���|�AU�	X��w�%)K����)JRy}��y4�/�*��g�>U �@��u��pv�Y���[��)J_~���JR����C�JS�����)=���JR��~������c����\�X�xn��$k"��նl��t�@z��:;2�%���3Z���~�JR}~����R��=�u�)JOo����~���)C�؝���4Էjӹ�H*�����/���*VHk�H�"i��I#M�Je�0�V��$@%XI�`�`��OQ%gr���{�%)K�߿o�R��_w�JR�����n�t��w#�R
��{��p�AT��r�	+)t�֫�R
����ʤH){��nGwn�5�c�5\*�){߻�)JRy}��y)J}��� mR�W
�K��͖�qٳF�[���)I��{���Y���\R����hy)J^���R������߁�<��O��%kXe���&��,�ӳ�&�N�Z,�ʯ&q]2u������}@ս��fh������s�ߵ�)JOo����~���򣋩JO��W
�H���QF�ۗw#┥'��wC�JR��w|R�������R��=�u�?��ZR����W�̸���-ƫ�T������R
JO/�� �CA����iWM�"mi��V`"H(���%�^���|� ���&S����z)�pJz*B4$)����4 �|���x�*/n��m��0�� ����	,� �f���_4*6Z܆2	�������2<��:�|=G�ԄT ��A14���A8�G��"��LLG���0ܧ3�w\TH)g�b�H*��<ywn�"q;V���9T��P���f�U©R���┥'�}ݏ%)K����JR��؝���4Էv���p�AT�}�|�T�'�}ݏ%)K����J� 
]3u��T���ۻ�D�K ˵[/bBѶ8�{��=��.��v�hZ�������wn��7*�Uj�+){3by)Jw;����)I��{���������R
��ٶ܎���j!��z��R��>�u�)JO/��%)Os�)I��wc�JS�������kFoVlӬ���)JO/��%)Os�?�H����ǒ��s��k�H*�*���˒D�.Ev�I�J��;��R����v<��>ϻ�qJB�����$���{��U#����"�4�ܻ�9*�U ����ǒ����{�)JR{}��y)K����H*�R՚���m5z��e��G-ݴ\�0li���s�n�fLʊ�$�N����Er��8��wn���R
�����E)I��{��)�w���)=��p�AT�y�˻��ڶ�n>U"R����C�JS��{�)JR{�{�\*�U/_�*��uHb��m�%�3y��Y��y)J}���R�����c�JS�����)=��t<��>�^1�;�&��qr�R
]�dU�JS�����)=��t<��=�{�ʤH){��nF]��ۊ���%)�}��R�~������R�����8�)I��wc�JS�!�
��?�h[@� ���y�X;S��-���,C�:D�8
�h�d�;A�C�N�'<m�:�����ձ��v�W=j�L��Q3�k�v�˳cOj�r�̻[�W 	KDY���}��a�x-�s�n�%�Hr�Y��諕6���ƦXm�.Y:����Nm��9mp� (nB�y�1�b6�-��]�[[���,nm�5۳��{������c���M��ۃ��uʉ���r��;,CK֚�m-�^..��L����^Ӌ�#?�{�R�����JR�����)JO~��JR�g�)C������������������)�{�R���ﻱ�)�}��R��_w�I�C���,�QF�ۗw�r�R
^�؞JR�g�?���>�hxU �Y}��R
�
�����q�f��ly)J}�w�┥'}��������\R��Y'���ǒ�����v9r'�m��|�AT��v�-W(�?k���┥'���ǒ����{�'�"��(J3�(J��J��(L���
�*^̛wjH��ܧt�p�����,v�]��-u�t��f�z8r���t/"�����fn޷��(J��0J��(H��(J���(J��"��(J�~��^x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B~�p��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bw]��^x%	BR�	�%	BP��%	BP�$BP�%	Bf`�%	BP�����pJ��(O3�(J��J��(L���(J!(J��;���Z�Yk5��k[������(J��J��(L���(J!(J��30J��(O�����(J��)�C���� �j���%	BP�%	Bs0J��(J��(J���u�P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B~����	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	B}���<��(J��(J���(J��(J��(L���
�*^����vݸ�܄�8�P�%	By�%	BP�%	BP�%	��P�%	BP�%	BP��~מ	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	��~����(J��(J��(J��(L���(J��(J�����x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'���8%	BP�'��P�%	BP�%	BP��%	BP�%	BP� *]z`��m��ˉӷ�ʐ*@��(J��(J3�(J���B!�߿lA�4?~�������v �D�%	BP�%	�w��y��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP��n�����j��{37���8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	��߼<�J��(J��(J3�(J��(J��30J��(O���pJ��(O3�(J��(J��30J��(J��(J������(J��(J��(L���(J��(J���(J��?}�߳�P�%	By�%	BP�%	BP�%	��P�%	BP���
�*_,�r���՟!	�6Ⱬ�ۃ.'k����	�:��ӓ����n��n�"�r5�ٳz5���f�����(J��(J��(L���(J��(J���(J��?�~���(J��0J��(J��(J3�(J��(J��;����<��(J��(J���(J��(J��(L���(J����8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	��߼<�J��(J��(J3�(J��(J��30J��(K�������av�8��
�*@�~���(J��(J���(J��(J��(N뿿k��(J��(J��30J��(J��(J3�(J����~�	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	B}���<��(J��(J���(J��(J��(L���(J�{����(J��(J��
��(J3�(J��(J��=��k�fZ�of�kֳZ���P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B~�_�g�(J��0J��(J��(J3�(J��(J��>��ߵ�P�%	BP�%	BP��%	I�H��F%����(J!(J��5�%	BP�'���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�&}�����(J��"��(J3�(J��J��(L���(�
��5;oI,i�n��\T�R(J��(J��"��(J3�(J��J��(O����y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	���ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�w�����%	BP�	BP�%	��P�%	BD%	BR�&f	BP�%	��~���(J��0J��(H��(J���(J��"��(P*[��[��n��CrF���RH%	�%	BP��%	BP�$BP�%	Bf`�%	BP����8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP��~ߞ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP�����pJ��(O3�(J��J��(L���(J!(J��>�~מ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP��~(	@X$I�����O��nŻnZ���u�6y��W*ڄ������:�-�ЉNMl�[7o5��(J��<���(J!(J��30J��(H��(J��������%	BP�	BP�%!��P�%	BD%	BP�&f	BP�%	��~���(J��0J��(H��(J���(J��"��(J�߿xy��%	JP�	BP�%	��P�%	BD%	BP�&f	BP�%	���ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�]���浭�f��[ߞ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP������(J��<���(J!(J��30J��(H��(J�����x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B~�p��%	G�*0	�`�%	BP�	BP�%	��P�%	BD%	BP�&~����<��(J!(J��30J��(H��(J���(J��/���O�hS�S'}��;�'{��t���0J��(H��(J���(J��"��(J�߿xy��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	���ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%g{���|��JO�~��xU �G�`��R7n]�rEʤE'~��JR��w�┥'}�%(>} Ni~�9��)J��ft��Z5��5�kc�JR���|R����a�)�{�R����wc�K{������� m`R*qZ;hp<Pt��t�
�j�۠���݉��sr�f���R�����<��=���┥'~��O弔�.����JR�jvސ�����\��H*�s3��?/��R�����%)K�����JR���]��(�`�S���j��X�cE�qr�R
_n�p�AT�{���);�u�y)J{����"�{�r;�v�ۊ�U©ɕT �7������)I���C�JS���8�	���jO�߿�<��>��Gg��m�L�'*�U ��ǂ�JPȤ����)JR~�ly)J_}��R���a�mE�����߫n����H  �+��9�ݍ���\:y�Z�	�W��V�#s�kan�X��[��lѹ-����O%�F�+�l4����Ɏ�b�G��ԣ��/l�O��Q�㛳��.{k[��no9�QQ��K���k��p�["�K��%���iז�\U�v�b�Xz2[i�*�2]	�Ѡ�Q�m, �k�����nK�/W0k+:�����v�wia�N9��37t�6 m�=A=p��+�]���\���2�{�����\�(��oz�?JR�����qJR��}ݏ%)K���JR���]��������Eiݹwq�*�U ���E\�Y���߷�)JO�~��y)J���\�[IR��@�}yw��m7]��[JR�{����)I�{���JS���8�)I߾�ǒ������f�ˁqKVݶ��R
�UUBVR�k�W%)O�~�ÊR�����y)A����uOw�*�U U�~N���M5-�n��JR�����)JN��v<��/��w�)JN��vJR����k<~a�u,ˎm'`��Zmg�ڪVQ�L�LI���4����ﻧs��\g���JR��{�c�JR���|R����d��L�R������)JRw���܎���Q]��-�\*�U#�̜Iy%�JN��vJR���w�)PR�{"�H*�����Km�F\M35��JR���]�����{��J�$�����R���߷�)J�����܊�\�
�U �R�n��R�)?w��<��/��w�(O�d���E\*�U#�0OB(�N���K�qJR��}ݏ%)K���JR���]�����{��JR��E>��w��]�d�R1�9�ma$��3��n��
ݫl��4�ΩMm,L��\���a�)}�{�)JRw���R�����H*�R�{"�H*������h���Z��o|R����a�){��|R���ﻱ�)}�{�)JR�/bv������.AW
�H�{'�)>���y!�	�<M�D��ʤH){|�U©R�-��vX�e�'*�Uh���3b�H����┥'��%)K߾���U ���[�ݻ���qB[��U ������)<�u�y)J^��w�"�/{�p�AT�c�m�EmH�3��N�c<l���c��Z��i:�bX�;tC\�z�^Ӌ�A������߯�ǰ�R�����R��}�v��%)�w7g*�U UՆ3nI$�܎=��JS����R��}�v<��/>�w�)JO;�vI�@!�K��	�Eiݹwpn>U �AK36*�)y�{�)O�$���~����י��H*�*��7�H���۲�U�JR���|R����a�)�w��P��� �$$XU���D<��7����)go1ݑ�4▭�nNU �AK;��R��������┥'���ǒ�T�w2r�R
Xe���ح�r!����8����6Lۚ�L^����m�����p������\��H*�o=��R�����y)J_{��R���<p�AT��a��F�vX�wm��JR��}ݏ%)K�{��JR���ૅR
���c�R�T��R
^���n�ݶEvℷp�AT����R
�	�{���JS�����);����TK�����m�F\M2ܜ�AT����vJR��~)I߾�ǒ�T�w2r�R_���2ܑY%Ȯ�k{�����߻�)JRwﻱ�)}�{�)JRw���R���4 ����i�d��$x54��0��y�04�B�a�XH�%��Li4�g��B1���!-����Ь AA�o�I��nh� xc �*�}�t\bal3�130�do��: RiM��|������� �   ����     	i�         hWP�\�9ZY�Y����6��F�͵U��zyCq�������p
Q˱ �:���5��m'"���I�;E���@wJ	c&�`㫝���]�xUɠ�[�y�i��G/m �N6����㭒 �3�<k���ng���T��ZV쭭�*]F8���K�p��z�m�Y�"�"�ՙv�vܬd����9ʍ;�S(S�����-I-��j� �f��l"��)zx��u�+R�O1E���n@ā��,�qƷ=�5�[,oݺ�j��$���̦vCk�&�]h�0�	vf=��ӣ��h�g�X:*���ѐ)�hX���8q��,uH�	�B湮�l�ÒZ�Z�mJd�:g(�M��1��%��Z���k�u�$oi HP��M���˵# ����Ө��e�U��y:��՞�zIv�h
]�m���)n�y�M0qdcR;��v��R^K:��F���I( ��n�{ ��gq����vH�`գ��75%�����m�Vp� O6x�ƭ�)�ag�m�Ŷ�Q�P[g�=�+ɛm=@=.҄ls[Hvinı�0�Y��� \��Am�!+J:Hry�6&��
��Xa�s�Aнi�V�*-���g !����Tr�c���N�l�ŗZ2&�rJ�1�j�����:�:E���F��m�ӝ���gpU7a-�.71����s�hb��v�<ҠJgRr�0]\��J��<[��y�r���3rtV��]�0�je^�Mv�v��Z5J�6�*�gs����kg�@���V�fܤ��@��VZ	�R�A;Ohs�	��Uq�b��R��ތpSH�8[��M�X���ʫ�L��)ŕ�֥Zz� �:���K�kƥՄ�c	����� �p�����#;h���{����]�XN���tC�P�EQ�͈�����*`��ww~��ߝ?����ݶ  *��	���o@��۲q2��:!'��#���Qң����u�$4]��C�AU�=K�Fbt@f�$�)<�*�Z���&ݝ�L��Ud�n�M�U�n+.�Ep=u]�9���q�u�t&
w��O�Ms&�[��%ITx�qJ����,W[�����nma"NS1�Ƒ.�j�A퉖r���Yţ�����wn�wz��~��qˎ�]�\�GE���i��ete�7	uٺZM��W�qK6�uN�7�Y��Y�ַ��)=���y)J_{��R����쟒�R��?w���U U��{d�m�X]��nr��T��]����JR���]�����߻�)JRwﻵ�ʤ9)w��ٙkYZ5�Z�]�9T��-��p�AT�y�|��);����R������)>;���XD�R��.AW
�K���ʥJRwﻵ�)}�{�)JRw�뢮H*��,0���n�.��T�JN��v���/��w�)JN��vJR��~)K�~�f9[���[ܽ:���՞ɂ�hm�4=���]t5.�W���=��u$�"끺�����������w�)JN��vJR��~��*��AKs6Up�AT�y����m�Gf�j�o|R����a�z���B��w��R�����y)J�d�R
�
�#��e�"d�"��JR��~)I߾�ג�������)I�{���JR����kf���f�Y�f��)JRwﻵ�)}�{�)JRw���R��;�u�)HU��@cNX]���ʯ�R
�g�w�)JN��vJR��~)J�{%W
�H��VբYl���v�\�X�x�bҕ�^���	�8�p6�O:�9���l��3[��);�u�y)J{���┥'~������,���R
��n��oKQ4Էw�O%)Os�w\��'���ג��߿~��);�u�y)J}�w���l�e��>U �AK=�\*�R_{��S�� d@jN��vUH*�o=��H*�R�Vc��ݻl���ݼ�ג�������)I�{���JS�����?��~�my)J�za�.�Wq4�$�R
����%)O��)I߾�ג���̜�AT��z�eڸ�\����눘�y5���D��GlJu���[��U�v3�:�^��K�D�.Ev7 ��R
����ʤ
Rwﻵ�)}��|R����b�U �G�|'��)�q��T��,��UpZRVU#7vr�R
[�{%)O��)C�~�w-�h��5�����JR�~��)JRw���C�2S����qJR��{�k�JP���44▭�䜪AU���+(���~����s���┥'~��^JPqW�AW�g��������7�)JO~՚��f7��ݛ�<��>���┥'~��^JR���w�)JN��vJR�����p��囵����J4���r��Y�wj�i9��{a�tK��҃��ĵ?{ݷ��{�?���y)J_w���);�u�y)J}y��T��.�f;��۶�E��-�y)J_w�� ����'�k�<��@�N��ߵ�)JO���%"�v��.�Wq4�$�R
�����R��;��R�����y)UH�fNU �@��=~f\�&Ir+���JR�g{�qJR��}ݯ%)O��)I�{���JR����kf���f�Y�f��)JRwﻵ��{�߿k�R�������R��;��R���������k{��3{�� ����d�k�:K��ٺ�]t������l���CpVN�����b�u�扉/#v�n�M���G-=��"$�L�ڶZxet1�5 L�X��:����t�rv�Q�,Rf7l�V�Np4�+j�ks&�%l����^F�\��rl�ӧ��J����Z�֓�C�m�/)m9J��ɐ�|/V�t�t����Ҫ<
v���yt1��t<ΛW]��+s*,ڤ�M��OSU�����ۜ��U �Y���R
�w���R��;���!.JR~�m�H*���j�ӊZ�n9ʤH���]�������\R����wk�JS���⟑�R��j�f�ٺ�F�Y��{����s���┥'~��^HB����b=����c�5�2,-f���~X?I�����)�߿s�R�����<��>���┥'���z�fk4ke�ٻy��%)O���R�~���~��JS����qJR��}ݯ
�K�~/Wh�₈��n��\�.-�z륉�e��Iv:טW�Q+*S�ū6i��|R����a�)�w���);����o%)O����R���fܒ&Ir+�p�AT�����H�z�f�rR����^JR�}�w�)JN��vI��`�R�g�QF�ۈ���ʤH)}������߻��JR���]����sُ�H*�*��l�"c�o�ۜ��)_�	�߿���)JO�~��y)Jw>�u�)JN��v���.���XƆ�Rձ�'*�U ��ǂ�H��}��R�����y)J]���
��*�Kٓn�6��.1�ȭ�m�Hv,v�g����t��7��)����8v�j&����r
�H*��n�U �);����R���{�)JRw���AT���v�,i�wm�#�R
�I߾�ב�@	��w���JR���諅R
����ʥ���R����ݻl���	nUp�AT���ʤH(��a䇢 �B@$�!�r����┥'}��^JR��o�퐻m\e��q�ʤH)gqૅR�;�w�┥'~��^JR�~�w�AT�W�f\�&Ir+�p�@�s��\R����wk�JR�����)I�{���JS���fk#F]*�R����ۃ,��-�%��8�mN��J��������Q�v�.;q�R
Y�wk�JR�����)I�{���JU���ʤH~��R!�9av�v��JR��߷�iJN��vJR�ϻ�qJR��}ݯ%)K��]#Z3F�oխ�{┥'}�%)N��)I߾�ג��߻��JT���ۗlj[��AW
�K/��\R����wk�JR�����	��Q"QC�N��vJR�u{.�%�0��n8�T��,��UrR��Bs�~��)?}�_��U,�f>U �AK�̸��w�lI�9(N���]l�Cv��i&B�-����nuE�\�"m�n�ݴ�-�	nUp�AT��d�%)I�{���JS��{�)JRw�d��T��v�񑐻m\e��q�ʢ����a�)�����);����R���{�)JP����������p����W
�K/ُ�H*�R�{"�R���{�)JRw���R��w�"�4��E�n>U �AK=��R���{�)JRw���R��*H�כ��H*�*��;�"c�o�Y��|��/���|R����a�)�����);����R��P<��;׽���~t��[Fv�� 6�ݧ8�}*K=$����Z�p.���zVyG�@��RG6�61u;��ȓ�� ���v�=nd�x���&��z���D�eB��4��b�$�#6h�H����J�I�vUf[�C�6r8�m۝'m�{,�F�c�[���\���1V%'�����dU�Vm�;[��U3������ty��oi����DF`����������_`<sXٷeR!s�5۴��n����c����WCP�7�8�Mp�٣]����ᚵ��~�JRw��y)Jw>�u�)JN��v���.���R�{}��ۂ`��MF�4
�k���s@/m���h�ړ؇�#Sێ�����M������d�2����Ŏ`��D�h�@��M������3�����<nr�2\l�`Mۃ �%�6���C�Q��&y���\�ֈ뇞����[��.����gQ�D�:F��wc-��	�p`d��p`��xHӻp��|=�:��iK)v�U+�9�� �za�2������r<c�~i� z��@���]����;h\@��A`�wv�̗['���&�l	�b�m��4Էq܇ ��c�U%�{||��M����j���I���9��6��U�m�^�L��feɤ�k�{v�'O�b�9�j`�q��留 ��h���<�����浴����
C@/m�9e4
�k�g�����Ɓ��+�PM�#Ǎ�&��]��]ϻ�r�q��|�0�+"Q9$�G_tx��b$�i}5�/������6AB�6b��o�'�Ԛ=5��R@�{��!ѱ>�GX�D&�\҄���A#,U`8&3k��C�
6&��<7��	%�#���	�&�`��<VbC���v�����UH��YDC�l^�RuT��w�� ?{�8�f+�D��%�����J������8��h����:$x�pq����&�l�p`E�q��͈�	ɷ��Z��u�B��4�]�f��$��[��m����˾�켳�?�� ��߭��.	��03%����f"��ӊ�9$��L9�UT�ٵ��@�}<h�@����J!�Ț�Hh�ՠs�S@/m�9e4��I�M#S܎-���߻��}��r�$tM&�W�F�Lҿ��>�B��i��9 �4�٠s�S@�v������m�=]x��j��1]��R�J��=�ѵ��v���R��p�P@�i���}����%4�j�9�)��� ���rc#p�ƣ��z�Z9e4�٠s�S}��t<?�4���@���`d�d�0"�9ﺀ�Np�"M�]�����>߾� �s' �fqp>T����8^�j#�i�C9wv�3$��03%��M�����-�bCB�s����z�o� �  ����K�E�u�uRp]U�l��Ҋ�k9�6���f�	����-΍F�)��[5#��u��pm�;r�Z3�M���:Ϧ�a�gk���۵�m��i��'�K�Zܯ^Cp��W��uV�:�-�5�h�ٞ�cf�J���ZW�Xe�f*�˕�q:n�Ie��"R�V�/Z���f�ga�ow�wwwoH||��\f��tSѰګL�#d�����<�f���)�m��CǑ4�rt�n��YM ��{�g��ޚ�|���L#Q�s��t�̗6K`�[l���
ֶ�9�rAHh�@9˓�����U$�����{f��쵒Z�6��Sqɠ�@��s@�,��^�4�ˊ91��r)&�6GL�p`d��%�1E�#Ýӑ�u�tn�����^7P�:�n���+<Kְ��[dL���nt��̗6K`�_�ꮠ���0��z��q������77g)	%Tm9�@6�[,:�P3���;6:`fK�T�)+��Պ���`�[l�����&�4��R"!�Țr94?�~���}��w��M��d����.;�Ǌ(�����9�)��� �-�����/�	 &��6��]k����C�h{k]l�%�v�&
��ۮմ��9�rAHh�@9�f�{n��YM��e�(�k�1��̒�dt�̗6K`��)_$�F�JB)&�{n��YM7ߌ#I6_�' =�d�t0xH4ڙ1AI�9e4�٠�@��s@/R��7��	?�=��_z0?-�z���遙.!�R�*�s�����:���k���ʆ�7AqDìR�"Y�Nʑ�7M��zi��$�����&�遙.l���%��Z"<���rh��h���f�s���'���BF�n'3@�-��M��d���#�d	��Ę���
C@/m��[4�w4�^ 8�̈0#D�_��۴P�d�9�o�*�=���7���1Lm�&�s��������{l�9�ҥ�2f�����<v��2�k#q����5�:殛�s�-�k�6�$"�h��h���f�s�� �
<�2A�jd�&h�`d��%�&����}���R�6��_��p���������\��S@�.x<s �c�M �-��9e4�٠\�	��h�]�&�遙.l��33' �WUT�8��RF+�o$����@ حe�jŷ�Tr��>���y�ٕ)ׯ4�$y�(�:ڈ��IS��;�خ��8��f�5A�Y.�ٲ�A�(\���v4f�I�2,ѭ��7�����͛�j�v9՜Ͱ�N�)�:�}YY��teٺ�n+���+��ˠ��R��.�Ԣ��-�b�t�����A��ݜ���,�N�y�����x�;7�9A(�{ݛ�j5��mj�تy黣�E���4�eq��i��΁�즀^�4��h��h�
ֶ&�9�rAHh�@3$��03%���b�v��s��#qɠ�@����9�)���@>�e���܉9�I4?�~��){o�L�_�7e��-�L5W2������Šs�S@/{f�s���g^e�UT�{�۶�ִ2�n.��Cq�+��Ւ���,�&]W��Ì�n0��6�,���s�:��Ӏv�k�/�@�,���z��A�k{�*�=�u��I(A (��H$)�GV{��9W�}��{�4K՘�<yJD��.rD�̗~��#�z����el�m��4ӑ���YM ��sԕR��I��;�w��wi�[�b�ݖ�Œq�3�&d�0=�33�-����L��E ���H��`y�gn"&"���!�5�0K��˜� ��#6����y��ՠs�S����h<y�����"��#�/9"`fK� ����N0	���J��xڙ1IZ9e4��i��}���
��)�8+�-w;�=��V�r���0m�!$��7O�䒥w��Ӏz���u�_ �ra�;_UM(Lhr7$�8�k�=���g�w��4��h��%���3.�9m��vL,� �b�[��a1OK�^�%����cjLY1�ȚR'�yn��YM ��-z�v�lDhnIn.��ÛT���s6p_�_ ��qsi*�v{��ӈ�$.C�e��,���:`fK���\�V$�)�1`ۏ@��@�s@�,��� ' t&��_�M~�k�_t�=�91��E#JG�v۹�s�S@궽�����bI���X`�0�U�ѷ`x�ц����,��iם�R�E� �<�2A�jd�"s4r�hY��o��j�_�3wx����Clr˻��p��UK_�|�������������ߒ;�W�J����|����=��\>T���{f�/w_ ��M:,x��M)�@�s@�.qp^f>ԯ�ۯ�f���7dhm��h廚U��\����ʶc$"x�`A�v�y������A�I��R`!�GI�S�A����E�1c``i v�D0@��I2�b�$`d�aɍ�KG� heiء�P��<�):�QHPx�f{�8"���tB���t�� �q=	1��'��HsK��/�>yㆴ�H�ٽ�F��y�Ou�����{�����������H     [F�      %�          $ �g[!R��J���Gf� �*�(\acn�Y���T���v��ێ��i#L�<��5�U��� ��(�
(�u3���6��PM�)YSa�R��f:\�rW; dS�5�n�6��#�ٝ�.K��%b�cSUkm�S�������$��I��q�i�N�( ��m���&����j6sg9%�-�3HF���ܚ8�[��rN��gҠ��.L�@G	WD�FH8,��0C�C��G�).��u�:���>D���Q�9�s͵Yv\�-�`�F�!L�vηy(�����P�wu��p�4!�ty�4�`J��mTL��AV@iA	E"j����a7泝Z5 ���;7L�Jָ��E�t�&�MR�p�&ע���R�[NRY�>K�#�A��z�z�T	!6*�v���͒�]��{R��Ӻ/R�k��6�)%���D��J�;�C������҄�5�F_S�T�̜�����]O����Djz�g9�g�\\�i�R)`V��x���)ېİ
Q[m�t�6���n3"We	�!5p�lݝ��[#�j��HC���s��� �PNH�r�n%���*�ݪVvYWm�C���\l�X����m�6�eZx�k�B�V���I·C��x��wm.�r�-� iJƦ�Th3盭�����v�Fs3�՝!�ZMe6j�)���,l���>�����W�m�,�#��EH���!�EԇR��F���F����R���u0�i@S7dIV�R�2��ZWp�2dkaVu �JԸ5�YL�d���׎�`L�m��Mn���K �M�q�S۝�n�I��+��%�as�nZ�cz��u����2lGDKS����:�ђ�I�6)h	v�!�>Ӭ�s�j�fjֵ���{�U�z�]��v�(����w��⏿ (���`	�"y��Vж�� k�䷐8\m��Yn�(-�ٜKЎ�1:�Tۘ�*�I��ݍr���y�Zܺglun�乎3h*�,��ce�m�(�U�li��Wm�Rp8�56���A�3	���Yշ"��P,.#�uqW,�N��:�>k;���)p��h�;�b:��r�̓��l����#��.y�î����G���%�t�l�{��{��M����r�'3�a^&9I��7j��⩧#G�s���8���sv������'d������7}�LU�./(4�)�1`ۏ@9�f���Z9e4�j�~��/3أ��N5$��v�{���ꪻ�{��{vp��Ǘ&H<mL���-���k�| �s'UUR����v���5H��.��9��{���J�����׻|�ɇ �K7w�wui�"[R�m5eN��v��/Z�Ŵ�7)��\�C�އ>�.���}���҄Ƈ �x7 -���k�h�L>�_�2�u��anޖ�����-��=�2��K�I% ����2����[4�R{ ����nE�s�S@궽 �-�k�h�
ֶ�&$䂐�:��@9�f���Z9e4�Z��7�c�X6���2p��f�����N����1u��]bGS�����NH�l7=j#�űI;I����k�l����k�-���큳�&d�����P�����d�S&)��s��hVנ�@�s@9z���BI�9��{����NJRUB�R�U\��U%�y�8��fqp���wp��r��ܾ�R�w�͜7w��{��\�ڴK۩0x�&��ɠv�遙#��'d��̊��D��Ջ�Dͤ�EƪG�^�L�C�&-��g�:j�cv�h��n:�I�������01n�0�-�ݗd	��ęl���qp߽��T��{vp种��s@�)XX�o��m��3$�v\�:`bݜ`��qI&2GmI4�e4r���������I�D޾�;�Uy�����S&"G3@�-��8�����hv����jX	��6F��\KS�s�/k%�k�э8ջV�)0i.�qf���c�6���I��*����r���۹�w��h㮦�&<NAd@�| �{'?���n�p�� �����vn�U���MKwn7' �n�pr�����@9{f��jOcY	���nE�=��.��������_/�Ɓ{�<����ȓ�	��8����e�;���ܑ�~��[[WfW.@ ֝y5�q���:�CI�kw�n��P��n���uV�]����+��z.�i�۪���Ӵ�ٵ��.�er�c�i��I�we�2�ZS�h�ع�'����;��o��a�h��q�9�mu]��s��M�7N��M �ٺ��`v�ʨ-/C�Y�B�jHÁιq�unz���M��m�ﻻ��}���N]�p���c�+��*��ҫv�n+ƀ*^c�LCa"i�Sb�� //���l���[��qw��Ԭ���#��r�v���遹#�-���e��J���3L�֨�v7qEd�.��t�Ż8�2l�vGLf�%]��	����o��r�������s@�}u4�CC�X�7�r��07$t��$���W�����˗9�y�y�)���t��Ub�2]y�$ӻS�݊�gn��<+��B��'��L�05I9﫨���'��o������㋀{��\���QI<�0L@��Wb\���u��������J����ȓ�.]05I8�2l�z�����t���:�8��yTi7�21�ۏ@9{f����h廚����V\�I���-]�큻��rGL�'M�@�ꪥ��fF6� �Ǌa�ȟ	E�0�=�kf�+vn�I�IzH�����Rg���X�遹#�T��&�`n���ް��BDH�����/{�@9�f����h廚�X�R!�r��q��̜��qp�i'J�J�|�/�H
8�o>���*����-k�Nb`�D�q94��i��#�T��2K`l�s��R�L�m�&h廚�����h�n�e�jK��H4�0La0�7Z����0�c�9���hj]��OU�����t�A�'Nf�� �-�{۹�s��hYN��4���mǠ���H�]X�:`����RA�N�ܘ�$"�ɠ[}��w��h+k�^٠�\yrd�����w���*�;��^����@�� ���߳3"�~� ����$d�	�
M�����M����遹#����x����o��҄��!��j�ё�T5z����U�9�xj��g��&�?����=�g �s8��J�Xv�u�w�?c��LȚqI4��s@�-��>Vנ��@�7�,�����Wt�ܑ��I��e�7v:`w�L��ؚL�8�s4=�����`n�t�ܑ�Cyb\T��c���r�����yn��{w�O������������m�7m�H  7Fѥ�bۉ�-e74x��q-�j%�Vq���r
Yꑼ���p$�Y�#�+seᴉ����"&0Wl�hh��)zWeJ���#��F]'7n�3@Nn��t4N����]-/c���I<��S�h�ӓC�GE.����2��iR�itu��#�uH��fӊ�H5�
��e��H�ng �A�c�Tv�G7����NoY���5V��g�W,0�+��L�`�^��7l\�lL����"y1����x�;�up�{�%����� b�Z���ں�ZWt�ܑ��I��e�7vqsj�*Wa��5H�#$�-�\�_�����0�-���䤞t���:`M�.6�1��,h�@9{f����h廚����}�qI��yN)#wc�䎘RN0�-�vH�Ә¥��q���۵�[�{���.��T��wi9�յ��F�u��+�lnH��$� ɲ��07*8�n��ێ.��1�J��K)*��$�� ��N���.��qsU]�Y�
	5�26���w��@�{w4����mz�R��rL���]�.�z��$�i�7�t��q�d�4�zc˓$hmL��I�yn���1�����qp�����i֛�'m�v�����K�Oc�u�,s��Nr.���^�nf�{f��A�l������'��?��&�`n�t�ܑ�o$��+.��Ac@�z��4��s@�-��>Vנ^`>㸜�4�h�n���{������x#�қج�J	��>���H@L�X�Bb�0`L�`�$I#)2�����֑Y����b@̅J�b�3��h�3�C+�+�4q��Z<���$��4 I"Y�jHa`�J@��f`�e	X!` h�d�9��,�
Z88�V�H@��[����&��+
	f����
�
Bb�(��@��? >]p��6��t��)��	��(��1Q��@)�{����� =�d�Ԫ����o�]Z�Q�ۗ"`M��0;9"`6[wc��Љ�ؚL�8�s4��h/l�;�����s@�;o���A��%�駭s�N\M��]�:ゑ�3Ƶ�3Lʣz�.
	5�26�7�r������;�w4��h}Jˑ�2<sqݰ7%���#�NlL&�`S�<�2F��Ȉ���w��h�ՠ�d��g6�%J�3q�d��'#������:�$��O�� {sg �{8�$�/R���g��;ܙ#q�r\G-0�-��c�䎘��=����~Û�����g/\y�aУF�u��Ɇz��� ��v�v���a���嫻`d�遹#��$L&�`{3.�"ujGcq܋�{��\�I$���ݾ {sg �{8���Uٞ�6����dI���^�yh���/,���[��ugJ�4�(���zM�06H遹#��'v���	9�C@�즁�[��Uˏ�w�0��]�iUڈTU<2~m�-�p ��<�Z�qm<#�8㑼��*c�a�P��Ͱb��E5�z�T.�%ת"E�'f덳pJ��&pm�`[��z:U�v�� �C��67mY�JМnϖ�sGPVX^R�9�Uܼ�j�eZ�lɯ���M��ۊQ�]�E��g=h�#�E*���k�Rj��B�fr[\s���q"�m����(���<? ������I�]v��pF.n[�-㥷9���WWL��B?L�Ǔ&H�ڙ�!�>ｹ�U�^��YM�����TI���璻u�<��� ̒�$t�̑��,�7�X�)�s��d���:`j�q�2��\��b�%#�#���^n���=��.����r٠}mI���d&F��Rf��Z遪I��%�6H遛"|�A|cs��]��b[b�	��v�96����m�s�J���V��Ă��n�m�??? ;���3ޘj�UJ�X{ۼ\-ik��ը�݃� ;��̪��J���ܲ���0"�8�0�NW˓!#ɉ���/{)�w��i���w��h}s�@.^����S"$4�02sb`6��7%��nN*�I�F����s�;�|���f��YM��s����$�Hǐ�1�5<���]��y1z�����x�F��oXCD��d��<ri8����w�S@�-��9_j�/0q�O"`�F��.����ܑ�'6&�	l�Qvc���hm�@�-��/_j���Q�����w��o�w�ە}�Ҧ-i4�q��h��h9K4�)�w��hYE�ԓx�21�O��d%�7%���#�NlL	_�����[<��Wj�z�)�p79nz�km���I]�O]���5���9μ�e�r\�:`E�q�fB[ �/Lyrd����yn�W-z�R���� �+U�$�������{���ᓇ�Uw����/}����Ɣ ��,h�@9�K`l��rGL;�UUw�m��0;���'�0y#NFI�v۹�w��hVנ�,�;�׭��<k�K$3���N��ćk��q����V����i�u��J�1d'���jL�;�w4�k�r�h��h����&�8)n遪I��	l	�p`nH遪��:�oFF<��9K4��pګ��� ����Nጊ9"��].Z��7n�0"�8�3!&�}N�yfH��ɑ�yn恩k����i��g�0��꒪E$>���0,�˻�fo{�fo{��l ��'_ؗ���:9'Y�-��+@���nh��l1R!�[o��%z9+O;!V�#;=��j��'l���s{k��l���'�]B��E�:���v�mL9����u��7C���ݑ�OO:#l�kf�^z�c��\��꧍�f���ִ�m���<�4��G-�V�3�3��FeT8#��^��.�kr���I�#je��:=�����o��q�g� ��v��Z��t��R��4���&�I�%�H,Xm��c����H����˹8������?ʪ�W�i���4ڪK��{w��yfM���r�����ᓚ����̚p�� ��c�*UWe�����l�ۑ�p	�p`nH�I��	l	��!?F���4����Z����ײ�y��ikM��73@՛8�3!-��#�䎘S�]�ټ�f�5p�����i�r��{6�:�N��H:��ы�bx�Ӟ�O�m�	l�07$t��6q�a��-\�&H�V��N�{8��}B^���Uޜs01l�`���;UʗW|Ck&LA$���s@�vנ�,�9��� �+UAE�I��W��IfB_z�Y���I~����ew�$W�=#q�9����Is���K���4�[�v�Ԓ�l|I/U}_s|yy��ܦӮn�v�͙㮢�]<Q�f��$3'�Ήۣϡ�����#N�Ē��:M$�䝮�$����q$�G��W�ɱ�!247�I�RIs��m$������]��ޤ�o#��InU�,J4�8)Ng�$�n�RI.r�~y���HVT!FF<L����-I%�-�>�$��VŢMb���W|I%�	}�If�:M$�䝮�$�ۺ�Ip�+&)$�H�bqBO�I,�GI����UT�{+1$�y�i$�r�}�Iu�UK�c21�?�� ���7�S�cQ�GL�:gI��lj��S�m��n8��]] ��M$�䝮�$�c`�I.r�}�Is��-I$���rH��q!��]��I-�lI%�	}�If�:M$�yo���$e��ڄ9�
8�IfB_z�Y���I%�'k�I,��4�W���\D��9'�$�:��Ԓ[�v�Ԓ͸��W��}U\�ꪟU4�t��Jۓ[bBdhmH�ǩ$��;]�Il���I,�K�RKT���I.���~�v������ \F�c��ba��N}k��m��ۦ�q��u��<kkf�n�]w�%�6$�̄��$�H럪������}��K��y��I���$��I,�K�RKT���InI��RKdl5$���VL��d�ɍ�	>�$��uƒKrN�z�[#`�I,�K�RI*�1�#Ck&D9�RIw���|�W�q&�IfB_z�QluƒInN"Uݥ#HO�Rns�%�'�ԒK���|�����ffg���y���ݣ�+G�#@0���ř��lۂ22BJ�3��f3�`���G�Q��}���3:�k�5�,,���4�И����Y	��g���Y{����t�I�<:uL�#�+�B3x��X<@w����b�/�#�^+�eV^�z���Bc�#����@"4�`�� �_$@~9��!{�=�绷{޻���     u��դ�    %�          $ 	9����)R��]�<�R�7Ù�#S�Q2n�6�n�����[���M[	�.������$�][ƦUV@Vv����h
]�6l��^m��Uط]�S�Sckn�&�m���%�������]yx��6z̪	�:ڊ!�ʵ�����\,l�Fw �����]8�K�ֶ�@ɕmZu;P�c��L�j��m��<q&��iȶv�Xn<�8�oj��\i���saX�<vV������(�ik.�ݺ�(N�u���|�|�p��<q�X0dx�N�۬��#J,\z�[��-���h�Q�28��G����}�cf���s��t��J��n�ӚGJ�����6m*e��e��"ʪ�]-(
�Fl�+(�.Dv���V��-���u�-����Hv�4���9��`�u5غGhU�i
vZ��ܻ�ZwXu����+��W�6�]X-��nv�;
�*0�����E���Etq��j�j�j#����PU�S��+-�X�9s� f#m��1Vٰ�д��m+[m��܁��� :
C��b��Wa7���[�G%�ݶ4��L���REx�6��+J1R�+�	�UD�(d
��)vC%*��U[&#j��n���U��e0�z�V2l���Ok�C�zV�\e��A�S�#s_Gn2�L��IFEkuDt4�mq�t(ngM��:�:@
�����7Ny���+d�\	�0��O�]t��#1��u�T�+=m�D9Ͷ��8+�� tv73X$��g%����D��t�p�d�kp�\Ds��90�R��UR��`�sj��ebؙ��M�@�[}4�x�J���l�$QB�F�v�)`��ZpeKun�ƤB`X � ô�����ʻCMa�W(�fGa�+[Jg�v��k[ٲ�j�[�@<@�j�<OE��ȧ�C������ b�q��F���[?�W.m  :ӃnD��=��b7ݾ�yR]�"[���� x�%ᒈ�����}n�zmۍ�Nu�lf���wӻV�a����t���z	뀶�uŻ`�U��S��[���2S8���v�b�o+�F% �J)�A��F����Hsd�g���&2T���Gmͱn��i(4���i�2�+<�C���{��|����˿T�Y	q6C��z��k��m���*��DF��@�W;�j���k�h?`�����I(�:�I%�'k�I)�q&�Jg軅�Ș<��#$�䒫�q�I.�߳�J�J���\�,�����������#CjD�=I%{�}�|�W�T�$��)g�$�]��RIw�
Lx�����%{%KRI.r�}�IU۸�$�yo���%�L���&�FF<��4�K2�Ԓ3n�InI��RK6��� ��/�?��F5���r��f^�:�c�+t��+�h�׭r�^.Z�t�y�&7$��9�I�$��~ϾI.v]F��\�,��K9�Y�46�a2L���33>����Ω��C�O$M �h�0��0<�Y���̹��������]ݝ��sU%UI�wy�vj��$9i��v�1$���CI$�!/�I#6�5$�yo���%��~�}#jx�$�-Iw���_z�F��m$�䝮�$���5$��軅cDhy#NFI��$f�-��#�n�L2��q%��u�$�N�Z���ls��'=n�vnZ��n��=][���\&��eQ��ے:`wv��3!/�_}��@d����6Ӹ1�n9n.�ޘsn���f�r�M��s}��"�g�KRM ��i��������8jX�Z��}��4v�Ö�c��$��l����:`w6��3!-����5�H�n�DR\��{��\ UJ�}κh9K4�v���[m�FVm��cZ[���pqR�!����{k����uؽ�Z�G��$	$$HO�Nn|;g�܄���l͎�ۛ9|��Y���B.�܄�ܒ��09�����]
Ĉ��F���@>����遙�� �B[��N�����v6ݹ8R��f�\���������P؁
� q9�{��y񪪄lcdI��h�n�}�Y�r٠w���oj��X���I�1�i�\��\�N4�����<�!�5�0��v7P��Q$�,��l�f�}�Y�s�h�n��;)���o&&s���`͖�Ig�03e�`�I�U�Ώ,�!�0�"rh�n��ۃ �B[ �l��8�WawvH����6|;g� ���@>�l��h�w��I�x��'!�r�p�}���p��À~i"��K�����c�� a�ã:���.v*v�p��e�����V��X�\�.��3��Ƥ�A\��U��NѶß6%=ur�9�`�ؕscR��ePz���,=�J�J�ͷV������r��a�2�t��ekŧP�<,=s�ON�8:n�d���<�X���ب]�-U�7�|r[9n0�.#[\2�9{�������8��ڽz����sy�t(ڱ�a�����1OC�^��e+�����rm&z��W�m�߭�nl�͎�r�)�8pymI4���즀}�Y�s�o�~�H����cdI��l�~r�se�͖���+ijI����C@>�,���8�{'iURJ��� 雬���$���ℚ�;f�w��@�����if��]�!���5�b�t�6퇣j4%���5v�����.n�'r�7���WQ�S	�'&�w��@�����if�}�٠�j�@�BD��5)��3g�:*�}��6�l�����`���I�x���@>�,���8}J��f� wٳ�g�߃w-�R5˾l�����`͖�;��������c����jI��l�=����f�_@3|z�se�7dO�T����9k-��kX8vZkNt�A��d���t-�L�"J\j���elT�_m��6[ �B[ �l���O�U}�|�6��Ԙ�F�Q��wǦ�}�٠w�������>\-Dƣ�G�ɍ˄� ��d���Iy5HJ�HH^1�-1x��H�%Ts���\ �x��2�W��)�����\�`�-����w!-�����M ��^D�$���jSg�s�ی�	l�����`E�	/��鵮$���t��I��X.i�����zËM�H�1�<sKs4�R� �l����}_}��Θ���4D��I�}�پH/o����nh.R���rV��A�hm�$�͖��lt���N0��`nW		qۻi��[��������ˀv���^{�w��@?,L�+
��Uj�eRT�ҹ�7��74�m�.��F�Q��>\�z�;f�w��@���.�Փ6���P"lP�+���˺:[*;WM� ��9fM���n5��;dY�rG�������M �;f��;w4�)^�Vs:<�$x��ȉ�@76[��� �B[ �l��S�� I!"G�i�g�s�ۚ�v� ���@/-���lcnx��&�0��`͖�&Il?W�_}T�l��=%�h���mM ���@ԕ^�v~ �g ;��p/�n�eR�ݽ�g���m��  m��]tW�����H�δ��r$8V��L�[-Vv;k�E�,[�z��ٱWcAfw���-��l�QB�����ѝ�X#��D+&�<�h��#j�ⶩ�'��<�VM���:�%�˴�P+,;�9��ds^�N��aac�62t�]�\kX�qr(9�S�,΃R9�kn�C��#�u�ge�ݮ�T*5���A߮�{��������I\.�Z��l��f���ۺ:�ƽKRR5��z�V�q��^e�Mg�ʥ������;�-�d6_���`{���FƓ�$q94�v� �;f�}�٠����F�Ա"���]� ʛ-�w6[ ܒ�se�>\)rcQ�#����rM ���@;�f�}�٠��4
��1�#�6����9v�7$���l*l���4���,X�x�<S8�B,M�:{W.��NU��նJLq-���o�����MumU�i���ހO~�v�6�sy`�{49���i��(9&�s/l��*�/�T���f� ~�����'?Į�_ŉ{�cǒ4�)&�s��@;�f�}�٠��4���^60�����+�`�[ �l��6[}�Ԗm��/r�OS�'��9NM ���@��k�����`�[ �͉/�U���f�#��-E�`���'b��]*�j�v��&�y�?m��A��j9�̽�@?w2p�̛J�����f��񦨝ǌ��1�4�v� �-�����e�YΘ�̑�S&)�B����*�߻×�qCh'p��M1#$m��7����JВ��G	'6�����}3E�� �b�	 A x�I,�$�ăH�3��2�,�
����l�&JXFcm���<O5�����}a�^!��[Qןxm�E�P$�` �  <� >�rD�@~�s\1M��C��i� dN��|����x*'��G�*� |�}a�?��0�����o�L�� ;�M ��?�RAď��fπ�<�eM��;6[�}�}IM���Z��1��cs4�{f�}{f�w�������Ux���cH�λBLU�m
�+;X8q\F捧I,�ø���"�()��X�<���I4��4�̜��qm*I%������:�֛A�hm�$��٠w���̽�@>��@�3�^��O�r8����L*l�ٲ������Z�A�ڑ��̽�@>����+�~��W�� �8 ������tB6#�Бw��������Lj<dx<�َI�^٠�@�;w4�{f�ε�R����'��5�l�:Rgd�L�ֹ-�'BI��[��!�r�۲c�2G�mH
G$��٠w���̽��33>@s��@/h�"B)28��8rr~=��ϕU*�������l�yl��tec��0Ę�� �M��;6[ ܒ��0%mb�������i�8�]�sg 3۳�{���̽�@�/rW�� �46ڒ0�-���� ʛ-�vl��k��=�w~r_���x�  �]iie����Y��\b�N�^t"��i.��(�nmɦ��uj�$�I��l� �v��n̸�4��_F*���$p�e��C�\n���`�|�I�jv��O^] b�n�]ƘD�K����luwbu�3X[���4ζ⮍�\"���.j5<�〷�4��G�y#\�p�K�����{�{w{������߯�ߠ;���]YSb�nɈ�lq��:z�̜��\��U�-��e�����C ��INO�����s@9��h׶hyl�;Δm�I� �mH�� �^�`�-�nIl͎�����Hŧ�dƣ�G�ɍ���_M �-�y۹���4>�\�#����lrK`flt�2��`�-�w��Г	&9?�M�>����e��-��[4V����Y�$5�k@�"����q�7-�=]2��TK�k�.u3���$O�cs> �z�hܒ������+h�\�|�K�y�a��|����|�t%�������I���o�����4��%x��#Cm�&�w������e��-�y�*z�1?�	��rh9�T�l�%��-�������a��&0�Q�#s> �z�hܶh��8{����T���/��W�d�|����s�Ճl5������L	N��h�[p��Y2cQ�#����rO�9�zhyl�9��� �^٠�2�����
�]� ܒ��0���rY�f~��_Lt$�I�F���fπ�{��*�;�w�I�o����$�W��ݜ �n� .�͘Ƥ��B�Ü�`Se���7$�f�L�ƻ�MD��yk�@>�@�eUR��_@ݞt�2��`lۉ*�W�qs�
K-n8۰덫�:^��@�ܴ˵]��] �s91��F�ێM �-�f�L*l�ܒ���\k�ğ�$q94s�s@9��hܶhyl�9Δlz&0�Q�#s4�6[ �IlrK`flt��ȪU�x��y1��@>�@;�f�s�������s��Q�ZZ��3W�N -�jؤ�2K�%�f�`~��=} ͯz�rK`z����ο��N�;���u�Vcm�����=�\j�S�&����a�gY�N�S��-�����l�R[ �Il3l��z�ƖH�9�%"�h��f�w$����f�����=R��xpoo"n<�h;�M �;f�H�o��s��M�;��la����C�}U�|������`ʒ�rK`s�J���'��INM �;f�}̲�rK`�-�>�_UW�*u%�w|�	  �.I��m2����sI�HLq����J�/���vmO��:Ws�-�f�@�k�̗=J�:�O5��������µ��mA/I�Un�uR���=m�t��g��t=Z��x�#^��\��e��V�K$Wn����y�����%��Q\��r˘�4�>���M&�N��M��[[P��)ۗI�����Zַ�2��E�E S�<白k�=[�k4�;����,]L�^.��%۞*C<k^n\�(:�l9�ِ�5�~���rK`�-�fl�VE�&52<Ln,�hܶh9�4���2٠�2匒bR`��ݰ͖�36[ �T��;�[ �)���$�#G��fπ;��s-��-��v� �w��3$O�Wv�;�%���36[ ��|�UR�����m8��(��ݵ�u�ήE*x��:��F�P�7m�ú�.����l�1���&9> �}��l��٠s-�nw%���#Cm�&�s߻�d ��HJ���`��@1VD�Q������������٠s�JޏO�8���c�ܩ-�L��f�`fip�@q��9�W;���@>��@����>Yj:�2LLx8�= �%�͖����VmN06�jGg��v�盖�].���ź"�y�n��O�mt6��6���v�A�e:R��;6[n�LY�8�&Il�)���$�#G�wfπ����:�ܯ@/-�����]���'�a�5��}��w\����x'��BK�z�nh��B�D��yC�W�2K`�-�7c��ڜ`m��u��A�hm����l�/{w8��X��̜�$�}��������m=IGlsh�3:;T��e%�vA���̬PBxƙ6��$q9>��s@��r� ��h׶h�QQ��_8��LY�8�� ��͖�����>Yj:���1����d��;6[2��遫6�HeʦI1)0R)&�}{f�{۹�}��w\��2_�1�E4¢qz���S�L$��h�n�����\��,| ��N ~�d�Ԫ�����v䶚J&u�H]m���y�C�7fnA����;M����k<�H�#�ۃ#w@�e{�d��;6[n�L	��иI��yC�#��f��$���=o�4�w+�;s�hmy|�]�͖����s�Q0	�[딭�m?�
H�rh{�g��}�h�疀^[4��4s(��La�h$s4��*�"��|�\���9W� ��ڨ ���**��*� ��B������
��*�
�� � ����Ȓ( $"�2��("�2*B("��"�0(��4 ���(*���PAW��PAW�UA_ʠ��*�
�"����*�
���*�¨ ��*����*�
��**�**��b��L���Rd�۳ � ���fO� �ܾ     �            ( t  < �I@  (Q� R(E(�@IU�����*�$   *� (� �T  �*�T�L    c  P B� �`P����q�힯3�{;ŕ�q�8������w�o{��-�i�һ�	����o����}�z� K�K��5K�(��_Usj*�k��W�r�{�=�}��uT��+�t�ӗ�^��wJ��� �(P  �h�>���/��>��Zzo}���>����+�>���W��{�Ҿ� �ܟjz������ޚ�&�\} �>��N[ͪrӓ��yp �  ��  ��U^�}=U�5��f����U P  �hg������z\Z�n,��W��ysn�qj�\ۥW����JR� ���   D5�)}`
Q�H�D��� �@@ �  � �� ���  
���C��4Җ2�z1:P4� t{���(0   ٝ(� % рi}\۾�O�ܾ gx��}�����>����Թ�_[����6�^�� =�]��*���eﯽ/���� |>P�I@P 6 �,��nW��qj��jU�>���r�Ū�-}�ܼ�y9:u{ϠI��rk����� ���:��{�S����.-�[��6��{{ǹ��x>��w����m>�׼��{�幽ڛ�OQ56�T� �?�53R�� �<z�U4�)�   D�*�"�L��%6JR�  "$5%)�@G�|	����_���s�����;�����w���^�2�� �*���� �*��@U��V  ������ D��� �*�-H��b%�
_�d�4��č����c�00_ 0��# 0�H�I,����G���H$}}�}��<$��5 P��ܖ�Ӗ4 a�$�#Oa��9�`W�?#�HA��Ń�.%��A|3Җ��}q!V�!!	�`�#�<bTr���0� �!�Xذ1H1�I�N{�Y�ϳɿI������J��H�dX HD��"�H+�@
+
:k��,�
�D�B2d�HD(�,����@��|'C��Hj@+
�$�� H�
B�Qƛ:D��hE b��jD�$FHH�X��`�
����ܔ�|�bY	�E��D)#�x{L����W� F%���`�R\��FLd`�!�7�`��	�G�!L5��,%�e�d�B]��w��6%�#!�H��X�X�l�߽�`ISXE�@�H%B#$T�� $���y�O`�h@ �ۘ�6m�M��	��IM!XX�ͅ��R[͵��I�JRJ%�#hr
�����Vp%	N����\��K���%�픞�
�p��	B%,
���$a��s|�s<�/���}� �X:@�>Y�	�B��$�dDa 4�J��4I(z{�J�B	�"E��"��	~
8C�IeōXĈ%	!�y��xJw�
�d
�k�næ�]�	�<�8� �H	
d66f��q�ε��r�p+��KT[tRe�R����m�)��� J@�)3��l7L�\2SF2f$))�()�c��S;�˙�ww	:w����a�S�	�n}����|x���)�ы �	eԃ`Ń U��!B0H�XL�ߎ����B�$!4���bA�T���H���L� 5X@ P"G �J8a*�#4}p���`�=!XP�C����"L���syp��l�
 FA F!T�� B4�RBI7NHF��L�`R�9�6hG���B���bВ0�q:�Ԫ��'{�BnE�qaB$�dX��턹�(B�$Z�H�L�	9�+�S%f�r��)�W`��Y���7!�1��!XB,$X�ag�j��t��>�*ć�H$ �J1ZI�"����SL��%"S��X!
1�ŀG�!t��x@�jF�����T��a2C�E$�D�bF� B"0w�����O3i�Je��$�5J��@,8JE�e����@�\�5p �4t��S)H0<��RdI{�vL�|� \	_�Ƥ�XW�ǐ�]m�e��L$m[]�"R �ƌ B@�22E�T2cF!��,F��
H��X�"$VHP�%�T���HF�H�I:��@�4�Y�
��Wa��g��D�N#H�� F#@8��p�B��8zp���5s���`�B)"�\d�$�IH��)��$,<��x"�1�i�K))�c�e ]��}O�4-B���Zԑ�w�g�F�HI$(�dB`x�HX�J!�1��2��	�	+Z{32a
��"Tb8Cؔ���	��p�0с ���F4�B1H��d���'��c�ύeܬ܈a
L2�8B�
	a6bVV,�$�CaB!��Ft��S�@�I	�,�d#
���K�%i�F#�f��1j]	����KJ�
��	l�|RŽ�cRV�x��)!e	�).s�y�`F1c�k���&C).�D��,<�r��><�Ù�I8L�ݔ$�Ѝ�+t����H*J��,��d��� I	I�b��dH�e!!`O����r6�/�e�`0"B����I
��@,�$H��4���#F,�T C�e��<�������g��cHP}S�"H��H� GD����D"�b-B��"0��Ӳ�L��u�d����Ysd04d=�A�1!�F R�i@��F@~5�HP�@!A��C/����q!VHЍ_$_)������۾k=w}c��I�y�A�G�
�K�B�!pH98��(B$
,R�	��e3y�y���C~�۳��)�a
�#�B��Fϗ58@���r]�և>��Z��1�A� R&0hC�L���#��B@�1�,"c�Y �l0> �`P�c�#
�+FbF�k�+�K��#
�od�0��K�Fa^��B�)��I$Ha �8B�, �
�B�Ê�I	 ���p�}c�|�),n%~�[�R�çNM{�^Ge�<+d C�HV$�S�
���%�BP�XC�#ƕ$\`X3,�K�X��{�nm�r�L��p�8�
� A�X0>,i�B�`Ň�������no���\�q�ŊW1�F�F2)�t"S1���)���A�O1r70��-�x��HFF�~9I�Bm�~�3��p��Lı�&9���i%'3:M��#5 "$$d��H�`I��F���0�	�$��%H��lԣB�(@�R9
0�!0e�0�5%��%,!8Jo!8M�s9�dHD��$��B�*��l&�K�h`A+J�X� H�$"1hF��
�8�$�.�6O�Oa��������ϼ<X��x�%RD�� W����E�p�4��ďR�s�s���gͪ�S���&�Mݖ�s���w\���h6��''���0.�y|����t�OHG��R]H0��S8H�y��F�'�M!�C~�^Kw>�%����ę����:g4�B�a����h�+�`A�!6�`Kne<���K}� C�R	�����B��.s�%��xk4#�z�{�F[���I��@����9O�P�G �-�Ã
1#�ҵ�a�\p� HF\0=$%04�6&���|s�=��X�+�(Ș�6!Y@ @��A� �%�\!m!��-��x&���� �"�d�$bH2A�@�$@vWWg>�qW\V_DBBB��`B�)������Lo�l<]�Tٔ����i�>����p䋁v��%��hzp9L3�}���<��B�r6INp�27S�������$�/�JD�V#YH��KJD���V��R5aX����)���}�P�L|I!FWHX}L�����ą� #�cL<4u��04����Ќf�1�M�᰸ňE�E�HC�o4�����G�˚J�t2�%2%{�c��B	B0d~|8�\4�	x��@�{�7xp���2!q"C��t��aN�������m��\��������|�����`P�\	X݄�It�O	ck)��ZG%�s�s|�_�	���s|�_������W�5c�S2�\Ip˾�a� B���,���R���W���  �    -�� �hH �`                                                          ��  l             H   ��  �`t�]�Jҫ��6��Y�VL�n�V�P
PQgm&�¥��n̎8KŶF���g:��n[E��m� &�-�gJ�i�:h��49n�\�5J�umUm&��RY m  m�  R� ��^vm��V�;Z@Ȫ�k@:		�l�ݹ�i�h��� 6ٵI��  �$m�f��&���p ��� [K���B���I�-  m��m��&�k�[�]3��Cb���m�l��8  ,$� mm����i��ӥ�H�  �| $ �D��Mm���Z� �t�m�#��[l�m� 6��g �]�h�L ��m$׭����lN��m� -�}~�| �ͳm#��	6�`-�   �c]p�: 	m�גm�Ͷ p lm� p�`�  m�m  6�ְ:� 6[:H�+�h�6�V��m��6� ��J֝ӡPi�M5�M� l�'@-�l��m� ���f�!�m�K2.��Kh��}�C����+t(�uP�S��+�@ ����6�m�6CH�mrM��nͶ��ab���6�"��͂tG ����qAJ�*��n��䗪8.�)�;VQ��7UmR�!+�A��gm�ඌ�[��-� m� K�͗[��A��D�asz�jP[��L�ʬjj�˸v@66��U�;�T�j�+� 0�+����afx%AY[#Ҫ;��}hT�v-����p�J�CWdm������|6�St�N;N-4f�l��`m�m�:�UY\aU�ppY3 ŭ��u� >7�&���]��]ѵj����v�5m-�F��-��Ԏm�m�@]�j� <�n���_�j��ki6p��lA!��jv��%�m�p]$��    �����h  ���S` �irN���� $�:���}�a	�M�!�ڪ�P �:ظ�UcV������ڶ�hI6�@-�  6��  ����t����kh $ �H�`8M�l�Iz�qm 8%�6�F�6��h)iYZ�Z�%�.˪h�V�t�H 6ۧ3���6�ıx
�j��C�jWf��x]��V�J�Uc+�>�2*���UPq�R���浯];.�'����[iV��T�ʰ
��MUUUk�=)-�d��� 5R���\�UU�Ҧf���wgvi�X4��u�m���4T�IÈ�n&��L������M!��l���l��b�-��ȫ+ ��m�M�ݶ  -��` �y�:�m3��0�np*pF���o�2�����  �6�H[�v��m��&׈ր ^��e�ݰ�Z�E�N�ebH�&�ۀf��H�dt��W,ҰA��$m �4��@ �X���ͱ�j�b�h8�)j�YZU����hH��zt��� ��f� m�� m�$,0m�  El  %�m��Mְh�hm��BO�}���E�-�	m��YV����ɳ-C�N*�̩=�j�Z����jͰ6�q�Ŵ�	 v��#l�F�WU�a��de�\�۲�+*YKu��h  ��i�!�l�]mU�T���[Cm� m�6��(
������P�`B8`*��ݩGH
��@��UR콂��U��lpD��^����� N[d�m:p�em�*��X��)�-��$c�A��HM&e:�q��i$��6�O@���7P $ [v݁�I�lu��	l[x�/i���8��<F�f�gl�$�/hx����ɒ�pw^�d  m��5�����|| pH;m�lH    � -���3k�ku��X ,5�6�n��!h��eU��ױ��e(5��^�Yk8H �9�l �i�]mH8�`R�� 		$�f�qmdMd �t�  �݃�p]���$m�  ��Y��-�[���   ���Hm���� �$6�~��m6��m��C $#�����f��lm��I[�u�i1Ŵa��	�� Y��d�!�R��U]�t���*��V��UU�U�e@jTz �Y�-WT��@\���f�ۤ� �� �8�[@�m�j��+j�V�܈qvp��V��k[p5^m�f�[@m��e���lt�k&�z9:I�[�E�޴[@-���H��E�(��Ը��pR�E���*;o;4�d��m��p$-�m�`�6��l�-�6�08sE<9�̋RF�ٷݾ���`I�nٷ2�  Hėm�� �iM,涀K(���ݚ�������U@��	Z�g( +[]mn�����m l��yL�mV1T�<ʲ��'l �ۋJ�@/Ihq��   �nu+m��GP$m�  �h�	������M������(6� ׋wmz��\���    �1�\�嗖��7#U[
Yi.0��p-�;����� ��Բ��]���}G�[��Y�q�<��ᆪ�(���YIk�W�7fRUTX�(t���1����S��ڕز'n�m�͖F��Y@ 7m��Hk[�$�u�uQ]�qԯ7�]1	����u����j�eI�T
uH1�}���l&
�)�sJf;x�\�q�5���[A�f\��5$ ht^5���$   8 ,0��G[yr\  	-����� � h M�6�@ h:� �D��a~�|��͇�sm��I@	$� �m���&� ��� l����E8 m�ۀ� �kYĀI��m ���ȐH mmm�s}��ٶm����T�$���p    m����m�I:ml-�� l[�� ^� �� 7mm�[C�6�ۖ�  �ﾶ�ԇ[л�H�m���d���� �:�6 ej��1��X � ڨ ��-�t؛lTVҷ*e�+)g`��	e�H��� Y` ���Y��-�n���	�mSs��Cm� r�j@�uT�!5J��5\�$�j��m���vBBD���mUԵ [�Xe�� m\�i"JU�P 8$�mm�	 H�    �����Y^����h�d�� m�[�]��}oPfδ��uܷu��.�������  �$dpMpӌ_��������iVCd"y]R[n �D��I���L  -��lm�`m� ��1��UW*�9\�2��(�6�]*�� ����m�,�  6�m� ۶'5�ٻ6��)� ��[t^$��d�+&�l �f�Ce� ���	  m��l- �I&lmm&1� �l�	�5�Ɗ �^�-�r@�kv�g:-��v$<  h��p �i�&�(�mݶ ��$"Sm�)<��mUT� +UJ�Z/r�5�۱� �Ci6Ze��m��� ڶ ��8� 6�� l�h�H ����YNm�"��d�����o���-�۶�6�P�����Tc<­[Al�xq�&�p��sl��l4��0��v��Q�a�y�f�����:2;!5�UobS������
�;��U������v�%��[[l����v��l4P�ͶK��� �$�a�ƻ���%��l�im��L-��` �`m�mmm�  ���6�m�|� �m�q���H�'G���Ì��m�äl$$$ �aV�l�p�Y�	�u�XnhH�l�m�7"�6m�f��6��Em�5��R��ʴ�)�����	շ  i1�����  �h�aQ�TmUG=8U�V��t����mp	8K/mٖ��  .� ����t�V���IU]]B� �����l�U���cF��۝eGTvm��$R�e���P���٪�Bj��
l ���jA��(m� l\�<�ԦPx�:V��6��� l� $֚��zVm@��1*�Q�N��v��Ia��l� sn�m6ˢ��jd&�IH��8 �����h�5����P v��[:z�������"ׅJ�vZY�X��HU͕j��j����*��R�������}� "*A���> '���Ab��B!P�I�ނ	�h���Q��=Rp]UCR�$� ���J:�����QR �郧qP~@G��N��]< ���4}4�@��>��D���� � ��������!P���X��D����p��U��PW��U|�B�0�g�߄I�CÁ�����|<���U|Q� �pE �Ё�$X ��#�@RAA8��!�O�ꀆ�h/�����C��ц'PpO�@D��G���t\ 	���V!�Q+�(A|W�:����N>ÈuhT������GD8	�WC�1t�*�*'�
|3���VuD�E�"� �1����@�A�=N�	�z��k�W����q��� 5GAh��,"�D�EX��[ 5�y�>��x&|0\S�"�"�C��?0�� ��hz�	0`x�z(�H/���D������"@ $
�U "1Q5> CUC^j%D�=@0D�WЪ��S�=�������;EL�TA�b�bT�W ���
. ZAUj�@!�� R.4@�/-����ܙ�&�           �p  -�m�m����{-�Zj�w3�WiT��9�T��*9ݤr�f��2ڣRN�\/C<��\nS[2�25-u@�B�m��:판uU \kh�/-�U*�,rq��*U��n�8� ��K�m6�@�¨�l��(؋<���֣v��a���ӷ���@�n�h�9�'%�F6˞^1�ʓ�ⱍ��Tf��!�d�فw<n�
m���I�&�mR��v�va�p�֗�a�;u���@nlXwn�<�ۛD�#�q�n���6M]-�	�1��6�bLK,8nq-��͗�+FP��C�^�������[s�PrU]&`��6��u�;i����A�	�x�hq�R���mQ5vv7�6�
�nq�j�<
�]7[�ݚ�
�yjYM6�%����=m���<����]G\�˺��.�ٝr3���=m�� �k����S���R'�D8���WGk�ݸ���&��h.���[�8^A9�j���p���d��*�q�KUa�`���\tY���g�����g<�ʵ]Zni�Zۤ6��
ݥm]5��!YYj1��ӎ�V�]\O�--��q��xɵB[;W(t��4i��/,�u-�r��+ ;6�A[!��V�fv� �PIT���̪�͠��9j\F�i�rʼ���HA3�QA�u�Ԓ�g$�r��Z�]�����:�r��ziѪ1�`��GZ�#�ha��ʽT�6�tF��]�#ur�-N�1��:�7s�G`�WcR+m��uh�r�����v^b!��*<L����Wg���{<nn����l	�����K��ѝH
��kѼsS����h��4�׵�:�+lP�yy�ʦ�+�"M��������
�P:�!f"��A8K�:�c�6YK%���^M��"�4�%��~GCU�G߅T<=@�A5�UY�S��G���oȾ(
�F�Y����zwwN�w~q4�  ֱ�|D�m����s�E���4	l
���P�,��薺L��F��]GN�']��{b� ��ѱ�fX�6�pj�������v��my�#��y&�+�)^l�����'��M��Ռd<5���zÁ|M3��eY,v�5{E�Q��H{�6�G��P.p�����9�0��/6K6��s	�گ~ qy��7�/+�����q�g���*�s�9ݹ8=�&ܞ)����*��V�q�3b���>A�{�`{t����*p�� ���m(I%�
*��ݛ�Of�m�Ձ��iU��҃L�JI`n��`w+b`I#� �l��6p�V���*9qXu�wv��>�l��UW�����5�䨓�(FԊ���j�>�>X�s`}�nlP�(onwo�Qs�p��wP��Ɏ���v����컮9�QKv�x}zL�q������$��R&�>0$6:�)�m��)�����W�s��QUF�h��p�����^[�D�����;�-�0�FR-�q�8Xu�36��$w7���<X��"Jp|ljE`ff�^�
L�q�,��KIOkՀ�I�:pQ�C�
qʰ��,�f���u`fc�`lD%��S�9ɞ*��M�i�X�<�`��+����Xe<���\���QS�Q$�iF2)'�wޞ,�s]���u`w6X�ҥq�)J�v��0:�e0$��w6[J�?s�ČY���Q'*E�#�=�z��O=�����@OB*�"��PLLB�*BWv���=n��N���429L�U�}��`n��`|����۫tݷNS �#�SI9,	*D��͔��G���l���󎥭�ݭ/5�bj�p���T��h���c��\����g����
ɣ6Ef�i�՛)�$�����T��%����#�7wn�Ԑw7���<X.�;��:pJ9B�
r��������}�%�}�`I<����[J�$�iF2)%������w{��}����:�)����wG��
�v��,Ũi�T�*I�>Y%0$��fl��"`{�o�+o�:%��5��I�
F+mӆ��^g����*v����v��^����@�E�,��7wmX{��t��%�g7j�-���F��)J��6X�uX.�wv��9UUč�6�9L�l�INF�7^j�5wu��Uq/{޺�<�|��m�6パX{����0=�y���"`n�"B.��I�n;wv������{��V���:����I$�H��'�q�3Hh�4]�qg'9�$8�5ڷG;�	ݴkb�1�loj�<�QT���U{$�>y�b��EƱS���^���=����U�;-��li����v������� 8��B��Y�no4�.t@M��khݩ�t�l�EAlL �������n�f"�ۚ:�����T�u�θ�m���;C�V�][��{ ����>���{�{��H;�U���q�	�'�����.�)i��5�WN8z�뮂{ ���:���hp�����k�7^�5wu���V���Ui&�	JDn;�nn��
���ڰ7smX{��,Ŵ�F�eJR���+���`n��X{�,׺���5��Q'*E	EU�If�`IR&VIL�[���4H���͖۳K��u`fc�`jID%��!�ÊWpN4�c��ͼ����⚮m3���1��'#(<`#;f�nu��W(5��~���K��u`fc��} f=����&fٛ2�f�ۛ9$����>W�`*����j��{�p�����I<�w���7Y�$"Jp|l����]X�e0;%��IL�\r�J���\r��6"v�ڰ;��,=n��wV���Ui&�	JDn;�٥�ILI=�t)=L�r��T�UKJI�=�.\�Pݘ0њx|��6z�":�x��X��җH�닪"��o��������[��������]��L�H7���u~�+�[�v���`j��
�n�O���7"%X���$��w���VBAa)����WUB��ɚ���X���ddj)QG���U������ݺ�7�5X�Q�%N6パ0"͔��G��ؘT�����H��=X�[j8�>q<c���vimVl�< A�u�k�b�lq��`|�,��>0&V����L��0&lȒ�P�r�ך�ܪ��y��̀�;W�%2j�Z�\��HIċJ��ީ���[M����01a�E(ӌ�JTr(�3^j�5�j��X����]�\��m��l����T��H��E`n��X�V�o��{��Vk�V�H���\o������']�=��n����9c����N�<]v� =�6	�r4ȒNJ���+u�5�wv���7m�S!#QJ���J�06V���G��ؘ5R��'�q�Ȭך��۫5�u����R$�'��Wi�$����0$�elL	���l�(�
�)�*��y����W�=��i���j��$��D$�%	A���ߕ�  [V�s��h�B[��X��#��uOvc�a�8F �j��"�5�mE�r�i��v�z�C	����%`��&�n���"m��H�su�I���%�7h��Pc��i��{,�ݶ�=�}R�A���Kf��X.�tU{ckӭ��r�.�c�mw!v�α�bط&vw�m����cDA�n�*�,�$t���&훺H���~=u��?fٺ�f���'=pz�ٺ����k=Nն{���p��65Ƃ���R&�ؘH���[Vb�T�N2�FG"�+u�w6���y���y���n�[
�C��v��M����06T��%lL���>o#@܉$�u�5���6%
\�j�x7t���T]]+媫L�0$������%f��f&�E"��"&�H�L����$�V̓UR�C�;`���s�v�=�8�m����y���f�X�5~�*�A���`f�/%H���"�Xyg{�ß� �X	\�4�A��.@j `�@�|������{�w���5X��8(ܡӅ8�X�"`l���%lL����!P�_iUZ`l���%lL��5X�ҥq�*28I"�7^9�1D'�Հ�c�c�R��a���㋮�&�]n�mlV�m=�J�Q79C�<YWI�UW^����q,�Т��OO>0$�����&��0�c���	9�%X�5_�#}�Ł�Of�bBR�����
d�n�*⣃l�8ț���l�`n��gk*��r�'b�hQ(���DS���"�H�4_�5��~x��s�NK2� ��B�8���}!� ��#(���;L�;]�I��� :���Q�K�C��7(/I��`C�����;z��>��J9 T�!�F�z>�(��<5��L> ���ur�(�6 �H�!,e�D������|Q===���D�>@>+��~�H(�S5�� �UN��+��'�&TX�a%�$�׹�Z�3kvl�*]�<��m�Q8X{�^��+}���7^l�z#�*�o�,���ʓ�U����9<���ڰ5BKw�g��i`7X����'bq��Dt҄���2��UV[��۬]�q�*Ƿe��{�����͂n�WW΁�T�`lۃJؿu��Ձ�����$�JDI��ܚX�9�1�`7X��/*�gv|�O*\eJ���X�?~Vnm՞�q/y�����mo5��C���H�6ID�{�7i��󌰥�
!x �E���(��D�(Q�w���^�D�j��f�ÒW8���-JD({z|�=���\�o���w�jN�\�3�;,�d@�O��v��l�.����.��pqL���ww��?.�������o�OŁ��U���u�UW�=�V�ʗ��#m�Q>u�oTB���`n�ٰ3���ȯ�l�?��T�)�I��E`v������/�ݧ�g�&^o4�7i���e����P�8�X{�^��+s�Ł��U���=����W�i4�)&�6u����{����Vu�l���w��׻�zI�?0 m�r�"��ݙ�:��m��,��x�m�ap�Ǝ���#���l�����ێ�O"�Ia).�X��H�v�5������5��.��lUh��F��m`x�v+9�Yn�X-�L'GnNfO#vkv��jn��B�U59�a`9�
���n���&вg[�Sɵ�t��`\��������&9:��[<�9D��P��D�g�%/�̅�lۓiA��,�M�٪�a�&7k��4EЙ�mt��`(ӌ�Q��I���Vw6���y���秋 ��	9L�Ij�02l|~��H��y0&��0$�����$��>{��'!�U��=�>��,���
!EW�[��Z�r[�NS �#�87��ʮr����~���}6c�V�
"����ܩۤ���q�,ך����\����utz��`}��X�F�(��Ep⮸�tt{J۔S[]F��n�����������:l~�s���H���"�|f�Հ�c��3�	yDB��[�����*p���u���9Ut��BMBIj�|o;ϋr�́��~P��D%To��
�j�	8��%W&���x��sd�
l%U��Ձ�[�`|��F�eJ��
HXz�U\���ٰ3ڰ�sa�$��6�����`�#$RE"�;�۫ܪ�G����:�6�B��sR�us�4$ke�7n���5�4��&��_T�CX{.�K���9�\���t'��hI�D��?/��Xu�u�w�Ƕ�$�^{?�Μ�A�Gq��w=<_ꤏk�&���,���ďBωEYJ��H�p�5�ٰ;�v���H��D(D$O�P��FP��z<>Wď=\���.�;3g�1�ԩDJp�TryɰԢs���ݫ�2�as���|����t��r�N�`l���6#����k��`w��XQ����k��܍�����j�e`l	�:���9Nǵv�,�&���6��c\kW]7��6�&f��Y%0:��Q�R�#����V{�u`j��;ݚX��l`�#�Ev��>0"�)��.	��0�q�|�F���N9V���٥�w�>���R��^�t��盜����ۧ)�m��m�`}ݚX��́��`9�u`jJ'��*vU[����+��$�a�,��I4a��%�;b�N�s�<G,'��6Eg������r��3c�,���p`n� ��ʰJ�T_�`fl|`E�S�.n��򪪸��f�:pJ9B�98���Xu�j��֩���mX��i6�D�A6�>��,�y���sn�=_�鿿;�� Q�Qr�W	�8Xc��<����z_�VI���I>}�DU������UT���˝۾);jɇ�yy�����[�6�r�l�U���5����8%-v��{Jsn�g���
g�7n[yF��Bԭ����4�rs���rh�h&-v͉�Kg�Js$�m��cN��vs����Ft7�F�5ԣMnځ�ݰ���Â���	�ƶuh�lS<a�] J�	Bp�5C�lN�-�Lg�8:��QʺwD"�R���έ�S�V�%Z��\5�j���؎g>�3�?�:�jP�$��R-ۿ��]�v�٧�U�m=�ejt'�q�$�	�qXz�_��(�1��,j����m���UI�y�n�㉶G�H���K��ͅ��c�V�nՀ��mЂ1�6�8X~U��\�r���|�6{�VKn�6Q	)�m�`7G�*Q��7R;�ͺ�=�s���<���w=<Xֳ]��ԳD�*3�Մ՗��S=Y]�q:�\\p�ۮK���M�~��rɆl�sKf�t�I���`|�:�q֨I/�=�`7�=�I�%"	�������gj��E��D+�Qߍ�3j��{j�s׮�Ď���
4�*Tdr'!`{Y��͏��^[�S�/� �o�_vQwv���]�f��Y%0$����fk����7��' '%X�%0$����F�`I��2��*�k��{Uc��>��ܻp�j�qh��$�1��w/=;&�ŷl����72�������u���5����ڰ���-�F8��r'*��fk�W��߷֬K���o��
dn�veO$��*��s�`n��`9�ug����!B!@��?������Ձ������Rl�(�
�*)*�b"v�v�׶��c�S���`=����ێ��ͺ�=\���/����V���ٱ�"��N��ѧe��h]����ڐ�&�͚G��Ve����n+�J4�*Tdr'!��{�`L����$�u�_��'�W�vYrDED�����_ꪮRG�{���l�`n35�wD�o��Г���=n���,�U{h�U�羵`<����G$m�a�^Ϳ���d������/���N��+��S�x�<�տ���`~��tR��ێ	��yF:�=�{�~�X��X���?9�\���QƳ�'VM��6�)�W�.W�,in{=%k��ѵ�b5Ͱ<�E�tl��,��v����z��׭68�nRC�E%X����T���K]j�}n�ꉑ��ع���I�������fk�ܪ����Ձ��>Xf�J4�*Tdr7!a��(U�}V��j�s��������ߋ ����JR�DH�d�����XI%	yD(��]ۼ�`<�X���u4�%��?1��4��5&	 x �*�! u� ��(Cj+�TtC��4�"��XFC��<��p ���Ӑ�:!��B"��
#���}���X��ߵ�'"��"N��ӹ�g�@}�s��~����F��           	  � �NSIm`J="j7F2��f��V�Y۩��X���y㵳�N�My���X��VUU4���,@(����ݝK>эe���WT;Y�5rJ���:*(��C�'4a�^8�W3��!����(9�ЀW�~���\j�u�	U�(pU=v��S�fr�K&ۗ����h� �5�6�N�Um�l9��J��i�g!MF��bt�zH؛�љ0��wI�L�W�={vݭ�n�(���]�E�5��H���-Ћ���v�	Z�%(�6,<�'cC��ﾗ]%��L�-�L��-�vؽM��tnD*/
�͑���Z[%QU��>�V��gf�c:��F[h�
4� ��tӀ$�Tm��i、4u��U�M���t�u&�u��Ry$��[��bѳ�n��^����V�]&w&�s둶EJ1���g�u�Sң����Ғ�Mㆀ�e��ꕼ �T��97.�-������t�UWk��A�Ƴmۗ"i�Q8��<5�Wj���Z�+��2���Oi�N�H��$u�K� �U�/.��u�`U��RNz�m���R[]5Mcnd�1;�l<d8�`�a[uV��vY�ݸ�����ÛT��[Q�a��VW�����n��U*�f�,�ٟ%��@�cbF+��^�Z��+�l�H(î�@�Km���jc����\��j�,9-���U�r�[���؜ۘп}����Ƹ�;u�-m/.�!��,N�F�(Vvə�nJ����+K+<��m�f�����ܣÀ6cR
8�nb��z f�e���jˌ۹C$Y���s�Ͳ�d��Ov�Xl<�- ��5��n��(*w:0iy��%\���I)4�'.�����U�b&C �
%��+4bȂl��fm@�����u�xH.�$j6*ܩ�E�#6]T���? x����b>��EV����::	P���A}O� �b������~�~����=�g��v���`gv��ssx;��mn���N�9�#1�]�̨G�ݭ�!we��o2�:�l���P]]f����w]7g<����.;jw<7-;��r�I��v��8�̏#�:���vt��[�8;Z8��Y�j6]a���b�{g��m���xP՗��5�m���<ݴF���9��Ύ
I�d�L�������{�����ͯ\��|=�G�r��9~����p9c��c.�&��ń߯w���_}�0Tb������V��,�c�Q�����i��(���H�̚_����7�`y�֬=n�fMM��J�1�I����|���՟�7�o�;��?v���%6!�dD�������6Sn�{��d�0=��C���$8TRU������{v�|���`own��xА����9N�g���=t�SvE*�l���+Ht�%�N����U�m��J$܏�=�<X�f���^���A�{�2t�!L�k�(�n�n�I;�O�����lz�0$*M,�rDo�߲Ձ��Հ�8� �3��)I"$n2G`own�]�vz����`{�v��7��hJH��Ws]���Kz��a��S���v�߿��N8�drB$�72i`j[���nnڰ�X=�M4�R��j�ɵmQ��"ݘZ���)Đl�u!-;/��:��v�3��~�nP����X�>z��{w�,k?�(�M�t�DH������H7�������F:�(�U�����UKr�*)*�?o�Ks&�v������)�����P�}���omX���$����MUs���KТ"����΍�X�ڰ�ԡ$���p��L�r�8���X�b�mW*���W����72i`b�5���Pm��,��u�n�z��1��[��랓5�<
�}����!	6�d��=��Հose���Os��o��v����+Uu|`6[��|��/��D�0&M��r�#��i��D�������`>ю�؉���V���Xd�B�TW(��W&k���G�yپ��޵rI�~��O����`+�b�EF"�@��� ��PD"N�(K�B^Y|��`k�{�
2Sb6DH���Ձ��S���:�z~,�3]������HtF�j�Ϙ[{%m窫�j��{u�k��CM#��>�U�M��r�uQI_ {7����2�}�j_Hnnڰz�VIS\i��rKs&������Y������]X�6X,3h���)�q9#��7�l���l��=%�`M�]Rq���m�H���Հose���K/d7��;�X7�r4$�"qʰ�|�<��{w�΍�X�ڰ�!#a@�E$>:N߷� j֕�4ݗ.��[F���&��f�;e%2�c�ɡ,�/n:<��N���9u��mntD�qN���HS�4d�+�Y̨�q��K������7ۜ�j�m�qe�&ǰ�r�͗v Z��2������瑈XH�aM]�^r�$4�4��x�F{.c]��2ݳ^��L��h*c��ce-��g�i��v���Vn웛��7sv�"�G�Ż�̎T�\%���e@?���c���5Ҽ�a��K(�n?>�ﮏ�a�q�I?�����u`>�i(K~�7���l�
T��qĜ,�3]�J�${=� �o����K:��I(�Q�t�h���͖��zK����=Lܭ�����D�2���<��},7�,�1Ն�����X=[%�\T��j����q��$��G���t?zՀ>���ɖQ*iX"�ԜT6��ꀄ����]��N�L���.���,?�ur��K����T��E!��o���ݫ }�͈P��o�X���j20m����ݺ���8Q�G9T
����~b ����9���$74�Q��В�P�Pg����G)	9�r����,̚Y�UW9I{Y�v�޺�7tSS'$N9%9,;T(��iޖ�j�}nՇ�T����`~�O�J�cn8����f�`L��L�l	�p`w	>Zu�#��󞍲u����6r(W�nN��7:�4����޾�}���ѩ�lnnڰ�|�g�}!�Cڰ7k|P�m7*'Q��`����\�Uʪ=����[�z�%25�l��&�Q��m�,n�����Us�����s�S�}V(	����s�V�����)(��J�Hڐ��J!N��`nnڰ�|�ԒQ:���i��m8�H���$v�v�����V��to�X�c��|�g�j�Ie�F� pZP��+s0=���)��˝s�`1s[�m;/�I�����>X3��h�Z�!B_Hnnڰ=��q2rAD�5���ɥ���BS&�j��ݵ`��~P�(�%����R��ێ$�`~�{�7�ڳa(�7��������1�<���C�ȉ�������`�zX�4� ��H���~<��O�����r�pj���{�,̚X(�V�v�%�ft�T��D�:cn�Kiz�q�Ѵ\�Z��	3��{W�uH&�EK�*�J���Cp��Q6���?���}n��_H�y`vY�
ySQ�*9#jB�޳5߹I�z��=��`nd��W*��������q���m�9ʰ<��V ���l%3��Kr��`V����	9�r�=\�K��K�_��6Sd��	�)�T���H�n;s&�����|���]X���	|�(�;�j٦�$�I$�R��)LSӎ��n�3��7X���u*�P'�89pb۸M؈��m�,p��M9�����$n�N(^�I�=N�+t6q�D���6�U�Z��'�Ʈ����oU���4t�]Y�� ��1w�5'�K��i�k�#W5).Vy�=�Bo8V�M�4Н�hmsY�]�"{.�Em�ö�p�n#I�'!�1ݷ-���W��������?GSrKn�E�Ω�Ə\n�5I6�7����]�2v[�Ɉ��=�}ͯ��cn9I8x������Ձ�����|�۳Ł����(�Q�t��$��ڽ�2l����J">���<X������J���F�j���]�v��,�3��l������Y(�
�5&�v�8��~,f�����a��"�Ǿ�'M��B��s��Wcf��s��w��g��7n�W*�sވ��tӔ�R��p��ѫrK��z2��\�\r��n�q�=#5ڍ�9�0m�!�{=�Ws]���O��|�ٰ�׵�|�#BNB'�o�w9��EA��`F��	�XD!F1"�2@#
A��,��#�1"�
��P������ǯ��`{7���}ݺ�s�����Ě�qF�#�R;ۼ��}�l�y(��?zՁ�{�ftR��ێ$�`}�V�v�����a�r�{v�X��B��)��WE����J�����0;6�V���)8��(���>5L�r=�5Ԫ���ڈ�'5��Q�������_n�-7)GU���|�̚XnCW�B^I%�?zՀ�{�d����MO'����v����"`L��6S�U�~�r��1x��)F�eJ�Hڐ�3���`>�j�"P�p�BĜD�LB��FX��Hz��a�EMD��U~B! �q�*�Ø�}Q|P����� j���$}@�z|�@�ȡAHH��A<=R$	��ثBB�� ��0��r(�>�y���T����>� ��=����z|? �>!�A鋂+�!�
�{��	�!�% "(� ThpU]1����:��O�3���$m	��"�؈�;��+�=��q��89���:��$ܡ9*����`z��V�z|u�ٳ�	%;����sd7��Z�c]��%���i�.�S��Z��Y�>�+�p�s��g�v4o����E�%�%:�!U��(S���`w_���[���j�~v�_���1���,�!��2G���L	�p~��$IG<y
2T���ڌ���{�V.�?s�����OŁ�����y���d�ڜ�qXj�.��X�4�>y�͆BK�!r���\����2�5%b���7WL	�p`{�g�<���|`j͔��\�W�Vy��"��TrI$m��E�e���&*٧��=�2k �١|=�K$e��x��}ۂ'!F�5!�?o��X�۫Ws_���n��7�JS��6��r0&H���6Sn�6ȟ���t'�q4�nP��`yf���4�ԗ�a�`{w�V58⍪��d�a�W���`y�M����qՁ�5mЁ��6㔓����j�?W���{�_`r""#��	r?��>����~j���W�ƘQ�IG
�̊�aMMq�]0��_c�zVݒXy\Bt�Ŵ�y�mm�v���p�Ӯ;2;v�N.�,�wO1����T����;i�`���t�R�v��ץR�P
u�Y�lܹ�+�i�t�-�փ�V�:����9!wl6���n,칊4���;t�����ue��;�P�S�a��%�Ͱ͆[�f[�6[����N���C�=Q�q������i^d���%p�,�Ks���^ù��u�"�UtZ��H���6Sd�0&m��܆�q�ܩMS�U������L���,��`<�j�)��S6H� 4�I�����`or��)/n���=��`w3@J&�	�ԅ����1ڰ�XlDB�ͽ,�o<��$m	6�"�73n�Us��<�?��zx�>܆�V�RBryΝ��v��r��9>��ڪ�cs��˓k���R���i�N4�M�#��Vo�������%
��ڰ��iY5ͷrl�3n�rI�{��� ���8�� ,AC���߶v���u`b��6��mЪ1�6�k��ל�1ڳ#b!(���ݫ���`gY��Q�*SI�mFEa�z��DS{��sv��8�(�
z��́���C��ܨ��� �����vi`w�VfmՁ޽hM�����:���i�:��L����6z�5;�1Z|������*�RV!�@i��RO���;�����1������H�
d��(��X�Vٛu`n�>ǚ��ă4�y)N2H�m�Ed����rI<���LCc�҅AfD�OkE�O�{��9��I����䁙X؟�nQ$�`f�>ǚ����a���ﾫ��o�d�FU�r�Wl�lLl��.��y�wgw�L:Q� �D! X) ��{ے�6�ݹ���M����:5fv.E�ٻ0�c%[��H6�8���e�4��c�m�	��ו���3n���?=���M��q�R�H��
�R�x�6َՀ}����+�DD}!��yX���r6���nB�r��ݖI���_'�m����x �{��|�����{����͛&\�r���A�66(6>�{��A�666?wz~�|�������>A��C�S"�C
���v7{���A�666>��Y��l���7s7.��>A�����Oׂ�A�A�A�A������ � � � �{���� � � � ������ � � � ��ߥ��nW=�%�emӣk#rm=�f�8������[��E��#���\֩L ]w�|�������>A�������>A����߹�p � ��A� � � ��ׂ�A�A�A�A����.9���f�wt���lllo������G�b��A� � �w��ӂ�A�A�A�A���?� �`�`�`�������
�A������\��۹�4�wx ���s�pA�666>�z~�|�������� �`�`�`�}�o �`�`�`������%�rf���ͷ6pA�66/��<*��A������� � � � �}��Â�A�A�A�A������A�A�A�A���~�|����﷭�d�&�I�fe�o �`�`�`������� � � ء��E\�����A�666?�������lll{���x �Ơ��D``�A'\Ϸwwwwwwv۠ۆ��=�.�-�eհ��ON5�0o�����\.���D؍���7��Ġ��^lv2.��aa&W�n�h�X��rxP䨷��D���r�;-g��Y�n^��ؚs�8��ag��I�g���9b�2\���#|d-��%��3��IM���� ��� �u�]Sh����8�V;;!�sX{D]��}���o�ѱ��W�m���OMI=�	í�n-�rZ�ٱ�CM#�<���?}�@���������`�`�`�����|�����s����lll{���x ����>A�������.�&L�r�n�A�666?���ӂ�@,ll{���x ����>A����������A�A�A��w�-ˆnɻ��fn�>A����oOׂ�A�A�A�A�������lllo���x ��~���� � � � �~���Lݛ��\�.�x �[���>A���������A�A�A�A���~�|�����, ����^>A����_���[nfi�n��� � � � �w��A�666>���ӂ�A�A�A�A�������lll{������lllo���_����-��sG�˵�2���<�\���/Xd{,��E�4�5ͷr�i.�� �����8 ���zl����	} w^��՛3�Hr�\cn8����yZ�W*s�v�Wf컫 �we��٥���R��*P7M�&�y�Հ|��̈́�)����kU���hm%q��.H�Xz�Sy�ߥ���x�3��͇�#�"����y
l��������������6���� ����J!%�3,��S|B)M�9����*�Ҩ撻7OF�L�/cժn��fԺ���%K�&��"6���ǵ�����vl��p`�O�Wʻ$��n���۫�W�},g��a���v����?r$�n4I*�;�y`>�2�G�	T@����T�<�o����շJ��6T� ���%����,���`<�j�>x�`>�[b�m��$�`b�5���_ w^��}|e���B�T�rUR��;�}�m����s��EE���lkh�ݫ\��Yr܅8���N��l����ͺ��6Xݚ~��j�<�W��C�*��I%Xۛ/ߛ?o���<���73n��W*�37�J�jj*j9,f�K'0ug�g^� ���RƉm5Dm�7!a�-{����o������Q_b�Q�P�E
��p�4`t{Uu_[�>,��x�)�I���<v�/D%Y��:��'0u`o���7g��k��f�Nx 
�[��٩+�)��<��E��v��6�^3zD�rU�}�������Řk�9U��޺�7�^�T�I�����ɥ��������`g��V����)�1�ͦ� �Q�I��պy�n�՟�����o����Ł����DtJt�e�t���vl���{�}�*C�����C��H�� �se���e���:�>mڰ2#��BDB��Φ���i�O�z��#ŢT��{0$� ��0�C�fs����0$�$�FZB���+``'��ł�����a
F Bb �� D�F$�t<N���$H҇ΔE���Q�==�HBIFH�	�!	�`�#		��C�zE��$��̒1�8~$dL-^@!0��1�`�/k�I����m�o��v�$            	  @m�n���&�֦p�u����>��� �+U)l�xl賺�E�t-�6�@��sss��ֶ�X���f�@T�UV���6�4Β3�X���=�z�VӮf��*�2��cN��gS��$�[`�u�1�\���S�����(��L�\��m�&n4���y���;���Y��kuj�۠��"�nM�M����t�+�8�G.趲U+�5dݶf�L��U���]j�	zU��f��&Gm�m�pK])5���6^�MY�Y{�a�C��nV�:�[#�t��������8(N��3��C=�Ɋ���ZA ��R�:����D�*r��^xK*+v˛&5i'S�! Q���.\v��	��qpn�@�Ӟc��=�)�Z��*���h�N�i�h�-pn�1mf8�������P,���P�[�Fڼ�:������m��q����T�6v�9���I��Mli
�$��۝���zH������5�E���0�7UZz"z@.֥Pz^mI���˵��bc=8( �F��N܈�uRq6�r��(n�$pU*����	���@��2R1T���.8��.jAIQ�N�L�Xx�7�k�1�]m�v�(i��u#����T�#�vfSlV�U[JR����mv��Z�p7�Y%�EJ�8h�����g"KÐ7Vymfnv@i:vں�P�v�HXn�ݫ��Ƌ/-V�
���[q�=N�[��6U�g,�SiW�ݒ]�i�n6	��U�
�+9z�l�m:Ʈ�9x����p�9C��s��@�[+�mT���K�N�Nڼ��@r<����	뵫�]�g t�Az)1$å�b�!
=a��*�҆p�w���u��9֐@<3НN3�Ҭ�8�h���Ҫ�Q6�p�,c���3m�@���L��*�"vڎ�9n\˓3!�Lٟ�*�σ �	��HT��碁�P�����G���N��!�h(�*�z�%����������m+W=H�GZ)�n��{'&y8�;p6ذ��:�Bg��[���\�s�1�h� �^���M�K��u�pm&� n�T��c��C��V�ySo���	��":�ѫ�NAVSu���i�͵�)�-`I���v�Rp�J4����!�^ɂR�S�^a�%a,tَ����s�%U(��/*F��kЮ�k����m�e��M��4�6���i��U�VV
Ȼ��u�*Nsǳ�sjڝj���{޾���YMBMEMG&�����Řk�>m��.���,:[�MT��y'*��U]�[��d���e�7v��}�?USa��/�j1�I������ٲ��p`j�%0�k�H�����R9%X{�w��`n��`b�5�yw���`o��t��8�d#�'%��ۃ�Ҥ=]'���;6[J���x��Ӊ%؝v�$�/�'CY�n:&�j��^a%Izm�[v}��g_|;Ojʕc��fՁ�7j�>x��IB��1�i`{Y[�DtJt4�6FG`}��W�T����ZQJ}|��,��Xc��`n��8�QT�!�J��607v��%��<��y�'3����QSQ�`fd���V��ݺ��R]���=���&�QDF�)��[Ș�>0��`n���n�*��+[)p�4��$�]�9rA�\&,r�������ՓYR�j��b��d������p`wky �&�C�D�jG$� �3e���RF���<&d��	5G�E�V��eՁ5�X��Xec&�J&	q(2��
�T��n��͖zn�dN��mI
I����M��޺��6X~�����`wޅ?*#�S��M� ��c� ��lݸ0;��L�)-]P�X�9L�y�x�GS��n���
w\[/j#���v�F��uW'$�H#]����lݸ0;��_��'��������q�SMiI,�M/�*�;�|+��]X{�/��${o�M�����Q\�`w)�6�ݫ6"���ܰ7v~,�Z)I�IM6��Vۻu`�>X��X�BR��A	D«*��\��`W��4=�I����� ��lݸ0;��L��������q���J����iקn���b���l�t�:���5�õ�s�b>��y�wSl]]�	%�`w+`��>0��ݹ���=�T��H6ӄp�>�����yU�z՝�I(�n��`6�����2!Г��`}��V�M,��n���`ekݡ�F⊤i4���'[�,o�X���)���X�x)YN:��DNs&���I-�='�:�mX3��.!�	Dg{��߻�{���i�  �6��fwj�[[[g-�Hm����B8� +��p����W[����a��C�$닍֋I���)��]>&���s�sm��!�ciTNɃ�Ӓ��ڳ����9+nk�0�4� &:�l���[q˰\��f͵+�TV�1,�b�N݆+�\2�lO���M��8���W`���
e���h�λV^-t� _���~���k�E\�'mH�z�� Z�i���fJK�`�k���Q"4����OI�>��X�c�yv���ŀn��
RqF��i�+�ݺ�72i`w2i`o^h��RA��t��l�H�X�|��M,��K�4P�v������M��(m@>�f��	�ݑ�6S0��U��vUR��
�`w+`����w�V�S7f���51R|��6�F�������������
q��iKg�ql ;��:3�UUդ�����ś)���s�3e�+k�ޡ�F⊤i4�����F7�,�8�l��W�Dz���)J�q�� 5#�7ޟ���Ԭ�v����k�7��A6��(�Dc���DD$����7޵`v{�����L���$Q�m�"Vۻu`v{���q���9��BI:��SV�9L��غ�>��߇����)����[9��v�c�`8^7�]�*n�����l�q��q��%�^�uϭN8�d#����d���ʪ�=��3`u�ڰV9����P��\�ɥ2��HN������n�Y�Us�Up�qJH�&�.�j�ly�,�Cj�ȇBN�q+Ի���`{vx�;�4��\�/fߒ�6�����nF�H�*��&��϶G�M��ٷV�xЛkI%6�q�R(0TA�ruў��{9M�=`��ta�i����^�[�����n��q&vG�}��,c��	��D�h�rw&���""d�nՁלe���2��<<��"�mI�;��Ձ�ɥ��ɥ��ɩX՘�4=�I�n)%qXl)�w����K;�s6��!.�
�Us�rw7�Ձ���ljqģ!$\�p�;��XP�;ٟ��ݵ`u�`�k�#�6M�D��T��&v�ɒf�Y�r����8��&n�ɺ`UUhX��ۉ0;�>02m����K�3uQ�I�c�%`}��VM�03v���ۉ?q"rW��E+�U#I�%X�,�&�w&�`}��V��YN:�1��$�a��w����fl���J">%
�_�X�[�i���F);�R�5(�{����,�8� N!B����w�}����9>j��� fY�d��V�OLtn룚7g��IJ�fwfX�O`Y���é;e�����-�u��m���l+;-[/X���kv뫮P��3�VLiw����q֝��n�&&ݚD�����]8Нf�t۫S��6�HU\t�H9�z��4�X�;[n�d�c��Q.!�ѭۧK���s��t��u��c��j��e�8�M�7_�������0����]��M�tmӛ�K1٪��PF�7�z�5�����&��5�g6ʥA��|��ɷwn͸�������\�:�fmݻ��"X�%��~�g�~9"X�~�͑9ı,N��~���Kİ~��59ı��կ�qě!$�/���G)����"r%�bX�{�;oȖ%�`�����Kı=����yı��5�����W�jP�W�)�p�;�y?^'�,K����Ȗ%�by߹���%�bX�w���,KG+r��2"P����9H�!,����bX�'����O"X�%��{͑9ı,O������K�R9]�jj18�h(�ʢ&�����Z-\�$s���$�5Rs�ۛ7&Ib��\�t��Kı<����yı,N����,K��߹;x�D�,K��ND�,K�~��7p�Y1�����%�bX��y�'!��m������%�bf�����%�bX=�xjr%�bX�w�vq<���L�`���\�f��.�wdND�,K�w���yı,��59ı,O;�;8�D�,K��6D�Dr��G)gL�Jrpl���_,K��{�S�,K��s���I!I
HM��B���KR�JxB׽=x�D�,K����,��m�L͹��jr%�bX�w�vq<�bX���~��ȞD�,K�w���yı,��59ı,O����_�ͳss(4��\��S8�*�������/���^�X��̽�ݟ�����'Z����w���D�?����Ȝ�bX�'������%�bX=�xh�<��,K������%�bX�쿹p�r�v[s.�sdND�,K�~���y�DȖ�߸jr%�bX���?N�*�ؙı?~�͑9ı,O�m?~)�6�%�\��6�<�bX�{���bX�'����O"X�|D�#�
E���!��d�:�n8㹳g�z1�'��$j�)"�~��"����"EC�� ���А�T�!��M���x!�s��4݊Xv4�����$4�����i���P�^A]0���0�ܩ�4T�֩T6�ߖ0b\�@����߀�=����:�AC��
���|x�<DW��/�����Sb{�}͑9ı,N��'oȖ%�btϧt�2�fݦ�\�t��K���Cb}������%�bX������,K��߹;x�D�,K��ND�,K߾�K�3p�d��nl�yı,N����,K��1���~�ObX�%������bX�'����O"X�<ow�w�?7+��n�	��J��2]���b��[]�!��3p]p=��*�vH�3�]��,K��߹�x�D�,K��ND�,K�����'�2%�b~���"r%�bX��~��l�7fL�3,��x�D�,K��NC�"�TB�k�.�)!I
H[�|V%�bX�{�;oȟ˕2%�a��]?pjFEp��9H�#��V{o���%�bX�����,K��߹�x�D�,KﷳS�,K��ݽ�2e�6�ɻwM����%�gၑ>��͑9ı,N��~���Kİ~�{59İ:
|��@/�S(�w4Q�M����yı�r�E����JF�l��U��r��'������%�bX>�����bX�'����O"X�%����Ȝ�bY�G+�+��GQL$*q��
)(|"n{h���v'1����Yyd�R�d�@��\wI�"B��2����}ı,�o���Kı=����yı,O��6D�Kı>��v�'�,K�����l˹�v��d�ݚ��bX�'����O"X�%����Ȝ�bX�'������%�bX>�{59�*dK߻����i2L6KsgȖ%�bw���'"X�%���s��<�bX����ND�,K�������2%�`��߉[MDICt��ʳ��R9H�nm�+O"X�%��w�S�,K���s���Kı>����,KĿ{�֥��6��W���#��R+�٤�Ȗ%�b{߹���%�bX���l�Ȗ%�b}���O"X�%�V�|@$ ���{���n����U-��з7[d(t��ܞ�ٳ[cC��Eu�ঞ�Q1��;j�a���Y׬�Ѝ)&�&�ʱK$Y��vWL��]
�qq�.�g�8�d�ؗ�����M]G[1FD��V�q�.��s�ښH�aM]�^r�q�Ӹ�udc�����lcF!v�ƃ��ri�lAE�X�:j{�Wg[@��O9In��>@S\�̤&y&���nCA��4FM�b�F���^fJ��t4��c��%&◫��e��n�ff�O"X�%��{��'�,K����dND�,K�~�m�~g�2%�`���59ı,O��y�r�n�ݻ��l�yı,O~�6D�Kı>��v�'�,K������Kı=����yı,O�/ynY�m�̶��\��,K��߹�x�D�,K߷�S�,(��߻����%�bX�w�6D�Kı=;��.��7e˶e�ͷ��
HRj�F;Ӑ��$)!I5ޖ�D�,K߻͑9ı,O�����~����{���翟�Ib)]5��Kı<����yı,?~��6D�%�bX����8�D�,K߷�S�,K�����<��L�3M&ia����R5��Vɺ���ܻl�g�t��7+�)v�i2L6KsgȖ%�b{�y�'"X�%���s���Kİ}�{4? 3șı=��~�O"X�%+�kޡƚ���Ԧ�U��r��B}����y R
!�Dȯt�SH"�|��K���S�,K�����Kı=����,KĹ�[ĔC�c��#��9H�#���~��ND�,K����'�,K����dND�,K�~�gȖ%�bXw�gY�w$�۳3f�"X�~D��|�8�D�,K���Ȝ�bX�'����'�,K������Kı;�os̙uͷrn��s6q<�bX�'��6D�Kİ�ǿw�Ӊ�Kİ{��59ı,O;�;8�D�.�����S0m�������v��<�M<�gv�o)���;w-m����h3΍Y��6K�"r%�bX�{�;8�D�,KﷳS�,K��s���Kı=�y�'"X�%�������lݗ.ܷ7vq<�bX��of�"X�%��~�gȖ%�b{��mND�,K����'�,K����f�&]��ww2]ݚ��bX�'}���O"X�%��۝�9�"(�P�Dȝ߹���%�bX>�����bX�'�}җ�f�ɖl���'�,K����ڜ�bX�'}���O"X�%���٩Ȗ%��&D��|�8�D�,K��߉w.]�t��I���"X�%��~�gȖ%�a�X�?MO"X�%������yı,O{��S�,K=�����~F�a�6��{���j�J`{�y ڮ3Ń"9�ې��WAE�/���3,����%�bX?}����bX�'}���O"X�%��w;jr%�bX���vq<�bX�%�{���2�䛻vfl��Kı;����yı,O{��S�,K��s���K�Es2i9Vr�Mr��G+��7��q(�ۻ���Ȗ%�b}�s��Ȗ%�bw߹���%�bX?}����bX�'s߻�O"X�%���{�f6���n.l�Ȗ%�bw߹���%�bX>�{59ı,N�w8�D�,/��(~T�j#�T�U���Б.��dND�,Kû~.��7e�4˛�8�D�,K�w���bX�'s߻�O"X�%�߻͑9ı,O=߻x�D�,K�ܷ��7M�Pm*��';�jc�#�݃V���(��^�ln+�k�n�aخ�CK��w�{��"X�����O"X�%�߻͑9ı,O=߻x<��,K�w���bX�'����nᤳ,�s3s��Kı;�y�'"X�%���oȖ%�`���S�,K��=����$�$�zL�e�[����A<�>���	 ��؛�;����Ȗ%�b{��mND�,K��޶�.n͙�fwoȖ%�`��y�Ȗ%�by����yı,O~��Ȗ%�by�����%�bX��K�\˺f��ݻ���bX�'����'�,K����ڜ�bX�'��ݼO"X�%����"X�%��!�pi�Ā{�t�^���ޝ��~�&�� ٖ_j�1-�[�<xƳaٖ��\ԣ�P��M��۲**u�+����.��:�A-��&܌�u�A$;e��������`�u!v:�+YNpnշA�W�u�/`�l5it�J�l98�ۦ�p�:�X��m�Mˈ�����;f���+S�m���� ��E��Ѱq�^�y�\:��� �c����!uW�(4r�c �w��mNv�����z�����ct����ŵÊ��$�:���5�s&@z���'U��ss��Kı;��mND�,K�w��'�,K��>���Kı<�~�q<�bX�'{/yK�M�72ۆ˛��"X�%���oȖ%�`��v�r%�bX�g�w8�D�,K߷;jr%�bX��NL�t͓v\�eۛx�D�,K���S�,K��=����%��a�2'���jr%�bX����x�D�,K���Y�n����˗v�r%�g�VD�~���yı,O�����Kı=�~�q<�bX���n�"X�%���;m��i,�6\���yı,O~��Ȗ%�b{����yı,s��ND�,K����'�,K���'oN~X��`��]#t�6���-l�e�v����CԜ����Q�v$H��gi�O"X�%��}����%�bX>�ݺ��bX�'��{�O"X�%��۝�9ı,K�{z�t��6a�fۻ�O"X�%��}۩�b(�����`$X �E���GЯ"r%���|�'�,K����Ȝ�bX�'����'�,Kľ����2wr��ND�,K����'�,K����Ȝ�bX�'����'�,K��}۩Ȗ%�by����̺�۹7n�ۛ�O"R�TB׿p!Y
HRB�V=���%�`�>���K��
�"{�s���%�bX���0̻fne�6IsdND�,K����Ȗ%�`�>���Kı<�{��yı,N��l�Ȗ%�b~E���_�n�ݶG]��p�p��[d-!q՚�N4�bS<^�g6�p;��6̈́��������{������u9ı,O3��8�D�,K�w� ~'�2%�b}�w�q<�b]�7������"b�D��}���,O3��8�D�,K߷;jr%�bX��w8�D�,K��sS�,K��~'d��i2e�.fnq<�bX�'�nv��Kı=�~�q<�c���b���V@Z!p�SX)���{}>��ns�jr%�bX�gw8�D�,K��3r��7I�t��jr%�g�U`dO����'�,K��;��r%�bX�g��q<�bX�'�nv��Kı/}��m���ن��˻�O"X�%��}۩Ȗ%�a���~��ObX�%��w?Z��bX�'����'�,C{������V�9Jt�����u�X�b�U=��׺ۛ8���5�r�8z�ۻ7r��ND�,K����'�,K����ڜ�bX�'����'�,K��>���Kı<���Y�\�w&��6���yı,O~���~c�2%��}����%�bX?g]ND�,K����'�?eL�b~�/�S��ss-���6D�Kı>ϻ�8�D�,K��n�"X�ș�����yı,O��͑9ı,N�{a��L�0ۙ�]��'�,K��}۩Ȗ%�by����yı,O~��Ȗ%�ЌQ�� ���!��w؝��%�9H�#��V��nPƢ�)#n�ݺ��bX�'��{�O"X�%��۝�9ı,K�wx�D�,K���S�,K���ܲ�e��.�l5h��k/\�ms�6��^�A��	��F�V�v���Mng��5�g�w�{��7���~��Ȗ%�b_}����%�bX>�ݺ�	�L�bX��߿gȖ%��r�g�C�5%�ĹVr��BXʈL����'�,K��;��r%�bX�g�w8�D�,K߷;jr'� eL�b_�~��n�7f�4̓ww��Kİ~�����bX�'����'�,�"}��֧"X�%�}�����Kı/ԝ�p�wLݻ�wn�"X�~������Kı>���S�,Kľ{�w��K��U�>����Kı=����ɚ�ۙ7n���Ȗ%�b{��mND�,K����'�,K������Kı<�~�q<�bX�$�,A�9�tC�:!�&�|Rp����	a1�wT��1V�@"�B�N��p��^sUHQ`a:iwl	�q���z��,0�$Ti�r�.�<ZP�0�
>GT~JU�'��j� "�� a ��Ő0�Q�>�1���F� }K�X� a���H�N�ee���规#K�@>�|����4( |����! �0>�������m�o���[x            $  	 ����f�JƎ�v�"Ssfq��4�Ueeh�X�-��Tvz��"r��m:+���s�͓q��$芧e��E��5ʸ�;-�Mn�b8Qu���pl��+*��s��x6���j��yAW��vP#����1V�D��=���;��uF�m!��Ʒ�YvV���cĖGuc��u� ����;	�Ĕ�R�JrF���Z���j8�TV2=�+�s����&��x{���Z9z�IE���C�m�������ιG���n�ֶՠW��pn %3�96�c#��(yz`.���ݖE���k��J�R�{��n���RY%�t�$T�Z��)p����!8�kJ�,�]��+Wg�ɥ{R==63]��1����͊�Hp�l�7,�E�[�Z�ZM�WYǕi���@�=i�$�\�K�:�HJ�q���1Um�*�u#�]����̃��O��d́��M��;q�dܕ��T�[���ԭ.FBݧ�;u3����
G��s��qB�B�UsYrB�ks�T�ڭZ��25UHs�qmn:�V�n�6��؎����͝6�v�pt`�sU�N�qMIm���ʑ�ݻT�Լ�N�3�#����9��́�9,P���+��)�b.�d�Ӯ���`c]��	�N�Se�L]�wc��(T6+�U�L���v'N�T�ZI{v�QOV��@�m��q��:��l$'dn$��m�rGHR�	b�
5�;�e�ꨍg���/Emi�eL�5�R^�3J���H]�Gp��keؖ����Sg&��N8�F{=���B�Nz
�PMR�� �C�������6��vj�u��N'd��II�Yf��e�c�6�E�����tP�]�Xԫc�
�]�D1���󣩸��m,�l������C�u�Ӯ_�`���A��z/� j��z)�� 	�Q�PR�!�P���#/����ڪ�%qb�̄kiIA83i쬧dh����M���9+���W��[sgL���^��Κ��x�֮������^nе&�β�� v5��L�g�����ӻu��rDL�YrkU��:��y�K.�Ӳ�����9!w��8���TH�R�й0m�w`�+��Y �w5x��<k[��m݊6�`���zdw�k8+p�&Hxܬ�aّYݛb����ļ�-� `;6�3p͖9�2�^w�{��7������wx�D�,K��sS�,K��=�����=��,K��~�9ı,k��E?"S��&�5$����#��R)�����Kı=�~�q<�bX�'�nv��Kı/�����'�\���{�?�~nNH���Q{���{����>���yı,O~��Ȗ?�2&D�����<�bX����S�,Jr������@l �q�+㔎R�b{��mND�,K��{�O"X�%��}۩Ȗ%����!v'�����_�r��G+{�8�QE)7GND�,K��{�O"X�%��}۩Ȗ%�b{����yı,O~��9H�#��W�ٚ ^�$*�6��Q��V�ř�{iJ$9C�<i���!0�����>�`��sr�5��7���{��s����Kı=�~�q<�bX�'�nv���DȖ%�}����yı,��w�E��Q\�IE��{��7���{�s��> ���
`v'�,N���S�,Kľ}�w��Kİ}ϻu9���,O�~����v]˻wM�78�D�,K��~�9ı,K���<�bX���n�"X�%��{�s��Kı:v���2�˹m����jr%�bX��{��yı,s��ND�,K����Ȗ%����X�f���$)!n튶N.p������yı,s��ND�,Kc���s��Kı=�s��"X�%�|���'�,K���f~�f_0�.]�8�:#�݅�ݞ�J.�9����Mv�n���4�Ϝ���U�J/w�{��%������yı,O~��Ȗ%�b_=�w��ObdK��;��r"9H�#����| ��TQ8��ʱ,K߷;jr%�bX��{��yı,s��ND�,K����Ȕ�#��VݡƓq�q�q.U��ı/�����%�bX>�ݺ��c����Q� �؞��;����%�bX���mND�,K���%�٦n̙�d���O"X�~@A�{��r%�bX�g���O"X�%��۝�9İ?/�؛�����Kı����&�=E:�J/w��oq����{�s��Kı=�s��"X�%�|���'�,K��>���Kı���c�ֶ���mn�;/NK� T��������X�{.��r��0����o�>�ޱ%�s7<ObX�%��w?Z��bX�%���x�D�,K���C�'�2%�b}����yı,O�����wM��ۛ���"X�%�|���'����ș��;��r%�bX�g{�8�D�,K߷;jr'�eL�b}݇��i�&l̗L.��Ȗ%�`���u9ı,O~߻x�D�,K߷;jr%�bX�ϻ��yı,O�7�KLܻfffr��ND�,K߷��'�,K����ڜ�bX�%���x�D�,�b |/���ME𫢎w�<�d)!I
H[�6O�+��VHm��x�D�,K߷;jr%�bX�ϻ��yı,s��ND�,K߷��'�,K��/r�a�e5��e3�*���4$�����=s�$;cզn�G��`��4��e��w��oq��%���x�D�,K��sS�,K����gȖ%�b{��mND�,Jr�nk%��6�|��R9H�X7߻����G"dK�s��yı,O�����Kı/~�w��O�����{���v�=E:��7���2X�'o����%�bX����S�,Kľ}��Ȗ%�`�~�jr%�bX��w��f�72n��s3oȖ%�b{��mND�,K��{�O"X�%�}���Ȗ%���"}�w��yı,O������p�����Ȗ%�b_>�w��Kİ�@ϻ�5<�bX�'����O"X�%��۝�9=�{��Y���~~_��  ��9�OlM�1u]�W۹T�[q;��ûs�n�7NPz�li�V�Ǝ�t����7[	���=�URL�iD�!��'4W���3���{l]��&��n4��v��;$P�r�:��k�Lm.��]�ݘ����>e윚2��ZzcB|]�#&��d愸"��툅�)�SuSvTL�cv��0��֍�^���{����o���u�2�h�{#���p�Z[�<Pu׌tVـ��Ӯ{v:E��5ͳ��ܒ����D�,K��٩Ȗ%�b{�����%�bX����S�,Kľ}��Ȗ%�b}ٽ�Zn��\̦\��S�,K�������Kı=�s��"X�%�|���'�,K��>���O�@ʙ��w�?Y���I�!��m�yı,O�����Kı/�w���%�bX>�ݺ��bX�'�oݼO"X�%���ޓ,�ͳvL��76��Kı/�w���%�bX>�ݺ��bX�'�oݼO"X�%��۝�9ı,K�~�K%�fn̛�2M��'�,K������Kı=�~��yı,O~��Ȗ%�b_>�w��Kı?(�s�Y�l:J�k�n���N+f�nj�^k���[J��ԏ\�v�E13�ow�{�K����׉�Kı=�s��"X�%�|�����Dؖ%�{��59ı,N�O���3]�r���s3oȖ%�b{��mNB���P�El�j�C�Q��ֻȖ%���<�bX����"X�%����oȖ%�bu��-���v�m�\�S�,Kľ}��Ȗ%�`�~�jr%��'�SblN���׉�Kı;�s���Kı=3罳L�3fe��n��<�bX����"X�%����oȖ%�b{��mND�,K��{�O"X�%��f��i�fə��Y���Ȗ%�b{�����%�bX~#�y��O"X�%�}�����%�bX>�ݺ��bX�'�v���,ܑ�G2]�uyy�h�l&M�8��5��<�ɖ{WJgN�'6vb�v�&>�~���bX����S�,Kľ}��Ȗ%�`��v�r%�bX���v�<�cH�#��n�h����AK�g),K��{�O!�9"X?g]ND�,K��^'�,K����Ȝ�g)�r��5��r�l#��_�İ{�v�r%�bX���v�<�c �(�@��b4?�� �T�ObX�����,KĽ��w��Kı/�>�2N��w&�����ND�,� dO~���'�,K�����ND�,K����'�,K��>���Kı<�}�2L�f�Mۺn]�'�,K����ڜ�bX�%�߻�O"X�%�}���Ȗ%�by�{���9H�"�ר6T��NP)RJ8������M<�[�b��5m;;���d��_�f�ۅ�u��jyı,O����'�,K������Kı<����Kı=�s��"X�%��O���3d͙��I����%�bX7߻����r	"{��ڜ�H'���j)"y�jr'��L�bw���IM�6L̹2�ݺ��bX�'�~��Ȗ%�b{��mND�,K����Ȗ%�`��v�r%�bX��ݝ%s6왒l���<�bY�?�����S�,K��w��q<�bX���n�"X��b�� 	'@"*��|��%��x�D�,K���囙���˛d��S�,K��=����%�bX>�ݺ��bX�%���x�D�,K߷;jr%�bX����f��gb���эwk�4f�vV���6����뎸ا��qn��8�.֬�S��~��İ~�����bX�'����O"X�%��۝�?��2%�b}�~��O'���{��?8��o﨧UKE��%�bX����q<�bX�'�nv��Kı=�{��yı,���ND�2�D�=���3]��7n�v�O"X�%��w?Z��bX�'��{�O"X�%�}���Ȗ%�b{�{���%�bX�;{�t�v��-����S�,K?�BD�~��8�D�,K��٩Ȗ%�b_=�w��K��fD����*�R9H�#�����%8�=��yı,���ND�,K��{�O"X�%��۝�9ı,Os߻�O"X�%�UD�N���������z�J�z�)���|�Q��鷚pΣD����O7�+�X<�ke�v.��=8kn`h�2���V��n5�ȳnT���C�;����꧕�!�����'9�.����B�+A�`��&�鶔�X{
��=�W �e�)N2��2۝�Ӕ�-��v�n�l�n]�m�O(�*U���;j�*S�<�-�;�d�UA�EM�[��w&���%�@�;���^V���p�[-<Z�l.�;I��k�n�c)�6��4�����oq��󿻼O"X�%��۝�9ı,Os߻���L�bX7���ND�,K����K�˳d̛M˛�O"X�%��۝�9ı,Os߻�O"X�%�}���Ȗ%�by�{���%�bX��E�4�qq.U��r��Gs߻�O"X�%��}۩Ȗ?�?�lM����8�D�,K��?�ND�)�G)osX�)I�BA����_�r��ϲ�+����K�#�6�&,�V�Z�l7�)#����wn���LY����0;* �Er�T;��F5����n]�xᮚ�a�l�{I�#�S�n՛l�'QS�b�H��ԕ`}׺���elL䏌��ҴQh��J�Y���Oo�w9��B0 :��%�Qq��+���Xv���L���쒜Ҍ���{�`}�۫<�q���ś�`f�V�� N���U���}��^�`b͔������S���R�ȩ
J�>��VWs]����Xwv���V{j�Q5�#�'6h��TۓNe�a&6N(6z!(z�q��p*�:"#n1A�G�b��;�ۦrG�r�Lf�RB�J��.ʪJ���ʑ01f�`b0ԓa��HƛrJ�>��Ձ�^���~�*� ~��z*T 0��e%��"ˁy�4z�e�D�#A�H�L���}|��x�I ��D��� �BH�	,��
@��=���CЄD��Z�g��<4u�C�t3�D1�Lú"z"�O���D ɡ�����x�OA	r,H� @�0��#ӑL��/�+O O�*�|�S�0=b ����~Hj!E���Հ����$�d�s��NrD�R'ԕ`w�����ͺ�>��Ձ��5��������6S3c��#��R&B��0L�S���;�WKRb�i�����
q��Nsh�s.{\��c\�6P��X��ʑ01f�`l+�D�VU���u|`w$|`w*D����`w��Vu��C�P�A
J�>�76g���L�=�`w7m_�Q�3�=J�q�8�8�>���r�<{Vc�V�nՅ(V�nC��wnl��ԁF��d�m)����X�������+�������4��ֆmź'rJ7�ѻ�R݇��{���^+<8�	N7��I+�;��Ձ�^�:����6���b�Z��26H�T�������$��*���U���Ձ�wn��q#t��&�DH�Q�E`j��`fl|`�-�ܩ8��)�pm(���?r�fo�� �{����uX]�vh�V�� N�8�0����~���z�����X! >@
�D���������UR���h{����\+�R�nj�jU��,#8,!l=q���t\#n̴Ёml�ru��"ǆ�ȱn��c��۷M���n0�H�iS�wi�vպzήٟ���p�L��a����˝�o9�$vE��&ņ 9n(�2�OΚ�n�ͥ �u�e�g���Rm���.���Þ�f�Lhmcm���ى7 ����q�fv�e���z��p6��{u�X%��xB+S�ݮtݹe)C�
m90��������sn��_ ;���3�=J�q�2QLY����ʑ0	6S@�I�2A�����sn���u`}׺���幡I��#r9R5'��B���7~Vr�f���X�;V]�oç9�9DjJ�;��V,�L͏�䏌v**Yeخ�M�<��njm4vIYݛb�F��Kβ�yA��V�1qL���&�h�m�?������kbJ#��ń�\n��p`�v{�uwK�9T��o���<�`uw5���tHpp�]_rK`w*D�}�Z�z��ό��
l��(t�nK.�����}�`fl|`�[$'E�UЬ�E��ŒS3c� ̒�ʑz�A�<!?(��H�P�aG�[�g�W=:�����\]����4!��eU%wL���d���H��k�>F�oa*F�r��J�;�۫�%2w+vl�ݫ��j�)��|ҕr!NP����������aXs��}b�(~Z&-��w���u`n�n��[m42"FҎpr+Q9Y�Vc�Vzݫ��s`uK�|�
��W@�遙��#���U����`z���|�ER�JirY�i[p��5�lRr՛sk�Mu;c����:3�j$� N�8�|g�u`}׺����ͺ�;�4)�r�N�IN+��s{
d��ڰ3ڰ;��^�J3�=J�q�2QV,������Y�K3޺�;��V�Y��Q��BA�����T�7�U���]Xu��9�i��*U�r݁�nV�F�nG)���03$|`w*D�ŒS3c� ��aP$��"*U8
��H]�����J�e���a�9���:�M�oX���*����^�`b�)����#�3V�N�D�I��X�5X�k��G�r�L�߶%tZ*ʡ]ZUi�����#�?s�f׼�T�`f�7F� N�8�Xۻ,�Ḿ�X��a)�{�7i�*�+����nK��`z��f�|f����w��I<@�#_��@�A������~z�w�J�v�  [`ۜ�{P6��˓<���sa�6�W`!6	8�V�q�mZ� pץ�����=�݇1v��{�\˷m6S��W4�آq��S�W1��'[m��$��G`'��4�:�����M����u��K��8.A��3vݰ�fdT��mV��[�j���':b��8�1�>�J�!U�����fUh�n�����~O�:{x5�qX�<��{�݉�ۮ`����#�N�v��MqW�O
�8�W' �{��=�~_ =������ �?yX��y����! ��݌͏��H'��`f׼�%����W7+x�	R7#�ӒU�f��v�L��������!_�+i��SnK�{���٥��ͺ���`w5m���T���Ĝ���٣7c� �%�;�"`wd@�vM�]���N4M���rf�jFȩԭgK�H����h�(H��JpJ8ۅ��;0�[�R&�p`l($)c�'L$r��n�ʵO�\���T#��U���K��u~�G���M���E��]02W��%�����IL��`�����V�%����u`b��a�s��=�`j���R�NB��Uv03v>0�[�R&͚X���@��"I�
Hr5(r��Uh��&�^hݕ�=�]kH�r���oۮ�9"���� �{����3vi��͕ ��t�S�b�INnK嘬ݽ6>0�[4��H��Iԉ����K��uf�*���pEH�A�p�5 �*�R!DPu(��E�m���mՁ�9�FD86�i)��ͺ���`|�u�z��.�oŁ�)視���%9�+'����K��k�;��X�v��������u���F:��9th�l$��s#�I�Dܲ�Ol��I��g��ݗ*Ut���)�ٷn����L�5���%D�>ܚX͏�Y��[%?}Ĉ���WB����
�`l�|`j͔���)�ٳK�no�T����NIV.�$����$�w���& M�qO���X�����AG$�*&�>Y�L	�p`f�|`E�Sej	|�WQǧlJk��m৶8��U0�\�M[`Ȍd�楍mR��-?m�?�ɖs��[�K��ݫ�='���m(�ns6�����`|�u��4�3Jɴ���	�I*�ՒS�d�ݸ03%���ۈ+���)��&�vWw]���K�٥������t�XF�b�L�����2��_`9�u`vz�X�K(����� S�� 8��x��'�)8�3��}`1>�(!�Z>@3U�))������@�  ,�R)�Q�ΐiH��ꦀ�C�)߾q�8{⧤��?E�}D��=W������!�R@�FH�bh$Q�5
���!��q58P@��yQ�R|Cρ�8����	�Ë!��{>�ۙ����fm� ���          �  &�RFJI�D�k[&����U)9;u�ȫ��h�V��FN�.��lZ���"k[��@�Z(j��^e�Ts�6�m�t��06��D�&H��V[/Sk����Z��۠��6)&�� {t�&Gj��n]���]Q�h���oh�c�����&3A��e�v��+U�M�n�$bv�(R\���Ny v�j�H���-���N�';����r9j���;����xx�޶��T��y>���LK�I�]��4�v���	�%�X��i-�~�x�����ۗmuٖ��!�=qa�ے�N�Ct�#�Cc��յ$�Mf݌��ʩu���j���P��J[H5b�9��7&Eؗ7/�����3�έP�쫔�q����n��rf��@���vw6�H��:�U��MFx�u���!s��;u�k��F��J���j8D+�o+��iI6[%����T���;4����"���2Bt��T�gA*���Yx0�Qm�siB�&\�+�^���s]{f������n�q5 �eXV��UYsg�n��͋�OR�0\��GB]�彩�]����];z��'nHn�M�I9�19V�):���W��ʨ�R�&v��W�v�t�d�UOk�B�,m�3m�"�H����E����������3K3���vܷ	�ݕٸn�U@����l�<]+����6�۳�v^zb��Mu����;	u/.��v����0�*�4�c�&N`�x�݁��6��We���㏓}Zw.Wi2J�M�Ǝt�k�p�<��Ā��K�"	ӱ�&E�vŤ��sP�x����H8��#AJl��S S�&��Ӱ�Xح������d��d�k�+�0TQN1Õ+� ��-H瀕[���DHNz�[�XȏFe�᛹m����ɹ%�P����i�>����T& �����_Pz
u��hp@���T�;��׿?n����o� �i�:�w:v���C�ó�6���8-L���$Q�8k��A�ĜE�3�@u2��m֍�&:[V̀a�+ԙ
��X��6��c�N�8�Ƹ��uayX֣��Z��eXNێleZ�Ӷ�zh�RI,K U6�/E&sNs@����2Sd�m�l���ŀ�!��s�ش�y�2Z�b�v����m�P��o�wu�x߫�]v+�l��h�p���j6T�x.1�&�Ȏcb�9��:w�Zڵ	U��d��ŒSn�#sx���D��SQ�X�vX]�v�M,�f���OD� ��S����,��v���Kw����03����!����v�M,�0"�)��$�sh�Į�EYT��UV03v>0"�)�ղSn�,X�hF�5Q��R1�ʏ��Ӯ��m��T���p����su�rλ��usm��	]��IL���v�������2jN��� �q�,�w��!���TY��"��Jr!J��|�`u�ڰ��{
""F�Ǒaq�2TN;۳Ł����&Il����W�^��Z*젻(J��w�|�|�0o�lY%0�����:���)EJ�95��ov[�d�ޤ��p��K28w�$J�ߒ��3Go
�֎Z˷Ok�n�8��Oj�)�����{`L���z�u6���In��ޤ��p��K�8{�}�I$�ޒ�In���d�D�r����H̚K�W8�K3���I,����]}�}��mm/s�DD84ۍ&�V�K7}�}���{��`'��"���<��_|�K�ۅ���^�d��$�I/��I%$�i$�/b�W��{�v4�Y�����%���6�SMMI%���f�ޤ���9��T��i$��w��I%6]�����#b�b�������w`��u�J@�6z&G%�lj��d���[J�"�Eծ�$���i$��w��I%6]�I.�f��I-OM�%)9
B��K�'y���URK��m$�T���I%7n�K�noaR�NB9%}�I%�.�I.��]�I)���IfG�$�E4U!�*I(d�KI%�����$�#����G�%_s��s�����}=v�If����#Q5�$���[�p��_n��I!M�m$�kvWz�YEmA+���5qnw,5 \�!���]Ӫ��q&�7,c2�''�3dVI�| ~��;��$�6U��]��]�I)���Il4���)�I��J�����UR�K*OWz�^��������;Ԓ�6�ӡ�)��6���I|�5��In�-/W9M��������-$�n���6�
�T_-]�z�[%�$�r8w�$-�r�Iu�5��I%��RR����%:���Iw#�z�B�*�I,��]�Il����
'� ĝ?Ng�����ڪU�^�^���u��n�p�!n�� �B6��ř]�n����h�1-��lǚ뀵gzɳ�[��Vě:�/W&mm�MgDi�_>}	l[W5���[r͂�v5��=j���I��,�Y�;���9õ�7hʰc�e� ��0v�e���QVŌS
�. ��N����s�V�Ͳ*��l�C&�H#�p�i.
�q/���}X�mt�MȇJ*Cc����薟�~�>��b�iM��-����zs��ذ7�ۮ������� c�?��� ����Ԓ�6$�r8w�$lW�\����$RQ#��_s_�$��ˢ�I}ݽ>�$���/�r�iny{�	L���RU���I/{��4�]��ޤ�RK��K����K���q%��n9�ZI.�p�RHRJ��K+6Wz���}�W����K|x�Rd��$�6���$-�q���͕ޤ��o�I%܎�InԤvO���n,ٸ���m��^z�����]�Cg��v�!M�� ��{3r&���$��͕ޤ����K�;Ԓ�����wR_m�(4�QH��$�6�/�������fbX��w�$)=V�Ief����RR����H�p-$���ӽI!M�m/�����z�Ԓ��`�b٪�aR�NS�H������`uw5�ܚXwf��r�����L�P'wLY���������;6[ ����pˋSe	8�IEQ�^ͱj��6�s�YBn��tr��P��RByUt��ۃ�.�e�1f�~�9�9Ď�ȯ[ID84ێ)!`w=<Xf�`b͔��ۃa�T]�Ң���X�,�qՉTB���B� �j1�E  *0�*$1P"A1#a�?� �dcGt_}����I<̚X�5!ӡ�)��6�vWs[sn�0����03��I��UЬ�E���076���K��l�Ws]���n�Q@$T�T��*�'�Z9k6,��*�I�$;��4:��ٴrl��ݸ#9
t�H4�`}ݚX,�vWs_��_ ����ž��T����&�`uM��ś)���r\�"7�J&�9��vWs]���K�����n�3sm��d�D�r���b���`w7�X;X}v �B�"�D��#�vo��j�~�N���C�M��r�٥�}�����k�>̚X�UU[��>Jr:i�&�9�}�m��k�&���OOYv��퍒��㧜�bR�$�'Lp���;�����2i`}�۫7v�:t8��Sj]01f�`wv���H��ܭ��#=�$�#n1A�J�G`w�<Xwv��μ�`uw5��͢��r�J�s\,��Ձ��s`}=n�6���]��:�����D���I*�μ�`jI.�n��n>i`w��Xd-�I"�D��e7��3��������+��YN��R��N ��ڧ�.��j��ڵh�Θ�������t8i�ntVQ�Ie�v�&m�#�m���K����D�-
��+�F�Fˍ�C�k�5�������:n�bs0�ؽ��좬�1�R0��`S�
��/e��ٌ�,;pyݳg1@�䫁�9^e�m	�lZx�ݵ����r���c!)A����*r�8��Y������k���+�ö�g���cTg��L�r,����7�4�;�ۯ�+�_ �=�7���)�R�Q�RN;f��sc�f��Vl�vqF�Q6�9V�ͺ�7��V˹�����X�Զ�$�'�J9V�)�{�;8���v�6{�~V�ٴ:t8��)�*��w5���V�ͺ�7��V�^�ZFH�H��1X�<�`�p
ClF.�]`B��ǫ��t�/c�j��q�2TR?���P��u`}�*k��1a�RR���JT�RU���_bȅ�����7{��;�Vz�Ձ���I:*TI�qI#�;�۫�$�d��Y����ʯ���W.��]_Y%03$|`b͔�̛u`n����T�D�nq)����X���k�37mXO[���A�p�K��8�bN������[��Z^n��K8ݎ��re�:88�t��3dVu7}������X�v���֨J�׶����%8	>6G`gsn�$|����6����k�I���t�r��9Vg��Տ���P�K!D^CP�ш�`E �� ��	�^4�E� �z�8 z����=R$�M�gġ!X�ƊU H�EJ^$�[m+@�X��%q},0W<���@|�|�>��
$�@5R��4 �}HA���iR1�%�a�n�B+"�6 ���G�����,@�0��#<"`!�S�Ak��Q(0J*���,A����$cp�Fi `��> "w�ϏI��\!$"��|�X��P��0=��HF63�=uS�_�A ��E��z�>	����O����g_��|�(���S�Q'������ʪ����u`g�}E��q�2TN;���ߕ���j���a��S��ڰ5i����r�J�jJ�:���͏�������K��3�un��"�fp5h�r��W:��Px˷k�N;N
Q!Q:*TI�8�����۫��u`|��؈��}!��j�4zj��%(���"9V˻�����VWs]����X��)�#Q5�%#�3$|`b͔�̑�ՒS�>Q��C�M�ڎU����`w��^�r�A�������U����->UW:�~ݫ��o�"Jp|l��ܑ�ՒS&��,�L��%�����㤑5���zͱHK�c&bاqE�vz�<�̦�ڋ�͉nˣ������`u�`v{��"!/�nڰ3����q�2TN;��u~�s�5l�0&�ό����"��%hr�J��J�1f���۫���`nf�X,µ:*TIʄ�1��쏌���v>01f�`٨�U}���%9H�U����73n���{�u`:���s���ԛ��I$�I@��a-�k�h:�ڛ�����&��]/Y�i2�򅶀�[$,@n��@-�+t�)�"e{m�m ���@�9R*#g�\׳��%�mN�ٻ4��,�;c�.�������|s����na�v�	�EX�Y�-�GH�ʴWX��[f�Q���-���V"���:�d^��]H�nz
0����,���q�S�QC�_Ab���Y<͛K�Ƹ�:�	3o;p9�v��A�� -p^AYp������HB��O�m��?���,�L	�>>�[�S'�^i%��n9�`uw5��۫���`>�z�D(S&���9�\	�����`{g�Y%0&�|`b͔��D��F��S�U����73n���{�u`wkt,�ӌpi����ݏ�Y��$|`ud��ݗ�i��(�3'\�qp�-�m��k�'h�5�Dsn�ݒ%�gӫn5��5J��,�L	�Y%0&�|`uf��R�NT��G`own����7�����DB읟���o�X���]�t�=J*nR#��Y�;{.Y��v>0$$uE�]��]�J�v>01f�`L��ՒU��r���q{�"!���r7+�1f���ڰ>��V�v�I%��ٞJ����`v����<\�:kf�*͕��4��Nn�NY��sc�\���]��w�|`ud����񁙱�$.
�PQ�CdT�`|�����VWs]���uuU�Uݭв6�iA�J���76{�Ֆ���.�%��.%j!qED%��}j����X8cB�9\���h����`fl|`I��ՒSV��V�EJ�9R(F9����ՒS)%01f�`E� ���^�wG��8}iK�c@f�f��l��{�Ӆ��y�x���rY��w�o������l�,�L	6>0$�5ʾQ���B����5�]�v�mՁ���3��lH�pi�i�`uw%0$�����)��L	(�\E�*�*��*�l|`ud���l�S@����U?
���W�*���;wjxN�nP�8�XO[��-�=���ǵ`7�Ձު���.��x��ո���<5�j��d�kX����&8�on�M�v��!du��J�01f�`I#纃�����RDr�DI$qX]�v��Ձ���7^�r�Ď��y:*TIʑC�W9V����:�T)��{6g�$�Y����˳4�sNI�@V�[=Lz����͔��G��F�W�A�(��4�7^j�>]�v�mՁ��k�9YUڮ5YCM�I$�I ��\�D�g�a��y�3�@��'_����;�۷)�����-�z6���a;FZ��A�;f�+�kK�1�����ŉN�f�<�="�N����<�,IYب#�����T�f��̰��m�=Ѽ�H)N��d�t��7`���n[v{n�u7y:)[q�r���]��v���y7\v�5������'P*�(��y�칛���MC-��ɩ�����3l��x�����[^i�:)�I��H%N6パh�ߝ����՛)�%H�>^����.�V	W�E]������͔���L����*h�8%�0��U���k�7jD��l|`I#�'6p�IQIYJ�Wt���L����>0:�e01a�E%��JR�8�>�mՁ�G�Vl��"`E���]�}VU)�5���p�$��wi��f)v7B�z��'\g�.*��GO��NT��%|��]X,�L	*D��l|`b"�8��ˤu�Y��$�_~�s���E�x��G@H��������^I?}�����ͺ�7um�r����ӎ���&sc�M����L����D84ێ�`}�۫w6���w5��uX��"Jp|lrJ�5�j��{��鹰>�;V�%��S���Ɲ�Ù��Yz�:��Ae��WNkdܖ��9�BV6�.\�y�M�ts7:-���"`w6>0$�񁓛(�	�(4�H�׺���u`n��X.��RQ9
��G"�o$�{�xrI���9><Ө� �(+�IB��D�v��6�f���	��D��#q���ݺ�>]�v��V�ɥ����>o#C��Dr��qՀ�76��2�m�V�%-�V�fsZN���5$�"��š�sj�=e�����۴����aט�L��g��ޯy0;�p`I#��6Sf����n89��riu�s����V˹���{���fh�S���c���$����L��s�Ĥ�������ʚ'N	G(T�9V˹��w���I<����U� D(�K~	���P4P"(����U����Ui&4��!�X�u0;�p`I#� �l��M'�%¿N�T��m�i�-�횺aɍ�U�٧80�p�r)J�E_�{�`6ݫ ����Hn���-�iTqZUwj˪Wi�$�����T���^j�:�ݧI�yNR#�`w6�T��ܭ��$��	"�QU�l�8�'%���=�`w���۫ �se��5-��!���pr+�s`V���t� ̬ɰ?J!%�`
�������
� P�@U��W��W���UQE"
	 � Ȋ �(�"( ���1"�1b� � �(� � 
���
���(
��Z �*� (
�� �*����� 
���(
�� �*��W�W���e5�%���0fE��?���������� �h5���_fF�vԁJ�n��k��0���A!.f��n�*o�  :�`�(($J�m(��*J���4�fTBMd�R
P��B@�    �{��z�0�P�x�浻|m�;�v�&������������z��l�uWc�Ϡ������R\���:\�� o{�l�kz���2�>���P4(�3t|X$=47��`���i�[z�t�a���AN���"�ޥ���� ����^��á�{��;� ��e�� {� =�� ����_ �����2�H��3����[=�u��\-��׏��\q罇\��
t���t��{B����ѻ@��������U^�-��F��{����ѐ.í�;����݇B�gU��$=� -�E�z*�J�Š*�R�;��%kA�:4s�zKB���n�C6(��T�< h�h�d(�`���6���E2hFF���x6��=���w��.h��H�ϔDa�4ģ�(7 Dmtg[��4�ׅm�sr9��    0�JR���@�h���R��#L �2 ��F�Ob�R�<�SC544�����@b��5P%( �     �&��4I�2��
yM� ==l��
���5R��&�   � ��}'�����55�_����������C���(� ��"�
��z�����6�g�.����7�g��� ��)
�����*�)���H��
F&����¾����8��~��|�wwwwwwwwwwwwwwwwwwn����wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww��{������������������������{����������������������������������������������������������������������������9�swwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwswF�{���{����{������U� �� |� |�>[m� ���A���|��|����� � ϖ��|�o���o�o�|� g�6�>[l>X-��,� >@� ϐ>@|�|�پA� ϐo�|�>@ϖ�1��|��7��A��-�l���m� >Xo��>@|�>A��6�>X>@|����1�_�{���{_ȁ������Re�/_G�OϤ��}nL�@�R��CPn����*M��tct8��j�4aƒ���5h+"´��H� �Y�D d.�l�	 3y"�Έ��f$�l(�w���oL�7CF�K$	�˽oN���d���N�F�֫X��A��xp2h�e��E�f#\-�kZ��5T���XHs��5�Z����7�̰�]��Bb���G��wX����T���Hro�.F�sW(��)�B� M���rj��׏Dq��T&��4�y��<��5���+!f�n$x-�ݑ'0`�! @B.�\�5��us:��6�h����jG��Y�?IF!K*B42c����V�7P�D��ٔ�"E�D�
#I�,YI�\B�&)��D�E߯�Ny�{��iǚ焽������-�=6�v�phA�0h ���	�8g;ս�00�5����lR1��S�����~9}�l�<�ǞK\e`��0n;c4�r���$���I!F�2���;|�c���KW<�o���;h�;yI���V�ц¯��Y�VR	I����߻Oe����;'H�kY��i(�	"��!D0d���3��L�'�sF�����'E��y����zj)���jvՋ--b�2X�R*~y\����+\ȼX$K`H�$	K(DÂ�5Mk:)�ȱ�ăg%��7����7��sǬ��v����O�[ŕ.x�[E����[����eӢ׿O"f�B�N��B���k�M&�y�T�r�,Tͭ��Sw	D�r۵��k*�5ӿ>�>Ǟ���Yf̄��
�b�gtj�A0a�ƫ�B��5"���$M�a��,2�д�z��� 1��Y�j�߾{�Ǻ�k��$�\�1C.�X�^&�;���G	�R�n*��yw}%�
��c-��q�U�)�	e�����bS

��֕���/�כ��%��ɖ��[�z��g�Ş�tI�[Y-��Y�kxE:iґ8�.޵��VG-kp��-�n���s�Kq�uo��Τ�	���רK��0�nNwK
ˌv�!�qu����C���-B2kn]n�b�I7o6z�g	�hTx���Ӑ�4(�%r��dռ�m--���
�ݗi�ʋ�BB�2b�JEhu�![���D��x3�u����XY	�����;ı�<}��J���dV9az��ˊp�q*h�$�%Xe � ��.�y��tL��&]�Z��{�X��IS�A�r�.^r�"e��Ύ�*�|�țC&H0#�����˷Mׄ��>X�6�me�`��[�뷈���V���['Iy�����9��i��5[9�ą�afGÚ�ܙ�2����#�{-�v&j��'�2�E y�`�@(��
������A�],ƺso	�|ui�h���L@��pl��3�\�pu<�m�]����  s��}HS��+��"L�k;dt�<��{ζL�D�0Jˀ�*�J�]t������K$�Q���UB�d�M���+���X���BOu�9^�.6�H\rg���'�FM 9�d9aa.�8��I�BC���Y�ht�R�=w�]����b�!�j�SJ�#�ޱ.��F��|�ՅYfd,��9yR��5�ۺ���뗷�~�"[�����%^�V�X�+�h�F&��$' Csq͢� �	L��%���+"<�4p�޵�V1zt�
!�M�k�g[�߯~��[Q&��ӳ�i;��<���v�zz8�����$%�̪���$����8�V��h��X����=>�w�O{#��[���莤�z���عs'&t�Nx����^��{����bJ����-�c��B�Љ���������Ͻ����JE�h�n����ⵑm'".B���$�:S��-q'<z9���IP�$)�#��%���#D8�3�H�ai�B��Vu�l��h5��pC\�2.7ݛ�ř�ьqe&y[����
�
�oI�ͅ�Y�S��C�}X��mʨݷ��춖Ы7)2{[�hc+#)�P��q%2���f�NL���Haa"\
&\!�f�h�mX��j�
�P�&��p�&4Ƣ%#0�cPv���m��z��nO4;[��'mz�ϭM�"� җ}�S;�0�B�4®�WLJ�%�9txK1/1%��ǅ�F��%�W�7#�C�9ڭ�K�)��y���t��{��z�t���NӲ��߷=���<�޴��	
��g0.�4� ���1�)�wk%�I��	o4������{#����r�n�H@!�՚濾��x[��%��^��BR�a��G���f>�f0z�h"��n2�p��%BV[�NK!!���E������S֖�����ſ7��v����,�����F���B8L���f��+&�XGm�囊7>��+nX������;/.M^<ے۝ێ�<[v��.N.�R�s�t��%s�ۼ����tZ9n�AӁQ�H6��H�4�	Q8p�B��aMg`����Ä%�s�1� PD�$��Y;˕[�wgm���'r	An�u��\-�Q��Gj��c	6��4�YCR�X1��1x��-��dY�8�e3�����=���t�Մ��9��Vf�����9��b�v���홺ܷE�#�@ݵ�6-ls�r��ί �l������=��='Ը��Z
�b�0hChT��-��.��2��F��$�g�,v�[nڴ�B��P�J�)�KMUi��:SL�b���UU�v�����O�����(���J��I�w�������7~w��o���        @-�  �  m-� ����  ~�z                                                                             =@                                               �UR� K�΁�\�7G�*��H�H���-��ej�$s�X���ѫjy@kH����]�9n�o<� h�vK[kk/lP�1��49f)PR«Pqm��vaz�t��,9j�	���u�B�oĺ�cj��*�';@UT�sj��7Jgyn��
�Z�]�%�s*ͷ`qi�[@ m�TUPs�����$�U -�h[@6� J�  �pm�ݻ`�iת1V5��	����XתN  �F�Om��Օ�U�8��d�m�6�p�sm�  2����	jD���m��  8S�sq��  ݖ� ��h� I�wv�0ni��Ui^�6�[m��6Ѯ�H � �-��0=$=� ��  �l[B�vڕ��8�`mޠ�mnk2�k[���մh�� l�L�۶�!���$�M�$$ p��0v�.�H2�V�u�vҭU@N�j��^���%yU(-����ng��Fթ���Qsgb[m6 �6��v�ko\�-����Hsmd�~�۟�@�7P=�S�g���Ȝ<�mq��u-'\I�s�%�w-�]s�B�BͶm�U�6���V� �m0�Ͷ]�cB�6��v�5�\ H�6�ְ9���J��
�5�*��j��k ��H ��ZRYVBj�4t[6�As]0n�vn(��fB��bĺ\p���i��}���]$�)��d�Un� ږ�rr군 �u�ij-�icdI�N�
[>InI`6��W<уv��8Hŋki���bڹ/��od86���h�`N�A�Cy,e�s���[ +UJ���b���[4*�@U,���6�m"� �`��>e���A[�W*�M���c����V�-  ��j�h�om�+m�m�$m�9bl��-�9�� $  v���  m  �  v�ꔅxx
�Au@  6�m�H]R��FD&�
�*� ;\�if�Z[� m��Ά�@��HO�{�Fʫ,UU�Z���h1��b8AU����R餓8�  � �;!�R��U*�@@mn�6�օ*�;Z�� ���� ���mUb�r�.�
|sU;����p�5�qkd��t�Ig*lym���t�� �~>��v�g��)�r06��"喒_#li/�$�  m���m � 6��[B@9��/5�M�jJS[��(-6[dHI�m��8΂յ�M%��Um
�0�A�;M��٫vp�j�����^�����*�*F���B���mMiB�����u����a��NPRř��.�Ye�a+\8�ݖ�m�$�5��Ammm����[N [@���`6ۀI"Kz�� z�6ִt� �s��k*3�wo�p���ӯM�yf������  m�N���V�m�2!5m[s���8@�
�9&�Ց����M�m��jQh��0&�M�94�L�豇p�5a�ckhd���9���9=1��Z��k��^��k��S��t]e�n�f���`��Y% �l�i-�����V�G �+��Ѯ�   �6�,V�zy�t+�jg�i��#,�o`Vn%�vw=uc=pun����ϱ�\"n��`)II�ն��v�j�8%瞭�m��T'[A��v� ���d���$'�ؖ�
�J�ԝ�Ju�Qd�Y���� $m�z:�c�/�?bv���^	}���L)��b�����L�y�r�"��c�Z��9�Pi������ �n��Ҧ�o],TuY�k�'��r=����V��&��ph���r+ڟ;!ۜ]�b�hZ�ͱŴUX 6�� H�l�ձ�<b⪪[Rs�l�[p��a���z�$ �U`ASIl��Uj�[N�'\�]�T;clWa�6.^�Z�i�타m[淴K|6���z��ԖM;` l$`*m��r5������o4�IZڎ��`(��ѱ�{g�D�l#����ې�r��J�:s5J����I�[p l�69��l�
�"��˰�3WmS�����|N`%eUn�U���Al��E�HH�4�� �k�+i6Sg���֜�J˝y:\��$^�m�{7��v�M�x�m �m���M��R��e�Z�U�	�j��R6�G�� h 6�� �`��*� ��gM�r��3K��A������   N ���l-s-e!%�pKh H R��h�$C��+h�4�b��jU���"Z��g�YV�3I� H�Mn������ ��	����F�r�V^ڮ���S��jڗvv`*�kR>T
U8r���쳒�5�T�-[���m���l����@l  � Uprw
���g��j�� m�  
T�6Z�$��ɬ��:��K,)r��K�������V�MV��탅	���P�K�� �[j� ��6�B\	C� �ʁu��6*�]���+��d�U;!�µI�Ӧov�� �d�Z������' �V$`4Q�m�I��-��\�+`m��T�WW@J�WU*V�Jt&���ڀ�
�*����A�Zڪ��I�rJ�*�UUPHH q�  l ]j�#)B��j��I7n�*A��n  �d�� ��j�;vZ��T��=��K�t��T\�,;(�f���I�  �6�-�m�h� �6�2 [B �ml��ے�8 	 6�6�`��K@�iLH����m�a���'�ۢж��m:C��Am�e� +c4�Rt�m��*y���M��pm��5@iz텚� u�2^�@ a�7]��  	lX����]ܕE]�Z�b�{�1UD���S��
�?{������2_Ş=���S�s��&��INi$H�MmN����WJt뢺:�-�궜��Vӕ�N�Y�:��wC�S)�T�͸CB�8A�8B����$�)%)l�R��%)l�R��%)l�R��%)i%)I)JIJRJR�R������$�)%)I)JIJRJR�R������$�)%)I)JIJRJR�R������$�)%)I)JIJRJR�R������$�)%)I)J)MJRJSR�I)Kd���I)Kd�����=�m�ܨ}�	Jz XP�5���*�,�X% �j�KV�	�t�����%6!�9EU�X���6�4`�uG	�����8X��I��,P�&1��&h�M(䊊�&��A �Z��M�V��Ңp��A�jE؏/�lE�8[��D(��r��'(h�h���'��UN�67�:���` #�E��iW<Cii��@q��*h�,8EH���M�]��8�v���i@,S16��
���)�� 8�: -p�]�ڡ�PX�F	�G@f�(�*�"��6N�)l�@�6�Ǫ�8�BQ(]� ФS�W"�#��' CgC+`��0�����ZF�ɢ!�Cn�U(d��� &�m�E@,@��!A!�tlL�� e�� ��(��mD�Ŵ";�
T:q�!�b!������//����r��ܼ��//�����^U�^U�^U�^U�^U�^U�^U�^U�^U�^U�^U�^U�^U�^U�^U�^U�^T6]��m�ۻ1�1�S1�1�S�� s����9ɤ��<�oꪫ��l���I$�I$��~����9�rI'�$������ m��8E��c���;7m���Æ�v�,0=�����.���ʓRBR��YI K��
r�C��x����Oc�x��9����.��v/}�UU���dn�l�               m�         �z�#n;�LLY�k t�jғx籸.i�.���p,
��1��pl:�� �<u�д�b�/WʛN8�v��T�u�m+���.��`nv�Rq�ڶk�@ڸ�L�2��2ݬK�wk]=��
��-�S3� Z�a��p���O\9�CJMTi��Qه`��v'K%:u���ZAde��5Ԣ��e�#6�ibVXژ3�&tUT��aic�rkq�\*��u��[�bb۞��b�Xkj1�V7g1͸���y� -+�J��'`"^�scNVX[%��������8p�PjF;yö��b�*�yV@��6��7dF8���f'�㷋x�����;)�(��Uh��VI텪Ս��3���MΔ'W�z�ݟd��r�Bq��<��`�,b�E��⺺.��V�ɛ�1$�Z�D���A���Kv&Z��2g���cs�	�9;LcKSj�p��Δ,;Zݑ��`+v+��gWfZ�ˡ=�3��V���٩*UK�[�[t��
�L�g�.z�2������5���v�A(�d4���4�<�si�]K�m���*�v��ԥ���q�6NSQ�nd� �/R��k4���GflY�s>Yr��e�ԸU^&�u:��@0�#���4�x ���[Qx�i�x0C*&#��P,R���rs�-����ʪ����l %k-s����H7X���sn�¶F���3�.]�ΘA�u��ks�[��um3��á�(�Ƚ��-�B^�)[z�'j�^���N4�s]�Sg��$��r5k��s��5�kM�)eH[�� �IԈ�Qp4�X��oX�1��!���������M�w̶N��!C�{d$��'�<�����'�(I�a���Ќ�3�M砗U�T���B���KT��HI�YbA8�q&�'��BOo$$�rBOoT�w�
xJQ� J�Nc�\$��R��`���\�vv �E	��	7�!���A	/��'Wq�I�U
�:2,��&X3-��Z<n%��<�5ɘ6Kf�2�o
\
���'7�BO/ ��ߤ<K�2BN ot����̓\�|h����!��L�Y�n�
`%�-/� ���2BHݼ�	7�$��X��cqA�M��I�fs��͂����!$����$(�8I��< 7���A	ʠ�=�I�����im&�&+�pBM�A	=�����8�� y=�tJ.�jʓFPR!��bP������f�Ѻ�-RM��G^�-#w3�$��w���^��Λ1�(�L��8I��9�OVb��^oS�;�� y��f��]���(�,��ѐ#�s\՗$Ѯ��7f�<d$�N�I��!'��!'��o���]퇟| ��t�z��HI�䄞���:��$�RLF�n��k�67�K���2ps��}��厉�M~17������	��$���N�Ld��
.p�wvN}Tټ�`�V���<��@�߱�Y��&�z�~A��|W����n�s�DZQQ�$I��M��"G��w�$%�CE @���`VU-�`�]kJz�0(Teo6BNe��&�`����}U@^>���6q�Q-d�W�\bc<�*��㳳�qYN[�4��sސ��Ü�&�A��M�=��������r��<��;��$���BN�ɕTEc�lE$�&'I9����IĎ�Ič��	=X��r4bn&8I���'���o6I�rRGz�&2$$(��N��>��������v<������t�L���U�   R��[�v�uC�]1�;JB�nb�Z�\��m+���:6�Eq�nce�xN5�$��:���|8�s�W��i���{<���7F�q-�V���Y9��ۇ��X���6���\j���qc�[������8�c���j����8́��tm��`�%75Ԣ���yYU�zI��!'��'s$$��(��68JWsH�S�y���d$����_��#A-gP>�@��T��!'�zD%��7��	F�G�|){��I�l���I�BM٭�)&ˍ���!'��!'�2BO73�$� ,I9���v���5�Mte�!��jݷ$�8��Pa�/ww,4���u:�������υq��!'���#��Lp�~%�E��W8�'D��.���&��A%w ��
�ȼca��)��O��	<�BO}pB��䄝�+j�
N�J���{��'��	>ː���G5���ě$��F�s9	+{���OsL�����E	�d ��Ń���^cPvpl`�Y�B襱���*����H�섞^�	=ۘxI�#boi(�D8��N=�s�PH��A	7��1+��I�5��m��o����	=˂56�Y ���&I����	:��b �LNorI�d���.g=͂z�X��1�ovBNeȒ<��{��$�}�Sh�CiYZ���
{W@a���9���ܯM�auz��P:�� w��@��Z��l��L,D@d� �l�$orI�l��w��+d;�<�F�2�	;{$�2{���d$��A	�z��`P�+�Rד�D�ᐓ��!9w�����T]+�c���P��(ˆ'�Ow$$��I�ـ�Ow$�D�v�I�eɱ�hE�2ipYm���ۂ�`LO��yn��7�K�o+��e�	=�u#��q�4�L����&�`�H�i���n�{��x�X�h��q�ln�I��	9����'3 ���2�Ȑ�Y��Gwd$�6	ď^A	=ܐ��75�Jp���$����>S��2�gmc�KT �>t��    ĭ"��t���R:yI���Z2�����b#��1���5Ɩ$ ��.��.���&:�G\ÛI����:�g�����)캊�5Ԉ��5�1�Z/��m���ɘK.‥;t����v�<sn6��3	�w�N�F�]P�]�$(���M��a���^��Z^@�w^m6WQո+:!������P<��ި{� ��.��F	Pp�{�δo2BL�o	<�A	7gL-�J2Ï��ݐ���!'�pBO;��r�j�y$���|$�6I��\$�rB@��$��i��	���&��՘�&���>b�x{Ү��b�p��J˹�6�'Fɽ�A�b4SH5��Q��M��	9ې���[ꮲvd�|F�Q��$�I�U�e���km��a��rro��!��щ��7��0� j��<܂o�$�rBN���%��
��� y� w��/nBM��4TD�Pp��s���߾�}�ן1�v_}�#*��%z6BM�x�$��A	9�����X�$���ڦ��k]k,���2�F3�
4nn���Ϯ����X�$u�HI���~�!'��o��b/�F̍���!&������	� ����)#���J2bpp��������O��>>@  �I'��9�$�I9��������I'�j�0*!*R�a�ú�8�B�&	0I ���>�>����ܛ��h��}*׌�E�L�axo)`�9��L��a$a1(Bܓn�3�'&ݨl[��$�NaL�j�HU����ǥ��t�=������?S�eC�)��X�A0����H�g :X%D��6�!���R� C� �B�\A]�7�7��署�+X�.�X�M��n.�
�y���O�􄟻���~���T���P���6�B"t@99�H�퐟G��V{�$�=m�O~������w���`�$�^h���`���f%x���0s��]�����,�e������z��z?d���U�|~R/������z���&�~
~��g��	?w�}����|*�6���IB6�;��r�L^����>�mdny"���x��b|'�  Ͼ�\��`��.��W%�RC)pAdC�R4R��m��{qZr�P ���N)�$~\G��#��#���j�߿U  ��Z�N�HI�m�~�xu�Vҫt&�i��%n8Z͐-!�m �ڵ�^m��A@N��I	�>K������NwϾ����'!�C�4J�H8ZW��}�
���$��'�v	���		���1�			H9�M� >��9�#�����}�$��������9)I�}������B	���^�M�{	?w�?7�G>H�x�'��_��]�}��c�9<'�x��}�	]Ҫ���  :E���L���/mM��6��a��H.�0!.;7h���dףh��]�n���@)�^n�R��sș�i�WBt\`�B ��.���t���\p�6sN
��Z(^.�^��q��-����Y�e06ؔ��rN�׮�\L������˭҉0�� z��X��Dn���Ֆ�Ͼ�=J�I���|8�V�D���a��	=�f���,z"|�|�Iڪ�o9�i��5�
n��'�}$�^}��� I��I��$��?R2���� ?O~
��ߦq��&���UT��$��1k1FȸI��HI��~({��?�a�{��@?}��O�����G�qVM����ˌ�N�o����X8�!DHJNY ��HI�a�{���@~�UW	�ߤ$��#%7�"�$��c♆=0"� �� ���;.I���o�I���!������`��'�>\�$��w9�ا���.�<��$��J�2$e&xO� U������	?c�z����T$����I@�1�􄟾�88I���I��HOW�s�����`�݉���@��[��]k�d�`�-����{���7.<$���$�_T%.~���D�BOꪡUZ��D�2�'Q_j�~o{ܚ�'���;�?��l��1k*F�m���HI˹���hRL�KliL�Mk�$��9W$�Cq�&%'/���������a�mr�'˿r}y%���%N}�2O�'Ǚ�&U|�g2O��ܝ�}�>���WD�SAA08ͫ]l5�4(�bWFjY�Q���RaqF�e$���^HI���﫬���'�ii�5%5�Ļ��}�~��!'���I���=��!�ퟘk����c�'�߷������UU7��(I����}��2�PF��>� P���t2N/j����.��NB�V8m,x43��T$� }��2���_b�_|7��Z8�󓋍}�2O߀��KnI$�õ��]t��K�Ɏ�����4������O�Gε�%e��?�s.g?�c��d�P�|G�~1� a)	9�M���*3��2N��|1.���mP���2Sk���$��2OU�B���9��	<����p��#xC+J�����Z��{�!&�r���$�f�5����I��Iԁ���}��3����j���$�L�j��"W��    ��:��jmc��B+Q�q�X��nLfm�q<�YxՄ����e۔z���XVR�X�̖�5p�\��5�]�f��� �@�f-U�8���^���h��tk
�����m��r��mh��Mv�Vm^w�O��z���LgV�XJі�2�MZ����'H�c=���+���E�Qy-��$�qu��d��HI��ϙmA���}�O�W�6qY�	7��%���z�#��%P4��'Vj��tn�*�k�vBO��BO���%j�_x *�3�\'{܄���O�B��jY���{^��@��$�FHI�(P݂{�f���wi{����Q��0���d��!�}9���c�I9Ξ�R���g�?~�T�v!<����P��^ܐ��je`� d#2M����?�(8���J0�A��V�.���u#�zBO���($^3x�*$�$�ސ��r����=�	>��IA 1�ª�x<�}�I��d��	�]��KH��י�-�*�@~�L�u����ߔ���;�T֙��]p�@��G	ʅ`�,Eɏ�s�u��$�J�}$�T+~�<�#��!'�s�D��2O��ȊJ6ы�����}C���􄟳�!'�k�`��>#�zLm�I���ꄜ���P�?U
�t6	�P�4Y>w���{����ܓ�a�����.p�� _z��n�$�ސ�wE=��x�^b#�4�	9�4��
�o8R�섟-!�o�|�%��v(��㞶�[�*�4640M����$��R�f�hB4S=%��U~�xI��!1{ �  "'�xa=���oi%���O��| � $��'>~��M��z��#�KX��ڑ��	>���}0�6�Sw��BO���"q��T�J2�'¨-ɦ{���y����K��D���& "q����t2O�!�c2�e��Ow����{��I?|�$�oT$��t��� �D���h2��	��%�e�CX���sS~�n�������Β}�2sd��"g}�p��h���DK� �n�<*�F�ℽy��$�2M�I�5��RIC��^��	=��s��k}�R�0�2��*��i&�	�m
>v���!'�t��UW�  w|�	k���7��iH|6�۲|*��$�� ���݆%�翟=��@   ?'��������;���g9�����G�7��Јy���F�X�ʆ��0�G�3�٣:*���84	�pv�Ӄ�r�2��%�r�U$�J�L1($ڵ�[��5�t���9^]�;w�w��z��:�ꪠ��lXkl�l                         r��f�V�RK�	�꥘�!�-[5��4H�6!�e	�݌Ii+�7gk�dcW��;�e*5�v��[j�\.��0;6�6�4p�.,Ͱ)l<W3Xr-����5�֜C2ۙ�l�Ŏ��'��td�a��r@0�!.��i�H��%��@l�뭹�x[�v3�-�Z8�
�/gF��{-�
��������mj�aو3�Z��U,�QL8trR1��s�&@�eqfL-���P[��g|�9�j�`֠�l�(�򪱬�8Q;�\+����7��ob7(ݜ�W����!m�cP,�(�8������ha3E&V����*ט�fk���Kj���`�z݌�ԛ���Ts�6�M�uY�'C���㣞Lו��f���3Ɲh�䆈AN����=6���Ν���@�օ�Th⭣GH���e�]Z���a�LD�c�)��d�T3���a%���i�,�ٵ�^�p ���i3Wn�I�6�ho5��@b�_b��۾{(��j��Kiƀ����m���ebP�ɱ8�"f��k/[�t&���US�;(M��Qv���Ħ�iV��p2˔r�0�km;X��3��X.��&�6qa4�mGK�i�I62��gB^� �����������x��=�0��P�@6|��&t�@K��0/�*�g�rw�y�;������    \�m�T�/km�5�3��s�x�/=s���� �*0���aBm�Tu�+:�_e+A��
�e�W���ev�䧎1vG�;V��U������CZ�`<�(l�������ۘ�Nڶ1�7Z[��'cv�cYmJ\�NN������T�0���s���qa�����cA�V���X5�&�uw��������f{랪�Y+t�I�o�J%i�ux�#��	>ѲjG���	�B�3M6⇄�����̐���!'�}0�� ��{^��B8 �Γ�=��BN����	<��$�$��2bi)�N��]Yj{ݗ�N��z���T�,R&)��fq�:]��s�������S�V\�bΠ}}�D��@��_�?�I���!'�|��hL���O�C�V��t =�� -�;!'�Xd��u|F����%F8=�h�^1����/��u���Ԏ�q��}U������o ���J2���*����^�;��~W\Z�؎�D�48�Ca�Η�+��㺱�ap&�e�W�1w�^�}C�~�]�y�ȘB�ۏ�y�1g�����ͣ�H7�-(
��5��k�{�P���``J P�
k����x���ihaI!eg3�� y���<�zsx5������J�A��1�
�]�#sY=�魻^�!a#M����D�ȂE5����ۊ�+h@�P��
�#.�j"gG���1�.�
���_��G��16�����UQ��5����(��G=B#|}�#��M `�Y�bUP�.���&�mH{Ю{��}߸>)�c@� �}�38,�h��DE�T�)��>@�1̔k�����8�0����]}B�f��+?����ݞ*���R���L�W�v��G��	 �;n�����4�
��+��%�����O^r�4��A��#K�oS��E�y���A�r��!Fd#72	�cǾ��V@��i�m����z=��_��p����<�,��9
)8��b�^N�������LC"S��B��!�rK���{��g��]�UUUUT  YF�u�l��ij&t<pV�86Z��۱V����dL�0iݭ� ��anM��cr��;
՚���6�v�������\35��<TN�ag��;=��Y}6�)��p��e�<����v'tp��ш˝b�uk~�I:���$�l~?+���Ddϯ$�f;�pV�;A�E�93�q��;�`]��n��/�c�婨SmF�d�s<� y������_ψ��P��E�o�	3}8q^o*w|�X��)a!@T�$�= <�4aeUP���}y+�����p����f�!$�UY��g�+���1x�I#r��:��y;1�v��n��e�%��q���u7][7I�w:?{�$������F�g��**"I+:�w�_�1Q3�t*AH d�8y��cC뽟�]P�H�i3�>�4ԏ����!<�f~��z�Wj���=@�sz>��Z��{����pv~��hyc1��m�W�z@q��'���	��K�$���5��luah@��N��u1G��΋Mtt6�������N�'�v�=~�x�s#L�`Jb�?���(i�ϥ��#��p���!ew�ߞ�!��ꡄwG�!����;�On��{�nC�kt��Y��\$�=!=�8pg���#n��'B��b�w�}�| �=!����s�_�$�z��67t�-�=hMۇ�����;X���$��q�P-��O���4��	?^}�^���3�^^
!hD�zI�~��$Э��,����?�PⳈj�d(�P����	˼�4O��7��Y� �!HAn����f�O�VI�LãOH"lOߞ�$�HO-�`�Pp���Z{�8}�bP�������0���k��E�*� �;cJu��07~;�}G�Bʾ�q}�	'��}�vG��BH�X-,�B�p��	/=�p�r�BI������C�����"�2T\��~q�zs�)�fy�	X����T��:H+��z�w�k 
���	9���Q����!��
@�f�=y0�o����d���|�.I$�I   Y$�v�g^�y� 6 $�m����{���[A�M`݂�6�x�Uƶ�*�T�l)"����c��OKƸ.�x�t��q�6��z�J��k�:`5��b�Mf�KC/��i��� nҌ�%v����(im�9$���f�*�L\0z��C��moغ�����s��ۮ�=�厏�X%HxF~�9ܐ�O�k� ���#�#����B��{��O�#}��B��ј������@U ��AX�z��_}����Y�}�8;�8��g��䐴��s��Owd����?P�?}��Z1$�3 ��EW~�C���=�8�᯹�Nvy���iP̠V��e"�Nk.���6���9h��f"IH�g�#s\<�=���C^g!F�c���?�C�*B��ili��4-�&��VhZ�6we�e��<�c�2��ZB�X[k�Zj�E��[;1�����0O�\��rJ�A�ۡDB�_zI禥�l����8|w��8��`r�m�xA�������؀y���{Xؐ��:O��	 n뀝~�4�~����w��G]y��PCD�.&�5Аڥ%؍�1a�ʡ\\�"䑂$P��y��[�!� �*��p��~���P���s��C��:P���zAT 8�,[u����O��������T   �}��@~~?{����9�n��ޡ��I		 �;��J;��tND)h�FT�J*�Q)%PT�P�v�j۝���WZ�s�]e��nMQ����o��Vw�0��S &T�F :a�k����4���V�g�mf���~�9�3Ȗ�����?N�gݟ~��}%m�?��8!Q��@WK����$�'v)BbI�!\�)����W���-6-"Ҙb)G�'�u���q腈x�zf@P�B�]���j��JR�*{�l�4#�h�R����0!�o�{���{/h�8~d��2�d� /��p����G|�W�w<3�CX�B����k���xa$�=���TQ���$�����$� �g�뎓��䱨��6�ۃ\�7��|�︺N&Y�G�,�x�w����*��C�oE��!J6�<$���s�+���s�ٔ�x�y�8�bPK��z@I;�=Ϫ� n<0���@�x���'����795����amB*6�>�A>��>p�$&F:>�OLe����${�! ��!?���I2��X�pە��Z�Xf�Xi�g' �������ø&�����S﵁睚��C̝
$�tw=���;~��=ׄ{�vd�;e�<R6P�&�I>���c�	��zBO��a@�{�D�q�����UN�=w�b'�}!$Z���
Q����8s��'�v�C5<�.I>)�D@ҡ��|�;ـ    62K��.N,�9!�o��]	Є�ey	ٲ�ġ��\��#�W<��T�c�z�nUr ��ä����Z��Ԇ9�v�su�qۧ��6�Vm���;B�4&��%��e�D�j[��!��TS4障�ݰ��K�zI'��M�:�V1�v�r4��X�s����)��ɠg:I!�$N(	��'�퐓�u���
�y�V�x����Z���z@}y!$�a�j	D䑕ܰ�/EisvC�T����"O�z@M���(�2�eBcAw���d�{d�֔D��N�14���$�G��B�A��T���ߦH?��U��[ST��gn�Dq\8=��A�ѬB�,&̉�68���5 o0�g���+4��J2$q����d>�\=@>qe�#�QD�����P?��r�,?{�n�f��%_�8V^A�  ����{o�BI��cdl(|��B���$�|�'�A�T �=��	=�-�$)\��pv�5|����u�
��������%LH&+���r0�z�9�C�L��h��?
���"ܒ������~�P$�=!>���8�e2�>�$���/�}���ۆPIv��:Q"�I>�!��?U�*�����n�!�S,F�� �"��X�/�A��p���-����z=�3�7�ᄵ���𽕞9��F�.>�����z��'��	�c�$bH�V)B���f�&[�E��	y}��ϝ�q�v]O t�僳:{3�����b��$���_��=2&	�t�o����9������{��|A'-��*a$����'��ĸI w���ܕ;������ޓx�a'��x�!��".��B�?��/��H66[)B8M���9��B9�.οI�Z��3��Hf9�>V����g<���p�.%C�:���l��8;��<��	|�yxH3�[Qț���������y��W>5Hߎ�%*5$1N�����#���f����h%���8G>�T���T��}����}?wd
��s�!9�>��	>����B�T=�����'�/��g✅�
��*?(d�	�i��.�    e�x+��N �[�vG,�;%*�n:I:�X��[������\�X��=R&<�nm�6��7\�̶�ЙQ�rf�s��B��ژ�宄i�6�r����I������^Cut�Bq�!��ù����vj���s���=t��mm@]�&q��ݽ�PC�8v8�����_��Q��	F%+���Xa����!;]���������
 �vC���=�<��Q�(���
P���e�{6x��>���Z:FBg:H� ;z��m�� �PG��Cc	�u�d�7�I��p�α�����8>�b�7��tٵH�T505�$�X� �6�jZdƺ��rW������e����Y�Bj�@ �uA�F5�?~����f5}�n"����^��0^%cw22
 ��=�7�)�`�d�
b"u۴A�P*>����  �xܴ${;�˫�l�dA���.��	PPd{�p ������A�dD�+������2�Gu7U\��ʼ��/P�A�|pdD��`� T����p �q���E��s`�" � ��{<���&*���"���c��QDA�CՀ��
b Ƞ�y�md�%A^�
�A�Pv�+\��.�]�b�*��^��&L�7��q�p=`��ƦK:��\z��LT�'\�����dP|ߘn"���s��\� �5<�
�A�y�NU���"��n���ۘ���^AEPA�>xyvyZ��"��y�� �;�7,d�Pw�PsMAV� �bs7b�x�2�2"��y���"��K~)�ql<P�%THP~E��k�A�~k۰A�du����[u����"� Ⱦ
ET�n�U��� ��<��pdw˰A�;� ��,���;sR�w+����̘t�k] �_���I"ڒ����1,��f8%v6)���u��C�aws�����;��!�� աec$��{��K1a�1�l=*��~���M�f�j��4
����X�?��}A�P���_��c��~�"�X�@E�O)GwB� ��E���N���
"�pwٰ��:oB���c�����@XpDbZWj�v!,�(�j�����c��6�]���~��tyz��7��c��>ؤ ��2>���
#{�^<#��UP6qo!aƓj5^���YUP#ﱎ�W4�c�	�O�ٯM��tݡ�G��<A�VV0B�J���yj��pm�xF������I   ��������׽�{�3�������2��rณ��M��-�O�z�Z7��Iֵ���3B��L[=�/��Ϩx-���Y��ȯ0���v����->~}����L�~�鳽8�-�����dZ�zVKYv�%�����㛸ע'�{!��uCǙ�����ߎ���t��,)Q)�I�������4yz���/�o��mt��Hk,!h������B��6%�nXH�8JJwY�_<�^�7չ�p�崥��6                         	&�6��:Lo&�ibh��ve�-Y%��@��hXBI�q�׎r��J���m�����\�-6�bF6@8�j	^�mUS�m���6�A��+rB�����P��dd;`2��[q8�J����⺣]��d��V�f�/TԨ��7�����[�\q�^������[s��1oXa�ƽ5��ɶ.�Bmv:E�h��4腪��<C.�5UJ�ӥ)��]�i�+�����
��ȸ˙ti	6��Ӛ</���#T� �1l$�M�VH�oI����ڻm�R�s�'MjM̙��Mڌ��V��Xjbyu�@\Ʀg�Pf
ܷ]��:wn�Z��y��^Ty�k�X�[v���ڤnA��0R��[X��۞�j�.ǲ�dsen�WO�S�ܷ�cF���+s�6�)�.]iy�8�	k��y5�ʜ��f8z���U��b�Ŭ��Y+b��N4�UF�X"VV��Ki�k�. l��p�h�cRqe�p��m�#RgFϥ2*�+�-�.�lUq��ݐ^�n�� 8wf��6vr�r�;ZNCYۣd1�\/(�B�K��.sZ�qŔؠ5\qb;
�l��( 4��#Sc�ЭKq��N-pu+w)r�5-��,�X3���?�T��!Ad�"J���P�G���F�+�%[���'�~��_��J؇�W�@�����oH� f�Dx��lZ)[��M��'�MCàH }��_�    d<�n� �Vy����K��qHoH���4ֶn��1�6��oc��; ���u:#�Dn�Y�n)�+�$A�Un�焈��qp���zJ�ͺ��;sh���e���:q�s��B� lC $�m-��s�J�DZ���g�����D�%q١l-S���:z��tP6
�i����9�s���(W�i߾bQ�H7���Qp�����woZ�P{��N�,I���]�c��D��Β��p�$h�8F�6V*�܃����û��e��g5W�w`��ׯ�A�W%Ug[i��ka.�K���۾��Ls���V��'Z��7߼�o��_���A�~D��( /�}���
 �V7���A��T �DU(4Sc�r�u|띷�5h6]�B���8{j���z���u�5`�9��9x�;݈��bQ�=-Xf0TU��9�vF��:o�����F[i9aƸz:R�j5�h�s�51�ʥ&�J�`�;�ߞ}��t{a~��#���Q�9	*'�t�{_�P6sUpg�s�u���E�#.>U��dg[�U#�];��^�1�����'#;�9�u�o��y��^�2& a>�; �\��iu9�$LF��5CAm�2n6X[+�� �c]p��ƶ����ۭ��;����XQ�\��~�cs=*zރ�=XP'��;�c������#���J4����>���k�=R�ׁ�iE�ҟ@"�����{���d��1��k�Vjn���D`\�m�@ZMB�	1�t9��dq�qI������q�r)QH�����Y޺��;U@���3Rbr:����U1��(T�{ޕ��4��<x`��2p<̓N溻멚�۸Hj0Br�u:�m�[ �Uߥw7��I-FXK���\�<�|�<�<�X|S��(�0K�
@�P�8��wv    T��y�/ue���˞Sv���jٖX�&0���x�D��=��v�*��
9���wR&�1�AEE
E��7��=p#v;(���uR/I� 9�-v�*4Z�̙ͣ�\�n֜l�7$f�8�F��icev������ڻq���+p�.�G��h�sŒ�LEu�7*;�bϾ�Uo�:���:�!����ݸ.�G��_ �	Gᬧ�F0�����N����޺�v�h�M4�z��-���o]p���D���a�ٗbJ��{ݕ�,�� JኤDK;$���iLa�����7	2�h@�|��F���c����^0�C.2�%9^�?�B��)�yt���v�3��?
B����,��K��k�o��3����p�Rc�eB�u�� {�b�g}�.���#�Y��f8�����;�ѱz���^�@Q��A�qfC;&5�]q���l�JE�£��4qs�X�}�v+xǊ+�c�:�
�Z����9�/6P�Ds7 ���=�~�hY#���d�vs����./�0.��"�S�y��09���1	�fgҳq��u�}�2}x��'+���6���X�9�I'����@�r��;W#k�;=��4cEB��IF6�\��ɻ�.��z���Ěc*ʌ�r�����u���4�dt�8���gf�����l	z�:J�E��f5wof��Y�l�T0�DTP��:��Z����a�C��|(s6��{�N��I�G�\�#7��#o5�����f�]�Hб�*�U��Y>���e��܂��ݴ=1�#�7t="�]]������5Q�X!9F�`��C����X���A�Q����1d�s���U����$��V1��P09�l�����s-��C�99��)'��9���ѕUUUT  �[�RM�ʮ����1�B��U�R�a���i)��v��H�%,��4ݺ��@;en�q�$��2�iPd4&��>yE8G�� �45�>Kn�oK
��� ��u�vK�\uq:&kk�pf��r��/�����II#ݽv��mI����NC�x����p��D��+M���w�n�}`M� �/Q� ьƣ;�X���K��0�E*)q�fk#;�s6U�X��F^2�(�r���;�}#��]�n c�#-k�3]v����I�]}�⪓Y�p7]r:w.�<ul�mf��N��P8�a�������0.��*�W~�;�F�K1�
���c� �ՀD�U���c��o�x�m7a�
���o���,���=��	g���JPp�3<��co��>����+'N3���������1���Ο>���ሖ�l01t`�ق4̴��i��������i��%$_�>����;ϟ�C�~�(���!�JE�op?� �:�{���x���4 h�#�<뷏�J�@r�����|    }��}	$��f�������$�~.���h��&����)zK�!@����d�V�@��f���i�A��C!�f�� ���q���ק���C���F��;)�u��C���C� P��۶���v�l�t�m�p�C ����Φ�X�i����Yc4�C�= �!uӤ���v]�m��o�_����Wn�m���^*�.��<Ǳ����=�!C��c��=���C�h��?i��� �� �C �΀���!���R}��z�0�P*�=���������w#`�\���-���w|${;�}u;�i��sN�`x͂���}�=:���SL��0f	4f�-���F���X9�,���\���������{�ߘÞM@�f@I�]K3үu���r��Α��l�䍵%s5�]�6���]w�N�E��h�x<7|������~�<h:������dG]ν�r�1Ĵ\bFg����M��̸xo^I$T$.��5��� ��k�ƣ��uv�κ']n�M�4����om�ߘ}�7CX\d�S�z3`���������ZDE��pr�`�~�y�ѿ{�p`'�M��u#�:��0�<Ǿ�����io�(���Ξ�}+��Aw�x��yႇ�A�w|N���    R���v��\������i��ݖ4���Ɨa�uv��ae2SvP�GT���й��#"$h�E(�/O9ӤX��f0�`F�8c���qBZ.Ûl����\s���p, �(q�K,�����v��S�wh�ꉅ��b�P[�����ݤ��y��̧"M�7���/�ߝ]�!��O�3��l}u��\$sm��)�kV�;�c�U M *��=���C��1O�w}+�5�{�^�Y��A����pt޶�_��g��1�<�9�w��M��a$`��j:mI[A��Q�Kb��7J�e�pL̀K˜7z�T*��c¥��]�2�Uᓞ�v�ˣդ�	��T�@�����ט�����/U��%AHAo�3]m��w��{=��y�����P �v�t=�pr���s,�؋��#q�e�:3r�xE��9�rI$��[b�1�u���~~����r���!�Cq�����������}��z��1�����a9�36U�woMKۃH ٶ�N2/l\���	B��^A����,#B,��+���\��3-�w.�	�f@�5���������g��~o���\�J�-��5оÑ;Z6����Jɦ�
"�1�e��lӅ���� 吐��f4����aTݸ/�v�-QJ-�a��ķR#�̟Ù����9�e%���{�n�V�%��}���
�@r�C�n�^�|�l���h����Y�c�M����gG�Z9�I�؅�\e ]%#LS�\�a���X��,I'��,�*��>υ�σ6|���-�J|oP��˂�{��C�+��l�G��݅d{-�O:��ެ-
&�D�y㸙�2�1gq�w���5\q2�u�z��V�͹�-�G�*��UA����q�    w[&�n�T�S��$�]q�O�)����vС\��^=����5��P���çm�=WB����:��)��ƌ�Җ[+Q�1���d��	b3nx�qh�˹��Q�'=�Ni��%rt։8�}կ���C2�yuǜ�
�Y8�&����msK6���ή�����Fs,Aw�n[�d�w��#1�U�ܕ}��H�ۃ�q9�5a��6Jq����-���Y����A��0Bp/�_�経;��������t�K1�R�ú�^fr�N�� ����.�E�S%+�K˒\��9a0sF6�lhb"7�F�a���LRA�}��22��w��U����'X���U��9��]��X	 ��� �
_t{�5��)�}ݙ�	|p&RN4��u���?�{ ��FE�C�!n3�yg���������P��k$���fBXm�7r#yl��N�W¨ U��IPG!	��F�÷$��Δ��	E��C��TA�d��
s�}���X����=�a��^0�i���ܯw6}�zV_�3~�]�u�"Y����W���ρ��i6	�Bр�P�Sv'~b�B�l�g�X$Z��2�1�;B����ş`�,��,�z���Ƃ��w]x~���}�#�]���s��I#N9ř�n-I�,��	4XҒ1�af5�.�)u���龠����; ݋CTN$fpa�_Qf�3��� �K� }h�����1��ې^[/��s��<�Î!'+4�wq���7�8�`���(�A��M5����2Z-��؂�g�U�ۂ��G��y$��.DA����6��Ò��g��D�1��t�0�щ�s�H�����7.H��˄ƫ�+�}�{��cx��;�5�EDL9�Y��[�ŞuVwo�g�R��ZM�
h>���s{��>�dE��D`A�o�M�U}ˌ��u����( o���d�H   �}��@~�?��{����9������8Hw<@a��3���H!(l�����jL+�:���f�lq�
,Hmu�a�sL�r��f�M0(�¦IfGi��P1�@04I���Oq&�"�F�`�'	��ŀ�+������g�B#�a%���.�S��- un!)i�Zq�^h@�e��$8��89e��o���b���˶�[j�`                         �IzEmJڪ4�hq�Ɍ�nL�{G"���FI�k���;���/!s�p&�Ί�Z6{�F�ƞ �F�QS��R��b�խ��U1��ɶ[�)Zɫfn]�m� ʥ�yN���z(v�b瓌[�Υ��'T�	�{u�#yLe��3����k��C��r��oN�c�Ŋ��ʼ9��<]�/A�õ�5;��\M��"H�������K;��S�A���c�ڶ1[�,[�d��A��<M��Iћc]�h���lm��%��a�:�v6�jl)����x���kJ5[rm��|�wc����J���󪮫�P`�ұ��h��8b����Cl�+tR�&p�p�ۭ�i9IL��R�Q�Wq���nr�)�`��@�����e�vl�.B{uq���[J�bђx�7l�͞"B3�y���:�.v\��� v���`�k��&�Dc�H0��J�:����r�T�[-�k5CAW���LT<��2�/[���:X�KU�l.�(��E�*��A��t�jZ�/Z�F��ciKf��`RkS�mMբV1 �`HV5�L�8��툳�`��䃔*х�UK����v��R�YB�n�5vK���b�I?4����@SB�}_��p2� )G}@�S��GV)0w/�Ӄr��0    H![F�i�as�k@ ��0�4lq�����Ô.*�*;uӳ6�*��gWJ�콶���cK{Bɸ�$躊NU9nxH��r`��sR�lMX�)Q�&��|Lh`Eӧ[ 9.��.���`l;�s�bj��-�U�ч���@o8�(ML�j롥Hj 9�́���o���͑��W�
~�]��/H
��N|�w.೶����U��-l��-�,�,b�����簰�߆:8K1�J�z��Y�p^�+{�4��j��p��G4��� ݕ��6׭
���$,$T��S�v���ۦ\ �B��
ڢ6l4�K��~�N�|�O�xP#ۙ)�^:m�aM1�����D&����+cn���	�o�M��2��{o�m�$��T�@�qV����o�t�R"�
��#���6���: W�^�ތ?bܳpwy�?S��Rڮ�k錓a���ݞ�!��`v�殠�#p2ܯn=6r�{�/�pg��_�:z�-�R}��;p^��6���&�@�V.K�=�9f����t�b �&q�b����8��!O��U[��#s��U���)i�4ӥM:��:n�����fc�]7{$l�#�BӀ�8�DUا��ܔZ6���,y��(��;��O�����,��n�#�b���a����;�뾶:��{���ȡaF����]��v� ���v�@�7-�[�}$ݧ���� J<N
D|��vW|<�&Fdh���qVe؂���b�v�䑈x�����۲ǲ���\N�]٠Y\A�0\B1�`����2펝WpY�Uޞ�	Q!E��n��>�c����z/J�4&����{s ����w��zF�I8$�8�ws;p^�
�}�b�G�~�ԐA#�H�=T3rW�X�>�� ����w�ϗ`    ��MeS1�=�;��È�C��\49�����i�a��ڭ�j	Ǳ�O���w�8T�yd�ZMK�j5�Ks�x�����vx���մ(,�m��a��*��j3:m&�\(��Eu�2[��S[m�e^s�~��I$�t���X�
��¦��Lc>m+�q��j[(F̑��ew�1Ý�,�k�C�y�airFMJ�ٸ,���sU�{��
���k��+�O�T̸/�����b��Q����f�ss`�Z�՞t!�����.(�n1�ylf-�W��>��x�$n#����0g��H��l�l]&؁4S���z����T����Ş���d$&�j>q�q<+h(i�`L9/��f��>g�.�vZJ1��\���E�gmn�m������;z�Zy���1c��[��lt�U~����=�H��j��k1���2ۇ#�ո�,���Il�a6p�*0��\U�5yۃ��+6�`D����Hh#�x ��W�vs�t����R�\��F^<��C�
 x��(O�B�b�X���=r�l����M��c�}�b�Z�9�d�u�U�#q�9oz4���  7���=�p�w＾���ٜ�;F\fЙ�.��n����dYH��^���s}И'_�yAyo���<꩖��rF9��pM�=�ZoF{��P?�c$m$[�����Z���{l�F�JQ"�7�7����x3������4��3�ryz�$��ቌ\�����^fJ���Z�9B���FG9t�θu�k*�^ɠ66��kCd�NN�n��.�Ѯ݃���:{�S{�s�^�d�	�Ss7��S�s���P"�H���7#����Z�����G��I�R�A�~� �l7`=^�c���	�bl�pH�Ỉ{C��xw�NZ�ܸ|�x�X�!RNb�ۻ��   o6�.��9A�cRc]j�jͣ��gr�V��T.=IZ����;W[�ղ��iW9r`uv�+El;zݤ���#���XM�&ex�u=PN���X��2Z[�xÛE|�݆�W�}�_>v�8b�M0t�3�1k9�ܓ��ns��rrt�s5�%X������y�8��ٸ<��
.,(C�Zs���0�P&}����ls<�C1�\�uW7rfd���Q�"��B̐�"U�{`���+���Oڵ��H���)��4�{���gP�;��.	 ���P�	"&�C�P$]���*H�-�@�D��w	pI׾����	"r%D�ͦ`�	��v$�H�߲�����05�+���M��ذC�;�N�I��jJ�yvj�z��!��\�A$L�[��A;�]� �'u�%�$U�d����.�uBH$����ZfI�1�)�(� ��5v$�H���%�$�`�hP ���l����P��T��$�H��p� �
�r��P�	"g�9eG0I�<��+���*b�Đ|\�	pI�;��P�	 \Ϙݎ`�	�9v$�H��B�@�)D���@�CRąEI3��2��H';۱$D�w0�G����-�ߕnΪ2����2��<睶Ԇ\�{uu���,�%�r�Lb�I�7�;i�$�o��A$O5�%�$uZ�A$L����qD���@����
HP�;��n	 ��7T'*��3��MA@�C4�ue�	��H�MwKK �	��U"�pP3��������    |�}��~�~~~~|�s����^�	�!*�V�M/X��aS�� ۤ"dm�[�>�-/^�z��:�s�B�$h��Pr#diL�&:9&�1K��u�h�kL�D���B$�qe.9M4Ji�4��B$j/E̍g�)hcBB��v�dOe���tglX��g-���9���'��dr�6�	0�UР8��Hqr��S��8�JE)�C��+q<�U�b�	����T$�����¬���W��A5�1ڡ$RD�5[��A<�.ӑ	����"�"���(���B���TMv�i�$�o���$D��L�$U[�E$M�o�������
q S��;y�����(ٙi�i�6f�b�r����9<�';wbb�I����	�����D�$��}��$A=�I��^
�v$���N�K�H'*�T$�H��n�0I�yv��H��J���R��j	 ���P�	"_9�L�<P�A9�nĐI������*#7�S������A�(,
��}�`�)���I�<�p��>d� ��!�1[�A$N���V1U��V2��H'<�ؒ'"T=~S�u��A;R��A$K���fb!Rr���W���f4,�])�x��R�.�n�[ W\�z�YM��N
�����B((q.�$�H����0I��.ĐI<��""9jr�H�H�h[Z�W��I}󶙂H����A$Ow�%��S�.)ʝ�I%�UYx��A$My��f	 ��.ԄD�]�\h(q.�((Bm��䑓��P�OX���6��H�o�%�$5Z�D�J����L�$q��LI�/���$D���L�$_D��\�A$My�X�	 �l�ؒ	&�|�<�ݯy��y���~/�`    t��{�<�ZA��dC�0j��4]v:�ph�s&uB��<��K ,3aS�n�$v�˚Hj4�v�ݫD�EeF^��,�s��n�Mk��L�Av{E�A5zb(�`+�{+Ԋc��ݻ1hZh�'�I��ܓuѕT�h����Mn�/3�!5qrv�g��[-�ˡa�������97U�P�	"_9�L���y�]��HF��΄5@�oB:҅�[HP�I>w����Q�T�;v��QI�a.	 ���P�y���k��l��M>P�	76A@��M��&��TaQI^_{��B����e�*���� #C3�%�'hNb�T��PI^y�L�5!�Csd		z��L�����$�n��BH$�{��3�N�s�' r}�ۑ' NO<<UIZ���`�[N+4�&�lW�t5��Q��5m��93���0I��v$�H��p(��H�ԭ!@�@��!��1�WyMA$�v�~���B 0"9J�\)�D�}�K�H&��J�$DϽݦ`�	�9,Ę+wX��b�I�;��.	 ���P�	"_{�L�$��ؒ	"o]+�+��Rʬe&�I>D9��y�*	"w�w��H&�r�I�<���Mʄ���2���Ek8Eh\Nn�,w��'y�%Ĩ��Vꇪ�C���͒$�E��E�#(۞��;`������2�n?��@�
���}�dP$P��HA$N�K�ȵ�V��A$��^J"�"���a@�n[pPDP�<�p���@*	ʮ�	 �&���L�$��.����LD�!�{UUdN��((bX�FdP&��q3 ��8
U*(_��Ƅ�RZ�!��<���v& �&9���	���$%�Kĺ.ꄐz�;�M�}��A;�݉ �'�鄸�����T		���-��Q1ȧ(�A;�݉ �'u;����J�M��0$�H��7i�$�x
O$��n� l9���,�`h�e�]F�;�d�mq��5/+v$�H�s�v`�%ĭV�P�	"k���0LU	���I�w���N��X����A&똥�5�3���0q��rv�I�<�p��"Th	�V#���x�F�Bߵ�%�*	���I�Z��{��$�McȅEhm�oBQ��i�H�O��{�lI�<ߘK�H$�k$�{$�]>��D�3��$��^*`�K11�O"TD�N�.	"�5�P�	"_{�L�$��v��H���ߕ�,fjk� ���s�0�4ͤR���enn��j	 �u�P�)"o<ݦbTJ�w|ĺA$N�K�ؕ�Nc��h�rk9|I)�ߏ�'D�	����I�;���$f��A$7�ky���S�:EE͒�C�*'w�%�=!QI��(9��'�}y:' NC���eU��y��8y��%�$f��RA$O�k��5@*����fĐI���I]��U]Ue5�I��(I�<�]妠�	�;v$�H���r%E>E:C�₸��LJ��.�    ݴ�;B�&��;1��%铷u�S�2¹�z�s�v:wV�2��vٶ�B�3���t�9$����8h������y��M��G��U����Mܬ����%����CM�y�u�l��۬����OS�������y�/��,s�qn��c�NɸێH9S���8˻��]J�9��'�ߖ��bT_���;�A$���Y�I��(I�{�7�����24�(t��� �H�M�.`�kx��$De5�1*	�N��*L�11�A$L�K�H$α�$�H��wi�$�w|.��P�&��U,��%ܻ�j	 ��1$�ȕ���f	5Bv�v$�s��܉9rwO7��l5m���I��-3�*	�v�I�3���1I�VꄐI nM����R�y��,��&�F�^]����۳c��h;5듲rH'y]����;�a.	 ���P��5�A�Co��8EE��2\J0[��$D�@>`ñ ⧀��pLO1BH$��;�j�0I��v'�P�'}䢧��IR�)�$�rw��H��o�MA$�v�I
��uЄ"���;����m�A$Mw|��A9�]��TD����$���_p%A$O9�vV<%^%�W�e5�N�bH$���\A75�A$L罖��H��s��t���V��c��:6˸�˷'[N�Z����bԐI�9�`�)ɼP�	��p hP�Xh
�#wQ�$቎ �t�`�&s�Zf	 ��.ĐHhn���	��C�x�DȌ8BI��D�;�L�$��ؒ>��\�QbP���KT"��S)�/"o�a.&bTU�y�b����7]���J���)�$�o��LĨ$���	pI�VꔑA�Z��0I�v���]U���WbH$��{��$��1�w�U) �&���3��"��䂁"�4.��$lBc�낻���!�����Y�P�H*YM���Gu��9��oڤ���7��Zf	 ��.X���M�t!	��}H[J4ci	"r%D�ﶙ�T�'7˱$Dn��H�λ���M�
�aOQQ6�aG�"�"�f�((+ovP�A5Tl�E$L�]-3*!PK�P�q��e�(T	��uЄP"	��U	!�D޻�L����vi]��%LeN��=�vđ<�Q9�{�Ԣ�c���SPI�W*��I9�-3�N����PI��%�$9<<�*�۵��ʹe�^S3��K`ݰi�UU��+��0I"B�"�"���(p��|�A$N���Rf&bTC�x��P��H���qw1%YWw��RA<�n���D��0��MUn�;����}�|��(((��@�L��5��n	 ���P�)"g=�`�	���I��w��Iܗ
*]Ue5�M�G*��I9�*�0I��v��PI����#�n���]Lb�I�5����A9�]� �T��p��L��I�,�5�z �m�  ����ۻ��s��IhDIem���R�z�"T�d�X-�	<�����"Ƚ7�g����ή(q0�0#	�q`��1Mk1m��޶���g�~1��>���w2M����h�&�!XW���ݐM�X'ٟ��s�'�v�{o<y����-n�A�N�U��$2�$�v��ٔ�s�"�`�A[c�ͥ�-�m��h�2S)��@Ƴ|�����
�BK���5���Ml9y	/1`@��( y,���LUM�6���                          �u��c���Ц ��������A���v�^[
O9�ua\��V.�6^��+hJ�ٺ�U ��� F�ڮJ%���㍍l���::�j�n:��$�5��e��v x�:�;�2Ԇ鍶u�s������A�0��c\�v��%=,�w������(�j-t��6V�1���2O͸kZ��N��	`7 $r���I���cn (�6�*v�Y�^��e�]sm!�����`�怎�]����9طm�����Rc��݂`r�".3j+�m�і��0�tYV�d��|}�*�V�f�*��*��k�iqn��F��h9ca��0��$��rc:5ɞ���L	�!q�Q3!�	��n�Z�a`�#�mʖ�� �鮶({]�u81���tqLu�S�gx���6}�"6MѠ����[=b��H�.(������c��mN�IoS�qW��zR��snސ�zY��J�p�gQ�6sdmZnɭe,0lp�1��gQ�T�n���
�hU�ѹ`�]�:pꗪA
��υ�OU��d��.CtZ.�(�� ]x
��1H= nͥ ���F�H���H�-�
���S�N؄�����K6�/a��!Z��݁�]��(N]N1VSl��X.��Jd B�<@��ʦͮ�W�=NXI`��2@��]��F�{�;���N��:��    U/,R'k[	d�@�ذ���n�͌f�8%{��|���gY�l ^8��L9��;3�s&������1(���]�n���V4Fඥ-�ֺ7d8A�s���S�FMN]�C�&Ɇr���s���GY^�ؤ���tu��Y]k34��s��(�t��W1X4c[� ��2�E����h"{�R�ݝg����e3���(~ΙY����((]ꅸ!Q��n
�'uل�$�gx�TA$K�{i� �Cqႇ�T	��G���	7O)�$�s�1 �&�TMo|��*PO9۱$����0��M��8Y*��Yx��$�H���i�$�s|�2�Y����z�L������V{�&c2J�99C�PI
� �H�Jw��\uBkxĂH$��ﶙ�C��߾�3
�ƍ�I�j��|�x
;:㜙|�n�P�	� Ehn��H���J�Ĩ<��Rs<զ`�P���A$N�
'1:J������	�c/̾ �P�f���� �w�*%gz�C0I��v$�H�w�K��4hh�H(�I2EEhg�%��BH'9vX�	"y��.	"v&�x�I�;����K*�x�SPI<���t�V$�H�y�%�$:l�@�J4;��8EE�F�1f&1bH$��{��$�gXĂH$��k��0I��v$�H�I�c�T�f,[sv�=L�Ǩ��4�˷�.9t��-�9sM�MA$u�w	 �&���f	 ��.��FA$O<���A9S^�QR%CEhg�e�A<�bB	"y�p��L�j�NU	"}S^��1�/urcb����@*	�˱$��);�a.��a�R�
1���	"n%D/��R#�P$P?��F
r8ؠH�H�ra=]��^�By�ө�i"8
Q%�Ӹ���]�poq��e��̒HݗGm���ᣵR�yd�z&��'�<��ɹ"1�H�{�ywn�Ö��	�f�8���#c�s_��Ϋ����6�
�Cu��p�Gv��p�����܎<d�7^v����g��r�I���:�E
{γ��`�(�j7�2�a���gZ��� n6�1Fde)@����Μ��Ɍ;aYb#�ad��:7vJ��!�Us{�H$bF�#!�+w¨Q��U�_���*��H�o)4�N�VGr�s}B��\�cĎ+	`Ƣ-���gq��.�'��C8��1���e�����w]��h
R���"H�$�u��    �Kn �f�W(�p��%�m�HP ��R�nm���^|t[[kQ]{����&���oGT�8�<�C�[=Br���6uf��ݢ���;��-ɢ�y�Ţ���VΌh�,� ��6�6��X��U��P��;�����~*���g;*�	���ݵ;e�����<~����*�wx��ǌ�܎7��cW���ל���fA�*���PQD�N*��=�u���y�S-X����nk��bj�}UB�߹+�jGRCa�e{u�yj������\�x{�I�k������4Ч��I]���P�&@�Q��6sVw��.�;�i 哈�D&_w'���  9�6>'�-W�zW�J0:����;��3��9�J�c��G-𓻢BO2����ŪIw$$����ܒ8��8��;�fd��N��I��;�M�sd�A臙��n�+�oe�9wi�[`Ҽ)R�k[�V��c�s�$$�d��-�=T( �]x���&7#<$�o�$�d���P�+�$�#6H�AmNwvBO2������)��0�>4��"T�b�  ���	9�2}m��0�2p��R�������}ܐ��Kۣ���F�A@Ƣm�n�x𓷲q#�ȁ�ޱ �9��Uv`͝u3c56������P��A��D�(Ͱ�����|�{����]D�<0����z!��o��n����n�p���o������P��=��j���tz��ވw=P:��z�&���T%$IC'�B�d��n�'��ܞ�� �D�e�R�$��:��m����ޕ~w�|�qB����<D��BNfL� �f����}ȁ��<=�U8]+-�1c�v�m��&ڑ]Àrq-�Ķ�)*�=��1����0���8�[qYx���	=܈���p�N�$'�q����"�5��M��Nc��Hx��%�{ ���eL	(��6xO����xI�섞z�Bv��񄜿FkB.8o��n�I�]���&��é{3y�H����'}y����<���v��     Ji%�͢[���`��x���_o��y:���2�RGn��Vu��e�t�sl�x��m]u�ƺh͒雫�y[;��M��95�}Vѡ'��]zWҩ[&��t\��d�,sy�m�.�M3����5���]ܞrs�������[��f�\���E�AV%1bf�lƫ!�S����L���~���	7oL$��'򸏑ݐ�������p��Nc�';�w2_=ܑ�����Pv�۠>��@��V���!%[�\$�#W���%�	�/{܇�-�!�w�o�&$w(�oDe"�	;y4�j�BN]�Ď�HIC��|��*٦��3()��pjK���"9S�]�"D�禦��ݴ�/���P>�`;�� gu1bb��Ie���B�R�� �*���X���!'����ߔ���C2~sV!cY�^�����~1���o@e�H�b��2D�	9�H�����	9w!>^��$�7�$�����%]�o�!'s$Ďn�':r<�H�4B\F35��ǚ[h��Kf0�]Y�l�˨;.:�6MH�서�A� Uqv�R���5���)�}������'1��O���#�h������.%��I��{]=��o��� m��  I$�I���n���rI&((jT((tSS)����XW���fȚl�f��q����,�#�@�L����!") �H�4^,�հw��f���n<ř	��'�)b�Sh!24)�d�!�t�s����$9�b̕
a��-�0�������PdCF�u�"�m���Ym��n$�&������dd�ſ=�߆ohf��r>����<�fy����	���Y�] �h�D:��@T� pK��҉�"���p]�0ف�m@>����\ �����Us�G�!'��ש��j&��:( �7y��'����BM��BNv�P�F"�M�wrI�ɜD���ۆyn��(�J$5Y+�b݌%��.m%��XM�MV�]��Kͮ����{�BOm�������nHOx��[�I��-��!'�xbH�\�����|�h�h&1$�?JW�\��^HI��H=V��rJQ�	9{w�����ԝ��.O�� V���` ��S��
H�"���a@ANp��ټ�������Om鄛�$�M���	t����֎pݓL�ZRZĖ���f�зWiF�U����P;�y��|P��ڄ�Ƃ���"��o\��P�G��a'/d:�W�O����0"˓lt�(�����@�����{o,$��}T���$�n(I�I�NIč���$�P(_	���P�Ֆ��Z�BOw$8��ǰ H� T=���˰    �g:z9%\�suI.������Z؛�D�|=���g:C�]�b�t�%�[�e�N�\\�6X�gٌ6���M�w��29�۳m���]5�]n��+
='b�h,�wRo:�gzS������Uv�R��&�S���>T+*������$�&�(9M8˄`L�������Խji�U�&\\��s#G-�������	=�'��&׵BN,C�끦�Q�	+��p�V�BM��1";�A�*�m#�
e0BNp��􄛷�bG���$�\��X�)`8�q��	�P�ݞ0���L%._�R^�	9�X���j��&�ᄛ���{�$ݽ����t�M)�j[U��$.EP�J�24h`�P�"\2�g�ޯV�����ys$��0�N&�o��ݓ�*"��ઠ;$޵򄟱��v���r�M�ڒp�w�BO-ᄵ����G�r#��Đ�"d�����&�$��Ry{*jG�P��P�ֺ����}�z���T}�X�כ��'9<ǟ�Vfv�e����P�R��`�5ķdp�!B@BNt���fo	���C	0l����)Y�C�'8A9����[�	<����rNP�IZHh��F5
x3$�1�rM�r�eLOX!ț^/�D���W
'��]�;�Y�Ԓ�Vi�eq���P;���>b^o�'�������&�d$�*�7�����D���] ~<�|��jT0�s�8�=�'�9y{p[��[�W�V[��۠=�� u��{���(��4;��{ڍC��y�D}ވϽS[�1����p��L8��'wd$�2g7{$��I:E��b��!�8I��	�w��yܼK�6�$:���x�*w��ː࿠a ςh�8I�~0�_� /y����@���w�������	x�hi-l�ll���и�����XјuKq���/�{��Ow$$���p�EYҙТ.�<$�섞�HI�zo����O
���a��(X����&���'3D�#���i{vs����.	$�5�;@
�d���GْOG�BOQ��Y�+������ {��(���<@���%����$�ܪ����� ^l���v4��ͱ�A�U �z!��k�q).��n���W:m��W:��˻l�<���wFi��v�d����]G9Z�%S)���ib��xn-i��p��e헷J���.ŀ�>�G0M���l`��Wx��u.�}z	�";Q�9��_�J�r��a�gB���6w��g	��@jNs���͍nl�+r;�m��({��DBI��� ��F!�!�ۜ$燤$��$�_�$�d���7��X�a"�$����x�&�d1.��1#��"���Sc��Z�P��.BOw$$��ݓۏi�c��>�}���@�͂O� |(R���$-"J2��gncv��-R�J���� b¥�l�]c�]��ߔ��!'���&�d$ݑ��	6�Q>I9����:; '���"�@��} (�~��Q"��>��88RY�!&�$$�=�d)��������	9�!�ro7rI�hjƤ���`��R���%m��	7ۂK� ����CÀ���&�d$��$��a�'wd$�.��d�%�
��ޜ�\�p�c`@Cg�l��+5X]YM����C�߹���@��T���U�.Ӡ;�`��W�{�!���sԑ=�53�:%�EY�';�ܓ\����6+�S�(�DZ��_���'��˄ݟ��m�#|�F�d'��x!'��BOo$$ݑ��	6�B'�$o6#'�p�I卐���	?��;�9�"F>�!�l�7q8������-W��]�+�~7�}$��BO}�{{Ԋǈ5�B�*8�΢q�B�6�BOo`��˚G	'H�-��B
�.�{��H���	,�!%v��$�ٌ��X�&�I�v˒g|�]I���K��R�:⨯ �o����9ﰺ'�U⮫$��A	=���.�HI��'R�Sj�%{0��ּ!H;Gܖ z�׬m�x.�a�$�&8I��!<]��$�l�<��$����Q�ď�굲~� $o6I�zI�Ič��RE��Q�lf�	<��KH��	<��8I��"JBb���B�W�����r{쐓���!8cd�⃄����$��jw�YrL�V\����IH}�I	 ��G�PTA?����HW�P(Af����{��]9�0S1DpATF�)DT`��"����T"��A�cm�k�k6�>䱼�`[mm�Շm�f��Y�6;���͞�!6����񡳛L�f�Ն���0��o�����[��J��Y�4���ܶ۰�-���T*Ȃ����-�P@�+�������0?��]��c��g���3���*
}��@�Ǥ  K���AL�� A�)�H��AM�c���� e�� �����������ߎ�z��  �f�~�� 4~'Js�1�����{�������(���!��QP�i@ݏ�?{����Y�K?��Z�A�8�
}���~��}���S�r` @?�DP�����(?�D�R�%(~C���� �X��_��J����jۜ�m�**�����*Fj?��I"�k�}����(f��͛�Օ��e����)�L�+l�,i6Dն���F"�1m�X��mmkf�cY�͢a2be��,��-�-X�%��Ve4ɴh�e����[4�"�CM5��PQ���h�Y�����""l���m�e��a��5�kb͘k5�0ՙ���,40�m� @��{
��W!�w�����?i��J
�'�	��QT��g��q��_������>������w�/���,?��>��DP�֟�KC������S��͓��{J���������-?�ԟW�{��O����A?DUHȟ�_��_�I��������w�c�M,��UO�?1@S�O�� a���,O�*������>�p�A�����Q@R��FpĒ��?q�`*�)Ia��H݅V�訪J��QO��(�WC�n���q�A�*�4�(
]��h_�?@S�~���?��>� ��w������8}}���}�S������~���������)�蟬C����"���Z������?�o����?�O��#�4�Y
G�ΊHG����7>��C��Ǥ�k��k&��h"�����Y��h|��+�d�N����#��
~�}��S����?��|��EO�`~��}��!��*�t�(
~��X��(3~MR}��,?��� ���W��w����)�k�H