BZh91AY&SY?��{�_�pp��b� ����a`? @�           )�      � �` �x  P�	�P P� ( ��R�JH�
P�
�R��(T 
� P�PU   ���   j�Q%H
 QJ� ���Ӫ���,��y�*{�B�yJť,��뗾���ۥ>� �>�ťv�7� ��۩P=������ {����8��� �
{��3�U����-(ZU ��*@ ��B�@�PJ&�Pt�Zsە��|]�NYJŕ=�� �|�W��ݵ�K�͕/p��Os��q���u�nR�eO>� =�K�Y���&�b�^�O�O[�]�sjt�ʾ���m�  �| �B��"�f )��Ŏ��Ӵܛ�o{��_}� ��nn�NN.���.sZ����N]��/�ϯ�o�x�W�ח�V�� n��']+��V�_[�痢� �yn-ҫ��^��oܽw�zj���R��%AB��b� ����[�==�����oj�sn�@��_nL�NN��<�]��/m�� {�J�|s=�:�/]���]�w�Ϟ�P���6��mx�Nێ��O�[o� ������Z��w��Y�+� >

$ 
(�� ���mۓ>޻��s��T�xU���S��Ů�9���}�O����������W�z�  nw������ {ڲ��Z�&���[����u���)@7��o�����n���,^�7�      i�	M�*�H �� b*ꙥ=�R�@  �� �=U*F�Ph�   ��R�4�SR      ��S�UJU#  � �$�T�h�4��=5���=C�3�'�����������7�a������}��"�����TU] ���@U_�QUq ?�*����EU]_����������EU[�%�r�0kI?�Q�M_����?ͽ}��P��Ő�`A�"�`6Γq�8�����O)��d%�A�[N^�k��E�a�F���r��ģTF�p��c�VÑ����)��),e��g��ރmY�Θ2���z��p��:�,�C#�Ƙ�nb2q�v�����g���7�VZR(_�QQ�x<��#�ѳw�����5B��¨��<�єM��U M׋����Ծu`I�2�6��!������ټM;Ѫ����3�}9f�~m��� Ժ�k|�?o0�xn#||7V;i�rՔZ�#��s�!�����y�ݵ�ë�����<��G<?�C,�l���!W�����%z+�J��G�콟�~�#�Ua��󇆆�! ��~1��硰ҧ�J�7��s79�xfN�f�	��D␘9	G�f.N/��6ay�d�1� �Y�v��fh���3��2����e��Fd�2�(�L�}�a�����Y��o.���%	�CzkA���d�y�kY�,փY�ve�X��:�
r=�j}]à��ki�E���kY���s�_�4{���k5'��r�Se�99�<v�8m=ۋ����`i5��BQ�d��\sY�����o���#�����g�k^h�{��x�'�J�z���^l�\�-��0�,���j4l�S��5�D��ݼL��<�M{F�G��K�`�%	BP�d'�6�r���y�v~�q�8{8u���7?�z���5�B�����MN�!)��}�O��.y.ER3$���s��\p��J4�0��y���X�X��p��e9�5�	3|Nn2,"�	�X'z�9��d�EF&&��Ų�*$�;6ݥ�5����ta�JxD���5K�P�3��5>0e�z��)xYg���4j�G�l<*����/L����M��������!?f*�ؐddAd�m�%�J����26�O3I��d.�d?d�����Ѱ��֍��牎�N$V��! �PNLc�� �<�!(J�L��(J��	��	���2!5	K�?n��{�}|g�~�O���hĜ�NH`ǎj� ��������=��c��clJ��J�(OqMH��r��Đ�(MfA%	Bj��� 4d��~�M�y������r��td9G�Ml�I�17!y!�@T	�F�WFC�Tѭ^n�}�N�F�fo��3�@zrY(NC��:�� ��h��%?���@sPz�K�m�rLz�����A��SBVߤ��20�ȇF��Oǲ���/'
#$��7�=���og�4;##i���R�}�3�2oT&� Ƭ�4r��5f8�u�1�FC:���%���37%1��ƣ�1��"�TU��kf��NTp��ԓ������������ �N��[w&7��S�������f�F�N�`�hv����X���P����V!�x׹�
,����g��e�MW�1٨J����MP'�^BjhJ��d4
���2#,b��1Ѿc�-�L~�0�z �i'��>�BrG��7!�Дz1���
� 2�r\�?k�(J]�>��4ddq��x�T���*�F�#���Q�É���[7o~p�(�����sn��Qȃ?@c�ٮW�q0��o����it�Luj'~[���xy��g���2LL��J��,X�Ax&C�HT�ZO�!(p5h�6��a�q<�	C��i�^8�o{m�o��K+=E��%AMG����%W����Q�9��9���y�!ܞ&`�I�������Iy��3n�sN�s6i�Z���s߶�������u�Z6oq�L� ȋ8x8���n繯��g�5^Dh�ڶ�۸��W��y�Q��s��\v�������p0\���%�ٙ�y��ǯ����:*�k5FBV��p��Z���I�0��J��,C!)O�m<���h��%�rԺu8�	X@nP�	BP�%	I��r0�-f,dcA����(M�P�%)BP���%MFɌ���78�)�ƣ!,vk��I�4�8i5�|�i���-$h�7��z� 8y�#a�#��V�:�f�K0J0k#52EV.YX�@l�%	By	C�ְ4<��7	C��J�����v	��#a�0�B ��Z3���g�?� &j"���M�3N.N.C���"�=ލc����	�L�<Fi�Թ�Jn�$�Y���9�Mu!�6c���0#���Z�>��K��<��cUO��B��^��$UiJЖ}bJT�jt�b�~M��4j��F�mڞ��kn�a��Y.9a�2�ׯu���o<s��c�}��w�s|9�9h�s��Q���!��>�,�$��y�3[��M�33Z Յ�5ZY1�Z
%�����J��(J��J�7syfk�k�����o�̼&�+�d%	q|r\k��NF�!����r5����ysķ2�K�6�8�`�h���?[C,�'!!���H�2\��(J�J�J�98/�������M����$9��j!=f&�r���A�5|kU������!>�M�A��	�L��F��V!�`����J���A�l�0J5�n�����k�{��_��zѷW��g �x�4C���%b	@G��(ۏ��ϭK��s�5���Q5&������f`HfA���"Ǟm7N\,��$�y�v~�`A���TTA�����Fd�Q��9; "���QP���(g(J�5��5-C�A��,ѷ~A�a�Zs+|2�eʒ�Z�fr�<�EF�l�Nh��Ho.���AF�7xo�MBP�' �Yd�x%%��sa�e�&���p�2��)8�9�%	BP�%	BP�%�5�%	BQ2V�?~��X���5�<�>�N� �O��>�ݨJLL���� �%Bo0J��(�	BP���	��(Je�B^	BPm,���֦�%,C!)�12�	�`�i ��@p����0Ѵ��pՋ�|ك&�c��3�2�t�ۅ(r�1�BxgA��t��:�	BX�������#Ȃ��	BP�d%�\��M�?f	B~�0�J��(���&���V@d%.��:�6���>ޡ���#�ӫD�����8�D&A��3A�sY��BQ��/��da��P��c?�`�2�Ѩ?k6�Nr��ٚ��������(�999lJp���X%	I�l
����2�TE[3%!j5��j��en5��k۟:��X�q�{���zw��z�^"'�jP�h��&J_���)58�7f�~�?��AD�<���23'��� �Re��2(�5�+V�[�Y�aZ����0�	N.K�BQ�I��%	��4d���x|��?F��k^5Y�l�%���}���Y$�p|5��^��Ȍ�H֭�8�r?&F�o'�����5	Y��W׆�g���x����Y8Y�XRR�ٗwS���rE��&)Z�Kߪ�*��Ŋ��-J�B��]��V}U�[�T��f��Þ~�~�����ɽC�d`q5!�dh�X�l�l�k��f��}�,X�pUe��5�\���&�Q�F�.|'ى�db�.`�%/�!+N���(J��!��%	G�d�d����L�?�L�Hş�۸�.����ŵ6�T~߼F�Kh���bT��۾oU~^��ݿ*\�~,��^�yo������&c��_o-���9�0���4��8���5��w����6�b՟o��n֌��#q���Y��Fx��Jp' ��]�p6�o�����M��n�7��1��058h���s���#4[�l6G��q�O��,�FӚ���i�k[q��8h-F�F�SEMa��Ǽ���:㉫Y�xm��4�A�n��(JR��(J��(J��(J��(J��(JR��(J��(J��y	BP�%	Bd%	BR�%	BP�%	H{��%?.���J��(J����p7���(J�7����	F���<���������4�5�n۝�vp�.��ǟn�w|��!+ 2q#,��E�o~~��kFFsF�����kPl<�\�E6fZ���%z�N����?BP�%����(p3#bBɕK���T����U�i���ڻ�:  $ ��          J     �p�   �� À)E�y��           �Ҁ���� �}�8		  �   �     J            �         |              �            �        $
P   kXs��l���(�U��mC�x�  YL���r�mIT(�����m�Ե��m��.�Ywk�I� �`      ��m��[��k$�����m��S�A��T�m�l  �ӕ�� -� �� ��M�@pI�Z[�� &B�Ӗ�   5Sl7o-sZ˦�i� ߛ>    �  �� p � gM�����l]؛�;m����"D���CS]�����@UU�:&�@Krcm��k�m���I�mH	nm�m���-��m   �-��m��x7m�f��UW@l�K�@Uu�%+5�-���U7%U@~�  Ԛ(�pz^�����]5�� m���m;����mUPuP���[Ļ,�*� �H�+� t�i[  8Z�T�*���K�� �`�$n��p٥��l�rKi�p��-j�21d���pq!Ӡ�p[J ���+��a�7  ۶kB�a��&�[m�� mI$���u�q����  �  ��9��-�8��9��h�[`@Hm��vm��"�0  í�����m@ 6�� ����8pڻa#m�v�8^�tP�`� �W���h m��[x[zBޠ ��[[v�*�Q�j���_g��I     �m6��l  $�$��%�l��ֶI� $p�6�k�Iwe� ܋@UU.�[WV�ԫUR �K8�]����UTk<��q�n�vE�e����Z$�`3��m���h u��-��{K(R���  7m�۶/Z�v�8������� ������6�bY"I��[ ��%�C�ڶ�]�� HH  )@ p I�m� j��m kn$�n�m�pm��� �l�%�ZlH-����-6t  m��T^�yz���U���m�hm -6  ��kI��o��oY7�t��� �m�I��!�m[xlu�[KhH 4P6�v����	 ��I��ض�    �   4m�h5�L��p  ���F��ŵ��I����   �� l         Ѷl�ڊ�Q��2t�UUM�T�Ev�m�k i6ڐ�`��m��WeJ
�T��(@U� �n $@6���Q�Jg���
%U6�.�Mt�" I?��^�[�� m��m� H� �I�mp  ;m�    	 m�2�wm����� k�l��  8$�ۨ]J�]u �ҵ�*Ƭ���,2@[A���z߀    @    ΐ�]�-�     �$	 �`�a� �m�a�� 2$�F������`� -7b��O��e�` �	t�I,�   �H          Am$[��Kht�S����9���KR���Z����ۀ �` ���[@ n��K:G mm�+���v�;T�p@iP���@�S�����j�������V�s�;`���2[��m�^PA�n�U�����6r�5���m��S����ke�C�����J�u�T���jRYv��PY�6�-�����j�%mV�$z�I�mm U�HVӵ��Y���`$� �ʭԆ�Uu`R�����n�nmm�t�`�6�'i�@�֤`◖�����t� ������m���am6Ͱ  �d��^�W���P;���YV��P��^��
�����@ ��l��8�� �nV�Rɶ��= -��  �m��v3l�W����\v�8�)%I��	0Z:ԋd�}��| � � �b�d0�[*��-e(���l6ۃj�f  ��@  6�@   	      lv�Cqi�ye��L�mKN�v�����9�����hq���@�jRZ���R�@�r.�a��e�4Rt ��^���v-� ���m��� I��p���[����U�v
[[Co`���N�i�*ඊQǲfJ�H [C�mf�Kd��C��[�M���6�S	e�f� �޴޶t�� $�I  )@ 		6�`  lh��H8� 6�n��5�wK���� �� ��워��UWUPR�  m�ɭ�"E�p��}�흕�eZ۠
��UP�m����YC��
���6�V��    k�%( $��[���m�H�)%�m�h5��u�Ͱ�)mW/;X¬�YZ�]�-h ��)#	Mm�mtq�$6�V����%Y4ѭn8	8۰�ۤ� n��m�R���m$��|m�̀               I�[@a�V�!�Ĝ �i	6�6�ufնݰy �m����I:l�`�   [G8mR�,8�mi������_^�N,�u6 p8rN �R���6�8D�΃~/�J�UUuԬ�*�
��    ���h�� �d�f8����l��`   �7l�lE�K���U��@)�\�-l�V� [v��)mR�� �6ׯ[��U�������+�Z�7`m[��� �F "Zjk )@  ջښM��^��l[Mk[[l-�   :���3�I� l   9���-�e��[��v�mSf�Z��[I ^��H ��Y�m���O������t���@�eU���]��ڽ�H	 oY-��ە�U���h����R�[@  � ��8�6�$��Jl 6�6�ֵ�r@�:�3J�� RK� [B�k�md������}�6��$-�����0���kX    l  ��k�m!��ժh�pkָ��I�p�`�I���`8  $   ��@��H�m�ڷ#t�ǲl� ������v�hеUUJ�  h6��P*�2t�4�6���	 ��1�      �շl����� h��K����tu�l���g9m� H ����ܲ�  ӆ�Y6Hl� J�e+���1��8 H�m������6�86��86�@��  8�@ �2^��a   ��hi0   �   p     SLm��l H�V�R�.�jgXT�h-�],ͤ�V�h�-�   H ���6�m��nݱ��  �[U�]m]@r�� ��YT��)Z��I�� Gj�XE:D�m�6�ݔ�I�l    ^�6   m��p�x    -Z�u�ѻc��+*��(p�T���$�d��at�� ��kh[Gicl � p	�  m�   �    �       ���7Z0Uʫ��
��CO:����m�BX�`� �   h -�Ym�����Ā�c9��U@�_�����s��p��z�@���U����[iW$\��� sm�m��� �mٳd[n� 8    $c�   �z�km�mI� ^��8  p�@ 6ہɷi�M�   �� �ȥ���$6�� �m�L.�s��$��D�  m �d��  rF�6���6��5P  �@�Ͷ $    ��  ���.���  mZۍ$  �&�96���rC��	 m8 :�(m�N�� $��n��m�-�o���M@�8�X�[x5�   ��~ݵ���[�� ����H pɗ\Wf��e퍺^_7-�9=�RL���������:��JV�*����@�6e��I�F� m��e�mb2-UAg��2�	� I ��m �����.��h�ڰHJ������ӛ��l ���QUW��EUW{��������ο��T�h/�PM���:S�	����B #���S��C@"����秠\���<G� �C@�
�6?'�
<�. ��>l�=�@����S���C���d��C�� ��@ا� �"��x"'?D����i(� H!H��f����%�B��I""�dX!�)V�d���P�AOU\�t������D�c�qE ������x���M|[0z�
/�U ���*��~L�D #���=Q<؀��UOA�H���E~B >��?�i�� #�|/ަ
��]�@@�T�x�� ���#� �/�����EU_��w��G����	(PY%@?��1)�I'����v������_���  � � �       6�    � ��U�6�n6Xi6��f�6N��D����� .�M�'jN����amZ��k��6�b쁘x�j!�Sf�5��=WNC�/K*k'��	���@=�R K����p\`�a�+vi�B�.�m{Ej�A��0�Q���kh.��S=N�6^w[E�/c!���y�e��F`����A�=tP��78h�vH�v3�����Q���:��%]�U��WV�U���۹m� ؆^ ��raŞ3�B���c�gY<M�/Z�Àʫ�i������(gJ*�T�9N[��eI�cvA���[u���S��b\�H�h&v��{m�#�eՙыY�B�@mm�e��u�i�f�����M�; t�-�����q�9u�!2�mM���#���uԵ��s�V���F;2�!7@5Ι��{m�$åS�;c�I�g�g��qЀPUd��q .$�]�(�N�s��gps$����;S����"b�ib��<�@UN�V�q�m<��.K�����e�q�+(x!����8�l��ʻ]�f\ ��y�l  �&ݸP��U(�%�͹�hc�� પ�كZ�U���ѭ��WFX�e�gpL���cTp�;+*��&�#%)�M'b�L�h��Y��#b��9�Z�]�v]cNŁĒ�Uڴ� �j���*@�ت�C��r&9�eiX%L�뙤�Ki\l��� m�%�Zn̛�]q��6
���X5 �9���bjU�����w.,)�ᕦ1*�Kh�l m�m�Z���N�E��^4�WM�c  `e�]���vR��26�n��m�Bk��v�k�8��VV���` �C����g��+	԰�,m���QW\���F�͔m`:�ݮ�Zԫ�觎	vS���ww������������*S�h�%�-�_�R����� 
�������yy}��y��c<.�j�8}sD�خV�%)��C;u��²�Y�^
9���֪|*]"���	ݔ�;�Cl�1ָ��̗HNgG&f�c���Qn�ۻ&�B�!L�z��:���Pp��J��89�tY\rN<�Az..�u�{;ɮ�ձ۵�6�LCЇ/:H��7u6�u��6�[��7k�n{��{���{�[�<�.{v����^^����l8<��evA7.����!�$�4�H�������ޙ ��O���p��HkĤ��	ɀ}�n,�!$�
$�f�^, �n��{V4��㙉��&�p�� 9�T�7���@w��s3,��]g�z�|� ���j�(��o�z`��j�tU+.��������|� 6� �5H��]������<���tDr���,{A��lw�ݍpXs�v��7=����u��H|� <b�5H�x��yWTqeU��UT�Z�7�3<�D%�P��V4� �<@wͪ@��N�����׬/0@|��@��|ڤ�f�߼�m><��crg 7��|ڤ�@|��@o�3u�"�0`�����p>���kӀ}�� �����Ee����`^e��N�=a�$81�FM;�[=���̚ғ������'#qϐ�<m��}�N���b |� 7�T��un�*��@]�{���@}�� ��[j��1��f�=�5��#�P��� �n���}Ö��"B!��b(d"0�
Pˈ8�
H+���&���o3���=�l��>�Nb[j��1��R o� ;�Sl6}�Lo���7}4������l���g �b��Fؙ���j5���fʑ�䞛���`���F�=�\g�[k��N��33cdH�M(,L�@���@���� �b�n�e�{��~���e ��[j��1�{y����&�jE4`��8wZ�}�EW���� ���p��{�|�I�M����p{����o�����AT�<�]ߧ*�~�z�N G�|�� ���� n�f��ŀn�z`!(R��*��UVL��5��c9�x��E��M�{��m������'�"gs32g>&L��G��s8n�@kmR��J��_��ۊ�GE;�X�����8ww��7}4������l���M���#�1�bnb�� ;��@���� �rǏLSc�ō����=�o3���@kmR�j��wk/fx��ae�e �>�mh8���R+�P|?``h$�5�?6�����k���2 Vխ�V"�Ω��y�r��k��@���x;R)(��v��O3l��M�vHI�ñ�ĎM��M5Z��Jݜ�Sb4�(v�Ϯi<�5���Vg�!�޹m7���n.��52�8��Bj笞0k"nZ��x�Vq�f�nJݹ�F��P����[�;H�f���z�X�&�^�#[f�:������@��3���4�J6��;� ��i�ۈ�q�$��!��P9�nuE����L�0fHؤLCF���o1 �5H��*�@7�R�s�~���v���]w��o���j��T��ۼ���{�1I�G�brg �sT�o����H��@uw�)�wXe��aE�R�j��� ���������(ّci���ڤ|� sT�o���WXw����;��b�����Ch��D�Y1������`u���mv{
j�����7��H�wc�T��ڤ ���q鑦���s8��{=� �H�j��T�l�^�=�⋫.�|� 5�� �5H�p��L�ؤL���I������T���b�j�{�����v�x�=u�]� �?6�4	T����8����-p�$0 `�OL��k���g���o&��������և+8n�=�@e�z�y����b�j���p�o3���A��j&V7��	C!�׋9(�Jd7� o^,~�����3dQ��NL1D����y�w�Ò��
~EO�w����ʾ���p{f&�l����$���7}�� ���|� 5�� :>�:�V_�������R�����@kmR﷙���P�mDF�
$�O�8�Iq�m��\�>0�G/Go��ײ�I"M�I��~2�,���T��ڤ|� =��\���&�jEL0`��ڤ|� ;���|�Ox�p/�7~C�<I��ݼ��?j��p��3�{}��N G�brg;��p�w�{wq`Z�ZD("}���8�����o!�E����ڤ|� _? >�;.����˧�cw87$��N
J�-�&�֞s�9�K�җ�7N�i1Ӯc�� � ��� 7��)7�gЏDēs8﷙˙�$]{|�$s�� �����Y~�����@>�~@����H��@{Cw�	��I�qpw�8wZ�|� ;�����wW��a^����1��H��@w_? �⫪�E!�������j���{ qVgIZ�������#bz0.&[mbW�ێ���#�n�{u�;;��:𳲐`�kqv�E������q�Fw�lL�J��Ӯm\IV�tTK��)��I%��M�X�!z�����ԻAm��6�b�uZ�v����80��|=�rY`��X�wi�	��O�a�d�e�g�3=�랚�#yW��۵��^���T�w��ذ=2�u��7F5�W��d��<;�N�e�S�)s���q84�Ong�?���3�{�ڸ|� ͪ@s���2�^ta�̤���|� ͪ@7�R��w��e�a������|� ͪGDBJ�z�`k\���n���fy뼤��H��@>�~@7��p{f%�l���Ș�ng ���8�ߪ<s��*@?�T����`R':�:M�f���Kn'@�tgfuۖ=m�<Ϣ7B����:�8v�@��˖�ϯ���T�6� �5H`ݬ�jdcXӋ�n�y���ϳ�09!��R��R���~���׳2�`Quy�H�j��T�}|��o����@c��pĞ��w�������T�6�>�=n�,�esJl��K~���q
!7���[�m��-��qE$BB�|��q��+vnGG�f7Sn|��[�%������n��XQ��R9�O_5M�ʧ�s_�}E;�g��ay�{=w�O_5M�ʧ�sT�<��۸�������&�3w�37߽�ϳ���$�LTMU���<����e��|,�
��j�fcyP�$�C6��R)������c$��b၁���Q��U�X���kx8�J�vI4ASF�Rdf�d�&&F.N dၘH�
�LHK(X,�6Xy�i��}�/����f@&MH��,�~�я�
#�Y��洂��%BV��sf	1>�F:4�H��4M@8)00MM@L�@L(P���&f;+�X�0_O��v����C�?"���S��:��!�����D�:~����xqiJO{�x>@#J]}����y�5��Z���R�P��������{�xq�);��w�� ��{�xqJR����욛�f��!$��^b�!;߻Â�)I����%��~�)JP��~�|��?�����Y�O�43�m���%1��m�����j��M�E'Iۇ��uW��q���Rv���R�����p|��{߻ÊR�/~׊<D �M�ő"B��X
]�޶f�����|��;߻À E$�@����"D.�ز!BO�׊<D �[/f����f��&�"��BR�=�߻��R��~�)JRw�׊<D �M�ő"Bձ�k*j�ދf�Y�s��)���R���������{�xqJC��U� � Rq�@�A�	FY@�~��w�����R��zG{��k7�����Y�o�R�������!=���/������j>�h���zE0�26ܒ���D��^���d�m�y$���IڸSZWp<�^t�/���=��;߻ÊR�=�߻��R��~�8�)I�}�x>JR�_s������f��kV���R�?{߻��R��~�8�)I�}�x>JR�����#�3�hn��jA&4qG9����`)���qJR�����|��;߻ÊR�?{߻��R���v7���n3Th���)JRx{��x>JR�����)J�����)Jw�w�R���}��)wsUsw6�n�x�A��fD ���������{�y�)JOw��������Ͼ����$�i���a$� f�n�7n-�[��ѮaɊ,'-�+;u��z��e[^#p�#�5۷<��*r"�!S�.P��ؚ�I��bku���yS[7�N�3>H�.Z:�AN��v�CQ�3�6zc���H�����Lq�Q�̓]t=�̌�U3�'������O��ukD~�t�	NR�l����@G[d�e0p��lA�cjZ��EXF��ꮂ�r�p]�q_�^�lvMmr���ϕm��Tժ���qsjl��=�!��}�<BR�����)JOw���)Jw�o��)>=}˽�����l��7�p|��;߻ÊR���w���)Jw�o��(}�����)w�;���Y�o7��o5��R�������JS��}��)C���%)N���┥'�ڙU-\QuJ����(��!7�̄�(}�����)���R������<D �C��XS�&iUY*���"
R��}�x>JR�����)JOߺ�(��!7Z�"D ��}5RSue�)t�j�*��z��^��Z.t�8�h�b{\e�����~��7�|U���ԥ)���R�������JS����)JP����JS����tZ���ֈѭ�g�)?~�{��7���1!�P���5��qJRy�x��B�޼Y�)���6�
z�n�MD�+���"D.�}9�!����Q��I���@D ������R��;��t��f���[��R�>��{��R��~�n)JR~�����)�����)>==�;�Y�����ܳ|��JS��}��)I��{����{���R����{����߷���߉qf���N�s�#���G�������mǍ���&'�<�k.��ͫ$���o5��R�������JS����)JP����JS��}��)I���Z�-�F��7���>JR���qJR��}�x>JR�����)JO߻��|��.���ݶ�Fky��o{�)JP����JS��}��?�/��~x�s�������u�s�R��_#uئDۘ�8���}��>�-�NKJR~�����)���)JB����Q�!B��1<�7wwHT��̈A��ͼQ�!K�$Gu�ND �@�w{�G��	�lȄ!j׫�������؎�>���{���.�r�x��t�'c7Ol>y9�P5��z���|��;�w��)J}����)Jw��n)JR~�����)�w�5���ѭ�֌-�y�)J}����)Jw��n)JR~�����)�����)>==�;�Y�����ܳ|��JS��}��)I��{����{���R����{�����H�m��o{�{�a���qJR�����%)N�_w8�)C�����G�S;�;qJR�ϻ�Z���������R��u�s�R�>�����)Jw�o��)<�����)}{�Z֬�kVtĞ8�]���j{3�su�׶L�V����\��mu��;N�!�9sn�თT}�v��m���~��JS��}��)I����%!7Z�"D ������m\�U��+9o|��JS��}��)I����%)N�_w8�)C�������K��h��{۽�[��)JRy����JS����)JP��w��)����R�����:Y��o{��F����)���)JP��~��JS���qPD ����(��!k�M5WU%�/Z0����(}��w��)��}��)I����%)N�]�qJR������	�k��` v�9u�ګ*h��6�hW����񱶃`�
�i�1��r���0��7K	��8�t�k�9"F����7�F�z�w�ܔ{:�*��H��T��籣�m�:�<=%�X��g��z+���lE,�&ț��ZGoQW6��]��ƺ�;n7Op��s�S�I���㗞�`��t���3d�ƼS�/M�qΊd�%����{�9xl��!��3�:�nZցj�s��۱ݸs�ۙ�>և78#\tk�~��8?�)O������)JOw���)Jw��s��\������%)K��+���仴J���"D ����(�B!)"uwND �@�w�b�"nّ"BߛS!MZSU*n�sW����{���R���������{��qJR����x>JR�_s��f���Z݆�o[�)JP��~��JS���qJR����x>JR���qJ�AMu-��ڹ��D�S���(��N���┥'����|��;�}���G�6�G���D�Z�YK�����F��gu�\�Äf7��Lv��t#�e��z��c8�Vv�g���'n�}�t��Iw��G��	�nr!B|��"D&ݳ"D �����s7wuq3F����)���� �J����JS���qJR��{��|���-ʩ��꤫VU*E��D �@��x��B�۶dB�B�$����أ�B��]ӑ"Bߣ�*j�J��n�f��p|��?w���)JO}�{�<D �[��r!��BI(���Q�JR�t��쵽�5��;ֶqJR��{��|��=�_w8�)C���%)O�w�8�)I���3��Q�u�Y:[{�ظ͛D<M�-�Eɫ��s'�gb�C�=[\���p�������m�w����qJR��}��%)O�w�8�*^���"D#`n��1TM\ʥ��y�)J}���|���)����ÊR����?�%)O���8�)P��R�]ͫ���M*��)G��_{ÊR����{��C��0Ԧ���8�)I�߻��R��������n7�4kz��)JOw���)J}�w��)JO}��������xqJR��O��gw��ozۙ�{����R����n)JR{�w��|��>�{ÊR����{��R���t��nټѫ�u�V�ks�$�ķG�����t*n;9��u���G%f�cr<lV�������߻��R����)JR{����PD-t��B����2�L�қ&m\��9��R����)JR{����JS���)JR{�w��|��/�%�����Sw3*��D �A�ͼQ�JS���)JR{�w��|��>�{�"D ��� ��ET��B���Q�JS���)JR{�w��|��>�{ÊP���$�F��H	�`IF�$dH����`�`Y	`��& �dE�e���H``R"($T��9�����)u�Ϭ�v-kV�h��y�)JO��~��JS���8�)I�������s�"Bk~�c��n�nEu7�݈@v��m%�=��-�n5r�q��thM�^��SF���'�4]݇#�o���{ݷ��w���)JO~����)J}����
.JR{��w���R����9�7����ѣ[��)JR{�����()"��Y�!/���Q�!B��.)JR{���Y�ٽ�5����|%)N���┥'ﳿwC���N�ز!BZ��x�A�^ʩvU�֭��F�5��R�����������dB��ߛ�"%Р����Ȅ!n�&{���R�KW3&^e(�)���8�)I����%)N����)JO�w_w�JSg���2	���1�+�_~�_˅���vf�WyU�a!!�3��LrM6VRR��$��@A���D4�1�!���P�B
�Y���~X(d*%��)A&�x	�8`�`?8B`%	HI%b�bS�@dT����xA�IWE� )�"׆:�E�����ָ6j�>`6�o18���C��l�y j@Ȇ2�Y��m`�K�L�9�8dfK'���]�~�?T�$��"i�Y�s5�Ua��KA-+-4�L0<$�<\	~DC��Jb��|�6�;�x=�4Z?���b�� m�a	��(fq��}���Z    ��@ 8-�Y� �a�C�           �I�z6�m�t��k���.�+UU[m`u�`��9�ѳ��m-8i*�4��V����i��ݍ��E8�fNՕX��h
�[��� �n�2����E� \�C��	Q8�XY�mN�:TO�/_=��R�t\8�f�X��ʹ�S��^�vx�\�5m��=*�B���8^�h�6��+Hbx8����L�ڒ.��z'kH/�Y���EYWk�kv��l�]v��][��lcJ����+ h^ˋ<#�����V�Ѽi��[k��	pm�y�oX�Bi��pc�%VG��[N���q�lS����G\���)�il�Wu�Md��%��[�`�I37P�Z�B; $�e��v��-�.-#�:
��ה�X�Kz��iЉ�"��HuT��L���[n�J��s�D�Kn�V8�4�s�^nK�u��{!ns�$��{rg�24�ĺD��:��۴��H�U�.���;r[-���@����26���g)�.8@8�Z�@����m۷R���.�Q0�0�����U[UWT�g\ h��67mb4��ڻ쩌����l i�M:t��	�H�U*����[�	���^9Pm���<�r�W5��@ݕA۴���L����^'3��X�:*�#�v]�5[�@�m�g�F�s$�bbG-��qlYy�SsL"�j�ʒ����ۃ�m$n@ :8 ������i��UJ�t��{A��xȵ��i3�m�:q*����ҭUU[�g��zy�"�N(���Alqӳ�I�r�+v�XϾ/����H����m$�9�v�[D� m�u��C�P�r\Fɶ�
����nz/�TZ�AA�lݖ��n$�۞�������.���४�UV7`��+s��@���nB���%��J�<��]��F��v�t���gWs��zvͣc*{T�_?N����{����b���6� �T��&��{�_{�^�������ƛ]   ѥzst��Wv%��g��ո���vۮ�S��*�����m���U�g`ș�w5�dٺeS��bt�1))[N���{n�!�N�^�),���}:�:]�|���v+v
��r[�&N�rR���R5Z�2K��9Ͷ��1��Dem�I�ś�`�F8܍M��$��A�Wi�<F����=���W�S�����΋u��n;���3�&�эݚj�&��Ђ��.�v�\ù���۸y#9qGUr��`�����WUV�!B_�}أ�B����┥'ﻯ���)߻�R�A	���WpU%��]�"��bK���D�!|��J�"7�qJR�߽�x>JR�[����bֵa�Ʋ�l┥'ﻯ���)߾�)JR{����JS���8�)_g��Z�S"i�b��Ϻ}��e߻ÊR����{��R��w���u�Tx�A�|�<�Ue�ҫR޷��R����{��R���)JR~����>JR����┥'��ʏ͇�%��wj�5�UH��<��Y'nW�LEIZ�	�T�����r���)Jw����)?}���%)��^,�A���x��H?K٢]�tU\�3J�5k ���צ1B�!$$!%!	T�Z����ʾ��{�w޼Y�&��g��j�%Z�s2{3+�sw��I��@|�9� ��r�޻�,R$�%!�=�����p�f����y��˥��.�K�"���t� >�{@rEH�&���wقs ��jh筙�vm�]۫�8�@�\�^X��q�-v���㛷!���6��8��tAV֭r)�4�	�1>p�v�8}���k�f���g�(S&�8�Ue��"*��X�}���ن���!f{~�:����e�J�7�&�$��8��چ�㊐u{�&�'�LV1��"x�Ng ��M8�����oz�j���݂RIB��B�L�F��nNln9$���4����B%����C�'�Ȓ$����g �M��<���P��,�^]g����{.��M��<���P�#ymʰ�&mᄒw�_;W ��P�#y�tP݅���=�x��@}ͨh��yɺ~��Sڸ[Z��LQ�`����9��t	��w5�=�,������k�0WV�Qm��wP��W��W6@N݇����������R�ݞ˼�t	����4	� ����A+"m��'#���j������)�;��ށ�]LV1��"u�2���jo �ߤ��N�<���ȶ$��S"X��΁}��zI�����ր�2�̯{/.�X{0@oI7@�ry����#�}�W�����H��{�Ow~o�����YSm�  r�V�kL����+9�$y�F�������.'��Kdz�љ��|Y�I�d,��آ:��ޱv�:ٕ W��s�b���9�kP�P�7N��vjG�Xr���C[��� ET���.�D��f��[�^{]
�ksѓ��!�įSE�3�0�vt�H����V{mze��5k�Gk�����1v�www~�{��p�s���=�[�W�WW&GD��UЭƉSi��oh�9,)��ã����>�#�	$��{�.�n��@����$��?ow{��]UԪn���U%���ۯ��2sw��{���Z�U��^I1�H1�9��e8t�t	���ͭ��A��3.��Eײ�@w�M�'[�@wt�Z��p�5P��I�'#���o��&ց9�}$�WIv��^��N�UvL�띝FTqc�&�=v2{Z��⎇ʶ��!Z\����>�wt�Zo ���&��O '�$�8�"X��΁we9�������W���M���k��$�G=�]ueU�{=�~���������s��sk@��N�r��O�����I;�?W�`}��/�m��Oﻻ��99tL�<J1�#)"����:��v�������ށ����_yA����;�0�(q��nzq	n9og������+��C�ˉN�m6:e�8�8�I�@xٍ������l��ny��mhG^�=Y�^]�����ߛ~�BJ!D��S��7w���o�S�w٪���7'�x��w�~���&֚�]��A��n�����a&xqp{��:�e8�Ϳx:~�}8i��뙫�%�j�T�fր����t���wI��n��?2��\Y�a7G`��;��-[��gs����n��m��n.�ßZ:�v�l5�w��{0@}��t���w9��>s��6�TTI�6�I'z�����mh�T�ߤ�����޹�{,�⮽��@ws�Z� 7�&��ڸZ��I1Ln`�s���̄�%��,�����ֹ�k�~Q{���t{qS��Ȍ&G&p����}-� ;�ͭ��wp�^�xK)l�����vƏc�p�s�'����{n���ȁ?�4�)ړ�5#���ڐ��ր��H�I�ޏ��L2�2�.��� ;�P�8��I7@�^��/��lMǌ���xt� >�&�Ks��4	�諗�Ln4�D��������\���t��g �sVTI�F�I'z������t�t�����߷��J�[$� �t�=x��m��v:�x�B���'[<������~�=���fcb��ࣞ����*v:�a��u�)"\�5ʹ���7-�+�8y�kcRP���zwd�އ��Oc�v�s�ix1�lu��9#v�\�&��m;n��#�f�s�;��5�8���d�[�M��]�U�㞙�u��ěD1ڹ�}L�׹�ߝ���w�w��+�s��c�3m�L5��Sή�L� ��{��C���^J8�\�LVN��fy����?��>qR�n���<��Q��&)�@x�rqtݔ��M�>�'�����u�/x�=�u�02��M�>�'����=�8���%a�bI�R9ށ��R�������t��ޘe�ve�fy���h�1�$��s�!(�޲�M)겦mMȂ� x��1�䙱p����s�k�a��ث��Z��Ȝ��I�K��/����;�oz����lںWp�\�m�*UsWx�m���&���� ��}> ��8ەarO�6���I;�?W�p�{@9��&���g�r��8�ǉHp{f�����;�oz벜�F퐘Lr�������byɺ����x����&I���mnݮ���3U�P���M��������m�u��p�|v�t�Om����~����� ��޹��	(���Ӏn�������'�r9ށ�� ��9���M�>���za�e�⛚Rv`���>~׋�k,I�� d���P-I3D�w0@mƕز�K$,�Q"H��)ÿ�?���PS�Q$D/����~y���w�@v�HJ0�L�K�2��$�,&��]H�����0�2�82I!IL�*
� �_��@'P�� ��(�'��8/�Q���gށ�v�}ށ����"؜���$�Խ�>qRyɺ��s�=�O[�:����s ����oz벘�۟�kŀr��2�U
z�b�S���kb76m4n�k� �'�	��`���p��&4)�a2L�yI'��{����>�4�*@}�M�	S�˻������~��e�s�� >�&���p
���0����Js�@�qR�rn��y�ↁ�נ��0�e׳�Y^��@}�M�>��s������m�p�U��ƤsO�y�����qC@|�����������B��ײRZ��mg�\;�qÙ�I���MǞ�'m�rZ�*f�^fy�8��>qR�rn���<���j,���X�ȅxt��g ���{W ��@��1��<32�z�s�t����ↀ�Ŝۚ����<0�N���\�C@|�s�tT�޹g���/<W��y��"����H�&�������Y	H�Jb����!0�� �W���}�o{�f�v���}�2V�t�[�����N$9�8�u�T�g.��mk�O��	�lc�l1��g�1�s�e� ��9nF�i��A�m���v7�ۣ��{:��ԇ4[�q�۲��>�;a[���05;F��6�r��ϵ�ێ��6�ncu�ns�s\;F^g�&jT����]ub����nj���s��7F{^^;;��{���������t�%.4��v�C��EV��m�l�ը�5t$�6�'1�W���	�@x�58P?��R�ɺ����E��C�	Ǆ�����=�o{�~�j����@�m�p߳U�5#�,5#��>���(h�T��n������6���H��o)�7�y�޶��~���=��"r7$���j4�T��n���<��CC~߶ߒ�\�<T��z1���[�4k���wH�o]��0�Xƞ=��r ��j�͆�m���ה��n���<��C@mŜn��˒`cc���I;�?Wj�Ϫ�U~��RG)ƀ��H�&�����Iǋ#&,NC�{��wo3�{�����p
���0����yiW����&�7��}�i����H��'ɂ�g ������ ;�P�qR����]Ox�e�uq�M��vFy�^θ��z3��	5�m��'h���5#&!�Ԏw�~�S�wH��6�t�t����L�]������`��C@m�H�&�I)�=��"r7$��S�:��g*����yx�� V���{�ܫ���:Wp�\�H����{���>� ��C@s:~	Y�v]e�Fff�I�@wH����޶��{�-�8�cȌxdX�F����ͻ���z�N�t�������#��1k�<܍H���1br޷�����=�oz�e8Z��!0�����hnb�I��d�(h]E\H�n0�7�޶��~�S�{�� ��8�٪�T�����e���A�"��F� _�W���7e���2���1��A�� ��P���t�t	� ��.��h�����3R���v.O6��w�ri{7lo��L��S����F�߭����n�:d�M��:*c�r�	�I�=�oz�)�=�os��n根&<o"�	$�#� ;��Z#���n�J"�;"�ᑓ䚐�����v��[{�-�NV�v�L&70x����	T��n�#� ;��Z��������a'HM��  6Fc8^k���WcZ0-��կ��ݯc�q�b��e�u�3��μ��LI��Y������v��d'eXkQ�޻bl�;ֶ��ે�V5J����[#qHELIgB��xƓ�<l���I�;*qm��v�m�9����F���x��Y`�-�G5V	���r̎���˶�m�
�w��]�A���]�U���SMZ�$�G��:ƴ;m`M�F{/O.�����<:���t��Y�-QJf���7{����`|�����p߳UX�$�|Ԏw�[���$�ɻ��^��,�~��jf��$�4�8�m�tv�8����[�����+	$��!9��8����t� >�&ր�86�6�'�ng ����vS�~����׋ ��⦤��*�j'n�)<��5����kj�7]��[o�c%�3�T��Z�j��T�P���߀�w����Z�*@w97@%�us3ٗE]57f��ߗ�$�(�J#�P���������p
��k�<&I����Z���rn�:dt���?n��$H9��JI�=�t� ;��Z���ꞁ�e����
�g�7@�ry�$��#qR�m�@��[�qdRD��G��$쭹�]�ѹs�6��ק��\sq܎�>�rdA�K=���uffy�$��'8��$���\���'rI#�	�1';���M�'[�@wI6�� �pm̒Li���=�oz�ڸw1/޷�΁|���sqe�>��Xa����8��<���%
N���t��?�PH�>h�.��yN�|����oz�ڸ�)T�1��={v㫰�����d:H�x�{V*�(��9R��=,j6q��	�@x�Np��o��t	��tj7�y{�ay��?]��fy�97@���5��\���kqĖO�(��@�܂�C@��-�97@�Y=~�ʍ4����I �뼧@��_ ���+E7)������~�3�y߳P�$�c�O�;àU�{��ށ|����yN�g�y\ƢS����hv��z�g=nN#�4��.������}h�pH��)&&�E#�����_=�@}Ѩh���~�Vg�ʻ������V��S'��8�:���k}�ʑ��G�&LbQ��?z�)�'��@w�M�'[�@Ow�w3�FU݅*�*�0�rP��_V�>�x�m\���ۨ��RF��x
G�;�&��A �ɵ�Os����ﳯĥ�	w>��fd��t���[�m4�(d�m`�YHHF8[��)�A���դh `(H��J�&��*�[���J����5����֊(+���T$�M)Md5H#�PQ��DME4~���Qn6}�f��"��l����'iUT�3�����4�\@<��9@RP�@R�C(7�%16!�/�"n"���#CM�D6*H�E645MfeF��9�U9~ ��1��l3Hh_B�i�J�|���BPU$�l̲�&"�̙�|S�_�`�6�oz��kf���{�   ��@ i#� kX          �l.<�/
�V�<Ut ���V����ɶ.�e	hT��5+v��(MGNcT��[�=��I�9�ǥ�Q,D�N�̝���kj�V�st�"�+T����.X{<W/U�����a�WA�q�s�Nd�����t��<OCJ9��ƣ*<;v�6x��$͵�d�l�T���f��3�U�	�g'j=�v�[3��f�W�s]�:��O%��*һ6����.Z�rUմ1�u*%R��;���ګ[32�� I�e��l�"Y��Y`� ��<e!b�d�@,�"I��t�ܯ%�i�q�k�U١1dh�v��T6�:�@��%�Y�;t�����k*��`��ss�s�bZ�y*�M�s�(��WQK���v�d��'j1R�l�Pq۶�r��l;c�4���n��^�,�̀Dyi%;m#lm�;�1C��h�$24��\�@ݬ`rԫU#�oIZ�|Ē�q�Y:�qyA�^˪tf6,��<�t)m*���U8�5j*��`�F�"<0��	g��ەT���ڶ�c��mS 9vwd�]�������	� UK��`7gmN۲*Ҫlni�v�۝@Bl5uU;ny��:ik���;�۶U��9J�{m���*���/X��b(����yyC�z���{u�:��x���<�F����&�8��.�r�sJ�U�"5�X�Um�㭛�I$M% ��N�[�Y9��8����ݓv�cf�g����<�CN�EĽU���J�T�qZ:TU��"I��޺�c��#�b�����@Z����;k#V%����lH��  m�RUmzܼ�0	GR[i�fL���@/�Ib%U�d�N{�=�,�[v�8�J�8U2>�m��@�[Ru��[��Q*����;c釶ܵp��8���yjs��G���[I�-l�޸�#�L�jM�@	�8 ���Ow���{۹����g��T�m&  FK�/kr��TsvmA^m�s��@nמq���k���񬝸㢐y����cp&6V���Z��lT�KN��i^P-e;e׫�:{�f{c�*�;nܬ:ۭݺ�0x:x
��T�Ep�ss�=N�K!R�i�mEɐ� Up�u�G���*��N�^t�T��!�$A2�	�źc-�@W���,��8X�^�:��37Pl�ۤǮ��a�\�t���l=�����<��h�s�4�F8�Q�R^�m����{�������~���w#M'1D�ǯ) �ɵ�O7-�rn�:EH�tI;�I&(�s��*ݯ�~�M�>r*@>rmh́32���ʿ]f{2�G&�7 96��۬�kT���)U+�"�����ŀ>rmh;s���t��_��zvz�=����X�d�Zki<��p���t�7�;����V/�&��I�5ق��w�m��g��ց�����97@|��x�w=H�waJ�Wx����8I/Е���H^�>������~����""!L��N�&m]]��*�����>�x m��o���@�{W ���k"�C������Д��� z��������}��N�hi�1�9��{�u���ɺ�@>�]׮�/�6�����͵�l���pͽ��3[mm����rE����$�"rX�
w�@�{V��o��Z�/H}�� �Xwx܄�cO�$\߶�����w���j�}���'�CyG'z� >��4�ߪ�s'[�@wG7@��qWw%\ͪ�j�D$����<���|��s�����.��eez���ču��|��s��z�)��*Չ�9�3#X,zfm�s[ۈGh�F���5��.���9�����[*B����%"����ށ|�\����ڸaCk��M<QIށ:EH�5;s��I��+�:U�3\����SSH&��7y��k�9(��w������� ���&��*�W5>��ǳQ�t�<�亂�>��~�~�qIB�n��x��ݪ����Tҳ3<�亂�>�tjKs���ϳ�K��<�4��5�fI9fL�f��#R*mf�E�s���bw\�ͮ.玺�����ff}��*@wF��t�<���ozv�w�La�� ����Q2oS��7����ߛŀ9�>���HL������=^��=��ށ����=뼧@�Ck\JFH�>L����n��EH��4���sk��!��H�z��g ���U�u�s�{���U��Q�R�;�iZ�d�  ݶ�%�Oj�#G�&�x��v�t�s�������1ǅ�<��7N�`ݨ��� �5j��
��!3hk,�RR���FKv�)['��-�K�V$n�4��8���Y�UZ�$+\�z8cW3UTR+v;VKhN��{;on���3��=�u����Fw]tT��b`�8��-�#ͺv6z��b��h�+d�\s�ә�WF�����m��?Mqe�n���Յn.��Śg��j��B�p�����維�Րn�#p�m��@6چ������o��� =���ّD��S�:�ڹ��يM�����b�?|����wJ��޼�2����rn��EH��{��A������.�/������ ;�� ;�P�:[�@l�n�G.���+,���Yw��m��[�@k�n�����/ߪ4��n3rdM[�VKԣ�9��"mٹ�J�����a6��_Y�~y�VW��/ىKs�rM�H����%�m���93v��&f�P䛠N�R�jKsʀߨ�N_��0<_��fn��EHm�h^��;���ێ�'r44�&��)͵;s�rM�'H� ��ĝ�!�D�����u�\�m�@����=���@���1�r 1c[��kRfq�k�Xko=��$���{��.A'�ɑ3#Ĝ�	>�E�;����y�ۻ�t�j��5aa1D�nZ]���?�Ŝ�ɭ���s�Ӏ{[~�(�Q�ꮑUZ���SEU�[yǀ�ֹ�a+J!&�Q�<~����y� ���&,l��:v�䛠N�R�j��q'��E>lIH�v��@����=��S�]{W ��@�	�Q����m�B�A��3���4��,�2Gk�v�317�Ƈ	4c�';�/��p�yN�u�\ݷ���I܍9���Uk o^3ܔ)��>���{�?�Ŝ�B�2=|�k�Z��\��ͩ���\��G&��T��������N��>�E�-�{�/��pu�<�P��l/gW�N����E�m�0�����8���^��;n��e-�8"2LA�5*�;�#ٶ�mdwfĚ��\&봱��yk�Rщ���c����po���^��5�7@�"���u/��eez���č;s�q��'H�Ϛ��W�Q	D��ꜙ�ut\�U3w8�Ͻ���Ò��νyǀ�O� ��'�Z$?�H��@����7}��@{Z��%��s��櫊��Ss55j��Aw��o���������K 興Ԉ���]�vQ7S52�]��݀6�5��r�ֵ���5v3��pgk�67P��Az7;+���l�H�WOgbg,�a���p> V�k��9ѳ�N��%��>سf�1�(�d�]�}/n�b��"��rdZ��k%@�N^\�65���u)�y,�e�׸���y�� 7
� � M�a^̆'i�<4�0�v&��2���Ëv�=a�c�r��X+Etc�`�4U�Wi���N�Բ�0]�Mł%3��Up775
����o�>�������?�ň�o)�5n�;&�N(��� �7@�"�|�4�� ���V`dM7&�s���g ����ڸm�ހn�a����c����p|�4�� 6G7@�"� �9��"�dō����u�\���@����7}��@��Hj�F�2`��1��n�m��<!��a�y2Sճ�a��Z���s�����%"��oz��X�ی脒�!ΟN��.O�J����7�������� x �7��C@�۞@l�n���=��_�,��.��P�#�<�����'[���ۉ;�c��O�S�:׷����'H� �5����u�.��ן�3<���t����h^��7h�̓ƛ�_Q2]&luH���i�*]�ۋu1����7�}�|g�ȚnL1��:�������ڸݷ� ݮ�s��	������=Д�9���?w>��7� 7��N�� ����ڸݽ���>�݀���!B����������e
�d�� ��6���i	�ac%5<�0~hJ1��
\Y`x-��O�H9�ppT��K4T�!A$#"$~7h�Y����*pDL��_P���E�PD����IG���ŀ~����������Z,��g��� �G&��T���;ڸaK[B��L1�����8K����9���=�_�����]��P�k��Q���Ř۲�\vЙ�uӛ]����>E�ȡ��9����m�g�C@����&��'H�9���c�,o(
w�@���n�ށ}o3�[��遫t���7Ә��I��M�'H�#�v�Wf�ܘ��nL24�z_[����<��k��+����$A"XR�	d(U���o�?7MYUV��UY�Yw��q�;s���N��(���㛺�(�S�w���*�a��i���sg��;L<㲆5£lA{OG!?p����-]�T����������~��y�ݼ�@�Ch�"L�A�ؒ�p��� qC@���~���	���i���y�n�S�]v��m�@��!�6��yHP�#�<�qɺ��������4��)��ڸ�|�BO�w��7݋ ׯ�:!$���ʛ] �i�k����v�Trtfc��^B�;]Gg��cp�mGZ�5����kU�L5�e{3�آ�N	��x��;2�'k�K65��2�xq�3d�]�ZlӍ��k7bZ��N4<n��3�	tc�ub���*��s�G;# +�ks���;t���-�u���-33���mz�jCg�Vq�;^�۱��x'�����w��j��7%�e�A�t:{=O����4sٛc�I,�6ݧ����������p}���<)EZ��� }�w��x�z��M��=��ܘ��NL1��z���^3�|��5�~�BS	Hv�u�UZ��R�EV�ϳ� ���^�ށv�g 7���_)�L7�99àW����&�ȩ ��6��)2cX�lI8�ݷ�����v��p�Z�r(I���z�ݡ�v[k;q�˸z��OJ%���[N���6:c#lP�K���@�o3�m��t���6���ZC�,m7>t��j��^3�
!~�7X� ��x��8�n%r9�H��J!N��ܞ@8��?W��T�q��Hax��� �8��v����8ݼ�@����\n{7�14��Vg�7@�EH	P�#�<��ɽ�*Ѷ���☜1|�A�$��C ��\çZ�{�����g',h�L���}��Z�*�`��x����~P�<�y� �6���L�`�1��;��	��G"��(i������)2cX�lI8��oz�y�;�%n�t�]��w�������t�ȩ ۊw'�I&��ZC�7�n|�6���7v��np����z�,�BI~��M)����ݺ6`�͘�n��g��׏:��rׅ��;�y��>�i2��/���m���y�n����P��(��pmH��� ����ϰ.���ݼ�@��\n{7�1190�G;�G"�74��#�<��I7@Wr6�7������yN�uڹW������&�)�@|�k�������ddP5�99à]v� }���$Zr*@6ↀT���/h���ls�V�;b���Fu��8䝣��n�Y�D�go����	����?�N.����������7u�?��/�s���?|�URQ9����@�o3�n��:�j�����3}��5PIb� O �P��`����R�+޹�$Kx�'��p�m�@�o3�����@�m0R69 �������ɺ�*@>qC@���$w~O���k��$  K#������ku�v��[���L���Z�E �ǋ�5�C��;=�n*V�0�@�=:[����;nܓ�����WOtC�MI�����x]�t[�n��WY�Ѓ�ͭ���wm��m��9#rێm�r/]Mr��.٢^��8�vN���8z���Q[n��^�c$'�Y���ѹ�hv�'f�:�V�l�w{�����~��,=��i�Ş�t�k�!uŔz��Ÿ���ќ����������2bӒb�)9�?z�g �m�:���?]�� �W�#&)����p�(h\�@}��I"�_��t�4R`�cXc��:���?]o�:)�}ذ������.�wSj�R�&f�p:�(J'�}���ذ��S�]{W ��)���R`�������T�|ↁ���ɺ{�n��~3Ŗ񭽚�n1h�]I�Ͱ��ۍ�����ڱ��=�wt�����������@>qC@���s�t	�p��W#���cl��àZ����rR��u�{�v�b���e�!H�܏	0n.}���[���/��׵p���N���$ǈR���BJD�B�����:�gv��}������Ɋ|c� ���}��9(BP��Ӏv��xͼX�j)��(�`8�Xah�H3X��m4�+,T�&��ۡ�f1���1����� }\�z�*�4�O '97@�"��:��$1���ƒN.}����������P��<�ߨ��w칫D��j����,���ЮƜ�T�Up�Ⱥ4�����D�0i ���i�1Q�d�ڄ�`�O���Wd�����~�eLӛ�TU]
��� '8��7ny9ɺ�EH�+1�ƚ"�������	L$�v����� �k�x��;e��c��Z��5d�ӹ��d̀t�-���Gv.'�L۴ɖ�m����Nnn���R|��߫���s����N�F�$ǈNw�~��8���7k\�����dJtT�R� *�� �}�x��8
G���?[y� �.���a�Ȱ�'8t�_w9W���|���xr���y��}�M�/)�7Ci���ěIL���t���P��<���c��'Ky���-�P���:�����a,	�m�X��ݸ�Ѭ̥�̩#l�k���"�G4��/ߪ���I{�?*$�Q�m8�x�I���yN��Z� ߛ~��x�BP�\̵nb�%�4D'�u�\}m�@�m�p]��@��ahn�d�G��t���P�+�����v�sٸ���RI� ��@�m�pW4�� I7@�������W��������!�������5�8`�j@�R�2��D����¥{����H�%L?�@&�	Lf6) `�K�!a,I�c�!Xm����;�7��hVqBYB ��I �D�����
�$B���2���n��R�<K�H��!���y�kz��   � #��ǀ�   `        *�y�$�����������9絉�p�KkB;ƹc%�e���E�T��V�R :Iq
��"��Y!��W��m�C��o5�u��ĵ�mιG )�k6�8�H���֠�.�ƨ{\d{v�����2��±�2$��#3�G�u.�A��v��9��H��bHRh�S�t�q���ݟP� �T��u�vY��n�	m8�T��͔]�8���ڹ��]����c�P�i	P;dR#h H��5UT�%�͝@K,�R�2��ʛJ	�,�D-�'�.q�V�ؕ���UU�xy�yhM5�x-�mMp��,�7Sl�d��4R�0 �x���ܻ��Sq-�'Z�f�u;$A��	l̰4T�a��N��j�9�&٩؅^�9kBY݅��m�j��v�N�˛�]� �]�lu��3�O*�xZ{���[��K��$��m��咷Ę��V!�ؗ����խj�]�zօx�̡4[�j4m[RD��i<ʽ�RP`�Z�˳��+(pͦ�}o(�kY!y�:4$q:W*�vة|�<�V��m� �ISN�t�Y����`Μլq�A=nV�c���{@8���EX�O�����T�"�v�����S7X�9C����;n��&�csIU[�ٍ�V1��n@iL�r�UV�98�>MD����^�����Y,�Q�Izi$�(k�fT�e��6k�@hGi��
�f^���)*�J��UR���N=	���q����UD9-�1�0m�l�kkź&�D�]u6�m�lH��  m۶�Vmɵ�bLQX.��F�����Jk[E,�jj4=��q5<�&�{M'�C��¬�A�Q��ت�P `1�ݕh�
3m��p��˱�톧��(��b=g���	����5� ��,�n٪��i{]hֳv�������P	 ��"@��CH�����}G�|A�]���w�ڳz�k$� 7%im��N�l�z�B^9#gu��A�1��ѱ�:�D1�j�+�n���qjr-��L8�kr��Á�Zw��d�������k���u�i�G�6^��uah7U� ��}�c�`��q�����M�7*�ma��<�����9��*q��K�+�u6�:7Ss�@�ܜ��%W!��̑��v
8�4v{9�d9ة�����m��y�wmUN��'<�`��9�.���=�X�l:y_PHPȖ651O�p��3��^S�7ny �I�����Z�EH��.�zńf"���u�\}m�@��X�^3�(P���݊��ڙ�*g�����t	$T��ↁ%���!��n��&n*
�������� �}�x��P��6��?K&e���(q����=v��j��oz��8�ۭ�%!��� ykv�����m�ȧ7@�X�v��m=)������������J@ƞ(	�@�ڸ��ހ�x�G�7�g���WRUYt���k[�U���|��Q�"�x�oWq�X��3�7M�D$k媝�BRI� ��@��g �����W ����Vn'qFb��m9���K��	�M�?W�EH��-�X����Rs�@�ڸ����y���S�{u Q�5�	����V��P�.l9�5��^^%�5���W.�73���ɉ����JE�/���H���'��r���묯{?_��7@�EH�P�$�<���{�0?*$�Q��q�ng ��弫��{���b�
��_���|��o3�n�ĬƜ��'�����u��6�,O��8�Ow!G&'&7N�pۻ{�-���ݼ�@��\���c��r"Zu���!��h�rq:���Puϸw4k�K
f;XM߮��9	�m�cĜ�@�e8wo��s�(�;��J�5�f�Tٞ�ق[���6��;��`�SB��f"Ƥ��ks��st	T��ↁ�$^����ĚI8��ݽ�� �ٵx?BIj��sv� ��4�USu4��E�f�<�\�=�Iny͹����0�}�@�>�#	�k!y�ŷ&�:㶯Fl���oa]�t]�<�1�����I�Ks�m��Z�!�7n�V18lS���-{W?�)�[}������?Km
��M��M��]��n���om�r�Q?�_t��}8l�4;..�U�ڥ3W�$��<� �����7Z����jˉ�J|�B R�e��r��I.�}>[}� ��0	����C�b��T�a ������{�&�H  3LFq��'`'J�-�)�I��tw�0n-�j�{:��gs�\noL�nc;�������Mn�F���Q���*������n��3rٱ�݆��ں��vE�������1��K�UԤ��f�)�I�]��d'l;��u�7���#]�ئF\ƺ8��22�5��k��hWwn6�s��n�f��r�q�w�{�/¡�_�����F�Ӣ�����<:̽@n]���]{OG$�>>#Nӻ=M�� �����st	AW�\�=�z��N}$�M$�\ۻ{�-�Nݲ��-v��a���QH�?�y��I2s$����Iry͹ށ�Q%���1�!�C���-]K��m��?~�$� ��^Y��r����s�!F����;���ݲ����x����24G#���qS�'����^�"=�8�\�e�z���a�I��!5H��v��[���e�>΁kڸ��Lw'ѵ�I��j���ftB���B�%�Q���O����>��� k���S7�ː*�� 5̓���~��snn�#�p~�W�D��d�rqt^��9�7@���I��H�y��0�4��I��=������)�;�Z�׵p�ku�Ĥ�71B,C_H���a�i��>	N_=;�S)q����T��睹*5����@����e��]{W ����*$�؛�8�<I��v�������9���5����l�6�.+�'�����^��=��w�/!��	�T|�]����O��t���$�	&AA�E��߿Q͹��@k�'��� %��N��F�I1��ށ}e8�-]��p���*-k�.(��>�*
�Έ8A�O�vj8�t���]��4h2!(Yu*�V"n%J� ������F�䛠N�ߜ�����.�i\����� �m��DB�����p׺��f}�bFз�C��EL�U�����;f ��s�� ���U5T��E"j���P�S�P�{8�9��O�{���!!BP$����!�No}�yW��3��֍$��5!�.�j�vS�]���?�� �JB���SJz��*���rv��y�][um�܇9�{cǎ��z���Z�;���V,S�U�5b,�t���o�`m���S�]���?+��L��73�]���_YNv�W@��DDBI �5MT�j˪Wwj���h�A�=�F�䛠z�'q)�A ��.�j��)�m����(Q�x�c[��sVU��f^,^�'8�$�t	�*@Ie��ngۖ�I(<M�I$�I��,���-l�v꣸�0�-r�qF7\^S�-�U���٭�d���ȹ�s>8δ�`J�Bۣd&\,�67\�]�T�1�N��[s�q���b�K�z��@ֲxݍ��f���䆪z$�P]���1�Q�r��;G*�"s�;�8`r:�ck�n��*���BY�L�&Cj�ͅ,�cb���~��w���nݞ�����$�No��ěk-m9I@�7\��;��'n�:��Aӛ.�h�_vϺ���F�m!93���?���o3�6�P�/ �׋ ���U7wk�՗^����T��d��'H�%���K-��d�!�M�pl�|��X	D!�߼�x�֚��6F���_m�pm���y��-]���$�	&AF��`���?�BP$�%��� ���}o3�{�z�d��&,��_cdcqf�tۮ����md�q�q6Ô+�.��/V��$��Nw�]����j���8���j���D�$ bs8{������)�2 HJ��@0HC�C#YL"jLcH�TЀ'����9W����ʻ��g)�p��S�+�j�\������݋ m�� �^,�mπ��˜Rm4�$�}�am����g ��W@����;쪕�8ܘ�+��#qRI�{@�"��M�;ߛv����,�q��Z�L���h^k�J�ᶻ���v����q1����u����^u���&��m���v�g ��ށv�g ݹqX8��F���]�� m�� ��Xn۟��zЮ�	&1A�	���{�.���̙����'�	��6��{)$1�"q�6��А�0�L��k]<��� � b���6iZ ��Lc������ @�'�h}|���>�z}}�r{��m�p�7ˏj8+�^n���L��r*AD�M����s>H$�ng ��W@��Xm�x�ŀr�4��6M�M��`��
�3��bv݉�m�cAYW���먟#��Qj��X���eI75U*�2�݋ m�� ��Yݷ>X6V\�6�HRL��{�.����j�m�p�*�m�I&!�$�zr*@I2Ohȩ$�t�{ɻ��E��ҙ��X�Owgt�}��m������i��bp�#��^������7@�EH�$] �C[v��I�"����&�Ƭ�v�s��N�mb�����۫�����8$g��`z��7@�EH�$��6�g �Sq���2I1�9ށv�,��u�O��݋ ��~���աO�	0ƛ��;l�t��8���@�o3�L���x�i��ȟ9��#�R���ȩ�d��	��rY3j��I���n�xP��K�w����}���� �Ԣ� �B��($�A�ƀ���B!�0YSf��w�ڕ-�L  n�M����������rnZ���-�]�
 ��#p$�
Ӂ���V9�x  kT��[xD��]m�h�W\�I1]v��fڃ�~�k�GI٭�s8kc=��le�6tʦn�F�R�I%�γ �cmRQ�ۃ�+�{r/������:�g��<�]��#	0q���-��y�֤��E�ǝ�t�#C.�	b�,w��������{��{������c����:����
A8�Y��.hbn[<V�Lt����[���E�p���'&������;l�t��8���@����bm��`�&���d��#�R���ȩ'T�Lbp�#�C���v�8���L�y���W@���2IH��D��7@�"�ɒ{@�EH
n7�2&9&$';�.����Z��T�m���	 �Y��^�e�еS�t;���
�ݍ�g��ib��O+�ű#y29���	0Ɯ� ���+qR����A FT~/Ŀ�z��F�\�3ʻ����$Q�`BEF��@%Z+����m��9̂d�=�>�d���(���b�g �ݽ�l��>��QU�����s� ���%�7wjJ�/޼��?G2�$�����{�?*$�ؓj<I�Yj�ȩst�A)�w0��+=]��`p��՗h-q8s�;r)�5v6v����%��4p7���}����n�68~�<��`w_��l���_t�����$�$�Ģ '3�]ݽ��S�_�Z��y�� ���yq��.�I5~�]� ��>��$�	��Xm�xu�j��t)��E_�0@O�I�9 #nn�� �]CEhDm}�]�� $�=�y��f �;n|6�Br��ܖ[�ݶ���b�z/�9!�ZtI�m��v���t-Z@�Yc��U߭��n�� '�$������KbRI�xƓ������ـ_�Z�ݼ�wv��yT���܋���Oق}2Oh��st	� ���%�WDҰWVJ������Ou�ʻ��w�*��nW��� &� aF�U �~מw<��~�*�vw%�a5k {���:!$�;{8��[��u��7�%���������d4��l�f�֎���ls��qh�p�fqrXS1���������~�l!j��}��N��c��#qR�����e�d����8�6��wo3�]����)��]CEhY_I�|�^�X���!D$�?�� ׯ�7β���(�������m�@�2P�#qR~��zz���̯������;f %
!-z��g ۶��<ϳ�/�m�Q���$8 4Y�"l�Nʨ<��<FH�4Rb�F��݊�y!W��i�r-"9y{:�X�
��s�]����\\�ަ,\�)���W�8틝[G �eC-L��h��;	����*r�O$CB�L�:m���Y9�b����r�ێ�t�`m��໧��sؿt����ͷ*.��j���=(K�՞��.���s�u�s)�6ɪ"^w�w{����w�{�?/ݦ�19�{zv�4�ۓl��jS�9��$ې�N�^���#7~�o�����#qR�&��T�|�{��&����S5�<�x�""�5�~���`��<�
�]���J-X]� rn�:EHP�#qRSM��7b�1Ȝ�@����6��<�x�$�#^�� k��踫��W��w��q�7 rn�}o3�~��|��n������H��bk�zK������H�\n��֌�Iq�z6��w?<�ǌ�������F��M�'H�DDDB^�g�ߩ�쪹W73*�]�R�&�x�H� �n*@w�j���H�!�hI���y�^�g��%u��5�~�H17s3WH�M������Q	D�}�<7ذ�oz����ۉX8����ר�#qR�&�8� �����/�-�gW`:]Z��D�n6m�Y���۷ہ�=s<�����ww�������`fg��XyH��H��(\��� ��qكpmE"����+ ��3@q�H���߿W�� �j.WƉ0���p�yN����9z
+) �����u����5�� 7�k������"�w�xz�`��xz�`D%�6��:�QX�FD�6���rn�㊐8��8����]�*������]���m� ^�u\s�آ�G1Ψ��F�<���<g���qR�4T�qɺx4�f��M���*�`��<(J!@8��M�qR��L/,����xz���h8� �tT�q�g���B�WawqR�V��X
(�k���5�ŀk׌�tB�"WK�,�cU�VYVU������k׋ q�� rn��g��U��#c��'V�3�2;������X�����]���&'�$�ɸ�ǃ��6��<�^,^��(���x�~���dm}Np��y�n�ށ����6��:����,�$�!��-`��x��X	DBI��<�_3�w�j���H�1�i$�z��g q����97@�L�����.˻�� qC@���M�>���ʾ4^(���Z:N��	�奍���#��<�h��/�z�$��o<� pw��}〘H�/���/}�'�
�(��`H&=����\bX��jBhĂ�����b��`F0��5�KN�.fI>"��z��׬N���qQ�U�eI�q�x�m�B�gᴧ�m�"I�X)������z��� ( P X-�� 5�      �   �UE�Dsɋf�5���+�����燬;�� �>��:+v]�Vb���h
^oY��҇��(�k�h�I��Q���$NĆ��[KlKwI+��$ɡݙ�]��H��DY�]\�,Uv�^��T��L�S6�k�(�0N�ayT���n�9y�S]+H��&�2�iΓ�Wf��ͺ2�F�M�e�e���ڠOoB�*�@J�O#u<&�6�����A�=6��� �&�d,�hr�P9�z���B^�pWY2�)�Ɨi���Ա:�F��.`��*�)�uUT��e*iI��ۦ��*[��I�^Y�D�jH�mp�l]UK����[�r-AK,n)Rۮ6tU�d�m9��d��[Q�᫊�c�\���[nV�v�^�e����X��u��\k����7�ǙvP��d��
�WLW+��7* @�Z���3.�Ke�Ef��&�N�aWZ�n+oIb7�^ �Ʒj"{<i�,� ��T�5Nf�n�8���4a���Y; ��e1�ya���V�	�]����ݎr�pl)�*K�I��m� ���7hV���(t�I�:�3kJK\�P;�غ��� ��J\@,��d8`7=5�>�n�`�,��z���<r���&#nlgvۆ�8G-T�뛗k9a�mE�9Ƕt���UU�ȓ�R;$[Umr�1�#�^W�m��K��8�^U-�jes�S�+.P&���)����YqIV�U�Z�Re��C�Y��jyZ��McS�^"���9d�hK��հ.��Ojv�O���8��
�  m�[�k&��mUT#�q;�xM��__m�;G�f)eX
�U�eBn�U枪}S��Z�[�.��(Z䕥@�.pݷ�h���\���*�rkl��+����/^����s/;$b�b��\R�9V�v��ލ�Y����o����<��QqD�/ ?��|�+�S���w�}��Y��k��  �X.u�ܬ�����֭�{/qL�z5䅌n���v۷]����&��gl�%�C����9P�ved�ٞ4&c��<V��	��#-j��[:V;(����7(�'��Իd�ls�Ŧm���vx:�-�c�������N��\O��y�
�d�^���xjf�H���v��#�bz��nռvP*����߷����p��mYt��\l.&�c��\�� ������v�m�� ��@�q>և~���������U5VJ���@��ذz߼��3�m��t�i��FI!�"&	�����D%#��X|�8�=x�F}��`�n;�BI�����X���"g��Xk}����Ĭ&���ng �����g ��~��(7� ��.h�W51t���<�x���v�߿�� �m�:��m�Q�|���'���i���6=�pܗt��ۂ's�~�r�q�˚:��3tQ%U�����z�`��g@�o3�w��1)�<M$�����g�CP�BN�(P�9�g��X�u�ܡ$�L�'J몪�U!TUV���q�׋ n�x����S.ʺ&����S5�<�%(]ϼ�����x��^3�~m��WE����{�yH	���$qR|ↁ&�g ��=���X2Lm"Ff1&��g�%Ũ�2��en�w\�1�k�aˊ8.���[.�E�bs�ݼ�m�:�y��3�/�oz׊��2ܘ��nb|ↁ#�����H�Q���QYg��31#@��H	����̣z�!��BP�D�9�%�p���tz���,�`�c$��X�!A
����ϱ`��g@�o3�w��1)�<X�9;�$qR|ↁ#�����}���=��z�uݦ����z�����rQ�<�ttρ��0O}�����}�<�.\�R|ↁ#�����H�?��j������bf���o^,铵����}� ��<�؊�t]�\�36yH	���$qR�D��G 4�Nª�.��D������� �g�x�*$�Q���_����yfC�1�m����S�}��y�n�ށn�g ��7p�8�mF�L��&�bw9��'m���ڌE��̝c�}��2�qw���qkS�E$��n�g ���G qC@�%��՗�{�e�.�) �t	T�q�G9����������1�	��vQ ��*@8����z��_���܇ ۷����p�oz�y���%n8���G�O�:��`Z����ŀk׌�	(_�����6�-��  6n�2͕:���Ǌu�P�pJ9�,�.�DRNN8K6��1��ˈ��(Z�[�-\��t\�okM\�,]z�ɘ�5��$�gk�9z]>��^WwQ"y^�t!p��Z^�ӝ.	�E��WX��@�a�55���7WKn���������y�ukf����
H�s�q�g��KF���C����l�����lݽ۵Ue����÷�-acEGņ��h9b%:����Մ�s�":{M������
�3�,x�x���;����@��HP�$qg ��q��p��,���v�9�8ↁ#��97@r�Ү�Vw���W^����(h8� �tv�8��ͪ%5�)�Ȥ���-qR�&�8� �t�,�����b�8ݷ�ݼ��o)�-�����+�u&,��xa� *8Bp��<q;��m�k���5���w@"+9�u�1��#hǋ��zݼ��o)�6��p�oz����NLH���k׌��P��!DU��`�w�ݼ��蕸��}�>��\T�qɺ�*@8ↁ��c$�DD(��p0۶��m���v�n�g ��q��p��,���T�q�� rn��BJ�8�}\s��V�]s�HvKn��DtkVN�WC��5���{<<�u�h��-�R�4T�qɿ�@q�H}�TIA�1L�E$���o3�lrn�㊐8��w?ŘW�+�ʩ�J���k���5�ņ��(J$�irYK$���9���mh9�� ����y�u���a���?8��9��8�Nstw��c���3�o뷹�6��p_m�@۷��7=�݂NdRdBp�p�[Y�����@l�^�q�ܚv�n[��X�g~���9�1?���_D�3�m������8� ��mh9
-VY����x����9��qR���qg ��A��8A�D�zݼ� ��mi���� :s��9u�tL��f`_����) ��mh8�Ӝ�-�H�E�T� ~^{�zr���ڢJ �C"$�΁����k������7����9(���̄�U�T�t�%�����\!�$�G+�����Y%�;�-nו���wx>7���M�1��@?�?�@�ȩ ��mh�T�QL���o��z��7����ݼ�����Z�;�X�6w��G6�n*A_�9��>r*�ڒ�bO�Ⱦ���@���p^st�����ց�8Qj���������뼤Nst�����ց��r���F�6`��4R�e���ޞ���߷���&���I���Gj�Me�q�L�s���Hڀ��<��s=,h �/S��s�pK7Z���X#�β%r'�gF
���zCe��*�����z�+0!�f�7m��X�s�7�g�@Ӻ��c���}���:]Ym��f�.�����ȵѽ������wF�{-@u��/+˹2�6���e��xא�i7ks���=��pܗ�$��P�N�TW�Qub�&gOk΂��Y-�a�x���Z.���c�<�k(ugf�4�D�"s�����8��{�۷��=}��k�^}�1�x6��7�����)�[�X}�����Y� {�-Q%��cD���=�y�}�n��Rw9��N~%�0�^~�_�y���t��|�T���mh(���� #������%)
SW~�8� U~����qV�㊐�t�͵��Ϥq@P�'�F<�&G02G&�I���C�t�N�ju�2� ���A�v(�.��� 9�T�ߛH|�`ݒuM2j..��\��xz�g�QɖB<A����{�{���ʻ��:}������#�GQ���>�7@q�H	��ր㊐8�wq��'$X6';�6��p�m�t�y�����^*��G	�c�ۙ�'s�Z����S�*@O�M�$qR ��Z6�15a4���28�x��]vo.�L,�D���5m�������aW�3h8�>�7@��H	��s�{����"��8��{�׋ ��<z�d(J ~C��#x��''z�y����t�C�����C����8ō�I��2K���aD�MM����BĄ��B�@�N�aJ@2D-x ��� ?����0�2	%d!���h<�#B�V8G�x�"b�K,D��C�I1>HK!0T�JFI��A)#9��0� &�PA�����,�$(���1BH?��,�[�b1#Z#	(�Ѳ��(
���Z�j�h���D�_%	N.�������У��d�	1�	a�� d�I� ���)_�?���]�H9�N*���-8�'�������	�G��22 z �I=�?:UOª~���~p�_~���ʽ�]LӺ&�	EQ5Uk�'�}�<s�H	���$qR[���=�����z��*@_���7�#���yN�e����RdJ$`ҍ�R��9:����r���n�fk���F�sO��(�ng ۶��[���6��:�y�n��i��&D�z��`��<z�`��{�(�R7֪�qeҥuJf��`�}��׋ ����v�8�y��Px�2�]^/ ޼Xۺ�������J"/g��/ ���2�SV)���J���}���?W�ӤT��$��#qR�����X�u�%��=v���+n9�.�i���&�+Ob�u�cu.ix�8����T��$��#qR�stk�4��N,Hng ��{�>ϳ�{���x�x��DB����_tME�)]+&���s}� �w_���g ��{��2����8%M��n���7� ����1��,m3����$rI��9ށ}o3�w[~^�Xۺ��9(��7��v	��  X��ˮ���vt��e)\���W;7^KV�t�5��dP����.5� i�fpt�=fU��>`��^�T�:��n{g=�vLѐ��9����p�z���l>�ղ�'E٩"�$��չ�)���Cb�.ㆨ<,�ŋ��d��.��yAc�mWF9���i���]l�Hc��68�n�n��S�q��c��q�s���(�,������pm,<���)���hr�A1����	>�x�7�&�x��?�����͹�� ����e{	�b�����=׋�5������6�{�}QY�Nx�!�3�km��?�Ň�D(�2����7ذ{
e��F�0Nw�_[��m�Zn*A��I7@�p���e���]���R�&ց��I7@�2�����*�26H`&���y�]hrdݭ�s�^�pm��{��4��kC�1\�q��_��6��T�rI��@9m�t�ʎdcy��I73�m���(U~���9s��N���:ݼ�����d���_�/7@�2mͭ7 5�7�nٍ���7&&cI�pn��t�T��$�t� ;Ӯ��]{=��e���/1V�����$Z�@{wos�|��j
1̍��h:4ڤ0n���/��E������:���������7&t�������pn��t�y��kb��C@8ӝ��T�����#qR\�t��9�1��bd�&�pn��t�y��"I>�߼��X��'Z��i`au���ͭ7 5�7@�"��v�:�eG21��q%M���&�U:EH��@w���cGgW.:�����5���qdv���2�p��ҥ��aˊ8����Y]SM�S~�	�*@wtT�}�Rd�t�U�c!&<K"M����3�o����m�@�����*�mL���%�Zn*@l�n�:EH�Q�|��hlܙ�;m�����^��xr�u����"z
r����=p�[���9ށ|�,��!6ݯ �^,�����,��{�,�n�N�aκ���r�s�c�֌qg6��ܭ�z�y��E�ɇ���@wtT�}�RI&��T���V�O A�7;���g �ۺ� mR+��S�,�²̒�f�� �o���,9)��ŀ=����sA�6�s 9����p��X�ۋ��������UA��̬�z��w��m�H
���j��=�׋ ���z�ӻ�$�)MR�  2��m��)n��Q��)��-VK�,�H1l;/%�.�l=v4n��9*��[v߾���":r\��EYʹ��K&�ל�i%qm�v�mk����m��I�m�]�2�x읎�lb�W%�ܒ!�`Β�Z�"�yI���g��9m;�tpm�R�#��wfsX��.�d��mI��^�8ěk�� ��^ݟ{��{��ww�;n�0JHzd��؜':����g���u�c�ƹgВ���k���>�|;1�:�/��`�ϱ`����x��"�9�b�>����,qƁ�Crg �n�w�[���=o���Ȉߑ�n����%H����o^,�x���(�o^,���[S�i��4'�ng �"�|� 77@��HoǤ��&�B�W15~^�x�([��� ��g �o3�o�ѽ�r%�$���yV�WU��qs�hݢs�\��;��Ҁ�>)��d��������ݽ���p���IG�׋ ��ºʪ.�n���f��w�w�?* �%H�	DE�����q`�����v����I2bX�ng �o3�n�y�Ͼ7۷�ݼ�W�]T���'eڭG 77@��H�T���Q��ǃ�hlܙ�7۷�ݼ�v�g ���8wRq�Zi9��h
�-p���8��q7"���Af|;���,F�~ϱsg8ؤo�':�yH�T�o������=g��~���vG��ȩ �5H���-����B�9�8 ���s�[��*�߾�[���YQ[FL�c��"r"���� ��ذ�`Պ�V]%��U�~��x����f$��{������l��!��s�݊�̂�j�97@}P��Yc��m�!ЭVϚ�Wkg9��i��8u�:vӥ��%u�ւ���{-����5�'"� <b�j�97@��H��r�K$��T�*UVY�׋:!)���{�w>ŀo�z`�l�U5����EPQUv���x��Ò�/]� o^,ߑ��J�˹��E����)B]ϼ��ـn���-��iBQ�,����U3]uWvD�)Uk �x�|� $rn�#�������讌`b69����㠵�� �7c)s`.���gyz��V�p��R�j����߬8�#�t	T��UP�1 �7�dcy���pv��v�8�������Q'o&��.�������������R�j��T��ɺ�U@�,��jeT�U�
"�w��������K��X �����cJ��n�g ��v��^��~ܫ����`j�����U��'���@@�����b ��� <�UE3�y��
��֏����"*����g�/����������/?�����������������DEU_���/����������ʈ��
  ���G������������DUU�{�l������_?�y�������������@@�TaEI@��HT�	% 	�H@��!BQ"UDQ"B�1%�

TJh@��)F�(B$
@�P���`%		FI�%�XB �"A�BB��!	�$�I@a �!A�!dR�!�	@BY�T�adFE�P� D�d� VQ�$P��f�@��F!$!%	FF ��d$Q�!a�e�!Td@A�	F@$�D$AHF�RQ�IP�`HF�`��F�bA�Q�P �B� �aE B �`E	FA�	 Q�U%@ BA�TeAP$FA�	PV�P@�P	FAT�aD�D�e@�`BD�a!Q�P!!F��%$ B �	$a!TeY@�VP! B @!QH��@�H��@��I!@�$�	I@��	@��Q%@�%T!U�I@�	@%AYG?�l�O��Uc��;�����g������wAEU_���?ݘ�g��o��5���*���������nU�����������EU��O�(�������Q��33���kg��/���p��DUU�������"������#���������UW�~�UW��l�/����?�/����Q�x�*���?�S��9�����"������6"*�����g��������?�����)�����.ܬ�8( ���0�?�  ( @ ��  @     �8  @P
 �   �
    � �*J�� @�      !
AB�   �   �  �� �� ́CN��NO d�{�:���� �|��k��N���zM�Ԧ|���\κg�� �sGO��z����ukۃ�n�"j0 �}��S����ɡc�N�� |> �T� QR (f��б_�14���g@�8�AJ>� 3�(�&�c)���::l���� �)@�h�)c4 M6`ҍ"iJu(gJR�04֌Jh���N�iA�`Q��J14iM1�M 1)��1��� ��(�  P l  -۔���&���v����=���;�K��[�97r��} �<��Z�&� ڻ����ǻ�o� z;ܪ�tqk���u��=��x�p��l�k皼�W^�9�f����$  ")@�	��}�|�Sɮ���oyS�{�+�(���k�۞�zl�i�m�ܥ�P nRž�:y5�^�n�n,�� h�)b��N\{{�;]�͊_p>�������[�n����frݴ� �R�R 
% l ��t�ŝ�j���3ɪ^� 9�L��mŝ��绚�]��}�}��\�}��>s���Ͼ���4w��T �S���g���5��g���{�;��=ﶕ��ק��NMD��  =LҔ� �S�P��R�� �<z�R	(h#&��Ob�@��1 �O�BSmT�* �"B��� )�'�|�?��Y���������>��}������w��*
��DQT��*
���*��AU��(�}������\T�Ŋ��"e�@c ��@�*��`,a��,���q���kzח�FLF,
�(B�)�F� B��R#�5�"����e��p	�"�b0"Td��sc���;�o[��c(�@� B0�H!��_?�M��h�NK�<����bc��!4�i�#+)
��"��!�!��z�D���9�{�\Ѵ(��vF�L"F;ѷ�+��M.�>pӸf@�B+�BI!
f�IC �2O���riaH��+���{�x@��&�	��R4#\ "�$1"Pb`�E�������Db�B��bF��"��@�F�
0*��u����)�A�M�
�h�0���<�9&������P1����bM)Jэ����v!5%��>��5(Ys38Hs~z�9y���k��]� W�c�l1�Ǚ��C��!%H�!H,�� ���w	�H��"CWg�`��Wd�6��iRR䆝���,H�d"�!��ӳI
a��c	��ЍhbD`D�(#��5�<�#\<ܗVGć<,̙$J��
���Ek�vI�戆��VN<`��!��"@�I�]�)��1#�1�q]��ݰ
g�͚�5�|�m�/�xrs|�9��cS5������&l��\�CQU�>�����������}�;y�<�����[�Y7˶<�l�*F�q.�	���|W˿�|������)an�%���aH��$�x|�H/�$��`he d�
D#�n�	.@��
a/��.i!%0���󛚺��	xp�3[c	�$��������<�i�l͛��B�4j�I
0�,�$��X�Hā���)������q�/<�I�H ɭ� ���a��ay�]�,ӽ����i�8�{6�����٦5r%�)�˷���b���px����������"'��/��*C�O^z���8Lt��HX4�D��V!C�C`�H�޹�7�w��K�&�F��i�4F�
����0���5�6L4�	p	a35�l�F<1�y�\Ѻ��	s�sS<8�&����B�o�y�;�..�%ԨJ�èqZ���\������l���*K�}���(�����H���.����3��㽞����ZB!��c��p6�O��!L_`W\�ܸH����� �_WD Eb�
�F��F�8�O~��xhhԟ\)��~M�DCK�~xH�p4�) �-0���)O���0�<|U��1*A"C	��H(�B	S��p���`���*2��	a1މK�	�٥�eb ��k���l�\�\��������	L��14�;�N�2X�7��[��AHcR�h�ɪ��j�!#���41BD(c.a����L+����#�k�Cf�@�-+���^�4��BG�,P��QB�-e	�������5��4lax!�nc.��
P���['̑�ʒR����5�r��)��w&p�BB><�cH���!th�'�Hp�ч�<ِ�M�Z&:k¼H1JV������h��H�"�X\.��<�f�o�4�qx��Ƈ�$B0(@�!�@���l� �P�@B
FFPL@l404�xH��A��hv�V4�I��$.���@�q�l�&�d#d0	��8qi�h����Ȗ\,Xh��'��ѳ��m�!a�gB�A"\tl�#\4B��d+�A�B�&��B0�� e�c�J�����$q%�Q��Hm(��h@"c��|�!L��y��5#�Ўy�Ç����ha ���t1jm4����"���4	[�9��s�8m�"$#S �[���F�_�
�f@��lCŠ�R� -���d���2��`���P*$B!�����k�@A# 	p�D�X�4�XoR�		 0"F$"# R�$m��hf�[$X���H��7��@K��A�@�"Z�4y��y�.P��fP�;t����}3�H-��jx�i��5d��|�MBS�����@��.�{�5�4y8�SfԎ�CU��<
p��&hH!� A�T�SwD��YL h�$���$�HI!��$�H!R`l6Ǆ4�0$�ٹ����.E�T�DY$�R�R��sGC,�Jl���Je4�����Q�5v!X�5-f�!���ce���1�FɅ���ѶBIV	�� f�l�$�����٧�5|J�Xo�����n��=��	��:X�&��	!\ �LCK�R+ � ��+G���� D$H��FD"F��=0��k4z��ޘ�1 $b��(���b�v,�:f����+���*a*�( i�4H��x�\I��
�6a�׷43[���4�`V�h�"S$��x��)�����N	����9�P=i�G7w�r�f�)�>�2�F͸Os[�x��5�S���]k^x`�]��njGw.�$4`0rFx�$[Wԋ��c�:H��j{�y��C�d"���0Z���(�b���h���� ��
D�k B1 H�"l�Ґ�L��4�Y"y M�$�B:vy!BRb�	$�	�a$,Ń���	$$�m<)L���ۛ�C"xH�h@����j�$��!�d�	1B�6�@�.��4��������P�$XJ�R��j>	�!����@#n}�~E�a���O  ID�U�BP�	$�J�(y$
�2�����b�B�����'��4d�.p�oi���1SHх.�xy��{�����	E��q6@��Ўݧ���N1�������.	$���P@�@}@�|h�,��%���9�i6L���1�H�����$#�oɐ�H�H1�`f� �/$�&�r8��Y`�	D��4i�!��pF�0����12L#%�oi$�acѺnJ9��]����kz�1� �����
@�JT�ũ�l}P� � � �s�t�S BM9ɝ3�9+���5R�ժ~�����-"�1�D F���!a����=���  -�p             m       h                                  $ 	                            �o��m�� $�	۰�lBA�kn��mm�kX 6ȣ'H�m�p��m� ���G`m�����9���ݔ��-��  6�@  ##nۣ�l�UŭjM�����j�� L[�U��m��:�d���� hh	v�j�6Zn��N�oP %�v� m��[@ �$  �5k�����ami;p�� rM�b������  	�-��K�p-��lդ�h	kY% ��6�iJ��f����R�j��lm��m�V��j��m� ��i��KVMa0  F��kF�z����Y�
U+JQ���v��E۷i0�$  �Y/0�a�����o�$�h������[hhm������ m��m�ӗ�� 6����Am� 8Hp �S]�!�'+m�m�*�
����2�ʫ�@VͶh ky�2qÃR�^��N�gZ]j�].�4P,�Y&��7[��m Tٸ	 5��a6�R��w-6JB-�hٶHr�m�]ʸ�f�	 6��6���h ��6�I&� � �I�[AhmU�흚�)�U�A����mB(SU�ʪ�$r�v]6���T���7h:��d�mC�y���s"YP�u��I�E[�˻gE6�  5�m pmٶz�h�m �`� [�I��h� �Q��  sZ�����  m� H$�j   �n�� �m��i5�΀H6ض�H�Бm6ۀ B� ��p���q �	Gl��� [%s��m�A �n���[p� �`Yv�����$��X�H[d t�� �i�lq���f� ����D��j$�l ��kp�^H�-�@�nݭ��[M���»u�\�I�  8��m�`���ڑ��[)�*�UUWU!<��� � 8�vYv�������I�� [R��ݻd��m� 2�� E���ɦ[���$�-�6��� ���y�� �p%�i��ȓm� HM�K�� [A�h  N�JHR���kx��U�P�W�   ��� mU�� HzY�-�Ǥ�@  "@+�����m�ц�H�H�`[@l�	       6�zX� H  ����i6� �6� 崃 �	;e�Y�l m   [M�a����A�       ��    m��q�A˾�i������@�� m�(��	        [@  [�����rBG�]7.�8 H� 6�D�� I'�k��[.     �2n�        ����+� �  &����}�   m���ݼ�@���$+n��� �IAmf��`��/Zmp  ���H�$�   ��l�([}�P �̓��"�+�@$���s;���  l$ ���ϟ    ��L�lڶX@  ��q' m���I�����s0@�UPc����UJD�3���&��:Q�lm� dPCZ�)k�iv'�tUJ��`l6�a�J��$��l� l���q�>��� �J�����@k�kh.JΠ-�D�i�ɴ�m̒-�l��M�nq"D�D��fꭁ&�q�kX �oZm�k���M��m($-���M�[v�6   p�j ���E�i��*h.���(������   �؎�ă�-͎&�[N|�}:6���M��i�Z�ye#6܅-[uW��:4͊�P��+hR%��@j��j�v��Vą���ג)�M�6U�j�ೝ���9%i$�ȶ�� 隻f՛` +j��㵷p�UK;�	en�ZU��s�HeRmm�( 6�Z�� Y�*	�i��EJ�R@ ��li6m� PZ�l�UT�X��W�iS5�X5;g�&�۶ �6����l 6��[@��� WUPH��V�)�V������N�k��lm�v�mn  i˶���gΝ�[��h[@ &��  Ҷ��v�h��y6X`   =��p  k5�# Ԛ�n� h�Y�p�� 6� m�mvkm�� � m� ��4u�e�m[`��hm�  ��m���,e��(U�6�` �`����e��.�Mm�  �h 6��@ � ä�����mĄ�m p6�� l�6� 	  ��E64YmX5@�����U�B�Z���F�kkp �$$m�!m��  �`H	 [@ ��I��we�����[�6� 5��Zl �`p3$a��T��VB2�<!R���He�^��A�V��t�T�^������x�VZ���&k̔v��M@(m���������5+�Y�C��V���EW ���:>|�����^Z4�� �ÁŴ-�$m�ܲ�$��m�I���yͩe����"�-��j�mp	��wρ5Px�������N֭Z��  -� n��u�  6�� H	mq: �Ӧ�f��4�9�vKYM�m�h �l    ��ݰ[@$�8 m��	��&մ����$T�lnM�;u��  ����m�[@  � $ �}           p�J�P�ȶ��8[@  ��-�m���[A"NpIm-������m�M�62󙴀  ��-��f�@�l.��$h"�� 8  @  p @     6�gY� ���6�	m!� ��    m�`    p���A$�l�\Y(�Y�         ݵ�`p�9��[[-*�U[ T����T텶�8[R � m���I� "���-����    8�   ll[Kh�M�;-u��m6�����%�i� k[�r�lm� ��%p�` �^�m�-�� ��l��   v� 6�  � <`   v�m���J[D���ꀎ8�(��v�l5S���        9��d��8u�մmH�M�	e��:H=m �j@[@d�$턲J  t�Ym���o�����%K^��� ��a �'[hR�q�ul9$�m��e�[��٭`   ��� �|����UaWev�UJ���*�˳��vYH���j�̐�((
������5\9evMW*�]m�$�:v  A h� m&m�&�5�lu�  p$e�頄q�C�jP��n�P��mF�N��l�g`fR	���!2V$݋���Z�� śҁ����55t�_R�Rӕ�%�m�;,�.�Aq.��N62se�첚@U@���T��4;��+�m�U*��5WS��Ӣ��6݀��0��6�� ���� �EkŻa��\��� �X` #!�ͪU���2�\�����Ȫ�u�6�6�Ԁ;m� 
���d�lҳks`8d���  @��[@ $	��e:t�� Wl�UP6�n�sm�  m�   ���h�J�� X"�� A��i��h	 �Ѷ�HnZ-��ȶ�h H ���[hK(  $� j� p� 6�m�� ��a�m�$ -;e�� n�ۀ �G�|   (I�� m�0   �lq��@ �[N �l�   �[\H6�\�PHm���8m���m��6�   N���[� m�� �-$��JH!Sj�,0��`  �5Wg[m���h6͛` S^�Ӥ�ۀ  �ٮ�koc�� �Zl�4�<ɶ�� �`m�������� ����]��ޠ	�mɲ�h�m�  �۩����6;v�R�OS[p�	VBi^iV��Vy_���� -��m:`]68 ?������w��w��w���J� �=Q

�P���^�/���N��X!�s�C�؁DѥE""����%-jPߨ���4"�F@
�Q�������`�'��J�iG�"�“A�@@H���� �hz�ꨔ~F�π�Px�S���%���A�
�Dp"�@Ҫx(����	  DH"D���+�b�EĪʊ�UO�>� L�1_`�a�kM���@� �<t>z�ɨ!��Q�E҅pX�	�'�(fǈ� m�0�"@A"EQ �X�1X!��p�P�G�z({ "@D�!��<U�(&�FPM�_P@�]'��+��!��`����*��"�B
�`
|��@����	_�7��*
��x� A_@H��	��~Ͷ               oU�h�(@�q�M,��6��W3sؠ�iugg���bO5΂���G+�6�#l�z��h`���a��ec^#;��v4���h�68I���#�h];g��f'�N�Ͷ�Zm���]Nα����D�]�{(�����z��\��vEt�m/+��*�Z��hԁU*�S!��q�2智��n6��C.=��)��T����&Y{`+���ز��KZ��ɵ�1h��)���f��.^����=��Bj(�;e*���P&��۲��vZ���W�8�3����{n��a&հ{��U�T9��U@U���ld�r@-k�� .�6�m��bw�Kk�ʽu�4.8z;$��T��2.��7l�H+ym;��Ep�l:ET���ڏ\F�Y073���@�k\�m���1���UZִ��#�}�m�m�X�"skS�9��r+��X[��h��.8�-x��� 
�{v�n��mu��K�l��.0���j�S�j�()�*�!@cR��vu'�+n�۱��mv
U������ڠ�8l`,5<��YP����UW�u��xݧ�Pm&+P�n�nZM��|n�ImlnSXr�ۙj��24����.�T��\�FBY涚@ ������@���ɰ,�I�-�Um��$�XѣSa���K�e�SKj�7Y'*dZ��)A��v��6�6�j�cr`���Ҭ�Nv�4��;�M� ���.�p6��)ʎ84��p��a a	L�T�S�n۳�-���P�������e^�s�^��t1&���<P�1��s[6�@�ܪ�A7�ohS���5[5m@�v�t 
��-jvV5D"@X�P�a���mpW<��V�6*���O9��j�t[��*��ջI2�3ʬ�2/m������n	X! �=b�0ݪ�m��f�jkZ�k-�iA��
� !��. i|U�
@<;�~]�q m��VuI�tZ��˖�|�E�h�aT��5��0F��ZA�Mgu�3�E�6��˴(�]�)��.�m�5�n��{Zl�ܝ]��}�m�Y6�#����m�T�U�tst��rǥ�t�N�۬�.5ʩ7c<<�OV�w`��E����@N��}�Iq�{l��
n7Cʸ�㮰lvy';c����ܺ��I��PAҍ0Յ��f`���y7+Ϝw����nǌ��d�]��ȇ�<|�Y��v`��`}����	*I|�{7��-aB	�ܘ�S�z��o�J���Rߌ����>}ݘڻ�܂�I�d����Δ�>Vנ|�נw>�@�U+Q���`��^h���1�rb�r�?�n��ו�6�I)2F��=�ֽ��Z�:S@�[^�����1�n)�Ɏ"♒z:^��bM�"�ݍ��em��n�,C��s1�#��D�0��)����ݝ)�|��@�u�@�wx��iֲܺ�]�<��_M�	��|�)X���i<^Y����*�W�w>�@/eT�xA�K����ֽ��Z�:S@�+�"q(dC��.��Ϫ�=�Қ����a�nLJ)�n=��Zq�)�|��@�u�@��7q☚y0h�P��X$��kq�ul���� v�.�X{�W,q��[�7B�I�d����Δ�>Vנ|�נw>�@�U+Q�	�$��N\��& �-Ξ�o�^�Gs��'z��zs�5�V]#��ּ��S@�mz�j$qD�0��)��9ht�\��& :d���19�m���@�gJh+k�>}ݘ{;� �U*]^����Э7���Κ����m�r����V.���l�>]��k9�n�-[�����������~`�u�@�}V��Δ�;�WVLN%L�cR=�ֽ��Z�:S@�[^��ì ��
9�n=���:{�I�[��ኴ��H%�$m8�vt����ֽ����P]��TU4��C���V�{�ƒx`��'�d��Ɉ��@s� 9�ܙ�{��۫`�K75���ۜ(c�o8ە�۱�0���Tv�MwZZ���ul�3?6>}ݘ{;� �Ww�RUU�?{� -��8�"c�Lx��@�}V��λ�����Z�WqQǋ��6�QŠ{�����ֽ��Zz���s"hH��h+k�>]k�;�U�{���m��Y18��j�dws ��v`���v���;�}�rN_��7$�#� z,��I'�;���ӻ�~����@�����ϝ�����8��dӷ^k%���1��u0.�F��r\��������rv���7<�۩���{\9wj�8����*Z�Y�G���P^P����s!����!W����Ʈɶ�c���%u�h�	q���d;j87�R��YP�Y���=Cwe�]��-�'3Xo[���Aͩo)�vy��|��R���=j@����z9��qenE�^�o$N^G=�@��g��u�{q�.6�f���������@s� :䘀��1軤�c�wv6�]���]�Y����8��L�}�w�u����7$��Rf��mz����j�;���z��9�,�i8��>V�@7�Z�qR�I��,�ͳLs	�q��ՠwgJhVנ|�v`���O��vK$��Zr�Z�x�:��Wh�/�6�n��^8���(�&�n��x�	̃m5$_nY��<��@�[^���� ���8��M	���wf}UT�T��UI"�sr`��h�Қ�cud��R)�d{�\���@7O`���1 �#�d-ːw-��$�S����埍�z��mz�u6R(�6�]���]�0*�Oo��q�0��Y�u� ư�Ly1Ĉ���/m���
{.��.ױ�N�'�9�ݏ7mm%$�x��Dk���^���^��}V��Δ��Y#�HŒ�'$z�ɋ��Wds~T߄�9��#�b&9�ǉH��Jh��M4����z*	�wn��nI���rN|�*8�b�m��4vt���^���^��}V�^���8��M
ʽ��b����@s��F߇���h��m��ɯDH�����vJ��A�W�=nR8T�xcv���.X�̍F�i���[���Ξ�뎽���N$�b�a�@�t����շ� ���`=ݙ䪕&��o���9�d�n�g�@�^�@�u�@�t��ު�#	�F�K0<�|��L�}�w��0˨I*T�ݤ�K���� s��r\��5v��7w�& =��6\s����z;$'b�@S���z���]�����3��^��n�8k��1���Nڽ����@>{6l�� =}k�>�⣏1��&�JC@�q(���1��1 ��p�n��v�DА���^����@��S@�q)�Z��Y�NI#pMǠ|�& ;��͛���<��ܻq&�J9�n=��M�Ħ����@�zנ����I$�I$�8��7gQ&�ufuWe�ݲ#]*f��3u��˥rN�%,Юˮid�����'���n��Y"�%�Y-�v'\\!�F�Y!y��;b�$[��m�m�m;��j; a4\�S���%_5���.���ɨOj��ۅ����A�+���і	���<��5��kk&u�vr[+�p[s����W�ָ�鼎����h8�YP8K7���,�����]{7�/|���lE�7$�����f,�ݽv�]d�V�b9�c�n��O�|�k�>^�����W\M<�(�!�@�������c���͂ �sv8�Y2c�&�z�ֽ�>�O������wK�q�}0��eܶA�[�e�� =��9�`�����@�}��<�̉6ڎ-�Ħ��c�g��}�v9h�����E�[s��lRi����=�n�<
�G�{Q�kp���$��BCJB&�I��^����@�Ϫ�=�Jh�6R!����r�ws ��vfU*J�*������%4�����둤Ț�Q�33q��-͛������\��ABG1,y#iŠ{���>^����z�}V��^��|�i��1X2�NY�6�^߉���$�*K����o�o���|��i�ͷ䪒�ﾟ]��؜B���b��͖������3�[	��[ v��ݻ/^ �!EQL�:�d���K�����$��V�$��;i��%�ҏRI.�Q#�(19�����Iy��g�*�7�nx������1��ӻ��mWة#����m��z�K���}�V�}��7o�ʏ� wLP�!A�R$A�أ,ޗ��!�Pp`+�����0Ü�8C���Ѕ��J<B"�mY),��B#M���p��a�!�$HH`�	$� �E�$�6څ$�!!�BBB�d"B$X��$`�HIBB���ň1A�n�z�H�@�$�´��XJ���2 �%T0�RD�A�$�$(#�H`d4.�5����Y �"�c$	Q�Q޷����NÊ1_�N�*�����C{"z��8 ��F��Z�g����|�-������fF����v)mݖ�lc����ʩٹ�cm�M��������1��I7M���g����왑�&�Y� }?�����7�;�cm���������zLm��UO/?��@����������q��p���u����.wv����qk�t� ܱvV?y$����I%�u�>�$��Q�I/�Z��$���
8��#m8ޤ��;�/��*UJH���Lm�ɾ��������6ҽ�~_A�	�����%���Ԓ_>���Iy���I.����$zݑ����@q�ۃԒ_>���Iy��ٛ���߸o�ݰX�ߟ}ZԒK��u�B	̌x���K��ORIw�u�>�$��V�$�Ϲn���~����54��BL�kk�sn����4n0lr�o
C�,�p��/n&S��7J�Q��$�����%�ҵ�$�}k����II:���m�／b��ݷ#~���%��o�o����R�ro�>���&�gP9�m���xs��s���3�����r�wd��|��O��)#��1���_֗���I.V~���V�/�9q��7�$������$����}����V~���?�I.��a	BǑ��ɍ�)7M��6�^߉��M���6�fߣ��|�I%����~�݅����ɰ�˚�E��:i�4�q��nhrq,n�m][���G��f��"�"�eV�ծ��]��|�v"x(��h�g�hJ�C&�v0욶xF�nU�+����ظjj�c��0����t�9{����j����uvõ(gA�u=��г(��!����y=�	�s"�͠I%�u��y:�58^d2���F� ��Y&�{����~Wϧ�*7C�������"ֱ�������w���_�$��'.��Z�8��F�W}}����������|��Os��ٷ��������l��%f[2
���ʇ�����} ~;~���{����;)ٹ�cm���2��1�ǉH���cms��Z�J��R�r6���Lm��Rr�ޟ|�o�S�#����m%#[���������$�+?RI|����%�ҵ�$�[�$1Ĥ�6��!��%�ҏRI|����%�ҵ�$���}�Iq��kŋ$�-v��=\�Sn׉�,Íg�cy�\�<������Η<��Λ5g���~��_@>N�Ǎ��ӹ��*�r6���Lm��}��A�a"�,�} }���|�{���"�0�@�,JEuuo�O���6�߉�����>��e$����KPP��,ymƵ$�Ի�����G�$�v���%�ҵ�!^�cLM��D����%�ҵ�$�v���%�ҏRI{��}�I/[�7i�$�q�K�m|�^}+Z�K�����%��������֮xX��c����OkKۜ���D;���ݸ����\�im����{b�GPƤ(�����ZԒ]ݵ��I/.�z�K��|�J��I����i)Ԓ]ӫ|�^](�$�����$��V�$���RCJH�i%r�������1��&�g�6��T��4x���w�o=��wm�ϵ�ٜ������#3��Y��{���.���%�ҵ�$��V��$��Q�I/�a�#Iē���8��$��V�$���v�o�I.V~���_�$�;�5��v�Z��srom��\�ny��΍��,� Zt�걝LX�1�zUdԒ]ӫ|�^](�$�����$��V�$��"��4��A?�m8��$��J=��3iyݯ�KϥkRIwN���I��(�F9�Q�=I%�z��I/>��I%�:���%�ҏRI/��$qEjA��|�^}+Z�K�uo�o����ߒIeTVw=��|�o���s��-ʮ
O������_@���{�O�m�ov}�m�v�<m��ؙ��$ݭ���c:iQ8�����v<J���s�.p�.�N�r�kV���/ߒK����$��W��%�ҵ�$��V��$�y^:�N4㌎H=I%�z��I/>��I%�:���%�ҏRI}��N$�mG0����%�ҵ�$��V��?�m�t�Ԓ^w����
�P�ı<���Z�K�uo�K˥���_�$��J֤���T�Ƙ���țN7��%�ҏRIyޯ�Kϥk@����~��>����V�UPU�خ�Ά�&^�<�I������8d.��k��[�[���H�^�c�l���m��y]�t�۵.*�5뢺�� ��]��L���d��)��X��۶�9ݰnr<��7��! U;�Ź%�G����byx����z�pƃ4�.p���.:^��l��6����V�!�q�F����������i�i�_��{�󗯌���Ah�L���[��ۜ(aړ��]��N�h ع.b�95�iX�Q��aCn�$�����$��V���{}�?*UI�W9m���m���e�PƦF�q��Iy��jI.�տ�I/.�z�K��|�J��I�9��ƤkRIwN���Iyt�Ԓ^w�����ZԒK��I��I(�|�^](�$�����$��V�%�o����U�lN	���<�\@z��@6�e�=�`����+7ƺ9�gJQ]2�����s���-{2�obK��Z�c�t��2�q��}���hs� :㘀郹���ܶԅ�$��w���9_�-W�I:��� 7g�@���|���"�EOq�k�#"m�ց��S@�^���W�wt�h��TQG��I�"p�8��0�;� �{{��J��4���H�5�dQ�=��@��Z�>�JhW��>�qD\PpX����h�x����vk�)�s��a�qy�1ZSE�w�|[��������������2��@u�1��1 t�Ct��K�����x���I&οo������+Z]�㭤��Q����<�{�nI��f�O@@����k@��)�}��L�q������1 �ٖ��=��9��5a	K"m���t���z���@��s�вb�6��p[uΗ����,򻷁tl��b]���3�aPӘ�'�#"m�ց��S@�^���W�wt�h��TQG��8���q�YWg����-�{�[�EQ�S"��G���W�wt�h{�4+�����0K�&����+Z��M��z�g���I��@=n��ppi��R5�{����1��1 �ٖ�9���@p�cn�k������m�S��N�����8��m���Z^e'M���8��0�;� �{{����s�~4W����ȇD��q�/u{�?�Sf�ߣ�9ݿ�f�S��c�G�țn=��k@��)����K����]=��S�i��16�v��=��9�_9�>�_����h�ߞ���p!ۆ��z�����;��ǀ}�ޘ��!%hM**�"��#r���Dhı� $U��H�=+n
kj @�+�b�mIjI#,c)-�,��!�4�R�fr @D"��.BBC¦#ZT�C0��%�HD>C1�� ��!��a�HE�͂ŉ��FH:0c���1Hb&��H1P��c�j�& Z�$$A*���(,4<H D�B!0�B,RA# '3Sh0�#���`D"�q	 ��L@�	�4�p`d�B$�	 x�]h���0B�B);��;�>m�ְ  ���     #m�    v�芼�mm�ӝL�r�E�MVm���@Y���<�:&�[�(1=���v�t��:�+n�^�e��&��#oOW�/=�X��V��k���,�؇k���lZk�ִ���.��Qwh6�큕�@�c`��-
s+�{uI>8��Gl�eyykj��( �����h��+��b�5jB��<��,����=��}�#t�Vk�k����,�!��/n��l&Hy0?����H�Z6��X��M���]�����YI�Uኪ]ɶ���*�n1�B�Tю.�V��r�V�KU��9,�d�M�`�Y-�b��5��� ��' ^�OP]V�2�L%�u��F0sl�F�AՊj���UVʲ�aĭۢ�2c�-v��ckX�
1��z���a[���e�n.���c��6j�ƺ6+��+T�d4��ǟ�`��D۳�wu�h�ĝ�Ɲ�Y�Jհg9����r�YB^�۬��-�@���dBN����5)��@n�e�YUiK�b�q==%��ے6s=���yUU@��ٳ)���2�I��ʀ�&R��!����;WXwG\�7�Ijht��l^ic;f���f\�"��6��ZT�76�<�f�H����PՃ��+v趘��� %dlI�m4���.��F����*�UQ9-��ʷ5lt�մ �9l��w۬�O���dµP�R^+"��շ
�Q�㵳;��eUZ�3��A��UUkRxÉN֍*.����wa�>7��@U��{�m��q�U�ID �UH��˶���ظ�-!��y�+궗��gUs��ځ�j�@�J#Z���tA�P�ٲ�u�5Y�&��v�9˵U$�]�[�:lO:�Ŧ�6C:#��z�`�a�f�ʮՓZmv�FX=�nx)U�kl[��W�J�n�@/D�뛲�g�r����tR���ԩ���kYn[4hz��wC�T� q3���@�����N�{���~��� m��5�]��b{T��G��#1�:qk��rݷ��y5��@6z+̴7�|�����u��E�CZ��"P�d�5ޔZ�el�M��;t�<[3ۮy�&�0dH����Ë�3n%�R2�m��bِ�mԜ�F�D��`�9{d�/�f�ɲ��Ycb]�c�Z�#0F�]^s��v��Z��-h��U·<Q5W;�����V�~���%T��&@��@��;-IbJ�����wk�^�cQ��	ɺ�	ywlsLje�E1b�=��ߞ��ҵ�}��<�W��*H�Ēs#m�H��̵���3s~�b��b �p��2'�i%#Z��M��z~���K˯�[g�
�+�m��Q�����z��^��ҵ�}��>煤i2!���q�/uhcٖ��=��9��y2��vs;K�G�������wa������s��S��v۞�X-�Zé��l�?6ߟ�fZ���� =|�#��?U����?\�<�F�Y>{�����{������m9�a! ��!?E(�P4ț�b}���6��bX�'s�{�ND�,K��r�9�&TȖ'�~����]R㚓SVff�ӑ,K��?w�m9ı,O3߻�ND��"}��ܻND�,��\�猥�I��I��7|;�nݐz5tR�5�ND�,K����ӑ,K���ܻND�,K�~�fӑ,K�,ȟk�fӑ,KĿ�t����-�4k32eֳiȖ%�b}���]�"X�%��o�iȖ%�b{�����Kı<�~�m9ı,K��wZ�k��x;y�ؤ�����gqͽ8r=Gy�;v�n��kV��s��yp�<r%�bX�{��6��bX�'�߻�ND�,K�������}���%��w?G��)2�)2����#���nB噭jm9ı,Os�w6��bX�'���ͧ"X�%���o�v��bX�';��)|R�Q҅&R�?~�c��[��K��ͧ"X�%��}�ٴ�Kı>���.ӑ,j@��)�(�q>���6��bX�'s���Ӓ�)2�)w���X�w,N)e�w��(�,,O��}˴�Kı<���m9ı,Os��6��bX؞{��XRAT��3�b%܊�nչ�bI�9�i7�}#�g�fӱ,K��߻ͧ"X�%������r%�g������Q��\�C��l\Xn������\&�n��d0��"%$"[��ꑢ�5&������Kı<ϻ��r%�bX�{�y��Kı=��}�ND�&Re.ws�R���L��Ow|;�nަK�WE-ֳiȖ%�by���ӑ,K�����m9ı,O=�}�ND�,K���ͧ"X�%�{ߋ٭an�f�d��m9ı,O~>�fӑ,K��߷ٴ�K�dL��k�ͧ"X�%��w�ND�,K�ޓ�Z�億m�ve/�L��L���x�_D�,K���ͧ"X�%��w�ND�,@E����}�ͧ"R�)2���Dz�	d�!wj]ٔ�)X�%��}��ӑ,K��=����Kı=��}�ND�,K�~�fӑ�{��7�������;$h��]v��)�^uÎ=!�m;�����[oM�{6�h���-��r\�_�I��K���r%�bX��}�ͧ"X�%��o�a�O"dK��5��ӑ,K���בּ��Xȥ�K���)2�)2�u}�ͧ!�@�DȖ'�w�ӑ,K��;��m9ı,O3��6��bX�'}흹�f��h�tj���ND�,K�~�fӑ,K��>�siȖ%�by����r%�bX��k�ݧ"X���]���,NT��dr̥�I��K���ͧ"X�%��{��ӑ,K���_v�9ı,O}�}�ND�L��Ow|;�nݐv��&��R��ı,O3��6��bX�#���v��bX�'���ͧ"X�%��}��ӑ,K��P"�O�_?À +�\�u[ymݫ���{?7J�T�,��:GF�V;;���b�i#V3�Q�bwE������e,�S�5�)�6�:��6�$�F.�R�9�jsT��s��[���f솹;p�%r�x��k�b+��mV�'0 ��ҁlB1J�ƭ�i�:�Z�,�I��P9c��z-�W�ݔ;cp���\�'d9]�{�7f�3� �xy���q����+h�.��^�㌮Ƹ���ۈmAŜu�M�wn��<Z��u"�g���,K����M�"X�%��o�iȖ%�by�w���Kı<�{��/�L��L���G��Bܰ����ͧ"X�%��o�i�D�DȖ'�k��ӑ,K��>��6��bX��ίg���I��I��:�<;c%���Zњ֦ӑ,K���}۴�Kı<�{��r%��ș��fӑI��K���)2�)2�퇽n�&��\�us5�]�"X�%��{��ӑ,K��ӻ��r%�bX����6��bX�'���ݧ"X�%��u>�K�c"�I.�R���L��\��x�_D�,K�~�fӑ,K���}۴�Kı<�{��r%�bX���ɝ+[t���tA��=�O:���"s�vM�w��!�zێw[Ksဎ���ݚ^��yu8�D�,K﻿�iȖ%�b{���r%�bX�g��l=Y�L�bX����)2�)2�;������4e�M�"X�%����i�x �Z�&�X��{��r%�bX�zw}�ND�,K�~�fӑ?���L�b����wnݻ �a���&Re&'���ٴ�Kı<���6��bX�'���ͧ"X�%��}��ӑ,KĽ���[tkYs&\�m9ı,O~>�fӑ,K��߷ٴ�Kı<ϻ��r%�`~��}��m9ı,K�߉�kPɫ��ɖ��SiȖ%�b{����r%�bX~E>뿿f�Ȗ%�b{�w�m9ı,O~>�f�|Re&Re.�+b���Waah$�=<���]��;�hۋ,��9U��n_]���:ylF��sV�����{��7�����m9ı,O3߻�ND�,Kߏ�ٴ�Kı<���m9ı,O�����aљU�Y�����{��7�����Ӑ��$r&D�>����ND�,K߻��iȖ%�by�w���K��K��}d.匊�I%̥�I��Kߏ�ٴ�Kı<���m9Ǌ#�"�Q5��}ͧ"X�%���ze/�L��L���<�Ȓ�V��V��M�"X�%��o�iȖ%�by�w���Kı<�~�m9İ? �2'�;��iȖ%�b}�e�l�0ɚ�Z�.jm9ı,O3��6��bX�'���ͧ"X�%������r)��I����K�)2�)wV����e��ɃZ�$��������w#�GnLY�t��DX�%ܝ�Ԫ��t:uf��"X�%��{�siȖ%�b}���6��bX�'���ͧ"X�%��w��ӑ,KĽ���[tkYs&]k6��bX�'ޟo�iȖ%�by����r%�bX�g~�m9ı,O3��6��bX�%�'f���h̙m.�6��bX�'���ͧ"X�%��w��ӑ,K��=�siȖ%�b}��x�_�I��Kӫ�ö',v�Wv�����K�Ȁ2'���ٴ�Kı=Ͽ~ͧ"X�%������r%�`x*����;���6��bX������k��Y�S������ŉ�{��ӑ,K�����m9ı,O}�}�ND�,K���ͧ"X�Re/�%U����dv�9b!mGe��2����v�ԮC;�q�ϛs1�6�a���]m�Vp�r�Ev��s�\)2�)2��{?K�,K��߷ٴ�Kı<����r%�bX�g��m9ı,N��d�f�.�V��w"�̥�I��I����K�,K��;�siȖ%�by�����Kı>��}�ND�,K�~��j�!���2��&Re&R���br%�bX�g��m9ı,O�>�fӑ,K��߷ٴ�Kı/�w�����jݰww2��&Re&R�｛ND�,K�O�ٴ�Kı=���m9ı,O3�w6��bX�%�~���a�����2�iȖ%�b}���6��bX�'���ͧ"X�%��{��ӑ,K��=�siȖ%�bqw�߯�����$ m����W	��Z�ߕ�|��أX��	f،�KՌ�b������<P�Ӎ��K��E[����ӖZ���ݸX{m����7�����CO�m6!:�^�n��-�� �E]`t���:5�BVE�����D�F�ܹ���ަ�`�������pJ�.��bVS`a��uϝ���cc0cc��g��;q��.4�����盍�o�$�Fz���8���bq@v�B���Yp���W`�;g.��s���]ju9ı,O>���iȖ%�by�����Kı<�{��r%�bX��nx�_�I��Kӫ�ö',v�Z֌ֵ6��bX�'��{�ND�,K���ͧ"X�%�����r%�b2�{��)|Re&Re-���8[%�3Y��f�iȖ%�by�����Kı=��}�ND�,K�~�fӑ,K)2�'}锾)2�)2�}f��8]ݧ0֌�ֳiȖ%�b{���6��bX�'���ͧ"X�%��{��ӑ,K��=�siȖ%�bw;�N�h���4[�Z�356��bX�'���ͧ"X�%��{��ӑ,K��=�siȖ%�b{���6��bX�'�;���٭SO6�Q���Mun��np��z��܏klFtX���u�ml�����N�m������Kı=Ͽ~ͧ"X�%��{��ӑ,K�����m9ı,O}�}�W�&Re&R{��.�vAڷl����bX�'��{�NCJ'�� � ?�]wı>����ND�,K߻��iȖ%�by�����JRe&R~���.!A�V㌎\�_�K�����m9ı,O}�}�ND�,K���ͧ"X�%��{��ӑL��L���#�ءn+R��ٔ�ı,O}�}�ND�,K���ͧ"X�%��{�siȖ%�b{���6�)2�)2���Oإ�-���K�2�"X�%��{��ӑ,K��=�siȖ%�b{���6��bX�'���ͫ�)2�)l�OY.r妥B\�͡�^۲qF/ �rCͮz�T^�j6cq�.6��k/BiI�3�������ow�����9ı,O}>�fӑ,K��߷ٰ�<��,K�����r%�bX��g�Y��ȮԒ�e/�L��L��O�ٴ�Kı=���m9ı,O3��6��bX�'���ͧ"X�%����;��殰�n�k0���r%�bX�{��6��bX�'��{�ND��z"b�>$|!X��2F.݊	{�h �< ����b< �"�e!BD!)!a	�)�IiB�)'�2>#P4� Ȱ�(`,�Č ���GX`�a������Q"U�� 	 �ĊU��WZA��a��!�*&��-Q�/�{�A=POD�V�ѣg�)ӱ2&��{�ND�,Kߏ�ٴ�Kı=�|O��$h���dr̥�I��I�������Kı<�~�m9ı,O}>�fӑ,K��߷ٴ�Kı������Y��pT��}oq���Ǚ��ͧ"X�%������r%�bX�{��6��bX�'��{�ND�,K)q{��<�)m9\Q��-�Xӣ���v�7g����x�9�Ynp\]�ۜj�eֳiȖ%�b{���6��bX�'���ͧ"X�%��w��ӑ,K��=����Kı/��;5�f��F�L����r%�bX�{��6��bX�'�߻�ND�,K����ӑ,FRe-���)2�)2���O�.�][�Zњ֦ӑ,K��;�siȖ%�by����r%�bX�z}�ͧ"R�)2�;��)|Re&Re-���H�r�\�����m9ı,O3߻�ND�,K�O�ٴ�Kı<���m9İ>D�����6��bX�'������Uq��U����7���{�}�w�iȖ%�by����r%�bX�g{��r%�bX�g�w6��bX�'�ߟ��kax:��N��/m���Wv�F�2m�&��[���%ƱS��bz�s3WiȖ%�by����r%�bX�g{��r%�bX�g�w6��bX�'��<��&Re&R�w���mƤR��̹���Kı<�����Kı<�~�m9ı,O>�y۴�KĲ�;��)|Re&Re'��.�vA�5�]kY��Kı<�~�m9ı,O>�y۴�Kı<���m9ıK����_�I��I�ڟ��ڻ0�.��ND�,�02'{�g��Kı=���6��bX�'�߻�ND�,K����ӑ,Kľ���֡���a.�WiȖ%�by����r%�bX~�����O"X�%��}�ٴ�Kı=���nӑ,K��߷��@���S���vɥ-�\6�Ϯp��<u�:�:�G!�;lNɗMqm;��=n�;7lu�Om�>۳۵v�9K�V�q�����ˣX��N"LN����ؗ6�eE���h.}��,��nz��Bص�ZТ;��]7*�Jm�8i^MV�`){��n㑃n5�'Wesu�s�d�
\7�tµn4sѦ�eH�oS�L�_���;����D��m�ͷk�8��'m� �<�q��lͼ������)&�<�#4�U�jz�D�,K��߳iȖ%�by����r%�bX�}��iȖ%�by���)|Re&Re.�}d$��.7r���m9ı,O3߻�ND�,K��w6��bX�'���ͧ"X�%���2��&Re&R���,����"�Y��ͧ"X�%����;�ND�,K�~�fӑ,K��=�siȖ%�b�;��K�)2�)zw����q[v�W.f�iȖ%�by����r%�bX�g��m9ı,O3߻�ND�,K)n��L��I��I����>��q�	d�[�56��bX�'��{�ND�,K����ӑ,K���_v�9ıL���x�_�I��K��O�DZ�6$[6�ċ�6�����C�y�uss��ɺ��zw�Rjb,��]�����7���=����Kı>>�ݻND�,K�~�fב,K��;��ӑ,KĽ���Ktj˄˭fӑ,K���_v�9
� :���
���q,K���M�"X�%��~��6��bX�'���ͧ"X�%�~���Z��V�"P��/�L��L���vm9ı,O3��m9ı,O3߻�ND�,K��ͧ"X�%������ �\M�{�����n���O;��7�O/�w6$�H�����pPR�K���)2�)2��Ѿ�I,z5��Y���fӑ,K��=�siȖ%�b|}�y��Kı=���m9ı,O3��m9ı,K����5�n;��-Ư���p��ݽn+rxh��ki�O8���Wm��t���Y���r��{���ı,N���m9ı,O}�}�ND�,K��{�ND�,K���ͧ"�oq�������]G-|�}ou�bX����6��bX�'���6��bX�'��{�ND�,K��ͧ"2�)2�;�'�[n4�v�m�,�_X�%��w�ͧ"X�%��{��ӑ,bh�B(B<��!��7�_o�iȖ%�b}�wٴ�K�2��їrݻ �hn�e/�L�ı<�{��r%�bX�}�ͧ"X�%��o�iȖ%�by��siȖ%�b^���WXC%�5e�e�fӑ,K�����m9ı,O}�}�ND�,K��{�ND�,K���ͧ"X������1��N�z�H�]:��ۑ�vLvr=G�\�M'E�̺ܺu�HtBr4k��Z�ND�,K�~�fӑ,K��;��ӑ,K��=�siȖ%�b{���6��bX�'sӹ�ufkY�V�ִf����Kı<ϻ��r%�bX�g��m9ı,O~>�fӑ,K��߷ٴ�Kı>�D���fj��Y���fӑ,K��=�siȖ%�b{���6��bX�'���ͧ"X�%��}��ӑ,K����^���ֵa��ff��ND�,�,��N���r%�bX�}���ND�,K���ͧ"X�� 'P�uȗ�o�������{���?������^[|ND�,K�~�fӑ,K��;�siȖ%�by�����Kı>��}�K�)2�)w}��˲8��;��;�aal�]�rp��:۪6{�v��1-Z
�րN�0#o���7���{�����r%�bX�g��m9ı,O�>�fӑ,K��߷ٴ�Kı/;���nݐv���̥�I��I�������Kı>��}�ND�,K�~�fӑ,K��;�siȖ%�b?{S�w cv��"9s)|Re&Rez}�ͧ"X�%��o�iȖ%�by�����Kı<�{��r%�bX������54a�Xe!u���Kı=���m9ı,O3��6��bX�'��{�ND�,K�O�ٴ�K�7�������R��������ŉ�{��ӑ,K��=�siȖ%�b{���6��bX�'���ͧ"X�{��~w{�������~O���H  S��uvuC��f#��4�c'�{1��6L�Xv3@狭����W��C5F��ⱉ��vK7i.�k��\�SqW�$��kWa�"�{7c�N�z�nӏ]���6�J�ǡp��Lo��:�<ev�� +�&���A�T���lu����%�y	c;�k^6������,��t��rDgq�97U[�Xā(�λ�{���w{��׋f�5&��:�[���)�^'��]�9�kv˰����>ѷm6-�j��]1��O�����{��?g����r%�bX�z}�ͧ"X�%��o�iȖ%�by����r%�c��~[���'���W*��w���d�<��}�NC��"dK߻��iȖ%�b{�w�m9ı,O3߻�NN������;��1=Լ�����bX�'���ͧ"X�%��{�siȖ%�by����r%�bX�z}�ͧ�&Re&R�w���m�#��v�ṛ�,K��=����Kı<�~�m9ı,O=>�fӑ,K�<���e/�L��L���6OKv샴]�乴�Kı<�~�m9ı,O=>�fӑ,K��߷ٴ�Kı<�~�m9ı,O¨w���kZ�$�kT��-A�u���wc���y�q��Wn3�U�qs;���|c|)�H<%?=�{�d�,O~;��iȖ%�by����r%�bX�g�w6�Ȗ%�by����r)��I��}��vB�,.(Нٔ�ı,O=�}�NC�5�I?�]<�Ȗ'3���ND�,K����iȖ%�by���6���%�bw>;��N�湛|�}oq������~�;ND�,K����ӑ,K�����m9ı,O=�}�ND�,K����YX.���O�w���ow�ow���ͧ"X�%�����r%�bX�{��6��bX�by����r%�bX��a�wn⻻b��I%̥�I��I�����r%�bX~��y�m<�bX�'��fӑ,K��=����K����������m�Χ�����gXݱ�V9�<�n*$"�M��MϚ6"O������2]�[���Wr),�_�I��K����r%�bX�g�w6��bX�'���ͧ"X�%�����r%�bX����~� ���|�}oq�������siȈ��bX��~�bX�'��o�iȖ%�by����r
�b�I��;���nݑ�v�%̥�I�bX�g�w6��bX�'��o�iȖ8��`��7q>�wɴ�Kı<�~�m9ı,K��gn��K-ѫn�Z�ӑ,K F�����m9ı,O=�}�ND�,K����ӑ,K��3"g�w����bX�%��I�kQ�Xh�e!u���Kı<���m9ı,3��6��bX�%�߻��"X�%������r%�bX��5a�zaM5&��-ˆ��]��.�v���ɂ8E��q��s��\��������H1:	�����{��7��������Kı/����r%�bX�|}�ͧ"X�%��o�iȖ%�bw����i`�i?=�[�oq���~���r�(�DȖ'zw�ӑ,K������r%�bX�g{��r#)2�)n��v�WwlQ]�%��/�,K�����m9ı,O}�}�ND�lK��{�ND�,K��{�������{���?]�����^[m9İ@K�~�fӑ,K��;��ӑ,Kľ{��iȖ%��A���G�N�2&t߼�ND�,S)ow���m�#�ݻr̥�I���'���6��bX�"�|���ӑ,K�����m9ı,O}�}�ND7���{�?{���ѡ�v�����kKۜ�p��gr�Ύܘ�՛�����F�(�� �-۲!�.��\�_�I��I����bX�'�o�iȖ%�b{���؊�%�bX�g��m9ı,K��<��nՍ��yK�)2�)wO�ٴ�?ș������r%�bX��~ͧ"X�%�|���ӑ?��)2�����]�E�`;�)|Rq,K﻿�iȖ%�by�w���KRı/����r%�bX�}>�f��)2�)zuzx��.�In�ṛ�,K?"�����m9ı,K�߿kiȖ%�b}��}�ND�,Di����K�)2�){l=�e�mڹ�e�K��m9ı,K��bX�'�O�ٴ�Kı=���m9ı,O3��6��bX�'��# ��ܸ�|A��0� ,RA�D��Hh�YRJHJFƐ%���>��ѩ�D��jf�6�6HBH2@��L��8 �)YI� ���F��� �捠��I()@C�sR!FBc)F�+�n��*�@�I0R!�S	C<�y����%�yB8)
A�E��hR"B(�	<�e� ��$�ئ��qb�t��������׽��?_��`  p �`      ���    �PL�,ڤm�Y�S[նk���������+���U���l��g�ZV�ݍ�w7�Ke��8�lӺ�r���*�3ujmF�ͫ`���b�/=���sdrɌ�n�c�s�=���*�c[r M <�2����!S�/[�����%屋]Qm'N�g4P�kh�59z��*x�:�$��y6�8��>�f��j�Xc%gt�[�)�m�`��Bfa$WcRsm�vz��9�a��h8�P��K) ;\U��:Ure���P����퐫mT��j�Ij��62��J�U@Th_=�Iv�+��%UrA�UG$���ΨDi��dd#9�[���U���Ғ�[���VRV�U�a��q�R�e픒h�X��M&�ֹ�N�r����6�c=���m�4�l�y^���s��L�:��C�g�'��c�:�l���1�g.�L��3v���χ���S��'f瀩H�GAv̤��US��殫v(�k�T�x�V�6$�荞�Q8�gb�^�UM�Sb�
���7)f�)� hZ�	Fإ&M�]zM�ny�ف{�������ꍙM`�>���ګ<���	��m�؞yP�U�yS)��H��9��j�vڜ ĝ�ĝ��.�9%m��mۄK*�UP�-�m�E�Zt렪UU0v�;`�l�o l��\��ARی��'���[��AEm*ʹF��od�9�5UUɴ��d�c�elax��e���
����"�����j��Α�Ԭ�2 �7l�j��Qڝ�A�����{8rId��ڻ89Q���j�bR�H�Rzઈɑ�2m���`SOa��H@m��]v����ڰ����@V� [Y�k������Yې�Z'�8��#�����nʲ:mt*�Z�lh�q[�;mrk5��u�K��숌�@<Aj������6
h�{����wsZ�� l�$��ج�����E���]���ɺ{S��n��u���N�]��ݛr,疎<�pą��-�g������p@]v�\�1K�׵vJ�9B����v9��Zw8��e�l��c�i�Tmmڽ�X�G;@���9{G83[�mNQm�A�2���#h���۶z�>��y(51�<L�)ѳ���n�Ӽ���k&�潺}���Nw7X$���Үq��k����5��%�\�[������|�U�{Z.f����,K����m9ı,O}�}�ND�,K���͈"X�%��{��ӑ,K��{ܝ����h�F�rfjm9ı,O}�}�ND�,K���ͧ"X�%�|���ӑ,K�����6����bX�{�fsSV�˙n�T˙��ND�,K��{�ND�,K��{��"X�%�����m9ı,O}�}�ND�,K��m�{��ku&�L��m9ıP�/����r%�bX�}>�fӑ,K��߷ٴ�K���{�ND�,K���;��cq8��)|Re&Re.�>�fӑ,K��߷ٴ�Kı<�����Kı/���m9ı,Oԗ��L���Э8����Z�m��W]nŹͬ\Ȝ�nץ��̢p��?;�>ΟBv��`;�)p��L��]�g�)|R�,K��{�ND�,K����ӑ,K�����6��bX�'s�٬���H]�r̥�I��I��=�L��|=S�LA!Ȝ�b]���iȖ%�b{��}�ND�,K�~�fӑ? �TȖ'�蟿j��պ5�k35-ֳiȖ%�b_~��m9ı,O~�o�iȖ)bX�{��6��bX����ze/�L��L���]�p��b��\�ֶ��bY�H�����r%�bX�����ND�,K��{�ND�,[����ӑ,K��{�N�\��4[�Z�356��bX�'���ͧ"X�%��w�ͧ"X�%�|���iȌ��L��7<e/�L��L��wg��X��� Ě���y1�D{m��v�.-a��t$���]և5W(N�+o����L��\���R���L��|����m���� w}� ��i���ӱ��M���sPǰ@{���b ��RF��RM�t����Y�����������rI�}��n�K��`�v`~�T��;�����b �9�c� :�˼"�C��9�mz����t����S@���8�&���f,�,�u�/m���\�]����az�7�Ƴ٣-ĦH�j	H��u���M�t������D�I"1䘛rhǰ@{���b �9�����U]��V~s"q7��"cp�=�~4���<�Sg;���m��9��2�H6�qcM�h+k���h�4:(n,6"�C��y�w��rI�剟�
�8����h�4�Қ�����QJ&����SvA�tz��l���:�׬#�k�7
�p��Ys�� �8���;���{�I�����n���(�r��;zg�l���0��^�:�h;+�i8��&7��h)& s���UU]�O� 9��@G�[ӂ�#��%#���h��s@���0<�S���0�Xz�ۅ��[�y���n�T��=��$��sw$��A>�$Ul�w�Z�Z��:���k�in��H��&�'G�G&��D�V��v�ݳ�B,Yvv���	����5�b��܍��Y�nu;����P���汧acqvݵt�qsS;pr���rp�QIc���׶�F���	�#K������FK�c��(5M��6D݆�8�ݠ��g�8N�gu+]��*v�뵷խ��m��RLі�5�ɐ�5�z���{<�}���.Մ�`��:^�{ vzx����̚ݲ��u����tq2M����u/5����_�绳 >�v�%�����^�nh���Dlm(�ƛp�>Vנ|�ݘz������<�%M�;�=e�"��%˘w� �Ww�o�� �[^�w��f ���M@����~���R������1��1 t���4儊4'-`s���\����:��ӊ�9�M�¯7h��j�V�ˠN۶4W����`m�tp����3��Y� 񼑴ȤKx������ـw����0�v�`؏z�nX�w����|�ݙ�T�ޮ�,���|��bE���i8��ɒcmǠIS�Hs� =rL@z��@F��*�qG��#x���t����^���W�{����uȐ�J8����& >�s��T�R��t�~;=�NӂU�6�<���;�ݵ�^9�۞�.w�ݛ�l��[e��NZ,�-����@z��@s� =�`���1 n�5�m�tZ�Gw0uwqg�T�g;�� ����>|���%J�)߼���h-�	hNZ�;��������%�X��J�IU}�}�L�[��N��ciĤK&7��h.��/uz�;��?UUR|����[��V��z^����bΜT��=����m�;���zШd��V5	�����wn�Ǌ�=�k�v�e9ĺ��;m��tl�j���ݵ�Y����O� =�`���3���[�L��~�,r��i�R�N�`s����v`>wf�WwR�_�7}��"Clm(���p�9~��z�ֽ�λ��Қ����
	@�����ـ}��ŀs��0J�%�UI/�_3�� 7�a6�&7tZ�Gw0:qR����s���1 {����t�v��\��.��I�8�I�y6^�v���x�юg�*XƯlujN�e2����[s��>���>T�>.~y�6�JD�1���>]k�>^������9�ޙ��*��gZ7�nX�.�c�s ��0uwqaꤕ7޳�y_ߞ�z�,�92H��&6���nT�Ԁno���������ܑ'y1)�7�L�=��?y�ޟ��z`����?-�)מ����U��&
��ml�\o{p�B�絨y��ݹ ���]m�]:t sklpP�q{r��%�P!�1��<\�]��qT���*O7��N���=�rD���ڧ����ʺ*22s�48�/@�kRg�mɲX-��m�AA�۩xE��f�.MJ�r˴�냳�m����1��qȝ�Vr�0=&�px�-e�ۀ�v���m��>|~u�&\����F�\�QcpOUm����d���`�n۳�F��ȋ!�6�qcm�x_���>^�������a�����S������c�G.`>n��IU6oM�,���|��3�a���!1���q���n��Xs� =nL@z�L@Ԇ�U����3 ��@sqR����Ɉ>�i}�������q)��4�h'& =nL@68���HT�WSA;l��uٺ�;�=��K�����u����ϴm�=��������=�4�K�Ǿ��;ӻ� �{��*U_0��zh�~�~��&I�$�ۏ@�:�jʾQ_�t��vo����<�w��'/���$~�R��"N(�%2D�&ho�Xϻ�ԕRo�}�n��X9�&H�6�Ҏ,m93@�u�@�u�@0=IRO��� ;�N��q[�;��|��0Ԫ�n��>��ŀ|�נ[��$XbqG��7$H�u��{;�p kc�u�����hWɵ������>F�BS�Li�#�K?��4�Z��Z��-$x��pC`)f����ʪ���UR~��`~��`�Jh;+�L�cCs4��}��r��ٹ��!2��bC�T%
��*g��"C�@�H��[�	�	 �$���1$����03�0�d�A��t� � " H�#�� �T�F�AD�O�(6Y& -�XEI��J�"�Oվ�@bC�����A!��z�n*��}C�Q��}47yɽ}7$��~ٹ';�8��\�H�˘J�R|��M��Ɓ��M�mz�adjI�q�jI.`��� �K����<�~���Z��c,���ĲI��Ok�.�cF�	��ɹ�����}����>��-�m9D��qG)�&'��g�@�[� ��v~UT���t��w��e�NF6�q�i�h+k�>]k�=�Jh�oL�$�M�{���r���;����؀�=��� =rL@:�m�LnӴ�m��U*T���	��k�rN_��7 
�0 +�Q(�
���6�P�������e��D�6������� ����>}ݘ:v��=I%K��7�۟���Gkn*v�q׷B�5�7ih��N7��\�q�������w����-�[f{� �����& 9�`��Қ�h�n$�8��)���^z���gt��wv�`=ݘ��6F���	16��=�Jh��������z��[�.ۖ�+Mږ���ws���z`�ݼ�*Y��w�w_�ܑ7�J2��z䘀<��1�����������  ���:XZ����d�d�V�B-�����jy��v��m�:s�ܮ��$�M5�y���v¶�)�ڔɵ���x���$��u���;K/���K�7��+8��q���j1�]*��u�F��훝��  �6�v!:˺6��W�R�7ir�)M���l9��qYT����F0��n�yY��=`�GM��!�$�Z�J�<�.�\�md��Q�����
8v�o\��ۯ&&ٴm��Z6������wc��9�ڗa�.�n0���Pc� 9����ӐՆĦ)�4)&��)�{�S ��v`���~��U~��UR|�~.�unXH�;� ���ـw�hqҚ^��Lȡ41�RT��'�� ����>��� ���0,:�4�I�q�N=��^��*��i���9�~0��f�ݛav�׵�CۮQקI�m�R�{����sn�`��KR��X�I=Pk�p���}~o�7�@z㘀��19��7n�]�C-Kpr�����I*��^J��j}�I��<ǰ@{�1V��Y�r\R9,�>{ݘϽه�URo�m��=l�h�D�p�<I�)��=����>��� ���0=T�'�����S��B�v�� ܹ�}ӷ��W7s��q�}0�{� �؟Y��h���c:��*�ż6�8�3��Dud3���	l�]���ͩ���(	���m���~�>{ݘϽ���U|�z��`}^�.4�$QcC��>W��>]�����{zg��6u�}��%��ۑ7���>��{y�����adj<�$L$�܏C�g�+�/�z��h+��.���JRD�Q�C��qhs�����uzyN��?%J�l[���`�V��n9p�������`zm�+��nh�,�'C�crk��;��l$M���mA��^�����.���>�@��U��Ƞ�'������1}_���'ր��@z㙠���0�%1Li�N=����>��<��� ������K��[���28���Z��z˺�����V# �VmQS�����@��W��&a"��1���1�nb�c����- �̚f�Wny�/=[��藶��7\�]����4�Ŵ����8�0�ڠ^~m�������N��>���0���`����⻉	17#�;����}V��^���{��"�Jci1�&�&�s���@5{���}V��u[$x�CiFF��Z��z˺��U�}Ϫ�z��㉍9�L��.sf9h<r��� W���U~�߯��H �`7d&j��UR�<�.wc�Ê9wg:��î�'m�۰5���d(��N��H��lV�v]9e�z�,��F[[A��cÇ�S:'F�V��uΜUY����.%繸-�m���6�49�g7m+GD���X�;�=S<���َ���EnѽR����٧��3;(���\n���V63���8�8Nq�Lc՛څ[�����z��F��ΉN��nK]�)8���X#\<�젦��Ǭ''n��p�bu���O����*]���g�Z���9�[sݖ�<_��&�OZ����z���^����*�WH�f(��qh+��.���b^�������ya�q4�m�	�iǡ�y��������>�@�^�@��,�G�D��L��p����M�z��ֽ��\&	�$L����%��t���x�,cpۓmv�/���r��Γ�"�-��[�9�&8��_��Ɓ�^���^����=�VƠ6�Ҍ�1ɚ���Uvu���c�����ձ�j�j`��@�u�@���i�M�wذ?o� s��{b*2Ӵ�n�q��6}h'ʐ�� =nL@vZH�G�I<Dqh�w4���.��p�� �Wa#I$�������]vx�&�A�c�=nO<wNۊrz<n���X�����z�˭z�>�@�[��ya�q4�m��Yy���rb��-�EH\q����҄�b�$�z�>�I<��ni�ج��@�Ņ���DZ��(�0�����|�I~�����u�Ly��K�廖�V��9f����� ���`]��qҚ��ljhmF8�%��>{ݘ�*��{�����`ww��z��1�#o$j(LlJ��;��q���'l۱8�}���ޜ'B�7$�.�h���[sc� <�U��Xu�}0��q��Te�i�ۗ0�v�@yȩ�b�ɋ��å}��Yn6�Lwf���`=��?$�}{���=G-���o��DĘۙ�|��0>���9IR���T̀�~@9����rO);�����fZ�M�N=����}V��Қ��zr�$I���&E�$C��7$�>2v�cb���+�N�;�������;.�$�C-K��\�i7� �wq`>n��U|ï���=�7~.ۖ�ZmZ�"�� �9h_I�\���_~��vI?-�@c��c��8�˿~z����%4��h֤Ӹ�522`��`)*I�{}0i7� �'u�~I'���������j�H��`3��r��� =rL@*�߫�_�Ah�
k�Ү%CzҺH8 @
��th 0�0�HT#H`0� �C��GJ�j��C�
l�3L<�j)�/*��)���H�(@�4R���w
�@�	!tZoH��q�� ��mXR��#T:{�wN�����#��6�  H        9��    ���w6�[���᎕8�*���+rmj�<�YB��$]��]c#��w6�sɤm5=��WH���Hqخ���`6��ڧ�@W��u9�;Te���۰Yic�����T	u6�!��[^��bڈ�Hn���g*\m��Z4t��*��ؤl���`Ɗ����R ���Gml�O>P	MРEʇ&���4�(�$�gE�*����n��� Bt3@��Nk�a��l�uĆ���\�s []m+K�&�؃��A*�5U\=���ջ/�jm61]�)�U��U�t�m�k� ���ȷ��m$���3`浒�6Ԫ׀�6�^�r��g���3��Z�#P�
��k���[�=8�v�/C<[�ìA��Mf{[����l�Xy-3�9�b�8�'���y�}���ް�k��E���(��YNv��*˘�+ma���b�JU��K��(WX�T�m��g��+�6�Fץ�����G4�<m�4�� N�<���v�+��mR��9#"�!<��[V��R�k�B��ER��SUU*5�[r'�"��nv����^W	1 D�.��
=���<�����Dp�l�J���<�'�8ɳ��d��v�p ׫m��;T�M/h�l�i�V��k�#^ۍ������T����UUgt!�<�ϰr�΁�+�Z�A[;��)�ՑZ��wim��[J�F��f��t�6��-[�g�6�nS��vCn��ףR����Htձ���ԗb�m���N2s�`����mnU6��z��Fơ��<����nI��p�2�=����p�b���q]l�4�9H���0
�Ya��[<�>����ѹ]�k���'K$���'Al��z]TH��=t��Ǖ����c�g�yU�@K*۱:Z�G0S)�<Z�W
ZV�ۗC53V�54g�!�H�b|�Z��P����@#F��b�i<EOAD6A牣�E��'�/����Z�Zֵ�kY�UNM���ဓ�#����:�ڮ1rY�9�sϞ��Ɖ:��Ϋ�"�%%Nx��m�z�tvݬ�&�v7j��`�ٖ�r��Bm��%#��[.�م;Mǭ�^E���u���<:�J���{b����ƭ���8��B��:��b��%1h�L���y��gk��.yn�5ٴ��wWX%uj�z�B�m��M��A��r�ઘ�V9;y��g\=ut�����q��;��B�ٸ��2۞�w힭O�ě^�;V��^����K�%��=������Kq�v���Kݴ�9��� <�r�y%��~�H��D��RA7�8�V�z�f��;V��^�oL,�G�D��49#���4��Z��z�>�����S�"N(�%���nZ������9���7Dή�K3�1pUk�z���.㕑!vѰE��f0�O!��_#��yIΕ�O� {���9�v9h�[�j��#�p�;���;����I	F1 ��H$#a	H�d @�X��_�߷Bئ�9㖀��1 wK���ĉ��ܚ�f����@�^�@=�@>촑���`��c�@�d����1 w9�>�wO���?Ì�#Di&9"�>W��{���u��v� �UŎ���$�]��!�*{^%N.�E�U�m�@�����3:���&��7j)�ō8��_�@;��hyڴ���zadj<�,Q�p��� ������9�_9��$~��H��H%��&��w��N_��7*���$$*�~����k˯�@/e�@��V������̼�@z㘀<�� ���ߪ�K�������~Q�dv��C����� ����Ih\sM��ιjMצ,�m^9�M:_�x6Nvl���5���Ԯ��7��|~~[��5�e����}�<����UU~���>�럿<Y@M��ɠ}�ՠ|��0>�f w��y��<��x�
.\p�������8�ݘ~����^��~Z�wTA��QH8����f w��xݛ�r��*_���=0z�?Hԓ$`�I1��w���>�)�|�W�ywW�{�2�FF�I���Ԑp��[���]�Ogt�sHU��>���k/�D��X���U��l���������6=q�@u�3���u>�I����3,mF8�Q�@�^��$r����^�v��~������d�;N�h�w0~������&����� >ް�b�-Z$m˘���o� ���`=��~T����L ����N��	�94��h+��]��x���g�b���4��u������ 7Me�L��nطl��mǳI�ʒ/�r\�\sθ���Y:�ٷ�Y奊9#i��Ӷ����z��+:��Y|�)�l[�7`]�j�5���82�Y����;��s�7>I�$Ůw;�㞧vȔ��%��C`.�v�]2���'V�.	^�ʭ0r��n{qW��`M��ʪ�����v���+�F9K*z�}��:��׫v�3��S����v��7k�v���Ŝ����kkr/0��]8(��8�hb�*�����]��x����_0��y�h��!%����Yy����1 >�5��-�bޘY�0S$��@;��hzn�=J�7����:�}0�[�.ۻw0��&��;V��^���C�%T��o� �w�.\Q��܍ۄ����f�IU$�7}> ޭ��vw^m��;�Z4g��&	gY��<�np��f�9�^Tfͣl�hG�mf���D��d�����@z��@��@{�����ް���`}�'�Ceթ#�� w��K��eq���Z۟b����R<Y0�ԏ�����z�?�%M��}0z�׀k��Z�.]������1��1 >�5��/@��7a$xӏ@�{��=J�{վ���f��=����&�v�U�φ!���X�{m�� v��]�{Qڎ
�Xz�{sv�[�Gf��v�$��9�v9h\s�s�6����%Z�H���'u��I&�?o������u���5�����`=������וR��R���U�轗�o}~0�;�;���.������� ��@{��@z㘀=N�ĉ�1���@;�f���U�|�W�|������\PpBn,`��1B�*�Ÿ�Pi�;W �g��F�N׋�������9��6�nM�>�@�^�@�{���Y�U��D`G2&^�����s4����c7��ى q'�H8���u���l�>��+��م��&8��]ܻ���I&������<�{�$碡*�
#U� P�o�s7��)"R)0y��&���U�yov`>wf w���yU*Uطg���(t��S&z�C���!��>���{��n�=XfN1�7���L=���叭����� =|� �j����e�񩈐$z��^�w���}V��z� ��5a�1dfLM����5�{\s�s�Hn�^A�(�ԎI�}��<�W�|���z٠U��Da��%!�z㘀��I�s� 
����%����sgK��IN�۝��-�ؗ�Nz=-�ٴNܫ�<��)Ne)3N�O0)�s����a"V��o!6�9�ơ;t�և��7����=�����.:�����=�HwUՁ�튶w[%r�*"v��y�'i�V�O �m���kN��V]�&0�a�1!�tv��s�π�6��)�z�v�qY������rPj�x *m��[M��K�m����ܔ��;6��^z�+]t��l��d����q�-�]��6���ּ�a�e�ڬ/#��;�� �j��\sM��ӓ�S$��@;���u��<�W�|���/�)IqI��7u��\s�� �j��q�lq4F�&hW��>^���l�>�]� �9�Px��Hn� =|� �j��\s]���o�>hWj���6�A�u�u�:�^�ʈht��xͷ©���[����u�^f� }&�=�*@u�1��1 }ԪG��cjG$�>�]�Y���*�K����#��0>�f w������ϫb�"')�I��9~�����W��f����h q&dMcN=��b }&�=�*@u�1 �Q!�y&6DHI�H��l�>�]���z��^���s��$i���%�^���M�ͼgI�����q��5�n�{p�lAZ���H`�ܓ@��w4+��/uz޶h�q�lq5c�4(� =|� �j���sos.�� rG�|�����G�g�`hb0�U%l�j!p�p��0"惘ȄЫv����h@*�B��
0�E(@�� ar`d��9��
(�
,�K9i!���Q' ~���CK�C���M���j��WJ�"�E�!��O��q T@��k��B���
�{��nC����!��#2bm'�w�����q�@zۘ��s3r�Lq�1�#�hw]���z˺� �7o �T�7��[,.!�Ev���]v1ܰ]�EvW�ぷ�+ۭ���S��/"��')�I��_��|����v�UT��9��Xn��Im��Wyu���[s�5��\s�Hӓ"&I1��w����s@�^���@��$I�&�Iwx�T���X_�� ���0>ƿ�1�-�uR��'��&�ئ��9��$�<�j��H���sŲv#�R[�k����;�n�gvy�s&���l7oe�^`Y�TJt��j�owm�nb �&�<�T�����j��f)������f���[�s@�]���uz��[�1�F�e���<�T������t����tq�D�!	9���h&� 	�j��HX7,�3o2����ʹ���t���qR<r�$��<*��9'��I�kZִ���IN���m�&Z�:�Z7f�ӝk9���)��zSLƺ思�\�/n
�Bgt���/5�b�r0�B��{[��tM�g.�%ܫ��[����d�	Н����f�F��s�k�m��h�W���&��>_/�M�Q�Ñ��
�� ��\K�\�]�m>�cc� ��l��g��v�H�8���pr�����tݼݦ���2��Z7uNM\�>.��
����|�%�m�b�m쫨;t��4��Bwmnqtuٴ�eѮ��v��}�7 #�- y����a���L$0pnI�}�w4Ϫ�����f��T�6	�#��F���G�Z �sP�5����ݍ�<jb$��@>�@/����s@��� ��5a�3�s4��	�j��H	��=m�@��ۘܵ����sH]]/g8z�<��ކN��8�"��n���,�ngJ)M_6<�T������s�����e���nZ�7����RK"J����@>�f�{����n$��[�$��o&���v��I$߷}� ���ZsîF�����Š��n*@N�-;$���̽�L$0pnI�^빠^}V�|�Z}l�>�GQ�C�LK����ئ�7�V<�edC[V4l	n��bfg��_�|q�O	m�I����h�ՠ�������=��X�k����%�]���x�n��RI*l=�z�n���ן�6��?YD�N]�oN���rO��훞��~���(�z�j�?s��hWUN<P�M����㖀��Z �&��f�q�����7-`��x�Kݿy���׀o{��ʒ�ח��A�ta�K�=r�:���]�z������&L���Bx�ݖJ�s�F���]	��������>`/����h��nFݫv�-��v��M���,�7� �v��r��7"��@q��h��9h[��T�}/f^�"\��7v�?/ʪ��g�<�߿Ly�� IR�R�T��q`7�e�q;%�˰�wo ��v`�RI{����:�ۚ��h���	�����8�T�]/gq�a6���.8����� đPpk�ߕ*Fe��eN�Z$n�|��b�=�w4Ϫ�>]k�>���x�c�&�M��=�w4Ϫ�>]k�/���*�Y�5�R�BNf�y�Zϻ��U*��UI�~ŀo�����ĘI�4Š|�נ_[��{��h�U�w<:�i�8&&��y�� �RJ����{f��>�̒��{������?���Me���ۭ�vn���5t���C�]Ͷ�ۉn���$n�����l'cY]䒳	�����ڱ<&�pu�
��V�%ׁ㡗j.6��y��@��6:8������SLn:L\n^A�\�L��d�Y���{!�@[mԼn	����Š꤆�!�j�BiM��fn���i�����Ц�1��0Aۈ曷l�����"�#LGj�.�&l��u�fܝY��n[��[��Ong�;&�ۗ]��w�	���պ�4��h��ٖn��~����x�=nL@N�R���{�\Eܹ�7v�����T�l��z`������s@=yW#O��)6��& 'H���H��@a�#�sґ���h�w^��$�7ޘ=x�VKR�y�������x�=nL@N�R�q��`�1 0C��X��:��M�n��s�';��kr�=4�]WJv��1�k ����>}ݘ�w�UK�o���-��7y&8Ʉqh�&'_�U�}=���R<r��r4�ȉ�i��}n��빧�T�M�f��{�L���.ݧuj\�-`~UI'��|�l�<��ـ_[��w���О8�iI��r��& 'H���H:{�7oAqv��7L��t��8S������ɺ�6mx	�i$M���=��{��/��uK�b�o�uϾ�� 9����ܽ �����S��JG�w�d�{�4����ٞT��6s���q5d��9rZ�;��X�w^$��IRP��@��s@���F�H����x�=nL@N�R�U~��r}�@yao�1���1�L#�@�u�@��s@�u��/>�@�ջ�1b�b��.⵬�̽��J�<����=�,�9WXl�u]?� ���amǠ_[��{��h�U�|�נw����&�Թ.Z�9��,�RJ�g�o�Ǿ��/���;�J�hOM
4���9h[��T������ܼN�-����yU*T�7ޘ��b�9��,˪�U'IRK����氞���S16��@��s@�u��/>�@�u�@�^.E�I��4�b��A�����X�(m]��u���>�ae����5<Y1Ɠi��h��h>��ԕ*_0�}�X��O#E���j˼�@G�Z���� 9����7xI���>]k�/7qa�R����X�o���wl��r
0�6��/���=�w4Ϫ�>]k�;�GS��I����q��=�*@G�Z�$�� =O3���K�+ǎ3vb�"�AP7��E�62��#r�?� �5D�!+<<��2$�"�&È� FZ[U.	U\n�`F�P���|H�`0��PlD���]M�VŊ@��:�`b��D,d
R$H��X@3HF�4�+������0��BX��Jb�x����V($�{���;ޝ{���??�  	              m���amZ�X�s�8�Ͱ��U��A�������OH���-������/����f�R�D<��M)���p�[g6���I�j��P�֌�q�����3u;J��[�$��l,b�gS��.�.�H�u�KKs�&�ۚ�G�W<ޖ�6Z�e�mm���R��g<=Y�ȵv�y�K�����y�EuSfw) �벍j���lc�=NX�n��ˀ�X�ښ�;j����<���`z��>|5�'�Ԝ���)�N�m�M���r�c+X�w`�H����uҤ�"� @�m�e�{Zٵ� H����jU��ۜ�=p��Q�!q�<�r�H�塈)j 3�j�����gq��{3��.�*^V�`yH��	�C�A�iA0�rs�,l�S�k��e�W"�Eq5xƋs��%,sk����o��xx���]�����dR]P�:���Çu=��3�ln�̆�a��V�:�J��F�j��'mˮ�:vUV�m/ϋ��GC�n ��ݜD��m�����Az&�M��e%c�5TU)����|�h��Gm�4�k[I��[��ٗ��-k	��Zһ7$�i��^�j���y;#�����U�_7�Q�kl��ۊꪪ����� V^y ��,�Z�t��Dؐ-� �u�[�R�v�^NU�m A�]�BȲI+%�[*�KT�=�,�qhN���N�jꭥZV\���]]� ��gM˲�e)���J��"n��U^V5nm�۝�]Cm�ʴ����R��#��%����q�s
�ӋsJ]9��+�F��ݧ
��)���@��L�@r5�жӎ=� �,�쫫�b{g�.��]�T8�7R�;S�)eq�٤Ȫ�KQM�pX�ͼ\S��u�{* �*���ldQ���%`Ŵ��:����	\J즭�WY�kX�@��O� � ������Eh`>���]���i��  2�n�΢�c:�Y=Z'����T'9�����,��]m�i�3r����`����NR��؎�J{f��2k��w<V�Id���t�t���bv���S�:�/m�1d4�Ҭ�[2��F�F�iw^֍���o,lF�0N�h�1%�M߫֟�P�O[v֐x��;<Y���q=�zeᣋ^GU� ��������{��}|~�h��Ѯ5�Y�t;m��pj�}����74c7n:J�F�#z�=���v�>$�<d`�JL���-�mz^��w]� ��r4�AH4��-绳?�$�7��X��ݝמ���UU)y��eN�-9˘�{�,����򪪦��|�?{� �a�H�d�1��m��;��h_U�|��0?*�J��o�X��O#E���"˼�@9�Z��}�x	��R�������mO�mǜ���K��e�䐺�9E{A�]��v��������3�z��(��@zܘ�q�Hn*@9�Z�����sǑ��z^���31J��u~UJ�<'����ߞ����;�K�H��LrH�hW�h.��z�h�j4'�R�wk�URT�R������ ���� ����=�w4�U��8��4��$�ɈT�����=]/M�g�Nv�	��º^�;�lu��p+�eΧ;����]�n Q�r��[��\��@8�7 �/���W��w��� ;��������؛I�3@�u��:��@�u�@��s@���#A		ܵ�wgu�>��%%U%*UąM�%R��H�B,B���T Z�������빠|���bpX�L�x7ꤩ~IN߿~��{�,����;��h�9܃pndc��n=�]��w}����<��ـ|�6lV[��̉v�K�����ǧ��Ӱ��p�an{u��Mz��������g~I?�����1�@zܘ�q�H��e�yA.��q���wgu��J�8�ޘ�}��{��h����()�$iE$Z�ɈT���v��R}��@��(bv�i������%O}��`��,�;�UU
��IR���ɀs������؛I�3@�u��?ٙK�|����z�h�������Ѫ�z���2]�DTtp=a4���'l��ODQ�4��s4���>]k�:���=�w4�z�A��8L��������ʕ6o�ذ��ݝV���-aB����mǠ_�ذw��ԕS{�x�� �:�mH��L'��$�f��빠u}V���^�׮�ުQ��<	��&`��x�M���o�ذw�� �����{��=��������H �`75r4Yi�=Jg�sò����98�4r�Ӟ��������^w\'[� ����'5�څ��!F�r5�,�4%u�X،S�p�6N�Y����;y�����k|��2`�=ƜfL\s��7���tfq�fx�Z�/p��������ܣ�3�]�W �{y6� �J.ͤ��ڶ���z�svz�{r��cn�>:���P<��^�8z��{�w{�fg'k���z�݋c�5-�7�Grm��9н��v�ݍ[mǖ�:h�QK�	"$iE$\]��=�]���s@��� ����FLncM%#�:�T���Wc��H	�O��rb�	׆F�I�M�������Z˭z^��]GIHE	9���=nL@8�~�nO�H��"ı�dc����Z��w4w]����Ue"li
dQL)�_��� �/kn�������_Fx����ao\���pnd��Cn?�������s@����ֽ�ʽ��I���$��X;�şʭ������{��:����;z�h�O�y&�)3@�������*@sqR ���ܼ����v۷woʟ&�� �m��9��-��ޢ�a�#&71�������H1�@zܘ�+���YB�6�[Y(뫥��nG�������a�UѴ��ݝkܚ�=�뫡k|�����=nL���a>�������8�,��s4���>]k�:����빠|�֢ı��c��xϻ� ����|*IW괨!RD(A� b�D3��6>g��~��?s�V�ݏ:���8����?����R����=nL@w�V� �Ra?�I$�4w]����Z��)�}�:��D�7;'%���(u��=T�l�핑!v��nC��P�P~�2��-�DȮ�ˍݯ��M�@zܘ�q��T�$w7w3*�Ra"J)"�>]k�:����빠u}V�{�X�?�D��4�R=�J`�w���o�Ǿ��>�n�qd���I�3@�u��:��@�u��]R�����`�M�.�v[�e�m �-�rb� 9���{��~���s��<uta/7�ˍv�K��cq.�m��lg�nz\{Gm��?绳�ϟe���M�(�������T������;��;�N&�"�z^�Hn*@9�Z���n�b�/v��uj������q`ٺ��*o�}�_߿nh�m'���$F���9�Z����*A�V��Ԁ>�_۱��
L$IE$Z˭z^����� ����8�{*�J�UO��y]��UJ�T�L���t��=������
s8���p��Kz�::ێZP)[F����c�4lw<[m�
�kz���O�[2�gj�q��
j]c��V��:3��b��ع��M�y������VL֣8v����#��ڣ�^^$e���l��Xi��
Y�Q1;s��i�_\C�]�n�S�U�<�l��Kd�5O�iܙ��/�?��y��.�Lq̓���w �Nۃ(���'��7.��΋�����\7��s����*@sqR̒��& :��ǋ�K#i&����s��$_��x�� �����IRl���w�B)�I9���~Z˭z[w4w]���n	�L�x9���f��ŀs��X��_����+�%�;�K�ww��RK���|��~Z˭zϽ��q)�� �CѰ�ܓ�[��Ok[<��ɸ�9.�J�w��=�S�񚻪����w�I��\�~�{��@�{��ݹ�~�J8�OD�"�kF���}wEP�E���Э%g�� �wq`�w~I%I�����mₓ	QG��~z[w4w]���h�E����LR	<JF�rEHn*@9�Z���L$%�ӎ;���$��s��X�%J���?���z`��X��NȂ�:��� �u\�������Z.Ɇ�lr�xgu�Yr�AB<��,�q�$����h.��m��=س�≸!�^ٔf�=}& �R��H2G��I$�;�-�V9nK�vZ$�0���ܓ�=�f�4��GK��0m҉�j��1Q�ā5����R^q�X$P�� ��}�8Bʻ!��_|$�@O@� �QM�҈dM"{@0��bh� 5҉=�(����OT�}=�((��
�
�I��,ER1$���5|* x�f:�}V���^��ʽ��L'��wwv�?�J��w}��7��xϻ� �۹�}Ԕq��!�"1I�Wj�?%T�W'}���{�wq`qm�h�qmd�7L�5�yy���x���<gn�Öf׶;�Ԓ&��q�m��:�m�����*@w8���a>Ͼ�;��(L����n�`��X9�ŀwf��>|ݙ��$�RR���i��26�m��-����:�V����@�n�^�^F�B@pI	��:�� ��v`��X�����HEQTU��� �y��nI�O;���j\�um���>n��J������;��,��h][�#)(?���F۝#�{m���>;���!ك�P���pjz�m�-�N&�	�n=�����s@��Z�ֽ��{�%"�	�$�I�9�ş��_��J�Cߧ�� ��ߦ����>�J8�O�L����h/Z���h�]� ���6�AI��(��@�zנu�s@���h��
����߮䓿~�'�F4]j[���@9"�s��d���������o��I  t�/2�ru��\ۍ�v-��R���ۮv{q�֎�3n����Aٯ4ٝ����i^ֺ@ܢY��ܾh�Tٱ��2G��E��:q�墸5��6�e�7,y����Z�t΀�\s;������b��s��S�v�ӦY�GQ9�ƈؖ6:U�J��*nnkn�U��|�٬47D�=*���W=v�!G8�e��w��8��6,�6�#0��c���7j�pYCh��<&�8`�J]F��#;���`z}�� �Ih_I�$T�'V�.D՗a,m�Z�;�u��*��l��0��� �;���\�Nܖ8�e�"]���ـwwqa�T�7��h���h�y����B`ۏ@����9��,�7^�T��'}�st��$JE&�d�I3@���h]�@�zנu�s@��\� Ʋ"bm똑�t���y8�����{���;8zJ�F�d.wNd����$��L�:�V����@�n��u��y;"m)0�%���ܓ�Ͼ��_PD�E�B����_Y��ذ�}� ��׀��LR	<JG�u�s@���h]�@�zנz��ǋn3$i&�4� �-��1 䊐u.#.�X���wf��=I*\����o�~0w�� ��f�wa%�u2\k��td��۳5��2�8:����H'�^�x�4b��(��hp�x9���^���hWj�;��;�N&��Ch����`���2K@zܘ�IU&�n�x�ۻwh��wwr����rO~Ͼ��C�C]O/��7!ץ4���6'��LNWj�>]k�:�M�Қo'dM�ۻE�n��xϻ� �T����,�h]�@��DX?��m`���X��Q���ճd�r*����×r�v��]�Q��濦GO��l���Δ�:�V���^��r�ǋn3$i&�D:{�%�=nL@96����I���?#.�X�iݘ�{� �u�@�e4vt���:�Q7cQD1ȴ�Z��S@�gJhj p`-��(<G�O��-�Ǖ܂q7&
�z[)�~J�$�*�����~8�Oߞ����o���_׭ �y�*^�K���`"�q��)'l�=�����v��Iڢ)�������d����1 �� ;�J8؞�0Dk���ڴ�wf��� �WoL�UU�UUR�?~�&��	QG�������SO�%�[~0��� sz��� �;�����woL�]�0��x�J��o�0�/x�d��]�ܗfήޘ�RK}~��=����ŀu*���{���W����nvΗU�T��<�7n���e��p)�;:�������(���cF�O4���i�ݸX%`�͵Z�Nɭ�Jv�ͬI<�ۢܙ*XM�P��ݶz��;�l�'9�.���KOO+j��}c�b+���Ѫ���l7&�Ie�&Uۊ����m�8س��<���d����h��v,5���.�(�\�K4h3�5�ɛ���f��">���;����~�	9gf�d�㢘s��;��8b|����b�WNW�ѝ�n1�I�j䴼tH	%�C@��-�ֽ����2��/�wVߌ�E����nE�d&�=nL@9"�:{�%����߳?�"�yB	�ܘ(L#q�����]�0���*M���x�� ���d �Ra?�H�p�=�Қ�h.���S@�U+Q����"5�ـo&��?$�R\��O�����9�ۦ���zƠ�`�M���`�%0J[lnڣ�[;'2���s�q����K�5Pj"�s�I��(��@�u�@�Қ�:S@�v� ��:��/�a1�R=�K7ClJ( BBE�2y�{��@�u�@�h�Ć�k$m����]�0��xyR�I7Ǿ��?[?{*�m$��!�_d����1� 9�� :���u���)2!��Z˭z��=�Қ�hʪ�D�
d�L#p��˾ �k�Ń<[y��v�))�Hq,@�K�?�UR�ke�9nK�;-%���ߞή��/��@�u�@������I�d��ݝ)�_;V���^�y�Zz�Z���b$��N�i'/�}��;�xD`#���`F�B I�$��+���@H!v � b��Qs�o��ܓ�O�ٹ���h�I��QG���^�{�L�]�0?�*����� n��ݻp�$	����U�{��4�j�>]k��Y&H����1�$]]/gq�zEP1�k�m!Ŝtr��ݻ�����|���bm�d�&���u�?�h.���U���F�B@pI,R�n��J��8�ޘ�o�ήޘ�gZ�F�P$ȇ��h.���u�ꤒ�o���`���ި��X�.�v�%�*���*�S��ߞ�^������R��S��ɀ}��&+�H%�$m8�vt��|�Z˭z��hu��
2,�����j�����X�K��2b�����u��9�44�jcǉ�$��N�h.������ʕW o���������n�[�n���ٟ�����wVߌy7^z��l7}�]�q�Z��Q7{��O�Ξ�;$��Ɉ��Iq4���7�x�I>���{��xϻ��IU$���x�^~.F�wa,m���y7^ ���zpl�ԓ�kٹ'�AU�؊����AU�����DT_�"����W�B*
��EU����X*@��
���  �B�*�* *�� *
���ET��@ �D *@`*U��B"� F� 
�EB� P��DE��X
�H
� X
�*�EH
�A`*@����A"*`*`*��*�AA��W��*
��APUz"���W�
���T_􂠪��W���*��AU��T_T_�����)���u��l�8( ���0���          
           =
�D*%P(P�P
(�� @R�  �P*@ (���     X   `eUP(	P C6
(}�Ov��k����{�gg��ɮ�"�2h^� :���o7�W�����8{�� ������c��1� �^{��v d  �� ��"����3eP�"݁���@  ����M�a��, ������8�����( x	��r�@齀�� pt��^��9�K�UE�v����@U ( U� ���=� 6� �� `�3A�9��H�@�hb `� @�l   3f��Ӎ�;( 3M D )  t@֔� *΀4�� J  
 a� PA@( PceP @  �
�wJ�w�w�9om+�Q14�n3J` )Y9r{����=�"��
)��o`�0u�cK� =g��Ę��&�ow� 8=@��EP���E �U,lT�c�3�Q7��n ��b�S-=��`�m�]�(�=%����  m\����M� L���C k�Ƌ ��Hr�X9��NMD�wR�   i�
��R�@ 4 �{���R� �d �~=U(h��hL�"{J��   �����R�  �M�R� 6S�O����?�i�����i�����{��� 
*���� QU�U?� QU��EW� �� S���������?Ѷb�!RN��C�I�GH@i�%�Jj�P��4D���H�O�cF�h!��-�C&c!�5�?o�f�bK�Y�4�(ƚeԸa$�RHH�dD�Fā�[5�N��D��D*������_��h�T"h�����6�4f|ʲ�K��aWfjă;�L�Z!�f�@�h1�֢���F�61�9�6�SՅ06C-܁1��.f��F�Y3r!�{�kSF;��Rf�MM���L��D�˜%��	���aщ�ʢ3G�^~����޻��0��X�@�D����?~�!'�Y� A#T���c�1 āB$a��c#�y�ɲ�RB�#��Z�q ��%�R�!MW���! ��H\޳������
W�H�|E-zN$��K���]f���[��m��
�)�!FM$J
1�B(!��WR�	��Ѱ�50�h"B��0�R�+n�f]$Zl
�biNɉ��ӆn���T�ҟ'�"Q�GKĪ8���ф�^HQ��B�I�$C�*JX�hĀ��m��B5��Ѕ.�˭��T�2���}϶�
B0#!��!P֍r�g�H�'��2M�@�,jD)
aB$�c5x}�f���� �X@�1�Ʋ��Z������4���X�Z��V֘�t@(i���D���8����}��־e4B "���$V&�}��Z�
D��0*��>�D�E�T4���?m 4l��6�x��)�� l�����HF��!3sqN?�0`B�p��s�g�$+�7�䌒�WLClx�(kp��u����*D�!!7XHGo5�0�H$w9����9�?�bos��#l�G��7y�?1hhɸ����t�n�WXϹ P8�F+%�Z�������8@6JI)��d#SA��)���b$I �`nN"��<4��8h��g� �X�6��U��"E0H%�H�F � ,�]i:�l?�?����c��D*&�$P #�A�?*EJ�q6!�\]��bAk���j@���a�|�O�]bkg��"44㳇��ц��?��:q۷�����)t���ߍ�%͘c��d��If�a����.�P�`O��ą�X�!B$*h�0ڲ�L��*F	�^��Ѩ[����$�+�/�B�n�$�����-�,
��
��X��f�e���rn��n_��Q�A�������1L# 6g~Ϸ2+������R�����5pX��b%���H=9HY��6�BJi06<I1�kX���ĉ���K�Y��ͻr����$���	I4S&�1�A��(}� �I�~��~�r�����v $b��4!F$ �HёBX��5�%�4�X�
b@R*`lٸ0���G�1a�����ߍ����3[8m�~4����������"���h����n�0Ĕ�fa�v��@�:�k�8M����k���SI#�.�1
�y���oؑ:X�,��~����"�]k�^R�� �n�����}Z0�������t�$�H'�~ؐ)�ٳ���0�Z2SX0֤0�a,`F�@�5 XӃ!i�#�B����IV�$1���L7Ga��%�eܜ�$)�ŌwM�"�х�$c�cB!ZkMI��V��0֯7�~�Y�H@�����^q�~ַ�6��f�s5�˚�Ӧ���&���DB������P�X1�l�JiX�!P�@06cF�kB-HR6�7)]e�ze4o��f��N�!���J���,�`h����BCXF2�h��J�u�=�4����~B�%T�aaB3�FVP��0���4Y�L�:�%s[	�@�*j-`�HWAo�[��WBD����f���I]�$֮CSJ�v+~x�*��uK3�<u�{N�_��p����E�BD�RF%�c�@��"!,�5�Sa����9��~O�'5��9�|%5�HB]�?k7�5�̟��Mf��74a�:���?d"�F-4a��BJi�� Ņ� VY�Mkf�6�K����!�
k]�'��`m�h��Z� �xJ���Ytļ#u.oV�"kC�?!��B@�A��+ �������n�X� L�~����	!�O��ī�~bB��E�bB�h��Yw��&����˛������k9��^M�s���[�u�
H���/8Ye���j�6;#2%M��7�ٲ2Pф7����7?k7x�߇�0�,�lW�(�����G��;t|t�3��˰☟"mH�BT!��6d��Ą����O��C�Bi�6P� �H���D���c�F^98m$��oe�L�71(�Z���E ;Hac��06�Lv,��ad©B;��JI���H쐉!(kS@�����F!F�7�rM��Y5�%��f��|F���q����I4L98�mٲ1�SN8��`M8ZKK�4`�X4t�)�ٿ����B����g��8���q��!����?$B��o7hi�b�!�I�� V�n~͘q�qv��H8�#�%pq۱0!�N8oq�l�Į��/	��٧����ۜ7(b�(C�!�"@��ٲ��4�) �6`q"SFÉ��٣�Ԍ#dю͒��L��M i�"P˸]����h��`mLaI �Ƹ�(�͡�;ջ>��ʒ�cl�u,u+-lH���1�@�cH0,�(0d% ��BB,ClB��~$��\7)�0�6�b&���_�5�g�i�6��2���m �5H�A��n����b @�
�@�1Z�F�W���l�%!e��m�@��#E��ҏ�E� ��
��%g
jSa@���B�j@`&�$^��!�&�a��ַ�H�b��pM0$����s�+�@ٴ�]�5�0�a�������%�3Fmv�F����m٩e�3�6R2+�c-���H	,�@b��_�K!��g9�$,
���a
,hŉ,� �B��C���"H$�e
��c�	��4�HA�d$,$u��nx8�xr\ٸ�Q�X��0ѨU)�i�����#ta�h�t��o"]`CFCa
i!]'E@d�_d:�?}��Z)������l���D�X'�#G���PИ�A�21/=���              �C�                                    � H                    � m�            ��z                            ��    �              ��� �-��m�.�& ]�I�o �  $�l��    �rukl�G  ���,�U�� +*���n ݶl��n��`   � �V��6�$-�$�f���Жk��a�5�m��*7��Ҭ�mUU�  [�m�m���Ԅ�UU*��*�+��U����zꥀ�2���V�
�%����[[j�5v�@v� �&�[׍��� �� �b��Q�9`:��Z��n祧��Fn��ڠ���P
��Uvp;5鼙���� 6�@ �`�I̵G+`[E�F�  ����=��  ���浛m,� �q�u�ܼ���`A2j��v��mPquUŐca]� 8ٕm'���ز��  iM�D$��jH�m��Y0[@dk��Z��:��v��.-:L�4R@ ��S�U����&��@ &5����m[&-���L��S�t Ġ�8�UK�*\둵-UR�P!��� �UUʷ�E����Hn�]��b���8$\�  ����P+�=s˘|��*�@pq'6�` Z���-��<��Q]�rU��[f�e����,m�	$tM��ow�rE��i�[�*E�`�fn9�y����%m�/[�e��jB�Kh$[Amm� l�T�y��G-�[��Sm�kYx-� -���8,�հ ��m�H�jn��ޝ=�v����i�� �c�-@@J�TU&����Du�sm�hݶ �H qm:Y[[��fk���I2������$��6I�m��V�U]�^�^v��$p��V{�V�%c�<�j�k�����n�L��r�m�b��^��%��WE�;Ut��Wn�F�M�a�t��ź�mm�ְ   wmɀ �M�Hw)j��6m�����`m��m� 6�.�& 'I -� 6� 6^�n3����8��              4X$� km� �n$[M��i+kl�ۛd�e��e6�` �4�$���V��]6b4�%+�6�v�ʯPq:��� $H]6�pc��m����Ih*m��pm���`�n�d�[-��l�nm&�m  m���ז�9�*˱��M��k����E�V� �u���:�v[�飞ذ�*�]V��輴�z���m���-�ڐ۶[[lź�nѴNe�@6؃qm�^�#&��p�`�ʂ��-����qs0����0 � $8�kW6٭�
ڸ�`  %�۫dmmu�@U��-Pv�������m���ܴH� �j�H��;&�x u���*�PUT��V���Mz�d8 nI,�am�p-�$m�/U�m�,����h$�t�-��*���mI�����	$�[ٶ�nE�8�㄀�r� ]J��]�l��ҭTq��ɀ  n��l  8-�qi�͆� 6�`ړ� �L����  ���mZk�n kXJ�ڪ�y�UeZ�J�hіӀ-�  H Ѷ� 	$�fճ�  ׬�&\�^� �-�p�m���  l      }���8�kh$�#ykp�         J��M��B�_y��    �D� 6�@$�T�y��  @�` l8���  6���[uU�pʅ��� ����#�l�     vض�� 8    �smͤ�^NN� �  �Z�(��20�ϝ�;�m���^���[A�zJ[\v�X5T���FH,�wNQ�n��,�� {e�    %�h$$��-�8-������d�     �6��`z�k̀      u]�]�U�"���UWR����2��+X�T�l6� �۴��^�s�:t�f�n T�U@U!K훡X��.�8  l8�:ͯ[��W\ Hڬ�� Hm�Z�횊�)g�`����s�`      �۴�l����n^��ݼ��>���L�    �`-� -�I  9m7m����j��ݤ��y�ӡ�.��|]}��T�k�r��! �kh� �  m�m@        6�-�  � �&kh  p[[l  ���$6�6ٲ�Z�"t�$�I�9m-��@ �7m�   s�  ���a!m�Ŵ�[D��[Wu,�  I�m�� �u���v�|�H[C�i�$8&�$ɶ��[m��$�@l����F���hkoi ڴ�6��2�u@R�\l.V��k$���bޤ��mm*�A\-U@.̭P��� ����ĒJ^�f���]R��U WUeq���    $ $ H6��d[��[����k�H[Bں�6�����ζ�e��   �m�m�%�  1\PBYu����k"�P
�3l����F�m&�UUU\9��0v� �.;s�U�һ��t���N�H����{�-�7Mڄ��`r����*�m� m�� m����WhͰ  $�� R��l��l�  ��:nӤ�b� 8*�i�m��`�6 ��i1�٥�6�$ 	�\%��d�[uJ��U@T+5��6�    �I&��Y/i��n�    ����}�o[%�[BF�V��u�rB� �Ûm�p   ��&�m �!�8�m����@4��  [�`    l�  m�M:��8�      6��� �L� 
���U�q��XV`� $��u�� �`�r\�g�� 6�6�F���/[m�*�YY[��j�F���ŶA�V���dX6�N��Y���a 	6[wL� m�m��έ� 9���Ͷm� -�ݲ۶8�f/[��kZ�  m�` �H6�B�ض�l�e�9h��  m�mm�����fZj�� ��  $�`�Ĝ�/��~�)V�A�ப��l��8$z��e����Cd7 �4�Ҳ��F�� m&�[I,T�\X�thVBj��t���jՊݴ��А�@֭�K.�k[e4���
Zڇ��+<��� �m���t��i��MvN���   	 kX
 �m��)i��^�����	6��� �%Z�����R{_ϯ��Ƴ\ 4Y�$H�H���@����*����],�v�0[*�W@�v뀶�A�������ֳm� ���  ;j�     [d   ��$��v  �  �۴�M�  pl ���Xm��ږ�v��  ��m��N��[A�m �@-�m[6�v�t��۱!�h �mm'l J m�m�3����:��C̛!�Z��-[.�v�1�u
KJ��     88]y[�[V']p   6�[qm6�a�N��6�nK����  ��d���I5�5�p   m� �����m�,�a��� ?�O���F��u�乖#sy��-�l�b3E���Q[4H��-�  l�hp m����p�� G׾��oV�h�6�m&         G@��7   � �  I 6���@$�k     � 	  m����   84ڂ@I�` � 9�� �      l   8  my� [E���i�l 5�t���jM�`���mؚ�V� �$  䉝`!m톝��U��g�'1d�u�<+r t�'FY"C��`���ֶ��2�H�m�N�� -m�7m�Ht ��l�\$Ze�lv� �k5 p�J�	����m����M�l���m�6��I�kk!�����`  nԴ	 m����`�� h �Vhu�-�Z@m*ѩ������T����W.ff��I��  *��D�D�U� ���|���(�
��D�(��C�� �+ �$X �(�� $1�+ -~U^< ��S ؉�� D@�^(�"#���������j�% �� ����U������R"��Q6
���"^
��`���| ~G� _�$�Y"u�"�����_�UC���@D���E�	c,�$Q�!�?.�zP�A@�����D8tv��Z" '�� � �B����4s�� ��#�E�� ��PB�XA��Q��P:��j,W@�`�UlQ�b� ,���Z"��$X��A��C E ���D�@�U.��%#6��/���@_ȁ�~�(tN� Ux���� A"D���  �Z��3330 6�      M��`  �@ ��    @  B�����&�v֝��,���2km����5Ս��g�gTH�,1x卂:�J���2�m��E� �Y-��z��K����Y��)#�����(j�LH�NGLs«�����Ŋ�>5;XMT� U<U��e%�I�n��M�RΈ�[C8�g&�9һ�-����ctck�Rt�F�]�p�/%�U����c-P:7jL� [�  ��I3MUnۖ\��b�x֎���Mq^MEl%ENv�م���BA)q1����u�2�9�s��T��Gs T�"�vG����P�M��VA㲩VV�ͩ���S[$������*���G*6R��6�4�Tm�m�9occ�j���i�R.{�����#3T�p�����̋I�=J��
���y[���W$#[URv|��b���mb�m�v���v��9��ke�L����J�r��t��;�/m��qm ��A��z��kY9B�Cmq������ۙ6�5%���gF��EI1��tP������2k'6��J&�T_]��LOH{\tv̭�&˫�;V�njT����q���3��uO���c:�KJ�R�!�6
j��4�*��/
�]�:���šn�zd޻tL����]ۭ��Xۼ�0��N���;�k-uX�g:k��J��pn;4M�Gd���Q;:��*�аy�,�J���n޻e8��3�ԭ��*�UR��F��:6k�R����ib'e8�5��=����ź��)< r�ĕ[K��<A���݋R�u����'6C/idm�� �n�M�Ha�hG���9�VU��ڍ% �i
���h�$	���3�G<=i�$Y|�KjUm�@Hk��UڮU��,ծSST�4]]a��*��`�D?�)��DO�6����矝�y>{���`�u��9WbW.�>��ɹz�-�`]��dV�t��6n�.	��v��4s����T�B�]��`���^�[<R��uH�ZL$�׆����#d�U\dN��֐,�=�i6	�ck��ce�:0#X�Yw,�rOa�X�d���y���׉����iN�y�D2+�Y�e���ܐT�zP׻�����{�V��Epa�vs�v�.ܛ���q�<`�v�dxݰ�`@�vX�<O�܏!˺���P�ӏ�?�B� k}x�ș��Ww2])�����s��DCP��Tk�� 7�^��@��Ԧ8��iH�Z�YM ��4/uz�Z.�c��)Rd�E!��f���@���C��3����[v88Dܒ<�)����ގ�����z����`?6�����s�L\���S��EQ�(�M94\`��ܱ8T��+��1)�oGV���S@=z���^�ʜ:�NdLDm4�qh�e5�`� DT��B�� M*BN"!dDBQ4���=>�X{t� �:�HƧ�lr!�h�Y�y{��-���?z�h�`��L��M��^�oGV���S@=z����%A<�$G���oGV��!D{^Y�z� ��]`��U2���sw%"<R9��֓��s��s�.a+q���X�QX'sg,3�S!Kl~���^�@��W�[�ՠr�f8I#�L���4׬�<����uh�e5fbG[v2'���%��������ۧ8Z�J!BB����g��S@:�4�i;�lq�����uh�e4׬�<����î4�D�F�I����S@=z���^�oGV��b�D?�m����X�;<�l�b����p���L�M�s"�Tbڟw���k�E9/K�2��}~����ގ������u��ʢ��Dln94/uz�Z�YM ��4�á���H�&�� ��9�?y�0��IL�z� ��]hx�z�dd��4�n-�������srO������P`+�H�P^��^׳[��z��a���.c�L���4׬�<����uh��DDDN�L�
��X*����zwJF��UN��$e'gVN_�����.�����m����1�$�~���F�������Q�@�}x ��f�ʨ�q�Ĥz�Z�YM ��4/uz+���aDm4�qh�e4׬�<����uh��R)18�n3�3��4��h�uh���=�E��UB���WWx�k��IGs������ �߻��i�~u�B,���P��0J���:�)��[pb�$4�Mh s;��l �aۧi����FE�[���ۨ��d������v��� �4䵩�1ɓ���;i%��\a�m���a=���u��rM�ۤ�v�'��gv�
��\����/	I�p�]PlJ[m���XX,���ԩ��<Tjݔ-�.renۇ��$N��ѣ���J�)a��q[ҝp��l����	#�/�ﾎ�ͶR�Ym�������1
��5ո�;:H�13�P�xܳ�ki��uH�\��UK�^�,r�e�a�I��������}���M ��?ff~A��Z^(ޥt]�uu3wUs�~nٟ(�Q2ϯ �ߖ�oGV��m��$�)2F���^�@�}V�oGV���M���I�"�ɠw>�@���@�l���K׬��+`�m�87$MŠ[�ՠ~�S@=z���>�~������y�ܽ��F�t��.���a�n=�0,�n�k�0��k�{3�#i�������f����ގ�������D7~����:�'�����v{�����c�h������,B��Q�����;�U�[�ՠ~�S@=z����&XM+��.�����脒S��p}���^�@�}V�ת��%22BGR7���M��現�OkoGV���IO���'L�ژ�$�t��J��U�V��l(qr�9�b3a-U�AI"�j) ��4��h�uh���:۱�)0$�<�)*� ݭs��$�L��� ���>�@?rJ�7c��qh�unI�뽻�J
/�
~P�:��f�k�W�;#�4��i8��-v� ��4]�@���@�<�E&'#c��h�Y�Z�Z�Z�ՠ{��$��R`�Ht	��WC���p�ȋ��h����m:�f���8�dln94]�@���@�ڴ׬�=Ň�T�"Dh�H�z:�]�@=z��j߽�w��~��~��t���R��o��z���ՠ[�ՠy[f8I$�Lq�8�>Ļ���>����-�Np&^[	(�
W��[u�73sI�"�ɠw>�@���@�l��z���`�T��ɎA��>������������w��2A�n��8i6n��\�WF�lq��"n/�}���~�S@=z���Z+���doM���v��%2ϯ n�N ��9�*云I�����Cp�^�@�}V�oGV���M�TX����#cqɠw>�@���@�l��z���r��*	�"4E$Z�Z������8���@����� l  �kb/.��#J��ݝ\�غ�y��ͷ%���t�N��$gf�v���jI�7H<�1���V6�y�������S�ώ��s���דW%r9�qςR�C���Q�C��kck<���;�%�חko�c�����*v�J1�n7*&�#]���c���4pB�Ygv�}8N�|��x�3�:v��3���;�w{��'���Ӈ�t��/]Yq'W�n�rӎm��hM����beÊ+<���V�R���������hϪ�-���<��$��E&8�R��hϪ�-���?[)�#��Z�I�$��wswWx�k���s��	$�{��Z�_��~䕹���䉸�z:�]�@=z��j�9^X�s#x��m8��-v�������_��>����-���-|6�ID' t��'l$�\���9(-����"��E�$&qd�[Ѻ5�S�Yͦ;R�$�?>=�j�-���-v��TX���j\��jkY���;�w�m�,�B&(�ۧ8t�����=�nbf�y$H�I�oGV�k�h�Y�Z�Z�^7��&HH�JF��-v� ��4]�@���@� �)ّ��$������������?��w]8t���P�{�
��WP��y����j���k�Ayʸ
�z$��skqjV+Y�MK�fk�.�L}I>����-���-v� ��4�$����8�ܑ7�oGV�����|��h}~��ՠr����F�5U5us�7M� {��M$�E�IB B(�~�6�UB�A�� Sʍ��tK4�a(���U�6&UMhNhD���U^�ڄ*�$f^��*$9n�<��> � ��H�@HA�!d�
FH��TlH���@�;~AE��4xT��:"�E��A����ʦ���PC���P}�k�� ',��s^�����^��L��Y���Mf��rqT~�}��{�����O{�]8~J"�uwN��RJ���f軣<��޳y�'��z�ʁl���z�qS=��8���(I~��%\):%J>�&�-�]�%�kkS�M��4���l���K�m��:
ŰIa�I����ww�믧 ��u�O��ׇD�uwN�='ʒшe�m��4��w����W�^T�n����� ~ۧ9�d���Ue]ʒE&8�Z�~��ՠ_tui�K��-���`I"y$QI4����� �78�"!z!B�_��T*���TM�}��'�֫a$b�$�MŠ_tuh�e4��4����.��K#� ㄪv(]�uq�W`,O[�R::n;La�9bA��X�s#x��m���;��@=�@�ڴ�Z\.�Ncq�ԋ@=�f�k�h�:�]�@��Yj6�d��4]�@{�Np]��?�7{�:)�_M�L�R����K������t������L��׀wWt��!��*�����컫�����В��� ��K�uww��b�˻���d���cm�`6�MUUR�իGi�
��ڞ����d��#�N�N4,�][:5��ī�H���v1y�0�Җ�N]��sɇA���X6��)�,՞K�����Y�^�̝���JCBMǧT�[l��v�"�J�9:�Z#N�.u'`2��ND�nܻ�>ΛJe�כ�=t���b<sbnI����x���v7m� 猂F�=�������v����m���cq�,[s�m٬�C@4�����l���c�HԒ)1������-v��GV�k�hmz�D�H�IRM�j�/tuh�V�{�� ��+a$b��&��/tuh�V�{���j�<�,vF9��DM�8��-v� ����ՠ^���*�u"s����ƤZ�[4]�@��ՠZ�Z�����<q-t*7�[��:�r������D�>��a4�Pe݇cq�JS�Z�m��M� �n���s�P�G�w��},�+�:nƋcl˻��C2���U�	�ȋ #2{���䓿��ܒE!�W�yAI�bm�i�M&`��8�k��np����x�R5$�Lq�8���4]�@���@�ڴ�\h�I�!�@�ڴz�4]�@?^�@=�%��o��]6��\v��')�]���η��z{W78.�aS��+@U�C3e�&��-��-v� �z��j�<�,vF9�<�m7!�Z�Z����ՠ[�a�U��D�71TUک�� ��� �785
�ZJ"�J?(Q3���0�np�S��;��FԌ�7&�k�h��h�V��^�@�U�Yq<� �DRE�[�,�9DDw_t��ϫ n����(~T&n���� ��v�Y�s:�=!f�Q=q95Էbw:^X��Z�rC@�ڴ��z�ՠ[�a�y[f8ԍI	&(�Z�z��j�-��-v����"$��D�����V�o]��k�h����$����8�ܑ7���p��� �/]`lDB�J!DZ�x������27���%&�ՠ~W��-v�������1�&���#n��^89���ݸIQ{qQ�h�Db�7�K��������ڴ�K��k�h��YdQ�ڑ����-v����Z�Z�z��c_�ˉ��"�-���Z�Z�z��j�/uxި���#q��0�-v��^�k�h���G�� ��8G��^�@�ڴ�K��k�h��d ` m�(�����:2�vf�[��ۗ�9�n�>���fZ���Jٹ��*��mN�R�u�5ѷ�H�.�6m��S����'3�Gm*����Egj� ��b�f�9��l�Fe�c�5M�ݠ����=�5��7-�#v	�n�d�h�`��ג�.��%7i�3�a�nv;�k�q�oe�+���G8������"=��}�����o�Gf�כ����'�t퐎�{rV�����Y9��:�+�n�@���j����n��}_}8�m� �ݳ��Pzz�������$pNH��@�t�gBJ���� ����7k\�����c��D��������s��K��W�����D7 ����Z� �m�`z)�y��H�]�Cj�i;x w>��sr� �%�_��x l��g��$Αb��6r��q���su�	<�!��:4k�W�=���Ӊ4Tn�w7(0 �2^����s�n�E�RX1���i�A�ɾ�r;5E��<x0������m����sr�=�<�@��Zhm�Mմ1�� �c�� �}��IEԌ =����@9q16Zwv�b�ݱ�x w>��.r��ɒ�@�ʪ��w��� �|�1��ۡ6ę�˜�`�d���9o ��� ߟ�c?��n^�U�uk	z�]h¾��a�v�0.莫S	x�����������:iQlI]��4 �L��~�-������F pt�7I2�i0I�����Uy� �ύ�����ɒ�@=�:�*644�ն�v� �}�\�#��*�yU�~W���2^�����؏,�Z�MX�lm��:��ݙ(0 �L��~�-����tT�:t7m&�m:F &K� �c�� �}�\�# ���'EX�
�$:E.��<����i[#�:��NC����թ0¬ٳZhm4ݍջm�� �c�� �}�\�# �%�r�bl����I:cv� �}��U$�\�# d�{��r� �$v���mЛbL� ��R0 �2^����s�n��mZm
���v7H�d�{��r� ϡ��+ʪ� ��P��F$)$d��ZU��%M"��G{>L�k?����_[���$˦���'{��r� U݊���F &K� �7i�V z6�d��1���gc�",v�"h�\���ss�f�luD�����s�n�r�) l�/t��[�}�G�T-S��h�6��\�#>��<�Đ{����_|���s�n�E�P��t�n�M�t� 6L��~�-�}筹|n�EԌ =]-KN�cM��[�۽��9o ��� ��R0����/~�~����&�N��lT��7o ��� ��R0 �2^�����{�W���%UWP%IT�B�B��*�"l��/��DЙ��Ut��K�$��kL���Ҏ���`D$$�$!$@�TC*��4:�ܤ���1�-VBؐ`ht�#����N�.��2b���A*B��`A L5�4-A ��� �(@dH1#�MB���!BF	`ԄRF2��`��+O@�W��b� 1�HЉ� �X��H-]G� �`у$X�X�4���F"H�� ���*@Q�p�� �#�>�"��`@"F,��a���?~�}          $��6ހ  6�`       @h  HSU��� 5U<���u��V���
���7@vP��vN'71mm�8��g�V�&h��8'وc�Z�M�c�cb��ӵ�Q�[n�,�fV�Y[��m�z�^���jѱr�n�Z��0��*�q�5��y%v�tl��ez�H���V�rkGNv����75�{�R�$��Rd��j��̲[qb���ޠ�������ɗk�k�� �m<��h ����8r�J����������<�����@#v{��і�@%�䦪��I�F$�$q"CN�҄d��<�����uu��JGK��7��}B�i�l['4KN��s*�:��9�Z�����\����6l�dp��-��E %鶲�m�MaxȲ��2�)��.�fh-�j���MSC��������mJ�R�fV㋶�hyH$�$u��x���o��G;ny	��ŮL��t�ܚ���[n�
Mͭ�q�A�ڧ�����ِm& lm%���
�4i��V�;�p"j[�ob�U+g(�l��2nƈ0[�
��[n�yઊG�\n���Wu
�, �W�TA��:%{U!]9�$¬\��p7f���Yra���%K�d6�&Cu�$�d��F6϶���6���8)��W)���l�4�7)�u��S�ˮ�d�Ҷg�=����]�vۢ��3]�,��=v&���wZ�r!�g�]���������݀-�Z�5��Tϒ�#A��0ãs��.N��v��cfU�����j�yj��b���Wv�#]7Ý��%Y2�]�I��-]묌�qd�)2�#lPJE����P�s���f^Wd���UUGn�إ��턲�$b���*�iV���p���[���b�Lu��\�����o�^N���]��<��Ҕ���n��JR�V� �(?� ��;��v���_(uO��>_ϰ  �`�x��=�I����[�k�����in{Y�	���k�ȵۗ�9b�6.�)M�v���홚�u���Y��VR<��Ÿ�K/I9b�s]Thm�{t�9�9�\J�(���(�}9�++�f�F9��q4�Iչ��:�c��a�B�ʹ�7e��gXR�c�a�n�d`��z[�}Gkqs���^��.��g�pq��u�H��x'��ȕv�r��}��k��>�ύ[�q�8u�q�2skH����5 �1=�x[bL���k �%���s�n�Y8�Bm%j�һ�X l�/t �8� ;�Ct�r�`Kct�.�V�����s�n����%��X {����{�uvTlhi�m�ـs�n�q�U� 6L�� {f �;�*��V4[��n�q�U� 6L�� {f ϡ��]25j�U��'�z���Y-<�ۙL���n���j���&\#qycF�L��������^��q� w>���Z���&�2b�)�}}[m�����O;��y���������<Ml �2^��x�"Q|�e�wm�*I��`#��s�k �%���8	�5V��M�&n�q�U� 6L�� {f�y甔�>7@,��M	���cJ�n�`�d�����[���7@9s�� $}��@�7^���v�\�Ș��������������؄,�z7F��Y�q��$�t��[���7@9s����Ԁ���� �We|���i�i��������F &K� �c�����)$�'�WŪtՍ�m��G�# �%��y�y�Vy�1ێ[��}��*J�Ln�E�I�0 �2^����s�n�<Q�-����v�n��ݶ��_.��}~��9V� �2^�#���3קgӮeڻ��u�� ��rb���5��m�D���A�#V�UY�آ������ɒ�@��8	�5v�v&ؓ7@/�* �%��3 ��� �qJ*�V��*�< 6L�� w8� ;�Ct�R�� ������N�V�����3 ��� �T�<��ʪ�%�tc���cCHm[m&� ;�Ct� &K� ;�f �n��]����u�b��{]�[����mz� 1�pW�]�7gt�b��S-S��h�Cl� �5�ɒ�@��s�n�C�i^P�ݶ�[bv� �2^���RH$3 	�� �[�������`�[�۽���`�����x l�/t%����m�RM�� ��� �5�ɒ�@��/���cUm�Bm�3t� &K� ;�f ϡ�[{����t���w��� m��
��_b9ؕ��&A�L�p=$枌u�Ͷ���vc[1���ۚ���	�F�幔s&�5���oc��m�����wQ�>�p/�:�k<l�"��L�6�Ր�<Q�at�\������r�Fsl�N��0k(U�H�q�
�L�]�t�ݿ������gj���5v�[���-��k���g�d�����&�]��G=��x��'wV���2l�D`yK�I��8�,qkv�GBG6N
�e�X�i�Z�:%s1��������������?W�^����|< >R˟[�եv7{�s�ϼ�<�ĐH����k���9yw}8uvTl�FԌ�7��Z/+f���M�Қ�5��ʇ�#h���@��l�?[)�{�S@�}V�~�.)�5�'&���M�Қs��V��p�V`I�4��&LyWga�v�`���j膹�PPљd�r�n���$�I�I!�{�S@�}V��jנ~�S@��uȢ�$�<nEv`��q��	L(�JG�6� �ݳ ��:!(�����n�7u%��]E�^k��M�Қs��X�ܑ��F�JG�~�S@�t��Z��%/n{� �d�����#��=�)�}��_��/5��@��S@/S`��<Q�� <s����c)�댼�׻*\����Iu ;F�Iv�5�FԌ�7����կ@��S@�t������eCɑ�4LRE�w�n��)�ϯ�[�0mk� ��Me�0�!#Q�q���h���g��ٍs}V�˕�@��T�	"�D��9Z��4�ՠw���}�����~��m�O���h�5P��[펮ՠw���]�@�t��{���v����n\���b��&�̸0��0r�ri��u�
��ɖ�j'�I3-�կ@��Z��4�ՠ�;&7lDQ�ґ�]�@�t���ڴ�V��ԑ�j##ch�-�ҚWj�=�ZWj�=�6�U;.�����B���� ��zpt��q
"!D/$�(J!���S�J�)Z�Su%����=�r� �M���ـk�� �IG��P�T��ݚ�ز�����5��7:��
]�ֱf�r�v�q��iƗs���j��(�~|�޲�Wj�=�Z����$RH)0�D��?z�h]�@�tUh]�@��j��D�'�Ȥ4]���v�����~�V�E
F�qD��=�Z��Z�YM�uzi�\�$N1F�ڋ@�]�@��)�r�@������?>o�   HM�m��&��7Lz������=v�=<h�'k��\豺9 �rI�	N�/�Ί �� �4�AL>�h�ͭ�!mf�X+m�:���4i.:X��\��l�*��K<�T0�TՎ,�֍��\�]a�����(����mL�K�.xǩ�����9��=�q�����Vx�M��7@�,�r��6ے�Fs����{�����3��0�sm]I�rP����%㱹S]o 7e�"ҋ��q�DYj��(�6&�"�/�S@��^����/��@�r���F�jFI��Wuz���@�v������j�*LSh�#�@�tUh�ՠ~���*�@?w	��0�!#QqE�_;V���S@�����U�w�O�E$���N-����Wuz�n\����%�=�3��u���v��]��T�Ӏ���c�n�QƔH�%�9�|�쮑�Ut���yh��m������wEV��Қ�YM ��l$Q��f��Yr�5�'��۽��*"�BBQF�x`ݶ`>n��i\�$N1F�ڋ@�v�����Wuz��o@�����(�6&
C@�����ֽ����z�����@YdQ�ۑ�F�r��@�>U��)�~���?[�T�"�)�t�8�hBN�e�F�s��ۜ���Z��N������,�y1LQ�d�=����z� ����
~�s�Հl�\��y!#Q�7�z����YM��z��o@�Z�=��
L���=��ٹ'��{�͛D�pX�KV]AO�jE���%6IT�D��� C��~	�j�dF,flP�Č��#��A���'��YH(X�E�-�F�
D!@i,��`�#' x`�
��
���8����L .�N�z�����V���i���*�i���qf���sZܓ������|�$N3���Ȥ4^���ʽץ4޲�y
�H��q8�q��ʽץ4޲�/_��﻽����߻���r�T�Z����gZ0��]�g������5c���I�'��cN7��ύ�v���zWkzTE��1FA�0R��Z/Z����^��?w(���N-��zWkz�Jh��h��*LSh�.��t�V����򈅑[%�@:�	��0�!#DD��ץ4�ڴ^��]���S)&{ʷrsѪ��n.�Mȵ��4���Z휳8���uڨ��& Jt�����Z/Z����^��;ϙd��b�4�7��ֽ���ץ4�ڴ���FD�H�q�]���)�~�ՠr��@?^n�"q���r7��b��h����9zנuv��UDZ8���h&��?:npI:������=߳�rM�� �t� �bH0"�b0*[�u������ɘ� �Ю��5�hdF�'6[tb��C�t�C�ṅ�����j$��D�1&ƒ��:􍝯]�ѽ�[:yKc������?[6�ivb����A�5�ˉ����e'�6 �éNK&ݪyR��7��<Fɵ����۷U�6�s]�8.�n�4��(�vkq��N�\X�z�+�b��B���YV�FB6u8쉻p&Gb-?�w{������~�X�.����JN�!�m`��`zi7;��GV][m5��B���7R�S��m�~~~���f��Қ��Z�5��ʇ��&H��*�vh�)�{�ՠr��@=r���0�!#D��@��M�v���z]���ԯ�BI& ����;V��ֽ��f��Қ�Yd#��$i�ln-��z]��ץ4yڴl�C��i��rN����\�>ݻ�����B�wc"��1C���s9�k(�h�)[G����z����;V��ֽ �y��B4�q�ܚ�Jl��}�У�D,ú�' ��u`wi� h��B���M
C@���@��^�Ws�@��MԱ���N-Ľk�U���=����ܴ�j�*LSh�#�@��٠z����;V��ֽ��ʩ�%21)�=t"�d�x]�R�'V�5H=��suk.Pn\cO �2"BF��7&��Қ��Z/Z�
���g�^lr)$�n��Zs�
����e4β�	�$i�ln-��Z����)��hTF~�S@=�� ��l$Q�9$R'$Z]������[4��h��ܓ$nbr9NM���޶hϪ�*��h�Th&' "��K��	�>������k\Cs�괛n x� 㘔�F�hR޶hϪ�*��h���:�c��FԌ�ӓ@�}V�W.�@�l��w����L�y1LQ�A��W.�@�l��w��s��(�2"BF��'&�ؽ�����hϪ�����Z�������5y��aWswv)0�4�l�;�U�^k��?[)�~W�ҹ$��I��%	0N��u��|��%�{@�lvI	sr\�Wd�7Y#OM94��h�����hz٠9
��(Ȝ�(&��/5�������@�}V�~���2F�"I$�4��?[)��f�����]^�W�8�%������v���Z溽���Z�,�(�#IŠw>�@��Y�[M���� ��E��GBJ/������ m� ��U����H�tt���#�GY,�v�x�3˹4b�V�nsV9�ح2�{v�{f��۷kv;տ���g�>Xݱ%h��7�Mp�b�m������\�v�Kӷ]heޝ�]�=*���X��Tn.���N|�q�V���:A��KF\!�z���gclj�%g�V�c��.l����A�݆y76�\�v�ih։�8+
<����c������%c.���{]��^�pp���]���.�v]�Wd�[���}����Ě�Q���������ՠw��@�ڴ֘�0�!#D��@�l�����#����-w�U�����;/���E$��5"�;��-�j�:���-v���:9	)#Ocqh}�ؾ�}��WuV �78�O��� <��=�ˬr)#PMŠuv��Z�Z��Z�ՠ��wbK����(9&!�lkF���]��&�V�h���{�e�X�k���6���f+}�?�����I��|�p��~�}]=XK$|Uթ��f���k2nI���n���(����w��8��u�6��D)�[�	U�]
26F��@����@��@��h���qr9)Z�WTeM��r�
u۞��������BJ{��p"��ɒ0��G�[e4�bI/og����=��� ��*�]���]î���P��hn��\k�h���K�7D�;8��_���v��ݽ��)�\��w��@�ڴs�ށm��;ϱ��H�Ix܊C@�ڷ����čt�� ��� ���:""�y9&{�����"�n-��7�[e4Y�����B�QI$�T(H��`w]`{N䐒4��9r7���g�b��ߍ�������
']���:zd;���3jK������v��
:���W~o@�����,x��ra�7��Rֹ�7)���&/v�����;Iuew�/~�IB����Ye�7E�wUg�;��ps�ށm��=�)�{��P�(��.��� ��ˬ���I$�Q���4���4
���?#���)�$$a$�����0�v�:!$��K}X�W�@��+ǣ�I ��N8h}���	O�������[.�%B���P(Q�\(�Nـk���v]ԗwsJ��n����D(Z��W�;z��?z�h�	*��0�bƟ�Ǌ%1I�<5�����y8kx�6^��Ln�T�nL�F�<Ƥ�A���|��/�����S���;ϫ'����{$���6��j�]���lϔG�(QTk��0����=����fbG���Ħ"6������ s����
g]>��;z��?n͢U:.��.����0>IDDOS}X�}U�y�Ł�$�w{8�=�����D̍��z��o@�빠{�S@���u�$��"$U 6Ā�H�&�Dbl�V�k�`jSU�>D�آ�4ȥ� ��PA����c)�"�A~%��B��dA�m���BO�]D@M����P$�Y	��="�?KKl-�a`T���!�)�BBK+a�h*1����,b)Tbj� �Ċ�$�FF#�� �2��Q� �Fo�]!#�E�"H��X��Jf�O�<����          [A��  �`       �-�  ����3m�����SiQl�$��X�1oT�u��׮�n8��e	�Umnz�HE�ً.���k�9|�m���������6��,r��c=�6XTbl�XB�nzvY�3��N�Rx�F٪�#�0>͵�1�*l)���v:��n�õ5����lq����]v��W ��V7f3�b"6��s\�k�8�vm�S�����!Ŗ�(���U���l[�4�`  �U�k�7&GJ���A��=t��u�f�.�n�'!B��m�=��mŧ#�Y�0�w�9m$�����8 �����ˤ����m���i-�ם�bư��� �RV���U�1���UW�V
'��(Rݹ\��,�zb����R�J�UӖ����r�U*�(&��� Z�����	ն�F�Hf�n��֦��Tw(6=*��G<k2�n�j7�-V�F�scj.���S$n����-�̐t,��Z�\sB)�v���UUR�R�1*Ի�6IJ�0[(h�*��sH�[�ѨU�3�gn��X��%��&�M�^��v�5�5QHĻpp��t �ΕJ�{���l�l�h@�ƃ*q�[j�kn�)��	�c�C�3Ⱥ ��UcQ��n���#SE��Փ�������Z)J�K�e��Y���2V6��y��L��+�˅��tb��*P��nf��C=5�WSq�MՎt��d�c�"OA���έ���m�(�h&�A(%e.����c�U��˶��6�WJ���R�J�Ա�qV�ujx^��3̡]��nz����Sn��1��ci�N��jq�S��7F�9wCL�P]N�m�ԇv��D�{1KC����e�56�:�!���-�B��T�fp���q�g����Kgn�H77e݅�Sl=%�9R�b��`��wkMe�t��@^ "/�6������	�D~�"�8#�Ϸ���������h 6ۭ��DhZ�滦�A��y^���5+C��.�Ol��)�S�v]ud)���Hj鴁��tvF��qv��u��v�n6�H1"/>kF��n�Fז�rrǶ��
�����-䀗��1�',��q��ƭ��YsJ�q�˰zv��ø��n�eC%�uu̷+�hxg�v�m���-#�XR�kV�r;�x�;@!M������ZRJ+(�ܲ��5��5�gpV��!�d]qt-ع��{��'��L���D����}���YMg��DD/���V �5ԫ
����I�'&h�e4^��׮����������$h�DۑHhw�=�ҵ�z���=�)�h�\Q��RF�ԏC���]n�ց�_�4z�h}��ʾ��}[�$���qȤ��׮��YM��z��kM��???q��<��F(����Ml��r�1� ݇�^�����D ����6����LDm��3�[���@��^���Z�=z�h�xv:ɍDF�27���o�B?�GJ� �js5�V ��`�lϔDBS'�pZ�.�7�4HǠ^?����sO�bV��U�|���1:
d�	Lq��?ؔ%;Ͽ,�|`>n�>R�����U��r)$�5&h�)�}���?�U�?����s@��IF3+0�ѝq�Ë1h�\^�1�^��=�
NN������F
+�CXlR{$��>od���}�{6��bX�'��l?�#�&�X�'���M�"X�%�}��5g��段�����W3[ND�,K����m9ı,O��p�r%�bX��}�iȖ%�bw_{��r�bX����0���ff�32浙��Kı>�}�iȖ%�bw���"X쨄50��Gn̉��������bX�'u�kٴ�Kı=��'�5te��ִkZ�iȖ%�5����iȖ%�b{]���ӑ,K�����ND�,K�w�6��bX�'ޘO���fkS0�fND�,K����ӑ,K�����ND�,K�w�6��bX�'{�p�r%�bX����j�\̹��ٻh�Ն�:�v�{F�5u�/NM�R*M	$sG��[ǳѫ�q&��~�7��bX���׳iȖ%�b}���ӑ,K��{�ND�,K����ӑ,K�������p�2fh�ff�6��bX�'��m9ı,N����Kı;���m9ı,N��kٴ�O�T5SQ,Ov[�5ɬ˙�.a$��6��bX�'���ND�,K����ӑ,KĿ��fӑ,K�����"X�%���~�k535ffeֵ�s&ӑ,K������Kı/�{ٴ�Kı>�}�iȖ%���H�qq�O{���ND�,K?��?FdY*K%?{���oq��K���m9ı,O��p�r%�bX��w��Kı;���m9ı,󿻼����ﮛ[�fM���f;��.�a^��2Ou��*�E'k3V꿞������ffffL����ı,N�{��ӑ,K��{�M�"X�%��}�kiȖ%�b_���iȖ%�b{^;tOjj�˅��hֵ�ӑ,K��{�M�!��MD�K�������bX�%����6��bX�'��m9ı,O�0�=��j噭Md�k&ӑ,K������Kı/�{ٴ�KlK�w�6��bX�'{��m9ı,O�N�g��Ma�ԙ�f�[ND�,K����ND�,K�w�6��bX�'{��m9ılN��{[ND�,K��{���ə�ffk3iȖ%�b}���ӑ,K��{�M�"X�%��}�kiȖ%�b_���iȖ%�bAoʣ}�fffffffL��  6�s��&�v׵���항��prlY��<��rQX`�zw�����ٜ�Q�i�r6�)])fM\����WY��Ӌ:�퇒�z�ۭ�m:S��Uj�]�����ۮ�m�//Sгkm��<�Vv[�X1�1��>�K+q��J��GnJպ#³���#��X���$�$�����{<��W��!ĕ�X��e�5e��H� Ƞs9,�5�r�;]�Rm�XbDx�e�rI��a���EƲ�k��Ԙ
�x^�l�U���}��7��bX���siȖ%�bw_{��r%�bX�����0�MD�,N�{����<�<�<�<�����`]�siȖ%�bw_{��rȄuQ,K����m9ı,N�{��ӑ,K��{�m9 �,K�ޚ�ֳY�Z�\��ɫ���"X�%�{�ͧ"X�%����ND��ű;��pIs�Ց ���UJ��d�����	$}�w�6��bX�'�{��r%�bX�������bX�'����ӑ,K���v���ї3Zѭk�"X�%����6��bX� w_{��r%�bX�k�{[ND�,K�w�6���{��7�����O�Fkn0��0�llq�"�n���Q/	"�4�.�HYk��Y��ѫ��r%�bX�������bX�'����ӑ,K������*��Q,K����ӑ,K���ɋ�7aV��.���!~!I
HRB���m9
��D�,O��p�r%�bX�}��m9ı,N��{[ND�,K��{�].fL�s5��r%�bX�{���Kı?}��m9ı,N��{[ND�,K�}�kiȖ%�bt�K�Mf\��s	.�Y6��bX6'ｿM�"X�%��w��ӑ,K��_w��r%�bX�����r%�b���~���I��n��{���oq��'���[ND�,K�}�kiȖ%�b{�o�iȖ%�b~����r%�b��~���C��R�9�%#�}}�Gn���Od�e�nS��蓞�Z��M&�$�Də��5s5��ı,N���ӑ,K���ߦӑ,K������Kı=����r%�bX����0���r�Z�5���"X�%�ｿM�!�
�D�K��o�m9ı,O�{���r%�bX�k��[ND�U5����=��G��J�[�w�{��7�������Kı=����r%��4���Cg"dM���ӑ,K������ӑ,K����٫��Y��ѫ�6��bX�'���[ND�,K�}�kiȖ%�b{�o�iȖ%��Q>��?�ӑ,K���?���3RfI��m9ı,O��}��"X�%�ｿM�"X�%���o�iȖ%�b{]ﵴ�Kı>�г�['�r��:AG��]�֧��tK�6N�v�(�M۪�a�9�I/Z]�]ήq�f����u�bX�����r%�bX����6��bX�'���[ND�,K�}�kiȖ%�bt�J{\�2�fK�Iu�ɴ�Kı?}��m9�:���'����m9ı,N���ӑ,K���ߧ����}�Os���~����S�5P��̛ND�,K�^�����bX�'����ӑ,K���ߦӑ,K������Kı/�����5�sY����5s5��K��>������bX�'���6��bX�'ｿM�"X�� �jnD����5��Kı/������6X7�w�����?w��Kİ}��m9ı,Ok�����bX�'����ӑ,K������ڀk�\3��	s#�3K���˸խ�X�͂��7R�e������z.4�ֵ�6��bX�'ｿM�"X�%��w��ӑ,K��_w��r%�bX�����r%�bX�w�l��W\�5��\ɴ�Kı=����r%�bX�k��[ND�,K�{~�ND�,K��ߦӑ?�j&�X���f��ᆰ�ԙ�f�[ND�,K�￵��Kı=����K䆢j'�����r%�bX�������Kı?}������d�ї3Y��"X��ｿM�"X�%���o�iȖ%�b{]ﵴ�K��ABj's���ӑ,K�����乗32\�K��M�"X�%���o�iȖ%�a�������ı,N���ӑ,K���ߦӑ,K����y�O'�wyӿ}����`�aUJ�s����n��vS<�v-;f�2��i����������"PR��t�m���홙CDp�6}M�a�jS=(2p�jt覵�q�lĹ"�u�-�u!�F�ʫ'*�4	[g��=:�۱J�a�u
�Y1�g��q�L�j��F���n�D�Yss�ٳeE!��Yc��w:خ�Œ�g���R�������]x�n��;Wa�۶�)^�{ ��f�a��Tb��b�\�S��kZ�e̟��,K��׽���"X�%���ﵴ�Kı=����Kı?}��m9ı,K�5}���\�j�f�M\�m9ı,O��}��!�+D�K�����ND�,K��o�m9ı,Ok�����bX�%���x�332ܹ��e����"X�%�ｿM�"X�%���o�iȖ%�b{]ﵴ�Kı>������bX�'��wE�����Y�֍kXm9ı,O�{~�ND�,K����ӑ,K��_w��r%�`�'��m9ı,O�0��&fYfkSF�d�r%�bX�������bX�'����ӑ,K�����"X�%���o�iȖ%�b}��g���5WMU��9�vܷp���y3Ʈ��t�����Wd�[����>׷��\�Nնk5��Kı>������bX�'��m9ı,O�{~��g蚉bX������Kı>�_jG�p�2fh�ˬͧ"X�%����NB�9I�1q5��{�M�"X�%��]ﵴ�Kı/��ٴ�Kı;���.e�̷3%�30�r%�bX�w���r%�bX�������b��b_���iȖ%�b}���ӑ�{��7���??Fu=5����7�ı;���m9ı,K���m9ı,O��p�r%�b
X�w������7���{���ܟ�4�E����,KĿ��fӑ,K�������~�bX�'}��M�"X�%��}�kiȖ%�b_�-�x����LԺ�kF�pSl��D[�P�F�&��0��X�g�y��{��8Ǿw���,O��p�r%�bX�w���r%�bX�������bX�%��{6��bX�'��wE�����Y�֍kXm9ı,O���m9� ����b{]���ӑ,KĿ{��6��bX�'��m9ı,N�a'|L�.��֦�\ɴ�Kı;���m9ı,K���m9Ƌ��BF�챑����B,Q) *��,��Rn�d����R� ��q$x��K5�M�!���0*o���2�K
JE�2��`K�RB3D���!2@�&�H@��5F�*1� !D%@ׅ\�x$ A�@� h��%])���+�@J�M�4;����D�F*���0�h�O�|!�E�pt���?�G������ ? ���O�����O����"X�%����M�"X�%����l�p�XfjL�3Y��"X��b_���iȖ%�b}���ӑ,K���ߦӑ,K������Kı?}������d�љ�Y�ND�,K�w�6��bX��0 ����O�,K�������"X�%�w�ͧ"X�%��]�֭�I��ՙ�3:%��I�@uv�q$ۦc0�E�]������]9��-���<�<�<�<�ϝߦӑ,K������Kı/��ٱ9ı,O��p�r%�b]�����ѝOMa�tV�����{��;���m9ı,K���m9ı,O��p�r%�bX�w���r*�c���~~���3*�DX)�����x�,O�ｭ�"X�%����ND�,K��~�ND�,K����ӑ,z�:�:�����������Sα,A[�w�6��bX�'���6��bX�'u����"X��P]�A熓v&��{[ND�,K��:S�TՓj���UV�����$-o~�ND�,K����ӑ,K������r%�bX�{���Kı?����������<�5�nŢ���l� �x�r�.����t��;N���www�����Eݩ��ꊩ�2�RB�����VB�Kı?k�����bX�'��m9ı,O���m9ı,O�N���a�̙�3Rf�[ND�,K���kiȨؖ%����ND�,K��~�ND�,K����ӑ,K���^�G���3Fk.�[ND�,K�w�6��bX�'���6��`�bX�������bX�'�w��ӑ,K���C�乗5�.fK&fa��K����{��iȖ%�b{]���ӑ,K������r%�`�X�{���KǍ�����ѝOMa�tV�����{��'u����"X�%�����������X�%���p�r%�bX�w�������������� 6ض���U�`��b��Ni{c�^�.�u;7%��&���qw;Zl�X�9i��:�i�Ó����Z����l�#=�qwb77!���I�ftl=0˪N;Of1��d�e���i�ۧqx��=m��\������.�8�����z���<������֑�u=����=c��M]�-q�2j��4���Ǟ��v�j�v{k���{�6�[y��خ܏[6��z�t�Nv��.����u�����=���}m�̫ک,���w���{������iȖ%�b}���ӑ,K�����"X�%��}�kiȖ%�b_{��d�6#7�w�����?~~�ND�,K���6��bX�'u����"X�%����ӑ?�P���w���������r6.t�+w����,K����ӑ,K������K�j&�}����r%�bX�����"X�%���{����,�jh��ND�,@������Kı?}���r%�bX�{���Kı?}�p�r%�bX���wg�̒�Lԗ	��m9ı,O�g}v��bX�
)���ND�,K��~�ND�,K����ӑ,K���zkW��Fis&)!��2����\z�/k8���k��0�6Ѹz��S�C{���oq��O��p�r%�bX�w���r%�bX�������bX�'��z�9ı,K�t��e̺�d��l��6��bX�'���6��PTx ���bw_{��r%�bX�}���r%�bX�{���r%�bX��_z�fS32��d�d�r%�bX�������bX�'��z�9�UlK�w~�ND�,K��~�ND�,K�ޓ٬�kZ�335r[���"X�%��s޻ND�,K�w~�ND�,K��~�ND�,QF������Kı/�w^ɫSX��������7���{������"X�%��G�����~�bX�'����m9ı,O����r%�bX���3�n�늸�ci�tn+!�[$�89��� n�ʎ��M8� i;/��Υֳ2�9ı,O���m9ı,Ok�����bX�'��z�@9ı,O}���r%�bX�za'}&fYfkSZ�̛ND�,K��}��"X�%��s޻ND�,K�g�v��bX�'���6��%�b}��w�\�5�f��5��r%�bX�w=��Kı=�{�iȖ? CQ5]��6��bX�'���[ND�,K��X]�K��3Ffe�]�"X�X��=��Kı>���Kı=����r%�`MD���v��bX�%����s.��.f[�s.ӑ,K���ߦӑ,K����kiȖ%�b}���ӑ,K����]�"X�%���������Vѝq6�)�F��G@uͷ`W']9���|�t�Q�w{�/�u=Y���k&�&��%�b����5��Kı>�{�iȖ%�b{���ӑ,K���ߦӑ,Kľ��{5��kZ&ff�Ks5��Kı>�{�i�)bX�'��z�9ı,O���m9ı,Ok������j��X���k�&�fk2\���fj�]�"X�%������ND�,K��~�ND�ı=����r%�bX�w=��Kı=��/��������������$)!I_g�,K����kiȖ%�b}���ӑ,K���AG�P������y��v��bX�'~�I��30��2�֮�&ӑ,K��{�m9ı,_����r%�bX��=��Kı?w���r%�bX�}���^d�..�]�&\7hف���ovc��xRΝ����#���}�b�Zv.������{��"}��ӑ,K����]�"X�%�w�͇���5ı?���m9ı,N�X]�Ip�2fh�̹�iȖ%�b{���ӑ,KĿ��fӑ,K��{�m9ı,O����r$(X$��t��MjˢkSZֱ7��y�^(@�'��
B��}8��bX�'��z�9ı,O}�ެ�z�e���7���{�������|��bX�'����9ı,O}���r%�b�w�ͧ"X�%�}�����{U%�_{���oq��������Kı=�{�iȖ%�b_��fӑ,K��{�m9ı,M(c�y'y�~���� 0  �۷e@��&�����y^�8ᢵѱϮ��]���pt�Qq8�$��a*�U�9�ƍ���f6a���u����h
�c���Y�<s�RӔ�On.w]��n���9���n.!T�|�k�뎢�6`������Ե�iNxB��A3ǋW,�u���bl�n/ �d��5u��$�fːmq��۲�ؕ��k]����5���Y:h� ��N{��*�a���x�f�}������f�F��3Y���,K��s޻ND�,K��{6��bX�'���[ND�,JB��Ր���$)!ur)�*j��3Zֳ2�9ı,K߽��r%�bX��{�m9ı,O���[ND�,K�g�v��%�bX����/����,ˣ5u���Kı=����r%�bX�k�����c��D�O�����r%�bX����ͧ"X�%��g��Is$���XL�kiȖ%��T5����m9ı,O�����r%�bX����r%�bX��{�m9ı,O�=aw�.fL�̺�kiȖ%�b{���ӑ,KĿ}�fӑ,K����kiȖ%�b}���m9ı.���������r԰�tA���v�mLv=�uk�eU��J�(G��w{�]��2��	���\˴�Kı/�{ٴ�Kı=����r%�bX�k�{[ND�,K�g�v��bX�'�����L�����kYs3iȖ%�b{]ﵴ�:5Q,N�涜�bX�'��z�9ı,K���m9ı,K���ꪑwj�l������$)!Iu����"X�%��޻ND��!���{����r%�bX�������Kĳο�7��*��M��<�<�?��`j'�w��v��bX�%���iȖ%�b{]ﵴ�Kı>�������{��7��������l\���r%�bX����r%�bXC����m?D�,K�������bX�'���6��bX�'�gf�}-і]k-��:����/g���ڡ��뒘ն�nr/Ll\붭��)��w�{��7�����{[ND�,K�}�kiȖ%�b}���iȖ%�b_���iȖ%�b~�u�<\�5�3R\&k5��Kı>������ؖ%����M�"X�%�~��ͧ"X�%��}�kiȖ%�b}���Ip�2fh�eֳ[ND�,K�w~�ND�,K����ND���"E��@9J"�"� 
?�t��(H(m�eC�?�$L��{��m9ı,Ok��kiȖ%�b_{�=�.e��3-��ɴ�Kı>�=��Kı;���m9ı,O�����"X�%����M�"X�%���﮳YsFfd�5�ə�iȖ%�bw_{��r%�bX(E�����ı,N�{�iȖ%�b}�{�iȖ%�b{��5�|kS.f�u&'T��B;wW�쯔Ps��
�rg[sC�AٺuG��+�n��O�����d�>������bX�'���6��bX�'�g�v��%�bX�������c�������T�T�ا�w�{��%����M�"X�%����]�"X�%��}�kiȖ%�b}���m9ı,Ok���M]I�I���d�r%�bX�}���r%�bX�������b X�'����ӑ,K���ߦӑ,K���	=�30��2�֮f]�"X�%�{���ND�,K�}�kiȖ%�b}���iȖ%��@��AM��]�"X�%���6x��k2f��&k3iȖ%�b}���m9ı,O���m9ı,O��z�9ı,K߽��r%�bX��agn�o��թP�B����v��:S��H<�v�hp���������S��[ND�,K�w~�ND�,K�޻ND�,K��{6�<�bX�'����ӑ,KĽ��|e̺��fe�fk&ӑ,K�����ӑ,KĽ��ͧ"X�%�������Kı>�w��E[ı=ܽ��k.h�f[�Y���v��bX�%���m9ı,O����r%�bX�{���r%�bX�����r%�bX�ݓ�׵��E�ar��ͧ"X�$D����Kı;���M�"X�%����]�"X�*�b^��fӑ,KĿ�|���+-r1�������ow�����ӑ,K�����ӑ,KĽ��ͧ"X�%��s��ND�,K�	$F�KG���&�2h"т��!�pS�F�b#��$cb��t#�k
��#��
 hJ%�&�shBI!	`�$!Ƅ!B���+F�!�Q#C\Ep�a�Z�`I�	� ��^w333333        ��   m��       @�����Cq�R\*�t��&�<S;v�`�U�FN�M�t��KJ$�,�IBMm����W]�3Ԝ]���Nֳ����ղ]^��\�\�k��)�lHD�-�rʉӪϳer�uz�v$���I u�M��5��iv�\qha��I+d&�}Q<�g���s���,[g��j�x�M���j��e�q�n6'\vӯ'[�u�ru�==Ӷ 5@r���E���WeV�|�s`  Xe�q���j��X:=��5���V�l�D��eL�;GU����eF�Þ6�d��$۳�v�$����<�uv�ui) �y�������n�6D&�&�2s�-��X��mUAԱ:�ʆ$��!���k�M:*�^8	�&�U�%��7I�*mm�Zt��a&�`m���^Y�I�:v�Yѓ"�wB5�T��e��H���r��P.��yۀa(- Y�kb����rfJ�P+<���{RnT��Y�xxL�ʆ�Z������c�k���S[y�kX`�q�c���`�=<���
�$�\��������N6���U���m��<���BngGu��a��C�+�(����a4]��q8���C@�.f\�I�l��5[++T���[jhت�>i��M��C�6V��Xn'q�d$�݂ۨ�Qw��ˋg�.� �r���v�If��:jw)Ξ�讣Tl��z̹P��]B��S��mv���,q�9�պ{��2E2N�p��I^�)ʰ&uk[R�J�UUJ:�n<)*�f�IP�M���s���X��̲�\�������d��v���R�꺐��+�&ڒU[$ꢗU��ᥗH ]�h���\��;f��\�s�[jU�e`*ڊF���P۲um�'-��k\�m�p�2�͎.�TFzxx�b�Bm09ێV��\���?�w ~J���&�O�E��� *G��S�GD�U	ݠUZ N����� �  l;#R=����6���=�ݸ^�z�4gΪf�vһ���4kMz*gV4��3۞ֹ�8�/�q���r��ɯa�zGi�"Uv$��i���Id�������WE(����Ǝ+�xs��N�(��0s�4�rt��t[Y��^��R�뀷&Kh�6.
���H��f�n�u[�����巀�8z��;�<�kT>����7j�i�r��\���6�97.�7�д�d!���	&rƕ�^�J5Υ�����Kı>�w�iȖ%�b^��fӑ,K����]��)?D�K�����6��bX�'��	=�&fY��ˣZ��v��bX�%���m9ı,O����r%�bX�{���r%�bX�����r�ؖ%����vx���d֤�&k3iȖ%�b}��ӑ,K���ߦӑ,K�����ӑ,KĽ��ͧ"X�%��g�.�32拙�̻ND�,K�w~�ND�,K�s޻ND�,K��{6��bX����s��ND�,K��'|e̺��fe�fk&ӑ,K�����ӑ,KĿ��fӑ,K����]�"X�%��{�M�"X�%�~?��C����Of�.��݇Gnٌ��^���k��Q�͆�Ʀt�n�6��w��to���3Y���k	��iȖ%�b_���iȖ%�b}��ӑ,K���ߦ��Q'蚉bX�{?��ӑ,KĿ{"?�!�B*�����{��7������<��>O�	���?D�=���6��bX�'��޻ND�,K�｛NAlKĿ�o�{&��ֲ�f��j�]�"X�%��{�M�"X�%��s޻ND�,K�｛ND�,K��v��bX�'u�=����a���d��M�"X�%��s޻ND�,K�｛ND�,K��v��bX����{�M�"X�%���w�ffj浖躹�v��bX�%��{6��bX�'��z�9ı,O���m9ı,O����r%�bX��s�����MLj���w=x�wۮ'���^�n\i��s�+�t-��=����������]�C_x�ı,N�?��ӑ,K���ߦӑ,K����]�"X�%�w�ͧ"X�%��g�7���f\�s3Z˴�Kı>�w��Kı>�{�iȖ%�b_���iȖ%�b}���ӑA�,K�݄���˫�&f[35�iȖ%�b}���ӑ,KĿ��fӑ,}��$��R$FHl4(~E٨���g޻ND�,K�}�M�"X�%��Ov��˚33%Ѭ�3.ӑ,K��_w��r%�bX�w=��Kı?}��m9İ?�@���o���9ı,K�������e���XkV\�kiȖ%�b}���ӑ,K������Kı>�{�iȖ%�b}���m9ı,K�ŷ���i�KU�q�S8����h�M�S�E�׵F]�����|A�?Yeb��������$)!H���~]wN����D(K��e���SSAv��˷��Z�����Z�YM�ff$w����#�<mI�˯�@�;V���S@�;V���D\R`��=��Z�YM��Z���wDr����X��WG)�j���M��\��e4s�h^��+��^��]���!R G�&���Z��W���CqvM��ss����\�-X� �Ss�z}��K�\�!~����|����$�Os	"�<����:y�`޾0�79�>J�����������W2M�� �����v�>JL�|�]~z��q�6�drG&�`r�og����u��(P�;���@�����qGL	��yڴ������<���v�:"!
 ���h�A�,", I@???~� m�l4�J��=@��1u�X�sm�K�!�9v�<=iղ�����'['h��
�v�o.��5?�_�Onؒ�������ɋ���ݶ�t�ܶKl@����I�׵�re4c<����rՃ�ɼ����wuZ�\�x�G'U	�56�oVʲ�q�e�hH׎+�l���f�#G������z�9l�h�=�j^v�=�{޺[��y�b��������o����{�)9۴��v��7�]*:B@ʹWmE���V�z� ������H=���:���g؜ �$9��z��ڴ�h�נ{���ɒE)q��ՠw��O�331*��=���L:�8�s�)�H��p�]����9%�����:Ms_8�#�'�9�qh�Y���������yڴ��e�0�Ju��y6���qv�4YEN*<Um����m�u�a�Kq¹�q�G"s#J)&��z���}M�В�_��׀�U�UM�L�fk0����~�{w ?�S�PP�y������<�W�r���s	0.����0�78�[�>Q
����@���hG�hI#��)��"�^�@�^��v���Z�����ҵWePJ�������"!'��?����h�Y�{֍�Q����)$hV���+nwO=y����sh�A5�֘K�0��ɒE)q���;�ՠ�٠y^�@/�:�8�s�M����7���В��%�P?��������j�*=���r$�G0�- ��x��)
_BQ�$��P�BȈ�����Ӏ7\� =�*j�Փuw5j�f���>��)��Հ=�:p�6�׬��+���$rI����
��h�Y�y^�@/Q���#��&!$��5����c{ ݇�㘤�f�ub{��{���Y���Wm+$�����- ��4+���
����$q��#RE��f�Ͽ�!B�6{��{�t��iB�������L��Lr�����|���Zyڴ׬�=�_苊d�"�H�]`rI|�D(�~>��}������*��X�E`D�`������R(��$Jd��@�6� <���z� �;�$��l �ܟ�ӵ�\��Z"��u!�=q��+�����Ͼ�>RF����ww�3���i�<�@�. �����<�W�w�*�;�ՠ�4�n̑(���������� <��rP�&C�O*���ؤ�I������@�;V�z�����Up�$pjb$nIs�o���=w�z^���DK�ç@��F�i�ڒ- ��4+���
��h�=k�$�I$UUU*�`�{%�n��b����z�	v`/<����,�c[��7k�";mB���xۋX��ƀӮn{7n��&]v-�v��iW�d,9NkO�|4�ݫu����ʲ�6&�O<� �����"3�U�j�lv�����ڹ:�<�<oc#[���!���<]�r!u�랞��8hg���*P�&�q�&J��d���'"��Z���n���l��Z�k�Iм��^�������y1u��]96��hD����	���z��s5�m��X��� �Ss���׀k\�菱L�!#����;�h�j�^�@�^�_a�`�Q��H��t\��np�]����J����`���-�ܝdP�D�I G�z�������Zyڴ�ᦝp��.�]�����z� �!B_%�>���W��- ��4��J���r)%.k=5������/u�Xl(u�森H���ڍ�H�I��w*�;�ՠ�f��z��\:�iO�2�3.w$���ۺ|�D�@���T9�z	���{9�ܓ���[��w*��$_����#R69!�- �}x��}M9�7����$��V��	Uuw��Q;\�����w��@=z�ݕ�ɒ<x�@�;�h�j�^�@=z�$����Wo���I�q�[�j�[�];mւ+���X��<+q7JN�P(���w5۾��nb�%2)�~����f�z��yܫ@��'Y#���$��=w�z� �SNp�79�S!�F�<��G1�E$���4�۹O�UO�§�@�Ba0^��h�U��@.�+�P�1� �D!b��Ċ@Ǜ!�+H��	u��jJ�)n��ҷ�n8���XF���HC
#�a	L@�"�!FR�YX4eH�\5��ZBN�!��b��u�������lK��U��������؈@N qL;�Q1ID&�5�~+չ8����f�����ɒI4�V��v� ��4>���K��M��̑Ɣ�HܑL�@�;V�z����h�r������~e?p�0�p78ɰ�6�{1<>/c���뒘��$�sY��d�������w7w?�7�^ y�}M9�I(_(�:���}$�SJ�&�U]]��Y�w�ʴ�h�Y�{���"�2BG�rh�r���Z}���_��w���gX)nb�%2����!B�{}Ӏϯ <��Q���nӜ��vi�wJ��Wv��� <���w�_��.�}M���6��Ȥ1(�bS$��4������=��r��\�v�����l��Z��L�l��BZf8����;���;��Zyڴ׬�ד�#�B�7	$�yܫ���- ��@=z��\:�j1�7$S"�;�ՠ�f�z��yܫ@�0�BF�l�BH�׬�wY�w�ʴ��Z����5eM�4��� =�� �P���˧�u�8���CQ/)Q�P�;�����   �j讝���e�6��6:��^�k��%�F.���-���(z�m���;+TlD�\����R�?���� ���tDt�6z��RH��4�L榡#Bv�d�on��\d�d8�c�T�h{{u�-I��0��\��]�*����[a��d�g:�!45t�;:4@�F=��^V3Ϋ{g���y�l`,q���zT�����T���d��n\�.d�iBԥ�׫[��t�t���H<�n�F��uEl���"b�2BG�rps�*�?s�h�Y��@/�ΰR(��$JdS"�?s�h�Y��@�;�h�.N�G��'�HG�z����4�V����@/vX6�Ȣ�s����4�V����@=z� �ܝ���Ȝ$�h�r��;V�z����4��A��q:N�%�\�2ۡ����f�z�z`�g\ܒg,H��ΦB�CQt}������^�@=�f��w*�:�2Б�f�3Y�&feܒ~�����,E!B(=�� ��Ӝ��s�{F�l%���c�M �u�yܫO�fb^�w��z�G�E�2d��8��;��Z�v� ��4��h��
E���L�dZ�v� ��4
�נw�ʴ
��dƣ&O��ݸ��%�F6ل��]��Ã���[1�st9��"Q8�G �I!Z��hu��7�Ӟ���u�8�β����͗V�����u�΄���G�˧ ���Z��h���H�8<�D�wX��s�=��
IzQ�(��i�h.��r��Y#�)���"��yڴ׬�*�^��w*�=��4�dr�E��f�W[X��s�y�s�tDB���I��]N5hj�.I�6�e�������={��:k`�`��зFƢ�Ű٘�k���??^��w*�=]�@=z�ݕ�ɒ<hr=��U�z�V�z��.����
E���L�dZ��h�Y�r�^��w*�:��:�G �I2G��w��U~���ӷrHD� A(�m������q`ۏ"�$s$��]k�>���I=�]?��]Ӏz� =���J�.k��=%$nt<T�g�B%���^������aw,N����2b��T����r��h�Y�Uֽ�\:�iLd��ȴWj�^�@�ֽ��U�{�3�H�Q��$�$Z���n��ID���ӀoWt��`��q&	�&�˭zyܫ@�v� ��4vTD\S&HH򤫺�7�Ӝ�z������6u�����w����  ���Z����n��^�Ě�m��f�V	�:�M�� �[s�6{k��$�QSќs�%�vþAX�F�I��6�f.�ۨ�c��ۻ4��;.,�:�v{ra��̊��t�U ;c���2B�Wt�$��u�B��;�v[�j{M��KZQ)]+�n���Sc.n^x�S�^yn�[��x���m���^���^���r�i� ��@t��Bo[�չ�.���tXs��n�mhuϭWd��Hm��o3��i����t�J����+��I������C׬�9u�@�;�hZ\�!�һ�wW8���
"dr�� {\�pWj��`�$jD�(��.���r��ڴ׬�ד�#Q�I�I��w*�=]�@=u�$�J]>��������U����)�h�ՠ�f�˭zyܫ@;�!��<Q�	2,J`�O�5�l1�Ix�q�ora#=��0�Tbt�#ڍյe�M�v��� <���������K�����:��`��8�L�M�Z�ر���ڴ׬�=�Q�qH<hr=��U�z�V�g�BJd�}x��X ���ɲ���\ڹ�s���;��8����n��V�ծj�B�'�L�Š�f�˭zyܫ@�v� ��%J����C�%��G�Mv�-����q���#r]p�y�������#��fy���6�'���4�V��v����\ �yXH��lRF�$�@��a ���8�[� ��y�
&G=,���h.�ꦕ� ��� <��
��D)�m8�����nIϵ�۹'�h�BA�5����@=z� ��0�4�����8��H�	�usbhN94׬�;��Zyڴ׬�=�F֊!�1L�h�
H�"�T=x�n7K�Ʌ��	�:���k��0�6���\V�x�@�;�h�j�^�@=z� ��:�A�LRD�E2-�M�tB�2ϯ 7�^�����3��p�r	�$qh�Y��f��w*�;�ՠ��Ơ��ġ.��9$�L�>��r��7���|���Q���_^ {��+�*�ꉺ��9$�;��Zyڴ׬�^�@/Q��9�2B@x��m�&!���Y}�	*��v,C^���KyJ�L�Ι�*�������� <�� y뿢"!~���ϖ�~hϾ	�Rb�- ��4׬�;��ZyڴsW0T��0N94׬�;��Z}����e�wN o>�ڜ�Zjn�v]R�Qɠw�ʴ�h�Y��f�_a�`��&)"S"�����@=y� {u������%$�P���)�RU� E�a%ѥ
6�+*B�B�Z�$! F1A15EB4$�	��R���T��h�e!H�! bRT�	 U� �h(J����"!��E`�a�Z��R�RT�L7��ţ��`�����H$ ���¼"]$�Bf�g��pF<XR	@�P�T"�v!�iH�;I j�H��_��	T��k/k>����      ?�� -�m��  ��        H�  i�����v��Ϋ�L�����a�\���㴷m�:��DL����闍��1qlh���e�(���\��c�[pW]��ό���鲜�� �������9��7 ��\�m����*�% ���eʘ�l����vu3ҥ�8vt�'4]u�X#�uҭOU�.��m�n�q�ۜ�wU���A��F�	�;�L���[h��E��qJ��1�rJ��  i:�nӦ́�j�wi:�LK���4f�x(��Su��Z��U���I9�`���x��[=FteJ:�^�m�&�u��Ͷ�֙[W*�t��c��4�M-4�j�ʏe��*nm�j�.+Eh	{8e�pC���ӯ%uf�i/^�!*�_}����T�/j��T���lv���j�B35U��f��<X�F�2[��ک]���,�\�Ā�%�od����'Y]�KwJe]�l��^� \�$O\$:�JI'���[F��j�
��kY�_fA�[yY�F��q�
,��m�d�U���+r4;'eN��ft�4�P�7]pMU1�W���5b[$r��q��s��f��Ō�;�+u�a��,l9t��9�@ ���P��rm�`j�GUU!��!Ҽ����lMU�Y��]��̦1�u����T�$��*��1]^�F�"p���k�%�i�Mt��rJ:�ud�+u�f�"n��j�l�p,�sMI<b�٫mѴΈ�I�E�q��=�]�e���ԵJ��T��pn�F�ƙ�qmWKP�*�"���]�r\Zö�8�T��&��5m/-\�:0�M�lv� �ꙥ�n�^[� �uu�@�l�3l���e�Z����+�@T��U���s���jI�n.N���g�nB-��H��B-�y�ݳ帛(���̹�j�.(�< 8��@6@z�&DDҠp~p�"AMU�(SH�>��o3333 h 6��*��i��v��H�b�j����ݬ�m���{i�4�H����er�Nְt1�6�t�0[�	��[g����\�knq��u�c=11�g�8C��,u1nt+ *�F�[�ʮM��&���Iq5萌�6*�{Q��[vL-��n866n67Lvڍ�Q�����T���ø*&a�gB�klܒ�n�C���{���w���;��FY�`B�Z:�9�u!v�δi�P�.���}o��	V�����󟏺me�=T��� }�׀�w�o��8�� /u��A�I��G&�{�������
d{\�p:� ��y�ДEPor쑍�أ���&����-�;V�(ID)�y���׀l��t]ժ�H��2)�h�ڴ׬�wY�����W����/��� �(���E�z� �S����r��?m78���]��л-�k�����n4;i��&7+gFM��.����wb�zb	�&�{����U�~�j�^�@�NH-�݅�wJ�]]��i�tD~��,Q�DGУ���}�p��^ {u�|�D(�;P�a6U�tU��ڹ�s�z��Z��h���;��ZG�\��*�ɥwv�����"���^ >� �;�h�ڴ�X88�`Ԙ(�rh���;��Z�v� ��4�ώ�[�L���3���7Q���x������tsb��u��I�җZ�겒�e��&��w*�?s�h�Y�g�[��*���$s��ۓ"�����@/u���4�r���Z	���ݗr]���w��w�J��!"�H(a>P���t�ܓ�k������	�ur\�U�]�}	%�}�^�Ӏ~�np��<Ӓ`�L������V����@/u���4^�Y���F��q.�h�-ũ�{n�L6Nn�IգJ�Y��d(W?��wE�F8�S"��=_�- ��h���/�ʴ
�r� ܂y$�]\��w�%
"d5����t���Z{�N0jLN94��h�Ӝ>Jgλ� 9�� ��T�ݕSuD�]U�ww��(���]8�wN =�xBX�!@��8I+TSyx�|�d�cSrdS"�?s�h������O�o�@�w*�;φ�I�!I��&�,�"4�>)-T�ܹ�H�݉&�qdڋ#L�		w5bE�I>~~|{ ��4�r���Z���*	�w%�]�� y��D$�N��Ӏy�t��w�(�7�I�M�We�*Uuw�v�.���s��(Q2s}x����3��L�qĦE2-�;V�^�4��h��Z^\\�E��*Wwh����� ��}��]8�����$�w��y����π ��UU!6�ۗ��Ύ+Gm�����w�9�$<�z۴61<#�WJ�]�v#��v'�����'�i�]����,p�s	�P�E��l@-�(���&���M2��J�No��\j*��r�;:�݃u��U�cج9�ͣ��k5�GK�9;OlH�I����g�E!�Lo7FiT�K�;6f䘽��=�lA,�v�H���l���\���
�%D۹�[�Rh̷2G<]_�d�����ƭ�^S�Kѧ������j�&��bd˚MN�s$�����_;�h�ڴ�Y��+����q��$��V���W��@>���@��qG2)���"�����@/u���4�r���Z	�j9	$Z+k�wY�uw*�����uى|	�q0�����:��h�ڴVנU��;~pD&nI�fV��O��1��\vF3˩�Z7#d9���w�l]ujyc�@��U�w��@�mz��hhZ�*�*��m\ڹ�7����DD%P��Rt��Հ���tӜϧG�ȱ��I8�Vנ�f��ܫ@�;V�^��0�#�r��w�^ ��t��np��`��`�m�8�h�M��V��v�����Y�u|6��ɒDb�V�v�.i���2��>M�nA�MI�ӮY3�$z�6�d�cSrdS"�;�ՠr�� y뿾�Pw���p���|\��+��BLRE�r�� ��4��Zyڴp�bYq<�"&�= ��6I�uӷs���! B��6�U
�I%�IW��t�w]`�N�%�ڵv]Ҫ������]8��e��׬�=pκ(8��JdS"�;�ՠr�� ��4��Z�xP���u��ٰj�b�m�	��=���9�m)m�de��d�o�_o��b�Ļ�#���呂z��Wr���Z{�RH�L�$���h]ʴ�h[f�~�\v���Ɖ$�:��h�j��H�}����4][���)���29�h�j�m� y�
X$�B`
����yӷrN�E��˖��)!)"����Z���Z�78�(���
�)L�Wv\�#{=��N�j�
�9���,�T =��'`m���Ĵ��#CRI�>_��@��U�z�V�u�h�j�
�p$#x7#�:��h�ՠ���Z��g]��L�dZ��hsw�D˗�X�r��6\��ՖU]��G0�- �h�נz��h�ՠ����$�	2H��h�נy�Np:npu��5|�G(�J�AV@dg�=�o�fffff � ����v�GD8��w+�;M���Mò�����yw�h.wF����JX�CAoF�R)g���[Grڥܸ�^�؛��Rt`��pN,Ok�Z^�ٲk�����i1���.�v��&�Lk�:�)�ݺ����tll+ul����]L�1�rB�3�������Ϭ�DO���c}�=lv���܅ּ�A^/�����u?�.k��&�E�y�x���"����/�ؼ\0��'Y��+��MU�����Šw��@;����h]]�H��Fܙȴ�o�Ă߾����:i�}	%2>�'qvUIaw�I�[��@=z��ܫ@�;V��j�
�pq�hi�4׬�<�8����$�����5�� �	�j캥Uuw�k���BJ���ﾚ��h+�Jȣ9��QW�G8x�;[��=nk��Q�)u�,��rƺ��\��L��ƦE2/�r�@wt�w8��r�;�t� ��y���˹$���ohA����	BWa���M9�7���DBP�Nw��5��H��h}~�Wr���Z�٠��:��lQ��D�h]ʴ�h[f�z��.��H��Fӊ)�h�j�>IBQ/������5�Np�$������O�z����^89���g�����8��TbB6�I�D	���rQ���l�^�@��U�w��@�5sA8565$���h]ʴ�np[w�
(�5�� �	�j캥Uuw�>�]8���6�RH�SʂkA� �Bs_Eڑ��%T��$U��z���E���, ��Ak J�@�(@!��(H��
����B��!+sW�@`%b����R8 A���:B]M:����	�*'~�9�F)�H��a�\؎$��b\٠��8��B#�
�� 	>�"�B$; J��4�T��FAv)�� �#"HȒX� R$H0`@� �]@�6��DF��T(���삧���T��;`�
����D0���b�G��(�D8��~��rC׬�=p������jdS"��g��IK�� }�x��tӜ���Aȑ$#�#�@:�4��f-����˧ �Ss��L���-]ے�\0:���)G�'s��p����K���nt��Z��7��I>�~|���s�o���~�9�� �ʺ�j6(�q�I4�r���Z{��^��ٙ������#q�c#i�ȴ�^�4׬�/�ʴ��D��	!�h�@=z���������
H� (
���'ʂ~w_���I�j���Y2蹪&���]�(��˧�k�p�Y�{�EY���FH4$�措kO^����}9�1�Z�g��H N��	sn'{(	���7��V��v� ��h�Y�w�������jdS"�7���(Q2�^ o>���s�Dg�$|���9�BL��#�@>���f�|�U�w��@�n���E#ȞHӎM ��4�r���Z
_B����� ߉�W�UM�uuWBR=�ܫ@�v� ��h�נy�y������  6���:�f�p��B�j׋��@��[r^s�u�Z��\��5�鍨{�۪.����ǆ����ώ���t&Tm���m��W��Thm��\6�z�qՉ���>X݉��ϫ1���<����z�Z^;����s]��,$Ѭ��M\e�1A�%C6x�m��L�
�V�0h#:ػKЅ�5�����;cX��ݧ���}c?�ܼݫ����X^��ˬ�>�It{���Z����Չ�mHΖqs�E2-������Y�r�^�|�U�{��H�MDAɍH��Y����*�|����-�ڴsW0Wp��6)�.����Z��h�@�c���d�o�z�g �� �J]>�����X���jdS"�=]�@/u�.����Z�PIO���'1&�6�$���z��8�W/\��뮛
c�LC���}�@H� �AȔRd����~�.����Z��h���Q(�y�sY��}~�u�#�U:":����}�̺���7��p��̖��ڍ�8�bR=�ܫ@�v� ��h�נUy:�m�SN(�E�z�V�^�4]k�/�ʴp��"H91��^�4�����s�>Z��h��j���s��м���N'k�n�]��n�ᵣ��.4%'#��N6�`�$�A�lr94]k�/�ʴWj��f��Ʈ`�'�$#x7#�/�ʴWj�^�@�ֽ��#�h����jdS"�;���rI��w70]mUp43>�w��?s�@�����J)	2G��^�@=z���U�{�S@�n��E#ȞHԎM��^�����|���|h�Y�[f�A�����jڳ���ܚ��6Gi��u�^��e��F�җW1�Q�G�JG�w�ʴ޲���h^��W��&��Fӊ)�h�e4׬�<����r���#���E"$�n�_����@�;�h�e4sW0W�Bln94/uzyܫ@��)�����P�: :Ef�A�
�w��@�����d�o�zyܫ@�D/�k��ǀ����k�ۤ�i�8{H\�`��
���mԮ�!ͱ�-諜4��8�(�kVl�N�K�ȴ޲���h^���V�˕��ȔRd�E!��f���@�;�h�e7�䏯�jppQH�'�u7uw�l���7�Ӝ>JϷ�� ��@:��`ڍ�8�bR=��U�~���^�C��ϯ�@���r	�#i�L�@��)���}o��:���i��%
×��������X
���W�۴�N�\���Uj@mk�������|�,��	hm�'(:�W+�h�R��r��s/<^��CX[m�:������k�8�x���e��x���V������m�h�켃�NV�<*mE;F�\�/k�=�Y#V�ۡ,/���9tm�ێ�}��ç9����e��u�j,��f�|s�Z�0���j2[�sԦ������->O&�G��k�I�dц��wH;a��Ș������#�ޱ]����;i��%���t��R�	�*�`����k���s���=�|`Z�0_`�L�hr94/uz�4� ��l���?�'�T����V�˪EU�`�˧ ��l�脦No� ���w�+Ԧ8��jdS"�?z�h�@��W�_;�h�Z��E!&H�R{��?�������?��~���?[Ҹ�JHd���|����m��,���)�ԛ�J�l���g��vk%
9�"y#N9?˯�@�m9�?y�?�	~�9�� }=%u�SuR�Z�Ks5�'k�n� ���$E,	$B��B*��P��c�`�w�z}��,қ�9��&E�~����f��3�.]~z��ϖ��u"�8�D7 ��h^���r������j�.'���M��^�|�U�~����f���VĢ�F�Nř[���ۣNB� ��گk&�m��0�$�B�œ��4�]�T����mr��?z�h�@��W�[�Ԧ522G�L�@��)�����^�|�U�r�jpr%��#QHh���䟯ﻭϑb��	�(An*@x"&� �A�\���'}���@�k֢p�9#y#N94/ux�4� ��l��"g����S5�SQ�G�JG�_;�h�e4�Y�y{��/���""�dx�0XbJ�a2�ۙ[�����J�郪�b�\�����# �Ɯ�x��c�"��������^�|�U�{��H�O#2K*�J�0�Ϣ&M�}Xmr��?z�h�`��1F�#�@��W�?SNp�
&}�|`7׀~�+R�a4�]�t���:QDDDW�>_N������c�P��P�G(Id����ޥ1�FH�R)�h�e4�Y�y{��/�ʴ
��d$jc��ٰj���%��nv�[5�U�(h�X��̚魥ɋL��=�O���/ ��]`�Ӟ�D(J=A����;���c��i��qɠy{���g�$}�˧ ���u�rJ!)�}�3]eR��8�bR=�g�@��)�����^�U8uƜ��"6��ȴ>J!B�og����k��)|�t�����O���Cp�^�@\���xꞛ?m�?䈈�
""?� QU�� U� Uh ���@����
*���
*����X@T$P$P�B1B �T  �T"(T"�B"�B 0�EBP�		dBD	P�DX��,B�T "@T"��T �DX��B"�EB"�P� @T "�` �T �P��B �B ,Q(,B�P�
Eb���B
#E��B#P��`1�P��aP��E��T"Q"�DX��T �A`(@T �`�E�1�`+P�)E�#P�+E�"E`�$B" �`(�
�Q"�E�*@T" E`�E�	 �������� ����
*� Uh ��� QU��EW��_�@U� QU��EW��_�����(+$�k&�2z`��0
 ?��d��-��PS�@�      t      �`  �@ ���@A���T � * 
)@  � ��( ) U*�P%E(��U( Q`   cT�
 

 Q2 ���ͽ��x�w�/&��yw�7��
���O-��W�}��w_������@toJ�n�m�ξ 
��qqQ� 
�J�x]���֜����M)�P������w6���[���7�]� υ  �h '���.m������x���}nR�= }>��[��u:��j�ê�J�ڪY�޷�b���ŪvruO�� �^z}<�].,�n,���g*��E
�=�^�z5�N^�^���^� ��(�P  ( �G�}���w�={��������:�w�P}o}>��RŸ���+qgU{��y\w}j�=�x Z�Z�o{���^ N������:�w:�w۽��wͩ=p �ܼ���ms�{ϛ����}}��^�Ԡ�
 P("`�il����w�W��r�}<�()e��>� ��t�� q �� lҜ 0 � �)@ R�� DҀ4J � 4�`t�w0t�  v��ng@�� � �q �@�P ��Z �ܥ qAF �����}�� >����sn�ۛ�d�Y�\�w�o= >�z�n;���^  n�7t��^��n��d��so�/x�y=�ܯ'.^���+���iqomOx������ϩ��z���  ����T�F�  ��jf�J� �@�=U*L��  '�U$�UA���ha������� 4�M�)$&@4<SR��Q�������������Tn�P�|��!% ��3/�\AES��
��T_�Ub��*��O�g�#Y�BH�3��Y	$u����7�xђ�������$C�H)�~��!��R05lI"�T�F��Υ�[��.I�(�	�i�l�����������J$�4�H�H�X�$R
���|���a��q���8�9$I"��b��"��I-��ֵhZ�����
������d �~�	�&���l�Ԁ$c�.a�҉�k_�g?}�~��m�9��~̘:bBjw�g���]?F�9qb*�c$��ɬ���
o��
����@�H����
��H��S�s|�|�I�j�J^u��]X��\|�ݷ�o�l�P�K ���?~0"@�B�B1� ��	#F����D�t�m �CN;�0a$�1�ٲ�#M8�v�0)�6�`�Rfݦ'�F(D�#H��rٙb�J���_w�=���W�㓫�c�ԺxNᳮ��|�8L,�a	��&�䛚?�p������W�r����0��0��K!���3�q8$CZ�l��l�aHP4�f�# �ӎ���P�I]�9�n?F���������tI%�n.1)���I&�Q+�pHA�(�U.6����-	\6Cz���v����,�r�R��f��+d��a5�H@�I7i��&�O�'��R��A
a�ы��H@l"%� X�@#B,��b����"u	!J\�d�@�t̔�$���jJ��a �S2��"�)$$ Ie���I��p�� �$��V[���6��$$!�d%�Q4�҃ E�¼zB*��r��vA�8��2BHF4��3rK!��ؐŃ��[u9ˣn�H�1����SHB�n��𳟿?�F�5��шka�Z#)i�?}��5?]���iă]�������6�:D�ֲ�������}�������cX`Q��f���G�O�220�X1cf�փL$��CC��	k��H�5�Ó�H��7��޹9��-�s��ѷ��%�������؄i����}w�R��N-�XaB#H�R�R:H��O�B�����8N0�!�2�	���!�(EEl�`�F$ h�x����T����Yђ�hCh�
C�(B��bƚ'�P"B:`m�+���	��X艁��"Zh1��q9���A6��)���7&�C��MD�I��ĉ��G�F���$lL���!a	Np9�)@�����qێ͘~�l��:��&9��l8�BkSh���i����0�6�y�5�a�d�ЅH�2M�rH�p8M�ȗD�$��pX�8Gp���#0L7ŃRH��$�!ty&��#yd6��<p?(�aCI+���!a?~�NkY�9��A$-B���"�?�cM�C�$(CDL6�He� NI
�B��,)�������d#];���Lk	`U��E�So*��7/
JD���
P��ۖ�C�[#5l��.��i�
���ėU֌b�@������ª�~���	J�*�a�D�D��E��Bƒ�aB��
� �� ���X�V�d�$+�H�8qՔ4��I�
�N!)�9ux|÷���� �*� v��� �]�ߏ�J�q���a�B���~�陁�k˼8��
��4�vƂE�h0��]�%y�U4�l^	��F�0�͘h�����ӆݘs����������]�ɦ!Mԅ��M8K�,�а����CP��b��
B����l���!t~Iteܘh��o!�g?�*B�M�
J�H@������l#M8��`c�V�bm�4aCd#�ƢhR%4��E����āMaw1��)��0H�HЍCK���	
iX]No_�q��s3�f���oY�S���!$#R��`F��V4Ѥ�D4���؜!SH`���~HsG��/�Hj~����7v1)��s3$��8_�
�����VB,u
i�T�E "Ađ"$v�BE((V!Z2ۛ�,?�aͤ�?$HP�D��1�$)(D��D4aϹ�M�~!������?3T�%���9����j%`@4���H���&w_�x~9��i�B��X����BP���8�]�X�)�w0�T���xp!!�(i�;!ͤ*J2聁f��ld�9��lvm����� s�ȅtMË�	u��!XY�p��rnht+ #��B3�M���Gd?<bR�5,���5
&� 8Gd	���iJB�u�������#�
�H��"�1ѦcA �tHq�e*���֡��"ɣF��%4i���Rt��	@Ө�5�.~�Ѩ�.�z��ф�hHj�@�@#4M]0��޻���ѣZ��K;�r� ������������фXФ+I�	YuYR�
X|�G<挚�0(�Y0�Y�X0t�����G��#]&!�"P�$hh4kI.����eϴ\�	�#��^hF���@#�]]�H�SF4�'�5�g �Fwm����$(��AMkY8p�NW��JwF�eщ�r]k%60��Ĝ�T)T�W�K��U�rQr�]������AbH1J���N��ꉯ͏�M,�!�7ZIL�y�R�n	��	L,*.�k�a��]� �~B� $i�����B
��8#�0�p�e�6s��ai��q�pcdI!IL�m8b���"h� ��<�F.�������F��8�a��0�)�����v���"�H��E��Wjp?Q���?	!
h�g��$�(iL8~?$+�a����MC;)��f�\�%�S�4Ҹi�1(iėX��
k4l&��ȡM\3[8~H$F��Q�o��%ռ!��1��p�l���,��!���Y��?
Ŭ4k\ֶ~9l���%6F�`h�9g���R7���O���^��k�`A�jOƉ�ļ��2���s�.�6�a��	 �.���X�w�e�cK�_Υ��pk�4�(s7����۬��f��H"��6E�#.`;�丐���@�����
�!����*��V0�@�Q:�B+�J�9j����FП���HJ�HE�����4o��l����M���%��:#�dYQ��!QІDX��!Mo����ԂV�ڝ����M1�#2L�e�B�7;~��)Љ��-Q�:rB��D���L�RBCbFWD ��#D8$	)UBƆ���o+YĤ�edT�������)'�,�Eȅ��OƒSD(]!��1H0���ټ])��(c#
��kF������d���5���������;I^3��m^$*O��g8�^	)�M��5ћ����rhܤܸRS�l%��g46<?3z0	6��!Ixa?L���s��l)��ƺ��k���Hš�8a�Y�����z{��ױ�k�ӯ�=g���� ���      ���       � �                    �                           -�ċn�cy�5e�m��;+�Yn�f�^R�$�:[�� �I��f�ݴ���Hd3d�Ʋ.mm�mpHR��e�n�zv� ׋I�`��ݲ��Pl*�UU@R�� Wc+�ĵ@�3���U-i0  u��n^�-��o�m�ĚmZ*���΁�� ��H�I6	��6ͰI���k�c�I6�hך�WeU^�6{;l����$��l��\�@V��ݺ-��2UUK�
�Vєx,�;��%��괅ʤ����WEp T��D\q'm�     	   -� 5��      K( �[@piX 	�kM�v� ����Iy� kY�X�944���� ��k(�dm���vc�	r������n�R]%�g��1�mA�`GA�Y�3��P�cR�J�U\�ev^U���@��l�5��W)�ir:n�rZ�!$ �ݤ�  ����`-�Hl���hH��mm�e�9  [E��iJnV��ʽ s�g-� t�r� ^��t��`j�ͶY�g�}�$Yڬ������$��U���Z�ܻz"��bۂ9��Kb]#��C��e^�3U+i��s�W]
�4��� [@u�mh H�   � $)D� ���    �        �            �����U[�[�8�ٛ�ϛ�|�c�2	\�^�f��vրHX7i�9NI� X擅@�3ΙV��]uWm -$��[W�@l��m q�ҙ���-�  r8ŵ�kn����k�l�����ت�X�k
���JD�S�m&� m��Y�����૩V��쪵J�:�-6 �/H���U��۴��m���m� �`  ��m����vÂ��ݶ)Im�*@pm�:�m�ړ��8��sk�ɛ6��A�Wl�+��ᶍv�m�K:��$�[C��u��6 �nٳ.��6�ժe@���[@m�ei���uu;�y���J�Tj�M�m�#�����*�U�Md�I��p����[�:�.#9�g%�����8 	!�f�Ÿ    p   m��P�m��`h�-  H� �H�Ğ-�  �m��lm��R �` M��     �	'I $$X���  [WM�t-�݀�P H �R 6� <�� �m������l�\ ]�[U�`N@ kjIY��˕���� ���[_p	6@j��}.ʱ�c��U@�V���H�`6�   [@Im  p$5�[e�6��&��ʷmlC�� p��  6�-�����m�k������u�'A�mT�0M,f'ʵuh   �n�@H ��%v΋�}��n�qͶ 	����h -�M/���^����  ��e� �q� Xv�[5�0Ӥ�� �md��.�Zl@ $  �` : 6ٵ��ŴI�� h�Nh�-������ӡvy��YkK����  f��N�$�o��� 8n���o` �m �n[d���ҍ�;n�뫥Z�i��j�m�kX�6��� -�� 5���.���5�쁷� �:���u��U��H.��m�j���p	 m��&ӷ�;���  �R�:I:�� m��x�]z�:���)�H:�:#� �6�j�����v�R��@'@�p,0  pֳ �km�mni4���kt��t��[DN�$��Hh�m��{Q�ڥZڪ�%���U1��V��/[��m��k $'A����jK�:��   �[p�c�h []6̀[@�Ze���oav��sl�X`�6���ZI�h�i�b@i��`�^/Pm��$���� �v�5��D�	6�:@�� Zn� ���ڶ�@� -��Am�nݶ�  �n� [@�3`H�a!m  ��ڢݵ�� m�(�5�U���U��[u� l��	lh    se궶��p�[L�a��]��}�hp �`         m��  mZL  [%V��s�� HR��d�   �8Ӷ��6ض�  $5k66[ @�߾�ko͝u��g	 	$������Ŵ  � �r����'[@ �%�m�U͋h[��89��n:R�-� m�  �������k�-�h���]�!���� mt��g8�2Fҭ+� ������U] l�f_	h � ���GY�l�co�|}ʹ�.  ��eY�Uj��q�ڥ@Kh nհ $P�0K��R쵻�ҭ<�����X����U�vYBn�j��շ�-ڶ[C� 6�%�-�� m�  ,��m�n h���n@�p��rA��	�  A��b��]���Yx
����i�6݀ 8�m�l�ׂ۝�    l� -$޵sI�� h���� 6��   kn  I)m�V�������	$ @� �-�m�  ��Yn�V� 6�g  ��@���N�)vݴ� ���J�|�  (Iy��l[Ku���a&�[T�@ �P V͗bW��6j8A�� :NpM�Ի������]f��t�m �[���WP6�5�a :v��+� -�)]�랗j�Z�U� l�m$5��t�_Db@�I( m���=,�݊j��Ʃl��C 8�UR����Omu��j6��-X�e[E� vq��6���S��g�3 U]uH�z���wm�m�\���6�[VȺl%(mt�2��� [m�d� ݶ����`	e	7m��9��|��sml���C�-�R�$,�nź��a��n��/C$�n��ͤ�ذ	   m���[YF��#*f��\r۴�� ieNt��R��+7R��O/`]��+`Hm��qm-��`���i���Pu Tf���
K�N6��yn��
��U�ݲ���]_A�v�H[@H �� a��4�mm��K�]�5���G%�%4I@����[]������6ۃa@  6�m �����kh$��X���%I��� �v�-KqKUU)�B��B@[v탚Ȧ�i���b�  �-6    H�� ��c#m� �����m䅜[p@�m�6�-`   h[@Xu�-����� [A��;M�m �ض��չr}��>t��5R3e�2�V�U �$Ͱ�[@�6�9�n�'MU�Cm�6������B�� 5O+\�U �0X���pp�[ŷ��b���U����%�|��>��Ŵ�m��[F�rޠ`m��m�6r��`m�;.��T�e[nګki`5��K֯Z  $m  ����`��ݷ`p�٠
+����B��T��<�M��I6� mRm�l��� z��m����ll��@�mR�*�A�T1I�l��*����8U��mkr� �Mf�U���۶�[@ $��TY.�6�U��\�P���h�\�m����m�m����d����K���b�
��^���h��ۛ�J�!3k8�ۜ��:%�0m�� m�vp�J��wgh
�@]m�5*��I�zvܭ��U��@r��c�]"jj��6�l��� �;I�֭�Hu^m&[W�[@�%���`M�j�r�퐭��#� d$٫v��m��[��      m� [@�W�8�         @        �6�  M�m�s���Tnc�  +����ڬ��\�a   �` 	 B�M�j    $ �     lm&��b�8����@ *��q��iתIlm�r��t�ʪ�������m��p�k�kkv�@��ٵ���ֵl pqm	�I,�  V�uUTUVvT�f��Hݤ�����Ci6�@H<�N� ���;n�l����>��[.���;$H��ݺ�b�\�,  !ź�,ku�6�iZ�'8�l����Ch6
�3:�����{���"�PE�O� �@�@�@��4U]�� A��W�8AM����pP]"b�F
�t���q��U�FEҊG����)@t
+J��S�L �� �/4��
��j��4( �!���^(!��A�]����:��b��N�-�E"�� ��F���C�@���� �S�~E6�����P�
LM�/Ȁ�� � ��k��(E �
 ~���@��v �������?���l�PD����t��"A��@x .��è�UꀔH�b�@*��DO�	�P>b �Dj ����� v��/�� s>C���lO�!cb�@!
t_��	�!�>Cb��@1_��'h��"����J�� @��Ê�~��)�H���H�:��S�!�`�����T��@����8?�PUx#��D���
���_���l �n    �ͮ     �5�#keeZ˵�!O]�j8�7�l/u�X6�˪�D,���nlfPWĠT3�܇1�u��m����j�s	*.���]`�+�mq���*��� �De�"�(s3]��̬�n��ǓbM�yvJ���w�t��[�MU+�2UUT08z�ڔ�zǎ�:�\�xiȘh�7m��n�8t����	Px�7F�5<�m��� b����w��c��j逝<Ɨ\��5GOB�֑j�h$ �����r�l��Ѭ˒%�5�^iV�n�"�Q��by��%fG�eA�x7�!��ά��#jt]�\���Ji��+�]�l\W8��ȵ\���&�W+Z^�܉x���BuOH
.nqI���^ȵnC��\��f�9xLmqsh���h����u��6l[�t!�
�G%t��v�B�bڀ���T6���eܗ�Z�T�T��nW�H*uh����[��)�Z 6����B۱�Y9��e��ш27^�jݵ������قj�"�vɰ�$����ʅE-�V����s�r����8��GEV�ܘt<.���v��❓vy'8!f�Zm ��@�%��	�!$�C��v:���٬m����ˈA�0�]v�m�3k�6t���4�����n�e��@�:�5F�X�N�)W�6��s����nZ� �<n[�����Q�b�0��'6C�gM͉�C�F�2Y#���df�3� ͷl#�J�I�0�Wy�B�.ݺ�=�틓�Hꇩrvj�Ah�v��Q�8��ۘ�D�`K0�{�X�t]��e64��K��������[�!e\��Q0����ǔm��e�ã.PR���е5��nv���w]��X;K*Jjm�@   n�m�r�KX�I�6�����'^�n�$6��@���]Ô�i�C=����S��#�8]�na��Ը/�q�@H����A ��LWg�������޾���jڪ�g��m�<ka.�WL�3�TTiy�0�D�NYv*��Ɔ�2�l��M�I������j��8��8�s�-�-�6�nq��l�3�< �Wn�9;g���3��Yj�1DB�\dxQg��H5=]�Ցl������`N�x�D�t�8��;Bn-�l���x����vv��㭎���4%��:qnP�������s������Gh��v6��dQ^7��q�\�n�����7.W��#��
HOIo)�{ۋ �����y��.%��~߱`���Q��HGl�����}�ns���lB�J����7w�X�n��?t���Y%j�l��:�Lގ��GLmȘ�����e,��S������5{w��u�w�Iq=su�����Wkh��^+�`J�0=�"`N�w�X溞�c�ƭ$�;	T��vn'ԂArޞp�k�D�ґ̖^+r@A��,�Y���܉�:�Lގ���� {��U��Q����w�P8�V!$@� �)(؅���W��`=x��M� ~(�+V��+�;�n,WH��uȘ$�O>/+
����^e0%t��ۑ0'\����� -���U�B;e$RJ�ݛ� �P�)��=�x���X�m"�	�3�e�z��۳\��c�R�iooU�/,v[�\/*��`����],uT���D����+�t��܉�nй��e��T� �}��^�ŀ~��x�n��qq&��jjo+��Z������4���>�78(J$ID!BHr�j�?"gu���I�ﻳrO�=S�(�n�ڇUv��f��7�u07z:`J�0
݅]ϱU�.�Yk/10'\�����WH�������s�F4KF���ajG7=/g�	�z\hەK\�) �FZ͌]�{�GV�v�m��߿�`��� �ٺ���x�v5���Dմ��V+�t��܉�:�Lގ�N��ee�-�����f��7�u�y����n,V���?t���Y-jڻ������׋ ku���
"�)6��D��������N�%��p��k�������۸�ݛ� �M׀|�\\�{��؛�X���q[�7	z�ݙ�6����Ru�ם�v��X�ջV�������j��\��|��ذݦ� {M�$����`�2z�Ss3���K+e0=�"`N�w���n�����V�dTv;-x�lLގ��GLmȘ�*�F%aZ����W�RO���X����?vn�}7^�ݍe�uQ5m#�Հ5���:"!%���u�8���2A �$$$�Y0� K�	FUЮ�) B!���(F	6,QjB���w����7m��%9t���k��݇�I6� )��-l�LSW=���X��'[`��9�]#�g��Q�σu&�b+-+ w�~|��^�H�y��D�i�N��Bs��3�(b�&s{:%�3J�"��^zn+��y��;:�й��`�#[�Lp�IP�i�G9�x�>ǩK��1������m���&�Sa:m�i-�`����f��n��(��dt��D�M漜.����ItMq���B�ݥ��o]�^u����8�ݮ���s�{��lBJ>�i�ŀ~�;���B�Z�K^���?��"d�}� ���`z�� ��;#����,���w��WH���7^��MM�v��U�Z�X��:`{nD��r&���n��0:�Q��d�7Uv��f��;�u�����X�t����¡�KY�lD�vK����[�:��cr+gX�.v�7C���5+*���k���|��GL����r&튮/��k5�˹'��wf�QN@�F'ً �[Ӏy�s���5�R��:�����j�5o���u�ٺ��ۋ =�kS+�ȭ��j�Ձ�>��z�� ����5kx��M�^Y%j�K^ݛ� ���Ku�����ذ�M� n��PTnzW-�m�s�4 4�A�/1��u����en��9"GJ��.B9������?1���t��܉���Lٔ��ْ��\�ʰ/n�ϒ�I6w����<����;�x{En�婺���s��۹'�뽻�P���ABĚ�P���˷�`��E8�Y���e�����r&�GL����f���֦���lUB�L��遵�0=�"`l� �J,7mQ�����ŝ�+Y;eݛ9�i�Á�=/��9�GB6�?���VN�{7[��$�x	S����Ll�07z:`�֦W]�Wm��l� �ٺ��ۦ�kŀy{^,�%'����p]]*Y�u��107�gၻ��kz:`{f�����Wl��Umv�%�⛯����,�Ss�(IlB�D ����]�&�}�)����I�f+�W���ގ�ۑ0=� ���� �|��b�TF�u�割�,Q�Vc�+�靊-$��[�d�q�ۧ<��]�b�$]�U��Y���܉���GL��q`�t��V�dTn��x���:dBUF��XO{������M
ݕ�,UB�L����:��ŀ~��x��� ��ڻ�UE��[2�[���r&�dg�Kw���{�kS+-�Wm��l� �ٺ��v��׋ ���X(�����=�Ҫn���׳��sq��,��Ě�h ���X�l]jXh���t��[��]߿�����v7������>5�7g#�Tf�1�7-\��C�t{v��@���s�8�˽���� ��볮�n����׺��6ms������,��6����lZ��Į�\A�	p��H(�Ȁ��V�ZE�Dq�.���nN�7h�\�ڤl�=cq�{�E��-=\���ǆܶ	4��Ħ��Nŋ�N� �',�:��ɠk��3�Kд6�����m�z:`moGLmȘ��>Ř��+0�������z:`{�D���D�g{�5���4Z�r�U�y{^,���	DϹ��ذ��=���c��%Uڰޛ� ���`����n, ^�mjVEF�w8�m�(Z�|��}� �i��7���&��X+H�NJƤ�+�v�n'l4�P�$�<����t{��'6�W�/.��Y�07�:`uoGLuȘ��Lۻ��UE���V��x�Q	}@��I$�+i��>{l�;�n, �|֦V[��%��V�uș�}T��GL	S���;�����\��}7^��q`�GLmȘ��>Ř�1b�ʺ���׋ �P�>������s�}ė8����5��8���j!*d�B3���=����y�H�v�6�	�N����מ[E��-r��|��`���}7\�����&�h����IUwk >�w��!L��p�ذ��X ��!7��Y��n���~��vn|#����� iq���#H&��D�$��j��ٳ7
M�V92B$�hFL�5)@5, B)��QM�,kF��>�$H'�E��Z8���8&��vJV-���SAH
�TMF5��Si 4�4j�*T����O�� ��#���O�(��R���A7�O�8�D�)��|.�A��� f�����(��$�����;"��2X���^�s��O�߿�xｳ��r�?}�f��"�����uʻ��X�]��""r��r}س�L�����&y�t���rK��{���~����وK)�
\�A�B�i�UcYu.�:炻hk�cf���5-Wm�)-_��$��{���$��o�?��}�IL�}ذ>I)�܋���*�m]MM���s��*�����$�.�� {{��ߡ�
.�h���[��]t*�W��q'����~�_-����}���M����}S_r���j�5�	fU��O�tBS!���P���^I�?� 4F*RS��'��o8o��~�����&�[����Z�.a�'��{9$�G������7_b��$���Xʦ'i�@J����ӎ�p��l0��	'��������K��m|8�n�c=bqU��������Ӏ}��_��báB�=�׀ޕ\�&��*�Z��P�2�~u�,9(Q3��b�ou�B_Hs����$�����/	UVЮU�|��g��I���ӆ��ϔ%w�?��t%2�Ңee���$RZ��K�w���>��8r����}� �݋�B_H{��E�utw6������""y�t���r�_Hs�Ł�>�����N~�UUw`2�n���:Z�M6�!K���9Ŷdw���9wΒ�8ά�n+
�i�̛��޵��;awj�v��:qTY^-c����uu��iBm�+�\;�GȪ�gRq=v�yu��:�բ���;)KU=��[n�Y�st8�psݪX��m�k��#F�㋅q	b8U��ͳ��Mk�rn��aY�A�:��NS�J�N��{��?{������n�pL��]D��j}:m$5L:z��t�5�9g4y0�n;�Emr�����>�?�� �݋�/�=��:��yD��t���5�--m�\�ʳ�ٿ}�,����_H>�������,x�OX�n]�[T��V}ě;��� ߧ�?������b���{��~X ��}EZ��Q���:!L���p�ع%H>�Ł����}�|�����,�%����rIN�� ��B��=��8��ѷ������lm�c��S*�����wg���q.|��ӫ�wi�:��^��9���ʻ�f�`}����`��:S/��� 哽�����I�����̳3T˙��ֳ�8����?��DA�(���(]Ok���I� ����w����(��3'������f�Rk.m]QWs�~���s�!B�7_b�wb�q%��;��� �ȚϹ,���B�%Lގ�$t��܉���Lٔ�����j��\� ����?vn��7^��q`���%I�����78vԑ��6�����7QgVTȢ�R9��\R���G[��j�[j�?vn��L�w���GL�aW0�Ux�Z��Lt�07z:`ott��܏ ����4YFKR9e0�ۋ~�����H���v��9��۹'��y�ѭ�%TR��`u..3�:`yl���L�w��'EWH��5]�BKV��u��..����{~ŀw��X���ǒX1�RY-�箮-����rknژV�����y��s��<+����Q8Ya��!-x�m� �}���0=�"`M�����^e�Y��w���}T������Lt�`��֪Wkh�Z�U�w��X��Lt�07z:`{���U�K-]ݪ�wv��M���f�kŁ�	�Px�}���rHw����e3,���^b`{�A�uUU����=�0?vn� �ᰭ}HƉh԰,.�������x��΍�U�´�]6Gj2�m��9��e�U#�S��ߌ����?vn���� ���[DJ��-��i�wtt��܉��2��0	�]2����,$�`�7^�v��M���`��ŀ~[7Q8[Im,��&��07{ �����ճ��e$�ڋ+��;�]0{ۋ �ٺ�۷LY��ؤ��ݖ����[4���"����H�5�r�ݴ�;tS���{cs�n���:�ɜ���&�=1d�O�Ƨ�9�l�=��C#@[0�::�[[W+�#@�v��֌����w(��]��jY�SsqF�U��z�Ma5�!��2�l؛1�H&��n�q�����D�zI1%v��Jks��ޫ�pݕ�!gi�9��.�˫����yT^�'�?�ߧ칣G�g�i#V���7[O�R�6���Hε���c�#ԵI�%u�[�D�'�I����>�78��?%j��7]�n��� �v9mR+mX��ן.%ĦOw_�0�x�{̡خU�W�,����� �������wf ~�jmYFWJ�e���������[	�W�-S ���j��QH[�� ����ϻ� ��t�;�]0��ֈ�j�K,�F���<=v��Ϟ����{t-Y�����8[j�S+-�-��KV��u��n�{��{q`���N�B�K!-x��3�BKTcV��[�� ~}� �ٺ�x�l�'�7��Ik�,�� ��ـn�ŇD%3���=�|`�T�ф��Z�0{ۋ �ٺ�۷L����ό�'���v;��u��LmȘ� ���������N�@��\�ձ��]D�6�GV�W§Ppj۵ 6�m�S�.�$�Na�b�2�
Yk/1xِ`n�A��Ѭ�f��ۭMU��0��-0{m�ДB�}� ��t��s�l�ѭ�%TR���7wq`�7^�
#���Suy8��� �uʨ��0��	-X�ğ��׀~ٺ���Lww�l�D�m$-�Y	q0$�v�&�:`{nD�6rqϷ�OC6���t&'i�]���U�lf���:6�d.��V���͖��E�&��L	$t��܉�%Șݩ�T�V�Z�-��wwg9�6{nD���v�&�|)XZĲ���wY����܉�%Ș��0$� .�Hmj�J'c�׀n�׀{ծp�ŁСRT� ��%)$D �AH$,H$H"�a�H)�`# ��X����),��h<�G��n����I;���*�eZ�Y^��k�7��:`{nD���L],�Y��Y�F�8�0<R!�ݛ,��0㖌J�rOmZ"�r�[��DJ��-��k�7wq`z���nyD$��ݧӀo�T]��a%� �ٺ��%�q���<ޛ��7wq`���N�BYU��� �78�Z�Ir�U=݋ ��t���5�R�I+�%$� �g���ŀ}�np9BIOu�N�֥WE�ZAy������GLmȘ\����_v�I�C� |�0zF���C�:�Թ�� �5p`�!( F!J��H �L�	��#F��2Yڔ�	 C�XY|�"hH0�c~�hHB&2��5f�@�{���h�&$H��  D"F	W6#Ab����A�4�ab���� ����iȰ*D�H2�
A�EthF��FH���"�!�K�8��!�,b��R"I,���X	(D	�))*J����BÅ��܃, ����#RQ�1
Np
��`�B�i���c D��R+!���kZ�333  ��   o[@�>  Y�v����m ڣg)�6vz�tKӞg؋�!+\���֪_i�Y�9jA�7n��l�����*�� �������p��G<Nq�U������Y�]*�j��0e��Ԍ:����U�x�R���L�s�M��|��v�t��W;st4�WUU+�2 gK��v����mu��[k�/.ۍ��@�������[uN��%�F�y�j���v�v����{j�s�;����u��n���r5�j��番������5O�n�검sU:�Z�,��N�r�J�[�-�3��9��ǳvU,����Fx.�t��z��E��<F�貱�[`ظ�;hbuʻJ�*X���<u����;k�tV��MO	�%�ɞb��Z��� ����^z�����E4�gu�ngu�v�q��)�;T��u-Q�J��W��^&�nѝyY��j����ƙ	�uc 2�o�n۔�����<� UT��ڤ�nz�%�Gn�������E�V����rJ�c%�P*
VD6rex\��9��z���0��٥tT�V:�FyY���BZ��%�e�U�fw���IdZ�=by���ݵ�Z$��D��ƓZ�I"s�M�JmV�K����I�k\kc �g�*�����mw�6�v(�u��*��j�s��������'P���qZ�LA���y�*��+1�4U���c@�{�|��S���e�2GG-��z�Vv�	��p�e��.��;tu�Z��8�v��<��+u�k�{ �' Y@�������nH㸩j�c���{i61���ՂkUz�H�*�zw3���ꚝ�dzX5%�]�����:"��o$��Uu�	�k%)s"M���ޠ   -��[m7X� ��� ��X�j�.�W ��]c�*�ϛ��J�c��Z��\��-���e2n�&�Z��ؾ�P"Pڨ���A;�EN�<0B*:rk��30�.�^s��}��ä�
�iͺ�N�!�ภle������.�K!ѷk�����1��9�=���ll�ٻ+���DHs�m�G<KkJv�t�(��F:��G�H"r3��u�j���-��9"XӴđ�&r�N��U�S=v�@=��X(n��k\Yr��v��n���]gY��坽,����Ye�Kz�(Ʀ΢\u'n]����غ�yz��@�N�J5�ck��F�nt���eC[x���-�-�ŋ��H͗�����s�`Ir&��L	$t�+vJ*�*�N�e� ݛ�?�s��ߞ��ŀ~��x������ʥ�\��k���a�BQ3���;��p?z5�D��B�ݶ�ww�$��"`w\��{�*����Tffe�y���܉�>��Ș��0$�� �}� ��b�KTd�6)k2�E'N'4ݩ�zr�❎l��8t뛡��]�j�uyyX��K�07o�`I#��n�����b�RHYB�,�;��{��Ad`E��I���ٹ'o�{[ �ݹ��I�wjj}�ei�k������X��X5$�� ݦ� ����H�v9e$Vڰ�ݘ��p�np:����`�⎱\�-U���e�$���L	$t��$��DoT�l�r�%cRD!�=�ۉ�i�5@Dr@�b���f�N�ť���R��U���zn�ww׻�������}ﾍL*���G\� ����=-��5�s�n�s�#��UE-��KV���L�7^�K��JQ�	(�_}�[��;w�`xv�30Wf^U�����r&�d$té�n��u��,�����W�n������r&K�07{(�]ؘ��X��-ԗZ���u���-ն���=�yu{\ަ8�4V`t���r&K�07{ ��|%�����k�[j�?vn��7^���{wq`�t��WJ���j`{�D���7ꤗtt��܉��kWTl�WI]V8�x{��{pܓ������l@X�#�����x�ݍL*����S ｮ�ۑ0=�"`ovA�6�)i^V5���RI�X�Ok8�Yu�ԍ��k��te�Lh�h�ӫvZ]5�6�]r&��L��o�^@�����1��qK*��^��u�ˍ�ݿ�~ŀ~��x�k�b�Q�[Q$�L��07�:`{�D��\���*jo-������� ｸ�ޛ� ����ۋ �f�j�(�q��W3)��}_lˉ����{��I�W� ,��!V�r�٣Z�eUG��`e�;]v����2H����'k�ԴT��N��ԝr�ٵn�=u�l��ӱrq��X^k�Dv3eU�m��L�v1�\�ynHІAJ��R�u����\c�L��@u�>�9�g(n� ��C�ao/Z�qI��m�w]�>f[��;m�y�g�����u�(Z܌�N�^�%��m:nV�x%П�|�(d��d���{��w��bb��Z��,и2;��Gl0��	'���բ5��K��my��E)T�v;-���<ۯ�׋�
#�:�ϥ_*�.�t���� ｸ��%����߱`����]���m�ݍL*���y�$��OW��K�L�����َ/y&����o�wkS��Km���ߛiuɖ�I{�E�$�tlI-y$��݈�-��YUv[f6����~m���4�[�=^�I-�2�I/I(<�anqpL��]D����5�$��0����v�$�8n�Ɇ�3Ѻ���^I.��4�[�=^�I-�2��W��[35���~��6��ZjZ�-r�6���s�T2�k��n�o;�����~��}�q.%$o}~�TJKY��3+�I%���[I%����]Ѱ��}�������٤6�]*�N�e��I/vH��I%����$�W������? ���s��C�f�a����6$��諭����I.�߲�I/vH������gc��sX�{�S��k<��8���|�s\s�1��ztί
[�u��̻�̼�K{���I%�&[I%�ɯ�����01��f�֧,-��I-_�6��ݳ>IqI�߾�6��ف����o���m�ݻ8[G���m��w�g{y�m���rn� D >W��Nsz��������}f6���y�V+e�ڋ��^�IwF��������Imɖ�_��\JN�}�����ma�-��Ե�Z��K{���I%�&[I%��IwF�� ~=���6��!:��LC���Y���!�v�����ʍr�(��JWuً�V��ffW��KnL��K�=�I%����$�[r�Lb/
Yk/3-���G{*���wF����t�{�m���1����jj�����{�%��K{���I%�&[I%��6�J��V�%��6�I.rk��ߎr�o���[��ϻ��r����T�DM���7m����e4�d5���]�W��KnL��J}_lN�IwFɻm����9�m򫯽�5o5���hɬW��ژfq]�f١��z;y�����`��/5=�f��S� ??~~ﯤ�I%����$�ۓ-���tqU��/WY�w���I%����$�ۓ-���d��I)#h3��X�U�,2��I-y$�ܙm$��$^��~��6��n�j���8�r+m^�K�}��왍$�����I%�w�����ٱ��Wk%��m��o�$�y$��`�It���$�[&cI%�����}����ݶ U�9^��is��
D�]S�&��^-:� �5�>��Qu����3o�v/�WkMq�I#Qc��v����n��\�Vn�Nf�';8�͞$\����P܆%�ɶ�Vk=#u�熡���:YN��5����ٱ�6��[�a�WL�u����;N6�&�<u��]	���k9&��O����:Ki�Y8�s�G`P����w}������R��Z4J���*h�V�x9�*�s�<*��F�եU�L���6du�C�k̳.��?�I~���K���y$��31�����ߛoukj�	U��$�Pi$�I�����Wv��3I%6L��K�sm�wv�9ah���Ij����왍$��&{�%��K���y$�˱������Ym��m�wo�ͷ�k`�It���$�ۓ-���H�բ�/������$�tlI.�z��[7l��oۻ~m����d�)��,P����mˋ�י��ms�'@΢۲F�p�:���/���>Ϭ�C/^�Fd�Ŷ�߻���I%�&[I$�I��IwF������������rZ�_�6��ݳ>�_�b)2�k����m�}�ɻ[~�����m��c[@��J'c��1��ܒ��I%�'��I%�&[@�����R]6i�L�}������{��II���$�ۓ-��ے_��R�H,�%TN+dvZ�o����~m�ۓ-��ے_��]Ѱi$�l��+�GV�J�U���@���-�E{;���ӹڨ;gȢ7 ��1ϧVf�Zﯠ�&[I%�$�y$��a�꯫�]��������~��8K[�[JՖٍ��7v��I%�'��I%�&[گ����Mͪ1[(�VP�K?~m�{sn��{Ü�6��%%ЉX�"A$l(X��,��q2I��Pb� ��:�(A��@bHR���� !� B�߄�`�C
��;�D4�W�)>>Y��E���P) E�L6c0�EH���J�е5��|
�'ȔF(&(�?)8��] ��A �� ��R�T|�6?=?
�C5��~�kv�~�~������Z�5mt���o����~I%�&[I%�$�y$��`�Iwg
�xJWv�-v�ߛm�nٍ��7v~��]Ѱi$���{�%�������N���ˀڠڻ8�w9��q��b�X+o�kBF�;<����'V�Q�q$��K�����$�tlI.�=J���޴��ݳm�|��#�R[)e��6߽�K�OW��KnL��KnI~�IK� ��q[#����~�����m�ܙm$�̑{�%��Jvt�Ue^`��1]�e{�$���i$�d��I.�ɻo@D@��s�9�m����4�en)m+V[f6������m�ۘ�o����~m�ٻf0=��8k�W,VB�ۇs����&a��Q<�ηS��[��\
F��Vxv���n+(Y%x��L��ŀ���;�u��]a���V�L���:`�ceȘ� ������(�rZ�X����7S�}_R[� �����nZ��`�h���n��_�x����=��X������T��\��Z�x{�L�C}�/�7{� �� 脔z�EX$b��*H�$	Q�@H����D�P����U�8*����ͳ��丑���`n�դ��IeFx��w�m���W8�FRG<n��mO7J�/ �O�����I��w]��5E�۞ٶ��v� ˦1=��T�;c��e	��h�u��kh2�[�I�yn�0���v��ֆ�-�$��%�s�3���یK�ɺp�E��<�o��=�/ͷk��;��xd]������w;&M��[s~}������Ӷ�1���杔2��!˻6[5�Z��i�����UN�彞�LGl�[)�>��q`{�p�ۦ��� �f�NU-��$�`{�s�	(�=Nـ{�ـ{��`��EA-n)-u�-���� �v�w��X�����݊1K)VP��`� ����nɌl�06vDT�V���Ye0�ۋ ;�ۀ~��0�n�{�VؤU��u�b�O�s<۬�m��6����y�[t�ݪ:,)xJWv�-v� �wn��t�;ݺ`��vljj+v�^7]v��9��ٽ�~ ��!�;��M�w��, �wn���Q���Gl,v�� ����nɌl�0'W6�8ZRF�Ke0:�}��{�pݞ(�z��;�합ʥ�v��� ݓِ`ñw�����]8��B�&����[Q�l�8��rK��)�W$��U�Liz��5�����`{fA��2ގ�����݊2YH�v�[i�w�t�;�n, �wn��t�;���*K,MI].��=�x��n��QiDB��B� I%*#�%d�_���L��D�qGk��j��v���L�ۦ��q`�fƦ��k%�u�n0=� �ݙ쎘���E��w�>�wVF�n݈:�n��n*#��.^Mt;=DƮ�
�ݒ`�I�x06vA��#��&07fA���[xZRF�i�w����ݸ{�L�����Z��Z7m��̦�&07nD���쎘o�"p��(�v+-�?z���=�ߌ�o\|�%
��� ծ�*�U���b//106vA���� ��7^��6���ʚ����z�'2�B�#�!�y�s�a�]�ն\۵���BUZj��m��;�n, �wn��u���0�h֪���K]� 7d���Lِ`n�t��m�Ur�K1�%�f0=�"`ñw� w�� ��j�B�\���v�vd�0�1��.�ŷ��$n���{�ŀ���?v���v��$�������~�UD�.��5����H\גz��]��u��蛥���K)A��=�ol�I:�9�)���Mv���;{]����(�F��{;�Wi�9�ط���qqh咮�9	��^�ީ��Gy7�k��ݬhg<��b'n��@��P#�wc�:��[�Crdn�7�m��sn�v_�m�W`��!�m�Ӳ�q'k�
��s���U�{�����q��f�v�S�'k7;1y�hڬ�V�z�u.�rm�-�cD�O>�u�����m�>����܉��2ގ�ΗE�^`��Ee� �ٺ���l�����b��v��v�Q�;\�v�Yk�;� ����nɌRK`l씪���Յ��)������� =ﾸ^�����ό﾿UIc�"�.e0�1��Ilِ`wH��_~��~��uel�$��/a��)�nu	q,���D5�i�뫯��{�t����Q�������:���`�`�����}��;��~W+�v�JYf��ٿ��UʼZ�ﹳrI����'绳?��l��_^���lvZ`?~t�7d��%�7fA�Ɋ��T�[e�Ձ�9�߽�� ������专���� =��8KI#r������`�"!o<���ŀ� ����J��n�ݩ�V�Îd�B�v�K5{z��QKJX���)��$��"�Q�䃵��g�=�ߌ��ŀ���:�v`�]ME%R����)�{[ŝ�L����6{��y�3�D%,��͕RX숲�e�`��� ��{��@�*QF�����>��ٹ'fƦ��(��u�m��.q'���Lw��u�X�"L��^�r���p�����Y�w�t�?��9��ߗ�{�׻� =ўd�
Z5k�J�F�!㜹۫M��>E��ѝٍD�3�u{��\♘Ae�iI��e��7~� nɌRK`ñ-�_�++W�uuWk =��?%�興UC�߿V ���`��, ��b�D��7+�Ym�=-��=�lâ""e��X��x˻v(��H;Y\�`|��$���|d����nI?~�srEU
����qs��{��&�۩���X����j�u�X%
w{��6{��y�>m���}��ue���.�)q��.�� Ap�%gV9�T�ʸ�9'��]l�",�YeX����wf����q$�0���XW��'ʷ�n����Y�%�DBUC��w~�� =��?���ߵ��B�R�k$��`��� �o�D(�7{� ����l�Vp�����d��8�Ow�, ������`~������ ���Q6�YSWyyw�LvL`j�[vd�:d�]����$Iֿ�>��$��"m��ف�X�֍�: �Xb�M�{� D�H0��ĉCk mA7�\��B;Kh��y�K�5�QI� ���ta�D`^�(x�*J~Ri��w5��
T��T7TU!A$Lx����4�hr�4 ��BT �@�Z HD ����KV�i,e ��R���'=��������m�  �   ޶�    $�S]����=�y���U�öQ�n.
W�9��복�
;-��
m���nX�Kn�m�j�V�����b���٬�ukn�yMeޕ;���n��IG#���v^��l�!��Z�5 ���x|v��[Rv����\���v����7@*� *�hm%��� s.�j�6�+۷f0lp�v�4�9Ŷ6^��vv�b��d���qi�Z�C��GYx��&;� �E�&mڌ��%���@F��j��fIj�)���%$�9�M��n۰6݆B�j)�W��2r�����]/l�6m�Ca5X��vU�����+�'�`y��V�"�˘�lȆ˳m� �J���N����X�����2���`�`��v��3���[����CJ �N�gۄhC9���v����C�x���`#4�� [�S]@uXɝ�%u��#����+4�k!Ԝ�b
t�Z�6e�)�!�Z��rJY 
����8��cs.]�������n�5^U��(�qT��4ǜ����l-���H<�pT�e7a�`蔛�3��[�s%JD�u�t鄳D�M�lɌhZ�c���t�anڃ��q�Z����(�Wn�i��ni�vv3����Y��u���N��ui**^Ρ���*p*�"[mۖ0=&�0vs]d�gbF���^����Qm�j�b�6���r7-��Hc9��0Ŕ;�ƞ2�^�#�jmN����\ch�$���L�n��+hw/	*�T7�xv��+�رԾ��e���0�� $�n[%���p���kg�����.܆N���)U��!탄�[u�F��ӦlONn��yDw�B��o��j��a�*м��T�+���a:.�lm�� 6� �*ۙ��6硛l9oW�uغ�����#J�Ar��
�T8�ٓ�,�cnƁ�[��J�+;J܂:z��W� �~� ��ޔS ��Cj�LD]�~T���>�ֳ33335e��僎ݵ�k���Mp�[�t�屻IlhK�������ҋxV�-t�v�u��, �aUhp`��ƪ)��u��n�	�\I��W*[i�7EX0qm�V�iS��lv�t����<V��١1�@�kmT��)�[��[q�x���W8M��}�q�a��6$���v{+���HmgV�h��gk=��nV��Wi���b4,��;�Bݙ�͹��qv���S�óћ�D7m���9�盧� r�Jۓ?��wk�̊1�HܮEe��u��0�n��x�!B�@���z��H�n檉�F+����0;�t�7d��%��I6{�&���b��k��`�}��7d��d� ��사�1b�!ڥ�U���~��\���`��0>O�߿,���व9x�u�pl�07fA���� ݓ��Ժ��`��f�ٸ:׌��sNq�M�s�<*�l%�mZ�LH5����G_6t1��e���@��_��=�x��n����x���Ғ7e���{�ş�K�\v�D6�|�?�N{{��9���;ݺg�\�l׿}b����YmrZ�w����~���� �}� ��i$nW"�ہ��.$��� ���{�Ł���ﾸW��E�������� ����nɌl�`����5�r�ʘ0N�|]y�&ў��N���2R	a���L�ѝ{v&nݗ�̼�0�1���}�������T��DKT�ʰ�����Lِ`n�t��6��_��Z��n��}���;ݺa��/ˉbU"�x�~������'߻ۀ~�5t�W+V�Y#�ׁ�������~t�7d���L��*g�a��fe������� ݓۑ0;ݺ`wV��Dt�[+��-��t�M�v^�7LU��y�p��<���l��2�6�̤�[l�U����?vn��ۦ��q`���b%��IG���i���&�_��X�7y�$���_��Q�䃕�e� ���{�Ň͞^��w������R�X�-)Wuf�kŀ^n��M���rQ�+�	@o{���%TZ��iv�3/)�ml���܉��2ގ�.%�n�Y>���m��l��0|�tʛ�V����m ���l��F�Ŝݡ�9x�u;o�;��� �v�w��X��ۀ��M#U�ժ�B�^޻ft(IG�T7߱`O���>�78�/F�𴤍�ae���q`W[�9(J&}��8�0ݙOQj�,��l� <��pݛ� ����8��'�oߖ }���b%��IGR�`{nD����GL�d��������{�{���~o�g��	��	��\��e�:��Efq�(����;�j&���l�-Xx��:�1��Hl�Ƨ�R��	*Ѯ��Ęҝ���k��SF�@r���7[�F4��fќN^�mӠ��MV/�f@���ݝq�u���s,��6[��R��!�=��oc���V���-�Itckg$�;����\�Y֒�nNx-�����I�� �@�4��3F]f�]s�ù���j������D��DF�	3��ε���%�v����+r�_@߶��� yy��J}!���;k��]E���JKe0�ۋ?��8�y{��O�x{�L�\K��ݿN[]r"J^b̦�߿cv�L߾Ke� ݑ��v&z �Nq9(}ē�n��>��� �wq`Wwn w|��5\�[WrQww8��(��������wf�� �ej�bn��,QWe����$-��C��4����D��Z�����I%y���wGLkd������%�������?���_�"RK-�Wm0���UIRK`{fA������}��Q���!%�*�� ���ݙwGLkd��̗V�����r�\�`|�~�|��� y{�p�wf����Y\�FZR�+�=�nS ����[��L�YWR��]����u6x�.�=��	�z	�zE��C�y�ǵ��-�-���TB�h����u�1��$��Ș�07�,���jr�+m�?l�y��Ēl��� ��X�u�t$�B��*�����Uj�J����=��8�Xr�J��Q|�I}
!I�;/ �W9��ڔ����2�e�`wtt�:��0=.D��������6���v[l���:��0=.D�������N�L�Z�5m�E�$F1���曩M])�Cѐ'�Ɨ��<dn,�e^f0=.D�=$�wGL��c�۱F(�rA��m���ݹ�\r6� �}� ��s��������jl���[�}��ذ/{q`�n� ��� �����k�DܲZ�X=M�� �Wt�ͻ��� P(^Z�DV��V�l����'h���V�f��=$�wGL���:�)E0��֬���)�t��w]��qPr��.USV�y�&5vh�Nl�3��ff>m���������0=.D��gZ��-)#v�,������n,��׀�v��.&Ͼ���*����+�XM�,�M�	$�\�u`�ŀ�kS#�9	,rU]��'߯�N �{� �׋�	D��X�_R�Q�䃵��k�5�v`�����~x}� ��s�~P�B�m�u�*�� l��iy�&'KQ�U���W�ӰmŮ��Kkl�ۥ�Z4[�UjU�ۜ�9�R��2�������软*�v��]��y���ŉ2�HXsZ�ur;��A����kl$C��Ͷ�Ux��v��'g%`���k�
�(;1؞��hqd�F�y�'v����5�t��"c��v�$E�a-�`��4�j-�T�$UQ�ݕ��n��n�9�j����OoJ����Y��ۇ˫���e�jR�e�w�b�;������s��|��� ����r��7-U�ݬ�׋?BJd��� ����=��Y����6i���'h���V�}��-���:`mN���EW��J����EZ��K`n�遵:5��8�~�|���𴤍�b�X���遵::`z\���d���?tS���DR읬���灺�U���G�'Q{N��0�p��{���>'?6�֜Ww7wk�5s�XΛ�g���$���߱`����#�9	,rU]� ���f�(DT�B+�� .�>g�w�}� ��n,�۱F(�r*��-]]���� ��ŇDD(S:��,ޟ|��n���d����o�u��=�np:!%
g��x�o͓��\��d�ڰ/{q`��B�ݾ����x��,�^S��`%�Y^��4����4�:��I<f�w].*.��V�\��������xl�Xg��S��r������06���ǷZ�r�Uk$�� ��۟���K�*���b�}���� {FԪb.�HݶKm���ŀuwۋ�K�Ib��'! �,X����H1#�@���U��R��F�lC���@�'�PNDn�##bxJRkȣ1�I,)F� E+FB��" mW2�.�M��>�v��0 �I#D��Z�H$�HX!��,)R�4i)
JL) �<U� S@ ~PD����D�P<��� �Ay�kf~x�n�ۻ�"UIm��V�%�_|�OwV��� �׋ ;�kS#�9	,rU]� ��v`�BP�k����ww�X����=��L����4�W=u�M��mۘ,�������z�*灶�Y�ܔ/%���}�l�7u��<��$�B�C��Հ{�_��Ie��륶S �����kŀ}-��>�g(P�L���d��-$NK�Հy{~ŀ~{�0�ۦ�{q`�u���S�KZn+eXq$��WwV��� �׋�K"�D#�0F(�x �6>�k�M�~֦�W+�V�����ۦ��遵�07nD���|���_�@l�:��V�0����S/�]�޻a�nM�&i�"f�M������ϧ���t"m(6&�'����t�ݹ�2�[SJ� ��j�:��şs�q&�z}��;�������Z�8J���������=�np��tDB����ŀy{~ŀw}u���E���^��� ��ŀy{^,����v�� �}~R��Sq�Kl�����?��(�կ�_�]Ӏ}�l�:CU���Rԫ\=�}l:��2�8��L&J�w�)�m;����;��� ��\�Μ����;���������8��g��][i�3�m��3n�������r�e��)�1�����ۨ���筃\U�\�5�	ϫ9Mmۜq��'�͵+d"��mg�m���ˎ 9�P5v�^��V}�.���!0��
����mUdس�Asŕ;.asY)�XqA4n�%����32�No
nT��GUl�@t��]%t�:\��BB���.s�,y��9U�q9,v�W�6���Lۑ0=� �ݑ� �ڸ�)S�KZn+eX{7^��t�;�ݛ�~?}ݛ�PD�T֤==��Ma��J�P�������Ň�~^߱`���o������v�d����%
��|�Z��Ss�}�l�7wcSJ�v��`]���>�-����{���k&�Ւ6�G�ŷ3vk�e���Q�k=�S�<񮭀^�䭹��N�9�\�-�]�m�ۑ0=� �ݑ�kz:`l슭�f��WYn�˹'?w;7׊�
��BI}��݋ 寱`�78Κ���Sq�IK)�w�����qa�8�M����}~0��['*��'%�1fSkz:`n܉�����]�}�`y�>R�Z���Vʰ�n��d�:`moGL��L�~�vh6nJX�z�Y�lq�M�w7�y�0h.���a�;Cx����+�����>���=��`^׋�DG���8:5>iIm�KL��ŀuwۋ �f��?wn��8ٿ}�j`�U"��^fe0:�~t�ݙJ��K{2���Z�8J���9*�Ձ���|`޾0y�X�կ�X�R"��������ِ`wtt��ގ��n��.s��},uN�qKQk���]{nf�Dg i�q�q8m/R;+E����~�6�C�Z���JYN���b�:�������2�"E��-]�e�ݬ���g(�=��8��� �׋?�a�k���VQIZVʰ�>��:np�-�ŀ4�b���*�Q��eXU����r&쎘]�����1�E�@:`�]N��L�F��-) �+�;��X脚o�_����� =��% ���v�q*OU��j�Q5^=4w
Vwk�SF��h�JE��mX����y�0�7?��$����� ;�J�	T��c���X{�L��׀w��`�^,�GBQG:�U"*�ff���,uwN�m����Xy�0���+��뮒�k�;��X�����n�$�}����=�~���4,�3e0:�����0=.D�ݓyĀI//k��)%���m���÷)mno2�]S�[+�b���Lp�u�$Ӕ�Mm3�ex�mu��!�r��cmTg��uFְv��9gl��]����5l�#�9��WM��1�:�ÑIl�B�F3��=����T�`p�K���+�'�#�9�������c��.��{ؘ����7];=�.��=�S��vy+\L�1�d�Ӄ{����޹�����3&[5��:�.u�lNv�z5Z�8��X�c�tan�=w�{�;��5�VR�8��~}���?l�07dt��q�*��1U�̫
��0=.D�ݑ���:`n̆}��6}����E�$��ex��ذ[��$�wz��=��8��U`���E]������IG�IW.��X���0=.D�ݑ� ��ʻ�w���fS�IlK�0;�:`u{ۋ =�y�]�W,VB��5�r���v��E��	���:z6�#]]߾�����,��IGU���w��� �wq`^���;ٺ����[mQ��׀{���GBJ�j�b�==�XΛ�ۻ���]��Kak�`^���?)%�=.D����oܺ�J�F^R&��Z���J#�N��Հo���py�,���X �{u�T+R�T
� ��s�~K�_��yx]߱`�w��??$���鎄g)t�*�.��]�sZ�sX2��܉t**�6s4k�:6ff,�L	�0:���6L`z^��=����Z�%��mX�����D�v�^����ŀ�S���UUw5Wdݬ ~n����?D(7���?�]TP @`����U��(�� �k���ŀo�b�;���b,�E��[q��wGL㣦�����9m�Gltv�^����?���\Q˻�����Λ�}�@�T�U&���9�,�r]�{]v<�f��:E�l#�<��Gn.ݲtģ�nE5ݩaN�I��׋ ��f��_H=�ŀv5򕔄�+eXv{^�f��7���5n�Y�dt��W2��*������o�(�3�_b�7���5�z54E�"��l�����~?}ݛ�~��ܟʿ "i 1�9Ƿ������F���-u�j�6�����ِ`v����+��-rDm�.*"�ղ曩x�����=��FQ�Lht�^ܹZ�`u�p����]	B��5k�X���Q������-���� �7� ���X���
S'mr��j�j����e0��b�:��ŀu�`��L���j*Wl���Z�X�P�V��`��p���$�K��~X�y�k�+)	bVʰ������ �7� ���X$�,��J��#���CKue�.��WL`��K�jS�j#W@A �J�`B`A�dġ �˰1At���T4��u�[H�j�*,H @a�a��E�W� �aK	)A(RA����b@aǻ�o�kZ��      ڛ\    
����Ӷ�K�g;��#X�If�n���E��i2�#Y�;l�����C�Q6��@�M��R�m&K&F���
&��#�Z���p�1F`s3�ge�Z�Wjȏeu@�g��um��5ۑ,�;i|:�Dں�B��/@*��nRZ�]�� ^�r�u������R2��(�cu��ض!�U`9T��͐���T��h�Ց�S&bEq
��N:Ľ7>Gg5�	�;����X*�*�lN���\����G/UJ��:�:�i\��re�8Իr��ٷ)�D��V� ����d��A�:�OY�X���v�s���)�d�b��3��W+�k����<c.zo5��.ga�=d)v*��m�9�Z�8*B��t�'x'c�=F��=���:�
�I�On��J��C����գV6�e���=&�\��-��D�����n�Wl��v
%
�;(�i
��0)UJ��c�8z�wi��\��q,��B�,���4��v�K!d�7od�&����%i�����]��)�j䪧D\c\�Ι1�֡�a��ChI�i�4�g`�!��U*骨��b����7g�LF�5�w[F�m簄�n��k����/[����<`�;j8۩�M. ��r�s;��ڧ���q�e��󳅋h���g'e�,�:W;��:�śT>ی�*�TD���k�a�@,�6���m�-v0�l��:�,ґ j�wi� mNEU^ڮ��Sl� ��C�5g���P���r�`BkgU�
,�gkݖ�lN�m�^�x�+�=\���:���T�q9�;x�p�1�*�h�����V� N��Th��۬����l�[@ m� H&��GAzf u���i�ѝrU�v�9�K�c�'Z�(6�&뫛��Qt��A[s[�Gi����������k��8*m@�
�h.�H�҉͈�R�D��Z �^(	�Qv ��TJ � �NTh�:\�w������[���x�N��8mN��m�flCd�i٨RMv�Φ���t,��(+�gR����vF"K&3��5�1qӠǳ���N��˫�f�`��[F䈮$-�魐��\��*�n�붧ԬE3gbvw6�6���۳�� ���idt^uIט��cn�s �$�Ԗyܻ�7mq�uZ�r��`Gϝ�{z"�`%��\��%�a2K�m.q�2�rs5��2e��n�Q;t�cn6-�y�Z�N�X���Jƥ��&5"Z�KkR¶J���m~��� ��ŀy{^/�B��$�����yuJ��ZR�Z�� �wq`]���<�ـ}�lΈIDɽ�R�Z��E]�Y�������gdِ`v��w����U ��Uv�����ـo�Ł�%
uk����U�]�#*�0`{fA����kz:`o���;��,*p��P�ʜ	yn��	9�N�i+D�m���F-J�u��5=7��{���}��9-��c������ذ��q`y�?BK�o_�إR���Uy�ff�ܓ����߁�J��~؂�(0u��k�f�kş��2���J�BX�VJ����~��0�ۋ �� /�jU(�\�v��y�0��`^׋�"v������O���Q-v�i�{۸���t��$��dZ(�k/�M	�-	�ꆽ1��R:iOa���PN��=)`A�����.\��"�\D��e��^ߝ05I-��t���U>Vfb��YyX�)��Ill�0;�t���}������eR)-e��2I��g��}����o�"��D���gvnI���n䟻��Yr�GK)�{۸���q`y�0?(P�~P�����>�إR�ݤ�[B�*�:��ŀ~��0�ۦ��q`k��k8
�IBUYcM��O]���i�6�\񛶑�t���қ�'���_7ɑ��n��+P�_�������/�8�K��ߦӑ,K�������A'蚉bX�;��ND�,K�������K5�X���˴�Kı?}��m9ı,N����Kı>>�m9ı,O����rؖ%��t�k��J�k�KL��q3��L����ND�,K����ӑ,K����]�"X�%����]�"X�%���S\��2�̹sY�ӑ,K�����ӑ,K������Kı?{=��K��/ȕȝ׷�i���&q3�����R��9-n�e�8�ı,O�{~�ND�,K��޻ND�,K��ND�,K�{�W㉜L�g}���VGLq�;��z� 83F��)4����q��3۞�E3��i�b,�Em�e����q3��L����ӑ,K��}�ND�,K�{� 9ı,O����r%�bX�{��tˬ։u�乚̻ND�,K���m9��&�X�=��ND�,K��o�m9ı,O��z�9��&�8�ſ}���T��E-�m�g�ı,O���"X�%���o�iȖ?�5Q>�����Kı;�p�r%�bX�㷺���rjk4\�kXm9ĳ����w���iȖ%�b}����iȖ%�b}�}�iȖ%�-�ӽ��"X�%�NϽ�kd�Yu��5s&ӑ,K�����ӑ,K��R=￿O�,K���p�r%�bX�{=��Kı0?��^�'��������������H�l���B<��x'�mʚ���i�J֨m��r���ۑ��0�v�Z����۶T��p{Gcv�ও�U�ړ{wf���=m����幺:�$l�#�sT��(V�����Sq 5��8�:��=�h�sq��/0��tX����􋰧.���-s�ζ���)��\`x݂����\p�3�6��ZNפȪ��$ɦv�����{{����(�5�CçU��JYy�0�s��>U+��kfUu�kQ��j[T,�~{�w���{�������iȖ%�bt�}�iȖ%�b~����r%�bX�����r%�bX����k��f]Y�.k0�r%�bX�;�p�r%�bX����6��bX�'�g�v��bX�'�w�6��bX�%�}O9��u�u��s�a��Kı?}��m9ı,O��z�9�@�,O��m9ı,N��m98���&qw�Z>�eR)m
�3��%�b~�{�iȖ%�b}�}�iȖ%�bt�}�iȖ%����o�iȖ%�b|{��t�k5I�˒�k2�9ı,O��m9ı,?�����O�,K������ND�,K��޻ND�,K��ޤɖ7.��5��ո��xzp�I!�����."�l�)��hH��nE&ݙ�g}��Ou��=�'N��6��bX�'ｿM�"X�%����]���bX�'�w�6��bY��'Ď�JBX�C�g㉜N%���o�i�!��N�n%���]�"X�%�����iȖ%�b~��p�r%�bX���}a�,�]f�\ɴ�Kı?w;��Kı>����K Rı?t�m9ı,O�{~�ND�,K�;i�2ܙ&f]k5u�iȖ%�b}�}�iȖ%�b~��p�r%�bX����6��bX�'��}v��bX�'}�j��&�D�e˚�6��bX�'���"X�%� ~����r%�bX�����r%�bX�}�p�r%�bX��{o�<cV�G�ڸ��z��y��)�۵��)͞z�[�l(�c���zm
A��6��bX�'ｿM�"X�%����]�"X�%�����"X�%���}�iȖ%�b~�;I�f�։���&\ɴ�Kı?w;��?��
j&�X�￸m9ı,O�{��ӑ,K������Kı<{��t�k5I�˒�k2�9ı,O��m9ı,O�;�ND��
�\@z���'A�n%��o�iȖ%�b{����r%�bX�w��FL��Z5��ff��r%�b�'��6��bX�'ｿM�"X�%����]�"X�%�����"X�%�~��|Hꤱ�b�N���q3��L���M�"X�%����]�"X�%�����"X�%���}ͧ"X�%�~����l+�������V%���/Y9�<������t��%�����zrgӳ�fˬ�&�f]��%�b}����r%�bX���iȖ%�b~��siȖ%�b}���ӑ,K��i�&\�&�.��.e�r%�bX���i�@"6	"~��bn	 �{^��)"sﻉ����T�K�������f]I�˭k3Xm9ı,O�{��ND�,K�g�v��bX�'��}v��bX�'{�p�r%�bX���<�˖�kY���36��bY�(EDu�����ND�,K����M�"X�%����6��bXo�� �P����׏s��Kı>�v���a�s��3.ӑ,K���o�iȖ%�bw���"X�%�ޝ��"X�%���޻ND�,K�]����^���zk�\mǌݝ9Y��Gn{v�t����1�vHͥq��w�����>�6k�.L�M��%�b{���6��bX�'zw�6��bX�'�����"X�%���ߦӑ,K���Y4d˙.��XL��ND�,K�;�ND�,K�{��ӑ,K���o�iȖ%�bw��� ���bX���u�\2k5Mf��\�iȖ%�b}�{��r%�bX����m9ı,N����Kı>>�m9ı,Jvw����d�X"Yl�/�8���.����/�X�%����6��bX�'����"X�"b}�{��r%�bX��mY��(K\r�)�_�&q3��[�}�iȖ%�b|}�p�r%�bX���z�9ı,O�{~�ND�,K�{~�����U[M�Έ;9�/i��'F��T��Cd�K����3��Z�c�����Y^�����#pq��p���q�\��qml5'cz�1i��[��ɓ�Z�T�j�vw����m�4�+��2ps�*�mړnz�5�����]����"y9�8�F�J6�3; ƫ�˺��'�1	b�lcS����M��{�P��'`�
�#
���ݽ���w�O��M	�i+�۵^d��^�c���W���S:|ᢟF�HV0̬�۵�;4j���Kı:}��ND�,K���]�"X�%���o�`��%�bX�}�p�r%�bX��O72�ֳ֭-�3Y�ӑ,K����]�"X�%���o�iȖ%�bw���"X�%���}�iȖ%�b~�;I�f�։�ɬ̙�v��bX�'ｿM�"X�%����6��b�6%���}�iȖ%�b}���ӑ,K���w�4�k5I�˒��d�r%�bX���iȖ%�b|}�p�r%�bX�{=��Kı?}��m9ı,N���FL���k5���a��Kı>>�m9ı,?�@� ����i�%�bX�w��iȖ%�bw���"X��gۭd�Fʆ�i[�&�iH�[�6Ր%�E+[x���=���sƌ-ۆ�.[,�4��h�%�6��bX�'��z�9ı,O�{~�ND�,K���m9ı,O���ND�,K�}�k�d�Yu����k.ӑ,K������9�Q���l�AF�M)�J�_� ؛�bk���"X�%�����"X�%���o�iȟ�ꦢX�ޞ����5&�.���m9ı,N���6��bX�'����"X�%���޻ND�,K��ߦӑ,K������fdɩ5�usY�ӑ,K������Kı?}��m9ı,O�{~�ND�,K��ND�,K�}�y��.�u�̗]a��Kı?}��m9ı,O�{~�ND�,K��ND�,K����ӑ��&q=�hD�\�Y�r�=Iḍ���rh.i8+�K������Ѝ����Xќ,�DYIil�8�L�g8����Kı>����Kı>>�m9ı,O�g�v��bX�'�۟2q�cV���e3����&q3���m9ı,O���ND�,K���]�"X�%���o�iȁbX�+ۿ~a+�p�T�s����&q1>>�m9ı,O�g�v��c��b��H�ѠZh�� �D�@�8��?�3J�0$�(@������$X��YHłԀQHF5RR$FVP�t�0H��-�t(h@��X1`�`�"�8�Ib�h
V!YYv�WKhE���eap��Û�l4A�HA!+)���e`��	H���ee&�WD�2�՗:�֤O~��.�qV����D�� v�"pDM��N���Q��z����N��}�ND�,K���m9ı,S��ω,))	b-D�g㉜L�q?}���r%�bX����6��bX�%���6��bX6'����"X�#8���
ZV�\�B�W�_�&q3�������Kı/�wٴ�Kı>>�m9ı,O�g�v��bX����ߤ����Z�����x��䂆u@"ꃇ< �[��Z"������Κ̺�̹���%�bX����m9ı,N��m9ı,O�g�v�)�MD�,O�����9ı,O{֛�fdɢfd�Mffm9ı,N��m9ı,O�g�v��bX�'�g�v��bX�%���6��bX�%;�S�̹u�u�����ND�,K���]�"X�%����]�"X�%�~��ͧ"X�%�ӽ��"X�%����'���Z2�%̙�˴�K���}�����Kı/{���r%�bX�;�p�r%�`|��n'w�z�9ı,N�w~�MֳT��\�Y�˴�Kı>����Kı:w���Kı?}���r%�bX�����r%�bX�}��Ք�˅���.NgK�&y�및<�,M��E�l&yGv�����*6z�@�ݪn�����{��2t�}�iȖ%�b~�=��Kı?{=��Kı>����Kħ����KemGB�KVq~8���'�����!�D�K�����ND�,K�����Kı:w���K�L�k��S�V�\�C��3����+�����ӑ,K��}�ND�,K�{�ND�,K���]�"X�%�����f�܅�ɫ�˙v��bX�'�w�6��bX�'N��6��bX�'�޻ND�,K��޻ND�,K����ɓD�ɚ�f��r%�bX�;�p�r%�bXG�����?D�,K�����ND�,K��ND�,K� ����!�D���fhֵ���5���]Ks�b�M��ƽ�s=tL�C.U�8�̮�vZ��&I6��z�lN�[�cvGb�87k�&�#]Y1�#"v�WGnܮȎ�Z��6�`���X
Q
��4B盭�A5�fm�p�<`��J�(��\pV�7J�ru�Z�Y�۳s��1�#�a�����\"{!���nm�׶�;Vx��c8�Iِ�)�������[����ettZ�"6��-�S�nEB�$�n��K��m�`"4;�:�D(5a�n�r%�bX�����iȖ%�b~�{�iȖ%�b}�}�iȖ%�bt�}Ŝ_�&q3��]�֏�Ya����nӑ,K�����ӑ,K�����ӑ,K�����ӑ,K��^��8�L�g8������K�WG,�v��bX�'{�p�r%�bX�;�p�r%�bX�k�����bX�'�g�v��bX�'��rɆL����5���a��Kı:w���Kı?}���r%�bX�����r%�bX�}�p�r%�bX��Ok�Z�S5���&a5�m9ı,O�g�v��bX�'�g�v��bX�'�w�6��bX�'N��6��bX�'�2����%2fM�E��ɺ��[W��Y�#{N|-��H�ڻW[��kA�gv3Q�������o����r%�bX�}�p�r%�bX�;�p�r%�bX���z�9ı,Ovv��3,�\̚�̹�iȖ%�b}�}�i�T@� ��SN�dK�{�ND�,K����ӑ,K�����ӑ,K������f�ɩ32j��"X�%�ӽ��"X�%����kiȖ?�
�Q5�����ND�,K�����Kı)���ne�uf�2]��iȖ%�b}�{��r%�bX�����r%�bX���iȖ%�bt�}�iȖ%�b~�;C�XEd���l�/�8���.�~��9ı,N����Kı:w���Kı>׽�m9ı,O��������(]B�m��%�@����Ͷ�D�Ξ�<�mٺ�υ����˴�Kı;�{�ӑ,K�����ӑ,K��^����UB~���%���]�"X�%������&:�2�]fd���6��bX�'N��6���uQ,N����[ND�,K�����ND�,K���m9ı,K����%P����j%�8�L�g8�>���r%�bX�����r%��� ���Ț����"X�%��{�q~8���&q=��VҶJ�-%�iȖ%�b~�{�iȖ%�bw���"X�%�ӽ��"X�%����kiȖ%�b{������ɫ�˙v��bX�'{�p�r%�bX=;�p�r%�bX���z�9ı,O��z�9ı,O����_�L2�5-"q�$���oR&��:%=�Gr4qs]X��ȇ3��"���v�+M�^����d�<{��6��bX�'�޻ND�,K��޻ND�,K��ND�,K����\�WW3%�WXm9ı,O�g�v��bX�'�g�v��bX�'�w�6��bX�'N��6��b���.��G�,���Iil�8�L�bX�����r%�bX�}�p�r%�bX�;�p�r%�bX���z�9ı,O�w~�MֳT��\�Y�˴�K���������Kı<{��6��bX�%����ND�,�O��T������{=��r%�bX���L�uu��33Xm9ı,N��m9ı,?�:���ٴ�ı,O�����9ı,O��m9ı�{��}���=w@�Yi'VE�K�n�M ���=��n�
�vJ�o����o��kjf��W$�&���%�b}�{�[ND�,K��޻ND�,K�{�ND�,K�{�ND�,K���32e�Yu���5���"X�%����]�"X�%�����"X�%�ӽ��"X�%��]ﵴ�Kı=��{�ɆB�d��e̻ND�,K�{�ND�,K�{�ND�� j&�}�{�[ND�,K�����ND�,K�i�3Xd�5�sZ��ND�,K�{�ND�,K���kiȖ%�b~�{�iȖ%�b~�}�iȖ%�bS��<�˖���d�j��"X�%��]ﵴ�KİP?{=��Kı?w���Kı:w���Kı?�v�����5�fd�������r��y�v*���z蚳��V\]s����*������.��ظ*4g:F�@=g�l�L�s����>O���8sjp� 7Ag�hw�w!����<ݴvnJ�ݺ�#�@���m��3�..�5md#j�͊�e1-C
m�E��Vvӭ���\XƸE��cC��l��gDu��	o[W8�t:�!��
��`�i`�u�fk+q��I\<��@v��� �M�ޫ����K�\ey{��N״�x�-�O��,K���3���r%�bX���p�r%�bX�;�p�r%�bX����[ND�,K��ߋ�kY�fjjf�Y�iȖ%�b~�}�iȢ%�bt�}�iȖ%�b~�{�m9ı,O��z�9ı,O��Sə.���ffk�"X�%�ӽ��"X�%��]ﵴ�Kı?{=��Kı?w�~Y���g8���ZB��,�j��6��bX�'�w��ӑ,K�����ӑ,K�����ӑ,K�{�ND�,K����d�f��5	r˙��"X�%����]�"X�%�����"X�%�ӽ��"X�%��]ﵴ�Kı/~�v�^ɖ��c�0��v��g�<�e����ڣ�4H�%�lL�4�[��N�k�_�߉��bX���p�r%�bX�;�p�r%�bX����[yı,O��z�9�L�g�������%�Il�8�N%�bt�}�i�D?�?+��q7�����ӑ,K��s��iȖ%�b~�}�iȖ%�bS��<\���.�fK����r%�bX���siȖ%�b~�{�iȖ*%�b~�}�iȖ%�bt�}�iȖ%�b~�;I�f�SVf�5�ֳiȖ%�Q>�����r%�bX�{��6��bX�'N��6��bX�'��m9ı,O���y��j�����5�v��bX�'�w�6��bX�'N��6��bX�'��m9ı,O��z�9ı,Ok�z�2��'VX��ܨp����K,&�������4�,TU^��{���>���[�vӑ,K�����ӑ,K����ͧ"X�%����]��`�'�wج./|}~%V;-�W�KV. D���q=ı?{=��Kı>����Kı:w���,KĿ}�k�2٬��B\���ND�,K��޻ND�,K��ND�����H��h�Q8 /��b~�����"X�%�~�}�ND�,Kݝ��	���ɫ�˙v��bX�'�w�6��bX�'N��6��bX�%����ND�,U�?{=��Kı;��o��4Mf\ֳ5�ӑ,K�����ӑ,KĿ���iȖ%�b~�{�iȖ%�b}�}�iȆ��oq����p<�V�G'�N�*/:K�۩ e$蛧6sg�r[=��F1�`�N��5�����p��ND�,K���ͧ"X�%����]�"X�%�����"X�%�ӽ��"X�%����G�,����XYnq~8���&qw���iȊX�%�����"X�%�ӽ��"X�%�}�fӑ,K���;g��\�fML̻̚ND�,K��ND�,K�{�ND�,K���ͧ"X�%����]�"X�%����O8ff���f�̺�iȖ%��'N��6��bX�%����ND�,K��޻ND�,��E�n%>�吾!I
HRB���U�]]U+��k0�r%�bX����m9ı,O��z�9ı,O��m9ı,N��m9ı,O��_I�^�32�V�\�a3q,���z����7<ݱ��@Mų�Ź�a��qU�������D����ӑ,K�����ӑ,K������yı,K��{6��bX�'���kЙ0�\̚��̻ND�,K��ND�,K�{�ND�,K���ͧ"X�%����]�"X�%����~f�ɢk2浙�6��bX�'N��6��bX�%����ND�@lK��޻ND�,K��NDg8�����|�vV�h�U�_��,K���ͧ"X�%����]�"X�%�����"X�%�ӽ��&q3��]�֏�Yae,�����ı,O��z�9ı,O��m9ı,N��m9ı,K��{6��bX�'N��H�#`@�U�|��£7>�ݤB�iX`XQ�RQ�X�R��@`�#�p����ߔ�u�6�5�.�:�!©�4 <1e+4J�0q�R�-�a*�i�H�+4�P��j[�)(A2��4i�"�!Q�@���H��4%�ZQH�yEpWY�`J�����������#m�      �mp    �d䤶&��fmm3��v�!r+l��I��gv* �[���K����Nvݶhn��l� I#t�J�9����sl�&�]%�g��-ڞݢ�8��w���2��G���f����N�+R^��1m�a��4��ZeV�Vΰ�J�,�5UUG3�x�f;H6��h�I`]LTq�ۄ�]*�c�'lR��g�\�+TTKY�n�jx�ү]��ñ\
�]=N���n�\�t��R5J�l�P��eRgm�;m&��M��tR4lA��蔹orb�rey�9 8{��dʀ��nv�WX�uc
7cҔ]J�mt\ulSJ]6��\���AZnY@�
E����$�e�o9�m	�l�n�F�����S�5)���7}�I\��GkKm/.Y���ѻ��[�n\�v]�L��R�Q�m��V��p�v$�ݑ���Ɗ$�	�=a�N�=yp=BS��g�%*��\C�F� UR��mU���x�5��]�EQ	� �N�m��ɻ[��"	��p����v3ħ&�<DĊ��Um�ٺ{n(Z2ʪҪ�䨮��ĥvQ���vV�nv|�f��;����Ql�f���bt��v��kHOn��۵.�=�Jo`m�k����I�g��R��cj���v�ݎ�y��x.m]^[��f�2�u�2���ֻ ܲn��v�[3n����45�rL	-6����6Q%Hi����\ݵۃ�Ƚ��J�I��^����ni�C�&,|�8H���ˉ2�Y'e�	غVh����mF�zI6�|�u��|&�)���fP�cn+l&ᚶ����nGPY��Db6N�h�(T݁m��ȩ�Ra 1���G2��8G3�vܺv� �:�)��n�  �` �:M�53�6���t��6���M��N��/N��q�f��Lڡ�R��u%vq�AWh�۹�� AC±:{���wy�EJ��B(��^����!�E ���P�U���UM����٣Z�����Y�\���8'���D���u�SIz�i�F��� ӓ�x8��1y�����^cs��]m���vV��stii1�����vN^�63r��]��b����;{+��G���j��? ���Ş-�	�a��Lu��e�LO	)��43rW#]�r7l�^A�+�sE�E1�l&ɲK��15�����;u�5�s�o'ﻻ����~_O�'\�E=5ٺ���\��Y�B�ѱ	�4��Q%"�]�l�W��{��y���J+i	k�����g8������m9ı,N��m9ı,K��{6��bX�'�g�v��bX�'��&�T-���v�Vq~8���&p����Ӑ���j%�~���m9ı,O�����9ı,O��m9�qP�8�����K�c�*�Z�j�r%�bX���fӑ,K�����ӑ,���j'{��ND�,Kǽ��iȖ%�bS�k�Jk.�P�����Kı?{=��Kı>����Kı:w���K�,K��{6��bX�'���k��a���5sY�v��bX�'�w�6��bX��|{�ߍ��%�b_����ND�,K��޻ND�,K��I=SvJ�L�\ܼ��:g��r��:�:|ᢞ��
��7�u���w��Kı:w���Kı/���r%�bX�����r%�bX�}�p�r%�bX���}L.\�[�W3&Z�iȖ%�b_�{ٴ�?���TW��yQ,Mw��iȖ%�b}��p�r%�bX�{�6���������/m�����;)%���㉜,K�����r%�bX�}�p�r%�bX�{�6��bX�%����ND�,K���u�Y̚��.�m9ĳ��w���m9ı,N�����Kı/���r%�bX�}��m?L�g8��5�m�7m��ʳ�"X�%�����iȖ%�b_�{ٴ�Kı>����r%�bX�w���Kı;��rkچ۫2e�Yi��y�z��beZ�ĭ��p�-�c�4am��.-�Ht��-w�w���oq�����ٴ�Kı>����r%�bX�w���Kı>>��m9ı,Jw�CZ�ˬ�%��fm9ı,O���6��bX�'��m9ı,O���ND�,K�｛ND�,K�kY��UD�p�S8�L�g8��}�iȖ%�b|}�p�r%����J�@�(~�"~�{��ͧ"X�%����M�"X�%��{ڧ1��&��˖�a��K��j'N�~6��bX�%���ٴ�Kı?{=��Kı>�}�iȖ%�b_ӽ�0�sYnY�̚.��ӑ,KĿ��fӑ,K��c�������Kı;�p�r%�bX�;�p�r%�bY���Ј��b�X����	�28�)e�ݩ��ڌT������N�#����a5�Z�L�fӑ,K�����ӑ,K�����"X�%�ӽ��"X�%�w�ͧ"X�%���v�:֦S3&�s5�˴�Kı>�}�i� D�Kǽ��iȖ%�b_����ND�,K��޻ND�,Kｲ�2L��չ�����6��bX�'N��6��bX�%��{6��bؖ'�g�v��bX�'��m9ı,O�=�e����������{���w{w95����iȖ%�b}����iȖ%�b}���ӑ,K�P��������?����r%�bX����ֿ���]f�.33iȖ%�b~�{�iȒB���|��)&Zo�`�u��hc}��Ց����dN׀Ѹ`��"�Ge0�^�5ES��{=4ru[�Y�������:`�1��r&�v5����%�7mX�����.%2}׀{��pn�Y�L���U�d�d��9*���\��ׇ�9�$߷~ŀj��������,���ˌK�07�:`uwGL�&07�3y$+V�Gl������?��߿/�}׀{�ـ~Y�j�=�UWww`Y"]2��Cv�j�bꭖ�9�I���4뤺��jݗ��
�b�K-������Mڵ�mS�8��u�]q��g풛��.a��ua �ri˰窜jٺ�{yT��ۣt	[h��=Vທ����ϛ�E�7k,���O]�v��C@�N9�y.�u��v�˛vp�v�2;9�{㺵�zvy]:�h:gi��'d&e�f�-��O�Aڊmd�jM�:��\��ɞ&y�벙�ܖf��"ݎ�A��\��i�M����ͮ�`��b����>t���x�i�I/%��Y(U%� ?{v���ߧ�8�ذ[� -�SVJ�����fc��L]�� �I��ͭ��D�r�k�;�n,V�ŀ�����_t��T��*Ք�ZY�L���n���Șٸ��7P��Z���k���nUV�iE(��TI��.�{�1�`"4Z�ł�k3�w��7zc��Ll��^���?zy�xY\e���� �����"Bq	/�c��b�9w~ŀ���;��3y$+V�Gl���wq`]�� ��K�0=& �����,��������}���׀|��>��Xtۤ���d,�*�Հ���"`{dt��j�*\Y�j����N�^��IO,tX��]{Nzi�x��hZ��ppR�V�v����n���ŀj�x�~^��׀~�_��V�0�y�10=�:`uwGLw���n���Ʋ�R"�V� պ�`�����%	�Q�D$�$�LDD/DDz�W�8�� -�)�d�2��:��`7�o� �������/{q`�<Ѽ,�2�Kl,� ��{��Wtt�=�cvJj�.n��LM��u͡j�QI�]f�މ���sE��/<��g��z�|�-XJZ^�����0t����vcT���v�JYV��n, ��ۀ~ٺ��ۋ �t��:셒�UWk >�� ��s�Dηذ�v, ^�mjWl`� ��׀w��`��X �H��B�$��K��ݸ���BK\� ��ŀj��`���t���(Is������6ug����K����p����X�s6��K�ѣ;d��{���ɑwe�������X��x�78�ۋ ��k(�amRJ���q���L]#�����/e���e�vn������z��`w����f�I[���K^�����t�=�ceȘ�Lv�m���`^�ŀ��p�78�^,��!~J!�!$
H��������!5S�k��V��ma`
�z�X����[;=��nT������r�׵���4dh0��t1Y1�\���W&�� ]zw6΍ؓtcu)L�z x%,n�lӱ�l�lZ�*l�<�.�f��Ȟ��#J*���������|5qs�v�[�5�^�%�N�TM��Yô�[��g�`���C���/���}q[+(B��6x�v�8�l�{���{����@���f����u�2kZ�LudP�NN���h��y����1���L��J}��d����\,�*��������ٺ��ۋ ���, ^�mjWla7wx�79�S&�ذ�v, �[��;���V��e�W�{w�XWH�{��ˑ0:Ij�|^VFf�fS��t�=�ceȘ}_?n��`����Gh�h�U����?%��?��,V�� ���d�\c=$���]Da��de�MZ���rm��k�w=p� ۲�k�a�KQW��:\0n��vV =�����n��eճY�Y�rO�}ݛ���R���IG�"E��� k�x��y�\l���>�������T��� �I��"`ott��L��}vB�B�mX�۷ ��׀w��X��q`�tSh�R�`�m��78DD%����}ذ�n�����l%�R�p���jV9��]��V5ǕK\4�n�L;0-fƫ����9�y��07�:`ut���L`l��ݍe�*�E���V���X��x�78�^,䒈����\�2B�Tܫ ;�}p��x~��s�EƆ����i:�I$��@8D�Њ���!>HY�4�x!�X�n-�,H�0H@H��$���c
A�@�T!B �5�H��$#R$�U�XaVHE�B4	d�5v�����a%B RXX�!# X��B!H$��>�j
H1"V����8���T$J�f� Z����IBT��Q���MM:h���$�`@���a
��i2�BKQ��� ��@���!E�D)H$� �F&�U;.�CB�օ:��$X�a������x�����L������ڌ�?& �4D? ~A^ -_�ZT���/�4�W�
��! @�AD$
"�A�@JhX �(IG�(���nb�m��>[[(p\��K]���$��~����=��,��t�=�c�m�'��-f+H��ws�{u��?D&�w��>��<��o����v�<C=Iqu�'l��u̗M�6��YI�cvM;m/����ٽ+0�2�]#��.D�����6�%�u�%
��`�n�Λ���,V��?(�СU��*�EZ��xX;m�7�<��ŀy{w w۷ ?wZ�u:Զ����kx�Z�, ��x�BHJ�@ �
���ﹿ]�9ｪo��m+rՀy{w��O�����}��;��X��qFբ�87lh�vz/5�;(Z4��k=�s�U�)u�>U�����j�Wh�iSr� �nݛ� ޑ���t����D��˱e�3�]�t��DB�5�b�}ذ�����q.6w��ϸܲZ�d��^���WH�oI��"`n�As�Y�X�3�fS��t�7��ˑ`t(Q��߿y`uqU�*nn���
�řLzL`l�zGL����s��7��m�Y���mpp��1�4��'m�Ѥ���ІWV3M]C2�;Ilp�Z<��m�.D��
MB�P�S�P����0�T{I�kd$�U������S0@oO]*�q��@v�76�3���[p����@�2	�e�׮[tWc-����v�ě�Ǟ��A�Y�㶝�ÃuX���R�1���̘��[P$馊���&�z&��ߟ{�\[�%��]'������*�WT�ٸ�{t�c��o(��cpz� &��ط5�:W]�`��;�O��w۸�/n���v���]:�j[BK\� ����Jdi�b�5�t�t��۩Y|%T�m#rՀy{w�Mׇ�K�7��<��ذ��kU�v����%yL�06\���#��T�����٭p��Y
[m��ٺ��u���t�޹ ��s)Y�2����v�򓐹�U��Bb6���.Z�\���U��ʘ��,e��^�n��:�GL�06\���1ϱf%b��5����w�7�P:TN�PGb��t@�����ܓ�k޻�s��XW��7���vJ��X��j`l������t�+w���b�ŋ>2�^b`l������t����x����-�֭��W�~�XCO����}8�78��ddn٭���sr��ә����ML�Âl���wX{e!X� )���gj�w�]#���L�"`ott�<wD�(�am*nU�~��xvn�����<���>M�[5��Y!Km�eܓ�k޻�~�����ڨ�DC��P��9Ӿ���=�}۹'��ΦIk���mr׀w��X��q`�7^ݛ� �v����nڬ��`��X��~z�� ��ŀ7�u�~.:��@��a�� ������7k��sŬq`���My,��	&�9X�)��T���0:�GL{�)5Q�Y/��^׻� ｸ�/n��?zn��6��}Un��W3fe�:OΘ]#���Lm�ۻ��UH�7mXW}����k���s��۹1�<��`DQ# #�P���g����ݥN�hʥ���V��u��.o�>��}�� ���, ��D��b�[yum��͐]Y��r�Sv�x�p�A=H��y���j:��E�e����+�?wn��GL�����ȟZ�Y�yh̬W�{����t��\���L�6{�V�WkpvR�[V�����s��L�z��5�ŀ|�L�qn�e��Wj�?zn��v�w��X?/oߖ -��F�d�v;-x�v��$���|�}� �i��-%�$����slRKm��!��hR�vغ{g�[L�k��3��Ц�ʗQZ�n��[&�a/S�y;��N�tq�7U��l��$mț�SKz��c{�IӺ�`��m�NJV�|�|��Gu�I7���I�+�&�tz�u�)p)�����n,� c]�냶���cc����6��ֳK�]�����6�[���ً/�vM�t�А�ɋ��lg�ٱ��{��r�QG �O�n�ƙ?j�WYs����'k��s6�9tV�
r���DW#u��[[U�Z��e���߱`]���>�n�}!��� o��e�V�������`moGLuȘِ`otu��`��k��v���I���>��>�a�)�o�`��,嵲��B�R�l� �ݺ`����n,����?tD�7��[e���Lۯ�j��/����>�`���\���+���3ř2���rY�gt��^V���\��a��j�&������x�����7?�(��5�ذ/���(�v7mC��V��v�B��:`�P�T�P��!-��IB_|o�ـk׋ ��n, ^�MTjVZ'c�׀o���=��a�DL�}ذ:� ��S��U�Z�Ў�^�{q`��� ������nȲ�R���Vս0=�"`zvA�����r�@�$rZ��m��	�Vp%U't�W7]��e�����<��8���U*���u�8�npn�XZ�,���F��Y
[m�����������r&������33(-T���׋ k[ń�%�!%j�A��"U| '?�������l�����E]���q^yL	]#���L	�"a�_.��� ��i>���cv�:��`�7[uȘ�0%t��j�*\Y�ef���q�ٜ�0tj�0�q!�={L^�n���L_߻��N��佖9+V/��/������+�t��\��n�m
Yj�A�ex}�şɳ�}� �Ͼx�n�ۻ��UH�7wk k[ŀ}�����y�t��b��ֵ:ݥ��i"�U��9ė�%���N�����=��`W�P��RJ"��J#]ذN�Q�]]QuE�w�x��D����+�t��\����������n�pLMȚ�7ʻ^vbI�t�	}��c����6�Sӵ�*ǳ ��\��x���X�M�/�BIz������������[��U�j��Y�DL�u�8:�ۯrQ
d�&��(�n�ڇUv��>�����0%t��n®�`��X,����В����N�� ַ��}~��}�_P��֭��W�{��`�9>�/���7ջ8�!$���ڀ���� ��� ��AW�A_�U�U� ���E�$Q(�T 	E��Q(�B�DX"�b�A`�DX*$!E��T �0DX��Eb � E���`�0DX Q"E�E�,QE�DX�$QAb�DXD(DX�DX(B 1DX�A`�@*Eb�E�1B �DXT"$"�P���bA`D�aT! T AdAP�X
��*���*�� ��@AU��
� AW��_�PU�@AU��AW�� ��� ��� �����
�2��w��,?�@���9�>�|� P        
         >�  �  J �ER��DU(H ((PE   �T�"��@ @J    ��*��  @� �HR��@���i�i �� ("  ��@�_[qg*㻟g^����{�^x �-�����ξ  �7��}㷍_<P=)��oKŞ���{��i�$(x���j�ܝQ�J��W��<� "  �̀w����:��u��Δɩ{�*�;ϥ�t�q۩��8�Kܩ n��zuqܾ˟}�S�U_=� ^�R�>쫌�֮-ULl*�� ��Ub�W�����q�P��;�>� $(� @͂�y�qo��o�ۋ+���[�����)��L���x��W�Pn��.]iɯ� �}���o}n�Y����{���ݚ��u�x�S� =8�}�^�*����wo�{�T��׶� �� �  �@c0 ;�i^�ϯ�O=zyi�O����� ���Î�q��Κ�ۯm|�P��K�����8����&�o}�h����v�N�zy4������y�@�o=}m�n�w��}��ivr�K���TP�*�TT��3` <�R��}����;�v�y� ���  
D %(� 0� @ D   @ "
 �@ ��  9�  �UCH Q���&� 1)@   z��iR�=L� �"������J�  �=U*�C@  ��UIR�  �*����کJ����d�aM�R�G��b2l��P������g���?�|�S33)ӷ�!۷��H�*�?�PUt*"����*���*��"���Q��Z����ҢiMGT_efX��{>����B Aia?���D�ID�����'�Z� T4#�
�*��0�$ ц��f��ѫ	�)�nؐč�!F� ER#��CD
�X�i�) ��#&�PA�4I
��� +�D�Y�c9�I5MGz�5"
�HCk,�+D
�H��Xm�� H�Ȼ$: VI�B1��M:0�GP�!f�$�H�ԁ�&�Jk�W�L7Ōu	
F�F�j�/T
;��?oW�߳�h��7���>4|��	+IbIÈ���^�H^}&:QI8�$V$k��6|j1���I ��5oŒ��$�J�.~�?ne>�I���|�'Ѭa����!?�����|i�H`^S�N
�%b���(�SFd�?��4���~�����J��k7���HWG�����B�7��k��_�\aV$Y$+
HŢ��!E�-�����!a�X�"@�H���:I�DӢ1�Z�>�N!B�sZ�֝0��߹~������߳_Q��:#]ֳa���M�@�|�,a�0���BHp�8<6D�!F^C�Ghp8���1��p9��`A�xh1#����i
jD�ǄX�n����8�f1v��GD0�ǃ���ӌ7��,)4C66��0�>5�ḧ#��EH�j�D5)��]���,%���ٓ5�!u�0�Ͳ�6��� ԅ�	u��t\)��RRS0��v`��̔�����m�����!��k5bRf�M�\�7�e4`B���Y3{��Fd����Jk�i!M?�Ą�0�� @� J$
|�� Dz!����p#aN0��JWI���$$"Y�`Wc���6`�I!SX W$�!u$
d�l�,���0��U�b�WK��H@��Fp�$������Y8�ރDѭ܆��!���!CI�$�!WK�F��$M�$�(h�26ۢ2פ8'r�!f�s YbP �Yы�������CS��	��X?I"@#�$0�6����p��K!�Z�B��9!	].;!NL��i�7�!�p0v$�.�����B��b��$H�
�p�h��~G@h$�٪K�p��CK�D�	��q$l&�$�HBI��,��F24C�#�]0H1���YHAtI�kaQ���Ɛ�jH�d�P���BP�]�C����l�~0�F2�H.�L��m?B���0M�$�a�S�ߠo�`@v$ ��A��Y+J�� 41���Ii$�� H�j� @���H'���!8�B���M8�(h�!��$'ք`H�bB���h��#)���7���ǅ� ����#]k��?������ XF��BD�GD"&�H�u 0+��A�JA�d
���b�W!W5o�摆8Cs�b� mH
��]E)� F� ڄk��HF��a��VCF6E!
��#"�`[��D������M�
�)�$�D�4a�&�H%�Forp�H�Y�H!
k6�"WY!�&�$l��gp$�*h�Ȇǌl�_߷���ֺ�C�&�<n��C����ۚ;���Z��y���HUx��a��A�%��]��$	�����Ap)��;	1�5�.ĩ��{]1ba��XH���Ő�F�jl�i]&j$C��������4}Nw??�������qS�,Z�r�o�s9���]81�i�Qt�B�h\R	��� @�b��d�) �~OɸN=v;��8��#j�,��b����E8�k��	��"Y06p8*h�g$X�у��)����!�?~�>�0�� ���NP٬$4�1���VЖ��D�+�������} º>vכ�4ou5�e����� WN(�Dç{����ֻ��4h:�e�)����w�p��� 3��L1"�R0Xt3S\�q �N? 6��� T�ͺ2���lX�N0����kS	�O�[&����!]��SI�i���&�d�9B���,� �YJd�`P��`�v����f���Y17�0�Cb��
10ZD�D�Q��"��X�� �! TI���`SF!r�	!!R���HP�	1aCA�
f�$�CNB���R4c��@(D(��v���	��8�3{�	9iɕ�@�Cu���G�l��MP�^�.��XO�!e�?sNH�a��&�_�!FZ[(���P`��N��?"P�8 ?$jh�06B'}34l6 �t�v	��]8od.nC�P4�4&���$H�$�"8\9Ɛ6h-�7]���5)	��#d�?�!��fHl�`E�!Q!���SF�zad�5���2Hńa �)&��WD�
~�f����7��H�5t$�YD�����z,i��A����a��2�����FW" ���s�D�R&�"�A���
i�o	��|�{?H%#�"�X��4X,F�������і�Ϧ|������Ā�Lʹ��8�HS���ͩ !�,H*�"�RT���� �"1?&�$$X���5�����АR�� Ґ���� �b@�$	HF,�F�f�J�I��9@�"F��Yu�.���a��!�D���bAH��X���@#YT�@�
~y������
1u] E�F��f��;�D�#����V+% �bĉ0��
�b�D�d���� �M��
�$5���A�7F� ��X�jl�s���6p�H���� �����YVk�.���
� h5 �]�$��)f�F:��OƗ�M����b� A�� @(F$H�)6 �P���H���hWE����k
I�4��U�0�g7���ʹ���i�������X��!>&#3Of,�`�b��푶�I$   ��                     @                                               ��                 ?�>                                                             |         6��҅*��-R�0�ͭ`� ��I�5� o@� 6ٴ�]6    -�/�۶��m��� �٥����8!m[[l�0(  ���`�  p[@  $  ��  �`[���z�8m6�  �q�� m����]68 p:N 	��*�R�-��m��6Z ��$��n����mH��n[Rp�lf�[@k�:	05�-��$�      ��>�    �i�  iͦ�� ;m�6�� ګb�pT��UUmT� ��ݲC��� �@�-:(�b��P
m�m%� ��V�,ݫ��p   �UFBZ������ m��D���$����i[�H 6� N�/-Ѭ�Mֲ�:�@t�r��٪M� ��ym��l�v�i $��5�.2h�\ p�ղf� m[^miD�D�[��� � ���Hrʀ��ک
V�Atq ���η��A� -�m��	 � ���on��umbe٪��jU�@5M�YЄ�v0�@-�Tp+v�ܰ��  8�� E�am�-`5^����v�[o�@q������U�`%`�����e� [է5��^k:[�eUXЭ/-UT�t�I*V��-� ���:@� Zl� �&ԫ�Yi�-U.��W8���Vݶ�Yն�   6�^�@ִ�,�]�g6��&���	~[����m�v�`9m�    6��if��qm�	�Pcl+++Ulim���m����� �m|���UeN{u��	 (t�dHB�TaAપ$ z-����W�N@R�Tjh��:�nT��Ggyf���.�6����T�t�9c��V�&�l� 6� 8m-��z�h�6ݴ�XP6��Hl�YA4�UWOh]�i8u�Nh���@[b����v�k�E�W���m�;l[NR�hH���ml� [@͖�;4l!�� �f8��r@�k �[tŷ`h�n@�X` �uԠ-�m��2�m�d�kn &�6�pV� �`:A�l�k�`H�z���A 0m��8�UԂ���d@���8d�mm ְ��.j�:U�V2���Kh�$�-�^����G /[\$#��*�!�+�j��PmT�*^�j��UU�W��쿚�|�	+l�� U,q*��YNj���
�:���V�ԯ<ʭ����*���qokpdYv�m�@$pI�l�qv�m"�-��@pH�
�� �p$� ��]0[E��S�V����AI$6�Tb�@j��*fi�Z��kX $	��%[�47�  �� u�     M�m�j� � Gk� [@*� �@UT]uT��-��    n�-���  ��/��  �t��w�o]g!�ɥ�)[k�ݵ�s���`���-�uĀ�[
$m��ղmp�����v �m��9o[o7,�0  5�6�`mUn��kp  ��p �I��kl�	���͛�l��۳m�� �%&�H3e����r�{Z�@�m�h ��t�`m�l�*کX)U٫��{�*�h
�U��j�]�@m�lp����(>�kgY~�.�5�2��Җ�u���Ͷ�6�
�T A
�@����l[@��$��lٻ` i� ڷa����mخ�i:��M�  m� -�;m��8�6�v�5궭a�|  �6�d�����ht�h ���ۀZl�vv�I���6� n�$����V���[m� 6��m���[{�q��}���-�Бm �h	�m���pmsm�NkXݖ� p n���\�  I �� $� m� @8� m�09 I  ��m�`Hhm�0�_����` $ �`  l@�Ãm�m�l���[n�   ��Ԡ[Cm�$   8 �i�m��(m�E ���i$�\�具9m �7m� � -���k� �HV�ޠ6�"�ݶݭ�4	�ݭ����ـ�ۀ������mk���p$��H��o��� "ʻn�]u*�+UJ��1���V��"Ll�D�c�We'�ݪ�βͧM���[��V� �W�Z�iV��usI��h[���[�e����nIm6��p6Ω )kn�h�᪕@�K�5Ԯ�� U�¯��꧕�UMMP	geRW6��d�����n������;lu�4�,�W\��̪���s0M�m F��f�b6���6ܩ.���{���n$mm���]m $  �M����`�iei5Ԑ�.ĩ����U[Kh[@ ��Z�m���^������H��� 6�$	�M�iJ�T���ƴ�kd H� -� kXp�I�[G֍)��k �a����ݤ�U*�J�@UU*��AlҋY- �`   ���u���6�*�*ʵ�U!*KTm@�`���p�]$� 	g�u���   l��Kf$�6٪�kiI٪���i�*�JH
�UUT�UPjۀ �f�   F�mk����#�@�ak���[)�6�-��:���l�lH   [zp���n�il�m `��Mn�(�Tu�l8�6��   m�m� $��t��m��M�kl  ZĀ7J��[@��   �m���&�m̀�ku�ݶ�f�Á"��h��`h �i   -�pj��8�6Ͱ �I�-�X`�v�m+��0$ڼ���Ѿ�~�|  j@$ p8    N���m�)��U<�q�<:�[]JZi0m� ���Kh6�  ��    	l �       m�$kX ���  Tݻq�N��;`���  H�����  -�       �h hl�-�^�  H$�[�-���m���mpd�P� 
��R@Un٩��-���� ���U���l�ְ �Ӡ,`$)���U�1R�J��8���X m�0` 6�  �8'@4P	�V�čm�i� ���� p  �    �  ڶ�`H;Z�� l Ӈ��[V�ڶ�m #m�	.�ܶ��d�"i�h,��$  �Q   8�{l �ְ p��e�aI�6�  m�  ��!��hhm�i -��� �m� M�@m�  mj��[Amh�kn��X�     m�   -���i �$�i���l �/i��� �lm       �  Y�  [@��W"����&�c,�@ ��$   �m�պ��$V�$m�� ��T,��R�`��h`�@   � �Ͷ�ﾓ}���i�� �[@  2s��m�[@^����QxH8j�I@9��H6���7m��� Hi"�-���[�	  �kJ��-�x۳��
jj���78�v`)�`�������1�2�8���C�ĥք���x9{U(]�J)v��GZ���=;-!=u���;����'jz�;;;���-r8- �̪�m���Z�F�$��:۶ͤ�5u�ڑnM"(��2+�*UUW<���,q%�텶KM� X`�-�[@�|4k����)���`   M� 6YV�U�^U��i	��   �� 8&մ��J\�K���1v0� h�@Zma�m m�� m&  �l(8�c��km��-���m�m� x[׃l��k�    �m� mi�@mٶ �f�8 �f�ۙ�������*"���?�?� !�����E@:L��QC���`�vU����Qq  UT'ؘ-!$,�a$H� ��Z
��T�cTU4��Q0�*P�S�@��:
	�.���( q@���Qn�b��M 0@
��8 ��E �G��@J����O����x+�$� `H2B"	F�C���J�(�Q�(� M�AF.|�ਘ�΂t�h@�j�m"�0��/G���*#�?|�J���?(����
&��(uPG`~ "��sb	�(�DN� b��⫡�$\ �
�? �_��@�	�!W�P�e`�@E�S���k_���   �        �l  k           m� -�k.�rU� ٪��S.�&Ia�Y�2�:��q�ח6p��.�x��]�h��n���p���n�c4��
۝�.4�Z�-Eu{m�݂汉�g6�i��((��� �ە܇cN�!2�4� Z,��:y]���3�V�O��A�@y��ke@dt�[v�2��y����U��@YZ�H{;n�)T��H�Z!b�JH9wJ�u��C�e(����NӁ��6�T�,Vq4�Un�֕{,�<�P�n���
���l��{Y��ru��m��� GY�q4��=-[D,al��1l��`v�-qm��gM���:C��Y�ɤUڕh�u�t�/Y�W%6 �ͳp,ݥ^�,bR���e�/FØV�GH9��D���Q����\�1:C$�/Aiq��֓����{l%�� 4��Mf�Iˌ���4i ���ӌ*v�f�v��,�h�kM�T1�nH9�t��P��pu���M��cX�{ojo�F"�����d��'-��Bq��t�q��-����+��f��c1�����R�l��X�ݙ��X��D�61 �7Cfx�VvZ�-�yL�R�mr��U=.K:�V���mW6 RɜcM�L�3>^���5��v*\&:v��ꕊs@K�7&Ӳl��YC]�b��ѥ������#{q:�IiV��VW�*ɑ��-��ac�^��&3E�Q;ruLR��R��gH*ۭهkm�p���z-���f� K� �<�[)��6��`[j�S��IAJ��@ț��\e�s�KvWj�mz��k*�3w�-���۵�q�ۍc�Ym,��{(ڜ�ֹЖ��Y l�yضQ�W2��K]=�V�	/*[Se��M��c�;V��$��S�w{���Ҩ����	�T4���>�{��w��}������À ]62�UUU)�3s� 'h1��q�wY�/G6Z�*�Fy�	^:tS����'A��I�m��ܯun�ytG%�y4�bN��Ғ�:j*�Sr�k2�Y�9��y���vMiBҁb���SՋ�t������S�ݖ�t�L`��*ݲ���2�����ݡ�����j.{FN�S*�����՞�i3R�K��W52IfE@Ё�`N=���(�]���W��=�odM�ێ7!��#�ۭӢR�5N��3x����dA$M��؛�H'߾�?�P����%�����ND�,K��Z�	���m�k2&�X�%�y���Ӑ� �5Q,O�sҦ�X�%�����ND�,K����7ı,K��:��M���UtU]�/�RB�����q,K���ͧ"X�%�}��Mı,K���ͧ"X�%�I�s,���R�ֲ�k��bX�'?}�m9ı,K߻�q,Kļ��siȖ%����띕7ı,O��~���	����w���oq�����D�Kı/���r%�bX����Sq,K���{ͧ"X�%����>1���
�E�tF��cigU;&u q:��S�9�tD=�@j�EЛ3Y��2&�X�%�}��ӑ,K����ʛ�bX�'��m9ı,K�uܩ��%�b}�ۆ�K�2�n֥��fӑ,K���u�&�8�~WB��"X�����r%�bX��w2&�X�%�}��ӑ,K��E��.Ja�M՚�J��bX�'﻾ͧ"X�%�}�ț�bX�%��{�ND�,K�w["n%�bX��t�a4K��kF[�6��bX�%��̉��%�b_�w���Kı?w��q,K���wٴ�Kı�޿`P�S&4���7���{��?�w���Kı�{��7ı,O�w}�ND�,K��s"n%�b#�>���mǀ��Y1�d��b�鳖�gI����+�F7�Ľ)\�Mtk�aK��e5�ֳ3iȖ%�b~�u�&�X�%����iȖ%�b_��dMı,K���ͧ"X�%�{'�̲�j�K�Z�u�"n%�bX����6��bX�%���D�Kı/���r%�bX���l��
�bX�%����\�j���k-�5s&ӑ,KĿ}�ț�bX�%��{�ND���F*�"D@!*�������wz�q,K���o�iȖ%�b��*��]�恭������o���m9ı,O��D�Kı?}��m9ı,K��̉��%�b}���Y�	p�ղkY�ND�,K�{��7ı,O�w}�ND�,K��s"n%�bX����m9ı,�}�wo����U���v�م
�i�F�+Q��2��ټ��SGYQ�j���������e�L3	�Z�s��bX�'���6��bX�%���D�Kı/���r%�bX���l���%�b_��ܒa4K��kF[�6��bX�%���D�Kı/���r%�bX���l���%�b~����r%�bX��>/r�j�&f�Rf��q,KĿ��siȖ%�b~�u�&�XbX����6��bX�%���D�Kı/���Iu�pֲ��ֳ3iȖ%�b~�u�&�X�%����iȖ%�b_��dMı,qQT�A�Dy�?o��m9ı,�N��%��.��aq,K���{�iȖ%�b_��dMı,K���ͧ"X�%����ț�bX�'����տ�hq$�ZTGO"ef��Z
�]6k��qmuÇ�S���ܹ>|pˉ�ݣZ�O�,KĽ�"n%�bX����m9ı,O��@�(3�5ı>��iȖ%�b_���k^�ˆY�jk2�fD�Kı/���r%�bX���l���%�b~����Kı/�w2&�X�%���oT�5�&an��kY�ND�,K�{��7ı,O�w�6��bX�'������bX�%��{�ND�,K��l�)�a�5��0���%��؟��xm9ı,O��sQ7ı,K���6��bX�'��["n%�bX_��ܒf1�2$�|.���٠z۹�{[ŀ|�\G��	�U�N���� $   $��3 �Y}Z�ݻ>z�n�Z��퍵B�\�iB�>��v�񗶶3<�]�t�1�8���7R:�oe�뭓uXS��a�hӭm�� N��c!&k9플Z�:�ۯ.{f�ykO���h��^�-�*������v3w:ͮ���8n)�=vBx{X�ɋ�c �mO����&8��뱷-��h��B�M�&�v�.�Y7m.-m�Ɖ�b=-���hʛl����ւ�h���Px�I��8ț����M�����/�Q��:�����Lښ�]Ҫ��ͼY�B��_v,�� ��f����o��D�����.���L`l�� �e�.�6�s	�8h�נ�@��sTD$�~��� {vj��Mͫ����-^[ ���:`v�t���[�������-Ɏ�s�m�SC&i�oc����m�k�خ%���im���\���r�Yw��;�t����ˤ���iIând�v�USsv���Y��DBIC�� �>�ͼY*"X�}��&����!�r�^�z�4[w4�)�}���8�iL%�ՕWX���}׀owb����5u�@>�I\�iLn,�I&��n�T$�[�/���� ��uSr�p�kmɮ�C�N��FFbm	>k�˷k
�G�nQ�Nɲ���q�5��0'tt���[ ��$t�<uu����m�&F�h�׿����wu��ذ�`����7d�MYsWX��6�a)D(�
/!����Q.���f䝽�u���q�E0S̊I�z۹�wu��9u�@>���\�"$L�Wke0;�:`r�-�zI��:`}�Įb`���&�dɃȰL�fXڢ-qŵI��d�aݳ5c��7�MY4n��~a����
c�dI��_���٠[Қw]���]m)��87�}d���`wtt��t���)R�6���Ȥrh��h�w4]k���@�P�`7�LX�r&�4D%;��X��`ͻ���!(���zS@>����ۈS#s4
�W�[f�oJh�w4�^��$�b�[�I��77�p�ҵ&Nvugl����3���1���vN��썺��ߟ��vA����)�����E͢mB�����g�+IU�ŀ~_�W�[f��/�b�$���fS���.������#����1L
c�ys4]k��f��n��{�٠}�n�ěJa#�D�-�M�vA�;��S��'��׽�w����������  -�m� 4W��K��X�Ñ��sJN4n����-t�m�]�,v+`;�=v+��e�5����٣1��M���{=q�h�6����=��|����6%�z�){R�g(k6���Y��z�k"(��z�/l-����'ka[�͚�y1>ؕ=�gn�ql�9�y��]n`!�� ��q����-�ln���n*s�D2Tz:iWv��0��+��n�<����su�Ώ6���p�5a�<���iLn,��'���O�^빠Uz� ��h+�'`7�LX�pI�@���)���1�'d�R˼�.�j�ɛWuk r�� ?7x~�P�&{��s}� 5�t\ݓ4T�X�^[ �&0$�wGL�K`wv��&
!���-�M�f~o�_�ϫ �� O�2���
"%܇j��v�u�K���7-�벦�/4�:�sܵ	<A���4�D�0l�$��]�.���1��GLkeL��]
c�ys4]k߿�p�l+�hz�h��hg[�q&ҘH�Q'�{�cd����tt���[-�W &Ҙ�Y#�94[w4���˭z�u���N�o��D��`n�X%�u|���6�a��w���{�ߪ�qU���m��j�쮪�I�y5�B�b�I�|�L�3ѪQe"i�S#s>�������=m�5��s@=���)���8���$t��tt���[������`�#�h��hw]�>�����4d �E ł��F)$�`0!�@�,$H$cĈ�D5I�LAo� T���8 E7 D$H*�-!i�����D�,Ql�HZ$��Ab��B���)JA�!P�D"�"� B"��]�$J�J� ��n�0�P(/�M�Z��X�����;��5��kh
' �`�`�`�{��f�A B����I��M[��3	�C30؃� � ؊`�����<����u�{[T�lllo��ٱ�A����{�6 �6667�z{��.��5�b�ֳf�A����ｭ�<��667�{�؃� �(�`�`����y��mD�A�R��o��V�k.�$�0�%�wV�q\����ZS�o�v���YN��XE8��
he�������w߿����i8*����~�}�s �����ℒJz������UW*�����݋� ?ʢkS�{�f�B�_krI����B_Hzt鮰�U7!75e�V�>IO���t���7׀y�� <����dCd�L�L�9u�$���N}�{�$��E�X� � 
��g�'����ɗ2�iR����oL`z�GLt�05o�w���?�V����CX��۔��Sۦ�9z�M

`��smUȬWB��R��(�̒I�}�w4��h�נ�1�Pı,Feb��ox�|a�	L�}Հ�_BI}!�݋�Q3��h�R&իUAe]���Y�	L��׀|�$���_���rI%(�_ߵ�$�S�M'����f.�����X��δ� s�m:
���(�b�ɠz۹�}�S@��+������I���w{�?�� .�   0kg]ͤ�ݶ\ڸ���9.	����㖺{��h̘θ*֓���,�N�FF�룯^�6ۡ+�&�?ϻs�o��
 ��W&
]Y��w�$,)u����m�쳬�f��n�N�x�Ñ�Y�x�\l�96��tl�N,�W��!<�����K#�v��i{S�pS��p�mK�:4�ur���v4�w\��*ϋ��2�{quC������2�r��8��Ë<�����d�Ú��B��_��r�����=m���ZM�Ȇ�m$�Yr����#��d�.����I��Lcn= �u�����e4]u�wC��"LCd�F�0=� ����`�1�H�J"L#��}�S@��^�{����� �Ա6���R�T�Wr�J���U[`��}���*<��u.�U��9�!0�<�����ߟ����]�m��$�_Hy��y7�D��T͢殪����ۮ�ҮP�����P����Phd�����?~�znC�\�$~W���Ɖ�<��rh��0=� ��ҥ�����+�&,Q8A���e4]r� �u����׫I���"�����J��=�1��GLt�0;k����W�[#f�Wh�2����R���ՅQ��"�W�H�N��"��漕�[ ���:`{z:`r�R�����F�
!�I&��n����h��z�����B�(��&
�.������6u�XZ�J�Q�s@��s@=�I���"<�9����u��loL`l��oGLV�u�$ƦH�&G��f��?����g�~��s@��+�>�뭷1�Cy�JCbwi���gY�r-��
C����<�kU�;N�"��y19$�=m��/��h��z}�h+�'`,l�ŉf+��ގ��UU$r�N�ޘ���s@=�kI���$iH�h�T�7�06H�7���˪�(�l�'�O#��@��s@���|( J�	�����Y�2njK�n��WWk �o1��9u���w4�:T����b`b�T^li�F�+1����>��vÆ���v�������"(��&	����/u��9u���w4zS@>�\�L'1���s4
�ez����)�^빠{-��cS	"���}n���0����_�� r�u�9�����b�$�s4zS@���W���]��y$���X�PI��;��S�[l��vA�$� ��  j�E����ΐ��3�=i%.�vX�c�����~Q�1�P%�m��`��͡�m��Ol��Ԑ���$�^�E��N��$�	f�.�Х��Q�.C���g'k�y����eջ\ў��`��luc�6�Ҋ��pK=�̦Y=Y�4�SZ+���{�mC�v76�@�=���'D�VS���)X6������҄��<�׉a]�Fc-2�E�N�Y"��<����X]u���m�������`�򈤡%�7ذ�����쪪]��WXͼY�D%2w;� m�,��� ���fꤺ�����ޔ�/u��*�����hv:�D�)0LR)�]�S�[l��z���Iy�1��s"Nf�U�@��s@om��x��V̺�A3Q%��*���h�f#�瞹���쯏.mq�sq��s=�EcS	j%2=���ޔ�/u��*���{9�lh��� ݬ��c��	CWe��XO5Հ?u�߿��1!+�7`<l���N��X������}� �w� |���ڍD6I䙠U{+�/��h��DB���, �D򮹹�uJʼ�J�-�7����`M���@�e���6�� 19�c���p�aJ��펶�K�o%��8h��3f��Z�0JhĦ��f�oJh�w4
�ez�]��eE"Q)�L�C@�׋:!)�����;_b��f {ɲa0`�Ɔȓ��U{+��ADD@��0��`ZǔM�4L�.dp�#��f�oJh��h^��
��Ui���8G�@��s@�빠r���Y�wc�6؀�gG���!g���#1s@��m=�v�	h��7aL���HD�n@x�d#�s4�]09t�ll���#���K�v�Q�FI&h��z}l�=m��/u���e��b�f91'���1��GL	�09t�l�Db�������]���;�ɀ�"�`��A#�$1 E��D��V��� �H�"1�!�Dy���|�G�%���19��L]*[oGL�:`{je�/.�.� ���vͷ�2�TE����r:6Nvړz�k��n˷|ѭ�W\ػ;�.����r�u`��`m�����C��,ɾ�&�RZ.n�f�� ��r���M��Xk�Xδ� s�.�f���7VZ�j���,�^,9D%2���~��s@�^I��d�d$�s4�x��i� ��(�;��, ��_��Q���#$�4]r������,�^,קw�!BT����$`!�|m�l#$�#ŉ2�+j�!Z��#թ3N�Z��0@� @=`1!*�b��l�D꿂R�#�XE�E"R,VyCCK���B��@#@��E`�$ ��G�,a�H�c!	��K.��M H@7J�ЉбK�1! �ʃ(�T �b@H4��L.�)bj�$B*�a	H4Cl4��/N�	 "E�X$FI$P4"�X r�H��[��    �         $�m�  m�             k�m����F��gCU@%�)�
.F*�)���Uu#�V�]�͍�f��Y����;m/ʂt���i�;m1&B�-��G6��*$�fw)P潶�������o�>ۙ-�T:"]�mI8�Vܮ�l��j�
(	��盀�:� lɦ�3������B����v�;�TΆ�W(J�p յH�GN��g9Q���H��ȼkf�H�b�g�LN�+���#S��+(�_����.��Jeez�Vb��3�7!a��Vu�r���Y̯U�cC�v�����v�U��jGKz�c����RY� -4���-��������K"N$[l;	#p�D�i�Yx�A�1a�Ѧ�[U�8�9ճvV�ʈ� �f͞�k�z֔��-��\��F�6���qy�N�.3�9!ܴ;M�BL\�/M�� ��ޓ��t�^mz�vC�Mt�R��ҥ�Xl�����vUx�b��j+j]�wQ``���ڞ	�]���"e��`
-��`�ͻ[e5̃��F��3��.s��ܵ�8kj�2��
*�ׇ33+��f�o(�<�T��ں���7@ʡ�$���Ԩ�H .���LbB@��m�I�%1��r�^��8{c��ق5�%$�s/:m�g�m�|%ɍ�����]���ꫩ�1Nh�z\��$��玬��U���T��<���*�R�UPr���崪y@�$0h�3c�i&��\ <QK�J�Wl�Q��n\]7sR���m�nk�-u.d�D
�T��J9r̪���Ʈ�L�öm��k�i$qmT����n�R\ ղ \���\�k�g;�Cm�ٜgNx�1�q��d�.�R�0��۠K���-���ݵmѰ����W.���J�T���[� 
�g���
�ʾ|R��+m⪡�P#�?�(��D�??" ^o��������   i��k�\��9���(<��]�V��z����Dt������r��yd�/���o�����;Y��L���t�p7�����N�6�l�'+����b�-J�YyRK/h+v0\޺�қc����m�bs�!^ޭ�[>�jv�V�U�v4Æ�6�6�nsI��4�E��u6������s�-s�N'ð�^)V��8���,���N��ٱv"�q-88����O��n.�������$Uv�i]p�ذ6�`�w4]r�����91)�p���#�ގ��T�ގ��*)�LNb$s4.�^�}�s@��s@>�VT��Cd�09t�l	�06H�7����V�X�0�F�S#�/��h��h�w4]r��X�cQ�q��\��z�����T���hc��lՔXӍ��h��	��=m��.�t��ҥ�&�t��԰ʻ2�d�ɭa�'}ݛ�;"���B$���/�V ����x�o�M��Cd��I��f��t��޷s@���hrel�"1�%u��wd�:`{�:`*L`wvJɎ0�Q�s#��;���>ʓdt�+w��������8���n��LY�g7S�ExW,[ڠ8��/H�xL�I�18	����/u�`*L`M���GLv�Č��S$�'3@=r٠_[��w[��^빿�#��O�qD�<�E#��I�v�b�7[Ň�D$�BQggf, �]�@��U������������wGLeI�:��� �ԗT�ʻ3�r&�h� >��z���������x5'�QF!�����n�h��wk��-��t����v�m<�J�l�27 ��f�z���������eL$�c�'�M��:`N����od����i7��u���)��l�/[��}^��4�'19��`*L`N���_�)0ܮ�L)��9 ��f�z���������sJ��a��bxJ��m=YQ�����^"n?�-�v�~s��k)۟6����#KɄR<o$������w[��^���������M4DG�e�S�GL	� �6T���#����,������/YM �Rct���:`���e�E٘�����l�1��#�t��$��w$�
� F#�<rh��`���<ݳ <�w�		/�BDX1 Iħ�g����ff -�  u�{ed^�e��H$�X��Nˌ�ݱ�tIDhv��9"6�Na0�m
ӐvMOd�LE���#�dd��K$���p�ע���y��5�̖�bX�1�!i:9zݍrp�c��Iu�̵�s��k�܅=����0#��R����zy^+5�t�tŭ���vݓ� m��c�3ɝ箹/P3v^t�)��{���qA*�L9�խ�mX�;nRJ�On���z�M
+�-���k\+j�Nut�{Nr�-ߛo�߱`nـi�����b�=Ԝ���Jbp#��z�M ��f��n��n�{ȴd��H���l�1��#�t��&A����[�%���)7�M��������h�[4]�VF�i�!H�.��:`l����t��o��~*�]�v�\���B�9
j�YR�&a��Ë<�]�Eƅ��=[<��d$�s4[)��l�;���;����9T��Q�)�n���J��o�o����72�?4L��r$�ɠ[����n��e4�-��Tl��#�1��w����d�0�&0�I�ަ�tK�iLn!19����?fN��}� �o j��U]*��6���Y��dyD��Sm�<\q������l��6:��eD�u��][.����߽��`wH��#�ɐ`{����Tҵs7v��������	B����X~�?���Ucm&�	�E#v���`ֹ��J�7xz�`/�6@Y�'��h{-��w4^���9T�&&̵���L����06vA�%�>m������8�\κ)�T���Y�Nɜݞ�`hat�̀��۫ۤs!;I��3�I�@����Қ����[4��لDx)�ns4[�_D�;jL`I����I�1���"��-}V�w�٠[�s@��M ��U2`�S$��C������xs�X��0:!%�Ewc��v�8��Tҵs7v�����ŀy� n�� o�w�t$���m˔;l��/=6���vV�l�o<U�M��b�k��<[R����L�`I} �1�'GL-��6LBLI�@��Z��f�o]�ץ4��U&Fɉ�5?�q0ړtt�����0	W
�2db1ȓ�&�o]�ץ4_U��h{�'���S�����0$���vԘ�����?��� .�  T㭮�@O[[c���$ɵe�`-d�M*G-סЛ�?��_O��ixɛ<���������2��ڭj�J��c2��d�8hxu�ٯN�7L��Ic�%'����x���盳��Řx��Ӽ]��4��RT�<b"<�v�ӱ"Y;m���@��܍d�=���X��m�r�nzD+�J.4�6G�����~u|�4��X��XӰ�RVc��m]g��73C��z�j����Z.XË`���&�RcN��; �=�Z2`�S��9"��[4z:`l�K��J��WfV%�cy$�-빠z���k������+#i�B�H��ץ4_U��h���>^uD<l�*�2��_D�;jL`I��gJh���r�i|�,J#���ߖ� ���,ZV^�Ξgk���"�Ç�
�Fɉ�5?�q|{?~��w4^��-}V�uEaZ&L����I�7�|�ItU�|`��p|������1D6
b����Қ����u��w4W�T�4�7�Y�0`I} ������Jh�e�&1�#�- �gX�����d_D����g
g%�n�mO[1���x�����9+�6o1N6�5���,h*^����׋ �� n��DD/��}8 ֊�����LJD�s4�Jh��@�c��Jh^uD<l�,�����>u�p�s��$�	T""B��FA�8tF	~ �	>~�q~�D�� ���F ECq�d,`E#	ň��(Ƞ�"D���`�Pb�U����Q���T:&�H� ^��b��(JJ+%�}���>{l�6K�dl��Q����@�c��Jh^��>���-aZ$��'�E�o�ـ|�ـ|�\��Z� �Q��}��VW5�A�>��f�ِs1�u(�+�Of�9�
�b��j+g�m%u�yWy��ߦ|0=/�`v��L	::�=_
��4�7�)��k�ھ��'GLN�06��YEв���9"�;��Z�w4�w4_U�}��Zɂ��"RF�H�z�0;�t���&[+#L�EҲ�bl&%"r9�u�����=qڴz�jI+r[l�A�5<I��N�]����g�k����Z8��p�m���ղ�!�d�d$�s>�$�r�RIz�{�%$lI.�=^�I�Rՙve]��Y�+�4�[+$^�II�K�Og�$��QjI%㹅h�23R4�^/y$���I%�'��I)/ �I-�-_|�^|��1�6
b��I%�'��I)/ �I-��/y$���I%��U�I�1���%$���%k�Z�W�L�o9m��w�7m�����qB$"t H�b�
���w0p 	   	�ۚ�"K�٘��M�#n�۶ܤ��k�l���9�v���v}z�/^6u��[�ه�s�C�q���]�U�������'��[�.�]���Pܨ�<�R�R�<Bݻu�$1,�OY�m-�jet�v��K���O�Wl��v�e�:ɛ�l�k<���ɋ�0��Ô(��:��v>@mf�l���X�������C�l����`:��v��Xn�k�� �u�';�I�����%�;�X�&�h�WgM��I)�����$���i$���{�%%����;��Ҙ,n"%$o��J��4�]�z�䒒�	���Y"��H�1K����!)��Ԓ]���|�V^A4�[+$^�II�Kס�!�d�I!ϾI+\�Ԓ^�-_|�V��Ԓ]���|�B�*�"yۍJ@��Il��{�%$lI.�=^�IZ����/Vے`�"�l��g7:j0�е�:+uWKu���}�����x��&FcJF�G�$��t5$�u�g�$��QjI/\���I/>R��	�%U�U�L���/������wV��Iv�H�䒒6$��4�b�)dCx��L�䒵�-I%����%m�I%�o���$xykY0x)�`��IO�}�&�JH�4�[�鴒��Ԓ_gu�����"R%�E��%dlI.�=^�IIy�Il��{�$~���*�ҜF���6y�+3W,#�z�p���ql�<��犱�u�Ҝ.�(G$��$���>�$�r�RIz�}�I[wCRI|�ح�x�0_�HG3�JK�&�Ked��I)#`�IwI���$/r�2'��H��
AjI/\��r�{��rn݈�;�o7�w�9�m�l�5$��%�*�2df4�I�$�tlI.�=^�I-���Il��{�%_GrL��L�7RIw[�}�I-���Il��{�%��IV�%.l�����k���Ea�Dƣ����N��z�W�����\��,e��I%�<I-��/y$��`�IwI�}�IZ2`�S�?�8�I%�E�$�tlI.�=^�I-���Iz���mL7�,�/�I.��K�OW��Kdx4�[+$^�IPY+.�&Ȅ�����n�߽�|�K�~�jI-��/y$�����`�Iz�:��]6L�����^�a�$�rZ��$���jI.�~ϾI*��m�&8��2I��.�uթ�euV�M��S-p&�+":♬�d�Tv��Jt2�� ?z��??�tlI.�=^�I-���I-�ҭ�&F1$��K������^�a�$�rZ��$��.I���Fp��$���>�$���jI/\���I.��K�ڕ"M)��7�)3+�I%�<I-��/y$��`�Iw[�}�IZ2`�S�<�5$��d��I.��4�]�z��[#�����׽���~~~~� ����� �^Z�Y0�N����8��g�v.�"�\;��.�]Sm�'Tܽ;�Ia�'\��';N�!f�ms��؍m�dX���t==#ucC��[���\<�XUn��s�$� uل3 #���t �\�ֈ;u�su���}�*s��7Lj�K�"�^��W=�SӸ�Q�s� ɻl�3���q�θ�&�X_c�	�n��q�tPUGV�\°�3WX�M��}�';��W���sֺ�U;�.�,�bU��ܒR|�4�]�z��[#�RIz�}�I��Ʊ<�J� 4�]�z��[#����Y"��K�=I%��b�D<l�/�$#���$�k����Y"��K�6$�t��y$�:���c�5��jI/\���I.��4�]�z��[#���[�u�.ɓ#�h�"���$���>�$���i$�Vt^�I*�~U�|���X�_/=`�4o7h�V{t���B�8sķ�٘m[t�-��4�e�[o�w�z��[#����Y�{�%��KԜ̰M)����I&}�I/[������~��b]+'���]Ѱi$�d�{�$xyhɃ�Ls�#�Ԓ^�:��I.��4�]�z��[#����oOX��<n"%"Y_|�]�t5$�z߳�I%�<K�j�]�����I"��>e媺3%�3Y��n�o߻���*k�{�9RJ�ٿ��I.��J�-����6�l�qL�&������r4�������.�R��w��������FD�g�D��� �}�������$�tlI-�z����L#	�H�R7!�$��m>���J����������L����3�!Cm%�*���2dc#�5�|�V��&���{Ü��� �e���M�m��M�~~ �����iظ�l�� �����{���fv������ֱ�}3?�P�U6��&���'��A)����I&}�Im��i$����I�{�u$�>u�$�H��?����+<�]q�n��r�r��Mf��g�\��&����:�b�GY�ut�e�w�Ӯ��:�H�Uh�����w~W��>�x�6�`.����CS����ۯD/������X�w��7Z�`g��Z��dȈLrL�=m��>]���L����<�b�>���.J��¢��n�`t$�g����_ۯDB�1��� r۪���Uwu77uWx��f�B�7�/��݋ >�@�gV���ljdȒ�72c�L��d�n�J�4�����,l����HK&L�dq��C@���h�w4��|�I}!���ϕ���]7U����=���Q	)��}x|���۹�}��$4�7O!� ����V�:Dϛ�X>�X�KZ��H�Uh�Auw��w�g��X�x�?BJg���[ݔMM�����n殳���t����06J�0>�w*Q6B;E����a@K����v�BE$��u��ʇR
��� QC�����H$�u���T5Qt	 �P�	iN!EЌD�(E"7�C0A ����Wu�Ď��"|� `�8a�� ��i!�'�����@    �         q��  l             
���%�-����j�܋Kv.���Z]���\��v^�����
�M�W�u��7��рI�;t��v�bd�Q���i��ی�Jnɳ$�m��jq��*�\8h�V7i	��f��sm�]x�G$�L�P�t���1�ۉP�u�h�*h'�E��ݽ��@p��ؘw�����+�%�q���ۇm�k�j�vo9UL��s��)2mm��zv_IF�vY�ivG�sٶj�ۢd�!sf�Kci6�]d)�7A�a���&䵝]��-a8��wgt;;�i��V�Y���n��橶��ͧv�[WV���6U�˰ԯ3k�,k�	�vL���*b*vQ+m�i�rhym��e����t�,l�Mȹ���5#�+n�!Xrs9=�В�]uI�ki�:9k�������N�>�\�s ��&tu�Rtϙ9ު8�1r��X#bȷ,�]	�n�𘦎��!+�V��]�:�=`��9���% �]\ۆ�gb������\�O/^81��.�8�,�jj�6� m��t��keڠ"c2�
U�N�̫���fLs���ؠe�%j�jdx�5[� �]�Ȭ���f���d�G
��i�
S�;v�5b� �H�0ր���+e�WT��"٨�M��Ҽ�j�iJ��تn6.ge�J�nι{.��%t���]V�I���d�����`T�5�P *�UI�q�i�;���w;��U��n�z@z+��hપ��T[u��^]�G;��^��%ڮ=7ik�1˚Ѐ�X�UU�Y��yz�����@eYX��L
@�nN�jHm٭�-�[F���S��X��Çn�j�McCm���˹��8�;��w�j�'K�7]s�r�C�r��ī:���yPn���mK$��,vveں�퉕T�誩Z��&h���b�)�T��)��?�@�C���z����30 �P  M.����q�<���l�����X�ӷpbȜm�Vm�q���
6K��+.�Q����P�P�m��rK=-�h��k�sĢWij_1�M������s2t,���0�	KQ�Ns��mͱ9#Vz9��R���<��Ö6�2Y9�Þ�G4e�m�8:�X��͇�.k��=L�Ogd���e[* c���cN�xK�8�&1��sb��8���6��ޛ��HYb����UjU�.��^�� |���ճ�#���`�Ծ.F� ?�#��}z�h�%4����n���H��e��L#	��آs4�W���ŀn�� �u��7T�Q�@�q����빠{���>�䦀z���0�#܉fSzGLwGL�Y�������~}����0��`�a��5���A�knz�c����oj#�P�a�B��j�f^W��>t�ޕ�`{�:`oI��_:�&1���L�=�%6�iC�|��K��ٹ'߻ݛ�s�,�	DD��ݝ%M��*����R�0��L�0=�07�d��L���UjU�-UݬP�u�|�7ذu�M�빠|���Q4d��/2�ҲwGL�0?���~��kXvx{8˨�jim$,�RvcZ�w@\���8{a`�Tv���B�yL�Y������'�� ���m�c�%2C@���07�t��tt�ޕ�`:a��veЦ��f�`��`n�X\DR���f�W��}� �җNh��mU\��]լI(�7�,�W���ŀz۹�_:�&1���L�;�d$t����J^�9�VS�m�u���a����]��9�;�����S���f�]�y�JW�|��#��0;�A��+ ����1Ʊ��&Bc�f��n��e4u�M������i�&?����dҲ�:`oH�+�J�Ǔj!�{�Jh��h��`J�JTD7�q��_+����#pS$4[w4[w4�)�n�l�:"�.}UUuUt�j�\�.�*)*$0�\�ml��2�ח��M*[��C,��Bd���f&��������e4뒚����y[��iLn&ْ���v��Jdo��k�ŀy���_:\��`�9�x���䦁��遲GLoGLV�t�eWW���.�����0=�0;�Jhg��Z��sL��$���X�׋ �jـ}�x�
I5
����~  �h  �������U��T;v.�m���5�u��˳��ՎE9C:���v ��t�s��]5ym̻[%�u�G^�K.�9��Nݻ8]�/KnG[:�j�؛�ݶ��Ge��Qt�q��:;m��:��Q�m�{l:��*cFLp�eF�J��ݬ齻1�,�m��P��e�"N���M��l�sv��y?��t��䫺Mm�뭇��:�]X!���[WY���kq�;q��&g����ț�}+/2���0;�dގ�$t�rj��Z��VU]]��[3�"Q�>t���� �����J˻�31�2C@��w4[w4�f${��w\��w7����$���}�ۚ��4뒚�빠}�+u�)���2I��@�)�}����=ZU�ldPn`��!��� ��2�E��\8�g��w���k2�m.���6��D��|�W�����=����g�<��z���bǊdjF�Hhގ�$t��ޖ�`z��Z�o��d&I&h��h/uzu�M�u��>^U��ƚ2c�&))��-��+ ���t��#�D�bI�Ǔ����rS@��w4[w4�����[n<R%Q����pt�-Z�
7%�]r,��.����$�F�d��L��>�]��n���W�{�Jh�XHF��3*�䛵�{[Ŝ�!L��}X|���kŝ
�<�uWUTͪ�������zu�`�[0�I)��DBJ=	*ʭ{�z���t�Ʉ�Lp�$�@�jـ}�x�6�`r���������1��25"o$4{���s@�zנ{�Jhgu���!�(ݕŭ��m
���*��ه�ql�mA�y�Xa�q��'0ɐ�$��{���<�K`oJ�07z:`y]s.�h���h���}>n����_+� �}� ���9%2t����	�Z�������՟ގ��:`yl��7���Q6H�8����s@�[��9~�u�+�"� U}�����$#Da����4u��˭z�䦁�빠�䫏�A�ƨxj�a�Ŏ��N��G5��+¹b��SvT�#")��e�B�wSwͷ����~�+ ���遽#����fQ�Lpf)#�=�%4w]�������9(P�&C�e��R�6���j�ـk}� �o�BS>��X�+�@�{-Z�k�d�LrL�;���>�n�6��
u��`����i�&<�Ƥ��ֽ�䦁�� �o �$�$��������������  ��u��4
��8�n<�cn��y�5�u٠���� {&礕�m�nvx�Iw޺pvۙq�5n� kts(7ny9�5�X�l,y��nb{M���k���nKi�N^�XK(��a��CD��q��պ�WT����v�	ۮM/f�N�]����j��mlo'C�����x�;�4�H�W������Z�۝�cp&��[���Zi7*k�%l롸�y♬�d����qj��&j���+� ��ŀn�� >�f�{/5rD� F8�S$4w\Y�27݋ <�� �jـ=���h�#1�Rf��n�}���䦁�빠}^T�BS��B9��L`l��`t���GL	��1�)�l��h�%4��h��hu��s�ҬA�4�!�$sZ�%Q�����s���|�|<�󳣕9�ɘ+J�x�����7�����;�ŀ}����J#��W��W&YJjЭYj��`���؄�bIjK0�{��}{%4w]���Ӯ64ѓ`��e0=�06J�0=�0;�y�Uy��(
a1��5&h�%4�^,u�X�>o�X�꫔��1��!�}�w4�w4����rS@�gV��Fbx���51G�$�i�4�<�s=q,�/<i�;�f�¶��W}��v�a Fcn$�π�����빠zܔ�>��O+�iLn&���>�x��
d��|`o�`���/���L �8	�"�4[���}ݛ�/t�AD�
�B'	9�֨���c(@�(�	ee�
��b��	$Eڇ�E�!$Fi�j-�H1aU4�HX!��e-�� D��	 ��H �Z�D���H���U9H)J��@��!�dX,����@D���0b�"�j��W�k�SB�"FB0���"D�RP� "B�H�b;m"8�B�h�����+ H@�4`A$R$X1��I�eD`��Ԋ~UG�ä	D] > ����� SoW�: �U�N*�&�7��o��ߺ�h�兠�<x�F�M䆁��遽#�������յ	&YJjЭYj��`��`
<�|��쟍�빠w��m�<���<���IfLs�̨P��i���k���]�ϭ*���r8�cM1��I���s@�\�`{�:`oH�뫺�eV�~V�)��+ ��tt�ޑ���� ����6��1�	�Š}�w4�0=�0:U�Lb����*��fn��^,u�0j������R���@6���������<��1��b$�4�l�5��8�x�z�`
Q�~��a[���w\�H3u��"`��I�ջ�l�n۝�˘�{�"��]u��.l
M�ݞ�*�Ӏy�� ׯ����Ǐ�ԍdqh��h::`{�:`t����D<.����U�e0:tt��tt��J�0=�w4�u�Pi�&<dprf��u��=ҲwGLt�YukZ-Tܩ��X�ճ �����|�[�XۯС$���]�ڻ�����-�m� l��f�$�5R��l��:�ݺz���X��O@`=�ay�k��ht;&g���&�����a8*pf�����p��@���㪞��ʼԉE�v������n�	vi�=�����Ļt-�,g�;� u�����T��V�c	u�V:Z6�Ǹ���]�W�v�'n�n��}�pZ��SD�˕
��s��Ǐ�|q�ԍ�p�l%� 2ef�Ýp��(�N���[���RF��F8�$<^���{��hw]��)���$�mĔ��{u��>�x���f��ŝ�
����Q��Q6�njiIwv���� �]d�0&���0YW�UD�Uk�|�g��X�^, ݶh�g���1��25&5����Dk}�����>֭��)������&}w;�%�k�� Ӎ[/6��'�Z��V��z��5�ݳ�9�}$��?�� �Ҳ�:`�L-aSR+T����� n�y���%���S��=�ذz�`^���Մ�2�b��f0:U�L�:g�O�Θ��M �Ȩ��F8�#�@���^, �n�9N�Y� =�ȻH�ۉ)3@�[�����rS@�[��}s�II�F����6�M�<��-Y�͵��ѹ��a���ś��P�Ƣi�$�4.��뒚�x��}ذҙʋE�j���.���Ҳ�07�t���[ ��q�x�L�H���n��sO���@�\��=��F��q�K�X:��X���ճ ��� -���hɏ��yu�@��l�=���=���?%��u3�(�xwWg���Ō6��33hqOGI�n,���.\����A���b�rG!O��V|07�t�ޑ�WIlNDFV��1�1)�����$u��s@�~z�䦀q�Ff6�sUk ��� ��u�B�����5�b�>�J�-Ƣi��I3@��^��gf䟾�vnO�_ȰC����KK�=�,�l���Y6��j�����ճ ������}ذN�X�������g[�t�֖4,3�ۇ]X�͑Ð��3u�����9��=7<�t�5J��=���=���kw�#�J=@��� �q�rniU\��.����o y�x��f��,؎I*��I1��X��y ;���@�c��wnh������L�a1�qɠy�l�7[ŀn���%;�׀�#?6F�9�L��;���;���[f��rS@�[�I�I$�I$Zl   �2ɶ�]��ָ�\��s�y�`��x���N�|z�Qy-p��v虵��֖Gk��>�t�ˮ@��5k���u:�e��]��N��4\�X��[I�N�c����Xj7..<��c���V.�w$kӪ�O�bc`t.ݙ�6{v1[u�IdA����d��5�5J��H[m�N�-�ٌ�n]m�h�t��5�k5�f�.�	�)2�ЈL�*�ckg�:�)f���[��C0[�w�6nF��3q
L�?~��4�٠zܔ�;���>��^Ƣi࣒f�z�4[��u��u����;�ڮTZ(�Ws4���� ��|`����S-�b��������6�Bm]M��+��Q�!Ww��Xw����e4[��gqQ�x�0����`wH遲d%d�:�������*�l��҃Kw=\�:9s+�n�ݔs��Y-̇n6��٥��������R��W7k�7���<ڶ`���;���*�N�$�Lx�q8h�[3�S#}ذ��`nـ�2�F�H%2C@�s@�s@�����M ��L#�m�+���DB��%]���`���`�[0�w4��׀�1��x)���c0Д~���r���;�~ŀk�f������Ƈ5���yB�/e��QOQ���#�ܻ;@鳮�.'_�ĝ"�;GD�E܌����Y�����Ӳl�����q����7��u����S#�|`��X�V���re���E�.�f��{l�>�x��J
��P�M�S��v�!b$�0@�0ZT`�SH�@�����_� ?ou�i�S6T�ܢ�b�.�`{dt��Ր`�1�Ӳ]�㤌#	�I�3@���h���S}������=��`Jzꪪ��Sp*���m����s�ҭaӹ�\��z�C�ttX�ksh�4�G2� ݓ{ ����ꪯ ���ɀi߿dm0�#܍94��>����>�@=�@���W��1��y7wV`y�X�s�D%2n����Ɓo/����H�ƔNf�}���{]��l��(K�J�.���ߦ�\3����b@�F�k#�@=�@��M ����U���6�"s�v�i{�3`x�#5S����xsY�#\pn�S��oQ/N��&���������`�n��Z�"����r���ME����h޶h��� ��� ���興�:u�)]w!t��!^f0>��`�1�7���hV��1�dqh�/u�4�|`��x�BSڭ����OK	1�܍94��>�]��ݻ�N~���&qF# ��
	(0H�!*`b�8`R���u�a�b�c�"0$�*�D4"(,U���Y׺{�t�'��/���~     -�        �m�  �             k;�Ή��s��@�'j�ƺL��]�$ m����`�V�j�ݻ�G*P�{b� ��:D[z���3۶q����UBjcv�lH*	��r['i�G��JK�G6ח��ژ�z�,�*e&e��iP��s�ۓj��v��>xw(��AWm+*�x��ݶ����k��h�+e��s(2��m���%���� �:���ٞ ��Qb}�[j�.e��C�P��#��VK<�ͱ�����/73��7k%��%qu��9Ҷ뺶�Ȁ��t�*�<���7m�櫫��QZB�ܫ�fa���`%^��4�\檶��
v(�y�&v6k��drh�XZŬ���� �4[.n�+m��d-�6iQ���K{j���ha���j��p V�nng�Zp0,��C�\�\�k����<�'���JT�/:�e=��V��gF��E�*�*@eT�[wMu: v:q�*Wg���k��v�er����a�޹�
痭��pnL�9tź定��ٴZ��P݋=�|ݰ<Pr[�����;9GV�����k�c�yX-�ӭz!D\��t*��ƶ\��VvX�{ �nSm�B�E[JuŹ�X�	�eh�uŕx|[m��z�	��a�ĝ�\��b}< 6N;A���̺geiUW�u:y8��;00 H-�{M&6�;i���-��@��m�5�8۝u��wZY���wb��m)��H�9]�Cb��h��2���٤ؠ����t[mr�n9z�e���ؖ��V�W��U�Q�WOQ��&�����Wv8ۋv���U�r�t�1����"��	/m�m��79���3.�[j�6�m91��c��v�9%��/V�xy�/l�c.�JKR��˳r�� ��9ыa+��5A��Y	x��ٚ�Թl�.�&��t��C�h�� �A���J���@��P���P:!﻽������~� $   $�]���F���w�B ��]�Θ��v�(������Y4B�.�^Mv���Ň�u�ݝ�Zd�n��z�����	��d.�4�dֳ��k<g�m�LN{,�N1���p�͝�y�[M�s�2��m��H��v;Y�t1�C�g[s�75U؛s=��=�1�h�|�*�E=���1����� �f;��S��{��{����>'	�:�́G/kss��XiژΒ�6W�����9J��2�b��M<Y$p�wu��/��Z���D(_Hv�� |���Sdڻ��E��0&��Lw�0&�A�����W�A�\����)���x�Z�7�oGL	�}ka��Xf!fcod��0&��L>�X��������Ġ�Q`��N���ھ��n����06T����:�v�SZ�qմb�g�N%l�nκy��M��|��;��ػ\��_ک���n��~I}!�� 3�uQtE]�Z������rJ-@,�B2A�(�@�k���%4s�� r���U�?L����~L$�crɠ_�~4/uz{U�z٠z��x[�D�ř�x05oK`v��LvLa�-�?���F~�s�x�r=����z٠}zS@>�� �Ա6�`�����S�aFj*�;Iy����_v����]�Wt��^�_9.M��)9c���~��cӲ�L`t��0:���!"$�@�Қ�[4����[7��Ar��~�!0N��{7$��ٹ@�8d�}f�}Қ�9a��
a1�7$z�V� ��x��`t����t����F9 �� ��4�)�r�@��S@��ZZ�Y�A���L�e�dZ�Nś�������ƛ���9K6��8�	1�܂�h���{�� ޫg�%���x�L����mR���H�r�@��S@>��ޔ�>��.2a�"S�G�[� �=$���`�1�m	WyV�S$JIHh�l�-�M �u�!""!L�V����*��J՗h�Mޔ�wY�[�)�u�@�u���m��&4/��CB�T@�T�mfٻ%G���L����
���ػL۳хЯ��Lھ��{���o�?�U�~�)�Ǌ$�$�;����2}׀{���w��L�:A�U
a䂙Z{��}zSO�fbG~���{���rl$�crbR^B�s�0y���Z��J&^�^�ߚU�b��CxI4׬�?DB�U����^��f�1!G���wzw{��_�� �-�l  X�+Ɠ4��:t>�U2�K�w��#ic94�L���O9g;����a.�u�m���*��e��oEąۧ��j�t��iՌ/FV皙�v.4l���G%I�b��n��΍�Zڢ�ɬqk9�ۮt�a-�=+<Q'k8�p(Mg�ݴ4�M��=8�5�G���og\ڞ�q=��v��Ȱoww��w�ݸ�
�p�;iX�Ƹ�
�v������/-�Y)z�ŮH�w+��5�Jd�Lc�?��~���- �h^��(Q��wV j;�QV�Q6��n�U^&�&0=; ��$��oK`z�J��MLY1�(����M��zr�S>S�� �^ |��,�)XR��D՘��|�\�����IO�����&�j��̕wx�}���B�/{��=��8�����H�s+[u����Va���#�S/M(���&�c�
p�rn�NӚ�س-�vɌmȘΙ��� ��|��r�l$�cr1�&��v����!BPD*��}xR�� o��y�Ƞ1F(��8�׬�;��?$�G�׀{��p�n�\U���WiLmI&�ݏ����@��V���s@>�ܬs�L�'�Š�f��"����7�b�7Uk���U6�� ��۹'WZ�8n&5�Ӎ[+��8��mٽvh�x����%�\�"��c�L`l���W�0�1�x�B��h�e�����<����D(�
"��Uߧ 9��x�n��w!6�j�������\������J��$��i$�I}���<X����AtU]�ں����BS/{� =�׀y�ŀn��8�ծh���NF7$���@�빠wc��m�m������.�ۗx��w3��-Y�M����85ն;з񩍩�^�}�������04�cxd�O�����ݏ����@>���蚿�b�L�)����7Uk��t(��P>�wu�ݵ�(���rU��M������ o���I1����u_D���D<-Z�V���������(IUo�߯ ��,uV���QP��QJ*�n��u
�&	�RM ��4�}V�o�� ��x�ICj��z�U̪�6u��ܴk�ͺ���!kGY�TO+Ր��զ�1���QL�Ԇ��K�0ѓVk3�ʻ������w�y�ŀ��F�H)�Š�f�}m����Z�:"(�h��P]��B�̤�1�o�}��0;��&�&h�.E���$rh�Y�n��8�n�9DB�3������M�L�)��$�;��Z޶h���O������I����?�� %�   �/\�[5-�5��m�Ԥ7]�A��{m{mY���+`�[&���OA�E�����ma���xa��q�`b2�cH�Kj9B�%G%�eWY	M^�E��p��h�"�08�nj{k��%]&]Ԅ�v9�q�qg�ѡ�t'k�%S{�t&tv��jd�<����Z[�n;|8��4�k�e��<���r�����A���|�����<�s[`:�	��,6uK/RW7DΚ�8�݁��v�r]����H�����߿M ��4^��$�/�T�p[�I�T�ڕt+�ř��L`l���W�0�1�g��:L2����h���
d{�x����7rA�A���v>�@/����h�@8.��Dcr%28����?��BP�~�~ �����Z� ӿUeKv"
��]����bck����`Zć5��S�Y��Ny�j�s�dcrM ��4�Y�wc��ـy�A�D�tU".�� 뼸�t� ��߄ءA< �Ʃ��ou�m�~S'�-WAjnT���nf���?ߖ�_[4�f�{��{���7�HB8�N-���%3��x��x�x��78��.ljb�̑E$�m���Z}l�-��6�F�(b�m �Q��S74�u��uwn]8��с�NZ��uh�)M+Dج�Sww��b�-�j��f�[l�>UlDM1�jI���Z}l�m��x������tuU�ItM]�ں�����ۼ;��iB��_B�sP�4��@�GA��`2b�,P�	A?QB���_���C�i��
"I(Q�BP�%w{�� ڦ� <���E�nF7$�m��Қj���>���7�À�r��*����0'tt���D�&ɌI1���}�C�l����h���v����\݇[(e�B �.��k|qz۶�7��Tͪ����?~U����w���B�Dz��w�X ��/ʪ�J��w7WB���	�c �L`N��%\�����3`�SFd�h����M�v� ��� ϻ�tlq��H�)&�;�8�T�p�7x�IL����D�؈� <�Ȝ4�}V�}�f�}m��Қ�^��$�j% ]{=
�j�f�.�������8�9z�S�DB��Ѹ�#�)�C@>��@>����M�:S@=�έ�DFP��誻� ��y�d�� �w� _[4V.
b�L2G&��vA��]�`�1�zI�wb.~�(���Ĝ4��M ��� ��4�w4춄sĜ�G��h�w�tDB�S��w���ل��B��EG�0u��fa�� /Z   M��9��5���j�Y��rr$�X�&�
W��l�s������ㄇu������%9i0=�=z��h<š��t�t��RX���={v&�M�y��2<���0(�P]&9n7`ܩ�n��:�c̏c��q�vt���t[�N���Wn��1�mf��5&�ω��VL�]N�n��z���\
�t)��&�Me����P�
�)��Ù�*�r݋=�QK��r#5S��z�<.o'\p�m#�s�S��vvz�%�\�%�� ���`n�A��]�`�1�g�n(��(d��$�/u��;��4�٠[f��b"h���fe0;��l��=$�eB�ո�Q�������f�}m�v>�@>˝["��f7#�h�٠^빠wc��٠��*��8�H�H%"X�Q۷Ea�����^zl*��[su6S�Ѯ�����b`Ȝ�v>�@/����hw��b�L�)��$��ݻ�iF��UHZ��&0l����� �uIY�����2j˕7s��� >m��B���n;�h�p\�4�œ"$�@>�c{��u_D�=�c �I(�.ڌ2Lc�hv>�@>�f�}m�{-�ےI	�	�B�ηVݕ�D��H���=h[k].xgm	��H��S�X㙠wc��h�٠{��heB�ո�Q���������DB��wu��b�7Uk� �;:�E�nF'$���@��wf�L �$�9�h��w$��f����@b��Ba�94w]�u_D�=�c �������X�������U�u�@>����s@��g~?Dۉ���D��Mӕ����2��_:��1�]��һ=%�r���1LĪNb�x���@>����s@���h�e*651d�BI1�zI��} �I���E�������ݏ���٠[f���$����0y�uk��RڷӀ}׀6�T(Ov�DE*U�s��ܒt�l�9����&��m]\����ġB��w_�k}� �U�pծ�r�.��ڵm�6H��Y�N����ɲ.��gk�,�l=�p/�������ӝ�]��6���ﱁ������`�1���pS�O�G&��빠wc��h�٠}x��Jd�LmI&h��� }�����=�׀k}� >[�䘞$�B'�H��h�٠{��h�����TljbɌ�wx�n�J!-o�_ ڧӀo���#����~?��    &��м�m�Uݜ1βr�㓞�mk[��q��u:8�S��M��M|3sx^�9Ք#��^�zv�[J��v[ �md���z^$���b͕:G�S6�M9\f����m�����!��v�9Mm�,.)�6)�b��L[��l�)����qMٳ�9q;W��m�8S�m���Ǯx�v�`9�T�OlW�dЀ?�
 ����z�kZɢ�e��F��]ף��"����g3ͧ�`�4�rn�*G%2LȚ`��4���s@���h�l���@��V�FҊ��U]Z�<���~JJd<�� 7{��=�w4�X��MF(��S"q��L`�c{����-�{y�D��nL�@=�f��빠yO��I%3��x��́D⩹&���y�Kd��&0�/�o��������	�nn�m]�j��ݺ����_�<|{)#Sg[�j皡��k�-]�ڪ�����{� >�� =���#��b�!��V��ͫ����j�zI�ԐuɌJt�ײ���&2I4�l�=�w4�B���wN y�^ yn���E]تꮮ�?�BIKo�Xr�Ӏ7f�z�4�bJ��ƈ&G3@0I1�l��0&Ԗ��2���]:����[++�t����6�Wh�"ڻ�5�c�������w��8���efb�����$�y��@�P�dQ����I4���{q`��8���	%'��I� R��&�D���� ڭs�����`	�P�*'���]�ٹ$���7֒�	�%2D�7�4q�Z�� o]�r�
���`���-�&(�1H��٠���������kmƱbF,hd0�%��NA�����u�&�m���޻5����BA��	��Iɠ�������� �h��,bbQc��&���,脡D�ܩ��}׀��bK��m�1�	���-��hu�@-�4[w4���1F7w2�]��tD$�e����׀y��$�@O�G-3���Oޓ�֦\�1�܌�I����)�[���z��Vۙ$��m��E�fB�aF��7���S�V�c��Kt�f��=�v��� E1)�`'&�oJh���w�J#����x�V\�s6��mSM�h��޳@-�4zS@=�ά�<Jd����"�z� o]��DD)��|`ʟN�X��)4L'�$�z�ޔ�-�j�z� ���X�651(���{l�T��m� 6��%?�`(}�yu�!t2��(�F����H+��D��"@�A�X��,a��� �)BU�Afகt��EH:Rh��D"�D�F	������N��8�Aj�0�ł������&��i*�[q�tf��#�4��DdX�FJ$DHD(@"�a&�F� ����@E$H�B�!Q ԪH�v����3i�i�� �޻����t���������    m         9!��  6�             ۽l*��6���t�R�Y�p���e@us�;Tڕz�5��d��0���M����m��n�y
vb�{b�s���7+�� �zIE�4�ҷ��n�@�\���� ���rw�v��X�d�	۪zrf�c�����kg�=�=��9y6��kt����	�v«����nqU�qڦ|��uY��lR�ͻ�mntb�j��ӈȣe�uצ��[#''P�!NͷE\Ĩ$ʧm�6� 8�l���Ɔ���aD+r��#KAx��7G.��\�V툛��wjf�p��*�CX`�s͑jWn����6�q��ݷ9 HI�i�`�va�ڮ��{	d�&���j��5�G��W����1-�3�]W0��s��v]=�s��
�gP.@=[V�:F��t���O��k��@�k�N�u�m�#]�<J���	�[n��KX�l�Hi$'@n��jj�T��9l�-oQ��W!�`NA7��Wfŭ���29ؠ�㍧���82
q�6����Ng�줩D�r�V֖i^��bn��e)���q���-6�=�^v:(�SY$��mAr�U�;vZt�T��Tʠ�gjgzNq����&̴�m�[j�V�C�{cJ[3�E��a+�]#��]� �n&mz+@ h�r��Z*��F�/�!��E�h]6�F�k 6Z'd�a�nm6y�=m,���(1 =��\�
���U*�WR�C�p�j
�/pv�%r���m�$[/N�]�l���[U;+��IU��2*cc��$�6�d1 �9ݮ��sɽ�	��SWj�I/;���A�n�;�v����mc��'r��5fv����o��vd����?�s����K���;2�l*��!���+M�,�U��(WQͩ�̺��ۚ,u�#�v�C��B"P ب�O ��|>N���o�  ��� 
�U�IT�\���{A��F�8�;�1���1�ƭ�F���(k�=� &�e٥ �cs��\�_��o�"62A�R���뜶�+���r�kq�Od�s7ۆ���0��6�'1+P��ȷ[��H�&%���h����+���k�ٕ^'gn�,�l;���5����� �������-CS��r�(������{���??%\`)烞��e�6���2������h�n�vWi�b��������<^�6Ҙ��8|��?���4�f�m���E��FҌnD�d�� m���I(Q2�׀wu�6�տ�����ă�/�Ȣ#������x��0�=ʻ� =�׀y���@LJ`�rh�)�[�Հ6��P�&}�׀n��XZ�&��Jjj��uV��?%	O��� �w^�Қg>J�	�c��G�H��,��-����gd��I�s���v�]�c&�&(�18��l��Y�wt�����h�J��M	��rIx��y*"�(K�J"�o/��Ӏ6�?%
S!��Y�RU6��Rf0$��������=:c	������ѫ�.ZL�M��S�^���8�����]��`�&Û��܂&G�w����4^��;�����Vۏ$�4܆���֥���ͮ�鹫KIPassO���a4�f6E�nF'$��Y�w[��o�k�_H�׀o;�� .mL�*��3�:`v��Ld��=:c�İ	����������[�������a��
"CP�B�6�^��� <����S5j�u6��p?B��g{�����t���}ռD<-Z2��yRM ����w4�>�@/[4q���	�89�S�"Q���^�i���ۜsHlm����ӆ�����%�lU$���s�ŀo�k� z��׬�>WU���I�L�;��&:L`�1�:GL�I��e�Q��`L�- �l��Y�^�s@�c��:�E�nF7$������ �*�8�/ءD�	E��� }��G 6�mH����x��s�䤅$)��y����1/�wٴ�Kı>����kY2j\�t���\{7j���jζ�v6X�T�˹��I� �R����w����Y��bw�;��Kı/{�fӑ,KĿ��fӑ,K�����"X�%�~'{=u0�-�e���.ӑ,KĽ｛NC��&�X���fӑ,K������"X�%�ߌ�ӑ,K��|zz�d�՘Lu�Y��ND�,K��}�ND�,K�{�6��c�(�MD�s��iȖ%�b_{��6��bX�%�����I�M\%�j˙�ND�,K�{�6��bX�'~���9ı,K��ٴ�Kı/�wٴ�Kı?kŷ��Iu5p��M\�iȖ%�bw��ӑ,K��｛ND�,K��}�ND�,K�{�6��bX�&�E��{�fa������t�  ��ԗAUK�q��N�rε��i����q'�m�8�:�ݯM����4���9Qֲ�4�\Ju�ΠW�B��n*�<F[�����Z�W�Jy�qk�$,ekK���3*�fz��=�u�ڣqۣ�츼�o<u����9�+�b�U{2pc��ۣS%��;p�Y�����W^��pm�g���n�kD���MC��E6�Ho7�kY�ԭƧ^�:"�vUCZ��i�f�F�nY^�u9�����v�ִ؝ _��x�,K�����r%�bX�����r%�bX�{���Kı;�w�i�����v���#Nw-9j����bX�%���6��bX�'���m9ı,N����r%�bX����iȖ%�b}��V�jI2�nZ&\��r%�bX�{���Kı;�w�iȖ%�b^��ͧ"X�%�{�ͧ"X�%�����Bar\3&���fND�,K�g}v��bX�%�}��r%�bX�����r%�`؟{���Kı/��g��E��	��u�iȖ%�b^��ͧ"X�%�{�ͧ"X�%����ND�,K�g}v���oq�������*��8۫k<�K��ʍUL[�۔*p=�\p�m�9^�M�۳�VfMkV�1�]ffm9ı,K���m9ı,O��p�r%�bX��;��Kı/{�fӑ,KĿ|K�=�5����Ys3iȖ%�b}���Ӑ�Q?�(dL�b{?�v��bX�%���iȖ%�b_��iȖ%�b~׭�ײK���.[�.a��Kı;�w�iȖ%�b^��ͧ"X�%�{�ͧ"X�%����ND�,K�}�R��j��ֳ!&fe�r%�bؗ���iȖ%�b_��iȖ%�b}�{�ӑ,K����]�"�oq�����>��ӝ�NZ�{�7�ı/�wٴ�Kı>���iȖ%�bw��ӑ,KĽ｛NG��7��㿟�������)�.�nK-���4��ᗮt61][su=+ƫ�.yT!�L�[�։�36��bX�'���m9ı,N����r%�bX����iȖ%�b_��iȖ%�b~�f���\�ɢ���"X�%�߳��ND�,K���m9ı,K���m9ı,O��p�r%�bX��w��S	��a��\�˴�Kı/{�fӑ,KĿ��fӑ,��dDu��N(#�M���������Kı>�=�v��bX�'�羜�u�[��Yu����K��/�wٴ�Kı=�{�ӑ,K����]�"X�%�}�{6��bX�%��/d�I�M\%�j˙�ND�,K���m9ı,N����r%�bX����iȖ%�b_w�ͧ"X�%��{�ֵ6�͎�vzsQձ�����l�ʖ�tV�-��/=�BmmU8r\q�W|�Ȗ%�b{��]�"X�%�}�{6��bX�%�}��r%�bX���o~oq����}߿w��9���Ȗ%�b_w�ͧ"X�%�}�{6��bX�'��p�r%�bX��{�~���7���{��ݿ~�����[ND�,K���m9ı,O���m9�,K��z�9ı,K��ٴ�Kı>�w�g�[2�n�,ֳ6��bX�'��p�r%�bX��{�iȖ%�b_��iȖ%����LH���ٴ�Kı>��~�L.K�d՚ˬ�iȖ%�b{��]�"X�%�}�{6��bX�%�}��r%�bX���iȖ%�b*�������vN[�^Y飞9ژ���N���>Ӿ�J�k0�Wg��g/�{_7��g�Xe�&fe�}ı,K����6��bX�%���m9ı,N����r%�bX��w�iȖ%�bt��N\�֭�a��Y��ND�,K��{6��bX�'��p�r%�bX��w�iȖ%�b_}�fӑ,KĿ�%�Ԛ���ܦ����r%�bX�}��m9ı,Ow;��KKĿ���iȖ%�b_}�fӑ,K���[}��K���.[��̛ND�,K����9ı,K��{6��bX�%���m9ı,O���6��bX�%�痢��չ��fBL�˴�Kı/���r%�bX����iȖ%�b}���iȖ%�b{��]�"X�%�P���{����?����    4�z5��^%��ξ1�]:yȕ�;0evv����Hu���Y6��w�:�#O<�	K�wi�ۊ�Tq�Gj2s�g��2U�Z��i-˛���.�/3ד���*�X����:���+�6/��o$���d{)�2l�c#\�sY�ݢ���&ܛ�'T���9N(���p�ک-��%�+���=�{?����{����˿����y�qC�W9Y�N��GT�Z&u9΍1	G6ݞ1��˅�Z�Y�����Kı/��{ٴ�Kı>���ӑ,K��s޻ND�,K���ͧ"X�%���wg�ճ.᫢�k3iȖ%�b}�}ͧ"X�%���v��bX�%����ND�,K���m9Fı,O��߲��5f�����Kı=���ӑ,KĿ���iȖ%�b_w�ͧ"X�%��{�m9ı,K�׾���an��3Ff��9ı,K���m9ı,K��ٴ�Kı>�}ͧ"X��5�����ND�,K����˗ZոL52k33iȖ%�b_w�ͧ"X�%��{�m9ı,Ow=��Kı/��ٴ�Kı"���~�*����3؉ĺl�3���i��cq1dx�Dmi[�0N�����sZ���$D���&��	ߵ�݉">�q7�,K���m9ı,Oޙ}��K���.[�sY��Kı=���Ӑ� .�C�?�uq,K��ٴ�Kı/{�fӑ,K�����i�"�bX��㾶��K���d$�̻ND�,K���ͧ"X�%�{�ͧ"X�%��{�M�"X�%�߳��ND�,K����Z�p��]k0�36��bX�%���6��bX�'���6��bX�'~�z�9ı,K���m9ı,O��ݞ.��p�].fm9ı,O���m9ı,G�g�v��bX�%��{6��bX�%���m9ı,O�;���]C6�2���p#T��닋�c|��"���:�0W<����ud�5��O�,K��s���9ı,K���m9ı,K����r%�bX�}��m9ı,K����S	���,�33.ӑ,KĿ���iȖ%�b_��fӑ,K���ߦӑ,K����]� 
�bX�|{�.��p�jd�ffӑ,KĿ{�ͧ"X�%����6��c@��? |DaE�0�� <|�l�h�B;�A(��`�`Á
D�I(��HB��h!�*D�(d�< �(t5� DՊ@� ŀB��F���B"PB0Q)�� ��ЃH@"AbD):b#H0b�RQ) �l+Q#Dt$A���Q	� Oͫ,�BRIE�FA�$HŊD�"D�H0#�,(Bdj,a�,B���B��BB��mA@(�(q�$TA��@pD�
B,@�"&�<~����7��r%�bX����r%�bX���zk�&�j�nS.kY�ND�,K���m9ı,N����r%�bX����iȖ%�b_��fӑ,K���[}��K���.[�\�iȖ%�b}���iȖ%�` �}��r%�bX��}��r%�bX���iȆ��ow�����8�[�Ւ�:��4ef��l���=L�^��C�F;/��u�֭�Mk2�̛ND�,K���m9ı,K���m9ı,O��p�r%�bX�w���r%�bX���u/�����ֳ-�ͧ"X�%�w�ͧ"X�%����ND�,K��~�ND�,K���m9 ,K����[<jٗp��r�fӑ,K�����"X�%��{�M�"X�%�{�{6��bX�%��{6��bX�'��z�4\��.�n\�iȖ%�b}���iȖ%�b^��ͧ"X�%�w�ͧ"X�Lt��'}�p�r%�bX��{�50�[��f�32m9ı,K��ٴ�Kı���m9ı,O��p�r%�bX�w���r%�bX�zL���kR��kZ�N�xLZκ�fc[��l�tZ2��.k����v�ù��tB�v�}U|�~oq����?~�6��bX�'���m9ı,O���m9ı,K��ٴ�Kı/�ץ��ֵpֵ���k3iȖ%�b}�{�ӑElK���ߦӑ,KĽ｛ND�,K�｛ND�@�G{�������p�����{��ı;�o�m9ı,K��ٴ�Kı/��ٴ�Kı>���iȖ%�b^Ϗz˙�[���d%��6��bX�%�}��r%�bX��}��r%�bX�{���K��T"�j'}�M�"X�%�{;�K��L�\ծ��nfm9ı,K���m9ı,O��p�r%�bX�w���r%�bX����iȖ%�b����333333333�  Mf��&��碇�g�عQ�%�`7��4�(s����dКu�i7���NI|��=m���m:[��, 1�.$.�8s1H��y�a��v�φL|O�<�P%m��Y���9-[m�m����L�v��k&õ�s�����N��ʧ��m1�R)q��Z�{G(�$��t�v�нC�ݸ�%@N���k�v�а���ϊ�U/lX�aI4��f���g0j�:..�b�&�6,�mKR�a�f\-�WE˙�'bX�%������"X�%��{�M�"X�%�{�{6��bX�%��{6��bX�'��z�.K�d�Ԗ��6��bX�'���6����bX����iȖ%�b_���iȖ%�b}�{�ӑ,KĿ���n�rI��iȖ%�b^��ͧ"X�%�w�ͧ"X���Q5����6��bX�'}��M�"X�%�����.]kV�2�4�ffӑ,KĿ��fӑ,K�����"X�%��{�M�"X�*6%�}��r%�c���}?x��p��-|�~oq���b}�{�ӑ,K���ߦӑ,KĽ｛ND�,K�｛ND�,x���޾��v
]�rF��&Q��C/X�z{b���X�t�(֜�%�K it�Թn��k�"X�%��{�M�"X�%�{�{6��bX�%��{6��bX�'���m9ı,K���Ys5�sSZ̄�3&ӑ,KĽ｛NC�/�� yT��x��%�b\��ٴ�Kı;���ӑ,KHZ�q��!I
HRB�5��T\қ��Z̷36��bX�%��{6��bX�'���m9ı,O���m9ı,K�wٴ�Kı=��V��e��5�K�36��bX�'���m9ı,Ow���Kı/��fӑ,Kľ｛ND�,K�{�y՗%�2M.L�M�"X�%����6��bX�"_{�ͧ"X�%�}�{6��bX�'���6��bX�'O�7�atj[��7g]h���tjXڢ(�Z��n��ûRn٭�]�[�1�i��g����W|�~oq�ı/��fӑ,Kľ｛ND�,K�{~�ND�,K���m9ı,N����˭j�&]f����r%�bX����iȖ%�b{�o�iȖ%�b{���"X�%�}��6��%�b_>���%֮Z���fm9ı,O��p�r%�bX���iȖ;����;�fӑ,Kľ���ND�,K��'u��j�K�Z�n��r%�bX���iȖ%�b^��fӑ,Kľ｛ND�,K�{�6��bX�%��{�\��sSY�H[�m9ı,K��ٴ�KıB���m9ı,O��p�r%�bX���iȖ%�b{G��kZ�f�j���#�civl��B:gjq����M�gcy\/7XZ]J�������2X�%�}��r%�bX�{���Kı?{���Kı/{�fӑ,K����oƵf\-�ZԦ\��r%�bX���iȖ%�b~�}�iȖ%�b_w�ͧ"X�%�{�}�N@ı?w�םYr\3$Ѣ�a��Kı?{���Kı/��fӑ,KĽ��ͧ"X�%����6��bX�%����0�-�Y.Lֵ�ӑ,Kľ｛ND�,K���6��bX�'��p�r%�`hZ��D|�����ND�,K��g�.]kV�2�4�ffӑ,KĽ��ͧ"X�%��������ı,O����iȖ%�b_{�ͧ"X�%����߲���Zr���۟Rq9y���2��u�Ύr�����f�7/�];
\-�W5�ͧ"X�%�ｿM�"X�%�����"X�%�}��6��bX�%���m9ı,O��;�՗SW
\��Y�ɴ�Kı?{���Kı/��fӑ,KĽ��ͧ"X�%����]�"�bX�%����.f�njk3)2kXm9ı,K�{��r%�bX��wٴ�Kı=����Kı?{���Kı/����f�2��j٩��u���Kı/~�iȖ%�b{�o�iȖ%�b~�}�iȖ%�� �D�����ND�,K���K�kVe��5�K�36��bX�'���6��bX� ?���m9ı,K��ٴ�Kı/�wٴ�Kı0�~�{�w��~��8 h ?���̖v�XW\�$i����A-ېڶ<=�5�2���u���8]��Rl-�k�hr.΄lm88��1p�]q�:�]Ӫ9.y�4��EÜ�5��ލq���إ��i�"Z�U/:Ɲk���T�۞���W8��1�)J�<������$�q�QGgm�8fx���N\3����*�xṸ����*�E�p�ռ�I��53	���9��q�tݦ��Vc(�܉�gU.�V����l��\��2M.�̽OD�,K�{�iȖ%�b_��fӑ,KĿ��a�
$�Q,K�g���r%�bX�����I��nɚ2�ɴ�Kı/��iȖ%�b_�wٴ�Kı=����Kı?}��m9ı:w�ח.��p�u�s33iȖ%�b_�wٴ�Kı=����K�E��j'����ӑ,KĿ���m9ı,K��=�.�p��h��k3iȖ%�b{�o�iȖ%�b~����r%�bX���iȖ%�b_�wٴ�x��{���?{~��K�!c5�{�2X�%�����iȖ%�`�}��6��bX�%��}�ND�,K�{~�ND�,K��w�ֵ�&��
L�	e��Fl4ݕ�P�nMr�+�k7k���d�lv�5�8�	�Gik|�~oq����}���m9ı,K���6��bX�'��}v��MD�,O���M�"X�%�����W�:.�3��{�7���{�����m9�Ȉ~>� ���,Mw9��Kı>���Kı/��ٴ�Kı;��T�5�2�n֥˙�ND�,K�{~�ND�,K�s޻ND��,K��ٴ�Kı/��iȖ%�b~�_>���ѣY�Y6��bX�'��v��bX�%�{��r%�bX���ٴ�Kı=����Kı/�}�a4[��f���v��bX�%�{��r%�bX���ٴ�Kı=����Kı?w=��Kı/�{V�F]K
�4�an�͕��}���VGm�y��;G)ۇ�gY;���^���]�t\����Kı/��iȖ%�b~�{�iȖ%�b~����r%�bX���ٴ�Kı/�x������Y�W5�ͧ"X�%�ｿM�"X�%�����iȖ%�b_w�ͧ"X�%�}�fӑ,K���I�fYu5p�˭e�Xm9ı,O�w~�ND�,K��{6��c�A?�%�b0d�dHă�P��D8�dO�.����r%�bX����6��bX�%�����P��v���w���oq�׿{ٴ�Kı/���r%�bX��}�iȖ%��!5����iȖ%��{�����t=(nZ
�{�7���%�}�fӑ,K��{�ND�,K��ߦӑ,Kľ��ͧ"X�{��;���>�[j���r��Ͷܡ���n̽s��Al�Mgd�I��r������_�j̸[���r�fӑ,K��{�ND�,K��ߦӑ,Kľ��ͧ"X�%�}�fӑ,K��ܾ}e�L3	�F�Y�6��bX�'﻿M�!�D�K�w��6��bX�%���ͧ"X�%����6��bX�%�ｒL&�p�Lі�M�"X�%�}���ND�,K���ͧ"X�
,5Q?���ND�,K���iȖ%�b||x߲�j�&f�D��fm9ıA,K���6��bX�'��p�r%�bX����6��bX�@( |dMg��m9ı,K��?��Iu��ֳF�SZ��r%�bX��}�iȖ%�b~���ӑ,Kľ��ͧ"X�%�}�fӑ,K��ǽ�kZ�͹uq��g�N[˴�SR���:���8��Gi^9�ι��j0�����%�bX��ﹴ�Kı/��fӑ,KĿ��h��%�bX���~���7���{��}��'3��x�Kı/��fӑ,KĿ��iȖ%�b}�w��Kı?}�si����wr{��7����/��Bl�Y�ND�,K��fӑ,K��{�ND�,K���6��bX�%���m9ı,N����Ƶf\-�ZԹs3iȖ%��6'��p�r%�bX��ﹴ�Kı/��fӑ,K��������r%�bX�{��YrS�VkY��m9ı,O�w��r%�bX@#}�{6$�H���7�N���ؒ	"�*
���*
���W��V��*��EAU��W��W�('�QP���P�AP�(�P�D�� `��AP� B E@���  EBEa T$AP�DXDBE$P�B
B"DX�0B�AP�����AP�B(�D
�P���`��(�B0B1BA@T"�BT"�P��B�B(�B*�B �P*B 1B*B*P
�AP�� #E��
���AW�T_"(���A�
���PU�EAU�B*
����*��"����W��T_�*
���PVI��u%�B {t7�@�����d/���2���,���kE� YX-�Q�Ow� zIE/Z�@� P�  )R  P ր����F���@ ���|%��Q���i�=�>��-�태'ptG�{5�       � �=N�հ·C��442}��p|O���$�͝M�t
 wWz:i����4|3��C�q�<$4��Q�}���h(��}4q��h!�ɻ�{�k��ѧ�F����
�Ε�C֛�t���ty�pPhh �l(S��z��>4P�
y�����O�����AA��qpkӣ�;:9z���ᡠ��C�(yz4:�� dP�w�W�+Ѡ�AqW�h47g�����B��������4�]����î�rhz�  @ @ 0��%*�����&�����R�=MS� �    ت�)�R5       ��U$�*�H��  z���  "�I �&���"4ښѡ���L��@� M	��z�x��=� ����?H�/��<.U�����r�(B�� >
�U�#�����K���� �lQD �a�5�l](��J����
 Ry?��G��O���_I�}7ϧ9�}�A �"`C �� � 9 '� S�/�T��O���� � #� ���PO��'� 䢡�QS�&�~H�|�;
�v ; �` ��w-�{�ѻ����Z�����̼���{�����{���y�s�Ә{����/���������������9�˻���˽]��{����ٻ�wwwy���w�s�����7ww.��7����w�z֞������n����n������y�fe�{ۻ���fb����X���g��x*�ϾKM��O����s�:�/���"���C��=.?`��?��Y�K�&�4�2�r��w�p���	�1�<޴�����<�e�JIM)4�t�Qo��3�l@��Mw�o5��4+cZ�Q�zR�`��%SOL�PQ9M�
!�Tc�����)����Oxтkg
���0:v��4�F�i�9 Uaj��^3��|�^�a��O�@�Dn;��.D�B��ސ�4���[ћ��� #�J#"#�1�*���a
�*�!_�Dz�CH�b��˾�4ba�OIBY�����efXIa%	\BW�!��#4ƌBD��HN'���}}4�!��,`Fj���N� d)�M���M%�2k	
���bgE�2U�IM��΍c�IE��`ΫAP%�A�7d�2h�0Y�m��(�C)Q�!� �/�$-��3F�4Y���<*<��y�]n����]1#p�Fh,�Nk��U��5��\���Ყ436���0#0�@[�$��a�+a�0�8��`q ���h��GHɘ"#N� �ݤbhcqȬb'M�E�4^
���qi�Cl��:�᠚D�e��V�dhȃn2���u�:�������~�dg��t|�2�q�
l� ��s;�Uɇ.� �	�����A��l��#�7�y�k~:x�Bo��sD�<Mվ1���� ����ju��p�I���ѓ�`%��:	a&���X`a����dL\CJ�$�xP�=|�4mt0b�b;BRt�2Nh6����������L��cKv�:�i8`ewX3�F1zH&�He ��KaВN(r\to����\5�q}'@�B#�XCA����I�E���7$%1:��ڛ!x8�D����aH$f�*��E�g���0��zl�HE�,�@���Dk�c�gl�;��i8���:rY�F׆s�$a�6aȺ%)ej��äf��b:ټxS�0!�&��8uX�N�0�&��k�Co����:k||�KӸ�Ѣ	b	'�&C@JH�!���y�������`��d�b%%a�B�,'%1f1i����l�,�kz �9�f�t���@|u��q�� �Sm���H-hh'�hG��jo{{�	����
����y���V��x��C'�$"�
S�ZC���l�ƕ������eo��.{�����,����e�/WŇq�PA�m���L��q� Ӻ�B�['rh Ѩ���D%�M8�����1H �Ƴ0՚�i*��
h�P�����P�oz�y�V�UWRVs΂	�P0�!�D���#í���NЌa�q,;H0;�A�%�����o�:�x���͘�,ӆç3q;:ٳ��kV��p�gO.�S��Y�|�ӺvֺY��ӭ����F��zn<#	������I,kda�%�V8���el��mc���o�И�K�/C��y�fK��,�'G��F����u�"+(C�F���SV�DH����oF�Z݉�Y�5�4��	 <z�I	�K&�q`�! !f\d�%a�HF
h./�.�&ǩ�_}��'�l�><OF3�N>!��H0tN&'0a�`"�� �A�� ��B@lxt�!�4)�	��14m8��hv�H	';^,a���hHq3�E�'�ۧ��'�f�6q�k0Y�D��x����(h�v �n9�|���0Ӱ��E�NX&˂oU�0��5x2d�02Q�cm��	2h�:��`��d�9�]U%�UM�T7ad�ucՔv?5!�Bo�T)כsB����ʶz������HU�~�Pq�rZ��M6"c癉����[�I�ck7�焤~(����`��|��m-��\���H����$jHމ�T?���R��|��l���D��͐C{��q�����}>>        � �    m       6�	� m�l              ��                                                 0�}�9X&��䭂g��wg'm|���l�i��ŵ۶-��� � ݙ0o���� ��*�d�éZ��a�tL�bXi;H$��Hv7m�m[��m����i-���[�Q�L�@OZ��2~�z�-�� ��  m�l�Ұ�Ö�ķm�I��1���
{+��R�� � 8 � �6ؗ�y;U�@$�O m���F�Kn���H�v\�m[M�@ �	ll��eT{2��U6�^U��g��[wm��H���X`u,��Ll�[l[R6����m��@���m�E�	�����m��/�i2N�Ӫ@�nn�US���p�+W)-��S`����]^yPL4����\g
n�(��n�ݶ�x�KXˉ��cHі'!��p�  ��ݺ�UZ��v[D�=�t;��Ԑ �s�$0\�t�/6��mT��m6�H]$��c���Hڧ7[n�m�p�� �'�z  ]� �^�$�g[˱4�;mW*�U �Ƕ��z ݤ��� �-��m�l� m� 	 p8h$��l5� ��m���FҫlH [\$ ������-����[@�� 6ۜ� �h �-���M��x3^^$ V�kn $�� ���i��ٻf�H�ݶ�t�D  ���j�	W���l�՞%��I&��o6�(Rm�m&�� 8j��+�ؖU�j�z��UJ���)���-��k�'s1��nЫ.�H����q��f뵵!  ��7��   k� lٶm��8�` ���v�%�K��0�}���=��}	  H�06� �;6Y,-Sm�j@�[lz��m:Tu��d���K�cvKu�,���R�`�[Uu�� ���mmηY.qr�ٶj� 	��/Y�fŴI  � m�   H��(�n�C���V��qrq�����U�hL-Pkp H]6Ϋh�A�.#��@\jj�
5�@'C� ���	 I����R�<���n�i<���l$ 8  9k,Y�*ډd-.�t�,�D�%I�/Cmm-�L�l�gI)sZI����	2 �k�;n�mm��mKh   i5-9Ͷp�9�H�u�u���l���ۭ�[y�'%�g��mo��6٭cm� W�8����B�l�T�j�i�I���$ �`�րlrKol�m���F� p�$:ս�E� �9��ٮ����%��A�U��-PR�JK $� 6�` |/���m&����6ؒ�"�x�H��V��ŀ�T�ʎ�e��� 
���\L��6@������m[@�
�R�U��l p&ݬ]�l�a#�9��Y��m[Hh''Y@ 6�[D8�$�v�H��t�-��Qm���h �  8 q��-� �N�M���xI�eZl�7�k�  ��n�6ص��n$�  l�&۰�Kh �[%�m�t����A� n��� �n�]-�i6 �@$	:�	����i6�@    ��F�5�H �� � �[D�-�  �  p 6�-�M�[C�zK/���-�i�Ŵ� [I��l�@t�kW���&����u�al�zA��Z� ��[@�I���++UV���sOizg( ���m�ඛm���Ͷ  K(z�m�m�� p$m�-�趀 m   -�    m� �@�` $z��  m��   ����� p$ ��`��,�l  v�/Q"�	��5Ś^��W*�n�* �k�Kh �۴�і�4�ְ��Qu@ ���X`9m6��$�YD�j�nI��m5�m� :��Idؐݶm� �kX F� �m,[�m��ZHҫ�\�ζO(M���N�l �V���%U�I���^im��  7]�$$m9҂@���������'ZK+2j� �k���#�0�y�inS�2u�	1����* �"	�"����\�U�@*���?�5h�
�ET��b��)�{(��Ih$���,hH�rʊ�*(k�E����"�,���Z�@�B��#��zE~@#�訞�E�6�,������tD�D0�HqDU��@ ��\(�m�hD4.��%`AiAL����lE	GH9T�&v(s@mEp� a@x	�z8 H@�( &r
�A6 ��� #\TC��l��@2R�>��g�����Ј�	dR� �A�T�BI <�A�*�U�tب���[P�(�@9P"�"�&�B��t��NK��� ���fu51SUUUS53UB����r*�����򪪪��*���������*��dUUA��  *�����<���������<����������<�� ����J� ��`qBG�7��~�s����f���x��w�$HH� �[�ws9���Y����s��s���=��|-����Cͻݧ'|y�W>> l  ڶl�  l        US�7nѯT�6Փ���/��Pe�Rm8�)F�a�	P[;�5�)�v��ƫ6ws�"���RlbP�ѐhKq��YwgMS��p��B��
�ۮ;GZ*�^0b�����܀Jn�i���Ĭ�..ЊN�:��S�D ;Xp�{r�p�]϶�Ä��{u�s��)k��ۢ�f�6y����(�lJ��z��i�P\�.����:[OJ���k�K�#OOT�<�j�6PGgV�r�)�쫗CǍ��'nm"�Kj��T͖vL��B^h��U���L�Lag<I���|����vۘM���^��]c���F⮹���rAmUr@��X�v�᭕u��X"Γ�y�ۑ��f�[6f���vl���%6i�3j�#���#�9��`�'�i��jMGMv���jt��B�K�R��ʽ�j���V��d���	7�)��3Ug�0��	\�Ѝc[k*�&���64����.�h��������j������,+,�i@ñ4�X(m��w�/˯�_���󷡶�7%��a.s�2	��&ֺ3L�Z�q�C���sŮM�W%˃Pb�j���v������㇌��f�	1�ɊG�ӧE�N���͔2���/W*��g��O	���ۺO�>���Ŷ��YI���SWM�Km�StP����Pl���׏�t*��α��Yw�[&#Cz��:�5�,��cOh�Uwl��Y]�S�$*��c��b��k����E�d��wlO�=����z&��a��::W5�[W[ �mqTk]�'�>i��㫾�d;{Q���wo�B���@�F)� �����w�p��`q������wl]۫��{L8���[b��]����l��Ho1�k��:��W{��bG�+�m��Vz;z��m�r�1���ݺ�v��
퍑�tX�%�V��4��w�Z�.�f%�U�K{r�Wm�ݺ��Ȣ�6cU��7ͺ�� 9w����ݺ�zY�v�<:�H��[�έ�٩\m�{b䪨[�@�)GWv놗m��`^��4�Y��1���X����)���1�����5r���1�4.��{�W�!�EGPL��X���f�]ܮ�nؗf�`�Yޕ��2(���K��ذ=	����z%H�1@b�gU=�ͺ�������kWlk�䫻.������ҍݺ�y�Vi�\=�
J09v놕���+�7��7dU�35��A��{�㽠^�t�9B B��C���$�� �!��}y?Q�  ,��d5��N�<j��2W������FN#�d�,M����7��Y�����N���t
b�)�3��b�T�(�	��H�U�.:�}7��~j�b��Ӵ'C1��uN��p���6�s �ߔ���|�t��|'������=
�r	�r�{ ��Ҧa�����fɹ�\s���riG��r ι�M�\�7�^@-f�G�����G9�j���ꈸ�9H�s�
��`Up�U,�VR!���܆S7VXM��.��3d�"-��U�L�Fy�P.�n�y ��P-���n��*n�y�P�RDP��"k�)G��`S��sEQ5�^@,�9�^s�|�(ߓ��kU��>�,'�~�G�=�/߾�%��N3S�s���!�9@� U,�6h
譣�n$�i�IF����j�Zl1 �5جg�k�M眠]@,�r�o�&,��.bp�� vQ/[����h�����kWW57U7Q ��)G:� M��\�p�����37QwSxQ��@�ި���(�o�&�.������&��uÓ@�9�9��V����v@q���j�n\�$ɉ�
�4*���]����Q�'��&*�"�{�Ҏ���u@��<AH@�:NuWS�^����{ ��P-�g��&�y��.���ùڢ#˺�s��e͑s�^@.k4��9Ƞ^sT��Fusy��6ni�[�#��NOH�l#B8�1�ل
�ݺ�Z����P/ ���5uu31xQ�9@v7�и�{ �;���3���E�7@���P��ҏ9�@�	ȝ��ɛ����qY�s���&�>Oq�LUD\�.u�Q�uJj" ;�zN䓻w|���|Q��UUUW:^F�;	jS3�0R���7M�V��˺�I���=�t�v�B<�Ez<���3�t��ݭ�j��u��=�瞫*gk\x{<��j�J���S^=3��v��`�]	Q�Z�c2b��ؤ������Lj��Wv���x����@���"�fɹ��
s�@��^W)G����p�.ɹ�/!5�ڏ9��5J8�uu�]T\�<�kT�kV�E��3WQs3u�s��P�����Z�)Gy��Ȋ���$.��-��wduƮ�:[���|�����\s��E�r�y�P/3�"ɨ���/ Q) ��R�9��7Jr 1���Q0���u�R����^@//��1u7�o���^B,�z�"��f�y�P.�y�Q�9J�	�
&�F�]��X(D�l�k�b�16��\Ǻa�V��������t�'�h��(�Y��uU ��(�(g{�y
�yH����殢�n���r�u�к�P�������W�k>��<מs�4������D�M1R�Q4Rbu_���&�H3d;Q@�)a
��+ �C蛦2`�"���	=O1��BL��4�.��緲���҈��`�	���� �hD#`�('��cYS�Ѳ �T$��tBH�߾J3j0(��|���{!�:��I���>i����ߖ��t^k�Gp4|��P�������C�� �D	�%	BR�%	BP�:~���{~b|P��!.�%6���r�`�l��ʸ�=N�:J��(J��"��)J��(J��J��JϿw�(J��"��(J��(J��J��(J��(J�=ٱ(J��(J��(H��(J��(J��"��(JS����J��(H��(J��(J��"��(JR��(J���	BP�%	BP�%	BD%	BP�%	BP�%	�%	BP�9���V����(J��"��(J��(J��J��(J��(J�ϛ6%	BP�%)BP�%	�%	BP�%	BP�$BP�%	B~~~obP�%	BD%	BP�%	BP�%	�%	BP�%	BP�'�0J��(J��(J!(JR��(J��(H��(J��ϛؔ%	BP�	BP���r��(JR!(J��(J��(K�>}�{�ن�G�(J��)JR��"��(J��(J��J����>�>�bP�%	BD%	BP�%	BP�%	�%	BP�%	BP�'�`�%	BP�%	BP�$BP��	BP�%	BP�	BP�%	��w�(J��"��(J��(J��J��(J��(J���fġ(J��(J��"��(J��(J��J��(Nt�=�����z%	BP�$JP�%	BP�%	BP�	BP�%	BP�%	B|��(J��(J��"��(J��(J��JR��(Mw��J��(H��(J��(JR��"��(J��(J����͉BP�%	BP�%	AC�%	BP�%	BP�~���x|A'��)BP�%)�}�ġ(J��(JR��(J��(J��(J��(J������z��o8%	BP�%	BP�%	BP�%	BP�%	BP�%	BP�'>�bP��	BP�%	BP�%	BP�%	BP�%	JR�@}�J*������wN��%��ī!H��]T0�4V��\ݳ�8�+���%	JP�%	BP�%	BP�%	BP�%	BP�%	BP�>|�ġ(J��0J��(J��(J��(J��(J��}���%	BP�%	BP�%	BP�%	BP�%	JP�%	BP�3��BP�%	BP�%	BP�%	BP�%	BP�%	BP�&��{��(J��(J��(J��(J��(J��(J����͚ެ��P�%	JP�%	BP�%	BP�%	BP�%	BP�%	B|��{��(J��(J��(JR��"�,��s�B=�i���d�E��NB	�A�j���� �����S4DXa���(@C�n�o��0��A�0N3E�G���No�!p���D5�w�M�&   ;m9ۋ���-�H��O���C�rt��qU�ܴz�-��ېm�nl��0���8m�cBP2�z�f���B�w=�{b�Ԉ�Ԗ���VM����x��ONZ��*%�Cf����C�/��d��ѹ�;����Z��_;*=�h��Gn".ɹ ��G��؇s�Q�{��ʹ��A{�Q�f��(w���-w�M�uu������=�f�eZ�n7���WQ3e����P��ʏ9�X.5�IUS5w�ӱA��C��!^J��D��Y7sxQ��sI�T�{I�EX��v�s�S4DZ/�r���;J�hX�(�� B���".�f���I����w�о�G��d��2%��U�̂�hP$
��T+3-�{���]�s�B̨�jﮨU�|"H�t�,�\�&*3�J�c`���d��{��"���iG�	���U6U�E�G}��{��`9ؒ��|�͕uM�/{�Q�+�_P�*��>L���Q ��u]�&�.o4�u�;#6a�>2�L�Whk[`e
�dk3{[,I"A�d��I�2CD3[]�噕@rC3w�b�x���.%f84s1���C3s{]6�@��Y���uwlo{V ���uv���]�uA��ǜ��5������u�5v�a&ݘ�A��ջ�g<-�eф׵u�QĠq�����:k1�uÛ�Q����0�=
�c{��\ζ�-�;���9�Y�c��G[&%!л�0��ÜU��K8$JW����t�bv��hr���u�m�  'L�[R�At���wJ�x�l��8v��c&����V��v��{cE����� ;R+��V,�.
ͨ,�95�W���9�����qd�]��]]�lیy7�;��ry��R&�C��@s���{n�=(�4�����[?�!��u���[� ���V�
\��c;͸ˌ���̕(˱�A��%��]�5v��cDf�oF"oKGc:�G:�sx��boo;�:Iĩ3r#n!��Ҥ`L��v(�������Vf1��b:Ht.��� ��̐x׼����@�``��:G���/{Ҧ���E��U�-�]�]7��7�`�	����ޝB=��Ʀ�yȑD*����-�-�n|���z��Q)e�L���X9w�T�o���RJ���(������{[����O\k|_ �e
�[���ۯ{��yƓe^Ň���c���q��#C3w�bϧ�}���}9i5�&�+T��B4٣@�Mh���I��>��:k1p�c����D Qh`5������kv �FsL�5�:�fA���b�kz�|>|������>�t�!Id"EM�d�{&cY�ŗu37N�����{X�Ձ�s�$�L�P�bnp��\Gd�Z�]5����Wv�_l�*�N�>:��A�Uz�v8j�:�zŚ�X{��X�(Lh�c5��«���9�á�(���8�f:��?�zn�����}�9�s:����s�퇀��JL}G�q'��Z�&�|��I�A&6Y`X�A!�eX1�Ԕ��"	�B��HL �lD��]�d����!�2�q I\�6N3L��0�l�l��D�L:�h�0&�D���a�$̄�A�� ��b A�	`t).����^�=�{��U*g7B�g^��/�О�ʪ�� ? ���            .:ڕ�u�aFh�[� �b�ȉS0P�m���H�,�ZPJ�,�mnٵ:}�3m�2��&u� [t"9DM��`�;n���=pL�`���]�
����j����m%���n*�0s��P�)��@�1ב^z7#l��ԦR�ѱ�B��ԁi�θ[�̈́6�u�36���e��v+b�f�� U��QpL��U�
h
��2v�p��dvP����0:�{�ҶZ�AͶ鲺�bW\l�G����Mjv\v�G8�)��l݌f�t@,[m�G\T�wg��.��Yv�G�"�ݻa��z��GRs���+�f�ޒڮ��=u:[���F���饨E�V�����Ӝ6ɱ[o15��и��m�]j�9����)O<�[f�n[la�r��:%�ԤKH(���%�[.�h�h�����.�o�ħU*�\�X��Q��"mZꋊ��������,���DWl6(��T� m]�D<�"'����r����F  _:N���r�-�[��4q�uZ�ym��L*����m�)$mң�-T����|A�]-dq:�e�{��ݱ��Iux�i��O.Uԭ4B�j�M��t���Ⱜ0�Z��<�ɻ��׺�M��9Վ&6t�\�1!J�8�T�O�&ơ23�{u��b��V��3_Ù��v�33˴d1����l�.�4(���gX�gb��}@=lx��x�s01g:�sϬ�Q����x{ނbY�7�	�D=[X1�En�v
�*�r ��f>�ׇ�;��q:����(>�3��� ��,�@d
- ok轞u��k[�HL����1s����z� ;�\;�w��#MM�ί��0����&�di1AaH��*�[�V��]Uj�Gk]�|���>���f:�n�(�EG40���wn����#_��l�Q��5��=�UP�!����~�^@Ot�peM^:�z�l֍�'GlCt�cb ]�wn�Ӿ<LJAB�%nu�X�1Ѧ%�f|�|4 2����ݾ�Vd�{�		����(^��R� ��q9�C3g;d���s5@C��d1�u��p�����*�1J�r�(�(�OOcǦ��34�3՝�C�E�㈔�&��($�NI#�D_�OL�Q�>#�C�ۯ{�a�Ά�Qf�fd�@31��� ༄D�q�v����u�n����[Mo�fi�'/ ��vBTh�b{uwn�����h����  ��۝d�F�X�,��̭͇��M�+YDV�9�Tc��zժ��݁�6A�C������K�h�.仑�[�q�ڊKS&ŷ$�׬Z�-+n�K��q��6��):c�U0���Y���Fqыb���j���V>��T���b��#!��䫻�U
=#�{�{�u���$��@�л�0�c�}�;e��lyo�� ����؊&�f:˻��`�/e$�-�l��R�憘j�Y#�!n	�*���7�fc��wg��*�'`�	Ҽ'{��3M��^����</P��y	��ݯg�	����fH���u���5�՘�:7�FC(�6s1��4-�u:wm�mo�VCs���2�����nm�ބ2��32V�w��M#���!��׽�0�}����A��wn�޿��S��L��1�׫�抹��=S���z�U�����P8����q�u��	���Y�8�L&Td͢�"6��$���]������]�p��ofH���fN���Mf ����Ҏ���vл�4oo�ɋ����<�����[C2
�36�~�\M�����3{�{ނ��WG������[fQYe�n�fsF�1$� ��&[��w�u���}�q��q:�fAMf!����7��-�5�!w��fc��fL��k1	����VjC�Xr"$��u�����}���w_�����?   �ֳvb0XL2�����.avGf��,&R�<�ڭ���e�-���C�s�G2�9�VzٮDw��7����5݀����C,`gZ,�Tpf�g���2��9��G�uY��d�$��d1��N��:�aC�n�{]�d)E5Vk[B��]۩����KH�f1�𺙎�ӱz1���}wr���f!�xx؉Ӊ:�]̂�Y�w1��UxP�^�PȐ-�H8T%B����f�����ߣ��熳1���H�0�b��@P�@��!����!�w>Qws��ƈ�z��]���ِ��i���5��f:�m^!J!5Vkh]۫�b����|X�o�:�젮��:		18_��Q&�Zf��7������P�xּ=�z"��z�J�Y�;Ñ��.7Wv�pd��S��k������z������t$���S��LUTQYd�D�G�!��X̨C�tC��}�O�`A1��C��bK�]�[2&2,�<�`�c!�X�IDM��e`%�b#�&p����"�"�(�G��Z��h@�% �����7�!��=�u�[�?#P8�Vk[B��]���A��G㘆��8s1�#4�� ��/�e�,5��b�K5�M�P#Q1p(��"�@͎{ޕ9v%x�b�1�m(Ǝfd�#�:�f�Û�&B���^�Xk[���3����4�g2~�ç;���ߺ?Vd��	$E߼z,E:��]�]Y��>��O����R���		�20�uwn�j�x�c����0��vF7�1��frs�HɄt�5�:��Xi��ԅȌ��Y��.�a����e�]� ����G�yo����"�*D���I���oH0 ͝u��7[^#����\���>��i8k��:�^�ei���]a�K�b�|j��WK��]���I�ͪ.��r��3�\���}���͙,�2֒a�ޒt����P��m^�"����A|���e�b70)�L�%��F���n�vĝ{���e#^���{�u|U.��R�:�u��՚�C�]�1���~���C3kWx�1Z�5����	�~�g��Oy���V��3j�K6[)6��s]����~ټ��v]Y�٫"3B��g�~�\�u�^��j�5�fCQ��>��t��.�u��&B�R�,�u�<*�}�HG?}�F�+H�����{�uf�
}*��Zٌs�c��r-n��H����$�CPC��.����A�u��d���]5��32V���a��Y�f}���vM�tz00�@AP(�=�ۭoloG�0@�&���۫�uf�;�ؐ��"ln����O��Y�o#m��c�Yl<N��71q�
�F��cj7Y���᫿1���/�Y��!�x�Cc�,�*�n�����ei�@�{��~���J�`�:��J#�����:����@�K~\��`b0���u�,�.�ַҸ�(�&BD*4�K�M��=N�IF�z��a�O�c3wY�k9�2a��&����Y�٫"3B��o�uf��g�j#mF���p苴>���|���RMV�y����O���y��&(*b�h����;��w72T���\ـ n�m�/ZmZY$�.����n
�9�m�K��{-�v�DPN5��>o�?&�R=5�ۭ�%���1۶���=20�gj��l��]���F���3�H>�mB�|P0��aU��,ey�Qg}�>|�����~�ι�_{Ϥa�fh� �Qhe��UD_m�p�b�dd��JUݺ᫴.�ֵ�ڈ��qj����Vf1�3�s�$d�5����Wv�i�.�D��LZ�[*8��\�׫�O ��4#.Df�f:�9w+��$��!��2�Q�f?��B� 5ǌ^q�P�C�����R�C��Z��u}�,~}�I���� �!��׽�%�Kf��%�C3a�(
����*��d�/����[VЩ�ᆚ��M�$�� S�M��fd���C3k]�R�Z�9B���:P�Ӭ�w� .>uA!��V��d�;������U���EFcpc΋������P��B9v�f �s��Ҏ��T(��B<��$�
��l��'d79u��%N*��{��PSZzfB�=�NI;(���n�BI�컉6V��>K�-~��hPZ֏w�	?}��&��[e@�:$�fkD���y�T*�8B$�(�^�d���{����Ϝ�*�,��e~��U�UuT}�I:����$�D�U
K��s2Bv�3P�� t����]p�C˥3��h���S�H#i2�:$�(���5�NfN�UZG�aD���`��	�D��I�xT)���	'�O���֕���"m��I߽�h�l��*�	I��1"���2��D�� K�O
$�d��
����$���"M���ى4O9�	>��$�(���3y'�j�s��{�w��{���)�A0!�R�CBHWI)P0��>K����$@HJ����'l���1�,32�"!�����J�t��C�z���0m�)�Ė�����{�e������� m�	m            ۫k�fv��v�i�]��aLp�n�{.�q�
P���(e)r�-.-�ݞι�`��[�Vm�m��A=���y�#�ɚ9�m����n5�t�� J�������cL
X®T�������x�(uu���k,la�n��X��{
3�7K����$`nx�;�h�*���x�e� ��Rٗj�T6g]�6j�T2ܱŔL^��,T��#N;	�dث��F�Ot�LpN�
�snP���cWD^-إ;"��.5�q��<��[�"k�GhE�5jXi�VɌ4i,�e���knǎ� ��Y���`3ă>V��2������-���+;������@L���e�b��n1&�iq���/*n��\��9��@�(8eA��U���A7-����g!�ɲ֭m���Y(��H0r^ɉ4nq{\�Vㅻe�����2���-��Ж�tn ��h�M�&�_?���}��8��ܺЭg�Ӝy�2�����fVn����{�XC�����x��DD�@(��'���<*�y>|N��y-�=�||  �ͽ��&��*s9T۩7V���f�Ձ�f�4[�[�����93Ԣ�c.�CT{�u�X�8�Ƀ�u��7�rۆ������/��K6qV�5�a�ᧄ��z��g�[���3�j���'M�Tъ�����<�f�? ��섞�N� p�L���`�9�NfHI6t�'
$�d�( �;�7��$�)vQ'3$$��։:����d�tNP��u�HI��	� K
%����fHL:$�d����N@>����o�&�ص���8�sfi�X̿gw���+v�_G��2BI�D��s2sH���<FB���k��W�>����GC��fv�e_}�	>�d$�w븓eiq|Q'���{λ�u�[��F���>��/��F��>4�p8]�2�`�u�C���NfJ�A�Z�4jAA�u�q#�(�P8����� ���y�{�3�"�3U��5�31�-`'Z�`�����{�эj�`�[U�U*�������4��FH�jh{��]�Xk3Y�uڊ$��Ν���O�y���￟�ō���l�gC+T�s�Tș�Ȫ$�I�V�+�[����]��4v���j�����j��
������CC/w���ݺ��P8�]��<�.�px"�
G�>�]���<�E��3@|jkl]��hz����Z s
�i۵\��Z��sǞn��b܇�ִ#.Da��1����Vt)��$RH��ݿUP� F/x���m�j(��:�U�=@P���{ν�~����������31��b�:��*��x{κ�U��~U
~+ͷ�  :�ӲN]u؛^�`���DY���P��h�0�C ���g�e�,��h.���ȴ��h�z�Y�x�1Fc�<��U�p��8�K(q6�.&�J؇I�w~����<������)�\B��jB2�ΏUT��zʎǽ�\�p��� ���[��0��׼�*����31���"o�;�`��68pַ�tof �L6[%��U@�c�:�VFy�xL�6����Y@ {j��f1�2�Q� b/]����t�u�KnR�@tQ��fg�PC��w���ein�/��.��h>�>�܂�t���P!��}=�X��U���a��Zg32Uڬ5�ǀ�]�0���X놳1������/��SG���m�2�c��*���p�tX1���|��ϟ�3�{�eȌ5�� �v�וx��TC�ym)��x�~��߀�: �@��1� ��IE$>�k3���^��{����ein�5�m��u/?6���b3FU,)K6��5�@�I� ��p%��ݱ����]Y��a�8Y�B�߀�E����fyb���1V�H�l]ۭo��"*���	��wl~LP�!�k
"0�e��P}\��{ʼG���6ڌ �1�l�uvwZ$�_"�č�431�Ua�31��W�(��1g��vػ��3���f6V��Ʒ���}���ç��
"8s1��vVb
1x�O��f-�uު�Wv���7$2�  ����s%�i��8�7�\ ���#`���x;]�n�ƍ��2�٭4`��&�\�wI��3p�X����8����&)Uk������
����#ܓ��ɯ���dn�ڢݎK�痩��|����9�\5��М�u�7ӂ2����( F����y׼�GZ� P9��1�s��"�>^Փ��4.��:�� ?{�G֕��F(�ثf�1�wn���������ܳm%�cj�K�#��� �~�Í����s|b{ή��"��a{L�g_��B�Uo3n��]<#����Y�Cu�������F��R�B(N���Y�ƨP{�s�nzE�]�^��
��[0y�g��l��
QQ�R&�e�:�@uv:N��%p�'}�c\��Vi\���4.��Dv¬"��įQ%u�U���UB�Bk3~��+�޵�kF���zֵ�& ��)H�*����B1l����1�*�$_C��Q��a�;��$���K0�f�R&(�`��%K�h�"�"d��$���	�I��ւ� ��3�1�5a��,r0�p4�=�!����|)@�iI�t�������������l���a��aڧ.p�e��ى�O;\NFG:��Ƕ]�+g�R�[��[n��,�御 ̈́�9��,���Pe��{�_r�� ����^9G9�y����WS���AT��G7�=�1��؄f�M��]���T+����^4�
��
DCPC1'�M��9��Lb0/8�oOc32Vb�<*�#3�/�D�R�:�d\�/V� F$-�46���36�1	/p(�P�F
#����;�=����)7�9�wً�cm��̶��UY��c؉ݴ��\:57<�Uv�*�e�uR�kF(��z�������]۫���q�V���UP�o�{�u��#4�aDj�����T 9��k�0=�#Qhfc��U��*��b]∙q:�C�  xk����+�O��B�g���� ��v[f�5�%Dm����q�q��,[���]�W����˫=m���6m&͉��Q�)pZ2sv)�n�=p6��;vz��m�.�Z�������2GŜ�L�gF�tn�.eX p����wI$����E.�2��ַ�;�|��kY�q)	5��6O:�f*���Px�o<Lf6�:�1�z��Yx�i+�IE������1��u{���q����x
���{�b�6ic�2'R�m�q��4�%�D&tU�3���Zw߸�{ΩY��J�&`|F�:��պB�U?B�C1W�#��D��c&@����dr� 9���+��FB�3B����f1�T(RX����G��6s1�;r����a30$	)�A$M��+v��X<��5lLi�\�B��s��� ��Y��Q%�q-�Y�b�o*���?_��$���x���w_���~��yF���a�GhQ����:]f!�����S\=���Z�گ�~��K��Q\���7�kG�i�$�k(޴c&A���f�3�r�J��FB�3C��
 �u��:�_���"1Ę�x��c����א�M,ֱ�m)�
��W��:�|@U@����׾1D�2:��8ff���[����v`&"XGH��&6�Ġ�#"F�E�?��q�����o�~��������[�I6\@��{�󮥡㇠3d831�8��w�뺻0A �A�.�p��ػ�Z�yh�Tj���ݓv����ꪃ,����$�I$�����^|���-��
�l=K�[���u�.��y����݇���*���[L��U6�kW�8�v��@���=�-۵:#��ݞ9l*e��R�S��Ƿ��/�ẅ&�V���]�i�[���luPsn�����7�:ˎ�Ӿ�ь�SB�n�:��]��͕�ch�#ա�W���}�1�y�o�|f�*-׍o[c3]��C8��e��fc�f*�I�Z���!n&̊�R��ʰ[p��Y���|�uު�Wv�w� bA�Fb��1f��ǽ�Z������55�.��5����b�P8����sa�}գ��4.��uU��lo��z&7h7�c�Cg��T΃-��K�!Q���Y�_�Y��f:���|\h����7Ǉ�γd^��l��]��(�U$�"|�<��W����=�u�n�����W�$�*�ު�&��v}��xw�#p�[��Bp�7b�5�n4m�Ą���Y�Z��o(P#1�9�$�5��o|�sB=C@ ��y�m)��y�=��
x���j�]�*"Q��b�5��|Р*�TwޛDz�����OOu�k|���\�cxv�|��8p8,�����LW"j�b;�����\�fq�o���Pu���8��2�9C3 ��V��ʠ 5{�	4��gd&�1��:���&3h~�@ pַ���y�@P ��oYȌq&� fc����q�~�����׵����<�����{7��ﾧ���;���0�[Dc���T%/$}M���N� �L�+B��m�&�!��8�H�&��"Pd���QQ6�DA	I0��0��&��0 ��	�0 j�W�&!!)�� LN�Bf&�!�:�i��!�x�i1�i��mt�3-���o}�  m� -�           *���o�8��'��s[3��U�j#vsJOIu;�<��Q.V�B^�KL$��f���*M��9J�&�sD9uV@����AmS�q̂vK������Pۨ�Km� m��v�2۴`�n`R]X# 1hn��v�:&f��Ƥ�2�J!�۫�T*�@�ۈy��@Yn��Y�'�]B��[J���&<�$ �dZf�v�2�Xњmԡ���c6ulU��<�$q]����r
g6R^©��H�:��@[cl�[v�hԝ��Ŷ��'GM6͍��`�i���֚ݭ��h�ܮ�xB�]�H�ݣ�N�l�n�έ��X��4Ξ�ծ;B�ϖ�A��=<�Z���[R)+���X9��W9ݸ2#h��M���8Rn9�dn��A�T��U�VVA8��4cT��I��U��-�W+I�Э��Z:ɴ�@!�Q��v�XN ��Ы'aΘ�,��f䪸�{�لC�/�,Aa خ���J"�OKD�����_���w��'}O�  }�OS��SF-�Сpق��kc����v�c����f�:�U�הXЮ�̌���p!@��Co\��X;�SBc[���'<����r�i&��Y�4���%�O�᪒7���vWBlD,M�����d��Q9M����g���:����B��
 !�y����4c�yVȲnػ�� g9�R�ch����do[l���w�gL8�0�1��hݡ�*����<E�f:�UY��9em S���H�@78�ٖ�6�4g*�Ajh�$�Ԭ�0���b��M�LeBL�Y���9:�f�o1���y��F8���1�u�b�4��h�ca)�wn��0��tY��ŝ-�
ꚕ����1���_�t����I ���H�ս�z��5 M�r��ϳ�1�ч�\��:�A�/q��J3Wv�@�d���w&�j-�n���C`*�.&�P��<��A�>zd��[5wa��T(������x�ʀ�>5���u��Щ�ِ�#A�'��2�0�vۦ	�����Qġ0�f1���US8G��3�F3Jho�����Y���^�j=J�
�x|}�1�y׵��XJ��_޶�f1�Р?S�����I҈�>�c�㫵Vp��;gF�Fʍ9l/d��֣6�f��O�~�=�۬8�ӆ�w�A QJ�U����;�O�iw��DT{tMMm���{ҽ�!��Jk���]���� �o]E�L�`�c��
����z%*�>�|_�Iz�(� 	y�������k b�5nN�ۖ��i��������c�;"��}'Ƿg|5�n[XR����=e�On�W��"s
���n8��ٲ���q��[S�rs����\��caӷ.��:�1Q���r�9N����V�}��P�3f��`J���x�7�=�:�Xa��S"f1�񎊣��w&�j-�uު�2�f��F$
)Y��j�l]�:�v�a&C*ҍ��E�����Q�+��s�>|��������mCY�� yޱg�4����ciMx�c��}��2�sXƴ�N������f1�̕�����in�l��y�'���B����qdYs��^y�k4BgEY�v`��i�1���ګ5˖�1��33$ .��#3���HR�j�A�Be	T;�� vjz��H�/��	@��ؠp���f:�!��+�8�0�ݱ�
��W��G�]5���	�bi$Qغڤ!G�d3)��:�G�Q�Q��:�U��Y��u��jB�Q�b�J�f1��WP�?_�	BJ�[��nkpwﾕ�A��{0b#�� /{�_m׼��>���:�M^oA��C3w���n펊�6�7
-&��K��Չ��v�O~@#�C�h����9���}�q��3U��7�33%w��*���&8�0���o�u�*�J��Q5Jh]ۮuU��@Pk35�^�&���[������믫^�&� 2G$�I$�I����RI��kv�m$:@�+��H���R�e䵤�q�VV�s5��4��s�1��\��re����ݍ����#!�5�
��n� g�HV:�{Q;�3�������XHx�Tk������/�$Ѝ������\� �?��UTE�!�|0b5��s|u��Xk�07�c���uެ(�#�����R�l�.틻u�7}k�$�3Uv�P�`�c�!�:�AB��R��݇.������4F`z�wlo�u}\"�;��D�m)�wo�(mO,��y�{�ǩ��T����K>��#����f=�3��+Kc���ǽ��1E�����ݱ���^�N����te�72�k�]��d$
")��તނz
[���5n��ؑ�"*Uڄl�ݺ����嫑%��57�u��NI'��{������}��}���NHPQU�e%O�������Bc�L[V����f`�bX�1 Y��֎���T$�)@�!�I�� XF1��8�$��N��������d�Ŭ�C!f�47-�-��7��� Pʢq ���Uǁ�h�"�����f8��s�k|~#3��@����(����31�:��=#1��_����۬o�2�@]e����܅�
MG^��{ª�V���^���ԣ%ila���u��'Y�B/o`�F��o�'1V뱏h��Z(���ݿ��}������MUTDL�LM1W�"n��l_|��3�W��ǆ�1�����s����	nZ���q[!��t���H��5V@��ѻ�W����r3$I�5��k|u�UY��ډ��SB��g�V�F����-"8#Ԅf!�f5���;������� > �;�u�d���C ��AC��������� nt�NG^K������I|��[�'��Kt�oC��s��ᆔ�P�h�Z��j��cE�pM��|�\hM�����s�J'5͒��GFT��3��03��Zw%���{���k��Z�a�1�	K66z]�r����]���1������헶Lj-�uޡ-wl��"f��1���v�w�u�������u�����$��3��e��V�mC�i�Ј4j!nb��
�)�dh��3!Ŵ.��:��_mԵ�-Aj:�_��
����� =�>#^����~��d�-׍o[���/{γdo{��Dk3����U���L�-�uު�W.��\!wʲڴ�lR���k2���&`1J�٫��B��{ސ�g�c������
(�v���׼ֱn3$I�j����8j��L�i�7�q$���y��#U�xv��j�Q�b��ݱw�_
(����i����.Lv���[�֜�8�_��Q���^5�m����Y�dAoq�0�c�㫴,���L�-a��Wk��fi��o�(`��>9�p����ϰoP��`Di�5�<�u<����JhYZ�໷R�.�e�"�����<\�g]����8@��5�:�B�
�l�\,���n��m�.��9��E��X��}UT����y׷��`����> o[h�c����S�/����*��`~����dv��F  uݺ�9����k!:%g^Ʒo���'ͰX!'�����C�<Wm]V��fзj��ta����C؞�0s���pK�;c�Tɣ�UxiUk��K�q�H�{�����MM'�ګ�+���Go%�m�1��~��]�.�;��GeD��c��2<'1�����0f��&��ݺ�B^��$�#�����p��8�SC1a�uU���V��^NN�[k�� p����2Bd�)PDZ���l�9��f0�k����OEn�W�1��{�u��#7��`�~#3����XF����E��uΪ�!���v#���[#�ձw�w�=���3m�Q���qn�����A�]��3��>wß=i���"^��$� ]��vвM+��Y5s37��{�7��,D�7�@}T=���&-�j��1qEC/�@�u3w�ci����F��=�:�CQcڑ��2��$�DnV�M��厛-.�����O����@����ɍE�����g���f!��+1�3��Z�`ꐦ#kB��v��~�@ 
~���fH����y�o��ʭZ��uv�	2��	��۩�wi��V�8�Qhr��B6h��%��ԅ$ܕv�f�틻uz�̸�m�=��k|c�����S#Ww�;κ���F��Oh��Z��Uda��.�v�_����9��{�kY��|M���|`"$F��*��:Q�!�#�k)s�H�v�G�3E��f���]hbY���`���}o<U@  ��            Y7iav�{o��6^K��!�1�h��=F��lZ�:�8]��!l����-���h�/;pm�m���f��6H�֍8<�i���t7=�$ʆݽ�X*�[utڂ���t�C��~'>3�G!v`�D��펔!�86*;-Xf�LXk�X�b��k]���Y^�Y��Te#�Q7���=*�ԭJ�9�`����i�m^�q%#��+"��1��j�"��bLk2��0JX�P�w���J;���EU�����(�n.��P���m;r�N�C)2�{9�֌�s�]�lF�����εqg��@+t�l"�3n�y.P���IvDۡ�� ��$�C	��j�j�v�n�����h
��:�9������n�]s����Z�-�\
� UTQ!!�JD�K�R���֩V���n��i��Mp�j+o#�U�q�O1�:$.��Y�lݬټކ�Xk2^���8"�:�e&�,��ZW�y܁��Y����.� ɮ�m����;K�1R�*�)fe�s�J�Hh#wN%���͢���K��M<w�*�	��CA�a�W�I�Oj�������P<�CO
����vm��7��F����X�\�����n�f�b�l̮zߎo�	sAƛ0�E��=U�\�c��f���R���55�.����@�9�Z�$�4s2o�t  Y��Ғ��\i)�{ι�u���bZ햤)5]����{�k�����~C����
R���.�8��pL�����P6���~5�m�����A����&���=���{���zU{�=��פ��� �|<���š����ӄB���f!����C��c3#J�uHS Mm�wn��t5��,,6^��,�����3�̍HaN.�o�".в0�3W�"�IM�uΡ��c �;�ԅ�cG1��@	B��<���:�s�L�/�> o|,{�u��"���`��ޏ]�,�!Ù�3!aFY�	d��pS�1�iZ�q�U���7������0�7v��]�!��*�~P>�����k^�J�(в�ػ�WhK��R�5� �c�_����]�UB�������|�qDdi)���\�@��/@��f�B0vI�CAmƬ1!#Q�ZGMGY�l����^���^��d0��>5����������Fm�$����Y���^���Q��-��7�f4G{�,Ֆ�о�Ԑ�DR���v��[�U�Ab�$�I$UUUZ�u4�h�·F��Rی�Yڝ�Uő^,���i�' ��y�L��K�2�&�i5!��s46�,#{ѭ��9�ˠ\��A�]3�.��S}�:�Ӧ�����'\^aȎ��i�q�+p�A�(����ub�Ư��8�p���5�:����UCV��$djևs�����؆�eGMGW}�:@N���+7���ai=���f:���z�����2��Jlkuz]�`l�$�q$�0]�����X��a�3B���t(!wla��8Fs�q��V���]�wn���J��Z@Z�v��'-���F� k1�o��wlCL�{{m��A�P(Cj'#�$]Z׬�������~~rWn���b�
8�b&����M�.�^��\1��[@[�U]U`�@UDP^KNGY�b��E0LY�}�vVe�1�X 1�f���w�b�d?�5<��ٰ2f�3)(�
�]�{b�^L��3���{����m��c��e@d
-VZ����lV�>8�q��j�o���Ő2f��L]��T�N���{���<}�����f�Ǝ�ࣉ&��z��]�v-�U �~'܊ ����q�^�*I���_��l-'�������(=��de�E�@s:�x������S�&4f�e��z�� <�W�Y��9�r G�fc����ɐ(�,���,]�����*�}��@l�jI$  ;k��ג�%Ie\���v�4���Kh���Lnt4��e�A*�B�V�F�S���D��n玽r�=�q3�W�ڸx���9!�y��u�S3VD��2MU�`Q|2��'����i���MV����$q)�Ӛ�i�M8@�xƷ�_}�paY7�"�1��Ùy*�d��ts0)N2�3�P1��u�����ZOc{c3��cDg{l`�c���A�`����Ē$ ��nF@���õG�t��TQ�>�U�p1d޺��&&R���W�T  �
�4Ƴ9+�C|̆2d
-����fAe���c�FS��1�q����n\d��wn��1dv�We,�U!�1�l� �V��HK��́)
MGW}c:�y�fc���wі��{@Z�c3]��E��0v���Ɩ���Z������9��w�|�i�#z����Ս�D�y��%v��#
ù6��SbA|Lp,0#�R1�]$!��<��٤G�D%&ńcb�����@e�^�WL��L`k$Z��ܷ�Dl A׬� �8Qv�T��K��"�D"�!��)���<�U)�G�(�/$�1u78�{
-y��r�3�x����F�)Y��
틻xO=�ߙ�e��.
���Sf`@�c1C��(�0���31��lo;�⑦!�f<;�]f[�=#��sE�R��+�n�if1�+�8�..�s�pj�(�W
�+#8Q�;��~��2�zOu�K[c3]��n�m�T�gRu�:��n�.��!�1p4�Ɉ���fu՚�cOh�ʏB�ݘn�:ѧw��@�`x ������	�)�A��>Ҿ��d�KU����s1�s-��{R6�5��5�<#2�+z��4h���)#� .��ֵ�����b�����!qD����3
�,m-�X76`n�)rE�T�A����<'�9�J���+�o&� 6�ю��2�n	�f�V���������v#���.mT�3E3�[��g4�sc��]�]a.�Z�$M5]��4���Y���F�L轏{����Y�b|�E�LWoy��Ù�iM�=�cQ��uѾ�dv�&��q&[�K�X+�˫v�bT�$D��Uݽ���n�T��2nɹ��=&�,E](�A�7G{ڬα�|�fH�@k�ƹ���lY޵n"�*=x�1�n�8k�{�ktd5f[ +�.���C��|��V���.��S,8���tvqo�|�4�zO��ol~����2����[ ������0V�m�3U���޿��I� �|>@MߛÞ����zݑ�M�v�j�2d
- -m��ce��=�D�P��-�MƢ���==<̺�U���c\㫾�d	��E�Tzv��۹XF��cX�	�B�Q�e���b��^��\m4������� @U
$ ��*�T �Lh����JR�Om�s���׾�s}>�ug��Mȫ�p�t�kmj��Fl�u'ϟ7�>[A!f:����(Pa��Ad���u�n�ɂ���������u�[�"2F�Y���u�la�fB�*=�u��Ր������!�9$ L˚�3[�[���n�]z�
0� *�Ӵa�	11b�M�݈^{<6ȶz��H�16�\���8S8� �&ŷ4�	G�jM�l��a��<�˼m���!�]��ŉ�Ws3uW� �T��2�F�D��2�u��z�'�fc���ˌ�^�������W}b|�E0LWls|uw�,׎k�1�431�;ޱ��7{��t؂(NV���V�1��u��y���
E�Z��ݫd�bFc�8�&@�гAkl{3%f[�ussu73;�� !��%� �-������>����
�>߸d.&�z��{�r�if11f�����if1����܌���a���31��_���b,�!10�E���xj�*0�����c��ΗVF�6����431�B��d3���w��˛"��g��!@&�S� dQw��Q|�7��uuv(�Vikl]�M���_"���n����Ve���Vm�bQ2�@�ĜQ��cTrx��D�Zs8���c������%��`�����u�J틻�^�r2�zOd����3]��E��Q�� y�w�u�׆�����E�lq��C3w�cy�{�_A�f������\���AFA#r8`�(R�-���ɚ� M{ι��5�E���P!�fc�λ��gb�(لp�1�����uf�toj2�)M�u��՚Wl{X��Fci�����'p��������*"�n)�aE&� ����/ִ����RDEH�g�����X}z�NzkPP���J�"�-((( >�ZUiD)r@S@b���B��y���h������� ���(����p¨�(��V�Y�/=0�ATE$�2�/�"����B2� )H"��(#�D�� ��&b
�V	5� �@P�7�$�H
,H�B�HH$��2@Q��%V�P�B�C���Մ�h����]@�����(�0(��v���ѯ١���**��U�N�fn�9��1���=�P	���*K��)k�H���*i�_�H}b��?�P��_~w�Cz(şB��T�hED ��߮?r~������H6d
(�U�d�<�����O�g�X���OO�
��������� i�H!�� �����TQ 9����_�G���2��IP����Ƕڀ"H�d����2~����cN��""|�w����=T�DA�g�q�Ĉ���� �R@�Ei!Z�X�P�X�(TJZA "E�hUiA�
�	�LTTIH�*-���C%R�

J�j�JQ
JPB�Q��TA�i@
�JB�)EiZF$) �J%���JiD� �)J�$(JJB��$JV��D)J��X�eV!�ZA�Z���!Xi$B�i��\D"� "��b Y?09�X׌K�7w���+c�����{�����B�)�8��������������xOAA�~���j����w��*(��J~�������?�_�O�l��VVFK��g�Ş��O����(��~_<~������ ~P���g���"?��|>�w���a�\��E >�ڨ� �����`?L'�3)�d�?�|�ق=�S�TT@=��0�"G�~cB(�����;�g���	ry��(")2�SkN`>�R�4���A�"� ��?��}��(� ~��}?���{(
?�����G�?�}�B���1�z����?��¿��������X����~A����Q >�"|����_�o����g���r�A���-a��rHA	PTw�a>�.���s/�<#�o��.|�
(���WI�=z &>}��gܟ�a�PD�=�Ԗ_�c�����!!QD ���i��_�|Q?��|��QD �����>߶C�fW��PX|�?���A
񮁯���"�(HUk��