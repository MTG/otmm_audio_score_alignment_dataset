BZh91AY&SY���y߀pp��b� ����ar� )@ $ �  C��*� �   Ҁ   t�
(  P�O�  zRR��E]�% %H% �TI(P ��$% DJ��Q%@	H�  P�UP�@R�    a��    �@�M }*ͯZ^�uzn-J�iW� ����oJ�j��Z�b�W� �-Je��  ��@�0�} ��LM=iW{��=o-Ҩ8��h��A]ޕ�\�][�Ҕ,�ӋWa�  <    	 (f���B��Z�|׍к���������� ���������y�=y�.�5˺V��M�W����ywo ���*�����}_mqof�,�5Ũ�siW�}�Pϩ��ϼ�_}ܽ�^/u�����m�7��
�     �JY�v�����ھ}�������[�R��uOW7_^��z��o6�^O.z��� ��m..�oe�� ^�˔��y5q�P ����wץ���s�{�|��۴��P�k�.Yr�v���Ǳ��x���  �>�H � PP>�M��W������;��Ÿ�� (w�^���l�,�m+�ͩKJ���\[�gO,� &��R,�r��|
���nn�-�Ú�j_o^����w� ���͹i�ξ���ݷ��^�w� ��   z@((�`���-x�[..�5�wm����՞�� �{}����qg&�Ӌ������������aū� }w�t�.�'9_y@O��f��[��z���W���ҭ�����*���iqiͯy�;�w�S�          4��iU* 4  ��)��M�J�   C@�z�RJ ���   "{J��ER h�  @ 5?B���*��0�  `B��*B	�D�=Sz�C�F�?Q�zjz��"~?������W����ۇ���:��u��  CW�@ @(  �DP  ��  Ā��  _��@ W�%�  7����  �������Z�s�_�m��f�aQEA�30��4�Fc��X[����;�w�Ha�"�6��G����͌HKS�F�ӳsI�dRvf	�cI���z2��4DF�i�,uHl�c3��ί��8�7A�X��h���GI�z�33Gp�z|�	BP�:���}��' �ʓ( �bA��h�I�h<�j�-2kPtA�3gF3p7�\3��%�(x`AIAI�gn'V������N��E��(7��Pa��k1��I�a�PV1��	BP��L�����2��#�ζx��k�ַ�<���0�f�l�\8c�|����^;�ć�&��p�o�!>��qTtڋj<3{�^6p�;�qѳ��x��d�5�c���i���{��s�D��k4w�9����.}����j7*z
ڕ��pZ9���]��YF��vs ��Z:�Aw�dl2=�;��2�3�	##�X�"�=N�# �դ����G�m�;�����Ù���C�:H�:�(�b�|���F�6�Z��ӳ]�tj��2C22�������25ݽfF������q��w��� q;L��g�f�q��w�ܺ�#0��"�xQ���T	Xa�e��Bw	F�a�JRg��g^������9�s]����4����:�M3�yf�3vt�)��[K:�xl �N$Y��uhJhhI��df�[��-�	C�PA�u�4В�BP��L��X�Ѩu����Ү0�������{�5�#�B�%�v|$!9�A5!�Ȇr�A[��d��8I��5Y���QU�随::ά7�£[�r5�<�pXs���u������,��0+:;�.����:���=��<hJ^�����0���ֽ�N�\9��]lxzw����A��0���s<�!<�'iG�����}��#��\�Z��k7��|�)�N<��^�y�\̭� �N���p#��=��z�=Nk�6���wĔ%��k�;��������a�3�u��MS�dbQ���C�2��E��d�9�3g�m��h۸��=�A�2c�����F��2��y��kXa����4\�L�klXY��]��d�&����
�4�\/���9����:և�4ؙ[cZ;�YìCu�۬u�h�fo��Z�U�w�UKHT+őG�a�aք���X�k"���0tdɐ�d5��u	G&:ѧ^���2����D��\��wC�J��i�Y��4��h��a�7�9�����Z���Q���j���Z�#�F�p�I��.������x�4f��r��=̷��K�L�"���JH����Df���[�����δ��:�!��0���RVG�f'�����L�-;<;qr1#Z�&�k^kW��5:����T��(J<)2��J��ݕ��(����;��ݤ׽��n�<9FC�dɖ<Z: �V&�����][*�5�]lI�Y�N�����Q��˘n4�fwj�E���2c ĳ��Yj��)	b��7(=6�Ӽ�;���%2EO	ʢ쀳Id;0��'��F�s1-�5���ސ���ݡ�����8.�B����j(,�f30ۆl	��ζ�ގ�����3��:��#d�Q�0��X-�G~1�p�d���n��1�Ն�&����a�x4�6���f	Yj%��>��V����SևV��5��a�ɛ#����~fxk�9�u�6g�鉢V�\V�w��7���4Ր�/>,���L��sA�0zu�0��e�kiIa�#�|������F]h�hֳF3Ứ�Ն�����Xj��n;�6s �֭�rِ�=�wK�q�8�K���8�1k[s[�Ֆ�P�eFi�ZN�4:�	�Fa�Da�3En�v�"�D�����u��gg������;��97�kD���еaEt"
	A�Q��ܺ[\�AmM�'3"��h�V���ٷn��ˋq��7O��)�(B/�+U1|�b��q?�Z�I��]߈����.������]���)�������u�=Ra]�xe%h�fF�Z�Z�h�C}VV����C"�4	��H7���'��s[�[.��z�g:�C�~�����)��&-�UlQ]�/`���V'Z�缻�Xu�juh#Z�]ֹ�gC�v�GIj��;���C�f@d�с�#&�)��Grd`XNd��y�ǹ�M���vhcR��Rc��9�i�0e�	���V�o�Xi�[��L9�98Y�<�v������sFХ���f	�0	�F��9�%��(dѽ�KZ�JF����td:���ّn4m1Ց����U���i�	z Ǚ���MC��CYɑ�.�WG{뮎�u�:��`�X%
.���Vp��Ga��Y���#x�D���{�/�����''���0.o�9���O<7	����R,Q�S��Q^�_/������g� 0�v�!)�l3bRa�w˭�n�'�k��λ�֣IFY�:w`�n5Ga�J��J��i�o����D�.k�p�3y���f��6��21�f�:mu�q�jN�.�[�[̠�5�t��g:}q�u]����Xe��Z��ѐ	�p�(������޼oq�ʴp�ݴ��WF��:#��49�N����Opah��*�if0F`�,�t���oX^����^s� ��j#���z�F:���ԛ
���0�q;�O9���{�!��vl��ך�"c 4f	�z��2���jz�21l�����=wu�˩q����rs�&�5��g��{�2pJ���ްi�v��u�����@fĳ6�[�Q�ގ:��%Y��e������F�����>�(_��%	�&A��!�bbw	Bj��7	BPp抱�-f�aя#1�J�x�������Rj0�4�U�4%�2�$�α#��" �g6O�`��@�Q�0!��rq%�#�0)�w�Oa�!3��gRdrM\���pf���z�[�x��پ�u`{�J��K���d�NX���O5��G{��m#Z�Ѷ'�p�W���fF��@�Y�|�n�	U	_4���d��:�S�b��F���7�.�G�9�y�p�d=�C�f.��v똆bzj5���jms�������Dm�Ӕz�K�z���:�:��$�r15[ۋ�`�I���!��j��#4�;�~d8㳑�+,M$`fPP�%$裝�3w9M&ykv��jS��y�0rMBR�()t��vM�E�;:�i��%����s�WF`K���FC�<�C׸���(�=:��v�n �a��9drgRl,1�ٳvv��d%	BPf`q5K��\��!�4vZ�3,%�:!��5i��X��u��n�K�bj�ٓ��2''E�����015�vp�%	BR�bn�YA�Plr!(J#3Ak0ք�l�(֧F���r�"r�.BRl�:�9�n7�à�`�Ի�ݜ�=�o��:�k����\w�dr4I���P�d$C��`�%	I�f&&BXњ�:7n#4Ն���4U�1*�ѽ��sd6X�v�A�m2�a>0d�,�!-�Ɲg�d��b2�\ؕ�XK�����f�V����TVX�I���GF���g[�͆����d8BR�A��i�f�4h2�Z�Z�M�2�#r�]n�p��	F�����r�i����9�r-�PkJ#5����r� �X��]	i}s�,8ttts��z:���T�.��+�\��l��w���U�Z6�*�	��o�a���k�ݛ�p�gq��gZ݆�3V"um���qm��/w�"w�V��5tKݎ-���;::M����9	X�'���^�s��1��*r���c�y��f��{ui�V��O�����zRga���ty׽�k]����u�124HfY����{��:�P`�c��p�[���bd%u��BVh�O�f�F��J��)3��Äd�s[b5��ש�49��Mk�dظn{HI�TN�i�R���H{�={�k:'V�&�F�t:��j3,CW�w��tl���}Br!7	�%)�s|<�Ox��������uy|բB�B�T#��^w�x��|w��0݁&g[����o������rL��Z�V#zN���y`p��9�Q���B�)xu�L5�<z���3����=4r��,u��f�A��[58�&Zu�f�Xh�&�)13N�y���}oA�wxa�tF��rLo78᫂d%	�%	BP�%	BR�&BP�	BP�	BP��	�J��J��!)M�P�%��NUtk�����X�Z�(u9	�&Bf��%��tl�F��Zuׁ�O3#�$\���ʊHh�8�8o�E7Y��X��4œ�����;g�̌B�{�٨4�c��9�����$WTF��f&����Z��fAQ$C�涛q�2V���ZF���{T_lA�ؾWi�ժ^|����NYWy	q�2�݆�37�E�:�\�0˕El(MGc�plr<BP���ߗ�3�^�&v�<x�c��Һ#Mk}�u������R�s
��Ǖs����Z�J>
J����jK$�5�v���$��Mo{�y�Ѯ�����a���cgHEQbi��w����>��(E��f����a��3|��u��6��&{ֺ�:'E8sY�������?�9�n�������    �̀ � ��@���� h        ^�   �$  ��        � [B� 86�v� �p �@
P`8 � 2 R���� )@C^���              (�� tQ�(     �@               �           �   j�m�N�   p		8�t�n�u��0n��2�UV5Av�h-�  �m���=-��ہ�ͤ�UUT�*�+�/� ��E��w�ƻ�۳l  @�m���岉�T��52��Y��:����Xd:�����l<��W&F����V�F�"��Y��`�$ �� �[pN����m�m�85m��R�m�[pp$lp�lJ&�)�u�崐1�.���l I�l��s���vN8-�N�a�� ����N��ybZ�V�M�+-U;g m�uSWN�͎ ��@��x{⯪WN®$�5�`n���,ga�v[���V���I.����kn�����nպ*�-�8ݶ -� Z�6��[@�kl�m��� 6�M*�BMR�K(^����Hi  ��檀U�ڪ�`C�*���kn����H�����ٶ�ͫjY(6֬�����K�u*����E�� Ve�3�ٕ��f�S;
���AP�f�[ Cwa�U��[,�7
�.̯�sm��J�mV����ɺ8�qt��uUA�7P �v���h�ݤ�ܒf�ݮ  �m�&�`�D�t�o��6���m�j�Ux�%�vj��l[���cͫ�5�Žl��$�  �      �S��2���*�ps��j�%d��m��-��Z��{m��*��u��������Y0�l����� 6����I\v�m��6�[Vq�Qeub�8m[6:�1-6݀�\�#\	2Yf�g���T˳��TSh\[wl�F��3��(6q���cr�Ɠ�k�]Aԫ�,R�u��:n�
����T���g ��]���HHu]�jva�P�Z7&��@m�k�U�m�@�k��]&�d�r��n4P�B�Tp�
��We�_#Pqk5H��$�� [S��zVV���?_|��V��LX���cr�J[�2%��$A�i���؎2��r��		kn6�6�։-�wl6�� ���"@   m-֏5Z����8lTe��I�UU���e�*���m��*�cK&�@X� UU�vYj�er��#�˻uR�V�\�U�iN`:���S�p�R�v�v��m!1��D��EUWF���(�=uQ���=�� Y�v�ۛ�������V�0 ��pq׭5�l��I��m�Z�6���cD��`Hm�5�Sni6j�`m�Zn�%��mp:m�mm$5��m(m�>���m��oa&���U�kv� ��A�V<�����pm�T�5F|/*UG����b@/Y(Im�Tʼ��UQ/] r� ��^V��R�^���p<[�ڦU];RBNr��eyz�t�[\ۨY{2�o0 �ɴ�8]xx4]�@b�;�=Ƶ篾�6�/'��Z���ܐU,i�r8�$��*��պ�o�	-��E��i|%��a!!�i�p�
l�J�TpmT�P�F�Yv�&�8��h���,2@[@�U�ku�m�b� a�m��hn�N��m��IN���Z��M�����l݌��-iV����3�mm�z���[d�$d��[ d  ^VV���@�*��s�P6ͳ�m������ 	$��m��t�ִ -��i1�͜���H��@ m���V���j��W{�$�T��k ,ho�y+J��@  'B��v�q��\��8nݛ� �m�	��u�N���^����m��,����*s��Ýit��=Kx�j��]����Z�:��cmJ�kjQؠ{�1Z�܂��7K��qq���e^rT��l�܌c�-�n�΢��IÚ�{*��k -H��i� ̰�6����iU�k�^��s�PV�Ty�t��ƻnY%��}�k��iV���YUZ�i,�J�5J� *���7RT�� p['9��ڤ�ۭ6�[ul8 2� ����͎��q����v�L�N��(�]A�*�UT���T\ Bt�[ �`�m"�I m&śi� �Z������2�e�̭R���e�}�Z&�jt,�k������e�  $nܫv�WE��m�`H [Rm���y�^�l��oNI�۫I��RZ�O*�m*��.Y��j�T�z�|��:T�#���Ip2MltX�ﾕ�u�jyP݉s�I�L�T���e����]+E�Q�^oX1��	U )oWm����s(�]ny���nڎ*F���#�m����E�f��NwaUVw"���/(�6�e�7Q�:S��#�%�����USӉ����*����N[J�ս�� ��d�	��-����&HY���[K{M�*� �Pe햛Ul������x)\��m��j#uJ�:K�����uj�ګmۜ��4Ji�t���Ͷ��}��6�z���JS]m��y5u�B�Ȱ۶��-�m� ض
]�
�mM+�F��kn8m�j�h   Wm�Ē	 m� ����vW�sl@UJ�콲j`u�l��[�	-����N�lm�oT-�� gYV�$p &�l�`m�r,l�%�۫�m�� �%U*��m���V��olUR�MTK*�����8mp��W�j�嬊t�m!rj�V
� 0�us�d�2U�y%� *��n��h��k�76������c�I@��Y�	�T�ҭU�\l0l��@ +��̓�v��3&�  �m��L�v��uUJ�4�n�6��v��)2���*�@mu$Q������)nwnݘ+��m*��Zt��6,+@[S�a휡�-��5����\�N�˻&I�Ȇ6��������������  -�i3m�[]m�p,��i66��z �`�@jBiV�
�%[h6�6���6��gs@4�U:-���-6 ZI�6�"@� 8m��m�l��:���[A��� ݶ�ම[��n�l�kh�i ��XV�2��6�-=ޖ�w��` �  �   m8pqm��	��Y5�mm�H�@�����8�Zll��L�B�|��}O�f���`��� �k��@�`h�� -�m����r�-�� [�՚��u���4Y  Xa5!UJ���D�K��M�*�J��ɫ��r[tu��t����!RFka誮�(�X.� :��-W@E����ͫm"m��m�tS�8N��n�$�]�� ���j�[��ҁ�-������z�� -�avÅ� �[[v�	-��m9��p-�l�ۤ�t�   ��f� 6ٶ�ր [@x �
��T8i&UVX:��� �i���m� �sls�lVI�q�ӤsE�#j� �m���PYV%i	U�j�iV��WP:�[�m�  -�v��6�� km��8 � �X`!�Hl�\�[@ �`-����h  �mm 	�e��׶�!�`-�m�q�lC�׾���m �m�Z 2N�	 �� [@i� ��   G z�h  u�-���m[ $6Z3�ݶ�` d�M��VÀ[Cm���ms�l�؆�� l�� ��MM�8�uf�K]J��nY�`U�Խ�v�h  $� m��-���@6�mԵ&��m�-� �v�P-�ݶ���6ڪ�  *�j���%�
�` 8 m�ŵcZ$[�Sm��ނ�m�9B��:�����vk-��ڵ� c\�h�%D�\�Gu-)F���j䅆qŶt�NpUU@U�*A�}}Y. *m$�m��F�u�u)U*�*�W�[��c��`�nt�:j�X��%��-Gt��)�U�i7;
��:ܕ<��d�v�l��U6�6{F&n�}��g�O*Gi�Uglʙ�e����G6��-[����n�B���    k�m�� � 	  !���ڶ�l  .�-nm�� 3��i!��\'E�TY%�2�z��[q����m�	i�V�F��5ki7`m�H<{�#����[M�M�8X`6��H 	�� u�����V�i�n�n��8�� 6Y(l ڳl < �[4�6�X`��6�i�` �`0U@�Kl���]��3Me:[:#I,���F�9zE�إ���gnH  m���`vʹpKQUmU��5R��m4���� A��8ur�s]ȹ +j]��`*sUIֳ[���[�� � ��,D ]u����'����;?ا��?�pI��m�Dڠqv�� �� *��`a�H8��g��*�b��H�� �OZ���@��+C�h�=Έ<l�3@�*
�*�: =L�$��8"<�������a�:B@��) I%�T%6z��:M�=�U����AC�S�$^'o����b'< H��� 4&���N�_zN���'��(�*����Q3��8*�P:�IK)��	�z�>#� :C�'��p�`I��A��T�H$D0;v��GHt�oH��҉��iA�;R��@����B4 C���W�@v�:���.&�G��@�8"���G�C�!��C��B���zDa��#��M�� ���8�=�
� &�FP= �d�
(��&&݉ةҁڞ
,
K v!��@����V@�}��Q��
`Y@e�)Ъ��N�����,`��ĸ)���,�9��!�`]��ઇKǽ#���lN6�B�N�b ��z�DS����  ��k3��(���_�hj��А!@�-EJ@@P�)^h�BV
UBR��!�K �B2& ( �)�?�kY��zݳ{�5��{�m[D� E�r� 2 R�k�6� p���      �[Uv��7I��\�� ��JZ�2��60�&.']�&��+f�V�����FBٌ�Bا��3���Ѯݺ���
s�����T�@�6�\[��k"�j�v�4h)��I*��/!��X,����ϻ@�U�&�ez݀����*�3J�UJƑ6i��哲��;�Q��u�C<uyB�V�}���ƹj�6���q�5���3F��6�x�Jss�I;a�d��+FVqn��i�ON��Ic�SM��aGh������6�]��j��ʜR�ڸm����T�1�b�Mb(��,V��
˻u�E9;Y;<n�Z��u.��c ��b��x�3���e���u���*9]�:4�GB�����һ2�M���m���Kӧ\s�G��#[Y��M�v�r�4�Өy`g�U��'�h	M�-HM���N�� �6�e����� �D��̀#s��vچ�B���/A�=�ݧ.9*����e�xRCG+�lG3�!\�Ԑ]#�银v�N�
A\�"��Sb�r��K47b���� �yx�^_E<��b=]����W���j�����V잃U�]�<Y5y�6gk[rpì�[��9�Ǳ��u�#*nvl�^�l��[Oh�]���֣�f�*�M���"�Ҳ�UR�nC�E*��/���X��I<��:�eR�.6���mm�ơT8�oh!'$[;K0�u�-���@���Vm�Z�u��8&s��:l����*���g�^����lve�j�j��_@$���F��`S[&kd��R�	��|��g`�4g\i95m�3��9�<���k�60�P9�P�-��ɝ��%d�n�3���٠6q�&��`�*]�������,���5�e��u7L9W]��l�6� 	 �lg]�κ�/[ ���We�8��v��{�߾�sЫ���qA]	���� �(/J�O8��f�C�H�{���7=�����UV�s��ڌ��v�Nz�QW�6۔���N�I�n�-����wZ:�'�l�N��ґ�;s�[l�M���'&�U<,���\ېvQ]v�{l��I�lgh���;��W��{`y�9�l�0Ek-m���sF-cF��mv+���c��7\�nf5�V�VB7Jgn�p�����i�ƕ�I�9ݗ �����t��䏄\������rq��ʼ�{8�89�m��p�p����q�r���?w���w���������ù���}�R=�-��m�o ;�^}��� ��F wr� ��ߋ]�7Aڤ��{����ݾ6���`�޻�"�����-��]��Z0���y+���ԭ|D��:�mZ���`�}vߒ�R�`]h�#��ș������+ u]����qq��E����u�kma�f�se���uJ�Vj��[���]��Z0.�`w+�>�7G�"���`s�����-m�i�6���%HV:T ��;�{�}\���}� ;��v�|�z��ETR��l�Z0�����&E����F �+��n��+Q�l���;��v=�ml���`w��jG�%��:Fܶ����F��0.�`w+���O��:��y>�j�h�4Bt�;S���%�7�)�W�3�
�\(��ɧf$�B�n⨚��ͼ�˭�����v<E�Km��ZH�*�{���;�^ w��RY}�r��zDU�!H���`�v߽볚KT֍,kC������*�7�ʻ�}�)�³V���݀w�z���ml���`�v�_yx#��b���n��K# �.�hrW�� qu/��~MtFx��l�/X@o#���^^c�x�:����umϨ��׺ϫ�i�z�*��n�@歘ܕ�y+�<�����s¶1�V�Z�S`�w�S ���9���yu� ��3S�UvB���-� �����}��I���w�� ����k���r�7-��呀yu� 7�^��""D�}��k�Z]�^�la�%���i"�� ��F or���V��# D�ߟ�~6�������ZS�uv"�9͞�S.���7�S��ym��c�����q��ۗ����� <����V��# ��F������F�����v_����,�˭��x��P��n"䂮�n��,�˭��x�J���ζX��"���[֓Z�s�� =�� w��}�# J�".�FZ�j9M�s�����^�e�������|߷*�������&	�"b$C
�8�$�A#��P��kGn��^���p�p 5��Ma�̓6YY���]!j^�5��\B.�v��s�����ۂ8�1�Z9VB��H�#"�H�f��u�>�8���&&��d��n.v�lʜu��Ѯ��Мm����9)�,.��[�d���=���w7�����3�a���x觞v��`�d�9�j�,G��D�WgX-
Gd�ꌳ�b�Iu��pl3��/�7�n�B�f���먌��X9^�Ճ���q���^/l�5���m���)r�vWz �w�o�d`]hϾ�}���_���7A��r[v>���ZM�ճ =�� w��|Tr������ɢ�&��<�р�W�� �u���#:%�
JFܶ�ִ�oܝ�
y��7�h�>���.�`�>O�t`T��Kv_��������ݾ6ϻ�3Z~<�Y�)#p�������ŭN��W&&�כ��2v�[�7%�J�]a��J���}�\6���}�\ִ��Ϲ�`������U�[��7��w������z��A�"���p�BQľ�;W��?7\�z�lZIh=���i
�R������p����`]h�7�T�UN)+ �����I7��]��}p�{������{ ����ij�Аv9.� ��рG��}�֌}\� ��U��}JQE4()#�v���J������W���V����Dl����s5��Ma7f�֌}\� ;�^���`wȌ�?:����m6>�����&Asw�{�� ��F��)Q�0*QIS�װ��]��ݾ6b�֒	 {@����W���r�=���*�5���7R�	Y-�`}�}��>�o��ϧ��߽�u�^u���UE-�j�˭�%X�J��0������ӅzK��g5�չ������-�vΧۉ�M��Bth����������1W1SV`��`y+�;���<�Ѱ;���#ڒ�b%��6_���iL�;f�[0JJ��L�R��Ywu�B�%�`{�p�{�����ޛ��zl�ޖ�h�h�(;M��yu� ��� ��U��A�DG�*�齛�DgA��Х�6��?yV �W7ZNـyu� ��L����p
�*����[�Ė�Z�v�s���xGZ4��˷^G�k��&~��� �K# ��F�IV i�� #�V"�Km�﯍斓�L�z�:�2l�{�`y�^u�b�*����Y�yu� ��� ;�^ܭ�/G<+H�a]�G)���]�w�z�����_{����{�ԏjK+�vff�������рyu� <��z�kZB�_��B;�[mm�Ӯ�s�7]���e�n,������]C��-�`�it��G���W9�����Q��1�l`�����v_Ud���1�pQڜH�ݝFv���U��3�v���kJ���Ʊ��8�ۺ�M�l1�kndn�`A��![��$㛰���ƺ��(mS�P��l�F�&��ё�{n��T��<Ƃ.	�O��w����{�1���8�q�n�IV뫬v]�6e�����r]��9�Om'��g��؋%-Dt�rKo���o�`}�� ����~����H��mv������� ��F y%x�J��h؃�A:Ό�n[M�}�z�����""e'l�9�f��)Q�H(���[�:�����}|l���`{޻ ᯼�u*�]��f��}|`��h6� ��U�<�Ag�;*�-�g����U�k�څ�(j�:���\e3m��G�}��s�@��.�`�W�t�*q�}��$���9����Em�9M�}�z�Z֮��߾�çR�{��Z0�"b�v����[n9n���ޛ���>�o��}�z������t�nKf��V�˭��y+�;��L��Gmn����{���������e�﯍��ZZ��b�6���	�����561[���管�:�Z��m��P��ւP��!YG��s2�����Y�Z0G�R�,�.")*%���{�x��i&��eK�����w-��_|G�`T�W�諻��c�������p(w�����К�*�QL�6f��(������4�	Es��QfD&AUf	I�д��CAV8dSE�Y�fkcm�8��-���_(�� ���-w�@B�ܓ�@S�p��̀rJ�"�(�֢���IX$��!�L��Cu��v�����-�!� Fc�A!HT{����1Ec�;�>�M�S���=֞��@My�! :t�C!(H�;Q�� �Ц�BBID�ZsA��9C,0H^�B�@�= �Q�*t��;�18���� ����O�"���b/�6���`'J `�B���@�G�O�j/����z���Mg�{� R��w��Z���kH�<�X�b�*���%\R����>��ԥ)�}��ⴥ'��|Q�@���r!B��Mlov��h���%�o��)N��~�)JN��߸=J��{�)JP��>D%�!BԔ(�a�W4�iQ$�Tq]��hy;ۃK�\��<�v���j�N�γ����lrr֠ g���m�v����߿pz��W�=���(z�Ͼ���)�}����������[�f�+{5�k|�)O|��A
R��|��P�)�}��┥'~����?2�5��L?9mr�mn��ʷ� ֒!��~��)@��{���)I߾{��S�=���)<��/����j��٫8k|�8=JR�����)JRw����R���~��(I��9A���F'I��_���R������p�Ӻ����);��~��)I"#=�҈�y�%�{.!G�x$��mo&����Ñ��s�چ�1˧;��vJ󵮌ۊ��D6���gz�js7����>�߸qJR��|��R���{�8�)I߾{��JR����z���֍�5��z��)JP��}��F���~��)=��~��)J}�p┍�b�si���6Yw���ig}������=��ԥ���ÊR�=gs6��I ֗_���ݒ�JVڎ��)JT=��~��)J}�p�*P���}��R���~�iJO|���5���Y��Y��k[��)H?y��8�)C��}��R���~��
O|�߸=JR�
#��@�
XB���w����{�.��S���ug� '�Fnvۗ�k�J�n�4d��8�WQڪF�6���o6��d�:��M�Ypki�k��9�V��mm��^��]�+vYގ�0�2H��Mٷ�>��~b���W��A��5P���ɑ{���g�ضM�v��{��I� 4f�l�V��ٳw ��ӎ�x�v�4X�;f�3�<�,E���g`T�6z{k�N�q�DR��~�������}߬����S4x�a�\��]z�WAu������t��p76�Y�r��N��R�ʳZA��-~��k]Hҟy�~�#JR{����R���skz�i�~���),���r�{�z��>�^��R����=��u)J}�p�-_y���)O<~ώU7��Z����Ҕ���pz��>�߸pZR��|��R�/�k߳�R���>|}V�a��Z��|�)O���R����>��ԥ)����┥+�wٵ��i��e��ETR�d��(z�Ͼ��)@	?��߳�Ҕ�}�߸=JR�y��8)I�������Ӷ�X�h�8�H�o.nAͮ�u�A��ŷ1���>)q�3����~N��zNZ�9��R���{�qJR��|��R���{��T	rR������ԤkK�3�Վ�uZ�mY+޴�ZA���߸=G���;X�!����:��?��)J�����R���k߳�~�R!<m5sVT͂�v����:D �[��)JP���}��R���{�pR4���6��ZA�,����h��)�qJR�����R���k߳�R����pz��>�߸qJR���3��*K",���]�{Z���ZY��{֐kJ��<��R���{�)JP���}�8kH5��?0�[�FH��{u�\e�/lt�.��<��qo4�V̎����+�:7�oZ����)JO�����)O���R����>��ԥ)�����4�'}ϟU��m�{ֳz��JS�=���(z�Ͼ��)J}��8�0�{����B�{%ú�M�T�R��5��┥_y���)�5���)���Hg���<:�>����)Q���Ȅck*i��$�%�W\�k���)Q	����┥'�y���)O��\R����>��ԥ)�{��Վ�Ut��d�z�i���k\5���߷��)J���=JR�{���D �Aa/�1I*gCJ��������g��׮��5GNh��o!n�s����Pnz��c�&�jʙ�Ue���⏈�׻|�@�'W�}�ǩJS�u���B����=�Z� ֖/E�n�H;k�K[��Z)JN�|��Q��@�?}�߳�R��}�߸=JR������4�'���c���+"�w{�Z� ֖zf=�JRw�����/����JR����V�kH5��k-��TU�!]��J��|��R����}�)JRu{��lz������^����������)>�}�}V��ۛ��7��z��/����JR���|��R����ﳊR����pz��?�}��G��"g�bj�q�p���v��9�v|�\u��^�7XlZDpY^��w���);����R����ﳊR����pz��/����JR���u��x[���F��ֹ͏R�����k�R����pz��/����JR���>�c�ZA�/?x��r��ki�f��Ҥ��=��ԥ)}��o�S!I����GH�	�7\�A�{���++7�����z��/����JR���Ͼ��)J}�����)I�{��J֖/E�n�n[\R��֐kH4����hz��>�~�\R����=��ԥ)}��o�R��>�X�B��	C��p���,~ֵ��7�f�� �w:l��B���t�4�!qqu�G��i���#���V��[���lWZ����\:"9��s��&���+��T����[jN�W#�qkv|��H���h�C�	]wWrF��f���C��9k��:�;nw'���:)�vyJ��l�{�l������n��Og�v�e;�q���\�.9{W�y"5���/��):s�'����}�������NϷ�����ĺ�i���@F�u���)�Z1�Z�U���x�T�2��X��9��qki�����������=��ԥ)}��o��f-*_l��(��!7:�"*�d��z���)JN��߸=G�I��}����)I������)O�߾��);��4���.%]�WW�"D!�wȅJRu�y���)O�߾��);��fָkH5�w�:�t�PQ[K%��R�`�;�=��Cԥ)�>��\R����=��ԥ2�{��┥���ea\b�+����i���2oZT�'~����)K�~�|R�����2-p֐kK��b�[q�Zr�YTh'��31G.�X<���뫋�e��	�ݺ�k
�\��Z�vY�i��K��k\5�J_{��┥'_g�}��R��=��q�i����r����8�%��iR��������I	�IXV�>R�P�ԥ'���]�z��<�?~��)=��~��$ CJ|{���HImqK��ZA� ��>�E��)O�߾��);��~��)J_{�w� ֐iw��C RYK"�o{�OR�����k�R����pz��/���BI!|�7iGH�#wW ��,���zַ�)JRw����R�؄D�ݾD �A�9�J:D �Nq�޴�ZA����e�Hڀ�E��QU�]4N�y.%4�:�N���Y��9��=�����{{8F��ۛ��7��=JR������)I׹��hz��>�~�\R����=��\5��;�i�dj�)k�[�i��}�}����*
�d�����qJR��}���JR�߾��(}>��9��q2��os{�\5����ɽi����pz��^��:AL�{QéK^���JR����~��:A�/?x��r��ki�f��Ж�);��~��)J_{��┥'^�}��R��=��qJR��<=�5�ѻY�F��-k5�R����}�)JRu�y���)O�߾��);��~��)N����2R�M
	��N�D�j�P�ɠ\�iڸ¨o7Tn�D�D���h��Er�j�޳5��JR���Ͼ��)J}�����)I�~{��JR�߾��)=��Se%�:[s{���i���2pY�);��~��)J_{��┥']�}��R����U7l�{ޭ�Z޸�)I�~{��JR�߾��):�<��R�����k�R���>||F��ۛ��y��z��/����JR���Ͼ��)J}�{���	�]�"��k� �Q<C����:�9�Q�!B3Ӌf�L�UJ�ݗUwȅJRu�y���(�8���~��)<�߿pz��/����JR���j3=��Ǳ��[='-��\^ثq/On1e�xݳ�ێ';=i�Hѣ���c��ms�?|�R�����k�R����pz��&��"D �ߧ�Ҏ�"N`�WSy��ލ�0����)JN��߸=G� R�!�o�"B�ӛ���B���ZZi����%p�v
+u�k\�>���qJR���Ͼ��!�)O����┥'�{��R�����/��5�Z���5��n┿���3�ߴ=JR������)JN��߸=JR[���4�B���U�R+��.��*��9�Q�!ByM�"D ZB����JS�߷�┥']�}��R����{'��A�ΒbC̱q�O���Oh$�����ύ�B�:��[�#f��A�2��H��rI ��H"h"��Q)���Zgxm٭]��̄���q�,�V�F��FD��5�u<Sw�&H��=(��нSH2zˡ�$9�a'6�a���F����l�!��D�D�gsA�<���.�H:'���,A Z�i��n������0L������z=�(bba�"�0������m�"�|������ǲ_V1�i�$�����AA�	��0L�B2!0#	����+��靲�^I�Ļ�}��n�n���0�%��Ɓ <X�E6�2�'Ee��B���_~�_��M�m��:�	8  (����~�M� �` ��        ��m�Yᴬݱ�e����xQ�ǒH�!p�<�}������s4�Ņ��eY��B��ԇ9m���&��	�
���⹜�W��������V��5Ӎ)�	z�p�:�b�G#�vL���n�P���,��Q�h^[mu<�UUU��T�˗�ݭ�Ş�]���s�d<���_`� 5���IH��� �Gi��s�=��z���|���S@:�:�#���ۗr���V�펹n��{gx��q;P�K�UE�5r�����89����9���֪[�Ge�t�R��StQÖR��m̝�ʒ�w*�-�>'m�WOյu���:�;m��N;a�vY��T�$e�N�vS�2��NM"����ݝ7b5O�ғ�P8��v��ZϊK=��/u�.��Y�u&�;05T�&��شic�7�P%�`�J�q�(�6���Hdk��C,��W<:vzی���5،���U*G$�s^�4�q��;�u���e0&(�������z"˞	�n�g�I5�ө>O����5�\�ut��f�3qbxMT��R�L��ͱ�A���pF5�����&�����l{�v�A�� �n����+<��g>�qͬ�ݐ7]'h�T�Ͷ_T̒�K�pl�nm�H��X)�V�U�������T���=�6�-��Ɠp�r�KZv�Ғs��rRi"gH���EvH;19�Z�[kh
�Q�ZŅwE��i�P��T@&�h��R���U����;-o$U�%��Z�� ��Aձ�z�a��6�S�9J; z�V�%���Wjܥj��j�9a5ۺ�55�nv���ü�#T<�lnMȮ�v�%w+sZsm�$�� -3lm��e����۬�+m��a%��(���j_� ��P��s���m�	����E��kiSt�Z�߯�������~���� |���J>
�^� �A���(hD�US��NwǾ>�n�Y-��$ 6esV6L�CC^�<�����Um��/Rm͜n��wj�'��pLʹ���9��)7giЙz_-^6	8��u�h��;�Kf����EHq�wc��+�[�q.��t��ֳ����\��z@�����;nѳ�L;aЛ]�j3϶`2����1��1@Q��$�^[�[6rH/nIΏ�����ݽ���������/�uјG\ތ4Fe���ᛮ�ܽ�h�i�2uA���=�j�K�s��d��}�]���e�n��D �A��x��)O��\R����5��=JR�e7<�A�|G�hUtE��t\��Ge)O��\�):��{�R����ﳊR����pz��/=���o��֍�7�f���R��}���JS�u��Ģ���A��>�߿pz����oND �A	���]J,�j��o\�0z��>�_}�R����=��ԥ)��o�R��}���JS����q���mY+޴�ZA�����%��o�R��}���JS�ˆ���/{�<�JԚ!BZ4�p��[���Ȝ�s��:�9�N�wc��e��e�R;-b�˵��ig�c޴�JN��^��ԥ)��o�R����mk���Z^Y<`�V)%��T�z� .��~��~;{@�@J���1�A		s���8~o{�Ss͈P�d�f)��+
K�F�7��?g����������<�ӝ|���������.�� ^��@}M��֜�~����W ~#5j(�"�U]5}����>��@�O# ^��@��,���bB�3=r�S�70�q��Α]�I�A"z���͢(�m�?=x�|��p���T(Q�yOg�l����E#`Z����g�kh}�}���<���=ԥ%l�{2���Z�.�jn��ٻށ�X�Z�K�����Q�����>ܽ8�^��eMЮ�
���CT(J&v�x�-���.!�������;*��*dUq7W8�\� #R�`���	Rs�=�.�1�9$�Q�X�V���,E��kvHnsK���6� ;p�j�-��MӭWQwQS5���y�f ��'83�����Ŵ"*�r��w�t�9�5��:��`�s�q��t\�'8�Zs�y�f��� =�ye�7\�U
�װ�Oۖ�z�oN�{z�
-��.)�c�8!*�"�J��ਧ�/��{��ʻ�����FQX����f\6 ����� ����go���2�eq7Ԍd�K�{�tm'+�	�p�!m�Z�I��Z�-���K.ֵ�wU�j�X*��n;i�=�S�*Np}i��}�l@nـr�d�*G`������=�Z5���-��nޜ>�>�J >YKuj�e�N)S������>�e�`��}�g8�=�`{�yLq��\��(����G�nـ/r{�%I�|k�Nt���Ј�r2�S`{��9�?kKOY��zۖ�z��8�*Q�by
���zt�3mt��˃� J�����<��tp]qɘ�veYC�v�N�f1���31e�|��v{vk����so�t�Z�	��s�t�c&���Nӧc��\	��
�	5;]�+���/��kÜi8ۍ�qP�z���m{��p��N�R��g���v�U�����Ѯ؞�s�u�vF5��i�W;Wj��V�v�p<�`#u������<�g-��4��������n����M�)�;m<��v���d�aPv���IgVz�F�򷾻�Ν�çE^0?u?�p}i΁���'� ��,���*�]u��3����I���� ~ǽ���x�ry�%Ԣʐ.*.��/'@�v�{���*Npgo��x���[,+����#���@J��_Zs�G��`���YSt+�B�&��2�� ؅nq���oN�{z�"�+���f��0[�Hj�kL���F���v
u��zll&nm���Km$r˧��^��v� �� ^��@J��y(�5$\]�U����\�uW}��m�V�N��	BK�2����X�u���v!BQ&k3�DWP�e����?s�{��8���@�v�x��8(�>�����t�9�5��:t��~�|��h,��M�F��u�k���c��n����{ހ�7<^��嫒݁[���7ɯi�ë'��vy��gq��s���f���)Ec�wo�7M� ����79�@�ӝΝcj��Y
�l�W�=�}�����1�go��ɘ�����w�K"�v
�P��� ̙�`s;}���IpKZ8����@����Ј��rf��ϻ�����i$�i�*rW��Q
�^9��s�3�c�CR������ ~mQ�
첮��*������ ">��O4��5�N���n�`�{[�Pζ�.
wa֮��\��S�t���@ݧ9���p��m�n�h�7W8�Ot��5�N�#@n����,D,5t�a\���1�̉:��� ^I� P���U1qw%�����'Zt��ɽ���`c>���a\`XY�w8�k��ݞ�{���s��N�D�)8��(Q�$�n����iәWW$ܔ\�̗Us�?&�@�� }I:��� ԡB�#P�V�(�E�X]���(�cץ��g��)���:د#���r��=rvŪ^�H��SD�����<�����s�}��Ցf;h���8�NJ�v{2���&�@n����M��"Ғ�] ����?~��=�����fLǰ3����=�{�N�S��r���{�y�f �I���� ||�b!a��
�� �2���2p��<��@�P�D�#��LȦI��۶� ��.ˣ�^f��`��V�SY+�J͂��X�n�'77�}v��x���ૐN�V��v5�6%���d�	�:���j;0��F�F������/}�?k������;%����������ܖ���-d����n�s�q	�F�a���NKq ��Ιv]nv�<X�W9'�n���������e�����'"B7��$�����
/��	���h�͢{e\7lM��9��>]�cq�ڗ;�"��Zn9z���2|���~N��9�$�@�v���<<�+�EQ[f��8�=�h�9�≯l��d��!�WX�!]��Us�>I���ԛ�*Npa�l���&�d��_f\6������x�PD�7������ج��8������d�����｜�7l�	/�3Cj˩E@��
n�j:��0N�v�[��r�>78���6��S����h���V��Tt��ws�3&~{;�g8��dG�?Rn���# 
�ȸ��5��_y�uך X���CC C@0�1��4I�a�4�lE!\���c��Ӏw���fV9�BQ ?�X�Xj��¹y�3&c���d��(�DDD)7kvx���@01cW*d��.,������&�@n���otii-fLǰ1�b��0�1Em����7M� DDDC��h�s�>��p�x��-����j��e'%�Y#��n�w��{��6.��ژ.8�k����w_3�:u����\�������2f=���n�
"!"%��zp�%���+*n��������npԛ���0���-��{����H�NJ�v{��]���������^�$��" MI�D�p�`����;��Ct1���0�b$4�[PAB���Cp:d�Fr٥w�K�M�;N�C˧���F��SG|�t��,�#jӑ�dL�)(���%%`���"F���"�$�B�6P�@��q�1X@�	����w��o�:D�:@�؇ht!iN�E8*�R��qt'_N���O N�#�T}P�&�S�G�!B�,�N!z��gz�nx{1P��WtM�N��h�y���>M,{;=�8��`���������|��>�*Npԛ��[0�{���v���x{q����&��&���/6�28νW1����C����Ͱ=�=���:w�8XW.��3����d�{��sI��{ހ0ku\�T�
Ֆ��n�vy7z��`��T�� ������TV������p�w��p���3�3��?g�׀}�!�[�!]�5sv`A�I��I��ɻ������!��\6�u��*G`�Tpr�yRs�F�ӽ�[0�Ot�D}�q������h��w���Ռ����ɬ.
i��ASy���h��:��e�w�uu�V�E梮&�� ������� �$�#��=�����2��Z��|��� �Y�5���M� �w�� ����eN6Wm6{���zf=��֌}�e����}�X�Xj�����6aD%�{��6s^�@�e��<�}���X�CN�]Z��W�>ɞ��6!�c|Ӏ7���ec��I-C(��-�8 b	 �J�`�X�i�n�2����۷�ޜ mݠ:�fܲ���k���r���n*�H�����9�M���l�;�er�ݶa��u��[V���ٮmg����V��9��X�u��	��Vp�s��b^^��l�-5c�s�Í��|���5��� ��wĚM�5t=�`;�kJ��;����l��lUO���}�|o��	M%�T��F�����ݫZ��5�"��M
��F�3i���k+���8�.��xN�{q� H<m�Wm��{tWAI�������{�|�Л��We�~������@J��Κu�{&C��)K[�ʶ���pZ�� J��Κu�y���}|��˻�V7X�Tv�y�=��{��?�B�$���������R�7WWsQT��j�p:iց��0����}�BS1�fyC *�e�tvr�s�w37�G���o4�9�9�N�T�g�~S�ێn�W"�\�K���:�r��i��F�vG(H��.���ɺ�kf ���*Npt����47l�K�ň��]8Y+��ޞǺ���UAd}��N����k@i_� ^m�s�&���������$�@�v������	Ss�>g�X<�����O{��&���s`/6�@��6D
{�^�ʝbꌰ�v�-���39�>��=����^��p��tߖX&�X�$��ܾ��[���ɜ��vWZηJ��s��;���w����ovȬn�X���� ��1�~���Jٟ|�ot��Nn≫��**쪻����Jـ?6�@<��Z���@UR�`��7w��>��������If�8���b!DFG�
������$�0 �"������������RN�������_{"����+��ғ� ����'z�'8�ot�����v��;!ա:��������,.C����k�ɚE��D:/\<��WWS7u�9I;�<�9��{���#� :�?M��w�����`Z��wx�'9DG� ���ғ��Iށ�L�ڵVXD[k���}���?{&�ZZKF?{�xޞǰ>�_�Q��X��:;y�5�����ɰ1����>���9^�n:�@���y�^���j����VK6?{�xֵ���� ����۬��A$(w7sS{][�ȓZ5S��������ۭ��Je�#�����P�U,�GH������� ����۬JIހ�&Q�L�N6[6>��p�փ癓`u����<��֒@u/����Uc+���@��� ��N�):�5�{����lv
�U��f�Ѥ����/ R��_7�Dz[u�l���&.j@�VQ����Nc��nn�����\����~�Us�����²��`@iTȤL %6�:(������7ie�ݧ� uh눵�)�X4%ـ۠���ude,�(���!�"w�+mĭ�a�EvFQ���N�5��v�J���u���J�(��e�Z<�^��,xu�L�mjD�#����4����i�����
���N�Pl6ӱp	ڗ$��E��:�m�j���ƋK�2�#�d��x�u�X�1��)[n6�l:�['*mD7���w{{��{�o�ߩ����n$SI���Ŷ�.����^���s=�3lvl���v������"�]�ٰ>�~���<̛���^��d�w��(�YYT�]�=-����$��f��Հo����.ņYu%�(E*�Y���|�'X����۬�&qd�VT�[�y��DB��`�����`~�I$D��=�@i�(�"�TZ��	���7�����`��性�������`,��M'QF�c��"�*z4�>��nD˓�3�޲��C ��>������n�z������=�x����΁��u��DuD�����\�j�S$�
�ڻ��� ���~�_(� !�C��~�Y���9&�@�O##�6Np�u5 \U��U�h
y:�7���<���{����ɍ�Ue�lv;f�H��Ǻ�y�ry�} �'X.�.�Z���lj�y�>�ͭ��$��}�������7�T3	�U7VT�r��&��զ̐I�y�z�n-�����.m�{��7��T%"eR�J����o�t�u�o���;���q"a]EYSenVff����|������ ���7�h;�ؙ�Dӎ�-��w��<���"��|*�w�qI�h
Su�(�5�����.n�t����0���@����|��f�� �;���7B�v���p�ry�G�GO7X�7�sy𭿯��;����Y�{ǵ\*�g[�� ��4n��[<3fw���o��<t���qXe�f���������F {�f�fY��QU�E���`s���?(R�JP��\ ���tO������e��q��/8{�����f�}������@LW:��&ʉ.*誸���" =�h<�`�ot�:��CXq�x?#���{����*g�T�JGI���{�}̛a%0�(K=�����. �ެ|����~0v=�ɕ+�tZ�*݇Y��.gLA�<t:�=�3M�\��W�ܛ��fBj��7�sy�4�����:��6��<�
�j�[�^p�3���	BQ��y�2sv���}�̆���4�I���w57k����@������" �s{�w7��l��%�L]T�Z�U×|�CTB��ݮ����y���KKH֏��f�fY��QU�mIuW8���y�x�sy�%I�U������#M>4,��e#{w�ztu��ˤ��f��Ia�+k� ��㤠���noc�@��]XSk�	���[�14':v׮�� �Ł&]��.�<8b�	=�H��E������'И0v��w��KSHI}�>��V[l�N�m�oQ���m[H08�M�   $     �  -��W@#��!l�UJ�*�l��[eMp�1j%�\Vx˝���sfwH��4�[�1�H]^ڵ���k!��۱nY&8�T힯,:bi��Z�b�z����%V�,�ݫ�r;$&�V,���]=���-p乑�ix�R˙�L�` -�i�,����,��lt
�z���ע�Guq��4t��I���1)���4���g*k�U�8�'�����Xʠ�K!5�x���t���n���;]m����5l�#��U:ȦMcO]";���.�GE�\�+��q��ʛf�+!�ݖKn1��#�4�Dgq	�!um9{�>��dV]�d�X,�9�V����u^J,v1�VU9�C����g��QnU�6�"`�- �W�۶�p�ZF*�ێ��ݵ�q�oc�#��e��u	�"�7m���+2�h6ʲ�g8���ڕ��{W@s؆�.�91����l�=)��Ek����\C�� �ٕ^mF^N[ug�Lg����`6z�tgq�#�f�d�S �V�[2]�VtdT����gv5ۡ�Z�tը��iUv��Md�ړ�Һץ���l��]V����Z�� m�6-$�*�e���n�熇='i��04k��n���Cq��$	Vܽ�5P,ق�!�OJ� ��8�LQ[<B̣�4ҭURc=�z*ò��h�/��컶�����պ�2�IqX�y㞆��琣`�$q�D�]����$m��n�VÙ&	ml�]���R�T�B�]�e���9,�4���R��^hZ�L��mN�e����6�R�1��y\b�u1�r쌎m�mP
��U���	lg[q�
�9�6�i÷����Ue���e��lG�T�]J��V�l�]����z��� �d���++�S\5\��`m�l���7k��n�n�Sd���3V��5ku�޺M��p�lD� ��=^ǁи	��}M��z(���hw��k5kF��RK�E �W#gm���#nJp��ݥx�b�L�����uv��&�є���n��D0V�qcst[@;�q��d��<�[��/գ����)�=Wu���l�\��ļʱ� ��u�l59Ƿ�n	�V��O�����X����ch �����t+&��f�x6z�ƣ\�K�	3\����ڹ�6���q�e��{��Ϸ}j.a��d��O^��sdR���'�s�kj�=<��iE^nhW�ZHq���
ۅ�l���y;�{��*Ns�� ����9⌒�:Dʥ��v���� �������y�y $�D�.,������+33@J�����y�x�sy�wǳOi���S��r���}�s9����{���J��Dy�pE��_�Qu7u{�m� {�<��� �s{��&�,Q�D7#������aUnd��b���F|��=A��U��0�;�����p�k������j���i怕'8{���"#�ۻ|�7V���]T���ڮ��:ec�oЩl)�����9*�|����~� ��{7�32ǍZ���Wke���7���6��I怕'8}׏(����c�B���&�������h	Rs�w���9�WsVLIqWw7w��O4�J�����}��`w�fJX�4(2D[d��u�@]"oe��Q���r;<�Dr]�k�Uz�Nu�Qw6V�ffh	Rs�w���6�ih�پ�Y���$UH�i�^���o�ԦCۻ| ���:ec�(@/��C�
��(����� �n��i�W�� �@{�CA��!t��Dd�;S@��G�>ַ�9G���� =��c"dj�U��݇��w/߳@n���=�otͻ�6LŃȚ�7[v��r�|ޞǰi}�o46�0���@��A�����箭<+Ѡ�uoF��\ulrw��{���v�(��	��E��x鹵�/._�'�������<���{�ȏ��� ��r��+nX㐲�w36���g�|����=����O-���܊��RZ���� ;�?٠$�FD�ot6�0�ҘE�w7VV�ffh	'��w���Uw��p�~DS�R�I�8}b��a N�Q�/���\��_���j8�N6�rհ;�s9�>�ͭ�}�c�@̬s�6!D7�([�JU!HLұ��ژ]�ְ�e�P�3#���y�V�j�<�ssl���Wv��RU!Se]���=��\ ��<��� �s{��|�$�����w57k�|��)D������� �36���yY��Tٻw� �'8{��">��ͼ� ��y�>˔�Z���WkU��~�g8ٙ����f���i/z{����L����������<���y��T�����@�C�Kd�B��L�U\����� �t�w��ze�t�����x���ΰ/kcV�r3��k"�	V˳�GUŲ�u	���Лɓ�]ֳj���]l���!"�F���Ǖ*�v�qjKT3�4fv`z��u��^��h%�L�X��`�jok��nm�JVrC�J�'����d��լ�Х��õ�B(�d��wV�5B=��1���[�� �R��������$��.����I���t��J�p�k����$���hm��n��Q$R(WK�(�*�U������e7<�y��"I%���\�O�+D�uINm۽�zf=�ִ��=���@�����<|�ʈ�Q&:��&����4ݯ`{����������g{�v�3���0m��7�4��(�K# =�h	Ss�os{�%J�!�F��Z�l��� ֖��zc�{���y�3�u���9ۘA�,�[q����x�eO;�ugq���A[btd�ֳc�adn��Sf����3��{�΁���$�
$y��@���.U�"�5]�Wk��s9�%� ��F�Kn`�hC�����*��߾�U{�ǽ$�}׎f���ܱ���w320�I急7X�7���1͗��i�K	*�%� ��{7�<��6;��ͼ����dM��UY[����%M� }�}��h���y'�m�����=���*x+���$�W�v.�`X�hob}�s����]u��.&jf&n� ���@��F {�<�">�=�����,B��dn�Yy�;��\�J�����t�vx}��݄�SI&fLA���5U���`�g�uW��ﳗ��<t��M ��~Jd$�F���ϻ�73x�d�9��n�)�{�� KI%�Lǰ9��s�y����S>�{΁���\��R�(������{��ﾈ�9����O4�c��Sx`���pQTӴ�W����96xrV�ث��u��Ӷz��ol�h0Cxd��¦���tm�`���*ns��Z��g8�"�*��ӪZIV�>�1��D��n� �3w�;.%�H�'�V��꒓�����=�8�7�6�0�I�ʥC�*��6�hv��������g8s3k`��s��_�G�>f��VM]�ڠ~E�E{��|�9Wi߿~���h�-��w36� �Z��{پ�Lǰ;�s9�<c�ME$�-l���:.�M����9��X���^묑�e�p&�N�dC,�Uj��j��g�|ޞǀw����>�@�o# ��NB�l����̼�*Np�7��y�<|��$���Mͽ��]���E�\����/߷@�o# =�h
Ru�r��3NX�,�R�� ����ml�:����)�3wii�e�*ʉ�V��� >�1�j�J	mk��^����uW�{�Uڿ?�L��1�$���}��feff���o{���BZ�-��ڶi,P���P�(�1n���f���=� s�`c99o'&��=S���mj�rss�u�rnu����0ݼ��k�!�Siهx���/=�1ێ�u��"�v�e�Ӯ��1��a{mZC��m��45��MW��p� n=�;!�5<.TP� W JڷAu�KH�E�l��aVv��&��U�ay��--%���.h��v���r:�e�3 ��st�����ǚ�z�Nq�k�td��:�Jն�,}������?M���3���2#� ��y�'R�ĕT�q352�j�w�o�؉�u� =�����M�KZ@{�]ȱ����^pi�`����N��otJ�LM�F��[	j��{پ�=�`s��� Zֵ��f���=�=�,���Z�����7I� ����y���M�����&��)7�='7�ܻ�d:\�A�2�.��N�f�_{���/��upT]\��]U��7�i�`{��P���w� ד�[U�E]���.�����~���@|�!c��o���]�Y�~�}U���}ߛ�uDBQ2b�Zl�j�������Z��'���9������O# I�{R�m�JI�����\6}��t��p5$�Q����ڗ�JB�Z���EU�����6���{��??{?^����w��1�u$j[i�!�suѥ���v��cng�1 �xD�F́�w��+�����D)-�|3ٵ�1��w��f�Q��f�z7t���uR�]��*�p>�;��%*$�w� �g����ͭ��fh�&����Rͽ�ހ�[8�����K�#�!i@!�S�����1#�ы�Ěx� @m��1�Y���2��.�!�a�{o�DA�qv'a���N�|�LX�I�y�*;}�"Ӯ�&Q��5 mw�z�Gzt��a����3�
�x���J���h�f-	IKH�R�AQ.�,�ǭ0�y�$>a:A�1�{��zx3��ϧ�t��qN��; $�hiJ	��=@�s�:|P@؃�i{0Q�^�D�z�Ё��@�޷������Uy�w2��j�Ue\��������w����# sܝ����5���Sst]�*j���@o �I$�-3��o�߶�}��pwQ �ń������nz�{,������v3'[�=:9f�ݒV*Wk!)�ʜ�l}���fF ���}�4�F ����*��jʭ�̽��0�ot����,�4�{#�i��b�6�j�V�ϻ����0=�ހӶ`�G*�D�R6U�^�4�F �;�v�W��P�T_������1��1$��^����5M)��LZ�WtU�`{���l����o# ����Y�7���ꮸ�Ӓ���+i��8-��>ţg�c[�˸I� <ڧm���.���o�l,#VJBͽ�߀���ml�����ͭ����^�{����JJ�]\`����|7��9�N����;�c�&JЎB������=�ޑ+f ������ˊ*�SrU����؅
v��@��N ��}�l��sw��7�\�˕Wv����/����-�R�f�������������"(�R|j���,��� �5�Ϋ���cG�p���0���s;Z����i��A֢Nx�f�M��x^K����`��l՛Sn�6L��`]m·�	��F����w/C#���9箢��yذt�"�s�;v	���us�+1=�{\퓦QY�F�hԃ�X�6[�P*"Ӛ���Ktn{=�
����1��^X�gNKh�Q�~w{���w�wN��ǎ�i��Z��p�)�4��^�d�㥶���5�a�Gg�����z�>���psD���]ݘ����7��9�N��� �"9T8*$��(����@|�F ���}�[8����BP������R��*v��v�諵�m�:̶p�Jg}����x��7r��*��o*r�4���|��ot�ml=�f���{�V"+)+D���{�G�}'��$�@|�m��?=���ߖi�U�H:���N�!�ն6cvw;��N�h\�������6ӎ�t�5}�1�p�c�@~v�P�!���� ��,?;Y	H�d�IV�=�{7ΐ_|qx�q��:��*뿾����{6�}���5h�����w{� ��f���}��'��	$�@9�Ĕ#mJ�q��`s33�=�����f�ֱ�2l�}�ka-��@i<�������~�X���r�w���e�*��Y�D�p�%�1:�a�:��<��u�v�J�5ņ4���c�޺��n� $�@s���7�F��{[ �Fbj�
I�v�|{&�֛���0rO4�I9��"��-R�ܳ`s=����ml�kR������6~�yD�B���E$��1�p=���>t��5(�?k���~_���Ԕi�KKm���f�Ƕ�g�}�w� ��|�X�ՖPTnw+��8��\�H��[��W�w8�/]���뜚�uU�9������}��}>���5��@N�rO4N]aS$c%M��%�`s=�� {�˰w��t�7<؅
d�^n+Tڑ\�J����o���ht��ɽ��N!���V�H� ��پ��ɲ��߾����(0�b@v����� {��u��U�~7��6kE�T]M���f�瓬�7� �w�ُ�T%�Ѕ�$ۺ����%½�v⵰�����~��}��p��y1�m�F:��DV�"�>�����8��]�gs?
��6q�p���J���.�EU�>N��O4<�`ɽ�	6cװSN��rP｛�}�-�@'x�r��싻���������u�?&�@'x �'���i��SvXӶ́���p=� x��@s��r"E�!(O{*zk�k��m� 	ӶNE�c�^l�=�R	t��7m0��\<�ed�r�)��%�����Ђ9gW0��H΃�;>ggU��bcE��p�R�#v��!>+3�9�M�Vrgt���3��)n����اDJ���ʐn4�X1ٻ���a�a�i��D��ׇ>�cn�a%�r�pp>P�e͸�s���=��S�����T�]p$�� �?���������`z\\��ܠ��#;��J�sV��n��];�M���.gk��ܯ������e�� �N��o4<�`�{�%R#Q���U�r݀wٙ���ɰ96�@'x �|7E�T]M���9��pco�5(�7� 1��8}�kv��Eaj���6�I'��߽���x����'Xy�vD�au2]�3w{��� �m�瓛��g8���d��4B��B��[e�c��C��f��H�����,�M�xv��/:���:�i-� �ٙ���ɰ;�7� �w�otH�}vE��q;yy��9��=�DE�}�ai�w@N�������4�2Tݖ4�`w��z̶p�Jdǻ��9�\о̊jmH�h��j���+[� ǻ��{�6}����b1E���[#����΁�	mf�p{�ހ�-����(���.�u�@#�v���2u�J��w��xv��-8O֟k�:��Ve��f�盬�ot�� 96�@���e��XZ�i�f��3����l�M���u�w��dIVD��D���z̶p���N���}x��m,,@I�S�p���/h�����5ʻ�7{�1:X9WqSd��*�U���
�=��@������z̶p��#h���Z�.������`~�ִ�ZQ����5�Ӏco���ț�S@JT�u8k)��U+ͻDa��CxbS��p��mp�3\�;�&N*~�_����+f y6�菢>���u�w��dSSjEr�bɫ�@y��l�y��:�n� �c}L��N�E51j�]��]� ���t>n�	DA����3޸l;����)$,wu۽��n�I��V��dz>����c�T�E�Y���p<C�־=���� �߱��+e��V��lM��V� ����7Xz���kv*\�/�r]!���H�]nԥ��=sgm�=�;[��J2��{�4��ɷ���g�}�� rm� ��]d-d%#��Ii��37��� ����l��">}�#ad\�]ܕd���f��X$���f }��� ���N%M��D�l?(���~�������@J3�� ��}N&�H����*�tjـ�y����ot��A2@|E��RB�c�I*`�����uA!�Ld8�DXRU�	�\��v#rS� ੳK��;�$�|��=Ks�(�I:@>�y��������.tX�8{�)�z vnE����>�Uq��#A����+ #)�'�D��9�!ܺ�����3���8~�l�!](��TЉ5$@������u�3��u�D@A#!�T�9�zi
��BC$�����b(b��m!���4�di�����B��hE�^���'f�&B�8�A[
�HHz�*z(�((�T��`P�
,�ȽJJ�u�y�{~ 	m���m�$l )��8���� �` �  (     kv����۳ۧ-mUUl�A���Kk$���:�c��HI!�'rfi�F�GL	�جc�ڽgv�k��[c�x���͓�IK.�諥��6�Q�X�;e��4%��]�����sD�f��!�6���])�+]mNS5�7I� 6��j�fU��&�\jXy�Q��ӧ��\�{]�ӒgL��pu�1I�V)�㓎Bp���-�K8�V6�����Cۭ�wC��;,	��L��]�k�3��z�r�=s��g��NҪ̑9u%�U����l��TI�u�^�h�Z�[�I"	����c�)��h��a��zd�`�n8�.�B0�*���0:�ٱ�^�We��9�<lH!�)s�)��2���i◵��>��4n���r��5�\�,��Խ�=��훫Y�#U���I�Y-�5�0MV������V�y�|�Tt����f�Y� m*�)�<E�RF��q���y�;����&6P_J�U�' z`tE��5��a˸�E;q��qq�`1�]6;	�k�`�ݓt�v�ٕ�mUl.oF���r��l<�jN*�%q�vI�;��N�:Š7kI�p�كٷo"���3Y5۔(�3(t��ݹPm�c�p���H.K��� +^�:jښE�,zج
<����x����tO2�-SUUUPs�{n{i �YE�.#mZ��L����v�-��ѝl�S�"�ڝ�^��J�(�ۦN&U��8��$�xA�����d	ۘ[n:����A���U^�&0PQ-u��v�vV�j�$ַ%im���rlҝ�.�f0���P���B�*���ƫex��ѩz���$K��ݴ���p�s���f�s�[wU�z7����pm��=�5A\�K��YTtlS`��q�C2+v��S�by�3�� #�[B	�L��=�S��F4ͨ��@Ml���Wh{���ï=ACk����x��t���x� $��"@�=����R��]K�.k����'�hYU��m��;U<Z����RN"�t�nS�at+��m��iQ3�^�>����D5V˫mO6���d�ָ�8.�=�vm�{`�h�g,múlul8�H�y5Ǵ�F����>^�Cۗ�t������K���������c����:k�d��V�>6����kJ�a�tH���m���U��%^���� ;;��Q.K���)ɗl�U�D\C���gU�YkY��޳���\G\0�vY8���ף��ӣ���vܩ���J"G��U��i�{�����v��݄DB_��N k�5j�j���,�˚�� \���{�sV� ��7�Z�{��Z+Q��V������`&�h�� �7.Ȓ�.�.≩���;�� 96�@;�����39�<�.�Ka	H�%NZ`&�hsw�rm�������oͿ2�=x����g�V�9n��C�g�kq�;g��p��'���ktr��N^^fhsw�rm���ɷ��z�8;vXKm��fs������b:M���#�&�a$�(Q
>��ק 7=�� ���(@w��vMđq1SU^��ـ�y���ɷ������\E�uwswf rm�w7x&��Gs�`{�1c���K����?{&���w~�ͽ8��s�5y��۫�D�;`v��i8p7�����#'#�:��ηluN�f�_��|�n�M:��~�O��۠>v����@r���ܻ%Z���gr�;칏�c��l�39� �̺�Z�r��J��pc|g@s�뇣�����P�-i+_�>� ���`s���jKBRj���N�M��;f�"S��uު�4St�U�ܕw\����`��:��`�A
�̛��D{3��!�î�4�>Õ��M��2��'�Y�B+	�t�����2���� ��g �;nz��Z�$�!�w{��Z�'h�\]+�����{�=�
!Dɲ�� ǻ����Đ�@�S%�����WD�8t9����ޛ	(��ͽ6����������2��kD�lM��;f��s�1��B�_G���ig.rl}��N<e�-Q9o8�l�9;nt):�96�@�}P?7��KN���۞�N��Ն6cK>�c�5�㞋�Ób�ݒ�}qNsd�7ـrv��Ru�rm��Dh�� ����
(ԕU(��� ��d��7ހ���v��TB�P��]�SAu7Jf�.J������?;gIBP�Ϟ���3v���'&fԊԪ��j�@�v���s����"%7�ހCkQD�+��ww7vp��s�6s7o�c{���p�!�D���m��H �
s��Y��V�)mt%��$k������3Ӈ���v�/���9o�Q��T���jKldm�3ִ٪6�N�,���wE�6έ����c�f7�۵�ov��C�ee��!��s���q[�5�Ɯ-��K��.PAf�oc�v7�(�v����L�����'!Xݵ�tn�L�'GYZ���;��K��J���xcw�_]�8[b�^��u��\[����1��ϕgjW���爱���_^�}���蜼� ���^�7�s�d|��� ｍn�X�,-R�$�`w��� �v���s����B�&��uUsqQ5Sw{�w;f���>���;�fs�yf]b����J���{+s����7�w;f��#p\�ԕU+r�oo��e��%��߾�fޜ�v��P�)�=��	��E������I�v��:�MA��y
S��n<��'f�\q�ʫN���P�[o �g����ـy;n~�����:#�T9�.$V�Y5}��si%
*&b6#�Q�s�oo{= y����@#14A�LU�v�����s ;�˰�>���ot�l������q5u3stN^N�w7x$���ـy;m������n��+rKv}��p�>���v�ɼf�w7x���L���;�6D9 ���Kd�#]�cua��A^�x��ȣ���ŧp�����J�_����ـy7��i��7�C��M8BV�*�9i�>�\���zZ�a����f~�����`s�L�Ej�%�+r��àx�{��ޖ����B��T�P48*I���c�A��_߮��ݿ��g�*Ӂc�;*����>���� M;�7��: �w�tG�*̗E�wU{�	�x��@N��Ot"a���*���ғ���
�#eո[��N|�[Q�݊���k[�ޤ[D��Y[��m���m� �w�w�{�	�x ��8�-9cu�`�v���]�	0�{7�g���w����=�c[�VF�e�V��� ���t4� \�9�Ӽ���&e,v��rG/8�����~�=���gU^����zHL��(
<����˳^Nd �nJ�-��ﯲt4� ~M�&���%��,��o9Y��9�x�g]����/"�nu�\�]�s���+�����L��R�%�+r��o�&�F ���KN��ӝ���
�bv(Y-�`g��� ��d���:i�d�P�rL\IM]��
Zu�>V��	���?&�@>�" �U���́���>��n0���)i� y���&K���������t���;ͽ��� �k�;��yG��$p�I%��UV�mU[��N�<`�v+�^�h�I�n�؀�vU靹.���)ْ�7�K0���s�ΧU���Y]D�n�c+u�����x ����/N����t<GK�:�*$t'i�i�$�{{:P|1�����i�-=�9���fJ�=�j�8��n1��
�8�����`V(s�9�����{eTH�!�m
[����۱��D���뎋�[�ë�F�l=�B��}�W�=��X���t�����������ɰ;ܾ�����={���t)��.�n�Қ�j���� �v�����;ɽ��G�L�?Mc�c���+!m�l�˟� �s6�l(Q1�{��:��|ԍ���UU�W3W;�:��0���-:�}}��w=qV�+��ءe����{�DӼ��@\�F������=����V���z�hx+���c�m��Gfv�]w/.�u����{�Ӽ��@\�F ��� ��X�<�en���ﯱ�-m(G���,��=��ͦӰ��|����� ��|�
"&C7cd�2Zr��R�������[>�g8��]����>���EdMбJ풭����~M�y7x�i΁�<�.�18�;UQ8�/8��.���� ｛[>�g8��x��Ԛ��Gj�JU�ݯJc�v��	�������gr���kZZUn�=�ƥnB�[e�;��|�y>otJn�����*�૙��̝�y>otJn�w/��KZZ�*Ӕqڝ��հ9�{�zSu�FD}�}
DT�_�8����ѫTeV�4���7q)9�6��	�ڇ~v��v��;��xy�����И$+����6�ᷝ ���OYqS����ǰ0�31�#8a�i�I(n@��H8����A���p$�0l^)�9�w��n ڱ�V���	B;��P:}S�F�8(#�����QT��@���OG��D0>�#:>�>t���t���:#�P�d��/�nn�tJn��ӝ�y�I#���p]�� �U��m�ٰ;NtI�`���=)��s�'rc<V�[:أ+�����.�yӸ�=Y{�8bv3�Y}�p�G3�����|\���@�q�ԡv!(�Ƿ�<3?5�E\�b��%[���s���D��{��1���@�c���Y"���R�I����ɰ;칏����ml�39�:�5�d%m���6
'�vz7�\���Cb8���	.DD(�Y�9���<Rf��\���U�W]�'�{1�p�X�w������o ��س���-U���N%�W�v*,���CGa�6����]D�EU�� �otJn�ݷ:}���K�z�*b�ph��|��`	���9'��&�����L��C����.P��ݽ���|\6J"e����z^�pNz��8��乢��4��0�{�zy��o�=��*��#�Z벭����p��k���y�@����>����GH�bD%U>����c�Z�����:l���	�����3�,C�<\\�`#X�-�S�@n�[�*�e&�lmzu�Ur��eݓ���j��݋���nc/�VM��b�@���R34[�lu���
Χ�����u��E�Tt��-ݬM���!��ӯkhun�R+Y�'���	�	�ō�vt�خ��-"M�7��u����n6�*��&�.��Nt�dQ�KI-�[�7v	��Û4Y�8��]ڴpqn!H��N��]Q�l�h�ѸH�<ɔZ���~����p��h���mW�\��s3V]��`7��O# i���3&��ؙ�V�RJ��^l��yM��=-:�o�&���M5sH�(���p?	(S�w~������h���tG��s%đvEAsUW� �w�4�3@\�F �ot�Lx )�����EZuXZ`Z�vR���׵��ki�,��eLD���ƍ�L�]� �x�rym���G���׷�2w#T�$⚛��U�5�=����Do���cM��
y��o�r�Y���;U��*���� ��p؄�DL�����.��)�r]M+�ET�]���P�կk�k��;������ ��^2�:۔!+����:��0�{�i�������߇)p�d��v3�3�����6�]��ۛu�&s�S���,p���3vN�N��<�����w����d5��N��ޫ�4\�u$�%�wk�6��vJ�{^� ���35D)��knd�"�*j�� ��� m�3�b$��"j*������@#�X�*�-��m���À{�ͭ�����ٙv^wX�!�NX�jZ:�4���m�y�xm�4�K����eC*�9�NA�:������t���#g'Qp�'��-���P�t8-Sv����@׻��ͻ��:wٵ�=�18�;$U�Hܷ� �=��Q�M��i�=�����1eF:,Pu�*q��33xpwٵ�3ٙ� }�˰9�&fѨ�	Ii/6t6!%-����w��m��

0۠qOHMΑ#Úa4lJ��oKKW%��8s�i¹\FYWwM��=-��o�$�F��z`�4ӱ�ʣ��Z�"�����f��cne�+YR���D�������8"������۬��I�`<�p]�� <AA��$�́���I�`6�@<ۼK&L��;��wo�{�ͭ����p�����=���5���@�1]1]R����UsWUq�4�� �n���:$�0�y�ǉ�"�2G%���̻��_�y�?�� x��@�D�(P�<Ke������ � ku))�[��H9�s��l|8�se�cq���KU`���ضc����ȷiwit���;dӛvb��_m��}��nN�S��qC��;�3�x�old�9�K4�f�P!j���%�*�&�;(��xώ���Zӆ� ����[mn; mS�Z�9L�J�![  ��n��9����2�5[;Möݤ^;]���w=����߯F6���)��c�v�ӧ�ˋ�%<����!�����Û�l��I<��!a-�������;�f��Ͻ���Q	} y�� ~�&�sd���l���̝�y�otɻ�+Ntj⭑�+���Kj���9�>~̛��@�F�J̗Ys\������`��:��0����刀�Wm��6w�������7�KN��G��#'&��2��zP;Y��6�A\�]�!OB���=��b����uY�ٴ�ƥ�����\6�ot��`��:L��E�D���Z����8��|�;�BH�����\��sbS#m̩��5wsjꊩ*�t~� |�9�;f ���垺2Y!+n��[�3����=�ـ?&�@9�x�qD������*��̝s�`ɽ�i� �^9��DN�t6�e���Sj��GZ��9�]���`x�y�&��ܓ�'f�c������+���-�����s��e��_c���Ծ���2��V��tr�{����� ~M�|�D�(+��l��_c��\6$ � `$D`�;�U�#�" ��>���:�@RӬ����6�[u�`�v�����{3� ��|�;��g�7���]R����U�L՜����l潾������p{^І{	l$�9$C�UJ����6r��wk��=��y|�[c���]C��棣@D�^�4� \�9�;f�7��z���u�T9l�`{����=ܶp�o� ��|�2k�#���)Tݢ��������Zot�w�.W�|�늴�nWAі[)�9���*��߷ʽ����u_�B�(�$�BK�
b!.7���>K��l��,���˻� ����h�� ֛��n���w����
i��̎0���c�62�S��+�R�P��\��u�볱v�$������r��@\����s�v_�x�D��r��,�� �rـkM�sN��c4�L�����T�7)�9��� ;�˰=�_c��\6{����Զ�7\i�y�i� �Zs�.v�[ot_�er
VJT�́�z� �r�9���K�\�h�
>"d�$)HPA��ZZB��a�ヶ�Ԟ!Nd��j�pµ����(�f��f�E���p��t669:��R�j��ېF�"��mw��ܹ�)C�(JN�-j*np�SP�Q2DHz�)�$�����;�M�*$ф��B� �(�SL�436ǌ��ܝt��ST��Ì*d�d�P]8d�!B�[�BtN�[�v�u�ٚ""֣ �(���DA1�Q$ A���n�7MA�!��n h��0I,h�I֌5�H���F@HE'�x*�TPѯ�]�M�Fbtn=B'�l*��\�!3(($	3x�0�8ƍz�1w�)��}/�뾀��n�� [Am(  �m�h0 9�� m����       M��$���r��$ K),�^́i�T�I�B��^��4U]a�"d��v��fl=r�6?�|d�����`�qz��c*#�*��3�֒*N�mI)���"f]Ut\��K�5hM(�h��ܸ�ٴL55:�M��)V�aԫUT�5qm��7b��n���_.��O��\��A�6�6۲������ؚ�z[6ݫ9m�6-H�Bt0����8l�w\1T�mv���ն��j�1����l��=j��x��pm�i
�Ã3�8S%��{1�z�e{[��y�}���n�(ܨ����Zx�4y��ܯX�!���.w]FA��D�<A)�u��u+�R�5 ���up=Pr�9���傛��'*��X	
�#��+Ciַ����E���kG�g�P��0�^����dcx�C�yY��6%�mxM;��0���
@�\�Me���*\�]�f\��i��kqM�joVFKh�ݻ`��v�(R�\�l[f��\Vmzۢ��v�����폱��JӘ5�V8nYn����fL�;N��VV�@.]��ǹ�u۷6��eQ`{-K�=��vVS"^�ӱ�zÉl���c�٧=�V���4]��I��$󂌎M��\sY5[j:��4���s��t�p&^v�6��+�8ԷV�al  D�i%�QSgҧ].��5�la�Km��z���h�|w8Я��i٢�4��tA��k�`������x��z����
y�q��6- �-M�> ��ml����%�H�K��$�-*�N6�Y0ɶâ�^�l@X�ŻX*�����
�)���3�����ťeT\>�d���
 Ҍ��A�8x�]�@v���`�m�`t�UA��:��t���&��';RԐ�T��D�f�
]���R�]�qBCr����U]q���V��F�ݢ���������b�{� �D�
$
b{���G�iu���q0H|^������x$�����m�]��_��|}���ӵ���5�<�5�8��sS�+S�<�֨3%XJ�#Z��������b&��A�U�Ψ���l�.�n f6��K	��<3�>.^�bZ���'1۫��g�G�Z�#�kxהل�]ɹ�<�q�2�'L6���9���Hx���6 ؞�e�8ۮ �s�D�!��d�ײ�M�ݝʹ�+7Z��_=��:���q�L�ֵ�o0��q�V���c4Ջ�S=gi�Ѥ�K9�e$��Eב�[�Qډe��oo �\6339�:��6���|�늴�nWAі]՘����#�O���ݿӠ.v�ؙ1/6�d-Ie�U�U�zN�����zl(��2�oN���z���_��e��]�`	+Nt�ـkm� ��d�zb�1D��r��,�� \����4� IZs�y������2�Y�c�]qbv[��ή\���[�n���tq��Mn�!0��Kؔ�a&��=���۠t�� IZs�.v���ף���Y[i�y����t��V�ZP�'�'��o��3��g;����b��~r�+"��n������� ^m�sN��T��.���uv_y��l(���8����z^:�lB�{�Ӡf��r������$���0M��:Zu�ro�)�� �Aۿ����,���;k�	�Bx�MV����X{��
�����y��5��M���-:�97���u�rm�k�X�5A:[l�́�fo~Zֵ�G9�\���z^:�z�1�*dȚ�.���k0��u�rm��!Gѹi
����߶���i�3����7Eګ�������ߺN�����Ϲ�`s�z<QKjuF^�K�\b!,{���V��co�6ߟ׃�&9}�G9�p�d��o�M�i��<9��-�1�]�����˞�]�nz�.M�4����{�t��`{�G��Z�Ij%��y��{�1���L��w�'^� �7�t<��T�sW4d������{�t�� ��3@�fc�%�yLaS)^�v��KQ
'+^� ǻ�:z���Kй0��!0$' ����������1�2�m�ٰ;�����npM��:Zu�s�0�
>�$�Rqm˭��1���=�ۚ���՗��wO!��ڶ�F�*ٺDٴ兊Y\�\Ϲ� ��� ���{L��u7S7j�jj�x����$��f���~����{�w�R<R[SUX�9y�<w�=�����%2�g�c����=1���V���[�;�������96�@9�x��ws1Uw]]���h���96�@9�x'�>��a�2A쿤\��}�a��v�$�o0 N�;fU�8�ʴ�n����R�$�ݮ���#����Qe��o:Rg=N狪�ͭÙn���<sq��c��ֻ<\�[���9zP��Y{M��;����m�ău�Xŵ�8a�}�R%9sG��<�m�ڱ��v�|k���.	ϕv���vx�c!n��#����]�礮Q�u�u�E�u9�V�<k����L#���KJ�G8ا��
��:�kL'</C�B�֪p�u�xbv�7>���Kk���3e�v,�4~����n�sN�M�4����I)�*e+ԣ��p���kI������n� �6�ݙmhT��`�������	����O7X&��4� �g���M�NXX�����}̛����<w��	)z��t��V��ɛ�J�́��g8��]����|���`g�{,�(A��Rҧb4J�+lpk�X�6�-܀����w=�(q�U%��;#/8?{&��{7� ��ɰ=��� <���B)hG,�`c��wc�y%	BWf�n� {�����6��y̵�Ԗ�YB^l�����{�9I� �x���T�Q.�l�l�����4��4� M<g ��d�K3�c
�J�+v�� sN���h
y��m��)gm��<m���i�X��5�5��'9A�^�c�[W9V����e|�l��m����o�.�� M����?׀%N0�H����-����ǰ=��� w=�`{37� ���0Uѻ�J�j�x6�z��R^BDW)%��DDq$�GTD����ώ��� ��(�)-���Iy���ff����{ٙ���zc��)X��rYw�&�3@}M� �ot�� P�~����.��s5��k��Յy[��\���덹�Z�^Z�d�{*�t	Y����4���	��@N���p�b���,�%q�f��fg8 �w�&�3@}M����!q%�1E����4�����Ss�6��@#10�%ł�WW5uw�؈R�w�t�ݞ��CIpY�LI�!%�y{����]le52�U�t�����������I� �x�������??l�F�����:��h�����*F:\���4D�뵶8��l�G0ۢ�37qW55W:��~� i;�O�>�ǰ=���1Im��d`�� 3���O�>�� M�����~����KX�݁��~��gfc�#ٙ��{�v���I1U[��YB^l����m���;�l���2�F��9\@��Z��39������3�?Ss�:�؂<�H%��|��|!� m�:l��4�pk�z�q�..���v�l���n��ne�):�����i�[��p$k��-�}�l՗�`��s��z��NHw\�ыF�K�sp/ E�:��?dݡ��+��fN��O8��_4:INN��9��k˼s��͚5�x�(������!rE��F�3����!�!�>�#m\��$;t����ܰ6k7�u��֧Yh�| �A]:ZZ���>�F=2���)Yju]����uc�'.��Ø�����uGc�/s\�++R�[.� ~�f]���7� ��ǰ;�fs���c�PevW,�`|��h���9&�@N� �_*i�{D�vW\�����`w��� 3�˰>�f����tn��R�䳀rm�4����h?���8Y�R?�Im,���{�v��2٠>�� ���c��&&P�&��"��:q�;6����,��C�a�[�<�չ9���2�J�qBV2R9,��wٛX�%8�,�ܯ ��@�������浙��uW�kﳟ
t��a����(@@�	AI2ҁJ�����)Ҁu}�}��U^{�v}��8kA��Q�<r���+�[��ot�� ��3@}M�脔S��"˘��nn�@N�M�4��`�{�%*Iq��]\���ɼf�������ot�� ������ɮ�Lc��7e�@н�����Տ<yH�G�)�v���.o��}d�}؜E]\�a�>o# ��� i;�97����te��V䖭��fg8 �w�ro�9��>�;��*��Ur��F^p=����2kTֵ�� ���iL@�8�l1��\<�N���p�TE"�4L�2������d�c��=�䩆ݚS� ����:E�.=�`}�&@���zދ�E�5bRR���I�Q^��E!C��=���C���
������0i,���Z3|.kj���z��J�̌�٬��O��흏��@x�������-	"a(�"	��P�:��}��$��&Bj�L�D�T'��G�8�+��r�a������H����1�� �HtIZ�B����0g ���;v�҆c�#�.�̀8zR�7j�Né��^���՝�Z1u�⧊�PٰP�hh�Q.��ڈ� m�>*:CZ��bP�=�<N*S`�qW�ֵ��9ܛ�{�� {Lv��+�UM]]�6���g7k�{}�j��&�f~��{�Oʪ8J���~���� 96�@N�M�4�ߍ/g�۱��8�V�݇	/]�Jj��c�3�������+v��<�He�O���ɷ� ���97����zA~��p���~aX�^�N�y�w2��������{�
"bBZ$�WN�W,�`{?~��c�d��fs��e�vyx��C�:�Ies{8>�\1�ހ<�|
���JT
"cg�.�%R Ħ$���14� �A	i"P� ӦC��66	� cD1�X�8�b���K$`ʙV�B��CP�Gb7��t��5���K��*�h���m�4����p}̛�״&�c���!T�����VΘ��x������ڮs�(M�k���$1�J�B+#C�� �{.��fo���`{��� =��:X���H���|gu)�6q�p��z ����L��7U[aeR�T���o�:�=����>N�6���2T����&��� I7� �;�<��h~���-�{\�6�l�Ȭ���uu}��;�<��hy:�M�~�����I���~��K,���B@�\�AW�&�a�oc�Yӆ�Gv�kFbT��-<�'Y�e?r��z׌I�x�s#�k�nf�a�m����ӳ�Q��v�:'a�[���z��e��nM�b�ܒ�u���<,\a'v��gأM�4��qã����ݱ�CZ� �bm�m�۝>xݫI��9�c*��ٶCm�R���\W���x����8�s9U����USa��#��ֳ5ff����[��C�m�npч��Q��.�'��.��l^�a����m������ ��d���9����b�1F��u����a�9��#�;�{�����f�������uZ�nY�;��� ��:�;��h	�s�w%$UK����bꤪ��KN����78;p�=1��X�$��́��o�M�����'XyD�ue�Q^�r��1sNk������kLl�`�u�j�mu(��Z�Q[�IiZrTՖ�y��}�p���):�=��4t�J�nX�bu�-{��g9����kI,Z���B���GK��� �����|���1�b�j�����d��<f��M�ܓ� ��0�\�sud�]`��4*np���):�=���)��:K+���>��{ J=�o�Ә�}��΁��-�hRw�~��*f��ix�8.�ֲ��z��������7����Ǫ���ȝ#n����#����):�=ͽ�ʛ��)$y	l�e��]��~�M��s3��}��{��p�H���Km�9D�]p����e7<1B�)�Bp5�!\���f�7�'�!�8�%J!t|��z��\�bn��+NJ������zf=���3���ɰ>�fqp��"x��[���=�o�b	e7��=����>�nx������Bi��b��I*��4��d�*a�u���J)�;Uٝ�]��F�.~������'X����ySs�w}�� k��#2�U�G%���g��M�ܛ��'Y�|�P�qS�Iq1ussW��ySs�w&�@�Í�s3��{���tc��+dr��ܛ��'X�����}��D}�@���� �ҿ �w�������r<��P��c�^p�{&������f��|�n� ��}�z&q;��U�q�7�u֪�Wx]�a��<;�7�K�%;����'c�DHJI]�(J۔rK6{��]��{;��-�ph��U]�15WWs7{�78sot�9�=��Wv��I�Tܔ�f��WJ虪������y��g3wz�m=�脔S��"˟��jn�@7xsoW@�s��9���@#5hT�D\��������ƁG:Np�{���f��Z�1G	����U 	���3��f�z�-��a$��ځΗ���̓n��]u�3�5셒TL�,2GiZ�ؚ�OMt��zKv8L7<n�����pZ2�v�v���LKe���u�6���`��K �x�n��=]�h��9�lr�����.�[�����m���0�ȎG=��ɷ<��8��ś�x�}�G�Ԯ��c�\j��35��y�j��  ��pL��7�v��&vZ�n�u���0j�
ܢ�Y}lg[<��Vղ�)��w��&>��<����t�W�� y����������pߗ���WF;J�l�W�3��� 7x�oc@�I�G� ��MT�*��
������������9�s�}�fs����T%mڜ�;n��&�4t��I�����8n��+NZ5e	o �Oc�֖���7��w�>�o��jt�E�J�B�����LA�p.�F��5qmK�8�ً��7=��*9��'Y��j�nK_ �g����� �M�h�9�99QN$.Cv������U^������6 �Ah�F�4��t`pHak��!�]{���꯼��g*���� 5�X��U�\v݁���ŠsV���<�{����(C�1�rP�KG.� �z�>��9�<��6��g �Y\�[۴�V��p$��
y��<�{5l�#�~L<;��n*X�J������2�$��v�[�WK�
m�/=�O���XS�5I3sWUWW� ���<��hճ ��g8���uH�;T��m�{ٜ���`I�����8n��˙*옪���4jـy&�M���}����!)*bЇA,��C�D���h{P�w��o�u������Fy3-q
�`ܶ��{3� ���<����D�X����$++�n[� {��`}�_�v��1��j��΀Y��RJ���/6.�v����uY�S8z�OZ�m��,����&�հ�u*�]��݁�ˆ��ݾ6�� \�����'	�����/0�9�f �Otsw�jV�%��lCn�T�G)�3��s��e��7�e�`w=p�����R[,m�S3W}�l$�D��v���8��Õ���R`!�	�t,J1'�E\�� ۙ��n�L�Mڪ&�� ԭ�Z0�{�)�� ��bń���ʋm�R���I� �:�ӥ����ͨ�v\nizA��J�R�A�������@歘I=��u�#~�0�2�=�O�e��U�r�l�'����~���0.�c�99j~L++�����~����>�o����g8�6�V
��̈́A�e��>�^�7ކ���7k���j�	�j��Ut_8t<�p�
!k{��nՁ�z�p���R��$� ��T  �?��#�l@A����7U@C@y �"g��PK��w�T  
�׼�?����������:���^׿�������<������q���k�������  ��������  ��QQ�?��?�?���C<���_������@  ����?������u�wa����_�����aBP&Q �e	����YD��P$�HU�	YD�Q %�J(T%�H�I	D�D�	D��%!�H`FD�D��F%`Re`Rah�
T�FaT�F� F%	���eD�XQ A�YQ(@YFTIYQ !D�H�%D��%H	D��B�ZHHRB$!RP %	I	H	$
�	�����d$E��E��Q��BB�%��Pi
B�(�"B		��RB��BT�!a  $!��BBB@���B	��(IY	B@���B�YAeQ$!BABBABD�$XI@�BFB�%�%���!d!!	%�HB��	@��P��$���d
BIIB	$	!��@��$HP�B 	@	A�!TY@�@�	@��	%
 �	�� ��$$	BR���YB@���%@�P�$		U_�1Q� T!EdQ� @�IQ!� @�% $PI@�P!XUB@XBDd	@�%B �XBIEYBQdV@��!!	!
BBI@��deBU�%�$dTRP�$	HFdR@��`�(PB� �dHBEda�aPV�aU	@FP!P�!HF@�!%		B$�b@�FYF�$	��d�d�)FA�Q�T�`R�$%$$eA�	FP!VQ�YTHFQF@�F$��@�@�P! B@�!V!$��	H��P!@��	P%	@��	@�D�P I@�!X��I@�Q��6�����  G�?����W�٣���� � �nS�^?��?���o������  ��>:�����  
� �������� ��g~6�@ �xk�y�8fgg�l��=w��o����Og`  ��?��?�  ?��O���_��`  ��  �Fy9G�����3���������x{��G?� � :.�����l�h��~<�� � �?�w_�u�ǜ  �������������������d�Me)�dn�f�A@��̟\��|>�@t�    � �  
   t�   �� �HTPP*
TRUTR@� R�*��U���J 	QEEIB�D����I�   A@�
@P*�,`]���m���֮,�N])y��y���.���y�o'x��ֹ�m[��ζܷjW6�  �^[�[k��׻� <��m�z�����u�C_^���{�x��5���z��e9nm�  {�P�  ŀ ���.�SM7}ǥ(���: q:tpGO`���(�s��bi�E8���� �� =;��(:oy΀ =.`��{�O@s� �:zR����R�h������� ���4�A�:\�t @Ӧ���H��    j��:R�z:h�(w��W���5v��(>��_O���}/-N��;�^��4{� ��s��i�;�� j�����=ݪ��폽������um�������n r帷R�׼��W�K����Լ ��   D�� o�����gW�N��u'nmƯx�=�ҷ6}���{��U�n���_x �^۝�[�y5�{���^���b{Ͼ <�Җm_Ys�]�-�o�^{R����+���sj}���t�����k����  P    ��N[��<��W�z�����8�����nN�m�5�z�5��Խ���ﾔ��m^�v�  n�n�x;���k�����6����j�׼����,������My����ɯ{:���m����J�    ����J�Pd21�����ʔ�A�F�"x�T�'�H   ��U)FMT @�����)P  �R�� ��>D��?������n�jN���;��_�PQU�]��]"(
��ꂊ���_�TU`�����?ْ,��xb��$g���j7z?�B,@*��qr~_O:�`�G���~~?|�p���#s6o#�X���I�}G��	m˫?0 ����NK)�������:q�u�������7�j	�h��q��A�%���_߿�K		&��g?||��]�Lk+��s��̃A�N��q�!�)��O���A������?' Sxa�u��n��I$$��$D(c
h�2\���.�6C HJ0,�~���d�3����8Jn,F$t�%0+M.���]4�J0�y�)ffa���y�|�������ā>l��9���џ�-n�U1SBi�b����WILB���'�3���:��~M@�
d��J�HD#��5$ 6
T`���r�	�r��͐�y��%L���}`��p��b�1h�c�%0�b��)���%y�!�3������˳8���$��;����ic��i>� ��{�ެsT�:������iW�^q_�̒3���	a���H��s`h6|���s���mN:�Y���;�a����
ׄ�h��C�5�A,�)��e	!!�V45���M�!�No��f�M����_l�R���b��"��b�#B��|%��~��B#	p%�I �d4�!F,YD��-Pvg�R�{S�l?g��;~%�����L���FLB���\�?��1N�/�O�?˕q&�Yi��Y @8/-��I l� �����f%��D�D�I H,x��"�ܒ��&����$)���r|���E��!Y_�	����<?2</�3��S�f���w�.�<;���4l��1M�K>ָs���ԊHI#1bH�w��1�0!�0��%0'�W$���j_���$���!H�`,"@J�I���3Fٛ��l>Y$�Ja F1J�c���tF4i&� �3X��v��a+7�w�B8ć�H�B�:9#dB�9@n!��a&���%���
J0�JI2"�@$cR���ap!!&o;�\��r���HFD���
��+���V3A4�JZdli)3[:r$IB0�L�BD���$RH���̻!u��K�+��	0�T��.���,,a2\J�f��9y�CY�|o����-$�y9�����!��6�R��|F˭�.�y� �"u@�<�)�4ə6�ra}J�e�|	\ �����H���-H�!!@�He20%Q �5�n�5�35�f�nY��H5�d�vr�O��S�IK���䍦l9Û�����'�!� @��M`B���G|���H�s���i�7lk(�?�b��$b��'I��p��$��f�S����)�����ٮ�+��\�+���MB�S�F�Ƒ�a
�&�h$&I.$���$�0�$��c)�
Ń
��
¤+@�HV5�T�� hj��u�$+A��BD!$!0K)B�t��6�6��Ѿ�~ѹ9� ���7�����сin����W�)�CW|�n$sF���7�t�sI
KV$b@����X�)�~IW��
aа��|}ƻ�f�C�,2)��"h�$����Z�۳��\5�I �9��h�G3�)R!i�D�#w�h������*bBl*P���B�M�$m'4��B�MN��܆.���`K�B0�)�L��ގ�T�`R2�'tkR�$Bj��?\֝�,�2�?p���4Y8jP�v)(� ��į�sP��z�L����!Yub�#�?~��k�|L*dJ�@���	n�ro� bI*,K�P�ti�����hH�P+�����75揕6wK
;Ir��*D�#	fn~�|����40#q��>�sFfgi��8d0�H,JZ$H,"����tP��B1ޥa$X�2qW��dJ�����5�6=&7ˣ�@1.���)�?�l���1!A �K�t'Є��41,��>��d�4BO��K�$�7��3���`5!y�ܺv�x�!�g&b'*� ��T4@�p�H~���d]5��#Y$�#S"P� �s�ϳNӃ @��C"�Ō�a��bB@艤��"ՃX��8�;!hF:eՄ�`��e:B� ��)*��f��.��0�.�HR�&e1%ѾI6Lw��iHۧZD97������[��"��
@!�7'����l�JF��Cqc�sl��T��C�r1$��˓HbMpU~��Wj��H��S�8�Ň�'�E�x�ta��Y
~���5�bCG�/�8i��w�`iRe�@�,�������	1���I��_�(E�2�;Ԍ��"I"D��"��I�?��~�+)�Vj�C��5�����Hʱۭ$�#�77��	0��p� �$�b�bh����n`��k?}iXBH��
F$.o7xh�i4U�4#X%RZ@h`�b�bE��x|x�J,d�������
Hc�fύ�ղ͋P67�4|��}��m�]��!��o)���d����H�5�&�0� "�T��G�Rܥ%5��9��a���
�H$J�7�]��H�Ja������_�I^&��^$a���ok{�X� ��D������@�����$4ϸ�c�Y�~>��B��/D8!P��D��e)���$Ja,0��u_���k[�1�`��������bCB�I�T�H0�����K�Ng��C �S��C�����3�fWx��ެ�ȫ]�ʼ�ר��BD��4!IsM�D�oy�a$�o|��5����ȽG�m����� �_���>֝��O�H?��(}�H2BA�@�Hl���H�#H�X�ލm���L���7 ����L]j�a���$��$.䦍�"�3rI?\���; ~����U��ɝ�u'>���#9օ�v$�A߈K�f�8�aR.��,�~$O�(�Bvtm����CVǇ5
7��5���9����m:�vF�5sRJ�/#&s��ך��HS�$9>I\ԑ��-�%N��/䰡L�@#����Z�2%IR$���0�d��T�e1 �)�Id	\�9�1�c��:~:~6������D9�|- ��3���b��Y B9?`X-���0���~O�ôܮi�@�D����a�h����l�2�4
��`G� ~���A#.&�����[�|�����HQ���͹ ����2Cn�p�:6$�a���@?��|7g\5�֍n���4��HJ$�����Ru�Ć����us�߀�CIx}�a.n��g6˭�i:S4�V�]�)�~n�D1�I���$�C5��|�8a�����	�ŁBA������ē��r���N��,9�_��]�gHH� �M}��� hH���}�2BE�ub51�vL��f�>1#���i�m�HCR�˟�o9�u�G2BHȔH	;�}��@���"ƒ8F㣌3[:t�`C1��!W&��~~,�����$L��
]�N0x�ͣ$����FS4B�$,BȚ4�R�Id�����Wl��Q5��Fi�1���Yq @�zn�w���Id���L��}���g�5����٣0�i�$"ŉ�
�B8S����H��S4��&�s��M��nz�r\~�	h����	5�y�f��-LH��j�U!�>��Ϗ�~UU�J� 4� �"�4���?�:O�ƹ��k�p!\칡�%u�H��������l1ևp���C��}���{��v��(0�
�&vٛ��R!F	�|�	P�LB~#)�0��IrF0���'��_\�!}������m��?�&\��m�� m�   �           ���                  �  ��  m  h    �`    � |  �             /Z  �J    �|                       �` 8�� �H�Pf�����ە�+i6�� ����T�^P�j55A��X��  m�m���m��Z�ܓ`m� ڶ� m�٭�� �[��?G ݤ�	v�  ��촒���bB�-�Mc��E�vؒ�v�^�U������:��U-E	�f�n��K+�FC�ķ]U:��T�)<�mT��ٻgp|/��*L	�\����&Δ��v�\	 ����6Z��$$8�� m�z�XkM� 	i�����ֺ4m�����"ى����a�ʶ��)Z�\��U�R�Pm�k[�,��m�m-���#�h���m��   .�$[Csk��m��Y,�^���f��kh�m�&�&�6�� �kd�� Ŵ5V�[N ��m�4R������-�	j۶e�e�j�(�j�����6�&m��۶�Ky4�ʵ\����k�m�)�\�`�`8�	    l����v֭��I&��J� UU@iY^�@my��l�m�Xkz�on� ��%���ݶ��mݤ��Ͱ 	-���Sm�[F�cX��)n����Ŵ;wn�f�26�T^P�t�7m�m� �H�q�kn;m�嶇i0�p�$W$��Ć�H��A�� �`Hm�-��ͤ�m ݫ"�m�u��l�l�UV1*�hl`
��
 ���ko[�T�U*�T	�
�h6.����㮀�V��������Y�Pu1�:���O��x�7Fِ�V{qXUָ�*�*��Kĵ��%�m�le�c�86e�흔�^s�ݹn�ȵ]}��n�����:��T-6�H�\Y��$p<�����KVy��~��[�}�� $�dΚcn�@-����]k�K(8�@�IoP6ۖ��]��*��1��mJ� $$m��n�2޶��h Vm�g�������V7 ��lpް�K�(���pʱ�4��cl K˒:8*yT:e^��K� ʫ���uWV�]�C h��mձmNO(l�2,�6ۤ[@ �kMj��   �  �@  -�ky4�:~�}�������I$��}��߀s� %����j��( �XH��e���<.�YjڨfȂ�t�UT ��H��m�n��#2� �T�
�vU�n�l� H2[���l:���UV��km�8�6ѭ`��-�m�%.UU��^[����j�<ؐ�@[@ [@ZUT�v�+pMJ�^��S
��( �n��Ov���*��Z�UZ�ZWA�n�Ӷ�n��`T�Jݤr8-�	dkh����E]�����ZWl$mKwi6���l7�k'H�@�m J�PR&��@eZA
�yN
C����MV���[���˰TY�RRڧ���X���8wj�{lU�����5�uK�n��z�jѧY�ّ�s�۞��<�J=TK6�X+����$&��ۖ��2@�*�SoQG*�P/���|��(�|��^�6%���A�UV�2�*�8�1��^�y�*���
�Ͷ�ZHjZi6�j��XrԪ�l��CZ�$�-��p�km��*U�bKM�k&Ŵ���֍n;mm� 6ؐX-`8� l��@������^v�n�4�Cm�^�	m�HI�� m�i"K�歃�>/[w� ��jۋn�4��\�&E,5�2��m�p����.��b�lԵ�[��;e�K��` [Gm�m�ږ� 	n��a d�,-�::٫l9��@k 6� 6�#vQi�6�e��A�ɶ��	�m����-�ڶ���-�� �`֛lm�v+U)�����Q���}?,lAm�B���ڤֹJ�,6m�JI�l[]T�YI6J��pU:Pp ���A���p���8`  p m�:� u�v�ii�W���?UgdWe�+V�YA���6��J��ȵ�����5mUR��UPqP3̪핐9�� j�Z��v�����vD1"Cn���Β_!��m j օV��Ypnշ$m[k���l� ��R��(&�ɪ�a�a��N	�U�h� �5^�X���R[nD�U�h��o@�\�ɴ����(l��V0X���&�1۶^9�S@v]����:q��Z�K=��I����˝�p# *�T� ���k�Hݶ$�k�u�t���	�� d��!5�S��Ŕ*��lԞ�ٳl9����r�h���ói$�[wm���  Zm��]'͖@  ����e�p:tmlN[����  [x	 ۤ݀m� 	8  �kgt�h6�+v8[��}���0WUQD���m�p��
���V�V���㳥̐�A� prdf�p 9�M�D��m�l��i�T�gd�m�� ��m�9����U$i. �BE��&�m�$.���*��V꠭`v�48K�\"�W ��t�e\ 
��$�v��N�6Uk��Ym`{[q5XC�������nݶQ�!Ƒ��U�RT*�f����ΐ����$��sm��BXi0H�%���u��Wv٪8 �#m�^�i0m[�k9m��l�������ɭbE�����q@
���P6��U�`%Z��Z�bJ$�:	7m�ۧbL�W[  �mp*+��쪵ʦ���T�P  �[V�+����m\�9^�W�j���2���QH!K<��in6�8�h$ �λf̓hP���<,�R�U*�=.�Kp#�JWU.�F�iUJ�rgd
�6j�6�F��ܫ*�9�&��d7'��.�*�ljzPb���g��y"����5�����K��;F�j�Dk<�nm ҭ��۪�V��������Mt3�Y�t�[�6�Ϟс�R@C�,� 7j��e�q���G<�؝͑VX*�p
D�j8���r�mue���`#���c�[h�l�UUU �u*�md�i[�lY#8m�� :x`vZBm�t�5[��@X���M��-�-���i0лg`H-��8;I� k��t�KtƄ�j�����K�09��阶�a�t $к�m�� ��cI��@:@�M��@   [m� �Kh�k�*6��V�l\=�W��Z�^\�UU�]hHmm�b�/a�X��uYӚUcv�UQmE�fݶp�v� J-��m�ai��ض�ۯZ�L   ��8*ڥm�ڪ^^����ܜ-4�t��m]6V�	��l �`��"Vml쭱U��.X�j���UZmm��Ͷ8kո�z�J��,P O+UU�T��r�*<��P���5Q����U"�YvK�)R�"Y&���[$<�m\ѓe�\�pU��m���K(�A"�;Z˄�Fۉ ��H�5�%V@V��L!Ѱ������RxT��*R�Mհ��ֱc̫Tl�\���T�-U������
(
�B�a����JV�wn�X��M�-Ss�se�]5�e΃:(ޓv��]���Mʒ��UU�j:��%��d[mY5ռ�v��4���`��\�� 9m��U��[@��d��(-�T�Ma�4R@q�v�m��l �6�sm�I%Uvk�v^kj����
�`HI��ܒ�	3�7m�����  � $�f��ݮ^����ÀH �ZbF �m��-$ �&Ӥ��J �+�z\[@�sl�Vj��kh�[H�r��R�U#�7��J;aV�R�n���R@�2��Jƪ�[��~���t��� m��� �ݱ������6� ��啪UU�U�]�r-����V��jUS'U�mm:l�Z` ��i -)@m��հַ[�H  ����` %��ݳm�,m�h�v� �I� �ګ���$��mm��*�n� �J�G�����8���~� �k�+e
���ۀi�rq��˵�!ݰ��8�q�Zn�$0�5]�2����J��4`f�Ȇ�[%�0.�\sv�x��d*�6J��p�β�D�Mm6�k[m�Jm��l8�n� UUU.�T�O@-@UWG���kmm�6�K�	 5��A�@�[H-��K+n�m� mٶzӧj���I�M�h]L9j 
��ӧ)��$��y�s�[V��;����k��"ղ�e[��T�3��f�i�'���:|/+R���mv^��6��c�mYm���ٶ zKm��ݴ�9"A�h����k�ͤ�MP!$|����\6ت��8*��W�W�|��|q� B�i4��p�R� ��i��w����{��_�*�-�������V�@�B?�S�X�V���8�A0�AD��pU:;),6�@"�6��AA���1��Gd[��:�|5��U*蟕�1@8����.�>҈&�_ɵO�0�.�%0P�	 XEF	 �P`�B.�:~T~��� �P੷����� ?��j~I����LL6��lOȝ������3":@U���Dv�|���ē��ç�'��"����(��>8*���cZ�uU�
h>$Q1$ � A�ɱQ� *tx��Q1	&*��pX
��~`"?�z*A�d&�H���;P�+u������D>/Q^(����@b|�u^!@pC�@z�zt?����$"��a���
/D 4�J H�+��	"��$���H��F"� ,���ƸW�+�M��� 8eEZt ���#�����:h�o㢀��:
 �X
��)�t:"��ވ�zh�0CB,  "��U�[ʂp^��R������M(�`~Cjr��_�? �D�P�b�H"E`@Lb��R*D��F{]�fnۭY@ l   .�8�[A����@  ��D�m�   		-�U�.��m>��aX�l0�P�UWdS�rM�Ō�u�6�n+�Xێ��)1���"�5���W��l����^���5�#��L��+���:m�34eꪇq:G�p�g����m[9��m�r2�Wt��jD�˷l��Aj;k<V��rGY�T�{':{PVk�gH����q��:��9nUUnT8j�v�rp���CX�lc�8�rG�g�l:�Fnwubז9���uWuͻm� �.��t�|3��r�R��i-�7��^<B�*��i̓ъu��h��BD�mFVF�KEs�h}�#O&<�]���}>U3� �7+Ul)�s�;1�C�y�kH�v�sϣ��g��;s�ʹڄ�� ���9pk

p�R�Ǟ/b��%��E��H ���m�"�!h��͐r����h]Ӯ�L�T]�z9�fg���5\�@pr�ʲ�E�J��k�<<NE�Li�^�Mgf�
�k=�p"ם���CQev^!�<�����k�G�M�T��&�9��t�NӨ�M�9"�3�&���jN.a�S[`��.��.Iֲl�����=���1{s�V�v4(h�W�d�]Q�X;���a�pgp9�$9�m�'�ݫ�o,��!�ӗ����tkP�ۅ�5�yz�/e�CG4�G�Yc^�r���5�5��*� �ٹN�8�^�Ul�rś���@	��2��=8�ո�Ⱥ*m<f���"�넻x��SF��k��8ܩٔ퇍9��cv�V;��[r6�Eܼ$�I6�SM,f�v��#8u����nH$i"�d�H����qR�e�n�g��b�d�l\�J�@ɶ�kj,-\�	�Z��k����M҆:����Le�Τ�Vl��`�^�8�k<��ꧥ�MOE����Kr��L�^�덎�dz<j��K�)AΓ"�J��Xڑm�_��N*�ȍR#�Lٷ����z"
/T���M>B
.(�p��ffkZ֮�˳ؚ���&�.��dyg�%u�Q��.����q�j��-p�vt�ι͋��.^�7�.{Z�#�����2voQ�����{b|�
b:G�u]����j����[Bp��9RQgh�Tݓ�r��n׌�'��]!Ԙ$b���=���*�g�n���V��F��tp�NmWf�5�ۗ�ݡ'+��fQ�t]�&Y��Ip-rB�ݸ1���nɞx"���(�"p���s�G���9ͺ`�hؾ�_���~a�mq`c׭��j���L��ٞI/|�6-�,���w�t��F=h��(���3qҜT��M��� :��@zA�eB�V���`��L�ۦ����ߓ�]�X�ǫ\�Vƪ���{� M���JqR�6�����ƅP�U�j9y�ɺ}�2�����{]�Nٰ!r��;)���L�e�^f��r�)�Ht� m� ��&��ڮX��m��j��Ϟ���R67����E���~U�E�{x@z=����$/�����RՀ~��0�n�{�ICx�zl�j�23[f��UU��h�����$� =�`����q�Jۖ�e0rw^����l���?��������y{���]�����f,�Z˩�S#�YܺF��fQ�6�e�;kD�jI_�;�ŀ{�� �l��=0����+v��(�ݤ�l��ݎZ�����}�)3�C�­Q���;)�N}�znI��}۹x �����K~_�m_���� 7u�֪��L������b�8����;�	���X��c�`��ŀ{�� �l|� >�UU�|Pm�n�ۑ!6�ƈ�L�k�.�h�]I��=�r��C������p��::���c����}6�s)�H�p��c����)�w�t�&ξ��-�,�6�q>��ߨ�V܎ID_9���mW�t� =�`�?wPli�~ 5NK0j���?sn�}���¨G5�D�����z����~Q�V��B���6�w�t�8�ݘ5wq`�ڗ�E=a")Ȏ��A��y����8,�x�˃�}�"nk,�7i��P�[��'P��V��RI�����@u��N*@zd��$�7+r�V����_{� ��,��׀w�t�?.G�Z��vƏ�n[�rS����M� |�'�!x��F8V��KV���Ӟ���?w�� w�ۀsWw w���֝c����ݴ�@}��\s���*@zd���M�IPH��Z�6DK0)X�p��Jh��sZִkYDF[��U�vyќ��pR�]�']�)�gv��.�.؛�m�ѝ9�cT���[J�l�6vn�n'��P�dzm�#�?�[|)����sk�Z��]��6h`2�����n���˴��J�a��퀷.��[9�0�7s������>���|�[>�f�EI//Aŕ{^����$��l�d:�[�n�$`/4ˣ�΃�s��64�5���瑹vz��w�:���"K
��חF�ɓg]�a2�9��������K�� ��� ��,���Ծ��ͺ`�jz����R�&j��fڿ(�l�����\X{ݸ穽��JV�D)j�?nIh�`�sP)�HY^dj�U$��^�m� ;���9�����_?�w^ǽ�lV5U��'�� m�@t� =1�@>���5����0tjT� �p��hۧ+uYC�kb�������5�%8�r�n�X������g-�V��`g�Zt~`ow� ����1���
�R)j�?l��[��P��R P0S J%6��2�s5��^oM����WP�l3���:ayZh{���M��9����w^�����*�Ic�S�}��U�s�@?�|��Z�� t�8'-��$� ��,�_%ϔ��?�� >sPLʚY{ar��V[��s4��+�[�A������5spR���1TʉSqʅj�
!KV�ge�M� |�:S���0�ʅ8��9��sN�϶���l77���[ذ�;� ��u��U-����O�}�nI���ٹ@]	�P>N�~Q�?f�ܻ�s���'�k2êI]e�7-�9��� �����n��wn�ou�uؘ�UH�� ��- �l�5ҜT�;���;�]m���]>�3�����uȡ؊x�z�N��H�?�ww���8����{��=�`�9����9hv>��PVW%�IL �;�=��6g-�V�;��϶��P�}��r'5EYWff��S�HLr��� w�ۀ~z��=��+@(�-X�(�IO�{����\X}�V�l!$
���W�������͍��W�j�&f�m�M� |�:S����?>�mmVJ�+��TO�'�Qr�	�vn;�8�x��˨W�tv[i�zι��YW�� |�:S����M�Žv��e�7-�9���<������`~ή,>ͫcs\ۧR��+n��+7i�Z��5�]�XދF�i�**��xzEH�� :S��o�=����\�T����>�f�]�X��`gӺ����B	C�������HV�޸[KY�֫s�D�X\��1팩ؓnn�m�������\7]�&��ֱ[�#�X�0��,n�9�Vj5m�O^m��-��f0�Z^|�M"�K�M�T�/O<.$ֱ�0�Z�nzz��/\��\�Ц]�x0cN�\��]I<�Q��YMC�G\m[dSb�۾���Ĕ�J �s�+FKu�B6�M�J"��_�J%�����lvn�"ۆ�:����-�;h�B�w/]�"��[��v~{�W�;��gc�03��������Z�Ih�r��d��UZF5-X�M׀w�u��������~�4$�W�j��J�;�Ӻ��Nk��BI��j��'y���b�*��D�ܯ ���0JqR���K@:��^i��8�s4Xj͵`t}�|~r{���v�9�h��Z��kM��갭�1��j:�n�nM�ו쑢s�Pj֤裼��
��UH�� ���`��xyۧB��~a���X�o�
�
��sD�[����j��F?l�"���� �c�&�Ҡ�,�vS ��ҜT��w��t� 9D�����#��9��� ���`ٺ��L�S}C�@��
!Ki��2K@>{�"��_�\� /)�8;v1�Br�K�p��n��ˑ|��yla����˱kem���3/sO>Ͼ��@9R*���=� ���*B�l�&(�xyۦxg;����[o׺���m���o9�~�I��Fx#������K�������[o���3v��ʼ��s�ІDM��^ZW�1 ,�|F����]���3F�J��D�� �bg�M	!�����M�B�H�bGϊ�;���&=7�^�(�&�	�ȕ]l�����5	Tt|~ �89�C`�C�?4@Ā�Y��b���G�����	L$�3�L׷�2�˄�.��U����(. ���h*1�w�M�� ��j&���0��|����*p�aqpD���2�Ԋ^+�@���`���f�4�i9����B�Px��H�*����v* Ă��>_��X�@���+����(D%)S���_��}��̞�W�̷ћ�~u�[j��R���o�N��m�Ws����3k���B�J��w~_�6���`�hT������Ͷ������FfY�u���L��{�9m�^��<���ߒ�����ST�6�d�&����c����y��:1Ѯ��y����j�'u�TT̔��bQ2���V�o�BQ����[o׺���Nf"�f{�_�ל����F�����L�R�m����/߼�^����z��M��$������6ٛ\WBK��=t�M&�ҩ�R
��~��ȉ���6�o�-��|�fN�o����~_�6�v�$�U�]$��̸OͶ������3,��um��(�]�/�m�&��C�3!\يG��D�?���I��~����	Sv�ߛo�y��~m����.I}����q6����n��m������ʆ�N���&�v�s�n�z�W6{[�ݫ�k���nn!:(�T���GZH���}����~m�>�&6������m����m����?:ڭ�
�^�\��6�^���}}���m���3-���p�-��!�o�]3T�	e&6������m����z��m[���ͷ�ۤ��|��A����+������a���ܩ=^���[�b���6K����5��*���L�R�o�o�����m���m��mn�ߛl�+J��y�i~�-�$@r	@" ��������� �.om��[��1��̓��I��V�S�s�K�`��r�)�ݮ��g��7k���c�p-�;<�ͧ<n6���v%�T�Έ���Wv9��5Gk#CQ�w=q4sbܝ���o�{��t=h�յ�O9On��^vq�[1�8�-f�:���̹z�(������R�q����sF (�j�Bv�=����&n��뫳mr-�g\��U������|�]p�e�����Nx����a���rǶ���g����v]���O]�����Z�u������o�{����9ۥ��}���~m�v�$ګ��6I#��+���_�wvs�j���J��z�ﳷc��}��d��Z݉�;_�Ͷ���v�o>տ��亮�����uo?ߛm����-�H��m��V�_�6�'nǍ�����~m��ݯm������m�V���W�ͷ���cm����f������m��V�_�6ޭ Փj^�v.��q��q��֓zڐ�'���@k#d2ݳ��z��njw������6��+i�m��V�]	D%}-���m���C�J:�+����o��^�|9B�y]+���[����9m�����6�^~��羅�?'�%U�ډ��^6���{�����;�m�ͽ���m�v�x�o�S}C�@�*
*ի��w}�,����/޲�[��]���S��1�2ͪ���b�Gm�6��������۷E��ϵo���m��ܖ6�B����Q�[B�A@��5��E^��&�=���z�_,�T�"N4�eʌ�nu��Q����;�b��o�տ��ͷ���1��6�_�Ͷ-;`hW)U��GmWn�J��z��ۊ�]��Mr�뻳�U���߹�s��P�U-V�ߛo���cv���ݼ冻�"ȑ`mz!�R���?b��o�5o���m����4j�J�[T��${{����9���l}���~m���Cm��}�

�ӮB�_�Ͷ��������^��o^���|��~?���������E�"���ڹ�%�nJ�l��a�r�;���0��m�%���o�տ��ͷ���cm�m�ߛm�w)��ޮ���U��(�V�ߛo����/��ͽ���m���q��y�/ߛo��ٵV�����T�ww�\�z���j���ҧ�޻�v�M��5��b���n������9����oߺw�9m�_�ٛ������8}�s9���m�N�ʭ�H��wv�T�{�wn������/޻�:E�����yt@o��J�tu�K�yʎJ��u�	G[RtWg�n
D8h6[�(��V���W8�{6�<m�ͽ���m�n�1��y�/ߛo`�63�D)e�m�ou���o��Lm��j�����������W����R؝r��~m��Eww~�'�޻�x�e���r���槮%�j&K*��o�������Ǖ��m����6����oV<�P�EA
ӵ~��}}�Lm����_߭�}�l���{Ü��"/b�?s��~ ��+gM�S�L馷9z|.R�j����,��9���J;L����kX]��t��:�8S;<p]9�;�s�u���gb�l]Yݱ����k�� �4j�Ǯ�)�W#А��ŵJ�%Z��T��Pv�n�$��n�Ͱ�ons�,�:n����t�t���Π�����돆����S��gd؝��:]V5ي^�.R-����qt���ww��{��ޗ�/�s�'9jV8(��Ӓ�R���':+9�{zf��ݻ#�Y�)sZzs��k��Y2�Ge'���}���m���q���[���_s���o����5��X�t,n������9��璒7�/{�������1��{{������4�ʤ(}#�����J���]ݻ{Wwv�P���ΑV��o^�ۜ��մɪh�֎r��C;��&�m�u���m�nګm���/ߛoX�63�D)e&6���i��m���q������������cm����s�Ӱ�v��[�V�����E���{Q����	�g$X2���OZ^�16�� ��H���ʞ�z����b���mC޻�i�S�%U��N���o�uo���D_��u4bX��"�P��(�qb:0�r�^&6���<~��|��m��q�=j�T((K�������cm�w�����/����m�|��~��|�ͪ�K#��{�b���mC޻��ww~r���m���&6���f�buФu�'%?~m���[��|�!B�yw��o�m�����:�]��`�"�m�������Q��T��sW1�v˧;�Lm�`;-��v��ͬ�C�y��TT���1�����jf�\�V�mB�K� ��6o�BI&�ݮ,�k��j�V�h�:٨�X������ ����ܢ�ċ�R�� +�Y������0�{����D�^�7�@yʊ��� 9�����qV�m����`��q`���o`��{���0!�[f��:��Z�7Re��+u���O�<�Y���q ��R��:��T�)V�������JqR�������e�y����|�	]�o`�� ?>�f��c�:�X݉��L�^��N*@zۘ�|����mn����������dܐC�{��t%[���CjV �!�I��7$�g�v橫v�����7i�nb�� <���Ww p�u��r�w�7������nf��ts�]�gv�o��<n'h�j�&���]�FfnU�Y���|�7�@zS��Ͻـn���Q���Er�`�+K�K�B�3˽j����3�/��$���#�"�Ս���L�[�V癳g(�M�mq`}�\X���֨%PR	%�T�<�#Т�wzlޯ������!Nyw�V�}��Զ2\˩��3�,DG�Fw{���޵`~y�6��	R�"J��~_���0�D����@H�@�!� �"D!! �HHBaa
�a�I�6�"�sX}��6���C���O�񮛖���n�o����P6�ک�u��#@�B�cD9 pc+Z�U(HB.�'?��Ő]m�T�1�q�)�bRH���h��) �ml�!A�0��F+�F'����bq����	�DHF/$��$�<B�2�$�I"�{��@lSG��4��,�	8��a5.M��?���=��A�$!`F"T�@���O�����F1"�"!B0�{6�ݐ�v���_��j�     .�8j@m�-�H  �-�     t�;Kv��L���L7�r��̒җ��c��b{j���m�f��pW 5�)P�-�8�M��IL�#l��fP�MJJ��)�x�^�k��W�D�h:�ԭ�=�k��@j���(4V��٩�u[�C���"�����[�݆A�-�9M�!�R�p$8�r��uưlv�A�dUDD��i�Nfe^x*�����`v��s�u����ak��:skpf06��j�UU�U�T������n����Ye���L��ʼ�g�֢Av�UQ�X�G���J��rI.�Y��m���-��dq��Ёs�w=�Y���y��m�:.�<�9i�λ5Ω��8#[C[dY��3�dv6�Ŗ��pSs9j�ͶA�n�Ζ�e�� �;$`��:E��Zʩ1
�:v��ڕ����
�)��J�f����Z�v�sۣh�`�^����{qWm+۞Ӭ^;X�l';0�n�)�b�c����琑�3���.8j�%��W;p6�M����ew�骪���h7Y$n��<cIE���բ��z3-Xx����y^r{����[Y�0gxAdv�9݊x�gm$�rU�F���u�Yq��,��v:8�cNd5�Q��ｻ}�v^Ů�1q�H�w����ᷚא���)�ݨ��5�i�zׄ�E���mʰ�3���@h��ݘ�#�����Z&ivx:C�-W;�8����������m\�ڡ���o<��6�ӵ�e�ٱ �����N!��b����;%ֱ��hz�L��r�mn{�\�̪8j���My&��d�lJ�Ns�y�	�0>���MR�Cg�!*E�t�̭!5*����J�j>��؇�UP��T��-Ǝ�v��ڹ��8��(��kv���j܍î�{B�qS�<��gؘ�bd�Cs'	~����[̽�\����e��:�����4\3WFf�d՚5�^�����G6&��!��q>x��� ��� �^*E�N�g5�.�wK(,��v�n�����N�ݳ���-��7g�k��qfv�#�
,�a�h��Z��MnO/X�!����q�h;u��?��>���!�\����M���An����	͡���.�n��	v�Ǫ���Ҵ�ɛD�mmZ��9p�z���Y�N�,�<㶭���Z:P��+��v�N�z�2c&+���M��FM�ۧ��w~s��{��W۷����-{:�x���r)����ƲN� E��r����O�~J�i�*�4��*@zS���� =� -9�ʥT>�v��ո�[s����#��u�{wjJj�ʪV��Vە���	$���k ��{�Z6u�j$�&�d� ��I J��nj��\����W ��wq`�{���������0t@n�9�i�D��0��)���Fs=�,v��o/Q�J$�]L�7�]�K-�yr����e_���{ w3j��r������j�9gJ5A*�D�5�3F��b^���Ӑ�� ��i(
�HD��"� 7L���'���6��bX�'��p�r%�bX��Ǹm9�W*dK����Q5-��%:��_�L��L�����ӑ,K���{�ӑ,K���=�iȖ%�b^���ӑ,Kļ��BV[d���L�~>L�3�ϗ�{�6��bX�'~��ND�,K������bX�̉��s�m9Ĳ!5�􇂪iMP����p��	�bw���Kı/{�kiȖ%�b}���iȖ%�b~���iȖ%>L�>��4@t�II�Ƥ�JF4��=nОn�i������*-e�yK�l�yf�%u�Z�kFӑ,KĽ�}��"X�%����M�"X�%��������L�bX������Kı?�9�y3R�&�j��!2!}ۿM�"X�%�����"X�%�߽��iȖ%�b^���ӑ?�#�2)���߇5"b�M�GSE��Bd&%������"X�%�߽��iȖ5���T���I"\�����K��=���~!2!2ӈ}=#��jKr�WY��"X�(�DȞ����m9ı,K�{�[ND�,K���M�"X�B�����q	�>���)�S%+P�BY��
�
A9ߵٴ�Kı?{��ӑ,K��;���~!2!2���<K�qe� m�2�ufs�h�!;�4ۺ-r櫱�������2!X�dp�۟/�ɉbX����m9ı,O�����Kı=��p��bX�'{���9�&|��|��H�Ydq��L�~>V%�b~��ͧ ؖ%��v��ӑ,K��u�]�"X�%����M� &Bd&Bxf�pUM)�7Up��K���}�iȖ%�bw��ӑ,���ߦӑ,K���{�ND�,K�Ov\�Y��CZ5u�Z6��bY���Ȟ���v��bX�'����Kı?{��ӑ,K��"�F��਑E]������ӑ,K�����-�l<L����j�9ı,O���m9ı,������bX�'���ND�,K��}v��bX�%����_O�^�)1�3\�<�C���u��.�ԏE*�)[l�w�a��Dv�����Kı/�{��r%�bX��o�m9ı,N�]��r%�bX�{��ϗ��ϓ>L�>u6��K`Pn:��9ı,O{��6���r&D�=�{��9ı,N�{�iȖ%�b���W�	��	��,�C�B&�R�Z��iȖ%�bw��ӑ,K���ߦӑ,Ŀ��kiȖ%�b{ݾ��Kı>��ˬ�i�5.�v��bX�'���6��bX�'�{~�ND�,K����"X���뾻ND�,K�����h�u%�ՙas56��bX�'�{~�ND�,K������m?D�,K�׿�ӑ,K����ӑ,K��&�!AQȅBB�}����ꪪ����V����qQ�
��2���HZ���3����̫l�]q��.��2���)6⤎0y�����m���s-�=�6^������R��V��
�XV��iZ�j�P=��/;m�ܶ�Sj%�Y:鈻�5i�92��c�}����9	��c�7Uls������%��6Nݪ6.U'F�ݭ���t���IlִK�V.��&����u!����x�t#��������:[�۝�v!��]����&�����h��ܦ|�%�b����ͧ"X�%��뾻ND�,K�k��D�,K���M�"X�%��'�,ɖ{2P֍]ff�ӑ,K��u�]�!���,N�k��iȖ%�b}�����Kı=��=v��bX�'��=m�l<K��SSY���Kı>����Kı?{���r%�6%��k���r%�bX�9�7�	��	��ݷ��S��s2�j�9İ�>�w��Kı=�w=�ND�,K����ND�,�k��ND�,K�����&�]K.f��Z�ND�,K��sٴ�Kİ�Tb�w��6��X�%���{��9ı,O���m9ı,O�t��7�W\�Bw�?|�pDnܾxn=`g[Ҽ׆�yp�H����~{ܜ�c��m�흵��f��Kı=���ͧ"X�%����]�"X�%����M�Ȗ%�b��g��~!2!2�`=�B�u2ř���ͧ"X�%����M�!�|@	:��AvD�,O~��6��bX�'��g�iȖ%�bw=�fӑ?��L�b_������r�K5�2��jm9ı,Oo�m9ı,O{]�fӑ,ı;���iȖ%��;o�����L��O�vC��SJkP�KsSiȖ%�X����ͧ"X�%�����ND�,K�w~�ND�,�HD���?�ӑ,K��2zRIg�F�R�Nf��~!2!2�wM�"X�%���{��i�%�bX������r%�bX����ͧ"X�%����x��:
I�u_�ӒPQ5>a�O�s�^7[R�3�kB6C-�{َ��v�v���m9ı,O���6��bX�'}��m9ı,Ow]�f�9ı,N���r%�bX����e�5uI��5����Kı;�o�i�*0Eș�����ٴ�Kı=���ٴ�Kı>����r�bX�%��o�I*�)�f��Qp��	����=�ND�,K��{6��c�T�� $@6 o�*w�*��j'���v��bX�'���m9ı,��Y����@�*jjn�!2" K��{6��bX�'�k޻ND�,K���6��bX@�����_�L��L����(TK�
\���m9ı,O�׽v��bX������Kı?w]�fӑ,K��{�ͧ"X�%���s)�33P��s�M<t�QGX1��ڽ��v�w#�6.X����2�f;	p�Z>�~oq��K���6��bX�'����r%�bX��{ٰD�,K���M�"X�Bd'�!�۪�j�D���	�X�'����rX�%�����ND�,K���]�"X�%��{~�NAL�3�ϗ��FzA��r��~ı,N���r%�bX�}�z�9�,K���6��bX�'�����~!2!2e5ͷ-�sBj�����K��>�^��r%�bX�����Kı?g���ӑ,K� ����xdMk��m9ı,O��&jH��4S��uN�~!2!2�o�iȖ%�b~ϯ���"X�%�����ND�,K��]�"X�%�����~��߷�wnW���5��V��{&m����Jn��^��w.���Y�3��Eή43Yu�N'�%�b}�����r%�bX��{ٴ�Kı>�^��r%�bX�����Kı/����i�P���.\ֶ��bX�'s��m9ı,O�׽v��bX�'}��m9ı,O������O�L��,K�R��
�t�K�&jn�!2!n׼��,K�ｿM�"X�%��>�����bX�'s��m9ı,K���fkY3T�.��ff�v��bX�'}��m9ı,O������Kı;���iȖ%�b}����Kı/���M��&j����~!2!2ӏ��D�,K��{6��bX�'�k޻ND�,K���6��bX�&�C��}����rn��7U�,ݩ�r�݁�Zn�K�*����4�th�f�3�<���ݯf�^ns���
ke4���:���#dۗJ�իE��O7f�å
ua��3��/2[�h���Rq�yu�,�yy�q�4�N����q˴�-h䣆R��,p�@̶nwC����X�I�T\�Ool;q�u-!R�;���%	t$�ì��MO�{��{�������W;d�V 	�M����a�5\a�e��e��n\��T��u��g2$��5-�k�9ı,O��}�ND�,K��]�"X�%��{~�ND�,K�}}�m9ı,Od=�̹l����)�k5�ND�,KｿM�"X�%��{~�ND�,K�}}�m9ı,N���r%�bX�{۾������&�f�Y���Kı;�o�iȖ%�b~ϯ���"X�%�����ND�,KｿM�"X�%�{�m��d֋5I���֦ӑ,K���_{[ND�,K��{6��bX�'�k޻ND�,�fD���?�ӑ,KĽ=��zf�:H$���_�L��L���Ӵ�Kı?g���r%�bX�����Kı>���[ND�,K�����"��m�
*�5������6��u��y}��r̻-�Yzs�.;a��d��fk8��X�%��fӑ,K�ｿM�"X�%��v����%�bX�=�7�	��	��f�ʪ�SC�I˖�5�ND�,K���6��	�!�"� "�b�J�/jȣ�b0
�V���"XD����bX�����m9ı,Og���iȖ%�b}�{ٴ�Qı/�vC��UD�A74\/�&Bd&B�>����Kı;���iȖ?���;�]�"X�%�����M�"X�%�����0�d�0�I�ֶ��bX�'s��m9ı,O�׽v��bX�'}��m9İDK�{�ڿ&|��g��^�$"<r��l��,K���{�iȖ%�bw�ߦӑ,K��'�����bX�'s���~!2!2��$��%�9a�z�*u-2b�M������Wpj��H���:�9���L}���F>�~oq���bw�ߦӑ,K��'�����bX�'s��l?���ı;�]��!2!t�����2�&j\�;�Ȗ%�b}��{[ND�,K���6��bX�'�k޻ND�,K��}v���*DșĽ=��fj�R%�Z�ӑ,K��{�6��bX�'�k޻ND��WGɶ��6_��%�$`@���"�Ҽ�h������ ��Z4$���H�e �R9����<�W� ��p�Ա��������8�0R�:��JB�N+�["D��F���aI.�i�
@��A��IE��s�~4<�c8Q������@^a@��u?:u��H�(JH��+�h!PpC`�i�E]��<M�U`�#��@? ��h`� 1π�@z�"S4b�E�C����߮ӑ,K��N���r%�bX���(TK�
Z�&jn�!2!��+޻ND�,K��}v��bX�'�>����Kı;��iȖ%�b^�%��Z!*���^|�&|��g�}���9ı,O�}�kiȖ%�bw=�fӑ,K���{�iȖ%�b}:|y���,����Q�T5�a�m���Z�S�iR,e�rV���v-����v�W:֩K���~�bX�'}����r%�bX��wٴ�Kı?{^��r%�bX�����Kı>2��&̒��nk6��bX�'s��m9ı,O�׽v��bX�'}���9ı,O���fӑı=���3&�KsP����m9ı,O�׽v��bX�'}���9��`�L�����m9ı,Og���iȖ%�bw���\�a�WT���.j�9ı��}v��bX�'���iȖ%�bw=�fӑ,K���2����ӑ	��	�s$�L����3N�~ �,K���ٴ�KİN���r%�bX���z�9ı,N�]��p��L��^I%��d�t�J�fGI�v�v�:�oNo+���N	I�z�\g�;�+a��tE
�v��p�3�ϓ�����m9ı,O�׽v��bX�'}����,K�����m9ı,Jt���jeՐ�f�f�iȖ%�b~����Kı;�w�iȖ%�b}�^�6��bX�'s��m9
|��g����-u:�#�F;%y��|�K���]�"X�%��u{��r%���bw=�fӑ,K���{�i���L��]8wHU2�L�A9�w�K��"��;��fӑ,K��{�6��bX�'�{~�ND�,K��}v��bX�'�!��2a}�P�5m�fӑ,K��{�ͧ"X�%��)�����~�bX�'�����Kı?}��fӑ,K��]1�`���P����9�֪�A��Uu(�a��K]�FQ��x����Ǐ�}o�	o;�КU���זu�̓�ٗggf\���\��i3�3:죸��UǅM�+-��n�"&�:s����:��b�m�xBͳ�-�� �ُi��ː�kOY�`^��y�Z�7k�r�f�B��4�[^UC�D�Z��5 e3z�)6^�f�8u�n�R՛M��@��߻���������~E�a�zo�]��%n]�.�n���۳M��+�n��k�y!��{�ݬ����[��ֵ�ͧ�%�b~����m9ı,N�]��r%�bX�����iȖ%�bw=�fӑ,K�����\�fM]Rj�k5��ND�,K��}v��bX�'�}��r%�bX��wٴ�Kı>����r"�bX�����UI��3R�i�/�&Bd&B�)��iȖ%�bw=�fӑ,DK���o�iȖ%�bw��ӑ,K�|]�z:���]�ٟ/�ɟ&|����}�ND�,KｿM�"X�%��k��ND�,D,O�j�ٴ�K�3�֠��!R:�F�$�>_��>LKｿM�"X�%�����Kı?}��fӑ,K��{�ͧ"X�|����y��Ur�턧�-�Cs����zg�%v���S&�b��ͧ�r��릖��A$Җɚ�.�!2!oV�_��,K�ھ�m9ı,N���<�bX�'�{~�ND�,K����Me��.i�K���r%�bX�����i�P1@���uHEP�@G�M��Ȗ&g���iȖ%�bw���M�"X�%��k��ND�,K���d��	#�j�ֶ��bX�'s��m9ı,O���6��`ؖ'}���9ı,O�O{�ND�,K�{}m���P��Y�/�ɟ&	#�X�}�i7�N�;�$D����7�}���6��bX�'����955uI����jm9ı,N�]��r%�bX����6��bX�'s��m9ı,O���6��bX�'�$��%{~wv� Z\�''9��N�,{Mxz�;�A��}�<�q��߃�ؾ�Ż,�{���%�bw���6��bX�'s��m9ı,O���6�"X�%��k��ND�,K�~�OeԗP�$5�35��Kı;��iȖ%�b}����Kı;�w�iȖ%�b}��si�(d&Bd&�oJ邖������,K���o�iȖ%�bw��ӑ,f�1]����ba�t�S�?��5��ٴ�Kı=����/�&Bd&By��抢�4�c��]�"X�%��k��ND�,K���fӑ,K��{�ͧ"X�*؟�����Bd&Bd.���,�I�C�kWiȖ%�bw>;��r%�bX��=�fӑ,K���w�iȖ%�d-��w�	��	����ET�Nk�s�.�xR�[��'1���T�n�3�Q�u�:(�L���;�v���ߛ�ou�bw=�fӑ,K���w�iȖ%�bw����@b(���,K��ޛ����L��^���J@�74��Z�fӑ,K���w�iȈ	bX�'}���9ı,N��}�ND�,K���6��bX�'����955uM[��֮ӑ,K���]�"X�%����iȖ "X�'s��m9ı,O��}v��bX�%����{!�7P��˙���K�� �D��{�6��bX�'���ٴ�Kı?{]��r%�`yd$RA$x�\����]�"X�%�z��=,C��d�ٟ/�ɟ&|������r%�bX'�w~�ND�,K��}v��bX�'s��fӑ,K��W�X���9T�Ѷ�
�MUVI��KcM�q�m�;y��49w��{޺���{Y�D2�����r%�bX����m9ı,Og��m9ı,N�ݞͧ"X�%���}�ND�,K���35u���&�ꪋ����L��]9�7�Pr&D�=���ͧ"X�%�����m9ı,O���6���bX�9Ϥn�N��L����_�L��L���g�iȖ%�b{;�fӑ,K���o�iȖ%�b{>��iȖ%�b~2��2�钆d%Ѭ�r%�`����}�ND�,K���M�"X�%����ͧ"X�؝���m9�gɟ.���]P
��Bv�f|�&|�	���.�!2��o�7��bX��x�ͧ"X�%���}�ND�,KS߄h!�Ѓ�P�\ A &gm��kU]K	*�Z�κX��Zo;dN���YNd;q�ld�i�[q�S�筆@�dN-X�f�
�:�v�L\�ɢˣ.\����Nv�t�*�\��y�R�@�M&|�B]9�犤f�{=���ɭ�bp@p��t>��H"���eĳG=��#ƋZ4E��:��N9���[F���V�����m�0�W��E�#nTڎ*��JO���;u�88V��OM; 3��L�<�n�������(�+n�W~���>�|��Dv�f�ӑ,K��{�ٴ�Kı;����r%�bX���ٴ�Kı?w_�	��	������*�Љ��fӑ,K��w��i��ș���{�6��bX�'�����ND�,K����N@lK���۞�h���$5��5�ND�,K���6��bX�'�{~�ND�,K����ND�,K�ޞͧ"X�%�O}�ML�D2�����r%�b�'�{~�ND�,K����ND�,K�ޞͧ"X�� Eȟ����iȖ%�b_w��J�
�r���i�/�ɟ&|���｛ND�,K�ޞͧ"X�%���}�ND�,K���M�"X�%�㿿��ǋnQ��e��7Y�nwa�>�n�=`;��9��m]�܄ge�����)��p��5���Kı;����r%�bX��wٴ�Kı?{���"#�L�bX��׿�ӑ,K���{�̙e��(fB]ͧ"X�%���}�NC��"#ڋ�Ӹ�%��s~�ND�,K���]�"X�%���OfӐ_3�ϓ>^����@*�	�e���ı,O���6��bX�'}���9��HdL������r%�bX���zn�!2!ou��5IN��幩��r%�`�'}���9ı,N�z{6��bX�'s��m9ı���M�"X�%��k���3M�R��k5��ND�,K���fӑ,K��#�{�6��X�%�����M�"X�%��k��ND�,K��=m���̎�:�N!5�N��/��X#�I���Y�N�v�l�������8ۥk?{�7��bX��wٴ�Kı>����Kı;�w�iȖ%�bw;�L�r%�bX��'�����S535�ND�,K�{~�ND,K���]�"X�%���}3iȖ%�bw=�fӂI3�ϓ>Ow}$���Mʆ�m�'"X�%��k��ND�,K���fӑ,t�؂� H�/��Qw�D�L�oٴ�Kı?{���r%�bX�Ͻ��n���sMr\֮ӑ,K,K�ޞ�ӑ,K��{�ͧ"X�%�߽�M�"X��2'����p��	�����%��2ҙTk[ND�,K���6��bX�(w���Kı;�w�iȖ%�b_�������L��\���*�Lj���Z��n���[]��=e�:�+��3X`�R��ľ_"��m�B�nT'm�g���gŉb}���ӑ,K���]�"X�%�{���r%�bX��wٴ�K!2!vm���IN���j���Bq,K��}v���TL��,K������"X�%�����m9ı,N����Kı/~/�$�k0�3Z�f�ӑ,KĿ�{��r%�bX��wٴ�K�,N����Kı;�w�iȖ%�by�3��.�l�CV��kiȖ%� 6's��m9ı,N����Kı;�w�iȖ%��Ɛ��� ��?����>�3<w��r%�bX��'��5�h�S535�ND�,K��m9ı,?�`"������ı,K����m9ı,N���r%�bX������;Of;v�s�M<qZ�#�0�krݍݴ7��͂�T�s��G��n�1s56��bX�'}���9ı,K�|{[ND�,K���6*�Ȗ%�b}�o�iȖ%�b{>��-�WE�5�sZ�ND�,K���Ӑ�R"�dL�b{?���ND�,K�����r%�bX�����O�2�D�?�������J%Ӫ������L��]���ͧ"X�%����M�"X���bw��ӑ,K��{��m9ıL�z���X��nT+e�>_��>L�D��;�����Kı?�����Kı=��{[ND�,���6��&Bd&B��}34�&�j��:�.D�,K������bX�'���kiȖ%�b{=�fӑ,K���ߦӑ,K��u��df�׀@�)����l�4��R�??��bB� o@�jy�P��b�,y��L%�I�41�`��9)H��F�M������6|�2'ˎ��܉	p��	e4	��B o[%	��
��l'�O�Y�:ǑJN��"�?)���Ҵ�Cn��� ��     @[R�	 �  :�8��    !�H��Q]m���&8�</HmU&�"��K�&vWT:�[��\84F6�0q���m�SWN4��,n�nع��uD��U.x)%�5�����V�e�))<��Z��Md��b,5��t�o%��9'6�n�۲���<F��m��Y˨Ѝ��R�&�6�l�#;e u`���k�ˎ�Y�͠�[��)vU�I����E��m�۶���M��i�p�mx��]�<n9�T����U@UҲ�U'ny����0�-i����B��\3�*guZl;��m�bۤv�#�$�I"'\A�[�։/m������toi��nnw3ܭ�6��ۮ���"tSE�\�ڝ���	�mSJe6�.�5=.̵ڹ-���iY���p7Ogf�lL��P�aQ��Y�e@]<t�x�!J��-�����5����J+�j0�� ����\p�
�t3�hܔ�Q�l���r8;u�z6��p��Ml[=fN��N�w �J{Wsu�e�fL���b�*���gs�Q�(���0�Z���څ��Ur�xkQ�u�Np����Q����uiQ�BK��v�!΁\�i�l�k�f0;-�K�v��]�c�����fv��S���,�e��q��痀.��[��]{�6�\�kgT���nJ1�����@؞��UJb�PS��]�1]l���]]M�A+���Q�vvW�q�-d�in�UyVy\�.�9���HF�F 횛���[�@���-�]�����n�z7�.�mج��funq���gp4�%��i2��6�bu�UJKJ.۔�hϴN�f��v�!��r��ܒK�UJ�ɂN�*Qa������-W, ��d�k=��<�����:0tp��3��Z��іi�8��nYR.Z�&z��
 �� ��٨+���Ԃ��nh�����H.��ϗ��LD�� 	�A�)ӫ���D�t àl@�&���ꈿ��V�Zֵ�kZ���3��O=�	�\�{+���n��x9Qf5�ru�\Q����Ng=I�����Iu"�*4Ug�����{&m��ۣ��s�ݒ':���$y�rZ�����ۢ�"A.h��ukaW������j�]�1�vkQ}�h),f�݁nN��!�= ƎP4N����Nr�0jp�9"��]�y�ޮ��khLssv��>WN���*Vk��믮po<�ܜ���BF{�d������������^��U�z��nL�����������,�_{�7���%���s��r%�bX��wٴ�Kı>����,Kľ�}��"X�%��>���a�DԶCZ˙�m9ı,Og���r%�bX�{���r%�bX��ﵴ�Kı=��{[NEı)���$���)�ֳ5�ND�,K�{~�ND�,K������bX�'���kiȖ%�b{=�f��	��	��wt̕J�4��6'3E�Ȗ%��%���m9ı,Og���ӑ,K��{�ͧ"X� '����~!2!2NwUT��)�uC���k[ND�,K��g���Kı=��iȖ%�b}�o�iȖ%�b^��_�L��L�˄��3L*P�[pm�3�0�O����
D�����r.:��4.�j7&�.���2��Z�r%�bX��wٴ�Kı>���Kı/��kiȖ%�b{;�����bY�g�a�<�2�nT+e�>_��>N%��}�M�!���Q����Q�_߁�%�b^k���r%�bX�g�����"X�%���}�ND�2�D�>}B�)�nX�h�_�L��L����m9ı,Og}��ӑ,Vı=��iȖ%�b}�o�iȖ%�b^�?H�+S$��,�[�/�ɟ&!(|������ӑ,K����fӑ,K���ߦӑ,K�/��kiȖ%�by�v���ˣT�CZ��ֶ��bX�'���m9ı, >���Kı=�w�iȖ%�b{;�����bX�'�=����u���tj榊\ԍ�u���l��u�x�MD�[�����|���gmg��kY�ͧ"X�%��}�M�"X�%��k��ND�,K�w�͇��RBd&B���7�	��	���c��)�:�nX�����~��9=��oM�����B��9��4�t�:�ķ5N����l{�6dD+�DDBVT?�A��a�LA��,*��(�
?BH��,��v��&{*\J%�sU6	B�O���=ޯ��S�ٰ1�����aHni
�j�������
uo?�r{�0{ݘ���$��v�` c�*u.�#���y�̽c��!�-,d�1�H�&	o��R�[�vS ݝ׀j}ݘ�͞���~a��ŀn.��̚L�#s4ꦝ�����(Q�9����\X�����g���'�Q�Z�IfϷ������DDB���y���M�-B9݀R'SQ�d� ��� ݟv�I������C"(r�b��E��TF��B��zB���ޫ �y�_QM��Srʽ�1�@J�& �j9�@z��6�t�Դ:ƦiR��3�44��ډ!N�x��ثõh�n�����w��$:�v��d������`9ݸ�n��m� ߖ�tcأ�":��`>ͫ�(�Q
d�z�X�����`|���m��Cr�G-��n����ΈI&�=� �ޫ�׎v"h����/sD�� %9 �j���$����ȽIS#�rUe�)ȩ >sP͂���T��;���ws��� %�6Yv�.*��1��r�p�K�{b��f�]�I٤�l�]-��|���\����L˳�U.����"R�)s�9����n��yG�j��n2�p���t�۫4�6iг��:p��-�^��)	.L����jϙ;�ۮ���6V�#J�a^�tZ�K����wY����f	@�{F�p��`g��^���6�v.�=[r�x������O(����d�f�Ytf.�4ac��b���r�3���O�݃uŷg�'��9��s�@�ȭ�V��jn�����7�t�3��^�
<�!B_Hyw�j� {ސ(��j[��skK�D$ٹ�j��֬�ͫ伔$�d;�b��6�9�nX�Mo�j�՛��؆�͚sn�9�`�q��*_/�I���R O�� H�?T�wV\�?�#�YV s{� �I|������ذ]�ŀou���Ȝ�����9M	՝d���u��"�8�:���բ��T�my�V^n�9�@>�RS�W�Т#�}ޫ�9�*D�MSr�U�rO�w�6�1P���-�>�vX}�V�֗伔(�j:eyTҒ\���TҰ<�޵`nmX�ZX��,S���Elti�+Sv�$��ޫ���>ݵ`j��V � n�R�I�j[��skK�B�����[�b�ov�| յW*n�6�svMɌ۶�1�v͡��ڏM�qD{[Fm<�]�	q�-b�����X���;��X�ݵ`nmt%�0�����:��R�u;F�v�Wwqg�I��� ��q`g۶��P�
"��^S�1�T��K�54�}ޫskK?+DD/"!/õV���� ���o{7$�~�`g4�m��M�P������$�w_�u�nڰ�o;z��=sЩE5M�n��>ݵ`yDDDj��W���@t��P3�Ue]_j���'r�(�N�x����z�7ZF�������]��$��*�pnJU�[�b��6��kODDB����u�c�\��m�4���V s{�?ϒ�6w޾0��V,ݵ|�/BP���X!{ސ6�5-KuU`o�^,�vՁ�n��ov��I�c��A;)��!C����ӺՀ}��a��$B;P�D��<��1"��>_#���0��v']NѱE]� ߱��(�y���ͮ,�vՀp�E�-���2(�e��'%�,��8Š^rj��bY���������y<�^� �j���U�U~�����ذ��<�0��M�n�ei`g۶��ڰ�6��D%I%2y��>�U*j��:�,�zՁ�ȩ tsP� z̩[�Xe���M+J!�iߕ�goU���ia�P��w�`tt랙UR�`ةUJ�>�ڰ9DDDz"��x��zՁ���ܓ�P���B �D�����O���U���suv��e�w��ݞ3m`Ѷ����8�p,py�VfӞ��^���+�����i�q����ۡ�{c�l���9g�\�C�rݸ��dp[L/#!�b0���q"0=��`�d9ܖ�8&'eȯ���h�;l�{p6��){.2����/J��9�k��vqu��<-��.���<�c<�k�p\B��ߞ�{�����׺�ߛo��6È���N�ͦ�͸�9�p��W�z�z��v��&.9�U_�����ϷmX�m�DG�v��;�)=F1�h���y��?�Bl��v�;z�ە��M���r']NѱE]� �o�, ��n�{t�;��X��Au��G�J� tsP�`�}"�UW�O�Ԁ�;���c
�ʄܶ���L��T�q�T�:9�͔r���QVt��ڮ8y�\n�cGm>�v���*��6���R舁ӧ6���T�d������Vnk�`nmz~a�mq`pl��eP��Bʰ�u��}�}����M:
������]I���ܓﻯM�g۶���6tt랙R�P�lT���`��`}�ZY�&�;�X�u� �|-�Q��h�nۀs{t�;��Vnj�ДB�%
g}ޫ ��ϨC������ϷmX�	F��z� ��j�� :��,���fo
�;]H⸮��ݕ�n�X7ż6�����k!E'��%p��n��9F��ڿ�ӭXۛVە��IG��֬�%���:���U2�XۛW���7�^0o��,��q`g4�m�5P9P����>ܭ,�v՟Dd�$+�A ���[���A1cB4�"BJt>^pX�a5y�kA�4i�KM���4m$Id@HܻFD���6l~0��َ!hOK��C{H@�$?Tڦ�� Fa�B!�RP�!,��7�n���,��g�h	$"��zOيe>h4�B��H
�I�m1?F!!X�%H�$@`Ȓ$#�!R}�$_�� �D���I�sqH)a�ڟ�C�Q:����2F�>Sz�0�¨�O��`�"�0�$��N��l	����1�a� #��T>���H�~T��@ظ��Q"��P\���4��tE�L���CnO���, �wn�׮j�}j���vS�K�'���X�=j�>�ڰ>ܭ,��dZ����(YV�鸰D����}�j���#[b��k�����7�J}�M��`�לb��뵻��MA��9: �KBA)#�DZQF6���~ ��`}�ZX��D/�7��V���^���ц]���� =� �&, �;�<�M�;�'=B4;kt�D}7� 9Nj |�{q�h�T�9F����������}��>���܀D!$v�AN��ڪt߷�nnI�镓�+7?hiF�f� |�{��X�V��j������r��u�Aĝ�&y;unz��l4�ׇ��:U��-�{�)��m�5Q�&巀{����?ovA�@��[�y��~ݭ�,�:�,ە��M�q�V��U��ۦ/�hl�����-0˷��?fmY脓}�\Xn���#ج��1�]Nہ���|�7}p{o�����	7˷�� gr�Q�D ��n��˛������rI�ﻭ�<'�ER�R Q�s ?%���U<�$�V����l��S]q��a\f'e�G�;A�7r6��c��02�Jr��B�m����{����@2���]�m�]j8:�ǳ��v]�r���ݺ�.3z䬸����n2�Ν�Upb��:�z��2mn;�9<b�6���rQ�Wdې�;i1�N렶��c�=t�q��rXǮ�/�K:i4�m�x�A�t:4��ђٚ�ٙ�n�~x����32��:��󫒣�.�O�v�����P��f���`�T5Ɯ��w���1�~��X����M�幨�q��nѺR�Z��S ��v`yݫ3kKrw]�"��B���=%�w�K�PP��U6��������(P�~ݾ0�x��5��]���Q�UNf��=	D<޾,ݮ,��`�j�;٠Un�za�E�h�m�,IB�������������(����rgkzMtA�1 t\ah�=xɒxt�]����ɜ�K�L�G�V@u�S����6��	&� >�}���B��8uJ��?n�]%	~D �����x� ��﹮��7�|`ٯf t@s��),lD ���6��32���Bo:N����wX��`�v��'e0?�{�|��;��?n�Xy'���X��P�U�T����v�vlBO������ ���n�Wk�4�@H��Y�
���	܍�^��F�ǣ6:�h6]{�;��ʽ+C
��w�5 ۊ�����z��<�i�m�5TnUSrڀnEH���	1 N�W�vt5�T|����C��ݞ��9�^�	A�J�nfՁ�nڰ�"�e������<�g�z`�}p�vՇ���������I�*��.��曈75�EH	�%�:�$�<�܉{dNxe�AUJ��mq��N�.�ҍ�g�:JLlĸn�`y����ݶ���Kݷ�o���`ɺ�=�f o{� 7������A;j�7��w�ُ����>��W�Cft����ڔ�]� ���L ��j�Bo7�Ձ�=���zĞlʩ�	*�4�@��r*@N�-~��UU�ME?>�#b�~v|��%�D/�������ÝUT��KsJ�sUVٻj��(���}�M�nfՁ���$���:X9S��4��H*�_jIs^�wX䤉V,�*z#���x� �`��sA
dC�����v�tٰ���(_Ho���`�9�G�aex�1 F��RvIk�~�	�B�����3475 �����@G�v`������B7m�;��H	�%�:a& ��T�W���W#��y7^͆���v����
��D�%
,ǵUUUT��C<�U��l�&�9�l<�`$�X��㍐.5�������幺n��ͮ��`��9�09xmvLG^��sҁl�O�) ���b�`O`ulj�+zͺ�!�X�Lo.���mQ�qC�N��;�'�a���XhN��1��i��%0�b=�;�g
j��+��
�*�{n���J�\�eݤzmvn�V]X z���U���@�fL�-�!��&n{gi��_l��ob���\���a��o:[�v+[j�
�_@�徘��@7"����˿�9y[��0�̽�@���T���b��1��c�-���r�����{��n͞ID7�=ð��>���ۅ5MЦD9�V	��t���; ��n�{����r-RU	"�W,@;�@��G %���v���]�.��<��|�k=:]{!����r�lu،v!'���;��\|�սrc��<��j��H�� �1 0��B�����p��ş���BP�(j2�\�h��_�^w`��`t�ShV�l�F'-X��L���Y�Q
;;���{�X|N�R��j�K:�,:=�߼� ���`~��,{ۦ��k=�+~�Y*0~ݫ�����_���`}�Z� �}���e�����7C��&%���Rj��F��^x�]��&����n�3wPr*@F�x�Z �&�'M�W���q��V���<�l���x��� ���X�]r-R��rje��9����Vz�	}B#���T�`��$TҤ8�"��{6�X���Mof`�"�)���v��;���z��72��9ٺ< ��v!RX؈I%���i`rQ�.�~�����>�ڰ1�V�\������1���&zK�vt��3����獨�`�.ˣ���S
	��`g�ZXd��>�����l���ޤ�Z�V��N�`���}��`~��v}���(P��oQ�Z��%�:��v�X�w]�Q	$�����;����ǲ[bj��R���@y䖀}6y!h/ߕm�%"1�m�������?������g�Zݎ49)�w�t�9ٰ���@y͂�O�(�0��]n;7F�]r��&wa7J;X�zx��lvt�e��Z��r*��#��;O�wg�< �sj���Zz"��s�� ��7�?�Ҵ��st���@y͂��`��y/��D*GX"I����� M��HZ ���֭T*�������_'��x�;�� s���'��x�9龵���ݬ�*�4@s�@�j�l�w]��h��,C��@��mSg���~�b��1��k��:t�|�q �E?'��B��]?16�6p���`�#��+��7��y�A�@���RIM��N�����Q�r��z "�4��A]
�?Ц��Q�i�q�ƨ)��tO�,�22*H�C���8?p	����t�	R�Eh/�Q�@�~�����ȥ�(���YY7n�2L��Z%�      l��m�@$  	!     A:[I26��I�G�*�v�0��i]�	v�T�fR�Y����6�̡��شp���mMu���2��8���v�A୪�6],SI;;;6vV�#��WT�k(�YC���!m)�'k��A��n���A���m�"J�cu��B�(!��h�1܃Ed��ج���mZv@f��OM�3J5��s5<;F�U��� ���G]�e��t�w&�S�Sm���W�q��'�d�f�c��k,�k\�vlhvZ�j�XqJ9Gy��m�A�;CRѸ�m=vf켓Y��O��n�8��r6m�<Uf훨��ɼ�q9�.�����wE������\�4@��V^��h)���O��㴷�cz�;2ڧd�Y�2�:�v�$VA��[U��9�^�SH�A�=[�lgpu�q�
(pR�l�m&86�*uD�<�22��/CY8#��g����l+���8���6:���s�Ea�tƓ��pa�Z����J�U��W��.ڵk�4�ZX(8�#�U���C�^�D������tm��d���4�K�!��:�ȲMOK�۝�jjSh��#�,�,l��ە�g��6�d��q@vڻ1��������a��)1�X1Ε��I�2��^��2ӻO{#�h�f�v#h��]�l���{u��Z��-&��.��v�Mdс��v���q�v<���ԅ�v�P�]JAk��Psh�\E����غ4��_m�� ���Irk�n]�ێѕ�Nm�N�A�n#�4��^��q��+���)e��-T�!l���ۨY.Yhrfj�"�ƃdi%RiflkX]U������a��l&�e���9*��7V����؜.zƁ�]�7$�8X�m�8�0]�30�K� �#Io�:t���Y���جXy;=i��P �Ȓ���G#&j��OfO{��h�P
��Q� 4��"W��T!�ꁥ@�X*E7@p ?��������,_�NM�ڭ���TH��Joa��,���RۥѶ����z�8-r���g!۬ݞ3��rK��s2X�0����.��	�&��;sIsp�b%6\�8wk����v+�,�(���WH ��h���:ʧc8;'�]�cm'��ޚ*���m��p���<�; Ie��l뮸
t��! [mxz�Wb�F�n4��q[r�@�~{���ES`�o��Iu5�ffMeѣ2��u�Z�-��� 9G��$t���Nnb�Op�Q�տR?��x����v�s�Zz#�HoO�;��O�5U)�R�)[Ff��l�`��6]��5}	6v�r�"j��r��X�\X�˴�&�<�T�:S�ʕ��x���� 9͗h�M@y��ߟ{��^5�I�h�4Yh���P�T��y!h�@)Vڛ�uvvx�v����x�-tr��*U�mu�C�E[e��C�直FfD*GX"9��>|��6�B������P�ǚ�ꪮ��d%� �6�K�_DH��@�,	S�pT脒������`�mX���I���g��J�V��N�`�� 9�ۀo7q`��0��E���~�Wt��&�'H��6>��W��}v�����-�5Tn��$� �n��9�`��l�@�j �eE˿�[�v����nݫ[���M���f�^T��t8��v�|�E*y���Zݎ5��{��@G6]��5:lJw�R���rY��ۭ�9�p��0sn����߷�~�;E@��[e�guX�vՅ��ȕ)*BDD�G{��o;v< ]B9�Q��D�.j�=������v۵��9B�D)��z����UEPSNe��R�;�K@t�2�t���R�¾�{.�<���a��x��{��9v��^��.ٻV�r����z>>�����m��?�gut� ��ڰ?f�G����%����jߩ�� �7ny|�_&Ϸ�Ձ�=���wnK�J9v�隶&���D���{�Mׇ�K��� w��oN�)kv9bsUJ�ϧu�n��`nmXJ���"6aB^�Fuw�`��ʪ�	�9�y{�����@yȩ�Z��5�}!&*18���3,�!�i��6��;]�O��[�yܸ�kVˍ�@���<Q�����j�EH<����W��{!���(�`T"In�����!���`gw\��f��(��IL��ǚ���*�����`gO���v��
!Cfn�Xou����j���m��e�e������<�T��(�Ϳy�K�G�H�TQ.&����5�U��^�}��:H�@}����*VY@���絭kZֵ���V��Uoh|�Gc�VvAz.�z���1��4�M�e��9�	��W��7]m��t��lS�����ݸ�st�����5�nd�1�g��u���g0�8�J���_������{�;i%�ب}�9��d����c���F�k[Qs"�F�g�<կ�b��tKIwnLjl�Q(c	\b��n�۽��vٺ��u�>[���[�qϓ�5����λ7WE����%y��-�jy�R�)T���������ZX��������\zy���
Zݎ�e��<�� ܊���=&� t������L���`��n_&��_7o� ߷F�|�&��l@nj�lo`�꫓�b ^B=�����D$r���� �9�|~w��`�6�IFf�������r΋�n��	.�l�Q�պq;v�5�f�lP*�X@�Id+��@��F'%?��Ł��l�ٛ^�����Ł�󮪚j���R ��f��P�DG��\PНUD�O����{��ܓ��� Ի�ѐjߩ�����ۀzM�?�]�����6�f��]me��V�y����R���V ����5�pU
�ݎ�e�`�� >�'�z� t�j�EH��ҞG�˲�����[�Eڦ�z��x=a��;]���%��;=�ի	����nEb �sP�*@y�� �m��M5HR��SL�ٛW�J�d�{֬�f����l�*QI�L���?n��eie���/�P1K5�	�h�^��ݛ�Ow�p{��oց]��NZ�?�|��	>�X�<�����=���[�Y�Y`^^� �X�<������ۦ�#[t�%`�@H��т�l����78�м���{X�4=VA��n��w?}��F��˭7v� t�j�loa�w����a�KlMU�*�-�=$T�_fgƁ'�+����Uv>5�p�+kv:ՖՀn�;��@nj�EH�𛻖�]�����$��;��̰��X�vՇ�O�j���sy�~7$�}������Z�ѻ�b �sPr*@y�ŀs�����%��O��l�@%�[smq]���ݑ�h����f�۩Z�`y���S����"�)���W�g{֬ّR�����<�L6�n���a�y�H7 9Ȭ@nj�EY�9����լr�@-Xw�� I5�"�n*@J�4�wF������b ��Ps`�m�H>�o}���5=��k�5Tn��$� �ݰ@6�9��M@>ʗswwAH\ݶ���]���o�k.29.wcuۚ [S���%�s���J;c�c1rRӶ7�c��'����$y��j'��3�^[�iq�f�v�e�K8�GR⹣��[{Y��z�.�@.N��=[��g��m�
�H* kp�J�s&�gsN�T6� ��*z�R���*+��ا��u�Eq��R���B�n;7"Vo���f��ŧ�N�����u��8�:�G�t����d���H뭑����%!n�,���b�>��e�~������w�ŀo��O[H��t�U�s��� ��� �ݺ`�w j���kU	��VX�ݫ�nڳ�$�3�޵`o{�� ����P����wq`n*@s�X�=$��ن�o��6��%9�Vfm��7��? }��`~��X��[kv�SQ�nJ��DE�[pj�m�u���<�r��l��#��e��d��t��,��@s�X�=$������X�ݢ��!o�[k0����C��*-H�b�����ͻ#�}���ܓ���7!���3����S�xv��UFꊢK��o�� 9Ȭ@�jYƶ=�)�]7N���BP�:��3y|� wI�s`�����3t��(��ܽ��TT�;��9�@wM��솧*�����s�b�=83�sǝv�7\ۓ8�X�&��[��gW~��w|�`>�Z��iإ_�;�z���0sn�;�q`z�>�G֢������ M������_~��WgO��\�Z(W������h���VV��BI�'M]H�P�ZK�2��' ��{�R\�N��� ���`��Ag�4���mSy�9$T�S��	����b�ٯΓ���p�"ja�v�*ͩ���X�v��š��?�!��Z'aXJ�&`H��b� 4��m�i2�k�%���;����1�)�����@x#��'O�~ M��ǁ G�Dҋ���N��䟻�v`���lT��v )e0wtŀnmX�kK��:��9-��&�����H�����@s�b�?����D��%+��>�C���G�	�l��b�3��מ��Hr*�7A)W��7TU[�o�� �7n��(^�@�w���4�c�P�L�:*jh��v��$ٛ�Z���?f֘�gd[KF��e����1`G5�6���$%��+wn�M��d*��M���s}|`y�p<�� �\��=�rI�l��=#�I�nG35Vٵ���O�z��˭Xy�p� յY*tV�"�@��[fvroI[���hk���5���`�)Y��ki�B����ov��� ;�ۀ~��0���ةA�\`�p�t�}	&�s����� �sj�!$��oP��55P䊪)X�uX�kK9$��ٝ�Voqj���4uN�j��QT� �ݺ`7�pwtŀ���5����>�Rt��`G5�9�ǫ����<�� U]���C#XpIDH0q`�_8�t�h�G�Q�
�����߽��f���.�9�c�n^{sԙ\���IY�nU)���Dڊ���M�,�e�u����:��X<��x���-���;�z^Bw]��Hf˻m�x8"EM��^f6Dp�=�d-�ֈ�gsf���Y����{H������6z�����\��"� "���r���LCd{uB�*��˴�S�%���vl��ؐ嵑Z
J;�]R���/����^p@<��U6�h���Z[F
C�u��Yʾ�8z덓D�b��v5{W�V������ �j�$�G�@Mlzյ�&��`y�pݛ����r
�K�y2�ہ�]�wy����-��� �j�v�+�Z�p��(�x�%��< ��R }&�<�K@z��^�i�{{y`i����� �M@y䖀����t[ҿ�-��' t8�Y�v�Ͷn�ֹ�[��p23ٹ��裸]����ۺm ��Ih�a����;�� �{����Q����j�$�u��WUW�&��AR {ݸ��{⢊B��;^�����7KVr�Q���`}���z̙[KD?�rUe���$��i�� 7��@t�- �� �r�wn���¶�ͤ 㚀��� �"X��+Ie,�@Q�Tq���f�-��M��v�!�m�����Yr&�KoN)���U���i`f�i`fᶺ"!/������B�~�D++�IL7+K�Q
6oi֬{z��s]�g��,T��H����7�{ f�՛�B���nw���mq`jY�F��f��·w/i 8�=1�@8��u��:�{��ؚ�7TU7-�?n9h� 㖩 8�>��U��;�g�6��]9yFۡ�a��6��I��bI״�R�aV�e��a�sˬZM����H�5�Z޳�-V�'�I*�� ��^,�l7��`}Ӽ�ܭ/��L|�U5Bi��y{H}>��9h� 㖖 oSGf�}`T7��}�����\X��Շ�JE)!BC�4�4"��@����t���"�*A�E��E `}���T�S����9�vʭm8VW*\Ӱ3r��:#{y�_�7�������˛����,����ʬV7fC�7`�M������h��ղ܄nyEzc�띚e��f��
��j����0K�O�6)o�
ʥX����9h�`�q�R�ۅ���]j��M�pl��ۦ_/�I���ŀ����ν�s�E!GK� }6�*@z�LA��l���'�[P��IS��y�� ��.N�����v�ei`v��$B!(@����N����߰ˮl���:^GZ��+���ۭ�XP;wO)u��xw�����SZ��I�.��(	��>no l��Z�YW�vˉ����ڵp1�F{S�y�x�6�N��Wrf�g���#/n(�B\��'.�Z���[J΁Tݜ��y���F��۬�9�Uv��[v�
96�ۨ�}��2��r�\���z�[et:�n�h�j���9k*=�ϻ�v^��+s�7S���F����;yZͫ�tC��5g<�\C'kV˰���|ӈTr������0l�����I/�7;�X�ѳ҈uCcr&�q���]�M�@G�ʐ�& ;{v�kM:T�;^���w�ܤ�ɈLr����u{u�fV�nf��*@z䘀��- �� 5.�>�6��8+,� ��v`��xo`�}"��P*m��nQ��r���/n|�R��2��Q:�n*��,toK(�v&�����`ٺ���L���������q����)�Rtܼ�@6�	�U~��c�R�$�I��>��h+((��ZKL���`~{�6tCy���ݮ,~�=j��O�W�V��H\�2K@6�?���`{����'h��r��;�������ݵ`~{�6B����7���*�s�������1�g�ү=j1v�1Z�D9PX@k�$���W-�4�S�*]S��f�������=�@?wV�X��Y)�s���f}�`}���ܭ/�J9,�G&���r*��VݽV�;�̏�!F(J(���t=O�k_����vnI��ծ�j��QTܷ ��׀n��`fnڰ�^ID)�{�V3y�~(YY��zn^m�${�*@9���x�~)sT���EH����Ȼ^ֽ)Y39�[�5��t�\@��n΅effn�� �R ��@9�Zw�L �jc֬�%�U�V n�j�"6oOs�;���3wmX撍�!Y[cpnKp��x�n�ww n�n���W-(ӥN����t$�v��u� �ͫ	���!%�H�@��UMwZ���}��Q֪dV +%0��, ����%�${���f�m���8���v�e�m�(d�@���;b�;=� �r2-_;DT�Rߜ�U��ۀsf��7r��
>��{֬'ܼ��t�k+j�7Pd����H� H����яEH�(�,r�w�L7v՜�6woU��=��Ǭɝ���
����3t@9"�#��s$��n��яZ����r� �sPc����8� �k��uZ+�u��J��b�-�"�L"�8�$i)A�H�0�����"�Qt�%҅Ϟ ;�qC��0����ˣ�af������	OƁ�	 ��4��B	�F���`U?#�4a�È. 0@�C�%"�
��(��(L\?,����� @�_�P�bJ(@��[��,�)��TIC#�V
c$(@�{�ӻ��w�w��/���Y@     M��-��`[A�  $     p����ۥ�۶��P�c!�(�UZ��r���z74(����˷D4��ݵR���pUT�\�4�%ֳ����vj�����.�u!s)��)�&eH�X�gky�J� L��ȷ�>ݳ�N�gv"�F���3˵���M��8�硪�De�[���v�t�n8�����ˑ���	��S�uk<}W��V�֣���8%�g`"E��8��8zp�n��X ��9�Vؙ��Y�T�\�S�����K2���
{`��26��!R�-Ѡ��ԧ]C���M�� �(qsB�R�j�.��	�E�:�eWj�i5z�3�E8���	�t��s����mMC��;;�����������Y�Z����ʞ+��t+�� ݵ�#��q̴^��D�"F-�[R0������ê=���h��2)d4�+೒��!�+�i�͞[��W{:pwX�OMկ.֌'�ה�<�|ֹ�n����̪�WÙCf�[;jgP*˰�aݰ��綾�1�l�9]s�\����Y�sve'3���v�n�l�v��Np�lM93�d�q��4���h�td��_(�Ac�g� T�kdwY�[�d>� �&��v�TkR�Q�c�y'Շc/)Z덥Ŷ{;�#�x��w����.z1[���ȥ��+l��oA�ʜv�k*���p �m��A��sC���V$���<���ps��*�i�4���Бtm�X�9�o<8㔥�ە�y`$���(V�]E!��Bns� 1��f-l�q���&j��{/�>.r�[V���X�v�;t,g46�[<������N��U�WT�9S�3QI'i����q��P��[��Wk]��z1����.s�@[��v6D���U�ţ7=;0ک�VF$�N�x��[��F�=�'\��l������CU��so��3��ڬֵ��n�T蟁@��!�ڈ'U�,j���Q�??UQ��P�P��7�B�����U<�	*�[��B�}�-g
��;m[����2n}�Q�i=��҆���=c�9��:�-\�qZwfv�s��������Wg���ݝu��nGe��(Rwh+Yv�S���Y.����s�سn��of[�u3�w��uȎ�m��/i�n��.ɍ��c�;:v�mL;��B��zֶ�6�!�ͱ���ځU��ٛ��t$ۑ� 7ce�i�����x�n��^��`��7Bެ�-�pmʃA��6���#;�����3��wu�g����`��3v��O�#� qR ��@w{v�ki��q�� ���?ě7��Xv�X���yDL�{���(T�*��U3E���Z��ڳТ7���{�|`�v�X�RQ8}m� H�9䖀��~��s�H��^r���*����������o�� 7{� 9��:XT��`�]�O�Kl6N=��I��rn��b,y9�$M��81�蜅��W�o&��<�T�'I�x�=rǙ6��Ы335��j�Iϻݛ��� �����=W�7�����w���1�WUS�C"jY*�w޸;7^��׀s���f�`��KA��۶�{�}������}�>��Vo3��ޮ��mm7]N8���|ݘ;�� 9�ۀs�u�����(&����A���ۃ*����=�9ӹ'���]u�u��챇i,ed
�� �wq`9�l�s_/(Q�����[���S4�$���`}�W������v<��wq`Oz�JH��QT� ���n䟯��78�����6T����ŀ�pb�Fle��t��v��%������� ��ڰ>��x��cd�G%q�0��ŀz"��O�3gy���́� �[5�`��c>+�;V��sý�;y�5�O8��=�VL��g����xb;}K����~m��� 9㖀��1�"���{`J�i�I%�;;�?�l���0o�� ��v`�݅r�1��Gv��I�9#���r}�2}hϺKEYTA�`%�K����,	���7$��}۹1��Xw�y^�̘�f���RVJ����Жmo?�c��?f� �f�D�j�<�Y��){k3��3��;s8��L�I��Sںsѐ��a������h\�r*@;rbYM�/p�J���;绳~�����`k��>��w��ϙ�z��iS34��M���Z�1����
"o6w����� ��ǭk��7�J�����9h�& <�T�:����tf֦��fj���'5�J2{���Z�1���	T$�B�"�W�������5�Rv+���b���v��F�%�z˻C8�	�{3˺�.ˮhݛ
\�����7�u���1-g�t�<�d9ݢ�ˮ.֠x�ɾ~����N-Qطari �v�u�M��^���7[zЫ�&ݖ��-���� M��u�z�dRِ��Ս�:KaZ�k��m&n��Wl*�qu��:��(
g�����\��@�f��[W.SZ���3&f���`��v�&���OfL��g���s�<n�)�s���)ub���D�gC] j�%����>����ܘ��Z ��%dEQvY�~��,��$ٯ}�wf��{�0���#SMHu[���v��<r�rL@yȩ���]�4�Fꊃ�`���wf�����?��^�S����b����y��zn^m�:䘀�Rۓ����h�O�?�&�M0���1r���d��9C��5��B�'���cW�dm�9`�$��l�7�ŀu�v`���wf�яZ2֣hn'+�X�vo�,�Q
?�*�zo����zl����.���KA��$�`�;���b?��O� %Ͼ��فy���&�fE.��yD<�ޛ�޵`c�v`�;� ;��X�dU�vـy���U1��x�>�\s�w�-��7lt���*�h��v��Q�kr̶!��{7V!:(����r�c�&����ٰ?d�繳�D/(�C;�j���/9�#T�n�RU6��`u�1���s��\�
��J���;��ٰ?fm�"J �� a�	��0\c��!CJ/�v��M����v�f9ږ��fff�^n <�T�w�b���ـn�c֌���L���X_��9h\sn*@7(�vR��]�{tur8;؛f�6�ட9Kv�{-n���}�A��\�`��[U��ߏ��9�7 ����0/2�����+/v�䖀�qR�I0ݝ׀~}����T�#�v���H�& <��@7�ZU_K��i����NiXr��{�l��v}��ܟ�8FA^<A7�w��|��˘�u��Tـof��;ٺ���,�wf��M ��`P�C�.����d{����뜼G�2N�b�Kp:�SV�i��J:��nB���+������ŀq���7�u�����Ӕ�Il����EH�& #�- �Ik�}��2��ȝ� ���0��h�K@G"�)���Fn�������K@7�Z9 ������m�"+j$R7k�;ٺ���繳`nN�5tD�!F�TT�8��l���MdΑ��[=�ȷm��R�v�V�ғ��u5e�
�<GF�3��ۛ�۝dNr�sζn��Զj�Pvnk�vM�;sK�Ź�K��7D�s��)����r"!9kr��Q
{u�P���o3&�%W'���;e��n���l���{.{�c��Mh�q�>y㥲4��i�X�;NR�U=��_��t��r�5�5�5���5������}�Y����=��5���6��r7d�lt9n���V�7��8�f�[9�����5���yAY{��?���R�I��K@7�^ԟ5�M�ԁG�rU�q���7'u������W��l��C���n7b�� ��y���x�wǻ� ��΍�ta!FV����v��繳a�
��`s�k��jJ�	�Y^��ŀ|�˳����{� �f��"��F�Ϣ�~P��ѿ�@�9Yݡ�v�CY��)����7.!���"ch����D��\ ��P;��h���j����Ҍ�ڻ�33Z��;�w�u�D�F� �P��T? mP&�����~��,�{�?�I����¶�j$Y�{���>��ȩ�$�y%�?>�h�u���q�׀owq`{& #�- �IhU�	t]�Y�m�S��`|�vl]����=���ݵ`j�5mr�X�ӎ;@l���CkkS�25�W�)�ax����e�����H����@G�Z��ȩ�nb�:����B���+�?w�L\���� #�-.Yəu�]]X�,��7���ϻ�ھ!|��D!�E2)F �S�z��̍���D�	E�A�D?[������	�S��| ~�D�~(�"$`%L���'i�0wz�	��h��-G�7 Cn�bmGp�1T?0H�X�H��?�?,�~a 5!0���`#"�	T)�I~`� �60cA����"bmX�%>%La�	����O��eC`��5$ �>� �??��9:h������xA�
v h�u� W�1$Q�,"�pS�ę���ʉF!X�"�*�pb!�:]*1t 0�"=P�m��*pD6
� v��O�Ѐl�@$AdU#$An�1郰��EW��`}�ZX�1�E�0��%:R��P��wzl��v���áB�����, ��Q�Q�i�	$� ��o`����Ɉ��V~�5��VvͻN�nҝ�i�#Ǫ\;m�$u+&V��s�;�;�b�� 9��9 =m���~���}��;f��7Z��I d��7���ϻ�`nN�>̭/�!�R��m��B�������}��K@s{r*@w���1�t#v*��0��x;�����j�bj�$�j� ш�����RB$�V(H�� ��+%!	V��1%�`�V$VQ*JUD�IZ�Ҥh� ��^�lP-���rO�v�=���J�/o6������&`ٺ�-�0�9� Et��_�n-٨�&�b����P�-lv��O)���
�2��%��i�������ذϽـof���>ݮ,����	m���X�n��gl�;sk�sv��g3�G�P���N�If���;��ȩ�b�فw�ݗ���VKuN�ϳmX����sfá(O��� ���n�S�� RZ���,��ٰ7'u��m�B�Pb���~�.�wK(Ѵ�̉�u��^����0�휑��6z��\��}���
V�U���m��֤�Ɉ��*s$���#nvF���ggKp;sv⺀]0)�r��#����z�Lf�P>�v'\yV-���G�Z��hV.��k��	n�ֶ�����k�
���kM<�ĻqQ��L� � �&�v��VY!�&+��`ғ�5ۧ�����������#���W+A
DJ�q���j�Y��'`nSʚl<4tS�������~��ݯ����y%�8�����וȝ:�@��n���T��EH\s����7+0�ͻ�ʹ� #�R��y%�5�:8l���d�`��X繳`nN��{�ߕ���4\�L&�*���@z㘀�$�� #��7d[[N��$U���Q.��6W+;d�;&E�U//7#*��y�y&����e镙���K@>{r*@~{ݘ7�`7
��S�Hݯ �;���?(�j
ʇ�#�9��{�,���of��?vl�Z��B@*�4@G"��I��K@6��ɦ�	�'[�YmX�ـod��|��T����x�.�C��jl��v$�so��v�Z�?=���_'�o��`9S���!�Mڑ�n��X�p.-�5���v�����Cp�����4�n��o�G7������7�u����l���\��r*@z㘀�$��_�������і�"��`����n�?@O�	���
頄�4.� j�U4mJ�lEC ���� ���X����P�Ut�9u� '=��� 	�j���V�J��Ge0�n�������������X�w]����m��S4�uɎx�۷;��ⲛntb3g�m
�H���NKc��:�;T$9)�s��`�5�Zs� Wd�y[�~����5�Zs� ;�i|�:;�sn�E2Jj����>ή,	�`��{9�@;)˺�V嗕��w�� '=����T�??UJ�D�iSg�%�}6Np�?=z�����7+�� �{� =�`����i[��~�.�ۃc^+�Ѯ���X8�κEx�;s*����8g���9�v�������>s�Ht� '=����� �|���R��:F;V��u���0s�Ly�Ş_�Cw��p��]NeL�T�oW�ﲴ��C}�֬�{� �݆���R8�9)�s�� :8���-���*�|f9U,�M�U���ڰ=�Ws��W�wn�}���U�m��k�����g[��� �&Z����v洪9{q�v�V������ �l=v�T]�_m�5�O�����ޭ<�8���!櫲��;��Wl� -R�\M��q�n��Ź�Ԏi$�9��ɓq���cـ�6<i�=�5�2�9`�d5�����t�Sn�>����un�R����k�հΆr����]9wC;�<݌����?��T�	'9��$���Cm��w�%D���������fޙ�\����d5�/�.U�$�y�c�RO������ w9��*@;)˺�U���if��f��`�;��G ?sn���ׯGAJ�Ս�����>��VBI����s���#֋kB���$� ��q`��L�ۦ s�ۀ~�=Q�Rь(�v��@~���^ n}��*@~} :����؉c� '!	A��vt�YT�*G�#�y%3ϫ�3D��;�qk������T�9��*@z=��6�c�H�� ?w�s�� ����	5����!�K�CN��К�k��M��U��e�)���>��V���΅�wZ��}p�wG1��Y
�RKV���`�T�<��G '�.��V��������T�9���*@y�� �7| ��6�h�_��X���r�;sI؇�g����H=��*	�x�����{�� �F�n[-�p���s{���ۦ�n��8���[ZMD���*@zM��nj��=�
Z1�-X��� �7qa����:ߏ��L]�UN"��B^��³����;֬��z��F�*r)��;ͺ`9ݸ5wq`|��}�0zz�V��	��h�;��JqR�6�`�8�lN�ЎT6X:ڐ������^:G$S�Y�l$G�����N��=��|�۾��c�U�n��O� =�`�}"��ݸ�����h��j��`��L�M��֬3z��fڰ����6��ҳK���T�;��JqV��t�8��8l+e��e��(��Jgw�V�w�X�����(Zf`!a�\8D�BP�S�`�F>h���)�M������l�T�;����klX�%�:H4R�B�ʷ#���L6^s����\C���m9v�I�utvڄ)�Vﶴ�3��V�ٵ�
=
>�����X��CpU֪r)��;��W��f�X�zՁ��/�l;���T��	�� ;���9��� �ͺ`��,�rh-M�� }r���<��XgW}����&�7� ����1��Y
�R)j�?sn���~������5$���nI�*
*��TU�TU�TUh���J�����
*�� �*������A@��P�AP�T#P�UT$�P�T$BAP�AP�	BT!BAb$�AP��*AP�EP�B0T#B0T#B,B,U��P���P�*�T �$��DT"���T �P�T$EIB AP��B
P��AP��B �P�@T"AP�AaE�B�T �T"�+B*T"�P�B�EB
� 0T @T B#P�B0	B$@T$U�T"�#B 1
0T  $B(�AP� ����0T )P�0T"�B DT"�T"�T �T �T �T �T"�T"AP�@T!P�B)P�+B$EB$B�B
 �T"�EB ��P�*�B*�B �T ,B
@T"��P��B	P�B(�T �H
"�U_��_�TU|�(��EW�����
����*
*��(��ʠ���J����TU*
*������)���=��~,�8( ���0�'�       P  U@ ( �  �    �  �"E*R�(*%*�HJ�P�(R� �
���
@
�!J( 
PJ"R+�   �	     � }�)�����ng�ӓ�\�� w��ώ�Ǿ�_Zy>v��^�����VmB��� ��=����>�ֳ��]���&�m��y����\�wϻ��t��͹��  �      l t{(�O@b9޳��r©� 4@�{2�yq�o�������p�����7��wg� ���'W���4��[}>��c�ק�W�{Ů���o%w��CK��׽��ܻy��{��v��,z��>�     �� �ϥ9���w�n�B�񲔡LM�� ;(,Ɣ�,f��,Ɣ��YJR�p�ܥ)G6QJR�i@ (�#JQK,�)F�r��,f�R�M(�14 ��P�� gJ14R��nR�)q�R�7Y�R� Â��    �X h�R���JR�)J)��_t���m�� �����+�]i�wm{����}� n��{��w+�j����y��_}� =��WWV��u�o+�ϝ�V��� �����g^��ϗ��ӽ�=���x(  ( P g��+�J�ﲟ{>��]��{�����n� \�./p9i�8������ {=�2ܲ�y  q�����'�[{�+O���>�������g_6�����x=;��=�<�����]�6�x   �M��! B'���)P  "x�T�$@ 4 ��U*G�R�	� "����ڥ)P  �� ��
@~?���GU������Ï2U<Ǔ�U
B���/���*�@S���*��QU����TT��$��Jz���M��0LM����k�~7�F#b�8g9��*F�,,-�B�N�q��I����L�r� 	`H�MB���6O�>�Ա��@�~S$&
W���D�A`Ӈ�Lq��C��.S��
�!%p��	"��
��)���HS�Q�C�)��ϭ�w��:'����#���V1S,��HG&�Ȑ�H"B$D%�.0䊕�M��F�M�����t�+��l�;�'#�5�.��.v����rv���$
J��
A(1n3�Cz�f5�$�e�����%�H���*`H����B��,�H\Jc�c,>Ħ�0$R$dH�%�]d%�����sp�,X�C	&WGƘ\0&y�C�y�#B¹BH�b_�`��I,.�H49ƌ
Bu,7�#�2�����B������$�L�	�VYr@�'����������>b�� 茗�.[��9����s�c!I$rh�N��i�%Cފ�� Q�B�VW$�X�|h�bC��'0|q$$#B2PĒ�0ZЅÌL6A�$B�$,\C�Ħ�a�#�bK�Lna�BZS�d`SF���\f�h�����	pM������)���w��8��B6�۔���0lk*Ak&��5.(I��l�]�!q���7����@��6��\�%�`�!��J�l7����K�S7��.�1���ape	V)���>�CP����/L	�D�[1�o\,�2]�lc��I$�`E�@�`��0�t��J@&!L�i�[��ԊH.F����BEL,�π����BD)a�A)����8ĵ�F�r���S��$aWL@�B�$��tK1 �MD�	�H�2F$$`35&-��2#��`F0盁�֭��{�.!pˌ�1��P�u���M��7&rq�
���@,��s��bX��i���c	�)�sht��gP�Σ�]��$�C�#�X)¦���P��0Lfj�Z�s���B@i�B�5�Mj�\C�3\�VƆi!�э0�ɨ���~!n\V�(I
�������@�0ʱ#�S!0�ɋ��a`(D�%�B�l)���IQ���F�q ���RBB�]�t�[f��\���-�<�T�
�m�@w��s�>����	"�+��!e�ѿ�Id4
�d�	��.�	 H+�B�as��_!Q$R�K�����		 �a���$\��k�7�@��V3$�`I��3�8�2@�(c!)��W�ԍFE��O� �Q$p��M$/600l>`��ۃ�:�@!����ƍb8�l%��#�3߸T`bF��\Z�Is<�w��&ȉX}���"�p��HB4ØX�$��$$L�-D��H}��6`�)��d-b�:I��3`�����@Ӡ�ðБ�@�ɫϷ.4I�툓K�n���}P� $$�	4ک�/�:1��r�D$dze�+�'5>�Ʀ��4e��pd։��~q7� p�$�ɶfow}�uv|B}�\p��H�ˌ�Ѥa!�։K!���fnfBV�VII^k�����.2�9�H�X�0A Ih��[.tљ6cXpH`ác1�ˇf>�^�)�$d�
�)���%��YI����)�9�l�p��4l�6#Cd"�R�RYϾ��A_k|��X� \�u@X����0C��"P�G�~�ӟ�4E��E'�E%F9j� s�i�	\�!Xцrb�ˌ�.f��K����1���&�,��-�3�`�sI�	@� 0K���	Wd�\c[7�w���ζd�j;���a"�a	 F
B���ʺi`�T��.(Kq.L�"`!F	R\� ���f��b�
��]J�DR�7h`�dc$!���H�BH% U�d^s9�Sy!�.	_���m��f័�cF�NϚS[
h�l���c@�2B�e� �C&�>O����2M��\a��4Đ@����B���`��9�X�a(D����Ը��Q�6#H�drL���N� �!L#�
Z"B1*Ja�p��yL�1��
F��8��$HH����}Lh�S��ҟ|!�!ϧ1/5Յ�#�S	��T0$���P����RS��B���%1�0H��:�w�A/� K
1Á�S0���;�l���U������2r!`Ba�k쐑̦Dٽ��a����
Ct}�댐�.�Q�#BQ!@��1���HS0\%�R��XX�,����۱��!���RVP�`E�>�a��d�����2j�S�s�GC�����b�X\�f��
d��H̛��Pí�4m�&SL
�P�0�$�HXVXG�)I
n�%*�bT�`X2C&�52����`S��\��%)�@���0$��S�Zbc2�h���L�K�c��j�RF���H�$���:Cr�8RQA�h2�x?0C�,4�Gfw,B��b��ŏ�@	�Wm�9�ЂGd77�߹��|JL���a�d����5n���p�8����I��j$H��&��.V�`$H�ष.S	� ��Nk��)�ίƙ���q�A��Jad!q��D#��d�7�$Kl��%1F�aFS>6@�L�q.�VK`���J� �$�~l� �//U6�!��H=�n���&3�جH̘� �BZTc,bFI1&JJ�e8� 2-�%2���	�� H$�l��Ɔ	0ÉfԃH�d�#	#ɈC���`�0�+"Œ���"R-R	BI7;	�O���B���*J�$I@�V!z��k��#pn1�SW�P��7"H) ��9%Y\1
�I�����Y"6�%�N����H04�h`�I1��&�0�50CF�)�$.W.!���X\�1
bg�L����Ld�\f�A$���]��tٞ�  �8�#N0,�k�0�7�<,Jх$�D��6��D�21��!���B��HG�WHWd4�tm�%p�]!���LI4�)��&.,	�����D�D&�� RP	�����q
ă$�@�Hč�D(�Q+i��*UԄ�i��7�Ne#S+�X��܄WX�]J"D2Yf\T��w%Ӛb#I`��J`!���i�t0c$m�<�BD�|d
�#�Y��H1 �G�����#�� ���Q�rR�FD�7�cY�ѫ�Cd8��+��B�A��d ;)��0�P��40䐰��#�	���	H�cHc#&��d��c�z+ӟ$���F��?j<��دzI�H�Ą04`Hq��)� hMԄX1��0 b�M�X;S��"�,
�&Lᄄ5��-�.&�3�\I1�:�%+���L�!F�!B,ֱ�C�aBA`��H6�1�fHd�\SZą9��ó��;X�`��%0K��1��\����B��ь�B��P�"C���G�s�m���s��b��L,"D��k��}�������iLVB�\��ϳ�rXof�@�E�:)�)$�E]�"T� Ek	�$�QĈd�Pp�N�Bd���gZѕ�"ⵁ�k1����,h`�$!F!��D��
be�m�f� @��I$*a@�!�A���j`�wd�v��Û�C~�6�
�kf
M��`P�MI� H�2jO�R%�]��'��	�� `���Ջ}�π}�E}D�g�$�D�&A ��   @  ���    $ $    m�        l                           �           �  $ l� ��-� ��       p                                        � ��� �l  m�ىIX�  ֶ��pj� m   He�
P :���6���5�6� J�M<���S��uU@�ͭN�RH�8�4�m�TJU*� 9�@�Z��U�L��z��-��[S�b��)>Lގ�� �y,	5!ګ�m����͖��z�    �[�m�m��j�v�j��Z��P�QT��u�荜QP\��pj���w�t�qh8ڻB얇��Hj؍����@��َ�/ѭ��ࢪ(�>��UAۃ�zBk��H��C�4�rM,���JSl�IW9�6��)�m� �@�s�մ$ƴ	$t�F�U���0��z�v��/�F���`�r�UV�U d� �    �p�`l H$l�N�i5�I���`[@l5��l��:�-�H �ؐ  �H����m �H�m��l��K�P�ڣa��d�mh�8�H�x p,�1I��
�v涥3@�UU[�JO��#�:��Vݸ�W+����6^m�s��E���l����8��ԯi���K�,��^�m�͍���}Z� �g I��N�H+=���9g: *�m�5�I��m'[k` �Sm&R���`ږ��Kvy�h	����j��� � lA�%��Y����f���%P�d:��� +�����,���\��%3�.̭,�=� �U\��h�m�mm�m� I�ۀ�5�ʪ�K�8U��U�m��A6P�0�@��1R��'T�/.�9�^��&�!3��꫋n3���$�UM����m=lF��N�C�����IƸ�D=�gmlpq�Vt ?C�|��K�
��*p�@U�(UTZ�^ܼ��7l�� Лn�3/���:r��T�"�Ѷ� ��b�Ku�b�I�$,��$6�E��2m&��K�P@�6��SS�%p+��HL�+:�5]4���bAmk��=��蒇�); ��KU*ӭ��ڪ� Z�ĵ\��]�2m�-�n��`:j��B���s�uU,� ��9��8��-Ul[@
�Dg��F�d�����q&�_�k樶ڐ�^C$���&� R��z��4�M�Ԓ6�^n���UU(
�5R�������'Xsn�Cn�i���I��!m8 $m��#+s��W�g;s�;��w�
�i���v�J�wSO+U[/�W�@N��y	�sd*6�J�f��MP1�� kh*�Rv����x�ol#��󍐠"S{uKJE�~1]�|�@�h0q���%�i�kn �c��I��kj����l sl��v  6�,����H��!���eu�Gki��^dܛ5M��]�WeV�
�]��������j8H� 9mHOUU[P�0�8�r^�v���Zlon�f��	-�G[�'ù �v�[�36�H����B[��7A�U��t��5�m� 5�D���  �lI��v͕^�Y�ʼ�+�h8[B��m��ky��M�f�Hm�Yg`n۰	e@wK�� pm�n $M-��:�X"��ԫ@J�*�!��_5QeR6��K��M*�-VÅ��u�Wl�m�U��)v�J&4^��^[������ղ�A�+�+���Uu\i�/UUU)+�vT�p�H��	V� $�OR�*ʷ��}���u�7m�S` �-�	/Ye�oP[C�C(�Pm����T�6�v�� �5I��u��ZU�������F����M�I-�����cIY$z�;���M�p�ԫ�k���!.Nzx=1��L�m��TVη �U�;`�X,bKe8ċ�evF��M�l=;U��@J��RlM@) d����j�q�[i�8�f��h����ȶLغH�$�Ă�!aUj��V�j���XGk�tVQ�j�0�nqe��  ��ē]�t/^��жJ�[��;� dm$/-U@/-*ղ�:�`���55UI�j�W��Z`:����E�h p  �X�g�/d���&8sm��˦�nv�*l��%��I!wl���M�%�-�6ؠ{2i
��� ��v� �6��l V�� ��ln�v]\ʹ�ݶ� ��Ӏe��m� 6��I0m�M�Z�k]Ws`䀐��m�:@�!JI�� $p�ػkh�:Kj�imm��b@��  ���������ݤ� ȶ����������j`$6�r�*�[R��Ң��S���WPm[kv6��li6����C�x�8�Eo<���S���u�(���(�wT������8�]�I��p��M*ܐWU�Uʷ*ڥJ�M�[A�uIpְ[gKf�$$	  q�YQ�vض�p ��}�� ���[zD�m �`�M��M#l-� ��R�K�M]UA8
�T8�hu���.�\�;m��v��-�sm��h��]W����A�� Z��Z�����J.땵�1  5�!����a�W��OK�Q Ue�g\�G!7@U[UUUe�X�cm�U��$p8�JH-� k�}'׬����k�a�H� ]�&V+��ݎ�ٕ�y��%d�vscE<�"�����:�(�]&��tv	�M�H�km�6l� ���P�Ğm�����/^���X����D�����5���[[p im�M�pnZ�b�m  	YRq$�mm�M��:&c�H-�;m2�m�ڸA� 
U8��� ԁ"C�]n[i@��l-�	$ � � L� ��m�� ��	$C��Z�*��^@Rm�E��@ h	��T�&ؔ�UP.m��m[ ��nݭ�I�l@ݩhq��Vatۀ $��oMqjK%��An�Zp
WA��5l ����Ԏ l[@Zv�[ն�ݴ�m�$�`8p |ݾ��6m�:�� pE�nl� ��`�b��Gk[[V�m��  ���!�m���[Km�dl� ��\��M�[vpm�`�\ +T`�)4�ΐJ���D��s]����$.x���J���nP��8j�^^��w�x X5l�h biڪ�b�P�25/+Z� p��cm�`�����u�߷l��[d6��v� ���K�dv��UUU+�2�l�RlM�d���`��M�  ݤ�[X[@ky��@	�z��   T��r��*U++Td�l [D5���P�K�ʶ�.�GUl/<�-�*�N�Z��H7#]�&�,�H�[|jZm�#�Nkn[� ����qI:�BM�f����mA�Zktt,Pl�L����K��n�� ����nXuN���� %Y�~��QY��yΖ���Zְ  m!n�.�m�6�	 ��� ��`�������E�(��U*�ժU%k@�km��NR�n�n�6������9 Hl  �.֍�` � m�m[E�  ��B_Z�]6m���f�p mm��� m� դ�[KM� 8$t� p��Ѷ�.���m���[)��&[\  m��(�g�-�L�f�`p�i0  A���ju6�9�f�H8�] ��G*� <��`b�hH m�@ ј�y�U��@�yZ�+�
��S�;k�.�!����Ym��S,��S:AcRf�Y�kh
�*�� m[:t�T���l�i��kb�.G-R��[@ �(&�[u�j�W5�*�	 ٴ�v��\�%X�cˢ�'�tp�q�jD�5+�g.Z�lj^��v4���q���@y��]�W�T���v�U}WmU�Ԩ3�É�ܨR�U[<��/��6�g���~�'�O+UV��T��I! HH9��@�ln��	�L��*F�H�  �VԎ��&��n 9m�$�9��[%� ��A �`��Khm�v�	���e� 8ɤ�e�  pͶmm�I& �#\tt�`5Mv��倛Irޠ嶠:�Tv�d���j%Wh� 𷍀I�m���&�յ��5�0��zY�b8RX8-�� ��k~�m��5Vm��&��v	��;$9�:�[[lp m�i6	�l�R��NU[�@UU[@��� ���L�R�Ua�q���S�����b�=m�d� `�v��p-�5ٶ� �@��0R��PK 8�-�M6� -��a"ƴm&�s��$�jj�r�::��H����eKZ^�gW�.eꪪU�m�O� �h յ�N݆���k-uR����@PX�뙌��.1s����  �� ��&�~Z��'��
��ep:"0 ٵ*\*@Ё��
��4D"��"&��CD]#����\��$2D4��>�$أ����u�U�t��(���.D��*:���WA�|�Pb�B$X,b�`,UH T:? ��?<���m��P5�x �T~@����� ���IDF<ʨe�@ا��z6�<�ZQP�<^	�8�8��@�dX�^�!@~z�<p�D"̓�(�A�*� C`8�(H�A"E"�dQL��D��� �0R`= ��O�"�<�@@~AJ��$Rd2(@�`��4��?1 :�� �bB���A0t 9N4Z ��N��M�: ��t��`�*#�C�P�q��8���/QH��Qȃ �@�(Z�"1# H�b�~O�t��J8�p���lT9����L�#$*�ib�d�c(�i�$b�[�~UʼȩP����Ȑ�T]��]!�@4�Uz�PN	 ��HA� �T�л �C��He<)�!�5�.U�Q��c�*/��?�QUv��@8��H��KPA
!��Pb,QbBI���B@8 H8     m� ^�nِ m�       f���l��&�W�o����s�;ktwg�E^�؝�{[K��W�c#���Z�М�S�v[�[�Y!�Sg��M�l;k&��n &��#e�I7��4I���MlY+���!���V�']���@���3���k�E��Wm�)m�js����h��8s.i#c(��}qY�.^��;��.�y���ְ�W[�ll�tҽ�l�E�`�7Z��"��ճ�c�dBZ�e�X�7����o%��0;����g<�ý��k�!��u��G�ʋ�Y��� c�e���wl�/KVZc���ȯ,��[�6�&�4ѱHu�#[aa��Z�;�'U� �2�x�l���˜�dn!�u��g�D�\Nks�4���4�vOj�ۇ�v���@�l�;q���9����w45�W�n���3�;j2�P�V��x���{g�G2L�f8 �[������.u�c]�q�C[��K,�|��H6[u�	e*��GiݳN
^�;�W����\F�a�
:L���m�]2gv���燮mn1 Lg+eNɩD��������̫n�y��iz�UE�ݎ$(�f��
ԯ;���		��N9�^���Kie�\����J�,�N4��`��x��]�&kpb�uqt���B�j:Ty2! �γ���֠�h+��N��c/PS(�j��򂒄��DEs��dv�
�-��1�(��<�#���X�aZ�R@��]mT���Z��ksL�.aZIH!K5��偪��@��us۩���(����8�Q�
��l��Pɔ-]g]V5#��bZ�=��[v�]���������t��74�\�(Ԇ��eU
���
��a�m�nwVn�He�i��w����=����ꜜ�ie�Q��u�]��L:)m��a'\9�yՙ�u&F�Y��m+������Ǽ@�%@�S
���>Pʇ8�l��J��w���N������ma������ӷb�,�{B�ڕ:#n���u���F�;0�2�����gr������|v�����9m��8(8��>��Ŷ��t���sh^��K����۵�nj����j��ѹ�������[-ζK������IK��*��ᛁ뜋u@iUH�e�{:����5�q����q�r�3���s��� �u�Rۢ�]�8�ێ��.M�.����<<9=�s�;�<9��ԟ�U���v�=�*����_Ñ�ܿnhb�(��1䄊&�$�略�8�*�����T �� �[�7X��'�$�.��}빠^�@=��hە�o\"q��1�@{�� �v�=�A��'�� ���Y#�jB9���4��٠r���=��� �ҶUc�̜�i���R�i�h��m���Hvh��7=t<O�F�0X7�S�rM �=�h>�Hy���@fCjffb�� �E�ܖI��q���J�T(� j&�""y�Dw��;��{�G����O+���7�H�}�s@<��>Ď���Uo�@��^"��Ě �� ��4��٠r�@��w4����BH�b�M �<ݠ2'1��mB �n��=p�u��a��_g����U�wF�3��÷\�R�<mfv����b���천�{r�xV��-��-�@;;��/\�z���n=�e4�l���4]��߿y�����E!j�6I=�vY$�w�,�*�$!+>��(ax�8��{���'>�i�{�Q�&�
$nM���h���<�S@<���Ε	,rq%&h���<�S@<�����I� W�:RГA#	In�N��າ�:����n���'��hZ%Cl�R�����7�H�߾��h��s@��^�W�D	��M3V ��o"&G����n٠\W8n�7��hRI�vw]��uzn%岚�f��Y(7#X��&b�f��ޯ@��M ���`��"�r�zc�ѩ'~�{1�k��87�!��-��/Y�vw]���^���ʔ�1�$��ț`�J���^����m.z�A9�Œ��B��']�������$H��Ӈ _~��gu��9{��g�=���w_���,�F]�ݠ23�z����^;@\�ҡF�I�'bRf�޻V�岚�h��s@�{��`�Q�
�����A��{w� ��@df5�j�*�׈�QLohĜ4�ݠ6!�{����:ݱ �9\�B
�X!�p8 ' �b	 ���%�1"�������m� T��5��@s����v��:<ݩ�go�o�L��#�\�p�vx�^�,Qݲ��Q�����w��{m
�sc����g�:�v�x��ܜ<t
�a�=�ֳ�L�	M��b���tW�F3k�[\.l-�u��v8����rcX8zz;J�,�e��y��Q���D����@���Շi��{�ִ��=f�xYI�9��vûs�rv���r)tj��[$rv�IƤ�v�Oe�C��������\���v27uB2��[�8�s�Sv��h�0��,�!	����=��Wꪤ��?�Z�_����w4��F޸D�xbjE�y]�@=�f���w4�ڴ�����RLmŠ޳@��j�nP.s�Ȟ�nP��TLX��Da�I�vw]��v����O�ܖI�*�1���dP��x#�0n�[��띦��[%�͈��K�^�gbch0b��c� �A�I�y���<�ՠ޳��\�����<��MG�c7%��ԓ}�{u��S�X.Sa �(�h`���H#����|���O��gRM�w�4I��1]��T�����0���!7r�3����� 3�ܠ:�@8l�Y�jʎK'E
�fo�^|�+�h���<�
\�&5!�����w�ՠn~����_��Y�\��h�P�Y�rA~I$dSH����ְ�c*#�q[Y�I2T���%��ێ8����h[^�{z��s@�]�@�x�Z�<HqHEr� y㵱2ln��ݔ�� <���Đ�1�R9&�r۹�s�w�R�Ƞ��T���ʁ�>S~z}�M˝*m<8���=M��n��;@8m�@uz����Y�'�U�����.[w4^��U��V
1H����#�y�9��n,;uv�c��{n
���Iج7��KL���3^�x�HL�hM�� �z��s@��@����ՖBbbB�e����832��PH���N��vI?gr^�H����q��R�
K� �v�[t�<���mB��o\"q��?'$��ʻk���ԓ��q�Rt3=�Z.��7�M�@�L���N)�nG�ޱ�����sv��� =��u3s5~;[O`˷XL�������έV�U�ٙq8��+h7Zs0�Ɲ���[o��҄O��e�H��:�-�6ڊ0In"R�$�}���T8?-�z}�M�^���sU��q���&D��<Vנ޳@�׹�r�נy��o		��M	��{z��^���^��^;k�<���$Bp��1�G&�m�s@��@�[^�{��d�TѪ�լ��$�I#J�� 6�t�C�vI-z?�}�ON����.1�Z�������[���u�%�{b��vd��'v�-����>�ѥ��l�۬���<rtZ\��q'�=�}ṉ̝�f�Sg�&(�q��.P^j�ݚ9͹�ӡwfV��i��;�@�����w��.��4һ���ͩv�z���nM�Nŵ�a��y9���ٶۙ�Y{pg?!� ��u�rI�L\��e3���z1�][�W4��ݵI@�0�u�:6���)1�LjC�e����+k�oY�ym[���o\"q��1G�x���oY�ym[�/m{��i�Qa	�!m�����mʄ}�DD˜ݤ���}�z�I!1
a�I�ym[�/mz��� ����:�ME �DUSp���t��z���k�@u�*����8�'昇�x��!���9��%���X�C'D+�7ju�Y��N������g1� ��h��F�9�s�AW}��=���񐐙$Л���;\���"."(�7J>n�����ՖH��A�1�G&�}��h��鸗��� �z��jJ\�7�Hbm8�h���.����h�^�}�[ْ87�!��c����҄O����ݓ��k���<'�ˆ{�6{OnrƮ1�ꫥ���m&�ۘN�Oe��[��k�@?7J>n�!Hvs ?w���
�l��rK$�َ��UTrds�������<����r9'��(��<��6�hw�=��^��l��f�6��uP1�.����Cx��ĬV%��`7 d�Zr��%?$4i>O@�0jiG!��$�9 d*�P�M-,���Ʌ�@�=��k0��d�GF�*H��P\|y��~��v&�`A��I ��(Y�pJ8��d�g$�t0�ې����!�TdL,�T������L���>M�$6�ʎ d>D� L�)(�Ȣ���B�A�#��ǨT��PW�P�(qG���,8l�>�Qz5��DW�*�<��s'�8���v/��?.�l�,�c"4�8�/�f�$��l�"w��Ş�P����zo��!�0�G�9.�	'��/BG{��Y�Kw]�~Y�����
^�|Pi�xȍ�S@�N��F��Y�7��a�:�4�4���<�W���ݬ@`LH[P6Trs�*�>�yزO*�Pǹ����f�P�/
�T��o���@PY�I_�N4�jB-��qnk� +�@�VI��Y'{��ms�Q�ll܊	��FH쟂���O)f��w��ŝ,[�쓛���B����&�׬߱#��繠y�_}�nM)�~��2��~8u^(�v��/�I��D��ɊG$�OV�v��9�[Ȏ�ombg1Ձ��w������|��[���]s^��N��bn.�z�d:�V���sP�=�[���/GV�$�ٛ8I9����[�׹�z��!4���'ߍ�_�����$sse�w�����s]������a��I�ےY$����I��g_
os_	'�͗�($tc�5�qc-�I�+{��8IŹ���P���3e�Nnl�*����RSIND�jB-���@�s]�z���W'76\� ��}���|!TB�DA3D(+j(x�C�1�BXƀh 1�D�]-�'[qrb�a�̜m]�\���s���Y��Q��}�z�.<C�#Ø�^^�O�䈕]�h����n���wTX���r�hë� ΢qN��1�������������9��&7gh�p���ͭ�d��)�fJ{nڗ<]:�تp^v籸0 �j��;u�+������Q�.D[�=�����@�M��,6�$� ���!�HZƮx�G����[��xu�Ί˷ks�t���h���v4���t�ә��5N��P^}���'76h�Nw5���~�{�쓛���B��NE#�;ڠ�/^���Q��:��v9��i��DJHa�$RK�I�k�d�[��W=]�vO%��,���EB�q�Kp!p^�G�$�w5�qs��A�W����=]�u����F�����:@~s�����=�K�H�aD�,f��l�8,hbO ��L�I�n�2u��xnn�X��]����6��n�����@����J���"9�s��������"I��F4(��;�w5���P`�����_��jI��}�O~̗��Sg{�)��"l5!	��@vu� =>�H�DL�7m ��(@\����'�poI������f���{�+��mY���<�ȢnI�z��k��9^�@<�@=8��J�#�����Nb�"�h�'�6�<t�q��k\箇��q1�ғ��R9&�}��h�W�wY�z�˝u
G �As4���s�x� ��(@v}�S�8�#NL�ǠwY�z�<�*0`t��$�1زN/��x=�		��I��$й�W�h�^���z�u��e,�$�D#*I��@?7J�^�@<�� ǎY'h`�7d	�!N�n�e"a�U������粯]<�fv/X��mRl46� ���g�U�����h^�@���4�ܭ��'F�d����mH+�4�s@�z���5�G�8܊&���4�s@�^�@<�@�z�#���RI"��P���t�;��ǹs9�s(����$�Fe�j8�%���,�%���c��?c��t���G?��n߼���T�8b�kl�a�G;�mNnΙ^��y�)���,�H���~ {o�@:���׹�r�^��{�^2#��CnI�z��k��9^�@<�@�̥rn!��
94�s@�z�7?$y�f�_z��jJPND�� ���f�����h<ݠ���uJ�\"q�oI�y�f�����>�z5$���Ƥ�o��E@�XU	,�@F��J�Bվ�����w{߃��qJ�U\Xj��(�6���sy��-��,Jv�9�d���B�;Jݮ�u�����Iv,�����w>�_v׮�v7`��N�<�=�u��pn�b|2G�%{��;�f�#۷�s&�yRhN,�/�5M%��O;	sN������y:�藵�[8̘.ٱv�
���9xu��ƹg����]t�����]�V�G!�{��ƀ��鉌}�������`�)Į�2��)���^n�k���8���"ݗ���ő�N7"��' _��}��hO�;��P��I�3e�{��n cH�䑹4�s~��H������4��hP�'���As4e���h<ݠ���dU9��pO#NL�ǡ�佷���h�^懿��!^�@�:ˌ����	����@�� ��(@z^:@�v�o���O��竭�����-��S��G'
ō��cl�6��әly]ۻ9T�7v�~n� =/ �;@���%() �� ���f��^��U��Fn����p�T%Ì,Shh5�3��:�O��gRN���_@�I�`X�4��#`�$v@�c�׎ѳ;��� ��$�y4�r(��h���/�����^���@�zɄx)1H�]����:ǵ�=-� �gd��ߛ�ݭ�)˞L@m=l����FK���n*R��]nv��6ߞ��ݘ'�q�n#n3Ē\w8�_'�N�B�ޯ�J�q�I/_\n���ӐF��I|����UU ik�k�K��Xv�K��|I/�L�d0F!n"��;I%����K옭�H�� hUTP�/�>q$�o1�I%���G#J2�R>q%�*�����Ԓ^?z�<I/[�ޤ��ޯ�K�����j'�A�f���ޯ�K����$����Ē�ʵ��K��C4�78jǌtZE�\[k�H� �9R��5hݎ�N��i��c���6�z^Ω�~�=o�z�J�z�<I/l�Y�$����ĒW��3I29�	8����ޯ�<�٘�^�V�RI/{��Ē=}TԒ^^��`1����8�Ē�&+f�I/=�y�I��jI/_�_�$��%^��qǆ71A��$���<�$�_U5$������m���}[�#���@i�g�޳u��m��{Lc��H�l"���9Ē?>▒K��q�%�k5$���g�$�.���	H��3�]j^}��p�m]�Z]���a��H�G&�:�˒6+�m����~ߞ$��U�ԒK�m�{�I��jI.���D�pC!j%#�K옭�� �I}���$���R�I|��>sh6�f�����&�ۊ3i$��ݜ�I�qKKj�@H�s_8�]٪ٴ�\`X�bB��DrNq%�^��/|���Ǜ��$��1[6��@��ݜ�I-æ�!	 �F�E'��Kﻓ�I- woW�I%�wg8�G��R�I]!���) �#Uk
��y�@�":�B�� ��.K�6Cp�3hc9�$6��3Q
�;���Υ����> $B)�||���#��rp! a##$d�(� 4�V)�n �mBp�d�&H��b�!A�!�p�R8s���N���R��H@$,�a���$G2@���%�-\��2�Б ��c,"���"HH�X�:W	�����cF�v$�
bࡀ1����1��8L�B0�1��	��A����6�7��R�!�m6	�$��bB�H�j�pА�Fw�n��Č�l%�FL�}4HEa��U�� _�B|�86!�D�͠g�c�#�.���U�0�B }�3G7$\�C�$�!�!���#�x�#	#?��w�w�~�Z�L�p �$        9,�� 6�       �6݆�M�Ή�`�b�!)C��kn����!�<����SĪ�\
��n���j;a��̥؁D�n+9,�=��qڕX����Uj��P��J6[" n�d����*��j�6b�*�:���I���ӵ���:kK;JCB�]�����J�/'��}�]�ٰ��y3����m���<nס{9t>! �[m�PWl	=n�n�9�.�h�*l㚁�y�+��X�YM�h�Y�&N����;�J����n5I�=���W6�m�vYn��rr��Ҹ�6����'<���;Ɨ�q2ԵA�=�+�x�9"2�l¤]����� ��Ȏ��q�]D��m`�5ɮ�zA˗�uώJ)���*�ˣnݪ�XW���Ia���e	N��t�f	�ճ��H���4EBr���Ma9@n
N��Er����WK�r���F�SU��.s�g8���as�XP�b�ٶ��ˇV^�Qa�S�Mˌ�[�N�Q�X�gY7.�J�����I:�T��Ld-[K��qrzx���v�G:��&a9�ȇ[�����v�sۏN�Nz޷e�Q�tM�G]�C�x��S۷e+�ٹ�#����D�m�1��ZڅIIo����O�����fƍv�����1vͻd�8�t� 46dR�Tjx�irjB`�Q.Q^[\�H����=a:�R^�-�upQ-U;���|@t���bb�#u/-Պ��r��z7NaP#b�^ݥf��vE�Z�/ YG)��d�)0UG����ȆB�SKƃ"Ʒa�Z7POg�vc���<���Zǘ��R���H,n]N�Xv:0�;c��{S]����t�M:6��ō�m��R��<]�Z�mKl}�����7b�n�X�͞��)��r��+� �n�d��I������۔�Ӝ�MU6VV�Jqmam-�4gF��78Ćd&q�fs�A\����%T2�J�)�p�0I�x�C����șy���{v� KX ݬ��08���f�V�[el�2�D�ϱ�L�iإo[��+.6q�#��yN9�ۍ.6����8x���w8q�vkl��j����f4a:�\x��td��9���bm������5��X�k�c�7Zκ����`�ː��}ێ;㾍^��@�Z���\ԗ��v��B�Ѻud�k�c���$�����]s�W0\-)(\4�qȠ�( ,
���� o��Wkp�����}mJ:�XxvV�<16���R4�u��ir�s�$��Vϖ�RI/}�o�$�}cԒK�'8�_cK.(�q�nji$��fNs�(~����K���8�_YV�RI{eX�I1B7�NDܞx�G��R�I/�̜�� So�5[6�Iw���I/�Ł���N�KIx6����$�vj�m$�����$�����^�j�Ī�XI�$��U�ԑ]�fM�|�K�6;I%��c�K�N�c����8ό̀M�TY�XY܋����ݙ�e	g���0��g�ƕ�;I$���9Ē_>�v�K��ǿ|�]תô�_�[�bF�0Yr>q$���s�h��@4��R�
���[���$�u��$�_{��ڠ�Gp���$�9r"���I/��q$�Ǌô�����|�I.���$�>�>#l� e�!���$��f�i$��k�I|���Kޓ��y�%�iz�'`���v�K����$������K绯�I/���$�{�ep��W��>�=��ۊ���R�g8{k���0f��Kڸcv��]o�_~Ať�����$��͎�Iq�c�K�x�?
���C�i&�|�Ē�����`�D�1�#��K��9���z�;I%�3_8�K�܎� H����^�6��D�&�m����F5m���;������D����)}���K}�9Ē�q+�c�6�(ۊi/U
 W�����Ic����K>̜�K)��
$�����FčG<�~x�Iw7Ivf?t�Ē���z�K�u~x�]]I옱�%��e!�<��ۅ��b{s���C��C�{4���յۙ��mWт�� �~~~_��Iuun=I%Ϻ�<I%�=I%�[�J191H���K��q�ʹ��_8�K�v;I$����ڦ��km��qHa�ji$��k�I|�#��P�H�{��I,תô�_vbe�M�ca��fH�Ė�S}���I%��9ĕ�qۣ����%(V� �R�F�`����P8(��������%��S�H`�7����Y���I-�U�5p>$�ݛ��I%�̎�Iw�aE�6��bf���x���<�n/+tU�Rw(���ک},�Z��޺w���Аh$��RJ��[�RI[-^x�K�l{@`��I-���I.椥� ����@ۊi$�&b�<��c����K���8�]Ǌýi|0j�H�1��1�ˑ�$��c��K��9ŠSo5��$�v���$��]i�#��	I���n��K5��$�_{��I%�=I%�[�J191��9<�$�+�IxCx owϽI%�ގ�I.fd�K� �@�o!Zd:_7$�A��  ۙyrۺM�:w\��i<6�^�i�Vy��Kj�t��c���c���s�'��a�Ss���|}�_�}�J.zީ��9�\��u�j�)�Q<�ڜ��r��1��k�l��q�ڛ�b�nY�^�7�&�\nD�YS2��s#=c�9��m����&#W��7W\�yT�ѕ9�F�5k�vbL���eCb��V��wL]m��L�D�*��P�-I"Rwe9�V^�[�6��L�y������˱H�!թt�s��{�ྉ�j��7J�?����_8�K���\���W�W{[��a�I,����I�da����Ē_<���M��ۻ9Ē�z�;I%����< ����"��n#r;I$����$�q��-�X*H�f�q$�^�v�KC�dq���Z&I9Ė�͚����ߟ�$�����^[g�$��RRҐDb0�M���]}�>q$�@W�_��$�}�Nq$���i$��Hw%�-cW<r9��ᠴ�Dְ]�$�[��h�Ÿۆ�Ļ�o�=I6����$��ݎ�I.fd�K��X}�6�o��<I.V����dr<r!)#ԒW}�s��*�a "S
[y�v�v�Kf>q$��2;� (Pm����JH�.@�H���I,תô�]}�?<I%�=I$���<I.�*�D'	0ǎdm��RIs��Iz�RB^\��v���=��y�'W���I�da��quWH������d��@�Nv�=��aD�&e��Ə��&=���n^K�8uщsqi]ͅ�,{��|Q�u�Pyn"6��߾�h��^�˺���'��d��l:�1��&I,��_V;��@SgVo��{��VI<��(RG��JjR	*#)���N.��ԓc���4#�2��)�_pV
UB����K$�^�vI���2FčG	�d��� �ݛ��'�͖I�����ª�{3|쓫�!��d�8�r"���'�ܖIڪܘ�𒮿=�]�@=8��J��M�ͧ�n�:c��[n/c���q�t�4�ї��p<^��J1��&!��'&�˹٠r���'�<ŠUq~��d��X޸�p�a��nK$�}�w���{��'�͖I��^K��ί/�R&�)�N4:��@x���N�>�HK�L&)��E��}^��},��w��'/��5'��Y*ҭA2�E
��}T(P�1��VI�)"I�ˍ$I&�˹٠r���<�ڴ��,��( �ۻ L9
qڢ�A(�'��ֶ�5]�tFx�=�u͝����]i�E PS""&1��W_���ՠ^�@����<�ʥ�����G�$�@��t�:����v���:@d�C�D�#�D���/Y�Uy٧٘�V��__���[�&��)1���94
�;4]������٠u|ۮ$�$�9�F��9wW�z�W�[f�U�f��g���t�F� 5� 	�M����w7nհ���w}�W��6�O��a�ʨ�!6������v�vnF�6���=���۫�=�ʀ��ݗ�'c6�a���u���!�ԯE�D���3[�zs��򝛤��ͭ�0-�^�Gfέҏb�s��^.����D�$#�a�+u�%i8c��+����N請p��j��g�먅�6�H5�H"衃)P��$?���S<�x���ݗN�4�qجYv�Bݘd���3�a2)@��������ݠ����-� 2u�"�y�rh�ٿbG����V����h\�X=�'H�M����uz|��_��{��MΩ(U&4DL"�ӎM�uz�;��'��,��@x?Ok��OF�)�5&0Yr;$���,��/�vp��q�OW{��> �a�,��5P(���	%{\Cҿ۫}���֌&�HMv8�f�j�e=I�e9QB�"G'ē�{��8�;4]���� ;���:����j$���1��N,��xA��UP� S�B��n�db����0B H#�XE©�� �&��]��UU��_��$���d��̗� :���'�C�rY'f�$���,���z��P��ޖI���K�Tu�ԉCxLmǠ޳@:۴����9�s�齤N�����D��I�fK$�
Z���ߞ�{z� ��j��!���rܾ�N�8I��ܫv}Va8:�{.��ؠ)Xp�]ē��I$�'V��d2s <w�s����9�P��Z7��&4&Li�&�˺� ���y���8��%��T���}=bI��2Gd���K$�grYc�!����\E��RH�	�HAbakb��!"1����HJ�H2&l��c���֋�!�L����F�	0b����ʣ�t0�P ĢaLK�1B1�
�Z+�P����@��#%�0"I�V$aFB�
G	5� @bO�W	CJ�j�ā��G&X� F9 2���"�v��6�����r��@�9Px�6�S�9���҇Q*����*8G����6*qC���3�o=��RM]�vI?a�2����l���O��6u��'�� {��1�7T��)?4��'&�Ws�@��W�����,�y��d�UV`ӧ���@��,燗n�8�7�l\����,��n�+q;V��`��"��I8d��p%��N��; {z� ���fx���M�����Ԋ?�<&4��oY�^�@��@��W�~�����@�A�pn IɠOۛ,��:�Y� � ެ�;$���Y'�;�q%#E��l�%���q�@9Ǵ���t��";��*�x��l���L�4��=_w�v���5����^S��Ȉ��B�7vV��d�������2�hB����-!�J3��-ڦЄ�
b�����I@Qr?�8��R �n�^S��G; 彤�l�M���7��@<��������d��w�
��sf��q����1��N�ǲ�=]�;;T(%�{��'�ݖI�s&Rp�D1!J'%���DV��Ԁݯ���ݠ�h�,�a&�Q�S0F�Oz��}B�@ ���'�W�,����M�@*��
�"�m�EN-Aq��D`P=}=��^���ēm���l �vl�G<��5�ht2D,�Z�p�[�}�2K�n3G*��.��}n��7v���8H޵��O]��S�/:��kW<�sv}��f���m����C��\�`������v�]��<��\.
��U�V�j]�rrp][���w=�ax�K�\(�.\��fRyZs����K������앛�@�6^��!�Z�����U�W+����2�DBS����N��R�y�q�-�䓍d��L�#������ň"#�8ʍ��I����8�[4]���ՠyr�cؒ����l�%�qufK�B���se�s�I�ْ�U
���:�I���`1Ji�ݠǶ�̦��s�'�v�.w�y���&�$�a&�@�v��mB�Kv�b#�3����gImIq�2)�y�e�$�
Z�n� ;��@�v����iD���,@e^m��NO����B�h��bn�rfF#2��jI$ԓ��\h�)�%H8IՋvY$��rY'�y�¨W?wvŒu׬0�*Qd�R��d����v? �@�+�P&�� < ��9Ɏ?�Z�_�����*���!�1
rY'1��y��VtURZ���$��}4
��"Dǒ��qh\�2"�ZX&���ʰq�n۔d}��IH��m��ŠT[f�{�@�ڴ}v���E�<i�@ό�7�Y��\��+[�:�=vN�5t�:�׿x�Ցf�ɓ������4^b�O>y�j���Gwe�~͉�$��b�M�j�<�ڴ
�l�~�K�@$N��:�r@�B6��d���z�I�;��S���0�a*9(N�C�Pp��K$���+$�2b*2�JO�< 7�Qm��f�k�4A}ٺ�����l��R�B�NK ���y���Zten��N;A����~+���5y9�����hT���k��ع���e{Wn�0��#�83IcM�uUv��;b��� �'����W̓���I՚<$H��4�(��w�ܭ�G9ɓe��@�m�v���Ǳ
D��m�-�.�@=�;F�#�ɟ=��ݔ�s%K
@b��NK'hP�Iw���9�5Y3c���j2"I��TL\����ݕJH�R<x���@���c��^������=�v�~�3N�5��x1��s�p��O.�ByC^6h3��i�cv�Hq�~���z���B�X��)�{�U]f�{�Y�u}V��̴�D����VIŋ�/�<( '3},��{�d�|���#��li�9�,BNM ���u}V��ՠUWY��ubC��"8(ے��Tl�VI��uY'.�v�	w��@��}�$Lp�4�n-�]��ml���f=�:�(����(����Q*`�@�h
�H`
�uk!�m�$�H�V� ���Ԓ���du�:��ᵶԭ�c�q�1�sH�v��W��n�-�ܖ���Z���s��bN�ӭ1��{s��m�,�U�Ob��|����C\���骞ίa1�=�zmS�W��D����#T�ÔLJj`�6�/[��]�ļ�d����\F���6�T�vmvì;��m�-�1k��hof�zX7'g� ����O��
i2���X��<��&������V�tn�'��R��+�Z��AX��v�R$\m�$q|I�~^�,��޳@����]�@�U�PY2��rY$��r_����=�Oq���8�w%�#�`�4��R0�`�$��{(����8� {�� w�&��72@SR+'Wݛ��:�f�$���;'�(Uy�|���{֒l��p�����*���=^�zW�hz��}Aié��H���[a�\Dȶ��j;i������IN��ab�6��\�8���������$��
���@����]��B�z�d�yo��}���2F�.B-�1�js��n���?�R �W��u��@v}/m��:_D����3�A!q�7��?�ZUu�%˯�@�;��<�.U�Z�6��Z�ke�2q� 1�9@w�ܠ1�;�XJ@b���rY'��q�'�U@f������UWY�x�K:ɋ�D�1��z^���n�ͺ�!
j6z0�t��lM��t�WfG��#�'Ww]�y�h�����W�uYSJI��	&�=�]�~���W�r��М_f;�#��i&h�m�	n+2r���ԓ��;�J��H�$I*�P&;y�cRM����I���;�Dى�hI�d� _s]�unk�O>y���=Y��;�f���6	r�������s���g�9�{hO�^�\=��� G�4#����]*ΐm��;�������CwP�Ag߾�w������@�F�dM�����r���=^�zW��<�-�G$�8�O$qY'�r_�ꪠ8�|����O>v���0eœ&Dcq94W�Z��H��r93��@9�{h�!ͳ#�H�����;T(
Z�5�'�۩'/o;�I�!"�E�Gx( ��^[�IϱM) n(d���vI��1Y'¨z�UP<���Oq���;޳@8�6$�c�����2,���k�l2�up7Ep�oV%� ]�v�kֆH؜1��@���hz�Z��M UUq޼�d�Z��e6br��RrY'�>�
��M����I�=�N/�r_�Gtn�#`�!��H��;��(�#�ɝ�������@<x���)9,�K����:�^���t��DD�Ƕ��F�LR*��8�O$qhz����W��Y�M����I���8�է�e��M@��5�.U8�M.���%�!��"� @`�� H	�d�A��*4*�h���i7��r����Ybl���,��*��"1zPZ��*���4I�#�r8�`E @�e
[8O�VA�>'Bh��L3ns!����m�5�I��8!Ā       M�         ����;n��KK�O;*c�+j�1���]�,�Is#	�F��Pږ��\kqlݰ$���[�b���D\�:8Ƴd�uq*�T��p$�T����&��N��kc��T�Cӽ,�'/7IWi��sYͪ�¯�DF1�U��sԫʍ��ul(�cmΔUC�`Sgi�qnM�c:솀l;=9�Yg��v{l籔�[VS�x��D,u�$y�ӎ-=S����+;.�B�v��5��SP�8���miA�vABc��jw�Lf�@r�7g�Ǔ`wZ.�ʃ����m�.��*X��V-�(n�cT.�v��29��\P�3�������J��3Jd��|�E<�Y�
BN�\�F�!�"�S���p��nȥV�=�;\G&�uͶ��\�:�����I��%��S���5*,��&�V�.�q�k�F��t���p$#�sZ���3[��smA���큶���s���!S�;p ��v��K���k��Am4�Bv凛CJ��+l�d��v� �@��nv�W�����K1�P�˝���Ɩ3��E�Σ��l��-�F�b6ܮ�v�j���6玀��=��2���t���W,��X�K��D��YRvo�C��̲T�\q�W3�n7Y@�]S��l.��dƬ�2���;�Y�.�v�2MR�q6��9N�,[j_]�l��p��z�uSr��g�7F�����yÆ��euM�؀K�!��j�*�xi䧋�AZ��,K ;�3IA�U�W���c�$��+�tVM�54g�ۛv�`{E�v��t���Q����&���v�Z콵�J��s�b��)��	�W=�z����1p��vYt<)�ZŬ�k� ㅝ�v@����v6���TF�v�5����D&�BM��q��a�7KF�{A�$�9.0l6�$��83s�H�8Źr\�3ha~7�Ȫ�G�a
�A�u���>t��:@U����4"�?+:v�l -� ښe\��m�n�L4�$$�B�:����ゅ��<��wc���p��y�)1�u�7+S���B��.θ�k������E��-Щ�βm\��b�J�&7c�����m>�6�K������ӕN�3�����.�Z�-�u��5	Ԧ#qc�gg�&�;c����GW]�[x�Ȳ6�5i�+v�X���6A����w�����~��b�*�	�M	���r�vy�	���an��ft�0��(����"�l!Q�NN�o�@�wW�y�}��g�*�~���|�Ď5#Ǎ����<��Hz��O��=>n��!��I��$�n=����9z����@�wW�[�Sm�ؤ��ăb%яm�����t�c��{����_�h���`���=^����}v���Y�U@�+�5�~�������׷.�u�b���ّ� d�-��tS���,Ihd��\�%�����$��ܠ2Oc����8���|��/�%�q�'�c���tj��uPu�J��*�B�BBї�d�[�vI����n|�c���6,�ŠTu�h���P	|�5�'�{��<�# h`BQ�NK'�T.��$��5�'�<�d� ��f�$�X5m�jFld�@vs 7��ݞ��%�=>�H7�ߛ��/�$DB�L*�%n�[���Z��X:��^�#����#������)x!SUt�啕@d�q���u�G��2w|���{�M�#*Jl1I�t8h"�%��r���n�8���'q�߱��Kı9�{�4��bX�'9�z�6Eh#A�c�
b$�D���7ı,Nc��4��bX�'��}�&�X��ܬ��F�lE�5P�*���tVE@����L�����I��%�bw��gI��%�e�;�
2F�.B��t8h#A��}����n%�bX��}��Kı;�^�:Mı,K�罍&�X�"47f��Ci-�AN;��Aб9���I��%�b��/}�&�X�%��s�Ɠq,K��ﱤ�K�q�����(~�FmzNn^c<t��*�e�vD�S��Z�pꮣ��O^@yv9�2Q��q]�F�41�fˡ�A�,Nc��4��bX�'��}�.�X�%��g޺Mı,K��{F,�,�!���C��4����TX�%��;�cI��%�bs����q,K��9{��7�b�"X���RFld��p�F�4�׻�tn%�bX��}��K �,N㗾Γq,K��9�cI��%�b}�Sɤ�\�&&�4����̿~�Mı,K�����7ı,Nc��4��bX��)  D�P�D@�xJ<� ���G�����&�X�%��g���L�2'm��N+��A�F�>��t8hX�%��s�Ɠq,K��ﱤ�Kı9���I��%�b~A������8�C��B�{n�y���*R��ݖV�z#���s۷~��d����7����t�D�,K�����n%�bX�c��4��bX�'9�z�7ı,N�6]�F�43t�(���!'�gMı,K�w�Ɠp��1��s���n%�bX��o�gI��%�bs����Kı=���	��ɜ\g�Ɠq,K��3�]&�X�%��r���n%���bs����Kı>�{�i7ı,N󦽙0g9��"P8[��p�F�4���6]%�bs����Kı>�{�i7İlNs>��n%�bX�vC�0�Р��	��4��hu�u�n%�bX�c��4��bX�'9�z�7ı,N㗾Γq,KĂ��=ӝ�˽��c�t�k�-`
�(N�\�W�p���{"D���C Fz�DVC�h�.ٛ�۠{^���y�:�/s�;Omxw�l'[�:�=ӳ���n4��u�m�]�`f�]3i���Z�9P�t���۝<V���C]�����D��kn-��S�/.��n-��ĒΊ�8�L�����fs��直s\^�t��n�vd�k�t~���z��w!���>��s�[%����i��-ά�"[��X�����u���u���-�$a��FH��F�47���7ı,Ns>��n%�bX��/}�� ��D�K��;��4��b#A� |�L�E���p�F��bs����p��1��;}�:Mı,K�����n%�bX��}�&�~B*����b~�?k�͙�d�ˌ`�%���n%�bX�����t��bX�'1�{Mı�ű;��)�$�s�����I���	LK���\e5�T}�罍&�X�%�����n%�bX��}��Kı=�_{:MĲ�4���W	FH�%�BQ��Rı;��zMı,K^s>��n%�bX��/��&�X�%��s�Ɠq�F�4;�u��"��%@�6L�M���#�lK�mѱ2�gz�>�ng�Z�pܽ���fc���:Mı,K�Ͻt��bX�'���gI��%�bs������1ı=�~ޓq,K��|k�dbH��Ep��᠍h#C_V��8;b�2&bX�罳I��%�b_��gI��%�bs����pP�F��H�!�A�"�ɤ�Kı/=�gI��%�b^��Γq,K��3�]&�X�%��r���p�F�4��6��0�`��Γq,KlK����n%�bX��}��Kı=�_{:Mı,K�se�᠍h#C��54�k�ᄕq��7ı,N�=��n%�bX��r���n%�bX��w��n%�bX���.�h#A��j4\�
IE�͝����/��C�Ֆ3����x���lNi6�a�s\�zpQ����oq��O����:Mı,K���:Mı,K���t���%�bw�צ�q,K(#C^,{LF���q��C��4K���:M���"b%�}�~Γq,K��s���n%�bX��/��&�~Eb����b~�����9�0I�d���s��Kı/����n%�bX�s>��n%���Ȓj���A�D�
��bj'�n��n%�bX��~��&�X�%��w^3��!�8�nK��A�Avn�Mı,K������Kı/9�gI��%�����{߳��Kı;��%�".@b��WC��4��|��t��bX�
�y��:Mı,K���t��bX�'�Ͻt��bX����I'J0��(F���B$�mV⧊��h�[�u�-��i9xq�ŷO&�]�e�3q��7ı,K�w��n%�bX��ﳤ�Kı>�}�Aı,K������Kı:���Lc7*H l���p�F�4��3e���8���';�߮�q,K����߳��Kı/9�gI�")bX�#��54�k�ᄔ��C��4��s>��n%�bX��/��&�X�%�y��:Mı,K���t��bX�Pћz�FFT����WC��4 lOc��Γq,Kļ�}�&�X�%�{��:Mı,�I��8D2	���ȏ�'����I��%������I���."���p�F�4X��ﳤ�Kİo{�gI��%�b}���I��%�b{��t��eh#C����\&8����E����͙C7[˶��u��OLK�k�jn���(�-��NK��A�F��͗C��ı>�}��Kı=�_{:wı,K�w��n%�bX��u�9HAӌ&�4��h}ٺ�7ı,Oc��Γq,Kļ�}�&�X�%�{��:M���1����~��$E�LP ۊ�p�F����{���Kı/9�gI��?����{�߳��Kı9���t���h#C�$e�PР����)bX�ؗ�w��n%�bX������Kı>�{��K���O���K��A�F��_�n(�@�/�t��bX�%�=��7ı,? �Nw^�t�D�,K�=�~Γq,KĿs�Γq,K���EH��c�e5=�W4�1�g9�KX ݬ���GN���n���=�추�v�y�l�g�R캶L��)qv��b�o/�c��l���i3�[�q簝���ѻYs���7T�ڱ9�&��٨��]K���p6y�p�[�$C=�;F;L�[nӝ���=A��q���4n����." 'm�I;�6v�r�c�_/Om��λ�%\��1sƃ]Ʈ�6��đ��P�.��+��(5(-�j����מ���N�8�Y�ŝ\#�."zs&�Y�Pi��R&\0����8h#A�͝�t��bX�'���gI��%�b_��g@�X�%�{��:Mı,K�6���))�#QH��h#A=�^�:M���1ļ�gI��%�b_w߳��Kı>�{�����x��	1r��R�]�bX��w��n%�bX��ﳤ�Kı>�{��Kı=�^�:MĲ�4��ӫ�\QӁ�ܗC��)bX��ﳤ�Kı>�{��Kı=�^�:Mı,D�/�ﳤ�B4��ݽ$$�i�r]�,K�g��Mı,K��ﳤ�Kı/�ﳤ�Kı/y�gI��%�b{������f�2Lb`�!,ܗ��[,N����i:7H���ک}���đ�&@Cn+��A�F����t��bX�%���t��bX�%�;��7ı,O����7ı,O� �h�FMZ�It8h#A�_s�Γp�>���b �DG��`�D�K�?{:Mı,K��}t��bX�'���gI���1S�����-����%�᠍h�/���t��bX�'��}t��`�b{��t��bX�%���t��b#A�CSI�.II�t8h#Bı>�{��Kı=���:Mı,K���:Mı,�11����8h#A���d�Ґ"ۍ�"��Kı=���:Mı,K¢�;���}ı,K����&�X�"4>��WC��4��d��e�R%$��ń1��W�M��\��m]N6]��:+�/i�#s���%��7��*�����x�,O����7ı,K�{��n%�bX�s=��~R},K�=}�7C��4��{G�(���
8���bX�%�=��7�@q,Nw>�t��bX�'�z��t��bX�P��5]�F�47v�H��\�f��t��bX�'��}t��bX�'���gI��4\�u�ކ((dS���.uJL���k��FLĩ�B0c D�D�>��nA�(��|�'c�~@ر�j����!!��� ����������ԙI��3�apd���M0�i:)�s��0�I��	�L��=��	!"@�!hB�G#2<Rl���$d�s�����2.��)(���A��)��^y8T �r��U�bτ �P4�! �ªpp ����pDv� Q:��17ιt��bSAs6]�F�4;���$��d��Lc�Mı,�$C?g�߳��Kı9����n%�bX������Kı>�{��Kı9��jJMZ�It8h#A���5]�bX��	�w���>�bX�';�~�Mı,K��ﳤ�KĻ�������q�Xـ�L�;���aؒ^�n�U��&�z�ح���F	7O����5-Ɍc�n�q,KĽ罝&�X�%��3�]&�X�%��v����bX�'��}t��bX�';�z�۹�b&d����p�F�4��fj�#Ʊ,O�����7ı,Nw>�t��bX�%�=��7 �,K���ܸ�(���qH��h#A�^ˡȖ%�b}���I��%�b^{�Γq,K���ﮓq,K��9{�zD�Iʈm�t8h#A)vf��q,Kļ���&�X�%��3�]&�X��WdD���
/t@����Nc�1�:Mı,K��uq�� �p ���p�F�4��=�i7ı,O����7ı,N�ǳ��Kı>�{��Kı?B���p��3�a1��D��$(ZG���]u����v]r�^�p\��+�,{��}}�Wn� �!n(\��|h#A��M�4,K��;�{:Mı,K�g��Mı,K�ｍ&�X�%��x׳&ȋb !��᠍h#Ck�t9�,K�g��Mı,K�ｍ&�X�%��3�]&�X�%�}�;1�uD�(�mG%�᠍h#C���i��%�bw����KlK�g��Mı,K����7ı,N�6���R��܊�p�F�> Q��}��4��bX�';�~�Mı,K����7ıQ�>�{��K�����������q��Q,O����7ı,N�ǳ��Kı>�{��Kı;����n%�bX�̄�Ă��P	���v���-�л��UWR� ͙ˬΒ��v���3�
�O\�"�i�}�9bĻP�K�'i�ֶ�,�;z�5��c��'�n��Mq����q�ɷ�:k�P��5��se�:���tM��³�'��H�Uv��{OMɨb4�Pgsi� �p��,x�M��۶��ke4;�U�����-���gv�+�-���#����\θ���x���x�{���}����w>]��6Vյʮ�U�WtP��������Wb�z�{���_��2dj@�n7��a��h#C_|�-7ı,O����7ı,N��4��bX�'��}t��bX�'q��cILD���qܗC��4���3V�q,K��;�cI��%�b}���I��%�bw�=�&�~*��A����yq�� �p ���p�Q,K�����n%�bX�s=��n%��"b'�����&�X�%���߮���4��̽$-����bX�%��3�]&�X�%��w��t��bX�'��}t��bX�'q���p�F�4���1$E���c7I��%�bw�=�&�X�%�
}���I��%�bw����K�#C���t8h#A�CsvD�2��� �+s>[۪
�wF�����9��J�wU�E��������)5�����K��9�cI��%�bw����Kı>�}��>���%��{�?gH᠍h#Ck���n"S$�wF�X�%��w�Ɠp�A! �AhQ��E e�,K�Ͻt��bX�'�����n%�bX��;�i4��h}�CSIF�qA	I��7ı,O��z�7ı,N�ǳ��K,K��}�&�X�%��w��h#Ank�L����3t��bX�'q�c��n%�bX��;�i7ı,N��4��bX���&�4��hc����JJ��1��7ı,Nc��4��bX��>Ͽ~Ɠ�%�bs����7ı,N�ǳ��Kı=�I=-�n)L��!�lmm�vۗN��C=l�Nّ� d��=�<LmۃDv3�[������{�K�ｍ&�X�%��3�]&�X�%�y�{:���K��9�cI��PF�43�z$H.[�#�4K������q,Kļ���&�X�%��s�Ɠq,K��;�cI���F�4;���$�� ��q]%�b^{�Γq,K��3�]&�X��1�0@#L��N�>�4��bX�';���7ı,K�Iٌ{6ܶ�14Q�K��A�F�{3U�ᠢX�'q�{Mı,K�{�Ɠq,K�31�߿gI��%�bq���jd�jEt8h#A�Ǜ��n%�bX~#����O�X�%�{����7ı,O��zi7ı,O�=�۾���	�Wpʩ���>v���:_��ֶ3mf`;[Vn��T��GBRCfKq����Kı;�߿�i7ı,K�{��n%�bX�w���n%�bSCn���A�F�ٺ�S&B�dG���4��bX�%���7�,K��^�Mı,K�ｍ&�X�%��;�cI����*b%��v��?�3.r�9��s��Kı9�k��n%�bX��{�i7ű,O���Mı,K��{:Mı,K����%���,�2Yns4��bX�'q��Mı,K�w�Ɠq,KĿ{�Γq,K����dDdQ�DB� |�؁�D�=��I��PF�43�F�D�����-�t8h(�%��{��7ı,����7ı,O��zi7ı,N��4��eh#C� g�K�(��Th$lV9��ڹ9��2�э����s��m]���g��U�$��"L0c���h#Aw���)bX�'��4��bX�'q��ʩ蘉bX���oI��%�b_�'ſ�m@Ld�$�C��4����zi7ı,N��4��bX�'�﷤�Kı/�����H-�H�<=�Y�����2��H'o{�hI�7�w)�$���{��n%�bX�f^���A�F���54�n'�q��I��%�b}��zMı,K��{:Mı,K��^�Mı,�c��t8h#A��7_
`�T����1��I��%�b_��gI��%�b}���I��%�bwﱤ�Kı>�}�&�X�%�� ��1s��~�u��� l ��tvMջu�*�og[�-��Wi.�r���l�q<Q�)���ثp�M^�p�����`l��n���eQ�5���u����͞�3J$k��f����ɰ����]��gN�{�qK��vź vSEͷa����OS�[9�q�n6}k����6���=bۜ���l�:mW�K�ï7Z��D�N�9���;ߧ���L�#�rnL��}��Z�y�n3�h��p�K��0Y�ƻ����m����%���X�GL�Γ�,K�ｯM&�X�%��w�Ɠq,K��ﱤ�KĲ��we�᠍h#Cs� QqDn[��&�X�%��w�Ɠq,K��ﱤ�Kı/�����KĲ�ٗ��p�h#A�Ѱ!$�#X�2Lc8�n%�bX�c��4��bX�%���t��c�@!����{_��q,K��=���n%�bX��M{2`�sqpfL��.s�&�X�~`���~��:Mı,K���M&�X�%��w�Ɠq,K��ﱤ�Kı/�װ0�jE$�4��h}��M&�X�%��w�Ɠq,K��ﱤ�Kı/�����Kı>�ߛw����V<ln���Й������í�p=e�8�,�X�L�[|�����ga�f��Mı,K��}�&�X�%��;�cI��%�b_��gI��%�b>̽7C��4����kh��L�$���q��Kı>�{�i7C�L��uı/}����Kı9���I��%�bwﱤ�Kı>ｎ�����n;��A�F��ws��Kı>�u��K�D�Oc���&�X�%��{߱��Kı:�jzJLD���q�%�᠍@���צ�q,K��;�cI��%�b}���I��%�b_��gI��%�bna�4b%E�JCt8h#A��w�Ɠq,K���9�{��}ı,K�߿gI��%�b}���I��%4���[ipER#-��`��/f"-���Ļ�h��ͼj�y�M�Y��a.[��wC��4���f���Bı,K����7ı,O��zi7ı,N��4��bX�'��^̘3��b ��᠍h#Cw]��ؖ%��{�4��bX�'1��Mı,K��}t��bX�%��=�x��jd%�#�4��howx.��X�%��{�Ɠq,g�ϔ�T���m�A�,P�\��=IWp$�B��j�? u�>������q,K��9���n%�eh}]z
fd��At8h#A¤D�{�4��bX�'�g߮�q,K��9�cI��%�b{���&���h|7:��8�a�ӑ��,K��}t��bX�����߳��%�bX�����&�X�%�Ǚ��p�F�4���xڍ)D���ȼ��/6:�7`ܽ�nXM��F�3�fl����n��ՊwK*1�������d�{�Γq,K��=�Mı,K��}�(��%�bX��{��K��;oQI����6��C��4,K���i7ı,N��4��bX�'����7ı,K����7�4�h#Cۧ�h�J �p&���p��bX�ǽ�Mı,K��}t��` !bX��{��n%�bX���t8h#A��f����q@^3�&�X�%��羺Mı,K��{:Mı,K���i7İ#�����	PĠH+�^��0�p�UC�=���4��bX�'��k�d��lBc"�4��h/�v]�,K���i7ı,N��4��bX�'���Mı,K�=$����]c��n^{X}����u�N��:i�D붎��9A�z�-�k�,�m[��w�%�bX�罳I��%�bwﱤ�Kı=���Jn%�bX��{��p�F�4��tm�I�q��j9&�X�%��w�Ɠq,K��s�]&�X�%�~���&�X�%��{�4���bX�'������rf�8���-�s�&�X�%��羺Mı,K��{:Mı,K���i7ı,Ly��h#A���0dJDDN;���&�X�~��~��:Mı,K�~٤�Kı;����n%�bФhnL�t8h#A��;oQI���3�g��t��bX�'��l�n%�bX��{�i7ı,Ow=��n%�bX��{��n%�bX�8�a�g�f3L�xtYr4G�S�c�;�Ő>:d�uM�`� 9�T��%�h@��
$,jO�p��ˣ�kx�@�ٖ��HL��v�4����;�rU�vJ|_�� ��D�De"�����НeI�IH��eKH#��a������O�����ԃ�v@���>^߀4lAT
��\� �9�cZSf�aHH@r!�
i`���&R� �I�]�ҬfCH?W A���� �b�;�V/�[8�2�)H���,�SU�|� �V1%�:�aC�[�����@�Q��(gE�39$��d� �H �$       �"��p 6�       Ѷ�m�K�c�/-��q	*��LA��`zK��ےZѡʯd�qJ��-�5*=s�`�.���p��-����X:�m��W!u�ڼˀ�s�6+L�X�v��&�H�N�FӤnR.Cl�r�\��Ӭ�֪���ۭ��q��t��C�����m����+U�ʖ������\s	����ݶ�6�����le���u�l�x���,���J��$@�ҹ�`OXYh)��E���Ʉ�R[�J�3[5h��c���r�.k{(mVמ�(�%��4�[l�Ә%L�m��1�{cS �M���l����X���5Ԝ��J���CTRd^C�qƱ�=M��rd��.ݮM�N����)v���뀬&�#꒸�)Ɯ���������2�v3˵Y��m�a�,<��%]�q�"@$!jv���V�e88���e��X&�,q��r��Sb6�\�� �6�nڡ�	��c��T��=��Ka�k�G��p��nn�a�1`��\ D:�XMq�ͳ�la#�f�+X+�6��#�����c���m��&|��g��5On�92��@<uU,*��(%�@.��W	V�k��ѣ����Ì���y
r�޶y��Mn�U{mt�e6:�Z�cm�y#�Ƈ��S��C]@�@5U��ô#ġ�ɕ�=�86�k��U����*�uV�Mpݍ۷&����{.�8�\"��ʜAK��SB�	��iF�jc�����s��΀�@�U������qPqA�jV��� ,�D��sk%.�ٸ�P=WFSq����bL�u�����;t�v���B�b/l�"^�_:z��m&Da�6v:m�/ �P�E��/��7�2F�Y";u ��l�+�jllHUt@�������#q�[N1U���]cr3���-b���R6Z��E�H-�U�  SӐ> b&��/@@�*����F�|��DٰpA"�(���3��GU@ B�¹UB�9�|Im�$�I�!Z���ͮ���Ŝ�qv��3�nyHa{kc�7.��N�S<fw,�ɹF�N�;n�FL�P�;c���;]���{g]�QON����!vMm�6�q��7������ ��������7i�䠙mumֶ.�\v��/���lřu�ʏ@c�lT�@�ɮ=��x��F��WZ�.-�=��^#;���fr��@�Qiww7�bg8ͥy�{v�D�외���|�۷d��OLM�n�0�kO�Gnn�����"X�'1�{Mı,K��}t��bX�%���t��},K�~�t8h#A�̞���q�[��n%�bX��{��Kı/�����Kı=�{f�q,K��;�;�� �h#A�/a,GlCg7I��%�b_��gI��%�b{���&�X�%��w�Ɠq,K��fj�4��h-�F���P*g9Γq,K??w��&�X�%��{߱��Kı=���I��%���~���&�X�%�����.&nns�3���g&�q,K��;�cI��%�b{�ﮓq,KĿ{�Γq,K��=�Mı,K�rӾ�Jc�9!��i����U����{V��m�Fvx��2��w�-��w���]��`i����bX�'����7ı,K����7ı,Os�٠�蘉bX�ǽ���A�F����	� I¢NDӋI��%�b_��gI�y"D ���� `,A��P�6'"X�s��4��bX�'�s����Kı=����n %�bw�����IN0ci�t8h#A�����n%�bX��{�i7ı,Oc��4��bX�%���t��bX�'��%�#b5E�M�t8h#A�ǝ�4��bX�'���Mı,K��{:Mı,D�>�}�I��%�bs�F�D����8�-�t8h#A��ﱤ�Kı/�����Kı>�}�I��%�bwﱤ�Kı<  g�A�E6�Kd��)b�^��-�m˭�jd���$��4jl�`���׽�O�}l��m�ba�wC�A�F���t7ı,O��l�n%�bX��{�h?O�b%�bs��i7ı,K����XQ�����]�F�4>��&�X�%��w�Ɠq,K��ﱤ�Kı/�����E,K�����S1D��@�RK��A�F�<ﱤ�Kı>�{��K�gh��j`*Ѩ��y��:Mı,K(-��t8h#A�����_$8�c��4��bY��������7ı,K�߿gI��%�b_��gI��%���&"{>��i7ı,N{����P&�Q'"i�t8h#A�_n��bX�%���t��bX�%�;��7ı,N�=��n%�bX��l���H�v�e��m� m٬i-�V��futceE3pOSZ������������=���t��bX�%���t��bX�%�;��7ı,N�=��~},Jh.�.�$}�䭅�Dn� Ƕ����D��=��ݴ[j� H�h������9�5X|ݣ�G9>��1�ȷaQM��I ��f��s@=��u"�>j��1��~��N�C�ǰ��D"94-������;�S@<���;=y�LM�'cKx�����[!vh㞝�BjN[9n�I/��Ƴ�י�d�9���4=빠wt��y�d�C���vŒ~�-)�r�p��r������7h�� =�j��(6w}�8�	�TIțp�$�=�@u��G9ɜǪ�� ��y��ڒh[w4=빠w{0�: �P���Y'ۧ��Q��T�\IuW��͵�@=����m�+�"�H*G�3{�S&1�g9�r�k [�t��,�f�ؼ�i���T���U5���n���8g:�N�m�ԅ�8��݄��i��!֫���M�;n�;����ndnO��b��7�g[8�5��3Nl�^���sm��d�;f4�gd:sʹ�j��S��m�W)��v޺��r���j�#�'vٯe�����͡펝�vj;f۔�s�/4K��]�x�<�ս���8.m�O��y6��g��9�u&1X��]u̽H7u*�}'O.ER�;�<l�y�d�O32�����slY'w�K����}��m�@w�� 32؀=˔n�(50�!ɠym��<��o"9-�� {�=̆��.bs"&9��y�]���4�z���T���$�����#q�� @fe���{}ۺ��cP���w��~����#�C��˸�ҭY#(�\�nF���x�y;V��\݇��&�`�[5WuUVt���m�@w��}���}��!'�R~Q�RM����?C�Z@c���@����=�4�R׊<�E�71���ơ���}���{hn���xP�a!	nM��4�z��n�y�Y�ZvJ��4������7h��n�c��m����ȓ�@Q�f6��ncBI�s�&�#tk�J5�gTtو�2h.:�F ��(�I&��s@=���;�S@<�٠y�ܲ��NdQG&h���9Ϲ�U��Z���&jx�̍ǒc��h�)�{�i�;@�	!QR)݁�L{�ɻ���4�vbq)��(����lDDϳv�����h̶ =�)b	'����<��h���wJh��4
��5���ð<q��E�ny�)g����Pf啮	J���pLl�ڢٵh(�F*M��nO{�,̶ ��:�P��u�
�	nM��7�H=��[w4Ϻ窀H����$��"Qc��&��@u�� w������pʧP�(�Z�K'E��{�$���Y'��{5'�N5�0�)���Yԓo�e�2(�Ȣ�L�=�4��>�K$�3,Y'¶��
͉��1(� /Ä�-@c��sz��fv���ki�y��MZF�6���$����{��I����n�{�Y�wZ�SȞ
LQ:���� w������h̶-H�t��$�JJq�NK$���,�}���;�S@<�٠^�X��ȿ7W]U� ���3-��n�m��=W+�2F�zwJh�٠ym��*�@��\u��~U� � m��*��Γ�n�MU�M��I�B�6�x�= �a�8�ױ��9��g=�F���S��pKɒ�'O��DZ=H	m�L�|�c<Z���ɦ�^��1S;J�۫Ւ�L�t��uXꥦ���N����ŉ���[.���֎і.m�2���g]��m�#y˂x۞��ܴ�1�.ٶM���;��ƨ��h�����x�wE�s�VNk\/W!�]���ֱî����/%	�������(�#��w�M��9��"; ۽��*��)L"�D�h[w4
���;�S@/�f���rˉ5Ț�L�*��@fe����q�=���L���27I�0R=��4��h[w4
������2'��nFۆ�?c��#�#>��G��^�H̶ �?��M[��|�w.�aLmF�fU�ٵ��K�'E���q��vL4 �^N����m�@9�:@fe� ?c���CL�ӂ�I��q��U\vm	@ x|����Z}�O�٦�?,�vI�fX�P�I���`@�!pȓrY'3&�$�}���_n��w_��i�+oFa$4>�G'՛����@�;@fe� zV��LjaF)#�<��h���wJh/z�˙��m<�_�b���=��z{6ضx6.�m��Ƹ�D�a��)����*�X��S1����rO�͖I�e���:��y�P���nWUu˸�&�����g���ڄ�c��@
H�n�i��*DanFۆ�?,{H��!(9�B�D7�b�����`�$a(���B��"}�a2�:����&� k?\��"6:��r5�R�-%cG�%�	i�%�#�W��[H�\h�S&��� � t1xKY�� }�*T�F ���Z.�І4A�Z�5vd��>�A�q�������N�C� r�)�ӥ~@���E�)!D�R1�`{s79�f�oJh�X�iĤ��\\�����B ������r#�����=����cîNf�{�[@w1�@v|� ;�� >y��T�b�1F�e�^AK��]��ă:�x�v�:a�_S>:�bL��M��GG^�ɐ�c�$����7H�5����9�� ��h'�vy��q��JHA�$�}��� �D���B �{h�[�!�ӹ%�L	q�w]� �޳O���Ľ̚l����O+�L�������}��Ƕ��w�����u�r8��Z�υ�s	Ձ[�7H&9%��e������}^7� {�/qu�Py ���lM���7�]_߹x����,��i�I�Tͥ%{l�i6����h�UwUUg@��� ;��@�;@{2٠u,��ӉI��5#�<�w7��r&C1�1����t�9'��T��@I8!M�d����$���6v����wu�'�ݱd�,�  �!pȝU��8�����@w1�@�;@_N�������C�x���߼��:���̶ 7c�����s����,�dN�vx��[q�� kX kZƒ��7b�+o
�>�n��bvۤZS��2dy����on�K���4Yp��p�/\��}��>뭬b������=�����V"6��ӫ$!{v�V�!Pۦ�;f�6أ���5�]�ۛ=@T�qtN��*u��2���p��4K!����u��ɇCŚ'����W7���Gf��s/C�Ua������?u���綋���uR;�8z�q��+�ڋl�#�����u�)&50&O�8�￮�{�Y�s��
�'���d���f���GM]� �������7h�5x*��̍��LxdrM��M ��f�~�K�~�����<�^��<JF(�]�UX��ȎL�7m��B��t���hK,m��R~jmI4;����ǵ�<ި@�v��1�P�L�헎L����7+(�=v���i��D���C��eݑ���7X���� ;�� ������;!��BӣX#a$.n;$��j�Ъ���!�ݴ��O����te��G!8l�y�d�O;ܱgª��K�_����@=��U�����d�
+���|,��7��<�f$�=�h~�,�&LQ�&��4W�Z����7h�5O�c�LU]�Hx�zyvNl ��]�Ls��n�㋪�F��g�-�߿{�jq�ig��k4��<��;���ƣ��G;!��i��8[-Hʉ9n$�}�/E
���ٛb�=]�vI�{0�Ъ�g���m�nR��RK$�w�,��������UHQLɦ�'�n�$��{	H<����œ5p��� ;�l@�v��cY�x�W�"�8H�q�wJhO�v���O���Fn�i5S~��<���n��c�ۮ���)r�L�X	��1��Eܥ�ܛ��i6���t�$���@w1�@z}��̶ FD�ܒ�jTFc��<�r��I��$��4�$���{@$~���
fe6\Uw�{H�[}���j�9�����#�t
����x�'��cRM�ѩ����F"P�P E�� ^�wXԓ�W�F�jLj4�mɚ^�z�g���x˯�@��h�E*cQH�v����5��#����&�7��tuȼڹ��u06'�;�-�ܥ&I|$���,��c�s��c�}Y�;� I�bNf�W�^���@�ޯ@��h.�xY�#2H�q�.��>�H����>��ߔ >��R�$�A$���RC��{��{���*���U/�f�$����Jm)FR��`� 6#������;�RϱҒ~�&b!V4!c������1��� �ɺ�����니�5�lhw+�&8ݣN�u5���j���sr�:t�T�iz��Aΰ�^M�n���'�F��8���=�W�b��Ϟ��3��ﱶ�뵷.4r�q�m����۲!��� 9瓬ي|p�0Z��"�8�ͷr����=�k�!w5p�v�fTtY{'9Z���ф����rj�gW�r��J����gwy�{���vwb]Wx]��L���`���qv�$�7.:����{W;Y���)��]]�m������;9��}���s���3T 7v�n�u `��vI��q��l�f��'���s@�ޯ@�D�M��b���ՎP�Bϱ���� ��qpn~Q�$�=�x��^�z����ϯ�@�������sIW>�H�c��c�}�P��Q.��2<K&��hXΞ���ӜN����GEnv�ҭ�n�E�zN��n��rDۏ@�wW�U�W�w�ug�>]~z��1`��Ƥz^�z���r9ȣ^�H��Ǵ���t�d2����LSR=��Q�U�W��	unk�N��vI�|A�`JF[e�Wr �v�v�:��s �x�� >�1k�����������v:@g��|� 7��G'M�SSB?�A�ܻ��A���E��Նp��[4g�van������?g�]��ĳe����Ҁ�cR ������z�����EZwD@9ws�*�^�k�o��?f$�\m!���N��8��z��Ƥ�^�Ԙ@#�E
����;�g�RM���RN_�cP��BH�q�����V���-�'� *����d��1 L�F<F4��-v����*���z� �޲$�pf6���q��$���:�t�d��@l�X�U�GLY��s��S&&��h�]F�U������V��\&$��C#���-��L�:����(�5"�"Q��~b�2'���#�9}~z�ՠw�uVנ{�D�+bpX�q��vO�-ٺ���Ŷ,��3���"�@b�Y��y �{>Z���i�9�F�H�ܮ�U��}v���h�)�Ci�ݬ�=�����]�g���vc762�*Wm=��cgr=�@I�����^:@{�ܠ�s�Gd5��.+ƾ�rDۏ@��j�-}V�{���*�^��DU�$Q�І��-}V�{����ľ__�����h�vp'piL��MŠ^�w4
�W�{�h��@�ɉ7�(�������Z���/u�I:Lc��؆P
� ʟ p��iU8DZ$�À�H��`E����T"d*�`���xA�b���68~S�1	DHBAB1�ϸ��; �{#3�'p�'=bd�-�	�P�1�`IA�������4��8����$��,A%�@a ��I�;Q�A��0T!VP��w�M V&�[������0� 
����CH�$L'�v�SB|HL��Y���w���c��3�����8H 	@       /Z  6�       �6ݍ���vglG��UnҮ�rlJ��s˶��[����}�������,��h������e�*��D���-�I�V�U��g:3��mqC)n�e�4ͫ'[���( �2� �Z����٘#}?|��֨kVƶ�ۇb�$����ڦ�U�g�.��8t���gk*�i6*��$3�0]l�u¦r�#Ɉ����mkH:���^�l��܋�0]�rA�EiS�BUs�6�f:݉��^�î�{G]7gK������ar8y�=�]�D.�Yy.�^VGf��&��&;+��n��}a�[u�#������3�`��8���ӧ�8V49Sk`�d�8l��Stb���{�-[h�nU%֝nV��Mi��]+�*ܗ1�H�<��Rڱ����g��n�x0bT�f��)*�m8G��$�hٶu���F���Zrέ��v�G�n�﫷kc�#�;!&��5�k�;i�*P�qH#�]ۅ:"����l�����a��/�M`��.Z������@��
v�L��T��6gl��Е�9K�cu�p��mۖꍊ�]�垹l�*��m�譊����9��e:�'�\�[UXp��Le� {k"��sZڇh3�	q4Y"�:��{ts\7i�vۉ�Gx�wj݂��z��۫��gA��VQ�i��)�8ʫ�2�q.�Oi��벛 �gH6�n��¢�N��vVwm�Mmݭ:�C���M��5,�l�e�
Ԩ2�T��օU�U��R��k����]�V��X*tZ�z��gA�&ơ(RKT��anc&��!�[<\mtț���N6��u�9��t(Y�S#'����C��[���ό\]X;pfxYץs ��ree��������>%@���u�c.)�k�UZ��ԯ'=7+m=l�gT��n��1��{�������=7�Cb =A� ElL��hA� (�����
���Up�Zl�7$�I!2� �#"�;%����Fz�-�n���J�p�7�kұ��gEE�g=��7���}�w��vN�a�\Fr݁\��m4�N�ڻӴ��v��V�M�3�6���MAVX�/�)k��������7Z���K�і��m�k���n��ƫ�o��M��][=����۷��;�.*^qZ�H\������v�<�#����{�ǭ���$U�����5�N,ߏ�����ޚ8���pj�답��<�l�3t3�<xA�����h��@���h^�@��	�b�Ǆrh��@�׹�Uz� ��7�H��>q�8'1�cREd���b�8����P�T���}4�w�S�$��I9��s4
�W��4_U�^���9tu���pBđ6�I�̖Iڭ�~^��幠Uz� ��i\$&"&3���y�E�V�ڹ �rl:�8n�CSv'��?<yIc�4194_U�^���*�^�[l�p��N�8b��sn1��'y���'� h���X9��@1���+fO`m�ɉ7�i�3@�}~zoY�Z����s@��i��27I�9 o��r�xܨA���{H�"y�bNn<�ɠZ����s@��zoY�x���C���M۶���$�z�`4�� �˪_f# ]�ie���q���#5$Z]jzW��z���h���v��p5��'w�UP�'w6Y'u���=��͊��8�,�&�z��K$�<�g�A�(�(� ҙ�b!�Eޭ���ԓ��{�g����"��SE��tKvn�$�_�O@���޳@=ó���PjIȬ�����'j�{��I;��@�ڴ��LOv
�M�9�\�r�ٹ�b�v�L�١��.��'T��dě�G��8��U���f�k�hu+�-����2'G�9) 6ݭ�&M�ݔ��i �H��U�n<�ɠZ�Z]J�
��@-�h�WI��"<j8�������d�[��y��Ɋ���J�x�8��}u$�g@_C�71�5&�U��+���V�{ܬ�=�+m-ȢD��+�r�mp��-c�x��"^�ی��o^:������0k$j$����^�k�h����k�<�`d�F<D4�Nc�W��	�Ų�:�u�'��z���w1����@=�h-�F��s�>�{H�ݔ|\&)�Lo��٠��Wj��Y�[V��dN<���@/[4�ՠj�@:�4
�P РHڡF7�I$�6� 2��,ף�'D��:n��'nmci�e{I�^6
��Vc�Y����w�Α��Wm�����a۞9����܅:��5���i7����<kq:���,
C�F���,��;j�BFz:�����zw� 7Dҵa��k.�7M���0��3�u,u�:��[Q	Ƕ6�l������+�u�vC!�ݱ��j�D�����v��$!L�T��ý���&n4@�e��y�Gt����7�ѹ!7쳷8�T�%umd䗲h�!��ǉ9?��9�����Y�m�z٠u��6���B��5� ������=ݴ�v��['S�`��<$��Ԛ~����Wj��Y�r�9�\���#Mɠ��Wj��Y��~���|�{>X$Q��Ӓh�c��˴g� �@w� Ʉy�s�n\v�yx���H�'����ĺ�M�&�n21�=�k�[�9+�����h�7H�v��V9@{-��q������<]�v�B� )�����=����VhՅil��#ǀ)�^�h���/�/���|�8�&��px�q�NM�}V�u-���zm�@��������d�8��l�<]k�m�����1��9��6��D�npv�p��=m��\0�-���D`���n]G��nc����zm�@����W'4��$�����Z5
I�@-�h���u-�]k�<�|U��E�M9&��>�@:��u4!�A��@(��6�P��?v��cRI���u$�'ڝ�LjA('"���@�u�@-�h��x:Q&�'QLOI4Z��f��>�@:�f�UG~~W���`@��5�B�\�<�雓�������7Fq�ۀ��x���<�G������ �U���z�>M�`(Ф�<Iɠ{Ϫ��Y�x�נ���Į6���B������Y�x�נ��������\�nd�jM�f%�n�$���d����ɤ��"� Ф¦*��rw1d�OF6VБ�P�8�z٠{Ϫ��Y�u�@� Uwt)4��"%�Sh�H�{-OS�r�V�%�bx���8�wd�"&�uE�8Xǂhi�<��- �U��[4��@<ò�;��ԂPNE�j�@<�f�^�h��x:Q&�G�LOI4�l�m�s��l�-(+�dƜy<0�M o�3+�f;@m��+&�Y���$��RM��Z��4�ݠ��ќ���������u6��m� KrmknGb3�\#�[�7�R7l���rq.�!
��kִ�f�ݧ/^��I�Ñ.,>N�/&�7[u�{�v#���[՟j���A�e�m&��l�v�C�K��+L";T:�	�8�6{=��A"i�X�x7E1����s������lF�\ ɮK��urx�����W����u����>���Y���3�L��ə�UT������E"JLbf6 �&4n�%ӆ�]�f5X٠G�y+����z�S(=���빺���}?��;�� y����(�r�d�nd�jM �{��=��h^Voٙ�"��ؾ����#�I�[��=��h^Vh�l�=�ů�E�M7&���2q��@G��;���9ɝ׶�=ϾJH���r- �u���ߗ�燎}~����r�-�� ���!�Rfn)�N��Mr��;I7.6���ۏj�i� ��H8�jbx"I�������6�=��̇�WqsW�80BgΤ���s��
�Q  AX@�C�;�⮹@�v���o""d��6�,NH�%$�-w�N�@<�� ���;���m�7�F�8����[v��h��(dd4�q�An�.K$�fd�NХ��8I���@:�f���q&�0��$	�i]�qt�uͻ�.l��$��v[���H��Y�0k$j$�I&�[�hϪ��Y�u�@�\Z��Q���rh����h�l�z���A�>�G#FH%�Z~/�BM�Χڌ# ��j=ޓ`iM��ɿ��ȃ� �a�v�w\X�C���i�Z)l�I(�bg;���i4H�˰,�8?����L'�Y�E�C"�»�$Qހ��0�่�DCbA`��B(E�$�g��g�|�|B�_ P6��|!���!&R.�1h���V�2�L�2��'�`?Y$�>2.ɖg$Yc�:��v9G�w�̺�|�Dp?#�Ҥ B!� h�$�S����q�!�&EQ ��*��`�eEt �K��TDjH��! H�q^�� ֕.��J�t ]���߲Y':��y�z&ؒFb&2K'�_f�I�͖I������PK4��$��H�7!��#x~�@-�4y�Z��4ζh8���6��ma���q�'4�9�.�%�k�wS��9#��ٸ\��^z{=�I"pmɠ{Ϫ��Y�u�����'w6Y'st�q$�l#5VI1�� w� �v��V9[�G"d�h
G�i�lc�@=�}4�f��>�@:��������,�U�ݠ۴��� �7h"";��p�ZBA�(8LIU01�Ď$U%�FE(�(��*)KEV���. � ��<�G�ν�I6_N{��Shi�4y�Z�+����o�M �٠fb����ģ�gga�{/O<�%ڈΑ�5���D7W��Ә'�j`��ő�D��x~>�h�l�m�~���4�����bPD�fId���K� �>��,�sw����@��U5�8���$�[���hݠ�v��2��b�2I"j$��u�Զh�l�u-��d�����R%��d�#rYݠ�v�n���&���`�+>y�_S1�g9�r�k [�IWR��ix5�]h�zYf�R�Ƹ��k���gs��[[����q�&��v�ջ�u�G5c�s�r�K�p�q���n�V�q7q1�y�;�>�QF��f����+h�x��0�5�k�n-��+�iس6��+�]�?c�L�&�U�泊������]x�)4���'MӤ��Hv�v]`��̕X�A.��c3���T⨇��57>���2̮��<�[l<�=s��^K��nlC�W+ջgigh��,�#��4�61����f�[l�{����@��rx�c���#�I��7�ă��h���m�b�ט���bM9&�u��1�G���v���@�Nв28�m9&�u-��٠�,�
	f��$���lF�J�,˴��@�hv�1��������f�x0�5;Z�,��3�6��gN�Z6�+�葘ݤkm]D\ɷOU��@7wm cn�1�@۴���W�G$mD��@:�7��ݙ�r*�*bM�}�u$����H�4:��	&��$nM �7hv�n�6�܌����/�Ә��&�u�h�� �l���@��rx�d�Ad����۴�"9�{����f;@~G{�������8��<�j8�3�'\[me{u���2�9u)',.��ܰ�Փu�M9'�z��= �[4�m�m�@;�'bFIoq�R؀=�� �HO���r"&Lf�¨��ĦD�d�@;��h[^�ً�oX�"⤊a�j���U:ss]�O>9��=�Bƛ��p�͹4+�h�mz�f�{�@�ӈ�y^$�50N-���������=7��}h�nP{�V�C��$����14��v��x]ժ�ÑZ�^�k���+h;u�3�x�@\��� �� {������ֽ�v]�Q~NA�94������n���kc�#��5�FH�I1����y�� ���@�wW�v.-y�H�&$уqhq�@��=9���r!��s����`Ch��z� \��=Zp���28�i9&�{�[@}r��^>����n�{x�{vM���S�uZ�Ԗ.��쎊[0�u�6���t�)�t=�]����tܠ�w��v@�=��}�67������<�ՠsv�=�;@zs-���"��itG��H����OwޖI?t�%�@%�o�@����@�ޣ�D�M�#Hܴ�1�Ә��M��DϞ�>�s��Q~�cLrh������ݞ�y�� ����K�����K� -����SL�#��箻�1u���@�>�R��,t��vMG�WlsnR@����td���u�l�;�y㺲���6�=�����]��
z�ʗm�ڔ�fy�w��kYTm㶸�4k$1qWvhw�1��IiiiR.�Vݗt�:'I6J擩-�[8$�7+@XH��C�#������v�axyҗ�6	Հ{Z��$&s&s�� /��@|�D��w~����0j�8��cZ�e������>z�i4-x�yNe������i�PY$Ƥt��- ��g��V����|�!H�&$уqh�l�x�4Wuz�ڴ��	�1�)�I�4�:���^��v� ����pL��JC�MӘ��v��n�a����R޹������<�)�u�@;��@�wW�{�k`��K����#��}_���ל���qg8�[��#X���&���9�4���呂wf�{�f��YM�z�YBLd`g9�3�I'99��q�E0p
!�%�#�}�F墱��Qr�@��Zax֤�7��IϹ��Hu�@�;.�N(�N1�94��4:�h�l���9{��*#n�RMβ��[4��4��4�ů��bbM���w��c���h� �E7���"v�S��k)�S'7�͞S���=�)r$j����ɲ��B����0�hَ��l@���q&�k���D�@=�@�빠u�@/��@��7�dn8G���s�'9��Ԓo��u2 ~D� � ��+G���HI5��gP:�4=:&��xd�A��h��xn�{��s������z=dBĘ��)�@=��h{�h�Қ��4}�5�D����f"}-��s�#n9T�{x�s���&��$I�IN��	2C��4�&�w�f��)�^�@=��h/s�ECmA�H������׎��7h�c�.-x�h���/Y��[4�1*����>4����BEIG%��(
	w�vY's]�~���Rk�"��ǰ��J�DT�+j�޾K�I��tME7A)��K�@d� =� �� {�w�U�e�b���< I�F���9��OT��r�F���M��cqe�p���f��YuIUt����@m� ���c�AU�=�,Mϙ�IR��v��!�n��{H{���#��3/��D�M��)�@;���.�H{��ݠ3!�I3vp	�����@d�:@{�� �� {�v��{��.&�mD�&	Ǡ{�]�~������w��̓���Ƥ��E_�QU�U�DQU�"���U�����""���PP?� � *`*b*���
�H
�R"���@�F�����ET *D`*��@�`*R� b*�
�
�A"� *R�Q��EE��DR�
� *P��E��"�
�R"� *H
�
�H��B��"��
�X",��B� *A��@A"��T
��D�"����A"� ** ���B�"* �H
�X�,
��"* ����A�"�H
�P`��b*P�T
�P�"�P *`��A�"�� ��@��Ab��F�  *V(� H",T *���E_�QU������*�U~DE_�(���EW�(�*��DQU�
"���U~U�b��L�����n� � ���fO� ��>       @   �   P     P (   *RB��Q@J�
)U �Q@(I $T	
A@ (
P�U$��$ HR��R�        
�E2�O|�f�rk�[�ҬfU���
��kq>��osk��Zr�K �s֝��io�| ��:��q+� w��;���δ�ez���]� ��O�žZ��k׫͕u��� �  �P@ZP=�/�y�˺\�盼X<���{iq����j��n��ƅ�͸-R�Z� w{t�f�����5�����y{��^o)�3��x }���o��y�h.Mv�o}n����    ���� ﾵo:[�s���۾��w��V�}>����}���׫�q�ݼ{�l���ﾚw���/m}� 7x��{��s�� wR��w־��Ժ������:W�� /y�g{=W�6��wo-J�r�V�� ��       a 
=��ӓ��O&��-�
\f�)� �:S ��h�J)�4�`t���)K,  Pb4S@�E�:S� ��JRݹJ ���e��h� : �JQ��R���S@( �  @
((b :R�f�JQ��1@�,�>�J]���ҭ�����ŗ{��r�_x �=��e�粽�wx �{����o�C� m�NO{�g���ݼ����9��� }|)��o+�wO���r�����m� OHS2R�  E?�5R�� �<z�U4�M@  D�*��j*D� �T�Д�R�)   "$!�Jh�4)�'��~���_��a�?�'�������EU~j��UҠ�*��U������*�PUO����_���Hi��s?����I.�^��!H`�����t�Fbg�y���Ӈ6l�4:����q"$ dpH�%!�81�jH�Ie�&�!;�R0Ӷ,Baq��nFP��!\u���7��4��-�5&��h��W�Bda���/�v��$\.ݧ�5p�ӑ����@
��*m�~��XW2Efa�I9y��L�i���B�22:�L4h����[��n��<c9����8K��=1�E`���V�)/���J"I��J4U�$p�0�YXL53N�4l����,F@ BA[! �$ ��fx�H{<�6ĉ)"�H$`ĐY7�u�F�d�N�_�X�7)�'�����f�F�Fhۼ��)Nxy�k�P<�����HB�0��! Hţ ���>�8���-�����w����G��M�$���)�sIĔ�)�#��n��	�-t��JxO�<�y�I�@.hÚ>���a��kiC@pZdֳ��b�R@���!14�ĉU���5[Iaɚ�'=�jl�CHm��HXŁ$�.�g���8���:SrȘI	 ��X����f�����g�1�i� �S`�{�����n���}���G/�Lf��b�H��c�&D+���zF�:�sXMy�Z����M,xf�K��F����%�Fs^\=���s��/<4��b@�Y	����<.�n���Ɏi0c�����\X@�m~U�R�H�+���H@���܎�����`@��#	!
R�����#EI, �4�L�50a	@ę�I#RY'�ܒ���]�!�mc\p!I2e��)Ť�(F��I ���:B61�6�'�h�x�10�a�ha.�I`�h��[adL�nI2R{��]�(�IuO|�͇��`Bᨑ"B�l�B�w8>A��`c��!\V\߼扜��gOo�9�S����.�h�|�#-qӲ	��rf��3�Yw8I&��I��n�c�\�=��sU!�����2�K��JJk[�߸zs9�� Q�H�p.,B��#�2�1!��m��ZI��2.$�I�f�%+X��
���X�Xa%���3��-	l�]���p�f�M�y�������bJk�$OdH�d5���4Թdѧp�#���O�(�@�> =��8�1$	#Iu��G�"rZp�]x��%3[����ܨ����Q��K�����$!"i�X�3�=4{��k���ל5f�y�j���4���@�� �t$�R�����d٢h��bj�%�p0�5�q�2�S�����5&�H�M�o�	��9�����!$�4S��.�ۨ�|Y=41d���a	�#���HYkf��B�1�朕"F$C��aC5r�u#R���$a�K
i�*Gw���a�1�$=aYSa��bE�xO=����[����ak��$�\I7.h榶cy! H�"P�#$��ǐ��sl.�ka87z��a�VRR]s0����CZ�	y,����В6REܐ�L>���p����B����$���	�I
���-�	�.�|�p"BF�$�_��Y�%�>6�Xl�7�0�j3�5q���P��.�! �~�� l��nm�@�G �Aˣ��	+6csG$����iw����`g�z�I�4s���a+π��� E�B0#@���Í<���$�y��g'��0�K<�u_[�I&��WI���2r\N&��8Ow��;��$B==�d�H���%��f�"ԑ �H%8p�w��ɭ�ǖe<HP0r6ID��`!BR��0$	��'���/�G�3!��.��H�B4�B�����IjRn�S�RE�e��8�����Ts�S�<0�Y0~bP%"Ϥ�Oa�ٖz}�r1
s �!�	�Pld�K�3nq<33N�2{#aO#���`Q��I#*c,*��R�HN{�~��}.�P�)�5��B,,��-RF0�G��ߧ/�����{������P�!HЍ�H�!H1�	#IC%2w� S�<"���`EL,:eь�5�8X=!�g�F�(K���.f��/����\����<��� \50d|rQq � X��a�F6&Fa�x���5��l)
ā,h�l��J`K�K�!L`�D)����{��#�$c$X#a��a:�bH�HĄ`HP�=���H@"q��=���rD��]��h�JF�,,�����z��'��@�P�Fbo4j��xb|�4��LԊnHYp��D���#\aR�	L�a3D���[��(h��ywc꾢�c�4�p�¸�
@��I�oC�dp\!L)�bSZfi���dRQd06��$�����3F���a��9km�d�A�jFols	5��.�,�ʸM��|%����x|���J�I�͛Sl�~Oa~�r_y|�o��Zٶ��ٳb_RY�6s@�;�4�&]�L��NsG�ۄ7J�F؁R- F���[n�~͍x�w3�!#`RYI-�).��`�S�_�Č<@!cK"S�3�M�q	 �Q=$Ob��P�$ �A"RHD�@"X�`E�C9��e1HЋaWЍr1�㣒,�I,	"`hv�(�oR���5��BB0$�H�dY��fka�����$#A���b5Ȳ D�.$I�U�Mp
@��=���2�BB2/|�I���H1,l
JBa$5�4a�E�C��=i��% �e�$+�e=�D=�@�!-i�k�����J�����N�|_U�t���B�'Pָ�8��ㇼ>7,4�� C�7�1�$�@�	����4�94�ZI	rS$&e=rh��kJG,�5���0�x[�|-��HāMky͘���tF��s#��2\4�$٢$���h�˿/�3>���H�)��h�d Cfds��$�0�d�hH��#(BG�>f���!LD���OB�a����!Bd3��Wd���B�!%��ݳ�������B�}����zJy�9�\���8���76�Ԝ24ċ'%��$e�|s&��2@�CBB�h�X�YM�e��x���$'��hf��8�p+!m��z�琧��\)v �3(L�kD��ޛ z�F�F��h�	2Cĉw5=���0��۽��$
��=9�0������-I`a�t�Ò��xr$,Il���z�8l��bK����~1��.�乭�(��3�+�� A��!ӟ��8c$F$}C�o�5���,��ՂC�C�w"��� H���x\�l��<4�iϷ��,���,��<a f��.�WRM͜qbRC\�(hH�A�a@ȕ26A#d4���D������Y!$�$��4�s�9��Nj�n��L�}�	
;�����]�Hc�Bx4a@�`ő
,)u�9'�q�@�I��.P2BMk��%i�6Y��L��A9�h���\ͤ7 �`�!SqY���B&����9�B �����~�O�x{�T�YB�]��/	I��6h��0����BG��y%\BJX��>+���Bțd�"B0���7�����h��!B)Wp�~8k��2�-���\$	�>J��R���=K�y���HCT��n�a0�	R\%Ĕ��1`Lu��e�!p���{<湫�%��Mr�R�/��.w�ð
��R�D��0���R �{!��)�He`�GC��C�� xk~@Ó�82M�۾�"F,��;d B-r67��i���D�|h�0"B��l(��lFH��
d`�.�Ray��#��,`ċP�xAdX�	�����<�͑)�窇�Ȇ�cQ�M�K���-�@��w
`h#HRSP�j"�1�O���P�n�2�@��F0,bc쑉-�i!dL�D�4Ĝ��kdf��	,�!M�f�X��IH$�~x�14n^0! E����%3[#C�/iw���� ��l   m��p                 �P                       m�        p  -��        �   -��m� H m����  � $     2��̽C���[@�6�jޫٶ�m[m�l [�� ���|  ^�� �fհ��K��
�'.)�T�Yz��Am��%�2ׂ���)ջU��P�^+��I]9D�m�%���U,�m�l0MV��   ��Q����$�pE�j�����Kʹ�Z���Xs�Tj�ష6��bc1��c��Ëv�`m� M�AM�*��N�nBy�-��N6��QNni��`��#�ׂD�n�,�����$�9�%��6͛e�@x�tΓk�ݯZxt�ȶ�	V���-�m�t���lm� l  ���U}T��R�;�Ȓ�Z����k�-�޻�}��>Cimnδ[Sk�ʕP��mǠ:�jU���T%F��eXXSU<ά�(�q��f���S"�ыVղԪ�d���uF#�UQ�C��+��OYm����BN�i68m�]�(=,�Cq\TvR��7:�R������6�T�JL쌃&F���[Ie�UԤ�
���p�UT��f�fU�X+g�� R��h �ny@U@��U]WmL�H� ���ۭL��Z[e�h�� �`k�-��m   �[%����� H�`�)������:Z�M+!�ں�w%���� ;(Y3@+��v[T5c���9l[YĀ�L����6�N���lx9	:y�ƚ�9��Xd\lG���Ԯ�UA��pmRNrN[��q>�+}�SlƜ��N�8�N��h�Kq4�n����m R��}����l[G
��6H �Mqm�z��f��]t�������i�;k��������r�r���*T6s�Ul�s�\N����U��������� +8]��3��j�jX�(S�T���^�-�UJ�l�Ls�n�.�[]PI��Io^]$�{m�`/-T�,#-H"n�m�ma�`���k�
5�U[@[T�M 5Q�cWP뛸��v���1�=S�
wk�nZ��V��gT�l��n���c�kj�ݮ(Pyg��*�ڪ�Ā6YҀ��K[m6͍mջ6Z�bR�6`�y��I@]��]�U�Kv�v�3mm�  �c���!J�UUHQP+Hu[[@r�/�٨���v�,4�o^h���m��(!N��SuT�n���-���H��8&�mi�]�l�@k�$i��f�x���9�5,����I`%K2��Ks��U�m$Ѹ��`�l��C�a5��I�kM� IoP��kźI�gk(��F�Bn��k/�Z ���kz�mԶ (�ZY��V����jc�y�W�@W�^Gs%�[m���r8���
tU!Ll2�UC�(��2�:A���퍻u�$炮���l�z�h˖�u-)WUR��e6'��̨}T[ ��;����f�3J5a�Bv�۵�Ս���<V��� ��܋+[UZ���v�$V�!��ܵ�U`��:�&�ʻJ�յ]U��n�����p��a�v�I��u�Ig]����p6�2m� ��9�­���#�$�)mU�(*[��j��7d� -�k{��􆾩.Q��    �!'�4�E��mm� ��^�֮�� m����������z��H5�Ke�����V� L�R�o�>��q�ٗfɕ��v���6)V�N�m��m�a�.��M. �k[Cvݒ�j����Ia��.�Lq%l@UWl����z�m��[@ � �a�h�p��;=�Qn��[��`   �cm�m��sm&D��   �_�|	u�6�$ 6۶�&�� kn���� m[[%�Pl��,���*�UR����N�6��ݭnI��
Y6٪�8p��m� �v�e�,	��태�kdj�   �Z�lͶċ�6Ͱ  ��8-�ݖ�@@W]@cJ�!�WUU<׭ݻ[Am��,]�R1�[��-��.����a�����m��h p���-� m���Z,��(-qB�M*�"�����	)��Qm�-n�$�=%�m��^�\�Z���o��k���l�  	���>��nUM�m����` �A��MSY��uO���+�+�u��C�[�j�r�������76���Ы!Qv]�m���e�@�n�[NL��V��������t�qֱ�7Qu��꣓��k)u�;V�����ۦ'���6�l�gy�+T�6H�)��lI=��î���^�����j�A�6zN@۪@YYn�7f�SUR�pv��'MQ5MM�[Ֆ�v���f�uM��C���#ulհԂL[�����d��T,ԫUTUcl/l�I��вZ,�kv�;N�"�jU�VH�63��� �$m&�B��̒�� �$��չ��l ����� ݶd$��m���t6 m��&m�<b۶�  86΋uUm�e[j��vUe�`�;�dx'�Z�}���Y�Ƶ��/@ڑ m�k�P �8Y,�%%� :��m�כ �a�a�����8u�l�e,�`|���^ ���m��*�m�l��i!d�/+K�+Ĵ��v���v���m� �մ���J�T�H���i�&�ڕ��#@F2�*�TpJ����0a]���Pҷ6�f�+���ID���m�j����	$���cg1�s��;Q�0�S�qS�l��5�۵��W5��7(R����E��d)6����x�Ͼ����� r�$��S��e]���8K-�z6*�j�m��VU�j8�pzɣ]:"SW�tj�R�t�R�]�j�g����uP�Ne*k� �ء���R��km�6l <��nޤL*��:)�x8
��V^���]�����-N����|-�l���m���Ұ6tH��J�����උh  �`  Hh %�h���Q����4��~U��8��ku�[`��-���dU�e_���YV������  ��u��c� ��6�l4SIk䓡������}�����$��Ik   [#Km��m��-����Z�� 6ٶ�o���?A��0[UL����*�U.�7l �f��n�h�.Ā H-� �V�U���ݹ�iM�@���,,T^���m�kn��-�[X�f�ۤ�m� ���`
Sm�e��j�3�R�AH�(���v��n�&�'�μ�P�[�6m�wM�[K�(5R����UTHv�kl�G4��ŉ��)j���@UT켮��-�3 �f^�b5'����	SST����m�-ָ�[z��  ��v��i�l!v�S��������ICÝ
�]J�+N���+�:M��7m�jn�\K)  �m��sk�a��Ƴ 4�e�Ӻz����J��N��\�	�ڻu֌Ù�j��H*�Woj�[[m�   ��o����,�`�9���M&�`  U��*��!��^�����6�� 6�� rA�����m��m��mp�4���m@:ޭ� ��	"Y���-��\� -�m��` [Fհm�m��   �m���ͩPjmU/,�ָ���*��P ڶ l �m�9�M@�N�Ä����l	6�m�J�VC ���m��e�66)U`�L��=<U*�W;2�KiV�}�B�8�m��t�����5rJ�M��[�u�n�m�g[wQM��vطeRж�n�8�`����5�i6 ��}��m[�^���k	 ����JͰ%����R������m�Y. ��s� ��eڛV�� 6���t�[:S�V���8���    ����[׀l��$m�-�ŷj���6���c �l�`��l[D�b�$����m��tͰ�`m.�� 	 ��մꭰ�@���J0�h [@ h�u�X<�p����km��� �6�I�m��ې�����R�U]��vvV�4$-행�j��cm��T�*�hL���A�����9I�) R��[uR8��ҵ@K�;=�Id��� sh�OYãF���:6��ܠ�&� "C^A����Y�[�� =T��\���� J�Y�&�t�I p�I4���[[?A�k4mU�=�(m��[�H7m���l�ML���@X�[h;�[z%�M�g"Z77�ҝs� �.iv#\�3/��^��ձ�yMzd`U(I��nm�
���[nԅR#�*u�t�� �[F��@���yk�j���B��А $F��Y-�k[m$��M�����F[���P� �J�UKk��.�]�7�V��� sX�e��f�PUM�?�8�j�?� l?�� 4!��W� �)h`b�������V0"!�
 U�p��آO]�)��Q��S��8�8|�y�J�h�H����Fx���=�F#��B ���`D�D��@؏ʧ���!��U��=P=TO���#�UN*!�6�?x�����B|ht�P���S����Av����m�0�C���D@6Q���x��qE�Dv��P"D��� ��E=Xb Ea(���ǂ *'��#�~�!�l�-a�� @�����z49�B�Fz?U 4*>���@(�.*� �
�b� &�D_����
�i� 6��
���� �� �#1*�bF 	*B HD �z��*���W�4� �A�P�a�|'�M	����h<@G O B
 g���l	*���>$"���j��(����A������CՀ
A �����=D�)�	�t�Q6�}`��U�G����Ȫ!"1c���(Ah%��G��0 @B��������       �a  $t�m�k�im��,���t�C#����ps%6�U2���vŖ����
,`�e�3�ge������53�ywC\ݵ�Z�Nu\���.�l�[]=:0ZaQ���(vE�ny�֡zd�t���-V�l���ا K]J���:wQd{���{2Z��o
W�Ӳ�(��TÀܼ�]&�Y�WN$n���v���c��q8N�in��D7]�v�<�$ׁ.�pw�/d�,=���U�̶;VgY��jD��;N$ .LVW���
N�V�b����`HƻsӴ�s�m%�|� ޶&P�W�=v�vd5��v����p�݀�9�4����U�y�Z���%U.2m�O�c.7<jg�n���e�g��m�J�mmKQ��`A����v���V��#8�����9�;)	�gM�(M��v�a�`ѣ,�8h�۠c�Q\d�r�p!0�G'!Q��el�:b��2����X�p6�tn��̶:�>ТWE���鳞8�ڸˆ8���XJ��O5l�j�W5]�d���ki�l��"m.�pr-v�6�l��x�	�5�t�J��*�#�����=]mK�	x�c)�q]�<8Wi�a�koV�u���3đD.�KP](۰H����t�m8��l�,�����Nf�ud�H;�a�1Xwh� �,��cQ�Wfލ��8M�<k";;[4+F�ƃv��e36q-�^%�R�SV�H���t�"IƋ%�d��XǶ��F�I��ӭ��V�e���m�i�M��0�����/);mHMs��x\b@ݻa)�d�8����jZ�Gcr��mUU�*���`&�N�v��6�7��
pGmm�F�7]�w+��S��k����ջA���#�gb�GL�cI�j�ȝ�Н�i+p��F:MS�{-j1��եc\)�j�%�+Tw���;��}�xSA�?��৊�x� z��@������֪��ɻ�]fm\��`n�K�ʖ]����i�K��^�֐�R����g΍�����i�E�$��lO��A;i˹��
v�K�Ŋ�t�"�\/p&&�n5ӭp���iK=�m8;35;��I����ҲXB�F��S����}mm۱�����d��m��}+��#�5^���2uS�� R�wlaf����5�ɬ�(�QѨ�m�
S
\�̂������r�nݕW��*g�\�L���:ߟ��H�f��گ񯾯�`����:��xX�����h�߱"�w4uڴӷs@�Z��dfHI�p���#��y%�T��ڱv�8�$�	'3@�]�@�T���2*@���n����fe�����H��@H�^H��kq H�rI���m�e���;�v�=��=s\v���,���&��FL�7wkLݤ\� qR�$��n��0��lkj%4�ݛ�o�	!j�$!(��W��%��-���;e4
�UlY ���H�&h]�����{�%���@���4+��Н��3cr-���@u͂� ;nL@rVJ�Uі���AI�;e4�U��8�k�-;w4~��}��BI�12cb� �ݝ����@|�n���w\F��û5�k�ZY]d�D�I�(F�>��s@��@����9�)�)�Y$lG1`�6��& $T���*^��3��$i������z�_nh�V%�P�q""k�q}Ϲj���d���v�S�I��f���M� ;nL@H8��(�R̟fx�Q(�v�M���@��s@�����J!�:C�l�UK���jˁ�e��eَ��d׋�[��;�x�jn�'�Q��Llo$qÀy{��@�Kw4���9�)�u\��4;�~Q4ۏ@�$T�UU��{| ��@;nb ��ehCX�!�d��4���9�)�K���@�Kw4�ծLSS�/7D\� �1 �"��T�꿳39�����@���PI�9�� $T��\� =S?D�n$�M��f���\i(3�˱�Ξy�{K�]�������g$�m	H�������;e=�� ��= �u�(��I��f�����@;nb�EH�Et��>�2�//os4@u͂�s�*@}l��Wꭉ�ci5#���Y�}�g��	EHɰ@u͂�ο�;�~Q4܏@�Kw4fw��������d���D5�B�,��@ Q ���{�{w��� �jG�7n2HM0�%���0���;�ԉ@�;)�*q�ԁ������ؗ�tm5��+�5�p�n����Y5-֗��N#R��`�l��{4��.�!�g:���_(ļ�x��Ep��Β���{s�c@c��d�օ�Ĝ87Z�� ��9n`Ғ�!إ{$��4F�-�j�b���G�竎۷QٝE�`y1����5Ӻ�[<����!� ���Tjfbpr\�X���n�u8y���%��7s�%��qt���FMu�^�p��s`�v��W�r�����cuɊ3$��q�h��BI6c�ٰ3�V3+�䍨$�Ɯ����^�ޝ��-��>�S@3�R�cQ��$��:� ;2K@vM�����91Q�[��1�a$�&h��h���:��6:fZ�6��h��C��͜�yyy��D��g.dݣV��\���1Ӹ[gl�]Xɻu�/&ND���m����X|̛�3-jI/�wg5��^�9��I�rUMM_3&�B@��PN��H���H H!�	��Djk���ڰ>��v;ܵr�_�#���<v'&a&	����s@��-�����J�Pʺ2���Pꕆ��B|��vs6Ձ����>�[��}ln�1Fd�`?�G���UUU<��:�EHLr�������,�����kٹ����3�n��T��Sk���������ƙ�[kU�A�@;똀� 91�@u�� WmJ�q�G6Г�@��n��?f$w��h�ۚW-zGQۂ�̄%)tJ��`s'��w�j�"!D#�.��r!?���6qwmX1�9y�k//oov�n*@;였� ;1ՠU��؜@LM1I$��urנqӊ���8�T�q��ywyZP�L�F�W[vq�^{���.H����vl�C'U��OO��q=��~��"�i����qR��느�� *�C,	sCr�J�Xd��Bl�͵`g]��/.]��G=���6dr`?�G-�<� ��ZvTT���- ��λ�d��"�ә��.�v���ܰ>��;����!B]X��j�X�T��b��48�˗s@�g}/��z�nh\���ex)�y1ď�K̾@n��\���t���z�n��\7Z�f�`�r	1���3@�}�@�qR�d�쨩�(�����f]cj8�Z�n��3&6U�y��˹�r�ՠu~�'LRI&h\����f9h�T�w*g�YStr~"�����.���V�{۹��.�Z��W(�<����2L�91�@F��Ɉ	�QR�U�VI�Oڪ��q*�!@�����,���:{��u�"7m��۞�C��8�:�M��f�ܘ�>�km�ym���	�F��y@��*�cn�m���+��UP9��anN�����W��C��a�1!�aT�t�f�G�p,�)��9.�Y��[k��.t��Ѷ5!�r�]���$���ݺ��p��7W;ë�f�{`{-4v��ۋ�dĹ:q[��{��wv���[N癅���Ë8i!5��Ǻ������9$�ok�&y�m��L����k�y���ʐܘ�� ;2K@I�g]Ʋ0�b�ci��:�k�>�[��r�V����kH3�R)#Xԑ!��56:�-X��vyDBM�3mX��zGQۄjF�cPx���ڐn*@;rb��T��WIys�CX�Q���9�����y�/�nh�ՠ��CO&�N0X�`n@��u��㺎��ۮ��8I:g�X�]6�H�\@6��I�z�Zݥ��9]�aDDG�33mX�dħ+jf�
t���@q�*EW�y�٣Y%�#�R��h��Q �i,qf���H�T��o$�\"�dܛ�[yf���ef��qRۓp���ՠUԳ��Y1��Nf���c�6!s4ߗ�wgu��rՁ�"#�������n��4c07s��{�ֱК�7"SuY�iVBK2]s!����̰36�g�*@vd��m�H�U�UU�a"�������ڷaB��33mX����Z�ID$����=���M����-���;��w<t xG�Õ�A5ѡ^�	��XQDO��p��s�2W��v Si���b���
�x�@x6�c���*|$ �hF�X��)>͡čw�D`I!�1 Ӷ��+�<L%۪��M�|�"���`'�B���QS��XB0	�] �jˁ$eX�B�H���"���h��˸�e�H��W�6��� �`&�))��0��B �P�wp �9��$2������ӿ����*t�OX0X��3a��1B���"�_F��Cb? ��@���z��ӜP�_����C� 1X���,��|Ý��6k�{�9����UST���vً-o�9���=�w�+���%�Lʠ�K�5V���m^�sgu��7��j�̜װ���P�p����y��]0H>�ɀq�jn�)on�9KK�D1��mtސmî�3��ܕΕR��!���y�(Iff��nϒ_?$�&��=j��I�s�
R�&����vfm�؄ٙ;�ϡBo��ڰ;���>�R�l�l�T�SN���4�8��{���9�o��;�����3mXs�H�Q�q�������=��H���33mXLvI��	.Dq.º��=����"r,��H����H|�U���� ���V�����V�-p��Lݪ����q}GW]����7l1���u۶Kk��@��[N���T�c������X,�͟��i�������q�ނqa���2G&���ק������~���o��W���4zF�Sn=���o�9��-8�3���[纓a��Z�U$���T���[���ڳbx�6lf�kT%�n��o"@�<rH�>��v��[���6Ձ͝�`db�(P��ȄDX�H� ��H)�"����q��z�2�UA��8���l�g�e�3@,����]����c%���cv�Xz �S<�8��m�Y�7[S��&spV�;1��^J�m�M���.��m�o	�n��v��.���ϭ�Ѣ�Vڻiv?����O0������]#-�v�59M�:1v�nL>�n6��nyI]Ė;[�LmY��uv��r��@p�O��(٭�h��͹��mҦ����}�ws��g����^.[�aՂ�A�s�Ëv�v/''V9��.���3t��vu)UM:��\�������63M�`}��}� �e�����7�I�k�vvx�}���qR nM@K�㰒D�0�49�����@��V���ڰ�$��o��� �j��S"��SNi��6ffڰ�����3M�`��Ͼ�yh_����D���$�L�ԞNń�.���_�;���{�����{����lu�ڤ�6�y��qg �\����2�\ ���U�N��z�.37q�R*@G�Z��^������a�}��.xcN	��9�L�/^c�N-B�d$Q��j�׹�`}ՙy�������~��M�@ŒI���*@Krb��T��$��e<��c�AH���hvנ}ܷs@�v�������(�5$Hhq�u"�x�dT���1�s}�An.�H�L�g��3�aͻn:׶�{��#Zp���n].'�(�ZXֱvq׻\�'� �"��Ɉ�qR���q���$�H�Zyn�W-z.v�h��h~���D�M���+3&��.��!.���}���m��*��j���7���T���{"��Ɉ�r�i�&$��I���Z9n�W-z.v�h�;���!$��܈��a�B��[�헏[k�{�����/g]�����
��F�]x������w�%�L@vS��M�L��@��ʄ��������ws@�yn�g��M���iǠr㊐M��EHrL@r��	�������^�M���]�7 ��Q;���9��|7$��y'����$�H�4r�hvנ^��;����	��!�6[��N���7����<�NN5�QSE�݊��v�ݸDcz�qY<���&�&�MD�� �^��z�۹�^�M���UX�:F�0$���@F8�� f�-Ɉr���Y�1%�
L�/l���YM"UvנZ[��r��o"�,'����`����c��͂��ey��R,B��*�@�;���Vy�����	(
� ����|}w�kZֵ	�dԸ��f��v)�N^XzS���;�&�%����̛�V1����l�sW�ӡ%C�ޮ2��}��wd;,'=&�=�sN��qZ�V�M�(bڈ��m���z�n�;J�lm��UN��Pr�]���	�N��ۂz.7�ô���s�PAlnA���g�*�6�l�W�Y<��u�ۣMm���;]:3��d8�5N@��vf�k=G�v�7�n՚̒�Y3Ν��
���-N�K��n���ٛ�����Ixpnm��DؠL�tt���/l���Oq�$�/�5�����f��iȦ	!I���;��hvנ^��؃�q���$�H�4��ܘ��T��l��&m� �hj%4<���t���>���f.��h]EX�:F�$����T��qR���� ��7�t�Q��]!���q���m�' �ۓ�Y��^�*�����׻HG ^� �b��T����D�P#_�s4󲚳7��b$�Q��	@�ҡT��!D��>h9ɗ��7$�2�s@���oߒ/r�f��1�
E��� �btqR��Hװ@mAb���L�z�۹�^�-X�kP��wf���355N�P��ꕁ��Z�6gr��}ݛ������`(��A�?7�֯nY�@(c���;UW5�8��[�Lk�q��u��m�=��H��L��\���n���[������"h�i�pQ�@��ɿBQ	%�2{5�Ձ��Z�9��]��!#q�^�sI>�߶na �D6��������P�\!�D���ݤ������}���rb��V�����E$��b�G�즁��1�ȩ���/*���m��z�v���@a��C�h�nX� ��t�����1&�rbq�R,C��>]��FEH�T��^� S����fY�w�e�^� 9+��#qR�{\��Gq�r(�
`�JL�/T��^�/�bu�T��XWjV_��$�I$��즁W;^�y�tܟ�A��,@�`��|Ey�f������h�i�pQ�@�����ҧ�g+�y�*@w�`�������C�T�=������4����<�.���;3Ӻ)zy�$��N��3k{N~��ȩ���� %�L@�����\���*����Z�K��ə��`y�63�Z�J!&����̪sUMK�&��iX�֖>�M�^IDL�����Z�;�JG���r���i�TXy(K�B�V��`g���;�j�УЧ3�x���'꩙M��%�K����-X����\3�����ɰ-W�t>����A.�B�������H���t��@$HA��0!�Vl	A<A�"A"��R(���k��H��s���'�ʿF#0	Ϙsh�C����I'�F@ ,��LV���HClc1$B!! B0�Ii�$���'e�Ӗ���@$S��3�q4DH@H��_U�*}�DҼ�of��P4�.�Ȓ����l@Ä��1X;��C>�7���+P�`� ��Z����	! $t� �2,1 A ���	���`V1X��BR�y�8q2���#!cfaC�<@���I&��z4�����}m=ֵ�Z�       � G/Z�����VW�*��cH��'[]mmԮ*k���ڬhPe�*�����8���E8�)MJ�s��MZ⋎!ջF�h\�Ǆ��Xy2����(V��TΉv�˰t�����q��ms�%��]�]]��ݤ
�ت\́���պ�rn/�m���r��RO�v1��"�HM����c��vW�4P��p��cZ�`f͝�wNW�gAd���iĞ�+�$��N=�<ln���[H��[s���Q��]���fEe�C�C�{n2�j�@������n9�*��L��%mc�k3�����m&�@w29�0��Lz�ӬA�V�=��LI0��prnz���#<A�C4.'"��qs�KVYz5�]�YM$��%Y�O
�R-\�-1�,�Q5uZ�dLsd�0�>��f Ւ�5V�������V˞Ŵe�f�<<���7l��d�s �6L�v"�W�\���e7g�W��_�{c���Z2]���� cn��-N�Ԝ�������F�@T6��4Db��J6i!�Im��m�s�t���NC�}��^��qAn�'p�IX)]�i�y�x����l�cv����#���1�\�;NWI]�3lv���$�:�{ñ��ﺳ�U�u��\y�!��i�n�+P]6�w������,	®1F{r8��7-���ә��`�z+
�n�8##/1��J�#v�uE�N4ݥZ���ݫ:��z�m�wb�#���8w4�^��r���@ܭk����"�����BtR:W&BUf1�(�U�`�Lv�v�m�B�f��1Z����N�)�PI(8����m�M3�Y�Vܶ�샲\涎
�a�BU@m"�Be�s*P��n�Wf�8+�e^��#�k.ɛ﮾S��Nny�WNXvU���8��=�8���u)cl#s��Ή�c^@�����M��mÔ�E�V^I��Sa��D.�;���{��|�&�-g���* lA�b;��K���kZ�-��[T!e2�jL[H�̥���4�9l�d�':w:A�wT��!y�O:E��o!��v�90�)Β��:�gMJ��i�KF�(��j�9*��1�<ٗ81�n��M� �k�ю	N�qŀium�G8��J��IL�-q���e�np��jr�12nFU��S�V��{mU��i��M�'v�`��mͺ��d�I�*p4*&I��	u��\h¸u�����=[[ޝ��uۮ�V��\/Ԍ��3m4U���7�o���߻�;ٰ@Krb��R�a]�d��q�I��s�Sf$U�^��K��^۹�u~��j,M������b��R?�}U����j�o��O �H���z/K�������]�zp�0xyXė�	��'d�{6	m�@v2*@q��׋iܡZ���7bɆ̂j�ޜ�y��8m�O��̂Vm��f����q�U��� %�1�ȫܰ<��@O{pOi�RJ�n��MQ`c�rn҈p�I���*�M�M�� w��z}j�>��X�V�$�.-��je�NF�HjG�w���^[4r�hw��:�B8�#"�ć3@/$�{6	m�A�~��HV�F{�c�$�d�M���{�4r����f�[ј44�\ �r27&#oA�;guY�6�v(�f�������L���עY�%8h�l�9˗s@/.V�B�\\���i`k��=�TL������@w��������� ߷� ��_��IL���S	�KrKq4���{=�9̬,��^:��HP�R���P�\�[��������ʜmK��r:B�檪�ВQ�%��X�}V9r�h\�g�o��_z3�ŎF�Ufn��y�O���T�p���{69cʜ�dy�1@C�M!
>|j{g��n85�;7��M�v�Ր�Y��߽�u��|��)"M$Ғ|{���^[4r�{?g�<����^�Ia�0X� 	�5z�����=��TT��Xg(�&8��@�I�s�S@�����{�mX��X`��g��D�54X{�)�{ޛ3�֬32������0H�jP�,@�V�x�P�(������s��5��F��#���ʩ絛����7����$�d��<���3�3F7/O7[�{;ѵ��U�=��ls���#k�^��v��������y�������l���	=IR�ѿ7�9"iLLrM�������/{�@�}���m�k�b�b�N,D��m�9r�h������e�V��rD��rh\���m�y�M��zhn/x��
�N��Ұ�ʰ<�G#���� =�z��w-X�� I" ���?o�꾎�Q�bfBmV;뛦K�!	�Ev������	�i)7k����	�5�歮5� �V���"��G��_UŻ%�ӫc|�0��9CX{8Pރ�w�]�v����3��Ob�r��Q�/,K�f�]�$�M)\`J�.ʅ��{I�4.5\֝��\uq�=a���a5n�ڃl�,]:_$�USx@g���u<��ƯGw���w�w�����������f�i�es��������{v�n¤S	ji7(���$�X+�M&ڏ�"����'�h��띻�����=�z�'~~M0nZ&�54X�j��T�$�P�`���]��W1zAD�M�$�9���m�jK�)���,wv�O���S�&$��Rf�����^��@-�\�=�h���o"rFҘ�&ܚ9����J�ݯ���V��VϽC���˜�ڷMbz�n�_<u��l�cy�|;.��ut��ص,�����N��r����n��{��#"�$����pd����k����nX�n���w-Y	�@�<D�N��&w�krN���ܐ��U�$�6��B��uJUU'CdҰ�ڰ9��;<ٻ�V7�`s����M��'&��.�_- ��Ձ�t�\���
%��ʭ�ީ�z�4��h�D���ͶfVm��"!dwt�.q��ݵV�o������k1�)�)UJ���mT9�m�U�� .'��ث�6:��rS�����s��YE�������~_|�ffZ�m��Wq�%�Ko^֓m����0f����,s#���$[w&�J̷�Y��o^֓m�����}����m����o"m��LLrdԒ\��Nr�~�k雷MU��Q�o�����OOP�)� =���o�Ü�����&����gi1��NȾ�%�ВJvv��m���/�m�3-U���Д%U��|������=.�.��,d�TU���3��ob!'��*���2�]�Ƌe&�%�e���Qx�H�Q!n��s���N�宓�y���ѡ�7.�͹�Hv�[jF)1�G�3�I[v�K����m�VS�J>�m�tߗ�6ل��	���'!�$���>��fI���Ԓ]�O}�|�J۰�6����M�	5��8���$���$�֗����m�{�I%�/��$��&<j����J��;m�BS<�7��m���m����?�m�ǲ=T�Q;�y�]�m��>�e��X�ϾBE�rjI.vv��m����m���I�ͷ�Dn֩D�Lr���j�՚�k�0�I�\�3΀c�P�u��ў�W�
��\�f2a[_�����K��-I%���s�$_ORI{ҵ����8���K��-I�o���]�ũ$���_}��?��b���JD��ܱ�]T�m��{�I�Ͷ�e�R�6�e��䒾��jI%{X�G�dN86�>�$�m�jI/�;W�$�]��I%��~ϾI"���&�x܁�Ԓ]�v�|�^�g��|�K���_|�o��E�ۈ�Q�������l���.�2Gg�˪h�ڄ4gmګ��&1�\�	�?��}۾��{7.���]��݃a�ݶv)�a�x� �l���Ө��*紵���A�����`�*p�r�[%�����u���
mL6#��a�0a^j
V:��ۛi��.��m��6;N8��Eݤ�vݝ��i	M���r�>�/9 ��1�����n1s6�JJ*��M:�I-_*����T�aH��w��>�<N��ql�E筭Nh��rs����r�;�=T/m�;7d�����ߩ�	}m�>�$�l�|�J۾>�$��O=�����֤����}��6Ҿ��RI[w��$�]��I%q�02"&$��g�$��-I%��i��ٍ��<֤����K��޷�Ln`�nE�/f~n����I+�<�������|���[�N�m���j}@MI15T�*�����Ucv�oR�n�s���v��|�o�m�$��\�ܩ�����i��^���;��rpvo�v5�l�����r!�L�&�FD�I%��}�|�K��56�;��В�%��U���os6��uRf��\֥���[l��kp�"<��"����j�(|���� �$ `T�S	*\��E�H+ `�T���6T9����-�rvӶ�w3��ڢ!)�oe��JfH�'2jI.�|��	v˨Կ�~��BJUWw��}�m��z����c���`I5��4���/e&�����o�$^�*�{
""&{������g$�.v�L�USE9�����;�����ԡD=�Ҿm��=���$^�MI%����I6G���4��=��n�xy�Ԋ��B��\X+�����:�(EbҪ%I-����lܭ*�m��|�fv��DB��9T���ߝ��������-ٌ�V�����W�$�{)5$�ݷ���/n��~������9�����G���~�o�|���s�Fߏ�}XB*k�0Pt렩�����,�׆a# 4 i�q�LR��@, 9a$N��C
K�	H��A�CTd �� �!E��`E���2B�(�޲Y*!�x!��NA�� c����1cV��(�������!�l"DGp�f�.���D6(�iOM��x|�*'�ڈ� �l}�*</��ۤ�Т�z�����x.Ԗ%
5(�i{�Um�������������j4�Ӑ���~o���}�I�ܚ�K����H����I^��0�4�ŉ�&�}�I�rjI/gn�.q$�Y�jI/��g�$�ӵc� (#p��i��A2n��k<v���R]�۝���c0V3��m��rNdԒ]��_|�E�aV�o���y(�{M���Um���=�S��Ě���}�I�ɩ$����|�E�rjI.��>���^V6�oÌ�ө������������̺-�%	z��}~>��߽��m��D��RKs#���/7�{�jI+}�>�$��Y�.������;v�>�$�ڷbxG�6(�bnj����r����Զ�~���}�ߗ�6�̬�m���(����S�NfX5TR���0���m�=�W&�R cL�ۣ%::��lq����}�c����b�z�_���Y�$�m�>�$����ٟ6�����Ib�=#XI#OCN3RIs���|�J�bԒ\��}�IWn�}��1���o�1�ĥR�����Ͷ�ki�m�s/�z�Q-�{�I%���g�$�ր���m��uAN�����BJ�3���Ͷ��]�k�����V�����u[�`	5��L�|�o2�����D/DB��=���������m�y���嶀�B1U �|U���W�ֵ�kZ���Z���S<�)!2&�^f3�F�u��O;S����kql�]v*99��q�\l��m�)g�<��=�۴���際��_�΁��K$���9����=���{mnt�nq�V��c�����0\^�c{�q�9; 7\�γ��� s�ݞx�����k�<��p���q����}�<�;��a�㷱���d�k�f�ǞLlC���c�&��� i2�×-�jK�p�3A٭p�.�݂^�t��L��n��ڞ�ѩ�7nͿ�{��q�ӑ�8(bV�� �����ϾI%l�jI.r�>�$��a�$�;D1T5$�%U/�m��YN�%�̷����Ͷ�v��|�g��(�2���E�9�2����~���? ��v��f{�ߗ�6�ݭ�m���x�0xL�k�/�I%l�jI.�߳�m�VS�ޥ
&{������kql�7#��I6�5$�{o���%�߿c��C�]����$���I��^D�1��
	yo*��n��@ۨ���K���y��v/��Ȇܐ���RL19������;ٰ@rH��}\�o�T�:@��ͬ�*T��敁�eav�Z]J�J&��� �Se�?t��� '��H�T��;���.��ͣ34@rH��ȩ��'� ��u^��؈����$�4.{��hO*@q�4%U�I�@z��(�׺gمỴ�m�H�l�*@s��h8�g�1��G<�2qdDaڀx��ȚР�Y��7Diһ����~�>,�dq� PrI���x�>��h�e�Q��m�{)�:��Iȩ�Lu��EH�EH� ;ٰ^��b�\�(���$ۙ�w�����鹵6B��j������w��rN[�������H��������T�m�H9 �}__}�r�e���6���rf����h����ﳀw��n*@8�(�2�m��w�G���V�����kq�M�������^���7��'��X9�I3@�۹�}m��;��(�D(�����_�Ir���F曧5UT��2��Q
l�͵`f_nh[w4��0@<VAdL�e���Z�;��6J!7��j���ڰ>�qۥN�ML� tMUR��JC���ܓ��vnIϾ�f�M�bEB1DW	D
�����$��%T�2�˚VgrՁ��"9��/��͵`w���˵�NL2<��	�8�'�agpc��W[�غ�\�f5懮$'ZE�fK�}���u���(��1�I��|=�nh���{۹�v��ho]���RL1�@ne���Z�y(Jd��Z�7��Vٙj�D&æ��SJfJ�.i��iX���T��R� %]1佺�Z&�:�V����X��Vs2Շ�1[}�h^��ף�����7&h�*@~���޾$��*@*��b�����E1	@�X��C�5��|��8ں8t(�{�P���ݒ�������ms.�"��6NSC4�����u��JuN�X5�����������܇��P{����}���l��r�.�B��֋[��a�x�C����>.-'6���]E�7GV��M�1���D�+=]k���2�k������8�m�M�*i�Gm-������۞L �E�J���~{��{���i�on�멎��Rm�&K<��=on5������Gd�9�ӚP��ww�?m�o�k^�:������ ۊ�H��"�r��n�nH!�H�w����߱"����9����r�����$�*��S��^m =��HI ${n*@:�\�D�o$&$����۹�[�M��Z���(�)���V���)�i���f�y��q��*@H�'rՁ�K���x�Y6�sM9�TLӣ6���l��o8�e����H��nvO���m��9��4��΁����s@��s@��-~Q�����Ձ��>t��D��ִnI����b�1bH��lTb����j������;���6�K���kqA��3@篷4{)��%{}��{�ۚqs���2	&9)랋�9�HT��U��ܤ�Q{jH�pCd��@�;w4���_OOr�}<� �� ;}tdۢ�
עS��j�.g�<	v7������K�X�#��ƞO������ɍ���m9�}}���qRǰ@>�� ��J��w�3J��sJ��;��T6n�i`gsmX��o�1 �����l���n�i`w��VQ	(HQ
�	#��BB��99v���j�9��	��]J�4�uSE��$�+w6Ձ�w-Xy(�������L�t��R�T�R�3;��BIss~_�����v�hw��q�9��<P"��� Ȯ�(y�۱�]ŷGm�cv\�+�mn�����x>���ĜYIɟ�_nh���;�����s@�.t�c�&A$�"�;��/�	y%
&M���}��`}����R�pr8�F�O#p�;����#�U_}W}���OZ<f��d�L�2敆�BJ����nm��>�=��M���@��T#��7���h���+�"G�$4�h^���	z��=��|s}j��w-Xr{�ZIC����ଭ���rWY��$r�^�4�,�4;R�jk�:+�˨Ұ3��vyܵ`g;��D(I/�s�ۚڏx�ڏqD��;��W�Q
!D��o�X��Ձ�Oqߡ�ߖt��0�!�L�I�=}��}{uY�I(I���;�j�>̗.ri9c������VQ	�s~Vvs]��w-XyB�����X�/J6�ҪT6���@>㖀}�R��H� 9���a�>D#YH�$�KQ����|f�e�v���h`.�N)pb;
:���c9�@"�! ���#@�Ja��"m3�l��ݦ�n3@}ׂ;�LEa�l!,��f��
>�xI�J��(k�l�h��3A�C �����{��;������wO�����N�      m� �n�h�I���r���`tדe��8m�����FKt�Di�t��H&F�v��
ϲ��+\���1Q\����p-j{]t�f�M@"�*�� ��D��Ybs.��47�-�e0�4n��l�9� v�P$�ˋd�ܽK˽h6"#v�x����Y���I�A���p� ��Z�1�4�X�IƮ6�t�l�X���mm��Kh�ět	y��@�DEH��)�X�����`��j��c�qπ��CO ��1�F�6�%g�[p8��,�Ȏ�x�ɞu�ې��"�2j3�o��諹���Oi7lF�ˤz�p�[��q��d�7�Tڽ��b��SŪ���=Q6��� WT��L�85�pO/6�Q���)l�D<�b�����a=�e�u�S�90����Pp��YcU:'�ML�dR]��ruej 2�zK���"!�md�iz���[i^��g���5q\9�m�e��m�ܑK��\��p�*u�<q�Qr�q�;<�q��cr:���/[z�H�غyvUz�[ڕ���܎y.�56e犜�-��*A�U�ur@k#<L�� (�v�il\�1��v}���0�Z��'&�v�zE�MTqX���s��q�I.�[�rJ��goV�eEZYŀ ��[�:�qd�P-j쬳�îGv@B�nU�{5�ä�٩[km�v�.�v4l�!\�E�烴|JDN��+��@$;rm�1wm�U/��` 1�N"�=��N��8�5���c	����l��ޕ����SH�^9j���K�S< 9�����-]@U$}�˥\$&��ˢ�>�8���{A�������vb(Hj)2:�m���UmWU UR��n�%Y1�%j��eW�VX����U���I�V�&���V��s������a�Dp��qv����v��ޓ��@�e��' M�I��j�( ]�N�i��M���Kl�5sWZ�xp5�Ux��||��hx"�>�x��j �"'��(��L��Zֵ�[%��f���2;rsc���c��׵>%�Je�$���[���v�y���n���؏Dx[�Uy�v�2���ri{�b���W���L-��tU���S���5�G[7ca��]m�M1�[o3n���]iB�ȣ���:.g�l㶪�km�	�ろv2^}	�<s��)�mκ�R=T$7]c'1uz.6��Ql�qp������;�{Fw/5���N���=c��A8�5�9�gD��t��Ӯ������V�}��⍤�r*ｹ�}{w4^孈���vs]��8I3�J�LT�S3�HG ;T�}�- �"�ꪫg!�\�%��)6幥`wsmX�e4����۹��ٍ����eH9�a��zX��V�ܵa����4�E�bmG�8�#p�;�U 9T��qR��s���ɶ��m�7}�s��������H�^zݮ3Ϯy㎑xY�`r�;��{���o��۰g%���?������9h� I��ri9c��UT9�V3�j���쏩B�I(��*#�,���7}����j��q���2,�I�L�;�ڴ�2՛	�nm���j��q�QT��Ӕ�e����a�
f�����ڰ9��Vي�_-���o߇� �&����HW��ܮOZ�EH	�/(�|���������K��(�s��+�Fs9�J���8�T�硍���7 ;T�}�- �"�Urþ�T�'��LldN#�h��[���/smX��V�ܵ~J�3Q4�˩R�5Ni���V�ܵg�
��4�X� )"#��*'ß���۹�Z�A��F$���ݤ��粒H9�H�r��*@Z�N���8�I���s@���{=|�yR��H�O����m�(amUA��Ntp^]�v�QS�.�MN����I�i�hnNT�r�8���}$��Y�@N����}\��T��۞�s�)�6��ȴ�����Ďz�s@��ڰ;��;�l�eL�3�J�J�������T��qR?UU]Ǔր�T���ʜA#�x�i9��n��w_M�>�߶nO�y��[� -��}�C
Q�b | P������`��ԦI)����<�@>��u�HG '\T��?�ӟ���-�-I����z���4�{[��=Y�m��>܁v�5 �c~���7�vn�L�3w3N�����qR9 ^�@;�p��	4�#n׷s}���H���4�<h�S@>���sI8�$�4�w4���=��g�_��z�s@�1�*��&@k���:�K@r8�����s�� -�~�<b����Q��λV��qR�EH_d����W�w7wwwK�ˬ.�.�5W<T�vu�
&���w��1�k
�3�m�ݭ#�l�m��8��ISq�\��^��xƶ�Ɲ�n���v�Z�D"!*�q4^�;@['Yu����s�"{^��Ւĳ�0bxf���u��ps�T����T�	jB����Z�q��1[��<;mۊu�m;bݝ�q�t�z3�8',�;���	ud�usY���# �9�9�2�����su���s�N|٢�z�q��/nM������`�g�5)�n�k��{L�l���̵`|��>���J!G$3g�vC�3�i��iR�幥`s�����}ݛ�;���;��|�$�C���&�D��<��hW����i~K�� ����'�5��n���꾽���*@uȩ�였��F$�6�Z9۹�{33?e����]�����Z�
�I�̡�ڝ��Mm���wZ�z^�oM\�ݡ�g,U��Aƒ�bi���ɚ{n���d���z�B��w���ꗠ�m,�Y�Re�u�rN_>�7�Ȩ�T��ϝ���Z�;��W�DBJd��O���ԃDM4���/���Z9۹�w��h.Z��H��`ǐK���}UUm�r�{ʐ�Ɉ�r���9�K��SmKsJ��3-X�%]��g ~��@w�*@q�fV�^��HЖ�ܦ�V����Wsnxܷ68��m��ۋc.���Җ�yI����n�m����`s'��s�kbG�3�����j��
"18�Wڷ��G{}��^�ڰ>|̛�QP�D�y �ޢdܴML��`fo�X�e�2���}��(��yۯ9��y���`�K��$�$��蚙�VQ�y��)�~� ;1�A����H	+/�X���
T�uJ���2lD(P�v�o�7<� �"�:��zn^�����=u�nh�p����@�=���dz���MX��ע��G�9�4�HN=������`w���""K�}ݛ�ҦZڦ�)T6��v9ܵ~I�3vՁ��ٰ9����"�l�>��f�]M2�j]��OyR��1ْZ�qR �L�*e��9NUH9�a��!�{�6vw]��w-Xy�ВD&���!�#D!�V��p�T� ��w��S�ܸ�&��Q�Ǡr�V��$��ߗ�fnڰ>|̛��K��9x2�O����p𧎞��ɶ��$��7�u{s��2�Ue۰'fR���느ȩ������X?g�h�4�z51�8�nL�;�w4�-z2s��w-_�"^P�L��_�J�by2d�����=�ڴs�s@�m��;����@�M!8�=���}o��Z��H�T��U_q�؀�ҦZڦ�R�m4�s�j�؅
�$�����^{�`s'1�Q�(R�T��"�B�@�Tj�ww��?��U�Y-���L�mI������B��.���P�];��)�u�o;��ݖNN�MG�m�r�;n}�GYƙ&ɱG[Y��Nvڔl8�ht���������v�n1�z�n܎b8��З.H-�9|���Va�D�[)p6p#��I8�Ɣ:�s<j�sNv֜��&L�*��z�Gۨ�j��`6����{�s���Ͽ�ww{��?=���x��v����ڹ��K����s��Wl��	֑z���y#Km�.@���$�T���L@vd�������*@)�cc�6���s4�-{����ݝ�`w����2��B�è��	��%�z|��s���{n���@.���&�q���9��H� vMAꪫ~�z�w���F�1���ɚ{n�}�f���V��v�h�L��Ʒ����Pԝ�'�nv]�-v8lk���^��ι'$��{�ww_����L�2LRg��4Wڬs�kоa�ݵ`fk��`���%��[���}��w=X$BυB��(Q#Е�ms����V�3*�	$��ʙkj�9��*D�;�ݵ`w����Cg{�Vvs]��|1d�S&D�D����s@9�f������
#�'3���{�d��S�T��sJ�9�ʰ<�!(��k��vՁ�[��s����&�H�&�"Oiέ0ͼJu/7���l�R	)4)D�R鰧�!���6�x�DƜ��?-��s@�-��(�0;�ڰ@.��2nZ&�o6�슗�����T���ْZ �+O�FcN%�4��� ��~��˰�I�Cݑ����"�Si�7�@B�ڱ0���L`*���&@�k��"&����l���6��A�J�]9�� F�;B0 ݦ0�X�q�	��Wܚ������1� �L�R�(Xx����`B@aBD���6Z�xm�R�.����+ŵ�Ss��B��8�ԑ)���A���i�|� O�Gi��	}@xQ|��.�~���q[�}~ CE�S�TL> 
�Q��誛���%���2~��vs2Ձ�)x
C):���R�ԗ�s7�`g��vܷs@�m��;ʥ���1�"1)5َZ�7�r�~��ɨ����m�wOD��&�跎lc��s�9S�t��;r6ص,�ZU:����f�;� dT�;�7�r��'��}57��:T�����`w�����h��h�n��?$)�cc�e�V�^m �{P�%�;� �Հq�*�sD��ҙ���}��v{�j��s-XT/�CDQ
 ��� ? '���Cj��|��`���1&�q�"�9����̵`s2�d�;b"D5�q�u�g˵�%'�E��Twp�]���j�^���Q盶�Y;���s�ܢQ��U�=�ߕ vM@vd���\T�}����Y�Bd��� ����~H���s@�m���H�mzH����ɚ��;���s�j�B��7mX;�4�ck,�dɐK����ٙ����X����fU��$����9��y�B�2$����;�w4�[4d�;��Z�=�R��B� ������8���XrD�u�%ȽY��ʋ��BXȕ���k���#�5��;u�٧cu�mБsn�+��9^�R�l��:��,ó\�i��=cV}��M�;���%�,����cc�'�.��:ݦ���Uǈs��=tq����V���r������Z	93�\�<s�`�5��-����Ih͞v�ݨ�����ߟ�����������)����O�Lu[�S�lx��M���okI����w��}���8���B�k����;rL@w�*@7"��:�H4��(�'$�8��@�3-X�e� �3*��D(^P�BS!�?�� �X�c���nh�y(l�wj���ٰ��2eTҩrꘪJ��a�!By��+ �wj���ɰ9�w4������&@i�L�rM@{ﾯ���޾ ߼� ܊���{mwn�iN.n5�s�dK�����:b�j^�r�v�@�,.��u�YswP�%�;� 8�U���X�ڀ��mg�ŉ�d�%�qh廚�fp�UCb�������f����>��Zߗ�Z�� D�9���{&����wٓրnyR ���Lb� i�'3C�1.wޚ�v9ܵa��3~V�`f��[�);�ڼ��-����7=���ʐ9l��_�f	�?��3rdm;����s�ͼ��ݮ{��L���z�v{mf��̺��3w8sʐn*@욀�w���z���!�22I3@����#&�8��@w�*@>�\��!2R'3@>�,�;�ڴ�~���3?f6�۹�}{w4���'T�c�]�Y{����z�#��~��"��`n�L��I�2R�Ca3N��\T��}�Or��Cڀ}�-޹o;�N1�\֝��`�|&��)�͗l�m��D���c^ex��\b���-HG FM@>㖀�\T�+����<���hץ�x�V��w-Xgr�ꄒl8,�S�MW{{W�n�#��@w�*@r8� rt�@;��[	��Hq�"�9���$����rIϽ�krz��1H� �) ���b+��(I.��Z�ss��N��K������wv��*@���}�-��-X�!,���mʦ��334Lӥdy��B5��}�I��{R���U��<8)�������R'3�z��x�V��v�{>A�_nh�UIz)ɓb���9h��HG FMO���̭����$�����>�f@���{^���Ρ+�q%�nf����ɨ[s느trV6(���$i9���f���k�9���rN{��7$P�b�b�F
��{�l��-��J^�\®ksql��,�//T2��%d�6Vl�{����lc�t{vsS�i�*cQn��1kr;�n�u�v�d.�,��Vyq[7\��i�x�e;�s�[�P���v�v�nn�!�Gl��K>��P
/J�v�h&�-�4l������p7���pfݝ\�Z�����t��t�,�������k����������b��u��ޮs�<�lu�EN�:���L���8yrMw�$�"̎�\�p[s느n*@���T��6���@���hw�s@9Ζh.���?$-`ߜ�8�Qd�j���ݵ`�L�=�o�3f��nڰ>O���IL�A.�f����C|r��r{r*@qȩ�;2G$a16!HI�qw��v���۹�s���׆6Ǫ4��D�ic��Cqإ�����ʙ'a)_E���ԫ$���1�Ɯzݷs@��ՠs�����@���P��J8��6�+��c���	r!,�QaYO�:�+�>�ô��#q���F��@>�^U����٪!�f��;��8�D"&%�!&����@����y%���P��9��|^eٛfn��EH�~��{��O��n= ��`�I<��I�q/Đ?(�{ev^�V�n��6�j{^��؃����,��@�wsv�x���P�� 8�Y�}����2RI�s�,�UU��Ob��T���-�;/&l̅'21�V{�`}��Vq/(�V����NGN�����#2���IN ���S��s�n��?��m���!&��	cN=������H��� w����1ϯ�FMI-�1�.iXvs��!z!B�o���*�����m��9����&��۬����q�V��vp�^K��r�y3���l.KԔȆ�ɍ29hl��"�s��{�`}��Z�!$�a̝�`��dF<��!&����o�G/���s'u�9�*�"M�@�͢���[&��R�9����9��BQ	$���`v�nh|s��?6,rI&hu�; �:eX�e����C���!�A��w�~�����m&����H���f��۹�}m��9�j�9�}���(��p�mqtWn�im��C�+��]�͎3�Zw:��%�4⑸$'�Rh���V;9�b!B����j��ڙkf�nd�.���@rH�גZ }d�;�j��l�>���cR(D�+��� >�j�EHI �dr4��#RE������@���4�2Շ�B}��v����mURooksou�"�$��y%�7s[�!�O7��x�@R& �+H���Q�@<�R��=6p�p2�W�M`8�͚�)�267�GDXI!�1+�#�Pڅ>8���<x�MP����TZ(l'�ʙ�=�ދ�9��� {�T��|�isϼ���<`�JkG��5���a�R�i�dIʚS�#�̨�|r�8<r�y� ��]�dj4/'! ��=S�@��%BE=�q0ҌA�T>v�ImBD�G\����w�<|HċX�>���kZ�@      �� E�h��]�@m��*^�䕖��V����㍛G)�a�S�^d9Zj�۞�����K�5VF��i�c)HOF�t�DH[�G��vIj�j�3�-l��K6Z�085�ku&իh�H`n�ۙ��qX4�����n���8me��^c�"y�+��	g��]��pC�\v˝1��a�(���!�#�k[&�s[\S�3]�;ce5�@n�R�tNz�{2��($ݝ��cd��G��Q����%��b�h6ض���h�s�g`���p�A�`a�%;w�m�m�`�ZMTӀ;mgu��݂[�N˲���1VF�7Y7X�;>!G���x�PWU�[,�z:nB�'9�lr�#j%�.�N�j���y^��-ٲ����]��O]ь�T��bGs�fĆ�1�1��ȏd�+��V�P�rm��Ke�`���8J�S9Qzx��|	�wY�#���V�ۏ(�TT����I�k=
c�ќq����wN�[Hy��u3vݟOr,)Vv�p1\��c4�b�n`�����3��bMĭ;��,�o=�@��E�@ΫY�SmƸ���#�:�dvy��5�g[�M��tR�Vu������6$�z��ϧ� t���O7��)ƈ�$�]T��AݱX�e��n��0j����`��Ce��*�Ұ=��Y�����b�m�un�&gjú�g�n�Q� 4Kx'n`ӄd�]�;,;h�I�������+�����1�G R�p�9���j���dz6z�Kx�S#��
�UfJۦ���
qۜ�u
���Y\m¸�viƲ��v�� �!I�g��v�x�wl[,�U@u���ʵ\X��a�ё��i���"Y�\�VҲ�Uj�Nc2ri�2	v���y�V��:�#Oh8q��f8����K���ڧ\��i@�:6��/S�V(mN'9 �N:l!-��̺!�Z�&? O4y�@��&��}Z;��>��b�"�A�Q����!�b)���w�u�kZ�&��g�H�├M�K�^y��^[���v��lj瞽�U��vݮc��e�m�[l�E�{�:��:�ە�����gS��,��G5�����\�󺰞n�������Q�pnY���;Z4�*�X�S���1՘��n+;ch���c��y֨��,�9e��\v�c [������6�{6�q���N&�k%�5��qO��rr3,�7�糚ѱ�����;&�秬p&��͞����v�u�8�7ld-�֫\�3]���ܵ`}��v�z򼗔%���� ]*�M�9��ic��3@��ՠw����Z�>��W��O5�[4�%PM����~�[���`���-�s��\O"��&������9�ZX��;$��cڰ7v�Z٦�l� �C@��S@�]�@9ޫ4v�hw�*�1D���3$H����D�����[�\.�$����JR��w}���b�@D����Z�z��9�)�}m����������mǫ�$�ߵ�¾���\$0HX%. 3m@�@jk�ne����~�ٌ�DԶ���dqI�v�x�>��h�h��@;��v�c��m&�4���^Ih����s�� ����g�~lX�rL�9�j���f���M�n�����[�4���EqȘ�iŮl �v�t���MQ��X{]��Z��%��w���������/�9j��9�)�}m��9�j�>G0�M���hDqM@rj�EH��������]��yg�@�F!1I4{���9ט��r �B!(J�}��`��X~\�T�)!nf�����Z���̫Q�
'�������䩤FӍ�Z�z��v٠}m��9�j�9��kqE%&(�r<O��[Wa޲:a�ɸM"F��l\�t�Y�~���|�|Q$Ģ�R|��M�n���c��f=��d&Bd'�/�)L73�f���m9ı,O;���r� �DȖ'����iȖ%�b_{��[ND�,K��{�� ��bX��{~�3�t�i��kZ6��bX�'�k��ND�,K��׺�r%��Q�Dȟg~ͧ"X�%���߸m9ı,OL�����E��&]kZ��r%�bX�Ͼ��ӑ,K��>�siȖ%�by���ӑ,K�j"�⡵�
����/�L��L��:��3���\$�j�[ND�,K���ͧ"X�%��{�ND�,Kߵ�ݧ"X�Bd'�ǵp�!2!2gq���%=-v��6 ��n9���"��*9��1q��V�{���:ca�v�������%�by���ӑ,K���w�iȖ%�b_>��[ �Kı=ϻ��rBd&Bd.Gk �t��T���f���Kı=�]��r%�bX����ӑ,K��>�siȖ%�b{���ӑ?�șľ����3f��e�ffk5v��bX�%������Kı=ϻ��r%��PdL���߸m9ı,O��߮ӑ,K���zSWV֋utk5u��"X�%��}��ӑ,K����"X�%����nӑ,K��r&w��5��Kı/`^7�R�nfY4ɚ���	��	����ND�,Kߵ�ݧ"X�%�~���m9ı,Os��6��bX�&�����=ޞ�??��Y�։� �:Ɋ�s�@����W� m����.p.�H�vA��Bc�w���1�ՍU�G�֕7B�.�ѥfRn��!����㳬�G�tCnv{ �61\��n��ӻL��Ax%��8�]Fr�]�B}/k��*���pݠ�ps����4n,˜5�n�"�<��gZ֜U�(�1�O�aL��a���qӹ`�vR2q�و׎��v�ô�3��uh�dUsطa�Ϸ.��ӵ�h5�v�g�*��+��۶HK�2��ִ|��bX�'���]�"X�%�~���m9ı,Os��6�Ȗ%�b{���ӑ,K����IL/t�2�.��j�9ı,K��vkiȖ%�b{�w���Kı=�{�iȖ%�b{��۴�Kı<����ܷR虖�sZ��r%�bX����m9ı,O{���r%�%����nӑ,KĽ�zkiȖ%�bw�^ӹL�HScR��|Bd&Bd-�ߕ�Ȗ%�b{��۴�Kı/{ޚ�r%�b6'��{�ND�,K����I#�J��&i\/�L��L�ܭ״�Kİ�*�?~����Ȗ%�b}���6��bX�'{���r%�bX�������肿�J炻N�qD��-b�sɎ����9��v�=��:t�vԦ���Y�5�sY���^'�,KĿ�~�kiȖ%�b{�w���Kı;���ӑ,K���w�iȖ%�b}٫��5ua��n��sF���bX�'��{�NChr*��>��y�,N�|��Kı;���r%�bX���Mm9ı,K�ϻ��mə�5ff�iȖ%�bw���"X�%����nӑ,Ľ�zkiȖ%�b{�w���Kı)���fgr��2��ִm9ı,O~�{v��bX�%�{�[ND�,K���ͧ"X�%����.�&Bd&B�z��V�K
	uUT���bX�%��魧"X�%��}��ӑ,K�����"X�%����]����L��Y�6$ۙ(�UJ�M)f`ג�yj̆��`s�<sz�K��E�U�Zpᐱr&��}����{��7���{��r%�bX�w���Kı=�]��r%�bX�������bX�'�)�[4��NXSn�i�/�L��L���xm9±ș��u���r%�bX�����ӑ,K����nӑ,K���~��kPˣFYf�f��"X�%����nӑ,KĿ}ޚ�r%�����  	9�@Ç�<��k��ND�,K�w�6��bX�)���R���aRMT��Ӹ_�	���}ޜ�r%�bX��]��r%�bX�����Kı>�]��r%�bX��ސ�Ն���]\��r%�bX��]��r%�bX�����Kı>�]��r%�bX�}ޜ�r%�bY�;�w�߷ch�?�W���P��G�B�՝^z�(9�i�ph9y:���7�ۏ_:|\��nj�<�bX�'߿~��Kı>�]��r%�bX�}ޜ�r%�bX��]��r%�bX��{�Y�ܺfsj�Z6��bX�'�k��NB�>��4��H'����	�<�ﴖB��
HL��M�%��T��r%�bX��Nm9ı,O{���9ı,O{���r%�bX�}���/�L��L���%�l�)�J\�jMm9ĳ������v��bX�'߿~��Kı>�]��r%�`C��*��&��vkiȖ%�b{٫�l�C��0��TӸ_�	�����iȖ%�b}��۴�Kı/�}٭�"X�%��u�ݧ"X�%��~�������N٤�-�w:!S!V8ٳ����H��u�W�Jv��\��]ND�,K��ݧ"X�%�~���m9ı,O{���9ı,O{���r%�bX���ޘ\5���,ֳ3Y���Kı/�}٭�"X�%��u�ݧ"X�%��{�ND�,K��p�!2!2ꧺ�N���7N��ѭ�"X�%��u�ݧ"X�%��{�ND�,K��ݧ"X�%��3J�_�	��	��lӘ�2M[sWiȖ%�b{���ӑ,K���w�iȖ%�b_���[ND�,K�뽻ND�,K��~�3;�L�.a�]kFӑ,K���w�iȖ%�b_���[ND�,K�뽻ND�,K���6��bX�'ʇf�ou�kZ֭�V^��n������ۋ\E�pb._AmJ�l��h�`j;G�-��R�V0tC�p��"��&�xyR��j��.
��{W�R�'Z��m�&69�D�M�\�v�+,��/�WK]�v^x��i��"=Zy\��aq��]��r-�t�)	ܝɭ����y8��b�Zq��7/
0p�κ(��5Vr�mp����g��۞^.�]���w��d����e����/�="�nݤ�+��r�]\QGW6s>t�TZ���51�{���oq�����~��r%�bX��]��r%�bX�����Kı>�]��r%�bX�{o�g�G"l5��ߛ�oq���{�w�iȖ%�b{���ӑ,K���w�iȖ%�b_���[ND�,K�)�[4��L)�U4��&Bd&'��xm9ı,O��{v��c�a�2%�{�kiȖ%�b}�_�]�"X�%���d�]n���s4m9ı,O��{v��bX�%��5��Kı=�۴�Kı=�{�iȖ%�b_'�z\2��Rk%�u���r%�bX����ӑ,K����nӑ,K�����"X�%����nӑL��L��m쪑��'A*�JR���WY�]q�����nQ��<c������j�s<���v캰�h�a�3Z��r%�bX��]��r%�bX�����Kı>�]��r%�bX����ӑ,KĿv�����32f�����Kı=�{�i�qO��#Dh��<|TW;��K>�{v��bX�%���kiȖ%�b{�w�iȟ�ʒBd&�͖L�]D�\ʪuT��&B�,N�_�]�"X�%�~���m9ı,O{���9ı,O{���r%�d&B�&j&e��)a@MUM;��	�bX����ӑ,K����nӑ,K�����"X�%����nӑ)	��;FKjZ��'H��QW�ı=�۴�Kı=�{�iȖ%�b}��۴�Kı/�}٭�$&Bd&B��{҅.byNeʧ4�����]h�4�n��
n��k���}�\�����n�����5sL��5M���p�Bd&Bd,���iȖ%�b}��۴�Kı/�}٭�"X�%��u�ݧ"X�%���I��n���s4m9ı,O��{v��bX�%��5��Kı=�۴�Kı=�{�iȅ�bX���ޗ��T�e�n���ND�,K��ݚ�r%�bX��]��r%�C��zS�8�x:�d+�p�[�4�1C�	� &	{��M�v8kDY�i=���fE����S�����o��ʒsJ�`+ �!�(��4�^��b����,��,iGt�v��Ϲ�y�Oܤ��JȦ��B��
aBIIG�4�'����|�:O\l���B#�U>��x�QpTc诨 	�UO�]�*!��ށh {�D�O>��ND�,K���ݧ"X���Ou�t	t�UHtRsTU����,K�뽻ND�,K���6��bX�'�k��ND�,[��ݚ�r%�bX��w5q�&fLշ5v��bX�'�w�6��bX�'�k��ND�,K�߻5��Kı=�۴�K=���?�����ѳ�9��uk�����1g�����[]��X���{:�*e�r̹��Y�ND�,K��ݧ"X�%�}�ݚ�r%�bX��]��~c�L�bX����6��bX�'L���r���a MUM;��	��	��{�u��?*)��,O�k���Kı;���6��bX�'�k��ND�,K�Mw2�L;��&d��kiȖ%�b{�w�iȖ%�b}�{�iȖ%�b}��۴�Kı/���b2!wJz��6��9RSN�|Bd~D�߿xm9ı,N�_�]�"X�%�}��u��K���1I���~D�y���r%�bX�s�ԝ�Q-�1734��&Bd&B̭�p�ı,?s��?ki�Kı>��߮ӑ,K�����ӑ,K��ޛ��ӷY7Z;se��0���=v�]����L�p�rl/\j)�2k���DJ��WiȖ%�b_{��m9ı,O{���9ı,O��xm9ı,O��]����L��O��=�)�U4��E��ӑ,K����nӐ���,N����"X�%������Kı/����2�D�/B����˒�sY�Z�ND�,K�~��iȖ%�b}��۴�K��ș����m9ı,O�k���Kı)��S/�(�7}����{��7����۴�Kı/���bX�'��{v��bX�'���6��bX�'ę��.^Җ�TӸ_�	��	�ߎ�iȖ%�b{�w�iȖ%�b}�{�iȖ%�b}��۴�Kı<x|89��AB�B�AD
�(��UUUUr�bT�Y(��f�stBB��X�u;nb|F�e���crD�nȦ
�!�h	�!%��/���F�7��w�W��y�+� �p�vl���Y(;nN �=k�PwFvK��6n�����kf��Ψ�ӬkrgN��YZ�U���^V^��f�k9l��zÓخ�v��q�k����.�;ap���8�9ɭ���95�C��6�F=x��^�׉jH���l��u�������Y��lڷ0��������#.Y.h־Nı,K��_��iȖ%�b}�{�iȖ%�b}��۴�Kı/���bX�'����sV˚�ф՚�j�9ı,O��xm9ı,O��{v��bX�%���ӑ,K����nӑ,K���g�w3D˭I��f��"X�%����nӑ,Kľ���r%�bX��]��r%�bX�w���Kı/�ӽ.d���Y��mֳWiȖ%�� ��3���[ND�,K�����9ı,O;���r%�bX�}���9ı,K�{�����f��4\ѭm9ı,O{���9ı,O;���r%�bX�}���9ı,K���ӑ,K�����od�����:�D�=���sŬH�;;�jJ�{v�ݹ�:뱠�m���d���r%�bX�w���Kı>�]��r%�bX��;���I�L�b�=^�_�	��	���ɟK��rj�5�6��bX�'�k��NC~y���ND�/���m9ı,N���v��bX�'��xm9ı,O��t�3����&�f�����L��O3�iȖ%�b{�w�iȖ?�U�DȞ����ӑ,K��u���r%�b2v������t��4���&Bg�bdO�o���Kı=����"X�%����nӑ,KĿ}�f���	��r���I��S�(�UM;��,K�����"X�%����nӑ,KĿ}�f���bX�'��{w�!2!l�	[5 M'M��M&��'��2ɫ�ƭ����C���nZ`ڛw��T�4�K�2)�3J�|Bd&Bd,�]��r%�bX����ӑ,K����n���O"dK�����6��b2!>��ȕ-US���m�M;��	�X�%����Ӑ�����,O�k���Kı>����"X�%����]����J\)!2�'��S@�i�.f�m9ı,O�k���Kı=�{�iȖ=L?S�����7�3���v��bX�%��r%�bX�����r[35��WiȖ%�b{���ӑ,K���w�iȖ%�b_>����"X�%��u�ݧ"X�%�_>�����Kp�&��Y�iȖ%�b}��۴�Kı/�}��ӑ,K����iȖ%�b{���ӑ,K�w�����w���������9*y�,�l�r>�q6E&�n31m�0.��N��v��yY�&��Z����%�bX����kiȖ%�b}�wٴ�Kı=�{�iȖ%�b{�w�iȖ%�b}��)N�D�ї,��k5��Kı>����r��DȖ'߿~��Kı>�߿fӑ,Kľ}�s[ND�eL�b~��zi9�t�Si�Qp�!2!2{��m9ı,Os��m9ı,K��w5��Kı>����r%�bX����N�h�u�.d3.f��"X�~U`dO�����r%�bX����kiȖ%�b}�wٴ�K��w��!bV�e�����TG�A �:�{��NOq����~������IU����ı,K��w5��Kı>����r%�bX�����Kı=�������L��]���93l���S�3L'�K�kGn[u�L㇝��dY��/]�n�{Uf�it�jhM"�R����L��L�����Kı=�{�iȖ%�b{��siȖ%�b_���[ND�,K�û���r�&j�f���	��	����+ND�,K��{�ND�,K��ݺ�r%�bX�}��m9ı,J���/�H�B��{�7���{���?���ӑ,KĿ{�n���c�"w���m9ı,O�~��iȖ%�bzd�Ip�̤�2�k5�ND�,K��{��r%�bX�}��m9ı,O��xm9ı,Os��m9Ĳ!n�#ԪN�2T������V%����fӑ,K���~��yı,O���ٴ�Kı/�����"X�%��0�d"�@�ӥ��z�y��q�kY��3��Sp_������q���v�7v�l���M�ٞA�Â����\m���u��"��"��@��%788�ni��.�nsp��aR@5�����3 g�On9�K��Zwg�d\k$�b�+[��ϥ�;k�����Z��"��Xl�mY�t��C�ֻ9�{S][g�%�竏u��g=�t�Kq��6	k��O en}���w���?���`qik�\����껎lv<��eݗ�]{v��U�[4J�7c����ڭ�v%�bX���w�ӑ,K��;��ӑ,Kľ���By"X�����p�!2!2)���j��P9�f\�ND�,K��{�ND�,K�{��iȖ%�b}�wٴ�Kı=����r%�bX���Γ2SZˬ�̶�Y��Kı/���bX�'�w}�ND�,K�~��"X�%��w�ͧ"X�%�|�rw4S55I�%֍ֵ��Kı>����r%�bX���xm9ı,Os��m9ı,K��{��"X�%�~a��m�lֵ̚��ND�,K�~��"X�%��w�ͧ"X�%�|�w��r%�bX�}��m9ı,J}=��;�2���y��2#��uu[[�8g]ۮ��n�<�yn孫o2+b@y7}����x�,Os��m9ı,K糽�ӑ,K����iȖ%�b{�{�iȖ%�bzd�I�.gi2MS.��Y��Kı/���[NB!��W�;���'u��6��bX�'{��ND�,K��ٸ_�	��w,Б��R�%�&�3Z�r%�bX�}��iȖ%�b{�{�iȖ%�b{��siȖ%�b>tݫ��	��	��)�٠h��I�Bk5��Kı=����Kı=�����Kı/���[ND�,Ē�˅�	��	��N��L�"��Nr�3Fӑ,K��;��ӑ,Kľ{;�m9ı,O��y��Kı=����Kı? u�ܷ2~����b�l4�W]�6��ۣ�M�Wk�IEďb��.fzzɭup��ar���{��bX�%�������bX�'�w��r%�bX�����q6	"{��I���svM�MM�4��UD�Z�
��}��Nı,O}�xm9ı,Os��m9ı,K糽�ӑ,KĿ0�r޶�fMkZֶ��bX�'���6��bX�'���6��c�Qz!��d@IO �tu��Ob^�>涜�bX�'���ͧ"X�%�\�s3��2�uT��&Bd&B���ͧ"X�%�|�w��r%�bX�����r%�`~&D��߼6��bX�B�&�#r�K
4�jn�&Bd'���u��Kİ�G�߹�m<�bX�'�~��iȖ%�b}�w���K�q��������hˬ������tnK����m�.<��iS������W<�q�a��˖MjkZ�r%�bX�����r%�bX�{���r%�bX�g��m9ı,K���iȖ%�bw�^��4a3Z�e&�ֳWiȖ%�by�{�iȖ%�b}�w���Kı/�ϻ��"X�%��u�ݧ"~��,OL��34��D�L��3J�|Bd&Bd-���iȖ%�b_=�w[ND�,K�뽻ND�,K�{�ND�,K�=;��2�k&d̶�Y��Kı/�ϻ��"X�%��u�ݧ"X�%����"X��p�$b �`�ށP\����ٴ�Kı/��a�I���&�SJ�����	��	����ݧ"X�%����"X�%��}��ӑ,Kľ{>�bX�%?w�q���v6�r+��ØdE��R/O��í^M���9:�4Vsq������u%���Kı<����Kı>ϻ��r%�bX��g����șĲz��p�!2!2���~HK&Z�k5�ND�,K���ͧ"X�%�|�}�m9ı,O{���9ı,O=�xm9ı,O��t��\��a5	���fӑ,Kľ{>�bX�'��{v��bX�'���6��bX�'��{�ND�,K��s��Ja�蹒�jkZ�r%�bX��]��r%�bX�{���r%�bX�g��m9Ĳ!>tͫ��	��	��)��UHUu��&���ND�,K�{�ND�,K���ͧ"X�%�|�}�m9ı,O{���9ı,Ol��d @���:A���v��BD��]�#���(�GH><��v`g�|]1S�E�D��#l'�#>��	!B�D ����G�";�:h�PH� 7�� i������=WӐ4-�Ѕ�B$k�U�M���_�ț
���� D�`iI�����p�K��,�ċE��"��'�+��Ԝ!��P�6��# BB5HT4�"���"q��t�U�CЀ��	�D)�G(iG@}Q9�́�xe������FH�	��ww��������s�      m�� [zt��5ʹ�hZUIk�[��n��mv�I՚���L� ��ʃa}n׋]��l�э̹I[���ӵ�6�h��ه�}��*�*�=UE ����h��We���\$:�m�y���v�sȘ͵�Ev�֒;4�^�-��+�+m�S��)p&{uEճ^;cey�ݮ���ju��]Ŧݸ�l���Fݰ=��w��C�/g�;',�ɠ�-㇟g������t�e�%�B��v��C�Ӹwm�iE�v9�{h���֪q!�][m|;��	"Z��бvvL�h�v�gN�t4m�re-})��q��ivt��Ӯ}��L9ݛf�1U�8.��h�8�ڱ�����N
��rn.��ø������%�`��vq�Uq�Gl�W/[xH�/-&רl*���O5��[!�������;2�}�e�h�L�B��N�Ǝ1�2�Ivw]�w����l���v-'"��9�6��2�B1̩sR��㧳K�ri�l[#�ۃ�j������ ��7=t���0:��͵[F�ٖ��r�;2�&g�IrQMP�ڰ��n���um�X�vӡL���8^@�,x���zR���u��'%�ӫ��;���RS�6	� ���q�	{�w�\0������m=i����o�}����eل]UPN�*Cb4i	��m�����]�nJt�4��-�9�`ॴ��b�X9�O0nӏ9i��1�$Ϋ��-rKcm�E배�յ�h0p�#CeZ�����c������o���[B��ݬ.�8�jy[ʫZi��E[s@l��Sf�Q�<�8iz����h\-��$���6i#��	z���;�ls1�:Ö�y�
Y@�\�AK8�&��V���&U�Ζt*�UlO�	�X*���it�:�P|�jӇd��mw�m�͜�$�m����
��ˮ֨	N�vj��ܭYxʣ�M;-Bh֗��ir�v�+k���q����5.kYh��".�@������ދ�@#��S��z�>O'&��ֵ�kT�q<�z�M[�iغ��%���M�l�0��X.�C��3B����}�I����vzu�愭�nn�v��'[���t��u��v����]�:�,.�û1��N�=Wl��n;i�u̦�7g�n��l�q�n��*)�n��v��E,���9�b���s����OOU;�s���Rsۍ�k��H�ܗd�_g�c�GJ��"�.���3(��[�?�����������p�s&d�c�vhݻ����7�N��v�;�\�b���ܩҷY�Zz����~�q���������r%�bX��g��ӑ,K����nӑ,K�����ӑ,Kļ:�S�GESr�l�����	��	���ϻ��!�c�2%���~�v��bX�'�~��iȖ%�b}�w���O�ȘBd'�zOM&��h�EM*����&AbX�~���iȖ%�by�{�iȖ?��Dȝ����ND�,K����\/�L��L����;��̺�uOiȖ%�by�{�iȖ%�b}�w���Kı/�ϻ��"X���u޻��	��	��f䷢�	d˒��R�r%�bX�g��m9ı,K糽�ӑ,K����nӑ,K�����ӑ,K��~�yrۆ����.���:�w�OM�o��zu������Ep2�w:Q3.f�K
4�jn�&Bd&B|��ӑ,K����nӑ,K���w�ӑ,K��>�siȖ%�bw�N����4]�l֦k[ND�,K�뽻NCB�C�|��K��8m9ı,OsﻛND�,K��ݫ���.���y�҅5U2�0��j�9ı,O�w��"X�%��}��ӑ,Kľ};�m9ı,Wv�]����L��]S����
���Mk34m9ĳ�@ȝ�~ͧ"X�%�}���[ND�,K���6��bR!ws~W�!2!>��ItUVf����k6��bX�%����iȖ%�bw;��ӑ,K���w�ӑ,K��w�ͧ"X�%����K�&��k���f�%�svo��Gp���5�!��rjƢ^c*�n9�vn�uf��~d�,K���6��bX�'���6��bX�'s��l?�&D�,K�g�ڸ_�	��T���'�9mL˦MT�9ı,O{�xm9��"dK�~��6��bX�%����m9ı,N�{��r%�bX����{5�ܳ2�ֵ�Ѵ�Kı;��siȖ%�b_>��c��N�	hR�ha���p��熢y�����r%�bX����ND�,K�N����j�]MW.��Y��K��$���~���"X�%��?~��ND�,K���ND�,K���6��bX�'{F�!I�r���j��&Bd&A��{�ND�,K��w���Ȗ%�b~�߿fӑ,Kľ};�m9�q���~�?/��q1��[�G\r[Ru��w:rSh�v����{x�S�m�4��Z�e5d֮k6��bX�'���6��bX�'s��m9ı,K�ӽ�ӑ,K��w�ͧ"X�%��}�^�h�3!��Z��ND�,K���6���DȖ%����m9ı,O�����r%�bX�����r%�bX���Ө�]U5D��SSp�!2!2���r%�bX���u��Kı=����Kı;��siȖ%�b_;�N�f��3D�h֦k[ND�,�(�"g�߿kiȖ%�b}���m9ı,N�{��r%�`m0��@*�}��#�=���kiȖ%�bxd���@�3.����_�	������Kı;��siȖ%�b_>��bX�%�{�m9ı,K�~��~��]���-��XϷr<�h�S���v�l=�WZ6R��mעBӅE9���r%�bX������Kı/�N���&&�v��;���L�D�T�JtS�tT���3*��&�ݭ,�m��k�/1�1,DL ��32��9��Vj�Q
׻�`�v�
���lY$#0�AHh���Vנs���)�|�Պ�2cfL���ͤ�*@빨	&��"7$�)a�#ҥP�;>��d�im�����M)�M�;J�l�0rm��8�%b��o/�/���G�1m�㱭�#��vX�&px��θ�*�X�m�NR4n�n���f���%���!�ˬh!��v���Wev�e�;Uvzʍy݌;��%R��� �H��']�Oj.9�4��/;m���M��۷63�몁,���L6B�&gF���lv�ݵ�o��{����)qӴ�vי^{rcG����mٲy��`a[��{��*�Gk�t�a,�U;� �����`��RI G�s<��̉̒)4l���m��33-X��ʿCf&-�{�jf]9����*@I"�λ���l�w�*F&�ŎBH�m����e������$�'7f���ЙzMT�"�ԎL���f�m��>]��۹�w����2�G&��$�:��ct�|��
����f��l���=�/���ɂb#�M�)�|�k�-�s@>�U��]��X�Q�B
C@�v�WU����0�"�λ���l.+r�27�I#�;��h��@��M��^�gs��7$�cW��f��w5�6[����}z��,O'��̎)4���9nL@6��w5�(�2V_9���j㎓��q��I��hYز��I:��i�h�S�M,m��p�>]���� �]���\�ｾ��0�nQ�9	#�;��h��@��M��^�Q��\�B/�<M�@>�o�ܓ�}������Y�K	���P�v!s�?��;̬,��K��m���{�I�@rܘ�m�9�f���n%1�E� �4�m�o`�9�sP�`��ٕ3p
�X�1�n��S�-���Cv�ãn.^&�&f�#�n����l�� u��$� 9nL@�ʼ�7$N���4�uY�}l����@�{)�^�b�2b�I��5�6[��� �G5*Âɗ�ܶ�eӚ�,6"!�{�6fWf䓞O~���P���W��7�>�_�����6,rG�w����ו`}�XX>�M���F`c�R��F$�zc4��K6:|�kt;Y3̗���c���[�v��9�n�#���m������I�@rܘ�m����Q�	Lq9���hm�@�{)�s�]��G:��qF1ȣ0���O{ڀm����=~T�崙 9}w��29�fF�6ܚy�M���hgrՇ���n�X��Nu��UTҗy�fh�� 9T��P�a`|��a�� Z�7Ϫ���EPU]�5M�%u�2L�e�� d��q�9��4n��+zS�I���v8�f�:�U���n�u�����SǷ*�N.�u=�X�-�2�0�M!���ۨ��m�+ �gn��W&O����p��ln��s���+���yź'Se3P�c�.�^�WZ̖m�Ȯ�'�n�E���ɬkKO]k��`u�0�l8��V�ŵ�8�~�v���sYu� )? � �$�}�'��5և]m,F���#��uv�D��=����데\|���P�<���g7j�+�'�� 䚀}{\��*ÆV���Kj&�� �h�e4a����w-_�P�5Ƽ�f�
T�:���@G7���#��rj �{�c�G2G�9��h���>��V��V�C���`s��m�B�G25TUQ`}��V�D=����V�ie4�|��$��q<X�G��m]!v���+v�s����i����݊1��WYn(�9f�s> ��8�ՠs�f@>�{��Uҕ�2DLn7���ܓ�s��M�� �V ��AF(@��>@��'97�6G ��着�¥?U�m�	�q����4[w4�٠w�ՠ�q�1"@c�I$#���"���o$�u"��
gX��4���nL��f���߭���Żj��fZ�Ӥ<FKdҙD��+g���#j�l���[��P������oZ�V��6G�,srh�h�n��n�^�4
��f'b�dP��e��:�R9 ��y%�W�6s�ul��!5-̍M*�V��$�{����%�l�y��"'"1���B.�mD�x6��D@�M!>�c��")���ۺ'���8��t���`�H�����(�B.2�������rA���0$@��V���kG��(����6��0CC�=���	�0�t8I�
��ȠQ���ބxG�04	�8��0�6����3�}C� *F	�U��`�(EZ�)�Oc�	�0�!�.ԷMzS�x�z� "p����@O)�a���j�z*>�0At���U�"�W�(H��*2
�2 �(�؀t�	��^j����I�3�s@�Z�n)���273@/m�;9��ά�VJ!$�7~Vy�I��n`�rh�ՠg���{��_{s@/m�˽M&���b�'ME��K��[c� ǯ=l�:n�GJ$�]���21�x���! �n7"�/r���2ՀffW�/�nN��)٤Ӫ9��̒f�{n�[l�/]�@��Z��	z!L�L�$�-��u35T�?{��@G�ZHEH�T���]u8�Ǎ�Ɯ��h��hO��훓�H�E�A��E�R E��i!j
��8 ۀ�a���1 ��[1`��X�J*k `HDȸ�Zk),�V�1��\��d"�֣e#�� ���a�h����
�9�w�ܓ�ød��Y�KB��.���e����/�77j��v��?gm=�#�$� <i�n4�Qrd.ݣ��=.۷Wc�]�ζ����N30��i hj!�c���_{s@/m��h�S@�Z�l����?8cn��gs*�$��2g��v��;V{�y�qp�nBH����mɠr�V�m�s@�m���f�e�p�F܄�i��@�-��;�w4�f���b識����Ȱ��I	&hȩ I&�;2K@88��}�ߨ��������?j��
�-����^ڐ���I}W�LƗ�

^6զs��?�[���ܐ�wI�Ʒe�N��s�{9ϝgV:�vx���J[��u�[H��;���ȯ<�'<]p�m��[�öy^ ���9���@���b�қ�����/,��L��+�:�-&��[�mҏ�˻,��4�ڬGH�&�K�]�x:ʾ�	�G9�MgH��g����w{��b�G&"<�G7w&9��'|�:7!iqg�&�Z���:\p�.�Z�x�����2��7k�����K@88��"���WT ��b�1�&�޻V��~�ٚfڰ;���3�W�6q��R9�h�����E�_ۚ-��ol�;�j�>�.T������h�*@9��KA����z��H������i��{f�޻V�nv�h��h��Cf�Dъ5:<V:�6;wI�6�^��Jv����g�z붰vV�8���F��&��{)�[��hw�s@-�hs���r�ˬ�ܓٿX�U��
.˫�V��V��a`q<�M[��ѹ��n� 8�T�$�Poa�[��h��ZW�M,m���4I5׎ZJ�R�EH	Ky.��254��U�����6��[�/��nڰ�ʰ<�GwM����P�Js�e)��ζ��{�����\���x�ٶ�Gj�zX5��d������{��nhv�� �٠s��hu�*I`Ǆae�mnm 8�T�$�P�� $�-_�D$�̗�*h�R�LН34���u�'��~�͇Ƙ���R#yAq¤r ʅM�Uh�QG��*���ݵ`ƞd�-��j]e������"����j ϯR,Q7!&6��H�s�s@�KС%�����o����rl��d���4cۣ���>svv+F2�ys���:�랺��ˁ��2��5�N^�z�F���"�#���1%8�ڰ��j�i���rf�[�4�{^�j�Z�>�r��DBl��;4Pӕ-�����̞������j�s�'�5#�cn-����>�n��'�{��&�CCH}@O��X�x��
 �_>׷rNy��mJ*A6���V��Z�<�=	O�ޮݝ�3��j���˨t�I��.���!���HHR.�9�l�`ѻB�q����ۀ'�q�D#j<pm9�yl�8��@GN*�U\��T�'��{ͼ�r�337Px�#� 8�T�3��z�B^J"d{[=N��:u3.e7T�j�Z�>�r՞�	�{�V2o��}�V�DD���9!�L�>��̫����Q	�,ߕ���;���rڙ�M�R��eX���Vk�śj�������!DR�anꪪ��b����+��cn�:�'=]9�ܵ!�S�k�$��Q��qal<Zܤ�M���l�%�퍞^�j�5��Q���&)�g�f��;[K.���VvwI�W�^�i�2�/"[h���x��k�҂�z��=Z'F�@L�]s�vt�gvc�[	[��6����p�������;{f�:nں�Q������/V�Y��˚4�@���k��ݓ&z6�A��^�� �!�e��]��ZQsն�����TM�z�mls�sr��{=-8��"��}U�ޞ�W��45�I��6��-����۹����}��ؑ��g�HxG��9���9}�� ��i��k�Z�_nhu�גcD#q1�6�h庀��-8��"� �չ�����$hcrh��Z��}�|/���[f��vcʜ�dy�d�b$K��mn��7)�v���\]���	�	�K��S6��CBF�qF�o�h�v�hw�s@>���ՠT[��IsF��߶o��_��6E��I���)�h"B�P�
��RB�M(\�J#��r{���Wn��a�*��Kj$�� ��4<r�ӊ�n*@K�\�zh]mf^Ff���u"���m�@�^�7�A�q����;wn*@�j�������)���\	��]��m��ԏ��:��ȼ�%,t�#+qI�5?(��H����1�����@vH��nb��R�-̭��!���3@�m��>]�z;��hw�s@;V+YX���&h/}�7$���n~>�8� "�T�G�D @B�W��tS�uٻ�޾����E$i�I��Rb��T��qR�EH=U�}}�=���_a&1�������hr*@rۘ�� 8�FY�mY}�`VC:�˯��8u�6'��v�u��vKi� �CdC��icmD���s��h�� $T��qR_��۬�/���@rۘ�p�R��H���>W����$��17��[��}��6�ݵ`q�l�vLX4�.QR��TLҰ�
�������{֮I��f���UX@W� a��Y�(K�:v�X�{��������r�i�"�-���EH774.�����P��!�ō��Y�[Mk�5�1����[;�d&�"���h�0�+wv쫽�@rۘ��T��qW���.Hw��� Y�l�T:��d�)���9ӹj����V7vՁ��roRM�3�����I�rf���nh�� ;m�@88��(�R̟ftf�U+C���Xy�6aܵa����@����E�#&&�7&h]�z�I,�7��wgJ��mX�D%
""?�����U�U�����EU�("���PEW� ���UX�E�E�@T �E�0DX�BdEU�DXDXEa@@�DXE@IE�@�"�("�������Uz���PEW�("�� ����U�U� ����U�PEW�PEW��(+$�k ����ȹk0
 ?��d��.�� }J�   �$� �    ����  @ @5�   >�z���HI�'m�D��٥T
R��%M�5$*�(��U*(��T!!   B$66̠F�*�    `�: ��(t��]G)JS�����)AGfSM�`���Bg��� ������7X�t�[�=�A�����  ��i����yԍ3x�@� �������u�s��{����p�� �>��)����ڀuC�v4ͷ�$��;bA����{�B��۹�ػ5w�<��к���w<*vӀ Fvz�x�JR=�l�#G{���t�6�U����M�^ͭ�n��W6.�]7��]��S�>���)��t �^g�T6_ ���=��A�]`4
��3ӣ��y�=��=7��h{xB��sk��p� C���k��th5������{�O&������}�Èwb�N]R� �Ġ�m����(
_ �g�5op���Dx\��{��pz}�pv�l��� s�:w`�^�=���x�[�H�Ǒ�r{� ����� ��I�;���Dm+���7a�g���ݻӠ�)����]� :\� .�i��g`:o���E��:i6h��:   ��
t1�4w�@{W�i����Jm� ғ��44�ܧM4p�w�0 �fz
iM��(�ܥ(S�q�M(  ��"�jRT� 4 ���R�j�a�2��U*Tx�H� fU%6ҩP  ��JJT @E�)"���6��?���������g�g���I$�9s'9.\��."���,��*���U?����� UW��*�EO�����BL"D�?�@�Tn$?���s H,�r2B�ZB(Ak2Zh��c �E�V`�&4�%�˔ɦL6M�r�E�19H��I�.�0q`S���"�J�9F�a��?4��Is�p��-l-$�������)+0bA#aC�$d��(T�WK�F�	!.�Cd�g�R@����Bg��!��2M�l!L9 �C3��K���!����$�����]��O�����
bI#';�D�	^Ad�7�l�^e�k-���7�e��Bϼ6�I�:2`&�3+�[��1
��hKH�xK/�A�#d�<�y-�_�����z�:_�뎸|���9L2���0J�9e6�$a�
nC&�8|K�2!�ٓ��D.\3��Ld��0.ˀ�Qdf�ѭdwv�d8�F�(u�� iH4B$��$
8�5L|��hq�4�w����0����6�f3�cL2`a��9��$bK����_Ƅ�q�Ͼ$���Ep���B��:$PÝJbW��0R���c�߃d�͛ј�$>FS��(g��c2��q]�o}aL�
�a_��H��0^|�\dc$5{󻤔�#�?Wt�.����+��Y���	>1�#D�*B�	d���xl�)�y D�#�t���(d�(|�`�_��h2jjٲ�4�LN��2i��dM1��e)g8&��@���t��r�%۬d%���{����I65%٪`	��Ip��1��$��H�XF葒P�9��v��"�T����ā��$$!L�I�Y ��0�fu
�u~�RB<yNH6Ɠ���7v����O�	B0	
[rc�	 ��l�$�K!$}rh��憤�q"r����>��XL��4���t�Ɵ�S9 h�z9;���s#k
0�zc:#S�$��c�L�������G39e>))�������Iߜ�e����8��B	X2�����#.��j:|�c� g���\�0c�8�Ĺ�5���]�S,��>.Xh���	F1���Ss5������k�?F���?kߓ?;'[����3�4���ă�s��L]T� �L��l��.��`��17��vˀ��ˊ���ɮ�CZ�Ӵ�B�T�cH]����
�(X`�Q��RaR,-�H�M��t}��d�`�� ƥ,
�i�YC$�1�F,@�����	�D�$I�`����C�hAa ,��4㔉h�	\$.5�c.>�z�h5��>�W1#-2��I[��`T�S?j�8(�,"A�I��؇����
B<x��B,Z�c"U��	M��bPē
f`Q�B�sBF�\2H�Rx�=��I��,�'y1�HB�B2GpS`F��#�*Zd�6Hi�*J��H�f����s7�;w!'y�YF�^��9Q�Ezh�d�H��p����,	I��D���e~S����7�F��89ӒP�HM}�2nH����B�tڑz�P�C��l�$6����4I*�𩐃	\l�>a�LA
���B�:h���Z�S�FɁ��H#��jqކ�C;p��٢f�$���F��,k΄�hF�M�B�a
��n��~!������ }���$��$)��:u ���;�m��\�fK�\98ߐ���$%��l��#bA�B7�*`3��1�R��"����Gƾ����ɚt�>��2U�!A
2vl��L`o=����bo�XS7�'�Ӓ9aC8�4}����5'�Y�72b�0�F$���!�#�6��΍��q�[`��w��#	rf�3i̧PW|5��J�!� W�-�"Ƙ`PvP���Lq��# A�FB��!$C�`��%�$bl�Rp$X���B�(dА�$����"[ad##i���*�Hp�p�F�3�dĸ&Nd~e�ҕ	Y���HS�8�;������0921�`X2��ѭ�{a
�����t�'�Hp���!0�C	b}+�2��B�B&3'���פ�a��!�k,�5��s�>'&d:���0���
`�e��	�:�j��/ƎI�w�29��G��p�ԉg�#�ð���HLD��p@���L���d�|��qu�;	���\��L����I�.Ct�$e'/je��%����$v~�0�fr9��$ �fۯ��	#�>9ϵ��4ۜ�}t�!����b
�pČd��C����x'l��n�zc�5�Me���C�Ϝ=��Y#lHtq�s]�XP�$�0A�M^ЏKn��y��I,�K4'^�����#�	���4Ft���X�E�R$0²�d��-1��.�RB�Rg[:�Ù���b��Y
���8'H�n2���m�Fr��S���!�������d�>d3~.�q�2�<�p\9d�ØB9!c#YL��C�_�
$)R#�3�����d�ʛ�����n���6A�9�B�V#SJ�¤�p�②H֒D��1�\d!�$�a ����@�Q��bA��a
!/t|fH��O��Ji�pf%�dJ�XT�kln�SO�@��d%pM�9�	�)	!�1�:�@��x�;�$�"HH���d�#�W�,�IyׁE%�e���C H��
B�q�?6h���Mh�P,+�HP�1�����VFD���WK���>g�
��~BL9��H`�evh��1�rjbM�1!���@��O�}H�.3M87��-q dtmń�.$t�
`!#HCC�2���8D$a��!L98��1���C�$#�kZ�\J!
�]�H��HD"F��,�'�l+	
�bc���9H�(��б���j%�!8$+�#��$>H���(a�!�%	 0Ja!$���)�C2I&��t�`��+dR��@)��t	IP�5!"Sk^%BJ�Y�&M
B�>n�B�,����뤔�G&��p\c[4�)��3�C	3Jt `�vHT�vL���Y�g�(r�J2���A'�'vha�D�W#�6s�H��	"P�*ka!F�ٮ����aLqg$3�'���x��Ń"B㬟
&���	n$΍w����u�w�B�1������$���&aI�����gR,����{>�x']��>��Bڝgư��t��9I�I���[��f�9�?h#�	��D,���*h���p1�a!�F�%��Ӳ$vK�Mbo@�
(a"ɦ$N"��"���0�Â���`2J	�Ȍ�T0�F�L�L��1(�`��B��dJ�V6P�&éՁR4>!T�L�����m�s��*���.�z&����e���R0Ϝ`"\b2aBE���q�d6E�H����b��K�X�5,Ri3���ڙ�M�h@�`�W	�4��5��^�h?@$l`${��@t�AbBHF+
0��2��S��C���d�I3�ă�"FYxK��4CX�w�kl���/!����<4�J�A� Lh� �W��@s�H�!��~6��̦�1D��C�{�Ғ��Z0�ss�vý�߱�~^�e�i�am׿�\	��+��2aֈM&��%&��+�S	#�|����L8qx}5�;u���P6`&%e�ٜ\K�4ξ��a��2�i�9�5�sﱗ1#-���1�����$܄���aL&C-�����	�d�eH�{Is����g�'��	��(���s\%q�J��%�f���/�u��X3�I���黭$�T�4l�I*b�`�	��vC�I��F����q� BX�"R��pHP�,���>����������`����_���p�Xu�s��te�@���tm���G�Ĳ\3��"P;bVp�S*ƤI�J,��(B�.��q)����
?"p!a`s�'���        �   ��� m�  �    [D�����  �                                   8�m� �`              m�>�   @   ���           [@     [@�d�*m�                         ���ku��Ջ�m����ક��#R)Z�o��	w��@"E�m�#�)�j)XBT�l�Qc]z���$��+Zh�<���pԪp���3�p�\l5�����m��Nʠ��  ���Ca�.�ջ e.���G��,��!ζ�6�CgR���
8+�)+R���x�	�pYz궍M��Am͒�,�6�`m�۶s ���jN�o   ֳ���i��u�{�&���g��mI#m��am[[l �a��`m&��e��N�dǕj^؉َ`7Q�)k8�[U� ���]ٶ�ba�`����F��)U[I����h^Z�ݭ�� UO[(��R�ت{n�yj�v$6�O�k�>�j[��+.�UA��qH\��������eUT���ک!
�=d�1:u�Ü�L�mŷ��r�Mn-K5ʭ��j�V`�sh���-U@�%���B�$m� Hm�f���ۖUYYyU�N���V�A�rIm� N�[�� [�r�mq����+m���E(Cm�Z�[m��[���&�6ٶm��JP�iKm�n�(z��� A!��  6ٶZu�u���l���*�U��Uږ
�j���`3m�K�h:�ņHI�V���J��h�"@H�L�VZ�W5T��Wfx+tAPAn��x�K�ڇ?}y���r��7���Zp�.ͦ��ˢ8��At�Q��h�i4W#�ەm5�j��R�t4�[p�m5�	��$�t�*�Z *��\MN�%�8i�j�j�9宽(t]%��lk�ִ�kq�յ m��i��-�c��b"�Y��C:z��j�R�]Tl�[m�`�����mU����a7R��m[ʡ�j�a���[��Nj���!�ѵM�H�[@i-ւ�"�UJ�9F�U�/���w���٨$ԁ��q�j��
CZ�k;.t˱�i'c>���^�!!"�Ҝ���"Ki�I.�U����t����,��e	qҤ��[oZ�B�$]&��d���=t���v�"�  �W8�[��j�����u(m�M��`۪�j�5�� m�M�`�m����!�ռ���UU�*�ԥ-k
�t��UG�����d����-�h6ۚԖ� �i� -��Z`�m�v�j/�А $V��ʕ���V�I�El*������~Uj� ��魕j�$i��yؐ)�Y@�Fy*�f����U@AH �u���H�h� Z�z^	�g/N�J8ݶm�d�r��M�ܒ6Ӧ������p �R�R�ԫ�X�W��	�7��AĪ�T���1b9@V��R%�� �U�Q]���&�
�E`�SJ����<�W�ʹ��\A�&4\���^^WR��T�&ʔ���^�ݙYa��Z����P�[��bc�l�vC�j��XY[hw*t[�f��K	,�݀ �-e�2Bki�7m9��
��2��gf��V�k´J�Г�m�-�0$�Bj�54� �մ ��l m~ϭ�|q�5� 6�����2`x��&�̀ -��m���� Hu)�R�  A�o][6Z  �$�����	M���� -� ��r�vksn�[J�O+�۪����&�.���ju�H��m�D�Im�� 	�H}�P
�+�Uu��̺���m#� � ���  UUU*�� F镗O�c�zPݶ�l.�tP     ���p[@���n��6*Rej^���7V�	$��  �4т�Tv�Z
�Ճ@���m�pqJ8#0,; �e	�m�]����]UR��Q�]R���lHp�ڷ[��6�UA�)-+4k�]�����H���R���$ɥҎ[��$�KA�] {E�V�S��T���HS��U#��檠 ��]R��Ü�M�oRE�m�+���(�.a0a��v�Jk� -66۶݃�ۢ�	l��e6ؓ�"[��(Ռb�h	m,FD�ڔ�-,�Og�w۫��w1�g���w8=�<F��N�+b��,�-б2=e�)#lm�P@Vm4U�'km5R@��ʯ;J��g\��l�҉�glXnTK�̵T�V��z��Xn�]�Z�T���9j����YzQ��T�m��Ć�%�@ �D��i�nץ�WR��:VU���mڔ��S���*�!���V�܈��%Ԡ� 6���j@�Y��	<&�z��$��-aJ8l.�[uǚDεOG4��I��sJK#�he�':���F�:���Ve�T	fiV� a�����OKf�9-�z�[e�*��IF�Sf(-�����]��9%F�p��=H�8�MsV6$)r��[yV�{Kb��Ԏ�탷Q�R`�������U4���-�* V55@V;�8
����$q�ʭ�s�j����.jR"iV�؃�!���UV��Z��3T��U����?YL���J�
�UUPJ\�u��:\,T��Z5�& *������ͥPبZ��2�#����Q��8n�+�e�i#m��l� 6��Y�mA"t�#h0H�f nV\֘إe�Ç`(�Z����-�����a�K����9tR����,�6�@&�w �wA�E*A���Ul�]C�`��5�Eq6ƭ��R	�Z�RX.�j�t�:UIjm&#	�k�۰�i�Y��J���pqձ�p�bLrԲKn��6� ��&t�2�J�t�Ԯ1Z���'J��M�!ʨmA�H�`�mV�H�Gh.�j��\�WPT�zm���'f��Ѷ�	m6�հ 	�޵  m�\� ��Ck���U嶀�j���W�h ְmz��ۃZ��m9�l kE6�Z@N�Mv�l;+UU[UU@/'fUB��m&��� 	$UUU+,�tĮ�UTL[�*�ʩ�kw�m%r����Z�AW�R�y�m��Us���~7�޺t�cQ:$�m�Q�UmU)Ӳ���A�[\H�Ys��Gd6Dk�����+[J�@9�	��W  6�m�M�ݰ	�d����$� ��h  m�[v��MoI���j��i6  ��$���I�h�lm&�C� l���&���Mj�m� ^����Z[%��l ��.[ L���P�~�}��U���~~�$�̲����UUJ�m�lUm��  ���  ͫ` ,;&��mmm�c^��v�n�6�8[J9�m51� 뫪U�kꯪ�(���T��    6�!��ڒ�8��Pٰ�X`O9����d��RY�KȞ��VXm� �A�ƞݝ �Ίy媫�L��vZ��6�kjӶ��l[BKh���z�M���> ��h �anV�a����l�Y�$`�m� � � 	6� m�  d  � �� m�[[l7GP9&ݵ�  �Ӕ���e�F�[C��mp -6m'�m +e�a�l	�P � )BAn�  kZB�鰶�_Z�	5�0��ld k� ,H ���h M� lh��M� �����Ul6ۀ� m�8��m �a�ѧ.@ �`6�*M��q��[Am	6��m�c7ge\�u�U)*��FZ��UU�v�`-��˲�UUJ���ʪX���UUV���z�m�/Bո7g�� i06ݚ^f�˻��o�� ��(<T�+�� �US�օkc��U@uMT�C���m�H�6��lE���V�Cmp�m 8�ݻ7�}m� -���ӆ�m�z��éY�m �
�ʢ�A�,-��d�kev\ڍ�V�U��O�6�?|_}�>�k�N�_ko�o��gX�#��k�m �F֤g4V�J	l6�[X�ԫU:%U&UA&��iVU�UV�ؖ��V�,sI�(� ��  ���`-�(n�ls��Hf�bT	f�6��BNڶ�ܠ�{l�H-6mn�@���j�d�0 � [A�����ڸ�\��4��2�h m� ڶ��l����h��U��v튪��8�IU]�V�@T9 60v�x :�Z5`�E�@����h���[r��������U�K̭! �J�Jh�P&�m�I'�h�)���[&m�`  ��  ���MUUU[$�� �a�@e��Yr�2򪽮��mT�mP�EL����A��Ї�o��� T���A�� m�&� �T�	�$�"�(�Q�E	Tv �M(qM
"�FWU7�!M*`:�C
�E:9�)�*QW*#�( ��d��uW���X
"Vb# ��F
�V# `^�i qb 	��`]#΀@ю :U��P�A`��v�~PS"�����i�% T�T����Ł L �R�@���/N(����2 ߪ�`~C"*d�h��
E,U"�P�U0�O���#�$HDl��mX���H(�t1�$�0������T�#M�9����G��0Dt =  #]`: �����0����Ev��.S��J4�&�x��X�EX� $HE�$d	�`!�:�GA���|�L�;C��a"P\�H�����c�EJ�Tp����T FYB����G�?	T�#^l�,`,b �H0�� 䊇"#���G�� ��@�";@ʉ���@@�H���q���*�@?�(q� "!,��|UOaF�"
Ȁ�`1� "�!(*�� �`���$���   ��d��Im  h�^��` H�۰    J$��^�%�	6ra�r���<�����n+�h(�qY�̘7�7��X.g��A���qj5�s��[�����\U�x�͔*Si�qq��c5��Ӥu;(��qv�MtN��6�N�d�-���ԍ�*��;����B�Ѫ�w6�cƲB�(+�Q�A5&v��\S�+�8���P`Ղ��V��'��P�9��1�s����Ż`��!b5c����{;�Ůy3��me������3Ö���S�<�N�.m;0��53�c�s�F�]��<t��hTg��6Ͳ���u��Q,ڃQle�.ƶA�{�-��i9Λj��U�ˆV��c�m�e��
,��^���cX�&�gv5MN4��Is
�mUK�m�c���ܾ�p 
��]�U�:G���5��]�6��ks)c4��n]�tODX��$��t.�[m��3u��]��O@�d=p��#�%v�;Z �V��Y�ܰ��P.�XQiqM�\�A9����zsvь1l��zs���n�ɴPf"Nݞ��+��-��;2��I �٫����;7j!�� �5��M6�б؍	������اTffnC	�
`��jm�L#]R�H�%�b�Х�,�R��g+�BL���1Rɗuf-�96$��K�)��Dj�y��%,HH��/[m����Y)��D����I��K���R�B.xԒƺ�vM���������|ܬ�mT��HY4)rҮ�J�0�V���Z����RZ��HU�d��HU \`bXe��`�[;dwg��I@O�/�S�C�/h�*l��"���l��y������N�mƴ��r����KÌt�Y��^��.w\�Z�������{C֫�tRv����&J]6���7e�Z�k����:I����w���V� �0�C
;=���/(�E�R��Kq�[����Ut۰�%]� ��iD���-�D�ƭ7d��:��\��V壢ܛ���]�t&��j�g���m��1�fV�6���1�.�x�z�rZN�x���l僧%��9��bõ�nU�xzc*mɛ�5���2f��g 5����-��W����̠X��GvP�	C��b8��$��w���I��3�IDh�5PU��RKl�)l%����ō	e!h�mo�>����j	�v�I�7�9��E&��d?� �1ı9�{zMı,K��G�Z��M�o'ND�ND����f�p��1������Kı9�{zMı,K���j%�bY����<�GL�f�F�w��Ȝ�����q��Kı9��zMı,K���j%�bX�w���n%�bX�!�MCm2�w'ND�ND��w��n%�bX���nQ,K����f�q,K���q��Kı9<�|��ԥ�w��Ȝ�Ȝ��nQ,K����f�q,K���q��Kı9��zMı,K�=���RQ���L�^�K�@�i�5K�˶�l)��Y�B%b�;`j�5K��)��%�bs�צ�q,K��w��j%�bX��{�&�X�%�~��N��Ȝ���'��&��\і���n%�bX7��MB9�R����`A�ػwq,N��vi7ı,�wMD�,Kw����r'"r''��Wɀ"뒮�s���X�%����f�q,K���q��KD�Ns�٤�Kİ_��w'ND�ND��<�{�U��\8�f�q,K��s��j%�bX�}���n%�bX7�wMD�,Kw^��r'"r'#���_�����q��Kı>��٤�Kİo��2��bX�'�w]�Mı,K���)��%�bx��.��g8��!�۲��ڮ����Ⱦ�tn�;j=�=g<s�A�EN�F�e2��t����ND�I��}���X�%����f�q,K��s��j%�bX��;�I��%�b}8�7�\cM���:r'"r''￻��n%�bX7�wMD�,K}�vi7ı,�;���x1S,O�@R|��֥�㼟D�ND�y�e5ı,M��٤�K��H�H>2b&`�s��j%�bX��5٤�Kİ{ηX��d0c$�0I�gMD�,K}�vi7ı,�;���X�%��s]�Mı,bN?yw'ND�ND�x�y��������ri7ı,�;���X�%��s]�Mı,K���)��%�bo���&�X�%���̳�nc��.-&�Kn��%؅8�u�,I����/�J�6Ve��y�E�Үl�|9��bw�צ�q,K��s��j%�bX��{�I��%�b_��榢X�Ȝ�~����J��\;c��D�bX7�wMD�,Kw�4��bX�%���jj%�bX�s���n%�gMzoﲅ4�l6ʱzyzk�D�7��f�q,KĿs�MD�,K��4��bX����SQ,K9����y���B�4��N�|9��b_��榢X�%��9��&�X�%�~�q��K�ʾO��H|����8Ϻi7ı,ON��i���<�9�9�����i7ı,�;���X�%��w�4��bX�'ܹ쩨�%�b{;~�0Bfۈ83V�#�':%bcf�4n��vV�4�Nl� ���n�2�j&36�D�,K��SQ,K��;ݚMı,K�\�P���LD�,Nw���n%�bX>�5��fC2L�I1��)��%�bo���&�X�%��.{*j%�bX�s���n%�bY\]�)�r��[%��4��l�s�&�X�%��\�T�Kı>�5٤�Kİo��2��bX�&���Mı,K��;�S$��Ĺ,͙�eMD�,�W9���I��%�`�{��j%�bX�|�s��Kı9˞ʚ�bX�'�N��2b�ݮ-�w��Ȝ�ȓ��<���"r"Xy�>｝'�,K��n}*j%�bX�s�٤�Kı0�CH��a��U�D#a*"�� �
�p��)��>�x�VˀGcbݲ��X:��P���.']'&y� *�q��7A�31��胅��sg\0nle��1q�kz��۰�3��ۭ�&Ln�;H�<���=��9[V��y�ף�K �sq�vVf�3X�����크����;7��]��ў;BBݱ� �w#�˝v�ݮ6(�v���j��1+79;9Z᭻�AB&�ˍ2f�q��P�MalIJ�lgJ��KȷMvu�%!�GB^�R�q,p���(SF�zň���������p�7veo*��	vG�uwj]�+� �����͸g�s�Oe`o���%�M���9h����ӳ �ٕ�j� >�^ٷ��m �̡[.�N��`�#����vm���R���`n�F;�:wE�SN� >�/ ��� �����K�=�}��W�M5IIm,����1�D8����n9Qv@n�V8�U��s��:��#����/��ٕ�l��I/ ��5R��lV��iـn�����,��"C�Xd� 4�\&-�r�ٓ�{YԒw�{:�}�\2뜤��
U�I7v�m�`{%��K�;�p�7�2�lMT�1;�Wv���{�\���� �/�;�+ >�/ �ݨ�����v���0Vr���t{�^v<����#t�K�RX�(AK]NN;E�ۉ�K��K�t���tGn�Y�G�HTy7U]�iـN����K�"�ǀwv�}]�@"s(V˱�WwX��y��W<�y�%��'ve`�)wN;���N� �{�ۆ�\��(�T8����xRI߽��I>���r��i�������� �ٕ�vK�"�ǀuw�eJ
-��"�n�wfV }�/ ����� �{���3V�X@+΁Z0��"0k��&�������#���D��K�΋٢�ݶt���� ����� �ٕ�TN�R�i;�Wv���wc��T�����=��X����l�;@��)���v��}=��N���엀Eݏ �v��q�����\�;�����u$���Ƥ�Ea�^������>�Ԡ9�+e�髻� ��x��y��{+ �ٕ��ll�\-����h��Sq��D*P��/[m��mc��Z�U�Yj%�&��%�C2��t����fV;�+ 7�^ v(K���I�I��ݼ�fV{�T�=��X;�^:�,��䠢���5wX�̬ ��x�ذ�p�'M�RYWI&ۻ��u�|�c�'^ŀ}�p�'ve`��jSM'|*����b�>ݸ`�2���x��6O��4�} -��I,�ΛlX5[6Sv��*AUS9θ��[�8	ʑ�u.SJ�V84n-HM1�Ђԉ�8z.��v�Q�Uֺ�ju�8��v�ʂu��L�"M5�P�32��M4ya���m�&c���t���U��x�l;f7F��v�f�y%k/d�<�2y�W���eL����qIͱ���b�{rę䚋�m2��i�iqF��$��N���.HJ%�V��KB���)@ƥ�Fh�h:m*�*X����U��wb:��cmɮ��nց7�wfV�ݏ �{7hQQ���,������'ve`.�xf�0���(NJ�lt�����ǀvm���*��v_�o���w�)�v���Cwxf�0�`�2��%�b�v��m�n�۳ �ˆꩾ����z�͸`�`�-���Eeմ1:.zV�=#Jt��R���>� �\�&�t��H�/]����ݘ�L� ���n��NI��{�:����G�E�vŷV wv^>W;��\ۆ�e� �ɕ����jP髲�wcwxf�0�\0�Xݒ�����N��]�����.�L� ��xf�0������,������7�e`T��}��9���RM��ԓ�#}�z>�ic��A�dp�إ�ܜ�����j�csY � ļ�Å ��ɩev���z�͸`�p�7�e`��F;�tZ����p�Us�H���M����%窹��A�^=v�v	�M�n�ـl���7�eaڕUϹ�Y��d�:T �A����A��$0b*�B��"K�h&M! �1�L$+��0�8� ��$C ���ȱ:!�0*2��n`4�L���+�;7R)� �G��� f�� 5,���r���ǋ���ؾ��W����:$09 ��2��L } pb�چOAƐ���8!�f�JE$�Y[�Bh�@"� 1 M��N�����G$*T2�.q�	������~��c$dV	`�QL�5J�~
���z�Q��Qv�4U� G��v
G:�S��p.�W�*u���{�;����y�zhA�lllo�%��$&2b˜c9�Ѓ� � � � ����;�����}��A�llly���B��`�`����=����wv~?K.̶���s���&�������t �666<�u�pA�A�A�A��צ��������i�lll/N��~�M$�7mZ�X�ɗ��;8�ct�6
��6�������]�3��]�F��v7w�ʪH����0��Wg���M������)l��:�h�w��̒�%!��0��ـvz�g����O߲����=�׀o�_o�>~�k����4�A�+X�
�-��~��`���;�p�>�p�>� jU�.�;�� ������Ԙ?rq�IB�����8��c����W�v�)���0ww�wv�J�`l�X���D��V��ׅ��f���R�Q�N�5��ѓ���u�V�v,�㓭��vT�I���.�&V wv^�ۆ v��� 	�)�-��0�L�?U$l��d��|�����R�z�!}WĨ��ݦ�d�竉%��>�g���v{���ȡ����,��%طn��rO�g�������ʮ%��e`���9\��=�����ta,vgc�󓓏�w���}�{G��'{�gRmF�צ��(��`%"���Â�0wBK�N�wIz�����]�����]��j�Cq`n�5�-��������Pm�"`�R k�``f��*mM��=4̹bn��me���׷E�Ȯ�騣�'f#��#3�cU�)��s�s4P2a�a��n�W\\l�(�9`.x3�am�HE2<�o>0tX�K%"C:��5a`K�� �u�#x����(��b�ܓ�ۀb)pL�ٹ'��>G�#��&s��Y��:l˭T��E!eЄB�&�׊�.�\�6�kYy(c��l������U.���ՀO_�ʯ�l���s���y`G�Sk�C��j���z���׀l���ϐw��XUR����d^�j�0`�T���z��6K�w��^��g����%$�����nӺm�m�wn��G|��v{�X�����0�um@����ݻ��}�e`��)'��6K�}� ��%�l����*hy�(��{oZs�nx�>�Y���o<n�6��W�(��ݦ� �z���0��~�rrs����t���E�Wb�[� ���/��z�Fr���s0�;��'}2�we�T���,N�QN���ݬ�~��>�2��D�׀ls� �� Ŝv�2��7v��L� ��xu�X�Ȱ���)�*�av�;�� ��xwn�Ȱ�L� ����\�k-Ҧ��+��@��ta������x^�1��yp�At�.0ݣ�;��;�"�>�E�w�e`���!�ݫ��1�j�N��r,��+ 7v^޹ v��� ��
��ݻ��w�e`���rW%g*�����Հwe� ���$���I��m�`v�%�/ �r,��XݙX:���Ʈ�R��n� �r,��XݙX���r���g������e�� ���QZB�&��1m�6֏�>a�h㈚=p4�;Tqһ�n��w��X�2�we�=� ��*4��Ӧ]��&��&̬�R@�e�6�}� �좊mN1+������ݗ�lۆ�r,f̬��V5e��'tZ���	6�}� �fV���W9^I����m�~߾���hɁ�Z}� �T�>��>ݗ�o\� �9��}�>�ᨻ3���hAB�`�e�k�M;C�5�[hB��bk�eeqm6`��ݯ��Oe`���7�E�}� ��Z$�QM+i�ݦ�� n�x�Ȱ�"�;6e`҅(��ݺUeڻ�z�Xc�a�es��w?{�V w߿^��0�]�\t���n��ž�y`�� ݒ�=\�)��,��W�Y�i�.��wk �ٕ�{�R{���=�'��{u$��H�,�$�r$��_%���,��nR�v��7a�����>�Ţvƹ"���0jз/C;n�솻��;';�	u�j�-�{����Rm�)���qq"]cu�N��v�i�X8��v�Zz�)v� 6��tZv��F�9Q)�Чa�&�\9�:�y���痋vyg�����8�@^�k��r�q��'Hc�;'$���e��B�=P��6�wm6�=��'O��q������Auf��C)q]��Ύ����X�kF�u[�oZa{�xW�aM���-�.������"�&��+���~����X���cV[mRwE�i'o ޹#�`�2���=ăHO[�v6ڦ�v�y�� �ٕ��//{� ���Q� i6�w�v����~����~����"��y�K�������W{	W[M�m� �H�T����{��Xf̬ ��~�lf�k؉(��<K�Sb���.H3J
-Ґ!��sۢ������l&a��a�5�� �Ȱ͙XRG�oeL,N����v��`9J����5U\�Cb�
�5	 jR����s�hԓ��{�s�wǿ�$S���-�6&�h�k�>��e`I�r,)#�%wh����BWe�e�����"�"�<Ur��{��6J^�,vڤ�T����r,��u������ݗ�}���٣����]��J��eX"�Z�C�2���V���%D�ط��:N����@4
jĝ���� �ٕ��/ ޹ v��� �mue�wo �ٕ���9\�$O^5�� �I�v�I\��J�;v��� ��x�Ȱ��r�,p�m�{�I;�{�RIߤ�F�i�:,v��s��.��0����L� ��x�C�ݺ|�Wav�ـ|�� �d��ݗ�wv�}��H�ԯm�ٸ�A3�ʒ+�6l �AⲖ���Y�\v���u�<j��;��}�e`���;�p�>RG�mM����	]����� ��y��W;�p�:�#�>�2��ҕ�'mRwB�H���"�>RG�vl��ݗ�)-ۻJ�7M]���:�XI�y��N�Τ�	t��` �r����X(&׀M��ʻ�v�͙X�UR7e��"�'\� �ۘ��|�#�����.X�iV-psGD���`�]ݗ�M�;h���n�	t·|�=x�Ȱ	�"����V��@������wx�Ȱ	�"�;6e`ݗ�od1X�����v��`�E�vl��s�ą�/ ޹����k6lM��۳������|�������"��+��.�{� �l�����B�jӵwu��/ �&߼����5$���I2|"|F0�!6�1��0XB!!$#B��aBB+ HrR�7�H^��HH,XE��JM7a�Ō0�0��a�2�z�C�v\pC��ŐX�ہC!���	R�J�!	$��H�Bx�G��B$`�0�2|�!��	"KX m*d@�V!��cl"E�aC<0��d"�`�c�mdHuѤ��)�Bґ�&C�;�[^̽L�B�c��|LĲ@�IA	 ����l�$+U�m��$�"��t.����"�t X�#T`�0�|�a��HDv����@�"�Y�)�#!Lh21�X��/�2j�9���t���$۠��# �C�2B�U������'I�~}��3� �89m���    ��z� ���  ��lkՍ�  �wm�    %,�K�k:�v��FV:�B�d A�5B���IE`���[�-�Y��R��i��r���Ù��ûF���0�8��ck@�M�H$sC4
F�Z���;[-P����}�̒��.�㣂����[��NL�E�V��v�٭q88���nl����H踕X��E��w��uPn�N����<������l�u�s�JQ��ܓ;[�鋉.c��i�A��/mÎ��
#��	�.CÓ�ct4��ʫNv�L�鵸�X;<�n�1.ʶrg6����Y���0�Q�̩x��t�>ōɵDY�K��n�K��m [�M�����F�@!k!�N �2�i6Gi.�ŵ�b^�l��-ە�V�5��X�d�d�2.ɹ�9'L'`� �2����q�2-�v�aF�Vx
�NnV���(�6"�j����IM�A��1*@v�X���<=Kt�]F�{f^P��.��G,�6�����F������0.hF �vͷG�6�N����n܈��HXQ\����]�#7ZT�1$�;(�Z�ʎ�]F�p;m�˗v���ր��.ˢ��+a�]R*$ۗ(���I��,���M�ɸR�'n�l$�1���:�N�Ocnv���gX���Wm$fMJ�݂
�ѥ��T Eյ�y%���6����Mc�x	V683��ּTnK�X�ز�@�Q�7"�K��+i�8�[eEh�����z~~�����B�JD�[uJ�r�H
fW�m\�<�P���m%өd��5�j��S�KG٫����n��)�+�nwf�"��b�?[p�Ѻ��J���]�qg�^w3�
�C�y��g�&\��M��키���Ɓ��t��^wNt�UWj���j�7��\vn�q�\��$�'	R�Jf�ff��rJv�G�Qj�Ы�CB$W��~Dh	�E��N����C�ڦʷ�R�QZ�ыg4*�:m���5�L�P��re�v�8Wb�rZ�� u]�7p���m��4ZY��N�;�u��=]��8�Y�a53 ]
����R(ƺ1@����$�/+��!���5xi��C�ݢ�I� �����2��\�4�GM�*��R]G.�&��zt�P�O��	��;��io<r��@;	m�;y�\�����t��+4�/1״��M-#E�)[�8 [��nS\�Ґ�3����	���n�;��w\��>RG�vl��ݗ�-����-�Mݦ���<�r�#�fV���r, �e@�h�|�����2�����\�q)��XT���w��pV�Eݦ��ջ�r,�<�fV#Z
����S�o ޹��WZ���2�������0e�E�wrHfJ'c�x����OGR�܉����Gg��VZ�]ۧUt��m��>[#�;6e`�ذ�`�E�R�]�J���9�5$���d p�@X��P7 1��
E�e�/�_���ﱨ��`-����r����Em{��nէj�� �s� ޹�q.����2���f���bv�RG�|�c�6I���.ɞ0������V�Wi[��|�c�6I��n��H���L���Li�]*VYջ�׶.�K�1cFx[vsY5�2����E�Ui]��6I��w^ŀj�ܪ��J�u���<���Wክ6�v6�ױg�$E���:��<�fV~��#|��!xcutYe�X[�<����<�W����I=�{�ԓ}�gŻhɣp��?��9$~�}����V��,��#�;6�jiҵuwI[��w�u`w���Vdx�lx]�ZTn�9t�&����ۻ8۞d��i�i��Ѷ�	.��hb�H� �7,jݦ���]��]��)���2��j3
M�wB@	��5vG�|�ǀvl��5wc���۴�V�Wi;��|�ǀvl��j�!we��#��wj $�E�J�n�>�tjI9�;�I;y��RlS�6@�*�, T)P! X��1���ڕ��s�N}~��o@�=��
1֋�[� ;ݗ�~�9<���� ��+ ���5��@q��]jB�ƕ���j�d:H�H���G�u6���f����M��֭t0�;���{ߞ�;&V�W�ݗ�M�b���Ҫ�Wt
���UU$z{�X�=x[#�;�E�t�v�!�wI7o �&V }�/ �dx�v<V�U�N:jݦ�wu�n��"��ݏ �&V��FaHe���h)'w�E�<ܮs��mO?�������xA\��9\�#r�;EV����M#p��$`�֤�V�1睼�jxUM�ƶ�H��9��K�=q<ƺ�n�l�d�aN��T1lj�֛����#Eݎ.W��
z��I]�#��6��c�ݺ�ƽ2K��K�H��������(ݠ8��=���S�ݪe�9�@8ͣ/��l�3gc�\��N4ⶴN�7D�W
��mXk�Vl�����|�����lI[���l�n��9�&FK̮xx�2lm�u�V�8�!ōg���u�e"˫����=���&ɕ�|�G�yOy�xo�� i+I�+�x�2��#��� ���;�p�ܤ���B�T���ڴ�	��X[#��U�n9~0O{+ &ğM&��j˻X�^s�x�_�l�X��X݆+I��*��w@���M�`��s����k������}��g�c��)H�A��(��Fؑ��8�YW�b�wF�s�-�v����<f�t�v`d��>�"�"���^̬V�[D�۵m�wX��x��"! �H��B ����x۳+ �&V{�\�+����)�i]6�I]�y�� ����6I��l��uAIn��"��m[v`~['��{���>[#���~~����_�Ai[C�VZ���L��+��~��	=~0�̬�]�F�M�Ycmվ�ɞ΁DE��pɛ[���l�%죣]"���%��If�4�Įէu�5{��nˆ�ٕ�s��{+ =<���y4���T�����ܪ��s������O߿e`��y��$�����:�Ú;B��';�hԓ���5(�b �К�Ur�G��z��_���,�������Wu���r����Հ�������'�9'/����tg��M_��ַwX��x����x�	��X�X���-��6�[G$�[�'9��2Vn��Ls��ۀ,fs�&�������]6��]��\0	ݙX�^�>A�� ��{�����ݫtӳ �ٕ��D��V�� � ���� -$�wJ�Wu�nɕ�Eݏ �wfV���T�ݤ�էu���ﱩ'=�hԓ�s�5&���$6!�� ~�}��M��/n.1j�iڻxd�X�̬vL�.��$���I�}�ذ�Gd5�P+m�����uE� 8Z6Ύ�ۜ���K�]/V�Ktr�]�Vۺ�l�V�&Vv<�L��Y-'Wi�]�!���&Vv<�L�wfV��V�E:v���wu�Eݏ �=T��{+ ����>��+U�4��TP���.�̬vL�.�xT�j��$�;�n�v`�2��2�	�lxd�`�\�9U�r%[BBr���������rƁq�A��n,��m[iΓ�=���.���p�G�1�$�˔u�[n����d��j�mi� '-�z���v��N�rn�r	�ZMQ�J���cG�;J��@���`�2��uf �{j���jࣩ#pt�"��&�ޓ��b�^p��n�:�Y�k/\���*�9,��3�F(����I��ˡ�(o$��ϝ�����ƴ�Yt"��`C�YHɄf^Yx�vX�%�(G B]���T�;��>���΁��lxd�|�����6��רI��I]�N� ޳c�RF��� 鱗��;;�I=�ռl}kk�f������`�2�����V�<�	��0�;tr���/l�ՀI�e`��yo���~���m������q�#5�vL��K�S���{+ �ٕ�rq�x��Xˣisv�@��.s/LTu�P��ݽ;r�gnա,�i�/0m��[��n� ������N���ʮ|�O{+ �^f�����j�Uwx{��kK�T��"!(J���Er �T-E!
�1�1 1�R�H""`TdE)��_*~ rk[ލ�����}���U\�$j�g�]ۤ�3�˜�ɩ'��hԓ��tj~ �o��� ��~��
��-�i[M]V�� ݓ+ �����2�=U�W*��{��6��רI��-�wX]�� �9U�V�����=��nɕ�:��12��f������(�/�B�����a!��y�
G*��t|Z�_1�=Z�U������N���7d��UU\��UT�C��{�z�����%��t]mӠN���7d��	��xd�Y�Uq#��E��6]�L-�!��'������2�S�W_uG�X�6	�*�0�	`&2E�p�$"�PI�-L!bB�L!oP�P� �Q�K�a$`�\��f���,1e�?E2�
�(:p%L4��,a&B2."�"A��0�f�R�H�#(UCbl(! ��|+����r�h`E %B�B�k��3�I�H��dL�Z�ÅF""�v|�~E
	�>mDب� ��T�P�v :t�| �YN*9����h��ڽQ<�o=�hԓ���jIÜ��T��;m����K�S׀o�~0	ݙX�X�Tf�����h(Uwxd�`�{g�������"�lx���I�m4fZ�].,,k4`A�ٱ��رm�#���Kz��y�w�P�m�m��@�=�+ ݓ+ ������WXO߯��<��i[M]b��vL�.�ǀvI��N���W)#k|!]yn��cWu�ymO<�L�?UUW�o������+ 7`���m_��x[�g��=��nɕ�9U�4�[��������C�Jۻ0	ݙX����}_�<��`��ʞ��Ԏ��<dM�5i(��3����[���^9�K�ъ��im	��������!j4�w]{��.�ǀwe�ܮs���T��׹n�N��n��[ݗwfVݓ+=��)#��{��j�4 ����y`�2��9Uħ���-��uv&ڔ�h�v+m;����r����{�k ��~��"�lxǱ`}]�� ���]��f�~Q�������}$��{�ԓ�s�5$ʨq1A�,��D����g�ǌc-�kv�~`��v�bc���Yzج��]��■;$m[[ay���IBg��Q-cc����c�����y����\C��uֺ�H	r]�U,,.��FPt�Q�ݨzj�V�Y9��.�-fș'lJ���Kmf59�QrX����)�M����m���k*[�l�/;T�D�,� ����1�-�7p�n�KuMxc��a��t��w?�?����o���[5�y"��f�F��Z��W:�(Ɠ;G�������Ӿ��"�����^� ��,wfV�fV n��4ھ;Uv��b�Us�ďl�V==��E�����Uq"J��-��;��n����6l����9T�����'���>��\�M�i�wHwu�lٕ�E����b��W9K�=�`�}��y�V�nӠx�����*�=3��{g���2�]:rF�@C��tonc\�����f-�U�m�GJC��+��8J���Ѩ6�>*���ر$��ϫ�Ke�G��Wɤ�����$��ɶ�HX;���1$��ϫ�0��b3$�H)U
�V�Q���p�|�y����)bI/�W�?�I-�1�IW��MNV黢�Wu��%#�KIG����z���z��Ē^�{�����"�HT��9�n�U��d�o{�z��ާUV�r�S���Ա$�݂t�!��ӵWo�JK��I%;'���$I2�IG����Ilv�-��.�Nꓰk/F՜��p/���<�u\3cZP0�m@�J���.�w�K�9��nO��������T�e^$��kc�+��I{��F$��zQ�Κ,����w_|�D�*�$�{[�$��1�JvO��\�mz��
U�9v6��[��U}�O=�>*����Ӓ*��ڐh��"���_(}�{��_|�D�ʼI%;(�$]�퉠Wo�JK��I%;'���$I2�^�+�o�*y��Ibm��X;��sf�����f�m�K�{y����tﱿ��y|�z��>�<��έvitVZ���C#.0+YLĲ���Z�YB��]� �Yn�ƺ|�����U_/���m��;��_� ���w��ݶ��D��F[tɴu����?y~|�NNJ������	��}_|�JI�bI-�P:"�v�j���$��e,I%;&��������[m�:w�����L�2�d��G���rI�}��gϋm����[m�8s����(�"��w|�U_����|*cYCmm>|RR\�bI/Ur��\��ޤ�����$���'ϊ��Y��[-&�	\q�M���q[���Bd��]�)*ܼxClP'�NFv���{�b79[����y���W�<݇U%;'����I{��F$����|�˺�4 ����II/(��UT�K��}_|�^���$������U��[-��SE@�Vڻ�1$������$���ĒQ�l�>*����ϓ�� k.�����$�U��g�F$��<��$���bK�K~��gϊ�O0��ŕ��\���m��wݶ�P����v�~���{���=՚�ۀZ���V���'�"R�C ��LD
D�� �h�����N�����clnʵUWO[%b7hr�g�7&�)D�e��f�X$�;R`P��c�`j�jkj�#����nxι�"�=e�&������l�nB�.�U�jM��eK�"=����al΁�.�xu��z�H;�t^6mH[Y��g�,3K�İ����(6eǊ"��=�u!p4�[H�F\�$s�:G����v���g�xrm����u�Nt�J����k.!^[��s*�0�aH��&��̚?-���t�X^��G�{él�iګ���K��הbI/��W�$��1U_�����_/��L魡2l��V�w��f�������ڳV�}����Ԥ��g��K��X߆�-���]�}�I{��F$�׵���I)&Y�$�d��������2w����nN��_�����^��έ����f�m����?�o��j�����14n�Pm~|U<�����䒒�#IG����I~�q=���bJ�9���&�K5�v�M��W����d�����Yc`��)�Ǚ��3�v����ݻ�I/����JK��I%����S����eG����<g����2�&�m��{�5�b�`�,�r���X�wY�����$����}���|�L���-�&����W��y���I
H�IN����$���Ē[�YAa�m��f�m{�_ym��v���=�_|�R9��%�q�^����%�+�Zv�$�r�]�����|�>*�rNs�{���$��������$��UR�eZ�Kr���T]4p�������� ���k!�Yۖ1���;�^�k�e��>�U���F$������I
H�IN����$�HV9n���I;F$�������M�/{��$��{��䒒�#=T�K�=B�&��j ͯϊ����WϿ��7��_��H����ֻ��Vj�|���_�_���`XmCL�뺒�+��g�_|�^~�3IG����%��\�����Y�~'��˰l;O��rc1$��s����ޤ���;ĒS������y�7�[G�1`�$���\)��j��|�?��,����є���Ӝ坙{@�]�u��U��O�ϊ��]�Vwg���%��I%� ���)7I�^��m������:w]�}�|��߿_�F$������IG�0�t���E�Iۻw�$�����%%�F%�Ur��~{<����>���U~O?N�.���8��D���5m����c{��{��:��U$ � ��t��~η~|U�<�8��&�����W��~�7�m��Lg������c�����{����U���Ȗ�-ΣG$�[����͚�cv�qt��]6]YaKeґÁ�,��v������$)#�I%v?�V��=՞DE�1m�8w������=�.�f��u|�m��}>|�;�N��*�~�،I%������$)#����J�Z)� 6,��պ����ާU_�o�����*���)<�IG����%*U�l<HZ��nN��99-��������}��$��#��ꪪ�?{=�1$���Y@��&�;C�V��$�r'�$�͘���uf����۽�o ���m��a�62���P����!��\�)	��s��0�H!0���D�G��O��>��r�5��޶�V�)Se�a,�s�;�r@�&�D60х	VS�at�P�];rA*B�M��r�����7B8�3!M��v��Ğ�������a� �N�!�   ��d ܄�h  -�4�:Fհ pF�H     [E��&:Vssv�I*��ka1t�� v��������z(�y%k�F*2�t���/Y=p�X�N���8������1�� ���Gb�v�V��\�Tj"Z+eI��Ԋ�0�0	� h4'G�M�3�����l��8�-��4t�+ݙ��v1�b�B)�:m����%W�e�Ir=�.O'�]�K�'�XN"`�ژԂ@��` ��e6��&\���ͧWC�Z���
�@,�͖�5�J�,��p,�R��O=]"�ƓX��m�B�{L�n�]I��Ɯd-,x�5� �&�Η���<B�ln1##{d�N�����XP#Y}�cH�Q��ك1Ó"[ `��m���2���h�-�'fl��9t	mm<�=�V���`�cDT-F��5��i�w3�@��Z��X�����읖�<����	��5��v.\6�܊�h�n="[��+��`�օ-�T�km�b����b�vt[�XHd�c0��&�3��g�ͫ��ƶ!�n�� �D�҉��F�9�-Α7k���!�v�f�e�l�p8�J������]P$
!��F�j�b݉����V"T��m<Wz1��g��xb�ۀz�놔�ݒ�0\����t���Su��dy6�Jt���[<���˶ۖ�I[i� HUH7�Em�[Gm�Cƶ�l�ʽ�(L�S�g��r�F� ]6 B��{j�]a���&޸+q��=���g�6���)��������I�1�ʲ��ڜ���#;!RrY@y��k��^^�D�˰v�r�A����7	�(K�noF��y�8ڕ����Y�ZL3N���÷ fQ�*Ff��j4�Z�`��49�%��j��vG�4d��j2���X���UT��:v7�]��3n��f1N���k�
�]T�j�Ne쎻O�������C�Tz::p\
���]"
uT4�~�?S�����&*��;M��j�Cq�mc\	/K�y�d(�-DQ&��1Vƶ[�y�lt]�ΜPX] �t�9�6�u�ڵ��.�XV[mT�	�m�LBdPSr���D���u���0b R��K�a����b�]�+2�w:%(�6����4"�]]\8nqnj7;���Ί�vsX�n�6��]�����nj�)n\����54G@��9$줝|lbK�qR�{2�L2��q���U%���)T��A���nq����I�ލ�)2`��ڀj���	�b�6=��\�|����z�*��[t��I��&�� ����'\� �6<�9T��8�ʷHNդ��y���'\� �6<kذ	�@ta˺.؆4�Z��UR�߼��<�	�b��U)��z'���t][i��5M� ��,cڋ �r,H!F���*�\-�۱�B�Na\u��4&�Bc^�d�G�V[�m��{:^�ص�u����|���`�E�j�<��b���������n���9�u�M�q���Go>XW��M{~H�xW@��6�v�nŀ{_��RG��K��,y� �jTN�7H�E�����W~���s� ���qM�y`�z����[�-�BN���,�U=s��	��X�#�5V�)*U|UhU	�C�	���fy׬T�v��1�]��Ŏd���#ٵ,�
nü��}?�݀o\� �6?r�A�s� ����×t]�4'V��`�ǀv=� ��?y{�}x���hi�n{$��}�I>�9۩��S$ E	(A$0@'�W �����N�� ޽��
��jU�V��t[i���W�q���� ��{��7�E�Eݏ �v���8U�uv[I��"�lx�ʛ~��-�xcذ�PIeZ�8�#t:F.��E�x�ᅤ&����!��b�5��Ja�a��nfנ|�|��"�ǀw^�������	+�݃|E��ڻ��}Ş�RF�<�������ں��`[����Wv��ذ��x~��7��,���� ݭ⁌��7uuv��X[R<�s�RN�w�ԟ�B�R@��)qT\�)��(| �$����=�z����aӛCj5 fנ}�E�E�<��,-�����zO=��3E�.�XVh��j�^��1�K6�bT�SP�Qhp����zǴbhji�k�~^���ױ`mH��Ȱ�kG*����WE�wo ?s����q���~�����`l� �v����������`mH��Ȱ�s�ļ����y`�
��awE��Wo �\� �dxu�X��8���� $�W����"�am]��:�G�w^ŀ����ȰU]�_���.ߢ{��P����ñ�U[q��Tdv.�yg�Йa�����AX+��͗R����^5�&LM&��{k"�jѯ��nm�ڍ�C<�A��s�`{b�g������O[l:��l�j���s�1"�,ɍ�<�V53p�ao[c�H۞|�]��z�gOb�k��RѺ�&�Ivؚ��seQ�G���찃����-��]>�>���g�Ns�|����r���۲��V��C�[v$�VV�oڑ|0��N�<��s�NӴ���wo�{\����^��ꮟ���?ſw��[}�����-h�� v�K��UĎ��,T���{��?I:H����K Cy
vh�Zo��� �<;UIjج�Ix˦��q>:�,=\�W\���y`t���Ȱ�ڍJ�J�����w^ŀz��U-�����uI�������}|�&U�=�[�w:���S��g�]�GM�9�6:m�C�p��*�);_ l=��>�"�:�����UUU��ߖ�~�:?Sl��2�����\]@B#��^�ԓc���NmIy�r�5E^����
m��5zy��b��Ix����ԧP���f�*�忧�;������[o��߯ ���6<n�(ʴ髫�Ʈ� ojK�=U��{�?����v=� 4��-k���n��I�|��J���i
�BB����J�}`,�onc�r�IM�����#�:�ǀv=�ܮU|��=��:�/4�0��������Sc�ܪ�F��� ;z�[#�s����'p[>����6�M�������Ԓo��Χ�.(����L�8��D ��u�cRN_w�ԓ��B�T��],�����$�_������zT��?qo�y`�:=M����wx������9Z�<�|� ojK�$z�]��.���ʶ�V5��(v���]\�@K�hb��J�M���ѕ'E�v�����b������s���﷠OB�v[X�S[��v9~�r� �=��"���:����NNs�{�C��b鱊����� ղ<�lxc�`�QT�5���qX��=�Ur�����5zy��㽺���hkA0��W+��r��{׀yCci�
�*�ln��6<�+��o�y|�{׀j�^�|��4XZ!橋5���M�]aVæsM�O9�j�i��
JF��K�3v�I]+��v9 }���j���N|C��ށ�~�|�eSX�� }[%��G�unǀv9~�r���N��\�IC���������unǀv9�6K�>Z�Q�:(-۷�ꪪ��O<|��|���?UqG=�ݩC�m�j�*-�wo �r,���9_���R�~�}�߿cRO�;�jI���J(-H0ΖI4o�zڦʶ\;jY�j�F,q0#<�[z9�D�t�!�O�x����0p��*�XdN����8Y\��e���XF�*�h�UD���H;����ۂG%� �X�W���8F�yư6J�0�l-fa�
�:��-�S@mR�tSK+���i��v�=v�-Fq��顙�3/2҈�գm�96��N��oL�7W^R�F(mv�!�Rոe������l,���mw*��Zٳ.)V(m
$&��,��.�BU�x��a�!�l]61[��|��^�dxV����s���,�<
��鬦7J�[��5l�?s�I���7��X��/?W9U\Hճ͍�QWe]M���5I�v9�6K�5l� +�֥Z��WCJ���E�|���[#��+����O<ki�z���+)%v���/ ղ<�dxc�`���%�lG-Ŏ��<&�7K���o]��r���_����ܙ�c�?�����W�,;F���Sm�_�<�H��"�	���|�T��+c&	mנx�痿yg8C����BT���>Ƿu$�秳�'��<��$������Z����k�z?y`�K��9�%�=�y{�x�
Prӧl�-��`�K�"ݏ �H�?r�U����g�� ��~G鼦7K��� �v<�UW+�~���{_����]�d*�4�n�Y۲�u��a��&zܔsI��m����Z4i1��'l����bhiiv� ���o@��`l#��UW>A�'� W��/U� :J���'\�=�����ߏ� ���� �H���Ų����+(I��"�G�Eݏ�ܣ����Q�	Up] ~B�Ȅ�ݸ�L�f�3 �NJd���.*BG(v	r�s�v�	8a�@�`Lڬ(@���,��"�m�E5�D�(���$�`
`@�d�K�� �$���4��	5���4�s��x7:��
nL�|%�m���1⚦6�J�@��
�P΀؃��q� ����Ab pDC����"9S ? �N�~�9��s��n���blDc��-]�-�z��?�=����ߞ:�,-�xiE(n&�:E>7v��� �\�W��=�t��� ��7UR�eZ-.:i������б.
��]n�3�x���1\K6�VX]-%c)v�n�] �[�x�ذl%�wc�"�<wB��bt���m+��a/ �����b�'`J���n�e�v<)#�'^ŀa/ �Wa�L*쫢��n������$s� &�^�Ur���@�@ �E8)��r/��!��7���l(j#u��b�	���I/ �H�s�\�}��O~[G,���CR�yˇ��
��w�y���>��ٛ�a����9�0��m̮(i��������K�"�<u�X��6�1ӷE�j˼ �Iy�URG���H� M��kJP�m�T�Wm;�)#�7^Ň������׀��x_IC��n�][Be����U��� zx���K��\�8���<H��Rt�Ӻ����	���~��{����X�ذ	ʪ���w[/N�^�u�wt7�>�mUvvJ
�u�� ���rKc��k���E͵Wl��G,�B�e�ffVYM�t� Gv]�q�]m�葇KI�:��5���1nے����M�Σ0��w<�;�9�������5V��H7pu\8�yhx���\��O!۳����κA�s^6�Q��ǭ;�Վ�1˲����F�v�h���k��P��c��F��A��B�̸���$��"��-��˫�_X]��e����q�"�Kq�X��%��~��$Ł�C)�yLn�e�@7���� �{ n�^��kg
AWe]N�wx�"�7^ŀ���I/?N�'O�:I�-�{��[����nŬ��, ݄�?U$o���<���>��|�@nk���NNIȾ�����޼-���"���7C�St���Yw��^��UW<���	��M%��	,��bE�YlJ�;[h�+5��Mz�K�����0��f��t�G���n��WVӻ�"�ǀn� M�_�r�@o���
�G��۵WVб3s�jI�c��¨d���eD\��Ur���=�z�l��l� ��*t�bi];�i;XR�d�����K�}�H��I�M�t��x�%�l� �r,r���y<W6��AWe]N�wx[#�?UI~��-�� vIx�i%b�Dʹ�m���'8� P�	aJZ��]hm�MЀA���P,,tMu��9t� ;$����<��x�1z��mZT��X]�< ����`�E��A��6�:=M��NՖ�}�^�r,7�uUT6�Ȱ]�<u��)[������w�}� �r,Wt��9U��[�z���Q봘쫥i'E�X�`�� o���>�E�{΢��$m�['x�n���ν!U]mcZ\6˹э�ʃߧwN��v�j�i������נ|����`�E�l��S���*e� ����`�E�j���Nr)����HD&����ݺ�o���"�5wH��K�
��ZwhT�J��v��"�5wH��ɝI���;b#
)������=�}�j�I�^շn���X�� }6^�r,z�,�U\�-5x��J��R�1�"ļu�5!.�w�|{v3Y�uVOd�R�'E�luv��-��O^�r,z�/W>A�� ���/+N���j����`ױ`��x��y��A]�O��*,�ذ�֫ �������T�V2�Ҷ]ZI��5wH����.��Xf�
)1��7J�Yo >�/ ���ԓ�c���}y��jH��t�P���n?����*�v��u�h3�ʩ��`�D��Xi�M�R A�Ij^B�̧��v�*y)��:�su��Nù�,�G*�r��ۊv�"� �'n��;&�XѲ,���ԛa.�2RK�u%��&�9W�1 ��u���4<uC[��c�t;%�HG<n��э�2Z�� \��qk��5F�u�Y�Ke��s���	c��;���R|�i��K����ʳ� m`�� ��	PB�k�i���������Pt�离�ݸ`�ذ�؞ }�/ +鰴�Ш��ݻ0��XV�O >엀w��}8Ԩ-�N�1%v��؞ }�/Uq-�_�u�, �&���F6[�ӵv��ʮ%��� ����;ױ`[�x�%
+L�l���w�}�p�;ױ`[�x�d��n[�;E4˶6���s�+�M�:V�R.X�:4J;�Eq	���c{��6ڧe:V�t�ـw�b�:�H���xݗ��T�V2�Ҷ]ZI�ԓ��N�JurQ���'}ϳ�'{���;ױ`�(�cYLn��� }�/ ����%���C� �Ȓ
T�lWN����U9?}��$~����x�d� �ͅ�v�@�t���ـw�b�?s�%������^���:�}�������mKf����*4&5��e[���+�MDMr�*�͘8f��t����~�����xݗ�{ }���(�ċ�v����%��*�#���n��uM����(�hB�T]ۻ�>�`�ذuNb�A4]!��@٢�fG+�d
5K��L�W#��M-b� ��(���>�q�$����v@��Տ�N�M�����qn���5zy< ��^�e� �ڊ�*�ZLV˫I;XT؞��*�s��m�ߟ@���z�, ��sce�-Ri�3Ƨ�[v�� ޻�hJh+u���0��p���Lj�ҠWi�.���\0��^�Ur��Ry<V��H)Yi�t�wo ���w�b�:�����<������zf�Vºm�0�<��؞���W9Iuo���_��ƥJ
�;�Wk �݉���s�'�w=��h:� ��Z�
���H@�
R����������=��I?��Ř/�.�ڻO >엀w��w�b�:�bx�8_7l�L�i����.��A!��_cVx�r[I��
�l���-݌�ش��n�v���\0��XV�W�$������t~���[�/4�K*�0��XV�O >엀w�ឪ�N)��'��vl���kn�@����ݒ��\0��X{q1��6�@����\�]�z��_��{���������3���8�j:Z�wx{.z�,�v'�vK��*������r5�B�9�!!���<��*�t�k�B����|�'�c_#�b i:M�1���7
|0~0M.���E���2"�Z«�r)�`R)R+�+(��U��e`Hej��.���r���5�����U�tC,B�hSD"H)"�PҘ9$�XB�"��(����aE:"E#���0�Q�#�pK�Z2 s��	b��H���ؐ���Ri��	RN2�I���0m=���~W�������~���H�N�C�   �������  h[�j�  H�    V�K�j�lr4�hv��͸%��Ѱ��4�^�K0Ǟ��B�Q�m����1��o n��QZ��g���`�y�k7N�,�h�.�,m��k��NK�qӫ(��ȏfj�Qȥ��Z#Pf]Ins�6�Ĩd���M��a̹����s��� �"kJ�%R�8���\0tv�v����y�)lv}]I�V�]��D�
�kX�h���;��[2)�콱lh2���n�8!SWi��q0P���ٜt�xG<�v�
��)�{`��@5�V���l�u����-�-�B�X��da�%hgie)IGb����ݴM=Gb3�,�;w3�ډ�������2F��iY�gv��9c���Oij՚1�m9���L�[�R\�M��8�Fvh�tͮ�A�i�
�,���SU��\�FJ�R�H���)Hx'�#��]dsݸ;9�j���e�>xnZ�DmiZ+*�C �e��ؔg�q��q�d@���%pn�a�\*�u�`��[���v��=�-�sb1�Jgb^��I�$;i�j�C����;!��e��Җ�vx��)�ld��t� CnnWR���HM�E��@���Z�B{�n�v�U�x�(A݁^Mڗ��<Tr���&��/R�&��!��a�-ɒ�����!;5�Hn�cS$�[m1H�z�yM$�*�W��貶ʲ��fp/-Ɏm�$�P��j[�'^(&�HB�7rlc//6��b'1j@��'��Z�(��Ca��mpa��!���	 �(�UC<�q��4�l;�y�5�-��b��z������]��N��*�`�:1�� �`�۞-c�M���j8*T5d�y�0s�:�sy��;�'�J��
���zea�m]�"/�lp�m5��[�;-��mFte��mޝ;��Ί�`x�/Ji#�SJ9A`}��¦L� aA�� L t�lk�zQ�/@� �߱�aŹ�s	p�vðU�1�sB���9�n�-bˆj�rGWQC�P�cVye97yޜ)���nNB�:�ԄNz���sm2�c�&���*�6y��I6��q��qz^�:��ݴ����p�wG.㎌Fc���R^�� ��Fm#]ex��ugX֝�;���-D��gR����bSh�Wa�I����g]N�9�t65�u�pk������$���N���h��t맬�ڰ��F�#W/Sj;�'��Z8ֆ��[�Q��ݵv��lM�ǀ|�x�[�< ��_�~�Us�$��q�߀(���)	+��un������`�b�r�� ݯ	��K�M"�]���k�X{.�ذ�؞:�I@V��ڢ�ݬ�ʮ-�g���ջ��������
�x=M�[E];I:j��'^ŀun��	ױ`�`�+J��ݪLw|v���-�;fP��I�m,f��\�@s�!ؖ�"�uSA�X�l��mݯ��'��'^ŀw�����<��
8�<�&�A���RN��v��'���#"�Q���#w���>��o�w�RO�9�{��)���=@��.,����{�0	ױ`[�<u�XSd�ݰT$���v`�b�:�bx˲<R��x�;�b��(m%vRWk ����.���\0��X��Ņzyq�e���`�gq�q�XN�����~#�ܿt4m!ǃ������"g�Pt��l������\0��XV�O �Ih(��� wn��ˆ޽� �݉�.��ܤ��ޣ��մUӫC���u�,�v'�䪔W(8���*����g^�e� �ڊ���+e��n�`-ry<�}�w����[�<��
8�<�&�@���>]���`�ذ�؞��&B����F+s�riB7[-͊X7Z�Y�۬p�e��R�(V�5����q�����]��7}~0��XWv�+� ��y�{��n��lJ�=���Ǿ�NN)���:��x��Y��I�1{�6�������"�xx˲<?W*��w�y`�y`��M4:���ueݻ�� �=� �^Ł���s�����r�W>��� IB<�!��wv��ذ��X��<��;���ktm��f�gp�%�چ�i��m1�SY[T%M�ZJ��`��-`ջXz�,Wd������,�^U�v��i�Wm���j��>]��G�`�س�UUW�l���(�`�ݏ �?~x��X~�Ur���X^�O ��*8����Վ��G�`�ذSbx��?~x_����킡'@��Wk �^ŀj��>]��G�`
���wؗ��hbz]�$�i�L`�]X�� Y�.�A��8�������T�q9��@�]H��W��a�Iɟfw^1�[��P���o.���.V�:�Q۸Hh�rfj�I�6�1vil��7&eH��CTcpݜ�8���j�6��%����'[x�=�Ƨ�x���C�L ��rp=Ai�l�nJ�����bq�8^�s�N�yD�����:kھRtYp�[w$�qM51�f�f��v��<�B5�&�l�0�� 6������ ��?'�|�#�>�b��s���`ڂi����L�V�v� �vG�}ױ`��0�^ }�#D�I!ۺ@�ݼ ��p�ܮs���O+�:�y�nʈ�j�*��&+v�	ݙX�د ����I�����'���˚�M��u����^{<��g�;�+ �I9���b[�v�&�&n'l��t���(M��9D��rY�����z���ó�bl|��W�[<��v<wfW�T��=��t���U��K1nƤ��s��2M��]jg��I�����wd�ݠT$����&ˆ }6+�ܮ%�=�ul��;)�⢁4��V�n� �lW�E�<�ݏ �.�y�i]6�e�m�W�E�<ܪ�������د >ӆ�*���e�]5wO��|�k5�ӵ�P�C@n�%L��v$�M�Ή�� A�m�(v���ݏ �n�د �lx[��uit�-�x�p��\��l7��+�?/����v<J�QS��Ze��+v`�R��ǆV|��?-¸�B`1�	bUJ�8���y�zK��ب����bm���w�E6< ��M�`�R����l)�eҫ��ݗ�lۆ N�/ �6<��IFN����7={r����x������lZB����7FSeX�^������V�gm�=�x�	إ��ǀݗ�l�G	�ub���0�	y��M��;�/ ޽/�*����ջJ鱦;���x��� wv^�n� �IA(��v�;Wo��%�z�	�_���}��u'�GgQ�cX��$>쨂촊�v$�w�lۆ }!/ �$x��x���	 ��V�M���n#�!5�I�D������Z6��(/[+2\˰�l����}=���ǀݗ�oe� ��TQ���)6�Wl��:�ǀݗ�oe� >���j��ZaM�S��U������7��HK�:�ǀ�ح;�T$�i�-]��� �B^�6<�l��z���Ei]��+n� �B^�6< ��c�`����튙����N�Si�Z��Ʒl]s���WN��8��2I���vg�8:ԝ%����8� ���W@���7$&J*\��5�!]-��mm7Z����9����9_�N͢FP�g[O<]&���ՉG�[�����T���S�GW�v�X����@��RayC��c��ݎ :=�'ۅ����J[���5�tʵ)Fؽf�+e9��5�], ^m �1nH<MaK�ѺYa��k�Qi��L��
b�a����{淪�we���|��z�x��!$��(v�� ��c�`��[#�
�eEE�؊t���w�v9 }!/�Us��ߗ�~x=�׀M�Ue;T��]]�;X!%��G�$��Ȱ��EL2�m���[#�=�S������ $$� ����MD����62�X��؀@֛	P���A%�K�oX�G����J�n� l���"�		/ ղ< ��+N��$�	�廻�;�/��0��+`-R�Nm>PG��n���^�� l���s��H�q�x��ZWe+I'k =�޼V���D��x��� ��8�v��cM���wx��Q�y���xc�`���)*Ў��v�;n� l���"�		/ ղ<d�n��Ro�c�L��j�n��Ȝ�Jv*Uw��	�� ���:�e��-������z{� $$�V��d��M�Ue]�v�h�Bv�BK�5l� 6Ixc�g���H�<�����Rm����� l��u���C�UU..UDNL�4]Q54]&b�<�P��#��
d@!��HH��j�\��>��a�Hd~"ҡ�)�+�� �m��B��
>���l��g�2��@��b�2�`�!@��:�&Q���0��!L�Z�!�ҷ.i��C!���D ����H��9�T�r��b�;�q �~D�aC �8mL"X��% z 
 ���8���b��K�>ZH�0��)�t�����/ �r, ��/���(���=�i�Z���'|�wxc�`���[#�	�^ M����*srg�OVt+؜b�E�V�F����;�c�Q�G�؄7bV����������/���W:�~�,/~��;���eݵc��5l�?s��q ��� �?y`������I$5v;n� l���"��G�{׀E=�ٴ@��N��;m��~�qo��Y$�����'/;�jO.<!�Q����v�W�e;T��]]�;X!%��~�����~����"������x�q��Vt��6�F��M����;aI��!t�ŘV.(���q1�)6>4;�V��d��v9 HIx��7wW˦�Ucv�d��H�?y`�{׀j� T��uj��1�X����X!%����ʪJ)�</{� ��RP+N��I��		/ ղ< �%��E�ul�C�J鱧v�V;�V��RG�v9 HIx\��"�b������� ��U*Ad[�9�`�%��:��{��Ut�+;#��-�����}�?d&�Y���{i��u�hۂ�XD���r�1�[h&��9כ�q��5�.�&�a���k��7Cc��[�k">g��{<n4v��*jY���e����\0:���!�mY]�=���' �O1m�<YEL��K�W@��Vz��p�eH�o��t��1�H(�h^ #�]�gYM+��Κ4�Y�:�x�i��!uV՝�e��'N�4����v�=�^��X!%�|�)�< ����uv"�;Bn���;� $$�V��d��M�PHʻT��v��`���j�H��� �s� ���ELfq6>4;���W)G�����ŀ/ �n����||v]*�]� ٲ��S�<� ����5M� >�������=k�և�3r5r�V�[���^��	Z�ط2c��4ur/.n���l{6^�l��\��O^=Ƨ�(�vQi$�`e�tUg%r����������xǱ`['�ҺliݻH�w�j� I%���ʪ��s� �==x'�-�i�ҡۻx�9U\�\���{�����`e��ǀ������t�	�ۻ�6=� ��/ �6< �e��T���(�:*��ެ*m⅌�!4m�NdL�\���p��;˛�����y��T��M����s��y`�yQG�M��+��5M�=�s��zz�	�<�������٫���݅_�J�Wo ?~���6=�\�s�*��
���V���ԓ���5$��&��M��un���b�"$��j� I%�8��ݔZI;X*Ix����^��X���_x�oV%�"!����9��w=�����
�u�<~�Ȇ�v v#%�.�
a[�黾���ߞ I���b��Ix%	m�I]�C�v�we��s��ߟ�, ������ǀ7h�]]��V�wj����X��/ �6<u�X�HY�j��h�Bv�?r���S{��~����<u�XU�p��(R#��wA�E� Pa��Rjp�S��n��>��i�� ���;�T��ױ`ŀI盠|~�5��e(Y��)	D0D6�uɠ�J�KnS �lD����-4k=�۹�`�>;.�X���H���X�T����	�e�m��vӵ�l{ }*K�5M� �{ l�[ n��	���%��Ǉ��r������ ���� �M�.�WM�;�����lx�ذ�b��Ix%	m�I]�j���b�?s�U=s������	ݗ�{��m}N�#�4�M{���"�ʶ\;\U�A�7˞���\�}��覰��zy�ڴv\����!%ټ/�<���+:	�a�s�nka�y/A�cNM,���,m<�*�k\ȁ������+�]�Hك�.�vsӫO�К�A���>��~�)��q�u�f���(�m(QB�bR�C�B�R2YR����@�Y�ᝋ��l��sB\�5-��)9'i��altt%������u�ImKd��@ـd��:�Sb�$����u��JЛwv��s���T� ���ʮ|�c�X}^^,��l�Bv��/?� ��^��,u�X���CYN�v>$�� 'v^�{:�, �eK�'\��݅�Ӳ�$���ذ	ױ`�*^�/l��C��۴]4�wi��:�, �eK�	ݗ�wve`mo&����\s�s�ɡ��gL7�'�|>)>�����'Aͻy.좄�;���|�������;�2�|������v+�Ɲ�v��� 'v^J����UU]���V���l�x�Jt
�w|)����̬u�X�ʗ��/ *M�Q|w˥hM��=K�s� ;=^� ��xwfV���B�v��j�v��`�*^ N���+ �{��.�_}k`�vp��[��P��Ӌ�'N&����c֑�LA���O��M�V�����~��xwfV:�/��ʎ��rZwv�Nˤ���;�u`w��X6T� �l��${�Wt_I�g7ɩ'y���I7ΝΦD�`D&P4���7�gRM�ѩ'/ċ` ��v��/ >�/ ��������r��{��5~�?�+C���v��� >�/ ����7�b��T����8~�q�q��f��$�#Z)��IsmCR�8y2�7Kz.[�=�]�����w�wve`ױ`�*^ }6^ T�J�vr��I����{{�Ig�׀���ݙY��#��K�YN�;��hN� vz�x��xwfV�{��@�P�ʰ�uw��_��gRNw�ѩ'>�;u&�C�DH�P�RA� Mk>���I�c���r]_;.�(N� ����7�b��T� �l�II(���I���O\�5ƥ�`�[�٦	C8�nb��[5�i��ƙ�����ӻN�ݸ`�*^ }$��ϐl���"�<PLj�Xӳ >�R��%�ݙX��X�o ��:mݷhN�����̬<��<�o�׀|�t�R�M�E+�wxf̬z�, �ʗ�M��ٲ�c������m�`ױ`�*^����ԓ�s�5$�Q�!P"@&0p'�$r��|� F"�Hb1H�k�fY��[R0��,
�:GS$B02��˜	�D2��Nb�"���P0�|51 �R� B�ր��4��t��e;Z�ٍƄ���!�����Q7�ʉ�i"Fgh\F��%	[��������aK �A�4
gc)F0$"�i5>U�0�@��&
�Q�`D�F3��WK>C�Ió�J(iL%�!؛L¡��ì�ٔ>������갌 F1,1�Fhv�ӵ���� 5�$�&I9�8    �`m��6�v�� �E��� @+j    %G��
ۥZۤI�].����Y���Qb�\��R�0\�n�+&z&��cqT��+�2^Ż*�38Y��}[`�av��g�y9�U�e�9����T���e�t��j�\Yl�4�핤&W�?��USo�b&`5!VPmj8
�\�5v���m�ŸE�q-Id�Ԥ��Z�N֧-�7l6�S�H��؟�v�ú��7s�ϣZe�#śV���c���=K��]-+e��(�V�6mV�gr�֝��˴xG%�Mhu�{���"���Q�#]u�72v�+��i��ۋ�-��[+�p��o���w�����Q���Ү�m���X����lci3&Vl�,��po��ve�*1���ǣeVBi��[:�_5T�Z����g��W&Ҙ+s��2ǫ'.�.\�F�%j�[�����[i�z�i8:�9�aEbrƔ�Қb���@u��SVΫ�(�{ �mLj^ۃ�65��լ%�D��㎷Z&���Z8϶�{u�9<v�N�n�<�b�2Z^�E#�C�앆���[��+��1���if8���+�d��&:QN}Yf糂��ְ�i�P�-�e��
bܙ��Ͳ�m��E�3��j �E2D�n�v4SV�u���q����kb�y����s@��jU����!lü�6�	��k����u���Te���bLg)�rd�nB�[�U�v6�	k��[VI�zW5X����R�h��gq��JG�N�pz�5��m�g(�	zq�E[mӷ1,�fpl�[S/���.Uj��� 8ll�U�Xӂ�Y�ZVg���h�Ҫ�S�+)<)��q�kmԡ���#�-���ʌ%Ne�����X�,m�q����5ejn�g%��-�UVRRw �v�6���\!�.bB�n�e�f�K�h*Q��@r�e�kS;)]�t��)�W��P:�� �<�d;{�諀5��������b�����m�۬���PuۮnS����ХlmAALŭ	qQr�����F�,B�) �wG`�3��k�֜��a���6e����F�m�ml�L�I#��v���sq��e.Xj�j�4fQb�tCj�n�R���
5Ld)
�׆Q\Օ��Ĺ�K�B"Z��v�`��e��*؜t:�uYEV�����K�O��O�<>|>J�m.9l�!�ڂU�ۤΌ��:�rmg�uֵ,z�ߺ,f���ɵ����~�^:�,��+ �{��@�P�ʰ�h��]��b�;�2�	ױ`�*^s�g��~������j�1$�`����N����W*�#����=�y`i$��ծ
��ӻ�u�X�ʗ�N�� ����'i�a@1�(�N� }����b�;�2�	ױ`u��n��9ujպn���������8�q��h;1���t��5ڣ�Ywv�N�v����u�XwfV:�, �eK�>R	0A(Cv �s��I>�;�XWH�E��DW��3ۀ�R�	ױg�
���m��ʺV�M���� }����b�;�2��D���N�m��'kܤ���x��,�fV:�,kt�B���av�C�w�N�� ٳ+ �{ l����+ce���m�wv�H9M#�$H��8lFiT�z7I�[6�v�ڨk����t�$��f̬u�X��^:�, �l�[��Į�N�;��'^Ş�r��RA=S׀{\��>�2�	�b�QE4�l��;Xݭ��N�����tX%L&$˗,"Q���jO��w��Z5$��箤���ٜ�L@��/���ӷ���O-�~���'^ŀ���)���7`��x�X���^۞_ o�^�/������.HJk35�LĦ��%bE��KTGJ���E���;p���#�`���+I�ݘ�ذ�T�u�X�`H	Y˴�5j�
�`�R��[<�	=~0	ױ`��
�K*���w�Eݏ ݗu�X��u�i�.������'o�UʪR{<`�<�v)xʪ�UDM+*=R�}Ƥ���;3n�%t�v��0	ױ`�9x�ذ�p��Guj�C�N�W���*�
��66z���k�^Bd���-� ʣ0�P �v�,��j����b�����}�M&�X�%��g��Mı,f�?��{�*�e���O���5K��}t���8���'��_��q,K������n%�bX����t���Ȝ�����W�cn K�{��%�bX����Kı=���I��?�!���~�?gI��%�b~�}��7ı,Jvr��̹��0\ۉ�g3I��%�b{�ﮓq,Kľ麟��Kı=���I��%�b{�צ�q,K��ޒ�<m�n�3��\��7ı,K��{:Mı,K��}t��bX�'}�zi7ı,Os=��n%�bX�U�A�'Y�t��m���k�vvj�Ÿv�V��7���A�b���`E�0%�ժֈj��6�:۬N�5������ȓ��M�D���c��n��������b]u�ɇ�:�� ��k'�_��}��	�2H �V�GM/e���9�ϳ���(�Y�jwR�W;&�,!#f��t0E����b�"�a2{h��]�rk%������:� �m�u�On�s;����� �tк���"k�U����M�HM��f�tr%.Qa�C�
P�
�fL���ϓ�Kı?���cI��%�bw�צ�q,K��3�]&�X�%�{�OgI��%�b{���q�̙pc3&0Yq�i7ı,N����n%�bX��{��Kı/{���7ı,Oc��4���1S,J~���Lc6�d�� �:|�5�Mz~=���O�,Kļ麟��Kı=�{��n%�bX����Kı=�2�� Z�Ha�^�|9�9��移��"X�%��s�Ɠq,K��}�M&�X������~Ɠq,K��?��*j	���>^��צ�=?��i7ı,N����n%�bX��{�i7ı,K��{:Mı,K�~���tˡwd�Z�pf��Іw0ܔ�����h�JXе�ub:%�	fs��I��%�bw�צ�q,K��{�Mı,K�Γq,K��9�cI��%�bSӗǮe�&a���K��i7ı,Ow�٤�5�k���b^�S��n%�bX��{�i7ı,N����n%�bX�{��l3�ٜ��nri7ı,K��{:Mı,K�罍&�X�%��{^�Mı,K��i7ı,N�����fd�f���I��%�b{����q,K�ｯM&�X�%����4��bX�%�}=�&�X�%��g����<A�	��O���5�O����7ı,Ow�٤�Kı/}���n%�bX��}��Kı/����$��ʬ�41�B�����9lr�+�8��۱nd�%�[e�x'vjś��Kı=��f�q,KĽ��gI��%�b{�����蘉bX���߮�q,K���7ߡ$�8��!31s�I��%�b^�ǳ��Kı=���I��%�bw����q,K��;�Mı,K�y�.��8���1�\��t��bX�'����7ı,N�>��n%�2�'$C�H���@�
���#��ND����I��%�b_�t�t��bX�%���=�,&1�$�9�n�q,K�ｯM&�X�%��w�4��bX�%�{:Mı,K��}t��bX�%=9|z�ٜL��ĸ�f�q,K��;�Mı,K��=�&�X�%��g��Mı,K���4��bX�'N���7�4p�<�S1[���;r[��ж��[�"�\f�嫭��1��ID�5y���bX�%�{:Mı,K��}t��bX�'}�zi7ı,Os�٤�br'"ry?{=�0�ɲ�^M���Kı=���I��%�bw�צ�q,K��{�Mı,K��=�&�Mzk�^���ﺃH�� |��%�bX�����Kı;�{f�q,KĽ��gI��%�bs�צ��Ȝ�Ȝ�����[��ԅ�:�7ı,N��٤�Kı/{���7ı,N{���n%�`uI���i�^�M{���n%�bS��9�'� j�a3]�y>�Ȝ������7ı,N�=��n%�bX�����Kı;��f�q,Kޟ��;�|�Ƴ~X�j�4.�+M�\�j�d&�S3B�?z>�u�_�v/,�-��.3�g&s�r%�bX������Mı,K���4��bX�'}�l�n%�bX����t��bX�%�d�o�a����9��n%�bX�����Kı;��f�q,Kľ麟��Kı>�u��Kı+��z�ٜL��1n3���Kı/y�gI��%�b_w���n%�bX�{���n%�bX�����Kı>�d/���
��_:|�5�Mzo~�}|��bX�{>��n%�bX�����Kı/y�gI��%�bx�$�¿&˵H\m�O�"r'"r}�y��Mı,K���4��bX�%�;��7ı,K��{:Mı,K���/td�����*����.-�d[�t�����''GkG�8�3�#=`7j��r�j�]�!i+J$Vl�f��3���۴qu���&4��;H�*���,!�v��:y�S:�Rm�����bj���5�L��]h���+��n���˧qű�m�0�:�l��6㠹��/u�#�A�l��ݵ*�m�>=v� �{m�9��F-/ka]]6���WozN�~���t;�N����˿�h���53@�^vp�iT���`�1������e\��c..�eƖ�[��xr'"r''�����xn%�bX��}�&�X�%�}�OgI��%�b}���I��%�bSӞ�-�a�`�mq�O�"r'"ry���ı,K���Γq,K���צ�q,K����M&�+bX�'8��zmԆ3�y>�Ȝ���秹�n%�bX�w���n%�bX�����Kı9��zMı,K�u�>SP�v�t�zk�^������&�X�%��{^�Mı,K�﷤�K��31�ߧ��7ı,K����_赍�[��O�"r'"r{�k�I��%�b�{��n%�bX����t��bX�'{�zi7ı,�9'�x���M���nр.��H�[/,�263�s1lRZ��:hѪ�ר�&�0\��9�A$N{��j	 ����t$�H?s��j'�X�'��zi7��Ȝ�x�>ski�s�y>��ı/����7�F
1D�@"�F
Q A��Ә��bo~צ�q,K����M&�X�%�y��:M� �,K�=�$��f1ns0�fg:Mı,K���4��bX�'��zi7ı,K�{��n%�bX����t��bX�'q�����I0c38�1�fi7ı,O{���n%�bX������Kı/����7ı,N����n%�bX����)*\5F����Mzk�}��_:|�bX�
����t��bX�'}�zi7ı,O{���n%�bX�x���ims���*����Z�'��]m��s�����E�|�PfYp����j����D�,K����:Mı,K���4��bX�'��zi7ı,K�{����^��ק���zo�SP�vX�I��%�bw�צ�q,K����M&�X�%�{�{:Mı,K��=�&ॉbX�ܓ�-�-�.3!3�c9�Mı,K���4��bX�%���7Ɓz>�q��a5��{0?7��E�b�� ��Iޘ/7
a��
`��!��B)Q��+�dpj4�P�D��`H9�fCL�Ez�Dp �	��\�p�b��50C)�dfB�Ft� ���@!�#�<X�n#~@�EL9��P����ʑ>@� P��"��+�%�pj�9@>B|�49`��1�jeP�P4�t:L��@ß�x��!�7��bF
&��LW�^���r�8|� `8b�T��ɏ����e҄V��p&$��#�L�_�����P���ʂ18 R���]@@$Q$��P���� ��U~�蝉}�Γq,K��}�M&�X�%�O��[�b\�4��I�q��&�X� b&=����7ı,K����t��bX�'}�zi7İ? ��O{��M&�X�%��߈o���I��.���^��צ����t��bX� ��צ�q,K��}�M&�X�%�{�{:Mı,K�x��m ܸ�h�Kb�f����f�3ӆ��]n�A�ZF���um�KX-:�3�&�X�%��{^�Mı,K���4��bX�%�}��?*O�b%�b^��~Γq,K��;�Ř�f2I���	q��&�X�%����4��bX�%�}��7ı,K��{:Mı,K���4���Eb�"b%�OӾ�(��d����:|�5�Mzo}��:Mı,K�Γq,K�罯M&�X�%����4��bX�'{��zrŻn�|9�9�����n%�bX�����Kı;�{f�q,K���B��-RT�Am^U����)���HF,� -���Sl��@�D"�B# ��%���DM
� G�܉���s��Kzk�^���ޛ�T�(�@j����X�'=�z�7ı,T��Mı,K���t��bX�%�}=�&�"r'"r>�$=�1Q��Pt�Ci@��l#C�tGTa�eE��!k�&,&n6xm\Ź-�.3g9�t��bX�'}�l�n%�bX������Kı/{���?O�b%�b^���:Mı,K����ꎆe��-��'Ñ9�9<���7�,K�Γq,Kľ｝&�X�%��{^�Mı,K���>I�Sh;m�O�"r'"r>y���7ı,K�{��n%�bX�����Kı/{�gI��%�bu��XA���;�����r'"HID�~��&�X�%��ߵ�i7ı,K����n%�`~��&=���t��bk�^�O����s- �%�O:|�5�ı;�k�I��%�b^��Γq,KĽ麟��Kı9�{��n%�bX��BE�SUw�b�V��l�;�媭h�9T�}�L�t�]�p��v�-�og���(�D����#s�q�IϱP�Ul�Xj؄{D �J&��k���盧.Nk��?)�n�~17m�r֎�9ԛ9�`��Q��F9ۘu��+;f+���&��E�F���Yݶ�.ֳ�Y��7nC*�̇'G�# <��p7�O0s3
R�[�M��H%),Ljej�7�9�}���9;��|�T��Jk�.�!hY���x�hp.HPnI��,ͥHJ��U�YI�YEj7ޟ�X�%�y�3��Kı/{���7ı,O��{Mı,K���4�9�9������s+1mۼ�"X�%�{�OgI��bX�c��4��bX�'}�zi7ı,K�{��>^��צ�?����o�SST��n%�bX�ǽ�i7ı,N����n%�����߽�:Mı,K�ߧ��O�"r'"r>�د�k�M��Ɠq,K�ｯM&�X�%�{��:Mı,K���Γq,K����|9�9��}��֎�e��%�s4��bX�'���Mı,K���Γq,K��=�cI��%�bw�צ�q,K�绯ge�c8����ɲ��F�gsh�SL�tmnp��ım�K�%���Ks��y���MzX����t��bX�'���Mı,K���4��bX�'���Mı,bry�|��|m�ڤ.6�'Ñ9,Oc��4����"� _�ة�O�X��z�i7ı,Oc��4��bX�%�}=�&�X�%��w�,�Ѷj�'�>^��צ�>���8�Kı=�w��n%�bX����t��bX�'���Mı,K�����.�-���'Ñ9�9=����n%�bX����t��bX�'���Mı,K���4��bX�'q��'�s�K��^�|9�9��==�i7ı,T}�w��n%�bX�����Kı=�w��n%�bX��$�����D�smk�&��Mqt���-�M�Lh��f����R�1�s�.�2k�m��M��,K������&�X�%��{^�Mı,K��}�&�X�%���{f�q,KĽ�����R�0�s�g8�n%�bX�����Kı=�w��n%�bX�臨i7ı,Oc��4��#bX�%>��nq�rL�q&%�s4��bX�'���Mı,K����&�X�z~T f2������SF�n'�k���Kı=���4��bS�9>��'�~I�.�6��O�"r1,N���4��bX�'���Mı,K���4��bX�'���Mı�9<��|��v�\�;���N%��{�Ɠq,K��=���M'�,K������&�X�%���{s��D�ND�|��{�"U��v�񒛈5,[N` ��[Xk�F8��B�k[z�XPh�5	nΟ/Mzk�^����&�X�%��{�Ɠq,K��}=�I��%�bs����q,Kį�=���b�B�n�y>�Ȝ�����q��Kı=�Ol�n%�bX��}��Kı=�k�I�#bX�'1�G��!G9��;k�O�"r'"r~���i7ı,Ns���n%�bX�����Kı9�w��n%�bX���=������O���5�s���n%�bX�����Kı9�w��n%�`j� F�@VA�	F�0�`P�DI�����6�x~�;��xi7�'"r?���Wص��6�y>��%��w^�Mı,K�;����'�,K�����n%�bX���O�"r'"r}�����B脣�̷e�sO6��q�\�j���P]͗1g��ㅍ�r2�R1��t�zk�^���?��i7ı,Ns��4��bX�'9�zh?蘉bX���~�Mı,K��7�sV��c�<���צ�5���&�X�%��{^�Mı,K���4��bX�'1�{M��NO���Ѓ��.��N�|9�8X����Kı9�k�I��?��"b'q�߱��Kı;�~�4��oMzk����V�A�(�|����,K���4��bX�'1�{Mı,K��צ�q,K�,�N���Mr|9�9��ǿغ�eemv4��bX�'1�{Mı,K�5��Kı9�k�I��%�bs�צ�q,K���7�Ǳ)�.s�ې�K���yV�k1��\�D���i���^��:���:�bl�8�n��t���s�ϣF�t�j��ġ�������n�$�X������w�u�0�����X睨@�Lٻ��e�j�#k����� f,��1�iYP*i�`
�Q�ms�lTl���H�,�(�u��Ջ<s�f)"Ӧ�*zM�܄�rd��C& y�P 	�<����7g\Ҕv�����9��t��p�aI�۵�ϻtn�.e������c%\�8�z%�bX����I��%�bs�צ�q,K��}�M��LD�,N㿿cI��%�b~�zF?Ř��q��13���Kı9���I��%�bs�צ�q,K��9�cI��%�bsޚ��n	bX�%�I}1o�qK��&l�s4��bX�';�l�n%�bX��=�i7ı,N{�^�Mı,K���4��bX�'��{78Ĺ$͸2d�.1�I��%�bs����Kı9�Mzi7ı,Ns���n%�bX�ｳI��%�bw�!}f̓P�v��^�|9�9������'�,K�9�k�I��%�bs���&�X�%��s�Ɠq,KĽ�=avu�0'X[�om6�;��EbY�7l��F]�K2�����P��M���Kı9�k�I��%�bs���&�X�%��s�Ɠq,K��5�|�5�Mz{����j�5�o�n%�bX�ｳI�m�����$E�! L*F��+ @
�,)����D�K�޿cI��%�b}��~�Mı,K���4��bX����{~���h��y���Mx�9�{��n%�bX����4��bX�'9�zi7ı,Nw�٤�K�D��|��=��ef˵�'Ñ9�'=�M&�X�%��}�M&�X�%����4��bX�'1��Mı�9=��v_e�6�r�c��D�bX�w���n%�bX�ｳI��%�bsﱤ�Kı9�Mzi7Κ�ק��鯩 G4ok��n���Nxy�!�q6�v�N�F��k�i�cb:엸��n)q�$͙�f�q,K��}�Mı,K��}�&�X�%��zk�I��%�b}�k�I��%�b{��s�:K.�-�w��Ȝ�Ȝ���{{ɸ�%�bs����n%�bX�w���n%�bX�ｳI��%�bw�!|�1�B��e����Ȝ�Ȝ����Sq,K������q,}�_���ʋ�˟��p!T�\0��(c��NDξ��I��%�bs��i7ı,N��	�y���s�&31���Kı>�}��Kı;�k�I��%�bsﱤ�K���LD�M��Mı,K����c39�����Lf�7I��%�bw�צ�q,K��;�cI��%�bs����n%�bX�w>��n%�bX���\z�����stH:�ܴ�\,̣^�����7�1W�c�uFW��:w���eemv;���bX�'1��Mı,K��צ�q,K������q,K��}�M�ND�NO�ȯ��A�Vl�^�|8X�%���k�I��%�b}���I��%�bw���&�X�%��w�Ɠs�9�9<��v_e�6�r�c��"X�%��s�]&�X�%����4��c�!����{߱��Kı;���㼟D�ND�x��X��vn�q,K?!;�߾4��bX�'q�~Ɠq,K��5��K��yd�+�J#H��� xPޢgצ�q,K9�����2��-�w��Ȝ�K��}�&�X�%���{zMı,K��^�Mı,K���i7ķ��?����Å�\�.�Ds۪�(Ua Ю101���I���{p���L̙ɛq�i7ı,Nw���n%�bX�w���n%�bX������&"X�'q���i7ı,O����u��.6�'Ñ9�9<���w��?�LD�=���M&�X�%��~��Mı,K������� T�K���݁�l ��w�>^��צ�=��_��q,K��9�cI��%�bw��ޓq,K���]&�X�%���q]����R�w��Ȝ�Ȝ��=�i7ı,N����n%�bX��{��K��=���M&�X�"ry����B.��6m׼�D�N';���7ı, ��k߮��I߿~�j	 ��w�В	"T_�PU��*��PUh*����T_�
����*����AC�A�A`*� E�E��P��B
�B �B @	T"�P�DXBT"�T"� `�T" ��B"@,AP��B$P�THBP�@T?�
����AU� �
��TZ
���PU�*����T_����A@���*��AU��
�T_�����)���6�B�/�8,�������_���0�?��  ��}�E4�  h(4 6�
� kTD ��Ѡv�h�    �H�$R%"�AD�
UH
U( D ��"�$D� �P )@%EB(�     0��A� ��M
k3[+��eL�].-(���y� �P�[��\ڥۗD��:����U.�zs��| �Q��    � � 4      
0���ũ�q�.�.�Q�o /g����7I�v�m^�u=Us��/� �� �E�T��5�}���c������/���)�<U��qN��c�����< q������{�x a��O<���}���O{u��t�������ow��nϼ�}�|�|��(	JJ��:���o|�s﷽}j��W����}�;P�����U�y�=�׶�=�w� ��y���ם�k�	x�����y_m�o�Z�������wY[��ۘ>�<�}����.U�n����}�|�� �()B�
P)U�0�o��n��K��{��]���[;����n+��}����c�p;�W;�s�W\�� �]�˭�������¬�Wi�{�i{�������vw�������j���C� ��*  UR���8���v���}�l���{���]�k���m_c�m{�P�ǀ�s_c�}������x/}���w zs�e�������7�_{���R��s6���q��\ϝ{�v�^             �MF�IUMOS�@�    ���)$��h�� M LE?���C@      '�T�)       ��i%%( FM4�C
D��f��T�7��@�$h�MO)����L)�S���:����ρ�'��|���#�b��,�  Q�� 	���"?���������,���SO�GP���ADF2S_��Т�#ԣ���J
�0:c��F��?�������?��[l6�m��~o�>"��{*��Ps'�Ȉ{*�슇��>� {"P젾�{"��Qa�G�TOe��=��U`�T=�C� =��@a�=��P=��Gp��!H P��=B:�� a�y�_d��T%W�=��`G�=�D�Q�Q�T}� �P!�E(G�P=�� }�S��Q}��E�T``W�W�POa���nT=�W�A}����D�@=�W�U}� �Q��DOeU�EC�=�C�Q9��(�G�\�dE��!T� S�A@�A:� e@N����w�[��oKm��n�l1	$�m��m��m��m�m��ۦ�o���o�>:I*r�|m�m���6ꔶ��:�m��)U,n[m��m�m���m�m��n�m6�m��ۺ��%$�6�|m�m���m��m��om�m��ݶ�*�T��e��o1��m�m���m��ۦ�m��m��e��m��m��r�o��6��ǒ�m���5-�b
I6�ۦܶ�o���m���n�m���[m�۪�i�ݶ�m��m��m��m�r�m��m��-�������m��n��m��m�-��o���2�m��7���ё���0�}{�j�np�}�ϸa�a��oVn.;�I�kW.v�n71�?}ܻ�����9�w'�{t��Ħ�M�۔ng�G�5ͯ����i��{V��s�>����|��;s�rm�n �{9ܼ��F݀ݞ^���;x�gt�r`{�7۵���NL���s�w�v�����F���	�,LR�D�Ag�q��Д�09EVh�W��<)B(S>Kn��	�p&�
����\}	�g��︯/_}�����4��|�R�ǾT��CHE Wى��Qi�E�>"�w��~���߮~׷o7,�WM���g�lJ�ɞ_�>�q���>��7n��>����}����3ߟ��ўVFa�&$�����Q	k��f��dWI���!F9=W��M+Dӄ)T��EZqs1*:�`a����і�Ғe�N: �Cƈ:��G'jl�ָ���Ű�Ra��G@pGV�4����vw@�E�]R�v����&�� Q=S���I�%sG)#/a�r�q��O.�i��]���޵�(��Ac8F�uՉh�5]u�����B���DZ%s�Wn{�U�O��8�<<��"�,5 h0��%�	I��0��[�;�vm�����Ǻ���^��݂4L�ӌ��jLK7a�E�碹Yċah�K$��֮"�;q|������w{wc�����uSUH������j����*��K+��5�=����|�T������`K%=��5F���q�Vqԓ����� )9a8�|s���s�pm�N7�&:MtX�2�0�3;��Č$ާa��f�[�,3�p�I C�1"��2�$ęY`� ti�k�bAl�F%��$�с�hf]E���T⑛�ۻ���﷭s�e(p�$@���E�pDNLc7�vt��v�&:6rlဈ�g�����딌-�u��S4PBh(Y0�筑�%Nh�6�k8�0"4F;�^puS�Q��f�5ifH�H!��HК3V:7��4�a��2��K4P�4��q�i���g�;����1��)�,�,N!�8�ٯ�o\LXkf���*
� �<����92X��A��z�[%��l"8�9��ڵ���K�l�PH�&�X�A�yރ�f1�M�wc{s�����?�˼���϶�4l �8<X�#DI!��4XN-%N�4a�A�����ѳ�3�1c	&s@F,$�TLXl�3Z����SD0U�jf�����Y;b4ml��y�����n�㞷�����i]�5f�+�y�`F:�0Ɗ�����M΍��l3F�4w�oZ֓��ċ9��96A'��8c�#4aa�8�`F�0�s���#���3C��îG�{�%)�\FDB�J�n ��p-Vbd5I�)����8��jWE��Se )!1��j)o����z	�1 �pѴ�2H�B�2e�4��b(�L����$8@�T�+&˭Ni�K�����3FUh��RYD�j��0&b����>F�g'��YL����
NkX�̨0"���k#Jt1�8#�0���λl�T�L��:N�;0��_�B\'# �|��u�������^�x�;x%;�q���Ǿ�¦E$�i�M�ȃs��Uܢj�%ȇ�vh�92+A��tOY��3A�1����a�e�ka�<<Č8,�p��i',7K��0MD�&&�Ji�A	� �D�r!��à` ���:�w�G�"P��t� ��Z^���ι+�f�f�]N�e<b%14l$����I� ���,M��%�y�Q&;����E'a�E���D��..-�0r�H���R��}��x�#4V��K�"	�9y;.7R���DV֤[t���k&�ޮ�D�k����)K�4���W�� Ѳp�6�0�5��6�'�M�q�lߙ֣�48Gy�y����;��_�~v��tNi��9zSRĒ��S�aѧ� �K�:;;Þ�ל��y��!B�:�q��5qD��6�u�;�Y̖�2SF�#N��$�0-�1���kC
P� D$��R�R4P�BSR� �y�M�L��8�-�t����kk-�f��&9Dˆ̮O�X�ʵ��q�g�@���rxA&ãf��i{�׾;<{�����{wo{}�vʌ��!�!�&C(�WÄ,�9�+��Ff�d�eA�1ԣw�&:g0*�$l��H�k-	�o�)Z�-v R)�BN#
�,�HN�/OiAlC5��sw�D�4:��g4�����������5$ҕh8�MT�� H3�œ���WI
U(&
b�&�*�\��K��w�cJ���c�ó]�����Cbt�%�$�/]o�25����:��F���P�y�:��brt���pro�H�R�p�MƒĜ�X�h�d!��$����"�P�q�����fd�����"Y�#q,��g^i��P����X�#C|t:���L���ͽbA�v��ٜF:r�#|,1�a��u����<c	YfH���g&�i��vq<��q2pI9*
	�è�SY��4X,Ն���{��ьaF$cCT@�$a#�0�  �"h�QprN,N1�@h:ULњ�f�d�|��ʴ��B(n_#��%
`R�$�43.I&J3i�!|AM�Q3k\�'�3�;�m�{��{��9�������{A�fV��pf��.xe�4p��
�g�^r�؋�6��SDS��.a&�'(&t�#��A�ᔢ�#�qM!�p4n�N�f��c��Z޹�\�l9��3�;�6�\d� 7ϙ��3[�7�'9�����ݏown��_n��ߎ��M�S��,:�ycDki����|7���f��#'61$D:9O{�u|��q���n���9��t]�pO M��4���Y�a�\W1�F�3�$�3�3XF`XaaP�iͪ�!�Xf^Ojڱ@�"20&r�,2��h��6�RDL�qLbS�]�\[�z�NkDwh�ќ�6s������Ġۻ��׃qw��};�[<{��ێNØ0���Q���%�YƮy냞fz�#�5��a�j������4Sk ��7�3�c:L�ʩ� �1"4	�kyd��#��h�"��I!�
0��DA�fY{�~q��V�߽!(��|�5�P?�5o=��1�=7��t~Fۏn��]yU������|-�oWva���2�=��pk�$���d� ��ЍcvQ�;z�ǿW�)��/��BX-3ZX~*���	n��X�_�}}��<G�7}�͏�Z��ߡ�߽F:v�?X�����r_g���N'�}�\���y���m��n�|~����6�dۿ�^�}ݷ~Im�<
����{{|}ȶ5�!�/�z����>�/������;�����\ǘ	�ogm��G���Hvw=���}�5O�TM�CJG��� hj��\X���0�a���g�����X��ފ����w���]�;�}��� m�      �      8      � ������0      �!�                                                                             �=                                                                             �@                                    ���f�ԭ4�6[��&�$ �Vʶ�H���|�V[�R���.D�Fձ [y���Wf�1˝��Nԫ*�� T��M���GV�m�%��A��5��� �ݧ(H 6���}�ʻ}��.��F�����[���U��!@Un��:^9˷UW]x�y�C�m��l8�[̛'NDr�#$�8K5�Yd�JY�����:�8�"�(jAËimԆ�ڶ�d� -��� H4\�$�B���6���d��+���6P�PA�1��{6�N���m��9i`��-���   m����P@e�`�@U�T�P�㊪Ѫ�l�ԫ�O6��P�-(� �5S��ۈڻ/S-`ԴR���u��<��۟���|$}����K[l`ڣ���^��K�
p�i/V�k�\�J���h06��b�-�.�k�Yt[�(�P���-U���U�f�q�K�j��Ӎ�C��wM�@^5�o&�UG��ӷ�ڧ�lF�ݝF�T<s��(p����b]��n�RZ��;f���$��7&�䁷*��F���R��I�M��j \t��*�\�P�[qtؓ K�r�����m�Hm�E8n��m���-��"q%�u��[���k]I�ź�R�����Ԭu(�ћnh�	f���lejX*�x�m��"r��m�h��-��Kh%�	 �^���v�%��i6�ˑ�̚]�$[]6��j۩B۷l	-�9t��,;d ���8 H�W�P�%�jU�M�^U� �I���`�@�m����%mf��)zc	�I�I�6��)YV�P%�����o��Ƕ�v�8�����M����`�ٖ��2�oh��f봓s�H�/U�Riz��+��Ét[��J�ᅺ�b����ygI[a!�n�wd ��JyC��kY���k���e�lհ ��h3��m-��-��ū�tm�m�e6��m��\&���l�  Zo0��Te@���Wfc
��M�$��l[R 8�ݗk&���ވ�ȥZUIi�O<˴�[��$��۶�9#�UpוUk��۰lJ�k��!�9z�v���ͺ77�]||c�l}5������������UH�ڢ���!�n��ڶlӔl��6�i;e�-�ɹֻD���` �4_�L�K.���HHH=i��l���tY$�� ���NN�p��n��Mu[�H�M�[ԶD:e�*��=iW��KT�Βl�ۂ�[�3v��e�z�d��;���)Qg��thr�HaM]�8�Tۭ�{"u-�����Ā#)�{e^kez	�Umr�)�m��!--��knnt[\l�۬����s���ҭ�m��Ɛ�����A��5�	d�I����]  [`�[�n�n��Jnm�%�	����mlp-�86ۛi5�����p��p�bt�-��ˈ-�c� �j�ݲɳ&�l�0�kV�l��Y!�R�ޮ[%Ӷ�6k�H�$ n�f��`��m��ʹ�6�j�C�+�P�~�횪���'�W�n�۟|�7�}��u����s��o����;�wn���Oyg��6��E��)vZ �km�d� �I݀'[F���o[n�Ze�/[�6�x�t�7��-� �K�0c�$[R-�Ӵ.�`6Zm�.H� $���Khm�gl���4Y��@�d�mm���m��	 -�fP��i+���� _*�» �a%����i,P۶�!� i��ܺܶ��m��i $u��䲁i���V�6ۍ�[v��+�F����傺Wv�
`�f�Z�S�W��(��t*^2m�*K��A�� <��yj��R���t�'i� ���i�S�礜a	�[\6�7H�e�mi�n��5^�����Ex֕�YUv@`�)P]/MV� '�o\�t��e��nx$2ޭo4��Ďz	$�Y:��s�-��InF�m��m���I$��R�޶����
�N�朧-��h�Lխ� ��:�.� ���[�m�@v�y��gE��۞���7tI���㗭G-�Mmʲ�UP�ݮڳkn�l۶��Fc��]��6��`�p5�#Em����d^���m�6��ku�p 	  ֛p-��Z����Zd�q�K����䕰 6�[%X�nZy�k����[���'2M�ݶΐmq��F�pxh��m��9�gfR�J�Waڸ�>��[m��$-�|�[+�I'@�U�ڦʠ<�դZUU�e��]�ڸ.�LB�PpH�H�ĵ[i.�y�̋.���t����I�jTn�t���f�^�OWl/�6�Ԏ�!�ܶ�,v�������rZx�@�^ԓ�uܷ�a���6���2;����HM�/Z�f3��	-�aQud��YPD��5�9`۶��������qԺ���y�k�$	 m�� m� �k�-��uWJKu����� �mm� N� [M��}�}��	�H@[F�lm�v�m��   8�l�L۶y-�
Q����v�
�iem���ٖ� km�m�lp�`�g$Ít�m� ��-�H[ԝ6�m�8�h 4���\[B@ ��΁�uWS��q�&�O��)�q X[p�X`ڶ  �l�~U}@Y�L:�p�R�*����K��8p�\R�n�ET�˲��.`�,��0��/��^y\ɡm��=�K�{(�x:@כ.�.55���M,a��hic mz��m6�ܑ"t���mH �[���d�H�mr� �e��m�A�6�mgY������q���;��{���Wk��'Vs�C�����ɷ�E 6�k3[A��6�c�V�n�D�p���G9m��h ��m���c 6�-�	 k5�$I�[M� m�Ͷ $�m�6�մ:ۭ`  mٵ�,Sj�t� �m�� ɶ�Kd�I    �ŝ�ͻ ��v�
�D���-���];��\�^��m�f���l����H�`z�[E*�d
-�U�`*�Zku�K$*��tͰ � ��BI�j�]l-�-����-h   l/Z  Hm�Fݴ�lm�h-��l l���6E쵮��U��    6ݸ�M6������yύ����6�qۮ;�=��=ߘ��'97��E=�sf��S0 տm���yU�'hȵUUՔ`-���mf�52��f8���Ѯf�n�6襴H jK.�u�hke�Ҽ�Qk<��ʵ'de[��* 6Cl��*j�
�Sg\2�;�524��Ԅ��T�^6�a=�����۴w�M���n�-��;���Nꪫ�Uv6�;M��O�^�� m�,��)�[o[�m���?-��Mfu��C��kI�1�����T���U�:F�U�mmÓk�� V�m�9�d��  �����k��-��M���f�o[����_Ҁ� �!���AQ��  ��~"��9�SO�b0�U�fPeDQ4d�QD�Qu�U�Zs(�+��ʔ�-h��4 "�"�@� ���  �0\  `� � ��TDUEEEE$EEEEEU4QUUDTDTDTDDDDDDDDD�EDDDDDDDDDDDDDDDUDUDUEEUQQQQL4D4D4D4D4DUU%ECDCDCDCDIDR�TQ�TQTQ�}�6���~c����C`}�xj���۹�4o���Њ#���"��(���<�.�����;u�H�(x'xQ�j
>!����C��Ní<�)���c��s��b`+"�2	"�
t!�lTM>G��@�D6�( ���z�t���(�	�1�
iP�'�}ȏ���X
	��I��H�� ���VS��<LQ�8� s�Pw�N�M��+�ۭ"Hr)�*��"$�(�9� �="��y�At��b� �r����AH�	�^���Ñw��b���"ʺOz��tr�H�ׂ�
��b��@:P|�(�x��"��B���	B� t�>*/*rn:G��^{-f�л9rш!�P9�95"D�8�T]�x`$и.��<5ښA6 �w�� =�C�U	�K�gJ��%� �L��;HDw�{���Ό֞U�^U�^�^U�^U�^E�^C�yW�yW�yW�y\��ʼ�ʼ�ʼ�ʼ��^�^U�^U�vݷm��h��(��(��kZ(��(��(�Z֊kZ5�h�?tAT(P!@����{���wwUV˻��D�RG$�J�u�݋�9$�K��|��@}y��9 �� 29�8����@1 �� �q��96F	7��)�e���x���k	�f��ʅ��g���n���1��{�W{2�P��*.C�������$��~�x"��t>�9곂�g�e0���!+�|*Em�Tw��˷VV+^�_����ϝ�~��	A  �G6 �`              �               �`      �K*�s���њh�]ONj��6����d[�;�0p=�q��e��l�d������m	5Ra�l��n=�B�E&�t�I����eyR�<J4�5�%�~�}��6�7���G#q]�Fv�M������M�j���;�vmi�~GV{a\���m�٦��[�$�C��U��*�l�e�A��}��j~��mߖ�����}��1����I[�LGY��6�g,��QX������6���� �RtS)��ic]�A�=��{����5�m�����;��͑~^gp���LX�(��l���.�\�*!dݸ����us��8�z�6t���j٭���}}}$uQ��^v&y|�Z�vN'��?R2}`[�m$`B2S�Y��������2��hsUK�p�紂jG�X�f�G9���i:�d�"v�czZ��5�l��sd������HzzmۧT0�]�y݅��λLa�w`�� ��Nc~aP���ӡ[�]i^��ʵ�L����6�3��b�Mu���.'�3ͻqͲe!�km��Q]:9<ɒ��/T�������cu�p�Pٗ���;\ᜧ���_�~�Ju�^v�Ljy/0Q�Z	�A��ݮ���aT9���n�ɑ�9��6�=�4���W2kNK,y�u�n���1|!�vĿϹ~��������.e�T�,",]:m�a�+U_�����[)?~
O1�6�$��K�Ѭ�4���4�5騗�Q�ؐym��m�[v�M�����s�趩yWh��3�e�h��Ԛ(�kLv��m�ۿW���j�Ct�/a�y�}�������-#��m*�Q�/NE��Vd�����ƞ²�!�h*�u!�.[�#!@�%�ӬrX��l��+λ7���D�;@L 8���9 ;лU�Q<S�@�Dz����0��eB�yx~9~�~%�N
�^��]�  m�  m�^"%Ĳ�SE�*�`\�OKzn0#���Rr;i���8��!��봲���������["P콨)���������?'���j���}�o�x�c?����6젴\�ƈ��#�vu������.��m[d�4�'W[W��o�<�!Cy�wޞ4�dsp� ���?���e�����y�w���|���;��.<�eN\+�s�p9rg˹��"(/���_]����y�w����;R/��j�����?&�!$�EՀ77��(����ޕv@��L9��Y($]&�N4}�d��j����r���s*5:��"I��6TNb0�� }�whA��s3H*�lLm5`w������#��v;�j�3T�km���1�G�Jۢ[I=�����swT.�[��һ�XvI� �Ad�,� �� �mՁCwK��y�H�� �i��p�nʟ�|=���K��O=�欻ӹP���+=�@ �'4��T�)Ӛ�bnm�@w��>��u㭻$����a��)m�i��TKu �~�tY��Cۻ 	+ܽ�Sp�j���k�-���{��������u���;߮���UUCꗳ@a�5v��c94G:��<Yl���$+���ߛ���݈9�zX���N݁��<�APa[�a�bz%���b���%��ݻBA��s.��m�[�;�i�|�]���1)(*q���jj�� }~Ǣ /wj4.�*p����܈�wU��zX���v����St�N��۰7q�`w��
���,D%�뙯6�m�c��)���\���>(ݮX�A��V����w��A�zz&�9t� ��֭��L���L��ݐ �nR�L&�iSTKu`
�k�xH9�{� w6T aß��Qi6B�v��d�o���������P݌�d�Y���$�	2�a�ۻ%�ӱd�����4E�@����#|���s��ju.QANI)� �m�@o3*Ձyܻ��v �b�F�ڪ��ϙ����ݧ�01�y���Ώg\�uG.6T�� �6�P�8�g�OCݲu}f�7�@vuB�i|.���f��P�{� ���ʀPØ\$G�$�&�@�� ��(��P��,��z�iM2��A:e�7'b P�׽I��t,��b�'�[� <w)m&M4��[� ��� ��;�h�}������\8�*�@�B�L��H!)� �ǻ�w��v��}��s����~\q�*       .˗5��N�m1fg��i)7Oa��Daۤ�Ѷ�v��ܯ=�N�Ue�&�U{&�u�]g�- �gN5�w@�C]^-�m�]l�;/<t/$���9-$/g=��mX�}]��u8<�����Y2��ƍ�t�t�yxț��]��~�������ʪ�m�;|�����n�q�F�6b���I��5��iIz�v��r�_s|D�M�IT��i@&/3# Ffg�D%�d���,�ŭ.j����]��[@�D@�Ƿ#l�F3;�!a	.�*<�LTT���J#wۈQӻ1
$���8��F4�;�͙�AT�(ݥ�	i��Q��!E�1�H���z�!Gwu9���R��JQ��T@fI�6!��b I���0=���߿���~��UQ0c����D�IGD�)5�,�$��1zR4�J����a~��߮�����w�3�Fgq@��3ܚlt'*��t�Dfw6�O����%%2�#Ky�Y��{�|���P0�F�u�d� � q��*UM��UN�B�م��Dgfwu�"-�w#N�HY57)*� z@ ��uD�x�G���=rG{��(���HR5*�Dx�`�׷��zR�ė{]iB��MHV6�m���x��:�=Om�[vW��{���f7�\g�����lґ4�@D�;8` O\��3��swG
H���34��M�L�w��\� Gd=�#�֠Dkx���h&QTKR50�3;�X(]�c��"2fݼ��ۖK9�ˈӎbL�Oj���*�ԙ�G:�!���pݘP��IOz�J�=ɦ�BeZ3n�{C�μߜ/p���{�}n������Fpm$�H�E�`�{m�K��Ў��vdԄ�ơݾ�~����m]�T�5K�:z�DG{Ψ���!���J:vt�ʝ�MU�l���n����< 1 c�(��b � p�� h��d�SU&�)I�. CoP�v",���Fgq}�C�$*���J#3sn!G�J#3�p�X�	�1QZ�F���Fwsd�T����J���n`�cw��ր���ww�����~�R,��u�a%�*^J�u�n������������;ww��ݿ��Q9̜@Dg;D�rG{�ʪ�.AJjL�X�h�׷#��"39� {3ܚH�!H�)��� GsDFg1D�<P"8��b�T۩�Jj�j��0��!fw�(����bN� GA��Vd�U�J���ߛQ����H�߽��/7�`/��߿����O?u�__V�       ]�VZT�u�r��kf�m䈓�-+�;s�`��7�y��t�oc���Y1��ԯ
��;;��%t˼�- ^a(X�E��g�0<p(!VN���fts� �@峌����q�� ;�;y��m��m�[%�:M5UM79��m�
�3�����������_ *q�\S��v�1�����byǌu�7'�{}ӏ�3sV�*j�҂��q:�@Df<w#���.�q��2"�*12�S�PH�Ǎ\@���t�@�Ā&"y=Ɉ_D&(��$�"�M��p�t�'r@���P�p"f�@D7�l��:�jfj�M9(&jb�!n�B�$������������ک�9 �Jj��\� �h@�׷$�N��޸�c�u�m��*jJu5R6�^��Ңk�ۜG:MmCvv�n�m�B���O_z>��ǎ���n`Dfp���,�#3t(� F�ʍ���M*T����n@9��T|W�v�D�λ�	̾y����6� GOe�t%s&j��SR#H�q�#��P"35��8[�";y#�p*��H��\@���Fcn���nD@��f!��E�ThE("ii "35��`}u���q�9�by u׺�S$C�Ͽ��y����y�qssh�%V(״¼��r�\ùu�;
чg=]��_�{�����Fgz���(��0!��ɡR&�$�ԁ�b l�d�t��ou�=s4� ���UM	r��������ˁq�,DY����ý��䒻�7~�����g��z{���������;����x��s����{]��| B@ �Q1H�AM4��E�0(��*2Ċ��&
"�����()��3��v�G\mCI�f�5����H��`�s�= �����4	dᤝ8�AgMC�kA�Zk\�il[�0�n�b��;���@2#,������P,�s�4"Fo�IH=2�@lx��� '���am��ٮ��0�$pM��#�i4Q�q���:5f�����P"hyW�� �CG��H |��:S��P�NA:M"q���5� P�Q K���	C�zP�Q?~u��^y�����_s�;2횑?�ݙ�ޞ(�j�@dk�@N`$A�yq$!H"9�9�Lj]	���f��-^y���S�d={��#Hy�}��9��`w�OU�qd@$�����6ʧ<��O|rs�%!׾�7�C@O�w�gM!T']{��*2������}���$�
i��o���o{��9cR�,��n�L�D_z�u�ۉ�G�f�_����Z5�����9��(�BP�%"P�$BP�%	BR�P�%	BD%	JP��ϟ=�(J��"��(J��(J��J��(J�
��;��88��(J��(J��J��(J��(J!(J��|���ʔ%	BP�	BR�%	H4%	BR�	M-	BP�%	BP�'^��bP4%	Bu��	BP�1	BP��	BP�BP�	BP�%	�y�yxoZі�n���"R�%	BD%	BP�%	BP�%	�%	BP�%	JRw&Bg~�����	BP�%=@	BP�	BP��	BP�%	BD%)BP�'���y�H��(J!(J��(J��(H��(J�����(J�}�[��(�(J��(J%(J��(J��(H��(J��;�(J��"��(J��	BP��	�%#BP�%	BP�%ߞi����0ַ����)BP�%	BP�%	BD%	BP��	BP�%	�%)@о����y��(J!)J��(JR��(H��(J��(J��:�ݛ��(J��(JR��J�P�%	BP�%	BD%	BP�'�y�	BP�%	��	BP�f)BR�%	�%	BP�%	JP�'={�D�	BP�%	BP��BP�%	BP��	BP�	
(@������@��e3W|�JP�%)��)BR�%	BR�$BR�%	BR�%	BP�{�͉BP�%	BR�%)BD%	BP�%	BP��	��	BR�u�|p%	BP�$BR�%	BD%	BP�$BP�%	JR�%	BP�u�	BP��	BP�%	JD%	BP�%)BP���H�/�8�zCG�Ϝ��P��	BR�\q��<�BR�%	BP�%	BД%	BD%	JP�%	BP�%Bu��fk-a���+�����(JR��(J��(J��(J��(JR��)S�=���(J��(J��)J��(J��))(J�� :��v ��|��}� �~����������o��<%K�2T�/bɮ_]�t�����ۢ\h���چ����%	BR��	BP�%)BP�%	BR�%	BP�%	JP�'}��	BP��	BP�%	BR�%	BP�%	JP�%	JP�%�~��<�BP�%	BP�%	BP�%	BR�%	BP�%)BP�%)׾�bP�%��(J��)J��(JR��(c!(J��hL��8�J��(J��(H��(JR��(J��)J��)Jz�g}4��C)5c��P�B PP�%	BP��	BP�%/3��%	BP�%)BR>w��y�J��(J���J��(J��(J��(J����3�m�H��(J��(J��(JR��(J��(J��(Jμ��(J��(J��(J��(J��(J��(J��|�(J��(J���������)J��(��(J��:��s�z����z���z��%	JP�%	BR�%	BP�%	BR�%	BP�%	BP�'~���BP��	BP�%	BP�%	BR�%	BR�%	BP�%)�^w�R�%	BP�%	BR�%	IIBP��	BR�%	B%	BR���	BP�%	�`�%	JP�%	BR�%	BP�%)BP�%	Jg~���)IJP�%	BP�%	H�%	BP�%	BP��	BP�%)Bw�緦���5�������(J��(J��(JR��(��(JR��(B���|�(J��)J��(J��(J��(J����(��<�(J��3�u	BP�%	BP�!BP�%	BP�%	JP�%	�~��<�BP�%	BP�%	BR�%	BP�%	BP�)J��(N���%*Д�	BP�%	BD%	BP�%	BP�%	BR�%	Bsߝ�<7��Zݻ[��"P�%	BP�%	BP�%	BP�%
%	BP�%	BR�'}��	BP�%	BP�%	BP�%	BP�%	BP�%)BP�%)�^��<�BP�%(Д%	BP�%	BP�%	JP�%	BP�%	Bu�ؔ%	BP�$BP�%	BP�%	BP�%	H%	BP��	�^w�P�%	JP�%	BP�%	BP�%	BP�%	BP��	B}#ҧG��C0�4��cH`�Hs��ެ��ی��f�yћـ       �E�Z�"+�W[b楷7,u�HD����s9���b�griGX��s�7=�Z��Mh��U���E�`���^�n;k2��3�=�]�鲅䮪�,���nu����nS6<���n�u�ه�jݹc9΄Yy�M�Μ�+�h��ڴ%�w=�;���UTW�r\�e��[�������]^��]v�c<u��Ѿ<�>��ڵ�n��t%	BP�%	BP�%	�%	BP�	BP�<��%	BP��>��|�%	BP�$K	�^��^9����;�h��{&jH�	:&j����BnP�;ڏ]{�ǉO%"�n{�|]%$G���MIR����Zׅ�5לy���y�~,��������	%�}IDYk���*M�S"n��3K� F ����������0 � yX�Dsfq�$UQ��UH��wyC�
�O>ZaK�|ڏ��h���~������*���^	��4��$��]��O5ͫvq�ݵ���UMIo���_����������|����pu�O��72���}�!�>���2f�J�@Dn� |�}�b{��Х�Z�������~�/��ȁݨ��nFEI5SR�Lҕ`� 7�!� q�� �B��P�Ȉ�f5��.��ZcpQN����9:�x"�� �@;�>B�����"!d�l��*��HL�w�D�@���)#3�q36�!���~�g���_����v��D�Zړ���ޭk�����6�P&N؃W������������G���j�!����C�9�:��$G{���r*hʚ�3W#�րف���4��Df�@D���Dl�9���B�QRR� ��y���3v�p�f�#�!�[@`� Woػ�"�v�@���@Dw���RJ��T�J���C�d:���O�qw��j=��ݪ#����\��9�3LRMS�����^w�y�c�)^�{� �PaꨁǢ �#kRI$��*�stb)G��s��nҋ֮H㍘��ڣ\��|��|�
B�R�V�b7� "u��D;�PP����w.!G3*<�7�ۦ��K�|��@�'B8�O3�=��5�!G9�8������fhRl���`Dwv��\Ψ���$D<�q8ܷ3RQ*����D%�#��j!X���@D_u���" �p  |#��?���q��y�Ё���4&��ԃ5`Dfn�;�w�#�wv���^(0����w�������E��N��ᶒ��N��z�NV��v�nPa�N�o%{�7v������� GwjE�:�s�� ��T���U +��+��0;�P"9׊"=�,�׻\�z@b�ۙ�FL�FUJ#�#��@ ׻ȁݨ�� 1��]f���
�X8@������Gݠ";׈��zA�I�A���J��ݽ�@��A�9����5�=�/�<���H�on��v?�s�����>-��j�      ���m��r�9��^���D[���{"��<��n�gذP]ɡu1N�vw5�Rl��n;m�/-4��Ҝ<��=���۞��Q�G�{�n{��O�ʝ!E����,��GFMz睲VrfG���7:��vӅ�kBU�Y�vښ.�fD��D.��/\G9��m�I���@��GK۷�����7��b�����om�t�Ƙ��<�g���`@�N�"9׎���[P?D �dD��}������ԔJ�a K"#���w`{n� nV�t��o�`"":C!�}��	Jpu�gz�E�[�aY�{��v��2y��:��/�'\�4�X��wI�R�h�*%��D�DD��؀4��B��@�� �aC0guΪIPT�����W�8`u�i��;�z��6�@��]�ＢW�|��~ .N^�v�d�]2f�X|]<ͦ�V�L�S
rl6113�����w�����~�:��=�`��y���9����(���C�����)U`C ����Fp��_�\CR�K�ӌ�������ǭxuk뿯8��6�H�� f6�@�=�D�I$��}{��#�	1��`��Ǌ!G{�iDw3�$�
�l��f���$ Gwj� �^X�s5(L� b<���D%��|�jJ���Sj�Bk� Y�dC��p�13��� Gwj�#��r���n[r�6�!A.V��n�m�ݝ�g��^t�ӱ�������nݨ,&�����}����߻��P=��=�/���\B�zsYNe�7#�2�J4H]����A>u��£�>is��lf";�5� y�uRJ��T�qJW��C�N�֐74�^w��H��0
���Hz �α�<����o�D�w=�B\�#�zI�I5N]K��^w]�Y��e0������0 �҉���	o7)C&�����B���@fu��p���� \��� y�w���S��<��I��T�\��a����s�)=����Q3.S5-6�Qb��%�������wuȀFf��� 1i���ķ��I4��6PL�j�	wޤ�B�^\� asR!�ww�H���3RhȪ(L�*�@f%�h'R}"��ϟ9�ʏ>h�y�;�h��!U7SK� �2}�����@��оH�_� �W������\<�b/���K�RS(*��*L� 	׾����<����B�]�� ��C ��G����I#!]:@'Y.��ؚyڽ�l���h1�gGb�v�p�sN�Ni�/�sW}J���P�;��
HN�:��6�H�Ͼ��"�K��{�Y�d�R�R���ր�� �j �A	HϾ��D(�Q
ȍ! �ݤr�H��5˴� ��!����b wv��\Π @̘�$T�jRIJ�G �{��߽* �0s��0 �Ȃ�����&�5A#G�5J�BQ�v}�	&$����q���s��
,���ׅ}_�3�k���݋�i+��Wv���������ػ��wv��b������]u������]Ȇg:1:9�\��B�6�����J�K�@}��g����=8�D�	K��'e�\�"#Y�EN�H�'R��;�A�uܕ��h��.s����`��Hh��A�2��T�L�h�bB	�����&�:.�{"!��$JT&�V-��13�<��a�T��^P�(`���I�z:�����美�����"8h%����&��&���<��"M�����D�I#7�*�T�pҞ�%��k�p�)زI��J��Շ��wl�B�?xܣ��Ѵ�����^��r�_�-�� H$ 8[%                                        ΍e"2]v��H�Yn.�X�8���z�����m�y;��)�jƵ�T˭V�#KlNݚd���Pkz���nx�&AQW����êiY�i��T���9�L��Q�}�۳w�����r6)����BS��� �ͲY�(�&�;uY�b�.Wr�#%`Ѹ��,������n��k�W'm�����:lm�w!m�7 ����p<�II7U�YV�]l��t�W��c��}����[�K`s$����8���56�2�6��j֛�I�3vB��=��p��a�n�dԛ'om�![/E�;��:�ن6�+�w Kp�sqHM�6Uc -I�'����Ƈ�+�J�Zv!0�ʹ���q�-��m���%�In��m�6��ظ_�︇����^�F�\���mؐۊN�us�9�ݮ)���Ĺ�H$���1�*��%��?���yG��h|��Bi�PvnM�f^;9�);��vӌieK�q3�y�]
�E��K��G��N���^�U��k�\Id��Y��E���H-���d�;!��R-]�nXp<͐�+��}Q�f�X67$��"�Rҵ�n��E��r�6ӱxC�ş8i�.��m�^���b�t��w�o��� 89�º��^�&�K����EȚ�U�T�\[
���rh�F���e�$��5J�m��m��n��[X����͑.iX拵,���Ѣ/M؋��q�[v��)q����T�AX��}�l��ŗH[Z�1��I�����w��ϻ����ȟ�W���M�*iM�ON{G^��x"�~ ���Z���\�����~^�}��wv�       	�,�нmoK��h88�v����~��\�ԯ=���v���T룖���6��\���ݟ�=7�;,t�W]T�ܩ���7�.�{%m��(��c�����}�����0�ulu�q��0�w1��0��IES���v5n���UxW�n�	�m��:�`3?���<1-���������ۂt`�ɓi�i7�{-�[�v�Iݻ3�<oo��|��9��s5%��� u
#��j~ý�`�{���	���^�K���U�ȴiUL��!�ǦP��`Du��"B�=�K�B�
/�Z꜎&9����{�(����	��qi��P�o�i�I6�A�N}��ܫEz�O{�U��w]�y�Z�~!0AI����N��~7���E������9�1��I%(����[��j�ƻ^�9���u�n{r&��{N��T�T*�f44����s��o�C������=�EJ�e*���u�����@�� �D��ͯr1�Q��s3,w��$I��UBT�(&i�\���}�S�vJ��of��ws%�T� ��-��Z_=��|�{����F<UUS��9�BJ����^f���Έ2��b�����v.�6����в�Q�v�+��-uˣ��m�[i:hSJ�D�[�B��;���q�X}w� �����Fg�>UIR4U �JV7�ZlÖ��̦��m퓟���I�d�R�J�ou�����~?z5v@���JX>���;�d|zۦf�F�Q�W'� ��}c��{}���g/)cH^Lf�*T�5)$�ԇ���,�yޮ��+����w���UT]z��7J���"��M����,��j�ܷ�!�n�z�8���o��4k��w�h��y�w�wuLԚ2&��2h���ƙ�{^���o]�u]�b)TL�AR��Z>�n��܀�7ێ�|vq���%3Je n���ז}#�;>��CL x� }D�z�<A�w��*��R% ��\���C��33Tgu���0މI$�T�YT�m���ۡ5ݢ+@	���!���sr��S���(���d݌K���\�c�Ϸm��Y�;�X��#"��ѥ^���_������O�g3��ݦ�D�I$�wL�_�}!�(Y��w���/l�H�U,r��\�rr���n�ws;���n���2&�
4I�0�q3�������|�쌪�(;=�����s�{[@      �tX�[y�G�m�6ë'�l�]�$�b5m�N����r����h�&�>�.e����ءْ֨ʝ�ۯd�e֫��]����g��-����Du���X�ԋ���H�i&d�F�7F�k���[v�I����퍹܎6���x]��uj;u�����������{��UZz�+��W7��Κ�,�{2GK��d:v��D#@��-|L�I[_�p��ٛ�+:�y]�\�;.��	�R4L����z9�
��~�@�y�s�Xc{�l�R�P��JR�whǙv{�Ң�^���q�ɤd�R�FP&A��u7vAy��h��&�H��UDҫ�C�{����ᷣ���?���l��I2AT�ԑ��y%�f�v�$�m��瞎�9Wn�9R������W���g�{����qPe��4��7hg�� p�y��71�8������ǎ��� ���3RhȚRd��|I�{P�[Q��;n���s�*���%E�.�<JwY�͊�oo]��_V^���e
B���A�d%��c� ��/���fO�I$��B�2���.��%%��c��zJ��j������?�}����'��|��f� ��C���{�;�3��f�	�UJ�J���S�u޶�G_������tRg�e��3�!W��?�����;�}�7�/jz�Z��� 럯4w��a�"��jRI � ����v��ch��7��y���f�%%�IX�� �u��Zdu��CwP�WU�%�l�j�:�^��㔶�]q-�:���H���D$U"� ��3ݮ���Eo�{���UK�|�8�[)P)J�������u��Gq�,��cU
AH�h�K�!��J��U~�?�����ͶKiQn�UJx=�(��=��F�Ԉ �$ :@��pO��3�|/����F�JUR��=������;�w���9�@�Zc_ u_!o4jI/d蛐��>�69��.=K���tRf�TYI������~��{���C��cR�5)$�gnޞ����,x���3w� U �M"Xi��2���M�9Q�{��5{�%g�� ��آH}�㫼��{7��s����>H�D��%5 �pfl�Q���x:�#��C�(�	<Ĥ����nQ��M+� �       .���w�yh�m���Ӈ�#s��9Nd&�:�N�'l*OO9�m�׿�︎�Ǝ�`ſ��g?v��m!,h�2O/����۷zk+M�����&m��%<h3Y��je�;��!��ޠxM�Թ�ƹxyf-�;/]��&���k�^���~F��񪪎��{b�=�.+�Lk�+v�<㫙}�V��9+k��辟7^mY�R�=�,q����P�(�;�uU!(*�)�R��wP�
���7棹�;�;�u�iUR�*�רs����ߒ{]����3����(1E��z���K��-�;�v㞁�徯m�zb��S&��J�=�a����ܒ�5�j<��3�O��s��'GmKjk�v.6�j�e'������
9��KT�A4ԒS|_g�4���s��� q��'F�ٚ&���3$�]��������dH�\�>���)��  aFA�!dn���5(b%���=|�� \��@{���n�� �vr�e�"��ԃ5c3u"7��y� �� ��� ���便T��
)&R��~[���Y|�B�D@��h��k�UJPSFR	*J�35@� ���B����:��\�m�
 /�JH�L0�A�[��d=��j�B<��f��)��C��?ao��4�SR�ԸӾ���w���gߢ舁�;@pn�5*D�J��4lw�j��s��j�6� @�ø���*$&�e����Wgk�:e�ۻ�wm%wwv��ݶۻ�b������ݫ��wf����ٻ��w�5�$}^UA��hxy��h��	��B��.�2H�i��	13ĐhU�1�4�L�P��TPAIȜ<��ဝlN�Pٱ���	H!6A�
����`h��pb����BBB1q  � �#�M1b���λ�k�=�ÑO@�t(��(t�!���4**!��8@]p ���
� p=�8��ਾ�h�~���=��S�'v��\G���Z̈9� s9�"������cQ��)ɚ� L�J�wP;�$�x��F�Fh�2&�̒��k֙1 f7qo��wv�H�N���������x�����c^��WgE��[+D;-՛����D��;ru
aߟ�����A׻zs6���Q/Z����(QR��e(���2N����=�$�N�ݞ*�)ML���v��3h��ߢ D�~���eW��3��^ׄ�5(J�Q�.}��3:�~�{�c��"�@& x�����6jT���4iU����} <ox;������;��%��I%(�fh�J��M�[r�[�n�1�ٍ�ׇ�ؿ���ݜ��d$���^ﷃ����D����/q�&h)�HI�IGwh:�x�<�J}{����Fh�2&�̒�z�c����}Tovw���UW,� qI�$�+�C~�#��x��u;�Hs��HТ��L�rG2���< #_��q�����y�#�^�(/��8�D�H��k�3���3����8��|���^��m�       ��SZ�����n�a�e����]�����w'k��n�۬�m�ϯ�*��fҹ�eˉӈ͊���ǰ�jy����ޣ��`�E�q��x�B���tS���JZl���㰧@=��b��ճ�����Sn��Vx�cF�BPK�uv�.*��U����}�}�w���� ��UYkN���աt�4`��FAB����v ��4Z���ww��ꠡ�uK~���?�w���L��]��n�g���	)D�J�*J�{ڮ@��=mY�m���b �1��UjeD��R�gt���g}U_a��I��uv~̠�J���T�Ojսr��RK3��a%+=W����A4�s4RW����2��u�_[���2g��\N��l�ttqm���4^"]���^�P-ּ�I#4J
hJBfITo[޷�Ge�ꫯw*�{�P�R`�J�����_S��O�|LQ��0a��:C��@Z++�+��H�̥#�9J�4(�H�2���v8�Eh����8�;�wvu��6�鶛��}U�҈���~8M(-�v7���T���J�C�n�ɕ��c?^���,<�I$�JQ	<�"�]�$d�p�LNj;Z3s�����������T�R���\f��c��͈X�0��Se�e��+;j^�U_�uq��l�oN�4L�	*F���ځ�]���=>g0�a�J>�I��O�_]ۯ1g>�]���tI��k�v;��ovƁ��:h��3�FY��B��&i�w7T\@�7V�wv�w��/�߬|UU��8�d�	��E�v���I�-u˷e�B�K1D�T�.� �^w{�^���<@��[ԣs�>UJR��(-�J�;�P� 1��Z�fk��'hII*�U(���`�=" 3-�s�{�@q�&�Jd���J�X� �7y�����m�#�b�Q(D-;<�n�4��; ��P��������1J�&M$�(����� :��޴;�� ���p�l���Y66�^ֹLg]n�!θz�X���"!�Yd�J[t�o���-B���t4�{�7wQ��D�@̒�ǋ���s7Tf�xzꅽ�іy;TL��	&	 �W�� �V�w����u^�݀sg)�U5(�	I��� �/v��+P���뱇�7g��JUJ�T��wv����w�j9��V>�" G"@����!������P�d�������w�K���ڪ��     a�0�n�{C�a�q�X��[V8{4��<b�"���R���t&Ԇ풞^�T�����/\݁�G�5�A������\�n�ҝe��%����l@��N��f� mӼ[��]�kqÜ�ь�Q��u�����c���\����ǻ�ߟ��v��q�UUE���&��_`����V6��XFnv倗x��[�������|�u[����o�/����c���ɠґ!Q�J�X�g��@��^�{kk�m�K ZnY)T��E$��}{c������u�oN��BRJ��3JƁ��chs�q @�9���{�Fh�i
�%C{��:�Q�f�g��D{����7;A��It��[^=f����)Μ�ۮD#��ͤ�M�H �Cw��O�v�P��o]���ڥD�%���מy�>}|GŔ��$~p:D���~Ψ�|�8�0�>�UJT�J�5IX����O��֢���~t��DR�UJ�G ��|�zھK9N�68{�@p6� ��34iR��y�.����@���^��n�|br�I$��	U�@����F�6��M�&����݇h랃G��~��2pjIRB�[{c�h23C�֡�6�e�B�MJJ�T���� ��j�j9��z��3RML�4��*j:[ԅ�1�<�"�d�$��*3J�J�(��~�����]�U]��@� H�HV 5�۲/�����G� �6����R�T��%&R�|���|=+P�6�{�q�KD	f�m��nX�I.�ں>�v��3��A����u.y����xz�������|},R4<��.���QӒ�(�n),�[��^ׂH�T��)�{�� | D	���Q�����Q��r�)���*U|/7Tu���`D 'sh��s�4��*�L�IRA�� �������C�a@ E��d���������t��e*T�5K����4D@%����j�fg�\��6'���+*5��ӵ��;6�wa�rz�=XӃ]��ZD���5w3BjdH�&d�@s[e��6���� �8;�@fd��.�5T��2���Z� @��ge5f��3z�U�L�TiP��Re-���-��9  s5݌�j,�s��JT��W|k=�wt!�b �B�ec�	#J��!2�����T�\ƶ�vG�9_O�W�K�wvm#�����뺿���?��{����ٙY���{����wwwuwww��x������㙮s *�&"(
`�F+��ʊ#�2��,�"u�1j�"

b	����#$��F�~K������~o�Ү����É)	J�u�=o�4���R΃j���6��s�]t��jJV��{7��p ��.i2M@<�.�� yӁ�m��R�VR� 騽) �!�	�=y�o�As�ۢ�y:�R*:u���Mjb�4j閈l�I�V,Y�l�Y�RFOс)=�;f۾��m q��m�                                       gG�l���'�t��D�m��Z�\��Y�z�M�<.1[����)Y�':5A�H�e��k vI�mƽ)�[;:���J�-�t�KO%��Z��k�Z��n9��ޯ ����+n�������Q�4�׶+v���]f��#��T]"fw2��XD3�R���r����<�������gaր1<�4�//���\+�s���h�C�)�_!.�m;�/�Vق�yv5�d@��j*�œ]QsZդ�)�hۓ��.� Yfv\�'�F�/j�ٶ[H�V�+�"U����Bi�!�,hzݨ�[���=u��\��ER̪��[�]2�  �Y��v�m-�`�Y�����n�^�F�Ll�ol�rsɮ:3#σ���t'n�#�d&�\�G<��F� �3Y�K�$�����#���`@����Lēϝ
Nƚ#9�6�N K9�994�b��5��P�댣�-m���p�󈞶R�7C)���F�Z��t�:�	DE���e��w4JP[K�IuM&`m��ċ�'d��s`dV�`l�zI��i-G�ZvF�Lmsm���PTT�;E�t�:b���F��m�ڵ�<�$ׯV�gZm�b�Un�*��v�iZ�K�d�i��e�z[RM�RѢ�HZ�fꛫk�Cc�x�~b�ɛeM�OkL]�u��lgcҷ���<T���u�]�U����El�1��˪����m���}�������?" ��@�>`�ݿJ�G���*��u�@N�/ <�>'� �?�h�"�8bjzW��7��9k��}��>�ϫ���^ǻ�f       ];����L��1A`��i�Ș�:�k$���7g�)��JY���F�M��Z�	��^9��cV�;`��w}�Ǿߛ�O�4�㧓���w��7`6�l�0��P����>���yk	6��%�'^������������������e �d�m��q�����??.'i���g�wǯ���zO/\]%m�WG���[v^�_�>�n`7�|m�i6���{���j�	&�hV�;�� ff˳Į�R��Ggv�0��i����3=v7Z`{u�`w�۽��TR�~I4�t�3O�w=�V�,g��r��͐�;�X*�&�dU`��t����H�ސ�,{��2��D���4R  �k3�@n��t�����
���m�i�i�It��v��Q��n�mۃ]��Kq�'�����9���a�0n����i��X~҅��QY�������)�U%*���W|''7l!��Ȃ��hD�(����>��]lLDP�O;�'��ֳ��o���}�d��݂O���ZF�)�D� ����>>��?}�#��Id�o:`;��RS&�S�
6O�+3��$���'kF�}�ar��F���:�K��n�2eg��^���Z�7kF9���y���s��D��eY��Bk��n��k���^���s�h�]&��)M1O�w�i��Y�c	�Γ��ȳ��p}�TJ�dJ�d�镰ɞ��p�e��d���y���TI�@)� �����79�F=7�b� ���]�W�;��w�(5`�&��E�����f���v{���;'���)I�m2�v�:��$mf�6�`6[A���gvB$�3g�&{�Y'0�ݩ���������öe����>����1�g��qZ�^��Bl���s���
�=Ve��.������0;޼,����u�>�'vu��HI4�B =��;塚ww���Θ-`�RCuW���-����Iĝ��c���{��f{o��պ�p%��l�Y�����0b�Ɠ�v� ���Ā�s�K�Q7#�(������|Pt*.w���'�ﯮ��?�z�TJ�dHj�uh`w��36u�O��0��|M��l��t��7�m	t�뗴�c>�1s������益��$� < ���	9�v@�փ LX W��j� St�@Q���<z]��(Q˳o��]ϲ�A�s�9�9�.�jJo����ɻZ2��'��EDn�H ��o.��M&�b�q�N�iD��s/ܒe��p�~��" ]�� ��<�0�!�6Ѐ{�� ����$�wl]��2�dЏ�"�@0`I^B�z����2Ф�ji\��m�      UU���J�x��9chUoV۶[��Ϝ;�����EM�{ d��eGQ vx�=��4n��iw&T�μ�;��rU5�]o.�l�MJ�c��\�W�Q��ۮW��ܙM0<e����3ڗ��E��EƵd���]�U��5��s�$��P�G���,[m�ۨh���bNN.�\n�-��$n,���������s��/��2�K��Q���%�ʒ�-�g��P�G(��}�X�||@S��DӰ8��mQݭ(���vO��Ϲ~�"���W4�$�rH��'���ժ�⋪���L��i�ޙ ��T)���"!DI��k���z�wZ`fV��'RԷ#�2N���e��!B��J�ա�.�����Mm$�4��a�Us��
�:�ѧf��mf�:;2t�P�,�Qwv���&�h��=����B[{�G�Ok�$iR��&P��Ͻ^+�@�	���"p
'J��?q֯���������k�*��>G�Z�i6���0�P���pp#7z�O��:��ץ�vW�)�Њne���IIB;�� �t�Ӛ�>�v�O��	T��%�&� }��Xk�P�ooK��m�؟t��F�����l� Y���k�q���VΖ�<�N�P-n��L���F0:Vzg�+�w��\�s=o�"(;�4�����L� �)�!4X�����Q��]�s�As+
��*�y�T%	E�&iY'w}vI�h#�D�xė�>��FD��^C���3?w����4��N�ԍ�'舀]f��m�l���7d�M��p��i��$�*ST�����ZQ'� �wyÓ;�����`_�^6�m�c�;�5���P�q۪�u��ָn8�\7f������f�-�&��F.� ���){ҧ8�����Fv��)�R)�[�������"x��yfgyZQɞ���
"#3n˫	cM�ӦM7�;�5����0�^�l��޺�wt%QD�Ӓ@t�=
��{����W,��W�O���&�y�O��˓���Ϙ�qԉ��(��P��s7�.��J!-��8��֘�����ꪱ�Ny�������ӟ^���lu��v췞����-J�&�	��9���q�y��^�DBW!��j�nz��i�n�H���i��YR�������]�	(�B�IO��|F�)���C�����$�d�| �]08<�!�M6��&@����[{b�<mO�)��ܿ�&�TSd�ۀn��H��UW�F{�$���f�{�;�O��� �������]������[t�Ϯ.zj   �   2�\�v�9t�v��!�df՜�b����'�#��z�T�ti[�b�����\u<E��tط���0�MC�4;�g�f�ܣlܙͱ�&����)N�d��/m�	���rۢ(}�w1��Z�� �{k�����r�{t&�`���ÿ��{��O���UQuG�S�@��Y3�G]������E�%���'c�����
uQ<f������s�;��s1ߴDv���]��ﾲiSE0nd��^��DU|�w_Y�=��w:{��n����X$HXwz@fl�W%��N4��с��8�KR��sA4�����t���O���d�[�2���H����{2f��)���n����8��i~|��%��mr^γm9�z.=�.u�#\nשy?�������3p~������۷{�vf}~	$�T���0;>'OK�y�kz�������}��:Td{^���gy~�	>ք��i�\�d�ڴ�A�U@�S)$�I�{�w2x�֊�+ա�/ݲg1����M���S���ݱd�m3d�ލwd�D@�+w}��G�}s4��USR�*�'��0>��y�w�����'��"Md4M$�V��7Mi�f���ns���9���m���D���o�Y��
�ޮ���* /u��%7A�Z@�z�])jU2�PM;fg��(SA�|�
�y���s�;6Io=s�h ��E	).{��.e�nl�(������������������o�˵~��������W��<�������I'���̬�f}�����]�����s���N�`�A�)L�1�(����(�j��2�;����)��*�bH����$��$�!�:�0�ӷN�f���=�n�;v�G  �e���]���s�F�<��ugA��$[I�Ɉ$�2����B��u����K��tx� q-<"v� � �фk���5�Wa�'��8C�C�i5���$�Ym�%$b �� 5��J����2k�'���A��и���|��s��_]��?�@�0M�a~?����34e����a�te��mۻon��*�N�7�K���ݻw�ny�y�}�u�w��v뮺뮺�;�ݹ�{���wu��w]ݰ  8 �0 ��� ��� `�  6 p p��@p @@@`� p }׵�O�T>�R"P�}�_�…���T�GA�?��yDCN;@C�� v ��8�� s��:k{4yݪ�����0��G-;��d�2@���� �i�x ��J��!vg�@+��̶�v,�˒���L����ST��#d�����>�����%אNd�_��O��7�� ���H:�ImuF+g���v7C�۳�^-�G<���Fey�ij�~���{��w^��� }� �p�Kj��lES�9��@fWO\�{�w޻��7��&�B��R�����Bm��X�l����8��<�&P�U,�	������;��87Za��]rȫ$�ʽA�.¾���r��%C�y��T]$�l019�����i��]�=�˰?!%	-]���� T�V���Y�u�ں�gF��������u�h��O�.��<B�M7`b���-�S�����I�{vI���x$�$�N�u`壧����3;���{�� {��$Y����M4 �� +3gY?}���L��0I�� &�L�R�J���@��{�I���\�eȡ(�Ϸ�ex�M9�b��U;����Gf|���	9�$�s�������>���T94|�վ.g�7���       ����m�[su��]����xD#�cm��tu�/F7����N� K{m���i��H)��b�/t��6%��g/.��#�����r3�WQ��s�A�����g���u	���sm��&� ��{
⣬��J��i�S�������������ꪫOfb�5�-������]�{;}�:.�e���l�m��w�د���,R�r5��@w��`gs���!�y�3�I�A"�H� ��'W�_D����;�9'�/�J�(�IU���T]$�e��, ���8����τL��M�s:���N�K�:��	*T����%�z�g6X��5N��Y'���4�MR+������> @Z���I-�ݹڜZ���=�"�?UUP�ܦ���g��xڵ��e۸�g�&㛇��P�	S��%6�l� �:@��b۰;���(���͖ۯ��T��T�R�K���i����� F�D �)Y��[���0;9�`s�e��%�Wl���t�hQ�S�����#�4���_7��@gt���J���
�`-��`{��� ��^�OD���^a:�&�
I�D��3;�������$�u���N	�i$�R�Iݸ퍻V�=���u�p\[�z�i�R�7�Jx�&Ka�[�H�޻��t�8��� �~'�|�!��tn��A9���O{��rNw6�@�=��mxR(�T��	�:;$�w҉3޷�vG�b�9ܸN�$�9rK�[
�����r���ͻ;�v7Za��	DY��"w�!��-��wH �F{�$콙RO9����IJ<\&�ݧ�\����[6箲�q�{nc{u��.�}���hQ)� {�Ӡ>���_�d�@noH ���E�I� �j 4�8�{v@�[��q#s�I����F5��0PI�D� w~� �� ���sK 
��u�h%A�� � ط7�*�~���9\���7\�Ҟ�J0!
��߆�DD  g��J��pY'��L��I��9h|��^�6�e���vw6�;>�%��_�m��%QR��7����]��v��tZ����	R��X�o�i���R(3�fg�҉<�e�=�M���N{Ҙ p��e���`���a�V=�y����u��cu@DPH��`�� x��<o J�d������-�ТS�H�w:`9��.�$v�y��Xd�gBQB�M J�>�l��	۰3��9���D-��Q���
��粄Y˩T��m�     k�Xn�v�a�Nr�!>e�J��N�6z�':��ʪ�8���Zp�����s�]�n_=�ۀ���<�[l��sg>嬙�w<ǜ:�ZW�6���N6�.��\G�vv�%8��ւ������`f��곖Hj�2���;�w����T�K1��N��u]�x:��'N@�ػCsY���d��,0[j�#c�>� sze�';�� q�2B���Qƨ�J�l
v �ΐP��0�O����H'8��ԝ2�	Ѡ۰��0�y���� f�{:A�y�I���I�L��e� e|�>�I�=7�I8+>�$f��3'�`��KSaS�����޹d	� wŀ=�m��_^�pY�vkv;e�mպ켫c�#�+��F̜F�m�{:@8�zS MY�l���wZӦe))U*"L��<����D	q""��97sw$�3��i��8x��ꄪ(PI��	T q�� ���@�����2s|�$�d����5R��%# ���W\�A�� ��l� Ӛv�ڝt����e"[�77s���;����G�ݖ��#�i0K��m�P��],S��5�n�ˢu��'i.d���|}���Si:�vH�T�$4�,oݳl����'���U)ST��$콕��O������`�t��3 lSJiT��g����&q��� ~@�@Np1RH�A �K�lP�}s/m�g3�X�O2���I9�� F�e��a�?}����i#:`}��%�� �q��Kd6�B�K���զ�>: �_�g��/w�d�����'�ܒ~��
��QQ�^�p��u���*<N�.٣�=z7aV����}���~�� ��R$�o+�}�}UtA>ޔ��}���%|t�#`����˽$cm02{��IB�����Δ�T9l�Kv�}���i��
!D��09�m���=3��l���T:}��=��2���8⾔��}^׼SB��5��`�>� ��V��"�>�v�?�Z��&e����s� �̐�gO�m���}���W��9�����r]t�1��KgWrn"�nwl�)��_w�;C0�1���s�����r�����P��wkF�5� M%��v �ސBo5Ӱ@�Ǵ p�I����T�ţ�-��E�JpY>;Ƙ�=�CM�ɶ	��@�޹�UEJ��l`:V�
��^w=�p���<�D�}i���M��@۔�E! �� �l��t�}��h��UU_௨]t��9�)$Q���IE)$�I#�]��]�$�I%�]�ݰk�uL���<��&U��8�u�8�gC�'�s�8q�z;�]� �$���`md��B��)�4��.s�;A�*��0��C��]r)����z5B�#�9!0�K���X�lW�9���s����
ዀ��#��������0gbt��@&�u� ܤ](���8zj��ح&"A+kT�,㉋HK�[GE]�j(Њ9��7�%֧~��K=)��b�R�x��r����K[ﯱ�w�w��6k~��|9�_�m��$ q�$�                                       �8屗��W5��v�V�8�XI�J�-��Wm��ƹ7����g�6ͺ�5Lm�vy�cX��P��K.æ���'D#�-(�סvݧeѰ�u�Ov*�ϴZ�%m���v�.ks�bލG�Z��z��Ji�a���n�ӧi^e�	��,k�.rKF�;N�T���[m�.t���Qk,{��u�7�v��:�uQmӆ\��xt��]�d�
u����n�Z�W�D��2C�q�n3�9�n-�ؘ�`ۤ�p��+���y�l�,�ɺi�V��k/'2����4�6�ȶ�&��WJ�dڤ��H��R�Lj��)d�!�W�Z��K%f�n:0lUT !*�����[i`"m�k��Էvź�-ُT�<Pt�m�Z2�� {��H�Y}�ղI��GE;��pA�t��y���8��y�������YCҸ�*��j���a5�Jݫ[����^K�Y&5�t����P��a7=��	��ư����%��s^�Ih�K�)��6��{J�VK�P�r<�
�͞2T���Y�mn&]P�g�Sy��%R�B���4�q×����}��~�������ERR��ڬZ��y"�oS�2��@#Y��ׯV�-l�h�`���nv��0�g�@�q���)be�]��j�\������gk[���e��v׉��]��.ճ��5��n�k,̱nX��2յ�ש�M��h8����{ְ�ky���$�W���:PO�3�O �>�q�a���8D�h/. ���\P��@���T��t����/{�����9��^{�����}w���       ˴��K����y�g�.kE���v���;8RF�kp�g{�8ۮ;|~emt��v�K�>����1hZ<��j�]Wm6������gw��ݧ6M�ْ��	g�k����|ci>2�Z�%�w߼v�h~�xkV�g�L�/�;����9���P�y�n|��BM�%YN��Uжl�� wX��w~����u��s���UUc�ՙ�y{u,=fKe�{�5�|(t���o=��
S��Z�-��2j�/]���Or��
/���~��߉�:��)�H4�q9��e�9D�w]�';�{����~��T��T�V �s�`	y�$�f�� {y� �CB�)�SE��p��� 77� ^k�UY�8��%C� Z($�)�� M�ޖ �t�}��%�N�$�����$��\4�:-9�����<%�]&�]���i1-��ТS�&�l2�OrS�29Ѯ��N���>��{ݙ�U$V���V�qW��y����?B�>0I +���� D�΍{�>s�'�y��#:l����_�"AH���@w6��֘=�`�ڜt��i9i�%��͗<H��* 4朄�l�|���+��ԙi6�dӰ��1�j��� �b���z�uz�O[m��:�oQ�,�sMtSh��m�x����N����~�6�I�.�	���C {sc���{0 �u���m��U {sd�A�i����V�uD��k�Pe�)T�IY$nnݒyւ?� 	�h L�_5Ծ��
s�����d�u��%�Z8�)��Jv��gJ`9�3��fβ����߽p��	H#B��*���,����ks]؃��j��Z��UUi��i^EMy�����sq�y�&�9�t��X_�P��A�����{:� 77��>����s������T�L�h̥{2���ߢT�Z�$��;s3>���E����Ӥv(�m�Ir�|" 	�n��׾�m=�PL6�2�:%Հ�-��+�)�{6��` 7y  �~]�Љ<�����9���U.x��;;�v708��,"E�43�m��o�"�=x+mstM��|�C�����z$��{vK�%��%�u��,�����4��͜I\�=�v�-Ǽh��I�ТS�({���"�d0��vI���=�o�s3B����j��};�D�׏�;�+k}v{3:��{	�*@� � _f� ���p�0�J�P��鹿B[ߪ}*���IUH��$�~�$�=�,����=�;�O��=����=�|*\��I$      U0Ħa�z��i��ҽ������d�^z-�7�s�����-��r;a���M�3�<���m���NӤ1�lD�������\�[ae�1!��Gx��u�B�^̧d6�;�nTAVB���d}���<,A�ֺ���Ͼ���k\{��w�����UT[�7t��&��%v��<���V�.�t7]>B�#���}������-P����OrX#���O�%����H,��ߗ�2�N�u`ǿ����p��n�&Oq��L�N�J�J�I��fœ�� szA]U�Q>�t�sK$ڮ�K)
	�KӀ�t�q�z�@l��J"y��X���4��-�D���y�ď��'<���<w�� ^��'�  郵�$�EP�F���'�-�=F�c�K�:lQŶn6�uÿ����<��k;%.����`^WrU�d�_�9!��L��ṚNUT�	�D��O ��������8��D������'{^!���X3��J�tʢ�H� �� �t�Q:sK _f� ߎ�#��l�t�NőUUF��>p��4� {�H��넟�OExR*���@�$코I���v ���'��1��Y��m��e0�M���7!�L�<]v�sv�n2��l��Ѵ3ж�V ��w٪�=���	�,>��Zd����Cݝw����D{:�@ӚX�f�č�À)��M�*R�O��Œ\�r��оF�� *H����������K��?:�8��^$Oot$�DR��UAB�-�����sz�3y��G�OD�(P)�h�e�Cݽ v�� �k���4�7�~�g�����&�ݷK��Mg%��[ӭ�m�\hj�v��d��G2/������ ��� 0�u�<�d �G��ؚsN�����۳gJ=����q/�?�c��3IMR��'f��@ǲ@��g� �:�@����)�US%͇���������և'�-N(1b��̷��d�Gy^2G-P�S�݇��o�a�����9]ɰ:�n�������>v��
�]u����6��n��n+s�&^�^ڸݭ��ů��l;Z�r%���뭄j�*3���@{6H �n�e*4BM� J�Nit ��H8��� �t�����$J
h
F /sz����M�:`q�[����Z�%@�e�m"���t�q�l� �9��/��$���x:M��L�; {�� �OrY�=�m�$'7�`}���RA���w�>�[p       	wGWZ؉m���H{d�[Vy,��tr<<�Cj sƍ�Vy��2iN'��z�[9Y�5�l�q��Ƽ`�=x�#Ӳ�+H�{�]���7"��waY�+�.y:�]��N۳6 *��om�1�#)���Ӧ顗�DY#T5��@7:�<\��w/~�+ꪒ�kc�R���&��t�%ӛKp� �*�����n>X���)I����&�u���~� �� ӹ���|����,���d��YM�x}��{s|��;�i��ܝ��T���T�(�!4�$l]I׾�$�1\�@���{4�L��n�/ٙ�R��@R)�g:`}��f�d�uv�y� ��B��I��ET i�,��6���?Y�Τ Y��-m��-�h4������ڹ�'Nv�)v�]hKͭ5L��vR�5:���]��ͻ�־Ut9���S�jD�TT�
UT��%����C�@���?n�^As��(��<c���"d�{�\���0t�i�� ������QݦV?_��O��wS$�s�V�
iTЦ�k��|��uGW3m܇3>���1ē�՚�Yd��6 �oH ��m�����K@rt�6�m���g��3�=�ݎ�4V��4���q�u�a��-��D��˚t��ɪ����wq�v��J.Jٲ��wBa��"��,�:SD��p���@I������$v�T!Q��l0U �� L�H��~���Im�$�HPJI$�H��wwWrI%���8��s�1(��QvI�D(�$n#�0�3"�ѭw"�xg�$u�;��0̫vH��=.��shB@t��q2D�hN�p�����c���w��A���͙�F$N�f�4(�%�����Ȱ�4�'�K2��1P��#Rv]q�͎	� ����:HT�x����Q �Aؼ�O�J����όW�^���zz�$�K���Vd5�|�Ʉ����W	ݱ$JF�M
 *Tl��{vN�x��$�wV�rN�@�kNY��Z4�h2鶑N�����֗]�L9;�r09�۰2=�m��%R��x��x�өqu�c�^�d�M�l;��nC}�G��0t�1���;/fE�Z0����(���2�9[��Y$~�|�xUIT� eu֕�D@�9_T��.�]N���$��pr�JT�Ll�2ssn��l���s�;�G�1p1���e4۰�'s~�X�4�̮��?��]h�@�9`o�[c��$��}al�! R��S���J�H�UK�6p���4�s~�s�'j�V����m�l!�j���Nu�-�Ȳl�GB"k����p��p*�g��Q�����ܰ0�칤��� �t���$�B�m*@$� _f�č�� �u��|�?b@,�
����E8���{��>� /)�I���(-��Ò��i�r����<�w\�0�f���o\ \�i~��M����#]iD�7��z��ݻ$�����,!�&��C!`IǞ�Խ���ӽ���f       ]V�X�l27J���v�d.�[���gr� )�n2.ԛ˸�m�v鮳��W�۝ŭ9��8����U�h�K�{t�M����\�{<v���zm�lV�m&�+/Eq�]��)֭^����QG�u�E{��;���u�:#Fl��i�&��Ӟ���������:Ź�������4��՜���v��|o���k�����ӱ���l�r�� S�zՁ�͐~�Y��t�F%]�&�&�)�ܲF��x��L�U��E���[���!�l�J�i� {9���wi@�ٲ 3��uX$oq�*($ZR��D%�==����߮��u4����$J
4耒ޮ޻'V�9�i���xXl�U#m��m��4ӟ/n�#'�Wg�૊�cn:��ڣ�m�d���AtJR�K�;��=�"O]3� 8�3��]�L����á˙�4�> ;�i�W�舀E��ڤQ;/3yg�9�n�d���*��J�h���W��r����ZY��K� ?��	F�m6�	6g�舀"o��Y>�{�_v��H#��ǡ�$n������i4Ӏ�� =��u�;W ��gY5m��n��v����gI6D����c�/M��.=sb�o���:�rڡT��r{���ܭ=}�:�_�� no� ���P�E��Z��šh� ����-�ݙ�}�d�� �=�r$�B�E�$ �6@{6u��?}�$�HF�~���ܶX�`�rr�MV �t�H�?77��7�}u`
��D _f�;_gC��e��I�$�`g�`gk��~�2N���ٓ䒟/��
 *rʺr�u뫬��z���R�F7�q!�u��%���I)X�I4���
A��G���{6�w7�6Zf�]^���]M� $�L6 ٽ$�B��y���P��0 �����L��a88��� �t�'<�0��n�[���(��	�UK��H���wZ�d�c�s, !�t�
2�bKր�q]y�,�B�+.S-��XT����R��t0sTX�Z4{��`gsn�L�<���{����*����e���u�Zc���۶vܯ[H>�R(�D�4JR�< �v��szN${9� n-	�U�2]2�)��p�����_�	ą��w���ΎA�e6��.��t�$7V}#�]�۲y7�}�3�S�^�RV۔� v�3�?YsK���H@�qjm�U6S,9=����B���}�ߚw2-�с~]IJDB���f�����޽9ڶ�       %�SY���EZ�n�fһ�V��v��[Z�v�������k�)�bܻ��	v�Y�X�ћN����w�Y�Ρ�ץܫ����]m�-�.�.z��E�\�<�7SC�W�Z$=Gո��f��œB�Gѳ�M��l��.e��V;wq��w���ꪢ�l�x+m*�Z�t��]��=t~>���ck��:;0w�d�4C5~���>wg��ejd<�~��'<�쓱�W~$�KtCb�N���}�j���ٶ@���#V�BH��`2� /�	�z�Le{� =�Z$���E
D���� ��8��\qh`?{�"B�!�閑N���
���A�.���=� �P�;
 /#���%����Il��*��F麫�Нpz�e�e��$�	�W�#<�V��h`�� ��:���K���M��	By$�S+�B�����'ۻWd��m0ٝ7�܅Se1�������l�P�vʀš�hx�b%��l&�{d��r��Z]��ux<'�T�~���ֽ�&�tۗ*���{����U�$��.�r��,��3cE��I$��NΝ��<>�]��{��LV^�&Y�,Bt�iqmݮ�9��!��g�ͻn-��|�[#5R f^�HPH�@$� w���IL��۳�ߜ07+F ��ȻQ��-9uSN�����V��I$%
q" �	���p�5�el���n���gG �i�I6)��:Qd�aD�or�| H�'��	?z�¾�M&�t	uxui��?�����d���]�s<�{� ���m��B��jjk2ֹ�k��+��U��i�n:$��ӫ���9�o�;����۰9�i�����;�םI-$�aSM� �gI���G]�C�n;�3���2(%JQU3T��&o�07+FT��ܻ3=v��rR�E��P��0^���#sz@-�B���)�PB���}i�|Ϧn��d�] 
O�#�ސ�����=�!~f���H��~�4t跉%���
�=�鶫m����t�y�\�ɿ]����sb�����fo���u�ۏK;�Uwٓk�t����� Ӱ���4;5� �g]�_q��|;53���W�Jj�4���vXK�d��rIx��$�5K�g���4h&
�� ��(q>�t��C Y��I��E�Zm�{:@�]0y``	�� ]�/��l2BZ�I$��I$R'뻺��I$�K���y�>�EB�IC@��TICIq�f94Dfp�|I���=<����F���ÏQBx��w�:K4@D�^Ր
W%�H�h����ϊ d�َ"�ؚZi��Y��C��
p�X�u;�Б�5Б u�&��a�bi#�e� 	�,D��LGvKr$7�NSF��NRq���Z8$�NJe�b���%�f
a�) DB��N�k;<�%eml���Dޏ�eck�w�l�E2�D�������r#ߜ}���o�s��5�WU[BA �I6�                     =                 �^hF���M���v��3��l����Y^]�7:1m�ѹ.k5Ʀ@X:ɶ�if�ΉKW^�ȋv<3v'Z.��b�9֢RLi����$�m6���鄦v6Fn�l�L:�yg�q�euNō:�o�}�|c����tY�f}�X���	Ӗ�Pgf�6�N4*غ�N�M�F�>֛>�|:�F���\kgm��
��@�]�E^L欸���D��`x�ӛ�L��m�9��ZL@[#pؓc�v��������nm���6���+�5\[x�{uĭd��T�cj�f�.֖]��6��R����v�P�@�]���#F8�h9;7;���c)Ե �����i����}�[i	�R�4p���K%ք��v8C���qv��l�7W@r�.�[s��5f]��3��<
�	��v����/��3�gy�g��ӸJ�ʁ�� ���jT��Ki�D�'J6M����.ӻW4c�;i�A8�����4��E����	J����b� 4�T��ny�R�c��}�WU�&����+C�v���VAZ�'����5�q:����	��E ]ny��f���ͅ-��P��v�k��ٶ�r,�U��M��X�2x[u�^��^������K$��*�/)ur<=8��U�K���U��f���V�E��s`�.�7����'�^�G����Kt�Vm6v���5T�Z�k8ȲW$�1W^�f����5%*�h=���w{߽���{�b�����D��pG��@�C�t�ȗh�uþ�+wqw��>�o�	ߒy}�[�       �t]v!��1��wQ'�n�R1��q�GlΕ�����>��υQ�����u���]ғ��t6:�!-%��;h�.~0��s�����q|��a�[�Xhr�v�����������}g.�u�ctp�$A�4`�9T��$��$�	�h�M%A�X�h�@o�����H%�i�t]_V8%Ѷ�m���k��;�+��v����ks�>�s�m�[f6ݺ����������M2�$� 3u�d������:�Zsz@{�B"�e�*����gy�j�u��'w=7d��PAh�S׾����
�j���>��`gsn�}�B�o7�zN׆r]LW�ڙ
X��ӗU4�<�w~큝�L����6���:ySҦU4� �y����6{��X����Q�[m��b`��a��]��������Q�dӬ+է��v��w�~�9��զU4SX���0=���ɜ���֘]���M�ce��ͻ�O�����_W�Wѯ.�6{��G��H@�ZI �ʻQ-$Qm�-�sz@{v} ��A���[%�n:� �h6*���
s~�`nV�������]�{}�R�U44܎iw�'v�0>I(G}�偹�]���L�Hr�)��m��l\�f��8]x���N���a���w6�5!*�R�*������2no���zZ`gV ㈐�(�]2�)��77���}@@3闩IyL�S7��߀������T�42i��-���4�ḓ��ý��{m�0�٭`lz9���gF��$���ݐ���u&���Y> Fӕ�d����	/�d�u�ےN�-�2U6�P����vЧsW� �7�r�`qO>m��m�7R��/Ska9�Ս�N�\�1��s�Ä�%�fI��4sH �-i;����YP�����]Ĕ�m2�$��=�I���D����72������$���5Fj�"�d2����I�d��� َ��rfꪀ����X|�!D{��d����'�h"G�9� ! G4�/>��� È�Z�At�H�P��R~$?gJ�;�N�F�e�A�_y>�@%���sY[Jp�zطV�z�Jބ-�����L�I�< ok�u�$t�E��3lz�'^��,�]I��E e�wP_&O�f�-�]�~�l�(�١�@I�I�� /�dN���瀀"(
��'wPD���ê�UB�M��n ������r�w]0�d�I5�븒�-�Y���H�s� ��Z�d��}�w}v��	T$��DA��������;�����k�6�j�      ]#��/%�ܹ�j���m��+Y��wk��Y]FR��|N4rݒ�����w������C���s�b�q���h��l-{-ә5�<kj���v�5��]�<�gfN�§1�Z�<ҭP��;u��n��fw��C,��ݩ$�l�ej,���.:�DFq*E �m�將35�D=��8��Zʽu����=}�5L��G��ih�i�s�2���ͻ��?���ؒ%
EH �@�zOD�l޻�U�PD��
�2O}9S%�2�PR�)���� �Θ�wu� _f���9�ʻvR�������?��̹֞���	�'w}�$���W�#I)��ht�}�Z�7�m����'s�2���?~u��Nu�1�xF�K�3�۪��zܛ�m9�\�M��6�5L�i�MV �f�ƈ�ސ��L#�u� �ʴ��I�ۦ�3=w��*e�J!#J�ȷ�i�]�J���������Ja6�f�N��y�)BM�Rٍ�w ��]@�op�R$UX=�)2�l� nV� �>Z�3�Ȓ%
EH �w$��۲O#�p�g��';ɓ�!��~UUc��K���J�N9�Ǜ���c= ��ͮ�S)�Y-��)�{yH���L��~��{��I2!�:}EhR���i��ζ��	*�6�i>���?m=�����@�'�|�b�<x����LAT�]��E6��{��9{��us��#2�`RM��u�@�oH ��&{:U�k��0 ��:ҋ!"�m����� و� �y�7�vĎ��m�h�R5T�]����a�p@�5�w����u͋��/}��ioͬ�:S {1� N�L� �d nn�J�����sJ��L�i��ͻٻv�]0mn��(�* %Wd�v���$=�N���%d���F�Y.�i���� ���I��:�zB�e���^{�;��.����g�6I�Zt�I��ζ�5]ve\��{w٪���I� ��k��I$�[�8NZ�G� nj��#����t�!'u�j�?������R4�����MT��G�<x��2|�o��@�N8��M�@RM��dX<������9g&NT�D�� � �$�|�J!�Qm��p�� ��0�0I�����]Ĕ�l��;�b�Ɠ��L}� sw�Y#��BRN�!�P;�`�ٶa;���o4��B���u}K|��k�3a?k}��׷ո       ]�U]�Mr����b^�Kz2�c��0��p�]��w'6�2��g��c�<����Z�W��6꬈)I�vw=����w1ӻ�Ѭs�]\2��x��0ݓp^�b�]��(�������c�;h�rl\[�=�3���@bF�m���׻���������v�������~���O]���k�ch���{���wb8:�-��t�S�J4�d U� ~��8��[� =��=��$}�"B�.�t��`f�Y3<���cL����J&IQ�9����9t�t�rg������v\�7�d�m=����M e��X˓���,���vI�ZfI��l)d��	��Y#ݽRY �}�n��ۼ-X��5q��m�ܷuJ��������n���s��>:��<v�O��4�]Q7� 35��t���ˀ�[����*,7�����~�����ww��{ǻ�(IȨo}*}@� 7V�:`]�����������U �:h�U@�:cI�͐j���HgJ`P�ñ 4h@J���o,�۰��=i��n�`�=����t�H�4��� ��uвn�`�ͻ f���)$�l���%Rl�i���vi��Kn�Zru�wN��
��r�yG�'��"�q�$sq�rI�ͻ'g�OE~��m����ߝ>$^� ���� ��|)1>�D$Nx��ml&�����g���H3�'��8$�(ْI$�RRI$��$ۻ�$rI$�wf��uϙ_�BB�!�$�����n@t�]��t�Jh�C��8U wܑh�&\4�[97`�vijs�
s��f��!!�!�L�`���u�:m��!�iP�,H3�4��ϗB;;z9yS@�67�$=)�p���6�f8�A�!�`�̨�y���j���aѧ�Sh�"i@t>�ڣ��֐�	Fd �f
�A �׾K���}q���g�ժ�y��g�5d�BI�P�,f��^t��Ǣ 7(��E�l������A�?X���e�Q>�'3z���w�
a6�	�6,�g:`	�Vnʀ�� ���@�ysm��\NI�qtn��ll'X^Yy���q��f�� 4BL! �:Td�z�n��:~���_�ޥ N��H�� �z�H+�^�:I��%��i���O䣊c+�Ԓu

��)��~�>��öX׮�6���d _��tr�S.�L��3���/�{�03���������,`F,�fD��$�J�h`�T�`� �0Űp�!��$ \C1I%D1�Y�A"d&�'�� P�Iy���2�?Y>�W�2�u3MK�� �6#�93'��$l�6���q$g���ni�'j�12ޭE�%uvnZ�I�:���%DK,��	6EՀ;3z���* /��t@f�!ߍv�CH��E� ��{������ ��L;�"$mV����l��e�`�κ��:cI�͓���FH������eT�$w]�M�>Y'ݻ'�� y=�]�����$F�L� J�d�C4�{�g�3��;3�F�K�1" y{yQ�~yu�D
%���]2Im��`     I$b����v�gaw|���[�����<j�9:�Z�<-s�7h1-�p,t��9�K�]8��3��a-9�[�H��b��G<&�mQ��W0��l=�������a2�̭v ������' �d =��i�Y�;�mٻ8����!DDND,�	(_Wc�S�m��n�jPV��.�|S��ms\U����sfy�ӫO&{&�Ȫ���P��s�I�l�~�L������ _g3��e��I�v,�g:p d��D\��p>p�1�ݒ|���m��а��xb+³$ g���e0 �:Yf�M�u �>9� =���<|u���Q�l�	�]��H�i�Ӏ��dG���<@�n�D��H8�9�.m��e�!���&���;i��)���:��Ż1��׊�������Vi��n߯���4��t��� {;n����*�J���rՁ��?b\/RQ	F�(K�*���Pa';����t��H�ޅPH�I�� �P9��\ oq��|I�~z�T�@�W�@�R�E3)����o��L�~A�ǈJ�\��|�K'���P��Ӛ���L��4��D%+k-09�۰��{y`}�����m�K!�����f�m�uof륬\@N�wV-���������l����I���"�o;����w�d�栊�>����4U&�h��v�H�u�'�����Q
d����#��%�lt����%q��
 "ET�Ha!�ց���'�;��TCb"�<ξu����~�v ��u����	�o'�gJ�@�� ��n����"Hwn�$�!�% �49ɓ���d�T@�[��6NH��yd��n���/h��;I$�JR%�eܜ6�Bk�VN��N�����Ւ�kU�}��|=��%� �@wt�#��]����C����* 0��ĒM
T�H�sI�� slY.[����o�D;SQ�K;EJ��5M��s�Lδ�绗`fnڰ2{��S)�_��h䇽�0/{�f�s5��g�l��1"�BL�}��D�(S
%��̹)�`�f�R�5J�*2��I �� ���Γd��`fu��!��n��m�P�H�TJmi:,�פ#����=��=�Nd	O%�vi��vݎ'6:t ��]P�k� ku֎��H�e�����5�67c� �͐
��wē۳�+�`0�eT v�J���oH!=��q��n�Yt�)���H	T fv� ����O�?D-�N�`rd����I>�*��M���q'��v�b�M�$�gp���Tӧ٦;�4۬ ��    ��WZ۳�^E�wM�ͩ["p4�U�:��5�Ӱ:��-��e���ՖY�5�⮗XYb�ZܲX�u�LR9�<��<�+�Β��1&[H�0�p�q�.��̩&��j�ȗD���ݏW���n��\B�kmy<�.Ù"ڳq����3�ۻ���wq�ww=�߿y>�ϼ/�PK۴�ժ��F�S��&=]7vܑӷ=^���o�h�,��N�-�߿:b��0��*�����ίm.��i��r��`�t�:�������@�>��!�Iz�L�T�	�� 3���F�t�v�`�lB 3v�ZJ�.�a� �� &�%1C��eHEvmH����SMQE*�R���kL�佞��L������~䆥�5���n[�Zt�X�&bn����R�6zݛrݛ�Өv�ʰl;�;i��o�s��nl��=?Y�=��/wa(�(�tHK�H<�}�~ۈ���K�mTB��nQӧ4`�$]�A�*@( ��7q{�9!s;�'7�t vs�ā����E��:E�S��޻O�]1v��u!ݛ ��ΎA�Je'M$���L>��ݛ �����t���l MEʴ��� �2]��s;$瓿p̞�Ay�'��,��6�V̒���u[[����2�v�,<c��8���$4�	��새wp���t��k���k�)"�6p��Y@�W9�0�6@�{t��n\�5L�o��;�i���LQ�Pw�ml@�F+��'b<	���џf{�s}v��}ɚ�*�e �p%���S�����w]����wJ���J �A&�@J�?oH w��`Y�Z�;�i�s����m��T��m���+��z���t��q���3�Dt����!���&I�S�${���~�`	�達}ٷ \>���M�d�L����OI�bŒ{���#���դK8�h�iR��X���2w|�$�qݹ�ݧ����j^�w2�Sc$�M��Z��
;V�}�����Ou�w,�u��	�h��y4��N�ݭ���]����!�I"�6p}��N${�ӄ����ݛ }�m��-�4~N��&�f�e�p�g�6�����=<�]Drg�k��Z��sD��o�w������>��ܢ J��U�Ο�a�޸9�:@�i�(�V�߾�&jJ�U:(�,g~�q>�� ��Lw��$	��"� M��)�3�g>� �k���c��~�9�u�@�Y���S@�� �L��=�>̗�,���z}����۷`~�K��Њ"���$ADF���@�߫�a����C������0����{ǎ�:��h�*((bT �VT �bZ)UJQD�Q&AP� UJT(A)F�TrUr@��T��UfU) � iT"�Q��iaT��T�TrF�D(�b�ԩ��B �*���B�"B�R�%
�
*� �3 SELT���5��1�P���i)h��j��(�����(
����
����))(j�h);l�i)����(��	���*��""
z�L��)J%h� F��@�R�N.{0AܢI-
�R
+H*4�J�H	H�R��@��4*�!q��JP5!H�H�H�4�(RH�\�X��Y�%�iF�%b&P)F*JUB�T
A�Uj� hA)�)ZFe ���x�iD��F��@�R�H�bN�@j����e����"QQFJ)h
����`&���� ��R��bd����0D4+J��T�Hb���e�*�
����b)*��jf�&���"�'�M��LA22K1,��T3�DS5D�@0R,H%DU-��R4��40M#$��P�+QD�QT+�0DM)��LE!PTEK
��*
b;L�Ƒӯ���o�P?��Q)>���_k�wo�D?�!����џe�
���(�� ����(��� �_�!�v��UU��ު�l��UW��W���Q��߯�O��%U^;vs����UU��<0���D5�j�����������_�((�����"
"?̘���������?�����1���{��*#������������ZB�S��?��������3�1�/����II������3����v��];�DQ����ƹ���*��|�������D2"JJfY��I!!��T!eEB TT�R�@iDaP�T"Q��@h�@h�D	DXDR��@`!T�$D�@`YP@� e�bT)��V�����(��%�)dT
��KX���(P1%4% P��J���ȢR"��RHRD��DJ"���H̨ȅL	@CMAD�A P�
��H3
�R*� 	�(�R�#H4�JP���#J	J�R"4�#�*,J�J#J�	A3
��ҩHJ�@*L"�H��J�TB�B%C0��P@ĤA@$�4�D�B�P  �H�L�P4�1�5DIБ3 ���D�L#B3ARKL%BDP-- Q%!KMAH�
IU4P+25R�(8�$J�H�$�C0I$0���"�J2JI0�I$PL4�!2SB:<rs���{����k��v�������4*���x�>��?#��O�:�}~����?A��w�7������������B����?�i6��?�����C������3}&<#��?���>�������_��WϏ�?_���"
">�� Q����������?��_��9��t��#/�TDc���?��Z���?���OՇ?�~l;8`�����0DQ�}���Xs�|�H�<~��7���7�f*#�Xr)���?��i�:\�厎Q��?��~��"
"?��������}�E����?������~��?��}}���o�?(_�b?��wN���`��!������lU��?�������������#�l�I���F�?l����?����|/ݿ����#�ADGp��݆���A�3��~߷�_t��Ȩ��]a��O{���?�������0;���_�� ~B����yȠ�#����4�'�`q�nq?.:���#���iO��/��;��w$S�	��^