BZh91AY&SYB��߀pp��b� ����a`� @�        �  z      (�  �  :$ �J�*��AA@ )T 
"	I�J �)@PP�(
�   (H(
(    (RT�Q@ QC O��f��Uf��k�+�ť;� (w�ť,��뗓O[�n���)@���\ZR��  9� �p�p >�=S�`�@z�Z �@g�zs� b�h �J  P
U�ATJ�U��3����|]�NYJŕ=�� �|�W�.]�[qt���R�
 n��z�q�| �]��K��� �R�}r�l����ԬYK� S�S�����Sɧ�.U�˽��� ��P�B��"�� )��Ŏ��Ӵܛ�o{��_}� ��ns�NN.��T˜��� �zS�9��g��o�x�W��^�[��^��t�v�[��}n�瞗x u帷J�{�{�ݼwr��-J����TQ*
@(D ���徳��n__O���sn�{��P>�Wۓ;S���O-���/m�� {�J�|s=�:�-\���wzl��E��W6�omx�Nێ��O�[o� �ۛW-�w_sw�N.v�g���T���

( �3` >�����v����\�����x>����'].-w��,���}��>���}_5Žy�  �y2����*�� w���m��sۭ��[����u��炀ޥ�o��O;��;�[�b��|t�     S=A)��T�=I�C�CF#��O�l���i�ѐ` 	��Ǫ�P�Ji      =��(z��  � dd  E?Т�ڪ���@0 � �!&j�(�Ҟ!���L#H������O�����������p���_}���h������ UUv���������Uq ?�*���r�UWW�����*�����PUU������4����5�����]��Z��&,�����t�������1<�?	��	9m9x~9�����I7����n��Q�Àg���[G��hcا�����8k��~4oz�f�w:`�ߛ��3���4ꨳ1�?bѹ�ɔO��Wk��՟��L�)YiH�~)E?����|r<�7xp��x?�T��G����o�ʨn�]n׏��V�� Ƀm�>2�a�X����ӽ���?o�>ӑi���޼=�K�Ʒ�	���'��0�7��uc�����-YE�2<|�?b: �癭�]�:�i����Lts����2�V�xo�	`g�zv>��D��輘����ѹj}w�'�,�X}~��ᡲHH##_�p�y�l4�����M��\��F���Y��w2�8�&BQ�نK����^k�:�a�6�hݪ#Y�,�q�����tc��Q�A�9��Ċ#5i�n=00|�z�bˁ��5	Bn�ޚ�~���kZ�f�5��h�ݙp�<�N���C��Wp�2��o��y�:5��g���rW��?o��I������n�Nj��NOv������kXM`��P�`!���k=�=9��������|����Zך8�~2^9	���d�d%��97�a:�"0p2�D�)�᪍m�<��o!(O3^ѧ�Q�G�R�%	BP�8	�ͺ\��)pǞ~ݟ��x���c�o��^�����g���r2S��JqrC!��K�QE��!�y�1�&2��L9��sA�r�+264>NG)�jL������|��ޣ�yEe�-�Q���6ql�
�'N͇7ic�`�20�j�:��(MR�T.���'Do��O�h޸F�J^C��2�����</�
��6y��� =22�z�(49.;��<3�Oنʧv$Y8�u	~�?j�������n��K���<8����?C��l">5�a�y�c�S�����p�4���`� �<���J��!(J��?Bd&Bd'�L��MBR��۴>��_������<�1'%Ӓ1㚱�2����~�����y�����3XÛ��2�
�SR%.܄�)q$(JY�IBP���0c�>._��~�h'f���\���A��Q�S[4RrLM�^HaPBl���ѐ�4kW��E�k�S�ѿٛ�<����G���5�(�3�f!7	O�2�����~\�ޱ����Py�ÆT�P���0!̌)2!ѽdS�q캄�(ċ��((M��nx�������F��G�ԹG����[�UI��1�,M��D��;�FeDG��Ψ�u��	d�:���IFA�Lp���F�a�nȇ1�d%ٲ|ӕ?o5$峄a��6�3�����?@h�1Ө0��Ɇ���>��y�,�*�{oDY�ѭ��a:Z��h�r��'�䫔%~��Ոd�5�l1�?���9��~�U�Lvj����p2T	�������Y��qrL���,to���G7��� ވ2C�AZI�}�O�P�����M�y�%�e�}�(��� ����(J�nO���A�k�^.U��`k
�ѢH��?rp�y:����ߜ2�+y���\ۿ2���r �����k��L0���.q�]:�Z�ߖ��j�h?Y���0�# ���0�?FF^	���R?����JZ1����d�O5�P�(�q׎����z��]��E��	�������>��}k'�iS�9��9���y�!ܞ&`�I�������Iy��3n�sN�s6i�Z���s߶�������u�Z6oq�L� ȋ8x8���n繯��g�5^Dh�ڶ�۸��W��y�Q��s��\v�������p0\���%�ٙ�y��ǯ����:*�k5FBV��p��Z���I�0��J��,C!)O�m<���h��%�rԺu8�	X@nP�	BP�%	I��r0�-f,dcA����(M�P�%)BP���%MFɌ���78�)�ƣ!,vk��I�4�8i5�|�i���-$h�7��z� 8y�#a�#��V�:�f�K0J0k#52EV.YX�@l�%	By	C�ְ4<��7	C��J�����v	��#a�0�B ��Z3���g�?� &j"���M�3N.N.C���"�=ލc����	�L�<Fi�Թ�Jn�$�Y���9�Mu!�6c���0#���Z�>��K��<��bUO��B��^��$UiJЖ}bJT�jt�b�~M��4j��F�mڞ��kn�a��Y.9a�2��{��>��y㟈w����s����sr��F��jC3B}�Y�I���^f����5ff�A�2j��c*0�Kk3P�%	BP�%	��%�n�����ב����ߧ�xMBW�J�����	����,C%ۖ!F�|����.x��^q I~��C���9�he�;��$2y���K��%	By	B^	X�' ���?�V!��{i�P���# 4d�?�@d'���U�h?��j������d'ى��8?�5	����x��2BP<�	BP��2��	C��ߟ>W��}�v�k�_oZ6��Z#��O �����J�2���4h�n<(���ĸ^W9SZ�	%Rh��O��1fd�d�+�,y��t����O7�gg��M0UEDi�N0d`�N5.���!��Y��	�J�r��8sZM`3Q��8�~r�w��e�2��*�&\�/5��Fg)#��Th��4�La�Ԇ��AYAYddi�w�����%	Br%��6A��PbY	�0v`Xn��!(J��n��P�%	BP�%	B\Y�P�%%i������o�_�̃���0��>�ڄ���q��L��BP`�&��(J���%	I������Pؔ%��%��L�q�j`�BPpr�2�̓!=��f֒��d�<�;�M�'X�����2h691<c,'A��R�(�d'�q���'N�(��Д%����A�q,�/��2<�,���%BX%�<��n�`�'���(J�٨MBo0�n5dBR���ө�i�J����`20��:�IѫC��4A�d!��4�5��d%���F��NF3���,]����hd� �N���o��o."�C����ħ,��5�P����)0����s+AEDU�0�R&��Y;&���V�Zq��;�>u�����t�7���qݿ�9���:�5f�e�۝�F��w�Y?�\���� �x|kV���[��V�2�e�a�畫Q��,�0�X��pv٘ڄ�%�!(�$�J��`2v���>~��Z�	5�����j�����i�v��r8>��CrdFF$kV�|9��#F�����kq^����٫������g
<��Ec��,Ѭ4�ٗwS���rE��&)Z�Kߪ�*��Ŋ��-J�B��]��V}U�[�T�Fh�|9���?L�����>�@a�R�F�5�&����8��k܇�qrŌ�VY�3[5�����j54l���}��&F-���	BR�r�4��JR��(J�!�BP�xHfI�8k �ȃ�Q/���Y�ݻ����F-������7%ZXDMl+�_���wأ&����}�
�O�����WP�c��_o-���9�0���4��8���5��w����6�b՟o��n֌��#q���Y��Fx��Jp' ��]�p6�o�����M��n�7��1��058h���s���#4[�l6G��q�O��,�FӚ���i�k[q��8h-F�F�SEMa��Ǽ���:㉫Y�xm��4�A�n��(JR��(J��(J��(J��(J��(JR��(J��(J��y	BP�%	Bd%	BR�%	BP�%	H{��%?.���J��(J����p7���(J�7����	F���<���������4�4l�5��f͘kv:c55�C!+ 2q#,��E�o~~��kFFsF�����kPl<�\�E6fZ���%z�N����?BP�%����(p3�Ϥ�w���w~����3�{�����p�   ��           �      ��|   �
Pa��޼�`           [i@A���` ;���  �   	�      �            A�        >�             
�            d        	(   5�9���o�v�)Rm��d.Sm7   �)� ���C�U
%꫶��`l 6���m��wM�˻\Hm��       �|��T ����ox �[j���Pe2U6��  oi��` � [@ sm��� 8���-�n  �!m �i�h  	 ������e�B4� o͟   � w  �� 8��tٺ
ͯ6�݉���]/-`$I�p擄��JKn�J�U]@B�8H	nLm��ۭ{-��Q�i0-�#mͰm���e�u-�   V�/����O+&��� �x%��*��F�1�gk�Y�m��� ?@� �&� �Tv;J��Ð���Pm��v1����6��
����UW��b]��
�j�l$y��� :[4�� �)�J��Nļ�J�UPm� ��Z�8lҀ�m��9%�5�J�̵���Ő�$:8��[�f��
� ��I��� 6�Zд�m&�I���u�  [RI/n�]s�m&��   �  -�m��}N$���u��uV� �v�jݛkjH�   p�i:m���p [@� ����$m�p6��H�d�ݰ�]6�$ l��-��  �m�d��ސ��  m�ݰl��@[U-�*�;8n�'RH     �i���`  �%%�8Y-[e�Ƶ�Hְ#�����\ 6�6Im��ض�m&ć�j�D�b��K���ت��g��N;���Ⱥ�=��8��6����m$�Z �kl��e�^������� �`6�փ� �ݻ$-�,0-� *��B@�`*]�������I���!�m[m��` $$  � 8 �ٶ� �kn����M�`��86�[@  mUu-mP����:  6�[x[v�۶�6� l �l [@hi� m���ZM��}�kzɾK�� -� �Pn�L 	j���c���[B@���۶�$�m�H 5�L��ŵ     ��  �nP�A��d�;�  ,55�p
4�-���M����   -� p�`        � ���f^��l��Tb�L�+�UT���f���� �l�!��-����R���5p
� m�  lpWR��S<U/(Q*�P��I���@	'����t�� -�?@� 6�� [Ԑ[f�  ��     ���Y.�v�mmL��` ְv��m� �@m����U�P
�+[R�j`k� -��}�o�          �Hq���     p�m�m�� �	 ���v [#Ywitr�m�m ��m�'�I��0 H�]	��C� g$       �    ��-��%�	:I"���9���KR�Q�� 4-�� � �m�� v�-�Xa�8 kn qUR�f��L� 4�M`U�d)��Ur�PR�V�JK+q���h���2[��m���[��N��� ܝ�M����6��)�az���2�!���O�Z��Y]m�),���(,�lѬ�UR�-W@����ďAq� U-��
��B�r2@J�U�U� �ܪ�Hm0WV+bvU`Mҭͭ�n�l�ڤ�2�Ԍr�UUVҎ�`ڂ����-��T�l-�ٶ  �̀��/T���M(��R��[J�
�R�V�V�T��� B���G�}� [�+m�d�kh���p  n�ۀݴ�m����m���*
@�)2B�A&GZ�l���� �` ��vm]B���eU�%��U�l6ۃj�f  ��@  6�@   	      mjm���Zj�Yq���#R��ջI���@		�m�U��L�8�[B��Ij�cIKu��]�&�m��Xh���(�i%��[@Ãl�	 � 6�a���!�kn�[�8��.�Kchm�= Λi�*ඊQǲfJ�H [C�mf�Kd��C��[�M���6�S	e�f� �޴޶t�� $�I  )@ 		6�`  lh��H8� 6�n��5�wK���� �� ��k�k:ʹ���-6m�2�T �khW���>�} ݳ����[t�V���
�bO��}��f���m(�m���5�    �JP IH�e����RK�� �k5��ٛa 
R�5�/;X¬�YZ�]�)Um [@��$a"魸-��0ăF�(
�UU�*�Y��〓�m��ͺM��f�u(	�N��mnl    �            �M��� �ڶ	�$��HI�$9��IW����uT�uʮ�tٶ�	    ��pڥ\Xpf��ammn����Y��l �p�A��m[:mpp�i��/�J�UUuԬ�*�
��U    �-�Em� 6�%�1Ĝ]e�e՛   mY�g+b.�\-��rꀠ�j�P�U�Vm�`6<��Jl
�j�YS�d��#U�E��{e�J�AV�ȴ6��H��# -�5��  UP@�geԄv�MT�m5�mm���   ��{D�m'  m�   ��d(����2�n�Mځ�M�mj��m$z�s�a  6�fa���Y>��O��[�	� R�A2���sO.�j�j�� $ �d���n�*U���h����R��  �@M�q�m�Il�6� m�m�-�k ��ru�f.���( ��  ���6�6��ׯ����}�6��$-���}��MAm5�    � ���5ض���j�4k����\�N$�d8m�m��l�     Am qm$m��m[��nc��v� ImwLmz.l�Ƒ��t�� 6�  ��"���[A���m��f@�H����      ���f�l��`E-�^�n�����e�f�9�h�@@ �����8  ��7ɲ@f� 
V�)] ,I��I�@]3m.� ���������� 6� Ē ��^�	  �[@�I�     �    �cl�$�aM�[UKĻ=�9�aP��ծ�f�n�I��H�   $ sm��hl ��E�n��@  �e�]U���+��@��jU�N )"������u��܊Wh�[�"۶m��)��f�    ��l  @�`8����    Z�n�գv�%�Jʼ�.�*�*p4�m�Sm��M�m�`m��-����� m�8�@  ��   m�   ��        �`m���2�r���B���Ď����m��"��n�� -�   � [D��t-Yq-C�#.s5J��l�_}���睾���^�� �m��� �H�i��j��`6���K(����ݛ6E����   "A8   
������� �l�� 	$ m��v���`   Im��l�[h[BCmm� ݤ��8m�Km�H   ��J �` $l�i8 [Cm�U   �\�`@   h   H 8 m��HH  խ��B@  "iC�k��}�$>�m �  Ӏ������HI-��[@�f����J����:Ŋ��S[�  ����_��^��l  8��ky��� '�uʹ�S��t��n[Lr{v+f�3Ks��UT�m����UIjCR��l�Em$ˣm� ��D��4J2-UAg��2�	�P	$ r�-���Y"���9m�V	 )R ����� ��su�#m�?���r����UW{���������?�?���������T�	�G��`����B
�& ��B! 
�����0����y���@�(���G�'�'¦�M����?�)�� �OEGh�+"|qધ�/��1& P�� 8��6)� >ȧ����OƑ$�)�ZJ!F�RA�!h�`e�	B���jRH��"YHA! �
D��!ih�>S�W!](�a��?�@�!�Q@ ��i( � "�_�ހ�'���@ �A8
�*�4��A��OTO6 (~S�~� �c�Q_����� O��Z@C��'��������W@���:!D <C�?(x��`= ?�&����PUU������_���������	(PY%@?ȅ1)��Ot������������`  � 
P k�       l    � dk�؛K�,4��IV�j�'F��͜Y�9`�%�)��I�Z�y���cPM/=�ͺ�� f6ڈC�%f�5��=WNC�/K*&�=�9��{� �3������� V�ӎ�h\9���� �g>a��e����]�Ҧz��l�X
^�C������U����-� ��z6�.�*npѶ���g;5�Q���:��%]�W86�0IsK�$�֤�P�bxKm�A�x��ԅ��)B�&βx�^�a� �W�ӬTp�����(gJ*�T�9N[��eI�cvA���I��mڝd��E�[UYv��{m�#�eՙѪ&�B�@mm�e��u�i�f�����M�s ��[uۢ%�.*�r�Be�ڛ��\G����ks�禬'b�veBn�(:k�3�3����4I�J�v����"ύ��  
�*��q��@\I̻�20Q,��Ynꮛm�u�ܕ��[�Dʹ����V�v�FV�q�m<��.K�����e�q�+(x!����8�l��ʻ]�f\�[�����` h1���,(�J.	C4snp��8*��E��`ֲ�y�8�4kaCvі'�iY�9j��@�4�U8nN�A�
��J��nɵ�È�Jp�I؆w%�%g�m!خ��y�WfݗXӱ`q$�Uv�6 f���/J�;6*����|��i�ZV	C�9:�i3�AW+�+UT�UcA9�l�aw��7"�F�T�����7!��,MJ�WUR��Ņ;<2��%t��Kh�l m�m�(] �5*u�-,�񥂺n�,��m+����m//T�SJ�I	�'F�M+H�l	V 
�8�تV{m���K;b��J��u��N�h��F���ꕭJ���x��7e>���ww���� ����A�
���8�~Q��k�7����V���r�UO//��O0۬g�ޭ\�h�;��cd�0\�gn��XV^�7k�G=�3�O�K�]�\�;��c6 �m�F!���9��	�����lpq9
-��wdۨ]�$)���]���[c�j6�];G#p΋+�Iǝ�/E��"n�Ogy5�ڶ;v���vI�z��I������s����27[��7k�n{��{��׽�-ڞs�=�l	�x�/gp�n6q�2� ��l�|bBMcLāq9>������=��,�_.Y�X�&n�J�*I����qg%	$(�Q ��0{y� �n��{V4��㙉��&�p�рr呀��.YOA<��&��.~��0�d`� K���F����-F�WER��ɛ
�� \��	r��%��%�# #�����9��qki�w:"9z�g=����{V��;�KnƸ,9�;YC���iua�ث���9r��+F˖F .J�{f6�g�n��s8�f��s>�썸�#�<�d`�+�;�d`�3
%D�6TM]��,� \���w��7�4���ki�䐟��0rW�w���+F��# �@�kĤPCF��wۼ� g�}��h�=ܲ0rW�trUXE��wW6wl��N�=a�$81�FM;�[=���̚ғ���$�i9�|���m���pw,� \���d`=�qSw UE��Uf�呀��RY�h�}����d�cy��0ng 7���W�}�Z`��&!����¸)C. �
)!��u�Wh�=�Y��R�ꋺ���.�j� ԖF �Z0�Y �+�=���A���&�p�M8�����^�,����UQ4EQ.�c=l͕#S�=771��s�!���{n6���ׇ���Owwq�9tȅ��ߛ	'��	r�RY]h���<���ɜ ������p�M8���p��L��у$�����F}��# �x�ƍ'���ͤ�4���� ����U}��o���>�AT�<�]߹�5~�z�N G�|�� ���� %��Id`	u� }�L.ETK�[^C[�.f3�׍L�X���'�����)�z�K�}�������i�[����� ԖF �ZG�l�I�`���7% `�rN���p�M0�Y �+�;���D��˨����j�0�рwr���^�,� ��<zb��,m��g��{y� K�����呀$	UeՓw$\�U]� �,�����6�F���9W���~���Ifk~g�&���v �[V��DV"�Ω��y�r��k��@���x;R)(��v��O3l��M�vHI�ñ���Y�g$��<�y�ẃb4�(v�Ϯi<�5���7U�[S��O���u�7H`��q�J�!5s�O5�7-m�ێ�v+8��3g�%n��#^�,�����v��.���fy��V#	�����ټ�N���gk�+���/0Z��Q(��l�ͧ8kn#��8��P��@�y��S��w����2n��_����F �,�w,����d`�RRƒosI<s8﷙�7��g ���8���p��ܑ�L<��0ܲ0�d`�d`	r��:;��QU]Y3dW\�0�0�d`.呀]+���.J�����y,�.Y�Y\�0Ȏv�C�9�w�9���ӛ�����#��cKt7I���8�덜9����.��/=5MUƀ�ywZ0�d`�����ǦF�&�����y�英Ž�,�.Y@�VM�7rAQAEUY�%�# ԖF �,���Ӏw�d��"f&<rL�Id`	r��;�р%�# �򐢦f�}%A55W\�0�K�6�3�wwy����O�L��0K�z`��k\`��=���y6ǎG�m�T��9Y�̑�L<��8�� ���8�Y\�?[�P�R\:*�˫&l����x�����G�x����7�N ~�a�"���ra�&�p����_}��9 � ��T�Q{�o\w�����M���#Ǒ�I73�n���r��呀jK# �QH���*ɉ����;�р%�# Ԗg ���8��������� �D*=Y�ZK��;ml��Y�ݮ��>��9N`�m���H&���mÀn�y�������g ���p��L��10���`���呀wW)��^9��0�Mߐ�Ong �o3�{�ڸ�������F'�#��X����B���8 ޻�=���-D-"��g�fĽ����j&k�G���p.W�/%��%�# ]\� �������\�x�7s�#q"Nm��D�q��2n�i�:v�A.�J^`�8Vդ�N����y,�.Y��8 �+�=혛ų�G�"bI��w������� N��0|zAE".���&*���ur� K���d`	v�8�7y! ���1� 7}��jK# K�F�\� �@��QSw6D�AAWw�jK# K�F�\� >�߷ʺ��dR��}�n�[ݭf�  gft��\�7�}:�UlOF��m�J�[q�\�\�v��n��gv�'^vRMc.���;9;!�#3@<n5���퉝�"m3��h��ը�MVu��2�i"d��I��$/T؀t\:�h-��fђ��D��z�i%����]2O���BK,��.�5a6����9,�l����g�}s�[Do*�м��v�7k�8��b���V���-�k�M�Q�f�ńF�'Y:u����m��
\�e� c�����<i����/��=��8\�0�0]tM(��j��,���ur�.Y�Y\�0g��&k�G���p�o3�o��XtD$�L�� ��� ~ߐ��n�n���*�� ^K# K�F ��N���p{f%�l���Ș�ng ����}�5i΀�y�Y��n�0Nu�t�l�OGf�8.�N�l����,zۮy�Dn�G1�tu�p�^�僗-���8\�0�0�d`�'ȤS �Ɯ\w����}�a�˱r܌{�F ��N����n�����0�0�d`���}����@c��pĞ��w���W)�呀/%����QwD��5d��B�r�}}���<��\E�-��qE$BB�|��q�f�+vnGG�f7Sn|��[�%������n�.,���N��Y	r����yt����*�	������B\�!w�d%��=�wz��B7�1$��n�ff��������H�M1Q5W��	��G�,?��!"�l ��f�&f7�� ��I�3h�e"��!�)�a61�K�.�
��YEY%��.����ԩ�`A$��@A$0P�`��&Fa0�A��bdb��N����Ą����Ca�����h '��"�JX�JVddԋ�R�������>5�J�kH.MT%m�0V`�Cc�c�H$�CA�ф�����$
Z��fc�һe���a:Gh�pl,:@��*�=U8 ~C�+�����<�a>@C��=���AZR������җ_s�����l�o0֭kg�T({��w��)���AiJN����� %)���R���h[d$R	1��ffb�s��O��S���8(Ҕ��߻��Q)N���┥~���G�JS� }��̬�_�hgv�mufJcO�m���/lհ=.���N����uW��q���Rv���JR�����p|��{߻ÊR�=�߻��R��~�)JR~>����޶f�����|��;߻À ���?����%)O���p┥%�v�>���}���'rF�ɐS�┥~���|��;߻ÊR���߻��R��~�)JR||��ݵ����n��8>JR�����)JN�����)Jw�w��$:(uQ� !Q�LD@$�e�A�<�}���%)K��w���z�oz�5����)I�}�x>JP��݂��~�~�߶����/bc�L>@̍�$��BgD��^���d�m�y$���ӵp��8��x9.��zS35��{)Jw�w��({��w��)���qJR�����|��.��sYwm���o0֭kg�(~��w��#���qJR�����|��;߻Ë�����7]�A5 �8���}�ﲔ�~�8�)I�}�x>JR�����)J�����)J~���[޷�4kz��)<=�w�%)N���┥����|��;߻�)JR~>����5����l�o{��)Jw�o��(~��w��)���qJR����y�t�����Ͼ����$�i���a$� 6nK��cv��հ��4k�rb�	�v
�N�he^��3�V׈��9���v��;:�ʜ��T��1��&�Rz}��l��T��Ơ���ϒ1�����S��]�P�d�뇍���j�R-y;rtD<�v3$�]Cv3#=�L���.w79�b��b+�A����/�D���&-�E�u����,YL1u�n��ږ���V���:���ܻA\c�A���צ��[\�x�3�[q�-*��WS4�.mM�ug�D Q�ϱG�)N���┥'����|��;߷ۊR�������onn�n��8>JR�����)JO߻��|��;߷ۊR�>��{��R�����y�޷���Z7���)JR~�����)����R����{����{�xqJR�ݷƮO���(��Ϻ}��e�)�)J}����)Jw�w��)?~��>���}���Pv|$�,lrR����{����{�xqJR�����%)N�_w8�)I��浖��nJ��:t�z�wc=���/nI�:�K��G�=�2�t��}?Ea�ɾ*��|��;߻ÊR���w���)Jw����)J}����)J~���[޷�5�l┥'���x>F����$2��Cr�����qJR�����%)N�������'�zr���Z���Wuw�<D �]��r!�>��{��C�2S�����)I����%)O��a��MoVhۼх��8�)C���%)N���┥'���x>JR���qJR����3������l��7�p|��;߷ۊR���w���)Jw����)J}����)Kۿ���/~�ś�O�m;]΄�^o!6�VÙ�6�۰�������6��[h�k{��)I��{����{���R����{����{��qJR���0��n[֍�Fo5��|��;�}�┥����|��;߷ۊR���w���)J]}�;��mf���j���R����{����{��qJj_A<��$��%)O�����)>5��2&�Ę��$�3�}���n�p"ZR�����%)N�]�qJR��}�x>JR��]��Fo{�����qJR�����%(�	�����qJR������)Jw��n)JR|}��/�措"�s�b;\�3L%�v�p���Y�s��n����=����@֯a��[��JS��{�R����{����{��┥'���x>JR�g~�Y��ޭ۽h�޷�R����{����{��┥'���x>JR���qJR����3������l��7�p|��;߷ۊR���w���)Jw����)J}����)J]����f������ow�)?~�{��R��u�s�R�>�����)A�T|1s�s��)<������a�ћ�o|%)N�_w8�)C������{��qJR����x>JR�׹��j�F�gxI��ً*F��<�7Q��{d��n���u�l��]���2C�6�9uG��m�v�������{��qJR����x>O�}����}���f�Z�ȦDۘ�����s��)����R����{����{���R����~��JS����4f���ވѭ�w�)<�����)�����(}�߻��R��~�n)JRy��,��7���٣{����R��u���(}��w��)��}��)I����%)O���Y��޵���֌-�y�)J}����)Jw��n)JR{����JS��{�R����_���J�k$� �r���YSG��\kB�<ܶ����XW����N���k��GmA����XN؜���$�c]�ȑ5\eW9��5��}Ӿv����TբDfʥ��=��m��A��-���==�s�\H��b)eI6D�npwJ�;z����쭎5��q�xÅ^�J�2L7</����ۧg'Y�&5�)zlk�tS%�-̇6{�A��e�Yn ��9�cp�ִ�V�Vݎ��Þ��ω��9����]c�����JS�����)=�����)����YrR�￻���R���	�*n�K�D���2!B_~m�G�)!�������)JP����>JR��wۊR��{ޙ���ְ�跚��>JR���qJR��{�x>JR�����)JOw���)J]}��Y��[ޭkvսo8�)C���%)N����)JOw���)Jw�����>�6�k�L��0Lk�s�Ϻ}�R�����)JOw���)Jw����)J}�{����\�����G���z��mm�w\E�8Fcx���jOWB<�Yۗ���6�J��K8�FN�;v�{����￿��>JR���┥�����)Jw��n)JR{��;Vwy������7�o|%)N�]�p��JP���x>JR��wۊR�������)]�f�kz�ZٻZ4[��R�>�����)��}��?�$��������������R��z��{k5��o-�����%)O��xqJR��{��|��>�_w8�	��������JR���7���h��X�Z��)JO}�{��R���}�┥����|��?}��┥'�k���F�n,�-��l\f͢&�͢���͹�۳��u�˞��M��f�S��}����m�����R����~��JS���)JRy����JR�����Z֬��޷�R����~���C%;���ÊR��������)J}�w��)@�4�ծE2&��1�|s�>���}�w���)JOw���!�^�
�jSZ�{�R��������)J{�}n�z޷�5�l┥'����|��>��┥'��~��JS���8�)I��ڳ��޷�m�ٽ�{��)J}���)=�;�t>JR�w���)JOw���)J{�:f��l�k��u�V�ks�$�ķG�����t*n;9��u���G%f�cr<lV�����=�;�t>JR�w���)JOw���)J}�w��)JO�=�;�fkz3vf����%)O���┥'����|��>��┥'��~��JR��3k"��"K#ng>��>�~��>�R����s�R������%)O���┥'��ܮ��Z�������R����s�R������%)O����&l%� �� �jQ�	=00%A�iXA��X%a��0Yp` %����=~Dy'>�<��)J]os�3]�ZՆ�3z�qJR���߻��R����)JR{�����)�u���):}�gn�7f���F�[m؄j&�\S�ۂ�F�W.���F��u��4mq}�}�EЍ�r;���~o{��}����)=�����)�{��P	rR�����>JR�|]��h��7�3th����R����{��?�	�����)JR{������JS���8�)I�s�gwf����4o7��|��;߻ÊR���������L.�ز!BZ��x�A�^ʩvkz��f�Ѣ�l┥'ﳿwC�)���8�)I����%(?�������"D �����*j�J�-\̙y���JS��xqJR�߽�x>JR��{ÊR���������C��d1Vc0V3�������ٚ)]�V��0��4�%1�4�YIJC��F! esv���20�
B	*	d`�%�B�C!Q.�$!J	6��L�� t����(JBI(���r"���Ĵ$��HҺ-8L��1��-.����k�f�C�k����x;�8pH�����c-���p������yc�S�Fd�z��U�l���uM�H�B&����3[�V�ҰR�CA)T��@���� ���A8���)�J��w��a�����E�� Jh&)�����A�� �g��/����k�    l� �,� m��`�      �   @%�t^���g$����.�+UU[m`u�`����j���l� [KN����H@:np�A�+v�y�ٱ(S�d�YU���f��u��`
6�c.���tY �=� �������Q��@������J�!��@�Ìfk����l���=���їg��ɓV��ҭT*�jC���j�2��'��;:�͍�"�;`עqִ��k:�]H�*�r�n�Y-�����9��wX�c�]�;8Ed�qg�s��`�U*�7�6��mcZ�[��ok��z��Lu� f;bUd{:u��.����:*�n�u��9�����UwY$�K��`"[��cBI����r׊L �5�*I�;l�\��#�:
��ה�X�Kz��iЉ�"��HuT��L���[n�J��s�D�Kn�V8�4�s�^nK�u��{!ns�$��{rg�24�ĺD��:���&Ŵ��%�x�����;r[-���@����26���g)�.8@8�Z�@����m۷R���.�Q0�0�����U[UWT�g\ h��67mb4��ڻ쩌���Sl�  �ɦ��;p�ۤF��Ulgt-Ȅ���m��6�T�n�	諚�	^��nʠ��quu&\v��UW/��f�b�Q��;.Ɏ������I	7Ab�٫��#���8�����)�� �C�ieIMWkum��[I� � *ꮠ���vtR��+y�gp�2-e �L�%�j�\J�dc�4�UUV��B➞xȵӊ*�$�[t�i=n]�n�+ 9���Y�j�()#�[I4�et��Kh�  -�n�t�{JR��K����6��\�{��E�J�\�%7m����mĒs֒/m
����n
Z��Ucv
��<�T
�m�� �,��[n���8��L�JÖy�c��A�������ONٴleOj�����{�����~|�|���A �A�D��w�߷�߷ww_}�~kcM��  hҽ9�`뫍;��]����N�u�jq�R�`�]���[�����=�f�l�7L��yA��C���%%+i�[/MӢ�8���ҥ%����N�N�v�>p9�݂�xD܂�5�jl-�^�k��R�Nsm�r�utQ[qR{qf�6��7#Sc��:A��AP`�j��7;3O`�rU�T����u���j�ێ�.Ĵ��Eɬ�cwf��I�5� �8K�]��0�km>6�H�\Q�\���3[��f�����l�R������>JR��{ÊR��������~�xqJR���ܮ��Zֲވ����|��;�{À�rR���k��>JR����)JR{����JR�}�Y��Z֬5��Y��R����u�p|��;����)JO~����)Jw������\�dM9�cL\�Y�O������w��)=�����)�~�)JR~����>JR��.��h���z5�-��qJR�߽�x>JR�����)JO�w_w�JS�}�R�����l~�?��[��v�#ZT��0���5�qv�q$��#KR!1ʒRQ���V���R���)JR~�;�t>JR����┥'�{��|��g~�Y��ފ���iR&�`�����(P�$��$�!*�"kW}�}�W߽�|��׋:d�ZL�T�]D�V�fOfexn��9s{�>v���s�A	���\)Y���[ށ}e8�j�rJy�� ��ҎWpU%�ww� ��0r��@M��y7�}�a���9�{u��4s��ջ6�.�m�ۜ� t�K/,q�8����bq�ې�� �%��O# �M�`mj�"�N`�����o3�w�߼��`���{��2n��ɥV]�Qr"����~����m�j���g���S�_[���ZĬ#qϒhrI�i�`䱚i�`tO�{�9u1XH��,���9���4��o3�v��]��z��v	HE$I2[y-3���9��䓗�d��F7pi�Gk�FD�("H��:�y����@N��ܖ3@��殢人�����y7�t��䱚J��-�V$���<0�N��j�䱚Jـo&�@	PU9�n��䊒�� �%��V�y7��3Oj�mj�	1F9�cLo�:�l�7ɽ�Rs�{�c472���Yݶ�uf
��j-��.��j�v�J���	۰���u�ժ]��Uf�M������3@|���f�	YnO��9�@�{W ����@��N������b����Y���� ���V�|���'8�E�'(���$�t��ͽ�Ss�w$�4-A�ʻ������&��7�{�>�� �I�h}�ܫ�����H��{�Ow~/���ʛm�  3�ʷ;Z`]�U�IYΑ#�P27�P���e%�q=��[#�ΌͿ���řT��B�;m�#�.�n���Px��':�..؎Ӟ�����t��f�xu���/��5�j���UJ�N�b�$NP/0Fh{%�� u�UЯ�=;I�r�J�4[S9�gO;������g�צQ,�V�m�v����mйSa۷www�w��g�9�j�����z�urdtH�%]
�h�6�����Ӓ�:=��L��m�<0�K@����p{v�:ݶ!$�!�{�� ��蚮�StU�"�.�p��~^铛�0������<��Z�I�2@Xَ9���)�;�{�>�� �i�h�K0��. ���0�otԜ���Ɓ}����Ta#R|'���z��8w7��>V��m�㛪�&�Ί���'c��&Ku�Σ*��Ǔj��=�v�qGC�[q�e�.]mg��m�����l�=������07q�"&D�7;���sٙ��1�ޯ���������IL�{���ʫ�����s7f�����V��>��~^�e8�ʊ�>�#�	$�@�^Հ}�������Q?���� ���3]Jf�.EJn�p��_���O^q�?{���w�~�j��Pn�1�N�0Juv��B[�[��#l�g��8PƼr�S��M��w�5�<�d��6cns:�e8Z�@�� ���45�&.˫�.DZ��0~m��	(�'�O� ���/��N�f��(ܟ	�r9ށ��s�ws{j���y[0�otKSIXF�Ɂ\���΁��N��o����N�l���j�IrZ��5w��.V�|��Γ�����7?��{�.,ܰ���hv��t���ŏ3��n{]7lq��۷i�ϭڻs6؋����� ��{�y�s�wr{���n�ED�mᄒw�~�j�ܞƀ�<�|�� p�T�Ӹ&�.H��������'��o�{�~�j�j7]$�1����m�gC��	DK��Xﻻ��s������m�����$#��L�L��m�@�� ���4��`
UL��"R�=Om(#��1��N�t�\O5	<��Y'n�<i�R�&	<jG;�?W�`ܞƀ�<�|�����˲ꊢ�.����<f��<�����{W ��72"dK}��7���=ͽ�<�9�;��hZ�)��1��ys8�[{�?W�p{o)�7�y�m�YQ'�Dxa$��t����4��`����������U��&  7k����Wn�����@s�R]��:���V�v����>�3ݯ��ܦ��S���/�'[�7m�I�]ѮU�Gvѹl9\���{[��V�+ӻ'��<�Z{�k���K��[`��A��5j��7��`[i�p�G���7e�����������u`;$�ݺl������o��ؔ묄n$�!��ϳ�fv�������{�˾?2�w<�r,q�m�Ɇ�Wjy��I�� �5�c{(vW\���@����	���wr���-�N��<����Γ��F뤘�9�`5���7vS�o6�@�� �V��j%�2]�wQ7 X]]�ͽ�<��;��: �l��j���n9�'�H�z��Xr��@N�������]�TU�D���ܭ9�������{W �����h�'���Ҙ�0 �.��`�&lF�/m���Z����u�u�*�>և00r'#dy�?s����8}m�@�^��=�W@���r�%J�j� �Ϳ{�d��Wt��o���g �r�.I�F�I'z���ܭ9������ p�Q3N��q85����ͫ��w����e8Z��!0����K�����y7��'8�Zs��2�rbk.[[�k����Ä�p�"�Ge�`F��7=77��s�����k�A��v�خ��}����0�m��%�@z�����3ʦ�I5Wu~���0r��@\�F������˲ꊊ�74�*��?}��|���X�bNP:�	$@�?�L��h�I�%C��h~4�Ŕ bY!e����E%�N����₟���"!|<Du���D4 C��� ��$a��d�	$eY�IBXMi"4��?�-�a�d�pd�B��?B��+��/ �N��@1RP�O&p_£���Ͻ��������y��lȇ�$^�N��<�y7���`�m΁U�c�	�ڑ72	������~��~�m����X(���.�P��f)S���kb76m4n�k� �'�	��`���p�"&4)�a2L�yI'��{���`����0rotÕEU9�����*&�� �'��'��{�{�~�)�*�n��c�6)�ry�7���`��5�H�R<S�&)&p��{�?W�p���t>�g�}���7�V�W��I?��W��'8�<f��<�ܛ���v���������\]kh�<��݋���L��*n<���;m[�ЅiS7I_U���O�.O# �&�@�� ��j,���X�ȅxt��g �ɽ�<�9�=��4-��ɺ���.�$���=ɽ�<�9�=��4��8�5�01��xa$���ڸ��f��<��7� �ʢf�6L]\�17W8��f��<��7�W����*���BR)�GR��%�dL qr 0U���}���jƻY��}�2V�t�[��1G^�Hs�2q눩 �]7����#�����j�cY�6cb�N ��pAE�r܍�6ӭ��p۩��&�o;�Fu�u�h���'��e�}v��[!F`jv�ٰmf&�;ٟk;�/7m�:�$�����v���F8 Lԩշ�����%W�N����\�uJn���02�v"w����www���?7IbR�Im�i8m�Q�n̆�pV���Z�sWBLck�{9�mq���v���]�~�`~��yrot:Np��5
�H�N<'�$��[{��{W ���:�o3�~���%q�Ic��u{�y�s�w7��'��w6�@�eM+"m!�?��pz�S�o��8�m�@�]��{�5D�n,I�rM�I�`ͽ�<��;��h�Xݘ��1�"�6���M�v�]�-��l��;�1��p=�$����3a��&�,���;�{�y�s�w7��O�V�M]�UE+�"�����&=�Gވ��;���0���­��Iǋ#&,NC�{��wo3�{�����p
���0����WY���Rysot%q`{�b:���H��'ɂ�g ������`��4���<��K	�s%̷uq�M��vFy�^θ��z3��	5�m��$"�rdP�Ԍ���R9ށ��N��3@I<�����je��T�WdO�7f��3@I<��������E�9�xD)�woU��|��WH@�'�{��}�F�)�*��:���G&8���m���sx� I;�P�]�EQQuw{�y�f��3@Vpz�ށﴴ�Q�"1�b�s�+i�'K{d��/")�i�F��8�Z���F,NC�{�� ��8�m�@�l� �Q�d&��*�0��������`��4�QW$�'��)' �������;��hI��B�,*�jfb������`��4��>�G�&���=�TҲ&19<b���x� i;�;�{�>v��s�vh�����3R���v.O6��w�ri{7lo��L��S����F�0'xsot�ـw6�4-A87 ۀ�8��޶��[��޶�:n��6�j�`c��,0�^��f����Ӽ��� �X�G�FO�jC�{���@-�8�m�@�e8Z��!0����`U��h���w6�@m[0����/{��_~����t���  �U��y��sU]�h��7V���v����݈󝗜=�8���:�1&�d3������u���`�F{z퉳$�;Z�g낮mX�+��3�Al��!1%�ێq�NXt�
˒u&��Ŷ,K�=�p�Gk<;��	��Ie�����XD&�s;��2:j[�.���4+��v�O=v�B��vuTn��-��,��"I$�5��q���7Hy�<���ª��K��(F�5f�KTR��������om��6���y����AV8�,�5#���Jd���/���Ϳx·52��$�4�8�m�tv�8����[�����+	$��!9��O# �M���0soc@R�86�6�'�ng ����vS�~����׋ ��⦤��*�k�NJڷd�u�N��/!n�Ad�6���.K
f;DԊ�Z�j��T�P���߀�w��m�h���w&�@eE;�����ۙ���U����`�����)�����@|����;����䨪��#@N������ �;{���*�D��y1�䤜��{�;f������އ,%�WV�J5�����=�os�]�������o�QőIF9f$��۝uٝ�>�n��z{\5�7��#�^�g&D���I�I ���΁}���=�oz�ڸ빨N�G�bNw:��0����9�;�{��q��2I1��ng �����j��Ŀz��:�ڸ��ŗ$�7�a�w~���8��<���%
N���x��-W]�M�%����� ���g��{W ����\F���}{v㫰�����d:H�x�{V*�(��9R��958����� <l'8t������9�=�c4JG92]�wR_�PL���M��[0sX΁|����P��8�K'�Rw�^V���3@s���M��C�������x�"��w��{k����V�nSa����Z��g*��j��LpI��xt
���~�{�/���?z�)���o+��JcPM��4;Oj=s���'�p[r��{v��c���t0$G��y"��~�{�/�9�=�c4<�`	�)����qU(E�߼���r�>�yǀ��Հ}�m�@.T��dR<2c�.��yM�'Xy7��Np='*w5��
U@U�a��OV��~}���p޻�tn���H9'��)�M��[0ɽ��'X����JZ �7s��fJ�PWL��)hu���J�L�)����c��M/8��t��-ZF��� J��a(+�廍!)�yx�pY�h(�h���IH!�e@rJd�B�!$�CT�b9[�D�SG��Q�g�6h��!:yϼ1-p6�EUA�#=_I(}SH���xC�%-42�c~�"Sb�`�&�(H��44�XTC`⤌0dScAcT�fT`8���AUS���S`8��4���/�����M�T% ERKV��+2b+ɚ!�?%�@F	kV���f�kZ��    m�  ��82��     A�     ����*�[ �UЃkÙPl�k$��ٵ��laݳR�i버�t�5M!hU����ԛ���z^�U�Kd�L��،��Hw[{9��L��Mn����凳�r��P��y�6�t�;T�J��{�Oc��4��[�j2�÷k�g���L�[�L���K�m�h��S<E]��rv�ۇhU�C:نj�y�5��(��^��+�j��
N�塺�!�][@c�R�2U �q�v�./V�Zٙ��� �M�.N�f�Ͷ�8	W���)[$�g�N�˦��y/KN ��d״��Bb��V�b������I,�ȗaۤݵ��YU�� p�nny�slKP /%Sɻnu%q�*�)s������a��F*Rm�j @n;vۮP��lvf�rZz��W�K2�`ZIN�l�r��P��+��*����P7k�*�#�oIZ�|Ē�q�Y8D���t��T��l<YL�y��R�Uk��q�j�Ug�J�n�:DxaE�Z�C�*�5]�m��c�ڦ r���r�M��#�7Y:  *����0���'m�iU674»{mΠ!6����<��4��c�
ٝ�m�*�v��^=��i�T�a��MV1UF�[<��ȽYH�=��gp�<@��S�T�rf�k�Yv�l�9N9�j��Ԑ��uQ�������$�&ڀvZ�F�ˬ��T�Iei�nɻn��@�����u�z!��p"�^�ӆZU�Z�sK��**�\�$ڂ�o]r1�ґ�t1J�U]\�-RGJ��5����v�$[I  ��*��n^T���Km6�ɃU\=h�)#�D�����i�bz���knڧ�@}
�G�M��( �kjN���kqS�b�%^\�\�lb�0�ۖ�.=g=t]0/-NsYɺE5���v��:���u�-E��n�G�N)�>}��Ͻ�=�w��q��*��&]�� 6���^�6�m���vmA^m�s��@nמq���k���񬝸㢐y����cp&6V���Z��lT�KN��i^P-e;e׫�:{�f{c�*�;nܬ:ۭݺ�0x:x
��T�Ep�ss�=N�K!R�i�mEɐ� Up�u�G���*��N�^t�T��!�$A2�	�źc-�@W���,���,L�N�}M���6Um�'���a�\�t���l=�����<��h�s�i��q��1����y�}��:[���m�@�qѤ�F�Nb��I��roc@r���7���0�tI;�I&(�s��*ݯ�y��@�o# \��������.�⦢�n� �M��F �7��zw]`kZ�5wJ�\�W~��^,roc@�� �M���G�P�T������kMm'����6{�f��t�W:���t��qK�5ق��w���?�͍�Ӭ�7���0='*�4�Wv��w��?�\ㄒ�	Z�-�������l�7�o�ܢ""ɯ��2f���j�L���s�����8�m�t�p�
�r(�?����x:�ל`_w��V��?=w���I܍8�<!�7�os�>�� �M��[0܊���ueBm{m��k��-��7�{!�f��ۃvCn�r?���$�"rX�
w�@�{g ���� ��sЗ�>�yǀs���܄�cO�$\߶�����w���j�}���'�CyG'z��0sX�/�+n�Rs�w4�@7]P��J
��UDլ�IO���x�O�p�ot��`zNUC�����b�
��4Ԝ�������=뼧@2ԫV&(�hjD�0�`�陶�lkn!��:�x�OX��6��_��?l�
Lr4O�Ĕ��o���ށ|�\����ڸaCk��M<QIހ�����3@j������"d��T�r����MM �� ��x��p��߻�������0�j쫱\����7�h�9�;ͽ�;f�}1�+��JSt���t� ��U]�wj���w8y���l�;��h�9�?��>�x5/��<�4��5�fI9fL�f��#R*mf�E�s���bw\�ͮ.玺����� ����k��# �k�s�� ��ozv�w�La�� ����Q2oS��7����ߛŀ9�>���HL������=^��=��ށ����=뼧@�Ck\JFH�>L�����sysX��'8����p��x�s�}o3�{�yO*����ʽ����*�(�})w��4�v�L  n�k�\��n�R�a�z��Mqpp�z���v�盧E�n�Z���i�Sم]p����5�b�)\�n�%�O����[��ƥ�7A�T�s�g{E��*��N��M=1����)���%�'Oc=���SV����ֺ���ƣ;��*N�10p�i�ӑ�f�;=D�1z�4v��A�9�i��+�qΏ����l~p���[���.�XV��.�Y�{a�F����.�
n���.{jܝY�27��WIc4t����������߽A;��I(�;àz���Ͼ�Ro��� �����6wD;�UWs5w�Yws�w�{�.o#��<�� �I� �B�*�*ff������F��3@�I���� Ӫ�WDV\MWIc4�I������g �~��+PQ��qɐ0m4AnqY/R��p�c���f�*�6�{q���������iZ�T7y���ֹ�=��x��\����5��x�T��ګ���h����56�@|�F�,f�Γ��7�B��J��$��.��t��`��h^��;���ێ�'r44�&����,f��'8�����������$2(�S���.���wm����8�w���cv4�<nD �ku�jL�:�s��m綒�#q�or���$��2&`�x��Ra'�H�v�ށ}o3�{wyN�u�\�f�,&(�m�B���x�x��B�5��xt�pko��
"T�}U�*�WBYjh���ko8�:�8L%iD$��#3����o3��ڞV�Bdō�Rs�@j��Sot��`��h`�OydS�Ĕ��wn���y����:׵p�
��5��!����)���;.I݃N- ��s$v�Wn:�1�q�hp�F<bs���g ۷��^��-�{�?n:4���Ә�xV���=�B�9���;�w���Y�(S#��f�U���L�ڙ�a�9���������׌�;�*ǉ86�$�I �m�@����-׌�r�BBQ���^}8w'(j�)����w�_[���S�]{W �{�=�����0MXԪt�Џf���ݛk���p������u�F-KF&�6a���=��S�]{W ����y�9MC����b�
��4�9�54�@|�F˖3#�Q	D��ꜙ�ut\�U3w8�Ͻ���Ò��νyǀ�O� ��'�Z$?�H��@����7}��@{Z��%��s��櫊��Ss55j�j�� K�3@j��[Ot��}$�������������&����� ��&��\�ֳ�8��x��L�rF��W���/F�ey�vӍ�i����L�%��#x����
ޭp��g:6vi�3ķ���l�&;��L��/�����V�[�DUz�L��Smd�I�˝�Ƴ0rn�E=�O%������]o!��`�T�`	��l+ِ��5g��&N��A�fUڻxqn�'�2l~��_��h��`ul�����
�9|��ù��[��ɸ�D�s��j���UQ3rM���wW9�<޿x�x����:��c��I��9"��^�������� N:�.�"i�0�#����8﷔�^��;n��v�M�O�&&73�j���� ����y �r�t��)�6��:׵p۷���g ����� Q�5�ɀ���a����������LcV��t
�EkOρ���DS�Ĕ��vݽ���`�n3�K�:}8>�*˲f�R���x�x��(IyBI/Е٫s�yRs�ki���d�7155tQPW\��T��A����y�{q'q�ri�Q
w�@��������0�c4)S�������껹�54�@|�F˖3@����E~l�4܂��(��ɒ�3c�D�usH\9R���[��\��v��7���~Ȍ�����s�_[���o)�.���m�{���171?�p�����^3�	J��>��s�x�x���X`�����.���m��<����	��B�,
HI����P��K+����k8�&��_62SS̳愣��K� ��	��� �"�
���	f�J��($�dD���q1`0��N��zx��z(������	(��Y���7�?0�V]�E��Q37s�i��7��6�3@j����R�С �x��z��������t�pk�����vtT3�<�a-Ʈ�f6����&lt��j��ì��z@�(f!�kr�w�o�r�hRs�&�ߴ��`���c��Ǌ���.���[���_[����:`j�0v<M���9�N �ot��`����� N;5��D�ra��;�2��g �o)�]�_w9\Tx� >�"	��4��}��߼�����k[5�5pQUq�&�3@j��4���ŀrJ">�8�*��]Ģf�J�Xnd�u�o7\���y��8졍p��^���O�9�~fWj�*�*�0�:}8z߼��g �o)�?P�>�&6$�\4�� ���4�T���khP�K���@����6��:�j�v��n:�Qci�1�7q�&�3@j��4��G�7��o��Vc�$�c��xtWj���B��>�߀o��^3�tBIu4?�K*mt ��]���#-�uQ��-���my
��t`��%���ݵk��׃{C��V10�ݕ���b��8&9�s����1,�� Wl˂���Tp͓�]vqi�N6M�݉k;u8��W<D�Z�%ю�Ջ�ثXN�쌀�c���\tK�������T�M�f8s������뭩�uYǈ�z4;nǣ��H��w{w���=�/|ܖ	��1����>GC���fm��$��8�v��ƼO+�kC��{��g��aJ*�W8﻽�7[ŀk׌�:mp���N��4�ra�';�7m�pz��M��[���JC�������
��(���>}�x��������8�6���L�`�1��>����M��yi�40�>�ɍc��$��v����o3�m��t���7=kuȠI$nb�v��v�va�m���'.���u=(�㧝m:vs���0D��BA,?�s����o)�.�W ۶��{]i�����Ҫ��X�x�l(���P�c�����.������)"Cm(�;à5M� �ot�>�i��4��لq�N&ԃ�㋀m�{�.���v�3��p���N��4�rAsW�M�`����� m7��*Ѷ���☜1|�A�$��C ��\çZ�{�����g',h�L���}��Z�*�`��x����~IDx��8|mMU����xc��:T����@i����}�
��)2cX�lI8��oz�y�;�%n�t�]��w�����M^�4�F �x��np6���ZC�7�n|�6���7v��np����z�,�BI~��M)����ݺ6`�͘�n��g��׏:��rׅ��;��_p}�t�eql_}����u��8�ot���9'���AN�&�ڑ��.�m��`]���=�yN�uڸ��n'rbbra�w@i���x�>��� �m�.��mLo�	���7v��r���{��8M�S�6����}9Ui�M�Ƞ<krs�@��\ �>�6�h7��$�3@!�	�I7T^�k��礭lv�ɭ���zq�;G��݌���:����W�*�h��کUD��π�����x��x��D%��p�#��T�N`����;�.����yN�uڸ����şf|�TRX�����T�W%�m�`	77#���cO�à]v����m�p>�>�}�����
F�$S..�� �M��y��t��#����?��\��   �Y���g�&�[�8���2��Ergv6�ע)hn<^��\����qR����������I�v� ����Z�{��jH��lg��������ku���6�Vmm��O�m�Cn��A���sl�z�2k���Yv������۲w&�]����n���vF�����!8����O@��Ϙ��C�a;7<�Ԛ���g���������Wm�`�)���N��,�k��\��,��h�-�7����>��G}�p��6���I����8�o)�-v�������1O�p&�3�.O�7M�����2>�����I��	�a�Np��W �u�x�P�y�b���<�̻�M��J������J�(���{�v�b�7�yN�u�\����ڍI�S�u{�>o# \�3@j���7�O�ݱ�&�g�-�[{5�b�.�4,���a���������c��:{�����3�/9oꨪ���rx��Npɽ�W��.ۉ\�b�%��<��kڳ��%*('_w�ov,���6[b���������oz�y��o)�-{W ۞���L@ڒLx�/��$�DLD/���>����q�7k\��oz�^\����<�m������%	�}8k�����ŀz6��Z����5�����1���&�IҲ�N�j�]��cQ>Ns]?�Z��k��UU�a�%M� �7�6�0��:��$1���ƒN.}�����6�0��4���7�1:����D��j����,���ЮƜ�T�Up�Ⱥ4�����D�0i ��&Әb� �9�)�D��?/��]��w����i�3Nn�QUt*TL�� �<f��'8���m�`�RVc�%�4D'�u�\��	L$�v����� �k�x��;e��c��Z��5d�ӹ��d̀t�-���Gv.'�L۴ɖ�m����>I���F ��3ﾏ���� ۞���D`ڒLx��z�o3�_�q�v����{�A��EO)�+���`��ǀݭs��$~{��������i+�,�rs�@ߵ�s�~��w�*����+�Qx�q�}��d�r�t6��ȈLI�����6�@�o# �3@J��Z�����-�oGX��C�,Bd뗣'/i��&շc�Wv�F�2�g2���^}��t6�0i�4�9Ͼ���sw��J��ӈǏ��뷔�	Rs�.m���F}}�ә��)"X�DB}��7^��7�����g ���t
��Ɔ�&I�q`�{�y���sO�G�}|�'8��n7r3Ԓc�7;�?[y��^3�nֹ�7�߼�G���	H��)�I+�1�Ƣ���BhjX&RB �H�YB"�U8T�rִ�	��g�	�BS�M�@.��&XK`��AAt��&����?��P�P��%bH!Q"t `��B�	�% ̩��۰6�T�F�������Cf�oZ޵�    `E  H�mq���          
��w	+z�=��1���F*j��y�bp ������X�pE�eg3QsU!hU�T��\FB�,�H��d�Hz;U�n��oF��8��oa�1-v�Ds�Q�
q�̓k�8R1tp5�;n˃(1��ݨlpm�̭z0�zL�-3��ƹ�]K�Pq6��}i`�0.���-��7�n(�7g�-�6�+2�nC]�G-���C�N(�*��etN1�q8v�l3Wm��TyBT���  uMUUjIy��gP�8���v�����Fz�1`I���bU�6%{r7UUm�y^ZMz)�m�[@F�\�$K,M��.�#m�� *��&�w.�,��KnIֹٹd�N�mk�[3,<&�{k�������v	��jv!W��ZЖwam�lb�����Ӽr���m@,�`� �]mb���ʶ����-n��R�v�=�[jg9d�ñ&:6��k�%�*g��ukZ��G����^0s(M�Z�Vԑ*�DO2�dԔ:���2����J�3i�_[�:Z�H^n��	N�ʅn]�*_<�bՠh�` !RTӵ�:lm�h�3�5k�z�O[��X�z:���P�'��QV=��ycy�9��:�ݩ��g`*���6�P�G�(D j�ۧsI���\�UV�vcbՌt�@�ېS<\�UU��N,��Q-+*�W��(1�<+�K-�pBޚI-��Y��'�{q����lj��������J�R�*�@T�0��Bb���i��eUEQ�@�lLi�t�!���n���$�]M���v�-��  �v�՛rmm�� �V������3��R���K)Z��l��MO �ɺ��I���p�(u�klv*�T b�eZ:���v�\>9�2�g;a��h�,jX�Y�m��n�f:Mt -�K/��j��Z^�Z5�ݭo� $(lG��)��� P���T�P�辊��>
 �.�}���Y�f��L ������M�h6j�[!/����� ��\h��a��F�7m`�8�9�Y�f��qga��-;�Ųmrpl����v�ϴ�#ћ/l뺰�4��W[�>�1�0N]����Nݦ���y������qq�z�s�g�8��%͕�:�p��� J�Nsa���ifH�n�R�;=��2�T�}��z˶��<ч;��*�N��m�Pv_ؗN��ˬV6<��$(dK���8D ۙ��ה�	Rs�.m����Dhm�`G	�I6,#0YNp��j��oz��8��S���}���Hd��ěS7s�.m��y4�t����k��������*�����,y�q���B�F�����,���ꨡ�cǈng ���t]��o�������n�`��RdBd� M���0Z�r���"��uc�l{u���s�p7�w�̎bR4�@O�:���7������=!��8�Ow����˥tV�Z�r���{��ҌI��Sz�����q��nr! _-T�ڒLy�z��8ݼ�@�ڸ��� ڳq;�3(Di��u�4��6�@�>�������b�0G�I��j����m�p�yN��ԁF�`�jd&��XeCX��粌��Iyx�L�,r�\��Ͼ|s�C&&�CI) ����6�F �x��np�N���j.&o�����o# i<f��78�W�3�J�x�����p��[ʻ�w��_6. ����w�*�v�8��J��i�0o	�}��-m��w_�m���D�o����rrbrcq��I ����ݼ����t^��.�_�;�7 ��%�\n͂�֎�'�a-m�\��sF�䰦c����ݹ�bg!2��Lx���� ���<u�y%������\��L�J�.@��� Ԟ3@n���'�j�9��e�Ьa�ȱ�9àZӜ�'�i�`��h�������CI' ����ݔ��6���37>��T�p��M��a0�,*��@m[0N۝�NpI=�76���s�"8��yL#Y�V-�6q��z3`�Pܻx3
�C�*��(��1���Wf��s�7I��'�F�ڶp۸���N��qt^���2ko��;��{]�>!�m�]\�$��
�pn��@�e83���}}��;����T�츺�Wwj��_��S����� �k�Gۺ���.'q)���mHp햮��"!$����m��{l�&�"��Pr�C	=~�����E	��  ��i{n�	�	Ҳ�vJgR_������lZ��ιú�����#���8A;(t�'b�Fۃ��h��gz�
�!%�(���LܶlfƷa�5=v��v�c9Cu�C���v{�(Uu)'c��k�x�q�Y	ƛ�FFcE�n��,����n�)��1���<L��MCc.��m��ۇ���-۸ٲu�.�G�����K��s��:�v�ѹt��,k��@��/GA��`z��^���/Ϗ��Ӵ��GS}d�?EO���Otճ#�S��@�x��I&�I8��v��[���e��Z�\��M����(*��@m�0N۝#npI>�ʉ,�&�!� ��j��s�rI���6�|�]�tMXҹ
�����?��[}���Àwl�t/��+1�%̍ �����\E����7=n�����m���9�v^��;b�d�a$�G�@�.�ݽ�� ��jϳ�Z��m7��md�e)��x�ٝ�� P�	D%T~}}��;�zp�u���54��ĩ��
��0N۝�Np>�����l��|�%d�&"�������rI�ڶ`��:0o&�ꫲ%���N.�ݽ�}�_YNݲ��.���\�[�%$���b�G����M�Y�Jr��޺�K�5��p�F�<���Q���x�''z����-]�ڸ�v��yQ%���1�!�MHpk��ܔDD�IΟN����;f��qX8��<�g@������yxpC�"?��� M�������p�z?��?+��L$��I>��9$�@|��m΀�'8��iܟH�I&87;�/�� �e��]�Nv�ށ�E�mc1e�S���AS��;���vN�G��b�rrƍ>�3��k&7��b� �8�-]�l�m���0�N\��
��W*�/'�=�f|��A�� ~��u�Y�gؑ�-���A4�S3Uf �����ـ=v���l�=�r�UEMU)-QH��x:$��$�.��0}}����HP�	%� .C���y��U�v����5�D�!�MHp�Z�ݔ�m���l�:��>'�Ҟ�.ʢm!\����l�^k�V�[vw!�k^���8t���>և��J�)�*蚱R�
���7ذ����)�.�j��ۆI&L��P��.�{�/�� �e��]׋""!$�m���Z�e�+��VU_��ـ4��V����s��� ����l�t�����HP�(���X���̹�
���������'��6���yvZ��}�o$�B���)$�I$����nn���Wn�;���(G�cu��8�ە[^���N�q�̋�+�3��K��04-�6B`����cuΪ��/�Ls��u�>gۛ�.*�����dk'����q=vlۮHj��N��ѹ]<cW!َӰ�r��'8c��#��6��LR�]�%�D�Rd6��,�Rΰv6.{_�C�g��v��w~�w]!'��sx�n�$�{Yki�J���6�ݮi;t��ֺ��t�G���}� ��X��6�i	ɞ����]��y��m�B�	x��X�NXꨩ��RTQQ3W���0ݷ:��0���YlM�$InC�[e������J!����ŀn�Ը8���0}�]�o3�[m�@�����j�Wn$�I2
4�'k m���%J]��������8��vI �b�5�1&F7mM��ɐ�&�N�0Gl9B���,��i�i�I�4�zݼ�m���}o3�[m�@6��N�M`�@'3�w��{�o͂��"��`�?�25���&��F4��UMx >Z�{Õ{�{�<���r���<R�&��ʫ�����ذ�~�u��v��a����!�6�HRL�g���{�.��pl�t�y��ʩ[c�Ɂ1�����0ݷ:��0�{�t����o�x��ƻ�ja0Vnn-�y�n-*ۆ��v�s����ڱ���{���`;�y�Ěs8�Z��y��oz�y�v��`��y>�.�v�,�߼��`�n|B���B��$���'3�[m�@�o3�2fg���`2HH��$\�\ڗ�����4��L��B@@,�	3 C�t��h,��x~��hk	1�42�_ʏS�h<`��y�U���
��	������ˠ]���6��o.<dM�દ���x�ݷ>�x��o� ݯ.G0S�L1��pl�t[ŀ6���m�X/ѣL]Sd�Tۍf����;���'m؝vۖ4�{P��n���;���e��MT�sUQr�k3'��ذ�~�[Ő�m�s�5�ee�)�#i4�$�m����m���v�g ﲪV�Ԓb1�Nw�4�F ۶�@i������L�n�Qh�4�jj�D(S���>�w3�[m�A���8�n+�0���+o'@i��$��7��kv��Z۰m�H�_g���7�5d�ӝ�w#ke^h�/v��]m�7���� �&ʛ	��$��7��kv��m�p�7ˏ$���m�Ι?w_t�}ذ��� n�M]Z� �i����W@�o3�n�����8t˸�W�F��<��]��0�{�4�F��s�&�Y*�f�UT�wk ��~��%�>�/�����=o��D(!BA�4PH+�c�AM�B!*`���w��{�*[d�  ݮ��m�3k9՛�ת�ܵ���[n�#lA6F�H=\�k��s��$  ֨19.���m��8�Bт��2�b��uv<͵����� ���[�p��{y��ˬl�L�\��z�N�K3�fR�ڤ�v9�X*V1v��_U���-u�u��u8y޻]2F`�;�'�[u���I�e�m�;H�R6F�]fŊX��{�������w���������G�q����ְR	�"Ηp�@�p����c��nN֊ܴ.�,K���RR��j�tݽ� �v���������K-��C	�Ěs8�m΀�yI=�o# o�Ļbp�#�C���v�8���L�y���W@���2IH��D�0�{�>o# ���o# L��yq�"c�bBs����e�@i<�$���6MTeY?Q]�-T����m��9wcD:Y�����X�9����lD�L�dm`�L1�!�;l�t
���I���0���u$��iލ��g�w�Ú8,(H����� ,*�J�G�D�$����`ݷ:�t;�"�)�&)&p��ށv�p��ﾈU_���|>x�|��]Q3wv����j�t�v�[��@i��$�z�D�[mC"�5!�/�-]��0�{�4���S�f�.k�������'{GnE9������C���ܦ���}_l}fp۷M��� ��X��� ��9(�}��>����2II�J"s8��ށ}e8�e��]��ϰJn7��1B�T�W� ��0��s�J!,BJ P�/[ŀ6���7]&��B��EM]���@i�����;f ]2�+B#k谏���m�p%	��� ��0��s�9�2�=n��v�E��+��x�q��ӢNSle��՗��j��� �������;f ���o# ޅ,�LJI1�rw�]���>�0��W@����.���*�2؛�}<I�ـ?;nt���I���0ޢ]�tM+ud��^O��I$�^,��}�|�����z��� ai`O�P��y�sʿwWawqR\�V�����J#����u�� �^,2Z*jJ)���vCN��ϖj�h�;/6�<M�����g%�3�����{���/�-�-\�o�6ϝ� ~v��'��&�� Na�YY>l$�9�ͫ�]���}����p�P�ZD��a'�{�����Q	$�l�5��x�n,�$�1�93�m�{�/;f �x���0�)d������)UI3W� �v� JBZ��<�|��m�@y�g�f_��$�I��Hp h�7nDٴ��Pyu�x���h��&�O=�p�B*���Ӹ�ZDr��t#P�����d�k�+7R��i�LX��S;���2q�:��A�ʆZ���϶vu'Q�nT�F�H���t۫���s�6���k��1���6�ۭ��wOb7N�iw݁��nT]=���=��zP�i�=��]s#:�V�v�SFl�TD��+���{�߾�^��~_�M�b0s�<��vi�#�&�ӶԧVsu�RI�!42� ��74<Fn�vߟ�{8�u��5�~���`��2쫢j..��3^��=׋""!(^�� �o�^3�~zЫ�]�T�ՅU� �ot��`	���O# t�q�Ę��r';�/��p�x� �^,	%׭���:):.*���`��� M<f��yi��/��p�V��8cmߔ�<1��,MtOIu�=x{)k��^�сti.;OF�.��g�����.�0�O# M7���9��}��`v�|�,�"�,��U]� �ou��<�F �x���0��TU1)�<m	9ށ}o3�k׌�$��X�o��&�fj���USV�?�"!(�Ͻǀ���m�@����7�q+�� ��MnI�`	��@m<�4�����/�-�gW`:]Z��D�n6m�Y���۷ہ�=s<�����ww�������X]�T�ՅU�^�� ޼X�x˟�]� �n;0n��C�9ހ�\X�b4���M�D}���� �j.WƉ0���p�yN����9z
+) �����u����5�� 7�k������"�w�xz�`��xz�`D%�6��:�QX�FD�6���Myi�4���suN��U-��l��`��V֛n�s��&�8i�uE��69�nG��< yi�4���M���'#�0llng ۷��f}�|	���&��4�0��˲�����&&kp�O# M7�i�`	����hU��.�*Qj�UkB��z߼�x�z��\�DB��}�wj�ª�*ʹ����xz�`	���O# M7�J%U1DL>��w�Q����z���,m{J�xۇ���DIǒC��I�����v�4�0�{G�}�.o# ��TĲ6��	'8t]���m�@�[��v�}QX�GY�Ӗ�z߼��,�!$�z�篙�;�5QTĤM�4�s�}o3�&�3@�F �ot�@7s5WP\EUM\`	���9���&���{���E�}�ϕ����٬ ��ZX�XX0ɢ?��ka��x��	G�2N\6��̀|���W�8	����H�r�݂z�����A�&�c������!��)*��4&�LH)�--Af+.Fcc\�Ĵ��d��)�'��Mz��|�UXT�} ׈F�D/v~J~F݂$��`����A`J��{��w�om� R���  E��H�Z� �          uTX�G<��iSZͰ�jb��
��xz���l)-r����e�ef*
����oY��҇�:]כ]sH��f�����$NĆ��[KlKwI�I�C�3�n�b;Bk��ʜ���q֘�(tT�mT��ڙʦm^2�lQ�`���>��1A�`5�H��L	t�"�X���e{Nt���7f��mб�6zm�.�,tV�x�z�V�U�*y���X{%�rOH�Kil��K�M�!�5;!gCC�j�l�)�7��	zX1�*�ɔyH�F4�N&�D���j4osnUiH@����'��)SJNl��0?�~��ҥ���l�ᥝ�HƤ��������v3�Ճ�|��E�)e��*[u�΃���l���6R̚y�j0�5q]P,v���}��m��N��+�̰s`�:�ٙn���p�U�F���.�0 8�[!U���y\f�@PUfe�Il�Ȭ�cv+i�K����I�ƩF�k����DOg�2� :�&�������q&�58�+'d  �Ҭ�3/,7���A3�k�S�=[��]��4��@�r�݆�  ;A�o:ۦ�B��dyC�JL��ZRZ媁ݸ.�е�(��R�e�<�!��虯Q�o�v��d�k��<��C�J�������n�P�R�n]�凱�HA���ҭUV�"N�H�5mU���h�v܎Uy^U�[m.����yT�y���luOl��@�֤��;��1e�%Z�V�j�I��
E]f����j�U5�Nx�כ�tlUa�mR��C�	=�A��U>�v �>��+�  �v���M��b�UP�	���7K}}�h�5���`*�V]�	�P9W�z��O'mkl�\�s�ġk�V� D��v�U��Cmr��bت)ɭ��T���z/'k�̼쑊����qK,�Z9�k5�ֳ3y����z	�� x�Ȣ��^ ���󠮅O�����O�Q��}���>  0,:�nVJ�EWn�lء{�g�Ѩ�$,cv�7/k�ݸB�x5���4�8�d�-b�� �9ʆs�+&����3�!�g�L)kP��mE:��ʰ��@�n7��@��<�N��&Cc��-3m�&��ԡn�Խp��m��v7��}T�� U[&���<3�p�S5�D�]�Doi{׏\v�㲁V�߽���}�w7�����՗N����m�9�5��\o<Wn�����w�hw���{����>�j����S5�h�{�[��ߛ��6��:���#$���p�����%#��X|�8�=x�B��� ��q��H�lNw�o��p�^3�DD�7ذ���])j��dMU�_TL�\`��4���$��DB����, z'�T��e\���.�0�u��:Q��~�s�X��)��KlpB�s�GF�<ݻM�\ɱ�����ۥ�phn�;�������F\��h��(���x����x��^3�[���;�
Z����&�NN���g�CP�BN�(P�9�g��X�u�ܡ$�L�'J몪�U!TUV���q�׋ n�x����S.ʺ&����S5�<�%(]ϼ�����x��^3�~m��WE���s3aUq�>I��y�x��������c�`�1��5�Ě�5�l��(�V���%�s`Ǳ��U�.(�Ƴ�l�e���TM^����?'��O#>����ށ���̆7&&c�ۙ���h���>I��y �IR2��>������0�=�ɔb@OR2P(J�9�)/3�w��S�{���ds������"�Ok}��� �k�xv�8aKS�<Cō����0��i�`�{�zX��~�Ş��wi�kp1��:ǆ����ܔb�>]s�l+���w��|v�}"�&˗-�x���0�=�O# ��2ګ�j..����a�׋:d�o��;�b��x���"�]w%�ͅU� �'�i�`}?'��O# l�U;
�,���UW�Os�,�}�x����P�MDB�>���S���b��SB�5Uk ��<Cz�`v��v�8~�Qģj4��5;��g�;n��V�%Mh=�f�k�<���G�fJ̒���
n,�����7��[���0��h�GEe�]\7EU]� �ot���O�6�G>� ��)�0r6�x��s�ݔ�	���O# M7�*�0�*B���� M<f��yi��-����q+q�'��8/�}��-�ŀ	k���7��^3�dD$�m~?�M�Ke�  ��I���P<CQ��N���	G7e����h�C���	f��37b��q��Pr%���.����i��%М'Y���d}URM�ѹ3�#�K�������$O+�.�.��K�zs��9h�]���3�6l;���؆��am�=��ޞ �{?O=��l���]�<�INy.6��t	hݟ0�hv�f�[,#35�[7ov�UY| ��;}��4Tpv��x��"S��Pݮ�n�XI�<[Z��/��ϊ�ݛ�U�Ѧ䪵�w����ŀk׌��ŀZi����BID�z�y��5��x���5�~��KT��Uܕ1Q5Uq�&�3@m<�4����p}�TJ<kS!�I9à[�# M7�i�`	���;���˘RbJ1�nL�v��v�8ݼ�@�o3�v�@�Ԙ�'1��*8Bp��<q;��m�k���5���w@"+9�u���c��cŃBs�n�g ۷��v�8ݷ���X��&$��k ׯ��$�/�B��_b�>�x�y���+q�'��8/�}��6���Myi�4&�+"�}����n�ށ�o3�m��t�y��M���H�r';�O# M<f��yi��=ng��9���+v.�9�;%�׋E�:5�'b+���X⽞z�ܴd�n0��h	���&�ߣ@M<� �yf�PkS!�I9àm���u��O# M<f�ܤte�w7U4IUv�z߼�x��t%	@�
!��e,�S$�
<����������`�Zꊻ�RR����x�O# ^i�h	���s��@�R���"�cm�����t�y���{�6��p�n�`�����P�
p���`�\N����0Mɧn6�ܥ����#�\�8���G�}�΁�o3�z�^�	���/4�4&�+"軿�K��f�� ��y�Oc@M<����4�$X9��v�8�����	���s��@N�]@��.�¦**��0�ƀ�y>Ot/�E"/dr��*�߻�ӕ]�f�Ph2$�tn�g ���x��,=~^��J;��NuX�1:Ik�r���tD�9-����dk&�If��K[��l�综�}[��
��]�/��7@�o# ^i�h����d'TU�TIQ!A5{�y7��/4�4n�g ����k�b�N,HUq�/4�4I�`G��=�<���/�%n8���G�}�΁�����׺�y�Oc@�&AYE]�us3u3Uq�s��@�o# ^i�h��ʺw�?�������1����޷��������k��` *�Gj�Me�q�L�s���Hڀ��<��s=,h �/S��s�pK7Z���X#�β%r'�gF
���zCe��*�����z�+0!�f�7m��X���7�g�@Ӻ��c���}���:]Ym��f�.�����ȵѽ������wF�{-@u��/+˹2�6���e��xא�i7ks���=��pſ�9��r�:�j׆�o[�l̶���/1=u��v��mmŢ�p�k�0Xs�v��Vv[U4���QWsW���ŀo���}�y���{�6�U�gЎǃng ��_����Mo�`��{�~��dDB�z�$���h�s:�o3�?s{�y7��>��4�GF]�5e��ԒU]� �����F �������u�����>�*�IJB��߼��0#���'��&�F ������_�7��b�a�nzv�4�`d�M�:�K.���z��8��e:�܃N�v�*��4��0\�0�Y�r呀{vI�4ɨ��W1sW��5�ş�!F�����w�;�<��~�U�}��:}������#�GQ���s{�&�F ����O# ��
�<�9"��9ށ�o3�_{os�m������@��W��B8Lk6�� ����>�>��4�0�ot��������*;�����l����OIuټ��08��w��xն�xz��>g��<l]R]�F��y�7�i�`�=΁�TVrC�4nL����@o^,�׌��Ő�(�=�Zꊻ�RR��5w� ޼X����EG�G�C����Rp%�$�1#d�03+	�"�0"����G�!�
1:�	) ����oc0 ����L�$`���B'��8���X��SA�O���I,�C)4C$�� e,��S))&#A��,��4TD�L d�BDQA�jJ�"�Đ��`��	 ����l[%�Čeh0�$��F�&��*�'	hC!�i�����|�%8�"V���(�B�i�$�p%�0g`��&4�FF*X,�	~�k�w� �8��(��`�(��
�`'�"(x�ȁ��E$<����U?
���o��Õ}����*��v*f��4XJ*���X�{����w>ŀ_n��v�8wP��1?�A�	� ޼X �$��u�o^,�ה�_Q�N��%&D�F(ܑIJ^\L��v��u�w87m�sm�y�kC����z8��&�p�oz�y�n�S�[���6��ƞI�`�Nw�[�� ׯ�׋ ׭��)DB���UH�.�+�S5Uk s�/ ޼X��{�-�����TIA��c����ŀ}�����,�!��"�z���zN�.�5b���$��Xۺ�@�>���y��ƀ�yG%U��,S:���z��J�ӆ�s�^]��l+jM�V�4Ŕ�69�n��\��6v*�@|�F����4�F�'�'Li;�X�6$��ݶ�:}�g��^,��~���g(��'7$�*蚋VR�VMߗ�����x�x�v���i���'��(�ng �w_���X����舉��\�y`i��o���H�"s���g �����x��u��rQ�ow��]ͮ�  j�n�]t핓���K)J�gʾi��Z�[�1�W"�\noL��q�\( �M��3��i�2��Q�gz�
�!�%�`�s�8	�ð�f������]�ۇe�w`��a�����q:.�I�'���Ψ�M�v�)w5@��d�,]g`�'��wef���j�1̄��MM���fzC�Q��Żw�pu�ۋ����>Nw�9�Lb���Y�].�q����]m�����*DkI)����7�#x�ng�����^�@i<��Ot��`
{����$��V*���<�x�([o���,m���7��������8�߼��XB�S/����s}� �ȦZؤoу�z�������v�8g��oz��N�&@XU5Wm����0�{�>v��Q\Op�$0�b�q%{5˭L����v+ێ�s����htF+��n�Qu�U{I�`	��@|�m��@�L��F7��	D�s8�oz��A_���q\����6���@����6�7�l�9
����;f�'��4�F�����>�rbf4�� ����@��F����l�:_T'1Q73DYSuw��4�F }�y�>v��v�:��Z����ۀ6��Ѡ&� Ƀtgix�=/Z.�d����/�m�e�
j˩*�J���?>���;f��g@����;�)��)�4�9ހ����Oc@i<�Sot���L�����Hě��=����.��p�
D�&}��x�x���N�WDҰ������O# ����yw^g �i��dcy�J4���;m�������F ��F�uN��{:�q���Ѭ���Z�#Ag^e�,�/��KgQ.ˊ8����Y]SM�S~~m�7��ws��r��5��@I�UPY����,�73�{޼����8m����g3�<��0PB#k �o��4�F�����0�yyI�|��hlܙ�;m����8�����D`�$C����������=p�[���9ށ}o3 �D)�M�k�=׋ �6��?K ��=��z�uݧ]0�g]Yz�9b9�1��F8��[qnV½r�<�r"�d��[���F ��F �ot��`)���y���@����-���>o# I,�#�ȅ&E�Ud]%��U��߼��XrS-�� {��ۚ��H��Ȝ�@�o3�n���7~�X�Oww~���������������K# ��K�F �Otv�8ٝ�>����Px��$� ���gnJ[��Tw;nJ{��U���&�R��g��]����@J�r�Vݷ����H���0mm�W7+��x�UN��.-��ح�s��7�-��:M����Xo��ڭ�\�m{7$�t�3��V�H���<��b ,Ṁ8-�q���
] �uV��n��k^CbE�L��9�wK���`�u�;@�Ru�۳�w�{�����m�f	IL�b����Vv�v�����,z��,�^r�8���q0PB#k �o��?b�7w_�z�D/Hs�ŀ}󑱾,qƁ�Crg �n�;�-���[ŀn���" ��h��&�IR"���׋ z�,9D(J&[׋ {o��jb�9&��M��m�`	r��$�@m<�R�[��&�B�W15~^�x�([��� ޼\���F�	ȔRD�6�U���j��\\��7h���3E���bA��%ϊs�]21��dDi73�o�oz�y��x�Q����;y0���������f��w�w�?* �%H�\�#ﾻ{��/%��.I���w]ڵ2�j�� ��X�ۋ(�}�{�-���ye�AA���lo#@m<�rOt���o# ����|x8F��ɜ}�{�-���m�p�o3�wu Wu���<7k@Tqk��W=��Ŝ��6&"3��.Е�bGСN"řTM�R��
E]�o^,��0�d`�{�t�4IN�j
�j�0���呀.I��|���-��Ӏ�Nw:�y�+�~��yo��Bʊ�2d3E2"���� ��ذ�`Պ�V]%��U�~��x����f$��~Xo&�UQwSWb.ɫ��o^,�l�呀6��t2\MV[n9�j�|�Z�[9�nٙ��^:s�m:],W]�H,q^����ܮ�^�]rr+w��� K�F �ot�����1JY$����R��� ޼Y�	L�ϻ���,~�� ��dک��U��*�����7���7��(�z�z�`��:U6]̕"(&����J�}�=v�w�Łm$�J�ԡgUw}��J��못�&�H��X��� �,�������(䪝�5qьF�52>�<t������e.l�;Z��/Z_
ێ�jB�m]Ϸ����<�������D@�� ]
�dcy���pv��v�8�������Q'o&��.�����w5~�ϱ`��,w�ŀ7���nٍ���I2bX�ng>Ͼ��n�8�ۋ o[����/�y`O��x�)�(,L�t�y�[����2��w�ʿ�����*����AUW�?������s���.���U���" ���}h�_���������������/��^����������_������������~��Q������@"������>���������UU���_�DET) ������������� ��D�����F�����������b>���K����?��k���|����a?������@@�TaEI@��HT�	% 	�H@��!BQ"DQ"B�����J �*%
� P�B�@! P�(P�JH0���#$�H�ʌ! H �!!CȐ��@�$� 0��J� ��2)@��	@�� !
,��B�B0��
#"���B"B2
@+(�	(B�3� A̣�����# B�2(�0��H2�J�2 	 ���
����" �# �ʩ(�$�(B0$#B0H�R#H1 �(�(	��� H0��!�H0"��
���	(ª���� �*2� �(�# �B�+�( @�� �H0�B"B2� @0!"H0��(�(��#@B��! J�0���*2���@+(��! �(�@��� B�JB @@����KJ��HJ��B�	(���H��*�*���B�� ����6����G��AUV/������i�+���٧���������G����*����a���������������UUϿ������������Y�g�!UW��EU_��#�������3���������h������|�ϸO�=r�����>��*����������"���|(������r?�����U���U�������/�6??���Љ��G�(�����^�O형���J�����F�?ϛ4?��������?���w���U��_?���?��UU������o?����������e5�������� �s2}pg�    h       �    ( 
p  <�(� �   P    %@RU%(
 �Q    � �"�H(P   �  � U@ TT �(i�S������Z��u�s���{� >�Ɯ�]=y:��[ҷU}� Ҭ��L�� �9���o=�\ ]Wa�{pp�lD�*�� l���r��NM�  �|@�  �� Pͅ�ϥX����QJg��)�AJ;� Δ���)��2�P3��\��M;�gJP8�h(��@ �M�4�H�R��@�)J1M���:(3�4�;�� :S��:14SJBS@Ji�����@ pp
(  U  f� `�ݹA@�������^�^�����G����˥�Ϋnm�ˋ�k}�����R�� W}���w|g�w� =�q��n-v70>�ǹ��� p	:�ru��^{��wy{�7�|>()  JMU �ﰸ���Mt�x��;�9U�P��M��m�=���O�O{ou/��r�-����k��w�vkqwi{�������9q��<��u����������ySɮ�r��m����(�B�� f� y���_6���g&�}� �=9=vۛ����k�qk�p�����=��x�y����&�� �z��y�o']+����>�ޑ� >�ުY�������/v�u,t�  zB�)P  "������)P  "x�T��SP�  '�U$�TUC#����Oj�)P  ԥ4� h�OQ>;��a�����?�jO��>��}���W໿�PUt*"���PU�EAU�*
�EES����Bz��")�D�ˠ�����T-`�X.��YL$��5����/
0�(��X P�|R"�:!@�	��F$
�k
D!)��˃�(�E(�`D�ɩ���5$'��w�޷��QL��@�a�CA�\���1d���ys%���ǅ�Bi �"FVR��� E�,%HCCA����):6s���$��hQ�!<<94�2&�D�w�o8W�7�]�|�ṕ��Wr��B�D��d�:7#����a�V!���P��cL0M��hF�@ E,HbD�"� ���!�/c��� �č�=�Ec��@�X`U���Y��S� 4�`��(a��~yfrM��$!��c 1M�����n۽�s�=����<��2�ŗ33��7箠!Ñ��xp8Ƹ�E��pѼ�<��|y�O8x�<R"T�b��
l @��
���Wp�$�!B$5vp�5vHskF�%.Hi�]�bāL�vB)��;4���M�1 �Jֆ$FJ�<��[��5���ud|Hs��ɒ@����h,�J@dV�d���h�l%a0�T��q�M��$4�H���]#0��#!p�޹.�� �xlٯ9�Y7�����ׇ'7�s��F53[ޞ;>A���f�lֱmY_�����]�gmU���U��=�s���xl�L�-ެ����s�6|#U�K2D�VTוz��_%T��_4p!e,-�\�����)zĞ��0 @��B$�,���H�b#�����%��B%����$$�#W0��ssWT�a/�kla0�Y�#6s�ớ�0��`BrVf�B�i!F"Ń����)�"X!�73���N<e�I3I$5����4�CL/4ˡt`�w���C:!��f�#5��X24ƮCD��5�v��\ьY����#s���� VSa�p���D�E�<"�Hs���^>}'	���1���(�`�J�(|B�b�@�	[�6f�.���s�d�h�M0���!R�S���Ɇ� XSA.,&f���HǂF7�8˚7RZa.s�jg�d޴p�HV� ���>e�0���zss�\4m�3��k<9�60�ho�$惇*ʒ��}��
)��|'��<<5˻�=ǀy������g���x0��b1�v���d�pS��W.7.&�$>b�<��X�����Ď!�߷�5'��
k�qߓ{�����%\&�JH��L.��JS�w�=�cF%A�@��H�P�BFA0B*E
%P�T�p�9�-��q;8l�7J����!�BLw�F��e6itj;$���6^r�p�f�k0ɷ;��4\x)�u\R�F&��`B���FK��vkt�tH) �jBB1`��5V4�X� �$}@�B�`���(H�e��1�|T"4	�s! ��$uy�l�e�r�bB8k��
$?@��'��5��� ���ڡ�^Zp��Y�^p��F��F�2��
��HL5�p<�@��%)M�#^+B��rgx$$#��q�4�><�F��0�{ D�]{�͙��Ţc��+ĀS��h��!L&��i��)�����&ay���M'��1�h}"D#�
J�0�� �`4`�4��CI�����8&�ocLt�NB��<�&�1�nFB6C �ٳ�6�)���8�a��ņ���p��\8NF�R&6p� �%�F��5�D x�B���D!��h���#		 BYv9�x��XRG"P� X�Pt�ҀMƄ&:.����mכ��R>���8xh����8�C��#L	�",
�S@@�E�����8S��R"B50Bu�p��i��M��fdn��<Z��+�!��M>�K {@����D"l0؞��X �0 ��	 �J�A����+���$bB B2!BF�l6�kqu�E�!�<����z.�������b E���sG�������.(ʄ}x�_�Z@9�Z����7Ւ��M5	Nj�jF%+��\ּ��@�YM�R;M�V�P�)�V�� � d!R]M�5e0�����VR�b,I!$X���"A D�H ����$d��[f�+�3Sl�IR]d�HZ�5K�E�!�5)�$D"I)��Sk�F��p�cdHԵ���jCe��$P��&c�F�	$aXL& ������� z�.�Gf�7���({�a�O�
���y��<��|'7��bD�O$d�p11/��H�D<P��ح�# B��#A�H0 @6��`P�[9�4L��K�szc�Ā������Aذj� ��c밮�t&��@�@�`��v �#K���pHIpM&.�80(bhه^���nW�x�E�Za�xp<�L�[1�@�6g$S8&�FG���@����޹�q��x�X�W6�q<`5�o9�8Jd��mLBu�y��vb���t� �р��E�@�la_R.�Q�H�I"S!�������`h0^R�j��<�{�<��/B�)1��ā H@jD��6OJB3[$�d��6T�
9���5	I�,$��`0'�d��#@h$������3[gnnM��#���2z��d`F��bŒ$@$dh�:���H@�C��LJf�ks{=B��a*�K�m��'�h4�ƃ$ � �����mU����=<�\�%	V%B �p�?4�N �S�bB+�bH�%��<�	�$�s�k{O�о1��F�)u���f^kܸ��x�ǀH�(FC��L��v�8�'�q�d<}�oۗ5��&�y ,�
BD D >��J>4Ȗ@��k	n�4�&d�����$l�Jc
���ӷ��F$H��03Q�B�a�K�dd��	f	��	�FJ4鍐�VF8#Xb`�F���&��7���	�t0��h�7% ���E�׀��Di5�@��ard`Ѕ F%*ib��6>�l�P�P�T9�]���M	4��x]��ޘ�_@�Rj�F�l�U�FDy�Z�"#Jc�h�˿�s�}殷�k@ �8              ��      �                                   �                           ?�o��m�� $�	۰�lBA�kn��mm�kX 6ȣ'H�m�p��m� ���G`m�����9���ݔ��-��  6�@  ##nۣ�l�UŭjM�����j�� L[�U��m��]a��Km �p ����L�g-7MW�@�� ˻l ��p-� @  m����[�Hm�������p 9&۱C[[I�[@  ��I�ָ��j�e������HN�i4�J��f����R�j��6	6�m�ͫI�@�z�6� HsY4��&��  �[�n���z����Y�
U+jQ���v��E۷i0�$  �Y/0�a�����߾IV�mi;nd����v-���� �/��k�/Wh m������j@p�� ���C�*NV��%.*�*��(��*��[[l� ��$d��нnz��δ��(4�]�h�:YD�Mqvn�[B� 6��p kc$�m���'@�Zl��[���l��� �-�q&Ͷ m�8m����m�nmf�MnA�@'������m$]$�`M�ev�t�U]/�ڄP��m�Uj�k���r��A��˓O8tU�8�9n��2�Z�ỈeC���]'mn�.��`  ֵ��9�f��\-� �m�6� n�&[m�l )G@ �k [G��� �� �M�  m�N  �K��֧: �bڑ [BE��n  	.PH���r��Ā8$	-�˶��l�� -���%��mmm�8ie۰�l[Ҙ8�ۭ`�!m��l��m��� m�`C��ޣ�H6u�H� m��Y��Yy  ��	���v��mm6ۺ�
���sm'`  �lH �m�.�KjF��l�Vڪ���	��(�P8$ �#�˶����O��Lm�ڐ��f�ؐ[%�lH�.�0 -���M2ܝ6 om�m�l'�I $�-��ְ ���-�M��D�m�Bm:\-��H[@  :u�R@/Z�������^�{     l �ZL �������|zI$   $�n�-�mv��m����6��� �      #mץ����
�k�6�n  m�m�[H0 ���[��f� �  �۶:�m�  pp     �l    ݱn�$����k�{�[d -�[@ڒ��l �       �   ����|l $$y��r郀�H m�M�H �p 춺Y���    s ���  p     m�"�-�  [@ i�oMp7���   �s'v��������۴�Y%�m�cm��p�h�� �[A l�H  zm�d�m첀k	:[r/B���N \�3����  ��@ n�����    [m�˦ͫ`E�$  hp 6� m�n�4�i-.��Nfj�v8����H��yYX$��'U��� �E5�-cm.��N��V�T���mR�'I,��6��;m-� ~O��m��vҮa�ks6���������h���h�m;[s$�h �5v��jۜH� � vٺ�`I�v� 8/[֛v��r@r�`6[J	�Gk��C��ݬ��  ���� �Ӵ���4NSS�Mt��)m�   d�#�q �sc��I�ӟ>�N��|,k{n�`��7+UO,�fې��n��^gF��\*2aـ�m
D��HUR�Un��Jؐ��V���L�ڃaUQ����9�[pX��Q��L�h[@ .���mY� mR��v����gv!,�ԫJ�T�v�l��
m��% �kZY@��"��V�[T�5R [`�I�m�
Ak��-US�0dMcC�^U�L�i`���t�kn� 6�H���vݰ ڶ 9m 6�7�����D�*��M�oNn��l���,�����i6���*wB�<|&�v�\sKQh� $�   �V�[n�m�� �   ��n  f�$`ړ\ m�  !�k=�� � �m��m�� �  �Uoju¬RV���U�6� [v�6��m�2���ěI�	 vհHJp���m�&���@  l� VӠ p  ��@Hm�mm��BC���8mt�	 �N�l � �l��,��5P �-���eP�m��6� H�mmn $���$-�6݁� l	#�h  86�6�.처^;k{� �\M��lfd�8Z�)!Ր��jOT��v�Yy׭��uէ,�&9���:9;^9U��)�I��%�f�P�mz��`݂��U��A���wD�UUS���x�Ǝ�>UHN�m/-vh Xa��� UU��UT���!��mm�R˵��E�[@nղ����j��o�}���9#��Z���  [@ ݶ-��p  m�  �:�$�t �M��WhhlsZ��4��l�n8� h6�    {m�`��Hlp �ii�M�ii7H�&�6ܛPv�u�  8$'m�[@�`��  � H ��@          ���,�m�mm�p�� ��[~�ci6��D����[Am�mmŴ; �v�nle�3i  a�[����J�]�m�H�E�h( p  � $ � �     mZγ#m�8m�:�C�m@   ۶�    �mĂI6�n��QƳ\  8       �k����si6���*�U[ T����Uv��I-� H 6�Yg$� @�g��z�    m� 	 ��-��U�&՝���`��l�	�}���ր5��9m��� ���ݰ M�f��Ԇ� mm�r�   ;m�l  � �0    �n6��m�-�@m�#�+�*����T�F�        ��B�:�j� ��m&Ä���H�$���� -� �n�v�Y%  :M,���l��� ��M���ko`  �m��h����u�ں��A��m���nlְ�  H[@ �|����UaWev�UJ���|���uK�,�\�ʵT�HrҔU[@A�b����	���A.-�$�:v  A h� m&m�&�5�lu�  p$e��B8١˵(h{�J���rQ�Ӫ��6�b��A7>�d �Jě�s�V��S�`�P5R��������^
Zr��D���e���h!�5�����Nl�]�SH�P ����1���5J��m�UJ��$MU��`�i�`�n�X�[m�NL  �`�� ۢ��ݰ�V.�s` m�0 	���f�*��z�H2�\�����Ȫ�u�%�m�� v�  8g]�ɀ6��f���8p�k�  �m��� H.�t�h ��j��*6�n�sm�  m�   ���h�J�� X"�� A��i��h	 �Ѷ�HnZ-��ȶ�h H ���[hK(  $� j� p� 6�m�� ��a�m�$ -;e�� n�ۀ �G�|   (I�� m�0   �lq��@ �[N �l�   �[\H6�\�PHm���8m���m��6�   N���[� m�� �-$��JH!Sj�,0��`  �5Wg[m���h6͛` S^�Ӥ�ۀ  �ٮ�koc�� �Zl�4�<ɶ�� �`m�������� ����]��ޠ	�mɲ�h�m�  �۩����6;v�R�OS[pG�!4�4�U�+<����� -��m:`]68 ?������w��w��w���X@@Y���A]��U����]��)�v� "$ !Nx �|�{"�4��DS��_��J���f�S ��`��]
1"<��l������PM"��P<P� z�������|��U=U������� SJpxB���( ��P(� �Á�B PUO�� �  A�B(�P�E`�X(��AyQR
��� 	� ���C��9�i��������P�51� |(� �+�=�E�� ��F��H �$H�$�#+�>N��(�OC�`H� >����E�(��	�k� �+���Ep�D>X�l�pQC�\<D]�APLO�](�<"����EAUڏ��"�	U�A<��� @       �     -�J��%.6i��݆��Z��n{�.�����I��U���x �لm�O\#"�A��[l<���k�gs�nƖ���f�	8�{m�l���)ә��M��k���2�v��(�p+��e�����/T�k�;NȮ���b�<�\�T�-�*�Z�d6�n8�\�7R�����eǱ�! �<�ꕶ�U��/lq�s�@6via�[;6��-�E7vlڛ���X���cg�;<(MEgl�UR��D�[vCqU.�UR���'�p�om�a�$ڶu��J�J�1Z��
�U�킌�nH�v] ���m�6�S��[]�U�A�q���&�;5H�"�v̀d���ӻ<�QW
 �äUI��n����nK��s;k�F���Vێ*�C��U�kHM�r;gۆ���8�R'6�;s�x7"�Ņ���ܑ��p2׈8\r ���l��n&�Y�$���N��l햮58Ʃ��}��5,�'gRq�¶��k��`�_J��ޭ�	S���S�;�e� MONZ�Ux[n'��y��b�v���n'��N�����5�-=���*��#J�:|lqqq��ٵJ���+Td!u��ki���d ��m��n��	H���nԙ٥V� KI��56lt�vQm �4���u�r�E��k7`ݭ�jCjV�7&���*ʹ�k�K-���4� o>"�G �j{r���K*�<����J�=��=��h�aU	�j�A�on���U��<�ꍷCri@0�����'5�mD�ʪdp�F��%8Xy�U�V��i��@ �<�֧ecTB ��u	�0Ầ��s�)ej�b��/.��^���E�<p2�Ay�[��(�<�̓"��9����v����-3ڨ��ѭfkF���ֲ�&���P�Q�����]��Cý���Ӊ lҳ�L#��O^\�s�,�;E�C
�]��Nɂ5����k;�`9�b.�ٴT�]�FZ�1O��p����n��\�t����gL����x����n�ɵq��sm��J�룛�4��=,��"u^�d�p��UI���Rz�S� 'Z-���GBv'���K�#�g׸Sq�U�u�c��9��7���յ�L��� b&�i��,4C0��.sɹ^|�\n0�_;v<`l{'m���nD8vy���G��ٰ3Ӆ����IBK�����k�N&�Ģ�F��/>�BP�-��6V��wM���ٰ>՚=�)�K&H�qhvt���mz�Z���h�R�<O&�U�\��& �-�V�� z�Fډ%&H�qǠyu�@�}V��gJhVנv|��&<M�1Y1�\S2OGK��p�I��\[���̭���ӥ�u0Nf5"$q5���%#�;�U�}�Қ���]k�>�⣏�:�[�Y��'����<"�@O��� +�M"���=��=�����Z{*�c�`�wwW� =rL@zܘ�o�:{�WVD�P$Ȇ5#�<�נw>�@���4+k�;�u���1(�����h���t���mz�Z�}cw)����5�E�NnIv��9�Kd��;]�@�=�[�����]�͛�H��Y2FӋ@���4+k�<�נw>�@歹�Ƅ�`��'�$��Ɉ��@s��[�����#����Ɠ�=���@�}V�Ы	
.��E	b�^z{�����u���1�cĤzx�9�� =rL@zܘ�钮<H��A���-�Δ�<��@��ٰ3'5�
.��N��Rr���Κ����m�r����V.���l�>]��k9�fI	y�8	�<����@��^�����Δ�;�WVLN%L�cR=˭zs��:S@���XA27s�zs����& =nL@zS�*��nH%�$m8��:S@�˭zN��M��TJ������h�)Z�i'�&�bp�<�����1 �9ht�:{�7oKym��	��sZ{/�9��]������eM$Mc�6t�I������������b͵�!(����wM�[��$qD�0��)�����λ����]k�>�⣏!9�o//smΜT���1�rb�r��*H2	̉�#��y[^��ֽ��Zݝw4l��ɉĤT�J%�M���ٰ:"������nI���f�y E���c	$��~{��w{�����$ m��n۾|�h�7F�IŽ3&���Y.ι�v���we:4����wN듵���	�F�N�l�c��˻W q���|���P8�Պ��>vڂ��e��<�`.q
�`�X����5vM�nk='(�+�kE�K��n�!�Q�����rȒ�j�/T����,���)n�9���z�.�mH�x9H��͌��.b�}���R�-Ԁ3�φۋ+r/\���y"r�9��8�3=�t#�3ۏQq�;5�04�ݕ������9ӊ�rL@zܘ����ڡ�:�T��\Ӱ=�6������/߿=�~zs�h�R��'��F�I����+k�;��@�λ���$r70Y 8�qǠy[^��Ih��H�& �w6�,��(��;��@�Δ�>Vנy[^�������?b��lPs���c��]v:�����f�-���>��d�-�<Y�!9�m����[�~4���Vנw>�@-�y!�%!BF)�9~���C��@�����rO}Ϋ@�Δ�-��&'�LS Ӎ�b�9h���� �:���8أ�D��������K�h埍��z���\�l �Q�IR��sN��YZX�==�?��`wϪ�9g���a0�6�c����/m���
{.��.ױ�N�'�9�ݏ7mm%$��#��N���.�����:S@=z�rF,�i9#�<����UvG7� �M�@z㘀��C1�&<JG�w�)�}�ҚO��=OEA6��־��<�}�nIϳ�Tq��72$�iHhvt���z�˭z|�� �EIq)�*�D�9�[���Ξ��~�?ֈ�۬��D��/m�d�\�ez0ps��#�J�7l�O�厌�խ�6�q�rb�� 9�� =q��;�`��NF(�8���7��f�������>{�7�D(M��x� �Q�K&H�p�-�?���.���Jh�WY�O�"5��ÒO���`y�t��,��P��=�ٙ��&OS@>�dn9#H5y�����1 ��ٰ@z㘃~~���Gd��X(
x5#�O]q�Y�y���F{�p�+����gv9�51�i�^�U�� =��6\s����⣏1��&�JC@����<�W�y}k�;���T��r��˲����1��1��|Jh�7VD8ӒH�q�_[��@sf���1�(r�.�Rn4��F��>��4��M��^�?/�����N�~O���   evy�:�0�3�3��/%����S6�����&]�$�R�
��L/?����m�\�$^$�k%���u���q�F�Y!y��;b�$[��m�m�m;��j; a4\�S���%_5���.���ɨOj��ۅ����A�+���і	���<��5��kk&u�vr[+�p[s����W�ָ�鼎����h8�YP8K7���,�����]{7���q��]��m���f㤓�6r��Lř۷�݋���լBG1,y#m��/����ֽ��^��Ϫ�;ꮸ�x'�PC����1��1��-͛���q��d�M��/�z�}V����3?�.���������H��ɛ�e�� =��9�`�����@���I��D�mG��q)�}����:��bݎZ �9���Qx��=[�z��;��d�����Q��^�v��-%��!�&������D����W�z�L@{��@sf�&C0�ٛ�j�]MUS`|��7q
��
&O�9�@������W�}��L����37�r�ٰ@z��@z�L@u�M�$sǒ6�Z�Ħ���W�y}k�=��ޤ�諭q4�O�RӚ>����m��%
�ot�ͷ�;�6�oز��������~�d�=��+��.-��m�ۭO]�>���Ųn.-۲��
�U��fA[?$���ߟ��_7սI%�gm=��t�ԒK��H�NdcĤ~�I|�V��g�m+K��y$�Y�z�Kϭ~�I*�$x#�m�oRIw}����}��7o�ʏ� wLP�!A�R$A�أ,ޗ��!�Pp`+�����0Ü�8C���Ѕ��J<B"�mY),��B#M���p��a�!�$HH`�	$� �E�$�6څ$�!!�BBB�d"B$X��$`�HIBB���ň1A�n�z�H�@�$�´��XJ���2 �%T0�RD�A�$�$(#�H`d4.�5����Y �"�c$	Q�Q޷����NÊ1_�N�*�����C{"z��8 ��F��Z�g����|�-������*�߽����Z1����?����|�m�ߧ{��=�m���ͷ�)��7�_|����wܙ��&�Y� ~?�����m�g6f�m��/�m�<�&�m�Q�����{d�Iv
�\Oc�}��th8Wiݺ����;�F���8�ںA�nX�-���%����I.㯳�I/�J=I%�ֿy$���
8��#m8ޤ��3~_}СD)�x���m���������V��6ҽ�~^�LB")3�I.V~����_��_7սI%�u�{�$}n��dly 8�m��I/>���[�g�fn�o��~�[v�M`
lP_����Z�Iz�r�s#%#��K����$����=����jI/>庒����GY���:gc[\���y^ƍ��Y��HsŐ�w������j{��VҎ'�$�}��I|�V�$��Z���S3�w��lo{��P�����[�J!�5k�m�{\M��)���t��m���3�̶����9�o�9�h���sYr8���Ԓ_;����cmsw�z�K��oy{ͷ�k��S2��#yT��njZ�a��I/�����I+K���/���g��I/�����%�l �#�X�6Ӎ�K�7i}��Ir���g�I|����m����m���K�����*����V���0�=��6���ɺ�0���N%��-��uz�՝�,�]�WdX��ڵ�x���G���b'��l����y6���2l@Wcɫg�j��\��X��틆���v9���y��OS��x�nɶ��Wl;R��q4gS���2�i�.��1�����G2,��4�\WP�=NW���QÅ�C+��Q.k�B m�Ր�j�����{��~?�qQ�,윖޸����нL�gm&��߿g���$��9v�=�נ�nG
�q]����_����$�w����K���ԗ�����y$����Y��V̂�~}�C��}��~ s��_�ͤ�/�g���;���$���"��rV\�S����S�������m�Уޖ�=�&�$�ϫ{��m�������i)���ʹ�.�=��g��I/>���%��ZԒK��RD�HB���K�ҏRIy���I/�J֤��;i�$����\X�L#]���W'۵�y�0�Y�X�Cc=�B�#��o,qs��4�#3��Y� ~?��������l�m��e���
#ޖ�=�&�m�����H0$]������'�缯T����(�տ|m��ͷ���m��wg�+��U=�:�PP��,ymƵ$��w��$�˥���y$�}+Z��J��i����(��=����jI/;k��K�ҏRI}�m=�_[�7i�$�q�K�������jI.��׼�?���������xX��c����OkKۜ���D;���ݸ����\�im����{b�LE�+.x��� �?��| ?v��$�˥���ޯ�I%_b��bnci���jI.�տy$�](�$���~�I|�V�$���)!�%$I���k3���/��f���{�s���I<|Aj ��7��컶������������FgM�����{���_��_>��I%�:��$�˥���L:�i8�q5�'��_>��I%��ݿ����g��I/�����c�&�#���KC��NnBM���+��� v�yѳsŘ�N��=V3���1�J�֤��[��K�ҏRI|�W�$�ϥkRI_�?cLM��&Ӎ��%��G�����_;���%��ZԒ]ӫ~�IZ�Ei��������ޯ�I/�J֤��[��K�ҏRI/u.H�ԃm
8�����jI.����6ߞV�m�I%q�������}<��{��U�I� ���������>�?$��ޯ�I/�J֤���?n#�}�M���v3�����l�kcĬ]�kG<��b���X�-���n`k
2��$�Y�z�K�z�y$�}+Z�K�u_������FgM��� �?�_��_>��I%�:��$�˥���]��A�e&��~ ���> �:��'����J=I%�_��]aV�
8�'�6�kRIwN���%��G�$�w���K�ҵ�$�܊���$<"2&Ӎ��%��G�$�w���K�ҵ�$��V���Uw$	$�H��I?�b�;:��{t�]&2X\lvl WC�tᐺ�����o����%��;v���.-��� �ۑ�<0��9�j\U�e!�Eu�k�y��:��ٺ��\6Sa�]�m�4s�`��y�tokjB@�vˋrK�Q���.���!�ݪ���i�\�7[�\t�/`��m;뜭�C�x�ń5cu�۱��E��/<�ؾ���w�^�3GC��2ںun��np��jO9v��=:���b之h��u�b"x|ݢ2�������~ ���-��ef��P���z�x���m����H����B�?y$�}+Z�K�uo�I/�J=I%�_��J��I�9��ƤkRIwN���%��G�$�w���K�ҵ�$���I��I(�~�I|�Q�I/���������'ս���u�8'dprC@�^���1 �ٖ��=���d����9�gJQ]2�����s���-{2�obK��Z�c�t��2�q��~���@6�e�=�`��b��^�SM�����M�������z�rI'?�����*���_u{�$^���5�`�DdM��=�Jh+��_uzwJց�ֽQE'�&�m�@��ٰ>~͛3+e�rQ	D?f����8��b�@��@����;�V�}Қ��z��Q7t\��u�u�n�q�;{�5�!<s��+JiLNg٭�ZH�,JA��ԏ�w�.Z���� =|� ��n��G�I%#Z��M���������_�@��Z�*�m'⌎Hl����f䜾{�np�
����U��t���xu��dC��&(�z���ofZ���� :`��
8�6D�q��+Z��M�z���@�g���,����nn�������Wv�.����lK��ss���q�(4�4ŉ�țn5�{��>W��<����z��<O���Ffh��bʻ=|� =�hs� u��QE�2)�q�_uzwJց�S@�^�@-�T��X'16�ԏ@��Z�=�Jh+��f�Ͽ�&�� ��)!����M$�k@�=���2b��b��- s�-5�۬��D�uv���p��øS��c6���"�f�E$և��E���f�@u�1��1 �ٗ�W�߽a�o���4��h�N=��g��$[g���Ɓ�^���ń$q,l����;�V�}Қ~���~��������EOq�,O�D�q���q�@z��A���_�H��@w~��H�X����4���/�f����v����P��$�	�DQ�W���O :#F%�i"�8�*DI�[pS[P�IX�ccjKRH��cIh�`�	F)�Ґ,(0��	 B!�h�rB�0�Ҥ�0a/�"B!�����$B(t�l,H��2Aу�G1�@�5�
A��F#X;U`�1�`��! z	U(��V@aa��@Y$���b�	9��A� ADlk!��H&*b@H4!��$b	%@0HĊ�D����1Hw��u��Ϳ�k   l      6�    �j�������9�ȣ�A�H���ʹ7��#�ف�g�zDآ��te'���.�N���[em��ڌ��$�y�Dm���ve᧰��:
�t�q��bŜ�v�9M�Mq�ֺ֑�մ�.��=�2��#�lWe�Ner�n�'�#���_,�/-mV�E6�5���8�n&,�V�+�s��̌۝��؛�ڢ7L�f����.���ɲlR���d����~ DzѴ2Ō�m��
�5U���*�H��UR�M�46�`�����SD8�lZ��-[)-W�䲭��6m��d�΅��\����4�{�z��貵9��a,��FB1��e�7��SUm=���U�k%n����k�@�{Z��Q��p�Խ��
��gs(.qu��+l��T��5ѱ\�Z�s !��<�� �ܢ&ݝ0�(�G�$藰v4���` 
V��9ϭ%g]��B����dXݠyl�'f�"p5�f�5q�Nrt�-jȊ�J]����-v�ܑ���ԫʪ�7V͙N�)�jH� fT gY0��!�vg�ںú:�Н�8䖦�Im&��3�h�M�e��Pr+��j�U�N3q�k��fn�t���˕�X;m��n�i�8٭� 	+#bN�i��6ܺ6�R��T�URr[%��nj�8��%�h�r�9$�Y��[��ɖ�P�R^+"��շ
�Q�㵳;��eUZ�3��A��UUkRxÉN֍*.����wa�>7��@U��{�m��q�U�ID �UH��˶���ظ�-!��y�+궗��gUs��ځ�j�@�J#Z���tA�P�ٲ�u�5Y�&��v�9˵U$�]�[�:lO:���N�!���v�y�m��٤r��d֛]�Q�n[�
Uh��8���ҫ[����B-�z��Y术��b���3��+ٚ�ֵ��F�G��`��t<ELBS< 	�@=����{�ӻ�����_����n����\1=�Ry#�m��ܝ8���9nۉ��u<��n�=�Z�|�����u��E�CZ��"P�dBk�(��٤�+Nv��l�n��<�l��#�s��.h͸�9H�N�z�fB�y�Rs��EGh}�B��Ծ��{&ʒ�e��v���j���t]y�S�yk8����W:�qD�\��7Si[e��DZJ!)�sr�D�H�tR��R��m�����DW�X�k��rn��^]�����S"��G�����@��Z�=�Jh+�����<1$���cR=��-~��Ü߄��؀��:\)!�����IHց�S@�^�O�ٙ�|��z�~k@������MŸni�� :㘀��m��@{����xZF�"M
'���W�s̴��q�@�ɕ�ٜ��v�7R�]s�����wa������s��S��v۞�X-�Zé��l�?6߿�fZ���� =|�#��V~�?W���G󑇛�Ы'�w���oq��{��6��ӂ���dD�����E�dMı>����ND�,K���ͧ"X�%���o�v���*dK�~�]k.�q�I��33SiȖ%�b}���6��bX�'���ͧ"X���>���]�"X���^;.�&Bd&B~���:t����K��m9ı,O3߻�ND�,K��r�9ı,O=�}�ND�,ȳ"}����ND�,K��������Ѭ�ɗZͧ"X�%���o�v��bX�'���ͧ"X�%��w��ӑ,K��=����Kı/�}�kN��g�����M=qk�w�у�#�q���ѣ�h��i-Ƶn�{Z�:g�I�9ı,O=�}�ND�,K���ͧ"X�%��{�sa�����K���K�_�	�����(�RI4M9���kZ�ND�,K���ͧ"X�%��{�siȖ%�b}���]�"X�%��m�p�!~�p���Y��S��L�r�j]\�m9ı,Os��ͧ"X�%���o�v��cP� �IO@4�X���oɴ�Kı;��w6�!2!2r��(rUM	ʚ)����%�%���o�v��bX�'���ͧ"X�%��{��ӑ,K!�ިVBA�9���5S*��J�ʙ�ĐI�{��pI�>f}�m;ı,O=���r%�bX��}�ͧ"X�{���}���4�=��Hs;����m�6�6��3�k��m�$�K�Ӧ�b������5�\sRjh˚�ND�,K���ͧ"X�%��w�ND�,Kߏ�ٴ�FBd&B�m�p�!2!2��S�WS%ѫ���Y��Kı<���iȖ%�b{���6��bX�'���ͧ"X�%��}��ӑ,KĽ���ְ��F�W2Mf���bX�'�o�iȖ%�by����r%��2&D�5��ӑ,K��߻ͧ"X�%�~�I٭
JsA2Km:��|Bd&Bd/f��,K��>�siȖ%�by���ӑ,K�u4EErĿs�iȆ��ow������sfU�[��x�,K���ͧ"X�%��{�siȖ%�b{���6��bX�'���ͧ'���{��>����`x쑢.�tE�{��x,e�8�m��"�r�wmm�6���٢ã0���������ow�����ND�,Kߏ�ٴ�Kı<���l>	�L�bX����r%�bX��V�9*��J�&f�n�&Bd&B�>�fӐ� G"dK﻿�iȖ%�b{���6��bX�'��{�ND�,K�����3Z�4e�5s�M�"X�%��o�iȖ%�by�w���Kı<�~�m9ı,O~5�nӑ,S!2gt�U6P���U2\�p�!2��>�siȖ%�by�����Kı=��ݻND�,K�~�fӑ,��L��w�T�ӢGH�Bn�n�'ı<�{��r%�bX|�~����r%�bX����6��bX�'��{�ND�,K=@�?�>���  ���:]V�[wj�����g��Y`*�Łغ�H��
�gpp�,PM$j�wJ5lN��q\�l��Jwf��;&�S����$���j]�6�Nj�<0`�vA��v���ݐ�'nv��^V��ۭt�Es��v��� ���P-�F)^�յ�<�^kP�I3���,cs�/E���[��`�n^�:�$�+��s���w �0�u�2S��em��WK��q����|:{q�8�����.��t���Sۀ.�\����,K����M�"X�%��o�iȖ%�by�w���Kı<�{ܸ_�	��	�r8���d��uSiȖ%�b{����r�Q#�2%������Kı=Ͽ~ͧ"X�#!{_�!2!t����4M;���5�M�"X�%����iȖ%�by�����K@!�2'�;�ͧ"�	��3o���	��	��h;���j��˗W3Z��r%�bX�g��m9ı,O=;�ͧ"X�%��o�iȖ%�b{���r%�bX��S��drUM�4L�T�/�L��L��]|\.D�,K�~�fӑ,K���}۴�Kı<�{��r%�bX���ɝ��A���[b{Z�u���D�웊���!�zێw[Ksဎ���ݚ^��y�N'�,K������r%�bX����v��bX�'��{�Vy"X�+)u�p�!2!2�z_�M�)�M������Kı=�_v�9  �]D�KY�{�ND�,K�N�iȖ%�b{����r'�Q\��,���~N�ӧD��T�i�/�L��N'���ٴ�Kı<���6��bX�'���ͧ"X�%��}��ӑ,K�����>����#?=ߛ�oq�X��}�ͧ"X�%��o�iȖ%�by�w���K��2'�����r%��L����~*�%9T�Im�T\/�L�ı=���m9ı,?"�u�߳i�Kı=ϻ�6��bX�'�o��|Bd&Bd,\���&��

A.��5���[F�Yfw�Щʮ�{r���8���b7�����w���oq�����ͧ"X�%��{�siȖ%�b{���6��bX�'���ͧ"X�%����~ŇFeVIg��{��7����{�si�~P9"X�t��M�"X�%������Kı<ϻ��r%�d&BΣz��SC%U)�����	�X�'�o�iȖ%�by����r%�G�E��j'����ND�,K'{��|Bd&Bd.�g9�52�St����ND�,K�~�fӑ,K��>�siȖ%�by����r%�`~AdO�w��ӑ,K������j٨a�5&�f\��r%�bX�g��m9ı,O3߻�ND�,Kߏ�ٴ�Kı<���m9ı,O~>�w5�&]=��5�1ROkKۜ�p��gr;$v�ŞgN�޺���.��N�UM+�ӫ7�Ȗ%�by����r%�bX�|}�ͧ"X�%��o�iȖ%�by�����Kı/{�{��!���\ɗZͧ"X�%������r%�bX�{��6��bX�'�߻�ND�,K���ͧ"X�%�|�I٭C&�3&[K�M�"X�%��o�iȖ%�by�����Kı<�{��r%�bX�zm�p�!2!2N.�19��r��f����K�Ȁ2'���ٴ�Kı=Ͽ~ͧ"X�%������r%�`x*����;���6��bX�B����QC��4L�M��|Bd&%��{��ӑ,K�����m9ı,O}�}�ND�,K���ͧ"X���_�J#k���D�a.hD�Ժ)�+e9�	7�퇩\�w�k�6�c�m��As<��:��&���a���gȖ%�bw��6��bX�'���ͧ"X�%��w��ӑ,K��=�siȖ%�bw>�'s4\ֳtkY�f�ӑ,K��߷ٴ�Kı<����r%�bX�g��m9ı,O�>�fӑ,K��߻3�M�HI4L�4\/�L��L�����r%�bX�g��m9ı,O�>�fӑ,K��߷ٴ�Kı/�w��"�.�ة�����{��7�����m9ı,O�>�fӑ,K��߷ٴ�Kı<����r%�bX���uMJ��S�,�57�!2!no�iȖ%�b{����r%�bX�g��m9ı,O3��6��bX�'<�w�����n$ m����[��c-_��u�9;D6(�;qBY�#-��c8ح�<�4�#��r��lV���t喺8-�7n�F[u���p��vv� 5���M�N������KG�Cp�>�A�X:�D8�vЕ�`�9{i�Q6Q�w.xy⹷�����a8 2:!���K��ؕ��gq�s�t<��X�����Y��i�ˍ/#}�}盍�o�$�Fz���8���bq@v�B���Yp��ݫ�r��tBv���Mm.�:��bX�'�~���Kı<�{��r%�bX�g��m9ı,�����_�	���O����5��jm9ı,O3��6��bX�'��{�ND�,K�O�ٴ�K�2f��!2!n�oQC��4ff�SZ�fӑ,K��=�siȖ%�b{���6��bX�'���ͧ"X���^��	��	���ޢG%UR�h��k6��bX�'��o�iȖ%�b{����r%�bX�g��m9ı,O3��6��bX�'s�d�f����E�5��3SiȖ%�b{����r%�bX�g��m9ı,O3��6��bX�'��o�iȖ%�b�;�����<�uFFB�5ջO�9�Or=���c�۷U�y��rk��sPe;9��#o�D�,K�����r%�bX�g��m9ı,O}>�fӑ,K��߷ٿw���oq����ߦ�"�.��i�r%�bX�g��m9(�*0�P��Ati�K��gw�m9ı,O~��M�"X�%��{��ӑ	��	�k:��
F�S�,�57�ı=��}�ND�,K�~�fӑ,K��;�siȖ%�by�����Kı/��;5�d��Fd�iu���Kı=���m9ı,O3��6��bX�'���ͧ"X�%�����|Bd&Bd.�]<:b��Sr��MU"X�%��{��ӑ,K��=�siȖ%�b{���6��bX�'���ͧ"X�%��}��k$�5�)�L�BٛC�L��d�^A 䇛\�����l���\m���^�ғjg��{��7�������m9ı,O}>�fӑ,K��߷ٰ�<��,K�����r%�bYQߨ��UT�*�L�T�/�L��LO}>�fӑ,K��߷ٴ�Kı<�{��r%�bX�g�w6��bX�{����n��.���w���o'���ͧ"X�%��{��ӑ,`���O��V)"Č���b�^��  DO�0��؏$H�B!HP��E�D�DXBD�
C��RZP�
I� L�����1�2,(
 �#*E�B! Q�*ED $`, �cH�qt �HB@#1"�s �U֐D��E��pE=�p���EvA`�����POT���th��
t�L�����ӑ,K�����m9ı,Osx���&Z$�
�K�.�&Bd&B�=�siȖ%�by����r%�bX��}�ͧ"X�%��o�iȖ%�c�����jb,��*~{�7���{��g�w6��bX�'ޟo�iȖ%�by����r%�bX�g��m9ı)˹;g*�4әR����(h����v�7g����x�9�Ynp\]�ۜ��a�Zͧ"X�%�����r%�bX�{��6��bX�'�߻�ND�,K����ӑ,Kľw��֡���2��SiȖ%�by����r%�bX�g~�m9ı,O3߻�ND�L��[�o���	��	��ut��U�un�kFkZ�ND�,K���ͧ"X�%��{�siȖ%�b}���6���L��^;.�&Bd&Bݠޢ��W,�˫���fӑ,K��=����Kı>��}�ND�,K�~�fӑ,K�O �����3iȖ%�b}�o��Z���r���~oq������n��9ı,O=�}�ND�,K��{�ND�,K����ӑ,Kǿ�~�?[[��ezu�/\�{m���z�s���6�m�4&2�d<y.5��-��]Fff�ӑ,K��߷ٴ�Kı<�����Kı<�~�m9ı,On��_�	��3x���ܵ2���f\��r%�bX�g{��r%�bX�g�w6��bX�'�}���r%�bR�o���	��	���zYU4��#�5�]kY��Kı<�~�m9ı,O>�y۴�Kı<���m9ıL����_�	��	�j}N�	��0�.��ND�,�02'{�g��Kı=���6��bX�'�߻�ND�,K����ӑ,Kľ���֡���a.�WiȖ%�by����r%�bX~�����O"X�%��}�ٴ�Kı=���nӑ,K��߾���H �`4��t�V�ٴ��k��������ǎ�#�[�B���7Gm��2��[N�m�[����eG��F2�����]��NR����V).�t�95���[�f!,@�%ͮ�Qp�h�`��ϾcuŃt���X1H[��ZB�x�K���\c�M��+ɪ�,/v��r0mƢ����n��a��K����V�Ǝz��[[���Y�/�����q�|~Z �cnvm�]I�V�;n���Ì�k`�m�p�&8��I5��� ��mjz�D�,K��߳iȖ%�by����r%�bX�}��iȖ%�by���!2!f�7��f�*j[��Y�ͧ"X�%��{�siȖ%�b}����ӑ,K��߷ٴ�Kı=9�7�!2!gQ����UU&J�335�ND�,K��w6��bX�'���ͧ"X�%��{��ӑ,K�^�ޛ��	��	��s��өT�-j���m9ı,O=�}�ND�,K���ͧ"X�%��{�siȖ%�H[���p�!2!2f�?QM�i�5&jܹ���Kı<�{��r%�bX�g�w6��bX�'����iȖ%�by����r%�bX�{�s�&FRiؑl\۳.��'ss��eE�A���[g'&�2���%I�����v
~{�7��bX�g�w6��bX�'����iȖ%�by�����%�bX�g{��r%�bX�������n�Yp�u��r%�bX�k�ݧ!@� T�A_���n%�bw�7ɴ�Kı=�߿fӑ,K��=����Kı.�#��4ܪU(������L��^��fӑ,K��;��ӑ,K��=����Kı>>���r%�bX�ϻ���R	�����{��6������
�/<ޛP�BX�6�X�.!{6��_�	�����B��.�k%�jk3Y��Kı<�{��r%�bX�}�m9ı,O}�}�ND�,K��{�ND�,K�}�wjڻ��-Ư���8|T�ލ��<4]k��짜OOT�����h��D��i��=߳ŉbX�;���r%�bX����6��bX�'���6��bX�'��{�NG��7�����}kOAu�����X�%��o�iȖ%�by��siȖ%�by�����Kı>>���r)��	�����E6�2�M˚.�X�%��w�ͧ"X�%��{��ӑ,bh�B(B<��!��7�_o�iȖ%�b}�wٴ�K�L����ʩ�N�"��M����N%��{��ӑ,K�����m9ı,O}�}�ND�,K��{�ND�,K�����-ѫ..k6��bX�'��o�iȖ%�b{����r%�bX�g{��r%�bX�g��m9�q������1��N�z�H�]:��ۑ�vLvr=G���N��u�t랐��ц�a��SiȖ%�b{����r%�bX�g{��r%�bX�g��m9ı,O~>�fӑ,K��zw;.��k2��֌ֵ6��bX�'��{�ND�,K���ͧ"X�%������r%�bX����6��bX�'�h�wPV��m,��~oq�����~�~{�ı,O~>�fӑ,K��߷ٴ�Kı<ϻ��r%�bX��S�҉�s�����������۹����~�ND�,K﻿�iȖ%�by�����K���������7����{��7�����Z��]K�m�"X�%��o�iȖ%�by�����Kı<�{��r%�bX�z}���!2!f��**�r厔��������X[�uWm���+#��ꍞ�>ݹv�KV��5��6����{��7����w��ӑ,K��=�siȖ%�b}���6��bX�'���ͧ"X�%����=4��#�U@�n�&Bd&B�=�siȖ%�b}���6��bX�'���ͧ"X�%��w��ӑ,K�>�O���Ҧ9D���_�	���z}�ͧ"X�%��o�iȖ%�by�����Kı<�{��r%�bX������54a�Xe!u���Kı=���m9ı,O3��6��bX�'��{�ND�,K�O�ٴ�KǍ������#4�U�[��{��2X�g��m9ı,O3��6��bX�'��o�iȖ%�b{����r%�HL��P�BD(_����UUUUUUUUS��uvuC��f#��4�c'�{1��6L�Xv3@狭����W��C5F��ⱉ��vK7i.�k��\�SqW�$��kWa�"�{7c�N�z�nӏ]���6�J�ǡp��Lo��:�<ev�� +�&���A�T���lu����%�y	c;�j^6������,��t������rn��:�`��s���ww�w{�+���풳���М��3�պ���M�6�aa�}�n�l[:.�e`�cM��������ŉ�?���ӑ,K�����m9ı,O}�}�ND�,K����ӑ,K=��~�������7=\�?=ߛ�oq�����m9���,O~��M�"X�%��}�ٴ�Kı<�~�m9����ow���}kOAu/-�{�ı,O=�}�ND�,K����ӑ,K��=����Kı<��}�{�{��7��������(�����Kű<�~�m9ı,O3߻�ND�,K�O�ٴ�K�,O=�}.�&Bd&B~�l��t��*�s5�ND�,K����ӑ,K�����m9ı,O=�}�ND�,K����ӑ,K��*�{�~ֵ��Jf�Lqڲ�']]/gv<1�����%v�=eP໷3���7��t��S�����%�b{����ND�,K�~�fӑ,K��=���D�,K����Ӓ!2!<�GD�9��RНQp��bX�'���ͧ!����Ȯ�D�K���ͧ"X�%��}�ٴ�Kı<��}�NAKı;��*[�u%7Jj���p�!2!2�7�iȖ%�by����r%�bX�z}�ͧ"X�%��o�iȖ%�bw��o����lT��~oq���{���߻�ND�,K�O�ٴ�Kı<���m9ıV��=����Kĳ������TOU��U�����7���'��o�iȖ%�a�c�����%�bX�����ND�,K����ӑ�7������᭺���tA�{Y,��4j�9ǞM�C$�[)�ݩ��F�I������;�Xbz�ym�������ow���}�ND�,K����ӑ,K��=����Kı<��}�ND�,K�����
<����w���oq������ӑı/���m9ı,O=>�fӑ,K��߷ٴ��L��O�͓�N��H�C���_�K��=����Kı<��}�ND��E{@�F�a������M�"X�%��{�siȖ%�b^��;u��Yn�[pֶ̺��bX6'��o�iȖ%�by����r%�bX�g�w6��bX��=�����Kı/ߺO�Z��E�)�M�"X�%��o�iȖ%�` y�w���Kı/���m9ı,O~>�fӑ,K������
hѩ4L�n\4�ڋ�]���n�@�90Gȳ;�3�nq�c������|�~i'A1v�|�~oq�����~����Kı/����r%�bX�|}�ͧ"X�%��o�iȖ%�bw�~m���]4�������7���{�=�u��?(Q��,N���M�"X�%������Kı<�����S!2!n��US�UULR�������%�b}���6��bX�'���ͧ"X��%��w�ͧ"X�%�|����w���oq��_��}kOAu/-6��bX %��o�iȖ%�by��siȖ%�b_=�u��K�ڠ�|M��G�:o�M�"X�{��������@"�a|�~oq��K��{�ND�,KP�{��iȖ%�b}���6��bX�'���ͧ#���ow��|~�hx��0G71F�����+�;7ܼ�&,�f�h�k��J=n�3SN��H�C���_�	��	�;�ӑ,K�����m9ı,O}�}�^D�,K���ͧ"X�%�{��uR�Cr����_�	��>>�fӐ�@W"dK﻿�iȖ%�b{���6��bX�%���[ND�8RBd'߿#�TH��*X��_�K������r%�bX�g��m9�T�,K��bX�'�O�ٷ�7���{�������u0e����r%�g�T��=�~ͧ"X�%�}���m9ı,O��o�iȖ%����������L��]��ʙ��VkYsR�5�ND�,K��{��"X�%�����m9ı,O}�}�ND�,K���ͧ"X�%����!0w."�a��B$�dQ6>��%�T������	Be-(���4j|�� ����̀�M���� >8� :
VE��@�`�!��Ѡ`�H!9�h)v�J
F�P�,�ԈB���Q�
�[�6�ʨP �@��F,T�P�9pp�`��0	@��GP��
FB�PjeFx���1O*sA"hI!6)�1��F�-'�����������`  p �`      ���    �PL�,ڤm�Y�S[նk�����΍ۉz]��pp��Cd��M؍���-+Vn��;��%��B�]�i�]�D`�x�����kfհk�m�1Y�ۂ�ƹ�9d�a�]��`�ݞ��c�{1�� &�vL�RI]�i��Ό�����mc���Ů�m'N�g4P�kh�r� +�T�u..I{l� <m,q��}^�����
J��V�XS8ۆԲ�Bfa$WcRsm�vx��s�"À5��p��+�j�R@v�
���,t���UUn�g���e�!VکS"ղ��Y�leY82�����о{P��Ws�J��&����I�ES�P�6�eX��F0sr�5ۣ�����V��7f��m[g�δ�I:㪥���)$�6�1��M��sʝv�Knmn�{m��ۖiv$�7H򽕉��`��t3;N�X�5�O=l�u��b	W�c�,�]����f퇊��3/3h�YJN��R�,���IUn��Y�=y�]V�Q*�l��� ,�Pl$I�=��qj�Ŷ�\����h�enR0�@S�@*е(��JL�D<�������i�A���۱�2��:8}�B1E�Vy��,	d�A�<�J��:�S5�6*�-�r'm���8 �;m�;W8]��%m��mۄK*�UA,[��Z�L�8��D�UU0v�;`�l�o l��\��ARی��'���[��AEm*ʹF��od�9�5UUɴ��d�c�elax��e���
����"�����j��Α�Ԭ�2 �7l�j��Qڝ�A�����{8rId��ڻ89Q���j�bR�H�Rzઈɑ�2m���`SOa��H@m��]v����ڰ����@V� [Y�k������Yې�Z'�8��#�����nʲ:mt*�Z�lh�q[�;irk5��u�K��숌�@<Aj������6
h��ww����ֿ� m��ĂF�+"�,v�{3�F�h�rn�������]g�,�g��n�x7f܋9壃0\1!F���EŶ��dmm=]��j�9�R��]��d�P�p:9ݎr8�V�Ŏ+��y�=�����s�[v�l�$���-gnN^��ń���[S�[k�x����:H�)⵶힥χ���gJLk<
tl�h�۳t�$��Zɭ��n�f!�ӝ��	=�����y������t��t2�t3�������m�T��&�\�k[O�X�%��g���r%�bX����6��bX�'��{�D�,K���ͧ"X�%����;�5sW0�n�j����r%�bX����6��bX�'��{�ND�,K��{��"X�%�����m9[ı<���榭��2�f��356��bX�'���6��bX�%���[ND�,Kߧ���r%�bX����6��bX�%���2�ST��Mh�u��r%�b�b_=�u��Kı>�}�ͧ"X�%��o�iȖ%�'���6��bX�%��s���*���U����L��^�>�fӑ,K��߷ٴ�Kı<�����Kı/���m9ı,W�K��L���hT��$r���72��݋s�X:<�+�9�ݯK7��D�c�~w�}�>��M�,T\/�	��7��p�ı,O3��m9ı,K�w[ND�,Kߧ���r%�bX�ώ�f��)��*����|Bd&Bd/OwM��>����& ���ND�.��u��Kı=�}�ͧ"X�%��o�iȟ�S*dK�tOߵffj�ֵ����Y��Kı/�w����bX�'�O�ٴ�K�,O=�}�ND�,S!z{�n�&Bd&B����䪪a��\�ֶ��bY�H�����r%�bX�����ND�,K��{�ND�,[����ӑ,K��{�N�\��4[�Z�356��bX�'���ͧ"X�%��w�ͧ"X�%�|���iȖ%�b{��}�ND�,K�=�;������ Ě���y1�D{m��v�.-a��t$���]և5W(N�+o��Ȗ%�by��siȖ%�e�߻�I=����ސ���Xo期����U#77��@s��{�I���IJD<MI4��M�t�n"�0A +�39~��ܒ{��kr�Q�T�EM�,TX~���o����b �9�c� :�˶E ���r�����4��M�t��˫�q�MI�?�8�Y$:��L����s�vG�ú�Ty�h�z��f���#��%#�}�hqҚ��M�����y$�ǒbmȀ�=���\���_W�ߪ�#����dN&�bS$Ln�g�@�����6{7���6��=��n��e��X�n�����4��M������b)�=ǟg~�7$�w�bg�E��&8��u��t���S@��n(��%XW%�����:�����S<=�u�]�XG�XnB��~����0���x��x����{���b �9����t��,4�����M�}�6�ޫ�:�h;+�i8��&7��h�& s���UU]�O� 9��@G�[ӂ�#��%#�}�h��r���ZXr����`n�USrUU1en��f��qR��\�����1~O�C�E	['��֤����:$�-Z�[�4�"�i	�I��ɺ�)�4��睱�lꐋD݆ݮ+���Bc��3�v���w#xG�x�۝N뢹��.s>��i�X�]�m]7\\������ܜ'TRGX��k��FѮgg�yH��ca�49Q����3�Sh ꍑ7a��6�7h9{�����Y�G��d�
��:�mÄ5klm�cq�RLі�5�ɐ�5�z���{<�ͮ�㋵a:�X:�Η�����8��;F�s&��l�t�v󵸝L�t0�p]K�T���q`|�vl�f��BP��;���s@�����#ciG4ۆ��mv�ٳ`f,�V����BJg4��)�(tH����7���Y���B_s������9��<m5�W���ۧ=H�o��$������I���o���{��?gϻ��<�zlśj�=�;E*�9�Cۭ���[�.�;n��\rc����Y�Wcl�7!g A�y#i�H�6�9���/f́��mw�=�\X���r���S���n�l��f�(���6Ձ�ei�y[^�ċL?H�qI�$�ۏ@��ʐ�@z䘀�󘀍��܂qG��#x���t���ֽ��@������G�$6�Ҏ,i���rb��>� �O� =�`���������;N	V�۲��j`�gv�ex�^�nzعޫvn����m��U8uh�ض����@z��@s� =�`���1 n�kj�!���*e�M��Y���(I�ٵŁ��`|��7Д(��C�r?5���5�'3@���˭zO��Z��(�%����lbݵ`b��N%"Y1�NC@��^���W�}�6Շ興OٷŁ�(�-�U:����w�st�����hgs�!m!��H"D�������۬qⱏg�����Nq.�,��G`�%ڤk�
�ݬ���ҧʐ�@zۙ�z×_�@���_�N(�bSo��{�X<͛��ٰ>śj��!B��&�~Ȑ�J8���4_������@� ;�� {���44�.�7h�56�۳`}�6Ձ�ei`�Q	/B�I}
�y{6���!1�����U�:qR����s���1 {��cv<����,닮��vN;#�{M���i��<tc��ʖ1��Z����L��ͤs� =m�@z�L���:T�R �\���m8��dc!�yu�@����śj�����СD$�1�{�-�QUM�MM���`{m�:!%wY��>W��^�#NL�#&I���A�V�O�H�� =nL@z�L@[�]�qG���x���S@�����<�سmX����}TT����IR2D�kn��^�6нƹ�j}w7n@.iy��[uN�����:�^�܃�4IA�n�k�6��`�U$f3ʓ�몓�gu�eܑ-�wmS��V�e�]9�8�/@�kRg�mɲX-��m�AA�۩xE��f�.MJ�r˴�냳�m����1��qȝ�Vr�0=&�px�-e�ۀ�v���m��|���VL�/��ލv�Z�����ۍ���������ݷg��57 �9"Clm(���p�_���<���śk���f�����SN�������vo�%ٸoZ�36��>}k��AT�0�%?�iH�K�i��[���u!������	��>�Z�.��~�i{4�s��Ѵ�R%��i��=nL@zܘ�lqR����r���N�6�m�vn�N��Ok��뵅:��n�vrr�(@��zh�o�������X�y�����M��fڰ=���(Q0����߿L?Hӓ$�ɒcmǠww6�|�� � ��{͛�y~�srN.���#����qG)�&93@�zՁ��ٳ�%����7M�V��=�bm�X�rf��ֽ˭za���BP�����3�9:����"]T�<ݛ�(�[����j���^�oK$�a��8ܑ"'^����7�0/9��X{Ik�v�!�|�\�����v��@�b��cM)����}�)�yu�@��^�we���NhlTX̭/򈈅�!DDɏ�~�~�6qҚN����"�X�Ɯ��߾��9}����|�j��1!�*�P�L3�ȑ��E� i�$HC-��A��`�H�e�@�	BCS��VS2\ �n:P�P�
�X��DV�B*P#Q �V'��,��,"��`%R�f
'���P 1!�l�@�t ���P=D7T����(��⾚��޾��y��l�4f����r4ɔ�jl9(�	�w�=��Ɓ�t���mz�adjJUR�
�33S`{�,Q�f���/߿=˭z���	��bqb]I��Ok�.�cF�	��͜��wk�>���n�I
G�61D��qG)�&'��Ɓ廳`|�v(�I|�4�����&�r�ڍǍ��y[^��ֽ�:R��ei}	$�a�Ó�*�A�&�sq�>�ǰ@s{�I�ی'hBct�'2۪��P��|\�߾�f䜿}�n@v`@V?�"�Q
bEHmF
���}�~z�촑�ȜО��>o`���1�rb���UU~�_z7ݷ?xv���Dl����^��� ݥ��98l���s���ӿ���|5��H0B,�cR����=˭z�t���t���íMĘG�%#�<���BP�l�6��3v��>{�6��,�G	&bmǠ}�JhwJiТ!7���`��71�ҩ��R�7Ji���7o�ϻ��>�ڰ�����Ի��;���H�Ǎ��p�=rL@rj��o`���U�~�G���  2�uΖ���T�z�c�s!��Xti5<�ӻYA��9�nWVn�E�&�켍�up;a[H���mJd���w<\�Ēbq:��Ý����LU%Λ����g�����ٵ֮�}q�:�#L�v���ِ ݛuP;�e�r�+�)[���]��ʌ�6�㸬�np���	ng�V������P&�L�I<�QJ*��nj��<[Y0Csf�������/nv�ɉ�mks ����z����|��?;R�7���`����<ǰ@s{�9���j�bSƚ�@�)�}�4�>{�6�f����D~��!��~*<_�8�<!�w���hW��wY�{���*�+�i3"�X�Ƥ,:��=�6��M��ZXfV���M7aCx��@��@��{M�>۵Ł��ٰ1���U-�{Y��=��zt��ݰ�/��ȸ�p�6��	�t��)����{T���WOͷ��{�� =q�@zۘ�����sN���SNG4XfV�I%�����C�>�$�Pc� =��v��j76����z�˺�?g���%�,�h[?��Lw	Ĝb�9#�=m�@y�`��{~�_����� �q3�0�%1Lm�8�qҚ�#۷��y���<͛�x�N�)�����Ð����۠���Ր�g�>�%�	v�oO6��Cl�&�ͷ�������́����
">a����9���L�E41���z�uz}�ZXfV���1�{�.f�����U�n :����Q��\sم���H�0�r=ٟدd����w��<�W�ywW�_�)IqG0Q7�Š{�U�y^�@��@�)�v�B���=4�2���n\��3պ��\lBm�ev���Ŕ��a�nMw_��l[	x�Pm'�r�~�=˺����h��h�Q1܊q�`�@��g�E�w��>��Z�����j�bSƞ$��;�}V��}V���~������vZH�D�6�h���=Ϫ�<�W�ywW�˿��F��(�*���;-��W��&a"��1�������ՎZ���2i��Wny�/=[��藶��7\�]����4�Ŵ����8�0�ڠ^~m������)�v�9���<�zl�uT��$H�I����c�s�+��]��$^�Lm&7���$��ܴ���
�� 'V9h7-n�U�CiFF��Z���.��p����� ��&;�&4�50RG�zۘ��1�@y㖀��1 ��W�*�ޛ����� l��V�*�V�K�;��a������fu��N���m������2@C'W\�Sն+@�.���=vy�-����a��a��)���+qa:�N*��kpz����6������ ������I�g,{�x���GV���C[j��O:|Xj�����GV���8���r������N6��l�f��V�����\���ߖy�)ڹ-�k��'u��k���ԕ�������XnLN��1��y5��bN:~��@�>�@�^���^�{��G��8D�I�#�@�>�@�^���^��U�U�WH�f(��qhW��<�����}G-���|�n6�I�4����v�z�w��=Ϫ�<�W�[fF��"DȦ��p���Қ���.��Y�:�0O�"ddM��AzwK�og��{b�7�6�i�<�˺.�z�V���Ϛ��9�&8��^�����z�Z�p����5�6�di�L�=q�]UWg[�f9hn*@&;�A�RL��]k�=�����޵`y��������N��IH�?��K�ho����z�Z�ݖ�<_��&�OZ�n��z��ֽ�>�@>��$i$��s�{]�����odܠ�>�v��i���q@nB�!1<n��F�Ɔ6�hW��>]k�=������u��q��n��Yy���rb��-�EH\��zadiBH�L�n=�>�rO=�훚C�6+!�P*�aF$) �����-L%HD$�$��(K��_�M������n��'sɎ&'�.��{4����.��qҚ�����ڌq�UR�>{�6~Q]ߧ�g_��ݼ�=��X<&5�`�M�C	��Cl�v��v�m؜o>�wl�oN��A�L�nE�� :ۘ����"��Uz�Ϸ��=�ܾ�,��9����a������ :ܘ���:W��W4S�۔�TX�֬��͟�I�W��}G-���_�j&$���繳`y���a9��Д(��!%�
���߾7$�~.\�fau��Yy���b��- �� =qǠ/:�D�k�dQH"D?�3rO;u��jx�֎�d�]Nt�m���j�z���44��Q��@�s@��������c��;9�⩹�SI�JjeLӰ�-��1�bs6��_��/屨xڌq�'��w��@��Ħ���� ��4�5�L��uU6�J~�ޛ�N�3Ӛ�?$�����g7/�D���̺����- ���9�\�
����V�z�@��S\��q*֕�A� P���C�A� A�bB�@����eR:T�TX Sf9��a�QH�yP�$h�H4,$ZD�BI���t�T�PI���zDw�F��j��mF�	�Y��;�wOt��_���� @       Ͷ     ^�.K����ݴ:��S���*��&֪���5� On2E؟U�29+gsh�<�F�Sۋ�t����Q�����Vl읪{dyh�S��c�F[��h���61
'6�*�.��D"�U��F���ض�6���c�ʗmh֍=�J� 66ST�0cE��qԀ9��Q�[��ϔSt(r�ɂ�3C��:
*	(��vʤ�l��2u����<D*Ӛ��x�9��A�!�nS�v��-�����NlD�PJ�UWe��un��ڛM�Wv
v�kj�A:H�Ή5� Auf�[�Ͷ�YRsZ����*��*���×��bB���z9�vmM����U�5�YI[�˞�e�n��-�a� ��&�=����Y�s�<����q1D�l������>�D�oX�5�R"��ji�,�;vne�p������1O%*�إ�w+�]�k6�B�3��ڕʛ
[�kҎXr�o �#�N6�uڀ�Kn�'vB�ram�A�m��^M��z�ej-�sYf�U�ӡ@Z����ɩ���筹���q�t�;�D][/+����"s[n�i	
^�UZL��P�8^6P�U�zo�d��v2{t��u8 ��ն�xݝ�t���H�N4�+I����m��H�hpӪN�FU�����p[g�9Cg@�ʭP ���S���ȭK�;���h��Z�m�u�OZ�I�F`���3�f�g�)�O;!�P��ѩB^V�$:j���p���K�X6���'9�V�n�S��*�U�=Yk�cP�y�D�s�X�$�Z�pj�nts�z1UQv8��a��v��Y���j����mtpmhܮ�5�[V��\am��iv�H�.�$t�˞�wv���Cs�1�3ȼ�͠%�m؝-N���)��-k�� ��+amˆ����m��3��E1>@��G�ͨ	�b�٠�AQ�1U4�"��� �s���"�E�߷��MjMkZֵ�b�T�خ�ɞ	;�:��\c�m��!u�c�w<��:�4I׷6uX�I�)*s��lc����fP�7;��O[�M�n�N�*lt�):�v��)�n=lR�,��胭%T���rU��5�����5nV���r�A�Uc�H9)�Fd��&k�m���;\�1s�t�ͤ�ۺ��+�W���cm�l��3�wT�2���͵�:�뫥�vG��n9��:���і��øol�jx��F$؈��|�Z���+k�$�B^��'�;�����ԐT�r7$�m�=q�@u�1�c����-}UUh��D��RA7�8�V�z�:���Z���zadj<�$Lq���{��@��ՠy^�C�b����?uJ~$I�Ĳc�c�@�ϥ�=q�@z��@c��nnJ�t�:�9,��h��U�n	����VD4��F��ɘ�<����$�s�Nt���O� {���9�v9h�]˝R�Y.�IHuU6��j�� #�H�X$
�����$
B
� H�V
p�߿n��M@s�-�b �ysJ�&��4�u��v���z��f�{��G��8�NE�MݒZ�������u>��ះ�F��LrE�y^�@>����:��;V�\���P� �n�e��c��׉S���y�c�iP�"��|k�Lλ}���7j)�ō8�.���w��h�ڴ+������y$X�$�7w�sP�r��� =|�/�#�T��D�RA,���94���Br��ٸ�PdE��! �U+����ƾ]|��[4}�lq��Jc#m8�+������:���f$�Nu���w�r��R�t�*C���nj }Nj�$��9�	&�ݣp�l�٣5T���{;��q/��͞:�����6�����������nu�p5��}�<����UU~���>���߉,�� &�x��=�ՠynl�y�6�Y����q<MIMK�\�UN����<�6l���z�k��h q���q�N=��]�g�mXd�舄�~S���`wl��I2F
d���}�f�����uz�X��&'RA�Ok�Mn6ƍv�=��Y�!W_�����IF^�a6�b�se�6�����m�z���_�3��M�-�<Cj1�ڎ����g�G+= ����>ͭ/�DD�g�r�Q52�:e"j�l}ߦ�3�6��	7�������^@�0F$L�6�q�~�įe�4oW�sfÿ(Jv��M�g/ߊ�N)��ԏ���hW��>]��yfՁ�j"��K��PUUUUP �5��2�I�bݳ�w5��'�*H���s9q�:�7/]d�f޹g��(䍧db;N�*'����8�뗬he�l�ͱoT݁w����^��f��^K���Mϲ��'����,�ێz��"S�g8�����a�`9tˈv�c��Z�%z_*��9ʖy�u��q_��<���5O�U-���3��;;uFW��r�0T����:5�u�ۯV�lge��kWv�g�n��-;�8-�ѝ����^ai:�`�?��I��H�����|����ͯ�B���{�����&jfS��̬��@u�S���d����1oL,�G	)�LrG��u��{�΅
���1����n��n��`��87�M��Z�����^������e�4��[x��m(��Z�9��~���>� GS�@y㖍�߽�?�3������u�G�8Qóx��ۯ*3fѶS�#ն�d�u"VI2\W������S���c��U_�a���`��z�16TR��3S`�R��Y\io'րv�؀��1 yԄ�A�$��#�&��}V��z�?ؒ���zlqoU���%k� ��������1��1 >�5��-��7a$xӏ@����?B���ޯ��N�>{�6<ٝT�5W�>��1c�e��<H�8v]�Gj8*	a�[ۛ�"��j;5�ð�I'��NjݎZ�����n͆��S�D�)���U���5��	&�>ޛ�������=�U��4�m�8�357$��߳rN_=�76i��D=8<??�4ߧ�@=Ne�Q����&���b |�=��=q�@�ĉ�1���@;�@�Ϫ�<�W�y}�����\PpBn,bfᘡr�u���g��󝫐Z	3���	s�k����	,��I�jF��=��+��_uz�u�_g<�#9�0B��@z㘽Wa�f�>�P�f�UT���n$�)4��?.���w���>�@�^�@��,�I1ƅJ����á$����;����ٰ�P��5����3rO��JH��L@pnI�{��h+��?f̀g�j���FJݞ�
a2Θ³�d�V�v���06��]�c:#ۧ���2F��RI����\����>�}~`��I�s� ��i��V^՛�f����b }&�=��:�W�^CV3Fd��n= רּs� :㘀��<�Cw*�L�Q���@��)�|�W�y}��}l�*�9�QD�E1	Hh+��s�5�{_�~�Uķ4���nl�uY�)�i9ٻ���x���ܝ��ەt�6e)̥&i���
y\�q���H�����M�Nm��N�9������~|�'�a�ó����V�A��zG��꺰6�V��d�WeDN���6��;jۉ�Ͳ��i�]t�˰#��l8�$8n��NxY�F�%6�]��n+;>�X;=�J\�/M�{ki��)v���w~����g`F۞s��]Ek��{m�Aul����6^�7%�����Y9zלl1��;U��g���O� >�P� :㘀�mcNLr!L�c�= ﭚ�빠|�W�ywW�_�)IqI���n*@u�1�nb }&������q����|�W�y}��}l�=�]� ��ꉨ<jb$ɸ���I�s��q�@z�q�Ϛڸ$⍣PqG]q�uθ���.�C�3m�p�bnA2V��:w\)���I�s��q�@z��@�U#�q�1�#�h��������� J��D A$�4	d�sf���ٰ��_�l�es�"��m�Yw�HO���1 >�P�wTA��	2&�����V�I�s��q�@7�Hn^n�a�n��{������8�����^��s��$i���%^���M�ͼgI�����q��5�n�{p�lAZ���t�4�����H�� =|� ��@������q��M�L�>W�@z��@����H����^�R�2�	���>y�6�ݫ%LB��D��@�F���m��D..�&B}�P��n��W�YHT�aF��.L��15�aBT!E�ig#m$7��j$�� <��HiqHs��)�uU`�Sx��]@$F"� D1	�� �<Mz| hPp�B��}���=�}^�}yX`�Y�i8���hn*@u�1�nb�m��ʽ+7ڑ�4w]��z�˺� �nՁ�B~ޞ��@ɩC�T��UKں�c�`�r��Q�n3.W�[u�I��OZ.^�D�E1	9�����]��}mtDB_0��Z�<�w�D�7!T��Sy����1 >�Pn*@u�1 ���4��ȉ�LnG���@�u��>W��<���/ܔ��8��C	����	?n������`|�6l>R��1�-�uR��'��&�ؤ��9��$�<�j��H�1`�l���+Ԗ�Z�ࡶ�[��ݞr��	��;&���w�G���<�����nb �&�<�T�����/h�D�&�2����v��6{w�X������^��b�Ǌ�#i�&n���H��@zۘ�'I�	Q��a�H�$�h�U�ywW��f��빠yuD��$Țʹ���t���qR<r��
��(�I�|kRkZֵ�j۠v�S�C;Es�gI��N�֍٥t�Z�nz谊K;q!ץ4�k�h	ݵ����`�&wNM2�]�)�w#�!�MW����D�8�q���kr]ʱ��U��k�&K@�	ۛ�K6i�lm�<v�6ލv��z��i����|nʌ��(�PU��V���\��r�si�C�l�cd��=�˶8�GI�^�Ã���6�ۦ���vj̅���D4�E ֍�S�W1�UrӮ�w����ۢI-�5I쫨;t��4��Bwmnqtuٴ�eѮ��������@y��9h��@>w{ۼۓ	�h��h�����@�W��УJL�/7- y��t���qR ��n�fh񩈐"�- �u�~�h��hאՇ��S��ӓ@/�j��H	��=m�@��ݬ�ܵ����sH]]/g8z�<��ކN��8�"��n���,�ngJ)M_6ߟ��ʐ㖀��1 NsP��(�4��1��`o�5�(���J6
�j�u�@��s@�uD�0�"�4��� �f՟�$��޵`v;�h��n@S#x7�_��n*@N�-;$���̽/6�a!��rM�]����h�٠{�8��8��53"��ئ�7�V<�edC[V4l	n��bfg���ľ2�<$q�F�&x���@�;V�_���(I|÷zՀgkꪙ�R�i2�)�S�7Ӻ�ICa��Vn��rs]�P�gk%�H�))9���`��nI����s�QO�T���s���?ߖ���Ǌ�#i�#�h��9h	�%�	�j܆Cw
�
�1��`nNk�?B]��� ��s6Ձ�BP���Z��i�R��]��q�=��sս���oi2g''(�v�Wi�$��q&dMqx��~Z~�h��h�U�w<:�i�9S)�&i��v����֬��v�ڴ��+PnE1L��q��/u�@G�Z���� Kٗ�e�SNX�[�V�����;~�6�vՀ���
!$�j�=��j��tMPʠ�UN������BIvw|�6���/>�@�W$x&��O))�/WK��p�M�2�ˎ!��ts�1$T����w�wL&聉�M"e�����V�6�@���˭z���,���I����@sqR<r��& 'H�WȒ�"�$Bs4Ϫ�<����(���������{�Z�>a�����	2&���.���w4���y�ZsîF���2a"mǠo�mX�����v��>y�6��{�������d��Me�K�+�[t��o)�j�z�i�Z����mJ*%��E��H�kK����N4Ʋ��%f��mհ�bxM���l��XK��C.�\m[L�ײ��ltq1q\A���t��ܼ�$���i��`��U�v�C���۩x�?��,��h8�ڗ���.�6�◫�3�9R�:ްvbbz��89�"�q�v㍞�V�xE>F�
��Sw7����%ִk,m�՞���	7�ۛ�3�ݯMg4��w������D���D����LS 8�s?��nh�U�yu�@�[��w�J�hO	L�ԷT���w�J!$���`vwZ�>��\�<Pnb$��@��1:EHn*@G�Z ��2i�#�sґ��w4���y�V�'���=�wR��iMKs.\�����㖀��1:EH���Ɉ��7��	1e۴���%��N.���D���k�mz)!e�y�����Ɉ	�*���~�X9nh �� �I��&Šyu�:�UR���� ='ʐ㖀o(r����DL#M�������sO�ff%���h+���;�S��㚚V�BI��|���v�7f��n�h�R��GB�)3@������� 9���Orf���awhLt�l�O{s�8^/m�.웯*3f׀0�v���W��=��{��/��uK�b��!�>��T��⮯XKr�������6��@�d�}ۚW��<ݛ�
"g�N�jSTMUH�\��Vn��rs]�$��IBRy����w4
�+�ma�	�I��/Nk�>y�6�vՇBP�y��+��C�<�d�8�.���w4���y�Z.�ܑ���p%�V�������@>G��\u��e���*���������Q�i��~�s@���h�U�yu�@��&�c��Ұ=����P�;gy�{�6�ws@歹�О8�iI���h�& 'H���H����yW��"�2�U;Q
?N�M���j��fڰ��B���(Iz��y��XOQ*��ڼ˽�@N�R���㖀��^�r�\��$�qdi���
���4��l9Cj��&v�C,��7!�3�A�q��i����s@���˭�(P�a��j�竧��h�TRcy�����Ɉ	�*@sqR��n$�"&Šyu�@�[��%
7��j���`fJ3h�f��/p7/37�T���x�=nנw�GS��I����q��>��绳`o�mX,��P������1C�x��(������
Cϑ�L��f h�O���S@�@� �H�a�d �-�����7 ��B0#A(dhB�$ְF�(6"P@�.��+b� @�
\01Va��2)$��C, ��P�h��@�@�BSFA!,Yp%1J�yv�D��+
���;ޝ{���~~�                �uQ�2�ڵ��9�:��6ªQWK�[n.�˹=#�W��K������_5ի�����X�c54���Iêmm������NгV�pX�ڄ&�`6s�dDv6����N�n8�Xf�����o��b�r�\	�܆%���ٓv�m�O#�+�oKU�րm�h�[[l�p���g<=Y�ȵv�y�K�����y�EuSfw) �벍j���lc�=NX�n��ˀ�X�ښ�;j����<���`z��>|5�'���m�d�֧L��&���;h�ͱ,�t�Ѯč']*I2.@ $��v]���m�\���H ejU��۲5O\6v�r�\f�7\���p��� �5Kv�kuJ�������Y�v/+i0<�ft]��� �4��c99�v�6f��5�VC2꫑J����cE�9�T�9�����7�~<<Q������y�s�).�G@Bp�ú����7dfCh0�l+[�b%q�ѣN5Tj���e�F��;*�^������ᣡ�7 C[n�*�{T�hq��[TQ���lsm�V�}L��LO�/�V�!��vۃLv����u��m�x^�ְ�a-��+�q�K֞M�릨�![�w��=�<a
U[��z۵�tI-�\kgN� 
���!����H,����RN��ț ����u�P n�K�ʻ-�4��(YI%dI��j���HۖT8�'�Hmy[	lm�`.NW�����:N�E��S�m��<JD�R���j�,�+�;*��ۃ�ikĥFG;.K9�;n�j�c�攺s�6� W���;+ջN2uSgy`��/P+R�*� �kk�m�{jVY�e�WW���@\B�p�q�n�@v��R��S�I�Uږ����*���x�6�����TA:U��)^�Ȣ	Ey�J��iG�uqV;kn���HWY�kX�@��O� � ������Eh`*��������@  ��:hx{Ւ���<���B�9���܇]AdWb�n;Ny������t��r���t�S�5�)�]�W;�+]$�btf:	x:	gyxR�;U��Kv�
��Y���H�Vxݭ�w�^#��N4��kF�\�7��#q	'N�k���&���O��^'��kH<\ʝ�,��v8�н2��ů#��z��G��a�����{��~|h��Ѯ5�Y�t;m��pj�}����74c7n:J�F�#z����w�|��L<8��F����;�Z���z�h�w4�U��� HҊH�+�7�I$ٽ�j��޵`f�k���!DD)����Q�%'2�jl�߭X�����"!���v�wM��ɺMJjd��I6�h�w4���<�ס�DBP�����竧��h�TUJ�m �-��>�<�|���H����jx6[n<�]]u�/m�$���+�8��^#���u��u�8�1��s�ўٛh[�8���H1�@6��q����c��n=�]�������%�(�
���Ձ��ߝ���ٰ3�K�H��LrH�hw]���.��z�h�R����uJ��DBP�B����ߝ���~�76Ձ�u��yW#x�� HҊH�[�8���H1�@z�^�4|��i�����+�룻V�\�G�f\�s�ʹ��ۆ��(�5���θP����V�6Ձ�9���J=!��~�?3��$xG26&�m��>W�h]k�:���*�:H�BBG��Vl�盳d�Q0�G�C�� �FD$E�! �!V@K*-P@�߾���빠ya��bpX�L�x7��!(_�S�߿M�߻��ٛj�͜�`w0�r����#M���w4�[���/�-˭z�}]y����3"]����{m���7���)84�+�>[��m������b�)�O�I�����:��@��^�׮��U+Px���-�+6s]��P���{���޵`}�w4�U��ɒ4��-ˤ��*G��r|�>�����&�1:RRs-�M��	({��+7zՁ�9���DD
#�	B��ڹ�=�7J���s#bm&���빠�2����+���:��������I�5S�W@����K�(�����&��d�yI�D�4��s4���<�נu빠}�w4 ��A��8L�x9�`|�vo���֬��Vl�����k�n̌pcn=���4fm�?BQ�N�<��l�:�uMȤ�LrH�hw]���.��z�h�R�'��8LH�)3@��`~���t����ٛj�����=�t���v����� 6��r4Yi�=Jg�sò����98�4r�Ӟ��������^w\'[� ����'5�څ��!F�r5�,�4%u�X،S�p�6N�Y����;y���w�뵾e�0Z�N3&.9�g��n:38γ<Y�Q��Bzۋy�v�jnQ�ݮ�+�P���pb�f�ty�[Yrs=k��=g=�rr��M�v��(Yn�f=^��ݻ��33���،B�Inű���ڣ�6���^�ػfN�I��:�1e�v�#J)"�*����z�hw]����������ƚJG�u빿�?�#����_��Z�Z�VZH���� �I�3@���h_U�yu�@��s@���#A	�!'3@�ܴ�ɈT��߭�����Ѹ�8L�x7��ֽ�]��빠u}V�\���M�!L�)��f���� �/kn�������_Fx����ao\�ڡ��ɉĆ�~���4�����Z�Z���{�%"�	�2I$�`{3m_�#a/⊢O~v>��l��Z}T���x$��&h_U�zܘ�q�Hn*@;�����W�ESn�U;P�;�6���6Ձ��Z��X�?�d��4�R=�J 9�� �9h[�tswk6�����V�J z��{8ۑ�83�e�;ysŕtm>y�fB	�Ɖ	d�2&�nC@��ڰ3g5�<ݞI|�{k���<M0�$"������.��zS@���hA���q,n%�n-盳`f�ib�P���I@(B��B ��1X��ꀛ.�����?�h�� �����Uϧޤ��H1�@zܘ�|"�	�2I$��}�w4���<�נu�M�c�,Q�dOq�9.��mC�n	�ggl��i��8�r�b��q���4q4<C�0DiI��w��<�נu�M�빠�F�()0ݻ��ݴ�Ɉ���H1Š}E����LncM%#�:����͵gBozw����`}�n�R�$�L���s4�����Z�Z�%����ٙ+��hZY�0�$"������=nL@8�7 ?�U~;����}��WF�p�\��GkĻ��7�����|v�W�Ǵv�,qs�=ݝ�|�k-��m�(�������T���������'r�n=�]����d����1 ۹��Kݽ�6)UUUR�=�����vt(o�{���߿nh�R�6���S#JL�:�V��ֽ����]o�f�~�W�#o�H��H�.��z�hw]�6s]���!$���|������V��ɂ�<.�]��[�u�paNg�[�;�o]GA�[q�J+h�65�lb[f���ǋm���S4MoV���I�Q�K�vv8�d�5.��͍��l`��c�O�l\��&�<��g�]��+&kQ�;t�OW�v�Q��//2�zn�pk�4���c�,먅������쯮��Ʒs)�*ޞ]6om�mnj��hӹ3= _� ��浮xX�y1�\S2OGK��p�;n�[��<��pܻK�:.�,s[ۍp�.
���� 9�� �Ih[�0����&��S-���`{3m_�f��;�{���ݵ����x�UR�UE:���6����@zܘ�rEHn*@y֢�4I�"�<�נu�s@���h�_���[�+��N&�T�fjl��V�	,���oOr�<�נ,�ݬw��q �B'Ѱ�ܓ�v�sv����웋����Wþ	��׌��!"�	�2I$��L�}Ϲh_r�}�ۚ���4I�$�$����*��,v(��P����́��ڰ=����I(M�v����N�&$��-�~z[w4����ڴ僧���A'�H���@sqR̒��& :a!��ur��T�nfiX��V(JoWs�+���:۹�}�(\Px"I���8��m��7'cĴ]�j���r���(��H�H8ВNf��ڴ.��m��>����Y���nl�!��m��1 䊐�*@9�Z��~��Ď����n@P�6��/�߷4��=�f�4��GK��0m҉�j��1Q�ā5����R^q�X$P�� ��}�8Bʻ!��_|$�@O@� �QM�҈dM"{@0��bh� 5҉=�(����OT�}=�((��
�
�I��,ER1$���5|* x�g׏��>]��ܫ�AH��L�I&h"D<��=���������u%m'�y&�Rf��ڴ�g�%������V��j���jvj�7.-��&���/=�/8݇���8r����b⤉���jn�N��Y~�~^�H�������>��Y���"b�I�R=����u��:�]�����/�%
�7���R�r�U-$ۙ�[����uv���^���� �����������uv��۳`f�ڰ��$�\4�DRJ!-I%����X��rt�hr�ӦJ&��?ń�D%��/��޵`f���m�?����qg�`�V�p��m��9�݅�)���]c�S�n9n���^�Ffn �R��H2K@z�נwr�rD�Ra2�I3@��!%�!$�&N�?�;��6n�줣���$��L�:�V����@�n���w4�VH��&$��Ӱ>~ݛ7vՁ�fڰ��B��DBS߯��`��'� RRuCr���� ;�T�s$�����TϮ}�  t�/2�v��Ʈm�ٻ��}���Wm�;=����z�G\�S5<sW2t围�^�Tm�W���7(�A�nf�/��$R�]ٶ���CYmێ�/-���ٵ�-�c�'^�tn��c�tz�ݷ/����{��ϰ!Oa�:N�g-D�#bX��V�+�����aV�[e�f������8{;�U\�۔��m�����|�7�,�P�p�t�÷���ݪ��e�[�p���Tm)u�<p��n��z}�� �Ih_I�$T�#�pܔ�A46�4���w�J!$�<�l��V��j��5������E2Q5N���vl��V(M�oZ�7��-�ǜ�A8��&����h�m�6w]��P��;������SR)0��$�I��u��:�V����@�n��>�\� Ʋ"bm��G��������K�{��gS�X���+u���9ՙi<C�0Db�4�ՠy}k�:۹�}�]� ���&��	QG�r��پ�+�����E����{ʐϕ �- >��4���j�K����@9"�s��d����נ}Yh�ŉ��4�r�u�@9�Z��b� �\72�J��c�Vl��%ӝ���?��s@�}��G�p11���6k�$��ݙ�u�q�����ܼG"A<:������&��"E�yu�@�e4����ڴ�y����0P�F�@96o`�s$��ɋ����ϭ?-��I���$��@�g�@�����D(�J�J"�=��7+K�IG�y&�bp�:�V��ֽ���>��M ���&��M�u4��ń�B����3V�Wj�=�Q��X(%"��4�Q���ճd�r*����×r�v��]�Q��5�28�x��@�e4�:S@��Z�Z���G,M�̑����9�� �-�rbɰ_~�ߪ��?\����K��?ߖ��ֽ���>��M�<�1D�I�E�a�����1 �� 9�� _����h D1A��>��}Ϲw��w �Mɂ��7���h�Q	%�DD%���ǀ����>y�6������/3�Kکy�����l]�6��$�������td�v��Iڢ)���Ξ� �Ih[�M�������<�F�8h]�@��^������YZ_舏�""�~��U9�D��D�QŠr���=�����u�?��~Z��5a�3&)�%#�3v��=�+K6w]�B��;�6>]�Ԧɖ�*��3TXŕ���%�ޮ��{�6n��J*{5�����nvΗU�V����1�۫n�Yu��\
i��λm�z��8���%�u�ѤS�)x"�lG7n	X6�mV�S�klR��skOb��&J�z�)77m��m�["I��q���6Œ���ڱ�`�X�؊���tj�'0ɺYvI�vⶻ/5��[jN6,����v��Y2���/93����kk�K�J/"��F�?�Y���)�VjN�#�
pN�o���I�;7K'�Ür�c�� )��qغ�ӕ�gv[�n�zڹ-/j١�Ӫ,��;盳`f���%��u�?�yLQ7x�Qr-盳`f�ڰ=�+K6w]�""��n<���nL&����Ɓ�fV�~Q�&�'��{�6سK��QI���#m�@���4�h]k�/t���U+Q����"5��@�N�?$�B^������,�,������`��+Ԗ�\	Km��Twka�d�W]�rn:��=n��`[
��ܴ�$��-˭z��>��M��Z��:��/�a1�R=�Ji���ؔP@����d���}7$���@��^��h�Ć�k$i4��ei`o�u��(I�=��k���F�B@pI,R�ڴ[����=����w[����L�x9��ֽ�Jhvt��~v� �UYH�6!L���n�ٚX�]���m�SHv�\hf72fI&�����L�0��Q�6n�	�ܘ(L#q�����Zݝ)�_��@��^��Φ�
E$ɒ7���=�vIh[�㖀U+S<lD�"5��@�;V������؎��#,$�0�HE!$ X�P� �A�����W���k|�f�z}���'>��#m)0q
(��<�נ^�Mز���$���`���:r8�TYW{����:{���#�^�L�$5#�cP$I)�+���<�H�<-v�-�8���^}��b _��{��ϙ�8m�d�&����~4�h]k�/>�@/eT������X�4��w�D6y�t����b����k�K#q(dC�ȴ.���U�D$�Cy�k��{����f�C�s5I�t��������u��`o.�Ł���`סBI)�f��b�&��ԂY2FӋ@���4�h]k�/>�@�X� �"�؛�ƦamѨ��ĽM�)�&)ڀ[�n�Z���CO @�s��I�#X�4�h]k�/>��(��DzCyu~,?s�US2��:t�i�<ݛ��&���vj����N뾄���UM9i���JSuS`}2}ht�	�%�=nL@uʐ͔ә�QU-˩�a�$��[|X����n͇䒈I����ϊ�h�T	%�C@�;V��}/���?W��{��{7$��*����
��W��*
�APUЊ���DT_� �*��UU��*�`�E
� *� ��
�`�H
� �D��@"�@H
�@��@*F�R"� ��@��E��EV
�U��
� X*
�B"�
�A`* *`*� *��A
����A��A��B
� *�E�T_���*��EAU�
��PT^*
��PUЊ���T_�"����W�PU|PU�b��L����5|�C� � ���fO� ��~ QT         �*�       �  �TH�%TJ�P�J�(
�U@R����
Q@� JH� UR�� $� @
�  ��� � �v�rO!��G�^�Ϸ�� �>�=����}���ҜGU� �z\m��s� �#��g��)@.}as>�=y=:�Xp��/�6�����w}��ǴO��^  �>�D����B�Aݝ(}���+��Pq��c��� w�=�&�j���<}���8<�r����g���G ��b;���s;���s� =�*���s�����Z�y� ��QUE �(U� z�f{����h���E:l���qTVٝ�r��.YJ3��$ӈ)K� �h)�Ҕ�;@ R�;�)@�e)J]��h)FvtR��e)JYe:h�;:
Sp
�JR�l�JQ��(R�&�����A��P ! ��Hcb��)JX�4�3eSH�_ms�w�}� �
w8r��W��2��1�{��9ҙ�޵l� m]���3�(��1eF{�%�]�4� u������bg�O��$�J^ PH
�U UHce��{��]9�.۞�$���\M6y��7m���� ���Y��\f�  �q�]o{9+�JgC�=�}��t1����s���x����=�{�u#�   4���2���!����S����RUM4�&C<z�T4�   =��I���  U?�	S�T�J� h ���ʕ	� ��|��=���u����?�����w�\�s��@��CY� (�� @UO� U� (��� �� T���������M��!
���Z���$� �A��@c0KR��RB �B%i���хkd֥�D55�B�p�����sI.Ȑd!�
�i��.�@� D���DH@�`@�H��5����-0��ɡYT���/_hi����
���Np�6�0־eYK%�qaWf�ăw&3Fa�n
���d\7�����dNa��)�5aMȣ|�C\��ˤZ�
�N�T�{��&wLeI��0����P�����pq!ФB��"���#0�K�߷�k{z�wXl�Ab�@��-�j~��BOĳXT��aR2F�$B#aX� F1B1�w��M�7���!��dj����`�P��+�)��<:�D �$.���꿞h�\�R� }"�� ��8jIi�.~>5sX����f�aX����aĉB �C=�E!q&�%�&�&�&�L��w�5
R%m͚�������d�D�"�1ѭٮO�B�8�)�~!��qcX�GL��0���anФ~��
�� �1 ic`�~a�4!K�r��\T�e�����mH�6h#!�5�P�(f˓_q �}��Ro��ƤB��! �$�!�3/�����X�+a1�R\����A)
`��5�!3)$�f0	1�C"��oz�����ۿ�ϙL!�`S$V&p�f��-F"Rd�	`��@�E��*�q����
l��6�x��)�: l�����HF�$BksqN?�0`B�聲s�k����
�FI�+�CD6<۔3p͸�np���R$��		��B;y�FI��6"�0xM���c�7��̑��I���7y�?1ha������q�	\�>�@��1X�(�H�3�����{� %$���H2����)���b$�`07'�`p��8aw~"�� @?$ �!m��W�1)� �"`��"Ap���M��c���75�f�&��TL�@��"��R*U�I�5���v\tl6�R;����%�! �l��?F�:vp���0ю�����t����a��)qӁ���6K��4��Y&LIfHØV4jB����+~���$,���)
!SCF՗$��ЁR0�$6��5���B�sG��Ip�
��?h��:n�$����-�� X�B!X�c$��j����\�����۫�J8�d,(�$�a`B1�SD`@d�w�}���?k�;>=��@�H�)�E�w(��Q�>���H=9$,�CA���bFP�����@��B2��~���"A���%���s�ݺ��>u�I,
0��#I&���$� �B�ߒ1>�ﻏ��W���.�Î�d�XcBb@�� ŉH�P�XP�!+�AM$"��f����h�/��~a���P���p����.kY�����4"W�����й��Y��k�?��$�!kF�۷��湟��n��0��q�4�bH��O�!@�o_������ĉЂ�ae?s�����Y��/)_��� �nfow�s�х����ħƑ�@�$"A?+�āL�͝@��Y��L�R���d��ab�a$�#R�80!B�a��P T(��h`X�ԕi����P�.I�tv�!.�Wrsl����1�7ċCd ��k�
�#Zd��-�kSFe��O߫5��Z������f��.sZ͜�r��:t��� ��E"!Go����;`�8�����D �XѬЋRT����j��e0�3;3{�d��I��������I��U���$3Dc,e�*B��}g{��q"SΡ85u
�g䌬�+aO�h��Mf��%u�	��Tȵ�I!\�����0epH�#2h�Ma:`Q���"L˨d�B+��U]�Cc"W�w�����rI��Mp����E�BD�RF%�c�@�����r��}�C�s�T5ߑ�󪏭s�S5��%Û'���ƻ9��\�	��C���QJ��wB���U(�k�jS�D�`p�Yf�36oA�b\9.���h��5?l�&�h@�F�.B�HI��,.,�ļ#r]o,)VD�p��W"`FX���>�w���	X� MO�r���	!�O��bU�1!@�D��i! ��0�Ĭ���I�?�8��|7����}���k�4����n����i�$)"��|��e�#�i��h����J2�e�n!�ٲ2P�D7�N�NN��[�W����	T�i��
&�����;0���k���f�c��vSI�&Ԉ� �@�4��f�xF~$$vH��[�d��8j�a����mJ���xh��Ç' M�ĂS[��[�k��`Ġ"�h@"8B)�@��\A�6�i�@�&���t;#0��#tH쐉!(fM$�޷c��B&h��ԛ,�f�K#����>#@�F�c������98�6������;0XS���L	�pX4q)�ٿ�Ï�5���k���m3��p]3}��l��;��������ػF5�б����٣�Ë�XA��nI+�ӷbh!�:7��;1+�6K�hv1��k����, B�4��r��kf�WQ�i����6h8�)����m# �a�a�#�0ӳd� F�&��C)��ȑ(j�zѤ��#G;jh U�LH65���7[Cpw���h������H��R�,rVZؑH%Ӵ�F$ �4�$`Y"P`�JA�BB,ClB���?\ծ��p�6ʹ����c����6p�ƙ�o?sT�~��T���A��*P�� �6 h D�U����m2�u���$�,�ۛtH�$h��T�Q�bH�  !�F�%g
d��
�����z�FP�k���F���L@��J�V)�1�$�1ֹ�HW!f�P,*��fI�a�l)�74����%�kmv�F�-a4mْ�4)0֍�6R2+��-���$ ��B 1Zį�R�FFh��e��X�B0� �4băX�c!�i�����"H$�e
��Ӵ	��1HA�d$,$so"0�$(�t�xr]l�k���+�цB�LÍ1$3{C��h�0�q�F�D������
bB��\ �S��P�l����aN�����f��~��H��~B4z��K����F#���              ���                                     ��                    �� �`            ?�                             m�    ��             �m���  ��@l8�v�I� e�e[�m   I:n�-�  �� �ܝZ�&�� -����ʵ�d�eZ�UVۀ7m�-�[�6�   m zմ p�	dI6��#���}{Xe�o�hp�C��>�U����� ���f�yt�mh��UU*��*�+��U����zꥀ�2���V�
�%����N��Xj����$"M���knh h� :��F)F����j����V�-��Wj���m@*ʵU���i�M���l lt ����Tr��[F �[C�O���  ���浛m,� �q�β;��5��cL&MQ1Nۘ`��.���l+��2���6��P6-Č  4��Tյ$v6�M��-����I��$�ۉ�^v�Zt��h�� �5���e'f�	�( 	�3m�9ڶL[A;���N�� s�����U,Bt�s�F�<�UJ�@�jWh �UW*�/=Zȩ����v,i��E�`  �}Uһ��<���[R��P��Nm&�@�uc�[�ny%X(���k�[f�e����,m�	$tM��o��rE��i�[�*E�`�fn9�{#[��J۶^�n���(ԅr��H����$ � N�ݐ`tr�U�*�K��`K/� ��E�ڶ  ���m�	 mM�]������А-4��v8���ERom��-�:�9���n� p$ 8��,���=��#���f8+j��W��Ie��&��![`�����+�۞$�4��`2�؄�s��mSmu]�N�am�H�t�n�
m�l\�`�½9亸
�6N�]#$�ۥ���g���:D���n���kX   ���d� ��	�	��-P� ����`m��m� 6�.�& 'I -� 6� 6۫ی�e�Ah%*��             ��&  [[l  m�q"�m���I[[d6��$��,��)��  m���1'n �����8���)]ٷ�nUz����u H��lJ�6�Kۃ�m��T����/Q��&ݤ� �[����M<5�p ��lH^[h� �.��	6�@M�v�	�[x�ַ@�e��9�
���mQm�yi������2m�� ��倕j������D�Z$m�7Ў5�R2m�m��I���U]8��Q�p�`  $HqT=��Z������R�6݀  �Sn��x���R
��+Z�� \�@4u��lm�&��GH[V�GA�6��[�k��`[@l.��m�N�k�K!� ;rIf�nC�mHpq#n�z�[nYe�����[A �Ӧ�l�ݐ*���mI�����I%��Ͷ�r-ać$ $ ۖ� ��YZ����U�U������L  t]�` ��ms�Mnl6� ᴛ Ԝ �e�� �  �m�j�^�pZ�����W�UVU���}�F[N ��   [F�8 $�7m�V�  ^���sz�t���I��L  m�      -��m���D��[�  �        �V�l-����~P    -�$	��%Ҧ[ͭ� 	 �  �a�-�  ��m�Wa�*\r�gEP �`mrڑͶp     �l[Kh 	     �9���m�''_ �  �Z�)�D	_��֝�6��r/[mg-��%-�;^� ��	�
��Yrt��	d�� �.�   p 9,�[A!%�m�m%��Hm�$�     ɷm&� [�^l       #����,�B���W�]Vxk)eI��m� .�m�Kz��'8��N�&m��  e���*����Ьl$� �  m��t�6�n�]]p sj�  �k��b�1K=�ק�ܻ�c 5@     �۴�l����n^��ݼ;m��K��   ��[� [D�  r�n�	m�ձ��Ig�s�C�]Z��.��
U�U5�9CX�����)@ pX` ��$        m��   ��M��ɚ�  ��  -�o	M��l�ֶ�8�$�A��[Kh8� "M�`   �  -66�H[d�� �-�@m-���K� $�6�l  �:��m�e��H[C�i�$8&�$ɶ��[m��$�@l����F���hkoi ڴ�6��i^��)j�6+R쵌�^�e1oRAi�� m*�A\-U@.̭P�o\ km&-��$����{l����T  U]U���V�    82H H �mѢȷ l$��i�װ����unlm	-�Ým��R� 8  �۶�hK�  �\PBYu����k"�Tp��Ift�#Y��e�����ۘ;q a��*��]��[�NYƥ�H����>����BFݰ9I�im�q�� 6�� 6��t��+�f�  �v )E�C{l�  ��:nӤ�b� 8*�i�m��`�6 ��i1�٥�6�$ 	�\%��lQ���ej��*����6�    �I&��Y/i��n�    ����~�o�%�[BF�V��u�rB� �Ûm�p   ��&�m �!�8�m����@4��  [�`    l�  m�M:��8�      6��� �L� \UT�J�1l���� $��u�� �`�r\�g�� 6�6��k�t^��\*�eenVU�e��� -�ڶ -�-� r��t-��E��6�	 I�ۺdQlsnؽvum�Ͷ�m�m�p �m��ݱ�u�1zݴ�Z�  hm� �@���6Ŵ�f�.��G   �nkm���g^�2�U��(��  �&� $$��~����!J��uWUp���@���6[EUUHl��F��VU���I��K6�3 N�
�MU.�||�QmX��K-	 [P`$ �j����SI�UUAK[P�Z�g�UW 9��p ���lm��s��'J]�q�   �5��om��)i��^�����	6��� �
�UP!������_HO��\ 4Y�$H�"jB��P�K�/At��ی�5l�U] ˷\��[9nNP�k6ے HkM� ���  � �@   |M�`    m��I��  ��hU�6��m�kWi�  h�8�-��� ^�"�ճmgh�H�m���:��v�Ԡ�6�aC:'YAz�y�d;a�P�e���8N�IiV�a�    ��ו�e�bu� �   k%��m�D�\�iV�]@�`�-�  y�l��i!ƶF��    m�  s���� -���,5���S�����Ѩ�@�a9�����-�l�b3E���Q[4H��-�  l�hp m����p�� G���෫m�P�]��         #� [V�  v� H  $�kz� Ƶ�    � � 6���X   mA �Ͱ  � �` �   �  �     6��	 -��V�m��� �:@�u�&�ā�mؚ�V� �$  䉝�B��;1ଜ��<9�%��Y�y[��):2�f�\@/Z�[d�i 8[m��:h l���ݶ 	�� m�mp�i�ݰm۰M����+ $2�m�$Xc�i6m�O�m��ĒL�[Y� �m�   [v��Hm���� -�m� [@ �-��C�qm����F��4r���P MT6�G���{����{����wp D�$��Wb� ����L|���(�
��D�G`���E�
f�
,ND~
�A~J�D�A_�W�  �5�#�6�6�׊&�Ȉ��|��_�#PP���A��� p���!�p�*��U����~I)P�Q6
���"^
��0_��>?#�/ȄB,�:��؂�X����ʂd_�U
��	�>������"�����E(����������(q����
&����D8tv��Z" <@O�;� ;
���~TTÚD�
|��>H�DBAF1aUG�@����\BqU�D"A��D����h�? �b*�TM*�ϔ:
��@��ʈ�&�@�]���1���q/j�D#�$C�p�� ����E�! EE�(���_��  m�      �m��  l� m�    �$  �5Y'[�M:��W�2tuT� �Q �;i�%�l훥�AX[��r��T�q`Ca6�T6�j�j����n��F:� ��8RGu���,P����L����W��+�#��|:jv���N@�x�<�Kԓ��06�ڦ���hg,�ܔ�:Wrbe�,�,��g,�9�P#F
ay��X�D��޵U�le�F�I� @ ���  ��I1�+�.aڱs�<kGW����+�QD�	QS���\�A�K�D$�ɋZ�\�*c�8<�J���w2KB.��dz��J5�[ed;*�ej��ڞ�A8%5�J���ꨁ�	p��p�r�`�+�t�說g�eZ�t����t6:Zq�UH��v�&�����Sq�����2-&�+֐*��i�nV��\��mUI��$fq�Ws��q�����P3�۞���m���2�;��(��Om�Zէtۤ�m����m�̃l�\�5���
�*&hVWOk��nd�t�R��gF��EI1��tIΫ�٬Ky9�/
P!7, Ң����bzC�b㣶emi6]X5�ڵ;sR�8�0vv�������(S�|�U��ZX�UڕA��SUmQ�AU��xVj���ǎ.-v�&�۠ze�v���n�eB���ـf8��u8�oa�KYhӪ�9�]�jW���{q٢n";%ϭ�*��՜qU����1eZW�p��v��)ǅ7X��ض�m�YVڨ8ڕm�50ѳ]�7`�&SK;)�y�\a�LMV�-�ՙI����&$��\P789�]�&�Z�S��J�ۥ�1�6���ɺ]6� U��-����0�jU�m���IH.�B���3�;h��c��L���Zl�	_7ڕ[r��xv��v8��5b9��g�n��w{��������X,Q�
|��(�@)�%ʪ���YI*�%Tg;ww$�HI.I*�j�&�:r�Į]n
}���r�5�[L��C�8ȭ��!44l�r\:3��h�-�J���v����M�#Z���x6�$�G:�a%6�5���f���r�"p��δ�gi��I�N+\�8k�(��р��b˹g��z\J���"����ּ��[�M)�o<�E|K6�8ے
�J�{�w����w�ޜqȮ>��w.�e�ۓq�9�1��������I0X�<O�܏!˺���p}���Ԫ��fl��2ރ�$l��ܗ�3=/5R��T��v{6p�}~�����oR��#$q�#qh�e4׬�<����uh�َD�qI�5��z�����ގ������^�hm���rH�H�rh^��z:�޲���h�	*��1�(�k&<QG9�7<T�g�CTz
.SNM.�aw,N)�q�8�q�H�z:�޲���h^��T��s"b#i��d���voO�"*@i!A`�&*!�Sj�ܓ��5�'��������@�:�HƧ�lr!�h�Y�y{��-���?z�h�`��L��M��^�oGV���S@=z����%A<�$G������]_}_}��$��G�/�x�����?(�sw%"<R9��֓��s����K�J�Af�uÖ5�V	�������JF��?z�h�Y�y{��-���9u�$���&H�R��h��t�II��-�qaU��P.�c�����$jG&���@���I��R�*�I/�*��& �fN {2ۻ�lq�����uh�e4׬�<����î4�D�F�I����S@=z���^�oGV��a����{*7c���x�q��^8[�3�6�̈;qQ�j|������俣c���}~����ގ������u��ʢ��Dln94/ux����[��Ē���%���|"ԑ�Zwr_ ���|��Ã���goY�y{��:�F�(��	iH�|��À�d�}�_S��J����������@s��f�䞾�8I#�L���4׬�<�������}ܘp���~�6�4Q�u��ݵ��K=;�#mt�����2���'/�_}�����{��}�EŰ.�Lx}���3=/ ��0���|���� _�i?��m�8�bR=ގ�����z���������0�"6�N8�޲���h^��z:�p�����D7����ztx�$��pĖ��ė��+q�Y.˹rpz���jI*��^����Ӏ�d�J��I���n�V�`D�D����V&\G�U�b��:�I֦a���w~��� �� 6�v��em(�k�윒�Q�1;u�8���]�0]��Y^�����7F92t�Q�m$��k�=����'���ζ��I�{t��݄������T���t�7e�):���m�Km������_Z�7���[���%�L�-�u^�v��D�i�dӋ�Q�3�ޔ�ŋg���XI����;{6�KUd5�r^.�g�l�*E�'X�gI�&y�+�=�K�然���a"�V�]�U�ql��l=Pi4Tp������h�Y�33��*�:�F�(��	iH�Z�e7�������w��Z��@���@��p�
G�#QHh�Y�w>�@���@�l���݌�I�$��H��;���)9�1%�8�"�=:<I)�I�lq��"n-ގ������hϪ�>����?��9��C�㊣T�w[pZ���0�7��y�N�j�V��$X�s�#i�������f����ގ�������֬��ܒ~����@��"���~���$�z;�bKdqa�/tB*["dln94��h�uh����p�z��$l��䏁�K31}����=���@=z���Z^�Ԕ��	iH�Z�e4�?�>�??$���bJNwIl� ��S�[�)prLWOP����Z�i9і-ӛ�!4���J��I��~�?����Z�Z�e4��dJL	$v��K��{��|�I%I�w%��|��h�Y��%l�����������;��n�%�?U%���e�N�~��<��^Ie�Kl����-�j�^�@�ڴz:��ΤRbp2691��z���ՠ[�ՠZ�Z�`ڢN ��@�5t=�N��숱Ola&��˛�Ӯ�a
�G���r�}���!�)9�1%%�bIztx��(��<�$F���@���@�ڴײp��|ڪT�f�m��6�HIrڑ���|�׬�-v�ގ���1�H)$Rc�š�%�_���{��fz^>��W�%V�RJ{$��:�����H�I�M��Z�Z�e4׬�-�Ҡ�N`�sY��}���{�۹�Z;'#��m�d���2p�l�9��@���3e�X�m�'���e4׬�;�U�r����F�4�qŠ~�S٘�w��Z��@���@���E&'#c��@^�$����)9�1%�8�%�(K+�!FF��@�}V�oGV���$��G�-��"E�l�1�`�uh���^�@�}V����g{ӷ���  6� �Yh����i]�����ѻA�5�9��6bSN����[M̦�j���+d�퇐1��*��RO69z��<�u���ᵃnq�ٺ�a��G5�9�J[uո�:��r1-lmg��7gt��yv��!Q<� �[]b�mԣv�r�`������5�IٰQ�f8.,�G/e�wnY�ӄ�WɘG��:�mN��#:�����{��{���~�p�.��!e�.$��mԮZqͱ�-	�W�Y,L�qXQ�g�2�!#�)�����O��f����ގ���1�H)$Rc�E!�%���K������[#� ]$�j%&�'�E#�@�}V�oGV���I7�{��������R�˗䉸�z:�]�@=z��j�9^X�s#x��m8��-v��U$����7ou��K��3/���@�5�K��v�N�Ș�����5��nGn����f�65A�{HV����$Z��h�V�oGV�k�h�q�5y	c�K��\�2�)�J��A��g{���rN�;۹$�߻4uQ%A<�$F���@���@�ڴ׬�-v�ޯ�F$$q�#qh�V�z���ՠ[�ՠy[f8I$�Lq�8�׬�I*ݛ��7r^��y��jIR��?~��0��y����j���k�Ayʸ
�z$��sjuCl�����F�� ]�E#��|��h�uh�V�z����V���pnH��@���~I%M�����͜2� ��5y%�doM�Z�ՠ��Oe��c��H�E��@�Cj�T.��8@
yQ�X��T�4D
 h���M�����0D���U^��BaB�
�3W������DJ�@�JƤ
D $ ĉ
�B�#$HU��
�6$c��@pQ��] �Q"~A��ȢQb��E~EGh���T�y\T�04����������|R���{�q\��v\�܏��URT߷6p�ݾ^Y=��=w8
����]�>��R�ۖId�IUs�9>v�_6��M�헯�ԩ$��� {ٳR���?$����o�v�x	��s�bIh����Sn�(mz� �e���[dnN��lG��z����I&�ٲ�>�[�u��f�M����|��m���v�$$�mܻ��n����IRl=���7ou�����_}��"RH��#�@;��@��>���|?7�{��n��.[$A$��E$�-v����@�ڴw��G�LTU�G���7v� ��V�HŎ<Iț�@����=��h��hψ��]��2`��x�%S��B�ë�ڻbzݪ����q�c��"����xЊ�d��CK���%%�bJw;�$���D�7��ɍH�޶h�V�{��@�ڴp�1e�F�jFI��f^c��K��5n�����9��6{5�M�Z�m������[�������m$���ݜv�^���nfڻ��d��-�.��}I'�7_ =�٩|�v�_繜�| IR��͒O�>-�m�m���mt��[��=�����7ZG��n�h0&Y�.��tkL�+m�I��.�/:�Vn�p�˴8.y0�74���:4e����uЀ��XX�@���;S��:�z�:���g 4��	E"Wa�׍���wYs�;�/Zr'5Cv�ݑ�t�S/N���E#�rL^��\�3�5�v+��lA<d7���~�|_e��%χ]slu0��q`�۝�n�g�`
��U��2k�Q٩�S�#/�o}4]�@��ՠZ�Z[^��&�'�E�@�ڴ�Z�ՠ��@?rJ�I��䉸��Z�ՠ��@�ڴ+���dom�8�]�@=�f�k�h�:�
�]H���2691��{���j�/tuh�V�~~?�����%��F��kr��TnSq�x�w���]�&������n:�IJd��4]�@��ՠZ�_�?��?� =���=��֧j)-�� �zgn�x1�@F.�=��� 3���f^c檪M������!#�'�@����@=�@�ڴz�4+l���$Rc�Š�Y�Z�Z�v�ՠwuz�D�H�9���ՠ[�a�Z�Z�{' ;�m�U�"���Q�.�q��v�u=�/3��=s������T�g
�F��rD�Z�v�ՠ�Y�Z�Z����1G�m��X���1$�tx���1%'LkP云9��DlrcR- �z��jӢ�|hM<�}�7��'g{w!���ŖE��$nM�j�-��-v��^��/��y2AKdrG�3=�� �UU�7_�u�m�]�@��J�C���M�R4��➮�+=ngX�"���'�#�"ƺ��N�K�j"BGI��j�?+���V�o]���m��R5$$���qjKI��%%�bJN��$��Iwq1ȉ0$�<rD�z�ՠ[�a�Z�Z�z� ��+`�m87$N���#�f^c�<�_�UJ�����2Y�����F�6Ĥ�D��Ii:^$��Iw��X�^�B0�x�����G�!�v�Ix��+���v�%E��F-��=���6�.k��ZN��).C]�r�$��Io5��,�5R28�z�ՠw�\4]�@��W�{�k�Yq<� �DRE�w�\4]�@��W�Z�Z��S�n48��ՠ~W��-v����yZ��R5$�G��?+���V���p�-���$����� ` +WECe�8�N�������rv��NGz��O��ƹٖ�pn��nv�ʺ�i�S�T�a�tm���6��t���z�h�m���F��J��;;��YڻH6�X�ٵ�dscM���Վd�6�v�{s�֊�ܷ���'��-�u�A��ç^Hd�"JԔ�]��ٿ�~/Y�K�Ett:�H���q���1�+�D�؀o$��M�T��sD�2�T�Ӏ�v�G@��+s�H�Nά����}��7W SF\I��7%�������#�}�0���������or%�$�;�;������J�gwf��so�{��hW�;#��"&ؔ�h���׬�;�U�w�\4
�]H���dlr!�h��hϪ�;�.��*W}����o��5�9n]�,�]�� �}��� &E� �e&���n$���!�����I"oN[���q���su�	<�!��:4k�W�=��t�����t��A�ɑn���RIwN��䒯���D��!���h�v�y�ﳜ�̢��<79f7�< =�n�w7(3�_}Wvr\jF����R�$��)5$�t�n��������߿g����lV�M�][i���s�n�u�f fs�m�$���y��m���݅�,#n�m�l� ��*� 6L�tz:MI%�:�ߒH�`�q�9��R6�-s�XK�l��F�3s�y�p�ָ��X��AG����}�����xЮ�r ����ź �O ��� ��*� %���r+��.˸��>�����sR���	�n�K��Y�ɑn�{�t��E��$nRIwN������[��@�������9�m����n�o;�[��e���[#�?�m�U~�9��0I�n�/G���7@%������v�M۫0 �2-���x w>��_9V`�$}-�H`r�'=Vyѵ�	�ҶGJu����-ӛ�R`�]�dɓ53�'��m���� �}��r��dȷ@9��C�I"x�Ȥ&���W���*����*� =&E� �O p5lv�m�m�훠|�Y�ɑn�/G���7@qW�m�ui��!�� �"� ^�'�}��y�oD@�Vi�*�D!� � �B	#��,	D�Hȣ�����7����?���h�X�.X����q< 6��.�|�Y�ɑo������-`�a��LCnv0zr"�Wlb&�uɫm�79a+v�TH���6��x w>��_9V`�d[���� �vY�*
�Ӵ;rG�ͷ���o�UUUwm�w�}�m�٤Ԓ]Ӫ��$���=2"BG$r��dȷ@���~�͹~7@#��kRIy��9&�C�䐽O ��� ��*��UUU]�����6�^=��ˀI#�wr���ϡ���U� l���q<@ �~{����D�[!BP�`6p޴����Q0M~d�\q��@8��P�dK5�8�! �$`@� 0 1	"����	��|��������1��B
�C�t��ũ(f�'Q��2b���A*B��`A M�е�J�pBP4@dH1#�L�2�i
 B0K� B��1�ha��J��P ��X�F10D�X,`F$�GDhX�ᡃ,R,b�TLF"H� k.1R B��H���U��`��@�3ޓ�Ozt��t������o�         O�l�|   �I�       	 -� 
���%�@j�y[���&�D��[%�`�[zm@�˗d�ss�܃���z�j�f��ڊ*�pݘ�8���6<�1[Wi��(�
-�	n�M3+s,�-�c6�=W/T`۵hع]�m�FT�Gt�k8��	Լ��sB:6Bz��W$@܋��e�5�#�;n�Nʃ���ӄ)R�v�2Y�	�r��Y-��I�ooPZ\ft�Qf
��˵�l��j��]�    [��Fĭ.�"�l={cÜ=;k�y	�I� �F��k�9�-��K�RE��m��[q�$q"B4R6�f��/]�t9�W'jbR�����ŏ�E�έ�d�iНv�b�R�R=g9K@q��U���^��,WR����`��E %鶲�m�GJ�u6���L��
p(I�f-In��a�N��qAm�g:�[R�T��g^�����2A X25��_ r��5`+Vܰ���&OQ�u��D�[M� M�+=(ٸ��mS�I���l�3�UUR�R��K��Fӂt1�U���8������طJ�ņ�.[=l�����|V۳�x*�����:U�B��4��z��Ή^ÕHWNv�0��$\٥#"V\��gp��ڸf�H�`$7Z�MNW<Tү����6���8)��W)���l�4�7)�u��S�ˮ�d�Ҷg�=����]�vۢ��3r��l��_:V&�X-Ӛ�r!�g�]���������݀-�Z�5��Tϒ�#A��0ãs��.N��v��cfU�����j�n��)E�&�t휫�Ý��%Y2�]�I��[Q�Y���c�j�\PJE����P�s���f^Wd���h ^�*!�KM5�b�V�C��V�`*کgڠ�xŸ;��-��Z��ݞ���v����|1e��٠�s�<m)APQ�()V�/X��ww{����q�����q��v��D?��"��V�%�Kԩ%�~�I$�I$�]�UU*��!�����9��kv�s�q�Ж�-�k8�;rk��]�z���,�hr���]�;�{ff�]n8��nկm$b��K�s�����m��*�b���t�9�9�\J�(���(�}9�++�f�F9��q4�Iչ��:�c��a�B�ʹ�7e��gXR�c�a�n�d`��z[�}Gkqs���^��.��g�pq��u�H��x'��ȕv�r���9�+vr�J���7c�)m1L���/-f��F@)xI'$M��$��}�Ԓ_�ڷ@G�s�n�"qW-�m�ڴ�v��+�dȷ@G�s�n�q�R� %�tLn�ةݫ�mn��3 ���?��뻄�^ ���߻�� �?�v�~Q$�:�� ��� 㜥x l����0 �3�EA]:v�bt6��9�W�ɑn��3 ��� ����g�t��4�]8x�%���s)��z���U���˄n ��,b�թ�7n���d[������7@9t�=I%��tpr(��BIߒm�&G�"�)!$R�$m*B�̙�� ��W�ɑn���%ܿ����m�Wm�� 	�n�q�R� 6L�t �q� ���c�M��.ٺ�9J� �2-���`ު�Wy��|�c�j�廒��#�`7J� �2-��q< ;�Ct�������r�����ۘ�K��48| vx�Zް�{^u\�B�X-���+b��7j��[���� �}ѷ���oU/��}��|�~�q[#��۷iۻi����|�Y���|�gra9�*�Wv�}Pֲ�R�؝�t\�� 6L�t���W�Ug�Sq�� �>����Wk(t�ӻ��V`�d[���� �}�'��0���[V��7I��[�����~�4�r�������� ~�P�������v�ã��ms/9����a�{Q*�gڤ�I,��m�Wm�� ��� ^�Px l����0 '#V�i7m�.ٺ �r�� �2-���`�W��$+�x����F�I�MIɑn��3 ��� ^�Px K�.����Tݫ������0 �}���UU}UA�d[�b�,�5R2H܋RIwN���w�ɑn��3 _�
Q�߆ke�˱D�=�٭�Wn�m	��m�˸+�.�3����%�z^Y��+X�/�@!��� �2-���`����+��:bm7ce�� �2-���U݄��0 ����8q</>�Lp�)$JL!$���$���R��7@!É��d[��]�lcm���`����px l����0 "�$i��&��m�훠�px l����|m��Oc���]�T"��B�͒I$���h 6�����J�t�t� �&d��sOF:���p�爻1��΍s`m�sr��#T���9�O��x���ɶ��]�ị��[����e5�6]PӦL���f(ʰ�y�A��
����N���m�n��5��*�$^��{& ��:y���v��9��ڽ�{)�]���'�n��&�Y�!�b��	��m�<���{��9��I�]մ�i���)QR�mvN$Zݪ�Б͓��s�$E9���Ή\�_������@��s�}_U{��7�� ?_�o��E�S�b��� }2>m*���o2f��m�y/g �2a�=j�,�5R2H�4��h����e4wJh��*L�Q�b�-���@�l����M��Z��l��DHH�FH���e4wJhϪ�;�Z�]�iY�&9.��E���e�X9��ں!�t�4fY.���nYk+�
�'�O����4��h�z�e4η\�(�I��� ������RN�U$�����>̘p��mRUM����$r�R4G�-�_|���h��;�U���d�䍌�6�R=�����4��h}����_|��~$p���Hh��>��/�����~�)�����(�ɓg���k�c)�댼�׻*\����Iu ;F�F�,r�ڑ�F�{�U�w�����h��?s]�,�y21F����v�e�j�&���8�&����@?w	��0�!#Q�q���bK��,WU�}��:.8��K�J�8I�%&���=�)�uv�ݷ�|T�<ٺ���{r9-�I��RWj�;�Z��ՠ{�a��~
�DQ�Weآ���Ex�7��.e���]n����M��T�nL��kQ=��D�qŠw���]�@�t���ڴӇd�㍈�6�R=��h��:�V��jנU�:�9�DdlmE�{�S@��Z���@��Z����5R2H�4>DF�����w����}��n�C�+�%j��G��pm���e��N["f$���bK��bK}X��r���w{�����ʗ��@��Q�]f����X�K�Z�,�����N�p����	�C�/�_��-�����ڴwEV��<zI�
L"�8�޲�Wj�=�ZWj�9{��D�$��r)�uz���@�]�@��)����G����Q8�K�̆$�\�$��ŉ.;��IH�˒d��"(��Qh��h�e4]����I$�I!$rI  kY�d^��麱ĖtǬ��*�.�ays�n��Ǝ2v�ݵ΋��$�0�����ۮ�RSI���&������n����s��Z�F�㥊�u�aΖˢ��ڤ��uC zMX�ʝh��5��HLNܲ�0N�Q^�������z�).�����ܙ����z��jo@4��Ifːm�q�ܕ	ue�RڪI}'�/��ӊ�H����8�Mõ�K�cr���@n˞E�m4㮈���	b��bh�.�e4]���ڴw(�j6�d��hwW�{�*��j�?z�h����1F��8�wEV�|�Z�YM����p�\S	�1�V�bJz�1%��,IC�^$��ʴ����H��Ra�Š~���(wKė��IO\�$�������� 3�mڻ]�v�e4$��./m���Tq�2��hN_��}��5
���T�-���?~��I{��ė�8�%��,I)�y���D�w�������R�^�����*�!!*��ٓ� �0�}�zi�\�$N1F�ڋ@�v�����Wuz��o@�����(�6&
C@�����ֽ����z�����@YdQ�ۑ�F�r��@�>U��)�~���?[�T�^ҺgH�As�f�$�_H�Nv���;M�R*lK#�^W���닉5���o��~˾��Àw�0��R��c�����y�)��	�D��ץ4z�h�k�=ϫzz����$�R`GrC�w�0�}̾\�J����J�UQ-Yr
|R,X�̑(ȱ�J��$6p?0_�� �F�Db�&��Bc2"@�� ����8�@��AB�B,4��!HK )�!��Fc�8� ��V$�U��
��R���SO�؉�B��T�#����
�z��j� ���ZiU]��3_��36^��;ϙd��b�4���Ǥ�I{��x���$��ŉ%8D�H��q8�q��ʽץ4޳����IU%��C/U�\Wq�(��k	[��.�a_`
���09w7Gj�V

3i.���h�#/�m����w�o�ڴ^��]��Q�8���Hh��h�k�:�[�=zS@�ܠ,w$n6�di8�^��]���)�~�ՠ~�]�,�y1LQ�d�=���ץ4�ڴ?*�\������b��bqHIl��7�z�����V��ֽ������]��=��[��9��Z�7@&�Aqq�u����p\�,�!���v�*�Ɉ�9!�~�ՠr��@��o@��M���H�f)#Ocqh�k�:�[�=zS@�]�@/![	dNI�7���ށ�Қ��Z/Z����I�'�q7#zf.��Ɓ��-��zWkzTE��!Lq6&
C@�]�@�3+����{3rO��]��m��R!!�,V#�E�w;�k@` m�hWj�0ȍ�Nl�낞�C�t�C�ṅ�����!Z�y�I��cI�^�{inN�7��{��t�ǄW����?[6�ivb����A�5�ˉ����e'�6 �éNK&ݪyR��7��<Fɵ����۷U�6�s]�8.�n�4��(�vkq��N�\X�z�+�b��B���YV�FB6u8�,!nY�$�����*㈁���e�=]c80��vC6�������nwM������k(0�e-�n���H1h+~z]��ץ4yڴ�k���&)�4L�ǠU���=zS@���@��^�z�ˊa2BF��7&��Қ��Z/Z�
���g�^=$��
L7�v���z]��ץ4β�G�H����Z/Z�
����Jh�hكiV	��x�5&}�I�0�v�{�;�M�݌�0Z��-f���1V�t2H�Q����4^��=�j�9zנ�7rHBF�#n5�@��NE�Uj�U���8n�8�_�o�c��&�qKGB���M
C@���@��^�Ws�@��MԱ���N-Ľk�U���=����ܴ�j�*LSh�#�@��٠z����;V��ֽ��ʩ�ӂ�	�N�u<.۩\���O��ݹ����(7.9��F�I�������M�v���z]���ԯ69�
L7�v���Z]������Y\��b�4�7�}�}۹'o�gu�
�$H�тR��*>̘p�̜ �1�BG,��H��hw;4��h�l�;�U��7rL���q��Q94��hz٠w>�@��Y�Z�mQ��kcFc���.G�f��(z��+1������&�[�k�7ƕ��n�]��Ĕ8��%�8�%�"��5R2cNM��Z\�����޶h�w�2���1F��Z
tx��X�]�$����%�Q�⌐�����j}�� �n��_��>I��/*��+�c��˸e��Ȥ�R`	�hz٠w>�@��W�~�S@���rI�����J=&��tvۨ���a.�n&K�$L%�M�r�q]��$x��<m4��;�U�^k��?[)��f�\�*�H�"rH���S��x��X�]�$����%���&H��I$�Ɯz�e4�l�;�U�^k��*�GĢ26��ėz�1%�}IN���Kdq`j����dl�'�����?d�����y��4�TIR���N�~@ m� ^��]5��EC���&�:�:0nw^)L��M�U�����ґ�N�:n�gd��ݎ��o�;[��֧��$�8��)�[�]�!��1�1��.�izv�k��Ӹ��UR6�ù�����	Ϟ.5j�z@��GA�0uIh˄4�Z��l�m�WD����luq�͑7Vb{(6۰�&��X+�.��-�:��aG�ߝ��}��p��e�]Z�k�b9�ۮ��뷐�ܕ�˶J�v�ϵў���R��_�����%%�bK�r���1 �`��8��$�E%ܜ�ɇ?R�����@�ߖ�Ws��H�<z9�
Lԋ@�|�]�@��@�ڴ����$x��<m�š�cݛ��f��� ̼���I�f��V!/��G�E$j	�����]�@�/1���|�'�&ޥz�q�+��(֌)q�6�'M��n�B:5;���˜�%����m�5��V6��?�����e�>�y�R���׷�5������b�v�!�;����%T�5UU��fe�_ �_�_ �ɇ5*����c��26F��@����@��@��h�e4q�*LS#a ԏ���'�����8�ɇURI����:��;�qE!%�d�_ �ɇ ��I.�y��n�����.����C��ў��]sѢ�-gN�ogIŮ5�4ais��N��m�ss�����ݾ�o�(
L��;���ՠ{�V�l���}��BG�H���R��ͤ�&�e���ݚp�&ڪ�M���/���$�	����ށm���O�p h�L�����;~�� ���$$�(��E��}�������8��N����~J�*~ɛw�5�a�\�����ݗ!�;ܘpʪ���o��]����hw��<�C�n�W@؎�&�;k��&/v�����;Iuew�/~�����ls����-��}���{�V�l���YM�_��e�qK��%�������%I~I%Uv����X�����$��/Z.�EćQHIa#��3�0�w&6�$�+~zWW�@��+ǣ�I ��N\8T�$���^f� ��/��*t 0E�q�;�w]��}�静�Mk)$��܎C�c���ҪT����o�i�>�L8ރo�.&��D��u�e=&g�N�&�������9��-ш�<q�#PjG�{�*��)�}ܘj�J�a�3o��w�E$���#��_ ��ß�W�*�=���~{���w����f�l7K�q2]۲�8��N�����*T��^m� �lӀ}�8��,�9d�$�p�~IUU=�;�۾��qp?RJ���Ӏw�TGȓ26q��ս׮�����ܓ����� �?"� t�E#d��#e��X�#%2�'Ȝ���_�2)e�/� ����c)���A~%��B��dA��� �>���	7�V'�@�SJ� ;�zE�~���[
���	65�B:�R%@���V�_`Tci�H�  ��H�Q��p�$V1$R0"1$l� ��mZ���3��?�X�R$����{�/>��߽�����         �m�  m�        �h  -�cq�_=\�U���,Ҹ�l�$��X�1oT�u��N��۶P��V��ĄY혲�pn������Vں<�9x.��sm���)�v0#ړe�F&΅�*v�a�0���0�:��'�m���0�c��YS9����'c�(*���;S[+�
�����mu�m]ur�cvc0���!5Wc�H�YW�I|9^M���BYjB�L�N�"�X6m�s��L  	6�H�Y��t��;Oh�7���72���'Q���P�9�n�m2�qi��b�����[I9��gg�N8�Cqvz8r�-.ū��eƮ2�Kru�yeĘ��1���;)����r�`v;q�U畂��a��nC�-.�'����mڢ���66��9Z��Pp�]ll[M�J�m$�����=�V�MT��Ply��-�7 �9�*�ۂ������g�tY9��`�)f�yZ�m�m���j�U�\�\�hE1��Z�r@ �`�iem��u&�)VF�e�%Prni\kpz5
�fy��۝��d��ة���.�F�f�)�n�����ҩQ�b6z"͞�����eN#u�mRm٥=��#��a�(pFy@9��j8��b�<RZ�ŷ���t������`�X)W�y̺8�6��8�J��QO4�I�ء�u�p���W�J�7�ӹCHg��J�n6ɺ�Ε܌��ydI�;�9ն�еX�M�3�%����64lt����t���"ӛl�ga[fも�Z�7n*��O+���y�+����V�1��m�ӆ4X�m6�IԵmN0�qt���.�i��4�m�ԇv��*��KC����e�1�}�܆�l��
�m�Pl�<55
�<σ��ݸ�n
n˻L��8zKr���Q��+���2�Yu.*�HE��P�6T0Q�@#�� l�?�@־޵�kZւ�[@��l�z#Bԏ#���]<�Odr�����[��R֔�ӻ.��	��h@�5t�@�Fغ;#{[8�xxL:�s�[�k
���5�BT�F�k�G99c�bj�{av]�v���@K��v�ғ�p��AcV�۬��r8���=
�nn��cm7n���뺺�[��<3˻f��C햑�,)Y��k��<g����R���v�)%�EnYtm��[��P��+Y��2.���]{J�r�A;�8����2Iw�f��p�&Ϲ��UK��Ƿ�1n-�z9�
L93@��)�r��@�t�|���檪l�^+��$�I#����W}��=�+Z�]�޲�֍�n5$jH�>������h��.��Á����v���z����qȤ��׮��YM��z}���y�2��Z��r6����Ml��r�1� ݇�^�����D ���� �s���CNg���?Ɓ�ֽ�ҵ�z���?p��u����d��ܓ������G��!�qQ��]�K������ ��0��UT�g|e>D�)�4HǠ^?����sO�bV��U�|���1:
d�	L�w/��%I?noˀfdӀy�2��Ο?��s��E$�������4�����
����=z�h�	(�w�Vѝq�Ë1h�\^�1�^��=�
NN����M�k�Evhk�O�������<Ͻ��ӑ,K������DȖ%��{�iȖ%�b_D��,�%������7���{���{[ND�,K�w�6��bX�'{�p�r%�bX�Ͻ��r�bX�������`V�����Y��g�����ӑ,K��{�ND��Q*d�B�ݚ���Ͻ��r%�bX���=��"X�%���ۄ�L�j�Y�ff��"X�
@Ȟ���ND�,K�����r%�bX�Ͻ��ӑ,K�����"X�%�����{dV�%�"�"�/�L��L�����r%�bX�Ͻ��ӑ,K�����"X�%����6��bX�'�{s5��+u��:E��E�BgnǴ/d�⣷Y�QZ-�$���u$�/��J��3Y��Kı;�{=��"X�%����ND�,K��m9ı,N�o��)2�)2�l�������5�ֶ��bX�'��m9ı,N����Kı;�{ٴ�Kı/wvr��/Ԫ�+t���[����r9&�։%�h�r%�bX����m9ı,N���m9ı,K������bX�'��m9ı,Ow��њɭe�H��G!�_�I��K/۷�_�Jı/�{��r%�bX�{���K���H�t��w����ӑ.��oq���d��d�,����ou�bX����m9ı,O��p�r%�bX��w��Kı;�{ٴ�FRe&R��U~���]����d�\�.5�fF�{8�х{ �=�g������mX��x>m�`��w�{��Y������ND�,K���6��bX�'s�{6��bX�%��{[ND�,K��	�p��f�0��ND�,K���6���E2&D�=���ͧ"X�%�~����ӑ,K�����"YI��K�Dj�n+q��K�r��&%�bw>��iȖ%�b_�����KlK�w�6��bX�'{��m9��I���(���E�.�@�/��)X�%�{��ӑ,K�����"X�%���~�ND�,D����O�L��L��3�jqE!%�I.NQȖ%�b}���ӑ,K��{�M�"X�%����ͧ"X�%�{��ӑ,KĂߕF*$��ֵ�kZւ  m��S�M��94���v���W896��pF}�(�0B�;���]\��s�ȴ�M���L����S�L�v�*hH5�%���[D8�t�V�:��M{*�잜���Q�l��L7Bͭ�BL��Y�o5`�g�c<�I,p��m�"V��Ok^�oh��jĝ�9$�%��\\����q^��V�c�-���k,���z �P9�K.���wK���)6�,1"<�`��ٳq���ʵ��R`+��{Y�EV+��F��Kı?w��ӑ,K��}�fӑ,KĿ��ka���2%�e,���\��I��I��~��HId��&�fkW5��Kı;�{ٴ�?��L�b_������Kı;���ND�,K�ﹴ�ı,K�ze�d�ܷ$�r_)|Re&Re'�ݜ�Ȗ%�b}���ӑ,h�lN���n	"�{ٵ$D�~�3��fffL���AG�>�}�iȖ%�b}��ͧ"X�%����ͧ"X�%��}�fӑ,K��x��{&\5tY��33Fӑ,K���{�ND�,K ;�{ٴ�Kı>Ͻ��r%�bX�no˔�)2�)2�w9v�n�c�;��	Icaf��r+��K��D�$���\��"0�Kq[��e�w9K�)2�)e�}�ND�,K���ͧ"X�%�����U��&D�,N����ND�,S){���r�%��._)|Re&Qb}�{ٴ�*ı>�}�iȖ%�b}����Kı;�{ٴ�FRe&R������������%�b}���ӑ,K������Kı;�{ٴ�Kı>ϻ��r)��I��n'��\�I"r��_	bX6'ｿM�"X�%���}�ND�,K���ͧ"X�%�ｿM�%&Re&R�ͽ$�Kd�;��9R�Kı=��iȖ%�`��wٴ�Kı=����Kı?}��m9)2�)2�wx�����CW�v�����}�wW�=�����NwC�NxK�hyh;7]4���K�˖��nK��JL��L�����K�,K���ߦӑ,K������Kı=��iȖ%�b_{��5�F�.�.K�/�L��L���i�9�*�r&D�>����ӑ,K���{�6��bX�'��}�ND�*���_���h�e�Q��www!�_��%����6��bX�'���m9��^����Cg"j&��ͧ"X�%�����M�"X�%��f���ˣ.��d�.�6��bX�'���m9ı,O���6��bX�'���6��bX�!2'�����r%�bX���wg����@�/��)2�)2��ٷ�_D�,K�{~�ND�,K��ߦӑ,K��w�ͧ"X�%��}=`m��{N�Q�Wu���v��͓��J<�v�Xʷ�����u���ܦ�m9ı,O}��m9ı,O�{~�ND�,K���6��bX�'��v�K�)2�)b�Mm�9�D�jm9ı,O�{~�NC�@�DȖ'�{�ٴ�Kı;���m9ıK}�Ӕ�)~�V�YI������Kdֵs3F��6��bX�'�{�ٴ�Kı>ϻ��r%�bX�����r%��L��o4�/�L��L���[ے�r�%�[��K�)1S)z��|��I�X�'���6��bX�'ｿM�"X�� �jnD����3iȖ%��=���v�8�Z�e�}��Ou�����ߦӑ,K������Kı=��iȖ%�b}�wٴ�K�q�߿��)�� �`�g���.G�f��Ã�q�[б�7=�n���q"==��Ț�,�fff�6��bX�'ｿM�"X�%���}�ND�,K���ͧ"X�%�ｿM�"X�%��{v�{Yte՚̙�Z�ND�,K���6��bX�'��}�ND�,K�{~�ND�,K��ߦӑ?�dL�bw���_��+�K	\�R���L��Yy���Ȗ%�b{�o�iȖ?���>����ӑ,K���{�6��bX�'����jqE!%��|��I������ߦӑ,K������Kı=��iȖ%����ȝ�}��ND�)I��~����r9$�ˇ)|Re+������Kİ�������~�bX�'s��ͧ"X�%�ｿM�"YI��K?UUR(�J����I$�wd���`�Ӻ��\䜻�NvS<�v-;f�2��i����������"PR��t�m���홙CDp�6}M�a�jS=(2p���)���K5��7\l��:��#WeU��m���힝[mإ^0޺�K����ٸ֦\��\�#a�ͅ�7l"[�,���lٲ����,�׊{;��lW���q��ݏH})`��{��C��Y�f杫����Q��/l=�K��3Y��n*1MF�@�J)d�����r��I��I��^����bX�'��}�ND�,K�{~�ND�,K��ߦӑ,Kľ��/�d�*K%?{���oq���_����r±ș������ӑ,K������ND�,K���6��bX�%�˽R)$��$���_)|Re&Re/}��m9ı,O�{~�ND�,K���6��bX�'��}�ND�,K��w�p��f�0��ND�,K��ߦӑ,K��}�fӑ,K��>�iȖ%�X�{���KĲ���7Q$N�%�j܇)|Re&Rbw>��iȖ%�b}�wٴ�Kı>�}�iȖ%�b~����r%�bY��������`�]5V�,��r�������w<��f�c��]��n�c�x�^�w�]s�I�I��m9ı,O���6��bX�'��m9ı,O�{~��g�ı=���ͧ"X�%��u}�v�'RZ�;���)2�)2��7��� ��~@SH��,L�w��Kı?g{��r%�bX��}��_�I��K7[G$��MND�,K��~�ND�,K����ND�Vı/����r%�bX�{7��_�I��Kv<�r�-K�wr�u���Kı;�{ٴ�Kı/����r%�bX�{���K����9�)|Re&Re'�����%���z���Y��Kı/����r%�bX"1����O�,K�ｿ��Kı;�{ٴ�Kı/��x�u��\r�h����
m��{h�vJ���״�y�+[���{���q��F�1��Kı>�}�iȖ%�b}���iȖ%�bw>��iȖ%�b_�����Kı=�'p�ɗ]k3�Ѵ�Kı>�w��?��DȖ'���ٴ�Kı/����ӑ,K����.R���L��Y�A��"w3&u���Kı;�{ٴ�Kı/����r%���"����c#����D� ��`�jiI��$E�"��|�bA�\R�І���#2�&���0(��! �$���Z�!�\%$#0�c�"FH$�R",�#r*1� !D%@�
��x$ A�@� h�@J��"F`@#@��*6ჽ� N���H�RUXFL3��>آ�"��@O��Q�8|�E�D?��W�C����br'����ӑ,K���ߦӑL��L��G�W��|��E�`*%��{[ND�,K�w�6��bX�'���6��bX�'s�{7K�)2�)w�����BKRGrm9ı,O��p�r%�bX � ;�s�m?D�,K�����r%�e&R}���_�I��K��]��!��MY3:%��I�@uv�q$ۦc0�E�]������Y]9��-����=�{�K��~�ND�,K����ND�,K�ｭ�	Ȗ%�b}���ӑL��L��k�d���;W,�C��ı,N���m9ı,K������bX�'��m9ı,O���m9*��L��L��t6\�ww��佧"X�%��;�fӑ,K�����"X�%��{�M�"X�%�����R���L��Ow.�H��6I$�	s6��bX��'��m9ı,O���m9ı,N���m9İ4"uAv����3���iȖ%�b{<N�}�.j]5��fh�r%�bX�w���r%�bX�Ͻ��r%�bX����m9ı,O��p�r%�JL���������Ze�N\��թ�E����n����2]�';v��v"�	������G��I��v]�R�I��I�{;���ND�,K�w�ͧ"X�%����ND�,K��~�ND�,K�\f�(�������&Re&Q�;�fӑQ�,K�w�6��bX�'���6��bX�'s�{6��bX���G�'kS�)	-K����&Re'��m9ı,O���m9�ı;�{ٴ�Kı?g}��r%��L���[G.A�H�K�(��D����Kı=���ͧ"X�%��;�fӑ,KR�����
L��L��k�d���;W,�C��ı,N���m9ı,?�V?k��ٴ�ı,N�{��ӑ,K��3~\��I��I��U*K��ߤ�I$��b� ���֒ħYy���Yz�]��ܖ��kgy���RΉ�j�
��jjA��NB/qjsW)�`��dQ�݈��<��۝&�Ѱ�D�.�88�=��#��ٖ*˹�v�n����,���r��O[t��6�Q��;�������s�ZF�����\V0����5vܵǆxɪ'ӇT3�zry۬I�h'�T�"�6�U�D+w��͇j�������ݦ<K�:�<]x.�l<�nx�ww�[}3*��K?{���oq��'s��ٴ�Kı>�}�iȖ%�b}���ӑ,K��}�fӑ,K���^��$���r���&Re'��m9ı,O��p�r%�bX�Ͻ��r%�bX���}v���
�P\��,O��'���2�ѓY�ff��"X�%��}��iȖ%�bw>��iȖ?�ș����iȖ%�bw�|�K�)2�){H�uD�2]��捧"X� 	bw>��iȖ%�b~�]��r%�bX�{���Kĥ.�7��_�I��K�2��d��%���fӑ,K������KİQO��p�r%�bX�w���r%�bX�Ͻ��r%�bX�}�L��ftV����Un�u�i���=B����\��5��˫�E�w:��7����<X�%����ND�,K��~�ND�,K����ND�,K��޻NE2�)2���-���A�$�r��X�%��}�M�!J e ބ 2&D�;�{ٴ�Kı>�^��r%�bX�{���r%�bX�sE�Ԓ7j���9K�)2�)e�v�K�,K�����ӑ,EVı>�w��Kı>���Kı/}��r���$����K�)2�){&��9ı,O���m9ı,O���m9ıE����ND�,K��{�� �]�nG�_�I����^��r%�bX{��M��%�bg���ND�,K��޻ND�,��O3F^�ENH��%���ٷ�ɭ�_��w 7a�GT�ۦ�u� 4�����Yd�wrG�_�I��KټӔ�)1,K���6��bX�'�׽v��bX�'�׽v��bX�'ޚ$裸'q��w!�_�I��Ko3o��ı,O��z�9ı,O}�z�9ı,O���m9,K�������K��/��)2�)2��n�R�Kı=����K�!�2&w���r%�bX���ٴ�Kı>��'�RZ�Gq��&Rb��K�k޻ND�,K��~�ND�,K���6��bX�"w����ND�,K)?ߵ���wrH܎G�_�I��O���m9ı,Og{��r%�bX�w^��r%�bX��^��r%�bR��R�h6��k���#,��64�-��{u�6�Di�\\�t���O���5G��菉.Y%�$n�˅�r��L��L���^ӑ,K�����ӑ,K�����ӑ,K���ߦӑ,Kľ��l�r��In�|��I��I���u�9,K�����ӑ,K���ߦӑ,K��w�ͧ"���,K�����Ī65/����Y��g�������r%�bX�w���r%��%���}�ND�,K��޻ND�,KoQ���n�Y%�ܑ��&Re&Q�}�M�"X�%���}�ND�,K��޻ND�,/�V<C���(~ȟ�����r%�bX��h�~	"w��r��I��I��3~�r%�bX�w]��r%�bX��^��r%�bX����m9ı,O��m�O嫌]��BL�nѳ����,��]&�;:9/k���Ft�7�%$��W1���<X�%��u�]�"X�%���]�"X�%�w����b�ı?���K�)2�)f���?�)	-I#��ND�,K�k޻ND�,K�ｭ�"X�%�����r%�bX�w]��r$(X$��t����\&d���n	 ��}�lI�;���n	"z'��}v��bX�'�׽v��bX����uܲKRHݫ�q�9K�)2������r%�bX�w]��r%�bX��^��r%�b�w��ӑ,K�O}���˻�I%�NR���L�b}�{�iȖ%�b{�{�iȖ%�b_��kiȖ%�b{��6��bX�{������w��߿���  �UT�۷e@��&�����y^�8ᢵѱϮ��]���pt�Qq8�$��a*�U�9�ƍ���f6a���u����h
�c���Y�<s�RӔ�On.w]��n���9���n.!T�|�k�뎢tɖ�����tK���6��B��A3ǋW,�u���bl�n/ �d��5u��$�fːmq��۲�ؕ��B��t�M%\�dmvu�@9�=���H�US.n��x�f�~������ic�Iw!._)x��L��[�u��+ı/~����Kı=��iȖ%�b}��iȖ%�b{<N�}��,�K��#�/�L��L��۳��(�,K���6��bX�'���6��bX�'�׽v��%�bX����.��;��Էrr��&Re&R����.D�,K��}�ND��Q �Dȟ�����r%�bX�����ӑ,K�{��@�����r�K�)3�IEPȝ���iȖ%�bw_��iȖ%�b_�����Kı=��iȔ��L��5��A����Gw/��)X�%���]�"X�%�~���ӑ,K��w�ͧ"X�%��}�fӑ�7������1�?���܃u,/]E�=rF]��S��kZ�YUn�tҹ
�����Q���۸�#r9)|Re&Re'��m9ı,Og{��r%�bX�g��m9ı,O}�z�9ı,Ov??Fu=T2�_{���oq���~�{��r��"X������Kı=����Kı/�{��r%��L����{r��E-��/��)2��b}�{ٴ�Kı=����K�"^���[ND�,K�=���r%)2�)>�^�HK�8�rK�/�V%��� "w��iȖ%�b^���[ND�,K���6��bX�'����/�L��L����Ol�pq\wl�֦ӑ,KĿ}�kiȖ%�a�1k��ٴ�ı,N���iȖ%�b}���iȖ%�b}��3/��jˌ� a�z0�,��|.����)��[h��"�,��:BA�*����w�{��bX�Ͻ��r%�bX�g��m9ı,O���m9ı,K������b�I���(�����"\�R���,K���ͧ"6%�b}���iȖ%�b_�����Kı;�{ٴ�K)2�){b|�qE!%�����/�N%�b}���iȖ%�b_�����K+�,"�
P�! P��äD�BACh&��E��D�5���iȖ%��[~���_�I��I��ڎGn�5�[5���r%�bX�}�z�9ı,N���m9ı,O��{6��bX�R��4�/�L��L��k�q�RH\3Y��j�9ı,N���m9ı,?�"�u����~�bX�'����Kı>�^��r%�bX���L�ytV�u&'T��B;wW�쯔Ps��
�rg[sC�AٺuG��+�n��O���Kı>Ͻ��r%�bX�{���r%�bX�}�z��Kı;�{ٺ_�I��I�^�{	%���D9/iȖ%�b}���iȖ%�b}����Kı;�{ٴ�Kı>Ͻ��/�L��L����Ol�a"	.�ܓiȖ%�b}����Kı;�{ٴ�Kı>Ͻ��r%�bX�nsNR���L��^� �	"�#�yu�]�"X�%�{����"X�%��}�fӑ,K���ߦӑ,K���8:AM��]�"X�%������"�%��.NR���L��>Ͻ��r%�bX�{���r%�bX�}�z�9ı,K߽�m9ı,{���o�c��BjԨQ![ukp�n�ѝ)юڤI�!K�oh)-�����\�kXf�s5�ND�,K�w~�ND�,K��]�"X�%�{�����"X�%��}�fӑ,KĽ��|j�V��I��R���L��^��|��Jı,K߽�m9ı,O��{6��bX�'���6���bX�'���\��-K��W.G�_�I��I�g(�Kı>���Kı>�w��Kı?w^��r%�bX�ݓ���[�]f����Z�ӑ,K?�D����Kı;���M�"X�%�����ӑ,KD�/~����KǍ�?�����V*Z�c�w�{��2X�{���r%�bX���z�9ı,K߽�m9ı,O����9ı,M�	$F�KG��O��a0"т���৘�M�����!�KJ���9�*
D�
]0P��Q,��6���$�$-�(��k�a
J��$ �hV�D�r�$W@|.�� @�H�`'�,��ր         ��m�  m         ��  ���f�W[�l�t��&�<S;v�`�Uarw:n���ZQ%�g�b�mm����W]�3Ԝ]���Nֳ����ղ]^��\�\�k��)�lHD�-�rʉӪϳer�uz�v$���I u�M��5��iv�\qha��I+d&�}Q<�g���s���,[g��j�x�M���j��e�q�n6'\vӯ'[�u�ru�==Ӷ 5@r���E���Wgm�7�nl  �n6�7d.P[�_/��1���V�l�D��eL�;GU����eF�Þ6�d��$۳�v�$����<�uv�ui) �y�������n�6D&�&�2s�-��X��mUAԱ:�ʆ$��!��j9�4Pu�k'k��Y)��t���ޑ��J�&l�&�-�me�t���i՝2,7v�&�R�m�^� 
�
��[U@����n����dwe��[���ə+��@<��[�Di�Hi�Rn	g���3�*@j���S#��k���{�H+!5 !���m���zy5[*�I��a����M��Μm�[��+aC:�I�y3Q���&�*�$���0W6Qa���h�e��(q)n9���6\̹x��#`j�VV�W����-�U}�&�M��C�6V��F��wvBN-���*eq!	 ���z��`�+��gi��n����r���N��5@&ɺg�˕���-ѹ%;6�k*���WlӞ�[��\�$S$�	�t�좑��gV�!�Ͷ ���:�ѵ*�f�IP�M���s���X��̲�\����^iMZA�ꎺ㍯h8Bs�ȯ<�jIUl���t��ᥗH ]�h���]�`��Laa���b�ԫN��U��7b��d��&<N[��ֹ0�v�Neٛ]l������Ş��`s���m��M%�g� ~J���LQ>�h P*<D hAO��D�U	ݠU08ww~������}�� 0 *��1u#خ�Si:[s�ݸ^�z�4gΪf�vһ���Γ^�);E���Hf3t���ҧm�Yċn\\'56���7mb.koW���q�c�,���3c��݊��������Et�w]���E��uf�t�N��n�k6s��r��\cp��m&��Az���L���a�{>��<��GX6rg��j�������Q�:�]�K��1F�c�&��f���̄7=��$�Xң��ԉF��]�K�����L��^ٚ�K�)X�%������bX�'��}v��P�"X�'����Kı>�"�In]�ڻrG�_�I��I��{[ND�,K�뾻ND�,K�w~�ND�,K�u�]�"(�b�K�2��ND\��8��/�L��,O����9ı,O���m9ı,O�׽v��bX�%������bX�R����8��9i�.G�_�I�b}���iȖ%�b~���Kı/~����K�lO����9��I��x����I��R��bX�'��޻ND�,K�ｭ�"X�%��u�]�"X�%��{�M�"2�)2�^�vި�qE*Z.q^��tv��m��]ƺݵ��n�jgL��#l?w{��F������T}��oq����~ｭ�"X�%��u�]�"X�%��{�M��O�2%�b}�]�"X�{��?���D�!�B*�����{�K��޻NC�������6���%���ɴ�Kı=�z�9ı,K������ؖ%�z��L�e�rK��)|Re&Re/fsNR���X�'�׽v��bX�%��{[ND�,K��޻ND�,K��{Yr�2+$���R���L��^ɺ�K╉bX��}�m9ı,O��z�9ıK��~�ND�,K�MwBI-˸ݧnH�K�)2�)>���r%�bX�w^��r%�bX�w���r%�bX�w^��r%�bX��u����;��44�ŝ�^2�����s׺�[�n��܈�����RI'�W��E�]��j浴�ı,N�_��iȖ%�b}���iȖ%�b}�{�iȖ%�JO��9K�)2�){b嚜QI��Z���r%�bX�w���r%�bX�w^��r%�bX��}�m9ı,O��z�9ı/}�Oa���r"H�%Ô�)2�)2��n�R���V%�w��ӑ,}��$��R$FHl0P���"r'}��v��bX�'��~�ND�,K�=۞�]Z�AڹqG�_�I��K����/��,K��޻ND�,K��ߦӑ,K�D!�;��]�"X�%������W�`���������oq��޻ND�,K��ߦӑ,K�����ӑ,K��>�iȖ%�w���x����륪θ�)�n��T�4e&ݩ�z"��ڣ.���w{� �����rK��)|Re&R}��N���:��ʩR_0�^��x���v�$A#p��@�;V���@�;V���a��$��-hI����$|����K�r��G$��!�-����=��Z�YM��Z
�#ު�Ung6���)f�RG-)#qh�e4s�h^��+�������ػuo$B�@��M�1�]�[K�]��6�!���'LK�s����X��\�$�{��K���ﾭ�}>4��?�Q�	�a$Z��/��g��� �i�=��|�_����߾m��r72$(��*�}�z�YM?%J��^��~; }�⼅ۗd�%ȉr��}�Ӏg�u���/���*J�~���1��W��D]�K� �o1��R���6��so�}ܘp
�R
H
�0Z"�b��	�%���?���  m�l��iT�g� v�a.���m�v�s�5g.�sg��:�T�������d���C��؍���Ƨ�+���M�W������y1p�^۶�.�[��bm���v��;���nL���g�66#�Z�s�7���7N�]k��H��5Ʀ٭��VY�3�b	��s�͑�9lݤh��2��qOBg-��ǲK����{�Kc6x�<LS��]������-�Yx�q�ope';v�0�j�t�aŮڶ�etEv䏠u���מ�����*K���-���&}��r�C��W��=]�@�;V�˭z��qL�$Q�'���Zyڴ�333����9}~z�ì�71I���{�����Nמ��jJ�'����|����P�D�H�Š�f��3������|h�j��T1��t�\�p���٥t�Sj��G����vx��.�l<�n8V�+6&�����~��c���?Ԓ�_0=�����^��˲\��D�|ݼ��$�%UK�I�T����| ���מ��y�W���K�����c��̜?*�Y�r�����x��8�"�ڒ- ��4+���j�;�ՠw��"��Er`�˓�u�����̽>�~����f��Z6�G��x�hH,�"�i��V��z��8/k:��Ԃk��˫�t{X��
�Ks}$��?��@�;V�~�f��z� �0��q9#qG#���>~��/ԕRWa���4
����ް�@��'\Jȓ�."\| �{' ��e�*I~���$�Ȟj�s���r�I��w$��}2��\��-��Ԓ��{�|=��h�j�^�@?T�;�l��&G�w�*�;�ՠ�f��z�6ߟ��g��F��lq1	'o�ɬ�>���<��'k5c��o�{������M���$�����- ��4+���
����$q��#RE��d��j��+��u�3�|���J�T��c(���]�W.Nן��z­��Z��h�/�E�2d��r7r��_�*�W���������$�߻��� ?E �@��"I�QR�y̾ g@�A���NH�R2-��Z��hW��;�h�IW�����XEv��v�]�E�'x�:C�z�Z5FWg]9��}|| ��Q�=���|g���r$�I8������@�^�ް�@�;V�{�4Ӯ	�G2D��hW��;�h�j�^�~����l;��{eۗc�\�K�톾�v� ��4+�����H���Hܒ2-��Z��hW���2�S�o|4��%�-ے˷$| ��4+���
��h�=k� -�� m��]�D�m�܌Vv��غ�Y�.��G��֝��,b�v_F�t�Ga㍣(Rܯqk���u��f��\dˮŸn��v*����)�o����M�ڷ]�<�.�bi����
ȉ� ��d��%�쳥�n�2�V	q�7�����s��cq�.ѹ��u�ON[�43�lG(q�W8�%Cf�]�WB-]���w~s6P��t��$�^F�T��{[x��<�����.��Fn4"^GLa���\=sYv˓�c����C �o1�T����6pb�Tf�RZ�%���C��v� ��4+����
E���%��v� ;�����%T��?�����~|�;�#��7jI8�׬�<�W�w�*�;�ՠ�v�.�⑸��=��?U*K�UU[���>���> w=��}�v�s�܌RJ\�zk���� ;�f.^���P�!��G;Ur%ݚm[J0�7�O�ʴ�h�Y�y^�@�W�K�ܫ�ܑ� �o1�R�RuHJ<DG?
�͈��O(�}'���`y�m�v�c��TٚZВܗe�ԑh}~�����V��v��c(���]�W.N䪩��>z��|��h�Y�{���"�2BG�rh�r���Z��h�Y�{�B��Px))�4�Y-$�n-t�=�Z���qc�\H���);!@�~���ȅ�A���NH�Q��g�u���4׬�;��ZG�:�G �I G�z����h�r���\�I&���ݻ�Qۄ��29' =��nI���۹O���*~c���~��`���@.$00���B$P�)�0B�05U��1�vB0	��"VT%��IP�"-�L�o6�:Wx�XF��n EGDa��EhB��)(��hʑh�3И$��4 @*�+�1{��<�"��*����U� p6" ' 8���M )�:(���>�ܒ}��[�N^N�mF�$rd�M��U�w����d�m%M�sg ǯ�$�m�d��ȴ�h�Y��f��x��ԫ=0�z;�1���w���m��bx|&^�jwC���wBI�m��]��!#N6G!"�/���h�Y�w�X��J��]�ܿߟ ���"���d��X�@=z���U�w��@=z�ݕ�ɒ<x�@�;�h��>M����nl�u�#�q9#qG|ʩR���������p1*��*��c��o���-K�v��K���d���6|z�k��j�?[Ҹ��%lJd��f���۷us����S<���VS�:�kAٺi�͑Ț�sDRO���h�r���Z��h��ܑ�q�I��M��U���w���f�ʮd�5��)�h�j�^�@=z���U�ue�#N6G!	$Z��h���;��Z�v��bD�wr���' ;�d�J�U����r�_ ;���2�*�UE.�������www���  UT�WEt�W�.�Ѱ��ѱ����\��.1u��Ah�w1Cգl\�)�Z�`z$���N�b���C��(�瞀Jm��\��5ܒE�ɤ�g55X��V�!�����49q�m��a��R���mր�'3`�ֱr��w��F��!ly��M6U��*՝Iv]sv�`�F=��^V3Ϋ{g���y�l`,q���zT�3/���T���Y)8[���ZUR�7^�nm�ӻ\v� �M�-�h9�c��Q�8���ի�'��^�|�;V�z����4��"��RD�E2-�;V�z����4�V�|���$y�y$�qh�Y��@�;�h�ڴ�e�n<�(G1̎I��@�;�h�ڴ׬���ܑ�py��I&��w*�?s�h�Y��@�>_�:�q:N�%�\�2ۡ����f�z�z`�g\ܒg,H��ΦB�CQth�ڴ׬�wY�w�ʴ��[�vK���> w=��RT��QJ�TT���p�x���y��w��%�Ԃ`��&�{����U��Ro�{�����;�Q��QHH��M��U�~�j�^�@=�f�_a�`�Q��H�ȦE�~�j�^�@��zyܫ@���VLj:�óv�✗�f�av�3�L6�lƙ˗L��Z����we�I?y��/�{���UK������awr�q�\W�' �����IRM�����>�z����;�1�K��D���x����>��$��-UI.p��8�n� �����.[qY#rE2-�h�Y�Uֽ��U�{��$i���!$�@=z��ٗ�=�ŏ�w/1���U�4L�ێ���5M�$ۛn2������瞽��5�g�Wd�[�cQwb�l��5�
��=��U�z�V�z���*?�.)�$$x��zyܫ@�v� ��4]k��3��71I�ȴWj�^�@�ֽ��U�uiru�<�A<�d�-���@���ܓ��ӷrHD� A(�m�;�@?{��yY#�&G$�*�o�j���zj�������N w�����v��B'\����m��S��E���iz"6z�ka�ܱ8Z�7S�Ɋ��H��V�yڴ׬�*�^�ʮd�4�2F�dZ��h�Y�r�^��w*�=��$i��r'$| �{' ��e��ISy�կ�{���@�5s���0N94]k�;��Z��h�Y�{���"�����%�v�c�Խ�u��͜�ٗ�?*)n��$�I$$�$�wuUR�\��
�7H`�h�M]6��rY+�[��g�v��̛ ���ɒy(���9�����	��q�n���Y��i��e��OmݚEb��mY�=�0��fEnh:{*����m!u�+��jt��!u�n��;-�5=���%�(�����7D�s���7/<Z��/<�Z-�g<Q�ٶ��p/F�Y/�wc��q��\ֵD��#�����u�Kv��d�tXs��n�mhu��:$ݢCl�y���M�8�X�s�bT5u�\��'����bIztx�㤼Iw�T1%�È����"���s�9�J��n� ��ϖ���Z{�q�H��#�@�ֽ��U�z�V�z����w$cj6)#s	#�;��Z�����N��I����z�K�s6�dZ��h�Y�r�^��w*��tx��d�L��'װ�q�n^8e[ܘH�m����>���umCdj9	1I�z��.���r�UUI|��{��{-�C�v���w�.��b;��Z��h�Y�{���"�$$x��zyܫ@����UU$�=���c���u�	-���8��R�~ٺ��͜�ֽ��U�uk����r	�$qh�Y�r�^��w*�=]�@=��~��R/\�,=�8wJk�qn�W��[�6p�����̭�_�{�܏�Y��v�0p�����M��U�w���~@z� ?^V1���I$�=��@;��π{2p��ڥM���{d�q��n�|={���d��T�*Dh@N.d��w[�s��*�:�e� ��BLRE��f�w=��{��j�y���ޤ=�8���M ��4�V��v� ��4zѵ��y �S$"�CaE��E�g6��˱%�0g\ݢ�Mqu����y1I��o8��;��Zyڴ׬�^�@/�ΰPq��)�E �o1�j�&�ۛ8�͜ݼX��+���'�L�Š�f�z��yܫ@�;V�^����7	.N�������g�V���c�~L�]�U�UT�e͜ ��RYv�b�7$�yܫ@�;V�z����h�!�8'1�HHr�����Y}�	*��v.�'k5c�E9�L��ے)�h�j�^�@=z��UT�a��Z�m�n����BD�@=z� ��4�V��v�����8�L�M ��4�_IU&�׺��͜�X�"��D�o8��;��Zyڴ׬�^�@/�ΰPq��)�L�@�����p��N��,|��I"�%�E!JA����,$��1B��
ʐ���V�	D�FBL��BĉR��ʩ*����"P��HR$$VP���*J�� ��b"X5C4a-Ib�f��U7�F�����sf�) %��	  �08���
aBkn��dX��BP!FT ��r��m��5F$K`/�	T��f�f��      �� �m��  ��        	 [@ m:�Փ^ۮҕ��P��Q{m0�L"B����l��l�A��]	Z.�x��ƀy^<��[r����n6[pW]��ό���鲜�� �������9��7 ��\�m����*�% ���eʘ�l����vu3ҥ�8vt�'2�μ���s�l7IP]sn�vc��w��䳺���v�4�M��rd��j�@V0�(7fC�T%�KrJ��  i:�nӦ́�j�wi8�fK���4f�x(��Su��Z��U���I9�`���x��[=FteJ:�^�m�&�u��Ͷ�֙[W*�t��c��4�M-4�j�ʏe��*nm�j�.+Eh	{8e��Wgj:�t��]Y���c��BU������橊^�i�kkkn��b�fj�q��ϲx�̍Fd�%�R�TY�
�kj�*���<��ی]�KwJe]�l��^� \�$O\$:�JI'���[F��j� kY�{m�bIm�7UTjP�����̆�6k��X�nF�d��\�7gf��J ����+�	��0�����Kd�nRZ�:]nv8��v���{�n�l �����.��#��X���M�In�����5���W��8!�-������4�K�������6��b�74���S&+��HդN?|m}���m>ɮ�t�vFت��&�bxz��V��@\m���Ni��'�]�{5m�z6���=(��2bg�+���ܻ��VU����nҋ����Rl.�Y��"�\�i���M\��1��mmA5�j[���5rX�É4=�ڴ�,j[��5�@ �'W]	6��6�i�N ��y_����6ڮ^vӜt�RNprtu��8m�rlԂF�*n3�6�-��G`��`�Y���֤�t](�< :Aq@6@z�&��"b�p~t~ �U�(S�}�ٰ m �zJ���GXw&�Gp��V�E���ecld�p+�Nq�h�EvtΒl�$�1�`�c�m���s�5��4�l�W@W�Ck�c��mm�5�n�lg�&5,�sv����-�.�@U,�d���\�7sg=�{E%�עB3lث��F#qm�90`�/1���ٸ��1�j7F.^�F�mP3�l4�ਙ���]��rK�a�!�}��ﻼ?l���غ2�cj�Հ�����vu�L
�!ug���}�@H�������~>鵖�y$�G _����@�;�h�ڴ�X8�`Ԙ(�rh��s�*�I�=z���� w=���~����ۮ�),�r�r��.I8��_� �ט�~T��M����fl�y뼲G1����2)�h�ڴ׬�{�8��y�_ ʹ�Аv�q�H�#�s�8�I?fl�����>��Z�`ڲ'$ȔdDI@��na5�N�{]���N����&�Xї^GLa���l=Q&	�&�{����U�~�j�^�@�ʏ�PR��8��;Ν��A����#�N�?�w$������{'?*UJ�7�Y�.Y,�q�������h�Y��@�;�h���.��v����mW꫼��� /����w*�?s�h�pq8��0QH��wY�w�ʴ��Z��h��J��s"q�d�&�
���) w;g=;�ء��B0r�st�ֺ����lQ���@�;�h�ڴ׬�3���h}[��9�LDmɑL�@��ՠ�� �u��V���-	�E���- ��h����0V~H�*$������Λ��;V���J�yDL�M��$�+���8����z� 3���;����ɒ<x�@�w*�?s�h�@=�f����21<�ҝH�խE��;m�)�����:�i_K"�YL�
��4.s�����.7qG���| ��h���/�ʴ
�r� ܃�$�� 3����R�l=���o�W�@��ՠ�������D�@=�f�|�U��1/W��@>�����I�.�.]�䓁��US�MZ���w$����rE����FL�vh���$s��ۓ"�����@�UOs6|�͜;x��v�]�n���N��l2Ͳ!3K��2�"Ż��;Z��m�륓j,�3�$%�Ոu��Y��f�|�U�w��@�5s��K����8��N~UI&�����;�����N~T��Z�&��)	-Z�rp����>��>�T��s6p��h�3��L�qĦE2-�;V�^�4��h��Z^\\�F���$D����N���fπ�^�|�^c�J����d�d�I$�H0�`Z��'m�/I{E�v۩�x^�{c�C�g��Cc�<ut�%��7b?�Wb~|��J�Bz�u�8/K��	!�0���5	�X���݂��\�ml\��+�cmp�=s��]laC�W+�����7\`i�^�=�Þ��;]��3[Tq�����Ĉ��ɞ^6{�Rt��tf��Lt��fnI���۶�͗iԏ�6٩��՗T�~AB�	Qv�f[�;=V�H狫���{}��xջ�r�z4�����V3C�A�5����f�+���IO���Jz�C[�!�%;�Ē�	N���q��$��V���W��@>���@��qG2)���"�����@/u���4�r���Z	�j9	$Z+k�wd��ŏ���&����&��q�0�����:��h�ڴV�����o����!3rN2�7]j|mэ���1�]M�ѹ!Ψ�`�S��b�$x�rh]ʴ�h��@=z��뢃��qĦE2-��|��URT%J�+f�߿_ 3����x��
�����O$�#�@�mz��h]ʴ�h�pqI#	28'#��.��4��>ZyڴVנ�W�q�8�q�I4��ZyڴVנ�f���ڿ�&I�%��K�r�F�̯�ϓxo[�bSREg��L��
���.4�t]m������y�e��쟿Wl7��_� �֙��I�j9	1I����׬�:��h�j�=ù�e��8��H��~����w:v�qCp� P�P�ӊ&� �����{�rN߾�nI�����)	-]˓���͚�����@�mz��h�g]dc�%2)�h�j�9[^�z��Wr�������?)']xsvl��أmBuv�n}1iJ[fͦ3uY�3�������Z	�q~ �}��^�@��U�w��@/u���II�Ĝ�@=z���V��v� �l��+����q��$�Wr���Z}�ﾚ�_��˫u�8�1��&G2-ݼ��fd�s�8�UT$�
�$`
�@M}�t�ܓ��D�F����h[f�˭z��c���|�J��f��
]Zl�Z��M�v�TxW�.�ށg8���;a��O�8�|p�a-�䓠k�߯�uw*�=]�@:�4v5sA8���]ʴWj��f�˭z\3��L�qĦE2-�ڴ�٧��U~����>Z*�� ܂y#�G�w[4]k�=]ʴWj��`��G��$JI4K���%�r��/K�Ē��K�����,��"����τ{�o�� A� ��������n�zƛg���e�Sv9���.�\��G\�G%�i!����VRρ�=����K�q�u�7m������AZ �6:�X��j����d�kq�8�Ld��0˹ݢ�ɵ��ζJ|�n����-���
�[=��ư��S,Li����G��:�t��귳�/���w��}G	�).a��-�P��P���$���<���"uɭQq�b�w3ȡ�-Ʃ���v/�.���B���e�$����g�Zyڴ�٠�f����Ԏ1LdmɑL�@�;V��H37g =���w/>~��lʹ��A�@��- �呂z����V��v�������Ӓhs�8r�c���>�I$�n���{eAڊB]��rpe���?RJ������呂z�����Ҳ(ō��*�H��'ktug��v�.��R�Y��p�q\��:Y�&�hf�W/�I������� �>�Zs��#��]�$� =�����QT�**���$�r�*J@�{' �׋ �o1�j�*M���-�-�%�Z�7rN {sf��ܫ@�;V�u�h�+���q��$�Wr���Z�٠�f�˫u�8�1���dZv� ԕ%O7v|�͜�x��?����g�.b�<a��FC�+Ix��+�ݞ;D�;qQ�۝&m&��U�H���@=z���V��v�������Ԓh�Y�uuc���> {3'6�*T��W�P����7����-��Zs}��$Ua�I��B� @�3���Ԉ-UH�:�"EZ�X����[�ϡ`%BX!P���IB !BE�`P�0%�B���Э�]��J�4����R: ��HQB\��ΨְNP�;�9��(@
1H�*D ���Gb:H	��ĺف�gD�i�\�W���$�"`0`@�U��(�A� 
�DƂ0"�N DX�0!FD�"����	"A�	3�j��Dj;B�Q�~�?Oʣ�`�P��@� �@� �@�&�؊=X	E�!����h�Y�z�������8�Ȣ���U$��M������pe�@���Aȑ$#�#�@:�4Ԓ�~�����_ �o1�������ے�\0:���)G�'s��p����K��nz�Б$S�z��h�Y�_;�h�j�g���4��1�q��$��V��v� g����d��ISf��{d��8���S"�/?�Z{��^�@�w*�:�ZEj,$�pjE��� w=��go>�䐕R
��J���"�򠟃����w$���n��ݎK���d��R��կ�/?�Z{��=�"��Hb#$� ��x1�9gYռ�u�F�V��R��B\�3�Pɒ�n94�r���Z{��^�@�a������9n(⏀{�����6������3��?UU*M��c�\��!"��%Ǡ[��^�@�w*�;�ՠ^�SQF���O$i�&�z���V���c�m*I~�W�N {��+�eۗb�7��@�w*�=]�@/u���??7�O���{���~@ �ª�ju��3X�3���8կ\������v��v���ts,����6�Qu�7]�f<5�`��|t�@ ��k�2�lWh�$� �u*�b�Z�t��s׳��Ln����L՞}X����)�L΀��j���u��ۚ�W!a&�e<Bj�.�I*�ųlW
fpVh���A���^�-��G��������;��w���͖���\Mdb���]d!�8K���]wdAz&�+r�5�4�N(�E�_����^�4]k�/�ʴp�I��H91��_{'?��f<ݾ��Z�r� ��B���L��H��9u�@�w*�=]�@/u��g�'�$#x7#�/�ʴWj��f�ي���@��>�����8�ȦE�z�V�^��%�Ix���PĖ�$��O�n���.,���`s��r��l�鰦:t�?��[�@؍nRb�!�F_Ԓ??����נ_;�h�ՠ^�S�D����\�k[�}~�s|G�tDpDv�UJ�IWꯡ�z����_ 3����Wcj6(�q�H��r��ڴ�Y�r�^�U�뉷1Ldm8�����Z{��9u�@�w*�=�ΤPN$� �ƤZ{��>���?�}���h�ՠ{���d ���[B�6��y8��1�v�M��֎zP�Д��k �]ظ��.i���ӭz�V���Z{��=����d�o�z�V���Z��h�׿$}�S��#�L�d[�}�����~�4.mUt����ֽ�>ʴ\�ND���$p�- ��4׬�;��Z��4��q��R<��H��<���^�g���ƀz���`�T���l�5mY�l��Mkw#��t:�/V�2��f�K����R\L�����������?z�h�Y�y{��9^N���SN(�E�~���^�@��W�w�ʷ�䎣���D�r!�h}~������U�~���=�\�\�����<����r����ܟ
%@b@� q�i*��gg �U�$<j)	v��/�{�� ��_�{?}��~�Ӏu��|���q��.�=��.g0ui��j燶�Wa���얌�U�KKVS��6K�QƦE2-����z�������U�r�jpr%��#QHh�Y�y{��;��Z�YM��#��ڜR<��H��9u���r�?ٟؗ�����hUP�Q�G�JG�w�ʴ޲���h}�����|Q��nA<dm1ɑh�e4�-���~;��X��J�)X�$��[@�޷�F�4.��ҪԀ��3]gqF1#��LY[���NPu®W.Ѳ�!,����^x��چ���nu/C�G4ײq�񙱺ˁ���uu:$�\u���Eu��#���e9Z���\IrȽ�v���md�[Wn�x��_cd�Ѷ�n;Y�G��/7]�G%�e��O-��i���k<�vJ��ɨfCJe����j��C��"b�������4a�����e-r&"hp�p9跬Wknm4��Œ�[ѺX�)rLI��p���8_}��3���*��}�N췩P�E"r�r\���^�|�U�~����f����v5s��E!.�w%�����>�L8~�X���M�_���8�R��#$q��L�@��)�����^�|�U�r�jpr%��#QHh�@�g�s�����ϖ���S@�lJ�i)-��@]ϛ|�^��Z���5ړpIYM����Pn����2d�n]ƹ�ԓ����3�� ��0��K��l�k�^��˱˗r����X�Ԓ_	RDP�`E�$��Q`UD*�%T�8w�0�s2p��/�UNq� �26��ȴ޲���N�S~~;��Z�|Z���$���@/u�����ܫ@��)�{���ˉ��1F�#�@��W�_;�h�e4�Y�yx�U���'#u�b̭�mj|mэ�!x��Y��W��r6�Θn0~��}�wc퇮�/e����ϖ���S@/u�����(ޥ1���8ԊdZ�YM ��h^���r��+S��(�$��C��d�}�_R�K��HT�'����P��0P�s���Z��?Ɓ�׭D�rF�F�rbKǺ^$��T1%��,K�����$�����أ��%#�/�ʴ޲�{��<���φ�ɑD�<e��J�a2�ۙ[�����J�郪�b�\������Y�����G5����ߧƀ^�4/uz�V��u"�<�� �Cp��f����9u��s�>Z�YM���\R`�(��rp��/�go>�S}��8��8?>{%�F�.����nO /���s������p=�_�RKԩR�T�5m�^����oR��#$q�ȴ�qbIN��%��/S�*���v��.|9�6Tbأd�um���f�ʰ�a����l�@��ALWRE �{' ���v�c�U��RU�g���������4��8��<����6o�V��lӀ�d椪�l3~i?�ڍ�8�bR=�g�@��)�����^�U8uƜ��"6�r(���T�}�Ӏ���u��|ʓ��^��-f�ȝ�R�w w=��=^�;��o\�zx��$��W��EW�� QU�� QU�����
*�� (��� (��ʊ��� *( �B���� `* `*�Q�V�
�R"� �H
��
�����"
���H��",H
�X���`* *Tb*P",TB�V"�P��A *`�� b*A��DF�R�(��P��D"��UX
�V��"�V���D`����@��E`����@
�P�"�`*(�
�Q",Ab*Q �� *b��
�P�"���`����@�"���@�"�"��@� `��X
�R(�Q�"� * "��T�"�
���T@S� ����_� U| (��EW� ��������
*�� (��� ��� ��� U 
*��1AY&SY�����Y�pP��3'� amσA�f��  4   � �  m� @�. T�(@B��(U
� �P �� P 
  ($  ) UJ�P%E(��� '   �P  �g` }�����������׷����}�(Uw��so��y���l�v��������
=�m��Zy����^� }���G�ye�u�N�[�J|��{�mO'�]�7zܯ���W  o�$  P D�jU>���g;m�y���e}8���@���g���t1v�`�R��=��`05�ϫ��T���^N�^�sﳼYr�{:W���m��ޏk�ܚ�8��7���Q@�  �@F@ >��������x�ի���������ju��U��V�ܪ�]Ǖ��^�Ƿ^ W�T��z� ���8�r����]��^�w�W��� s��wR�����v�j^��{�׀��PP  
PP(H� g>���{{�)�w��뷝��6
 ����3e M )�� �΀)΀  �;�� )L�: M((� '@(� 4�`t�w0t�A`��(�� �gJ(;�t��� � @ �@�w q(Ҕ��P  l��[� }7�O���j���sw�+�Ϸ^������ɷ�o7��x  	��W���*�@7��s>���y�ǻ��s�������in}�}��_w�W��zw�o�l|  ��қ%I� Ѡ������)P  "x�T��   ��UI�UC#�����!ꔥ   E4SeJI	�ġjJ?��������C�������uF���(JU�f_�*�
(���_��*�� ��DU8?�'ѳБ��!$k��,��:����	���
h�e�d���͒!�$с?s���c)�$���G{�\�!s��(���B@3O5�g&�~����_�>�Q 5`��bD�D��`�"�hP4&&���8�h���A���"H!#� ��>P"H�ql܆��@��
b)�U~�<�L� '�_@�}5d�p�d�� �#�fYs�T�MB��������j�d��J��cQP$*W�����n-=uX������3S$�6Mg/`S|��T4���D�4�m`T4�D�H�����bSI�v�8�)V��k��b�y�$��>�¡ �@	g�~�`D�d���c A�F$,���Ỏ���@#��vL`�Id4c��dF�q6��`SF8m����ͻLO�� P4�F��)�$�2(>.�z������g�o��ד�NƆ���u8S�κ!�l�0�,-�&�� o�nh�k���Sg+��
~5^�k'ߠ#����x,hh�xsa,�J��v����ja���HQ�!@ӆ͘r0��CN;Û!C%t2��ݸp�;�?�RC�$�3��Ħ�1&��5M$`BM�ђa�ݡ�Е�d7�Yk7iM��a.��7.�a5.�vm-��L�ؖXD���v�^�k��~Pz�(,P����$��!ZR�1$"�H�*P~�!WP���!Id�L�I@�:M1֤�n�l�3+2.R�BB�[[
@���� 0x��"@H��au�ڏ3i�BBBaVBYEL(0`Q��+Ǥ!�� ^o9�dS�͓$$�cH�37$�]�X0��E�S��6�D��H�0Ԅ,��Yo9����`��`C_����5H�Tʦ��m��;��}Q1I����z��@i���!u���u�����xo�!�@~2~�Xa�Y�)`Q�,����#VX٢�u��	%:�遠��D��C�~%Ma���0���5w�N~��u��~tm���	tt�8?!�6!h�{0'�]𔿶S�`P��#���%tS��#�i��,HC�̆��c,tHE�
B[$X1� ;$hic0"l �B4d�"��$�������`� ر���������x�
�0�nBpcV:"`l9��c�NAk�d�M���JD�(iǉ��#SQ!�C�E8�"A�4�j��$A�0!#�XB@ӄ�DdJGP$p6��v�f�4qN��tI��d?8@����,-����B��xD�ƌ4�ͼ^q�tm�7�!RtC��|✒:��i�%�0	!��7N�$�8@�H�L�`��,4�.�]�I�.��Y�"�
;P�F��Ġi XO߳���kd8IP� �d �����C�6�I
�� �C�9��B����9�
a�#!xA8�Y�N����Xc,�u��ʤ-���$�*B�%'6�����[/!K�aZjB�,d�%�u��x~i�t���x��=��*�~La��ԑ�(�"�B�!cIR0�!XхX`R P�	H�H+��2I ��$n��8��Ee�Յi���ќ��>�ۋ��AҐB	H�;P�SK�R.�o��%t����ٰ�!Mf�?St��޵���xpRDӃF�cA"�4Ji.����*�p6/�l#]of� �4``�vZ��n�<����A����4P_¯��:����M8K�,�а����CP��b��
B����l���!t~Iteܘh��o!�g?�*B�M�
J�H@������l#M8��`c�V�bm�4aCd#�ƢhR%4��E����āMaw1��)��0H�HЍCK���	
iX]No_�q��s3�f���oY�S���!$#R��`F��V4Ѥ�D4���؜!SH`���~HsG��?+UTy������[���	R%8_�
�����VB,u
i�T�E "Ađ"$v�BE((V!Z2ۛ�,?�aͤ�?$HP�D��1�$)(D��D4aϹ�M�j��|.��ߋ�*E[�۬��Z5� H�B$SS{�;��<?�a4�!HV,YYYu!(Cpx�x��,b�;�s�*B�d�8��H4����%t@���hl62J�a�;6���MHd9��B�&���?������ �,�8~�974:���b�@��&�s��1)V�� �H]Y
�B��#��q	�4�!N:����Hq�c�`@$c`�X���1��H�$8㲌
�t`l�kP�JdѣLF	�4�@B�:GA�i�u�X?|���ЗP�E���P4�5	k i �&�aB��Rj�]��	F�ѭJω%�揹
�al~~~SFB����h�,hR��������D�,>R#�sFMCq,�K��,
�:LH��c��𑮓ڑ(h44 �5��Z	B^D���.f��M�XB/�#FP�֠�@�.��$B�)�n�
�˳�J���6�nhy��IK�����8K'+�sL���w��ą�9.���UPBS^��MU�_"�ǅ�Rs��106���xuP�zA��}�W׷��j���ERN��E7T�$�Cv�]�%/��?9��&	��:���WL�%����"@$H�Y��+��8pFta����tl�#��4�1����ȒB����p �!�
D�
A�.&;�y.�]Ͼ?)I���.$)q�É�aXSi	M�!hE����
���~�CF8~Bю�?�LH?�PҘ6p�~HWN.Ï�_��.��vR5ӎ��K���i�pӴbPӉ.�!�h�Me�]�B��f�p��"�H�8��)�K�xC/c)������Y5�CgƳ��~4 :(>�Xhֹ�l�r:4�i��Jl�4�цr��k�¤o�Y:�w�/½M������ ԟ�5�y�xe���2���]m$$�d)�4"04L]� �d6�:74˺ƗZ��K�4��6h9�P�oAw#%�Yɬ��Y�H-[�-y!�aY��ƑW�Z�`I�*:y��r��c��D"��������� AL`M	� �X!�ĩ�Z]L޾�F����]a.oD���r^!Yc�"?(vE���b`$@ Ŋ�"���쿭H%j}��~�4��B0!�!t˦]d.ss������b�5��!�)Jh��˥$$1�$et@
i!4H��a�!JO��&c��֩�%&@��m�%}UU��C�B��$�i �4B�)���Ji��	�pI���Ґ�.�620����j,^np��k6I.|s_�<.�O�Mc����9�Ȇ��B���;�s������m�]���޷ A���Mˁ�%8f�_�vpcCc��7� �n���"�������?0ћ6?,k��V��ڟD�ZS��R��{��O��A'R���SST)�"��cm�����      ���       � �                    �                           -�ċj�C�Y�,n���]��5t�-���`�``*�6�`9`ٵ�m&�rUڪ���4�C(Vж�$)Uɲ޷n�;\ kŤ�m�m�b��o,Pl*�UU@R�� Wc+�ĵ@�3���Tڴ�  :�]�/C�O��6��M6�Jpv�g@�a�[@$m$���l��V�<UF�v�j��hך�WeU^�)�;l����$��Wf����,���mU)���^XU@�����d��ݏ-�WU�.U%tUWm*�+��R"�ĝ��     $ H  �� �k�      9,� K)m ��` $e�6��` �6�fm%���f�`2,���4FHwcYE�#l�-+�@K�p�uld@,�v����,�<��kj[ j:z��9��ʅh��l�v�f�M�m�l�d��&�:�M�K��vh���m�`	1 ��&  8 8-�$m��m:@��g-�-�m��6�[[n�mH ��B�4��+Tje^�����l��N�N^$(୷j�v�UTJ�������,�VE��H�L�īMR�	�v�E����s%��ĺG	r�k�Ux:��T���m΅]r탚]�� -�:ڶ�� $`   m �@ @qm   �H        �            ���|q*��-� �el�����>n%�d�d�n�}|� ��n�r��  �ͷR�J�L�U^����[E��ۋj�h �m�[@-�6�S5]��  G���mm��up��`�m�t0�vV���7¨�!�ґ+��m&� m��Y������WR�A�Uj���ZŦ� [%�Y�[J��v��-�c��ᴛ����l   |��m�� ��"��p[]�۶�) ��j���kv�VU�����$ m\���fͫ��v����Jමm�]���`μ I ���m'M�:۶�WXcj��2�J�T���P�l��Z�Xԫ%F������r;�
��r�uQif��d�m��o���u�\Fs,�KS�	 m�p Cnͥ�p    �   �`,�&����6Z  �-��(���<[x  �cv��m���� �kp     �N� HH�#	$  ��� �[��m�,� �$ �� m�@yÀ -��`�kw6+j	[�5pv�5mWm�y9  -��%gKC.VX. h �{ﭯ�e@j��}.ʱ�c�� J�`q��l�   Kh	-� $ d��+l����d��yV�:^�p I� m��([@kX6�&�on��oG^�tVյR��4� L�O�j�[@ p  vZ@ Xvn�+�t_���e�v��m� M��'@$ [@mi~�>������8 ��-  -�s�p �ö�٭I�Ν''@�k%t�t���`8   �  	��ͬ�&-�zM	 [@�p[G-9h����lksN��檥e�.�^��  �sl�:I�IKh pݶm���"�nܶ�Y;e�F۝�Cu�ҭJ���(5V6۵��l
R@��@�	��`]Um����@ۅ�z'^�[Bιj��ieՔ�mS�� ��$�v�g}��_  �[GI'^�  m��/�k�]��[_7E:�	Cu�Dy@ [FݭU�[^�N��Q�H� �n�  �d �-`m���&�q�Mn��n�s`�h�ցĒ	m �m��ojJ�T�[UT����6��޹�p����`���6ۀ6�mIa�gZ�`  kn��q!m k�ٰhkL�p8�.��m�kt� rt�I6mm!�lH6�l�K����d�z^�� n����\H�A!��H� M�  �WcP [V�h ���-�m۶�   5�Ԡh�cFl	l$-� ��T[���  -�[%
����������ۭ ��k������   6^�kmm�	������{w� �� �         �  դ� �Um\8b�(�H   	�-;n 9�m�h   �CV�ce� $ �-�����[�6p� �@kY �J�8[@ ��` K�-�p-�u�  [BYV�u\ض��@8��l᳥-r۰�  	�i[ �h�:v�r��i�5�ۻl �Ki�s��Z6�i\�.��/(꣤m��l��!m  �`�H�3m�lm�o������  N�lݶ�`u��m���� ��[ �j�e���]�Z�e��}��hy�v��܀��0ć&�m���]�kY�C�KV�l�j�m  ۴�ܷ[���  ��[A�m� -�zK5�	 [��O�۰'@ sm�Pm&��ٷ[u�m �\j�`m� @$q"�+��o��:	     �h ZI�j�s� �pkm� m��   6��  �R�	���km�m�H �-� �[@�` 8�ֲݔ�� m��@m��m�	 $.��R�i$ �秊��l  P��m�ض��u�n�M����z�A�� ��.į1�l�p�Pp�s��lN�ݔ�޶�r�0����h �ި�wdZ�����3	Ӵ�\�m ��wg�z\��j�W�`��մ��c%��}��$� �ֻl��%ئ�y�(�j���t2��U*���m�q���] ��iZ�ՈVU�[ ݜmkͭ�t��>vzS2U�T�g��: n���PZf�kj�M�$� -��bF\�Yx�m���`������l,�&����6�C�tm����H}���P���ط[��`,5�-���E�d� m�T����!a��   m��^Z��5VyP�5UN��i/6 $8�ʜ�-*(�ezVn
�%��w`]��+`Hm��u@K�UUWU*�R����*3W�� �ku`��so-�`:B�U���[�R^�k��>6�	h	  �c�<B]&���Izk����(�$����( Rޒ�k��V�p ���pl(  �$� -��q��6�mm��k 6�]$�6[@.�AV��������!^U�����5�M&�	l9�Ŵ  Zl    �$�"v�F�mh����8������m�Z�   ж�8��n[[i-� ���nv�2�$�I�m�m��r���|<��j�:f˲eƭ��EI�a���lm�sv݂N����ۤm�h
�n���
�Ā�<�s��T <�c
:r�I���l�m�i��U����%�|�������!m)�z�A���ݶ�<�8IʚM��l��UI�U����] nz�/Z�h  �u� [#;m��#v݀q�]� ���0]��)yeJly�mv�I�  �j�ne�$ 6� �[�m�n�,��8�aV�H��U�Z�6*�)8-��%U�V��� k[�p�k6Ҭ�,�ݶ8r� %�UA���k�Yy�����-�ms���k�ݶ�Ͼ�ﭒ�6�[�EK���b�
��^� -�6ۛnnY([4�ͬ�KnpR� ����� �m�IÉ Z���[FE��:�� :/,�D��[kr�e
���J�SUU��/m� -�v�I�[��:��L��Z��	����U�6᪩�C�J�[D�  9��f����֝n��     ��m �_,�          	         6��`  6ͷa�^��Q���  �V�j�j��msm�  m� $ 
u6��    � 6    ���KՊX� [@�  ��M��9�^�$q��I�G-�᪪�,b�.�;��`�&��m�zɭ�� 	 2N�f�gk�Zհ�Ŵ$�$�8  �[[ck��-N�V���I���IͰ-�5�D��mĀ�y � �-�`vݰ6�UU@@�
�ǆ��m�Me��$[On�H�\�U�   ���n5�ՙUċmm�WuU�!��l�l!*fuU+�w��{���T��*���T�
��@uU�A ��|��؟�:(�&)`��J.(	��Ydd](�T~ڡ��������A@P�"�D�i>D�@�
�>��H�p��6���SB�� ����� .�(�ʯ���TO߅��: �G�������U�� J� AN��ڈ~���B�)06 �"��� 
���,A�(l���>MDA؂�DB*�� �������qA��*|DQӧ��1� ��+�~�W�PM Dz��� �G��?('�1@������l�C��4b�ڠ~п?(����V*��>P ��U�I �DH)�~'P4�,X<���u �~@C�@B"$�,b���(#�?
(/*)�z ��#���"�TDX~D�O����f�_��|qR��Q�â�S����AU����	 "tB +�{��~F� m�m�   �6�    �������k�d)�t�GF�<ͅ�eV�f2귑.�B�63(+�P*���C���h���b@�/$ڻj��J�����X8��\q2�ʼ���)�=QA�LΨ�35�y���v�;y6$�J�d5�i霷]b���� 5UUC���=�K��x볭�ͧ�����}sv�n6냇O��� � �3tl�S��F��`�q�,a�x�{\f9�`6��	���iu�;Tt�(�]i�V�2A	�{l�7;n�h�Y�$KDkcW/4�Y�J�]��m�<�M��#��2��<�����V
�n���:.ڮNz�%4���.�6.+�A�dZ�Yv�m���/cnD�\��:������tp/dZ����j.k�S�O�&6���4F��\�zm��M�6-ɺ؅y���ae�q�X1m@lf㍪\�v��K­uF*k�xsS�7+�Ӥ:�i�n��j��bɭmm�Z�_Qd-�u���l��t�1F�ܭ[��7��W�V70MRDV��6�z��P���j���n`قVqt��h�؛���ֱ�]�`x�dݞI�H�Zm ��@�%��	�!$�C��v:���٬m����ˈA�0�]v�m�3k�6t���4�����n�e��@�:�5F�X�N�)W�6��s����nZ� �<n[�����Q�b�0��'6C�gM͉�C�F�2Y#���df�3� ͷl#�J�I�0�Wy�B�.ݺ�=�틓�Hꇩrvj�Ah�v��Q�8��ۘ�D�`K0�{�X�t]��e64��K��������[�!e\��Q0����ǔm��er��F������;u�vN�vs�`�,�,Y&Pl    p[wcn���Z�m�M����L�):��t�!�-�	؈5�9A��摎D3�]�5;=r:ぐ�j`[�j�5. ���D��"�����C@+�SV-FB���%��������sN��"��nx��]����g�$���Na�X�윲�UQe��e�X.�����kSg;��;Bq��q��[t[*l=��U.��g�x n��hrv�7)�g���զb�������m�j6z��"�˃1�'������d���p!��v��[8�5r��m1������[)��h:Ki�t�ܡ��C��������ގ�9��m˔Ȣ�o㲹@݁6�s��n\���F7��cl~nO��{�s@�_�z�'�)B_H{��X�oJ���*[�J����[�|�$�"BUGUwM���j�՛���VR6N�uNSm��`N�)��Ѧ]#Lm�L�"����ᗋ1b����F�t�0=�%0߾I|�U�Lي��efU"�*�0"�`{nJ`N�)��빠qgqTV�`�Y ܍F9�L4D�p�>�����X�\r&��6��d��[�$�L�L�9�j�/��@�}w4��s@3��7rD�(�r-�]�ޕ@�EXt���iBJ2!B�D(�����V�ڰ>�n� �j�
2,�@JG����ht�0=�%0'\���%�y�x�V�0���L�F�ے��J`n�����*2)5#�xۙ�s���Ծ_|�rSw�L�F���'�Y��y뫋n�r�m��iK5���W<p���n�p��`n݃���t��SSu�Lލ0"�`{nJ`�^E�ゑd��Z{빠\���:�Z�l����;�1c���,$M�74Ձ�smXz�f�	D�(�( r�j�?"gu���I�ﻳr��+j$�$�)�I�:�Z��Lލ0"�`v
�}��(��e�^e0'\�����.����Zي���O�Ac�#$͒9��{<�LS��FܪZ�F��Hj2�lb�{ނ:�I %#��[���s��h�h�ՠz��l���b� �rc.����뒘�`
tYq�ȣ����v��ڴq
&}��V�ݵ`}ⲑ�:uC��f^e�0&ܔ����.����`Q6��D��������N�%�~$�Ȣ�1�����h=n��V����6$�(��8n��K�t��%�nD�%�vft�k��YI�w^v����b#VὋ�jU\9ne�曚k�r��Vޭٰ7+vy$���޵`g��KID91)�I�:�Z�h��s��hw�����<��G"�/\�����.����픮"%92bR8�&f.�י�\���:�Z�h���?52�H5��՛����I{t�mwM��f�ܓ���@�H��1dH�0/T%WB� ��"�#�$رE�D
������~~ߖ��.�3���ٌvn�դ��X���ۖ�q��)����m�S���t`�㮑��֨������v1	���;�_�>`×���=�}v3Zy�Ӯ5��P��L����g7��^��4��/N*U��q^�ʹ	�����)ܚc�zJ��N9̛Ź�=J]/�7�<[l�8�Y6	Лh��V޶
�p���&i�&��,!��GK@l��k��Ҫ�2�$M�5�V��y��8[Tu�ա��WM��3+�l�ݛ�͵�	(�CV���9|�xO�q�7F܋@�v���&f����Z�>�ǹ{Ȝ�`�7"�dcqh������:�Zk�h혱��H�d�Ȝ�ˤi��)���$��ޞL���ƢJ!ɉL�L�9�j�;]���Ѧ.���!��_���EUA�lD�vK����[�:��cr+gX�.v�7(�(cs ��L��G"�����7z4���4��ܔ�=���²򩙣f�Yw$����߀�)�� |	}�Z��L�ߩ����UGI-f��L�,�G&h/��λV���Z{빠�YqE��I�6�:""'����ή�=��V,ݵ�r��'�8��"c�h�ՠ}$�f�����֬�[�`�5TҞ���u�c��M)Pu��F#i�j"ꅻY[�f��$H�V<��G4�~�n�i�ˤi��)�����J�7L�6��ni�nھJJd�Wr�=���w���|?
��F���.a�'?k���~�۹�
� O�IB��8P��}���gZ��iElE�!�j9���Z{빠{=n�λV�s�c�K$y1��h�`jލ0=�%06\��6B꾑�j��v.n^,��Z��.��ͫLn!�}��q��:�����du��W��S�Lm�Ll�07z4�;�,�����RF����v���K�͵`y{6��P���������ں̻YWy�������F���L�[�`�'$�r�S�ƛr�a�\B���+V�Z�>�ǹ�%�		���5�rnI��뙬���2�2�V�i��)���]���Ly^5���Iǉc��Y�����v(���k�<�H�-�s�l��+rAnLjdRf�λV���M����;�����h��$C�%R-�ץ�(������V�ε`}�ݛ ��c��%�<���4��s@�w�s@�]�@�l���y,���CI�e�`jލ0=�%0=� �>J�zyh��#Y��2G3@�]�@����=��V��mX�":"t�ι[������s��c9�=��&�y� $a:"�X�4OL�F��y.���g���v7������>5�7g#�Tf�1�7-\��C�t{v��@���s�8�˽���� ��볮�n����׺��6ms������,��6����lZ��Į�\A�	p��:D�t��3��.�,�s�$Gr鈚���v�E�=�F�#�7���^�=���5ɫn�xm�`�N�<Jjn��X�t�Rr��Ӯn���^�<��G�m���_���F���Lm�Lu�O��*��1f�07�4��`{�J`r�S^f$w�bː��a&H�#��b��V�[�g脢gݯ�7zՁ����F�����s�ՠr�Q��Ѧ-�� ]�W0YJ�XU9r��n=,P�w�_�7�XemZ��۸�23$sqx������@�7��r����DW-��w ��UYxQyk���{�L[Ѧ��Z/�4[Z͟�2�H4���|~��70��4�����n��Қ}빠�\DD�dRF�����뒙�|�V�F�N�09ڥ�O�q��L���|�Z{빠\���:�Z�་�)�E1��s`{ٶ����|� �w;r�f��ID,Ͱ��J�5Dҙt�[E̙��Fp���rY�o2��ap�ƭ�ۋ�W��q�672��sM�5���Հ}��`n;S���Pw�����1��i�1�����n��
d��37�X�n�g{F;�,� ��$��nI���ٹ���H~��t���@� ��e��S���f��(0i6�X�H��c-�0rԥ �X����45E4WHH���W �P� �  e�D41h��Gh��`BA�)X�#�/P5MQ (�Q5֖ILD5� ��!���P`�C@�A?t @@b����B�Q<
�J(@b���>���#��;TSH�����g���,����|P2Ε\�K�IN�U-ӛ�!D)��nI���)�$�����B��WMwM����SpSLT�g(���v���Z��Q2��g�3�]�`foZ����{�����ˣ��&Sl�B����&ӊ��&��]tu�v��$��9c�4f�S��U*��ވID�f����I.��?��j�IL���V$���܇�AM�N���`v�t���(UF�~�gВS?�~�j�=�ϢߣR���WI��4ܹ`�U9��BS�߾VЗ-��|��vrJg������t672��s]��;_�{�_D%2��`}	=���$���#)�������7��[?MK��W&]M6�SN[V�B��w?��
:���_z��~i��J���j����_�JՕ�Z�qn؍��C!$񞽡�9�\Z)t����Á����3�'_���po�����DFf���9ou�:)�����ҫ��t�)�j�!B��s��֬�D�ou� �w>�K����IN��r��M1Rm��j���}��=��6bIL�BQ��O�foZ���&Cݽ*��F��n���V�
�>����9BIL�oZ�;{�r�K�q]�p:tܴ�nl>�����6f��Q���V(S�}�`DdDo�ΕU6�e�4��t�ΚmjB�9��Hs�l�����9wΒ�8ά�n+
�i�̛��޵��;awj�v��:qTY^-c����uu��iBm�+�\;�GȪ�gRq=v�yu��:�բ���;)KU=��[n�Y�st8�psݪX��m�k��#F�㋅q	b8U��ͳ��Mk�rn��aY�A�:��NS�J�N��{�������m�Ų�b��+��������t�Hj�t�	}��kZr�h�a��v#^�"��c���o���������Q�<�y��39�]�̡���sM_)�{�Ձ���_HoWt�}	Nf����+I�*�2�i���m��Jd�Wt���=
>��޵a�Jw��V �8������u.���2oWt��ֹ%HowZ����B�e�M�ft��J2Jt��n��rINf�����У�ewM��]���6�?��?X�����:��2���[��v}Ol��Ⱥ�:��v�a��*��9S�ٺܦ�2ꚰ�!)���X��:S;�޿�r����g���$�����fY��e��jkY����{ן�H�" �J�b ������w$� �������}
�P�l���~E@��SrӪ)��?e~�7��L��֬��]���=��6b+d�L�n��N��w�L�4��ܔ��rSvbYHH�d�Ȝ�����v��ڴ��s@���u�3Md�r59�ö��mY��t��\���:���Eґ̾�~�!�D�NI��f�λV�Ι�F��`v
�)^Qx*ˬ��`{�A��Ѧ�F�ۑh�d�XG8�ci����П���7?*u�]�!�Ns9�v�I��zX9�+X�i��n�]SVJI�`z�K`{�A��Ѧ'JW�X�Jr۪*�Vޭٰ?$�{z����s@�w4v֐���"dnLO=uqm�ܕۓ[pF�·���s͞[�.9�\�e鹃�GԎdlr-���{빠w޻�:�Z�ȿ�pNF�FL���ѧ�|�Q]Ѧ���d혲�"�,$��9�}빠s�ՠs�S@�}w4xtV�J4��v�3�rS�2ލ0���%�	G�B�O5���-�(�')�)���/2��`ZI-ޞ^�Ѧ��Z��dY�Ac�#!8������x��΍�U�´�]6Gj2�m��9�m#ɍ�8�gƁ�z�h�h�S@�����cd�(�4wF�ے�� ��� �ҕ��H�Icrf�λV��e4��fb]�4{�s@�Wn�$$���D����d�`{nJ`yK���q���G����S@��w4uڴ[)�TZ��rF�rI>Sj��I�/b*��d��,q��-��:F�t��������M�:��n���2n��cM��jx������P+��24�����yյ��r�+�4gk��h���r��U�Y�����70�iE^݇���^�]� ;V͉�4��nݶ�(�ݎ�K�����ة���qb�n�Y��1��YBv�������f�5�U��������.h�n�-$j�;;f�i�jB���=8�ֵ�;Lpdx��3����z����?�����rS�d?���_zúg�п°b�F���$��v��?f~�H�s����Ł��j�����1�b���̦��07{ ����ղ= �����1��h�4�0=[%��%�յ2��0Ĕ6HҎC@��w4.��[)�w������$�Ci���M8�y��<v|��&��nsۡj��mF� ����Ts��4Gܙ�s�ՠr�M�����z�h����$�d��ȴZ���	,Qz����,����V���(Jd����tʦ�:r�`{���33mY�	L�+�lw>,{Z��H r(9���z�h�h��a�
s6��=�q<�%Ժ�tʤ�b`{nJ`zL�w��0;����u�l�m[9�\��Ocn4unpup*u���`t�N���wq��;�:دYu��^vd��`wti��V�rՎ�H�$S����R��S&����]�`n���9�+a��l����m��:�Zw�~ȏDDBBU[��l{��fʨt7H$�1�3Cs�����V���Z{�M�w4ev��A�G269�%�L��L	$i��)�l�J����3a���Bbv�0��t�*ƶ3D�K�\�Y�����3e��VX�����4��ܔ�����J�$q r(9#�@����߿~H�]�@�v��~�@��\�Q(ӎ�����ܔ�������4�3��,2,��Q��Z�ՠw�ݻ�w�����M��_�0�� �`� �  0`@��HF D ��@��h Ecb�X�����_u!�����$�﩮Ndt��t�́�Vl�wmX�h�V������2H�7b5��I��.��d����bW#�z{h���ӉF�C2�#JI�m��:�́�[��!%�eoM�{w�T:��:*�Vޭپ��"d��3+ztm��9�ۃ�I���Z�ݛެٳ�\�UOwZ�=��6�_�Tc�����;��m��>�n͇(I)�}�`fsR���s!N(9#�@����v��j�;��w$�!� >P=#J�M��z��\��K�0H�	#��@��� v�Z��M���C�,�JH�����,��>x�4$X����Q4$!a���P A=�Q�4a$`� � "#�����B��] Ěh0�1	B�ST�UHX`��dX"F$p �"�4	��#RQ#$GHB��֥�`��1`B)$�sl�B,�"���%V
E��!a��`nA�`YJR��(��'8CP�d�t@4�EX1�$$B"�0��Bߜ�UV6�m�� ��   o[@�>   �A�+�+=�j�����-��y�/Ny�b.���r�χZ�}�gQd����:�[^I��,쳵� ��ShmÛi��q�U������Y�]*�j��0e��Ԍ:����U�x�R���L�s�M��|��v�t��W;st4�WUU+�2U@=�.M��^ҥ�ק�I.���n7,gu�����m�:{0����B�I�B���0@��q�����N^3u�n-�B:y�֝��X
�V��ںT�>������T�^�j��֨U;U��+9ndd�$�;Gl�gc��T88,���,g��G@;-���$P#�n΋+�����'\����� nڼ�[�K�Ӷ�Aea�kP���]��&-��ѵ�,��	K��5�y:��dSH�w[��w[�nG��s�O*n�R�Ԫez��k&�ו�@jv�XZ�i���V0!+�ۖ�I�^X�rn�$��mz܊N6窑�\�v�knl���)h�PlUoj�:W#c2���kF{��>k�ݽ��z���0��٥tT�V:�FyY���BZ��%�e�U�fw���IdZ�=by���ݵH�dI(�i5�Ē'ns6IM���ip��)<�k�ld��V81ӲM���f���Q���a��]]�W�rY9��|@�����]�.+RɈ4Vӯ<3%^q;��f3�f���vt1,h�|��<݊u�#�`�,��fH���Q/Y
�܁9��S ,����9�n���U��@�ݶcv"�]vn�mt�`d� �(���a�M�w-@P,z\�4Om&�%ol�s�k<n�yH�`=;���kuMN�2=,�ˮ�\J�j�
\�7�Gl���赏�����@��ޠ   -��[m7X� ��� ��X�k�WN���zW.�� ������%e1�ܭP]�ygWYL�[�ɣV���6/�uH�6
&�<PN�S�������\����332@]/9���}��ä���\KNm�:v	��c(�n��\ݪkyd��V���f�鞍���q�n66f�ݕ��΢$9���^�["6�hȥ�E�/�G�H"r3��u�����-��9"XӴēE��+t��u]E3�aބ�;u���z���ŗ+ η`�]v�m��u��NYϱ����Ye�Kz�)�΢\u'n]����غ�yz��@�N�J5�ck��F�nt���eC[x���-�-�ŋ��H͗������_��K���ҘH� [��`��S��Ḿ�[����3+zl��ցλV�s�c��E��c�8���f��ݵg%	Dϲ�����2s��cd�)$Z��hVנZ�Z��Z�z��$k	$�nD��ܔ��|��L��L	$i�w�����u=\�����e��N�<Ni�S����;�9np��7C���>�a�n�9�k�h��Z��h�h�eY�86��D�zz�V��3��QD@�(�2{�Ձ�����|�%2n�R���r�Sr�mӛ��4�ڒ["���&0;�J`o�E�Q(ӎ�f��mzm�@��ٰ�J'���`3�9��cT�.���`IrS���4�ڒ[�gpy��]Ց�X�+۱����#TG$�/.T�F�qH�l���zh�yYÎ-�v��w4�k�>ΰ���Z���郙l���@��s@��ڰ3kvl�ݛ舙6s�ʨt6*m�ESj����3kvl��B�JQ�	(�_}�Y�;3�Xx׬�d�x���)����d$i��۵@9�ʲ#pm��Q�����j���`z\���rSw�R�U��=����.x�ѭIu��k�Y�o2�[aN]K�ۇ�W��q��c�h�Eo�o�߱���K����`N�)E�pQ��M�f�λV���Z{�M��� ����ȡ1�j9��\����7䪫�4��ܔ��JYH�"��di����S@�w4w]�ܜF��;J�!g����ֱ郙n(ҍ�@�w4uڴyڴ�Қ�^U��G �j! ��d��8��p�6�J�q%iԺ������d��$�ϧV촺k�m�?�ߧ�뒘ݐߒ�wF��d�_�d�ȣ�h�o��#�ύ����s�ՠs�J�#$pM�Lr-{��0=�%0=�%07f*W>�ŋ�C@�w4yڴyڴ��s@�]\��MH��$��rS|�ٗ)��Ѧ�F��_|�@�*�w��^�4kZ����À�u�2���wAB��V���+��i���j���\��b�YI㧣�IRh�n�4�����.���fʫnہ.�4�c�:�j�ܐ���7b�v��g˞��Z�y���}rs��P:ݼ�ևp��^�&�[ۜ�d|̷Khv�z�R�7f4���nP��8���lK[��tܭl�K�?���|P���*�{q�����u���펵efY�pdv���a��2O��;�Dk���N�nh���6!�j��Ժnx�_ߦ��fڰ=����D}!��=�)��r�n�SR����WД(S&n���]έ$�=-\�IWkX��̆7i) jI.�י�$��=J�co�m\�Iz��Ԓ]vر�����ɜ�I/;cԒ\��s�%�]�Ԓ]��3�I%����H'�9�G$z�K���q$���K���s�$��RIrہ������+����mu>I�I٪a��%�6�I�r�ld�m���M��vV�����jI.�י�$��;��q��lڹĒ��Aa�8�c�AȜI%�z�9� PLPD˖��{5�m��{ל�g3n��"���gq�+�E2�MKsU�I��I/?��RIs���$��wCRIw޼�q$��,(Lp��H�$�=-\�I{�t5$�}���_g��ߧ�G�$�o��҉�pr2	ȹĒ���jI/�߳?[�s�I%����I.zZ�Ē�7����lm�c��3Nf%���D��Vι�,i�q��Ƣe��:�<�V��n]M�#��$��^g8�K���$�=-\�I{�t5$�]�,�$1�$�rg8�K���������g�.q$��t5$�}���Igl���	�G$z�K�����߾��&��@�}D�7���9ĒU���$�=Vב#�O$�6�\�I{�t5$�}���Iu�����3�c}��˜I+dA��"�9��Ԓ]��3�I%�lz�K��Nq$���^�~�Do�Yi&!��r���됂�XJ�A��F�WBG%+���ّ�y$��$��=I%�]�8�^��I%�z�9Ē3����p��H�$�=v����m�z��y��I.�cԒK��ƔO#���RC�I/z��y��I.�cԒ\��s�%nT�t�̆'�6܎�������[��9m��{٭�m���g9m�(tM1"(W[�๙���s�P�lT�n���q$�]��I+�?v��8�^��J���Ü��*��ޓV�Z�Yf���kD��S��+�bv��4#v��Gc/6�X���L�e槳��<բj ��ߟ���޻��$��^g8�K���$�3�jƌ�ē� 6�\�I{�t5$�}���Iu���祫�I+n�	�H�ŎEど$��^g8�K���$�=-\�I{�t5$��(����ƚ�7�I��K��~m��5$�}��%�]�Ԓ^��9Ē3����p�RI5$����%�]�Ԓ^��9ĒK�ɩ$���������~���@
�'+�ܭ��H���cU������ŧYA�&�'�j.��Tm���Å�
�i�7	$j,v� ��U�:��+�
����ܤ�g���䋝��VѺ��ĻY6�j�g�n�<<��=qP�k����cY�:-�2�n��<��p��(p��Zی!]���m�k��[m�К,p�6��n~��O��[�rL�Yrj��jK�In�k~?��Q�����"A`�$��LX0�I'��9⫗:�­�h�ZU^$�Y��fG\�=6i#q��RK���jI/[y��I%�dԒK���$��Rɿ�2�H�r8�K��g9�߳i.�&��W��q$���K϶ŏ�d�9$�nL�I.�&��^��q$���K��g8�K�W��9x�Y��I%�l�K޻��$�m�s�$��RIs-��$pI�p��I{�t5$����q$�]��I%�l�K�33�7쭴��>N<��Bcv6������x6�든gQm�#Q�SZk7NvEӹ��9R��c�L=33=���q$�]��I%�l�K޻��$���c�LjD܊L�Iu����~��X�DBL�Z���r�{�orn�o޷��$��u���C�(�rG�$��I/z����s�$��RI._&\mF���d�8�ė3�f?z�$���s�$��RIu�_8�U�36~�by#j9RI{��9Ē]vǩ$��I/z�^�ʱ'�,�s%
ܪ��٠q�ۖ芢���Gei��T��Q�Vi��ӫ3P�w���~��$�]��%�]���g����V��3�I%���r$���9#Ԓ]v��$��wCRI{��9Ē]vǽ�����av�h�y���I/z���xs���u��+$H$��Q�����X�/�@�I#4�JX�|�B��E#p@��P�X� !� �C������h`�@�|}h����E'���� 1 �H�a����$����,bFH���)[Z����_���� ����':��6�!��� ��R�T|�6?=?
�C5��~�kv�~�~��m�"�,Y$P�8�K޷��$��=I%�m|�I{�t5$��<,w��ƤMȤ�q$�]��I.�k�W﻽ɻm�}���-�¢w�M�������S�s��W�+u���ʖ���$lc�΀[�;um�MO����>q$���K޷��339ƒ]vǩ$�|��ڍ�����|�I{�t5$��o3�I%�lz�K���Ē�љ��!O$mG jI/z�g8�K���$�l�s�%�]�ԒW��ŏ�� ��&ܙ�$��=I%�-\�I{�t����D^�;Ü�����L�e���#�=I%�-\�I{�t5$��w�����2P�T-Ӛt�P�@�s����&a��Q<�ηS��[��\
F��V{�FH����F�Z{e4z�� �m�k�h���qb�"�q���#LvL`l�)��2���ÄO�7"�4��h�զ����UñN�0<��Ҙ�+2��S�t۰��}�`fs���ݵ`��9|�q���H��N-����#w���gs�=��6D$�В����H�!$T��H"� ��!!#��������U�UE�m��7%čn�[v��$OjK*3�73�]l6f���5Z2�9�u�[jx�TyRx���/7=�MN�˺��Ѫ,F��ʹg��]1�y�u�2����7;(LN�Eۭ��[A�P�*ݺN���su���6۵��7m!n� 4ta.C�������b]ɬ�HWIR-�v���t{o�ݮ���q�wk@V��[e���&��h����{�����Ӷ�1���杔2��!˻6[5�Z��r�oI�T�N[��D�S]�e�~��`�c�2ِ`g�v�����]6檛V�n��BJ*���`ñw�LgKE�^eU����Yy���̃vd�`�f����F8����9$4��07z4�7d��d;%�3/)R���//�F����̃���{�c��`Ҙ��8�Y##�.g��u�6�M�:F��=wkn��۵GE�of<jD܊L��٠s�S@�l�����hκ�;�JD9�(��h�.���$$�ED(�J��o�ٽy��@�L~ƕn'##R8h� ���� ݓِ`N]T����iIr8hw}w {l�9���zx�;�����c�JInL��1����07z4��_\�v4�ʋ���I-W�X��q9��ONSF�H'#t�`���3��k%�W�=� �ݙ�F����ْ���)��;�)�w�����4v�h���8�ō�	#�䟿}ݛ�O߻���+��b�8I%*#�%\�>,�^��ZJ�!�'�H��I���4v�h��;�]���Z�p�H�?%RM�2ِ`n�� ݓ�d���>�wVF�n݈:�n��n*#��.^Mt;=DƮ�
�ݒ`�IM����`�cvd�u�Y���iIRC@�m��v٠w�S@�����\X�Lr	I"�I��&07nJ`l�vF�N����&�M9t�6�:st����=��V��)(Ten�k�U"�L��Y�^^e06vA��Ѧ�&0=�"�;�pi-C&1LJ8����dlyz�'2�B�#�!�y�v�A�]�ն\۵���9�X�8�$p�;�]� �m�:�Z{e4��e�<jD܊L���`{nJ`ñw�L-�t�#)H�?%RM�v����{빠�@���A�8�JDF��h��07z4�7d������3�!Ғ5�����h{l�9�j�=�zX�$���DD%���:UT�7U	��ǳ�چN��&�vs���k�n�6^�3A��=�ol�I:�9������Mv���;{]����(�F��{;�Wi�9�ط���qqh咮�:Ӫ��J�1�Y볮�:��\5��n����{pS��D�� MƋ(�;��jn-١�27F��6΅�9�g;/�|/��#<�dW��e��Nפ���El���;�����q��f�v�S�'k7;1y�hڬ�V�z�u.�rm�-�dERG��d�5$�7&x���snJ`ñw�LgKE�^aWe[���`}�ݛ�2fs���޵`��@�v���6�"r-����F���ڒ[gdT�]�,�)�ܶ��N�w��3;����ڰ�
s:��;��)�S�uHt�t�V�&06���ݙt�0?�߭uC���n�����7e�7s�8�Ρ.%�3נwV���b�;��������N~v���r��:�������`fn������VO��8��nǠw�S����UC� ֧{�lܒw��nI�����%
d��(\�leT�n��e���j�7d�Ԓ�� ���e+�,ŅM6��6�:"�gs�2{��{^��%;��+ �ޤT�US4�:m��ݫ�DD,�>w�Հg�]�������B��	��y먀�1G��ݹ��^ީ��^֭i��y{��;���_M�B�H����{�>4z�� �m�U����<nc�FH���n��B�2������=�z_B�Jd���D�8�o�8㙠��M���T ���m���ܓ�ݛ�p����9�dӉ�.[v�BS���`fs���ݵa�"!D�gs�=�)�P�S����X��,�DF�w����u[^�{�<�
�c�Y#�5Z��P$<s�;ui�z�ȴ�Z3�1��fuN�~���s�tfl�HA���G!�-��� �m�U����*�c��L�NH�m� ��]�J!/����߿U����,z�� ��xу�m��o#�hWv�{^�tDDL��Z���`|��iT�����[��S�Q��ξ,����'���nH��T`��$z"���Ձ�תU*��Ҥ�n[t�3vՁ�DB����=�V��K����l�x�'VZI�r�H��@��Vuc��M<��!#�z�5�͡�2���LvL`mI-��2��$�A/�nh�?�?�$����)&��mw�%�DBUF����;�~�`��Тd�l��C��nJ�:u`fs���ݵg�Q
&L��`d�uX��
��MHۙuL���S�����`zwv�?DDD�u�`t�s�Q-4ʚmӪx���ڒ[vd�4��|ӈH�@�$�k_��`oH�6��l���L�F�R�x,�`&�=�"A�$`�bD��!��6���|�H�!���d��H%�֨��� mpJ�����"0/M<F%?)4��A;���*H�v*��*�� �	�<�@`�W�@4�9EE��* i H�$"H�p�%�+l��2�XT�)��R��=�{���?���   8   ���    ��k�#]�Ihl�i�v���W[�DgA��)\n,�P"k���((t�/)�j˹�c�*uע���6��K.I*�Wf��խ�i�=4��S�Kyf�z$�r8�(m&z�ɳt�Cmk��<v���۷]mI��HK�r��s���7[l� �耫������ u�l��NպmW�n�`��N ��\i�s�ll�=P��*�ö�e;��J�T�a6���a�Lv;."A��vL۵[XKMg��m���
���@R=%�Q[pݦ��m�n� QO��I��-v.��{g)�nR	�ز�3���`�����^�<�z�l�b��I6dCeٶ�o%k�ѧUPNS�]\�ˇtU��h�\u�;V��l�-��@��v!�xN�g��m�4!����ag�`�!�<k������l�v�-ѩ��:�d�Ӓ���n��zGl�y����Nj1:A�P2��ǐ�\�	-R�%,�UJ��Ul����.��Us�lm�	m���*��S��*J� ��U����
�N{d�v�*U����0tJMۙ�@�ӹ��"v�ݺt�Y�R�&�6d�4-N��NѺs��mA�v�8ԭp/+��\qӢc;-��9���qГ�r+9��βi۬�:
-դ��xS:�/��<���l�m�nX�������u��Q����xV����
�g=	$�L��6܍�@m0��xG��1e��`1��������ڛS�t�6��* �� ,��+�������J�UM������v,u/�7Yevx�L"&�	9ۖ�pv��)4v����.j��!��6��U|�H{`�/V�qсd%��ӛ���Q���6���"�ڡ'Bcʇ�/.�ų�J��dXN��� �c  � 2
��h:M��f�[���l�v�9W
6)g<F&����� �q��'<Y��ݍl�Sʕ>4Vv�����/T4*�t @O��D�Ҋ`� �mT)���O���{��޹�<�UU&3���k��ej��\�N��cv��ЗIuW	��٥�Z����-�ݧv�c�룰�nڣv;Y�ݻ���v(Mj�N�ڹR�N�*��C�o�J�M�c�;���v1����	�zK[j��	M*ݵ�یC�h��9�n���ۍ�dٱ$m�[�ؙ]���ȚCk8ڶ�D�c8�Y�r��һLg�{q�g�a�pr�θ�m̯K��0͒����ݚ!�mg���W<�=�rVܙ�;�ݯ�><�� �I��G$�V����h���!B�@��v�s�U"�nj���sW��ݙt�0�1��$���I����UMS�JZn[t�w�Հ{d��d� ���,Xeb˴Sj�tՇ(���v����KS��s4���&'?%RM���ِ`n�i�nɌ��ʺ��ʯ�@l�;7�Z�]�iÎ9)�.uǅ^m��m�P����?����4\�qf������������� ݓِ`J�,Z�leT˧C���͵�,�iB��P��BP��Q�u۰>�>,{^�Тɳ�ΕC��U:m�Sj�3;�����g��|X�֬s6UH�l���sT�6�?D(J}�|X���=��V�g3��YϩT�����[��fِ`n�i�nɌl�0�q�������uv������]y�&ў��N���2�Ƥ
H��gM�<�g����x07z4�7d������;�g��g�ǐ�A���f�w���v����{빿��?�?�LND˗-��ϋ�ץ�����P���z���~�}�f����nI�䧥JsNSi�*��saДNg_t�� ݓے���ό�
�32�/0`n�i�nɌm�Lِ���Ͽ{���KGRZ�&�mC���b�W��C��y��{e07�9�f5�s3/2�0�1��)��2ލh��ƌ�m��c�h�o�3�f�� ����%�O,�ԩԉ�'qȴ{��w���|�����Wt��z�R��t�F�St��F���ے�bK��/��bO%��,�|J�i�M"�Tۦ���ے�� ������/{�ߧ|PR�6�m��&.�2��k�E��9[@�.0<����g7hk���+fg�޿ߩ��2ލ0[,�_,tk"qd�"$�@�l��
Q�DU��Հj�ߝ���vl�X�Y���iG�����hs��>J��ewM����3&V؊eS�ۦ� ���`}�ݛۏK�Q�޿s4��0r��ɎI�snJ`l�w�L�Ɍ���ߗ��������g��	��
q�sڈY�4룶���:Уxd6�,�7e�����]�\�a�:��@���dq!�C���mHg�$�F���cJvr���M<= e�뇤�n�شI�Fq9zٷN�Fd5 �2�6d
H�-��XK��2�mSe��u,l���{&�9,,elNaz2�đ�wF6�qMø����a�i.����n]n:m� �� �~��2�4f�3�n̈́�[T�����[�"4hI�.u�V8�m��#ƌjD��8�]�g�w������Д(�C�]�`vW)T��M�#c)�e��fڿДD�b��`{+�l{^��BQ2f��UCn\�"��ܶ�.���%3~��e� ݑ���I��)���5L:S�=ٰ;9��ݑ��d���\.�U�,řE�6��K�Fgw��Y���v��`ő8�)�����`�^;<䅳X�r��Bݲ9ȕ�kPt�^ո̺���`�L`z����I}������h���g��2d�IRf�j�1��*��$��d�����,h������ɎI�u}��@�l���z�hs����+ƌjD��9�ua�}Ϻl��V�3]����X���rcD�#N-����]��%�=.J`wE�Եt�Uq3��l�r]�{Wn<�$d���<��kў[v[��>���0�]�m�������[��wF��_E�*�Ӊ��m�mn��Q	%2{��l��V�3]򈄡L�vʮ*\�:T�rS�NluwM���j�Q	TBYj$�_B�Rr��`{��l�YR���ʪ�̼���wF�.�K��~I(�s���WX�i�Ժm�rڰ]��%0=.J`wti���U��<���M[lt��n��9��SWJu��d	�9F�1��1���#�5�K�������� ��1��2�hƤM�H�$�h-�~���m�s@�oۚ+�o߿�/����rbCc�n���֬Y�j��kvl�h�T��H�oq����o���]�`n��� P(^X�DV��-߫�ϲA8�HbO$s4Wj�I1��Ѧ.��r,U*a�+VF�nݺz�;�.�y��9u��*��O<��4r�6H��336���߷�;�4���`z\���g])���$n7&��z�h�z�h�ՠn�IB�;�eu�M1�-�T�`j��V�[�gBI)���wzՀv՗Ә��72)3C�1w���@���`ffڰ��BQ9������ԪEJD��rI�Wmz���߹��֬��f���(����ΩU6��ۅg��s���kv]���W�ӰmŮ��KkKۥ�Z4[�UjU�ۜb�4�je�;u�����{^U��q��G82󵣍�eN���#Å8��wD�'#!ۖ��H����mx���4)��N�J�V57X�V�rPv8c�=+�`��Ɇ���LN�s+��
k�1ND���t�XA������d�Hv�ջ;��{.�>ez���s��u��gNi��k#���[��_+#�:{p�u{BܻF������������;����>����3u��Pۗ5Jf�Srڰ=�m��	)�3�NwU��nڿ�&N��(��4�Kb���5`fs����-��#LS�L����u�W�f,������-��#LS�L?}
}Ϻl�6�s���S-�T�Ձ�Ѧ�Ѧ��L���۩R�/E8;QE.�����^x�[�z�u���*	7~������s�l�i�QY��r�?4���)�ղ_�_$��$��4�|��CNbln4�Ȥ�����@r"��]�S�u����Z}�ۚr��h��F5"o�:nl�nՁ�nڳ��P�qv���|��ˍ�q�C�27&���j�ř��z�fâP�}������%Cn\�)�uM�j�ř���
#1�O���`{۶��yNV��M	�^��4����4�:��I<f�w].*.��V�nn�|�{���;�V�����u[ �Ɍ�05oF�%+t2i�7%U7V��]�/В��Q����r����q[^�|�5��HA�-���vfm��ٶ��G��%DB����ňE! �#��k �Hā F#�,t��T�! E�� `���9P>CD	�T����ă������(�yK
@ѽ�Jđ��b�H�U�̠�����i(��� Ō0�H����%���	 �@bA0��T�4MJB�����@ �Cf���+�4�Q>T |"�'^s��˰z٠z��=0s ؤ�I&hfBJ'o|�OwU����`ffڰz�������i��I����߳?(Y���x��j���m���W2:��|�4�W=u�M��mۘ,�������z�*灶�Y�ܔ/%���o��ץ���j���m�I(�􇧻�����6qǉ5$��빠w;빠};�V�ץ�
ɽϦJ��ʤ��H�������mz;e4{�j�>�Nj��ʦ�L�n���I$����`{9�`ffڰ����Q�`�Q@� ?(l}��C���Y�8�2DBI���M��s@�w�s@�]�@��~W�*/��@�Oa+UVR��)��j�z�µv^��ٜ����I��"T캕V!��D�۪l����05oF��%0=� ��%Ҷ"�eQ-�-��/fھ�J�3+�l���w��h{V_Ɏbln4��-�ޭٰ>��,舅3��j�ŗ���ҬhƤM�R"dr-�����j���m�����1�M��ϕP:�M���,m�,{vՁ�"Db���fWt�{^�B��Y;ΕU6�Z����a�u���ŵ
a2WC����N#i�ԴV���7XW\��nt���š�n�N��d�����<s�N�z��n�۰88�:0q��{n�n�zn�qAp�ob�v�;v|��`�t�5�m�s��S[v�l���3mJ��;n��Y�5�b�{2�N|�]�ע�h�#�(HL&�¥n6�UY6,�P\�eN�\M)�XqA4n�%����3&���9�)�R#�U���\7G	t����r�m	��yDBJ���J��dҚ�Rܶ�V��V��Ll�07di�{�,��VR��UV�/v��d�4����ٿ�O�AjC������Me�T
�9�3?Ł�nڳ��,޵`fWt��eJ��ʢ[m�6X~�J*���Ɂ˧��%0=� ��%һM2�Kt�Ձ���VD(P�t�����j�=�-%�L�����Bڸ��n�qa�\ݪ!�mg�Jsg�5հ�\��<<�ׇ7�E�+�m������l�07di��z4���)]�˽��p�f]�9��پ�UxT~�{�L˧��%0=.+��Yx��K�S2���mX^͵gD$��ewM���Ł�ǳ%CM�iMS�n[L[Ѧ��Ll�0��_Ww��L���ϱ�Qc�bO$s4�ڴv��4�ս`��S2��e��6nJX�z�Y�lq�M�w7�y�0h.���a�!��X�2,qI�1� ﾟ��j���m��HfWt��mJ�!�$����s@�w�s@�]��������7��UX�i��[�-��]?4�ݙE���{2�`핱4SSTU:�����:'3���ϋ�ݵa�8�{�`gk�U")��UU�fffS�2�05oF��$�
"�mu:��-�sJ�CmHN�.���3F�3�4�8��6��������?~�;i�q91(���p�}��������Z;e4[*C�E#O#$Rf����W�&OuwM���33m_�2�Uk>�n,���?�Z+�l�;�֬[�j��*��ʧ9��]fK���4���a�}��Q�;� m���ܓ�teJ��ʢ[m˧6��j����~�p{��r�V�w�r��8���uĩ=W]V�����U����Gp�gv�e0VV4�C	<jG�f�������K����%����Հw~��&�j��q��E&h��9]�@�m��<�6��#�(����UH�����j���_�����X��i��fA�6⫕W��(9�@�m��=����;�4��S�}�`f��U&9l�Kt79��˺4�ݙ��L�`g���ww{����<�ڪ�Ęød�D��l�X+d�M�zq&]p�4�=[L�^%�A]`��x\���U�+Q���rNY�1�WA�u��.�F�#��g�{m��g��i���R[*�����ka�/�3���+�J�I�jH��x-���9x�x��˷�^�v&0b�,��N�m˧�Oh��/]�DJ�A�;Le�8��������{��;�������$�4kA����ys��bs��Ѩr��Y�b�X��v��{��^O�f㈃x'�9����r�V��#L]Ѧ ��)^+2��f+u�0=.J`n���ti��2���N�6�WleQ-��ӛ3�Ձ�3mY�Jg3������ݩUbH���m���~���r���`n���ڴ��� ����1�m��M���LT���%0;�4���f���7����OC=.��㜐��5b��g\1i�t$�m\
F���}�w3|97i��U2Zt��������mX�6Ձ޻V�z�'D�cR5#�h��W��IU������`}��6n��ǐ�F�FH����]����Wj�=�]� ��/5�D��<�����J#�Z���3�~�6��j��{�s@3ǭX�2,qI�"�M��́�/�~����9w~�`��`n����m��R�Uv]�7l���@"�eQ�3�K�QT鳙�^�Љ������09wF��1��rS=�R��4��)�r�j�ř���D�vw;�]�`nfڰ͕�4SUEU75M�ڰ��>�ݛ?D(3�Q�A6�U � "A �!d"�*'������7!�����V4a���M��)�;�L�L����\*�m���Y-�s`g�mX�%�B�]߻��}?��ڴwхx�LiP7<stY��t���&y�͉�t�`�G�y�Ǝ�\�� ����"���H���{=빠{q�`}��=��Cs�Հdl�J�Qc��G3@�~�@�v�ݷr�ř����-7�U5NeS�qP6���s���nڳ�%�qf��:�����y�t�B��܆��۹�w;�䟻��w'� �@@�[���Ł��uJ��sH���m��ٶ�/�0=� �푦��X���:-\�`����ul�9��^&�z4�n'�l1ׇ7.V��+�m���S�2���_/�A˧��O�4a��19���Mݷs@��m�ӹ�|�BJd�S\M6�UY�XVx0'~��V�i��:[�ץ���jU&9n����n[V�P�o|��ޛ�k���)���XyV��qc��G3@�~�@�u�`g�mX^͵`B[Ȋ��>��ī�$P��YtK�$��$�%�İچ��ڈ��H�R��@��a�1(@:mr�GP]�����B0g�,ځ#��� D�.�D E*hU��6@��JPJ�`Ab�o^�_N��N�N������8�`      ڛ\    $��h7N� m/!��s���i���/�m���U]�i2�#Y�;l�����C�Q6��@�M��R�.�H,��l(�'[F7�$'f��b���gF��r��F�Ց���m���uRj5�"Y�,v��ul��u���n^�TGܤ�T�E 5U{T˥�#kK���e6<3Q��8�ݱl8C���r�[�!aej����5�#2�L�:��٤�u�z*n|��k�w[v-U �U@T$؝���yyK�^��3:t5�t'ҹ7N��^q�v��ɳnSn�+<�� ;c���k�u�����4[���5���U���E�n�1ػ*������Z� 䦏˞���`����}�Y
]����n�n��
���];I�	���Q��Om"�ΡB��{۵A��q�y�b7CuhՍ��m�u�I��W8;l��a�Q#�mn3���.:݇��B���-B���
B @UR��j����]�j�=��K*%ЁƇn�.�WN!��Q�^�)g�g�����;yb��Zeb�g�'WI�"�knB���6��2c3�CKS�j[�Ժ�Vwk;uF����6���`���*8�ݞ�1�ץ�lQ]�s��������c\�oT�;P���n�4������J�j�^
y�m������-�PI�����t�\�6�4�,�ڡ��f�U�$��]�:fq��#l�k��;fސA�9f��VӻMXjr*���t��g��]���<-mʄ�[��[[:��PX�7f&v��`�����5�ǯ�W A��ᎃp�=e�%�DD�m�0$�LmJ���78Ab�}�ս��d�<:6�C��m��6�� l I��Q�^��mㄫUYȺn�=V�),m��k�L��$�K��n�=E��m�n%�d��e.��-����N
�P:���A�� t4�sb�T�Q'��=W�uT]��A⮕�+ >�*�������k��33V�32j�!�tpڜ9[��D�؆ɖ��5
I����W���Z�zL�A�p���Id�qw&��.:t�qr�	�89uvlۃl�khܑą�]5����[mҝv�����l�N��ܦ�q�{9�vp�X3�mv����n:d�v0��$v�������k�ê�㗞k>|��Ϣ*�[Y�ɺ�]�tIs-��"~BC��Nf��FLɫ��AD��m��ض��5k:�c7�)+�g���٢ەN�2S�qP6� �c���nڰ<��k�P�%	%����`~�]R����̬˼���#L[Ѧ��X{^��	(�3��UX���E7.[x��~i���l�0;di�n՗�c�؛�G2)3@������M=�jÒJ��������^e�3�d�`jލ0']�@�m�4��2%0Q���̉5m���d���@�����^t�X��\�g�����ϟ>p�M�1)��p�_���;����9���	/�=���3w�J��-�J�`�k�?������K'�!Dͮo=,{6��J�z2v�r��1ǉ�nf��}>4v�h�����g�ڱ�pC��`ԑh{^�f��ٶ�:"'+����խc�"�"��޷s@�w�s@궽���EU�BX2CpZ[�zcM$�t��+'9��]rzR��	7t(v�U�i��Sr��k�1f��jIll�0;�i�n�S�0�*�2��ef&Ԓ�ِ`wH�V�ھ�'�_J�骥T܍�n�gg��}����o�"��DBX�P�BJ�X�Ձ��vln=S_��x��AB8h���s���;�K�(_�(���~,��jU&9l�W�������z4��̃�2�]��;��#�&d�n�h�u'��[t4�Q�i.x��H�]T܉iM�����:M̲�t�D���^ξ.�)!I
b~����r%�bX�}�p�($�Q,K�}��iȖ%�bSӿ����f����v��bX�'ｿM�"X�%����6��bX�'����"X�%���޻N@[ı=���=���r�Se���$)!Iw��p�ı,O���ND�,K�g�v��bX�'�g�v��bX�'���Mrˢk2��fND�,K�{�ND�,K��ߦӑ,K�����ӑ,Kȿ"T"w^��"X���~���nmK��������"X�'ｿM�"X�%����]�"X�%�����"X�%�ӽ��"�oq������~(�M$���]Dh�y� ����S�;#ֆ{s��xm3G&��UI���m����$)!I����}ı,N����Kı:w���,K����]�"X�%����L��h�YnK��˴�Kı;�{�Ӑ���j%������Kı>����ӑ,K�����ӑ?�j&����߾���-�J�`ۦ��)!H�'�{��ӑ,K������K����g���r%�bX�￸m9ı,K���S�e�55�.a5�6��bY���O�����Kı>�����Kı>����K������ӑ,Kħg��5��Y���B��iȖ%�b~�{�iȖ%�a��)��ߍ��%�bx���m9ı,O����r%�bX��`�	='��'�OO������.����#�nW�{vܩ�X��M�V�Cm]�̥,���i��۶��H����ݲ�g��3�;뵷4�r�Vԛۻ6�8Ρ�lE��]/-��Ԙ�#f;��WiB��Ů�Z����]�ƹ��y�F㛍-�y��+��v�>H�]�9wn��k�Vu��v/L������֧�q¸�|P��@I���[8D�4Β5�������8�3�p�b����mr��^yL;a��uϕJ�t�ٕ]sFZ�n���ڂ��#}߻�oq�������p�r%�bX�;�p�r%�bX����6 ��bX�'�g�v��bX�'}�j��&�D�e˚�6��bX�'N��6��bX�'ｿM�"X�%����]�"X�%�����"X�%�{�S�k&]j�k2��5�m9ı,O�{~�ND�,K��޻ND�P,K��ND�,K�{�ND�RB��죠t�R��:�\/�RAbX�����r%�bX�}�p�r%�bX�;�p�r%�bb~����r%�bX���]3Z�Rk2乚̻ND�,K��ND�,K�>=�����Kı>����ӑ,K�����ӑ,K�����2e�˪fMk.\5n9r��4RHl��t�K���%�B��Z9*�!I�[*�:hm�W����$-[�p�r%�bX����6��bX�'�g�v��%�bX�}�p�r%�bX��:����L��&�-���
HRB�?}��m9�D? <"�i�Mı>�����Kı>���m9ı,O�;�ND�,K��3%�ˬ�!��6��bX�'��}v��bX�'�w�6��`
X�'���"X�%���o�iȖ%�bw�m7�f[�$�˭f���9ı,O��m9ı,O�;�ND�,K��ߦӑ,K����ӑ,K���S\��2�̹sY�ӑ,K��Ӿ��KıD�{~�ND�,K�s��ND�,K��ND�,K��I�1�s#�]m\[s=sFp<�\��m��n���=d�ێ�F1��ꎽ6����a��Kı?}��m9ı,O����9ı,O��m9ı,O�7�W����$/c�G@骤6�6;�6��bX�'��}v���1MD�K����"X�%���p�r%�bX����6��bX�'�w~.��f�5�r\�f]�"X�%�����"X�%���}�iȖ0�@����P_�?��?�ı=���m9ı,O}�޻ND�,K��ܲhɗ2kF�XL��ND�,TB��Ӿ�ӑ,K������Kı?w;��Kı>����Kı/ޞצ�Ze:�N����)!I
H^ξ."X�%����]�"X�%�����"X�%���}ͧ"X�%�~��O�
��f�k�"s3Չg t���Nn(�pqh�]�X�Xv�����{u�����a�M\̻O�,K������Kı;�{�ӑ,K��Ӿ�ӑ,K���t�/�RB����e_!�X��̹�iȖ%�bw���! ��$���}��$�}�{�hH��Ͼ�&���SQ,O���O�Ba�u&�.���a��Kı>���m9ı,O����r%�bX�����r%�bX���iȖ%�b^���s.[5�f[���r%�g��N�o���9ı,O����6��bX�'{�p�r%�`u�H
�@�B�G7^=��ӑ,K����O35��e�.fL̻ND�,K���M�"X�%����6��bX�'zw�6��bX�'��z�9ı,O�w���YL4觡�U��x��ӕ�m%zv�cH��Rp�&UY��Fm+�w����v��]�^��Q��O�,K�����m9ı,N��m9ı,O��{[ND�,K����_��$)!ow}!I�[&�t��5�ӑ,K��N��ӑ,K��^����Kı?{���r%�bX���i�")bX�%���zkW��SY�&0�r%�bX�k�����bX�'�{~�ND�,K���m9ı,O���ND�,K��3%�ˬ�&�Y��r%�bX����6��bX�'{�p�r%�bX�w�6��bX�-����kiȖ%�b{��߈���r�����$-����Kı>>�m9ı,O�g�v��bX�'ｿM�"X�%��螿g������vsv^2�5�N�1���چ���5pv����̼�K�H�����N��Y����ˇ��%ӌ:�'(3�ka�;��O�B���L���:�sV��%��m駱\7i����U�nԛp+�����/K��v�v���ĉ����-�(۔���;.�ԜZ��%�e��Ns��q7+Y�K�Bg����+��*;��v�{��~m�	�un�v.�^H麩	{	����^v�L��}e!X�2�sn�P�ГG��%�bX�>���"X�%�����ӑ,K�����Uyı,O��m9ı,K�ާ��r�V�Y����iȖ%�b}���ӑ,K������Kı;�{�ӑ,K������Kı?}���3XkD�d�fL̻ND�,K��ߦӑ,K��}�ND�T������Kı>�{�iȖ%�b|{���n����e�rf�m9ı,N����Kı>>�m9ı,O����r%�bX����6��bX�'}�rɣ&\�u5��ff��r%�bX�w�6��bX��E {�����ı,O�����Kı;�{�ӑ,Kǿ~�;�����F��j��yn\�V@�1�m�[��p�[c��0�nl�l���ͣ0�0�r%�bX�{=��Kı?}��m9ı,N����Kı>>�m9ı,J������e�j�Y��ND�,K��ߦӐ��FbKE�_�E4��(#� �bn%��{�6��bX�'Ow�6��bX�'ｿM�"+���b~�~�
c()���.�p�!I
HRB�}��iȖ%�b|}�p�r%�bX�{=��Kı?}��m9ı,O}�j��fL��Y�W5�m9ıQlO���ND�,K��ߦӑ,K������Kı>����Kı)�ާ��r�WZ��p��ND�,K��ߦӑ,K������Kı>����Kı>>�m9ħ�G�V������N<���18'+sԖL�;��W&�擂���9m���=��E���MU!�)��sp�!I
HRB�u�pr%�bX�}�p�r%�bX�w�6��bX�'�޻ND�,K��ߩQ5N�7NY4:e���$)!I3{�iȖ%�b|}�p�r%�bX���z�9ı,O�{~�NDı>�}�&9l�)�@�n�|B�����;�ND�,K���]�"X�<'(N��������
�H$ӎʌ����4��KB�����]�+"E�i%��X-H�TcU U"D`Q�`��N�Ď��ٗB�f�YqU�F l��.��@�aR��a.�t��Y�YVV
�L9���@DĄB�b�Q!�VP����fVRh5tJs)� -YpӨ�jD��n.��Z�:��@�||��6U:/ChiDN����;���m9ı,K�{ٴ�Kı/�\U:L��!�Sj�|B�����޻ND�,K��ߦӑ,KĿ}�fӑ,K������Kı'M�69��ӡ
�9�_��$)!~����r%�bX����r%�bX�w�6��bX�'�޻ND�,K�=����c��iքa9�%C �^;qy ��P����;Z��ES��{=2&�WY�2�?D�,K���ͧ"X�%�ӽ��"X�%�������E ~���%���]�"X�%��z��le!�:)���)!I
HZ�{�p��bX�'�޻ND�,K��޻ND�,K��}�ND�,K����\�պ��tj��"X�%�����ӑ,K�����ӑ,KĿ}�fӑ,K�����ӑ,K���v���a�u��L�e�r%�g�Q>�����r%�bX����m9ı,N��m9İ>Q|����=v��bX�'O��Y��Y�fk.K��e�r%�bX�}�p�r%�bX�;�p�r%�bX���z�9ı,O��z�9ı,O���Oj�ae���[�j�:\�3�6�]�y�qbm��-�a3��;��<׵AQ�֊f�Sw�w���oq��{���"X�%�����ӑ,K�����ӑ,K�����ӑ,KĹ�WN��̪���W����$k������uQ,O�����9ı,O{���ӑ,K�����ӑ,KHR�8U�s%9�B&��W����b~�{�iȖ%�bw���"X�%�ӽ��"X�%�����ӑ,K��gi�3YnB�d��e̻ND�,K��ND�,K�{�ND�,K���]�"X�%����]�"X�B��̫�Hm���j�|B��X�;�p�r%�bXG�����?D�,K�����ND�,K��ND�,K� �������w��;����_ٻl5��[�nv�5���fr�H��Ůev��M�2I�&s�=�bt�����;���]�7!�ɍ�����8v�vDun��6��m�����F�sn�l�4B盭�A5�fm�p�<`��J�(��\pV�7J�ru�Z�Y�۳s��1�#�a�����\"{!���nm�׶�;Vx��c8�Iպd�kE��h@C�	n��K�5�h�-rDm��[��
܊��TI��/F�3�
�(�DhwLu�Pj�������bX�'�����r%�bX�����r%�bX�}�p�r%�bX�;�p�|B�����{(�:):�Kct��r%�bX�����r%�bX�}�p�r%�bX�;�p�r%�bX�k�����bX�'ǻ�Y��Y�fk.K��e�r%�bX���iȖ%�bt�}�iȖ%�b}�{��r%�bX�����r%�bX����&2�[���35�ӑ,K�����ӑ,K���{�iȖ%�b~�{�iȖ%�b}�}�p�!I
HRB�㫊��t�UK�Y�ӑ,K���{�iȖ%�b~�{�iȖ%�b}�}�iȖ%�bt�}�iȖ%�b{�+{�]2S&d��k\�.N�M�m�bڸ�mb̘��s�m�2E��ںݗsZ�;�������7���{����v��bX�'�w�6��bX�'N��6��bX�'�޻ND�,Kݝ����23&��.e�r%�bX�}�p�r�(�H*�TӨ������ӑ,K������Kı?{=��Kı=���s�2jL̚���iȖ%�bt�}�iȖ%�b}�{��r%����MD��?��ӑ,K�����m9ı,Jw����r�Y�̗F���r%�bX�k�����bX�'�g�v��bX�'{�p�r%�bX�;�p�r%�bX����y���S%�庸_��$)!{�t�/�X�%����6��bX�'N��6��bX�'�����"X�%����-�r]b�����@6m�tIk�:yvu�m�Q&v�ۇ���7U�u1a�6��bX�'{�p�r%�bX�;�p�r%�bX�k���ʨO�5ı>�����Kı?����d�Xf[��̓35�ӑ,K�����Ӑ� ��j%��kiȖ%�b}����iȖ%�bw���"X�%�~���5��t�UK�M���
HRB�WwU�Ȗ%�b~�{�iȖ?�| r'"k���6��bX�'����N��$)!N��c�)�:�M���%�bX�����r%�bX���iȖ%�bt�}�iȖ%�b}�{��r%�bX���=�d�!s2j�2�]�"X�%����6��bX�N��6��bX�'�޻ND�,K��޻ND�,K�_����S��KI�q�$���oR&��:!���h�溱�g�gU�nD9����VV��=���7���'�{��ӑ,K���{�iȖ%�b~�{�iȖ%�b}�}�iȖ%�bS��<�˖���d�j��"X�%�����ӐlK�����ӑ,K�����ӑ,K�����ӑ,K$/c�G@��J]2��7���������ӑ,K�����ӑ,K�����ӑ,K���{�iȖ%�b|{���n���f���f]�"X�P�N��ߍ�"X�%������Kı/���r%�`|~*�D�����ӑ,K��}��2f[��fY���iȖ%�bt�}�iȖ%�a� �����ͧ�%�b}����iȖ%�b}�}�iȖ%�c�ǿ������^����"�ť�ٷn&�J�ꎞ�ݷk�n��?ӛ����p����Μ���3	��i�%�bX�k���ӑ,K�����ӑ,K�����ӑ,K�����ӑ,KĽ�}̙l�]f�2MfkiȖ%�b~�{�iȖ%�b~�}�iȖ%�bt�}�iȖ%�b~�{�m9ı,Ovv��2a���5u�s.ӑ,K�����ӑ,K�����ӑ,����k���ӑ,K���?��ӑ,K��ٕ}4�E7.��j�|B�����{�ND�,K���kiȖ%�b~�{�iȖ%�b~�}�iȖ%�bS��<�˖���d�j��"X�%��]ﵴ�KİP?{=��Kı?w���Kı:w���K�RB�
"�$���W�J��`�m��t���f��U盰��5g�p����5l5,Uy�!j9ձ�]���pTh�t�j�z��X� �:�	?��>O���8sjp� 7Ag�hw�w!����<ݴvnJ�ݺ�#�@���m��3�..�5md#j�͊�e1-C
m�E��Vvӭ���\XƸE��cC��l�����%�l\�-��yM�T�H� w���3SZ��#I%p��Q�c���T�q43{z�N�Z�/=q���6�E;^�9�l�-?}߻�bX�'����.ӑ,K�����ӑ,K�����ӑ,K������r*HRB�Gm򚂩Ԧ�Ӧ��|B�,K�{�NE�,K�{�ND�,K���kiȖ%�b~�{�j��$)!I3{�)�cd�T܍�j��Kı:w���Kı?k�����bX�'�g�v��bX�'���7����$,㯊l�әc��M�ND�,K���kiȖ%�b~�{�iȖ%�b~�}�iȖ%���ӽ��"X�%�~��ײe�Yu���e��ӑ,K�����ӑ,K�����ӑ,K�����ӑ,K������r%�bX��K;I�d�Jk2^�çU�C���ɖ��U-pӭ�U��FZ͌�Yo�9:��)~�~'��u���{�ND�,K�{�ND�,K���kb"X�%����]�"X�B�f̫�)�PSsUM�W���%�ӽ��!�����K�{��ND�,K���]�"X�%�����"X�%�N���r�ܺ��.��iȖ%�b~�}ͧ"X�%����]�"X��%�����"X�%�ӽ��"X�%����'���MY���Zͧ"X�
D����iȖ%�b}�p�r%�bX�;�p�r%�bX������Kı>~����Y�fjjfd�e�r%�bX�}�p�r%�bX�;�p�r%�bX������Kı?{=��Kı=���L�kpN��5�P�[�떖XM��a.!���\i^X-U^��{���>���[�w���Kı:w���Kı?}�siȖ%�b~�{�a� �$����&�,�өt�Rs@�)�j(DN~�q7�,K��޻ND�,K��ND�,K�{�N@ıRB��s�NiЉr�w����b~�{�iȖ%�b}�}�iȖ?�ة�m�' �,O�<{���Kı/��iȖ%�$.�e_cLR�*i�nn�)!I�����"X�%�ӽ��"X�%�}�fӑ,KlO��z�9ı,N����5�MY�5��a��Kı:w���Kı/���r%�bX�����r%�bX�}�p�r%�oq��������[��6-��Qy�].�I)'D�9���6�.�{e\�c��ԝq��.�fK����r%�bX����m9ı,O��z�9ı,O��m9ı,N��m9ı,O�gi<��#�:t:n�|B�����}�p�Kı>����Kı:w���Kı/���r%�bX�?gd蚩r�e�����
HRB�f��iȖ%�bt�}�iȖ%�b_�{ٴ�Kı?{=��Kı>��)���պ�Թ�Xm9ı�����ӑ,KĿ���iȖ%�b~�{�iȖ%��"�������}��p�!I
HRB�����:uT��6��6��bX�%����ND�,K��޻ND�,K��ND�,K�{�ND�,K�kW���̶L�"�	��g t���Nn(Ѹ��펶n-��-�h3�ӊ�����7���{���z�9ı,O��m9ı,N��lG�,KĿ���iȖ%�b{]���	���ɫ��˴�Kı>����Kı:w���Kı/���r%�bX�����r%�bX��m7�k�&�.kY��iȖ%�bt�}�iȖ%�b_�{ٴ�Kı?{=��Kı>����Kı)���.\�[3S3%�WXm9ı,K��{6��bX�'�g�v��bX�'�w�6��bX�'N��6��HRB��죠t�1ӡ�w�ı,O��z�9ı,O��m9ı,N��m9ı,K��{6��bX�'N��H�#`@�U�|��£7>�ݤB�iX`XQ�RQ�X�R��@`�#�p����ߔ�u�6�5�.�:�!©�4 <1e+4J�0q�R�-�a*�i�H�+4�P��j[�)(A2��4i�"�!Q�@���H��4%�ZQH�yEpWY�`J���;��������      �6�    ۲	rR[5�[[ff�Ѓ=��p�m�"��j��6q�b�
��A�T� *z���m�f��m[�HH�6��'m�{4��/DI�WE��l�ڥ�S۴]0'Z��i��.�eڎ9�`��+Ͷ���V����$bێi��4��ZeV�Vΰ�e�Y@j���g�j�v�m�Z��8���68�s�	��U��8N$إ����VV�����6ݎ$���^�cW�b6���z�uO.ݐ���p�j���j�+Nʤ��-\��-��U��V�,�W��)r���t���r p�-C�ɕ 689���Ю�\��n�9�(��d���ئ��m��p���%��ܲ����-g�Z�U���A�K˫vV�n�F�����S�5����7}�I\��GkKmm˖u�� tn�V�ۗ-�xbS61FԷTc[l�ի��:杉8Ʒdj���1��(z�XsS�^\F���q���J�n��T���Uo7��^r�vq�d�TBz�0U��^4�7kvۤA ��4�z�n¦x���g���U�*��[7Oc��b�FYUZUB�Է����63�.��-�@�ϝ����gv8B�� M��� ��N�Wp��}խi	��5�v�Շ��	M��mpB��ݸI#Y���j[>�cm\u�n���ۯ5WO�{g[�f!�m\_:ٕ��.k6���퇮]Plۮ��(�o�KM�%e��덄�IRz�:8t�7mv��/etҪ�c1׮*�g�eP�Ƀ�+�${rr�EL�VI�CcBv.��5A=��Q��M��#�q��	�
{��ٔ;iXۊƛ	�f���#tۑ�tt���v�8I�Z��}�>�,�IgB=%���gd����r�ڴ�t��k 6ͻH m�@�6T�δ��
W�窕j��Vy8;S��:�yƑ�Z�3j�aJk�ԕ�Ǒ]��n�N؀y9
��}�{�{����*����>Uz*#��	x .<DjUC�W�U4�Wf�kXffffafa����8'���D���S��3��w5-�w[�x8��1y�����^cs��]m���vV�����0�c'gm��:으;tlf��޺)���Aqv�*Wj9�'7`��7�~0�/!�A�<[d`��ޘ���v��S��h<f�$F�2<�nٔ:���Wl:拎�c�M�d���.����SH�b��ɹӧ���!��5�f����3F]�&����qr�n���bHi�:�JET�,ٴ�9���wy��qT���QM�77�RB���g���r%�bX�;�p�r%�bX����m9ı,O��z�9ı,O���x�33WV�3R�]a��Kı:w���?�#���b_����ND�,K�����ND�,K��ND�B��������qN��',E6��,KĿw��6��bX�'�g�v��c��,5Q;�p�r%�bX�=��ND�,K�}�k^2SYu���\�ͧ"X�%����]�"X�%�����"X�%�ӽ��"X�!b_�{ٴ�Kı=���^�S��ɫ��˴�Kı>����Kİ�#����m?D�,K�����r%�bX�����r%�bX��zI����ع�x!��t
.�ML�� u&t��E=��:�5:of�=�%���̖%�bt�}�iȖ%�b_�{ٴ�Kı?{=��Kı>������oq���}��u�L�k���D�,K���ͧ!�l8(b��cȚ�bk����ND�,K�w��ӑ,K������O�uSQRB�}(��E)tʧC���)!I���o�m9ı,O��m9ı,O���ND�,K���ͧ"X�B�F=���Sl���2�|B��� �'{���ӑ,K�����ND�,K���ͧ"X�%���ߦӑ$�$)!fu�\�6�je�E74����ı,O���ND�,K���ͧ"X�%���ߦӑ,K�����'���{������6]�`Z�j��z�^�� �ؙV��+mx=�k��[l6ˆ��K�S��W����$)��;��,K���o�iȖ%�b}���ב,K������Kı)߽
�L�NiЉj[n�|B�������ӑ,K�����"X�%�����iȖ%�b_���iȖ%�b{��_cLR�*hn�p�!I
HRB����Kı>>��m9��b�~�e���?�?D����ӑ,K���ߦӑ,K���S��a�D�e�s0�r%�g��5���ND�,K�����r%�bX�����r%�bX�w���Kı/����\���,�fMZ�iȖ%�b_���iȖ%�a������i�%�bX����m9ı,N��m9ı,K��}���u=��v�m�c"\:R0�;��S��3��ɛ��5ն�|G�����Z�L�fӑ,K�����ӑ,K�����"X�%�ӽ��"X�%�w�ͧ"X�%���v�:֦S3&�s5�˴�Kı>�}�i� D�Kǽ��iȖ%�b_����ND�,K��޻ND�,Kｲ�2L��չ�����6��bX�'N��6��bX�%��{6��bؖ'�g�v��bX�'��m9ı,O�=�Mkf�]LֲL5��iȖ%��D����ͧ"X�%���]�"X�%��{�ND�,�C?�G_�x|:�'񙾛ND�,K��v��ˬ�%��fm9ı,O��z�9�I
H�������V�Z�os�7*g�϶�g7$"v���Up,a";)�2��l�N�8-�����MqYL�09wF��L`z\���6�[��e752�V,͵���C���uwM��͵��x��NFKd�)�R��������f��	L��Z�.[���?,/�8�#p�294K���`r�0t��߶���l�$�jF�Z}빠e�~�p���{^��q	F,��:UT�m��Y"]2��Cv�j�b��h�t��l=�N�K���6��z�@��-$�b��N^���ݫQ�af�=s��X���p��)�P2���V�&��z�ƭ�����I^��7@������n�y�ߟ>|�/\a�Ye��xz�"rq�d��t3�F۷n\۳�Fx+�I�����ծӳ���A�;Le�8�!���̶[->j)�E�Y�7�J\b��+���3�� �]vS=����;�[�����!�ӫ��:2���]h�#;�?/�ߚ`�1��rS{�L��7?8�L���ܙ���Ď���h'���Lv�]Ņ+ʼ���3�%07�4���`�1�3&V�
����T�r����V,͵`�k���>�3w�U�)�P6˪�����`�1��rS�#L��}�~�D�KBP�`eV�iE(��TI��.�{�1�`"4Z��b.�0�Wx��L`z\������z�h����#��7	#jI�r�V�DB�[��ٽ��V.�֬��v�u��l�$�jF�Z;n�����w��@�v��� IiI�����E'�&�?c���F���n~j(��1�3@;�Y�rܔ�����ti�5]P��ς�df�n�a/�뤧�:,Ht.��=4�<[T���q�1�dX⑘F
I�r�V���mX�6�����~v����S-1U�W�Y������ti�n��+�h��Y���A�$"RL�=��ٹ$������ H	��(uM����^���oW�6��j�f��-�:d�SMX~���v�����۶�g�w4y�a�����ɠr�)��Ѧ.�� �I�������17#�� 6���E&�u��z&�ҩ��P��󒽟������a)h��t��`r�0t����)��2�(E"M)##��{=빠��@�v�����;K(���Q�7crc �I�K���ꮓ�L���0ݦ;�R3�$�k�h��恋7mX"I>��J-(��@���piL�' 7"qh���.���.J`/��/��~?X�PcgVz�Mqk��+qq��Wjp��E��3mn�	v�4gl���{�}����97@eVf-����� �I��%07�4�3ޫ* �$��� 筚˒��`r�`yu�"|e�]T��n�������VrJgV�Z�߾�?u��n%"i5#r-������4�=�ce�Lٔ��&)$#��{=n�s���ڶI�ﻳrO�*� �@#���Ԅ�Om�{=[�����8+��b��l��ݪnT������r�ײF���������Id�qs�.�l]\�k�u�8U��:7bMэԥ3�������;N�ly�I�jt�����i��"zj�(�ۊ�f�����j���@k���K ����s�"2��i@��Z�h-n���6_>3wl��VP���.�h��Ԅ��3Z�K�]�y���w^����~w�?3w(�YYӫ"��ru��8�FV����ݱ�u�"f��S�s|�s�D��	�I���>�&���Z{�L]#Lv�\�e+�̱ef7`{kvo�L��֬[�j�>���&OgJ�EL�NS�M�9�3w�X�F��L`l�)��K����ah��*�109t�0t���rS���}����"
A�ALm��z�`~J3�t�n��nڰ�7B�O�\c=$���]Da��de�MZ���rm��k�w=p� ۲�k�a�KQM~��{w�`j�ŀ{�����˙�V�f]f]�?}�vo�+�(I(��|�!$3o�Xnk�=��7�Də�C���3D��LtՁ�{�0t���rS{�L��]��YQ�7c�f�s���ڴ��s@�z�� �v��2,qH�#�h��6DD%����[�j�>��`���ހ٬s;�[s8�c�M��-�c\yT��N��dó�lj����.#��[*��`r�`�1�����f�Ù���I3@�z�� �v��f��fھI(���Ҝ��d�Cljf��os�=��6}�%L(�hiYa�a !�C�đ�@����An���䅚#H���@Ł���!!"Ĉ@�#� ��BAH�X�1`�$B �P#X�P�"B5!RH��XU��`T�XD#@�H!#Whh��VT!a%� Սbb2�!a����!R�H��f���!�h���ÈNA�1b@!t�j����{T�%HkU
Q�D�Ӧ��~O�	�F�@�!(Ƒc(� ���Q���X �~MbXA�"��AX��bh�S��4+�hS�j1bE�� �A�����k� ~��YH~��Ὠ�s�b	�D��W�W���h�"8��!U���b�A�"D�	��PF�P Қ ,DJ>IDC��]�V�ڰ>YY(�:�]K��В���>�3w�X��� 筚?u��n5"iD�Z�6Ձ�!j�����`{kvl�}�v�<C=Iqu�'l��u̗M�6��YI�cvM;m/����ٽ*�x��F��L`l�)��Ѧie���6F�LrL�z٠v��`{7mX�v��Q�B���U��ʧ.\�m�W��`{7mX�vՀw�� �j�@jb��qŠw۶�Y�j�=����BI	@��@�T�<�}���I�}�Sx�a�Hm�f�V,ݵ`~I)���]�`w��h�J$��LJF�d�'g��\㲅�M1[v�ۧ9�[r�[s�\����j���H!�HLI���٠v�V��[��{=n������#��5	�K�[�}
d��`j��V��w�DBQ2z2�N��uM�L���s`f�Z�9t�0�1������efUYY���Y��ˤi�oI��%0���*��������W�r�Tr�`�ce�L�`r�`/����m��ww`�m��h��$��u*�N�"�IW���X�5t9�P�$m�����7h�Qr%�m�Rj9�5۷\c����;Wl��z�i3�l��j�[�"�<���WJf��\n4t�҃VvNt��� �I�-�i���@�2	�e�׮[tWc-����v�ě�Ǟ��A�Y�㶝�ÃuX���R�1���̘��[UU�g:""��κ�������������w�[����O�`5A�똹df�Y�m�鎰sѼ�\`#���딀����b����!����=�_�6�vՁ�7mX�l�9ڲP���$�N-��s�)�V�Z�3k�lmń��R��M2��T�6�Y�j��V�����s��l��V񙲜������i��rSe�L�a�QO߼��Շ߈�dl��G���Z}n恋7mX�ݛ �ɭjF�[��;�u�c�NB�f�W\q	��f:��k$X]rˋ��"����rG$�ȴ�����w4�ڴ�j�;�;�)b�dֲ��|}����@�Q:�A�Q(I-P���~�zl���f��;�~���F�pȤ��~�@�rS�Ѧ.�� �xW0YJ��.��)�����L]#Lm�� �j�@��I (�@�}w4�\�}���-�ڴ����3f�Ks����KNf2c�{=53�7	���8i�a픅c��W�u���U�6������rSe�L�0ҖQ��Dd�����s�ՠv�V��z�1f��2yml��t�T1��9�'�׽w$���ٹ��Q�����%Us�}͛�{���rN���,֤Q�$�ȴ��s@�z���v��ڴ����D���$��yf��^��?�]�`{3mX�)���:��@��a�� ������7k��sŬq`���My,��	&�7E���)��$��F��F�����!��5�@궽����1f��پS!��\әsR�6�Vf^[����H��rS�rS�ֳg�̃	 Ғf�����>��I���n��N �V�D���C� ~�y��Oӿv�\��#T�)L�V�[�`~K���O���֬Y�j�=�b)N�n��m���v63dV@�0ܫ�ݫ�,\0�F�R9�^m�n�I`��~#���IZ;e4��s@�w�s@睫@�A��R)#�U�����V�i��)���L���+��s4K�:cmX�zՁ�V���(S>�|X�֬��J���3�LȤ��v����}빡Ӌ7�V �8U\�*���]K����� ���%�~���~i��)��-����������V��݂�;sA�b��qm3\i�J�ά/B�w*]Ej�\1��il����N�Y�t�N��;-��@�Vێջ-�Dmț�SKz��c{�IӺ�`��m�NJV�~q�|�#�׶ϗu�m֨���p���`����H�k 1��u��N����J�N֎�Y�����ZЌ�G�-�L�ً/�vM�t���<rb�b[�lg������{��� +��-��2~�3&���Mg'C�`N׶�d�l�r��x��-���F�,t�,���I�t����w;빠}��?�}!��Ł��T��M2��T�f&����rS�2�?���$�U�b�H(�$�������=� �䪺O�09t��˯��/.̻0����`{fA��Ѧ����v��0~E�ㄑƉ"p�;�[V�Q�7�_��>��,{l�p��.	��9��<Y�c-�.{7%��wH�pa��l��Wm2t�Ʋ��J��ؘ��Lu�L	�%|��z��������J4��)�I�<�Z���DD���@
�R4FA�B��$�/�3���3smX��j�3ݦ7rD�(�r-�ڴ�m�?(��[�j���t���Z��sS��3�2��`E�4��\�������Z�l�9�a$RL�=��i��)����F���-yv$rZ��m��	�Vp%U't�W7]��e�����<��8���/-��/��`N�)��Ѧ]#L/?,/�8�!$�Š_;V��z�h=n��;V�Θ?"�q�I#	�4���fڰ5f�%y/�	(�� Px"H���_	���u��@����w� �ȤI�9�^&]#Lu�L	�%0�_WI�Ɂ����j%RLȤ��v���L�0"�`MWT)r�ॅef���q�ٜ�0tj�0�q!�={L^�n���٣��{���n_�c��X�h��~�����`E�4��\��7`�T�M�-ӛٛj�)���Z�=_�-�ڴ[Z͟�2$�JI��ݵ`}��6tD)���7zՀ���r�ɚ�32kF��7'�P?�X����l�_�M��͵a_�BB�I(�J9(�wZ�1md��t�T1��9`N�)��Ѧ]#Lu�Ll�o�k���܉��p�����I!���/��6�u�9y���zv��X�d�]�����.������/�Kl?�_���-��?��H�lL�f�s��o�=��6mwM��͵|�B�3��z�IDI0S"�4���@�v��Ѧ]#Ln�]Ņ+�1aYu��l?BJ���6f��Vnڰ�
'����=�+�1�K��a2�9�=��V�����f��fM���%	D+�� ���ʠ ��� ��AW�T_�U�U�UE��Q�E�$Q(�T 	E��Q(�B�DX"�b�A`�DX*$!E��T �0DX��Eb � E���`�0DX Q"E�E�,QE�DX�$QAb�DXD(DX�DX(B 1DX�A`�@*Eb�E�1B �DXT"$"�P���bA`D�aT! T AdAP�QH
��*���*�� ��AU��
�W��_�U�AU��AW�A_�PU(*������)�����C&,�4( ���0���         �        �   }  R�(QT�!DU(H ((P(�
@ 
UR�( �  P ��  @ 
�8  1@(
�$ +l(�i ��������� ����mv�qn}�{������h�� ν���Ҟs:�  ������x�� =)��m=��mnnU�o/N���=nf��5N����y�]� |� B�  P�
'��q|�.-�NM*�4���P�|�&��_N��j�o�_8�t����qܾ�}�Jr ��  m�C4�`� `�}�ۻ�ٵ�7,���|PB�    ͂�=��\O���6��\�����y�B����7N�-�Nv德�xW�Hn�����rk� ��ە{���ϼ
�z���yO-Ů;�_[�ut�x �;��{={j�n�n�����7�ԫ��=T�  UT�� �ն��}�����c�N��۔�����d�,}��g�QX���	�JVOsS����m>[ͭŔ�}�<L��NO�^�Y=��������}����n��w�u���kٜ����yJ�TU**EP� ��){���w�}�s>OK��� �Y��   "   9�� � �    � A@ �6 � X �J�!� c( D � 
D    ����T�   ����U&�0@'�UJ��%LB'�T�IUC#����Oj�*� �M�)T�HlM�	�g����?�?�FfnZ�����������IWAg�b*
��DQT������������*
�ES����Ժ.��Z������~�_�����ʑ`� ��q6#���"i$��]`jc�R�-N*�v��iI
h�vo3fnhՄ�p�ѷlHbFĐ����n"��T�!�C�a��f��Eđ�p(��$�`VH�"K�����$����\��y$!��i���V$d�V,6�Ȍ $Ad]�+$�I!��&�[#�D��3DK$hj@ѓ|%5�i��n���:��#I#a5`����PП������au���n>�DBJ�X�p�5~����I��P����+5я�>5�Vo�$�|j����HV@%]?k��2�
h�݁��D>V���0�GLY�����k�����>4艤0/)��']	�Hk�e)�2o��C�Mf�?s_~ύ�Z�SY5����$+����s�!G��f����.0�,���$b�taHҐ�Ж�����M���,F M$`�i$�D�i�˭M�~���9�rkN�k��ܿsY
~aaq���ٯ��
~��kY���|�� E>X	0��HB�!$8J"J��/!�#�8D�QИ�d8�P�0 �<�4��p`R4�5"l��,F7ND�
B�]3�S�@��Gc��E�Ji���c�!���n?���S��Ji"��T�5tA����.�XSa�Zblɚ鐺�w\��u�e���ZjB��d�	�ӈqaM)))�@ػ0fkfJh`U��l6ĊĈ[����C5��)3P&�.h��2�0!T�c����K�2o`��%5���4�����bB��AF  S�>WN"=�[J@��8���f�%	+���Wi��,Ն0+���MI�J�0v$����+�H���2G6RBIMol*��c+���$ HP#aI�i�T�DO�٬�r�oA�h��CFi��H@�A���I������#lu�&��H�4͙m�k���l��V9��,�(d��h��U�I`��u!���B������� ВZu`GY�BF%����C!\N������&R�4��W�tF�;BFn	X�R!A�1�l�$RM8n4B�?#�4Z��%�8a�!��"V�a��6F�$!$��PіX�#
!�`�J.�$�Mc,� �$�L�����IcHE5$Z2E(HF�!	�C.�~��ԉu�g6m?F#K$A&f�6��ZT�H&В�0֩�o�7� ; Dd �H���%BF�BB$���ei$	m��I s��$��𐀜d!�@�B��H4c���F�B0$B�!FH�4~@����T�a���rc��O�@��	���~��Bb~��� ,#CI!"A��C$�:��a ̥ �2@��1[	+��������H�	!���j� 6�p�k.���X#C��mB5юؤ#CI���A+!��"����X��Q0-�ta"F�HF�X&�Cђl"B�0܏p$ɣ7�8V$k��$�5�N�+���|�6CK����H�4f�Cc�6k/���npk]\���Y7Nr��_�u������q��%a␪�W�\�!�$ԖC�v<vȐl&�n;(#M���H�$ �4�l��,#t�!tŉ��ma#CKCCi�1��ťt���� :�����s���9���\
�r�g��N$T�jD	�Y�e��[�!t�Ɖ�#!E�A
��qH$BD�a��!�k��!�?&�8��|���G�l��D �R��~	�1��v�'#�dh����D����bSFǀ@��k�����"PÒ��r�9Cf��Ӵ��p#d[BXj��D��~�����
���^o�ѽ��n������s���]8l�F����/�Z�Ѡ벑�`���QީÄ�,�p�su0ĊEH�`5��Ms�ă]8�< �@
���RS6�˼6Ja�c]8�	�L&m?l��l
 B�t`K�YM&1��v�l�͒�l�	
�sd�<d5)�hi�C)��E�b.�y��o	d��l"���b(� �i D"��F�B�D���!c#@�B4XT�`PM&B��Ml��$$��H�"�I!C$HŅ)���9
L6mH4ю�$i ���$
p&����|$�dK&V�Y�O�N�]I��K�5B�1x���a>�����9"�3h��~�il��"�
�A�Cm8S���`l�CH� ����0H(��A�	��Ѱ�l5ӵ�&�%tὐ���@�f��x�Z�H�"�04�jh��p�@٠�D�w6nP�,�&�����4�d
��!�-��aD��*9M酐7��B�n�8�#����F%]0)��L"kS0��Q#`��d�]dij��3�!�!#2Y�3D�[�Z�\�|�����H� �TM��)��';�����u �48�ĊQb�@ �`�5�W�F[�>����j��P" Pb�36��|h��!O�7�;6����� � �AHAR��F�ԃT�T`���@� �b�FH`�BKH"GBAJb�J@B"D"����E��0 h�$a!�]1�8I+�&.��	�@�Z�d���L
���h���²щ"DcbD"BH- �eR!L)���(S���0(� q�w
hH��ɚ��4�� "R4"�X�����$4��D(djŋ�q�R�6�X%4`GlB+ ����	H�`p��c����,����q#FR�`B�7�dY���s|+ā�ԃ1w$���5�]��?_�7������D� ��#X�@��EB�Bi dV�#�]6��B��)$��^��WH���&��*�o�!���l"
p
qbH�<LFf�f,�`�b���#m�$�@   ?�>                                                                      -�$                 ���                                                            ��         q�l���T\�J��K�6����6��kX �$�� m�i6�l    [@_Z�m� �c�l �-�K#m�pBڶ��`
P �m����  ඀  H m  ���[m��p�m� ��m� �:}��lp �t� k�U��[A��uhl�m Hm��S0l9�ڑ%�ܶ������&�pt`kX[@�H�      �|�    9��l  6ӛMRh@v� m�h�V��pT��UUmT� ��ݲC��� �@
ZtP�UJ�:m�m%� ��V�,ݫ��p    8����UUE�Wh� m��D���$����i[�H 6� N�/-Ѭ�Mֲ�:�@t�r��٪M� ��ym��l�v�i $��5�.2h�\ p�ղf� m[^miD�D�[��� � ���Hrʀ��ک
V�At �@	]�o[N�H [@�i  	 A��v��m6����ͤ�ګa��n�YЄ�v0�@-�Tp+v�ܰ��  8�� E�am�-`5^����v�[o�@q���)mJ���J�7UWM��oV���my��n&ʪ��Z^Z��:�ƒ�V��-� ���:@� Zl�pjU�,�薪�e�.�-�mշm��um�   �mץP5� V|���MrUW@��7k�Ͳۖ�&�r۸    m����]Ŷ0&�A�����U��*�*�|�UUW�/�	��VT�Y�,���L�D�*�A6
���@ OE����zT�4 �,F��m3��K,dvw�j����i<L�HN�KӖ8Z�@]$�m���  -���oQm �f۶�K
�V���(6�j����@�-'�c�Z-����ئlKuT�l��E���)!�l�m9J-�"�E�m�kXm 6Qy٣`��H ��1�Vu� 6�0,0mm�݁��� ��a�m�R����l�m���m�� �l�a�m[ m��-�Y�m�#m�[%���֑�ʮ�V�"T.���J���kkE�mTJ�*�W Ҡڴ��rI۵��($pp �b���"B9��U(�9]SU�j���j�1R��UUr��2�6��e�k��%a�=�
��%UZk)�P ӡ�TR��*���U�YKj@᢬,����E�k��$G�� !v�8'l��- A��  m���`�k�7@M�5��[@�%9ui�Hڤ�CmA���*UΉS3N��Q&��@�[l�U��C|   H m�[@     �t�� 6��  v� ��Wm� ��*몋, r� H     ���HH  0[B�[I� �I>�|��rl�Yb��\v��o��\Yol[�$��Q#m��6��k�8ݤ�ʹk��m�I�z�y�f�� ��a�� +j�uԓ[�  v����:N��[d��MT�t�ۖ�_,�5R�����R���� ͖��K)�u�k� k��-� 6z�u�m��l�R�����]����,�sj9�m8[v�v��m&� ;n�c���Tp:*���n1��B:M�`�])i'ZlH�m�o`mj�n�[Nmm	�m�h����� m�7l -0 %'��j�SR��vWi�l�f  m�h�a�m��$Ͷݴ�z��X|  m��6�0k5��$�� �,���������}����  [��-�-�հ m��j@M���ay��W����_���� 	� ���m���kn��6�$浍�h� �� �m��  � m�@m��  $�8 �c�� -�&ٶ���ݣ����^�F @�  ��$ l86ٶ۶�m�H�i5��   [��J�6�"@  � X֜6ؐ8R��4P �im6�M��nX[s��	�v� 	 �m�V�m  [D�mm�m"(�a�m�ۃ@�]������ـ�ۀ���\����5�ku� �t�`$[@����h TdYWmګ��Uej�U�i�m���l�`�g�k��U�I�j���#N�I妷69!����yU���m�9W4�V[Bޠ-\��\-� �rKh��fہ�� -mҭ���5R�iy溕�]`
��"8U涺��eUSSTY�T�ͦ�Y*)�;5[����my���ۚM�v��ve�UQ��Eù�&ƶ�#Pʳi1U[FknT�l�j���m����ru.��  ���|pm�m�����k�!
]�S';h5���-�m ڽhm��Az�B�'A j^kh �`�$[%7m�J�T����i��� �� [@ ְ�l�l���Sl��Á#m��I� 6�m"��m���ݐ[4��K@6� � 8�>�l�+�A�ll�c�k[j�,�l �{Y.k��`,�`��"@6�   m��6�lěb��J�����N\B��m��ڵ�m� 6��Z�� &ٷ �  ��[Z� m�E�ŲP6�Z� ���v��n$N�඀���6�   ޜ0 �jۀ�[.[@0��S[�i�&�n�m��p   l �d��	,�� p�nnScZ�� � �Ҷ�5��-�    �cm� I�[s  ��h7m��Y�p�H��Z+j��� 6�@  h��ڶp�ͳl 6�`Kl�.��[J�	6�#tv�o�_�� ��ڐ	     �m�P�)��U<�q�<1v�����`�  	 i��m� m     6� l       �`Hְ!m   ��v㶝-�v����  ��m�?��  -�       �h hl�-�^�  H$�[�-��T U@*�F��1U� UU) *��l�嬖�I�m �dq*��ڶHkX  �i�"0��U*��V��Z�g;Y+ � �  ��;J�vؑ��m5  ��@R����    �b@     V�l	kV���m��p�8j�@[V�-� $m�"��ۖ���dM0m %���d�  9J$ ���m� �`�� �]��l"�=��  m�  @pp$:ޡmAm�m � [\  ���a��H�  m�X�h-�Mm�[�     �   �p8m$�m6["�m��6��$rCm�-�       [@ k5  h 6��^�p���le��H ��   �c�Ͷڷ\;d�j�������RZ����ـ�UBl��C ��  p  -��m��}����n��Mf� �  ���m"���m��ڋ�A�[VBJ�6�A��$Ht�l�i �CI9mm�z�pH �ZVo �m[�ܻ-@��1�����s��f�V}��X����+s�9��D:�J]hI�뷃��Q҅�$��h�tu��{^�Ӳ��[^����{�\�v�������[��#���ʪ��ݞu��
t���5p
��W�]h��[�H�m�e؉*���]XV�8Z��v��%�Ā,0�ӭ� �>5�Ll����հ   &� 
�� �\��*�A[   [@ -�m0qR�-R�;s�]�;` ������ v�m� 6�`  i6�R���8ڶ��I����v�v� ��x6Ƞ��    6���֛$ݛ`�m���٩��nffff[���(�*�DP� �8���
�#�� �Q0
AE�.E�DA�W���E� ` yUP�b`�X���E��Y"��h(R
�R1�HQT҆�D��AC�Oʅ 
~P�('Ȼ��������E����4�� t*~@���Gm A* +�~>D>p@� �AG𮄐F� �,�$QB���(��E@#�P�P �v��\���Q1�� Ѐ@� �ED`� ^��:TGj~>�f�E>?"~Q9,{�M��Pꠎ��@D���Q(���@�C��WBH��~�(�� 8����W�P����X�"�F	�{�ֵ߯��    ��        ��`  kX           l lKYt˒�u�U@-ڙv�2K��ͩ���{�������9u�ĽZ��#Fg�;t�	8JFL7k1�X�B��m��&�Q]^�ew`��by�Ͷ�vB��
&�y�9���w!�ӱ�L�M*�ք9��Wicf���S�rPj�m�i��P%Vݴ���g8v�j�V��۱JU;cF"�aKD,WII.�\��Z�<vR���,A(��8��k�KR�UgJ�V�iW�ʓ�u=V�I�஭.�Ɂ������W']���HPu�K�s�հ�B��!������v��j�{8�l�$9����M"�
�C:ܺD��۫���� SfٹQ�����J]<��̼e��s
�h�:(���j1t1rb�[��2L���jmJݕ]�����a(��g=i��k4�N\d�0g�I�7fV�aS��7d7]�;K8%��v�qے{!;�#��c�n�fwAb��j���6FKm��h��K�	��m���38��F�N̮ґ�wM�Ʀ��	K���nI`Bvd"7McJ���� ��!�W�Y�Õ8���xl;l�Z��θ�r0[U�M��g�mS.�ϗ��;��l.]��	������b����ɴ셛$�P�C�Ҧ��ip��i9h��V���[l �6z��HBڸ�<�!�"c4Qm%�'Q��.1*�Vt���ݘv��w�����xk� �T�B
��1u�R���V�j���q�*�Wf �^Dݮ�*�/;�୐�[�
�V�k�ԫYW�s�In�@�'meݮӍ��k��id-��F�垵΄� ��e3�Ų�B��v:Z���ӰXH�yRڛ-��m%ٞIڰ�5	&������=�*�� �/���ECH�s��{��w����w}��~�� LҭUUUJc���	�ml�n��i��͖�J�ўzbW����/3�	�c��f�v��+�[��]�e�&�,I�ӚRY�MEXT��n^�fY�2�5;6ݝNɭ(C�P,[]u�
z�t��ڞ�1�*q���n�i�U��[�R=�]��sB^wc7[�6��>�E�Oh��#jeS�����z���$�8�H$�lk{�׻����������l����� ��{lsۀv�Dܝ��r�=���tJ[�F����o �w�̂H$��~�pI�����J�5ı?}�siȖ%�b��=��V�35�-��fD�Kı/?}��r@� &�j%��nzT�Kı?}�siȖ%�b_�w2&�X�%�xl�:	��UUr�誻�_��$)!=�D�Kı9���iȖ%�b_�k�Sq,Kļ��siȖ%�`��}��.���u��Z�&�X�%���w�ND�,K���D�Kı/?}��r%�b"b~��eMı,K�������P��q+}��oq���/ﻙq,KĿ��siȖ%�b~��eMı,K���6��bX�=�n����pWj.��5�K:��3���%���k� ���P�:.�ɩ��u�q,KĿ��siȖ%�b~��eMı,K���6��bX�%���T�Kı>���W�ՙp�kR�k3iȖ%�b~���p�Q?+�TL��,M}��m9ı,K߻�q,KĿ��siȖ%�`����%0�&�j�k%Mı,K���fӑ,KĿ��dMı,K���ͧ"X�%�߻��7ı,K�ߺa0�%�Y5�-̛ND�,K���D�Kı/���r%�bX���l���%�b~����r%�b��?޿ P�S&4���oq���/���r%�bX�����ț�bX�'﻾ͧ"X�%�~���7�G�#�=��ͷAd��q��l��ml��f
���Ų�/JA�5�]��upֵ��kZ�ͧ"X�%����ț�bX�'﻾ͧ"X�%�~���7ı,K���6��bX��w2˩��.]k%ְ���%�b~����r%�bX�ﻙq,KĿ��siȖ%�b~�u�&�*�bX��_��R��`����7���{��?���n%�bX����m9�*pA� `� �@`���:2&�}��dMı,K���ͧ"X�!�������Eў�h�ﷸ��x�/���r%�bX���l���%�b~����r%�bX�ﻙq,K���7�Z�.᫫dֳ6��bX�'��["n%�bX����6��bX�%���D�Kı/���r%�g����wv��ϿeXxGkM�P�6��j���qqc-�=�ȋu4u��V�����{��YrS�h֮\�'"X�%��}�M�"X�%�~���7ı,K���6��bX�'��["n%�bX��w$�Mᬚі�M�"X�%�~���7ı,K���6��bX�'��["n%�bX����6��bX�/�MR�f�f�wWAuWd,!I
HRB�ky��Kı?w��q, �,O�w}�ND�,K��s"n%�bX���tոkYL�kY���Kı?w��q,K���wٴ�Kı/�w2&�X���(�| ��<ȟ��s6��bX��'u��j�K�Y�ְ���%�b~����Kı/�w2&�X�%�}��ӑ,K����dMı,K�~��j��pYēd]iQ<���Nu뎕��d��m�Mk�>��wwr�����.kXm?D�,K��̉��%�b_�w���Kı?w�����D�K�����"X�%�~�{W.f����u�q,KĿ��siȖ%�b~�u�&�X�%�����ӑ,KĿ}�ț�bX�'�}�R�֬���j�Y�fm9ı,O��D�Kı?}���r%�bX�k��n%�bX����m9ı,�^�����֮\�&�X�
�b~����Kı>���D�Kı/���r%�bX���l���%�o�~�HL
c�dI��9u�@>�f����o�Qq�$D
!V];��@ $   $���f,��0���v|��ݬ����j�n�҅�`}w.�)�/mlfy�b���cnqg��n�u���d�[&갧i��F$ѧZ�]6@�#���BL�s�)��6:u��^\���֟ԥN��#���!��}�q�}ɛ��mt`p�A�qM������L\�+jxΎ�Epn�1�l^']��l��Egx�Bl!7��awɻiqkm�4L3�m��FT�eͮ6n��G�rA�&ҘH�"n?�>��M�n��־I~��/�&J��}�������Wt��� �o~P�d�݋ r��@=�Y�yP�`7�LX�rbnf���F�n�Iy��kL�t�#i�0����˭z�u���X�!%����۳UT�nm\�T�q����/0=mi�=+L	��a�?;���[�[������L(Ӛ��Q���n�V�c�\KY�f��;�)8�MbU4M�]��v,}���� |���j���ه.�j����������(�I""�s]Հ�׀y��%DB�ă���0�<��9�Z���`z��K�`|�N������]�ՕWX���}׀owb����9u�@=���`&Ҙ�Y�M�kL_�I)�~_2[���`H���U�m�5�u	�z���M�'�t�v��a]h��M�*6��6Z�y.8������V�%��>���֘�WX�l����dnf�˭{���?� �w^�݋ �;f {I��svL�T՗5u�z� �o�B�I�'���EҨ�~���rN�����%��h�`���@�۹�wu��9u�@=m��yr���2L5n�gr`I+L	��`[y��k���J�&��kL�<��Ό�TE�8��2�l��8����ٛܦ��7
jk?�����s����s>��� ��h�����s@�;���M�0��������uJ��X��]�S�"�ɠ}m��;��h�נ��ʇ;�jb��7!�J!)������ >m��		DDB��4�Ucq�6�q
dnf�U���٠[Қw]��/Vےrb�[�I��77�p�Ҥ�9�՜��G�t���c����:���t3��-���uJ��X@³vK�D�*�swx{l��(V��}�@��~�@=m��y�H�&���L	%i�2[��o0=mi�}�vY�`�Sȓ��r�^�_�������_f���u�$�S	j$����@��4�w4
�W�?=�����zz{���o���� h�` M宅��i�sa��y��'7YV�sv��^����.ܖ;��k���m�܅����Flј�{&���	����v4dZ��Ş���}G;DlK��rR��(�P�mcC��cp���DQu���^�[mQ%�N���]�5��b}�*{V����Rs���=����CӺA[�㣵Ӱ[��+���T�Ĉd�.�tҮ��aq�WK��8y�����*뇝ll,�6j�y3 �JcqdN9>���?Ɓ{��U���l�<�$���51b��'�Z`\�� ���Σ �ܺk���܂S$s4
�W��f�����Q=���9�ŀ�Ӻ.nɚ*f�[���/������V�,����u�"LCfɠ[Қ������:y�`�w�	�f]]YAB�D���]9�.�Iq�3kr�.�*l"�N3��=�Q$�K� ҉$��$�4�Z`L�� ������<�U圍�Lpo"Nf�˭{���?�
�^�����8�iL$q���@>���֙��IZ`L���N�M�1��G�rh[w4w]��Z���h_;�jb����}��`�DD:}�����<�ŀt(��K�����M�إU��] ��W7euV�M�ɮj k�2OK�gA��R�6D�R$�F�x
���@=�f���p��r�v(�c�$���������V�%���p�l$H���@�۹�{��i����~F���H��X0� Ē D"bł�D� ��a��H��1	��!m��D
���6�� (���� �A�R�-3\U��[[H� E�
-��	D���H,U0B(Qu%)H:D*�H�T$V@DT�@K��$�P�UA���M�F ! �C�� �U��+ T4�O�pA�A�{�mD�lllo��؃� X � � ��0��rنa5�ffy@lw���A�A�A�A��kb���������6 �6 �� � ��{��A�����Oap�%�f�lQCz�l؃� � � � �]����B�����}�y,l~���b �`�`�`������r6([����j��e�$��$�wV�q\����V����v��<�����j��q3�.��?�������o������D$�{���o�a�"Je���$�Sհuu�Lڪ�V�������UZ�{��78
����[�O7��!/�=:t�XU*�����ʫX$���� �:}�����<�ŀ|V�q�!�D�E&h�׿���7$����rJ~D_���	 ����_fpܒ~>�̙s,�ŝ߳7��}�y����0>����}� g��s�@Q�<IL�� �nm��$�T��N^��B��&���Ur+м��ԡ&
!�$�h��h�נwY�{���D�Q`ؿ-ٹ�<��â�r��������$���߻��g[��h�M�V��ʻ0/�VtDBS!���%	-���y���ď����q&ҘD�i<�@���f.���7��`k�`:Ӭ����)�LJ,��rh[w4u��9u����4��ٙ�ŖI2I$�I$��   0kg]ͤ�ܬ`��N����pO���]�����Fd�u�V�����	e*v�24�]�8�U�X�*����/���>��(��{q\X�)ug���	
]il'<[k��,�=��i�[��Ӣ^;0�pVs�$�= NM��]7S�5U�`O�#=�����Ý�y��^����=[R�΍4�\���ݍ=�� l�ʳ���iL���]P�z)�iy��ܩk��&���(�v��B!*BcQbQ�A����~4]r� ����n�u��n6D6H�i'�v� �������^� ���QH$��&1��}�f���s@�YM�]z����H�&
!��������^�ݻu�zK�v:�D�$��9���h������>��hΥ��6b��}+�m�TJi*���n?f���*<��u.�U���Ӑ�L
d��A�xߟ����]�m���$��}|`M�Q73U3h������� �뼴��$�)"P����Phd�����?~�~4]r����_��&(�b�ɠowb�>�l�6u�X��x��˰6LX�p�s4u��9u����4���׫I���"����d�� ����֘K�`Ow����r�^�l��=]�`�ΪvyJ��.�VG4n(X�V�^�"y:h�ʹow��]��^`z���J�d������H�#�D6I$�>��hzV�%WXޗ�E�)ٝ��.�4IwV�����:���TB��_u�^���u&���x�$�0���l�� �����������.�D&%0�G	2= �u����/��}� �֝`hkʪ��T����!�;���t3����s!��bk�^���,##H��q�cD�LNI4����Z`L�]`���36�b�8ŝ�ݛ��Ҵ���Y��S�~�4����u�&�dCd��#���*��/����0/�i�yL�v(�l�'�O#��Y�}m�Н��vnAW@������nHۃ�ɹ�.��*i]]�ͼX�B�����9u������:T����p�b�T^li�F�+1����>��vÆ���v����X�"!�LR`����]L	����Z`[:��J���46Nf�U�@�[��[Қ�m�(�ĦE2%2=��X{l¢"�~v��i� 粡��y$��[Қ��h^���w4+�'`,l���3x`Y+L�+��Z`[:������ �� ��մ�����n.9�!�9,g�z�J]t�`�+�7G;��G}�,�m��c��mkn�{f�&���6�FK�v�5��Xۮp��B�wiF���h�N�<�7�h#h˫v��=sl������Tlu�P'���{1�L�z�5�i榴W&0�<4ڇ��=*:������Y�&����A�%�4��MӛZ��f�95�XWtQ��L��b�S��E�H��}�"ƻ8|*���F]Dfn���u`����g�IBK�o�4��c�R�c�y��n��J!)���o�`^�X�`u�1�F%1��ɚ�)�^빠U{+�/��h�t)�LR`��R����b�����$�Yn���b	��46D����^�~� ��0��`୙up*�f�K����4q�&���x:9�+�˛\l��\h����BbS	j%2=�n�oJh��h^��
��C�&)J�ʫX{l�
��˧ذ�k��/�w7��٘��䛰6Ab�AMY�?kŀ9z�a�)��ذ�|`��[M��Cd��I�W���^,��`tB��S���ȞU֢�L�&$�=��s@��4�]���^��e���6�� 19�cf��)W3���i{-䶝���l�փ�]�%DbS�G3@��4�]���^�~빠{�QH�Jb��"�`��gD%2t�]Xk�X{l���I���s"Nf�U�@�������`u��<��(��hJa�dz~�h���{��U�@�쪨�M4LQ�8���֘Ҵ��*��/���m��q��6����wY����\�,��GOl]�Z8��S-�\ZZ����Zl�0,���U�}o0=mi�|�+i��l�2I3@��+���@�۹�^빠�.�!��rb�]���`z���Z`L�]`wvU�dm�0ns4����7$��Ӻܘ�(� |@J$0H�"@�Y�Q(��"�"@#$H�c|�U	G�^�X�'3s6��D�uk �V�%WXҴ�����W���]�]vѹ��oFe���]����tl��;�&�����"�d�0`� ���9|���x�6�~ID}!����[�X�4L"������]����ɽ݋ �}� �֝`|��UL�Ԗ���VMZ�<�ŀ?kŇ(��Ug�~��s@�v�ɂ�I
�X��Xδ� ~׋�B��u�/�M��Cd��I�.�^�}+L[Z`_J���O$��-Ib�,bF����v�2O�<X�,R���%��=Z�4�Ū��b�F�V)6�*$N�� � �B:E�4XR!"�g�0�4�*H!�ND4�PHV"B	�}R�ĉ1"``����P���t�M���#,�2�B$��J;D��b�!��D"���D6�LPM�����$XE�A`�"Dd�@�B)�+D�����     m�        'l  m�             �^�lm��20�7CU@%�)�
.F*�)���Uu#�V�]�͍���y�7\�߫\�>�Rt���i�;m1&B� �ƎmmTI���R��{m �����{}��s ��J�DK�M�'�ە��SZ-UE<��pR��4�Fr#Ӳ�t٨Vy��v.��A�s*������]��� #;H������*8�P��6�y�l�	�[,���%b:�#7jvր�e�K�0\��IB,��\��Vy��,5�Jκ n]�b�9��lhcpn���9@:�ܪ��V�H�8C]��C�X��j�����E�X06�6��dIċm�a!c�n���嗊p�C�mյZ#�C�[7&Zc*#P���6xw����ZSsh�ssϡH�vkY���:Eu���r��6�	1rD;,֩�,�n����)ŧ��hs� ��6�.��d-��[����Q[R쫺�D<V��N�-]�(6v�k Ql�6m���)��M1���n]c;.B�>X�-�Y3����C-!;���-xs1��2�K�m��ϵK*=����cp��ML�YmJ�$�� �mT�$$
���ܤ��S�g)U�Ç�;j�#]��ğ\�΁�[j��6�|K����8�A��WS�b���8��6IT-�&!�Y���U:-�
�P%jyiG�U��Z���9�;S#�iT��:H`��,fǎ8�L��� x��X
�@��V��	Vܸ�,n楍���<��Z�\�j�Z�u��r�U	�ɍ]Hٹ�������㴒:��V�v��^�m�.j� .T�@��a�س�ڡ�ŉ��3�<H�8��2WA�)dF�vm�%��Ӗ���nڶ��RUge��b�e�F�Q��-� A��fv�T���K���-����T?�@1�x� �A ߄D�??" ^o��� �  M`�s\��9���(<��]�V��z����Dt������r��yd�/���v�fn^Ll�gk�3�������nnn�;�5��0�Zۇo1��+�e�I,�����Lusz�wJm����t\�m���{z�X@�x�yGm�� Ht��a���M�M�ۜ�s�=�:��`�]M����%�e���\�S���.��U��N.�$T�y΄��]�b,GӃ�:�E�kHo+�{:�x'�B(��c�y�?~��s@����V�%WXEY���;L�F�w&��0/�i�2Uu�}+��ʊD�S������s@�*�������0���3�����q�Ɂ2Uu�}+L[Z`_��h��BƉ�R7��~���֘Ҵ��*���[/n�F�=W3� ^�Ff��lrU9/6�Z ��y�2�5b�r2���M��m���Z`_J�d���V�eɻ�B�Qh�eݕV��x��F"��I��!B�(I!]�_.��[07w4��M��Cd��I��α���F��0>���$�"��ga�r$�I�{�S@���=�w4����VLq�b�����kL��0Uo0/�i�/zf]��<�	�qs��!���:�n�\��X�3�@q��^P��Z.aƦV����ִ��֘��ԉ��L� �� ��@�[��n�� {�r�=ΜSs*iZ.n�U+��;{�`���ˢt�(��� w���h}�X�h����:Z��Z`��aYZ�>�fdU��ɂ�9s4��@vwM��s@�s@�-��I��Q�m��Ⴌ�WUi��y5�B�3է@�=/8�Q��kf�ƛQ���##p��[4��h��h���w$�*a F#�5��-i�%�0,�F����c�h�#I���;���/YM ��@�n����I�18	�wo&���=U���֘{���-�����D���hl����[4-i�%�0,�F��]�Ԅ��x�!��z��5KOmN�dx��o�n���xme;s�Ք^=�N ��S��6߿���v��n�z�h�-�]�U���h��73@�s@�e4��������,������/^� �V��Z`IkL�\�25�"��\�h��h��h[)��.´H��"O�����֘���=U���@��H� 	"!�����0� -�  u�rőz���A ��bNh,];.2�vǝ�%��*8�8ۭ9��a�+NA�Xn���]?�G���u��m�n�p�ջp���ͮ[���j�%���v������Nlr�I.�ٖ��sq�v[�����;�r]q�R9����O+��f�n�Θ���������۲p���u�y3���%�n��.��4]�w��n(%\i�'>ڵ����m�IXi���\�]i�Ev%�76�k�m[I�ή�Oi�[f�|w�ذ7l�4���K���`~yQ��4�'19���h���Z�KZ`��r5˸7E��0Uo0$��������������a��&��n��n������f�˲���M4D)���;���>�S@>�l�;���>�-�ۓ&GcM�Z!�SPХ��ʖ�3�vY��Z.4.ga���ɂ�I�h[)�\�h��h��h�9T��Q�)�n���~�'Z�z֘�����Z�a��d��c�'�M�߷4	-i��z��[��p}�7�v�n�n�`IkL[�`��a������>���$Ҙ�Bb$s4_Y�:!)�]��ϱ`���[��Vyͱ���o%Q)���lf�G}��l��6:��eD�u��][.����x�x���`nـ}�۲�ц[���ff�}����6���`�|`�n���.�f��-M���Z�7[ŀ7Z�!(4�����<��`<l���N�.0	�o0-����0��s4��dj$���-��w4�Jh��@����ňc����)S�)2����9�= ����3�1��W�H�Ba&L��9x��-빠}zS@��Z�e�@��q=�DG����n�`z���e�<��������R$Ҙ�Bb�Hh��@;췘���u��.i��g.��.��p:!(IL�]׀w>ŀy�	���{}�ܓ����.Z]e��kGw0-����0-�q�O+y�����?ݿ?�����}wZR[��Yn�q�+pY��u��*��j�o��Q-����_?�v\`��`[+L/���&!&$�Z�� �٠[�s@����{��I��bl������y[�ei��:�vU����d��c�'�M޻���0-�q�O+y���Y���v�Lcp��}zS@��Z�e�@���>邏���?�� .�   4��ͮ���%��N��&M���-�+k&�iR9D�]�=[M��x��c];Pu6[<���������6޽2+Z���:iĘ̰��s�%�r�kӤ��66����I䮸9^.�Ʈ�����f884�i���!d��;O؈��:�]���H�N�ju:��=�7#Y-Oh솆i*�j�g����
�ҋ�9���{�����_C�t�m�Y^,i�E�+1�`��.�������m=y�X��X-7��R���Z�e�@�����M ��Z2`�S��9"��-������F�.0=��q��cdȔ��&�o]��Қ����-�W8VF��"�����0-�q�O+y�l�0>�ۑ&!&$�Z�� �٠[����$�}S?T�S6R���'�7K�H-2������s����w@uȱp���L�$��16F��N/ ^�ߦ�o]��Қ�����+Dɑ�7WD���׋>I$�*��0�}8�gY�{��LQ����73@��F�.0	�/0-����2��Jcq	�E!�Z�� ﳬ�-빠z���|}���<�0l�H�yK�ei���F�.0'�`~7e�)��=�ѵ=l�hXf#���듣���l䮸ټ�8��ף$k���zj� o^,����=��z����+�#ka1)���=zS@��Z}���;��>_:�6DJ��L՘ε��U�p�Ę�*�+����0g.��"/�!'����`�/�H�B X1H��h�n"�E�(�a #A#�� �H�x�,jP
��Tj0 3b�QT�Dآi �#U?"@u����nI�����>�U�Fɍ���8��U�w�)�z������ ���@���"y$Z}Қ�Jh���;�}O�߾�{��{���Y\�m��3͚�fC
U���uԣ<��=���3K1Hʵ��j6
b�܇�������Z}���-빠}_
��4�7�)��nˌ	���Z`}gQ�x�s&1�#�-��j�-빠w[��Z����E��,n"%$o���V�Z�ݗ}�����둵�������h��h��@��i�V��ԒV�6و��$l�!����b��Y������<v=�br�L��!�d�d$�s=䒵�-I%��j��Jۺ�K��g��B�i��cmF��NRI}rZ�䒶����$��QjI%��´L��)y^�I[wCRIw[���J�(�$��%��I/�)rLm����7RIw[���J�(�$��%��I+n�jI/^�^D�S�oRI��IZ�����{�%m�I%�o��IX.(D�N�@	,V#Bt���߀�    ]���Uj�I�W��*mX�tfݶ�$8�]�g��\i�^۴��c���az񳭝����>��یg7��⬭��m7q=hĪܙu��uN���D��ڔʗ9������G��ٶ��2�l���a�%�P�ͫ�tx;k��d��6z�5�M�����Q����v?�N����6�h�C��p��~n�wwqt��l����`:��v��Xn�k�� �u�';�k=�>����bH�����]�6G$I%�/�{�%m�I%�o��I+\�Ԓ^��iL7�7�E�$��t5$�u��y$�r�RI}rZ��;�R�mby ����jI.�}��IZ�����{�%m�I%��s�!�d�I!�y$�r�RI}rZ�䒶����$���ZdO#q���Ԓ_\��y$����$���{�%k�Z�J��[nI��1wgss�6�-Z3����͖4u�r�6򺓳���xFɓ#1�#O#��I+n�jI.�}��IZ�����{�%��.I���S��jI.�}���������Ԓ]�KW��V��Ԓ^��e���oRI��IZ�����{�%m�I%�o��I#��d��9�drAjJ�7�պ�V��Ԓ_wnn��s�-I%��Cj`�����d�{�%m�I%�o��I+\�Ԓ_\��y$��lm���mb���d�q��͡Y��a�K���`�匏<U�۬6�by �#�@Ԓ]��=䒵�-I%��j��Jۺ�K�>�lC�ɂ��B9��IZ�����{�%m�I%�o��I!}ʴȞF5#s)�fg��s�3-���k����/���o��$��n�I}�sJ�L��)�E�$�u�I%�o��I%��I%��j��J�����n�����$��݆����{�%�wCRI���~3g�箧�>�\�B+:&5�M�*p�X�3�ʼ@ݲ�V�c7�$��$��݆����{�%�wCRIw[���H�yhɃ�Ls���5$��%��I.��K��g��K�v�K��|���cq)�"��K�����$��݆����{�$}�R�mby �#�@ԗ�����I%߿�33=W[�}���^����y����#�!�d�I!�y$���5$��%��I.��K��g��Ue��rLq=���˴���4�6�#ί<]L����h��s�f�	�Q�v�)��[����j��K�����$��݆��_r\ҭ�&F1$��I.��K��g��K�v�K���$�|��1�6(�np5$�u��y$���5$��%��I.��K׵*D�S�oRI��I/��jI/�KW��]�t5$�u��y$�����<�0O9I%��j��K�����$���O�������w~�???� ?���m� �W��L,ӫ���Pyĳ��;Z� ޮ�s�v�.��ؓ�w�zv:H���N�gDN�ݕ7=�k�8&���kl["ŭ\����ǚܦ����*«u�;�n�&xY��!��޳�Xآ�n�A�s�ms������S�NɺcW*\a4r�0���ڞ�ƚ�� �M�e9���ӎNuƁ7"��HL�v�狌ˢ��:��5Wl�q�?}��6뾲�{k	�=k��S�NR�cq)�"�$���CRIw[���I}n�RI}rZ��3��Ʊ<�J� jI.�}��I/��jI/�KW��]�t5$��}���`����g��K�v�K���$�u�I%�o��I!^���0��E#r�K���$�u�I%�o��I%��I$�乥[&L�b��$��I.��K�������n�o��o9m����޷��H'���L�7��vI+=�z��i�9�[�sl����U�up]��-�$������I%��I%���{�%�wCRI}I��Ҙ�M<D�g��K�r̨[P�B�.gZ�������������y$�����<�0O9I%���{�%�wCRIw��=�_[�Ԓ^Ϻ������"R%���$�u�I)�7��陙�yfL��J*��>�����;G��A(G$��$��}��I������އ�I[�7��$�u�I%~�|�p}*��-��)�$�03P�֮F�[\�:��y��jW�.��������FD�g�D���]���RIw\�{�%�wCRI}m�{�$+ն�F���nCRIw5���J!*���02ffw��_}33�o(����yP?���C�u�Ntȝ[������ݶ���xs��̿w{ɻm]�ͧ��K�nH�)�np5)�
�{���fv������ֱ�}3?�^��O����_ ��_��B�x�K�f}M�33?�(o��{�$�ذ7w4�б6�ƛ�&,c��ne�%5��m�]s��7�/�\�R�=��������u�}��H�Uh�����w~W��>�x�7w4.��g�CS����ۯD/������X�w��7Z�0>^T�s�V�˰��r`z����u�$�e�W������YrTԖ7suk�%>o� ����>�x�*"(��G��X��UM�Z��������=�[0Jy��|��� �u�}�ZZ��	���"JL	l��+:��3��Ҭ�l,���x}�G$�l�21������s@�����]�I%�W� o>WwsatL�WS7k ���9D$�C����0w]���YbCJcq4���v���láDL��ŀs�ŀ?��-��V��Wx�{�q�y�ŀn���$�|�^��D��*��.g�7Wp��J�KZ`Iy��WSrO����ʆ�M����B) vE$$�CF���am�]��I0�i�tE��Ԃ��HP�A+�� E#	#�s|�UT]C@$�%ZS�Qt#2�H��P� �H$�j!�t1#�t��!�'�Nl7 &�Hn�Ow_w}�    �         $�m�  6�             e�K�N���cr-,Yغ�&�ivZ��s���z�W0n�+��6�^��N�޶���$��K[�m12q�۫n2e)�&�T���ˍ�m�NثmpᣡX8ݤ&�<9��QͷUu�7I��3BmҪd8s�Ƿn%Ce��t���%��v�����ba��2��������;j�n�ɮA���hI��U2�	�v��ɵ��a��}%��gm��5��f٨�m7D�XB��Z���l-���S�n�v�mˣg��uvb ���H4Hiݝ���5�
�ZUg�ɸ{c���og6�ڕm]Z6�8�V�.�R���tXר9 �m��T�Vۤ������W.�+[G��Xݒi�6�=@&�q�mѤ+Ng'�;V�K��M V�jݮ�skoR9���(v��IM��n`#4��Ύ��N��';�G�.T��lY�ˡ ح�C��ڛ�%yJ����Vg����8��d���p،�Q�:��v6yXA����G�`��֖l�5Kb 6�Ӻ��5��P1�X*��N�U���3&9����P2��u�2<b��� @.�dVyb�p�W]�s���Zb4�)��;p˚�H\�mk@W[r�����C��l�	K&��i^O5U4�km�U73��%P�g\��lq�`Uj��j�]��mS���R�UPr��@ ��U'�ݧL�JB����yV���:U�讃m����
�Qm�­yw-�v�z6�j��ݥ���.kB 2�b�T YV�drkQ��x:�Z���ec��0l6�K���[R� m��C%O<6%b�6��i�y5��;�.�G��,�ݪ��.x�u��mʝ�˶�G�Ꞟ%�A�J��,�3ı��-�j�s�&US#���jf�4]]i�E�ت|e��
�ؠb��E��}�fg ,�  �#�&6�y���h�Se�=\h7��F��k�D�n���m��U@Q�X��Yvꈤ�L���j�أl-��Y�ynP�EP�r\�(��B��kSd�vtb|��̝i��6L5�RĔGj�����slNH���@��Ԫn:�;g�p卵L�Ny�竑�z�v��V0�3a�E�����S#���$8��Vʈ�}wXӫ���+��A�E�ح�N9⵷M�%vC������}n�Iyn:�N��ͷ��v, ��ͫgDG�_b�=)���� ?�#��z���>�%4n�X�x��d�������-U]�s����w���J�KZ`}%i�z��J6H�9Y!�{��hu������\���XI�1{�;��֘IZ`zU�`}%i�����~}�u)�Na�d�-Y�k-���.���n�t49<��GR��Ì��w�swo/����0=*�0>�������U�#Q�������0=*���CJ��r^����>�����^,�	DD��ݝ%M��*����R������0>��������y��M�*�R�Yj��`r����y���uIZ`}�۝���o��7�0>��������J��ך�c�i��(�Cd� ���"HYz��Ƶ09uvp���̨�sܷ����LJ����0=-k���[�s@:��?F�d��L��=%i��kL��0=*�0Yx�ݺv�h�w�3�0=-i����w�ߵB�Q	R�_+� ��ŀ|�K�4IS6��jj.��$�O�� �+� �u������U�#Q�������0$����J��֘^��6f~6�.��YNٶ���F��LGQ�[���l���V���)�u�ճv.�<�%+���֘�����U�`yvqtq�nbɐ�䙠}m��;����\��>��hA�Ψ��2c���ܘ^�Ү��֘������%BcɎ5���>뒚ּX��X�����`����d�゙!�}m��>��h�3 �jـtD%�\������ڹ'Cj)��l�QٖD���.]yz��ҥ�k2ˍ�!2F��3q�L�����u�M�s@�<���4�7U
�`�l�I$�F�_��X��0/��q��g-�f�;��J���+L[Z`}�Z`|��*3��V�����]��J��֘zV�U�`|��^�n��X�q˻�0=mi���i�%]Fޕ��������w{��� z�  271�5��۬�{8�;v.�m���5�u��˳��ՎE9C:���v ��t�s��]5ym̻K`ۊ���8�cm֛Ӱ��vp�	$<^�܎�uu Sbn8sv�{O)�zD5�lQ�/<t��l�aGe�1��s�,���1ikX�:M��͎�e�nG�Σ-�t���3̀�nnܽ��'���O}}*�[`:�a�zN�Vf.h��g�|Z�pÎ�c6�����n��b2&\��f�ܼ$������J�������P��c�d�M��tDL��ذ��X��� {fu���Ӹ;M��9w�+L[Zg�Y��\�䦀}��6������� ���	*�0>��0>����0iLn&ْHh_uzu�M�u��>��hY�iW��A��R`�v�0�j���Qg��9��]����~m.����������߀��w���Ҵ�����	B�Cӯ� <�P�*ԪSj�n�w�+L[Z`}��XU�`|��ǻ۫w�.\r��L[Z`}��t뒚�빠y|�+��4dǐ�3�0>�K�	*�0>��0=mi�QnX�a1�Ƣ�qǠw\��=�]��n���W�U��mǊD����]ך��Z��nJ)���X��]1͊`��s#m�@�qĦHh����kL���Ү� ����кU\�v�kx��D)�ӯ� o��}�x��P�O:]U�D�3j�榢�`�}X�V�&Jr>Q��BK^�0'�i�|m*ӑ��[�����7Z�`{^,ͼX�%>���1��V��۝ٺ���+LKZ`}��X�uR^���Î������P�͡Y���]C��{0�.-�8�1�) �� �Q�Na�!2I3@��i��z�`zU�`{Ҵ�����Ҧ�WAd�7k �|�g%&�W����orJ"d�e<h�Ss�ݬ	�zV�����=n���wM�c�%2C@���hu���9~�u�+�"� U}���BB4F�ۉ)3@����>�n�=*�0=%i�)�w��q�ܔ<5j0�b�Ea�Dƣ��b�\�lg��*n�����!r»����%�����������0/��ZL"S�H��䦁�u��;�ŀ}:�g%
D�yl��U�T�����R�0o�`��Ò�Jg��� ��|`^M�M]J��+VZ��X�x��[�ͫf(��:�|�H��H��FLy�I��Z���Mۯ��,�IBIwe������݀��  �ۭ�2uJ��8�n<�cn��y�5�u٠���� {&礕�m�nvx�Iw޺pvۙq�5n� kts(7ny9�5�X�l,y��nb{M���k�������q�/Y,%�BʰPj E�k�wn��:����4�ӷ H&�ri{5�w.���tkb���,�t=�<�p�ǋ��COd�5q?���~�V�6�n��	�nm���uV�Mʚ�[z�n9.�E8�k �, 䰺Uu13Ww��_�^,u�� �[4���d��L��=��gD��v, ��ͫf |��HF��3q%&h��h�٠}nJhw]���N�!�1��d;y0	m��]F����֘��q�)�l��h[��[Z`IkL��0
�72��-���3"G5�bU���7;�?��ǝ����Nu�2f
���İ�Ǐ�ԉ���o��u�X��/�$�>���|`�q�e���
Ֆ�����,��J$�������Q��+L�Mͻۦ��j��r`}%i��WQ������`[���U�G�)�Ƣ�ԙ�}Z�`n�X�x�9O�� o:��l�#q)�����n��빠}nJh�uik1f'��\L{<����Ӵ�u��Ĳȼ���m��
ڶ�]�&�� �@���II��߷4w]��rS@�u��=^T����n�.�`n�Y�B�2or�07ذ�w4���Ʉ�6dRf���;7$��wf���*Q>B�Љ�DNl5� ��1��"J(BYBe��#�dIv��b��A��t�FD�!FUM!ViuKB$!"� DH$$1ր���!$"�&�3GBD�
A҆#&�5�!A�A �Yb�&��� C�`�H����@��B TЪH�����`��� T�"@��B+0��H�N0���Zf� � �6�����!I�B(Db�mYQ/�@�"��Q�)��Q@�((&*#����� ? UD~S��ɰ�����u��g�A�x�L�H��������0>��������yR��՛�\��ܘ������z�����OƁ�빠w�n��F۷�=��d�=�ʅ
/&��P�]�x�t˶y��V1L��⍍4dǎ'&h�]F�V�����f�չC9�;?f�r`zU�`}%i��kL�������6��1�	�Š{��0%���V����J�@���II�^��u��:�괕
G�UKb�~ ڣ���� ���'H*f�U�U]ݦ����l�����������ww�;���
ܼ���2A��6��*�m�\O���//\��:�b�DVr������d�Q7Svx���N��,^�Xu��a�\��<x�F�k#�@���YZ`}%i�*�q�����7��q�{�0%���V�J�����w�X%�2c�G&hIZ`}*�0>�������o.�Sa6�U7*jn���l�?DBK����5�ŀ}��`
Imou�ݫ�� [F�  �Ӷ�*m�MA�$��.v��wn���8g���;q��OcX^q��mZə�kɡu�+ci��B�
��gc�vᛔ���5��U=���y��L��ۣ�%�N�	vi�=�����Յ�[�X�nwD@뙞!ɛ��%y����"�t�m͏q�5�l�@�:��Nݨݗ����=@�.�՗*��s���!󌦤n��+a.��+0ն뇦�F�p>�h&bد/�H2F�1�F�9����߷4��L��0>�u�J��C�;E����Ɂ�+L��0>�uIZΏ�T~u���H(�U754���X�~i������J��V��
��q6�ɚ�K����>|����,ۭ�%��>B��Vr��帻��x������}׀}�[0���[v3�����D�PU�7�N5l��c\�s�kѼJt���i�&�y��r`zJ� ��`zU�`z�� ��eM�5"�J��*�`�w�i(QK�+�>��݋ ׯ ��-GL&5I4����n柒���� ��������c�a298�x�z�`�w��u��0򿰐a Fcn$���s@;���rS@����=s�II�F����(¨yc�Z�X'�k]�s�]��t5���7�7,�I�Ƣi�$�4�Z���f��.�C_v,��r��dګ37N����]F��0=-i��� �ʪ���Y˷;�uwKZ`zZ�>��J���WQ��!p|jݹV]�ݬ�}�,e�V�jـ}��h�w�M1�#��4��X��f�o�o�(���_�~�o���r�x��֐ffm)���2�ŕѠ�˖R��`�3u�l]�H[�ݿ/����kLKZ`{%��>9[#�ĦHhu����H�݋ �}Հ{Z�`��L���UU�MU���,ӭ�
g_+� �����T��b�j&�,$�4��X��f�o�W�Q��Q�"~ �;}��s��5<ja2\3&j�����ճ ������}ذ�Z��>J���)�ģ#��icB˦#����ś#�!A�f�Yw=c�s۞zn{Vr����]��֘���=-�����J=@��� �q�rniU\��.����֘��������֜���$���yL�SR)RUMR����=���}�v�����*�d��F(����<ڶ`���7[ŁВ������UAtUթ�Wf��,KZ`��֮�z��ܻ���M�  fY6vEU:�+���cnu�6�]��Ѱ)�/�OX J!�%��.�6�;z�����x���Α�u�vƭr��.�\�l��k�]2���Ƌ�Z�i6����u�<׫F��%ǖ5�qԡ�J���zuRi��Lln��۳;�c��+n��,�>��y������V�m�iץ��1���HkS$�4qT:��ֵ�ֳD�Y�����B`)W3[=iԡH�4��"�Lj�߽��-��J;NӹX�w������0[y��WQ�%�0>�sn�b��M<rL���@�ܔ�;�ŀn��:!)��ͪ�E���w3J����W���,?%2�v, �� ��YSj�&����R�09%�w~��w~�� �v�ͫf�tre��NG.;���KZ`zޣ֮���n�{���X��NF�v����̮ŻsvQ��l�����c�{4�7~��~��%���'�I��~���rS@�s@�s@��:L�a1�ɫ06���)���X}ذ7l���FV��1��Hh��hZ����u�J�w4;C�UUrM����!B�����~0���0���u����׀�1��x)� �v��%�(�ܾ�x�߱`�S@�ϫJ�����_ͥ!%�ݪ)�0W:�u��ghݖ������h.��h�\vj÷y|�����+L	gQ�������q����7��k����2>w���ŀk�l�<�ʍ��Ʉ�H��hzS@���i����C6AO��P�������iP��M*#�%�����_� ?ou�i�S6Vnv#V�j7x`}�Z`KQ�{���ץ4
���IF(��f���\����S}������=��`ÿ?��Z�����
�y���aa�k\�t�Xt�n�9��n7�̺:,i5�9�i`�{�o0/�Q���k�$������@>;�썦c��&�~�F޵���q�{���ܻ�Pi��njiM�՘�o ��\��	L����?u���&_�1AL�'�(���V��{]��l��J%�D(]
{�׀WO)�2j�n�U�� �����0�o0/�ˌ)?%]C�;��Kص��ő��FG�@�Úϱ�vڟ#���۵�Vyu��PM���l����ʵ�DD/���@>����J5O��٠?*�8�k��m��2t�R��a1�NI�~�w����4�Jh��4����da�28�?)�k��;]�{]�~�	Oj�Ӏuƿ&c1�rh��=�\X�s�{]��Q�QJT0 �(�*���R��
B�.�& H|�G[F*@1�#AYB�H��4CA 2 b��X,A�.Ņ�%$D�3w��fffff   �         I��   m�             �7r7ky�7��UU��rJc]&h��.� 6�Lj]��`^Ul��mPӧu�9R���0�B��l�oUӗ�{v�9ظ�\�*�MLn�m�eA7ayKd�!��㶐IIcx�����S�R��BL�̰=���*�؎{[rmT����b`�g� ����*�%eQ���K�*v���8B�[�2�T9�^۶��s���zj�n��gi��� K�(�>��-�P2��ԨIڈ��s+%�U�����uv͗����\����Tb����d��[u�[Jd@c�͹��7jI3����WشN�$�GI��]�T��qtݍ�]��#�N�/6����v,�nM�X��r3q��e��m�2����*6�tiom\��Q�m9�S�[[.��-����N��� <�x����mv0������X�=��J������PL���C�ݕ^,�ٚ(��U�H���n鮧D��N3%J���2�r���̮P6v<��<\�����ɓ.��\��]��[6�Z��*�g�O����Ks��gg(��^��qlrO+��u�C(��َ�eZ�8�˞�*���d��m�h]��iN��=���=P�N����m��Q/Q�a#�vl6X���p��< 6N;A���̮n��iUW�u:y8��i2� 	�/i��ؕ˴HMUP ��@  z��N�ɉf����,�݊ʰ]��Ke"��v�	(��ٛ/RMmu�1����N��m���9���MPc�sgbZ�yZy^�	V�jm� Ul�T��e]��n-ڶ�UW��U�TƶB���$��1�2`d�����<̻mm��ʹ����1�[��8䖬t�[I��t������tq)-K�W.��v��T�F-�l�W<��d%�:��S�gp��������www�P� Z(h >PG�?<Ҥv ��6 �hTB(���;]�ow���33333332@  M%ѫ�nt<�6Є =^�;�1X��Q�a+��9��h��>]����Ë��;ڴ��5����۫�����\	ri�Vɭg:�x�N�R���Y��gau���c�;�󢶛��e�5n�Mn�e��v�l�c<�h���nj��6�{;{rc\�2�nU8�{�c��-��Az�wql.���{��{���g��8L�Վd
9{[��n��N��t�Pٲ�8X��u7)�T�prQ�1Lj&�,�8P;��h�|� >�����|`��jl�]ٚ���L�� �����0>�x��(�C]ʦ�HM�����Us����Ө��Ҵ��[.0<�K����	��
I�_�S@=�Y�_����}�� =˫�͕57(�eҙ�ޗ��e��K���`z����l<"t�u�MMjA�Yt�5�-8h��f�u�:��s���7�x��q�}k�Q&ԏ�~�w��}l�/�)��� 4��_�͑�c����}no�E��FH2%�	
��BR�$��w|`_:�5�o� ������@�f7 ܚ�g�@�z]`O-�޷��̺�Lks�sV.���K�	�� ����}�8�;��jl�Ws4��� �'�h�[4^��[f�\�X�r�+l��	h�갣5P�����9��H^wJ울���������غB��<�߯ �� >m��U� լ��68�d$D�hzS@>�٠k�l�y�Ή�i�S<T�`R��D՘��^�f�K�BQ�$������0>�1
���G-Y�7$z^�M ���^�����ߞ�S����0�rA)���4�)�r�@��S@��ZZ�Y��g,F�e�-�"֚v,��=u,�W�4ݜ��i�Y�ģHb����nAI4z3 =�� oU����@��Φzzp�5O��@��^�od��z�4zS@��q�����r6�u��`[:��^`D���5��"RH�C@=��ޔ�n��q	
e�`^`�YTU�ɐ�I�[Қ�u�����h�[n6،p�cB�l"vYyU54[Y�n�R�v�^�MօH���]� ��A��4��Z}���u����|`����&�j��̕wx�V���!��x����y��3�_�͊a䂙Z{��z����Jd�}x�O� >��.�.��U]�����S�y� o>�|�\�~K?�����;�J��S�o	#��y��D(P�[���u�=�`� ����=��������ff[w��  ,o�I��v�nԽπ�UL��]����X�M)�0{p��Y���y�q�K��]@�[n}�����Y`���q!v��9��<<�Fuc�D��y�z��:vDm��Rqظ�8�����m����.rkZ�{v�;�Kv��f�;Yě�Bk=���r3c1N7Mn��B9!p�Y�6���Omw�;r,������wn-B�-��V ���j��ݺ������/-�Y)z�ŮH�w*'�0�L�)�q��?߱���@;���m��
>�����Gr�*��&�Ĥk�@;���Jh+k�=��@�}J��MLY1�(����M����ϔ����׀!�K) <�	�@�^�@��Z�[x	)�<� ���w\��-R����� �O����P��u���� <��~�ZZ�6�#�)�6���C��Y���r܏L�4�^����I�v<)õɺ];LrBdR= ﭚ�v� ������q��@>˗�a F3���4:nsQ�"%B��׀5/�`�l�;�\�b�o	�@>�f��\��%2=��]Ӏ}�uR�Jd�LmI&�ݏ���٠z�V��빠�ܬs�L�'�Š�� �
}���ϱ`�������⭻s��<6��I�ֺ)���g��V�� N9s[vo]�7+�&��q�:���`[y��+L	ˌz�`��T�����wx��Y�(��DUʻ��?߯ >m����n�)�Ly�9�v>�@;�f�?ٞ( ���s���3rOw�ـQtEU�ͫ���D%2�����x��X�s�-Z拰�f7#�h��@����;��Z�[4�YRSjdi�6(6��gcZ�X�k=�pk�lv�n9�SS���}������J1�7�H������;��Z�[4�٠{�&��S$JeUk �U�s�ТU@���=�׀}�2��?�anT9��H�������x�n�=x��Z� ���eMMʵE����$��BJ�~�x�߱`����B�P�T�w�;�Thy0p�Lb�h׬�;�k� �7x�n������L�L�98��{��{�@336�-a��=���z���������{��t�n��ػu�Y
���;�w���w�6� �׋ 8.��F�H)�Š��@=[� ��x�s�
L��jz�.��U]����wu�z�`��� w�����PQ�1�2G&�y�uV���w��")�wu�v&�)�%2D�6��@���h}l�[f��빠}���l�I2I$�H%�   �/\�[5@���\H�GR��v�Fy��f϶d6譃�l�2�=���a��[����k��3m���3,k����t���牲���0��N����������i���
̕t�wR������iŞ�F���Н� �M�Й��Ν�����g(N1io�q�����vl��g��>�Z5����;��w�}�|�<�s[`:浄�,6YR�ԕ����9Rn��C�q�9&
d��7��"n3�@/~�4ֻ�<���	/�T�p[�I�T��,��RM ��h^��v>�@;�f�g��t<�8d&1I4����Z�Q
d{�x����� �2c�4ԓ@���h�٠�� ��h��V�h�nD�J���� �D/�	B������w��7q�Z,���m�`��H0"b��h0�ؘ�禡�X�!��b-���a5��eڂ1�܌nI��� ��h��� �[4�-b�o��߾�ot� ��߄ءA.I$��Ʃ��ou�m�~S'�-WAjnf��ͪ����w*� ~n��f�{��}���sĤ!fM\�~���{{� ;�� {� ڦց�}�s`�SFd�)&�[l�/u��-�j���@�X�a[��[@<n�e������]jz�]ۗN66�t`y�M6?~���t�M�s�NGj�'���0-[n0�y�[o0>ˀ[FLy��f�n;V�_��[w�=׋9(�GGU\ԗD��M��� �� m��-J�(������I�4��@�GA��`2b�,P�	A?QB���_���C�i��
0 G��A:f}��nIޚ�n�}�gVȢ#����m�@��ـ6����Q3��y8
'����&�{��n;V�_��m�@�s�ե��h��@�I�I6.�A�a�TSG`�ní�2� y[��k|���m&okJd�Lq73�?�������@-��(������ذ��_�U��3j�n�����/��m���V���^P*|nnr��.7���[o0=���-�j�}l��v��0P�rQ7w��N��0�>� ����ľ�f��D�؈� <�Ȝ4�� ��� ���zu�e����A ��z�����]5-k�.%+1�q6r�>��ыg��a4堸�����������0$S��<���E�nF7$�[f�ď����-�?~�hV.
b�L2M�`{Ө��N� ��� ����D;��S$Jcp�;��4�[4�٠^빠�hG1�Īp�UV`�w�tDB�S��w����ٹ'�P�`Q��]{< ��  ^�.m6Miwiڲc���-�:ɧ���<�.��kh����	�;9{nJr�`{>z�o�y�C��u;F���	f����z��Y$�j�i�dy�Af`&Q�t��Lr�n��S��+�u6Ǚ�=8<�3���p跶���5̮�cz�ͩ�j:Mϟ]���^r����ӞI��c��$�՗Z�&�Me����P�
�)�{�]�����-سص���"3U9���S����u�
v�;�<u8۷gg�"\d�H��x�����>��4��M ��� �u��`��c�@��s@�Δ���@=m��@[D�i�&h�Қ~�h��@��s@;*���ҌNF�G�_[��o0,���e��]ӔDc1�ܓ@=m�v>�@/�� �}�V���ĲE�A)���v��Xi�k�t���
�{,V��M��4k�8hb�L�@��s@���h�٠����w���S$Jcq��>��ݻ�iF��UH���y�}�y��+L���f�Nd"p��@;�f�z�4�g�%��ۚ���}�p\�4�œ"$��>���V�-���`�n��8d��$�>v>�@=�� ��h�[��$���c�9�n��+�����i[zжֺ\*��.�!�"#iLAc�f�ݏ��u�@=m���s@;*���ҌN���� }��tD(���w^��,�U��έ�DF3���4��srO�}ݛ�A0����}��Z�[4��cQ	�H�`zJ�E�� �[��o0>��w���S$Jc#s4�}V�{���l�>��;��&�L72&݈����ʌ�U@v��o���c�!v^wJ���M��X�2LSs!�X�_ w���h�������e���.���X�i�ww0�������e���h{��1��
&1�4���ݏ��u�@=m��!%lDm+E+%Uլ�IKj�N y�^ |۽����j�DR��Q�;���\�%��8�Q������u�@��P�D����5�ŀn��8��S9EÊ�$�,�#]�l�cf�;6�OT�[C�tܜ��ij�m���w��w��M9ܵػ� ����0=%i�"�q�}-����@1Lj!?����s@���h�٠��׈��1D�H��Ի��n��8��xrJ"d�w^��f�{;-�1<ĪNb�h�٠[y��+L	ˌ/R�����*�r]��ͻ�9(����|j���f�3?��=gY$�I$�I$   M��y��.!���:��ێNzM��n*pi�Tg��<���L>�s�6_�k�77��#�YB:��7�i5��m�e���In�հъ�h��<S]��C���k[ j:��똫r�7nӔ��2��Sb�+&*;d��5�npf�Ҙ�[P7ݛ;���y��nC��>vۋ�,z�7n���uNx4��1�&��P��7�ֵ���:���u�v�8�Z��t �g�O^.��i���hT����&\�Ź�����0$[.0���>���"3-�.�f�Id����yO����$��y�M ���hw]� �+�SQ�1�.��`Ky�{���V�Y�u�{�Em�4F3�$���hv�X�����Q>}׀=L�-Ƣ�dNM����/�z�l���h�б6�<8���bqt�$:]pZ*t�GT���}����I�:ܛW<�W4a1D�H��Ԓg��]���u�@=���#��b�!��V��ͫ����f�����Y�6�`zJ��/W�}�e*65Ld$�h}l�=��a�B�-�� �� ��U#*��	�U�]]�����|��O��z�4�l�<�U��ئ4C4����m��>�� ���J�6��;���e5!Z�uIR;��lˎt����6�Wi=����C�ﻻ���`���1��$^ ����@-�4<�����U�(��cr`��=7���`Z�\`Iy�/�%�0��? �Q	���>���n>�s�� *`	�P�*'���]�ٸ�٠}i,0��S$Jcq�3@�V���]�z��(P���� 5��d��S$�f)�w[4޳@�۹�[���=��m��,Hōg[�v�O0E9�c[���\,��]�˚۳z��8w8�c$j ��$��oY�}m��-��hu�@>�챈lq�D�ꮮ�6�gD%
&N�O� � ���9v$����S ��ղ� ��`��[Z`{��M�7EU�ʵws������� ;�^��,В��J:"\ʷӀ࿛"��f7#"�h�f�oJh��޳@��+m̒D�6�s���2�
4汸�Gb�����[�c6n)�k�M�� �%0L��-�M�z� ��$�>�;�^ ���e�7*d�Lm6�[���z� ���-�M ��Y0x��1G�E�� o]��DD)��|`ʟN��Q�i�a?���&�[�h���n;V�[�h�g,��ljbQcI�4zS@��@-�h��!�r)�0>����B�eC�(�F����H��D��"@�A�X��,a��� �)BU�Afகt��EH:Rh��D"�D�F	������N��8�Aj�0�ł������&��i*�[q�tf��#�4��DdX�FJ$DHD(@"�a&�F� ����@E$H�B�!Q ԪH�v����3i�i�� t"E"�S?M��fff`   �         ��   �`            
����o(یO+UӡKh!dNi�hV���Ӵɤ��X�B�t�C����j��5U@uUW*�+�S�S�ۜ=��u���U�$]P�.����cvrb��Uei���;眝�;N�,E2W��=93^1��aV�s�5��=�=��r�m8��%is���W3�&-���X�L�Kb곞1�إi�v'>����&wV�FE.���56�u:��
vm�*�%CVm��F�c �j��CJ�rk0��]ˑ����@P��dl����΢ۧ^�̊�וk��0b��ȵ+�[`Im��m�=�nr ���
�Q0P���mWH����P��U]T��.�ɫ���_u{�8S��#<�ò�	';NEt��5�h�AR��
��b���M�M:8���>��"P;Z�ۗp��4�vL�+��3��&�����&�,IZ���ڪ{K��yP�峴��F�m\�!�8��]��'k���b�g�6���Vp��)���0J(b:mq\p�e%J%0C����"k�ölB�жL�4�s\��4�r R�oj����0��I4n�nUJ�tg`n�A΀�7h��A�������A�M�h�62�`��:�؇�
�Ɣ�g.�N�%���H�8kWr�6���v�@ h�r��Z*��k���}m�zZ;���M����Z������a�nm6y�=m,���(1 =��\�
���U*�WR�C�p�ih�[���\�q�k���n6�Z�U����vW��ն�m��S�Q&+�c	S���j�<�ݐ�oe1�%v�;$��Z�t�#��i:j���0ގ
2q�.,�Vgo]��)���fO��}���s����K���;2�l*��!���+M�,�U��(WQͩ�x	�yN�{���{�{�{��>�q@b�m<O��{���{�;����  Ѷ� �/��&�mv\C��:7A��ݱ�d��5m�7�m�1C\9�P5s.�(���J��~�v�荌�pT�+h�zv�n"�W(ַT�H�3pݸj�8�C ���kBs��*<�u��)���b[�Z��=���\v��U�vv�2�)�ûo0\ݎ��.����O+۝�P���58��G/S��3��T7�|�kZԲۙ�E��4C-���M���=gج�{Dt��Ok?����w��|�9P�5���ͷ�������f�[l�-��s�_�m(ʫ��j�� n���JL�wu��|`�ns�%2�����.�U�uw��׀n��3ܫ�p߿~�צ* �bS��@��L�M� |ۼ�B���w^���ajl�We)���0�Z� ��%>���߿~�wJh��*�'�I�C'Kz6�"vHl�
����,ݓ�r�&��Kێ����Lq��L�q��Z�l�^�@��M���h�J��M&:��ffnI9߻����̝��� �S���w���	)��S,�*��
Ф��~4�U��� ��4�ė;�51b�a4?D/�(�k;����׀=w�o�ـ��T��܂&G�w�� ��4�Jh�>�@�>��q䑦���Y�9*:u�p��1�k�h��65˴��򸉉�1���DF3���4׬�7[ŀo�k�_H�׀o;�� .yfr7Q���	-i�<�\`�� ��4^%�L �H<N7&h�?�w$�����Ȕ�؀#�$"*H�DK��wy�'>�vl���h�3V�Sjj��(J&w�� =ϯ �o�U�p��re��&���h�Y�^�s@��Zz٠[��m�Hp`�����Ԇ�Ff�h��k�/6��c<Fy;4����kƦ
Ф����s@��Zz٠�f��q%]�O��D��&��q�Yo0����֘���m(��0&I�^�h�Y�^�s@��Z���DF3�����>���Z`O-�b_��5�D�	E��� }��G 6�mH����x��s���$)!O>��_D�,K��}�ND�,K����M���t���\{7j���jζ�v6X�T��Nͫ�:D��WuՎ����bX�'~���9ı,K��ٴ�Kı/�wٴ�Kı>���iȖ%�b_���]L&�u�u2�.ӑ,KĽ｛NC��&�X���fӑ,K������"X�%�߳��ND�,K����9�WVa1�]ffm9ı,K���m9ı,O��p�r%��CQ5��]�"X�%�}����r%�bX��{'�&�5p�!�.fm9ı,O��p�r%�bX��;��Kı/{�fӑ,KĿ��fӑ,K������%��-5s�"X�%�߳��ND�,K���m9ı,K���m9ı,O��p�r%�bX�Q��ٙ�` .�   0���8UR�usӺe���L��:�g}&�#�S����l�n�q� �NTu���-���z3��P�&ۊ������#%ֻť��kZ�	Z���,zʴ���C'l�k���v��;./<��v}bzG�o
�tسU^� ���b����dy���<�i:1G<�U×�j\f����5�䄳Z&��jJ)�BCy�Y�J�ju��â.�7ap.#�v��&$��Z���Ӎ�z:-'jmkM�����Kı/���ͧ"X�%�{�ͧ"X�%����ND�,K�c��_��$)!N�}T\ܗE
���fm9ı,K���m9ı,O��p�r%�bX��;��Kı/{�fӑ,K���ޭ�Ԓe��&�L����Kı>���iȖ%�bw��ӑ,KĽ｛ND�,K��^B��$)!I͙�"��6�ʒ��a��Kı;�w�iȖ%�b^��ͧ"X�%�{�ͧ"X�����ND�,K�N�z�a4[�0���Yv��bX�%�}��r%�bX�����r%�bX�{���Kı���_��$)!KZ�ꪕ�T�
�t�I.��*5U1n�nP����x]q�H�{7n��Օ�������7���%���6��bX�'���m9ı,N����r%�bX����iȖ%�b_�%�Ԛ���\������Kı>�}�i��(��2&D�?��ܻND�,K���ٴ�Kı/�wٴ�Kı?k����%��-ԗ0�r%�bX��;��Kı/{�fӑ,KĿ��fӑ,K�����"X�%�{>�nf�njkY��32�9ılK��ٴ�Kı/�wٴ�Kı>���iȖ%�bw��ӑ,KĿw��ٗ,�MCZ��ֳ3iȖ%�b_��iȖ%�b}�{�ӑ,K����]�"X�%�{�{6��bX�%?}�}�iԚ��:Յ�[�%��r�V{Ip��:
��������U�<���p]��U�������ow���m9ı,N����r%�bX����iȖ%�b_��iȖ%�b~�f���\�ɢ���"X�%�߳��ND�,K���m9ı,K���m9ı,O��p�r%�bX��w��S	��a��\�˴�Kı/{�fӑ,KĿ��fӑ,��dDu��N(#�M���������Kı>�=�v��bX�'�羜�u�[��Yu����K��/�wٴ�Kı=�{�ӑ,K����]�"X�%�}�{6��bX�%��/d�I�M\%�j˙�ND�,K���m9ı,N����r%�bX����iȖ%�b_w�ͧ"X�%������n\��`qǧ5[
jZ6�ܩk��Ek��\"�Ѯt&��S�%�i�0�r%�bX��{�iȖ%�b_w�ͧ"X�%�}�{6��bX�'��p�r%�bX�Ӿ���kV榳2�ff]�"X�%�}�{6��bX�%�}��r%�bX���iȖ%�b{��]�"X�%�~����2�sR�Z�Թ�ͧ"X�%�}�{6��bX�'���6��`�%���v��bX�%�}��r%�bX�{�ճƭ�p�]kY�ND�,K��m9ı,Ow=��Kı/��ٴ�K���� ���L�}��r%�bX�}�d&%�2j�e�a��Kı=���ӑ,Kľ｛ND�,K���m9ı,Ow���KĻ�����?�~�w��vN[�^Y飞9R�J�8�Wm��W�ﳱx�a�t��It�_�{_o�L&�u�Yrff]��,Kľ���3iȖ%�b_}�fӑ,K��}�M�"X�%���}v��bX�'N���˭j�&�5����Kı/���iȖ%�b{���"X�%���}v��bX�%���m9ı,K��^��I�M\-�j��ͧ"X�%���ߦӑ,K��s��ND�D�,K��{6��bX�%���m9ı,O�����Ժ��R庙�ɴ�Kı=��ӑ,KĿ���iȖ%�b_}�fӑ,K�����iȖ%�b_N�z[��[���d$�̻ND�,K���ͧ"X�%�}�{6��bX�'���6��bX�'����r%�bX�:���ӻ��ou������ H   D�e����x�����2(*%v�t�+Bv`����N��m��8�m���uTF�y��$��A�`�㎎�d:��<7Td�<�{@�[�7;W]P^&g�'au���n.�9� ��x�������2�-��kL�1���6��k7h���ɇ�&��/;7S�''8������ƕ�E��g��<�~��5o�atkWF��.����r����+F��l�L�s�b�m�<c踐��_{�w���{��?���ͧ"X�%����6��bX�'����r%�bX����m9ı,O�ۻ=f��p�]kY�ND�,K��m9ı,Ow=��Kı/���r%�bX����i�"6%�b~�f���\�ɫ55�ͧ"X�%���v��bX�%����ND�,K���m9ı,O��siȖ%�b^�����u�Y�35�iȖ%�b_���iȖ%�b_w�ͧ"X�%��{�m9İ?ɨ������r%�bX�<�N\�֭�a��Y��ND�,K���m9ı,@_��siȖ%�b{��]�"X�%�w�ͧ"X�!����������VϠ|� y��N%�g5��gmp�%�O^#��#�"#kJ�Y�ul<�[��kW38$�H�w���A;��۱$BA���&�z%�b_w�ͧ"X�%���/���u5p��u.k6��bX�'����r�Ш~T���n%�w�{6��bX�%�}��r%�bX�}��m9A�,K�|w�ܹ�sSZ̄���iȖ%�b_�{ٴ�Kı/�wٴ�Kı>�w��Kı;�w�iȖ%�b^��_kS.5k�f�fӑ,KĿ��fӑ,K���ߦӑ,K����]�"X�%�w�ͧ"X�%��ݻ��Գ.᫢��ͧ"X�%��{�M�"X�%������ӑ,KĿ��fӑ,KĿ{�ͧ"X�%����>�����ٔ�5����Gg\\X��7��}Ȯ�1y4�ӷ`�[�',�\ɫ5.����%�bX��]�"X�%�w�ͧ"X�%�~�}�ND�,K﻿M�"X�%�~;}|ja0�2e�&fe�r%�bX����m9ı,K����r%�bX�w���r%�bX��=��@�,K㯏reֵnL����r%�bX��wٴ�Kı=�{�ӑ,h�'��h�(�F0� ����m�Gr�%!��p#!H��%	U"�R"T%H��R,�4� 4���:�H"j� U�b�!HT#X@ҡ(!(��c�`dhA��  �"�1�$1`�)�(��U�����: �Vh(��� O�VY�"�"���� H���D��`FXP���"X�RX�%"1��# ��5�Pڂ�P <�P�H�������,�X��DM�x�q9�o��Kı/�wٴ�Kı/���ײMh��ܦ\ֳ6��bX�'��p�r%�bX��=��Kı/��fӑ,KĿ{�ͧ"X�%��^��ٚ�SW
\�D��ӑ,K���ߦӑ,K� ��ٴ�Kı/��ٴ�Kı=�{�ӑ,K��O{V�V�5�kXf�fD��f�Y���r�/i��S"���P�ю���F)Br��o����7���{���fӑ,KĿ��fӑ,K�����"X�%��{�M�"X�%�~�wR�Z�p��]k2���r%�bX��}��r%�bX�{���Kı>�w��Kı/{�fӑ ı,O{�ճƭ�p�].fm9ı,O��p�r%�bX�w���r%�bX����iȖ%�b_���iȖ%�b~�w�3E�p̒���6��bX�'���6��bX�%�}��r%�bX��}��r%�`t�GH��"w���"X�%�~'��S	��k&h�3&ӑ,KĽ｛ND�,K���fӑ,K�����"X�%��{�M�"X�%����{Zְ�--9S��o	�Y�U���ku9m��FT�e�vٽX��8w3�.�T.�Ϫ�����7��,K���m9ı,O��p�r%�bX�w���r%�bX����iȖ%�b_ϯK�I�j�k)���fӑ,K�����"�ؖ%��{�M�"X�%�{�{6��bX�%��{6���'����w��������Ӈ%�0-�'"X�%��{�iȖ%�b^��ͧ"X�%�w�ͧ"X�%����ND�,K�|{�\�j��ֳ!-�ɴ�Kı/{�fӑ,KĿ��fӑ,K�����"X��Q;�s�m9ı,K��j_�je��u��s3iȖ%�b_���iȖ%�b}�{�ӑ,K���ߦӑ,KĽ｛ND�,K����ٙ�����   �Y��;5��P����� ��6����F��b�<���T����]�����c���۞ݦӥ�m����B�Ӈ3����V݇o��'�<�P%m��Y���9-[m�m����L�v��k&õ�s�����N��ʧ��m1�R)q��Z�{G(�$��t�v�нC�ݸ�%@N���k�v�а���[���V�탫�)&�Ö��7l�V�E���W���e��jP�!��"��w���d�?��{�ӑ,K���ߦӑ,KĽ｛ND�,K�｛ND�,K�{�y՗%�2MjKr�ND�,K��~�NEFı,K��ٴ�Kı/��ٴ�Kı>���iȖ%�b_��x��h�d�$�ɴ�Kı/{�fӑ,KĿ��fӑ,�a�������ND�,K����ӑ,K��|{ӗ.��p�u�s33iȖ%�b_���iȖ%�b}�{�ӑ,K���ߦӑ,K���m9ı,K���}�5�\.��5sZ��r%�bX�{���Kı>�w��Kı/{�fӑ,KĿ��f������ow��_����K�nH��d��
5he��Ol���ų�9F��i-zY�K���.[��Z�iȖ%�b}���iȖ%�b^��ͧ"X�%�w�ͧ"X�%����ND�,K�|{�\�j��ֳ!-�ɴ�Kı/{�fӐ��| U:�p ^"~�bX�9��m9ı,N����Kı>�w��Kı/���{Z�ˢ�u��s3iȖ%�b_���iȖ%�b{�ߦӑ,K���ߦӑ,Kľ�}�ND�,K���l�f\-�ZԹs3iȖ%�b{�ߦӑ,K��}�ND�,K���m9ı,K��ٴ�Kı?w�םYr\3$Ѣ��d�r%�bX���iȖ%�b%����r%�bX����iȖ%�b{�o�iȖ%�bt��~np-�nκ�9��Ա�DQ�:�aLݣ��v�ݳ[t��c��s��ͧ���r%�bX���iȖ%�b_w�ͧ"X�%�ｿM�"X�%����6��bX�'N�z��ֵn.�Nffm9ı,K��ٴ�Kı=����Kı=�{�ӑ,Kľ�}�N@ı/�Y�ڒ�W�f�\ֳ6��bX�'���m9ı,Ow���K��M����K���iȖ%�b_{�ͧ"X�%��^���Iu5p�˭d�Xm9ı,Ow���Kı/~��iȖ%�b_w�ͧ"X�%����ND�,K��=�.\Թ��̤-�6��bX�%�}��r%�bX�}�{6��bX�'���m9ı,Ow���Kı=�����$�V�ƴ��N�K����B:gjq����M�gd�.�����K��Cr�Y�ND�,K���m9ı,O��p�r%�bX���p�r%�bX����iȖ%�b}�l7�Z�.�jS.fm9ı,Ow���Kı?{���Kı/��fӑ,KĽ��ͧ �bX����ά�.�h�sW0�r%�bX���p�r%�bX����iȖ%�b^��fӑ,K��}�ND�,K�v�ŘMᬗ&kZ�iȖ%�b_w�ͧ"X�%�{�}�ND�,K���m9İ4
�@Ң>Ur��]��"X�%����ח.��p�u�s33iȖ%�b^��fӑ,K��A�������~�bX�'�����Kı/��fӑ.��ow����쫴�֜�e���ԜN^fj匽<�]p󣜽Aǀ��1q٧���N�Z�]k4j浙��Kı=����Kı?{���Kı/��fӑ,KĽ��ͧ"X�%��^'}���j�K�Z�5�6��bX�'�w�6��bX�%�{��r%�bX��wٴ�Kı?w=��U,KĽ���P��v���������oq��~~�ND�,K���6��bX�'���6��bX�'�w�6��bX�%��֟�t=(g4}��oq����~�����Kı=����Kı?{���K��f�k���ͧ"X�%���z��5�2�n֥˙�ND�,K�{~�ND�,K �{�6��bX�%�{��r%�bX����r%�g��s���ǻ�������p � `��̖v�XW\�m�.@Όà����m[��E|��݂��.��Q�b��P)���]h[�f�Ӄ���p񝣬��wN����ҧv5�(��zޮۥ6K�cV-L���	cN�Ê{�۞���W8��1�)J�<������$�q�QGgm�8fx���N\3����*�xṊ\.�X��T�.����L�I��k�]r-ϖ��L1kƬ�Qݹ$Ϊ]�V���n�/F,uճ�(��~�q��K�{�iȖ%�b_��fӑ,KĿ��a�
$�Q,K�g���r%�bX�����I��nɚ2�ɴ�Kı/��iȖ%�b_�wٴ�Kı=����Kı?}��m9ı:w�ח.��p�u�s33iȖ%�b_�wٴ�Kı=����K�E��j'����ӑ,KĿ���m9ı,K��=�.�p��h��k3iȖ%�b{�o�iȖ%�b~����r%�bX���iȖ%�b_�wٴ�Kı?k��V]M\)r�Yf�&ӑ,K���w��KİT��}�ND�,K���ͧ"X�%!v�q��!I
HRB�.}UUt���J��cgћ7euT5��\���Z���$�;�&���qN)BsQ�Z�{���oqľ�}�ND�,K���ͧ"X�%����]���Q,K���i�����~�E���C9�k�w�%�bX����m9�Ȉ~>� ���,Mw9��Kı>���Kı/��ٴ�Kı;��T�5�2�n֥˙�ND�,K�{~�ND�,K�s޻ND��,K��ٴ�Kı/��iȖ%�b~�_>���ѣY�Y6��bX�'��v��bX�%�{��r%�bX���ٴ�Kı=����Kı/�}�a4[��f���v��bX�%�{��r%�bX���ٴ�Kı=����Kı?w=��Kı/�{V��7�cK��Q���ً�5`�v�g��S�r��{i�۾���Ů>��v�\���r%�bX���ٴ�Kı?w=��Kı?}��m9ı,K�{��r%�bX���<{R]j�u�ѫ��fӑ,K���ߦӑ,K���w��Kı/��fӑ,KĿ��iȖ%�b~פ�,���R�ֲ۬6��bX�'﻿M�"X�%�}���ND�᠟��12H�$bA�J�K�O�"A2'�_��m9ı,O}��ND��oq�������P��v������,K��{6��bX�%��}�ND�,K��m9İ?�&�}�s�m����oq������N���AW�Ȗ%�b_�wٴ�Kı=���ӑ,K���w��Kı/���iȖ%�bS�}o���$�ˣ3M�Zպ�F�m�(Ea����/\�PSY76��*j�'�{�ڬ��SE�r����7���{���}�iȖ%�b~����r%�bX��{ٴ�Kı/���r%�bX���Ϭ�)�a4h�k5�ӑ,K���w��?�c���b_��fӑ,KĿw�ٴ�Kı=���ӑ,KĿ��I��nɚ2�ɴ�Kı/���iȖ%�b_�wٴ�K�E��j'����iȖ%�b}�o�m9ı,O���[�[���h�5�ͧ"X�(%�}�fӑ,K��{�ND�,K��ߦӑ,K����̉����ͧ"X�%�~��{��)p��寽���7���{�{�p�r%�bX��ﹴ�Kı/���iȖ%�b_�wٴ�Kı=�~��jۗWv{t弻H�5-���*Z�c���v��,�kf�K�!ku�6��bX�'��m9ı,K��ٴ�Kı/��� ��bX�'��p�r%�bX���{R�kV榳Yl�]fӑ,Kľ｛ND�,K���ͧ"X�%���ߦӑ,K���}ͧ" j��X���ֿ�52�˫&��-�fӑ,KĿw�ٴ�Kı=���ӑ,K���}ͧ"X�%�}���ND�,K����Y�pֵ.\��r%�b �����6��bX�'��m9ı,K��ٴ�K��A&�k���6��bX�'���?�\��0՚�j�ND�,K���6��bX��w�͉ �'��M�$�w�6$�H������aW��
���节�DT_�PU�AU������
 ���T"�� T T"�$���B* �@(�T"�P��P �*� P�DX@	T$P�@@� T AP��P��Q"P��T" 0B*#T"�P�*�B� T (1DX(�B
$AP�P�AP�P D�P��� T ,AP�$P�$AP��P�$T��P�AP��P��T��T  �B ��"�������������V��*�PT_�PU�EAU�aW��T_�PUЊ���EAU�ъ
�2��@�8��>�����y�?����G��5���4�@hTUuV˻wF�e"�{� 4�
��4  
 )E(   Ry� }�����@ j�nw^��)�������m����pI�Ѿ`�^�   t   � 4#�|}O���oh�4(����S�'լ�(4Q�ʫ��4ç�O]y��^�G�Hϣ_F����!��������������|>@���F󻢯�^�4Ѯ��98((и��F�\���}�HࠡG�x:
@�����h��{�aA�MC�p�PQ�C��	}Tǣ���D�ףA��ڇ�r:7�j�( �7;�+	ܫp�hd(7qz�wcG�B��_B��8+ѭ:5��<8k��N����D   �Pd���=OD���12d �E?���MI� 4     ��T�Mj�bb #!�@  �Ѫ�2��P���d��M b2d4!��Bi�44�<���&M�jMR"�H�  @   =)�����}#�G�:��G�J���ͭ~��l��a�fl�����\�6x_���u����j��l��9��:�^�3`|[m�Pf���o��c����.��_�}~����= y � ��o m��r��,ym����ym� �y�f�yp=�g��fyά-��l<�c�m��yϟ<�
��j�333����]����w}��������wwww���������������݋���������]���������]�˻���훻Wwww˻�www�����훻����wwwwwwww��wv���}wf�����������{�����www��Wwww�wn�y��hEi�_��(_��?�aKU��,��״.00+.���7VW#�i7��)n����A��]��!n���K���&<{�%�M&�`�I4��&�Y6�=��d��hy�؁̓����փAljJ�p��kcZ2��4}y�<�'��k�:b�&��΋��ףq�B�G�N�d(K�D�M)�ہ���25P���D	$�\��]1��55�n�Zd��6l	VC!��ɡ�"5)-��#ؐ�\�+4Zl��Bq�,���'��8�iݕq�q�	�*�TdW�۱���j��2�7�Q������l[Y��,#�227f��mki��-�6�C �@�t�
�l,�"��I��t����cHB�Ryf��=A��:0),�6�c�gZ4���5�ou*�0cE��-��;��Z0�``i֍�}���1�,%��:7�B��A�F΋:H�E��Y�aҐ�3[��,�e�,�Yxh�А�����z�f�Y�F��I
�z���%�����<��p��HՌa�%jM�E�f�"E QVI��[YFh(4�^��;z�{NZ�$�vpz{�!I`1�CR��]8U�
�4\��;-���L`�-�q�w8`&��ٶqu��������&��0�3�4¡]1�lz�1H�cAnӠ05��}��4����t�(�8�0 Sy0֘U�CF�z�z%^tl���m6Q�&��#@�2I�aF�aA��J�o���U�+�Oq(	GY]�tl�h�L-�)�����d-��4,[B�D����H���1B:v�
,�H����b4���R6���B0(�F�!W��Զ5�0��QN,B��čJ0�U��z7�ѭgI
�4��LaN�$M(j-6f��ޥ輋K�i6$Bݬ����8(��Z(���%�R������d^�c�4:G�8R(j�]�}L4֋	�Q5[vaE�	�\�F�ZГ��5���n:�rx���V�6j	7b��m'�z��V˕���q�f)�)�#�`B2^Q�jp(��J]
o4�X�[	W�	��Iٺ
�,�XA6�-�YɤB�f��p]��A����H����1 �%��Mdk��6��p�R�
YWz7S]�&��gD(��Pt�K��>:����XT)��!W�&��h�W�L�/GZ�o{��''#�(v�Ƶծ�N���ޟ#��/�4qHi�eg]V��Nu�&ccJ���Ӄ�7�]�*s@�
E��Zr�/��6�����̅Lt@��4��+F�%nIB@�#�, Yp��QdU��-��K���\�4�ȋ8�◂�1q^�^�!f�Cy��_8���P�oz�{�!�i�{!. Bna�{-�m�B|b�|=�-�#HG�0a)֒P[���$�]�HI�Z6��7�	p�U��\	(���f�!6��Yֈ]�GA�	[:�7*㎝���ٳv�w�U���m�J�l�D��
4��|'�W]�w9�|[Gv�z$ZnQ���8J�d�XQ��2��h�#	�U���t䑢�W/�@�@�:��;]@���ni:��֫M����"���f�R^�jU�C	DG����!6�)- @H���2k[sY�lAi����H��ʁ%[Aw6wSU۪��o.�&�Xñ�i Ti��Ȑq�[����8��m�!�M�#����4:ɐ�=�ptvz��B��t�4��,q�t����.�`¬,H4���V�·6h�AӴ��YFvnkR��`�K����w���h%�֌�͍Dh��,��-�
�!Y�/�B��W�6l�`�dp]���XQ��Eu�2�ѵ�����\���Ƌ���d�.Sn}K�V���@a�.��٥�YI���4��wTk����9:��۵࣫f�έ��:���NA�����)|Zm�6r\��g��3�+iF�i��K�z~��������'�<� k�YC�4H�?|������I$�@      ~�    m       6�	� m�l              ��                                                 .�:��1V"��Κ�Z�Jm�h���K�(�6ӱ��k�l[]m $n��L��?0J��
���VNj\:���vDʶ�jv�A'�@���ljޮH�m�6��IkT�[(
�l�ҙ*����M�z�-�� ��  m�l�Ұ�Ö�ķm�I��2�{U�[M�m,�l� � 8 � �6ؗ�y;U�@$�O m���F�Kn���H�v\�m[M�@ �	lm��ٶ�{2��U6�^U��7T�����s�� 	���⍪�KUAī@[J�̐p;v��m$ m�h�ݤZ �\p��J̀��[��I��$�8����L���QT�vt�<�J��Kc-�T� �`*�{.�W�T%u��@����b�t�����`"Z�];bō#FX� �T6åʪE� 8m�n�Ѷ�b�]�dk�hB7���  H8rCZ���H۲C���l����m���Iq��7e���Nn�ݲ�h�Ŵ lO��  �. TU`�`9�r-m ��I��li����m{o����M��h 	�l�� 6Ͱ�  ����Kk��[� pm�ۜ$m*�Ā���@	;m�,�H��z�m� Hm�m��-� m�� �b�m �ۯg�5��@ umA���N [@z�kV�Zݛ�m��m�m�I�@  ie�-�	mm��M��<Km��L	n�l%�P&�۴�M�6$� p9m�)�t��l�`����i�#�SO([��N�cWlݡV]��q9Ij���Y��mHH-�M�-�  ���  �6m��i06�  -����zR���Y����[}	  H�06� �;6Y,-Sm�j@�[lz��m:Tu��d���K�cvKu��i���ᶽ-�9 UR�g��a��ԁ+l�t l-�^��͋h�@ -� �`   �m���6CceZ��Ųt�kv��m�m����� M����m�����U�.v�j[]a�[@��H�p  �a 	26���U�Ym�m'����  Ut2t@Z��8{%���,J�1�^���[:�
٦ΒR洓m���d�� v�t6������   �jZs�l�s`$�z���wl6���9m�[���"NK(�}n��[ 0m�Z��x .�.q�--���6�,��V�j�`M�H��-�� 6����z�7_4�J �8Hu�{f�� �s�i�]i5�Kۀ�ޗ`9j���RY%ڪ��� ��}�I��-��$�ȶ^$� �V�f�����T�ʎU��� 8p�� �hҳm�k&��m�D�հt�� *�Jc, �M�X�����G�si.��7�8ڶ��NN�� m���q�m��TN9��Ԩ��T�-��m  �`  6Z��%wf��P�n��)j�Y��\   okw�ŭ�[q p e�6݀ ��[@ �.�m����e�n  u��  �kv��m�I�  I��L�$�m&��h     p���f��  �  �  ��h��   [@  ���hz�Ie�<��m6ض�� i 6�m��ڛU]�� ]��J�x9�YvM��O�۶� )%�<�N@m�`YgM�[,�I*��. �2m��m�� 6ٶ� hz�m�m�� p$m�-�趀 m   -�    m� �@�` $z��  m��   ����� p$ ��`��,�l  v�/Q'k���k�on�|�W�8`m��* �٤��'m��^�K;N���NF��  ���8�i�� /:�$[V�p�N�ki�sl  	�g�K&Ć�l CZ� ٶ��X���ͨ+i�\�tKu���M���N�l �����IUy�f�W�@U�L  ,�vH����J	 #��{�q�����㞱lH���nr� QsZ	Ű�ׄ�\�m��.��(���^y�� TU����APP�)A�?%����Gq�e�ՖV�sj�����9r�r���mO���s�n�+S\�-�-�u6��A	 ��ED�E~`#��TO����[B�p������6"h]�� �8��W��*lJ � 4�W����-()�@�i��P�{Aڥ"i4+�C`t�����'B�\Q8 R�@�h��F	�����K;MZv��*!�w��4��b P:G�
�@҃�Q��B��͕����&�؄$�#�*�U�т�-����C� � I�b�Gj!jZ�%�p�,z-@` ꁮ����m��m��m��m�UW*
������ʪ���������������򪪪�����<����������*���������ʪ���������򪪪��]��Tj��>� �"���⅏�w�Z����9�}�����x�˪�b�Cz�@
R$�1E �ˢ�B�� ���JY����!���O��jR�4<&�����UWm� �f�@ ��        �^��l�Y)b �aڲw3��b�V
�`*M��(�l7a*gt&�e7nҰ��f1(�V�;��jB�J�=�`6�w�Ȳ�Κ�#��ȅm�3�\v��U��`Ņѵ�m�� �ަ4.�7��l��B(Y;`�N� �5aÙ��%�mt<{>�#����eΗ���n�n�=������l���+Ǜ�e���u8�+Ǫ.Ζ�҅�z;Z�e���yW�d+V���;:��AL�e\�<oW9;si�[U͚�l��f6z�F� X����e�c9�L���/��l#���ll�����^�.uY�s��w^U�ځ65������[*��:�Z,�8��M��v=Q+fikjWf͎�Sf�3)3�׮l�U��d����t�am�)Z�:�Э��ԧt��j��쨭m��s�&�Jen��Y�*�p%sGF�����k�`STh�MQF]�cUU��^��'�- SJ�4�'j��h�v��)5�����6� 7&��{K�]\�tdg�M�tf�3�QN5�r��nx�ɲj�\�;Pd��3]�=��"rx��;;Y�$Ƴ&)�N��8��l��@�v������g����wn�*�--�B�8ܨ�G�񲣜/��?�N:���=�?�P��3:ƿ�eޑl���냼��X�e�=�c
-Uݰ;ޱdw�+\�!P�n�m��u����2��{b�����C[!�hC.����:x�:��m�z`�QF�Wlk����d;{Q�ˣ.�G9���M�#�@4�� ��v�����^_	���Q�n���b��^�ﱔÉ�Y���.���X�Y��Ɉ�7��7�Y�`Y�~�z��4��,�lۍ2CDS���8IH71���ݺ�v��
�s�o�X�%�V��pһ,]�%k��q��
-V�-�� �uwn��r(���kWl^�؈��V@r�h�c,��/���uf�ۮ]�	0� �̄��j�+G��2��H2�8�:��\4�ػ����L(���-틻`]���;�"�0#[�c�㡙�Vj��Z�&]���r����j�����QРP i,`sV0H�
'Ywp�nػ6�
��e��&�[	P��u1�� 6�v���^�}�{����Ʒ��(�f���9*�ˡ8�����4�GC�a�;���f��ph��2�u˷\4��M�t����ª�@��>�o��G������x�;5�<�nw�:SI]�ӧ����Њ0 �\�mI����sơ�Pc%q�l�lZmկ:�gX�x�`�zp���I�ءj��9J�����8Y;2�ֲ�5J����E����窃s@F�W�l�+��4���c�#v��ى���Z�-����T+���=݂��8V�$˩�J<�,aQ"'9���<�C;��U�\��9`�@Z�*�y�X.��\����+*��{�Q�9`�9ݨ�|�(��˲d�9`���;�^@\95�J�]�4�ͳY���ϪN�z�"d��˗���y�X/]��/ -w�Q��8V\˗Y`��,�vA-b(S���Z�:��pS�N��%�2�@�����y�X.s�Q�U�}�ܙPCТ�:���{���]�/��µ�&]Lҏ\�����`Ua�f:�]�4�d��-��"H����w]u��1..�eV�`��,�\��\�}r�&R��� DK�V��Z/�wj:�}e�]e�V@^��Q�]X���s�`������.f]J�(�^��ǐR@^_Q��8V\˗Y`��v�@��+��Ü�^h�빒�����v@q���k��.^fW&U��W�Q�9`��V������K�&H�^Z�[��|��S�
Dk·ԓ/����}X/���λ8fUaFU���/P���w]�!�v����V+@����ڏ9�E�:��u�VK/�����)n�G=8==L)�yys.e�2TQ��j9�V��uh���޹�˙�US4��r��!�S�r�|�� 7�X�"nV��˘\���;�^�//�j<�-�I�u�0��2�@�����/9���wc�Dߪ�;�K�2�/�yj=o��ά�׉��/�$Q� ����#a-Jfc9B
YwQnc�5h�����{p^3�WLm$#�W��z^8C;7O��q��Z��M-�&�&�*V�j`F^�j�(A�+���������w�]�����D�-��d �+��U�e^I2�%mG����V����]�Lʬ+*�pS�����j<�,z��	�VUi�Wy��s��uj:��ˆ\˹���뮬���E��7yrfUV^�y�X/]�`���߽�;ߣ׶T	dR�V�8��e�gV\9�Í]'w�~���-�-G���s}s*ref�y �#Ђ�	}uh�Nn�y}uB�.gt�d�@��c���U��< /3�krL�U�Q�9`���`����ZE']�C2�ʰ^s���r�y�Z/�N����ʼ$��� �-��c3�Pf&љK�􆻘a3
��/���Q��,���u��Xe̻�u�X*P�}�/�r�|���7ys2����r�z�b�*���{{���zֹ}��{���{�w�}��.P"�VԬZ�[[ZZP�KZ�I-ng�:���u��P�zQ�X@i���0"��
�#q�+-�4]�"	fD(@����U��)�~p��()�=*��t@H'Ib;G� ��`�������
�	~r�=��FϾ�Q��Q�4@�@��!�:P��!~yh9<��ȯ�N��aW&�5z�9����Bk���)�[��y��Y��S)�e2�D�K�A$A$ྃ�;�Ù�s���6�2�-�����)�qtz�t	�'@�t	�e2�&S)��el�S)��2�L��g���}��L�S$�e2�L�S)��d�L�S)��e2�L�����)��el�S)��d�L�S)��e2�L�)��e3����L�S)�e2�L�S)��e2L�S)���L�S)�q�S)��e2�L�S$�e2�L�S)��d�L�S)�z��w�.��e2�L�I��e2�L�S)��2�[)��e2�S)�y�n�L�S)���L�S$�e2�L�S)��d�L�S)�__]��e2�L�)��e2�L�S)��L�S)��e2�L�2�L�S)��e2�&S+e2�L�S)��2�L�S:���e2�L�I��el��nL�S)��2�L�PL�A$A$o�=T̪�4�e2�L�S+e2�I��e2�L�S)��2�L�S>��}��e2�L�)��e2�L�S)�e2�L�)��e2���L�S)��e2�L�)��e2�L�S)�e2�[)�}}��)��e2L�S)��e2�L���S)��e2�L�S<����)��el�S)��d�[)��e2�L�S$�e2�L�������|���e2�-��e2�L�S)��2�L�S)��e2��e2�L�S)��e2L�S)��e2�L�I��e2�׿��e2�L�I��e2�[)���L�)��e2�L�S)�y�n�L�S)��e2�L�ڙL�S)��em��y��}�y���Ke2�L�w���L�S)��e2�L�S)��e2�L�S+e2�L�}}|�zw��]w�L�S)��e2�L�S)��e2�L�S)��e2�L����l�S)���L�S$�e2�L�S)��e2�X�� ���U|󖢯�E^^J�r�VB�S,��a�h�z��L��3�@�t��N��e2�L�S)��e2�L�S)��e3�<�S)��g�8�el�S)��e2�L�S)��e2�L�|�w�s)��e2�L�S)��e2�L�S)��e2�L�S<�L�S)��e2�L�S)��e2�L�S)��e2�מw�)��e2�L�S)��em���e2�L�S)��bA5]�ʬ/.Ue�I�I�I�S)��e2�L�S)��e2�L�S)�y�}��L�S)��e2�L�V�e2��͍�חL�y����^L+$�� � ��h<�-���<��ח��Y& ��-�(@�}wh>y�1ȃ�V�$�3B<�-���
�@Uڠ+�X�h�wR	$�I$��ӝ���^��ƶ�ӡ֟75n�f�靔�.	-�h�/[S�� &ۦ���/4a|;���c�%(�fa�
�����M��ΤFv�Ad���s:ww�<<B��-VP�롳CL��!�.�z7f�k+t�ߏ�V��	��(����'�$�++J>@]n�y�X/��y�(�~w0���,�)G[Ձ���,\��s�����+/J>y�y �|�nw�*���Ua`�y��y�Q�5�N�>ϯz͵��{[N����֦�{UGglj�*|��I�w�Q�9i�"��=z��w;�|��$��*z���%(y�,~�-G�S�@���[�I�UY�"TJ����_b#����9�Lʬ+*�|���$���(�5�|��3�ZQ�@���J<�,���sP�uf[y%��\<8���)�4�Q.��ˬ�^�J9��/9�Q�����ax\��O ���9j>@^y(� ��Uayr����-G���i@3�:ECH��Q��\��k}_��d��j�V�q�b�l��Yl�e]��m� s �WXw��Ē$�HJ@G�vzو��z����ȝ�u�u�8Fb�n��3��c��л�Z�:m�E��[�v���ַbjWh=��ݱ�7T�<w����b:�:�z��C�zuq �I�!�#9�n3.�8/j��h�(e(�����C3f�oF#Zoh�Dr�ַ|m6P0hݡ����X�k���ɉHt.�:�z��Uک,ؑ)J ����Y�fc��=��n�  N�4�����4μ���q��W���	P�۫D��lj!���nF\�1����Lq-�[n��i�WP�+6�� h��e��*ٕ����SW.�Pj�����n'�~��3�x_<Ί����ł�����2Ѡ2Tetx�G8��au���[� ���V�
\��c;͸ˌ���̕*���k1{x�2�uwlp��v����Q�����Ρ��/�,�B�>�6��fX.�+E&� �
pԍ&�0���9�J��3��X��R3���P j�̐x׼����@�`]�c�|b3%Me�0�ha���n�􊽿A��H�Ux����{���U�<�(� J4���&䰛��m���.q�������X�Wh3��P8JG*��xP�xk�B��K��?�f)�f���
��U
�Oz:���{�i6Q��Cz۫�b�vZ:HF�ݺ�ző�Y�h��G"!��-V��*�i�F�.�4�R�D�������fc�k��Zoh]۫�cZ݈ ����	����,ӝը���4.����,���Q�/e���ϐ���{�=�˷q������Vqc��3`��5"H���0(�Z�h:;?&�Q��S`�m�uwn��q�2��O7�W�b����v8hš��]�X�Wk�8!�S���c���U{ޕ�ݜ��a$oh]۫��s��^�o{�����}�}��}������ E�`H�H�B0.�,�u �"P�8��s\\�p�X涢�79Wsw��|��&��.E1 0J	@i0"MڮbL[kZ�M!s�6���m�'ksZ����/n�gzŴH��wE]0�ȄV$N9����k�ŶX�kh\��GX�V\�뛡u�7��J�2��3ذX�Aڗ
������  ���6�$            S%���Za։��� hl��3���.m���q������V�"������Jl�LP���B#�D��	���/i��Z�ET�GGM��<�ڠûer��@�6*�n*��<\��&Jk|�Ls��&��YJ`�(-�*�H��vxL�Z�ۜ�#�f_*�b�*�j� Y
�L��U�
h
��2v�p��dvP����0)wMؖN�ڮ�{,\bW\l�G�aYZ(�6,Z��]�cf�c7��b�or8z⧳�8�n9u=�
˰^Z=YF��Ũ`��:�����V7=����u$	�����-�6��j*N',˻([NpV�D��+�=%چ��/IpEmu�u�YZy�r�4;r�c����4���/]��5�v��3���+r�/s�]:(�����.�o�ħU*�\�^�eJ&ծ��^qvI�z3���b�O�j� xz>B)����W�ɕ�������U\sn.أ��m*���,[���M�pn�!È�!�qt�Ė� ��nJ��O#���/[��n�Q1�]���v&i<�WR����</+\$�Uػ:�
Zk�{��n�
��=�2�b�-������f���ڌ����îq��m1d��FT�����!��c�3��d1���m��T(���`z���Q���P��ǈ��f`uwn����[(��7����=�,���@X�MҖk�dZ��5�&�0A�fc#��Y����É�ݿ�-A􁘆f�� oyg� Qha{C/]���&FDU��C\��d� *��=Σ�DN���[�X�8Go�M��b0����E��]|K�kͅ�m)��v��3��+7�ȣ1���5�.��ݿPk�|��:<���=�
@=O�����׬�t`fh{1����f�ni�tv�1:q1�8�h]ۮt��YR���ր��c�M��1��n 2�������*�$��v		��5�P�sr��@o��cq��.����^4�b�*�#!��e� ]��:(
��R����8�1M oh]۫�cVv��C�"SD�SO�op<\���c��~?��g}x{�s�u�y� >��؊"�л���]��b����N9�3 f!wn���b Qh+\5�!w�<r��d%F� f!7�ݱd�l`٠M s��  ��۝d�F�Y1����[�-��6�Q�lU�x^�j���v���~����^�F�w%܏G[n�99M[�͗��%��l�d��Q�k��w�7�����m[�.Mb�Fqыb���k�]0Fd�.���%r폈����2�nJ���UP��<G��=�0=�y�EQM 틻ub���sYl�4b��x
����؊&�f:�zŐ.б�/e��[X�eD���0$��H�4�DÉ�ݱ�Xs��SWg1@���?ʪ��]��u3�*��s�z���@{�M퍟{χD
�݈̑E�=V���X�^�������ce��f1���wn�N��m�M�����C�������&#!J=��q�u��	����iW���7�^������f�ݺ�z��(
��Pz�?|ƴ>�!'__θC31�P��32x���pC-l������Ϛ>��3{!�\Ժ\W]�k@��ͭي�v��ݏ����Vi�Ո̑E���eJ����	����d1����u�]�.���d�YY�����9g�v"��\��[���ții����Y���f�UB{��Q*��\pP#�۟F��z@�LA-�{λ޺�Wh>ٸ�L8�]��'����Z՛�a��͚����31�U�c0Bdd�Y�M��ݺ�NwV�H�3B��o�|"Έ���/��I���~�  �k]�Â�F邆W0uC4�C���.���6ńί�r7h����e�-���C�s�G2�9�VzٮDwѾn>[9�j�	�y�P�֋+����6�;d�N��#(�f5�].I��cM��_�놽�]���vɐ��Y�m�uwn�g{m-#Y��7�S1՚v/Cb&!л�]�]Y�f!�xx؉Ӊ:�
�b��Y�w1��*�������ʋl6�fJ�K�ǮըH$�l��([�5�������0̹2<�{���DFA�����Xi��̑�wn�޺�Wk�:����i�s2WMf!���[]�d)D&���m�uwl@o���$����$97D���q_y�I�V��yV��d{���P���x{��E:��w�uf��}�q��.7Wv�pzr������s�����z�����{��8E'%\�!5Z�Uj-�#�^Z\ֶ����t�[!/�yo���X��f�]���'��q@��T#
���НA�3��-95�C���qdB$�-I:���̴5�Ҵ@�
c�.")b*�x���@�@��e�U:~J��!�wߺ��ռ{����+�U�Z�v���ַb$d�WhM퍛�vF� [¹������*���nP.7^�n�]�[��}�u����ά�d1��5���F�bz.�[]�d)�4��-�u�����l�"<}�87�^����5F�#! H��+�z�S��V4w����5v�=V��	&ڀE�(��&�ePB\�aE�7L������Wkf:���b���a[B��vXַb$f"F�49�Yx�>�]H\��h��̕�۬<#1	իfCeGW|��	�|�O^�[� v8�(R��:�|���?` �:�K��=[6m��\&ż����d����5��n/c2�4�E讍�����b_�F��WK��]���I�����C<g��[D�wPw,�e�f�����N�37�ڽ�E�l�	X�d�P��"։���sU��������{���e#^���{�uf���؊`:v��5v��2c
)Wv�GMf!�����F�-U����t�I���}|>�ڛei*#6���e��B�h�s]����>Y���v��>�X��B��g�~�\lg<��_q}` �׾fCQ���@OH���5�xL�(�lY�\��c�T}�>��}����>#���^��Y� �[�Ml�9���9�m`�^�r9$��`J�r�۬5��΋��*��WMf!�����F�p-9n��J������$J ��
旝k{�5�t���k�Bkn��Ց��^��B��v7��|�%a�j��'����1���.u݉���Y6䑲d��cj7Wv��᫿�k1���Vx�!HE5^5��fJ��Z���i���^!��ׅ{�VmU����1t3:��:�����b�����2Ww�x�^c��[��1(�&H�D�UЗ��l'S����'�g>q��u3��( ��]�5�Wv��>�X��3B��o�uf��g�j#n2�]ۮ�C�n�[�d)�O#���s��G,���a#$�*i��A�����=|s�;��  ,ݴ۲^�ڴ�M:\8�	��9���4s,�<��3��[c�ܳ�(�	ƾ������v�G��;u��>;vݞ��FL�\��9�+� Wd�sTѺ85m�?}:G�y��[/��m��[���W��,���_#M��k�Л�����Fg!��P(�7x�UQ�u��w�#&"R���]�wn����D��Ug�o�fc�s1�g:��FL5����Wv��&E�̅	np\ŧ78ѵ�ݲx���Ќ��������U@���=�FC*:���Ъ� a�c�~������R�C��Z����l]~}�I���� �!��׽�%�Kf��%�C3#?
�/5^�y�P�\�ڶ�H4�l��젒?U *&&�����`��B��k]�����P��Y��3` K��PHc&�/g5����(P�T&w�-�n��F\��3G�=z��\�Xk1yv��4ێ��T(���Dř���� ��a�l�p@ۍ#1��y)*�meW�R���:[�̅(��$�D���9�!&��$�~˸�ei��V�UT4(
�u�	?}��,䎎�P8��9���&�r��T�'
$��2EE;�O@"H��kY��rT�y*Op�V�W�T}�I:��E�=NI�UP�\,������BOp���t�,��B])��U�F�=7U�i2�:$�(���5�NfN�UZD�(��g5Q�!0蓙�}^ U
l�2BM�I>*��mig�R&ڏD�{�OJ6P#�9�!&�FB�Q�P�	x�I�D�̐�UA{��$���dI�R�;1#�;ޤ�G�􄓖�&Ws���{��w��{Ξ���{��wd�@���RDWj���A|(�@�����׾c�zi�P������;`17*�TTSTJ*�j��I�ZF�V���i�8'�|���He�X��d��K�-�w������� m�	m            ۫k�fv��t�jmWg�S0[�^˨f�9�u�J\��K�f�g��wX��V��f�p��OCn`��u��0�f�sv�����p�=���lplm:�����0��*���ۻXܼs`:��X�����60�,L�X��{
3�7K����$`nx�;�h�*���x�e� ��Rٗj�T6g]�*�T2ܱŔL^��,T��#N;	�dث��F�\�J��`�.m�є�,j�!��Ŧ)Nȁ�1��s�m�O:Zkt��Mcv�����BK6*¹1�ƍ%�l�A���^�m��t��ř<H3�ks/I�k��R+���4��+�����Y��-9mu�bm�I�=PP�+����.�l�m���,�Pl�Y`��9h&�嶖�W,�66Zխ������%q�IK仺l�Fq{u�ڵn8[�XY[�>�,� 2��=	az�A��	nwb������_W�~/����6�k��<�J_ӧ��e�|	K��hT%��u�}��Ab@��|�>*'�*%(�(6��>�D��jwy�O;ϙ�[��Ӏ ��9cvɵpJ��U6�Mխn�l�C:�0L��z�w!e��!�L�ҋ��9Pe��bd�&y׍�ݡ�44����^ؓU,���0Qs[v4��$�$�τS�7<��Gݞ�X`gF+��wqE<�CF��?�@�;!$�r� 4I30f�����9�!$�:h��s2L H���E�=N�'es2BK��h��]�H�A蜠+$�|����` �KZ�sb3$&s2BN��	'D���}�v�k-�\mmS�G6f����>N�/��V��V���N�$�(����D����d)j���7$�J������{�R���u���vBI���]ě(�q|Q'���{λ�u�[��F���>��/��F��>4�p8X1h`�u���f1�s2(!	j��AA�u�q#�(�P8���j��� C��s߄E�f�Ʀ��f:�X���2䩓P��<îr�p�\U��Q� 1q�<k�Dd����;��U��5���IE�v놻��N�o3���x���;^3i��R�iR"f' B$�I�V�+�[����]��4v��8�]��]���*�#�0>�!�����Xj�� ���@�uwN��<��>�"����О�ُ~�'���2�D�ػ���P�+XW4Qݦ��]��W#�<�vC�7^����r#������^�4���$RH��ݿUP� !x��׽����EQGWj�G�P�
{<ǽ�^��w�ein�5�m�x{�J��b�:��*2b5���a�_��
���m�  d�N�9u�`��Y�	ZX�@��@Kl�mA&��D2!nM6q�f^��ņ�]sA��i.;v�G3� ���ŉ�3�%�����9ŒYC�#v\MX8�s�t�s���$���������h-qk��ːA(��k@ \�z�Nǽ�S�Y������o3��.7^��8k3��� ��|�f�Mm��b����L�FUU��o��1YB/4o	��Қ��� ;n��f1�23$�k4`�l<���1*T�fCI���	٫���h{�u���|�l�-����UT \����*��@�l�%��f>��a����,Ŧs3%]��]�xF��b���1V�fcv�}<�QbTn�HHL�!A�f�M{h�vѺ,�WϢ{;|��uv���j��"0�ݿ������:��
��z>�2�SC���;k� h >�	�����^�$��yT5����T �{ҽ����Q�V��Gƹ�1��WhK:m=�M����(6䊋IHi9B�n�Q��9�:��5�,=�1h]���C��^��L�#P8�f*�����u��r�EA�Ykl]��Ӡ y�ng`P9��-��P˽W���p�{���&LB؛%�]�։0�ȸ��$��Қ�냪����m+�IEf*��m��~#9���cein�kz����γg��P(����'y�Y�}T(W=��,š����	�Wv��0+�9!Q� ����$�K8�-�-!�gr��@��[���v(�4h���ݮE��ڣ���.���u��˪Ԧe��,��1�
s�LR�ׁ䛪�+
���E���Kӧ�E�z�ͮ��GmQ��%���N�[�!��7�\5���9�낇����"!j��( C���Y��u�r�k3�8�1U�\�+&3AM�uΪ�����8}Ի�E��yV�fcv�u��[-��%ԁ�	��-�)�$' �_��4�oO��*�����]�E��$���8*�� Я����m׺���������2�2U��T�Y��]�E��bxk3� y�;�]̙ׄ�f�#�
�w�f���\���!{�B���TeF�����l :�;�����Wqfc�f*�J�l��m)�woP�#���37q+�IEf�n!�aU]�����n��{��w��{���3�=�?n�n��U�5�!
YA
	E2���Tś|����_��﬑e�M2�W:�Vg)���̫n���SIk-�ŔKV�Z�i�Cn�*���9D%%4��,"BPSP��H�[��;��?_�(�)7���%�<%4��'���ފz���e%�a8��$ѨT��M�Ɏ�&�P�kn�<�E=��V����ۣ=If4��U�M�T+~�=��(z�(4��> ��Tڀ|~G�:���v����pq�ޞ��(
���7�1�y�b���I��5wl��U
�oců8v|j���U�Ո��V�r�3�֤q!N0�b5�f:�UY�B�31��_8��(�fu�[�.��U
 ��pH[&hl�o�fc��$���1a��AI�Y�����=�`�tm3�<<Z�#��4;���5wn���P���.��a*�cXe�UJ5��KT4�+3t�cv���~�h����T'����f ��=��Q��9�p��U b���a��Z��Ude
�G3�Wx�&F\N��@ {�cc��{�s��`�� gJ��tkJ��GzϤ�m�3�x���g���m�&���SD
�˃vX7,u����@����uQ���N�
�\��2�B��\��Wl��a�+�KM-v�o�ݒo<]I�����.���̫  ���$�y"�q��&�ǽ�P#1k9�%5�����9��¨
�@5�牌�҇B��8OV<k/�%xb�(�@Q��p�f1���{��.4���a�UU��{�C���V�>#"p%)��1��I�[4BgE_�6gy-Ҵ�1���R�f�tL���Dt;}��!T*���@!����u��a���Vb��� ��� ��[����г���1����
s��JBMfc��a�3@��q4BD�m*���T�������m໷\�> 31��m^�J(�1V�gq��yUDg9��\i$���Ʒ���ԏ�:ߐd{Oh�Dv�{��a����,�5��oժͪ��3h��P���Fᱍh���B�c(޴c&@cr�l�f1wn���ѐ�:6pP ��;��K�޽Ȍq'	#����X� 4��0�K5�F3U���|��y����{Zp
��l}��Q �����Y��31�w���0S�7d��mb4l#d�B��h����x����?}��D{�xi�D�e�{޸7κ����D�	����\�5�ۮ����5*�V�]�v�Z�-
��U���v�������I��}�  S7o5��	lu�T;a�^j����	v�\̨<]�����<��aW7�J�g7��ЫZ�	���Ɗ���0���nݩ������aS,`gZ,�S���6���7P�ۊ��p"��7`��B�RI��g1�뎲�Y�}գ�4���ˮuU���;��f6�2?ZG��@��c����>��4T[�޶�f1�s�gl��}�z�a��}�yх�l݅��-�+��D��ƒP8,��.��z��]۩�؁�jU�?��^�����Z�yP5Vjkl]�7ho[�Lq&!
���>����x���#��4.��UY��c�Wv�Ln$Њ�A��0�T΅f�uiq��
.�~�z*�ݓv��~�+An��������9�B3��6\F�1�o�~   ?yT5~���8�Z�:�UY��w]�ԫ�?z����y������<���t�uN���I��r3pG!2 3Uv�\��<�@��7��F8��^1���1�P� ��#�����S��<@��/E^�%f$F�]��W���y�Vw����E==�Ʀ��s{1���i�Rt�<�ݻ8�����r �j����$�q��5�:�ʡA��h�<E�fdݪ�Y��T �w�A �J�3���.��[�,��d��� �Z���=@P ��oYȌq&� fc�]��a���`�TחI'�~?~�{����{����I�� Ih�MS
�TT��P���DzL0O�	�"1a�W!x�H��#�b�e��ɹ-�gX8g�;w�GI+"i��htNs��7M5�q8G4Z�s��5V[oNg1b��,L-%��0�9�B���&��S}�$���]�Y��ix^}>��ߏ� � �            �t�v^��[��BpV��lϳ�We����)=%�����D�[�	{u7\g[��\���a�jr�@M��,�r
ꬁ�����.ڧT��-u���¡�Q���:@�(]*��/�7b����m�1������@ٮ6�b̢��j6��
��P(6�{��[�� b	�P��V�ҩ���AI���B
@5�n�j�-ō��JNqڶ3gV�]n�<�-qV�%]�AL��K�U!�
n��c 
���q-�[$Ȱצ�W��x0������l6@6�z�[��<�-[�ܯ�Z˰� �۴qA���A����f���ex���Ѻv-q���}�
�	C�����	R��T[[h�P���e������F���ż�$�[�qY���lU:A�Uy����N*7Mմj����H�=�1D��Э��Z:ɴ�@!�Q��v�XN ��Ы3�*�\X#�~��{�z����� د�P)_P���T8 ��M�$\�H�I"��i���hP�l�hk�t�9��e�v1�V��d3	q�����WF��*���P;�wP��<��ѝ;�SBc[���'<��h�v�5��6ˮҬk�;�1���]	��6J��$6QY�V孛9��j��|��uU��B�  C��Ş-�
h�^򭚻�/�^P ������P��x�7���y������)�&�cz㫴2�Q��h�<E�f:�Ua��9ez�{�-���s�M�na� q�������R���J�wn���&2�&j��
c}��cǞ���b1Ę������Y��һգ����ݺ�UY�� �bp��<�m�V�Ԅf*����3~����I ��8�kp��[���5 M�\�I���+K�ƹ�1��uv�"^�	0�f�����d��a���K�1��3:��M����j@��PJ���8d�u�U����?UP�>��ڮw��c*4,�ַ�31�bUSD7�X�N4��әmd;mш���h(�PCY�Ʒ�Y���XG����Қ��wTGmV���u���)��0*�����ǽ�^��}a(
��|kz����:*��O�Cdk��'J#^������U��Iց����Q��NF�^/d��֣6�f��O~��;ݺ����8k7x$���9��36�Vs'�4�;�x"*5^55��}�J���^�c�A{�c[㫴0Q�R�	���l�431׀��۬5��|��Uw}{�O����}�Q� ��B\�Okv��1v��'e��v��h3L��6o dg�[p1�E�G�|{vw�Q\�嵅.pzL��^����|2'0�j�v�]�m��+��2���5��99rvI��Nܻ�<��N .B�NBӁ&���U�_}�� ��Y�w���-׍o[c3{1�;�131�o�tU�Xk�07�cQhfc��U��s0�5��1 QJ�U�W�b���<�O~����
9+.���4�\�X �s�F��;�Ϟ������k[�qF�5������Xie���Қ����;k�TF�c�i��Q�sp��31���e��(i�Z'Ā;�����B����q`�,�7W�p����Vb]�]��9�:�Uf�r�{���̐ �۬5��	���!��[ �v�%P�i�P{�}#|�P%SCb��[���Y�j���pGf��?
�7��Y���*�N�&ɉ���6SIHBpkAc2����o+uv���:�U��Y��u��jB�Q�b�J�f0s2xP�#��߰%	+An�5�����}z�����S">����2�����rH���"�<�z.�&f]V��c��V��.�ixcP��r�67�W=m�Մ\�c��%��C���f�1��u���c)@a�Y���wn��*��[�Lq6a��c[��Vi_uj&�iM�uΪ�0PfH5���)5f*�U���g]x��?7|�  vi�[�^��GH(��WmTrm�\��R�e䵤�q�[���ܻ<���OQ�F��s�vf����!B�l�]!�5�
��n� g�HV9��Z�r�\����s��XHx�Tk����ܗ�$�%�V����������� x�#6�
`�Mfc��u�b�5ܘ�1��.��z��P$�fc5�C�Vb��Eݱwn� ���Ȓ��Uڬ@o��Y�J|�g�=6T�Q-��Q\��`�1��p�&Z�6�����9�u�\#;��D�m)�wo�Uڡ�g�hֽ��( �^��!I�%f/{�c3���﷢�	Qlz���\���f Ƚ=��1��9�:���&s1��hn.�waW�wn����G'U&��P8���fJ�U��3p�,H�)Z�[5wn���
j��Ȓ�)�ò6�β���$���{�����{����ϱ�{���n*Uqg�6�a���F�bR˖B��	d�6���\9���eN�z�w�"��JR@*BR�hN��sNk�n�8�9�M��
AB�Hı�����d����[ �P1Q����� ���ohK��1Ę���1�����6e �f��j6ܚ��Ug�<c�
���Ln$Њ�$��H��.a]���)�����~/>�ff
�=Z�{���R������o�{�N��f��L�]��vsa�����E��P�^����y�#���	%��ԭj�$��W�ٝ����f��><5��fc�����S!�uIr"�:e��C%M	���H��5VjkoF��^�cY�Fd�:��1�o��
�4ﺵQ6��v�<�5wlN.�hAʏR���X��W���
2V��;�ۃ�ۻ}z�׸lP�"�P��   ��,��#�%�1�~|��� [�'��Kt�n��r�9�a�.(,ֱ1��Z�����n�Л{eu���ДNj5�%'&���,�<6gc,`g�K�ˉ�&�a���H�lE�&`��cg�����U��#��2��|�7�W�I�>�{dƢ��3]��@fc��3�Vg��n�Ȉ�s��@f��k|c/f!&mFd�8kf1�u��a�������z㬶)�@����r(ԑD\h �л�\�5}�R�l�a�.��r��@'b	�u���3��{�u�}Ϭ(�Z[�7���@Q���1Foq���f1���ګ5�}��ɑ��.��:��\���+��HR"���b�\�r��Y&��C�	��U�Ww�*�A�{ސ�g�c������B��w�{�u<���d�1X�c[�c� �P�q���M�<�N$�z�0'UY( s1��W��"-GY�3�Wv��}@P���4�	ő���m�����{+3�9�W��w�o[c��Vb���)�`��7�WhY���kl��B��w�-a�D<����P|}�8hfcg� 0�B�p
���*�-Z��I�@��v��W��E��pN:x��λ!�H'�'�$������� +��q�л�\�GH�A��w��"-GZ�6kꪠ}�?{ν���oM6�> o[c���f ���"�&��s|uv���~d���w�~=���UUUUe���tی��k!:%g^(������kut�JM4�R7Y�j��D6��V�������ნ�	y�v�N��\	�W��V�hz�DgF�ǽ��D+Xc^��t��ɼeMC!2$S.2cQt~���z���`wWlGeD��c fc�sk��:�)�4,�5�.�����̑&�5wlo|h����M�ف8�SB���:��]۞��>�[��Y�5P����d��R�
���jƚ������>1��#��=q���[��c��c�۬���S#��p_m�iV���2QkC3s���n큫݈��*�V�]�v�w�q$ِ�L�2c)4ڛk����Jf5K���{:kl]��ٲ5|�fH��屃|��0�Y/	Ē�Xs1��k�J�B
/(P�(
$����-A��!�!�e�c@
�*X�}sm6��<@��c����H�Ef	q�N"nV�M��厛-.�����Û㫴,���/l��Zv�B���f���b���x@̌]ۭj�uHS�- A��wl|� t  ��!�]�d�8�����졫C�'N�!&A�����2�;u!�.�=r�+@�I)�swa�Ҥ����e�
I�*����5v����q4�Z{�55�31�����)�M�`�:�ٻ�g^�m��C�y*�VÙ�]���RO���9�w��z���s�U� r�J(��S)B
D�4��)5�"�"��n��]��I��,�����y��u^A����z   m�            U�D�q��Q���2m5fz2SƉ-#�a,�M �T\�Tqv�]j"���rd����Z6�A��%�2����,3�օ��4��N=�x&2�g	gmhC�T�P�$X�[Yyt�C���g �B����e��(B'4plTvZ�ͤ�;"�uuu\�ǲ�D�Ƭ�m,�g*2��
GV�t:����W��P'7�O����9�ڽ.�JG]�VE��cZՊE�=�M���NiR]s��m�q��x�ٴ�����tUQ�M���∶���i��ӷ)T�t2�.W��Mh�;��5�f�k���/1m��P�z�B�H��*s6�`��Bڪ�%�n�r�^���5
�2�MRݴv�-�RC�}_A�m[+�s���-]t�/#t��f���- ی��R�Z�*�(���"[��p�KkT�xs�����$�55�Q5\�:UX��B5ֱ	K�lMXԛ���*����=��O ;�@Ђu���/h�-�矃�����=$�o��A� 	�,@!����g1�QՎn�)b{l[��Ѐr7t�\�l���t�Z�𙩴4���j�.��v��g�[t�%�u��U�B6�2�,]ln��Ǔ�F���p���f1���I惍6QQ��g��^�w���O�2V��-HSj���ػ�Wk���!jH����5�1�  �Xid�1Jk���ڬ�1�k�Z���uv��<5��fc��f�˱�Z2Q,�SP�=nn�o��ͱ|�}��ֶ��|�� Ƚ�"�j3Wv� �PCt �v�����C�@=���P1��=�uޡ��`^�̐�R��ᡙ�fc�j�uHS Mm��uv�5gn$����Es6�,c-�M�(��MD�]���D]�daf�Eƒ�x�Cv�P�xZ�����1O�lP (?{��{��_�ہ�V��7�1�y�b���)�`v�x���!da������,�݂�6��A�cJ�ڰ.����Z3%s�a�l�ْR���@U�=�1�yֵ�t�"�� M틻uv����!��^��f1����y�wU
�����5�Ȣ2&ښ���P�_��ϋ>z�ψ;6���L�n5`�Wl��m�Wwϟ4�$Y��3f���@�I�x��ʠ)	Ά>��^��F�L!�ݱ7ǲ0T(�F0�n`{�����ƈ�zŐۡ}ݩ!��*���]��̕��@w��$�  +�u����4t�78����م�%6
���h��AqdW�;���p����9���u�'6R�L��:�I��]s���a���)�n]�Fi\����!k�������y�7��u���Ȏ��y�!�"n�2�����f:�}cW��#�'�c\㫾�dN�;����uΞ�dv�7�*8�,�]�c��^c3%f�w�L-'������W��O=���}81��c,��^�����Bqē�5v�7�W}b�凸La4.��(PCwo��ߘ�y�)Y��
틻u��T@�в�ػ�W}u���F� j�o��wlBg��؉D5�6�r9�Eՠ�zȸ�a�o{����;�,��؆�(؉�#3�Nc3f��2�i�2����Ք �@U�*��u��!�DS�5����ef[5��3Uwn�ޱdY^�����y3m���lR�-x+3��������5�~��� �ػ�5�o2ʀ�Z�4��31��X�
ٲ���5��5�:��
��{�������\�X�^��
� �i��}�I5�lp��ػ�*�\=�3�m��m�R[���Z���9 qĿ=j�'I��d�}��@�z���b-��Y�G�������t�ɍ�wn�ޱ`���<E�Fb`��s�f1�����c&@�в�ػ�W}};��*��D� h�nI$  �]֦���*K-s�<u�:�ҷ n�-����cs����+-R	V����"5ژ��R$��Kf��)+�Z,�n�5j��h�e�kvmuT��UԩU�v(���@�k[���vwFg���d��Hvۧ��¨	�4⑧��k|u��b�4�Z�q�����W��6@y�C��Hbq�Y��u ���o�;�ai=� -��c�s-���E�I�k1�o���9�{޲X�D����h�I|��õE �u�@uS���__S�]�o5;�I�d�ǜ��� �"]�F33��U[�d1� Q���NfJ̻�y�����1�q����n\d��wn��1dv�We�	ʤ42QZ�۸T2	HRj:�� +�.����;����{@Z�c3]��E��0v���Ɩ���Z���9�g{������:£B�|鵄��ڮk�Kq9|O��AĀ@!I��r&".��D�������'��P�H!A]:���-�4�D��e,�
YD�U��6�5�4i��vt���{b��a��E� �(��j�i�m��f�͵���
m,mOT�ҥ��Pu�\�dM���c
-p�B��}�Vf1� ��E��Bb`��fc ,�.�����Zl(Y��n��6�, ��j8`bJQha���31��lo;�⑦!�f1����]Y�%�x�.2�����]�u�K1��]�1��f:�ۮ�r�J�U����T_<�o���߬�V^��x�����W}cUU�|�F�!HB.:��n�.��$F�lשl�b5���7�W}uf�X��&2�л�]�S�4�ߪ���x �������6h��31�u�}b2d
-U�[�ͬ�cG7lo;�⑶a�f1�����s�^>:I�ΒI�}>�Q� �f�$�7`�hы��I/]��˵�B.���؛c����T,�07Yv�թY�2���'�����9�X#`퍶{RV�Ќ�c3�e��fW���.�qD���Ǟx݈�4�6�f��"�2BL��$n8��������{�XF˻cV���^����駙�31����I���<|i�{�u��!�D[$D@����w��1�0i���X�u��� +�!7w�2�r�aȐ�KW�l)�b�c���c��໷Z��2c���d}C�"�J&�|6f�fy�<�6s}c2F�]�5�:�b���qQ��3v�Ä�ĵ|CGWv�z@w��^�p���E�Q	���j@JfN6x��]�o�玷]����I��?~��3�B/���A0]�����r!���w�I�S4y���w�OjV� �*�x�ﻪ��A)\��#���33%ky��d�Zh-m��ce���c�F��e,��.n�+AJ�8فI�bY�k�uw�,�ܵj"�*=�u����h��5��$-%f[ +�.����e��OA=�![ݞy�P(� l��9�Y�.�"�)J�=�9�:��@r֭�̙�wSr*�(^�mՐ��q3B�߈��0�B�u��P�Ù܂�#��j�2`�E�d�����-��"2F�����w޺̶0��Y�!q��л�\�]Y�v����g�_�� � ��5Kd;`t]�tmu�X(�4��J��m���s���[r��.�s�r["���#H�p��s�ԝ���3�	�mbۚX��F�˶H˰��1krی�6Q���'t��:v�,<PvK� �T��2�F�A��l���]�>f^��	�����2�-���0���31��X� �Ȋ`������]��5����Lh��:�{�0��nV��b�1J��
�驘��u�g|/�$��6!:&�͹�V���gM��� QhYkl{3%f[�r(��D�k3��}��ڂD)R� �A ̙��j����@'����ӏC��v�W�,�&,�`�4�xFf:饘�f:���r2�zOu����f?�lo���7�LaA�,R�n�K�j	�$��$E0b5��9�:��uf����&���p��u��c�vpA+s���`��6(�m�{u,o�q� Qj���ػ�W}c[�E����7���;+2�a����fpz�ܰ1��5G'�=%rI
���P1�wn�޺�Hvؖ���FR����+�.�:��ݽF[H��K[c3v��"�Ȋ`���� �c�]fu��
(�oCo���Z���p�Nc��N7�!!E�,*�m�B�\܌b�1J̷\4�� fc<���@��x����=�:��;�v(���G3�{�Yv����F\e4.��;�Vi]�-]��ƛ^#3�R�S�{�u�H�~ʤ��j�h��?��/��?�m
W�}���V:��������Mww�5U�����u���`�6�oWwAml[u8k�'�'M�M��me�w>/��=be�l�m����M�6��͌�e	��`�X�E���͹ӛc����l6�����cql��lZm��0Vg-��Ŭed��\M�B�ޮ���

6��&� ����`������" 怲'�7U�?�z�_�����V
~��Ȫ\U3����Z���G슉��ϴ���3���TL_�~[��tY�>�=��"�^� ?r����'���G�����S���`~v�7�����_����ҳꔟ¼�(�������}}Oȇￅ--��Y5��`l��o������0�Ҕ����~ˀ�C�����T~���k��7Q>���1��M��u$�����c��f�EKUT�"3Y�-�3��'-�����`�����2�ڛl+m�I�چmM�ձ�)���V�%k+3V�ձ�3�6gb��Z�����l�1[m����f�6+ڱ�նbLm�f++fڶ՚X��Rj�i`��+fQ���m-�1�b�eb���fV�BM��V�aL)��+fSb��Ʀڌ�+Jm0�C&�lFB�ƙ:� �ALߦS�;����l/�����I�� �����ED��k��?g��g��?@0=���t�:O`��?y��j��?�� �耢 s�����83�������.�����}_�����?��O��I�O����C���  >�� }��������/�oz���?{��}ʈ����@�������~���U'ͣ8~���٢{���b�@>Hǲ�?��@
HB�_G0+]�*$�U�UUP�z6�õ�p>���:Ja�aѰ P(�_�ؾ��  ?g�>������"���_������������~c��O����>����+�JO���ـ ����?7�܀
 |�ED�h����������?�����~�}�k�Ѣ���D�\��b~ d���m����}[i����  ψz��|�oh>X}���'@QUC���ި���k������`�(��������!�ED�k��Ѐ(���>���Y�n���`}�?�6�B+������"�(H(ޥ�