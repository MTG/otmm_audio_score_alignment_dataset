BZh91AY&SY�5٘��_�px����0����a��      �su���J�j�6�*�  ;���@P *��Zv��V@ 4  M4[4#����   ��*
�����%T� U(  (	@BB �(P�)THQ� $PC�A�     S� ��4�(TU� ��Ը��Nl�g&{��=/� +�,��97l�7[��� ,M�r�&�  T���W{�OT{� ;�iM^��8��{��T�q4�������h�Y��XP3B�[ۀ=4p  
��J	�AAӛ������^-^��6W=��צ���{g�J�����ܜ}j�o�����n�[�O��_-swz�uﳽ� O��j��6�������_M���S����_}����ũy�}@=���w���^��w{V���v� w�|
 QT�(�pwp =�ꜵ�m{��#3Ӿ[��Z���v_5snl�mϮ��ۼ���ޓ�} ����s\Κ�  )��o�on�jW��>����q>����g�m}���ww��:��P{�nNug,��Żmn��OZ� {�   �( $+���󝯯Wo�ޏ�w=�үzۻ�k�}j\��n^M���m=���[��k;y�yew� :�q׮�ܫ��� ;Ԧ__y��m���[�|�������(�z�sk�8�Nnv�o���-��� B � �- �}m�=��}g��o/-�9w=�>�w��{�R�o/���n�g��R}ނ���ڶ��ݶ�f� ;�]:�x�N��z�=/)Vm�ʻ��֜�]��ys{�����vj����}|�z��<��m�               =!&eJ��  0 �E?�	��JT�@���d���z�T�m5@шhhѐ hh=��$i��      S�2I��%Q�z��ɑ�� M0�!R�MT� �C	�4z��h?����x�����_����}{����(*�����]*�����T_�PUp	�0EV��*�EWQ����gP�����?�������E<��U�����?�^@�� �젿�#���� ���D��A@;����P_� ?��P�P>��G���G�Q�Q��Q�D�C�D~��E>�S�D~�W�T�DG�@�>��G��PS�~�P>�G�@�Q�@� ~����C�S���D�_~���!�D#��p>J�A��H'�Oҟ�~�>��C�Q~�~�~�>�~��S�G�O�~��C�_�>��C��O�~�� ��'%y ~��"���	��?E��ҟJ}(����Ї�?@�	�/���/����E)~��~��S��C���Cr��܏����E��C�'��~��>���>���B�H��?H}���/ЏЧҔ'ҟB�J})�B@}B�>���B�E)�"k0]@��Ч�)�>�� � ��>��<��B���C�_�~����?@� } �=��)�I���"}�_�~��S�D�!���}���d��O�9#�G� �yrw)�H��O��O�<�B~��!�W��H���R��>��C�~�G��G�~�>��O��z�ܧ�?K��ҟ@}*u+�	��H��O�C�_�&�@����?B~���O���+�	�'�?B}�?B�@}"'�	�} �+������?J}
?BB�'��!��)Я�B?�����@�%��@���П�>����O���O�~�>��E(O�~��W�S��G�_���T�G�r_�� ��O�>��G��_��>�7np} r%>��S��>��C�O�C�O�>��S�O�~��~�)�/ҟJH�J��+����H} �JBH?H���*�J/� � �������������wt;�����;\Qۛ�F;qg @2�C)���qF�	���.R��O����e�I3.�5�M��R�@(i4�cC�D	�L�3I/��ݤ�ū�A�fi���k+I�i4�u�R�^ݷ]��=\���<v=�Wk��v�s2Ի���G�7C��^;�Ck�L�1R�)5�����޿.N1+��20�0�C!(J�̃=>=���3��k����Ոd$�Z\,�d��FF�F�0�y�rvf��26xѨ5�tF�,�$2��������KȂ��t}gݩ�~]r�'��Y�ؕ5J��C
���2�٫C��z���>L�G�1�t���bP�	X�N.BX8Fp�:@�K�Rv�����-�
*�F�c����[I殷8ٳLu�tO<�|޺6v�!"�C6ePP�������Ϣ���� ��R��Y�i5�l�`���C3Y�3Vh�Ծ9��7��j�F߽��������ӆ�7� E�(JLL��d$BP�<=5닖]��GP�l:F��H�	N�%k��{֝����h��LkBQ���F:��]k�.9<���%���׸�J���'K�u1Rk���Cdhٔ�˾&o�.E8z�K�@a�c�����yXƝ)Y3A�u	c�r4US!�CB`�nmU�[\Q$���&Vx����u<:�F�t[�6�tE:i�)�Bd�RwH��A�s��]�Rf�-\;H֌t�!(Jp'0N%���%,_!�Sĺ9}諌�>�vd����]�6�AX�s��7���p.��#[�r{u���e���7�F���7�TvĠ0��\�H�4i4IHff!��hc4������jp��}������f���5��8h7��n��&BP�%�d���Aj^ܳ�N�@e�d%�$��]tAl�Y��r���iJD�r�K��9I�ګs�uiS�˥hd�h��;�9wֆ�_zbhٸ2��f��'[�&�6��h�ti�֐̵&��8�Q��jLj1�K��C�0��6���u)Dw9A��(2p�u��2�O^��
��iM`�N��݁��X�����ª|����r��������贙8�{xxy�h%�/������huM��� �Bc��e��	i��x� -�v��j%�q�>('jP�BT�T���E���,��!(t�Q�6Xof�F���:�P�%df1�c�nSR�TT��5�'��b	F�rY@��֣Нs�:i�������d���3u���h�4%m5Ǿ`�c�d�4y��c�j�5�p�8������#o���/b �ùٽv�n1'	*����㖞��ǆ�%N�(���g,�sa�(�\$�(JfBR��u���&�ɍm$��TQ'�5'�:<rK;�p�:��3���	��4�����vym7	BP�=��I��	X1��O^�kg��ʠ�2�5A�%9�.b`Y8�kX��|�f	���s���02N�)2�����q�08=�j!=�!�aX��`�'3�1��֭�fo
���Ѩ��  �����j2��t�Q�V6��)���y�enq:r;�N1�k}�͆�(d%	C�޵���������jN1��}w�����[ϼ.��p�cߨo��m�{���Tڿ��ꐯ��E�q�T�4.�w�L'#R��t��c,46���t�Gsx�w<n={s����5V8i�O��?�[�0R�&���4j5�MNF�s���&�Rh���F󝼏@��6=c�`f����;|Ci��LQ	9ܲ��KR����A��]�o<��f`�ն�l�f�e�5&Nl�vB]��a���We��h�:3PdA���Ǯ%����I��zR9�}q��K��
� �)���#�	AӅ	����l�5�Z����pjseF���c����`��:����ޮ�tl�ezW,��1�td�BP�w�=�x���u�ysF-��=|w8��N6HfbPV.�FP�Y���&����;�� ��U�|�L�T�Tȩ%j'�w2�R_�i��:(w��%`I��%	ј�r��3!(01p{�c��C%��ؖh1�0Ӥ#5k���I��c��b
P���C��h3�����u�K<s�(q�3A��y	`�Ԙ��	�JMul!)121u�69	���fÃ��D�d��BP�f���f������%	Yt3��11gymk��l�H���u�0�0z�5.=kO5'�>��P�������!-����ˢ4��`v9tS9r��H2�\���ƈ��	�r2�2q�!(�a���Q��hӋ��2�j�4�'Sh�vA�r��I�В�G/����r��NC���Z�.�5f��Bu��=�ti|�u�wö�]��RA�j��z�z��{�H9/��9��l��<�클�`p��q7N��o����;�F\I3�� 8'�Ot�&I�Y�5�<�w��6�f8�ӕ\`}ٴD��8�Ġ������_�k�|�K�����ל��~���̜Op�{��kg �Fw�;ѼMh4�v�+��C��r.	�Ֆ'=MJH����G��a�{��:>}�n�
!�h|��RqD�&�6."p�Ӂ9:��7�Mk���JN��y7��R�ugU�ϋj��Gޕ}|�߾WO����e�:�>H�������$ۿ��X��BH|$����Þ�q�f�PaA��n\��Xkr��r	9>N+G!\����������M}�
,�Br�P�ﺽC��m�y��`py'��z�}�Nμ�q��]���:�$��0JI��p`�OS�1<�;��GBP�㙉M�`A%=��u�o6bFj�$3�����d�Z�L�cK�b`Y3��XK�a�F�����i��R��/�t�\��rב��
W���s�����j��H�B�!GHh�Vٳ5�l+ ��C�٭O�r{ӣ2p�2�����>4��S�mǔ�6�;<��1I�ᬵ�8i���,t:��@�.X����mE\����J��|M�"��t$�'.ڝVsYgY6f�*	�g��l���,Ċ�89	BP�%	JPg�G9�>F�0�f�t�]j���lkXi<7	JP�%	BP�%	BP��	BP�%	BP�;��!�`����(J��(JI��|�.�|;�23��r��(J��;��;uK�!���2��!<������2��P�%3�%�u	BRk���m�fai���l41�;�;# ��-�	L�M��3m��r��9	Fv���3���.��b��&Y��$�	`cFBQ�mZ �y'=߼>K�ݫ!���-|$[rG�Wͪ������ýxtx�ݚܙ�	N��L�3��#�C!��zl���&���O!-8��:�_!:��X�d�&&a��5c�������,!��2p��,��@�|�]���U(O�rW=Ú���&&X��!����,vk4���f	�A&N>��OY����lǼ4C�N��+�� �J�����4y�o����7�Df��#ABP�8�	BP�Bw�''�NBPuM�%9&��y���G1���	#�Ě�b��H*� �Z�X%2p&���H�ָ`e�f��Gg<����(J1�3a�2\A�8����'p����(JNz�1'�f�͖D��y��ޤ:��ѳ�xP�����;yӁ���ќ]�	N:���O`u.9��Ѯ��J15��:�k{�t�Ѵ����rM��A�Z���06j�����r8Id%�y����00�5�^�A�"�%��U��E;�v��ugv�.�G::yi��^A�.�	�Q�O�O34��C��'fGTF�`b��Q5��@e�X%!��]��o����ŎZ)��5i]��I�>S�4�S9\�\������}�R�G�*MZPQ�qw�HV�~�U�Je!�K7Ʌ�2��CQ�M����Qe�e����aѢ��CI�N&%�%"e�WmʯL*�.Hw�a8Ld����Z�i�[���� 3��WPcFPaM\��u��W�#����\J��PvA�i�!(Jl<7 �Nj6�+X�E�A��;�a�J�m�Q�%a���Î�N��A.�I�*���]�ZA�'�CA����t���s�l�Vj�:�%�fe��Lc��n0Ѹ�8>k4����&a�6�˨b�"��+Ds�#B^�/����\�ln�kV:N:�h7:5l1w��^E�q�0����+(���t9��f����BPd@a��4cjq�f�2Lz5�D�;u�늬�Feڦ����pi�I�c^h�uI��㐵���ʋ�;Y_-9k�],q4ITd�Ti�������o����X;�Ϭk��(t�]�*��:Ar���LCli���ε%��e)4�5j�Y1L�K����uH�(��wuaTBJ8	��|��|`�UVV�-��P�UJ�6۩�V�44���nI�������n�߇�?.�}���������8�d � p��� )R�� �@
\ Am�A�������� 8�� #�@
P`8 p�Ȱ� �ߧ��@
Pb@�J  dq��@   ��[pam �8 | �J����  �m�  ��@
P`8 p (0 g@��H�8�d �   m�  ��e0       ��  p            �         m�pd  t�    -��6�d �R��:�+�@
P`8�A����� (0 8���J��u�H-t����[��6�sj� [Z*B��9ό��C�!5U*�T��UAK�EYZ�z�vj�s�#�ٮ�:ڨ ���6�m �[a�m� 崶�]��v��ӡIUr�U�T���(   6�6� 	$$Y=l���8��Ҽ���KhhW��ٶl�UM�Q�PRRu�6������� R�V;s���+��pQCD����6���`���zГm��8$[� ke]���l�[J���6�� ��׳�H�X>�������|���{}�C�t����vŔ�w-�$���th�M��-�m�K	�w6gK� u���Pz�8�Sۢ��z;y��m[;���l�}V�V�g�����X��r�z��z��E9z���=*��stʘ��n���UuPg�Lū�̶�vF�Y3���R����l��gw�?k�����]X��{��?l�
�Zl�m�| �Z�ԥ2�4s�z
vy�J:{s�v��ڨ���k)eB;JN���+l��c����.�ڷ?J�p�k���N�nT�܄KIjSm��4���UU}_�aȒ�Hi  R� 	ֱ���V���6ض�@^���ZlH�kV�r�sm���&�`�M�n�H�۷nqRE���Lb�;6�@�P�[v�8 ���K.y��z;C����2�~v;?�L��~�֫ʶ��v�p�7K�H��j�UX.����^�X���T�UuM�`�	Vz5� -�d��T��й���g�&��zS@[��uش�k��a�����Wi瘲��b�E�-�$�^2Kө	:�ki�ٺ��
#�6�l�m��d����q-sj�hp���s��.�U ۝h$��kYa�+�[V1��r;K͵J�P�bkt�$k���
v9z�t�eC�;��	�Zq������ܜ����n9�j��|�l&}��vR���C��_ǯ��_��� ��65\�F���l[�m�d�H8$ݶ����#����j��U���Z��J���N��Vl���A���I �Z@�:Am 	�����#d0��/���-�U\�AKHN� p  �h%{h#U��ճ�v2��s�ց�c��ْ`$��L�- hV�j����vь��.�Wf<
��hg!�gm��G��6�nq�<�k��6�v
�����8ꊣ����_Ci��i�;$�n.���v��9K��v��f�nv��R8�n�F�vZ�eZ�[%��xt: ��� �M�BF�mZqh�VRWj�d&UQ�N�L��UU�� mh�����d/]n ����$6��$���  �u�s�*��e�6���k�  h��nͰ��� �`�����e��gu�` [@�N6ݤ$h����h�t��戝����л��۶h�ֺ��l �$n�gL� �J����[]R��=,�Cm$� �`[ӧ[/M����)��i�"�x^6�ڶ	��N�ѻj���$��$Kjޤ�Ei�m76�gUj�M�l�� �f�9'Hh�8;i����v�`D|��m��k7V���3itm�� ����  ۶[@��  �    �)m ��[     � H�`�v� 6�x� l  GӶ��Ӧ���� p �v�����d�v  �Me�l�.�ku�		$$�6� ��I� �"l h	ѻlz��nX�լ �E�Q��� �����tI�mzkXNۥ�*�G]v�p���J�� m�������kYgk��eRܭc��v�m�I���[�6���pօ����ImȗU�ܷ�N6�m�H   -�hv�ޡH C �m��5���h�< [   �ifV�T�5X˕��;,O3j����n{��<��x7���/^$ H+j�l �l�h�m m�     H  ��:@ �e� 6�m%�      f�    	ݜ`���[L��3F���lE6��ڴ��>l����l�8m�G $�m؝	-6۶��[\�m9
� �� [G   �       �� d ��ͩ��Uu%VԂV�3̮�9J��
�T�#�����.�.����	W����@J�s�C�f�q��6��ܛl[[m,���Bm.�isa��4��S���g�Kt��uƼ�$Et1u�6�6�<�:�T����	�&�����)R�� �����%�  
Sf���mm���smi�ϒ�8m� $n�m\�mk4p4]�ֳm� [@�j5���` :F��   �6� �[,s�����m�m���m���qV�s9�nr�M����d  �k[� ��#FmÜ�ְh��[�h���Y��H �`ݶ9 	lj� ���@P�ɂ���$��ڶl en��[\J�r�P�P �b@ͯe�������          �- I���o��9#�o��RP�A��U�U� �^�[E���޶��c���n�m  m�%� �6������` �U��UR�֡ek��� �� H  �@�ӗ�oP��j���;� �����X[s�6Ͳڐ�������lH�v-��W'N['K- ��f�  q��s�ͳ�  �6ےi-`m�kz�u$	 7Y�0k� [@m��� m��)Uu[\qŷN�©@HN�F��gd66�k�%n)wjͰH ��UUU.쪱���p���U]P�(]� �`�˧K��i�
Q�@V�� ��A�Ugukd�گ)j� �Z�=��#���=Z�{� :�*�X)��Z� :�È�_]T	�R��k�#`��U���UV��`�WZݶۉV�j���A����b�n�6۫nS  R������}V��7n���f�5�sNT�\�MT�&"�$�n��z���d���uN�UXdq&H۳Jؑ���ٍ~�M�:#_��  W.�$6�m�Kh���=�{�m�   $   ���`{m'��6�[A��h� 6�c��   (�Rޢ�U�T궩We�Uٱ.Kz�	���C�T�XV�j�*�
U @ ����@'Zv�J����]'l�f��h :�M�nZ��V�X8|�շUR��[T�/� Uiu�mmUUJ���4�\�����6Ԑ�Q#�ؓm�z�        R�� �gRmUV1*Ԫ�tn���<*�UJD�R�5@�*�쨈=�5uU�� zY8 -�==�ym��� ':^����  [DN���m6�H  U UU�+;*�[Y>��m!�� N�  lH�h͖��8l� r�       ��6�#i6��h���HZl-�  ��À� p   8���Vۏ	�gm�Y��<7A��pVk.��e��l�n�q6�   ��|    m�ŶB�$�  H ���;Y+   Z�t�pV�mH��m�v� -�5�p�b֛l D�m�  7m����i �-�  �dq��-�&8�mqm[% -�y��U�H7 ��Pm���� 
(ک@ؖvVmPH �C��`���_x   	��G^�kd`�_��{�j:� Ljl�2�PN�Z�  �PH6� +km [�Yg����  �l-�[Rŵ���$6�D�m�i4� [@ �n�I�F�۸��BC�m�-H    ���$6��6��l6ۀH�[@    � � 6���� -�i� (
��ql(@J�+6�	� �   p:E� ���[- A$�8��`  � ��{�o{������*������@ :����@_���UUUUUU@           UUUUUUUTQEQQIUUUUU������3������|�		D��PīC�B��A�DCDLBPL-������?����2�9�(�(����r�9�9G(���r�Q�9G(#���r�Q�9G(���r�Q�9G(���r���(�#���0�a2����08{Ç�Ga�=�xݷ��G�w �2�8�(ڵ�ֳV������� ?�~��E4�1P�'@��|�I�2��Jm�?� 
$a	t'OJ!������i�+�>� ����U��P���VY� خt �x��W���z�oI�=] 'H*
,�hC���'`p �nP;6��"�0��'�c �o��z���/A⯈��>�ǤN�zq�G�_'}���/i��o�Aߝ��- ���=X"���0�!�߾�t��A�{E�p����h=M���ߨ�@����Y��B_T��4 eN�C�N���J'B�gN�� �4��S��L�AqS�]$(t��(>=�<v�A+20�!
!<PC�(M v�JeL�OQ9�*�<]�"J�� �.�^�Ӎ� $�Jx(���(@�;Q����8�":Q�� _#]��!��Ig�A�%IP%��(<Q��{=W@�t�|�ti��vT�)��) ��)aҘ:�<A��~*b�p8�Ɋ/�@�T G�T��U��OVEb)Dd�� 0��(�b���df*�bJ�%ך�<T�HP�D���p6���DL�Bm�S�"$ `�@+�H+�(@����P�6�+�����PU������o��>Q���o��������˔\����������~n�7�����
1HD*d�z@(X$
TT�S�('�I$�o�wh��d��B�|��<r
��J)k�p��+�Ƌ�Z������'v�_��{������ߎ�qm���p�e,� 	 �=�{:>[@s��-��p �$ �p� m�L    ��g mS[n0R�0l"�b��mʶ�f����.Y]���&w�i��;���c�rXl[��p���y��8;]�zO~��}��5K۲��;+��G��o���}����-o*�d�My;;�(��5c\kͺY\�/����gC; ��o<۱�!7Q�d��.�T ����ѿ;~v��s�����%-�����>�Z� �a�� �O�֪[uM�̷Bm�(��Nܮ�L�?Oܸ87���X��mU(;���:�H���JٖɁغ�Jܛ����Vwk�۰�{�U�v�j5(���}����:B�jո�ͼ�f�f6kY^������h�,0i)�dȲ��n��Zs+ˈh��{HmY6�9��$��C��2�����G	4�T�UU*�'�J��p啸8If%�N*�j����l��\S�KP�9kR�Z̈́ɺ��bMF��H�X����6�"./-����� h���M���kU�"2�.+�n�JR�UUR�d/ ���Y�&�o9v�z��ЅԜj������@�s1�=��.T܆�\����)��ۯ]p�9϶T�:�#�:ȳ��;Vɝvs:�Wd
7b���VUc\�2�T����q$%,��*�7f�v�7"T��4��R!5	�;\FF���)�^Z�UU�����R���s��d2,p���!�Q���9�d�;^�n��ls����i�S�N(�A5*�j�@�SPm�z���Y���=����v4�H�ւDt&���m�����{�CG]Y�u�I��+4��u���m�V�n��� ���r����ܠu�xWE{u���p���N���|K�V��'Yu�ϠXc�M���m�:^�jI���V͵H@1�U]���t�^Ĝ�I	p�E��z;b�@$[9w]k��q�yZ���z��Vo3y�ٖ}��
�"v��<��D���
<8?8�?���B��T8+�b����~�?*�RS����E���Tk��@[J<���跐[���Qљ���X�-�t/&��]��5���d�?EV�m���UN�w̗������qk�]�����}���@�v�x�m!f��Qi�<�q1"�J����U�7m�9�f3��e�6��n9��x�b�7�c�f�=	�0��sm ������9�:�:��Wh�)j���v�k{��1]#�W�7+�c��q����<�˝�<�L+�nܘۓg�3�^9�pl��Jp�UACJnR��Ʌ���� G>������ɰ1yy0� [���SUf o�^?�����N��j���(ci�R�RK ���`l��`�������P�1wTԔ�U$�����]���j�>��,W��,{�cj�QTC��G`{����W������ q0Ĝ�L�{j嵓7�c��'���:w=;�ŗ&{[�"Mci�n��Ӡ�� r�x�R�aʹL`ޞ�H*�)AR��%Q��KԷy�pi��}O;:P�\|W��}k����� ���`ƫ�U�
�� ��*�9W)���}��� ����'q���8���~ʰ�+Ϲr��}�!GGD�� ����j����,�W+�����м��&+:�'���O����jQ�	!�)r�,;u8�X2��&H(�eT���Z^�d�r��<����do�D�~����*&.���������~�{�|����rNk銸`�D�KY��W=����s��p\����
�(�������~�����=�j�홐E�E�us�{ܳ���j�y����w+$E(�Q���9|ϳ'=���Y��W�}��֤���hja["m�M����d.8lP�lf�9ͦݶ5���ɷ-��W�i������L�R�I��m}�{+���g��{$����<R6�U2:m�_e{+W����˛��{�G���AE ]TŐUU\���Y�y+��^G�򟷎D*��f�[@R&�\s���/�w־��D#�$BC@���S�x'�B�fk�qw�U��H��t)$�W�{-}��{�{/��2s�߹���U��t�*����l�^t���RH]]���i̪p>Y��W�D:�:����6���촽�dԒ໾ݴ|�h��H���
&�G+���e��fN^}�k�e(}�����Ȥ�\��P�����^G�����H���q�� �T�o8�h�n���ms�}쵩$g�g;�1=m��dtۖ���W5%�O~\�����0���߾�}T�**�{��gmzK���m�������u�-�Bh���g�V� �9un�s�S�\�j�<�1��z�L���NTn�$�9��K��3�`]�u!��tmmչ�����Q��	n����⨊�D)J�[���6�\ڜ�e:����G]Z��V^�\s���wV1k���e���/;Tl^��M$���spp��zɋUt�NC-���w�{�����y{o��x��՚�vEnVe�h����G�D��mq].����Kr���aR�S�E6�s����̜���k�eP�w��c*����/��d��s���^�ͮ{�{-w�U�t�Pt:	�w�/r��S�o�g�r��yp��*��������!)�?w��>K���d!qS*f踙��.�~��,�.W�/r�J}���K8��jn��m�ET��b�Rs6�#y��1�C÷l������w ֑�Ȥ���n��^}쵙^��.>�m����q�A�$���Ͻ��<_]#���t�v����	�5������e�3�4�qgO[n��6�!�N~�{�d�+�w|���tH�
	���n��"#�Os�ӿ�y,���r�|#&UduH�Zfg�s���]�o*���p�َIHI)ʍ�|�q��	�uD��]p1��l\%3K�m��[ ����)�4H��';�̵�^���������^�1�N!F:��-fW�����O��ܻ��g�t�%T�E����x��~{����va	��Dz��>�.:���ϫ2���{!")7"�DGs�r�f����yN�t��FL�ܢT�W7EM]�]���9O)���Y�.W�{��?�x���]�pݵ�VX�v���۵�$Ilu'�5�uV�������k��@u�*��9O)���Y˕�X���P�HP3Y�U���rϹr��y,�S�Y�C�(�wS0\]��ɧb�Y����}�-w�TfURS�h�T�-H�ۻ�߳߰��]���u��ݮs�w.r�g�T��T�$���K"9r��W,�q<TQSJ*¨�����i�bl�G�3����q���h��9�7��r�UrUQ����2��{';��Z�W���{�	���I"
#��.W$n�Y�)���Y�w(�qtT�W��U���ȮU�~��+>����G|tR����,��j�#���%�r�p�z�Z�/*�%�r���fZ��q#w{�<���?J�GE3���.�U-���\�j�5۴�C٘��z�nuk�������wZF��۱�u�7��sn����S�\���^2�$K�@�gn����B9Z���q�݉%8a���1�m[U.w�Ut8����=k�N��^��ckJLg��D���v���9��-%�y����M8�t
ֶ���;>5&n�S�mb�<�F���b�K�N�{��ǻ���{��=����
�sj�s{{͓�յ��G�~�D��M]/F�4j�f}���'����Z���n�Y�����Y��I�jJt��Nw���eP��ٗ�fd�,��mB�B�uRrײ��ϻ�e���5�}����>2�*�(���������K>�%q��DyO)�ot�&����������������dyO)���Y
=ԭ��ؘ듡���۳mr�7gT��m���ȕ4�ݹ_K���9@���\]����oP�y[),��J~������6!sw�9D�z�uTȇNN��������9_s�_�J��S��_3����+�pY�ʝV9U T}a5Us�o�dGy+��dyO)����btP�)N���_=�d�}�<����R^���]�f:�RS�N:�r��fC�I� �'�w��!�B���N��e���zg�&��vy��7(8�ܻ=��ܔCO<���62A��v�/m��NB�������ܳ��W��u>��*����`.*.���{�?����7a�'��<��D�fV¢)7$r �N_3۱Qy����w_���_���{�ݶ�k� �mt���~��:ס�g���K�@�`d�]�a��$f�|ܜ8d�#�M�����h���?�r����U���3,��j��@��0؎�=�!���O3��)&�J&X�J�	BA���F$c�-�CY�X61c�`�A�8%P``M�N8e	P�hA99)WFf���+��Q'#,���X�.ÄU5Eh�)(
Y%�	Z�J����u]��k���qc1�\��,}P��ꀡ������Ud��{�HMAIM��GD�`�i��vJ�@�����
h6���b���}^E����"�ڀ�1@O_:P�S � }PڠH�a�x*�*@?��e���Q����9Ɓߝ��R�������(�����rJr_8�� Iw}�k�!Jy����?I�}�u�蔠W�ݗ� �.w�U'��UL�q�]o|��JSϽ���(�Q��w� �R�rg�{���)K������m�w��~��y�N9쬯�vX�`�\phn'rڄ����txj�7M�;s�o�����J� �@��r拈@�/w��Q�JR��~��iz�Ͼ�Da��w+K�A�WV\�^�r�b�T�ԥ{�o�~��;�����h?}���)=��~���'� u�j�F?a�mn��5��JR����~��)Jw���┥'�����)K�=�|�JO�~��kM���5������^}��p{�%(�~��s�ԥ){�o�P��?�a����&H�1)�L��UH15�B���}���~}ݫp�~�����������U��r���,�ۥ�v��$?(&�s��7��~��^��D�ϒ��dq6*B!J�(%8���mV��A��Z���ц�{v�Y[�����],f���{+7����){�o�P4�_y���)K���|R��`�����R��|>����f�j���7��JR���>��ԥ����)@������T�3ٲ������,O[n���k{�8=JR������&JRg�{��J)K�=�|R����>���)��cnAب���A
��e��R��~��)���=JP~�;�������^ZK�	�T��ETՏR�����#JQ�U�������R�O?}��F����=���)�a��+�
`	2�~��̟�[�?���
�U,�M��%�,8�;'M)��
��Y69�G��2�����x��[$w7mWi��M�7H��q�g��X���`�T��=l�f���� ��qt��7�}�{"p�8����;Il��^��� q ��Qq&�r��Z�l憍n��cf�uκ�qԼ>f��0ь˭6�F��kzs8�Y�d��7j8	{-֝I���v+=��w��w�w�������9��H�k�I4���w�]:K8���;^�7n>��W;Yێ�r�]9�'5Y�!F��˲������)I�����JR��~���Z�w[|B��$�[�k�9�N��\P�i=��~��)J^�����!G��eZ���,n!˹�T��f�E��g�(}��߸=G�$2R��o�Sҡ������JS��V��A�~��St�Nj���:sV��J(K�=�|R����=��ԥ)������&H�{����ԍ)�| �T�lc����� �$��͵ΜJ�
����┥'�{��R��#=�-.8����`ܪ{q2�@uM9��{N�/d��rM�5���f����i|\L�Z�uTȇ��wk�9�
w����4�'�����?F@�{���:Tz! �5@w�߿pz����ծA۩@9�P9��q"(��{����t�*�ʜ@ ����o�R������JS�����?��BdB[�夹�
�8�U5j8)@�{���JR���>���R�g�g�)/|�ߺ�ܙ)ߕ��0־���Y���|R�hN���=JR���~�)JR{ߞ����R�/u���8��Aū7u���(�JKH�.�:q)N�׿g�)}��~���)H�{�7�5��!�����)�9�W���<�論-��hƣe���i�Vٶx��u7k.L�3n(������˶���)JRwpw�)J_}����({��v;�)Jw߻׺��)=���>�t�SUT�:sV��B�g}�W�����c�JS�u��)JO<��=JR���_��5�V��y��R�_}�ǒ��}��{�R���=@���T�~Ax�g]~�ԥ<Fg햨�Ts�8�yb1Mm��dC����lz��;���qJR��<��R�����)JR}��I�rR��Q�c%�H����%��e��{�o�R����}��)׾oۊR����=��ֈ�n�{ݭ�6����5�rGM�9�K��Y-&]d��F7��*g�J�|ua��8��s�8��F���R������R���7��)JO;��Q�!�_t$�NBri�1�UZ��_}�ǐ)Ju��┥'{��Q�!B=�ʴ�"B��̙�&���F���9��R���w��(O<��=B�7�}���)C��}���q�Zm����UT��9���}��R�����9����}����'��3�(�� �	�؀���=��_\R���߾��f��5����Vo5�R������JR�z��<��;���qJR��<��R������k�����\����Nt�3��[��si�ݺ�'�9��;e�#*�+?������}�w�jխ��k{┥�~��R���7��)JO<���Az��/|���=��q�(�Si��㺐�k�9�Jy�������JO}���R�����o�R�_}�ǐ�J{ߥc<K@\�T\�i@D QߺfZ�)������C!����JR�g��A��]^%ȥ�:�e۫��)@�}�)JP�߹�ג��~��mqL�� �9'�{���JNJ<�(�S*u�T6�j�(�
���^JD	�~�ۀҔ�w��pz��/<���R��'H~�g�V�o{��β�� λf���5էh��.@��[��g�t!�uX�$J�n���F^8�:�2�.�m/<n`�:��Gd�i�N~���o^	2YBt��nrk%�%k�Nî�@�u�d�k���\\3���W��	��g�tr�Ob�c�%,:�f�Q\<�go�6D�-��Τ &bqv��V��L��t7#��5�cj%
�����7,�{���n�PO��.W� �+3Z�W]tMNd]��g_׻����}��n����ǩJS����pR�������)K�=�|O�*d�����@҇{�%:��́J�m��(]���=G�G%/}����K��ly&ᣜ]�&��T����͌n*�܊9e�o�ԥ){�o�R��������%:���pR��<��P4����ŭ�3F�m��[�����.�{�J,J!}ܬ.! P���M���+��o�Ҕ�ޞ鿳zֳ5l��s[�6=@ҝ�}�)JRy�}��R���߷�)J^���%)N�o���g�/ML��Ebz2�1i׫��GgT�FI�o���;U.2rȽ7�������	ַۢ��'�y���(�}�|R����ڼ��:�|���(}�y`�㥵(G"q�\�� �����_�M��ti01Q���_%G�<L�t,(>|�&iuߪ;���{�[JR�w�>ָ0�{��Q��BJ"tD��eN�j�J&j�!Bn�(�(���zmJy�y矾��JR�~����D ��31��ln�S#UV���"*)�y���'��}��JR��~��(���%)Os��=ћմ�)
#��q���tK��U�?}���JR���~�r��F}�/�A� �����{#t�|%7�����Iđ��#i�sm��G6m���9�٪����,�U$RE[�.�:qAr�/����Nf'p����y)J]w��)I�~}��JR�>����fhխ�����JR����c�����}���)I�����R���߷�
P8�b�b�M��"w��v�|r	*�����)JN���=H�
��� I��0%	p�ȡ�w)?����)C���v<��<�����s5�국�R���W�o��pz��/����JR����f��{߾�R��w��ٽ�o7��;7�o�ԥ)}���┤H���ly)J^��┥'�y����9ū^��	%9Q�pM	��;WPnvWe���:�-���]��id�1O����v��h�3xo0Ѽ���)J���c�JR��}��)<��︇R������s�9�Y���$L������]�\�)}��o�қ�O<��=JR��}���)C���ly!�9)��{g��ճZ�[7�zַ�)JR{�}��R������J C��߶<����q8���{4�RH�EQ)�/R�!3�}�|����>��R����w�hO��@4#��O_�� �9͏ҽ�l!0�����U˹9����(iI��~��(i�9rZ\�\�s��,�
@���u�)JRyߟ}��R���ߥ�9�]K��jj�NI�Ut�(�R\�z�7���7/nqb�8+I{n�և��F���ltȉ��.t�s��n�AMI�~}��rL���߷�R����~��R���K/r��\�a��k{┥'����^�UJB���߷�(J���~��R����w�����mk�l�o3vkz��JR��~��(z�߶<��� �Jw�����'����߸�z��;�#_dkF���n4o5��J_�B.AC���lyJ}���┥'����R���	B���W�D ��ٺ9R7H޵a���9��R��Ϸ�g�h���翿p{��/���|R��:�߶6s�9����뻻ln�v�$�*I$z֍�{��|�|�|)'�͹�Ɣ?lM��g�=A*:[a�`4ԆԐ�#��8tw٥6�(4�p���؝�����p�C ̅N��u��<P�-�d���1��e�tD���ͷFf�������|�%���}ё��sHD��	M&�4���׻g:��o�R"T�~����*�ET�T���?>�_o@p�-��6]n+n�#�?@�F�u|��Gl�-qm�0 +�s� )E� n�  � x<  [@ �,���8 �J���e�4<��B����$*��ԛ�N]I�:���XqOc�j��mq�	������l�X��rՎ�x#֥1���\[u��m���e���g�ɰ5���ü�vq1�n3�1llD�ϛv)繞cF�G=Y7M
�������b�Y�mX�B�Z��V�7V�#v� �l�i�T��m�VѵV��'6g=��W	��5�jH�̕e�7$i�iI�c�;���T������6��$GY��)���c��䑛j9(;q�R�4���Yt�R�)�Mvj���;0��� �4��T��l���7K�7L��l�xg��N�K�`���ӯ[e��` kM�6�@m��$� ++��b���%�n�vf^z�bU��s��l͎���^�Bpn�3�@9챫l���B\FH�GNv�d��}�y��I$��h��   9bJ.�/a䇂#�m���V�` ��=˥�m5�q�
@�cq�u�lgm����m��]�Yɀ2s$�gT�p1����+��n�$|��KѶ�$VK4m�%��3��*U��p�3MUT�p#��:�e5��3�@�LT�&Ir��ZT�ke�l�Diy�8`����٩RX�˸�]�"�V�Fg3'@;޽�y7gMNY�S�=r[mp��l��d��l��I@�ԑ�[�k9.�%� M+5����c<��w�eRy	�Z�]��\�]�.�3`�2�U-U�.�ylƓ��g!u�����-'[nS��	 �*���^�>؛�'&Nōשzv�`P uL֙bk���$�V��B��ѽ��t�������c<j�@k�m0Vʸ�`e�u�=v6m��F���Z4f��#UT��sOa������#8�5��]��^���J�i��^��5�C�Sb?�]�(��ᣊ�
��UN�G=DO����}~���?~]�U-��4jn�@:Ē7���ꛛ\���$�������\�
oWԡ{[�l�o�������?�����:z�=[�:B��bs��]e�P��+���+��-�V͂k���D^�Il��L�霍].��qpm\mR:1��.��	�!�ܭ�#��-ɩ�mr
��)�4d��0�&r]D�1,������][����m���8�dLt�8�&�O�0N�b'j�G�3��-�a�:�x� ݳ���z~,}(�j��ݙ���>����^����R���߷�)J^���{�Jg~�ۋG��h5T��J� �9ހo��lK���\�����G�Cp�T�!JeNFT��;���Ͻ0��K��%	���� 7ٵ`�yyU�fIrR$wĜw:8��&��=����}�,"�o��w�@��ZܵB�Y�w���"">���6d%�x/+E�>���ؤ���(qEH܍U>ܲ	;����]#�eFSV�6�j�\!�%����G�;]J�UȜr��3e�wse��d���{�n��/�B{Bm=�A��[�+����������S2(�"��"��w���.U�~�����6X���Cb������ws�o�ipx��t�� =�� 5"DM�qU@]�37f���@N�s$z��В��s�X#w<(j��)Ҥ�������O�?׀>v��;����翏����{v�bܛ��:�]�ŵ�X���t�ם��*�l��{_w���ػ�RTQ7����L�G�W�2/+F �o����ڰ>~X���]L��MM����d���5	� kn�?G�}�{1F���f�������޾�/��'���P:DL�q��� ��XX���K5�m8�55���B���m_�=ͫ�z�Xu?�������8�**PMJrX}���q�?s{�@Н�����3Q2UP��OT���Q���D(��d�t�q̤�����sU �9E6TD��I���@�l����7� �w�F�� 5"T��Tݓ3v`�ot�� ���3�_.����e)��
��z�� }���#�yZ0�ot�B����-!S%H�*jj�5("$���Հgrp�;��s��B���\R�Bd���?�� ���s�o���sG���Sltȉ��s�{^��..r_�g��?7�� "<�� oA����۫��X�u��(�N溝{G<�'Е]��!�|e)/�K�m]0���҂���� i;�m�DF˦р/r� �Ԫ�\��;����I�t������v��;��g8B��I�C�lj
)NK K��,A�d�����zks6t�f�!�hRu�z@>v����4��)��r���2�FD�	R�B�����@�ġ=�[\��{�V�ޯ�
R��#��T�&B&.�2*� �b��Oަ��l��kz�X�V֩�Tk�i�����&�����=@�ny1����T՞0#�'!������9{\m
���ힶ�"�f,��y�e�c�I�����3h�R0N�x���뤺|�
=����6أ�N�nT�,詾���:�ҝ��˽6�%v�]��$t-��3)^���z=2�N����ڵ�oJJ�0N H>.�I.s�s���&ä����O[�u��?fǆ\e�n�`"A=,R/\�m�g�1=�[<M�.�cM��� �Ӽ �����Z7d:�����Ш��2� ��͗�!Pg�3 \�~� �N��

P9�����Gi�s��M,ｻދ���� ��˜���b(0t�t�(!6�`���G7�� y�x�kN� �>�u� ��Te'��*�\��!ހ}�����IŞ�_����;��9��?y:�tJ��s{9��[�w�+���U�Nj�KT�wӓ����i�9ՏH�� �u� ��{h�w�8I�S�)�hD�uw:{&��./��K���
!|�_�?}��� ����`�2�b"!&�x�s��J�́U@�TX�n�y�xy��;�h�=�L����TS�HS\�kO��V��Ұ;�kņB�I	>�7y�Y�S��U$�w��wy�!M��!r�h����<�`g7�6]=�L��4*�!ARdGK13N��,����
�^�I��6��MΞ�t�2"Gc�:{&��f�z��i �e���Ja��)I҂�����fs��BQ0�H�VN�l-���������p�$<���M6�Ci�)��p}�ʰ߳*���KR"$!e%��$;�`��J":�BI�9ZX��s�/�cN�M�F�c�"��V�.�ݖ������fs�?$�(�k��V�7uӘ�!%���=�K�P$��y�} �sj�;�eM�Ծ��N���n�jP�f#�:̇B�l�9a�5`�Gb t�i3�͹���R�TQ6�T�6�� ��߯��x�n����呀4��k阻j��Ds����8�9�}�,��Հ}��-sb"a^թ�1�d�u��wx ����呀{��� m;�;Y�F)��2"Gd�:�M�`{�~�����߷�e�@"H!��),Q
=�G/;���՝o'�a�Z,j��.�0���@N�9�.�V�$�7�Щ~� ⡍���#�=�F��uі����[�����o-�1\�UR�����ڻl;�ʰ9��Ձ�w���vUA�CڒTg*'$�����d`���i�~�>�&O��~��dT�*�77\w6ՇY��9���`�l���FR�QF6�)���;ɽ�Ӽ ���"�.[-3�i�#P�
 �z��,=�n����`w��� ��w�m(�Q��rp'�V����Xzk�.���^����`Ϯc���6�۶�Y�/eӂ�::�k�'c��U`
ۮ۶]ْe`0cSɧ�(%�\0[r����Q��/m���<"vSbMS������J�S���t�*��]�b�z�m��u�㖁�i,A˴�lM�^�}8�k��~�}�}=hsv�%��Z�YqY�̹���ٓ��cg7����!����G[�}V�V���k5�v1c���dK�z�CY���m�Z��,�d�MªN�s�H�"�cN�$�'�{ے��}j��g?�����V�D�O[ltȉ�.�f�ڰfn��o���2���B���b0$�X�&((�������i�l��^˖F�S35��~���� M;�6�}�qX-{wy�7u�%̍몧ʊI%�%����=��V�����g��� "#aB�<٤�iL��J�󷃳H��Ʈ9r9�%`�t��$д���\h��� ��*�?K��}�Z�>i��Ӽ����V j�T����2�34��ٜ��P�G�ؔ4��#����T(x�
0���1�}6 ��V�"}��
qԡ�q�J�Ts� �͗�PQ��f(��L�/e�����uw0n�)F4�rJ�Xq$�v��j��sw����Fnl�;_/#�M��"��˭4�0#舉�M�N��ێ�^�T�Vr9#��qTp��v[p�Ҝ]Om�cGkSOB�vMÂ���E��s����D��`�E`{���ހf�`z���ĕ�T,�eڰ;�1	��[7���w{�	�xK�X.Y ��}���p�a���.I�UU2�Ҫ��+�k�=��Vb���^�n��mۄ����m���N��Z-8�BK�8G>��B1X5�Xފ!H���:aז�������!N�@&�f�\1�w��u�A:������3NaF�kQ������8��&�?�S=���3!�� ��(Ă�4�����4�b�|��D����<U^ 0D��=���� ����"|�.)"B���{:S?�y�.׈h{Q<�Pv�="���5�u����o�j�ݍ�J�P%vӷ�Kw6Ձͧ� �w�Gu5U��U0M���R�n+�Q[���Ip�͖ �}�;3�j�����7T�I%H�:Q��b`gE��l\�6�$쐥���眊m�����QV�r�SR��*������m`/�`	r�{�G� ���f'��$R�i��"��}����Z�=�s{��5K�8����-��c�R*��U\�g�Ձ��g8j�I�����V?ٮ��<b*�TYL )$V
Gw=��g�����~P�&�E�S�8�}��~�ʽ��=p��k�MU��w����8�9���eF��Y7)������_��˻�.x��㍰F��z��^�n��#t�`n�K-a�x���U���U�Kksj0�d`��� �w�97wLR�TIWn�n��͵��f��� �͖�}��K�2��������U\`�{��xK�X\�0��SjjUSr���p5(��%?�?א ���	r��;�Ot�L���u9%I,Po����n�qZ۹��g���,J?C�������w��
�[R͐�u��j�R�N�lڗm�X!�����X�r3e��`^�ɞ����#�klt99uk
&xŰp�ݗ����ƺF�ney0�v���]�6:�����=���Tb�HJ�1��1�q������*=�sR��1���Ӈ�����u$���A�� B�0�xG�8��浣L;6����K9a��7�ff�5f�[�{Ё�;P�.���Wy$r�=JYn�R�"	��0N�N�#�����mӰW=7U�/(N���y�wЮJ.
�������L��Otˤ� ���X���!(�N��
I�Q�p���I �w�L�SS���O#"  �[�m���EQȉ'z��,y�U�����̵`wws�{1�&eN:���R9,y�U���*��ww���HݬҬY��d��)���ݜ �6�hm��MN҅T҆�$���|�vz$
6���6|�V�v�Ժ��,�٠�Iغ�碲�}��~��� �7y wSSfJV��5R��j]Mʠnf�� �̫��.E�Ȅ�UJ�H)�b�W̯���g ]��*�U���z��{�"�cN�.���Z�*JpJ�<Ǻ@�vk��<F�m1�"'r롪��ڰ<�{�	*�=�]9�';LL�I&MT�}a7s�y��@n��Mց�9���a`���UD�UM2i C�K��5n�9�EYɜ���`*.��C.���5v)���7,l�EU_���`w����� �i��&�ꪢ����Duw�2OSS�T��m���U��W�v�T��i�S<�|vw]���}�]_�4��R��f����1TD��a��Ձ�/*�`{��:*(�MJ�nIV߷w� �7e��l��T��2��2�[UI�$�j�U�6���р%IN���yf��M��)!BlcU��t}d�rVӒ
t��G�h���p��{[���ݎ�ө�)��;�S1�U�>���󋐡	}��umՔ�ϫ��Z�T��K���Ss��D��� m��;�� �B��*L�����.n� �m�6��}����Α�%II�
"*�fT䱲)U�p�'��j�=���*�=��r��p�P�^�AR���{�3�U(�'���E#��s�`}��U�:����̃i�@o���~�e�n�yۂ�8�DO�\����wl��N�I���<���=W�/���X�}Wuy��[u�m�Ѐm��}F�,��K ��iUEi�RI�����������/�� BJ����P�骤�I5��ހ���`}�0�M�Vf;����%��4uJ1�Q@���.g�Z0>J�i�����D}3��V���f0j�̩%�H�2�� �s2x�sw�ݝ�`}���Q)1�b8��օҚ@�~���S�����-��n�a����a&X���$�ӣv[���i�z�����n:����G�P*�-�x��	�GtR���s;��4l�v4[�F7���mok�
\<QA�c��l�3�ݦ�9�m�N��g&%/%*��vLݵ���*ث������Yq�=a���[D��ntDজm�U+l���|]EɚM�q�n��uWg���سћ���ym�o��6ó���m͹�����[W]���Ii�j��O\��u0
M
M}a��;��t��<գ R�;<��m��UG"$���v���;�`[u�w���	������UWeO���\�jрIV��{�6�j�՛�*�%B��T���f�ڰ9��@N���DDO~x�$*y�&�˕JeJ�T9���Gw���	Fmn΁ߝ� �IN3��N�*����K�yݺ<��ɶ�U�K4��c\Om�z�xD
�JPlR�UIҒ:jSs�|�j����`w��=��.0���8o�ۣt��IR�QC�v~�x����M$�H�f�����y�=���?�Q�YM���غkݫW�7{���*����`{��,��ݶ�%7T�E���7�t����`T� ϖ`���j��D��5����G~x�:np��� �$W�L:"�ա*�Pȹ����v�]�.w���Z�W t�15�ڡ������_�}����A�7�t��n�j�ɉ/깫�4��<�{�t��y0��fRn�t�m5*B���no�u������_�?��HbI!b��d%O� ~�~���k��Xϟ�*�����*��I5����J!�mn������O���9���dE*m:�
�X#�-�}ʒ�9��4��=��A/~��q��<Z�ӷ,r[	ZS���YϴC��4���s�V�RU�Q��i�J!�vt2��� ��:nl�~v����L�2�����fs��$ś;����XǙEЌ��t�Ӥ��9$� �Nc�>�W�f���d�;ۿ�w�n�R�cڎA�	%9V	$��'��0T���{����ѿ}�B��/%���%��g+�`uo�
d�L�Q8�I�:kݫ \\�K�sv�kݫ�Ʌ�||{%ER��6�M
T�!v�s�ƣe��F	���7V-5����Gt�[*R�(�&�)
rJ�=��ށ��j��r`���X��*���h��I5@��.pd�;��J"wr��=짎�����@9�ʣYJ�N��)�V�z|]��~�y٭(I��ms�f��>gW��8�T̵H�2�����v�7y�=�����eab�����3TM}ad���7�t��A����3*�ؾI}�M˻���U6�w&��kZѭk^�rt�����::Rd��&�� IgWg��� �#!
��	.-6+�G������q�:H:_����bIa&T`�$a$e(���i(�&�!s�wk�tBF�8�%Q3D�SD4�k���������vF��Y�� I$0teH "b К	��(J�2���P���OL���Z�����sh�-7�F��tӨtx}tJv������A���fCe���P� )@@��� �-��I�rր �� R��
ڀ6Ѯ      ��,��� R�j'YG�(�C�ĭFq��D�d�ۮ�h�t�xځn�;�vdЈc0�	�I��3���Cc`�u�9���s�6�W\�P��1�!��o=�mit�5��h�GV|�v�g���:�y��^���wH�T�q� H�)cբ+T'o���ਘ,6�*nm�FZ��5m��g���x�-�h݈�T��ˎ0�#mljTsF�%�A����We�@":������l�iA3�n^���F�қ`2m�vQܵH�3�ܯ]�<��W^�S\����M��@{5�:�@��Km�ٶ,7h��hUT��GP��s���q-�7k-�WvE �� n٫v�h��I� �n�$i:9�gH�p/d��M���lL�S�\��ݳHB#h��-d�%-*��k��ӡ�$qI�:��Z�$ 	�0 ;�A5����a�2۳n�t�i� l�Y����˓Y�79�qIn�qƔ���9��
^P��M�r,u�[M����-���⹙VZ��w
i^��E)<� HO��õZ����[��x�bq�n5�lcU�����e��P�l�Ilӛt���U�:��JJ[۰�YѴJUnN���#F�֗�p
ppa1�5���p��j�ƕ���̑������Y��ѩ�-�k �و�McR�ڱ���&ҤnCc���ݶz���8�&���`nĶ���ɝ�*,hg1�P-]��iu� E�5�V����].r�q�9��6;v���� l��b4�\�� (����P�ڞve�%[�Z*8v��T�*K�msՊ�)�9�*�j���rIU��Y��*�j�l{��WS��a�ᑛ��\O���A�QaA��fh�#�0,�̬����|@�b?� @��	��ZO�(�e�����HE�<O�zC@�q�Ј�@��'a� ���1�
��J���-��T���mjg`r�ڤ����8PwGga��:�q�_J�Ód�i���<�M�c8�Xͫ+��C�O�ݐ�c�@��U��훷���@۳�1@�m���^���a����~�v��)f����Tqv|<W�N%0��mg�fʑ�\���Qu$��
a+;k�v��v��8�u��˭6�a`wg[Ӟz��9S���q//a��J�N�{���~�n>�4N��+�Vb���m3��C0۶� #��ۃ�;�%9Rk��
M��5Vr"I~��4v����0~���Ba���p���b�#�(�I)ʰ>ܘXǙ^�nn��f�ڴ� �f%!�qʗ�F��784��	�s�y�D`ؼc�TMS�*�!NIV �H����	�s�O��h�Gܩ)�!�nk����I5��ށ���X�XǙVnn��~^[�0�n�h��r�������f�3�]������Y^�("��O�\�W�.��DRm��)ʰ?f�0�`�ott���!��8���n�C�N��36i���=�p�	d	(T��PE�6�y�l��ĭ�)���ɪ&����� M��:np>�����iZ2�N�h�7���˖���E!MW8��ku�#s+>u�$�F~���̪Q���9E�M����%��}�D}��T��m���v��5}���T���'E�8�t5:��LȖtۡ%2ȃ��Y8L��m���8�rutA��ڰ�[��3���
��s�Z���K)RsJ�j�SUN���g9�C�k2w]�nw)Xçiq$���A��)#��*��� �Ә����Y�Fµ�	u��
%g�������s��GLm�53*\�Q5N���(�
w1]�s&���w{��[�`v�/'�m҈uN�������I%�����ݫs��3���U��9"!G)Tj�=p�׆�v�uI=���Y꺨�-���_�xd2��ܧ*�!�O ���p��;=����!X}����|6�2�ːx�E]��79�"""$?*Np9t� _���jl��j�S;5T�$��;}>�`y�ޛ2B��?�^�8��#����"����mf�3}�ށ��ﳅ������W=�5� ,u�pL��x�g�ֿ�g*��_�ƪ(��*� ���{w�q�Ձ����Ͼ����(��%L�;U$�ϡz�Lt�n�b6�Jع�m�M�!K^.��s�E6�䯗W	am�)#��US����_�p���U��|��}�B��*CNeL�E4���x�If?fM�o77y�7'u����8�T�%�S%f��`	��O�����7�0�ـcU[l���T����{�kV���рD}�%X�uN�0�
9��׻V�g���U����]Ti��_(H�����I�u�o�H�u�l�u�,�m��qLӬ���9�#O�)#�n�H��W��´;v�7,���˪�͕{hSKG,	�qf�1@c��Hs��ݝtQ۷b��6:W�һ�<�΁�rUv:�K�k��O6����uC� �1����c��u^юx���è s2�i���C�����q�<�q0�2��-�L��C�V��N����$�-�\J/���~9!$�Hꪆ7���i��U��p7*��s������F�y�{!ҝ*t�u�I%Xo����`{}���DD%�:�ֻcsuQ*��SUU�8Ǚ�z�����8 �S�����%	4�w<,�R��&�YWwu�?������}��T���� i �(��&�fk0��� MZ�����Ĵ���@//b��I��j���� \�B��`	��@n�j������U8�q��qҧ*,��n���8=d�ۮ�m`�zj�ɅP�_���7�~K������8��a �ot����f��Dk*���T���`g���FP��
R�����|�vga�?{��!�s���R��dR&������p?�Z0)*�9��@M�Ŏ�tۭbU$�*�p�ra`efc�>���z��j��nn���	��Iؽ�۬ ��i��78�Y��=5����U4�T�R��58�.�e�$gy��zݭC3���YM���i5њ�%YWwu�/������ �K>���2�1��i�5UӑӁUNw�fNc�[2zs-XfM�;���5'
"f,m�53*\�Q3N���� ���k��?����������^���>�?��:���MNTʖܔ�q5yG�9m�@�{�Ct���-Xf�uUchp���^�ճwOL��DCt�r�G�d`
|�`�q{L�٢Β2o��X�)�ʎS��4j[���]\!�s.���a֎z{�f�t����Y��g�}�@	���f�T&�m֪9Q�r��,�����3&����pd�;�DD&�����QCSUU\\�́��g8kݫ}�j�>��ʨ��"I�K�o�k�f�ڰ7ٖ�?��$��]�P�y"/�����M��n��&�S.���5���`~�q�ٔ�6��1�g���D�渚h��(�*T��ri�:o�7BE�g$ɶo7����������!2"�m:q(ܫ}�j��fc�3}�]�9�F�ڰ�x1=��Tڈ�E^F���X&��:np&_%����"p�� �%�d�&�SS`���思78�0��a�@�f��*A'�]��;y8�0��b��}9��� ���&ӧN�!�Ӛvw޵`j��#ә��&���Kg�_}���| @�\ ����w��w��e��OZ�&�c4lζ�H��9�^�4巙q-cf�j�ce�ގ8��rF�9���O6y������Vc���ק�]����t0�V�}	\.5�m���jq�s�ݱvl�6�5�v��{a�s�y��c3s��njT�Yh2�ny��6�9��;g��3��L��� ��p�Z�zFͺ��M!`eX:y��&(H�tB�Z?���������w��>O˱�.��g� �ջQ=8�������n�vL�ڍ���3-��e)8䟗BW�����3w7�@f�ڬ���eaZTQ��T89$vo�9͈�̪��77mX7���6g�m>*4�G���@�{�`o�-Y*�Y�����@3Uk")6ӧ����|�����4��	�78���bz�N��*�-t���������� |�F��ۂ�*ʲjh^Ʈ^c�j�����溺�ٱÉ*��i��O\�H�T�)��[tL�h�5<f��8t�����:RU�{�B�&���)�)U���cw�ON(F'����#a|��	k�_V�X{�����q~Q�f-��j����d:�sN��2��:RU����=2�<���us_\�
Rq�:����`f��z �{�a����?f�y`��E�C���lo�9�5$�{ku��̵`u����sߑ��GaDuhIJpOjӧ&ۮ�by��Y�=M��͐\�Ȝ�������J����]U��w]����X}���T��nn��X��&Թ��E�\����>�J��{�s���B�ؾg���vfdc��M�V� Ǜ�`�g�9��P�g�~����7s)Qʪ�*������v�Ƿ��ۼg�	oa��MChq��w�J�� �V���y@�`&�D����p�tYaj4�F$�L͓�5Ak%�p$���`@̔�[��"'	�Db�X��4z=i'I"#��	�p3#I�.��ad;{�Y���$�M8K�Q�F4��CN�����k'z4D�1$�	�	0� ��^�glf��BFl�!�Lf��h3M������:'�z���]F&fL3!I�vl��C!2�A�QCYr��̱j��	���	2[)�'1���`A�4�K�9��T�I�D6kXb�N�8`A�&�f�RG4P`��Am�A���M,��4f�0��T@��iG��w������)�?�����#DF�a�FFF	a�A;/�p�h�3y�Ve���-:i���B�*%ƉTp.աRQ�a���Fa�[�s6l�aa�0сF��hV�E��i8i�1��&1��4ƙ��e��S� �a ����?���ૣ�^�C���< ���<<҃�Ё��w�_w�pDG�W���{}j���@zImܺ��> ����M7�:np�d`�r�c�>�ōU:�5Tr!�ށ�{�η�TD&�/)p?fM���g8���w��e�׉��N�Y�9�g�[�%�n�[�ԛ�jt�I�+�,�9R�x�c�%��t�U�&���vA���X/<ɧ,N�j����\�~̛�ٛ�����vw���}}=4KT�f�$�*�� M7�:np�˥h�:}����i��Jd��N�����c�3��_}���a([��&�P%*h�A�_7�˯���@�-�hqU'LM���*�7�<,�L��V�����Ss�>��~_��c��}���n�����v��5�oo	o>y�(���NӀ�N���mE*�{$�I�h�C�=/���1��9�s�>V�ٓ܀�:��MS�T������I��Հ��I�GD�U�{�B���(w'�]�̦� *F
y*�M�@��Ti��M�*9NU��s��fo���M� �s{�}Λ��>n�iP�MSSSS\\�ٓ`l(K7ۿ|�w]���X�BK�BI	FB���1$���>�_�V��kv���a�j���6L�k�i�eѫ�t�gY {�+`��!^��z��I9���:�����i�+i��L�[tG#��u���۵��U���G�a6p|Y�Ӡ�K�H��N�u�lX�ۘ$z�U̩��tX���ۀ�'*�F����wiImmvب1�lnA����D��aR�FSYivaө/K�#Bi��A���0�/ȳ���t�eK�R�</�\-�k]�',5(�E��y�Mm"&{wTSW9˒�j���Q ��q��{����n�8�Y��R�� ��0�>UB4�L��I}��k���LV�'�zlgs9�N!Ba�X��&Թ��T杂7��V}>~�q∈I7�{����vή��93!$�H�r��p�)����@�M�Ẽ�Wy)c�[w3#� C�����p�(P��[����,�:��M��_{IByU���(eC+:n^��h��t#s���MKQ�����Y��P�ήx�����2s���g6߳'a.0�f�8��tLʒ\ꑉ�Ӛvw޵���a	B�	
'�\Ͽ~�(�g����j���ڔ�BR��rM��n��{�$�T�������ҝ*S2�TMMT��77��ۉ�8�0�W+���5�͗QE�)̺�p��Nc�ǩ(�ٜ\f;?f�W@��J9#t�E��%��4�13��7i�8y�[��ۃx��Ja��R�s��*��fZ�2��������v��^��l�DJ��#@N�:�$�H���o#$��g*��������M� �>g/�|�B���)�)��3߾�>��V��V'T���T�
���np�d`����}�ѕ������UA������RJr�.�ٝV�}��\w7y�3'1��G����MR���+t��>����ە
n�\S͹�6�U���7UR!�2��R����U_/�{��\����r�By,� ��T�Ua]�UWi���� ɽ�32��&��k&EJ����]W8 ���~��YIdVH&����Kc��:Lm�B�� �fE`ffZ�??~�������I�$,>��qS��G�	G�S���]M�O&d$����J����0�{�7M�N��V�.s�f����V�q�&�r���It�N��d��n�D�]7ۇ���n^ok�SK;I-��R��R�����q�9��%q�$�F�×31S!��w�)�T�����K# ��~����BQ*C�1��ަA29t�fZ�;��,��n�ȿSs���s_qe�U���h���	��@n��-n�X�wiUET"��t������Sv��?%��jK# ��_�}jb%	4�����3/�*�����nSs���Ac��*��[eB�v;+�����68�6]Y:��g��p9 	H�A�^،!���{r���&�S`���m��q�l�6^Ө���v�oV� ��s�ׂ smS�F�8�zNۙm�ۇ[��n�쐇;�7Z^�$��t�������qx�!�Ḅ�6�h9��]Xt�2fCFm��q6�-�a�L��\{���ww/o�����ϴ��:{}�x��ڌK�q�bd0�n5���x� N6̕M�U	ʨF�)��ԛ���j��K# I,�M�%
e���T�梉�v��y��+����V�s9�b��z�(l>��5N��I-R)�j� [����fs��P�L���=��`s�x	�[w2��)��a��$�s{@���~�rY� �Y����f�2}a7{�sv�
��l`�K# ������G���IHI)�:Bhl�61���8P`N��v�j�dJt�Ѷ[3bX��ۉ�U	:�ݵWA�fZ�3��{��l�����P�JrA8�\�̵�W�$�r!�(_B��}9_s�p�kKg}�V����74�ɠ���ݐOs@��H���g�o>�yj����`t�T��2�����s�~M�Ւ<�`L��?h
E
f)�UI�c�8Jp�7ٖ��?dvnn��{vi`w�fjj�N9��5/Yq%��Ѻv��8=d���]dZzn�P�"�����l�DJ��k�ef�3S{�sv��YHPT��TUU�EU� �otnِ�0�Jl��h���M��U���eaa}��9g�_8��*t8����~A\����<���IB���zl���pf6�E2��D�e�Y��g�n�I)��~M���,�IS�P �8�'WNVn������� |���8_L����z�GQ����e�$n�s�m��A��<rÒ�7e���m�m���	��B���d ��E�S��V �c�s�J�2S%7Rw�{vik�^e���V�{3���B�X��&Ե$�_��Y��FҒ�~M�	���;��+T��c�*�-t�����{3��̬-��J;�x����9��ޯ����TdUTi�"�vi��v�!�YJJ��T��ͦ�^��U�T]mͻ&+*9q�M�5t��5�:j���qmlv�q���`��*g�$Q�	�{�}��=jJ��uJ��`�Ȭ��b�%��@M�0�9l���*�5���en�nn��ݚX��V�f���r�C�r�v��f��7kE`g}���l����6����*Ti��)�q����٥��%��t���{�w����>��c_�������*���m6�m�7]�/��ė��k}��v���G$	��5�� �{W\lt���=����!�A�t�����z2B���hJ��O �C�j����C%5r: 8GOn��!�CE]�
F��)�(��Nv��@m�o�=6ڦ�^�6�"�xlph�/�kZ��ā=Ys�6c���0�D��\6`�5^*<RP�A�׀�� MCԯx� ��e���8�;��T�7}r�m�m��2q���k&���5�dp�t�l+�m�� �8R�pp[@v���`8��H�  �v ���� �    �A�I&˔ �uUPǶ-rU�iɄd��^0�
���bɃ@ج��ц�Sd&��6�<;l��(K�r�ە\�@1-�t��*<Ds����E��v݊���r�uҮ��p�N�K��Wm���=n9�O=^�6����Srn�bl��S�c�W�MNz��U\���0u�VȨL����<Oo�V�t\�D�ю�<Fوg�@��dv�qA��c�gq�Ө�!ni��WaŮvӤ�`,�H�q�kgeC �{n�g:ӱ�1p�>�9�6:{v\��F�r9U4�v�ŝ,���R����h�\�[�U�ۢ�B��غ��s�������G4�N��,��24Y:k3�Tu�m�l�l  6��k��%���l�t1[�n�z�%Z)"�TȻP�m7mH�q���G�<vK�Z{F��m�H�4��v&�f�W&��6t� $$q&�  ��q��M��v��}!=Ъ�����UjZ) ,Z�Wq��%��CM�x��8����t3��t���*�@�S��@uR���=s����l%�3i��Yizʛs3G2l����:Җڬ��� 6ٳ��Kn$=����)l��eke^�t-J�`�� |���"�:����i�qV�*�k��A=��*�Y7 ���U\� �N(���(l������v�$�l8��z���ڊ��^A�O=vG�	�V���ొ��8Ѷ��ΡN�Enw�ݬ\��vz��d��n��ҭUuW:����	�cl2HB�UQ�H9��[S�\=Sl X�>rn�In��d��:��u�5ݢ�-  m����8�lV0++t�ګ3��#i�6�t�����7 ��+�R(�%�^K\s��l�M��Ơ;M�j̭��[�=Ӽ�Ī����j{�kF��!�:gH�����"�1׈�p�E������"]@	�f� pPH�O�:A_Q^�ww�j3��sfĜ
�YV͐f�^$e��WTWeD�H\�����c,F����mv���6l�q��-��/2Jv�]���Nح�����6�����ne{!�"6��ۇ�ծT����Lڒ6�hu�'\���>A���3R�,k&�5q�v�����d�n��flqPj��(0�㰏h�I�쑺�����.��h�E �P��:q��yqq%W��^�ݺK	Α6ͤu5��]�M[�$U��qd��ۧ#�jw�P'��E���V��՟�sYJJ��{��nـ��g5�:Q�*�-t��vX�~�v��YD|	+��33uUdM]`@�oM�ݳ |�F���h��H���Q��'zn�0�g�@t��>��4��!��U:sJ[N������֬�����������8�+wu�0I:J���Wc;�Iр��k7 ��s�3e���uŰ�$�
RO���B���������vl���pfV�DGo�e� �3h"��P���3�n��qq#�=ET�zzPOU��o˕u��Ձ���is�w05�TlDtF��t�[0�das=)*��6�� /,6�
�6�*S���̵`zRU�i��>�ﾄݳ "﷣��Y.�Ij�t�Uk�y�d�#R��߾~��V��V :��U&�r:�rl��:u[���qΝ�t\���ٮ��q��:���\Wn�]��4ۂN;=��tݳ |�G菻�
]�[ ��j	N��Q�"�]7f��ݐ����Y[���n��Is��5A�RT��U	,�饙U���.q�.(q.G�P�M(�IDF|�g��p�Vt�����h�j�ygbN�́�w6y��+!D$�{ⴰ�솩Dۀ�qT�«��wvi`}��ӵTen�U� 75����#������g\��mv��-��X�R\�3v�س�۩.s�R�UJ����ے���4����X+����q�ۛ�����R�$�fj9��_tS��(P�g�fM�>���{'." sˡ���L�����癓`s�fr���o6��`��OŁ��UUUm�����L��̬,�����A�	$(��'9���{�H��j�r'Rn��y&�]l�:RU�o6�@����{q߷t,g��j�q�I;�m=:ݙ� ��:�h�9iZ����qn%�l��0.�`)*�7�{�F�Jo`{A{v����#}��en���DT���w�7ե�}��B@}�|�D�7P��;����i�K������c�7���ʩQ���'z��oK������6
�;��p#��؇��m�T�������y�<�n�8>�]��J#�� Z��w{���?Ռ���U-��%+��a&X�F�z�%�xk�.G�7fsu��*�=㎩��C��������b���gk&ɶ{`��I��W��~����L/��,3����س�g��&�5ڧ�V��&��䗈��zή�-�^�*Z���&���h�����p=��g��mל��M8۵�Z�b�pC�.�vւ�[]���l$�l�ES���o�cL+�w�QR=_}w(�֜X����g&i��:I�ɔݸc
=�+���)�/P}�P2�u%	���?>��9��� �eii }�zX�B�����6��7+�C�۽�9�f̴`L�rU�ϡ6{<���Ԓ┺�pn֖��da�O%X�ot�c.n��f��"l��0&|�����V����n�,��ӧ��#}����ݬy��@sv�˞F�">��ˈ�v�	���+lc�e��-J$�e�]�0Zkb<�<�n�7n��m��ٮ��/߿n���0(�`<�`}��U*6":#�'z�f��%��&`����گF�C+>:�V�{��ۻށ��tR!�n�s�)� .yO%X�o}�����ֱ2�FAS��Vn����@���<�%r��&ffl�� �j� �m�ݳ =��0��v}�4*�F�rU2�MGB�����jfw��t�8��CӺ{;�E���B�Tc�D�N��٥��ٶ���c�h>��{�3�{"���P�5*�y<��%[����ݳ �oi�RSc�A�NutA��u��w{Ӈ{P� �?J�n�)CC��4҈�z.��`y{XX��Հ��]�(�m�T8��H�BG~��ށ��L��3��0��`>�L�.��.�����6�2 ����7����7�w�=����F鶅Q�H�]�=��͡����k�ܱ�^{papr)��G�}���6�*T��}�j��fc�=��gz�������Z�
�)Tdr�@R6�=�m� �y��/��Dȗ�6z���6�h3S`}���=����͵`z�f>���QQ��V�F:�R������wx�[G��j��g��a�A��_1��-��u�s�u�^�OdRU8�R�I"�>�6Ձ��c�9�fs�w3-ZT$�z�nmU5U�c�۰��7%�^��ʜs#��l3ԇC��(�^�MG�*��ڧO�%"�-|�ݛ�fg8��SkaBK�G{�j�=��(�nD*C��`w�۽�ۻj����V�َ�}啴�Jb#��j�tm�`�a��V����Ń�EAD̺�N�Z�}�^�Ҫ��}����1��F@j��.$�f*bn�"�0��� �6�@�ݫ�i`|��^<�NU&�T�G!I.����嗵IAc�LqFrv�z���M�H�QcnM�SՋy;��̖�ɹ�nҗ�a��M�e�fȶG�s��f�U ��뒷l���p\��	�����*B��Ssc\�����mö7\r7k/%�V�Vd�j�\�c�O�T���u�ꗇ��Hu�Q6�%��݀��<�هJl����{,�,��ubWҒ>�t���I��|�:#�k��I�\ټ�ɷk���[]c/n��N^ok�S�Q �aE7
�~7���ށ�ݵ`}��V_}��]MR���M�qSw�6�0 }�# �� ^ml��NB�P�(���Ձ�ٟzl�
!D8O;�����V�3t�A�!)�տUUml�`g�w{��vՁ���,*��!D�n��9WsX�ot��y�yO%X�MLt�8���U1B�(��R�.��y�z��� ��5���x� Cv� �G:HwF�.���t�w��y*R� ^{����J��u8TrX�m���[�_�4��@iH�FRC�S�mz��}�o?
^�sy��uz�!����%K�Z�N����\�ڰ=�fs��w=�g[יj��g%Q�q6��n������_~��t��x)��da or�zR1ln�UW"u'z�f�}�X}�r�Ϸw�@~�����AHI)9
Fr���[^wi����g`Jq0І\-�����p�IT�(U�K�g�V��x��{�Hw�y�8n&��,��˚.�4ܝ���n�{��}�g ���4ۀ�q��`/6�@=��֊���s��32ff&r�*��L����˟��qj�Z��M~k�ʨB`Z!�����a�<E�Ԉ��&�E���IJT�Vd��NbtI�d���&���t,�fHA$! D�#� ET�0������T�@fk4�tnt���2� �]�Z�)�2�4��@PRTAxDY!fTFI�Q�L�9V5eI9D��a <��^4�RSALM4[�Q�h41UT���C$IT�$�L�Ԛ�p�Ȏ$����4LG�t�����"��	"`��$$����"1��'#�RÈ��+�/�� �~���X��8�p;أ۴N� {R7>'򈊙��{�}i(�_+-X���ϵem2:��P莜���͖��|����8�_n�z��Z7U81�7�sW{���`�+��{�ܜ�;��ST�q�%&�)I�
P�7��ыj�v<��m��7<�xn�AE	������h��M�e�]dh����<����}���V�b���*�A�3@MMU������a�fՁ�ܵ`�ޫZ�ެY)�-��n)9��p��U��g�_]�˖{s{�>� ��IT�(U�Uh5=���}�ʰ=��s��j!����t�
������W_����̴�T�SNf����Z�6��f����N��YJ�*	�����OB٫]GѻU��n����<n�/9�xᲄ� �pA�QIq
��:����uz��5ow8���Z�=�k9*[���YR櫜}�V��{�j����V{�oz~I$�̦e=_��N��94X��V����2I����y{+�hw��Tʌ����>��F �&n�ܭ��0 J*byA7T3UaW7q�&���&��l���9W]��Qf��_p�L����K'�e��� ,s���d�Xڪ������9L:�,Y9)����%�S=OE��Q��8�2e�黀�˶�.�u��^ܡ���]�=�������V����<�q�e;��۩��QN�iT+���'�&�G
�@c)i���Kkuu=���csۇ�{.�u�t)daX�ks]�5wg{��eǜ��wN�9��Wjp�QXZ���V;w�w��}�ׯ��ʃ��]=��ޢ�ݹݞ�&-tT���]�\����]d2�CV�Y�r����૷��l����7�d`	�����'�U9
I����3��;���4���� �m�SPQ��WeQ��ڰ3ww�;U�ɥ�߳-X�ـD�r
�:qX�'� Ӷ`�d`�d`�9�V7U#ӓ�=�K~ܵ`w=������{�Y68�|
���*���)��u�9�;H��Ѵ!�ՏW��Z���/g(���n�"�r�`w=���Ձ�糟���,1���Mk��Ԩ�A��� �sm_�А�! \$E%SAJTQS�A�XX�����r�`�<����'�A7T�M�w���r�`��0~�X��]MR���M�)u\�jP��e�`}��Ձ�w֬w}��t���*S��*�&�h�՞��ffF�'��l�h��)�M�TL�p���8bzp����1����<��Ę	"�RD:��Qu'W@�wmXԞ�	+g��%�,�ÅN�����@�iXnfs��DD6fei`}�m�s���ȈI6nyk�#�T�I,���� ������r՛�,�����Um���w�z�a��n'H��8����}<���&�0 ��OtJـ��Zڨ��ԧP�R�@�7mX�Ot��E� ]�# ���Tʹ9E��Ŷ�+5�Kv����!�Z�J-�,ٷLs�M=���f���Kn*�ͷ������v�w<��K# J:&���M�)u\��X^�%��mŁ��j��3�؅��ЧeU:sJ[N�����.e!,�ӕ����߿_���{0$���:*����!���+@}�������""T.��IDS��$�0JJ@!�������z��S�瞑JT�P��&\Ұ9��� �������V�2Ձ�i����UT�G��H��	�ZٝI�e"��G��֞v���g�Ŭ�Np��J#ӓ�7f��3z� �ݵ`w7w�uA��":t�MY�/sϲ I,�[otݳ ;��+Z"*�R�A��������s��I�ݭ,���`�m?/6�+�ʚ.�0���Sx��ݳ�(y��Vb�h�-���R&�����������;��V739�l�65(Q����������ܙG�'�Ur�,�fu��@,�������`�����T��#��V쀎2u�]�W+�+����R8��\��W��1�g��ceۙcmY��M���\��AY�.��N!��:�T��d���t��tiZ�l�R�l�]�ie�7�m�[N��m��]I�5�y7kj�6yɤ]�Yǰ�tv�%,�m�c&�xWf�3�c�$E���Z��ϯw����n;�t��H屚��qͣg�[�R��7$���]1&ddeE%Jq:�RF��Fo��>�zՁ�ٙ��DG�=���t�˪��:*�g �-^�$���� ���Ձ�zigj���x�M�
q
������:nr ��f rJ� �1V�R����ۓ�f�ڴ}�X��j�_��{� F�R��-.\��U�����,�56�@�Mՠ3}�L+{w���i�S�"H:��2]I�m]v��f8����SnJ���)����������(��@M�� �ۭ�<������3ʩcUP�Q�`w{������ �.D��p{��$�/b3�F)m��F┺�pͭ,�l� <���56�4c�)�]�Ӊ��#p�1{�K}��Y�����rv��!6]�3d�E�{��ɼ�[otNـ{����O�=)�� 6".܃���6�1�^+̵(�k�.�s�,��<�<�E���ﯜu�-�����	������9;f�SS���q ߼�J*T��1�rut��@;�]8��F ��{�DG�қ.n&`������`{ޛ*�{2՘��s�{��ry>ɽ�n���`��r�u�3u56D�d�̑ɼ�ϛ���`~�%��(}��; �M��bID��4���3�W�oe�w���w��`}����B���2�'#q5ܒ6�7�lγ�.rs��
����g�9�zlq�gd&��૽�9;f�SS�,��nk�@�6	�RTn&�T��X|ڜ#��ܖF@|����?}�L��7^��PڧMUW.� �nڰ>��s�{6i`}�ܫ;T/'��M�
q	�\`}�D|y�{�rv�ަ���}�#�$t�*��O�߹�G*�ߏ�م�܄�l#�'z�f�~Cݫ�fZ��{�{ހ�b�C�ۤA�|�$�u�]"+�Ƴ�#�m혬�v��\�m��v��)U"�r�A
p��X{2Ձ�nozq%�b٥�.��7�*"�����*g,�97�d��?x
ic4��K �G���lBl��)�`gͽ���aS�����g�Cܳ#�J�uZTN�D9;��U�4�7ޘX�fZ�3}�ހ�M�֚r��*���u� �%��'����0�����u@�G�UU_��ۊ)*��/�3vI[�b���B������O�߀���8f�Ć1��{��V9�uK�7��!)A�` d���$'��5�P�!�\3c!ٱ����M��g�[@ �p\Q�.(x�lxX t�HK,) I!�ú�<�x!���H{��=�[]�S�<#����
� �|��NFT��*T�Y�XF�B%OM��2P]�]�
~��]C��,�6���郪�����zu`�P��l��6�:� )@����@%�:�-��p)@H�� (6�R���     �$ �I� � UU�3��ӰB�s# �d ��v�1�$��h�恝l���h�ۊ���d�-<d�(���Ɗ�T��==��5j�v���2]��w3���	ݛ��'��7N���y;9�N���L��L��x`l�.��fXM���n� qw`'\<�qQ�۞(�㤸��ӫ0�7�9�5��Xz��m�Sd6�p+��p`�ܦW#ck�pY��O��p��&�? -R��Va 2*��3�'m�^��ۇ��b���A�톺3Wjb�َ�@[p�����un���ۮ��y#!�V����͵Ҍ&G�9:�δ��i���_b�l]Hl��ś���Yzۭ��� ���� ���3��x��ꦌ�����N�3U{Z9	����"a�Ŷ�(�5vG���*�.{veM3�j��)s%�&:�m�' � qm��^�ܜ�\�l&4�4��֫k�` �Hݐ�Se��H���J��l�M��
I� ��E�#�tqSlhG#T�kaup�m�s����e76�]�G)���|7ۗ}0� �m4�E�/m��\��q�eb���ٔ��K[*�b*���(S������I�.�MBC[I�5ž�T��<����qpg�s'<L�
=�����s ��4�����bw=���#qh����m���!j�[�uA5*�յJ���kv6�y`*�T��%S݇pڔyM=� ���}�\���V�����6�ab쓚B�FEH�x��j�X��d��Z��+m�A&�Hm��q��V]�t6�s7AU 	�I�r�Y����kvK�m��&�����e��E�خ���تK��f1m6ԵO�P
������0&r:tպ�·-P	Ʊm뫏7�Z��/b��f��Z�����Cj�� :t�آ�@"������g��D�J= '��v8��P�z��ݿ,���}s�CjYn�;g-�2LR��Ѹ]��&n��<���Պ�]ד���=}v��;��zղ?n�X�C����}�Ux�;�n^���շX�����t[�oRMn�eb;q���s�e��%`��*�7������\@O7 �s���E�Lml��V�90���!a�e�;�ga�]�$-�7q:�ji���U��v����Q&?��DF�Ƭ�ƚ^l��_Ϸ7�U��K�vy��D���IԜ:W�c�H��OD���a��#����v�0�9���nfڰ=��� �l���za`�=�
&��M�M=�9;f �u� �rY|-�,҈ې���rIށ�٥��w����D){2Ձ�no9m�~�)�mWW5pMY�?u�rYM=�8��٥�ߖekj���ԩI�p����9=�9;f�� �\���W�æ��v�,Bk}nq��z�î��$�p�lX�����{v��]ۗY*j��k��n���0 o��U9|�PV!�mTM��T��͚^�s��,���4|o�o�*��6Ձ��7���$<����V�r��U%�`�+f {������� ��䌚&B�5�8	C��������@Hv�Kk0��9T
&����X��ށ�٥��酀}��`{���:z�M��*�(�˗g��H�pX������p�5�H���(�h�F܄�l#�N�f�,�V�X�̖��{��|Wۤ���$r�A4+=��z�"!6#�̫7sy���eaz�a
>��7�����5#�8*�����~�ߺ�� �J�J�*�ȨN 2�o@#�߿u��U�~�X�@b��r�T�K#7q�ӛf���`�+�zO�
(�U_�]���� ��汚��3����/nM�	�II���U=`�Νu�,��.K���dS�iq0ІP[3��;XӕNDP�H�,�	���y)���6���;f3��EE�!T*s\��y�oRl���pA���������y�Ri��QE$���i�3ޓ�(�F�J��mTm�NF�7$�C�f�W��?nM,���	�B��*糼<�d�u4�h�n ��e�����\\�|�������=�4�:�����>9$��J��ҍH�6x�Wh1�f�ۑ����7U�'9@��%'*���**�#��p�mc{���=�!'l���� J +����uR��M�g�39�Q�#�֖�e���zmDD���0����T��� ����{޸�R����2l���Zlӕ*��*�&�`nfXXRJ����
��3����%E�e�\��V��۬���}-��NّW���i����~O~�sA����i��+e����[b��zz�n`�+m�D�.�v�N��L�w3��Zcy�;6��뛞Ų�أ[W pYͦ,��X�nx���11�;)�xgt�-�/!�+�Y���8p�*��sj�j%�E�2���3������ݚC���}�o��B8K;G��ϟX�;�R`�l<c.������s�^�}Yua�zY�Ѻ3mO`�C�չ�S;ǿ]׎���r�z�l�=t�ץ;M�6�v}Dg�D��^x8l�d������蛋���`?5��'l�	+�=)c�7ڱ=m��D�l��;�,٥�}���g�����`�ot>Bl���G)��k3��fc��J�7wy�36��ϗ|<��ܕRՎ���m����P���w;��,��`�H�Ԏ����z}U��s$�� �\��<��L�*��כ�C'�[˟n��]X�s,���\��F�t]�˹���("a*�4�$��3f�����JJ�m��9�,�VE��U��7wUf���x���Ȓ�-V����fl�����cP�I�N�w:��N�6��	C�d ws� ���M7��"9Vww{��٥�{��`v��;s�(�Q��'#dmK��ܭ��""y���N�6�efV�O�T�"S���H�RтC]�mk�c���NGц��M6��G�=讷�G�%P�`��]U�������$�G��+K K�`�PSrUKV9��>�&�����p�ei`�r�b�l7P�F���#����������k9p�����*Hb��B!o�DB�J��\���mX�=�`y|��m�N�QC��d��;��w�a�"!>�~�����&����T��Z:�>����}�v������K����c���ETq���G���srN)�O93v�a����`��gS����U����e���� ���@�+g����� ��6�Q7���v��{��l(�lﲴ�A��U���}6�~4[�UJ��`�R�'z�ɥ�u5xx�=5ʰsOtO&\��UU�L�
4Z�Q�f�X>�M��w�� ŤF
b��B|�m|X [պ�J	B�d��Ӓ.��y�v����{&��ܖ䏗��:M�0�n⭸n��ѝ�l�:t�Z�e(;5�6�0�%���B�T�T�;�mf�t����+�6}ʰ��AE��������ܭ��C���>�X������*��E��XsrX�r�����ܭ� y�rsSL�7���e��N�sOtr�`~�����9�Y�
&��UE	N;���~��@��4���ۖk�c�<��I$�%OϢP~ښ7��sJJh �ǿ?q��ߥ{��n���1[�kĀm�s��E�VB��\Yn:��7K�pv�tn�3\�u�5u�����g�& ԁ˜p]I��ô���,�3�[���g�X��j��sm�xyb�ӝ��;\r^�{j�v:1dx
�2�̀=�]mm�N��FWv���.��(8h6ԅu$��mȼ@�����֍0�[h��K&����t
+S��9ϒ[Đ쿾n&ꪣj>4��ҳ��3����3/��l��sgj�����1n�D��D0Q�Dp�@����,��V���J#�;��p�f��6�����&��#ɻ�=<�a�>�x�@_{&� ��K1V�ES$�$��O'XSɷ��[0SW�	A�����܎��ۛ��>�M,����	B}�?d�#W�R\�("f�u̜����gܫ sOwm������w��#;��z	�E!�6����̝;r����a��s���[��v.��wUf���'}Հy��}֌���t�*�S����@����.s�
��N��U�{�]Y�y���Wy���s�꽈Qٍ{S��*S4���.j� ���� =�ـ��6}����DuQjQ$�D{&��g���������߸_�Jt�C����&��M^t���c� �����d����"a["m�O�FӪd�a�$ٜ��n�qGps8ۖ���ܴ����|��ES$�$�W�]�3ۛހ}�����~�buձ�:N�#���'��� ����6}ʰ�ТBT �~�����:zS� ~j��?�~�u@ Yr�*����wn�4T�fNaVYU��#IY�c�1-��&	Ȳ5�h̲�Q�Gë�����E�o3h�9ǫi#�h�+������It����f'I5���z���H0���q�p8yУ�!+H����|S��'-i޽{��h����j���� �e&v$0�8�zP2#������ 8��GL�5B��8K�rN �	�"�����)�1/P�iP� gM�z�}t
�@�ITx���@|]�iUt��jA}.�%hw
%�o2��wٜ�7��c��:��T�X~����U���lwLÜJ!�j���떥Q3E��W��zy:�fW<{��� 7�,�.��U*��$�hNGFG�e��Nt�euQ�k�&�(Zs*���pDhQD�%TP�����ހ}�ج>�V�	DG̛wE�2��D��J$����,~[�����@�7�8�f���EH�qJrZ ߵ^�� \���� #T�%��Z���
ܒt�{u��i����������qX\�W@��Z }@�"��y����:���7��c��6��7ۛހ��#�͖ ���`v��v{գlhU��H��s�u&��^��[S�kX�v)��"͞�l���Y��q��;m)�n
���o$�&_��}I]~���?۠G1ض��46�R�U_q�ٓ�V(P�[�Mr�sOt�;��DL����L�Q{�y7�t����=�$�TWے���4(�r�(J��>��(S���p��V�g��mDB\}��ߴ[�JTC�I;��f� ~j��O*��\����G������BJb4[�N�E��[������N[��ް��I#p�JGZ'T:$'�ۨxVv�H�.���4��"��z_�Aq�m�[�!z��Më��xj�,#�[�b��[.�6J4�!���-c6	��<�t�U��{,uq��72��x��n"X#\��ؠ̮a]g�R���e���y6�<�D�k�+��d��v�܉9�1P@�au��Q*����U�7C	�*�%���s�Mw�4�S�n�
nE�sQn]�:Mj���\A�َ�[mɌ���٣�p�R�r��$���%��������y'x�z��Ȓf���˻��ғ������=�$� ے��������7Pq�ܗ]n/ߙ��� ?5x�r��ТAE :���&n�@<���� ���V����������PD������LǕ,� ]��G�'x���!�$��F�"�)�#�㍹6�V:�CY{-=(j�m�3K�m��K;uI�QUe�W�w��A���=�$� 7۲���4(�r���>�?g�u��*eC� $ ��q�}�����y��ɐ��x�!����jP��@>��`��`}�r��{7���i*"�Q�GQRK ��� o%x�Ot&g�w��5�k|��1�$�$�ٻ,��Jry��;����?G��Ob�bo4���l��K<�m]p7��걚�h�K�p���)�����^���e�KR������t�w�������10Zڮ@U$�@=���7۲�;��`g����.%�b�Aki�E(T6�K��,�̖w�ȗ�%J����T14
�DC?v}�����} o��`{C��Rp�p�s�%΅U|��w'��;����7x	t��QE:pe9,��{�3l����d�;�bc���m	�iG\�/']��W�f�{Z��ǁ���p<r�!�f�wQDuQjP���U<�`��`��̒�3���@�f�ET�H�qwx ���� ]��rN���u��H��:d��$� �7e���oz]Q�͖���^���c�H�j��ܞ�$� 7xDWD��J�� T.�����WǇ�W�C&d��Nj����V|ި����q�sv��s9�5DGVm�U
h�)����b�.z؎8�D���u�*��Lk��D2�ٞqֲ�X8����o���e��W�.��t�v�A0Fb�hnJ��.t�ݖ��m�ٛ,}�,�feG�E`����3�=�HJV���D}��T~_�^ rj�ق��[�J
�L��p7����7�v��^�Xd%;��� ��iN�j��G"8X�vX}�,��{}�����r�w縳�th>��L���?\����N1)%�F��r���Tk�iꌦ7����m;n[�n��!,cu��]����}�Q/I h��i5h�@��5�*���F
�PZ:&�[e�${v�nx�q���ڥQ�56�]9�"�$�qľӨhM��;r�<=�x���^��H]o6���s�'�:���J�7=�cHdM;�Xi�L]�:y#6	w���T@@; N�e�o}�[4f��{���ݵ��gc�j��nvX��.מ�OWh.suUM%�v�R�ڐV䓠���ܞ�����}�F���׀y��vJm6����,���W@���,}�,�̖��&� *rn�ʐ�S ջ��G�'�w�4���=�(ki�HU*�8X�n� w'�%l�a��Yw77d�^e�^�y7y�"�Otݳ 7}�������σ���Wн3��a�wj�W�m���1vࢪ�r�8l�<s�y�{v���MYD�ހ��O���`@>n�}�,�mkq�
&���U������]l�)�8'����Y�^� o��ܿn���ȹ����������� |��<�-����`J��6���͠��
�i�[�N��cu�.��@䭘��\��Q[T�A��;｛ށ�ɥ�}�����6�
!unj���I�sU*d>m��:Uέ;\Ӧ���iv�M�vC.���*A�3�9>�ݟ� �3e��fI`w���@�5A�HU*	Suf y'x�OJ�X�'�%lʚhx�i81�U�R�t6���h��ߺ���ҁ���^ i��*���A��� Y���"���:vEM�`�Ot�;�rw��������]���z9�����)T��s���2d�rw퐙IV����p'�gn�%#�CE�Π�C9e�l�#m2��6�Dr��jw/g)��#Z+/-t��wx�N� ��U�op�� z�`z��n�*1����������=��� ��^�;�5G@(���A���vW�w� �3e���l�{j����6 ���a� 2�9��TD7�ͫ �{j���}6�B�?2~ �L ���[�}U痦ﵣUT��A�%�{=���{��������͖�ٯG���)�unG��7d�[���zq1�D\[q�nzp�4`bL\�d����JO��΁���`wٻހ}���\�����-���(��8Bꮳ�!�_�4ܝ�@r�xϹV~^�6w��%!��*����6�.g�;�L��U�o&�@>JS������U3HSUa����j����6��ǟt�͖�b<��F:c��ܝ��� ��߼�Հ{�� �r?������uC�EW?�TE����?т��﷮s{��P(P$H*H����(�(�JP%(�!JS-
��%B �
�F!� �!J JR`�����P���	�
i�
� ��JAZYiQ�b(T
(�@iP�)JF �(V�A�
�fJ�UU�%Q�A�VFUP�QhD�A
@T"@R��ER�B 
DPYX�T
E�ThF A()Q�UbE�PZE�Q@&E����2P�D� �
�-H$��҂�(3*���!J�PP��P
Ҫ�0�R(D4�
�J*/7�@��H��
 �J*<�2T�D���J�P�TiP �T�H# B�J����R��(�P*4��J �R�P"R�"-"P (4%"%H�
� B@�
���% #�-� )(- �J�R��4���*"J̊
P( �H
AB�+�
�
�@�ԣ���0� ��hR��V��:Q��ˆ�w���T) �������������P?� ��(����"&��@��|"?�����".�_�� S�����D����"�P��?��'�������������������������������
��]�������gP&������?�)�ߑ�����Q����s�����_�_�g��������r"������B *�H���{�/����G�C���|��U����?��?���CDD�D��DT���?�?�(*������o���������>�o������5���q�Á�݈ ��?�k��7�DQ�TI!D�BAIPFI	$�� (Q"JTJT �)Q"Q��@)Q"H!D�!�P�VTHE �aD�!D�� ( �@	 ��R`�HBITH�RP`��PeD�TIHFAI	Q$!� �I�R �Q ���RBTHTH U�TH FH�RP�HQ  �Q !D�D�TI$�Q)Q&H%�R!�H@�RT�T%D�@!D�YQ$RAITH�RP d d%HA !UBP�P`a%	D %A��RPd%`%��PIBT����	$&X�� �$!%��a ��@��a �d$I
Ad%$	BBD��P��T��$ T! @! ��B ����� E! @�QI	AXI���! &BYB`&�BXH$	��JB�i�i�)FI �!E��X	���$��BD�`%U�!BAY�%�$IY	B� H ��BE	BF@�Te @��a	P� !	IBUYBQH $	�%�� V� �$���P�B I�
@�@��$HB`I@a@!T!	T�%IT�!`H� �&ZP�P��$�h!�)B	FYB� !V�H HHFXB�"@i@�HBRE�`	�XIDQ�F�@� �aFE��� ! �RdX �he	�i� ��F$I�e��$Y�fE�Q�Q�Q���aa�aR&!%T�`�	%@e@`XFD$`YFT!`YRP 	P�Q�P$A�	�	VE�`BE�
 
T��	�	AV�H�d�	!BDH�V$T$RT!�	P&Q� 3������I������ *�����?�����Zצ�g������_O��_�EW�3�Y�{��������?�֏��G�������PUs��"YTF����>���I��_�PU�?ğ<�t����y�� k����J�
�g��;�������v�:��¢;��
?��������^���xtY����?��?������P�_�u�����t�"����`"���O�@�w��8�?��Y`���o����8\���߇����?���O/��"���.����&C��y���-�k����?�{���EW�������������\o�c�������*V�����b��L��a�E�ٳ � ���fO� �~ ( 
	
 *�(Q  � �>�	�� T� ! P@� �c	lԚ��
�*�(�M 4@ ��U ()4 d�b�j@�R����$� PP      F�ںn� Z��:��9�=��GW{��j��*��t��U7!.�����֧��W��ڪwz�ɻ;���� u���`�
��xfz;Cݝ7�觀�^g����;��w�;l���Фh��^�P �PKŽ��w�R����Z��@�gA�M���H�S��۹�������((�u�JR�s�AK�PR���)@  6P�����19�(;� 
BS�A=e)GK�S�(wO@�^zR�\�ti�/]�@iz�i@� t� ��� ����$ 
�Æ�J��
f���Ñ�08� � {g ��m7X��#�l���>�/g���׽�<5@ a�������Y��-�|}��=�O{ �����=�p��9�� 8�h�����a�0:u{/��g�;�q���wB���x���!��n`u���y���(����PT�l���70<���BI.l���y��  >=���
 �`h 
�w�:u�g���w`t������0	��9.��;�(�p	��2  !�2wXる����9��70t��=�Am�]��������    >"~���IR&  4"x�T��M0h�'�T�P��#@  j{MTSzU*   z5RSm*�@DHCR�� ��=D�����_�?��s����3��>��k�PU~��EWH"��uW��_� ��DU:���_���	HP���VP��]�m4�c$��P� "BI��xhٚ�$@����O=<`h�{9��C�L\�!�!]�yu�D�.����m=`@� �&ݜ��Ǹ:xE�!$����Q��B�# ���C�C�i��L/<���I!0��Qʏ1tx�(�_WsnJwn�"����	H�0�%��[&nNi�l׶杄a��j�ȐZ�4`�.�|!��x!YYni�>kA����-����I��rp>�'�"��<%aR\��_W	L3�2np=O��}D�	d"@$�I�]��5�'SрT"c\|80!������{�L��$b�"V@�!���$�y=q`XE��H`P��"���R� 2I �a�a�)��>5��s����,B ɤ�t�e=���!��'�8,=Q%����x��+9
�))
��JfK�K�e�V�~�Ry���R��u�����"(F�,$yG9�������e�xdff����-�(J�S��X�ۓs���SZ���`��;5�i��B2B��kϴHF���a��7���M�CY�`p�l���S=sK�q���yn������}��L���j��\(��gnB��.@�8�����/��5%�.h�M<dJ�*8F��B����!.�Å)���O�h��db0K�dt�,�ke����~k\��!p%0��>�[�sR���U�L��m�j����t|z�~[����&s��9-�'5f��熹��=&x�!u��By�9����!�(�/7�5�,s���:I�����덐��͇���dH���e�����$,hB�i���t��$B��A��\��SI0	���� �Dh8���v�b$P�HHP�p) �$Vdl
)��Al�:��i)��JO�*]1쯻>EwpU/�*p\uv���Ma�8S�%���a���ߛ2���e.�:)"�����e�� uB��9��y�ߛ%�����ۚ�W�"b�Cy\#t�)�R�`�I	$L�-r+b��(h�ZJB�����1$k��S)8sy�g2���NW79�K���].�(m�$bP,"B�M���6R%-�>�>�i��h�\
����ϻϻ�}�(��P��UE��YR��s����.f<��lᇰ��1��{y��r��{��r^F���
�\S����3/r�W���f�e������
�s���VRϮ��pNV���H�:�I�:�Ԫ�������p���)}���լ%5|o�9%�ЅM1)��ދf�w$�.�q�rK�>�Ω�y���>ϩ�|S������K��O�2�AT�9��i�T��W�΢���_0�T*�Zr�J�,.)Ѭ����0��a'����e�z�66��a\`T�\YCLXU�6%U�!@�XaR)4�8�`hLB,1�$P!R!H�ċd�`P%,B�
B�#T 1	B%XH��'�K!���g�g�L�����nk�6E!
H`1�/�x�@��d��nk|��Xߕ�����!����B{)�x];B�H� I �2.B�'���[�"OAe�.Bi��0�Y2q�G��Xo_]|}�7�5�L[�f3�\5�$�޼2!q��$zgSa�q����`l�-�&����7����B���� HY$`��rȲ�
RjB�Ѓ!JF�\��%1��y.r��VV$Za�٩��0���K�ɼ�o9#�xD�'��e
�Ϻ����~���_*�1哸Lw�Wut,�K�l���:����U���bR^0����)��$H1�K��ߑ���$H�����I7�������ɿ>�;B�V��&�7��N��,Cs�t��כ�]����t�����%w�s�C��|W�*Ő��H�e	Mp����S�s�z]�8{�n�h� ��L�_Z��|N'���H��_<�=��33Yy����~�7v��Q�.��_@��Z]������6�J�]����˨�|�Q>6B�:>IsN�H_7�F����Y3�!g��p}�+��������ܺ����w�S.���Ą#OD���u�s��.�hߍ��).��CI$�A�˓X# B��E#��A�
�#� ��E��"�@! *�
+
(IDlBI`�hF�a���94�?$���"�ʁ�I�[��������X�ʾR���y�{,�7~4b�<`�F���kX��H��i$LY!�iBd3��eÁ�	`Na�d��nH�H�~>���8s)
s
l�)@�M�lhB�D'�|M�R�DA#쑦xC��_r}�7z�'�h�D�aXa�X�Y��3 �,��BCqf��H��@��@�!c�A��܎�S�!%��`Jy�E&�$ui�/�E:�y��.�)]$>._}�;�>�:�1*��Mrq�O�`L���H��L8�ۙyg$8�
a����a�ӛ�ͅ�����oL`�	p�3\6E����$Љ�9�c
|h��M{�Yu��
[+��R��2�v����S�Y}�>>;*̎�P�s���_s��"���_��/�7��bk�䔺qt����I�!S)
fM@�f��1d`T�Ն�e2B6B-33������Nk��sgQ�
_kj��V��P.>bu)�g[¾��|e��|H�J}��Rݞ�ΩI��)}격9}]s�����*�B��OIp�Xyt�Y5���s�>�9�,��p����\���3z�eaYs[HVBЅ�S	#I#cR.h.��SWR-�	\b4ăHi���cB!,0�� ��a��H�-GL�H��R@�D�$H�0"�"���Ŋ���
Q�$"�a`"�$@�C[Jf�P��"B5�H�"�Nk����1!����!Iy�BHhi�(� 0`Ƥ*�H0�(d[�+�AHA�OM������ۘ�_(�G>>t}EP(u3s+Y�g.�K�!cJa@"P�H�~T!�eBcVXi�0��sl��v�y�=��1$$��h!fk[��{�Mᆝ���6�
C�~�
�z9�y��[u�5Oi�7����u
a��7��=��������Hp)"����>����?�.��Q�}O�<���T�^'x}���>��w�T����ǒ�,̺�d���"D!�l�*�
�eQ]W���]���Qt�<�XE���p$��y���4cߗ�h_1��� �&�A���,C��a��񷥛�4���"�B0"���ZDJ�  ������'�3�	|��<p4m�!F�B�-��
�:�|�A��xT�n�KĂ�sLk+�d�i۳����b1 A"����=H�y��N��O�E��Y,HX)BZ��|l> �6���,c!$dB�����|`D��r�

��Y�X���,T8'�8Bs^N���$Í�l�oz=�\ɳЬB9�)��ON`i�vd��0�Cn���6����7gƍ����<���f���2_8s'>�Jg�)�y���D�.�B� X�H�Q���$crHP1�����+���~�f�U���s�.���Èl��+g��_\�R����E�.�b��㖉}ۺ�_
)��7�͓f�9Z[�fd�3z%ѨI
�`@!cB5�HT�ڒ�kp�,шF!��$��c�1�72�s�s4y�n�u|޽����2�Zx��gN�˻ϻ�Ν��s�Gp/S�>�����0�.!r%2���\��s/y�8�e��f�#�j�h!e���Ox{�򏇥l� �y�ɻ[����Y�{ﻆy)&�I�4��K�{�o����V��(_	L*����2N?���@g������<˾0�*����`��D��np��9��h��n�͆�S!F��4!R-#@�60`F�b��� ��FA�X$I!h!a]��B�E�hܑ�,X� 8��0`�E�EJ�$Ġ��$lX$K�A���)p���0�1���*T���o\
|g<���X\�=9���j��B����Zp�w���ܧ	��L7��=��(��զ�
ੇ$|/S�U%ھ�[��������]VEܧ��k�B�+Zњ�%�����HSg�sMSg���h��".�][�'������1�9#!!"z��F̒Kg�.K���e��	�Ұ�������$�0!5���
��a�9 ���=���  H   �                                ��m�  p8 	�   p         � 	 �`   ��      Y��T��DJ������"��@���,F��nP�?�l����h^ݰ�m������u뜃d����S̮˸�^����	-����H���Ֆ��m�$UpWj���l;aU�n�8�½��X�{��9���k�35:�|��?+V۵UA��[�dFn���ٶ��'5�:��ˋ�b��f�����[\� ��r�8�M�G1��5�p:�g����#��U�[+�Q��J��� �mךL-[��p�m :Y�c��7M���kn���@���mm�8�C��`���Z���V���eUj�� %皪�j����6����l�m��J���`�m&�  	/Y(��k7�I�������fܩ�� 5����r��WI�5UR�ҭHMT>���A�ҙ��
[@�����i2x[v�*�lIe�W*�\˪*�ͶNM��q��6[[R�n�nj�9`jږ8��f��1��9#�J�Z�=���P
���a�]��@;�ϧ��k�Y1��ڹn����Ep-���Z	 ��)�ru�b��Z`l�WGWT|�9���Q�mk��%���XD���*���;������\�z�1v�	��4[mҞTz���h�nAݻ����UuR��^��ȅX�����	awm�!�[S׊x��-�dq��"��  ��U�V�tk�AP����)@YV���X��vp�D�nz6�J7˻?+��>�����G-���-K�Xlnٯk(ݻ`p�N�ԩt��� U2ʻUTn�0�*�cE;i�cl� ��m�tW0�ⴃ�z�d�Ɲ+!�դ��Nf�UQS�zY`�pVa���'����ꌋWmO*��]]r�W*%�f�ڠڝ�m�n3�p��j�V���V�F`T��.ʀ �&�l��6�K���K�V�Bv��p�OV�L-�&��dL��r�EU-�����Q�>ݞj��X��V�W�� �/�qìn�ڋ�-�mϤ ����Z���Ⱥti�ʼ��T�QѬ6�2��@T�*�T���bv;��l���Pͫ�o��7��m�i���s��K��In ���.�שÖ+.����0Ԫ�4���q�;`�nι՘H��mjIA��]�T9���P{5���6 �-�� -�1����ҙ����#�W���.��nj@� d%���m�Kn�	�ʲ��jm�E��B�ҙ8L�j�"dv�.��'0\i��%^���;����춝�z�ŵV�`z�4�Nv�*�']p��j�ɸ,���7�Om��畀U�uI��;U�L.X�˱��v3ųK�C��� tW"^7�i�6{W_A��T`ęD��/����%�g�U�y�ݰDl�=v��MC[��j��m^m�6�$.�'6V�גĳ��m&�  �+㜅�����V�=O��z�4�*��m�� ��i�n�	f��O-�f��  m�����m�pX6×I�@#m��-��Tub�K9�m[���8�,�l 6��h��Z��ݦ98�UvZ�[m�� �� �  	eH0�L�J�P�y��!��AͶ	e�'k[�;F�t�`�˯�8��)�ܶ����������6ض�i�6�   ���� �m��V���p�mu��m'n�BA' [A���ۤ��p[A��lq [@-��	 �6Ŵ��m2��UT��L�V�V]��4�m���q: 8n�@��(  $     ��d�l�p�� m�� ��jG-�a��9#���c5���n�o��Y%�}�k�� UUV��7	! ��&�m�[F�m��� Hm�$m�� Hm�m�kh lm  ln�m� -6��� m�  �&tRɢԛn�h n�G�m��$�� ���'�%}Յ-�ж� 	 6����ko,�l6���u\�J�m����  l$m��    � �6�U���`��h��0\�[��*��U6�]v�CNR��`��۰	 KlN�-������ �h (U^mU�&���E���H[x � m��h  I��ѶƵ��`n��kKv��tnZl�6ؑ��H�m��%�*E�pB��hH �p  � ���l��  *�5�*UT
mPY`+j���N`�/Y(��I�T���9�w5�5UT   m��m� �m�� $ 	 �  m  p -� σ�-�����l�K���}8���ͰH	��m��m'�WY7G$f�;E��� ��`      	�������Pq��kY6�����Y��a�[Kh    �     l6����GY!�֤$ r��:�-�H�m��
�T���+!r�;Uf�p,GkD�m    R�Y˭�.����qZ� UI���L���;V����vv�j��|֚�-�ibbbrA�"�2*�7G8��G:�Aǩ@��s��I�%Q�s�j�s�+��A���N��m�Vګ�N��9ylGn.�6ـ����)8��y˴;t�/k��UJ�UU��ʁP�V��-��]n`RZګ�ejU�.��Q�Ō5gp[/
��pܯ ��T[�e�c$lm����Y-��3�[v�����A: m�N��Ɣ ^�6�PA��V����_�/a�V����p5[mQ�����˽�	���ֲ�ģU�]�]���k7������-R8j���� H/[,��2v��l�^vݬ
����Mp�r{p�l�⫆�+�9by��ڢ������{��yV2�.��9��W�qJU�j[`��d��WhڳpfҖ9h�W�.Z�D�{B�G=��B���E��cC;���\O\���V���ۍѧ�[!C���R�64 v&69
2��ֆ�L�2�ux�
��(M�"�s�ݮp�<
�J؝�7%d��v��XJ�7S�3�İ�3eb���l5،,8ڵ��q1v��9,ͱ2Z���[5Ǟŏ8�w���wl���e�6�K8�!g8Cf�g��%��E��2��j�YWm�4V:�^�Y5���Z���{p�8H��±F6�V�ca��Ss��Ի��$ �R�����2��UP�cW5 T��U�Ôp$�Z��  �kn@I&�m���a�׫l k�  7l��Q��I�m�lÜ�N�5$M���ċn\��}=-tD�m ���ݫY���-�P�8ɚ����n���Q��U���g�&���:e%)�\l�V�<��V�E7C��z9�v[ l�6��m� ck��m ��&h-�I� m��V1�`�V����^��� ��~�| l m� � ��U�Um+� v˖���J6�ms� ��ے��6�[@&װ	��ZmSlp���$�Pm�����Hi�G_���m����	V�$�T+,�K�cIF�&� (��Lh���6Z �E'A�� 6ѮK�++��S˳�XUUTIkp�ݻsf�Ë/@!�4E�\`ͮQ5��w$�m���ms�<�`�o m͖�mI ������z�-�6���~0�����ۭ���kh��mm$�  H�9�m&ٶ9  �m�7m�,6[@7!����I#�p�lƆ��Hl�(hB˙����$k��#�����rÈ���]��ҩ�@  ���H�ӶΧ��I��Ih6FZ��ܐ�ظ[V���Z����}o�w�L�hHd[���p-��p	5�m�� Zl�Xqm8��۶�I�`pاIf�5°�jUUZ��UU�f3lҬ�p�6�X"�5�u�Hh�	 w�����N�N������T�vUjV	�3���S ��g7*��H 㶩����d�"�j��-�d^�Hv��R�$5���r��k��	{K��,7m��mm�  �u��ڶ��Z ��6,э�����_������ed�;^��R�n�2gC��Ŷ�v��Ļ@ ,sm��mp��z�l.�km�9��m�	��6�7m���:F�:uU��$4�AL��ҩ&�/Zs��� �]mNu� [m��l�� 9$����ݣ��-Λ�m�6�/R��mI�.� vݒ��6���&ܴ ?�7�2��9#]�� I�Ɗ£�h��-��6�  ���6��j��ـ�몪VIk�W ۵�u�  	V��I�^�_\d��UzR8$8v����@��� ��8��WlA&v�,��8		  ����	p[�m���m�m	6ؐ�P�Hl8�u���p����w���yK��!�C�S�_�6
�� O��Ep� H	��B��i��l�P8E��! `�ߊp=J���#�k	�*�_q`��<AOA �@� �iT+�] �/��U�4(�b�)�4�p��;8�6#�M���KB`F2��_W�@� �4 DpP���@D#�`�}�t���y��S�b�ϋAx����Ҟq=}M�����q@$bEY@� dO}�'�<E~DHE@>L�OTj�cH�� �H$HA ���}�����/> � )�����V�|"b @>���+�	��A��%Q_��xP����V*��5,�A��H�(z!�@� �lI�#��� z(}ChA������L��8��]�b�bA��S@|�`DU"AA�1�с��@<��8���U�/�h� '�
�`�  �}qУĨ��FDW�O �8�������_S� ���ʴb�<6}����]��#���x��EZ��b�T��P4'�mjA� ��J���M�� ��}|*�BXH�"��$J>=���bB� �������p}A���Tһ =�=CB/� m�A���BZKYb4 ��P��R��bYe)(� 5�ZRQ����Yd��T��ŶZ),�HB�Q$ F��R�"R1�B� �����VRX�zBz����hv��BI$ �0�B2H����	���Iq�j�@�����a�@���F1�I	l>J���؁�ȵ�����`�Gj���� ��G��h?8L �`���!Q"�dbq��eJ�A�B�4��������     ��\�i6 z�n�i��P�)(��3�Q1pl�c�64�ب�1\g�B����%֥�kkV�r\� 5��5ͷ����J󲂼�f���]i���hMI�n-�H�h�&IZͻ���!r�u��r�������9lZF�Q%�A!s�4�4��Q2�����,����� @��Э��ZT%z�c	*�2K��n�"����&tK�tp��p�ov����vч�mm����4f�T;sn�,��E��.�+������nX%Cf��C���bF�����9� �x��y+�xW�ڤ�ј|8[�� "(Y	��K�v�\�#�M��-��l\��m��s�@J�6]�ڕj3�9����
!*KTVpne|��f���J��Y3l���smP޻'�`G$��/- �J�t��*�O��]�l��\@9��.�V�nݎu�=��qr��R��5�-HL;�F��ΊP2�J�vb lH�1��d,]vAns�q�Z���8�1�ˣ��\�*�UT�-ǅ5�RAJd�51JpuO-UE����`f�qA�֑�u
��Tw���+YP:�b;�ڛ���1���	��[��e�l��m�F�&�8�s�c��2�5mI�\i��&G��W�mQ�bP[{^�*v��c�[�C5��54v��qGm�،)dy�ܢ��yI�m6xZ���^�$5،�� v�0����%E�.���������B�%]����*ҭ,��2�Uv��'7M��j��b5�1V�V��*�9�޹Jx��H�L�j��c�V��%�4J��8-���I��b�����٥9ѳ�4h4=К�ڍ������b�We������ʰr�L�n�N�U*��۫m�V��s[]-�:��Zl�BC��;��5�s��vEQ��j�2�[`�6���ga���m����:�ў�������|� E�hTz|0x(ǡ���P|O h�"��.$�N�t{�����UTqe7g2QT��m����˭;�����N]�܍40�F.�`���Z#;k�tD�l\w;�q�c@����c�Bު�+��9i�6��·�#�v�:�����,���-��\LA���y��f"8g>;F�:R��n^��hM͘v��XЋٻ@V��U�V!0�v��k�3˷?�$�����o�^E08ݔ�{��˸M����{m�"<(�=�a|�	��:le�"�|�u��� ϻ0�o�w�|�Ƿ�&�:MD�Q�����~H�l�`w�|�]�v����oP�PƤ��&���U�����3����;�5��i�#���>ך�]�v.�{�K+��cI�R�������>��`ori`}�5X�r�{�1ʈ�>Gr����^Â�^���ks�=�i���s�����g�T)�Sh"I��w},�M,��Ww]��kݥ"�7"�Ӻ�nI����z&�+�@��B��XE>EĲ���ܓ�����N{����+tBڑ�F�m�B��j�5w5��%ջ�`{6x�1t�I�H�p�q	Ȭ]�v�3]�%����>��^�> �;�M;b�Qw�$�^��Ine���$c�R�Ik������Ϳ{�ԙt�,�Y��.�r1[C�X;tv��3۠�Ĺ ؼ�i�7.����!C��ϒI{v�}�I�T��Z����$��m��K�wh4��ӀG	!��$c�R�Ik�����ݶZI-̾�}���N՛�덖jl������r�|�_n���>B���0�g���g9��7��[l�=��v�xzI��ڃT�����Iu��-$-̽>� ~ߺ� ���{��m��5�Dn���������Ic͎�Ik�������7����h1���nqH����-�VƌEd��I-Z�;J�$Rы����"�} ?o�w�w�{��$��n��������%��I=���BA�'$v�K_s_�z�U�r��F{�R���������� ;���X�	�Q��I.��i$��z}��)���� >߻������^K��Yp[I%����H׺��������*�}Q���NC���| ����c6��{���G������@��� {��w{����L�(Sh�Y�ЎLqmѦ�zN=iz]�E�Q���(�h�Y�6��l�ѭ�G� �߾}� ;ݒ�Iu���W9����?yKI%���5�F�ص�W�@��� o������w����}����������r�Iu����Kwd��\�mf�Ͼ�S�π�տ�J1q6�s�����m���� ?w�} �{�� o�����_�7fF�Ƀ+� ~�_} ��}�} ?n���� �z� Ǟ�%���74�{[�-l�2м��FŹ��̪c6x�v��]Vy��[.V ku�흝�Ԗ�Bv�(M�@*v��]��J�8���DÖ��"�e]�)w<��ѧd�@H��:��ֽ5<N��U��<�nx�7]ż�õ=���#n�6ER��V����\;s�x<OW1�]���v�X�	��pV��	tkV�G.]q��N�9��t�,�ͻTL��MW]�x�FW6�����=�����/:�j�
hB��0;�1lnW��S�}� y���$���-$���ϾI-Э�9Cw@��$�r�Ic���߹�m��ޒ���}� ?w�� ~����������@)��π����� �ޯ�������~����M�5������9����>� }�� ~߻����-$.�Pm������@rO�I!n떒Ifn��$���ZI%�ݗ�Iz��I�~<�ɥf�B5%ڜ.�nFiStֺ@��<�E�=��3t�RQ��s�;߾}���s� w�~�r`�_ ݭ�ԣlMf��[l�}�k<��k�5C��nHlt��/<M���k-�����Z���$��ݟ}�r�kɛI?L9ss2`�| �}��z�< ߻��@)��> ���鲗`L[���>��$�}��'������{� ������[�B	.1�� ?~�_} ���> �{��@��x {��нi�L�FRjYs�hb&����P&\��͕�PF�@9�ϖ��.�m ���{�(�����$n�%��Ǜ��B[XIOxӤ��A'$��K��>�$�٤��X�5��I%��ZI/�j���M���[m��}��m�������TM�,���rߜ��]�߫�K�o6��!�#v)�� ��~��Ҁw�_ {��}�I�Ii$��3DG�����_} ��� {�����{_ ���}��C�Yy�Y�bd�x4��Bb�Ti�G]��cN��!4�;2�5��Ke��-> ���{��^�� ����H�۩i$�q#\F�M���޽��m��{����> ���{�{l������vk� w3g�$���R�I}��W�$��4��I~�{�h��u4B���c��> }���-�}��5�o1�{ �P�L�V8�]�&�Uw3�o�s��g곱���6�K�> ��}��$��Vm��|�If��$���夒�J��t%�x�ML;,UZ�q����.UM%c1(��-��!Z��f�h&]c������%ܛh��K��>�$���-$����=������Źr7k����fk��n�i$��߫�K��Iw+v�R�96�{�?w�� ������$�v�i$��5��IcfROjFܷ3%�s������{����5��Iw\��K��ޅF�M���[�p��^�ɻ�ޤ���9i+y���s�����YbH0�� ���k�m����h�W�E�d�3���T݀��Be�̺��sF㩴�H�'�{Yo@��C�g����D���Ő�KJ69�m�U:��΍��e+���{QJ�ٹ-�`E�b�A����@�n⌔�q�l��WDXY�,��Ɩ/���_mi��4 ��b nx[X:.��е�N�C�I,�Vy���]BeR�J�����s�+��q6�|�'���j�Z&:{m��0!�]��׶��!�7+!w��?bq�k>�Ec��D[��[��������RH[�夒�6���[�p��K9��j���h�{�;�������RIn�Ձՙ���鲶�I�rSd"I�`}�4�7wn���%�w��=���>Z��S�22�D�$,�۫�3]�nn��٥����u*A����`ufk���`}�4�3wn�Ǐe7"H�Bq U qS{=l���/m��O����Fi䳰��%�.�lj�=2mƤv��,�f�n�׹��9�[�v�ͤ��F�r�CnK��}7�W��0@H1���J���I�����=�{�n��,���
�J&���X��VVf� �ݖٳK��G,RSR�B"����v��,�f���Հg3v5N7#�EIH�svXf�,�۫�3]��U,�x{vZ����m���!8���mJ�ֺ)S��7F�\kn�k���J��,t_��O�6�����`��`|��[̈́j2�D�$,�6�����`��`}�4�s���)�Ҕ%J�IGr�[�v�͖v�8�VQU��\��|��W�~M�H.i��[N��41� �T1%�5��sqOp�w�&���M�5�ӫ�n�L|�9�cxR�2f�D9�ʩ�gO����ք��!��3=Ĺf�-bbI)�Cc��)D29�8����7��2��~��CP���uu�=4		=ɽrߚ��,BFO�<�ksy����S	s[P��������|u�BB�U.���fC�kK���M�7���k�y����'76�G���nsF�!��0��3L¿?,9�c$=:u�0���<�˚�6
r�d6C[�/��I�@�&��l*ľ�}�X��ܼ�<��7��H�_p�z�q4 �l4�����@� :Z�� )��CԪ�"$B%�m	�@���DP1��P�� D9����4A҃]]���Xwv����$IEM�Ԏ����Xf�,�۫s����{ߝ����I���A�q6���٥��W=�����|��۫�*��(�JI�Oi�fR�#e����� ��tۄ�ݗ�T�9q4F�����4��ku�O�~�u`ufk�37n�r���ΰ�~��7�K�R��j*$�`ufk�s���Ձ���`wwn��+���M��߿B��F�'R�%#�=�߮��f�{�ĳ}�5��%m�ے���ԕa��R���X��Ձ�y����U9���8�Z&�0M |i�R���_�M�����}7$��ğ�����9NHX�۫��ʪ�~����t���Vْ���tJj65�i�s��q�q�$y�[2�Ge���6�R��>Y�0k�����o����X�۫�٧�ϐg��4f�D�q6�9���u~�$wޞ,�z���y��r��Sg�O�'��n9)�ڒ���~,��՞�Ku��]Xq!=EF�MU'!a꥞���u��ua�]��Ł�Х�,C�C��D��ǚ�ܪ�+�s߿~�t��~,�۫�w+�9U��\�HI�>f�0�m(^��9����C�9����/T�P����s���g�2х݄�Sf���&aH�l/A���Yx��lZ�	\\m@���@h��g�,��/;j���Z��[��鸆q����:!��賎��q�� ��J�ϭ���H�vv����hQ�P��4tfMCM�7�]�b9�5n����kZ�e���a�P����$'���
�2B���jx�2���]#4Ӡ�T�ݪ�	�1\�����b��Qv)te"��߮��f�n�׹����+Ճ���&ܔ�U�V۳K�8�����׾Vn����T��hW�#����)�w޺�3j����_���������ߧ���
{��%H9UJJ��URݛ�`o���٥���\[�{�3F{ԉ*(�Q6�9���u`~����s������@��߮�ǚ������6�e�Q�2�F�*�3��.nq��t%Z]�X�.��)��wH������r�LrW�wޞ,�۫1�ܮU~�*���߿~���!?Ȩ҉��r�{��lޓӊ|M��Ti���C�yX��Ձ����r���UU��x+ߨ�*r����`f��Y��s��OŁ�߿]XVf��m�IԥB�Xz��}�}Vw�Ł��ua�r�l�+Ճ�y�ے���9*��6i`z�}�}_�w����۫�9�U,�w}�Ԩ�6+l֎�j�-ڂ�	q��1��Yb��CW����C�tQ���n�M������Ձՙ����ۯr��A���`wJ~�DRTrH��%XY����RF��������ݺ�W)#)�G�n(�u��{��`}�4�n���f���Z�ִL�k>E>��G���wݛ�{~���'���+�F��r�CN���8����޺�:�5�z�\K}����y��JRh)97v���9�s���W���l������銜��(��)�6��hm��3��W��aQ)�6�f.H6gT��1����#B����I�Bb�W@��~v�����6i�Ur�� �{�V���?P�j�Z��'�|}��Q�
fO{�_���߿]XY���U�r�;�:��M�)��$�I`w}<X��V{��)/k���o�^��B�P�Sh�䅇Ao��xnI߳���O~��[���~��\"a�ڀH���=P:������g�{^���*�mIV��V��T�ޯO���y���V�=��i����.�\��\���
g�crJ6�0��Q�:oӤ��Rx�vR�f���W�`j��`nn�{����=��V��н
���r�CN��5f��U��fO��훒~�~�w$�y����[d��B��D���Tr;پ��7��s���W?o���?/~�����,QJ��t7J9V�U/l���nmzX�w7'�D��g����rIӽ����&X\�I��`ܭ��s�_��W��ߟ@�����՛����9�PUsy�+�$�*~9cJ�א�m��rh�f�����0d�y�i�<]F�f䝋*I�`љN�F��ȏR����j�{:�[�Ξ9\�."jfv�-�hʢ���i�A��3�b�Ү�Ev��i��\ҼQ�U&"+ab���8�͞�@�$:uN��ԛ��n�x����rn�k@�	��4��0���{y�v�����s�H͍�ђI����{9�y��Ŧb����$��*Je`��CXl���X�Xml ��@�M?N����u�gM�n�����v�ݺ�5f��W9_ 36�,#�Z�T)F�%'#�>����U~�9M���~v���,Y����*�;�?W�G%G$�����}�`�V�=U�%��;��Ձ�F�"�AF�t(�?
~���'��߳rNy��7'TQy���~�z#���8��I`j��`z����{�W�yo������u��i�&K-\�i�b��n,,e6�%���ū�˗HV�Sis���Ns��"Ro8��h*9�w��Vn� ��l�*�U_ ��y��o��T�J��Qʰ>���n"����V02SY�%�VCVFL6�Jh�qC7R�0��a5�x2␈.��B`ׁ�aT(��}^��2X��v�ݺ�W+��$[�C����JM��f��`j��g��UT�s޺�<��v����6$��⨒u%��ʮ/=�������[��=�rs�;ޟ>[~/e��ѳ:ٱXe��ݺ�?UW�s���?~���y~���vwJ���p%6(�$(lT&�ɯmr$��F#NJv�e�o2����MPG��N9�>GhFI�89+�<��; �Ų�ջ�ܪ�9��u`e#ը�H(܂n��v��e��r��W9M���ߝ����Ձӽ���s��{پ��1fd���$��{��s�~ٹU�� EB)��"���b����L��&P+�OC@B�r���?/�|����Xueҧ �)4�����U.�}�X^���w1l��+��^~����W�%J�T���`j��`z��ž���^�����������>���5r����3�ܫ�r:Jݱ�,�m��V/km�hozwN�����	Ԥ�q|���`j��`nf�z��_ �����>k��t�AmI`j����r�\l��~��?~�+ �Ų���q#����q��%'#�=��ٹ'�g�]�� �� ̟�v��䟯�߷�|��}��p�T�Ug���"�������`j��au%Ps���r�"H B);f�S�ͻH:u��5]"q(|�
�UW9Sn�`e#kQ^�Q���X�-���s��?{��=��u�-��ýYx�3fh��+�m^�nS��uqs��e���˩�f��wI�&��G*(Ӕ�jO������۫u�ި��O���nI>��I���.��*9���u~��s��q#�~������w]����\��ҽผ�*D��(ܫ�~��[,�Us��K���=��Հefhڐlt��Ri��?W9_�������$�~���}��lܟ�_�<�������>y�@����"m�,[������*�{���@�����7V��a�M���Q������7�@���U|G(�o�<�_{!�Yxe�P���!��$�$���0Iad��$�����\�"�j\���y�T��X�#��utHq	fY�`�'5�! M`���$�$&�����`�!�t5J@��Y�b}�%ڦ ��dU�BR��H��0dB	��<�">���$�Ie%��$e�Cp$�&�$ B��<�����MkZմ     ��itٴ�  -�	zW:�\ґ�P�6��A�WG&��&ܥ�O9ȝWT�unl5��D�e��¸�7� U�Q��h�Ƃhʯ�:l���.&�2鹧Jv�}�ۋ[":K���� �Fz�s�ni�+t5�4فc)�����4#E1V �gv����|���"��hGl$.#Hi��"�,&��[������f�0ruͭu�$2�f�./0�<��U�s��-i�,�x��vwd���s�#7O��m��2"�ˮz�b�g�ܦ3淂�8�&(-�� �E����-5%�\�����C��E��]+���"M�e�<e���U�r���g� ��X.s����_	�E69��/l[p�`Z��!�<��P�ɩ�a���̪9S|}���J�啕S!���u�wk���@�X'DFPaבctmS�6v�)�k�VH�H�UYh�K��9��ڣ\h��WTr�IO�(ܐv��O+J6E��u���\��^)V��4�j�VV��Q�7=V��>�M�Z����ћ�E����f�p���(vl��Z�%�z7ID���tm�"��zwg[��
���\az�db�K��@�+���_Hr�w#��r���H�l�T�0�D�X�M�����ˌ=�t޻.j9��zbd�8]�2i��i��̭���u��$��zfaG�lxU۵w]R�-n4ਖ��Y�i�ۮ �����n-=C��ݱ�V�\�B�M�[���� T F�q:�q2Y��НS��[K�)[���;J�+@=��!Z3�tR�<�뤹��Ve�É��j��\����e���Wf����K��m�-����niX��GlP��-vlnY�����֪p$���s���#n�nZ�L�m6^IJ8s��Q��m1WT`���-Q����l��AaZ�e�v�[t�P���I�U*f{<���?C�?&��.jf�[6n����}�ğ�����
�A�PS���L�@t.Ө�����*Q1x¸|����|�g�gt�(�ˍ��da�+f'C�e�2E���b��S��1T�6�,_��:л�L�ӓ\98�p�)��s���6���h�m`C�ifɖ��mmj��{:xl�ԕQ��;[k�%R�t���!q{�ݻ$`F�9�_6%t:XVT,Ŗf��q��[J���ݢ9(�Z���{��5��e^�gp�����s�rZ��	sg��n�֚��N��Iݺ~��#��џ���z��F&R賉��˗YVJ�1(Ƭ�B�!6�I'�7��B6�I��߽����{��3ul�+���K~>����������w��W8l��m9ı,N�]��r�b�"X��������bX�'����m9ı,O{���r)bX�'�N�o� ��Z)�'�����/!��;ND�,K���6��b�ؖ'��xm9ı,N����r%�bX��{)��fJl/���B����;��siȖ%�b}�{�iȖ%�bw��fӑ,KRĿ}��m9������6���1lr�9=��K�����"X�%��w��nӑ,Kľ���m9ı,N�{��{y�^B�}�&� ʹKuk�1�sy#ʏ]�g�n�љM��8�R�&�_:N���|���hW3Ο��N�����iȖ%�b_~��bX�'���6���DȖ%��߿p�r%�bX��{���j�ae�E�sSiȖ%�b_~��'�Bq�E(�2@#"$��!H��$B-$F�`!;���E�'3�y�ND�,K�{�ND�,K��}�ND�c�:S���{���et�`ݵ_:|8�,K�����r%�bX�w���K����fӑ,Kľ���m���N���}�}���P�Q�.�9ıT�>�{�iȖ%�b}��iȖ%�b_���m9İ?E��~��6��bX�'�~;��a�f�j�C3.�m9ı,O���m9ı, /��f���bX�'���6��bX�'���6��bX�'�k���h��2�\�k�Vaa�.;b�\Kc]m�䦤,v�j�]�F'��&��[����bX�%����ӑ,K��;��ӑ,K���w����<��,K��o��r%�bX�t�I�fk5�4f�˚��r%�bX�g{��rؖ%��~��"X�%��{�ND�,K���kiȟ�"&DȖ%���'���e�#�y��ҝ)ҝ=����iȖ%�b}���ӑ,j����M�D�K��ɭ�"X�%���﷜��B������>�����.%�kiȖ%�� ����~��r%�bX���~��r%�bX�g{��r%�`D"�'���M�$R|}�I/M\�Yth�.�lI�=�煉pI}�}�m;ı,O��y��Kı>�{�iȖ%�b^�ٗ�L�i���j=pMp�Ͳ�G@N�E�rC�0�:��M�9��w7�;�-��a�m����ҝ)ŉ�w�ͧ"X�%��~�6��bX�%��Ȗ%�b_���m9ķ����-���[a��.���^B%����6��%�b_���iȖ%�b_{��m9ı,O���m9�,Kק�30�W5n��5��r%�bX�����r%�bX����[ND�[��;��ӑ,K���w�ND���N��ϥ�Ob�K`*���ҜY�X!�3�w��ӑ,K��?~��ND�,K���m9İ?/T"�*��
8
����p@=BD�o�5��Kı;�п�nW\��\��>)ҝ)��w�ͧ"X�%�� �����6�D�,K���kiȖ%�b}�ݜ6��c�^N�o~�fٔ5͕NhGFk�a	�8��le���^zL���q�Y����w�^���!t\��k6��bX�'���6��bX�%���[ND�,K�~��D�,K��{�ND�,KϡӼ��h�n�s<�������;߾|����"dK�w���Kı>�߿fӑ,K���w�Ӑ[ı/��i�.l۔c r����/!y������r%�bX�g{��r%�ؖ'���6��bX�%���bX�'}t߻MftSRkF��"X�X�g{��r%�bX�����r%�bX�����r%�`����vp�r%�bY���@�.���Q�.�å:S����ND�,KʤS;���m<�bX�'�����Kı>�����Kı4��1"A)e6HIgG����Uv����9-�a�G�j�h0v70q�t�7�a99��Ost�V3a8��Q��o5�fLe�׭�paX6����jI�4� �a��[�dL\�c!f}�k���k��˴ݦ���g�B�ݯ�鼫#�1�/Z���j	+hA��&�V��@A�nj5���u��CÄ�
xk���
кl�V��e�T-u���h� ���̙Z?���$�������y��A��t�ee�lY:�#f�t�,
���;,�v�:�Q��=�y��v���RgU�t�t�Jt�K����iȖ%�by�zp�r%�bX�g{���bX�'�}�ND�,K�ϥ�Ob�!he|���N��N����iȖ%�b}��siȖ%�b{����Kı/��u��ı,Oݏҟ5L�32L��r{y�^B����6��bX�'�}�ND�Bı/��u��Kı<��8m9ı,K�i�za���d5��m9ıF����iȖ%�b_���iȖ%�by�zp�r%�b���w�ͧ"X�t�O���{�B�����t�t�KĿw��ӑ,K��( ���O"X�%�����m9ı,O~��6��bX�'��ҝ���sD��ZÝY���}o�s�WoU��5Y�%pv(;�li1\����Kc�	�1�9|�����/!y?}���iȖ%�b}��siȖ%�b{���ND�,K���[ND�,K��C��Ik��]#<���N��D�;��Ӑ���KH�ρ���x�DȖ'���6��bX�%�{�m9ı,O>�NND�(�"dK��g�]�]�\�Ο��N������iȖ%�b_���iȖ+bX�}�g�"X�%��w�ͧ"X�%����}�;E�ͩ3��:|:S�?q!�3��~�ӑ,K����8m9ı,O���m9İ?�ȟw��6��)ҝ)���=-�~F�L��>	bX�'�}��iȖ%�b}��siȖ%�b{����Kı/��u���/!y����녉�m\�PV�{yѷv�73a����J��e�R�l��y���)�T��9&�g���B�����}��r%�bX���xm9ı,K�{�m@�Kı<���ND�,K��g�������y��ҝ)ҝ=����r�"��L�b^���[ND�,K�����Kı>�����@ı,O;�乭�֬�u�6��bX�%���bX�'�}��iȖ:4����ȡ	��b!�"��Ȃ�"�E���I		����
��@5Q>�����Kı>����{y�^B���lWCr�`_99İD,O>���ӑ,K��;��ӑ,K����iȖ%����;���m9ı,O�����Ʉ��f���"X�%��w�ͧ"X�%������Kı/�w��r%�bX�}�g�"X�%��G=����5�ZE��W�XG����OD��ý�V���8�@���m�t8��ڰW{��y,K�����iȖ%�b_��u��Kı<���^D�,K���ͧ#�^B�~�����*�]fp��Ooı=ϻ��r-�bX�}�g�"X�%����fӑ,K����iȟ�RdL�bw	�v��~���Ԑ�ֳiȖ%�b{���6��bX�'�w}�ND�,K߾��"X�%��w﷜��B������>�֪��6jh�r%�b؞���m9ı,O~��6��bX�'��{�ND�,6��N���dO{�'�ӑ,ay�}�v}q������Oo!xX�'�}�ND�,K���ͧ"X�%���vp�r%�bX����m9Δ�N��������lYs��.%��{aÍ����,6���Ӎr�[͚�0u�:	V\�Mf��3F�Ȗ%�b}���6��bX�'�}��iȖ%�b{�wٵ�Kı=����r%�bX�����e���.�[�fӑ,K��߻8m9ı,O~��6��bX�%��w[ND�,K���ͧ"~I�2%:}���v߬�Ƃ�g�>)ҝ,N���ӑ,KĽ���ӑ,ș���ٴ�Kı?w���iȖ%:S���a�]�9�-�fT�å:X6%�~�bX�'�߻�ND�,K��g�"X�%����fӑ,Jt�O��Ͼ�ds�	1�_:|:S��b{�����Kı>�{8m9ı,O���6��bX�%��w[ND���N���<������UYM�̩vmN�`;N(����m�����f�Ԇ,�F/;��J����*d02�n�y��|�65��������5[�n���fO:=:���7��R���K@�o:6�2��HZ�)������N�9�q���M�*��T�,�ܩ�ѥ�fiI�ێ6��m��D�p�sAӶm׮�7U�\ ��ri��e6s�'$�9$�NOӓ������1�A�30�F��!�]��-IU�V-���ؗ��Z�����g��x�n�l�:|:S�:S�������r%�bX�{��m9ı,K�~�/"X�%��w��ӑ,K����ҟl�iV��Oo!y�^N��Ϧӑı,K�~�bX�'�߻�ND�,K����ӑ?��S"S�����u�=Yu��å:S��{�����Kı=����r%�%��{��iȖ%�b}�wٴ�Kı<�:K�F�ղ���kiȖ%�'�߻�ND�,K����ӑ,K����iȖ%��VdL�������N��N����~ڎ�qX�Uw�r%�bX�w��6��bX�"{��m9ı,K�~�bX�'�߽�t�t�Jt�O�޿�w乎D�X�٪C��>m��vm�ݴX�Xi@��@�M��en�xQ�:���N���߷�m9ı,K�~�bX�'�߻�E�,K������K�S���a�]�9�-�fT�å:S��߻��!�����(@�	 J(c0#c(�����Jc9�Q�Z٠ȫ�|FDȖ'�߼ͧ"X�%���ߧ�"X�%����fӑKı=s��5��\�&6��O�Jt�Jt������,K������Kʈ�E2&D�o��r%�bX����[ND�,e:}��}�ٽ�M�&˼���N��������Kı>����r%�bX����m9İ ���[ND�Jt�O�����f�\�g�>,K����fӑ,K� �w��iȖ%�b^���iȖ%�b}��p�{y�^B�|Ͼ�\��
Q�dlq7k��D܆ݛ7�-���c-�E�C;t�wF�<�.���fV��y��ҝ)ҝ/���m9ı,K߻�m9ı,O�����&D�,O߿o��r%�gJt�����卹Խ�WΟ��N,K����r%�bX�w��6��bX�'{��m9ı,K�~��I���N�����6K���Ο"X�%��߿NND�,K���6��c �wda5:ec	�0�}L�� ��^@�g���;Y;~%o���It�!cF��oz���a���vE$�"Ǟ2� ��InG o�I��d52]z."����s�a��4��Ⱦ��Ғ����<�����p���4�K�m!��O�ᯯ�:	Mx���9��~���+
E��A�;]��	aP��l֖ Fc�aBHB�cq�n��&<˚�|oW7D��y�qs � 4�b�zJJL����u��燆��i�׭�͚�a�>1��1X�}R!���8�D1]?�4�
z��S�������(��~@Mz�
��z���m����Ģ��v��A�X���{��"X�%�~�{��"X�%���7#�;.�Mj�Z�6��bX����}�ND�,K����ӑ,KĽ�{��"X�%��~���Kı;�Կ:d5��Mֵ6��bX�%�ﻭ�"X�%�y��siȖ%�by߻8m9ı,O��ݻND�,K��{o-/�.e��=;������`W��F�n�ι�\h�I��~wC�'�_8[�0�_:��%�b{��~ͧ"X�%��~���Kı>�_v�?)șı/{���O�Jt�Jt���zYg��͐��ND�,K����iȖ%�b}����r%�bX���m9ı,O3��m9Kı<}5�;-2�R�-�Z��r%�bX�}��v��bX�%���[ND��\��=�߿fӑ,KĿ~�魧"X�%��t|v\�34jf��%ֵv��bX�%���[ND�,K��{�ND�,K�߻5��K���E� b�B��D�y�]�"X�%����q�&�1��/���B�������'"X�%����vkiȖ%�b}����r%�bX���m9ı,O����0fi���6�\�Kn�Lrt�l�+x��KE�)X@���i��:wI�s��XXۘh��kY��%�bX��߿�r%�bX�g�w6��bX�%���[yı,O3��m9ı,O>���Yp�֩e��r%�bX�g�w6��bX�%���[ND�,K��{�ND�,K����ӐBı,O�����k�[j�]�'�����/!����ND�,K��{�ND�Rı/��Mm9ı,O�ﻛND�,KקK}�u���å:S��8���~��6��bX�%���ƶ��bX�'���ͧ"X�%�}���iȖ%�gO�{��k����t�t�Jt�ϻ�[ND�,K�>����Kı/�}�m9ı,O3��m9ı,O}C�zAO��� ���uU�X6Y�Q��Y�pS �mn�� <c��$�ޜ�2�hT0�m3��Q�5*�f�k"�nY;P�`�Dq1�g+��o�����Ԭ�V6���6�W���L�v�Q�Q�j��9�c�@��u�H�N��2n<�%# �м��k�l�0�#:)i��n6	�ËF�6H�s���s��xh��3D�#qYa�K(�]ic"�ll2��7��O�������Xr�a���2Ҕ�1F�4+�;Aή�^<i��ziٔ(���}�ݾ��Xk3F��ı,K���siȖ%�b_~���r%�bX�g{��r%�bX����|���������;>���X%��k6��bX�%�ﻭ�"%�by��siȖ%�b_>��[ND�,K����Ӑı>���eִk35�.j���ӑ,K��;��ӑ,Kľ}�f���c�U�dL���fӑ,KĿw����Kı>>��ֳ%��m9]�'�����/!���_9=�bX�'{���9ı,K���bX%��뽻ND�,K��܎gu�L)5�Yu���"X�%���}�ND�,K��{��"X�%��뽻ND�,K��zkiȖ%�bw�� }��%/-��J$6z�n��P�2��β�%&�D��jBl��fQ5%�96��bX�%���[ND�,K��{v��bX�%����Ǒ,K��{�ͧ"X�%��ӥ�3��k3I�k4m9ı,N�]��r5���$A��H�=_��3�=Q,K�����r%�bX�{�}�ND�,K߻�ND�,K�'�i;��ֳ5$��[ND�,K��zkiȖ%�b}��iȖbX���xm9ı,O���iȖ%�bz�k�^�&�.kE��[ND�,�@,O���7�O~��6$�H����M�$^ľ}�f�χJt�Jt��Ͼ�`�1V��x��bX�'�}�ND�,K����r%�bX�Ͼ��ӑ,K������t�Jt�O�O���7��[�ak3j��V��P�X�D�@�K1���o+5��R�&����M���5r݇M�u��t�:S�:S�����ND�,K��ݚ�r%�bX�w��9ı,O~��6��bX�t��Ͼ�Ņm�F\����ҝ)Ҝ_>��[ND�,K���6��bX�'�}�ND�,K����rbX�r~���8m� �RZ����/!y����m9ı,O~��6��c���)��H R	�|�F���&D�k�ͧ"X�%�|����r2�)ҝ=��w�u%�ʞt�%�bX���xm9ı,N�w6��bX�%��5��K�K���ͧ"X�%��ӥ���s5���֮�m9ı,N�w6��bX�(_>�Mm9ı,N���6��bX�%�ﻯ:|:S�:S������#�3M]-�n�a	��Q�L��[o9*�����,�g�
�c�.��t�t�Jt�K��禮��bX�'}�}�ND�,K�������Gșı?g���ND�,Jt��c���	p��-�|���N��bw߷ٴ�,Kľ��u��Kı;����r%�bX�ϻ�[ND�)ҝ?����&�GJ��O:|:S�ľ��u��Kı>���r%�bX�ϻ�[ND�,K���ͧ'Jt�Jt��=�{��t�$L��>D�,��L������Kı/����ӑ,K���o�iȖ%��`>xC|����[ND�,K���b�BmM����^B������ӑ,K�>����r%�bX���m9ı,O���v��bX�%��n�M-�N h�$ܲ��F��v�n�wX[j䇹l��f����LE��
U.h�ӑ,K���o�iȖ%�b_��u��Kı>���~T�DȖ%�~���"X�%���R���ʆ�ՙ[�'�����/!����'��"dK����iȖ%�b_�~�kiȖ%�b}߷ٴ�O�3"dK��?[������_:|:S�:S�����iȖ%�b_{ޚ�r%�bX�w��m9ı,K���bX�'���{����+|���N��ӡ�DϿ~�kiȖ%�bw�w�m9ı,K���bX�����iå:S�:O�/�~�F�r�s:r%�bX�w��m9ı,?����m<�bX�'s�fӑ,Kľ��5��Kı<j��pH��.��I̈́���חfgu�kZ̑��4�Ժ��9���wjGV�LK-3�E��o
�NO6�sla���X�vF9��\�8��v{yZgQ�^�Kd�幜����ҥ���v{]a:��f�t2����EM�{���N������I��vǳ�<�-���9ݸ����:�\v��.M�k9az����|6ʡ�5�\���%�[f��X¨:���:�	�K�9��4'{$���՛f�0��B��b`�!vj�X,(���݅�&�W��x9�k��1�c16����t�t�Jt�/���[ND�,K���ͧ"X�%�}�zkiȖ%�b}߷ٴ�K�����ϔ��t�!+�'����K���ͧ ؖ%�}��5��Kı>����r%�bX�߻�m9ķ����^���i�0�]�'����K��zkiȖ%�b}߷ٴ�Kı/�w��r%�bX�g~�m9�/!y?�>�]� �!L��Oo!Rı>����r%�bX�߻�m9ı,O~�{v��bX�VdL����O�Jt�Jt��ۿvn���3*x��bX�%���[ND�,Kߵ�ݧ"X�%�}��5��Kı=����å:S�:����fjgM��3��^�չs�2�q�r��v"�nT\g��!�hg���|����������ӑ,Kľ�ޚ�r%�bX����l?
�<��,K��ߵ��K�S����~�c��U�t�t�Jqb_~�Mm9D��@i '�+�D�,M���m9ı,K�{�m9ı,O~�{v��bX�'����~�DZe������/!y����iȖ%�b_~�u��K���>�~�ND�,K��ߍm9ı)���{�65�&Ҳ͔�å:S�L��w��m9ı,O��߮ӑ,Kľ�ޚ�r%�`~fD����m9�)ҝ=�?O?-2�ٶ%WΟ�%�b{��۴�Kİ��G>��ƶ�D�,K�����Kı/�w��>)ҝ)����<��K.t��X���V��n�X����c8;�[3�m����	w��j�0���'�����/!��魧"X�%����nӑ,Kľ���iȖ%�b{��۴�Kı<���gm�Y���4kiȖ%�b{�w���Bı,K���bX�'�k��ND�,K��zkiȅ�b[�޴龍n1���Wy���/!y�߻�m9ı,O��{v��c��$E"�!�D 0"�	b��?'�l�9��?�r%�bX����ͧ"X�%��Ӷ����f���k[ND�,�"w����9ı,K�~5��Kı=�����Kı/�}�m9ħJt��������.�E[�O�Jt�,K��魧"X�%��{��r%�bX�߾�bX�'�k��ND�Jt�Ow�寧ȍ�
j\�0�Gmn#9y�e���6���u�m��l�m�ws4�@"-2��|������������Kı/�}�m9ı,O��{v��2%�b_{��"X�%���O߱�Fmv�%�]�O�Jt�Jt��}�m9�2&D�;�~�v��bX�%����r%�bX��{��r'���t�O~����E��m�r���҉bX��~�ND�,K��zkiȖ?��"}��~ͧ"X�%�~�kiȖ%�b|}��N�-���4Y.j�9İ@lK��魧"X�%��w�ͧ"X�%�}���iȖ%��5Ш�X�1MHDg���&��D�w�.ӑ,K��۶نw32�3T��m9ı,Os��m9ı,?	C>�ki�Kı;�~�v��bX�%����ӑ,Kľ{��V�qv�R`J��.��΄�%4����2�,3
�pm�<v\#u��F���Kı/�}�m9ı,O��{v��bX�%�����ND�,K��{�ND�,Kקm�%�e�f���ֶ��bX�'�k��NC�,Pșľ���[ND�,K����m9ı,K��w[ND��2%��ڿ��~պ5��d��Z�ND�,K��ߍm9ı,Os��m9�lK����ӑ,K���w�iȖ%�bzzj^��-��-�|���N��!&:}~����Kı/���m9ı,O��{v��bX�%����ӑ,K��;ܷ ۱�u�U�r{y�^B��ߟ99ı,O~�{v��bX�%����ӑ,K��>�siȖ%�bt'̃�<�uO�A�� 3]�8d���yB0�!$�'��Z��0��������I�,����w��X�C7��07}n���ߢ�bR3�>5�|l6�'�h6q�Pjk���n�܄��|�}�Dd��!��iQ>pO��=��x�c$&�c_�P����}~�xkZ֭�ִ      �  	 ��[UUG&Hم��z��J���\s�<��&jVL�ڧ�֍��٬�I{N�l  �Ʊ��]��-ue���a[� ( �2�p�rm�p�%����2���p@�a-���%�ѩ��ʜ��C�!�ӛd�7	�9�@�]V�պ�$�'\��n�n.��6�Ͷ�u*���=�
�;a���&VE��Ê�p'j��!�]�2^����Mi�ۆ��ӯAq���bֶ�Hqk����D�kʈl�;�<`�P���ȭ�i덞&�X3���kV�+�^\��:@�6�CT�Q§g���X9��ƲrJ�ݶy@$�#�vh�7U��v�e���D*y ���cr�l���M͡m�s$q,��[/T�����3��:�N&���m��n�*�J��Ȼ��˳��E6���B<R�@�T�Pj2bVkTь(��0����\����	�,n
<�sۂ�J��Q���.��!>mQ�R�R��45�6�ok�vn��H� M��ݧI���6�[wH�g�2���-[�l��^��;�'�n�p�n[�a���F,�5����c(�@f�gtr���x1��,qJ�Wg�Vб��ηRF�<(�w[��M��.���n�=�l�Ss�[���$��8��]Z�	�f�8���l�)BT��14�%̤6�s6۴Gě2��*�U�5��QNh�*چ籝[mu��F�
PΜ���K@T�f��Jz J��laB�7hi�v�@`��d75�m6�Ґ��k��M���؜s�g\�F�oN:�L2\��X⧗�x&����m���n�S�F4l��U�vh �w@�n�[n'^�m��I�1+mZ���R/-��@0�[�T�\��T��]�[h9�^�d�B��%Ɓh��-��z݌�� D�(
�+)e��t�l6��u�L�A2gZ�X��:N�d�Ҩ����<M�h B(��ୈ���jp>��J�-#�
�
}=�S���l��Zֵ5��n:l!A���sA�
�<mۛ��k&��ܦ�
j��� Wu#��>!k����ez.�
�3���f4�b���*� � -�����ݶ�u� .����q�h�4��-���;�.�Dv(7x���J/T93���xŴN��B��]�a��3e���J699U��V�M�n|��sx��a�bSAOVl`\�nfY�����t�:M�|ی5ɮ�"w"v��r�b0�gpf"Zh�ev�f��)��2��$g�(�M��_9?�!xX�'�k��ND�,K��zkiȖ%�b{�w����șı/���o���^B�������	�ai�iȖ%�b_>�Mm9ı,Os��6��bX�%�ﻭ�"X�%����nӑ?TȖ'�?n�g��3&L�,��[ND�,K���ٴ�Kı/�}�m9ı,O~�{v��bX�!�߾����B�����N�覦��9��m9İlK��w[ND�,Kߵ�ݧ"X�%�|��5��K�,Os��6��bX�'�N�ӆ��ˢ�I5��m9ı,O~�{v��bX��9�~5��%�bX�g~ͧ"X�%�}���iȖ%�bw;��ˆ��lv.̉��N����a�9f��İBh���
 �y9+��1�-��q�y��Kķϻ�[�{�w�rI�����rɚ��`ee1y��*��NJIʖq��{E�4���5����w;۹!�nԿԑ�u�4�(��2�9"����;�uY��UĎ�R��~�3��6E�#��j����T�g����T�;�uX~�s��n�XZ�!x��Q&�R��v���r��g�� ��K��U�����9Qȩ&��.I�[o ��{+\�����av�ش�e�[h���!9R��=�`��`w����s�r����~�R������q1���e7"��l�ܮUr�3_����T�;�u_�H�z����Rq�H�F�3��n䜾���
#B	4�Īx/��K�|Ϲw$�y��ܓ�2���Q�Q�ع���?s�'�~�`o����;����8�g����/?!%Q9IȄ�;��U����n�|k����n�[}�ӽ�a��ţ.X�(��q���`��N�F�K4@�0�]H<\6ۨ�T��;����=�`}�v�����+r�S���tۉT���=���r��<�~�`o����;����c1%�M #*R�>ǻJ��=�g�U~�Sf�ߥ���+�[H�
t��+���,��+ ��K���>�=N�U4�m��`�h��1a�; hD��z,A?~�~~.���ϳ�uX�i�R�X{�,��Vz�iXǺ��U�Uwu+�	�����m�{=���b��3y��s/���[�4 ���9��M'R�'��RO��~�;׻J��=�`��`gZ���nF>G"�>ǻJ�\�+���V���q���bרIQ��I9J��=�`��`w�>ǻJ��ҵj)CITe*rEaꤳw���~�>ǻJ��=�`gkjlj@r:mĪ	�`w�=����|k���w3e���ns�����UZ���6`�Mx�ʹ�$L�:"����u��q�.'�ms�6xκN��q(�sjq�<����(�\����"�\-,&u�-Y���eJp�Z����j�=C#7#��Vuؠ:��1و��kx���#�Gj�1�K�Z�H�w.Z�l��@]��S�M�ɭq�����8��f�+<y�v���m��u�&Ð�V��w���$��4/�`θ������n�+zԘ���(S�Vy�=X��@9�j�2c!�J��H��y�Vq� �f���U�ܭ��-cT�ܥ`w�r�ʤ�7},��+�{���\�7X�~�M4JCR+ ��K��U�s�bݥ �=�`w�eJhc�`6���`n=�Vq� �f�:��ި� ܌N�qXcݥ`w���`w��,�
��cht�ݴ��qۄ�m��/hR����q4���H��&qυ@�(�8�NR�;�uXfl�;�u{�\�����~�`~ZW��'JP�U2�kWrI����*,Q�*��=Ϸw$�����I����O�&ǿg��L��ͳlm����~����Vu� �͖k�'���5��IsWr~������]�>���]�����{�����zRM�8���J���`{����O��~�>׻J����?��|�� �����
�ӆ5ڸ�N^��]L��s�U5�h��HL�%�96�h���_ n論��U����_��_ �?yX�W��]G#�0rX�u_�RG|��Vy���37e�����cߺ�����M�#��oߥ�ϳ���><����B���I�c@�!���g{��;���'�j*�Tr$��a��UŞ���zX�u�~�Y��R�5a^�IҔ4�FR�$V��,��W5����vu�����JI��NNAS��ַ�ؚ�WM[�>��o����D��e�$�ui�)%6�U�|����ջ����_�ʯ����2���~�4���J�q�wv��s�I��+ �����w]��t�c����.�Kn���]�������37e��w]�wwjX�Flm4�)H�=ķ}�`j�����ZܐT�?F�j� ��/n�t�����?��k�.���VI`b��`~�9���{���ߟ���37e��͵��J'Ơ�t�)"�����D����X�����Tc�gl�xQ#�5$br7�wwjX�uXf��>A���;YƵyH�TrRNT�3^���`b��`�ڗ��U\�\lե~�7M�J�)S�+ ��~�-�v�ݩ`f��`gka�RP��ۉTJIa�����?~��~�R��{���s��%��K)hj��ЅnR��v�ݩ`{�����_�ˠ����Ż��=���i"�Z	{���U4($&Q)�i���a�7�����5c�XRֶXd#�u]d��m�P��d�v��(�������c������&u��dZ�ĉ�{T9�Ms��g��@D�l��"�iă��7�5�V)�.��y�\b�c/�,���]ĭj	��[UXc�q�4��psˉTٜn�df^�/u�aT;CCA���]`i�ң���r����k�����s��/%݅�= D��3q�)d.��ok�u��6M=�f��^vԙг]-�cQ&��}���ڬ3vX�u��W���R���*o�Ci��P)��fn�� ��԰3^�W2�G���)�7$�5{�v�ݩ`f��`���ε�[��I$��m�`�ږk�V��,=K_��`v��j���TrRNT�3^���`b��`}׺� ���ߦ��0%�#����k�O<�j�sm����\�E���r�v����쮐J�)S�/�7}�`b��`}׻���U�����Ȓ�Sn%Q)%����ٿ<�����IL(P���7!��!�iBB���h�s��'����I=�ﵿ�T���7�I(��M�T����zz+5�?W7}�`j������gM1D�9"�3^���`b��a�t�������zٷ��k��MdV��,��*�������V�ޞ[~��''���s5��Xe`8��[�&v�l=���M�$(�ZB�Ŷ�]ӣ4-]��Pr�ȓrN��~���wf�`n�������K���� ) ��ۍ����b�ܪH����7ޖ��v��bרJ�G*9#nE`n=�rI�}�π�B� q �2Il!�|����Z�����ᥞ�K�F�k	��(aKhjE�#	p�0.3-����ν���Hq�ۡqwM����\-��
4%�UYA����� �d%�$��!�U���fq6�	Z�G%	BQ�!Ձ(��"�F*�cX�"��H� ]�3��F1; �ǁ/�>�����H�I��hi���f0���P&f[�L���R���%�VD�h�Fc]0sO�l�]���.��� �!��<(Wa��.s34e�K����4K���a�h��1Vb B�S3%�\�AD�3�kn������(��0Q]/�P���*��)���Uv�����!A���t�]{��̛���V�M��4�F&I��}�`{_����b�7�3���E Ԓ�q*��X�uX��m�/���yXsvX�*�A�J"�Pkj��>�l�v��ە�&kRKBFЙ�Cf����nBQI!�R�8����X�uXsvX�uXei(�$�b��rE`n=��U\H3}�`{_����b�7*i�m��P�V�ݖ��V�ɱX�uX��c�M�)�'$�7�>�M���{���<Sap�$�@�`��FI�l�'�k�nI���k$IH�������6+q� �n�q�ܪ�==�
#�X㌘Hc'k��6�.�a䭘���vx����A�9i��3Ox����+�[������svX�uXw&�`b���d�M%Q�ԑXsv_���~�;�=���U�����'(rJ�Ī
I`n=�`}ܛ�����V��K���i�$�jR�8�?s�]ͿE`{_����,=Uʪ�UO����`g��(�RI�(�$V��V�qf���=��W$���]�>�`E*$B� �w�:y��&ʪ��9,r]��+�k�� 05���L�U���d��G���\��,�Ȑl$�L�
�Z���f�i�#��Z�j�l�����؂1�.�qd�*�l8sm$�HŰ��vP9�Q2nv��g��L�����V��x���;��3M�u�"ޣ�fw�mӊ�G	�q���n���36Q��fCPM`#�(R[�ٶp����=��nNIo��Zf�p��A�=�:MR/fw@�E�d �k).z�i-SK?t�ٮ�6�i��)��zX�uXw&����9�����������9��D��X�uXw&�`n=�`��~���g�k��$Q��䡸7����+q�?r�Č�zX��+��3^���Uv�|d�������������V�ɱX��hr�i*�'#��;������_�_�.����+V���O�q94�+����ۈ�c;!�<��/jش��J�^&^�Y��p��rH�AI,ך���c�5nk�_ 3}�`m/Q�o�đ)P�V�y�7@؅����Z�d���F�P�$!_��52m�����(�
�Z�$�F3 P�FHe�AI$�ۆ@_Q䜜�o��$���[�}�5Xv��$��&1D�I#�5nk����I{�|���G`w^:i�m4�R�I�ꤳ���<��v��c���/?o�������Lr�Ȓ�KV��r��پ��<��v�ݞ[};��4�qk��\зk���!�˲[�;0����Mk���N
 ��y��D6�J�8��f�`j��`��`j��`v����Ѓ�$�M�,[����,]�vVf�`ut�6JT�UNG�wse����Ü�r��+$@ �(
��_}�Zܓ뙮������G%I"U	$�5wu�Y�%��3]���{},��4m�8�#%*M�`ufl��ʯ=�?�3��`j��=�6��)*9$��U.�B�cy�nQ����^֫��(�i7i�cA6Ti1�&H���<�|���,]�vVf�`f�t��bi4�P�; ���Ww]�ՙ�X�5ߪ�Č�Pח��c��D�rXY�;�3d�5fk��l�7լ���NJ#����͒�ՙ��;���j��/BM�	-!l����`\�V�e$��15q
K[�`�J��}W��{�����:xd�2�z��I!rKVf� ���Ww]�ՙ�X���+�+|����6.����)���8$�\f5�����L�fPp���BR����r8� �o���������=U�-�;r���GRJNF�I`j��:�6KVf� ���ڪ�+���R�4����b�����grX]�v{ZJ)�i�Q2E$���v�͖���3d�1uV����i��RR+ �����3d�3^�r����
��$�,�^�4��в^��?�������7�$$Y�Q�nz��3��q��Yl՗4�F,U�鍽P�=�����ғ���0�b���lT�����Q��t6�Ѷ�7BЛX풹5��+2X���Dg��KM�
��^��b�'kd8֩����KZk`�;.��)hBN�6,N� [/�����:�:h��]h*X�3�^9t�6�CUn�X��`��G:��9����6RT����l<��e�V��ݩBm$�j��D.���̼�E�2$�� ջ�����,׺���,�X��R9(�6�:�6K5� �����9�$em3ͪ<�9RHDܒ��?yXw6Y�UW)-[�;)n����j�a0�r���9'9�����oN����,�vu��Okc�1I)9�I%��7]��Y����v�n���J}m�h���B�h�B	q��V�S%��c4G[i�4ҫ.���R�	�`v�f��3]�}�����;��P�66��%E#�:�߳~!� $L��q���5�'���`v�f����{&�M��#��6Xc�Vz����K=�`b��>���Ckx)HdI�%�����Vig����v���\U#QD�87��.��3]�w����zym�Np����,j�X!���mpL&�	sD��k�cQ#t9�n.m+'e�l��V��ԩ%&��[�v����{����w]���F��ԥM%Q�F��6Xc�VԻ����vv��q�II��D����U�����8ެ�)hA#��	�]BL��9 �Rm�BF�&��O\j�.����$�~����kh �(�J�"���[�7��Ż�`nl�3�uXmlT'�M�M(�J�+�s]��W?r��~���=���`gi���@	l\T@�ۨ�[Nų�	�������h�T�9�B�!����Q&� SN+ �se��{�����^�Us��V�hkQI���C�I,��W�#r��X�V����r�Ď�Z��n(��GQ���{�`unk��9UI��X��V{C�M0�F�D��Ȭ��v���:�V��xiD1����Ъ����+ʰ<�Jt�UDn; �se��{�����VV�se=p7	�n���QG�<AգD6ۀ��f�ߚ��~˜c�׬�%j�liy��Hn?yX�y��������}�����^e:�0���8��<�`unk��6X׺���z*�mQ0�V/o��}�����%���`nS�+0x�EJi4����U%�o�����`gi�r��?o����7����C�I,��Vv��:�77$�}��ܓD��r
D��`&��h�=�'������>�Ҧ�޾�ɚ��x���"/8fqi�T}�Awx˅�	sW5��oE)u���%W	���JBU�CÚ�5����ȐcA�E�bE�Ă�8�ۚ���2�VE�H��i��~�k{�.�� �!������7��d��sD��FA�n��mz�i��M���df�6x��x��')��	nK��s~�9)/Zx'�"
��8�!�=�u8y�WI�-�h�߰ѭ��{4s=� ��$߆�Xl�#�-%��
�h��K�8k|e���ow[߆F�$8��!M����>+=�T�	>2�fa����֧0�Z֛l      2Ѵ� 9�-�ٵ�ٺ�Y��.�s�;��g(W;1�
8- ��y�P�yl�nKCE�֦���"/�z�iY �� ���Bl�� !`g��r�M�j�ms�n��3�R6�8�����q��]S4F�+�H�8$.��7[
�J\�C,��� fj�[u�0�v�]�àM˳Zk���*�5��F�M�Zv�x���4����!.)��â�#j�b*7W�Gm�� �պ��G�3�]��՗�x�9�5k#��MQa��k-�msؤ;+���#��ښ)�8��6wm�%�����)�T�F�q�曵局3]L@�b�[K��@mgvn �%���v6˲g�ꃩp��x�Os) ��M�\	4�9�CW]/T�=�F�d�J�HT�nE@IW<Ә�ڒ�k ����4]�YP+ڎ�:Y3��ᢀ�/iVBiV�*�K��"\��\��*�M&]�@�Cge�a{���p�6	�Y�Vɪͤn.������JK*��llY���c,��a���]�n�v�.� �t=��:as�Uof�ٺ��6˚�&��eѧ��K\�G����Sm�u�b����dTؙ���]uR���Ø��G�vGMaJ΄�D�(�˹WC�B��[v��[�n
��h��2���aMT�ƽ!�9Ĝ=�K[��Rp�Ȇ�cl�ٻ�$- p�ֆ[�UiVs�iT�*�Ε��^U�VK���&.*a��P��z��F=It���V鱻mٶ$`�v�J�E�eZ�1�[=�s����C!����.Dὰh1r7I� �+\\��I��p�:��4�#�zؐ����u�[��D�0P�.t/5��U3��p����5p�� ��Cg�-�lI�R�Q��R\��]�eZB.���h�A�#p��ñ��!�
�wF�C��
��Th j�hv��50F�f�[vQ�A���T�Ӥ�7u��w"S��� Ӱ�&���͠����(h҆@��I��F�xD>pOA���~T����jd.�cJ�׳<Hb�r=G,br3e���n��1�̣���ᔶ� �e�nx����8mvؕe0�;7e�֞;\f�U�6J�s�Nv�8�l�%-�579zi��(4.��4;�d���v��E�YˎZD2�׬{//Rn�N
ݽB�B�mtom"�](�B��y+92�0����ϭ5�F��V��e�6*��GM�s�'$����sVM�D�؎��\�'Y5�������w7MQ����Y�LaȀ�++��ym��n����w�� ���|�q���̡�b~&�"bt�VV� ���:�U�����](�[D�M%Q�F��l�3�uY��[�������`w2lt�D�Sr1TjIa�=�`n?/;�s]��q-��XK+R�Q����H��ծ����s�����X׺�rt�}��b�R/hЮ[ɥ��9��z_7<����6"�:78�d��wy=F|*�(�Ԓ7�5~��`���ν���UU_ �~�v����JI��73rI��}������f��g��ǻ�չ��UURG�hh����D�X��V��c�:�5�n�>�X��	H��F�1n�;�s]�f��Ur������Mh��*I�E�����v�qo�����V-ݧ`{���J�F)J��Z3mՋ3�F:�Ft��{�%9`�/6�N�w�y�����Gg�=����׺�[�O�s��W�1{|�͞��ێJnF*�I,��V,ݧ`unk���ܪ�$m,�I��EjU���_��7$���ٹ���0 �Y:j�B&Z�Q�@"	�
��M��d���[�}�{�ܓ�͈O��7LqS���a���X��v�����{���W9ů}�v�Z�z%���(n; ���:�U�wsI`unk�>�ǬrR�u��	�8c95Nvl��Wn#F�k�� ��m�C�;�4"/����5$���+ ����������,�Z����9(��qXw4��s�I��v��K:�U��W3)�)��H�@�BX��v��,�ķ��=�%���F��)��4��v��,��V߽�krz��(1K�}���ܓ�}=pn))��5$�3�uXw4�V� �ݖf���'9ĝ�4\@��_�}��^~{;�mĖ&L	!Iv�[�i�7[Q7*TmĢ� N/�3��X[��3v~�9���+��瓤�8���%���U�s��,����wsI~���g�ם/�(Ll�"�{��`w^��*����,��+��Ax���A�%��{��;���3���Kwޖ�zy�	I$rQ%F��i,ܭ��/�7}�`w^�&��	t!Z�@��v�~3;�U.�ֱ�p���N�ζX%,�*�e�4�G�i�]n��E�P4�ж1A�6���D�T��-�lv�ͥ���d���6�2���9�]��{(��7�>[S�3�ja�p��u�V�
q�3M]��2���B�ǁxؗ�]lڻDݩn�B �2֛]�M�(�H(s[�k��/b
+�5��S��k�u�'��sg�#r�n��l���y��j�v�9�2a4΄�u����U�e�d��7M0�B�����i���l��q�h܏�~�Xf�;�ur��{|K� ���jSITi5$V��,��V��%���U�s�ʪH���i�9N��Q�%��~��i,�\KW���7}�`e-���q(�����;���1nk���a�qo��X�=)'��&��Ӑ�-�v��,ך���K�s���砜i��QԄJ����Ƨ�ۦ7iN� ��0����@��M,6�ґ(Ll�����K5� ���U���<�{�6�P?�����Nɩ5������w�1H���HbB���"�P���#�-�,	������ߦ�$���ٰ�l�7���QFG%�n+ ���Ź���\�Tٿ��X����3҆���m��"p�-�v�͖nM,;�KW@׮)"�Ҩ�r8���,o��|��%��s]�������2��cC�AD�!�v���f6�B��M5_+q4I��ѯi���E���nM,;�K� ���o5���ۉE%	��3���q#W���3��`f����y�	�A�آ�Ӑ�-�v�͖]'��UU'�C���B\1��De!�1�!�zQG�|ϻ��ܒ{�~%���:OQ�1�RGa��,��X�V��%��s]�ݠz����`f��`��X�5�w6X-רL���`�D�T�|y��#�u
�c�ŝ�4���A�&�J�(�R����7���X�5�w6X�5X�iCz�'#i(��%��s]��\�a��o��Xw)�1|�(� �U��; ���5� ���Ź���rjq�$�$B�rX~�W?s�߯ߕ�{}��-�vGM�@��=�[�{d��.gĹsR�%	�`��X�5�w6X�5ym�$�߻�Es�0�W��u&���6����S��PqP�<������}�����b��NBt/�����,ך�s�\���%���S~D��l���w6X�5Xw4��ݗ���� ~����l G%��{�`��X�vXw6X� �TrP�F���Ks|K �{��;�����o���? o�m��J"'	`��`��`n<�`��Xʪ�*=�HI�<flt����u�_%l�ԇ`7^��6-����WV��+e��ͧ���nӪ0���In6mh���	3���U׉I��f.�����n�*4kq��^4k�4Z��y[�Q΍�2������4*��-�D�KV�#(KT��Z�,q�V]rB
�Xrg�Y\���� ���-��7���ق�ÍZ�m�ߛ�υ�fI���3;C�Ֆf"ee�Ś)���src
 TA�m�d�:�J�4"qE*D�UQ�'����7j��i?�������,���u)1�9��`n<�`��X�vXw6_�W9ď �y��Biĩ�BqX����ݖ{�ʯ��6o�~��?~V{͕�J��B����%�owe�wse���U�gsI`f<Tޢ�): �,��,r�����������$������ M�'W9�aR�j��zt��Q���ۭ�+Cl�cm��7j��i,]�v�͖p{��l�$��#qXw4��0�A@*6 
 �X�V��B
�xq�����qt�c��,ǚ��9I���%$N$�"p��{��;���%�{�`��X���G"�(1(�v��r�UW9T����`~���`��X����6㎥&8G#B9,ǚ�3uKWw]�f���W9X��~Cm�[U�eKIH��+u���G&u[סa�M�<�u�T���t��s��B괇%	��{��,]�v��,�����ԥSm!JTڎ)`|���76X]�v������H���7�Te'M5�#���X]�vJ�u�D�||����>XC�� #������o��O�5���s�	<�߳2����]ї!q��s�(�2n	%�/% ,�u\a�����b�<8�>2�S�����!I9y2k�t�T��DI$�6�øhVWZ%�@�$38+����������2{���9��Z�LF����y���W�Cv�ie3VetE��h�eN5�"BD�T��
E�(]�SdFC�Tb%�T�����6h�d�]�a(ar���-���Q~�⡇�p�>�ϑ��&�C���*@��_
|1 ��4@���s��UUUUvv��1wu��A�[�M�#����k���,�w]����o���?y�F�%I%$�R; ��R�μ�`����nk���}XK���vⰬ%Y����ySl�6�=�id���öe�L�˩%dM�μ�`����nk��s������~R�š�5��H�JB�+ �͗�������yK:�U����qԤڊ9��`|�5�f�~�[�|�}�� �1'�)�")�'#���%��)`n=���a��K�x�*�QDd4H��)u }��srO�:ŵM��NR��qK:�U���U~~��Ӡb����37T�;���O_Gn���]���N)�z�F��n�vmcD�+�rS#T�EFRlM���V��,�� ��R�μ�`f�=�o%6�@�K幮�W8�n׽,��+ ����UW*�I��Mʑ�$r�nG�n׽,��U��r�#=�K1�=m	����	*Ia�w'��=�K�y��ŕ�������I#JIG�wwe���̛�����'�g�]�<3"琮I�
[! �)��O��+t��R��G�nF����*Н�� vNq�V�V�8�Sk�7E#��uƮ`��u��ֹau�,��af�lů.�g���x�jΞcY��Y�ò�$�0[lLS"me
�M�et���Fudl�h,�]�����ӟk��=1�Y�4�6�noX��lé(�DiAFK��ٵ�n�Y�s�ڗjԩ���X�u˷w��$��ņ�՗f�$mi	H�!�Ƈ����YW�e���b����1�pe�h�S=p$�F*�r`��+V�;׺��@g��`m*�jO�)�" IV�>ǚ���,��K�k�[T�i�T�)�`}ך���,�]͞,v��`o^�oTT�'M5�qXW9Ig��`w6x�>Y�����5X`�U���a9,��K�u�ן�w�Xٛ,�m��6⤣t�]
нkh�p6	��%Q���뢨���� ^cr��6ڒ:JH�,�ek�>��V�f��U�|���Ł�?6�O�(�k.I��Zܓ�g�]�*��,tf��al�;ݚXw+e�Ձ����H҃���>��`}�4��UI�^�u��wJi�⑊���U~~�}��o���>ך��͖R��{R�R!����V��y��>��`}�4���H4T�|q*z�`�*�.�m�e�r�,��lv�rCX�b�nw&2c@�af/��o�<��{�,�&�����ץ��z��(��M��ӊ��ri~�+�Ď�����`}�5_��H���^��	Q�Xݞ,;��¾���EPʪ�B�ʮD��+������<�nS���ԑ�X{��UR[�^�q������4�3��S�(Ӎ0�T��y���ri`}ܚXw+e������U����J%f؉�\L�Fduinݽ��x���.^mȖ��U)A�Q����q� ��l�;�5Xw59
�HH�b�R��U���ͯKu����ʤ��:�<��Q��9 �V���`����ri`}�uXqa�T�I�:r���9�%���}�Ł���a�U_qПHH���C���d"�X�&����WՁ�x�zEC�؛�5$�>ܚXk�V���`��`�Ǭr�*�3�`R,/�ls��vjpm��
�K�YZ�cwRڛ��(M��h%F�`}�uXw+e�w3e������ty���7	QF���3�[,��,�&�q�3Ti���F�i�R����>ܚY�r��~�ͯK��ֹ��(ے��ri`w^�1w+]��T�o�,=�NB�HF�b�Rq���kͯ?�7}�`}�4�'=��Q���GB�3z3:�hPHL�n�i2m��ֻ���4���tsr��m/Ɇ�e���H!��b9|<���+ݺ���dd�+�W��v��n��l�����r�:-�
��㕺��t<hP㚂jӭ�Ó���X8f �u���Ip˥�������
���2��:Γ)1��۶��lt��nC�[N�����X��-P��L�A�l6�Vc9u�$�&p.�,�y^��G�]�>6��?)�Zu����px^��t]��LM�6�G7!�2��?/~��`f<�`}�4��s� ��i�q��Ӂ9RX�5_���_�?z~,��~V���`w��F�*N�i7R
E`}�4�>׺�;����y���@Л��h%F�`}�uXw+e���U��K���`e`��rQNBSQ���V�1��ɥ����`j�4�I"bdJ:�l�A9Ҳ�A��F�n�y�V7�c�ȋ�ɐ�ʛ�����I`f=�`}�4�;�uz�@nmzX����r&���WrN}���|h� ٹ~�}l���`f=��\H3���H��D�AMHX��+ ��l�;�uXnM,�x�GQ��9 �VKsk���{�`}�4��Wv{�����M���iʒ��٥������{��3�[,UUUR����q��H��"\�]q��u
oU�v�+&7SU��Q .:�54�Q�D�!�6&�!�|�o����U�gr�v�A��}�i6�y6�rX�߻Y,͚Xۛ/�*���ާ 2��' ����O��_Mϕ>jB�J�W*�����c���>ݚX�]4�7��N4�)RX�4��6X�4���N���ݷ�}�� ��e�휵�1eR���u� ��l�7vi`w�O�ۖe3B�Lf!���eU�NUu�sӃ]�\�>3�^���e6�I�Z��ͨ��`n��`ܭ���,�͖c1�JuN�E`ܭ�ꪤ�o�� ����{��UURGx����m��GCNT���ŀ}����{��3�[,�z�[ lN�ʉ��T�}�����`ܭ�W_���Õ������C滽�nI�$�:\�^�t��`n��`fV�wf��f��ŨL��q ��BRY]�������1ۉ*�����덐+�'��:ndFF(�qXٕ���٥�}����W������x�B��"6�L	*Kwf����ww���������`b��L��D��IHXٛ,׺�������{ޖ�̓�T�)M#���{��3�[,wvXۛ,��(5؜V���`���>��`n��`}_r��}�-������{�8�a�I*�51�n��w�f�1g�5�w�'���I�3�`ܗZ|z���z{�<��\ѾK���5���(�E��!���Ci/�ѭ2��A4f��|w�8K��kЗ���Y�9��3��������˜�S~�Ӹ�.k{�Q,a��~�Џ���.����o�I�O u�~����7�� F���|5�K�hA"y��y�y���1'���z�߇>|���w����V1F2%��{�J3^ku�$f�<��E��H�0�ys[%�Qjt�� ��B�<<��^sz����7�� �!(H��:#�d��>��wZ׀ͤ�̅�5K�%��g���y��=���9�_w���H�Q�A/ލ�xNa�9�o��-��h�l��/�9G��ٿ&���?W�����      .Q�� 9�/Z �aЕ�%���6�;&8�r����ՅcPͷ^L�&���ߒ��6'`�3.`�����.J�Y:������0$
��R�[/�E<�i���g����'.Wj[�i,�e��y��B#������Q�wOF�U�h仵 ő�!��g��sI��<@c˕x�sU��c����Ƃ�F��r�ʵ=�A9vG�ݑ��v��ݢ'lPp�����)&X��ݶta��n�ۃ7��|�o�x{n�yx�P6�ݴ��;�6.��zE Jx۞��2�S0";��ݎ8גP -�[w[eA���c�hX�C�%�N�<g u]�кV�������<d�^ vP�����r6�\�P	�ms�j���dڔ9�
+�i�;���;m�r1B���+*�+$��Z]K��m���J��h�Z� b��Z�UV�d�m��P77 Ϛ]�B�`�w(�J���f� 
l恲�la�2�f�i�)%�UUy&V�S4Oh6��iپ�خ� 헬;��3�� ZUvWn���^������*���7*Mn%�Y��b�bB0��F�v)n%Y�np
�˻	]R95�:��m��v%��nj��k6{��NϱZ|���I���p�鍷;#�p-�<�]��㇙�kq��]���7����˕��mG 
�031E�!@����Z�N�g�m�1KpJ�E���;��8��:���]Y�a�pW[��L�kL��.�7�Q�)���c=�����<���6����Ie���VT�,�������� �����TYrv4���4�ܝvd�&��6����W�e$.�e�WBۧӺ��
D4������u��c+� r�^<��ke.�J�9F�Z��"V������D�X�S�N5���ɽ[�.d�0���ksy�p��$�4��*�P��\�@)6�ɀ �uc
�۬�g(1Z.j2��Yӻ�=T�����"� : ?�R*`!�=A_ O�����&��iA4��|
����rI��;�����nܨW4�8�.C%�p�7hCs��l�6��t/)z;t�oKSpp��G��g`+�	�Qy���^l���nN�+K�2��H�u8�$�*�-�-ڵ,��8����+0K��W��9ȴ�P/u�_H�wm+4⧬$�s�Cfkv0��X�gg4�Ss0�4�je)�*��m��0��1�$�Yf2��^G&P��b�F���I$d��k��īs�fT�`�-��|�i����ݮ��%R��ZM�m�31M��A�*L ��e�}����{��>̭�z3AmJI�l�&��6X�uXٕ��7we�� ln���h G%���U�}�[,�UI��,���գݧ ���4(�qXٕ��7we�}������=�`n�ɤ��%q��%�n�� �3e���U�}�[,�KvJ8�RR�)�q�Wj��Qŵ��	�x�l���Z�N���ٗ��ãqȢPb�rXٛ,׺����`���;����5�&��rN}����P�HĀw�n	�=t����ޤ�_�5�$����rI�se��9I�D	�)��'"p��ץ�ff� �3e��������bM8�jT��W?7�{����K�٥��K���`w�</H��N��A7%�}����vi`ܭ���,�I	#Pގ��
�1�(M�mV�������ag��Ӹ���#L�	�X�d�����#���vi`fV�3&��9����k����8&�M
$�V�el�Ur��H��x���X�5_���RF��b?TQ'`IRX���}�[��D#�D�pE���ww$�}�zX�6�֣�D�Pt���任�`{�|����`n���;�����QH�h!���V����z|��ŀ}����f�bM�D
�9%8#��Z��0�n���̺3�GWZH������ABN�lR/�;�^��M,�͖��V�U���&�pԒ��ɥ�}����y��>��`}ј�����'L�� �3e���U��U$no�������@6�{Ʃ�#���y��3����ɥ�
��"�Q(՘� p�s[y���t{��$��I�D���3����*�� w��`n��`b͒�u�OP�&'��P�8�ou'�^3ؠ�n{x��'e�۝463�)3�Z��m�:Xۛ,ܚX�5��6�֔�ĜQ!' �͗���q#������y��4��H;�~��R(�I4�Kq�����UIw��V��K�� �'�I�����չ���^���`f<�`}�Y�HBi��q�k�V�s���O��{�`j��`oܮs�p�_)*���I����
���@Q̸0��MlG��<a<�Jyk20�k"�n�3X����h��t2�l���ӳN�T�դ�9z�&�Ҷ.l[�'�,�'����u��4&�]��V�+\m��p�b��,�I*$Y��\��l��������:��P9�-�,�5y8p�� !՘pac4�\��1SG��@)�t�.�sZ�gv6��u�)���mV���I��I35��v�:ѶK]�lE7+/;u��"�77P1��F�+���MVgJ�˦�߀?{��ǚ�[����t`ڧ�j�A9,ǚ��9��r�?/�����~V��/�W2�?z��#nH�q�Y�;�{��73e��3]����IS�(Ӎ1(�>׺�w6X�5�{�U������������S�8ґA�r+ �͖.�V��y����]ۆa�sb7R�++a�M�D��Й׻�i�#�u�ˇkF���9A��Y�v��v��U�n���� �'���H�[�틜��ڮU&-sU�n��s]��f�!	��I:`�,�� �͖.�w&�`�F� �R��D܊�7se������j�>ך��j6����@�Ks]��ʮUwf�||���>��`fnڎRn��Bx4��5�F��a=�gmqh|�hh���6�@�k��vW%5��-��ߺ��� �3g�U�Y�v��?AF�i����^j��6X�����WLB{N9#���X����$���ٹ�臙�ib0�A��	�E�ǠA1C�F]�>�>��� �,�7"cN$���μ�`}�5Xk�V�UURכ�`wt��$�pPj��Xk�V��U������fk���H4PqqD	9=&��j���]7�9������گ`���m�gݩ�I*mē��"�>ǚ�]�v�3_�Uϐw�|�V���QB4�2(�V.��s�\H���;�Vu�� ڍ�{Ʃ�$�>[����:�U������`�j8���BtԎ�ܪ��UR�M�7�Y'�Ͼ���#�=@0sS �">��@5��'~�p�,��]e�e�iH���V.�幮���`{?7�Uck��R�p:�d�C$�l�&I�Gf���U\`��T^mȖL4D�r/�՞�>[����Vu� �,�7"m'Q�G`|�5�ך�]�v.��+�����z��Q4I`g��X���]�v����Zem5E4ۀ�Ȭ]�v.� �se��UK�7���k[M��$j!�$NG`j��=K��O��=�ܓ��f��H�P#�T��v%F��d $U*�H�:q4�I�S�)�'��b^fɥy��=�5[9(��v�>�ݵ{ҷAt85ۊ�+�
Bg����
�b��Gj$�n4�����.[�R)@]BH[�.��7���4Μ�x�8r�6�U<�A�vW��s�ZBlJ�XS\�����&��4�s]q;�*l�`�(��s��s��u��y+92�����lW>�`�m���xy<��fWS	+5˫�3���� מ_3y3F�kU��-�OK�<���7g���v�q�a��;a���	Q�R�6�D�}���;�5X���Us���vV�ި�7q��R;��U��������`|�����MoTiƙQH���w]����;�5X]1	�JD��PI�������՞�;�5Xz��,y�v����$jD�@��.���U����`b��nn���^q�<^2�U�����ۚ+�uD����1�CY������ix�A�J�b�>��P���`b�(����-2��*i�uC�X]�w�r�U�(�]��T��2{}��ܓŻ������\��W��oԉ#R�r;V{���wu��5X{�,�j&�aQSh$JG`|���ǚ��͖�W)y����Q��j8��v��V��7��<��v˻��Ŧ�ԅG:�(�AGAU4,���,�J����i	�a��IIc�QKff�t�Cr�iƙ"��6X����w_��A�{�`b�P��n�cqA6����幮��y��3���;�6����H��R; �se���U���xV	��H����
_U9��$B�&�L6I�&?g��o��bx�����|���^�$ќ�]Gʲ�
�_	ZB�>��o�\�6���.�b˄�RS[�033|MK�s	1.�S���������<�ӞiT�3xrpތ<7��n�9�Z������X��%QX�l6bR�i W������4�����>޵ɘp!M�i��]�9�D�0�)� �S������5���6���_M��� 3BnGT�����|��+�Jy����a��BD�kxm��h��ADaȔ�LN�s~6�f|�#�M��C�P��OAQ���> �i�bN5�Oq�|>U�"�A!�4]��S�=<TG�G S��}�{��<]�vۄ��'Fӊ�m!�,=ʥ��`��`j���+�w��`g��5I1�Rt܊�3������`nl���`n�`��c��9"��hX��5A�����k3¬��[ .:�54�K���D��M��rKWw]�}���73g��U_ 77��﨣�MW�QSh$JG`wvXw6X{�,]�w�U$g5�z�n(��16G%�g���;��`b����,��MoiF�i�$�˹�����`uw5�z��E~"#4F�G��!!5� !��&H(US�U�R%������O�7R1��Br+ �we����`�����uX���_���I n�.�ˑ�b�23flR���;F:;��ٱ���
mv�����RP��O�ś�`�����uz�@w���;�J\tz�T�j%#�33n��ʤ�����w���;ך���$o�^j�ct������`n�;ך��۫+Z�oQJFJR�r+Ur��}�K1��u`}׺���6	��TT�I`w�4�33n���n䓟}��$���T�C�$�׳oUt(��%2�h�5���5���6�g�� SF0"�v��4�&Äδ��]X�J+��;�v�;&a�8���?s����E�'��v8A��j���y���SWFi6�b��9^m�����t�q�<�mS�l=��`���Tк�Z��;!&[�m�͏q<ss/M�F^ń]ټ�D�<���]"[�.SE-�msE�V��;����t�{����i+��BjB�M�7��x"�Y�;1ٙ�o\m �9���s3�b �7qX���Ձ�=�`n��U�׾Vc�6z�n4ʒJ�>Ǻ��ݖq���u~�UU$j��O�7R1��Br+ �����<�`wj�>Ǻ���j)*(ԉ(�I`uw5�ǚ���U�}����0���m(�4ԍ�`wj�>Ǻ��ݖWs]�ՙH�'#���JD�@�ݴ��ڸ�Zu�m�[��[m� ��:�Ę�)�nE`}׺��ݖWs]��y���ֲ��Rq�JS"nEd������C�1aѶI$Vb!�)�hjoY�]�=�7U��^j�>�(�&�aQSh 9%���k�;�5Xu� �7e��kմ�r5���R;��U��<�`f��6X��MoiF�i�R+�y��>��`|�5�ǚ�Us����òՙa�\��BP����<W�da����K�Z��I��.)cF���a�|�������`wj�>ǚ���jG*8ԉ(�I`fl�;�5Xc�V�n���R�Ru��Cֵ�'��]�9�{��:ΝQ����PF�4�G�+�0
�q�~�K �{e��Ǖ�P�n��7MȬ�� �7e�}����<�`mcYM�!5�)�7"��vX�^��f��>ǚ�㤕%KPގ��n���$<0M��7.��2��K����lF�V�&�cd��&�je|����������j���,�^�7�q9�5#�>�M,�� �����fk�;ݎ�ޢ6�Lq8Xc�V�se����`}ܚX�e$�F�9	���>�l�>Y����K	H{��T�&E| A=��5X�ݤ�RF�APrK噮��Us����;�|������9�{���F����
!�Ī*�]�hc��.�\�/a�1
F�q�պ�e&�#�����U�}���U|������k�5�4�' nB��j���,��V�ɥ���H�ֶ��!5�D܊�;��`g^j���r��l�`w�|���2�ڃT�Ia�-ɾVsg�幮�>�l�;�{��R��ct9��ri`}�5X���nI�s߮�|BD��!8B�!	YA0�A�A!�`�m�Uv��3��!u�ncs�|��1�(87s[�t�"�C\	PX	J�i�wR�'vˍZF�sۮ�s��v'��KG8{��Q��p-];1d�bv�gD��g��9z��]���� �WghU
�z�ؠ#��Pr�v��XZ6	c��+�V��+�֣h�
T��FM�Bd�Bo��xK<���2K3KsWZ	sV�	A2�4��/N�w��CB�	�y�u�&j�kW0�%��7�Z%18��.���n{r�ͥH6;fy�I6!H�c���>��� �����fk�>�M,]2�{#q����>�l�>Y����K�y��4��NE$i�D$�>Y����K?R]׾V��K�%.=�(�:����4�>ǚ����噮��c�V���' nB��j���,�f������UW}�y�#���#BP�0�h�h�VV���\F�J�´�\�d�fa�[�l������>���`}ܚXc�V�E�mA�m$�>Y���\�ʺ�]Wk�E���D2�����LcB��U\�Wj��l�����|�����׻M�!)���v�ɥ��<�`w6X,�vz�-���M'���<�`w6X,�v�ɥ���ROb�$�c�NE`w6X,�v�ɥ��<�`z�����5)7(i�#bb����	��R��q�a:�~Ƒ�28�[��v��'8��t≠�9'@��~v�ɥ��<�`w6X`a)p)�B�������K�y��>�l�>Y���d�m5I����>ǚ������}�$�	 ������R�������Ʋ��M1I"P�9�}��`|�5�w&���U��QF"�cT�I`|�5�w&���U�}��`~���Q��4�h㋶��u�� ;����h�<8ۆ��Csl͑R�F�0��o����U�}��`|�5��T�B�D�i8�,���A��K�w����4�1t�I�Q�R!9�}��`fl�>�M,�� �sx��t≠�9%��Iww���l�`}�5nM|sI�hHeL*�`(n�ߥ�������Qp`��ɥ��<�`w6Xٛ,W)niMR� �sq�E��s��u�v�u�\z��5V�%w;v��97%rkF��5M�&�ȩ��ݾV�se�}���ϐw6x�=Z=����%9P���}��`fl�>�M,���8���j�LJ�AN; ��K{�K�y�����`w��iH����cR;s��/fߋ�{�`j�k�1w5�kT�Bڑ�F�N)�y����W�o�@3|��f�~PU�� ���U� ��W�*��AU�Ҁ����AE�(0TH*H*D`�AD��
�@B
�A� �E
�A �D
� �A*F
� "�EB
�T�� �@
�����  �Eb�A`�@`�D �D �A`�@ �E �@"�E �D`�D �@ �E`�D`�@ �D"�@��D �D`�AH*X**"�D* �@`�A �@��
�X�V
� *** �DX*b*��*�",H��� �H
��"�������E �E �E* ��@ �ED`�@ �@E *E`�DV
�����@ �B
�
�`�E"�F�*�� B� *"�EF��� �E��D��"�
�X*`* �B"� �D��F
�*��B*�
�`�A`*X*X����
�E`�D
�*��H*� �F�"**��� ��"* �@��F���b*��A
�EH
���D �@
�X
� **� 
������TA�@AU�� ���A^�*�@AU� ���AW�*���(*��AU�@�
��U}Uي
�2�̵��
�"�����9�>�!�4A"� ��% U*�ID�
�P���@IB 	A%H	HT��  (�
@�(�D�*� $�@( PT(
*�H��

���%@
��PT�(Jp       @@  ;�}�]�Ҽ��c�ꮷ��{�מ�fϟs�ŒX��[��Wp �{�U]�>{Q�� R�j�eW&��U��@m��U����j�mNo:ם�^;c� ��}�o��^<��ݼ�ʼ��=�
�   @  Z h���w�|�_o.WKru<ۏwT� Ԫͯf�yq�;��j�[�R�� ʾ��><���  v���W��ԫ� S�T�����x���YD�݊���篬��{�=�&����r��� >�   @���F>�P,z b 0E� 2= SE
S ic4 ��JQ�� "@  z��
P�&��}`t�,Ƃ���(b(F�@8 �3� �ΊR�F����� 5@ ���R � ;��(4��x��NMWNN�`��B���u/0�5�����Җ���ҽ��>�^m/  6�����Ω{� P�қ�{}t�e{�=/6�ە �X�vU޷/l�4�Ͻ��(� �� P p�@���[�>�S��{|����t1�Ӟ��5K=�{i�����}/x ���}*�wɽo-< (@��}�{k��6���>�}��|����w�-ͥWp S:����7m=��y��   ��=��J@  0���H��<z�UDg�  تTR�  EO�	L�*R�  "$!�I
@Ѳ��:_��X��������}>Ͼ���g��ʢ������Ut�

��U¨������S����H�-�b�������(�X�v5$O�M�x��������ɛ��Gq��cA�$���Eg��R�P�Cz4˅�!%bM#!V6�5\�������JC<����3-�8��c�`��������Hۭ5�)�L2و$M�$\�d��=� @��T��$Z���@�wz��;�z����J��^��UX8<(�'�bY
 @1F��	�x����k6���X(e,r��x ��(�Df�2d�>e��37��<�)Q�4�"V�k��5���y�|77	˗f_�i�~�9�,?���4!/�_�����ȯ?�=�솅�4��8%�"� �yC^k^�'h!V01�d� 4@`������Th��;���pk�0�!�Zt�tw�TZg�)�ԁC+HXc	�)�� �!��4b��Q�V5�!�E�aLQ"��5�ъ�Q�b�!���'	B,�����юv���>X�G�� R]�����J̕c�?{ˮN����p��Q���@B$��P!�d 6��	���g<��=D����ٷ�m�~�
9TC��1�<hbr�,,h<-�D�!\�HQ �APP�(ș�!hF��
Z0)�E��&���,�A`����?{+��h��p��eo���N�B@�[�,R.*n�7t���A��T�p�ᦥ0�)LU@�!&)~6��Z��q��b拿;����R�'��1x�6�9��!\g����n��	1���\���#|4wH�(Jx>ܐϑ̜�=J����.]�XJLu$Xbn$�y���XF1c��S����޽�)�i$p�q����O7�H�3\�Í���H倣�kwGh�`�q�؇��{jx"4�0Ѧ�%���dSbO�j
���cq�#XYV$3R搀@S���G��_�s9!@ۼT"傺OY�0k�#k¨ �X_B	C�(D�RA�I`�-�`�,dd������F"$�c���&�߰��1�*B��P�4�6�ݚ.�o<6[���CZcB$��"%t@�X�4B��І%�  �H5�����@���ㆶr�fL�S����F��x(�qd���@�@%�TD*'���ۤ�=�^v�(g��Z���T�W�D�A�^>�cJa^Y�F���cTE/qg��� Y{��$\c-i�\aef)eQiy�{+���L�G]�+(�@�K�,5����5�Jj��xE����,^���tm� ъ(Uŭ�eM��=���h�&ڄ�4�̻Hמƛӌ��l�K�Cd\l'4K��|�K�F�մFP�E#D�&� "H���L8}�ޡ\�s����%�	Bp�!B4�D�{55Xh�)��RѾ�BJ	��=���C �^XK3�fS�^LG=@P�	U�*�!�(�:X�5r���׾��S9&����  �tE��uz�L�JɅ��g*�Wt�02�rŉL%BT;��؃�<��{KA��3��l݅��\�І�SW�Q1(�H�c(h�|!���D�=��ƈ"h[�S).�6���5 �@4lH 0P&4 ��������M�w�i��S�F\ѹsCY��f�0���#F6H!\�YI��%ā��"P��	�H$��#D2�B!��I�`ň��I
��LJH�:HA�R�q�h�a�&�a��x�q�9��*d<ω�`�q�`z�ނ�
�9^��e� ���eٷQ�14jkL��h�c.QB�%B�6�T.�+mаBbV$�!$�$)���%C��81#3�ֈ\�8ĕ&za�V<=��	�퇙��@
�"����'���O�ƞ��iA�4�cSWxnB��4�R	!"0I�B�符�\԰��=<<.��s��l��h��GP
�14i9�sN�GHoi(�of�s�aK��ǉ�C5���:v<$�b��"Y$P��� !�m��)�!���=@�^�����D4�A&�
�)�L׹�&�%c)������<Th5.MF�6��Y#/�`Ij\ҧ�*�I	Cp@�'��߂
��D��J�Ԕ��`b&,��P�2��h�%�uf �Ҵ��@����3�<��p5�*?qN�4|�K�w�ią_H�'���`�D�� �h�`�<T��r�T��ր��$�n�pؘod.��.S���4 �� 0�1$�8�B�B���yi˙��q�O4`A��ȴ���0nxX�m,�HXj��

��$XC4��`6qOJ<缌��}8o] x@b�x�u�!�Hv $�;�`�4\�����iO�]2�I�)�I������$P� 6h�E0�t&�i�0&4F�"``�5@�Y)�4kc��0��Mh�w�F��z�K�a[a��2iXv�]�v`��]���U1D ʗ�.sdc�e3Q���1ӳ���$����F��B��#��A#f$`AP�@ѓƈ8���}��p�r��Uii�Sq'S\^p��^��~$pAf��f�̼hH!d�xs�48��ܷ�½y�|Ά }o���|Ͻ��1/ �r�{��c�zP!=�}D�M'B�)6d�(F�`@�c		M0��%m�����Bd���Xy � ��V6`�C`d��v�����		�q@CA�K�	i�B45��J��tF�WfLɼ6�s.�W��`�S�'(�~E4�^`!<t$v�b�Aԫ��(��n#h$ecP2��`˰Ppl�! �A�Q�,�߾L8ksy�Ȓd��
a6�	g��VPщ�.����%p�!BBD��H�62^I)��CG��3D�)���n�B�����h��ݹ�.��r���XD�3������zي$�Xdd$��/hr�� �ŀR����YM����$��5�~o�4s[%�_|)��g�&�Z�
$�B����lKf�rh��� r-���ƈDJȑ(� ��(Á��@�!�Ra��F�`��0�J�f��A�K!.&XQ�	B@t�	#)0sX��%�A1 �5�@��h��of�.e��	����H�H�(��V����.�\8��ë́�L9h@�� aB'"]	|xq߳ɗ{U	� �@F� �6,[�yJ�@�p � �2w�<���dT!�h��Ͼ��	>!��v �5y!$�Cc�e���c�͒;�$�p!�h�����V��AW����J��fkFӇK�	
f��5�M������1��"HR�J��	`B�����מ�j��\�_M�
ZX�S^�!�˹tìH
�%H̍JD��Y3Ӟs��|	�ߡ,��<}�ĸ�ay�0#CKL6F�!�!tC[�p�� Q!HA�"BIMl���I'&h�0 F$`-#I�Hp3��{G�^>��0��#Ҟ�J�4B���� �t0�*��1^fm�u=J@��X/�F��,Ç�n BrŀBKӚ� �
��X^�۞׾+�Y  �
0B��lL$2B��¬���-t%��n;���A[v��\4�̢�@�Qtam���!�yh�عV]��vz@7�.�4��6.�{�L�!h�$�j$H�`�0d�J�@NQww��tAVȰ@J�x��Ÿ0N���)㱀Wq:6`�L)�TH@҇�!(8��qb(� � �:Br�R�Zf�2�1j0���(c�!F!B%�J���Ч\�aG|0�G~ ���i��q���0��Q�R�j$)�.s^Jxi0]	H�5iD$�A��S0Љ�t&�� %	�B�233SF��kg���"]��tC,M�%�B�rkI�����Cx��l�"ŋ�#�x�`B�Id�&���$B1!L!��&}���@�#nh�l�c�p�&�n2r%�$���oF���I�!I�0=�E��$HS7�}-ʑ8ф�ǉ�®:��>(�T�@� X�]�kcج K�H��!$&�4q��j��V76˚�cJF���4}�l��K(@�#�H0#L	Ip��w��o.�Ʃ��\%�����eL�f�c�z
nHGF�h^.��a����K/��cv,���<2ņG�H1;��4��zb�x���R��jA��T@TT*����i8��%d�fzZ�����,�2,I�@@I�荆\3%���ߵ�@�D{H�)$ *B�aP"�
iZ!
�B���.�Ow5�|2�@�8VN{��\����@F��a�Z<Zx�ЅpѺk��Lޡ/�]�I$$D��Lcp]��ù�O�M���P?��xל�z���=��#��w��H���h��I�,�c �RZ �pz��a������i`Uh�Ԁݛ��<��[8$:<9��v��9�$��0��  ĤJz�2��Oi��S+
W��$�D$H��*��� a
�+,J��@�@�i�aRRH�H�BHI4H��"H�B Q�@�X	 #CoӚְ����<+R2�/� ���Uu��A:��
�ɻ~ ٭������}���ޗ������       [@� p2 vr�pp���mm���c�2F�[Y��2�����}�A!��,� �XM�H�J�MkN��U:H鸣ĭ��n.��u�f\��0�U Y��ϥ=����7S����*�4�	!����x���ʈJ�<Qtt
⧫)�2��G'���)��c\1-T�^��]ib�bܛe�I��Q��5Unǵw͍������(��2��Wj�ګj_@�O�U��ҫܬp\����2"������3�[s��\I`Η��c��� �v��~���^�p��s����b��X�|�K �S�.۟g���&v(�mS����c6ݢ�+

!�j��W[8�2�b�vn�GRa�n�Jt�ˍ�u���kͤ�K�rB�ZI��x��US[�o\�VU��@�q��O�;Q�>�á��ݝS�T�˜��#I�k,��8���m��4��U�m��/mq $6�,����sm���z��$��.���:�8t�CD��ֲ� �X6�
A���m��lA,%��j���]��;&ALg������PR�[��h7"UUUA�	�]J�v ܻ�A���� oi3�-�#/K�]�Ia#f�m�����9���S�F�ʠ+����)�v@,�W��݋�l�  �R�pm���E�^�Y�IO5ٵJ4��k��^gg����C�[\��n���23m�Zl��E��+b�r�]T+��V���L�N����G��pZ^�öVCr9��u�S��:�VA�@�������X����~U�æ2 �^��Q�+̓��]�x8���p���'e�.=���u�Q��4�-�;z�ʫC�j�p9���b#��`���j����쫤v��;!�UT���0Z1j�'h
�h
�:U`*A�m�Y��uEˋ p�BR�2@���-��*�T����ƺ�\R�ҹ��4n��fN�P�#���m��m����{i�� �8I���y��U�	X&sـ�Lʮٶ�]!Ƶ��d)��<��u3i]�u�<FCx��+m��Rϻ����'�*��k�iy��pp��@ m��WH`s'K��\�esA��Zn�����6��M��m��c'	
��Fw��I��s�ť�k5�� �!%�D�@�R�۷�}��I:m�!t����gE-���{aV���V��@Z�l�AE*�Ǯ�+`*b�M'��[A��I�/gY���js��v��b.Q�`�{2
�T�$�v�h��\+ .�t���ݲ��n��)���A{l�kk��]��`�{��䙮t�{���e裂�Ɯ�*0�V݋�m��ҺŸ�c�q�w#qm�]�jt�u�MLb� �\8�KĽ�׋Ý{�M�rq0n�ku�^r���h'�݅�6yn�g�p��n�h2��']6�0��f�B�	=n�6S�'k<ݴ� GY�NC�[d�ŻV��b{K�c7/O*�G�dʖ���9�<�Y��c!�;�X��{&���J�O������\*x���r\�` ����(N��6�T@ca�A�U>�ق��l�tT9�n�R�q��^T�q��@y@�r��m4���'tLi�l�*���*��Z @��ZE-)��n�g�:r�ql�[	i1���c�����M#T�#�;qE��Cf퐚��ȴa[��\�Ks�YҮ��n�IiV�j<�q[e6����׺�X:V�,LRt�Gn�In��$K4��oB�����U�U۴ gW q��ut�n�t9��NB	�M��Z�&0I.�i�wl�s��*]@gcg�sq��Ry�tn�7xx��ڥ[n�p�sCve�j��/U.�J�����j��(4kp�ș��> ݶse勒	7m��[%%��u���$` m $�"G\�Ͷ�I ��W phA�l�T�,�UT.����ɤ���x-�6� ��Y��4P�  p8�ڶ�Yjn2�N�+��*ʽU�v�M�6�m�Wm�6������+;@�*��m[Ip��qn�$ �-�"M����m�mm knHh    �  � m� [@6�` oPH��#l�,,]��n�Omt���m�4���pct�춮�p�r��j:�d�d'Xl -�6ٮ���S0 �m�������u-�$��i H֭�� 'I m�m� �$ �$�-�   [% H [m��l�Q�,�F��lF�.Òj�k��d�< 0`������  ڴ��KI��7��!�-���mwL��ŽG m�$`NbkC�X:��V��\�nۀ � mm�o�m���  � m��� m�p-���-��? ��Hm� -��,0 /�l�<[&M�>�H]�l�)��q��'� Uu��t�uDѰT�	    �b�I%R��fW��h)�j9 `H�`����Km�n��r���i�۴�gE5�m�ŭm ��  i%�`p ݶ&Z�[�  � �`����ҭUuU*�K&��2  mdv��   m� 6�8 �` ��hHI: %�p�U�kwE��;lݖ��h� ^�l� ��~_���m��b2�4nY�ݣ(P�ŵUR�Ƌա��۷Xd�� mRe�#	[@m�v�8�rI����.^۶ ���i�5��Mm ��v�  Iĵ����&�^K����7N�ebA�oK���opY-�� m�  Vɑ�1�N�@@UU[*��F��2�7��vgk` �Z���Yj��9�W<�L�$�`����(
���<�q��W�)����Qj�.�uKn�b�����*�A��K� n���P�y�[rM<��!�4mcT�k�8�M�i"�:D�܋k�nҽ)�.��o�� }��k�Yؖ��0�R����@���-���ֶ�L�pp�W8�n�nj�f���p �ٶ�F�ÔFP.���[v�1vݤ��8� @ �\V�� �$��-�@���6�@4�n�m��$��` Ҷ���M�˭�-�  8 � k� 5����   �l�[EUJ�U++Q�:���N̅�S+*�T��U.�uԴa�	VRZ�QjU�-%R�r�;S���`(ZŽ%    -�   �X���6�%�K�� m��FPZu�UR��`)V�i^u'����Z�k&��uX���4uۖ� [M�6�սn�ݥ���H�Sm���G�܀UU�9e�Nۤ���I-�B�ֺus|�t}S�(�ʲ�[\KZq��RY�V��/Q���ݕv��lvl:%�(��NY�=����26���wG �i��c�
��YY	�kO/�U�Z�ƪS<Ƞ�UU^Wˢ�P6'���y��8�k8��uU(���S ,�زv�.N��W9o]�`-��M�5vL1@�*�ʇ/fVyS�p]�` [RkX�R����i6�  ��	$J/V݀  [@q4��6�D��ِM�T�YdБ:[%qm����Awm�n�,S��0�-6�m�Xpe^^�+�5@mV�Se^΂D�<qd����O�﫫m��i4����6��#���tv78��1%�[iV���[�����f�:n�FA�U]]�E�6��kmp h�`>i7ܒkd֛l��  a@3Кb�9�yc�Y{s��8Cm�[�Ŧ�66��Ҷm<�Mm�Ɯ�n�8�`���j�QR��U�n�51�P-[)-�I�@�Q�:�\ۖɎm$�PT����Ҹ� 5Up$  m����  �kk�km�@�n�	6��m� #]� m:l�hD�Bl��[oV �knZY�� �a  �����p��6  ,�9$���6��m�8$,6��5���̜��;�|��!����E[T�Uq�T&ͪ��0��v�n��n`pkj
VU��eq+�V��c��yk�MPS�	Ba6�Իeڪ���k/Elpuu�@�Ѧ�hɮG4����t� כ]5� �m���t�;�AU�����]��$�I<l�2Ye��t[N�d�H�^�z�A�Ͷt�N��7`lG�e�ru��[�v�` �)��(
�����P�\��cd0�"N:�m�W[T�U���v�ы��UUA�̪�4��#��C[XYݙZ��Z�
3۵4�I��
�k����,�0���i�n�n�v�m�{Vm͖�h�A�����N���
@�a�Ҷմ�m�l���m� 8��� Zl-�ɀ��m���[F���ݎPuY5�am)V��U[j��1�I,�m�X si�m&�����ݰ�e�m�^�|�}nҲK�d`�i����f|���id��9�ې�`E���m���6�$6e��[m�� �M��E���F^lHu�����WUYv9��k�k���Y��f�n��mK�I@q��MT�uUK�T�ە���,�Ķ��x�iujV���؛�= �����g�iV���7��j���Ν�� �Uk�3Mnr�� hݚM���-�����%��UUWdan�Z� ����� �m�mK\HH��Ͷ k2L�k�� ��mCB?Ț ��*���"`'�@	��L@���B�]ՉD"GB�G`�(�T��ঈ�4�Ū�|�a�� G�qS�	� �x*��*��@�C�
 ��O
��j:�T☦�B,X�#�)�0�>!�Si�"�H���J0
�Z�x�,�IHҩ�4	��X	�ͪ�(1_��YZ 6m�ziT����FH�Oa c�b��ڧ�8���T�(z!�����AU�HC��|��=�* ?���0R
�`$��] �}���~C����_�6P"��9��W�1�1�1 ���~8���C �G�������0E)"�1�W@,8"iW����( v|��> � 6�)�� ��J�j=������Q�4|���*x�W`��S�W���BT�B+F DA� d���DOQ`�M!��W8�O�0H���� |>Q�"���T�U���0�j�$b�Uh QB �<v���>���mC@ ��������P�! �`B#Hd�$&!�
P	�J�W�@B`�⯀�"���d���`�6*:6�O~T�H�*�| }G�RD"�	m-ZE���!m$)��eIiaZ����#O�OP=�!!"� �		"��F2C�]K#F1H�ER�@U0 ���!�d	$�|�TW]�� ��4(% �>q�}!��EE_���I �@�$`���<�n{�m��{?���UԦK���ے�r������n��^�N��[9�S�	���햌�*7/�^$ڗ���մ���ٗG���i.5�l���z�6��%���,����ɑL&^���������魦,�Uәe����9�W!{V8أq�.�&��3�;���97]�[q[�s&9��+$Z�T��3�u��\�y�5m����WY<�#{Z�� ��ƕL��֧��e�ݺ��n�kM*Ե�Hg��K�5xg��-�8����NEU�v��:y�����0Y�)���g]�PX1��b��pc�+̻5u�<�9��s&������z]��=^^·V�]���}m���F�չ��Nw��u�m�c��+��o�
�tڜ���';bWې�t��]�ܘ6+.úL��֒#.j���u�[���z�ւ��n�­V)]���x��@*�՞GF�ܞvy�FPtHeG�M�����)-uJ��ꮽ�T�gs[�l��݇bd�\gT��GjdmPI�����m��Uv9 �4�$!of�c:Սz�\�c# ��YeU���u�8�LP������m�lU<�`8�m��P۶Uxր�v媉W�ێ�ɸ���VS*D�{s/�_O\<�Ss���{;[&U�v��aV��,�5����Ĝp�UI�mEN��K�s�z�ZK'���va����c*�a6X�vN6�U�u�ڳ�&K�	�85�7�[��3�ק�+uW! g������9��̙7�`1�J��[m� �y�V�b��M>���z�+;iһR�-6yVږ��J�9Y��]�vv�nkKv�u�v	��8*��vF3۠6�1-�i�]­�ht�����tJa�ع@5�NRZCj[�\GlڝS���.��-�����c�� ؆��-��H
�R�ŭ�P`*q����[A���V�(����i۩9ޫC�ۂ��;8L��7i��)nf��٬�[�[Z���Y�����EP
��S�
�©�pL<6(~�)�b��|$P6�|D�_�~t�x*��HK��'"��Imr��\�nݳu�]����9��������r�pD �q�Q�ۗd�q��∸5g�x��N:��18]C���[�����QǵKiφnN�}ٶ�a6�6�\�7i��)e�m�g����m�����A�8܋F��CC������ɍ�-�� 	�F��y���s�(DJ_<�lF�1$�Hp�{�߾�w�z�w���=��o���˗�1�ϻ_;/<�=�>N}�o)�2�l	-�1ʄ��K$�{\$޵ο�����_{s@�p�q�����@;�٠}Z�z�n�^v� ���&�i�`��@������� ��y�4�2�Lkx�q����yl��٠}_]zXR����(����� {��;�� ��,�(��qU2��O��<�W�k�/jp�rX�[N�	���w�R5��E8rU�t�~�[�^��Z廚yl�>�W�� ӑ�NK$����"+h���5�B�j? ��榾�6nI9��M ��:w%�ә&L�!�9�h��`�w�L��� �Mt�:��	 '�JLds4�٠��@�}ʴ=��}�h��8�$N0i���]�kS��^, ~n�_����@�?�0�"X�r~$CY�i�.�.T�Wkk+�{Dc�լ.�/��-�#"�������yh���yl��٠�*�"�ɍ�E�^v�h�w��� {�9�ID%2t��+�Hd��D�� �}���I������K
1Q��	�RH�6��P���Oou�$��ur�4�RLJdmɠ��@��*�/;w4�٠r�^��2BLp�94�­�s@/-���˝��if���3:��#��E	ݹ�U�7�N˝�q�8ގE����n�]1�գ�������yl��l�-�C@���L�@�ELݪ.�`m�r��)��>���hh�n���]qDH�`�� ?=w�6����ذ�����uPbi��Mɠ[n���u��ۼ\��SqR-Q	TL(b�@2�ޖI<iA�0�	a�۰�7��`m� ~z� m���w0�������l�&�����2SXqSJ5�!�v�� �ۏk���vwk9�un�1%�V���}x�����/�}�����hR<Jdmɠ��@����s@-�hZ�͍� S���h廚{3�${�����h�;����QB@��	$��w��׀z� m���]2)���)3@-�h�������݁�o�ŀ+I	�<�G�(*�);�C�.%BY����}��p��8��zwk����l�x([=eХ�v��NL�f�I���/on�ѱ� �x��3��_h��C!ڋn�+p��X8�����]$O�|���/5�rXě`��o���6�"�:�T��t��\g;�w���Td.�ϗA4�ۤ1ڻ7n��'R�lf�c�'g�ا=Z̝�y4�[O4�n���Z�s�'��w{�w���u5�8�'\g�m�R��.NMB���"��X�]�']�9y�s�QfviI���M�t4��� �٠wt�CN6�hp�M�k���ș�ŀ�׀���#��"�P�ۙ�w���m�@>��@���4�)FUX�hH�s4=��L�w^ {�^��X���X�Z�W�%#ĦFܚ���׹�o���ۼ�BI{��蛙������SRo1n�&N�粺J�4b'u :��=;֒$�58�hd�|=�=��׋ n�BK��}x�]Z���Ww77WWV��x��yrD"�rJi�#
�i�,$������ji �4��	*[[�>��VU�(d��,�s���Nv���<��tȞLo)1
L��f�^����)�^[��w�5�dQE5%]�(�3����7� ��, |�hŝ;SX�i&�"rh^�L���������w�{V̩k[����;Wn��+�.�c��D�g���tT�ևnֱ{e;;��n�{g������o =�x���{6���*�,i�$dnf�^���~����@��x�>������	�%#ĦJ������5��0��.�B"�I\(p�����ͻ�=�]"��x`�q<qI4z�4�n�^�� �;f��㿋2D�L�F��8h��X �]��]��m��Ӫ�M��a�5��7g۰�Lv��q<,;M)5��&����8�y����n���7}�� �k�^ͳ ����7©�r(��Brhy�7ؑ}T�s�ۚ{�7ߒ=��_6���i&�"���� ������ 7�� ?��0@��JCd���I=��rI����=A��D��~ ��@!UN�+�O |x��(�M��W5k ���}�|���?=y���l1�x,qG&��!��t�F�q	����m�z?�Z���۬���k3�Ӵ�)%29$���h�e4�n�s��@�Ԕ#�c��h�m��%2{�b�o� 7�� ��p;��2I���@�۹��l���h�e4����㘛��O�I���x�������,�U2쉨� 	!94��xYM��b�'۽,���	�T�44$����v���2:C�cK�mv��N�.nN�֭4�$+���Z���{qq��ng�9���u�:�t�Jqt�t=l� ]!�	���m+u��m=�Uo 팻��:��bͷJ)Ǉ�֔��������?9x6~�]��xe��M�Ս����ƺ��������Żu�uF�	���i;)ʱ���(CVAw3dH�
[��e�ٮ䉚�\�kV�)�Թ���1SIO}�9ŊMx���f6x�.6�v�N�l���u�.�Z:^��iz�;�tN�t&�����m�~m��n���w�a�*W2<�9�n�{w��N����K|z��$�@���2�DF�v�I{w�bI%��ZI-�-_|�\V�=I%����\M�9%rI��In���K|gr�I/.��I.w�}�I���`�s$ǑI&���ܳK����$�[���I/7�ޤ�]�ʤ2~��	Ɔڏ���kE�swn��v$�0��:_m��I���k���o:9��"�I/-��I/n��I/7���UT6��3�bIoO�����f�M�ћ��|�ߵ�=
��R 9".%`��R�;G[��moRI^��}�Iqv�=I%xdK�F�0�II$�I/7�ݤ��ܳK˷q�I%��ϾI+��V�!MD�̎7i$��w,Ē�ް�$����bIy���$��k�.#%��&H�K�zô�K�ޙ�%�����^��1����δ~~rdt�`��K7\�뢽�/<F7]al��Zr�Vغ絞9;`�=�nmƛBFF�?�I.��}�Iq���$�8KW�$�n�Ԓ\�:"��lqA)��'�$��o}����{��K��q�I%�vϾ�g�m��������Ldq�I�g�,Ē�޶m-�Y�|h:���>�|J��L����#�����.�l+9���S4*�`hJ�m�ϸD]$d
�J'5p�����H(�<��0�_Nd_de��I0%�L߸h���\b�3�x���d���p!s�D�5(M>��fg��O>��w�Mhxp^�\��لD�M��yr�^<A`DcB`�"\v@_B}��uo���=��41��HF3F.1�{d	���C��}!qy�r\���@ F$�XX�&�W�(K�?��'Bh3q�߉�i�0c!� |�6�l������XM�p|5�}ˇ�_d�{hH�b����T �7z�%�2���Ux�`�R�J0B����8M�-Eo! 1p3s{��q���K7chP ��! �'7�WsH��S�hO<�|�4��h�#�
� P�c�|<_��C�UE_�բ1�RAd�v"���} `��h/��P�w���|���u�T�O�=I����c�%��K�zô�K�ޙ�%������T�7�/�I.��Zc�"k)1
L��Is��1$��sV�K�3�f$����i$�������\����Q�p�k�m��<=v '�m�˺5v5Ʈ{i�ݳ�jS��a$G'8�����$�8KW�$��n�߀�����}3K�#�lӎ8�h���I/x���Sm-�I$�{阒\]�{�߳1�����{Dx�IbI-�I$��阒^[8�I%���}�I%�Jc�QcLx��5$��;�bIl�-$���r�I`P *�="\Z�(�"G�48+�!&(� |�� 7m�p�I,��%�.(R�7$�I#�e���|P|��[�\6�Is�{�$����#M⌘��L2NS�6b�{�n��Z�C�Vw�8����b{g�a�HǓ�RRI{9-_|�K��I$��g�$���MI%�俇H(d�$J ԋ1$���I$��阒G�8�I%��}��k�������)!i$���LĒ>��ZI/x�嘒K��I%s�K�F�@Dr}�I}�ZI/x�嘒K����^���I.�.��8�hqGԒ\�-_|�^�߿U=�I$�{阒G�yKI%�� ��<ʘ(D�%ϲ��kF�a��VXn2;8�;IR�L�{h�exӣ�U�Hvv-�.2N�!H���ùL]�m�_�)d���y�.��ѵbN�y�����SQ�x5�£=���2�Il�j��������m�鵷��M���7OE��9h�S�Z��g�kn��ԗsՃ�%#e�X��5�X�W<�k��g�/gm�bMp����Ā���Q:�k��\�̓Y��.��E�v��.�uN�C�m��*3�d�6�;��5���]�X��=�����������	$��阒G�yKI%�ܳI t�t�,i�$L�ԒK��}�6��|����I�/�I%�݆���i(�26��S#rO�I#��MI%�����m��I$�{阒K������(���^��1$���I$��阒��e�J�'���)"QcR/�I%���I~ U �{��$�ޟi$�rZ��$���ra�d#�&)�,���pl���o4��;d.�GT�M:z��Ob����T�$6�I{��1$��q��K���
#�ۙ�}�Y�33ɗ=_]�HU��I$�I#缥� UP�*�P��{�K��5f$�>�ٴ�K�ޙ��C�������x�L�������嘒^{�ͥ�����1$���KI$�{���00�-�d�1%�
{;�f�I-߾��$|�����7�7��1$�����BD�5$�ϖ��I/~[;�1$����f$����i$�UP}���r��n����s0����R-�TJ��i���=�n�k����~͌}Ҏb��u$�?�)i$�L�Y�%�l�B�|�K����Iz�Ǧ��)��)i$�L�Y�  m����i$���bI}�o�~��^�K��AL��B�f$���ᴒX�y�,��@�� ����Ff�-�x�p8(|��]kS��.�m���_|�\븴�!X$��)!�/~�o����$���)i$�L�Y�/� 7��CRI{:E_��7 $�q��I{�ZI/�� +~9�庒K��p�I,}��K����9	�:���TD�ڟf�v�(�Y������{	�6.�&�/��w�m���MH�x�n)Ē]�=���$�;vh��P�~�������O*�.��U �����y�J>Q
�����]w��9��+�P��?_�1Zm��� �S��=��8t%3�S��ot�9��B�ڑA��N=f~�]�}8�O� ?y����$�	JR�B�W�)X�M�+R����>=@�9�n䓽��L���(	�+$旼���A{~�ay�-�}�@���;�l��S2,*N�!'us�րuٮ���ݧp�\oB�����~��M��BDL�(��\ �����Z� ��\�I%�ÇӀ{_)�U]�T���TM���k��(��$��n���7�� ?y�Έ��NZT�뻩���%'#��;��VI�/yY�B��B�l����W����s.q�R4�27s��%>U�Հ���=>�XBI}
")�wՀ�|OʭM��
������u�}�P������ ���� �P�iA)�n��j�d��]���j�;Gm���7F=Op�\p[������<��s�s�5�4�#́Lh닜��8@�����tۥ��ݭ�մ��N���v%N'�'vz��KX�@"T�A���w��i(iN@�7�=I�s�h68zN����=��̫�`�۶�y��gv�3(��'�#�u�3z�N�.e�\3�LkZ�ԊkT������A�G\�a�L�9�oz�>"��N�̘#f��\�թӓ���u��'X���2<ՐzDdchH��}����Z�u��O�����!�}Հ>)t��*���T���Ӻ�?�}�Q�_�V��}X�Z�:!%2�R
U�D���h����w��ӭ��&wi�����/1��Nd��9Qaz߿g��Еm��V �wӀ{k\�tD(�*���9o�i��&�II����>ՠ{?f�;償�|쓋{��wF��В8�1�N���)U���؝�X�ўy��k�n�8�qÝW~w��ݺ���H˫`i��ƺ}8�+\��[��
�u>���I��!"��&*Ed�����Ex�#p0mR6��U8 hF�����������E�8�mSN+�T�&���nI�q����9С$����O*�6�$*�]����X�Z���϶�N�;�:���� 7��~�Ч�o� ��� ��k�J""}Z����Iz6���Š}��h��|�B�3������?:�8u�8p�� Ţ�����tQ�s��fmr��^�g^�c]��~ww�\��}m�b5�V�}����8��쓜���X�����'����H JD�L��q{y�� �Ԓ�7�� ���~[Z�:���ܧȇ�JO�H�W|���M埳 #@�P\B ����l�)�*&0��LR���`�4"���{3����{�7$����$i��'#�C��3��n��<�}8�����I)�[��9oؤ	I0�N$旼���P{�<$���hs���T���H�����c=�x���9P�sնݺ�I�kX����#$�
�!P:D�	�,$�o|��^��?{m�
�!�S��NW�ɑ��"q�+��߿~�H�l�r��h.v������Gh�0m9#ƭ5u�{]�~ҵ�DDD/�"V����:��������	`�Q�49DB�>e��ӯ� ��\�8���X��X�h �HJ)D9�5S��ϊ�0G4��$�\�BI���� ��U\]�	��.UM����� �!|�BK{;����0���h]�b�7���D�'�=�nú�u�gѮR�i�V�T��G-�v<��绻��&-0S"R~JG��x�>�e4�k\�DDB�!��Հ8�u��R�Wa3w7f��l�P�$�O'O� ���d�ݜo�  ?����BMAL93V`N�N���aВ���w��w� huKWd� ������
#�	V��� ����?{m�(Q�Jj�� >]+�.EtQJd���`�m��D/�!-}���j�� ��x�Z�� �r�0!J��su��a�M�7�+�ɶ�JR��S,-k��5�h����R !c@�`�bFP�!$�3� Z�@�;��v��3���~�ͧ8f"�%k�M��]Q#�v @#<��H!D!�d<}b�$��hS؉��ҙ��$$�l
�y`�� H1bF���d�a�����4h1+�c��BF�0bD�b��"����F�B0$�������@��I�����a͓"�9�m��`A�YM��9���SU"���x��V3��|T���jT�ꉨU����� �S"�f�oF��>>�=	:%Ͽ��U*�3s^6Ne�㐸48F��T��}Ӯ~Ba�j`����z��\{JۥP�`����fۨ�3�¶Bq����h��ܽ\��)Ӝ�D'���v��$�VG�t��u��Μ�h{@OF4�Fy[c����Xx�6�ۋu�� �1 �qnz;	n��[{k��^��ݬ�=v�wK��aj8÷3�m�L�::zvzF�r�gAˈp������:6�1,��86�9��ѲZ���D�K�x5g�����.ma��g��;�ؕ��v<l-�Ο=�<�;s���Zڦq�̍.y���C�p7U�Їn=�/Yw��qѠs�P��і��@ٛ/;۷iqԵ��E8�ɷmrm���؎1�׫]�\�W�/P���s���vp�Gs��5c]����7l�� ��(��w0���N�Z���x��]�D�w>��;s����(
UU�e�D t��[�k�WcGe�ɷ;-mj���v����S�9�g������Į�h�� m,�ͧK�YB�=rYnܝ����{d�Mk]=i4���:�q�:�S[U��]!�I�Εvd��H��V��8�-��IWj�@�k �Y^�w]�/祁ŵ7g�^�Eմ.J35<��u�vحj^\s�wg�7���]�sg�0JN�:���5Rjt���N�V8��iV]�Ks8l��%���5[URM2�m���r`­\On�8��X��+9�r�Ol����i��5�����'0d�viۮG���vT�u�=9ݎf�U �:�X�g�!�v��v�|��κ2���X:Wk=\�3�Jַ+�.���k���x�#�!���WH���*���CJ��&��  EfXazፊWH���L��q���gjsg����}fn68�B��v�Fzb�ua�m��]����iܛ�b�q�/��.���@�����7	����ݎ%t��I��»����9K�';�dշC����<lvx�7���Rhnt��]\v+B�	é5r��f]j��5�&(p@�|E<4�t�x�'�qB�|�@�u �4����b�}  �A<E>���~o2\�L��=���v����t�t�r��"�=�'V��k��\<r=R��{��1�ٻd�G䰱[snÊ�g<u�h�&�sV�]�cv���\컇%Y�m9�6�4�64"�b��8x�`�A��'��j�5̩�O���5x�����;6^���/W)zݹ��z���0�t��MŎ�Q��M��n'E�N����:��Jq��\њ�;�&���re2JkH\�ևZ��rں���3�u]�]=�?o�����D:;hZ�{�㯺x>����r~lw�嵮p�׋�P�Ho� ;�󈠓�#(��pk�W� ��T*�}�, �� ��g(IL���uU�ڠ��Sb����� {u�/�P����4����>幯��II���$�L�}x�����t$����f�VW��1Ǒ�JG&��;)�r����}� =�� 65ʩy'i�Ӂc8G�2�gZ�G^r�#ky3Z��ٯN1�/[k�������x�06~��t��� {u�У�
=A��� 8ܧ�w3t��������ˀ@�H�H�H4hЈ!I"��$V	��E��DJ�	D�k}x�|`��s�B_(IU�J���R]R��U7k w׀~��0脔ϓ���=:�����R�l�<&4�����s�|h���~�k��Jg[��|�u�*f�mEHl��_r�O�
����$�w��9��h��T�!8���'ܘ�m�Id���L3���4/�ۘ���w��}����1��"�$��.�= �{f��6��DB�"�5u}����eAt@L��T�� {u�tD)�����t��;^�f~�����g��q�Q�$�rh��0�i���a'	
��-B\(
��>�d��w��9܉�F����F�f���$��V�Ͼ�e�Հ�w���%Z� `1�+TT�N/j��A{w�}�O��pk�VC�B�c"d��""nI��?L�ݶ�Z�:z;I��k����5�t\rv�o�{�Վ�k�r���� [}4��M�;W�f~�o�����yLL�&1I4����P�Oq]Ӏzu�`�w�	D�z���$	�?
C@��-��ׇB��9��]>�|���.�ݫ�$����D%�J��� >���m{�ܞ��Ճ!J�B#�(eT��݉� |)��S[�}x��f��xLx4��ԏ@/{f�DB�$�}���������u�l�?���t 5])6�w#\n:#��F␞y�1�n�vn&���%�v��{�Ｘ�̝(0��L$�>�Y'8��d�[��(|�����{Q�b�""9��t���/�(��g�������Z�9,����C	�4�E�q_y���Ô(S:����N {IL�LD���&���g�Ľ��v��}Gڴ=�31q�y����&G����=��p�"#�[�}>g�����"��DB������ST�ju�gt6K�\K�����	���]�ر�.BEw^����e��;v���Ěcf��f}]s�4��Eˉq4�ݎM��� �,lR�n�yau��͠��em�Q�D��v�����v���Zen۷S���:�%���N�v+�,�go6���v�a����u��Q ��unҁ5[�<��i�rwvcY��-S���׽{��I�)�Yέ����9�V]�ۦ���P�;���c�7F�������`���0@�Q]�W�8��� 뾈I~��O� z�3�BD<���Z˶��?$�׀k�Ӏ~e79�27��	�H�������o� �ֹá(S>⻧ ���/��V���F�rh{���:���⻧ �:�`r�Jg����G��dDC"�>��Z�fg�I}�o����� �ֹ�?6˪�f2J#5�L[vP�x��|ڌ��'<-�<ݹ�;��<ۇ�?~4	��@�i�$��K� ~�x���DD~���p�Y�z!D6�(17�^v��߳�� ���B��Y���=�gݻ�r��g�(P�I(�W�%���,)Q7w�>��p̭s�(J&}/�������BBqE1(���f~�\�N�}Հ����$�T�;��9�C?����r6�"�>]���l�O��+$�����|�ph!��
q�7.{�&�O\1q�دJm<�������뷟������``�S����$����O�������%�C��� �tOr��.�
�����mk��#舅	*�~+��g����]�DB��L�}2Y��̐�`�Z<���>]����P�b�A�"�*4 $d�QQ��A�Z
�
d�#��{�':*{gy�5�'}ϻvI<I�@��D4Gd�(UK��� 9���Z����$�U�d����g𿉊!��&���٠rJZ����S�X��� �"!J��r��n1��eq�s�6[����J7�h�O[��ۛ�����Ikg�5�t�pΥ��?N�_(P�����_z1!8���qhV�{��ЦOK� ���mk��%脕P��3�I" �m��������I%3��N��u��%��Y7��H�=���o����k��DA� 1�A��^�ϼ�|z�y���F���$�9�ڴ�N��?N�X ����(�˧���}v�ԝc�����[��[�Z��ێ8-	�4�XP�/��{�w�c�ݮ�գ;4x������u���G�t�p�z�= ��ƞ(�z˶��g��ذt�pΧ]g�(_(U@���~�M�(17��}���s��i�ىs�_=���@����*��� ?�8�9%:����Հ~�n��x���ЇX�N(�%Zծנ{���}���ذmk�+ �!~[��wvrUv�v�<��X[�Dӕ����t;H��^�7k�u�֍�SH���m�qm\��<F�x�{/k�ݸ仑��u�Nܚ06�\${\�N�
v%n�u�fV��Cقn7�K1k����"m���N5���oX)4�eݛ���,e���x����:�:���q�y9n��t� �'h�v�Fy��s�<��v)�Vۈ�lA�xd��y�?���z�~�P��ŧzAL]rw!nwj�Z�,�pfL=�]�k':�Ż]���O���s�fU���������`��<�?H{�_V �+�'�����I�y۹������h�W�@�v׿����#߫��<��#*�`����N���3�}Հv�ŀ}����L�E�ȴ=���=��=-�`��`|�K�og}8�� HPa�CL(�vIŻ��? *�k���t�pΧ]`B�s�� �T�7��|G�{Rގ̘#ns�e�,ȱ\��e1�u�����^�ܞ[FvUŜ4�������Œs^�Nq{��
 ��.��d�.�译PF�����d�k�W�(!V }+���+i��l*�6l��!��[
rw�a�aQ1Q�!�v�ۢL�@ء�]ro�?yw �~���x��D(�2�($��ff�nmL�\��N�u��䒈���������|���w�Tӟ�<r5��� �:�`��`��8	O���@���g�8)15��=�s@�Dk���qO� ������ۣ�I�1��'c�n�Z{�Nݫ8K=�.��c��u]���wn�_s=m)j��~]>��)��?m7?DB�(����ŀj�Ϧ
EZ��䠫��?2��ޭs�?kŀ~�79�B��QT�J>�R�R�H.�p�� ~׳sET(���G�}��n��:��Ы/���5 X�[��
g�-�Y-�����3��^ii���"�[c��</#�P��S^����T���)>/ O	d�Zh	�T�i�Y��4�����)"3L�@L�� B"�"�����Ą�R��p�b@"���>��|��_m�I!A"lX<�Ӝ e���#����#BZI'�OM\I'�E���VL��ɪi�r�۲�	�`i�������q�"B(���C8�.��4\`�!��0!��L�Q�;o��>�xsFV�H ��O|="�"I�y�}�|IB����TE�P��U8���M*iE8��.*����z)� z���`�����
p\� |���*�����o�Z(��ί��"6�(�n,J"{_~X�wN�2ـz|�`�S��jK��I��r�O¨��`�I���d�ou�$��F�4D�݋C8|���C�
:��:T��'mqJu9:�]�!=��2-�4-�4�1���_+� =�� ׯ�(�%	z�������?�Qd�1H�jE!��@��ŀ{����ͳ9$�L����Ur*ɻSR����>ŀ{����Т"�~+��@-���α[�B7 ��������}Ӏ{�}8�7x	lB�$��2
@ ���O�@�ʡW�2	D0r-�>ՠrJ!)���v�ŀ{���B[���c�[�5S8�&z�.�ˬ[%�؎g\�'�h$۵�/l���t���<�T���������`�7<�D~�皾zܫ����`�x�#rh�x�z����X�7y�D)�ҵ����25�Nf�޿yhV�^����#������nh{�`���QFU]\�}���߲{������x�qڴw�B��� )�6�z�7x�D%�＼u�Ӏ~u:� �QR�����{e-���їST����W.���$ɚ]�z��Zg<ۙ������7al.׳dN�G[z�76�7#l�Q��]�{N��X�]qS�u77T�v"��n�N��Aƃl�=R�R�]��:Jwhu'g�t�vx��f�)`�4%�̗l��H�r��=�]g�[D0:q�j�Ͷ�����@m��jC�x�؜��42�K�cL�v^�f�iY�/k'�_	��4��9拭k2Lђ�WZ3��>;��Yp�]m,î�b�݅�)�`����d�k�&nG0�X%$�������@���h9�4��]���#jbnf���}��$sþZzy۹��߱#�|���c��Q�@�}8�Z�ℾ����ذu�ӀՅ�1<x���-�}�@����?z�����[��NW�-XUK�nE�^v�h��g�����9�ڴ*���$LSq��(��'c�n��f�������>7�;��Q������tA��'3�9��-��k�9�ڿ�3����^�`���QF7Z�L��|�"r�����,_BX%�/�W��Vl��ذަ� �{�X�yĤJ4���9�ڴμXr�3���=�>��7PM]�HA"�p|��BO���Niza=_�.rv���W�n�mLM��>�78�V��=��8��X��DS�����1�=���sQڈ�{XٻY#]�����m��ﺋ|s�kX#;5��=�>�ޭs�?k��􇶻� <�/c��E&qh��Z�n�����?2��rJd59\u�j©0��Ȭ����,��}�ʡ@D���j!�4�Ap�^�����.�}�v������t �X�F�hqڴ�Z� ��\�tB��ߖ �����n(��-�>ՠ{������������@>�*ɓ�`Lp"�O[n�����zQ����MF��㞤�r]������n
cR%cqh��Z�n�����(�^�ߊ� ���	��wav��I7s�?kŜ���OmwN�)��9�ڴܰn�d�F�&�h�M����p�D��>���,�sc�(��ɛ������BU��N �wӀ?kŀ(�1䒉��s�	��+��3$s�Z8�V�����}�οyhQ���B��LpMd���x���s��}�s���cT�u�f#<��E�Lp[�i�	�Oq��{�ۚ�w��s��_�
1���d�!��W�͓w*��`�M�tBK�~+������/;w7���ċ�P�z	����n8�xw�@�j�>����v���B��cR%cqh{����w������}�ռg}8�}7PMcq)15�R-�۹�fs��_�?�w$����&��_V!B+C5B1���K�b��޽��w��������2�gO8��5�ɭ�[7Qv���[���0�˷B��ѫѷ).��\������g�!X�NKd�^�n{a��YЯ�m�@l��=�e�Y�F�S��(;�v�v��iJX��+uM�vȱey����b��6�u�Ý[`�m8�0S g��b�HsJm���k�V�mgs������'I�&�T�N�6Y����\�±�[�NA�O���q�w�{����08y)nM]a��u5�u�Op=lܑ]<���b�=pW1�8�n���}���$ 8������>��V��>ՠ}{w4��c9%�˜���s���T7]���}� ��ns��z��2d`̑�Cqh�Z{�ŒsϹY'<^�I�:x�$�	m<Q��Z\��h�����ڴ?�B��)�� �O�*���l��U%�լ����?=�f�V���ŀ	�NQM�[�N+����s�f�4�ԑ����E���8�]��#pF0R TNY��?=�f�V�����D(IGޠ�������a�#pOyJE!�s����qR
�E "� �h�\0
!}�d�y�+$�j�l���:�7�X�"�/-��>�i����\�SƁ޻�s��7P�! q��3@��ՠ}z�4q������KXŎc"��@��Jh��!n���s�X�Ss�~�T�E�fBr3Z��\��7�>mN�'3�N���󫶇�m��Ʀ�@̊L�Hh��Z����v��T��s��	�Oq��on���@��)�s��o�G�J�	�&�X��h��n��믦�������*!�a$�BE1WG �   �_��?o�b�:<�R��L�]��Uus���ߏ�|`�}8������yh�zE7
C ��]`%Ͽ/�{k�p�;f�q\�@I�`�pbq#��x�M�er�k��+��v�jC���ǟ�����o�p�$��_nhqڴ�YM�}�@�s�n���#�G3@��տ߿DD*�x��0/���^,ƻ�*�A��P&��Y'4��d�y�+?�_�(�T��`�� d����
�ڲn�Q	%;Z���ذަ�$���p"1�	����X�bDB�٘� �x���*���\��`z�`(K�ID%�>�||O�@��k���"���G1��V�k�����C��P�ւG����F�'�t��6u�4����q�FD�hqڴ�YM��u�
G��ذ��g�T����]WW8��9(�&ξ�y�f����?$w-��IxH(If��� �oDB�3���5�|hԡ�yQ)15�)�����{�f���=��`}
��}Xi�U�h� b��4��Z:YM��� �׋ G���_�bJU7�12m�`�`{�=f�\�/�i<<�k	A��1��GY���x�"N+1����!#�}[�Ӭ��04��j|��
�Os���:�� �@�dH�>97�|fc)(J2�2���>5L�f0�l"�y�ʚRI-�`"Ve������ל�II$�I�F�ƺ�m7�A��j:������ڭ�����n/v�'z�5o�Z�Kgr�T�f���)cF�ΰ];Z�ᵡɎYSe�Nq����`�b�[T�k^քP�mAֶݰ�Jҽ,��Ys�s�(����lK�N���F���y�ۺ6�Kgw'�tE9���2�t�d�餦�m7h7X��ݮ���;n��ݑ�U۬���Ǜj�	Wn �c.�[l���u�Y���UN��Hq�u���٘��\��
E�a֧�Jٸ4 py^��<u��c��+��[`(���;En�(��'������n$�����Z�&��!�J����3m����˒�u�v�0�<m�G����<��/f�؆��tp��:�f��Fݳi����U��`�c=��Xƀq�����Wu���q��;n͢Q�I��8�Ɛ��5�&��Gh���m�Zk˸�ɵ9�����76^$�v:孺��j�YUM%����q�ղ���m���vj�m�B��7GV��%1'M7�m6�:Z�%�y���--��;��P9ڙE`Ne&ɕX%%��l�U��Pt�cs��n^��eUh5@�3���3ۗt=s�t� v6lX7��j� ; ����]������c�Dq�1�#ּ�1h��d��B�*q�H�IVntևg�e�`ڮ�)Z��I���'q3H;��b�j��vl�6(3����%���Vһ�[`�k��jY̴��9a)ںy:��ݢ:�(��a�u�&س��s�lO\*���g	��l���yy�+�n.V���C���W:uk��Ω6/^�[d�I6y.��������Cq ��2g4q�5r@�F�k�8m��HUEp�!=L<b�H�s�`�;�=��GmP��&^n�\=�6���������n�����ҚG)�\p]v�[��a�]����\g��&�6��-$��oe�,�l,����!k�Kh���Ѻ�y���97d��8U.G��p�]�Mǣ�XzvnE&6���Q�O�����T*	��PЍA�([T>66�_L�U�WF� 4 �M.���{��w~����ԏE�x�ul�����8q��8k��uĆ���G���g�Mر\�s��[ۨ]�f�_Kf���0F�Ax�c���6���\ݔ�W�u�7=���.�����vVܜ;c�]۝�
J����+�ۣrFew`:�!t��A��6蛣�ۂ8.z\b7U�s�e��b�\\�{="n��]�nQ��$=�6�^�g���n�����8r��I��tC-�kU�34�6J`L-9խg��p,D/k���XP�O~{����:�bC�Ȧ&�"����@��k�<���!/�G�5��N /���?*�n�L�L���8���^���;V��KlϢ#�QT9:~>�-XUM)�������,����?h���� ����q�FD�h{3;=�r��4.v�~�˾��4�P���Q���-�S@��k�9{w4��Zm��?��c���½���w9��T��ڢ)�.õ��gq�:�q�������Z���d*!�NP׽�h#A�߻�ND�,K�u�݇�I�L�bX��~���Kı?~�n�?a5�V�E�[u��r%�bX�����r,+��h6&�X��]��r%�bX�v}�ͧ"X�%��{�siȖ%���:�"�R2YRCh"�'�뽻ND�,Kϧwٴ�K��=����Kı=����Kı:����E�4d��r�֮ӑ,K�����m9ı,Os߻�ND�,K���ND�,,O=�{v��bX�%;�~/LԺ�,5u�R�SiȖ%�b{����r%�bX��߻�iȖ%�by�۴�Kı<�w}7Ch#A��DE�X_H[�3(⃳�ي4�ql�Wb�M���SM�P�n=����e3!&Ki��.Gt0�F�4��w�6��bX�'�뽻ND�,Kϧwٰ�*�șı>ϻ�6��bX�%�������5.�����ND�,K�u�ݧ!�D#�2%��g���ND�,K����iȖ%�b{߻�t0����h{��QI�ZiGF9��ND�,K�N�iȖ%�b{����r%�Ą��Sh�1��E�:��Q9��8m9ı)]�NB�B�����w#�vU�Ҫ�u��5�M�"X�X��w6��bX�'���6��bX�'�뽻ND�,�̉ߏ��6��bX�'�߭�%�Mdչ��-��m9ı,O{�xm9ı,W�u�ݧ"X�%���wٴ�Kı=�~�m9ı,Ouޖ�λ;�"��^ܬ�LX�zԺSn\���r��k�8s��r匑N�+��iȖ%�by�۴�Kı>���6��bX�'���͏"X�%��~��"X�%�׽�v�,�4d�ђ]j�9ı,O�;�ͧ!���2%��}�ٴ�Kı>���6��bX�'�뽻ND��TȖ%?~���u�Xj�Z�֦ӑ,K��>���r%�bX�����r%�bX�{���9Ĳ����2����$-��`Z���]f�kY��K���2'߻��iȖ%�b{��~�ND�,K�N�iȖ%����K������b+ B"�=9Q�Tؖ!����4MaVВ�tT�'TwA~�O5石iȖ%�b_{~�\�K��Z��j捧"X�%���nӑ,K��ӻ��r%�bX��w6��bX�'���6��bX�'�{�ߖ�~�v{IC�=��O�7jb3ێ���hg�����:��k����u���F0?dBur�f�Wi�Kı;���ӑ,K��=����Kı=����Kı<�]��r%�bX��w��֦kZ�3E֦�ֵ6��bX�'���ͧ!�H"X�~��ND�,Kߵ���r%�bX�zw}�ND�,K��oܓY5nh�Kn��ND�,K���ND�,K�u�ݧ"X�%���wٴ�Kı=�~�m9ı,O�>��:fj�Y&K�Y�iȖ%�by�۴�Kı>���6��bX�'���ͧ"X�-��~��"X�%�׽�v�JCP2T��a��h#C�}ND�,K����ӑ,K���w�ӑ,K���w�iȖ%�bA|N��ow�O�͑]��덗8{����ޱ��1�Y���E'E�ݳ��w6r��,�A�mΐ0t��۱�b��/:ws]��W&�˽�m���B�<.�;p�U��i�<KgZ�+:�7f&;);f^�RF�L�G��{v�;u�A��f�6�Q�ά��"'P�˫n�v���Q�q��[ fʐ�nm݇9�h��'B5�uv��؍y�[�1j�����﻽�{���o��|~�VT�Cv�<g����]�r[�sP!��)�G=�y�l<����n���]jm<�bX�'�}�m9ı,O{�xm9ı,O=�{v��2%��5�|d/�)!I
HN����.K
���k5��r%�bX�����r��L�b{��~�ND�,K���m9ı,O}���r'�VdL�b_�_����sR�X[\Ѵ�Kı=�_�]�"X�%���wٴ�K,[�~�pI��wfԐI��d%��\�)�sI�$�؟zw}�ND�,K�~�6��bX�'���6��bX�'�뽻ND�,K�����5��a���SY�jm9ı,O}���r%�bX�����r%�bX�{���9ı,O���6��bX�'���Eֵ3&�0�-uƸ8ό:�l��5�FB"؎�pb.˱�X��Dѭ\�r�kZ�r%�bX�����r%�bX�{���9ı,O���6��DȖ%����ͧ"X�%�ޏ���ː�ʐ(�h#A��뽻NC��_@}Q�R���ND�5��iȖ%�bw;�siȖ%�b{߻�iȟ���,O������)��ԷFIu���Kı;����ND�,K����ӑ,K���w�ӑ,K���w�iȖ%�bS��zktK]kR�SiȖ%��D�_w�m9ı,O�w��"X�%���nӑ,K����iȖ%�b{�w��LF�aG��4��ho���"X�%���nӑ,K����iȖ%�b{����r%�bX�����֐�sD2�s�ܶ����<J�mf�O������ۛ��1�ۈtO�u�b�ڹ���Kı=�_�]�"X�%����fӑ,Kľ��u�yı,M���t0�F�4��3�@��I�E��f�ӑ,K����i�9"X���[ND�,K����iȖ%�by�۴�O��r&D�>�?~'&�9��1���A�F�����Rı,O{�xm9ǚ��eb��Z,�\bH@�8��&Aq�N�Ч�C�ؙ�k��iȖ%�by���6��bX�'�v��ކH����JIt0�F�4(#C~�]D�,K�u�ݧ"X�%����fӑ,K��=����Kı>��s��rYRCh#A����r%�bX(��wٴ�Kı=�{��r%�bX�����r%�bX������p�9��8{��籺�Z�ٍ�u���va{r&�p�V.�5�;v��bX�'��}�ND�,K���ͧ"X�%��~����bX�'�뽻ND�,K����Қ�D��ֵ.�6��bX�'��{�NC�1ș���p�r%�bX�}�߮ӑ,K����i�X�%�}'{{���Ir�u���ͧ"X�%��~��"X�%���nӑ,K����iȖ%�b{�����Kı/g��gMY���al5sFӑ,K,O}��6��bX�'��}�ND�,K���ͧ"X�zA1AX��V�RHb�O�"����{��%h#A�rH�2㈱q]�bX�'��}�ND�,K�0O���ٴ�%�bX�~��ND�,K�g�+���4���~?!30HJ�p�����pX�\��X7r�[H�p藝�v�.#.ֹ[�k���������d�=�siȖ%�b{߻�iȖ%�b{�۱9ı,O���6��bX����ZA/��"d)��q�4�����ND�,K�u�ݧ"X�%����fӑ,K��=�siȟ�dL�bw�w?h���f��]h��ND�,K�o��r%�bX�{��m9ı,Os��6��bX�'���6���h#C�����H��)@Ɏ����`'��}�ND�,K���ͧ"X�%��~��"X��T��s��r%�bX���������,5u�K�M�"X�%��{��ӑ,K�������%�bX�}��ӑ,K����iȖ%�bt�,$
�AH1+�"�H�t�|��98�����M�tv���;p�ƸB{�6�{Xō�ɸԩ�З=�6�tP�G�hu�m۪n�+Fض �+v�v�Z�	�]������k��S���
�
���%Yl�qi�5��ǔMt��[����@ml�ɶu�Ȏ��hzAsJt�K3�};st��^�J*��v�]�l����e����u��Ж��5r����,T4l��H]F�\e�:8j���K��5�^!P�ޮ��]��Ϣ�<�sڊ�a&�����bX�����"X�%���fӑ,K����h��bX�'��{�ND�,K�{�ft�˫���Y�6��bX�'��}�NC�1ș��o��r%�bX�g���ND�,K���6�"�F�4��3�@��I���Ԇӑ,K����iȖ%�b{����r%�bX�����Kı<����4��h{���2�G��$;ND�,K����ӑ,K�����"X�%���fӑ,K,O���7Ch#A�+H%�2�4Z�m9ı,O{���r%�bX�{��m9ı,O���6��bX�'���ͧ"X�%��{�ۭL��5sF�h�YtӁ�s�xܽ"��+���q�vz�����n�����[����Ww�����o'��}�ND�,K﻾ͧ"X�%��{�siȖ%�b{���ӑ,K����;u-�f]Kp�5��ND�,K﻾ͧ!�6��	 x�+@JBDꯠ��8D�%����ӑ,K��߻�iȖ%�by�wٴ�OȎTȖ%?��~4j��Mf�f�6��bX�'��fӑ,K�����"X6%���fӑ,K����iȖ%�b_I���d�R\�]f�kY��Kı=�{�iȖ%�by�wٴ�Kı>����r%�`~X�O��fӑ,KĿ�߱����e�\��Y�6��bX�'��}�ND�,Kʠ�{���6�D�,K����iȖ%�b{߻�iȖ%�b~0��ʊ��7�����)��<V)t{�kZK�K�c��k�U��t��;�(ֹ�+|�D�,K�~���Kı=�~�m9ı,O{�xl?
O"dK�����6��bX�'ߧO�&����Mf��Z��r%�bX��w6��bX�'���6��bX�'��}�ND�,K�g�
HRB�}93ER�vZ.�[�fӑ,K���w�ӑ,K���w�iȖ4�0$�3��������50�"n%�5�J.a��� �bm����̙g���4�si5����aIIxX�s�sS�@d�!�4�x���6�a�36��Z�6�vGFfLm$�q%1C ����! �K7��&'^��d�
� �j[I���VYa@d�Jow�h�"��!tF@��xR5�pf�[�ֶ�I�=��IH��RӇ�
B`�����-#➀sP$��"�վE�pR�0�!HRP�F%��7P�@�H�[l��Y��nh�:���`�*�Hox	�� �1֝�9���)H`�����a�WP��򈇊�H#`&����~v���� �U��X;<@� ���>"E>~��� �Ȟ��]ߓiȖ%�bw>����K�F�p�/�N8�EHp]4���"{��~�ND�,K�~���Kı=�~�m9ı,O{�xm9ı,N���R��eշ%֮ӑ,K����iȖ%�a�`����6�D�,K����iȖ%�by�۴�J~�~�~�z���aLb�69����� M-w6�Etd�am �ǭ]`�r6�Ԛ�h@Y�8ː�4��hk���4K���w�ӑ,K���w�b�bX�'}��6��bX�%�I���)n��p��\ֳiȖ%�bw��i�~P#�2%������9ı,O�~���Kı=�~�m9 lKĽ;��8�(�YN���4��l�nӑ,K���fӑ,K��=����Kı=����Kı<�A�S�ې�`N8���F���{�ͧ"X�%��{�siȖ%�b{߻�iȖ%�ƾ�@$�FC��BV!�E�'����<��s��ND�,K�ώ��2��\q���A�F�����AD�,O{�xm9ı,O=�{v��bX�'��}�ND�,K�ڟ_���٧6��u�6�Ov��/Q�m"�:kk'3�Cm�!�������	����f��f�Ȗ%�b}���m9ı,O>�{v��bX�'��}�ND�,K�����A�F���-��N8�EHz6��bX�'�뽻NEı,O���6��bX�'���ͧ"X�%��~��"~ 2�D�??��?f���˫nK�]�"X�%�߿o��r%�bX��w6��`(ؖ'���6��bX�'�뽻ND�,K�=�Y�I�D�5n���SiȖ%��dO���ͧ"X�%�����iȖ%�by��۴�K���QS"~��?M�"X�%�~�~�]RSE˅�j�Zͧ"X�%��~��"X�%��>��]��,K��߷�m9ı,OsﻛND�,K��A0M4 &�ja�
cD �n��%�{��w&l8{3�g�'�DD8,��X�9y�5�`<;-�J)m�F��\�S��\�8f3Oc���*vr[����	�x1[c�m�����K6ڥ���j�������[�շY�%�ʜ	ey:P6:�s����\96�b�6T0r!,�:n溱����h����&75��1��pd�
I�[J�����ҳo]=��V�'kV]a�LֵsD��: �^�a�k��gS���\�1ڴ�3�	wWL�E�)��)̉�v��o�{���g�����c��O�X�%��u�nӑ,K����iȖ%�b{����~y"X�'߻��ӑ,K���GYs�˙u��M5��ND�,K�{�ͧ"X�%��{�siȖ%�b{߻�iȖ%�by�۴�O�@ș�����0�[���.8��a��h#C�w�m9ı,O{�xm9��!��=�_�]�"X�%�߿o��r%�b#C��m2��H`.CJGt0�F�!A�=����Kı<�]��r%�bX�{��m9ı,Os߻�ND��F���-��r(�EHp]4�ı<�]��r%�bX{��m9ı,Os߻�ND�,K���ND#A���dlBHII!Sd��`��r�TQQjz�2�H����ƌ�+�{�g�f�5�\,�Z�ND�,K�{�ͧ"X�%��{�siȖ%�b{߻�a��DȖ%������9ı,J~>���	�щHʐ�4��hk��6��F{hB;�a �-!��ƃC$��VEZJ�\X�n�KD���YJd^��"dK����"X�%���nӑ,K����iȖ"4������(FYaG��4�ı=����Kı<�]��r%�ؖ'��}�ND�,K����ӑ,KĽ���Iu�u,�sFӑ,K?
2'�o���Kı;����ND�,K���ͧ"X�	b{߻�h�A�F�񃨧�I����q]�bX�'��}�ND�,K�_~��O"X�%������Kı=�]��r%�bX�g~̝�R�YL���s9��z�`��B(������v��[�`A�NB�Hn��F�45�{�ND�,K���ND�,K�u�ݣȖ%�b}߷ٴ�Kı>��n�t֦����5�ND�,K���ND�,K�u�ݧ"X�%��u�ݧ"X�%��{��ӑKı;OYD��FJ*@���a��h#C�u�ݧ"X�%��u�ݧ"X�p���"@�>e�J ���g��m9ı,N����r%�bX�{����nk2�ۅ��WiȖ%�b}�w�iȖ%�b{�����Kı>�{�iȖ%��Y�>��]�"��h!�w��L��JF���aKı=�{��r%�bX~#�߿xm<�bX�'�k���Kı>�۴�Kı<�֖ܷ,���w5�T1{Pvz�k,M[�:ⶻ8��g����I��5���ڏ�ز9�ag�w�{��7��;���ND�,K�u�ݧ"X�%��u�ݧ"X�%��{��ӑ,KĽ�}�Β�R���e�ND�,K�u�ݧ %�b}�w�iȖ%�b{�����Kı>�{�iȖ%�b4tE��m����a��h#G��{v��bX�'��{�ND�,K���6��bX�'�뽻ND�,K�V@���!�)��a��h#G��{�ND�,K���6��bX�'�뽻ND�,/�N�,"Ye�S.
j���i��nb!w�[+k��U>Ȝ��9v��bX�'�{f�K�Mjh�k)��iȖ%�b}���ND�,K�{�ͧ"X�%��u�ݧ"X�%��{��ӑ,K���)�g�̾��In�����c���㒹��Ɩ�"!�Xӗ��v��g�9�^4�f�te�Z.�\O"X�%��߷�m9ı,O����9ı,Os��6�y"X�'~�ͧ"X�%�������E��IR+���4���}�Rı,Os��6��bX�'��y��Kı=�]��r$� \�H��>��)PT�USUp�P�Br���B
D���n	"~���nӑ,K����nӑ,K��	;�۫%�˓����m9ı,O���iȖ%�b{�۴�Kı>�۴�K��=�{��r%�bX��ﱝԗZ�V��.kiȖ%�b{�۴�Kı>�۴�Kı=�{��r%�bX�w��ӑ,K��B�KA>�����8���	�:��4�>�U�N)��R�����z�ѵ��/�l��'����l3מ|�|-��tm�,��zH��g	��-��z�6ָV
xq�K=��j)9�Smv�UL��q���;l�ݽtW`i�k�7d;n�+܇����L�:�O:곸7e��E�[s�*�.��)5�t�۵k$ג�^j�dM���Y�I�����w��;����֩6:)\��[�#3��V@8�X��&��V�}�����u�~r�j����}ı,N����9ı,Os��6��bX�'��xm9ı,Ov}�h#A�ߏ� M�B���f�ӑ,K��=�siȖ%�b}���ӑ,K���w�iȖ%�b}�w�iȟ���,N�~7r_�&�4Mh�e���r%�bX�����"X�%���nӑ,,2&D��~�v��bX�'���ٴ�Kı>�}����5�tK.�]f��"X�~D����v��bX�'k���Kı=�{��r%�bX�w���Kı:vk���K��]YrIu���Kı>�۴�Kı=�{��r%�bX�w���Kı=�]��r%�bX����ݷ���L��j��^x�G7c��	�Z�bVA��:���:z����9��#�k���ND�,K���ͧ"X�%��{�ND�,K�u�ݧ"X�%��uߕ��A�F��O|�q�i�q<�m9ı,O����r��
ix�9"X�s]��9ı,O{���9ı,Os��6��bX�%���}	r	[p]4��hnϾ�ND�,K�뽻ND��"C"dO��߳iȖ%�bw���6��bX�P��u�E�$rR���4�ED����v��bX�'���ٴ�Kı>�{�iȖ%�b{�۴�K��ߏ�"i�Cp���t0�F�)b{�����Kİ�;�����,K�����6��bX�'��{v��bX�'�{�߳���u��&��r��q��4�����'�igWE�N�2���yx
��sJfkD�MZ2nk8�D�,K��~��Kı=�]��r%�bX�w]��r%�bX���m9ı,O��Y���FJ*@���a��h#Cw���rbX�'��{v��bX�'��{�ND�,K���6��bX�'N���)�e2Lp�4��hwӽ�ND�,K���ͧ"X����F� R�[�$�����S@m�`;63A�1T@�>���=�����"X�%�￷�m9ı,JyӸw$�Re�Yu��֮ӑ,K?"}��~ͧ"X�%��߿p�r%�bX�����9ı,G��9�
HRB����Z&ʚ)M段��r%�bX�w���Kİ��W�����%�bX���߮ӑ,K��>����Kı=3����	�i�r�`�u�U���{'S����vd�7�c����O�f�2�}��oq��Kϵ�ݧ"X�%��u�ݧ"X�%��}�sb"X�%��{�ND��F����[�4��`M�n��bX�w]��r��DȖ'���ͧ"X�%��߿p�r%�bX�}�xm9���2%������\�����]k3WiȖ%�b{����r%�bX�w���K���ٴ�Kı>�۴�Kı<���33�f������fӑ,K�����"X�%���w�ӑ,K����nӑ,K�]ܐ�O�5`�"l���4��hh߬��Iȣ%!u�6��bX�'���ND�,K�뽻ND�,K����ӑ,K�����"X�%��|}���e֡rK��k
�}����Z�Xx��������tɆ��6ۋ�$�p�N�]�������d���nӑ,K��>����Kı>�{�`��bX�'�}�ND�,K�t��0ԙm�]k.����Kı<Ͼ�m9ı,O����r%�bX�}�xm9ı,O����9ı<�N�Κ&�˓��ֵ�ND�,K���6��bX�'�}�ND���2&D��~�v��bX�'���ͧ"X�%�{>��MkV���ffh�r%�g�D�����Kı;�_�]�"X�%��}�siȖ%���N����iȖ%�bz}��̿����֦���M�"X�%��u�ݧ"X�%��}�siȖ%�b}���ӑ,K���ٴ�Kı0�!�;�:|� ������>\gL���!W����sd���[��<��-kA$7���:���Hm�A�G.陠�3Wj�CSp���jSL"��P�we�*��[V/�,�u���ָl��jR%���B��l�=�D5��'(g�����/��$��uc����ǉ���(��
���&of:�Z�4�7��T��=�d��_W��6GDf��=�Y\�����#�7�.l�I�"�1�H0�C����xBq9.l���$4y��TM+�I'����<��r���p��1bJp�`P�����B�m9�B�̢(�{�D��H$�2Y!�#FK�V,s��E�������ܑ���nu���Z�h�1�z�Ձ�r����ڜk�j�J�V�J�nw��ۧ�7E��Kd�F\;��N�.IGs���2Bk`]O<�J��7tu����� -M�9��S����\��i�dMɘ:�����u�����cI���7]hz}g*�*�v�Ri��2^��8d�&�J�T��7Y6S��⮁TZi:��g��t�}Q�5�sM۴��E�\�� !B�=��pgmM������랮�q���%rJȹ��A��61؍+�S�'�v{s�m��=jU��6�q�n:�{��6�*�"�ۢ2&{pnG�<[��yvt]�v��V�*63t.x�e�(�e�`�-�;`��=�,�d1*�n˴��񒧆����Li�um��wOh$kjVuī��ךک`RZ�!�y0l9�yѠw*֬�R��*�R�PUދ��ڕݳ�̛@1�����J���am��^�6U�R!{$H����y٩۶�$&��ݽ[cT9u���aieMMU��6Ȝ K�pX��;^����m�ǭ���n7 �Ӓ5��TG,�m���n�����:Y�&���TT��%���[�����O;v���ت�j� ��[�k$LM�d����8�vqξ��g*�.��3�U�UҮ�tE��wiwv(�� -'6���vX�#^���⸘�nʩ���vm�[͌Oeۊ+��+�s�5+X�;lD*�sf�An�=��ў���M�q;Gj������Y)�ge��]�]';���Ɩsp�OH
q��)r˻2��U#���˺A�(�2�c��Q��uHh7;lI��O[f���F(z1��[��;u�%��d�H2�[t�&gGZ�!!�U�˛��j�\�0�6&�㇇)��Y�.m�[ٻF�KM4��RƊ�Ԟ��x��)qu	;Mi�qn�<����ڬ\P��b�Z�Y������w{���^/��M�"�(x��G�4��O@] ��z�:*���0	���"�C�Zx���D��>Ge��J\�7PF����<e��vҭ<��6!���T�,n��:nal�����/g��k��5�����|#T�΍��i�W�k���1�1A�:)�H�u=�S�0�Jf�r(+�3Z�ŷt�w:�H��Tq�\a�Wp�ݞB����[�)��)ӵ���������w�1��j�tn4�a��2P사1!0a0�`����U.ݔ$$�:Gm��\�gkӄ�4��D�۪b��m��v�.c<����lV���w�%�bX�g��m9ı,O����r%�bX�}��6�Ȗ%�b}�w�i��4��p�းYG�Ȗ%�bw���"X�%���o�iȖ%�bw��nӑ,Kľ}�u�aH�F�48oY��FJ*Dc�ӑ,K��߷ٴ�Kı;�w�iȖ?��Dȗ߻�[ND�,K��߸m9ı,N�MN�4R�Z��K�e�M�"X�%��뽻ND�,K����ӑ,K��{�ND�,�<���m9ı,Jy��:a����]kWZ��r%�bX��~�bX������O"X�%������Kı>�۴�Kı? �����m�8�BGOl���dH�"roG������nS߯tv�|o��<�<N��O"X�%��߿p�r%�bX�����9ı,O����?
��&D�,K�~�ӑ,KĿ�{��I�j��al�Y�6��bX�'��{v��@ =G�`����܉Ȗ'|�yv��bX�%���[ND�,K���6��#A��zz�c��-�",���Bı,O����9ı,K�{�m9ı,O����r%�bX�w]��r"4������&�$7qH�WCı/��u��Kı>�{�iȖ%�b}�w�iȖ%�X�w]��r8�؏؏�}��m��9��0qɿ���ذ�������uwN kn����?
�=����uU�j�M��##��s6�]��tI�ǳkv����}X�@�;��uk�w��Ӏ7M� kn����C��nh�3�s�F� �Z�ՠ�4m��-v��ă9s��I��QI�h��M�w4������`AX�0���@���)q�CJ  �>���'���-�TX�7�d�M������{�,��� n���K��ﾼ ����$�8���nf���Z�ՠ���w4-��M&��氘�4W�r�>�w�E��o)�KQ�	yy�nwncj�ߞ�}�Ǜ�
9	��/������٠[n���/�����lM9�7⑸�[w��Q'wv,�wN �79���H��P6ױG0�f94{���5�s�Ц{��p�u��Z��3W`�"#��v�V�k�hm�@�%@~��Ͼ��>>�=�4�D��L��Z�ՠ���w4]�@���C"�F �d��1`^v�Q	�n�Av4�권�ǩgvP���st��2$�RE$Zm�@����j�-v� �r�� Q��bRI&��x�t���s�ۼ f�C��$�bB���k�h�V����$_{�@�����\;�o.7܄�G' n�� ��������N�y��NcX�$R7�v�4f{������8t��"!�s�R��U�w/nӔ��och�\˴^��nzΡ�l�K�v�<�&�n���t�c+kz�$��kלV�t�닞nG���y�c���ugq�ضٖ��8%�D�$�M̄��s���6�e�ez�[GFĘ;���Ce���m��Nu!�m6[DV�5�Wql<�^�N9N�ׂ]�r�= <\�����!�u���ѳ�	�#v��Q�E[�+M��v��{�O��w���u���4w^���m"8w,Ň���6��ۄ�Ǯ\�9�s1�8�������Z�ՠ�����T�9`�"#��k�� n�� �����>�
������EfG"�=��- �h۹�v�V�gxWX�Ʉ�$RE����w4�j�-v� ��*��F�ŉI$���h�ՠ7M� kn��	)Lit̪���Epc���Ŧ�ms��p�p�"X;QEt�/<{Hq2�(�HD�oM����-�j��f�m��ظw��V8&�03VI�t�~B�ꁠ�HP�HȄ�#F6 �)H�		zb�P�����m��5�s�{�r�ؚs�2H���l�/{w0��U�W�N���0thE4]Z*c0qɠ^��h�ՠ^YM �hξ�I���f���ZGog�w^ �^,u[As7r�w/�<��X��s����|�n^�FN�OR�FC����F�pJF�ؚ��Z���f�{۹�v�V�gs��&�bP�
C@;m��n���Z���ʲ�,Q��bRI&�{۹�{�}�����r�BR��&HCa!�t+"�)@�G�RB����U����x �:�aws5sD�75V�>�}}Ӏv��ۼ����\;�o+pm�Ldqh�S@5�x�x�t���v�t�B�	9қ\�o�8���7pQ���@�h좽x�ƻn��C���4�5�d�G$> ����{۹�v�V�ye4�t�p�`�P�����ōr�:{����� 7�s��bG3���y$@�"#��_��-��hm�@����.u�^DIT]Q5*��p:S��� >��7'��0~B**�5�r�Is��y$�)p��f��۹�v�V��YM���3A3���sc쎯	zn3���^�ԛf�닫d�SM�rY;v��X�����6AbQ5��I:����s@�M��v��%��׀oTu���q�HDnf���Zye4�٠r��o�bG1v��ͨ�rZ޾0[w�y�ŀk�� �58ˑ��d�$Prf��bW���9�{s@�v��m�٠_2����s1�8��?6�`��7u��m��(_��.�� F"�pq�2q�e��˗v����=��8,J���ˢ�ݮ�I؞n�N�'6݉��9nP�X1�Z�z"���#ճ�z�n��h��p$��ݖu��3\�O5tm�m�&�/Y9�mF�t�~/�}/Y�س�g^��<vt�p:@�E����j�a�x��4lF��x;GZ��g�:�I�����秊�3l7�`<��f����R�kZ�Ԏ �C��P��5X�.����kۅ��܁�Xp�FH����x�{Ycl���kx-�37j��x�]Ӏn�ŀۿ�D�>}� �:����ʫU$ԫ����ŀl�� ~o�]�>J�&����7$�)$�4�|��w4�fc��� ��� y\�V�M��)S5wwX��`��`[ŀl��^��DG�x��h[)�g�f{＼OwՀ=o��$%J˫�Z�ݗ��;V�t�L��5tm�]���m�y=lp�"h�����r�4�w4�������e4����K$5�]MkF��}�7��� ���A"*�`�����Pؾ�'��D׳;�74z��z�`�M��cQǠ^۹�}l��{n���פ�=�I�"%�#1�d�����������ذ��X��`6���c�H����{n���נ^ۋ �ݳ �[��gR�Sj��n��s�lZ�������*i�8t�Ύݻxm��ٙ�HǨM��,�I$���=�x���0���B�)թSu-�Ĝ�=����e4�w4�������x����8�$A9�=�� ��XR����"*Z[?�DUT(� �̸��c U����(H[Wa�,�
�'�1��6��F��u��,pZ�#58��t��[~��<Z8HD�FYgRbHCЉ�>joNh�$h��kGƢq�%0�ZM	���'ǖ$A�E&�,<*��\3��i�/����$峅#|������V@$d1�0�H��H��"s��f)VBh�:�$�d���x �P6+���Q�B�H�y�����QF!���.0cI�	�CpwhS�Q�A�^*l]���l�E�D  �V z��=A(|� S�j��ھ
�U=N�~����'��w4�s�ƞT�I�	���{n��X��`tD�_t��9usW�d�$Xܙ�Umzݷs@�ڴ�ڴ쯾~��#0�1�1F&q��=t�ť�㣠��:m�u�������ۋ[���Hc1�����s@�ڴ�<����ﾬ�?r>.f���T��V��\������ ��Հy�ŀ_�j�iĜI5��;�j�*���w�b�;�����f���Z)7737s��)��Հo>ŀ7Z� Z�@j��b���D�X-Hz*��P	n�۹$�;=�sE.�fL���`z�`	B�����8����r��\f4B5���RH�v���stӡ�ԯ9W�q�b];[`��>���Ĉ'3�=�|���ZW���n��.u�ˉ��!?9"�>�o�����V��,��9ВIL��-�'1���nE�yz���n朒��_S��<�pt1C���s��M����;_j�>�hol�;��
D�Ȧ)����������׀{u����B�R1�iA�Aa!D��^�����_��m��YwF��S������$�䴎���zu�qܼ[[�s�v���R�nL��s]�^��n��ŧ@��� �<=���s�e�-ءm\m�v�K�Tl��nm�Z	ʝY�ix�i)�t�ӳ�:!���jz��eN+[�\�;l�ig3^%��nո#v��yU5�ݱ	��a;fi�d�t&vN�K�q#��1֤���\�`��HK���{���������}�+s�Vm����..f�u��ۋY�t�,�g8�n/�8)���Tr���4w�s@�}�@3��ctj(<�
8h^��=��`ֹ�?k�`��N�,Q��bJI����h�ՠ}�)�U{^�p���R&��"	����Q=��p>�0/]`�x���&4�	�#r$Zݲ�W���n�k�ZUv���8�Ls�8�Yܾ�]�vm�F�t���]wD�g+��N��GRcY&9܋@��������sВ_�<���Q�*�Ue�N��˚��{��7�%��(���ڴ�e4��q^�H���#1�d�缬��Ӎ���	��X�ۚ�_]q(��Mdn-g�S��� =}x�^,�s���Cy\Q��
8hy�4w�s@��ՠ}�)�s�k�m%7�rBG���[�y�ә�DƤ졆ގwi.o]��r�;�ne��X��ǉHܚ;۹�}_j�>�l�
"����7�:nI���T�K&�`�k�脒��ϯ� z��w�s}�����j1���F�&2H�>�0}����BF@��J�AB t8 y��ٹ';�v�{ہ�8��!$���f~įo���}��}_j�/,���i��q�Lĭ94��������h�l�=����ƣ���6��I�9����']��Fqٮ��Œ�4���:�\�'gF�S"x4�ds>�w�@����v���s@���%�H��F��/,fr�Q2_^��,���t(��^��7�qF �Q�@=��^��h��h�S@.ڲ��,Mɪ���P�{���;i���ـ�,��x�d �('�P(mM:3M�@4h�v�!�
� 0M���ߦ�p�_���<H�������g�;_^��, M誥^���=���yU��hN��3Z��Y�j0����n�ȴriVv��h����&�`���<�ŀ?V�����w�Y#$$�y�4�w4�ڴ�)�Ui�ƮLĬ94����\��)�}|`k��<���Ŋ9�����L�/j�/l��?k���y�~XGS뫢n���\�YUs�=v������}ذ��8� �I" �BA����S�N4v�x^ְ���\P��v_m��{�1M&�]���J�Pn� �n��G�wcۈy�O]�ձ�RCb���O���f��6������<�*vE�S\�m6�:e.^k[b�������k��y�Qӆ55�nB3C���4�3�Y���s��Bּ��b�K�^o29���[���F<�[��<�mm�D��u�BY��J����~{���]�-Ӎ��ۋ��`ֆ�cJy���N=J^G���]9zbv;CD�����������`ծ~I$��!ϯ� �'ҽ�@B��Mɠ^۹����#�w�@�����@)��X48��Č��`ծp�l��w�y�� ��q;�fHԄ��@�l��^v���������H��QI.� ~�x�x���8�`vA�덵\�l�#�6�;�^ �50��gY/-�cz9F�����%�\�;�94[w4�ڴ��h�l�9��ODp&
*@���=缯��UH������ =����,�J"d��w��b��M���}<h�l����}�nh�Z����qF���� ����,���СK}�h���S(	!7rh��hծp�l��w�tB�[�GL�ԣ�tW-¤��35f��.�����:��87Cu��rqu������}l�	g�4�~��:� �v� ~�~_��V�uIR�	���	����>��s�@����/j�~�ċ}�RB	d�(�������a��R��""RBS
*A�Ҁ�}��=�l��u0x�Ȝ��$�/{w4q����0>I(��(UZ�����}r��ɤI7r]Z�=��8Зog�=�נ^��h\;.$�R,f"94�x�.2X�GHr�<;WFN�Oh.�;9k�-4Rd�F�Z���l�/{w4q�� ϻ��ydQ9p��n��S'7ذ�}8�g�(�2�/�zcX@I���@�}���}�@�즀}�f�S���hq5�M�V�>��}87|`�7x$���	�|��v��׆�^�Y����$'�Z�e4��h��h�h\�ex,�D���	�i��lI�t��$�˒�r���z��]�Z�wh�B	d�(���[4�w4q�<���C��0S�E*�VU�V�A2M����}�@�즀}�f��\�:��	��"JL�9�ڴ�)�r٠^۹�s�� ��$ț��h�S@��@��s@��@3��q�d���h�h��h�78�l�<�DL!��ʋ�%�[�#�-������}��70�t)YQ����9@��҈��`�?jSIЙ�p6\1���F���`��D�n��׊�y�������9��	�z�e7OD7H�)��^mk행ŰI�!q3A��jk|��3��{�p�y��L{�!bCm�/9���״P��Mnl��Wm)�n��ZA �V
	B���g�=KgM!�5�Hzcqf�Y������Ӄ��C�C^P�{O�|��C������izb�T�*ł�By�\O��uc���Ghl#�|��)�|�x��Hk���+>�H�	M�B&j��k�8gp=�c�7��������3ﻷf����x���X
���i�v��5a�ۻm-�0�۲����;;�g`�m���M��\��ܻj����k�K�ۃ f{2�v�]v��ƛK���lO��s֞�k8���Xz�-K�S�Hű8�ޗWu�'��P���n��u����=���2}��:}`.��Q��ù�7o�]e�q���W��rp�=kz��n��ScFg��\C�s�1u�JJ"���܌S���e�v�]��Zkl��,bX:�ty�WG/���o,u�	��mv��x�l�2�;'b�qZ.��]�i��f��$��"D�"8���4[�N�m3�I;v��F9ӎ�]��;C����q{vB�]+7t�ֶ�h�[��a�����[w˝��1�>�
[��(�v�7k'h�v����6W��g�k�v۲te��pd5*ݓ���k��b#�Q-��NNr��[f�rr��C�^hj�U�Z�k��9�}iW�Y�9áE�c�U�V��j�.UQW��ڕ���9����.�lݶj�(�M	9��K����α�ӗ2 �peuf�)�����&�#�sbRW9�[�Ħwj������ݜ�y��rx�<��2U?\��ii��-��o$���Gmù��㠳{;)�Ep��@�7.�l�[֧�l�g����m���b+G�V�.�Α�m ���6���O; �\�dޖ�ɵU�T�f�^[lJ���g�f�g����c�h�;�!)��+mb������vت4�@mgeڧN�5Yj��UT1�}��g8���]��*K4�a��Nb%������kB�7K����Zګ�Keh;
�4.2 �v��������.1����qUm8�qۅ�h��P��7Vx][����5n&����Eof�:�A.�cm��;l͈ՠ��%����/5�qg�
G����m�Z�ȤlF�-���k�KY��
�lR��wY��z��v�@�d�8{J���#�<q٭��ak2�Rf��jkZ�fj ��xz��@@���|� u"�
����Q��D�R"����@O=T �����՜;����tk�:�Hۓ�:�:�w���&Ҙyx��i��]�K��m��0#-с����b����t=k�ڕ���1\v]=p�n��8l�%�;d�m+q��[<O�z�)KU��Z�^m5����n,~u?'5R�s;��P�ai���W(k����n#N�Փ=c�6��.ofz��Su�$���tm��N���8�)#N�
UU�BL(��S��]�I�v��=M§X�K��wLu���KM�u<��J�2�a����Hm�q|{�nh�h�S@��@)ο���,Q�3@�j�/l����@/m���"�\C~�l�2Bc$�@��� ���8tDDL��� ����=��5L��Y#�(䆁��k��f��j�/l���V���D��F�
]`�� �m���s�� �>�X�����t܇Զ�c�����][l%��M)V�u��ñ��΋v]��]em�4��V�{e4�;^�^�4~V�&Fܘ�D�F��/l��E��2��F��&��x���Հ�u��Z�9%	L�mO*����4rF�qv���@���h�S@:T�0aaZSϺ�m>��`r�
}Z���_�B!��`�c�=�>ՠw���>��Z���������&�9�u^N�՜�;^$�M۠f�l�:�3Ѹ�ɀ����)�d��I��vS@���Y';g����}�Oo��iA�!.�nn���?z��rP��=���=��h�e7߳�䋋���"ps#_���I�{���9�{��� v*R,R
� }� ��s�޵ٹ'�����qs�T�L���q�$Z�}�@�{)�|���
��@��k�dmɎdM�n-�)�{3����<��=�>զ߯����9���K���6-v;t6i1\���Dz����a�F���n�yx甥n �ؤ4��Vנ}�j�-����Y�X��'&�k�o����]Ӏwu�zOk� c����R'#�9"�>�h�M��l�-v��ۈn!Lx�$��"���vq�l������D�@$Dʡ��0�ik�����|P�7�)�s�SR��GR7����W��r�h�ՠU��Ĭ^�g4�)�<v�륞9���c��if�6�:���K�5���v˫Ef�8����{^��YM�ڴ��@�s�T�L���q��z9e7���~ďy�- �Ozh^נs��2A8��7v`ֹ���9(�=<��޾4;�Yq�bn1!�����[4
���r�hs��*e�0����!ɠ^�ՠs�S@>�� �9l�9�Y�_�/�4��&dL*
GR����|���V�œY��P,i���ڟ+�=E"�q�#9���V�3�\���eF�-���jt&�I����g���q�A�Qƶs�T)������ەk���Cv{�F�mõ!uל%�ݶ��Hz�ݐ��,��S�S����+��Y�m�cr,m�]��4D�&�I�ͭ��[#��I5�|���m��z������G�0R�h�^f���e���4&k�*��n�ルaݎ�(��u��A�ѳ�<��kl`�BH�q8�������� ��4��@�_j�9]���%18ړrTݘ��y�J�-������3?${�^5)��K$qD8��-�e�X��� ���O��q�dk�I�u[^��vS@5�x��O� �k�>wd�$������e4�٠g-�U��r��6���q��9{f�pu�'W<���t��%.;8�f�s{WYnѸ9 �h��f��mz9�M ��\o�$� ���r٫�C�	T�i��=�`�� qS,��,m��@궽��%2>� �����;�����ǉI��vS@;m��r٠u[^����9�&��&�!����!O��_��u`��0����=m�@�k)�Tp�`�ml�B�n�1r���r����Z[\��2�c��������m��H�׀r��c~��!̍`�I4�ڴs���l�����̬�<��.�p{m����С5$(����A��L$ؼM��=T5���y���j�9�w�Ɋ�Lpr�]���� ݦ��!$��� �Q�����Ib�Ȝ���l�/]�@�����f��r׸�Jn4��*݉���e��\��Õln�\޴>��E'��C$��LB��A�4�)�}��h�����8�}4ǖx�'��.n�p۶�䒉���x��^z�Z+����R(�
C@/m��w�h�ՠ}��h�]H�(��]��wuw��	%3��^λ�rN{�� Aր�Q<Qt�)���������8�25��$�/]�@����[f�~[�����Z�Se\�mM\��&{���z9%m��%��n��.�Wcn^����={y�Ӻ�Rb�E��x�[f��;�4�ڴgG�\DQ�Lx���y�x�n��7i��?n�3�$�C�Oh~q%4�#�@�-��;�yY'7g$�wt�N/���% [�7&���M��S@9m��ً���@)�="I��ǉ9��Sd���I�wzY'w�$�ʺ� BH�D� 2I E$+�>����.�<������:�v]���s��qۮ��ع��04�b[cwt<S���<�Kv��xvMc�R��-���W8녷���x9����[�0�v2�)
�U۴��i���@��s秣�'s��qt�b��uKknݸz�����8�U�B�y������gtl�6�3!*�%G7[�į�I#�;�kړ�l��ɴ��s��������8��s�f\̒��WY�Mj:�*�<Pn���#n�ZV��M�m�$M��#lv�s��HȢ`�N{勒NޖI��Ɓ�{)�^Uu"b�0K$q�&�~[���l�?n�0ͻ�<�ND۹#�r5��$�;�)�}��h-�@>����̬�<����vـm� ~[��>Q-�q�j���"9 ��RC@9m��w�`�ـ~ݶ`��2�h��.e�6��5q�@C֫N��k�����;Z1����$z��q��oN��3��9�Λ$瞘I9���8�
:G@]@�-��5��=��}7�OA "(�<��<�/�M�����Ny���8��K�����!��I8�a����d�oO��Nn��N#��d���I�v�Ɋ`�q(Ƥ4����f��?n�X�D��q�>�$�tZ%d�"8��:���@����ײ���,���S�H�UL'@�A�;� suͥ�x.��.{\�Sz9�ױ����B�i��sw�Y';g$���d�\�נ|���A�'���s4�e4�sw��uxo;$��X�N˜�8�p�.Cd���,���y��P�hf��x��0��q9��E9���)��IL<�3p5�L6��
�!DT ������3.����H��3.���
&�q�	�6,C�N�<��*k���:X	�C^�`�ȁ�i.I��&BDʆ!� U�O0f�%)L!M�y��Ҋf(툛��f�l�y|7e4b�Ԧ�I���4�}���"����f~5��}@Ѱ�hFʑ�,D�I��K�1��}#�R��hQ�@ ��aX8p�b�֪�.̈L6G�x |��!$%}�
��d'�v�K;}�%���S��L�2��ن��h֪X� �! H�ؐaH�`C��#n�\�c�͠J.���@1L# ���7���ЈF�ը�J5B�4��ɤ�CѵGh�8J[n��5�~��x{��*�}�f��6*��>ڡ ڔ`iBʈʺGb&����!���Oj�!P�E_E� ������̀+�'��zg��{7$��h�(6��F�ē�rhyWܾ���,��fDD$�|�^ {���K����'7zŒs�q�I�ޖI���p� N��/��($�Tԩb�epW)]�su��t7^ގ׫��Ӣ�HN<x/�9�ײ��{f���:脒�!�� �>����EM�F2Ԇ�'7zY'W��Nn��$�l��31"��zb�L�%�H�qɠU�:�ۯ�m��u� שȪ��!��Ɯ#�>�n���M ���ܚ�z�1����E�3�e��E]�$�J kB��a�
D�E95�g��%^γ(I�<�������M ��� �z�`�m�DB�Gg)%]Uܪ��l�<Ol��:��nml���\7�+�Gk��k��nL��9q<s�$> 徘��� ��l�I~�|� ��k�G���oaV�?g�[<`���]�)��)��]E��R�P�@�Ɓ��M ���@��*�6S��aur��R&.n�IBR���}4�­��S@�_n!�
cJF�Ƥ4�����*�>�n��=��}7$�x1`�!FJ�������G\�0qr��7=����웃�n��n�v��[;�"v�Kyݭ���KR��g[��ƹ�6KLv|�:�<���q���]�-ݭ���ʝ��kg��1�X.��!�FmF0ܝ�0�=fz��Ƕx�u�=
&$�N�t����L���ΞW�7g�g�ۈ��Nܓ��͔���۳v�����ݱ;5��{#��w�NM4NN[���������w�����.��'��u��m��荳�f�4n(�<٣�u�:NB6N�X�oc�I�����'7zŒw�q�I�ޖI��_ͻ�8��3�@����m��ۮ�����(S'�WQ�ujiSUq7V��0����N�י�s���i��,rC@>��@����;�����h�YA�dR14bp�M���@�;w4�)�^٠w�ԱL��ݙ�͒$!�k���u��m�Ճ&.�]�St�wkC�j8���wV��LknG��ۚ���l�/_h���)`G8��	��-�_M�_VHċ�"'��A#*�J���*��M*�f�ɠ^vT��s@�n!̘�4�h��!�^٠[�R�;����)�[k�#&)DqɠZ�E�w����S@��@�w���s$d��1� �^���)�v٠Z�E�f~��u{=Ɩ&�MI"v}�-r��Y�Z�3�"j	�{;��ú,����A<#M�Ds>���^٠Z�E�w���;��F�H	d�����N�׋ m�0})�jȤbx��$�oi4�sN{ �v�P4v �UP��Q`  ^�z|l�s���I�	#�%�	cnI!4�s@��h׶h���:����X�ǋI��-��O��� �|^�׋ ����h)�3�Y�Zy��s$�Nl�(����z4�Nn�3���`-��닐�Ӓ��m�� ׬�}���07.�W�?)JE$���h����S@/;f�ޝ�4�HɎA��@����-��y�4��4�3�����71��-��y�4���[��� B0 �R@Ta@!�E� "�׿of䝸��pY %�Hh�l�<������,�78(���8�76����]��-��ݔ.�GL���I���ƍ���2 �j2��Hh�I���x��X�nz"� v�� ��������6�r)�^v�h�ՠ��@/;T�fg�,<x���<H�j�λ� ��
d�����-�졒D��ԑ�8��h�e���`i��<ܺ�Z�V2(��I����/;w4�j��~���S ��IG!C3��r���u�+ɵW�;��.���x6��x��l:��Av�eݮ���k/<t�=�m;)�#'
j&!�����)�#�nW�\�l^�n-��P���f7n�u�c���A�i�w�}�:�ZV�s��Ʈ�Z���vv�k����a:U3�h��ֈ��8ur��z�1�Gb��˸��ʚ�0y+�@�:�t�=O%����Y;��c�r�V��������� m���D�Z�h��kZ5�������l֬/��Rn���������{f�88�W��1�q�����s@�v� ��{�M���(I��71ŀ=�� �� =�^ ���@�D����Zy�4����n�z�Z�.�q���hh�I���h����h�l���ʢ��܎E4�����8 ����\��D%��e�rT���κA&�Gi��:N��l�n�N���x�=Qc�8����u�i�g�8�����~?� �� ����!�� ����i��"j8��k�~fc�3	�X��9�M"��R475N$���o�v��z����h�W�Ls ~R(��I�9�e`��`]� ���5K�ndx�8�5$�yn�{e4��hw�z��J@O	�B�X�l��� s����ŀ~�����]Hg,su���ø7DF�q׎�\W��t�́Jl��6�v�M�V��$4��hw�z廚���tˌm�cX9�@����/-��/l��^�� ��eDʚ���+ ~o ��0=B @��&�!�! J��&g�krO�{G�U�)`G8��D��^�� {��;����X�m�]���ԓҐ��٠U�����h�S@�f{�{�d�q� ��Lvi�k۬��Jv=stt�!׊a���1�l1�@��DR''�y[����h�S@/{f�Ν�̏�Ƥ�`����f =�x��V yoJ����9)3@���{�4
��=�����v�$mAHc�f(��L�}xK|V ��,	�	�7�3#R��-"c�cʱ�BЕ�p0�R�e*�C?_���_8hx�Pcițf�94;����X�l��� ��󿿟��dV�n9�v�Ol[��l,���2W\��7u<h��k̓[�[rr�]ݕ���X�l���G���=�=8��Ŋ&�h�վH=��sο=����졑H�Ƥ����4��hW�^������f���^�!��""�94=�3'�n��s�X ����]��U�i̓$cqǠ}{w4��������}�sRM��g��'�QQW�������QQW��EEZ�**��QQW������U� �� AH
�U *@����A * ��E`*H���� * �H����B�
��"Ȃ"Ȋ�X
�
� ��D"�
�U��A`*b* *��F�"�  *",���H
���B����"����F� *",��AB��T��AA"��D
�@
�Ub�� ��D *"��
�
� ����F(� ���"� ����D�"�`*(���E ����E�"���,T��DR�b��R��"�`*"�� �� !E�ꨨ��¢���Uz�**�QQW�����UEE_��**��QQW�
��������ਨ����e5�-���g�� �s2}p��J���E�R�	 �B� PP D(""���R�E@"�R����R��B�%E$$�$@J�@(( H�DPUEJAAE)$����R"QUp     ` d  
  P� ��3݃�݇'UӗJ=� 7B�y�W�q�c��4;����-�w�nB� �>�/y4� =���3o���wO�8ϒ����j���;ٹ��h������\]iĪ� � (� *�`Ob�e��4�aU�C���1���*�n�e�����/��jU`�)e��������B��^ZW{�ɥ^�
<�F1�;^�c*ũ\� {�����W��ˈkӝ�W�� ��)@ T�F���M�uT��C�ͽ�t, t9ҙo��,>��������"��;Ҧ�{�W�.  .#.�w�J=�}�(͟��u�ͩ\�sB��3�X�v��q�,�C]����J��|  ��  S�� }�FO�O�}�����LO�� @ D h�h�   @ � Ъ Q�� {� >�E� ��q� "  D�G = 'G���nP � �`���)J�    � �; �� G��bt	�Uӗ*=�@��g��qe�,���2;���'�S�.|�����<Y\��X d2rGv��q`{� p�r�}�<��g �  4�M�%R�  $ I%R ` O�����2ddتT���  E?Е<�*R�  "$!�J5�➢]��m�u���d�O����s��***����QQWB ��B����
����TTU� ��x���ݧ��e$%��Ѡ���<?�?��ƞ�R16��c��z������9E�V��w<B����fL~��ՃE,
��*��6�Y��xuYاW��Ōys<]Tb�c%���_{=w{~/x�Q&;d.�F14�J.x��G)l���w=��:�9}G�:��?�ۯYv�`�^CR��b�jbB$�\�z@�(H�Z�M<`274P�}��&�<�y��ga�,!����l����7�o����%iVO(D�"M�I�62 �4�X��J��__�2��y3OFw������O���;�5+�i*�s��5'�G$�P�,���&B�3�k��{kY<fI���|\�,���cN�m�|�T�<�uJgx\>dJ�<5:Ǆ�U�@�*��ʽ۞޳�{��^���ى��>	$x/ V,�D��(B���R%ą��P�Q�%	V4�@�B)��bX��Q�aQa � � �H��! "A� ���"�D "���eX��$40&��10��@����N��oW	�CeKͼ��mW6��ѳ�f��r�w��u}C3�do�;{��J*��D8�d(�$��p�K�H�����>=%d������\8�<�X��CF��L�	��anRFʒ2H��V��I#�����ѶxYF�`ǅ�ꋣ�P}zu��4�j+o/6v��U��輞��(�=Ճ�>�Ӛa�A80�c�O0d�zh�5�K+��<���Ŵ<ޟ�dT?`��{�޽���<4ܢي�����Vtr.��7w�4�Բٓ�S!Uq��{�dٓ6\����W��gK��cs+6��3��o�$����̙oТ����7�>H�!XU!��4���aI\cC!X`E�r2�0T0����@yͦ��9�iN�g{���h�[3Ϋ�̩��s/�����+
M��݋���N�L4F��! J`B�FB�K����T���������􎍓��y���m�`O+^��L�����~���7��G�"RH��# D�i�v�ev<���t�����%��>�3�1��y�{w�.����vQ�[Xev��#	i�B�f�g���SN�乻W�����y`�C�lJ�-8S%�?��h5.�;��x���X4�*rm��B�{6�����o�!���;+��7����N�����{Z;��_�R�Z:�/=��]�i�����t{�P�b�zӫ�]�E.�.�	RQ�	t���Є�q"F#bGF�P1�`����D 4�H1d!2A4.ص\V��!�KC�#\
h7!����*�(o���R�TRwtV��z��뻴�_�����^����)�t�V:�ɷR{N��ni0�S�#~��^�Z�	�.fK�.�i�u�R��ld�K ʪr�K�+_>q� �ְc��ZF�4<&�Z^�H��[A���<���d� P�Y"%�%�@�R�k�V�,[�V߸��(��ۣ���)&J���s^r���F&v.�o+���	����J���;�}/(�;�%.e��j�aC�	J����G��^���o�����T�ޘ��J�C6I~��g��U������ǈ1�t<��N-|F�=I�o3���=[����f�?W
\��vVNI �T�B�hƐ�|H0�B#X	E�,t���Yׯ�mܿ�t���u��dy��/��ו�d���Iޢ���ިrLM�`AAEIӭ�o��,�zaɐ��-R\J����`i�����[��w���l�����,eV����x
]n��+�򅏢`�3}�i�z����Q��ʝ�*9^�4�z黽�ufv���ۙ�c3A�%É!�����0�l�B@��(Z�PMW29F�����N��[xmof��x�i� 0~�B�a��H�d�J����b�@���H�Y#H���@�"�	�"���c$Y�I��8o�on����f���� ��$!������ӯ��7/[��{hĝ��Ũ'Z^�C�,���0��M<��bm9�m,;�W�D\R�+{Տ"d�g�(��<jhm]�'�*�e2���7�T���/sܲ��8��U����7���UY�g3΋I�+��+>$k�&oN57}�8���4��xx����4�ջ]�Xxl�ܿ��EF^Ae����ӛj�}�^vf���d�dJ��5
-`x��6��+������f�D�=��z߽�mf�}|o�x��4�5'%Uܹ�D+ $���Ź��2�D���>��|����/����{{o���o�uu6���������0'�o'0�D2Qx_c���w\�=�c���z�2��n��u�w���tc�2U����ΔO^b����"p>-I�Wc���N�%��b�f�����!�,%p#HV5�S VH\���x0�!0�&�<u�4E�zP��\�0�4B�4J
�
��
0��
���$X0¸��0b±�jF�c���HH1 `Ð�j4��i(D�
#�H&̼$"Y �FCL�v���`�^(�����''+z&�I�b����(�nm���]�bh�ͧF�F��D�r�A�� ϗ���<���D�~䜫��s`�cdZ�OW'�S�t�c�+��	�c@���D��#�j�����@����A$ b�@����mU��W�b�P�"%0g�Ŋ���vf���L���+4ll�dL�d)*�e*8��.�	��i�]�k�J��Iz���Y�ʭ�P���@�b��K��7��xB��C!�T��<�.l~>��ZD�%Z�{�v�L� �1�I�}Y�D��M��F��}��oi
m��*��\�ɑ�Y���%�s����fc��?�U[��l���� ȋc��Le�c$�0�\a�#aH2!��i�2\cRSA+�.H�Iq X44l&���6#r\��~�u�_����T�7���o:e)*��w�s��P�Wy�q���%�"���˔j!�7]�*�+�.	Mo1ĭ�Ď˔��!�$#H4�F1�4%"���٬���L�L�vC�W�$lmŮua�����]�(B���bB��KF��L��J�2Sv�\ꇚnc/�isI�L��%SM�(c�U��ܰy�
��'5��,����EL!���]���1�aHԍ�`P�Ӳ70� �ddR������Hk:XQ�%e�@�#R,����aad ă,�`V`4��q`GQ�a��H�5�XS �H0#R$'!�Ldxݪb�VK�oh�x9�q�Ձ���{\��n�u'*�,էwǴndN��i¼+�0��q:��Jٕ�N�zg������������n�D6d	�:)��&B��<��f�	����E��L2���M���]���V�9Ȑj����p������pv��d�����U��������֦(���g���[{J]�]�UZ��$�ILM|NA+�g�Di�!A��N�0� �i�81���$�w ��Hqy��4��{�.sDܸ[7�5��fP���A
0�FW���~�l��Pꈡ5��-�*m�V场��/!p��ۏ�I�A�xx�a��FH�__�&��A�w��tN�{4>���'�S�e�o'��r�g,�vEF�MLj����h�H�gBS���m��3U��L¶�
g�9KU��|��h&�Ҫ.�Kwt`ۚ%��<CI�"LL�e��$Sai�����[<q�z,�6�xi��pdli��Z�~�pӌ��{=�[�9m�ƈ^��l�L��h���w��,��D��(J����g���a�UW����-�E[w�|��ɪ�n��>#�A�#d�H��愉dHF*Q��� ��4o���ѩ RL��Z��x���+,i�pLtD����n`���p��l�;܄�xC6�5��MJ,d��&�<�P�����z��C�+�X[e�"��B�9e���ׇSLV��������2����1���@��5�L*Q ��-���
�#0�n�����<�q�V�7~{�Ziȹ�C����̿�e7��҉w�w����}�)>��{���u�>&�GV�g����m�2�CI�I��&CF��E���1��dH5p۸F� M�(jh�� b@�;!�����m�Os��2B�q���J�a6�4��]j�Ťtq!H�$i�L3�sڥ�_�X:yX���1�����j@��P���<���&{�6���R�QR��8�gU��l�lo��]r�q�p�Ѡ�ͱ�B58~Y#L��U����ڱ�V���112�G�9�-�*��ȝܴ�0�aMa�=�I �I ���|�5���w�Ώ�5mڣ34v��)�B���lޞ3�L}}������q=�oD�$��20���x�:%HGL��4 LtB�n۞l7�-*���x�0���s�&@m��P�2HR�d�\�Zј�� P4���@��f�%pB��4�N���%cVQ�Yp!�9MM�2�5f��9��%��
c�j«�$��!�03�9�h���Y����)���qߞ�^$���&0h6�`�N&���6��G�״_��    �l   m�UJ�A�m�Y[dP[z@82u��H$e��NRImm�@$A�-��I�m�4PHᶓJ"�(�G�
������l.��ŵ#�=Z&�VݵA�"�6��6�X�eg��ŵیT�Qڷ2+u]��f�m�L�q2b'W�h�U�ԅ�U�1�k%��H���g�T��ٝ���+��]<1b�3���5�P�I����^_Y���u�[Y��WH�Y�k���jh`�r�u�7n*��f�j�b�V��C&�V����Ln.�	���OZ�U��-�3���W�r��;+U]�k�*^Z��Bf8�6��֝��` H�8��km��md��zI�$�m_m�O���Cj�`+&����j�<8��q��H6�t�m�YR��XbN;]�;���o��,6�Io	 �BCZņ8��n}7�h -�;D�v�m�%��t�P��K-��`�N��]����qUU<k�{Z�����O<���ca��7�:[�gl/�ɻ+���[:%5�&�a=$��I���|�~h[(��j�&���ѷP�@�Wn�\MR�U�]�r�q��9�.�ش��M�u�UNP&R2�`U��'�9r#^�d%�c�=�j6�/�}T@�tcv�X&���pV������v;/BL+\p�4A�c�mg�.ۧ���]�re�\s��2���*�Q�|������շ(��1���h��o�ݹK�4����n }l�Pݻ`-�l�;-�ƀjnS��` X
��8���A�	yP����A�� 6��U[���z���i��-S�
�m� m��=\�Mʁl��6�-H�\�J�-C��UJ�R��l�8:������,��T��,BO,ԓT9k�s�-9�l�`�l[xZ�:��m�%6��)��i�ݶl�	$H�dh�n�m� ��76�P��S�v>�W�G] �+�vRej�U��� ��hq��Y�r(R��z	�
����"NbGѵr�k��[@-�Ѷ��ؐ���!8���l��8<�:Am9S +���T)`)"F�	Vj݀  �ڻv8�m�[|���t�Pq�@R�z�VWJ���UPmP  �����md�A�������h��մ��`�� iӶӶ���mX`  ��N�l��e�ݳ�l��� ڴ��$l  � ���f�ۀ��8 ���Y�l���"[-���]UUP&8�
�U+����� ��� 6�A �d�ڝM�� �����E�w�Cj�Bz]�e��h %'������Zm�-K5 m��f�I���ޠm��~������m���l-I����p$mm��8 �  p � [@�X��s�5���]4�8�x��P�C���E�l���m��l���hV��mճm�h��G ��m��n���ۀ9"@p-���  -��[�$.r��,���� n��T�ΏUI�O���g�*���Bn٭ts� \����٪6��v�][����A�[Hs�U�^v걶(9ȫ ]V�;�q��\�Wa^���luK���nL�K��g=6���кcc�۰�C�0�Q��6ۍv�;�N��k��V��G�b&�ͧ4[�[oR����K,l孶���l� �8NB��V�z[�q1J�=b5ɐCr��f�v�\-��]�\t:M�1�`*�;7��x.wN�uֳg��	z���x��c��@�]|*��yza:�:z
l�l����q�HsΩ��z��=8��y*f�T���F�Eu�4j������{U���VsSh8�)��m�WjtN7���r�Iv8�vy:#l��K��U�P9ݶY�q+ �<v�孺પR��j�vU��J 6,�TO[�B�pU�=���:7�dp�V_*�rt諨�,dvڍ�b�+�����O`q�nY�ю��{�;۷kk��"L����KW9pA��8��8�,6��E���[Sl�v�����`kC�I
:��n#v�ک��]\��]Ylx��,�v�g8���&n�k�X�pn�ё���'K�Rd�q��Zڹ�g�����T����n5�Ŵ���q��
��t�s���u
�l��y7��]�Hڴ�3Li�����Z�v�ej 8��]���.C)-T��`�0tc��"<u�uT�uU���e�jev�U �S<�m�IA� -6&7�*���i��<�y�P�z���Obq݋i�ۅĳ�W؍�U;�@pJOZ���N���v��\Tѡf'Y�]�n����N�9�vA͵��Y��T���˄���rD��4\�ױ�Rsk�� ֙�'a�+�#�ny����b�����Y�)�<��v�W��&�ki��A�*��u�];�p�)�5�s�����u�{�t��;5)-�=�7]�"����c�[��&!9�N	����,����Su�]�3�C�f��tݍ���#���/v��l�֏<s��:��Z�I��ɷI'8�u������v������������ir��J���`��.�ve�9��(Y]���[n�n#���D�פ$(U*mHf�
�v�i��Qٶ��*��5��|X�*U�΅Z���$`�$���t�����m hl  sl�,�Mu8�hԃ�ڪ�z��Ch�٪�iIUj����8�mٷf�&a@�c�Ͱ -� -�	f�\��"EͶ	�p�m�m6��m�m �b�� I��6� p5����� 5��@ f3�L�TڪUW�^�
m�Hl���dTCQ�4�ʫ���6 �v�ZĀ�m�HN�� ����m[m�[v�@$6� �`$ -�6إ7m�(��`  �UV�V���nUyZ��m�H  -��p��p�O��~��z���j��e*�m�-�mm�  �6��  lV�  6�@ $ l�i��Ҥ�U ݶ	��ۀ � v�X :��꣊r�Z��`�.���+[��ʼ��ܻUl��� $$qmv�E��N�鄃m�v�����`8 m�7�Xy�JLD�u]Phm�e�G  HM� pm  H��oCms��� 9��]��*�@T�UTZ�r�0��m�kZ�pJ�ڧ�o�����[e[upAo]�m��� /�u���m�� $�gqr�\���UR�TI덶���N���5�-��b@k�d`=O9fB��^U��5�U���o+��@�@]�U�����v�Ƨf�M*���;v���4qWHf�c�j���� �5T[:�k���s$��rt8c�eYINKgv�ض�	�q��4uv����En��ޝ�jU�wns�l�� ͇Ɣ���Z2�F8bЯ��;���ka+4�t��8�:��z�6��f���IN��`^��Ws�]���ź���|�n�8���j�C(m��il�GX��&�ȫEF��#rmU�O���%����_w���y3<�u��ԨT:��;!-�WU��]�[bF ��]�u �j�� 5R�; T2��pt�@l޹\�5U\Q:Ν��N�V�kX۫` $�`m�mN�I�����n%Q��7�R�U��Bu�*ԝ�5N[ptIv؝6�Kok9�� 4Q#�����S�T��$6�Cm�jMm�j���jB`)�ͫkh  ��n�6�բD։:N�`�;ug7d�y�������-�0Ⱥm p���j��;G#��zV2��S`�\F�lH�C�̭\�n:���v�;l�u���8	��T��U! �V��a������%�rбzӷ)�m�����ӳlp  �f��ܪ˳�r�����O%q%��p��{qq�DƩ�)�P;��M�Rn����n[��u*����j�+�Y
�[�I��R��I�`��:<��WT lRUJ�H ��23(
�̒0nG m��m�հH�  f�杗z�`�r�pLP үU*����e��M��Zm�qm�a��mH�U�t�5*rT@6a̴��4�WJ�%ӝ�U��X�
���O1�J� ps����wL�m&�$ m�,�m�ڐ   h�,6�BͰD�檮��V�����-U�v;!J�}�GԫJ�U]�U, ��P
�Q[���U�U*U[J�r���*�K���=J�J�Uu) 6�D	e��[%$p�K+���p����jNZ- 6�i&�b�kn   ��� F�ͤ��OB��E��n�U+q��4��RҚჀ�viv@�v��J�8����l  ]z],Ҁ rAm���[�  -�[p��u����v�` ���ܪ�Uҫ��*��U[,���`  ��
�٪�U�*ye�� ��K�$�`H�6�, ]uU^T��@K�YB.C��m������S�CؘiV�n��|jj�"I,��m�(�� ���Z�x�j?K�/Ӕ���#�tk��6�@�J��UUu* @YFе�ռ&��<�N;�e�l�l��k���-�Hl���h��Kf�̀8-�ۤm�8��[tݮ8GH�+UR��*ݵIU�t��lհ6��>�v�!j�kG�AAT�H�����B���S�
�_�:L<!d�F ,���4"�P�E�����*|/�|:hSh���X*>".�P�(��1C��EM*!�� }P|؞���pG�a�bH$`H�%��$CB.���� "�X�#�T��"`'���U���?(�|�z�ৣ�LUB(� �����x*,P=>A��I"AH*B#����
|�ꉂ;��͊��06 bz"���H�B1`���B|��G�R<SI�C� ��'�(E	 Ab$)ЀE*��}O�T�	���"�>0H�lDM��1��(0�x�Oq|\E��ר�(
'� 6�Q<Qxъ��$��i��>��G�}X�ShDqQ}E��LV��O�x���W)�+ �| � �
⥈���$ T %U"�ETׂ.�C^A|=b����������z8HFF	���
PNTKX�xz���⯠�| y�h<�@�I!2) �Qҧ�?���|�"<=m�	JTj�JXR�B��F�@���a%ed Ĥ*�F, (J[-�Ս���[XBB%��(����	%�HR�)����H2xh��T�v�}4�H��(&*{�A�gȿ@@0 8��1 �� �#�>�B#�⢢�}$���!"��PY��ز(R����U��j�"�m˲��u\ uͧ9��,pi�!!�z��X{���[��g^��ܭ��f��klxrҽ��4��qZ�ls�l�u�Ny�F��:�g̳��hz�Q1ݻ=��frX��=����`�F�jڸ�շ=���5�B�8]��dR�Q��lH�X�����y� 8�)�'n�@�1��tKɭ�mm�d�"ᮆz�V�K�'ذ��p����ں�mb�z��ru� ���K����h����	U�j�lM,�M��rC�����vL�O��M�YXMex�m���IT�!�% ���]�v0�5藩���j�O5�n9�F��ώ�7`���6�zp��	�{=x{�h2�p����Փt�&C���d��W��b���8v��<��9��쌹Z5J�vF�)�rb
�m�x4R��mn6N�\����&���3��>��[�m�s�,�;X��q7f�c�R��<���%�\ে6�<Dtna0�n �8�!�$���r�(z���z�����g�������t,�ݳ��y�]���ݰoA��W�/n�\�V�ٝb+C:AdZw=a[v�gv�̼�Ev;
ʼlrS��e�1���]p���sۈ2��vz�v��v��Y K��(+U��d`���` ��I6�H �d �]�nEi2��Ujک���b�RZj���6���W��d�fx��[8��ǧn�m�;��]��8�3��ջ�ɫw[�F�[4��B��x����X���6���*�r�`���B��u��cl�����w�p�^�cg�js��T��:7`��{陹�d�|^7�3�G-�����ccT��Q��N�r�6ۖ�'\u�������Iv2[&�od�]p���kf\j���$�mY�N���s �.'�^4ѵ�q��d��M�N��`��[ט㵔�˱*�ۚq���2�f���[��xu�g��KY6��x���[�dW�/G'=Kd�y�q�Map˚��n�kZ�ji@�\گ�O�+�?"�6#�;�PN"�6�%^*/��U�j>�/��	���x�@�=����&cnN���-�`Ѹ|$s�u���gg=��$\���'Xݥ't9C�9ݪ�H��rntk��Ζ�c6\c˝ЇZ�y{<{v�;���thҼ�Y9�o��d�����u�c�#��Y�+r�Ft*�A�\�g-������\���u��vc2s�;\�nc6gg�xy����'V�/]6�{���P�4�KT��	��T(�6^də��3»��"���{��)�ʇ7 ���xGdT�p�AnT'�ի~�}��ߧ����~�H���Ɓ�?Q��acY0mŠ^;E�^�S@�즁x�Z��@'�'�DڐZ�e4��h�ՠ^;E�w�U�V��DE"p�/;)�^YM��-����αԦ�@�m���h��h����l�:F�YJ�ɲ��Uj�L��K�\�m�6�.�bR�
ŭ�aE�6�Q���V�F�i
 ؔ��=��@�즁y�M��h�\���S��'nj]�>��}7����ꩈ�
a(��3>�`�`�l����P��4c��4�4ײ��i�Ī�=���,�����/�@���/{)�����w�ǣd�2$1��4�U{S�/{)�s�S@����r_H,��X����+r�籛�e%J��T�`�vƚ\��.F�i�mz��C�����g������8�ڞ�޵V$��$��@�,��ye4.���^�S}�fg��+��cf@�b�� ��� �w\��Ȉ�B(� �5��,"�B�T\R��9�)�qr�;!�a�lJC@��jz�e4r�h�S@�˹q����'�Ln'�^�S@��)�^YM����w����$
<�R����v�ޓ�G$��k&�����6�_�o��u�OX�Ğ	�i8~���^YM����^�S@9ŝv<q�`���Wf �v��B��ɳϦ�n��?r�h��6L�"CɃN�������z��;z��>������"5$O@�즁�YM��7'�t`��ੁ�����<��z|��6����D�s�S@���{S�/;)�~�	R�IZ+�\�n�۔�p!�R�2�,a:��=rӱ�r|�H��0�̘D؜��y�L��sXݶtBK��_��*�̈́21�)�������9�)�^YM�w/ʶ���y�n'�=�f��هD)���e�����:��%�'1�����]�Ɓ�yh]�O@�즀~�Υd�)�(��/�@��|�o����4�����h �؅1w���x]�wf����V����q�㣜 �]���HW�5��g��ʼ.����5�T�@V
�M����'C�ݷ��ն�q[��z<S;�M�:�-����u�㧑H�dV�up��lp�V����u�etn3&Nk���kZ�q�[myC�s9��X7Z�������ɝ÷^�f��u�.w.%�ㅉ�\�;��fWGk]���E��xgh��{����}���c2;db-uY�������'Nq�y����nH��u��l�:�]]ru�X�vߣ������h��/�@������w77w�=�fyD���������٠w�QbiS1B�@�,��y�M��٠^vS@�gYb&ٓ�I�h{�^�����@�즁�YM��1�3dcbR��w�?�ـ}�`��8$�;�����az�Q�rZ��6ʯo]��ud�vGh�{^�I;���7�W!�8�^A�0�������YM���ffg���= �s�̘�%�'2D�h����d>V�I$)H�A�YYa1
A��1"B:�������t+��"6J�ݜ��/� ׯ w��H�L���4�ڴֻ^��n���M��U��$�,bYh����	%=�/� }݋ om�k�h��8����$nH��q`����}]Ӏk�wX�Q7.z�H���!].X�;����k[�@��8Y��Rܘ��nFz��]n��qb���k�h��=����gYb&�sM��4�)�ϒ/��z����^vS@��u�`I��6)�0u�� ��,-!"@�(!B*&"W�P���\��0��`8m����!4�zm���e4�j�;_lz�;D�LF`�L�����0t���]���X�m�ckν�fsmm��4D��s���u۬�u���rH�I(����[�vͭON�l�C@�v���Ǡv۹�^vS@���c�2O��%��Zk�@�s@�즁��[�H�_��j|���n=����/;)�v�V�W;^�޼U&�Ld�#��^vS@�v��>�{�nLG��1W�@��P�W�("y��xnIϳ�����jI���0t���!־��>�ŀ~��9��4�Ɏ$c�h�$K؟\[��qƪ��pq�lz7��R3\쁻@=t��3s	1��F(��8����w4ܲ�k�h����Ǹ�<�R=��Y�L�o_����]`��85�d���~��;]�@��k�;m���Xu)F	@x�����ZW-zm���e4˽V<rO��%����W-z����{�~	�~�f���}w$���U*V#{woo~��]���H��۠�c�ۉ��-�s���]m�Ǌ��#����a�$���u�8-Y]mQ��X8�W;�D	K�3nyo��ر�&�,-zl^p;q�)�z�{C֋`�\M�;W�>�g���7�Üt��V����Tu/3;ûJ�����]q��t����j&�.�[�W�=p��^5�t��m�ف[V�Չ"�삜��3��,h�����{��{���}�O�r�ͨ�n�g���y^}����1�� �H���+.�T��3�12$�z��M��hs����Ld�	��y�M�ڴ
�����h�]e��(܆�x�Z\�z�e4������1Ħ#��Z\�Xݶ`��X����M2�U�U4�d�n� {�������mwNW;^��p��m}"#A����,yZ]9�B���n5��6wn�r�&)n��78l&FcmL����n���Z\�}	DB� �� }���黻*I�
+3F���}w�L�T�b���B�Hy#5��������������UA�>k揦8hW�����y۹�v�ՠ~��8��FDd��@����;�������{^�޺cbyL2}1AE&h��h�ـ9z� ׯ�!�y�M͙;e���U�Zø�6��얳��\�i��a��76R�>�}��퓂�����?�Z�{^��n��v�hV�:�H���219�@����;��������H�w/�cǿ6�D�)���,~׋��
N%b�����x����9{\:������'u�ʲ��$M��A���7L[�gt�@����RI/%�H[R�f�.�����xI}x�߳Us�;�39�;�v�P ���k�f�o\e�7��	͌$#���^[9Ծ4��|��J�B���s�2�%�X�{s�2�%��+���!�n�|Vm��lnT,�e��Z;�H�:�����^V���yYw٘��t�F#H���ɢx�O _4ˡ���K�fVdz"B���� r�6OD �������h��/�Hrߋ������Mխc(��Z1譤m+��.��K���!��p#+�
w���] m��3[!� �d$XX��v�#�~�xXO&�I�rRqN; D��?L��\>1��P4�Dு����>_UG�S ���'�z�T�HA��B�"���;A@8��ʤC�UO B��R
�_࣭{����W�zèh`��6��ۙ��JK�ߖ ���z�В^I%����hj���G1�(i��;{)�r���}_�|��kŀz!}\�S�r]�v����g��/9�5���l�n�D�lM�,�ә��k�g:a? }<��z�`��]
#��ذ����$�� ���;{w7�6z��V��b�?K�Y䒉��p��P��E��7uk z��^,��u�k׹�~�.�f?����k�4��h��~��{��lܔ�b�1
�ŞDȸĄL�БX�])uB@����^}s���{|�w4kWDں&���s�|�DB���~����} :���fLB���Lx8�L�v 7]�e��P��������î���9��:�1�6�D������s@�;w4�ڴ��� �w�(5��26�h��X��8�Z� ׯ ~�Q�:�sI@CNf���V���ՠv��h�n��s��Rc_4d����ֹ�5�ŀo��`�\��7E\�j��e]�SW8�x�DB�������pε��F"6JB�����9�p{�o}�o������OOn�^a���[&؝���p��p*QnL������lXa�x��y�n�r������C\��r9p���j�8e��6sz���;݇�#��.�nn�^�9�,v�R瓵gY��ۊtf�� �.��ۨ�)���pquˑ�.�]�V�7n,q�\��[���+��W���$㶻KVb:�9�WMu�ke0غT�ט� ��^S|��պ˒̚v�77.d��wk��h��2���\(��9�N^�M��6d"���̠^z�h��h��Zon������4�&Y3v�u�pε��^,~׋ ��u�r1��db�-�}�@�s@�{w4��h��Ǐ~m6F����^�X�X��`�78�5�6T���WSV��x�(�|��}��8�x��N��R+��悲�s�^�6n������ 9�y��n�7ģW�H�O!#SI@CNf��۹�~�\����I%�A��XδO]Uݪ��L�Ի1��W���(I/ .���ŀo��`�Ŝ�D%2}����f�%�	��}�nh�n���V���ՠw�(��

)3@�;q`�\��k�^�X�[U)ڨ��&X���v�ՠ~��h����XDD%��GR*�f��UwswuR�9Q}5�G�Qm�6�"Ћ��.+�撶?��}��dx�O��\����h����]�A�>��q�Ԩ��SJ�$�_������-���/���?Wj�}��~F16L�9��ۚI���鹉k�i��"B0"�R2@����dd�XԔ%� ~}D�U���<�ܓ���7$���~���h������}wƁ�?yh����R��� �֎����%P�Us�~t���>}�~�ذu��m��{���z���ZwH��#�Y���c��5�嚍<�+��LB�<m�.F���VJ(�	d�i��=�������jI.�ڽ�}�4�|煩$�����D�.]��I���O?��wr~����vI>���s$�{�}���U=�����R��:X)�$�����$�\�Խ��۾����$�w��I$�\��rH6,S#rn�?^�y�̒I��i�$��}��H�1&5�@��EJE�	�C�� 9�9�ݼ��d��36S�Eʩ$�s$�{�}��~H�����D���_�$��z�K���	��1ds)�{3;�RȜz��غ{v��[+��[���y����u��S�NI�݄�d.dѬ��ﭷ�~�e<�I��M�$������RO�}�M�":�/{��ƈ�Ԓ]��~��g��@ֵ~���f���p�-������Q������L�4�lɃn/ߒK����$���i�?�������O$�~����vD�d��)"QbY ���%��ﯹ��I�}�)�O}~�n�?�B?������֤�����k�c�!AE&~��]}�͒I�$��_���������βI'���n����~��2Ơ[��0;cN�QJ���>C�Wk\wSn�v���+Q�a8�Z�"x��He��`;n��Z]����v��:��Yy�]�g��^rn^n[�/gַ�ۍ����33L����i���g'a�[qt��%-�R9�h��x�N.t6�G��GXfsڵ�F�� �`�8ў^�L�3��X�t�Νz�e2��q�F�Y5g��������Ԑ�.�K�u.�[��o��F��</�ږI��5vN��\�� �����e0z,m�LCX)RIw�����ⲕ�I=��������W߲�I$���~���BYt����$����?!UT�~����I�}�)�O}~�n�I
���~��#���&��ԒW�߳�����j^��m�K���Iv�n-I$�N�Y���Y�F��r��T?����dݶ���^r�;��$��J���~�vI���*��S���U��$����ݒO����=�E}}�?~I.>�f��]��\D�c��ǫZ���43y;
\#���[pfmқ�W��l�ڿ �����.�T�U\�O}�<�I����I�ﲟ�ک'߯��vD���"r$dFH(�F�������a�)+��x���!HІI6Lİk �I0	M\M����HK	�M���o���pT�'�({�/s�7�v�~�_v����vo��fe�}5;L��0���K�f�?Wߥ�O}~�n���������K������$�k�`豼xL�*���IW߳��vI=����I'���n�?$*z��/$�z���e�.�!,�r���w��$� �~����ޒG���K�v�ߒH��m�&H�y1��9��;�<�����hK���r�ǘ�n:����.YDr�*t\����=�I��i�$��;�$������.�{����I��}+�1©�(��U��H����H?�������M�$���dy$��{�7 UU
З��LcDp��J�_/ߒK����ݻ$�Eh�� �"��P�J�1�!�"� ?�K�?�����H����y$��~��]�B��\���$��z����I'���M�$}���I?
�}�=�$��?T�Wr2�.ܗWS$�w��M�$�����%�����Iq�V�$���ְd�d@�ʯ]�����mU���4	R���L�m�2��?H�*9���w�.]��H���w�I;�g�vI:W���	-��{�ߴ��$��c�cx�bcr-I%�;f��*�zWߥd�O�}�M�$����~*�����W�.�v9	eӗW7d��_~��$���i�?� /�	]����;�$�������%�u\h���Ǒ6�$OR^�@_~���H���w�I=���$�#D`� �(��V�Pt� 2,RI��2��ӄ!��
u@����k�\ݶ��ퟯl��ˆ�˚9�m�{���m���;���}��~����$�{�}��rN~����*�R:���н���s��ݮ��5������0���ݯ�{��x>���K��؉�� ?���n�'U{ꬒI���� .�?}��I.��=�#KlɃn/ߒK������U'߾���?}��O}~�n����{ܩ��P~$4�u`)~ >���7d����y'� UU����ݒOU}��$�x��J������-˗f��G�u�w���m����ל��3=�3v�ʇ�Qֻ���9�m��љf~�R�D�.L�Mn�o�k߯9m��_ʡ����|�������>���$�Y���������J�#Jg��*Q@]�ە
0��^:F�^h�s3\ԡ0��~(�U�|`����$�5�\ѧFc�H����a#	ϵ�QZ'l�e�T=��UN��P�n���Ӹ1	\�A�!�%�XsU��z���E w�����0�H�	l-���M��q5	)h�l�|��W^�J찌�Y���͚�@�R�s~�8k[������l���S<6\#=6Hg�D d$F`A���F	Į�ib��@� �zz��FI"��BH�0 ���B0bD�XH��0���!�@?k�T6��֮���6C���ݪƅ�ʢ�鎷K��N{sw[����t��'��`-�#���qD��'<����/��d�<������L������y�8��k�u����{��N��p�]�:n����LQ�;Dt)�MӒ�;n�e�Ѭ �� t��u�ck��nc�*㜶	&�g;CHE4��:�K�7*x�;�����\��G���W3�[V��l`1@ ������Qsl�<����PٛmĄ��+!5�i]O`�S��jcm�_�3�3�i��]T�K�h錛*�;[��u�䉗��y;`��*���h�8���/sMh�{p� ��A�󗜓���>~�;�}:t�4q��Fb�e��m�o�]��3[�$9�!��,*��Pqہ�a��x4d�\�RE���=M@��z���;�\v̮�[�n�;e�l�ǥ��kD�N3\U)�V��N\�طkoX���{u�{�(�/hU�W��9���ؽ���^؇��,]r�n�.����Yp�g���s��*[�����:쵺ΧN�g�)휃v��Ŭ�ه��]���V���T�,�F���;�7-̤��p�iJ�+n��(
d�ڗs�٤
]�S3��ñ�ScHI���Ɗ6�;r"�X6,�*��S��ȵ]�Y���Kyy�p+mP��PF�%����Pg&�l���L�[[/nKֽs�i�[v��<�q��()��gppu2��RMl������9���c|��l|��KƲYY�6��z�Jzzo9:m����V��r�t��uԬ	'n�_.X�>F�F��g�dݻmp 
�2qp�y`��T�ۄ��S��W+\�=�f˷l�%�@{[b�c<FaN���1D:�mn��E�����ͪJdcKz�ѷ�me��Sd��W74L��܉4&Z�Hƒ�s��!�E��kr\��p�Zk��Ut�d��8%:�N��i�$]ݸ��g���;��H*u�f�f�U�W�=Px��TҀx����G <*�>�~1�E��T<T>Ah���[�*t�Qr�U�\���E����3�N6G6�9�z�!҈�&cM�kX�ƺ���;2l�l� �@eH�`j|�x�y9k9��!��ֶ�շ࣫��Iz�&�ܑ��{�m��دl貋�㕶�f�c�x�.�C)j�@ڎ9밯:�!j̴gg����e�ڭcgm���d�㣭���](�kv�R�\̈́\B�G>ç���b37j��/���wz���A{[���,��we��K���	��k���bf��:@��gW
�ux��v�z�;����/L{2LNX�F(�$���kRIv��7d�����IU$����n�'�~��JTEʩ.��d�O}�����wq�����O����n�'W���BJ���|���ĒO&&��ߒH�&����n��@�W����I$��ߴݒI���cMLcDr-I{��������Iu}�d�O}�ݒ~I�����I$�{���e�Ӎ�L��U��$������ G���g�;�<h�ՠUn&�D9$��	�y)��;/>�j�l�ۜJ="����*Iv*�d�f}��7bZ�ND��������,~�f��<��(P���e�Հvy��i��0�PR9�9�My����+�B�i
RR�����b)F#I��R�� ���]no����=����'�7�<�G{�E��!jKSEU�{�� ��78tDDL��ŀn�� �7.;2LN`�S#���}��.v_-�v,��l�興�ݜ`��ED�<�+������5�� �Ku��}��@��ڴ���k�L�1I�)��m�i���q�q1�\<u��[n�{s,�Y������< LI$�bm��;g���h��s伢!}A���`�3�*�&�������0nٝ	%2}��p�ذ�m�=J"��|�\ڻ��P�5f��Ӏko��"�Jb!T%��m�����@��Ul�8���*�p=�=
���� ��� ��,�����_(��$�,= �PR9��K�B������N��Xګ_0�M��\�nw>Fݭm�k;͖.�hڶ8���"��~{���9���q�ƸJ�? ��,�ծpz�tD(�!���@��{�I��K�2173@��ڷ��IL��b�>�|`��Έ��ɪ[UQ*���]�M]���b�?}��:"!)�ϱ`m>��շ*���V���`zG��Z�����b�?}Z��H|vLTc�H�1p��TA�*~T~�y����-�ٚ,�qtsuf��X�(�DD-yޟ��{ذ�m� �-lӨ.��n�J�]�����&s�^rF�V�����Lj퉞c5���	e�.YwtȪ�c��5�����^�X���
�ϱ`:����Ȯɻ�X�x�У���__���ŀ~�^,�D����5JQ��6M�Z�>�|`��ÒJ&~�}8�ذ{j�EIȤ-Ijh���P���� �i������J~ל`O.U\]��S16�����~������{��|����`��V|�������+s�ꍎ�\=�]��շ\�[�7���H��+l�k�����t��bN$�Kbgi��=:��C����zk����+��vDC�F��Y�c�ɳ����{��q�ܻ^\Qa�N��G[?�v��۩�+�T��s�ۭ�y�Q�*�m�u�U;Z X|HU�M��"CI�ظ*�'-��:�B^g3��3��I�ƓLm�4º=�{���{ԛ�|΍���&x�cH��۰@��J��}�.ß�v.1�Դrn�?���{㟝�(�s�7���,��l�5�g$��!����;L,�� hy1D�h��M�VbC�0��N��Y��󩖺��d����R-���@��ڴ����_{ۚ:�ޅ�d��lɃr-����y� �����8
"_[��9_��"n Ȍ�RHh����BI%�^w��;�ޜ�� ����l���ש�p��@��;t�jw\;���/���zq��u9zO��������o��pE\ݯ�|����\����(P�H>~��;�14�瑈&"bbqh��i�/В��D(�Q�Kά��,�ֹ�%	%脕P��ʫ�ڛ�f.��n�p��V�^,9B�3�Ӏ>�Ӏ|�gQQ*�(��������%��|���N����!z!(U����7�u�!@�SNf����h��h�{^��۹�~�o4��!�dM w[���y]�<��5�87]�wR�]�ΣJ6�o��wz�R�H�d����R/�_;�~]�z�x�B�K�ΟN��uͫ�R�K��pӺ�=
�$�UG{�ŀoWzpu�s����>u��E�U�Y2�ɚ����X�s��
�D@�$�1U�Z���A	T��a�P��~��������rO/�w7$��ŷ*�;$�W.�o��'}~��}8��u��P�
!$����`�jJ�K�)
RZ�SW8��8B�I}\�� ��,~�s�y(M�/�5r+�T ��Nu:�5������M��%M�:dr�M�&$÷l����+/����^�X�k�D(��A�>�T��TJ�U2��n�� ׯt(���Ӏ>�Ӏ~��g�%�
*��]h=&,hjb���=���v�է�>�./{�@����9Ɨq��d�����X���Ӏ}=�X�x�*	,�!I�h'T|�|��rO����Z$`ō��Z�mzon�޾��5ֹ�=
O��&ɸ��E��s�l�[�zqsW�k�
k\�.�/#��b�h�{�}��m�I2#$r>��nh��8�ny%�>�}X[�j��:���Rf��>վϾċ��-���@��,��T?u�*U/H�)IjUM\���� �/]aТ&_wb���@�q�I�LK�db�-}����}X��X���]78�\�*%;X6�����hϾ������ޜ����P�BHɆ�;��t��\��X�'v��]C^l���hj�͹�[l�`F�lTt5�̔%����v�r6�Hff-$�0$��p��4m>n�۲r\���Z�v�I鲯���5��m�Ն�N����I��b� ΃[�i淁�[`����!�����=
�DͬgL��gԮ�E���@N:z��/T������p�lV�������w��{��>���o��N�i�2n���=m�g;\��LmЪu�k��\�;Q�Ϥ��? ���USjnj��^����?O��Q�A�v,�*Z���|��N-�ڷ�}�$qv����{�ŀ}��s����Ê�vT��T�����>�}X��a�?m>��w������q|@���Cٙ�+�{��>�}8t��y%�"+m�� �~�UUA�H�3E\ݬ�ծpJ!w_�����[n�n�,T��
(�ٮ�:�����7���&q�6��:��n�i��^+�DэcȄ`�mŠZ�Z�\����DG���N�˕u�ST8���.�coz����@���j��i1�34�4�J��4i���>n��{X�Z�K�!(^IDF�/>�,������9B�
dj\�TJ�6��T����݋ ��k�<���%	U{��N��Ӏ}�.LEB���(���j�-}� ��k���!Oww�|��]4\��*K�n�pt��
#�y��>Š~��Z���\B��@�s�F�_Y4��a$_<�]�'l����xԫ�ֶxl�{����G2@5�LMȿ�g���s@���}
=	%�z�Ӏk��P\����)$���۹�~��Zk�Z��S}�z���򰪪*D�Wuk ޮ���\�j�ab�a	$
���I�(e�C�+��������!��1s���$y��j�I�0�չ�R1�w}#��%�^�؃Cvp�fd�5Y���%&5�&5�ӯ�+L�����ʄ��c�8w��6JESr�6���X�m_xQr���P��%����*T�ѩ�b�2YIF) 2V2����'�D��e>�r.�cV�#A1!$)hK�,H�84!�L��_ a��ֳS�Ѣ�
�P$ A� �dM,! 0)�	�*�5[G�K����$1Otăd��1|B�a��
�$�HA�H��
�(
��|�rl�Kr���+�t�@8��0� vDH�T8�|*�"}�!��~P=	�J����O���t����_kɹ'��{w$��ȪU'$��%�����舅/��p[<h�ՠ~��Z�r�&�_D�ـ~ݶ`�!>���ΟN�e4��&ᑐ� �! �a�m�Ʃ�-kq�'ϳ�m˺�:���P��w���g��y� ���܇�*����}�@�v�$�z">����l>V���!UJbrG�~��Zm��?w��U����9G��d�L�Ģ�Š_zx�?n�0�DB�U��z���N ~�
���<b��&�4=��.[�4
�����=��MF+HA 4�hB�}����z�>��]܌�˷.��e�X(������0۶��3;��5�$���9����Y6N�۴Zܓ�1���Sۊ&ζ�宻���w�t� �Ę�p���h�S@���{�������@�� ��� x�����5�f�vـk�� ���s�)���{�<m�_�Ĥ4W|��k��g�r��_zx�;��u?�J0�������K�]~�� ޮ��ݳ ��ڴ�s�1ژܒh����!>���:}8���<�
"/V*(Va����k3Z�]hֱ���������gd[�M\]/��6��N�������= "���!Re��qX�;o;��ɤ}��cv�^8=J�����]�R�Xzѣ�#��ˮ��WO�vN�T��ZNr�٪N�5 r�-�� �9]���,?ԧ��gg�v�dpv�� [����6��E�=��%!���VxEy�ݯn�'N^Iҫ�w[��=�����?_�;^u��9��ֽ�uٻx�ݷ��i����*V{�2ݟ���|��FL�Ģ���9�������hm�@��ڴ�zV�� F,m�qH`���rJdw^�Ӏkv�䔣�u/a�|�d��E����?u������޿�w� խ]D��	�`�@��ڴ�)�~��Z�į��^�cl=����n-��h������4�}�@�;(㛣u���,i�M�>�{��]g��4v3�(#:���v�=tU�ݜ��zpV�m��]s�ۼ���ߤ;����S��陴 ������ۼŊЈ�	!(W�)!V�(U��<X ���h��:T x���7$�y۹�v�M<�<__M�Z�ߦ"d�%�rf��?]� ����]�o���y�LP#6�8�4��� ��y۹�v�ՠuv�lU,nQDeӹ�N���Ǵ�ǥ��s�����*IlL�-tQ}]!+�$�o��|y۹�v����9�|�}0c�<&$��&��v�h��h��Z��7������&"$ԙ�_;�'>�~��t�T6�a� nZ��0A���L����{��܇�L0���FF(��?Wڴ����^,�}o� �&��WI4��Ӓ- ���o�g�/���?Wڴ�C�Y�dX�<��bΛ��qŷ�=�3��or��bY<F�#����M�U���kŀk�s�~u�|�����w� ީ=^�VZ�D��5uv�u�s�L�u>� |���^, �t�L��F,m�r8���� ��{>įo�4�|�q֮G����r���|����`�\�b��D4�ϟ�Z��ŌEC	�`�@���`�\��k� ׮��V�E��tg���l/lGQob�u�/b��KS��k�H��ܮK����m����s�ۿD$�_��ŀj�~�1�Dcb�-�}�}���E��X ����Έ������Q]3L0#m9"�/��� �;f���Z��V�ϻ�:\I4,M�Nf�w���k�� ��\�tDBR����>u'W}2#1(��94�j�?Wڴ����'�{��$��b, �ք$A�x��ַ=��z��S3d�5�%���VeǇ���&��q�2��n��>h6��:����;S
m�s��<p��^�s�.X^�-��v���h��h��Tr�&�$t:9=�-���|*��]8{toOoj�u�����P.��rn��D�HJ��vt��߾��8ۜ�讙6�[,]'5��'����tpg8:�k�f|笹�l]n�
��nX�i��g�=�V���Q�����||'۴P�iқl������ے��gsq��U^�s,��e��SJ̘�F,m�rH��Zm���v��ڴq֮F}2`��9���Y�A���Wt��k�W��c�&����l�;]�@�����w4ܹ0cW����kv�����m���Q?k��:���S��F6'!�~\�zm�����@��h�"dF!��x$Sp��ۜC���WϚ�����y���͓"Y�x�&�6�n?�{���~�]��g����!����69RgJ$�ۗ*�m��}yC11&���}~��&��}7$��נv۹�s�
܁���B��nـ~�������ŀk��w:�d��cXә#��?.v��w4�;f�m��9�Z�E1�$��*�� m�XBQ?k��w_�j�9����q7##�D�<Rb�7;F�u���h�e��ʺ��8��r����`�&)� ��٠[�M�j�-���?r�m���&!�7&�oe4�}�@��s@����˕�S�\��f�����8z�`�@D$�B)H �$	B%K�H���Հwob���OFV�m�Z�/z��h]�z����>ՠs�:\I<Ky��`��u�r�Ͽ/�}��pz�`|�y_�����'��m��w3���䧠�clg�.����9�Ԥ^7�{��7�x����j�s�X�\��ŀ?�\��i.����R�j��U��Z�<�	EQ�w�`uޜ�x�ΝKAv������UW8z�`��8yDz����ذ�����s�&4�RO��#���J�Ӏw>ŀ?���P��Z�	�H����$w�i���ŷN�ҕjJ�����x�/DD(��z~��b�ֹ�7��D�Ȯ�K���O��˙1��NK\��9��iL���f�E
���)�	�G�ȌX6�h�ՠ[׋ {Z�$��ϱ`IȔ�z���US7w8�x��P�UG��Ӏw�ذ�79��M��3��ҙSTXU�Z�9���5�Ň�D)�����Z�4a�A�� nE���}�����:w��z�`z!B�v�p��yL�&5�9�73@�����s@�z� ׯ �����,���}�	�4jI! ��8$R�֣./oF�c��tv�����)�!�}6�d�e�d�|<��=e�����L%B&pw�e�Ixˉ����la�@m�!9긚vOG�>@����0##v�HM�*>X1������x�L>%y	��ݻ۾/�����Y�EضF�j8�j��l�#v���RvQ��=pt'��"��CA��k�<���6{a_k	�����'���K��H��=�rZ���f�
��h^{���&\�@8i��>���� wg����b����q�v�nŸ�Q7Y����Ղ��=�$��u�-��\s���mT�g:��;/f�3�m��t��j���mn`ص�U��\�g�
���vj3�i�ͻ��N�[U,��8m��F�U��Bved&�RMč�
��
�N�� �I�S,ڶ� v���n��,�L ��;q+�{nz� v-H��1ӥw]�$���Y�=k{{v��֍�4��&^�n��=�n�8P��ɱ�=ƺ��w�s�'<<;�֧\�ђK�뇞�i���Q3�vj���#>��ַ���GH�佶��ɒ���r�E����M�^$'Y�uI�D[�˦t��.��w'd�/0���7+��К�������&S�C83���n�d�u����ೃ�)�Z�x���{u-q��o=���3��q7��Ų�۱�RSl^��ɸY��s��`�t����]��}Fq�8�������EU3�mh�
��ɻ*�ڶEN����.���2���`i�'Z�m�*U@@c��x�4h�	�n���lS�!U�m�����gl�]��H��+å�Zޱ���p��NV8����$F����5��3m�s`�)���`u�K�\�&��E�Z�� S���s�<'6N�9@�f��|n�t�)np�i�p���t�-�p�3�uI�C��f��H�����m�<sK�7u���\�m�*�yW\�S���ݩ�M]!\�g oj� �M�Ye�"n�+��KH��N�9���wY-��*Ί�mrV��n�@ݜ������Gn3 p����];X9�op�5f��Ӷ��t�s���jn�tGk�	7N�2q��v�t�i\�$���ƽ���g�dV�l�:���a�x�35�Ԛ�kj"���*/�£�B��@D�t)t��_0O�_�p@<D`)�!���]�>�{332�k2�354m�םk�k��e��콺��uv�8۫�;i{��;YRa��a�,hn$�t���Y[�3�z3��]���v�6:���ypq��.���g��h�������k���m���Ɠk �&�M��9ss<ˌ0�&��]��;��-����0�`��-fOB��u�n@1)��)�Xl�d�$��ٝ�ػQ����ߝ�������iɷX�4��M��f�%
s%��LC��W#��b�h���1kַLi@CS�~����/^��׋�
�G���V���*���a��s4�ڴ{w4
�k�׋<�G�U��.f�D�B�%\����{ ��� o^,�k���-���ҥT\�QUV�:OV�V�� ���$��}�`IȔ�x�����������h���]��yh��E�51dqD��&�5E�:�'=��k[n�!:�Qj���S ������CXn�nJ��EQaWUk�=��N�^,η_ľ����s@�Z0��HO� ��z�a
�2I%�?=�Xovf�z�Z�
�"cXӘ�s4:�`��âJg�>���X��WLi@CS�zon�z�V���09$�z����E�U=3T$�7uk {Z� �Q�8�N�V����;���Lc�&4���XId��v�N�v.K�ӲM9+��e�kd^+�2]m#ؒ�*��[�`u��5���!G�P���z�`.}�\�r�U"�S7f �[��(�#��X>�0ݳ=����WL�Ꙁ������;��ܓ�~��r�z1#�;x����Bp%����>����5Z0��&T�+
��X���� ��� s���'����>ڑ�U+��d�*j��l�=	u>��wv,�`��c]2�푼-�ܡ�-M�mۍ�a���:������Y0�ѝ��u���Ef �[���`]��� ���|�װ$q1	50NG�v۹�ϒ=_���O]���ؑr� �k�6fjf�`�pnهy*�O���;��,wZ˙�Q6��EW3W8Q������ ��,؉N��Q4�%%
�R$��&h�14��c�A�S��}��rN^��"��"1cJC@����w4��5�f�B���q5wE�W6�Iӳ��ti�_PL���.�x��ܰc� x��F`bō,#����$�����U���S@����wJ	<h��aWUk r۬�	)��_OwV�n���vŏ$�Ĉn=��h[^��n�U��xw*q2dXә"��-v��w4
��@�+U\"n(!&�Hh����� ��nـdG�B�_���{��n_��\�g���n����Ś�rs	��
6�W[V�Y��N�Yq�u��I�jF-�60�g�G#��v�=�nd1�h�-p��OFp7=n<B��u�b�qsn"�j!ۦ�+���-\��g:�$�`m����;��nҜ��<u��V|��t;Fy����n��ۜ����n*fu�X�m�I�u��r�WK�P��5��{߿w�{��_��V�F�y���ץ{v�M�4*��K��/λ�\�s�t��iH�p.Z��)�[e?� ���4o�$ł��Dc�q��S��	L��|`��`[u��DL�N�r"�6��XҐ�=�Om��_�H��m��;��:gVI&��:�����[�`�f�5V�xщ���4
��@�������=�Ooi��qw��#>���71��v�y�ё&�8�:g�xǰpj�(��{7U�l�9��z�S@��h���
=����`��MU�7E�*����o}����E��ԐPr�n��ً �?k�[�g�!G��~�T�7W!6��h���U{^��e4{)�w;r&�T��iE	��b�(U���X{�� m�0z�Xu4���Ud����0Qݾ?}|nh���죎a�7$�v�d7(��b�۬`7\�l"�q��ɗYȢs�,Q�F,iHh�M^� 6����0�\�tʞ������0z�Y����_m��P�
�5pW	�U"��®h����x�l�~=�R  Q�"2U��$�ܘI*(�	@^�:~��a���~xco}Q�]ʵwjI��f���"��� ����;{M� �٠����d����\ݘm��:$���~ ����h���u0Ɯ�$I&@rGˁc�e�؊�:X�:{E�H�%����pL�L��ژF�h���U���Sٙ�����nh/��y��$�QYk r۬�(���_wv,^�z""dm��f�B�!\�����;���-�s@����*����"Hȕ�\�Qsv`t%=�ߖ��ŀ9o�܃�`�D z���X1�HH@��
������!��oݯ|Fq�'�&�j�� ޫf�J=���_���h۹�qq+���A�(������]Nz�n�q\����+'���q���4bl����k�;{)�[n�? ��<hU ���$������5� m�X�V��n�В�BU@�{�Ss3t]EU���0{���;{���ՠv�S@�tvJF/�j`����}s|h��Zoe4?�>�z�߳@�}l�,hmD���78B���{�x�w�� תٹ'�H��PJ���R@��GZ)� !"ϋ;O�d�&J'�N�����A�%�n�4F�mv¯m�p �������l���4�E�3U������n�ft+۶�gKr�d���$�褈��ݬ�RCi�ڊ�Ķ0d3���t'Lp-�gj�d�!�H���#ۙy�.�7`6���xq�V	��v�JpG�磝֐헵��m@��e^6k��`J��7\���n�\5fa��>
&��<sY�\xb�BR����c�h�-ƷE��9�e[a�mͮ%/h��7v�������?޶`[ŀk�l��!λ� ���W)D�%!�^۹��bE���@�]Ӏk�s����.�3!�S�UZ�5|`i��5ֹ��� ��ڰI�B H�C@���k��x�9D�k8�>����Wv��@p�;_j�/m��;{����9��M�"R)�C252Hd���u��n��w��̺zG:�D�(����}���"�Y���#������ܔ�/l����V������bM)ۙ�v�k�E�	)�0K���1sԏ�_�f ��� �oy%�F�\�3<��8��p�;�Ok�Zm��yIM���܋9�dF27]k�[�`�-��B�w���U_��DH�"1}���e4��!(Q�������?k�`�DF��6齲�Fx��ז�nq/%p�A����y��6'9�P��:���{��|�>��7f�������0��ė��|`����OK Bm���H���_zx�9Β��Ԃ���&"d���� ��ـko����1���$۟6˸��m�5��ɒ�0��Ӌ�!��� �"B�K��!)�����)�J�B�$#�4�vs[Ѷ\&#��JH�bD�H���p��2oK��ʉBfI�ܰMf�]�5��(H��cf2t`�	�v�Mn���
nf�ah��b2`1���f�@���q����kd3	�X�3.f3d`���c�� �&8A�	+)tT�@�I��&jՁ76P�d���R�Jd�1�H��Ja.SI�!�������X��̱�5B��)�ƻ����e\�]9BU�L��'"X�vq�T��xHK��M�QN*��R��'�����_��(�X/U=j����ڟ"QP�������v� �\�E�����>rCCد��٠w��4�)�~��9�GcX� 	� �s4}�� ��]�~��޿��`�O���s$��.�Mn{qX�5:�|F�)��ж��8q�������;!t�ʳ ���v�[x���_o�b�R��Ȩ��0��興�wb�7Y|`ݳ<��6w����#�_E!�_{ۚ9��h�S@�,��qr�YS_8�&�hz!N��� }����ف��$BB �U��HB$"E)jR���>��m��_}%S$*;n�f����ͼX�U� �D}������md&Fa� Q��5>a`�{�j�3ڨ�֙�<�9ڜ��������]Q�5�MY��ͼX�V�u�0��� �Db������n����5|`��k�fy(�����T���)��E�Z�;��0�l�С%+޳Ɓ�{ۚs�bo�H��dq�v`yDK������`t/$�{ܿx�;���6)Wd
�TWX{l�<�}��~��� ��� �
�	A�X�hԋ
ʑ�$���G�����H����*��˦Rf؜�g��{�kN�2$C�-�e�/e���Muλy9��\lx�3��s�iu�6z-v�#M��>���ڵ�O9L��]PY��ܯr��	�� ��nS��/u��ȳ��y4�G9.��F�sIv&���7N���fx^Y6[a:�k�� ZYG6ۤ���bm�� �N���N�1	�x�Z76��4¶-�������;r��ݮ&��X�ջX7'�����9.:S���CU��7�����ww}6k܍b���#D�:ｹ�[�l�6u����|`�Mu)�3ɯ�Ls4{��U���S@�ot$�z%F�
�J&j�2�K
�Wf ����f�IL��ŀw�O�Ă���&!"iɡ��f|�����Xz����x��.�r\�D���W7f��� �z��r����z��ـ|7usRZ�ʨ7WGX`3��eױ����3�� zs+��T7����F�(�M���f�oi���� ۶z��C{� �}Jj���(�.���� �n�4" ��$��B��!��!2���0$XV�dJ 2CIi��U�"�(@�B�|��5".!R�p�?�%Q�o^��ذ_h�w��Y!�DcĤ��3 ����
g����^�~���Sd�ԗ"�s7f�DN�w�wS�pu���%=ݜ`H��S2#������Xu���"���wu�s��h{h��D&�!#���N)$���s��Gk�F������^'��qڿ���w;}G`SƈG��ޚ�S@�m��3��=�|-��a�dI1	NM�)�s��h��h;l�f$yu{ͬ���Xۙ"��;}�����f�H��#x�T����>�h�S@�tv5�EbMLs4:%��' 5�^ ۶`!)���`�x�3� dfGpZ��4g�}�����|`ֲpQ܇�)�֪Ǎ0]�ݍ��c���y�0�qv��^KF��N���Ǐ�>��DX�@�
I�?��~0��`ֲpu��?N�K�LDPH�Y��9m��f${��Z �u��fyB��5Ԧd:jbnh*���O������&{��`��`���X�l��@9�f�[x���X#\FB�f$���OF�M�VRH���B2��� Lo��cZB�����P���X��(�VR��$�a55w�6�,�k����O�����<�B��y�r\�i�E�e�����k���긹�5p�d�]f��/ZɆ���G\Z&��2'3����[�M �m��3�{���-~�X�Q�$��� oYx��x��`k�f�t%��X/6�1�1� ������d�;:h�����Ḡ��#�I4�w4v�h���s����[t1A"!a��s�S@��5`����ŀB�H@�D$Af`?����.��#s91� ���&�W=��x��-�<V���\t���m��[ӊ{%���ag���[���˄U��;�v��Q�Mu�3oaգV���tv�GlJ�����%�!��st�#bYI���al1��lXk���1O6��@���um�KC.:��� 7n�J�p�����z�TN	$���\l�l�M!�f����������w{��>�lx�$(Ċ�]7M�ҝ�j�-��#��[a�Ɏ��mJ6��n9x�v(�7!�;{M� �m�m��-��?ej�&���ɚ��0m��>nـk�b΅'ӳ+�]��FbD7&�}�nh�SO}�|�����@/-Md��Lnd��X
!(���0��, {��m�h����Q��j`䆁��nh�w�ko �v�������Uv�\fg����x��÷m��+�kp4)�ssۂ��`���8�6�wT����ߟ�ߦ�on�ye4m74w�DJIt۸�E���o�}�������G�~�_~���� =�x�ݪ��(F�"D����h���}�$ww^�݋ �H�t�d%��UZ��E{����z��ŀ6�,�t��0cD&h�����/{��|��b���,�M�\�����T��mtdp�U����YH{��q�sW4kw�p��9	ƝlIn�������[n�yj��m�yjk&(D�cs&D�h۹�ىＷ4����m��+�u��Ja�50�����, m����a
��PH�(�$Y�	# O`������im� �P�{���� z�� 7]UI��*�d�qL�*���w4m��/-[�{ہ�Q"0"0pN=�w4Dz!{���y�Ӌ s�����W]v�0�������d���h'�1�0]��X�]�lm�e�A�Jݷ�M�����X��ŀ9��#�wv,T��R�����	���?��Y�Q!Ϻ���X��g(I)��ï��
�T�]M� ��xm���	L��nhＷ4˩e�>���NM��`[ŀ?��X��)�J�"�
D5�w��䓾��.�u5k�2'3@��s@��nh�@�����u���&,�����mɛ]�+�U�M�v�&UF�;u�e�%0s�6&(Ҙ!72(�h��� �m����Q�C{� 7�UT.����]�W6���`�� �[ŀ?��Y�
Q�_`lH��NL�=�{s@�[Ň�L��N,_v,���S@�QtR�%T�Z�����`�Ӌ �[ŁУ�{��� jE��S2� ��j�� �nq`���o�o	4��}��ݡ�f�P�p�zu�R�	Jp�c�4kɛ1EsD��!fR�"��fl�£-E���n����W�Ǩ	r���YM1��$u\���&�&̼ڳ[I�%�tBqY���W��SÔ1�b�L�DpZ�x�fa�x���c���.h�F����'0-%�aj9<�Ga�����/G D�)b�b��lB��6@rݗw�9V�
󯼏���C���j�4m�]� ���.�T���rۻ�Sd%�܁����p���C� ye@(AT�*�z����֟� }4Od!����ϣ�X>b�q�O�sf���F� r"�)�`}@��$��$I�8br �a�8�v����Ӷ�h�.;-�{n�8��ŕ�-C��Ѷ��X�݇����Ny����(6��E4l�\�$�����P�On���v;J���ѹ��cU�"���'9�a7Ҿ[�n�[t�*�O\;�Ѝ�w<l�\���@d��5O�lh4�3k�6�J����Yocz�/��:�5��<aݤ��ܨ�[C��-U�Cd�l��9Uq�(G:1�ncmZ w;t�]����� 6�C��g��(��J����U$�,;�::WV�9)��N@LGm�@�֬v��p���PS�Pn��K����݆�F�8��Q���FM�94�uOS��d�i��vոW�w[��Ϫ۝��ͮ�3�nQC]N��t�i4�|�Y�F�m�ޝ�W�^����D^N[ɺ9�)�%]2܉,T�]>E�|]�����t��7.�ι<�u�ɵ��wi��q�'�nƥ��;���5{g�V�x�T���]7nێ.�����^����`����c��rgv;>|::��F���on�͙;SГ�>kp��Ln�^�V���-��j��I9l���X�n'h��x'U���5GR�:�4&N�i���@��m��g�����2nRș�m)<�U�+��!6��QUm[J��l(L�bɖ�F��YU�{F������q�W,�t�ɘ5��u��T.�=��N <��)usΒs��s�q�=�nG�i�\ְ sEc�h�mݬ��9׷��r�i�.nٰ��2����r2�9�;�ص!gbLg�q
�Dc�̶ڒ;���\A��Xq��7
�܆�2��Cl;��cjPyLa�|iG{N�$�me�ۄ,Eç*����@�'sۀi�
뱵/8e���\�Cؔ�Qڔf�;"�)%O7PWm�a���5KU6��� S$�Y���*�qڞ�۲�K��Һ�oYp-��kΜ*���i��D��m����K������f���u�5�3Z�u����Q6��W�^�"|A�]�|�"�j�b��0"�H��� �SI��@<E�G�~�	��/�m��#z�է:F%m������,k�����-j[>I6�JѬv�׎���0�j۠t���t��n��Bƭ��bO=v��^6k�F]q�Z�8�l��X��g5p��[���!������=m��k<�Q��^{u#4���N:�Éٗ����\�p�1��B#��M�A@��xn�=���T�b.*7.����^��ww����N�Ѭkv�3؎F�=�;�a&"�z�Ɍ�KG9���;�ܜ��.���}��Xm��5���~���Z�/��#1b'�I���h��h������ ��50P���U�W5k ��,�����2�����4ו;q�0Bnd���/-X�m��o��, �sSD�J��we\��>m��:!$���/�k�ŀ?��X(IkV�*��fbn�K��a`'i�[�7O1csd6Qደ�\i8���̻A���K�.DQ7v����`kx��s�Д%�C_v,�s.���Ӣ�9Vco���`� ��$jBIJ��k�X�^,�x�ЦF��<�$���&	���|�4v����������R�/�f5�u6�z�`6�`kx�:%�����J�˕wB�%�M�΅$)!I{���r%�bX~?~���i�Kı;�^ND�,K��ND�,x����������`��Ϋ�NF�z�d�ہ��k:8ΓO�\GJh�ef'i�����}�"�d0��Y�i�Kı>����"X�%���v��r%�bX�}���~TI�L�bX�~���ӑ,K������]7$���՘�h��4}�M6��bX�'�w�6��bX�'��xm9ı,O{���r"ؖ%�}�LG��q�$S7��}���#췽��Kı=�{�iȖ1�>�H����%`��a�"!�8���7���ND�,K�~���Kı=��p��Y��j�d�֍�"X�~Q`dO�~���Kı>����"X�%���v��r%�`~ �N����"X�%��v����c��MY\��iȖ%�b{���ӑ,K���8m9ı,O��xm9ı,N����r!���������ۦ��}\�)j��=\��$.F�]՜P0�8h�+s�]{�{���J[���33Fӑ,K���vp�r%�bX�}���r%�bX�����Kı=����Kı<>���T���e��殦��"X�%�����!�@�DȖ'߿~��Kı>���6��bX�'�}��i�6%�b_>��sT��B�i˭ND�,K���6��bX�'�w�6��c�!�2'{�ӆӑ,K����p�r%���~���v�EYm�Y�։ı=����Kı>���ND�,K߻�ND�,��x��D���ӑ,K���'���wR��
�]Y�ֈ�#G�}���Kı=����Kı=�{�iȖ%�b{�{�iȖ%�by��y�N�snσF곷<q��&�n���"Ø)�1�r����	L��;fwT�Ѵ�Kı=����Kı=�{�iȖ%�b{���ӑ,K���������$-o���Bɺ�E�ZѴ�Kı=�{�i�~E#�2%���߸m9ı,N����"X�%�����"~\��,Os�_���k%5e2捧"X�%���߸m9ı,O����ӑ,+��;�߸m9ı,O�~��iȖ%�b|d>;�������34m9ı,O����ӑ,K�����ӑ,K�����"X�%��{�ND�,KÿY���q�e���5.ӑ,K�����ӑ,K��G��߼6�D�,K�߿p�r%�bX���ND�,K��v�wn��������Y��ڒ��SD��{u��[�Y��+�nw]�;D��aX�-��8��S���SK��{d��r�8�GM�L�h�n�ء5�D��.��<u/.�=ح��R98�➮�Lc��)��FC''/F4��WX:q4�?߾��|p�����*p�ݎ�]�8Պg'nB��mҦ��Dv�ݘ�����m�{�E�m��S�����������5q�	�h�'���}��n�m{sc$���K��Nmx�c��OS��^n�z�D�,K�߻�iȖ%�b{���ӑ,K��u�e�r%�bX�}���r%�bX����SD��Y&hї4m9ı,O{���r%�bX���ND�,K��ND�,K��xm9� �L�b~��?j��d2�tL�h�r%�bX��k���r%�bX�����r%�bX��{�iȖ%�b{���ӑ,K������$�d.�n�.ӑ,K�����ӑ,K��{�ND�,K���6��bX�'{��.ӑ,K���N][5.�I�	�u�ND�,K��xm9ı,O{���r%�bX���ND�,K��ND�,K��w�2��q]�Y��U�3r�����9.:Sڇ,�v��f��0��>ӎ�!�8�D�,K�߿p�r%�bX���ND�,K��ND�,K��xm9ı,O���p���3WRff��"X�%����˴�8�H�	�Y��A�$�B�H�=QL�)�ȞD�;���iȖ%�b{߻�iȖ%�b{���ӑ,K������q�e���5.ӑ,K�����ӑ,K��~��"X�"}���ND�,K��~�.ӑ,Kľ{,��tf��,ӗZ6��bX�'{�xm9ı,O{���r%�bX���v��bX�'�w�6��bX�%���&dѓ	�5�3Fӑ,K�����"X�%��u�˴�Kı>����Kı;߻�iȖ%�by����	�u����d�,<��c��r�۫vz�dn�\��� ��\;Mn����SND�,K��{.ӑ,K�����ӑ,K���w�ӑ,K�����"X�%��{wr�ِ�5��%�ԻND�,K��ND�,K���ND�,K���6��bX�'��q9�
HRB����72Y7@\���Z6��bX�'���6��bX�'��xm9��t���H����Z�1D:��+|=��O���K��Kı?{��6��bX�'����fK�Ɇ��s4m9ı,O{��iȖ%�bw��e�r%�bX�}���r%�bX�����Kı>2�Rw-f����m9ı,N�{ٛND�,K��ND�,K���6��bX�'��y��KĻ�~����/��(���`�f1v��2yH<\bTۖ��@u�ynw���]�v�}A��ɬ\��L�yı,N���ND�,K���6��bX�'��y��Kı;��fm9ı,K簽��.��[%�r�Fӑ,K��~��! ��-�녂�
Ow��D �����;ı/��3&��Mjh��ND�,K����r%�bX����6��bX�'�w�6��bX�'{�xm9ı,N��w;�kS5��M35��K��"~��ߦm9ı,N���ND�,K���6��bX(� � �Aꮹ�|��r%�bX�}�7��.en�3D��\�r%�bX�}���r%�bX�����Kı=�wٴ�Kı;�w�6��bX�'�������n�]K�\�&E�{\�q���sc�6�F�1��d��c�^��kd>��&��u�O"X�%���p�r%�bX�����r%�bX�ϻۛ�+<��,K����ӑ,K��;e�~�\�M՗W3Fӑ,K����fӑ,K��}���r%�bX�}���r%�bX�����ı,O��ݘZṊ�ԙ���r%�bX�ϻۛND�,K��ND�,K���6��bX�'���6��bX�'�gM�Vۍ.I�n[�\�r%�bX�}���r%�bX�����Kı=�wٴ�K�lN���ͧ"X�%�|�ΓV��d��N]h�r%�bX�����Kı=�wٴ�Kı/��s[ND�,K��ND�,K�����ݿU?Ve:�kw1e��g.^췌p�'ƶ�.�9u3��n���jR"eSə�5��q��W��a�kv;..���#Zrg���q�޶W��82�>{�{]7<��b�6�v�o��}��:8N;lʽ��Sg<t��:y^9���x���։vm��4�F��@�JXv}�vn.f�5��
��:v׫�f�hsZW����;����s�/���홎kaxӫ�Kۣiޗ���"�WY^n72����n��u�.��j�+���%�bX����M�"X�%�}�{��r%�bX�}���"DȖ%���p�r%�bX�����چjf�L�&��M�"X�%�}�{��r%�bX�}���r%�bX�����Kı=�wٴ�Oɕ2%�߿y3��+5!�usY��"X�%�����iȖ%�bw�w�ӑ,!ș�߷�m9ı,K�~�m9ı,O}웓-�D�LԺ֍�"X�%����ND�,K��}�ND�,K���5��Kı>����Kı<��zvs-ԔՖk3Fӑ,K����fӑ,K��{��ӑ,K�����ӑ,K��~��"X�%��~��zu�Z�����ɻv���g�v6�s\/=LNz�ԣh;�㗱ۧx�e���Kı/��s[ND�,K��ND�,K���6��bX�'���6��bX�'�Ӧ�\�[2�Kdֵ��r%�bX�}���rE���@H�X���:�U��D0���K��6��bX�'��}�ND�,K���5��O��L�b_~���j٣4L��9u�iȖ%�bw���6��bX�'���6��bX�%���5��Kı>����Kı/��/M\�2a5��.h�r%�g�E�)�>����ӑ,Kľ����ӑ,K�����ӑ,K�����"X�%�ߴv�Kun��P�c��x�h��4N���ND�,K��ND�,K���6��bX�'���6��bX�'�_�~m�S�r��|�k�K�1��ZT��3�32mc�l�}7�,���z�׻��}���'m�:��ki�Kı;�߸m9ı,O��xm9ı,O{��m9ı,K��kiȖ%�b{�dܙoe�$�f�ִm9ı,O{���r%�bX�����r%�bX�Ͼ�kiȖ%�b}�{�i� X�%��v�Ӱ�2Y����\Ѵ�Kı=�{�iȖ%�b_;�涜�c�k��^�3&��'~.�@0) �j�^�ĜCd��6$�RH ��X�	�R�!!tK�{��ڻoTwP9D,h���Q�����G��JV�Fo{�.�<��a+���QmX@�_�%ipѶf%�bBaN�愳Adq2V_a�c��`�]���V���Z\��DcM4��%1!9w����ɚ.GaHm;����UNY�Ac%b������S��;�hF���ZB�0�
��C��)lq7)͞h<4D�������"�4�|����(�jH���!�	Cب�T ����|L@*(z�Q�؛��w�6��bX�'���6��bX�'�C�%){#uu&fh�r%�bX�Ͼ�kiȖ%�b}�{�iȖ%�b{���ӑ,K,O{���kDh���?���J�Q)�n;���r%�bX�}���r%�bX�����Kı=�{�iȖ%�b_>����"X�%�����55r�5nI-�V�=rn}�.G�F�Sl:�d���<75u:{�庲kf��f���N]h�yı,O����"X�%��{�ND�,K����l?	�&D�,N���ND�,JB�~��E�)e�U����$)!X�����?+��,K�����r%�bX����6��bX�'�w�6��bX�'~��Κ�Y��SDֳFӑ,Kľ{�s[ND�,K��ND�lK߻�ND�,K���6��bX�'��w�;m�I��u���r%�g� dN����"X�%��~��Kı=�{�iȖ%��x),i�#?pbA ����7ț�]�u��Kı?~�M�v[�I�j]kFӑ,K�����ӑ,K��	�~���%�bX����iȖ%�b}�{�iȖ%�O����Ǔ	�<�bN
bxk.������snm��˥0�qccm�\�@��{f�Ք˚6��bX�'��xm9ı,K�v�iȖ%�b}�{�iȖ%�b{���ӑ,K���|w$�/I��33Fӑ,KĿ{�n����9"X����6��bX�'߿~��Kı>����Oʪ�S"X��C��O�d0�&��kW[ND�,K�߿p�r%�bX�����K���;�߸m9ı,K߻��iȖ%�b_;;3���ˣ0�i˭ND�,K�w�6��bX�'�w�6��bX�%�v�iȖ%�b{�{�iȖ%�b_���4Iu4d�f�d��iȖ%�b{�{�iȖ%�a��~��뭧�,K����p�r%�bX�w���Kı6А�� �s�#ϧ�{��n�a�WK<����ag8v#p� ݉@^w-�"����K���v7�0�3�Eo�ŀ�!Qv�x��4v�%�W\���[(]���y��H���ζ<v�:;iک�V>]l8+���`Ӹ��2ŗ4��ղ�h�6�e�Y&텛'4�]�>z�{5��l���u�W�sf	��\�>++��a�fp��:^�l�.��,3����>����{��9��{e���]�x��ͬ���"����d�g%�\�/%�tt�9Û9+,2�M5�>Nı,K����m9ı,O~�xm9ı,O����r%�bX�����r%�bX�}��彷1�V2�kY��Kı=����Kı>�{�iȖ%�b{�{�iȖ%�by���fӑ,K��ޒݒvK�ɦj]kFӑ,K�����"X�%�����"X�%����u�ND�,K߻�ND�,K��as$���V\�4m9ĳ�"}�߼6��bX�'����ͧ"X�%��{�ND�,K���6��bX�'�{O��J[4X]k%�Ѵ�Kı>�]�fӑ,K�����"X�%����6��bX�'�w�6��bX�%���`,u۫�>��s&���cK:'�Xܚݹ�'3u-��u���892kCK��Kı=�{�iȖ%�bw���"X�%������Y�L�bX����ٛND�,K�w��ڗ-�ј[4�֍�"X�%����6��A� ���;U�o"r%���xm9ı,N������Kı=�{�iȑ�4F������n[����r��kKı>�{�iȖ%�bw�w��ND��!��;���ND�,K��߸m9ı,N�Gs���Y4�2�&��M�"X�~����3iȖ%�bw���6��bX�'{���r%�bX�w���r%�bX����grɘɢ�.����Kı>�{�iȖ%�bw���"X�%��{�ͧ"X�%��ꬅ��$)!I	�o����d���sڻ#;3����"��9�L
��1�W�ۚ0� �h�\m{Zk��~����{�O����r%�bX�w���r%�bX�{��3a�'�2%�bw���6��bX�'������$�d��幣iȖ%�b}��i�~TB9"X��_�fm9ı,N����ӑ,K�����"~U2�D�>3�t��,�S+u����iȖ%�bw�~����Kı>�{�iȖ?�!	�� D�a F0�$`#G��,Yz*>
DGf�r'�߹�iȖ%�b~�߸m9ı,O��xN��2�M\ֳ6��bY�U dN����iȖ%�b~����"X�%��{�ND�,K����r%�bX��L�s3Fal�3Z6��bX�'{���r%�bX�w���Kı;��ͧ"X�%��{�ND�,K�����w����Z���Lf��"��\;�m�á��̺|V��I��5���-s��5��'�,K���߸m9ı,N���3iȖ%�b}���ӑ,K��{�ND�,K���Κ�Y4�2�&��M�"X�%��u��m9�,��,N����ӑ,K�����ND�,K��}�ND��S"X�������L�Mh�u�ͧ"X�%��߿p�r%�bX��{�iȖ?�XdL��߷�m9ı,O�k��ͧ"X�%��n�gi.M3SY�ND�,��L�����ND�,K��~��Kı;��ͧ"X��zuYA��4��Y�@L���dN?$�&�"���{��xm9ı,O3�o�as$���VY�4m9ı,O����r%�bX��]�fӑ,K�����"X�%����6��bX�'~��ܲ���)����s��j�h94<�"�;�=��xlK��^F��"��?ku�ݍ&Ĺ[����d�,O�k��ͧ"X�%��{�ND�,K���6��bX�'��xm9�F��Ǚ�?�$*�Gn�]�b5�ı,O����r%�bX�����Kı>�{�iȖ%�b}��fӑ,K����!��fh�-�5.�Fӑ,K�����"X�%��{�ND��
�ș�k��6��bX�'~��iȖ%�b_���M]Md0��S.h�r%�bX�w���Kı>�_w3iȖ%�b}�{�iȖ%��PE���B�B��������M�Ȫ�MZ�ND�,K�u�s6��bX�����xm<�bX�'߿~��Kı=�{�iȖ%�b~�;�sǽ����[��;搦�>9"!l�N�
�Nv�E���U˲��'mŌ�"c	J%ɻ���E\"C˭�mg;��[��/�G&N&g�ќ�Eų����Xlu�fG�\�ٺ����8Mm��lT;����� ��b�֨"�8R!���0�=��y��
��Ca噻IӋ;D�v���f)�&d�\���v9�������('p��۽��w�����0�l�Nݍ�g�n��8Ѫ����,8��jj�9G=�18zH8jv���5���}ı,O��?�6��bX�'��xm9ı,O{���@'�2%�bw�w�fӑ,K��������%��XMK����Kı=�{�i�~9"X�����ӑ,K����xm9ı,O��}�ND�,K��as$��&���Ѵ�Kı<�{�iȖ%�b}�ݜ6��bX�'�}�ͧ"X�%����ͧ"X�%���vt���Ym�]fL�Ѵ�Kı;��p�r%�bX�}��6��bX�'{��6��bX�'��xm9ı,OO��xN�̙f���4m9ı,O��}�ND�,K��}�ND�,K��}�ND�,K��g�"X��������_���n�<�
o�q�;��ۚ"7x�	f��弪K����^V���jj�SiȖ%�bw�o�iȖ%�by���ӑ,K��{��iȖ%�d&�q����$)!K���h&ˡR+F�f�6��bX�'���6��C�O"/;���'{��m9ı,N���m9ı,N���m9���2"4}g�[�.�2�P��ݼF�F������ͧ"X�%���o�iȖ%�bw�o�iȖ%�by��iȖ%!I���]�*h,������K��fӑ,K��~�fӑ,K���fӑ,K��L�����ͧ"X�%��ߍ�3�h�5a5.f�ӑ,K��~�fӑ,K���fӑ,K��{�ͧ"X�%���o�i�
HRB��m��=wT��mZ�`U�wPnVu��/��:�y9�:�α��D�.Y�u$�ߞ}'��
j���XIUvd/�RB������iȖ%�bw���ӑ,K���ٰ�lD�~�pI�rvtˬ�u35*n���1B!6�p���)�b}����r%�bX�����r%�bX�w���rbX�'�Ӳo	ܶ��,�ֳ&���bX�'�}�ͧ"X�%����ͧ"X�� qB�0 A��8�E�br&���6��bX�'~���ӑ,K���ݳ:�ѫ�,ѩ��M�"X�%����ͧ"X�%��{�ͧ"X�%�����ӑ,K�ȝ�y�m9ı,K����ԅ��C	�5�5���Kı<�wٴ�Kİ��߿~�O"X�%����ӑ,K��~�fӑ,KǏ��ߟ�\�I���x�,�9��z�*p"�����Ә�&��xp9��<:kX�ݜ���kSiȖ%�bw����Kı>���m9ı,N���m9ı,O;��m9ı,N�����!4I�kZ�6��bX�'�}�ͧ ��bX�����r%�bX�{��m9ı,N���6���ʙ����f_ں2�f�&����r%�bX��w�ӑ,K���fӑ,K��{��iȖ%�b}����r%�bX�d�흅̒f�MYff�6��bX���{�ͧ"X�%�����ӑ,K���ٴ�K��iX � �B|V�௨<v�'�����Kı;�~�2�0�-�5�2fkSiȖ%�bw����Kı>���m9ı,N���m9ı,O;��m9ı,���	��``�c���h_4��1�{q��5�=��k;��i���z�yv���4m9ı,O��}�ND�,K��}�ND�,K��}��,Wșı?~��p�r%�bX����d0��2�����r%�bX�����r%�bX�w���r%�bX��{8m9ı,O��}�ND�,K�=;�Njk!��ɚ��r%�bX�w���r%�bX��{8m9�,K��fӑ,K��~�fӑ,K��;�5�u���2�&��M�"X�%�����ӑ,K��>����Kı;߷ٴ�Kı<�wٴ�Kı;�K�˵%*h-vZ�_�RB���7ՉȖ%�bw�o�iȖ%�by��iȖ%�bw����Kı<<�4���6D���M\�[uċ�\��%���e�J� �I��-�%^o�,��6��E�Pqtou�p���77�����%qV4����2��&�ѻ�Õ�1�mЗ�
M�y~,(��MnL�]R�!j0�=���]�s�������|�u���xc(r�5�I��h�]�C��K�ChB��ʑ��:�AX�XJ7M�1��'�"˻�+;��N9�8h�t�c �H$a�`BL_|�Qm�n猬���4X;�4L#��V8[��1�|39��4��j��zF��.$�"��A�[��t��ٹ��bBD�f*�[ӻ�b۩�9W��;��+�=��#�O>�}����	��A ��(a)���{��DY]��"�9��իG��M���P���7���oe1JD ��w����o���T9k�g�v�5س�2<tx{6� z��B)�'�����h��kV��3�����\��[wn����s)�9Mb�qÏj�m�ڠ�ZL/;[k�nܭRP�nL��n����k��g���d�w�i�m$MeBӨ��|���ׄ���g�\��.���ɸ׎����k��S�[�;n�Ǝ�����	�v��/]�:�ml����+��˲�Ҫ���7�= �'v� 2W������tʥ�2f���Q1�gN��+�vw�G���#�m����NWXgD�I��4�R����3��U�ԓ����L�E��.^]���8۠�w"�<�)nh�:훷u����%�hヶ������&�:�{I��
��k]WU5��3�D���f�G���8����gW�y�� i�݁�x.r�g�%�Z���rݭ�ݝ��Y9���%�q�T%z}'`oI��aS��h��b>����՝��n�ɱKӺ�)�3�%us=��8�+��H��m�.����㬑�v^u۴���il�[���@�|��Cl����e�8�l��79�E�j6!���9x1�^Tb�UY���|ӱ�0�ʫ�[�l���xyV.� 2�y5�k;$�"E�{j�<��ضWj��c"����Q�dT,�F����+�����t��@��J��l����
q˂9ݝm	0v�� (��ަ�۷3̏]��!GL�΋��.{i�cKg�w��^z�m����6�Y���OE�ݸ��`�	�s��7n�G&�lB;t��ãn��k=v.�V�K�쉎W���ɣ ��������y�u3v�i�s�LM�(��ݍ�uq�'6�r��X�e
��^Q.psP�ȷ1R����Q�t��-�ڲUq %�;`�jve�I]Wc��}���W6M���!&����@E+��*Uq��ĸ��"���5����n�U�,�/"��\��\�J�.4�͢�:���8V�9����Q�C5�\�榴j�TE�<@*��a� �� �P��)��Bp�ȋ��)CBx0<T0���ym[�G*��ʺ�Qwr�ݺ�&6|'C\ul8ݞ]�nqk��G:lō/b6�v�������=�i@KVz:�P��0���#W
����J0Eb��X&�Od�m��X)��;ֹ������ےݸ�B�s&�1Ӱ�ƞ�T�Ul��R`���71mGpF:h����d-�<p����s�|Y7Wd�u�@�=[��n��N�'nhj��X��3&|�}]�d�,�wEԦ��VL�S��Y�!���kx�ڔ7N�M��.FMm��9�Uue��R\�����B�
HRB�k�M�"X�%��{�ͧ"X�%�����ӑ,K��>����Kı<��佥̒f�MYff�6��bX�'���6��bX�'~�o�"X�%��}�siȖ%�bw�o�iȖ%�b_�����,�5�3,�jm9ı,O~��iȖ%�b}�w���K�	��=����ND�,K�߷�m9ı,O^���wf�j[�u�iȖ%�b}�w���Kı<����r%�bX�����r%�bX�����"X�%��~�%�ѫ�,ѩ�ֳiȖ%�by߷ٴ�Kı=�wٴ�Kı=���ND�,K���ͧ"Y�7��������^u�1q`�E���teKq���p;q맛��L"��0ݝ���^m0�h�5�M�"X�%��{�ͧ"X�%���^��r%�bX�g��m9ı,O;��6��bX�'~���kV�5X��,wwo��4F�{��LF��~�P6P>���ț�b~�o�m9ı,O{��M�"X�%��{�ͧ"~Pr�D�?}���5��2D�35u�iȖ%�bw;��m9ı,O>�}�ND�,K��}�ND�,H��}?i�ֈ�#G����ջ.Q�j��Y��Kı<���m9ı,O{��m9ı,O}���ӑ,K�2'u�߳iȖ%�b}��俭��K��VY��M�"X�%��{�ͧ"X�%��^��r%�bX�g��m9ı,O>�}�ND�,K�����kխ���-p�!Ɲ�s�T���� �9�롺Ꮆ ݠ��<C���9S5���bX�'��{�iȖ%�b}�w���Kı<���l?*�"dK�?{<d/�)!I
HN<�}�S5%PY2�֍�"X�%��}��Ӑ�
�r&D�=�w�m9ı,O�~���Kı<���ND� eL�b{�we��.�\�r��f�iȖ%�b{����r%�bX�����r%�x�_ԯ��4�'"}���6��bX�'�������vY,踛.�H�R]ـou�~�G� ��� ��l��nʈ�#5�	$4��w4������Ɓ�e4��F�X�H�i��ޛh�6���}���CY�X�(�U�nJ�]��O\���&��&h]����M����t��yre�"hȌ�	����:!L����>mv,���@�9�*��
< !�������`N�X��f j�uS�Z��Q�MHh�ܻ�z�Z��S@��v�b1���188�O]M���`~��>���0l ��L�8��@���h��?w�w4.T:�y� �0�1X�����ֻ��Ѷq�n8�U���˙#�bS�ai��R=�{)�w]� ���,�z� �t�\M�B�Z�.��7�l�I$�O�]� ����?w����܍L�#5�$4���`O���$�^�� ��� ߜ�u�_0��&h\���e4r�h�r�h�˹G�0Ȍ�#�;��h��?^���8�k�/�ؐ�d��ܕN�%�Bʻ.1ܷXs��]�q����Bd�=d�nxr��i�-��^�wF���o�wd�h��Z��O!���֪윉i���l�s랹�)�m�[�O�vq�>�b��Z����ǵS�W,^;n�{��Ƹ21�u��pE
F��<�P�8�� �^�[<웁�[d��tq�-��6棳�Vjj:�Ɏ�/g(�h��KCv�����.*�TG��53Xh���,�Zr܃�k�u�ne��X]�lvy�a�����6k\��آM1", (����zx�?^���8�k�;��h���:�����SSv`���<��2l�u`]�}�x��L��]H�EPY%R�X��V�m� ���`��� ��KS��#dmcn=�즁�[��~�ǋ�!N��V���WeЩ�M�h廚�ܻ�-zy�M���|�<u�v����ܙ䗄v�=I���۳�چ��6ˣ�:p㚹�t�^p㙠~�˹�qrנw���9�)�w�N�	�b�$����Y��v"6D]��l�>��0�Sŀo���%dFE����e4r�i�ϒ�{s@���q��*�X�C(܆����o��������@�;)�Ù�fY �Ԇ���.���D-�}_�z���ـ}-UL�fqm%���'��ܖ$��v�t<�L��4v;\@��h�0�A�ؼ���v���������7�`�v�Q�C�k�`q@��,&�Q5�����YM��]����@:vԲ|�����I��f��x�Ա	!APB>�$}���"ib������=���^��#S#���d�����`N�X���IBS����آ�l3	�1I�f���^��vS@�l����.������"�l���v�..���ތ����a�K�m�H�JH�(�"2,�@�;)�s]� ��<\�%�Ce�V n�ˢzdUAb,���0��3�B���k�`������.��4�21�i����`N�X����v���R⚵U35E�]+��Т!B��}Հ=w���fP(@���"�)Sl�A>v����z;�r�a~���$��,qǠw���9��~z�,��� 腵�����ɻ��ˉ
7J�m�����Y��b�N��+]��n����P1C#1�1�����w�����^���M�����5�$4����8�k�9{)�s]�:"�򛞺��H���V�}ذ��0��0��� ߵшD�)&h���9�)�w��懾��v�߳@�[Oɵ��0���h��;�ss@�m��9{)�~4������ 
�#���}w����LT֮p�	�f�M6�&6�:���^-����Ы��{t�`8)�aM�Sv+�f�3<�+]P�ϐ��Ym���NCk�\m�	�g�����U��=u�dH��bz���I�t�s8��ٌ�vM�s��� 4�L���ֱ��%�]��{^Q`��(�0 s��[}t���;�2&^r�e���JSZ�ӛ��M-lPN"5jɫ=������w���{������.:m��2lf�\\�:C�hvR/~�}����6�y���Ü�]s�H�-՞19
����;n���M���>�5~w&6�l�jL��s��h���9�)�w����T��q�0I'"Ȝ����;e4����9�w4�;R�����I�����ŀ}����Q<�q�s��e��Ƀ�幹�r۹�^�S@�l����'k28��A��!5ڐ��a�0�̨۶H���vWWaG=�1r4A�0x'�L	��&~�̀w��4s� �����ۏ~DYDdY��_}��)��ā� �C�Wh�����y>�5�ܓ�~��h��o���#�iVy��6a��`��?�X��x��l��\VFǂ�H<br幹�r۹�=�f)o��c�OEr�U35E�Sv�`6�`vـn�f �mb�o�����oA�2M�u8)���m�u�����*�F�ln�����juv�nr�n��v18�uk {��u�0�k�o p�Z�8dc�D��;�)�^[��-���e4^v�ɉ��c�h��0�k�o��.[�Q/��wm�PH\\P�V$��z�>��i��ֶ\��.�C�s����B* _��0
!CT����dBV4�PG��6�M;/7����q��% [�� e5��au�}�_�=��I
�f��^
[��3�vl(IY\cIkji=#��G�=�U��Wپeʣ�Nk�A�Ă;�.Mc���R��}�ff��8�f�1�%Ec���ĸN Ŵ�.z����՘�	�Y3>�>ߥ����!V'�N�3:�\I�P�A�Hc� y�K�c{{��T\ /����(T)jE
��І��ieڊ����c��Jd.�Y�m�S��ں��C�� �iN�Ɣk�X��P7�J���xa5�R0+�
�R�2���RWɅ�D�,i����XQ5���M%�߄��04���'���+�/�	υj�)�E�H��Cj�@N+�`�G(U�A>CG�TҠx(lv)��w>���%4�j�/.)\��f�Z����� ��v��Q
����`_,�&�r
�W*��`vـnֹ�ͬX��,����o�ȹ��+�s�/p=�]zX�U�Q�����5sζkny`]"�Gk��cv�� �mb�?6�r�����t��/H��P��QŠ^[����h���-v��$w�c^��#I�
��Z�wb��f����k�:�q�0Q�܉�����;s��}����@���X���&�f���#3e*��:}�g��������u���x@j)]78�k��X��0Q	����L�c���ۑׯ(�� �ˢ�� �ԍy"��k&4sC��g'\UU��9�X�m�����	B� ���@�n)����1G2f��n��D)�����wN �Zŀn��\��D1)���h�ՠ^v���n������ō�XdB����� �|�`�ŀ?�ـ~�����P�ǌJC@����������[�`�G})DB��ˤ�����B���[5ű�����83�e��N.�J��+��A��;���:.Z���A-�d��؈��;O�)2\�,[���v�N�+[�8��˝ƫ�G�\e	m�#�S�e@��b����!�;<�*�s�S%����jnZr�g�`ݣ�s�GZn���U��-�HvM����9�Rn�V����W��{��;��w�}��\�ہ8�sa���ۯg���۝lb,>�9�����C������=�|>�95���������74��h�S@�����u���(�nD���m��/5�X��g�D�n˪�T��tR,*nn��_�ZŇL��ŀv�� �ם�2by0�Lp�/;ss@�s@�즁�e4��u�`�xO��&h��h���;]�@������(���&HS≱����c��n�m
��C���ym�뙮���6Ɉ�H�h���;]�@��������iwM���JHh�հ�"pX�d�*�U!�� >�"&����4�w4��h�ˊ��ġ����@��������k�h���1���MI�4��h���/�@��74q��W�(�r$�^�S@�v�����/{)�{�����A>d��24|�)��q��Y�mlF�9��4ү����K<ۦ7�D�����^v���e4��h��F�'�1�d���y�nh���/{)�^YM��\&������� {����0���@��O|Q>ASx ��M|��9{�F����D��D�H�4��h�ՠ^v�4��h�K��lX��XdDr�h������/e4�XۆH@���c���'���P�;iU�anJz�v�fD������C#��;��F�{�M����h���2�F! �r#@�즁��M��h�n�@���ڸ�
&�i8h���/,���v�4��h8�ڣ���(��/,���v�4��nM�A�I$RE	Q AAa�E�US߾����w��F�<qƲ`ӆ��k�0�l�>{l��ـrP�}߽�S��Ө�m�6����<�}�՞����p��́�#&������=�;^HZ�?���m���9%���&�m��C"���N/e4�)�w���������#�i\~M��Ȱ�br���@�;u{�K��{��@��VF�y�lJC@�;u�e4r�h�S@���Y�
1yӑ�e4r�h���6���G����К`��H �#�Ga bV�g�&��+�agu�	{�E˷F.�0�m�t��ܸ�gy˃����5���r�"��������c��c1ɝձ;��g\v�t�1��Nv6\�LsIM�d�+����us]�Z�-c�+p��� ;cN�^G�]�"��md:�M�G�'5���W��ʆyq[�}� ��գ\F��z��ve����$��9颹��Q��]�5��j٬�5�dA��� �_w������u�88s�sէ��i���ƺ6��I��Kî�EM���X�9m����D�8�g���h�n�@�즀s���<pɍ��9��h�n�@�즁�YM�Ҩ��"bY0i�@��h���h��/,���:�`�a>j&9�^�S@�,��ye4.[�@�{w��b"�8h��/,����q����?��˾��6�6�t^K�N�i���G'�m�]!��lm�f��X��Q��"���~���qr�z�e4r�h\���<C$�nI����4�J��A7Ǉ% "(j�\�LE �5��srOs�Ɓye4��u�`�1$�	�Lz�e4r�h�S@���r�ˍ���i�p�9�)�w�S@���^�hn�n%�PG!�w�S@���^�h��8�����cɆL���dQ2<yGv�x9�V�۳����H�tI@��4V�9l�\�4�qr�z/e4r�h��9�]R,�'�D��=���9e4��h\���۹Ȱ&IsW5f��l�7�l��L�" HI"��D����|s���nI��k�@�X���1'���4��h\�Ǡr�S@�{)�qs���<C$��:�ۏ@�즁y�M����ٙ��\c^�d���a5���<ۀ�˫��歎͎�n@�9V�G�\�O�O �������e4��h��Z9R�q�0�,x������ye4�n-���Ç]��@M@h�ye4�n-����e4uҨ��2$1��4���Q=Z����0�l����T��e� dJZ�`E��	H��d)d�0��-�0�HR�!(^�J2D��}�:}w6"��j&9�^�S@�즁ye4
��=��%��9�a��H�)��0&����Z�@���ήu�^;gW+�F��90&")��=l�^YM�v�ٙ��z��@�X��� B6܆�x�Z\�z�e4��h\���0C$qhr�����/;)�^;V�ߕˌ�J|�y���:(�o8�;]�?�����89Te���D��sN�e4��ｾI;{�u$��5�ܓ�***��TTU��***��TTU�����ʨ����QQW�(�"��XQ �b�B+E�DYT�1DX�DX�DXE��`�$ �Q"�`�DX�AQ!E�DYE�AcE�T"$AP��`�@��EE_�*����TTU訨�EEE^"����Ш���EE_�**����QQW�QQW��(+$�k=��W`:��� ������!�} "T  �ʐ��W�IJ
"�; ��   qR�(B�U �T@(��T(P��QD$�"�A	 �P �  P P( 6 xm�h�(9�,t��:��`:p]��P ��r�9�4�8�v:4Ԛj��v�
r1;���U
8((  ,\��,=��;a���E�<x�����NC�n��z3�1�wg�j�� ��9�r��4�����{�%{���v��8��и�@ }��=m���{{x�����t�*�۽x��=�w���{�x��籸 ��Y�� <=2��wg��zw�nW<M5Kc�ˣ�{� <�(   &&�y����^�������{=�;�tփ��������:݃�����M��݇g pm�@�
�� �  \n�MCv $ LQӀk�:�� un�7 ��0l� �� ;{� ������݀� vv��F����A�@( *HA
xM4����$ i�I�j���J��      "��URbR�`      "{J�<��      "��2�T�P �    !ԩP@     �|8�Ts�Jk��6l��2��#R����"B$a!"H�B$uC�(�"E�S����jd�*�Pb�A�ʑTA�� �*�*M�5�S�	$"�Ǐ,���~��t��wVYMU2�����*U������[6(�2�&6�XB٩�e0oQ�&�SF�ވ��ۖTwgR��	�;��c��d0��	iP�.���ɖ���K�U]�!z�Q���%U�
���2t �HQc*����$��$�F���j�3�����&�XN]6-�DHX��%,e�(�0)�J�ae�&YԣLZ�Y	 F��d��L�r��YHT太�[�wZ�)4�Z��D�a1.�v.u�y�$��U�f��iв6��v.PJ���j�q*���[v(��5h7$d�&� "AA�#�T�.Z\	CF�8�!ԄG�Ql�$wˢ�:HM��ەݕ���"@�l� �n�6��bfà���֌YW5;K-聁0�L$�`����
e���]HֹdLs�F*k(`�@�K.��\�gT��۳ek��*��Y%J�B���YX�5U�E��24�T��PF�[��eU���cԮ2��h��F$�7���:Ԍ�8C��BTh$		�#P�b1�zh7��0��#�析�7�s�Rs�>��\H1[ ŋK�%�
e*41(FY	
�-n��
cJ���\a
B�E���!�eB�DV����H����ĔB�q4F�Z0�I��މLj04_�$�r�Xֱ���P$aM�q T(*�c�@ą^fA(�w|�^H�S�i
���b%@�
�u�)+zy�(�D`0��h�4��(�a�f�Ua)�<�!	��d��#!�B2@�:��X�4���nVs\HA���u ��)tH���En�_h�ea�4Da � 2
#M����|}Zf���[�(�0�r7��shu�D�br�h��e���GL*�PJ,�$i�$am��{�=a���s�^�}�w{� �J�d�M�<��x�W|�ڳb�-�&A���Ճi:`(ʻ��n�@�6 �S:h�a�R�(^=�1HY$*5�U�*5�v��0ͻ$	E���;9s��,V e�ȣ"�R�Bۻd��C�4Qĳp��4��'���9s�>AA��t7���dҳu�wuY�N�+cu�7�5R{����`�A2��Q�i�*��;@�jl7!x�Um�3(�S���o
eT�B�aVEƥPi��4��d2�­�tBY*2��Li#
2&����֍U���-�R�n�ML�[$�n�YB�n ��e����"BM�rt�#e1�)�C\�e�]���A(6E(,!V�!��ٻ4a2��r�w�6B��>���h)Uk� �@�XJ- D��!N(�)@D�b@KH�$`�F�-F�0�)aHR�c��$$H�X�"BB7 b@#�N�2$
9�ą��Fh�	t�L�ٝKwe��:��2H3Ri؜c���^����/5��1��	DB�$�9�]A��� �%:IMIb^Pࢦ`���7�^{P�s��Л󗞌��;s^����t��@5S�$
1��Sp�%�����F����p���5,��O.^�TdiX* �Lқ8�H��I�j��	�"XUJ�!�I�z2k5r�ٜ�`�$F�T��*��An�̪�&������[�T+0h.�t��р��^1���A�LDh�L��UM�9�I��L��ݤ!
0ĉ$i�,d�[�ɒ���m4�*rN`�A��
�&2�eD�7-��R��tQқci"O���;�#���c��A
�C�����B�L��[�9�$6o�2��92���ךe
Uu7Y���"U���r��++�Yd�doUz�u��б6)#��d*��:9
HI &�bH^=�6����L
��@��0
�"�M�*@!)����\t�).)PZF�4�,bbB�!�F�t���DcR��/,)S5"��u��:!�)�o�ʜ�gm���;�kq
B�M,�E����m�*w|%���A
��{�V�*v��U��֥ren�,�A a
-�
#.���2^�5�W���V<F�R@��f0���!Lj5
�������zN��Z1#�����@�h�(��J�V�!�y"�[�Gf�Й 1��9�\��`��3lؽ:$&3Bݙ����4J�f͉5�w���00����
b�6������RH��7Y���SeHI��D#)˫��spm*� 9�RM��u�aR9�^e|�}��Sd��-Ԃ	GU�X��q�_�����"��H1$Va�ݲ��e�KÒ��%�^��Ad#L
e�$$�0��e��aBI��^*�E(�CV�%^:)(*Cf:#L(!M��$ Q�+w�-�o�����'Ƙ�H��4��և��;*BBJ���u��w �Uc���L�e�M���^a�����1I!	"�I�THں8Z^��ˆoBVQ*�U����hsV�Vl�I�R�j�"�2'q�Y��uݞq��9�y�׶���+l�5�UL�t�a����*��0�a�h��y�ޓP��HU��N����#5���Xe��I7D�Q����W3��e���(��)�E�.a����	RF��l1!D���bCn�[�0��Uʺː�Y{�"PơVf
$�H���(��M	r @�D�!#P���J!.1!L�0��P�Jmd %����,�RX��� ��V�%2�B��ȭX�Ȑ)-@!0�F#Q�p�)-�i-3AD(*�B)$(�lV6qI�{Õ�h@�����b]�.Ѭ�DgS�˲���].Ĳ�8�F���Ã�&7�׎1�b���`        m�     �`z  @       =�                                                                            �P�                                                                             ?�    \��+o-��V�<��l�N�5X��[l�m��hSl��Ji�Bj�ڮ�y]�X��u�ؠ��^�Yn�[NI飪OCjRw3��ۖ;V؀��m�ݑd�]��`q;/:\G������I��L��ê�ggRj�v��Y\ ���5R����x�1i��Ҫga��6�����A�+)�5*�3�1ue�.�(�R�H<�h �B�uk3-��$�$�YM�ZK:�۶�3��n��|� c�Up��Pq*�
������  I'p-�k�� ��h-�m��L V�JͲt� H�m$���VUUU�
���;i+6m��`�H'Ju�TF/Z4P s�V�Q �`�n�f�Z�B�傠y�hc;Y%vVS"�j�*��k(0�;q֮����t�U�"��W]�+o.���ћ��(6�n��:\4�`�R��A���w6�i���<l�nҫ�$�CuUlI�lܐ�^���� $�m�Y��,�b� �`۰p\���y�MU*�@R�@�6�05�ɰ�T�d�ⶊXWX���6��\,Nݝ�Ul�J���[x�6*"�i
�z���[�櫩M���RRK�8R��b��]�%�l ��` ���;dn�s��ɪ	�Uc[l
Yаܱ�ӜY�׮
�MU*�նRu3c<y&l@��Kulٶ�o ���j W%Hͷ7^�� �檪UC��z�vv���=U��sv���tXw?������@���<[�<��!��ѵK�E�؊���jvWq�Qǆ�Btc��Un�l�n�*y�Q�	���Ůs����4�Q�;�W*�=q�43e�,�n�dL5U�g�RCcm�h�Krs��ĠG8�]��᫝ �F�,��St��]C�2J�@R�E�A:9#m�l)��A��Y�*vFW��s+R����[���(�M�pmU����WT�p����p -��:P��&�]�[n [Am m��.�9�N��Ca���1� H��NQ��m
��� ��h��}]�}ee��)`����1��l�*�
y��4(�� ,b6�V�����Ik��&�K�q�����`۪c�F��G�GJ:㊬c<;'w�5���(f.v�S��>�F�}��y�e4��:�	���4ʕ{Yy3�t��z1Davi`�omU[.��B�>��I��6@��ؕ2�l�g�2BD�ɠv���ّ�򃍱�g!�6�j�#-�6�ә���m\],�^�`���jWf�����:UZ�����[A��i��Hp ����m�j��֙��h4�^jTۍ��j�ꀯ����KVy�e��x���Ut��m���zk��6�  ���gm��l�8� =&�[j�U:20�WB�5UUTݣ��Wf��v����R�*�]pP�X*���A��� �\�֠�m��F�$�o���ꪥ�Td)YZ��s��L�k��앸��R�V��!K�,�TUUt�����Ur�l��3�W/p]U*��k�:��6�GiV[����
��j%�t��9h�v��JD]�Fj�P,v�q�M�8�5UP
kkpl����gӃ��KU;�/b����x�x�Icn��tݣ̸�Ĵ*�[8���T��b�[C��g�V�������3�����n
n�Ʃ���P Kun�K=�+@b�g��yGm�D��TN5���R�vd�i�o��n�n�G����{�^K��9-,Y�[�e�Ī���V�)P]��[ se��-�hS�u���W��-T�TIU��컧�VU�t��P�P��ݠ�;N�%.�� 8ǩWT��j�������Z�I�� ���t��,X�U�AWN����f�i%���z@�@	�m�m�  m�m�-hdH���ѮƋ�����R��¬7F���pl��    $ � 6�m��pH� ��  �eλj�vH�)v��^+i6�� -�m�  l �[�ޠ ��bڶ��)v�   $^� ����N�M��[\ ���,�Ā��[�ף� m��   
�,*�U[J�����,d�fU���Z  m�^�gtmǓY�F��3׍���mҽ���Y��u���a3�t+z�p�������Q�`T�UOgPtk���H�bdB��
��u(�U�X�Xg��]��ح��U%w���V�VõP�Clj�a [m�Cm�8[@��m�h 	   �\p �-�+k���ԙ,�dnL�K[���ɰ7*�J�R�J�UP�H m�5өX6�HYBE��)�+� ��݉Z��Onb�k��K�;�51Gf���n�����p��#m�vR���-��JH� ��L�u����`�VEe��Im �lI��I���%M�H���קz^��nө��ַ9����EG��^J�պ�n��{W��n��Ԯ+m��*�;s։mH[pm�m��� �$m�a^@���A��ۮ�k�n��R�c
��*�WT_-�Ip0 6ݼ�-�:rŽt� i�:�&�	8 �`���o���36瑨r��]mli�[� �  l��   [D��lm�[u�2I�@6֭Ä�Hm���d[IbM��l�j���v�V�U�d'���]����b���;pr1U>e֊����ҧrt�x6��i��ܝ��Btp�m�R��S8�I� �����r�ܵ�j�i��FEz��S�U�\�*�� ��� m� 8��6ۆդ�4�� d  [@  H-���XySI�Ѷ�l��mհ+m��� �%%���k�k_F�"F�ń2��F_ğ�>G��� #�i*�M�Sb8�_���J)Q��"�/E�dA�v����[C���k�� "
b;N
�@@�U� �ڽ��N"��� HmӠ&.��6H�
tҥ*��J��L@��A6`*O�6$�:�j�D���=-��;�4���]����$�"A`@=W��S����* O�A�������@�|�!�4��I���-,4�'%!�hX�T�4�v�tP8�t� ����iS�9�R24,I�H-��lM t>��E�]��T�D苴 �c��u'Q!�z��4��|!��	�0M�� ��`��:��P�
�
НPb��+����j��B���D$ ��'�A�U>BА`��4��t/�(pC��[�T� A�!,���նp���'���'$�0@�[Ch|�����B���
�RP,@��B�R�(`���C�B���8�R٢A�`A$"�#$!H��H�&}F����G`06���G�0V��>`Fd���'ːF�R��S@l�@.*����]�"��¨�"I��>T�~�#�@�C�R��P8AD�J�5�������a�m���               m�              �2u�R���km�����\�n���n���4�tY8�X&6���f��eFz��2F�蠁v�o-Iy:��*�K��\9�==)Cܕ��S���upAҜQ�̉{����6�m�$���k�K�5ض�'��̹�� v��coWlQ���\a�,�t���m��W;V�K��-�&-�99-8v��.��n깤��м�ˮ\A���9H೶�ӗ��gT�ڲe+��\��V�0!k����H�gI�v��["6'^yH�T%� �]��C'�-Ջb�-�e�.8�	�
�U�VZͬ#k�jvV	UmR
Чd������ݳn���Fd�jvӝt�ݻ*��(���K�Ωl���v�LB4�Eq�q��_h��n���I1��97U�]��-�Ё�\AӚL�N�MїA*:A�D�N��l��l�풪��N�փ� `����;#%���v����<��v��N$�s�6��HMUT�P�]=r�=*���kf��'X�\q�FuJt�N�K]�O�D�bܷ�Y���H����e#�P�,�O�G�:)Vx6��e��1�ݼ���B�+�MS��Jae.��Ll7ltOMV�Y�]J����q���| ��¯�@�h& |��ڪ�����N�x(�C�P�P�!���EC��y�?z��� m�UUUI��MF@�Z�̻kjI�\Wn9�	�n���mtσ����Z��넺�|7���mie�i��t�i8bL<
���o캓T���]hs-P{WVغܱ7\\.�X��¡���n֗�+����=����o�}�eC�M�&����r=����`�{g~I���~?������ �^����s%2�%��������q[���)�%�xì�+�\f���ʒ�)�$���Vn������Q�\4�T/��f��]Ͽ|�;�����K9�)2�ۣv�yA링����j��ٲS�ܹi���g:����q���.n��d���H^���Gt�Pm��k�� ��$ �-&�^w1Y��7�goT�eK�Òڡ}��7�g�����m9��Mӌ� �u��wk�@���6�e�m)A�hL��m�@�w.a.���yV���AH4Q-�����{\f���ʒ�Ԓ�^w1Y��7�g�����zJ�����{��Z턊G�#"�8t�o[s�Y)̉n\��7�g:�b���^wKR�r)*xì�+�\f�����m��L �6L�e�R�1�������^��� �HA�ZM���b�u�o �ʗ%�%�B��� D#{�Q���y��s%2�%���8G�W�b��q[��P% �D�B�u��vsQ� ��6����ʗ$4ڒY���+3\f�p�Q���m9lJM�	�9�N��!�ڱX+��fHn
i�dˆr�_o8��(��@"��b�x���Ȗ�̷�B�u��vs�� �RT0�W�����{�1w��6KI�47�b���o�goT�eK�Ò�о�q��(�������w��~}~��o�     ��i�]��]mF�:�&�����I�U u��וٲ�s���3p�ܙ��\Vκ�`������@=�c���ɻg�.��H9\�in[Bt��TŰ����M����9@��.x냧"-� *�99}Zċ�M~���}���WW���������M�;6�n�sE����m�e���3ϙ�3�w1]���w�@��e�<| W�����7�Vb�*\��jIf/;���q��3�u��.i�C�@=�Toypïy���̔�D�.Zq��3�w1]���D���6�l�E��2{6�6�vuY8:�^ŉ�VəX(�NZ���YIX����{_� ��(fhrB��l����!Χ�Lj���(<C`����-����uM�FT�,9-���3ypî�y���KaK�=�P�>O�C����3`�*j$��0������
3��m��M73$��Lu4q��ϵ��Ɋufv`̒�M&ܩrCM�%���b�5�o!G:�A\0�j��s��B��u�1W<|�NdKr���8E� � ���чb��c/5�^w	jRK)*xì�+�\f�]�rB��l��s��3yp�q���l6)�����u�_e��R��x�un�.��.\�Z��2��a�mX�{�3ypî�y���KaK���4t�_��{���w���Ph�e�xü�+�\e�1{�\�.mI,��s��2���� ��4�R5��{��Y�V8e�^��s�Dnw�Y���X7�6�l�nCN�a�'^�ױ�)�{H	f�gk5BL��U�{���ާ��q���Z����)P���1]��3y����d��1{��f���(鎺�����Xr\���37����8����6�Zq���0������9� �	A�=	$���m��`   �/]�"s��n��[��:�U��ը�Iq%ː�y2s�l7.���Hqɇnn��*�����!�c��n+g���닂���:�9ʄvs���F��Ş<V6I}q�n�1�ӂ�h�3������f\��U�/3b���҆���᪩آT�4��a��Wpp�j�l����2�E�-����1[�q�����mI,�����37������.iˡ}��3y�:a��s��)̉n\��3y�:a��ݮ33�KR�rYE*xû�+�\fo1����a�Km+���*<e�Ԡs�.��qz�b/g\坸��<����{���f��" ,�e�hFSS,9.]��:�="���!�M؆�CF^��S����~�>3-��,�Zq���0�������
FJL�B�wx�wk���/u-����i�^�1Y��3y�:cѕy��mᎤ��9w,�r+�n���X��r&�����]����3y�:a��s��)̉n\��3y�:a��ݯ� ���&fYF�G'���3��Z1�+���,^�w��J���9Zֆ�N5L�.�*k_��F#aH�$�A�	$$�+�-N
F���9�Cw�o(k�Q@bS���箳�t�C��+�b�L���恂�Ka�K�Г��IT�p�J5��[É����"�#Rĩ*�K*Yl `@$$Z�<�Qc�M,���6�
�?���벳De�@����k* �T�^ 3A%Ѕ2Ј	 �e*�����|)���=��?~eҊhV
%�"9BO�D�:$�,�R�6��4~�@��A�Wy���aC3Y�6KI���+7\Vo1����˜Ќ��Xs�˫��qY�b��}x��~�Fº�*�n�{
�u�l���g�j���i����l)`��y�:a���"����{{�ʉA�d�t,����b��qW���y/L�Hm��f7�|�f��|Ş0�ւ�a�.���*/;�Y�4D|">IJ�������Rү�v�`�����z}�^U�YYx���g�@�5��}�b��Q���m���N��՘p��g%�������������\�9��<�b���DA��,n�3!�i6b��� 7��/;�Q���	nN�FSS,9*]��U�? l��k���i��,�� �w���{������2�PrY2�<c� |y�c>��+7�z�'�'��ϛ��߀     Il��/�Gj�2F�T�����0�d�r��O]m�K��B�ۥY&�tRH�m��ç�h���(���X��ힹծ H�^4�uδ��K]Lltcb.Ǭ��y��U�����J*���!���ʖ�1-Ď���@@$3n�m�mCV��m��@C�s�V�kc������?m�JIf=�s��+7�D,��bh-�E:�s� ���xïc� ���Js"[�-8��1GH���� �}�g�y�f}�Z���e�z���+��8@��y����A�ZM���1�@�g{��|�1U@���m��i�חn��Wl<��8��nκ#u�~}��wp��8d.����{��]��jv~@Ȋ4s������yU3�&^:�bAO�	��������ww���	�B�������L�CO�*�����_w��Զe0KM�%�������q[�c� \��bh-�	:�s���P��*��www��} ��IU�+1�;n<��z��b:��m^{����L��D�.Zq���Q�_g��B��q}��&fYE*x� .�X�{�VA���Ȑ�d̤cw�b�u��(*��y�t:?�T��}��Lz�o2��a�)�� g{���(�" �k���m9�2Ĵ�|��>�����s�������6�e�%�)'3���ǵ=�l;�u����
	&�� 	m�2�PrY2�F�1U��}��  _w���e2Cm����?�? �s�{{߱�k�E����Y�e��	:�y�n��@�"�b���\��%�fVV^ ������:׹���*)#��@@��h#���p� ��/;ޗ)Jfe�R�g�x�w�B��q[�c�/�m�JE0��ܙA��X�`5��<���0X� CUFD�&e#�|�f����E<c�s����AN����"�G=��rz:��gP���Va%�i��y�:G�= DNg��}��^f�&��̹�Vf�r���^�p���X���c}䏥2BM�%������ 3����b��Y �>I&�m��m�    ܵ�E�k��v��N,�C��s�;�F�qƖy�K�A�AA�������-��xָ�=C���H�����e�۫u�u*�x�,)c<Ӻ(r�iƬV��9�[���utVۖ�8-� Hw�^Ud.��Lʻ0��S���.I�{ ��M�Yf:hYV���K�ْ�n�q��m]��{�_|��%�a'����+w����"~�/92Qrr�����1w�b��} }��R�S3,��>1U��~�8��1C3Y�!əH��Dz Ow�1��8�ߘ� E��\�e52ÐS�~�8����<a���d�m�Ĕ��(,��Ê�ۇn�q�N�u�BeHr��@��te��2Ĵ���0�y� B��q���2�4Y2�=2	�К�.)�2���)�B:e��\���l|��7�s��8��? �H��HM��f3��+7X�" y�b�w�Aa%�iK�� @�{���(� ��f��y2Qrl��|Ǡ@<b���{��d��m�'���l#n��.�g�c�{ٓg�v>�}"�(�c�<�b��~� ���7y�l���_���舜�y�o�b���#��
U��\ʗY�������`��$G���� ���4���U�U�7*�l(�q|)�����}�g�km�K`�� �w�Y�׌h�~�TooxL�B'&[�g�x@�͡~�8����޻�_� љ�l���/�ϵ���b��m n��}��#R�%6�%��w���qW��B�@��!��4�п{����������z�|�̔\��-���1[1� @o��3��>�L�fYE*�Xk�������H�j�����T"@eи' ����'�f��8s��E^��7�����s�z�7�1[ }g/m�ؔ�f��9���8��o�7��~� C�5AML��x7�qW��l�@ @"��Ǐ��l�[,�UB�7����{������2�B�K`�C�L<�z"" 9�s������Ly�veQ������;������~_��O�b��C�%�iK��}�>��  f���v���aG_m�:zȐa$`HH_���$�Z=�M���q�譑[J@�@!��c���UH�٢�؛Hm��t��n�G����I�S(
����Bђ	�hH[D�(��Jp2�t��$�!"F*\5�, @��a�	�H�f�X��		z���;�ny���|�z��_�o_m�� ��                          ��    F���'m�pXxqj@��)�{%�j�Tu%[n��{@�Q!��ֶ�Ue���n
�N��j3GIV:��\)T��;19Ys���G�\�֝�n��4OFt�lviM���b���۶u��v��Z�]n�wV(�r�'��pj�۹]=Vf�u���%���b��hB���ܻ��<]��X�F�ã'W��ʫ�c5WW�r9�L�n����Zy �'jC��,u����`��u�ٻm���L�����l��;�Dn������>
/L��t��qS��v��h��5�-`<���Z/*Ʒ�;\�h	�GM��clS�қ}�������\��{6ɤGb��%ۣ�9���D��ŜVG;�����f��}}���Re����b|�I�͑�A���Y�����3xGi�Ђ��N�A*:B����&6�Յ��meZL𽭓�0Tjj�ΆBu���FA9��Jd{r�=ix�:�	�f;#�U�����z�=�]�����pqm�r������p[9�5jۦ��=[��v�%�����ˣ"[`��vwQ-�Ɖ:W[:���a�n`��i88������ո؎�9`�B/*��
nK����j�.Ix��6ۃV��]����CI�?(��_��W���
Z?,G�q��T4'T>���� ���؀�R���m�     
�y��z�;M���'X���^�)a�S��5�i�\�(\s��Z^�]]�UM��:��۶���ڞ]hĘ��N'^f�9�s��KK�]ve�gk�<��vnR��@��\��o�S|���T�%�PN�U��v�C�E�W��ffd��(�ɓ�'	p��W��=<�ə-�*aMD Ѧ)���[e��|�na�y�C=�qy��R�S3,��Gd�H���"�y���8�ߟ��̉&�S����p��8����e52Ò���"�ި��8ۑ�"{5�w6�d�&X-8��~�x����Y''zY&��}z�~u��}���]�e���ҍmҡ���`�V+`��>�w�'"�T�Ix�h>�@{�� | D�{�O}���H9�$��VZ쌊�H�"iIA!#�#L �Na�M�P�2��uQ'w�TI=����$s��� ��
�T�7��́��l�铲hM��Q�(SHI0؉��� �ϮPd}��v��y]ʤ��L�ER`s@w�z�%�}�����<n���3��;Z/�l�m3l�k�%����G?�{������2��$����o7j�7���| �C�� e�lQ4�eB��K�~���K���;&�s��#c�?O��%8L�ԓ�{��$�r�l��ʺ ���#��W(���2�IT�I0�" �!/�Q''zY&��j���{�`gr���%UP�X8P�G�3����-ݴ�IB�STMMD��G@��lPs��ƭV9BL$���8h��J\�'}�Uos[ ۞��!sy(Y�9
`I	&�9����ɠ.o%��o~�d���RT�&��i0ɠ=>�F}3}���́���L�E �������r�Ҥ���֤��kR~!�< �#b|4�C���W$��}��]eL2�J���l�DG��3������I�z��4l�ӓU�f�L[��;+q��0j�X�?�w'I!(�P*^�y���=>��rݭ�noH����)I�m�~�>�	��d���Uow�D��y���UB�`l�JטٿD���`\�@z���TBAU*Xd}7��`^�6�J����٫�%
`I	&�}TI�DG�$��K$��mQ&�B�(M,�V���!����Wٙ���    �]5%����z�d������D܂'�fj�$ω[gQsU�K^�/[=ic�`�.j���ڜh�E��������}�F.��ٶ��$:�� &C6P1V��ٳ�pc��s8�Dܻ�\2�&��w]Q�ww�|����z��7`ךv��m.��hp��9g��g����}�:I����L��ip<P�\����G���3��`dw~d�TR	*�Nl��6�5�=:W}��{�yM*�B��K���=����}3s�sy(������L�&��M���<P�\���}ݾ`��$����
R`nx�O�"G�kޛ$��z��{�U{��*a/k4�y�K�q��L�x;=�FJ�L���~��_M%U@���(y����}��(���p�����M��T���E`i��P/�{��~֤����7[������\�\��-�$��Q'�J:#雛�@{�[�]��ji4R�蟇�-I�ޖI��ڢxDD�w�`^��&B��C'6P�۽TI��5v�m��E��$8i�J�D7kpzP&��0a�%9t�Դ\�.l�����7����Ӣ">�!sy(�ͤ���L�ZtI��U}>" H��Q'gzY&��j�"  L���	l0XA0�$���f�|���`�D�B�H�P���$i�!�N�����~ʢN��TI��)q)��,�> @�]�d���M�����|@_�w���%Cd�.h�}�D�@����''�no%�~����m��-�ܲ���U�<cnPr�p�X��d������ �L	!%�/w�ӥ�����!�{�[�&R$�$�LN��}2zo%��l^s���#��}Tg~d�U ��`l��@;�l�g7��$���I����M&%54N�\���I;߽�I7_K��18�<���Ҁ���I)DʁR`]�6�JϮPo[�}�D���I(I�T��@,q�M��wr�;i������]Ntv��{�}��ϮP��DG�/7���WT�����C�6WDL�y��y��8W� }9��\D�l���~�}TI��l��Ҁ��J�5EtH�(T�����02t���޾l]n�L�D�U&�}꼖^s`z�%��ߞ��ݶ      7/K��I�I�[v�ra�2�%v�e������F��v�v�6�AF{^�n��������\7��<D���-*���9����[t�o���}�+�+���ܝs�*H{'Wm�:���8֭�r��;]�!�����{�����;�磌�\�׫\�ur�A�e<�jD�P�Q���2J	��@��Ҁ�^6�?>�Hd�@鼊&�J�AR�����}��y��:P}r���"&O���m��`˒ӢNoz��s��&no%���^t*P�P�Q)&k�$���$���D���ﲉ=�_T�����C�6P���y��O��i'���|�K���`�V�����)�PecM�;q�iUJ��_$R��vw6�5�=8~�����Pf��"�(I���o�S����	("Y�1�(�bHH23B����h*?}5_K�~���N߶��@�2sWޒfXs2���rx�MM��D���߽TI���D�hf�d*�IT0.se~�l^kd�@qqD��9�MK	���}����舼����Ҁs����I.�2ƇkY�b�7�m�<]:1�� ���ww���G]D�K�^�6�
�랈��_k`�ЩB�B�P�&�
������{�U�D${�0�)�M��f�>�},���Tdpޮ� ��N�� [ ���"�ByG�T��MA�Y>S��C|"�$a
H� ��E
�:6��)$��-s2�ؑ�cZ�D�ҧ�A�q�5�rV�#Ԣ�D�+kî|U�2^!2���A��h�H!��C8'1v]��j�,�4���H�%V�R�hM�
z��FJe]W�l)�[E8B1 p�V�T���u�8ā1�j0cj��k�v��W�K@�Q�6��'�tHU:=U��E���W��!�6I�
G�b	@l]!d@@�̾�$��D��hJ���R扑��wy�{���(O�P��AJ�`{3[���7���w�^����_ߠ%�bk:u�;m���Ҷz�vn٭I���>�I̓*��54�Δ��(�c�"#�}�]w~l���!T�J����(�c`{3[ӅtDDL��7�D�R�d�sD�o�TI�ު?�� %��;;��?O٩7!���%�D� Nw}�I9_K�n���<��"�P! �o�tI;���,4Xi�$��D;�>���_k`{3����IT꘠3/<����sѝ���]�m�y����w��?f�i�X=�P����g��DzB�J��D�K�ET�`u���5�=8P�\���.�U�E"�I�{���(ﾙ���_k`z�:d��$�3SI����}X��7kD�~����́��L�R	*��h��������tI�҉?� �U�I%���m��    7]�y�6T	7���,O)�]��5T�g:9���ϖ���pG��2��q���
�Ûn΍�Ɖ���3�vL�����8$:�H9]�n��$�<�g;JV�(5Z�!�a0�s�S���L��͒�	!��JP��� �j�WW.n��`�U�}���%�l�2�Z���'w����%ԅ*��g���́����(�X���ʤ�(R T�y��DL�:Pu������!��
�((�I�s�r�$ D%���O��Usy�i�RH�07+D{1�2�[�"n��=���q}J)	*}���F���Δ��@z'��$�	H�$"Tʉ��b�^ء=kg�)��JQ5R*�R!J�$�y����U����l�ޙ&iI52I�n�.�z1���#ݍ
��}�� =ۭ������a0U"f�`nV��cg};�́s� yϮ(�U*)
U.2>���sy�$7���@l�uRS
)*L�����@_���q�2&�I$���Jj��t��b.��.ϵݹLh�RKק���L��I��?$���@_��{������l�QSP�*�����l�����]�����QHIP���l��ȇР~R��q|;�ץ�9��d�{���"�(I�����(�X��'����ޙ&iI52I���������l�n��P�D�Jj%m�|a�Q�s<�(�S�!I!T�J���Z /ٵD����@�b'g�N��e5,&T�����}�Dɻ��:P���וIL(P�A)0/3[�
;�"f�@u�6��	R�(�
Ra�9ZP����`�>�{쇓]l�Q[K�R���ͭ��7�7y�'��i'�^��/eUm��Kc���cb�� =ժ�<扪�qP�}I
i*<��`^f��� D9'5id���x\��r��Nn����	��$�.,�_g�^'uw�f��S%M&O��@>�l�����L�R	*���G﫿>��No�TO� @�.I�[��)� �C߳�`~��7��'��^'���R�X�"H�0�<��yӻ����{��m�@     <�w4��5ds��{d�˜�J5t];���Y�_o&
kJ�9��3ķ�.�6�v��� ���6�NR�ՈM���s�N�ɻu�ꀤd��&ҖR^�7Yvs���t�Ҵ�`0�2����*Ȥۆ���m�N�\��0��ü����ς+E��{����X�Mq)h��6Δ�� ޶���Jd��*L�+�Kʱ��l���d��Ծ&�MP!��Z ^6�k`\�@z�EX$E$*T��5�/7[�J���"?Vk��WW�$S*RL���:P���{z�O�'߾��uhnYʋ�[����C�����i�ߟ��L�&T�I;$���M��5��| � �t߿6�w�L�R	*�m`�>�� � ��8!�O���RN}��ԓ�� �z⊡T��	P�����g艜�({ :z�"�R`{�[�J;P��'ݝ����B��T��I�s��G�����lvk`n洒IH�P��*%Q��Ԣ&��k�#%v�"]�R��/��ST`z�B��`{s[�J]��*WԨUICۚ��K�����R�VDL�emt(��
�'$���$�}.~O�� (#!�(H�HED�0���7�+���l]gL�4���&i0菾���@zoe �_��������L�R	*���PG�7��y�.t�o��v/ڪ�u2��JxY	T�$����OTOhM�]��{�_}UBR��T���́��l�?DB�s�Of�R�P��PJLvk}� BG��79��5�}U�d����`�l9a&蓳�.k%��Y�}TI߽�Q&��\�l�A3D� ���K�o���I7���IbCb@�g�B j�(�٬,*\&�R��&�z���@���	=?Is�,�����m�d��,��k�nPr�p�������Y����0/s[�JK��"!�{����32��s&e:$��_ >!#s�,����`{�k���47�2H$�9Ҁwx����"f�o6O�z���JTR
�,vs`{s[�J�#�~��ͪ�0�TL�%&�5�.t�c�]�TI�1F�@ 9���"�
�~6yi��̭xT/9�N��@b2��$տ���	E�K"ٟ^�ݲ�Qr�$�ɝ�!�(y�"��Б�$$#�t%�$���T�b�X��# �#Ȓ�"RH�X�@ d0�BN��I}{��6� -�                                 ��s���M'Wb��!�mԼ�t��s�1;q�<Μ��m���U�6�F�˱�UJ�]���N��wH�M 6
�3*��ưD����TI�ݹm̭1��
���AJS��ĝ�n^��l�4qo&nSf��ًy�l[V�R��(���իb]���k��v��[y����6�*47��l�j��.iݭ�M�v]����kn���V�;�+cFs�>���0!�̽��=;y��红����:rb D�]�V�p=�Č+�d�Y�YFՋ��9�t;��[�,�
CcV��G+\��9*X@����Ň�M@uκ�ɗ���h��^�N�3/&�I���7\���څK���b��"�M��]=j	�z4r\ѵk�m�6�6�C1�8�r��v#u���]�����kV�%N�k�ܭGRe�5�� J�+��r���KUF����-�gc�������>��[ka�<�<q�D.�f��:�]>t�A7VR�v�쮳WoaL뵡��L�;I�`�s�e��<���=Cam!V�F�(uĪ�W�<��n���vA��V/n�@
Z:1<���fw.x�@�K8J�(	{D�ۧ�`�ܒ�i� ����Ϟy�y�~y��8���$f2b�D��,� ��CHlȟ%����,F��B �K��Z���>}��d��     ��v"/X��β2.�명g�l����e�{v���s���{qB:�pf�:�Nn�:�hŸ6�Գ�l��I/OE�`쑜�v�9aI���Z�d�yɻ9t�����˯6�;1���՜�z���]�L���o" E���f��l5-�k�D�8���ws�Di�r��n��w�zJ�+�>�>OIu�2Mvz�>;���$��0�O�R*j)^�@<�lnk`\�_�|F��\T�M�b�;���$�oUrx�K�a�n����d)a���s�����W�3�}��`fV���ҒT�3I�s��!�`{���5��{��+��\�U��]vʣ`�Mx;un���7����2H$�<��@;�l���>�䝟I�Y�)Kr�g�B�9�}UI�!�b�&�>���I>�K�f�����ʪR�TL�%&�5�.t�����P��g6��
T
iB�I0��� ������D���0/�Eu(	HSQH`z�B�#�no���a=߳I=z�߰2�cM�n�Y2�by�k��{PEg��ub�QH�_$R�J�����Ο� | �M�0�;�y|�B�M�&�ު�&Nϊ$���^�U}&Nj�fe92�L�tI��D�X�8�`H�����"��k)s`]��f�d*�IT0��&�\ =���}��~��'+��W�5R���)%Cݜ����{�f�={rI��A�Y���6A�3q�M��kd��]s�(�I��I�XR���}�TI��N� ޶��
T�
j*�`\�]L�ء��lvk`^�iM!ME!��������N��QVT��R�U:"o;����l��ɉ�B�� �b��62͙TI��T�m�xux�R>�I]��WVA��P�$��f�N�v� �q�;��/!OrI$�j6�e-�ɷ;67Z���v�jM�7M��1�m�x��ݍ���lXf�d*�IT0=z�tDD���l�����@?W�&�R��$�`{w[�5�=:Q%��;=��r����:'�;��0.x��B�c`���𒊚����(�����l���q���|�>}�ߛl      nZ�6�i	'i�Z*�9�4lV�=�p8�u�/3����{c�",�.��NNv�u$�����O$�!�ۮ�ѩC��p8�^W�a�����OO<D&:ͣ�whˍ�ڶ�ݜ��s:��cd*��X%�v'l:쭹���y���ߝ맯�S8��#�:�k���;�Ɉ��H�<&lђuȻ�|�~|��׼����lN��QVT�IJ�T0=���D}2_w6�v�d}�DL�eut(�T$�`_w6�J.>���(���齙��
	�@9oT �6�u�=a�ɐ�PL��P�~�ln�`d�@���%	QSJ��?{�}����`8�ë9�N[	�6.Ԯȶ��I����R��N���w�2OO��NX2+/5$߾�ZâA ����hT֥�I��&����&I��.L)A$�<P�� ������{���5	��}��k��5�/�['Jݨ�)Q	)T�����l��D��(�Yl2O�#��m��婤��q�hz�����)7n�:�euN�~I>~��`d�@;���`]�l�Ҙ%L�T�:WG�'�� =}́}��DDɸ�fd�A%P�������ꊊ#�# ��ڡ����jI�����U)J�B�T0={��{��:P�����T�J���0/w['Jߔ �[�`�ԒJ�f�
y� u�]��g��wnSqB)#�N3\�y���ԓ��(~P�~�l�����F�	*R��tDD���l����Ҁwj*�T�SP�����`d�@;��n�M0�J���u�2t�&��2JG��,"+
?�m;�NbސZs �3):$��D;ｖ���l���0�ԒJ���r�&�n��29�Fv�ƞcf�5F�m�m������l�(����J�EI*�����l�(~P���ʪS
%DʂR`^�Δ�(@k���'wx6�-0�ۢ}"ux�Oe�@>�l7��s�����]4������(@<�l����Ҁ����!	$"���r�����    
�n�<�FM�:���7c�N�qFd��4z�;Z�]d�tg��r\\y��Ev���b����Z@n2�Ba۲6NٺY��㵞�`\vQ�7F'+vƭ�1���nL-��pT=tH���E�[��D����ww��wsݻ���_����8I¸5���1����g:��sȦ%)�a2S�Դ�$�oUs���\��)e�@z�y
h���URL���DL�<P�P�}|��ḓ�0*S0M5I��� �����u�/5�̉
&j��(@;�l��ã���wW�5R��J�����l����Ҁw�0n�I%
T*笐痋��<
����q%�w~���z�*J�])�$����:P�� �����J((���3RNW���$�H�Ԅ�IN��?o���s�{��Z�_n��Ul�
*R�� ���g;��2x�ڊ�H��U)�`{���u�.t��}��뭮�4L�Դ��N{z���@� ���5��$׳�D���>���a�%�܆$�ne�8���u�p����_L~���)��*f������B����}�����7�ʪ%
&j��/�'�5�3���J��q5R��J̱D���M��Q��D A"��-@��f�`E�!��7Vշ>(�<M���i�I(0a!(�@�BHF)	 @c)�J$H!)�+2�`hHD&ٲ�-ͦ&��le[��1�l�2�#%�%�,�p�je,��p�j�l��J�D!Q!�f�����'+,�cr-�]1(%����d%mh�d��� ȱ)$����Ԥ+\���H�����%1�D%d+�	���X\�7
�Ś�z��6�-{E�i���m#	b
F*����G ����~���mT_�O�8�����F� &�$����٩$ԙaK[�~����'�;P�}|�^j$����&Δ}��8`{��ݛ�ԓ�ߟ} �̍7J�u�6�����6��tj�+��gc$��T$(�0=z� ��=���s� ��U��%R�Unk}�}2_o6O�(@?V�B�&a*�T��5�.t����P��g6w9�*S0M3I�s� ��o[� ���K���i�)�^}sRM�w�UVT�L�n(A���/s[�J6���b����3^y��[��e��>W�����~y���)P�)%G���l����ҀN� 6v�T���A)0=���}2d�@?b����G�2��
�QSQT�'�;P��L��~l����ꭚAE!J�Cת/ۚ�~���D��7���Xe�-�o��������ܓ��rL�0�&�#�͑*���Hء�F�++�n������   ��]� }l�A�,7iZ\�)��!�\�]s���e�t�9��Uv��.�lWl����	�g#=�n*�MX�񁸆x5�&y�.Krvc��SƐ6�L<e��j�<�V�ԁ7G^'�,���pOn]�G���û��ww���UQVg`Y�\������놳�)������w|Μ)�f�UI`�́s� �Y����{���T�`�SU)0.t��o[ۚ�D~����;�S(Q3T03k��wx������l�(]थ�a�%ʚ'DD|߽�Q'~����ҀR�P;yUU*fTT�%&�5�:2�@9�J��`���J��+�ҙ.ܜU�˻�z#N:����U����\�@)w(����������]4��y2����n��e�BQE,�2JJ[����$�X�ԃ+D�E��w7��$�f�Δ�QV
�J�T�=�����l�(.� �Y[
J�R��a�}��Oub��`z�6EJf	�5R��J�>��ݜ���Q'4l�m�ٙ)1)Ĺ�R�zqCcc���n��1���pԒ�"�
T���ֈw����l�(�\:�JT*Q"����lnk`\�@'V 6v�T̨�PJL&���ԓ���g�$a ��ň�nְ�9y�D�����e�2�M�:P	ڄ������V���)QH`z�B������_o6ΚI�M��N�M�o(���nz�;/cUn:퍫�H!"�	Cۚ�����ҀN� �+aHW�)UI0=���s� ��@=�l]fȩL��*e&Δv� ���=����f�TԡB��h�y�2MfmQ&�z�� z�
 (	po	e�(�ID�UbP��  ��D���IKr�LI�(�{��$�oUrx�K�a�|"�ʹg]��6�'�����V�Y\�E�.6ڭ��)�$�����J;P�{z�^�D)�L�U$��ҀN� ޶�5���>���3��j*h���@^r�����`\�@+�`�	�J�����Δv����R�JURLn�`\�@7jo[DQ?DG�a-H�" w���.��33333     ܽnZtY؜����mX�%��A�%x]���y�:�;�r�.�C'i1��Z��٬�1v�=3l\9z .�B��u�X�^��8m�s�.u��!m�1.��f�,�����Y�t�j���ҭ���T27N��(��{���y;��IC9�����$�Y;I�@�|��kRl��mi�b�J��2t�������l�4r��
T����w����l�+� ������,4ęb�;���$�wU�	��I��'��Ԓ�K
\��� > -�ﲉ=?I��&��̀e�TB�D�E$�:Pڄ�������[�$�	M(Jf���:�Wm���;�Ɉ��L$WG�&��R��x�P�yx�����Ҁwj*�")P�2M��R�� ` @1B L�vUrx�ڄ�ml)
�%*�&�u�.x��f�Xd�����x��4�I��ʤç+����́��l�4r�j�J�h`]������Έ��&���a�SNe����T()���1峪:�[A��*�T�P*Q$�X��6�u�.t�������
*T�)0=���s� ݨ@=�l/uJ�Ғj�$�}.I�s�[>�BJWĩW�ZF� "�DJ�R ��Y{������lf-SHP���ã�3� .�[ݺ�:P�EX$BE*���`w�_w{�t�@7j??��[t�(��P6<�8�"zMZ�s�n�tb�IH�&�u�6t��{u�7�O��2��ӢOO�2n��I��lv�}�}2gÕ5T�USC3� =����f�w6O��R��U(�j}́��l�(1lLL�o�L24Kx�h��I5[�n��$��L�ۺ�:Pڄ��������5�6��-�Ub[V�ݏk�s���ю���3�&�I06t�������ln�SHP�����������l�+�K�QX
�J���}���ڣ����D��a�j�/$�m�I�&�{��O��d}������q�)���*���Ҁ�������~�Z�c�1���˚:B6��@uh.`q���|P�Q���� �!D�U�,� r�E@���T:0�؉��4Z��B¬�6o{�2̂Q���X���vU>
J�,��Z�*�0��54BW �e�eh�6�e,*1�Zd&bc[̺,�HXAl����p�DH��"Nr ¹��@n��m ��}��
Ε�M�P��h�3�k5��n��� 4��I�G����~����m �                                 	,�����i�O2��[IZ��7O6�i�"���з����(hw]4�v�F�Y��nY��n$`m�]�����↌![�j�csg����Au��i'�*��:�nz���u��e�L�oJ��q�,ۧN�٣\��ۇ@���m�uԁ8�AN3�s��Vc�!���5�!���l�s���gq҉����Fz�ضd�3���%����cŹXu�[n��Ő �v�wI���h�;&�n؃`n��	�fۂ����S���l��5u\�Y�"q
f@��gF[*ʴf�'�#�xԺ���1�؊���� Nim�ލ"uv�]��On��c�\݆�9�Ѷqsv�^z��#g
���g�u��\���r�\�@N̒�k�-H�q�LlZu[Q��leM���J��Hgp�٦ڀ)bl�ʖ	����4;$KRd.�]�E�c�჎:81����=.�e�4�[r:JҮ�J��n-�u��JZvɑ4l�������2�1��8}l��Mg�V��[D��d�۪�Z�����$F�s��M�:��
�m^YS��E�պ�n����-ϛdܒW.x�#JE��E�r꽸	���!�vR~}����;Ώ�qz��B8� �<~Gh!�A�)E�
$b� �&��h@��o���'T��^��|���_����     qf�֖�.��2L�^ �g��p��LM�:}eڻ�����Fܑ���c�g���^�vv*mv�e��G�u�8r ���rG�Y�A��eaK%b�=��W�pv��}b��� ��]�Tn;v��y��<��<��OO@q�e��rM>2�dĹ�g��ZGK��"��+k��'���@wx���ސ��~��T�(�J&�����lf�`\�@z]�铧�j���*I���́s���n}���g6���Q
iI5
R`\�@z]���a�o������i*R7�����7����.t�:>���%Uc�t��+�]�j�\b͞pl�Dp�9�7��y_��i��NT��N�憎7��D��? 9&��Y&�r�rJ�ܴ��M�����E0DH��;_K�r��d�\�u��T�kN�Jd*��R`d�@9w(�́��l�4r���*�h`\����`{w[���(w��%�D�P��g6�����'��P�sv%U�qus�H���BdsѼ/]Y�����W�]mB�$�^���.t����r���7��$B�RM@�`\�@7jo[ۺ���d���i*R���k��"��Y�J Hu YNOI���*R%?D}7��`_w6Δv� �Y[
B�IJ�I���l�(�B��`m��$���)"H�"�T5����cV�%�Nwi��!�c�Jd&��T�Ov� ���=����f�T�R%UM�P�DD&�z������9<Q%�चlJ�MCۚ�����Ҁw�����@�J�e&��`\�@;�M ʐ� i�oY�sRI���fL�iL��`\�@7jo[ۺ�'߿>�W����K�o]6��{Q�]�%{<��d���HQH`]�������O�VD$R�(`{��ۺ�:Pڅ�2z�k�HWԐ��`_w6Δv� ���=u�¥2JU*L�(�B��a��՟�~�q߇*j����ި@~�fo��s`rx�K��@� 7���Km��m�    s��w&:�0�<k�ܷH�S"6UY][�;�K�<�ܲm�ջ;�l�ˤ8���yݙ{��M�Qt
1�f��4;\:��u�g�vl�p���[����q�c+��='��G�-Eɮ�\1�չ�ЗR��F��;��<�;�ҽ�/^]���Xҝ����^W�r�uY�s��l�]�d�=�����l�?�R�(@t�mB
T�)0=ۭ�s� ݨ@=�o���"&C{�$E(�3TJI��� ݨG�~�́}���Z��"�!E!�w�/ٺ�wӕ�y�+"*SJ����l����Ҁ�����";�ߟ����K�aH�<���PTr�a���oP�Ѳ��i7d��z����nk'�>�D���Q'yx�s �r�N�9<P 0D(B+�H$i"�2��~�������~�lf�`f��5T�USC&�P�?}�D��s`d�@'�I%
�J���9�=���s��w(�����
��������Ҁ�ߥ �����I%	}))����v��ׇ�y�<�&.�玷U�0N��v�z�{�f�~M�Po[�u�=��MB�T$(�02w% ��/7[�J�j*� 0Ӕ��&�z����TX���$� �i ���
T���i�@��3�==��5k�C�T&�I��k`\�@zoҀ{z�u��B�P�M&Δ��(���y��O;�}�����u��F��X8��	ծlg�����*�h`d����`{7[�J?\8�I(T�T԰=���L���:P��L�=yEP�BU32����.t�=.� �����D%�f�M:$��D���d���ri����z���{�T�T$(�02oe ��=���s� ��]��T���%E@W��KA���;�0Un:�f���aL!B�5*|��`{;��9<~�!�97��7����T&�I��9�.t�=>�@=�o�L���B�3�*I&O��(�́��l��2���J��~���v����lfsa�r��=��I%�
jX����f�Δ��(>��s>��I      ��i;8�^/-��,�stʖ��I鶷"��8t>I�)k�����N�d��=8͵��Z�
]����{$���u��ͮ�d�F�.�����9��&P�r��tA���n;�|�]:���y���/i�9��=������q������Uuq�]��(�W	�#��n#�]x�.��s
TU%S3)X�́s�����Ţs����}��&�&(9N�9<Q'�ܠ޶�u��}��}��HP�a3D����MnmQ��-��Uz~(�y����C9R�7������B��û���*r�t/w�| �#~�����|Ńkm�Km��(�T���;gl��[>ٶ�&M�Ҋ�Xĩ!4�q}�Y��}��fs��;�V]�䕕uz;;�.�H
�R� ����`��9��w�ȿrW���lK`�S��Vf���,�Lu�j)K���C�#舁�����,�L?��٩6����܅�ɇ��Vv��"0`>��m�[M��Ye��=Lm�G<�� Z��;Ce| �i�2�r�e��x��sX��\_r��XJp�NT����+7\_rk'� Efr�rJ�ܴ��y��-Q�#6�m~G�ҋ��.ٔ�
�%�"FA�"E3HS�wZ7%B�C�:�
5F�n�h8EVg4��2���2�D��H�*�R$mSbA�K2J5���!8#�!}.����Mj�P(��a��I�}l!3@n5xklh��C!@^q%JT�6J����M���$��H�$E�_ �mA؃`���o��%��R�i�+������\�s �M4�_rk&g1��uFn��e�,�r�Pӝ0�5���ܡ��m��s6.l���v����l�c�(�s�XNٛ��u:%L_��Vn��w�DCof=��E"�a�32�^����3�C���y�{6SrlL��8��,�L>�b���no3,�Pl�y���S��p�>����O�}�vb%q)�9R�+w���"���=�?'�w������R��v����$<�8Ⱎ�Fɮ��\f�̴�4��t/{�_rk&g1W8x4�A��i����p��W��V{_DD�3w�3-)d˕*��������8�yW���l4ĹS����/�5�}�I�,)s2�^�8�{�a��~�a�`�L�թ#"H�b@��:���     UO@��z�E�v����σ�������ɴq��t�2[&kksu�P^��v�L[I��L����iۦ���[p��k9cg4�N��u��Ax��^�e�ûp=n��۔�H�~��	(A�{m7%��w�����}�v����M%�Z�GU���@7\n��ū����4�NS,�ؙa�q��,�L=�1Y��7��K(6XN��釹�Vv���/1��ᆜ�s��Vn���,�L;�\HP�R��w�Q��k&��U�9�d&�n/�5�����q�{������r�gU<�k�.rZ�ܷRk��i�R؆U9�3X��~��#=�(^ha$�I��t���q58�9��=��nk��d�BN\�$�B����!f�a����l"�be�)� ��a��w�1Y�q{���%�˖��:a�k��3���/]EK��k/:iq�qf�86{V�k��9�P-�-�nT����+7\gw�@c��fyx8����t/}��@o��ه~�� �N�2S�m7�!g.G�8�C�)������9�{o��Ue�d���P�����+;���8�r*�0���-)���/3\grs&=׀Ϲ��\�W^� 'g0pnWsѼ��Q�8��t˝�l�5���~����,�L;�q��-�lL��q���û1Y�1y�} ����0�e�	��ޘw��fy�w!yh�����R�z!&��a���y��@Hb��B1���ӽ����K����܅�ɇ}�u���m��*[d>4VY���v�g	�[@0�vݧF���$�z��~���������q���2ҖL�R�iޘw��fs��B�^�)�.T�gs��x w�Clǽ��	9rT�����B��D�y���[E�ؙa��=�xFNlƹ�a�s����!P$�0"$쿽���     �����Y���K4Ĥ��ɝ@vl��TvN�ti�Cp��6_��Mnv��5O]=aD�*�{3���;Y$t�i�I�y��z؁pY����6ԩv�K���"- :F�t.͑�Ʌ͌`����D����������:hG��c�8�'b�z���m����M%$Ð�-�,'��>�w��f|� 7�C6p����R�+=�� ���!f�a��y�$(l����܅�ɇ}�U�d�2$&�n3�7�����q���2ҖfYR�iޘw��gk�ﻞ���`$�I9�����v%h�'ks���=�hϮ��a�L*b�����܅�Ɏ�ЈI˒���^�;`T@� E��`P��,�L;�~�o���Y-��N7�B��ÿy������a6��<a�ky�xD��͜il��h�f+=�*�\grs�=:ϻ�m��3-7()3)c,��vv�ȣ��+.��0�')���P�M���܅���+9
��̔�D��m���w8a�s��2�zfZR��*U���]@� � H-�By�����w���@����Vn���=-i�{gx"rXR[T/}�<7�c.tÿy���m��e2W�p�ݹ8hׅKs���&.�玷U���:�Zy���ߞ������q{���a�˖��<a�k��3�x l�+KD&�EK1{�1Y��=�]Nw|��3*)�B���w!u8G��q���c.t���Ȑ�I��rS��1Y��,d�6�lȖ�ē]�ui�P�
k�ɣ7\�AP��T�f\�fe�*���{�Vv� ��������@������3����9���ڡ{��;���0���l��ؙbZq��]�w��^s���C�\����7X��q]�L)(ı�s�� a��A=#��[4fp �'��\�{*�p�Y�u��y��D�'��F	"V�4Fb�kZ�#p�$ vF0LՐefH� �����wT�Y��3Dt����{��[
Rޒ�8Uf��z�ϴ�	3f�?wD�r9�
�0�UɺC�0��) �w�E�{���|k� A�
��/
0�Qb��D�����Z�I�I) ����?!�
���PԪH9 �$ `j%���m��[` �`     �z                          ��^�;&��iWT���7����K*��G�z�:�mF�2l�$(}�S�h�d$�j��m@7t�;j��Ҭ��JD�Egz�N�6�*Ƶ:-s�g���gj���v�Z��ݹ]�sH����-/���][\;����'ժ���8E�����yR��*G5ۚ�6�^'��z����j�v�u���9���gHb��S�!q�$6���%�����v�5��u�2�<8��6ϒ9`M�A�1�85��.�`�;��z�Z�j��F�8v]�V�T�Ncby����� �}%�)����Q�R����*��d5�I3��W9�5����'8:yPI��6��C۔��w�Nݹ��k�'S����vݮT@�F���U�X��b䉷���W��/��S�5���C�8�Fڭ�����V�UU��-�h�s��n�G����R� ����E�]��eV۴�Z3O�^�G^\A���)�\��fzg��������V��iL�x���y����N�t���ݛF��-�L��#����n�[=p�mҐ�[^��:y��Y��� W] �k6ڈB�cۥ��/� A7��G�+v;tVGv���P-����ۤ���SM�8m��j���e
�'���j@�*D�Z!�5��P7b|���m�v)�`.�#b�ztFy��w�����m�      9��f���ZM&�ck�:�~�$ܳJl8${7\)��q�6x�؂w!����ك���T-'MZ�=�'e�*��ŉS����<�Ѯ����ܱ��Ѫ�^�Ct�\�L��,nsjݺ�
�p�:r�����:�����4��\�	�&�g�����9܉�������d�Z!6�*Y��y����B�p�|�����y�⻐��0���ogO�)̉	�ۋ����#`�������*Y�eJ��<a��y�+�
xR�)�h�wsy�+�
���߳�πq�u��t�:�^m�\�v��qc�/��Z�W$$䰤�t/7�Wrs�v��͖�fXe�:���HB>
c
(4H#� ����1��b�<�#{{���-�,'Cz|a��y�܅��8�E�EK#� ~����q^�=�i��^peCE$�^o�Wrs�v���kmձD���ф���k�5<��j�5�3�rZ�`㪤⻐��0���������eʖfYR�^�  D]�����{���b�CJU��q�}�5�w�?;	B������~�#�0=�;�����n	 ��ߵ�$D�i�I�/��I\��5�I�w��0�*�˼В	"w޴�$�o�قH$��{ؚ�H&��kBH$�Ӥ����N��Q.W������w]Ӧ�:\�^�5·U"�4��H'~�LA$Ms�bj	 ��}�	 �'}�L�H';|��V33.]dВ	"o��&��	�}��$�H���2	 ���`�	"h�=~�U�r�3I�$�s���$�H���2	 ���`�	"k��&��	��g�Kʢ����В	"w޴�$�k�قH$��{ؚ�H:Q��IJ�Gx'�pf�ϴ$�H����U�u��%��7�N}~�$�H���bj	 ��ք�I���A�;Ξ�� �H�st���K9ft�%��8�����^ά2��x̹�$D�}�MA$w�hI�;�ZdA5���$D��]��r��S2���H'=�����j	"}���A$|��	 �&���&��	9��VfC«	��A$N�֙�M��0I�1j&���&��	����$�H���0��ɕ��pI�o��I\�ؚ�H&���В	"w޴�$�o����V9��uY4$�H�ｉ�$�o�ք�I���A${��A$M��6F")���������   ��������&۬.8�G�J{S��sǗkur�uαq��܃���Y��J;<ݹ�:�f�{-��:Q7I�����d�zrWhg�vm�s��i��̵֦۵cW��n�nb7����\�����A�V��A���F�DD�A�V�m�2��U��(�Q�s�;&�V9�ܛ�k�}9����;��w����ք�I���A${��A$Ms���A7���IyTQy�y�A$N�֙�BPM���$�H���ؚ�H&�w�hO-P�'����*�%VK��n	 ���LA$Ms�5�M���В	"w޴�$�l�:j����	�4$�H�ｉ�$�o���	 �'}�L�H���g��I���E�aImT""}ު		N�֙�Mn�0I�5�{PI;�������4`ξm�[�ۄ�yC\nܼb�ںv�3%efC«	Y�A$N�֙�Mn�0I�5�{PI߻��$�H���ؗ-�-�P,�����X��r	"w_kPI���$�H�}�L�H&�}�eˬs/.L�A$N����A7���	#���߭2	 ���� �&����*�+/4��H'?}�ZA$N�֙�M�e� �&o���A7��{$��.�e�f��I���A$_���,I�5�߱5�M���hI�?}=��333O%Cӽ�T�v�N�6���cX��-�	`�?&��	���$D�����H&��kBH$��z� �	��髻�+����I}��5�M�ߵ�$D�i�I�l�$D��\�r�2�e�7�N{�kBH$��z� ��B��@�b��`�	`���e� �&��bj	 ��{�ɒ^XL�В	"w޴�$�k�X�	"f��MA$�)��{zA$N���Lʙ3&V�M�$��ĐI7��j	 ���ք�I���A$����@-�VT�K6�c^�%Ȇ$��=�G5���(Leˬs/.eA$M����A7߾ք�I����	�$�M�V$�H�9���U�V^i7�N~�����H�D���L�H$��bH$����PI�/��IyTU�˼�	 �'}�L�H$�jĐI7�bj	 ��}�	 �'y�x���%VK��n	'�U�}��I�5Ͼ��A7����$C� �!���� �0/�P	({>�H4[�4 $����&��	���ZA$N�֙D[(@$@&޼~��l6ږ�^]��8Y���D�n'<Yt�;#�\�6��Xo�;��:A;���hI�;�ZdA&�V$�߼�Q	g���%�2�iЀ`�'}�L�H$�jĐI7�bj	 ���ք�U	"w���fTə2���n	 ���ĐI7��j	 ����hI�;�ZdA7��k.]c�yrdВ	"o��&��	���hI�;�Zd@��_�ĐIG?v�c
�
��&��	��~ք�I��~��A9_KA$L��ؚ�H$�C��$G�� ~/���{     ȫ�Eҩ�:*ܖ��,Nyy+���L^�	���bq�.ƒ#���ڎ���WE2�Wr�6Q 6���e�Z��q�z^݉���9��<���­r���8�^�V
v*��[#>�fz�sȝu�)� |�6 &�m��je�C\�4�k�{u� :��������2�)̉E����H�L�r��I�nĐI7�{PI߻�hI�;���VU�J��W��A;�$D�����H&��kBH$��z� �	��髻�2�J�	 �&��bj	 ���kBH$��z� �	�݉ �'���K�uXa�3/I�$�s�{ZA$N�֙�M��I�TMs��MA${��32d��V�4$�H���L�H&�v$�H��{PBD���@$@& voy��r�4�R�i��;r��|=����sog��2�j5�E���w����w�o���s�'��'}�L�H&�}�]��7��2�$�H�ｉ�t@�FO�4#� 	�7�{��$�H��2	 ����5BH�9���++/4��H'{��$�H���2	 ���A$L߽��$�o���IyTU�e�f��I���A$u�bH$����5�?A��oBH$��~���ʺ�U�����H'k�ĐI��>�pI��kBH$���P	/K��m���Hp� ��Ќݝ�g��{L<�g�0��WWFTɗ4$�H�ｉ�$�o���	 �'}���A9_K� �}��Je���@�  g��hI�;�ZdA7]�$�H��{PI�s�K̬�0��Vf��I���A$u�bH�:'�U>'�t�t#G,n$��o��2(lβ����T�P�$������Ba����,	(S`����Z-%ݠIfs5�fr@�)I�X�0��4��ul�!��hQ7p���v{�w�bA"a�՘J��C%b��
/2�,J��'ȴD�O���xЍ�e�B����(�0ډ��c�D�넵S��l/�ol�������t�<*|'ª� G�/��T�)/e&q2j�Q:����=��  �TS8A9�GJ��>]���kPI��}�	 �'>��+2�Lɕ��pI?D>��ĐI\�ؚ�H&�w��$�xTO�~��$�o��컫�o/*L�A$M���MA$}��В	"w޴�$�n�,I�>��{ULS�K�a+\��� pf��u�h���nj�^���I�$�s�{ZA$N�֙�M�e���PI\��PI�o��IyTU�e�f��I��i�I�vX�	"f��MA$~ﵡ?U	"}߿~*���Ud��&��	�~�$�H���PI���ք�I���A$g9�Ut]S&\В	"o��&��	����$�H���2	 C�4J �}!,@�"�@��U2(7(��S�����bH$��_W�.]�\�*f^�pI��kBH$��z� �	��$Dw�8DD�����n%'%J���7nNZn��nv�]�$c��%��u2b�:�J~w�'y�y�~��$�n�,I�3�`~�� g��P�H�L�{�,��e�	�"H'k���1�$��w�MA$����	 �'z� �	��{�uyp���2hI�7�{PI�{��$�H���2	 ���A$L7�{1��³3I�$��!����	 �'߿ZdA7]�$�H��߱5�M����/*�����В	"w޴�$�n�,I�3~�&��	�w�В	"Z/�~H, ��a߽����������    �:u��H���.w)u�ã�]���]���/�i4�/�����[�I�ę�^wl��'k	Hj�`��J��\��]n}u�W�xl�n�7h�a:��溵mJ�:xšLmnK�Ӈ\VR�۩�K®fV\̺����/ E�=��⪬N+�l�\s����ح��u���WY*�]_S�$�r�,I�3|�&��	�����PI�߭2	 �;ߍU�teL�sBH$������$�o���	 �'}�L�H&���P�'�v��r��S+4��H'{��$�H���2	 ���A$L߽��$�O��fL�0��Vf��I���A$u�bH$����5�M��ք�Iw��̓,��n	 ��KA$L�;��$�o���$�H���DDV�m��MKmL���1�M�gӝɞ
�Lmv[)��JSD&��������
�H&�ߵ�$D�޴�$�n�,I�5���1��³3I�$�s�{ZZ|� �D#!B`A!� |�%��w�3ܴ�$�v�,I�5����$�o���IyTU�e�f��I�z� �	��$D���MA$~ﵡ$D�{�YWY*�]ޓpI�zX�	"k|�&��	�w�В	"w�ZdA6s�5WEѕ2e�	 �';�bj	 ���kBH$�߽i�I�vX�	"~���~ʫ��T<>7ŗ�ԋ㍸�$/H\D�%s��tL��r	 ����В	"w�ZdA7]�$�H�߽��$�O���2L«	Y�A$N��L�H&�ĐI[��5�M��kBH$�ϻ��̨fdʳ3I�$�r�,I�5��P���R�E�@�6#b 5�߹�	 �'?}i�I�V�JSD&�������
""�ﵡ$D�޴�$�j�,I�5���1��³3I�$�s���$�H~#��Zj	 ���� �&���&����{���� IK�O-�ۯ��=�`�'�� -ԙ�ܙ-�%�QW����A$N��L�H&��ĐI[��5�M��kBH$���ުʺ�Ed��&��	���$D���MA$~��В	"w�ZdA4s�5wE�ee�	 �';�bj	 ��ﵡ$D�޴�$�j�,I�>��.U�T�*ef�pI��hI�;��2	 ���D)GdI�T�"�ʢ�����A'��̙&aU���	 �'~��A$_�Gw��dD�=�PI���kB		��Á��m�[M��Br����m��)w����m���yUxLʆfL�36��H'k��$D���MA$�}��H5�>��L�H'>��˗yP���2hI�9�~��A7߾ք�I�z� �	��? �	"o���+.�I�$�w���В	"w�Zd�,*	��X�	"o��bj	 ���~�/*�����В�D�߭2	 ���� �&���&��	�߾ք�I��U�u���wzM�$��bH$��󸚂H&�ﵡ$D�޴�$�l��#�Hmc,���M�V�333333     �.�{8�^��.@���#�L*�/��\������gV��R������e��kV��xxθ'�N����[����Ǳ[[�"�^K*�6]�L5�U//j�ݱ�����]-WJb���r]�˕Yd�
�,���P� &n�m��$$�B�*�"H�����5�3��[����xe�fI��>A$O���&��	���ZA$N��� �	��$D�ۮt�WYS���M�$����$D�޴�$�j�,I�5�{PI�s�/2�L«	��A$N��L�H&��ĐI[��5�M��kBH$������*fdʳ3I�$�r�,I�5��PI߽��$�H��֙�M��ܫ���ʓ&��I���5�M�ﵡ$D�޴�$�T�B"0?e��6�l�m	i��_Y��8�n����V�2$�ACᄜ���@$@߾��@&��tïy����Js"[�-8�~��t,�=A�����P��N�NT��^�^�q�9者��QXRT,�W�Wv�����ґ!�\�b�����8cz��#*\��.��s��A�0빊 �km��I�,He�`�5S��]q�t�WU�����;���3�>�OsǮ�+�\V��-Ķʔ�g�:�b���o!Y9�),2�rK1y��f��A�Ph+�������k۲ޕ�	6�_��3ypî�*�O2S�ܹi�o �u��wk���w�m�Z
[c�;��P���!��@��=v�=��X!,qe�o���c�k��A��)%�F/;���q��3�;�o2��a�mP��q��3�w8��	���e�Zc���tï{W�� .�,I
KH$@_ r�3�x&T�[�g�:�b���o!聻�M�ۙ�E�,�3! d�I�* �Z�pg���c�-���nT�M�%������q��D(銿b
<%�I�B��~#{�Q���o'��)̉n\��{�3�{�Wv����*Y�,��z"2|b�u����o�b�JD��rы��;�"3���zB6c����$ҕ\j�UUUQ$"֟�$�$x�Oh���˒I$f�߶y�i��O+-2ipN�"��*?�����
�
#�($������� "��DDJ �HFt>�V$a|\|�(�eSg�߽��{3���e���YW���N��u\��~���s&'%3jZaf3"G�4mk��vI��$#ꦲD��uȫ6�����w��M��΍ܛ:A�I �<�ܧ��J�0,�X9�_�cY�L�%�b_�c�q����=-*l�K�?�������(��-Њ�%I�UDZ��BI!؊����)��p�+�,����C���2~���$�$mp*�*�[�'��F�^M����m�7C��+���<J�H"G5��0x�~_�s����s�i��H����/���>|�����9��$#l�:���s�W���ٮ�k�R{���!:;�H"G�����sd�T��)RuY��7^MU$�\y�"�pQM-'��̑�e)y��bl˄[SC���?��hv����I �=�jo� ��y�I��n�����?�4�|�I;g,�OV��맶I�<����Z$�$w�xI<� ��}��n��s���u�ܙ�,�wv��R�WWe;G_Mڲ�G��X�}[�H"Gqs.-�k��׽ɼ��+L��&H�b&�ޒA?�Q�]�]�Bޮ�RH"G)�˺:-a�3�82ҌN4�Jx�#�J���f���H�
�� 