BZh91AY&SY__�*��߀`x����0����a��      	 }�>��(�[ZSf5"�[�ݻ��J\ԫb$�,�� �E	*�P
�P��4dY�'�j*�        R�R�$ U  � ��"�   
   @J�@�P�     fX� :�� P�� W�1z���͒�x� 8�m��2�۪�����t� 8Y�&�   
�jU�i֎ 7v����U��aN�s���3�YQǠ'T���馷0t�[�� �:P �  B�$ (1�� �׭<�Uū�\��zn�uO�zO�|���h�����j��e� Gt����:��۽|���u��s\��|���,��U㻊\����j�� ���[����y��ֻ���}��z��o �� )@��� :^�Vۗy���-Uӓ������p>�Oi�k��w��Uͩ[ڬ��� ��[mͻ���sǠ �q�齷�wV׼�����>{ݫŹ���ҽ����{�Р�ҩ���+�n���}n���y����J�    ��
� ��Uź�ۛu��x���y=T�������}�i�kֽ��]9:�����V����m�j�  ��Ҿ����m�����}5snf�-sg��ۼ�W{� s�,[֕ͮf���g�����z: 7Ҁ   %@V0����x�k5ɧ|��jOs���ҦO��ͫѸ����|�����R��֪�k�  μڧ�r�K� z����yy5��x��n,���S�>ۓ���k�����q��    =           ��R�T0 !� ��&����&RR�	�� �&@2'�UJ�S&�L���hѓF#0"{JQ�(@  4 )���T�� ɦ�C  i��`B��I @ ȍ4�ޓjhG��`�����~߻����=/����}{���A}H"��?r��@E\E�����`(������N�PW��>؊*P*�U�2�@�
?�E���d ?��� �Q�<�� _$�$P�E��TaP>�S�D~����@�U>�� >�O�W�U~��T��Q�D�UO�O�A�Oe�O`@�O |�O!@�T}��Te _eDO %<��|�<�<�<����V�~�>�>�>�>������!�_! �C�_��~�2E����O�~��@���>����~�>�>�~��O��>�>�>����ҟH}�)��?@}	�/пA�ҧR=Hu#ԽOR�ҟK����H�J}}(r�!��@��:��N�:��>���}��=�!~���Oe�`=����~����O�>���>������C�O�� ��a=��_a�C�d}��S�O�� d<���|��G�C��`>��
>����S����O`=����S�_a�C��~�~�2U��>�>��P��O�>�>�>� 2C�O�~�>�>��O�O����R��ҟK��*})��@������Ru�'R�=J�K�/��?@�*}JJ�� ������:���>����>��O�~������O�>���_�~���C�P�P>�>��>�����G��C�O�>���_�~���y�s�|��rC�J�����!���?B?J����+�}!�'҉�����/���'���{�HJ?B�"��'�}'҇пH}	��'�dH}҇҇��@?O�JB�JjCR���~��O�~�� ���>��~�>���������>����D>��~����<������/V|!�ӳ��:�ô16b��ə��ʛx�P�]�jM���N;���<���m���X��d��JJij�
���JS�رfc[])BD��rT�B��d�5��ighd�l��ex�V�.s�6�	��RM>oyVM8(��6�=��bl���kX�c�殷�����i�I"�&�Kq�?7)��CWr�ĉ:ʡ
�(T� >*��u��[�u,��'�C�:71c!(�C��M&F��BL��%��y�h��v{ݽo9�98]ft����XK��d%&&C�d��N.��
���錀ѐ���DK���mk�b����.��:�o �'O�=A�7��WA�����-���b%�xF�Q�%������#����I��d�9cF�Yy��83�4%�1�ٖN6Y����dg��y�Ğ�/FB��f��=މ	Y����վ*&��C�մ�A$D����a�"viz���O�8g$gr��p��9�8�S�'������'!H������թ��K�'�-C�H��l�˰���x����|ʑ1[��XB�6�Vˑ�w5>���w�ɜW/��C�A�u��}��Yu6;�ڇX��T��Y
1��:ߛ�`�f	���a���nL�AK�_�8�T��PQp�T,���Y*D/Sġ���K)�i�DU�T4�B��0���nG�Kh��2s�u�5K�H�{D��zv��r�0�J�=7eԏ	�omn9�q�݆�q�u��݅�1��t���R��$�$����2X' �r��<u�e��2�p��%a1	CHC��%L$y�MCy�N1�ŪJ���:�P��)=!���mEZ�3Fڝ^�ɠ��w�P��	���㲔��*�c����"��O겮��}��RAle�oA���ѳN�J7(T�:K�*���N����R�����ݗ�+Y��򉺱�&�=�}�5�}u�C����%�Q�vޞ{��dc÷x��Z�푎��N��,a�8����4l��cĽ�pѳZ��g��.�*JiX�0�;;��1JBV�Xh�3�8�`��8	ݩ�vy֍f�xDlK�e��kvV���=�i���{�I�"=�֮a���:q'�y	a!�.��V��:XA���h���1���S���z�Y-���C��Ē�K-���O/l�J�D��ԩ��s�3����.\�z�u."��U�%�<Ϻ�L�M�o�g�dJ��3��"�>b��(I2�0!�ᙤ�Ĳ#-Y�ɧ�	(�udىԀ�ѓS�ԫ�uO��D��/=�[%Q��B�hu	(��j2g>,��k����D���Bx�@�,�1	���U��*�nQe�y�QQ~�>����FR:$h��

b%
q$��aS	3�����!Bxc��ʺ'_.ȝK�,��J�is�.�	�PJ̈��JEP�ɴ	�Nr����3��e�F���f��8��3�JU�HL������MZ�t�#EHy��C<�U2!L���y�٠�=ђc�Rp�͇o�9�keR�$���'-���֣.b�&�".�AL��q 00!>�l�菩|R+����|���� i�j�Ӎ��T冋VFK6��K+XӐhr\���
5ڵ��D�׸ɱ�pJg!3�<!�X�>��?���/�5
3V�q<Iy����C�x��E*�����(F'ξ���9��DYO�%TꐔT��Y[��� ��إ�㏾X�S�QJ�G��M�M*�����Hc��I}O�_�>>yZ�"$�T��ѻ��)x���'�L�y���X��:��<)t���2�_�"G���>^D�ҴB���/�����z�)?��$g�S�j��V���q̳,�JLc!�����^e�d��_.�i���g#1���%/�I���'���f�/9�h(�x9�͸Hgt�Z'|�P7��i՞OhP8�˨���%��W=S�Zyj��[����8C}�S��c\<����i�ATQ�P��wwTU�~�����oq����B�L����U�B���i��A/uT�L�ba�١ӡ6C�Rɍ���}���[�s�]�;�s��Q�~:�V�q�5�]ov-e� 2t�!:	v�<�o��f�兎H\��Gh"��]&�Pꆩ�M*{x�����ϵ�?Ə��AiDī��M\Y��u*�q]E�e�4hd8�"��b{X�+�]<�û�8�kvh"5f������]����1��@�B��2���7�uc��wN�)�z�e�����%c���A!pBF��w@C���&얔�d�r��޳�yrtfalu	�4k5Ӭ�w�A����s<�k�]����}KT]�(��Y1J��X��&N5��0BƵ�N��R����7��h�5��`�dh���9��;�&��-P�!'�B"UQr�e��]ګaq�����G��B�BC�����((��lʫ3��ͺUDWJT�A>I���~���A3�|ϩ}H_B�*��RǕ8�@Q����Z�U۴5C;@�M�z�)EYR�H��;�'Gĺ�ʝKr��*�uK�B�,�j��l��ؓ̽������u^!�){a�P(h��ٝ����S�z�Z�|�|�%�u}Ӆ��NՎ�U'۷!R���������k=YRv�V<���	�˘o<;c�Q��{�ӫ :�.���+�1�Q*�"�i�O�)�<&�
rlD�S�V�)]5�y)b���6	�&@W���w�b�< �0��#<�茜5�ӆ����`�JL'f���u�ނ��}x7q�a��k���%!�v��OjE`���D"q,uL
&餖����OTMTBW"XE4�S�0���2N����36kWY彻O9�Ӣ�h�jp��Z��Fk'�p�%.��b�xSY��F	<J��8#^q�C.������]Rju&�h�M����jrR&2�������	9H ���ޚ���M剤UV����`���RJD��*��f�'BN'&�L[RAOsN�
�Ny!D�Z�MFMk@���ĳ��xwy٪��lUo1�*��ē��*�j]9�����,5����Y���_r�����2�D��ڜ��8�S:E$��>qfQHU��A��QJ�T"'��i�-�
	�2�s�y�tce�z���U��J�o�w��ZxWW��i���;�P� ���k*,�j��ESۨ�J����QhQ�F2a�j�k*��׃��eJ�7&���^��]�Z�%FA��7�:A��l#F�(p2��%	BP`�X��# �0r���d���rLM�����O1�#6r�)��5l.��VHԸ�ޱ4�N�֡(J6�:�48;�r�����u��2M@��^��P���7��'p�2��Bs0�N�<�s����&���w&�2]��`���BP�`��I�z<d�BX�M�L8Ɂ�o:��#@d&�)4H`<�IBk�Oa9	���a��20b�Ho.�&��y��l��8A��*�ԥC���"Bb�U*��>m�SK�ݭ�O�^&�h5bEޠ�;5f���%�sQ�'����ON�y�Z8�n��t�q�ta��'5�o$n6I�ֱ�V�؆F����d� �ͦ�4����twF���&��BP�>��C#JP�:�����R��zzv����T�bbdbn5:8�����C��d�`�����y���y��S����86Fd��: ߼+q��G�8��d��	I���xn:7�	X���w�:v�d��2�F4����3F�ݏ�A�MXi��xO�gA�Ō�:�����I����J4j�Bk14��� �h�(�c����D��	��=�a����6E����=^�{������&BP9�Cy8o\�3�j4�v���Έ�s�0-DFv�	`�y֓��bd%'I��Pew�X����S.ȉR�دҝX��^QhI�PU��0�)�%#3��5�:�Nkk��;�K-	h1�2�A��e�4��BD�y	btJ ����a�����C��U)�*n��+�V'A��Hdq�'2滷��=��7+�x�D�:C�D� � Ţv�=Nf�íɸ���h��J�1�*�j�g�)�5u���6	A��6:�4�C�=�X��S��a���2��Z`�Cy�t�zw\9��6j�cf�4t�`h#!(Ka(;'P��&�ѕ�I�fv�3���C���2��̃�dK�2e'7�o9ߙ�:ٸ���&��xY��F4��x[Φ'4��45���bj�2YY�e��P���NZNգGp�Ր�`��%�2C�%���f��VᗇY�ۓ�Y8a!�4�0�Z�zf�/࡟�dL�D��2N)f��y�a�k�1��21�)�q:b^;�ՏMަ@�k�3��[2�D�R7������P��vB"�@(�vǘ�2ڕ	�-��)���q$�D���������M%WO�w�GY���	b��A��R�zG�a��sX��id��g:� �Ļ	�Д��i����
�����읓��5��W�R;1��d�S��Xh��p�v�6bc��f	I�=�:���xa�ZsE�n4�xx���1ӨKoK��I��f:�S�ה���V�s#��S���#�n�̿^C�<$8�Y
!'K#���R�h5e���04j0�����ѫa���MBu��'r���&�S��
����D���P��u	���+c�d�f��ѓ5�o��p2��d�����\����I�d�Q�bd���X��Y�t:��&�8��5C�AS5<\��&*�fd�rp�.�yՅް�xun�j�NI�f8�N0e��wsV��oz_+# ˆp�[{�+ ��,X�0�kG��s���p�XQ�j����p2�0�_ͅ+�a���|'%yR���"U�G�W�X�u='f�Z�0ӫ&��kz+��"(� ���J�\�0�\r����;#�Q1�wVG���'��N ��4��ژ���l2t���	J��Z�%i�u1��%HD�s"g%�P`���&&I���r���<��;�&����3q$P(I8չ��3�ӫ�ח��A�����s����>Wt�uD�W}t�C�t�D�ʄG�*�>�EM�PS����	�p�7%���g��|\��[}���[��뵑@�\ݞ��^v{��y�} �E NGq�ԋ��Zi��ev�s�ĺ���n��6]���w��w��}���G��Bj:�PUq����!/�C��]��Wt��K����~����>~?�ǿ��FےI$�I   �@  �_�� m����@   2  ��pւ n�    �� ��     $�;tq&�$�bN�;��.xm؉X�C��3L�4?Cg�7�yV\��t�6]���s�K��=eܫ4`;.���	U�I�qG7kL�u�h��L�a\mu��qf�UG$�\��N��i�7jjt�M��Nv��,����Uge��vuu�[o`
�{-m� ���T�'D�@-P �;�q��v�މѶ/Ak��̓�r+�xY�+���;b"6��68}��*Z�G�殃-�K�O��]g��+
[��(�[���������Z���k�����gy
�.�8�e�������rlu��dNt�<��v�:S��۷l:��1ZvXϭR�4F��p�*�+�h6'Z�ү<������\^OC�T��}����V�^aة��}��{U�a���t{��w���q�~U��|��>~mXۨ@�g2�u�<�x���+wC��PΣv�*s'^;�q��i�@8�F��|:wU`�<njM�me5֪۩UT)���Ԙc��s��d]mU���!q[/& �1����ɧ����;ej�ҳT8�m�z6�S�L[����n�6��d���x�	����э@�݀�`SIPVp!\�܃1�CE��xy�=J�s*�����Z��pt�n?#���fm�u	���UmYFuӶ�Ĺ]�^�� &��m���ܑ����UW1���G��ze�:��۠�5g�Wh�;W��;�˗����q�\릪�k��B�P5$k��d%��26]�v �4�6f9�a�vcE�D���U[�!+λ8�w*ЛF�Y��ʪ��F� 6�FV��W�� ����!���U�?|��2�O���Q���Ng�9�Vͮ1#u�F�ۨ�3=�v�����<�6s�A����\�̦R�r����6�ѻ=�m��n��/0�nj�\<�vs����{5�1c���&E]�g��f9�q'Ol�K%ǔ����n��Yv��G,�#s�f+�켨L�n�c �l���2�KY��ŧhjڪe�� ��g�v��jxK��j�;���=��qס�5Zһq�nMPYj�T �{4�y5kv�jU�ۍO]T�K�,��T�R��:�wV:n����õbN�ڪ�ZB@.��UƛT��v�6a�ɻ�+�ƶ,�o)s��MT����v�1l��L����T��W��$�ڪ�om�@|tў94F{/@\��X��9���f��s�V�#dآ�|Ak��2��c�]�cfy���4���+v��'�]�����M���(�q���ӍQ��jx6���1�W�ت�.��ENk'k��۷]At�:H\��Vӳ$.5�A�`�a��A�;t�� ��hy6��zN�7��z�a^y��`���lЫTN��g�1ѵY5(�Xm����m��p. ��/[KoL��k:�M	�^��m�e�m�I�  m[m����z�e�ssIR�F�R�*���6��mTG��\�u�N���V�{V�&�S�(�<p�UWT��� <`�=ĳ�gGU�ڤA�"fv�m�U)�Pt�U�\���yUE�N8ej��.���̨�jp�=�����||�����0�x�
v�uӪ�k��g���yC:�6e��٬pP���J���Ae������Unk`�õ�p��5U�Z&����֪�����]e����V��r�D���vQ	�lq{	x�B�2�p^�Y'Ki a�������j��R�j^@�j�R�5D�ml8	6݂@$�[f��*�U*�Ye�Z�K'5\n�ze�yYT8��UUP�b� �d��v�M' � m�m��M,)���Z��UY���H[I�f�`ڗ�h  
ڴP�M��"�@�5� 6Z��jکUV��0V�f�8 ̌m'哾�� m�m �f�Am [B�m۫I� U,:�݅WF�Wg��J�//]R�B���9�'���5N�H)�'Ju�$�ge�:�@y�m�  �p ]�` m���8��ZE��}��O�/m��T�ۛl�i6   ��		��4��3f��� A��m��l:�'@ ۭ5T� p	l�Y[,�-��v� ��U��Ke��]�;������^��A6շe�[���UF�jUUڀ+q-���nݰ	�[%�6��m [v咤6� [Rʑ� 4���ӷ2�: [@$[@i�*�k@���m������cZ��&�K��v��k� pm�d�p mZۆ�f� H �&�f�-���-��[x8  6�m��q�@{m�Z��m� m   �� ��l  sm��5�/-�Z�[BC����l�LigJ���f^��`
�m+̵*ҭ�IaJ�������W����U�Z)^�\�5U+ӻ$��@ � �mmI ��%��9��`���'� ���  G �  ��L�m��,��b�8 -��m��ՠ���e�E �m�����I�'IȐm�8�����U��N��YP@ ���-$*�];u��>�u�q�+7��(�<�A� �P�n������[����f� ��l E��`�U����]nG�ڻq�q�[f�� -��kn�i7�v�  l�T�m�	�\[@��I�vں�.ٶ�-���-���nٺt��L��� ���ֶݶ��^Iu�v��am�,�e]��c��hP6:�j�݀��\���`�f�W�7<<���v �W[Yp㎃�]0&��)%Y-�-�zM���v��E@@mF�Ts�Z�T���ל�5��%!�  ������q�����5��v�K��� ����   � �lm� ���d��ll��nk�l��-�G �I��кU7�O��	V�Zlk[jͰ����mm����$  @h     ��  u�   kX�m�  �� l    6�z��n�L�Ž@5�Uf�h�s�m�  �m�� �6Ͱ {e��`4P���Zl-�ll6� �WkX/U�p��imlm�@�   �m�  -�4V� 7m�   .[      �[p   [@[@S[�m[v�      	 m��` m�  p�pm�	a��`�m�   M�� ��   8`�
U���Y�&@e�   -�mY�`z�6� @���`[x6�m�A��n��  ��6���  �\ mHA��m�����Ht�  ��l  �  [F�� �n��$sm� �H     l.� l8$�m��`  @�l.�h5��  ��� �oW��【m��k͍� �� �`��V�h    m�j�cm��f M�  %�L�ll �H�d����-�����`�{ �3v���     l� [G.�m�8�W�@H�[_6�| -���l���i0SI�6�d��Q��g �#�Ӥ -�5�Cl��]�q۶���Ͷ:Hƨ�
Zڥge!���ﾪݪ�Y�:��������R�j��8W��,�( rK�\ �/Z��[�  [Kh-ַv�$�&�  �-�Nݴ�8p -�  � �%�I���^�s�i�I�#MH��� � *�z�le��@���T$��ػ+.#���Ƀ�u-�eڥJ�)US�h	��T����m���]/�� ��_V��:�ȸ p�5��d��p�v��.�pEmv[Kh ��Iz� �$[\�s���UUYZ��������t��:蝚��j��	�Pܦ簦�����]���`�r��]R�tpTdU��t�
�H֭��Hj��>�$}J � H��&�kn [u�"�M���Ԓ�d8R��ksa�4�;6&�Nۺ.� [m� -��ռp�I�6(�L�ڶ������Nl�n  G�ԍ�J�t���P�$J�/_,q�t����bЇD��#H,VSF��Q��)�5�.����k5� �_Z8�һf�  ^��� m�����*YnJ[@	 $ �H��b���m�V� z���m�G[�ܑz]Tս��`T��8%UYUV�����j����Ca����m� ,s����B�,�d� [@�`�e��l��m��  m��@� hm��PlJ��enT�m��*       -� e�D� *�l�mm��5��$m� ښ4�[x� 6�i0�����|I���v�Li��J�bI m��� ��L 	�H��$N���lH0�s[p m��z�o���{������0TU?o}�(/�?03*�#�����G��: ;`�&VfF@��&Vf�fa	d&Ba�fBfefd&a����X`fff`��� ��'������~J��*bi<T6hE!�8b�� ��0����"N��/Y��*�.���AE�q}@4(�D���.����CB'�CGC�^�0�9
�@zA;�c�P;Ux!��6&�YJ��!)��b8�2H���M�:�	 e ��v�
��II8 L���CgJR�B� �@��` �Á�:8����w��`xB����D�D� ���#�� @��^�����{�z�OE����P|d�N�]���"�w������B�8>���`��T|@P�"2�D��D��@�����>�L
v����&"B�B�`�Ҫ�[<8�!����W�4"� <BTSjhA<y�+��T;���a��p�(�
�j�4�v�v)��;H����lQ�@� h6 '�@���S�z7A	�'�z��&'4D�!#B�J�H5,���8�@��� Ĉ8���}=OD���G�]R���$��怜	��>����P{T'I������N
�{�`�@eE�d���J3���$&c�a8UVdI&A�3���> ���ZBI)�H�� �&&^�v;�G X�BJ����^�& pʅ���A���;�P�t����� �Cb`�B�x���ff����US�L�dS"�����@ ��m��]��-����h-����h-����h ���TP@UW35�k35�k35��/��������z�� �{�����{��{��?�~;iNܻ3�Ba�5)��І����j\���h\)lt�I�&������IRB�!BD����e%I��kp���FUM�ou�u�����[�V�H�S�
�X��s~~*�G��uU�*�u��ڪUUU�U%[n��nwTn�?gݾ�U����G�b5��b�#k9+O5sS�i봄��)v,1�����j�tsƱ��gv�i���q��e,�rv��<�On���c�S���=�|��n@�&۷ad�6Wh��C�7Y�c@'#v�g78�MXz&��M�����#)hkZ��.�s9;8�g�^�l�ڬ��u�4c&ة5.v
��;W]�Rc���u�f����s���3¿mb���Yu](<����::�6�4�ۥKy��%��^��k�lDۊ��$��&�3i,t����MINI끖�-�p�n��Ϝv�o�v�;w��7n��b�۰��wt�r��z���!7l�Yv���[I�Ɩ����F��]���]U��<�\Lbn;k��F:ЧH��<;g��%�r]3���\r�b�$�*lc�;��ݍ�CZ�$���^3T SY	�G��ml$���u��9RS��qؙ�Om�W'��s�8#��^;e�6Վ{u�$֍u+�*��gN.)1�,����5���vU��3;J��&�x�E���rp��&p�&�BtҋM3k�v�X-@����9���z��&q��Ge��wk���=ў��t>���22�g��F����`��.���E�ۯ]56�-�$�Ͱ�v�%�v�W�ܹ��n:umجh4+ej�-@@E��kb��
��j��t�r+�S�÷L[l���xUU�um����^�T�	��Ⱥ�`��vzY�-Up�p�plj�)�v�5T�u)��%�(���0[sC���r����}�����%&ظ�vPU�\�۴Q�9��ų�=g[t��l�����p�6S��9�pK��N��GZ�t��:5e�:w[[l��ָ���-6��k�.	�vvm��>�%�d�7�E��jd�	�O6���/���t�ak6���� C%�ԺI�IpS,m��6ay���#6����{�`(v�z��B�*��4)أ�!������7؀i@<{߼�����;2�F����u�z-s�q��1ݡ{H�b���̲��w[�d:��I�~�qmn����c�M��}�|�pL�	%t��ix�fȷN.��ez����x��Ѹ�864�j�GX����з��j�1͔d":��fv�[@K+K��{ŷUM�ż ��o�-��s��E��Ĕ����NI�u�6�^-���wy�w��>��<�;!�y�W��Le����m�q�vy�W�鶐�Tr�����W9���}��U�<�s�+#R	��N
9��w.��xp��Wz/b���`�q$G)��u��h�{���wo^n��z5��L�1#̒�3"�-j�<����W���w�l�2���P�������^nҽ}�m�l���w��U���۱r9-�a������B'X��훋��G��enLs:,D���w���m�wR�}�m�l���ΠYm���Q�zѽj7��o�~�����J�2@6��Đ�33jIM���[�����ڮ��U��5�F��k���W{K�U�W����v�n��+��qE$��;���;i����ot27WOנ��0�#�LK�K�y��}���ن��J�|�$������]Mln���֝�v���<7+��c6I6���Q��0��d�lr,��w����Cfj����;^��,���`O13)�Iwx�l�����;^��+=�̐�{��1/)�b̸D�/k�;^��k�2L�)4a���{�~�D��K�92�;üK�n�iY��l�����;e���� bfiY���{v��?��77n�:��m�$pj(GI"���p؀u�+�K�E�RQ5<�웆�\w{�wV}s�P�2�0ٛ�W��v��ҕ�݆�^�dQ�#�ƒi;��?bگ�����m�L�t�z}}�M�#R	�#n(�_s=�J�n���{�Vy���ٜ��D10�/��4���6f�U��
\�ȹd�̾�U}��v]��Kpj���(��'��zW2�G��;{�Y��ne���t�(L5�ۍp�������+'/hpkX6-;��JyL�]F5r��[�)˥B����~�g��n�/l��3$'��`�ճ	�a��2�;üK��nҳ۰י��<��l�F�@���!@���g�a�3g��k���R��u�xy�3.�"arď�i+=�b��ٗ\=���v��#�G#�$6�g���ɓ_ou�7�36`d�&dh%HCB�A��¢:�VSE��6*&4����ۤP �G{�z�:��7��[�ԛOn���mB2��[h0�i����f���l�u�n��ջN����㛇j8�l��:���y8gJ�Եɺ7Fn�m����<�&6�h��;oh�N5��a�b-.�kFԹ6;�ٶwn�mIs5<����F�j&j�n����_|�5�7�.I�u���V5�c �i����{�6Qa���4��ϥ��u�|���w�~_��<u���{\mrn��O����*��am����h��r�{E�F�QH���m�f?���uw��VeybH�ƔN2	Iu�,���������_^�e���$��J��r�$"���J�<�V��a��.���e1)�a���L�z�;8��M����nf�׻�1����I4�_s3�.��Y��w��ު�&e�f�DG<JD�%�e!��ڵ�� �F��y�[&�[���Sw��T��dBs������W��-������n�Vg؄�jP��2�qW��~o�:(d�_(M�_�LL�̩7z1�����f��]�]�fffbfb&܈�[�.վݥz��י�Հ�^�8'���Wꪯ�9��u�[���{�#;��_w��(�(�b��A).����$ݻ�K<��qWn�+�̢"5!��^4֡ܪ�;,�s�
�kv{=��˛]4�K\�i���Ů!&/�/�����yڷwi_�u���[(��O2C�R�^ťswv븷W��rW=�(�Q�$A/)܇�v���W���I��d��ꪻ*���y!�y�/��w�#E!G�ҿl>�^f��|�I����m��mJ�l��_s��^�����ٗ\31����x2�DiJ:�Rt�)1'��CڶCRL�In��帷O'c�Wi�[�܈�^��]�}�J�݊dl�-��^�q�8�m�ԋ��̽;�u}�n���,+�ݭR�i��#��R]wV������y/b���˪�RY��)#r�IH��fʫȏ;V�v�yv �����d0�A�84�4THR(��UP��w�t��`�����v{�VJj9I��QF�����_mW=�����_w��]{��D�A
�:�B�:�����t�]qs���v��6v����tн{�Ȥ�PN
St�q}y�ˮyf/���uw��v�xț)����#�\��[�}���{ew��/�}�~+3�`�R�8�!2�y�+1��վݥz�����'�329�I6����_^{2똳��r}}Iw�I�DܑH���e�1f/����w�{A�'��R�x��tsE�ތJ�ͳ`��t�f]Ӊ��c�k{q�6ׯ]�<�7Yr/g�Y�^���̛��<��;SHd�,�pv�:�v͜c6r�4.3V��<��V�N{a��;rv,v�۶ڎ����lr2�m���������@�Y�|�4� �vA��p>.ZRCp�c����k��\1���\�	�WF@�.�����dL�e��&mʶ�*K�{��{�x�ض�M���N@6߻�m}�5մ#���pr��-��� �tKH�AE$RF"8�%'�:���rC�]����ˮ�I{�9�! 9��rU�睫}�J�����j�P���
^a��,��]�}�J���׾�����#�&Q
�]�}�J���כ�W��v��=�1rb]�bi_�u��͞�k�_{e�xEc�A#	Q�7�_*��Jy���٧u��9�ix��̎�1��^��q�v�36��K���U�睯}�ɓ2V����{R��9#q��w^��/}�y�}�%_|���JZ�%�B۽��7b�y�-X��^O18)���)��f]s�1}��s��_s�^�RF��DqJK��<����!ή�}ܮ�]t����Ir���+��J�|���ҵ��v�d֙���w�PVg��%-���4��Mʔ'��Z�������q�]\��Jh�?������k�ݥ~�҅��+=��""a�x��D(w�v�����3&c;����ef>y�&�^7T��ډ0��un���������zl@  ����  *���  ���gI�<�Z3�ֵߓH[�t��JKz�o�t��:��)V���)�EǢ]QD3ZE�,�F�1j�q��:�����V���H��o&�,-Grt�a``m���̃Z,��0��E�o2�dA�a9nw<md�ð�8ff�Y\y��bd�ˊz;��gn��0ȯX��n�Yv���.�D�6��ޅ��28��$�\��y��ȉ)��s��������1�-M�֑5ӝ�������	u�'[7sRr�+6�F���U=s|f��4i4�y����P���e����.��,!��H�5���8�):�*:w�޴�7kq�E��7��c������e�E2��#Z�LM�%���3HRgk���4;`4���I>��
�GI�]�d���!g�t���6 vv�M�i�<�z/*���hC�= |����XD���1R  ��r:8B����C`/D#�A�C���@��5��z���)��k���R�������ԥ)������fZ��7�E�o8�I���<��<�^{�R������ԥ�(������┥����~ٚ��5�����`�)J{��8�(����X́�	����2^��8�R��D��^k_��n֭�-f�a۶����8k�T�hJ��sL�Z�K�ꍬ)^����qH���}A�W=��믹Hw�>��g��)|�<���R���j��������ߨ�4�b#�����┧�o\R�����JR�y�=�)JP���}��O�A�%1j��*RFܨ�q_�P}�}�1��%)O}מ��):���=JR���W��}A�{���jSu�վ`�)J}���8�)I�{��JS����(I�&�� ?DziBD��iϴ�y�0�~���}�~�����MA8�'M9/�>��������R���\Ͽ6�ߙ����ߛ��ߟ��?���&��#[[��i3rx�.5�X�\�s�ڷ#m�DM*�̻q��\�k���JR�}�~�)JR��{�%)O}��qJR�����R��޾��-���{��U���R�=�����JS�|��R��뿾��ԥ'%����s��%����6�M�d�ȓ�7r*���!�O�>���){��~��)J{�{���)I��k�`�R���9��Y�7/C��ʚf@�+���$�̵�{\R��rN�����JG�|��R������O�i�Dr��}AU�/��\R���<Ͽ0{��=�s�Ҕ=w����)OЇ~�ҚT����$�F["f�V�?�;g�x���;sO^���|]�h�q<����E���i�u���wh�[#t\{6�®�Ir�z�۵m�bv&���r�׮[v��=@n�K�{<.!��{��܍j�۰!][	��v
��%���=���;:sm-6�R""�P���:C��������I�r�@uʇd`UT��kVj&U/a+7k\f9��m �%(����}�}���}W"�$7̑εP�ϫ����s�ɋ�]�t9Üt�ƥ&3�y�Q?e���`�V���޸�)C��y���)���8�,����Ԛ�d�_����3 e��#�����	t�v��}A�՚�U�}D�']����(L�ߵ�)JEﵚ��*���=��m�N'(u8��);�Ͼ��)J{�{���?���X�>g��<���=}�~�)JRy�}���K��q�i5��M��fT']����R���y�qJD���7�5���ۭ��R�!�^b"&)�R��w�{��J�����qJRӦ���Rl�3-~�f@́���(뵷'=��Nvzܶmkv�e�nn��Q�&��N�4u0����u�5Gk	����u)I�����8)I��{��JS��ߵ��@Y%);�?>��){�-�LR'��E}A��W{6�������'��+�J�)���渥)C���<��=�^{�S�(K��������$i��:i˯�}�Wߗ����)I�y��<��=�^{�R����6��}A���0�{u���I�┉K�~k�z��>Ͻ�\R����ޤ�3 fn~ފf@́���t<Ģ ���K���:k�3-�}�d$���~��)J}�{���)I�v}�%)O��{h�ٽ�y���7F����lQ�"=�[g�����nݵ1�^��7[-��C�N�/��́�/}��&���g���)JP��}�!�JS���u�)J{���ݎ[7�z�e�o|�)O�׿g�):�>�������R����qz��#�_K_,���n "^��3 ex�����gH�ckc�S�]"�nz$z?	���'�s�{���)J{���)JE}��h��F% �V�H��}A�իs�qJ�N��߸=�R�}�~�)J�s�qW�}�W���eH��N�#&��)JRw�׿pz��?I	����3�Ҕ�ߙ�� iOs�=��)9ꯪ��g�Tn��t@�"���aH��fϝ=������R&	�re�@�����w�_}��yrb\��4��d�;��I��+�>������뀍)C��{��k�}�*V���r��"���������py�!�����)JRy��ߜ{�)L����)JN����a�l��^]�a��i�X́&���d�g{߸=H~ d����.-)Iߙ�U}g�P}�{3�CV���u4�W��@���y���)N�����(z�>����<�b�wu��"z(�}�y�����Ϸ�rٽ�FYf���R�����2rR����JP>y�=�)JY���{��J~��������o�9�'Q�'M:e$�� �jU�J�ܪPZ���흸cI~{�ܞ�b�-���ֈ�[��)Iߙ��%)O<מ��);��߸u)@������d	���:I��%D����t�3"S�u���? C%)<���˃�)����.)JZ�����+P�vA,��SRJq�E"��������ۯ�)Jw���Y�s1�U��<��ϰhf@̷To=3 f@����13/2��Ĺ1I�I�$�gGs�2d����)�oۊP��*����&��3-tr��"d�Q��%3�']����R��=��}pR���~���)Jw��p�4�'�~�_%1�!�����~kxj�m��P�1�b��v��%��j�qm�9Ͻd��vi�7\;h��kb*r����$�zv�Ҫ��b�v��h�n�q�sv�3��N�q��^H��ڃ.۶M���Wn�r�+`Ř�M;��b��]��b��9�)�帒�����ؠU����tRN�j������&#��s���nzcq����>w}��L�vaL6N�֍oZ�h��Q~OM1u\ֲ��3�O�v������VN^����ˬ�=,r�u�߿{���|�n�B����?�����w�qJR�����R��~}�
�)Cߙ�<��;�̏ukDQ�!B�QRL�vou&��d���~p�'��`�R����Lə��-�-���TÒ�@���=JR����8�)B���{����y�p?��%)?<���ԥ)z��[_�TԊGEE%_�P}���W�f��)���┥'�~���JT�.�T́�l�;DGA*�Q.�53�ԥ)�ޛ�┥/������2S�~�)@�w�y�%)OOOp���v���x�ƍ��Um�ч���N�����7�͸ۈx�w�ﾻ}�uBTΒz�)JR}߿}��R���~��({�#��y�pNJR�{����>�d���>$qȢJ@�'.��U�}�g�n����ڇ�=(}��z�Ϥ��RM�2��FRfE�8�+�1�ޛ��@�a��A3 `�Y�#4,��A���R���;��)��J�`f@����Mbfe��r�S����kf�޶qJR��3�py)@������HA3���~~~p{��1O����>����a����D��Cԥ(w���8�)I�}��JS�=���JO<�=��)�>���x��!<�ʦd�g{���3"���~���~g��<��9�˫��
����w�g��$ģ��9N;s�l.H�s犡sF���nثg�5c�ۊ�1}�O��:��U�F��{��)J{�{��)��);�>����~���4����pz��.�k�GŚ�������qJR����py�$��=���8�)I�翟��)O|��A�(z����J�"TK��L�k�3,��T�c�2$ϼ��R���v� ߬4�N��`&k���~~���!�/�Ѱ��$�̳<��&!�b&�7��������pz��=�߸qJR����py)H)׾oۊP4�=��r&�Q
@��.����}Y�ۮ)JR���}�%)N��~�R�Y���3 fZ�Tt���8�bf���rdk��,YZqa]�l�$fmЛ�WY�
�5qUz8p������٭lݛ��)JR�}����R���7��(N��︠�R���{�G�);�̾����LI$I.EM:k@��e���$�HfE2���?8=JR�{��)@ĝ��{��QS�<}գ9oy�ַa���qJR�����R���{�)O��� d�y��`�R���~�)JRy���_c��7��Yf���R�Q��~��iJ�Ͻ��)׾{ÊW���pqH�LMF� J���(�R*a�� ڣ~ ?�_��}�R��v�E���,�f��oDo7��R����{��X��	T<��uO��JOu��~pz��=�߸qJR�����_ZѬִ��n\xj�+����=\��]�$u�El����n,�Q�}��{�||c�]�3�G{�{�Jw��p┥'y���)O|��B�����JR�y�f�M�z�oz��o{�kw�(9w��}���>��qJR����py)Ju����}���f�{�(��������S�=���);�>���R�{����)I��}��JR�>>>��F���٭lݛ��)K�u������������)JRw���pz���Lݽ_́�/x߃�&%I2o5��0z��;���k�d���y���&�0{z~(y�Ao�Ջ�O��TU9�q�UT\�9ǕUW��W�B� $�$�H"	$	B	Z@�$���� 4~�l�]:�å%�I$�J}:�����{'[6w�� i�l7�=d%���s7���"���Ͱ�$�G*�:L����֭���Of�|��� ��4�2�JM,�x+N�![�FcJ8�&���7��H.����9��O�4lJѤfZ��5�:��̈b�P٘�{�A{QGW4`V�ƪ*��ø2�y�T��3[����>�mh�@���:��b	�J��R�9H�=��>k��G܆S���ˑq�=d��U�6���[��m��!�Nu���qK�u��;i r�R����\�����ust��k;���fUL;P�o��6ٷ�d�p��;75����v�ݨ�q'aŸ,xCr�m��D�S��<h�2�>��.��S�tّ�n��Ltp�;�!�38d��õ�Ǯ�k��ṡۀ���u�mH�������J���Kg�z�[�J�g���q��K�k��t������[J�̄нsآ�7[.�N;Y�ۇ���0>�A�v]�3�[�$�'N������W��ܕ�6M�C�:��F��-�d沭�`��5k���`guS���ՠGf�(�nj����]�/6�1�F���[f�;j��]9�����v��8��_��9�%n��٦j��N;sl��9����v�J��v�s�p�N�9ΕݺۂD���̪�;p�[^�K���V�)��5��K&"Ü�c��jR�7�|l�5T��`4�m�>�[*�ۧ��`�(J7n��R�ܤn7;�N��	<��B�h�C ��r�z�^�\=��g[x�#�m\�F����\�1�N
nV�ǂ��z��c.�6ѪRL��͏�Cg�z3�.[#+)�Ŏ6U�m����m�U��-i!�Ӓ]�E��)V�#��J��s�e�&�j'�%2�ʰ��c�Bj��(4Af���v��&�J�»MZ��8N��K<UTms� �ĸ�[���ڸ�lu�#����.���Sy雛�1#��ݹ5�����f�	�ȗ<���Ψ�<q��S���5�X(�XvD��Gu��@^���J.�2%���l�+��N���;f�g\tZ,���XTi��S��N��L��|����Ӥ�ћ$d�1�y�����]Z��&��]��)c'3���;����.���v�ɦ���w�	��Ў*�~/���(�(�� �[Q4��C�?�F:I �{B?�@?����kk�{��)����5J�J�*mϢuv��/��g[��c���v9�	Þ�^m�;v��';����ɧI:ɽ��-$�N� zu��� �(vڮ%yͪ��t�sQ;]̆�X�*�yup[q���R��:�BoA9��Ŧ&ݝ��n��r#=(��  Ҁ�Ʀa2"��
��uN��źU��e����ݛ�I==-�� �J��7��P:�VC�;����w�������'k/!nd6��ɀ�9v���ٻ��{s�[�$���Y�)ϻ����u�@pT�p�9�����9�;�X��_UU���atxզ���:R�)D�� �t�L�y�@,�N�������3^����КR7�t:���<��������~{��]U翟�9TΆh-dcr���J8�������=�޻=�J��Ax��@_�B��q�H�d�ȋ���p����v���^�;�L,W|k�$T�� �oV3�����V�� ƶ�rq�tc[��n�bu~{�>�vӑ6' ��/�}�u`s�qX��>L����﷾�]r��3
fd��kf�޶r�����?g���0��YJZa%�����e��@&�d�� t꧷����>����u*��fL���_/�^Q0�^eK������=/;z�I�}�u`r��U�����J��ੴ��31k;z��u*�7��L��#ج�M_(�GJ4P�����Հ$ɕ��=����޻����q����fL�����g`�g�N���kU8�e��w]nrݎg������n�;���ۥ�U��s���zfv��ə!�d�tg��V����"!ۋ�{Ѽ��f@fv��=�J���篓'���Fx��$�#q�E"�=�����>��.���v����<
�ֿ?3�f?j�3�W�oZn&��1�9��}T�$�����)�=|��e��5�����`yVVVȪI�B))Z,� Mw��ޫg��P�9�<Iuvz�lZ���c`��;F��-;���"kV����s��G>���r�}��ē=�@fv��=�J�&�;����5q�H�M���n�8W��f�XL�v;���������#�(JNpf�Ձ՛�Ϻ�[�+���v &��6C˼�ḐSJ�dɌ}��=�@g���G��ɼ��gK��(i��	Ӣ<��ҡ�472��X~W��@�=��L�30�S�ŀ�Ѽ�ɓ3:oi��V���T|�u�3JۥnRT
'%N�k$�����z�9bZЃV����Ź5���&>�?l�%nI)H�dqH�D�{��n�X[�������OZr&���35V �өW���N���({g�ޯۼ��nfժ���D22T"r�8���Jd{��vyoR�3[���
)*#�-� ���]�n�8}�uaTun�;�X�c���8CDDI@n���o}���1��m@k��(�ӥ��'a ��̙~���#蘀7I��cP[���Q�5�mgI�ҭ�)�q���d:n��6����'�sm�8Q�����أm��w,�6���]�r[Ӷ���]�mgٞa�*�����W��zD�i~^�6���V�
�u��ح�η1�E`H�^�`,�S`+e���6�bN8:�t�t�m-V�{c��[��V�mqѺd.q����^	�C����kz��Ѳݎ��nyeL�!��ˍc��[�B�m(S�X���6�8����#�(JK���˫8�'/#Ɵ�fgA���]������E8�ۢ�r���~�謹�sK�;��]��ʚ�37�9L�Ò�O3oJ(ԕ�������wt�(xh�2H�8��r8\J�x��pfmՀ}]3q�w�,���z�R(ǉH���3ySPffݟz"���E����p�+��݊�mD���R�&��۰g4nu��ӓ���fَ�]x��.�9�������)�9VV�;������w��;�۫�6�G�BE%Dr�몎��\��#+�}��I���	}���r��^����ݱ_�$̝��f�W*�(pT�p��߿_ �iQNϏݱ@g�t�-�b�x�h��xD�C�f�Y��T���ؤ�J�$&O���]��Q�'qDđ���t�(͞(ԕ��������v�h{Ov��]˽��M�
�L�TV��b8�7Ow��P�}���ݛ��mL�<�X�w�=��{�ԩ��2;q�u����:N'!�@{ۻ�~Nə9�߾�`k���@fvӔ� /7�����#��6�8}�u`un���?�u'``��D*ш|�'�$����3��'‼��=�5��^�p)�R��a�|un�;�L,y%v�}�3�{��������I�����j,ޔP��*�3R��c.�6�������,�G'��l������
�[k��p�B.+v�6�tu�����0��7f�,D��J��}���t�>f�w36x�;���>M����jNp�v���n�Q�����M�J��|��3���U�H�$����`/?ߵ���?&I>��]���R�0F�w�"I��	x���2��������u*�i:>S��C�
������뾭r���fyF�'��I*��n��w۷V?v���@~I�r�~���eȗ~.�l�!�����qv��^��v�b)Ɇ���b��|��7iIdr�ܾ������:wlPc�^�����jw���bACʕ�J�1��(fH�l�#���p�f������^Ix�[��r�	�w��� �^�u%mc}�f�E��<���h`�(J��m�t��J��(�w�K��37��nO�~v�R��T5'8}�u`~���U^?~���oM��}�v�ԙ&�ђ>����%vݽ�ݠyc\�6�^�"�켏lm= :9�n���<�ۃ��+�K)��[d��k=����d5��Vt����˛�sd��s����Ѳ����7b�(.���4n!�M"�* �n59�݁�){mU�Z4��+'H,Iݗh�e�H�f�F��D��0y�̚���4q݌�WfIzlo-ۛ�ˬ�z	8��{��w{����=��*4��t�r�C���E�0�F����r��*��<gn��%~���W`�)�)�E%%XQ���
�3=�hf�u����@05e-D�R�#�uR�͗_�n�8�nʰ:�q���}UI��6H�8�e�ff��������SP|ź]�X���JH�jF���q�ooU���N�#3�43&d$��~�������
$%"7*�8n�d�g�h{����wR�>�$�\����wZ��׭�v)��^Wqx��a ��X�)�"�:����.j�uMX?����m�{�=�޻=�J��2�;���t� R�J�
]��f�����bK���`g�A�g62l40a2�X�%	k!T�@%��G�=AC-�p�_���qPg�i���ktt�
&`�xtC�ڰ3�Ԩ��z>fd�I�d9�ޖ�߷�8�իlE9%&�RRU�y�B3�4go]�̙��t�@_CR�e���"j�\(I{ٲ�>���1r�5�aJ(�I�fޘ�"]��^q�����s��|秤���\"j��iДq�]զ��{�S�:|7\c;��^��T�������k �H�=_�S_��(�q2���l���_s�g�h�֬L��x��3������Gz=�`y{��)�S'�����8�����8������̐ٮ���4E�|�����B5�gi�C�<��5�����¬.:C!-F:�]��i�R���@�
i��>�Î>�'�Ό�Cp��ތ֛4c��k�^bF]t��5��" �y�b8�D�p�K\͇dd�09���Aj-���9̫���]b�8oF�@���Nø�R�	����Q2�z��&��3	=�OW�$�jKy�N��Ę^#�=M�.*b�В�v,��g��a.
��HS�4�Ba1h;�ґ�W�{����]�����gh� 8"<�i�C�BТ�"�+�D�<� �|xzEOq�4(�:U�^������=�>@���/uϳ��x}�Ձ�֬[NIB�#�	>]��^ͧ@f.V�jT��$�v�?@=K�*S���qX{���3�4���{����c� ��[[{M���d�6��*d���3�|�T<�d�:m���y�q���C��ϛu"�*4��ٳ�i*9׺�|ӣ�|����^���􃻍2�t�'�{��F.������ͺ�U �XƯaul�+��8�}��@f.Wg����=���l{�@g�JX�r��H���U���p�m�*�}�r�O�thIHE�n�<����=���I�8�ܜ�A�ޥ@
������lP��v���N�{�]�}�{�kpd3�T��9F��I\XW�l�20��
�4b5v�z��%���k6=����z)���+k}�]X�tq�$RA'˵�5��S��]���5y	=����
℩N
�JG`v����U�۫
��{����c����[>mԊH�av3&go��R<�Z��3��vpʁ��2�!:w�T�$����f��Q��)�����ySP��	s!/�^�f����w�e�����t2/m������xy�l���8�65�M�!Λ�vu����[���X$���m�d筹T/��v�H��/s�؁�b��n��/�8�}���ڶ��(b�c�E׍��D����������*���Mq��+���Ge��h�ol���Gm��0x\vw�m =��c���U�<x�Z7g̈́�u������=';��Y���Y��h�j�<z���sv�X站y��!6�2nҜ]//Yrt���!j�R��qG%�\���~�?j�p�mҴ��Vs��X6�'�Ԅ�����bHw�oZ�/#����/��x�c{$qH�nK��*j�r�z?o��5!M0�^�kY�H�G r��&�X��V��&���vd��oR�/9���bQ0�^fGx��V�ޚ	&fY��Vn�u`s�{��f=�F�%62�1�l��ɞ��q]�z�8�#�.m�o��+�JM�)%JpT��,�3y�;�۪�Gs�fM@�٠E�����0���tHD݁�ަ�_ƦfJ�$��C0L98�����+�����y����1��]�6�wb�'N�*����Ty�L��޻�^��X�卫ڗe����ݮ'd��z$3����l��2�7_��2A*�Ԥ�*�$���w7��͵@j�OK��hfK�/!lt�366^1�:1���k�k��\���*z]��r[�X�Jߞ�h����Z�_~m�ySP1y	=K�^oM|�n�W`����Jr��%g)|�Հs��`fv����T���"TJ&����T��ޚ3����e2f�z���$�|�)P��y$����Q.������SL�	R� r��f�w՝J����&E�hzw?LD)&f]�7`g��Pfex��An��`w����[I\�)!��`�k��K%��Y쳋v;G;��\�4��κ���m�H�t�'-.u� �&q��w�$�fL�����Fx�~��UUO���E=�g���L�fv�؃=�Łν�V{�BX�r��H�T�Kf.޻=��d�W���y�@s՚��R8��������:�/#����4���b@�	&fd	2����k�yA��beLD����#�J�/#������l���|��۫�0�����4�Q'Oׄ �k�F��-;�ݜ�:�r/W��L7o�w���ڎu�	;�\ �ah;�����P�&ff��}�Ѓ���;�Լ��D��"&hϷ��Ja�2���R�G�>����;|�f%�>�����$̒�7`o/PSy	= ^oM�����XŰE8���IIV���|����3yM��Ovfg�������{��T��#IG%�\ �e����}�}���R�3��� ��L�%7�a�G��s��	V %;�+��>���r:J�ܟ6܎��2�6]��zM�ݓ<h9ӛu��l;��"�6��F�N�\A��68��<p.t���O0<��l忺_|��J6��p�;���N�yF�.�vԼ�l��:����u$f�_���؝���kvN]�b�z�b�d��9�l�Y�(k�K/*����p�6���qv.�霺�3�n�*�"u�r4��W���{�����w���w���9N�^y� g����z펮��:�4�]q�K��� ]$���V�nhfF����{|����M@�란/=���P�I$R8�s��ͺ��$'l}�@��F}��n��["��9R�ܫ�{�É.�%�#����;�۫�՚ە 7Q� �e>���3�����*�2I{'�V�R�
�� nK��U�����\�{�Mk�t�0>R��":ۅ�6t�=�܅�#��t�'YwR��. u��� �t��G���[[ nl'z �ޟ33[8o��v��A��n�%%X��W�}����ȴ������o��}矟�uW}�u���N��KQ�(�k�����4-�v~(�S�j`7���ݑ�nS�9
�$������ �{6����(�s%��j���'qB
D݁�ʚ�<�}��y=�f�4g�+�A�u�-r:j�����T�479�y��ӓ���m�y�tl�]x��.������5l�*%K�D���נ�[4����/f�X��Z��G)�A'˵�mJi���[X����\�0n�?@+�E�r]��Ӝ�ͺ����� %�	|2��=Q~W{r��[ 3d��,�-��jO��� y����r���O@��@���޾�F��AN8&�RRU��=�`$^{f����3�Ԩd��b6C�N�n��i˞%�y$d����ܬ��u�+=�����g]��}�ѹ���__���� ��4.J����M�sz<��]��7)Ȝ�J�I`w�n��W�|�f���ޏ'��� ��9
&b^&f&$�yy�=�J��Gk�>I3�{vX���s�{~y[��9Q&�X$�$#<���^n���u�~o�$�'��"�����ۿϾ��מ@��1Q��$�:CpI��p�ݖq�����3%��w��@g���X�[��3�Mמضǔ��������x�eZݻjcb���7ZR�	�"cV<-|v�]�=�����L�5 ^n�N�[��ԟE!J �� ��n����6= ^wM����|��w0�Q�N8&�!IV�_�X:���}��}�]��ʚ��G�"�EM<ĸ�5���g}�zi��/z����Lc���><���o���rGND�*T�K��֬��@g����v^�-��ס5To{�����*�_��Ds�;���@o3���$%%ABt~)+	H`�Oǽ0���w���A�㐯S��T�L��@��(w"r@�FZ� NBP��HR L0JRa����@	J&�J��EHb&���	��� a� ��zLVA25��D�� ;j"�X��$��]� I�S��,�	�VIc���NBt���U�}�Rf��W�QO$��J��Q�9ͭ��2��T�\<��k㧆�n܌�>ѭ�vͰ��v���-�k���#p)Yi�cm�&��5�f�vwmصȏl�kq̖OA��秳m�jE���$���G\w��sݺ�n�q�y7TG[��0{�<���'#��uv�;�Żd���;cV�:�ⵛ#��`�M��s���]��]dqoAlvy���� [�s��϶��\�&CI��7C�#:�a�ͺ�ٙ�{G�v6:$Z[D�]6�a&8�7:^��u�9��j�I�V�'[`e�P�wG��b|z���ӣm�6�.���<m l\�r�q���뮅�l��紗A�Tp��E�<����gI��{q3�J��1ׄ���WcW&LמW͠�i9�&MC�p-���c��hȏLg�֝d�]�	�sl�Ir��f�:��i�N��T-���ٚy�F:�C����Z��m���-s`��%��V�ёs*ø;k��v�ػ�&��vNSu�T&����x�n8�6ƶ�J�����;v�!"zv�V[U���R�#�h͍����cuS��C�Ձ�wm�d�Bq�n�Sv�7s;m%ogD�m@�RٙT���Uų��mtt����n;65j��vz%�-��k���;kR	1E��Yy�X�[t���&!�`����۳l�%��;]n�+l��.*�v��E�7 2�nж����g6 ���'��j�
U�I'��HJ���Q1���`%+[��!5K̷	(e)%yj5;6��B�Ì��:�(�b3���V�6e���lm��8��۷$�t��q�����`4!^��PKkSb$�4��R{6��s�F��`��D��y��F�7Psݤ��j��ά�<@9�tn�*�t�;0^�r�)r��ޒA��Lk�tg�oWG[�Fsu[�̪�<�˳�m���dvIj*� �'E�ۭ�p�u�f����-��z[B��\�S����[y �[�Ə�{���������������q��ggC`g�x��>��P��A����v'�Aq����`� v!Ӄ�z'��X��j��W�D���0L��$S�>�{���wm����������p����gw�O.�9z�%vG2	���w5��Uű��<d��ݬ^3v�L���|��A�xtn�J�c��6��M��tF�z��I�Z��]z��Y�6��vچLv�[��>|&vR���n�I����W<�l Ř']�]��PlTH�Dgs'n����\�i��ΉAnڦ^���m�eg<m�绫󫅳��$�a)O�@�B���������>����W
�=�����.��4�L2GH�r�w���_�w�qX���W̙�$�㿾���Q��S1!*%K�̻P���|ފ%vӕ5{�ﾯ�{?-�䀪4�|�\Vo�@f.Qv�T�f����e��g�x���T	�a������y�[�۫=�A�I3�It{z(����D�v���@y���o*j����}�E w�n� ϑ�HӒ	SS�qFS�X�ɇ]�P/4:
mju��l�[�vḇ������Z��H�J:HRU��=�`b�ܻ���v ��@	�,���=U<oY��s��s:��<��s����R�!�O��@�c�{�z�˱����M@^�.z�5�: ������Bf&h;{���oR�I���v��w�,{u&�H�RH��s���>���@oG��8�������J��<f����b�*Dܫ��b��$^{f����{z�K���1��Xv��s����s//+�ݡ8�+�rU�����x�G��b�9E�?�|~m��zh��g��|�$�����폹�fV�Ҹ��"ARjE`w�n���I����P���P��zd�k~~��nQ	R �� �n�x{������2I�<��I2�:>��;�z��ĶȐ4�j:HRU��U��=�`^F���+�3ySU;�i��D����J9-��Ǻ�������A�ۿ��oqX�S�	G	P����T}�Azm[��||��7/b�vD��jwN�����N����ND�!q�~�߹�;�ͺ�;縼}_W�����hk6��(�rT˼�݁�ޥL�$z;^���k�{v������#ߩ��U#�T�J�7*�ޏ'�/#y��f3ܕ�����oJ�jrF���q�k����o�`{�}��=�J���̳���2Q�y�
Rar�3g~;QR��]�*��#��QG)H:MH���7o���Tz;^���k���j7�$���q��h�r�����>LҼ�	q�N��W*[���V�=��{�÷-و�0�Ձ�r��3as����.J��������B$)���aG�>�&d� ��k���]�3�z��+�^Իv����p�� ���Y�&ffsѽJ���zr<��)Ȝ�$n,�n��wٷV}�X�W�W�"���V��[Z���$��&&��eM@-�v�/#y�\������pɴ��.)��: �^^@��Fְ�C	ݺ����A-�M�Q�܇gk���W`H���r=·d��.����e�W'�a�8X{-�ݱմ�q7t��e��v�맓v�c^�
�o�=�G+J��&�y�K-���ֻX90�(R n�-�*�Փ��l�
�6��.�
���usìatP�:N��8z=���n64g���f]�̀�A�GO2���I6�JZ�2I^@�����r]�<<�;l��3�m���(ˋ�"m:���8.��Jr��R���r���_�^����+���ou�2fa��l�wԨ_w�rI��p%����W;����ͺ�;�_���UR=����hr(���Hx�%�Z{�`�f����5KH��z�n�x����fI:d^o[P�(���#y���]��p��R7%$)*��a`}���Vw�#��W`f�	�K���03��v�y̹�Z�5�8��bt�#�P��yl�*�+�RM5QPKD�TX���I+�3sn��ﾠ=�م��~M�m�r'!RKĽ��֮���^BL�v�2[,ɒu�3$����T�^��%yׯ̙����{O�u���F�R��'8�z���Uq@^l��$����T��JR�nVq������~,eB��1�I]��ʚ���8�e�B!�%ț��͆��{爈f���ަ�7����f��f�*�i$$�A�n�ǶǸ��/�vm�`�,�u�#$�dnK9�◬��YvG)H4ԋ�{�����f�X��+ꪰ9��V����O[��S LM؃=�J�d�w��x�w�N�������W�H�a��iJTm�I
eP�O��k��j�7�ܱP��I�����ɿm���˰3�J�����.��)D��y��,��=�@gwu�C緮�?R�~�,��r9ND�*H�V}��b<�2��R�w=�(�n�7���r��:Hm6���` ��C�k�mr�[M�s�WY���n�bu+k�X����f���*��Ҁ��k�d���w���5�1�F�Mʰ=�P[������`g��S$�n����j�qr���Vwwy�;�۫�=�X��)�pp�"A&�^�3$���1���J���t��ح���Ē�kLɒ�7�@_;��̑2����
bn��oR�?&gL��z8�;皬���p�j�V� ��(��N�Y.��N�cks���o���������iJTM�I	ʺ{�^�~Ǡ;��l�5��ޥT�n��?+��������z��ބ���])]�ټ��w&�����}L�0Y��r���T�8�N^�]���+j����/#y��k^��$n9%)II�~U����ܫ�J(��z=�"�t�4��1#��J�x�T�gJ�2�Y��z>߾�0{z����B`B����*�"X���R�HB�ʟ~~�f[��ݽ�v��sG\q\j�Grz��]g��s`3��n���Г�eo1	�Y2Y��m��]#�8�!�t�ÐӺKmsHQ�K;�.��jK�U�
jwZx�!꫞wA6�荖�Ͷ����5v��=:w!��Z�͟!Fږ2/,���p.�N�M���x<܇����uG5v�V�R�k��-�V����ww���}����w�7�c�(�o,ix�;����a�=�!�S��_+�i�m`z�k��<��T��52��3����Z���3ySW�7�n��a�j�n�R���$jE`s��w�3&=��*w���=�I3��k֒dq*��L�9��f�X�L(��������8�A0L<̴@�*����Ҁ�F�����JL�o*���[\�wr)M�"�8|�= �%vo*jw��4m�"����'$x}�s�a��Wn���ZFsiuù��v���G���m)m�)ȇ!ND�7ۻvo*
w���7���94(x��������n���U�k/�%�̄�3(TQIM2���1"���9�3.fd�}=_M���@w�w����U_$W�3��q��)NTI�Tr�P���{RWco*j7�)P�H�mP�jNY�;皋A���p��*�$����Y�u/�T@L����L��I]��f��ܽ�r�y��d�����)��"8g`�x���
g��=c�䜺s���O��*�:+V���HT��/�f��X�O�o?����=����7�y�`v yi��� x��w*E�����Αv}Y�W@fx�k9j]ȝ7���'�N�������JW�o�y�U&�UUI�UURj����&��F͟�\큙��h��fw��C�� ��MI��K�PrCzӎ�9Yh�0��_���F���Z���hey��k��ǌ����+{�Ï��M�wk��|��$�Y%�31���X��'X1��c�ޫ��3��+�8	�8cTM�g|�;P�深6�k��Z떰|�
��Xb �F����I�E�A��=�8v�i���N�@���NG|�.�k�	�� F��P�j\y���Z�3��J�@��6w���Ɲ���&�,޻�ݾ�����J�g��	����g��=�Ӧg=���l�Ӄ3��1�C�8��2;a�:v�;v�fCL�2��8�3�fqӎ���� ?p���p�(~�N$.�`qOވS�m `N�eU��B��' �t*g�<;E����΀�����\����{���X�~���δ���)ȇ �2�/T�߬����v�r���ޞ(��+�ͦ�1�$nI%9II��f�P}���y�@-I]�29җ��s�����ck4o0��rt��+��3ք�\k`��<NA�f؜������Δd{_��;z��k=�J��X5{)*��`�jNY\�y��}�}I�w��/E50�<Q�[�f�sK;$#��M��7ۻޔ�۫(;�X��+�4״�M8��*(�8 L�{�R�p�l�@{Ѻ��17&L`BJ��(/��b+�mZ�K������6بddj86'*�Δd{^���ou���T�7m�v�N�:�<�c�����r����	��%��l�6�P��d��3q�{���>���Q3�Tbw��� ���5*j}�
3�^��$��Tdq����&A��@{�:QC��퍿�J��Jo�RI�INRRs�W��뫴�{&"�L�����{`�%䙉�"Z]�%�<��?r�P�����<�~�_U}^�߹V�kW䤎'M�ԛ����Q@-I]���50��� ~��82���HHi4������������3�zp���s�s�.�@�:���5�s������m�cnf47A��C
 ���5M�'7���t��	x�r;�#q��sn֓َ���saٝ<�:lk7I%��r�O�6�/���J���H�v�kb�RRu�a�	�����r�FVP����͔�ݨ 9֞�]��]�nh�r�#��N.�(��m��ɻ�9�t�w?{�����{����c~�dk���=�[i��Q�V����es[�m��gqu�.�w��'��ui�&G�&b��w~�=�J���t��2\A���`w��LI�9REO�� �wR�=���ؠ��ws���3����m���)Q���'*��l�����}�7���v��MLgrxx���t܎%vp�������f�W}�u`s��E���x�$�rv��:Հ�6{��~�Ҁ��lR{��߯ڝ�{RWg��r�%q{b�G7oJ�D9eb�e���!#&A墪Z�S����ԗ�n��^�K,���2�ɛ��3v�t�(�*$ܫ����O��}�Hj2�`Xa
)1���x��Y��N�%�o*j���3������0�7B�w1��(�;��	��z�����t�d�q	�a�g�y{,K���Os��6?OEږ�t$��"��s�{3n���}���?%{W+�3�~u#��g��L��Yص�6�^$��6�)�l�q�ۆ#�^��8��M��m�}��U&��䢀Z��f����M@��ڒ�r�N���]���n�}�����T��ޮ/�I'I�s�އ�rfH�&I%�f6�>����ޥH�֖&F�?1�M	�Ͽ7�r�����\�s3i��I#r9)�I��������ڀ��‷�����fg�/{,�x�Dn����D����&꯫=lX��]��ʚ��s�?'�~�6���'b�S[{N��^x�Z2�/U��F����]�RI���q˳�GVf���Y`gr��ct���֗�a�	�\D�D�����5}U�����X�L*���w����;����i&���!���kR�5���330[��E ����+6�
����t�����˾˲�܍م@_{znÙ�4�Iq��!�fWѫ0�&�B�iv�L�-iL�4����;�U��%��m*@w���E�MR���3�TX;��ޕ@	��{{���Ԩ�Ζ�������fkIB	�D�%(�CT�z���G����nk����h��P��%]�-���	Q�I	y��?�?.���M@�35k=���mkzԒF�rS����A��m�����ފ`-o+��ߍ�3D��m�n���@;쟋 �2 ���s��ͺ�����JI"q�܎9�,�P1ky]��r��b�e�F�q�AH4I�7ٷ�6�6��y��4�lPƦe��2v�!0$H����>���fkv��۳�\d�E��]v;��A�ԛ�m��ձ��]�]��.�9���L���<H�k4��oo���Ջ�9RgmR�*潡$&C@�8lg�3[C�磍aے05�ǁ4niѵ���t������2v�e���ͥq���A�g�霺X�UWt/G=���GE��jܬS{�ۻ�i&6
j`�(K�Yy������G���ߝ����;��S�Wn���������:�Crd`g����W9�m��i+T�"��MI�C�9/�W�~۫3e?oEkR���Ԑ�ĺ�Dt�ܫ����Ş�e�s}�|��uϾ��g��/Թi�q:NG��}�E0�+����;�����O����(ҐT㈄JGa�U}�T���z�yz��͔P����@n&%$��� ��5!nmՁ��i`b�c�9���pG�i8��P*JjQ1n3���{Z'2��kK q:أ�����4}�j][�rJ��A7*�$�饁���@Z�W`v���y��x�5��y���*�>��p�:<@��l��� �_�v �t�P��(�����		 �$����7�=�K?��U}��̟��s]�G{�岔I�"rt�'8�}��K���8������o8p���� ��RN;���30�͑��@g��]�����2���~+�ꔡ$�iӔ�2��7�pstz�5k���ph�t�6�ٺ�^��U����ݾ��뙉�^��5��n�]��(�36U����%D�����JG`s}��	���}����‷�lP�����$m�%I���M,��K?�t��Fk?2�E������ |��iQ�QJ�{��W�~�����ͥ��nIBR��!�X~�������c�Q��+�;zQ@[n��J�Iێ)�+�unk�?UUU|�L�l�{�XoO�y��m�f�R*e=�����l�½��8��L��B�����O^oE�g�f��6�1���m���]v�g�@^vӌ�ɨO�ؤ�庢MI�C�99�3ٷW��#�����s��/���y�f���Cz�q��]��t�2��� -�v(&E���p:��n��=�Q�I]�i���%vX�� ���X��*ʡ�&_	�0; �F���@6�q@�e���U�νXBHG��8���f�y{z� �=<P;��7f��9<H������6�rF�z��)�4��p� =�v�=���*F�%*N	�#nI*F7;�;�Y�(|݊`E��`g�O(���(��*	�X練s�s}�|�ɥ��y,�	�rH��D���c�QL�J�oϝ����c7��ۭ�8DHG 'R;]����3[P"���̙��#��@f����xy�NA�N>W���۫��������޻Z����M�����)5����1\�8<���C�;ahJBHSõ5���[�}�9�k��%&R#�͇9��MD��gQ���Bx$�t������խbk-�ۡ5y�8��hyQ$�w�gYg8x'�NQ��)ǋ�I���(V�y(�d҆E���G|^,���秺t冽���nv�\<��G���KJ�wBX�3Q�ڵ�!��=��İ:щ��נ���[A�!ҫ�������o�pb���d�l5�pӠ�l$1����eF�̵a��E�0*���T|PP���U���Uj�$�14�-�6�%R�@m�i�U�T�î��,��+�]5��Yۣa�-έw^�yѸęe8��86��e5u�r\{<���z��n�W���ۃ�v�pX�:��jěl�;B�\��ygJ������8����wh�@0�mҸ��&��5&��s�7j�zf��|V���v�زc�wJ�
F�n}NW�We��[��q�/�q�V�7;���'e��!Cs;�p]�v�Tq��[�iݪB�`vȽ<�G������%6��'m�V����f*e����s��"�v�npћ��ȍn-:^�zq��f�۞ݕֲ1̝���sV<:"�x7L�iU:0���ɋ�Q7M��N-��iW��Ǎ#@��*�ga�M�ʗeP�2�βk����	��ZR�{v�}���c]��n��^�睽B��d��%VY��"��P
�pR��-���T[]��i	��E�tVq���tx��W�mv�ftH�S+�;t�msn5J�v�)����b�W0���Q�@@8�r��*c2P ��nR�@!'&�cn,�;mV^9z�U@�b��^+S�Q�!ð<[�T,\�nH'tWOUi�P�]�f7&+��4�-�=�0��b�N9�ݪ�a�I�45�6Mu�P �l���vejt �Aŗ���3�nF��$%ʃS���� [Bޡ����%�g�ձ6����Lj��m��[sen�)W�
���:1�
�^g��"�Pp�@�`�Zt�N�i�#U���q��5#`:&��d���T�s;n�ٓm�뫕���7b�a�g��^�p�㰨t��g4�Ό����7����P8$�����4P�e@x��蚴����9��g�r��ޥ�����isJ�L�����@�6�Ŗ��%��x
T�kj��dԀF��rF�)3%r�� :m��a�
�DM��f�����U�	��:X��ֻN#����Vi�����q��ݢ*��/W~����@X��'����"���G�;N��L@�HPG*���e�ΡS����6��FTT#�kk�Mv��$mI�ۮ�91r\�B�F�N����,g�K�;U����j�D��>�᠇;O��a:A`wjp�:�d|��-m]H�g�όݽ����c�L4���՘۫�g�,Q��͗fJ�(e(�L���B�9.,�ݪ������N�Ӷ��V�Ǩ�pW=��3�7M@S���jtnϙ,������}�u�����-�b�"wg����cĸI�6�<Hb39�]nqtXp��h�:�N��W���J�7b��޳�πfo�=���J�;r��Į���QT�f'�v0w%M@^wR,��D�!q�%q�Q��[��f�Y�.�'�����?o�R��FܒT�n��w�5����;���[����J��$��n2HX練꯫��Ԣ��r���(�<�}�2��y����{%ek��������v��r�S�:S.�+�݋���0ܟ�6���b��+1w�o�c_��([��ޔy���3z|W;�I�Fԍ�Rr;����eU}�Jd��3RM	2T�<P�(|�w@sږ�u�8�b1���d��͔P����X�r��Q�Tt�)*��}4�8����9��� f[�Ԩ&K��\�T�O�fb]�R���^��z���ix+Հ��
��**$�����*9z ���.��'7Y���n�n0.������~`���$��/.�LP��]��ʚ�k��皾��n�
7�����䑷$�#����*����נ/��v&f1n���NJ��� 䅁����u�/�zO���F�ү=1BB�������ѳ��7c������"^^n�3?�W���r���QA��������`f�["�"B9JB)#��J�
5u"��ޔP��@ww��������w\nͰ��6(�����ȶ���U��n��7J�_����ܠ�f	!D��ՠ=�<R3������M�g�޻�x8C�H�C �%�����|�v�O@g�޻WJ(sNe�v�'nS�2+��Vy����p�_U|��������x��9RS�0�^e�_{��v�g��fff����A�"h1W|���r���0�V���6䒤cr��&�<����^b�9[���A�U���1C��
��q���\�a1t�z���wfu`:w[^!��ϥPI�B���jHXQ��i`{�1XZ��7���4�=������#r%��;a'�/���Ҋ�e��﫭��-�G��
B)"����w�Ԋ<�}�|��^(�I����7B1���ʚ]��i`nG7=y��ܽ��7���y%�$y!�x��͔����ky]��ɥ�
�����koGC)Pܒ4�ᒷO+B���K�v�OEץs�;��bg&Ր�z����ʋq�ɖ�Ł�C�쎗�x��&��ɨ���gsg���Oh�3h9�XA��+�@"�i�vݷR�7n'�J���ԓ������u��:�9��9tX����(��$���fJ:Ŝ��'IN�v���2��VO.κ�ݭ0��#2�gc^��,�.;;ߛ��}��˓~p�^�v�݇����ò뵃�\՞�-���X�qɹ���ֺw�C�4L�K�Q`%��@^�uv��W�C���i`s�'*JrF�����7���Q@^l��Ξ+����y�$������g�w�K*������o>�����)%%��ԒPS�ή(��z3���[�<P����Q�$�m����U���m�y��x��������<���K�F����Sh���Qs����}��Z�̊��[4��I��r:�%!%E )"����� ݼJ(�(��n�'�;|��@�0LK�Bxy�V��\S��70���L����`|�;:���s��1BO@-Ԧ�m�MD�IC	�e��27^��:f{���A��~V�ڶ�9j�*�8�]�(=��f�]��	=�Q@n���2�5%9#	"q]�w�����Y�5X��,��+ۆ�Z���7�J��^*ڌr�N�Ŕ��%��-T�,@��XEɞRRr8�rJ�4�8��U������^b�����p׷AZNJn6��z�J(��2;���\��݄�����'��8䑍�✲�W�]���}�V���	�.�����5��YĖ��U��~O*DHI 7#���c1�+�7a'�����}ފ�����bd�H�����=纬�����ؠ3;�����xb8�q��[,2�ͮ��B�H��':؄6F8���)R��*E� q4�Rr*�;ݚPϝ�@f$���I�����X��S�2+��y{u�RG��v��U��xB��U�'��I"����J��I��(�3#���3�NGNIQ��� ��i`s�4�;ך�̗	B�I�מ��������e
7P����f�z�1X���{�4�H�V���U�@�mW%g�����nМu�]��S9K�ͧ�#�.�k��"8䑍�✳�f<�`w����f�/�}�;���`��cz��$$��&^���+�7T�����̎�3��뤓R� 2RjNp
��i`w�Q@�dw=���N8K�I/�2�f�����/a'�3<��纬��k[Wj˧r�5vp
��O@�bJ��I�N��(��y69zgN�9#sV���gs�7�{n�g�lq��3pn�v�8v�Y9�tr�O���F��n�n64s��(:^�ڮzc��E����ϺN�%�c^7;D����I�p��K�z]�N��<`�Le{.�a";n4�S �`X��{9Ld8�[n��b��6���7+�<ZQ:1�����m����uګIa	�؅Y���m^��w}�|U�#'H�n�~��m��]�|�ܽ[���g[���+���\=53�s[Tl�.s��ߞ�[a'�/����n�	=�?R��7��$�Ns���l5X�x�3#��q�����3����=;��(�mB�`wߧ����ٵ_}I{߷�9�o��`o|fȆ�)M�✲��Ԣ��\��݄����(j{g��"�) ��v{���%���=~,�O�;���77r�rd�X��<]ƶ�aHV�Ӹ���s�ܑ��-9':��5%Ii��MJ��I�9�(=禖���͏>�3;��A���I�O9�n�k(��w*￷��	��0���Y2J����獢({����t�_W�W�K�g鿣o��r�һ8c��3+�7T���R� �3zxi�T̸DLK��2g�w�bߧ��٥�޼�`��29SjӍ��S����3T���R��-�z(�If��~�v?���j��%�����=p������c���m��gX����5�a䘉{7�‷�:��r��;U��=�GM�$q�9g
���@f.W`v�'��J(�׎��]�D�JA9#����f�:�7\�e��]���9�s���9������X`��5J�#)��Y^~~�Zޏ+��:4'D�2��kl� ��3g���,���n��X��da�f�;:R!�[;R��ae��&Y1j�A!e�F1f��y��y7����fXY��5�f��`F$Y�����ac6�:��"b�¬�30��+33
�� �,2�H�K{�A�1[���#(��22��l,b��+�a��fYX�j�e�n��neİ�0���231��A�[�(�vAC1e�X�cb�a�	�4ń�Fl�Z݁�Ae�8�DNK��f���c3affSgc�]p4���i�� ��$gw�dl�N��e������Z��f���d�)^k�c`a�Z!�6��A�0�g;����#;6dT���0Cۘ��Їb��� �,ؽ���p�v�`"��(v ' T�|P}�)�;�oo���ky6�^y��wV�i&�J��"^�����5o��@f.W`v�5�6R#pi���V��8V�7S��;c���|��C��܇�K#%�Ӻ4�۳&r�/a;UNFENM���9���yI�6�b�v�#-�8�Wg@��EK�.Y`f�'�3[�ǧ� |��B�*H����f�#q��V}�~,�����#j'��$�Q5`��<���R� �ޚ1r�2�)"N6�����T�����������o]�����b�8��$�a}_}��_w�&�V?_��28(4�M����������{ـ.��3���Ֆ)*P�6�4UO�:z^�P�@Waަ8uB�<$��u��0�l13.�wKL�34bJ����b�P��%��կZI��r��6�� �<��fI�!���@/?v���u��$��/hl�e"7�
NE`wߧ����dP�����w��`.��5w��	�"`��w�,~ފ@,Y�z��o=ޛ4���cBt�����w7� �F���<P�f�DJL�S���S�L�2�12�,�M���U��**r�R���Ƥ.3�<lb�6�<$ɱ�s�
�,Z��lvѬvf�mr%�z99</7��x,�v�uҮ��k���\]Ae�6R-��ݩ�n6xص��O"�`�պ�l�Y'�g�������ڔ{]`��N�����
a��v7<t�+K��M��m:랟h���G5t'Yt�*LN�ՙ#��'�Y˞.���E-��{����a�j��}�\��_v�x:��dն�C�Oi�� �=���p8.�����Y��^%`�O=x�1@v�E8�b�� �{+P�9"MFB7�����V��1v��;���S�w��)�Ò�N8�,��f����p��V;�K(3��#Q�Iԩ�H�?>fo�w��c�^z�J*��|㢃�s������'(i�jN�
�{�X����x�1�(��r�k��~�y���.�&Q[��q.R}��N$1q��n��q���I��6�Dn4����f�}�4bJ��33}��y�� �g�]<�RD�ː�EӸgoMZfR��2R��d��lv]����t{����Ą܃R"�X���g�j���I{�������,w�֧��$�x����|���y�}�w��37�������t[���In2����'��:h��+�;c��[��z�h��mu�#�v��&26���7*u;b�Tt�^�3٢��"ᛚ๫O#9����m���i��I]������[��;�@-鍑GQ'R��;����~�꯾��7�y�|��-�z)7���:�C���KD�^C�݈;c�z:=�G�w�0&fL����%��|����o�v-���Dn4����UR�韕�չ����%vlrzV�C��x��be¦����t�(ĕ����g������?�>�#u��a�%��<.�=&+�b������Jݍ��x�u�,�o�-:������8/f������<�; �iڒ'��N���3�׾gs}�j ��h�%w�sY&�@�$Di9P�qX��� �{%����p��Vw՛(R����q��j��3}��zh�{�clrz%���������X�$	hI �H��0������fjfRҙ2;=T��r闘���xR�H���wR��;c��1�5= �����^3I$j�)��b�����M�6����>�t�،�u�-��t�u�}���.�Q��I��y���j�g�]���8�k�B�Ӊ����Xש�`����p�T����Q@��4��r �k�unk�'����_��睊/c7�=���`sǫM��"D���p�W`7>�����ϐ�Ah��K�~MI�IJ&��X����K�N�������������d�J�	B�)����f�o���)	q�}tۊ5��Km3���)Eb�+�3�ă�	�����=��C��|-�n�g���s��~�m��f1)-֊�6l�tj'��Մ8'��q���58��W1I�7�Rg�j�>8�f���[��WA4�+W�,F��x���u��8�����2n98y�������4n�q��N��z�Z-��NR�\w�������[Nv�[z��k��`N7�x.��U�5$��![�[���<\��T�!919PLq��?��g�XQ���o8b�k�����e9!J&I��{r���������vt�k���̸��$�T�rGt����P�S���_#�C���J�D�'8,�v{�j�8�1����pz�i���M49�7T�{%n$����Q@_ȏ������L����{ n�]���#m2��k�O�����N�.���q4M=�s^��7W`��ܢ�Q��>�kՔ�nFI#R;8����9�64&vL�eL�9O��@�.�k�����*G}��~mHӎIJ&�� ����5=����^$���Ԟ��`؜�CN;�����,�v����~������=��t~e9!I�K�\%�J�P�E�S���殺Q���lB �p��PJ)'L+Nz�v�D�9v��Cs��U`���gquʝ4�LD�#��Ł��z�~�ft�~kp��Pf�����J�4�'8�dHќ���q%v|����SDC����:=�@[��Q�`d32Rə�]&�z��_w���/��]K�J9�\�%����{w���5�~����?*���i7#$������7��[�������߯���������F�q�ꓖ�;�qe.�C�!�LX0��8ؗN\���+Oj�x&�~�tjz߻���I]��ܚ��$Di9P��`w_�YAŝ�@n$����Q^��o�a�[�1�&d�hx�"������J���Q@w�X�V;�8���T�rG`{��]����H��=Bd���2fe�fP�оh@���ˬ����_��L�"PӦԜ��5���Vf>����p,�Obm���RAJ)����6��^$�'�';������S6�󹭍�$�������~�`qfc�Kݭ՞���;[�t�b�i��f����IE�����E�5=EDׇ�NH�q�������pY����� ᙎ��ukSR�$���n���Q@b�O@[�tP�J�e��&)"#MʄR;�������`{;��_w����}��I*��IL��.*�<� ��ȴV�1�Jh�
)�212Z&q!̢s���b��JB�bbhl�H^�j\���������o�vv�Z\=�d�ș>�y/*��w�W�R��)Q��	�/�H"�C&�5N<ZE	y�fKz釵���f�c��������o�do#�����,̚n��\̠���g�QΌ"�uf���~fV�� �(�`4^E
[}atf]�'��JW'�w����\T۝�F�;փ��3}f��13�l,��e�ww��۰��8{.��;���ճzw��dM赣5��l,x->�$:��b�����4h�-Fh#]�ٶ4�A1�S�*�Z�"�;�㧄@�!:wtHty��Q�ۥw�xl̠��xhCe�\K��;�o7�-`cl��`�r�h�k3D]j�=�5��ּ�ḏ����4h��Ɓz�iD�h��&������2�*u������3|0Ch��qW (�|�DDt���ܔ �9Nc�A�!��XML�I�M"e�f1 {~�W�4j�F��<�;����7m��`�[U+�a�$٤��d����خ��A^L���g���k�j�s����.c� ��$�@�A"Gb��ZUºJ-��4�����[nv��t�v�G�,�� 6�ښ��3#��؁Fk�Σ�7�q�Q�&�:{�lg�d�(�q*���lS���gl��}\+�;��i ��qar��[EnŻN3�7oQ;s`4�ذ�֥.�,�{(���m�����];��cn�=��9����jz�I���p�;�h�
g�9�r�������;dӎ�M�qզq��ª+�ͺ��I����n�s�v��ci���<�vxn	.��m�@c:�\��r�r�!ֻ��u��RP�H�	A�ѣm��2u��.���S���¯l�R��<�x�́hqq͕ ��g% �GEJ�L������PX
���3��?+���'�{8Rh)PK��p����m��-u�3���\��sj���1�b��ײ]���v����93d�Lf���Y�j�F;7�n'<k�,��l�)ق4�( ,� �љ�U�Х�'��mΜ�N\�)�s��Ma��;Y�v�˅��g��=��^�H��M�lF��ݱ��^��8��ca6�ِ4��݃9ή��5X�Tj�.E6�,3e���V�@祎��n�G*3��y�����iN�c4kB���WI5 ����"��b��4IW����^�N�u|[j�vY
� ����[p6Z�*���6�� M:v�[l*�j:1��!�%��n��H�j�
��+��l9=366n`%]�̖���_j��%�@�<��M��˴�8`G�'\sM����J�D���� p��έ�lm�P��C�J�vC�Ʃy�9ڢ�5YxH�X���m*� q�3g��t��t�ί�b��%y��W�D`
�W1���8�7$FJ�9ܢM�o[%m������ �vU����4;U*�bg�&��I�)�\�����ww{�@���� ��
'�����W���CMϭ� z���K����A�����\6=��~���5�t:�s�6���7�lBn��7+�F-�H<[vڶ�.d��ZQ�r��u<��[��k<8��n������s�ٝ��2@pH����\�a���Κ���A�c��bX��h7&e�v�Z�fQ����W%�Ʀ��t�n4�Yl� jC��� ��#)�S���-���첏Z��5�� �Zh��d��-��\�9����������{�~g�~~iHy�o=8��wc������Nv�9�8�[�����Î.��y���;1.O��)�����@v�W`s�(�1F�`s�X�TN!��T�jD����9�1{5���V{���ORI�DJt�qs�b�k��w\�g��W�unk�3߿~� ��JH$�����Ձ�5=��oCP�+�9��P��%��r�˦��jծ]y����+߿~�@՛������5@�R
I�!:p�e3�����枞��h��T�]2Q&[%u�J����F��) �o���������� �~�`s�ImE �331//v��f�ol�J��(�t�7&LaES���;���뿒gs������
&�A����?+��c+�����p��V{�l�n����0]S���������z����o�{����$�mkucN"A�T�rG`ny+�+�y=��;�����3��o��
�z��׶���U��j��,�[j�h9[�	����[��길G����9=�5=o������`j+��@�DR&�
NE`w_�_ꪯ��Q?oE���v�7��I3;�I6�h�ɼ�S�Q.4��4�J�L�&M���32Vʞ��ߣ����,M9N5rK������uY�/~y�X�l�9�Ԗ֨���ȥ�n�[	=������{ ]�h�n�j=����A��Ө�87L�On]�q[\C�ڂ �3 �7�u����$�(�dqX��VK�X������V�׳e&���Ȕ����S^���@���<����S�;���ݱ�J���rK=���纬��� �{%������Jr�N�R]�ə$�l���.��7��٠�J�+�`t�Ib� h�ѥ5ш��(�x������^{o�������pg���#�{ �ޚq%v	�{���+�R2"J�Tn�*�)�梗��3N���kG��@���5�:�z%s����}��p���ܦ��I]��J(Q����=�NS�F���ww��I����Gy��zh�0��̎�̼MD�8�f�u�U����H�͖{������n�Ғ!D� Ԃ�ש�~}�7W`-R�1���3-2LL���=�.�4�$��K�t{���k_!$�d��̸b�8xخ���_l�m�MǛ�8�����"���C�;�'_�Z��rަ.�h�p�2dݺu�v�+�Q��<�۰��ے�s:Y9��<;�ݧ���1�{C���G\��݃v�k+��۬W/��vc��qO�՛h�GJ��d�A�<fM���;] QP���<d�k�ֲ��m��4�j�;�+=tF4��]�������o���`�sg�\\�up��lr;Jv�nGu�:v`R����w��-�.�s��334���v](�1F������5c֒rH9J'M�9�7^j��ԑ��<�:P����B�����6�eɘ�"fe��w��;��-�w����y���v�+h嫻N6���%�/M��z����~7�3�����hn�NS�)A$��������[�7�ڬ;�}�jm�B��8�|�˱��j��ti�ۛ��r���y��.���p0(�EQ9���X��V�̖wwy�;YOu��$B��A9
�篽TP̼��5�fL���4���� ��X�fj��) �>\��-Jhĕ�����Q��Gy�v���t�$%H8�w��3�7vYVן�Xw2X��z�M7)K�D<���Q@{��Oy�jS@g{��p�V=��E)68��ʦ��S�rq���lm�q!���1��1�b�
��`7�"!���(�����hē_�fj��?mk�Xz����wc��[���4bJ��(�Ƨ�Y�m�u(!$��3��y�72if!B'�$
s����]tW���ӷ��� �%����7Z��TGn4����K:��;�,��M��߻�=[O���F(�di�<�=��4�J�SE�	��9������2w<�0c%u��i�S�������جX��8>��U��j~�?6�M|��wJ<�}��.������WN!�5*A�$�9��y��I�g���y�Xw2X��6�Hi��J&�3v�P�����h��љ�E"G�
��ﾪ���Ϟ�����~:�)���rf�d�H	M:�H�0p4;�(=��}]��Zː�QDL@��{�Ԧ��I]���ljz�s��Wčћ<e�=��)�=F�*�\/gIw'c4.��"z��4.9:�4�th�? b��v�P�����h���j�AQQ�Ӝ��4�3�ڬ
3����n�9��V���J9�q�RK�������4���trz3MZ�7JH���#����춑���p��V��Y�?+=���CR��2D�I4�%v���c��jz ���-�z@�"H.j~u�y[�SI�up��T+�s��Br�l��/.b��=��dɟ/�]^WF�	tW�<W]ub��BI���}�>�/���KA˱;�փ��Ę![��v��v��Wn�-�n��v���M�<�h��fs��,Q��ZeCeh��+#���$KU4�(�<r��koj�rny�h�q�V�僶�-��9���L�����$l�e�bTN$�mI2��L����d��K�Z���K�:�m��m�G����JF���nsu��t5mJ���73�~��U��O��>oM��K]���҇q�����$�/�S�f�����zi`{��F֏��Zq�-���l�/W+�p\���5= X�ϼ;�̏,���z�]��z�`_F���Ϫ���f����~MH*#�7)�9�����6)�=�-�4�]�M�n�)ʉ�#��AL�H��EI�����u�Ԓn��Tk��<NG�44��"d�1�<�m��kz��:g� ��cZ�RD�"wqp}�/j�漢�Jx"�
�*��W�ﯺ�:���矵_����6.�mF����0L$D́������P���(3��`gkVV�hi�*":9��Ҋ�5=S�voN۞f~^�e�pM��6�D�ep�9�ڬ��r��\����E�n��S/�@���	�<����î��\ԛe�T�rg{l���m|�`�]
���h-����9��� �/N�y��8Wif	5 �����/W+�5t����O@��C˽�-�mH*$�'��=�K���FH���D^�J�����)@3���1��'��?*!��=�
����\CK��fh&�-�J����4�`Q�af�����v�����v$Ed�׽<�2������@�C=����l��vu�R��@XZ�V��<����"n�D����DI��j��P�.�ps0�6�& �orq=�;���K��z#0�S,�h�:M�Dބ�;0@��b �����4A��f�:Sti���
������lI���ey��#�:���zo�E|�`SM1M����`�

B��"ZjHdL�2�u��4�T����a�<ِ��f �F�Le|�CL����oI�=*8�$Q�1.�� >t.� >����T�m@��Ҡ(�r���WB��T�gw@,��2hd���՝4K�{�����T;�r1D�#NB��?j�w0�=���>���~w����?3�j��(��R�9�M��`�Q@_F��
��4���Ӑ���(�A<)�rr����b�l�4�ƺ�V��c$�L14��w��%4P	i<{�o�kp3۲���~�CM�Q�Ӝ�ܔQ��T�@��@�tr��|�;�ޏz��#��@�,��4�
�s%���W`j�E n���L=UI5�ýI`']
hm\��\](�=�|?%TKMBg᎑��SB��J�]��t)I�#�hB�!$u�$ЀA
��sP�P�UK���.Uy����ܒ6���`fg�|�[�M�ݘX��,��+���$��T��>�ɗnNj��Ŕ��r�d�Qn5�"(�az�u2JQR
�"�Ƥ�A�����7�0�-�����[��^�xިwg���a�d�x�(�<W����sR�y/]��ɥ���k�YNH)C�S�� 3R�r�y*�����Ao��EK�r%q5#j���U}���������`s�qX]� �kW�)D�MJ%7Cx��3���/�s��tH�z�aG�QОǲ!����ٽ�y��F��7ݎ��j#]jV^S�©C';��m/N]F���tgu�7��I����>���mƭVoR��*�Y튁�i�vV)��N3e؎0���۠ͬ88��3�S6��}�a#f{]��Q�7a��ij�fꕉ�����b ь�ü[�u�x�-ԴuGT���c��Rzl��	T%L+��GFKUX��{������w������8{;MŶ{n��6��G���s���À���njź�v�3l�̭��� {6$����͎ﾪ�W�?���[$Ar. g��/7�vou*^�k����0^]�;�ME)J6��X������K-.c�V��s{HYX�q*JBG������/�s��D�x����\����r"4�#NB��=�`�8;��p��,x���j&莚�Rn&:ls͋+�۴�cu�6{0+i�Z�p]#W�u����48E-��{_�s3���٥��=�`w��j�N$�ddC���{��u�@%�@^�Ĥ�㓓4P����ؒ������4��Jn���������ң�� ��g8v�f�1�*����gޟ'���w���������	���&��p������]��٥��qX����f= �q����
d��W�m��]F���%�5��[�eHT�����)J6�����8sf�1�+�w��,�n8�%!#��7`g)E|й�s�@�[�`�ksElJ8�i�F����{��+��n��x���G�5ڠh{?s�8d�X��l��9$C�����3z$Ż�`g�x�3c������jD�N�"�����~���z�X�<��/z$�|�}w�4L��2�ռaC^2��ayRmt�]qs�+�m��6�m�m�7Mn����ḹ{%~~m���r(�\�{�T�_����H�PAH��'����{��9�p�w'8}�K����и��\#Ar. w�H��vj�Pй���n�%E)J�v}�����A�{���v�A�׽" �]�Z�[���-�n8�%!#PNs�w�4��~��O��r����`&����=G��a�{N�0�������um��#jM��}V0�<:�9�B�$bpL5�k~m���w����@��u�7���8�o<�9�#Q5-��s\8��fs�w�SK����W����36��jD�ND���{���8o)��7��<��w3�H�W���9NStSNs�wߦ�1�+ ��9��s�wq(-e"Gx�ǉ(�\�{� ^.�3SJk�c��RT�d������Y7I��a ��v�P�s�;Ol�p�1&��=�;Cs�iw�:維�>���>[�h{|[�[�q�zn2���6�i//Mʺ���}��ڱ�s�1�#�m�%��ـsNt��4�:^N�����W�]��˺T�m�۩��%����9Z[c4��li(�uI�	U�/�Ol�ct;9%��F�;g���u�a�n�dqs�b�ï��{����Ͻ�>�;~$pYy�IN��YK)z}c�N��s����N�k�t�q�`9ڶ����Y�
�{ �tH��vo���n��Vҷ)�I�$�PF��=�ۼ���,�Ŋ�9�poP�+�$�q�Rs�w�4�K�7�{����9�A�ٴ�ҍƑDi�X׸�ٱ fw��szx�/��s˨�y�3174�ڢ@���|�H�-F�?/{V�H�*E*DO�&���J�`��4��[�ֲ�H@�Mư�^�n�ZB��Ȕc����s�w6i`s^�v��q�=�V���DJi��8sf�u���?��C�2�	#+�T�y�� ��&P̅�}O@{� f}�4����!8X׸����s��`f��@�G��C��UL�C�L�����3����R��.z ���'(��@�&�{sy�;�X׸�/b�s�֞ARP�J)Ӊ ��v4�zɫ�\!t=���t�y��"]+Z��5 ��5"�Ns=�,�9�pV�@;��s��~�h.R�ƔN24�(P���s:b@�[�`f�E���EJE%H858�p^���{9�*�1H0RTSB�2�(b@�JI@TEQ8PP$Q@�D@�XQQ%D��DDT���4�.È`2� �2�� :-�߷˕w���X�e;�IQ�Q�F�{sy�;�X׸��� �[����R2Z�n��R��.z ��3���U{�?~�$*|����
gΓm�3rq��˸��nq!���.�]���.�][/C��r�$�|�Ė���z ��3=�vjWV~�{����܉�5j.ZA����I_c��j�.z ���x"%���	������1�J�������(7�$ed�A)i����W�'����w�‷����|��&��2e�����X���w��w&%ɇ���/����y���vjeTۛ������۫�p�Y<����&�˺�(�Ss����/0��??	�m6SR6f�����^ww�$����|7�N�ypQ�Q�D��ٷ�*�~�u���_=�q{2�["��4IR�i9u�����Mz2���]��_���[�ڒTO�B��ə2^���כҮ�ݦ��z�6/-\���܉���WN�6V��������a^�ߥw����o�Ff�As�������e����E���s���T��V%A �iF �iQ�@TbUh�R*H- ��1 ��""�C%biE�hJ
AF� P��TA�$r )�$E�P���IH�*P��QJ2J�H�4 2H���@)@���Ў���( L��A �% B " nU�B��@�E iUiD��(T(R�J B�P�QB�A� �	Q@F�)D��F�JB�(E(U�A�2%E� (�P(�T� (��UR�JD(�Y��i"���iP:@��>ߟ�EDJQAh�7k����n��P� )�?�O���*�������������?���(hhJJJi���(��Ih
U��(	V�� X
��`
����������A��?J���
�S�����D��B*s�����I���������/��
򪪪�*��������������            �����j����������� ?����w������#�����A�h���a���_����DU����@PD� N�����{�aC�P?�{���#�����?y���'��@E_����[3��O���_׳�}N?����~����A~��� ������?�ޔQ0P)Q"U�D��HQ%�RFHIQ!�I!�X&TIQ �TH�RaQ&TJ RIeD�AI�D�I��TI �H!AI	Q%U�I�YQ%TI@�RP	 X �RHQ d�$�R	Q&TI�R	Q !D��eD�� ��AHIU%D�BTHQeD�P$�D�RRHQ!�EHQ�R	%�RQTHYQ �RQQ$�@eD�IRd 	��!!` H@����d!I	D��I	��Y$%E��E��BT` ��$ a$�!"BHI�� FIHd$����HI &��!dZB�i
$"B$ ���%	HP��IBB@�	��B ����a!	BBRFB@�e"RI		HHBP`E! !!U! dE	I$%HIIFU!��P�JBa�(Bd&B J Id!HE�$ ��T�$Q��P�!%a%!	H!	a 	$!R�BRTe	 d%@ HE`$T HD��$XD�� �")B�h%
B�)  $I��P�$���X@aVRU�%FP�I �%	�%�BBE`H� �BDd$ � P�$T�$E`ID�$EV@�YB ����@�@� P%Q	QIBT!	�%	 �%�XBHB@B`I$E�!P�IBD�!�a	F��

@�P�� �$	F�%B�Y H@�eB�e	�`I@�$YR�	B!� �E�IBYT�
�H	FHHF�aa	QIFDD�FE�HBE�!X�iT�
Q�HA!Q�%H I!Y�h��a	F�d�A�iQ �!D��m�o�����(+H ���|8}]�hv~��?������?���ts~�����>���������8��濉�H "�~�E���_���G_����t�*�W�������?�@E_�y�X�PW��sF���3����xo��@�(��y�v���G��]@E[��_����?�� ����?�v(A��;���Ӣ��?N ������󠀊���( ���������g�6Y�3����O����:/No���]~��??q�W��U����?q8��?����W�~��������?o�"*������O�?Ȁ�?���O�ע "�_ч���c�������PVI��VF���/sV` �����d�Ǿ�TU��*IJ! �A@�(
:�S��f�5J��Z
��zzPh+�!J�UB�m$��ݺֵ�z�
J h  *�T@ 

 T( ��� 
 @   �  &�@T
(����      n�U�P��)F����K�z�]����U�ۗū�k���j��|�	7�j��|���u����w���l�w�
�{�S���j^�u<{�9P ���u�'T�yR^��+=����޽�t��+����u[�y2��wԯ�.�J����ܽ����﻾�� ��� � �ѕ WB��Y�頽�( )�f���s� =�p)Ҏ��j� K��F�i����y���P)�wUE�p)Jw,�
S�� t � ==� =�zjSݽΔ�Y� w2��l�OwqӠ�T!� �� {3@4��Ҁ��  {�^�w�[`hQ��W�w1����ON��۽�>�����w*��޷J��k=;�W�o=�w��]�u��=*��S�{=�NO��޷W�P�=����u]��>�;o��NZ�j^X���x|�To�����+�X�|Z��.[ϳ�^(  ��(4(-�Em�n;�
6y�+��}������}�W�NP�>mB�yS����Kf�{r{=��Ҽ5z�eޔ�>q����_   ��ܧ��Ԯq��	>�*ž���uxm^�u/3��P��ljK�R��������n�_w��_ ��)}�R��4�((���-��4z{}T���Wz�^������N�J}�<��V,�i�ʹ��R�����K�=�{:�   ӓK�w��_z/gz��{�j|���^�:^��ܩy޾�v�����.m\�{���w����_     �m)*��db40�2� R�  Ob�QQ�H0@i����������@ OД�RR�  "$)��(�=@ x�����������9�Rw�gG��w��tW�wO��T](�����T_���W�PTX�"����_?�,��SJC����b�W�,�~v�C=����>\G�/��/j���s�$����'��Ë��{|���S����YΉ��U'�3>�-'���lW'\�D��~��
�0�5�����yw��� �̲���CTX���qDG�x���#'��s���$�h!KwMB�a)�]����.n$!h&�����B�}Ȑo�}���~�3�e�e?����\�Ԑ�*GI�B�'�������"�Q`�W{��I.YsD��j��9�p���V}��	�}m���#� �0��^B�T��������_�!e$�b"�U1J�˜3���#��ǈ�,
����̉q"Id7��mc	��}߬�:��"ȝ�Ͻ�Wn)OF2]���-�M։l�v��2[t��Y�w���m�vg��<�I��'$%/v�w��w��`�����;�~̘��3���;�9��^�]�˾�7���q��&=�+�w��h{���'ڗlF�S��U����ȇ����m!E"���ʅ��G���e���o�f�����Z'9��{8��I�g.o��u�Hl���b_5z��K;z�{�NT{��p^!��=���>�u5���x�|��q>R���6p%�~?��4p�Ó�@����ZC�:�}\�����V|�:B�"�v4���Pe�'z����J���(�VBu�n��>cB� ]��6Fk&ἆ��4,�ȱr��w�TN�HI�,XF�k|!L4�lBD,H�%4c�MMK��$��i������^�v.��8��q}99���_|��Μ3��+y�,��Ϭ98�&r'ٳ���w�8���޳���2p�ӭ9������X^<7���W�w���W�>�âG��[��9p�����	݅�0!�@��I�k����F�1��K0����3�NE��E1fpk���Mp�JK^��R�J`����!��g7��e���胭��v�~��Zf�!$����A7�N�[e"���'�9��׼zg�]�&���*�������W��$p��V0�Y�D�;췟tO�H����r�� /�c���ws=��S��MT!i���Ms3z����L�Nd�0�|�! �0)��I54���5���08�KVa-By�!bPI�2!J�9SG�|���}p����x����������C]��Ļs�O��8���>þ�#�A�%|��l��H�~���"V��ho�
"HG�����s�ː�4: I>ie��=>�[����z����Ufȸ4sKs����</�ϥƢ��gP��ʓS�`Ԝ0�"��q���E��bu0�[S>�u�f"}��B]�u��Ys��MU����B.}rq)�7���,��ɧ�_�Q�~,ľs��g���~�lቴ�2np泓�H[]F�(I��+d%l)_ѳ?o���h��GG>|��,��|�H]�0\"���/��}Ԭ2�|���4�T���u���������jT!W��	�&�N4�%g� BjT��r�g*M=��t��W���U3��A�����u�)�WW�����0arH�ܩu��b�&��T�}�y�rw������A>C��׃���$�g�8�}�Nyj�p=�G�S�ŪNg1}���gWG��"@�h�υcs��'c��_	���U4���:|���]�ӌ��#�����~�K����W�*��0şB���ᣟ��d�[Bt��d�B$X��4�Z��0��$�%y�?CI kW!?~�K1Dr�f|����_\�N�軝y9b��-��}y���i5j����q���/\�k������"V��Ω��B(�w�CN��;�Ēu)S��j��u�,lg(������^s��>[�}��3G��%�0�@$�F�B��<���b�~3�������ڮ����{�H�W˾uv*������ߔϗg�!�����QF��y��}��m��D�̧��A��
�|�D�ۍ�q;��*7���KRL�j*q��G/��]Ć�&���i	󘠓I��߽E���0ь?FjBYN���>��{����|�~�!6��b��%��->_O�w}��B����5J����S8��Vbjq�x��!?�P�Ó��%��_�#����bqQ���by=�`)z_�:��u���	�|��y���
㿘H$�?(O�O�=���~�JK��ß~�;���Թ�I	��ٳ!R0�a�$����=�|o��$���m \VEj���)j��g�.���"C@��u<��B���|�f��#9����Ј߰�%�T)�a�3���v�!����DԘS����>�#�9z���eth�}�[�xj�N8�{��. �ky��������:�d����<��i����17a�ލ��!-��Bu�y']��V=ۭ����.�\�R�n�4���Y*ۡ,^B�����JFƘ���`e3j��o���C�X�����y@��Rb�[�7[��e�ʑ��vC)���)	c������rl��ͺ��%&oy��!#��X��C���ݭ��7G'Ϋ��Y�ۉ,�����m���5�3�|���BK0O����B�S{*�qcJ'rW�r��_&O.����.�7�Νi�3ٟpU,���2����@��#�,Q8�#�Y�)50j�c���)�g&��ϵ~N�{1|�/'ܪ��9D�Ȑ�u0�FDthaB44"�aƟ�W�	,�H�O����޹?}�.Y�{{9�����j���xq��-�������_�Ԥ$����N$��{�ׂF����x���3�wZ�}��߳�;��
Á�A��f|��_�A�K�$���utj^.���&�Eg�%���(�鞥���:���=*8��8�9�ߎ��}�~���+�|}����|[�Dݚ{��ޤ>6@�O�	�>��5���X������4�I�q��(�oM5��/���Zgge�M�]sW�JŲ�.���8K9Y�M�}>G�����,'��!T$ ,՗���J�Q	��8����a�͛��z�>�'�J�Ǥh3��W8>^\z���Ǝ��߆<�os���5߾.p6P#_���%��#L����!�#�c]����i ���I�u�Ş1	�B��TYZ�<�%P{�]]�P�1b�����>�Z�};�bw;:y.)��E�9z��_\�|=n\���_q;�������#>�?r�,��S
��T�/uj��{����"K>��X��"���˿Es-�T��b&&�pycHQ����Ò�g:�C}��|�n+{�A���LM9��*H�-ou�B�\�Is=����Y1�\�a.C��ĩ��XL��v�u.�Kw��A:)UK2�� 函��K-��f���4�7;D	��O��`�����J���~&���\��տ]ݍ&�p�%[3l���q""}����^�
��=<�9�:��7���~�cϖ��z��Z��>���(��!�$8�4 ��5�Sܳ8H�+s�2�gq��(؜���8�~�=׉��8a[�2R˼n�\���q���0UV�gL��؏U�|�jI��5v1(�܄	���:1�1���HK� F?	��@�ũ�Fs���U</s��Ʈsy�"󳀅�p�=�YyX��1��hm^��FY�b{۫�;�������/�X���侬pO>߻s���W�u�k��s��Dz=�����9�pN��z����/��cO��w���%b��q��t�������� ����|�����\5�@��l�g�h?F��e�(*q�U̕�dW�k���^+_��G7е��{��I��L0��c���C4\y����dj{���Fp�W��px�F��̟r ����m������v�[���h���σ_��?�!��jk|3��g6F�2��j�a	L4`oY���>L&�亽�Xw��~;�ל(]�����BI O̤�a�����W*�$[=��z������>�����D��LNU�OR�ϵT���K�qO�U�q�fJ�����{��|�'���#�|��B.���,D|j�-]�]����.��U�>h�w�xOU^b��T)v9y�ﾚ�<&����['1���q{�hkȊ��38�IO��.�4s0Yx��E~�����4/r24�P��
UnDr���<��n�;,	��]�zg�\�~�]�>�yiw'��8y�M�1F���["8��Npi�r^;���0�9u%�ՙ2w�}�LFO�e���B��Y+,d	HL���V�Dթ�.��|=1�89���c٦B�-���Y�V%�8q��z.%�G��Y	q.FG%�Qn+r4Wy�Ͼj�g�	�`|a����=f�{u�������^	qwU3�|��	��$s�k�TŖ��&�	FH�XK!m%�#i.K�i�r�8#�t�8�m��S������D�Xt�qc��RZE��턲�!)KQ�O��13˶|�x��`���E��y-*n�E�{}����S�"�-�e�	1�ioé�VTG�>�;�;��;���j�q|����9�x2Mg۸���&�d�,(A�!H��2��PI��}�{��+s��a��߅8_���(C	aH��"��B�J.0��{��a,3'�˿|��z����w���yR��!lJ[s�L���d��|���X7����I���rpn �*Hߓ���������F��TGM��P��$#e���.XC ʵj�qf�KH���i>��<y9��E������9��I)YP���U �Z夳*y��#7�'��q9��:�!��
79߅2K������In�m����iܲݱf�N�l�P��)ae�w#���	���b���	�W����G�����+�,��F�1�\��â��x���.���D�(U�C�R�����������7(q�2B\�{/>���p��C��l\@���O�Й�FDA��Dݙ�� �mtmj}�->>���?��h��zZ��������!
FÇ�WO6��������F�l�mK'��Ϗ�}�/�y(���&�~�������s�̲�
B�-��,�4�BjK%6Ae�J���V�Խ����w�C����1�4 H�w�.k���t%�go��?�sD�h��7�]�������|��;]�B�Q8"@���!���i �$)���cY�r	T�R*XS���<�8s�%Dqt���c�a��_p$�m����į@��DLA�q����L��J���8\��;�w�:�Fy�d G�qT9S�*e��&,�)NF�����M��K�������y�g�}�l���Q�Ad J�B�u��6f�_6[�MfVX�\u�zSm>�<����{}��N��16�ؐ��KwR�e���˳V����I�2f���@�c�s�!���Ɉd���G/�3�Bq�`�SF��'�Ba�b�;��pi,ߞ*�%��+Vu!�s����aMF拠º&Wv�+��ğ��_q��Q-��r121��Ŭפ�[.��zbz�l�*6������B��Y\��J?�ߔ��"��s���g�s�g5�Gw�Nr#���\�����	�Å�TgҜ�a ��i}���X���������UUUUU)-UUU*�����UUUUUV���ꪪ��^P*���Z�����Z����Z��
�����*�����������������UUUUUUUUUUUU���UUUPUUUUUmR�UUUUQEUUUR��
�����c�UUZ�����������*UUUUUUUUUUUUYi��A�3�/L�,�����Wiwe�lgl�:�"���� ��r��98����uT�h.vZ���
��Hc��w.���C@���j,�@�j�g��䇶�;Z��ҵ]j��KѼ�� puԩ��mt�v��ڭ���,!���+��xȝ���f2� �F�:k�1�tSq�:\��="bV�т�u���Q�]����it\�ڝJPUWF��+"���y�2�!r��ګH�g���7��N����'d���6r�r�����Ö�*��Q����-�<P�̧	q���x׵ʹ[uV��gZ!!�-���)�*cS��8��$ݧv\��aݺ^��(���)#�康����#W��[��fl���j��v;��5����h)փ����q�c��(
͆�ZmEOk�qD�n�����h��yj��W��-ME`��L���6h��k�0�����p��mg�+u�嫪���
��� ���,7�c�8�=�n^�9w2�VR�x�x��IC\gQ�I����v��Zۖvn��.�[a㊱�K���M��]���(��6���6�x�+˻n7L�zI畕v۶j���BЗ ��[��U�Hv,���qƇ(ޗ�uPq��ۡ��(H�]U���ܷ=[=�*����Ee^�i�K�5��m۷X�n���u�`;<�Kh�k�d�x�ڶ)v�m��v�
�[K��۝F'�lPp���b�'��m�nכ�
�-S�漫��6�ţ\<���m5P��ĘZh8�q��UM�q�� �j�_`�6Ȯ���0:*�Q����U�L���d�`�Ӱ�E{9�J��;<�c1��D�/r�l�r�,k���VQ�cyR�D�*�:ٺ��ն^��&����VPmb@�2mMR�U@Fғ,'�M��4�Y[3���,e.�DL#�1�G��L���:a[���NiWYM��r���ԇ�f��H��R@�U�P�:���&�a��g�����U��	�tL�1s)Y:5�b��U	Dɥ�;8�gvK�z$�w3�]�IQȘf��K�Ksv��	K!P�����
�&Kx�1�e�n� Tr���k�u��Zd%�
�;C��[���喞��X������7����f0�0@�u�|��ޡ���lUUUC���3���;N��`n��{2a.�R�d��(U�vZ��+*�;���3۶;%vLO���WV�3<`���]�t�3���l�4���t��f:�𫲧n�W�q�k�&�u+�ʵZ=����h�ٝ��a���������L�UUm����J.4��ip
��Ғ����kU�ËGcnێ LgF�k5]
�<��H�dr�z�p�Ğ�h9{fj�����1�UUu�X�m�ڪ����!Ẫ���Q���]���O4M�%X��<�V^�)�&l�t+4��K�Y�������euG���y7e����{��;7:z�l�v��=k>���SOa��;*H�n��R��w�3�[��' g�S�3Q�-D�f��4X��jM�˞�$�6�ڲq]�;BbBݍ�F��]��A�rқ���T��h�g��j�s.7!��ŝ:�Wi;��Ț��<�p�U]�lm�!Ŝu[p����c{fᭂ�B.��n��y�wR�R%�ɋ��(;mY��i�9�h ��n(.��l;Te-�<sC��h
@�@*Ίq3l�����mhlr�M����ˠ�ն���:�<B��ò��^���2<�+���C�V�v�쑔խvb�E����z{�y5��@I�X�`��+�j�j��㎋��T�=Kmfb�]m�W ������f�k@�<�Pj3�����_e���麷s��S\�-J�<1��0���mX����N�nD9U�R4�ZǶF�v���u"k�J����A<����&qy�M�ܹ}�X�g)��%�н:ݷX(�p�T�מ(�7wd쑭�G���r"vZ���UK\�s� �FC���\��Td�K�ԪK�F�\���N�;��cc�Ӗ��XЀ��/�{oo�����Y@).��t���
��m]��n���m&������.� 
���2�$aڄ8�ɛR��Ra
9�l*�c��������N�&O/!qͱ����#kr�^��c����b7MT��iW��ɥT*��*�k7Z�Z-��')��{��=�;Ud+������U5N����d��F��XF0T���e�%֬GlnwcMt.z���]vY�����5A�(r��O9���.��u���^x�M�����,*�ť��A�%X�+���M���mUP�	X鞅�瓄#`����Ax���P�kg�M����jyХN�B�t�e�9�n���A)!��՚�I��X�N�mɞ�
�]����o��ٷdStj��8�U\�T��eۍ��q��iJm���n�d�ɖj��P�.�ڗ�L�c�KR�!���]��9d�����J��vٕe�R��%g. 㥬ĸ�C�3ۿ'W���7A^�1�IlcJȣ�5�X۶�)e�L=)vm�UE�{GP�@�uh����t��"6A�5T:��&yq*�֢��ƶٖ��lZLD�P��l��]���G]��MT���48�)V�xg��^�خ��;v5�؛K6�H���,n��
�����*s2�}:C��*�T V��Ճi��Z��vw(� G\`-�A�������km�&6�L�S�t�-ԫ��d������-����m� 6�h��ߊ��_��Tv�ꕔ�UWU[WUP�eY��l�b׶�]5�d�A+Ǌ+�ۂ	[�6:j�M�j��[g�s E]@n������vx8�j�Fـ-h[n*�X���	nƊv�V\�I�;%XK
l>Uoe�ؕ��f7Td���S��Lih+Se�VKr�(��ӴQUb�ƨ�5�Y%��a�
[/�+�E�Q�(�j��7K�vdCN�n���.S�\Ӎ\���A�+z��ڒ]A��T�:)V���v��+U��dy�j(8׍O*�� sR�Rp+A����W`�75&�+�7Uj�]�rT��fG��A�n��5��6��C��=��t�=T�vX��+l�Mٕ��õ֩��v���Ӹ�`!�u�m;)�)�\kM*�t�MP��f�X �vݕj(V�b�l���X▨3�ӝ����b�@^��x۪� ��o0�K�gc&�v������[-��j1�G��-E�.����ܸ�&�b%cU�Q�) ��;�]PNW���#'#ۜ.�2@��b�n6L���hSz��8u�\a�R^�7��]����*�%���,m�b \GW[f��������=UUe'�U�;�]��;�j�	]�T9
�F_U@v���W:8x;�5v������ by[��G�WZ̑$Ѹ��`��vXN��1�:���:�V�h;s,���ﾗ�9�/#&�	٥2S����s��@Z��.h\�=�
�yZ�Kn��N��9�2<��1ƙ��p��P��]���yZ��pj$�nݪ�Z���9
x�z�fUUT&��LXvԻ�;A^��9kiЯ1vYN�m(tbv�@u�jǎl8P�Y�].Y�a<�.�/i�%�y#Q&�p�FS������{�+S�^�v�r\�n �=�
̭�����H�%�o 'LX�,�:\�Y�v�V����.�fv��j�s����$���t�n�,]*�>�DN@���5���<7j�l+�R��UUU�����=���'c�ku�ŵZx�Y�Lde��:���#v���lڎ]��nH�q`��=�٣l����14�  ���F��M�4��E%�\7�
�⸶M����p�;�����i]K<�����	՝��^�L>��햝r1z1��!��Vԝ�D��6��
�V*�b�P�F�+��(MUUUU]R��ڮnոFCm��Q�sUc�����.g���I�KV��V��hk��ř���)��h7`ڔ6�ڮ���U�R�-T L�m%\k5�'����=2�*p6]��j�4���Ef�7a�5P��ح��U���W��V��
�����j����8��8j����3m6���51U��l��AA+-� P���@���-�P�����ibW�V������5������BZ\6˵�BU��UZ������	UZ���j�[�T
��;U]UUK�KUUWUTUPQ-R�U[��7P VԻ-uUR�u�[+�5mHPj�k����s
#�b�;d6@8��p�m/m2�rCWZ���r5R��+T���m�s�=[GkM��P���X�i)mt�׆�
�56��ɍ��UW//\��k����*����r�v�˝@j.V���Āgl�P&�:]��y2v�z�[��)���>&Cr+mZ�Ʒ!/nbv��EU	���Mp}�͜m�lՊ���V8r#�(㡠%Ml2���ںb����q��UUUU���^j���5 ��qc5�аQ -V�neZ����*���kn������Td^�ub�x�0EΠ^���o-@Wl�A~,_*��r����7����*�X*�����x´�e̻+��ծ�MI���X�-�[UUB��J�K����UUUTT�5�)j����
��W���U�*�P�v�V�M��7<N��uQ���m���j���ꪶ�j�4K��u4\���"(�z�y�"�'���@
	D6*`��,�ة���	���� ���D����H,,Ji�@B��ԋ��D� ڜ��� �Ҁ�@*�d�W�T�� ��uj"�64����AP���(q:� x���9���� �� HŁ�X��I ���Q�
Q�� BDA����R�!D��(����R)���т	�'H���(Db"#�WH�@���V��m�:�X$�`D"@@� � ��O��UN�u?+z)��0A��+I0 @����J�t��Q�<UO��
D�@�'Cb ���N5ht��T���8(���@O��BA�"i@N f�^����	"�h�ȧ~P�1����5�aE ����� �8�EC���Uڽ���O��X�H�� �ҨUG��(Ū~A!�_��(�W`��z�=@Jq��!$X�:��C�H΀ZB�����
+j`��U� 4��{���H� )�S`�Q�
=�
�)"�`��C8�AL@����(~T>0)�_�#�/U����Lһ� ��S�:*��4���I	$E�K
�XZFP��P�	Fe�l%ih���	#kKJB�Y$0ؒ��R0��0R�P��0�!!I��T>��Ͱ�		!��B	�$"�	#"�1��$>IPJ$Sl�$�!���XȌ���/�nB$�#$�""!�PC�hmM��?��mChP"�!�E? |���
���G�А"�B��h���H
�@8R�T�)sL���J 	 bE��T`T+Z%�K"���)++PcR�6\�$�C��^��M$��?�V*�j���_J�UP*�h
UU���X�UUP*��̘�n���m����<ґѷJ]3���%����U���rt���L���p�ܝ�Dݧ�i�1{��3���S�������eԛ�l��n^JC���R7�%ڒűsP���%, �Z��%�N-�ۮu�s���[.��
��LK]+/�X�vE�cĩ6�W�[Ԥe��E�-��M���D�I���s���v�m7]�.��WZD��u��-^e��'�J������a9����&d����=��Ƨ(��#���%��d9`�J�/cd�"��O9Bm�!���:��V��6+fįm4���!�`v2��ڻX7[�}���Vxڠ�q��C�{��t�3yL����Y�d�pt6+�c��	ul<��{MI��ڽ�!�;&,�_;-����J�
����/Y�g����t&�-�3�lL'����\�Z�*�na��Ѷ�m�3��<�9C]�&�-�H���F=��qõ��#\HN5���@�Ve(V�X�j1+e�R�-���8z�f���t�YF8��r�^x{nwn���Oj����݆.&8�ù�rY����V� �r��`v]A�s�v�Br��\�.����gN�S�FU��{kM�n��G���t�c�6������ݥ�sQ��[F����וte��.�j#�A2�u�m7ctj���n��3b�"��=���ɘs�u���i�Ų&6KZ7d�2�ϲ@h�ʖTU�Gl�m�[�ō&��t�E9�΂M[bղ�z=�]SF�+���� �F���V�ݶ.,��]F��c4��C�Fv�$�v��qe�bЌn��fD�F#���sh��N����[M�B(xu�-:�^7#(ר<���c���;������ò{�����cSdB퐦�f\w^� 5d]�;uP�&��q��p��[F	v��䴲�,��ۛ[�{,��b�Gf�l�nV�`��뻡�K�;�����Q�U4!��� �A��j(�Tz����D���(�Q��o�gufK���)JA��\Ge+5�vV.��:s������(8<ދ��������<<���#����mfsNK�2�9�`ؔ�9�.��t�n�v��LX�J�f�l$3(c��J%p�Kaf���X$���Z�v@�t���"y2(�۳v�:�X�]ø�{@t��#���r�RV��ژ�������a���\*\��'}���'{�p���l[�40��[��8�s�n�d���q����� ����")�� V���}�Izr�I$�9����{Ғ�:ҭ$�����ܮ��*�� ��}�_s����{Ԓ�:ҭ$�q�;Ԓ���*�a.: ?o<�w����^���;Ԓ��9V�K��+N�T*UEL���%�e2�$�q�;ԒY-��I��{������1T)vk��;gz�K%��I%��sޤ�!�*�A�����{����զ�uD��"s��q�k@�:#%S71.���.JL@�YY�˓+~ =�|�7�{���ۥ��n�|�g���J�Ⱁ�f6����}���8q#�&�N �H
X��������mo����m�nٍ����-��WH䨂����$d:eZI.�l�V�r&e9ߝ���߷}�~����mc\(ETU���v��bfRs�Si$���ޤ�c��_W����|JnW��j�o}��Ku6�K'1�z�FC�U���v�� ��C���hK�����lJ���S��3���9:�뱉�rY��am�F�t�t.֣3L�a%�w`��~��|��נ�v��$�Ku6�K��
�I!��*f��I,C�U���;gz�K%��I ���������������ڮ�F�͙��m��ߧ9m���u���S�(Q!	 �@ILB*���1@y�u��\���������Χ�9��K�V�����t ��I#"[���^yl�RIf'
&e�iMvz ?{��`����^yl�RId�Si$�1�:BS* au��ㄼs�\2��n9KMs,�2RdV���D�6��`7%�����o}�Iy峽I%��M��Y��I/L1��VX�W
�� ~��^���rI&ғ�ڛI$�7k�I#"[Ui$�ݦ����J�ﲅ�{�� �{��g�3)��Ҵ�Y�zw�%�Ԩ&�R����dz ߽�����t ~���9�o�g���@ۡ �A^����� ���-�o�
\5���-��I/y�;Ԓ2[Ui$���w�#��>�W��k�V�*ؕ�Θ�Vm���2�SVj�Pq1����WI��ObӇ��P�6�
=�y�_^� <����7[�#ޔ�q;�6�I�Ԕ�I�+�ɕ��|��= ��������f6��w4��oǵb�ITq7���U��^�uޤ��t�Z[ə��ӽ ���|�����Θ�,nW���9�ˍ��i$�6��RH�mU��?~�׾�?�wZ��:�P��@%�;gz�[N�Uu$��ݮ�$�:sS�m�tM�5�XP�E�A�/+$ǁ{���1t6�:傒�.�֩@m�Z�YM�!W����:um�ci��u��S���:�G.۞��`G=f��A[��N��L���Z �����{;�m��ۛu"�jg 0�o�c޾M.ݐ�Q�ݲFn8�fsr�aM��Z�8�kd��S`J3��:�8݋+{^X���#n�����vA���1��;R���7�X�Vn�@�Q�A'�ӻ�[��z`��Z���f#b�	�)[���]��%��O1����h�˴nP��������� ?~�׾��=3���i�ͷ�[\h�[��q։-��i{��{�92�ީ�I%���z�K'O@~�Il�z!Bl�8W��)瞓V�K�v��$�N:�I$���I,t=M6����k�=��9�w��$9z��I/y��RI,ƪ�$�s.C��et�2���/��G� ���^�I$���$��l����"9.66]�#���E�uiv9��0h�ٺ�{v�����n�;���u�+r<�J/�I$���P������[u��9����{�� }�~��:"��,C/}��~��Z߾
A��@��+t���	��8��P|���7���-�{=�� y�}�~=�㩠��չs�^��}������ <��^� <�^����]�av+vW�����Jt�U��M���$��j��I.���6ߵn8�9B���J�6�~���ԒK1��I$���z�FN5V�I��˿!�u��%�e4ystd�c@�ţ��,ٷ�a�� �/g331��� y�� ��}�_7��@��={��{v�,�P�L� �q��vfRr���I,ok�I!f55i��:���ysK�*�����t��ﻮr��b��
������.6�o���m�=�@�TH�)»� �瞽�P<�^��=������ ����������K1��I$���z�FN5`�u`wŷ{��4&���"C���)+�+2k6�#l��&��ٞ#��[d�i1t�sSST��;���y8Հw1Հ<ƪ���h��b�KQQ,� �Ok��X�j����de)PL�R*���`�u`1���:�N7�w|�e#���%�W%�������}�nI߳������l�A���P,E��H�����nIߏ�H��,�R�;]���p˜_��] ����5V���*&e�Ĺ��Ysme�\�-KQ�BV�^�K�Р]De�oMKjc��FT�%����x����c� �n��F95D�%)S*�Xf:��BA�Հy�Ձ��� ݏd�cn�Geb��p}��;�Հ�-� �c���T�(�*��e�ۀ{v�ٺ���� �/m�>�CaS��D[m���`�u`#Xq��=��[��#)B��!dP�y��[�aM�p��,I�lY���:m��u����uX���_����!v������6����GQ����v*"���r[.c��V��m��,�ٰB洰�@Ͷ���n��Q�m�Bf��#G6��56(L��)+.�cv��P]���9q�^�Km��c]�s����l�v���h)�m��LsZ�]9�C���1nZ�k4��a.
���l�=����g�[���z���V��a���˸eٗJ�&����<ݑO7m#q	�����&i`�~� y��;�Հ�;� ����NMA��k�� �/m��u`?Kj�=���n1���D�(�+cV� �۷ ��׀����{n���m�Uu��p춬َ��c���:����$uH�
������ �/m���p��xW�X��$�m�;t�b^:bR��D.�FBU��
�l�A��[�]�d%�n�F�[��z�� >���������ڰ=��;*�j`��SZ���krO������-H�8�h��`)���7f����}�p�~ۀ}�4F¦�%��*�l�mX|�XMc� �Ձ�W��k(�VZ��`����^:��X<s`g�!�e�IP���3U`bkX^X��k�̀w1��9���"�H���j*����dB
��-ƅ4ѥ]�A�P�iu�XE Pn�$QHIUW@<�Հכ� �c��_���n&۵�E`Y)� ��s{�y����a�K��_y�q ��$��Gq�[0���ׯ�p��I��R��o/2-��#���b_����T1<�`RM�ý�ۨ�ZP�&�Pk�����
��t��.S��o��أg9��G������/s2�Hܖ�k�Ζn��cq���g^�u�������aT�"D� �!��7�Ė��執��0�������]��H&!�S�hx��iM%�$��Tg.�,�Ss�̛�s���$��jܰp�޷~O��T��Ç>8����R��R���N�]k��$��"PJ�3��$�����(~���h����a��)	�@���q����9R�Dg%����|62�29?�#R��.h�t�s���$'��1�0
8˘L�d�٢IƤ�,ӶX��]���I�C�I7�\Ձk0��Lt�����ۦ����04�$!!0�,-������ٮR����3QZ��������VN�S��a$I;u9a FM�m�(HI!§�W��~�����*�T?<Q�+���>E�U�D`*�#�F� J��񨸟8�û��Ͼـo�d�l��)J�"���ɬu`�:��sa��$��{�շ���}�u�ȭȵ`�:��s`�:�<��V��(_��,x��m����R�^+z�e�:���Z���)�5ѻ�cjT1fYYUU]Vǹw����kls�@{Ձ�-�4E�2�+-Q�0��n��:��Xy���rj8����We��� ���������� ��ۀj��䖍;H�ݷ >����0��nY�	\H��� R�!4~v���ۯ�ܓ�w�-��+YdN�p}ݘW�.s���|�翮 }�J.���"�ElD���ܦ��q��Wjw.x:�k�p��Zڜ�YvT���RXH�
ㄶ`߽� ����}� ��ـo�d�]u؛v�P���ɬu`�:�1�5`�;�}��u�XJ�ۀ~O��נ=���;�u`4�:�:�J��-EEv��=� >����n }�m�>�mE��R��I^��XȈ������{V9Ƭ�(����s�8q�&n�`&K�kpe{��:�vv�"��M�]���͈��E��lۍ�j��e��)x�P.�LVg`�BR��k�[8�"��U�:��]Ie�*BrcQ6�5�n�	�=^}��-�V�5�sw�t-�K��]�mN�!{Ǡ˲�v�0&nn�����Rql#	�������ϓ�3�Fk	]�Q"��0r�xC<��嫝Sʸ|*�9�љ.�%nNf��g��a(�k�9XZ� ���ʜ��[����mmư|p�TQ��er[�~{�����_}� >���n�ǖ�8�HĕUX}����5cٰcڰ:��Vwۈ7/#VD� ��l����Լ�=� �=� �,I��I3�JTʚV���XZ�Հw���~�׀}�vH��e��mܷ ���Ձ���t�z�������"�!�k3a�	b�j������+����tx��M�rU���;�Vy=3����W���XӍXs}�G>�Hb�o�`y�����N;QQ\� ��k�$���Tr9��� }{VMnՀw����G�)�~�QE���+-D�����u5���ؙ=��`k��`6��R��H����S5Vȅ����ٻV��V�cڰ��)
�*���$$���;�����z������Ձ�I9=�}`�K��+�xL�7(41��%��a����cc
��������fβʚ䨩�U5^�;�{XMc��$�`w߿\������IT�V�ʺ�����q#�Sڰf�XӍ^�p/�z7�9�l���o�߷�VN_��nu�1�>"c��j! �H�$H�K��E:E�G"9ݎr8�r|Հ{wj��R�*�2�]�Ge��\O�߿LM����V�s��������T��TIMM��q�b9��,ǵ�<�=���ـq���'�?ҡ[V�KT΀m�F]Յn�偛�Ȗj�[f̈́],?����{���e����n����_��^nw���#�7%�=u.+���a�+����s���8���s�C�L�;��^�BC�7e!]ET%1D$$����ǳ`?N5f�9ďcڰ<�=�p������Tj������=V�{VSX��a��p9g9!�$H� ��؀'���ov`���U$C��$r� �Ձ��sө�t,{6��V܎s�����R&�"t�$R�4��.�0��mH�FR:ض����	��:Hf4<邦�� �5^�~�����~�����e�����m�����`�fE�������9Ȉ�>s���ߪ����^O�''6��~����\�ΰ7'uX������G��r9ɖ���l{��0觛QE��Ҳ�I^��qBY�j�̝����͇܈�9�"9ȉן������Py[���+����6l��Ds�s�̧���5�����V_�$���99 !=�]F:��@���m�5G�y��'sz^�ĺQ��k.��QT)i� b��:�Q	��
0���P�*b���d��e%(�F�-��gՖ�`�r�4k"�!��5��\Zv�޹[�[����a���볲�Di�vB�%�$/Yt�a��a\������ڜCe]��I�OC�V�j��\���2�5tob����kz�q��z��|�qy	�[xs.���sF��e �ȳ��6Ay	nƩv�b��b1ڶ貤��˓�o*�7ݒY��Lޜj�=�u���s�3'gf�͇Q�()1J�Ձm��=�?�Ŀ�IHk����n~�����s{H=�R�&jL
jT�ʪV,{6�.\ټ�G��ـo��x��I6�Kj��9l����9r#�M���l[��`g���s���{�۫o�v�`X�W0\X���s�򞮁��́�K�6���[�`�k�0P@�+K1�b-�[`�1lc��r$,,!�t���'F1�о�,P%5=�V�76�.\�DG:��w��?x[X��P�iYj$� ������v���,��Z���BҮ�ʬv�	��B��
H@ґ0+\�ް�+���3BQX� �E�4�6�`�X�M���$W �h'���5&��*�ݫ=8��"#�	�R�&���EvZW,�{��p�{n�ˋ�&u���[�M��1�	]M!LQ	T�R���s��/7���V��VI7�~�����"*b����-Xzq��s��r9��߫������ŀ|��B{���؈Ԯ�Q(J�,^�6���5J�B79�A5V˓^>䜄0�M�
�ԩ�&�zО����[Vq���qs����� ����$V�9%�rT��ӫ��r9�L���Ł���`uf=�ܒp/�O��XA�+��^����nI���sso���C�L�`�F��R�	P�I%�2 B 1C��v�s7$��ݿ�ܓ�N��&�F��*j���ĸ�{L�w��y�V��9��b��!�"cjEQH��SS`uf9�7��DB�յ�<���<���^�ޡ�������W��:�klMSD�5�^m����҆@�}'9'�c�2*�h��J� {ߟ�}�w/c��"#��&�l�艙��#���K]�������9���~�� �of�=�^�9����`�*
i��k5�rN߻�ܓ�ﻛ��� ����� ����X �7ڤ�;�[J������Y-��f����Ł��+�
�!_���� @��BHI!6NJ�b�� ��|�
�f����'���z¸�K��A޶߯��������ӻ������j{��O�����$��On��jb�[����D��F�m9ͭ(3�r��izwN�;��L��G/@�ݸ�1{�Y�v#��GP��XM~��2B��%� >���Ģ"17�`�ڰ;��^�9č�6�#�D)]e��n��`z{n�r"�ݸ�cڰ;�jHW0J��H��a�#��Dr"e�~�7�,��VG#�����DK�ߦ�ߠ߄
mRRJV�)m�>��,���$���������{�ٴ�Kı/�N�[ND�,K!���`|�$�B�����!,�"B����gT�%%R�"XFR�Bb�j!u-��o3�2_,�t.4
ц�01���B��$H�Cc.&?k�Ѱ%(�΄�������:L\M��hl`n�5
� @�@FF0`B�T� [��	h$#���;"�)�}Є�CDbD�A�I�\uS��:���&@��f8a����M:�+��"�Q���d۹�T����R�ޝk��*�a͙Ðtq��ߍ�6�X3����Y�㉵��:딸��$���I�Ѝƍ��GZ��>��lMbD��&�0Vd]����W�����*���h���P*�h
�����4��UUUU�@T�.�FBru��F���}�lt�nr���4�|㋆L�m�J����B=E�r�����l�tk����7<�cq��U��&�/���)�&�1�	r�<x��ՔɖM�����K*�@V�wkv6�۷l���A�\WM�v��,�7c�����:�w����K��%P�و��h����c��Ksd+� ���Fۘ�V,�l��q�%��-�4��ҷa�����b:d����
6	��ix˻nQ��j��6���cq�M���{rZ�G�g�7�F���y+��8�W/.�Con1l�k����@g��(p�7���9y��k�lh�l�>0�z"9G��$"���s`9�˫�س�Ϸ�u)뀃�=C�;0fHD�&�ir:��]���J�XYL5M�#k���&$���fx���x.�.�s�X�KfC㑷h[���n�v��×�:	��s�&9�n:ks`�l'm� ��ϱe��s:����uJn��	�^.1qZ�u���nz�6�m�]=[e�y�����[�:�� Vܢǝ8�X8`��#m���8����]��Ya����S�l � ���a��)m��M�	��_gF��ي�2�f��m�\�� �i�["ɶpZ�l�ӝV�Y��r:;���8��bU��n���fM<��O��:(�@h�kaUȒ��T�{O)m�N���ێ�`T���um���`��9{h�;X��z2gZ�e�Vf���T�mm�e���m�b�GՕ "iyv�y�x�;m�I����0)��֣ф��qWa��`1��v��;]+�.�c/:ݜf�[�ݝTy���U��;��	y�B�V[E���;, ���Om�N�.��j-:Z���)r�r`Ý�g$��V��O`k��v�ج.CZ9��@�c<k��8$���&v�P���CAU۝Y�J�,hCP��m2K�F��ϚC7G��Mf��ֳFfk0�:m��U�*�x*� a�
*��"�DCJ��E\6 (��"��b!�Es��y,����a�gƝKM��:�d�jK`��f#f�fxN��I<���f��i�3Ɣ�쫼�p���Ƀ9�����IS�=����!�v��sŻt�M��Lݸ��bذ�lB��ì�Y��N�K�;�s6\���9���/��<mr{?[N�Nl��<�U�r�i���D�a+a�f�L�i+�+I�TQ�>k�u��Z�1�A��x��.CjP1���rǢC[,e����:#nv�%�ܰ�"���t����'W��������t�ı,K������Kı>���Kı/�N�[@�,K���{��'w����/!?_��]�m!�g5��"X�%��u�]�!� AAșĽ������bX�'�����Kı/��m9Vı,O���s&��W�����8���'����,K���{�ӑ,�`*�L�{�kiȖ%�bw����r%�bX��}Ѿ�a2�r�U듻�^B��}�ND�,K��}��"X�%��{�M�"X�
��~�{��r%�bX�zO,�e�I�$�h�r%�bX�������bX� 	�{�M�"X�%�~�w��r%�bX���p�'w����/!��>�"Z+��!6�gs�Ng';1��x��Um�hZmWe�2�ޝ���Ժ{�0,Z�g�/Mzk�T��ߦӑ,KĿ};�m9ı,O���l?����&D�,K�}���'Mzk�^����]�\Ԇ�Pw�|�bX�%����Ӑ�����!
�AJA�@�H� a-�,����H�$��1"ń"$
@H����]�,�Ȗ&��p�r%�bX��{��r%�bX�w]��r
��bX��;�Is��2�[u0ֵ��"X�%�����"X�%�}�kiȖ(	bX�w���r%�bX����[ND�,K�{�Il�nfh�Z�ִm9ıT����ӑ,K�����iȖ%�b_���m9İ?�"dO�����r%�b[�O����Pf	��Y�}���MzX�}��m9ı,T�w��r%�bX����m9ı,K��{[ND������y-��/650k�@��e�E�]M41����K�0�qG5nm���'t����v�qL���N�!y�^C��}��"X�%�����"X�%�}�ka�"�Q�L�bX����6��צ�5�������i�[Q��O�,K���{�ӑPı,K��{[ND�,K���6��bX�'�>ﵴ�O�`�DȖ'L?��2���sRf�3Z6��bX�%�����Kı>�}�iȖ5 �Ey�\*�� dL�ܚ絴�Kı>��iȖ%�bw��/�h̆�5f��ӑ,K?�`��N��ߍ�"X�%�ܝ���ӑ,K���{�ӑ,K! ���{I���t��K�܈��I$r�\@�������� ���ٴ�Kı>���ӑ,K�����"X�%���&e��'�r�6��V�Yc�ҷ�4�X�Kp�x�]lޝ:ve���=v!��MU}ӑ,K���{�ӑ,K����ͧ"X�%�~�}���"X�%��O��_L�g8��7?N�q���M�"X�%���{�NDT,KĿw��ӑ,K��'�����bX�'���6���X�%�N��34\����֮�Z�r%�bX�����r%�bX�d���ӑ,Bı?w���Kı?}�siȖ%�b~���j�]ff�IsL�f�iȖ%���Aȝ;�]�"X�%�����m9ı,O�{��r%�`t����--H�P'Sr�^�b/ ���AdK�����r%�bX����ˬ��JSF��h��k6��bX�'���6��bX��(AQ�^��m?D�,K����ӑ,K���w=�ND�,K����H�,cH�
��`��0[;���[�e�x7�a;]#���M�}o���k���f�m9ı,O���6��bX�%������bX�'�k���Ȗ%�b~��iȖ%�b{�қ�٢�kSVf��iȖ%�b_��ki�(���,N�^���r%�bX�{���ӑ,K����iȭ�bX�=�z�B9�T_t�zk�^������Ȗ%�b~��iȖ%��;�fӑ,KĿw��ӑ,K���߮���mF�L�u���/!d�/'���6��bX�'��}�ND�,K��}�ND�,��{���Kĳ�߹�_ZB0��D���N�!y�T���iȖ%�a������i�%�bX����ӑ,K���{�ӑ,K��ԀH� ���3,l͟��d#]�*.�ǯ1��.!�b��L۸���y����0���d�˲�����:��5n�Mm�3e�#`֘��XiL0�,�m����O�i.eM�{�9vN�c��GU�v�p[A;<�I7�G���Y��=�sz�ꐊ�ϗ��	%n�6,��R�P��FްM��Дf�� n��v��e�Aŵ�lc�l�4�t���N���23��6g��Ŏ�97:P'���]���9J�l���s�b'Z�J�hW3�t�o��q����ͧ"X�%�}���m9ı,N����ND�,K�}��DȖ%��=�fӑ,K�����պ�f]\�晚�fӑ,K��{���Kı?w���Kı?g���r%�bX�g{��r X�%��{y}��JSI�����r%�bX���p�r%�bX��wٴ�K,K��}�ND�,K���fӑ,K��$<x�o���Y�,�h�r%�b%���}�ND�,K��}�ND�,K����iȖ%�'���6��bX�'s��"q�c!]d��3�㉜L�g���Ȗ%�a���?��?D�,K�p�r%�bX�g���r%�b3��7��r2Q��d�*ܳ�Cq��j3���
Υ)�����ֶ��wOC�ޥЎA��'�}^��צ�?}�ot�x�,K�}�ND�,K��}��Kı>���Kı:x��K���4Q:����������w:��h^�����T��C�K��s�ͧ"X�%��k޻ND�,K���ӑ?�T�"X������ҽFQ΢��>^��צ�>�����r%�bX�w]��r%���bw����r%�bX���p�r%�bX���}�V-Ĺ�s�������9,O����9ı,N����ND�,K�}�ND�,��9�{�6��צ�5����w��e 7[����O��ı;����9ı,O���m9ı,O���6��bX�'��}v����/!y=��}�G2GLd�dA�Ms̀��
���<��sK5bU�k����Ͻ�H�4#kGQ��O���5�O���6��bX�'��}�ND�,K�u�]���bX�'{��]�"X�%��Hx����VY�h�r%�bX����m9�"X�g���ND�,K�����r%�bX���p�rI�L�g�lR)�+��9fq}ı,O���6��bX�'{��]�"X�܏"�q`62��V0b�c2B) �  C�� P؇��?w���Kı=�w��'w����/'�߹���֣����m9İ@�;����9ı,O���m9ı,O���6��bX��\��{�ٴ�Kı=�'����n\�u��f�uv��bX�'���6��bX�+�=�fӑ,K��;�fӑ,K������r%�bX���^��~�FSh�-s�.���y�Xm>��
bp�f60I��fb�l�ڲ�Q֎'�%�b}���ͧ"X�%��u�]�"X�%�߻��yı,O���s�N�!y�^B~���6b��k5�ND�,K�u�]� �%�bw��z�9ı,O��m9ı,O���6����1L��,O�O���[�au�$��kY���Kı=�n]�"X�%�����"X�bX����m9ı,O���6��bX�'���S���Ɇ�\��B�I���~�m9ı,O���6��bX�'��~�ND�,��)��dM��O]�"X�%�ܐ��%���5sF[�Ѵ�Kı?g���r%�bX����m9ı,N���]�"X�%�����"X�%���9��e&s)��:kG!Z4�eE`qɚ9���q��j[gm�hE���ޡl��΢a=�ꥉbX�����"X�%���w�iȖ%�b}�{���Kı?g���|�5�Mz~O����)BU2�3�9ı,N���6��ؖ%��}�ND�,K�{�ͧ"X�%��{�ND�T��2%�����Y��W.e��u�kZ�ND�,K�p�r%�bX����m9��`Dȝ���m9ı,N�{�iȖ%�bw݆�2�70���>^���I���?O'"X�%��}�ND�,K����iȖ%�b}�{�ӑ,Kħ�[��eM���+��'w����/'���fӑ,K�O�;�M�"X�%��}�ND�,K�{�ͧ"X�%��O����mu��)imy�]�dK`ͩ����Y�� ����*��v�:"�v$܄�QM����[K).a�hd���=���V�`ǎϠ���u�u�R暰�{t��87j�X3��n	`kkF���&��) c�� b�݂�e)G�����<�v1.�_�&v⦍��'��C��f0��۪�tIne��2z�Kt�#����I�
�&�s�����N�}����!V{V�<qP �<J�Hm���4(�J;�r�ʵ�4�w䜷��U��n2�4m9ı,N�=���Kı;�{�ӑ,K�����`��bX�'���m9ı,O{�����4jML�fkSiȖ%�bw���"�bX����m9ı,O���m9ı,O�;�M�"�	�2%����o�X�m�{���^��ק����{�D�,K��޻ND�Fı>���6��bX�'���m9ı,O����
:���a=���Mgtק���]�"X�%��gw��Kı>��iȖ%��
�������i��zk�^��������@L���O��ı>���6��bX��w���Kı?g���r%�bX�w^��;���/!y>�_���v�f�0Χ���ؖv���z����t$��+t]��+i뮄�cj7Uo\��B����{��m9ı,O��{6��bX�'�׽v��%�bX�vw~�ND�,K����sQ4�\�듻�^B�?g���r?u�^�J	!QM��ҬiSPL�����@��0!)JȲ2I b[C�`�c�|��؀��&D�7���m9ı,O����M�"X�%��}�NEı,K����f�5�k5n�Z�Y��r%�bX�g}��r%�bX�vw~�ND��b�Dȝ����"X�%��fӑ,Kľ��}��5��,2��N�!y�^O=�ߦӑ,K�����"X�%��=�fӑ,KlO���m9ı,g�?|^mk[�̷�N�!y�T����"X�%�����m9ı,O���m9ı,N���6��bX�q{MC<��'?UJ�M�Hӑ�X��Dc�Cj�$�3+�H:Xmr]7��z{Y�]e֦��Ѵ�Kı?g���r%�bX�g}��r%�bX����lD�,K���6��bX�'��}�S2�2j��]f�iȖ%�b}���iȖ%�bw�w��Kı>�}�iȖ%�b~�{ٴ�O�dL�bx���� [�ʪ����צ�5���?}�6��bX�'��m9������d����) ��@�B%�������80tG���A��-3_�-I�V~�d�%6F�d=2f�40�4J%�Ӝ�X�?���kan0 r ^%>�}����,J!e�,.}h�K	͘HC�	 �ն$-l�^3	Ҕ��J3����4ȕ��b�A(��q`��P3Nc!��aD��fkR�$����Ԙ섄�)�B$�l.a�G��,K�P�[dt�-�B:��)
C�B��'�~��F�m�0ǐ�		�j�1e���seT#G|�d,����˕RXC���l%���p��1�'xϑ���� ������C����!L����il���4���	4�!n�i�a������²0�R�iN8�~"��4
���f*��:"�|�����E��TM���Uꃂ��j��� ."s7߳iȖ%�b{=�fӑ,K���w��jk.fL�˩MkSiȖ%�X�w���Kı?g���r%�bX����m9ı,N���6��bX�'|z{�Zk	�n�jMfkFӑ,K�����iȖ%�`���m9ı,N���6��g���;�p�r%�bX��ϻ��{����s�g6��!��Y)�.<���Ɏ�S��0#�ݝ'��Lܵ��6�Y��ı,O���ٴ�Kı;ӻ��r%�bX�w���@��dK��?���iȖ%�b_�����5�!5��.kZͧ"X�%�ޝߦӑ,K�����"X�%��=�fӑ,K��;�fӑ,K����[��!lѩ2f�3Z�ND�,K���6��bX�'�k޻ND��dL�����m9ı,N�{�iȖ%�b~1��%�u�����[�6��bX�'�k޻ND�,K�｛ND�,K�;�M�"X��,!	R)$Q���|6��bX�'��}����dWd듻�^B�����n�;�bX�/zw~�ND�,K�w~�ND�,K�k޻ND�,K��w�����Z0���$ڱ (�W@e͍E�9��9�e�.��Ҷ���z� S.��ֵ�O�,K�����M�"X�%����M�"X�%���]�Ȗ%�bw>��iȖ%�b~��_Kxj�tf�]JkZ�ND�,K�w~�ND�,K�k޻ND�,K����ND�,K�;�M�"%�bwϽ��5�&��5��M�"X�%��=�fӑ,K��{�ͧ"X��bw�w��Kı;���iȖ%�b~�S�35�u0�e�Z���fӑ,K?�b�����m9ı,Ox���ӑ,K�﻿M�"X�%��=�fӑ,Kľ���b�:W�˺����������_]�"X�%�� D}��M��%�b}���ٴ�Kı;��iȖ%��/�ū�BI|���j� �����m�+N��;S���c�-,^����a*L�csT�������5YT,�5��	l�]R��#tWTM,�n�C4�mɢTSK
���\q۝�s�X�Rhu�L��ʗD�h��-��bS۵��5�nGN�v�=c��-)��=;f���xۼ]��j��ٹn�+sd����H��3��ys����m^�ǂ��Q��5N�(mD�� �533
a.)�o���,KK�5�g���Nl�k���gk8����\̄��6EB�KL���bX�'���m9ı,O��{6��bX�'��{6��bX�'zw~�NF�������O����-pfu��Kı?g���r%�b}���iȖ%�bw����r%�bX�w��N�''�^B�{��Φ��R���fӑ,K�����"X�%�߻7��K�
9"w���6��bX�'�����ND�,K�}�^ffL�����ffh�r%�bX����6��bX�'���m9ı,O���6��bX ؟w���Kı>��_Kxj�tf�]JkZ�ND�,K���6��bX�(����m9ı,O��p�r%�bX����m9ı,O�<�u`�X��YJ�����4e8���u�v�4dG"�FX'�F�M(�6���r%�bX���z�9ı,O��p�r%�bX����l@9ı,O�w��\��B�����o�M���*�sWiȖ%�b~����(�/�[@�x}�4b�Q?(�%�bw��~�ND�,K�}�ND�,K���]�"X�%�}�K3�Z��Ri����"X�%���o�iȖ%�b~����K,K���]�"X�%�����ND�,K������\55Lՙ5���K�V���}��A?{;�$D�ﻤ�D}��ߦӑ,K���<d��SV�kSW34m9ı,O��}v��bX�'��m9ı,N��~�ND�,K����"X�%�}��<j�SW5O�5���ظ�fc�ndRR1l�B]�.J��F[��jk�Og�� 
��A���zk�^�'���6��bX�'zw~�ND�,K�����%�bX���z�9ı������o�ˁ�`}���MzX�vw~�ND�,K�{�ND�,K���]�"X�%����6���%������S�;��0�V����/%�b~�}�iȖ%�b~����K q4�#��`p ș��8m9ı,O};�ND�,K�>ߥ�W
e�3RL�h�r%�bX�{^��r%�bX�}�p�r%�bX�w��6��bX�b~����'w����/'�7ߦ��,v
���ND�,K���6��bX�
����"X�%�����"X�%��k޻ND�,K}����)&fT���^-G<�e�,s���lSӛ3l`������۵ژD)�h���;��y�^B'~���"X�%�����"X�%��k޻���ı;�p�|�5�Mz���%��5�u�g��,K���{�ӐQ,K���]�"X�%��{��~��,K����6��bX�'�!�_�?�e��]jjۚ6��bX�'}���9ı,O��p�r%��bX��xm9ı,O��m9ı,O��{Y���VjjMdֳ5v��bX�b~�}�iȖ%�bw����Kı?w���K��~��bf���ܻND�,K��ﬧx.ٮ�fu���/!yý��"X�%�?��p�r%�bX�{]��r%�bX���p�r%�b3����@p	"�����5j�!�m�r��)Xͩ\�)b9��	hXu9:өN��.їR�f��"X�%�����"X�%����ӑ,K�������@I�&D�,O{���ӑ,K������vF�T�Kj�/�&q3��]�w��r�D2&D�>���m9ı,O{���ӑ,K��{�ND����^����o��Hƚ8ڮ\;�9ı,O����m9ı,N��m9ı,N��p�r%�bX���z�9ı,O���s�u0��4Y�6��bY�9�;��ӑ,K��{�ND�,K�{�ͧ"X��C"w��ߍ�"X�%����{�ɬm�M\ՙ3Fӑ,K�����"X�%��$~����i�%�bX�����"X�%��{}�iȖ%�b~4M�@�N�مJR Oɘ��������@���\2�9�2�=b^˦uls��4p��لq��LB3�X��t��ݑI��@�i[	cR�,���m�D�aB�[��Lkѹl��o[N�iL�)�R���zr�����t�m�c�7�7	5���{h&��2���6Z�t+ۗ�`Î^���p���
���fe��{;K��\;���;�ՠ�XG:,�ŮM���S������O�':i	���|�t���`��U�R�Rф��kK��434f���bࡆ#Fc6k�t���`0�Z�����Kı;�fӑ,K�����"X�%��{}�iȖ%�bw�{�ӑ,K���]d�,ՙ5&�j�5�ND�,K�w�6����ș����6��bX�'����iȖ%�b}��iȖ%�bx�}	y��5������Ѵ�Kı>�o�m9ı,N��p�r%�bX����m9ı,O��p�r%�bX�<v�R�-�Z2��\Ѵ�K��;���iȖ%�b~�wٴ�Kı>����r%�`+"w��ߍ�"X�%����Œ�$�h��.kFӑ,K�����iȖ%�b}�w��Kı>��m9ı,O�{�6��bX�'㿾���,"F��ʓrC[�ڂÅ��y3�M�0��p6��mP�ԕ��==�%�.[���m9ı,O���6��bX�'ݝ��"X�%���{���F?�dK��?���iȖ%�b}����k&����[��ND�,K����Ӑ�䊌�x@�'�"X�'��p�r%�bX�g���r%�bX�}�p�rbX�'��{�&��L55sE��6��bX�'��ND�,K�{�ͧ"X�
C"dN�{��ӑ,KĽ������bX�'���g���Y�MKsFӑ,K�?g���r%�bX�{���Kı/������bX��߽�ND�,K��g��.Y4jjMd��k6��bX�'��m9ı,?�#�z�~6��X�%�����ӑ,K����iȖ%�bw�<�%1H�0�Y�k	b����hZѡ�R&��F&�[ilތ��6�!��j 3�r%�bX�w��ND�,K�w�6��bX�'��}v��bX�'�w�7���/!y����}I�r����;&ӑ,K�����"X�%����]�"X�%�����"X�%��{���[ı;�G|Yn�5��L�kFӑ,K����ӑ,K���{�ӑ,��@��))�R ��� �$ pN, �br'�����Kı?����iȖ%�b}�N�ylqr�ý���M�Y8�>����ND�,K���p�r%�bX��}�iȖ%��L��{�6��bX�'���_�d�·0�k.�6��bX�'�ﳆӑ,K�{���Kı>�wٴ�Kı=�o�iȖ%�^O|��|^�f��-30���;t��l��@=��zӍ��+X�'����z�:�CSWZ�.h�r%�bX����iȖ%�b~�wٴ�Kı=�o�iȖ%�b}��p�r%�bX�d�ǲ�2�f�533Fӑ,K�����i� r&D�?����6��bX�'}?��m9ı,O{���Kı?{]�MD�mڣ��'w����/'�}��iȖ%�b}�_p�r%��	r&D�����"X�%�����ͧ"X�0���>���i�[�\޹;���,A�>ﯸm9ı,N����Kı;���iȖ%��0v5J;h�W�V�XD ��'���D浾M�"X�%��I��r�Re�k���h�r%�bX����iȖ%�a�E=�����~�bX�'����6��bX�'����ӑ,K��'C����A�̶�`�pS`c*�+�����'�܀p�z�tɆ�rz��	ܓ�fu�iȖ%�bw=�fӑ,K����M�"X�%��}���,K��}�ND�,K�t��F����u����m9ı,Ow���r"X�%��}���Kı=�{�ӑ,K��{�ͧ"!�2%��=��]jh�9�u�Z�ND�,K����ND�,K���m9���{�ͧ"X�%���~�ND�,K��=��3$���-֍�"X�(@ȟ����m9ı,O���ٴ�Kı=�o�iȖ%��'���ND�,K���3�CY�֦�fh�r%�bX��{ٴ�Kı=�o�iȖ%�b{����Kı=�{�ӑ,K�����WM�;��n��k��,�H�����މ���{��k�l&)�1xh�CL�֟�H/���p�~$���1c�6�>(d���!~�@�D$�E�	$ ��0$�F)���H�2B��ws��tZ��J�w~p������,ިL�L������~Ù��Č\B�^ዯ�|����h[l+��
����b�� �� *�T�l�[UU[UUS��<�jՋ��F{U��LF�ᐞ�l*X����l�3�&@�㣄�9����\l���1�F�� ��l8�-�eP���F�F�*u]ZY8Ꭸ�uRŚu���[��e3eR���[�M %#I�f��6���8A
��'EF8�x6
�w{'"k�mi%s���`���Y:x�{q뛰���N��D3��p)��k��x7�,����h��ER�ե+Z���ذm�v�<�q��)W�mi6kKj:n�iط �F���i$83�aFM�jL5�f��ۉ,0�0"l!ZE�uv�r�[�n5� 3kvϭ�������A��9u����ր�t��������y���N�f���t*Ѧ5
���°1a�ci�������g�'�5c]��<���֖��K�vqc��mת�0�Uܣi�!!�s��3���I���A�s�d����	��������<v�;R6�1��S�=��c��=d��cU��Ų�=!��re�c�;q`1�8��:M���<;v��륉�N��ĭrC��N��g�:�ɼ��^Õ��D�ՖY6kVX��3f�	��G[rsV�|#qFg�k ׳�}�q�]\�e�8���g���WYXЎ�B�X�X��{5��>�m�佋G\\-�ϓXIҙv��V�.y�����0��v�s�9{�x�*W���m�8��,���,XKw	b3\�ܖ7�^���@�^Gۨ(�8�2I�s�6�v���8z���P�ۅ��3,��Ҷ��ꕯ\���nrX�1.Y����8].:�7a��s�6��;�%���\�`��/4��J�R(�i6�듫�oZ�^�=���.����b%9w
�ۛ[�����2nDb��v
C"��]ͮv`�N�Փhx֦�v�y3v۲��n�)����:�mXt-pu��m`�jh����� �V�I���V�ӹ�\pm�E��T���xrh�FY�`�#����$�pQJ��
u�K����h���@
!���]����)�N���� j�� ���G@P�⢟}�j�Ÿ��d��<mZ��6mr	5���W�tn���5`<��:m�jR��f��q6:�4�����c��:�͈ƌ{H�4�ꅶU*C�G�{/Ec\�r�ÜA�5\��g�Gm��F��]�ڦvK�@	�cF�X�*L��f���@җApR��M���W5⒓�C.g�Q���,�Be"[),t��p3P��k`@�+�0�4t��'�wKӤ{��o	�\����;��#h�p���U�b�f3r]b�M�斮��:lz��ƕ�m
�f�i�%�bX�w���r%�bX�笠m9ı,O{���Q �dK�������r%�bX����y��J�%-�9L���g8���7��8��bX�'��p�r%�bX����m9ı,O{���r'�0ș����~�\|+!��3�>^��צ������iȖ%�b_}�kiȖ%�b{�ߦӑ,K��Ӿ��Kķ���?_�Py�u�ȳ�N�!y$��{[ND�,K�׽v��bX�'ޝ��"X�'}�p�r%�L�}�F�R^Z�%�Y����y��,yL��s`{�`8,���f�E���ճ-�u�T�q֓��4]�=�m��l�LD����z��c3`�������[q`<�e�ױ���9��Y�6�?�i�@vW8�j�7޺g�q$$B@�	����	�DW"�">�G<�Orlr�X�����|�{�7��\���`}ݘ�n�7���׷�ZX�ƨ&$����*����[9�6F���e2���!9�ٰ67M���QS4MQ*j�C�q`ls������`�Ձ���"{�*����2�0�M6 E����5���W��nn�;Li��V�*��8���S,�w ��}��9�G#�>߮,����@�qJ�*��Uy���"9�<ݫ#^�XyL��#�����*�[���-X����[��r�m�C�`1T&��u��wۋ �צ�+U:)j���p?q$�5�b��u���n����$��Xg�J�e�vW8�j�=��`���w���j��y���@�ffe%$�c]M6�8GPLAB�Y�lf��� �^I�;r�����V
K�\�Ucv�{� c�Vc��lG#����n^�	� �(�d����1����Dɐ����߿_� �}t��6o�����F씖�J�ћ�<�Y�9ĳi`^Ձ���<v��Ecv+%Xˋ�q���,�ZX<ua���q� Q<9�F�##.1��b}@�Gj|(���O�?�o���w�~?�+�;X��`ﮘ�����,<�XDz1�bTL�T�)�O��,br4)W)��4Q`��bÞ�k�gI��c��tf�V5�nh�-��߽��;n���e2����`5��54�O�ER��p�wqg���I)������7��`�j��&i��SSJy	UE��S,y��>��$n��#7�,���Nj��e
۔�;��X �:�=n��b"�,��L"ӕHJ�X��Wwq`��`��,9Ϲ��݄V�T:КA��L��:]j��]h��KB0GA�1��Z�"�v�Ή8��v�j(��{ m��\:�q����e���6sv���9�'Qp�7k�l�^�)�1^p�a-\j��G���;4� ��h���D[��83�Pj!P���AXp���ۚ+�[ZD�bָ6y���6�NȣF�s%��y��k�pnpع�gB4�_�@_ M~��Ԓj���5Ln�-�I�$z��n��Q�W�Cvʦv�s�1[!`�"�7%�W��,�륁���r9r= |����߀��&�	R����e2��Ff�ŀn�Ձ���Y��;�~���'J�,����q`�V>q,�u7L��2y<��T����,mՁ���7L�;��X��6�b���C��n��w��:f�ŀcn��`����� 1=�<�/6�t-ֳZe�]�ڮ�n\����k&K�ȸ��rέ�{��`w��X6��s�H8{�Ł����#3�����-���'?w�6��`�"��`AM�(��}�w[�~�}ݬ��qs�����b'!]|�B�j��j���w<�X�;��зR�Y��-���s�����`��K��q`�Հ��I\T��J�D�E��)�����1��ŀ}�k�Q��ۍ6E2�6V�L�u"�薄-&L�F������7�m���[i�w��X�����Xﮘڶ�ET�ʤ��W*��m��r=��q`j׳`{��/RŤ�IJ��9-�����, ���>��EI�Aia���`E$�B!	@`@�b����'M_���ܒw����v�X�VI,�$�j�o����c�V0��X�*u���Jj�{ŀ<�V�7q`�Հw���ƚ�J��Z�|�r��_bsВM�"�G�[p�]�*Q��B�Z��T���ɒiUG@3^Ձ��Xy��=�w�X�ȥr�$r[�w��,���y�Vcۋ ��V`cIR�q�G]$� =�ۀw��X����7q`�=�)t%Q�m�;�n, ��nޛ��>��!$��E��T��u���nI��tt��C�GIl�U��m�?q%�/~���}���;��X�P�^RLr�� �d����9���:mn�i�fV����VT��h�n(.�)S㲇$�����������ŀ{v�z�\��W$����TXf:�=��,^nlG����D6~O�Z���m�J;-�=�߱`�ݸWwq`~��ޞ����I&�TX[u`{�w,�6�B�?�,ߵ��J�d��nޞ�V�C��z��ŀu�V�s�www�箲�՛b�	S"ԙ)@u�C����+78����AZ\u��+��ls�[E/^�0��dK٭՚�uy�4we(�k(�.I�Cc�����Ќa%R�]�]�K�[0b�m���Nv�+�b���g·0Ҽ'#Q�j�x�����Ҕm̢K����.��:�J�ؠ�(U���-�v+�ef+����ve�h�ˌ͡"�i��:O��i�?9�s;�b7�R1��Y\�"�;���]`���K�:ڕ)zq�&QE8��s������D�QS5�76|�ŀu�[�/M��{��"MUU��f�wr/��$�ڰ22^�c��������n��Id�� ��߮���x��� ��������j���C�T�X�N5`b�s`{��X[u`cպ�ad�Y8���}����ŀo��]�� 7Z~��j[$���i�h3^Υ�����;.L�4X��`����#��UT�J��Ea,� �wq`ۻp��׀y��0zn�(�J�j�%wF䓝�u�ʆ#G�����#�2FI$	�cc#c!!Gj�b�MM���ܓ��������;�bْЌ���#���%�`b�s`{��,���1�`��� �d$� ���`� }�� �M�`�=�,���+v���q`}��ݮ��mi`b�s`oI��_����0MH�3��yMCq����6��]-�8�`mR��UI\�L�\2�)&�5U �ݫ�2�k1��B��=��� �����j�q�C��n��`5������oP�j�{&�e�[,�1�`��{�Ň�/��+�� �����Yu�s�����@��B1���4��B_�	S��P��%3y��RN)�RIf�L�uh��XJ¤�1���P����5�D�^w������*X��<�ن��qdkyL�r��8�!-6E��Z�SQ2���bA�[i Y� ��#c8s��\B\Y��G7�Ї�}^k�||�
<�3�䵶�ZKw�Fn��~P�K5!Z�R�y�@ԁ%O�����Jat���]s����L��M�9�>��&$��)P�f�3$���K�qTt@�Q� ��4�u�v�'�R�TC�"PS���΋`� �g5�zܓ���rN�Z��j%�����������L_wf����o���J��c�b3
�]Vń�c�����f�`��I��5.�h�xf�H­45%�K���pB16���_>,j�b"�gE
�������76����:��{X�����V��)dl��ϻ�?��s�	�n,5�X�-��=�{a �i���[�`��ŀ���;�n��۳ �V�r�ܔp�rڰ7�	cݫ0��`yf9��p:� �@�Ȭ @!"� ��B� H2CZP⎔.�}ݛ�~���N䱓����p��� ��`� }�ۀo|�7��N8K)-VP�d#A��xsY�B%x��4�ѕ����������쑖�Ҥ���o�w��X��nޓu�'Χ�#[F䢰�Y�=�w��$׵`f��^�7�BM��~�Y�TWA�]� ���� ��mY�Gk́�����jDl��e-�9� �����<��{�Œx�PϿ���ܓ����\ދ�d5.f�J�V/c��s1�c�{^�X�8��'b��^�)�������h��(0�'7�cfI�.�(�E�$.y^T5����u ���J6�X5�lMqcu�ʫ�#ĸ�1�}/k��M;d�Uэ���n�A��8�*�Y�J�td���&�cT�@��6�{I	.r��	�w����bݎ��5�r�Үs���gq:��s��6ϚN��Ӊ�mru�;��{s���6���ٝ�Dh��d����*��q�1��;+�R������b!5��s	�f���R)mU���"�m��E.�>s����;.Mu�C���Ć�q��+rπ����<��X�8���s���vl���UG%%��{�� ������́��q{�s��#��1=��BUIOMSQ`k'~V���>�G^o{�����֥�:�ciRZ�?��rN=���Ł�7q`g�Ƭ��B�ERQXKl�>���qq{���/��<�۳ ;����QH��m�6��3 `S0���ˇ�7fk(�6�E��9K 1Z�(�!mX}�� �I�,n~��7ZX��7UH�J*��vՀ{���|Ax���)!>%K�-��(Q)	2 V�W[�j��E�c	! ���Q�=����5?]�ٹ'�w^0�ի�ӘT���Z�^nl�S,�r!,׷�^�=����:��,��I'���`׷x�j���':�l���
j(S4*&�U4X㸰>�G�tZ�L{�� �Ax7��7%��dv�����g�ۖx�a��v)s*���3bE���s��9d�`�{^��ـo[��9A����y����
T��Ԋ"��Vz[V�w�;�̜j����&)�'PTL���V��Ł��vnR$H0�D
0*��{^��׀|��dM�m�8�Vȅ���`f��X�Ƭ��,�6'v���Z���V�'���(��z���Ł��\!(sqS4T����d-��mVʖ��/X �&�KqnZ:h�!��v�7l)շ�7���w[�Xd�V̄;��U2���24���/脏n֖F�׀{����j�9h��r�����,C�j��M��n�X�;iثs��9c��:�{^�M׀{���5%������BHK�$5�	H�`B2HR�L��HЁaА�!M0�@�!"dhA��� ��
X�hB[BF0i+HVH�P�B��$l�@�hc	�$�h�d��b\�,�3j]V��h�����!4Uh��#���u�M�=߮��kA*bbjE���,�Ƭ�w{۵����e��s�݂6�fQ	)��JT(3��,N[��9�s�8�A�γt�I�Z:N�Iس�P���E	-��~ŀwv�{̦}���56l�$���T�����<�2��2�`fKj�ǎ��D}�Ds��O�R�aB����_�y�;�{��`/-֤�Qb���
h�3%�`y�q`y�e��n6���ʿ���K^��ŀwv�{�n��7^yp�J��M.I>$.w7Ěہ2�֜.���Of�%����lm�Wh��M����ɶ�X	����n(�e(�H����������jأ�k�^"�����찼4�&�Xs����Jh�`m�3[0��K��o70[�s�v�Y�l�l�v؇�g��L�7���a᫋�kk���4r
ͶF�z�׎LORm�q�t���]Z2XJ ���&����ӹ�{��b�m,��7(��u�x٭���8�*:�$E�sV�i;`��p6�p�3B��(UU���3!�,�m���X�^��;Zs��
�i�fC�X�ڰ<۸�<�2��G#�5RKj�%0��'�4X��<۸�y���i`7ZXɌ	�Z�H��&j���r97w�`c���̇L�;��{�dM�ee�8�X�X��Xcs`cn���1�H:�k�$O^����x�;�����n	����u�.C=G��Pfq�ʋo��ZXcs`cn��x�r�&ZQQId���ٟ%�.5��Qq�r Fc�ŀ�)����3!����dl�Y�{۸���0��G8�8�����́�N4%5$T�
j����,7�������ZX����X�^��J�8젬v�|��`b�s`{��:�2��r#�ǶDĻ/r��+�k��`�
	���=��b����S�8�w&�f��amfߍ��ٰ3��:�2��2�`y��Z�����`�n,��M����0��,�mXff��*�f&ڰ��0wU��%ƒ�9�q���D`��f	B�NTā�"%cFQڻ.)������
 ����*���� �����bwmn;�RWmE����b��1f��x�,����k��X8�"��:���s�C�~�x}q`g�X���LB���>^N9��1vq�ͮNۮ �s �u�]T��M8�e�q;,���0����:��;��X�l���D�+%�;-� ������&�����,{6}�����5��2��yS4J���̔�l/c�>�^Ƿ�w��XM������0�{^s��ٹ'?w�7%@
�@E���F�`E�d%@(�F����`i� �іGZ�����q`�w�+���V�	�QS	c����T�ak��q0�ru�Xa�׬#�X�qfe�����Ph�5�(��o�=��`w�76W�́�c��bD*uIJ�&*�d��������X�l{Ł�}��Z�lreq��jH8[0�c���qf�8���Ł�vl��dH�@�Y�}�`wۋ �I�l69�D~���M�������QS4*���f���q`{$�6W�́�wL)L|�#�N)��nLjۊ.����� Rԙ�Ϗ�D��.1! ��>�.@#��B�J�e.eād?s�B@�ذ�����j�n���{E8(���BƇ��>���?0�w�[Y�BdY	�Fh�>.%��2����/��B25����0�@�rh�`�!� HH�쭼���OƉ�a�Rە��� �$��&L�fN�N;�8�Ca�3��d"�H��S!"bn)I �!m_�������������1�! ~�;��F���5��0aBI^i`l>����C�~MK�M��t~� BHĄa	F"A�dئ��_HL�n�~K��~�h�>���d�z-ނHh�I!��i�Ӈ�C�oF���|E��7o��2���������9aC��T�p��qwkq�v��ar�n���)$)��I�������]ݚ�*���N~Ki�����Q��	���6��������>ag�Z#	�ݿ$���GA(80bBE5�Ľ�v.)̝'�,��v�J�UV�T�*���K�U@J�UU�X��N�]UUUUR&m[Ka�	s)�	ٽv
�RGg&NeQx�sp���ܶ�Ś̘sR�^�U�͠M�V�S�A�V8���ۢ:��\�TK�:��Ӯ.X�d��S&Dk��W�\�9y��^-�s����1����bU-Ғ�`�Y����&����8���+H�60���p�z�{/m� ��P�,��n��噣��5�9J&��r��v��ۨ9=�Q�GUN���uz�<�T]�[�Q�Wm[D[��@�$%.���kc\O>����y*y�n�n�� ����VS[�v�Ƴ�̔[v\�6|���q��2�6�/H��h��kD�#�l�x����
��6	Hp��sF�re6Ň�r\WN�t�+(�˓	���"e��7@�n	�`����ܜ�m�ST,�t[�t=�!�"�hf�DҖ�vbRa�aay����8) y�[�[X�ѻ()�[r6��F	�ns�0��;�gY�����z\xvW�n�(jKݬ0x��M����*��J�J65e�8%e��#l;:�YՕ�Kk�Q��.᳅�&�nM�c�28'�t,Wg�jMT��ɧ�k=�m��dxˊ��+���q�+:G�;Y�G/6ױ�����P�H�^1r�Pn;�M�*�N�Mn�,-t,j�,���4J(tkv�+�[��+ƎÊ�<㱻#�K�5s=�^�z(#ַ<��qx�iV�0i�f��W%���Ll:el��EuӋ�cT��	M�N���'I����W�/Y�9&M1a	�I��ٚ(��[9��劙�0ۦm��:��z�k���@씘��#!�5E�@)��,[-�u���lK�M��Z4kKOk��6z��s��۰�8�-��O�b���;@)��Ŗ7*`8_]'�mkF#06ϲ�ų��<N�ruC��wmBjݤ������#H�1ؙ0鞖9Ԙ�w1�B5���7)xڪ���C��0ص��0�t�Bt�Γ��G��x��� /Ȧ�:��j�O�� �h�P6��M�'ȇ�?
p�*����>Ey�'$�?~�'�˩E��T%�̘�^c�Z^9��&�E�91�.�=%�#���n�j����sk\��(MW\m�#�q�s�B��s�Ш]�K��\����+5 %��0\��:萵w1j"�[���ڑ��.t`�]U�b�R�E��R�`6#4lg`d"4���T�*ڛ)�4M۳X����R�A6��f!I�`�K���K��).r�%�;�<��3M:	���)��Zl�ټ�\,�����b�]���sٻRj3�!�ä4����+�ݫ ���0�}� ��t���`{b�?��O�䰖�-�Bـu{��L�;�w�Ls{	��Ȋ?Ҍ�;�`���}�n,>�K�f��ǳ`u{!9�%ULȦd���a{�,r=������:f��c.��*�V�-�`�=� �s��s'�@������X��9�:�4�4ғo��ѼH�j�AMn�.�YP��Ā�D�UT��K���H�#<�J���{�X�L�;�w�Dur�́�aj�H�D©@
h�;���~Ev!�Z�O���ܓ��~�nC����l��y����%�7d��=��3%c���e��t���E̾U9dW��V���x��� �v��'���s�o�z3o�g\���r�P�e2����oN��q`dd�V���o�dk�0���-��`�ŊC��A`�6�M W<`�;���Ґ��J�HL��3����7q`dd�_s�Π���`����F+	a�S ��ۋ0�j�ﲙ`w2��D$ki
��V8V�-�`��� �}t�uE�� �	��3 Ⱥ���D!4֚ 6���rnI���,�#��dR�dl���������<���;��,6>�����l���Y��MX:�v��ۦ�wq`O�ـw��Xw�EG"�Vq�¬�d%�#%������@�d��n�ksڝ,�~�[��Ա���F�,�{��X��s`{��}��-ݛY��jTP.T�W	���2c��s��Hy�q`yn���n,{���U��x��`�wSnly��!f9�;�Âb^¶XZ�� ����;�n,�����ä�J[�ٹ'?gl�L�uJ�D��f��q`O�ـo}�����}�Tbr4�޻P�r�ws9`2� ��=k�!4�2Ѿ["� ��xf1R��
�c�jJ��5=�� ��q`=nu�ۋ�52��R��TTʙ���Ł�ۛ�Ł�1���dߠ���D��mڰ?���o}�����M���ۋ2[���QJiL�L�U5V����Ř������x6��3ʅʙ��J�,Y�l�w��n�X�;��!r9<�@��.�Z��qQJR�����F�[��۵B�;#�z^.+��.����@k�r�-�U+(0��.�����h��%K[� B�(��K B�u��Ѹ��V9ffނ��ֹ�ڜrq�L�y������)'�ewVM��� z�;<�u�n�e9w�u3e�"�Xխ�8�����z���ԒeV�8c�����ӭdȉ�
����'�t�om}�j�,0Զ�#;^�{2]y���d���n.�,<��U�ʘ�e?-�_��� �n�{����ٰ1��LJ�U�e�ڰ�ݸ}�� ���`��,�K������F*����[�cݸ�1f9��BX�n,-ݛ�$�4*��
Ԗ[V��l�;��Xɷ6�b���F̩�T��Tʙ����Ł�ۛ��Ł�1́�#�ed����b��6ID��<\![33f&��2�-���)q!��;3���K�����{wj��c��1f9��<�n,���l��d�Kdl�������$ڔ	J�h%b��$@�G�V�.!�~͘{� }�� ����(��x۶�~���z�g��9�"g�}6�~��T�5U9*���p�=� ��v`��� ｷ ���QG��U��Ik�>��,�B�{] �����V�,D� ��oT���v�*d�ak.-5��#�\��I�aB���%�0�!A��ߙ��َ���Vq�,�"�*�aZ��Kp�����l���`���{�p��[#��c���9m�N}�v�Iϻ���?�I ��i^-�,RI��H@�Ĉ�|�"	%�Հw^Ձ��*E.bI�T��5J���B����ݫ �c��7^����-�r��S =��`�u`c�Ձ�t��Cb�S�%7f�9��,k��n=+�Q[i��Z�$�O��zcǍU��q�W塍�X�`w2�1�V�Rjj�V�*���pl�y������������M��y
A�,Ee��UM���i`۫ �c�nl�q	�"�MJ	��f��{�V��nI��{��:A]�����f������ʬ+Rq�n w�ۀy���>��0ۻp��Hf��h�t�!�F6�pι�oa��
����r]r�yŹnI��Y�c�s��G-����� ��t�m�܎r9�7�`fCU&�P�H�J����:�2�1�V���M����w���p�.�9�[o�}�մ��V&���L�y��EU")M"j���q,oj�kwf��:e�܎�~����ާ�c��c�
�m�y�l�X[u`�u`v#D�e�f�̂���9u��Ŋ��v�r)�VLFwe5���z�sj��X����f#�sǮt�c:T�t�76ܱ�-�3ǰ���#�>��-g����eo) &嚴ѱZ>�l���ִs�R��7.׉E���Fp���[��F6S��[8]��,�:��>�i�x�����.^�.p�tc�[�	e��ٍt��؄��$�O�I��E�˜���˾e8�:�$�*��rV�ؔ�^�f��x�sK\�K����&fXܬ�{ZX[u`�u�������X����6�NYE	)�{v�}��َ��_܈�$6�"�ʊ��L�UU�c{V��Vl}ȉ�߫� =����i���nY�$rۀ�u`w2�;�Հ{1Ձ���*D���j�UU��t�y��] ��� ���`��`���`�����k��0��2���^��Y9�����a�P���F����p�����ـ}�`]ݙmL|�PM�u�$������E�yR�EB,S��?�!�j���rN���܁�n��$fɫj���R�RW))��17�`w2�:۫ �c�<KbS��*�US5Sa��r9�D��ߋ Ͼ�������ـ}��=��S��H�3E�u�V��V,�6q�,�9�}���e���"2���unu�L�s�j�L0�Ι+�r>� ���#߷���}��4Ҩ��5^ {�U������:e�u�n��k[�a	%|�G-��}� �:e�u� �c��BFl:R�U)DE�O��0����n�R���n,?-���m��F$��PoI �"BD�!	@���&X��B$3T��13�HL2@�G�/H.��)�)FKK*�+k&ëM�X`�)Bђ��I�#�0$1BHI$f�1%!�e��%q�%$&K��120�V��u�&]M�'�
g�҅.�$ddP��B �������m�,�)�ߴ�BBGD�9�C0�a20��k�4`X�8RĶ�M���K)-����,��F�m��m�$!HB3��M�c��I�XRHU F�����������*F2��B���JJ@�
a
����L%,%� ��!R����`GT�aFIjVHЖ��B�	i��x�Jʒ���!%-	R��$#HJJ�JB��l
@��&�d�B���T��(�D������&���,-���J�%��c#KID��l%�� ,c�hT҈~>8����>S�EE�E�SC��O�?*�C�
"E�=Z���
�mM��������}4��Pn��Fݔ��:��u`b�9�؅����q�[u-����	�m�{�p>�f��� >�m�?������E������Ե� 0֕�7�:(�����t�9����JZ��L�����~_���>ݺ`^:�r:�m�X�RDĩبD�ET�T�n�{ă�����`b��`vy�H�7Up�ʰ��� �c�>I�{6������vU�UE"�����3Ua�rx�����x�,���n�C.BڄE�[
O � ����[�w����.na*h�Tʚ��3ӍX����:�{p����y� pq	ƣDc��y�v��7m�K�����svu1Ʋ�Y�c�="uN��eu>Gl�>��,ϻ� ;�m�:��0��F�cuW%�7m� ������>�����ߦ���sr9����c��'��ܖ�w\�1͛Ȉ�%�f�=��`u���R�)���RSUa���l,{6��X����M�nj�uKU�[0�nl�y��@{V�q��D�$Ud��i���XU"Ed�� �߭;��d���չ:'2v؅g��`
�t��P��ۋ��-�v����ϝ�{��v]���mcJH4�,�MkM�[֚[l,�5�a�t�э�$�/�dZ]�fIf��KUu��`nu�cM���hde��K����u�M��k�T�X�p��v'a�a�ϓ�v��v�f�W�D\m��H��e��JcXk���6����ѱ��]R٤�4J�+�;����Ǭ�GD��{�.��n�vӐ�0�{k1[�vr�upuJ\b9Ŷ�t����e���9,�����{m��k�:��;��{�j�*��D�SUU�{����N5`uy���u`{An�s��E,�[p�{^������p�����"�:ZH\*�X~�DD/N=� �ݫ �Ձ�Ok�7�Mb���S��H�x��j��8��k�c�����;%9	�x�mԇH)�s��B��q��[kAE��3	\��]�s�:�7Fی����c��mX^�?s��GP��`{T����U,��*ܷ ݛ�5qs�� �E���T�~�w��$���[�>��k�\M��N�l+r׀|��6 �u`�:��Ձ�N!0���JQP�UUM��9D��}�X{�X�׀|��0n�:����K�� ��Հܶ��76 �u�Pf>T\Š[)�h��K�HWL]'0ul���2�u*�i��5���;޺���AMUt���VW�� m�����1�`~A���"��p����ٟ��s���wv�1�X�e�9�$k��m��uJ�)a%����� ;�m��� ��@�#$"H@�$"$�!HB$b20�Ec$1$���!�Ѭ#YFI�WK��!-��ɹ'׾�nI���v�����SP���؎s�K1�X�_���ـ�ۀwT����Y��X�2���s`۫ ��Հo���!mR�DBT��!Td��պ�{���yn�6PQ�(ma#�R\��0���*��:���f:�{Xm��>]�cЊ�-+$��0�����DBA���kۋ����9Ȅ�7��V��5j��m��o�}��Xϻ� =�m�<�i��ca%9d�[V�����XY�6��V8�Bh ie�"�n0�S0�)c�X"�̽�5�'�;�N�V�5c����ـ��{�ۻ� �t�r(�s���m��rg�]j���.5�'e�U�jf"mX�ʥA#B0[j�;
��2�0��� �}� �wq`>���ƽ�-�O�ʁ��`�:�:۸�:���f:�<�p�%�
X�U�n����>}ݘ~\�!!��`�j���C�tP*�U%BUQ`uy���u`�:��DG9ۻذ:%hLRTT�2��l3X�rc���ۋ��́��F�A��������D"����J�0m+p�Y�����<����v[&��c��ф����:��N�#�!x�m�@��4���U���ih����1]�n�ZihV7�j�a+PĆoSc{=Dp�c-۫����k�v P�vH6�N�@`�+�/^M>'9�SP]t� ���HK�bg��
����uj�^��H��ړUc10�[��A��<Vm2أ3��H��,���;��v��(M8��x�A�rsc��ܞK�l�7VƊ��Y�����z��b뢖�5U] ���Xm�X^ns�Π{p_���M�l,��n�����9��G�ǹ6����V�#2$Nab�FZDՎڰ�wf {�ۀu��0�ۋ �M�kn�7*�2�0�����VsŁ�����`�2[ �G*� ;�m�>���������͗x����J�z8��F���Z3g�#Y�k�5΢Ҥ)e�S�����X)c��V���L��ـ�ۀ��|�k�mu�l+�� ��vg���.qT��zo� >����3�K����?�n�2�#�� �ݫ ��Ձ��W���*Yʪ�5l����n�m� ��vl6"9Ȅ�wj�q�F�)��IT̩��1�,�76��X����I��J��v>[�����^Q���5�S�v��v��<r �n���+��Ġ=TT(��h��v�ͺ�{v:��ڨ�mm�㒪�Q;-���@ﲬ{)��7V�$�UETH��q�p��f�m���8�%��5�'9��rI��{��?t����V
X�u�0{n�ϻ� ;��������<������-�vZX^nl�rn�t1�X��`_ߏB��ƾ�e�˙����z�LXeNٻsh�]�=��79�8㞘ų�
�̪�� �n�/c��X^�6��X��ƭ�)m� >���L�:��lu{��BC��jB�P�D�T̩���֖�c� ��X�����{��7STvS ���lu`�:��s����Drb�/oL�?U���%C�F[f wwn��s`f:e�w���~��b��H���۱�j��Rƺ�%�Mzw��d�pǢ�*u���7 
,Y��fZa^����z�m�t� �7[�r9Π3wj����viM!��m�� ���{�p��p�{n�Χ�l��:�dvZ`��V��XsX��`w%�0�S���B[n wwn }�m�=�`�����jBjcV���ۀ{X��`�u`mՁ��PB�(I��h�O�߮�[�h�d֭,b0	!B���H��,R��0! F1&1� �BJҰ�B�ʐ¦�2�C��L!�:#��A��gĨc�7��9�ZM;�d$��ɡ��t:�����e�2~����:@�`ȓ��-xJK?h�O1�I�o�X�X�����d������ؐ�D9��tsl',�I�b2ђ!ĩJ�b5�c,"�en��?r��d75�SL�HS�&g�8f�\_�w�D�Y�ľM&�^i�rjx�����J�z���s��|ƺ�4����L?Mo��Ns���}Sd��<r1pO���i��I5�H��&�e&�B�9;Ri(O����b^���rcGy�N>#�X�uX��^��X����Ffx �( \�s�]�p�>�>��p�g	:~�~�9I��Q��n��Jc�??ӭ�2��%�5�S3L�).����Sa��G?9q���@P��Ԛp�������l�y�M�J�M���N}VR���M�$��I����S[�&�Ɩ;m���9��M�������#ȌDs|'3p����P/�}򫂮#��G���2{N���&%�%��J|=[�s����+[UUT��+U�R��U*�UP�
ڬUUUU@@UX�u����ݠ��݄���q�
�a6U��(1��n�ɬT��嶐3E�
E.b�Ux:�q��9�C��S����1�n�m���qms��vb���8C�,��Gۍ<Hzi�34#cͥ�Q�\<E���	�Iu��,j�ęև���cvN9�ϭ�-ifvÅ��ytH'n����H(���s�\�U(</[�m�S��x�_T:u��R�㳻�΁��cغ�o1h�v�Sp!K�X��CͥKj�y�kp���O�P����@��r֞�U
��כo��i�i���=�8�*<����;LW>!)K��4Ֆ�����h���[Vd
���5��<�$�Պ�`�Gm�pM��YBf�ʌ�;XVQhYA�Ca���^k!��u��-���;vLW'+�rgJk��`U�-��sG��<,�rqڈ�4<R���2�M.�e�BEQ"�K6����i .յ��PxXC�k�@��g=��6u��o6�Z�d�]�,.Е0�ْ�FX�l�,��ۡ:���(:�%�<�;a�{Cɴ�ld֑0n9�(�.|�9��회=�6���q����m�j.ɮ�ػѝ�lnF��)��a�0�:JIl+�v��M:����m��DN�t>klv��S�*�}����]�E��q�l
YR�Xf�u��B4c�PKKز���,����kɻl��Y�c4v��5㋥��b�e�6��S�#	�\M�0݆	j��n�p΃�˶��vy]![�J�&݅�Z��7��>qqf��s�s��V�d4�n�Z(��.Q�jEe��هt�3��%\��u�.�[.�7#`Kkh�k��1r�g��w����b��j�S��j���g��6�0����Ş���`�Į�Z���F^!)L��.���<21s���v7g�.�f��9f���+��i
��.��!t�֌ـ�8�m�<�p�P�])aX)�zwt��I�:I'��AC��R�*��5 >>G��+����>`�~_�'�F* kZ�v6d�.G%Մ)9�K>�9���e�H����ў�;L�:Bٖ�8�3\��M=/�U��mۭ����C�ӌN�^Kl�zt�ꗔ���;`�:�&�kn�c�q1m��u�×��t�Ot#��n6M�t��7 p� �l�	�ov�v�P�8#��0v�V�u�s�X;��+��h[���$l�1�88����p�ʳHYGE��R�ˈ� ��S��OG3�Է=`蘸ʹCi�Խ�]\0x���b�tb���Bj�m�|�������{n wwn }�m�;�-�3d�Q*�T���V��X{X�t���q)�?U�[�cuT�Q;-���U�g�՟s��I��,���<{r�T"�T;n {�ۀ{v�x���I��X�9����h�5U��X�2�������Xs`��AȤ�RM��q;eM4J�0"Z0hY�+F��J�3��<kE�FN���u2�T��� �c� ��XsX�� ��X�%�JR�k�ۀ��?.Ѓ���Qq�~(]�b��d��7��9���ܒs�w[��keR~Pj���p��� ۦXY�l���nƢT�2�ETʩ���[�zXM��mՆ��}��pyMr(��I[�j��`Y�l���;���m�,�q��ɔ�U�Di�6�k�32&K���ZYX���]�[�:���\/&�����;���m�69�u�ݛk�r�T"�PN;n w�۟���ǻZX��X6����q#� �JST��[yG-�7������p�q~I�S��cCȩ�MI}��ܒw߶��甚�Ց��� ��v`mՀ{1Հ�wrZ	�S4T�j�fjl����B�����ŀ}�ۀk]��+U�H��e(���X.�a`�jw.���d}O �	#���(:X��n w�ۀ{wq`�ݸ�ݸ��S%���l�In�n���	�v���X���z%��3I!\cTvՀ|��0ۻp���ۻ� �OU��e�N������Հf=�w�9�b�)BI$`��(�J��]�JW���;�=����5�����{X۸�����u`v~}���k
\�,I��Z�9��t�\����<��b��8�ܶ�r�M���Z�D�U����;���3�Հ{����Ũ�Q$�U�;*���s�\l�� �{V<w}-	�5J���MR��� ǎ���VlDBO^�X�v�x��
��J�55V�c��w�7V�n����ښ��P�[$� ｸ���� �۷ ;�m�>�.%���� ~�;�kN�a��.�&�B�, Z�m�����O9�j8�6���#e6�d�qӵ�e����Y��+U�hhٱ
��K��RM0[Qx5�ڱ�C-����v�Sh�f�;!u"f���3�w �7a@�����n�fF#JC2Ys��
6י\��4(��)���w	�5�&��<٢z9-Bo=n5�R�^VX��`�2�L+2O*"�ڕQNN^9#3$.S,�9�ڍղ��5�� �����4P&*��0�iBi�B���b�2��Tv����ۀn����p{ۋ �OU���ʝLL*�� �n��s�cڰ=���v�丛=�[���,�(�ۖ�cڰ3��,�n��:�:�2YC�t�[yI-�7}����� �����I&���p�Z�?��uV��j,�n��u`�:��q`�I��Q	[b!��l��<�M�YҦ�[[��M��G4��[�[iw*b��Qg��L�tu�X�X㸰<��l�6:��u�J)e���nN>$���Ȉ�
q�X��x���f��TXղ�%�� }�ۇ��$n�� �{V}$d�f)
(��� �Հ7����Vx�,��ZWZmT�,Q;-��m�?.s���{]u�ŀw����yԹ%D�RR�ͼ��]dWa��e�g�z�"^9V�svKP��K�ӭ*�6�a������V�w�c��Du��VlK'J9K���In�������ݸ�}� �^C����uZ�qʲI9���rI���n@SI*Ԡ�X��5>X(TH ~UF3=�p��ŀ}٬z��v�5-vZ� ~n���V�;����%�{V��`Ӭ��댔R�p��n�����������*rA�&��B~<�Ֆd*��lXL0�5��vK�PLb�-�b����eR�ȭ��-�;��X�c� �7[�Ds�cڰ<�2�S	�*UUE�w�����D$7j�;��p���ա`�U�;Nʫ ǎ���V<w�c�<=OE��PL���\����w����'?}�nN��H$,���Qx�7��u�':g�;5.jk��TBSQ`c�q`�:������X���Ԗ�!*er�-��X8M���nuZ�V��k�Q��vb�n}uح��
*��ʚ� �Հ?7V}���y��f��"��1�k�ۀ�ۀw��,��,��W��C̈́
-DK��,� ��,��ŀw�p�ݘ}�6+���VJە`��ŀw����m͆��B�=�X��2	��Q��,vՀw�p�n���ݛ�~��ٹ'�&�!�k�!@B0��!! BC_z���s�tM�$�-�f8:������k�WnÇ�z�nZp\��ӝ���84ud=s%��y�gv�.3э�2ۡ�!Mnb��l�ˡ�b�����fjB�6�.M�s��6��
s�D�`�i8��v�[v��	��"[`�jn�;��]�$F2�4�m�l轍�4e�sbj��3�wt:�on�8�X�ۣe��[�g��v�褹�J/}t��ﾓ�A���fCq�uR���t���x�l�c��4�GEXg<��S:�cjY�neHMUU��}6�����e2���s`f�∴r!�
�l�;�n,��� ���0��f��Y4���;*MME���e���s`ucs`w��,.�z�Ym�k�Ii������0���`w��,7�X��`{'P�	�UR�Q5U3U6Vc���q`w2�`u{�{ǖ(�܁��,䅴��p�	��q/7��l:�T#l�������&�Lj�c��d�to����}(��Lߖ��xIr+%mʰ��hc �h �E*�̛�wٰ1y����/�"#�H�$9�!j���"*T��{6Vc��Ł��� �|�аe��)	l�>~���Ł��e��9���j�lz+�c�PLr���q`�����n n�n��b��r>V��dWLV�\۵��a)u[�kH����)�����
KdC��ܫ ��� >����p��ŀu�C򚥬N+\�v��c� y���ŀ��}.�"�X	�H������qa�����_'?m������B1�&�-�P��q
!�5������0+1�) D�[,��]�"�Xa6sG��3	�1cLe�#�b�&�N�6�M�#~$�>���O��9���bna @�A�$"im��,	r܄q5�B@�}gS,������� FH2��z���:���a���ci��d��� �pHA����|�_|���E��&^3HKI%�@�eHh�bF��D����i�@�!	�e0�%9�~�?mG�����A�~%�� R Q��Y%xkLdf�.��$���A����T��B�RXЁ!H_��S����g	�u���O�J�H E�C�7��39 �?RL(�t\� F$�Sa��Be4~f����?��FH�d�~
Eu��b��8���Y1��Q�����z��`T	�k��"Б�ֱ��	��J�:4��1/��\�;�S��BG�ҖGK�9&�CnHNF��8�A4�h��6�ظ��Hkm)�� aCo0X@�ZA+����T�r�+�ɎؚC� v ���+�i�	�?��m؉v��> x��?)�FE�����ڢ�Mb��g�ק�,�����䟴�?��T���ۀ}�n,{�K �Ն�9�%��X4��7R��b��`ݺ`��� �{n�}��y�����UyTu�Q�Jd�V�y��p�=��vŜ��c��]���$�jP,���������q~\����~����W౵b%E�'e�玬�Ł�8Հw���"8��o��vI%�-�;��� ������n }�m�;ݣskR["nʓv���N5`�:ޠ<�Շx��
"1.����#MPu�*E��XI�"hUv+{��f��H{#��M8�r�����n own�|�,��X�Y�(S�S$�BW�{6��P$'U9���k����XæIfŘ�HM��",�R��~ ��߮�}��d�[����1�P���U��%MU��c���Ds����<�������	4����j�R����5�i`u{��u`w��,��L���V�T�:�?s��I�{L ����wۋ �v�x{�V����*,Q�jl:��X�RՁ��s`{�������6�����!E*�BfE��h��]���0r�@��x�L9�ێn����4)�K٣����@f�R�FK-���Aĸ�0-Ŗ` m;#(L��uK`���6��Ӣ(�s�mzi�ر�M%�jga񮂴Kn��U�/�ZH�����sq�iK�f��Ō�ƺ�����Z[(���ge���������[
2��Z)?�zwN_ܜ�;�N�d�mEm���.ۮ��4�n��+Z2[<�,�E��;�gA8��J�&b�����cߪ��:���c� ��n���Z���v^RKp��Z�:��<u`�u�Ȏ$b���v�qZ⩻+�:�L ��n }�m�=ݯ^�a�`8��BjX䩰x��;����:MXY�l�pi�,��Qۀ{�p��k�>~�� ��n���@���F�G�,k�*mk��r��5����b�,"�r��7T��[{��zum��s`�Հw1Ձ���050L(�kW35w$�����)�" X��dH�Ԍ$�)������9�9�~����nIϻ�� �|�б���b�v� ��n w1Ձ�u-XY�l�9	�DҮ"ESn[�{�p��k�>~�� ǎ����S���*P��r�����:���6�XsX�f ��),��Ѳ�P\�-�Q��)t%M�FREI�)h�H�5�%�c��KMр�]ɽ� ��XsX�RՁ�I�bRҡ5,rY������}���>~�����x4��ʫ%���� ﶽxN�%�\�ěI'� 6���  �����nI?���lC*-t�j[$� ���xVc� �n����N0�b(HDU)��`�u`|�ݮ�{Ձ��k�=�sT$�#�E�eV:�,��Ե����X��U���f�E���a�C��	-�RIn {۷ >����ٯ >����6�)Ybr*��� �����:����V��Vq�*]T����yI-�;ݳ^ }�m�w�p��n�ٲ2�+\U2����V��V�c�B�8D�G;)�ڿ"�7�]�?_t����SPT�U�{1Ձ���t�� ������r}���[lb UF���=@�K���ͱ�9�rch�#ƞ�
�����6��䬭�FJ!�~ ���>� ;�u���,{6n�Z�nJ�R���J���"�`�:��9��^�.&�=_�?6�:�d���o��9�b=�j���j�;�P�T2�I-�R[n��ـ����L �wn��&1J��U$�`{X0�X^:��9�3�8hA��k�U*HXJ�BB.R�/y��e��ԙ2AYs����x���2�ce�[e�����m��մ���Fy���(a��=έ�̳]ah��Z�Z÷V��%�V�7������� �n��;�ᡌ�K���cr\�6���R:�1��b	c��k�7"'r!D��x�7*`6-y�W[v��6x�g�L��ۛ�JE�.r����l�IU�c��ݔz(��rk5.�O���P3��s�&I�ɔ X�J����r`���X�*�<;�b�::��o1W7\�46K�������� ��V^�6��VL�u*J������ �}� ��l�w�p��׀|��b�T�8J[m�5��l=���	kt�X��X�Ą�&������`����[���p~�����l�J+b��c���M+ ��VY�l=���ss��kyM,4&,۝�Ы�-�!�t֕�5ta�v�PҍdPtU��q��&��� �N��K�׵`5���3��z�q֥`wv�ջ���b��ۀk��d_�~Q�š#�mX�F� ���b@���T�@�h"��ł�`!8��{����k��X��]%J��3!3U6��V̧*�:�Հ�c�۶G6YUTnJ�I-�7޻ }���k� �c��Cu*J(�J��&�U�u��nl=���w& }�-M�|����3*�J������본�-����*\�K�F�-�:��^��໡�UUTtOvl=���w%�ה���l�1E\�d�� =�m�����)�X����R�QQJ��p�ŀo}t���s�BHH��"D`�``V(T %(�H�`łiR�I?��~��o�|��b���*jJ��;��`5�����s`?at�>�յ�B�XYT��L_we���̀��2��:e�����e2vJXr�汳k`Wf���[�M��y��t�dg\��B�D�,�N3�^���������`g�2�k�*m���rV"�f�g�����n��۳ ��l�5�7l�R��X�L���L�:����,S�l�r\�>�lC�I�[i���>���`_wٹ'?}��ܘ�+i
��`S* '��%�3��ܓ�{d�͘W)Y)Gl�<��0��t�=��`?nǍ���Kj_)����n@�}c�q�q�9�bu؋�Fļ�J4��(2�,��f3JS�L�]������z <�-��Iz]9[��;2�s�g�I,�*d�I\Cj�IK�����>��?M����Nu���%�e2�bfR�m��U*I����+{����: <����Ş�q�߷٧�6��lAe��H�	��V��s��D˭{=�IbiV�K_���?oq���C��T��,�5=�IyL�I%{Ȉ���3I��)[o3��g9m��
����
��������ꂠ��W��T_�APU�PU�AG�� ���P��B(��T ��P��B ���*�T (�P��B �*�"!BAP�(�T"" B AP���T ��P��B�"1T ��P�(AP�
AP�AP�B ,�0T  EP�$B	B*�P��P�B$$UP�AP��P�T"0T")B#B AP�T"�"AP�0#B�T"B(�P���B(�P�DT"T"AP�AP�T"�T �U$�T")B(@T"�T 1T"�	P��T" AP��EB�T �B
�P���B+B$U�AP�B0�BT!B0T �T"�$EB"�P��T")B
1��P�0�B)BP��T $B�P��B EB ���"T �B(AP�DT �P�P�		B0EP�B0�T �T!E�BP�AP�DT"$B"�P��B��B @T"0�P��T"�B ��B"� � �*�� �*�􂠪�AU�*
�W�PT_�APU�AU��W��T_�APU �*������)��d\���,�8( ���0����*|�nX(*��s^ƑW��Q�p[��M��J��[5"R��m�S�l{�z�/G@�]{��QR;4��iU�R��Ka�� �V�4 @Phd@RM�:
��E@ )@l*��EP 
�R���$4<      )�۰h��UMhg�j��T����W�n�&��t��ޕ|��$�=J���ڗ�Ή���_��ޚ��%�Ы����\ڮ �i����x�֯��﹇�X�6��{�嫋T��[Խ���i�*������G����z���}ު�� >��ml%�4�e� ݆����]��*������ە�����T�T@n�Wsu�=�u�j������U�$��uU�xZ�}�< PPM��=��	X=Y�.�w�U�[�Y}��n-t�w�U����^���f��\f���W����+�>���>ڄ�����3v]��x����>�w�t�zo0B����S�I���l��������=�=4�== /�ܥ=4�� ��iO@ ����z�@c����J �ܠz �g�z1 � oY� pt*]�ON���(��� Q����JB�R�p��ѧk(���cZKǻ���t�@��F��n�篖��u=��<K�&�)nn�i_{����(nܩc�>�;Җ�|�S�gC���f��ry�ť9
=�ݟ^��g^�-+�\ڕs��U�q���R�����u}j���z��R�>�����vi@B�P�JU�e�o>��}i\Z��ﳥ�s�J�P}]{�S&�}����O�ܫ�{�s�>w�Q����K�n������   5ϷKů}�*������=��쫞��Ǿ�G���}���]���y���y5��y��_v�+�   ��B6��   ��*Fʔ�  "{J�'� &&���5Q6�U= @��Jf�)P  Ԥ��������Z����?�_�3��}��>�>��TU~e���"��DTU?��"��ʀ���TU`�**�?���!B~��փ�����"E�OVYXN`��|�C^��	|z�����P��9*L����}�^Ł�����>�!���v}�b�:�N���s98�pN�w��Яp೽�/�AZ`(1��&�ry�E���,R����JC�|�K3�K�ۚ2�R���%�n!sD��ާ�^\^��ĵk7~����p���=��Nk0��y�%�<]�)�'E�CȈ��|"Ug/>��J�N��.�Q����;����!-`6�l����!���e��U!^Zq���cn}�`��R�������/7S�)~J{.pg"�Ƣ8���X��Ұ����rϧ�߽���dgQ"D�1xNa�"�(Z��O�B�ňX��r��%���G�E�'"�B��>�ŧ�y&6u@@�����"��*�5����w�:�3�.�!�8}>��q&�Jɧb�-��k�5�<Iӛ���ƈ.+�dA�}���p��Wbp����v�Y9S�2��}�˭ǈ�j����G�o=�o[&
>ɽS�]m;5�9�⹾��'��Gj��'{۱.����}�>��x����5C~��%(�;��O�w��k�7ݬ\^B��m�h��S.���ڨ��r煂R�>�e��F>	��
��B�}L�>�=JM��K�_]|0<�c���zd]/{ӭwW8�ġϾ�Zn_�R!�NbM�D�4TBBD%J+����ö�>�#�|x�/����s�!&��D/��y�ć>�ӆ���#��'�P�!"bC�����;�'���th|'��d
�M��Þ ���m�ɥ�s���ޝ�.�8��J�<<������@���&}}ڑ��<C�<�> �\H2��:�Ј�/#�V�qTT����zg'����9�X���)B]����t�}(2�Y��	=ۥ�/M��,��Gq�z�=�8:����a�sG.�C����e!cX��Y_5rj��״D��gb��9�;�qU�N�~�o/��k��z�<��,�w�pw=���x�9�#5����uLA� ��D,�m�8'/|�:���{��0O�#�+��߹��##�*��B~j҉�S3��TI�Ϻ�����{��C�Q�X�T7�!/f!9�P���$�|�s���g<�ѳ<#�|ѳ���o��j���EֳS\�"gE!Ȏ!A�@	�ƲU�1�O��}S��3�2Y[�24�����!L�!��=7�xFƜ��.�ޢPŐ.�!�2��n;HC�Q��K
f�bP�c�U_/��#�!�d^�8�P�p�u��I���{�������<[�\)p�%e$�n�%x�X1;���ˋ�wdE���r�O��#=��*�^�xAgH�'U�>M�1,wB`�4��rS��]�BpQ�zF�w��5�\6��"�׻����)����LZ�sI�&�j��PA3S��k.� �x8`�3A$�z�oh6Kq�>����22j�XQ&�#��&�F��޵e�����g#�	�erW.��)�2u$O�X�N�wFa2bd!�a���7��x��k���R��~��]�f]l��h�r�N�l{�� )��S۞Ք��s5��'�/����p�f2z-�[�� �C�&w^ׇ�/q�^��f#�X��~zO'8I��p���G5YX��|'��B�j�f-O�W���!��Q:�v�f,>�xN���|�kTƟ��6uN��(g��9�/����>��2��?zη=�̶3Me��M�і��ya��{l�O��۲}���/����b߁Yh�����>������yNCZIMCG�ͅw
a����o9���x���C5X[�wu��M��$	�C�`I�0k�m \����h�B�4º
���W)��q�e�f�[>i��$B�*�\��w�h*�{�Ժ�Օ�T���i�Ja�$,��X��,���N+�X�#�ȸ9�=
{�S���'ӎ=<=A�)�x���-s�"����ƴCo��S¢�}��ώ�
�%��W!�T80 l b�$IE9�Z�\&}ȓQ�~�1?�y#��!	%%/�ZD��\3L(4������BK��չ<D7ψ��[�y�}���1)��Ɠ�ĩj|K�E�!47���&/��rV&���#��<�FA�b�G�������"��v��)W��h�5w�s P�c7�Ӛ�2mx�)�2��	jc�g"E��4��\���93�x�Lߘ9\��7�}�S�7OYsi4C�Saɘ��4qa����9EBs�xQ7�N�5��_F&�m��>�{wϹ�}���<��W���{?��7��򵒌�j�A�w��	�u.��u�#�w�B�pw#_r �,8r���j�{V{��]��ƞ��~���./"O���UA�9����M2���~����I���q}3ʉ��<�oj��&�Q|����1X�o��|êAj���q�{��f�t�J4a	!HT�Ғ�1�
I�	"���8z������1�s�.0�x�]H�%S��8�}�a�VS���g�ٶA���/D]���\�/$q��X��R�Aī""z��`����G�ݟ^EG_:'{q�x��o��ҡ�1�$aY�aƒ�ޘK���H��B&��]���T���Ssg-V�����U�ˑ|�C�t�Dg'��%�����<���:$#x4MМR�֞����>]ߖ�ϖ �U�����*�X�d�/��/�o{K�����8p�Ce�;�f1);WK����߰�N"���FD<���F�}�ڢY�U}���K�R�۝�DΡ>f}30_}&s1��Ng�;��p�0���nÔ����`kV�$d+i�$ȔM"W}�pB>�ru,\k܏$ל=��H�%1���g���I
D�52I�iaS�M��b �R���<�B�յ�g�x���w�]��a�s��Z �H�%8&���� s���y�]K���8B�`xi3�Sr@�3���h��]����f�1�BČ���T���$�eK~���
c
��p���\ֳ|!��JἻ���}���1L����pz���	�W[�rc>�XT4H�.�!��L��8Gb9���G[�7bS��!{n<�e/5~NO~�se,���$h@�1)<1��nf鱈� Sщ��m�xy���[���wpԎXq��>�.}���5�5�۫D��0���!/�В� ��S8�v��2�v�� �q	z/��;|�9�/N8�o�{u-�g���znd�����@���}�y���Bq���=�焾�g�Ow����%�-�-����(����.رW5'��<��u8�� >r�sv}���h���]BS޽S%ƃ��>�\뫿v�j�|���}�w�>��ާ�ޤƉ��-X}����0��$�R����r�y���J|+�r��'9L�4������׌��L)�6��}��5&�S��:��_�Z�v�j���1}�z��:���H�s~\W�ꌉD\�=|�����pp�(��O��,�س�.O��iy�ʝ��j>Q<X����ꐂ�����'�|B��fr"�dJ���Z��{-	t�;���&�{����/�k�zyq�g=��A߽��v�(�K�%y��� ��|�2��2��/}b��9I~�用��o�yMK8�⻏�2�%�ƽ̡�;N��&��b� ���	�Ӂ�B���Da�l+���4�d����.�n:cH�Xj�L��Vb_/�qt�u�*CHA;N��]X�}��x�V��(p��~�3�Q�K��E�r'�[����+�ń�2l��g>��g{ߟUI��Q|���RS"%+��$yY.{��Ł���l���G~��菲����x?��κΑ1|�"���
�quv��Ȑ&�$��p�֭��<�3��Ѫ^x^J{M�1�l��)��Y �Jf�D�i�v�*`9���G�����2\��mD}gR>1��x���m����i�����o�y�h�>/�!��*�rE>�.!5&A4�r��N�Ng�#c��/��݊&�)."Չygw������Uc�z.�}�^��Ş;9}]���7�=W.�}=��h�Y~�׾ʚ�fN��7����{<���X��G����\�#�ɇq_����?����<x��R���y���5'�Nw'jS� @g�Z�J���1�����%��]}^�{�9;|v+��`]�<�8�	58��� �|P�4F��&&��W��{57�U��}|��=y]~�2*�4��(&^��fj���֏%����זpH<���N?�9I�^�oD$Z�nH]��WiHw��$�M�H��G�׋�A�;%�L�D�T숨#}�W����q �$dv�\�bS������v�!�IӾ|�w�3O���C�Tu���2!�K[=�x����ڱ^�;߼%���j!#��*,���X�:MuV�)7�y��R{�˲K�}}߄�c??԰x�l����Oø�O��������!s�ߗq�!�q1^��O�2p
�����
%U�|�M�g$O��"~\/���3�s��1lL��Ȫ���/<{�{��o�%��K �!,d��҄�����6��f�<�I�=�[�|8���C��萱�M`6��1&����}��^ָ'Ə���/��ÿtk3�噜BE���4B1!(\�[�I�%�y!/��y�|�)�,�������I
2JFK#H��I&��e���+%Ƅ�,�>���o�~�f{��w˟3��|b���"h��3x�awC&j�m簾�C�N<$ �{��:rf���Y�,���<���b B#22G	/3>Qr�.Ϣ0��,%���}�ھ��Q�&q�Tj4�p s�3�D�@>I~E_V�����J����a��g��Ő�0���.ZYƆ5��ߟ����5q}�W��6���l-e#@�%e��+�9,����Y�$��2��J��C�M�˜�pL<9_����'��nN�!���7\����γH��3(�x���TNǚ����m͏B~�i���@��� K隺	�DC��߃�!L�xz�B��ńhAlϹ��Ɛ��
*��$TE�;+E��6�������ϐ�������9�4��ˏ��$(F��)�Yl��M*p@��	<��!�&��pr�B�ʯӟ?g~XЂq֜�q%�BJ�A>|�n9���5���dC�,#{Bn���z�,]YHsˈ�y�b;����5jN�H�8�_.�w1���M9}߻����&|�K�ʔ��|��1xBں)���Ϯy�g��B0\a�����|BN(�c+�q��|���pqr����Vy
^�}=�<z g<���\\Bh�RQ#3�|uD�}Ə�.Z
1<���P��l!��!/,����;~D]3�懻���4.X����)�l�q����h��<<���3����.qyC�ǽ��rV;k"[����_}>�y$����B�i��钬���	��)�RML���JHK%�8�'@#����G8��e$��k2��a����y�I�������� f[��wm��UUUUUUUUmUUj�����������UUUUUUUV�UUUZ���������j������������UUUUUUUUUUUUUj�V�UUUUUUUUUJڨ
����������*����UUUV*������*�����UPUT�UUUUUU*����UPUUU�UX��UU@UTUUU�����������*�����������W�YV��b�V��!� �1ò�m�6���ż��$i4�16zX%V��ܮˉ�¨p�����xc�3T�\�(�24�նB���gON�Om�Pc�U�k(��6����vR�ʕ:+��.�/�i��p�2����`9H�<�Sk�88���KV59�`n��vq��`7��lX�q���Y�\f���g�.P�%�0'����|�C�P�iImn��E8|�8�)�k���3��l������»{MW,^�e�-�۔X�m!n��D���`�(������BV�n9]�n9��3�:����h�5��j[S��j��5v-DU�guo�IÖ䒔T���T6�\v��"�32&���K+�W'ݹ�:���s���mKZG��� ��^ĝ��Xf�-t��G�
	���ۂ�g��5ʨڤ��iz���j��6)CEi��t�]mPlU���]j�vԫAwTi�/ê�nZ���e��6�r�����B�/T���[\�yU]�Y��&9�Q��㬪+�-[X򻶖�jCl
6���6��*�j�p�T;O��u�k��u&;t�p5�S0�u<۷*�HƇ<��������TS��[�!�Ǝ�J8�A�[ٶ��l=q)6�`��%ܬ�r��A�R�0�::���z���s5�v�rVex���5�`S��A6��vmC�]�qr;�@��������m(j��q�`vnU��ۏ&H*4�v�Uj�j�8�T��l>8۷k�ثtl�zb�i����bw8����� � m5�{Ts��Y�l��������40�٤-�ڌUB�:ܥX
���6!)�z�x�%�f�m;:��ϵ�YC&�Y�����f�6;�)®�ȫmLN��#��u*������u���O!r�dv�7N��q�|\������[��a�]���J�El��@��X�8��%p��rQ��qь�]d6MB���[b{&�m2Al������9Y�l��r�;n�X��Ÿ�Ѭ�}<�JzDM�L;v�� ��oY�uMmUK��T)J+�մ��)̷�u�]��)�=W$[7P]nĒvj���е���b�9PF�� \k���m�Mm2,u�^UVe��m�;n8ڬq0'�H��D�+�-�LXZ ^��<ٜ��ky� u���݃ƆM��plF�x��iUv�����UGW*�U�H5q8ȀX��+ ��;v�i�7�g��*7b�IU�&,C<H5Ҿg�Mv�D2�Qko(6��2�7Un��v�wMv۰���n���w���B.mbK��^K{m�^�s۷!�
a�lݓ�,^Ձ��m9ܼ�S���Ə��
S�=�՛J|x�n#�|g磷4(���3hBx��u�����zz�kK� 5̫�*������y�݌˶�x�k���҃U/���j�i�ó�Q�u���U�a��Ue�Uf��-J��[��3�p�1&�wqXs���؛K��c(1;�<�J�dp��!;��|:�cs�g����!++	JM�WmeŹ^Q�Qj�\�whb6�-KU	h_ ��k�!!�\�+�r�}JO�(L�;lup��U���C��c�NX�ե�h�:!�Mm�����f΋��ki^f
t���P�tٲ�v�Wl��k�ܗ`�%΃��vڻl=�KqƱhT��c����X�ƪ*�� �t3��d�Éa\ڳaxՠ�p^{/oe08���F�M�Ӝ ͷ6��C���e�f�;^�㹻r![B�:)Wnݛ���j�SRśm��u�q�`��9$醵�ۢ�%%x�iT�ݹ�[l��U�����.�M�J� �6ժ͈�M��rq���l�pWNLM�Ip�*�͙&ݥ��0��@¥���b<+
ôֵiT�끪�t�g�v�cYd�u��smܜ=����\.�X���ksB;F�U@�KJ��0C��ui�wO6�$l1Wm���nn]�[��uJ�U\���Um��5�U)���f7��v�^֐t-�� �fH���jɩT�\�r�+5�Q4��ڹ	Vgqϕnw����+^(7�Q�n#nfvQ��=��x��-r�/Cs��ݴ�Y�>�X��v�����b��,l�vլ�ι��1�v��N���M�մ�<��@��D *�k��(�:�*v�"հ�Y���a0'3�5�N2VD���2V3��N{*�i^�3�u�kb�8N�*�b�T��v��-�4��j��'l�^4p?-�+�i땶.(EZ6�,�
�!uFꓧ��n�ńբ�b��(.xܱ�A��&�mU���c��k������v	��cm�\��\L=6 N�qN:o[:�^cm�i@%�m̖��SBYh�� l������v�*�]�kUW����'��]"E�ꪢ�:*wQ��UT�^Gn��nўT^�QUmV����*�R��!7S=�sr��*�Z����*�
�j��� *	M
�fP�sf�@:3­�$KV��%�C���_5�S�ʅ�@�!�,�z���%�m�M������݀���Ss�dq�.�s:D��̥ki�������V�*�;e�S2�r��sم^�r�*�{m�M�����>ޞ������j� "o5s�f�0���g n�5UUT����%,J�ܪ�t�VJ�i��ʫW�)V�-���@��	`�Wl�������l���\vh��@`f��	c.e2� b�W\�!���~[T�i %�`��#���H��2�Y�rP����j�{	ZZ����[]犠e3\�&]�NR�x8Y����Ts��;OA�d"#N�'�A�U�F���rA[��S&�Q6��X�mQ�i�-���P�A�:)��X8(�F�b[e��6̀��v�V�En�]��@�Q6�I������yT��^;8v��˸6���j�Ca���X��T�d7�g���uջe�*�-�%.r�⮝N�*6�ih�+�f�8iTY{d�k�(n�`���z���,��<Y@�u�v@9��f*@-P.IB,3�[[M����K�,�xȮ�`��(Éj��U]Q�9{�`뤲���t���5%�2lضZ�z��ڧ��UU��h� �ݮR�ZbۜsfI�������ɒ��"�-�sM[UU��h&�����٭����(�����؄�\��0��ļ�T����55 �T�U�"��{t���`�C��Z��uOy�{[�U��`��W��Zt�5WN��d˹6�-���`�UE���ӡ���6�*�n�{v�EY���*����� �cV��.��q4ue�ZEV8�[�
�kj댵�d�`�h��%Լ���E,J�MA]pmU�	=�UV��Ŭu��VE9��U�{i�p�<;c.��X�]B��,3���!j�TY�n�7���F��`��k�T�*��p�ʽ�����P������Z�M���eW\�v���Θ�qU�֡��F�tj{����� ʻj ٪^U`�-��.(�aKn�;UI����E1+X���Kc�7���UP\���,��V5��/A��� fwTҭF�R���6G���d�2�ij*Q2��<�h�]������{�L)���]K��N�;$�-�N&�3��Ӽb�z8\�md�F8K�f�G����̥,&ګ�:۱r�PlT��b�B�( 0�DXѱ-+׎��g;!�6�5V�낮�j�nڻo]���[��˵�m��D�ۀD�V���24$5UuUU6�%. �+��K�H�(����gtUA�������[<ʵâ�[��uR�UUUUWU��\������K@*�EPU]P
�x�"�;����2.ܣ�(��+*�'D�Uy\lr�V6��)�fiVꪩVڪ�5gs�z�����@��8�9e^��0��E���
*�����U[A�lfb�AUU���F�Z�v���T��P' 5R����ɕKy��U򯙴�U 8�g�V�N�Z�T�`Fv�Y��9)A�՝���!۵k`�j� �N��뭍[ ]�"�����{����s[��*�8@�%����R�Ma�ڷ
��-����p}1�`�̠�	u�����{35(�=T�U��uڴ�	�=�F�k��)vݹi�*:#Z݄D�v猜��Ԫ9M��,�f�F��(�nɉ�B%����t̠� *���kV2� ۥ�C�sn1WZ�P�m�E)Vh�;�R]��*���'�1I�Ͱ'��:R)8�y��/#���L#�e�#(�b*��cn�g���u5NW#��O+妰U�c�*��v����媎��24�zŅ�ų� m���[��l�) �6J��P�4��P��рk*8m�mm�"�M���U]m�E���u�U�Gjv! �.�Keu���jG��$�5UR����P
����8�h@�5��/4k�P6����8@�T8W��(
l3�UUJ�UUM=oh����	j{jn�c`� ֞�N����ev�����V꫶��T8�ڪ���Xeo*B�.�F*�R��]�@�d
�Z����I�wEA¬ UUUUV�N���=�-UU[A�UUUN�v+�� r5UV�QUUl��0ϲ�J�j��ڻL��[$�BY�薭�ռ�-�5�kj���"�Y��5ڗn�l��Y��}����cm�J����(<@Z�W�
`�E��#�<B$ �����"!H
��X!",!+�����!�j���(������"�`+�W�"��!� lX��
z*�>QpAЩ�����N+�i�pP��k�8��"�`����m�&2-���P,j�J�H,dB���D�=�"�@b�����X�p�$	,H!�#D���D��H,���F1UH�D"��=��E8 A�_�p�
��!Uv�� 8�#H���E��b�R	�< �D�O�*�
b&�OD�$", �d C>CB��!�=���)"�qC��5ϕ_y���",``	��{s^'���#�U��z�φ$T���ET4��q�_�F��	�#Q�Q�"
�q0A6��2�"��N %qA1h�N	��GZ�<H� < ���Ԅ Ă2>�@�����pV��,C�� >�>>[�Sh��>"'�-x i�A"�|�x�o�FP�  � ��Z�m�HXH��b
x�
;�	� ��@�� ����x��
| |��.�"@"�BP�Cuj�V#RDGX#}E�8�����(x�N�4�D4��Ҟ��� �~ _�T@��'�"�H�1䄨�إH��m	��F��HZ��$KX���$�d,*�h�H����� B%kU��hY�2	�_DGA BF�	I	B�`�$��X!.�d#Ǉ(�A �Y$�����l�����d��"2"��>4��@\R��A0pZ.���y��u@EW����J(N.�1�@1(`�b��$�Z�Pb�B��0"P,q1*��"$@"LC)��*ңE+�bL fX�6���i
�� aj��S i�h��kRkU@Tv�T��UV�UpqUV�RۜMF�T�*m!sA�U*յW0�$�:-��3���cC��emFQ\��6Z��5)�n��[c\�b���y-n�E��A�-�\���x�km��i��H���-v��Lq�p�g�gx�c�KeWu����S��8�unc&Ս��� [����hV�X4Ƅ&2� �d(� *���&n����nzݍ���B%ҲR[Z6���t��[a��2�y	�б�j�E��P��N*ۨv;%��$An-���7A�/W[Il1�bWE�{U�[��v���<E91���v}S5�6 <)�r*q���:tt%fz�_Z�S��|��x�n�*Nt�ĕkcn�:Ժ:�`)213u
�q��X�I��w.���Be}nd���z�㮎#!��l6�����\�F�bǛ��[��<''V��t�S��ruF�W\dx��h�q�sI�m5p�)��lHM�542�]Y�@�5c��˂GZe;��pz;k-"�E�Q,&=m&շ\�=K�;��q�c5r��!��1�������3��C�`mm�<T�䢝��6�Y�Q�P��,��,�Aɤ'���&KQ�UVN����<;[[���eJWT�T��Y�*���m:���;�1�[@H�v�1�*�)7"�9m�˱��6�5��a����fJƤܖ��[���Ewc�e�3��d�E�� ���F�a33i��ׂy��s����n�<��[P����\��T�9�IGɲb��7d�	s����8ٷ<f����cUy��j\ĺ�3�e�V�$)UIH�d�XƮ�65ۗf�n�4V�JViT�V��Z�k*��D�����ϝ)�[.��:Qܴ��]EձӢXH��v\5�d�:A�ֻ<�ʦ[���vz[�N�ǚ;Vlj��6;;Ɛ��v����`�2�u%e�I�2�nk�qs�k�9-��0��Kf�r%��C����ؕ&�2�����!�̭B�r�gK�]h����N�N���Q�~EtVm��*h�� ��M����� �g��T�M��]���~�*	��6�"m�q��Ƭ�r�f�\��\��ܱ�<Ҝ�JV�Ս֧X�u�1%�rY�����J��L���4�t��.r�y�V�ق��hUm.���\�}�G���ks���(�I2ƅֹ&�enl%�;g	�ѓn�F2V���Y:H��+�����I���ˆ0�X\�[�"���ٚ�R���We�����$�{�s����N�1f����e�vx3�S�n;��CM��ڟة��ـ}��s,?#��q�XZ��)�H�IR�UM��N5y�H^�h��:���������i�%x���`�u`x���N5`6N8��j����`��� ��n����k�m�`�5�=XYlu�p�X�Ƭ�;E�w�y�}�-O���v	V�UI-�R��m�RVS<X֬<��)�5#+�TҶ�YP-��U]�Vc�Հw1Հcn���S ��XIf�mz�O-�L�H�".AQ�#����ڰmՁ�1́׎�TF�ԪJ� >�ۀ�ۇ�qri�������(�Hs
fjB�����m��CX�l����%��������	��p�vۀy��0�I� ��V���7����w#h{ �ַ<�;�%�� ����=�v�º��xl�:9c�A��@V�Ý����:�Հcn�^�6P{!�d��� �}� ��ـy����W�����5(؊�R�S\r�_�ߦ��lé$��.p]�IB("� ��6�i���X�q w�k�_���=�[�x|g���%V����f��l�=�^ }�ۀy���7��PqL����`����t���u`c�Ձ����}�&,�H��|�Glh�X(2�N͙����6̂ũ�It��݊�ф	�����V׎�rڰ1{���V�5�u:
�Ue� ��ן���ǳ`7��X^:�<� Uĥ*RT�US`b�9�3&��q#����~�0u�P�Q�hӎ�0�I� ��V&��v#j�'��9�3&�������l��(� �qՁ��6/c�1�j��qn�m�jD�L�ta�[mR�к�ݟ~���_��w�F�ړ��3����	Y@�b�Z�1�����1{���_Ds���v�/�o�a*�Rm�0��f�mMX^:�16��q!��N&��T)�&jl�I� ��VlDBOguX�����Y���lt������s�{^Հ�wU������t��1��1�8UJ��ۀ{f��?.l����}�u{w$��ߵ�'���C�8<�Ud(A��<�2L��Z�M2��vjێptq\]��;'R�y��j�v*���b=�R"ݨhkFfX�t,�}���6��M�Π�iwh[:ݺŎ�&
p�m��(��nل9Ѹ��;�[��p�!���*�<�(
�eT��G�nw@�[n�!l���h��s�,˫��A#��Wicr��S�ڱ�sLWm�)�`n�C�M�a��齍h���5m�c�wN�z��z8�+in:Ġ���.]�x��s;��N]���p]^٫���p��k�=�� ���x��n훯 �Q�����8���t�������������P9��������ͻ������t���I(�J��P�L�U��"��Ł�́��5`wv�Z���ꎫ�+-� ��9�<�+ �;�y�r79�ް].���6��(�]����D[��n3 q��a���u�k����o"Xd�����V�7V�w��r9A�́�z��T��U �������?HO�Q>�M2 f�4�t04��0�P�Q=�y�=ٹ'w��5��L۴�M��*�U[j���,/c��c&�;����uT�W���;eX���O���`��6 �X1�X�JY:��D�*jl���V���;��c�k��� �{ɡ�Y�ۉ��M���3k���@�5�,�ez��R�I�%�{��/"(�F�& w}� �{q`����I�}�M��j�b"N6�����#�^́��`�u`w�9,B��X'YmX��ـkﴘ$�ĳ��%���ǼI"s.��������<�#��V;f���`����;��1́�m &� (���TM�w1Հ�Ł՘�$��c'� ����<�JTbl�5�9�d�l��B�!4�	��D�&0A��un
�^%��a�>P��}�� }�� ���n���{�| =������J�\.g���u| ;�}۽� ���� ��}���[��z�ں���� ��=�I/7tZI'���I%��ZI"w�e���mE���w�7�-��~��[m�����m<��XD"��B1"�E����.s��K�[o���e�����*j�I$�c�I-�D�n�u$��=�6���)����|��,cu�/�^����kaf���@�`!�T�閷;(��<v���h���T��߀���� ���.�$�c�-$��}��$����tpN*:�-��o{}����$�$o~�ZI-o{�I%��ZI.�iA'JPEU ���RIcwE����c�I$��� ��ݧ��_���b;k6ct�5TZI,m�;ԒI㪴�Y/7�$�{�|��{փ�ĵq]g��Tۚ��Y/7ԒM���Ico�ޤ��_��
Z@�FX$bB �#�I9�	#�6�D�kDn��f鳦f���%�
����jI�[-�9��e�M�١(���[!��&��]YHˊ��l���ƥ%�T���6�M<�ئ�gr<k#�c�u�۬.����%����y��Л�@]�>3��
�v��;�\%#�m˓��j�N�˲REa"ޤ[�Ħh� �ՃUr�f���;u��9c����͘6��L����zI;�4o�k)v(�&*��ƍ��f!iõ�ձ��n�7Y��Uh0����6�ͭ��X����߿��{�(��X��w�$'�j�I,<�U2*Ќ�aɽ� �{�| >�{��� �z� o����>�����l�9o���}�� �W����7���|o���v�Q���4���}$۪��Y>mOz�I�qV�|�˖���{){<��FW9� �~�Mޤ��w{�!=��w�$&�դ�rY�[�K)��S8��#JЪt��^�qs۳��@�$��Y�H�SA�&ҕ��5�P*iOz�Cn�$�6��I	�5���w}��o} >��&#������ݶ�~����R#� F�VC��`
y�֬�}��������= ;�|o������#�P���ޤ�OU����j{Ԓ^�tZI,m�=���wR��ʥ+����v;Ԓ^�tZI,m�;ԒK��$�K�v�v���nl��} ?w�7��Ɵc�I$�U���6��Io#kt���^ K{�,+5
r��ڻXB�`�uj�26ޘR���Z�h�a]�hV#2��)��	'����$��uV�K<��w�$���h߾�u�F%���Y��z�lG"&e'���ޤ�{�E��e��D�|^�S�ʜ�Ѡ�U� ;������~�z�������l��{����(����� ��rl�$l�y0�0���$�2$�]�Ky�9�b�A�gi�.�����=#���_o��<Y)�d��<��5F�!#���R�&!�����@����!��\��!��}�`,0<�8l8xr$�A��X�ǳ &0#$�	�ddr�L��~G�O!}�&�ާ�n�=�)=u�`�� ��*R�<��PL�ȱx:�O��!�7�s).V"!� ��]���Y!A��.�*@b�B��N%Ϸ�/����L�<y
a�rg4xo9<��p��ơ�!g0�1���q{�����9J��AOD�ĳ��Ls8xO!�����gc�
0�7��;�|��f���72���DՅA"��4k$9&�<��t�S}O� K�.��1HBy�Fkd�K|���i�<w��t��h�-O�BO�9�`<�����m8#�|�!���j���HF��.�r0�0��S�P�����|�������5��Dd�`D�R$L����EO� ��S��|PJ��`)�s;>�>�z�If:�I$�{0EDUF���}� �{�| >�{��� �zդ���s���y���I!��f)H
����[��{�g��{�� >�ޏ9m��ަ�����L�\&w��ݵ����kX�%����g8"!�]�^�!��-9h-�t�
�+?~ ����| �ڮ�$�n��DGfROw{�I4.B���)B�\� ����@��7�����} �{����9?rK�A��@���ф0���@�����{�g��S��| ~�s����;<�v�� w��{� w���5�[q<<����TmZ��5%!���g~�ݶ�=��3F�fh�0��Z9�m�;�s\���⋯���$��ۢ�I{2��$�����Mr�Q��d�*��\і[��x�q��X�Y�)X�� �����+)E��	\�� ����ޤ��wE����c�I!f9�I$�[���E�u��}� ���� ���;Ԓc���K�nk�ؙ�f�rL�(��@��-�6���n���޶��K� ��{�} ?w�7���z�c�ҕ��Y����� ��{�= ���#�����J-��f�L���ĒK�mWz�[Ȉ�{�:$�{���s��o��w3v�z�rDK�A&�:�~}]�`���IPp�d�,��\����rkh�;;�0`����1h��&�ZJ&�{C�4]p�7� �s���T�y޸4�h�=JAvZb-Ҙ��¦�$���K)0=��j�7=6L��8s��v��B��,u�&�z�g�SR.^�75��h
�9wN"��:۫i±]���h�رW 2�!X�W�c6�.3X4�4+f���,L�~��f���+�aU����!-�\��/���1�P���t��(V��s)�:��2\.����#����������@?��� ~�ޏ��wꔇg��d#D�����g��?�� ���= ����{���登1,���;Ԓ�jm$���Uޤ��;���^��=���JQ�Nhh�h.� ��uWz�G��U���7��RK�8�m$�6�k�2f`tʏ��|�< ?�Ϟ��I,S��Ē]�9��$�F*��\g���u��A]g�"�8���N�(���6�P��Ȥ���g�Bӗ��
�=r������z�IcuV�I{��lG#������< ?|�2�y���\"�} �۲���%Ĺ�{��~����m��o}�����K�RG�!�QI�mJ��SV�I{^�w�$�7UiL̼o�ޤ�}�������F�va;9��?&e��ZI-{���$�ۚ���f}�f��ݸ�?����#D�+�����ޤ��)�ٮ��^ǳ]�I$ۚ��_rs�߾����))^6C4!�h^N������99�Г9��Q�:5>Γ'���A��(���y������m�����ձ�Du=ۋ�p!n�.L)��UUX}�j�9�$n����Xm���l���4�t�9j�ح�\�����O~�훘�&� {IXDA��p*l��� /Pu�������p{Ʃ&&ʣ���R��r!=��Y�G���`7UX}�!n�ߞ�OߪW�J8B�� 7۶���Ds�:��W��g����dVƶ|fїi��YKHT6LX�%�eö!a���T�#)rDY���}�v��b�jکU5^ ����X۸�r"9�������?ȶ���vK.�����#����7ﾸ����;��^�	��Fj�i��:�`�~�� n��s�KۻtX�vl����4UQH���UTXls�n�Ձ��uX6�rq�"�\�H� �b�	���T�Z����}gH[�ܜ�S%H���;�RՁ�;�=ۻq`�V�Ȏn��OC�$H)&E-.��jDnz��&�M��[sk<q-Z%�{]!��:N0�}�˯$6D��o�����:۸�ۭ�r#�<�N�6&f����D�`n�,�\��K����}Vn����~�F�9ȉ�SݨJU䒎��Հ�~�p��5�����Is�O��������� ��6�Ȝ52������r8���U��wU���œ���QL����[�{{zY�e-�G)l� �M׀$��9�/������~����g�rJ� Hȉ	 ��>-��ձ7]E$	jv��qQe,jË�Z��n֐�F�ˠB:Ǎm�Gq�.z&�3��1�!�Kp�pu$osqf�5/�XF��:u�u��Q�8��sk-�t��A�m8���q�w�Ů�sQ�x){��BX[L�c��Va�2�&2�� k+���fۮ�%Cv����pZ�����ӈ�@Gc�������xn�&�Y�\��ղN���NCK=(�����+sM��R�����x����k�S[��<�c*O�wN���k喷%uQ���~���ŀ�ۀ}�Yky�Dr:�\�Vn�n�5H�)10*�� ~n���9�9�3v��`}��+��ş�Iq6y��_�ȜTm�<�N��Ƭ؈�B^�ۋ �{V���X�(�b��c���$���%>���`|�����V�Dr���1����X��T�-��w�%ķ^�@���VO�s�8�%)A�r`M�.��ypy훳b��L�'.��żPl�'t�2�=���I������ڰ:���w��s�77n,Ɂ7��E�2�q�n���y�C�7�H�<�a������JD�!�E�@�b�HD�F	)��PX��1.`U��I���1��,Íԁ�T"��D*̤��(TB���@ Z�5@*!���2n����}��ܒ}��k}TBو���T�P�MSJ���f�~n�ϣ�s���>߾�#���Il,�Tq�,������������vS,7���-��l���D��&��	UTX�u`}ȎG��d}���l���wۋ ���=����q��R�Y���vITZkca���"ʜ[��jVV	O��IBn��"qPt%��?����g���=V{��ȎGP��`k�P��2�v��0����\�\\�����`��\ �o���M���92(�UGk�7�� ownB�\��#2F���
bE�k� 2XET�Ȅ�����������5��e%%!bvՁ�(�8���X�^Հ�76Ȉ�ǽ������cv[�.���r"6[���n,'�l��B���,���&�5��P�Q�ѧ�x���kn7P���T�1I�N�:{��}1�ms4�b����=�=����x�y�G:��n���f����U*$rK0wۋ:"���߻��O��nI��߳}F����~ʡ]R��M�V��L �o����@? ���f����nI�=���5(�Tm�0?.s��7��߮��w7$��~ٹ�����"�yL�=dSC��,�E"D#	���@4B�pP��� ������ߚk"�,Q�J�� ��5`}���G߽�}6�x����	�J��MSGbe�t��*��9�XP7;<����)��M�f�B/|�:v���Hbf�&*%M.���Ł�ۛ �<u��K��<��ߨ8��JJB����x����"9�	�{V�z��n,����������r��$�`c^Ձ���͈��$��Ł�f��jyTlu4��p?��K���w���7~����x���G#�Ds��q��U��~�??��*,rK0{w��?���z�~�� ����p>�fI%���_�Q�)�+fF0�[e>��Jͮ>j�0�N�vc���$ �)o�P�!D������a%ٴ�4T��	>�ܰ���#�BsZ><�V�%�am���B�}@�^sҶ�T�8s��"�a=�p�p��m���#m����֑���̆�j�{��2։1.���A�K�ĉdHi7�Ɉ`N[���5 H��X�8c�ջ`�CSf�kA��"E5��tHf�Y!B1)�$���B�x:�0~߁��̌�L�﭂���ɏ6����]�(wY�[�M��rc#-�xp�����v�PPe��Ub�����f���T&5M���u�Ur�[T�U�Q���V]l�A�[=�O:7n�R���
���Ȩ��c� <���5x�
�'����P��7])�rd⣞gK�=8�A��ˮ�nzt�c���J��]��X�̖�҃vqKtі:�`�-܁�j�l���в�KmVYk����zs�mJ̨�&��v�����[\T��4y�]j0�n���#��[9;@��]d�0-��0m+4��]J
�.��"���[�/��#���t�[{GSs��;�bJJ�[̈́�iv�2�{�R��}/g]��ɷ����@ǘ�e�u�YfpY���dۀ�2���{&�̦�C$/��:b[�+Y�qm�W2hJ�ҌU}n؇�C�c��'���6�Np�vN)ᗞ.{=�l<�FC�D�]{63�F�$۲[] !b�
��g����m�]�>���c}�U��fD��.؋q`
�ٌK�2bF Ny͘\C��{6�SӴ� bsIWKl�\\���2.pt�sє�Lb�[vM��q�77�WH`�m�m�1��/ob�2h&S���\l(�,��ڭ����L�oR޳c�ݸm^��n]�d3u�Qc��s���LYն��k\�"���[r]B�Q��v+�����p�R�%"��d�X6���&��>�-\I͠t+�p	�s/7����	0��A�j��񹶆���FU��2�ia�J��v��|:cV��#��qBt�Hs�c�W��A�2��X�3#ȣ�Ҫ�Z��,�'kk�9ؓ��x	��px���Y��t�-ó���m&����ip�Z�ufHkt�Q,��=:���1�ץ�l(���nvK���fbW��}[�J�Gn��,�l@NM�rlnn��G�dr�3�X�X�G��[[F{L�Ef��+���.|�'cf�I]eu�bzY�r6�ղҲ<AVŞ��ݞY;FQ��u���ͫE���̆�֡K��_�4;��M(��!��U�@nH����P� �+�>���`����"8+�P />�.�,�5�j�ܤ�:����e%�hz9Ė�qn7K�-�Q]�9��5ۃp[�r�@�	�m͓oft*���z-жf��/n-�u�3�ݵ�M��0\M&�	Բ�c:E�ͥ� ��te����^�O��؂���pn��ke=��r�,��ם���rQv�T]�.�H!ى�yz�v�q��Y0�!�V��i�5��(�9�(�E��Û�0֭�rj�c`~�k�<4l,��\sb`�ŵ�,f�[��F��J�I'��ʙ]R�� 9m_��߿������w��un�Ł�0I5?%����f��3�K��I.H~{�M�������r9H�z�E�&(c�m�U,��\}������9'������������!�E��������s��Z�{�=�����c���������ߕr��RRW)eXW�́���6\n�@<�Հ�}�;z��5t�b��GHֈ6�@�kZi��4�]=�)k��ޱ�$��m��i洤T���O@2�XsX��>�>��qv���� �~�_�%R1�ӎ�m�$����#$$
H�`�MQ�� $Ta"1�a�@`DdiB�@H$"`� ("�AnO~�vX=ٰF7W�}�Ds�'��(ߥD��TY����������9�q&�-����\wtYX��ұ8�-�a�Ȏ/Kݛ �{�`yf9�؈������/ɷ�~J'[v� ������9Ȉ�og�cݸ�:���'"u�k{�.3�S@���l�����6�]��h�m,�$a����'N�:i}D��bRTTL�x&�lcwV7?G#�_�%������� ��?�!�DG@�JSS`{���s��!#��̀d=ڰ:�����ĒR����U��II\���{�?~��O~�[�(�x���r#�mv�l���,�|R������?(��\ώ����;{�ٹ'���,�ˋ��߳�@�7�������i�P�����*�9�G���@��=�p{tDiFr&�e�@���Ce����`�4���z�6̺d�1�����/���%d���#�߀���� �f���n���9�oj���!Z�UJ�
�0T�TXrڽ�9�D$v���`{ş��gX�&ޯ��NPu�,�Cݫ �c�6"9Ȅ���XM����M=��*�l��߽:}�N������������`%�T�BA�R�1	XI��EOȣo�Ͽ����C$M�J�#���w܈��}Ȉ�en�> q�}VVc�-������(�)I�`�I�V�Z�8]�v�ƛ��j��R�1���Iݡ�z8mŵ:J�,��:�L ����>~���q/�{~ŀy���"�JJ��l�F7W�s�G""dŻ��~�����ٟ����sW�/�J�C��Nۀu�ٰ=��Y��%��̀d=ڰa*�R�ei�H�������:�L �cua��%���װ�+�SSH�Q[V���`�\\K���W�����~����� \J��8�����r��4��wN4�@y4IB�h�M�9�rOFo;�Wg6Ѵ�k�K
1me���]u!m������2.�״xlBs1Qz+n�j���<�-�$mX笖���.Q�Jh�G�Y��<��ߑ?��|K�A���u���5���m��2F�U+��RX���3kI]Sz��.�j�K4)YX[r֭�kkx��@�X�n��N���;��g�=�r=Rⶶ�ˢGFVm����KM�����ұŔ0�/9���s��bmՉ5b���,����� ;����n�� �G��y�~�~ߔ(��E�6�T������f��ذ�ڰCn��s��l��I�LMB**R���ۋ �c�7�����`y~�� =����VYF�u[*��ēoՀdn�XO�o#����X���"��u���V���.$�����=��\X{X�P� �(#p�'q�#���Ge}���sW	����\��ej`������v-���_�i�{V��� �c��s��ݫ�$k
J����9-�=��X��G8��"=�s���"�w�`�V׎���>�����k��u&*+=m�?~}� �cuf�#�׵`7�q`w�%,��"qT:"Kp?.$������:�o�f7qa��$��X�T(���"�&TTL�XO���X{X���m�ӽ� Z���8�+�	�l�nf�<K-I��֛<��C��j����{f�D�R�Ucrπ��� {�ۀ[�q.q|ï��������!\�t��U5��W�����q��V/��3۸��9�q��6
)��W��n zw��rN_��7*��H��$6��c"H����U�=E����f���$���e�Qd%M8�r��\}����;��\X{X}�s�r"e���XA�UU���	%�}�� �����z��ڰ:�9�>���(Io�T��;��n;=�9�\;rY������ͷE���^2�Ym���e�|��� :�]XO��u=ۋ�ؔ�lQ �*D5V����#�Z�l{���ns�\_�\������YIA2�t�������6<wo9	Հ8׵�w��1H��TʬnY���=���V ��XC�VʎG=��"�7�3�� w���k��E]�U���C�VS�6<w܎DG�
|��P�����k;�Ү�y��mƥ�H��!4�HÒ"Ͻ�e��`{V�8+� ��~���;��:�x�����g�)*i�U��=���ě7��ŀ<{V�nj���9�92liO�r���TL$����� �c�7�Hy�.��L���f^[m���l�`lq'�j���XO���X�o�U�*�r� ��e�?.v~�Ӡ<ݸ��:�/��e<�"fp��"�m�*&)��#�a��f�+m��%c�L�C]��]��a�L��7hT]��N���1�	�dD�!�FmJ��=4֛B�� �f��������YLR$�e���r����ջr덡�#��I�wf�aq���5
QB��phYne�d�K�7���f/���~j�� [�3M��&��.��n�8W1��L5�����
 ��s���>I;��������P(�ml��O���孲�c0��� Z.��qӧHK��a�O.f��6�Q��������,=��#��f��-���&&EP��E56y���q x����.��l��q.6��[$+�WF;j���=� �c���D%�f��{q�u���$�)+�vU��.q������׳`{��,>�9����N���`n��n?悰��,�Yp��f��s��{�ۋ �c��>�pC��X��[�;f�v�PbkZho��z����4d�Mpc7L���f���BP�'�����論�c���s_���:��7f���F^[e����j�;�n,9��_�ĹV�ܮ+n¬��(zVLVl��fB��$�9�搒A�
5�H,J�2��0�����g�p��5�'׿~��<�n,��ě;��=���7I%� n�X^nl���G܈��׿\X������[cCv�ۥ�ˀ|��{Ł��qa���٫3M���PLJU�$SS`g��X�{��ǳp��� �v�z*�mF�iG�uR���R��y�أom1���mh�lFf�� �3+l�E]�U���� =�l�Vc��>��H7��F�y?M
&J�S)T�Xf9��1́�7q`w1�_�I.H~���9�p�U:J�\����{��Xb�>X��椟'D>��6Bd.��a�K/j���A�/\�8RZK� \)��if9����Vl��F�pٱ�9BB�	��T� y7�`XCV�d]��,��%,`Y7M����� A	�(O<�K8z���^	���>>/�"FB�B���a%s[��l8�+�&e����4��,%(jkFY��aᚪ�Y/�� B�iK�a��dE�q�������h@��d�b-(̚`��J��.�&Y�XB���d�F�L4��i7���t�P�jB�{]�& R�]����ev��MS�=�r{�u�k�����M���a�ލ��ˁ$!�>#�k/�R��k8Ȉ����h��`
M�K��7H����W@����&*���hO��D�( �ꞈ�"���x��� ��C��z�����;1 8��Q�k�o͛�O{�s[�|{!3��j���$�����,���`}�.���`{�yx��m� �c��5cݚ�M���q'�n,�v�^�u���j�Y{)���У��(8,�.�lF�խf�uefs���oC�]�*���y����@�of�ǎ�b9ΰ���X���i�m ��.՘��ǎ���c��csW�Ff�/DR:�U��0���`{ۋ�}2=����`ub���D���BEUTXj�{ذof���6�9� 0`��`"����䜤��f�5aer7eX�{e�?s�w��׷sŁ�#���P!Ẻll�6}���nbJ����>M�v��x�]O�g1e-m
�I\���<�~��^S,�;���1���6A/�UQ3J&$���yL�;��,��ՁՍ��G���⪚�T)T�`c{q`m�Y���ݛu֖��VD�7��.%������p?߿�������w��R�[j%��:��s���:�ۋ �nj��rߚS����8o�H�S��ŗ���G8��M9V��u�7q�rlƝ�$93rn�Ct`62��kw:�j�e�����9|���Y��sv�g�� ���5�7$��)bFY���c�&%����Z��:�q��g��ԋYq�yհr�5�c���\�z5�U֦0sp��B�����=GSRij�YV���F4�-���'������۰a�:���'����'u����;�lG��l�6Zȭ�X҅ Z܃�{���^����)�X�����~�����>�� w۲�?{f��O�X�H��V�`�w�H1��Xr�X�{�q#\�����5!h�vU��ߥ�>���?9G9ɝ�k�����Ł�:J	g
�*t��l��{^��� �������7�����
?��+,�ctrW�y�2���ssw��of���X?H:�-[d,��Y�O8(^#�v:܇hD���t�[�j�f$4e�f�s1r������5`<�k��G:�5֖y�G���F��d�`}�"�3��ťvQk�C �C�S�C���p��V�u����ŀg�BN����PJ��\}=� �����I��~ŀ��.��L�n(J��7)Xz7���zP����49	�cx_���a$U���e0��, �nj�y8Հ�S,��:E"&f4��α�ve����#Y�GYbj�V���ZL%��������f9�Y�m�ߛ�V�Ƭ�A��q`f�B	�EB��W����o���w w۲��%�پ�~����7G-x����7۸�kB�.!<�]`���u�滻�nI�����<���y,�A�%�S �n��䶬7��q=����lJro	LP)*f�,�ӫy��W@{�����ŀ{�jDO��#��uT��۠+[��'#u�n2hFb�"Fl�\kk��PZ�%��n���L}���$����`����������`�$�*IJ�Xn�{�G8��v��1���9��?~x�Og�\b��Ki�{1�X��V}�r!/9�V{ZX�4oxZ����ܕ`~�M�~���}��ܓ�~��rO`)>���׋�ٿ,�[	�
(��+-�;�ڰ7�������X��Vq��MƼMe����!SA����&ٮ�1nJk���K�
�f�'I��=ܸBT)�] {�V�ŀd6��s��#�����?n���K%PuH����w��}2}�X����1�W�D�\����z~n��jK��֍�'N��Vr[V��X�;� ��ē1S*e)�
�����Փ��`��`{��Xqqq)?/��� ����&Q���T,j��=�Ձ�9����dn�X^nw$��N'�����.X����*�1@�!���\�.��I�8	j�F�f���j�V�7n2ngU����qs��v�m�^l�����8NgIc[]u���ơ�dʚ�1��#��S]��e��dv��׋�n�@Q��n�����v�d�vc�g���SZ�+�0v��#l�i��n�X��,�n�w2�]$�]K��,J,�[i�a��9�i-Kip���8�/�;Z�:�Z5�պ��Ҕ��d��Ѭ,��Q��J6�a)!��9ݒ'
��e��ں���2{:H�휂�-��~�Xa���̀g�Ձ��`�����##�U�-���8���ߦ o���;��Y���G�#�
�N�W���vl3X�w�mՀ����NW �r[0�����ŀ-ݸˏ�߿L��~��y,�A�"�5V��ŀvu`{�ڰ�u`~��i��+es��nf�U1/V�q�Cˎݞ8/e\DIS�a�5��=���vn�m�)�����X���َ��9�}����X��)$+�:��l� �g�]��Q�~= �'5'��5�'�n��;���F��4*JaQ%HJ�V��X�w}�${^Ձ�;���鬤E�������, �qՁ�Kj��I�ڰ<�`NuEEUEJ�MUU�u��G#2�W@=� �wn�z��
�6Xr:�&���Z��ԝ��V�xg;��\���h���{��쁑���Pr��������p�ݸ���tQ��P���� 3����ڰ�ڰ=�m^����x�%����]� =�߮ wwn�j_cU�1�da$��"� ��*�dB$��X�!24x�[ιޫ כV��)d8T��(��j�>�BY��`f���3��z��w�m��M�ۈ-U�po���{���j�<۫29��	J�iZ�]��*4KGvޝ�(��b#.Q
�kd��̒�%-$��� n��V ���ͺ���`u�KE%���]�� ��nq/�.)\�_� ;�m�>Z�6kQ[U�A�쪰���~�e�G9�#��7w�>{�� ��dlEi����~�\�ޖ �ڰ����Dr2 �p� �9��X�V>H�b��&ߗ��d����4���RA��Xf:�>�D}��G�� Ͼ�����A�3x0d����;%Q����6�ͱb���.`
��5ZŖ9��4��Xׄ[
���5V��ŀu�V�-���s���psToW��c����Հ�DBFd� �{V�����BA究�X�(�Aj�[�{��� ;�ۇ܈��n�X�ڰn��D�Q%HR�V玬�w�n�7��m�� ����B�-���%�`o����X�X����'8A���S$!��&��4B���d��?E#BFK��H�z%4d������`ptz�#	�y)�$����"kABHH� bJy���lL�m��8�1D��	 ��(SZp�`���+�c��4�VV�'���zf�3��0�H|����oN�ҩ�Ɂ ň�-��r�sϧ���e�w�
�
���U�R
���� *��p䊂�T9�.�Vθ��Z��V�tv��V�|�-��qHi��eJ��yͺѸ�I1�trN39�Y.��%�۰���@q64��PlV%�ʦ�����(�m�⑃�X�mK�lK�[@K`cYh�`���N�܂�H�8���=,j�jJ��T���x���'-q�H��g����[v��9���֭���ۍ��Yv�XYu%b�P1�bG��qd)�.�{�[`5�`J��CY#.q3rQ6��t	��Yלs�pq*�F0�J�l,.@m�:XJ�q��}� �x�Ĉ�۱�'�屳<�e��X�	ci�$� |j�Q�SEʌ��mKSE���Q�9�b5k�kVԲ���ˍ�5-���X�s�UNX�gB&0��<���U���O[����W<a�_
j��X�d@�v<�pL,��cuH<��T�1�B�$�ـF�6�u�	l&�SXH�y��ݎ�t�9G�8��\�=��ŵ<JM��qq��n@�������8�i�7/mpvg¡Cx�����睉|#�Q���Ru�<*�x�ۙMm�^�z�+n d:N�t��+FP�*43,��t�����4�n4v	8�c�D��[*�&��3PS�����������݇ԛ�x���\۠��N^�6�y��s��+�w`5�qٽ
�,j�.9�ۭ¯;t�ݻr�����ɛq�z7�C�x�QP��L�W���k�6f���+�7��ǫG;{�qHd9��P�J�v��7k��������Z�6g������@�G`�$�Y[2R�	�/m-M54Zq�uڍu���DM,dr�kͮH5pU�����cfpr&�F���nۛn\Fۖ	�wUS��l���l�n�!]6z��;sn��q���m�ۙ�nQ��#��;2]a 9�g=&��a�v'lF��R���\�ҝ�p'6��J��Ս��l�\v�a�\鲷`Έ���Mp�B���ece�-�)�`e&D��$�{��0
��)ꋈi���@*� �E�� �	�GB��|(��4�h�%@�]��J
bUS�S�/�k5d��M�<`pa]Ӟ��c\�A��g�n���q��\V��-�,�c �s\]�i�Tⱺ�+L�l2�sK��"���g<�b3��x� s���nʆx�[Cʘ�nK4�:�l�eI����\GX�7+��������J�K�϶�7<�s�4�ֶR2�Z�z�ؼIhN�\�)m3�ᵛ����MZ[sRd�kF�|��G2$�0����Z6��qu{v.ݞSX��L�kgE2�M��$L��q==�����0���ڰ3�L�1cs�G9G9��}���?�H&����E(�nY�{��`^�6��W���#�s��3�$/��SB�E*���i��`y�2���s ｸ����ay,�EVB�0?.r!y��`yf���wȈ���f��z�jޝ.��Irj�56��bX�'��{�ND�,K߾��"X�%��{�siȖ%�by��iȖ%�N/n��O�P����E(ө�!*�pV���c�[��)�h�A�1k)��$�ŀA�u-�&�fkY��Kı>����r%�bX��w6��bX�'���6�g�2%�b{�~��ND�,K߿~��	�P�n�g�8���/Oo��4��B�Q"�X��Dh�,O6�!�6dL�b{��iȖ%�b}�}��r%�bX�����9ı,N���n]Mc%�DWd�����g8���~��q|p�,K���ͧ"X�X�'�뽻ND�,K����ӑ,K��ng�0X�d�7�?/Mzk��^�����"X�%���nӑ,K��=����K�����iȖ%�bw���VТ�R�,�/�&q3��^��۴�KİD�=����Kı=����r%�bX�g��m9ı,g~�@��7�����XѨ�v��i�5����;n�"L+s��	k�#
c����ֵv��bX�'���ͧ"X�%���fӑ,K��=�sa�Q(y"X�'�k���Kı>����h��]���g�8���/{�~3���ș��>���r%�bX���߳iȖ%�by����r%�bu��_���*�L���g8���ﻛND�,K��{�ND��q8p"�'�Q`���&g��m9ı,O>��6��bX�%��$���R�$֬��m9ı�<�����Kı<�~�m9ı,O��}�ND�,�"{���6��bX�'���o�Fm�*V�{���MzkǙ��ͧ"X�%���}�ͧ"X�%��{�siȖ%�by��siȖ%��.����਄"�9$�l$���]�m�x2��G[�+�FYy{'�M�m���i歘I�e��m9ı,O��}�ND�,K����ӑ,K��;���D�,K��{��"X�%�禋ܹ�S5�Y����jm9ı,OsﻛNC�E"dK����m9ı,K�~�ӑ,K���ٴ�Kı;���2N�a�:�eֳiȖ%�by��۴�Kı/�w��r%��b{����r%�bX���w6��bX�'���~Ϛ�e��t��5��'I�=����r%�bX��w�m9ı,K��w[ND�,ü�~��)C Ȓ#�`P��g"8&U�;���P��tF�?��~�}�NFk�^�����οyf��j������bX�'�}�ͧ"X�%��}�siȖ%�by��siȖ%�b_;��iȅ�/!yO����!��Z��N�͸��`��.���TΖ�\�kYpX�39ǻ����bem�A»)�_L�g8�n�ͧ"X�%��w�ͧ"X�%�|�{��"X��;����r%�bX���v�`�f��D����zk�^���;��r%�b_;��iȖ%�b}����r%�bX�g{��r%�bX�ϟ/���0�Z���5�����r%�bX�}��6��b#bX�g{��r%�bX�g{��r%�b����gM�i�����/!xX�}��6��bX�'���6��bX�'���6��bX�X�����r%��Mz?��Ꮞ��m(��?/Mx�,N����Kı<�����Kı/{��iȖ%�b}����r%�צ�,����|��7E&�kH2[5�B���׫[M
X8m�`\G,���gGD� Ҭ&1�#���t3��X1Y��0e[���������h;;]�'�`M� WR��+KJM��
������@�kT[x�,��;v�lpe�ܚ�L#��Ɨ�� ��k��j��U��;���\O[�k����֝\	��2�.�ˣ�q�X�١r�#�H���eK����#�w'wFx��o�q^V���Oa�]�[I,�'c����79���/��1q�;u�9-V{���צ�5�����r%�bX���u��Kı>���l?*�P�&D�,O߿~��K�L�������p��v�.q|q3�ı/{��iȖ%�b}����r%�bX�����r%�bX�w��iȟ��z��7�߽~��QP�!��O��D�,N����ND�,K�߻�ND��ű<���n	"���ڒ	"|�I�����.e�&��
����ͧ"X�%��~�6��<��,K�����r%�bX����6��bX�%����u-�&kWY��r%�bX�w��iȖ%�b��~�bX�'���ͧ"X�%���{�ND�,K�}l�/�\�M*�֢ ,� ej����̆�C+lX��6��[Ti��F��Mm9ı,K����r%�bX�{���r%�bX�����ND�,K���|������������8X�lM���"X�%�����!��1�D�	uE���6؜�bfw}ͧ"X�%��w�ͧ"X�%�{��[ND� �\��,O~ԗ�_٧0ֲ����iȖ%�b_߿~�ӑ,K��;�siȖ%�b^���ӑ,K��~��"X�%��f��m����-�ֶ��bY��dO���ٴ�Kı/�߿kiȖ%�bw�w�ӑ,KĽ�{��"X�%���jO�hP˗y���/!y�w[ND�?eL�P�����6��bX�%����m9ı,N�~�m9ıL�k��6(�~��C�����e�l�
���anنr��K"�fr6fJV[*uyf���k��q<�bX�'����iȖ%�b^���ӑ,K��u�n�yı,K����r%�bX�zj߻-5m�R\�Y�ND�,K�����L�b~����"X�%�~��[�<��,K��߸m9� "X��ߒc�5v̵U_t��5�Mz}����"X�%�{��[ND���	�҃H� ��)# ā$$8�U�Z"b>Q|=��9�?p�r%�bX�߾����8���/������uUe�8r%�b#b^���ӑ,K�����ӑ,KĽ�{��"X���~�'�~^��צ�?~����nvYs5��"X�%�����"X�%���{�iȖ%�b{���ӑ,KĽ�{��"X�%�{�Ӳ��[l�0�������srU���lС�M��\k�@̖%&���&����zk�^��{���r%�bX�����Kı/{��j�%�bX�}���r%�bX��k��-:j��d�֍�"X�%��{�NCՎDȖ%�w�m9ı,O��xm9ı,N�����/!y>�[S�#B�M��'����%�{��[ND�,K��ND�,K��xm9ı,O{���r%��Mzo��%�������4�>����Kı;���ӑ,K�����"X�ʦ�	 "�D��� lGr&�}�bX�'N�R�v�V�4Yrj�Z6��bX�'{���r%�bX~ "}�����,KĿ�~���"X�%�����"X�%��Nܡvi(��2�7e��y��ɐ�h\�l.��U�<�[V���ٞr{y,K�����"X�%�{��[ND�,K���,K��{�NE3��L����X�݅L��Z���,KĽ�{��"X�%��{�ND�,K��xm9ı,O����rt�$�Kн5鿿�7��k����m9ı,N����ӑ,K��~��"X�%��{�ND�,K��w[ND�,K��^��M9M˘[nh�r%�`؝����Kı>�{�iȖ%�b^���iȖ%��dN����iȖ%�b~3���~-�Y�:�3Z6��bX�'��xm9ı,?��߻�[O"X�%��߿p�r%�bX�����Kı>�AN����D"1F��fd�xkCR�K6��ۭ-�)���v9�M�{k�i�t�6ے])�E����أOc/]�ځg,z�ZRBW��T�f��5$�b7T��n���rf3�G��7]p��n2���.�jN���+�]@�f�{n��{9���ٷ���X��Ln�v�`�1X�4>�v�͂�>-an�`R���n��҆���S�f�\ֲ窇�
Aw�j�ɪ�4��f��;'gkL�e��eh\/��Z�$�f��]t-���kB�M��'o!y
�%��ߵ��Kı>�{�iȖ%�bw�w���Kı>�{�iȖ%���?v^�p�P.1C/���B�,O��xm9ʱș�����m9ı,O�~��iȖ%�b^���i����/'��Iُ��6aMQY�'�,K��~��"X�%��{�ND�,K��w[ND�,K���6��L�g8��ԿIT�Q�PY�8��2&D�;���ND�,K�����r%�bX�w���K��;������/!y������°�1�r�<ND�,K��{�ND�,K���6��bX�'�}�ND�,K���7���/!y�N����������1Ib5�JPo9�로��v:+&`DÄ��З��~�|�F�b8�_t��5�Mz~����Kı;���ӑ,K�����"X�%�{��[ND�,K��^�4d��j�ۚ6��bX�'{���r$!�2,HĐ HF�c,`B�D�X
$ I	2$c#D��P��[!$$��~����5�����iȖ%�b_~���r%�bX�w���O�eL�b~3����K.��d�֍�"X�%��߿p�r%�bX���u��Kı>�{�iȖ%�bw���"X�%���5N��SR�nj�h�r%�bX���u��Kı>�{�iȖ%�bw���"X��H��~��r%�bX���f��
cmp���zk�^�������r%�bX~A#����O"X�%��߿p�r%�bX���u��K�k��t��~�}�m��J֭u�ĪK(v�\Aq��tf�5�E��S5lt\J�M0�j��\��kGȖ%�b~����"X�%��{�ND�,K�����DȖ%��߿p�r%�bX������1ve���t��5�Mz~�����r%�bX���u��Kı>�{�a�y"X�'�߿p�r%�bX������f[�c��{���Mzk�|���iȖ%�b}���ӑ,h������]M�L,�������IR�,�NzKT{����}ا*���"BZ���k�0˅���h�\��l��o�	m%'�s�t��'�`b�nD؎�QuHaLK����r���$��M�SX�x��S`�y����f4�)���F����H�pP�5�>�o�)���6�b��sX� JM��u�Ц��i91d!6��e�T���v�8BBC-�5䌊Tɽ�Kc����D������P�����l��!�i� ���Ą�o����v��I���J2��"y���B�<����Xxa�nWJ%�;�"���@ҡ�_��>БP���pT�x�� �'�>*��v��X� 'L��L��8m9ı,N����r%�o!y�t�qs]Qq�Se���^K?@ȝ����ӑ,K�����ND�,K߻�ND�,K���g!y��S���� � 3<���,K�w�6��bX�!����"X�%�{�{��"X�%�����"�����?���J�2X�/*X%{ium�C2j��t�ػ�T`@q��� �Lۣl��a]d�֍�"X�%�����"X�%�{�{��"X�%��~�fӑ,K��{�ND�,K���>�ִj��r�3Fӑ,KĽ�{��!�U�L�bw�w�m9ı,O߿~��Kı>����[ı/����Ķ��G r����g8�ſ�?ND�,K��xm9ı,O��xm9ı,K����r%�bX�|j�ܴչ�,�2�jm9İ���6��bX�'}��6��bX�%�~�bX�`D �	"��@ @����0 a��+���w�o�iȖ%�b^�׷4f��n�5���iȖ%�bw߻�iȖ%�b^���ӑ,K��o�iȖ%�bw���ӑ,K���N�����˥ŭ%9#&�Q��L[k&��n�EE�9�ʍ�B��u'����6�kTO"X�%�w��m9ı,N���6��bX�'~�xm9ı,N���<�������?w����t��:�5��"X�%�߾�fӐı,N����r%�bX�����Kı/~�u��O�eL�b}�K�-�ę.�j�2�SiȖ%�b~����"X�%��{�ND�ı/{��iȖ%�bw�ٴ�Kı>���]I]\+��ZѴ�K��@ȟ����iȖ%�b_߿~�ӑ,K���o�iȖ%��������r%�bX��GT��]Y��5nh�r%�bX�����r%�bX����m9ı,N����Kı;�{�iȖ%�by��!v��X	%J i�B<�Ӑ�ܒ���5Im^ۭN�Yj�j�`X����W,�ZSSK����d�������[�&.3,�0�X�y��Z�+e��U���x�1u=ÞF�5\;*Z�z�h�u�29�շ�f:ViAlm��������;�£@�.�2�V搤�36��U�*\gh�I�s
���`M��-���
�VV6�0R��χѲ�v�4kfͩ�4	���
+���l��e�LѩEMd�rv�h!�h�m��.�Q�3�SP0-b�.��B})�D�˚�̒�35���,K��o�iȖ%�bw���"X�%��{�ȣ<��,K�������bk�^�~�O��m���7�?/Mx�,N����Kı;�{�iȖ%�b^���ӑ,K���o�iȟ�Yн�^��ߓ�s�	�-@��Kı?}���"X�%�{��[ND�����������yı,O�~��iȖ%��=����t�sRjkY�Ѵ�K�lK�����"X�%��u�nӑ,K���w�ӑ,K��w�ӑ,KĽ��;�.���֭��K��m9ı,K�~�bX�!�~��"X�%��~��"X�%�~���ӑ,K���I��0��2˹�r���-�����kk��3ѴF�{���12L쯺~^�%�b{߻�iȖ%�bw߻�iȖ%�b_��u��<��,K������f�5�O�c�}�h��&l�ı;����9�	 ���"��#	P��������XX9��$�1̉LcH0 RR�&�Y� � �d�`��:�z x�Ȗ%�y�bX�'���ͧ"X�%��~�q|q3��L���U��[%����Ѵ�Kı/����r%�bX��~�m9ı,O{�xm9ı,O��xm9ı,K���˚�̒�35��"X�~@��>���ͧ"X�%������Kı>����K��/{�u��Kı;�t��ՙ�K���fӑ,K��~��"X�%��=���6�D�,K��kiȖ%�by�����Kı=��vg$4[��F����V�N
�	�c��n�3q�t���RV܉t�5Kk\3�?/%�b}����r%�bX�����r%�bX�g~�lyı,O��xm9^B������ś����o���Kı/����r%�bX�g~�m9ı,O��xm9ı,O��}�N@��/!y�ٿ����:�/��Ա,K���ͧ"X�%�����"X�M�  z
a���߻�M�"X�%�}���iȖ%�gO�����չ��a�O��^��,O��xm9ı,O���6��bX�%���bX���~���r%�g8�����6��R�2ڳ�㉜,K�~��"X�%��F?k��ٴ�%�bX����ͧ"X�%�����"X�%�ސ��o.K��qˑֱ���*�ŋ�7�5�}ok,R�Z��\�3�&��/{�Aqv�O��Mzk������9ı,O3�w6��bX�'�w�6��bX�'���ND�,K�z�Nܹ���,��iȖ%�by��۴�ı>����r%�bX���xm9ı,O3��m9�S"X���j��j��%�uu���Kı;����Kı=����r%�bX�g{��r%�bX�}���9ı,K��M����`�*�/�&q0g�{�iȖ%�by��siȖ%�by�}��r%�`E|Nu��jT�Xe�Ѕe�W�ҲC4J�,	)) ,B�@�A��#Y,�[aKZ��1��FE��lZ�  Hf9%�%��B$h���Sᄤ�m"���j��&9\�C5�I�y3�V��x�����ډ��s�ӑ,KĿzw����A�&Mk5�ND�,K����r%�bX�g�w6��bX�'�}�ND�,KϾ��"X�%��P���~�ɪc�KeEou��dc���O���+�#�<����Cip�t�^��צ�{����r%�bX�}�xm9ı,O>��6���,K����r%�bY���;v�й6Q�˝�'�����"}����Kı<����r%�bX�w��ӑ,K��>����H/����j	"w���RRaYL�\�n	 �~��ٱ$D��}��D�D�>����Kı>����r%�bX����f���fK����Ѵ�Kı<�{ͧ"X�%��}��ӑ,K����iȖ%�b{����Kı/��t�rf�3$��ֶ��bX�'��{�ND�,K���"X�%���w�ӑ,K���6��bX�&݈EX0P�$!!��|�)�[��s&��u͎bCM�Nɸ��3U�ج9r<u�@���O;r��wX�\��w8�f�]�����=mq˲TRe���v�#�cp<�z�Ua4�ڦ�ԑ�f%�K�0�턍�=pN�����lT�h��eA!/[v�ÅB�ټq\8W7n�6�ӗ��Ęͭ�ͳ�r�A�b��ˆ��c��i��m���y5�VG��'I=$�ѐ���T-D͚��QCG[�c��alփO
m;v��TV��R�\j�h\m*U��]����^B�<����r%�bX����6��bX�'���6��bX�'��{�ND�,Jq?n�ɹa �Z�ʳ�㉜L�=���m9ı,O3��m9ı,O3��6��bX�'�}�ND��B�/Mzo�������.�U�}��bX���߳iȖ%�by�w���Kı>����r%�bX����6����/!y���(mXgaҙ�r{ĳ��EȞ뿿fӑ,K��{��ӑ,K���ٴ�Kı<�����Kı<�e��Η.�f�u��kZͧ"X�%���w�ӑ,K��߷ٴ�Kı<�����Kı<�~�m9ı,N���Y2NKL���.t�]m*أny�i�[�j���64h��3f��C	b)E-Y����&q3��~�fӑ,K��;��ӑ,K��=�siȖ%�b}����Kı;��c�K	ku��i�_L�g8y��si�z �����Gh�&D�7�w�iȖ%�bw���ӑ,K��߷ٴ�Kı/���w&K�K�Y�[�fӑ,K���}۴�Kı=����r%���DȞ����ND�,K���ٴ�Kı;�^�2�uf�!r]\��r%�b%���w�ӑ,K��߷ٴ�Kı<ϻ��r%�bX�{��v��bX�%��٭[����*�/�&q3��]���8�ı,?EL���ki�Kı=�]�v��bX�'�}�ND�,K�t?��}�i���V]� ���m��u�G�s�ۇ�] �����i.6��`%ak)+m,��]8���&q?~������ı,O=�ݻND�,K߾��"X�%��o�iȖ%�b^��t���f]j�5�\ֶ��bX�'���ͧ �b~ʙ����"X�%������Kı/�w��r%�bX�g��fgL�L3Z���Y���Kı=����r%�bX����m9ǥN�Cĺ�X FE+��D��\B ��Z(@"��k����	�$��s A�]�z/�1�EȞD�ן���Kı/�{�m9ı,O~��씙��j\֍�"X�~Q��>��~�ND�,K��ߵ��Kı/�w��r%�bX����g�8���-ը���X� ���r%�bX�߻�m9ı,? �Uϻ����D�,K����iȖ%�b{�wٴ�Kı;���)��L>M� 5��U�]u�uP�՛��T3k�䱙�ٙ,34i*KJ	L��~^���,K���bX�'�w�6��bX�'�w}�Pyı,K���g8���Ui��$�����8�8�K����i�~Z�Ȗ%��o��r%�bX������"X�%��}��ӑ?�2%�~�O�kZ�\�e�e��ND�,K�����Kı/�w��r%�X�'��{�ND�,K���"X�%�{ӹzh�Iul�f�����r%�bX�����r%�bX����m9ı,O���6��bX ��
�U@e�0� D+� ��x��UM�"{�y�8�8���&q?o��X�H�-vX5��"X�%��}��ӑ,K�����ӑ,K����iȖ%�b_{��iȖ%�b^���uHj�35̺��f���R\dFk�̷����3�^hՐ�^�.���D�`�8Ot��5�Mz~�xm9ı,O~��6��bX�%���[C�,Kľ���iȖ%�bl?H���!�E�����g8���>��~�O"X�%�~����r%�bX�߻�m9ı,O~�xm9 �,�g��c�GH�l�E�S8�8���X�߻�m9ı,K�{�m9��ș����"X�%������Fq3��O�Ƈ��D���s��ĳ�"g߿~�ӑ,K�����iȖ%�b}�wٴ�K����"g���[ND�,K�I�~��]d֤.CZ�kiȖ%�b{����Kı>����r%�bX�ϻ�m9ı,K�{�m9ı,M�	�k��]�4d�zS�T���<xl��A�	$��_V�S=����E�\-�x%�� �_ �w���K��T�2FB�f�#�7p�h�:MЈ�<��|$�@����\���c
͚HE�!���,��I�� BB�ը���Q���D��sӄ7o��_i�4�>ͼ��K���4��0���	��A�p�����!!�ZHKe�E�h��"Ou9����W�螅bm�H�Rs��B@#!p!@�!�xdU�0��
g0�Y`'1՞�����S2`��ӆ���$���B_�B8L�g�Y"i�(�H��"������	�4�;���		(��Z�%�疐��|o}�& l�-���s� B����e���$l�K��4{"�g���+pqz��O�lh|q���ϏaV�g�ϫ���=֩,������g�
a��R(h�LS~{��>�F������.x.}��2��B�XV�UKs�j�*�㍊���9Yh)e@PB��V�J��WT�W0l@��ۊ�O�gì{2H6�h��mf[�j�Vʽ-IZZgrRFLU�΃\-Q��ٻe��+�#Qu5m���Ӧq�����s�x���`ű�pOO�2@�Oa��Z��Z��-�Q�8uds�;�\�v˺�kT�lȲ��+e
i��ib�nL�ɰf���Cn�>1�U�����I�k`W��m�BjT[YX�Af��u� F�Dݟ)�.�:�r8��2���:�S���Z C�O�-���l�*S���X�ϝ3��a 6�	{H��6B�{dMŎ�h�Fmih�[0�������L��9nF�=\��ű�n�F�������N�K.FR�
1�l�Y�B���#i+�mt� X�H	D�h[���n^���[B:�@3Ge:�)Jٝ����\���Y��\��4z���j7Mb̹TS����컦�P!��/n�.ym��7:�9�*jzɷ5$�9w'��O��[3(kr��M�aj�@#+�sl�4�q�[^5�f؀jMrzUt��ޭ�F�6(VN]��[vnc6�:X�Qb��;�J�Um���tA��lA�.:#�NӍ���`v6+:v�uk�g-���s1�u�[��u��BxY����6 ���jH%�i�;�1��l�y�C�˞!�d{S:�%<�s�-Уc�����o&�i��&�i7F[l�9LlZ6���ݥ9b��.��{Hv�8p6;qlK�E܎.k�c�<5gn�s�ck74q�ʆe�9g��m	j��0yh�K6�d΂�%�aA.KY`��q���c�=u��Ԗ��V�ш�\s p"�l6�����^F�W\�(�6.�^��cu��'�4�N���<������K`k�{s���kn�փa�������m�t�A�YܯP&��eZ�0Ю� �����[���s=�����ѩ�{\��"S�l���Y�ff��05��:N������DG��< |���ȼR�|(pF!�8(��H�Q�mE�D�U�5$���.-�I\��v��]r"�ٮ�w�O:�uڄ	�F��#whڻM0��A%�a������/Nцm�X�D�B�{�dx���╻F���v�tu�x�M+��CɲI�t$oY7-m\���6�ؙ��Z^�P]a6�:�p���X���N�qɎ;[U�O��n�9��˜�KQ�T�)�F�f��inciϤ0>�ncpd7`�����t������x����6m\�+���qZ8݊��p2�yyS������)U�rsxF"*�k��ꙟܝ���/!y>����r%�bX�ϻ�m9ı,K�{�l?Cșı;����Kĳ�ߓ���f����Q���zk�^�'���6��bX�%���bX�'�}�ND�,K﻾ͧ"X�%��~���� ���@��'�����/��u��Kı>����r%��a�2'{��ӑ,K����~�ND���ק����̪�@&@_t��5K����iȖ%�b}�wٴ�Kı<�۴�K�������ӑ,K��;[ܒu��jfkFӑ,K����iȖ%�a�E���]��,KĿ~��[ND�,K���"X�%��w��O)����0�[�q�v,s�<�(�;���z���]j2���uB�J�)�Ȇ�����zk�D�=��߮ӑ,Kľ���ӑ,K����a�'�2%�bw���m8q3��L�z����V4�,�ל\�bX�%����*���p6�ND�3�w�ӑ,K����iȖ%�by�w�iȖ%�b|����!���(���zk�^����w�ӑ,K����iȖ%�by�w�iȖ%�b_{��iȖ%�c���+�#�<��9=���/!x}����Kı<�۴�K���ݫ�o{��[4�U��UQ`w%�`}�"wwk�c{q`6�Ŗ߿[����)u�s6�j7\���F�at �4�M���l����u���K%�;^ o�n�{q`��_��\��v~��������b�ȋ� ��X��;�ڰ۫\YLԢ��V�{q`zn�'*�p���A�j�"@�4D�@L�v�:P�&��zܓ�n��=��U��eq��ʰ?q'�պ��v��w�ŀd`�Uj	�W;^ }�ۀ{��X}�ŀ}�u��֧8o$�2�R��eG��R5�.��{s<��ˡ��Lձ�q+.r"��૶����{q`l�x��n w�Zն��;�cr�َ����G�wU�y�Ձ��q`6�^:��@��KIj�>��x��m�ı���1�������
h�%L�D��`����c��=��,9Ȉ|�J'��B>�+������r�~��,���EQ�p{ۋ ｸ��n� �۷ ��֘i[J(�Tǰ��[B�=�m[��Nt�X@�k��ltL�TѕDT�&�d�`����׀{v����/p��U�Ց��YQ`u�j�;�Ձ�����f;��DBA��ժ���)���*�`{�`fc��c��%���X��V��jd�C���ۀ{��XW����n�ϳ~�����펷H��ʰ�c��:�`�����q`w�ōҚ��Y�J�m���e���ut3�'5Z�õ��7W�-�Fs�NČ�ڀhj��f�]�llt0��㴵�sD��K�;rX.#��y#Q�#��O3�wd���7G[��Zb�&q8q<�X�r�q�۝��cn.Ɋ�H��,���nM�����O2�W^���t����.�.�m�aL<�bkl�3P]�����|A�U�P5c� �|�N�n"z��(�G��㸴Ҏk��5�l/f��f�C�^WB��n�tR�(3\�埭�~��ŁՍ́�����f;�=���LӲ+%�;^����=�n,���X�7^s�\l����Z+ac�Y�6����f;���6V769Q����j�FKV��n,绳 ��v`����y���Չ�"�ʋ��6Snl�w���6"ݿ�(��°�M�xqCRmi"=��iC�QɣR�^+\ݺ-��q����D��T�-{6f;��c���-ݜ|���B�]`�(�}�Ň8? 6� I	��H�"����c�T4&��7͛�y{�0������Ȥ���:[,�=�;���>�s�yn���ٰ0w�r�;H�X�۳ ��`~�����X��=U"Z��j	����엻=[q`ycs`w��k���JG* pIn�]aŘ B
²�5"�M�Ѵ�:�0P�鴩�*E56�c�ى�X��V\�^�F��Q�5h�� ��ls���X�z��76x��UQ�@tE�ʰ�{^��k¯�τ�~,`���1~A<�G#��U�l�-��x�����%J)H�f��������7f��bw{=� ���ݱZ���n׀|����N�����:��:�L\T	>T����Fٵ�M�D�srnq6�r{.����!�m�;�_3��R����mmŁ�N5`u�5`�u`7��P�y#�A�Yj�;ٺ���R{��{��}���k<�M�a��)�`wg�y��=�;�ޖՁ�#�T��[$���^�߽���=��ŀu�v`u.%ʒ�|Jwv�`�mh@����p����:��0�n�����hM�p6)�jhR]K��&t,ug������bH��/)\��$�\E*�U��ae]v<�ۥ��c���G9�Ƿ��ը�&e�S3J��t� ���21�X��x�͑���N�L �wj�̌w�-���,�p�bfj"*%�e���^�X{7^��� ;�ۀn��¨H�!*�Z��[V[w�7Vdc��=���LlZN�WG�vA,�n��\eg&ձ�8�����,�ە�����v6g΢^s�K��Qv�3;D�Ў�B'$�u��]�d�N�.^.{k���sD5vM�]�n�JX�9���,�X�f� =�cugm�7����g�-���rѪ�u�a���[�6�b���lJ�V[U�F�j;"�v8h�Dv01�@x�ݳ�k��5F��x�ķ����I���n���������X�պ��4Fh�L�ٷk�q`�Y0$�q�m��u�ձ�]s������,�n���q�":�2w^���'�h�UY$E�Z��ݸdc��=�mXm�^�"1�5D����Q"SU`7n,z[Vj^�ۋ ��~���aS��� �� ���`u�q`�u`fI�l��r�H&e�S3J��n���,����L��� 9��6UR:�$��[e�};y�9b��rܶf
�f���x䅺R����-G]�`{�pzـu�v`n�, ���E$�*�^Y-ܓ�r{�n��bń`�A���@H���N��\�ٹ'�n��=���9H�ݹ�+�*�"j)S`b�ٰ:۸�y��3$�6��͠�8���k���I'�߿}��Vd���掠`y�d�)EEi#���V w�ۀ{�����׀}���ˋ�������D(�mZQ����.�3�[�u�Ňۺv$�[
3c@F	*ubmLh堅e$rK~v�`vn���ŀ���]��m�؀uYV�Kj��n��=�u`fF;� �<��rWmW	$� �wq`{�U�M���&�3�K��hHЛ�	A I�MC�� c�"!�H�p���J�,i1!aNw0����c�|Bhנ{_`����b��d��0H��$�eeU�
XL�d���cp�X��S ��H0�!����)xL1�M+I	�ه�&Y����Hd�!�Bn��G[_*�!�fh�yx��)hR�P�eebYº�ŌHB�1��D��p�����S��o=�3
&�kdh��BH 3�
�H�М�tc���wM����	�!�<2�Fp�C2`K7��9S�/�4D >�}Q�{k�)Qm����t�Ku��G���!�I�Y����HX1�Ќ%o5p�,y��j����)�a���0l		IaHZ�)*@���������֊J �K#�]h"�XV�r� %%�$a1�"FHŕ�
pm� 8|�*Q398�O�HVNk��6��u���B�	!		��!$,.�2H䥄+���H��T]ϐ� ��'8�;�QAY�4����OQ�y� �"`DC�����W�9�b}�ws�^�<�D�eJ�*�
�UE�{Ձ��,�q���� ��["rT�MK��e������8Ձ��ŀw����d`�^�)�xmp
7`�z���\:h���uҳV���c��l�����f3,���ۿŁ��ŀw���9��ۋ[*6�WUU��IL��ş����n��� �}t�:���Ք�Gc�� ���21�X�Xm�^����Q4H��Xu7{f֛�s��ܐz� ,�`� �br�,�� Cꠗ�]޷!��/�U`��U�`l�x�G"76��oj�y�,X��%%��֟A�i�L5�n&"]��QkaYf�䱙��V�B��
�Sb��.]�m���ZXf:�F;��[Vp��DK�2�L ���?�?j�ذ-ݛ��/y�B@��bfjR
�k�ML�X��ŀu�Vo9�^ݭ,w\wn�AD^2�)URՀn�Xm�X�X����y�C�U2MIP�j�j���n���,ok�7lܓ�߾��<�H� �E⇌��X0� �H�o�.,D�t�l�f��B�陱��բ���&�'��ސ���۝%&;*��n�.]5�v��8�b8Fָ��N��+ikQ���kat�]��r�u�c�d�����ЕEc6+�Q��ڀ��Ƕ"��c��ˡü�M�C��V�g�6�������D��r$��i�LE��Ų�-Hlhu����{I��v�έ,j:�2�::أ�tņ�ⵚ�.�T�d������maq���2%.{v�e0+�}���4�*���������tr�{T��<�ݫ21�XX��n�`{cG��#�Z@r��^�X�۳ �v�����]�UFQ؀U5V76[�X�X��� w�~SX�bl��7l���I7�߶���`fF;���6��P��D���D�v� ��� �����ـn��5v/(����Z"��8Ks׭`�1�0��H�qȤ.ݕj�:9�Ec��
�7l������>ٺ��ݿ��K�����?_҄E�n�)USZ7$����- �x��rI��� {�ۀ{�ۋ ���h7d�:������u�V��Vo!&��Ł�;���7G5V��r8����~�M�w����r[V��X�FB����Ui�py{q`zn� �wn w�ۀn�ƥ8�l`�i�ӕW���Rf��.KV6)e��8��S�HC�J9ݞڝuQ�vVU�}���ݸ�{o�$�a���, �<�C�	bj�j�1y���#��$�Ձ�n,䶳�\M��5��,�1�8Yf {~�$��߶n}��X�B@ D��I$��J5+Bb�$�c!�dB�"�2����!B�D�Q|CRM%���3��:��� ���VUbTBT�j�7��,�{ذ<�uX��`}����T�IS��j�;�ڰ;��� �c��Ls`���l��j륰0���!9��۬��Om���1���T9M�I;��uэ7J�V/76��V�����Kj��7^��NWd�"�K0������3d{6�� ��W��D$=��j�����5V�́ܖՀu�� ｷ ����Pv;#h���G9ηU�n=� �c�.�"M��R)
�Cr�ca-jh8M&�.�{ĉ��H�5�q�K�Rn�>������㊙�U+�[V��V�1̀w��#P�a,��K���6�6�&���݈������R:m]u��:2sN54�!L���=���~���q��7}������U�*���� ��Nl��X㸰f:�<�*$�!�T��Y�{v��n,?qq$���� ��~�0���QX���Uf���L�f:��nl69�B^�\v���E���Ie0���y�ܡ��'�6�;���DD@�iRP
R1�R�"�H�������ܖۣZ�M2��F��ɍa�v�ڬ$3O64�Uv��r������dn�rY��� 1԰�M��YÇ��Y���J!ۭ��k��6�If5�qISgm��ӛ�C����G ����t���K�CL�F��v8݉� �GE+x�rM�J�)X�ғ,s>KA��g��^ 9�m&�e�x	����4=��X�닭��:0!�+��"���BH^k�t�զ�s#&�`Gj���I[s��f4��5u.�a���GeckUƋ�Е@r���S���?�vn��Ƿ�Du��X�����)JPMD�+�-�؈�!#q�ŀc{p�=�=���zU�69��`?c��f:���6r[Vp���F[,�N �Հy��0�{f��׀n�q`�嶧U�*�	�d��Ɏl�mX㸰f:������)7�a��%�@4�6�]�i�.��^8{8� �	���t�\�-x�lX�3`w%�`<�e�{1Հܘ������q�c�������j�8�s�s�
#����`nɛ6r[W���l݂�?+#�-n8Pr� ������mXmՁ�Tb����u@r�v� ��u��v�~��8���w��7 ���b�WDԕS`w%�`۫ �c����~N�&���.�o����)D1����,��v��s���Fe��V��h���װ�.�HB����U.�=ݫ �c��寘wf��M��4�~��#�Q�p1�呙6ru� �7V���m�NV&���W�`zn�>\E�����������w[ ��߮��u������U,�Fz[V,�6��B���^��ٰ<۬���Q�:�r� ��� ��?~ݮ��l��mX�TÒ%(Q26ѣ3p&�WK	�4�X��&�s��T�x�؋=oeC��q§e������́��Հ{��X��
�1Q5
j�&�6�n�X���m��K�l���?aeM���Gif <ݫ76玬,c���(��N���t%� ������~[�� U"�B�= )�賚������_��eq��2K0��rF��;�Ձ�́�8��PML�Q�a���j�G-�\j���g9�/=�n����A�Ԋ��U;�[�w�ݘ��XX����GP�����*R���VK0�ݸvn� ��� ���0��^������[�y�j�31Ձ�#s`mՁ�$9��aep��L ��� ���0�ݸwn��3�F��B��U��#s`m՛�n֖��X'E�}�{�$%���s�5��-���s�������FRS$����b���<Hjb�$��P3���y#9̈́�<Mo,��i=޽����f0�6l}p=�V,XF�ح���_'ҕ��	8X���Č� @����R4 Dx밧�7�J�0�9��nz�!$��n33<c��G5�<�F�h���r_)�<ٌ�a���>�Hn-��k���{36�� 3�n�#%$H�! �s+	D���І�3�H$- y��Iѡ���A�j��F	/�K�!#,����D�h5rEU��Li'��|E0��N]K0\Q	Y094K�}˛��%�f&ص]�A���CA�}�(س��w��}9䳒����&���y`y�G�w#Yu���vI�	I�n$��H�v��]ĸ���8��H�(�3��9D�����b�Iί��!0�����
[9s��9�%e8�4/9"똇Ŏ'�2X�bE���R��Lמ��_)<�}�˄�xp'�d�xBjh�B$�.$�0᫫��7��ɞ<����&�Q�Cu��fǘkF����	�[of?p���5���2�+3{%�.eiy]>J�B�U8�R��Q�(��<2��Ȱ߳�C-����V�US�i�����b��l����,�
�*lr�T�]Ps���ݓCM��KY�s���]���f��2Rm�]��X�k��#�GL)�R�$B�R9���77C�nQ�i-��N6�U�d,�kpKvi��T�44e�����C�A���Gj���f`�-� ζ�n��N4��`���o�dޘ�Y�m�ɣ�S�c+r�&��b��f�� �m�J����#b�g�qy�S����rV�n��x�����ti����i�S�.���r�4l4FջLd���b6����@���az�U<��k7Dv�6��ʔR�N*wZV�2\=Y�lci�^ C����s����wa\����q&����V{֔���w�eSqǝ��5�rF[G;�H��9�n���c-]s��p#�vnB۰�ma�@�d�v��8㗦�3��vL�l��\k���kZ�wt=Cy]y�Җ!��M�2X�5�̱%I���ME�n��κL�m���yOg$��x��)�]�k[mLV=�w;��x�C�9��G�`JW��"[3l��4��[�H��p�7WkaK���/'�st��Ѻsiv����k�Cj���Q�\�u�p��H��GS���k0�Wp�ֶik���56-W-��<�lm��g�0k,�ĸ����Mf�&�@��
�cK��.p�K.obbg3�+��"��X�q����F&�Y�'.�.�������L6���.�Еc���hR v��逆�v���4�L\�P��ɓYܟ?s��TM���.5��X�VԲ�2Uۅ8��kW=���o\X�<���Tj-�C�ru�K�Ƃ\h�\���k�QK0�q�0����浌c��5�a��"��`Qu��;s�dV�v'D�܍�.74����["�`�#��H���<��s��c�#KӺ��h{p�ey+a�I/.d&�� �j���,b뜻����`��+Ha|](�G1HLb�.�*h.�S`�P`L7�w�G�!�*�� C��@� ~QH �O 6}�s�?"� @6(`@�<>�{t��{���-����Jji��f��ģ�T�P�m%5T"��.��K=���D��[o'G*�R�MI�t�ưY�+b�74;]j�btb�[{�������m�3gn,����+)v�����<n8l�plY}ۮ�2�m-di�L���Z1�j)2�p�+pJ��aړ*�tZ|��F�������A7�ՠ+!V]a�ūm�ˌ�Gf�ۆ��
4v�a��E�:OI�'d��?K=�o�K��ƛCr�X̒����|y�,l�d_X�J��ˠs�v���t���Kg@7\��L ｷ ���0����ds�*�Kn��玬�� �7Vp�Pڰ�Y�CrS ;�ۀ{�ݘ�M��߮�߯� 7�[+H��R�X�-� �7V��X�:�3چ T��,U9^ {�� ��׀�m�=�n����	����]��)h����{[9��&�g�a��F��f,�n��hqq�Inݛ� ;���̑���u`fI�
���&VMj�jnI<�ߵ�	�>Bؐ<���G���Dg,3�/����7L��8�g�њ�?(�[H[�n�������t� ��Vd:���R��R�jJ���u`y�e�y���ݧ�� �7D��S�WB[p�X�:�3$nl���:a����>��Nq��ȡnc�u!�j���'�� �E5��X���nbtR��-��<�Ձ�#s`g����G9<�Gd3v�����H�;�-� ���3�""N�5��<u{�D$k��M�+/!j��`����7�u����
����|��_��䟿a��}�wc�ګ�Yv7+�7�u��Y�Z�ݛ�wU��$c�&k�ML�ASS`�u`lk�[=�wV�wf��nU �p- ��T�3qL4iB�a�2��i�cFlb�e`�us�!FF2�:@v�}5��=��{�0��p��=UH�dm�ـ{%�{čOvl�X$nl�0�T᪣�Wcv�_�f w۷ �Cv`}�p�(������ ��69K�X�ݛ �7VDz"H�X�EƱ!	�;E���8
�
�\�3��$󿎗$֥�R[�{�ݘ�n��7^ w۷ ���7dh%���Z*�ruq�3T�s�5��KXŀ��,�hK���p���j�*��M+�nl�s`��n���v;m�`��J�,�5�����$�j�ݓvl���3$��*Kƚ�HPv� �n�v��I$�=ٰ5n���LD��RQU"�UM�܍̀{�������[[�TU�F�,-��n�^�� �7Vr76�z8�v�i
*a*�L�Lf4�`4IL,R�W�՛�D=q��*�z�v�Rzz��]h�Cf�4i.�,a�o,�@�ɶ6\oF�ln���cнy�f6}<(s`�=4'gv�0um�j1��Ǜ���ùγac]y3ݱ�0�+W:��[H$̰���x�F�3C�ۭ[�N0��\v�<���svӆ�S��\�Z�Lcɤ��ֲeִj�i��UMs�&W>P^��R�ep���<-��Ϊګbh�5%��[)<�<�Ÿ]���5����7�� �7Vrӛ �7V|D��XWllR If w۷?��������M�cݫ�noyĆ�l)���!ISU`nέ� �7VX�����n�q�&�2��VK0�ݸ �u`���b9ŻF����RL��(섩�n n�� �n�ـ|���-�����Ҩ�e���g��s�9�m�mʯVS
��3r	��6a�x�)d��Kp��n����>}����v��N9�M�*i����M_��s�9�C�r9�b��`�� >����SaTRƋ#h��^՘��7V}�$y��wij�;y���(�r���ݸ��� ����?{f��=֬+�6)j�������7v֮���̀<m����}4��@��V��b�n�l]��!
}���8�\�F;Dk�X@����X��e��ׯ ���0}�$�>`ww��?~�U!PӅ�-C�� �c� x�XsXc�6�T5#�ZZ9*�[��ۀ{�p��,dE)a��@�pj�"�qQ��u��ܒ}ｸ_|��;�K$��[�w�p�Û �Շ��G!-{�`c$�R�P����[n������� �n� ��ۀ}��ƭ8ө�C�*(�(��6:H�TCFݡ�l��U��	�W��䎝T��F�$�� ��ۀwf�����#��P7;�C��P�LJ�SJjj�9m^�G! �=����`����b���ؤ%��}��y.��Xcs`<�I�J��r�8Yn丹ğ��������f�D�� ���a1"�Br���Dg�/��w[��Y���B�QX��� ��ۀ5�̀w1Հ�\5`}���̮�x�r���&�s��Pc ��r��νF{*�G\:�̕eM��mJ�/�����`�u`<�XsX^�!���%��5R�jl���������?=��g��6n����`+*i����cU�w���k� �Հ�dk*��"��$�W�w�p~ݘ�c��G#�e�l��1El�S��Қ���nl��VX�̀w���$�M�E$dH�$d� ���X X�����SZ�JдX�n�X-Yq[I�B�q��Iݚ���C��Z�C5���q-��ѻaH� 82d��Y�Q��ݎ����V�r;z��=[���V��v�ׁlO^�=�d�KI��Z\͂����إ�kc"�h�H��i6�5�az �m�rWi�3궲"ny�܏Dg�t3Aui0�3W�XM6��W��Ґ�
U��!�^�s����I%�����z-��[��!m$�i�e+�T )���V��V,�z��4^؝U��Y��o���l��VX��1Be�ET�%�p��_�l����n� ��ۀn�;�B���(�qـ{�VX��sX�Nl�RN��	��n�۳ >����^� ��ۀw�~��dC��K0��Vn�V��VX��
��E�B2���(�+�Z(��7f͹��2�ƅLV�^3q�k�:���+,sZ���@b�d����;��`b�!��",��]v`~ݙyԑ�/..<QC�1Ar{�{�ܒ}��krO}�n��8�<�ѫ��r�G%�K�`�2q9�����%��k���`Q�0}�pzy��5�v`~�����������%�p���32�VX��O������g��c�[�f�������4Ip�)���l���� ��+�Ɋ�6Ê]�ٺ�=S*��{1Ձ��̀g��3)5`y����H�j�-��}� =�����MX�ut��H����`��C��l���p{��ýRq$/�Ô�%KB��`F�ف�M�t�a�X� Q��*QM���Mj�[�I����fS<�Z���6���ŋ"B�i2�˷M)!�"Z��4��a����i��a6	i��E�)��c�>c���lwA]�TȘ	��y����ŖX% �I�ip��em0�	µ����krH1�w��H0~ւD��]x|�0"�H{m(M��0���,�&��|�o�B{��9*_8B?}����B%�$	KX����hZ2�x��.OBĒI
R'��d�ZR�|�[!$���1k���P}���i /ĀJ�OM����Ռ��a2;�c�$�du���F���Z��-��6�{-�-��i!,K��`c4Mz���4������y�0��A�$���-.��ޓ�.�I���RR��H���͗.$L�&YI�l��Jhe�8h��!KYH�X4��"������1��^�3Й�Yu���O ��������R�	���l'r���	�d�<��{���h��P�W�=���v'�>��!�����`���Dd5����H�l�����@�_�`���U�  �}GbmV�;U"@��D�I�~AMlٌڂ#��)�=���O+�GPj߾��J�)�L�(E)��32�V��XO�o9�Bow�~�7�URDX	�x�ݸ^�6����Rj�3hs�7cNzd��b4U�Lp�I�Y{`���d��V����]�P(��mq�&2�m�����,�I��9���X�	��'m����0�ۋ `q���s{č�QS
��ARB�SQ`f����u`5����c��7u��B���QYBJ`�ݸ���t������>D
t�9�Ԑ
�%ԃ�,7��dd�
$a�bX#�a���!��?.q)��|`����KknF�����76d�V�8Հu�V�7 ���GƤ(���\$�q����9��5j�!�N%I�[�4͗#H�iq�J[f����������'���b9����V�M�� �&j*R�<�Ưb9�A�ݫrwU��8��BCٿ�UT�H��%���~�p��x�=� �����i�7H��R���c���ܭ�`7/U��N5`n��>�����m�um��=���'����k�̀�D����u3KX�j��U%�-����,UЛ"fh��֑#L\ٳ�Z����ǭ�b=���N�i�mR�p㤱�k�Q��=�Vˑ��D��1��25�.�s�k�de�͓eⰭm�Au�M,. Ď�̬^��x�dE�@r���OX����{��d��a�x�D.�y��ϟ.ͭ&+��kr�̵r�M��85��:ش�l�	3Mp�QLo�rNN|}�"8�8�>ꍪ�Dܲ|�E�N^��M�8�h�pVX�3un���mlr�smu<f��QSK�?�_��Xy��3'���wl!F�J���%0�ݶ^nl�Ƭ3)��Ȅ�n�Tî�\�YV[p�߿L��ـwO]0���݃���`Dԭ�Km�<��l3)��7V ��X�MLڄT[F�%� `�ݸ�ݸ_}� ��^`�q8�!.���є��G�}���]����u����Ȑ9�����D�A-$������ۀu��0�=� �t�OV"�I\�.k[�O���oǈ�>(B�Fŉ�B����ČB�(EJ�)��P����G<���M���;����-�e-�A:�N�p�{f�'���ݸ�ݸ���,R;X�`y��Xq������N5`~r����T�+NW�w��6���N5`fD�V�CoPGB��d��[��c��;n4>�\ca 9p��6#v�Ժ-��q
��L�W���>mX�ƬȜj�;�Ձ��c"j�5R�am� 淋��=� >����v���G��QA�F��ׁ<�g�]�'=��np�æ a#�G�p����CP !��~�����0i=�*�W"-A-$� ;�Հu�V��V��e��0P;8UIR�R���:۫�X��@�:��;�ՀGO&I�H(�)$���ݻy�qA��9`RV�m�l҂(K��-���J�m�	��[������ }�ۀn��7u�b���]*���=�S,��X[u`�u`{wr��X���������p�n� ｷ ����vn�!J�kvX�ۀ}�u�����^�`u4�	$vU?/��^:�k��rO~�~襵5R�e�׀{���yz�mՁ�-��DG9퍍;P���D�Vp��`�.�y�]v#pf���lѴ@���R�V�X.��ЫQZA���{ٻ�ym����:�s��#����zK�
�SB�U@L�LҰ����ḿ�8Ձ�S���8�ě:�kh��^6뵒[�yn��'�3"q� ~n����t��a$� �Ok�=�=� 7�� ����=���L��Y]p�9U���X�u`u6���j�#�B@���ʄI"! BF�9f��W%�+�mX���n��ƦՖ��LLXRR��I؇��l�;�����w�Nc��p�Ʀ�X�ӈ�c��5۪�e�x[๷��֍�Pe��U�CA��٤R�bMi��@���Q+R�7Li��rG������z�-�6@vi�j8�I&��G�b� 1��uv��D;t�����ݎ|� b3�Ӽ멌���0�	TvR�5���b�t�� J�Cq�L�Y2IsVJk,�\�e��*$���8���٣$���D糓��u�P�D�(��SI�n}�`u6���Nk�;�{^����~DT�����U���wf��N5`{	Ƭ�X��E%�S�Jݕ�f��k�;�{^ }�ۀ}�u�t#�ʹi�h�U�V��j�:�Ձ�-��́���V� X�ZI^ }�ۀ}�u���la8Ձ��l�$�2���e.f�-�ں�A��sZ[������]NcF��Ln��GaWk���=�?��������}���XdK�)D�R�V��x�=�K�$$���J��(�@(@�;6�&;hX��� �0k�G��WqޏI���g�:�:�s`?5�1*ԾY]�W� ��x��n }�� �g���ܪ�T�Լ��rY�<u`x���N5`{'%́���KE+u[-�>{��=� 罹� �}� :��58���Z����z�9�;�8�9�0��]+P�*;��NoX��%P�erـ{����zl���p�{^�Hިm���F»^�8��q��:��=��X�ƫn�)
�d�Gf }�ۀ}���� 0Hi @�B�4B���H@�AeR�D�@���Zk��}w$������8{�h�-�qH��-�;����{^�Ol���nފzi\%�����4�d�V��3`���y8Ձ���՝�_�`��tb)c�Ŗ:��:��v�ɉ�XR�weY�GE��O9�zb�jeM.��^��[u`<�j�̜o �n�Q2����,U�& }��'�3'�1�iX�aʘ��������x�=���[��v�={�nT#�,vZ�?.q�OU��kR�������9�I\H�ZTE��8.}����>����eU

�X�4����1<s`g����9�o����բh�Gd6ŵ�[XQŲ�+�q5KRY��s���W', u^G;�5Q�����dr��@=�߮�ـfN5�����Z���֔t�B�Jj�O��$4�̀�kR����>�S�B�-%�ـw���n�V��X�9��j$SrI
j�jI���9�rݽJ�<�j���l�>�����̪16Ԫ�B�J�;�����qֽ��:P�e��_����TU���@EW�**��PU�Ҡ"���@@_���@ *��@R
�D"*��EX
�  *��E
� `*��D ��EV"�`*��@B�H���A
�@ *F"� *X
�
�B"� * ��@�b*H
�B���B"�
���H
�"*��F� *��D *���@�*��F�"���@`*��"� *
��, 
��"�
�`*�"Ȋ���0�*�"�
�`��"��"�
��"�� X",b*T�"���D�"���F�"��
 ��ED�PU���"��UY�@EV**�_����@EW�**��PU�J����TU|TU�b��L��x߮*"� � ���{λ �������B�R���݀ �P��K�J��V�v�($lĕ$� �A��d�@  /� ��QUH�AB�R)EPPRR�( *�(T�@QQ%	U$���IQU*�T�(�J�      `���P�S�}�}���<�s9t}^�>"�ٞ����z�y��y�y��x�^z��>��˯�� 7�ӽ�x��z{϶qzt�޼\}�r�'���>��o}���o}��ڪ�j毻�g���w�n�� Ϩ@J��a�
h�>�8N���W���8��yۥ^��(8�YoX��wo;��g����N���y�>�k��{��E����y�����xz2y������N_v�[ͯJ��R�����������{�yo3U{�)|>�  �P ��`D��R����}���b��&�-�z��>���Qf�{py5�g}����{����ԧ'������@\�Η����^x�ǽC�g�aq�z�}>��m^i���y�O\��μl���y��gU�T�U�> P  
� 6�����N��}���7�pz �:����N@��� bt�:;���SӉ� �Ҕh �1 Ц&�J0�l�J
bz:� ("  ��)������`����OG��b*�@�<8A@  *�)�c�5�=�/����{�/��g����/���&��w�O=��q2]p�O�O#�� @9�q>�z��z)O�ϥ7�ye<����8:d�� S��NA�1�d��q�@    i�
l*�@      OHLR�(i�0  L��=UJ��O�j hh   �*TM��FF2`�h�2��2R�Q� 0  &���T����4�=LI�����2����/������Ma��ݙ'�����8N���PE�kU?�'����AU��PD_����G�[JS@D]��?�?�q����$d�G@ ",+ �AAy�@�DX�9���*��� �����baO�S����������e;��Q��C�߹5��dm��f�.���3�;���ӗn�:U)����z�.��/��o������*/ =n�a����zq��S��%�PJ�)d*0sH�I���
�����.��"my䄄CŃ�P$"CGn�OM�\{�1)���P5B����2\���x�VZ�����H�	��8��B=�8p&�,%_�嫺xg2�����55�r�'���M���lk �n`�JHM�[oE방%��55�}&��#򺔔��b;�9��X;C�^�H����Ҳ����iK%;��v5E�՞3d�%,�\ђ`J���P�A!40AUEݻ�r"R��g��x<r�srx�}_q���i�I�H�ƞ,��z=*�:��2��;C�(���T��4R����:�AS୤&��E:7�!��yR� 3��&�1����<p�v�����C���J^R�#)�fV��Ĝ5�f"C&�C��N�\	�'K�D���qHy��t��u�?�j�s��G�j׌�ղ����	�6l�i�y㨙�D�V:-eE�Z�\�Ș.�sT�BO(�֥y��-18�BM\M�9�7%� �eK"" �$\߭1������P�;2�cFR��9�fx��2ܖr���*��+��UmD�Hm��Zl����,�3,���V�$��&313�CUԦ.rovQ����p�"! �D��{š�xlb" L@ЂcSU�BKo�ش)�$+��6��vR��u�N�C�8��>�d��7���IǛυ.	JP��&�촆_�̹�}�d�t�}'N0\8��\��d.VY��-(I���#V-!�$�M v�R����[{֋���֓! �G�����.˺D����K�B�Y��6�be���ܹ�)[܊�Br���{9�O��5����&N�����U�{�)����_�F�X���&���R�L�q��UxEUC������d��3/�w{jM��BJ��hS�������7w�(v�:�'��"|C����{/k�t�xV#�/�*�I�{¹Y�Y��(��VC�9�v�M S|�+�^Vx�Qc���/�s���5�툕� X��j� �ZDj+ɍf��Z��L5^&�D�D!bW �VB	�O�T�B�ƶ��y�2l$���$=���z�g�W圗tZu%�V���}����jBja҉V��BbD"���}�Mw<�p��9��X�+!/*Dtz��T[�ɧ����d|��#��h��Y�j�"|���O��E�L�2�a�V�ת���%e�:�E��^N��ego���yo�,��[������d)�޷B�����CZ7u�U�.&�l���9����R�r�}\�eP��7.�3ٗ~��	��&<��zP�mJb��+Zmb�{�V��Jt@Xɦ]\�?e��jɇf+��r2Q=K�M�U8��@BwP��}+�<{��sD)�\٤�4��&�^�j���^�3j`ku{ޔ\��A�CQ*$��ǻ��VN���fݛ�"М!���T�z}�(�.�"���Kf�1�\�
����ceva���<�8JnD��^��d�{�J�.}$��s ��#Fv�"���LGAwZ�&�� ��mg{��w:}������Cz�ӗ���7��\�ˣ��l��	s9��#i�ۗN[�L+)HW1+hN$NG.��e0^��	�uAh��/2l�.@��O�UˉWj�r���B��e�\�j�MZ�TDl$$�ލ��J�ݤ�n�]=*�ς�4RF��$�"�;�f�]0D& �1T��R��}0?+���9o&y1�{�ވT%�(V��[z&�C�`�1�����u6��	M:VئQnRh�-
P����ST�S�����p�B�#�6derU	��-��ىr=�3��e�NjP�!H�	B�´�3#��r���%I�Ni��V��/5(H'QU\��%X	���J.�6'5�R,�^J�����sBl+��`��;�<��k�V�#Rڮ�HML*T�"<�UӧJ�=Z����U�ҁi㫮R������{�h��h��&}���%Hr�u'0L�ф�!CE�w�}k��=��Լ�v��Z�~�T�5(|;�~T��	�@��y�w\�p�З<m�1c�p�*RK��y�sZ��S�w�Bh�!F2S��KjwTB�.�D�&�h����t�Ǉ���CA��\�2��ys�Sm`�z��4cp�"�I12�$:��ٔ�2J�[��{�۬��޼�X�cn%)��b�-��7���5η�}e�e�{��9�\��^,!΁/��rs܅׎n��ky���k�s�Lw�0im��f��9P��� r�%����<��4�rjeN�D[sK�z)�#%�Y}��_��/MŎb� FSδ��
Ӂ"��$c�-b[�tk����H$"抨µ5i	����sޡ��%>n�#r�s�9�9����j��яw"A�{��a�١��e��m��j�����w-�^��:�w�Kq0FE_��V
@��@���� �2��hR���(�\�\�W��\�a�U�õ̷�b�=���#�Ų��F8R'R���"��wҕ:z���w<��W�B���
�B^nj�!)�]�2��:*�@$��[�[��a
���4xxU��QjR���׏{m:L�B%߲�4eߪW��y�%
���Bb�3�{~.j&V�%P)��+�!fא�j}h ]�!�
��D���3R���v��ݴ�0�k�Ԯ�3��}߼b�YL��
��M�[�Y��=�w�&��]�!���i��^�<�[N�����:�#P�l�?{%Z��:�SH�jM��ô�O'#�rۧ/"��b��Z��R�[Hx�$$�D+�a#n���i(jg<$|"]���̶�����],�M܆zh���k���Wn��$Sy�T���HwwR�S��1+�o����i")}-z���6}Mr)E��G��J�NI����O�5��)s9��2�Ѿ
nM���"SfFhcT��B�s��R���=�T�f��JR�����R����j�j��MLo��w�����FU''���Kv���۵N�`.�BqNBd�s����3y�w����Em�����G�!��0{�Bjb���]1,UQ��*��bzo�}�P
`u�q��ǥ'
R�Z����0��h�0��6l�-2H� �5)��h Ԇ�)�%�!\�%d @�aT��.F�.OsP���%ٶP��sN��KB ��cI���4�3r�wN�'�\�����t��O�U:xt��{��9.�@�ۢ�kFH@���IS|�������m�ʀ�%��-!����*�sw���՝��cѶI�u��Vc%��\	�m��1%rV7L�CG�6{������'=pG���!��9���=Uz�)��@����HC=�g�տG���W�[]b�m@�!"P!45i(D"b����%g�N"T��ȴZ���e)�3�/��V)��N!L��)�n=���%F`D�x4i@�$HǄ�(0(D�ˮ���ok���X�'*���U��=�W��B54� $�e�1�g����lA	�C�8CT���HUX�<m��I7'�8��>�[��__��,H��c��f�qe�r�j��yn�B�T��f����+�I��-�F��ܓ��j���uR�������6gdy3�`�=���
�A�%>�C܄��J��%�7�:�Uw��9/��1�)�Q��y)[�R!Mq�b��"S-�$��{�'��ʧ��4Zm��r�0�#��������N{�쁧2�J��xf�(�6�׭��I��"���I��+.T�i%딜)e��	�w!B����9�<6��-Hv����Lz8�w�:���!
�]��1�ٸ��5TZ�)�V�.�D�����`MVJZݧ�zڳok%/b�<��y��m��tjmYM��S�I:H)7�*�"t��2�K���T	��F�z�����[�Ǜq5'�-Z̯bn�ؓ�eԥ>�E473JQ�Իݱ��,[Z!�`�)բ�z�p{��ӏ{�e]�mMZ&���	��SPY��4_K�2k���̥S�����7:�drR��&�h����0�,.kd.1	��I��j�JZ�[���n�G!j=�Zɚ\��Q�.��^"bv��o�S��� ���>�#�$)��7n�+�r2��Fc�޺�b�8�`������f�����P8�zf�gȼ����Dℳ9+���s��6.�����|ڜ ҾI)A.yQuv�X�O-R�IE$�cA�o�w��/XP��DЎ+�1 B�*B��*�iz$CX���V<X+�
T���\5"!�1 Njk��X*M]��T����m��P�日��E+P�7�c�\�IEp�W�����,�CĄ��)Ϧk��NW�������v"�糃���YH�S�v�h�ՃĜ�.�Nj�:[lL�	��WA3Q0J�eM�>���S�4uXs%��5���3Iw�]�_O7�LU�rͮ�l�����O�5���X�I�jZh�a-
���&h
V��@�H�!��%��/ҨQ㪗FH��/��\�|��������9v#Տ�
М
�����Wm]�D��޴�~�"�	�é��Jwx��U�� =zb�S"'�5t�QP��*Q5W
Rm1j����Jf���B5BV�o�cͶ�T�ʖՐ�;��Q74�2�����"�u_��<�XX��'=7�f5�'��S��Q�#W��Y���Ԩ�!4&�PM%�$�T�HJ�^���W �擥�yT,�<��!h�ZML+�۱�h-*��b}���i�DO�5nBU�6UxJ�h�ua�sy���k��|�m�O��$��z��E�Y���k�*�5���_�>��0T�\�&3���_�	�53������DB�v��T�Kp���S$�j��(�kF�;JK��Į�nZ��Dd�!R�k�����*���^iB���R�E���+�064h�e礟y�� 7�+��z�6�m8\z��B�R:sm�	<Z�^�6�Vj��[�WwUb=�6�Pw�B�F�W�v�	o�*�
%�e\��$�+�Q����D��Y�s�Eh�=�yʜ���Ycm�N�o�7��r�CJ��D8����b��9ʒ ��r�#�%GUt(�R�X�yW\�kb�隢��J�U~����
��[[*A>�{��w��2�2��h�M�K�bE�w~/��������������`       �   �      �    m�  � � ��   l      q ��m?|�  �6��` p  ���( 	 �  � l�  h�        6� �|  $	   ��  m��   -��  Fɰ�:��1�WX��ڤ�om��sn�k)�m�-�wjt�8�v���+����Th�����,�^l��
����O8�I`�Er�wP�p�=�l�c���	�����m�:�m+v�f*����ۉn5�u��I#���l�ի�2rGH��ͬ��`�o[@A6ب�g,���P&:8F�j*I-��i��z˛$]����pqv]ZLjɴ��&8�J���%;U�ݙ֎����n�;V��Γ�7:A{s���m]=f{.��!��ص��s��jIr���ț$�Ş�h43+k��ח��e���S��1s-\<�7G%�{�ci�Tz���V�:���%=���>�v]Z�&U��va�9�k�O��eܞ�:�&��&9;��5x�up�?b���o�y-�*-��9��:���`<Z�J�n�t⫋���l�v�C�[q�c5���u==�Z͖�T�9��"d��R=�:��,Y�m���FCCl<˹]Fݬ��u\]d��Ȏ�����b�Br�6��u�e���,�͂C*n��V뵛���7Zt��m��O<6����UnsT@���;�$����d�L�J�l�6�8z��\I��8��:�&��ݺv��mB�Z�Z�J�]��]�f��K͸�|	a�AQal�[�u���㾷b�Α֋�e�s�������j����_>�2�^͛��V�S1��������*�Κ�o'4�G=O�Gq�]��Әƃ��Uĝs��P3˛n�]�w9�Ngg��P;!y۵F۬q�g�lְmm����^VGVc:�`�Sg{e�dv��[En�N�M{h�:ν4��[d^W`��8�Uږ���ƕ�ka;kp*RV��PVݯN�5����zW�Z�����ɱ�!��8�m��Q��8�����ӕ��#�v��d�v�����.�<�К�kp`���ݴ�����n���&�\ l �f�  � .�u� Em���H�f�f�����<0\^�l۝�v�꣊��u���6���>�b�`�{":���v�l�wd6��{F�^��:�x7fv.���r���==�C�h4h���p�6�s;�),�Mdt�V�q�Y�ƴ��wl���MM6y���W��Y��8�L^b7m��$��^%���[�7��	�v�Lj�2����ˊj�T�[�se�V�z�v+)�g��mc{]e\w ��v���6�Ʒmm֘u
�:��I���!��͒lP��|q`vv2,��2{F��n���z��.��[=���<������7:��mڢ��f[jU{k-iؙW�w!Yu�2G���ul�Z4�㶸�셷mm�:{sՊ��ݱ����<$b\��,�@'��b���8�WԖ7Ol�At��H*��ժ�hݎ�9�{�a�6L=���}��Q���U�K�����n'Lݯgm�M.@����m]�c���ڢ�X���{Ae�rm&�V)�eT�,��A��Y�1׭@��D�NZ����ۂ��Ω�n���u�㎧��m5��k�ĝ4/K$�	93:E�a�[q-!$��n�FU��]m��H[Qsإ��6�3���z����q��c*�g�;U���wSmC��ԬGv��j┥vfh��-���˕�)����H��FkPݶ�.�8�/Wc^Nw+v�.�+Wc��2t��y74�9��[e�t^x�v�4�Y���6�4�F��/���ʶ�$0[B�v�ݷ�]�n�04�Ja�Z�T:���ό���l�L��9�ا�i�ō����qv�˅aqӭ����f�L��xuӝ�ʩԬ��uM)y9:P�[��n�sT���z�8�\r�55�}l�xu.:{�#�i6�#�íC��]��>�cکL4&Z��ˍ��.gW�G������*�\�nՄv��5��e�r��6�6��mz�0mdP���-T˷�Ϥ:�MW�dm�'t��Q���l�Y@4���ӛ6Z�����yu�%H�r�/nvڎ��ltZ�ksYwb�Rx��kXwm�+S�(c��ƅ2�<�d�z���XG�����yz���wk�8�ioE��f�M[�u"�4����k��SK|/9���.�~|���zM7}8����ۃ��m�s&�]'D��H]�mi1�v�t��p�@�@�pg���7Q�Ԁ��m���G��uI1j$��5�=$�$�KS9r��i٧C&����)���3l�q*�9���6�t��PF�95;���v�c�-w^�frF�6�ݰj���Y�@�R�j�'GBY��`�a�v�+��\�m�iuVUԇ �#�A8|vūR��y��	 H۬��I�CA���i��&̼�wa2^��؎�Jo^N�zJIklD���.혴�D�V�Q,��Uىa��/kU��\��v�I�;ZFö�ٯf�I2�T�9�$��gMv�L�l�[VK�[-�R6ݶ�%�m$6�[�����+��m�nn��-�4׻P-.��Os��&�8�.�4�k�R��M��.��
]��m� �2�],�e�m�Bt�\g����kn�:�Ҧ�ʴ��Hpv@c]V;s�ڽnm��HN��e��+�7g���V�tvʚ�kճb���4K@�ydMd�\H6Ӧ�f$�Ry:�^��X��[9Y��V���]ڷK���u�ֆ�$%���W#�ێX��U�S`�m�`�fw�j�g;�m�[�S��-E�r�q�6�l�se	�skF�N���)�D�A�ݶ������A4�oM��Uu����'�J�n5�3n�t���q���i��\�`]���}�tuM����9:fw�x�0k+`��Nܾ����+v��j�����~��~���c����Z��]aV�wN�m��!�{�j$2��q�&np�!�e�gYu�õ�v3�L����sVY�U���v�������n��U����Z���'�iP��0��3������o`]m�6�>k�N|��a�WT:���Ә��X��M�K����x̼��m���v�T6�m�n���V���&�ඈ�*M�|OglC��8�6�,06��g.���1�m�.k<��c�U���(;l'���b�j�%��l$��x�l	 -7key�� �.Y�B��yx۵���s�2g���˶�<�cm��-͵��m��F�Ӷ��p�:C�7:^=N�v��l[i�Ӥ��h�Aì�"�u.�W9��	�t���]Z̵V�x��#��G��vJ �0ps�w<���'.��0`��|jը:�ڎ�Aɚg�֌X�Y�\O�m��f1��9�0:�)�z�>=�|�a3�3i9�]��Jx�^�w[Kd�5��;`q�c��/KmN���Xû�>|��g]�ݒ6���e'	��+Y��V춵� �I��:�2��[k���O82ǧk\%m]��v�bi��N��i0�cb(@ ���jڕs�^˥Q#"�i�m�.��Ƴ�:�d�8&I&��s�ں��̻����r�v�q3iu�͹�`-��W��:f��ܳ.�A�E�[j���ڳ��k6��a j�6q!:���$��n�vݝ����KN�F�v��h(K��h�%���1k��qN�� ]a��«Ɩ�Ge�v]�,]s �����s۞�;g=m�5o#�]�Gu7NN5�Խ�r ��4y5�1M�*�ݪ�n�Y.��u�/mض��yv�
�,T�v�j���]��K��m��Y��YX$ź�Ɗ8	�Ukn�*Z�[m��)��l�����Y�$-��@l��W+�mуDŀ*��,��aWm�y�C�:ͧ�m��lQ{+xł����C��)��l[[^��v-�-�8Һ�-��gZ��m'a�6b]��Yуs�(5m�U�d�[:SZݐݱ��o:�ܨK��ݬ�w-�V��m�1��[eN�,���z9.��M`�c;emI8�U/r��<U��5����O}*[����fݺ)����g�v��[WW6�`b�gH��Ȼ_�˞v�s�1[W0��u�A$�ڑ�U%�`-"�Vb���l�hїv�kb�U��Tp���ݺ3���)�[G[A��.�.�	�%�L���J���i��q����]�(pc��Um���%���T��ʡ�v��	eN��������6��YJ��)�Bm���!�X�������f���l��r\��&�^6ۍ�K��ko�I4i�Fmcם+v�6[96��:$��t�.Wu�S-�WZ��Ӟ.��m �]mR�5����+*��N��N۹VΒX�.��ۮ������[m�k�R��W/'Slv���������3���J�	���p`�]�;�mm:I�[{s�T�[v�-�z�ՖI����a:���h�k�v~���Utљ^e�ʵ�YgO�{��������y�TD^A��y�:������|�"Dv|UJ���J#6��O�Ҫd#6E��V+ @�`@�h@k�	�L
�����% �^E�މ��)�_( @�'�%�j�B��8��(p�&��Q�bO&�l@�E���}S� z�����z��z&��}@ 6�2(�B�V �H��Px�F,�6���� �H�	�4=P�=Y�J1!;z��+� Sެ H@�"N�0XB ��E�j����`��h���z��x!�N�������z�ᰋ�N(ld`H��b�a �j
��W�⇢>�A��	� ��↍�:��M	'�у�4' � C��u��P;#D�H����<�OEC�y�����;W�1�ǡ��R)p6.���_�B&�B: �P=ؘ(S������= ��b!1uBhPȌ��v"G� �"������=^	�iUS�"���7�QEa��S�8#�GK�j��GO�6��Q0*�*x�D�(�(p��"�`�R�� ` h<S��*�ы�HF��`�$A����0��|OX 1"� �ꣴN@O}
 ���6 8��	,H����	@{�51�@�,  <\4����@ �A�0^ qiriCÁ��"��Fm@�(z��	�CpAS���`I�%���I!B%��F6++Im���IFZ���,$J�J2�imh�1@�i(��`H(����*� ��HB2H@�$!$qE���P��I,D�A�`��\ h��'�$!�I&�H�P��ƶ�+�b���)�<6��C��z�E�}�� ",`2O�!�@}- C�	Q�R
� � 8!@�dS(*Tj�q	UȄP .@�0��j�%�X�R�BA+ E���(!�(A$P$<�u�kZִh�$ 9�Ü  ��m�m��-�Hӄ��h +� �f^�:�:�������f.4
�D�%��/[9��&gi��N�e��ͷR ����ɴ�<l<�8|���p�s����Nw=c^����XT�kuŰb���������a�tb������\�!.���f=zc��]kl�ܷ�	{o[m�W5�2�P[�[C��B�hwY�{m{K[�[;:�7j7k�b��$�����	�M��s���`��J/]c��*v;q�/��ɺ��e9�zI:� �ݍB�g[��	U��[�e�h��nzYu��v�-��k�u�/�g��5#�j3��p�m��nђ&��r���u����jηNzh�;���v��{�z�0-g�.1c��oOk=*�sD1��\$�����sʄ��l^��n:z����ɶ7k%�:����[:'D�k/D.��n�۵9n�<7W&<V<ɓx����s�VU��U��=��r�Ki���1#�!��L��Z���s�.X������cL6Z�����kZ&� X��Y��:'J�V]ɽӒ/I�1פ��Ae�f��j����ud��۞��سc�ڍ�n.u@�Z��;v�(˹n�z5'@^��#��8�9�5X'�u�m!�)���՞[�^A+yi�ɜ�y���㇔vj��VЭ�'���M��u ںƷOI�{u3�fvַ ��m�2�;�C��pr�C8�ҽО�ͭ��ח�N�ڎ�3��Mc���\���Dӹ��9�m;������O>mW'Z�\]mE��T�lx���t��`���!�����X����m�6��띌��InN���n�����S����-vi^]C{Onͷ71��A˛�˧W��G*�Xܻ��vi	箴82V�ӵ��c#l�.M�	F��{�_�w����� �T� ?�҉�
���B=`�����D<P��Q�)��Q�NTGQN�Өx$��(#��շ<Ըfk7.�[����q*]�Nb�i�3r���Xب�W<�=Yۅ�;z��݊��nh6{unV �+<W�8�'h����cg�
Ѹ�퇳�1یs<M��;��6p;��p��봜P��F�bL���1���{n�u��uӍm譓;W����9������kq�uv��;vݸ����A�t<���mv��(uM��s��e�2Yn\2�<-uP�Eǘ/��	ⅺ#�����_�so��w�=�E {2$��m���뼚�uǡ;�%m�������|�#S� /��`b��;�V�J�8���ݕ /��`b��8�5��"aC$���)V�͖.��3]���P�b���A$M2'%����`��;:� ^fՁ�P�Ϗ��?����U�*s�;;8t��X���<m�<��c�k��%7#T�P):�I%*���zXݕ ��q�����v�Q9p���k[�w����pT!�n�%��E��>����s��������,�z��lI���iՁՙ�����g��H������T8WhKt�L�PN;s��9����l���]y����$�t�Q��r; �n����\�;����~ww��ǟ��{]��9�vhӨR5�K�0Ǻ�)����c�_\�ۖ����L�n>���;����k�8���f
��)�>JU����`b��8�lΥ_%��])m�UN�ә��9��M���fD%H�	���RD�
"�*�؊����qn�8�Z:Ф�TRJU�����`ovT�{��ν�`n���R�7���P]�;:�U��y���Z����-�q6ԩ��:�Նv��@o9���=��v���չ�w5�bZ���1�}6��;�;����T��r�i�@�sS`nOs�Ȉ�M��������{���x�T�j��M��9�uXݕ}T�Vf�q���4��R��q���ʀqw���y��܏��;�Q<W�����s��D�)�>JU�ՙ���d�����`f����X���u�jx�v�Ě����اj�=lN�7vi�|��n;=�4�JQ8���f��`qf�3v��	E�ǻ�`v�/�T	ʤTʦ9�����`f�{���<�`nf���Ȝ���G����\�;=_U%����;���;�x��pnQm5
�Y2gȼؠ/#5�켚�%H]2�X\��d
�q�ǚ�.�v~7eH�q@k2�Lμ�_2P����������L�I�Ʃ�K��\r�{�0�[�m�����<�o����y���;.v1��Hz��\L�nvh]l�¦�	;h�V�Z��۵��=�5�<ps�M8����|��0����r�ל�f�zƽW����ܝeӧU�d��:�!�GV͹5�L5��oYFsu����<lC�ٳIj6ܨ�wZ�v���o!mٌv.�ʱ덶���w�篗�ut�Nwj*9*�юu��&t��sq݌ãhX�j!���h�N26�rE$q`=�K7e@:��vq� Ӹ#dFDT�I`f����3^�Xw6X�EZ��ʑ4��:���;�5Xw6X�*y]S)����(�I%���f�����7vT�s�޼�h��u*$ȅ"��6X�*k���ݝ�`}�%����2�T�mM5.���Q�4�����U>�ף;����u��g�,�eq�NH������f;1痫ꪪ� 37��̠{����m��������7�T�ºtBL�+�"�ID/�%k'&��y�M��ԫ~H��i%��l�T�$���{����k�7vT�3��+t"�j(7#��K�jI�=������
��]�����Ī8��#�[������Ws��޵�qҊs5Ҕ�YN i�T�ZzB��ѡ��]̮���d�INMR��hu��:J�{�n����k��*�{u6�R������v���/3in�%7�^���S*&JTܔ�T�sw�wt��$�>P�/�?Ͼ�6{�����֮R�N��MTծ3v���q���Y�=�9��Nf\�J�{�f���޵�җ�����@�l�U�̛���v����_�gY�u�zm�x4rD`�ҥt*P��Q*����n����u���w��]2�h� �"Pr�����76���Vz�5�����F��"Hr�R]{|�w2����ͺ�`�Zu(ST�f�]E$_ou�7�csw�
#�$"0A<�d�f x�vT�J��]�9�{�Ke�֤^34��d6��/3~[{	M��ד�~l�����:�;s�7ltdބ��f0��iήx)�!���:D��TI��#�;��[�uS;�u�w_��k6�N�E"tܒ9K=��3-u���-2���Wldb%E*u32��W��kL�����Δ�bƇ��%Sj�*�֙�1���]�)Vf�2�h� �"Pr�q���ۭ�s.��w��_`�����H��Q!�N��53VX��A1����y*O1���t3�&�n��<�z�ɹ�s�[p�ӛa=��9��6�&���x�h��s�ŷW�8;���p\�ڑ������Hf�Bv���p���a�n$�/%��ƙ�G���N(U�Wcb6#K����%���s];׶��Tf��v��.�"��H�����3�jn��s�����l�^=�뻻ݹ>��;E��Jvn���m�g�f����'k2J���q��]1��������4���/�e+�ݵ�}�����WJu(SU2梜����ZgtǷ{�vs��9��_9D�]a���37n��)^f�͓�����SrR*�cs{�vk���e��w���"��)��K��B\ɗ�y�,/v�y����@D;���D�l�۴�!�vyM�N�-�v�(�NIG��U�9T�ҪDԓ.\����Zgt���|�^_oҖ�F��d�mTUZ�>��Ixb�)����1! |�)�eI�lo�K}��_��x���.�U7R�K�����]�)V{6֙�1��G$��SA.�U5k��*�f��;�/sz׳uJn�C�HӔӪ�����s;�u��Uﳻ����>D�}!*6�Ēi����졨�9�g�=i"��e	�ݪx�`sq��i�����ۭ�f]gq��R�ԉ������yZ̙������J�nF��o�"��)��$�^�:��̷����za �XÝ5���5-���B0�Y�����o>�(fa-i0�5�H@�2�ܲ�4p�KR�$yU�Ry��iʑP�^Y0! (�K���,,B�4�5�2IBa	|����͢l�*2.C|�0�E.����<䆵��!@��<���@�ɵ$$1t`xp�ER���(�5h�!ia눭�H75{5Jj�5�`���Ȅ��72�%޸��&!� ��2]9e���!�8h7�f@�Lq��fcmā%~0LL"���$�!	��}�v���H��4
�Q ��a�	wjP��rM���S@��<�LMzA6�y��ɘ��^���$��H;�	 ���{ ���i>$᠁�l�4_P"P���(]�bowt���8Lю�-d�K8rh��bf��c�D�*]x��0���4�Hi.D&�
�{���$WR�ܺ�.�o�a54T�&��޻r1�w�G������׎�xV1�m���p%&�~xI>F�!!6�g�sa����.��O^��> H慇�z��z��x� ������"�b#j���D=( ��"aAR�z �U|���#�D��˿���;�����t��Է.�\�J�;�i����k�(�	/��K1N�)��PUkL��73z�gMT�f]z�����v�i*��M�/�t����6�o6��XR�O g��]��P=n:�Se�yP�0�w�K=��U��/��3�1�g�t��8J�9u�󭢹�ݾQ�{ͮ�wR��&���/)�y�w&f%C�|]�u,/v��e,�BS��1�Q2/:�Zgt�{;�vt�$�("����@���2�0�a�GJ� x�M�wD�K���R���wPJ��v�~�ߕ�L���K���]�x����x2w�P�s�- ;=�نۓp�2�sz�G�t?s}'X<���Ch�TBD�	'+s]U�w.���]~3��]{ޠN�I�����*��o�M3�gs��ܯg���h�XkN�Q'.���o}���se/{sk1n�D��0���~��Y�����½3"֕2��&��m��I&^���yi�Щ"�{��2�3��g@���_
��^]l�p��Su�I2k����R�)����y�ݻ��綦���j탗c� {d��w�/]IɐN�d���#�YuJ��읓h�q{t;k0X-��k���f�&w���vz�t��:�I�sU����'mںM�b���:#�rX�X���w��H��L���6��vUn���۝I�<v'�b��8W�Q�k�ƌu�L�.h�/�����rd�]���!�Yz����{vEJ��Gy���Z�/b�T�6Ԥ�R�RF���������֙�F���i|ͷ��x�� �N�d^$y��dn�k���u|��R>�/)e�-��%�6��S��7�v��I���^�y���o�"!H�7!$�U��}y���u�]RFz�ifj���������G�y�����-�ޥ���$+�꿖*��uX��rl#ۭ����ȋ���<T�u�r.�[��֫����[��{���������B���n�|��܅$��K�us3X�<�����~��U-�2��0�ɫv�����$̫��<<?4����4�z3
�ٔ��������빾")�!�n{꡹���n{��a{3e���Z�3fl�X^d�C�Q2135�ٛ-I��^m2�fl%W��M�~�����?��z��:�S������[:��N\LtZ���-�Gn���y;ݾ���r3.�	%�e�5�o|�6�9~̟������ϩ#����H�RU���U�M���Xw}_(K�3����!�s�/]	�ۑ����+���`o��{ߵɤ>H"���@!J��V*�2�jذ����G��T}Tҏn{��ܓ����n�=�t�T�J29,?v���U=��8{}j��Y��2L��ٓ@y�n�L̑���3@{2p�]��C&f[�����F;���@u�N�8r��u2ЦdO<1�9�Z�6�k4�ݵ��E�q�������{����j~������q{��@��f�Fn��fI%�gJ�u�hrGu/*"QP���&d��2d�!��M��F��*_��Ԑw�^��N@Q��K �͚2/~wfI;�� ̼��-kQ���J�����^��+�F�Ҥ�w��[�A"H��CڃC �?/�'����o�krO=��3�H�#r+7e@7��S��Ӡ�zX�5_�H�[�ο��%�RT*:Y��B]�[��rhӝ�K���ns���ܛ�]77����E+�M�&ԍ��_���g�#7},y���K}����*�I1(�L�P��k��2�fMwF��-�`j��{��I[��*�
5ڜ���T��f��6nң�I/�fQ�������x��M_Ҝ
�)�$��Ji�;��yy�4jOə�:feռ�����S��(xT���2I2^I�Fot��.���Ϻ�
$�zC��3NT��)R��ɘ%wv1g�6x��&��ls \Hmu��FxCud��1�\��,��r���z�t7��u�r�m��c��ٮ�v�����{n��ݵ�d8�.�ct�3&���9�=y�(�6��.��şa�����-̻�B�rJŷ;^Eˣizcji4��B�>��*�Fj�wI�U[=o^�P9P�Ij������2�&��M0SL�W�s:�&��H��\�auɽ�Z�͍�{��??}،@��8�������7ˀo�gAO� �$��߳�r�����]�̘��"���v3^�	7&I(�z4�5�6(��;���_2ffw.�͙�Iu2�e��`y$�������g(Q���s�����{�`nz�^�$�Fґ�2�̓�&P�3GOoE f�Mɓ��f���� ���jM����}m��[a�KA33@��@jfIn�k�li ��{UT�����t�(�ERR)6��Mm���Ks�ݗ���U��ؗhnv�߃��{�׾`�PI�NN�=��}T����������:I��3f��7\�)�D�"MK�]�=�vkhH��R�$l!�Qz��I��v<��W� �Z&Z!��a�ik Â��H�0f�;d��Di�H�a�Q�jWh ��b �������$��<�����[��^��+�W�Wԑ���tTe5R���2w�͚ �͚9rd�DwF���o�{��@�nӉ�@Q��K߾�I�33��t�����l�҂�2fw�͖���Q�CnF���%˜�{�92K��m���2d���٠���X7����%L�⤔ct���6�d{B^����rqs�F��?_����>�~��q�٢"%�li ~��]��32_8n��7<��&��$hL����Mə(��ޚ�7����'Y3's3T*�$����Xn�X�5X�_ь��!@�y�Lk`0�hG����`���Ǔ2d�$Ι�{��D�{w&�/�O�k-�ն�շ5��������rN�i ~���d�=�f��n�
)�=&����J��!BI�oW�ǽ�7^j�74�AnTB�7P�%%v�9�f�s���=R9�i��d^�EZu}������_�**2���Bu�{},.�{�OU}UU��� 3�v��#�(�����S���2Q�Δ�ʐ/ޛ/~����3לm:R5Pdq��N��%I�$��2d�72t�-�z(����qT����,=_W���7�P�,<ߦ�TB�D@�� "9��	�J"41BR�vk�tbC
 ���Dv�	+�Lɳ�e|P����`&b!�P˜(dܙ�.l�������PVSM �I�ۑ��H
����=��3��qvݷ,���;��W�w��}���ȵå%4x}�M���Ł�ԾI%û�K �IyJn�HJF܊���ҵ�L�ܻ�R��
n�
ԒI���'N�t�P�H�,�ʀg{0�RI-J!�'JogJ�fO�0)��ʠ�e̙�;w�(ݞ(�N�d�$���~R������C�)y����2I.���{��̭,����DG�� �X��&�)��D��,d���R2!'��fɳE�k<�&�<H$��&$1�iF���-��[Zm��"���|��� �`MY�`DـL%l�� D���Q�J�^�<���,��@�iuj��d��!����Ǿ�=CF��4��$i$k6�I�Ǉ6xh�0�ѱ���_yAa`R�_i���I�y�����>/!#��7Z\�.�H�'��ș	 B#a���u֧^zG[^kXhyFej-�ïC	���w3�abk�&����ݐ$a΄���l.����ް�礟C�Ϧ� ඎ 9�Ü@�  ��mj�����_���_��m�VWv`�6݃m��\���.�������1,n��1�Yu�7�.�6 �t	ʹI���囲Ot��i��!]Vy�M����my�L0�tF��[�ʆ9�A��ۥ݋r7
ڇ>7R&�9�+��m[RO��݋��s�\Q�]n_F+�,���{���r���;�y�k]hr�[n]�N�zI+ȩos��+M�,ٳ)�����إ�����f}om��1ڳϯk��(����vz�y:u-���x帮�ǵ��+��u�s��]܏l��۷`����E9�yvɲ��6v�$8�;h䱣������\3�o8�ڌj�\��T����М�4�g��t[<m(s���{x��=vv�3S�ێ�@�㵾{t�k����5���\Nɲܽ�nHu��[I�f�`�Y�V��V�N��e�rc��L�mt��ݦw�Y��uq������mulp�bmvdg��)�c]-�&R��e���Aln��H؇�]�`L]lDs�	�����g�F�����0=bM+ոr}'��nS��x���s�mֆ��ֳuz2�un��
tsۤ���m!�8:8V�!G]z�FY��V�zN����2��';k��r^��.Ÿ�t�5ۣ�q�$�6���v)$�h@�J��	XӴ���.GwMv8��N�R��p׮��:��N��۶�AƲ:��[v�f��f��;<�,��:�7`�-���W^^�N�t�99�UJܜ�*�i�It骺�q�l�Λ׮N���v̷�����T-Tv��V4x���[�Iu��]8��&7P��\t����l�j�����Ǣ���k���9[	�	o<GU8�zɸи4Nخ��M�=�:nݮ�]����m2����w$�"�<E��)��؋�'L�,��n����������w����ώ�9��U4��AH�l<Aq��P�"�
	DC_� h�E��t���:
�A�
s:O6j���A�d�wa��R��r6��� �ɝt�#mɛ[������[�peg����m�-�J�,�^t�*��V��ҝt; h�j@{����9�M�l�x�v��#K����P�ۅ��a��u�j��4��}�pc%��q��f&��:��r���9vY��poT5�4i��9��jr݃s<�3aA�h�Ŵ�W0�rLԺ�5�
��p�t~�{eg�1�d<j�2FO�܊��:pv���gW<�T��{��n�u<U���~������T�~�٩�%��N��>k��0(���ffbJ�S�	���L�2wl�@{vx�3.p�I2N�n��C��T)��xT�N��s��f\��h��(Ε ]�n��eK�
f$�ē2vV��N���R��|�r��񴗔���4�`n�ԙ2�C2fW���ܝ(��
�����m�ˉ�{k��c�n���!f�g��u,��oO�P1������1nn��[����.�T����@}�8srd�z{g��;�$:�`�R�˜+�`��A�	$�d
�@bA��`�*�
I	c��T�l`2 H���G�D�U����������(��<�rLɢ-�T2��C�H�%o��@_�p�Y�Iy�#3f��,�CG�7$n�Q9,=�32O��������ejffM��,Z�~Q�RG"jE`n��IBKwo� v��`{����UHL����D6ڒ����v1˸9=�*���]��}��o��UUQv�6F:���pݝ(�y4���&K�$�+fW!�Ҡ��_��@��d#��gse��d�'s��@nl����X��&w5�ͤ��7P"RrX������������;_�*��{�M�'��Mx^𞘉%��^��L��&ff���H�:P��h>Z�34f֒���nfh�R:T�X�J��Т=͹�3ޞ,͕ κ�|��hƎ���y��mM�xp�<�D���8�vۙ�q�a�n;���q]�ӎP��7!�5f��ݚX�+��}Uh;�4�76�ܑ����`gvi~����o�@;�4�3�<��U}UI�{�8�"H�H�`nl����F���2Q��=���~�)��
b$��̙Fv��{�@_�p�������xJS�C�`@=<4�b(�%�wʀv̦�IEM�w�@s&L�$�6�}ǀ��R�����h�ö�B�)JT_*pu#(T�K��=��H鋀�H�6��!�X��{��'ܿ;��SuM����WŁ�Ԩܭ>J}b����|RN��8��`flSərd� ��Ҁ���/.p�I3��{�ҩL��D���l�`qfk��UT��g�wҠ8�>i�(NP�%�d��L���z7'J�%Hk3=�^���ÃT��7Pdq��4�9�d����w�����w�@E4B@���!�ɪY\��j�X�r�����u�·Olm�*�@��uD���7Kwkțoi.{fi/��G��'�V�L�P�)�ܬ�,m�J�Fmo=�#�����;��K� �u/tv�f\�bu�'-n`�G]g��ݺޞ�u�1��ެ���M��Cn�ν�-Rn�I�y�ݺ�uuq�����Um�mĺ��~�v~�>���3m�ww{�]�=����)ͱ��]L=��n�g�i_Gld���r}��`���s�k��q�wڛ��*f$�;�T����@}q����ܛ��<P�E'xr&aC� /.p�I��Fk��:Py*y$�f,c
t$�%)��u��K=�v��zT}�Ł���H�MT)�V�O���{����I��s^���`O����$Ĕ�%H�%̔g�Ӡj�~vnM,�%ڦ��Z��xۡ�]�N4m=��������,�2�����)r���JC"jD�p}��Ws]�ys��e�{����Z&%����k[�y|���A�1 	�}6��L�&e_=>(wJ���5�3%�W�ٞ�_�Q�M��8�V���XݕUW���`b��;ַ[i�$��q���}_R�z� wse�޼���h�︠7�8���D��D+ �ޫ�-��v�W>�@}��U���WF�[�Zvu9^�<�Y��m*-�R�u�r.�no���|������;��U^v{�`nuq`c�B�����V�#i!�j�AH��9�4��~��Q?s��l��_=jd���xE�T�M)�4X����6��H"�"Ec�
U�n4��a�H��a�s�������s�~Vo������N�*1�m�T�'{�٠.�5��'
nJ2{�@=�����8n9%�޼��W�����-�^@>��hI+�SƼ��6�Xo&�s�vH{cs�������Z���4]m��$Ppb�ԩR.���`qn���'��� �~�3�&܊������`qn�����f鹿n祁��¹$̹�(�{�tS�$&ü= f�M {ٓF�fw�l�@y�^@����`m�n�(��a�	7���`g}_$��n���~@5��|��~~�yV��z���	9,f�,���`c����?!([�ቿɎ?V@6���b�;��6�[��g��y�tmest�E~��\-�unD�Jq8t_�(ޏ[���:�8{6t�=����J���rFՁ�y����g�,溜����&nf���Z^"bB������>��(�f���y�3^���ߞ5M�ԩ)�%���|�������+ �s���G����@�FGE����B��ޟ n��`{z��^�;��w���_��u��p�<-k�_��q������Յۯi��ilC�q{t�N���B�F�K���܊��8v�zI�{�4�[���'ŋB�X�}Y�/f�aS����9��#�E	���:�x�nm�ź���&-O 4�� �˞�絷>��v�(Ƌc�i6���3�E���5�4V�m�b3�OCV����,�q�tr���߃�F��n�s5�0��&���MK�j�8�׵'�q-�d��n��7n1�*�o��h>/�t�Ҏ�I��?~v�����O}����� ̭�&�!4��D�v�^�;6�$�fΔ���?�q_��;��V�C��Ј$�X�OV���.��vs}u`w4�!ҹ�#��y��Rd�� y��(�{J��$�.L�/{�(}�OCJy�P�31@y��(d�z�~_��Ҁ��@����m8��1�S�Jt�		 	�Bn0������J�{1'%��~w����f�������Ձ��Ł��!B�a�����z�)��"��J�3�4�_��ʋ!$�6��k#$!�k�`FI��(o ,c�$��El� �M�g!�7l�l��Z�"�0�a@�A魪��2L�9���@��Ƞ>�e*�ɒw.��&㔉)R�p�:��ŝ�g�d��h���T�Ofȡ���S-˰�����`f�Z�7:���$�O|���*��JJn�lg�j��d����>k�=���l;��#t�]!�)�,��`ۦO!�δ	%�h[r=��u)�o�U)u)���Ј$�$������<��߮9�䗠/7�P�����9�HXY�ŝ�`s��T�'
�K�����Ҟ �$���"����>��*%��a!$Cz,T"���ҵ"�h�� ��ܓ!�3�����ֹJ�r� ���T�EB�DK�+j�"�gpӄ�������t��<HE��F���o����$�àfyD�EO�SN�v�!$����BB<�!6d6z���1%O��OO|=�-�&l�;��&Ed���o��=��d�:I�Q  ڦ�2�%d$�Y!_Mx!���%ަ�KG�$.��L]SD�%<�	'��M;��"@�@!hIxk%�a0A��N��j��6#%Z<�oY���"j%�8�ܦ�5"�q�d���A�&��$B!I%CE(�e� kC�1�I���>D�
P���������6�6��_@����*{�>�t��Av�PZ���Et��1OW��h6('��M}�דrOo����>��Dp �r;���r��OVj�qgq�ǋce&JqB7%Xך�c�+�s]��箬�{��w�����9qض�M�uuZ��Պ�g׷gxf纇LQ��I��kv6�ݡ����?޸�>��.I����������B�:�86S��I��y���oZ�=���{ξ��X�
�&�-�Q2�/@z�iP�^=̹�1��@��yX�k)���Ј$�$��y��y}�ԓ|�}���'bň� U}U���l�X�ҧJ�n��F�v=�@}ξ<o}j�̝�`~Gw��q_���,�����p��<����h��@������T�K�l*T!�����?;�u`g^j�b�(�-ߢm�8����箬��VVj�^va~��;�<�E&JqB7%X��z�x�jmf��d�@^nR�<����^T�0*`x����.e;� {2t�9��u`sj�7p+]Z)�I���\^=ɓ%�y���/cy�=��I��r�_�w[�᫫���f���<^�3��뭷�����M՝���8�.G��-�˞���=q1nX�b78��&i���+�Gt�{�pY+N�{s
 �di�?��cpG�LއY\�u�i�x$kwd�zZs��+h�%gA�����5�n�;nۏ�C�W�672��u��ħT��ո�����
�n#��.2�=W$�抆
��sW.d�5fC6��5�N��esM:�8���ځ�Sv�<��N6
�7}��I!�JS�H����Ձ�y����P��+Wk)�e5�"	)I*��<�~���f-�w^�X�m��#=��St�F�Hڍ�`b�(�����jQ�Ԩ��z�ȗ"T�K��ڰ9�5X�mՁ�y���,{� 7�QTG)"�9��Ձ���.�|���V��,�)2�#��gsܺ{e�k�HrbI񃎲u�:����������!��R(H���U�՚���^� �o��+=�$R�#*9sWrO/���G8Cqj?��p�q,0HB1><^C��̾���:�iP\^=�l�( ��N4�j��<�`s��Vz����5�΀��j�73 �M7T�1rK��ʀΞ������Vk�_/#Қ�R�r�c�VVj�__qX�mՁ�؞��n�e9ʫ��t�w:���Z�óts��W]������s~y�ez��:$mF����}}�`s��UWw^�X���	�>cR86�c�v�zՁ��`c�u�$�S!���M�#�#���۫��U����"W�>:v"b������ԇ���V1皉&�q�(H���]��y����>��O7���寧��H�J�N+�5@=�}U\ɚ�s}u`sj�9�#��L�J�QǮ��,�rv�vs�N��ѓXL��Q��j���[����i�Ձ�y���sn�c�_���32Jҹ}�5g�)ǈ�DJywT�f���D(M���;_|���v��y�*�EC%8�Xǚ���G��o�;����X�19���6�qXz�����Pc�V{���	#2D�bB `�� �X���l�(�8���9�5XBQ�.���gO|�}΀�J�����TsY���pۋ�/l�f_\\��]�v]����n�U}.
S�m�H)"����;�����"""-��w���=��@�N2E	�`sj�}�Wﾦ�_�(�3^����W&fd�� 3�y�S�1B� �V�~P��+���V1�w��'h�i5au��}��+�v�����rff�'y�W���i�NR�H��?]X�������ԓ~g���>P�x1	�<H6:4U%C：��3WYa%�����cv&��z�x�&�]�^�_V[��k�i������@���7ks�:�Z ��7٥�Yq)��ֻ�uE�+,�R�/i&�گ	�Y�����[ʅ�6p�m�n�Cg����E#�,�9���[�[�T�wQ�`/ ��޸�i�(l�6=�x���Ƃ�`�
\��zӹ�P	��G1Z�����.z[nD ��	� �9f�s.��L�3p�a�1�����8�ӵ=s�U���#]m�����"ԥ�"����������P��+�ͺ�;���葵����S�$sj�37�V1��}���N�R*��Ձ�{�`w��V1��u@�Y�G���׻��P����1�?�r�n��~~��@i'"��J�3j�:�T�&{�u`ecOU4%I�R%.����ƶ�3��Nv�-rW�Mgd��7�����[��r���HJC��*A�t]����٥����+���7^�X�OP�d�8�Q�ܓ��7�	 `O�8,C�z�r}˫���`uwu��#sǕ
�MF�R�m������̚Y���K{���<X:�R�Њ�FG*����Ҁ��ؠ>̜(-���Ҡ>��܉:$n8�X]�v��_���]X�۫6��]8����P)Pݨ���ml=b{
�q1kv��m�-N�y�z�Yw8A���͚X��Ձ�ݺ�:���:,��6@d�V{�u�3}�{���<�`s^k��9*�f��X��V<�?!@�	%",c��	�2#"؉��1�W�W�ߕ����)	HqХJ�2�9���b���נ=��T�ٻ�7����*|�Hq�`wj�?}��r�w޺��vX��7�	��Q�wmE�&�aL,��b6�t�8i�q����j]+"mGIJQ� ����f�ՀfwU��;�����DQMS�S*���)W7%i����1�z(z�����HV�I�#q�*�9��`y��(�.J#3z���J���<8�[�I$���,~�;3}u`gwlܚ ��,�؃@�1�]D�����(��w���$�E�m�!���sn�W�~������wt�fExc��8���m�۲1�v��k1r��l��l�n��Gn�{�ӑҀD�ܒU����XwvX]�~���z��7W���8�R�LL� �fMr\� ���7{�P��������E�8�JC�9,���w�J�L�w�J�/wf��`#9-�D�J�a��o�ʰ37�V�ݖ��&�M���Qa���
$"&U��j�3{�����3{�X��s��tj���,c���f��X���Z���	"�HJC°��O<�E���B?��7�ڏ���zSn�$C���BD�V���!ͺ�\z���'�
biD�f��㛑�њv��Wa$� �H�0��c���4��Z� �$H =酚%�vF�HȠ h�5_=�!�`�!��5�����$��Sn���*c��t�W)]	�4+Un�A_e��$	 �a��#n� N<���t�ޢ�$�  -����m�`l��ݳ;cg%5F����6�N͕�]��ۭ�_D���m֭7&k�����l���7m��mV����5����:X��Ӷ�f,�[�'h��`����tu�����\��9���Fs۵���yvb�)�<�S^�-��{wn�,.�'g�{g��<�`e����)A��@v�I�+��m�W��h��SͫR���Y�:8�{Cϲ��kk;�7CG�x:�t����:9ǞnroZ�f��#v�ֻn���^�Zg:�;�����\k�"W�f�H����2]��tM�S��M�	���'=��]tq�ŝ�-���Q[\s�GFu�]]���='��s�G����ζ�o,�.�IHnMֹ��+<͂h�]�X����܋����7N¤���h�ڭ���g"�1���ǩ8�pnz����7-y8�2�]��釗�}ѭ�F�����:���'7bvn�9�!w#���ǻK��я]�7�������r�ǎ������\�M2��<�t/g��e��,i�����7Q�=�F ͧ�m��8^d�P�Jq��0R������y,'�F���[�t�X�L��Ǳ�S�T������مӞ�s��):�5gL�Z��h�7�<l���z�0B݌n���d9�b�76$	�MӃ�6|�F�Y��nݹ4���t�#���xmZI�F'���Y����xrf�7V��fxK!0l�V�+`8��f���Yޞ�����Ѻ���-���"]/B�Q��0�&���)ݪv�ۭ�<�8�[-[��<�҂��X��x�S��]���n2��gNӫp��"��I�:]ʹ��Cv�����굶��1m��y��;��p[��w]�؋V�:�tv���̺.�_��?*���8�莁B��@�U��J"U��|D_D��D�G��M��ODN���l i��{���{��Y�j���K�[r󋳒WN�͈�B���i�o1Qz݇o[&�s��\�Z�S9݃�	���yy5�EHr/;m����:z^J�wn�����p�G�Њ���:�w;7t�մ��Ne�-�i�q��l�ȱ���.�gi�M��%:�9��7\���#��U�癙��nͻ�}\\'�'(+�qrv���O��������Q3g%!s28p�Y&�SVi)n�ݴ�b|�"M�ۉ�����-����'?߽���;-Ƙ���X�ݚ��dP��_�d�.MU���u`g��4'_��4�ܖ�"���R�=��T��Mre̙D��$@d��;}��V{�u`��`qwu���u$L���Ȩ%��E�o� {7f�����3��V��򺎂G�J�J�f�<�l��V�zՁ�:Y�Ϫ��:t������y�]}����v��e\m�K�u����꯮0QZr�!ƈ����=w��z��&M��ݚmkC��KE*N���7zՐ�$�$$��(Ŋ���@�JSZ��iMɓU���ٻ4��Ȭd�Fm6�B**@nJ�9ܚXs���BI�{�M���֬�bn�Sn�Q8X~���}�`uf���۫��|�6�X�y�g��rXfE�$�7~_��Ҁ=y�@{?�����\]�%�\��j���]�7	�ΧĮS�����D��AB" I�H��܊�\�@����2T˙3zB�7��ձ�	Ԅ̺y&eə��\�\ə���vh=���ȮI$�e���]���n��K����__����8��U=Ϯ��nI��_M�n�J�����DNK�WԺ�|�|͊�\�A�'f���#$5�]L�(���<�y&Iz��ٻ4s]��֖m!R�J}���2�lN���lcF�=&��"�9�-)v���=n:1�19��������`qw5���� Ż�`o�E$\������ś��2\�%[��P��޹¹��l�ߑR$�m$�vVo��ՙ���}�|�f�V���3���Q$HL��332[;��N��y�@�A��P�Y#���4B&ȯL�F0�d.����@� l��3rfIOmm�ˣv�	�t�f%&�;ܚXY��.��3]����?�~9�v{Z��������ݡ�����۔�Lj��Q�����>����kv��:/~��.��3]������ĕM	$'�ĢN;����W����l��~vo������v��(���EQ��SS`k��=�\Y�J!7���l��;�Emm��DDG`s�0�>{̊���Pk2f{�͊7C\�U�ӢF�RU�ś����k�:�5��mՀ��Us�U/0�����$�\��{��ĩ;�c��LݬTl���'s�O@%�g[�v�;���]GVy�nQ�ε����N&����9T��w��5�C�ca�]��4�8�[۴e癞�	g79���ngg���]�K͝[3�N����uֹ�^4���8uAr��rmm���A�����U�F�e��v�vף^�ž��&SE�z$8(~|�^]�s6�#�=ۆ1�����F��nֽ��v��8���IQ�$�4DH�q�n>����vU�E�^R���rI7�-��(5���S��	$vVf���l������ؠ>fEkrL�,��N�����f%ݸ��OŁś����][�ՙ���P�>CLJ�4����Ǜ��������v{�u`n��D��J�j$�(�^=��\fl|�6���dP�:��Y܏<ٝ�����Q�]��q�7j[۹x7BR�{J�*XYFO�B�p[������dw&o@nF���\����aN�MT���W�P�	��X����H�$�}�nI�罴��"�32\�(�7��	�L<C�1
)*���ߝ��y�����`ssn�nM�4JR97�ꪯ�UU?m��5{ߝ��ɥ�ś��;�v�c�T���+�3]������.վ�3j��R͑T��LR�7	I6�.ϭ`�s�;�f���iݸ�mu��'��3洆3��h�M�`o^�8�u��5z�� Ż�`nh!J��rD�J�E`qf��|��܌נ�٠3ј����� ���a#r�N5q����Xs6Y�0� Qa@�E"�V
B��[I	�� ���(�(�!D����v�}�`n�5UjR:j|�����RY��`{�XY��.����ҨDEC�Xz/�������=�� z�&���>\�k%����X��t������˂v�v��$W]��G�ٹ�%�ڨ6�V~��u�]�v�͞�� �{�`{_�DD����7��������3�XY���|�ej��6�J�!!$��7���;ܚXY��u��ך�B)*��7%��������`s����X�+e�,H�E1�/B�u����A��C&��ʥST���"��L˓^w�x7zhz����փ��i�uuI�I�8�Hv�7eŮ�%�j^��HȀJ�kCu�,Wh�m���{:����=�־��}��`}��jW�q�Ϝ��,��,w6����dPz�
�e��h��w�K�	z������7]�����;����5jT*-(�5$�a�]{�;�3b�=w�A̟כ�7#v\�)�Q3
!��b���y�nL�w�g�foR�N_{�ܓ�� Edą"������q��6q̝��,9��7np����7Xs��ǠD������q�I��j���Վ���·��iy�$^�9��.�X�۟j���W@���'g:����@Oa�v�X��*q���Z[<����[��Α���N����ւ��u��ծ��	73��c�vs�7Q��4a���a��`��x6�c8{U��=C���{�����������߮�萃�[gl��[&�Bu����{0���CT�WI�tחq��ĈfLX�����*���L�p���P�<�2}$�R8�q��M/���$u�v(=���Ȯfgs/AǕ��L��J�����y�]�vVf��y����b.���c�$I�`qwu�{��޼�A���3v(�F)Z�s�"N;�3]����XY��w&�w�-���DR"	F�Y؏N��mw-d㣗�$����{����>G�� ����������`s�4��l�3MZ TX��4�rU�ś�����IF�	� !�#!		#
@ZVA�!1C���l]� mv��s�|P���z�s3���<)qJ��M��v}����l����o����8��v�ŕ���R$r���,��J���2(92��37��͞�'�JU#�nK�ݺ�?UUWro� ��X�z��P�������6Ɯ�;�絳��a��7(�g�[���[sk���I��z��c_�s�WW��n�9%`_���`w��V�ݟ� �{�V��iUԄtFF�����)W&w^����T�ב@z��i���`��9ܚY��������d�XL�ay2�� ����c��L�U����)�,l3p%.�30J)�A�����Ma!1�3�CNxlBDA�c3ZX�D��-0�L3�B���#ӳ���&qj����0���˿��
k��w|�����/��0�e,�M�E�oy�]��R�����+��t����⛮"D�!&��3�k�K&T̎E�#<�$P��[�%s&�Sc�0�	�!G{@���5H8��¬�i�����~<�d�t��땟H` |� N$,D�.  `���uB�x!��ڼZQ=]Uʱ���8>��_b+�@} �<� 0������gG�t�Z�=�Z��Ш��SUVra��ʀ���=w���fM�-�ptP��x���@y�y7%����o����n�X�E=T�$�@崷c�W;:����%�۰�N�[�-8��m�ۥ��})H�ۊ��n�X;�,��׾�ǾV�յ�6�N$�X�̚�d�N��m*�3^���)W$���O���Gܖ�����^j�9��V���wA
V��!�șT���5�nm* �ٓAml0�����(��BF$�A�$	$I�Ϟ���_V�>��n�J�H�(�H�qX�۫ �we��ͺ�;ך�}�<&���Dl�K\F��k�=$�4��ۮ^77�ۏ/)�:�K�T�m��$���ߥ��޵`fN�=�֬b4��QJ����sn��$f=�;������W�|��5xBAdm���ǚ�޼�G&w���P��T\>`��(�(�q�~��w7ܫ��R��̒�J�I��1l-]$D�	���3]����XY��wv�rO<Y�(�(V�7DcD�R��P*)�A��}󕚸n|z��ˍɊ����V3ֹKG b6'&�s���p��2qqݻpܻcbO�����l7<������c�s�oe���F�7 N[s�pm�d�;lR;�v+���E���3u{i�BY�l{L��us�W;v]j�rWA�k����v���gv��v����9" q=y�zM��ll��vҮ�ff[�\�*"S���o(?�D�]��A�kq�e؍ �n�an�����v��������v{}�N�s�Xx����J���2(��K�2e�y�����+�!�F�SrU�ś���)P��hz�
�\� ��xz�y��GN84�3_���;����UT�f�V�����J�#d�:m�����o}�f�n��{���Q�5�}��Q�,�&���7ˀw'�v�ޫqp4��HZ�TU4V���=`�oH9�;<*^�E�&�/;ƌʢ�9cn6�`s�5X]�v����}\A�������	�J(�X]�w�y�I	ĒI �J! ��"�-F3*�0��	���!��`F�BFI �H02K&��̙r���4�N�ދ�`v��V��jTC$$q�;�,w&�s��ǾVVo���u�R$J���pM�a����soŁ�{�`qfk���s},{��k�!�F�Sn:���ɽ� z�f��\�@yײ�~o�~6�vx�<��]��a�6ڹ�tq��hM�9o66gE����6����?+ �oU���j��N�3@7�9�s���w6XݚX��V�� �s
&4/�>�I`w�4�8��ssjz�7$�A�@ �S�� ;��`f��$��$m�,.� ����;ݚX׺'�(�R��; ��~��������]X]�v3V�)\����b�Q����+�҃���<v���l��{i�B�����ѐm���͖{�u`qw5ʴ�1�,T�"��TL��`gsn����ؠ͉ ��s\�N�^�Q*!�M�VVo��n���33n�w�c�lQ��#q��~ͫwzՆ(�GD�)d&�%7*H�BBd��$!eF0�P�
Z$��HH�,K#!H5�@�ĵ,!-#,��E!"�R�(A��%�%)dm�k-!!R�-#i`YM�����S�z�v0ҷ戝O���9��`r���|��b�2�$L�/�K��ǃF�P2��ͮ6�	n�hǶ��fw;"�9�D�ʪ*"�dt0�����Ձ���P^F�o�^l��?�r�e(Ӎ�Vs]�nk���3���ɹ�nS!�?'x�;�<�v�H�&��g���zlZ�w*r�2�IC̀{7���޵`y���|��L�|��F�J|���nK;���<�zl���/ٵ`dLB��KȈ�

��w�L7ST�r�)�����-ug�W#v�@� [ �R��Q�gv2�v�LhU螗t��{r�v��΄l��N�cc���yb����ZD��'N�Yԩֲqek�8��ݓ-d�À�!�z��w;d���pz�J���-s*�u�uI�	��Ή��[�9[ny���Ÿ�+��I�p/(u<`�8ƺNmPW�;D��37f�h��j�%��}Mʤ���u�L�>nҝ�C��Q���l��r��DnS�V��ߝ�n���37n�w5��:n(�v�q ��h��T��ȮfK�D�+�e�<�P�oMw�J�w���{\��(����rKI�.M))��@|���q �\�9��IRE��F�rJ�8�5��\ ��%��ݺ�3��1��{f<��,u�l�Z^}��mqr;n�	���\ߞ�|�W�I2��'#��� _{����n�,�v�[ި�t�# ��	�|�~���u��D����f�����p㮬T�Ȓ%Q27&���R�>{��9$̾fQnĀ{2总�5R��D��&U�&Qs���=����;�����qZ���'��}� �U_r��}����Ԩ��"��ɛ�,ODA�$�N[�dъn��v�S���P��ږ����`k ���pU$| �論�ݺ�8�������&F�d�S�I���R�L�����Pݕ |�z�'r���J�$J4�U����`svT9��D$�d��jT����q�u T�b�"5L�SiK��@&��M��J�;^I��%�䄚&�d�����@uV�l�$�S䤎��Ի�]@:�����u`qwu��a�Q4�DFB��@y�y�%ənwyx|�=�������l���ܻn]�)�6�h�������s�V�srOf �n,v�M����M���j����;:��l1���Y��ߩ�ԒS�U�������|���R���~ܥZ������y�y�0E(����=�p.w������� �{����h�C�	Q�G`uw77$���f䓞w�ܛ 
�Vq
��!A��-�b�4R�0��2jL�&e�ʽU� ^�'\�A$v3��X;�,;����37m8�DJ:)��6A�+uNv�{\�����'���:{	����y{�M����{;��7:h?f�	}	zC;ﮬU��A�(MR�	�,�����9�۫ �we�#��=ꉧJ"2B"
��b��ٔ��gs׻4�4�-t;�F"��Tm�a��.�ʰ={:P\a!�����b�ū���Hn!�9%X��,c����=�֬"�"$bY7)J&��i�	|�v�d�l�M�dp�Ɯ�����JR�QY�A�-4�|�D@$$n��h�d�D(��hB�@�^��/]��L-����e�d�P����+Zr�iȔ�t6p����#��]C'�'���{w�������a���Č�3$$$d�kT�2P�D��9��I�FH�������R�0�ĉ @���a`��WaI#9��5a MO/�q��s�"���K��D(��s�Ӎ�u�EX�@G�FIi'R�]D4P��|�����	�����!�����+�mی6H�c�lbH�H^��$�!:�{���%ak[b1��y���.�ǆB�l����atvf\�W�C��D?$�<�t[^m,�juy�|�k��BI'��8�\�x\e���B%k�p��P��	P� DH���n�/�f=�\	���P�O�_>dU�3y�$���� I�À$m�m���H m�.�N��$�m� ��ڐ�M��6ڵ:ݎ�t�,�d�G��s�u\�A�g�=�w59��m��F��5����0u���,.�5��:���ܩ��ח۷f��ָ�H�ò�#��`-�A��4>��cW����#maD��jx�;W8�s�x�W(�[�ӭ���+j����t�h}]�\�s僳�������v��� lی�{>r�k`���ͬ���]�8ݻcl��<n�ˀ����\Z�p�n�vu7n��s�O�=�Gg'���q�o+a���s
���s\r,f��nh�'K�7C�n�=��zݏgbs�ݯ[]q�"�j�{v׵�� ���CpN�t��M�׃4��6�ѹ�m%��s��%Rcl��N��V��-���ڵ@ssU�{XIl�ݭ�IwX�l��t�e�e76�,�`��>Φr�C��n
���!����>5Od�v�V�3���hɵ�Cny؜��t;�A��֫]v��H����j97<�A�;F�/L�i:������\B�#[�{r���swY�[huOGi#V4�H;6㵍�
"h[Unf��ۮ���ƴ	�'0�Ǖd&���G�v���:8�������a��۬��-g��b�[��ʚ��=����K�fł�-�( �sgzK���;96������s��wiI���L�E���rJ��ijw ��)��a����Kź�9�!�y�{.;6ºڷNꭐ�@�vn-g��a���4�����ٸ��[�́�ݝJ6�ݷ��b�6;�u�67g۞5�|�`2��f���̩���&s�]&��Md��s�e�'	mmt=�U��,��#m�Z�u�AS����x0�!q�FM�k�ΘM��l��F�\���5 �f=Fs�;Ej]�;S��N�����-��nyiwg��V��gu��~w{����^����]���@@�G����@�G�N���@�C�DD*�N��@}] �x!��x�>k�>�vg6�e����u�8�7M�vR�lNNwm���u�B���<Ih8��%4�%�wkg�ϗg<O5�V{���ɼּ�.�u��vx�3V�t�f^�ֹGh�ia'��a9����:����Ż*�;���4f�7��Ԛc]h�q�ݻ*mkm�mv�hK0�1l�G�%v�tٛ����t����V�jd�W$�1D莆�߽�&���ۋi�Al�[�������Og��K�IE�I4����֖�
�m�F���(��K�/@^t�@f�^��t�:p��Ws]����X��,c�{�;[�6�ICI��={������;�#I޹�m$%V%4�U������= }鲃�Dz�|�u��d��L:yg��(�0�9�&K޺��={�������2ܕ�(�C�C�I-�"�krd+n�f��sH��e�gm�\A����}�}�fns��D3g��fR�>�N������ņ��	*�%Q5����vm>W�S���sr��}7$�������ez����:rJ�9׺�c��va`s��V��(�9DR��/�s&��&���}�iȖ%�bw�w��Kı=���0�\5tk&kY��Kı<���m9ı,? G�����%�bX�w_~�ND�,K���I��%������G��X�1�ۜXPgA�϶n+t���d�D�����.��n��ѷ;X�9ı,O=��ND�,K��]�"X�%��w����DȖ%���iL�8��N2���;��a�a�cZѴ�Kı<�~�6��bX�'�߮�q,K�����ӑ,K��߾��ı<���5sX]e.�u�fӑ,K��;��n%�bX�y���r%��Y���>�S��R���z��D8yȞo��ND�,K����iȖ%��Y��N\�L�4�3%��	����$������Kı=���6��bX�'���fӑ,K�"{��M&�X�%��v}~5$�ֲ�W.��6��bX�'����ӑ,K��>�ٴ�Kı<Mı,K�;�ND��=�������-��^9�y����\s��]��͸3�筻m�ޤ���kJF��:��o�Ԙ^�kFӑ,K��>�ٴ�Kı<Mı,K�;��O"dK��;�T�ᓌ�d�.�w��.�"`r_Z����r%�bX�w_M&��#�2%��~��ӑ,K����p�r%�bX����6��pC*dK�������WF�5��ND�,K���ND�,K�~��iȖ?�"w?}�6��bX�'�k��n%�bX�����Q"��KC��W�&Bd&B������%�b{�w��r%�bX�w_M&�X���@���N�_D�j&��=6��bX�'�I�ŲӚ��5���f�ӑ,K��>�ٴ�Kı<Mı,K�;�ND�,G]�iL�8��N2ݗ�˄�ʕ�ۍ�,7�v�<^7h�������,uT۶��N� #ב������m}����'�=߿��d�Kı=���Kı<���6"X�%��{�ٴ�Kı<���W.Y�Fj�̛ND�,K�~��ӑ,K��߷��r%�bX��}�ND�,K����O����d.��� ʩn�3U4��L��V'����iȖ%�b{���m9��șߵ�i7ı,O}��ND�,Kӧ��Ϝ���kT�f�ӑ,K��=���r%�bX�w_M&�X�%����"X���=��~�ND�,K��[���5��-ֳWY�ͧ"X�%��u��n%�bX~������Ȗ%�b{���6��bX�'���fӑ,K����^����T�]e������݉����w=`��W�8�.��z�k;����VG��v��8WY��"�4q�=Q��F.���A�]�&�N�-c]#i�G\d�5v���P�q�5;Nc��1������0ɧ/+���+P�N��>����vׇ"��נ�����	;]�FMݮ}z�0Z�XȤ��l 9S{5���"Cvt�������_3��<���$M����d��+kegp��s�ݸ�vw<v��"�F�k5:�D�,K��;�p�r%�bX����6��bX�'���f��K��>�*��	��p�NE%Q2K�֍�"X�%�����i�z���,L�~�6��bX�'�k�I��%�by�{�iȟ���2%����ŲӚ��Z��sY���Kı;���6��bX�'�k�I��+bX�y���r%�bX����6��bX�'�}���(*Zt����^!2!2}\T+!X�%����"X�%�����iȖ%�%�߾�ӑ,K���I��k&I��Fj�̛ND�,K�~��ӑ,K������Kı/������bX�'�k�I��%�b~Cߤ�s-���3�[���ɺ��谽���a;{���cujIݎ����[�^���Orx�;����ND�,K���kiȖ%�by��4P�r&D�,O}�xm9ı,ON�f|�ѭkY����ND�,K���ki�m�BI'��@jK���H�~��]�؞ı5潚Mı,K���6��bX�'�wM�"X�%��{nϝ5S4�uUU35W�&Bd&Bϫ��q,K�����ӑ,*Dr&D����6��bX�'s��fӑ,K���6�]�C�/S/�N2q����xm9ı,O���6��bX�'���fӑ,K����n%�bX�v�-IT�ST��L��L��u�m9ı,�=���r%�bX�w]�Mı,K�;�ND�,K��W�.���'l������E�����n�e�'�(͐�6ct��&�ދKn�u��2�e֯Ȗ%�by���m9ı,O;��&�X�%����"X�%��u߮ӑ,K����\��4k)t[�k6��bX�'��f�qRı,O<�xm9ı,O���v��bX�'���fӑ,K�󦏏�d�5���Y��iȖ%�b{��p�r%�bX����v��c ���#�	B~��_h��l:� �zv%����iȖ%�b~�_M&�X�%����T �6��i\/�	��d����r%�bX��}�ND�,Kϵ٤�Kı<���Kı=\�e��)ԕT�i�\/�	��	������bX���o�IȖ%�b{���Kı=��siȖ%�byw�������?K�=b{IO��À2�7]����n�ʼ�Q�9-%��wzŸ���6�M���Kı=����q,K�����ӑ,K���~�ӑ,Kľ�ߵ��d�'8�u^�0�
^f$�_	bX�'}��NB�$O~��M�${�~�БI��Q?��S"X�=>!�&��5�d�Y�ND�,K���ͧ"X�%�}��kiȖ%�by�v�7ı,O|�xm9ı,N�w�Ym�ֳY2��k[ND�,��2&w�ߵ��Kı=��]&�X�%����"X��������}< k7Ț��y6��bX�'�����5�h�R�5�m9ı,K���&�X�%�}��ӑ,K������Kı/�w�m9ı,O>�? ;�]���;\n:�]>����Og��8�Ԏt��0�e�fݷ�����u���w��X�%�{��kiȖ%�b{�w��r%�bX�߻���y"X�%���P���L��Y:|�B	�m��MS��Kı?w��m9ı,K���[ND�,K���q,K���w�j𡐙	��r�ܓ�ULӪ��sE��%�b_~���r%�bX�g{t��bX�'�k��ND�,K��M�"�	���:��MK������5W�+��"{���Mı,K���ӑ,K������K��3�٦_�d�'f�k֠ �%�&bM�"X�%��u��iȖ%�b}����Kı/�w�m9ı,O;��&�X�%����{Y���.S5]�kbarcs��S�j�G1�:�i�nv�gv�^Ʈ���Z1���j7S�<ώ�q �\�Ɨs �9��b⺳�xU����I6k��H�=��u�ew�u�Is�y[��tt��pJ�ly����5u�8�6�9� �W�����/N�z,g��֩�u����L�����ېy��n.1�9m�ʦ�N��Sٹ��e�k-֭��M��;���"g�j�C��1��ݛ'=����
��I�� ��/�V2q���e����Kı/������bX�'�k�A�(NDȖ%�����Kı>;��)m�5��L�sY���Kı/������bX�'�k�I��%�by�۴�Kı=���m9�TȖ'�����d�tj��Zֶ��bX�'����n%�bX�y���9��Dȝ���M�"X�%�{�ߵ��Kı^��y�.J�r"
e���Nk2B2'{��v��bX�'�wM�"X�%�}�ﵴ�Kı/�w4��bX�����(DT�C���p�Bd&Bb{�w��r%�bX~��~��Ȗ%�b_}�Mı,K�5�ݧ"X�{��������s�ݜv�s��y�����S���o[��.s��3p� 5Ts�S��VwkY���D�,K��~�ӑ,Kľ}��n%�bX�����9ı,O~���O�	���:��Q.�r�j�\�\/D�,K��sI�b�r+��T��-L�>�OT7�H�ı<�\��9ı,O=���ND�,K��~�ӑ?"eL�b~�$�w��Y5&��ֵ�ND�,K�����Kı=���m9��dL�~�~�ӑ,Kľ}��n%�bX��Nü��D��L���ӑ,K?"�L���s��r%�bX���~�ӑ,Kľ}��n%�bX��]��r%�bX�=���m�5u����f�ӑ,KĿw�kiȖ%�b_>�i7ı,Nw]��r%�bXd}���m<�bX�'�{�?�o����2��\v.l\���Z��f{EGm��:
���x��_�7&�v국m<�bX�%��٤�Kı9�w�iȖ%�b{���m9ı,K�{�\/�	��>���u"2��nfv��bX�'���]�"X��2'�wM�"X�%�}�~�ӑ,Kľ}ܨV(d&Bd/N����C�USiȖ%�b{�w��r%�bX����m9�*�O7	���^�(0�uJ�j���8��$-V���a�F$��Y$#ZJJ��)�$cm�%ek�K-��ZV[KaB�B4�%	IH�{����W����x��+�W�����D4�Ц������R�۽��5�5�ц��jn��@+���dd	�6GP�	hQ�J��p��L8>!�e�B�Ą1d�F�(JZJZ���]��	�6Ä��=��!��!zV�T���b�#]IXZ�� !B��n��0a�q�<-6���!�omM��+�P��ހd�6�-�@!�f����Z�#C\���l0͐�
R;#%K��sd!�aM��WĚ d���u<�)��,Lv5�4�6�JQk�b�!ZhR�F�-��%,Nx�����Y�ی�~�IB�$���JJ�!
�!�*Ldѭ�'E=AO�M��@��R���'<}@C�WB�@�����)�Z�A��R�"::'�)�8*z��M���"n%�f�q,K��}�siȖ%�bo/�e�B���J�TӚ.�L��L���~�ӑ,Kľ}��n%�bX��{��r%�`'�wM�"X�%��:ϊjjU9U5U.j��L��L����q,K��{��ӑ,K������Kı/����r%�bX����R�k$��-�m�ɷW6�SY5�֓��@ݩoo/�9�0���k�w��'�ı<���9ı,O~���ND�,K�����凑2%�b~��t��bX�'OO��30�55�$�\��r%�bX����6����L�b^���m9ı,O�߮�q,K���nӑ4+�2%����m��ֲ�.fMf�ӑ,Kľw�kiȖ%�b}���7ı,N{���9ı,N���6�!2!2þo�2S(�"�.j��xK��2'�w��Kı<���9ı,N����ND�, ���J1Jr�T�a"2�#��(��S�by������bX�B��;�-�9t�s2��L��N'���]�"X�%��X���~�O"X�%�{�ߵ��Kı>�{t��b'�=�������g�L��Sz�m�5�#�j����.�T��T�Of.+�.�'�l�9�֮ӑ,K�����iȖ%�b_{ߵ��Kı>�{t��bX�'6����	��	����*_ʊ��uT�j�ӑ,K��=�ٴ�? �#���b~��t��bX�'��~ͧ"X�%�����iȟ�*dK��O߬�]I�5u���fӑ,K�����7ı,Ng��m9��D�Dȟ~��ӑ,K��w�ٴ�Kı>�C�!�SD�:�p�Bd&Bd,����Kı;�w��r%�bX���6��bX�'��n�q,K����&ePS�$�57�&Bd&B��."X�%��=�~��O"X�%��;��n%�bX��^��9ı,M)�ސ�aV�*T���N��uϸOw�;��+��a���U�p��yk\K��Nz;n9�g[=�<Y^yr���s�E���,VVd㴼T�nȻ%õ.�]��\m<�`��M���y�g-�u��[�x9�NU�%�������ŵ%����y�X��O"qc�#n�����9v��^��}�j�꼳��vEIܛ+u�f"�s�}�o�y�;۳ֲ�A}�y�/6�%�*ȅ�%*}�S�A5ETԖ�M2�ݎd!zu۶l�u���.q���z���q\��1�����=��Or{�w������Kı>�{t��bX�'<׽�ND�,K�wM�"X�%�}�����L����5U7�&Bd&B�w�A�t9"X�{���9ı,N���6��bX�'��~ͧ"X�%��|�L�*JT9�w�&Bd&Bͮ��9ı,N���6��bX�%��[ND�,K���I��%�bs<���k!f��IsY��ND�,�D����6��bX�%��kiȖ%�b}�4��bX�'=׽�ND�,Kܾ�	�IT�TӚ.�L��L���~�ӑ,K���vi7ı,N{�{v��bX�'~���ND�,K������i�ݷP�T��<[΍f����p>�ls���d@ ���ز=����M�����bX�'��I��%�bs=����Kı;�w��~T/�5ı.n��/�N2q�����C� �,�36��bX�'�߾ͧ!\�1�8*�x�Ȗ'>�|�ND�,K��~�ӑ,K���vi7ı,OWlw�ePS�$�57�&Bd&B�M�"X�%�}�~�ӑ,)��?w_M&�X�%��w�iȖ%�bz{���l�5uunfMf�ӑ,K?2&w�~�ӑ,K���}4��bX�'3��6��bX�'wM�"X�%�|�}g��Yu�u�kiȖ%�b}���7ı,Ng��m9ı,N���6��bX�%�����"X�"{����ď~v��1'��ַh���Z�9d旳������Z�. ��`�ڔ6��j�ND�,K�u��iȖ%�bw����Kı/���l?!�o�5ı?g~�Mı,K��}a٬�֭%�f�v��bX�'{��NC�șĽ�ߵ��Kı/���Mı,K�k��ND�r�D�=����?7Y55�h��f��"X�%�{߿kiȖ%�b^��i7��1��"A�`$� �H�,��`F2$�d��#�I	*A!"Z�##������"y���fӑ,K���p�r%�'�=���c��Si5ٶ�o�ߣܞ�~>���n%�bX�g�}�ND�,K����ӑ,Kľ�ߵ��Kı>읷���,�u35�ND�,K���iȖ%�b�߾��Kı/���m9ı,K�~�&�Sܞ��}���+��X�8ݷ,v���zm&��ǃ\��k�$�N���:6{��)�b�պ2jɬ�q<�bX�'�~��iȖ%�b{����r%�bX����Yșı<�{��r%�bX�;�Ŷ��j����˭ND�,K���fӐ�(șĿw�i7ı,O3߾ͧ"X�%��}�iȟ�Pʙľ�߬�n�3Ya�f���r%�bX����&�X�%���ͧ"X�%��}�iȖ%�b_}���r%�bX��R|e�3-�֭52�ͧ"X�~AbdOu�߳iȖ%�b{���6��bX�%���[ND�,��=a�ϒ�����kc��L���_=�s�]&�X�%�������3Y	r�Zͧ"X�%��~��ӑ,Kľ��kiȖ%�b^��i7ı,Ng��m9ı,Ou>-�ǲ��d�[�Ź;=v��ݰt�A��n-x��+����7���"<�\0�:̺��h���ObX�%�|����r%�bX����Mı,K��{�ND�,K�{��"�	���>�O��&�U3U.j��N%�b_~�4��bX�'3��6��bX�'���ND�,K�����"Y	���>n�T樖�E57�&B�,O3�}�ND�,K�{��"X� 	��/{��m9ı,K�߳I�!2!b�N��*�JJaSSp�%�bX����6��bX�%�����"X�%�}���n%�`~AdL��٦_�d�'j�������Iw���Ѵ�Kı/���m9ı,?*1����ND�,K���kiȖ%�b{�p�r%�bX��CBQ�Q�
O"�1��E`�T���o}��{j�'��s۱1m�;<�pW[��er���n7Tqvb�l���7E���x�k7B�霹����	u�{v���ؑ���BE���yO/0����Ձ'&�ٍ�x��m�h������<t�۞{Ol��i��Ϸ�m­�m]'��[��\���s�C��8�1h�"�L[f�_7GM#�u�^Og�^k�r��q�qw�������������V�y���Β��c(7+�=�K��tά{�`dոf��Xh˭k^�bX�%��&�X�%�y�{��"X�%���8l?��DȖ%�{߿kiȖ%�bt�R|O�̷SZ�je��ND�,K���ki�~H�L�bw�~��Kı/{��m9ı,K��f�q,K��Wș�����MUU��	��	��{�ND�,K���fӑ,Kľ��i7ı,K�;�m9ı,O:}���e��kE35�iȖ%�b{����r%�bX�߾�&�X�%�y�{��"X�%����ӑ,K����̟'TUHT�:���^!2!2߾��bX�%�y�{��"X�%����ӑ,K��=�ٴ�Kı=�R�Ϧ^��u��u�Q��v���\/,�t��<�&�v��ͧs f�iݫ��V��~�r{��ľ{���r%�bX��߸m9ı,Os���ND�,K��٤�Kı<;����f]5r]k6��bX�'���NB!C���x�E
��ND�5����r%�bX����&�X�%��y�siȟ�S"X�}��n\�qֵl�ֵ�6��bX�'���ͧ"X�%�}���n%�bX���6��bX�'���ND�,K���>�2iֵa�k3[ND�,K��٤�Kı=�=�m9ı,O}��6��bX�$��������'8��X�!��&k2��nfӑ,K��{߳iȖ%�b{�~��Kı<��siȖ%�b_~�4��bX�'���7{����Գ��m�U4��r9�J��,��'��qɻ�U3����Td�y���ŵ��~�r{�܉����ӑ,K����ͧ"X�%�}���m6	"{��n	 �t�XL�ֲ�f����ѱ$D�}�q>�bX�߾�&�X�%��y�siȖ%��w��^!2!2��O�uET��5m�m9ı,K��f�q,K��<����KQ��)(z)�8X�D���iȖ#!2���x��L��]�_L�ʊEj�&f�iȖ%�bw=�ٴ�Kı=��p�r%�bX�ϻ����bX�1(��T2q���ej�
���x�ђY�k6��bX�'����"X�%��~����yı,K�߳I��%�bw<�siȖ%�bz~տ�a�����=h�.�G�Һϣ����n5-�q˵r�]���[��~�r{�ܞ����m9ı,K��f�q,K��y��ӑ,K�����iȖ%�bS��9��*i�4��U\/�	��	��f�q,K��y��ӑ,K�����iȖ%�b_�ߵ��O�&TȖ'_�'����]L�52�ͧ"X�%��;��m9ı,O}��6��bX�%���[ND�,K��٤�Kı;�ܜ�$N&�C&���x��L��[���"X�%�}�~�ӑ,Kľ��i7İ?!������ߑ<���[ND�,K�O�s?d5�]LִS3Z6��bX�%��[ND�,K��٤�Kı/=���r%�bX��߸m9ı,O0��}��34D���=g����`ۮ��v��qy�F�䴗Pፑ�\��[o�ߣܞ��'���?-&�X�%�y��ӑ,K�����a�A'�2%�b_~�����bX�'ݓ_�~5��SWD�3Y��Kı/����r%�bX��߸m9ı,K�{����bX�%��I��%�bz�@�|�r攂�����!2!n��6��bX�%���[ND�,K��٤�Kı/=�u��Kı;߾%3393Xj��ֵ�6��bX�%���[ND�,K��٤�Kı/=�u��Kı=��p�r%�bX���8s����ҧUUp�Bd&Bd'�}5�X�%�y�{��"X�%����ӑ,Kľ��kiȖ%�b|m�>��V��Yh��t��L��Ĳ*"��+y4�1�.M���h�M�g±���g�^SY4�V�N���e¦$�9���6f`Je�p�Á���7d�	p��W��R�����4y*�M+M��C~�d��r��1��Q�g=���(�p瑩�'dķ�����)�&�!y��~y���C�oKP��H1 @��`a �$	��,B��-%��B8�|΅���7�MKY�a6�Ƭ0��e,�t����׾n$�&��k-���L��n�l\���w4���%a^5������ffS�K�5���8r���!����'���z�w��0�--�$:>55"R�$a`�z��@�@� ��0Ɩ*E*�j@��w��͇��!X5�ԟ��J�V��ڡ��)I�HU$kH��%�e-$�3.�ǟ�U�M5�R!�@@�2�2�U�I��%Ku	Q���h��<��L�Q(��1Pؚ�:��	M��>�SLs9M��!�V��<S�'�yh�c��&����k�9|�=,��'�C�s^�$qc�iZ[���{�gϟo�	@�� snͰ ,������:�u�� �H����[���6����u�E6
���6�e���+��vI�Ε^�Ј0mY�y4m��u��ť�+�q����l���^ۮZۮ{U���mb�m���ݹ�A�n��=��u	Jnu^`���� �\: ca�����w��<��=�F�.:�n�.ܮe�q�9̳W]Y]n�f�^�$�k�]KWE��6�ɠ�gNn@݌ak�ݱN�.p�X;^���!�K�wl���˫�z5�tQ�b�냓���k�p�^�u��[sb�&�%�sg﹍��Wv��t��ѧ%���޵z���F�qt������rn����td�;ڡ��wG<m���u9��^���r*+���2�od:D�lѸm�x]�+�����O�.��B+�j���ֻ����p�����FJ��b���P�GO!Ӗ�3u���!��g�6`����O)t1��'���Qxz!�>��ȇ�k���n��Ӹ��(���y�T	�jn3v��n]k1�ӷk��<WV�n��E��[��#A���m@� �`��#���@��X�͑�vl�hc�<���n���k��r�xœn�֞d���]��r�3��Z{�u�����G����NK���[b�XN�Hh�2�}��wu{
��un�������Y�:�r���(�\kn#�%�3�nܢ�+�\L�l3�n�e鲯3�ċ��N����р(3-���8N'R��#'&�U��W��&Z
��ֹ���nq:�hY�m"Zyѫ��gr����t��#Ozݎ^8�]����sZI�����u���Ff|��|������۵kU�_�������T�\�[[��}:�SH����}7M״�=�3�����=v��%�Yr�WX�^�n�SNj�6���]je�Y��k3H~T�E�� x�т����@��V�D��h}�{�`��G�A8�:W��S
��rHJ�R�G�|����)�Hn&�����s�R[�ͫ��;\�QV�p��@mu�
���n���Ur�퓪�l<D�/]�s/�^���٭�v�Np6�tq�d���U�CWڸ����[��z�^q<�<<9K8	� �v�X����69'�Z9ۏǮ�&�m�]k��Φ��V{�(���v^ٹ���lc=�틛�P%2l֨�B��	l$�%��0��
�a%J�|�{�p<����'	�=[)���Jmy��d��L�je����Kı/�{����bX�'���ND�,K�����"X�%�}���n%�bX�����d+�j���ֶ��bX�'���ND�,K�����"X�%�}���n%�bX���ɦ_�
��eq���$DI:.e֍�"X�%�{�ߵ��Kı/{�i7��ș�����"X�%���~��Kı;����n��Y�Y�չ�m9ı,K���Mı,i.fl�;�� �f�zڑJ)Ԕ��v�͖�����p�����t�fSiҦ�$C��"�*Un���s���1�nwf���H��{ b��6�;g%��ͺ�fl��p�ܖn�mL��)�33SJ�=��(DB^����ʐ>D��/��I'|�ܓ����U}�y��4�'�"�%NTRI`�p�ܖ3=u`��`g��Q&D:qD��fl�9��V���UUR[�p܌5��A$T�8�=��� �ޫ ����X,oy���^E�+N����76��'	<l����&5�<F�e7J4�)�$�ڒ��͖w� ��u$�|��ͥ@f���rF�dnDܖ��{ꯒwvX��* ��&�&L�Ͱ�}�&\IC���|y�4�{J�ebM�C��f؄�j�
|u{��f����ԉ��0�$�3=u`�l��p��,��J�M+�EێU�w����}Kw��9��`s3�Vc5�6������6��e]rg���C:on8�	��v݇	��:ܺ�7D�ʉ�,3\ �fK��u`�l�3�aY�j!Ӑs��&�7D�Ԩ3zh�"@����i$IS�K��u`��`���2X�-iꊚ��RmIT�3��l�fĀW���M,��D�r&!�:/�qD����Ձ�k4�N527"NKV���`ff�Xs6X�iA��2���u�+vn��h,N\��Ǌ7\٨onG��;YZ 4�J���)�s7e���u`���� ���+0>Sj�i�aRI(��U��4@f�M���^���yIRi��6��`��`b�P�ԑ�ݖn���05`�oё*r��U������X�֬7z�����"MD:q��s7e��ͺ��uX���B� q�xE���u5C�r/Sd�4n��89�yynw����h���Kh�ۤ��U�^���װf�ۅ4.%��nF�z��xB�>F�ı�B��,[\�:ɲodv9-d��ښ:�z�m�6���b�;Yu���{c8����Ů�),YoI���g�峑�f�s9�ۤ�Iv�c��m����e��:�g�UH�1�ݠ�	�5�g�4U}��9��d.���fش��O3�]9�M���`��i)��;1qV�Fg�l�ko��~~w����պ��d�3����P�JM�*�33e���H7�p��,�z����T��kk�%##�F���7�p�2X��Հw3e��mm(�'҉Q�3vX�۫ �f�(J}��@j�@β&e�)UUVfz��;���3u��d�;������kΛ���-�+s!3�')T^=�^�D7M1�I!���m���Xs6Xn�}̖s6��05`ӭ�2$�UU`�5)Bq	lDbP�N�6�fmՀw3e��nDV�$�C�"��י4������٠݉��c)��q�`w3�V�͖�� _s%��ikoQ�$��RU ]�M�$��v(�̚�{J��s�����Nwn7l��L�V�]�v�m�ke8�7C����9�N���'u�ۭrj�m��"@+�s@z�)k$��fl���W�F>�H���9����f�X�4��p���e&�� �$�n��wk�9(P��Ix�Ą~P�L]�}AB�y����I'y�,�m$�n�UM6G*��ɥ�^dH]��jL̞�7�@�C��ɑ')�!`���d�;��VfM,uֶ��П$��
c��$�����sES�v��cb(��e�$\��Nє�]�:��wuX�֬ͮ>�`w�0�da�� �"���{n���W��<X�\ ��K���jԢG�r�fM,7 ��%��ݵ`oKz�:�5)�*i����D$�o��n�X���� ���4�����V�LD�*d �b�l$�*�J����=�'���Jb):�v�͖s6���d��3u�=��?��X�K�s�7F�kl���b�.���E@���^�.���.�)�c�'r��������d��7u��rX���)�c�F�dr�fM,�� _{���oZ��!����K��Jn�ꨰ呂/3j��o֬n��P'�RC�R���`��`s��V;�KU}��%�� ͬ�5����D�ܖ�~�`{6��ޚ �fՁ�a%bB��
T��ii2��U�!L(��}�uNj]�J`KA1�L�/n�}�ŷ���ٷQu����I�QwG��z��r��c�M�rj�':ہ�E/`�rj[(�c�':��^k�zwll�d��m�;m�u̸���"Ba�I�F���,[���W��c��'����_Nv�Mή�w$��S����c&�q5�ށ�7%�v�Ѻ�u^�]��l[n���7e�)��w���DC`y����2���anI)�'lK��bmvD�����p��ǢN����E�ٍ�jQ#�mI^���`�p�ܖ;�u`f������EGN$�,�� _;����k�9ܚX�f֨�	)JD�v��������ri`�p�E!ؚ����X]�v;�K �k���;��AM�M6Ԏ��ri`�p�ܖs]�������ӭ��]v�mT�\���;e�GT��R���3��[;�t���ܦ�[�� �eXy΀������b|�;3SWWZ��nI9����c��!D(��{�ݵŀ{zk�DBl�R�v�R�H�dNK�=�`s2i`�p�ܖ:Ŧ��9I�ӑ�]���H{�4̙��{�@^�׬q��#�R�� /��`qwu��M,�*ף�����2}��z��a���b0��݄T웝��jչ���cSJR�8݀s������9ܚX3\���v&�� ��w]�����9���,���%&\̹��=�\X���i	%�����`l��HB� `$	��MXl$ L4;!��l�_�( �~^c�ҡ
�4�"�n��D�yJ��i!��RbBY���a��BRV������c2X��|���Z��C�Kr���61���H$#\�8M[	���@���P�ɉ,�!�$g ��BH�a$� `kA0��]ظ�=3���	"A MJk B�D4�0Ĥn��h$B>��#���<5���f�Oo ��	P�=;�� X6�����@ J�
ƌ
�b[||`$�j5�	c	XĖI�j8B�vx�u���2ѣ-c�3GV��l��
6Ґ%�t@�.��[X��xg�=P���6��B� ԁI#mᐙ������H�a5�e��r7\��M���N'�!��I��)B�T�cz���Me�ӣ��h��5;�
��X�"�l�M�Mw��C�ԥ���"��HD�+���JJ�ͦ�f&��1��F��rp�Hf��K�H@�k3+I���M8��9�	��w぀�"i"���1��&�[��F,��:t�9}�肝G�q 8x�_�4��A���'4�hM�Oi�
A|8
Z�W� ~L]tL����5��8u}Sy;�o[�y|�r��Վ�z���)7!a��K�� ��k�9��V��]Ϳ���Ji����n;�������w6X3\�u�,R*rF� �6�Ef��&N7 �펎#���wf��͍㧍�N}�se�l<� �ޫ ����B�y�6q�u�1�(q�4�v��� �k�Z�c�8����Wԑ�׬��D
F���� ���`qw<��͖���$%Jr'�8�����[�Ny�u�>�X_0/tԑ541p� H��ʰ�0�	�i&ک�a�J� ����G�<�v��_;)JnR7�޼�w6X[�k��`z���D�KͲ�O�i��L�٣H��i���B�k�3+�unu4b�9���dQ4�. w7����P\�?UU}��|��j��G��I���1�:�DDCg�oM��=�f��$w5���4�QJM5`uf����v�ޫs�=�Z7P�⪝7��{��fM����:�T�3��f��1�(q�SN+ �f�����vl��v(�% �/�jft�R��.�^E��zr�rIRC��> ��vW�t�QX�җ�����GF�,y�N�V.���o*ț5��G1[���X��	bOm=�6�g5����:Mm���E�Ž[7$�HF魸�q�Ԏ�ήp.���W]Z7�7U�+���h-����9��6��r�ݻkn᧜t��ɫl�Onw ����N�7�*�ˆ�>G�=A�G�''�k��6[5��m�&��r���<��
=���p��ՖJ3#D���0����;�y�V�͖t)�m%#cR��Ƭ,�2w��foU�����Q	6f�ɔ�"�"7�����;��g�K��]�v{u$1;�#��$qXn�X��o7f�̝�`y���[
�h�����P]�vz�U�w3e��4��9�(����+�/\�ų�.�(�rn����B��)�[7Uu��)4Ձś���^j��l�:�T5KF��MQNi���36��(�(Z	 �� R`E�e�UX���>@>C����<W�`s�]o7f��������(q�Sn�͖u� ���`fd���ijF���,]΀���`n�q`��`f��#��9#�XY��̚Xs6X�T�U�f��iҡ�(4�r|��<�9;Mũ8���svl��n�d�P�W��Z��7' ����;���պ��2X���1��$��R9V�͖�� /����ͺ�8�7O~�h�UX���۳fBR���DB�"OUS�i�	��lܒs����sq��I��Q�M5`��`ff�X�5��T���r��B&E34��*R����}א�\�Ӿ�����=�1�����Ye���]	�.Vx�`�4O���Gg�N��jz�Ŭ)X�[��[� fw%���K��j(��
8�v�� 3;���ɥ��s]�ރ3i$ƪS��M� �͖fM,{�,[�|����j#蜖fM,wvX�T���I�!��ڒ_3%i$�]�]Mkw�cwR)"m�!`�������wvX�<X����͞O��iģ� �<A�ϱ���H)���eU�zp\3�����>� T��y{� ffK3'�W����K��J^R�Iȣ��j�ޞ�`fN���ޚ�D$�gb�Fm	 $�'�:�|�;�,�$n���U���󥬦ܡ��q�3vXf�:������`wCv�DF���#rK �k�s���,ޛ ��U�$� �4�%)R�"�� ��;�}�Vj�K��Yу��Z�&»q�e�N�m�W=e�=�e�����r���7n{5���YH�&��m�%N��90X�)�F��1�Nz�<]����:5�^5�!�lBt�k�ʜm���&	��s�]g#s�8cuڤ���Ǫw��Ô܌g�a�O{nn��pb�m���_�>����us���8��Tی��`�)��o	nkD�� �P�o$̷��k*�m=�.Z���>�2x�`l�7�sģ�e��P��Q�o�~��U����`��`���TTݤ�qF�`g^j�n��p����$�N�E#Cr9�swe�nk�w��Xך�:�$ٿJr�ʑ�,s]�����;��=��`{5��:N[r(�6��32i`w�5X76Xw\��T�ܭc>D��(pHlJz���<�\�QWF2]�n��D1������Ul���8c�+ �f� ���ZfM,��:^��R�4�fl�꿾��T�RBA(թh����]a�ZD���������y�X��Z���Lr6����+�y��;��`gB���CBm���Vu� �f� �� �(�>�bq��Q������;��`j�P��V:f��4\F���m#N׋Үwd�lG\�\������PaU��Z�6��������5@/�1X���L�	��*J*G$�5f�yم�����9��`s��H�N4�����&�.�ss��"2# 3J5J����)���\t}_w����<�� �VGFSI$Q:���0�y�76X�T������kF��H�n; ���Vj�w���]�v��d�yH��jJ�*9�7�I��H�F�8�V��ۑ��g�y�N����ܒ�Lr6��[� �qX��v�͖t�BM���Vu�;^oM�{������c��7�D�1w5�;�,Y��>�;��T'q$�����z�u�6Ͼt�9�¾Yjb���p@�ˤ ��'>���ܒ{<�Ϥ4k@9RG%��5@/���]�v��π��~~~}�t%���q<ntxv��ywa.�Wm �W��DlPZpe�3��&@��-5��\1����9���U}�Y� ͭP6�H$���1w����,]� ���}_$uexu��D�R��������__qX����v���8�(�q�z����y��3]����`��`fմ�5R�I6���,���l�y�=� ���@��ɿk�C_�@ I$����� ����@�?����*����s�h~�����Ȃ0���*��
�X��"(��(#b� B�!�ACl �UP�ѽ�I@t�ZDA��D?���] h0��G�hE ��:'��h�l��M��(��G�Դ���ߜ�/�p�:z���a�ԑ��U�u��D����'�������h ��>� ���������1�J�[���� �i	��O������]?��( "/��������I m�J+�k���}�H���Q���a��_�㣟��A�O�ڲk���h����w���$$���-F�
H ��  ��T0 FAcP�QQ,BE��`DX$B#E�E�Ab�DX!E��`1	E�DXEdDDYE�DXAd1DYE�QEUEEVAP�DE�DX�@E^� }�ԛ�����3�;�O������� D_��"F����?�������(A����O�N���b���O����a����a����D� "/�b�!�?����p?�G����'�O��
%M�o�����/���?�a���|��?����� ������W����?�?�3��g�����1_�EA�?� E�z���B�6���$�ڿ����h��}R"�@�?���@_�,�OC������T�#��	Bssz�(h6:`��ī��W��� �����`�� ��c�h��~����������?���?������&�?������H�����<L � ҋ�K���` "/���h��?���>��?�A���?��?�f�i���jF��?��?��?�}�� �{��t��~ ����D�����%�V��������x��C��?��?�� "/�,��'��?���?���� ����Z�K�����٧��T��ߐ�Q	�uC�S׫�����)��T�@