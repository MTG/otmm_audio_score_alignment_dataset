BZh91AY&SY����߀px����0����a�?       �I@
(�@  �����

 
kF�QE�  U*@Z1`  ���UD�$�(�R�$%*PR��� �����JQ*�**�RRU@�D���ET�Dxl�    �)ITR�I"�Po<�w�Oy�G�oU�y���T��f{F��p��`v=IN����A��(([��MP^��C����ms�
��� zx����5A�[�{�QUs�T�ЯJ�����:����^�Ъ�-�<�J�QE"%U*��J�z=�y��j���q׾��{�w�U�J)���e��u/��w<��[��UKu(��Yo������"Hйywj�r�Uc�Iv��U�n�Լ���כR�����x�R!�{o-�U�[�ŗ6���ҥ���E�ʔ��JB�����N5P��W�]���NMs��S��޷J��].U.o��S���Ͼ�{O��m*�ETӽ*^���Wͥ�Mj���_�-�7*xoz�>��ҫ6�ZW�;j�w)���r��TP��MەKvu嗽�S��o)W��ABR[�(I*R���AÒ�}�*�{�����מ�*wnR��UTܩqo3O���_w��Vl�q��9ԭ���;ۓ�|������|���+��
��ʥ���j�����y�W��ۥ^{�J���Yw��W6���{��w[�/�AEO��BURT�U(�F3R)/��;��ʽ���i�Ε\�q����U���.MR�O6�y:�Z�Ү�}���J��W�N�G����t���wT�E}��*[��Y]�u�5��y����EO�y�+6������.M.6�ۥ^          '�yRT�� �0  b0�2�% ��0 &   "~MT�J=1M���z�4�	���A�"{J�m)�@     ��S�JR�	�	���&��)5E"h�
y2'�z#M�MG��?A?��?��������v_}������UDU�5�(�� U?��(��TE\P������` (������3�@U�����j���p �� C��)�r��"���\�}*��)� U䪇$�r@�O�U���>��D~���ANJ��^J#���^HrB���!��9 �!�r�QH*�
�� �*�S�dQ� �T� NH�rE^J U�*��� � �rJ�� NH!�9(�%�rG��H#���>B��y!�G�R�!y<��$NBr �%䜞A����=@B9u�w)�Hr��!䜑��BRr9�W�rC��S� y#�NB�+��S� ���W����}/$���܅��9)�^A�^A�C��B#��{ �����rG�>�u(���<�NO$9/Pr^@� 9
����rC�<��%䜐�!�^\�����C|�y	���_��<��M�ʄ9 ���?B�B} ���H�)�����9<��!B<��<����<�� ~��!�~�r_�~���_�~�����iO!�%9+�^@rG�����rE�D�^��;��y#��#��М��y<�9<�9��C�'$H��AG%9 �)�^B��:�+�C�K�G�^HP�%yr@�@�NK�J#��G�<���C���伕䜀企���9��' B��.@ryr�/'������O!B��$9!>���%�rJ
rAW�$�*Ј�
<��"��
��ʨd(��*�P����
rAJ��NB�%�(l��ݛO���M�&�_ã���X���i��ђ�^ɥ� 4k��Y�`D��&;6�I��6ᆭk1�G[�m�ƒ	�b��Ӂ��htc�	��8�k���6lqٷ�^u~v���	b��ic)���8o�ׇ}�F�z蝼�!{�d3;�_��J�oמ�������*��;��$0����4��a��]�:#5��K�F�h�a��*_=���۞K������]��'A��Ք��k���Hҧ4i�Ѹ���$�~��S�F:Mu}�>�Ϻ �0��uA�Ra�j1��j�	C0D��X8=^!��j��i%D�.�!�!�t@#���P�z�w%��MDf�O�j<E�f9����\�)��#�J�x,�Jyر%���v�@��	K�ђ
����0[����!E��u&͠i����j�t�LAl�	±56Śt�^ט��ж� ��sJB���!�"�N�=��Og���.�\��Nn m���N��H�@ﭬ����o;�~��G&�#
�	��1�������rg�r
��<��,"x`��4l�5	��%	@�u�v�REՠ@d)�O�U�̀X���6P�H�:R��z�= fP$���-�PQ
Llm֎�N��->��l�Y�a����FF	G�S_2���u��y�x��� 4� ��`�}F=�TH;̵�_��H�MS�D{�j���&�O�g���;�����4h+[��>��
%\AA�^� �VA,Hp��=�<$r˛z>4�~����Xn�(�R��@��'/��d��{<4h���#��4�aA0����5a�;z�:37Ѩ��4j&(���jgqLs|)��,��ҝ�������c���0hg�`�E"��QG)MUt�ڄ*�K�oz���ŬTVe�.�)?_�����`�Qc
��8܆�4aH����C�A��:^-�+���D峞!����@z�K��n_����n�WZ�r{�� �@m2��|IS&ޅz�h�9�PLJ!�
s	�y�en�y�r��5�@��`�>�D�-T�,�y�ڧb3^Z��DM��,��KW)�7wc���/��X����kw�<�#f�f��j�v]�X����ֹ�=,{Z�n��)����F�(]��oI��׮ǀk;��k�����C|�:�L4���x!Tp����@Y<_�ܲR�(���4p��e4l�!Y���(zzM��ǓQ�f�T�DD���Qs-dyv��,'�}KH�%�7��<�lV��,���̆.Og��HB��fs h���Ϲr�y�}��V	�2;���y!j��m%r4�� �k;��CM�4�(����E� >�r�0��Hѩ3�Qw�K<(+W��֡рM=�CQ+�,X�`.�M
O-1�Wy�Y� &cS,aNYC�+

,�Ƭ�'Ǒ��l]��AѭS�F,�����NL�D���k�����+"9+�l��^�q4��z�֍��h�8h?a[{��x2�p���h������8�E��-zH4�pB
Gn�+�w�5�y|��ݝ��8��Y��n^\��	~�aT�S���	��Kٯd%���&�LK�D4�����g�2�iAn�.�K3I@��n�&�Ҁ�L�,�6�.�=��@"sp�0P��n~jǦ-F$��iz0M2��"�$��@oc(��H]�]�g�YNJ�o��~*����n��?x��C a��Ѝ�+H�n�������TNV2,�zL���G?��ezV*ٻ���/HY M�;�΋�|GV��5��0�fT��]
�!���f�N�5z]�c� �A�B4�2%���~SH]�<���ǔTA������{@�� �G�
�=&����4��Ӧ�A��b{.:��H��ē�|�_��Z�>ʢ<���_�����P���z����YY���`�f�Y�=ڸ�
ŇOWƳ��Ʃ	�SK�z`(��|N���ԉs
dѣv��MrWv�>��P&Tq�-��:!g��_���x��3G�6A�-${ʡf�8�5뀥�yE!�F��Cl"�T���x	�đ6�C���[3�^����\:�h�Fw8�w��ef�i����b�k�r��Gf�[�ބݡ��\��J��U�<oP��l�z�x��ݍ��m(�`'F�ɉ�*3H7/��1�n�\�������0o�ӹP���s����5�D�H�	̂rə
Ԛ�3�CP]���G�Ab��1��4mV���`�.Գ�r��dq����׍R!�'�o��f�,3d[���0��bC��MaD˱�`���xq� +Ч�,x/g�A�4��Z�풥�!DG(��6�.�tT�(n
1�lDG���<X�*-���e���A�+A-�}l��J,`�y~�}EQ�F:�wxB(�K-�1<��%�� ��E@9Z�C���B#6�s�4阮���=^#�Wy�Bu⎴���;�<�N��D��'�a1^i�c��6���3ƍ @���E@n���x;�9qV�&A	ow�Nz���P�IXQ*1�t�^���Jv2��	4%$8�1�nP��t�S����<�(��K����ېzn>�>�5A�F�4,�UE�U��<�F�\��g7�#Å��Ս@5d���*��TrOJ��fH�$ш h@B��� � �j���g��
߉��\.ǐ5f�*��cJ ��YU��]�B�$9 A��A�B�DI-��F�Af�4P�!���+�.���_^#3<�$�>��C(�U4�/m@	��v����s|�n�|Nر=�X��m�t���1 |Q�M8�%�<�h�@&�
��TI��Za
�F�L�;�#��L���1�4$��vuH�L�[.��B�'��W����б�������'�����@0�#�����O����[��
i����wO{���7�昞����4�I8#��@P3�&��@�ԛ�R5wt����潇�Bzރ����A� �<
��",�.i��2���$����y���s�}�:ɜI����23�YP ,�!�#$����t �K�#\4���hlK�)%4Q�5=��3<,�ǌF�ж���!�~I���C�@L�//�@�Ke�4��JՓ۾&�E������p�����Z�cMy�}��(�վ�Ox� 91j���K!x�yx��Ļ��ʴ!G��	=�0Ԛ���*AF1(�P.Y���\�R8"pѤ��,�}EN�$��0�QD�]�,�������N�J�oQ���%��7�3Fy,�+u,	��(	H0�aPd �ʄR*ᕦ1 4�<���K�{8.�k���6��R�J~� �t�v�=�	-� 3T�sE�ԅ�l��H����!Lc���'�|)�0Gt�Ȑs��v�ôxՋ8��r�Wo��{|n�
��F��d%	A�n�;ߟ鞾y=�=�T��`��[�_(l�}=j{�,���ԝu��Đ&�^�����k�3Y�����B��(��� =k�*%x�!qQle"j��SB�iuFB �D��Q�����پ�������y����g�aCM̐p!ת����v,���S(��ـ�s�	2�-X� �Jb�����"��ϼ/mέ��#_gBut=	���ύ��6��Prr����m�M 0Y
�v'f���4DP�,��+�fAgh��Ȉ��z�GF�	�v� ���z�x' B{�È�q���
�bO{��G�ݚ��hL;�;���E�C�B��k1��40����D�1a%�w��,����c�+��EV�-�zHV�!�5�K9�q��z�Q�T���PnH
�ȃ�i@�I���P��0E]�uE��.���k0et	��;n���4�9���\�xZ�M;@�r�QV_H}�[ �6�v'ا�)��$�Vi��0r6S!�htg�C���C�S�����0�j��-�w"�,�����x<�(1kk�]̈�v���Nb�!r\�A�p4/�$ �i��i�9am=ҥD��bX��}(�K�0{`>339y"X�/*��!j1+�X!�(3}���y�dgS����2p�Ni#4ƴ�v�4���>�M���S�ELX����^4#l]�%�N�.׉�	(C�z^���6E�L87��M2i�0�tl{}�#g�kx�����<%����^!9X˘7wVx�G��1�&l������r��݃��e9v���j�x4�.6h�aW�{���Л��:��1��eu��,�{zq�X*�P�7p�l� )�|�k�Bh�������}D0|}�lOJ ��1�>t������CD �A�^P	9D!,� YJ	���E�@A(� �)lw�І� 7��$B@M�� �tS�|��	*�C�F}aN�2X�Z]B-��3j��x�m>D��4nz�KUf�+�o��nxo=gxgj�QMz�ߏXm��rbjM8n�K�L�U��l�*�u���3�U�_Z�6m81V���^e��20��v�v�fVj)���{<�L=l"n3�C88P��~*!�E�U�����t|i`��s Ӡ���&}�7h���jà�4")�����X��l�{�#�����5tÐkd���"��H��1�؇�0�W��G�<�a	 e�摦��aA������@�vl�,�%EV $����e�� %Y@�ZSg�`ѼYU<d�f�T5J�b���� |6ǲ��A0.fh���9n��GĦC&��FI��`9��$�����=jy P��z����rH!xM�kݻW{yA5��Ve�$�:h9d�@��{�
<]���枈ѠԸ��A�7�Xf�4i�Ga�6u���]�cSZ�]�k}ZƩ�z0 �C�4lu8�ٹ���`�}v�'7��գl��3'L�HYF�g3A��f��sNi˿�i ĤA�!	k�hM54��P�sID�5*�u^�+�W�ٯQ�H)����Qҋ8��kt=� ��H�j�ɀ�.���1Xf�;���"�
a�!;НI��Q�����^���c0�A{n��v�GrI�d�dw:{߆���F4h݆�Ν��K/!ȞeA��C�%��.�S���١�&f����
�4��yl��O�E&R5#L�)���U�1�7'h�~=�Ra��1�y�8���Q�g���`5�A�Cx@�+D�,��4J�c�w�అ�+)�ui�;3��4�2e6�wn%�<_�y��4ߥ40A�ݚ��-	~����@�ˤ �7�4'����V���D�hz���9n֥�3כ|7|�ܓf �w�`qVT"ĝ����.ם��{�=^.�ˀ�
��������Aq�Yv�pH�D�AK�h:�M��x2Ĭ\�Z���X��a��ץ�,;� E��p��ᙉzxz�a����V��fmQ�0�׃m����]��{�}�Q�a�Q��(�=���`���qS�栲�M��38$�7�3r�Oh��s!�Z��)�`'�{{�h.K 1
�eD 1�k)a��V�?�$ p�|���Pxy?yx
s9c$�!<�RhB��=e��ՙ=�(:6�ˠ�j�tA� �9���^��
j*F>�ڱqh-�hN�'.�#�ŔH,z�G|��+��e�<��;��3ד�66 �9v<�X��wV�Ǔ�x�qԞx%�c���9�rq�`9��
K���Rt���m�l�'�������l��'�\H�e�`����C��ۮ��%p�W���듨�	��`�Q��2?��?/[��d��ۿ?����檶���������������^j����.����������UZ*��������������UkkT�P*�UuUUUUZ*��j�*�U�UT]U6��*�WQV����������������V������UUUV/E=��������5)[�3�ͭQ�F�ij���E d�uҹ6͆���fjQ����c]WC�n�nG����� ��[--� ��΋�Wn��X���L�36r8�KYtn��W�:���ѱ�!�<=���qli����v�Us�hw��*xb^k]nĚ�:�q*�x77�������tۢ�*��#���n0�[��c�T��3永��!�!6��n�`M��#�E8펜�� ��`���u���)^jۥZ�T㊮nڪ�Z�S���\���GUUvҭUURZ�y�:X���t��iݴd
�Ut�<iˠj���Mj�	+����
����k?�_��qN[HK O=/��T[������`~B���P-7b��ڦ��D�9��ydH:���ar�+�.�/����h�^�4�m����nR�)0I�]rm��Rvg�g��UF���]ny��CUuTY��,16���9c��K�����sA�V�m�(p�M�vʵR��:ܼP�xv��z|l�Q}5���Ð2f�j�S�g�8Zk���9U��h{v�l���n�Uh�᪓;���T��h7"�R{*�KZ�|��5mK\nYg`�U�$��ciB��DQ�n���m��
�q�8��c!װ�"m���U�j���y��Y띍ڻH �P5;d�T�S��9煗�L&�4���Z���[E�`����e9�rq�!��sc�1�Z�UP�G�i&25r��ع6�2Š�xgUFO�ˇv�rv3�BHsi����ݽ�ɸ�.������<�T��uOMV���@t���ReG��ʸ�{v4�)�L�{sN�.�l�[*�w�����\m�i0W��٦cgv�A��5\���Xf� |�[���7g�X�=d�f��M�닱�� ��F39n9wHvc���5�9�um�"�Jt;�q͜�J�U*�ĕ��5#��(���cm�e�M�*�=0��l����S4����s}�ۈ����˒KtB��)��H�V�X���T�ʽp捣qƺ8Z���mD�'GcZ�s�ZwHU�W/8��ꌊ����ԅ��E<�j�z�mC�Qj�p�c=6���9���E�cЛ��Y��-�`d��݃�f�ds�x�R9\����9kk����eur�u��ƺ�pOm�w�:�m�3�qƻv�Y��*ѯZ�ZxϤ����g]u�������[��.LH=P�-��óW\nxv�w=��m 8�W���V�*p\������صHRIDk\�����Y�V��8�Z�*���8�Xl�f��t�t<Y�f�Nd'�̓)3@���q(�\��<Vں瞸k�=ĳ̠5��R�6�V^y(��0Zn)!�Tu��<��j�<*��l\��6��k���h��Ze���͓[�T->Z��N8�1�n�km�U�d꓁����<��'�'n<ఱ2���5 Q�kk�8웴�}l��SR�8�4��<v,d6x�SGqe������w<nڜ�[��A���r*�;6I���<��/���>�:�u��'o�b�Q�X*���"�;�n[8�"k��;F n9J*=�/L����I�4��C��w7(kc��n;X�Âe�4<+�qk�R'�ie媕�]��������Q�M�!���jÝ9�1�姱�M�	=�@v�x����"6�eu��Vb+2O.�8�F9v4��}�^�ύ���yBZ`f�b��$�Wf�I�0����l:��� 0��n�'5UK���ĵ�Ş�a�UU[nc��2y	
%]�3iSm����*dz����*䰑T��y1�,�z���3-J�j���&�,�J����:���f�����sƺ���8����i�� ��]��9��P��/�;�+غ��Ǟ�uP�U���t�uV8�F-�,Z�r�m��D�*��뤫��%^y7c�٠*�����u�ԐE������*�Π�骨�+UC��.��kR�N֫e�娭�81�s��bݶT�O��Z�U@�D6zyh6*���A����^v���Ik��]�2�ʙ���j� �9����$n0�7n�;	�dOm⣞����䓓��f���:����T��O��<��y�Ɍ�k�������Yj�OCUts��N.'n�T�T��}��c��U�� -��
��)iV�*��NvG�I��wNLb�zデvU�X�`�W�!8�.�:��ꪪ��{�J��[[<  UT�e��Vݷ����/��2�������u�6��Z�����]uUUYv��ّ�u�nX������;k`)V��UT���UڪꕪT*�(�6����OUUUU*�UT�[=mPU/V�TTAh�����Q��<=���k�]�$�:AڵWnez!GMUJ�5UUUiM]� ���rn-W)U[E��ZU�[M]��Ac���Q?n6L�۬��W�<*�E7B�]uUP媐6�s�JU1��T�^ۚV���l,�:��tWUnќ�%�]����
�-�)�UG����V�ڨ�)l@p�z��E[Ur�
��Ut�����M�;��	�c�WeZ��U-9y;I�2h@6U;bT=�ڮ���ڐ�\G:7oYPz")d��mə0��7j��v���Lj��^ݷ�i[g���ꮛ�,*��@ ������
@٪�T�<�Mu�����hv;s@��֊��*�
����	��.�:�f�����;�+kmW\ 5u�R���CX��ĢV��8f�4��ꪶ^��H�UGg;�Y��d]U!0�z0<t[7�UU�T�zv�QS�\�+m/-���� ����*���d��{PWBQ���9uum�r=T���U�>��p �&��X��8\�m=�>Д<UUF\���' \]�*�Pt)ų�lL�UQr��-&^��S��[��v�������)�W ����x���-ˈ�C��G]A�SN�y�ij��g��\�F��l]�V���c��꧐�E�������q�ҷ���ۏ[m�U�q��{�p�9Wțm:-\Cb:PF�N֊�܏rn�]�Oϫr󶤪�A�֜/����2X��{-�fx�lQ�O�}�}�ˎa٨�Vk��'��k"#WK.���vkS���C����֎2��Q[��P���ik��8(39��|�`��k�kV\�7[�De
�D��5��ˢ��^N�
56�T��dr��J�WHN��-Ͱ�@�\��ƍu�<�t(��#�N�q�����R��Wa�mWkp4x�Q�[k�7S�1nK�Rr�U���%[��`�:���N���kP�P ���(Ӱ�y��d�;m^(���[��*&�����[�U�=������tR� m8Wi˱W<9]���s)����j=���i��$H\�vƔ1������]�۫8TPW�5�WgR���\�G�'��9�U'n�ە�$��z3\�;���	O,{�*�*6�������|*��F�r��H��A�r����D���n�N�mYH��bۂ��[c���i�s1�
��\6�t��.2��v<Rl�8�����=���#�
uN�ݶ[������;�s	Mgn�E��i��V8�j��,t�Pu˃/v��#�۠�M��VX�Z��雐�M���v�٫��0N�9K���$E�+�x�D�+��8=��s�T b�)Y�V��ˎL�����W��g���S�UUX�����;�6W����ԫUJ�P��4Ke�t��7j���Z��,�N�uUU�V�����ynI�bWSL��hZ�d+��s:敺���ҧf�����}W�$2����SUQ���jBj�ڍMmJ����,,\֗�\e����m�4X��`�������n;���UUR�ԫ�[UT*[S�C٭'2�r=mPUӱ�ꗝǱ+ҭt�UV�UV��{-���j�3WJ���vي�f��� ؇T�v"Wt-T�08m�@����m�������w.�솺#geu�(r��N�*��������D�L��AU@��Z22�ZU��� �U*բ��rQ
%�PRU��Qі�sUT�*ՌU� �a ��3�&m���ЭU]A�J�.�BV�+8�:�@En���U[JcAUK��?����]mʳj���WKUU<�uj��*FbU��g��f��l��'i\=t�UJ���ERa4�W��]6��9j.�1F�-<VsrWa��.ك�Ln0nDv��聬zɝc*7jdݙ�J���m�ڧ�T�Oe�\��-����z�m�J�	�5����qq���4����Ƀ�$c����y�v��oG���؍��ll�!T�`��#n�ܻ�ZtW8�jUZ���xk�Aƺj]�u�H�p��ݹ��^��WX�#������	VU����G7qt����:�U�t�Öy� ��ȵ<g0��]F��+O*p hӃnni�Kn�-�؟T�p R3,k��UU/-��&��EUvW�ȁ*�KsUmUA��m۵UPUU��-�NVS�@�
�UR�UPUUUUZ�/.�mpfܫ�����
�q�8%��[�w�}M����
�hZ��U��8�M��W
2펂P��:�g�v9�h�헑�-ؔ�9P�N�IY���f��PpXx�A�`��ۋ\3�,����d�����6)��j^0���ڭo��AE�<@PU^��m@G�8���?��/�k��g랥MO�EEe�H͙�%�"T�a�"b2�$������}�����~������%mc&5,�1�e�O2�ƥ�v5,��Բ�cRʽ�DK���+�Բ�5,��K*�Rʸ԰� c#�w8�au.5'{�R�Rw������Ըԝ�n�Ƥ�su6Q��A�#e�������~*�� �_�p@�C���r!�&	@Q0�(�
s��T��QLT%CJ�	ڢ�:{U�E�PqD�D4'�
�P{Tv�l �v ҁ�T�$RHFN�TXQ�A\:N�=]'���$+D�
mSH��� S0���UN��S`�(��mL�_GH��C�J�x(z�z�?" {H�>@4/��N���	iH��� �ڨit�v���W	:z<DECb��N��E�FQ4����(����z��ڨ���=��	ҏ̡��.*���J��}=��E<�O�>T0T��? ����&� �_EQ�_T��q��	%�!)�U�1h�
(�A< D>���x�x �"��>+��U��SԱPQQQE��AB�LIMRDA	��AD�D�i �@M ����\A G�^�O�;�l��D�2Iad��a`Ēe8`� �f!�@X1,DX8�L�DdFEQ �z |��eX��W�~_���;��+,�rb���
�+%�bD��S)�2V�`�� �Pp�JBH�!p"(�à���]��|*��P�Epѡ@�ȝ��A�C�T���R*�����������՗�#�9UETUUO���_��y�=��?�]@ U��E�E)M��Q4��r\�D9�	���Na�NH)�j�#�2�,���3{��n_(lx<���8{=�]Ƕ޻�����55�}�*�Bg\�UU4�-v�WT��g^�L�ۉQ�T�$�8x8��������cz�s��n��)=��y�dvND�J��n�`	bۚ YYy]��;<+=��N�֑u�2�G)��<]�g�쀝v���۶�8,e��<1Ǯ��舝U;���C��<ظ;��x�h�^Ě�y:�r��p�dhE��p�1l�S��U�RL$�ַ.8�p�)8�[�$�9��/<$v΋u�EbS�ܞՆ9����^h/���U��c���CQ���=����y�ż��dD����I�4�pr��Nפ��8;l[�9q��>Ty�U�9�����6$%H�r�1r�y[F��p6F}f�+��Y#�g݃���9�'�©����u���˭��9T�y�7R��I�;u�g��2�B��
{1�)���&��S4n�%�m� d�=vC�̠:���,�^ۈ�m� �n FM�U����^8��e�ru-�K+ڈ�\g�#���l$<�v�&vnΌ�lf$��esf�"�g1����J������n�]��"ųrk;�X�b��3Ү^pXl��q��^�AUaި�gY�6Mn�wU�
#�1۝y�[ݺ������ʇl�#��t�ˮ�ܱ�[H۬:�J�F݈�`���v�"$����W384�t=�1���EU�I�Z��OnM�� ���Pmu)���g��Cb�R�:z�ŜZ�r�<�v��� ��q�vP;/�ûpl�{=rU^�Zl��l���mZ1�-E;���5Y;*n�v ���5v�/Z�KL�ݹ҂�����-�*^!�E'2�ی�[*�6�r���7:��������9gi�Be���ϑ6Ne�gK��m��x��ُg`�p�dQ�qvyGf���z}V 3��v0�&ێ]�+s���&�l�r�[��M3q�ѵ�L�7[92�m��=h�Tf�[�;1��@�����%ֻlEѓ�D|w�:G�UM�:A0@M����������SB� �_q6�lЎ*��n{ַ��k5��;\9,'l�ܽZ��ϲq�����8϶��dZ=��� �E�����5΅���L`:h���QM���m8編�;��ӈŬ���qK<uv[b�s���In;rak�m���v)��\ԵD�ꛆ��7�Pۖ�����mvK0a$K#۵����/������y1�iwQx��DpLv��ww���#u]gDf��,0̴�5�qݻ9퇓vW���A)����l�p�A�pv�Oz{�����:�~��i%�y�6��U��r4�.I�yos�O/o;$���m#�{��9��3i��i&��O/o;#��X�-�]��c|9�ȗ"@�m�����[ʻ���o:�и�C�E�%���Uݽ�8�y0;����^Jw����襂�[+i�����U��:KӅ7;]p�^��C�zV��=�z�����y�qu%��>Sdu�"x��-�
!��>�s(<h�mP�tj2��F��E����fBY���E��� ��{��=��]��u��,�P$XQ%(�%w���v|�84��?'|����j�f�j�r�yo*�oweoJ�ou��7��E NH�.Gw���;zW{{�o�r����/)Pn� Ui�X����[[cp�ni���$Nz{>�y��mkvjr�t<�tFy2�V��J�ou���^#�����-B������{{�o�r���ׄ{�O�
�3��G�,'��ܒ�j��]��D��(R)��d���\�v������B�$H�����lx��u����ܫ8�Z'�J$�e�nX���H�����Wow]{�sq��q�Pa�p3�/M�K�㙳��:�S��z��o���ow�Ւ��i"i�]��cuw*���˻�{7��I����
�v���<�KKB��3k�fM{�{�n���n
jF�rH����Ǐo�Ť���f׺����<�#*�7E9cǷ�w����w!t M��A��`��"�)�;����=����&����:�ou���U���cǻ�F�����$��T�%��n�k�GzP�i3��J�ٳ�ƮzSO�NHq��Q�Ip JI,g�r���X����P����x��p"P"M�����cǷ�w����w*�sG�ED���nX��s�����@oou��������(a���U
�=�t��U���Ǐ��{��q$��&D�K�ʽ��x|Ws���SIa���	HZ�U�U�2W;���7�qa@�@�Lk���6�g�f+/l槮��	۳fn�6��9])�ݺ�3�ڳ�{
g+p/T]N�9�\U���i8�f�\p5��d�O=�v�\�l�F#h�����zP�gp�g�c� �]�4t��c�뚫q�
n刴q�(�-�ict0�I����9K��z������ ������^�w{�A�c�#����cd�e���A]��/�/�||���M��YQӛ���3(\�*���x������uVw��96X�FS$�w?�
 ���yw*���ctsC��c06�jG[۱ź�A�ޱ���W�uh�r����yw*��u�y�[ۢ��"���!L��qW���{��u��b�U�@m
ǫ��q��Iw[dR��;fu"-�A�p=Ub[E�p���;���7*t�� ��;�������}@ G{ﾰ=�&�X�F!�8�{vxV���Y�k+M�ʗVkXL@T�n�{�C޺G�!\p� ,�&"�F�ښ�3�6F�m,ff�['�S$�{��'��(:���x��9Ώ/w:���MZF�K��U���>�u��ea��&��8�M�$�}B�{ﾱ�~����su�w��8"�P(�l������[۰a��^��ù�胴�J�O�&х�(��
�
u+�S�]�_mԖ�n\�ۣ��D��{v9��۽���;���(�Q���s�n�K�{�����F누�FHT"6�n�]{��JD@�&� �P���Wl}�u�>�"���`d�����ov�g7]{twX�=�I�,X�F!NI+��U��u���>[��O�y��D�-�taU�Oc�\d�'�
�r�ۢ̎�e�����gw��ν��c��η�\p��A��6�q�[��Tf��w��,����284Ӂ&d��o:���n���t����6d ��8�Q�]��Y�}�瞟}ӵ")��|TBPs��^��G�(��iGc��|(Un�gN�'��j�the�UYd,Kpj}\xz�FɁ�����[����Yƺ��;k܀��Yl�d:��{��c��νݰY��^|���"bl@b�,x�y��l�uW����W"��$$hB��W��ź���u�oJ�wĒLd[L%���U�ou�o:�v�x����Z��E��{{��yo*����;� (�%�r�S���Y��fgn�7���[O��\��2X�`��cuú���F�����r��6��ɞ4�Wf����r�����M��_}�RȚr�q�7Fڛ�4���cr�>��-�¼������':m�k���� �Vp6���g�r���ҠF��qD �� �ZE�	�g�q�^� ��3��n E+���T��SO<�L�S<8/`��n2�� ��J��%[�Bd7;�Mv�Y�*^�Nj!@t�>CҼ�ϋ���56��GL�X�&�L0۞��U���n�����4��4I��q1��ݰ^-�^��X���Ѻ�4P,8n�v3˹W���=弫�����M��n��*���Ǐ��{{S��n�чV�OblA%�bx/o:��^/j���X����zwQ4KU��T���H�ػg�������`�x��A	��}Y�"Vz1�nw����O7�K��G9�F�O'\��)��V�Z��}������B�Ҧ�E0�wX���[��^!�b!��FH�EȤu���0����l�ګ;��|FD�M�ۖ0�y֎��{Uv�>��<G7 $�`.6q����{U{w��o0>��8
OrTWѴ�2JP0`a�r7+βZ��x��W��lrv��ݍ��<���%�A��!�Q����W�{�a����/H�qi�$h�㊽��UZ������Ax����4q�9#� �$BNX���:�킇�?a��I �I$�I�_zn�۸��*�j��~5�AA��2�$9�K����S;�& P-�* 
�3��|�,��vi ��s
�8k*�A��Y�d^5�߁^|�-A�U�����ntޚ�Al0��3I��BS~�EA�����R�9an��lg'�O�� ,8Ez��Aj��xg;i�`&C����GD-hx���X^���u���fFf��������� bT������@ Ҥڠ4 P� g�����]��&٤'��n��i�~Z%0M �{��MY�@:�p��`mx�l8.��'���v&��2k� ��F:�2��=��=�}��!F�:2W�����r�n`5��<�r�J�b��=@�h61$g�^��4�DI`i�@߽nҒ��1h�WY�f��8c�$K�&5�{d�5TU	N�l� ����P�˔
c��N��[����)��{;��d.�;v'H�蠞Hʂ&�j(oULBH�0�2�v<P8
�8�C �?��S�@��rS����:R���Ϲ�b��@�=�/�H��.H��#��M%����)N�׿gJR����9��)A�*�����'��9�կ��ekF�Z�=6u�ǹJS�u�3�)JO}���Cܥ)�{}��JR��{��Y���x��84�-�ّ(T+�d�&���䪻v���n�e���mT�zvD�h��1��.I�j�47��V�MP����Ҕ����O��R���}���i�~�5	�N֜rI.ָkJ���}��JR����R��~k���JR�����{��rS�_��k]1IQ���5@�_}��U��MP�=��H�����9��)Jy���t�)�#�E2����rAXj�5C���t�)I�Ns�p4�����JP�������f;�Fa���I�FD��8��(�"y�?���cԥ'R����]�o2ַ���y��JR���s�t=��`����}��Uo}��Uy�B��G�\"�Am<�ć*rwl����ͫ�A3�'Z_\f�ű(j��F�+q�: ��k�ZA�/����JR�>}϶R��~{��JR�������i���<�1�N[��޺R����}�����~�)JO}���{��<�y�t�)C�y�\-�ZѼխ=]�cܥ)�s���rR�߷�t=�Ҟ{�s��(~�>��4	���"[d�"H�ܺ�HM��s��R��|�|�t�)C�9�ǩA5C�޻��ho�p	/�3i��Z�Cܥ)ﶹ��JR�� 翟�����߹�JR�����s��R��G���2d���Y&!"tG�����y��}/-x;�d�B{\���
�s�6\h,�c���t� ]�v��'d=s������:�훶f�%ƀҒ޻ў���6p���hD������%��<�{6�.�9���7m�`��X��W�cS��݋��	n��WB�G=^x3͹|�K���k������lt�"M\@���q����8:��b��h�P����!-ik䵢+Ìn
����&y�]:�֗nNz�����8��q�Ľf��/[�����]�o8�)C�￻�)O<׿gJR�����:�(=�9�)JRwße����5�rAXj�5Cu��ꁵT���s�r���k�Γ�rR��>�٪��;��(7��Q�n�#TR{���Cܥ)���Ҕ��r�cԥ)ߞ��)JO�p��j���7�o�����}��R�߹�ǩJS�5��Ҕ�'���t=�P1�.|J��hI��MP$V��\��"�����t�)I�ߟ��/r��/Ͼɽi��K�:�d�
�dD˹�Or�#�J:���آq�7^:̘z�S*��˅�0��1��Y�pV�MP���t�)I�>�:�)O3߹���e�J~��ǩJS�ts\�V�����3-o{�t�I����C��D�T�E6�R����])@���y��R���w�ҟ��b��~�p,ֿ�y����[�{��=Ϲ����(|��=JR�����R����s�r���G.��jލ���3z޺R���}��R���{�])�����Cܥ)�{��ti�1{�I-5eSwvծ�<�_s:R�������)Jy���t�)C�9�ǩ7J~*����p�z7f�X�f�s�z8���J����R�.{f�=��b7��0v��'�<S�������Ry�~~t=�R�g�s])JP��}��R���{�t�)I���ٜ�a�6nu��Cܥ)�u�7���(~�>��)Jw��:����·�JR<�2&��v�5,��-��kٞ�[5����{�t�?�� u�fcG�Fj���4��4M�X8E&�sDAZ�a3�bqP;�5��y��)Js�}��)@�?{�-p�e�j޵kOW[�cܥ'P����t�)I��s�r�����gJR�<�>��&����9�D��rD�.G�h
F����]r���k�gJR��s��kԥ)����JR��~E~�5g��%�����ln��Pغ2$`S�]��n]轫����s��aoL*�9�R��>���JR�<�lz��<�^��C��&}�9��#J{�s�ֳv�37���z�JR�����)O<׿gJP4�}�9��)Jy���JR43�܏�4� ���*��j���gJR��}�9��)Jy���JR�}��*��j����h��J0�"8��R��~�:�)O3�s])JP��cԥ�>��	2���U�{]��<Δ�?��'����
��f�-��y��Cܥ)�}�����(y�}��R���{�t�)I��s�v��Z_�Ik&}򤌖�ME*@�xU6�L�`���yJ����b�u�8I�ݚ��"`; �j;,洃K�����ֶkJ���{�t�)I��~s��R��=�5�@��H�����Aٍ��˻R�P2������9)I�y��t=�R��ߟ��R���9�ǩJS�5�����a��yek{��(~�$Ͼ�:�)O0���JS�@d?�����)@���t�)I�ߟ&f��#Y�h�Z���=�P�g��R����cԥ)����J���~~~t��R�r??��a�1��F���JP�&CϷ�ǩJ�D��w�3�"R��~~~t=�R�{�s:R�����A��i� b���
BbJ�@�5Գ�77`ܖ��,��vN�\�;�hK��^�k��g	Ϟ�m�荮�� U���E渄:����a>K�����0n1̋�����y\ͧ�Ma����p�K����o���';-WFT��!�}8z�]�w8m�ʝcFڣt􃇮��7k`\M�KZ4��P�!�N�7b����;=��z;W=v���̅�;��Qm�+`�j9�{����w��:��e���;�v�MۖW�#��������"�)�prC��z��sh��}o{JR�����t)I���:�)O=�9��JP��}��R�����i�:WT��U+޴�-�}�3k\��<�\�t�)C�~�c�:�%<�^��)��)I�/������X��f���=�R������JR����R4��k߳�)JNs�9��)JG����B[#���7� ֿ�ZZHI�Y��=JR�����C��'��r���>�M�H5�]�dx�L�+!&�M�[�(}��Δ�({�s�J{�o��J���cԥ)��}F��i�
n��zٳ'��a�(�{0Jr{tK��L+Ν������-�kIɪ����'9�\�{��<�y�t�)C��}�z��|�^��)��}ϓ���bM6�i�,V�MP�߾v ���Z=0��\��!��i�N9���@���f���*�f�J�1;��R�_�y�Cܥ)�5���<�%)>�:�C�#J{�s�+N8$�
	�j�"���eJS�5��Ҕ!I�s��{���,�2oZA� ����f8�J�*��v�]ù2�߷˥)JNs��{%)K�s�Δ�J���R�����}��t����Zm-��Kٙ�k\5�@~�����Δ�-`�s���)Jw�����	h4��/�[��ա������a�y�Š[��r �DV��ʪ]v�o��Vn�$��jDm���T=��(y��lz��<���t�R��{ٛZ� ֐�`��I-d���If��9϶=@)�o�)JO���:�)O=�9�"Ҕ>��5�n���{խ=]o��r�����])JR}�ܹ��!���@�FH��,����$@� D���S�k��:R����߶=JR�����;7�o[�-o[�Ҕ��}�߼�rw)Jy�s:R���=�cԥ*y���t�ZA��g��r���H9v��Z@���Δ�(�}϶=�P>����R��>��s��R��5Ú�k3y��7;0��.�Ge��׃�}h���[;���2gg�������v�~s���`-O����>��^�)O<׿o]JR}���H=�R�����)JRw�ό�f���L�rAXj�5Cu����$Wў��t=�R�g��R�����cԍT=���E"d0 �P��T	Ns�k�r����9����!S!���3cԥ)���Ҕ'�G�k(�?7[�z�fZ�Cܥ(��9���(y�}��R���^��)B~���WދB1���3���W_�8z�w&���އ�JR=�9�o3{��Z֭���z�R��s�R��!
�����)JRs�~~t=�R�{��7� KB4��-w�m�[�Zꉥ�y��ʮ��.�γ%8v�=v����k��w��i؍6�R2�Y�pV�MP��|�JR��}�9��)Jy���Ph�����5@�+���u*@��"��EҔ�'�}�t=ʊ4���9���(~��lz��<�^��H����sן6%l6q��T=���)k�9�ǹ )N�׿gJR��}�ͭp֐kK�17�H��nAYk޴R�(�8~scԥ)���Ҕ'�}�·�J�X���~gJV��K��c>L����7wmZ� ֏}��Δ�h�!�s���R���s�:R�����cԥ)��Y����bI"�I �K�n����*���?Q_���n#:x�;<-�����ɨ� ��`��aU�<�{�3���
��e���=,�#L�w��}c�����7�B���/$���Ɖ۸�"1�o-��5=���"
��������{ @��
���DJ fW��e���7�����Qf^&�E� �Xy���Z��tah���j�("�L���L3g��4M$�G���]vF$ՈN$PfN��æ����v��Avk�w�m7��vF����ю)Cٍ�sv���@�ѫ1�tk��/];��5h��gy��Mt`c�T���K�� Ն�^�3��l=��-���:�! Zkf�v�q�.ȋ�ѷ��c����V�0  4�(�]my���@l���&�߭y��A=f���"��mQ0��(��k1�"�<as3�=I�y�זkμ2��AXH������(�h�,�2�H �0� �ߺ�I�-i �ʲ�D��� �Đ�0&Є�t�U�7�;���u6��k��B4h�)8��������{��~i�k����0��J�	֫i�]�ۻ��Q��eJ���:�*�U]UPM�U�)ZY�>��n8� ����n�<顷C"�7&�e�U�M���٩�/]�s��m��z�兂	݋�!UsFu�N��ŵE��遺�dȡ�=��OG<��\�d��9苮�>�<W��ۥ��Rs����[��۩�=f��f���4]��z��ێi����r�����u!L��%�q<2��n 뜼.�ȵ��Vz�1�N���1vWGGQ��t��0I\���<��lk<)�K�i$L�&6Gh�0vHmg�<��6�3�>{�{o��9s C�\������z�I�y���G�9����<Ls��dNXz��3i���x�y�.�g��;l�^�{�L��y`��˘��3�sk��5�Fn�l��|�\�@��u��ٲ�a��^�����-�����G&�,[�i���.0iֹ�;��x_/\0���K;��s}>΀��]<**��p"�8��=t�Y:������f�֪Ny����6M�q�p�K�zu礸��.�hy��`#�[���<����8�+���z��y:��q:s�ڸ�mp��,���l�qs@�'��YZ�{����E�J���7WWL��x��=�^d��Z�uIM@�*b��Kt���w[7�Wr��h�;¸��V�.��<u�	k��`�&�\6�aM����p%�##���i�\�Oe�&��Q^�&�ְ08
���
9ɺ8�z�����=nʞ[�A�����E^��@���)�Qmݤ�x�7+�5Vp
\�@�/`n��͔�]��[i8x��+'.�)�����;�L	<�$\�i�f���{,��(�x�f��47��&8�v�� |�N��x#�F�Nr:.ɞ��p���9���qp񣮭���l���cI�٭����%��ŜML[�C\���B�\�g���X�`���PQ�G�h#���6��k�o����޵��f޷����)�y��i��i��i��i��)��i��P:?A��� �� �IA;�@ |��
?�`ڀ����v �����@�Ϗ;	��Փ���:3�4<`�o<Y��s�!s�Z0vx�<�hJ���K���͔J��F赑;���j��U�I�
;c�[�����A�s�ÆA�8�O~��|||�mC���	����:Z��rXջ=n�vg�x�O7l��vm���\9�['l�on��g�=�u@��C.��rR�ی9:��Wd�N�:��=2P]q8�Ra�RUUP���P�<������q�`���J����hѠ�	n�0G:�%j�}��o�����EMUk���H5�_߾��ޗ ���{ i��G0�yN�%@AR⢧��*f�t����� m��Rs�M��K@/�/`۶Z�au,��=��{^S���"c��i����O���"M�VG$�%��7wxK_�=�`$��@��ӝ��G�+�{IM���5*��������3�kK_�=�`u�zl~�}6�d�)K��'l]����'1@�pC��Z�ne&�5kg��T�Wn(�PH���ӗ��-uwʰ�yO��r6""C����	���3�2�UG�l�g��ĵu��4H4k��2lZB&,qă!L210*Ę��Y|�DF�9�3Ԝ��}���7Y�r �D�q5%��Q3qW����{Ԝ����9�v|�`�5X|�%VQPT�e������DG$���7X��`~�Z�KIw����11|��]2��g�� DDD4���yI�	&�x �S����JXȂ�
�Wu]��-p����Nֻa{�z����x��>�{�w��q5ue]�\����i��;��"M�夒H֖��:���h�ϣ�Y$�v䩮a�w�{Ԝ�Ns�A)7�}M�$��Ij������Μ��b"{�uW�}�w�^{�s:�~�⡈;�}r�z,���u`�
�E$Q����ZI5��}~��3����=���%��}��������⅖� K�`G9��N֥��#��� �����;aQh��Ou�j���qt�Q�ꮖ�n���������p�z��Q9ywz�I��&�4�n�#����Z~�]��w�?M��ڇY]������9��y���j����9Ȉ��!��O/�EM^��7X �W�9�ה���� ����P�G]��Q�f��-�Zg��`.�yfuW�}�����UU�
��8"q�����u�W��f~����Ml�ڼ��ǰ>Z�M-k]oﳠzW�V $��`�5%��V<i�BN�gJӞ[�=u��]U�U7�=T.�@�V  GvnT&����N����7X �W� �r"4=�Np{���U*���H����}̛�G �9�H�� ��9���|�H�G�Fb�z%Q�+�ٰ{=v�ӾO���ԛ�{^n� ^��Q3sq3SD��]��9�G�9��{�v|�`-ih3��?w�^�M����װ�{�}��9�+�������k�{�-sZ^Iw���gҲJJ���4q/ms��2r����]4&�Dܹ���d��^�b6�-t\f�<u`4��m��e�,ph��)�y���cvKl�ӷ��:Ӻ��(�-v	�ӂD0֞IZ+��e�G���s6wEnkc�����xw���zu�<�n5k/ r�c��l
�-���ь��n�*r'��Y%�B�kW��-e�����~b�s��s�{۴�����Aoz�R���Р��a��s�����y��;#GF*W�JA�*q�iiiS����/�T�^0���`M^�ה�KZ���g8���GK]&�r� 5x{^S�(�ot�[29���o:!��Ml����o�� �&�H�s��;f 4����WW137Um�e�a��${��� �ܸl�5q�s��w��8~㚆qqeM�A�y�7���8�%��$����x{=�`{��9���x�7%����R���79�쾺]g�n}���� �A��w���7u�J������?~�N ��؎Dh�f��N�f�d��6�y-�0�����(JB��]B����w�u�~y�G��o�ꫜ��~�)���a��7����]�b���p�[0#�ͼ�=�Nr �q�RF!5eӎ�;y������큞�^N�����A����fdr�$3wSʹ�0��*d���� ]M���p���18e�$lR��h�x_5+t���R���	e�3�C� �y9����}�}6M�M�0�ˍ��� �y���l7�kZ �g����d��V�h��b��� ^MG ;�l� i��;�w�kZI =��8�2����A����GU\��o��N�_�	� 
(��Hj��V���@<T=^�˜���]��ߝ�W�E��YpG8,�@R?}:Y'�{Ӏɼݙ"9�����{ʇ5M�7�����f=�kKI{����f��Ffz�w�c�,�[(��|i+/e���Eܸ�2cdr��8.8Mx�]g�`�=V����RW�=�fs�w��[ m��s��2G{IN�)!�AEL���7���9 �m^��S���7��kI��`���cu��cJ�n� >��x{IN""��t�������䘂� �N�l���	-.�\�{�E���;�}�::���Q���ֵ��v�vL�V)���[%{%���o# j���;IN���B�����\��U�r���44f�T���]W�����8�!�Կ�{��ϡ���/b*����̉}�F kj����#����9�;�y�h#r�lj�V��j���@w��8I��#�9�Ϲ�"�.����1ڛd'&�w��L������������s�"��KHZ�v�����wٜ���������)�:�(!�AEL���y��CM^�ה�ɽ��K������[Y�I>�)]��4�D��r�������\S�ƺ��r��3���{�q�.M�s��������`�\uC]��\�	����j�:��8��H\��[�kjR�)2�9���7pU�x�v�����o��>w/XWqY��O����7:z͉���=§Eg�3���c��l{vYd�}��.tU�s��q�/�Su�窎���u�I�������J�qpq�k�j)P��J�(��!� {g��0[�&--�5��2�%U�����͆�Ǫ���Wj����K�?~�����-$������?w�<L�v�f�o{�ޤ�9y7�|�F 4���2�d�^�&�"c-�����}����[r9�m��;��K�j�b��͓TM^�Ȉ�;�o#�� �k�p>KZք����Ͼ� �?�{Р��L]��@j�G"9�yI�	&�@�ܸm�kZ���1Kj���-b/b.���n�Fc��'	P����Z�N�69�V�ܪ4㜏v��{��9�;�l�s��p�� �"�&�
�(���-�]U��s���'��+�'�`g�U��u�eGdl�U������p%�f�zkl�D�&[�`l�C@.�!�p�\ qA�US�]u�� ;ߕ��z�DG9 y
PG�H\S5���r�͙3�l�Zֵ�#KKI-3���h���p~��3Lz�;��]�Y��x{^S�%	��9�*�����I���(�E))�Ve��O�i� s�ȎDjM��;fm]���^�C�k
�il�	�㕸����+��<��\�������q�^��e�{���{�-c!iX�l�́��}��޸m fg��I-Z��\��ǰ3�k�+n*�*�j�j�@ ����� ����}�kI�IkZg��Czq�R+m6��e؃���=���U{�.6�m��I�I$�S���j�UWU@R��G?Gm� d��Дh��v�����O�3���ƌ��5��X����.$�V[zQQ � ��!&`���Pb��Qbו�2(��L�UP@LN�� ެ����O}<u�&3#0���7�,�m,뮷fjO	�M��#D�:�{:��e��PƩ�)v.Xk��X���f&�@�!� ��@ ii�'�`c���ѽcI֍�ޫ�N�����t�H{m5=bb��w�𝑀��zڦ��,�ٓ��;:ن��M�g�Ԫ� iq� ����Z`� RA;�P�,ՔD���!�4Lփ&n�3���f���");@΢3�:#@Suhу�N"`�l�P`@
V��)�U�)Tq7�#i��S�T����
x>�/���N('`ʧ�/b'�_�D�=6�h|N�;;(�P;޻���W���.��|{���7e�Ds��� ����a���{�w�ِ �W�G��UY5!WdU�]M��	&�@�r9�xv� �ڼ���=�9�/RBB�M���4w]�n[���9�lF.��!���w��w͸�p�7.����`#3=z���7��� ��W����}�����byqWu<��� j�������{�g�7M�-i ��LM�4ݩ٭�"�.4z��$���G9""9�<����}��v��c�lQ�:�M�m�a�	/��jـ�W���9����@+����Ϊ���Ȱ���9��;�������[{����������̸���j�)b��"^ݼK����`�[��\�i�"��p߄������m#%En��l����8K��s��u�f@��P为��.
���̽z��$���\6����Z���&ԐjZ)j.��p�{�u�fDs��x�]��^��E-��R������G�y���;�=��$_=ЮL�c<����ǨYM�ff]��е�kݩ�g����t��V����9�܇�����!�1:�����4�9m��������G0�Huf��<�3�g�W�Ck�$��{��1��D�[W �n-c9�
�dV��yB���p:��j,����v7V�+!��j��yCugr�q���6��=4O��7�su�Cx)������[����ql��Q�����ۛ8W�I�3���v�,]U��j7�����$�J��[e؀��=h��m<�p�43-u�d�v{(Ȍ��+��bV�r=�>���������O����`���XI��:ճ j�;��űGD�U��[f�����	- �O# j�O|�9��	�4�b��I���?g�kh3=v%�����M���fs�g���V�������Hڼ6{�XR��@�DG_�k`ug_�2�IB����o ��a0�Ȅ�y�u����W�jP�;�N#6:����m^|l���O>��L�K�xӵ�rcj��e��	����/(ot��2 j��=>� �{�`La!n�(ܫ��{6���b\I/�|���`a*F�� ��P��ʿ?7����?��Pf{&s���31��m*[V�3�M���`Dr J<����F
dJ�n�n�Uw[7�x����{/&�@^W�@//^��TU�AWˊ*�� ^M�֞F@M^�������bjD2X�)�ʬ8���6�ݲ l$8}nj��N.��5kg���u򍷶����89w�?g�k`��==��G" I7���S8����j&�� jo ���+ ]I�֜b�ֵ�:���e���r=��wپ������w��N�R$P������qU��;���Ύ�'�Y'w����j:�Id���H��� 6����9��`�%@Lc��GE[�����[ Z֖�6���ʰ�{�4��XML�����;�n�4&[xS��8{v�V�����-�jyi�����T�5
�j�fe�{�y %�����s�΁���澟���er�ɭ�v���&��֒����7���x\���E�w5E�ww8���o##��r���9�w�`{:6�r[%��������Ύ���9����{�u_��|��������di�N��7���l~n�s�����{��ԞF�y�k-)l�0�VZ� ��%�].��d���륨�f��vt~;���s7u�..k+*���Np����<���G#d���`w�<joBsU��E]�`{��ۿs���9��o쌀��^��)��D#ZKI�p̀O���U�W%� ��# N���RS�%��@#Д�&XU,�P������;�v;=粷�����I����Ϣ�sؾ������Da�w]78��D4�������{�o��x��HH%'FA�Rʸ@�$	�(�
��B���Q�E�:l�fk7�ӳ�\v5��n�^;5ٹ-4
p�vu⧇GtV��� 㥸���i�5���1��u�g�v�8ㆵN����vx�y�;����K�ܓ�u'7s�9K!����ݵW[ak�$Y���9n��d�|`��8 ��`4v\��U���x�lsv@i^�[�����Gb���x��QM�u�.�Z�i�%���nܖ�p��uQ���kZK���㩹�ېRB9�\���g\Q���`B'9ӽ��#�L&Ꭾ_Ͻ�ﾻ�lM�K)l�Kl�`~�￹�=�\0 ��U%�'�a.�f��j�h���!%l�G8 ����)���\�kA�<ѐ�Ct*�q��h���S٤� ^�'�Jـ�9Pd�[�����o ��_�{��{���
�߷˪�A	W/�}���=�,��5˒J�������t^V� i������u�Ԭq	ʛ�´�E��٪����ui�:��'�G%����{������9+Ev*ݻ\���`Y�˰5RS�9�r9 �n�B���*b�,����z��W>�7����W�<{���gӀ}߾{�$��� �)w51:�u��l����f=�=�{9�ii&�2�l���~��l-���ws���}�Jِ �w����u�y�αcySu�$p�������^��M� ��۠zaBf�O�ڳ�Q\�Y�4qv�s0Y�$���v�r볘�4���g��_��ܸMQ�7x@j�)�༓�y[0G��l���M�x�Ǵ����y[0��DDp:�7*�4LX2TK-{��� �}p��u�/! %)H��2�rJh �0����*`�
h	����f���}�s�{��U����/��9@���o8�K���`��b�^S�$�� �%#&�	���UՑ�w�s���^S�$��y[6��ֵ�;1=L���ѻK�M��jGT���,�g�#��-0ݶP��N~��v���*�ɺ��0�˽:�9��{�/+��{2�߼���-e���W��{�r""y4�� >}x���G��,n,���8F(ݼ��0����#��$�� ~N~�'�9&�ܶ� �-��ZKZg�*���~Ϊ�߾�}��`"SH���Ȅ��+
�s[�������`���ܷ�~��{?䴵4���o��;������D�*�쫲r�'lCb���0���[�pv�M��/7��o��A�,�V�J�{3ٗ��V�����r9�j�)�:��3Q�,j�[�����zIi g�.��|���}��>IkM��cGƁ؇S�Uwf }��^���#��(K����`�|��e��l���~�ͳaI=��V��r�� T��������"��������`m������׿�m��i���m��s�o��T�B�ST�%AAUV���`kZt88��P\��~�k3vf.��4k@��soe�8��FZ������0wh�|o��Xfj�,.�f�"d����Q�&%���gF�Y��	��nJj�.��n�X���GutcPkCHKz46��o�Ʒ�s�zB@HM�
�S.�l$�Su7�-h4�#���2���{�7����kc�әY���ޭ�!&��q�����F��hCA��6ަ���,"ll,��ٙ�TN����0ʩ0�a�Dya��4xb��3���[�����=�&�[ �:IdQ��q�۴����e�W�j�V�YZ�gHUAU]Uh��]R�a�q&��`��U�%2��z�y�Y<f�
.�-����j���Sut J�*Ś�5s���x兺�_DP�;K�=Y!��u�7I�������6d���[����z{JM�)���ەt
厎��y�ɻm���/�	{��w�����]��U�a�qk��0�ۤ����e�R��hm�Y����{qr݅:&q���%�Ln��g��<77n�X�պ�f��Y;)�'���\tdm��ě�&���v8.�t�z�>]���v1"��i�c�uk,yk@J�4��u�']XVT�D��»�\��{C����bxs�+���9&���;@�J��d��l����B4Z�ls�8���&t���B�s�;r��i�V�ΏG����t>Q��u9����>laK�t񹅕V�I������>�O�̠�x��t���(9+��n`��0O��Y����5t0�Г��Ü�e�pQ&n�:��x�`6�<yp���!����t�@!�i�*+��{�9O<��շ7���W7R��GggiеD���q��u�Ó�`����7q��UV׺Z$�Tnn�֮��#x�ݘ꣈Wu����F��{�eM�v�d���҃=�v�6�;��fy�л��8ȅs�&�Xy��R�v.r�f�N���Sv�':�����`.�ܩs���nݐ׮_GG��I���S��R��C$��۳W,��Zl��.�;`��ݢ .-�I�%���=�d
�P𶍃�����1;���Gs���,�0UW"��փ�Ca)��k-�҉ɝ�;o]�r�.���vy�Wn�f
ܦ)N��'*/-���l��,1y�<
�l�y��������<��V�g�۫�.��9K���s뛇����1v7\��zxKv98�J�&� �N���˴��f�.㞧H��u��&�J��p��1u���y�c=T��{�������Ƶe�d`�8�a@G�U;A���U�H���j�'J�?���j��z�)EM�D0D�C��:Ow�~�ߪ���]Ua玦�Q����S������γ�in�1�Y��X��m��Pg����wu8��I�k��;��������=���xxl�猽v�'֎���B�*8���i�y���3��y��7e�#�^��M�i��y��sv#��.��pq�d�쳺��n���G4�v��v��	�4�cu{s��'���!�rM(j|ߓ��ݽ��r}�ᇚ+S���q��jn�Vֺ�gb�#g]u��m��)w�;������0;����~�/��33.��;���$��L33>� ���މer+%�26���RS�$���O#>�G��&^���n1��&��#ݼ����	$�@�O# n����(�I�.d��4(��%��Y$�.�Z���}6��F6�Uu�B�w�@u'��@�w��{ʰ��}僃���R����T���Z�R��V��jI���z�ڃgu&5�����}����7S�Bʶ�̻q��������}�[��KI{=���F��,��ﺏ3߹��yЕ����1�+)��@^w�2�w��R��b���n�(�����{�w��a��n�����M���̎d�Ӱn�p������g�U�༓��nbf����nj�V�s2�k��}6{�g8 ��,����9�T�Z�����z�4�(�q��}���fB	m�I[U��zK�"����n�x��d�#�����?wٵ���4�������1����WAW]�`�_n���92y?�0?���8�w�ih��������
ݼ����U{�9�����4�1����
������]U�=���uG�pg
��f�jb���pn�ϒ�:�{���# <��D�
��$�"�&����� #�ԓ�<��� Y�v�u{Mh,�������r,�����]�l��!�lo�y�/��x����k�+WaE��օJm���:���۸��:��E� �u3�LQ�7Spv�y���	�x��V��4����Z��t�hٙv_�*���'��n�����T"���	��.�C�s��t�Հy��Ɓ�7������~lpH�)��q�-i��{hsM�8�[z5��cCYeY1M��%$����ʧL�X.�T`fVA��f�& (0��[D��ְ�l#Y�u$�#vٿPS�M��J���������:�msh�/۠g�{�n���V^�~QwA��g����!��#\�uд�����^+��#t[[����|��\���U���ydȼ���%XW�� �ֽ�h�E �L�,��w2���l�ʰ��{�u'��^N�n
��.���˸�;):�=�'�G :���~������v�J��́ޯ'�|�D�����;=�J(��n*�Q�����ͭ�~�{6�g��`M=�7���ȸ�G9�ɟ��Ȫ�Vi�����A#n60�Ԟ��܏]yŖ�����x�7!�v�#�v�N�a��Nr�-�TM��cBv��	ٻң�C��m)��k)���&s�3�Grj^�l۫=r�D'����ӗ�qΎv����ty��)�����hڎԉ��׃�����z�<-��N6�v��ρ{\�^��#L���%�u+�mr7AUIj�M��\X^�7D�K�H�OgM�[����ѓ����xh]p�+��#qGl[ ����q����%�~��9����(�˃�.&��
�ܛ��;):�;��Jـٗ$����yfd݄Q8���l�m��R�`�ɑ�Vϒ�=�8��#	7�_��|l�̻��Vԓ�4�����.�&n$��f�������U�u$�@�V̀�=���ڪ[-���m���"�:A�'��Ӫ�ƛ�wW%�~�����}}�@������ٜ I��&M���#Q@�1GvI�w}�?.ꠄ*���V�?7������͝U�{����4�����f�ΨE*�:����y�� $���+���'�i��S�ҹ�Yf�}�I��}v?w2��/�@��Nc �5(M�ԗ�j�2��@;�� 9ԓ���� n� ���w�p�Ճ����\!�Ϝ�A��T+��h^ݹ<��ޣ4�v�nZ���T[���WxROtϓ� �n���4P��>I6����j%&LD�w|��*�&A�� :���K���\�p���d$v͂�2�����亐�ĦeXY$,Q8�@B10beA��2�S��FF+!(�pQ�C�9��?{;�����`��ɸ.ʊ����2s/@�ԝ��Ot����G"e}��� /:�s.�-E
;e�?6��}��Oc� �f]�s���#<��	l��ʮyu�(l�u��Q�S�ax���+�v���������ZƉt�P��� ���-�wٗ`��,����0���$>B�ICi��]`�w�J��	��+f}ȍi�>+�nC��������J���`i��IV]UTMQqs1\����'�|�� �wd��h� ����"&�&2� -i%�.s�����w��VQ�XT����Jـ~�DO����� ���=�Y�Ց��JG��P6yc�絗"X�:'2n6S��A״�.�9��J(�� �I�Ѐ�R��({�y+��{��IP�-��x�ٗ �I�䭘 ����iL͔pXY7uw�y$�4y[0&� G?{�`s;�S*�*��;�[0�;��W��G9�8o���r3���WTr�l�̻�?{�t]�}�;�}�|����B�E$"FZe��dP�a��
F	� �@�y���ٰѝ�ѕ뤎�=WXF-�g��m��,�pbB�q�κ�s��N��̛�� �]����؋<�v׹�LBd��h��	�!d�S�����2X�%�A�,�e�k����q�G.�������طF%��Kפ�,�<�T�ghr��:�+Xw"����u��,��=Jָ��aM�0��y�5�ƀ�Hk�)ff�����/H�@��e��0�4C�B6wq�3)q�>ٔk<�wZ�GV@�K��� �p-�v������������+f ��X��	V]L��J�jj�k����s�KZM����}������]����ڤp�#vK��=�l��:��Qx�Otw�i�:�t�J�����6�����{�{�ـ�C.��j����d�րw��@I=�<�� Rۊ���&�R
HI �Ґ@E$�p��F�́bN����#a��,��i��G�{ITM]]�I=�<�� ���hl�Sr�>���?J%'*AeI�I�������P?�Q����_�꫟��}[o����=���m����!\�`w�ԯ ^I��'��������,��2����n����x��M��?����n68GiEue�`w�}���#�K�4}�׀A�J/ ĵ���Ԗ�2�R�+j��h3�4�ZID�yG�����Kll���c�k��n�����j&D��
g��� oR��������p{����T������B�w�;����A�۠y'��ޤ2�.梮
�e�]�Sw�v��?�KIf�?��`�6���m�������#��O��r��8�J�*����'��TXD @w�T��čj��`#��Cf]�GH�zl���X�5�ރjn��wN�`r`E��M�ޑ��r�h`4��M	
�2L�Z;1��a��#U�D�"� @�b�X�&��ɠ"�(�G�D���u�i4D{-o��-"�������	�� @U�ݢ��"&�,n�F�a�3n�:w:�WZ٭F�Y����#�0���%`ܑ)yЙڒ�h{�hd*�Q#HM5*4�N!�1!5�n�z�������ԗY�;�{���j�,�5�6�c�n�`:���vvc:�'!ں��&D�ʭ[A��I���� U�`�P�$����-�������1��I�H)F�K����|������������ӳf���fv�d0t;pt��t���`�0a�a�&a�"4l Ѡ�f0�Dq|?��~(� QCIKT!UB�
D L�T�UM*�� �� �������(?�A��C�=���Ȉ��n7������T��uEP]qWx��r9�����# �K�w޻�{ы,�d�Z���^p$�0y�����xROt˝��秞i8+v<O��T�Cd���n�{����z��g1k�̶8��-.�F $������ROty�� q�y��X�- �9ݼ�e��kNO6����0&� ��ʙ&*���/�Uw�u$�@����� ���`{�~k)d����:ݳ��}�O������U���������%4�L�S�GB�C�m�>� �cO�[����U�w�����'�|�F�R��e���B<����G[���:���5�E񲎝7�q�^.����8�.֗\W�����;�<����y �'x�eT�U��a�n�6��g8��6��3=�`��]�$�l���E�[�7.���.�t'�F 6��o|� K��m�[M;j�B�V��7����|�� ��۠w��d v<�jBJ��fl2�.�̇���K���'��W9�7�_���
P�UR)%z�4��&E���TH� F"H�3�D�e
h�2�����ShA� A�3I?*72VIc���k�t{Eo	ېMC��
����k�t�K�l�:��݊�LG����7K��Nz�l7f�l`#���<��C�P0F��}r��$۷<q��FY�=/)Y�|�_$1�QL��>�t[�Hfɹ6��7$7W
����o[��F�5ˋn�l ��7�K)��V�O]���� f������
��&Qt\�#e�B��z����wv�vi��|��i���a��:��&f�4S�^q׵؝g�l\�xd�.��n�/�>���|�F 6���#��|�����Ie�W!n�� ~ﲭ�7�x��^ ��� ���扛��WU ���@w�W���:�K�D��ml���ke��uv����'=� U��@����� �쪥u�1�j��^��{�9�?vf=��� �k�p�(\d�]MU�]UE�r��Z.�jY,���!�س�銫0��烮���))�ӕ�B��q��&c�3�/ �k�~��"#d_}�nf>�ȮM��-n�Ͱ3�e����A�֑���?JhY��:-iX�,��0XSIϐO}�޿=Ϊ��}��rݙ�`qw�q���ͻ�;�Np����7X�|�5	Me&�!aJ�^��ZI<�����u���33�`~�;��7�猒����n�tϛ��D����z�:�_g8 �I?}����1�J�I���g��-uЗZ�Vmsu8{j�r�n�]��Bj'A�Yg >��`~�;�=�ﳟi~a�ﾛ@��|X��	Rݛ�ޤ� �{�v|�`[U�v{*�Qe]Q5˲����$���'X~�.-2�I@�7����k���\���ǈY�IPW\h��/Ͼ������ה��N�@iLé�-�UvI#�`c�=��KZI~��3d}�e'Y _��4�ˢf�BnFf;E�l�V�#m!�s�.��y�̖�U�_d��n'e��7?��ǰ�=��@��� rڬ�Jb������������M��I� 6���Jw��fg���nW�HG]���y�}6 ߙx��� J{��)���TM�*��� !�� �W��	&�t>_��9�fY�p23 �s ̒04��f�1�`E�ZG�҂t��I����cV����f� �g��@�ot�N�6� ���#���ώ��n�K��Ļ�tf��Q��E�`,=o�{�|�o��v�{a����غ�����~~����;)������)�:Բ+Qʁ��,����ǰfz�A���O`w���=�4��6�+$i�`�ڼ;>�����۬P�cdQ�F�	6�\���`s��� ��d�s=vg����*��u���&�@��� <ڼS'�Z�����hI|�|�>�8��Z��H�m#��8 �g���\F��k�:`�d�SÝ�������i3/l�
���r������N�\ړ�ܺ�K��8�ШY`�!TƦYG]����u!�A�y�bVn�W�C����!�
xŸ�q�/Eqn��'�qȘ[xq���9�����7S�l�%R�O�k�m��G�
U�@cs��a�����w{ɣ�wAѴ�n����R�v{8yR���(s�}�<)\�pt����(m@�S���):�6� ����=���w�mcl�V�If�;����y��otJn�{��.B���#2n�@�*np$����`m^?>�I�%��DꅲW�斴�~���� ���`@jn� �)�2y��U�)T�2����ɰfe��=�;�{9�?39i��-��OU�ќswoh�(��;S�1�9�b;h���D��e��Ƞ�f�ͼ̻���=��� =)��;�s3Uܕ35$iu��ySs���8�9͈�q�6#I�����Ͼ� �g��]��574�J�kws�{�=�=)���&E��^�M��~�&�a]j��.��M�w1\`�%8��� �yLÙ������UM�d y�x�IN���OtI����|��}�6�݂$����E#m�c@7X�`%u��7����s�����?����@����w����G;��p��&�s=v�?z?Aʠ8���s�{ɽ�#��� ��� ��S�s��X�*�pn�y�:���3ӫ��>S�9х���4Ɖ�NI`����3����Ϊ��~w�\����m��NH�a��$����~��8��{�z|�`��C���.�jf+�Wyzl�}N]`y���:�=-�����Rn+H�bc�UD�����ޟS��E��%�'���YqԵ�sٲ�������k�&��� ��{�z|�`��X��{�<�0m�Z@pN�o8 ���"9"��Հw��������G&Br�é�"�RKl�{�?~�����{�G��� o|�v��Ur�˝��� �S{�z|�`~�lD_""�

Ĳ
P��Fdb
j*I�*�P W�~gU}�3��r�'T-������9�:��6rw���/y��^~�8�c�'M���uc
�k]r��&����#����&P<�: j�%q�`K-�}�s`w'���RS�{����L�+,�&*n&����삪�ݤ��u7���l~X{�j9�|�|{�1�v{�z[u�yל��yLVAQ$�ĕrM����ot7l�<�����c���'ͩ+v�;m���\0:jp�))�=�����r#��s�Uy��cm�m6���m��������it��鬢���B���z>��3��s�sq{�z�;��B�R�:���$����*��E�Hgf��M��ִ��vkSKL���Ivy%��q�u�{�Р|M�:� I&�t8��{c���}�a{!�l���4$h����(���I�_x�̌�ù��Ljy+@���tQd� @(���}���>vYd]X�c�fb�M6��Զg{�Z��w����n�/��׫tEHCIU�aF����"���4�e�Ef`fdu�'rR^���e����i[%�Uq� ټ1a������t�jvX���MnC(���]h5��e��Ѡ���4���&My�6f�3�G���^���4E�u�RՌ&!`�%�v:��(ؔ.	T��Q�{��2��RAVP����j���f,�[tWJ�Y�y�u���� ����$��]��@X�D��f��S��!0T,�A�1L�@h@g.ir�]��t��M���N��G ܦn��"
��#���{=�r��PXG�geCIH�ݭ�n������Qu�E��o�O��5��	�U�
���()u��W}ؽB�&�����bof���yGf�@N]�*�Q�Y4�	�.��D�x<�ĉ �r���'��	aU�	�e��Kn��wtBq'��ao,phrc�p�L�}j �N�D���,Od�-UP��S[@T9�V�����7MWU+Sf�3��ƽ�����U����d�˺�;��$[��z^|�X��T���i�� b%�T���;��k���nzZB����\�n��^8�6嬤.��M�l�p&H��$�""<Om�j]9���cV�R��9zvN���p%2s���N{&�^�n��/;n�z�k��ǧ�t� �su-�ͷxCuի���[=�ak�%���űv9N��jnN������<����4����4˃�P0����S���ܻ�����r��,t㺵���0`Z��v��A\Ӝ��nwv�n�(�..usn�u��'M=�<���{I�<cֶ��q�O�J�{��=�[si��`������كŞ.N @t��c�y�1��cpN7#��Nx���R������'������`6�-aNN�<��m���9�O7R���z՝Zx��BL�9ڜK�v-\b��=��{����к+�:�ձaȮ`ꛒ��w�V�t�K��tn]Ȟ�քڥ,%r���sF½q������zs�5!��m�8鸞��˄;�k��|�L@�E�*�Z#��y��^��zQ�i�q�Lt�E��Qu���G[����l�8[��q���/;q���c�U�nC:�p���)ûoJc�/�{���t5�讦M�K�u��x��;��`5��ձ\r(�k���L�����ͭ�q���3�5���.w-�g�=/a�2��p¶�'e��On-=ƒ)��ȻY��}i�i7F��g�uӆ��,�\�I]�fs�g(�d�B�z����W�l��ڍ��6�lnή���v�
E��/��q�]O0�<�*V8Zۤ���)e4n��sq�nca�o[۞�B�]�vE݁(�1ˁx,����w9â�M��i��l�j�K$Y���k�v���s\�AwRCv��͘�ݬp�Yʀ9��mPs��E.��u��'����/��Sht�z(��hP� |�m�P8 �	@���+����E||T;@1j�
u[B�㡭^��%��E��mv�η�&R�x9�ޫt].ۡ�� �4�>͛�ԛ��:N��k���:��7`���ȷ�Y���]�H�̦��܊B�哴x�L�q�J=�,t����.ƷR���Oq���tcr\]cV���B����z�:�ܕ�7�)cnbS�kn�yK���3̎'��6�<2ݻGf�]G=�`��]��#C�M'n��;ߧ����{���w�ބAKJW9�ݹ�q�����v�f�M�㬧R��n���闢ðDMw��~�p����_=�^r#�Ͼ�����}@ma&�������A�M�M�`t���ҥL�]6DUd�`w����ͭ�ܙ�{=�3��b%��"��^p�o# � �)�=��� �&YvX�:��;V�ɞ{�ﯱ���n�����!/���15E�D]�{1��@�n"5X������u��n���l2]���%lnQ�H���6����w������p�Z�}>ǳ��=�M�&䰈ҍ8��w��>����J�
�h�y�}2 �k�8}^S�y�}3AvUEU�������A�MN��)�=�fs�y5�cj�D��NS`w&zp���y7�S�`s���̇`�U�������=���3�~�\6rg��?/�ɹ�
H'"n�wn{a�C &�q{/<B=��*���mn������dE��Z�u��fs��ˆ��L��֖��w�����}�ρ��
���t�l�Κ���)�'��<��vyǆ����d�;V���=�W����:�v}�`X���>r"9ٽ�>��瑐�1��.jn(����;Y:�9��� K�����ld�簯����8�ۅT���`o�{�u;f�;nt*np�#�~���&�S]s���n�zP�����\�^�,S�g������ ��m�U��I��mT`�Jpz{���59"
��%�`w!���Z֖�:���}��!���!� ]ܓ71Y5��uSs�{ɽ�<�9�=-�l�����(��R�^��}�9�<�9�=-����C�s�;�G"/�����x�	A��
�/8}=�`y�zlv{�`w�����^Y�-m7v���ң�%�B�1��:������f��E��J1�&*�adnG%�`q�zl+�)��Rot="V9�=�bd�wse]W6�+@^��.d�M�`
^zo�6~�<�!�Z2�Wk����p4�0ڬݤ�p ��\ML�TM����Y�)mV �^S��ִ�Ͼ�~�I/f&"&�@��p�|���k �i)�5&�@�O#3��U|#���n:�R.��[n�w4���%���ک�ݧ�]�y��8��n;���ݎs�Es�y����pe��ZN���/��w�t�ָxЦ�]*g%/�9�꫓��!͖��w Ж��Z�r��G.��<�k��/s>��#ֳ�2v�`kI��:��q�V^�3�ݰ�E4�wu���{vGB���jm����O"L��ӯ��+�߈-�Ύn5���8Lg�ې�p�6uI��V�lQ<�IU#�&������n�6�� �����I��<�� Rڬ�vT����j�.,�����7���3�)mV���{��>���A8����Yy�d`
[U�o�)�<�{�$��D��@VF�rʶ�g���g��}��p������+m�KM>M��Ss�y&�@�V�2e:jp��r=�����疺ⱅ4�
[�6]'$�ѷ���ˮ.+��y|�6	�}�	Q���1��7s�&��_dw� �58�����@�U%jD��\����JBII@��%@0�0�0�3�@@4���v�5���^s�yG�{��2B�%�Eő5rU���\��Jp/7[�y'����cE@W]M֡�����1� M'���`	ל�L����MM����U���|��ԭ�u�8k�*�;�:�-�R)*G-�Ѕ��6�1�1�=���,��t&�e#��^�Gj�2\MIrW�Ry�	���p�%8}��p{�x-�-`Y�rʶ��� �E%8����<�݆7$]��XH���' ���=��pk�$���R�)T��`��U4H:�` ���i�H�EI�[������]����:����
lm�*�㖻^�ﻙ��z�6S��@�� Q�T�b��b�.�t$�0:�}IN��C��7�$��t��x+�̼&���N&�Smv.�EhdԽk�췚�C1��Muq�yל��Jpu7��y���M�4�C{��~��{����y�y'��uR, �>�U]uQW˺����{�y+f�^s�o�'�0���EH�+eer�w޸lK�}IN�Ȏq�9���}����㲀��[M�םY6;;�����[0��D��]TRS2Q��hLul��"�g�jS7W��1�I]�
N`N�V+l���ݜ������g4�NDs� ���`�D�5TLQWsW8��{�uRs�z_�`����1�)+��m��@~�ǰ=/ΰ�yN��@#�d�.�d���"h���=-��7��8�	��:�1����AF�C ������=��&��Cέ��mV�����u34�ڸ˪�Oc��X���<&��ؼ��M�Sy�d�pe�,ܕ�m��]m�ݘ��Yte�=���l�F��v�+���u��5u�Rj7,���lv���m� ���[��ҫ�^�N��-sO]M�/d��F<s��>�{v%�m�3�x��ˋN�
^���^'��{L�]��1�C�O��.:�g���yx�{i̱j�x�{��������x4'Eg^�+$���-Ќ6J#p�駮ߢ{�}���.����zWeq֍Iud����=������3��L���kIq�}=�`}���T�Z6�%�^�T�9 y�S�o��py7;�=���%XHG$��̙�;��=���T���ܲ�.j�袢����<�Npw���t��y���]�~�r1��G,r��ަ�@�� ��� ��p��uESts��h.w3r������I���.�8��1����m�Z���]]�MS~?n�l�=-��;���m�G|�*y��[23vkwUy�����qA�U*�Fd@XSC⡂=j��y8����:��?DL�R��.H����"jk&��S2��$�������:þ�vWCR]X�6-$���|w@O���6[U�wԄ`@�n$"�VV6VY/8}����zl���;�fs�}����(|�-AܚnV���:|�m�pZ�<����u8���RT��Kc�V����}�`~﯍��/��Nـ.�r苨��d����YZ�78zf|��ʛ��ښ�;���{�@���;^��}���Lǳ��D��1�m��M�}��~������C�qq�00�֓N���Lp��
"br	�ӠɈӂb��޵�5ظ|���{;:� �m������Z"�L4ae��։��R4�tH@G[�!ք���U�D�K�Zk�!h�Q
�~ǗF�J�E{��*AP�J9M#V���5K#䨣H�Q1�'��l��Z0g���r���ްMXQ��YҺ����ɝ�CD�bF�ʙ�ׅ�^hq3}GY=��2&u���r;�zr5u4$�-�w��F�h|�xu�7y�� ����avN���բtm��
2Li"h�663���Wp���D[6�:�IQCIIn�܉4m�B_	/K$�F����$lߊ�T6��Ѭ�c��*����]�<�+�@l:��ڀ��}�>PЉ-%���kZ�����S`}�_��;���DMPǗ����v78��X}IN��}�� .�#�x�C�LN�W�=-��;�Jpy7��6N�h!�^ݵ����!�ҭ蛤���7"���^m����x�ٱQ�&���'��0y7���'9ȍ�S�ΰ ���ӗV9M�����>Z֓a��|`
~���+F�P�&*ɂ��I������<�� ���  ��{�{�a&�P��q�)�;�<���]U�s��_��'�"L��Ù�`�ȍa4i��с�F֖kI_��׆����?璸K����ڹ�#��0�8������# ���}�^�E�B��,��&�vg�k۞��g�ɽ�ۧ9�]
<�b�q*�B.(�����=����u��y�S�~������2ؤ�ֈ@���8M�g܈��;�|��}��`	4�~�DF���d"7$�!:;V����`u+F��s��m�����F o|�a3u7pD�ѕ��y�ed������-��Oc�a�y�Bj��$���|��	7��2j�� �U� ��s�q��ba��!� �����~�<E'����Bø3ջn����P�)pN�7��0�uǁM�y�x.8;^�'/Ӳыn����!�]ۄ�ԁ����mFSu�S^���\�N��.U&*�ɞq�<���1�����q�����#٬-�|P�C���䏓����=/Oq�;<y"�ƻ#n뉒'�礹�OJ1�.��<s�.�;u��i;m۵b��P��*�K����[{ڎ!��e��R�U�n�]]9�k�胢u��Bh�aJ�eU�n��[���G�8��F�I�ԭ�!�䠙eVE\M�ATU]��I�ԭ�<��{3kh��y�Z�*�����n���yU78z%1�Dr���M����-'�/g߸g�m`T��Jрy�S�����,�.��@I������Z0����ٽH8Iv�.��Br��n��wAOt��7Ns���t;z`n!V�qi�������� ＞���o�� }���;#�4��_ ��p��Ե�֖��Ds9�L[y���}w�uSs�zC˔�6a4�"�VI��}�I�}�䟦c�������f����UYv^s&G9�G%�N �_}8�h�;�/�@＆�I�)b�n29G�?zf=�Į�w�OtS2�9�;�LsT�X��g<�e�<�\秧x�V;��;.R��:�,rWD�ȝ$�V1>n�m��e�`y$�@J����0�K*
�����B[e6����}��Zl̟|�V}~6�z��%�i����V(��H���+� �v�?8��@D""�(��)�I�*���O�Ȉ�9�����?�_�@!y��O�T�'I+�}����o�`w2�;����ޙ�`��2��Q�	��p�[0w�78Z�`r#�>K�&���w;y���:��lI�@�gn�g{]8؍�m�6���N������6Njـo�� k�ą+eU�����Lǿ�I&�{��;�l߽�ϖ�M����9�l��J���p����V��_=й�ǰ=��yc���	B���}������t�����8��"(��$4�h0t�b-�ְt���Ii4�{�q����E�RV��ޯ��T����X�������f�ܱ��1�6���;I=A��`ۑ5j�J�q��ÂHm������;f ���a��%1�uy����h��8�U��l?ٓ`w��xW����0z�K�&�5aSY�u�R��8�7�~��"&W�_� ��}6��޶�9m"�V�^������<ݳ S���DDJV��y:�nT�*�6�/8s.���߾�"��s��^}��;��Q�&J�$�?Hrb`l�������Y���ˀ�:����p���`^;`�>��h{������i)䃣rl���&�un*�&���].����]��#g�̗ ۭ���!��nps˸�^Pї��!M�M�8T��<<j�6x;��6�m���1�v�h��!�n6�Tv8ţ���ȱ�&�)�A���K�n69Yb�u�O8n�H��`Ԩ���y�l���s+�2�	�Z�����I������
�6�x�9tJ]Y֦9�=gY8p��ܻC�:�9��y�d46�v�ثԃ���?��l�{� �����Ds��� ���?]HeD��PF�]h	Ss�s��<�n����0/}��;�\E�SI��d�� �&��)�f ��U�dJ�N�UFWE@����ˑ�>�&��g��=����y��܊4�4�r�O��ޤ� �m����=�X�v��n�m���nN�*�z�9�lbi-$[���vƸ���X��}��%���wՠ$�s9!�������T� ;��KH�Cr��)�?{39���i-~\�EȾ���������92~m��PZ:�VF���ߘ}>�k`y�6R�`M��=	@H�r⧕1TM]� �%8�%8�ot>�9/���=��?�l%#��96��f=����h	��`t��G9�s��D������ ���Es�96NjuH�(!�n,-���y�A�7.X�q�W���'\��{���6�0:Jv6Cʑ`yN쉺$��@���@wު��ӽ{�gq����&���\Ys7q�u�S�{���:�~O�	)b�fT�X��uk��������󣪮����̱6�Ac���ɘ�sٜ��2fml?�������sl:�fKH�-M�yd���&�@�����=�78�{�`w��/�",�ۧU#��R1B�����1���K�ݸ�@\M���'a�����n�QuS37W�m�d�IN �%8��9�:������V�-[�=��� �M��F}�DG"d^���U�J7P��|��=��{3�33k`~��=���~�m9*RJ9\�4��m�`�ZS���9��r"�I}�kKg������ַG"�j,��6�F�v�p�� �I��Oߕ��.ꓓu׵���(�p�j����k]��r�]b񲗚'� ��7G2�0t��H$������Gd>��0�ϓ����:�c����1�������k��>��ʡ��	������"��p�n��y��*^{?{�Du��#m�y�336���ɑ*Jp�{�z��$���E�U�����c J�� ��{�f{6���y>��@m 6�`߿����N��aDw!�ߤ��Zk]z)�AT'mf!����F��e�Tfm�ARJL�[ƌ&���VDX���cT�ff�grf�Ѣ.�뻾�%�@�Bh�Ph>9l~u���a�VY�w��L3��iԑ&�LwQR,Vؒv�ۡ�����P^.�J��z�c�-^��!q���Q�B"��]`���V3hq\ ĩj^����"HY���FKq5�z�mw֝�u�E5#�1E1D$D�A!]�-$��f&Xt���Gġ�ؓ�v���a����a���z� H�C< L9\>��}��ӫXc]S�"
e�L�f]kE�w!�;�����l3���у�ԛ��u�����^���J�84��`�Wu$WF:'�g�Xa%�aoN['��X3�sZ�>�$���	(h((�X$�+bI�%+F�������tE�]i�z ʃ!!j�J	� �&���������nс�u�9""ۍ�5��}=ctSuca�E�	�!
���&���6E��U��TUQ$h��1��a���Y�a�Y��2ݔ�h�)�ш}˸瞀��86��	Z*�������sMu@�[ڠ��a�"�X1j.u���&��ez�:ؽ�L7)��l������6Ǝ�ܗ*��a���%.��)��a���{�t0�����_lYcfY� ��95h����P�f����Mԝ�C��$�q��a{s���2;��v�)�g�����i��}�G�������}�	l�Ǟ��ۭ��O�x��%��6t�z��o�Hs��Ýnz��$m��t��Ƣ�zz�㖻d/:�-KTZ�징��$�nni�<��d��v�G	�[wm�!�tB`#\���%of�Tc����g�}@�u�a��ѹ뙜cn���<�/t��77��v�\��u�
����a�g{&u,��z���r�	��k����Ʊ��v�|\H+��"� ��.�6|�U4��a9�'�M * m��P���r���s�}nsi� (=�9�볅���G�d٘���6b�b�iW/A�AV�9<ݞd6�������:�e.� tg�M��4���ts+Z�l"�ݐ�`ݬ>R��u'$���4a���چ�����Up�[h�;H�a��*�NI�p�*v�6�"�2��YH-�����N�#7U@:���pA]n:/Kҧnܡ��NѶM��<�l�Z���٬]6�֔dF6z|q�c�Zfa,s>�Kg��]�(���Xk�r�]T;��_q�`x������n�BI`�Ge�|���V�E�-=��ԦC���G�nf�&��k�����C�ݠ�;�-0�Z>�[b6C��g9b� ��Ѷڼ�����,�ݕzM����p��F��;=
��=V��I�[�*N0ƣ�ٗ���˔0�M��LE ;+K�o �Q7Kx6@6M��9�p�\��;�.Ÿ��먖���;!\B={n%��ӭt�픥�R�{@��c��a朻aطG � mr�e�6�� h��-���X��-hݍ��I�!���s�k��`���f�o_�_U/ʇO��(p?�!�N׀���A4
m����+���w�o[�Z�kFN㌱���q���Δ�`vu�(�!u[t�bF G]~mv��M�}�ǇԻ��in�5��E��ud��;G�S\���s��r�<m����5h�c�m�[�6Nl�R����[ڶ춃h�bDy�nz^��{n;f�%�{�f^���X�V�����r���
ۆ�d.Ƹ��l�$�9��S�j��D���ێ�䛒�oQ�vg<~��}��v���
������ϴn�(�� �t�nk��N
}��F��)n�$�ٲf��+�r�@n�~�����u��s'|����##�'%���������k�"p��'?���&ML��bn*6�Ye�����k`s'q���pu��l�� �DMMId����ـ%IN��@m�0��<�,M�Ye�� ̙�`~���p̸l~ˆ�h�dj��%�a������璲��v�����{����(��f����A�أv�]��w�g���p�0��p�������~ʚ���I����9�����z4�̱$�;P� � �N����.���s9����Ϲ�?�%�ً�4����TT�1�E�?w��%IJ�{绠7M� ډQ.˂�&jn("�l��� �\'�t��>KKO��<��<�1��9,�8{�{�6�s�w�يdU^S�v�	��J���HV9)bq+&���U�aӇg�y�p���뒁�%�vk��u��]�U'8{��`U�?s������s�6'�0	�UFRZ���pϹ�r9"t����}�t����D�%�w���F�m�X�VY�p�}��y������L@�0���"��1 �LE�IX �����/�����:?z���޶��`�v�Q�߿7�t��L��3�.ה�ޔ��*����e����{��=��|�?fg8��d"��S���%T�8gU��.�9�g�+<q�L1��N�+�����TvE���߲�=��=���fs�fL�6g��K`Z���
�S@~�� �Z{�7M��v��R�m�9t�-��߳���3���lzw�`~�����EX�Wc���9?}o��;�� P��p~���8��-%t�^��߽���0>VI$�V�*�p�`	W���Ot�9�;�`,�M8��+����V+�[�r.�^Sp�n�wA�n=���(��_���\	��5�h�s�w�=���0�`��@Pq�Ґ�VI���?*����|�����|����^eB�T5h���fOc����6|�ZM�Oc����8��'6����@ŕ�v�*��i�fe�Xj&=�X�� �����7[?~Y��
�{�5�]��������V:ʎi����Z�z�<<H.yo�|��&t����L���;0v�[zT�|ۋn��e8���m�yݴn��KB�:���!�+�m�Wns���M=n)�m�3F�yG6���hΞ ��d�M\�W�:�f���S��I������"zkD�<Ã�M�;]�\��o/+�P�&+�n}�/d(6$r������Vze���t!ѫ��йt��5���DYWJ�!���5h�l��4]v猝w,�O�K���w��4��T'�g���&wa��+S��o����{�9i��v�J�����ܖF*�B�/8<�M�-kZ���~6{&����g9�Ii�־���򤄊U$ŕW1�w�_� �%�w�'�Nٰ~�L�n�㬢��Ӏ�˰?u��Nف�Dr9=���yT7u!R]Ma3wX{�q�nـF�ۃ`u�ޛ:���[X����(��I�6y����ã	�:�����[77dkP&��G+mZ܄V[��e�`s�\7�ο{�`w����f&)6�,
��rS ޻f�O9@�7U�$�{�ue�`fbg��U��K���8rc���{��s��o���:���}	Lq�������;�}�p{.�ˆ����=���;�u�au�[%� I�0��u}��78{�{�{�ߟ�ބA˒��훝���坻l)�4g�����i��7k�m�x�[�5+��lz�U%8z�߹��7��S�ﾓ�݌r�૖�{|�=�`w��n���`�l�=�J������� ���;֞� �y~�bGy���ra����l�b�j�  P6՞�o��~�ǰ>�יB��T���p�VF�v�*�܉����t�}�I�m�b,6\pݤs�O��s��O���p�\6�/�Yi��X5m�1��v{�m��Z8lD�R�	��:��4qX[kl��-�8d�{���s�b̸}�?;�~6|�nA��6��w8{�{�L�}����>4��<��:�Ղ�k��33k`/ߝ� ��)�7���m�a�E��܍Z�[��ִ�߷�ٞ�ǰ;߳9�����J���A"3-
%V�洒���|��=��; 9k�"��.�@p�;��M��7�����kO��516�Fj5�@�}��[\&�n$
ݗ۳�м�vj���KJ`\�jxĶ���Wk��}�8{3k`s�p�}�����y�������[��o# �;f ��V���߹�L��DQ���E!l��������}6���9�3=p���d-��ݰ�2�Y�9i������l������� �c�H�URK,��w�� ��� �;f �yV��b";8 ����R"�������k3+1n�<t�	�>{��Pu�fU�T����`���^+]��q�K�D�����鶖�PM���$�c�7y㊞(�s�w@���b*��]�L���dv�
��|�I:�OQ�ʯ[�{��|�݁�ی�d�\�s�5d�^k=u��Ō3..�<�u��M�Wt8���3K^6�xLD㓈C�"n�67lW��`0�[�S��^�E9b1�4�u�Þ{�Du���s�m3�=s�x�. �BN͖9S��&XA�_p��_�`s�p��*�;�7���vEU�ՕuS%�V`�`
W�`�ot�l�~�G����H���c�d�w���S#wl�=�l�#��Jꦨ����� ���;���;f�f �%�w��:V;jv�y�32�=�l��*�;����9(w1Sfȑ�l��eNmY%	Bj۫�(�:yڸD�ocY�*�4�d����v��=ܱ`z}�V�� ]����m�SR6�8�� ��ɿֵ��ZZ֪�9��G8s��������pu�3����&���"VFԒ�.�w�������M� S� �<�U�UtE�U��7X��0>J���� f&��Z�eq��lvf=���V������ <�#��i���`�g$vC;=����dAgsV���jK�����S{����#��
�7N癓 �Z{�'N�`�l�7�S4L�qP]IuM�`�Ot��;�l���������#eN�ڬ�[o8�78z�l�� �� ���	]X�=ߪ�b���>&��Y��BZ�tӚhII�QQ�Iw�q�*��9�>�܈����BL������&��k�(ds�u �kFA�Hfâz�4�b��'6bl�7�FhՆ�����m���13-�8�3%�v-��P�J�����\�N@m:�8`t��Uz�x`@Ku0�~���YEQ�F`�6��y���+=�f�!Z���F��5�Jn6���z���w��tO]���ֈ)
R&�Eb��s�f���)tG��B����5��Sz��ᇤ	P�5lm�BK�̕^��O���Bˠ�	i�`���P��@�%��֤�"�ȉ9p18uoY�b"-�rbX�����Xh!  d�G����Ն RKd��.��^=�y��#�UC�΅B�1���^�4F� ��`U6}ąO�����Y��h���FoH�K�Sv+���D��M�K�4-
j����un��B�Iv��<����`��y8���qeǒ�:��=q���soq�nmnѭٽ�/K^��X.�ɹb�*����}EpU�@~P:Ҙ|;�hUP�b�ib!i�	"&JH���T�U|0G�W�v*����}�溫󟟜ﺽ��2�\	n%"�O����'Ww;$�ݙ���������`f/���6�FR��Kn��7���`�78���/��R�+��ϥ��Y�r�E�r��
+���x��i�6D���&��UM�`�ot):�}M���r6A�s&���|�d��G��/8?{&��Ss�)�U�v;��@�T8�����������}M� ��V������`�ܘ�bv��Ywk���^޴�@i[0?o��3�<�&b'�92fN�g�MI%"a8ȡ(�U+�?|Ϊ�潿5�f�ތވ*���{�4�����OR��-kZ�e�jH;I.�
�c��%�燛���va�p*�:F�k���kb�Y,q7E\]�z���8��0=J��-.0�~Ϲ��ϓFԩ���#�����""&G>n�{���Rs�fy<�Y(0�G[�p���`~����Np�;f���(�I���&��������Ԝ��l������w��B�Y#�l�s�gg�̐��`
|%8{��@��9�r'��gM�4:ێ�+�de������]I����7#��"�Pvźâ@��W�V�|��y6n�8�1�Y0uњ����sf�g��t�\�=qΛ<�U�3�1�YY�����Yx���}���\#��1��]4�*n���n��\��{j&����\fm�hJ�ۮ5�q�Pal�<��B����Ůغ���ᇎ.�M��HI$B@�x �P
B�O�|4�7\f�y.�Ÿ%����:
�&�z��Kjf��V�=t�Ju������v��*g���t�l�ｖ(�eN��Yf��3�1�߻��y�o�����i�ٕ�[i�P�E]D]�������v�z�^�;�eq�`[S�������޻f	zрw�=�N$��"�&&�h��� ޻f ��F���ݙ3�p���-i�-�X0��F�q�:���r$�D��'g���m>^&��oV`䉫M�7U4w�h+f��������w.���0�8�pp�J��=�;��ш��L�Y�,"qx;N��5ε�^y�����~��`w������4���fM��v�$�0���3̨YUuWutE���{��R��;�7�@9�ɰ~�I����pV=���������0��`G9��Bb���P�-���J��n�n%�c5b�^x9�r��u�|���nn���F��3���\���۠&���-:�V��d���(�V�Yo8f\6{&�^V��irr�$���*&��n���]U������:a������	��" ���h�*� &(���?|ﺼ�s���둖;,e�8�vpɘ�g��2f=�ǝɰ9�{�7!"r���8��=�?s������;?/� R������H�E�BЀ[c�'�;Bc:LW�<O.wh�Nλ6�Z٣3�YH�����npu�8��-�^o���b,��d�S`s;p�
RU�g�����l���Ӌ�bj������Y�9M���@j��z�}H�p�	�����n�0���W>�9�Uߜ�.��<�(�)FJ�(J��*"J�*%� �i	}Q:��}溣;�쐤��m,���p��{��� ���i��9��*>	���;=��W��[=�kpu74���p�g��+c�U��J�ju�,#&����~���^������r;!���0j>>>���]�ET�}˞�?7xz���p��3���M���[����F������w@m[0�� %�x���~�K�4�/8d�=���l���0��� ��	����.�,���7�ـ�^޴�@r����N��F!�9X�~Nv��i��<��v��k�vޞA�Nm:�5s\�z�Ug�s��<]��<<t����8���j���G�5gzaG��D��.��o��o��e�V���D�3���$�Gj�Ȓ��c����c�=�Nϱ ga^���q����;��WUtY��dw4���#�A��T!� q��1�l-��Z��6rT�����O�(
�
t(U
p�?����pz�r��+nwY��!\��2q�W��d��C;������m�k+韭�o����i|�`;�`�"Q��n�I��M���Ot�Ӭ���w޻;י-*��I	n�t)��7�ـ�^޴�@��b�������́�'^M�{����fg9�̓1�uf5�YuU�9�W5��x���t��=�n�����n��-���TM@eJ:�i����M��(gyx�9�v\Omn:]Ú��5ww�{����� �:�������,���K��3��KY�N���i�?t8�lJ�cD�����R ly��A���� N�w��@��p|"�f�戲j� �:����m� Ǚ�`�r<N�HQ�+w7g n�$=�����`}��}X�1�"��(��Yn��{�s�c�ɰ9�1�?��<��r`FI,v�R����pv��k�1Ԝ;������K�m�VPM�l�6']t#��!o8<ɕl�&�줫 ^�{�&ܜ���..K����� }�� R��{�����X������$r�W�1�d��s';�b�J|��D�y�s��\�^��p�Y��R�r[f���>p-��i���J��`�asRU]T�]]��[u�k�� R����g8�KKـ�棰�j�B�V�=��1�8znl\7��wϴ�O-";u�;׋1ʬj�,���/�����6u����py�6��#���mҊ�u��r� ]m��X�y�}ȉ�<��Q;�U6}�� Ǚ�`c�M���zlA�b�U-�FKc�%]^�̎[u�l�ʰ>J�-����0Aa���k)\f�a��ֳT�!��f ��2a�I��200ѭV���(kZU���/������UeQFIf�s�*��)��?7���`��Ƚ����Ts���r��&��ZA�n���{��7Jőn�sq�W*����� O���_r9 |����1$�Q��ٰ=���s奦ϟ�}X�_^ �%X���9���j��`.l����� �� R��쇻��p�=ben9h��l>ZI�I}X��`�7���`�¡���R��E���o2\{��������_�������ϵ�_���������TE\��PA��W����� 񷮺��h�� ��� ��������� ��$(����1U"����"�$ (�ʪ�H��of�D�( $��(�����Pp�	QBP!DbR� :�W% r 1�H (��(ʢڢg��w��A(Q���k�����J��� ?����E?�E?�D����� ������QM���
 ?�?�QHР�w���'����@������(��(���
(��(�Wh���'���� 	���������������O�����o�������TE_�v����ӟ��������UDU���DU�����j4'���k��QS��������������$�`�$I#������O����������6�i����ύg�g�q:���D�7k�b(.*�L2�L�H�2
C �J�$�"��� ����ʉ0�Jʉ,���J@))*$,���$(����2�B���,(� ���)(@) J�B�

@,�� ��B�($��*H)�ʉ�#
$�ʉ �
J��J
�!!"JJ��#!+!+!�H��,��@J���H�$�JJ��*�H�	 ���*�H�$�@�� @J$"�+! ���!(2#	
�#!
�"H@�H) ���HB���BH�$�BJ$�@H$�HB$� �0�!$$���� �J	(�	���!*�@��HJ�� HH���H@$��HB$��	! � B,� ��(����(��*�!*��"(B
���BH�0����+	�	"(H�	"�(0���� ���(�@�	�!(�� J�
�$�HB$���!"� �J!(��!"�(H@! H�$ ����(�$*�$ � J�B������(�J	@�����(@��	��"BB0��"H2��"H��	*���B�!!*$ $*�B(H�@#! $!0$�H�	(��J$�(H�$	JJ2��2���)	K!,�,�2���! B�JK� `��H�(CI(L�$(D"�R���5����?��/�������+J�6�G�s���WY���������O���%UW���g���ߟ��Y��G�k����3�?ן��UDU��(�TT���?������gv������TE_�����x@U���<�� }�?��i�<}��* ��P���?�w��ч�����>�<Qc#?�������*�*���*������D���ઈ�����TE_�ED�W�3��ՠ���W�g�<����:/?������w�a�s�c��}
���+�+��zN��O����|:@:%EOo?L�^��������_�UDU������ �{��{Qp��M��_���3������e5��I�`^e� �s2}p��QS�݁EP�PZ@-k2�Q ӹ�R4d"KML*�^څE:Y�hj'���hQ�!�4
( AJv�t��: 5�Jk@Sv�@P:Jh�F���;t4hk@�  ������    ��=:�@��j�(�&���N��nxګ�7W�W}�U�Z�Y�}���P���j�#vjv���o��=�_l������{�<  9�����ק����|���}���=7��x�W�W#w���׽�^�@v�@ϟ-�A�ww\���JSB���x[��zzP<�zsz����N�>ץz���@�� �����o{��y�w6�s��ݹ@P)�{��  J]�x@�`�Ψ�罽�((���6 ==�� ���=4�4=��:��O{��S�z�4� ;��z=��(  
�� ��rY�W]��j�o[�)_{���{���>��O�j�=��m��-�@�Í�y����^Ʈ��@�ނ�{��� {����0>��F���ϐ��w�N�� ����{{>͡ž��}��h(_|{�u��t�`l���������>{�������2=��na�n�3`,/m�tx����< }�;��y7cC�}��ۡ�kz�u����8��0������C޲�9� z =�y�u�R�킀�Q�֡����$�����<���
2�v6���wXyv���6y{������^� <�/}�}��+ϻ>��A�bL�����c��}�F�u���oA�      D�&��IR� �D�*���( �3*RTߪj �Oi��{R�@  S�j�2�SM�ɐ�"B���b��}����/������Y�>��~ϵ����
��w� ���AO� �������X ���?��$����sw���z?�H3�fyy_-֍�.�{��1X���I�������2�'F�P� Sag����ٰ���aą�L��[&�1��ba��²��٩�3g!M7|�\��n�_G���E�{����k/�B�fV�ǯo�b�	��]��u�k�ܢ��2��5�߾rh���\���P��ǉ1�5�����B��+��6���D���{+�Χ���a���8V�mw�wo���R�V+�x�QW����iZ����*��}Ɇ���p�)Jc���y���ת�t;����<6����-Vs՚�7��K�	����Dn��M�F��zI�ӷ���)�;�;��6��B\����5�!��t�&�,.��<�,��n�B�dsVm�t�z���7�e����>���>�þ�k4�@]^mf���eU���:��1�
�
����CԋHI�F���y��%M�af����b4�c
�K���0�����w��.�k�^xn�߾�59���ZGm�ӿV0X1I|���Z拇�����rsۼ�e1� �t��
a�q���NQG
��W�[��z�Z��=�V ��!�A�H��{���D��xF>H`0:�vߟ5����-��f�L��f�P�ߧ�&��q/%"8B�t�|	L�+ܵǕ�o�,5)	
�$��W��+/��i�kw�9����xK3�`IŅaB1� \���s��rx�Խ����%~�u_N���R�T���{~.�<O�f���_��\��a�233D.�ؕ��Q�=s8k��4��!2Nhن�n��`I�����aj��H��v��Lۺ������^�ˬx��S�o����{�'��ef�fdM^r�XK�;�h��y�oVo�X�ff3 �}ٓ������a�q��ὒ��qy���jˣ׎�d)s[�ߒ�F�zh�7�����%2�,)-X̉bm�z��(D�x���S�h8�2��f�92����C�$�tB&:�		L31������ᤁ[�ב�����<c��]�~O%���=HSz��h�b�)������t��~��3��z�{Ǔ��ᴛa�ԲI���BB�w����B2t	��:��=�oS�#�ĉI�0�	��^���ą�б๋�T �#&�yy�4j<�@�05�B��!8�^Yo.��E.YW��,׷�^���
����~�T��jt�3��6��ͯr�^Y�t�߷*��ek�ݻ�<��N��].��ꫠ*��;]V'��n?z�].�s=U�O;�Y�W�w�8�����;�N;�pW�޽���E^W��^�]{j�q^�ݧW�Å)�}y�U���V-v�Y�R���z�/����=t��𻝯w�n�8U����~~Y��W�Z]��_|�(����F�9��2�&����|�*@���u��p<��-yN�r����������C�C�=G[&��9~Q��ޘ{LϏ!:���٢n�:ߞ��o�~��
L�.{�c�|��l�y�a	��s�1��f�6ƬK�W�L��y�o�%<9=�P�d���7�04m6�Ca�.h��.�	��a3�VMS	r�E.X7��'!����J`��,��
@�
��K��K��pϲoy�Z��cj����Z�	RKh�+��+���VVr�ߺWd3	A��4�����ā*dY0ٓ~y���:�x���s+�=bHXd!�f�Y� BB��T���\%=�
�.0���!cHX��!e�(d),����~���<�i%(s���ᴃ,ry�D�'�������<��hA��Hh1ه4y�g���fb��j�gx�����iw=��+��?>p�8}���4ٰ�v��wa_���t�>�JE�'�h)�yOo���>���ǜ��u�FQu��Yy������TPf�}��-�kI���Y�K�o���p�]������_��JUB^�����Ȝ����s���x�bh��$����]�S�-��zx��
2��*��,̅�af���<,�at���(P��+��t��:U��/[���k�I��I��SS8灻���B��YYp�F�a�aB��M�$1%㏮�g/9ׄ�����!,>���x�_��N�%��0�5RC!�8�!�,X\IC A+.!�B2��Z4F���,�o=�{I$��7wv���+
��uu�Vc�]�{®�ݾ��_�S������fs���ם뗞�]��[���� V]�K�<o<��'�Ǟ����������
U?9:[w�w�+̫ ����fQY��R����{�y�/��q�o�l����Ѝ�o~k�(��J���ݺ�,A�]+��y�HwK9uv&�{G}Y��w���y��w8W����J�U����}�I?{r޵[J���)�!��3���{%Hz����y�k�A��rՃ$����_�3�r��'֡䯾�x����w�j�_�WY�>��(�_����PP�1T�)�k��M�[���q���V��͑���)�0�Y�J�),޷�Pݭ���t�Å+\
�]�YA��o[�	����]�afpF�I�M������Vu�o)sw���)�
��ow�$�U��ⷉ+]�=\��*ԋ�.�ݣ��9�*��M��8���An�V�֕�}ܦ�,t�}�3��p(��ܣkǕ]�j�}�;�#+�]5c����x�j�<�ַ�������W*��i�?3��hр���4W,%��X^9 w٦��w�c}�gޟF?VD�{$�pu�m����/v|�z\����l����cM!�d<�<!!��B�̜�����VJ��|�����L���\��.�zy�{=�C7�*���g�{�j�g(����1�%��O��+��g͘n�K%���;%�����*��t��>B���	f������kN�1�}��C�>}��ά���)�3�ͥ؆sR�4�iჾjy�rkwm���FY՚:�QO���k�{ù�����Ev�tU�u���VW�E)�஄z�)�᭲S�0�
a3y�g������:�]w=�G �jz�]U�vnz�Ψ���s��4�fa\�J�XU��~Z�WxS��z*\��s)���+��kz��A��,2�M˦fx�1�F57���6�c�t;�������/]ڬ��J^)X����*���
�)���]u�m$�]ٰ�=�@2��D�\"\	HX�F�#y!<��h�<X�b3[�OrksP�W�]i%�9dɹ�%/ ��nk�s�.`^k�x)�ߞsC
��of���Ja�kNs���{�K��7�o��y�$I�˚�<�8{㎂^C[u�r��8{函��T+�13f�P�T+j����Q��w�O��nS�QJ����u�7�/�H͞Ʈ:�C�Jr5 A������[�Is��.�f0����)�,��|�3[��2���nY��ކ74!
!%8r���)�{��v��U�.Ow�/�����n��o��[�Xd����əUV�s��U���ﲊ
���w��ꢪ�+������.��)�$1c3[�z��80�<�p4�ɧ{ԧ����g;~������pV���e���N����w�wZ����QG��_���{��WY����Hy�e�/��!������R7�f��t���6��iÐ����$HD �
B!D�K>3̚OH�`K@��:)f�s�WPok���
Un���:��������'z��x� jGi�T�#��	�\�8���%HBP�_9dO-�d�	HF2a�\� A�#X#`Vd�0�W��Ip�[���pHŉS  �HR��}9�P� ��g>�Itz�޻,^�!�s��i9$�q�r�]xj�sF1��eI�1�,��!r`JA^����U�)s���?^�=y��:f �tz�{ܤ��{{W���"����M#h����L��y��q�x����⭺V�?+.��ޗ]��%^�y�V{w�[��L����yn�\�d.��wj���k�ޢ�׽���{���xۿ��א� �d��7��F������s���4��S*�Z��Gt�WNqr�,�{<��=EfWk����N�8�^��͵��n�3����|���Vx3�qͅ𙙍����B�1���5�|���Qӎ�W�6�(���ee��T�p=��=����]�Q�Uׯi��n�%�M�@��fb��L�K�J��,��
��p{|�%�;���n�<�[U׭�����Yګ1�8F]�`kcw�|����Bs9��6zY[�=��Ww��*��͔�Э�S�R�0���n|l��
sl�Z����F��w�K�.\��z6�ha@��P��e9�?a�N_�6J:=r����K�.i9�A.kZ!7�ߏM��|����u���y��+Uo1�\8U��Sc��������8� XGp�r���<֏Hz��4�ח������K��I���ܑ%�ї+��,���g��*��Ӌ�.�u����ݬr��+��mv��W��D��ݔ����m����79��!��I6k��hAH�i�ἁ!���q�0Ұ�5�޽�;���ͪ[ۮ��3���
�b�M�o/j�{=UE��߽3k7��l�U��z��.��r��)U�Ｍ��W�>�v�ׄ)��8��<�CHl6:$!LuLv�y�X����YS�]��o(�y]���Q�'{�;�̪T���WӕB2%�%�>�e�?/Oܜ���Wv�=��y�Qu��������ͭ+��i*�53�]��3ςG�L;��ݎ�ۺ�
��ۥ+=�x3޳}Wy��QH~������z�.�B�V[�jΥꥹ�o�y��%0���og=���y|��M>l��d�R�'�/�Y��^��d$������@/~�l��84����f�Y�2�����%�q�ω�ٗ��d�=��h�������*�k����c�ĉE(F�=)�a0%�.{��B���7�F$�����!	󄰲B�t�B�f�,M; #pf�Rs<�mzަn��$�]]Q�z�z���n����^�Cu��ڂ�^R����\;tm�<��~8>�4z�K�F�]s�������8C5�s ��.��9���i��xy9橽��6��	aŖ�e��l�tp�U�*����:�^IuB��r����zY.�.n����W�Z�K��Ќ�@����!�&�܌�7���!M�+��g<nxk�v1���4ąH�%,�|i�}/�}7��"h3f�槹�޷|�Jp$�~:͍)�B](drB���.��Lfe	i�(B���d6��c�g���	�g����hRʷ������Z�k�&�����V�i�0%�X`OIy�'��g��YxK�s��J`���4l�Y��!�$�e����c���2�uҒ˱gY�:љ�)�.%*`ap�==�O�硷Į��*UR�4^ҋ�U�L��$�\��mʞ����k� ��#f���ذ7�[䬺�@����q��z���f��T����{��s~j�w^a
g�<�o�`n��\�g�_HP����p�%�9�[�i&��y,9���۽n�(k��\��)a�v��7RPϧγC�Jou#H��ў�璲�0�.B�7��7=��Sf���2�t;��;�&��Y��)Zڡ`���*fL��I���<�6n<	!JY�6���*��V;�Uv������C�{��Wz׳[�����W{tQ��iU�u�VS�<�߷o��e+tg:���V��tR��׬��-$|w�nsfnS�-20�P���\��9�!�!��_��g����/,8I)����UUUUUUUUUUUUUTZ������������UUUUUUUUUUPUUUUUUUUU�_*�������UUUUUUUUj��
����������������������Dlr��;�Dn�Tr��������u��uqHa� ��bէ�*�E^� �BY��oR�����L�*����4�HJ�؝�U¢�K�/�V���g'ge�$At@AF5S�Y�6/�E�8�m�V�[Sh��QVЕ��&0�F�]A�:��U[]uW��0�9�e�0<
���ؠ)�{N&|���v3t!�;������P۵Ѥ�R�	e����P���Oz�l�dskJBX(�W%�jf���w��Z��q���NXv�B���:�\��[��r�8|�J�팛a�:��«	f�B�m�9���ª�Ӎr��uյ�
��p;ګ�r�c��ـ3TsN�j�瀶���I[={�A۲8�*�nGD��@TÝ9YĖ�v�7#�9i����WBax	ĚAl���8޳�xF��`��0n ���
L�D¤aL�����N��WYEV�k2.��@*�Uu[==ilv��g��\n� ��i5k���k��"��PXעL�@�9P�qѓ�#Y�x����ge�;B܏7���욞�G�hSq���R�xT8�%ck��]���5���:^=�A���Hp�#�U�2Zs�\g9�Y+��T�v� ����h(��� Ү'cm�[\����1��h���vv
�'Km�u7P���줩ڶE�Ǫ�Y��x�+lN�b�/%˲�ٛpA��r�Z����H�/�t]�.| ����j�tR&Ab�T��*ڃ �f����n�llr+d-���lܹn�@l;n�PM���h
�s�E,�UUUč��.�`wS��0w��<�t8�HU��8��X�NMe㴎��Um����ô�*F�P�ӝ)�쭈�lC0.,Ԡ����ň�:oLd 5���m�ӻ3 3��=L��cI{35�M��Xj�3XZ��u�m�n�UOK�t�ד����z8;kyQ�.q}�J��n{N�����C�'v��8�v�U�3����`g�n�cu[q��gR�&dR�d��`���:7A�ہ�U#�U�tmR�%�[.�Kv3j*R[�$�0��űK-Zp�ʱ:M��6��j����N�2r5�U��YV�œ�G\�lU�JQC�Ӳڽ�A´�xc��U�8�'gjv@��o1��x��qK�E��c�K��Q-:^�M]+@e���L2�\�#B�y[m���6K��� �8�'l
��QP0
;k�P媪�WVG�Ռ����j��J๶Լ�"V���{&���ʺ���f���C0 ��Ӣ�Tʪ��v59��WUM�ܗcUUU*���*�UvUX�VUK��tu1���^Z��
��j*�Z�I)ʴ핋U��%� �+.YMi�3��E�A��U ]�-Ce ����]��qX��)թ;R�u�C��ܫ�j��: .�v�U���[sm@�dl��.յW9tl�M������Vt�J�<��F�᪮�X��@UP�Ic��^�ڠ��y�K��ʐ��,�%w�UuRҥ��nں���Gc�j����6a�tj�U��b��K@��^ԅl@\6
s�����W���c�UV
B42��m�R�g������k X�X����f�J���V�j6�I�m�Wo������T<dx�j�e�_[����: z���R��v��
��vHͮ9W)�UU�r�]YnX
�:��U��v�CbV��=jB��L)����B�8��#M'\n����;rn��Tn����g��72�!ݶ�y�)��j�c(�:�^U��EF�jX⪪ݺ�WfU�g 5��m�8�! �;v��+@$յZ�57����cV����<����#+��-ЬHʱ��s�����Ƕ�nQ�v��'^��5A�0�VS�b�1V���$l;���[y;O�k2����=6�;���E;9Z����[]Qu'm��B��SqCO��Q���T�m���h ��e2L���K��++W]ej�k�:�:ֺCi�@�y��F0s IuݐZ��n�j5��y!V�6Sgvw��D�Y�`���{
f���L7�A}��`K@��[UJ����>��m�"6\+�,B�\�qP�U�"��l����^�m9j���{qnҬ��!��[�ڐ�NݨkR�U�u�c`��y�#tV��U�U��mKE�� Wi�핍���t�
��yb�56�(�[;��UUUQ�����A� .z�(;U�2=��j�k����'�jT��7��rM��If�#lae��m^6��fU�@#a�m�GOA��j�A-l�j��2�Xsq1e���3*�����O�sp@�!K�����J�cAĜs�M�L�x�Q���X�X�cU��F��+�Y$�P��6q�Zt��Z�5�iy�W%�\g �4t9�Ƿl�հls�"�f�����I�n�K���V��AmUw:np+Uҳs���N���^$�h+x��36��5��:׀P�f��m\��'S��pv+�z�s��.dU��v���y�����U[<�+WR���&Ih�5#���5;�� �i U�V��UFt���q=YB��*��+�t֠�j��7j�U��lvy�tP�K l��UJKQ��맙5#uK/����Wl�V���kT���*��M��U@!�ck��b�)E�a�Tj��PW�$�UV*�eb�K���u�U@UT�UUU@PS#�RV�Ì�I���j6����[I�EU����q��J�S��ٺ�x���r��U �Zr�~}��[���6eUUUV�%x�U	��ɰ�_*k�v騇,���A�#f��,��ҩ�֨�ݹ�Iz�<#U�UUR�UZ����j��vQU��\�uJ�0���n�R������mUUU�[���7R�䥨ڥ@�5]U ��*������cV,��ԫUPqW ��%1��j�i@PU��	���dtN�uUUJ:����)UT`V21PH�gM��u��KjӰԫuT�;��mA�]R��u*�d@�ڥZ�@�Ѻ��Wj�ڞ�.ZJ�EUP	k[WU��F��U ��R��ZB�	��Φ	��.�&��	�Ԏ�T$�iX��	�G��Y��eX�X��j�،�u��]˦�k�����9UZ�ڪW���"�UNK%��8Ů�UU{�_+� �y�^���T����h׭����U���Q���Z��*1�91�E:X�@ Q�>P9���v0����l�����)0���[f�!2˚XH%��f%���lc��LVY�PJ3\n�;SkR��J�axp�/b�Yi�Kaf�Y�Z��uv�AB��.)nx�T��y��܍.���UhX��^[��+�WC���d.�������p�yX`M���p�fqz���ƭ�uH�Nu�j��ؘ���3��XZ�R�a����#�s	k�lݳ�ӎ�T�ct�lGZݶ��kJn�)tf
�!HG\��c	�1:*u�n�hIQӍJu�QIң���t��͖���Ғ����m�$4#P�� lA#Uׁ ���-D<�M� 5N���@U�UU�l�jB�]�r��XHW�خ����=q�U���+�<,@-�J���� U*՛lv�j�i��'�G��ga)�W.���s6�yj���k�w��/Z�e��j�ؼm��jy@٪����27-m .�j�� '��`
�g�)�G8��媫,Y���xZn�'cUE�U9HHː.�VU�
�5Vj��y���ꪠ*V �ڡc�\�m��d��`��s�0T���pq[T�PUc����b��[c�jw`&
��S%U��8����:�)Uln���L���V��o�炱2�Zkm�5m[]UUV�)Jd���	$[vP�]]T�v@�����U��S��e[�M֦ۧ�j�'�j�����r����e���m5�F�����R�Gh)j]�J��;/t3��j�Uc�WnV'��>'�����L�1�Sme.em#+�UU]UT��r  �N�H��wgn��s�m�*�Q�nhGPY���UUR���u:�#�mzѹ��g�/`[0L�����&�yj����
�6�ul=8>Er���5$�t:ż��aݖy=v�d���NX��������|��8� �*�ؔ���� ֛�9�۷�i�o�M���xgoh�L��m�B�G�ʨj��@�e�ڊ%q؞����s�v��e�cf�0VC�יt���m�)�lǲ�u��K<�m���]t>�Z-�c��I� 2�je@x1U1�!WV3f�TZ�[mdR��ڬ��%�K��Qt��n�t.�;*qV(�n��Mcr4�BR1�ej���"�kpM�u/T�E9%��q[e�5/e�9%��V^}���Ux
��qt�:3�������O]n�\jrE_�_����qV�*�����Z� ��p��s5 ��[�v{f��X��UU&�Z��TT�ɐeuq��&�UUU/<�W#
2�MJ���F)�1V��qO�5ur�t�d������lh�շ�������k�B�Um�]&XU[H&����j�0TUTøUV458u�e{<�O5R�Ak:��5ːv��U�ɝ&�떀�0+�v�����!����ݤmlPl�[�V�U]��w�[c��,�=�U)u�����zS�������y(*��旞9��C��Uc����PY
^�Z�y�����,l�jk{�\n�፵�V��뉴0�%�mb��t��N����p�h�
���	� C舾"bD��Qz�qB"	�pE�"��B��U@��@���@J
�qH�|
mv(� ���>]�UD1"�Qڂ�A@ـ��(|$��<@i� ������ >j p 8��i�	�'��"��CDڟG��=QM��F!�|��C�_���W�?"'�.�⮑Sj�OE~O %Ex)�>P�!�0=P8"G��*��DH�� �*�@���!�E> ���� �VqU�J+�࣊����(b @�B'ʜ UU�PM �ʂ���$ "F22!1"�)
BXH1FDaE�X��a$B@I�A012D�T" � ����$ �*��E4(@}W�_AG<��F20�!�IB`H0d!	H���$��1��<J p`����1S�C�U_�<QP���)#a@�P��!-�Fʕ)%X���F1�B6�Z�j��I$kb:6栋 b	��|����Є�Ŵ-�BA��%$�6�z�OLa`�@=���c�D��:���#�E�CJ��Pb~Q �S����@^�e�~*(LH�DB+X�LL��^�����wI?�m��UUUU���V���U�p�k�ц"�+lf6�45wm�S�r���7d����@�tP�,ȅ&��4��fJ�S.���@�����\��R\к�&�.ܸ�-C�A����۲.���Mϲ݋��r���gkbP�ɜE�LW��b`�H��#ʇdB�r����Q�)���g`̹�u��fY��.�g�L�m��aY����8&���uk���*I���]�r膔KMq"�M.�S#�Z37MtZ��cD�e� �<v�<k��>�nSs�;��̈́4(!U�b�"�Z�1���@t��l n{th;��ts9\��؅�&���ljd������q��:�l�[�܆焨3C�v�Nu�e���Y#2��y�Q��i��$H1�iM���B�J!1�4E��۠��^�/m�]�gN98�]�`@eڻ,+m�J,&�)��k��m�pgP\�B۶�q@r9�g����M�Ŷ�#�.$k-��zL�ٯ�Ƕ���1�U��ls�X��%���S�p��[pq��0{u����٦кku�֘������x'�5=�E���!:��V�E jǔ�;0
KOr�u�mR�pb�� �l6�@::ɑr�'�G ��ãh�7l�9m�Dl�(�]����j�d��v�Wm�����糍
�5nv�H�a��!!v8���9ۓ��z�j�Ԗ��6˝��[v���e���N����_ �kaB��t+,B6�)��L+u��>xw��F;l�zd�����+q����+tm�cKkd톹�t+��@3����F.�u�u㒹�9�J�*UX�M D�;KVg�b��3K)�#-3���w��'(�ɞ���KB碤��K����0�0�!��f�fT�M,�ؙǃc8�\�۞�qLf��V�؁�3-�N����c���2V�ؤ1�M3�!-��lAW�<���!�FJJM�ػ6KRjЫHBY�LZ�֔�B| �h/�m~U|D	⾠�(���WJ%�����Lϲ��g������jl֮�\"�5�8�Fq5�&�n�t���r� k���6���,���C�lh���l��&n�6n,�Y�\���!�b�IxI�1��PMXZz��H�;�i�$��rk�'��{pX��{az�jZ�<n��`[bVV���&+��uhP���P��;u�;=����jL%��5&h��fYf�)5�+�;:u���ġ�6�u.!����\n;.�w��.;>�(g���B��V��M�L�I����7<���@yd�����S���0��2�c��X����,�r,}�+ �Ң�[����m��{���Ē[흮�$�^�x�K���\�\r�X��=��n�o ����@>7�7��~��۵Ӧ�kR�]�n�$��l�w�%��+Ē]�b�RK�����O;�ͳ���t%mm��X`�,�I��p0�S$uk�۲.n���<a�+g1���
8v�����M��_�{���.�$��gk�I%�2Ɛ�o����Ē]�b�\�UTE��9Đ
�jZ��B�pQH�I ��5�$R�+!,�_se,IV�Pv������fn�o�{�'��|o�o ��<ٮ��.ew�%�ZĒ[흮�}\�������$������Sv���[2l��o�v�Ԓ�{�I.��}�Iz�K�I#�>>��6mu�6�=��}�x �se��%�ZĒ[흮�$��9U[(����d�Bf��P��XM(!�_!��۟0��;q�9��)������;s6�nzm�}I%��ﯽI/\r�$�����RKM�M��S�:�q��cg{���-bI-ݝ��$�^�x�K�$���UT�oҺ~��K�E�ǀ{���r�}���7o��(D���v��$�w%�$��!�$��؄-�l�} ��t� ����@?��v� �������#�6��ro%ے_z�^��I%�l�w�%��+Ā'��z&K�ʑ�5�N[Fd�����'B�f仅�q��#e-%�fm�F-�����
��RK���$�흮�$�^�x {�����||��]n�`�.<I%�l�w�r����W>W�$���z�^��ǀ�N�6�כ��b�I%�9z��9w{?�bI-��k�I�,%����qf��� =�{��B�>־�v�|�߸s����@H1	�T�(xb�mS;��\ݶ�~՟��ی���c;�@?�� ���w�%��+Ē]�I}�II
ʼ�m�J-b8����\�cW<r���#u��ݡ�Zۗ�����h�Q�����z�Z�b�I%����W+޴����b �o����� �����M�I.ߤ��$��bI/{r�I-ٖ:6Ų��ro w�{�����1$����$�^�x�K�2Sv��t;�.`g{����o�7��x }�|�}��}�x {���� n�[�&x�Ll�I%�nC�I/�[�+�I/^ϯ��wW�x Y'9=�����͂o5K�Fq`GK�kBn����;���n��л
X�q�tP˦�&����)0����2� �6�
��r���Jpf�K���	��Fa��1�A%�^����]���.^�םA��1�u�;:t�BW7#�s%.6�Қ��62<�\���s�:B;=���V�x0��f�#V�әm����l�D�&��%�XE6�/��������`�1�vi[��Um֩�5�@y#q7$�y6��˛���\�t^h`y�+|� ��� ��yԒ�mK�I%�nC�I/m��n�Z8�EWo w�����rrs�c��~�Ē^ٟ�Im�˼I%�4.��"�"�]�Iz6��I%�nC�I-W�^$��!ޤ��P�aa`��ڴ�j�$�}��$�^�x�K�܇z�^��M�����3WW�6[�m��Ē]��;Ԓ�c��$�}��$��;����jJ@xf��Mq��pmW��:�ۭ�f{pV�sƅ͉�U�X����I����RI{f|w�%��-bI.�r�99������ �~�F�K���Y��[o�jk����! S �1:i*i!	])G�jBFI��`f���	�HBHDe��u4	B���a	S�1�$$դ �J����=�
f[u�o�|�߯��w���y�� n�ئ�ၫ/Iwې�RKV�^$���ޤ���n� �O�׺/4د6o�����s�.gֱ$/^ϯ:�^��w�$���w��Ͷ��h��.< =��w{Ԓ��~�_]�$��g�z��k��I/M��~�x�p����/I�q��9{t�Vz�1ۃ]Χ���bm�=��V{&�s`F�4���%�mEx�K�܇z�Z���$�o�/�I/\��ua`��mM�Iwې�RKV�^$���e��%4n%�����3WW�6[�=����<���.(#"��҈I���r�$��!ޤ���b��i4���$�ov_z�SF�X�K���ޤ��=��ߞ�x���.c�{�u�-bI.���z�Z���$�u�]�I_�{.m̬��c��1��.��eL�Q�AH�hk1+6��<ޛMm4B��o.'m^$����w�%�\/Iw^�ޤ��=���O�׺/6�כ��8^}\�r�����ޤ��c��I%����}�_�ā��V��4\��߿��z�Sm8^$��v�Ԓծ�$�揎�!L+k�}���=����}Ü��o��f�&Ё�Hv��W*�ir�����ԍR�A��+i��&��ٕ�}\�T�>:�<������;�m˛,��`�!�޺/-��]��!n�9�V������i�k���v� �� �<����l��7��!>��[0����0�̬w\0��I[�đm��;*8`ݙX�`wc�=��Q��V�񴩶`ݙX�`wc�;*8`U�b���ڡ��'n��p��ǀvUȰ�͛����Ou���h�)��LղW(NF�DN�'c=���3��jk.���ZщB����8����(gh �n-�c��Ѱ�.ǷT.²�щ�+4�B�)(K���*����i������Ú5�����ڠǶ�B�����y&{*<OY�����/��e��r��g�͎G��kl�M�� ���&�j�B�H٣zll��f�:� "Fe���hZ\H�;�������؛��X�+��P��̌�F�'���p�[w��Mw�L�m� D�3�WghM)����=����+ ����Z��+i
�l�o 쫑`ݙX�`wc�:�"|�
ڶ��l�;�2��p��ǀvTp�=���e�:Wv��X�`wc�;*8`ݙX�8Ҥ�]>'v;b�`wc�;��0�̬ۮ��N*m����fXI��iuL�ֺg��{f�d�R3���-\�,�<f��Pr�����@����=���UUs�Π='� �_[r��e֡��SZ��s�~ٵ8�@Ůs�#Ӯ����N�nժ�|,�|�I۬�\0����NwfV��Qj]5i�WE]7m�������&V��j�Xۢ���ӷm��NvL��\0۱�Ur����%��!ի��wh��.ТԸB�b�s���j.-��[Gg�C0�^ll���O�}��{:�?8`�c�7Ҝ0x��*�˺t%wwi7X��gܪ�) �>xߩ�`�2���9č��`���>'un؛0d���N{�]O��m��@�}%�yg9��瘄.�	=vPq��o�$�	�e'0�a#!b�Re���;�6�Ɇp��4���@� �@��8:�Zi++1��������3��e��u��ӝ��g�N��C3�_�Y��Z"�燴f�4H$#	�N�'���W!~�4)�}�hvk76����5��9�N;�^F��Ù�Zb&��aJ\��5�<�e�7���<$��	2��k|y�8��l��7��9N�z���櫘e����y��p��b&����SEĊ$�$p�;I�IK�̪�h%�Jh�8F(�H�D�1�n�����oZ��)�s2k'�^h9�d�
� �nH-��f��eͷ4��֎y�M�9I[�{��7��P�Zu)��'����љs�0�R�\[��}���]ƾo3��R]��1��a6�K�.�f���]�ki4�Jj���A���4	8p4�	�b)�b���j#��B	@��+��� � /�Q�`*�M�y��X�8`ے���VZ%v��x�S�ݓ+ ������>x��+v��Ֆ�M�Tـwd��=5� =����z����+I�y��<�;kҝ)ќ��Q��s4��m��ɧ!㺻��V�ڡ��$�`��ݏ �Jp���u��e`[�Akᦝ����� =����wd��=>{|�9�p/�bt���X�9|�����ݓ+ �� ��xT���%].�mS�l�;�e`���ߵ�0�:"x�
h� B%�D"@�PJ�2-G"l4Ic��>��뽕�F�΁�k�W�|�ߩ�`�t�����+�f�*��1@���1�b�lHik��AĲ����h�*���V��5{�x�S�=&V�{�%e���IЮ�J���N��X��X[��n�Ct'j�v�� ��+ ��-�x�S� T�m*�tU�O�bV��\0�e��N�p�:�
-K�ڴ*�n�0�e�T߫>:����=5�$���a[B�"��f	� ��$�bQȩ��L�s�r�3md�熱[Z���ۇv�����3�	s6�3�KZ�vܬ����u�B|2��lۓ����h3TZZ������ih��6�[����#;F�d�Z�մ�9�*$��sa.0�di���l��c	�ª����d�/��`lu�D�%��)���T�mf���m�\�J��J�c �`Cm���RXL��֎�5=٣���3$�$iW ]�� X�pm��8�pm,��g��]���'6&��tڮ	uX̹� ���`�ذMp�:�e�R���,C����6`�ذMp�:�e��N}A�Jwj�	]��m��\0��x�S���� ���	>]��ˤ�V��fV���o�b�=5� 쒲�Ltˤ�Wm��`�N��T�>]~�� �ٕ�i;a��̮r�(KM��X�3���v�#25�.�uC�x�Q�bz���M���,�\0͙_r�UU]A7�^�����wI��+m`�ᒹUJ��UUʠ=re`�N��]�rNZ�!��j���٢�:�}�+ �Jp�7ob�=5� �$�Cv��t���`�N��X��`�e`R���.�t;m��f�{�d�X�S��Ur����b�`�%���V.�7��:f\ީ�<�K��D�L�ꜗ]��J��-~�� �+ �Jp�7ob�=�r�'WE��˧lV��fV���o�b�=5� 쒲���ˤ�Wm��`�N��,
tW4�U.*�P��i�XF��$�aT�W�\��v8�`�2�n�C`�ݶ;LTـo�b�=5� �ٕ�o�8`vJ�_
���j���Mp�;6e`�N��,�r��E|��A�L˕��8��l���۷ ve8�����<�R��t�t�=Mo͏}>��7Ҝ0��X��`�Q)7aJ�7MZ�X�S�={��̬�QR���N�m��l�'�b�=5� �ٕ�o�8`�jRv]ӡ]ݪ�m`��Ol�������� �D��o_r���-ت�>2��� �ٕ�o�8`�"�=5� ����|���\EIpX��v���S�;N�X��tq��n����D�
ћ��V:��]Sf9g����?�z�X��`d��=��M�it�v��ـM�}ʤ�#��>�}��vTp�
ݭ�W/�+�Wm`��Mٕ�vTp�'�E��R�'Nӱ*�n�0	�e`�p�&܋�r�ɟ�����&�9v�Bwn��8`s���?�]d����0�B D�B )!��� #�H�a 0��HBOOK>2�g2h	"��e��s�-�W[d5�r�hAz;����n.ӱ�sx�� >l�M
p��ǭ�%e���U�g�e|�gB�����n��,"�Y0a��ـ%�p%���jUu!J A�@�^;&B�Y��QՂZ\j(�w���F�:���u��1U�2��b��3/-�vTl6�pu;�p�������2��N7���p*�s��NIɼ��5��l�]�f C��2�Z�3h'���xFP�lhJ�R᝺z0m��FWGJ�@�����?~��t	�e`�p�=��)خ���Wv���n̬���X�*,��� �ٕ�vA� ��� ���&��+WI����u������3� �o���n̬ۮ$��it�v�cf=r,ۮݙXd0z�\�i�X�ɛ�"�\���4E����s�뀮"�.9�h�&�O��'����G��������&���; ��P}��� 6J��mt-�r��߼��$��9�HI�0��DфA#���X�BHB��P��I$ctB2"��;2s����7�,ۮ�)#���R���n�պ�=�|�0�ذ��~���|��{���>_-��_0����g%��|���`�Xr���}���֞�Fku.2ށ���àI9?��}���7���0�ذ�\Di�Wo�6y�ysv.WAt��%SSq�T�Pk�k,6��H���3d��\� ���+ 샆�{�\�������jܛ]28r΁��þ�KO��=X��0�̬��I#�'N�T��ܹK��M�<�}۹'�������/:&��}ݛ�yߦ�7$��{%2_
V'�Hm�Ur�l��M�e`�p�����|`_]��N�];v� �l��>��}��G�{uà}�°�]`����;��ա��rU�j�M�Jۮ�s<p���e���S�N3e|׍�t[V�{��vk��ٕ�+����=��o���/�WGQN�ٮ�*�6O��	����*�=�|�}N˱եhV6�d�+ �l���s��ʫ����|��
�A`��wV��������k ��� ��}7'�� ���P	�F����s����:�{�F�&.2:���; �~��~������>��V��;:�ߟ)2
��eBk,�Ie{4N���z���|�kK�n4��� �5�ӗ��KX�n��V�1��{��0n�`�_W9Π��� &�+�QJ�>]��`�pϹU�RD��V��ٮ�I$�?xC��Æ�p�5S�y��{:d0���q/}s�l�� �٩TFY�]f�����r~�.{����'���� �����_���_��ެW���E�n��0�ذܮW��O����O߲��8`ʺ����Ӷ�̢���8Q�Xl=�o��+ں�Z���0��������H@!���$BcB M�H��(�����e�ɤ�e��L���d�R!S8fe����W[q)H��u��6���l9�g���ow��=��U���=<INY_o��L��פ������W�0����Ö��Jx{3G	�/��t��
�ZI`[���.B�5�\6B@��a@��)xeL B1�B�`��l�<Ѯl�	��ti�u�$�fT�s�#KOt��|	V����o��99.���H��޳�$.��r�RRJN^lCq��B��i)(��p���BW~1�Bm��˿����E#� F��F2g�$�5��OGfL�1��3;r�ri% xž^BYai��ԗ&�s	��Id�!�.X�L2f�5��9���{	$	Ng(��P��m��[�GF��	C]��5~w���3K�$?�
����n�m�c2	0���f��M��0�fB�LZ���E��^�>���>���g߼$��~~UX�UAV��UUUT �P��+c$�g�ج�(n�1:j`��U*Ye�3
�saL�q�TV�%Ѥ^�ݳ�"흓q���`�!����B^-��MfXlS� �����ù1�JqM��R9 �y��km�B��&�Մn�O`�n���TpX�f�b6�a�5�x��R�P��ա.e3- �&̅��%3�Z[*d��a������ ���3���0K�0R�V��s��]������g�&��z��ܓ��Ĳc<���>^��gu��b���M�&�o	�Nv�Nyt���KÉ-�KWU��+s��K�B��+5�8��l�SY��	��Y�;Z�u.��N�aN.ړ��i�a��>۶6������d�˒aFم�i�+E.eKrfm].��)���`*�M��E�Si���;��z�Ŧ���	��3��캮���n���t�etkt���	��4�[*T)�4̀�6��%�M3N�eqv�9��(Y��镄Z��k��#�'�c3U���H3��\�*�/j��iB�@���h�M	t��#{gB�xv<V�2q��Ak�av�{n]����T����
�	��I�Liշ1L��onJ�)�v݄��<�h�sU+.泂	�j�9Vqe-!�����쥋,�k�h�33YE����a3[[u�4�;���ݑ�zޅ�q2���@�ʥŜ��n.D$�?ko���cV�[K�TM���`��K]�L���Ȝh����e�EУ��ʙ�Ӭ�TЀ;����`)V�zӴ�z�����@�a��0AuN�l 6��R,��D�M�,�kU[�'�+��ma�8�W]��x����STļ\S����M��X$��ݬ�ԿЯ�ێs�M��]�k� �n9J�Z�8��[V�;pN��6G�,\�C��l���ۀ{	�9�-�v���*�*�M��b�[v5=l/�cn��s#�k�1t�Nx݈��C%,HVk��h8��7%45fjL,�32Jf��U@Ҹz"�U�x� R5A~SǪ|������*�~U
��ܤƟԭV��`#�E���5�6�Jk�4ԕf,ly�\�J�]֌�e�����h6�Î4V}���({�l�8�0�S$�a����/%5LYl[�uҢ����D��"@�s�wc:�շok�����n-�.u�'Y��݃��Wl&덬�9�D��d�O]��Σ�6ĲҼ)��m����i1h��
��,5�@���\�$�{$�y�I�o=��ڽ�ZX=z'���+K�E���]�%�[f�m�K4��ٗ���� �Ƹ��N���gyı,O��xm9ı,O;پ͊�%�bX��_v�9ı)���;�
�A���mY�O�%9)�b}�{�i�bX�'���fӑ,K�����iȖ%�b{�������/'~��ډ��a�eʳ�Oo!Rı<�f�6��bX�'��ݻND��"� ș����"X�%�߻�{<�����������`cb��b֦ӑ,K,O;��v��bX�'�}�ND�,K�~��"X� X�w�}�ND�,K���ٝ�%��5�5�]�"X�%���w�ӑ,K�C�~��"X�%��N�iȖ%�by�}۴�Kı;��-�љ��Պ����qv�;�\���ᴒ��x���qg��x�C��Qҳ�XE�b9�/Mı>����r%�bX�w�}�ND�,K���݇�`�2%�b}���;���%9)������20[�6��bX�'���fӐ��HA��	��� ��H��Iq,O{��v��bX�'���ͧ"X�%���w�ӑ?$���'��B�T����eY��Kı=����ND�,K��fӑ,Q�,O���6��bX�'�;�ͧ"X�%�����^乙4d�%ɚ��r%�bb}����r%�bX�}�xm9ı,O;پͧ"X��V ������9ı,Ow���Lі���[��ND�,K�~��"X�%�>w�}�ND�,K���ݧ"X�%���o�iȖ%�b_'���BV��i�R�ʜ)Tñun:��	��2㭑1DUj��4�S}�������Ӭ֍�"X�%��{7ٴ�Kı<���r%�bX����6�P )�L�bX����m9ı,O���ԙX����*)�O�%9)�NO��{{�� %�b{����r%�bX�{�xm9ı,O;��NAı,K߻B�����r{y�^B�}����r%�bX�{�xm9ơ邭P0Q$K��s�ӑ,K����iȖ%�b{�R|w2h�4p��kiȖ%��"�;�xm9ı,O~��m9ı,O;��v��bXX���t��H��e�Y�eRd`�3��' r|��Ǔ��p}��v��bX�'�}�m9ı,O���6��bX�'������r�F#30YLn
���c7k�e�ږ*�u�X�5[Xi4��>��y Z�u�/Mı<�����Kı=���iȖ%�b}���S�,K��{�iȖ%�by�;w��\�h�p�2�Y��Kı>���iȂX�%���w�ӑ,K��{�iȖ%�by��si�"X�%��{���d�4j�h�[�m9ı,O��xm9ı,O:w�6��b#bX��~�m9ı,O������G)�r���F��X��j۽f�m9ĳ�Q2'��߼6��bX�'����iȖ%�b}���ӑ,K� Sm�	�Q@N � ��H�s��m9ı,N���52h�[&����5�6��bX�'��ݻND�,K�EN���6�D�,K�w��"X�%��N��ӑ,K��z{N����]�T� i�],+Lh�2K��h�Q�)�I�6�d�΢�}�H+poiHcY�kVkZ�ND�,K��fӑ,K��߻�iȖ%�byӽ��,K����iȖ%�b_~g�s&�3A��WZ��r%�bX�}���r�B "X��?~��Kı>��߮ӑ,K���ٴ�D,K�w�/C��A�5���9=���/!SΝ��"X�%��u�ݧ"XbX�}��6��bX�'�w�6��bX�r}��}���f�7E�3��JrQD�=�����Kı>���m9ı,O��xm9İ�<����r0���/'ݗ�����қ�����bX�}��6��bX����{��O"X�%�����ND�,K��{�ND�,K�=���2�v���%r�ۚ�#!P�,��\� �b���0Ͷm�� 뱙[�m�B�f�3R���{�����n�e�m6셜��v����>�p��F&�N%����*2���'f��V�Ɂs�1�ɝ&��0Y^kx�9�C�ņ\u݆��.��O���-���Y�@��q��=�jcB<�84�b�1�Z�����5����e6U�X�l����$�# Z����:��)�$]x{Ol�������[���!�sSiȖ%�bw����Kı<����r%�bX�g~�l@9ı,K��w[ND�%9)���}�
dŗ2ܹ�;���bX�'�;�NC�G"dK����m9ı,K������bX�'�}�g�I$/!y���{��k���sFӑ,K��;��ӑ,KĿ}�u��K��߻�iȖ%�byӽ��Kı>Ͼə٢��j�՚�]�"X� 6%�ﻭ�"X�%���w�ӑ,K��{�iȖ%���u�nӑ,Kľ�ϻ�.����u�ֶ��bX�'���ND�,K��P=�~���%�bX����M�"X�%�~���iȖ%�b||}�?m���ӊ�'${��1��sJ	i�*�s��6?�u4𸺗�P��!�i}��msfk+5�6�D�,K����6��bX�'��}�ND�,K�����yı,O��xm9ı,O;�K��$ї2kh����Kı=����rT���H��bX�o���r%�bX�����Kı<���m9�	2&D�;����n��h�\՗YsSiȖ%�bw����Kı>�{�iȖؖ'�;�ͧ"X�%��{�ͧ"X�%��{���d���!5�R�SiȖ%��'�w�6��bX�'�;�ͧ"X�%��{�ͧ"X�*'�}�ͧ"X�%����$֦jd��浭kZ6��bX�'���fӑ,K����fӑ,K���ٴ�Kı>����Kı>ó�/u3F�[4�x6\=]��gh]��h=��5kfk[��҈R��n�I'�{Ѣݴ��&j�'"X�%��{�ͧ"X�%���o�iȖ%�b}�{�j�"X�%��{;��O�%9)�NO��1��.��6-.�6��bX�'�}�ͧ" X�%�����"X�%��{;�iȖ%�b{��i�(ؖ%�~��w.k&�ӓ2j�6��bX�'�w�6��bX�'���fӑ,pЌ�0� �Px(�"{��iȖ%�bw��iȖ%�b|g��ܒj�MY5�4m9ı ,O;پͧ"X�%��{�ͧ"X�%���o�iȖ%��9����"X�%���_��K4a�-w���NJrS����iȖ%�b���o�iȖ%�b}����Kı<�gxm9ı,N����`񨍬c�Ј١2���9�n]i7#�d\��GhJ���]dl��:�,���r%�bX����6��bX�'���ND�,K��w��yı,O;��6��bX�'��}���lѢCW.�֦ӑ,K��߻�i�#bX�'����"X�%��u�nӑ,K���ٴ�O��2&D�;�߹5u����4K�֮��iȖ%�b{����iȖ%�by�}۴�K lK߾�fӑ,K��߻�iȖ%�bz}�x&R�2���'Ò���$�����nӑ,K���ٴ�Kı>����K��W膀CH��,O{��ND�,K���3;0�e5���f�WiȖ%�b{����r%�bX�}���r%�bX�w��6��bX�'��{v��bX�'� =���\�6n�%�; Z�ў|��6��$3�arL����&�>ww���u(W}����,K����ӑ,K����Kı=�۱D�,K߾�fӓ����'�~��_p�G�gy>D�,K��w�Ӑ[ı<�۴�Kı=���m9ı,O���6���T�"X��ԗ��0�&fMh֬֍�"X�%���~�v��bX�'�}�ͧ"X#bX�}�xm9ı,O;��ND�,K�gn��h��2kZ�u�5v��bX)b{����r%�bX�}�xm9ı,O;��ND�,K�뽻ND�,K�{��n�Y4h��˩u���Kı>����r%�bX��{;�iȖ%�by�}۴�Kı=���m9ı,N����/f~�5���K���=�+i�#n-�����z��p���:�e��Hł�FЭ,��/�4	|Ul�ʄ�����qS�h��0��ڲ5�%тZT��8��Ԏ�n��s/X�`è,��sf�a����bQ�Rv�hj�d-s1X	��T���6T6e.��T�X�V������:���^���a�� ��c�k��bZa`�rNs�$�>|���gOQ���v{�].=.HL�L���˘�����8a.�'v=�U���ֵu�ND�,K�~��6��bX�'��ݻND�,K߾�f�yı,O���6��bX�'��w���M%��&��6��bX�'��{v���bX����6��bX�'���ND�,K��o�iȖ%�b}�|e��ɬ�5�5��ND�,K߾�fӑ,K����iȖ(�%��{7ٴ�Kı<�۴�Kı/�3�ɚ�\�r\��h�r%�b�b}����Kı;���m9ı,O;���9İ?�#\����xm9ı)��<=��ڀ�ɨ�3��JrS���{7ٴ�Kı<���r%�bX�����Kı>����r%��%9<��;��6��ݶVҹ��^�3]�V8��p�G���єIjJ݇BY�Qb�'y>��%9>����'Ȗ%�bw���ӑ,K��߻�h�r%�bX����m9ı,O>����f�0���7��JrS�����xm9A0� ����a:JB$�d
���#��{% � a�HDn�]�6Di$Q�(�(H!���DH�D I�ы�8(A!!�b��Q3�WJ��
Ȗ%��s�6��bX�'�>�fӑ,K���nӐ�����'�=秊-��%ungxr%�bX�}���r%�bX����m9��UW"dO�k���Kı?~���ӑ,K�����Z��]J\Է5usZ6��bX�'zw}�ND�,K�뽻ND�,K��xm9ıF�����ӑ,K�����sC1�S��JrS����}��9ı,E�{�ND�,K��ND�,K�;�ͧ"X�%�޽7�f"�fS&kj ��FF�\Q4ݺ.A�[@��&�m����&��oT��.�WZ�ֵv��bX�'{���r%�bX�}���r%�bX����m^D�,K�뽻ND�,K��;ܙ��˧%�j捧"X�%�����"X�%���w�ӑ,K����nӑ,K�����"~ "��#)��==��ƀ�T�3��JrS�������ӑ,K����nӑ,`��V�����Y�8nFw��)��"ky�g�Ӣ5�����Y���������$����$Hd$/���JH�$�"F���]ae!�j���j6l�0�0�	1Б$H:��7H�HD� ���!�Z���k1$7�x����Vk8@�a\��Vrq5B�s�_�a$��RV���,,8id#3��L�vM��ޥ2Q�B�O=��^RLiI$\� ���J����JRMMD�"1f�x��% �%eۙ	,F0�%�T�b@$�yv�	9u������fbZB5]h֡7�HB�#�\4)I�l��	��e�2���p�aCWl�0�i�I�Ą�R0��\5����mjVDx��-�b�x��E� �C�%�0�lA}�lD|A~D|"�*	�H5| �P�6lQ⩰S�+"X��~p�r%�bX�����e9)�NO}K���fHmuj�gy>D�,[�뽻ND�,K�w�6��bX�'��xm9ı,N������rS���������l3
�]]]�"X�%�߻�ND�,K���6��bX�'zw�6��bX�3�_}���rS�����������DV���^��豺3�J���
襷h� �s�@��x=ӧL�ޤ��U�֡\3�>^�%�b}���ӑ,K��{;�iȖ%�b}�w�a�A�)�L�bX�����"X�%�߿~�֮f�R�֤����h�r%�bX�����r%�bX�w]��r%�bX��{�iȖ%�b}���ӐD,K����嚚ɩ5nh�af��"X�%��u�ݧ"X�%����6��c�@H "w���6��bX�'�ߧ�ND�,K������J��'�����I
�����Kı>�{�iȖ%�bw����K��P� 0ȟw{��r%�bX�����S.��!��6��bX�'��xm9ı,E���6��bX�'��{v��bX�'~�xm9ı,O�����~��0�a]c�5xM��@ctWd��3��=����Vء��ӻ�]7���k .��6�D�,K�����"X�%��u�ݧ"X�%�߻�ED�,K��ND�,K�Խó
kL����h�Ѵ�Kı=�۴�Kı;���ӑ,K�����ӑ,K��N��ӑP,K���۳�j�ɣ&���Yu���Kı;���ӑ,K�����ӑ,TK��N��ӑ,K����nӑ,K�����i5�$5��W4m9ĳ�"w��xm9ı,O߿O�6��bX�'��{v��bX�'~�xm9ı,O�������C"e�r{y�^B�w����Kİ��@>��߮�Ȗ%�b}����r%�bX�}���r%�bX����fZg욳!�͗w�^Q����M����1�ݨ ڗ��>n�����f��Đ�d���R�Cl@�TA.ѱ�V����z��#���e�!!�&ezے�Yx�G�ݬв�P�nݏ[�\j�3FN Q����H�%ʗ*s�5�GnNs=�cY��V��f,�-`�*��]o1v�d����7��y���
ʑ��K�Mb�k�T�c�9X$cv������&�	��㚚��FLɭ�2+d��X���HFX�cYa0<1)�(�\���I$g{��m�v�fw���NJrS��濝�ND�,K߾�fӑ,K����iȖ%�by����r%�bX��;	�Hl�IU�r{y�^B�{����r(�bX�}�xm9ı,O;��ND�,K��}�NAV�/!y�����l�0��r{y�D�>����r%�bX�w��6��b�X�'���6��bX�'�k�ݧ"X�%��}K�i��E�.fL�ND�,K��w�ӑ,K���fӑ,K���}۴�K�@�>���������������E�6��U�p�Kı=�wٴ�Kı=���m9ı,O���6��bX�'����"X�%�|�^��Y30֦LMt�P�{lC��+�4[�nn�s�BG��v\�;�uuR�l��t�zk�^����ٴ�Kı>����r%�bX�t�xm 9ı,O;���9ı�����Y�a�]S)�O�%9(�'�}�NB���
"��%�0��@����bX�x~��iȖ%�by�_�v��bX�'�}�ͧ"X�%����&��kZ��I���ֵ��Kı<����r%�bX�w]��r%��bX�}��6��bX�'�w��r%�bX�����`�i(�%��t�zk�[$�N�^����n	 �}��6$�H����M�$@��{�iȖ%�b}�_�gu,�35��Rf�v��bX�'�}�ͧ"X�%���w�ND�,KΝ��"X�%��u�ݧ"X�%�����蹙4\�n]���7OD�*��a��A��}��wËlJ�%˟�t�{z6x��m<�bX�'{���r%�bX�t�xm9ı,O;���9ı,O��}�ND�,K�����.Hh���ə��"X�%��N��ӑ,K���nӑ,K���ٴ�Kı>���i��%�by�[���)�2�fkZ�u�iȖ%�by�w�iȖ%�b}����r%�!H �����H1��B@$�HD�"��������]��EI����ӑ,K������B����v�<����]U��O9=�,K���ٴ�Kı>����r%�bX�t�xm9ı�뽽��rS�����������;&Y��Kı>����KİO;��ND�,K�뽻ND�,K߾�fӑ,Kľ{~:�MjB��LK�l��\vb��V˸��#���W���F�Zʍk�mH%ag�|�5�MS��w�ӑ,K����nӑ,K���ٰ� �D_"dK��{�����%9)�������晋����Ȗ%�by�w�i�bX�'�}�ͧ"X�%���w�ӑ,K����Kı>ϯ���L��]ְ˭fӑ,K���ٴ�Kı>����r%�(%��{;�iȖ%�by�w�iȖ%�b_�os��欺m�usZ�ND�,�>����r%�bX�w��6��bX�'��{v��bXC�#!"�!�c�A�@��j'�s}�ND�,K�����\!�ۗ32捧"X�%��{;�iȖ%�b����{v��bX�'�}�ͧ"X�%���w�ӑ,K���� �z�M�%����PZRE�i����p��cns�i��ڼeن�[�;�v���OhL���V�;���%9)����oy9ı,O~�}�ND�,K����"dK������ӑ,K�����42���q��Oo!y�^O���6���" �"X�����"X�%������"X�%��w�ͧ"~$�$��&9)�����6�42Gff�6��bX�'~��iȖ%�by����r%�bX�g{��r%�bX�&|g+�)�r�����-'mYj�lN浭ND�, ��w�ӑ,K��;��ӑ,K���ٴ�K��$������Kı>>��_��������rS����������Kİ�������%�bX����6��bX�'����"X�%���@`�"D��$��
� b� ���6�$���ɴ�m�6�x{k����u˰�� �����C�6��֢�&��]aVDu�b�q�0)a	�,`ٌdЍ�
��]GVR�K����a^{l�K�bs��O��X}S��c�[c��m[�T���;�fwW)�Sَ��ϛ!�ɻ��١�i�0�,���J6D�9���n�v2m��7K�1r�
�[uuK%33Z��~EJ�*h��G峓�KJ���L:�L[LfZ&�4b�tu�"�F��s�t�깘�ii���sY��Kı?{��ӑ,K����iȖ%�by����r%�bX�g{��r%�bX����V��K��2��6��bX�'�}�NC��W"dK�ߧ�ND�,K����m9ı,O~�}�NA �,K�����\!�ۗ32捧"X�%��{;�iȖ%�by��siȖ%�b{����r%�bX�}�xm9ı,O;�{�{a2@���Y�O�%9)$�)��{�siȖ%�b{����r%�bX�}�xm9İ? �DS"{�����JrS����?����n����'Å�bX����6��bX�'~��6��bX�'����"X�%����ͧ'!y�^N��g����v��i�Ϸ��Π�6���;v�X͚��-�2��D���=�{ͬ5��2���rS������=��Kı<�gxm9ı,N��l? 0E�&D�,O����ND���'�����7T��)G
��|9(�%��{;�i�h@ ��D6(m�,K}��v��bX�'�}�ͧ"X�%���w�ӐE�,K�߷r�c����w���NJrS�ﯞާ"X�%���o�iȖ?�!�2'~��ND�,K�ߦ�M�"X�%����.���pl��|9)�I9$�=���m9ı,N��xm9ı,O;پͧ"X� ���u�ݧ"X������(�aKsr�9=��K�����"X�%��#���?M��,K���~�v��bX�'�}����rS�����y<�ԩ���x�s8q� NV4�u!�*E.�LR3vI�>�7�ı�c =���Mzh�t��6��bX�'~�{v��bX�'�}�ͧ"X�%�߻�ND�,Jr}��ݧ�'
ګ.N�|9)�N'~�{v���bX�'�}�ͧ"X�%�߻�ND�,KΟw�ӐB����}o�?Ta�5W �<��%�bX�{��6��bX�'~�xm9�^ń! $�	$F�I�-�� �(� �H"HȬ" �HE�AN*$ND���p�r%�bX�����iȖ%�b{�w�Md�S3SY���M�"X�*��߻�ND�,KΟw�ӑ,K����nӑ,K��߷ٴ�Kı;�zsP��j�\2h��֍�"X�%��O��iȖ%�`���}۴�Kı>���m9ı,N��xm9ı,O���>��mD��mlš��s�Bv�\�2�iۺ9�<�v�5�ĽOL8�ы��a�ND�,K���ݧ"X�%���o�iȖ%�bw߻�iȖ%�by����r%�bX���d����L�I���5���Kı>���m9�)Dș������Kı=�w��"X�%��u�ݧ"X�%�~��p˜VR�L�y>��%9=��~ND�,KΟw�ӑ,!ș�����9ı,N����ND�,K��/gf\!�ۗ3&f��"X��X�t��6��bX�'}�{v��bX�'���ͧ"X�~a"��M('�w"w��ӑ,ay���~5��3yDc��'���,K�뽻ND�,K�)P;�y�m<�bX�'����"X�%��O��iȖ%�bw��,ֳSVc�:�<�z=���;8��ܶ�p�xb��F;V*J]CfՕZj����^B���w�6��bX�'~��6��bX�'�;� �Kı;�۴�Kħ'�=ﭬ4�F[��;���%8X�����r#bX�'�;�ND�,K���ݧ"X�%���w�ӑ?I9�y1�NO�?��č��f�Y��Kı=�~��iȖ%�bw=����K�,O���6��bX�'}�xm9ı,OO~ٙzhɬnhְ��Fӑ,K?2'�w��iȖ%�bw���iȖ%�bw���ӑ,K @�<����r%�bX�g��m�r椹��u��r%�bX�}�xm9ı,N����r%�bX�t�xm9ı,N��w6��bX�'�d�s�j� ��w��Z�Kz��eh[V�4F�!0%�Ғ�[,)aIB���eIjK�%� �Ba+
��J�-��st�+q��m�HFgϥg��8B���I!�9k,6�B2@�FB@D�2@�BL�٫H��K���Z��s7�-Ќ��(J�3AZK"Ô�Y�6Q!HRR��L𕨄�7B �~o{%�3Z�hp)xr��90�$���&�U���l!�Wd&3��G�a,�!K!�r�}4�<��9iaI����UeWUUmU*�UUUU**��5��n<��շ*�6��O�(��,t���Ľp��qk� �Vw�k��U��hE9�Lf]P6��v𝹮���L�іx�H�ȒaL�t����iَ��B������[K�Kœ\��w#� V
���Z�-ЌL�)��tv��.h0��Ѳ偺�\�]�,��,����;q���R8��,���<���YN���룚�����9�8��/�vܐ�C��ېݰ ��^='�=��8n�Z�{*��� &�K ;Y�Uqr��:Q;I(.5e.�����&�4c��m:�hm�-5ue�wJ���^�U�F=v4�N�*rGL�v����s]� �2k��㘖��q�N^��=�*q�9�����:�lqXr4f,��1�(B�k�I��^�'el������A��93۞���Ӝ;�\����[]	63O'ev$<���r5Uvd.'ۮְy뒝Ŝ5���b,�%ڂFh.��/V����WO�#�-��H�@лL ��Lݳ;�=�7U���p�` #��hx`�pv�����+ �@1�[5�)Q殣%�H3�D�Ge�ӄ43*�E���U['��Z��铍��I��m���Y/2]��[���w�ԫY�x��e['G�H鍠4�k��_k�W9����
�2̬	m��붆+	l`���
�7�˩ڄ4I��u���h��;N�sڡ���n��5�7�����k$,m���T&�.����b�5�ڡkcAc�*�nA�eX��m0M��s-�(Z<����q� 98��BV�m��,��î���^{�x��G+�=�t<�^om��)��ܝn���.9�CՒT6�ѳD�����lu�^@��x���֮x��N+ca�3���3Uqbݹ紪nrZb�!�K,U��V�Ҵl<��]',��x�me+�@a�9-��-D)�D�i+'`D��K�����:3"Y�[�M�#��G�I%�F��U�4_��(	�B"'��6 |(l4� �@0�@ڞ��7�z�%CL�t5�T7.�p.6�����y�&rJ�]�&6l!@/(�x���c�ա�D�k�^1^�K�i�7M�[*��61�yKv��m��6��2�cPe�c��c�kJ�$��9���<$����	)�wƌe����:$�% ��9�%�3J,�R!K��U��F�l��.�&13^�/5�'gp�3n���Y��d�a)5�ҫ���[�-�f�u�/X�\���T�ci(i�P�6�3%F� Z+����I�}f|Va.u�Ѡͧ"X�%��~��"X�%��N��ӑ,K��{����|��,K���ND�,K�v���2�Y�Z�34m9ı,O:w�6��bX�'}�{v��bX�'�}�ND�,K�}�ND�"dK��W�h��Z�e��'Ò���'�����Kı>����r%�bX�����r%�bX�t�xm9ı,O>���2
�
�kV����NJNs�Q>����r%�bX�����r%�bX�t�xm9İ,N����9ħ%9>��}�h�ksvgy>��,N��xm9ı,;���w��n�ٕ��Z���S-Ӵ�[���,�uv���Ћ[���n�hV:�0�}��LfVU�Z�+�!��ۮ��>��'�E�{ve`d��=^�WjS��ۦ�53F�{�}w�m&����y�b#�e`}��Xd&V��Ww��`��[k ����&�W9\K�|{��=����}�K|�Mtuq˓ft	��weL�z�XW9�-������w��B2����?y<��������t��n�`t�tF�t�­A�^�[YD�`�nոA�����b�EU�@̓�5�@�r���}��ٕ�M�ܮ~�W+������o���ֹ�
��[�>���g�'9i�� �����'�E��ʪH��������4յv� �G�weL�/��91�l �Z�@���ʪ�R�go �ɕ�v���cV�ݠC���0>�W){~��X�|�{fV7\0�k��O�2�:i�U��'�E�}U\���k�}#��;�S+ ��|n�jf[����E�[WF`�r��U=t\��7��(-��I�[+�m�����l��&��Jp��U]A���, ��	}�;�X��j�`u�>�*���������,�ٕ��>QR��5Ќ���e:���Ӡy�y����9ķg�X�?������e��c���\��_�,v}��M���駱֙$	R�Rւ+��!JA0��*`350��B0�����l��EdBnCWHD��Ӏ�%t�X�A�3�/��i
7��o�'�����bN�+e����I��M��G/Ix��;�Mڧ��
�7m!��4pu�NΉ�ud�\Z��'^og99+����i�Gg\π{珦飆��ޓ+ �I+*ƭGkY���|�>���KOo�}�wﲰ	��mn��R���L)�`zK�7���\�)/��Q�`�l����v���i��7�� ���k�ܪ�)}{�׀!B_}N۫��j�0	��zY���%�'�}���|}HB$�����-���[�l.�-�ؘ9R�iP�p;�9x��<z�eeNy�<{Llt�E�8�b�b��8�[���q��'l7A�*�g5f��)E[Nlr���ZC� KKF��Q��xq[u-C�U�j^z����ua�)���n9Nq��gqms).#���f���\��{I[�s��r�ٗ����=[3 i��f50�퐓��9�'9����>
L��WbM�Q����,S�7c��ye��ƍ��#�n���35��6�B�5�U>��y��_l�}?W9\���r�����J�gʮ��P�4��w�E헀o��=���/?W9�~�Us�d��t_�-�E��hw�}??�=�w�K�Șױ`��VQB��H.�����J{r��}x��X�8`�%eX;)�T�uvճ ��e�W9\��}}o�� �� �ԫ-�V�����1��)qu�TrAtt5��9}���/=\��+2uBS���t�Յ���^����}\��Po�O� �%ڿ��*탷f]k7$�ϵ�؉H�- Kg�{���͗�E헟�ʯ�\��W�~W��۫��j�0����=/T�/l�ގZ�nwt0N�wi�ꪮ-����-�^�G{\0T�U]�	�m�0����\��|���飆 v$B�q��[6���S�H�o!.W�uAi��v
h���.�Y��5c�Wt�w�^�=���W9Π�l��o����+�V��6�{\3�W*�#~��X�s�{�"Ϲ���vm~�����V�$��f?|~��'�b��+��9ʠ`�H�-$U�H��	2�ĴB��4��ڪ�}�o�rN��vnI��e��������s���}��߷�ށ7\0?UW8�~��XR]��n�˧M�m`�Ȱ��W�g�@�����;7zym���.��p��l�҆��Xqʉ�q6�ħ�����|��pb�f�{;��QՎ�E��]H�0zT��:������߷�ށ���oIv���M�������v\� ��E�n�}�RF��E`}e�ӱ����\� ��ސ��;#,E���t�i6�>�q{_�,H�0zC+ �W## ��HE	�
3&N�v8]*�V��6�w\0�_��'�ǫ�o���`�Ȱ�[l(K��$c1���ˁ��^#G�X�J�rK�.�d�\=ON���.�`�V�r,���Π�?�H����𲝵M��u�v\� �E�n��Heg�s��\�>_}ww�7e��|m�m�e����p�=����X]Ҡ�5iՎ�E��XqI3� ���+ ���W9�^��� �E᧥�6�6�S�}��g@������3���6_�� ���UJ+��PUq�1�, ��?J�`�:wnt�m���jj���
ƕT��	!��2v�M�@��"t�Q�v�9�[�/�		�F�tYɍ\X�V�K�v��4 1U,pr�h���&1�chMlkL�y\Z6����^�N���6�ʶh��<ϴg��u��H0�)��N늇ή9K�)�.�7��7��k�iݠ�r���Nq�=�5(iE#/n�X�a��t`��&h�Z�k��C��l��?;���N���7��݄ܛ�ͷp�͝5a�U��
-���ZK��.AQ+]�E�w�"�&��s�7~���=視}�kL�45[�>}�y{��I�Q�� ���+ ��~�H���t�h��uwI�۶���!��v\� �E�v�J�B��n�$��v�ސ��;.E�w�"����$όH��_S�e[iSi�`�"�;�`u� ��2��Jww)S����7hl�� {6�`��1�Jn%�E��i��mG�ۺ]��Y�4x��o�>���z��>�ŕ�O\� +�V�[uc���]kWrO��_M���T<t�)�Y�>���X}r,���$}-A|R��Rwv�ݖـ}>��	�a��z_�,��ꗥ]�G*J�i۬z�Xdp�&���9���~�~�~e�K�&�.�ai��vG�(����rI����rO�Ͼ��uSܝ���rtK��7�p69�ۃ�kq+5B(^f���$�0pL�SI��4�I�f���O��� �)��O\��*�Π߾�ﾬ.��T��+� �)���>���o�?�n�`���(|VU��7I&� ���v��ҟ+UVRW����wI����yd}���Ⱥ�����j�2�o�������H�
����֡5_��/ۃb�y%��O9�]@��	�9�JJBa�ĉNJ���6n���]�W��!�Býz�o\���c2=׬���ɭ���&l�J�JD���$��BF"M �B�BI*KXY ��HH�J¶�a,��hj�\��(Ci��DuM�NL�Y����2���_u�9��K�f�	��9��.�:�%9GJ9e�%�1!��O	E4� n�<��e���1��.K�-� �o�浚#t{#%�dְ�����)#/5��bs�S�nO�[��.dH`ș�P�(e�k5ulf�o��6F���L��XA�30���|��''-Ԟs�n�t7!r���7�$����0��fk4s^)��B�B��$��@���o�	�X�p@�����K	$�H� ���d"�"�Ba�������"b'��"��O���	�� �	�>��jy�׳rNx}���=���cŦ�G�͖�?�9�o}���t�}�I��O\� 7�l�C廢���� ���߫�]���7c�@�}��<�t�����\Wv�f]�,���Xj�'b��d�L�nf��76af��n�Ym�~����'�E�n��A���m}p����Hۢ�u�O^ş�s��'�� �c��=*L��I�]#��Wn݅��'�� ��Ҥ��'�b�=���4Uպ��t7m�R�f|`�}�V={Wh�*��0B)�dDST09��H}�_/��g{����"F�L�i&V={�0	�p�?s��}����8���4I�H�ֵ�Z!A
69��0	o4�C7�t�T#�B���.��ln����_ߖ�0	�p�&�e`��]F��J��۫���3䏶?��}�V�{~�*�	�O�t6�Ym[f$�I���K�X�?�m�)6�ӷb��0?r�T��������,v8`~_I��\)Q�j�BB�­��'�E�o��7\0Jٕ�g���\�Q��UY�V BR �?1�FbbAhDF��mշ>Ӗړk��nQ�U4��-�#"XK-V0�:�@�"�Y�Z4CKĄ	������ERcl]4t,�P�%P�u�Y��WFs�]FzS�U�@.M�mȈ�����Xf��x��Х%�`.	�O�Ľ.U��#m��)�LZkh�5���k�����/
�O=o��� :��Rg�n=6��r��a�\�Iv~wt�wt�6�a��{>�따����8�0�[�l�\�cX�s�4l7�/F��E��pj�����M�Ҷe~��P}��� ���CuiI��;��l�&��[2�ˑ`��U$z��VI�ST�;�ـo�>��;.E���U%7��I����7�Ĭ&̢�9��/�_}�o�� ��Ҷe`�Ԯ�n髱�۲�X�8`��zV�`��/@��߼�l�CfD0l�a��cX�q�9N����P���L�P��ٳ�)t�Ym[f���k��r/ܪ�9�~��_*M�)�b����'���?Db0�+��FB�@(`W7�����:O_�XϾ��7u� �/JTF�H�v���X�L�>���� ������'e]7C�:v&���R����$�)��R���ށ������4q�t[�?~��`��s��V|t}|�z�X]�V�fc<pM��] �Y����4eV[�q@�8�j�A���)
�SL�&�c4fK���{Ҝ0ˑ`�ȿu��`���N�vm�m5M�eȰz�X�`����.%u�n�t��j�֮����ܓ�}��p!�{Ҝ0Kذ�V�WC���[M���)&|`�S��;.E����$όKEE��l)6˲�0�Nܪ�=����$�� ��wJv�t�(�����F訆:�CZl�@�4��A\¤3���
w����Km.Q�3�{���n���d�����St;c�bm`��U$I�ﾧ�v\�?UUq#����vU��wN��0	#��;%8a������X��`�����ҰN�c�`��0ˑ`��ڪ���QW\

(f� KJ��@ $))+���A�� �Ͻ�f�y�I�Md�aM�Si�l�;.E�~�$���$�� ��~�9\�T����ƭ�X�#���"������aA�a��������#�v�`L6����J�Ս��]H�0�p�;%8~�u���X��W��v6"˦�0�p�;%8`�"�7u�;UI���tYwIc�S�ݽ����0�QTP�nƩ� ����`��0��>*n�m�Bm`��n�݃��r,9��8���j�W8�G*�+
Z��k(��a�ón9]�=��$v�'��K����]8�ن�e���Ƿ��њ��,өC��̲��$��zFuÚ���;��wA8΄�D�On���v�����2��8x:�#��Q��'����S�xݽli�.KY�d٪���"5ƶnv��I��I�S�1l�)��8���`�Ύ������%%Y� ���+Љc�\k^�ςI��-qB�`�]�:W2�q�P��>'e*NҺj��k�I0M0ˑ`�Ȱ�ɁWc�t'b��0M0ˑ`�Ȱ�p�=�pt˧�ؘ���eȰz�X�`����+�m�.�1�[k�s���5���$�� ��p�;.E�j4�]��e�[M��n��Z�v\� �\� ���Lo�	I�mcE��;[�16ֱJ��%4�ۧn�t�Z˖"�,e#U62��\0ˑ`�`��zZ�J��ZLֲ�Z�ܓ�g�]������9�^b�7u� �k��� �ձS�6��Ȱ�p���+�}�0}|��w8������@۶��p�&��v\� �\� �l���+�;�ـM6e`�"�7�"�7u� ;�R�e�J�;Ǘ��3� ���D�'���Y��\H�ᥢՋm�����۬��X��X�`M�X��+���J��X�-��j���n�4ٕ�v\� �i�Wc`�.�i��7u� �}��ʃ�=b,4��&	Ձ��W Bo����>��ٹ'��B�i�R5Sc)����%���~N���﷠j�^�����e>	PۺBn�ˑ`���n���� w�~����e*� u[M�F/5(����ݴc�K49�[�
��
	�8nK&��Ix�`*8`�"�?���bv4a.����=�~�,�����X�%��\�$z��`+C��'e����eȰRK�7u� �f1۫�M����eȰRK�7u� � p9E��BB!!$�"�D�IKE	c �d�"@!%+Y"I1���7ߏ���'���}sYqUӦ6�m`�K�7u� ���}��O-���v��2�.Vjhͷx�Zx�渞�rcD��D�@���%e�d�taJWa�e�e�t	#��=*8`�"�7c��h�*��E4�.�l�=*8`�"�6Gw\0Qm���|��h�l�;.E�n�w\0J�dQ
v5lT�M�ܥ'��I��Q� ���ڤ�v��ݵ�n��Q� ��r,��*ݢ���-.W!!�I,�A�@]�޺54��9x[A�ܻ�\#�	�!	)JJ0���̸�>s>�3�!���x>��h9����cf�%�������D!�-%	w����VYÇ�ќvI�����6lK�.+�k)����)Rk��-���Z̒$��� fd��\z�z�=þz_ɦ	t�L|�]Ms	���59���|�T�����5ag����߾&�&p�2c�'�"h�4��HR�a d��-%��v|S$a3��4Ѿ2V9dJB0X��a۶f�i�7�xK9;�����~i�� @�-��l�;i(b\~�S��Є'*D��s[�f�\�q�0���Z��fFa�r��Sa0�iJ7X����}���5��<��7.2�ğ]��5���VE��Y��^H�p����k�u���� h�������\�_�JXBcS	���^S7�9���f����g�Mxܛ%�ֈ:�ㄯ�Mow�p���\��4��3���y���5	|�2�����߉�P����Hb�		 �<�"���"�P�5�~R���8B�\$ �����@������X@a6�b��u��K�ƙ�B�L��f��7L���p��|�>����V|���!/9)�����UUb�����*�UUU**�2�*��8���=�2��2`C�n�iڌqֻ=B:ZD�s�K��Վ��04LQECJ�� f�$����,ZiL�W
XM:i`VRTj�͗�����M��X�m1����cn;]r���N^<\MX+]�c;�2\��s�f�<��2R���3���<ڭѸK��fs�s�y�E�%�
E�n����m>���Ǳ�\[��Ę��ā.@bťY0�K��Ґ[l�������냬mt�T%U���h(Zg;B�h�����ȵQ,H��xM�O� Yزv��	�)��C��e�D�٪.�Jr!�|n��{Z��l���)0�`��t9(�8Qr�^�C���6v�6��<�6��.1���V9����vā��w)��^�[�YJ�;R�s�F�� �u%&d�A��ٱ�J3�F6������70H���2�K��N	�u��iDf��cS�8e1�v�t{��&�9)�lʏ���`��H�6]Qn��h0�#k�]4!�$��C��G'�u̶���Rcf���g.�p�@=x�n�3�����ñ�]6t��Df�Ә�v�LÚ.��i|D^�,��Ez:�Mh����P�"[!s+����ZCG.�7.cbA�"ݧ:�g �@tʲ�t�0�u(�]Ev�|l/��r'�����:�^�P�k>]�CJ9݃F�h�13	�.���8 ܤ]�N&���K.Q�9���t��m�������ė�F���n����H��v�Nw�5��gyh�m�wY�
@�U�n��M;r`5�=p��Fr�ף�ۘk�	�K��t�K�.!�Ue�7	CBW���0��1ĺ%�x		�W
�VYr-�4wb�Ս�'�Ѣ��
3n�o۠���X')W��H�Zh�bb6JV�er@�n�,Mh`�H���l��b�ڡU!W�)IrGcT`�My��qX�:��ۍ��
��=G3\�X���u$�)�"m<E�G� �D∞���.�A~U��Q�%B��iUX�x
x�������Ӱ��	��K��i���N���ѷ"�F�7���Pf�͠ p%�-BVe,��gL��8��$C-R�!���]T7^�m׀V�� n9��&ZJ5��ď��鵍�+��2Z��:�n�Qs��br
�8�D�I�������ru�ڔ�4���H���p�k1m��A�|u;�u��R�9�8;Pj�(��v3c����]���W�:t'wr�Ov"�3f�+iaM1.�P��5��i+]q* ��(�䋏QT�(^�:I��� ��p�;.E�n܋�NN|��>��<��s5qa���;.E�n�w\0J���+��ڵWN��-��n�w\0J�eȰG�"VƀN��L��w\0J�eȰ��n� �6���E�l�=*8`r��?�]K��n��9^���;��dvE��MgZE��v�}�����0'6�%�g.⋦�6��H�
�K��}���ۑ`���:�~����Q�a�չ�L�u��'���]���"�$���Q� ��2��
�ںhv����G��X�Ȱ�Z��N�����v�i0ˑ`�"�7u� ��V�ӫ�;�`�"�7nE�n��vw�O-�N��7f�nv�"�+��h2����3��& �.�m��q<L˛���ŻV���-��n܋ ��Ҥ��������� ��_����V]�[f���l��;.E�o���h�Q@�n���0Jٕ�v^˹����Qq�B��A�}�nn��yE�J$��ݴʶ��\�/|�� ����7���-��|`���wWN�V�Wbm`��wu� ��p�;��`G��-��v���^�+�����,4`skto(Jb�;:���ŗ],v� -S�|����|���{��vJ˵N�ht;nݵl�=+\3ꪪ��K�,o�� ��=��ui�IՎ��0��X�8a�q/H�0����&ޤ��Z��ch����w\0J��ܘ�Z�s���'�y���Ժ�%���2�0�`��v�,~��t��߱�M�Gfk��5jד�w<Fܧ��⠟���m�͹�l댥�0r��B�l�B�� �ݗ�o�����-�Q'l*Ҷ+T���:�e���wu� �^ş��\H���E��m]���&� ����;��M�����xv5����j��M�w\0	��^ջ/�W9�7���>���h�h�+U�:�����[���p�;��mh]m�V�EWK�l��2�M�����4`�as�V�\n��l�[��� sC:LͨVe���R��ml�*l�N0]�k����&�f�m�Ĵc�M,X�[��k5k�&�Sm֎��'���x�i�L�3;�f���� l�t�W���x5�-�i^8��n�a�b+,&�v���`����,�ڍg;��k��j���4�%c�f�c��˲��iwUuɵ���Y ��)���1���&:�r+s[��;����'׀o�E�wu� �ke�oRWN��,mZn��Ȱ�`ml��v^~H�ؾ�t�@[���i��=#��&��xV�W��v��6����B�l�&��xV�W�����[r��*-[T�n���x����`,�x��9ʪ�B����M;��%�sN�e�K.�w3��+6^��Lph��`z!��κ܍r�:�� ��绠|�p�$�����xv5
I�*n�,U���χ{ǀs��9�rr#(�	��G"K>���j�^�l��"�+l���c`�X��^�$�T�x��X����պe�Hv:-7xT��Se���`Z�x��
����n�Sj�w�j�/ ݽ� �f��:����?O�߼�9����i3��z:x��[Xx˖魡��� jw\R��Xzc�+�v�����6^�$�T�x��m)���Vـl�e��"�5M��n��-�j�n����1��;.E�j�/�\�V�  D�1�R
H;R$X�`�b��%E'�����{�Ixd�J�Ӷ�N���5M��n��͗�v\� �ơIժn��v��w\0�{�r,T�x]�Di�][�-�0�[�K�'$�lc��vUm� L����c��b�f�կ.�(Ut[�lf��b�;.E�l�w\0��.��c-:C��[k �v�6\��{j�`w���j��۴���X�p�7u� ��ذˑ`�h��|-��۶��{�W�`�"��sJ�o9Wz�,v�Q����-6��W�`�"�7�"�7ob�$�;�RG����^�}�,ďDZs��:��Am犴�cj���`\�ԙN��r,}r,v�/��]A�T���뻶�iS���}r,v�,�G�Ix}�,����un��m`��`�8`RK�=�`�3�v��Ut��v��=4p�:���{�"�7u� �V]�M�-�:��6`RK�=�`��zh��>s�~����^�\\9�^��u[��)���Kp����wof�dU�ѩ�+܇��^۝v=�g����rP,��S��©�#��n�vW�e��$�0(@�NZ�l�tXa�8�4�Җ�ie��mɱ�T.5�o9�'l�!L�M���KFl:��v`�)����f�\�\dceMq��t>;v�5�s�vYx4���L�*!sY���]S��|�}�٭��T6��UΊ���]a���qv�|��x9p�<4d�v'ej6�)�7o��������Py}�׀j� ����.��m�w\0M0�%��Ȱ�EW,SNݖ�� ��� �^Wݿ�X��`Qluav�I+n�e��T��z�X�`�8`����Z`��*v�w�{�"�7u� ��� ��{���zz�a,R��!�����9w���&�����.��1������G���V�v�����eȰz�XvL��v�Uui��� ���6*m mt+�,�ϳ_]�>�$X�g��W7g�;�N��n��hcf���\� ���G�{B�Z�ն��m���-��� �?��Z� ��@Pv]ZO�ݱ6��p�=5��ˑ`�����O}���/h:6��V9�8��rs�`^u뎻T+� q��4�
�,�3.�14�m�~�|��%��Ȱ�p�<���uv�I+n�e���$�ގ�`��Xd��D-0N�!�M��Gw\0U��Q�4�|���D��,!�B"dހ���	Iq��8��hh������a�M(8B0�(��@�Zl�򰛕����1�q��l�RK� NJW�Y�DL)D7�P�Q�Rda	�)��1�#6�tJK�p�eLd�#F	$.K��{&�����D.���1N0jc}Ӣ[<ւ��@!���'���;7�a���`K��	,��b1�c����Sm,a[q��K�P�y7%%"NS�j�9��B��&O!���{��M�}�e�-˃�e]��y�aKHL-�$�.���@�l����?!���4��!�EqO�<>X�z� .)� �E��M�k=��x�e��ܵuwM6��i� ��n���$���vL�5IUՉ��v�m�XT��	��n��/j��CMؚM��AV�; �³RةZ�{&+�ݸ�r8պd�e�mΓ�&���<����'�����NrO�=�y����y=f���fp�X�pϹUUIG�}.|�ˑ`n���E��]�� ��m�XeȰ	��n�8H���7bVف�Rߜ�`���`�ၜ��:�iB�P#6�Ą�(�,C�Bm�;{�f�_m�)񚔪��k ��r�Jo�>�$�Ȱ�!jR���j�����h:,3��1�8�7G�@q������q��]�hN�Rv[k 7dx�`�"�;.E�n���WWt�n��&�w\3�s���_�,�_�, ݑ��URZ}��{)����V����o@�s��9ĉ>��G�{�0�t��i	�.��;.E��<w\0K�`^�Duh,��un�������Ȱˑ`���#B�)a$
@�b���#$ �I�#̣��g�P����	[p���M+v�+6�"�4�R�,̀r���{:�燧Y�D�;K���&<g��EF�����2r2=�v�.��.���9Ϩ�2���R������LkSJB*]Q)�!���a.�5R�ZY�����b��Wkc6-���H |�׿}�G�n���vA�R %�[�Gv�5%���اsI�8�Y��̊�b�Ž�?}|G�
=-���[&Ȑ�ZL�S���;�X�>�|��c���ۈ	�r�@���Z|��o�M�� ���r, ݑ���!1!�Mؕ�`�"�;.E��<w\0(�*]Ҥ�ۤݻk � n���p�=/b�;%�K����������r���߾x��`��`�"�7�j⻱S�l�@����p�=/b�;.E�6< �ԥhl)sf	�A�ڐ3AX��h�GI٧�ۈBnL�cv����M���`���?y�yzeȰf��Ur��$�� �>�v�������wzy윗��9�q��W����7��l�� ���[���-��[���fǀn�%�XeȰ�n�A�tZ|�ݷ��9ʮr��>0	�ϖ�$� ٱ���wI*nĭ� ٮT��fǀn�ݠ.A�Yv[*�+���W��`Sp^Ya���N���n�o::C;8�ҫ��$]��[�l�:���6<w\>�	�����_Ym	:e'v�� ٱ�ܪ��8�$�?����y�N@���I�Ԥs��nE|�$�p��Q ��9T�@�!'Ɉh(��O��^�|���bVi�������r����<��������f[�Wt���m�� �^�l�w\0�~|:�O'��﹪��;aKf��\­�J3U��D^ˬm�j��X�� �vZ�T�l�M�M�@������l��Ix�ۡ(��E��]������*��'��`���`��Ϫ��i皐�����e���{｝��Ix�`�U	t7Ii�V�[������E��^��6��# G�d��By	*""�1Q%h�F�Ԅ�Xt�4�s=�����ߥ��6\��j�^���2�ˑ`����eqX�i�F8��s-�$.�9�-�Om;N����������$�:5�zn�kk ���L���X�%�vF���);�:� �&V�r,eȰ�p�7�0j�:��m��lM��r,eȰ���s�I�>���ڒ��$R�@7cm`.E�n��L��\�^����"�t/�4]�v��X�`s��T�}���w�rO~�~��t脈�@�b����P�	��w�ٌnR�s��98��;SH��vwG��V�b{=P�n�=k��v�	9��R��5*vۧ]�]-Z�e�-�Eb�]��LXj�h�v0����G�)ϱ�l�u�*�}źٗ+���kT���|���������;��d�a�F^:�i���M�w8�1=���Pl�1�[V���/..oSF)�5լz[��h��%�w~t��R���.�gh�v�� ��B[�R�TK ��OG{)b�/)q�����l���6߿���XeȰSe���u��`|�|/��H�M�۵n�ˑg��&��,H�0M�Xd�2�m$��We���Ȱ�p�=6e`�"�7�j�'��n�۶��p�=6e`�"�5zK��Z)�)5i:� �ٕ�v\� �\� ����Ӯv`��m��&B��a��KY�epU�l��L`%�HX�R���/*�3�3Wn�ˑ`�%���`�2�/jJ:t�Un�wcm`�%��S��S�U2]ά�fV�r,���$E%����tZ|�I��$���=6e`�"�5M��nڣDZ�E� �v�X�p�;.E�o�E��W*��|�_%_�m�����l�;.E�o�E�n�ŀzk��W9����]u��^�h�͵���vi�#���j�f����=���+n���&2Sd����߷��{����D�����
v�`;v��z0;�z`\� �\� ;��vS�)ةЭ��\��s����+��T��5~�ެ}�������n�I�-��v\� �\� ����\�[�,VėΝ!*�]��X��XܮTٟ~���;/b�6�V�X
�c&6�Me��ж��r���7�7a��g2�"�����:��S!��!�J��~����r,��,v�X�6+n�b��j�0K�`��`�"�?}��w�'9-?_m��{�.Y�*�}s�n܋ �k��r,�A1�i+mp�-��n܋ �k�����rt �8�T.{�o�`H|�JO�;wWm!۶���`�"�;/b�5l���E�պ��6���K�;��!��!vxd�:���5���
�xn���e�v��-����巪l�V�r���c��7g�5m�t��;h�k �/ �$�}�ˑ`��Kt�Ī�𻶛�T����`#��6^��t([�Nʵv�ۼ}���uM��j�^���M�ب.���dp�:���6\� �k���G
(�P��&� �0�!y
�b��(B�c#�D�I�V1R5ӱc�E
x������FH� �M8�m�f�P�`DD��� �*J�o21&�]f�o	�����RBP5���D"�@�+	$$H�<��r%�si�)a���ʄH1��#$"J�"@	l6��l�C~７C[�q9�@�iKFK�!%VP%-����f�G�}׋Ĭ:�o�̅���s�r��3s�kf��9e�I�")
E�9���dQ�*ʮv�}��B�
k���m9�#0�>F�74dU�I��"45Mj�f`K�O%id �����3|RGfIVa��p!�В�BV%	XRBB�Ō�O"�A�8H�j1 ��
J��vۯ5UUUU�TUUUUR�5UT�O�\���q�����S�L;���<mcD�l
	y����(f������JY�W^ df-l4q���c�U��<m�8aw;	�+ǚ���˗F�h3F�]�H�1B,o�b�Ƽf����5�l*X��M���E&c��ԕ,QqOL'��E˲���Dk��v!K��
�@�=�,E�G�T�4
,YS��轎�L�`�54-��n[���X��#g���XZ�:K]�Z�Ęd�J�vs��
([���]�F�©�K��t�!p<�6�7�h�#�/��l;K*ƽSQ��^-��QR	h�=����-1M�;�hvf�e�l���˴	���!���ź���ܵ�l�m�c[0�qJ�SB��!l�6�U$Mc)�]&��v�L4�MsR@�J��=Piٚ�#'To.t;q� ��06	^4Y^Q�]j��%n���VLְ�u[t�̅Ľ��[�mav$�Nb�����aۋ۱�*ck��`Z�r��>˹L���u�h�e'8qX��;\��ۈ7mM����rnȱa�6�Fk@�i���Spь���n�S�+�����3���u��^A7F�9wO��쪪A�lYs�Fx���Wd�;+��6�1�a�u�3��/:1�9ϓ���eݮ�r��v�����SYfc�6�)��,�tΘ��]chy��3�eM6�u��ذ�\�nl+�8n�/H�&��G�lN5�t���=�#�����Q
3vl��4�j�f�^�mn\=uX1���J8܏����9m=fx��r>�q���]k�ٟ�~'���˦���%�ٮB�s���B4�1�q��$ͬ�:K+T�Ă	��&&ͱ�!"�f:��I�@��f�0�t�H�U.G����اg�qKײ�)���m1ua�ޖ�Ձ�v"[�.�b�v�C<d`!��s1�����V-[����کz,���ǎ��rۋ��Q��� #:Ђ>��)�h!�+�1C�S�V(z��/�Рlb�*y�p��~˼ө)�M.g4��Z��9��m�7Z�±-֮�D�g�V��tgWe�:��^B�*�v"�}�J�e��1������V�u<RP��h]�D�!ζe�]����tC՚z�=m�Ts��M xC��t<��x�Te8Ɍ��k��\i�O��΁�۬�vtN�=����׷KE��B������n/)����4�F�#vm��ͱ���='v��	|�W�r�R��60ܯ�\�)�C�<�q�h��
w<;ҭt8�l��t���P����.E�o�b�6I��vh&�K-������7xˑ`�ذ�e`Se��r�$>k�TS�uv�M�ϯ �&V�6^�Ixݖ��o�tSB�իw�lٕ�uI/ �6^�v^�ٍ+v]�ն�C�XT����`�e�5� ի`Sam�wv��n����5q:�	鋦(�
��0��6�+u�Gg�n�!*�|.�� ��/ ջ/ ���Ix�m�Wi�ջ�V�ح��=���o=���P�,��l�+��\�*��s�f��`���7�"�y'-?y�_o�.��	����|}0�%���jݗ�yD�Je�Wm�n�f�$�}0[��>�9/�|�@��[}6ɶ�˶����/ ջ/ ���Ixؒ؝��x�/"��{��W ��ݨ+e"��tՐI���D')�Q@��e̚�~�5�/ ���IW9U�o� z|`��X�f���'9�s��W�}x���jݗ�UU$nϱ��.���ҫhm���}x��XJ��UU*4dX
RD����) ʁb�`�(�+QC���U�a�x��� �����H�𻶛�}r,V��\0�%����j�n�U��+k ջ/ ��ߦ|t/����Ȱ	�Q�iy�n!ZbA�1&ɳf������ϛ���[�1\+LBV�4�M��f�`�"�7�"�5l��yD�Je�Wm�n�f�r,��&��,)�׀zk��4�Kwv��m�}r,V�x��`�"�7�j�m��n��uS��$���yﻠ~��� ��r�K���Uz�n�a�l��N��$����z\� �GV�x�l��UՉ�6**��7װ�p:�9퀽&�<�K��<���V�wv'n�[Cl�=.E�o���d��\0�jJ���O�ݍ��o��}��9�$E>���?���X�m���-ݪ�v˶`�K�=5���r��o��� ����=�QR��t6�t۷x��`�"�7�"�5l��yD�
�1�Wm�n�f�r,}r,V�x��`�ˠ�9|�?Mm̢;�b�!�f��Pr���̀�`k.1�6z�K�u�㓏\�^�{#m�;q+�Iq�-�jlR%�#�)@�sW!p��e�Z�j�Zl���a9�\��z�k�k�qaGTnS�J9"��UF�<t]��AR8W����b��֜(�e�KL� `�U3�%єjZl����:��h]:3�`��i�Bd�S��M 1CZ���$'y'9!�A�c|]eD;%�ú��.��ȝ�\T<���%���pGh9L���{�ձc�Qm��m�m���5l��zk����\���M�v;�۶�-���s�I�ϟ���}U�${~t���S'`�&� ߣ��=�� �\� ��/ ��c�]݉ۥcـ{c����ܮs�[�ό�bJ�+J�|.��f���^��p�$���.Ҷ�m�騠-if$���tZ:?�OOz`��ڮ�&��0��b�I�Z�v�ZLM�)�׀zk��0�p�=�QP��趕t۷x��a\���#cp�7�� ղ^��*��t��hm+u�zG}0��U%���7��V��""���n��������I2�K�`�j�]�*vաݎ�f�d��r���t���`�� ;��9����A8b����jݱ�эn�,:7e^GShL<�*�x!(�e����X�Ȱ���9UΠ�}����b��nv0M��r,v8`�K�=$��:��+���]���Cm`�� ջ/p��PU@��XD�`%FB0h�b1�+�x�Q��B_>���6^ŀj��E(5j��Ui16`�e��e`�"���O�� �e���N�Ң��m��&V�r,v8`�e��r�Wv��e*J�n���su n�;���5On��l�;�Ds�Ș��PbF[��3�|�y���GV��L���DE7J�we����URDR}x���XeȰ�5r�X�[�Bv���V��L���X�p�=�J�����t�w��+��-����<����7c�r|"����A}CH)��2�{ec�[wi];+f�$�v8`�e��� ڄF[�K%��ո�]3��v	Fj�+Yi��*`zĎnk�̃�5�a��E�[~��LV��8`RK�5V�ڴ�*���0[��I2��%��x�w�s�Z~���Vf�EWt�ﲰ�%��� ջ/ �Z(�T�+m�2���$�v8`�e�}�URߧݬ��Б��v�;�M�����x�̬�Ix������e��O�|�	��Q4f`�������Գe4��\�L� )]�X�����;p�`v#����sN+���%��z��-n�X��5����l©)�nl͙�Rј8�hаv�P0��u�F�y^:ݚN,R�mF->��N�m���*fJ��xY�ز��7g�n �v��doi�(K���Wum�Ѝ�u��ʂ�Xś]Q�,�;����'N$��'���>p�R��	lb[p0ɶ�'bh�f!,�X^��p&��Ba�I��T�ա;N�g@����=6e`RK�7�"�=�K�|R��&� �ٕ�uI/ �\� ջ/ ��p�lv�%t�`���$�}r,V��\0/jJ���[��M7x��X��x��`RK�5W��J�Zv�ZLv��v^�T���Ȱ����"����M7�-`8kt��2p]�K�`��@M,�]ޏ�j\��\�A	�30R��U�@��������7ף����>Q(�\�t��N�w�'/�}�� lU(M* G�"�r,޽� �/ ��Б8�%v���w�o�E�n�ŀyM��uI/ ��N�R�n�	�v�v�,�l��Ix��X��)po�
B�	��yM��uI/ �\� ���O-���:�d����l���ZC�/]��{!�&����x���dv%�)��\�J�6Zn��%��`�e�Se�^ԕ�ݪ�V®�M����v^�{�$�U{m#��;J�M;k ջ/ ��!��
*�� g�e�SQ)-�m�Ϗj�z������w{��a�9<LbSI�ޑ� �	�9�X\��`hL��`0�!F25��At�V�3ZR�Ɇela-�M\\}}$�m���Ɛ���>	���M�p(�R�**�=}g��T/��;�gM���y��r�y醵�'��XE%伲���BJ{ᮎ�	�ٳ߈_Il��޽���~h<ׂ��@9��{ȼ9d9�����5�Nj�
���B����2�	�.!�!	�O[�0�︦2o{�� ��!LVŁ-י�TO��d��!.�)�p�t�팖�t�HB��y�0H21)7	0�cF0�5��F��&��"&�854�e��3	0͙L(x����1 �5����|��y<��=`H2>:�!�4L&������8h4a�[�0�P��$	�����2�p�8H\	\!p%ˤD8���W����@ >�m
��t �X�)�RH�!!$��Y	c�E$$!!HHFH���BDXDXD�H$ � I$��C�ņ)�#�j���]g�[� �r,��QW-�t�J��m�x��3� ���� �\���qK���5|��QU4+ӧi��;.E�o�E�jݗ�yM��Mҥ]cI7v�M�]��i�#����ٶ�c�͕�U���sa�a�,�2R�\e���痠jݗ�yM��UW9����`O���e�ա;Nݵ�jݗ�yM��v\� �\�>�7g�I�|���V������"�7�"�7ob�=핉�LJ�b�M�����X��X���rC@ǧĠ�(�!�����@!h �V �X�JfP&I�(@�@� h4�!ڢ%���3rO���s�Y��c
V�l�7�"�7ob�=/b�;#����NNv}��[���a%�3 Jl���˘��bi�&u�����nRV]%̘�v��Z�,n��\�`�ذ��=��|���﷠}��Bor��G6��>�s����z_�,v�,�R�Qr��X�2�Xdp�;�"�7ob�=��`���)Hi	�n�ـwnE�n�ŀ{ob�;#��#R�e���M$ݵ�n�ŀ{ob�;#�ݎUW9�P.�ҫ4�,E�SX����å��k���ջ)�+R"K�'+�To1°e�˅����8�'O+͘:t-�� ��y�m��ɺQٳ�c&�7cq�ϓ.z����ѨN�9�z��3�ꃃ��9�'��8]]�:9�����t,e�n,6�0���glya|;� v�Wb�b�p��/on�)V%Z�Ҍ�e(��2`�;8��P�.��]kH��
��z������3K¡D,-䶗Ut��K�:�,Hka2��\Pt]6Cjmr�R<�p�no@��ߖ�0�p�7ob�=�0N�1]ӱ]&��Xv8`��yn��=��g�r�5lI|�Z�v��X��� �ݗ�{ob�;�"�5W��TGiZe��ƛ0-�x��,�r,}0��n�iQWM�� ��� �܋ �G�v^$)��S.��C��;:p�:ٻtR1^06X�б�Ζ�nR�J^AJ23b�cE��r,}0-�x��Xv��!�I�n��X�8g�\���UDh���
�̹�3rO~Ͼ��sܑ`�5�E]��I��6`[��K�`ۑ`�� �l�e���R:t&� ��ղ^�0-�x}�j�.�6m`[%��� �ݗ�z\� ����ų�o�#(�E�l�͜�o,3���1�* vͲ��W7]T�TtvDn3��ğ?��v^�r,�d�U{lJ��+NҫI� �ݗ�z\� ��/ ݎwY@F�t�E]6ۼ�y�}�ܓ�߾�Ά�#�X�"1<!	X��%A�
!H���&�A�/�w\��y}>��%��
�t�m`[%��� �ݗ�z\� ��jЉV5I7mۻk ݎ��*�nO��o��� �܋ =[����;����t�c��@h��[��v�H87;sw����QhJ*���M'i� �ݗ�z\� �܋ ݎ��c
|��%N�	��=.E�wnE�n��v^�l�Z�˻e�t����Ȱ��yn��=.E�y{P������ջk ݎ����X�«�W(�*��@B!� �O@ys��5W�Ĩ��-ݪ�4�0-�x�Ȱ�Ȱ��}UϠ����t5��Fe���*F��+�Oj��0mę��-���v���t]�	������� ��/ �G��s�A�O� ��_%E��E+MӦ[k ��/ �G�v^�{}U\��O��h>����m;w�M��`[��Kذ�����+�*�.�i;M����l��d�}0ݘ���!�w�yM��ul��o���/ ��	 �*#���Z&CF��챐��6zm��6�BAn�+e�!�B:h�)�X�Ӹ�X:��#�A�[q݈Ӟ�u<�n�IE�5cc����!���;��sf�÷�s	�mH��.�t�\���+	�(Ԇ6��)!aIqe ���`�[�Q��v q��^ᝀV�Srv\�L�t�i��足ѱ-�8�F�y���t�A-�Yy�1�2k��|��U`I9��ɪ7=����ˀ2^�I�����N{`/��.�y��ε�,̶�QT�L��m�{� �\� �ݗ�yM��y{P�����t�i�w�o�E�yn��<���:�K�5V킢4�i>X�v��/ �/ ��/ �\� ﵪ�n��J��m�x��xT���Ȱ[��(�J��tRt�Zn��%��`�e�^���!~�ӄ�s!v�7�Y�\��d�n����P����ܽ۳m;=�tjP� ��E�jݗ�yzK�;.E�{��Bf:��o@�~�u� p�!!$I	E�!$#�'�I
l�R��D`�]}�nI%�X�r,۳-�C����x�����X�r,V��م41���-�;w�v\� ��E�jݗ�yzK�<��W�jպE�6��\� ջ/ ����v\� �oղ�+p�tk!���!$i��A'����❌���	ģ^��v;P9��Y[:R}xW����X��wZ���N؂��m���/ ��k��v^��Qs�6�ҽf�rN}����y��nl|"�b�^V'��W�^݀���cHvۻ� ��� ջ/ �E�vG� �YwE���4��f�v^�\� ����UR��_R�v�W��q���P��V������
�	��g]��Jep�<�m��w�>���zdp�=��jݗ�wvaMڦ�݊��ݵ�vG۳+ ջ/ �܋ ���\�EݴU�[f�ٕ�jݗ�ul��vGʷlD�e���j���R���)�׀v\���f`d�F!0�m2��#edI�+(`LL0���b1AMg���rO}�T�}������t�n����ˑ`�̬V�����Y�w�]�K�� ����ѻGs���i�y8��Pn3���w�r�/]�mӥn���"�=�X��s��>P�}���>�=pz�p�9k�[�7�2��Us�I����� �^� �j�Z��I4�ݺ�5n��;/b�:���o�e`ݙ`�|���M�v��r��s�yO��}�+ �ݗ�w�0��N�ݤZ-ЛXV�x���~I���I7�y�ܓ����W�h���
� @U��� _�  *��P@?�A�0T"�T"�,��B)B+BAP�T �B �T"$�B(�T"�B"0T "AP��T"�B �P��U�AP���AP��AP��	B T"�B
�P��B
T"�B0T"�B"���P��T )B(�P��B(AP�T"��B �P�B T �B�T"B$
�P�(DT ��B	B(AP��T"�B+B#B!B AP��T"B �P��T �P�� �P�,� ��,��B��T �)B*�EP��T"��T"
�P�P��B"$U���T �B(�T"*EP�!P�B$� T" DT �B �T �@T  AP�!P���@T"�AP��B��T"�@T"�AP�)P�AP��DT"�T"���B*
@T ��
�EB	BB(����T �B"���P��B*�T"P��B*�T  @T P�B*B�B",��EB(�P��P��"�P��T"�0�B(P�B*B($B �� �������W�  *� @Uh��W�PU��
�� @U��� _� ���`W�W��(+$�k;�� '^{0
 ?��d��0����a(�tAET�-*�w   P�@��N�����0�h ;�����|�� !�U2 `  (�( >�] � .��    � � ��:�  ;�   ���GN��V� �@�x��:u�C݁��檞�}�6�|@�h���k�ܪ���}-����k�U\ڜ  i}\��^�I�&��}�O��޽j��ǈs�t���<�<m�v�NB���T�`uy�+�� x���]�  SAK��v����7w>��ޕv��p_3=�P���M��@w��s��{5�;���}>g[ww���3�U��ְ v�g���>x�}��>@����{� �����6�>������a�@Ő >�=_Y@��� $dx��On���� i�{� g�zhw��7}6X�w��w4 /w 
t������p 5A̸()�`t�w���� ���(�  Ow�tr�
P-`:�����P�@{ޅ���͔ [ۂ��=� Y�@    ��SѠ� A���3��{�t�Gfz��o�� �ϖ����m����`>����[[8����x <A��Ψ�>�նx}�'��3�C d�`�G�ݭg�=�@�����:|�`( ���)o�u�N@4���{�π�g�2jGy�}��w�]��z��}�py=�s��(i����8   C��3�^Y�ί �� ��p�=�&{:z>�5{=���}���6`�� O�%ԥ* �Ob�U��`LʕR�{�*h��S�j��Ԫ��� �Ѫ�6�T   $�B�*R�D 4x�Ї�������I���?���׹��L�s��p��N���� �I��H���O� $��@I"@BI?�d I'����?�S�͚AsY�o?�?��7����'��ü+��������0G?n������'�`�G�s���G�ɋ��OwwN=����������Y�y�>}�s�~��.-�zf-ְ���������ϼ���u��o��5�H��Z����3�ܙ��M��Ϸf����1b�����}���)�hfnsZ��o�7~�?���~7�nM��J67!adr�bT�w���6����eݟk��$�M���(}�k|�n�a���~����
����ύprͱ �eu���~�>`p�q�[y���M���<��ߣ��\�ߵ��*�M ӃpDDJ6�8%��3�E�J����#>o}�{����ϴVl�� �������������C"�c,�PM�l?}�>�|2�5w�޾�R��&�}���nQ� ���f"9���0X�Q�LEj�H�I��},��}���XM�y���/���3��K�6)m��e��~5��̕v���9�������~�3���tg?~�V�B����������_�����Ux���No���m#YźfL\���^,_o���>���χ�=�Z<�s=����=�o��߲L�cO_��]��=���_d>�jǈ⛇�g�'m6���2�ٹ�z�����#��!����_�~�w�����9ːjn:7�A����ˣXQ����m��y�%������b��ջ������w���4M͊������o��m�^hsfѾw�5���o�{�Z�a������M�8ϒ��|	f�@Դ�`�7b3e�%�b��9y�O�~��#�R�D��o�S���߾�K������y<�����y(}�����W��̦k2�?o�7Z�Cy��)�$J`�%�	nD�M��6D�u�p֢	rhK�$ٜ��X�x7�?<3��>��l�xs��˯ܹ��3�����_������c����6�|�?}��9&��U��5�iv�56j9�n��Ʌ�ˮ~���-���y���R�z)��MMԽ_y��^������{�>�!�r?�|ϧ4�k��4}7�����L5��4.}�.\��+iq�]�k�`��$g�:�����S����MT�M�t�����^A���.k�w��8lώ	u����8������T>�a��oko܌�~�5��4�s����g'�\��d̩�6���͸����˟N��cKf�SZ�G�f�f�R���
 ��# �1�&?��������hw�&�����f!�{灾�}��|rq���|�Ǩ�5��t�~�Y�꟎����?~�k����
a��|�e�L�ᏜSfȣ+5������s>��4�o�������L1I�d1;�/{6����<�ϛ�������߳�~5��&�zy�ٮ~���Ƀ0�"JpJ%�.��ݚ܎��-�d�adaA/#��ё�\6Z�ky�4�j�f`���~i�_��[n���jS!�hK�n忣cL��5��:�4F�.�.��%�pe���6v>鸢�	2O��~733��W>�s�~%��n������c^ߖ�x9��_�埍�9�.�掇 �f��h�������'�W�x��A���q��}�^����\��\�m���j��\��qYrջ�,�kPBݴ�M�oe��=,,_��Fo���8#6�J%Дo�de�*,�h�]7��<���f�Zj�������Bј]3����s����8�'����|����{�]�noǋӉ�18�4{�߳�{����f,>׾�?�o��y����Υd/%����橈��q�aT�a'��4�x�Y�1�`]ᖱ���3Y�嘄dY��X$L�f@EB!QDB��Cg�n���:����7�x�Ò��� �h)�����F�2�A����\�5�����~@��H�t9�F�`�O��Gs�`��֜NnrSz�KT�fC�0`�B2��R�|?[p�G6o�o���u�ю�o1��5�
�����hɃ+us[�.i��M�vZc)�)��\�q����7�"W�EȢZR��gd���tȴ�.	62�FT��ýs�b	o2�9��9nNJg�QPR�%b2��q�e"Tb�%�tF�Ħ����F��2	5�6�!�ZF�MD�H��%����.kh��ΒC����L0�B�K,���F�pl�\n�0F)��ۚ�.j7Q���JD�@c[8�jnF��D��F��uu������i���ыw��9&��Q�0lj�n��|4p�����cn�y��v7���5��ZO37�HD��y�f�p�0��W[�MV�`��Q-#%�X0�%2��쫮�f�#n�E��8d�\Ѷ�{D�nk�8�s�X�[�s[�i��!.#s=w�z\���v	h�\F5��p��r��%����`k>�<ֿQ%h�T�h%4���k[mޟ߆������\:~�w��}���}��M�1�9��(�;�ކ�j�eX���p}�Jr0.A���9��7�0��9=��i���Ւ���`7H�7)T2%i��KA0�`�4�Q��6f�pqL��	%�5��փ��N%24��:Ӹ�r��!�֛,�7�9��)����o�t�d?S~�����&�oaq�v5.y,ʴTŴ�ś���Ї��ZYD��  �c"���)��'] ;���d���z�
@v�즍A��&��.��K���	L��(s
��&����)C T�!dJ	FFA
Lٳy������&D�	A� ��.M&e�	F����S&F��pf��
�!21�J2ȑh�4K~�8n�ҷ\&���4�6Ln�PK��e��h��y��g�+9����g� 4b\�w�Ә��*��b�b�`�mh���%7�%3Sm��c��5����59V	@�����ѯ�3rf�n�CJo%�N�]-Ǆ�����f�]��ɂ~��q�"Ze���#L�&7WS���Y�'�R�ʖ��62�5��ϓ�2�e}'�Zb2RjA�H֩�2��L��5���vZR���V�r�K��r3q�����0>/�O�S����3��"#?FDlS�;o�~�A�dd ����|:�4&�[(7#q��13M֢#�b��Ӛ�ٳ�.?_�4�3M�y�Tl]�Vce9��`٭^!_���sТ��p7���������+���ߧ߮����4�eHH2���ټp[3�8�٘K��	n�&��� ؕ)�m�܉A�Dno�O�ώL&�3_����%�n~���#?�	�5���K�A\9�4_�{�AO5������t;�}�z�~+tJ��y��}d�[�?�������o�Sw,�ܚDD˷*���#Ŗ��7�kQῂ�H���1.Q���ˀ����#2�20b���rD�P�A���d�	p�R����K��y��G��玹��؏Y����sf����}._xJ9�`�40[������#���gȜ���FK3��ô����d8���\�7S�\5&�����\8%�J	B�J�FY�L���o2&��~������l�������qr�"�P_پ|a��o�4~�p�U�,nb�����57p��j�����i.hL��+���9���%L.�͜���o��\�t�-���񽜗��O��=բ���E��k>��~���{�	L�w�l���+��|7q�����l�ƪ1�X-?O�˖2��2�A���c�x�noSy/��)|�|�@�߿o�f������%,�`��`7�#a�5���3��?~���Gr�o⟎ �j}�?p9r��IG.�L]D���������37n)��O�����&z�{���M�|��#�S��>��}�{��X������7T���������y�s��sAdr|<瞽2%���?��s�~^Ś?}�s�����ѿ�ϗ���?r˽o��Mf��Ø��̺�����tS�a�ύ7�]&<�1����6�I��+ɓw�d�ｗ3���7�h�b�!�f�j�cs�#�[�����f��;�5�����7�7[���Y���՚Ÿכ�}�~x��}��Ͼ�\�8Z����~l���Z�GV1־(1TϏ�~�����u�*7G"9��?\���k�������?~3�o�"JjM�74���F���$df��)&q`�L�\�K)V��.���55��jF�7z�������Ⱥ>�V�w:٨\�Uiu�.DnO�(ꅌ����L�Y�4�S5���l��^}����1.n	s�"���4o��� �y��7��G�s�����>��O�]��0{���dli�>NF�L�3�3�9�V���� %�XMm�LO�ǧ�i=�Ś�J���I7M��J_/���X`��	J�̱N�n�ʲ�1���STR\5��e�]�]����	+D,`$0��K0��s�������d�h���S$��A��fj�n���
;�nkZ˽�4�T���h̺JF�[CI�B�zt�}%�3�g�8n¶�7#p�n�n�`V�3�\?M�"~��ì���������k�f���Īԅ7.i��IWq!��2�I�5&�h	���~>p�×�7>�B����kSJ߿ni)��m��[�#sg\v]�ˣb\��4s�0�s��}���O�m�2�`����ễ~����j��9H��4ȗs�İ7�I�yH������W�}�f�I����cn�~�<�L$����s܏ߏ_��'�0���|�\�|��g��Zk�n
n�Z>��S|9�j%Ԩ���[��o�g%5����)���O����乡��JR�f+L�CS e�υ��0[����܃sw�K���t���޶͜#������7���s��&�
s7پ��w�?}�� C���?~|y������9�ѿ/�g�sw��Au�f�p^�"}�߸]��y����_�mX��#Z�jF�K�A4T�4$�b3:w[�1���hxo_����nq������W��{�Z��?;?"�كD�(�B��$�Kd�{Y���-���'Zw���D�h�3LǼ����r?�ջֳ��n�.HŜ��f��������%��Z���57�*!�	rR� �~&�~����g ��	L�����:4��ne�B���g)w��,ܭ)�MB�%I[�wu�n����&�%�*����@aDX5A2#-�"X�����5?R�ş�B���2&0CrQ��V=~��b}�]V^�P�M܍��}�>����h&��~XT��@��%sdH��Kn���5�~��Y�S2�~;ϞF�����>-s|���n��~��0ϒ��8��g9�&�p��o�_��o�[��55ĺ��61Ѳ��o�^g�۟!����h�H�B���&�I����~�*���*����UUV�������������������������ڪ����������
����������Z�����V�*������3
�=��U�M^nJᔻX:ËU����,�;orga�K�J��`��][�>=m(�ܘ:/ �sؼ�PR�/5v� `����m�R�.��*�x.XXv�S%��Ͷ+�cS=�UU�@m Z��]:*��5Q���U�`
��R���!P �]~����kf �hb�jK��K����.\��<x�۪��.����X�GU���QD��U\�m�[,Q,ځ�[7f���(��%]�����\�S5uR�fؗ��i8v=����jR���M���ҡ����6\������ү[<N�q��[e�w�j���h�N�v[�qltX^'�x�X�-(���`��Z,#a!ڌ�9yBa���(�d��H�s�-���ٴ�ٓ��uR�L6����uu֧�H�3�M�m�*u�(��UN��g�=�>�㟝ˠ(q-+�Gs� (
)86	Z� ,k��>��pce&sƞ�@v��p�d ����r���z8�ΐ�UU`s*���0n�6��Q�UmN�h��*�u]UUT��)@P\=��c�Z ��-+շ0N�t����ET��.l�M�L�H�W`T�5ՙF]2������l*ѐuմ�����>ک� ��3����Μs����z6&�V�DG�8�b�e��:j�ڧT����k��Maګ�o\Dqog�;c�ʼ��b땖g�����Q������7Q.�Џ�&]��*t\�	��^7,���[+�B�jRXL�+�i�"�.���RR�\���G9UF�\�a5]$�;�w.�L\ЗlM�)H\`�Yl�*��l�0^�)�r�2�j�L�uV卸.ћ�Dz��vZ�� �� �,ݮcj4������讙 ,NE�ؖ��Cb���`-��Q�����b�뚪�ڨ
�ȭ/pX̸��
+��a�� 5��
5	W`b�Ijٕv6uL�UU.˵tk8������������[�_`�A��U�8�R�6��ٻ.�+҃�E.�n��E�����H�u���u�"�.�kʖ^��m�,q��OnX���Zr��.��k��۰�	��DJ[K�US�����y3M����j�ێGi��N1*�i��\�d�V�؄�fJ��6&v�wI�7ST�#�az�=j9C�Y��,��i�6I���>y��`���oy]ڍ�ϼ�_S�6M#��ӕ�Ѡ61u]@@J��eH�Z6��U娥��r�P���V\Y�lUTt��C�g�s���*�sS�*s"ð5\�f�m�}��w���S.pA ������"Y��nUڶ��R��U-�e��Ek"�qZ ��[)v�PQ*՗ns�p�7q�r����ԯKj`��NM�a��V��*�V��c�m
��Q�Z�V�^j���[{F)pml�*���d[��#! ��p͋��S�\m=: �sGM�������}Ej�e�3*����W�{yլ����U\4�غ)R_n*���ggeZ�3VԦ\�GUj9@�6ʃ/l�%q3�qR��}�B�N�=�r�[N瓂��8�n�@ T�+λdh6�ꗲ����G9Y`j�*�:	ڊ��O#��9���\��m��9�s�2��Z��h�Y�ncr�)�.��vEVWt��N��m����\��7=eV�x�f5dݔj�r�J����a�UT�������kNܲ�=�����y%��y"�q��NQ��Y�єJ���sZF��m���ĎZȫ�WW-U�O3���8I�۵9���p�8���b��ݸ�\��>�!��G-�n�&)4�9�4	�x�gp�����lu �����u������f�v�"�F
��xN�C�$2��d3k��Ј\uٺRoP��^��
��u,A,�\Z$�K(�E��<�Ed�Gjy�����m]V.Si]��"2)�+n��ò%*��PX1	�Z��y���j��<��`[��4�&N�i�]��òL����Oi~+��V�z�IAEV��\�îٹ6wP�N��=m��$Y�A�v�j��Z��*�%t�cH�^(x9�5�&�	㌹�tEj�mUWPp���b�7������*���j85u�6�����/sv�{'='Cu��H�3S�bu�ʽ���f���>c�a�m���hG�.˹��z�c�N�ٖ�4,�f
�R�8Ë��c\aa��Q�+��Ҽl���imMT��:ɱ�N7N�j�N�y��{�3�T'����Pr`���ekq.���H 6.ƛ�8�H�ȅ��[q��\�)V ���l"D��ʭlں�' s#Y�-��Nm�aq�	��*��8�h-�۪�ī�`x�R����5�;�t����ǳ����x}j
˹�h�f���\dR�m���M��� �U*� �hX3a�A
���O�ۅCL���� ��ͫ����ĄRGL����� �g8�^����ŞMۘ�	�l�Uݚ[B�WR��{�`؝qU���R6ڲԲ�[ہ���zn5T�Z���v�'����P/9ғ����/��m�aBG�@lV�K��i��`�8�p�:B��U�k�c[P�����NP��YQ]�).�5q���UPx�j��U6w�*�[5V��f;p6���A��UmPuWAv���a�e�⪪���JJ�+<TYZ�^m�j�Z�*��(�YV���D�ı��j�p�6�m�V����	V�d�h
�.��6�t��6�`�Yz�6�:�2*��@[q��U:*�m�
��*p꺪�aY�\�����E��ͶQ��`����	�e	�2%ǒ��U���.Z�j��7eX
U����mW7)�j3�ڪ�������Y��޶Pj�4�j�U����S�UU�]�n�y�l\۞]pJ� ��$Z�
���,�0pݘ�ŔUe��^�A�k�G�i۬����l��,.������U�AK6��U��	+C5]��.�9B=Ex���� �j��bU���r���2�让�um��E+���(Y7��|�M�$uY�%j��+hU�yU[��V�yk]dq��e�䑎�*�Z��Ҝ�@V��@*��-J����Ԫ@�NyF��uUR��ŖT���� *1��h��t+k�S� mKQW@�;�̫�u�g��۶�j�����0t5p�0pV�@���������ks<��^=��nG��t�p\7��jYո ��ڀU�\�+����� ��ѥV��u�L2���AK�Q]�b�]YeUn�VV�8j煬v	��WӤ��tkg]�����M�ݳ.�������U�<Q��]���nݻ�uí���r�=a1:�Gi
iY@ڕC�ժ�Pmu��������D+l�Dx[8-�vڍ���+��`s��V�)�P�^m�떓;']ͽ�y� Cȱ�)��s���G�B�cMy+��}_U��E�@�j����}}r�+d5W7S��m.�ৱ4E.��ڪ���GQ�x�2�K]R&:y^��f��ӌ>f��z�a*Y�b��UU]���t�̲��T�-v�uUIPL�t���&�=�dvݭ�"j�svsi��LC,pQ�<a9�T�8㑦�UpqVyك��E)�f��`�*��F�T�Nr$�U�URMUlp&`A �U@�c.j��R��3uF�WUWUT���bڸ�F�\�����s!5[.���iv%�#uTڵ[m�.�ٌRg`4�1[K-:�=��m#�ĝ�P&���﯀��u˱,�Wq��Oɷ���Z����tv�.�`뭓�ب�+A��mO�ҽ��#l�"t�v��ʫ����օ �!��-�.�@b]��n4�#�m�����^O]/2��9��e�q���tէ�
�閊nqn.���G7mO,����X{z�
�U.[�؛���i)i�=��;m�����m��mȵ,: H�F�U��+���b�39�ؒ}aK6녏KT�I�����r���-�]��O#�IWN<�{Z�%�J����UP�]#�Fe�%O��~�;+���l�W��� ����\S���Z��:�����1+J��p�d��V.��J�Q�۷T�USr�U\�Q��\�4��UT��Z�tItt�UT�R�5˷l�UU.ĵU\]Tpdҡ�Uʮ�p�K=�wi;5�T� 譪�{5*��v��
����z��U��m��nl�5T�f�*Jǅ�;T6� psUT��2�d�kj��
��-FՌe��UUUUUUUPUP Td(�x=�Mn�I�U䍊���*���U}�ly䲐b��U�U*���U�ڐ�:��������<rn��������V`*��˱,�@��_G�}��iV�T�*ʰ@U*��:Z�
���6T����Q��]��[��ڕCg�R!��U�,x�YE���V
ڭ�=�s5Z�L������[�M�3WT�1�-�-�%��-�h��l��T6�/<�J�R��lJ�pf�mr綹
���(';����{i՞�n����U*����k2��
�4/vต`-�3�X���]���v�+ə�dj��Y+G%�-ѧ�H�Wg,������8�A�<>���i�3���ݼ�8ke:�r�vƥ���7�j��Wn�ԁ;m���WLi����]sl#K.�4کgX�<���X	U2N��U1D��-��R�T�{f�U5@U����mm+*��A@\�+��mX^��Mo.7�:Z���jN��[G�-���W)-^�7�+�Wha�];���wtz{�|��n�� R�C� ��B$� ��$@�d!2v���Ir�	!�X ��@��I ��@60$� � @���B�'�L?A!!��~��$���$60#	 0BAB�H�|
B�!�#A�$�u$��(A�RF��N�)	;$!� ��I� ~@?HCp��O�'�B |'@�!7>AH��@��6md�@�  
BrI'd�$���Hn ���jHnB�� 	@�O��@٩$�0��@
O� N�M5 ~�XI&HI|�6HB�� �	d%:I��BO�$���RYH|BBE��|HF0�@����B$?B@�Ą,���r5d��	;$	>�I�u#`"$b �Eb1DAI"�E"0*Db2@P������	�$`B !$�v���dbX�DDQ)A��Td �0$RY!�� 8I��Ȁ��N��D����gc$�# �E�T*IVB,#��>I��$HD�#'ıI����$�� �� �|I0��p� � � I$����HF`�@B�RBP�����N���Iӿ���UUUUU��j���[38V^p� �c[l�ۈj��q�X��
��F����+�Vd��WD�8��օNy�K�w
t@8ܛ�z��AQvK�K���'a��;]��M�ε�!�a�:0C=�
s�Z�0+��2�!�M�Rr��7ݬ01������o5�����d��8d-��n�9r��Ş|�p�i]� ��m�1v�FolRʒ����t�
 j6�)t
�(@q���m�nw�Ÿ;\��n0�l�q
#W���Y�q��j@4�%�]�ڼI����bS45�R��Lm��-˖4r�y��Ӽ2a�z^�Yݎ�D�2\ܺ+5/V�m�����î��MX�@����9�g�k]b��d܆M�j.�ئ/RO8����ayݜ�ӣQ�y0��xVmq��^'�a�5n ��+�3�J���tW�-#x�47Z����cT���6y�s���
�4B\j
���G�l@(2�0�͍̥KV��k����:�u���'�9��Ջ���uaj+2�ç�Y�^&���㔬��Q���v�۞=�������/j�H�K�n���9v�Z�K�ݼk\�p��G�ue�#Q�و#Kvԑ�P&�P�K�R��QsP��q�Q�%�Ӵ�y�6�t<[�]vZ�H�+.���;� c6�=+L�@�����`^��e��eeѹ��u��hKf�[ll�b��
Ufnˈ��,g�g�� ݔ-�8qbWsv&�eWk�@��@m�	��h�|�ˇiv/������M/��kWn�ѭ��m�ŻT�\�u�V������P�f�m�f�M'%V36���HX-��D!���em�ַ��S���r��@��ҍ��Gh��y�q�WW*�=��>�մ[`�h��@q6���Bݖc<v.�Ρ�;��8�h\�q��6�N�r	�·�M�)aeh�[	+��S���f٪,)�c����Qm��Sz�8'���ʖ�	�kX�c����C�@&��`HH		� �"�@>�� !��$�$�&�B!�[{�G7�݄�EG���/S̼��c�0�ӧf�$7m�.��X��ܸ�]�HPٻ4ŌԆ�BX�
��Vܨ�
��;S����)I�K@�Y����T�5��E)an(B�v��p4�P�*[6�ڛ8���m���8hq��ln^\��gn�r7DqGe�s���I���Z-�r�g��q��JݣuW��*�-��p$&I7!5���8�Qs.aW	���;o&˔���y9�t��u�4)�J�vto~����� 9��O��=A�{נ}Z�;�djDLM9�Z�Ӗhs������֞8�$܉����NY�Umz/%4
��@=��N�$��r$94
�+�/�S@�� ���@�>��RJda0�1'�o%4
�+�S�h^W�w�2�g����k��uJ�m�WZB��kv7H�r��[�Ƅa.׳�:-�3��zuNC�:�z���W���S@2𵵉�Lrdn= �9f��	N�0����� �;��sj��k��U�z�>�D�9�c����*��@���u.�w�@/K٠}��;�Q��O	$z���*�נ�,�*�+�=�\yqLD�&��nC@��^�r��@���@���s<̿���{5�:m�H��9�4J�
�7�wdy���g��(��aX�D�#����\�z��h}k�s�u�%�1!ɠU�W�_���U�z�9f��31#��u3ZJA�a2bR=���Umz{�}�g�$YE 	 H��iλVנr�+�kQ���H���U����Vנ_���e��_Qdœ��@>�,�*���e4
��@�aEh&cx�&C�- `X��HZ�J�c:�b!��74�طi�@�ЋX'3p ��Vנ_���U����>b�8а����@����<�31#���@/K٠Uy^���ˊb��LF7!�Uy^�r��N癘�W{נw�t��kOɂ�#bb��)�4
���y)��)0&� �>	���mW���]dJ'�#�y�4y)�U��@9NY�{K�&QD6�n1Adm�k�F�x����b[��L�ƃn"�%�L@�X��ȒNcD�dBrz{gM��z�r��g����h�z�Z�d@�)�G!�Uy^�r��@���Jh^���y1d�&F��S�h^W�_���U�z}|��R�A�94;���b����;�ΚW����>b�8щ���@�YM����r������4V �9�qw0��(j.�\ܲ��$v�Lp���s��8@�#k`�o���ڃ5���ʓ>l=cXE�.t���-������CC@P�seܺ,=��F���pb�j@���-�	��*큑:�P`�˷��`8!{L웢)��j��kR�D��Z��5Ƨ��k(�/�.ݸ2�#ډ��\�U=��.h�-�In�|�׻�>w�x��1s��U٥�N�n�,���ZT�.k����(&�Eɳh�2�,2��o㽯@>�,�*�+�/�S@/V6G��F�M)�}NY���1#�޽���U��@=ϸ
Ƣ���"X���*�+�/�S@��^�}NY�s/^jI9�	�q��)�U��@>�,�*�+�9p�B֔ȁLS$RC@�� ���@���Jh�;��Y���	rk��BջK�m�Rl��HL�[���	�@���% �e���$��&927����*��@�YN��瞠����*�w���Hxc�D��&��߻���>y�4A�MҖ��(�
����Q����
b�'BvI��}��~�Ɓ��נ��4|;��� ���$�@�YM����9f�U�z�k�`�	2"��hw3<�]}�zۗ�@���e4�kO��bdq��h^W�[�M��z-N9y1�$�" x��tt�:�%�ٱ�����pݴ�c��H��çਢ�2B`�s@���@���_Z��k�2�U椓�%0��'�o%4
�����4
���n�Zڙ1b��H���Wֽ ���1��NB�Yۚ�m^}���W.s-bLY1ɑ8����W9^�y�M���,��P
d0�0���W�����*��@/9T�o���u�\��vs�lW	U�
<Pi6j�J$�H����ڻa *XXNH-��RG�^rS@�� ��M���|�15�1'!�Uy^��� ��T�:�z�y)�[Zx��dQ��q��h^W�[�M���ߎbVD� H@bR)�[߻�W��]v�o~�mK d$�A'�O:�o�ӽO�YY�go%m�{�Iw�3�역��Iw���}I*����߻���j0V4���֥�e�؎��t@ֱ,�2�K�M�Ky..�`��h�������� �w���V�[ԒVݧ���˗%bN���I%nr�}I*�+z�J�m=� ��wo �?���V�3*cL���U�V�$���{�IV�[ԒJ������bV��h������o���o��I$��Y�%[�oRI{ȸ�h�:��l��@;���� �g��9m�������������I:��qowq%��)�Wl7CT�&-�V�Z�Y�
�Bd�\�!��直��t�<��;a�!K��\�X�2��KV7����#�R'&�%R�FJ��BVic
�E�#/9�a��l���c�5�9m-���ye���lUm�؟;���M��fM5���Hj��l����źADkq�j�:��mi�7Hc��|_�F�Yq�����{4�|��ݺBwOV��p7,��Z.�A�ǎ��-<�����Xр���V�l�@R<��W�� �O�>�ݾ�� �|�����v� =���bj�qQ$�Ԓ��$��O}I*�+Z�I}�޾������gZ��v�[v���U�ZԒK��{�IV�oRA�e�����1*�o��wu�<��9g���n��$���{�I,��UK�7�bg {>��۽�RI[ͧ���vV�$��9r�RLD����H�lA=KR�����Sp���4��px�ͫ�`��nfeLi��@;�kz�J�v���U�[��y��g���n^��~���X�M�h�;x w��u�?�!8@$�j�3��ݶ�ޝ��۽��ߓ��]M�uֲ����n��$���Y�%[��I%~�v���׸�Q��T9�� ��l�Ԓ��ޤ���O}I*ݭ�I%���˱5Z��W�@;�{����{�IV�oRI+̶{�Iw3�\�f����Eh�����m�<\A^�m�n|u�P�=���*��ہ�Z�U���<�������Ԓ��ޤ�W��=�$�v���g�lYu�J���@;����n^�}I.�޷�$��i��33l�e������ ���}��w�xrΟ�s�,܄�x�G�m^�Kr��@1	g>��2	��o��f����AD`Ōa�p��]o��)�9�A�׉'��f�e��r�8e�g��{�^F`�s�?E�,Eu���5���fܣ�c�\��a��w�.�;��"���	fkz�����\9���.��a9����u��Yw�`0@`��F"2B� �$�X��@DP"$c��!�3;%��$�8-������A' j))!h1DgF���)lf�(�pkl(���ab%�1D�#�PвfC���7&��2������	��9�'⴬������R�f���fƛ0��f��^s�����R1XEI��P0�'&��g������ka����hY��_�g,�Ѳ���?��9	$� orO�$	���zX���r���$$HX�X@6O�$�$<Ͻs�_s�RK��֤��ϹB<M�9�M<r{�IV�oRI_��=�$����?rNI����Ͼ�|k���&
f�&�z�J�o��%]��I$��,�Ԓ��ޤ��SJ�m1�����0�T],n!��J4��aD��є�kj�����LD�������ǀ���_} ���߹9�v�߿{=� ���j"܁�q� v���@;�{����=�$�v�������#k���'���[�[ԒW�}�}I*ݭ�H�ߺ��ӷ�O�-���o��[�{�IV�oRI/��=�%�{�w.B���! �YF�D���$����y�f�����OY@ұ�s��۽����$k��~�m���k7m���l���'����2���[f�"'����j�]���WV�h"J9%�&%[�9!28���$��9g������$���s�RJ�������u)��3*cL�� Wlz�J�o��%[��I$��,�Ԓ�&�@��%��Z.� ��{���vV�$�����RIWlz�K�E�q@c# L���}I*�jI%�9g��wz� �w��} ?����"܁�;x ݿu���ro���� ���ޜ��3��ݶߡ��B��DH'w~�(~��&�����`MkN�aغ�l%��C��4�;	O\����+���q� �m�l��Wuۂ65\s�0 �v�7g�׎�5��(&kYt�WF%ٌ��$���W�����e�6D��ϑ���n���\m�z�0�&U-��Z.;)ct�p���V[�.��^V�֊Ba�ҵ��[ڴ�� ��0��s)��Up6R��zӤ���{}�_V�!��������s��uV5d�K)��X"��	xu�Oj�vW�\M.9�6�K$��U�ǩ$�-�=�$�v��$�}��@>��q<ɶcY�+����群�n��$��9g������ }��t��f�+es=��w�x�I[���RIWlz�J�_s�RIe�xm��Aɢ�� {>��wz� ���=���q�����CJn93C�.�s��{��v��$���� ~ߟ�� ;��_} ��R��#�q��&���p��&�U&�M1��%��bESc,2q.u�2��w�{�}��$����$��l�fg�|�K���RIr�w�Fc,F�M�=���q糒D������ޛ��r�os��n�o{��翤�9��W��
���0.< ���{�I*�RI[o��%]��I$�����*�ͨ_} ;��x ����Ԓ��֤�V��RK�lK5ɶ�ѕ������}���׸���9f��v����;�������J]-��-(X����cK�Db5�2\�ӑ�\��[3�k�r�� �������h�ՠ[˹�\���Lc�Q��I�r��@�v��]��ڴ�}�x'�f8m�M�ڴ��ٷ���3c����PYD���@�"��D $D�dQ��� �F����y^���٠z�����n`$�Z��h�ՠqUl�9]�@��㠞8�$�3s4Wj�9Z���ՠ[n���33�:��qM��ɗOt%�X���e��!������W�D���Ce��hʃ�n�O�~�]��9]�@�����h�9��XL�,�0JG�r�V�m��+�h�r�켉eq�ɏ&�@��s@�v���W�r�V�˜�����d��f���Z+\�E���ݩ'd$a@@I�jd�1�}���Rc`��L�E�r���Wj�-���9]�@�fy��_���ma0�M\h݂b5�ǌ�v�V����� v��Yb5Ё�6�&�~�z�ՠ[˹�r�V���+�=Y�RPk	���MŠ[˹����H�}��/Z�z+�h�|yq8dq�f6�h�ՠr����f%z�ՠw������ĉ�q��qh����ڴ�]���b����̸.��ŋ	��Wj�;��y��������]��s��m^�Y$D�`D@�0�FAI�Bg�K{��=��`X��)�*p�6�
6){.�r4���`�.�98cz�&ph�:�\1���z!�>x�Ki�$�l{Tv^�R���qۿl�c��].]ץF�8��X%z��M��˰BV*�4�aҖʛ�u��h-/\u���ZJ�1��vvܝݶݻ3)��a�aXs6�-�Hq:W��+�N4��3����r��h��.e�O�ބ�&�1�NRi� )�o���<�lΩz���n�2�Z�n��V3�K{i�:����w����ק��v�����3�P^��h�^��3#	��9�+�oq"��נ^��h�����Ď�n�ciL�)�ȴ�_^���ZwĻow4�ޭ�r�(5��$ۏC��3��c����h��ۚ+�hw<�W�^�嗽I@Ǆ�50n-�]��e��W�^�z�Wj�*��OǒA�2E2��m(��a��f�Y��@�J�j�2X$֋�;�ך��7 L���@�}��9Z�z���<�{{��^t��D�"˗Y��~�_���D"0���"�5�H@�� Ē�&jH�g������h�V�33�H/2��$�G,`��޾�h��i�<�<Ļ�ޭ�e��>����bNd���Z����{{�h��Z��z ^�^�ڽ��an��&hth��k&h�ՠ~��y�y���w����~����ܸ]X�C#O#<�7�����[�h�{83:�6!I�F�.i�Y��t�=<J�F7I��L����/^�r�4yݞ$$�^�=�~���NSN��\RjG����y���{��^��h�Z��y�$|���(�di���rh���j���nܒB'�B�Y$�� �I"$BCP B׿5�����f���H�J@���m|H�׽v�}��ͪ���[_H��}���:<Bd�$�MG��U�@�y�+��z{��h�ՠ|�kp��s�*���R�1@ka�A���S$b��	�� �^ �wI�OOaG68I�.N?@/{٠[˹�r�Ws3�Pw��z3��u��x�Ĥ�����<�H�}���/f�r�7��E�^�㌙2b�G3@�}��s�i�<�<��獝����?~������ڊ6ڙ$ȜZ���K��٠���-���| �'!�����MI&�����h,���Y���4�ɠ��W� B�������]�����������%Űt�ђ�s����
�p�4vkl8)	����j{;�Gɟ-�`S�	��;����ڴ���3�3��{4��<�6H��H6�h�ս�33<ă��٠���-�����;�=��}4��W�5����g�_ 9m�w����ow4�ޭ ��̩�S�$��A}oӤ�����}��o߻�s@�v��y�~����~������8�'�c�h��h��<�ٙ����/�?~�ߦ�r�4�_��3"^���Z�f�0s4��?\N[�������7w�P��S�����7D�>�5�+�Dl�s�5�cl������aJ3�Ս+,BX��V}��iGe~���]��7c���d�]s�8<C�I2e&�98�`]g%ERn<���[�ɒ��K ���怛�0ݤ�t2,��+U���H0��� DC9K2L�+0���$� ��Ob���p*P20�cA�U�DQ�k��SAX��6UDa�&���DDb�$A�<�y�L�5\�57��!u
1�,�liAd��C��亊(�H��2�\���j!"(�����s+��h�$�Є�!�q/u��ͷO����Ut�U@UWU6��i&:n\#��5�i��'�M���C���F�#��%u�!T���[b7�!N�F�vUr;���9�}C@�c/[mW:�sv�����/�u\�Qk1�&fQ��la��10f�`��H4�eֶ���Y}�1�\M�B^���ñ��q�J1�'�;��w(֫��l��Y`��nm��l;�6�D�ݡ]�L$���jgCЋX�mhz�&����s�Ý��r���#ksZ֊����X�I`P��m<谦�2.*�h��{t�16�Տg
\U�
����Nye}`�S��L�ӊ�����]���;(K�UI�e���p�O�mu��ŵ±,a�)ol:�w0��&ȑ7�b��`|��j����,�'Eb`��d�=����m��Q'�w�r
s7(q\�7/b�)�����`���v�mm�	�Tư���J�m�@����Uy�0R"�E�Ж�(�;J�,�q�����k3ف��� ԉy����e@N�W�W",Y�����r�ǜ�OnZ �66bQ��شl�N���M�:uii��mА���|w�|c&1���2����ɴ��0�&�g��8-T�+q[C��1Ɔ	���[�Y��٘��X��n���O���v�����;
��Ϣ�����<pD�з��+�ٹP5�7Yyű�V�kAfl������F�V���mY����I.x;]�c�#�^l:;[�b��a���XnL��iݖ���md�S�(�.�h*�j=J����fԫ�j�t�,n��yS���QtS#��{=nN��Cq5��nzk������X�ʱvR�Xg��~�)XA��bQ�Wgk\uh��:�J�>݌�����o/HL�BG)�o1�=��m�K=�1��B䎛JQ�%�&�:����{V�'���lڬ�J�/�)�4}��N7��r�٭�1�Q�Y:M:I��z |��!I�HOH�$=�! C����$� O�:N�o��~��ZT̆�d�a�[w:�69�����=�+���hR�g@5�4��ٚ������,��aǶ��2j���k4db��h	��m�Ln�ڐ�s�����[qT3���GN㋛ev0�4��4p�n�$���M'BmӴSՍ��Z��%�*ŶS����MR�L���K(^lTM���Y�sJ1@,cIp�1*�fn��'I�?�NO=�� fY���`����Z�`E����m���F��Z���t~��z%ބ�22d�$�g�?~�- �-�+�w<�Pw������u��m9�<�Š�{�bE��V�����+�os<H��^�G�C"Ǔ�ǒM���@���?��������߳��z���K$i� 7�|������z�ՠ�C�g��e��9Gq�q�E�@�3@�|�@�g��N�z�Z廛m�ݽ���%\P�����!�H]�$����j�*1���np�'��_z�]9�x(I����������y���<�����h)����G�N<XЉ�m^�>�ރ@A"�(�Y,�IaR ��,�`%��XI'�w�ٵ}����u��߂�3��KsTsѢ��ھ��ٵ-|�N���{4�ޭ�9Z�d�jd�#�f�s��w��h:^��ʴ?y���<���f����	��A��H�'�}NY�w����^�@�;���}��o��;-�MX�k�ٓa�P�ah��U���1W`�5qi�M7OΒq�>�$��O#hrzz�V�~���-v�$?��+����m_���������&r-�˹��3�Ď�ޭ ����-|�{癞x��ǝ��H�ɓ1\ѵ}��������� ��I	�w�z���s@�)(����o&j��$	�	$Ͽ�}��W��=�v�}ݞ�쓻����}����+��VX�'��>�y������]��=�s��o���;S]2�)��l�����u �;t��X�l�ڠ%u�~N�OOC��q`�9�qzy{��Z�V��k��333��Z�^�-�� 9��%&h�U���<�#�z��z�������1#����I�H6���N-�j���էs�3�K��w4�ޭ����:��t�m����:w�ӧ�{������ͫ�s��_�	? A$Hv l�'� �{����ڿ����m�"iHMŠ_���?g�~�<�<�����]��Wj�/ԅq&��c��@��a��.��҉���U�q����5�T������+��ɲE�l�m���V��jנr�W|�<�3=A���h�I��1bq��
E�}Z����?y�&c����ڿ���ͫ�s���	j����E8�ɂR=�ޭ���=�����_���ͫ��N�75GC�2!8�;�y���{�s@�w�@����;�癊�^��;��� 9�d�9���h�<���y�������~���h�w4=�
ָB`9��xғ"Y�⥱c�ks:c�����L����攲1eKmK52O��;<]p͝YݝϩB�l��u8���w7'J�z�AmHi�/4(Qu"�j�K;[�g=0r+�Vɝ�7�W3v^�s�H�8yËX�K�U/f�n6�v1��(�M��ISLfӱOclnXFۂK�v�8v�!�� �cL��`�,)g`����@X2�4
�Q��:I?N�3F'��`7L�qc��]��.&8�jͳ�h,���j�kE��U~���o�14�8��\���נZ�Z��g�*���]��׾4�sX&iMU��k�h�]��j�=�r���,�z�,�<N`4�Zy{��Z�Zw��ľ�W�@�_z�}���'�q&L��4;��.�w�@�Z�z�ա��<]�w���t�#(���$ZծW�3��3�����������s@�ڴb3��Y�,I�qF��ҥ3Uu�v�Fq��i�vMHRU�]��q燓\�)��E�LJ9=�w�@�r�h�U����U��9��|�qa1㙪�j�^��vorHG�� �=�{�j��{�m_�������L�������4jHc�"�f�����|��w33�}��;�����]l�)�<�š����o\�/_z��]�癘�gz�
���m&�xc����+�h���+�h+�&��υ��Vx��v���<�fNE�N�>�v���I{vK�ٟ�䒓>ZTISEa1�{i�{��r�V��w3�<�z�ՠ}�:g��uMK���6�{��߈@�����Z�.��3��;zN����BH�.�ɠr�U��y��VDaY$HD!"H�I'��$�=$ ����W��v�����\��!�U|zN{|�{��r�U���������4gq���0��L�N-�s@�y��{/W�qw��@�|�@�.s.�#m<�Sx�VT%��I��Hn��+���e���u��R)&FL���$$Q��9_*�>V�4Wʻ�y����ow4�z�m�14�8�'��ٽ�<�/]��;�����ݻ��HC1�=��\���`��5�b�@����@��sN癘��Z�z��m�߻;�B��#��[��������j���]����!$�A	�x�y��oV��c�����f$�h��h��4Wʴyw4�gq�B�+��3S	���ҕ�1Hԗ5�@YK-��vf��T�G�
�:I�_z����R]	"���ߦ���V�yn�|�3=Az�V�}�����fHaE&���V�-}�}�j���]����u�����f?c�~h�@�D)������ڴ�fg��{4���@�i�5�p�䃊9��<�{;ՠ�{4Wj�/��h/���&�qL�E���4���{;���{��r�V���߯š݉o�!7*Zꠑ�D�e"�.��WM.���j���\����[���Ւ����L��Ű!��`V��kAr���k� D4
1�
M��׌� �M4�ZY�fe����8���Շ	ඃͺ���x�n�7-�tZ�%���BB��$ԮM<Nk�&����lKg�:�"Mn����6��23gRg�V���s���_�CbX1dl����!.���V�w,��%Z���q�5ڠ��K�_9%%�lX�����uh�w4Wj�ffz��������A	AǑdmŠ_����fbE��V�v���8��@���:4$���M��9]�@/2٧|�<Ī���;ow4n]��H��1��z�_��}��ڽ��j���ͯ� ���1�����e�~Q̒Dc�a�&��y^��3<��o}�@�w�@/Գ@����ǛM��4���M�Q)w�>~�2�u�Mȥu��3K�"�ެ�x��k��&D���;�z�Wʴ�K?ffy��
�z��w���<�q7�˟v��k��$�L�d��%��0&�����`��İ0��d����#!	�H֗���������ڽ�}ۿ���y}�m��R#�hyӳ@⼯O���Hg��{��_g�����}�\�����0��	4+��_*�9_*���}��kj��|z]i�]f��u�G�Z�Z|���32�^�@;zvh����ޜ�wt�L.)WE���-�e��"�,Ų�,��6��`�
�ٍѠ蟓�t��:=0$���/@�w�@���E���o����g�v����2Z]bf�ŠU̵���h�ՠr�]�I��� [���|#�At��+�;����*����Fa�dƾ��Ɯ���4�bL�d��X2DM��F�%��i�w���/&�(|OП4�� ���QO�o0�����~�?~r����7�K��e�蟦�"����X`"d�A ��`a��Zi.hnC\�06R�Y���"(������@Ad١� i��� D�c"P���H�0%6.V�J逃��$Q#KJ�,e�iXQ��L�H����2"�;,���81�~��(�	#a��'�V
Ͼ.:��80�",D3&�����~�
J!`"��!�$�	����� �!���$� ��HMHBI' �6H`@�6@� !�����Ϲv�oO{6��|u�b�Po"�C�g���n��/]��*�-z+�Z�L��c#�,�pN+�Zs��ξgz��ޭ���SyM�f`1�S[���.���یuE��Ư$���ӽ<[�J	����ɑȽ��޽����$�	'�_g�������Z���STвcx��9]�@�䦁��Z_e��zwt��g�g��u)T[�|��ם��s����?�$��ק��m_g����g�oƤe�)J����'u���]����f����ݯ��BF2D�y�x�o����q��)�s8G���+�;�y�y{;���t�9]�@���S���L݅vq�SM���E������*�΁�,���*�����I�o���6��I�IB?�����@�䦁��o��9W��>ͫ��:yu���j��4�"�9y)�r�U�q}J�Wʷ��fx�ܴ��ٌx�D2'�ޭ��W�s<��w�@����rл�03�1zߺ}���������㿖���M�����ۏ��cp�@�|�@���<����;����8��W�~��<��Ѿ���?df k���ƘK��*�44\sG�	��	s#�%s�i�*�7l]aAm<z�:��).ۙG^�1-u���m�lۂˎ2��S�t£���"*�K��]�5��ͱ3`[(
��u�5i�� f�f�[��+.�m%�A6��nw�!๨殲�\e����Q3V�][�� �d�h������Z�N�w;���[w���37m�,&DlfJ)MX㠱l�t�+f�-��HĖ�?�z�s51a0RI�"�}��?����V���r����g �� �I�!�r�U��31"�gz��ޭ��M��N�<B�x�8G�W3�z+�i��3�l�^��h��ǉ�#�4�H�Wj�>���9_*���e��>���&)F�!8�o%4�y�^���r�z+�Z9q��i,���&��ěl�E�V���m��7���2�.�\%.h��ܑ@��D2'@�w�@���z+�_�3�=A�{�����i���'3F�5v����st���#!�I	 �,Ha �B<@����r����h�U�p���jLy1�G�Z�V��sN�y���Z\�^���\����)"@�qh{��31��� ��h_pP.ff.Yʴ�����$LF$�h��h}½�ڴ���/)A��9!ڎ
Rʑu�� ��.�^��׊��{\�f��D#�'���l�!dF71��zW/S�-v��)��3=A޾�h�P�Ss��=�j�/,��k�Z?���$�/����fsDр��}�k���s�ݴ�A�@��O��Cz���sj���]����ۻ�Ǐ dC�p�-|�@��T�_*��g���{�4��ո�D�72dr-��S�;�y�^����gM��� �x����%vB����-vF�b�����]�Z�뮲Vv��Y�歋S�yN�G�ƤO@�|�@�������3�3����{�=�;��",2`���i���w7��y癉��ZW/S�9]�@��|�G�"H��I��9]�@��T��y�g�bW��Zo{��_�(�&!��#�C���y������ޭ�w4�|�33Ö]Zώ*�C�̙�r=�ڴ癙��w��^��h[^����T����5Qab�
�Uњf�Wc��l	s�u�=�Jb{]���{��O7���f�tF%2{m�����i��ZV��3<�=Az�ՠw9�;�A)���sNf���s���?��3�����;����m���g�~���������ji�9�䍑ȴ����@�v��w4Wj�P�����!��r����}�{f����ݯ�������,��ؒ��(����/-�ڿ�'}�z�_^�ٵ~�w�j��$dH���@d#!".�N5T����a�����a�D�a��+Hx�)k��2�7%��f�SV�D��l��.��-�L�����Nۂ��W� a�!�S�c5�ҩ6�4��Ձ�HZ��]ba�x��9l�ҹWvb7f���9�!�-��T��!��uЗ��!f�lH�8��K����m^�/	��s����=�q/�� �b�����eg�99�$���o�܂;�狮�ź�&�Y� �)9�5�ฯ#�%��R��m�y�)&��U �`0����
��@�v���h�J<B�y@8G�W-{�3ċ�ޭ������[��H/
��M�2<��$z��V�ye4�٠U�^��X�F9�ɓqhw�1v�zmW����{~�sk�I�	������W��2/�$�bɉ��h���Z�]�@���˗˸�Jy��)H$,(����`	x��\��f���
5Hf{�<{���L�$m)$��޽�ڴ�)�3��?g����~���Ėm�yѦWx�����N��t��ٙ�����f�W-{�ď�v�IG�Gn-����m�~�����;�ޭ�c�:<I"H�L����]�w�������V�s�]�{�h�G׀��
C@����y�w��^������S@��-�A[4�9lJ$1ΊLԨ��]9닅�g��:��� ��7MZ�2dy1����}��-�s@��h[^��X�F�&L�R-�w7��$^�t�:�޽�ڷ��$w9�'Y�<��sZ6�}�yڽ��sn�|����$" ��!�Dd�5>	޺��@����rۋF�dɍ7 I!���<]}�^�z�ՠ[n��n�p��&,m��G���Wj�;�y��w��^���Vנ|���
���.��:�6�:�ܸ�ֶB�̡z4���7M�q���+���(�ɉG7�w��4[)�U�^���Z���tx��I2<<���e7��y��3��˿�=����@���~���X9�&�AHhrנr�V����3��g��������OƁώ*�ci5Q�b�=�y⽝��}�������]��H@d��R@> ,�5��{�W�\�;L��4f:��V�Wj���n��!�$������˿�=�ڴr�.�"��6��m���z�2ް��	�P�06k�h��2�E#�q�p��c�N-����k�9]����z��}��;����jdƔq(���k��瘑z�ՠw��Z-���<�<H)·I�nG����ޭ�j���x��gM����=Y�*IFa0��MŠZ�Z-��*�����w�@���>�Q�&9��qh�S@���Wj�-v�$�}�jۃ���1�4�V- �[����,]Q
[�"���PV�
���DSt
1��l1�lۤ8R��NP�A̴#D"9 %���!ąc4hD�6��f�XNH	1����� �itj�h�FG�'%)K"���E�P`� �0`�$0�R�(�)�K�n�śa���1�0Ԙ�bA��A�� �,E�#��ý��6Ӫ�����UUb�`��b�L�ӻsѴ��au�W�6�/nzm2�m�x�|zb5L��7%�,���lu7�\����
��k��[���y�vB��I�51=��T`�ƢDf5#�զk��dR�"�mn��hz��sPZ�& �Q1��M�j�`K�rm�,�/ZC��#�v
����V�&e�����u�E�r\Rh���Dl�R(��l����6C.��nҰ��l87B\t���݂�pg5�n��x� Ln'<�3͐��/��;��{�J�Up2rfz�7 �x��E�tM�֚\��:��n8�v���x����hVҘ���JS^\�0�B�-�%��F̺jh�mmP���V������I�Ll����.�Av|a{%�`↫�\vU�c��I��=v��:�n�»��9C$���;��m͉WkZ,����x�:׋x&�o]���c�Ȑ�m��A��U�+�	SW�7,�.�·E���4!4!h��b��͍c`��j7=)EFj뵞���[�=-\�ˮZ�)����ռ��U*
$+ �l�E�y0�Mas�w"lxŗ��TkL�I�݇Zm6:�m�au˜i�fB��f���v���"�vL!�]v��f	',,��96���l��C`�lď�;�����m��$g9����nt9\aw-�!����o�z��Awe]ݬ�bQ^�[�'��糢�FT�qeΥ:f����������X�Ca3�#�P孒�8!n4M��)$6s��GL���uM�S<empk+��I�h�c�,6.C)��l�\[X�np7Vbd���ԅ� �׋�ZC��
���.�:��f;\O!w,��:��7KBl��r뇬;:"�B�J�Ts�TV����x��b��>zm@�h�e���U��A�f7`˭�ת<X�:«۱.�Yz�A��,���7V��SSWm��89o8�79t�ԭ��(�rb\; l�8c�wp� � �I���	�	�!�}	��	��r@�� ����HI
@0 ��l	�U�g٭Y��!5"�C@��`���vc*���q�e����Ԃfa��X����L�Xꔰ0��0h5�)��`�1����Pky��[v���q���P�瞦l�#H����Y�Ԥã@ۘ�%�tv{8��b��q*�;c�Ld�ў�r׭dK�Ȇ�l���JZ�r��7,ؔBݻ��:�stٮ�{k�6�q`�{�9	9Ì�x�[\�e�Ѫmj�Mc��4�y����ŁV�Tjq_�2=��x,C��AH|V���ՠZ�_��3�����?i�����j$����z+�h�V��e4
��ffg�31��E�	�0�2!H�ߟ��@岚Vנr�V�s�W �2!�� �4;�����:�޽�ڴ;��n��;������F����^���m_w������aX{�ߝÌ+
°ｿ;�V�d��߿d�"\ȓ]�Ĕ�����a�*�3jHU*�$��e�I����LR���U˚�Ì+
°��]Ì+
°�{�;�V�a�{~w0�+
������V�a��妌]�4`��w0�+
�����FN��d�a��}���8°�+�����V�a�k���V�aߍt�8]f��pQ�Ӹq�aXV�w�p�
°�=�{ٸq�HV�}���aXV�����8°�+��Xڙ����sF���aX{>��p�
°�;�w�p�
°�=������@�;������aXw���T��Ks����N��N��{�q�aXV����aXV�}�p�8°�+g��naXV��~�OS���]K�ݡ5��4�hհ���ck`�aE$�C�H��5�7KXG75w0�+
�����aXV�}�p�8°�+g��l?��?0��a��]Ì+
°�?���Ɯ֊h�FkNf�Ì+
°�������°����70�+
�������V�a﻿;�+
°���Z�]2�ӫ�70�+
���}��V�a�k޻�Vl�@`HȄ��@0���w�;�V�a����V�aN�w���Mb��kY�q�aRV���q�aXV���q�aXV���p�
°�=��p�
°�/���i�M.�������8°�+}���8°�+'}�p�8°�+g{��8°�+�^��8°�+d��\2�5�i�j�=2��cb褷kW.;]�28+�n���meE2h�6*�t�t�Jt�N���q�aXV��ٸq�aXV���q�aXV���q�aXV��X�㩬V鹣p�
°�=��p�%aXV���q�aXV�^��8°�+���q�aXV����f�.J�V�w���B�������q�aXV��z�aY+
þ��naXV�s��naXV�ޏ��j]��4�|���N��'N!�>�����8°�+p�8°�+�{��8°���H��H!�v�*�֌��n�r;&�F�nj��@��w��!�X
��jE�QOBN�!>�}��߳p�
°�?��'��0bd���^B����~�y0�+
ù��70�+
ù�{70�+
����]Ì+
°��ݿ3����s�\�������H1Hg���J����W���޵���c�n�h�8°�+�{��8°�+���8°�+�׽w0�+
þ��naXV�=��9�Mi5]W5�f���aXw=�f�ĕ�aX{�o����aXw��Ì+
°�w��Ì+
°���ᦥ47Y���5��8°�+}���8°�+���q�IXV��ٸq�aXV�����#�G��3�.���c��H�Ӹq�aXV�}�p�
°�/��kp�
°�;���p�
 V���q�aXV�y�diu�b7Nf�Ì+
°��}�Ì+
°�{��Ì+
°��ߝÌ+
°���V�`�~ w����%�J�2�TK+)�KQ<�3��u��r�`%4���������DW��X.k��;P&'�4�ij�WvyB��S��7>�<Lj6ZJJ�Ж6��,e�0Tz�!���- P� �Z��6¡f-⎥8�c��`J��R��Ƃ�`���A�A^7nt��ɞ�p$���z+f�#��,�����jL������Z���������:��Ճ��˷g&��
�U�v{��ú���"��'S=Se�3J���_:}:S�:V���Ì+
°��ߝÌ+
°����1�aX_�{�[�V�N�����Si�+4i�Ο��N+}���8°�+���q�aXV����q�aXV���Ì?�$�zc�:����㪺۠�.O:|:V�a�����V�a}�{[�VRFJþ�����y܂�Xv~Ꝗ�7��m ������8°�+������aX{�ߝÌ+
°���V�aN�wخaSF��:�kp�
°�;�{��V�a��޻�V�a�{�70�+
�����0�+
���S.x��\tX�3z��4O]��v#�s�j�
XU��Y�k��bh�.����,+
��׽w0�+
þ��naXV��}�naXV�}�sp�
�N������2c;(�Û�O�JqXV���p�}�#	Y�aX_k�����aX^������aX{������L��������Z�5�sNf�Ì+
°��������aX^������aX{������aXw��Ì+
°��[�hˣe�b:�Zַ0�+�1�{���[�V�a��]Ì+
°���V�a}�{[�V�a��wɫ���sFmֵ�q�aXV��q�aXV�}�p�
°�/��kp�
°�/}�kp�
°�>��|�F9m���.+s2���TR�3!�Z����G�"Ze�H�8�ch9p��J�ݓ�O�°�+{�����aX_w�����aX^������aX{�ߝÌ+
°���߅�k4fk�W4naXV��}�nO��3c
������8°�+�o��8°�+���q�aXV��}�f���t��k[�V�a{��[�V�a��~w0����%��Yc�`��)$X0a),�"I# (JP0b���)���0d��������?0��߸naXV�����nOo!y�^C������6ci�|�V�a��~w0�+
þ�naXV��}�naXT?��3���:|:S�:S�����9\8P�w0�+
þ��naXV��}�naXV���naXV����y��ҝ)ҝ=���m�v��u�l0v�v����\���s��m�D[�&N���O]rL�f��+a�fy��ҝ)ҝ/����0�+
�����0�+
�����aXV�}�p�8°�+�t�oMY���U|���N��N�����0�+
�����aXV�}�p�8°�+����8°�+���#XY�,�-WΟ��N����w�p�
°�;������aX_w�����aX^������aXx�P���34����^B������V�a}�{[�V�a{��[�VI�@� �A�]0���w0�+
���W~��]�c��<���N��N������V�O� �������+
°�����Ì+
°���V�a��{1�"�6�^\�Ay�-�n��K��Ʈ�j�s�ԊLY��D�յ���Y�naXV���naXV�����8°�+���q�aXV����q�aXV����u��T��K�u�naXV���z�aXV�}�p�8°�+����8°�+�{��8°�+�;�<�֮��Zu���V�a�{�70�+
�����0�+
�����0�+
��׽w0�+
���s�-ӫ�ZևZnh�8°�+����8°�+�{��8°�+��z�aXT?� G{����q�aXV�|ۿ�N��X:�Zַ0�+
�����0�+
��k޻�V�a�{�70�+
�����0�+
á�0�@�RH(@	#$`� HFFA���YnhQ�rHs�lTd7q�3�a�7X�!.쭘���Aݥ�%3Gu�7Y�N�B��5䂃 kSb�BV���asWAI����u�Y�iT�Ai`�Y���:e���ں�l��6����h�Ν	��i��Z���\% n�H��2c�ꮽjNy�l]�)�6X�'�`�Ľz��ʤ�ɦ+��*�H�3��Ӻ='c�V��L��A֦%X�+@KH�3�8����"���4�Ζ`�r��.�_�>�)ҝ)����o�>�+
þ��naXV��}�naXV���naXV���żr��ә�њs5w0�+
þ��nO�1�0�?���ٸq�aXV�����8°�+w^��8°�+Ox=�g5�[[��O�Jt�Jt�~�ٸq�aXV����q�aXV��q�aXV�}�p�
°�)ߎ���UӢ�3Y��8°�+�w��8°�+w^��8°�+���q�aXV��ٸq�aXV��ﴵѩa����t�t�Jt�Ok޻�V�a�{�70�+
���{70�+
�����0�+
�������iY��P�Ar;�:k�	��[a�3)�N�s��T�`ѦQt�Ylu���V�a�{�70�+
���{70�+
�����0�+
�����aXV��ǳ�[�Z�ZևZnh�8°�+g}��8��F��$>$!N0�
�����Ì+
°��ߝÌ+
°���W�:S������C9A�.�åaXV����q�aXV��p�
°�;�{����aX{;�f���N�������aVQX6ܾt�t�+
�����aXV�}�p�8°�+g}��8°�+�{��8°�+�x�\���Zs5w0�+
þ���aXV?���׿��p�°�+����naXV���z�aXV��O����cun�SYn��HR6mvth�K\��h����1r�[]�mK�p)�Bf��9O�>�)ҝ)����naXV���naXV���z�?���0�+o��8²S�:_O����jA�s����HV���naXV���z�aXV�}���8°�+g}��8½)ҝ>���+����A�/�>+
°�u�]Ì+
°ｿ;�VP~
�������s3����P)����h��X����¥/��k%�4�x��;��Yn�LY8��[
HK$��^��ٹwX$`�d�X��nL6iG��%�h�`1�65��4���1c o#��P,1������H���B%8��A8����-!�)�i%��b�@�B�(l�Y�PPM��
��X�h$�!�0Ab��#�Q�`nCf��2AX�@Je09�PjU����kd����0�!��C���N	J�0TBԄ���	>��	�l$��| vBO�� �<ù���p�
°�/��kp�
t�Jt��~�ޚ�b]3�:|:V�������q�aXV�����8°�+�{��8°�+w^��O�Jt�Jt��zot
����L���
°�=�{�p�
°�/}�kp�
°�=�{�p�
°�;�o��|:S�:S�����ܶQ�K4R[��D��4��3KQa��RūKESa�s�Xf�7e�t�t�Jt�K��{[�V�a��޻�V�a�{~w0�+
��׽w0�+
������`��m�|���N��N�����O�#1�0�=����p�
°�?����q�aXV����q�aXV>cp�L.�i��p�
°�;�o����aX{�����aX^������aX{�o����aXx=�=�V��C�a��;�V�a�뾻�V�a{��[�V�aｿ;�V�ĐD$�f���f�w���p�
°�/^���j���Ο��N��{�kp�
°�=���p�
°�;������aX{�ߝÌ+
°���&��f���,��I�Y�k�^aGš`�s��c8�L՛B+B�����-]naXV�����aXV�}���8°�+w��q�aXV�ﵸq�aXVt����7.�L���N���aXw�ߝÌ+
°�{��V�a{��[�V�aｿ;��������-��f���NkN���aX{��70�+
�����0�+
��{~w0�+
þ���aXV�O�ۿsZ��]iur�F���aX^������aX{�o����aXw�ߝÌ+
°�}��V�a~�{=�KsV����ַ0�+
�����aXV�}�p�8°�+w��q�aXV�ﵸq�aXV��d	���`�D�dK����	 �0d� ���,�bI�ξ��p�EX�ڕ-��$1D���E�����1�C\��}Ө�*�����G\��D�
��[h�%����t���e�.��pJ����a=Z%q[ٞt��l��a��qΈ̶�61XΨ�و�B.#���R�eK`i(J�vc��(�%��ڬ�gg9wf�v�np4eS�^�$�f�,u�\Վ����SlQ2�~�H�I��w��([�BY�)6NV*ix9�6���XPkEUp��0G$V��a4�R�����N+
þ��naXV���p�8°�+�w��B��0�+�o��8°�+������un��WZw0�+
����naXV���naXV�����aXV�}���>)ҝ)��Og�,ٚ
��aXV���naXV��{~w0��c{����aX{����å:S�:}�����4pb���q�aXV����8°�+���q�aXV�}�p�
°�/}�kp�
°�>�ݹ�\�m3B-֝Ì+
°﻿;�V�a��~w0�+
�����0�+
����]Ì+
°�Ǻ�qӚӫ�[AM���<� n�E�5u�E���l�]l�#���2�t�t�Jt�O߻�;�V�a{��[�V�a������$#��0�+{�����aX�n���5���i��w0�+
�����'y�A%�]ғ�#DC&��2ĶH[H#(�&��q�a��=��V�a����V�a�뾻�V�y�^�5�L��+�'�����~�{ٸq�aXV�}�p�
°�;�w�p�
°�/}�kp�
°�<w�a�iј7F���naXW�@�����p�
°�=�{��aXV���naXV������V�a����][��㫚70�+
ý�}w0�+
��������~aXV�������V�a�{�7)ҝ)���8���e�\���Sk�c��p�E1zRyr��e�
,++�K��m�&�!q�u��浬�8°�+�{��8°�+�׽w0�+
þ��naXV�s��naXV��}�Z�:�Ui��YsZ�8°�+����aXV�}�p�8°�+�{��8°�+���8°�+�k�ys�b�4�ni�8°�+���q�aXVg{��8³p� ����m�s��naXV�~���aXV���sإ�1�.�4�Ѹq�aXVg{��8°�+�]��8°�+����aXV�}�p�9y�^B�~�~���p�T&���aXw�����aS�￹���V�a��p�8°�+��z�aXV��{ŧ5r�.bkV��w\8���q��8�1�d:�*���ۇ��7gj�Ԙfv�Y��oΟN��N���o��8°�+���q�aXVw��q�aXV���q�aXV>c�X5ѡ�i�8°�+���q�aXVw��q�aXV���q�aXVw^��8°�+O�.��f88fj�Ì+
°��ߝÌ+
°��]Ì+
°�;�f���aXw��Ì+
²Y�������SΟ��N��}�z�aXV���{70�+
þ��naXTO�C����T��h�+H�� �2,H#&2a(�d�d$�g��]Ì+
°�{���ֲ�t���5w0�+
�����8°�+���q�aXVw^��8°�+���8°�+�@��������ez� �N�1��uS�v�rP�t��5n��.nٗL�l�d����ҝ)�a�����V�a�u�]Ì+
°�{��Ì+
°���70�+
t��zopK^�
l�:|:S�:V��q�aXV�{ٸq�aXVw�����aXw��ÌKH,<}��V���s5��o��� ���{�m �����q�aXVg}��8°�+���u��Ӭ֋�m�f���aX}�{��V�a�{�70�+
��｛�V�a�k޻�V�a������5WF:4:ַ0�+
þ��naXV���{70�+
þ׽w0�+
�����8°�+4@;��h~���JFd�Z`�P��&혓F���d-LV�@rl��j����k,���3��aF�:�[M.�3�Y�Av#v3˱�^�!�v����69׈�*%G�C�x#�!��!�Ɔ��77�*X:��B4��+,3{��F��qll�(P�\�8�t�6+I������m�� �&ݱ�o\��rέ2�E��wI�[�69f=�rs̜c��#N�&,m�
��XF� ���+X�0[�ڛ73�O�8�+��{70�+
þ׽w0�+
��{~w0�+
þ��naXV����Ɇa�(�Q�f�p�
°�;�{�p�
°�>��p�
°�;�{����aX}���p�
�����}��F����gy���V�����aXV�}�p�8°�+���naXV�s��naN��N�����[Ee[�Ο��� �����naXV�s��ٸq�aXV�{ٸq�aXV{��q�aXV�{/��tc�]i�Ѹq�aXV��ٸq�aXV�{ٸq�aXVg���8°�+���q�aXV���f�����.����\6J���7>s��&��i�Sٰ��<\��ڸ��.[a�y��ҝ)ҝ?o}��8°�+���naXV�}�p�8°�+���naXV����H�V�-`��y��ҝ)ҝ?�}��8���d���;�߸naXV�s�{70�+
ù�{70�+
��{��1Ժ�u��8°�+���q�aXVg}��8³���1�����70�+
ù����8°�+N����WL�f�h�8°�+���naXV�s��naXV���{70�+
þ��naXV������4Q�:���f���aXw=�f���aX}���p�
°�;�{����aX}���p�t�Jt�O�>�u�3]�f	)Xlh0�J�ҳv��w%���`�4V�]vħPh:�-h�
�enwΟN��N��������V�a�{�70�+
ù�{70�+
ù�{70�+
ÿ=۞���4�u����8°�+���q�aXV��ٸq�aXV�{ٸq�aXVg���8°�+ｯ�vq6A��3Ο��N���~���8°�+���8±}c$c=,DH�B�B��"���Hl�0�k��p�
°�;�{����aX~��n��iu�֭ֳp�
¿��0�����p�
°�;����Ì+
°���V�a�w��Ì+
°�y�Z[��т7Ο��N����{��V�a�{�70�+
��｛�V�a�k޻�V�a��/���(.ϟKI�Ѳ7kU��Nɕ�sմ��:�V]
�4�F,���`�+����aXV���p�
°�>��ٸq�aXV���q�aXVg���8°�+N����WL.f��naXV�s��nO�H�a�+k���aXV�s���70�+
þ��na��aX_����јf���Z\�k70�+
�������V�a�{��Ì+
°���V�a�｛�V�a�>}�m�u��Қ+���8°�+���naXV�}�p�8°�+�}��8°�rNr(�ȉZ""�)� ~�w�{��8°�+��n{Ku�t�B9sY�q�aXV���p�
°�;���p�
°�;�{�p�
°�>�{ٸq�aXV��~�z�e46�BXYYZ�-/��S�g8Q�[qG.���(n�0b���7&ә�p�
°�;���p�
°�;�{�p�
°�>�{ٸq�aXV���p�
°�?x�~�4��kV�kY�q�aXV���q�aXVg���8°�+���q�aXV���y���/!y�}��~EEqYt�5w0�+
������V�a�{�70�+
ù�{70�+
þ׽w0�+
�Ǻ>㎋�Fath��f���aXw��Ì+
°�{��Ì+
°��]Ì+
°�{��Ì+
°����/Z�50���Ѹq�aXV�wٸq�aXV���q�aXV�wٸq�aXV���p�
°�6|p�7�M�xf�é��w����{9���I��T"VY��^��I��nO�7�h.�b޷" ēO�D?pn1#�-����p4k[���L�c��:!8��DQ�E#����
Ql�Wt��F^<�v�������[�����pe�F���ӓ`��b
�"*"�X�L����p9?_֣k�%��nsqѢ����F��#���Hs�
"H���c"���1��d�b}Z2�0�@���1��M	��62$�$��#)
KH���1��AF1b��$DQP`��N�+TDD$��X#�(�����)"D��Db��KJ�h�
�5����AL��XS����G&C6F��j�ۑ-h�j8e0�G�Ie�b�hˤ5��� #]�F`���1���})�D���V1#����lQH�F0E��K���h�dDX�
},���~@��0�\��C1��� �F1�b,�b0dH���)!�U����7(�h@I̘&�$fKek4M<6R�`1��VP&�8!�P��c" !���Q��R"�FNG��6�uUUWm��*�
��K�ka�m {s�[��1��lڮ�;6s@*�������:��7X��cP��ih�-�z�k�i<��Q�1�9�{\j�c&]t��e)3G0�K���Xkv��1atT9�����s�jR�`�i[����$u�� ��v�ٗǑ�;<�{+ړ�'m�Wl8=�u7�M	l�7nP}F� �Η<�v�)j�Ys���4�%p.R��$Y�0<i{m��M�n��M=��^^�ơyqqd�*j%�	m�c�pq����y�-�A��ܝ��6����!�'q)�Ygzbե�6��¹qu(�B)J��\����%�ua��qs��6='`��7e갷�=9N1HOa9T�6�-�W&�w��9�-����nç�����v��u�([ 㰻�t۷a��.a1��\q�Vj�#Nq`�[�Zg�6m�hMO[�*�3ric�]&�Yuh75�;<�]���c)��[	�3�
�N�2d��.m;:�Q�C7JK��&��I�,#%kk
���^7C�#�#���@��Gb�R	k3�]�턅P�[l��l�p�N�mˍpLyP�ZpҔ�;�,4m3�oF�5���q�]hv�̖���Ò"<p�[��e���<�b�%��G���S[5Í�8����]�6i@ZH�m�;M.�j�#�㵀y��K�\��r��Mi��:�;R�:�^�ۮ�t� �&'4a�;C���l�0��f-��ct���k�،����(a+�V� ��〃�We^�z��[U�cqqO	�s��T;O2v�Zv�6�-<�حc��2�[���2\n�����u����,��ax�v*ցSkA.�
�0s��1\�̷6���m�L����:���e9�S�XY�8"+��#��շ�6���ܕ+�Olu��klQp��fhP#Bh¸�j�j�T�!��S\Z��%�8K�9"4�äpݵ�:���h����n]i������Bv a	�	�$�p��FH�	!p$�?I�I' %������x�}�f�����,h��Z�lA2i��̦ ��]3`�k�p+Z�P�u��X5-)���T��*�Om�lF�$<sn���q4(�)�!DekI�ՆK0�s�V2�ln,��H�B��2��oG4�8�!ȱ����a��pIR�.�d1���ywc]�{v��ѹ.��9%���M2���[,C-\��a�Z�ՈŞa�sLt;]nm+'��G�E�ɵ�!r�@^�pxj�U��t�\�s<+�Og�h�fa��*�]����۴�Dg~���/!y{��q�aXV�wٸq�aXVw����aXV��f���y������@�Z-���^A�a��}��V�a���70�+
ù��70�+
��{~w0�)ҝ>��7��uE�5��å:V�{���8°�+���8°�+����8°�+���8°/!y��ߦ�͕l�o���B�+���8°�+����8°�+���8°�+���q�aN���������.[`�y��ҝ+
��{~w0�+
��=��f���aXV����Ì+
°�{��Ì+
°��>�ك���.k��r�m���=jY����o`h27iX�����J�Q�r�a`�����ҝ)ҝ=���naXV�{���8°�+���HH?�c
°￷��aXV��}��~Ԭ�x&c2'�~צ�5�}�o����!'��FM��
�y��70�+
���~w0�+
ù��70�+
çS�ż\��SE���;�V�a��}��V�a�}�;�V�a��}��V�a�}�;�V�a|�w�0���Zp���naXV�����aXV��{׾g�G/{��q^����ZJ2dI(��%!�|�k�>廚˖��e4xemj�dm$��Ƅcf��[r�.x5�72á�c�M�3@�WT�͙�
BD�`ۏ@�9w4�-z��~�3�]�^�s�}�☛�O�9����)�qrנs����*J\o�I$G�{�)�qrס�Ad�w	��!&��u�ͫ��{���{~�L���l�[�s�����z������mz�p�2xئLJG�s������mzֽ��\��q9� ��b�v��3gOoF ��V�V�9�ģ6��Z@ZX��,by<�����>W���j�8���廚O�ن7�ɐ�x�q�Wj��y�y�E\�^�o{��|�+�=Y�*IF��J#&	Hh_Z�s�s@�^W�{l���� �!"p0mǠ}�]��y^��,��ٙ�f��33'7o�@9�2�"�I#O�9����;V����@����1��jm�����GS�X�9ke�yB�f�u���j��7@7)�b��tW-z��^��9w4�ֽ ���S�8�d�m����נ}�]����@�rנ\��\a��ɉH��˹�|�����h/�^��e�n�����f���נ{�)�|��z��������^w�"f8H<M���e4�ܯ@���h��z�k�/U�����dt�m�kGIn��V"�Ma��W{Tk����q��4�6���B�����78�9�]j�D����p�-��4u������*=U����E�"����e!��L��5�t��X$ͤ���Vμ�n���n�Z� ��UAH�C>�ێ���ɦ���
HE�*����B���Tmb\�X���m�n�i'P�Z�찢�3����찔{�^��P�,њ�[yLM,��n�Tc6BƉ�l"��D��%��>�ν�[��z���r�h�A�$$�i��nG�}�w4Wֽ�YM��+��x�[YׄP�����������+k�>_r� �-��*J\ițRH,�@�[^�����9l�=_Z��s,N$�<��cm8��ֽ �-���^�����y�;������77Zh -v)���J&X��kPeT4Y��2�L�0�#`�0�hWXf�zo{4��z���/�z�0���F�L�2g/�}���o	�Ӊ�'�6 �FH,�ĀnAy�MV��.Z��f�_�^_��� �6��*�@�}k��f���נ�k��Q��z��^�^[4���rנ}񜃬HI����ۏ@/-����
�k�8���/RጎA��Iڗ������9����N��5Ԃ�|�:R{Ep��m�&�궽�Z�.r� ��h\�)q��#��r=��h\�zyl�=Vנ���JBa��@��+��l����<��I�� d���� �a>����m^~���^��u�$����q������y�M���@���.nDǎy1��&�궽�e4.Z�����e,ո狭�=���o=�@�D�ň��̂P)�+G`���V�+8��ڳ�S�m��8�k�s�h+k�~\�ő�(̙!�qs��ؐs��=Vנ{���?��	9�x'#�>���=Vנ{l����W�Z�xE ���q9�mz��h\�z<�<�c���{r���G�Ń���)�qs���%4U��_{���<�ݭ�b�2��0��y���i��i�+�!h1.��\�3`T�8�d��R�$��Uo^��rS@�[_��3�w������w�#�L���@�9)�z��@��M���@�0�F�M'��1���z��@��M���@�9w4긝lR&c���jG�{l����W�s������ߗ+B�PS2E�qs���.�궽��ZA[��� ҃Nic�EÎ6�&,\�"�L%����.#kB�8ѠY*ݳ�Z�q;�$�;�2�`�����<5�f��u��݁5`�!a�[8�V�>�1ڋY��s=�������:�U�ăv���]��^.�g�Մ�z��s͗-�I�u���;Xui4��X�Sf������o
;s䝗^V�c/�CL�J鞄�gI4�[1�)�M�+��6�x[n����ӗ���M����)�sq@��<��B<�	������=Vנ{]���g��
�z���]xE2''�h+k�=�ՠqrנs���Ϩ�Ѩ�6�sG�{]�@��@�9w4�����U,r	��8�k�9�]��mz�ڴ��\�%$ƞ'2bR=����>Vנ{]�@��@������I"��Lm���a��t�[s�xzB��,�@QH��9�ua*(��Lq�&h+k�=�ՠqrנs���N.*�r(2)��ԏA�s���@2���H	 ~���<Ǟf���@��h+k�~\�
4!Ld��@��@�9)�|��@-����� REO�z�31w�zh]�^�[�4.Z���W�R	�G���h�ՠUy^�W-z���;�fb��iv&�qe�8QWxng8�g�Jc����*5���\�M���<E(��\�QOm��߿o-�\�z�S@�;V�}NeNLX�8�a0N=�r��)�_��@���e�5��`�)�q�۹���w�n���3�>����t��W�E���I��J,���n�.�G���!��#�3DM�kH�fddMmh���0�
�A�Q��NFҕ���S4kN�f�	b@`�C��g�f&`��;��Y$D�X�* ��DX���"�`��(VeQH)a�J�0P��F""��h��4��A�
�1RY��`r#0��� �x��;j�kLb����J!lԆ��l�`�vQ�	'�$� `Bj�h�?�$�l�� 5@�>$'��I2�C�����w�W�߻�W���.�&LQ�&h�j�m�\�z��h>\��F�(��r- ��4
���m���ڴ����]�v��eݠ�պ�:������A"�(���k�v�頤ų�s�m�r��n��v��g��;����1�}bX��G�z����g�u��@;������@/8�a	�#�����mzm�h\�z����(+�"LiI �r= ��6��ﻛW��vm}��
Ќ��$��2Q$,�(I%@�2>t�k9��6���O\ֵ��Ӫ��8���W�w<��������z��s�������C
3in��*Q4�1��3[j����k���
��B0�*J9�d�2bN?@����궽 ��4.r�ۅ*5��ɓr9����� Z����ڽ��j����HIj��#L�"!��w��-;	$}���j�����~��V�t�	O�)�8�k�/��hWj�[\�>���u�d�c�`	������h-�hrנp3qy��'~�=���<l�R�qh�f ��V��eɕ�\
�,[٥ֲTBb�v��C�s��h�ۤ�����u1�v	�{��luaGk�f����nkUj4��iH��C֙�Ejr�8��I�]\;.��PX	1,b�Yj`*�hZ���p����[�{
8+��'��ȘZ����}�i�sSct�4�ɬ{�à���ZT�����'�t��=1�L�P�V�p֤�^����v����V��籩9�n1�U.m�CfxzNg �}�@�ɠqs���w4�������I�H�+l�-z����mz�eNH�c���`��@��@�[��|��@�ɪ�����X�EѢ��m����{����z�+�&���W�{p�CA������f�궽��ɠqs���]�����FG&<	2	!�Wa���x�FqeΎ���vb��ً
���h�&�G���ԏ@⼲h\�z��OHIʿ���گ����Ӫj�tWS35�m_��w7Ї��rBI����ٵ~�hW�M߱�bY$��I�'#�/ܻ��ڴ+�&���W��c�^b�e�%��=�ӧK�{��=]��@��+�=����P�����9���
��h\���)�|������t�i�V�d��˄�
�a	��.�j�(%��8{^ N�����On�uk�ӹ��Da0RI�qrנ{l����l��1\ׂ�)�dĜz���$��}�f�����m_��w7�HO>��4�LM�!�|�޽����ޓ��AU��� ���YDU�T" ȓ�@'�	����=u��@�y:h9�ǂ�<dDȆ�z�1u���@�޽�n�{m���*B�$��O�M���@�۹�U��@��&��g+�k�5���;��&��{&�%�0^jPX�C�	�6�f���$�nܼ���$�$����w4
���[d�*�+��uyC����U��{�y�g�����4�z�m������;N�wRC�Ҏ4�R=���\�z��h}k���WcƤ�`��C�f.�z����h=�����?�d����	b�RT#H�L��o��9�m_��^��ɏ�2bN=�˹�U��@��ɠU�W�{��K|pm�&
0Ȑ/��I�2k/o;�ۦٶ��`X<���t�	��+&HОLQ�!�U��@��ɠU�^��䦁���B�b���$�*��hrנ{y)��� ���!d�K���nI�U�^��䦝���<�H�{٠uv�M߱�,iG	2c� MǠ{l��}m�V�4;���*�z������� ���$Zyl�;�g����O@���=�S@�0�@��$	��7Z�sFR㬦��� �r���nhSqv�6��Mu%ݠG�R�!Ɔ����L�:݇�����ۨ� =S���bh��VO.�ĥ�\�/��,À��(�E�3hQ�,z:ݎv�M�M�lr�=�mn�"���M�)l�_e��P�\�X�b�	[��͖����:��h����fbł�pr	n��p%;hpV�)�H�Q����'N���$�xx��S��Z�N�qk�u�i7�Q:�Tu��v���<F;utL�HӄC���1H�����@����e?g�g�z����@9��vLF6)��'$�*�{��w����{נUm�@�9��JdŊb�1)��\��[d�*�@��X\��,O"#���*�@��ɠU�^�������D��1I4
��hrנ{l��^[4V�����F�<��%�Fh%f�b�a���
��0Wjl��#�sib��ֈM�&�W-z�����h^Y4~��?:�Eb�x�;�>~�}�gt����@��4�\�8�k��癞x�w�����	�N
C@9��h��h\���]��ԩ�I84�d$�y\�8�k�=�����<�.w���v��1�N8���s@��@���h�٠�w���3��w7��F�n����(c%���^�Ju���\�H�&G�sJ��]�`��m>���^[4�\�z��TۜX\��$<��73@9�8�s�h\���w4UЍb�1I6��������{�X�22A$"0�@�6D5����j��{� ���!dq	�Bc���Z�m���f�s�<�3�o\�9��;J8�y<q��Jh���v�������Z�
�>�qc#�c��P0���2:�.+.z�B�Cj����e%m�31��5Q�dmE����^[4�W4
�k�=���/ŭ=�G1�55$�y\�*�@���h�}�:KC���}t�st�π{w�@���h�@-�s@�8����1b��LJG�{yw4�٠�m}� �$>	�s=�ڿx|���BǑ���h�@-�s@����˹�}^��b�d�b�����b�zp�f�Ы���չݰ�΍	s%<sA�l�J5�jdx�$�y\�*�@���w333�o{4�/RH� �9�Ln9�U�^��䦀^[4
��h|;H�RG&
d�QǠ{l��^[4�\�*�@-�UĲ&�0����W-zV�4
�k�=�S@���l��3j!�#�-vǠU�^��\����=��)���?Z��*�a�,�,��	� ���7��0��D+s3�s5E�E)�7bZ2 ��D0]��`�R,Tld��و͎Ĳ9M��#��H�/�+�AG���������P��0��`���;�F͌F��%��4�[������,~�}��x��G7=�s�>�Z�}[���#F��D�5j
����A�`���1`�"��,TQ���衩�DM�\��$P$B(�PX���1�X1`��@�a�&�2(	�lԒ���P��@pB�Cd�A�"FvE.He����c�dX@-�QPR"�R`̀&# b(�H)�"�8l��
.�����))Fƚ�pdH��LtJʍP�6DEPP�z2���C�n$g>��d�b(E�u 2�`�H�(#�
!*""1��I&��Dn��# �ր�,dFؖM8A]G���$C�B����>�}UUUZ�
�ڪ�����I���HB��4+�+�+k�F����y�\�ۍu��,�����[ ���%F.�ݑ�	j7juAL�-qY@�m��ե��gr��tEtq������+�1���&y�答��pw <�8��˴��s�/(�[.�!�I���t�묽䵜�'VY�=v:�6Y��tG����Xbm{>�V�Cb���,nΰvt�Bq��s�gx��5��r�a�c��m�.�1��!t1H�-��M�9,�&kB%Ֆ[X-URM��.n6����_7�� ��oj�G!�D��.ð�t��il�f�l�,mC��0c�*69+�����5Ѽ��8]f���nݪb0Ԫ`�-�;F�.-jaqȺ6�y��[N��5�YM	�԰�m��Bq	w�����s����#�Ki�a%��\e��d�X����vCr��W��ֶWeb�X���:&%KR�Ps�ns�ۯa���&tSFg�aKl:o`Z\�-�q>�rB�����n#n:��i��k6P�;0IU,Y�J��m0�Va�j�k�4`�n�Wn�9)v�a�D�I
r#��6��!��h��M�P�wcTgF���<�;�!�L��#	�z�IDn�0`m�������n�iP��dUq��9ۂ���8��m�W��r�V{sl�@7*t�Y��feخ\z��oK�ÄA.v˗��n#!�NH�Wku���7�{85�`���]��k�(XR���n�km�W����u飵!��Tp�[�B�I�wTn{oMGQ���9�`�U�b�\m�Ʀ+e�
��]76]N�C	�g Z6̓f���	"Nn{oV͢�s��[�Y�^;S��J�%v�ݲf�iG�zX����sȯ:��7����lݶ˘b~�0������S6˔e�b����q�3tN�,u�%�x ��Ⳑ�Ѓu��BE;��-�Y�OӢp=jwF�a�s"tG�f-��mZ�8P����p��`���NOd�Ӱ ~��BCd�!� �'ВD�|@:�I'B@��k���P�Փd�S�n�,��A���'<�c.�N4[t�:�rD�m�՝�wl��B ��5Q���&*�ݦ��Þ�!�`��JS8�s!\R�O3�.�m�I������\6���Lki^�7.K����']<<�:�v���v�퓎3����5�F��}�'.��0{\�d�7��5��h����P�=��S�����n`�u����C��_M4q0(k�� `�X��}O	��M���"Re*�L�2ј6aF۠�c�`�n2�+�v����z����Z�]���p�ې<&LJG�{m��*�@�v��U�^��<H����Y��`��dq�������ށW-z���՗�RQ�cS#�)&�k�=�Z����yl���I"8��brG�U�^�~�s@/-�+�@��o��\aniWM�
ݗe�Fc�dӺ������Q��y�aJ�bq5\^q��]� ��h��=�Z��WF�s	��Nf�^[4�a�H+ �CRO� ���;�fի���˹��<�#���'�F�1Ƣ��뽏@����˹�U�^�{�Ù`���I�&$�z\���]��Z�;�g��+�{�zU��Ɋb�1)�~���*�@�vǠU�^���+ha�7�x(�h8]���B�a��k����4�9����G,�Q�%��1��<��s4
�k�9]��r���33�w���>]Ԕi���]k6�{��~��k��{6��{�6�yl����^��A�p��=W׾�m^w�ٴ�?,�a,)$0$��BH} p ��o�����c�>�v�4��LI��QǠ{m���f�k�=�Z�yO#M��	��9�yl�-vǠU�^��o���o�7LJ57:��b�lؖ4�SKG\\9#.���\��	��pq���&�k�=�r��e4�l�h�I��Y&H	I�W9^��~�h�c�9N*��6�LSɉ8�m����@��&�W9^��ʲ��r0O2H�4
���-�hs��,��'��L�̞��4URQ�cS#��rڦ�W9^��_Z�W-P���W:@�,��-��Z��ڻ�t9���N��Gcyᣖ�]c-4aq�|������e4
������}��E#���H�m���癞x�����{޹�U�W�[Ȫym4����*�נ����1.�z����@�̴���Q(���@-���r��e4
����܉5I�)�*�+�=�S@��^�[k���N���o�l*[ղˣ�����箄�����d�f����c"0��n�����Ŏ5�H�{p�:�ᶙ�*�i0TbbY�2�.yK75{u��k�� ޥu�X��&M��ۆ�ʠ��g�s��4#i�cHi�ͲnC*��,pDIs!��|�i}�i�m�Kzڂ�5�c4�,s&��KXuȔ!�lX⫀\�����Lc(�v*�V��l��t�wNd�d��B��#�b"жӴ0"㮺]q�U��f?	��L	���+�mx�@I�b��' ���h}k�ms@���@��X\5� x�2H�4�l��y�fbA{ީ�u[נ{l��338�*5�(�1�����{ީ�U�W�{l��_����*B� N`�NE4
���m����C�ffy�^��h���P�,m��rG�{l��_���j�\���ˮ6Q�����s�v��ԾwW��i�e������Ƅ��ɮw �[��b��b�٠���U�^��������F���߻ޏ���=�skӗ^��䦁W-z~��"MG�Rd�%"�\���)�s�<K���@/oT�9C�\�6�@�Lx��@��S@��� ��S@���ۜXP�G�	�I$4
�k�;�y��;��V���S@���E�Lm��I���h.�a�q�΋�bʹ�^�C\fe�q�����n= ��Y�U�W�r�S���w�@8s�X,�"x��&�I4
���[)�U��@9r٠}�����y<$���S@��sn�Pdj��F@"F2_<���2y�d�.m�\�z劰q%�����R_Z��-�\�z����w���w�l��q��JG��l�*�+�9l��Wֽ��&�ٖ�Ys�K��q��$ŤR�-�� �Vl��[l'7l�Kh[��M�r���h}k�y��/f�zTgscM�a0��'���M�y�y�$us�zޝ��*�+�9r�(-��bxFI��Wֽ ��hs���S@�Qg,X
a�DH�7��HK}������}�W��]v�"2����M����}�mW����ɘ���$�$�\���S@��� ��9�KQ�",I�Lib*�J�&�¬��AC�s����㑏`�] G%ۖ�ą ��a#�@�䦁W-zil�*�@��\y"�X���W-zil�*�@岛��<�H����8�dX4�z��vhrנ}l��W-z~��"@�"nd�)�*�@��M�Z�;��y�]�z�zTgt����ǉH�m��*�@-���Z����g�b�D�I!�x��1��Vk5kP���Զ,(����ZB�q��FY�!m52E)(�XT]�M�D̶��f�B�XT�*eōшSJ)�X�\�ΰ����c �9��p9��&�kc��.�ʦ�vɸ����ϣPZ�� \���M<���Gu6rs�u�.�W��)�^:ɞ��}�8���Ņ�-�z�a�,k�m�m��0l�$�vr�Ѻ��t��w<���1+�ڌ+4����{`LJ)��]��u�P�]$=�.���ꎎ���,L&8��]�����U�W�{l����X�Jb����n= ��4
���m��*�נZ�Y3�pI�#�\�z��h}k�ms@��v�@XHbra��=�e4�l�^U4
����E^1�������@9yT�*�+�/ܔ�.ecb����I�&���I���a5��N.b�ut�6��s;����J�5�RO@-��q}��Ϲ2 s�rh�U`�����SE�����$�C� p�F���5M �٠ڦ��qt�6&<��'�~��~�h���U�W�{r�,Kr<X���$�~�h���U�W�_�����R`��p$pnM ���r��e4�l�=Xe㸣�<�#�� �9�v�s�f�/Q`{t�$A��pMm��9�9����	cNE4
���m����@9yT�=����	NL0RG�{y)��� ��S@���W��@�"� �4�Y���if|y�
��:v�nBT�D,��.�Ś�c`�����C����JoZ�׽�lc�f����Fvt�D@c+PEI�$s[`V���w�[��uÎ��y���5��G�� N~P�u��S��E��E�@p���R""b*�����sZ��o�w���A1ĩl�R�����#��$è?���(�1(6Y��c�D	5���1Q�NA)���~���XF0F"F$D" h6��c	ڠ8,K$d�(��^�����MЁ�\X"���-�-�W��"�K�G
|3g�p�`�_��N�@}>���Dwh�F(�����j	mN��Ab��,H�ԕa��$�HM�"�&���H�o�"�]�S�Y�u�Nd̄1��
��,���n�l�$4�~�`g	�Vh�
�s� jh@AMYbVIM�Ud��5�*p�C�L �$� �$��O�~$7$0�M2�!}�P�O�!:I$� �@�!�@'��y����ܔ�/Z���'�8��^U4
�+�/ܔ����g�w��@>�w�dN8����S@����M ��h��h��reJb�6ԉ��&*�c�J.��m��Z+�n�z$yK��:l�2B4�1Ly2bN=��M ��h/{�n�9W���m_���ݚʴ�c�I ��h��h^W�_�)�|����",#�rh��h^W�_�)��� Ͼ�!c���Kn)�Uy^��䦀[�4&g�'����$� |BH�}��m_~�ކ)���`��@��S@-��ʦ�U�z|�3οg{�C�s��s	�vE��9��y��ok�u=I#n#���jUc��1�vseR���{4��M����fg�>�4ӽkd���1�&�[������<H����>�4�Y��-�##rD8��h^W�{y)��� ����
��NbSL���@��S@-�o+�W���9RŬ�`���$�o,�yT�*��@���x��N����~V�.2L�\��5R�Q�"31rՆ�m�e�:Q�����`-�4�k��ͺ��$fLJ6ScK��U1�ԥ~��o��	q��rV����ؗ1����h�t�W��.IW=��U� }�6�ɨnSu���9�::��vN������%�ʭ.]&B%-P�(4��T���[ly퀶�J ��-3n^���v���I�C[k�u�܉:��?n���Gޭ���yM	�8 px�áh����0u�vd Q�W8B�\1���� 2"G�����\�zג�~�h}�*Bǌ��pKx��*�+�-䦀_��nr���y�$}�}�b��6�`��@�l��� �9f�U�z�k�*#27$Y�Hh��@-�f�U�z�S@�-kd'�5��&�[�����l��[�4�^��$6�Rr���x:��]T�d�!�uQմ�˳VP�6kP3��Z(B̿ ���נ[�M ��h��4��Z�Z5���4[�ͫ�����~�~�H��I�	���[޶�Οw[B���\9RŬ�<X�d�I �[4��\�z���>TY�u%�Q87&�[��@���@���~�h}��ŏ$X�8i�@���@��h�٠�@���g9ߣÿ�lgVkjm�-�A�Ha,h��0����í��Y���2�J��i�)#�����[�4ܶh^W�}Ƹ�3#rE��) ��h�l�*���)�{rֶB'<q�b��nr��k�s�y�y��a�R@�H?I
BHs��5�j���h���"na��&�U���S@-�h)�4��Z�Sɋ&LJG�r�S@�瘻{��z^��Z��qTLX�mI������٦nPp��Yu��܁��v�:�u�����%�2�cɒI$4�٠�,�*�@�����9��y15�rh��4
�k�-䦀^[4��X��ȱ�cO�\���S@/-�nr�ܾ߱Fa� ۘ�=�Jh�@-�Y��,�0�A	�,b Qdb�E ,��(�(�$� �$$�����=�\yq)��8��E!��4��Vנ[�M�����}/O���[l�&��^�O;��;�����V�P�B;UF�F�g/�}���Vנ[�N�y������,Y ��,rh^W�r�S@-��گ�>����Ǻ[�wZ�Fɉ8��:h��@9s�h^W�r�ʖ-q3�&H��yf�r�,�*��@�䦁�ʳ���&6�pnM ��\�������m^��H�1�!�.fw4�ѫ���WPnW� �+:��6bU�1B9eU�M#ѴV�+z@��Gh�a'��Q\��ìr�X�n��7�T4ݹ�wY7E�ŷ��B@�Ȋ�I��(.�1fͥ�d&ZCM�6��lA�AD]���s��3��qm�.��؛�1Ժ�;�'��ڭ����F٪B����Z��&���Y�T":+�LUR֩31�L�:��$����i4k4�jc�xY1{\΄fv�my95�E/-�)�tt� d4rэ!3"M��������m�@9x��=�;��� b���=�m�@-�f�U����\Jd#�,'�Hh�� ���Vנ}y)�{rֶd�#RL�!�&�r�@����%4�f�{N!X�Cn�$�*����M �٠��h�e3R��--�.�S�q��U�\L[a��.�<��Y�V�T���`mX�f�`.��gM �٠��h[^��Ö�|͘,ы�O ?~���uモ�.�P(	HP� ���<�9n��|��@��S@�eY�TKȆD8�ܚ�ʦ�W-z���\����(�9�8i���W-z���\����h����L�$�2`���%4
�k�^W4
�k�/8B���d񰘉�J-�MfP�7i5+��Ka��b�:�W)�Y1uo�=bS!q�9�Z��U4
�k�=���/ŭ=$�$�����^h[^�y�M�k�xq
Ʀ��&I�Umzג�o���y�0���*�^�_�Y�}��*jO&Ly2bN=��M������W��\⠳\Y0X�c�I����h^W�^rS@��y�wO���]���`J��Տk�$��3�w&NӺYM[��J�k\�4�X�g���{N��r��_Z���H��4�&�W9^�y�M��zo4���dI,Q� �G�^rS@��^�[���r�ߚ�ˉL�j@���4
����{�����ͮ�OŲK��F�"a�����8�B`�bb� ��7��:�_ߞ�.mִi�֋�j8��h^W�^rS@�����C~!��8�.�Ie��Ü.��V�	M����:�\�Ife��(��*أ�bMI�Umz�%4
�����/j��9��]5	FLS	������瘑�����]�Vנ}s���qdHO$�C@�������k�>���=YPr�XD����z���j��:�޽��M�Z��}̠�Nf�A�Ԛ\������y���{4��߯�ڿ� 	$��� I?�� 	$�� $�X@I'�B I?� $���@I'���O��@`0�I�@bI��D$��IBH�H
I�!$�I���$��$!$BH��� $�� �I�! 	$�� $�X@I' @I'� $��@I'� $��@I'� $�� $�� $����e5�y6��}��?���u������� �      � z@H	1�JQ�*��@֢j�Vf��bj�V j�LZUMh1 6 ` �2 3 `$@$@n�F (M4���D�@��  Lښ�T�M@ �&&�da�i�L� `�  OǪ�52*      RPL�	�O"Ch�@m5MB�H�i�I�驠221M�ӫ^ʻ,�*|;	���H���E�)�����%K�F+$�@A)��0�Cl	c �H,�C��ꟿ�������bh�8~�?���!ʤ�����$������0F��^�

���/��Yg�*2�!B(�(�R�QVaU�e����{���J
�ieJ�+s{���SMf��k"UkZk��%��0�ʼ��m���)�#dJ`U�`��%��2 ��Ē��L��Vh�h%55(� ���R�U.��]���I0�hK�@�ouxUP1��5p�w�P0�j��*��$r0�2�����\�Z�B�D@
�K/�^@���IWx�K�aq�$D�Xي��i`���W�$�*	@�	LR�&�ֈ�	R,"T�1���B�w��(���?�,,�w���w�ӻ�+���޻�����                             �=                                                                             �@                                                                            �=               -cK�6i�.'���]��/�[oz����"in�@X�v�^:��ם�m5�5�۬\K$a�x���9z�f�A�6�.�m��6�^�ܶ��@�u��.���N� �@�mnl�#�P�u\[F���m�d�[�m��^�3mJ 8%�����4[n��i{M��cm:`�[I��f6�n���'kh6�c��Á&�#]�k[l�cdև[@s�� 5���m�'mp�h��q�I�c��Y���$� �Ӥ�.��l �[f�$�j�f�M�^��ޡ �������n�ٷe(��j�n 8/Z[�A��۰i�+v$�t�:ie�sI�$bKk��e�.ۋkn�I�%�mk�ȢI�B�ImH�ηkf�.tۋ�k�_,���~��$iK��H�cZ��~���%ɦ ������] ��ɲD⤕1�(j#!%0�,�z0>�@A/�,1���	RB'��Ϗ�    m�              6�              m� �jU�k�v���&���dƐ5V�-��wj��eЭ�sIv����,��ʽ,ͻi6�m���e�mv����M5һiӚv��:XMx��+�r������ �@    m�  m������+^�%�5��P����uf�m�����~��~Z��7���_}���$���雹=�� -`$#�����UWʳ/��mn�e��<@ 
(�
*�{���o��7R�&=��{��< x���=u=6���\�S_}���Ͼ�ڽ����=�� Y�07~^>��䘌���=u����c�          -9�v�gO
�����i��.0���$���!�{���o��7s�L�ϹU]� u�b�'���=u=6�rI���!�{��@ �AF+�O_W�n�T�����#.w�z�~   U�1n�e��Cj�=�F�y�/L���@ ��YbX�^I���{箧���I6[yڬ�M            N����/��V:��6��P'2J���y$���雹�&n�罈��� W����C�S�kw$�-��n��{ލ�� ��3ś��&n�罋�"��B����}�m��|C��m���������S�| w�`����}�w��z6��3w��}�s�� ���A�-����]O�rI���!맫���� ��     6�,kkU��Kv�B˒J s�i+w�^������)������|��� `+A���e��Cj�=�F�T���J��r����  Z�Łk:��|WX�˅��]�;���q����4�al���:8Ì��V{3330��2V^
f�����q�N$�z�i4������� i3]�alĶw�kٙ���Ve�b��3i���,����}�����e��Vh�S4����Ì�q�}z���    �� :�$t�E��n���5����0%$c.��w��i����p��ү�L-����|�3i����u��W�<� f�$���u���f�
��[;��3�ė�U��[�w�\3�����;���@ ����fSf�J1��}���N'X?}�Y��XBY��o�G�ڇR����Ӭ�:�Y�t_>��  ]�
�{��HgY���#��sn����'u�!���%u�J��I��D�i52CK���}�/��Wr�u˛�  �HX�*�^f�m4��"c>����נHf7! ��l�Rj�;Lg���B���~P!A��*�PT1�z>>�_p                               ?�       ѥ��\k��rT��%]�T�f��;q$�o6�j�ŗ�g�-�u��R^K;"Z6qi/B	[���PjR�q6t��i%�R�Z�U|w���Ӟ�=�      �����v�v�K&�$�o}��נ32���4����������%�K�=�fӬ���f�L-��w�G��{�i��� E�3LK�Y��y���q�	��L��L-������i�}��v�'i�����ҝq[=fӌz�3I��{�ᣈ/i��+/�t����]�v�ʿ  �J�2�i4������-*�t�ىl�o���m8���z�3i��&����� ��++k����]}�n�r������q�N$���i4�������i�_��       5�6rmk�撍z��͚� %����Ke{���3i��z��g��p��e��Z�P�i-��{ٙ����e�Y���q%��sI��g}Xm��iW˦�Ke{|�3i��}y�fffc�幙�x3i�Ͼ��8Ì���Zj�A�c;����ė�U�&�+���@ .�%�kmv�]�+�^Y|-������fӌz�3I��{��z�s��<ӯ�|�r�])/�g��[;��3��? A3���l-��}X|O;�y�]�Y�i�v�_~��       M�\Yi���wm$j��v�ՙYX�y���q��^�i4���{�4q�i�Vh�S4����Ì�q��� e�]��ͺ��+�OL)�)�ү�L-������fӌ{X�I��W�<� b/+k����]IY��L�[;��3���<�r�8ts�;yW:�al�s���m���� �
���J��J����\fӌ{X�I��{�ᣌ8�z���m�+/�t���$��Av%���ͧ_�W4�al�{Ն�m��|�`��Ҿd�}������          ���I���-崳����L0k2�/2��f�L-����Gq���kMB���w��g�/ޫ�M0�o�  �ai,���|WX��ꉛr����q�N0{�b�f�[=�{��O;��N�g�TeY�u����<�{�8�'_�W4�al�{Ն�m�����J�]+�� W�B ���>��f�L-����Gq���f���ͺW�{Ю�;u��u��  Q`a��usi�o�F����a�u8�J�]3I��c+9�ގ3i���/﹋8�g������o���       ,��4�:رd����@ H�gkxh�6�f'�Y���ٴ�{����1��Uͦٴ�s^�a�q8�O_�y�w� �bY|wE���=趻|w]f%{ױ�M3i��{�4q�N3ެ�gҾ;����  Q@P��������m6ͦ3���3��bVz�t_6�a��mv��|.��  ��ܼʼ��6�����G��1=�ޚ�KO���>��u�N%����si�;��<N� ]��B��6�|w]�Xz�Lf�Y�v�q�N3���ͦ�;���N��o����+�O���                                         sM�ե�K��XӷJ:i%N�uY�kt�F�#��&�.i�M�I�dj�ɖKڮ�I۵i�֝�FT���l���Y#��+�Ŷ�-��Y������;�����ww�������      �R�յm6I�*�m�V�M�+��%���(�;�Θu�N3�}W6�f��{Շ��1+;t�&3I�;��  ^`,.�-���o��H���q�3��W����3i�b}�oMM��wE�I�+���v�]KQ�$�^�wW6�f�Q�w}Xu�B	��4��]3I��c+;�^�3i�bW޽��i�/�^p �@RH����o�׽[�Sil�c=�pÌ�q������o�|�Ʌv�ۮ��{4  �"�m1����G��1+޽��i�Le{�ᣌ�q���oMM��T�i�}|z��       ��iy��Ydi�Mc��}��O@vh�u���>'}������m�Lg5�Vgbgj�����E���k��u��|�D� �����i�Le{�ᣌ�q���fʛKf��{�g��g�W6�f�]�  ���%�]�;���<���C4���w����q���^�m4ͦ2�������v�]  x`�.Ċ�4�m1���a�q8�f{�si�m1�׽Xq�N3��L�c4���;������3/-̼�fӌįz�3i�m1�����3i�b{՛*m-�Lg��q���x���wo[� 6�     -9eB/�7T�ݧY�I� 9Z���6��kެ8�'�Y�i1�Leg9���m8�J��c6�f���v$��V�o����LgҾ;1���a�q8�fw�si�m1�׽Xq���s�����KDf������������{f��}[Ȩ��b23�hJ)(��*������A�#	,jDF25R�#�(5TD�(1�Tc��*�D �##EȒ#H�%�,�Q)@c$h�@0	�~H@���{�����w�t�� E�-aOZ�鍵�Lm�^���]�֔�  ,�V �S֮H��RA�Ƥ���t���]��     6� d��S-�xض�&U�vL�D$&��z����������{�=j���֮H��W=� ��w���IO9ʪk��6�I1��zf����� x�����:z��=�jH:xԐt�� ٘���X���cmZ��5Z�|���'k��s� � H
S֤���vA�ƺI��	1��d�          �U�H�[�,����7K`;b�Xƭ{�=j䎞�rG_r�\�:�}�ç�(�� �����5�Lm��cmZ��5Z�|����� 
�b��OZ�#��IO�t�cm_�  ���%�Z�=�j���=j磧�\��֗�� *�$SƤ���t�k���V�3M^��
���"]B�B~��y�                                      �e�N��v�[{v׵�Ӕ[�K-��v���]-��Dt����6�.��k�[wf�%�K5�.�\�/kn��IinܚSt鳚91���ӷ����Ϟ��[=       \��k�n���֥�4i;S :UX����{�OZ�#��IO�����Ud߾  ��(�1gw���7��}�k5m��@�cW�}�P'l	��Ͻ��333�[��@�`M�'��@�`K`N0&0'�}��8����`L`N�� N0'�	�	�{���	��cv��3333��2�.�q�4��`L`J�}Ym�4��`L`J���P'l	�������N0&��	�	��k��N0%�'�������0¬����	���cw_}Yq�8��`L`N��V@�`N0'��V@�`M0&�����6��`M����=���{       �Yj�i1�Yy�,/Y�`hً���m�8������p�	��q�1�>��p�	���c}����	l	����d	��q�1�>�}�����31r۫�@�`M�'��V�!$�4�Z�W􎞵H��W=� � �� ��]=1����g[V�3MO��  .�/�c�#��\��֤���IO�Q� ]ш�K1cֺI��k�4�i�4�s�t����        ۴��]��Is]�E�&�,�  ��*S֤���IO�鍵�Lm�͚  ^^�ծ���+��k/ǝ=j䎿�u���O��  ��Aff ��W��6�I1��@�1��������KB���~�j���5<�� V,H,����:zԐt� ��]=1��Ā H�,X��^����9\��ó��#��_�:z��          ��'K��m��:e���l ��f^,E<jH:x�OLm��cmZ��5<� �*���XƮH�v�H��RA�Ƥ���_�  (I,IcֺI��k�4�j�~ϹOYH��K�| V,�F"��$<jH:x�OLm�*�K����g�  �B%�j�fi���:z��=jH:x���       i��[n7]�E���˻*�  �(G"�5��k��6կL�U��4ԧO  ^����\���q� ��RA�ƺI��<�  �(,�,zծ��U��4ͻ��\��֮{` @�� ��]$���鍵k�4���� �і,cW$t���:zԐt�{ٳu��#���e�5AR�у(:kf�L�21ČA��t����t�y�����         ?(=                             h�u�z�$��ͯ��tkb��j�";\��]��uś�v�\�[n���]	ڋs���I�v�h�N�5Y�f��x]f]aT�]��F��iBN����>=|{        �vMcY+����vU�ܘ �2B]������~���V�3MV���U�y�ֻ�� H�P���${o��IO�&6�OLm�M�  fV�կL�W��I;]����Ξ�${o^R  ]Ҡ�3SƺI���Lm�]���U,���S��  ���"��rGOZ�=��IO�&6�}          6�*�b4�4�n�wE�H��� �+�,zծ��U���U�y�֮H��K�@ ���X� ��9�y�Lm��cmZ��5<� ����1�\��֮H��9Ƥ�m�RA�ƯĀ %�j�,z�I1�����f��vg���W����GOZ_C� 
�e��1��#�xԑ�k���]$���r�u��OF�          -�Vks�[*�T���:o]�y}zz ��hծ��U��t���:zԑ�j�  QFXs[ƺI�j��k����]���O٦�:x �!"��rGOZ�=�������+�����U_r��������۷1�}1���` `X0ǭZ��5Z~�5\��=|�+�:z��l  �,Ł�-SL�=��x�k���V�3MO�x         l��zL�jQ-��)u��;�  ��5rGOZ�s>���w��{o�=��O(� .�E�icֺzc��v�UΖ{sMV���U�y�ֻ�� H�P���${o�=��U\�U;��[mt����h y`abXƭzf����\���|�r��I5�Ɨ�� t�e�E�k��m���jצi��}�j�^         m�.%T�mm�,4Ҫ���ם�s�� U��`�E=j䎞�:o$���{ލ�� �XQ�,�ίL�ʫ��r���s��]I6�s=�  .�`0)��W��z6ꪹ�雹�雹�� �^ �HX�.w��&��I#��U�Mڽ��d  ��ʼ��L�Ω3w/;���F��ޏ_���Z��� !U?� ���|����"�;>�ِτ�b�,rV��?��I:��AZ6 H��(��i-[��J�	*_F9�߉:+b١�	�K�Lʸ$>FO��(���j����Y.YvI $~q��v]��'�8��2����%X��S����:�Y�|��e�8����;)��T��V�T��	�O���,Y�)����?M���?{����v?��F2g������`�*��BI �	�H@$7�0�l�:�k�Z�y\����}:O8����F�b�s�e�	I��f�kO.���+��v�$��K�1q�s��<[�˥w�]�Y�f���O����:f�9M�V������g?���zxc���jv2EI�"	�q#�}��Jn���;e�m���3�bb��KS��d H��UR��,5z��$@HP"Y��yh����.`�䌩|�vغ $`o�_1� $r�Ryg3�7�ہ�n�^�QbN��S~�>�sצ;��p[9�tw�"F�ۏ���&�^�^��g2F��dQ׶�)J�WӒuoэ���z�vM��F�u��Վ˜t�iL{���%��:�$���Q#��zOZ�rt��66˅Y��Q5��u'�5���?���'}��w$S�	��� 