BZh91AY&SYy�u��#߀`x����������a��          � � T_mv�J�) "����ET� *QD��8�"V��U�v��|  �J
�P� R(����TcD�@h�	P
�֐�� ��E%%�    "� /     .�<� SCР��  t��=htΌ��FG;9� fk��te�� ݎ@Dw� AL�Z���]�U�3�e���y�U��nދ1���E8����O��ԭ7�ҝ+s�a�8�j}ڮ�w ���     ����У�Vw|���a�3�ǽ�˻Rp �w=ir�f\��;W�n����oMkp ��T����ַ��/ b���^�9�my�G�yN&�dכ�{8�^Ǐ �EY�YN6]��5�s=���| �x0     [�� ���Yw^[���{��z��x�Ϡ�m����&�{�.�\p����O��m�ݘ �y���.��uW� 9�����yv�y����D�����ԧ3T�;��˼�U�w��<�  ��   �E} u�Wչ�Ԯws姖������>��}���{�m�o�v��z^ۋ^ڸ}�r|{*��}���Wͺh�7Z�� �{�e��J�k��y=�y��oZ� �W.�\������۵-�  9�|     �N{� Ə���Sɾ���h��:� �����3.����^oR�{��5�Žc�ϼy� ���K�y��o< =.��s��η�/1�-Woy�׸ Q�zq�����o����>�                P4��)J�BaA�bh@�2JR���M�4�h i��4 �EO��IS52       ��R�4� 4      O�$2�%( FM4�C
B����	�$�&4&��h���?Q?��k��P�O���?�o}�5����U���ޢ�*�TEO��*�DAW �@� "
���V"
���J�u""
����`d!�%�!� �����!��'�'�H�"}
}:���>��~�� ~��O`=���e�S�O`�_�>��p'�-(�ҁ�"�JP�Ҩү�@
�niT��ES�R+����%�O <�Q>���PO`�`P�O�MB�Њ} �Ҡ}w('Ъ}�H)�j9 'Ң} ��+� ��P���P�P_�S��Z
E;�C��T���?B��(Ђ?I��������J)䈛� |�$DN��Qi�!6Hw.�}���S��C� �S�a���@�!�?@��} HB��y>O/ $>������G��>��O��_��>��5����'�'ҿJ� }���!������пJ?O��}��nU>�>�>��>�>��%��} }P��J��({*nd}��e�D��pQII�{ �MC��{>��L���|�<�K�\���=��C���H}!��b}!��K��%rW$���~��~��@z��=��D�{(R{�>���} �BR�!��{�|�������w!�P�})����� ��O��Q��@�!|�<�<���d<�����!�쯰��>����)�y y#�	�/��҇�>�B���ҿC��j�����\����O��C��_�>��������� �P�)�NC���)�} ��H{/��!�|��� �#�K�O<��Od=����C�~��_���~���\��_�O�>���>��@'�nW�_ddo$�S�|��'�'�Ц�>�}����C�w/�}�����w����'�H}	��?F��O�>�܇��?Jn]Hy�y�I���
^�@{'��>����>ǒ}!��D>��d}�w�>����'P�'�����~����N�~��_��@>��:��`�M���/�P��}�_��=��}��}��;�e��ܿJd��'���>�Ԟ�{	�`�O���>��>��>��>�����>���Oa�a�_a�7>��K��J�w��J}!�G�}/�}'Ё����I��B}�^A�A�;�����>���@�Oa�e�}��=��=�$�O�5(}�����J}/�}'��@}/�}	��B}��*��{/��짲���>���y)��;�u��;�� �N�~�����S��C�S�W�~���~��}+�#�~�!������C�$i}��e}���OeOe�r��\���>���_�=��C����>��_�>��
W%rW���>��>����);�
|���C=��¹��XA�s�'�쮻��)�G᫡� �u�j��*�+,.�Wf
���%q���;�`�B+0pXq�!}m��T�C��7C�$����8M�Y�ծ��s���Y��\��|< �y��qK5��ɓ�L`�8;.�QJ�U�9�wW�+��8/*�B����`b�t�/���L6Ia��V��T!��0��$�˾��/��}��^�[fӻ�n� w��"�J_Gjû⸣�ָ��0�!��!J#�I��ޕU̫�Ev��*�
,]]���w�C5˜�(�����<#���9y�ʊd.A�%�[��d�|�9	ܛ�,{��%o0v����8�K��9h��� 20���Hk�Ѡ����i�����Hy.9	A�ܺz֍=GT���-jM���
68u��4�8��������w���ýk ��Ek��ե�Жi������ל�ƫxT:S Ҳ��Uf��+�9\�=Hg-VۗW@��!24BT�2�-W�=og �3�>X��w;$�i%�Pc�Q�7�7Q�q�[à�sp`��F�XN��=8j�}F;ѻ6i`!'���8��m�N�w��l�q�Vb��17�:�r���9�~���V�S��^�a���@�0$�0�!�2Ɠ�Xhc$ۇ!+��m��rsO2��:�9�4�9���4��Mɤ��l�i:�A݇[��=�(=����g:�{��O���8�QI3�`.=��r��cܜ3a��k���c ��B�M۫%B'x0$r�C�������1�'����0+,��N�3^�!�n�T��\FC�|�o7�Y�	U�S�j�E�!7H4&�Wzi��%	 ����J0����C\�����zn8�ͧ��[��j0�겥��(��,�QY#���o<��>e��m��6iP"�Y��%/��DFfMj�-Ztp��IoE�rH�.�l��pD"����_]� ���W-�鄐�יu蹾��y�t��:{�F�c�P�AǨ��n�2aZ$�N�A��cʵA��%)BP�%	Br��(JR��(J��N��*�`=�dYa\MJPi<���(�^�3p�:��Y��I� E�b��o�pr�k�0P{'�l�ݲ:ٖT�����ܤ�GĘz ���Ɔ�!�Pfa�ᅻZ2qr�	�|rL"�g�:s޵�'!(�26f������.Q�x�9A��(Q#��,��Վ���,z:������ 2�@�J']w�X����׉��Vc|�� ;.#k�ɼC���gA"�p�5��P�����G\�/c�ҠJUJ��")���w�g9zx[��ǣ�@vd��fh��`G:O)�c�v'�����Ἠ���	�шqa|2Qz�ȠM��,w7)�0�S�����:W:{�\bm���Q@����is4� @(Ҩqe+ӡ��g
t@TM�EFl�J �%���맮c���@�4I"$����@�[=��)]�XF8�3��h@����cVk��5�fo0d�d%!��te�[��{׽��xh�׶�	��58:՜<藐�f!(Jl�L���n%#��q�z�G���Ru	�a�;$��79Bj3�d�>f	BP�&��d^{��Xp�358fb��h�̞ƖD�LhJ��!+��������H�{�)�� �4�H�bZ^����s�=�r�p0�V�i
�F�S4'C�Fǭ�Gl�&�������� D-"����&i̹�5	왭�j�Te:��oD@1�a�J�yƈf�� �������3�[�I83mKW���@�E�] �4�Q	!��;�5�LkFPxFn�w�l��}�I	4�U�r+�=I�rVN$f87Z�N`��^u�:nZn��C�Dq��{Lt�Z����� �0�t4��qe��C���ۜ�Rj��r��TBN� h��L@Ds�E��BX�Έ)t�]|3W8H];{�5���	BP�'r�'�a��8�-��W��Oc�O 4jH���
����+2H���Xo�0,��mF���4���H�����0,�K�
���".�q�A�	P	%��8�����B4S� 3(�!�(�`!H��XO8�5�u]�=bń��@T
7�;k�ܢj���/!K���B\����0!f�:LL����p5a��ޠ0�[�w��֓Gn���_3���b�e!�����<_V���-�7�Yj�΁�@�D��j�V�8��z�f���l�fܐ�4���,_* 
��W3y7 �J�!Ґ� $H��D�l'
v:�v �m�tŬ�/��nq��1S�	#�j6��ʡA ��Kݴ�˰������8��&�Tb�,h�8t���H��Ɗ!b�Zd��8mx��DX��8�]�1�@=,@�B�c�BZqjth<����u3�A��(MK��!�����F������n� �l�Z�l6����ӳLj�q5	`�ދ8��24o#d�q���c����=jv�.=�Á�`����A
}�Sp��t8�%_N��B�J�A��e{�0'�t�F�'m"���I�&�����giN�����m[�ݹ27�
4:�&pˡ�f�2��:�F�1&�#Q��d�´��ɉ��5����0�p��&�Ɠq��sL`h����TB)�k��}�	w��iΌ��2�̄���4�!���"mꦜ/����K��Aka�{x4_t� 6�t0�*�� �e�d%i��֠�����	�&BR��5s��r����9E�4gq��<�M��P�/�����1���9b�gk�a𓸚�17�b=X���A����LPy�>�k^u�κzIt�����MD�A�lrM�y��nmf���n6T��6�;3aHE`��7�f�3�ͼO,5ֵ��54��	`�`A��'Y���w�Ɯ᧸:��2�i3��0Jαv����ܽ�K�%��NM��\�׻]�nM&I��[�g�VvÎ�TC!Ѣ
���΀��s� �8Ä hG��`�E�e-I.�$ �j��2W �h��o��}�ĉc�2c5���dkfT(: 2��_:�ɀ��a�vX�&�m'!²TPE����Fxo�y�m��̌1c01h��
@�f����)M�	N/m]E��q��[3���lr��cQ�S;���2q#��e�p�@Y�����u�m�(M�1�۱�\\)U�Z%{۶�)��Rq2t�	B{�%�#�<7Ӣ�AàՋ�H�*c2����Y�8Ɇ�b��d�! �d ��;���v��ȃMe4�J�%*b� �I�`2Td`�6�	TVu�tp��
��@`FQF�T���h�������hw2u�&����t7P`�2��4�5fӒ��7�d�1�v\�P�k�(J�JCV�hJC���Ѭ�c�6�XÒdg(�<���,%�N��%	N� ��̓sd%NG �ȓ�f�7�.\���$7�9����剷��m��z�l�Ԝh^��#g�I��k�T3�c#&�3#qߜ;�� !/3�o����8�$�#���ŵ:B�`��Hh>�F���
�A��K�5^�Z�FN/��]��bjv��a�B�:3S���#F�z	���u�.���8�(S*�2L��pְ4���U�xF�sG!)���Q�d%�="(`1�^١ٿ5&���)��jp4�x�g�!)w&1�bN�6f��r{��Yy݆�h7/m	N.X�'	5,�<�'
�bh9�q���-�����
'���[x���I�N���.��9�f�hѾ������]�f��PxД�zhFr��:��WP��!Ԫ_1QTSc��a�<B�HO`��tz�oЕ�SHY�C<�uߴ�K�v8پĬ4�f�w��&�Ԝ7'�d$EE�%�
av���V�b�,tEj� ��R
wb1v!5 �N@d&��!�$W�F�(t��J��(J��(J��(J��ӗ�w��^�`jP�%	BP�%�ay�^���q޵�M�i�f�g\�	A����8k�D9Ld��Ho%��9׆���uNo15���GSR�P2�2C3MQ%&.�y�����پkҙ���Ƭ�cĚF:��t�F��z��)�G@,� Uڴ��f�tCu��ǛC$;��J�DG"�'UNNѫo�VɈ���P�Fg�m5�Y�d���3��p�v�9�'$��y��uգGln]��Z��O�\��b��bU���rFw_:Y��˂��p�`�*�t"�R���n�� Z�#F��g1�mu�\��9��z<t.���80�aA���PH�]�v�d�p�C��5�*sf��k�5������`dF,p�E`E?��u	X�D�'�&@ȵ*����$�r�?L�\]�	9��d����#̋��k��w}��擆�[�.u\����F`�F�c��iٜ�d�1�g�20�FE��T��5�V�A����Y�,�@�f=.N�$���N:��i9�N&Xl�;Ѵȳ�=��}�J�\�N�C���������]�@�pZS���٩{r5jNZ��S �@(bd�)������!-���|@����wه��� vB
]�0�	
�>n��ֹ���w1����-��╜c��G	Lz;��H�T�|�ہ&�<0��HJ����☪ڀF���R?*��j���X8y��'G��1�X{\V@8�߼��͝�������cۓ��%����O�=�:��L6�E�Vs�z9�z�h�t�eA1���@D`���K���Yh>SD��r&��BZd�鵫��	�s�����w}�l�	ˎy秮�ú=2�<f-�B}�?����}���}/�$�	�I$
l -� k�    2            �  � A�� fYv� � h�8 �      �   �pl Hps� ����0�Cm� l9��l��  -��A� �x  � 
P                   J         ��  4�\ )@@��չ��$��k����gtpTlm��^l�n�vu�{v9�ٚ��j���C�`펀�%8���cs�q�|���9�%vV��u4�k����,��3�`�zv���r������2��`��Vѩ������:����� ۤf%˟%�ס�����&�ؓ:�I�us6�M����rXs嗖�z��f�mzѭM��Ȣ�xy5i{n�'FI��11�͞���{8 ,]�YM�a�s��� �e�m+n�PT9��B� A�I�Ӷ��  p�l���m$�` ��3Wn��ۥP�Ԙ�@��6�Y����s��%s�  �M�M�+vi6�knZ 6�(l6�d�W���T��@A&p�Bn��ŲPH��M�4]� �-�����u�^�m�� H��`Ѷ�zѴ�N� ��*ݱ��S����ol�Ke��m�tUZ�Y-�j�
�n����]2]� ��;vZ $�p-�$  6�m�$�h��γ���H�a��� >%�moP��N�M,����J� m��� 	�	��4�0�i��El��U�N�VH��� 7�=�.���ln��7a��9�'5
;��WPF�q��&q���`}�G�|$7P[n�A���6�f�@/�Q|���`�e�vI��[Bڒ�KmW<�*�-	��m���m:$e�9�����۲�.Z�L�n�R:���@UMڪ�P�kѸ0�Ү�.Fu����ki^ݞ��N���Vԓh�n��[)uJ��ĽP��GiV�sM�ä�'�)�PJ�Sj��ͪ��W�ڟ UR�)���;�V�Bڵb�Xn p�y
���ہ�mCi��[��hݸG�j�fv�P�.uЗ]m�A��!āJ��@��J<��s�w���|�kpTm�e�"D�li
�<���+n;�
�V��{-�M.���-Tk��.@5i�j��gC���Q���>R8*����u5�����l�{"�ո�8�Ba۞�I�	�x��@����[\8 8��Ӷ��� �`6���\��@R��[rɱ�H�lٶm�l�kuu�m���W �J[@�v�t���u�EU]�԰U��+r����s`ݷk���(H}Oy��� m��F�޸�mmH�uf�p�gN�`*�VƳ�ڛBD��p �hņ2�е��ObƞnÁ�^�a�=e���zK�9��E���t�'JrnĲ�P!5mUAKE�l��^�[��M�M���
�]��iS�p*�KUW�����F����� �QER�]slY���,�bM��R� �r�Uj���^��-�4̮�.��F�X���/�6բ�)�-�05m�&�SjVV�s!+.��+;*&�4��U�{(v԰V����5��Vp)�nZ��Z�V�@��z���b�m�[B��"��t�b�!'H��	����嶺�;�հSiU�-�rM��� R��J��V�:ت��u  �	��:�Iv����6�O>k��Z��I&��5���L�  8�ꋛ�M[6�m&��m9�.� ���k^��> | F@H�K֋@u@+�URŻ��{�[�pT���TTP�*
����M�*sY�9�T�_���=>i�t�<���uP� (0` ��8�/^�@�6@b�y22����i0o>F��zܐ٤�[m�G�;ͥu��nÛlmm�m�[@ � � URŤ��j��%[d�j��)YZU���i  m�[[l��UU]Q�d�>`���:���Зu�)-U�UUT�� Jt���]��L o���[2`m�[%[�
Yf�K��L��[Mj�^�T&���x�L��������5S8�۾���ˋ�q]�z� �ɂ��>k��R�em�^�%��!*�`�Y�������:��v���P�� m�Bt��P+uS�q����/	��	��<���;r<d�%�pRU.�	ۮ����s�e�j��,��.���re�&Ē-�N�6i��$�-!�Bv^�78�{c��f���Rt�ȋ�p�)�m	C��
Rx�3c��X܎Q�Y[`Acm;vT!�n�`tr�EUyj�n;vວ��l�*�E�Ҥ�6��. v�
�U�P��l��AKk�6�p6Im�R�$	e �9$�a�m�Ͷ	�6Msm���$n��)@��mmű��ͤ�C�f�@Z�� m�C�%�dkNؽ5	V�6A��X��v j�]U6�K.ܶ]:YӰ �I���6�W��-�3{p�uR�(V�%�D��:�H:@�J��scmہJ/S`��	�[g	0>��ޖrѶ��A�Hrۭ�P9m��܇9#&� -��lp[@p,1&�6�m��p$�À  8�Z�UJ�*��V�+�T-����H vY�n�J�� lU.�5.�U�]J�[*յ[;-�g��X�[m�Yc�����T�\�T�Ѹ��}�� *I$m�A7,�o.�ذxݷ���a<g����m�+�` Hչu�i��q�n�K]���&F�ݏfK�2�N���n���R��A�%�T��	L��&I"ZZ�I� ��n[���݆�m�����WRUrIZ1��P6���P�n�՜�`  koi6h��mwm�@� ٪��� m�l$�`*U��:�z�UQ\Gi��>���`6�d��� ͫe�  $����'-2@��橒Xu��kh� RJ�/Z[v�&I�@ [G m�kn�8�m�f�	����m� 6�l�ām[@�$$-�  [@��&I�Í�I$�$   �ޜu��m�s�����-;E��l����r@-ֶ���   p p6�$�  k���jV4+r�j���5@[R�4�ԫUJ��M�:U���x��Ҭ4WYS�����[R�5���`��qoP�@K( ��܅[��m�ث�)k��,�ΛxH6��Y;e��:  kn�w@��-u�on�:�m�`����� �E�k���u��Q���UX	Pjͅ��$   
Q���M����v�d�-I  �j��Ij�IjH�%کV.�݁�V�F�� '7E-�n��m)A�jmT��m���y8�᪪Gá	�n�$�.�I$�@R���9V���S�Ԥ� Y"ZyZ��Z�kv�@$gM;f� �L��5Vm� -��mr�2UGQ@Pm;[lm�8m  >m���.�r��  [A om�-�������UV�@UQ�ʪ]�6�)���-�iJ  i6 iۤ���ȶK��   �o ֱmA�������` �vָ��UHlq��x8reU�` &y��1�.��Kv�Y4�ݶ��xn�E����pkk�@��,*�]Y�h�(��-�l�<�E�I.�u��IŲQ�h г�� $���m��zi�썳*Z��  ۶��� ����� q!m�k�l�4���   �al�&���Ѷ� 6�bC��I�lH�����@.�@$rN��l$8 ��[��M�[A�5� E�4���}�N�i��G [I��۶��B�����`   ޠ	5�Ŵ��pn�l�  9z�m��� H  <�j@h$.�P-�kk���[CF�\8 @� ���K�m^�-�l -���� ~ x�i�H6� [RmZۀ��ۻb@6�4� m�-��6�[@����  ֲB۶m�p�6Ͷ@ l[E��Ͷ�p�O���-5ܠ ����6�t��6��0   c� k2�vm��ճ�lh 6׭�m���m�i8 K( �J�ր�^�E��,a!zս��  ��,$��� ���(��J>үO<�(2t3:�ۈ)����Z�gr��.�.�K\�R�k�}&�$�v[/L� �a�T.��&�vj��Y2$���v���m����`�5�d��  ��[D��mt �z�` ���6��V� �@���8m�     �ѭ�]5�M���v kV��v�l���y�{l-��[@ ���m�� []��9�m����7���f�k��Ci6$Xam�c� ��im�6�h ��Z�nm��-��` ��K�$����\lڭ���{��o_�Π�����x����>�ڈ����)�7���p?�@G��FVNf�X9A�QNfHTHeU��$-X�5Zʭ�1:�r*�2"C'3V�FfUIB~?����#��R!�?�~���W���ff� pwx���p��݀ ���� w�1� ow8 ��� ��� ����wq� ��`� �1�``� 6 ��` l p  �� p� v7l p�  p�  ��� �0 v�0l � pl��lpl��lq��m� ݷv���� ��� ��� ���` 8;����t4O����6��'�?�����c�\5���Ǥ	��%X!F	7��p :Ѐw �����pB�'{���Pd��x
���+֕�ڐ�
���x�y�ޕ�M
h/Kӝ���|v=���.� �Pt�lq�{��z��Y���s����Ez�~
=�b��	꾨���P9ׇ:P��&�	�P4��;�@.��6`�)á W�B��v'�I\ר�lxv����ীv"�*d�<��� Q4T��S���b����T�<�4��1� R�0XA�!r�z!I!I� ��eSЅ�(��G`H�GC���׏�m����Q�(�OF\C�J��[�����@�q������!�ǣK��v�K! ��P0:T;�n��U��D
H(>�!δ��ؽ�x'Jb���1;E��pP�;7���T�WF!v(<AךT=DT�:AU� ��4$I@@�I")�I��(� p��f�pM)�{k�(ɯD@��; =WO�G5)��J�$�JS@SB3 �B�� ���΃��E8(	�/G���H����T2 ��;Uӷ��M�׆��'<z_W���_T���H*{�4 ���+�^�1Mx0!��<�+��x�(���kBkX�f���=�+�r�{�}�U��W��{�E�*���������UQUUUUUUUr����    S{��ʽ�U��kZR��ꠂ�����������?��B?������#m�!�9	6�۟����ٻ�����y�o��ց�%v"!�8e!)E��3R�C�a ����C湳��e������u��k��]�}�B,��w��`}M�䮌��]���(h��g�2��e��x��S���6��-���{���  �|��&.� �*薇qD�J�jk��Vm`   � �T,��<¬֟N�<5Q���\t��<�i��DD�q�����}����=N,=�*�ә�����Eam�gWkϳ�J*��ss�wϱ��2��=���v�7������������w8z���
øN�VrY����n	Ctc(u�s6�<~nc��뭛���<'5���`PY8u ���n~�&{>48���n�j�3qgvU"WF�~e�d���5JD��P�>'�eH��$+ ���������[nͷ�(�d�8P^��\+S�ձ��3=$S¸�A���>^&�>�S�k�E4s�%�F�a6�Q��ēoH�r}�su������]���)�n�k�x@v�& �;ume� ���U�vʼ������5a��� aK1ȣ�F�j�M΢P��wkz ����������������t��+e�"�����N>y;��%�����V�g��u�&׫0�Uv]��I���9����F7ns�;����)6$<K���Ft刈0��n�K�:r�xN�.ѫ�3[l���;��4�g����rtl�L/*	�LΨt�t�7Rǣ0;�ΐ	U5�m�!ME좛��*��	cp����!�L��7e �1�.���K|wy8[�	�xuR7?;��N��n��^�u%"�S�4nR��U�Y�����k}�IΪ`�L���lLrs��)V�^�Lܺ.�Mܖ���. �E�<�S�;��i�u�̠T9��9fFWk����2�4 �;<肞jY�va��5Ѯx��Ӆ��л���=�t�I���UKj��V҂V�	��h+���l���j��ɴ������b�]�1�n+<�VPj��Mp�$E��O<��u�l��Z
m�p	9. eYA�p��J�O&Iyi-
��p<�[��W*��
� �ZxQͳ�櫔�j�� U�F9�m�َ Cv�s��p���\�Wk�ўA4��rKn�Ën��ǅMi��A���݉VV�J�/��&�s��E4�fE��oG�������y�=�/� �${C�o�ͨ!�x�(�/���>���:$UT+ )*�<V� �4�Տ�� K`䪥C�\�LK��ᵑ���ۂύ���ۆ盞Yeڱ	�n��[=�v;^ ���:fz?�ۻ�hثm����I����F���aCaR2 AϚ�9X�_�_m����Pm��\�F��!���Vkn(�̲a��z����g�p�3��;��ٱSu.ڻ�ݥ�����ulۭ&�`�p���	ļ�^$���sc���	@q�:ѽ�<�ڎ�|yN�ލ�"����&v<r�ǰ�ʽ�86<<���`L��l��yDܙG7]s��W���2��N8���-8q�9���U����z��Tfk+jD�n!D�빻*���\#��\�sn����r(�A�
R����,���m�f���ml ��qDm�w�b�\�sls7`��U��3��Z`"����K!�E�1=:Zݫ�gl�7��	I�Dq���'$#��{�m��ѷC����������$��HIr9$�\=��
�т�h�(Kw�Y��\�sl27�6����h(JN�n����{ܛc�� �bñ�Q���������u�w6�3v��ͺ�G�M�b$��M�]�n�s7`��=�:�}����Q��JJ`b�b�]Ŭ���8�ʨz�x�^� �TWT�u�ޝm�<d���	#�݃�3s�͖:N��%�m��)Hy� ��q�y��g���\��gГn(��D�o���g36ŏ~��(��3,C0, �!�ρhh�\�a�^���eޱ�
��
rHc�;����n�9���{�u�����D�BYq6���n�;���{�u�w6ǀ:��4�N�P�Jsԋ�vC��q�-έm���=�X�q�8W�+�)� ĂI"A�iBS�;��=�0;��8;����>�"��%d.�s5��������3���wr'��e*�@�I#����́[U�۲WO{
��Q�Q���Ia��d��{ݝ]��}�QA�S/�@� �C�U�UU�����>��%�i9"J@9��p����ͱ�Ѱ���w�x���6���0�Ny����0�YR��V|m!�#���j��:7l��V�[�`w�ͱ�פx�o�sǭ��Ɯ����z�0n���8{�u����8D�BYq6䓜���nl����Y��Z5�Ѳ#,2�m(Jr�(Q��o�����]��X�n�;�sIL6$!&� �c�3]3��o�3<=(ss``4������E��%�F�*����\�T�푱%�n�1���12����Y|ܽn�u�7:�yGrXڥS����a��m��\2�s��[!�0�k;S�g9wn)�qM����9u�;�Dx�8ݶ����Tڲ���C�Ȕ��kJ�A�Ëĸ���*�䶙�sY<��F��n]c^�.����nC�D�t���r��˸7:���v&䶹z���x�w���˃�g���g\O>.��l����.�;��k�����}���V��2X͙m%�!rG\�o�s7e�v
6���[����D�QQ$��݃����������h�����%%wv����m��l�t�3��n(��7c�Y�u����3v
����}O�#TS��x��c��r��������;_e&�>���k[���U��-��7@�Q�G���n�������bn�� ��rT��,��rI���{�{��A�������l�DT$8�b����/vp��#)߈�Tڃ��n�/����ݔ;�E���$�d�.�{����N���fϺ��e����!8�  5�����l��͈�o7i��!T@�,s7`����q���7��ӥ�$���@�Km����o*��Ps�n�ꞩ]���D;p]O!�{m��̠\jÒ$���sD����Y���<��t�Z	�7P�#��[��� ������l{�,�����I��Ĝt����w`j�� (�HP"�IG'��x�G���\�6yy�}��Ml���%nI,s7`��8{�zF�66C"2D1	N�͂qw��w&��n�;�:��ӎ8X�(�q��׮�Əeׅ�vqXn�#�l���:8S��Vz�cg��q�\�ә�������l���<�eXt�e��������.�j�3`����m������$�H��`�,w��΍�{���ͱњ��Q��D8�JJ���z��n�9��Ժ ��ܠ��������z[͚ͨ��7c�3]xW{�������x���F���ˉ��KpB�v5�l��-���^4v�vΗV�09�:����n7]�f��n�8;��V:�wC�1�J26�rX�n��C���0���s�[�$2#Sf��̓���W����seaŇ6B@RrԱ8������l��OIú�0��)9�:�sv�;�(pw6<�:e-�d����v�M�f�q�Z�T�p6Cv�3ו�����Y6�=6m�][���v�q=n���Ѣ�M��t������v��h�۶3O�a����+e�F�'�֘�֪��<	�Y�'>۲����lB��{Bf^ɻk��ko����k���vb�f"�qF�:$b��y�'[GF�X�۳���f����5�u��I�Ε4�E��oe���[7�����]�����ۍ�v5۠^h;�'e�v�kp�i�MlNwP�Wv�7)�]�m��ۂv�h�} �pl{�������{D`��7 �se�y�u|�m�w6����6�l�P�|��_;�~�(��@��h��^@Њ$�M�I�W��s��W;����5:�Ł���1Tm����s6���X��k��=cw?�\r��qk�\;Ua�ն�'7�(�W�1��ۭ��v�j:�[�곢77�X{��w�����
 Wo� ���C*I�CR�sX����)�H�@�@P��@o0'����{�ŋhb$��m�W��6;�+�3}s]{4����!(�r]Nw6����g��!�fh���{D$a��'*��l՛����c�� �� �hP��߲��&v�P�5*�ì�m�k=m8��Gdw��n������9n��m�������;����`o76��݁(T.&�GN:�����{ �������G����dm�$���@;�ث��|������������y��m�n�f���fn�fe��mr�А�� �LJ�y���	��C�}��{��~�����~y��_sj�p�����!t(t�i��Ͻ�!�I���{]��H�w����L��|^C��ͬ�4��5��|:�� ���84%!���SԚ����@yvaǰѯ:5��>�]��LN���v>F�1I "X�iY!�*ezD��\{�;��B��͇A=`��(*H���F��ˊ�А		l����Q`1�����HB�:M�H�^'��e�b��Cv��Ї���ؔ4��퟇��mK�~�� =D�M��`!��l�H�l� �� �S�5��m�	�/���U?���翙���}�GV��T`T�]>u�����k�P;�O|����B� (�=RZQ��6b-�`Q ��p5/�~��y)@��~~k��4��￼N�����?M�qg�;���&Q3%2I,�2`I���́��7��ԛ�3kf�Z�h_}���G�w|]FX�m߲1���k$m��ܯ!�ۂjj"EC�s7[���0��q�V�M���ݷ�ԝ}�ߜ^�i߽���iJ�=�j���$��c��RL�v�jpO9Ff�V��R���}������T	�x�)�f@�k�tS2d�3?S5��	�e"l]��1(�Q2�Īd�(~��͏%)O3�}�������Mc2e��J�P��d	��d��	�/$�Ț��	�FwE2`e �=��ߜ�7)����\R���h���?��2``��t��� �g ���ݩ4����~ ��7����}����j�3���B�Y�y��[�JR���w�~�z��$??DO�����}���`���D���<cߋ3�
d���ˊ��my3�[n�Ħ�T�!�YV�n�\t�m�\�֋�k�e(�??8qJ��Ͼ��R��3R\38͂N2���MbL����%��!�l�ۂ�5@����#�I8̳wj��$������3,wfO����s�2ݼq�3 �2�y�4�1R���9)����8)I�~�����V�u*f@́6gt���2�G�!
n�zٙ��_��<��R���u*f@́7��)�d�N&�7v阥)?>���(�_�Nf��޷��R��~������Z�����R�������);��x=JR��d��|�j�}�g����Fq�@cM(�R�ڹ$�gC��#�[X{����8���LGc��L�F���;�<3�@�k�#^ziK�.��û]��ҜXf7]F����gf:6���;V��"�ϭ�N��C��owU�g&��>`�O��O�8Z�3Ë��V�o�YS&!yl=h]�Aa�����e���^Y�mkg� e1]mmk*[��ww�����1��֋E�F��D�l"�`������N��=�b�����3�t���Z[۳X�{�z��/^}����R��>��qJSy��}����޼��0;���޺8�U|��~c�J	IQB][�+�}@̱�6)%�}́��w�5�&e�˸pR�>��$��%<����Y�ۙ�{��5�pR��>����)J{����p�q�ݯҚ�d�wb�`����s)����6�����P~��O4'�����������c�S��2)� %�˹Ԍ�;�Rk`fB����!RTE9�d��*����������?U���~~f��C�4�k����ԥK���gG�)?y������_���؏Kz�.�9� {d�)��ٹ��阂n[P���!HR	a)pV�MR���)�2_}���Ę�n�*K�;4�o��)�ń�%����D�o[4k[��)<��s�8=G�/�وb]#�Ý�ܧ矝�┥��}��)�{��~�.��'�w�?'��;�K�M&��2�߿R��)J>��$?pԧ���渥(	�;�Rk�$�8nh�28;�3�g���!���͏%)Os�~��@��fu&��S�\�ͽ�J�`f@˷�1��8�%E	wrM>��}A�խ����(���>��ܥ)����)Jo0|�߶��rd���?=�3W�aj`"����藍$��ch�u��|����'�Ͳ�6ټ��W%�/��O������翟���(~��R����~��R>���د�*��{��S�H�&&i5���nm*I~���3 M߿T�P��������pR������ԅ���A�FC�����V�P$V{~�׾�JS�u�s�S��^��1�`y9�M,�L����h��C��}'����2N�(???8qJP�^���EHR	aGpWP'�T;��ޙ�3 e���Mc2e��J��&\3�����Ṕ�nFD;�(Q ;����O�u�R��>��Rr�������??|8�@'���JR��k�s�P4���������֭ff���u�d�ۧ��n������iP���׶q�j���^�x�D�a9���z��JS������(|�߶<��O}מ��S%)=���WP&�:���B�&"�6�c�يd>}��G��'P�S��_~g�(z������)���Ê~�JP�{����TP�w$��}��V��_�;%)<��~��!�9)��ߜ8�'�H�ߧҪ�P&�wwn�AJI�*L┿C�{��~pz��>����(|�߶<���S.�D}�<�$�2W�gʪ�~	ߙ�ϑ�Ϲ�]P&�C�o��A"b����]��NK�����8�)H{���yJy��8�)Iߞ{��JS�>}>�~:25�����V��B������x��,v�Ҝ"���7绯�S<5�|=s�w��P4>}����)���┥'~y���^�(������)J�>����i3{+[��\5���)J{���8���)��R���}���R���߿��8�)C����䟽ຓp������f�n�z�Ykz�)JP��~pz��)��{�qJ$C!����c�JS����!�.�ժ�BA��*���5�0p��O��o�8�'p�>�o�c�JS�u��hO�Q;қ��?O�P4�����% ��9$/�>�����6��������`���~��R��������ԥ����R���e���@~~~Fg��ew�G�����j�wf�����iZ{lJ�l୛�'���OE���=��	^9zl�;ڒ�7W<��TM�ؓ����B����;��ȖW�712[հ�����AF+l�۰�XN��ƣ>�=�����Y�����B�k�Sj���m����1�kל3�'z�m���Fa�Z������#��3��÷ �'��c'#nv�u[rћ�oY�~ v�����[��oИ��mitvױ�K�6�?w�}�9W/�&eٵgĒC/>_�5v�L����9���;��ߙ�hO;=��ԥ)����Iw�3'd�I��o�MC2e��;-�����8T��5@������}�5)����qJ���6���3^j���UAf��J�31��y�|^�)O�?3��(Sϼ�c���5)�����JR}�翜�)C���0�!�LF�p]P&���:�߿~�y��J}��?3�R�>w����F:_�$�˧��3 f@��qߦaC<ʌ���3z�ǨS�u�������CϏο8=��d�����\R����>��hT>��Z�^q�#1�A3H�#��n�ӏv(�\"w=����ֽ缿|��w>-�{�f��┥�N����ܥ)��o�┥������JS�~��qJT�p�xw�""i5��on��~)��ϼ1&���7�~ i��D��_�(z��ly)Ju���:�S��>vm&��k�2hl}��ʷYk{��7qJR��=���R���{�q7.Oߦ:������R������Uj�49�Z�.2��8eܻ��TW�*���?3�R���~}����%=��p�'�"��{���)߷�sZq��(ȑ��WT	������\5@�??1�??:8�)K���ly)Jy��q�Ęo�7��K�D� �0�tS��\����dL���;[�x��\ls�l؛j5tUw�(�%�q�㺬5@���wR�I�q�l��)�f@̽��zK�b�J???~�{��rR������7f�ۚ7Z��)JP�ߟly��"b��~�_���)�4�~~�~�z��=��X���h|�"����$aҐ4�Ԋ�V2e��I03 @
�si5�~	���;Q$���W��t	
B�$�DIREJD�4�_}���_���)��w�`4߾~ly)Ju��ZDe҄�$IȬ
&�ƀF�}����R������)J{���ԥ��v{��`f@���w���o�ԥ)��o�R�~s�=?6=�ҝ{���)JRu��pz��;<�~񳍳���Ÿ����hD�_�jT��baЫ��x�x>��{m]������)@�>���JR�y�}�)JC+�ͦ\/�d�;��I�&_{_`?B\j(#�]ܐW�4���V��Kx�����{��;���qJR�os�U�DQ5C�w�ۈI�$bf��R������ߜ��2S��.)O���(=>���R������qJk������%L#n5%��>���S%���2��d	�'�5��df=2P�!��?	C�A�4z����)%N̽ח��e�z�X́���fo-ѭ�ճY��R����>6<��]���wWs�2d�߻�&��2���u@��MϨS>�J?�N8�%ơ\vZͶ��i:���z^���+���T���Cg��(�\�:*J�@�[Wa���}�R�����~��)J}������pL��0&��Ҙ�f@̻#��"bZ {�f��┥'�����=G����<Rd�Κ3$ǭ�d̓@v��������v0ob�(g�����陙%�g~{)��v��}}�tIn���k5��y������Ϻ��*�����ٷaɓ�d�ouqH���#�'"9	˹' �{�����}U�Ww��|�uqh>^٠5|}���ULʗ%�l6�n��m�����{���,����<��|���cEUy�4V�r;؉�C��K,$���$�Ӛ�`!�'M��03?p�rZ���_xiڝF`��<s�[=���/f�B�N�c�(�)�`F���DK��xt��D��\���ɡ)
Y�"&������HB���zu���2w%U$a峏�Zpw=��@� h*� �M���$P�Ҍ��d�!$���)�
�'	t�$0@@���!,=���SZ���ax+����ˁ�v�v�Ӧ��4IT5!%@��������N���;��4rW�6��E�Ѯ���Q��3y�PA�oPFĪ�{�F�A���u���D.h��'�[�X���G��%�tʤRTA�������c���)Pv�Mld�9�|__w}z;������    m&�ɋu� nL`ӭc����    -�l��/�}Dhc�����R8ޘ��u'�%�g���`��x�}l��3ںۖvZyu�*��v�D�Ý\$l긻Oln��	6Q���ke%�������g�Ć��f��ںݶ��,�;�c�awn�곕�{:'8�����6۞�ps�g
�u�a��3g���^R�Խ��p��p�<k(���E��M�DQؐ�u��s��v�u�rkd��z��z��
��.Ζ{�kQ� Ӳz�0��E֦����f�:u�İ6��������/RӍ���њ�F��'\�jM�$G�f��9�m�0t*P[6N�Ҝ��U�O�Ҷ����.-��`�cF�v+�ۑ�	(<N3#���>>T�fe."^�nW0h5L��8��᝼X48�Np���zݬ�Cw�[u�\�f��-��hm���x�̈́*��&�9�����m�KYq�8&&��tu���K�T�Y�z��&^��7#uùZ]n�Y�v�����l�N�FT���j`�z�N�\#���mq�3׷d��*]�L��<�ҖlS�2��j7j����Q�JV���j�X����5NQy�S�W)X�*V��h�Dt=��5"�� b ik �N0�mc<�<�w8+Y�	�H{h�9�6�Z�e�3�;@+H�n�@<ڹ��C��z3�'D҅�ز�Ivyl�&�5��r�]�W�0� �](춉ދ�#m�[Uq�kH�q��
�(mpv^�ܱ,�;sR�2�U�k��Ж����fs�Z�����p��z	9.9�Z�,���ٶF�6Qd-�۴e��n8m����E[��R��(�;��8`�� P�(������B��lc@�9i��Ɉ��1 S��k�F�Ԋ6tWR�-˲�R�hVb��"�M��*P�,�8حt�uƹ�t~?{���?�=@\����M��Lΐ?G��D���}�zM
���^�A=tFb���P�ʡb��8�4���@ۈ��#m�� �r^�\h陧noniD�����7���6pq�,]��[��
y�s�c��x�+�Px�I�����϶�nx��o8�u̲����"亻D]D��M�����gbfD��r��q�N�9Q,�6�6
� [��F��[&�\`v+n#�����.��M�#�5�0�80:�{%��x��n��ċ�-��q�����7Y^�5i��@�\�>:��Y�U�P����m���r�K�Mrs�}�_c�c�k=<�;ʼ'A��.}&�j�{���}�Ptnu=}���6�ݝ(>��e@/df=�{i����m�9��4�������_/gM��@_{6�I f�� �8�M���,��l�=�V}���o8n�,�����l���G�rR������fnޥ`wۋy�3via����~�f�zA�u
t�$�9��/��wN�ɓ-}�(�f�[�����tH��Z��*䃧i�=ʎ]�S�73��{F�wP�n�r�c���{�/�q�(L&���/�H�,�$.祒FkY��}�fL�6;�mX}~�$���k5��]y���
W@p&� 1�#i��dL%TC�y$�Y���f��;^���`o�<lP����a�����2�� 3an� ^�mX�nΔｳ@{�&S��T�*A�r+���wvs�f��@�ϳA���gLٳ��{yGL��ę#j
Npݚ] W��X�uč�{��GI=��%aԌ4���9u7��l���L��f�cmɷ\�q��GV2�/�r�B�*R��1H] {�6Xǘ�����+�ul�X{�3dt꣟9%m����U�UI#��{�u#6�Y`��e_�U�tff��N�Ĺ/@}ݽbݝ(����p}� W��A�UlXo;�d�u���ۛ�!�HH'yq�n��32vK��� {����Fc��3�u����Ȁ���9)��`�p�w��X�f󚑯ei`o�yV�T���9P�{���m۶�M�65ma6��1^ۮ�fQ�W�%Ӹ$�QJ���+�m��9��� �nޙ��Y��`{1i��m��*A�r+����|yf���}���Čo1_���e7��(Q&8�Q9�����/��4p�3���z=��`	��5i2'�S�-L2Ps	�����3cvb)�>�۰�̃��d3$&EL�쁈.�+��ڡTL���`�������Bd�$·3`f�����32��~���<P��,��v�`�U�ba�!ĉ;c��8��E,H��቎��v��{���?k4�MPIr+�9���f���=���
�R͛��>����� i(�v ��ҙ30{�*�̌ǣ����+��_|Y�c�"�lR!8] g��B̌ǠL�/ͻwgJ���oi&�d�!9w$�_WMٶ�f����,+�J�}��Fw��q2��DȦHi���Gٻ�`s2Cr�(}�4�1�E��L��䗾vJfQ���?�O����a�3сf����4��q������5�0�89�n�ex��w��[Q�]qc�$�݇VGa�N&���m�W\��kB����1�Kq�6S˛�umg��^&�����cD�J�z�;�����w'q̆cceL�;�u*��kWf��Lq�n�;���t\�k������
յ�$gq��*����ݷ�����oU��v�qlѸ����@����������+ێJx5ˢ�yu���hk6����f�ui��ݥ̙뿷�-���d�L���_�o�4���6X�1�E������bo�tȡI0@���y��/�ٮt��n�>�w]��vt����C3��5a�I 7i��Oގ�/��{��ΏN��5���S�dM��'"���9�;P��(5��f�ߝ�ݭפwc��! ���n���Ҁ9�3k�bΛv7U�����~��hֆ�$n��;s����6�6�wg�V�����n{n�u���W�s��rP�p G�Nb�g�e���U�/ۻ|�0��p���=����q���L�SS2���z�3'K�	73g�ə&� +���]�:R �=�_��LG٦x8! �"B�r+$�~��p�wf�A�����1�+�U�R͈�Lh��s�
*�wf���԰3�/��9$��'���`��Y��0�����J����ͻ���۽ָn���Δ����J �AI�H�m)7(6���w��&����b��������]�'�r�$�vܜu�������.�� ��l�3�(���f"b^���w�ə$�34�<P��K����WUT/��/Q�!�J	���o�M(>͚?&N�7$�f�
���A,-)�
��Q�7����^����pٚ��R!8X}_U}�VwS@fFc���ݫ�'də.�(�3ڶ���荍�K����uX&L��ݫwgJ �ٳ@szqB�n_�]<����[�;�k\�Og�Y�+:3h{�g�|�O���{�f;n�gs@����`n��B����&�w7cuբ�x�Y���D1��m�pܛ�����6��̌Ǡ/��6�$�����6ʍD�jSR�����n�����vs��O ����a�)��rS���_V��V;��p��٥��HB�v��ȁ�>*>�'~��9箶&��I�F�qY$��nՈ7vV��ٳ@fFcЃ�kn��W������D7�u������ȁ�u���eC$1��IwmQ�!0�J���~���@�l��d�=2��۱�͈ �QQn[NXZ��6_�?���^��}��|�vt�fI2�s�GK��L92M�T́��@_ۻvs����I���Os�*BXm�G��2�1��v��S� _ٳ@�by���2�i(�H�Hڍ2s�f�ҁk�l��K����n���ɛN�D�����H~�.G)D�QDc3P�	v��>�6�9��x9���mћ ��۞]&7뫯'ckq:��h�{t�nè�����[n\�keŻ5�a�Yv�����qv��nT�����9$��.Ӻ]mrӏ8\���Ƹ��Jg!�]�b���=�^1ʚ������Z0���6�A�nnR��n	�[^�tu�[��΀?�~�~1�5;>��{�����W/�X<.R�aL���ȩ�����vu���l�a�S۵Ɣ���Sڿ�u��})��j'MI��D��|�Nk�VH=�Ͻϧ��������4��|���s�n侽2ｻv7wf�w/۳_���u뭉�

H�qX�~�� n��@��١�3�w77n���BA���s�W�[���$/n��&b���!����v3w�@"E.���q�J K�n� ̳윇�>����:P*����喬���X[޳[��]Ѷ�ӻ;5�l�T��]�]>�tGM�6���e�"F�K���Q���~V]�n�V������-{������\N6P�D̼'���=�ͻ�3 �1P����Nf;��9��ѡW~�Z��~\��^��3b�����s)f�*!Gb�"n�[�:P��SG32HI����ޞ�g�c��s��[��i��N���yz%��۳B|=����Jݵ`&dʪ�v=VU��摧�s��e�	��7^�w$�o?��W`o�t�����OV�)kP�mĊJ�@��m�U2E�$��]�x.O�<�	�i��0ʉğ(UUSwl+�*p����G�����Kwf�����ffHL�5��Tn�����;�K��M�pݚX���Fc���}�s�B� �-���I���L��	A�mn}�$�^��K$�I$�I$�8I$��rI$$���������ٙ�-�h�<���~CMP�HEQ�����N��џ�p-fTŅ�ŔfBx�x]�·���ͦζE><ѶS8��Qk�<�uR��؜Y$&5��;eX��)�Q�bh��s�<��9.@�5��}��n�sLy�8!s���ӁWc���7��8���(0(�^��9щ97�o��{�|�����W1T��p?
|i�[�Q]� N=�#�Q;�I^��Ы� �xv��ч��y��b���SW���y���R�Lй�3RL��̖��컰>�Ιn�u��q�r�ܜ꯫5�h;��� �}�K8��=�g�,q���$��r+:n�8q*���vi`�ɡ�3���ob�9�yR'���;/:�g���a�ڶ��n9�;\luܼi���] P������a��q�I>�����hg��5�ɜ>��k���(�������H��K"�;�uY�wy��f͚w�W�U +r��G>q2��<T�n�����vs�2~s�Oŀ{k?K1�%1��(��2L�>�ݷ`n��@�٠�̀HN�B!#�S��\P�.��[��<��N��C;ˢbo�n� ̙�_�f�^��zｻv�/a��ݹ���ƣ�r�v$^�u���K�M�J��x":�z|��������|�m=�K�!t�������w�ݺ����ܚX�OZ)Q#(nBqK��f�פ��{v�ݝ) _�f�d�H=�&�$��H�NEv��{��'��҇t̙���6i=�������Q%76�nr�iW��f���;���$f��d���_8Iգ�ΓaF����Ps۲������bV{��s�lk���_�_�� �(����&(�;�pݠa��~k��)5�)n�/���ݐ�k�dl`�V��l�:��]����t��rmw��p��*N�[GaH͌G[�?ț���'F+�W7;�:^s�lpl���nz���>p(���\bh�����G��J��M<9"��R�A�î�iƝ;p;��\��\sڋ���O���4<��nc��)��^C��8窝cn�8;bܶ���k6f[���ٚ��hOԔGl(���r�3=l�U�1P^�N�ץ�8�у]J�힭t�qû���?۽��}�E鼴�������v�[���m݁��� _���9�]lL�0#���#�=�rݜ��Ҁۆm+67^�9O�N����P*|��9��٥�swe�Ef��`�Y��
�n�@FI�%%%{�4���z��۰3vt���f�"F�nBZ�'
�� ���wv�nǪ�+���x�T��+��)�tY�:��͘n���8��N��yW��6��uc���R:�2�˻T>>�~�_��pܚX	w���{b�w0z�Sp!#mE'8f���W����t}K^I�ld�3��Q=�@_�:P}�����յ�F�C�&��+��we��Ʌ��ww�=�K ����jE>�}$�YnJ�z��ͽ |w���^Ǆ �3%��]dMS��Sn�罻w`>�����t�����-�x�����H�Ң)|�r�0���	���q�R
L�4�����.B�s��������n�����A�٥�{�.�;�]�����b��FEI7�HXP{ے�F�fΔ���'����Ҁ-n`l8�KCrԹ8P{6�{������G'�@�J
"�0!F'"P�!\�D���L���1�fl�nC��@�d����8�CeD�NB��n��f�`���`w�0�7s[ E$�6��|A�٥��^͖}� �wv�I�Լ��B�-�S!��R8S��j�ɉs��z�ѱ��[-����r��W��;�6�� �we��)�����8n�����ԊR"�7"����٥�@w�[��(=�4�
�se��Y#N)��,�o9E�f���]��;�XVj׿�O��<MX	&eͭ,�ݚ�d�@���}�	�? �N����]u�~f_fO�P��7�HX���ꪮ�&�w����٥�F���5'*�1#���u�ݑ*��bP�6��1^ۮ5���3����m�c2e�|_WX͝(�ջqnٳ��I��w|�(3ՓiGRR�B�"prup�ۼ��d�9��� {��@}�+Raût���(8�QI��[�~��;��e�v;�Ng��p��B���%')�Ľ|�/�vj��fN���a�2m���\P �ݼ�fdIh���TT��:P}��`f��@������2s�J	@�~/`�� X�8��&"��!���3��_��FM-�w<��[����)W�2�J�l��=W����rVȸlp�]��1�Kx�6���;��>m�h{�m�I[�p�8������n�ƕ�3��lF�!���U˶�u� ���ƴ�������{xܜ�Q˲񞺇��:z�v�e[m��ܖ�"�'��P���i�Ut�0 V������J�8��V�����?m����m�h�ң��Ywk����������n^�.�;WmBn�ۮwcfv���R��%:����������\�ƈ1!8�i��?������K �we�̘X5��i�5L S��\y����t��q��7gJ����pٺ��PI��
B�9��`{2ag;Oso�H�٥�z��Ї�rԹ8n�,�sy�=��JF?&I$�����ql�y�"H�)!`w���Y�zXPw۲��b�(f庇9�)w�C�#��ۮ��g;Fa�Z����ڴ�&��+z�׽��d��j'/�V��?@\��=�8s$�[����b|����x��y����[λ>�} ��*J���������vnɯ@	}��L�
��V[�7f�{������{����/�����c�U��pb�c�(vm�ݝ(_ٳ@A�aXQA��^�"��R��I�{�3d����n� �f�.����-���1����y��d�\\�zuu,n�=n�aV�(��l�ۈB̀*.f�i۬7b��mf��d�@��sn�_۵�?��b}MD���Q���]��o8�T�� �se��ɔ�`���'Q�P��݁�����c/�3!!��$��'^��.����������xX�=��(I�pq��s�7f�f��fV��o����R���s��r@�l�%F:Ʌ����8��,V}��Pf�i�EH�C6���"�ܼ���U�b�t�iAJ7m���M�������(O��pWs�ջ�e����8�������(;��EM7!�7��Ӝ�қ��� {}���Ʌ��Դ߄Q�!F'9�wmP�6Uɐ�nΔ{����Z��pS��$�XW����ٛ��V�����A�蒅�C�e�	Hz��U�TÏ8h���w��Y�KRCQ&�%��vn�,�K=����t� �٠=�b�H��rF]G%��]�z�����3�V�ٶ�vu�O��H�� �(�'Q�pwwyޠ�{j� ��ʯ�����Ƭ���@�fH.6�Rs������ 
��Kݝ6o�J�v��'�6����I8j)�H#{�K?%��6Rnb͜[�ٺ���1hH
�(����Yz+�=��`f���0}��`wαSƘ�I*4�,w4�U�y������4�'[��\~�����p=ޞ������7����{������w��Ϸ�ww'�?�� �:֥H� �A�P���
oؖ@���$T��:��]����<����㻶���]�|�/����JN͞�����3�E�|%:cDI�рzRq(���;O{{ 챈�!nx���X<�{�O�X`z�d����c|�T�����o����h��P�z��b��C�0�[��l����#��:��8)&��p	zF��NDv��n\&V�J�zzt��ǴR"	��m����鳷���
�pc�I#|H5a@AQM�0
a�^��{�N����v���o��s�3�)�����X+J���O�����k��{{��I��e��l   ���m&�J �ه[ �6��m�l    m� ;m�����Iɻ-*���p�x*���[]g��:��Z ��:1�n��p5�m�h���Mm����"Ke�2�ۍv�tΎ�΁[m���rhΑ����Ӏ��.˶�g�����]�m���!�2�+�r�(�a��Z�b{uedի�*E�qHiD���:��1�!��e�J�պ���שHt������T�����v\mB�/Ip��S�.�nS`�z �l�@ѫ\*���Uۗ͡HڍN�{4���n���j;4Y��dS8�^�U��&�f�j�1ݲw-g�����{m�MM����F.㳎�Jgn�҅#6惇t��i"��[f�;�6�]mfʹF�����68;1��:%��fѬ/!�*l�+lܑ�Ճ��s7>��!�V��awn�e܊t��{qm�S�"2s�.q�ݲ%��F�����^Lܫִܕ�R�	��Gv�����pp�ܾ�c	�u�^��l9s�5˫��raq&*�d1���j2�F�v�`,�I�=��Fv��K�;�>f�ݷ���ʽ�V����F��v�n�t1��r�jMO)�K�@Tڕ��tC�ϩ TVR[R:^kR��Iɰ�v��yܻj��k���k�n�q���u������u�ܓ�g���h#�� Q�5!���ng9f�[I���%�ru;,���@�	�TV1V�u]T8�UFð�:!�)���3�T$�mt�k2K�n��P��ʋ��*]��b�^e���N�P���A�=pR�.pM��VVV#N�Vhݨ
'l�/WT�J�����
R�iV�b�-��P)Ke+Nʫ�+Zx����V�ԑ�T릤��ѻe��$Q[(���i�K.�l�MN�m����+ �r��D!$��UQ萋���������@Q�j֫�0�X�ʩ����
 ��|�b��+� ��/dtoAڠ+:{`��� �#����@�y��*R�\��	u�D2�@+Z��$(��A�j�$q	�(Ty^qm�8`5�=��5�1��5�B]l�u�7��7pg��6z;_��!�>r�qѳv���1I=6�߂ݕ�����널Յm���m5An�y6z��F�����s�lxy�wv۟��v�tZR��hP���ݼ�t&�M�v��]���Ƃ����[�Y�»�yb�<�g^$�z��C0Z��'�{ZO�T5[��<��+̞�7k�=h�T�lNW�n���W$�S}��XTE(����@���`�l��32��+q���� L��2��^�>�l��2p�=����8f���3;�,�S���2M�*��p������ �{�������Q�A9�N�����z��5� ��Xq{2찣wpkg�MS���I9�$f�Z���&����������i���8����z�Xm���OD��^�<d���!�;qZ���ev��l�˪��nl�ٓ��K��۷��~ފ j����o�T9%4�nJV+��7viϾN[h�I.M5�<W[݁��tPw�/�_}IW�V��� AH1�Y��۝v���;���4�e���� �!�L;�݇$��LwE }�}�3'
fc��۰�b@����çxx���q��4�ZP��{�	n�;��!��U1*�'��W΍qM���Un��h9�f�oo3[qnߋ���C��KWrpݚX�n�A�}o�8("N}��I�j�
6�2JRDĉ�z{��w�̒J�~ފ �ܚwf��D���!�DL��n6R�q�W���k�W�{��~������,`͊!	����q^s�w���̹�e�7�p��5��	M�-8܎Ga%�d��ٳ@�ݝ)?�ۿX��ؠ��ݭ�#��S�$�b��Ƒ��h�nn� ջ���얒3�0Q��66�l���t$�X�2J(� :�Ԧ�ێ�պ
b��͸�]NJ��;�ߛ��F�]��}=��H@{1d��+
@f��P�%6�Ɠ���u�Pw}���Ʌ�/o�y���_�T�r ������v�n��G'O~�}�������*������EnBZ���̙��Wvw]�F���۟���_��w	����L~:�K�k �}*�á�<�;,���h��a�R�&$���ݫ_wa���Od�;�z��>�P�V��> �ڕ
��m(�-�����Þ8���q)��;�4n�\�=%T�GkYka��C��L������({sf�����w�T���5�ԩ��N7#�>�d�$�'swgI�;w���y�m���PGϣp,Ws�������n�*��N�u�Y$Pr��$�`{s7�(1f�nd�3�@�3���!�N5��7b�/s&��0���Ͼ	{f��M�#)��M(P���(�t!$)����F�[\���T8���t�a��%��C�<= �͍���srb)ɳ]v)��(���i���q�I�S�2`��[:c\�4pѨe=�
��9U�׷7F�;Z۫q���܇Um�E�z��K�ݬ�N��65r�=n(�K�k��gQ��\�W��K���t훎�ē[͢ۋ��v�ǈأ7	.�i5��p-!�k�x���u`X��ii5����~�� �J�����cgqV��R)��MI��&�<n�ml�	��ۏ 73����~%��g*�P�<�v�pՔ�	Ɔ�%��8��32LÇ�p۰�{��>�d�̓}B7�6�n*�|���l�3�~���7]��֙�c�g���y��):>i��+�ێ�k��8c�PZ�c� �<���m$��RH�o�X�<X�fs�b��`wیz��<L\��W�.ۣ=��ts�"�R�l��ҥ��N�髟Kr�rRQO���H��u��e������˹�f�{]l�"�ș����{6�~L���i��n;�\P���>;�G�����=�	�6��ۏ��������`f?8���Os�?$bjZq��q�?
O�f��H˾�U����@�/���iD�#����N���~�f��|���XD�{6$�'Bղ&�B �#����9��5o<���U��_*�j��i6�f�F��(�T���'Q����7���c�o�]����V�7��S�\&&�A��\���vl���C�>����P��<>0[A�F��1/@��@fG�?&A��/������FF
��0"�m��?T�%���缻�ޅ�^�}���&Q�9(�]�jG�T������_,ɺ��9��`sb�1(J�R+�o�o�}�wf�`�d��1��>W~��R>0��_!�K�TT;eW�v�5���L�!WuKpN4a8?G���v6���Ɣ��3�kU�7�,��}_P��9\ ��Rz��4�Bn+�o�n���L�wF�{ٷ`fGk�$��2P{5~o�6�$cq��ܜ�?~x@;�������|��{��^�u�r���7E������pǺ��Gvd�y�y���G@'�$���9]��w�}��$
���#e�D4'��	��27^����ْ�oM�;�I}�{.�����ws��ܹh����i���U֎��'h�8��kN!�uVxQ�d+���/}�@,�=S��g�l��7^�+�=��"���8�U�� �x@;�{.�̍נA{��dəӞ�Z���-*I��P��
;7���7^�I���͖U�"P~=��)T4�Rn�]�1�@�ɠ3#ć2ffI�ۛ� {?$�
��A�F�ӎ���̳gJ;������[��B�(�
P �(ѱH�	&�D��p$XX�H��F?L��F��0O��f�\�c\�l4���5�u����fcE�:<���Y �i���m�sZ�F\;ˬv�yn�죰�m�N��p[f�c����jU˹��Zۗ�<3�;m6�WY]^�>��v����+����m��@.J���ǒ�rq۫q[��WG#��p�9ewn�]Y��̒����y�8�[�����ְ��-�;���a��K��u�	�Ñ?�P�=��4:A��LjH[A ;v�^v��Û']m��-��خH�#����q�K8��6��]ա4�1��t����x@;��� �ƿ����ϳ�8RI���<ļ)�,n�۾fL������}�6c�+R?eiJ��P7��@�� 7_�� {}�@fC������j�&1�A�%8� �o�����@;��� �Ǻ�<��wC�5	V+��7^�{9�3�${}�����C
���ht���Q!P:I�b�Ř8v��iܚ
�d'�����
�����������sU�s}�,���h�B�mӍ79�3��Ԍ�����!��l<�8����>X�Nxrbzh!��Ny��˿���/�g:�IԨ�q�7�osg�c����g8c�V�=��M(ڌ������g��(;�uXu/n\�3�t�9J8���$罾�z��B�ޞ�P��t�S@n�36j�C��YG�͋�������=����F[�kd�[Wj�q�����F@[�$4��D�;�O���Py���4dx�p�nm؃�5t��8�4��v��K�_R�n� �����?k�-��ۺ�� P�b�6�0��g���;7�����`bb����������o_���<�ɵ�gW{�Y�^us�31�w���ٽWv��}UUSo��3�S��?��_��������4�������_���֮���_���t�a3��N�`5<��E��n�cI$�_�n��.�׈`�`A�a0LA�$�@-��@�&B�Hb00�9�ܩ�t4�8�p%���|�: b�<)$�)�������bc�0���)!:D������Rff� F�+͎��c#Dj ՠ$���%�K ��:I���4��/�]A��9UA�&�(01(ie!0�	R�31��N89-���<ੈ[۽��S6j�Y�&E�U����u^��T%>��psZ#�` �Ja;���m(�S���3eF�������t{v��m��6'�(��6��,tBJ8�F �w��;��N1x�`����L$Q�FM�7�
R)��@  Ѧ��A�a��К4``���	��A��L`l4&�A�`h6@OTS�� $M?�?��J���/�����T��R��G����A��\U
'����Pp�{�_L
�c��W-�$�۲�RZƧ�2���(XQ���pY��-�;1�P{E���P#MҌc����]�?�I�gӳ�����>��������r�iK � �m��{i�-m۳��+v{g�SԶǞ۱;Z���u<�]�����#�1���<����A�{�V�=�_}
�&TiFa��	"{gJ�L�^{v����F;�O�e�&�R�&#g�#����	:��v��Gec� �V2�Be7CQ9�X�u������ >��>J���/F�s' Іa)���_�kη�7���U{����:n���D��rX���
����r�3vhL�|��gr�B��9�ճ�7r����b:M�Z7)0m���̖(D��v�	*DE�o�~�x�;��s���X�ծ��:�q$Ԕ�ԌBe�W�6������[Y����~��;���H@�&(�s�w��@�nl�$����}�v���I�Dr�"FĜ,?q������f<���}�v�̒����1��"RCQ�FB���7^���Ws۽�in��@��b���w�a	X�`d��jZ
`�-6�3�sE��=�_س�$4u�����5 l�h.&�ppn�i�L�<0u��7�]Y۪S=�J[i	�t7R;kc�ڴX�8�>�q�v�O[�n��$�u�%An,�<z95�^�a�N�v�{ml��6c�9�;��\���b3�;vSUɹ�Ã&f�fɫq���Gv�G[6��]��6(N\��g�'QmHل��[��/j&������kw�^���~{����cX���S�-���7I�뗱��[����\P�47�ȊR�D�)����뻗Dl�7>R�N�e�����<�l&�c���[�?�����l��Q�������J�s��܌�|��/s�w¨
@UU#����Xl7�� jCd�v����ak�O�v���(g��n�r!B�%"���}�Wؽ� s3�k�;�4��rX�X�h���d�vv�7������K�=�*�8�T$�����Q��n&a
�^�S��:��gp�8��nnT��1m�ۜr��*K���;�(JR���M��͚X=�=�	���L�8��3n�o;�;�
A93fkw*�>�����G��p~��2�)�kM� �n0a�c�C�]�z��:��w����XfΔ��)q��ݹ	j�N���@w3��Q_sf����d��ס��!'J	��`���ݽ�����7=�@/?���,�&��n��$�@��i`��`yv�@�۞�p
�z�YF���&!Q#G5$u�xW<۪k�${ �۵�C�$E��\-H:n��BPiIN�� 7se���Pn{9� ���,5*�Y�.�(R"�Ws���t�syۚ�����ʢL�Z���IL�2P&�����������r��%�0���fvjȰ��SB�&]���*�"T�I���~�]���`Q���A�9���p�D/|��E',��w�6�92|�� >��۱�ӥ rI�r�j}��s�C�y�$w^�X��粖�U�ct	�jW���ۇv��~���*$܄��o������p�����v���7���j�$M����t�݈>͝>�}̊{ئ���!ml�2�������٥�[��=�p�9�5mc7M�"))��s�{����g8������H� �kKU����ȝ�U�
�9���;�d�h~j߽vK�B�(R!�v��k��sٝ�w^�u{u�'�U^�[i�|ʅ q"�1�\�'�c�um�n�r]���m�|��l�9�oi�.��1�����P�Lǀ���>͝(�ۑ����� g��k��Rͤ
�Q����_�եc�a�Ƞ}� o�̻�7&��~�Ǆ�
A����~xr���;ٵ% +�v61.�D��Wc� n�p�9�;�4� :�����Q>�&���}������@|�̊ ��!��K2�2!�(%R��|<}���g�5�off�5�	p�j��2iLݵۤz˪͇=lb'6ͱ�^d���K\뫭�m��B6��A2t��7M8�8�Mv�=�o�KjG3[�pW=-v�&*^���&M�IKÞwd=��=A�=v�"����O �4F�!y�^G��ا=u����)��s)��{E��[�ہ0v��h۠�:��� �yƮ�9e)F�㍨%���
�
��b�J+�Jm� ��;���}�f���nnq���g�$c�;��n�#����\	4h��xI�ݟ$�f�I�q�7��� յ��:T�mA�iIC�(�svo���ؐ=��.��vt��Á_�f�����H�m����p�>e٬�3������@c�>bw2�3.�S��32fg���wO�̖/y@/�R�ϕ*�LMA8��3VΔ�g��lA����{.��d����;�NAp�re�r�8[��v��d�Cvz�Q�=��5��ɹ��9�h�P����9�f��+��Mc�����ɥ�s��X£%$܄�N偯������\2l�����a<Pnn� ��{Dl�)
�b��&nn��nΔ��\A��4C��,y��ò�P�(�*��oԑ[���XP{we���R���fp�YZ�5M�"�0��(_ّ4&lf<�ٛ�`,��K>�G�6�
H�P�IJ��
�����l�T�h��R�m})S:JJ�]���$n�".7s�}�w_x�rn�f��6H'��j$��ReIR7#)&��!��ݻ���Ҁ>�ɣ���� _tA�ߚ���&�8n�,��9~�� X��?C�A�W�t���5�C�� �@�"����P�Gv�}o�C&f����M~��I�y�=�`c�Ɂe'Q�N���`b���G�9��zX;����8�܄������@�gdۙ�_��� }���"tn��6�lG	�\9�'m6�FzZ���y��n�!MSuB��]컣1T�X����k٥�w3%W��YA��P̬3'�t��99�3viK��=��@-|ǐ/��.�$Μn}�t�7�(m8��X�n�(&?yX$̙�̻�ݭ(����T�T��H������]F{2�n�9_���@��*�y��� r�ݟK>Hj)�����4SVI��۰'7kK�|��y���c8�s��vz|��2�^nؼKE�=��T�fqp���v�f��4C��o�Ϳn�>Δ[��������RI2_�.�0��Qϒ�Q�N�{e�E%�(�{3��v�����
�5�E9Cr��pY�����f�K ��%���6P��R5`{}�v����p�ɠ��:d�lf<K�n,6XxgQ.3v�;jJ@��&���������V��l BC	X����0�2��0��LL�)30����E�?��������M�z���o?wvfr�I$I#̻��I$�������o��n��xffD(WMUD�@i @��ҏi0��=<�1Lj�����K)A��G��6q'��Z�:Ӂ�L:GtJ��vo�f85�5�;0��lL�"$�fa���C�51�|33jn�����i��uޒ�l�4�b�ox�v'^$�D������ ��Ѩ�ߍs2���G;�s�4�Ul��J��f�:�LXa��2�A�d���c�'�(�5�KJ��]�u�1�S��~sWoq�L$r�N%�s��	)���D��2s�s��%)g�Y�`"sr��2� 0�1���2L�ܤ�l"ׁ�֓�z�J7C%'��8�[���t$m<��:$|S�l��&6�z��zb	�l�8�T��ˍ%--4	ю	M]��Y�&�c�$h�s����,3���A�n��^>�u�ް�l�|���v�?<���v��h:�bіc��-sORtfa�iֲ�M����#O�s۟x8��6��   6ۃi6�n�[�� q���l6��f�l  2 � ���]�OV3�2�B���%��7c=�P.�^�k$<r��9a;D�8��Z�g�-�8b3�����,9�벉���'��Y�M�S=�
��C��c�X9ц����-��M�y���jrg.�8�l��뱺1]N<�������Ӻ�b퍎�t�j�o;�9��nګ�&�E'�4��̹�oA���֍�����l�W k��pr�mY2t�&����
�Xî*w,p�Qz�������6t��mFxU�s�;���� ۓ[�Q%s«v�zs���I�v��4G]�m�j�y��>*��y�.̯�6n���҇V�e�e��ű%H:��Ed����c���W���_B޳8�*��ec/VHAQ]��Q8�Lr�KSc�z�aę��z�ҜX������:��s��[�%�ZU۔S��T���)�{sq�`,!���j�*�u<�c5=�'S����	����3�8.��Eӯ^Yb"��GD��i�7n�K��EC�A�Y��6�iJ�;���@0��:m�@�mV���x�;��ٺ���3��u/p�m*���8�G�l�� �P�r��\,��] 7
t��Y{iN�vYS���gI��^1�4z�<:튃�֞w�D8� �Е�v�j�Q�h[\i/n[֋�a6�PnaAt&�)-�7M��um�B���)��b4Ù$dge^k��݂����"�h��JF0J�(��#;�����e�f��@ݶ�6Z��ȷ�ghs�tv`gf1��j�1,��J�*��@��S"�V�Xm\�R�[�m�Y����ke��ZT̮�<=@ig5zvV�(��N0Z�m�:p��7F*y��t��!\ӥ�s�����6���ɳU*��-.�(UP����0m�+���Z��,ݚ���=8'0Gj)�%��/jz�C���P��iP^�1|M���	P��"�)Q`fF�)Ief�*�R@��H*�����6 v&���|G�������o������5�)mr��]���ۏf�hz���N�hI�_��<|�Kn�a朮���㓏��?nwʝzu�d�����'�j�r� ʀ��@��IJq���o��Ŷ���b�w �n�̯��k8A3�۔�\q�6Z;S��<(��j�c���U�����]��#̖�������y�g9�@\Du��t�h��ۗ��z��7n��^�.&�
,Kv�7k��������}���=<�Ż<�ss[R;��,��$$^��l����*=����lU��#k�e��'��3��@c�� W��fI+f��@g��n���$�
D]ۓ�V�� ��2�ݝ(�4330}����@�HܔК�;�͜���K �%�H���&��$�#���i��wvi`{K�Tb�P*��;�����|��JDl��6I9��q"5f(۞˰3vt�?��vD9�$�y�e8����8sv��c���a��������N$u�8�ЪR��,�A�2һ�$����'�fe�vΜ�2�3vh�f�TB��R��H)�n���Y�2C&\�:d��%�&g����/}�_:s<���T�>�����I������J@��h��_u������f�(z[P�&7B�33%���P(���p
��٥�Z�UUR*�,ۺ���y�(����c���w|y�{'��@{��`~����!�7AZ��!���۪2B�sf�۳�X;N�<��mu�����R��%F܁���O|>?}�wvt��dO2Vᯛ�@n�'����.&6������4�Ԑg�_ ��T��=��_UW��m&|�
��{�y�g~}�U�y�l�۞�N"y
K�;��*��y��_u�^~}SK�9��Tq!�	�����א>�v6��(9	&^�̞�o�6�/�j��F�g�7�7f�q#��,^�G|m��F4܀��#gYrX�ϋ�4v9`����ڱ����,�~w{D��6AԊ r_(ݚo��pw������sn�\��
!?)%D�"d�ｳ\��$�|ǐ/�6�-󶴤̒ [����L���e�&�l|Ǔ]�w6�����<P{:U�F��5T�#r2�j�/�{}ޒQ��Ҁ=���~3�݉��U)fI���&����%�x�=\#L��M�p���ΔS��Ђ��y�=�`|φ����D���]�)��E��Tlq�M�<�Y���u�lGQK��X�q��]�J�f�X����=�ɒk7v���7P��(��	j\�Vb��fI;�n�݁���ہ�ʚ�2d��.�)�i�'�T�X���
ݚY�P8����Y'�V�I�;�k��l�ڈ�'8q%����Nfz\H��P���g8UU�-�[%7R*��!`��퉠8[� }��݃�v֔��6${Z��MX��4}����_�?�G:��s���U<��tgDrz�έU���܆��qaog� :՞�ad�Wg\.X;��s����h�v���4�ݙ���ʎ���ƹaW�9j��L�ԋ��ۣ�����U=F�_mڨ��1O\w':��oa�*�[���츅�"7@6�jh�j����(u%ηktFv2���%��/}�NI�v�Z��6�v�@B�X����[}�p��n$�ف�p���ۍ������u���R`$�nӍ�Wm3�).���*Dl������>�̻?l�I�ۙK�p�P��!'�7#MX��\��4����VIՃ��H�~!xx$��&SQ&�8I���������s��o�.�����3J""`����۱z�)f	/}��U��K �t��!*q�܄�f������f�������)Y$}@UUg�e�m��B��z8�:�ۊ��;��"�.�p�"�Y;.���:}��YuƩ��SHՁ����8n�,w=t8�:�(I�wH["��e��$k{��=��}s�Η�8*����E�M@�7���A��	|=wu`u5@��W���k��[P��S�!�h.w=b�'�f(~@ϳv�Ύ�(<�ͥJTJ�.D��!�3@���vnΔ��J��^b)�>q��j��y�*�f���=�m�$�Y�s��<�J6�N!y������[lpt�.�ܹ�`�v����REnJT��Q*ns�f����}����(I�w7�#R(�� �	DDL�w/=�j��s_��{�e�3IҀ+�3u>r ܄bd����R��}��]X~�;T=a?I;��DH4�N � `@�?}���|��~�.�;�~��{K2�bn�j�7RE`s���pͩ�����ŞP(�o��G*:��p'8f�,(�k�u`b��9���Ԇx��-B�ATA�R#G>ni� q�q��t[v�N7���j{W�~8x~�r:jB��wn�Y� �7����4����WQ�4�D8�� ո��N�eP�:P�<����2:�w��>q��j��n~� Ś��9�۫�w1#�V�-`9�Q���9�d�;_�P��@��H/�x���d�(������P�k5���3m��8�(�T#��wv��������Ȼ�ݥE;�d��mU���k��s؝�}z@�`��le$콶�]Y%^��D[ۭ�^�=���پ1�5�,��4ݎ�b@�Y���\�ɇ��u`�[�):lT6T���Q���� �7iP�m* ���32׀��L���M��Rs���o�/��]�$��8�}��׸�:M�$�r8�4�X�ܕ@�"@��e�	���T>;����u)ȉ���\Ԩ�w6���T��J�_�S7�Xɵ�o�:~���R9&z0e��4��\V��nM�SZ[���k�cv{��d+�\�մ�=wiy�X:;	.�n�Lc��n����Mv �眝�-��-��^۬�m�5un;X{V�����m�H��v�ư�'s �g+vv�B7��~S��3R\7v����*��Ҡi��II\]�L��TEՔZ����j�t>.N2�ˬ:�z�Ͻ��=�Ҏ�FՉ����6乽t�^v����g�#��v�u�2%�\+�����߯��?���ͥ@_ض����|��ltH�!h�!P��m�p����X�$��z��� �=��|��}��N ���D<ʠG��T��z$�L�����u�O�Yԏ^��Q!��Q��I9�p�s9�+��ua��_;��I�D�_�)��v=��p
����u`gsn��Wq�9��e�JCpt�!Y�dnܽN��u���uUt�s���;F�s��'�;R�eI#��R��-Zm���ͺ�3��V,�N~��7��T���P�����[9W���+���H� �X�M9�T��2� 5YX�&#�8+�����z�d�G�b@���˿����_�5D������!u)ȉ��~�(�s9�j�,��ut�]X]=�#'�I&A�"�k!&d��������f�,{��+	�D��r�;�ͪT}�J��3�@W�ܻ�V��~�E j�42�&�:��L�w=vN6bny�Ԏ�����n�0�xߞ������/X��"]�J�F�WSP}� �*��n�Xs3>�Q(pj2;�F�\�^�2Ձ��T�}�Ԫ�$�3���eDA�t��M��=�V�8{v���{�|���}[� 3m�T�A����������l7@t�T<4	�AN�^��BYH �dC��胂��ٲ�v�}�.F����ξѱx�;���U�m"����2�����jH"!��c���!ç\L0�ނ5��٭���d	!�.Q��09�M��!$2�kC1A<H$�h*�q	"�8�S��3C�#5��0t�t$�sw}��x��M��=��s��@	Sc�{������qt�6S�A@P��@Pt<��O{��N_� 9�'�Հs�p�p��TLM��i�p��*~ͥ@�D�&I��ۗ`k�-�H�GBr�;��\���~Ί��۾w7'iP#>�w�	��;R��d�ل��͹�=v�n{T�m�Ve��sط*pr�]��d�өNDH�� 7��~�2��f�*ff@g۴�:�#�⨜���=����ߪ�G��Y!�@gآ@�zpIO.�L�D݁�ݥ@o���\$��۱%����
���Lq��RU��߶+T��I��˰�z��/��L��Δ&d2HI��O�@���9.�����
`�D�+ ��P#�$�-����W@o�.�}�=R,��ER:t���C 7
[6�"@�תw'�\��ru�)U��C���4�JnH�(���{۷WQ#}�u`�8[�aY$l@鉵��n��ݥK�	�;;iPڶ$�~��=B�
H���4��d�F�pY��R�y�&��=<mX�ԩ }�}�WQ�u)ȉ��~UZ<�gۻj���iPy�Vb�T�^�ЁI�NIR����� =��V��uu�a޽��cv��Q�~U%BaO�Qӥ;a6B��??,�kY�N�jw�G%����T8��m6y��B�i�N�ݳΨpGV�s�� �U�-=���)����(��m3�.;z��Y6�9��P���R(3v�R�jL�˧��f���#<�v8��Tm�
9���M��v@'2lmN�<˺�.Z�<��$񕌍��1��u���pp�W;��`�p��ⱈ�l�u�J6�n�$%��18�-E�a�ԯ
=U@N��̡���������m�U��t%��~@>1�*�Ĺ��8,���a2����GO1��}��T��M@��^�]��n��B|�Pn$IVo��� ���ng8xݺ� ���m"*��ڈ�R��ps38o^�ݻ��}�8��yQ8≪��ʍ���y�=�۫}�-�� �w
�#��'"�$I��n�] }�����wVs�wshEҨ:e	�ܢ�M�]�z�Ͳ]�i;/l.�@cɣPAvݨu�]u�M��u )IcNU�o����9��ZX���=$����)-_o�U�#Q� re��u̻��o���G�$B����*I�bh�s{�����P#s�J��������$�B�����+�{۶��2I;���Z�wD�f`��!�9�<M+d� ��� ;s�P3
=�~�A��VS��(��q*p�7=��+̉z��v��� 1��~��)�u����0��cH:�:���]�a��yԱ�Q�Զ���n��*�̏.<��<��ؐ3ٻv���&I[�n~��:�P������$r7`gL���d�N�ŝ<P��T/2'S329�D!)��Q%�	;�O����~�×�p�����F�>� ������2�ϫB"j�3$2RI��:� }������{:�t�}�WB�m�C����r�+��e��SK�7��Vg�����ў{��b��V)n{lmV)�t#���v��1МEF�SRS�S�GaFwۼ��텁�ͺN��� =�<�$�p"[Q����<o�TA�=�� �v$��>�Y&w��D�C�����y�Z�vuR�̈���eX����nn��D���J$���/���C�}��X���??&f�33s7�2_�!��K�R@rT���%%XB��ۂ���X�1�TQ4�ʐ��݁�{���̑��j��oR�̉@}�?��{����G.K�wk��N=y���۝NWj��In���pf�X:�~zo�[�˭Q�^��Ӵ�۫ �y�H=\��8��:���$r9V�6���3���8P{۷V^7۵9�A2K�DR��bA��.�d�0����},Y �=�D�XQ�H%%6䁁<��{�ՠ>��T��J��g{b f~V�$�r�6�i����t� ɷ��T=�@z�ܻ����������}���ߊ�Q때k��j�wm��N�ݺ��i���t�N�nΝ�;u�0����N_�7��:���"�mYp��nZ�n`�j��)T�[	u��9���Sj��Y���kF��8Ƣ8��;��6�9�.M7�]�@%>�9���m�b�!����NX7U[��kt�NzAw���ٻQ���Zwir��꨻��*a5�cؖPBS�s�	�w�ߏ����k�}9��X�g6}N��v����M�s��6.ȧ��ۮ�b:�vy�)ng�7/mi��&���J��ȐG�����d�̾p��R�;���f0�.�6�@g�'�$�]��>���7���fҢң��)�l�R9�3���r��f��(7ۗV�����/�(�e�S7a�4G���H�6� �}�T(�����$yxj���r2ܪwٶ�1�3bA��n��wiP�C��]Bi0B�8Tm��0��� ����blG����m��	�j��e�����V�E�$��7'7���)g��*�!o}�V*��5'͹%:vm{6���vIX̩���Ԩ�r���>�"$����� �N伧��x��{��P�����32N^�%�;ٷ`��>���H3L=33?{6���������5?���;w��L��w�w�V�lH��߾{z_��߽�V~��[⑂�bjJn�E�V{)�<7�c�P�<ݛGhݳ=����{�}����H�n��ٿ��+�w]���]ew�(�L��+U)&��D)9�+�r"@��ԫ]�{���e���&����u���G�� ��.����2#I]��$�H�(���<By�]�y���+��5�Q��Y�unT�%&�%w\ ��$���vϻ��2I&�L�&Q���V:܎2�3*y�o��v����tX{6��>�"@��;��"!�0Ź��:�����M��l���4g��q� n�������+��h�쭰���ݿG���vZ^���=�8o3����	AI�Q%@���<�m��`UP 2_u�O���p�X�<��A�s}���q��iH<�_�,���@߽�vS���n��{Ϝ���*F�!�F�+��ꯍ�c�݈��d݊��J�����0��	|�˓2I��ͨ�+��
:GR���d�)9��f���u`�8o���z<Z^�N8�!�
�ȢV��x��7tcm�{mF�x-��v�f{W'G=��ۉ#��H�feՅ��""��{�ʪ+����x'1-~%8"(!��R�>k�@g�컧s�פ�f*T*���F�Т�s3y�;�5�&L^fR�����GŌ:���m�79�;�5X�˫%�c�V�f���jD|�@�	�`gL˫ ��o��Ȼ=��?�أ<�����2Hm��mF�RI&�߿/3g�ᙙ����th�R��y�uy��*�=���AiL��0���`��H�Q9�]I����H�`łfL��3��n����#	x��A��n49�rٛC6a�2�l�#	!�T�6��db�f�3M�"tO��(�����������d+��Q�7=���m��(Ñ<wպ1��f�z-.��ζa
@ٵ'�`��0Iav��D�X�u���H ��С�1���=�nBe04bvn�1<��1���/�(O��А��P���8�b;v!�	�����+UERSDzZ�DG���J�BR�q/e� F�YTn()��M(����6Y�$�`�Z��S`$�.���A�a?[(�!:
�()�����wk}vzq��=�jv�. �*���Q�������O�[���d+����B���J��`1�TΑ^�O��Ӭ����:6�  �����zS]6 #m��v��c��3�m�܀  �`�� u�l]x[yG"'����������9vu;�j���u�$�S����{|�ݛu=��@]]�s���Q�	��=��_}b��`Z���T�*
��!���Z����
#�+m���7/I�Fغ:����#����=0=Zݤ��'luζ�s�,n��rm�;�����lti{�e�FY�mT�Ӷ�!�-�5���-۳��h�;I�t��۷`�g�s�͍��xxہ�l���4۔�ˮ*��cB��@�S.MC�UoI�H�=�����»/.YQ����۳\��a�nļ�nv��콝�Ps�ss�m�禫ջ �(��c��CVt��*hW��v��eE�`����U�)��$J��)�g�UU� �n�R���DN)V���še�ۧ�O�`���L��۪���G���=�/5��N�s�� ۬��cr��V�n�\[�C ds��]�̀):�(��g�0�h��&ٛ����2Ô�b��="�0�:��K�۷8���d��=����5Nkf����[�3-��n���[<�����m���V�ff۵h�v���v�b�n��we��)чl5/*�/JiX��ӭ�v��W@s�`�Z��d�F�ݦ5 � �Tb(�\C�z�č����ʗl�l\	@>��WE�t�n�ڜ�'Q�
m�h�<�RyrL�v�����DM���i�:tr��g��)��*�*� 9Gv��T�
t�uu�U@�ŝƨ���6�-p�H���;l�W3��`�+eKE�H����6��9Y���Ũ^����~�-���eek�F\V�J"UX�l�$N�V�U]�c�lT��T�,���E���[ J�Į� !�-��6�At���nhЂjv��Lt\��Hn�o��i 8�$Pl���� �l��vճ��n&�e������| �#j��&��Wk��&!��AM ����⡂z mYuB�]��\���oy��}�ψ����> �~4s�L�n��;`���],����tt��f�)�v�5�qAv�ٷō�]'!O�qR��rGC��(d\Z�.�t�p竷m4⌔`(��q�5��`�ҍ7�!��:��z�;V�[F���w�V��x9r���ewۙx6gcnR�熻C�����l7���6�򵬦|<��M�Iʜ��h�m��d6ܷ�랻
K���`�����o���}��v�(ݘm���=����/�̡��fڎ��9�����w}������J�������7k#�t32���Y�&�:h�QBF���� �=ԭ32��(+=�%}�6�� ��(4dI��Oq���<���*���}��37�(
�mb�M����H8�+��u`�|�Q���p
����V��n��R�4�BP6�nG v�f��r;���̥T�g�c�><���g.�n���Hrs�<�������\}��Ÿs>d�.�ÚY���J�RO�������F��}�� g��5�c�ҡ��\�纯�_�UW����>T�'	L{���C�����ȫ���H�{.��ӝ�'(�8�e��y�"^�>�[*�3���e�=�@��f�h��HF�\�O��� ��ڰ3���I?ۻj�F{u�ɒ"P�(H݁�37�<�U��X3��]ŹP�
T��P�q�jn1�8=�d�un�v�e��NѸ��:I�;W���T��6IB���F㚬(�f]X��}T���p[X��Ғ�(䐑��
��J�&ffȀܘ�;ٛj��Gy_Ա�@
þ?Y	Qہ�I���Ϸ���~y�]_��Ё�~� �+��>��{��r�����9�n��A8BnH*;��wn��F�Ђ��)P~m�lH�>�@��J��s�<�j�9�˫��8���ށS=�"�@W��@x�S҃ɷ��vO�]�]-2`������H��}UV�P��IM�`w��VZTgq�7ٙ��7�+�9�͔5#"M��1j�36'�!>�3n��c��~��T��(�(pl�(�M�����Ǻ�*�����̺�<���|W�%!��P�� �S�Y�AܙX���~�ٯ��)0޿�ߪ����
"[N9$�8��̕`W�}��{�����p��W@{ۉj8@q?�xtU/\;�\��<^H��T��&�鈜��Dv]	��^��jT��M�d�7u� �k�����pk�V=�X�Y����Q�%:�N#}���&fIޟ�=�@{��T��U�W���e`�R��ܾ�{���}�V��kWs9wb�@�	 �m�`w����
=�� �w���{��9�͔5N��H�iX�lH&fl���`/�7^����9W����+�c	~w��6���s�����D!4��� `q�$n�t,��gC��HӞ�`��Eq�ӹ��]s�h�6���z���S��r��vCK�a+�F\�z�l��E��eruͽ�:��Q
�F��qۇwFL��Xu��6�y�.����q�.�A�3u�\A���;q���}����T�i��`6W*v��N�k!Ҽ�����m�ɳ�s�F�Z�c��{��{���?r���;��I�GE3p�e��D%��Ay<��u�ۓ�K+���uv�_�[����fm؃�נ=��)P�dH��+�tJ���]�uU���&n�=�Ԩ�t{�$-���w�;�f�k[�o�(�(�3ض��=�p��;��{����G�y�nm�*P�J�>݉���y�6����;6���vR��*7$�IG`{߱o8|�U���[,�� �j�iBM���tX6�r��b�&N��D���gu�����6$���*r�Ns�|�U�Iwr����� ��3�(+۱�H����Ȭ�r���U]}ﾪ���5����V�����,�=�(�!@�@�L��ڰ��/>̻57�#��{��Y@s�M�(dM�E�;�g���=�`{��V�9@�ms(�dJ����D̼��`/z7^��d̳�֬�ؐ.��vn��N�� ��.:�9b�k�sgŲ]�3)��ڀ�8#V���jvV�,��!E(�(�=�6��9�s������[j�޼ݫ�*R��!R�R]pٮq*=ܼ� :{5��mՁκ�Q)T�F��(�${���G������?P�����r�;��C;v�������ﮮ�{��x�c�AB��*r�u9���M {}��{�I�#���x��~�� |��Q�`{}�V�9Ď���p��.���t��.9'����+\*��F��C��}M�n�í�'�Q�����W =�p^f]�}���-@gd�@��hA/L��@{���3�{���� ��넞�ú�$�E��s������l�@�� ^�f]���_�QHI!�$�)%��
���=�$��}����~��U�xw�BD�Z{T]$�_���O�y�����܍NՀ{���.�>�٠��g�����WF�����& [&�.$����L�q������=��q�����^�d]<��LJ��1`ggu����f���}����׽n��Y�BQH�P۔'9����o��W?�lՙ�|�pΎ]R�H1�RK߷K� �V"���w���`���"��N��4��ؐ>Y�e�ۻ4�����$CQ(8�=�sy�śQ@��z�p����ɛ̒��K��$�D�pqWU{�%��~*Ȣ@��չ"�[Sk���J���͎B���n�2��#�F͜�:;��6l�]\Ku��&qَ�xzNޛ��F9���NƎ�n�ss<p����v��鍍8nؒGm�P]1ʩ�r�&��`�Kk�����^Cd�E���.:�_�u���I��f�\v(�v�ъ8܇I���T�V;��F9gkY��|�<al�ڷ:�!/�(P�z_8
0�Ȥ����w���e\�N����n�5ɶ��h��y�uA	$��s��_�]���¬�� �����+�EI�I�)�r�� �q�;��s�un�7�+6�ur@T��E�����K��[����k�;��X{ν�J_HA��:J;�>vo}`y��(�N�\}>}�]t��B�MDnP�� �����K���"�:�wz{9�H�-�0�h����=�c�ݝ\�����n$��1�	�j����:�p����k�X�Vq�rS���w��� s�p�}n�qfc�=��MS{	̏$<�j�=��>&fe�&B�! D�2(���::RfI�d���}ݗ`c�lP��+�2tfb�{A"I��t�(�ٿ��:�7]��=0�wk���"PT�m��8Q�i��;�0��'��ϳ}��G����*)P�d�G#��<�L���lP���/���lP����ؕ��=H�)����n�t:�1m��,v�����a۱�n�{���71��/��I>ٯm��m�,�i]0��a`wν��H�cq�t(�o�y�ۮ���a`Q�c�{��`P���m�������y�l�s�.~�nH$�HYI�"�6����������}��������ܚ�VhՎb_a��\@8j����!����
���@RGà�'�@��P��;MD�IWZH�h�7��������zQ���o#�{GI�<|]{<�ˀ���}<�s�(@�e���B>k�@���9�N�p�:������{������+��MSQ�PbA-gAu<; )7�c� 2_������ N=i���z���<��8�׭�ü ���Ff�Ёo��� ��D�SOPC���l�T<��P�A�&�^�	 b�R��hmM"i133c$̚�JcA��}�����{^�T
' �~��g]����}�]A���j�!
R�;��~��K ��f��,۰�L�?�;�����0��%&�r|�%��ﳜ(:���o���˵��!����	N�En�;*���jSۋt����f�m[�5� �j#"�F��Y��s�#�w��=�L?q��D�ޢ��)�:m��,���(�N~Ȑ>�=�`k��=R�I�G#��`ss.��� �����Y����Jͫ�**m�T���b=� g��`|��a���͉#C�	٭��Nm�1x�Et}�w�zYio]{�)}!��(��f�8w�{����t�}� k^s�;�<:��0�G^1۫�gv3�qm!D֭�.W6-�����n�D6Ȝ @�@4�&�z����	��ab���jp�{6�3��\�1D�*�vI�ri���'3�j�^����n�tD�ܤ���D!*�{p��9.g��`O�۱f;�c6���ꉯ0dE���5$vO�)/g����|���
$���_|�������s�un�9��X��P�ߞ��_�׼Y�
G �0 1���r?a�r����+y��{�V��Q�n�j�S�3E�[����Ѻ�˳i���k������ʐ�����Om��.8�DV�ݸ�Μ7dՋ<uw�04냣J��*�����@䫎\z얂\v��!�`ŷW[�S>�We=��Q�����r��ln���<V��EY]�[�WiY-Y�6�v9:��0��&#rv�v�
���$�,<�`wKN4Z!s!D_�����8�
9e!Sp��wL�-�K�8ۑ�oGck<Aml`v�rv�f{W'N@��S2G#�G�I��r|l���P��}��[����+6�ܩH�U(�c��Y�*���g�}��	՛�`��隯�$w���q��QY'~��������G'�'Jy�� z�`���)79��~5�ט���P�UU�=����?�B�E���b�:�X���9�3]��{[����'"�"���s��΃`��%Cu=q�d�{y{o��}�q�F�k� ��y������lr��7^)767�j$Z�ȣB5g��~������}U"�*��Q3��L��?��@oޞױ>#I�s���� �m�HG9�ٮ��b��ء�{}���0oF�� �#�r8�I�j6��3B���o8OcOw��7�+6��*j8�|\��1f��I2�ۺW�y�oE�{�zp�L�o���\~�jm<��z�uHz붗��Iv�{P��{k�v���)��Y��}�m�Yf�wy(�����3b���k��z0�3��4>E9N����3_ ��`{�{��sUUW����%�wyO31@��gJ{���ek��L��'��
�+2�~�T��� �T$�o����;������/f��"Q�ڔ�rr(3�p�fw�y<�t��z�n������Q�����p����5����Y�D^��$�LDIH��h)�4�=��э����7K�4n:�l�qk������<cI�"r����;�@/�ͱ��}u�м�u�@��I%�;�m�^�mL=�e؇�����Y��.��h ��3=���z����[w\��Wܯa��n8J]`���]��s��_��*���T(d�&�=�P~U=3���_�� ���i�U.���m���Hf�ݯ){۲���e6�I��`�!�G��b6�ƫ�D�1�s��{s\W&�k;��t�D6�1FI���C(���:?�c�%s�������{�����$�i�cwI/��/{�u���h��>� V{55���)#v3���\�o��*�.�ހwN�a߽���(YI�s�����_{�[�}�ǜ537�7���'��%<(K2G#�K�w�(gNl�{��\�;��Ǣ|�N	����9�����"L�`Y��1�5&R�[��-��7�}�V�e��\a�3�	&�;�*#�����F��aͮ��M���h#N�k��b�O�y���{'<��5��wSۍ�2�a�N3˲�7Qtۍ� �9^�_�&��$ۊk�z2f��٠��-Ü^ɤ��W/f]�a�*,����˵7+$��gt�zː�Y�z0e�vh����]��m]���Ѳ�d�ˇEP� ;Wn�B���u���xl�vi${mֹ�o����������W7��\����Ur��zP�h��Q97�%��~�/�a��\���ssg�C��(�b8�-8]^w}־��R�L}����f�w�V��d�q��X������9���s3}�~~�b�6�r����J��m�3��ݔ>������)����V��ED v�Fv��θ_dw��nμ-yXu[��<�������ަ�{6�owvҿ����G�ȗg��o[�����=���4(`,3Ĕ	S�SzPLU=���h!T32I'L�7�=��,��zW�g�����$N�BH�rIu�̕\��~=�3o��ﾱ��-8 L�$BQn�����o�w}v9��]<Y�cH�-�%K������X�{`��]���d�<wt���܎C��Z��i�$T8�3;�pY;���
.�D��	�u�þ������9�ͺ�o���!�$QQ%�g�P����fm�9��]h���B�J6ېw�K�͖�����%�5&Z�$$���$�0<�q������Dk9���Il7PȠj��}��s}`s=���=�����~*L����s��X�}��76{wU��>����)��j �R�����2u۲V�T�!�S]�W,��I{n�ud.N0��I8;�z�̓�fm�����uh�VeD�!)�a��o���o��7�]sے���2����7��S������X~]װ�vVg�"&Z�"KNܱ�k3}��߶WL�ݱ�����T�]�P� |��~�������ɩH��2K�o� w���;�����ޜ��E�҈��a��aEV�v�݂v�`{j��U�4q�ۧnolW�_O��L��R�C7����r���\�l���m=)#-Em�-��������}u��(s���G��/� Je���',����G}�wvwٷ^�x?:�6 �H�fjfd����*�vU���o��u%��+D��Q4#;��A�f��i:=�9�l?��g���f� Ds��E������E�3z�7�M�(��*�dd*	�)�@(� ����B�P��@�KH"�@�J�%%�
P��bP�A(�P� �!��Q)��P(PhThD
E
TZQ�B� 
DT�ArA ZAJUR�")QBX i���_� ��iQ(PZAD�f��JE�D�`!iR�D��QE
)
 ��	 F�i(P���T)PJ"(!��B��H�0�C �L  ҊS�٠T�$H�T )E((� �� ��(R� ЌQ�@��!�@��҅!H�"P�@%�3+@�4ХJ��B%�-(Āj$V�$@��X� ��
Q�J �J$���X�X$)����P)�hXd��(R�P��ZZ@(ZZi & )i"JB$Q��bJQi� �i �EbEb(R�
 "
@bP�(@�iDh&Q�`@�T�%�D��R$
Qi�i!��! �R�
AB�b���dh
bQhT� 
�h)V�D)@�AD^J��
�R H!J��B��Ҫ(� ���H4��P�H�4
4�4�P�ЀP�P��� 4� t��p��� ��O�
Q�����?��]���P?��)�(������4 M���ꊒ ?�@��E?���(��������?������������*��������� ��?��o����S�������A_?��.}�O���� �*���C�E�UQG�����C�����⪩�����?�����?�O��BZfR��p�3"� ��Z����%� �� � ��˃��PAW�?��?n�������ލ���?�?�����'���o�b��������{���F�D�
U)D&@`�`@�JUR��E"TI�R"TH�R�R%D�TI�RBAHd�!D�TIHQ!$�TJAH��TI�!�X%�I�R%D�Q �eD�$�eD��I"I!D�Q"I�R�D�Q!�RTI%D���RE�RQV$Pe!T		PPRA	H$$!$ %d!a$	RBBQHI! B������������R ����$%���bBA��X	E��RBD��X ��$$��	d&D����I��RHH��$��BYBRP��YT! ` Ad E		$"P` Y	HHa$$!�&	H��	!$�&BH��@�	!!$	BT		Ee Ua	 �� a$Ua$A�$@��	�$B$%�BAI	 d!!$	IBUVDVRH e��"�	H�%	THH��e��
��HBBQ	Fe��d(BP���
AS��&@�@@�	�	B�@��(C(P�*��*4*P�(P�(�A@� H�+(�+!!	
�*2�����	�R�
��P��)@�#H�°��00$���(�B�H����2,, $*��� BȰ$,�	 �%@$����� �,0�(���@��!K"�
�(��"�%*%� ,*B0�H
$�**ʀ�P�2,*J�*� J�-� D���D�H�ĂC��� ��+
B���H��2
B���@�
�J��R�2�J�$#
�� J�J2�J��2"�"�0�"�+�ʄ!"��@� �$�J�(B��+"��$(P	������?���O�k�]�"(���_�����M~ן��lx�����AW����k��y�_��?��g�'_�M#� �����UU ��_���u��՘y�_����*�EPAW�G���v"
���3���a�AW��xh���9�Nރ_�QD�n �3��f���� [������@AW� 4�o�_�i���H?��n� D�����TUр ��/�|�������\����������)~�?�̞_Ӏ�����������CZ%US����w?�����[�_� �*��:?��J���:<��AW/��G�l���g� ������PVI��W}ߢ)�` �����`�}( hiT �� ( �   P �v:p ��@R@ (s`� ED�TT$R �  dP����B�T
 �IT�H�(�
E��((
 � �@p     �  
 P � s���5NY�a�`��=���ϪY����N��a�6�� 4�o��f��\ 5�}ީ�n�r�� {�x+;q�>G��W6��*���Kå���s���u/N��   o��� �� [���)JR�ܠ)K,���t�7]�JQ���9�)nܠ
\�Рn���s��R��LҖcB�1P  � 6 � W�� 8�)�M��B��`t���
��y������:)J]��QOM唥�( Ǖ@h� h �q�@+�=�}��WsC���m�� S��+�+ͫ�J&�:��� =/Q_u�=���  ,w��{o�n�^����u��ۼ�.��n�t<�ť;�@}/�K1�����|ǧ�9�p�=���   
 Ԏ�����Www�7�ν2��Ꞝ�X ����[��1�y���;O{ܥw�PV��Oo�C�μ 	������{��L��3��飭\��=g�5�u�-��_st�wr���7K�締x  ���   >��B��:�Cs>���z��w�}�|J� ��ڔ���W}�K��_<�7y2��;�� ��=��JX�l㡓�w,q�j�k�������Z��WA�ˡ���w��|     |D�&��R��  D��R���	�ɀD�*�*���� �5=��&�)P   �Х6ҥ* �"B���➂}�����������R}����k��TA_���QUt�*���QU��"��AX�*��~�?�/p���
��,	���a�M����/��g�.O=��HR���-ך�)�D'�s9��i`P!�8�5�xs���"M칅�К��`0QF�o?~_}��9��?�~�{$H@�#[e J˲7���}�D� B!$���"����j$xd@`�#8��o^���S�C^��a����HG \t� HB���*�$Ő��>܁���f<��dՓ!�6K�
���0cl��lB�|���Ŕ��q�S�cR_Ys[%��n�r�j�P�%�3r�8|Si����:�Bji��~�j��.�fh�aCg4z�6����5Y�q!�JR����0b���n�纞��B��	&#IZkÞs�����
M�6_#n>?��Q�_P�㮜��1*��İX�j�py���g7�.sd��E�2�0���d#�v���<�nA��ltBdB��_�^l硲1M��	.6��>W_oЅ�e��b�M�~z	�����}��4�ܾk�m>r�T�&z]q�<��;�����"���SÌ�֎37�cJs�B�/��\G9�Ͻ,W�^�!_`I���C���y��GL#�)����qw�������������2�`EK�(&�@��
)�AJ�H�
����"������F�s�� ��!\��� U����"B$`cčd\H��S0�́��/��'� �g=�GVp��3��}4�{�!&"G��B���$�C
A��ŗNo��s��T��iBV-�BX4�k�:��"�%�sG��xp�N��Q��M~�L�qN^�M
��o�%u�O��b�$%\a���4��6Cz�$k�+H�1k�����.�59��=���~G]�n'Ɖ"C�,&`�aB4��h����D�jb��D����/��HB�� bE��j@�T�"F25q�4� �aD�X�Qc�BW�J��q!�
~�ߎ��6��y���ю{�d���S�� Y����v�g���ӏ��K�B�B���I�j䎸oBk)�ѻ��ZE�XV6%D��v���� ���2s~��\5��rS�f�Uַ��.][Iu�<�o�LR��wd�[�4�$'<!#�)X��H@=).��8�����Ә��
1�c�BCy���SÙ��0��|�ٻ��z�]rni�X��9�(Jb��%"H�b��b�"E�Mt>�p�ʸ�TZ��ۊ܊��?�xvC�9�#�e?/Ԝ!5��<6=�8Iw�˭p�q�j�ɒ��!fͱ�$�H�+�r�����novB%� \6�����w{�ӵkBx�宮Oҵ�'f���o�x�o�sܾ���%!Y}0�~Ei#JU���+k���A� ��ׄ�ٞ{��	XH@$�@�E�dd`Fb@a	y��3�d��C���S��yG�5@�B��'������<�L���l�$�s�<5{�.��1aH�]A����L5��B���$�a(! �BE�GF8��`�H$�#>���o���a��$_yMm�R~�s-\��8�=!L�lЕ��&�З6q')��0�aL];���jEHHL�_tMj0�漾^��N�۾�g�>���H\[~>�$�ʯ����|��1�Ce�Z�)S�ٔԀH���!Pi��e�K��ōt��Jb�6�%CK�$ H�\5��o��]jB��4��
Ѝ,3	�^k�ky
Ǒ�	/Tˌ�-�y�ߏ�S������YvS�E�.!Mn5$tP�hf�L��e��ֳˮo|䑑$b� ��N�p�.:7Î�I���%3F�潚s\��ci�@�1�4İ�
HĐ�@Y�I�||l�Ƶ~�@i @��}���@8���m�>6I�2B��P��#\!$$\4�؍p�J&� P1\��3K�!��BH-�V@)! �q�4]���ٮ]�]�A�H�42�d��jA��}2"cE&��I#���e��$��> ���k B�Ia1`@!@��I��Lt&�5�q���|5����ݘh�x@�D#,�E I �DY��F��J��8bE@kme�I��Ѓ�x��\�`�& R*�S�Ȅ�~���W��98q^Ж��q�Itr�[�Z|>��诤i�Q�@>,!-r���4���$(�|��0�$4h�5�k7��f�n�	�=<�~�,=,t�K�JCn���i�D��缎�6}�޶B��l�f��B����k�B' �o4B�!�406@��<�^�8Ԇ��ύ��D�S1aK���=��4D=!}���I0�C�ɐ����h���k����˿&��O#p嗚7��x���
�Hh+���a����$.3���}R؋�d��0�_�˰���SO�ߞ����1 A�5��HV���r�0��f��(@�����@�{�l������%h��Ò�TD�`�1Y��4Ig�~�N��U*�CS�Ag��-�����F&�t8���p��@�Ʃ?�Ԉr��>B��D��\ ��͉�c4h M�S%Y�L�K�o6�n���@�� ��ɼ�d=�-��ڐ��.���XJ�0��d`JJ�L�C ��6Fz�zH�a>]�gWL����}�>̻)YE
�i�~_uW�s️���/����)�%�%A�;NN#��0/��5�A��.DOÂQ(�$�8�G��=�W�ټ��O'��<�o&#��ʿ~��~}M�%�b'qL�?��DT�3��`�?ݵm���`A�d+5��B��1 �����(�0 ���(K(S%hJm�P�i�{�X��$�H؄s,��d#����4��}����x0"B��.��aN{�*E#�)̓߾�xH�`��@�K��)�[ H@�`�(BH�"1(�"A���� `��
��F@!�3����	���l��C˚"�ȑ"A�aJ2)$�bV6�d�r�+HO�#ie,`A�c��qxu��L5��:������=�<7�y�9�x\2䐧%�$4�A�&��߆�筁$��d�1C���V � 4�5���2aN���1����g�K���_}6C�� �3�M�6\�<���$8�}C"�9���W�H��Q���!�7y��O}}!w��g���m D��Xѐ��x�jM�v�{H���@��<��8:!aA�$b����	sM�0��&�&�BM(a�w����~��%��LEƂ�Q]�w>��uzI]�s���$֙�cs�G~{��z��$o��^>�Յ�Ě� ��f�:39s��U|&�5w�q.33�߮����@��)	|3��K����#J�!
�|g��g����x��������5w�9���m	�a���߾owV{�ߊl D��)�/<��O}\�1q"h��f���9�6r��AB1!����q"MM<����}g�!4m�oՙ�h_�,���=J��{�iY�i�j��ysM�e�YYo�:�>H�j�d�`�И'մC���^pDu��#���5��'8��d���o>��t�[��=�ޚ�Lp�h��!���B,$9rѣ�q4�RkF�WZaM���b\���(Fh��ߟb�xr�bD
A�M���y�)�	X�CHi���\����l��������FJ�MU�3�# @�=aP���"�p�/a�
l�34�a�H1���
��h�@�ma-d�/�0��B������Mo�2�˂A�(V�	r{��=܉
F�
�o.�ʔ#Z'�#�P۷�eL�lܰ���k'��OP#��xB��$i,z@���r3<2�s3�
��#�{7��I&�)Ij��6���$#�U4�I�~��H1��Wt�_&Ӟ�Q��R12�#�xz!�T%P�c���������S�1v�%�C�&�fs������[���SY���߶_��Y�����<���K%O,�>��3�����a=���|?C���ݙ��"~}�}+6��\1�4��I]�:�4ԩJ���X��Ɛ[��Mn��L�D�k1�,�h}����X��,6_g3w^�	Hf��%�q#�dI�f�1����Þ�$!����	\����6��1 �n�edpM��zx@�
`jP�а�5���8F�$��� �I�.���^~��w򪪪���  m� H�   �h                  	�[_�> 1�                                      m�  $         ~��   �      6�`  �    �� p$ ����     s-�ÂE����Z��Y���xF���,g���:�Z;/*� ��c)s�u .���X��0	>_��D��JV�靍V�����y��7bݮ�Z���j]�Hʻ@x(�k�4m�P-��m���`^"7R�U�;[n����)-��V�V��v�fF@��m��@m�  [�}�~��7e�U�V{"ڶ�$i�����<۝�k����S��=�q<����=r�ƞZ�$Nݫ�� Kj���6^�*|��(sѩ�*��hㄓ�E��X�� ���p�q��� I�̪�79�5l�UT��uY�M����T�6�ZLu���`�`m�k�k�M� h�v!��   �
��[��u����m��	 $h�  [\WS�A�X
����
����m�%�2�5�g�MuUT��p&۱�*� *kח/�`M� m��H �;m�Kn�H���Um @! �� kY�dm�ͤ ��
����e���5��o�o�[wÉ$��m�n
Z���O���Ly�$����m�˭���V�tPY-I�++RtijCm��  ��H>��]���H6�Ni�� �  m[H�m��rL����.��uH V��jXWM`���ɰB09���� m�D޹���� ��
S��Y��ح�U�O,�ѡ��8�6 d��m��m�l]�4�v�I�o�ed�:��U�`To;PQ1���[|���Kt̢3ˆ��-��y[��#�z8��w��3�N��Ғ��Ʈ��B�ig7)���Jw���C�H]c�Gf]ؠ�T@�2�!��Wm݂qe��!@y��a��S��4J5P&��HH��v�m�"&�\1.�4-- ��i���.V�T����M�z���r��c�V�y��:��3���]J]GG
�mJ�瞞*�v�l������5UH'�}��|E�Uk����8FK���ҳ̍v���)�t�]Px�0CU�;Î1�gB�Un�J�Үյq)�ګ��n�Ն;�'����v��u�e�o+@T��9��gszw�vy��M�pm���7b��>g�6T�B���/<�,C�b���AC�-���-���@�`8l��wJ�uY�µk����;����!�ds�B�\�*�G-�����R�6��
�6�]��,1�V��tM�1�y�M��2!i�kc�Ø���Jlm F�*q=U���@���'�6�!@�֗�zH�M�O-��1�.�W��(Sӱ�e('�I����N�l]�3ܯrmm�j�	��uN�k������pj��ݔ���M���a6��X�!&��ㆫ������U��V'GR5PP��V8n��[�H���M� tjis[ ��R�D�UJ��Dh膺Z�.���cJL�W!*�Л@@��l��6xSj��@b�����+�
�I�glkp
J���猁+ ۶��ꩳ�e�0 �v�Ӳ��P@k8�8�1�V6n��/m��(��:�Sl�i:���r�ܖUvPxyẜ�=���,�̝y{PM�K�\�\��uk�$Ŵ,�]G�W-�&�
��][*�k��Ҭ�/[��!]�m�8-�$� ��m���`q��k0 Wd4��vj���ۆW[�[@Ht� �[T�����M�	 �I�� �JM� ��/n˰�[�
�
p8ګ#��m�`n�[�E� �i	�
��UKqd���VR@V .�*�r.ҵTtdeeZ
%�B
�@R�]�\Q*�GK�I�'` i����`H�a�Q����3`���Uj����iZ�%W�$Ұ$�c[qm/�s�c'�j�������?@��M�I	 -��t���^YT
�Z���P],�� �K�E��oZ�0+�=�M+ܵv�Y�g�j��L�PF�7UH֐r+U��nvr�UV^4���4��g��R��e�G=���Ywg5k���P*��붍Jm���\۳�:svz��^Y-��2�[xkWOמ��r�z�v)���[�7!Ƿ5�zrt�����B,�y�!��ā[��i�������U��m[N�$;"A�  郎6�d�� ��/�$�m�mu�r�H�z���.H�Ӣ�U�U�&�fYd�۶��ֱ��k7�>H�[B@m�O7[�8
�"ڐm� �`m�0��h��0�h ��I.��Ͷ����[Kk��Ce����m��j��j\v6���Ҧzi	���R��R����w��"�  m��&�6�h��[��%AV��` ��V�`[��6��M� I%[YGh�#�Sy%oV�PJ�#����)M�$���n� �;l�lCԤ��;ck���!���%/Pu������V�![�[l9~������]��`[F�Xm]�bͰn�-�D��[Cma�U��	R�'I<�l���4���m��VQ�,� mns���8:ImM����I���:�JI���A�� F	hr�J��S��n�b�m�jA���]@��K�0B�l �d�Z��� �vʻ��͹*�]�n�p5J����y�-U�N7Ұ\�L��Ӭ��hʸ� �XI�������̔2�US��Q�4��WT�r R�W)W�kh
�4�5��i�ntW�n�v���m�dF�^V����ٜ	�:�e����6j���t�	���1���iscK���g����]9]��F���5�i+�GT��Ȫm�D�f�{<�A��muV��m�te��
��[[�����饵i�3��VYXjn(=.,3w�'u��vշ�L�n�$2c=��-��THD7<r�MU�*��i"i]��Wv4�z�OT�Ʃ�]`��luˀ�IꝐ:ꪔ͔�a 
��]�ճUl��6r*��� -Md��v{vH�i�BF�-M�h��F�&���h�U\�ehA��]�u/e������9�zc����Z�%��W��W��H��-�����'l8[@�l��PUm��q�����c�iY]�*���wg�J��R�+�� k�ùZ�e�.����6�iKg4�U�R���[];oB�ඃ�R���Nu��n�Hc�-��oIh3��UU�T�r�<�i[-�ж�H ڷﯢ{�2daiG�Wv�yX,�h,��pe�%50����[u[U�uWB̸l� �m�I5�ݷI�_I��  Ƶ�m��nm�� ���Ͷ$��D�m��  �h��b�S0 �( p$ koŧ��  2��l �-t� m��.`�I�� �kY�Ƶ�	Z�jU��vm�4�Y+*p�U�8Ӎ\�Y��66�b�Y�M��	�@6�g  -r��{�8����e���V�ej�U��p;P�+Ppp�� rޣm���&YC�H$p�c�   ��s�kX6�mMk䭩K,��F�*��V����SMn���T�[d�j�p��}�#m��/Mnq�R�A�kn[M� $�p	k�Ë%��ܳn8�zʱ(�/i j�m��m��I�   .�qmm��5�i:� H���-���� $�n���  �� �A�m�ƶ�h�m�` M��ͳYg� �[f��S�]���m����8
�  �����p�kh   (l�v�HHu�J   �L��$6ض�M���5��ũ�$�b@m͖����[dӝd6q�J�v� �i��3L�^sm�5Mq8ڻ` H�A 6�[R,3�h � ��3`Reh *�����@���@"LuB�U[A�R��5����8�������kg���v�������Z��sK����0�qm�U�%�Rմ F�L�L�	m:�	�l�8��4�r^�#Z�)�F���h6��	��ۀ � H8 �� �`!�km��l� ��6�sE�WgRJ�l��Z��C��\�5T�[ � ��iX-�m#A���6�I�m��   �oP�`KI6  �!V�M�[6�	���@�`H �Ŵm���}�m��m�t��M�H�I�l�`;m��
.��
RU32��4�����`�v6ٴ�
��u���� �.��jk)��·���;-K�K���]AԺ;!;���T4�tͶI�6ͷ��$�[��K$��Ll 2j��6�H���  $� 6�6� ;k� �-�kGH ����knݖ��Vs����n�d[�����k��� ��g��@?�Ҿ �� 0�Q�uX���g��E�|�S`� AM��P�GP��")�� H$.z�p�6�1C�h]&�7SN	�� >�PЮ�Ri4:�@�iE�!�C�
H(�`b�1@ *����E<D���z>���S@� C�!�Sb��=Qv'���Xp^ ���/�?UA�|�x��A��~]�lU� z����� � >!� ;`!�D�i�E*'�����]
��O�T�X0؃�"� b|�O�X�X�Eb! �����^ &�>@��`�� �����_�^*��6�GXA4�#�*p���^Qvx���	���� ����>4��� DT�Q�>�S����~���c`��@h<�M!��@bc������>(>���PJ�a)�@ ��S���_Au#� D=_���hM �"F0�a"��Mh�$!E�FdHFH�dXBA$$	! � 4� �
�}TI��$��C�| }�4
̈́X`B!A!"H�B HD"�H1�H����B0��U�Cc������v)���"�ȧ�$i
F�RńB� D�Y*�"��_�}�� ��@�IO�T�v!�&� �����	�~_��@Tt ]�H�q8���1D'�G��T!H�O�QUx����(�% Pb� �6� [U;��u�kZֵ�J�   m��      $� �	 :[Gm�-� Y��'h�:_��y�r��\�f�:M�<���b�����g6u\�WF�:��{m�N���۶V��T�Ĝ&���R�y�v��X7;���]�M�z����J�(��:�sqU,!�uӼ�83a��J�Ѣ孺U�OD�bN���g3p���y0����ݲ��H8(��mX��XM]\�8��'��l�MO�nqbx6��n^U�5�.`�Q�H��K��[{^��3��� �⌴�:f�l����಼�Z�#Nӷ��8.��������:������I��6�K��[p�4�yݳѳ���ڻy���nv6�6�ml��v���F"�ck��X�L�u�t�m�!��/�FqGpq����mf��u@�WkE��j�ِx\N��䢸�jg� Q��x�����"�Ge�`r�a*��Sqmj��x�n�Ӱ���t�)9൹���&�#�C�N�*,�H�J�����`�&�c���]e�8�l� �ݪ(�˝��z�Y]1@��S�Sg��
�x�Sݭc�{<9Y-N+��uZ�gz(�.�D��t�:�5eɰfܹ�j�C@@KͶ��ݞ +.+b��cY��1ԙ��i�\8͓���n���O00k���9��c6vG����Nv	��؋v�g���ĥxL�zU�eg��X.�d�vum�i���8�%ӫ��9��]r�á��<p/]��*tJK�UK��uU��5`��tT��f��k294m��T�&��!!l��kuH��:S�-�=bѕ�e���%F� �մ�*�۶n9.-d�a`��pN���[ �/nl1�$l5+!��Rv�l�� �f�[Fx 4]K�j̄��Û����,�� [���	��6W�,܌�-��B��x6�y#���:ι�P��f�&�t��ꗁw ��NyB�lh:M��X"�.vW�Co���B��e@u"� �8~N!�P}���>LQ|D��{ ߇�0ְl�uݢU����5�J���s��M��\�W��㶨^^�v
��c�3��y��<�9Tu`N#�-͜uۏ������;���K!q�w��z�Jv:W#k��<9�u۞���.�=��	[�A:��{-��Z���m;v8��Z��Wixk�A=�ƺ�k@J�[�ڵr�`Z&[kn�l�m]>��e�n���&�ṵ��3,̹�m���0!��Pɸ�q�]��g��g.q��ls���j�����~��@���o�����u��� �ӽп��
� ���D�u��z�˻J_���H��CĒ[����//fB�-�+� n�/�H�CĒ[}���$��ı$����]�Ⴖaw��_�=��
}�v_�$�v�$��͗��Js[S��`4�+� }��}����� ���w��_�=�� ��ݘ�n��vhp.#�	J�2��v+A���-v�s�z���.�i6+H�v�_} ���< ?\�|�BݕoI-��J@�I\(&Y)%����{����B�x�3�y'9쓒!N��π�����^�����ي��.]U}�����I-�Ww��bI%��|�D�����[Yvg� ��z����-��,I$����H]�V�$��ݺD�aX�_} ���< �����_���� >�޾� }����\��iۮ:�;V�痪pȸ�����v77ny�۵
�u
4�w+3J[�����x ��_�I#���ĒK{#���Đ��.$_��2�����O 7�<�t��ݼ�f$��鴍{ƛ�����x�t����ԑ��Fb�#�"!#Q ��&�w"s��)�v!��t�һE$�M��� vlx�지E6^���%l)v5vـlx�지E6^�c�݀��Z,�i����n6��s��v� �vx���w-�
��CKY%x";Qm��wU�����0M� 'kaC�	�:.�M7O �l��Ur��;�~0ޞx�지E[�H��J���N�n��0M�U$l���yzz��>��H�'C�f I��we<)�ٹ>'�8� pA�"���p����Z&�����we<)���8`� ovYbHI��`K�2��f�:��/Z����}��������;�<���S��]}��l��0M���$�<��1W���wh����x�8`� n지E6^45�ؕ��]���f�x��O%����;<�`*��rW�#�
[g�,o��W�y�z��p�"�/ 'jB�]	�:.�Mۧ�E6^��}���^�� �}���X�F @F����>����$0�l�/BY�sn�'%Ļr�ݞq�湵μl��.�n�JW�6�n�6��W<��sl�0m�Z�]{b������s�͠��8�E���`��.�q�m��Ң�n������:7Aɖ�m�v�C�N�?�xq��њb ,�E$=��GQ�M.f[���q'vv�c� ��p>1Ŵݱ�7��,:6��k���fU~��������牝��Ӯ�^�ьݶ����۝rȋG�k#�<����(�O�pk��t�����M��ݔ����$֊��@��w�E6^~��d�>�����7_ ��כ!q��tQ7x��O �l��Se�|)�6ǩ9"n�گ٘�=����� �l� �지}؆*�un��E$�ݻ�>��E6^ wvS�"���=����l�NxUEk��A�뱣x+��0��t�g���ܻsrl��:h�`gm$���i[g�yzz�we<-��,K��=��>k��+�څ-���u^{7 @��X#c ��$"���, �B)D'�]�� �M�LX���(�ds������5�vs��{��H�PTH�Ux��Ӏ~ٺ����ݔ��V���I�4����{�U�.��� �����[�"�/ �5"�:'i	w�E6^ I%�)%�)%�wnU�+&	Ң�L�9�e��e���.��3v�g�+vƗ�"�N��ǖ)r9"�tQ�8�%�-������K�%t��i!�RH��m��of��>~�� ��zpwv^��e���17m���9~��ܓ���f��B����<"b�s*�\*���ğe��{�Ԧ+i;h�;��m��x$��	�"�>�"�5T�U��\(��m��ݔ�	�"�>�"�"�/ >ݻ��a̹��R]�Z��q�D��9���7`]]�=DW2{p��KW7���M�6�X��X[%���xU��)�t��SI�ۼ�r,)%���xSe縑��U�x4$�$��<�=x��O �l�����6+H8�tQ�8I&���x���7$���rz���*�Sb�}a��}�י�'ǰό���h�-�O ��� �Uv��׀�u^���sJ���&�2�$F;ݸ@�n�F�y^��v�Č�.�.z��n��
n���춊I��X�Ix]�x���;{٢�v�v>!ݍ6��we窩 �z����^�Sc.�k�i���x���;���X�����M�u9rʯ ���^v^ wvS�"�U�L�6T�n�%8����<�;�O���x�p�6��;����m�aw}��+��݇\CgF�0o��v��
�v�P����Ƌp�t�랐�b:KJ۝ãp:5��g����iv�����Knz�c�!�u�;�Sm�Y뗅^��ծ#c+r7OK�a;B���<��Ҷ˵�,s���s[=�u�"$ݶԄ���X0�qvs���J�0��hȶ�C����ٸ4�t6G����?��Y��38�~���[Nc3�����m�뉝v��mE�����uc���0��k�)m���(���o��߯ ;�)�u� �c���\�����BeZn����7\0��X]��	ӗ�i"����&6�<v�,�ܤ��z�d�<��SU)U�.��e����x]�x��O ��� ��/-4���Ć��x]�x��['������^ ~������3X�%�ܗ[m�Y�mId쑳3�l<\�{u��l���*�MIVۼ �지M�� �l��W9\��}��:��y���#��U��߳{O���"XB�p�v�آWx#Vv^ wv< �지j�U�N6$:T�wj��>[%��G�ݔ���g �za�����r� ~� w�)��K�>�Ȱ���WB�uv&ZM� �vS�5I/ ��"�wv�bğ|�"���Z)%�����Y�g��OFCH0���ӺvɆ�;j֩6�%�:�m7K-W���N����G���x��SU*�+�E$��w�}ۑ`� w�)�����I�{�ӑ��-hu�k��޼y�������&�+�<�m~
�֗K��5�p5��37��Vh�͠TЅ���)! �vi_� �{���>2�f���cWA�9����۔*��wVQ��no��DJ� @�H�!�@�/�=�{}D��6>/���� }��&�:h�p׸��0�@9�8t�����zxk�s���x����|�:�g��`�<�[��G�3b��&	���P6���E���:��HO��c�:���8���I�	@<��|p4+���+�H" J"�M� �P>��4C���0W��9��s� ���ulQ�V���Zl�v� w�)��ذ�r,�UIv{׀u�T�+��E��]���;� �U]�����y�we<�s�����4n���ӧI|�Ru�l6x�x��Ct76pݬ��ifZ�䜤��<�@�"�mt^�����we?ܪ�?s���������5X䃬r� ~�?UW�]���O ��ߖ�엟�ʯܻ7������c��[��+�>�a�K�}�����'Nk��*�*I�ۧ��-��XV�׀�����)���5@(@8ia���Kڠ�l�z��>�������v�k��۳�u{1d�z~ ݞ��un�}}���V��M]eKG��	�����&�ƤF4Ϟ�y�{fw��뜽��n�P�,hu�l��ݼ ���v�,��/ �lW*��ݮ"�e۶�����{��/ >�<�SQdh���*��v��>S޼ �H�����QV�Ҥ覓m[X�d� �H�����{��%*hWv&�n��#�=\��=O�$��|�K�>�Wj���^����u�~x� V��K$mk6�F�����2���|��I�EϮbu�8zz�;b�s{f�Fu��|])���m�`u�G����Y6�S6.��a۶���Q�8�#p
�55���/d�B^�vy�6�63.�M��@w��s��u����n��Onv^�z:v�N��/gWg-���ͺk�Z��{l[�v;����r<�S����Gbm��X��+L�k����R�K;���C�ܢ��$\Dj@<�X�؜d��k����t�[����=:���.�i<q(�qB�d����������K��� �+F�@�Uv�&6�<�{�^ }�< ��O �j)��7E��)&��X��X���we<�{ݨ��Bm��j�Ҷ� }�< ��O ��ŀ}.E�}�́)j����-�{�W�fbY[����y`vG�}��TZ-K�T�t���ly�ۓ�f�9�
4��$ƍ�l��e�Qnt̮֙�1�.c��b�>�"���\���OS�5W��B�T*ݵ��훯����%�X"Id�Y��>�����U���|�,X�5�A�ɪ�$������� n짇���y`z��v^�*W
V���5n� ��O ݹ�� vH�	Ҡ�h*��$�ۧ�n܋ �\� ;$x����rN����;+fg$ZZ��ж���te�3�(��ٚ�i�%��n9s�ɻZuv줘����� ;$x����6^�凘�����M+m|7�x����6^����其�_,��Jݷ��)�Se��p�p�X�����P�@%.&|������?����{w$����rOoޑ��n��X�v����`K�`�G�䤞��j�K��MP覓�V�����������{ߩ�v=8�X�޾��T�%����z@��И.2<CZj��I��+m*�PŇ����n��2�4+�I����I�� 7vS�>�n�I~a����{<���ӎ)u�v� n짟�_�U˳g���7�������{1cg�g�F�y1A7KmW�}�?��Xz��Hݞx6z���{+�r8&�Ӂ���|�����=������TaF`{TP�"�OD:������;�>�sU&�*J�X��x�M�����>��vp�B���YcNT;�)e��y��s6c�m���`��3�m�Pp�ì�ߝ�O����T�G]nYo���^��p�>��{�����E�^t;@��)Z��n��c�~�~�9˳W�~� ��׀�u^u{Hk^�O�u�����ݳ ���x��xz��$���w|�p�j��
������=�����	��<���\�~�.��~x�k�Nʚq�"n�� �۪��ľ���5zz��v^)���wq�m��2���K$����T�c(	�7!D�*�U�.ƹ�i�^؋=:'a�C�m�mEAˈQH��`��Krt���w��v]qӛIzí�E�y�[�u���`n�Øt�&��k�����:���#<Om!��m>c���.����+۳y{4��@Ir�Upͮ1�t݁��3��k`9ؤ��҈�@�%�<6ƌQ���g'd���I&�����m�cvJ�8�w��>Q�<�D�q����V�F�p2�B�k��d1�X�m�~~0�%�.��{��Ȁk�݂�VRN�l�:���ԑճ׀{���{�V�M%|i�J��ۼ�ݗ��S�>��XT����ȉk�d#��,����X�������~���%�.�Wv���M�J�6�t��{�$��ݗ��+�;�k�6�%,�#� �
�e�X�[\��1u�F�i���5��r�J�s�}���m��i2յ���x˻/ 7d��|�����~0��NH�N[x��f�����A��,]Q���K*Ʋ�Y��aB^y^����ۻy��I����+%Q8�7T�� n����{�r�˳��~x��׀}ӗlmjN4�,���,v� =�z�����{3o۫׀}��},�$����k 'dx��?W+\����{�x�u�ϡ�19��+S$Q�G=v6��Ы�XG�����grl�F�ۛ�#v4W�{�{�14���@ջo�?r��_��� ���~���o��Z��m�W�-4ӷn�nǟ���s�9vl�~X�~������<���0j�Ӎ[\��y�}۹$�Ͼ�� PX $*�Q�� "�T�\ �Ē�ru���{����{�B���I���s�{}�ul��ݏԾ��>�^<�y�S�7T	m��ݗ�{��/I��۞X;#�5Ir� B9u���m���u��BE�])�l�c6�h-���J�l��e�9����fhcM��[n� ��xݽ� 'd~�s���� ����"my'n�Kx�u���o����� ���UI��-�$j:����=��??����b��������;��πw�M�[s+,l�n�=\������� ���`v��7�(b��6���u���`y��_,��Nݻ�ݏ �\���l�~]_�� �we�wcm4�.`a4a2��]�b����W����;t���X]L?�Nm�yk�H���m�v��^ w��W�r�]�=�~x�_�t�S��1�m`)%�m��~��ı/�}�m9ı,O}�{v�� 6%�by�3�I�$��e�,�k6��bX�%���[ND�,K����ӑ,U�,O}�{v��bX�'���6��bX�'��t���f\3u��ֶ��bY�(��3���m9ı,O����iȖ%�by��siȖ%��D���L��ߵ��Kı=��3,��)n��5��"X�%���nӑ,K��C�~��6�D�,K�����r%�bX���bX�$C���ĬBx�j_�1~���.��#y�5|B>e���!�H�@_H�zJ��b�l	��6�<�{��C���J���G%�2 B:
r�1`@"A!�m�6.��cf�>�< �5�;5Ğ��8.ͼ!T�xr0 �i�IA1 Z@���B���<����a	#�d�HHH&��aF#�����`x@�(V�զ��4h�1�K+a<6��: ���zlyI ����&�b'��F�O��M�	���0\CPB٣+*l��L6�����/�C���������Ӟ�����ʮ��UT  l�h      ,��   mI7`�q�ӛ�tݺ�禓���VSw�����Fu���]X�
�9.�t�!J��ف����7��K^�9Nj�j��Gޭ����AM�ذƳ�2m�Ŝ�w4�讫������J�ѥȷ6��($*�5��2�$ՙ(z�T�6F��2�OSY���^x���&�Gf���N�8�tIƘ�n�w	��[X2��\�p+ϳn���\��qΌ<�;l�Жx���.k�ЇNΐv��nwh�F7gm�2�sـ�`������ʣ��v����3��M�� 絶k�����XP����6�F`uĦ�v��p���ț؞[m�Y�r����F��.�ú8�b�xpq�LɅs�����������
��h�)���A˰������f
q��*Mˁ�襭���g$�董��ͭ%��v��'}ų�[�ʽ�<�#V�<�P�)z�Q6q��u�M8*�U�!�m���Wi^6e� �8��ݠ}in:�bծ�I�v�%y��"Р��©��%ۆ��,�̏h�T=�"Y��s��{s���;b�__.{c}s�:F��mr/g|q-��d�cu;��枌c�I���m�n9���� <�gn���+v�Y�=En�m�/�'O:Y�f�vw 5(�;�p��vb��O=�$�����땣t�w�j���Ms۪Нi-�;-ۢ���s�q���
�nì�&2�\d�u�+��T�YX�<[AW2+v���
!Bv�me�#ՉTf�T�6i:���8s�mű��'s,\��Bl�R��oQmr�d$d�^�[$�t��6�m���=���N�՛�iS���Y��9�J[nM[@�uT�u��޴v���,]��ӎ�м$�\�λ6���p��8�Ie�CI��+�5�K:݁���Is��vq�$�,m����m�6܋��������V)�u����s�I<��	9��I�P"�*��/���AL�Tz
!�� ���.�n��-��Uu�d�-[5��y����.7m���v��m5m�q�'pE���ny ���/�����&������oXj�4����S����8vS�7y{2��l%)R�	mYF���=FΕ�hƶ�zۡ�Yϓ���:��J�7R��rR����C]ud��M��c��ʗF�p<pn�-���',:�SJM�J�u�Xؒs�s��P�*s[5�Ys�Y�Y�p���ۢ�e���yM���F�4 �>]�/6ۇt����r����$�v���_�L��Lž��|�Ȗ%�b_}�u��Kı/�}�m �Kı=����r%�bX�zMwҶ�*�l-�W�_�L��L���z�9�� 2&D�/{���r%�bX�}��ӑ,K���nӑĳ1v�0��Ldu����11,K��w[ND�,K�{�ͧ"X�bX�g{��r%�bX��{�m9�f&b��SŐ����m�/�&a`b{�wٴ�Kı>�]��r%�bX��{�m9ı�/����p��L��]Qy���[dMV�rS��ı,O��{v��bX�*�}���ӑ,Kľ���iȖ%�b{�w㘿�����}�OВ��*���YH[`�V+i̍e�h7�؈�p�iUa�ش��,̲#�WT�7lv�b�bf&ab_}�u��Kı/����r%�bX����l?P_"dK��߷�m8bf&bf-��<���R8�M�]���D�,K�߻��!�4D�
�x\L(b+ < �Z!��9���wٴ�Kı=���m9ı,K��� ��2%���jt�-��Ku5��m9ı,O����iȖ%�b}�wٴ�KKľ���iȖ%�b_{�u��Kĳ��������������LŃb}�wٴ�Kı/����r%�bX����m9İ?)r'�~��ቘ�������ֱ�UV�Um�1~�bX�%���[ND�,Ko����r%�bX���xm9ı,O���6��&bf&b{��Э�*�Ryo5��1��㠛�EH�v�a��˹������p����K�Yo1~1313��bX�'���ND�,K�{�͇䀞DȖ%�}���m9ıLų�_�0j��4[]������b{����D�,K��{�ND�,K��{��"X�%�~���iȟ�,J����E�ן�m�5[��W0�Kı=�߿fӑ,Kľ{��iȖ5���ș��涜�bX�'���ND�,K��N�Ք�]�3W5�m9ĳ�2&{����r%�bX����m9ı,O}��6��bX��{�&�)���R�(H�M�]��,A����\H����iؖ%�by���ND�,K��{��"X�%�~��a;sZ՘�cU�i��WK\İ`M��=;��e�b��;d�v�Z�%�@��ɈB�!�v_9=��%�b{����Kı<�{ͧ"X�%�|�����Kı/�}�m9�����?����Gj�/�%�by���NDKı/����r%�bX���bX�'���NE�313��"p�[amr��,Kľ{��iȖ%�b_����r%��b{����Kı<�{ͧ�131}5��,%&2X�r�y��,K? �������r%�bX�}��6��bX�'��y��K����H��T��##D:E(�*�ŀ��=H��P�.w���r%�bX�g|����TQ���y�񉘙���߻�iȖ%�a�"}�߿f�Ȗ%�b_~��[ND�,K��{��"X�������۶\(*3E�����ץ���ͻ��-H��+v�̭�#��Z��9�Ny	�)�m8�[��Nb�bf&bf.�{Ә�ı,K�{�m9ı,K���
<�bX�'�}�ND�,K��N��iL�3Vf�]j�9ı,K�{�m9Rı,K���bX�'�}�ND�,K��{�N@D�,Jb����R�c�7ev�b�bf&bb_~�u��Kı>����r%���b{�w���Kı/��u��K�3�2�6x1ƛ���b�bf&,���ٴ�Kı=ϻ��r%�bX�����r%�b-�~���ӑ,S13������+��/�&%�b{��siȖ%�a�H�g��~��Ȗ%�b^���m9ı,O��}�ND�,K!�t|�{��ֵ	�ha�t��Z:�sj�Ů�M�N{rPc�j�|��C���-�X^u�A�����y�=s�M�A6�v(�]z�/��L�sr&,�k�{l����������KUt�;�8Ze��m�c�I=a8�:]}D��E��B��!
�a�3���FF�).�NB�#�	� 1�n�x�1�^t�v��7X�q[5�X���O�'#'��9�.g�,������v[��۝�(n��\K�Jyϟ\�&�w
�<�K0�{��k�'�ywk�6�g��Kı/߾���"X�%�~���ӑ,K���ٰ�DȖ%��=�Nb�bf&bf/�^�5a,bqٚ˚�kiȖ%�b_~�u��?���,N���6��bX�'��߳iȖ%�b_;��i��%�b}��a�e��
��ie�����L��[�����bX�'��{�ND�U�,K�{�m9ı,K���bX�'��ת�c�U�l��/�&bbY����}��r%�bX�����r%�bX�߻�m9İT,O��}�ND�,Kݡ�<�M�Yk%����������{��"X�%�� ���w��m<�bX�'���M�"X�%��}��ӑ������Hy���(��9`Ȅ�Ձ�3��6[�սn��a[l�%e�n]���s���9KI�D4ݖ�y��131=����r%�bX����6��bX�'�k��T9ı,K���bX�'���6y!ț���b�bf&bf.����=��p��K����ݧ"X�%�|���ӑ,Kľ���iȟ��"X������&��p��u5u�iȖ%�b}�~�v��bX�%���[ND�Fı/�w��r%�bX���xm9ı,N�j����&�e�kZ�j�9ĳ�ș�~�ӑ,KĿw��m9ı,O}��6��bX��������Kı=��H���'��[Nb�bf&bf'߻�m9ı,O}��6��bX�'�k��ND�,K�{�ͧ"X�%��w�h���UdnR�Ҋ��gm�kn�X�ɞ0k�4n+0�8Rì��{��>N����n����k5��"X�%��w�ӑ,K���w�iȖ%�b_=�u��,Kľ���iȖ%�b|a���55p���]kFӑ,K���w�i�~E �dL�b_~��[ND�,K��ߵ��Kı=����r"	bX��ݡ�<6��:�\v�b�bf&bq/����r%�bX�߻�m9�@��S�V@
� @#��"�0#��(dL��w�ӑ,K���w�i�131}���J��CM�l���	bX"�b_~�u��Kı=����r%�bX�����9İ?"D��������bX�'�G]2���.an�ֵ��"X�%��w�ӑ,K�=ϻ��r%�bX��{�m9ı,K���bX�'�����
T锺��q�:ݞ؎]�L��f����0�t�1��x�vk�qv�7�h�yı,O���fӑ,Kľw��iȖ%�b_~�u�A�Kı7��˘������ګ~��X�]f�Y��Kı/����r(�%�b_~�u��Kı>����r%�bX����m9�r&D�=�o뜳#�	�d��-�/�&bf&b{����_�X�%���w�ӑ,�,Os��6��bX�'s߻�ND�,K�~�xb�6�a��r{y�_�K$���w��ӑ,K��;��m9ı,N�w6��bX��(�
�@8��C��L���bX�'��OʔC��ܮڹ�񉘙���o{�ND�,K��{�ND�,K���[ND�,K�}�ND�,K���ߵ�߻S�����w��v��p����G7a�\dݞb�2�0�dC{%�ɧ����.�fkY��%�bX���fӑ,Kľ���ӑ,K��߷ٴ9ı)�f�Ә��������<��I�D4�m9ı,K�{�m9�,K�~�fӑ,K��>�siȖ%�by�����O �ș����[-�X\�]K�ֶ��bX�'~��M�"X�%��}��ӑ,
�2&D�?w�m9ı,K��ߵ��Kı>϶(?�8�j:���/�&bb��[�w���Kı<����r%�bX�����r%�bX�{��6��bX�'|�~�
7cal��b�bf&bf/��w6��bX�+}�{��"X�%���o�iȖ%�b}�w���Kı7<����y���eM��UGeق֕��6[�͚יА�+{(x$89�>��K�%ps��1]\�2�hS�m]�^*T؁�-
��T�8��ywI���=B��g���M�)vÖ�u�Λ�����K�66�裮i\onn���A��@��'�\�.�Wk����iεUi#Q�\�x �O<����J���}��=t�]3Ȅ�F9c�Xٸ��m8O�{�}9�m�b�]}r�1�̬B2�y��2�N�&��m�:��3�ۇY��~�'��.�5��ֳiȖ%�b_>��[ND�,K�~�fӑ,K��>�sjr%�bX�g~�m9ı,O���p̒��їV�Lֵ��Kı>���m9�,K���ͧ�|��,K���ٴ�Kı/߿~�ӑ?TȖ'�w���%�&fjm9ı,N�~ͧ"X�%��w��ӑ,Fı/��u��Kı>���m9ı,O�ԞSʹ�T�-d�s�11f3����r%�bX��w��r%�bX�{��6��bX� D�����ND�,��[��_ĲɎ@hv;m�/�&bbX��w��r%�bX�߻�ͧ"X�%����ͧ"X�%�{�{��"X���_ؒ��m��I.T6��ܮ�+ˣ'�SW)�'<i��cn+k#Z��o
lv���e֮k5�'�,K�����6��bX�'��{�ND�,K���[E�Kı/��u��Kı;��9�$rQ�m�1~1313���1~���%I�HSԍ��\��h5�p,B�@L��!` �BD�K���kiȖ%�b^������bX�'~��6����13��~�AVڶYg1~18�%�{�{��"X�%�}�{��"X�Q�)�2'�����Kı;���6��bX�'��v�ۙuq�u���3Z�r%�bX��w��r%�bX�����r%�bX�ϻ��r%�b
��}�{��"X�%���wa]:2�۬�ֶ��bX�'�w}�ND�,K{�w���Kı/��u��Kı/~�u��Kı;���wV�0=�[&�Փ�۱�A�<�]sg%Wv0gy�BE/nQ�_���wy�����kv:+���Kı;��siȖ%�b_{��iȖ%�b^������&D�,N���M�"X�%�����~i%R��[g1~1313���_�L�ı/{��iȖ%�b}�wٴ�Kı;��siȟ� .DȖ'�{��9��e�������������r%�bX�}��m9�T�"Bh2�Rߩ�8t�M�~���I�{�d��U(�	=��x���=���&D�
���a�&�`��O-(eO�5P�e�Ǎ���&�R,��1��H@�XBh�$##8^F��=�V�$$���L��ja���e�"�r�j�'�A��1��� j�k`M�1 ����xM��p��i$4{�$҄.ª���ФD��|N�4�D �J��x����> �>�>A=L�Ҡ�}QS��D��0U�A�(t$O�k9ﹴ�Kı/����r%�bX�}}�Jt�\�]j�Z�r%�`(X�}��m9ı,O���m9ı,K�{�m9ı,K�{�m9ı,O���;��f\3)�F��M�"X�%��w�ͧ"X�%�-���bX�%���bX�'�w}�ND�,K����w0���m����3Fd(kh� @C��V�nvvܶ�>nL��t�_��{����p������Y��%�bX��߿kiȖ%�b^���ӑ,K����a�
DȖ%��;��m9ı,O���ɖ��cr�3Ys3Z�r%�bX��w��r%�bX�}��m9ı,N���m9ı,K߻�m9Rı,O���p�
�їV�eֵ��Kı;�wٴ�Kı;�w���K�EL��/߿~�ӑ,KĿ������bX�'�vw驨K�5nL���r%�b�'s��6��bX�%���bX�%���bX �	`�x�'�w�&ӑ,K��tό;a	��5�3Zͧ"X�%�}�{��"X�%��^���iȖ%�b}�wٴ�Kı;�w���Kı?�����@�\lфy�ݏ[\Q�wg����ٛہ��ݵ�,\CE���s�q<���p��Q�kZ�yı,K���kiȖ%�b{�}۴�Kı;�w�� yı,K���bX�'��_e%:KL���ֳZ�r%�bX��_v�9ı,N���m9ı,K�{�m9ı,K߻�m9A�,K��q�ˆe2�Zֵv��bX�'s��6��bX�%���b�%�{�{��"X�%��u�ݧ"X�%��I���d�&�Զ�k5�ͧ"X�~*�;���m9ı,K���kiȖ%�b}�w�iȖ%�bw>�siȖ%�b|t�����X���131?o���"X�%���{v��bX�'s��6��bX�%���bX�'����C��b�������N��M��m�-��meXٟ+Ǜr�v���kkK�;u�#�h���/N��9� Fy�1�'$#6�ەYw��Eݩӻ�-������u��Ml��R���[8�ݍ��;r��z�Y�Ah��+˪���5���iM��7	&�	��uv�bfx��B<�.�[���^�Og 0#��� ɕ��]<؝�*��GE˥tw��'�}�C�S�{�����������ps!������x��R�e!�f*��X]2����y�f��0��ֵ��ı,N���˴�Kı;�w���Kı/��u��Kı/}�^b�bf&bf-S��<�D8���˭]�"X�%��}��ӑı,K�{�m9ı,K߻�m9ı,O����9�,K�i�0�&�f�֬�k6��bX�%���bX�%���[ND��	"dN����iȖ%�b}���6��bX�'�v��2�0��Y�f���Kı/�w��r%�bX�w]��r%�bX����m9ılK�{�m9ı,O=���m�d2d-�\ֳiȖ%�b}�w�iȖ%�bw>�siȖ%�b_���iȖ%�bw>�siȖ%�b{���,�٬Ԡ=�7vŶ���|�l=�1�3��b�/�kC�Ͷf�EO��U�^J�>�~������}��ӑ,KĿw��ӑ,K��}��ӑ,K����nӑ,Fbf-�.��F�Ee��9�񉘬K���[NB���E# �Hz?�H�x�>>D�,Mgy�ND�,K�u���r%�bX�ϻ��r%�f&b���~#r���;!e�/�&bq,N���m9ı,O����9ı,N���m9ı,O���iȖ%�������f��0�"�9=���,��{�&��	��{�A$O~��&��'bw>�siȖ%�b|gg�O*Q&�rGk�/�&bf&b��zq9ı,O���iȖ%�bw>�siȖ%�b}�w�iȖ%�b~^�����T�?���|�$Kd��VG$�ִݨg���#3��m���j��<�=�n��j3k<ObX�%�����siȖ%�bw>�siȖ%�b}�w�iȖ%�bw>�g1~1313���<r!��^'"X�%����ͧ"X�%��u�ݧ"X�%����ͧ"X�%��{�m_�L��L��EM���&�r���Kı>�۴�Kı;�w���K*�"$P`�E" Q��
!�D�Ȗ%����r%�bX�g�w6��bX�'��>��$l�����_�L��L����r%�bX�����r%�bX�ϻ��r%�`6'��{v��bX�'�&�^�6�Ue��9�񉘙����޻ND�,K�}��ӑ,K����nӑ,K��}��ӑ,K�߄-���G%� �6��ff�C��-�ٞǗ3��uջ=�u�q�8`����K���\�ָ�D�,K�߻�ND�,K�뽻ND�,K��{��"dKĿw��m9ı,N����FSN����]k6��bX�'�k��NAı;�w���Kı/�w��~'�2%�b~����ND�,K�;/���@qJ2H�|����L��^��fӑ,Kľ���iȖ
X�'s��6��bX�'�k��ND�,K�k(�`�Yk%�������0X���~�ӑ,K�����6��bX�'�k��ND�,���@5�w��r%�bX�}�v[����R�dֵ��"X�%����ͧ"X�%�{��۴�Kı;�w���Kı/w޼����L��Oz�"<嵒���]���i�p�s��k�e��t�X�vͬ��ěH�o�!ݎ[9�񉘙�����nӑ,K��}��ӑ,Kľ���a�y"X�'���ٴ�Jbf&b�ֿ����R4ݶ����ı,N���v���X�"X������"X�%��>���r%�bX�����9�.TȖ'M^������l֮kWiȖ%�b_������bX�'s߻�ND�,Kߵ�ݧ"X�%�����/�&bf&b���~#r�2Gd��Y�m9ı,N�w6��bX�'�k��ND�,K���ͧ"X���3�����"X�%��w��h�
iїV۬�fӑ,K���w�iȖ%�bw;�siȖ%�b_~�u��Kı;�����Kı<��yTz� Z!A=@,D�5WI���`�8�b�{�����U*���\mJ��euȒL�T��2Z�!)̚N�t6�dMx���k7��:ن;�f��s��J�Y�aפ�v���U�����{Y[�d�Z���nEyz]xT�����Xz����&��%��򍵗�Ĳ7[ro<['������Q���vw	�����Y^k��:z����q��ɧ1b��/����Pb42�����14uѢK0-99'��r�O.�h��l�Ӥ��<��a��v.4��]d1�v�Z%��BWXq�ζ�R���Kı>����ND�,K��{��"X�%����ͧ"X�%����n�~1313�p����-c�sD�,K��{��!�#�2%�~��m9ı,O��߮ӑ,K��w��b�bf&bf-�Ó����am�ND�,K��w[ND�,Kߵ�ݧ"X�%����ͧ"X�%�}���1~1313�T�c�q�&���r%�bX�����9ı,N�_v�9ı,K���bX�PfD�߻�[ND�,K����ɟ�fJfR�kZ֮ӑ,K�����iȖ%�b_~�u��Kı/����r%�f&b��y��131o���X�IjZ�8�vySke @�B2mm�+�㞶]���ʃs�+��M2�-cpV��9=���"X�߻�m9ı,K�~�bX�'�k���Cșı;���6��&bf&b��^������c�[�9ı,K�~��� �� $_��i�7�޵�ݧ"X�%�{���ӑ,Kľ���iȔ��L�ٻ�B(��Q�$�Ky��ı,O~��6��bX�'s�w6��c��Dȗ���[ND�,K�����/�&bf&b���A��HY,�ӑ,K��w��ӑ,KĿw��iȖ%�b^���iȖ%�b}߷��_�L��L���5D{���X�ND�,K�߻��"X�%��~����yı,N���M�"X�%����s�131vk�,G%�Ĝ�o-����0�X�m�H���+ײ�N�X�I��G,�$�����_�L��L��ﻭ�"X�%��~�fӑ,K��w��ӑ,KĿw��iȖ%�b}�T��F���r�b�bf&bf-����r�bX����r%�bX����m9ı,K���m9ı,OsZ�E=	&�Ә������{��v��bX�%��w[ND��'��E`�
ā �U`:$MĹ�����Kı<����ND�)����ߐ�ªF�;l�/�&bp���[ND�,K�߻��"X�%��{�ͧ"X������ٴ�B����ӿ��=�p���aw���Kı/����r%�bX�w���r%�bX�g~�m9ı,O���m9������rS��:ݣv�E��^Lcŵn�Z�]�\�:7�h�)�:��}}[=P�;d�Io1~1313����_�X�%��w��ӑ,K��;��ӑ,KĿw��iȖ%�by��+{��7l,�S�������g�Ә�C��2&D�;��~ͧ"X�%�{�����Kı>�wٴ�Kı<�{P�WQYh9g1~1313�{ٴ�Kı/����r%����2'~��iȖ%�b_�w����bX�Ż�<��&I��m�������%���[ND�,K���ͧ"X�%�}���ӑ,K�@��ODɐ�/�Ҁ�剞�ͧL��L�ފ����A&����ı,O���6��bX� ��w[ND�,K���ͧ"X�%�~��|�����������`E-2�m�k{q
O��vkZ'ZK���<c6a�i�Z�)$qKI&�Ә������ﷺ�r%�bX�g~�m9ı,K�~�"�bX�'��}�ND�,K�����+Gm�����L��[�����?
���,K�����"X�%������Kı>���r'�J<P��^Z/��;f2�d�Y�\�bX�%����ӑ,K���o�iȖ"ؖ'{��v��bX�'�߻�����L��]���$
�Tv�$�ݧ"X�~@��;���6��bX�'�����Kı>����r%�bX���^b�bf&bf.����Vq�s5��ND�,K��ݻND�,K���ͧ"X�%�{�{��"X�%��~�fӑ,K��
����<�� �:�������u����A�ip��H'Ҟ>�<��!z��6m�@��� �9���/��`� Y D�a/ bx P��|>� h�5��ՌR0��5<x�`�!#��Ia!��{�U>)�Y	���x�ҘBE���~FFL��� a�<-�Ѱ�-J�!�͵�2M� 2)!{�4��C��fՏ�F��I�K8I/���UU��j��� ]0�\       �Sm� �� pBC�UU��Ll:�<��ۜ��g�k�]�3�٭	�g�$�d�t3�����^��q���MV���Z��ee��TI�j-Z�]�lY�kc��Gjr�ݥ���(�Dh������+хsy	���Gh�eo]n��.rmmj�8I��r��W�k0)�u���^|�웞����uF��l��&sؽ�9�.��ia�Eƶ���)cL�Ƶ�Rǌp���\��l�⸒W"H��c���z���K2Þg��)۵Ҹ�- ! 4Ԃ4 ��,s�َ!b�kVŴ]��1�;
��@�m�Wi�'���ix��!�qm�kf8w<��r$ΆtcE�:ۣ:���夒�x;aW�v�.U�'f�ڗ�ľ"�Èl�q�p�IIvt��ki�����&Jz���{j�ðҗd�vC1y����&��
��ͷ��m�va��;� ��1�j뵶Мn� �m��U�)�˸��][��-�%��^�O���p��b�Sg��5s.y{mdcF��t�G�,1�t�iЍ�%�)��8RZ��0�vbR�:�G1�; v��:�*�x\��)����0-X����ϳ�uqq�/,��s�ݭE�{Z�u�m�H�+�Y6Ki3Y<i�0/���vݵ�a숐���ݵ=s<�Ƽ�#���d���ø<�Z��yN�Nڔɫ8�c���p=t��`wc���f3��^Q�)V�Z5r�Wft��Zg5��)�y��Juؘ4�ӅS(+�'�6�ȶ7up͞G���<x{a�v*��UA��55�a�Ձs���on;��k!�
T��
f��`��8��C��m�@W2�4��"�ʘ�ͺ�r���i��IrU� �u*�g؝-�6�vMf�%�E�U9K4[D��k:�Tŵ�⇀y�jմ����y����$�ܚ�t"��E �Aãsuv�(���8oF�b�c�� �����>g����@��U4D]Ü���N3�ۭ�UUQ�t���Y�1�Q��F�)�qcH���F�����{mكa�^bk�f��V`m�K��.��֞ͷd0u���MuӰ�ݹ,��������jwmf�ʾ��5[d2r�V��z�+�3&����/�&{}l�ɳ];&R����kr�j�u3����\V���5�s�dA�X#���;��5N�B!���n��3)�[�m����{��>]���uf��ٹݲ��/6�Y#���T��:�bGQ[넸���}��������Է5v�D�,K��{�ND�,K���[ND�,K���͇��L�bX�����ND�,K�����k31�Ƈm��b�bf6{���پ|v�,�6^~�&��i!���I�v�6�6�,�6^ N���U���Ҵ���m]��M�� �M���<{{��(�T>4!��x�l� �����XT�xvZ�]n�tbb��ZR�2�2�M4R��b�$�z��xF�:��PI��U[� �����Xٱ��\�W�� ���T8��Q-rH��N��,0Z�b�LĖP;n����8߷o ��#J�J�i�V� vlx�l�?U$M��6� s�Jpt41�V��r�o�׀g�����1&�����կ����hv�l��c�=\�������>Se�����Lg6�xie�&֊�qDR���p�#ڌlWm�i���x�(��;ٳm�f�`�c�5M���U������E�^�v~iZUv�&ݶ`fǟ��\�) ��< ��<w\3�URD�y�~�SBM��E�������ih�B���."���8`d� ��Q^!�t�&ӻ�n�?r������ߧ�� ��?� vlx�����:J�vS��Wwi��l�� �s����� 7dx�.�4\�K��`x!H�g�RX�jCKe��Toa�w6骘��1*<U��j�>��<T�x�#�+��<���,^�Lt41�V��l��	=�O\���~��<�=v첕�	�ۼ ��x�ذ�r������� ߌ���ނf��\$�=��>O{��rOo������*zu�(�W�ED�6f0��bM�.U�������'���v�Or�N��j�*I��X6G�j�/ �L��;��y,KgCdbs���U֤����k��ك�9�^�u{���ۋ�����颃��e	%M;m�^��)%�/b��<jj�x�vª�N�ջ�5I/=\�r�'��ܤ��y�zz�����մڻJ�X͘�G�j�/ �r,T�r�T"�n�m� 6H�Se�#��LF WN��L�t4X�+o �6^�8`$�`�uU�UT�������󼜼�N��+Ar��U�]�v,m�����J<u��OY����ѭ��:��B�z�m�;t&��ɖ�A-�Х kt�^���E^)�#v�q���������w8M�qoh�m���`���n�#.�V1�+K�a��m���r��堞�
T�Y�Η���]�@���Z����Dk��h�cj�yW�8��.m��N)-�c�6΁���T��s�rH�o|�3P1fٻLKl���g[v�Epsn^�ָ�m��u�x�˧Iֻt�*��P������`$�`���=<�i˖�����V���1���RA=�< ��x���,��׻$=F�M�\����x�cõT�����f��;��TU�ZWv�;�׀v^ŀlف�nǀmCe�B���Nիo �ob�6l���c�� wdvշ@\�x�0p���3�7eB:#��ٖ������evS!��cr���o���[�nǀ6?r�_ ��l��[����)]�� ?w�y�HY�,���r����l��ˑ`6`g��U���O���
�9m����x��ŀlف�nǀnƪ�	Ҳ�;m��j�/ ٳ ;$x�c��&�	�nX䳀w{��-��� ��x�#�>]�wH�����=��m��a�2:�Z��l[i��h�yk��
�A�T��i�l�8�� ٱ��e��_ ����$�ww�eЁ�
���~�H����'�� w���,Y��d�����1��(�v�[x?{��6l���W���\�'���"ʨR1²%`X�H0���C��6�ɻ7�w��'~���&�("Z��x�b{�� &�� 6lxٱ�ۄ�[����)]�� ;���I'��_���wd��f����Wt��X�ã��9ݮ�l����X��V�H���ݠha�ٺrI��dj���!U��������xvK��U�|���<O5⭺V�d��x��o?�HB��l��Ӌ��z��ݼ�ēf�
z0My�n2�l��+ 7�< ��xٱ�v(HM�����*�yfc{�z�w}x��o ��b31#�0�$,/�0X�BXvm�\���QK�B��ݏ ��~����ߟ@����{#��e;hwI�cO�ُlܣ��v��N�c�[�e�c˥��fa��r�1�n�U����� vlx�K���ܯ�g��y_�ҫl�E�wm�w�أ�� 7v< ������d���Y�2X*���u��Oߞ n�x~�����	��xɱEmRPd*������o��� ;���w^��,ı��x���R�:�q'n� ���UU~�+��ߗ�����ܒ}��krO�",
 ��R! @ �H) `AH��HJ!D�0��s3ZՒi�4�e�d'hKz���H�Z8W��v�XlvA(E����Ȑ��kV{&���UCc�����L�r;��u=Dk%���/�v�;\Ai��b�K(ےx�ȦA�6�cg5��
���m%���;e�-M�+Y�m�';\��͋�FDt0�ud� v�7;�t�E����0�x{��Xu�WC��^��Y\-%+��%Ջ���X�q}">r�����������Pѱϱ�,�`����˷nX�l�)-�0��
�A7)%��=�}��M� $���U|�-��-P���68�Pv� ~�����������Y��$Iv��eЁ�+m���<Wv^��+ >�+��1nʫm;Wm�Wv^���������M������y�ԗ�ݶ����+ >� I#�>?}������\UڳA0�c-�;^��sg�O7X2MZjaZYZ�Gh�+������%��)�.���m���� $��vK�6e`&�K)����Z�krI��}��Ċ��,�+@Ŋ`h@�v?!�B�s��.�vw�7 �۷��f6{v�e�n�8vY-��X�L�?r��&�� =�y���p�����V�X�L� ݑ��<�����\���,�*����pT�uAڸ�����,�O����;��>�7x��Y��۬�lh���x�۱���<]�a)�nӣ��}�r#9㑅�s�6�Z�C�ն�@?~����"�6e~��'��V��bN��m;Wm���Y���'�{+ $�� I#�"�WҥV�Pƅn��7M�. w����s����f\KSUuB�C����#q���X� �X��	�pH��U!@#YFI%R%�(f�C�+��Y�$aR)��H�q���X�RN�1�.B:�b�]]��a�� �b1 ��H`�� ��$*���1`1jB���LM�������@1)��@$�R�m��Ҹ��0����i�y"���s{	%dH�T�V!B A�7���a�����������49Aʣ���la!diHѬ�T�a��-!Kt�)�[2"�H�Z�@�B�
�]!��!"b� P$�B�c �R\�r�x�5 ��6�6(�6���CJ�Z�� (�E��J�]1
��)�T�8�M(����G����X��	Q�S�R&�T��z��<E6�� �C�be��}��<�n���f̖
�D�)Kj�{��� {���;.E�l$��n襔5v�c�V� I#�?r����?g�ˠ{���V n��RK��?���������X�{
R�e\H�$D�W�e$��2&V�q-��n�	�%��識�t���{�����^��O�A7n�6���Y��r� ��x�{� �����l�ֶ9	��uAڸ��� I#�;�"�6e`v$�n���m�q/{�x�����l܊���!�*����2?m�gN�l�'Hݖ�ݹ��+ ;�< �G�~�Uw��R[��5B��Z�,�Ҽ��T8A��ܽ���3;�δmq��f�����~8�ݻY�[����e`vG�H��ȸw��2X*���-��wv�عI��<e�� �I���UI$���X�VR�Kx�{׀}ٺ�%�$��{+ 6{� ��T�;V]��ۻo���,x����#��+�W*�������ZC�5���n�;_ �e`vG�H��Ȱ	UWEQ%T
(��Z �K2
`r^i1�/$������UUUJ�#�.(y��@2��tP	�$����jK���&e�\���桨�z9�������ը��x�	�Σcv�t��ǔ���g�aV2Y���l�ݚ�[6v:q+g<������M��j���7v$u���9]���p��ڀkU���D��gj���ʬ��,Y�d^���bof�N�abX�mӫ�A�SA��93���sZ�L��%�$�d���F��¼��B�%ҥ0���\����9�H���N`Ԁ�����z�Iݹ�r�A<{�Xw�{t�BT4!��x$� �܋ �I��'�����?" fO�ݿ�ܗ5�B�ZN�x�����L�?UU$��{��o�x_{"؄բJ�,�����U)�/}X��x6G�wnE�l�Of;Z"r��ڸ�wo �K�fb���ߟ@��ߖ�)��n���T��d�nI��۟V�s�5��)�e���V.���%�)�qtyD,J�]��m���wnE�l�e~�W*�@l���F��+���,���;��Y�i4�s0�6���	���#�C��+���''�����'��u�	�<�����r�"�M�[X�L� �dx{�T��{� �s� ��[��q
:�v��%�������xv�,ܪ^��}X��+cm	PІ�m��ݽ� �+ >���>�B��!�*�J��X�؜T�xE��r�)a%XMn�^ײ�`|#nh`�� 3:�cI�o �܋ �+ ;�?|������]5WI�P�+v�$&V wdx6G�wnE��������4�r�����z�{�x$�fDƬ(�)(�����'�{>ٹ�ݥ,�LE41�V� M��nE�I	�����%��<ލs�ڵe���v�o �{�s�������x�wo �,M}���peM�q���f�M��5���&����5��Yml�@VB��>]�P��%m|�=���< �������>}k��M����N��	� N��	��`kfV��D��c��hCI�����	��a�)*{+ =���'7e��JݕC���6�,v�e`�s��*�+�$�Z� $"|Z�列-�HI"�Ʀ0Kl4�nI���#��vo' �����)1��r��z��X從��z��Ȱ��9�W�z��1��O=���/N�;�mn�<��:L�05���t/nQ�.q֌�.;��7�� �I/ �܋����z��+ 3���q�:1V(����wg ��u���+ ;6<���s����9�B�
˻L^������{� ��e��#:�P�ԣ��wWw��ݏ �6^�nO^�B���+��;)7X��x�����eo�7$�:#�
�>�f}�֭� V�ΤK�܍rf�k���<��iV6�n�n[��9�q(�����U۶Y���q�h�ٽ��6�j f�f���lb^]	�[�2���%�z;C�
I�tv��5oE"���t��Oc�tm!�cb`�N���*��H��	�3��I�Î��*�M���rpNK3�΋m��kr ���|�H�j�M0qIc�(TI�K�.����#�\�Vg���lk��ᱧ���t���v�ӛoV��7a�N�IG�U�:�V;n�����-�x�ٕ�nǀNl�,V�Н��>[����+ >ݏ 'f�b�Ϟ��X�V�-	,��{V�+ >ݏr��^�����:�rJ��q��ԕp<�f%�'}���{��>�ذ��+ 9;�+��؆%WV� �#�>�ذ�&V }���M��m�A�JG�!�UNI�nL�. `��sZ��m���y�Ӓ���̟mʼ]'�M�@�_�,�Re`۱�[%��DQ]�6�m`ړ+>���(���z�=����}�ذ���H=����N���wo ��E��K�s� �^�V�֨^;N�J�Bo������ߖ���`ړ+�$����%Z�ҷePƭ[k ���`�U��S���k�����Ȱ���&R����f%�NY�m��F�ק��g]%�&^�;;V��n2Xdn�M�	,m��Re`wc�;�"�>��}�܏5�V���Ƥ��w�y�f������ �ԙX�����1*�i��wnE�}��㯫��ܪ��vpR��;�8g(P8/
���k�s�T���r�����>�/m@�.Һ,O����8`ړ+ ;�ݹ�A%%eЊiݳ �ԙX���U�{������>��E+�Jt��%�n$��6��m�xډza�l���$�OlZ�.�u��^��;F��`wc�;�"�>���r�A������w�:І����ȳ�RGg��e{�X�����s������`�J�-�����>ջ���bč�� �{׀|��ull�!���0ʓ+ ;��d��Y�
�!!� ��w��n�w�/=mRV�N�]��ݏ ղ^�^�Re`I/,V�BM�$�v�=����t(�me���Y�F+7c��Cm�Г��ȑjeQWm���� ��vp�n�ff/����w&���q�"N�M��]����o����ݏ ջ��ٙ��fk��"�knW�;��e`�c�5l��|���"�|V]*�i	�������%6y�Oz���x��U\�_�v�	(��^1�hBN��5l��|���&�e`�c�MbF� ���R]!�!�c�$d� J��A+/t��1G�\!	�~dxa�3H�2� !��A��T�h4@,��	�(ˡ|
zI�y���%G��y�h�+���`��5��hJ�H$`��a��0$H��譆 L>���M��H�2���R4tm��l��ff2��L60�&�������0B M~_~ WZ1�8�C�
^�Fx�fb��Ф�D���)���R���`�]�9����A�!6�!�#���v���ٳa$ ��$@�4�M�	�1� ���B��Z��o�j���he 10թ+���4u��	��y�9d�9�^s���r!�k
   鎶�      �m�  ����	���A%�z��dkf2��[9��ٷkP
���Bm�l�<���RMղ��_W�� ��� ��g��C��MlD�7i�[c3lA����ձv��UA���9��:����;q�i"��m�,j�Mq�	�&\�rpMq��jgf-ts�����9رC�csc<��]>`=��l�����M�<0Ԍ�n/=����ug�A#d�a����<n�Km'�Y�	fV���2nw�f9*x��c�v�bwj��i[���<sA&�1+��qg�}�X�=e-Yj�1Ȩ�o]]��tz���'q���fG;�8��g�ǥ��S�Ū�g]l�ښE3����k�6�7!s�3�6nu[sG[�VÍ:���h�k��bT1j�yDؼ�a�as��*[�n�K����ݫ=9	���5ĮΪ�Li�3��n��]�8�`ܬ�<ivV�P��Q�����\�v�$�m�hL+#cni�+�=bkA�v�s����! ��6S<C��Sg�l����S��R�%<�tM�9Q^�Q�^�T�k%by���h�"n��c�g�˛������2=ù��2�Iʛ�a�;��V�s7n�<�rn��GJ��Ƌe�k� k��[se�۱�4�9+6�`mx]�9�!�{`��bɊݍ�����d�
u;�:S��PL#n�a�CB��K1T����⠂�[,C����B�TR*�W���'T�ut�:�=�E�P�M�M�����bP�8�+�Cn2�v�ۨ���5&�
�ŭp�\���$���=��y��C�� �2�X�p�=�9�t5����Wm�T�l��R���HV��������ix��s��cv.j�QXB3 m���$-��O문m����t�9�����:�k
2�W)`��'�մ��ӻ"�.����1H4��2kSY���*�M��#�m6(x'�!��H��q}�'�����j)E��A�E
D�+ �$BX*�H�8��+�����O}��4��M�e�wn%�҄��/ݰ�#ڷ�L�V�ݷ�(Ej�YSP��Xy�Dq��n�rѣ]�B6sPq'SU�+�ɰ����d}l���u9q�<��g�4�a\��m&�i��%)�Wt�dL�؜gB�Z�7^R����{�c�h��񉫞$j0��f��e�a�D/Vt�7*s�����Ν�.�4��9c���I'9 xy�fJ�F�����fQ���P�9�R�f�sts.����SA��f�A�Nl�6��D�)�ym���� �I����ϐE=��:�Eu롖��
���&�e`fǀj�' ��u��g}�A�ei���jKX��x����Ȱʓ+ 9��nD�S(ڊ�o���o�8�{π}�w����$�o�Ӏ}ܛ���bt+�� �܋ ��s}^����=x_wg �{�#�[^�2�9$�طb�)��rr�{I�XU��c6�Y�b�֫��9|��f]+�E"�ݷl��~���|�K�:��?�3?0��y�?l�����V4nI���|٠M" �7=�;xT�xeI���#��Ǖ��4!�ۼ)�^�l�����5M��NnԳ Nʦ��[w�j�/ �2�Se�z���z������Sl\CaNۼ�+ �UR�=�{Ӏu�vp/��G���K`:�S�M�m�v��p��ȗn��E(�ޤ�vsd����{}*�\%�i���J����Ӏ|�vp����Y��o�{��}��;*؛��Ix����S+ �;��ى��d�yǎ8�:�%��k��7$�ߏ�nFUJ�E��u��+.$bLM%�'^�g �wx��:ε�6��;h��X�|��p~���L�s�W/���^�����W���Ī�`���;$��5M��l�x�vwcn�ƣ�� Q��U�P���6h�p�2晖X�R���zrR<r0���v�?BL����o��T�x�L_�g����s�= �2���ʸ�����9ʮ$Ox�V�� �+?�I��y�O&�.2��Yl���� �6^�IO{�X��,v��P�cT��-4��0Se�$��5M�7'�x���D�*��w�&��vxM]RLCE[w�vI��j�/ �'T�xV�v5g�2�]�J�^yݲ�v2�j%3�n��|
nl�b��S�-f�T�\�<q�A�7e_�������T���������y���x)&�
��bp��RD^�� ��e`{�9��I6{�����`8��i�"��xvL�?Us��^�� �x~0�)K���!��xvL�T�p�mӁ�����zpgt~�	�c-۬T��վ�g�������� ��b��dX��������Z���^6�lm��C3�U���r�gxu����pl�nuc���n;[��v�ݝ[ITq��L�P�qm�1�5ݺ��,A���hx�=2��Z3�Q��AҖ{;\�ֺ�n��#Ŝ�mƀz�xZ�N7�����WǂI�n���F�禲#���b��0��c��b�4����t�0�h�D�]��9�7XM$�D�̚��γq��B�[�k�ˡ,#5��嶠����f��G-����5E+�P�~�T�x�_�Y������{�P��,+c��ƣf�l�vL�f̬i3��ăJ�y&��;�4U�7x��V�fV�UIz���/O^��"�+*�]�'BN�`6e`�8`����'���.�gXh3���mNZ���T��	�e`$��?W9ʪ�پ�P0峚�����'����yuRjf�
𛕕 Z1�����ڶ;�g����/o�����d��6I���_ �W����~��n����p�n��2� � 1D)I����<�j{��ٹ'>=��p5I/ ��`�q�vZ-�`$��;*8a�%���$��wmEWqc�,j�Wn�ʎ�%����;��\~�֎�ZnB;���%������'������7�[;�t2���m��l�����c�"�X^�t�u�n�P�	n�ob����7c��fV�Q� �6^���{[���A�7m8w���,l�W��/O^�0�jT�(v�嫀}�n��{��O,̙s��!H(�VM���?��+ �W�ҩ�V��)6`z��O^'��f̬����b%�� ������ ٳ+ �/b�5M��Iݢ���;m+�S�ݸ{7�7���F�z��=�Cׅۣ>��+�qTIZ�#��p�w��uvw_ �6^��j*��h|E�*)]��6��,���y0;�?�]?��H��@U�CI]��N��"�=x�8`6e`[{ t��N�;@�V���z�ʪ^�g�z{+ ���d��E�D��5�����<��_���]؄�N�0�2�	[{�l�v8`�URݞ�I�M'v+u������P�$u�X�5��9nƝ7n8��Œ� x��daA���;jr���_�����X�����r�A�{+ ���W�)ZB|k �6^;0�2�]������|��,�Z&�Q�g ����6l��&��`���>�DR����c�l�6l��&��`��8O{�x�l`?zRc%h���	��XV�{0�L�Us���;��UUTL�5&utZ���1^ܜ�i�yv4S0�%���.ݰZ�I�x�j��H%C��
���+#'mӜ���g2N�1g��cח\6�R�D7a�b�a�gv~��尯7en��'�"���:����\-D�\b�q�3��q�X��=��%��W�Tn�`2��u"-4�["M;-��������v�&,��3k��[���U���O9��h=X�r�1�b]��L�f��5�&Z�KH�j������<u��`W1��5I��7�� �d�����=�X��� e�[-��7�� �d��&��`[���\H��yxj�E��'Bvـv{�X��,=�븽�׀z~� ��F��8�n�n�	��XV�{0�L�i�;A���m��v^��+�����@�~���J�ذ�ԻB�>_�wLou˸׸3g<���0�q1���/[zu�{��:h�x��T�M�Q�g ߶��?ww��J�ذ��x�(�+(�,�;�!�Z��s߾ٰҤ��G
T�V��sA���P#Q�0"�r��@8+�<}�H�w<�)�^;3�+�������U���BJ�����>�g ���+ ٯ�K�4%wc);kܪ�Uʫ���x���0�L�i{ B� ��X>
������&V+ob�:�e��ͿK�X��۠��G�w=p�{.l;�eMR�1�!�-n1kt��u��rs�͸��5����o�n���i{ջ/ �� ��F��8�n�n�	[{ջ/ ��N���\�f$�=����<�c�6��O^;0UߘU.�>U}ʪ(uXG��L:���CI3��!P	��O<��l``I��ie0!���7�T��
��H,`$������L�	)+���CƁ	)�ʻ�|��`x1R"�c���ƒkjF0�� Y  �v����<Bf$� �H��o�X��4_6���e+��e@�B��X��ئ�	3[��"D�!F��CI����!���dHC��|S�S��x+� ���=�Q(������@<C�#���, Gb)��U\����e�,V܋ �JR�ۦڥBucۼv8`mȰ	[{�,O�wӀ}��qV��m8�r, ��ջ/ ������!�Wn��nv��P;�,�=,b���e�D\מ3�BA�S��lgM� ��ջ/ ���W+�������Ȟ:¶䅭Io ���9��ďo���{׀�c�WdN�4��V�n�	��|�K��$z���:�}8݂�Mq�DG�Wi��X�n{׀���:�e�gy��PS����i$$ "��<�ܒy'5Q��
�ջ�	�ǀz��'��7��8����>z�D7&�m����,	,eͰ4�m�-Cf5%,Cb/.�%�-f�E;@Ê��m��v^���d�V�ŀ}%)�ۦ�\�1]��'c�{��~��}�,�=�� ���9��K>��'1�AB��m0�����/r���=x�����(�j�ؒ�Zl�5J������� ��� ٯ�K�5C��ۺn����O{<|w���T��NjC��yˈ��}ϵ��֤� �)�Z��N��4�>z;cz�_�}|8��bԻ�c��ׅ[WR���t-�,s�N���qp����'D����]!k���s�h�*�>4rL�@&�S6Y��C���cG3E��- i5��0��%WM�i�\n&إ��g���n���u����F����&�^��i*����{FH�k�)2�B�k��ZܷMV.5	?rs��y��
��Z�x������;&�f�&J�F�ѭ'�f�ZW�,�Kr��9K,�n��ȰR��-�x�YWq4��-ZC�jـN܋ �*K�"ݗ�l�"\��U'��:k �*K�"ݗ��S�~0m�� �sS� ��i	����W�O^=�� ���T��}�)L�m;����#����{}�>/W�x��xwuqJ�G$�U�b�dDl��s�=��/:v�{b�5�s�&�n�����uv��0�0R�� �v<dp�;K��[��'wE�ـj�%�x�$��`kh>�DԜ�}��=#�}ۑ`5Ղ�C%wm[T��{��#��ʮ%ݿy`z���N�k�dYpqG-�yg�%�}��6_�� �T���ǀou�wH�-!�jـ}ۑ`J����x��8��"5�UuY ����[\�x��{v�-�s��*��'V'����ŉq�F��>`!�;+����8����$���UU����!PN�A�⍎�Գ�}�y�Y�7޾8_}��:�n�yf$��Hi����lu�X2�������=��ؗ�1q$c`$~`U$R|��9A�w����;������'2J��de��%���z��^��ݑ�#��]����ȋ,��u�ݜ�b��}���~0���9]����I��Qlut��vݱ�k��]5eݺ�pޤ�wmI�m���t��i�8��%�&H��m�������w��`�Ixۊ���4\D����9噋?�%!�=������� �����Y��ݢ�ζdR6F����,T�/ >� �0�f�I���_�$��z�/�������ݺp7���"�X��U�M ��#MT"@�n	(�y��M.,Z�~7���7�h�#V��j�� }��8`��X�	x��I4&;�T41�G-n���MY{.6���ݷW\O�zvg�Zj�����&����������� �!/ >� �	.�YI�v�ݫM6`��X�	x�dxdp�;K��E][�2݃i� �!/ >���*���w?~�{��l�˥Ȇ�wm[Lw�l� �w\0?bǳ�=8 ��~r̀�."Kx�8`�Rg�.��������x��.W�������Y!�4�e�d[���??k�!.#��%�	㚨(U*���D9 @as+�p��]���^ݜ��6f��'X'��J����,��V �ZiGn4�N�[m#����n�Θ]�՝ntcɭ�Vɑ�n�a�wf<�:�|���ͥK�]ngr��t2be����4*�.F�a���c&|c��!{,��E���.��c9�.w!b_fNr�@V?�rʤ'li��9�p��s]�86�9��nc^y�۷3��m�o]� um[>e���?�K�O_����,K�{o� t3�����cvU�E+e竕\����	=���y�0�r,�)#l���V��j�� �v<Mp�>�Ȱ�l�t�PZwE	�cM[x��}��E+e�{}���ho�|��Ide����[/ 7��\0	��E�׵\�k�lѲ�KX5���I�s���6�Ʈ�):���gtf��V֦`�l� ��x�p�>��lۑ<�PU�J�Y��ݼ����f�3c�\0R��9��$�E�n�`�ui��o��`v8`�M� ����}�(��!���`z�w}�0��׀�ǁꪥ��x�EA*��'i;k ղ��{���� ��"�=�wHg��IZ���q�rwa.�l%C���\I2�Z���;�h���fm 4���I��G���"���~xdp�>�Ⱦ��j�I���),MQI;�V���}{� ��Ծ }�v��1��z�V�,��Ny�w�rOo�f���!��@���*� 
O צ�}e�:�	��}Jq��o�I�m�X��/ ;ݏ ��ʪ�?W8�w����=��<�eY$�[� �� ��o��>��� �!/ �W�a܋� ��u���͗�E����d":�,��v��7CX���!�wb5�y*�;#��c��B^ w���SiqA�R�N��s�bl��� ݞxdp��UI�"��^����$ـE�� �v<�8`v]8�],Ѹ�u���ē~��u�'��7$�k�?!ċ��R!�=_E��u�w���'>�/Iwf��I؆�����}ۑ`�%�[���|����]�:�L(��J�������c5�M/(z�[.���U���zn��whm� ��T�� �����f/�o���8Z������7h'm0R��RA�x���;��|�\�aMvյM� N�x���W)/l~0�^��TZ��3�4:զ��8`��j�%��ǀou�VR���jـN��T����8`N��8QTUT CmR�`�x�]�ݫ�|6@��Z>��hR�|�d�xy�11�x��=H� ]�!�@�� H�"T����",aVB�0����y�I�g	3��|�E�6m"ERn˒����!&��׺0�d"@�X& �(@ 1`1.�OU��p�p�	���0a^�Ċ@8��(�#j��kEp��I4�(�jHa$s�bFД��:�x)����qA��FF!F���$�c�3L�@�P�		��vm�.�I��L$�u��fx����JHC�5�1�
�eD-!�$���
�4�}�{��,X7�}�s�FNOx���U\�UUU  k�4ڀ      �   A�h��(�UUv��(Ùǂ��W����P+v3�$g�-�sX�6G1f��kvp����4o(ly�l�Q�bS$�	��n�h,����.����s��^w:�r�f�*��r��z�L�: �y,Fj8Uw��:��r8*C�y�V�R�� �Ag�r��1��m�(B%��iX�B��L
'�Ԫ��ר��	�v�8\�SFE6�a	wl����y�y����̫���3�sM���H}�rg����4�4i�ne�v�K���;gs���;Z 9v�q	֜�36�!ع��M+��k]��lq��8��m��ݹw����k�7U�l�X�6f@y�ns������.m�G�6�[�6��ak�%�W�l�u��pxq�3ۊ6n�Cb,�zd�pFO�����N�K�����&�u�mۍ��k���)稱۳763��v=@��9�nLg\cѹ����nۦ��Q��V|���dFS��܉��m��9Dq ��p�nTA�8���9q6��g�ه`���[��4'`������&I��u�Wq��6c�6i[q�V�bm�r��u���Z.7bs%�Q���"�by$QAƢ*���+«�z�kYN
�덆y��#mi9B���N�9�P��`��]Vl��ݎ���r�.&1c5���j@1�zEyCg�%vc�WqՀ�'�4�Z�/<r|U��ێ��Sin��������A������H�{T�y��{#��ь�Q���]r�a�N`	�O;n˹۝��Ẫ��J�:њ��մ�
�\>����v��ըX;{v���DRt �����͝I76H���9n��۵��rC,��0ն�f0s#HՓK�#ќ�6IͶp*�J�ծG�&�t�/�e��j�'d�9c;]��v��\���y�;]�v��˜9K$)�X��pm��P6�5*��{�/w|�:@�q���D`���(�!�Lz��u� ��rs��I�$����������UUVvW�ӗ<ݍ��7s�4��w',n�#H/f�Ȼ��{d�l��ٺ-�E͉�������{AVm�����
���[�:8K�qݓ��[g��ao[Ӌ��P��	�U�ᐌ��v��DF�;k�ϖ>76�n�' ��Q����grr9R��R��j����0�N6��PZ����F��g����vqt6G�uVc����<}t��l(���^H�(E�Ivf�tQ�SQ��[m�p�@4o���R�!؛��?i�8;���� ��iZ;TN!ZBi���ǀvGw\0SM��$�>�'�>2�Ӳ6ݕ�x}�� ��?��W)(��׀��N�����M�E$��0	�p�5HK�	ݏ��{<`U�~��()&l�5HK�?/l�����w\0�����i�iul"C�JC�k[I�z�;sF=DSۗ� j|�����ڶ�� 'v<�8`��`�%�TZ���RM�ui��vG���#�k����d�g|��|��Ӏ�v��1���(��A8A:��ـ{ny`�%��ǀvG �sPV�K((N�;k �!/ 'v<�8`z������T��=ĕ�M5c� �����N�ŀj�l�?�dc�U�rJݘ��^B;cGQ� �0uф	h�oV�O7o驲����ZI'm[xdp�'ob�5HK�W��l�ߞ��׉ݡۻE$��0	�س�*���H��=x�xdp�U&|׶z
��ݠ���~����ߵ����EL)�߷���oӺ�w�"y���$���g�$���<}�� ��� �!/ ���,Ht*Q�x۷N����{�|�/x���ǀ|�.Z�n�+I蘧%$ц�P��ڴ�-)�B�[��v�N�Y��ZrU��) .C�@���Q,���7πj�����0�Z$V��(Nӻw�j�����n�<}�� �vK�&����T
�MX� ;ݏ �~�R][�^�z��Ҕ,C�*v�I�V��0�d�����ܖo�aZL�(�~9�~ǀwCe��!7i�l�>�ȰUW%�ǯ���vG ��v��4a��ݞވ�Ϸ;BgIs���=����Y�K����n.����ZQo-�����ޒ������|�%�5Ղ�E��],��wo?�I&���� ��ޜ�t���X�ּ���ćB����w޾8�����1$޿x�����:�+l'�;T��ـ}ۑ`�%�{���� :�F��4v7e|�t��?�$��w���?ݹ3����.ݶ�M�lnΤK��.A�����P�M��Gn�����S�-�6�����1�#�d�Q�s��\�ģ�Ks���Q��ዝX�<�vx7�s��ٝ�j�v�U1�.w^��	ʕ��m78�w!�-�)	����COf����$j��Ͳ/M<fc�T��S\pNع�@�v�A���8��K��\d�N���6��o��o��$�؜���{����[�$����ۑv:�ə�Q[N�u��^]��\vͬ��n4���;�a���I�vG�܋ �!/ �m)X��V6۲�o �v���%�b�R����<�~?^ w�~�${C��ybv�	1���~��5HK��c�;#��ˈbg�b�m` ��ǀvGs��������=�ά?!�ۻ,�X��xdp�>�Ȱ��XdS,M�i�����}�v�u�˞ݦs�x���2��\7k52=�kBOnn��bC�P������ ���|d&V w�ա[a8�N�rS�~�n��R�]Ř�&�x���׀vG �iIATLI�X�L� �v<?��o��`���4��H�'n�������}x}�� �vK�6Be`M�0���BI�V��0��s���=��X����>���+�G,��"t���8�:�s͇�:[�.˰<b�nn:�-��[E��M��$��0�d�d0����ݰ��?�w��~��bg�b�m`��� ;ݏ �0�r,f��S�b�ƥ� >��xwn����J$>*�_AN"�v�����_ �.�8�k�6Yn��≷�l�ݹ�I���Uq-��jЩa�q	ڤ�v��l�f�+ 7�<�\0�˺"�t�+�v���Ͱ�`vX��zy�;�n�z��[.�Ɩ`���jgym��^�0{#�;5� �/ �s]���
V�'e�� 7�<�W7���5zz��L���)��]&�Nڶ��p�	��I���<@�w�-X�%��y%��7��^��r ߷o��Պ�"�c�X$�����~Ė���u���Q��ݣo ٳ,�	��� ������}����$a��"�� 56�۞���Vf�{��i�"�j�c��%� �z^����+I�V����<�7c�6l�0�V�[\�'C���6���`n��6l�0vG���$uo	�f9u�N���;��C��<�V�*[J*�E�i�ջ�6l�0vG�w��������'�����q��$����x�׹'��~��=�߷�rN�TR&�X,F(�0Jc^�$�ж�m��+,t��=XpQ��jP6�ظr+@s�v���۞�,nE1K���jƪN'�qL�^�����1�6�l��-�5�ܖ�Y��N�k.�]�W���NL����)&�̜�����i�Ժqus�Lc[���۬��z��n�ٴ]��5�f�գ,�/��&��N63[F���8�N���q�.gA�%ð�N(�j�Y5���OȣA��~y�-��u�9������,q��ϚǗm�CFk+YF�M�-�ۡ6�*�t3�4ͥmɗ�����f̳�>@{}�{����j��ul�m`n��6l�0vG�}/b�>]$!7TRI����6e�;#�>��`n��'c���'�t]��+v`� �^ŀE�'��ߡ�<ֽg�yu7Tv���� �v^�fY��<қ6��38�ɘ�iM��tʃЈ��jٸ{s�֍�1[ve�Qa'�{X;��k�������Y��l����}OZ��E\��w{��;��,�DD���,d(�T"�R P`��D(�T��%ĒMb om���|_{���1&��-u65�	ƛ��À����X[���2���S��N��&�����X�p�6l�8o��� ��ޓ�H�X�$��	��sޞ�� {}�}/b�;�-�׵\R1i��Ì�-��2�{n��lp��[n[f�Wm��f�ͫcm��V孀I���<�{7\0	��R���v�j�0vG�}/b�&���(�U$yTQ��i&��ݷ�}�|{ۧ�	!��B��F|��؈z�]l*h"S��y�M1��y��A�#��D����C�R(�#��2(͒� ��*O7q�����ఄ	)�B�9�'
.ox k��Nc	�$ �#6���(�,1 `���HD���@�"�F+-������i�z"m�B$<��dҦ�iFB,H$FBF$xr�O�_u���2bB/��/6���@��7�����&����"��oG�D M���u���<a	4p=��C��� �! ����GZ!縚G!&h�k6�1��p�@�޳��ġÂBF����8���	��Ls�=��}�p=|�4�j:`��|���xX��{ =GH0����C�""�.� 	���@�&(��X�������F�� > ��]	��(�
 z���}־&䓞������Ѵ��eR�_�$���l~� 'dx�9��.��,�qqR�^Uj�He� ��`� �^ŀM���˴�M�-�N�3���I�[��)b"{��J���mm�0�L���T�)Z��ݷF N����Xݺyb_�ov���:�R�� �m[x��,n�`�r� ��竉6{����$V�,R�Z���^��(�	���� �t����RI����ou�0vG�}/b���ŝ>E�0�A�������f&_~�x���S�b��Z� N����X7c�7�����w��充#N�{�A�����s��`t�����k
�7n��P�:c����Ui����, ����G�\��l��>�<�I�U,��~��yeRD��F {g����<�ݸ��]/*�E�2�m�c�;��Kذ~����GTm���M�%��{*���<������(�>�Hr�U���j��>��`ݏ �ݺ� o۷�%�1���}�F�j����\mt����������&�18^Ć���n��#ۙ�6�R磜�Pmc@�9��Y��x���f�V�fKB��b��ùܠ�m!�a�6�rF�����7h۵�qsŋk���v�\��s˸� �@еFgV�3T���[�[K<l���t#���4��6
����,&v9�Vt�� ��k�Ph��H�XY`7�YH�Y�I}�I�O3o�=LU6�*�[���*�sM���#k��<�=q�n�wdmæ��б��ػ�e�k ?{<{�Q��<�{�� !Z�|)$����7��;#�>��`ݏ?s����J�N�b��Z� {����w_b��n��c�Z-�F�:$��o �^ŀv<{�Q��<��WUJ���ݵ�v<{�Q��<�{��I+T���ӣ��v�=�j��q-�g�]�'6���q'bN�k��8�]&����o ��`� �^ŀv<s�����"�)'woDܒ}��k{����|�:�Uc"y��۱��r���S�J��h&�����x7c�7��;#�$�^Qj�(.�m� ����r� ���Kذs��^BE�\*�n�6��M��`� ��������ŝ��#�m:����8]v��ϣ6wf5�G�M u<=]�zө����8��U:�C��KQ���� �M��v<{�Q�E��tY���'V�x�l� ������ 'dy)#�xJ�IU���	ۼ ��[�{|��7:A`��|
��`�`T�<�E�q��hEd���5�'��߳rNy�֊�EV���X�x���	��/ &�x����
��Ye$���vG�|���	�KV�E�I/����7k2�]�r3iKBnnY�b��׎V�Ӯ����pe7S�6�m�De���^�� w������� w���w���y.!v�2�� M���$���w�I)��$�n9kI{�t�B윳��_} �o���d|�]��I$��|�D��P)Dc�69�� w�z���׸�-��}�\�HX�V�d$J�,� tڪ" ��]a���| ?=���bKX0�}�ێZĒJn���$m��$�����A�Ns�N����eMYMvU3��a9뉨;rl��M�l�%�ܴ�l�uƍe��	k)Y�2�q� w�Ͼ�_�݃� ����ř�ѷ�����o��x�x�+ur���精 }��@?n�ύ���ݿ�{2H��V��?&B	�Kn��$�������-b^�9wk��<�P����ߺY�t"���;/�$�n9kI)��$���5�BSv?} �m{����av��i� ;��}����_ �}��@?uz NI��K�g'l�����ʶUUUSS�&a�3��UH���n�z$hS*H���r�ᤶ�y��:P9��s�]�y�;���Z��.ԫ������i5�v���e���rm�����i�=�7h���$`��us���Z�ru�ny�k��.݌'�ͷy�\�5� Xf[f,�v�F��&Y֍��]��C8ƌ�����p�370��q[]a�f�ɬ���4�|��ʢ�=rI��俏�r4��E�	,�ݝ��u���N$9�O�7Q��z��|�TF�k�yf��_߀/�_�W� ��u���^��P������G����қ	��� w���C�W�� w�z���精 ��0v-!X0�����$����ݒ?P�$���|���/ӭ)i���S4� ;ߺ���}�� �����~�{� ~~8KN�+u����c��{�_} �u�� {�_} ������JaP�.%���{W���g��m�+qe�Oi6�;d���mU���lͺau�r�} zy��IuGĒJM����H�=I�H?}�Y���Y\�L������"�v�qsN�X��'`!�خ		"	��@�~ ��@�����?k|�����Y�m�ϻ��@;�^��e�٪�� ?l��Im�x�Kod��I.�r�$��ޗ�.��0,�U����c� 6�K���ܗx�IvH��$��|����i���w����{��ݼ d��Im�x�K�zy{�&�n���W�åe�ZH��lm�cTԶv.LZ0pݨ�Q��a�&ج�!X0��|ݿ��o �{��@�ݎ� �}��} �n_�P��K�2��� �������c� >�w��@?�7��~8r�x`��W�@�ݎ� �}��}	�Y�
��<7��s�7m���{�r�~=�7/e���X� �{��@?�7��������x {�����6	`7e=���x �޾� }��w��=���������Ș2�/s�'l^���t���'c�#�N˻lγ՛���bf���1�lf�M� }�����$��S�I%��_|�]W"�I%��)H�o,���]����x }�ޞ��n�o ۽����G����%69�� ��=���x ~��w��o���>��0�a��巨(����n�o���9�m����r`61�-K �A#KE�J�! X�)D�2�
J
�}�:��^r�|n^��!n��̴]� ?n���@Koe;Ē[�E��%۹.�$��.�X�n�D[�Y6���8+I�Ao1:�{����I7vmf�vt���nJ_�$��S�I%�6_�$�n�ĒKf������ZN��X��x }��w���G�=�8�m�����}��g=�H���R,a�K���m���� ���$����Ē[���% \ƚ.��:䤖��߱b�&�}~m��|���_�{��}�x {��vK.M�cm��I�(x�J���+��O-ԕ���j�m��=�9m��EW��A_�� ���AZ����EW���EW�� ���T��D��E`�AH*T* �A ��`�DX*
���H*��E��V*�X*U �A
�T �@
�E�� �A"�E*
����� �E��
����  �D`�@X*  �@P��
��P`�ED��B
� `�DB
��� *E���F
�A`�ED��B
�*��*
�X*R
�
�E��EB*�E �E �� ��  �DD*B
�E"�R
� �DX*
�
�
�� �@ �@��
�H
�
�X�`�A��@ �D �E`�@����B
�UR
�@��@E*U
��� ��D��B
�T
�`�@V*�Q
�H*E �AD *PH*�EH
�D
�
�H
�E�� b*
�*��B
��E��"�
�F� �A��F
��� "H� �H�� �H
�X
� �H��X
�D�� 
�b* �AP * �H"T�TA_���*��DU����EW��"��A_�����EW���*��DU�� ��� ���1AY&SY־��/�Y�pP��3'� a|� J�MITP�� �)Q* @�
�UJH�(U44
< }H� �� @��I��� 	HR��* $�D*P�*�!@ �B�U P	H   ��8   �@�a4	i�>���C��l ����h2w8�E��N �݃�þPT@���ې���|�LO��#��<̮�yz �&O{ܫ�˙�X{ۼc#ި!T�|  � �(q 
<}*�}��<�zg6����W��
O����M.,�aϰ��̪�A�If}�=/3Oz:���zy��U� 
8�Y��Ξ}������w��W��T�Rf>�r;嫓S���
��>|     � n0 �JR��E)�#J� �g�� =
14R��i@SӠh��Ԕ :0i�9((��T �@��P�D��E(���ҫi@3e(FA�s�)@� � {�zj ���   P ( �� �򃦎w;�Yy3�'�� �Kݑ�rڗ{�͠` -Ig��질p����b��2� ﷃ�/�)��Y��n�X }���X�T�o�\YE�J8�U��  
  �J b >�!����˳8��ؓ Ct��B�}�'���� )��' �=�Pzyr�l�� (�A��2;����h� ��{w�<���!��8À  =&�6�R�  $���   <z�TTm�`�`=��#ҊPa2 S�&��)J� h ����AH��z��w��?�`�����L�}�}�Ͼϵ�"�*����UҢ"*��*��Ȩ
��E@Ub�����UEN�_�C�a���V�3P��O�\�����oFȖ%	#pѴ�42��������L4Մ(����\�q��0��# ��_��*d�V�J�*S�}),ÕO6y8��1�<\{�+C0;Tc�ӝ��P���^�k���!��L�4эJ	�HR%XB[���IHEaHËZB����S�0C�z',��7���QR����n�rX� "�&�S1�1�MsI.�*c���~�������`�r��0`��Hb��"Qp���%!T�H�1�B#������;]�������]�\�¤J"Q��H��v4Ⱦ��� �6逕�~|lX�=e�#�iW����}�gz*^��*�X'/7|��\�m��3�ˣ�]XP���w�J!h��3Z�I��DAF�"-c�� �:�I�`Ō8Z(UdЍ�R
2.(�ľ/|��!H����@k;B�D�Q������np� ��IL�1�#@�P�UQ:��`�X
QHXI4|m��K��A p}+`�"�X\�\��0B0�,2 ��\D`�
"%+X�2/9����X5k�*J:�°��XS|g7.5Ʀ�j�^����9p�,�ت�(J�����5�0�/��w����9��]2�<j�gO�;�t�A(���}��֔YBU^g'*HX�ߎe�W7�2�#�"QfM(�9��R���9+�Y*��xw���wM<44��<c��ˮ��6/6�ܹVK}��O{�x5U�9w���Z��5�����s>�>펧ҕ�pU�\(�_eq��|2��Jƃ�W���h�E������T�0bk/���stss�Ýkz��9Ga���H27'k�>]��a�w2�R�����x�E�N�I8�b��$�"� @�"��!� ,2�3=~ֽϽ��{�|%g\6�ss'D0(���넠TC4:�@\Ѱ�a�XZ�D(D#�0i �WNn����eY�5)�C�DĔ��0�f�!HR�.�%F�9`Q��X_������� A	�PP0Q�V���Ede�����G�MHj-H�ԍ�L]	x
��\,�� �%�PD�K�|Ncvd�\�)D���w�^Д4���hn`h�V�wЕ���7:OMes�NЕ(l��L;�,��a��dy��*0�0T����Dc����2���Z�*8%%�]�	��4ҋ2��,���j9z�Y�M2&�cVD��m�����eĩhU�W�iq
�FX���B{��C��p�M���&8����p40(@* P�Q[0�Y@�p+�*�(S
�X4��@hS�X2��� �79�7fJDQ��J���2 �%DH���p�p�� "H�B�h����,�2������n:V藪�E`�*���ա��j0�,�h�6P��p��a�8���\�%��H��hP 0-@���"$U�Q�l�E���+�T�d(�� �4$F�������|t6�2E�F���20Ao�@Ij��k �(bs� +tӒ��R�M+�
E��� �
�
��
�(�ސJ.sh�,��6	E��,��U�y�1�f�q'D
��l5T�߻�0Fl��A
���᧣(�D�f)5*��BP*�*"�׈����'o7�������M���`Qؒ$��B�eIi06��UpB�
6��LJ�`�Ns�����P	QSd�)A�DҎU��/��4:`
��#��G	�I��$�&��B_5��x��4A�cM4�rD�u��C�ܦ��)sOx;O7��ZnU0�	r��FT�	

`P�D�������0���\(����/č0(�(�Ĥ�q���)��`��5
F����E�(�#W\��<DѠc�E��0������5�A������:�f�"P�(R5sP���&�HxV4��B�׉����^�.�l�1l/��q�Ԡ�*bS��l$C�A�I����
j�7�8��4e�q��ɫ5bT�df�ĔX8Y
��R��L�D�����n凑�x3���F�5~l� �F2��#@�KV�`�P*��Uv�}
�����O(ߧ�>�DR/�$Z֥���7T��2[u]���>$��0)��@�� 0l����������64<aL)���Lk��B�º @�.ʒ<NJc��F�  ,�@���󴩑0�<���ن����5a�9%F�l�F�eJ,j�k2o>��l�Й]Ve別%6����
`,�M��o�s��cw���B|X#*̍X�V0L*4V��*��#
�pJ� ��g��˿z���%K2�U��J��qt:%s#E�+��Uxlf�CN��f�j���3�l����J�
�D����׈����9���=��WY=�v��V��Ԭ��aMl✡c#K"�yNst�̀��<�s�� �PT��c�/)��k�����}�c4eQ�ei��2J�ͺ�w3�[���Ԩ1��bQ�m)/�oN�ٜ/<	W �ʰs����´Ѹ5�J9���*\aA��
��b�0U�H)S����5"K����g�,`�U�b$eW�ꨫ�{����1�zq,��PD�S(� �JR$`�$�XTCF��4X���RT����h��,�$�X�@�`X]��y�S��s��n����a�z0(F/�����X�c4o�}�����&�
%��	��V#@�B��F��0��n��03�f�|8�S���K�֙K�DG|Ձ���#v����zT(W�R1eK�V���^2,��j����M��9W��z�k���`o�hO�(ȕ.	Q�d��	W��s�ϙ�=��LcLa`T�L)K���bi�^s2�"����.@�>�\b:�U0a�4���E��vdH�B���"�Pȍ\B�A�BYp.%�)p�;@�0�00X�1��B!\b�P�>
}�c<��LЁF4�A�!L aE�q��i����ĠJ���XF� c0�0pЇ���ݫ����Dc(��AhY��jcRl��p�˷�
���V{��w��J(�$R�ޡS���y��#��AT,���e�����5%���H��tj��D�^�Ž=�n����l`՘�� �6�7�u�ry2DZ�4E��7x��a����L�D��/�̅���妽]�cc*N���<J:��9va�A�8��r,�ٝ���e�i��F;8�@�ʂ�@J͉p�9�!L��lhċ]0���Ky5��@2�g�D�J���B�
ĉ
K���f�K��0�Hq�t&���ߍ`���3	�Jӊ$����")%s��_7�	F��1�a��"M�V$'���^�/&A��t�5�J���u�J��Q�D���^�y�^m�*���gg��V��ʣ��q�{(�8rjUɌ����A�]��Qӕu���FPXMB�(Y�7�,����`�KOl��K�J��h�K�N�o�4�H6e�d��k~{Vf������Z>��r��7�@��`܃^�g����1$�0L������7����WG)ӭ;'/�����jd�6(ʼ
�v�t���(���M�ߺ��nB��TJo�z���b&�kV�.�Uc�5���_�!h&g�(?o� �ґ)ƣ
T��g��<<�P	Fw*�����7�D�1*0�J�܋H�'�H�A����(!DC�gyg�C@�����Y
0�ɳ�δţ������XR%���H�F��h�m��V%��>4k��R�+"P��(�0{����<ZU�@e\����6��^���%��<4]��L���ff   l   �    ��   [@    �C�         �   �     �m  �       � -�m �� ��9qYj ��j� t&��i$�[l0����"zH4�5Ycm��im�N\����ݾ��|�1���(聫hȲ�<�ɫ�H���f�"ީČA�e_[�ۓ�k�@�ת�f��W�e2�[j��B���]�ڥn2J�T��%��j�Ͱ�`m�B� I!{wH,�����ūY�빤��ԲrW�CZ릠Nb^��Aԁ�\��V������m��m�3֧j�y:�<*[E�i�4<����+�n���.�A��)7�1S�ܰ3MO
���,ժ��ۗ]mքI���2�/9����]#]Rr6�m^W��:�25ŷ=%F��3��N�4&��=����=Xk�]a��`H=urv�BbH���j�� �.��[���%�v.����H$H[�l$6� :�9�]ڭ�]���6�V\:].�t�n���6q"M����m�s�� Hh��lp     ` �K:@6mےe�m�j��-��붼 ٲ�IÀ$e�'[,�t��K�ꀪ��U���Vו�� kKX �  $�p��  �^�IoUTݪ�THH��=�4�V�O���~� l�I�m�1�l���@8����媪 В�����p��඀�O@m��ڢ�U^8636�W�w,�n�L,1�� �H�i�#I�v�	z���  �      �Z[��#��]�� �a��a�o2�m^�N[h[\�m�P  ��m�����$-��ס�6ئ�m]�
 8�'�G(MU�+��b�A>ފƻt�Z���.���;
f&��@��Z�vVf�Dk9j�a��,vjrbe��r�5U!ל���o�R�D�-��*�ĳ��N\^9�U�mUՌS�6�ϲ�h�ұ��� �U���W���S#��\�!�[�ms�UR�j�^��n� <��[u�&4�i"�;i+vIm�����k�ϟ�
�[f%òlJ�7U*���E
�WWv
�8-S\�j�  tE�vvk����t  M����$��k�uPm�b ^�e����(/E��p/(�  1�]���ݱ�n�VӏgJ��ɝTY;jzی����q�2.����b��ڂN�uv۔��;5̍�!�'Y54����ң=��K��ޢB�1 N�S����jꀙGm���ږ�������EUU\p�8�6^P�d��5l [Amn���v�ֶ������c{A�n�@l8uU�7z�� &� m�5�ݶ$5T�X��޺$���Z����ָ�� X)���Of��R��E+m�1�9 �Ћek{ﾟ^��Ii�o6�[l[D����-�-���ݺN˸a5[��k��v���n�53��J�yی�*1l��-��� �u�g[	+��ռ]	r:�2?�𸢛d����ƿu��kX l�it�z`p��f�IKR�[m�! m����7�U��*�m� -�I�`�k�Kv�d��^yAʛmS�� ��m��ӥV�<$[y'�[m-��e��m���Md�qͶ�i0}im�l�p�l�#�ݻMg��Gӡm[Au�p��h�ٶ��M�4�hl�:�%�N	6ط&�� X/Av���j��lrtv�[m�n�	&�\�⳷R��hJ�m�Z�͖��6�`�P��U e�����ڝ5UTf�����Ш<z-���l ��
�UUu�\��6�@���h H5�V%Ik�tn�C����q/z�l:�)�I���kn� �K���A�m��ΖID���v��&� �koa�m ���X��w4%6�۰p� m�� � j��m�f��#��E׮h�kv _C$N��չ�ېmm�}O�z��r�Q�-�UT�zG�6�m�P��ۯ����m� �]�ݶh����  �p;m��� �f�ڶf� ݳWl9z�n�/Nڶ�E	6�m�m6���JU�<��]V�U���m�K�հm�5��
��Sl�m��E ��I2���eZP�TՇbPUӣf�OjIz��[@ �ۛl�4���:D�m�h��I�Ŷ۶!a�Yd��� �k��$�@���mT�����jv��
 4���v�2���U���d���m  
��6$'(�m +s�8Ή$H�[@  �ll���&㶭�F "q4�^���rI�٭N�Q�P�*��f���ctҚ��ͫs^ma�^PA��@�]��mm���{e��Ӊ/n���i�{i7���\�T�/m�*vڒ�U����eۚ�õ�E��]����]gt4R��UT�%eh6�� �t۹�Um\qmk�ݺ^R[v�` ɭd�C���+�Y�,ɑ� �Bu�ճu��7-H�u�\��m��`�֭���ƶ�χ�߄KZ� �"I6��n��n�g   �Ƌ��[G�mt�"�6�*��f�Hu�6�@�%�m���m�8��npi1mp[M�a"�   :ީ+g$ؐ8����p������]UUm��Kv�l�b��^eZ�T�:� ۷l�`&׌�-^�K.7&p d(P\Õ��@���m��p[d��6�u暭��Ɛa:n���6���Y3��6� H��h��e^vYI����9��4�=�S���5�4���D����m��1�I��[&��A���ٻlH��6�.�'@�x��W���k��[p�e*�*�
��ʣ���R�V���j��Y^�Gn���@�
�U$̣�v��������-��(UJ�*핐%j�Ns��:r�䍶��n�`�G ��m[Ԑ-�ݖ�:�l�M�R��̀ )I(l �RI���]���]�Aa�6ۍkm[ �6�"��(K$-�6͚E�!tۛn����Z���L��d�]�v �ծP�I��ݶM�kJd6�@�al�l���� � �na5Q)wK��6RڗaY�5���u�i��:�/^�lXe�l�(l�[BAcC�����~�����%��h	$Ӕ Hm���l��amm��  U�l6��t��mY� u� n�$pn�� �il lrSbD�ڷ���[Զ�m�oT�R�F�(�eZ�'��%� H�P�y�78�WJ�m�ආ��v��Im6ٶ�ƩoF�[�ŋ��e����` �f�[� �jY�}o�ݶ�ԣ�h)[m2�+-̧4KcU,4Ԭ�J��4�UK����x�ہ��&�Z�h�  p	l/Z ڶ5�%��� Ұl/Qi  ��l6ٶ�r��UzV�%:�j������I� m&-/6l6�m� ��7f�oϕ����m�`h '  �(hp�kX�8[@m�mY��#m��  ����	KhM���0"�&m�-�,��pR�Aڕ]c������` ql�@4����#� H�ؒ��m͚�fؐh3f�   6�l	 ll�Iefj�*U�U%�	@j��F�%�L�-*� �HOR��o�ěm�kn� ]+��\$�KF�[[M�l6�pm[&���ċz��`m�sm�[R$�����RK{^�j�,���6��(Ԭ�z�h8B�5� H6Ͱ�i�$l �7lԶD�lP����+�5UT;�VYZ��R@�9Uj�^��  ���5��g$8T���$H��u{5�gc�ݭ65�� Kii�>Ym|5�m��ق�
�pJ��J�D��a��g.ݛm��Ͷ6�� ˩nٖ����R�O+m*��m m�Amp�bƷd0   	   5�m/ZV�UR���N���9�m�j�l�{]6L9 ꂪ��OO(�R�WV�a6�� %�m���' ��e� l8 �ہ)m��rF�6[ ��ٍ�� �m�H �}o�hIʝ66��   ��@  �6� @$9 �m� �EK�*�U*�+T��P 6�v�� [D��޺L�l �p�v�6�Qtۀ7m��   8��GV�m�   p� �C��m�[A��` l�6��	 �D��nm��K9@��`�	��
U�JԬ���p[]]T��8$  �il�kX�6(i6j��m� j����f�l�K(�$��d�&n -���R��i�V����F[�[�[vۀp��$���AO'մ�ʪ�e�8+eZ�ڕ� ��f�  6͛b� im$��$6�5��nu� [@m�-�� 8� ���� ��]�m-��l�� kZֳ3_�DER(b���?�x��1؅���]
DdQ"����W@A��x� �<SГ�J��_v�*	A��NP8��=Ђ"T�EY�hР4��L|
Q��8 �G�� �@������E8����(!h	R���(!(�6hX19��)���"�TBQ*���>�'�qP�}�1'��h	��M+�!�D/��h|���A�}�=�G�@Q=(��&�8"|1j8���J�Q��|�@��z�!�h��T��^(���S���B���D�D~�'�� ͫh�H��C�1����>��E�B*�b���lE1<qb�
�������}ACԊ����E���t ��⊄�hCi��C *�|�Q�}u��0�0H���AA<�C��L^8��!�8zD0�@"�� &Q��
;>N>�_�0��p� � ���� � �
�@�0P���Q	z"�
|U>H�x��`���� ���dQR(�$X0I0�$` E��I0�� P�J �Z�G�F��@6x���O
�$a�"�!�0E��pWI�z$!���m@8���$>(�P�a�"�b �DW����șȑH�1dIbF0"E!=�P�E@g| k�1p<P>	�R�>G�`��\^)� q4 |�S� ��
+�g��U��G�AHR�-DbqB�	Q�,�����ޗ����?Qi��Il�ۃm�� 	6�� I��Ev�Fֹ'�d"{
�nM5���_]p�q��xEc��6�5,�L��8�<��sl���Wm�R��uM(�
�׳ەx��+*x�ָ�oF� �;��U�v�1�+��t��[u�+��P�@C��	�)d8A�f�Ґ�%��C��u����M��*��	�E��<�0��P`�67JY�c�]��of�nW���*�ܜ.�{S
J��Vs��u^�����M���eu��Q�u�����`x�z���'Z��^��]��Y�iR�vZ��uqƠuԬ�d�Lv�6j}ֵq�r�c�"t�j�U�#%�cu�X��L����'mKdDv���'gn��5K�0�,�C[V�n���Zc��g m�p鎮	�<ɪ�Է6���K�8	�bM϶�Y�������sRa6���]��uA��2�P9x���TZ��h��E�MIԲ�ɢ�ö�$�S�s�u�����/i�:kO:ȨH��L�;F6�a{W2��ذJ c:�p'���-����]��`��Y^��:e�cvв��m��^z� m���z	�����<ݛ��y�;vv3�]VּCv6���K6���oP��\�� ��WY��<Ps���ځtRb�+���g��n�`W��q\�P��f�l�ѶHѶ�G��*�ٻnI�UK̯V2ϧ�K���7m�Uԫ���f�]�Z�[�u�)@��u��B;s���+Ÿ���.�F����V���G5���E�ۍ��n 8���k�f.#n	4U �fG�X�=�jc 2�]4V&�e	�m��4�=.��d�k!�f�E�����Wq UUU��UW�Z���.8���I��.Y7n��Tnm�(l�ZmԬ�v]:�m�Q��Ӕ���#m��5��3����V�V��������n�l�sr[:8�ҩr�Am+v��SXd�54[�&��*���?"'��� h�S��P�T��ڡ� '���v�� |%@<> ~Gk�m"
:Q�/����Tt��ݸ���OAہ��P��5�r�ئ�Fzt<��-�:�Zq,����&f�����;a�t�E�ӎB�x�`vm��c�aD(e�����ې�z����3n��&Z�ݝqYy!�m��$=,	۝,2�9��8l֐�<a�.�"қ�"�&Ν8��;Gn�F�	�mԁ'���/K�U��d-��J8�s�ՖkU1ة�j;��\�,��6ܹܣ�܇/�;��ۃ&^������!�H�+�t�lp�9�� ��_��\@o���P!j��]�n�� 佋=U��$�� &�<v8`�)�Q��v��Кm`ݏ 7�;0Kذ�J���J�]��V�x���	��r^ŀv<��թc��l��N���, ���~�N���s[��4�զ�4]ȱek �0W�����ڎ-�0�u�A.$͵a�N�۫AT�g �y`ݏ 7�;0jV�v&�ӧUwv� }�}�^��b\d# xzH�����p�9/b�5D�\�n�cEڤ���ݏ ��%�X7c�"���+wbm;��Z��	��r^ŀv< ��xZQ���շV�*lM�%�X7c��ǀN���<��˳X7� �����j͵۳��r�l�=(��+S�N�0.ں�Cq۞vՙ��t&�\ ��x���	��r^ŀ�lZWj���$����$���q$�w��I)�9����m\jת�1�64�-�x�K����+o�����|�X$��#ȩ@�U��z�h�<�=��[l���kv�}��;�wmա���s�%۽�x�J^�q$�ݖ�$���s�$J�ڂn�պl>��wx�J^�q$�ݖ�$���s�%۽�x�K����y4]��J�ãZ���[t��6��n���P8rQGS��ô�Q��ӣ)�� 1�������q$�w��IKݗ�$�W���(sD��� �~}ߟ�����T���]�I/\��q$��-�I)zQ���շV����$�n�ĒR�e���݊O[Ē]���Ilt�(��v���I��$�����H[��$��̇8��@���%D�Dڮ"8!��Ms3�ͪ���j�����ݎScn�Ē췉$��!�$�ۑ<I%�ݗ�$��Z��RBU~WM�*�h���ھ$%��t��r�;�i.D[G`�ȸ��f���)�64�v��K}�?�I�Ē]������B���$�����wv�Z�j�s�$v�OIv�e�$-�oIsd�s�%��ڂn�պl>.�$�{��Ē췉{���x�Kn��I%/Vڸ��j���8��}_}j���I%��r�Ē�ܗx�K��/����W?u\�w"�| ??�~�W8�^�o޻�I-�=|�Iv[ĒW)	8	)��6!���~��̼̼�r\�vmH��p��3��+���@+c�.�qI��F�Q$�|WF]��EV٢8����rs֓eb	�8���@��=���M;c�a��n.��G��ktq���ɗc�͜:��7tcs�n��4�\�Yռ.�]�,dګm��Ϝ���A�* �%��;9��2�XL�n��m��Y��quc�DΊ�pf�x��?�������ܧ]�]�<k����y����p�\����٩���=��"�컣��䍮�wߠW��� ����H[��$�����Kc�	F7c��L���$�ov_9���Ф��I%��r�Ē�ܗx�In��c�.��w�$��e�I%͓��$�n�Ē]��|�Iv�Z�)���64�v�%�����s�%�~��$�����H[����q�痢k�G�7~~ ��ĒK���$-�oIsd�s�%꯫������ �:@��s6�*=Lm��5��gq^܇ �3��[(�sƪ�y���o����I-�ϜI!n�x�K�'+��w���_���?]����Weє�����k[�:�%�N��1HE�;b��|���P7�m��+�I(�|�B]ݏ�I(�nˍ7H�ӻ*�ݻx�K�'+�I.��w�$�wc�H[��$���j�U�n�4�n�ė��ﾫ���I$�O>q$��-�I.l��q$�:`�cv;O��M7w�$�wc�H[��$�����K�r]�I.i�+�Z���LBN� V-t�[���0�팝,�� m+�6�qrx����]m��$��e�I%͓��$�n�ĒK���Ē�^�jSmS
li6��I.vNW9ﾯ��m߽w�$����$-�oIn�I�t��5�պ�W�Ͼ�ݶ����r��E64@CK�����U&'2�$�����HڸJ�'v������I%���Ē췉$��r�Ē�ܗx�J_R6���h�T���Ē췉$��r�Ē�ܗx�Iwv>q$��YB-]�I����[Q�8\��F�ׂ�\t!��46m�e�l0p���n�����v�$�6d9Ē�ܗx�Iw�8�Bݖ�$��V���n�4�s�%۹.��]�Kvy�$)=oIs�!�$��L�n�i��	���$��v<�I%�Ē\��s�%�r+� ������s�^{FsO����y_�wZݶ�=��9�m���\ݷ��@�a�QL��v�ʪ�쫯��S1ċm�I.l�s�%��~�$�����I-��$��g���T�P���ٍ��n:t���P�gq̦�Ѭ�t���Y��f�iZ�{Eo���?��� �?͗�$�[��I%�̇8�Bڗ(���[yV���~����w����� ����Iu\��$��ꭅ�t]�j�v�8�Bݖ�$�;2�Iv�K�I �?�o����T�Qv��K7��̇8�]���I.�c�H[��$��
�V�-��M�m��Iv�K�I$�ݏ�I!n�x�K��q$����_W����1��ʔ�r�Z�H�z��"�]��&��Ru�6�cH6�v�B���ɔf�+v�j��à�.�u����lv�Ѓ��wU�$ug�e�oV�#e�aݷg�s��̼�+Wjs[Μ��_�'��K��6�����6�%�U���:J�����j�_6�t��yT���N۴T��v�1жbP�nɖ����j�Gڦ��̶�����f^R��$��rM��l�i��ZN7uw���0��ʸu��6ĳch�g�*g�	uد�
�&��:M��I%��>q$��-�I.vd9Ē�ܗx�Kk_�c�-]�WBE[m�$-�oIsfC�I.��w�$�}�|�Iv�Z�)���i6��I.vd9Ē�ܗx�着���z�ĒR��I.�'�髶��g�M��Iv�K�I%�ݗ�${͎�R�hM[��뻷xV�ԶO>��� ��/ ��_֮�^*�_6�I�*T:�Iͫ�r�T6'��iW�h�er'gDt����v4]��x���lp�8�K�UR��0��m��˻z�8��6��3U�~ϝ�= ���$�@��}[�^��ݗ�ݏ ���
[ut���0-���� ��x;0��RQ��i?��4��]�x���v8`[%�[h���j�,�� ;����<p��^�ݗ�~�x������UX���m�Y�zNn�g��幗���8D���gGK75�]\�s��Sm����ql��uwe�wc�;�JO��VۧVφ�0-�����$j����� �c�z�H$�_��5n������z�������}�F$:����\�8ױ�k�O�p H�յ*&�+���`n���V��o��Ç���V!�I���a��ڐ��:����G������HEa"�X; �bU�Qcq7��i�#�HI6(B�$?mD�P�! �B]�X�6#�	��rc	$X	^�o70K���Ѕw�cAH��F,"�T���Ӣ<�;����Xs��d�� a��J�nd��F �hK��ܓN��CK�Ξ ��e��K��|��Ij�G! � H;
�j�uGJ>��4x�U�Q<�*�(� ���@��!A�0j��9򇠠z%6
<SP/�kT�8��_~漛�l�.��]7E�բ�
�� wv<���x��m���=�v���Av�_]��sc�Ų^ջ/ ;��ר��q����,�M�u3���Q�n�:��/N\+:����i��K�k����N���?���:��xV� ��ɵT�0�6i�;�Z��[�7)�&���v^z�H6O<���Ų^mRI�[lR۷"�6Y$� w3^���xT�x)wU�I�S��Sm�{0-�����4tC�F'\"��A�aU5�!�����O��w�nI�0}ʗ�W
#���s/�um%K&ypRz�m����$�V+����nx��-�{;��v�n����GG��Vԅ�Ar��4�T��7bj�6]ݻ�:�����x68`[%�^�F]7B�2�P���:�e���ql��un��${�.�y6����ۼ���Ų^ջ/ �ݗ�IAS-%wM5O�`[%�[����x68*��7���/2�M'�`��x��[rz�*���_�/�w}�.���ݾ�� C��!gi{�k2̷3&�ja��C8v�.{n�dm��뷢�ql/Y��g��-�Z�\�U&;u8�����ώ7=� �7���m�;q{iA1Z�\;�Ӷq�8mg����@<b�m�ͼ�Z�q=����3ch9S��R�Z;\�,H��rX"vvtF��x778�eM���m���l���s��b\�{u��,s�H��͹���l�H�͌D�k�34�C��k���vcCX��n�Mr�B���&���+����f{Tl0�RY�q�M�t�W=�:��m�}����sc�Ų^ջ/ �.��L*�im�͎�xV��w/�M����KQܑEp�9����>�/��^�ǻ���O �Ş%��t�}wv�<��O^�O_����?�I�y�|ul-H�c���r���{��<�R��w�~盷�>w/���������f�qt�W�6���7-�����i����bۿ��_>U�l16�K����4��{��>w/ԩW�%��^﯀{}+�A�.En5(�$��߳V �B� ҧ�*U�J����{|�wo�~�&�y*��=u�ߡn8ܧ˒�=�_ ���|<�J���u�|�����[v�WBE����Rۓ׀vy��8�K�:�e���V�he:��ۼ�0-����xV��}�UV��p875��`�]�e��|��{F���[	dX�4
�3&���]soh��T�� �ݗ�un��9�� ݫ���ڶ���뻷xV��v^͎���䈷��]7B��7WE���~�������ăE�����6�|<���s�y�nI����e�ݩmӠV�J�ݻ��.�� gwg ��ܾ�}�;����c�"��I w���<��f�����?}�ꪬ�Me٬�ӂ�ݎ��m��4�ݔG�����g���F]�t���vΒ�Zhi�l��@�{��Se��p�}��y�����M���"˒��3/��+�������>�/�J�>]�-�"���r섹|�٦ n�x{�KT�������R��1ܸ��Q�U&�7g ����wﵹ<@<`�xD�
�� �(���� ���/�䬬���M���>}�_ �I=����f� ��N䪾�q�v��-�.;#(Ѕ�3g7iH��������Z��ٔFR�绻�9�r�C��Eh�%���� �ܘ`�����Rz�	�v���@���K�' �ܘsԽI*�v�zp{�� gs'6�%M��(�F9r+q�D��{�|�����z���vn�Ӏw}<pݼ�㉹N�%�6��>�f� 37g �ܘp<���IR�����j�L{��-ȭ�I/��d�^�]�~����_ ���|�]BI}IV��;���{��w��_���&A�n-�^�nH�kg]��e[c��ڤK�ZT+��<�k;h,�닒,����ƥK��1�[v�;n�[M�k4�{;[9���Gn��d3��2��pn�M�v�*��l�g�l�t:;S7�6��l=r��c��6��\�ѱד��,�{�wn�-���Y㋳=��ݍ2Rb`N5X���{mǅ�nFn{Z�i�LuӢk5�x tEv)�K�rK%��y�˫YT�;W��lk�3ӻ#�������E�p����U��Ƞ���˓�{�g��>y�|�����^J��7}��7mz�E�\���Q� ��e���+�﯀�����mRlޫ��YqȤ
��w�j�׀�<<�g��W���:�)jD88H���K�w��N����>y�|I��6���ݽw@��J��m���z���_ �'� 7dxwRI�Uܫ�;�ݤ|��v���͗A���\����٩���{֪�x�@��V����8�{׀un���������~�i����'m������%��V���d=��4KUH�q8Ut$*��j��w����4��f_6�����y0I��,m� I<�lp��UR]^�� �'� �v��M|��N�W$�T����8�wo�|�ܾ�RT��� ����h�n�[>l�8���^��L�_����?}���M�o����*��8zi應*��*���\W�!�4g5��D+�M�������6��V��[�^ suG�w����Wu{޼ᰵ"�Ԋ�rK����窪��I]���8_���?�/���v��ו���IRe�o ���qI/`+�)"O��ZD� �0��l��}���܁�ǳ�g׆��\��jQ$8Iq$U+�n��y�| �޼�����e��e�N���'m���/ ��.ȼ��Ix4�eb��b���kVZf9�mP���)<� m*��n���h1��.Χl�?6۲/<�0)%����~0��K5�n�v9v'q��?}ه%*۳{{��w2i��ד�I��koh�+�W
#����|�ݘp�R�%vw��8sg��W�NK�q�"�wi?���uW���٪�ϝ^��|s���Nj�(
��u���yw$����L5�p�Z��p�u��UIz�b���������w\0	"�*�E�fTg,�I�h�\�q��^'����k��l[,awl:7]��揊�*�-�Y2����ri�3��|�ݘ{�J��;�~�_�]�۹�ԢHp��<��UUU������N���9�*��gr����Iհm`��`&����_U}[W{q��=��,Q�`�7WCe�p�z�$����+��}s�w}<p�gԫԕ$�����/�y�-���Z�;�� �ܘp*IyU$�����~��?����W٪�w8Fv�!�O���y4i�YY
���Hp�}�ӰH�}��58`k[#Uk�B¥HI[D��vB��Ĉ�� �$A@d`"g`����Y�����4�@�t�I�1a2$H�+�� 0;"	H��^z :{�4H��ݍ@��R!r0"�b��֟��x$T`�"D�<C��H�$�յ}6!�%�8)��! ċx��$I �o �	���v�� Ca F\D@E:]F��t:�xH.Y�������CT���MF��c��}P݃*<X�!+���s2�3333�i0    A�� v�a�NSK�.�5�̼ܠV�e�4<u�r�lnf����h	v�.ܻA�zz�Es�i��d;=g��5��k�-�Y�۲��L�,b��P3�Cp���L��9v��ضx�M*g�7�3�<88��F�γ�eX��Q�1oQ����yYEYekzאu�ׯ�a4�T�ún�͕�Ij��l��c-h�|������i Zu�"X8v�3�5oE��=��v�M�0]SX�r��LV�����rSQ�kq��mp락z�8�r�.q���vB��=�%s/>S����/��6�	̖v�/\�[I���N�/^!��m���v�ґ�����&�Y@۝)7Q���G;�n-1Ɉ6��g��d�.]C͏pݢa���ez�v5�\�xsD���hb�B�<y]��� � ґ�M��m�B������3��ܘ��m�r��(笺c\fZ��d2h��7i]�͕��v�8\��I�nH��v�r�捬���cv �18��s�chz]�ݪ��MW|�)��2��zvv���#��*dP���N�4�r�,�0>��m�q�@�JO�cgfb/@�
ر��>���ɢ�wC�X�BqճC�ۍT�����>z��ջomVc�J�v״P3��k5��c+�h��U��m�*�
�i���ۛ��r��j��+.7]$�t:%[����S�Ѭ��4v��v�J�����j�Ӣr�۱PAd� ��{a{X��^
�-�(�UtUk�lG��Y]n^�v-6���[R��t�Zm�H6M:�lt[tN��.�����U�<���<
Ծ�uUg5�����R�Xh���@:��`������V��vh�J����>~m<;Nf\.��;�ɷ�-�/2�:*0jP�خ�B��<4�wQ�E��v�䃓��f���i�j�<�*�2��݂�98�v���ݴ\�fқt@{;�Nˍ��Y�'�g\ڣ��\>z��v(b����$Q1:� h�>T"f�@�� �+蠾
!����7����p%.Vwi�:�p�	�f�^��'3�[��ʴ���Z�֠kp��1��<r��Ny�a嚎��v�x �xMC�[��>sΪys�n�����ŗ�u���;����n���М��:�-����7�h;��+7`���Б�ا��vÛ��ԅK�T���Wn�'M�w.H���[�J���^�&CB7Zũ52fj�\ֲ4R�#��
?������Ï���vz���c?-͸�=H���N9�2�<F�u�҈Q��~ww{����W
#��7w�\��a��ܹ�*_�}�4��{��w�(�nE�>�f�^IU�w��8w�� ���\ԕRD���T�
����f vE�~�L8y/UUU�}�qpݞ8e���;�X�&�-�r�i$��7�p����UW�IvO[�<��ߕ�n�ƥC�}��\iRJ���? }���lp�;������V�4��ךr*nD�>|�Ny��py�eU�b����{�j!��E�I�Wn���`7e��ra�UU_�wwx�3h�,�X�7�x�=��7��P,*!��EC2P)�B��U]UU�����͝8s7��}��9��&ϗo,�#�D�����f�8$�X{��Kv?�=o ��K�Z�r��D����T�ww��fM8��˜*��I_w}���~�9.��p��&� ���]���d�V�&V�(���^*�_]1���Zseƹ����n8�^8���	��|<��~���o�,up�Ln���p�z��ٕ�vI���$�������=�{o�〝�ۅ����9�2��_$o���?��o�U�Wg��:��r+q�C�p��Ū��ϝzQ��&��7�����W��~Ӏ~��2�-��7wʕ*^J���� ;�����.V�����δ)�:,n����l�wU�'�W;���6G� �u� %w�)X��i]�'l�nZ�&^��g-v6�72�x'U��vWM��f/RMrr�HKj'-X��s�w7��vk��뇫︀�=o �u��Ŵ\���Q.��gfڪl��4�s6� ��s��T�g�^�H���(V��� �췇�������7���;�� ��;$V�Hp<��U$��w�8w}��>��8J���$$�ER	H!��F
 |�?"U\�ߺpz��k����ۅ��\�����K�U$�����wvx���\���ｿ�x���zzgQ;�."6��R�^�k��F\5*�9j`�e�FVD���V;T�z�[v't�u�7���9���Q�������{+ �~�yj�i�`����ه<��%I]�n�N��qp�\3�U_$JZ"_�tX݀�[m��/<��+U}T�}��?k��!"prՉ�rp5US�3.�G� ����-�y�]z��m�(�K����ÀyR��$�����w��[�s�~ٹ"#�"�F���������ݏ��S!��SXRu�^g�I��H-�'Z���@���?+t�l�����^�9��;�i۰�]�ܻv�����G�ֻ&�L�qu�����d�s��]���on�Sî��6���#��!�,+��nk�v ���-�Mw�^��;[�����]!�FĩBuA�ëh�\����g-�r�N�۩�s�v�cQ��&.vڧ��N�r������3�u�i���˺��,��*�������E�x�X���#���V��� ���ys�禇i�L.��l�����o ��qz�}a���o�~���H�l���x7fV;r,����#��=u��I2�v����X�Ȱ��}IvG� '�����}w���-J���$�&��fM8�Ǐ�T�'�X���cV�L:���ه �UU�J��~���qp��X!�ZD�e*HjӤ��+��T��A��cL���[3k�a�=�6Dhl���q��o�,�����J�l�����ٕ�M��i,�÷�N�/U셖D��Վ�fj����n�XI�O����5��M8�Ǔ��IU/Uٻk�� K��W
%�\�~���ه��=��vOe`���hv�t��wj�ٜӀ��8��8��^��g=��7�=�)�p�Z	!��e����I�W �߼�n�`hTPs��[�pTE�u]�p��g��8��8qvd0�7��K�Ǿ-m�pL�� ���"�^��}_q�{��xcb��n��R�"��2��J���T���� ���{�\�I*l�]z��1��0Lۼ�?�&kr��X���A" @�����D4'��w͛�{�}۰:ϛ;�n"��;�C��UUT�n���f�p��ʗ���_wx����~�[�'��.pٙ��5R�O{�?�ɧ ;��8�'��^�x�6�F{p��{*�lN!��������ȶ�ۚ1��cn�H�zs���ѝ�����3��8�̹�T���{���>��jFKrE�n\�>�Ú�$�f�����. gٓ���^J��z��
D;�&��8���p�����#�'u� �.���Rt�v�]�x��s. owg ϻ0�Z�J�R�������y��$��vW3�.kF]*5n�vG�ou� 6Io �ٕ�<���a�f��e�PW�m.�7k��l���G��ϲڝ���쩹�󽋮��Y��0LM�������[�96e`� �ԃcuj��+�ـ�˜�I6}��\ ���߻0�*I/$���/KW襻"p���K���e`�UU%6?=�[�;�R��	rZ��A..�I7�ݜ;�N l��ɳ+ �.O�C�ۦT��8~�Àj�I����ۛ���2|�^����q��Jd��������cl���9�[j�(7b9�ٱ��\��L7���6�B֮{<��)��\���D99�K��љLV�u��AѴ��r��{b��;B7�9�IRT9�^z4[a�9۶���4�\3R�ˑK>ؠ������4e�G+��! ��X�{u"��oh b#�x��;�fL�\�d:{m�*�Y���M_}��������?6߇~s;F��ا�����=�2d�z8��\��NKIj�/$��b-�{���|��8
D;�&��<�͹�?gs���rm*_�gri�:��$@��B.ݼ�fV{�H=�� �� ٹs��*lצ4˽v�En8
;���� ����"zz��Oe`�P�(�n��+o�}�3� OO[�������*W~�����_��jEcN�Hp�ܹ�6�-�o��{��	�p�?}����@�H�:bNׅ���_Nz''O6����N��.D[Gͬ=�n�7U[��!dN��s�;�� 3������J��76� �^����/�xj���ٰB�� �����*p �Rc�N!2l>�W*�%�T�~��ߧ� o��p����Ҥ�6wKݩvII�$�ܚp�ד��R��T�U�}����}8�R�)���t�i� 6j� �ٕ��rp6��RO;�Ӏu��[vH����]�8��qpIU*Os6~6?�Tx���U����bN��v���9����eQz�n�N�l7��[���y*I�q�]��܉��(�/����w��8����IR򤪾���\�k�
�~M7i�覓o �� l��;�\ ��'<�z�I]���_����;�!���N�;�\%Uu,A�0Rɐ^dȱPDb�lDZR��7`��� �|l��>�����) ��D~�e�|Ϥ��Bh7U;.}�` ��d"B:0Y`����0'bN�y�Dc_8�U�Pa\�3@�ʉ��ã��E�����D�Ǡ��A�`��a������I�S���l�B�詁�|>��)��ꠚj#��⯏��j7�hP4���~T�E�}D}A �@����[�¤N.��EN)�dL]
���C�������x���O�2]�V:Lk�+i�}��K���`���7��5G�}�� F�ܖ��PK�����UU6g� OE�rl��?}]��]���]-s[�I�W6v����Pp ����9��9������~��z9��*�9&�?2O՛<p�ד�~�����I/�n�p�R��)�V]6�P�f l�ɳ�������m$���n�۲D(ܶ2���>��. g{�����UUJ�sg� o��pxu�]㻹q�Q�\IR��3g ��Ӏ����$n1���5u�������j�F�-
7$�����*O76��>ݚp>�N�J��p)�[���r��Շ�+:q0ʜpvtvVxY@<�T%�K��w����l��ֺXv���~`����2a���6�UR��;�N�}<��c�ƾB�������� ٲ�{着�"K��4�w%�����l����USfl�����;W'ͻV;t��m�*KʩU�o� �o�p�ه 3���8�)�e�n�l��-��RK���> �o� �ݘp]V�*\�GB��@(b�^�}���k|ď58.�s�ta�6�^ү��v
�S��S�-�:�U�Gmi&"�E����N����kqY( 2��Mv�Vێ����2u�خش�-�b��&.#�s��{����y̘S���ã�*�D�\&�(��6x��\d�mϜ��+Z�\��Jv�b���q)m�b#����!7m[]�ȝ����LUɫ�uY��k0�ɚ�~��pDr�2\�����9�I�f@���۱ׂ�\lOkp�Ӯ-��C�^����^�=�uv�cI�v����?;���p��-�i��q'n�v�_��0wc�|�6?==o ���RF��Ԯ��li�!F�;�N w;�8Uz�]��<`��� ��Q�N����J�l��-�������M�� ����\�dM\LN�\�����=���	����[�&��X���:�.��k�#�}����8�7J��hs��=�v-9qf�aڒ� ����W
p��ݜ{��K����;��`ڹ�MY��-�Vff���>wL����#2P��@�㞂'U{'�����;�� N��)JO�e�n�l��[�95�W��G��x��`U2��d�2��Ū��� �u����%�Kx�"�_�v�m��� 'dx�\0d��I2�����7ݸ�r�u��d�K�90�<�Yۃp��"T-"[㌋�Ҝ�λ��* 4�x�`�-��ez����� ���Zt!�)R��0d��I2�vG�n�{�=���5"bwr� �wx��fN�U+��
0@���	��4��RY䒹{�� =��8{xd2�;�Vρ۬ �����$���T��w.�W�+$�II�$��fUU'��s�n� 3���?f�~�m������n���se�k�l\�ۂ�x�z<4#�$n�+�r0/P����sj�Hp��s�~��. gٓ�U^T�}a��� Ƽ�yڑ�d�2��?I2���URA���$~0d����H���t����պ�	���m$�6f���n� �n�;W�����F�T�S��i��ۜ�fqq~�N|HI��Bf�۹�������H�iܒ �f\���_n�����x�`k� �J�
P]�۞۔�(y�P9�V��N�fܾ�&�#�$�A"KQ^Ҫ�u�Xr\�"jD�����}��X;#�7u��}U���o ��y���j+����fNjU�+�wg� o���fqsԗ���د�ۖ�0���o ����Kx$�X;#�:�K����-��ZM�ߪ������{�\ ϳ'ʕz�w}85������N�NЋn��$� ��⯽�U}��^j�$@�vI@O1 T�P
4� ?�gx~�K�
�Y���f#�uC�l���I���j�;�-\�F�.NO8K���{v�i�l7��<��:�����>�v#U�O����u��I�ct���I��n8�f�aΑ��n���n��zs�����[_5h)��)8�s��e�Ixsh;� ���q�Wi��H�����;w�r��΍���F�IT�=-)�v���w~�{�볷��~S�H���җ4�J���p��xsїKV�M�b��Kۮ{�o��<,��g�=�� 7v< ٲ��$�UJS�HG	�rN w����U�o��8_���}ܜڦ��ݸˉ�K�i�x==o �^ N�x��xb�v̻�dMILw%��$��ݾ osg ��r�IU*^T�]��8�����j�[>-7x;���e�͖�)%��tpI*�b�=v���W6��ۊ���α��Gkr�
ٝ�XG�+ĵ=UJ����,$��ܒ|��_ ;�˜����yUW��}8?/_����Ih�%��ܹ�UK�",�@�$���>������|�e窾H�^^=v7@�4��n���z�wc��}IO< ����E��E�;n�ۺ��ۼ�{g� I<�f�x��U(R��i��M&� n�x���OO[�^�� 'v< �
���!ݧG�4X'WV]��6��	��ۧ��6�v:{V�aQ�Ӗ��>F�>3��n�T�m� OO[�8���� n�x��Z%�U��7��o �^ N�x���͖�ԑ%��(`�F��QnK��6p��N�T�X� @Bt�!@a# ���WV�wZ�krOo{�nI���Uۖ�i7$��Kʮ�wӀ����)%��ǀuJ�M��[$�m�8��\�T��ݿ����ݏ � �Dҫ��Eۥnĝ�n�׍��xջvE�����L�rJ=�n��{����t�E[���"���^�� 'v< ���f�xZj�\��]���w/��rsʼ�+���N o��8癗�j�B�(�i�7E4�x���s�s�������{��f�p�g^I�l���.I8�$�nm�����$��~��:8�U��TB ����O���'�w9���ʺj�XD�Jc�.p�3/�y/UUU�7��{ߞ l�o ;�EĬ_$U�cE�r�a�#�bm�T�1�p��ձ�E���Њ�hx���+mS�gŦ� 'v<V� w:�m*U���wo�n+ݫ.XII�$�}�_=I*��7��p�{�����*I��Sյ ]��KE�/��l��f_URM����c���:�(Kcue�i;C��x���owo����u��|R���6��F:E�Nۥv�R�w��<V��U�}�ת��T-PeJ���sd8+����?F N�ӄ��
�p=Α�׮�,Z� �`v�&����R"k�G���6����B�υ���X�B�	Kv�H	#BX��M� ���(y��@�!�0@A �K�2�D:|`_�� hOP�^!E=�	����d�"_���ϵH���;��
Nh}�
��#�DW�C�	�u��%ʯ_>��s3m�D���  � ��@ �i6rU;�*s��j��<˛]&�bٓ���L+lň�]JH�X7g���vA;#��	��=%v:���70aa�	s�,n(�����N�z:���h�;�e7=&F"i^k9�O&2�����v���J� �钚:�������;ʼ۰=̛f����Yk��vymSP��H^Bm�T܅����۟P��9n����ݩV�R\�=vݎܱvV�	wR]Y"������M��<��q�>���K�;cPv�/(Wn��.��^%���t������6�y��)[ �k#v��=aݎ5���R��e�5���
;ga����njJX����	����t���J�� ����7]��-�Y��윳���9ȸ���e@�HX�.";k��d'o.Ig؟EÀ��gyj5.�V4$p���6�T�	d�m�W�e�Ѻ#)&vX��Ǉm�"�*93TQ6�-iݻj퍩�`��=����qV��&�Q�υ5gt������
Y\���8�i���7%*�s�L�y�tSf�m��xg��e�.�,�14��t�;gjmH��a䴡5�K�%n�������t�)�r�i���m�m�tG�uuu�4���<88�����۶���F8-���i��UM�v��=����ۡ�b�fᠥ��J1M�����*��v�AĎ$+G��(�e�
'n�����L��G�P"r�N5"���5��r۸!�V�M�ga�P�t���Uk�0�J�R��pu��V���#m�k���`2t�(v�j8)Qq����]�bq$� ��E4oV�������e1l@�M%��U�ۨ8�AXb^z�c���iܾ̭�R�y�{>-�t^�c�1��j�\��ʑ1U.�.;˴��ge]qekcn��֚�ζ�q�
��������Yʮg�����K�	!�k�n�qmS��}�( ){]�nl���wx5���nSy��$������O�N�:�X$>�|��!y����C�(>��T>\Sux`��c��)��t6xc8sA��ڛ���WDf�嵛6�a����ƜUu:���F��m��Vױ��ВK��'$`�ڸ.ήxw-'cup)�Փ6�۠:�ͭl��ڝ�]c��M����v]��D���vi��E���7b'�UeC����b�)��M\"�fㇰ��pU�a3t]�Y���㣙Nu��KiJN;[�C��n��������~���`��p7j#Y�����vS/i͎�l�E�ጻ+'Eq��.�<|)�Ӷ��N�������2�癗�U%������_����biے_L��y��w6��bX�'���6��bX�%�߻��"X�%��}�siȟ�*J�VRe/j��՞#%4;%�"X�%��~��6��bX�%�߻��"X�%�~���iȖ%�by��w6��&Re&R̚l�wq��*ےr�D�,FĿ{�u��Kı/�}�m9ı,O3���ӑ,K�/��g)~)2�)2�b��r]�.(�wrm9ı,O�ﻛND�,K������Kı/��u��Kı/������I��K��#�\�	vFG�v�5iN��;n;g�TX�-r�99(���x$NF�_�n�Zl�[��s,n�/a�Ss���ӑ,Kľw��ӑ,KĿ{��a��DȖ%�{���ӑ,K�Yk�O\$V\Q�l��/���Iı/��u��1[�!�!Û@6�șĻ�{��"X�%�~���iȖ%�b{��w6���*dK�t��/×"wm�.��/�&Re&R{����"X�%�~���iȖ*X�'��gsiȖ%�b_;��iȖ%�byk�3I.]�Xܓ���I��I@ș������bX�'����6��bX�'��{v��bXX����m9�q���_��~�)���������ı>�{;�ND�,KC�뽻ND�,K�߻��"X�%�}���iȖ%�bw������ˆ��ٔղ���z2�Cʹ���s�i.L�������c��ոLu0�i��5�ND�,K�u�ݧ"X�%�~���ӑ,Kľ��u���Q"dK��}�~ͧ"X�)�����DC���|����L�Ŀw��i�~�DȖ%����ӑ,K��}�~ͧ"X�%���n��T�S)2�)f)�W%ݒB���6��bX�%�߻��"X�%�}�ou��K�b��&�B���	G�tp�M����nӑ,KĽ���iȖ%�b{�KӮ�&d.Z�\�����L�J������=��m9ı,O~���iȖ%�b_���iȖ%���>�����Kı?b��넊ˊ7-����/�&Re&R�;��ӑ,Kſw��ӑ,KĿ}�u��Kı/�v�[ND�,K����>_�|H��zv�j�3GX:B݅Q�q��-��]���ks�{G�Uʄ���m9ı,K����r%�bX���bX�%����ӑ,K��;��ӑ,KħI�K;2�S552ɫ�ֶ��bX�%�ﻭ�"ؖ%�}�ou��Kı<Ͼ�m9ıL��wg)~)2�)2�_G�r[��ɨR�ֵ��"X�%�}�ou��Kı<Ͼ�m9ı,K����r%�bX�Ͼ�bX�'�=����R��˙u��"X�~T��=�{�6��bX�%����m9ı,K��w[ND�,���X��WQ������2�z��tT�-�3�����L��_dY�Q6B5�5��r%�bX���u��Kı/�}�m9ı,K�{{��"X�%��}�siȖ%�b~^���Y���V,
O\��1^��p������tvs[U�!\�l������cmI����w�{��X�%�����"X�%�������Kı<Ͼ�m9ı,K����r%�JL���j@�����')~)2���}���r�BDȖ'���ͧ"X�%�~��[ND�,K������I��I��ֽ6Ԅ��7-�n�G"X�%��}�siȖ%�b^���ӑ,Bı/�}�m9ı,N�ݝͧ"X�%����[2vۭh��d-ֳiȖ%�b^���ӑ,Kľ}�u��Kı;�vw6��bX�X�^f�)~)2�)2�Z��f��.���kiȖ%�b_>���r%�bX�ϻ;�ND�,K����ӑ,KĽ�{��"X�%��R0������?jU�X����B�b�����`�A�ٶ6nx��I
�wM���;c,m�N�(r"#���Q&��n9��W;��}��Y��YhM��l��s��9��3���1��� >�tw8����Fu���qAy.,6�`:��2�{d�e�z�B�ݼ-�����vK\z-b�p�%9��V&�����یpVP�%�f^�e�f.Y��!�&���7�o��;2�!n=��
]V������ru�,sj6�	uv��{6J�,�kZ�{ı,O>��6��bX�'���ͧ"X�%�{��[�@�&D�,K�{�[ND�,K�[�����n[�m9ı,O3ﻛNC��"dK�������bX�%�����"X�%��{{ͧ"~UH�2)��b���d#R�(�%��)2��~��[ND�,K����ӑ,h�lO{��&��!<���jH$����7-�3
�i7�Nľ}�u��Kı=�oy��Kı/�}�m9�e&R{�����I��K64�vL�ְ�u�m9ı,O{��m9ı,R����ӑ,KĽ�{��"X�%�|���iȖ%�bw�^�$�b���Z�
�N�-��x���bu�)y�Ѫ�xC=[������Y��������b_>���r%�bX���u��Kı/�}�l? �<��,K�߿g6��e&Re/^�Ze�nH��c�r��,KĽ���Ӑ�Wc��x��9ĺ���ӑ,K����w6��bX�%����2%�k��&x�!p���\�����L�Ľ����r%�bX��]��ӑ,Kľ���ӑ,KĽ�{��"X�%)w#ݒ\��[�M2���_�L��(�D���~�m9ı,K��ߵ��Kı/{�u��Kı/�w��r%�bX���ޝ�NKMk)����m9ı,K�{�m9ı,��w[ND�,K��{��"X�%��u��6��JL��[����p���G�8�p�;��xhl#���k�lj�:<J�nէA�=U�ε55M7V��Z�Ȗ%�b_߻�[ND�,K��{��"X�%��u��6!Ȗ%�b_{��iȖ%�b^�_��m�!�n䜥���L��O3vr�!�+��,O�k��fӑ,KĿ~��[ND�,K��w[ND����e&R��~�	�.Z��NR�Re+����~�m9ı,K�{�m9��=��,$H1U�Nd�J�1cDi��G��O�}翽�ӑ,Kľ{�����bX�'�v�v�7F�u1�ֵ�ND�, ,K�{�m9ı,K���m9ı,K���bX�D���~�m9ı,O^���nH��eܜ����L��>����r%�bX*_��u��Kı=�]�iȖ%�b_{��iȖ%���v�~��nizv˪��\�s�)QsўD�^����%�v���n5��jje�5���r%�bX���m9ı,O~�{��r%�bX�����	Ȗ%�b}�����Kı=�W�ֵ���Y�E7����
aL)���߲���@#�2%�~������bX�'s�fӑ,K��>�siȟ�`�aJ�L��cz�K�Ԗ����|���bX�%�����r%�bX�g~�m9ı,O���6��bX�'�k��m9ı,O��L�)��i����Z�ӑ,K[���ͧ"X�%��}��ӑ,K���w�ͧ"X�����>T�4�������~ki�S|a��yUM�8�w�{D�,K���ͧ"X�%��}�����yı,K��ߵ��Kı>����r%�bX���2�3��i_-ڞ�Ӻ }qr��r�q=3�H�VW.�`^���
s�o����q�0���k��m9ı,K�{�m9ı,O��w6<�bX�'��{�ND�,K�v�v�7F�u1��k[ND�,K���[ND�,K���ͧ"X�%��}��ӑ,K��>�u��"~P�VRe/^���nB+v��ܜ���ı,N���ͧ"X�%�~���ӑ,�!YJ�Y�ޗ�_�L��L�����/�&Re&RkQ�����-�˹|��%�bX���m9ı,O~�{��r%�bX�����r%�`~PdM��_)~)2�)2�l�ߥ�"� ��5��ӑ,K���w�ͧ"X�%��9��ߵ��%�bX�����ND�,K��{��"X�%�� } H����PX�"��F*Q�Q �`��Ð���k2LiPkv�c��Q��\�V������n;k3i��<��`��yCrS�.ެ�q�q��B�΋
m��\c������gu�"��(�n6K�p��#����;f�If8z�[7=�X4rN����uc�]��V����{N�7lWlĶ���w������]��q�Ӑ�v�H��Jx�ծǬ	�F]�V��$6<X���o� O�A��R��m�V��1��n`�q]�mrv�s/G���ga�jٌ��4Z�9:��Z���oq��K��kiȖ%�b^���iȖ%�b_��u��Kı>��fӑ,K����Қ����Y�u�m9ı,K�{�m9�șĽ����r%�bX���ߵ�ND�,K���[ND�~�ߥ�U7���Uffl8X�%���[ND�,K���m9ı,K�{�m9ı,K�{�m9�L��]�[z� ]��KV���_�LK����u�ND�,K���[ND�,K���[ND�,K��{��"X�%������MѪ]Ls5�fӑ,Kľ���ӑ,KĽ���ӑ,KĿ}��iȖ%�b}�w�ͧ"X�%����F��fI��K��M\�iK���ZZ5�sv���(4�[Y�X�������[u��.[-�ֶ��bX�%��bX�%���[ND�,K���l?O"dKĿ~��[ND�,K���ɞ-�\!l#rNR�Re&Re'��6��|��S�(�������o�؜�b{�w�ͧ"X�%�{�{��"X�%�{�{��"~P2�D�3g��7"$V�L�rr��)2�(��~�ٴ�Kı/��u��Kı/~�u��Kı/�w��r%�bX�d�ޝ��d�kYL���fӑ,Kľ���ӑ,KĽ���ӑ,KĿ}��iȖ%���;���m9�2�)m�y_�	QYc�%��ı/~�u��Kİ���{����O"X�%����~�ND�,K��{�ND�,K����e�rc���`ݧ�\����S��ܺǎ��[����ٵ�y�[���:��f���_�����oq���߳iȖ%�b|g{��r%�bX��{��~	�L�bX���~�ӑ,JRe'����Ium�9K�I��E���si�~��2%��~��6��bX�%��ߵ��Kı/�}�m9ı,Op����n�R�`\ֳiȖ%�by��siȖ%�b_���iȖ5\D� �=��)(B������
�hf��8�9���D�
�F3X��H� ab�!!1 sN�iw�&�wMP�B1e@�H�V��e����T%�M��` ��FI���RC�;	�Ԣ�S��>�b���RF�QB]�����$B1�}%(�`��KIT�HPP�%��Ѹ��̓Q�U�vt;�����jk),������H� sy�e�X��"�%d"@�V4R6V1`H�e`�ְ%�������a�(]��.h�M�N��P=P�@+T 'C���Q<Z��>����@~<&� P>�������B�¡�#�q=�w����"X�%���siȖ%�b{�Y��N�u��.[%��m8Re&xJ�W���)~)2�)2����(�Kı>3��m9ı,Os��n��)2�)5��Vۻ��B�F�ND�,K��{��"X�%��=5����yı,K��ߵ��Kı/��u��Kı/N�}s���Y���1v�jx8�P5����-��n�jykl�����q�
�\���3_=ߛ�oq�X���6��bX�'���6��bX�%���bX�%���[ND�,K�=�w��92��S0��]�"X�%��w�ͧ!�D�DȖ%��ߵ��Kı/{�����bX�'�u�ݧ"X�%��w���ɭZk&�e˭fӑ,KĿw��ӑ,KĿ}��iȖ%�b}���bX�'���6��bX�'zh���e�Z�сn��m9ı,K���bX�'���siȖ%�b{��siȖ%���"� xZ(@�@�*�����O<�����ND�,K�w6��\$���NR�Re&Re,�{��r%�bX��{��r%�bX��wٴ�Kı/�w��r%�bX��UK���󉻃.�d�r��Ŋ�;wvA,=��9�-6�ظd����7^.�.�7.����,K��?~��ND�,K���6��bX�%���[ND�,K������Kı<��S'm��ї-��k[ND�,K���6��ؖ%�~���ӑ,K�����m9ı,K�{�m9ı,Jt���[�\!%�K�)~)2�)2��ݜ���bX�'���siȖ*%�}�{��"X�%���}�ND�,Kߵ��j9"� �e˓���I��%e-��ٴ�Kı/߿~�ӑ,K��{�ͧ"X�����3���[ND�,K���i��M9-5�[�sY��Kı/��u��Kİ�߿s��yı,K�����"X�%��u{��r%�bX�@=DA�b����$R�4�(fv�_�ֳ,09^Fz��ٽ�ɺ흹'E����TY��8��S��5�v�`��Ͷ6A�Ϩ�%Cml�mF6���j6���8��l�ע��;��d99m�Fm���n���#������Q��n3���<�sE'S�TTIkmbk�H�QYܹ��\]�q�X�@���GE���!:����f�B��f��4�
�uif���غ�YҾ	��W#��5nJ���ݗ5�{9x�[a�t�{�^����"�u�͑q���w�w{�����ڃ�GKY��Kı=��}�ND�,K��{��"X�%��u{��~Ry"X�R���|����L��^�}N��QZ֦ӑ,KĿ}��iȖ%�b}�^�6��bX�'���6��bX�'{��m9�*P"dK�;����Iumܜ����L��[����r%�bX��{��r%���Dȟ�~���Kı/{�����bX�'�N���7F�u1̺�m9ı K��{�ND�,K���6��bX�%���[ND�,K������Kı<;��k��Z�e�d��ͧ"X�%���}�ND�,K���bX�'���siȖ%�b{��siȗ{��7������2���óƣ����n-Z̝v��8Õ�9�l����p����\<�n���BK �R�Re&Re'��9K�,K�����m9ı,Os��l?
�șı?~���iȖ%�b}���D\�V�r��/�&Re&R����m9���"%����`.�J��\4�@)����dK��ͧ"X�%�߻�ͧ"X�%��7g)~)2�)2�i1�zY*�Ԃw2�iȖ%�b{��siȖ%�bw��fӑ, �,K���bX������)2�)e��a#jY)e˭fӑ,K?02'�߹�m9ı,K�����"X�%��u{��r%�b6'���6��bX�'zh���e���fc��
aL)�}��ٰ�
abX~����ٴ�%�bX�g�߳iȖ%�bw��fӑ,K��ޒ3}��#vp�t*��iz��l�ڶ�ۣ��1ۗP�U��O����{Vój|�_=ߛŉbX�wW�ͧ"X�%��w�ͧ"X�%���}�ND�,K��{��"X�%������MѪ]Ls.��ND�,K��{�ND�,K���6��bX�%���[ND�,K������ı<;���w-�L2�\�fӑ,K��{�ͧ"X�%�~���ӑ,y���(B%U`!����wW�ͧ"X�%�����ӑ,��L�֣��D��!%�K�)~)8��~���ӑ,K�����m9ı,Os��m9İ?�"~����)~)2�)2�l����\���"X�%��u{��r%�bX~D+'���/�L��L��{�9K�I��I�~���ӑ,K���Ӷ�B��ë��K�C6^�h;K�mK���RxR�csiS�ܱe�����<�����bX�'s��?��r%�bX��wٴ�Kı/�w��r%�bX�Ν�m9ı,O��;�JkV�ɪYr�Y��Kı;��iȖ%�b_��u��Kı;�;��r%�bX��{�ڿ��[�e&R��^��.B(�$�iȖ%�b^���m9ı,N�N�6��bX�'���6��bX�'{���_�L��L��f�	�.][w5��Kı;�;��r%�bX��{��r%�bX��wٴ�K��O�Ԥ��q/�]���H
ke�v��k���<��k���Kı>�{���7F�u0̦��ND�,K����r%�bX��wٴ�Kı/�w��r%�bX�Ν�m9ı,OȂ{��3,���hK�O����xbv�/
���kp�5 �	�u3�G��!jݶ��K�)2�){��ӑ,KĿ}��iȖ%�bw:w���$|��,K�߿siȖ%�b��3W�.��!%�K�)~)2�)1>�]��r%�bX�Ν�m9ı,O{��iȖ%�bw��fӑ"���H)f�~���؇n�.
�*^~_�fĐIϾ�I�$��'��xm9ı,O��{v��bX�'���̝�4�֡r�ͧ"X�%��{�m9ı,O;���r%�bX�}���9ı,K����ӑ,K��;Ӻ���CY5K,�kiȖ%�by���ӑ,K���w�iȖ%�b_�>�bX�'��y��Kı4q6����{���������cg���ϗ��v��/[�뀮-���&"�I��4�1�՗��96��c�	����9l�;]l����qʋ! ,�^H�;DE�9ݰ�֩�l7g���5ɺ��[����y�w4J2���#������V�g�5������-��'�z�s�B�>6��͜�t�C&B�헮���ݶ�Fnŵי��>��������^qg��Pãj��[�8��됍V�틣dkj�+ϕ���nm-Z�4�Z��}ı,N����9ı,K����ӑ,Kľ���ӑ,K����"X�%�N�w���3$�֫&f�ӑ,KĿ|}�m9ı,K�{�m9ı,O;���r%�bX�}���9�̉�,Op���r(�Q�Nڒr��)2�)<��9K�,K����"X� �Dȝ�~�ND�,K��kiȖ%�bxwW�\�[��e�e���ӑ,K?(��Ȟ����iȖ%�bw����9ı,K����ӑ,Kľ���ӑ,JaL(�>���Y��n�U�l8�,O��{v��bX�%����iȖ%�b_{��iȖ%�by���ӑ+
aL;��Y_�������%�f4��"+QٳQ�����u�P8<�W�خ��̿! \���]��_�L��L��l�.D�,K���[ND�,K���6��bX�'�k��ND�,K���fNܚrZkP�0�kiȖ%�b_{��i�zs�`i�"dK}�6��bX�'�뽻ND�,K���u��I��I���V���!K#L�rNR�ı,O;���r%�bX�}���9���2&D�����r%�bX�����/�&Re&R��n��q�p�R$Ѵ�Kű>�]��r%�bX���"X�%�}�{��"X�%��{�ND�,K�;��kD̒�Z����ND�,K���u��Kİ�������yı,O~��iȖ%�b}��۴�Kı?w���Ja)s+<{s���$�Bm��x�����nTM:5F8�V냳�qtqg��=���7��b_�~���"X�%��{�ND�,K��ݧ"X�%��|}��r%�bX�Փ�gun�a�-��k[ND�,K���6��%�b}��۴�Kı>Ϗ��ND�,K���[ND�Q�}��ʬ�m/[��6abX�'�k��ND�,K������K?zu����?�wh���� �a�Ԅ�l(��|v'"^�~�iȖ%�b{�p�r%�bX�߉ܽԚ3Rf�.k3WiȖ%�����ٴ�Kı/߿~�ӑ,K����"X�%����nӑ,K��'ݹ��֡�)�B��5�ND�,K���[ND�,K���"X�%����nӑ,K��>>�m9ı,N�{��;g�t�=����nX�\�YLv�F��T���=*ڶ�E��lU5�e�n��˭kiȖ%�by���ӑ,K���w�iȖ%�b}�w6�r%�bR����R�Re&Re-�Fm\r�;�Q&��iȖ%�b}��۴�? G"dK�ӿ�iȖ%�b_�~���"X�%��{�ND���L�b_�~���։�%֣�����Kı;�;�6��bX�%���`"X�'��xm9ı,O��{v��bX�'�O����E֥&��ֳiȖ%�b_{��iȖ%�bw���ӑ,K���w�iȖ%��U6_���W�
!�8��5����m9ı,O�ڲv�[��e�e���ӑ,K����"X�%����nӑ,K��|}��r%�bX�����r%�bX��u���o�4���ͦ�sJ�"42N���g�*�Ky�`Tm:7On�ȴ�N��&]h�r%�bX�}���9ı,Kߏ���"X�%�}�{��'"X�%��{�ND�,K����5&��asY��ND�,K����iȖ%�b_{��iȖ%�bw���"X�%����nӑQ�,K���.^�1-�3���6aL)�0�~��6�bX�'{���r%��dL������Kı/�����r%�bX�g{٨\�Bf�feֵ��Kı;���ӑ,K���w�iȖ%�b^��u��K����G"g߿~�ӑ,K)2����U�.�E$��K�I��E����nӑ,KĽ���iȖ%�b_{��iȖ%�bw���"X�B�p��=Z� ;�D���
ԑ��A�vgЌ@�DwwX2 �Q"��Ș4�6�	6"���a5$���^t��ETG\��7s[�𠯚@"D��`�N8N����Fx!T��ķ��*��,|��Z0!��x���C�<|�Ea��mv�(�~R��F80@Q���VPU�r�ә�q=	�ﾆ���@,Z ���>�E�D1�`�I��*#1J"P�F �,(0�hM0�i!�(�S�	�4J��y��%�K�"�ϫj�:튂0Fy$�`9�>��@�	� ������ rE�%   �6�	��� &�lE<�����1�($g<��Wd�L^]Z�-Vѹy�gٗ��FK�����̧!չ�qs��mGL��S��P=���]P��ͮ��mhۮ'X�̮�.��DM+�����>�T�T��.q�V��h��N;0�X΍<ő	t��b�("���5*�R����n��^:�7�L��y9��,���Cn�([��9�]Zv�����ێO<\��yv�O[����;^��vy�Ƽ�gN�[8sٍ�Rs����O39����NL��nɹӧ/k�'�`{2��"Us��G6�P��D����m��B��EP��.a{����͵�!)��
\�D��]�8�����ά�Cdr����@�d�ncڂ����wQ������撞۞@�#p܊�3���n����n���M��&ˈ�8:�
%nI˝lF�hQ��,�PІ�6�Ӊ ^�nP�:ح�Pҙ�u�bI��&�t�oA�W 407�������7-�en4�#�e-��ZWFƻ"�&3`�.x�7Wmƶ6]�{U��A���u�������h�źdFG�\:����[��nXm��V�4��cU��s�S�zjv�O-v�%6к��l���wm�m���8Ӥ3&��=w��R�o]bv��g�N��.-�7(-�NK,��6R]R�m��멥���s�QQ�����&t�:l�\JtԔ�F���e`��If�մ�J<N���c�
��ST�0˶�	^93�]rQQd�ݶJ�YT��sO �
fz��eS.z�*uᐝ��5���ѯaࠓU`9����*�:%��55m�	�Yk*����H��r�5J����s��V-ؤ۵��9J(�p5WP�+�8j��\vv��A�un�m�a ��a�p02�#ȝ��u-V��,��gś�Nm�f���9&$��)�6<pR��ѻp��Yjشf��;ݽ�{�w{�{�p8'�h=A��T��Fx iD�ER(@"�F0HA�ň�Z�!� �� �0D��"`|��L>OHs���w����˫//.�[���v�Ng�W(�i����dM�ْʻ���׷m��ζ���\Fy�zw1�w�\Cx�
��c=l��I��`�w:�&˵�-d��Dr8��%�0��=��l�ݗ�Y$۳�`��I@R�	n��J�]�0��k���9�2d��zq�@��FE՜C�q�bݍa�'������e��ogD��Z�Sr�􆄹�̼'d�Hf-�t%�u�it[T[tO#�pi�I/H\=��y�z<5ʶ��VW>`^����H��r����&Re&Ry�{��"X�%�}�{��"X�%����6���DȖ%������K�2�Z=��qD�!i�RNR�Re&%�}�{��"X�%����6��bX�'�k��ND�,K��{��"-�bX�Փ�gun�a�-��k[ND�,K��xm9ı,O��{v��bX�%�N�[ND�,K���[ND�)�0�����Yw�M�����a���������Kı/�����r%�bX�����r%�`%����6��&Re&R}�۽���Iiܹ�,KĽ���iȖ%�a�9��ߵ��%�bX��~��iȖ%�b}����r%�bX��>>	g�W,��jh	ٸ����8N��]\��\���f^&6[#7j��J�6��h�n�Ħ�͇XS
be'�{Ӕ��I�=��ˀf^k�07V����N�Wdi�nI�3�پ >�B���x��y%�:���x�#���G�����v5lt���%�, ��x�#�$�+  I�`�>e��J��7c�$�+���s� �G����NA���$���' 򥻻�~���ř8�_Y�И�r�ڎK�K<��R�y%��rob�FPYq\��
n:.ݧm�R���7,�n�rO����.ͽ� $�������6W��n��릒n�m�X%H������\��gA��E�$�r�|����5W��٭��Hu�B�6�N�T�4 �y��暯�~��^�;wo�[R	�j��y%M����n��pݾ��z�7��g Ʒ4�wl��Ʃm��I&Vͽ� $� sv<�4v*IZ��E�	�N�2��;�.�0e�G�l�!l�C�U�O_���{f}c�lLt��� ��T� ?w�<�~a�����B&]�Ĭw 3d椕$�5�v��� �/���T�g]�Yr'pj;Nڒp[�^$�X~K}s� =�����A�\i;.�Z�v��$�Xe�X!��܀��*	��h���{�9��:��)^M�+�餛���, ��x��x�e`Em�%���΍�.�O��gY3�C-��=�Ժ���Tdm��<-v]����m���lWd�I2��}U\A���Dz]�֢�յ �v�N��e�ʒl������| �Y��^UJ��5�����vF����{�\����&�ջ8>�� ǈ�T-��Q"K��}��|,��f_j��*�{��p��ߊB.���j��"�%��%�}��j����j���� ��`B���s�=绛~�~��K�)r��6"��9���k�=�������0�t�����ƕ���vkr��gA�ȅ�ٻh+A�i�������v��"秣�`�DGns�z7"��-�H�|tܕh;v�aѭ�s��zN���ms�xM\���iЕ�[&�<7lsM0�&\�h˰N%��M�c⡝n��c��m��?�8L�YV#��Z�ͶǴ�]vu��n��\mt��m���7�hqHm�JE��g���@xv��}����t���7p�o��$�+ 콋��}U�^�z��h!W擲�դ]ݻ�$�+ 콋 �T���:��)^M�+�餛�e�,)R^��H�7g ����˩��E�m�i�r, ��x���	$����R��xG�ݯ&���H��o ;ݏ �^����>�� 3d�J���f��x3�k�؍�{r�,����/h���wV�aۮl��Mɫ����zۇGF� �����ٗ�ř7ԗ�f�pyZ�T�nD�..���|J�_@G�J0�E|�iځ�"��� n��	$�����"�.R��1�̾������w�{�\�=��:3'r' �v�ڒ�=�x�e`vK�"�%�]�UƓ��դRV� �L��Uz�޾���� �v^$C�v�I1X]&���:8n֘�΃l��e�q��l�E��{+%�㳫�:bn�]4�u�E�/ �B^�l�X+iK����n�heۼ)	y�#�O^��e`vK�5n�D��)Z��n��O��훛<C��B��/�� ��i � D�����@����\�/ 9��t�2��0�cT�ݻ��K���`[�^ I��e��]ߥ��;:��u�E�/ $�x[��	$��9%Ãl�wV�ЁL;b
N���sգ��t���֫g�	2ACj@�8"F2�.R��sM�-�x�e`vK�5|H�+n�bQ�v�' �����vn�P}ݾ wM����Hڮ�-.4��V�"��x�{�X]��l#�"ݗ�qT�1�,wV����*^I_�{��o��ܓ��f���J
�����᪽>+���UVa�Ӎ�^ M�x[��	�e`vK�?}��R[�\�j�`㸈���as/| ɭ&�n��n9���6���h�w�[��w��ܓ)v7�����&ɕ�E�/��R����������jp�2Ir�	�e`vK�	!�m]HS��j�t���d�TR<-�x�e`����"�-�Bn�<��{� �׀I&Vd���E)[t�5+M�-�x�e`vK�5E#�;]����J�wh����nhF˱�;:��N�V�ʃj$�m���d3����Q��e�,]d�J�m�mu���e��۰��^�g�Z8z+�a��Lp �7\�����˼�Lq�9���OFۗ������God��8M�G<�ڹ�鸳�ɥ�����u�+K��qśQ�݌v��+���5P��]8��5��3����v�:�e:�9�]����XB7]�^O{��d#>xٹ�l��v�;s��K�\�s�U{N;[���e�dz��;��e��՗We�[o�{��V��/ �Ǚ<���3}8Z��rK��I7Xd�TR< �v<I2��M��j����mȡl��>�^���w'��]��� �_��Y�wf9BT�)%j���c�$�+ �nE�j�G�E�Q6��aVƩj��338���*��=��������N�>�w����-�Ҍ0�b�������B3ιغ�d�ֳ�IvT�q�g%G*����܋ �� ;ݏ �L� �]���"�-�I6�QH�꾪���B"<��)�Ph T�D�L_x"���z"�����n�p�^c�*M�tn�N�ة��Zm����$�+}Iwo�X^^��6��KK�ݫ.����וR��{��p��πu�̜ ����U([PC�Я릒n�v�X��x��x�e`���H#��Ww0�h��7	2uFsuj3%S��lv]V�py�(OWb����w�����!]d�#�_��� ;ݏ �L������ȝ	RLh���o ;ݏ �L����)z�ꪤ�-��we�
�5H�V��{�X;r,s�Wܥʮ�CZ���a1u�\B���P�%Rzo`a����]�<���ĩ��^����f��P�r�a	�R2$.�y.���8`N	�1���;` $��1�� ��#*^��`2#� ���tO_�̆ב �l��8�Ve۰t �$7wg�iW��6
 �pA��h݉���Wd͐����(���4���>OA"�#SkUQ#��TSh� � ��}Z(� �5U*��ڋ�ǀ$xda��L�:uCv� �nE�j�G��ǁ�R{��� ��%��������x��x�e`�Ȱބ�]��xsۿU	:I�:�b⭀��.�c��[��iѪ0�gj�p{1p����U��}���338�ﯸ�U/*_Xk��� Բ���%۲��c��p��.y*l����"��� s��R��ն���i&� �ob�5E#��}I��{��V rKH��M�-P�[X����ݜ ����ffqp"���BIZL"!�X�7�mj�+�]��m7�۷rp�{��m*T��{߿v��{����x6�H*�i��p��:������3z��׏�N�Ҷ��h����m�hmݗL*��"˶���V�ݗ�j�q�;��SiG�llj$Iqp�������vk�ߧ ;���3��.y%T�lWw@��]��C���/� 9���������:���_(�n��SW��?|��� ����8���j�q�Uۥ���՗We�6�7fV��=��z_� ww�nHg�O��b��q��]���G������t����V��\�ԁntu�9�dy{\��N�un��`�6.u�(���X��Avy�/9��Ѻ�St�;�;Y��������c0һ�=��2r�Um�v���mE��!��Wh2rn'���\k�z :��y��h)�Tk�l�Y��[ی��nvk�k3�9�u��؟gO�)�m�Ƚmn��_�� ��zNs,�qL�Rڭ�Isk��@L��,�K��v�QMkf�-�M�<�Zk۟]�f�������15m�:�i&��uw}x�� wv?��A�=���Qy[���Z��n�Sn< ��xݙX�xқj�&���I+v� wv<n̬=IuOz��/� �����t­��]������Os7��<ݾם�� ��x�Q��[:��u�ql��j�q�wc�'ve`J.�����_g��@�-����Z(�g[<OG���Dn�
�����M����7����ۏ ;�;�+�_}�S޼/�y��*�*���^����7�l`�k�T����sx��7o�}������-.7m�]�$�x�̬�d�?UW�_%��~� �<�UmAZ�К��r.�J��}��_ �^߯�w��	ݙX�В�.��n�j�]��;/n^ wv<wfVŲ^ n�Ug}8�l6������:�y苫�{̰n�$��v["Ѩ2�~��?�p:7n��d��'ve`[%������5z_��iںaVƩwm�vef�T�6|�v�=����ܜԪ�^���ڟ�9�@����:�޾�o>����DF*��0#$��# �~�I�?��sU���i���}�,e�\�9/��*O2n��s6p�L��d���bR��V�M_��w�ݏ �==��g����� �;�n7o�9��sg���]��n��g=�Dќ�.�4bnz-�N��qf��\��m�{�+ 9�<{r;��ǀuV��j�Bu`ƛ0�#���}UI�<� 6O<��ﾪ��-�$��ۻM�����=.y� wv<��͑��`���J�+�k��/U�n�p�g� ~�d�}IR�E"�G�6!Tp�J�BQE�P�.�ﳗZ�;~_�,��	�4˻�8}ه �?�v~v�n����M��V��ՠ��V
�Sa΀-ڧ�����l����eYf�Y�ٷ����c�7CV���i�����6�`wc�$� �]�v"�-�	6���Xٱ�k� odx_R�mҶ*j�e���c�$�?|�R�ٹ�N�/|�W֟K�$�We�6�&�`�G�l/b����Io��ݺz�+�n��� 7�' Ԓ���?�3���3;0�T�g��;���w{�~��r�̼4�5�/��[�w�M���7��\���1`�7>5��by������:64�;t6ˌ6!�%-����lp��5���Ύ^��6ҚE�t�Och�tq�v���Ɲ�gu�m�nZ�;88Mok��t]���ܘ���,���L���=:nخn]�������{u��t�/qux�\��b�#����j�6�\��eq�Z�ɝ�n��iւ�4.�0π6�*�6�Z(��2�[�/k�G�����y�E�حOT]�aS6��������7�tRv�@���E��&�<�$��;�83�Z��c,mH1��| �;��UUU����l���zp��X��#L���;�;�o �\0{#�6�`fǀE��&�j��}m6`�G�l/b�͏����sN -]�#r��8�Nٱ�u� 7�<�(�\.��Mn��θv׈)�Os�q�<�n��%��]��ɞ�r�H\����V�ٱ�u� 7�?q�O����{$��j챹$���9�*K�����#�6D��~��ꤎˠ��ȭ��D��wvp�\Ç��}<�H�`�CB���i�N�N��y'�����͜>�Á�T�wv`����wISb�m`fǀN� odx�q��UUKtQ+�.t��/n��=������gum$����͑q���w���6��5ۅ$�-��?O?� odx�q�\@n�`j�j��nݍ���f��L�^���<w\3�}T�C�<�n��ci7w/�f�������UKI+�N��PV	H�����'V�/��J��[Hj�m���#��f����=J�%�IRW��ޏ�mz���$��j챹$��f�*ۓ��'��X͑�؆��v����ְ���h26z��x��\=��e�u7n8lazd�;m��+\�v�|����l��l� ��whhRӶ��N"˒�s�#�*J�a�n��ɧ ���|�*M�����]�j j����'u� �ݗ�l��e��.;���i����z�����y� �����̗��$�RB��T��\UIuVU%���NN�ݩq]ː�>��0��xˑ� sdx�s|��x��-=�!k�.&��[���x��t����s[<�$�;=V�k�6;�J����w��;=_}�ꤩ}a�w��<��G�r'q�;�w%�6G�N��v^��w�o��iq�ݲ��&��'c�ջ/R��o6�e��ݜ��Ń���J�� �ݗ�l��6G�N�wh)i��o��ۼ-�W��;0��x��*��_�V�FH� I�n�k_i�8kQ+&��$!�0Cl6�����0M�j<�fV""2eTVSB�j�HC9\��H\��I�B��A��_�ξC@x�!�/����"�H�'�ӈ �(ݐ�)�B D�b�(m�>��⾛ТȬ2��0Ơ�`U�/6�
^q��}��=@�=�
�����1�0�����A�՛!B"��h� Չ0a#!4J� ��Y������_6��`&Ь��|8	���JH�P�66�n��*Q�<�pٰ/���j�k3Z���  @ ;mm�ě)�WmU�J��t����ֹ�7-����S�l^*�k���`��y��C���ղu�6X짦�۷/k;n���;K���=��t��ݰ[U��ga�n��I���M+�\��5_�|��5[(��ؠʨB�\�������˰��LN��{[n�`e����*�^�8�,��.�,vgL�'E۵�b�8���q�c(�H� kȜ�Kr�N綃uͶ�{=��g�i�ʥ�7e�8q�ǇYj��|�Y�&`v��/b�E�uպ�- P�c\�d�:�r�v�1:�r�L��n-s�	�6�Rb�:9�G%�y{ɒ P�D�����N���;/8 V�g�I�.�<�A�WF��[���sF�t���Gq���v�{���N�p�U��kn:�{v�ذ��A+SM�dnN�WZ��fÜI%��B�Pˎ�A���*��J��r*8W:Sb[�;���
-�V��5m�CP�:���M�p�E�t�ݍPJ�]�/ �u��kcu��rkh;c 
��Gm.1FN�]-M�����._e�j�ƪ�i�JtU�݄M�F�F�]5��X1�b�R�j�J�t���ͧ��'����GP��ۊ9����F�8�:��֡Ħ�Cq:C�
�c@e1�nY6�@m@^�sv�V��J�cs�ېv�l=����qI��"Yz]���8U�ڮW�?�هe�tY��%���\vv�j�'�ő��^�%� � )�ka��T`��\��B�3+_
!�'Ͷӝ��b���չ-wl�I%�6٥f���P�(��W��.����m[n�p3�t���v�ذ*�y��+���e�.���Y�� R��%vd�]��Ef���`����n��y���EN�UUeܫt�\MG9q�Q�UuS���G�m"��Rq#����U�9�ذ5T��t

�b�7Gg �f�t�:��z��1�t�j�5�]\�K��(4enj;�����������*��!���'E". mQ�U4��h��? |*P4 �|�}��>�X��fe��yY��6�۠\k�y��usr���L��u�pp���n���;s�-��6C����j뎳�[�;g��θ��t�[˓����1�nP���K���ʧ���B�dp�P���g��+�7C���G(�Z�u5MNHG54;��T�=�%���Χhr<EQ�h�0۲e�zy��8&����B�S����/)m�6 /[i5J5wM\XnO�;W/�I��Q�L���;�9I�a �i^,�RU\�i�E��m0.� �~x�p�:�e�nʼ�
��TRv��ݷ�N��v^����N*T�J�]���ܹ	�9 f� ���T�6}���o|�`��0�4��P���"ݕx͑����UW�l�x�yAz�ӥm!��v�^ sdx�p��ǀE�*�u%����\��0�t4�ն͗�pvw^TU{N;[��he���<xx��m�.�ʴ6�;0���nʼ ���۠�+�n�:T�m�$�{����&
E	qN!��NҤ��$��y����}�8}�z��7�
'�.ܲJq
�I�5�j� sdx�p��ǀj5R�:.���#]�|�Iz���N�����ܜ%I=��/�u�X�Ƅ�i����'c� wv<-�� ��~�>�x���[��[0�ib��Q�9R��[<��v�ќ76G�.{`msv�M�3�>��0���l���%���}�l=��8��z0����w' �����T�Sf>�� ��Ӏgrsj�f���[�J�CWN��x[�^;�� ���1�Aȏ��TJ����>�_ۥ����^I$�Z�ݹ/��O{�Ӏ���1�0���/ ݺ�B�[t��N�ـv<-��.�x�p�;�`��U�ϫcg����	��뛑�ダ�;.��o6���`���weۮ>2�����W�S�/ ��^;0nǀn�(ڎ��uwCE�^d�v8`ݏ �d/ ���M�Rv���w/�g�0�w�8m*I�y�_ ������w*\N帤
��8J�����'o����<�=��OW�z�jG�n��|I�� lD�P�I���v�����*�]ٚ��٧ ?w2p������<9�7<z�M����H�4cp=�vS�����:3YW�gDt.z�4=7l��{;0�#�"��2���y$��j�V]�|>ɇ<�%T�}���k���ݾ��R�l̴���܉��"Hp;�8>��ʕ|���,��� ���IGi'M��v��"��&�ŀN� ����.��]ݗh�Ar�3��|�J��w�~ ��������)UBJ����{��8��Jd��g���mٌ�v[y�m�ӍcP��f ��9.ś��+�;�F�X�� �ٺ͚�6�\���Yɣ�ۧ��y^���et���n�ok�F:���ut�nRU�c2�n��n�7.z���gt;��*�X�S��El�]m��N�Nk�b�!���]=���$z�LN�n;[9�������K�f[v��Y��O���uϏ�l��(@;�|��-�Bݗ�VWZ��YǍZW�����h��ݭ��VF���:d�=}�N gٓ�u�!x�ذ.�gͺV�:l>m6`}�9�U��+�^���m� ��0�6[��q8�$Hwrpy�_ �{�0vG�j���t�ն��S��^6�,v8`��}I���|+m</d�\.�j����3�� 'dx[!x�ذ	J(.�mV�`SN��nK�h�M8�9��"TU��u�頴������\�ڭ��<-��m�X�p�;� 7��qIN!]�8>��W*���w�h�{�� ���������ݗt4P[e�ob�'c���o��)��w��剴�U����k ��;#�"��&�ŀqQݔ��ܸ��H�8�fN�J���t��s� ��:H	wV��j�r#v�y-��݆w3��vx��(�RVU1�8�e�V��M67T+���K�&�ŀM�� =���<�U{�t�ն��S�n�	��`�� 'dx[���]-.6۶]���]��N� ��}��L��2B�zUM�&
h >��pCH����Nz������m�N�:f N���e�ob���T�����:+͡:o�tU�o �v^6�,v8`$� $'֩K����'\(`�����Eێ�s,�ٞծ��jv���j��t4P]��7ob�'c� N��U\A�'� �/���n�j�b�G�3�sUU6���5���	��`TweRn�����ـ�<-�x�ذ	��;R4X㐒��_j�������3o5�_��|��0�A��FOB�I�C��s��~��}�f^e5�F]ۼe�X��j�/ �d���w��ߧn7~���^�v�v�Y��䛫q2�}/��FYQ�L@�����'j���Uڻk�zy��5M��E�/ �{���m�N�:f�l�-����`c�{�6W��^m	�+����S޼��,lp�5vK�7m�4�Һ(.����`�� 9$x���O^�\����][GͶ�	���<-�x��]�>7�:��x9���E���n�=���~���S&{37c�OMs��-��t��[OX��;_�|����<��ۑ�]�[&�5��xwb��Y���+�����;�6.R��x�r�u���v��bk�d���U��6x�Z��]�
T�N���M���`��㇮V�É�E"��5{�>S#�Fm/cv�M�9�-�5�0B[�PZÌz4Hm��s�v��s{t6�������L�{���C���'�䥶\�)�̆kE�l9ŀ��U�x�x6^�qm��I'f�\,O�خ�F�����ۿ��v�,v8`ԍv&���x[��	��`�� 9$xUvTwM����S�n��ذ	���<-��	R�iq6��]]�v�������x�}ݾ�����T�{7_ ��եڶ�'J�� �엀E�^�܋ �0�߂}�dIRv��}m$\9�7k��u�8�ҏob�=Q�e�M]F�n;s�ڛhN��] �� 6K`s������������6��Wi]���>���P4�$V"���6A0_D^8<T���'�����"�^�y꯫ꤎ��k�m����4����O?Wd�-�����TweRn�����ـuvK�"�/ ;�����յ�44;M��4ۼ-�����c����o��ݻG���ƪ��Ρ\G��r��1��%�z^�L��.ӸO]sHN�;�w�� �0��x[%�[t��6��]]�j���&���^�x�����"T.շI:T�m�Wd�-���U_�]��X
H��d
i)� a�!UłsE�df��",$� �2�O�71���L�aL|_�m]P��B1C �r	���`.�0��c�O�y�}��ׂ��$>�rC�A���`W)��6�E<9�.�D����>x�	����1S�B��HF HA�Y�� �#1�A�<P�8>FX��3O���PE��^ a� 1"^M�饛Cf��Q!F��@ /���K�p@|����8*;`��9�k⠆����!ኁ�C`l�)��DH"�������nI�8`ߥ:*6�����n�<�s޾ w���gra��T�7����FW�ZJ�t4P[w��68`$� �d� �R�RB�ӵv�h�{/n���{Zlq�8{#��[Ir"�;6E�Wg6[�M�uv�T�o �0�G�E�_�磌�	'�����MҴ�46�0�G�E�^ odx����Wf=^�q�,q�H�wrp=����68`fǀM�ZGt�ձ�v��ۼ ���	�� ;6<	U�?�}i��O6�����\v! 6��ҫ�|�$���o �m���6��]��զ�7&ԓ����k���~̜�/��|r�����Z��fУͮ�׶�r�{N;X�h��s�`{�%qؽ:Q�K��M� �O< ��x���︃����Zdqے��;�p��'5/*��zp硫 }���$ٌƞ-�;v+���m� ��<�0�c��ǀw��qZl�Wm%H��UUU?�y� ;���w�8���=��5�}䜉ۑF#���ܜ ����w�U�ϝV���&J����;~��q���K�)r�v$�m�[�"�]^|���)vγ"�Y�Ӗ�{������ڰ�ŗ�.�u��v��ۃ��gg;��n�o�Si^���WD�g�s�c��u�Q�&��7g�[s�
����N"��e�6+\���q7d���d�]Yz�m,U[��mm�mr��/�������[���Qs��pFg^�&@%g{\�\�-�[��e8�ES	�@�j�;G����h��l�Q�Չ�����g��9lg5�͔B.ƪ��	�Vm�ݷ 9����G�sc� vlxۥ�wN�['j�V� ody����? ��� }����*lն�[�Ir�,�V�6��?ٱ��䍓� &�� �j�T�V�Zt�؛xٱ�wc���%��<mx��V��]���ݏ 7�< ����c�9�����+�+�F͏�ac�]y�����)<� m+�6�t���Ej�t:E[m�o���#�͏ ;�ޗ��i��]��*˶�	�~�[�q�pTO���آ�﫬;����������[���7m�fǀݏ 9�< ����R��M��v� wv< ����#��ǀM�ZGt�ձ�v�%m�6G�z��v{π'� wv<�_U}��J���SV�����]�#�s��:�Nӎ�᥆ضX��$G<qt��6��]�h�� ;=�ݏ ;� sdx���J�ڶ�ӥN����ǀݏ 9�< ����W����y�զ�WE+m���߾���7T
�o�6&�Tꨆ������;��'}��ܓ۩Q�Z��]�V�x͑�6G�ݏ ;�ޚ�&�Uv�H��rp�s' �*����7}8���������Ï��2lt�a�1�ij���=�P���y�#�=r����s��\��t�|������wc�l� 9�<�T�Кltꋻo ;� sdx͑�wc�$z](_���Iڤ������ s� wv<R��Pm۶:�*Э� ���W��٪����VI���HNA��@�|D��W�e�x%�KJ�ڶ�ӥN���}ܜԗ���������N�IW��w�o�ߪ.���;<���3���d��ۀ�6]6#l�6�	��^8�������m� l�x��x͑�︀��< �J�^ui]�t4Xۼ �v< ��������y��d�y�����+�lWr��wޜ �����7י���� բ���5v�4&� ��xV� ��x��=�uz�y����V��ݗ�~��<����5W��٪� vFA�WaCU���r�U��N�T���2��ul��`I�x�x�̞�nNu�xt`��M��*�����˿�w��vD�[�]�H];@6^�>��5y�Q�r��v�m�ּ/�a��]�s]�êc��S[G��z�d��I˛�ڍ�;���^�s Nӈ	�U�Se7����۞:��[k�\1���b�e�&]�	� �@�'!�$�	�[�ɐ�[]j4�	(Zq8�v�W�n����.ӣ5��	��*V[�l'j�v� {� s�< ����[=x�AK^v펮ʴ+o 9� sv<��/ 9�)#ʼү]�n�:T�M� �xWv^���H�x���%J*������)6��ݗ�ݏ 9� sv< �R�j:��Һ,�� 9���<��ݟ�>�l�?���<��Z�c������~r����pb`ǍX���I�\���u����Zt���A���g�� 96<��/ 7�գ�-Gw"�*G!��ܜ��.�*��1�ȴ��ZAb:�6P@�d	9�W��z������;�|�[R�	�M��Qwm�]�x����%������&�-.]7Cc�v�Wn�{���p�M� �ݗ�JSU�nݱ��V�[x�p�M� &�x���T�C�l��s�t�c���r���'q�ӞFbh�;u�j�%�4]�T�U���&�Sbl�}<�nǀݏ ���J`F�V����J�x[�����	��� :D�ڎ��ڻ�����{�U��gΨN�$��~, \I�%D�$�*U56l���5�6���IfY)�E[E���'c� s�<-�|Ro�͜�4��;�`�� ����e��c�'c���������͗;��ݠ�Kvyvjˌ�|p����!�(.r����u��S��u�]�}���^ ov<v8`Se��-�n�m%v�J���c��|����uzz�nǀE5]����N�ʵj��'c��6^��='� N���t:[X�ݧ"l�w�UJ���=�� {wӀ��8t&��/�#(a22
P�@9~��w�)�ݧi���� &�x��x�p�8�%��>�J]�T��\�e�s,M�rU��+��n�2�1������4��QE����m��rp�&��2�����}8Vi,��HЮ 2I8}�yUSgϻ�������NmRlƌ�)ڎ�E$�f�\��	� ov<v8`ԭ�&�M[�N���|����	�� ����9�E�B�t��J�RJ���ǀ?}�{}�}~��u�'������*���U�tTV��*��U�(�
���P_���"� `�BBP�P�P��AP��P��@T ��T"�BDX@DYP�+P�T"P���1�T ���B@T"�B ��@T �@T �P�DT$BDDY D@@�EB	P�B
�B �E��
�B DXB)P�E@P�DE�E dBDXDT$�DX�P�$*�B �E�	P�"1DX�P�0DX�B+H��'�P_�E@U�*��TV��*�P_������TW�"�*��U�H�
�􊀪�������d�Mg���0��f�A@��̟\���     ��9H    )M          w� ��"HJ�(
(QA*U )E(�JH�
�T�R�BU
(�� *"@  B�'     ��P� )@� k\>V-��ŝ��a͹5u{� ;��s<�qy��˛'!˻��}�-E�5\X�  �O�=�x�w C�_[�>��ޮ-^fq��w�սݸѣ�_GyzMsg�`�mŪ  �x    ( )Ea 
;�+�����Wqa�[� ���f�=�=�uy��e���-� �w�X�-Uū�}w�J��Z�s�-����qo^���!��+��=���_[n]����y5͞�O�T� ��    ( B��}�q���ם��s�ڝ��ӭ�� �=�=�W��i���nkݯ=�U� {ԫ����o�  �׎�w�x��^� {ͧ6�7���^��yn=��x} ��nY]����{y:��x�:^  >     ���}�;�t�q(��� g��� �A��� � X� D� `=
0t�@=(�f�  "t@�P G�'�&�@��(�wJP�J8�PQ���cN�h�i�:DiҎ���(  \@    @��AE�����ɡ띺�� 5�n.�NYy��W6�ҽ�>��ϫ����r�M�  mw��^O!�� �R�n����\�{����Z� <����^�y5�w^,���6���  ���©P  "������*��A�!��=U*B�Q�����UIRT��d ��)�R�  �A1JQ����'������������|bN��=�����^�s耈��AUO�U�dEW� "*�AUM���X�,,���?���L�L�]S�?��I��>�38צń&��wu�x�b���sZ���A&���h�Ӌw&�q�E\I�A�n��x�>������F��ș��*`ΆS	�3�e��M�j�)�X@�k�%1K0�)��Q�"|l6B^���4l#RCjs�k\�W�&�f����6nm��փ�	w�/7��*�ҹXQqd$!l��&4�HRB�3y���zoy����F�p��.��,
Q��
������d�la$
Xa�nc���H+��e��5並^v��\S:Iu�"��F��;#�!,H�H� �@#@>a t5��&M1'\d�����\cR��h��!�,���!�a�3I)��,�$$.������ D�Sz�.1��2q \9u��ٛ�c�i���)��Cf�P�)[%0m`��-Ø�kG�q����X�{�a���(ZbsJd޶Q��T.��Z��g'��2Ip�\�� �X�\h�B�@"��,�F�
N�,$�,0�  ʓ���q��#!�	+����;ap\�����&,�HmvδMJ�&$�%�B�w������>O���P�i�:!IK�7�m���>C,i��\$. 0D�D�0�bA���Fc8��2��2f�R�0�) T�`�p@$R�o7�}��ew����d��0���2��R`5B��Xfu�_h���-H��2�)	�i���}��`�E���!1��ִBa��Y�b���X-�[s�}�`�1�Fk89��#��J`�%�ֹ��?h�}�p�����$�LeHW! �(�a���	�,��L�?��'�BBt�����<(V*_8T�+�B`���Nr�N�������v���B��M��:�����'�U�LT�T�
����2�#bLl%i��.	q��r:�$���ή r���}w���a��>>�  N^hP���t�B��t�td�&�pH�~�B la�aɦc������ڨm��W��g�ZՏ*��uQTj�Ȭ���#HH�!	-��:.�����.	z9��#$����y���;�td�!BB!1�c;9��֍;�ۢH��a�����~�ζB�3�5�u��+ �?Z��ΠK����ě1��� �$�h���~�Yr�HB@�3�}5�6ʘg���>����@D�ƹ��Ln>�>��̆��Eǲ�-C)L��Hz�����0T�Y4}0�쁁]�ΩP�a!��z�c,��l�2�)��p�����>X��h��!LW�����0�5_��~���Q��(�������$�DR$ �X1X��Z�B4��9�ԓZ~:�@�B� @�
�ʑ�Ao������~���CF�N!	0 �u��P��k��B�R�o���� >9���F��-2@��)I|�ݘ�}�S ���$>Փy3�0�a��d$$$�0��0Bܘ��ːR@���HCa�ak�+
1)
SARA��A0�P�R�(Š�18!�뻮cYrŁ�dq
@�ɂ&F0����C)�~]Z�����Gr�B��$�>W�aa]��M���@��pȄ�VH	 I�C,$i#�HY��:1�`�����02�7L,)�4��1�$�D�a�bO����HY%��cd���5w�C�%B�Pi�	"%HH� ���G�h@j�d`I!jbB�l��4�̤�� Fs���6h�9�).sK�&����4`cZ1,b[όtp̄(��Y1��~v0�
0�l�\d`aWgF�d�BHJaĒA	�$�K"Rb��d F(���a$`��d��q�$r�E�Z��k$(�hHA�b��[3�� |ٮ���6C��BY��0���~tH�$HKA�y�nFqYn��7��f�/���u�D�w��:��I]�i�k[ �� ��'�HfS&P��0X$~���">)huIH�yڪ�*%��c��D�
�S'Rߐ=*�i�Id���
�	!��Ah	BvuR�*�I���V@���ƛ;�c�H�(BȐ�)$�n���o��ᔖh�ݽ)��kd�l�WTZ���0}7��t���(�Qĉ���!����!�[��5>X0�Ţ����#pb4p``l`$F*��	ɘt�5��%HT!�L
��^?0�Ω� ��@�P��@e��O�゙���$���C,@��͒2ۆ��`�@�d�1BB��������a3�CFYBT�#z&3������E�J�3&�
�ă�JM�c=��$B(sd�ni�u���bp���J&!�͘�ٟ�XQ#RQ�$q���܅�ahBH�1�!~H�B2"P��(B�c�\�on5�D����b��M��$"Q�$#��9&�U���)�"��z�$@� )	"�Q�1!�jR48����B$i ��P�"Hb\@"�$����>3L�A
I�Z2�H}2����`k�d��f�Db�E�Ks�0J�`�%0��`A�1�}�b���Ѵ��D�"�bX�HWi��aN��t940��s\�X�AaB�l���C�H}y�Na����J$�a����2�cy fD�D�!�g�Ƅ*�
�XT��O���f>�� �H���k#�&�pl�qi\|��$/��iWP!4d�L,8��$1u�c_`�̥vCI�B����"d��>4�D�d`�����~������F9�'C� �M! �GN#��k��&-�d&NŮ1�ȕ��L�@�&G�#x�;����p8Q�(V�����c`ɭ��\�����&5 �0H�7���WnO�a`S�]����Ml��-ɢ�,����o�7��}3�2�#de7��gCD�N����@ǟȁ/��*~��&r��	�\��>����o���y:A�@����y��RY�39���!`� R"����*D������CrF�0isy$�m�%�pv1j��L露!ؒI�$*Lh�>��Wn�D	��X�HI!38��7�Ć��w.>�²}�*B��c�r��B@��7�ݽ"U��@��G'BcLو��gvHt���5�ֵJHW:�S9���	�M�/��m�Cs|�,+�
CX�2o��4H^$�6�W_q�I�@n)�6bX�$�l�b�)�\F♐���/؄1�l�S}3
?dӦ������2h ��2�H1�j%�`0W&���&��I��0A��Ja�7r��6��e�p�I7���f1!���!��cq���d�]����x7i.,�Ƀ)�ލ܄l����ׄ���!$��c	�+�C
c.�F�,.x8͈|C
�dd,�0I\�'�6���2#�b0\j?|���%�7���9�
$
4�Z�n�I��B�#"�I	�B���3��`��e�
k)�0ŨB�C�+�	c (@	)q��'
��^CJ�LB��B���"H4�2��+V�\�Ѡ�dC1_��P�$i��� �S���ܹd`�)�C5٩�!�$XaԌ�)�Ʀ
Y�Ȑ�ѐ���!cvGN>�c&�V��8f!k9�}�n������~�Hۜn��d0W��p�1�;��1+s�<��R�)�j!c����B�H`��S+
���r�F�)
�ξIL0%�#52.�V%���k_�,Z@$!%6�4C!Ht��]'�\���fw���roI
�7�z�O��&�������R����.���dɈh�B��@�+1�w�y�ԥp�6�g��xS!x��1����Z��9�0�)*P�(���Bu�7�˹$�I$� ?h|  �      ��8  �c�l                         � �                            6�     	    �` 8l       �� �   m�      �` mp �	��ъ�l�!d1;�Z줦�p�6�L��f��l ��ۖٖ�����c4I��� p/ ��R�ԪqUM�D�?w�|�I�'ᏔSeg�N&�޸�sS��=j��;[Q�U�����:�;�獶YV�
��eWgc����M^�^�������p��f��.Uv�P�Z�v��I$���@T�	�Z�1���i9.$�z���f�I�ID�igG]4�n��9:Hc���[�$�ؓ�(O�O2�*9j�GO.(*����U�^�YUoY��>�W��2�n[o<����E����`��	M7H�<�zY�YzgPl�U��� հ �����ݣ��Zm�����`��s����{��`��8G�U��m��$�i��հ�  ڶ8���m���l ��ymH	l�l��` Xg;m�f�ݶݶ@��T��?���4�ZT&��ک�p[ �1@m  ���m��*�k�ؠl���Ѥ��-�  �� m��&q�"M�C�E� �J�mJ��AKTmU�[A���i� 6Z��� 	 ��[@m� 6�ջcv�&�<���UUS� �Z�>�'O���b��� ��amp��m��$ ���Z�� �6�˹�I��p m  $��qmu�[m�%�`�P
l*à��,��[J�]U*��vb�rĥԨ
�Jܳ:.��d�v��<��j��U]��`��͹m�V�u�n���U�6*�&9v����
wOd�i᫪�e�݊��m	lR��nJFu��r�)x���'mp-�$��&6��'e�T��W�1v:T��30@��/E�H\	��U�,ln�� a)WTŮL�m�N�j�UW��Kk���˰��5MK9�y0T��
38��1Ơ��*��L�s�'k'V$�q�Tle��]���+���D��v
8�`���t˱�� *�s���*KGn��8T�UUvOD���$f�m[�Z�Զ��ӡ��Yv]��VӚYwm�Gݦč���@n��F��`�d&\�{�U��3W��u9�����������[�W��q�A�~�|�'MR�ͤm�֛�kiL��K.�*�J8G:Ȇ^�
Y�]8�.1l�V�9<ث�4�n���y��T¼�[[u[t�v�#�n������zF���$�E-��iY:8 �n���Z��	�*�R�@P��W �[M���n�mUS��l��G��љ�����ʲr���t�6�m��H �5uJ�]SH���VE�f�4�kh�e�S�p�ee]����5U�8�y檺�N������[Pm&հv� �� $�t�  a�mK%�e�kv�m�i�� Hf� sv��8[F՛T����l��� �k�ԭ�훖� A�-�ŵUUYv R@G%�5���$0HI:`���l-�m$ҍE8Kl���m1��{5v"Jܺқu{&�R\OU��h��q�՘�(�l[85�B���̹ԹN��I���;T���@Uu�mg�n`�m�m�n�I�� J�J�mN���M"�ppI $�e��D��$5�HkX䱣:�p �i�e����ҼUUE�) �e�-� �I�H�.�  6�6�gauu�WU*���¦dԁ��l�{`6����m�[�� ��  ll�����2�1u�d�f�
�Ysl�I�l�L $�N-�1R�; �UHMT�NVV�-��l��m��!����8   ��4���p �i˒Se�� 6���ە(��]٫���A�  ������}�� �.�UU*�z�c��jv�l�I#j݀J�k���[(�vf�e��R����OPQ3�.�sl�h p��RޣŦNkq�.�[[- ݻ'*B@H�j�IY��05�ҙ*�8�b)؝$�
���aZ:���%X�Ɗ��5��Ӷ�쯞�4;-[Kj[���	;�ph�#�C/= c����q(�M\77N]k3��al�mb�{�-�lA�8]���!=F���^��
��d�n��a��HM]�`ت�V���β�mt��BI��U��ݱ��� $ٵ�X�^�j�v��^��v�x� F�$ [I�9�<�h�P�� �e2T��BCS�B���UW�P����U��[UԼ�-r�*K^�j�5���l�NSm����U������@n��6Ͷ۳�Im�Pv������T�X)UV[v̫UR�q5Eqr�T��hV�l�j��y��5�%�׹{�P sn���[Bt$d	6�b@�&ܶۆ��[F۷�l	e��@�ZM�ؑ�E�6��r���Qs հ�m�A�.�5[��Æ�bڪ�`��
��)eUZ�`�%Z�6֠R��#N�2�K������S�p�I���UYW�uJkt�Ϩ��sk�V�Sj�*@�M%�ڶq��($��K���4���>7��7M��Ƶ�ں��xN�k���mր�m��H5T R�:ۡ�R�p�dଝCl]h���EM� �ۖ��i��A��+��2@T��j�l�L��"� <�6�r�l�ee@���35��Kg @l:Uu���[J�ҽ�m���o�P l�o-Z�	�,��e�l�*�p�j��l*�[-[���\��a,� --��	6�@��t�A� {lհ m$��ki�mmĒ6�||	 $m���6�h $ M����߾��UUU]R�������f�p[Kh 8 �t�im�ְ���m��k�  d����A̩H!���h
��%#�ڕ�ب
�;5T��[��� ��R��vz��`6���m[p�nkn iͻc��dU����!�<���$Ct�-B�5lu���j�� ���K]�]�ޯ��-�6��� �@�]$�&&�m[ ���KCm���H�[r�$ ��Z)�m  -�m�m�S[pH�|!# �`�t�l�  �� l���0Sv�n��R�jg��]��������ƽM��}����K>�ﭮ���l/Hк�s֠m����2�`��M� $r@�7M��:۶�C�]1})���nh��H��)EUZ�+Uu*� �P 6�M�l  om6�5�nm���[$K%i�$��Ā6�Q"��@R�yw`s5J��\���� hT�  		�����sd�ͧg�f��\�n�s���2�d��*nJ�#��UA���y����^l]6�Xa�Ė���9��ն@6�Hnͳ��[t�m���-����n [Z� e��m�m�  �-���V�ڛ]  z�mm� [E� E�A� m� lHΚ(p l�h��mmD�0UUm�(5YF� kX��Ό��U�tN�̫T��jj�����jV\�ؕ]�
�F�������k�l���}����B�����I.Mr�� $��^ĳ
{�H��(
�`�n�T�@6�nUT���R� ��a� [@ -�����v 6��	8 �n�մ ګ` l�p�� �� �   ���q  k[: �;l   $ m�6Z� 	4[j@ l�h�!���J�]eeiV�A&�P�� �  6Z  ��l�P�,�l�m��kh �h��$-���h� �n� ����a���ְm�    �ņ GPm�e��$    V�1����mm�� 6�8,�n�El  �;ZŴl�>6� �T�C[oV8 �a�m�mp		8H��
�x��;���|'���S��-U�u [j�Q0�Um3����0C�r9�D�����SP��:6�L�d�V��������Rݕ� �K�-@c
�� -ڪ���.���`�P*�Ren�X����#*�U+�5A�j�sE�lPEJ��s[v6� 0�bMk۶�ֵ���gm�$ �`My@�6�m� �Hu��@�����KUUT��H[[l ,�d� l  ��   [~�}�۲ݲ�amsv�4��[p �;!T��
��W�`kiV�x)R0� �U*䊪�� �T��$+dn�%(��U���������D�� !���pl�� m�k4��q�UTU4��)��ؘPȘ (�C������#� B 0�B
�)��BE�E*=/���
9T��\:���L��
��a�0"Ax�'�hQ2"�X&C*��"4-v�F�A��_� � �p��E�	�N��ρB!H���VB Ȩ�	"�(7R0�Mg��i�(��8@��"���H1F) ����'M��^*���D����d@����C�N���;Pڃ���~= �N��r����622L�L��ʆ u�:M��)�ht�AD"�!�0�.�  �pB�~"�@@4"��7��Ga�c�I� �(*@�D�.U0'`q~��D� ��"iQɀP�� ��uL��� &xl" ��@4�B(dr��� u�M5\+J
u�Qxq��P:'@\#����4�H@�A_�8�`W1>@p� �^�*��h��A��
��i@�՟"�u*��v��A����;D��>E"��@��(��B��P:�Q�p'$���H0� X�b���c	! � a� @�V��(1��X� t�ZN����U�|�\� �BHI@I� �D�!��X@�M Dt�8Q
��|��9Pl$PlPiB@�|!�Px�ndH#��*ȌD�D���h�M!�҇X���u��`ҺWj�j�t��D��J	�qCb�|��@DUx�� !֤���D!Z�!,Q�po��x��������W�^����jkp  h��ۀ    b�&�' �hPcg6��8.v9`6�/] p��S5۰�k��@5{	]�mў�=��f:����yռGGYU�,ͻt��j�d��F�NFs<u�΄�@����p%��:�E+M���X^I�N����5X/@ږ�K�V�I�2���p�8��b���u͕�<s�z�#��A�����0��� T�l�B���l묓�Nڱa+{=n�^pm�'�N��up��̓�)�9��چ^�K�c)�]�-�lr��tMt+�^�b�е�ä�6�5�8�8-����{31�<Z�n'(�'[���3\��^�#	Uሑ�K�D8��6���Ӌ�q���Ҁ�;m6��;/� J�&�x�pJ��+�v*�9,�1��t�ޞ���f�bۇ&��
�N���9�n�����t9��<$Y����m4�=��m����VzZ;\g��f�ތ��ME�#gӳ��9����Ӟtٗ6�98�9���
ܰse��$s�����1��n�H�{/2E5�T�u�"pH�\�2���V�Q�c&�/;&��[��;���&�\�SLΆDZ��l���m�H���bn�X���ŝڃ�o]%Nn��.��S� �n�����M�� 0Q�e�ڝ.wVe�����i�V4��.:��k�qi�[ ����6&7R3jy��pװ�Ju��I��f4s��sUT�bt�	yl�k�6�Pɋ����&�63�8i:8�n�7V�g���r�r��]��\�-͛.6�lVl61�VX��ubTt�P��E&�N�e�i�X���V�q5үRʋ� �;�l�uR�B���@RڲjY+F�� .��Ͱ����FښU8"6�s�KVc�P@t�9��S����7[O݆�T��m��
�ƥ���Pm��綍���MKΒ�]�p�y��\����ڬ�7�՜\���:  ��'�@��(i2*4���A�@>�e]��H��T�rtx�4'ɶ �Tb�^K�c̙3��9�L��v�
�������p8�G�_7[6|�Fp�6@��g��k�Ů���k��6���:˶�@�ŬYg���p�S�Nu��c�yQ��y\Z�6��M�;[{tv�}˨:z���'�Y��v:�M[]�A۶�g��9��ѓ�e��!�N;<��wE ��:x�Iփ�D�"�lNi����+��q��z{���~w��������.䅗���1,f'ls�	÷n7��|n�&ᤇN�E&�t m�Rr^�vW|�]�y��U|�}�u`w��F�Ca	��`uw1��9I�+]��n�X,�v�c>(�
(���]�-��#�����K`{�e��uw�X���1��#�����c��.�̖q��MrHS��U��d�������Ύ�}�eN��sІB�V�:���\�eEN����N�:sۧ��km��2=��*�I	�_��������Ύ��K`{�X;R�q���Ԓ���f;��s�d���}d��d��O_�J���Ƞ��,��^�1D�hrR�v}캰:���Ԏ��<�[����
���+�fb32��K`jޖ�յ%�g����3p���h�F�q����=[j���GL[%�>����������I�n�=A� ��K˞b�(�)���d9��r[z�6�m<Bk	i^_�;�ﱁ��V�l[�������*n�ctS�����VWs���c���%�9T��^�MrH0�1*���ؠ<���<ɛ̆d�f�H�bH�iU"� ��32�M/D�̚יJ��ֱ��D�̫X��-��z[ ݩ1���������V
Ԥ�n))��q�{Rc�#�������>��[t}���K�#������ϭ 	���>)���kqv!kwZ�1^볹�	L�qU��?��05l��ս-��jK`o��Te<I:8���U�������)#�ٮ���n���]X�a��P�I#q��̖Wk1ٵWʦ���V,�vq����EMI��$�<�Y�@z�)PfE�|ɓ�gI2P����4�3ZI/;���{#��|$���.赕yl�K`�1����v�U�TY�'J�`H�6E�î:�tN8k�d�Xx�ݖ���h�u�~��.��5�5 �N�#��1f���,��cߐ{3n�*=��4��Eyke�t��յ%�7�:`j���L��IH�NShjI`uv�����V�l�&0
��Yk.�����I4^f�P���I�[R[�B+?(G嗔�fS��Ƞ5�ٻ?okv(]�*ē����A�AH	O��_�k$UWG.�R�S7,M�%����Ԝ)�����E�X�.�:ۇ�i����0�t�u���gų�)���F�7=[]�-A�=��?zMGi��&N��=���n�Q�4�c�5�����Ѕ����M=7-la���	ɉ�2��8H�8�J�.^L���;�7/n�ۅ��ݳ �Wn5(�jݮv\��`�70E���M�+����ww)o��7"�US�u���!=���/
-�=c-�m�l�{>K�oI��t�\l�L�Y� z}�05mIl{�w�߫�9tv��fc5�m�9%����v}�t�ղ[ �I�w`���0���.赕yl�K`�1��a.����mrH0�H�X~�,~�v�ݚ ��ɠ���]�ʀ�E��v��Qƛ�9�}��`uwv}�@[�2(d��ރ2 i*A��L��ṈcF�㳰T�3<�s]�7h�b���#R�q��JmI> ���`w�˫˹�j����,��-J5,�s1nLg:�}�wF��|)��<!� U g�Q�@6r�\}�(�ܚ ��dԤ̓�y�8��P�/)f^]%��1�nԘ�ݙ���f�6��n;�9�K�ݖ��u��L,��;��c��Q1(	�$�:�Y��ھr����M)���&0;J��"��E�����Y����O)��M�Ϯ0{.�x�-�ҏМ6�7R1���;ܘX]�lvL`jڒ���v�`^`�WXZ��K`�c�jK`ñ����7tH�M���;��`{�f��%@��*Р�aU��}(�jh ��u�MI9}��RO�3jRUq�M��%��?V+�Ƀ�IlvL`mpU�bYv��.��b`ñ�IlvL`wv01{����6)Q(�r�D�����br<�Y�C�nN9�ɵi����wRcu���o,���xxRK`�c�����3�3�ȣb�1B'�w����#<��`{�4�:���R3Y�h���JnTr;<��`w�0�:����̖��I
N�ct(���5%{��>�E��dPy*��̓+I2X�&M��5�1�̈u""d@'Pi������\^����we�����Ş�$G��("��:�l/X�9w5�S׷:�ێO��v��ܺ��i����{�,�����ra`y{����"�IP�JmI,�������{f���vWs�x�x)��Q�9��{�����ղ[Ȓc�B+?(G嗔�/.�l[%�<�&07fA��f"��CaD�:����7v~�gJ��"�����&��j�_�Y"���8��ZMi�(L�9R��/ib��V�b^����'�[�֮m�m�&��餳�y]�W�͓]�������9���a��@�&���K!cLTۨۮylw����pW�>p��=�lNm�Л����Xz�H��K�^vs׮���|p&z��2���.��;bݎK��˱��s��D��`���������1��6�c2`���&� ��h��������[��C�SA 񲹻�M�o\q��7]�K�F9}�6K�:�՗�l������09wK`j�-�m�7R1�"��ｗV�t���L"I�-$�U�Z�,�9V�����_�Y�����ݖ}�u`yQ짔�D܍D8G#�;��D�j$�cI%��/�I).!�˳\!U���߿�������?��I)r}~�IN��I$��Y3^��'� ��=]1�u#��x筱�ݍ���ݲoD����: ������ ��ƒIwt�y$�F�����W��[f�ϾI#؄T�ДqG(��ZI%�{���y�*��9���kPi$����I��Iv����J���2�W��$���4�^�I��I��I/{�>�$�̕�"pk0I/Y$�y$��i$�wL��J{.��I{�V�o)�������I)���I.��$�鎆�K�I3�H>������l.�B�s�;=,�8�m�.q+���q��+�Үű�į[�Z��]��I$��g��S�0i$�d̟|�F{.�����O)������}�Ig��/x�K�����$nmԴ�K��O�ڪ�6���X�6'$�5$�ն߱=�g{���wFuoD�b��P��kK�	��z�*��g��N�H^k d"�Y��q8��D#���8p�H�&E�N�+\`@8'\�^'�X)%��g��&�v;"��*�6k�eX�#�����A�H|g_�0�����}	����	$b�t���"�S�چ=�2FJ8��>GB�I�K!	���e�t���3���$ ��:X����r�p�H�apу��<C�fC�|�A��>S3��>8��c(�������U����A�O����Dc+��x�=��)�3c�x�({*��4�MiB��E: ��#�gTJ��4�	���(A�CX>������"a��7��y�g{I-͗E�m%����%MJ�!I>�%ڦ�7ꖒIffͮ���6]���ޙ�;�~����q�,��P�bV�z���$�Y��﷕M��6����)��n���76�mW>m%��?&�Ri��)�4�9v�:��(;mq���m�Vn�{=F.ƺL�4�e�t�k������O�����v
f{���[l�}�?��1�1�]����w�2J;d�ȗ�S �DD�)�����wg�2e�$�e�ޥ4��J"wz~���r6��_rf��}�zw���B�ctO�Iy���ꖒInfϾI,�˥i$��fO�I.�,m�Ԃh���cI$�t�y$�\t�I%�I��I��\@J�E(K���
ڔ�P���jL8�q@M����{�:�ծ���n&�$�Ȝ��K<��ZI-�Ds�{}m������m�9�j�n�X;�v�:˦=��n�\����r�['"6�'v��)�s���]�>Y�nҚӗ%���6R�I/��}�{�$N����S�g��S�.���^;^
mc	jTQ%$��θ�4�JwL~BS�:M$��)3�I#�B*qe��r�rR��K=�|�Y�&�K���$�뎓I%7��I*2�2�X�3�I)�&�K���$�뎓I$�t�y$�Y�(ŔaYWw���M$��)3�I/���ϽK�$��{;ݶ��m�9:��� �����ꪪ�g{4��T��V�M���5��=l3K��뵌(�T�t/!o]�l�^��S��nM���7,u�݈�ՖļZ�5��WϘ^�`x�;c��;j�m�]��<�D�����ZSF�;u�m�#Z�k=fݣ��[�^LZ8�	�B@���ŘGn�n�s�����u(�%�C�ʞ�\�������޹w@�]|��gc��nf���|�{���������|����1\6�a���«�.�����IG�m�«�VG>4�v�S"Ph�-$��I/y�Ҵ�K=�|�Y�E����̟|�]lX۬(r�n��R��JwL��Ju�I����&{�%:�bIc��O�tHIMHܓ�K=2�N���c�M|��~L�lu'�ww~����w|ǈ�1��NIHj9)X��}��g�$��>hi$���$��G���I(uM��d�Ѫ�� ��߿� �{ܓ.���ww힧)����3'����1����d�������\yzu�>�B��7kM��op]l� 5�}? ۯ|�]����~[m��}���{��Rj�n�����~=������I~�~K�%D���9���{��RkO�P�)!�* d
�_��s��7�m�s�[�m��w���{���w�����ݢ����l��̞~��ww˜�)ߒ�}����w~ުI%���i�9Ct8ڏ�K=2��I.�3�I)Ѱi$�r)~�Iwfcmr���6�q�I{���K=�����ȥ��%;#CI%�������R��z�+�e����Kx}�s���7t9����k�����!+Z�)j�K��`�In�R�䒝����]�g�I,Ɉ�1��9%!�$I%��2�䒝����]�g��S�`�I.7���Ɠi�Q%�$�ze��I/w���`B�<P,0`&10,\Uht^*oW]ֵ&����rw�I-�~�Ҭ�)e�f^bI%�&{�%:6$%�I��IN��4�Sj5�%C�
TpNO�I,�K��Io+���ޤ��ۥbI/{�>�	mr��o$���̊���nс�M�\�vx��CqTw�r����m`.�{N�t���$�ߏ��y$�\t�I%;�{�Jtn��K���4�2��CtO�I,�ˤ���ݤ�����K���i$��&{�U~�mnɭ5U*:#6�r���[���K�simW9M������%�{t�$���x�Q�!%5#rO�Imr��^�Ҷߏ{����c�.��`�}e�PK���+pT]�L��-d͗wy�������Q0D�!v���I%�g��_~��3�R�I%&l����ZI/�\��7X
�R�t��I�OFY�t�j�kn?�k����]�	��1�ۑ1����[�;��K�\U������J�I/{�>�$��0[ʯ�I.��ϾI#5*\��d��r�r"�I/{�>���̙�e�fyޝ���wt�󻿮r��fJ"�V޵$IP邕��K�&�i;���2~���$�3�=NS�������[�h��}t���}�r����������ն��s�����{�n���6�i��#�7A)9>�$�開I'��ӻ�7n���T��������wwI��P�DX�$�
1�{�_�Ӣ��:[k9+�k���T=�h*0=�H�rh:y���g-�1��'kn�j�$t�6ݬ��HƯ`���ZRYS���神x0�m��g0Y[W]���d�c+��t����H��[�8���6�az�S��W:�Y�%t,�׮�+�X=�ۮ��v���&�eZ�mܮ��Ϋ�`�ۍ�<N;X���Wg���[�2L��)K1sL�g*uS�r�����ӻ]V�����i�\�V�ێ�n��OnB8���f��>q�;��@�q�bI%�o����V�fd�W��Xg���5Q���M(ے)M�ܒ���Ǯd�.L�@Z��3�����oyI�ilm6n@mF�V����޹ ���0
�x*˗�$%*"R�X~�){&���`w�1X~�%���`ԐVsi��JJrH���Ky웫�����=����m��F�[e+;-��6�΃�''ck��uQ�n�$���vB�gt}�P�v�^
�<��ɀz�����@I>��D��Jp��Tn$�V�fd���	 �rrG��0|�)�:ҁ�W������I;��:�}�w�������oh#�7A)9,Ǻ�wy4jfd�{�� {M٠2�V6UJL#6�qXmW*��͖�f����k����M�`j�[OTJ6䑍�ܒ��a`o+�����c�V��K:<aK	Q$�tQ$Ƹn�myy���⧟na��M��Fݰl��}�{O�Wۢ(��q���,��+ �{&�s�͚Xa�
c�HJA�\����\�7%��@f��@a엩�$��d�����+ �w�ԓ��{5(�� �,EN0���\h�X�1B��|	7]���hdv�~Y93.�PpnK�����;[�,�����͖{ ��Jp��A�����=����f}����07� ��:�@�'+��8v��-�]ֹy`��\�\x�we��-��U��{����~[e�/mp��;�uX��|��k�������l��r�F0n8�w�/��W3^�V���K�<�{ČU�M�Fܒ1��Xǚ����gꪮ~�7��+ ���Xǔ�1�DQ��ӏA�;���hdn� _�&�ҥ�;)�$��b��W��S�W�'k�����`�߂��8�BR�$jK�Ǡ9�&����������h����3kg=�W
;�c��7`���gFyy}m.��ۃ��E=����l}�� m׾s��<ʉ���/vh\^= }�|�\�M����7+g椉*:� ܖn/��$�2��~��;��3ٓZ��s����Am�(��A���Xwf���1��fd̝ͽ٠/#5�z��2 x�D ������ɛ�2L�{]�@��@z���9�e��ɢ/��hΔ���� "&&%�=�4&e�̛6�����4��@R�fX���a@"F
��W���� uB�B8Ӭ#�"���km!,#0���g��p`s\4cb?|b�]�/јd������"B���.��C�)�_�!�.�)(� �ŧ�p� �Вd�@��\@"�D�"����S�Ջ��)���y�2���.WO8�X@�*F!�G� I#�v�P�iØ< э$Δ�q�)�:rhQ����)Pˁ� ,dH�p��R�>�t��`O�I6i��>�\�/�ލ�"�$P6�L.��J���.Mv������8�C�a	�7۷Ozv{�}���  ]6��   ��kn�`    E -��m�$�6Z�+��%v�������6%�-�B�(G��\��\�.���ͧ��&��`�\��am�����lǕ�\�n��7[���������o���c7��ԭd�H��Pp++��V��@;�&�q�����=�۞g�keh.L\�kPY��\�Y���]-�P]&�fu�%!�=�Fq�+�[�m	n|t�gvζH�lqɮ1�<v:x-��,�^�lj(-;[k6���7g��Σ����s��$��t�୬g��<�ٸrΓ"�l���i!,�[@�F"�۰��T��x,�n����c;6mȫ�t��ݢ���\9�3���ts!�������æ�6��nX�<`�(G�oHe�z��ݨs�ԕ�%���/;N�!.+K���9�*�\��]�����_�l���e�e��wH���&�j��4wJ�:�r��d��(W/a��*;�����Z ���vʦ�<�u�T�[N�X���v��gm��ݻ#�Y�t=n�RcT�">�re*9�k[b"[X��sЌ[@2��rF�Pn����+9ٝϧ�4m��Wt��W%G*8��+l���&:�+ٌ7m��-p���2]�����B�Kl�K�o�m�E�PR�rnU(����ưR�#�F1a�h՛mc�m���Nҭ6��A�u)�k�<�����:���p�&���B�S�ݹ�pӀ*���ݙ�ɛkk[���'v�ӌ�]�R�aL;26E�x���Vi�<���-T[@�
յ� �*+e���s�*�ÓV�����:(��!�C�#s�"g���8�͚�+�m�<\�8�Ö��U���ත�u��Ͷ�rmYmJ9ѶR�eZ�˲�ld�Ř�f���s[)�t�g8 ��b�5\��۝��3�93w+���f��WX�M�� %�@cC�B������d�&�%Π�^8Y*^��'V�ѩ.q��6˜�8�@���aGJpp��~C�
��*@>詔z�N�p��B
p�E�S��� �5!�{�3�*������H.E��i�s���]�1WR��	[iQ9+�,�[j�/f���eM���`Ӟu�(�nK���RK��|l=��%�V.,p;���r�G����+`*�U�a]S�䛒Lx�[Om����*�[<�um�G��{}�|X��[�#���j��c,�f����Y[`9��zeF.1���hyb���.l11f� ���
5��\n�7h��8�֩:�� ��.㒮�:����n�r��769獾w{|��ݧ��-4�������h�������ݚu�-�MҊ9�#���%�?q4A{�����@|�y�$��ix	�dBBR�$jK��K{��s�o��@��4�wpXؠ�'y�$̔̙�76(>f� }x�4̙��zX�ɲ9"T:t)R8����@k&fO�7g�=�:P|������K����q�79��g�.�e��m��.�n�7F9v����w�>v�wFz�������vh��(>^Gs3$�o��@s�9�2��D��`��.�=��RL��Ej�a"& 4P���A��0mB�" 7&�҆S�.�9~���'���<��"��3&Qn�w�i�L��@[�tP>fE�d�oxlP�4�<�����'C�!H)"�ڪ���ؠ-�5※��2eɚ3k��״�F&�E�ڂ��]����I>�x��Ɂ�$�:U�1�"��ӹ:�:j˸�����>���<[���^�n�t���*�2�$% ��ff�P\f=��ds&eɽ��z(9��sr�P��Z&%Pz3��;�}݊�٩���������ɲ7 �t�<�1/@y�v(?�(�u)&BI�䷜㼼۫��U���X��j�:�n^f&(92fK�FNo<P�Ԩ\f=�x�7TW�44��T�Jr����������殺5oEl	%g��IN�zk��ɓWGۋ�إ�=$���n�,�\�nC���m���.���t�e�e���Ɂ�$�����^A�[fSz�$Br��X,�w�UI^�N�ř����c��U${)�lB��Q�M�)���5������s�uf�:�u�x�F$% �*LPrK�&h���-�(�3"����>��~��`BB0�(@��T�_~5�jI=��!���2�1*����2�L�\�txY[���������8��JQ�8Kb�{[�kn�9w�\�;y8ݺ+7b��� vﾮr�ʒ�nAP�Ф%F����v���(��Z̙�p���P{/�*K��H�y���<�W�]�ɔA��J���ߝ����{U\��^��b�QR��)��۫���f��K|�U���5���%������ʰ��qu��;�uX]��k�K37�:��7��rD'R;�y���\�����]wz���dP&P�|:t$�#T�EfG��1�379�s��JY�t��mW�ʫ��Rj�k m:6��9!�j�xN���pY��BR�$U�s&=td�"j�Ѳf���gr��'4���n��]��d���0��y]V�u�[csD��NΞ��u�l��ε��i���Q��yIpK������lµv;S��2t�O;�Yr�n�m�#����.���-����=��۳��,]	��������t���d��6bܘ����ujq���=����C[�����o��~2Wn�n�-����:��\�h�� ��m�����wyJ���2?W/@_Gs��4s̐HJA	ʎ����W�#�7]��{�@y��Es3;�뻆���;̴LJ`��0"�-�URQ}+�`}'Θ��\��*:���,7���ۮ���5��eՆ�RY������Hq���H�����-��E�3%̻w��������,{��IQE|jA���8v�qЪ�u���GRQ��np�Nz�Nx��X2��������	J������;��`{2o�1z�]���KW Ӫ���1�RI�y��1� }��'���+nh{�b���R�fd̹D�u7��6��G%�{~��p�f�/fmՀf�����X�6�9)�S13A��"�ؠ/3iP���rK���� \g�y���w�y�x�=w0?�O��<�ﱁ%� ��*���tOV.P7nJ��\t�-v��z9#{[�M��oqsؐ���mm�9�n
�k� 7wf�.�&�̋��$���:P�͹�T:tӕnK �ْ�W*��rd�wF��n���5�ə's�{�"JiF:�nF������{=��-��5Q���	 "D�TI:}�:��fI���ߦ�.�f���D;�DL��w��y�b�Y$�'��Ҁ=��@^d�r����9�E�;�4�:&&J �3&��Lɟٻ?�xlP����nT��m'N��4���qK{.�B�)�\�n5����w@q����ͺ��{fG��T��7 '!$� w7e����{���U|�����[6�Q��M�M���`yw�;��)#3&��ݖ�fMrL��� ���.�;̎�����<P��4k$�{wf�=f���H�RRS$���{۲�;��RI��{�I�(J.T8!�W÷��,�n܉�*:iʎ7%�}��@x̚��
 ��M�$�����[�V�Gb�� <\�q��˳g�q���om���^l�����Ԅ��)S�úh��(�y;��ݚ �֓��H�R���)�`{ޘ^��٠n��ֳ&���7(��w�\'xv��N�fd����2h乒�/k��`n��X��̊����9$��%�ݖܭ�`{ޘX}�s&Sj1S���R9,�Vd�7�������@fd��L ЭY�DF[]UU��ݪ��A�\�GC[��ݸ�iӓ�Ҹ���m���+��M`@���K��jL�݄����;!!��[�X:��H�+f�^Y;hv�v�0vG���y���qƚ�ۈs�\`�ֵt70�lvKo�>;g�ǐ�א�.�B%]��嗳ǯV��k�5ڼ.�l�km��mq�/X�.ѓ�a��i�2͞�C�B��6Y���p�B��E�O"̓����.r#Oج�O�[�<�3�W��$��׵�]�%��qv���y�lo�iW�����<P��h�̝K�ڳe�i�4J��(���I �}���wvXv�e��za�RF�M�ӐT:tӕrK ��� Ξ�g��Y�4��l�;�AeDFیm�Ԓ�Y���٠32t����re��/��+ ���I�j���)JR���酁�$�����vh�Y�@^1T����vi��
�n�ɡ]q��d�m��1��.��f.�s��v��C�s�V��z�&�>�ɠ�fN�3|ᙓ� n���Sn����I,�̗�+��WP��x�2U��P�\J'A _�ܛѿgP;�4���/k���H���mF*q7$"L�� {�����ɓ733&hfn���߿K ��a$�6% ��������h�̚I�&N�f�5j��N��5$���,fL���wg��vh��hX`�\�4��[��nv#y�ҋ�b�McM�m�h�<����[����������q�瑕133? {wf�/�d����.d̕u���������"������%�_�ɠ�ɠ]��ٙ5̹�$��w�M�L�)JPҔ�7w�Հ}�w:�>��ۙ��-���A�&�	�&`@"�������"���4&����"D�	�d��^�8� ��dFHH@�2S\*pHB�"�5`��� � ���3%�	��Y����>"I�ڐ�	�$���Gn���@�� �OE���B�ۇa��2���7�ڃx=S$N�dG�̀3bc=M&A��8�W�H |��2qX^��E��qQ���Q�P٭��h��立��RCr�e���<�\�!�N��U��*�.��`��c �T�����IJ�x��I�@M�I`fd�6�\]�ݟ��ͥ@�ɠ92J�J��J�wCa�w��j�Ap����%��O>��m��k0���ܻ��ݪ��Ne���k��׫�h��T뼞f�/@��@���G�IM)U$�=�eՀw�ɠ�2h�fMjI�w5��k�S��y�PLʠ�٠�2h��̙$�<��~v����3�e��b�Ӧ��䙚L�2w����Ż��*d�m"16�s�c�Τ�����rD�R��7$�>^��`o9U\��߫��٠�2hI��5o�'�����R�t�Si�ƳV4!H�6�=�;.p��k��U�{���|�|A���Ƹ�8������R�]��ٙ:�ɒ_8y�n��hX��Q��H�X}��fJ絙��*��ə�7S�x�O�96I%�w7e���f;7�������V�͖s&Sj12���IA�����s��(��T뼚 �3&�30i�9#M�H*R�v�캰9rL������>{Y�@rCd��b�F @�� �`&"�	D���>3�Oc�2fb�7[ͭ�6��]Y��n����7N�Z��%׬P����,�F�"��qfn��Lݹ:���ab�g�(#�����,��g���6�u�K��y��=��<y�sO]������9e����ӳ����<fV�։f�q�<G!1���L�N+����ɘܦ�ۭ���m�n�ѻd����~�o�����Id���M�qeq)f-���?!�"�Ԛ�>�̶s�m`Q�Z�[F� �|�BAL��-��`���`d����w��n��8׷s��� ����zI�]]-����ef[�Ɛ:m')9$��{%�Ur�-�f���J�>�ɭfd�e䏩�<�x�yQ134�,ؠ/ה��L��$��t�����p>K���"%w��lގ��L`�1��_��\��`wIe*Ғ��ur��fJY�nl���f��^R�1�����/6;z��5�F���uM�jz��Y��+����<q��p����ꯛm���@��4�2�����6hܝM��d�i�#��=]̖�>UW�AG�JP��_���{�jI>�����Xfs��Ĥ��X�:`�1�W�H����}��
�VR'
Q�r9V��*��� =����G�W���X�ͷ� t�^ay���7d�i2�0�d�>�q"� �@�DS��ϔ��'�M�o\q��ș���M���?,|����R�q5$��K�̺���7��6Xs�*��:�D'ݑ� ��gL`ul�0=��]K�	6�:�IV��K �{%����V(�"�b� �Yaj�A�R���G�ʉ����7��jI�n�X��bx��I�JD�Xs�,Wra`{��V\Kۛ,״�6� ܂m#���w&�W3ۿW���`�d����RR�� ���3��΂���]v���[Źݍ��I���LϷ$�2���ؔ��I�̺��X��y�.I�zVt�@s��'%���f%P��kY3$���@b��X�eՁ�e��j�:m9Q�$�e������$��^�* �͚�d��T�)�e�&f���nI�h՝��u* �^M;(_&I��$�9U�<�K �ōBF�:�JI�fR�533'�͟�/sf���(��������YJ9u��ڻ�G�"�m����ݹ��J�t�$������{�ǉ�|���t�5%|�͖��K�ܘ~�s��۫ ͥZޔۤ�%$�I,�y5��̚ ՝<P�Ԩ�y5ɛ��7����;�$D��)���5gO�0�1�M�HZ�/2�"&""G�L�AܔvoyPv��z�h9&K�Vw�P��9���a<Ĩ��T켚�?�6~��@_�)Q&�0��J�z�h��D0�Š%
�s�;�1�ə��UV��֡-NTF�^�����&�錜M���Z�(�t��ݦed��Q�J^1sǗ��s��n�ލ�6���^���'OH�D�s�OL�1�c!���p�5�^��;@@�TZU6^��	k����5��\�=���z���Ĝ��t����8�ڭ��zl>�u�lŷ=��e򛱱@�a���'�e/��0.���'b��t�m.��׻���Ϛ߇'��zN�i�D���;n�^C�v��������Z�+�s�91;9����]��(�M��9������w&�캰�X�X�J��n19���-{'
�L�(�sz� v�M }��� ���'t�r��,�m� ��Ӧ0&� ��R�U)TQ���jJ�Գ3e�wse��2aa�ɓ2����Tܝ?G	��)��Y��=:cҦA���� �������
�D�nS)2#�����'Y��m�<��r;��|v���H����������q�:�M��$������캰{�?�d̗$��������1//S&s��'>�tk��Հߓ&������h�d�Zəܷ�A���N���r�ٛ,��K�VL,w�u`gJ3-��E*m7)���U%�͖r�i`{�˫ ｒ��{��R�m�'"�I`}�Ʌ���t�����`�1���Oٕ�^_������!ʜ�]a�k%kx�ۜ&��wv;h*�lp�IQ�D��I���}�V���L`zT�0;n����*ŖU��Z̦���L`zT�0;{.�1RǇt��BdNK �=��7ӹ��O$�@��BD0��� =���jI;��:�s�)b�L�r	�P��.�m�`g�n���K�����3ti�r8����U���������L`zVL,���ŊTdJ
B��R�6�[�c�%����s���n-6[����g؀�'l�5��yW�yL��0N�����`v�u`}�f[�LnSq�`g�_ꤎ�l���f�X���ؕ�ʔ�D<�/34زp�/ה���ɢ��,߷����'�SD��A����~T��4��A"L���
B��J!�D~~"e�*�Y?�	�K�y�B�0�*�.�&��2M}[��/�O��������Q��#�����۠��6컶���������Y�u��c2�����挬�y�K��2ގ��߫�y��,״�F&A�m�R+쬜+���MnoR���>ȼz�K�mkOaq6�T��3ٷVwy4s$�;�c5�j�Ҁ�۠��R'G*H�X~�RY�����`}���UT�ٿU�ݣv�N (7*�/1��}ҦA���� ��'B�d"5���!tn�H��$n~�GXs�Y[]}�kA	�S� }��i��h�S�`4�b�#�|$ҟt��]Q�����X����4S?&x��%�����tA#�)0�z�Bp'�N�98�X��΄���M!�t�5!�)�CQ�m�B���|dHM��Cg�� ls�0@�0�	��}d$7�!)�E(`2Y�07��Ā��� �+�lR_{'ϒ�32�ffd	
kp  h���      b��l�8@j����Z�rΒ��Fv�f�z�������XH��;�%�n�"����l�(�2��5p���ucZ�7r(8���'�ր��6�W6��y1��kU�z�!i��E6�-��`��Z��l*�J��F;k�`6���N�ۇV��m��zӹ^u.�Z���'pt�,����q�l�ڴq۔��d�+�O=;0���ݹ��ڈ[;p��ns�t������E��x��9�\Y۔� �]usrh��b��[s��7��5ӎ����#vt6�)M��b{c[���s�8�-�g�����N�;�K�U��$puI�j烞s�v�]�ᣱse�m�FzE�ҖR�⍹�X�.��mH�� H8��M�U@���fڡG� ]\��i6���]���#ud�ۥ�6�m��;2���:�9��z;p��9Z-��5�M�����A�i4������i��8���ѱ��nw���pNG��t�ë5US+<��m,�4��%U�g�U=�݈�,����\WM�g*\؎{Wv&��'7+�щ^�R�a-�MŶ��e��vz�K��JFC�۵��r�m�ēimc��^���2�\��4�Yҥ�����I�3=���#�gv�O;Mn��k9���2p�c��0����t�(S�����J�ق�kAUTt8Ye�@m"��b�p5������F��[1�i�P�������VL�r����6x��ٵP�w�;Q�ʌmeh��Y��\�v1pd�6u6Sf��$2����Ӊf�{v�vZ6췘�ȓ�Kokzt��k�ܲ�� [d�����٬��.��:��
Q{�l���v�m5�Ψ���)Vy4�[�Ez��M��>�����G��$�����9K���V��U.�-ۗ��H�R]�uu�sq�g9�fs�d�E4�h�c��"&@�]"9L"��#ҋ�~��8�6��N�� ��@v4>L+7��c��9�WHٴ�/S�«��v����(���4K�]3Ù%�
j���������̝\��ɺ��=X�]��$���4�t[��d�����
<\�"s�n�F�q�4:��;m���C%��a�ld.dM�b�n������甗��tia�n�sFy����4�^�9�Ŏ��ջ;�^ ���R*A���s���Yr�9�DGzc�׽�T�N9g5�F�\�mp<��ĸy���p���n�s��t\+ٰn�ڪqĬn@m��NF�� ��M(��* ���K�}�@����ʼ+�*є�oGL��0=/��>�Ʌ��$g�%����EN�F��$���0=*d�0	,xq7I�D&D����5X�٥���.���K��ڌT�q��f&�L��������0!����ߥ�D�8��t\�i��֐˜����$��׵��aɳw@@vD��r�2+�YX�ԩ�<��* ������M󇶶i`z�*�m"pBt�r���K���ުh�������I>���jI�{.��W;�� N�� �rX>φ�L�?�~K��� �}��������,?r��]�����f�X����]ͽ,������E�Jx����R�5�'�͟��l�@}�L,��ʶ:eEBnF�!'s�.���Jh���ܽl�/�<�nܘ���Ue*ŖU��Z̦���`zT�9��%���T�7�g�OL��.<L�^Nə&gsڶt�=y����K�U\��fM��b����M��}���ԓs�5:Z�U# �0�����0��7�l��@}y:P��#�D�DH�T̔ɓ$��(���`}��0=��`zT�0<�PJD����,�̼�����0=*dw�u`yw���*6�F�(�;1���E�����[���m���>���G���i��+�.�+//1���ҦA����~@ff�ٚ���	���H��`zT�0=�0����A�zu�xH�I��M���}�d�{�,�Iw�4�;��K ���tS�A13A�&w�͚ד��,�(-2� #�S �RQ�L`c�M�k3J�I4�oz�h}����Ay�W�W����A��S �=�1�{��`~��UVx���T�HI'���[�#���\��h�ۘm��h�6�;r�Ǖ�Tb����M��;��K ���`��Xw� �`�x�j7n
�I% }�ɭI&nQ��4��زp�>GJ�,�|�r�{%��}0�R���,�&��f[��������`{{ ����`{{ ���ff���V7Ni�)R!8Xed�@}�(��h�s�,�ɣ������N�^����lH�@��:#����j�;N� �˹�Q���1n�D�vx����p��Y�u΋kr[����a��ع�x7Z�-�`<� 2h��l�y	ą��ckY�����J����<�w�I�Q�k"���[<#�]�la�:ٸ��湴�-��a僶�^���k�q0�z4c��U+�N�.��5I��d�k�7���u��y�@[�g��w�����w_��~8����ΜNz+64��N���tm�i�&���n�YTẒJE��M�����a`��Xw��v�i`�-��QR�>F�`w�\ɒfw=y:Pճ���p�d�%��7�
"L��L4�������g~���� ;�cv���)4��	2�}�����l��=�d�>�W��7��ۍ�NT����A���ˤ�<�φ�VA���.����s�V�������\q�趷;���[�[ƹ;��M;u�������I>���z�
�Z�9�e���<P��W ����Xw�U��Q�	3*j��jp�.�p��y5��tA���pMQ���ڟ���A�{zc���jᘳeѕh2�ߖ�z}�odީ��wԖQU�dtS���,��%�޼�>׊t�>��\^�k���ݒ:5uP��}������k'�O]۝f��+��)�c�<m���nW���k�m����Pz��@}�92�����y��!�5N)@����}S���U$w�4�^l�z�
�eɚ ��QG<�#��2P�<P޼�9�C���i�`�(?�l���I2��O���:P9�bsLð�1%2d��y�@z�t�>��a`}�L,�� ���rh�s��̯1V���Ҁ>�ɠ;��\H���H��cJ#�����λo
���o\q���{-݇�\<���L(�1;\`��VA��� �I�~���>,ڒ�$R!���:�����L��wf����(]��Z�rh��q�	s�/	�(i���/{����8P�Q���
�*Յ���������I�yZP�����p��d!F��T�.�b<����9��o����6���q8���J�jp�7���~����@}�(̩ٔ)RuD�jRiӔʌl���k��u��s�X'����[x31�g�CϷ%˖#+*�����&0=����Uyz�i`���#T*%F�,��M��p�=�s���p�LɓrM_~U?D�tr�K��~V{Oج�T��&��n���%�����0LDĽ$�js^���נ��4���qw�uX�%�H�I���鸬z/��f\��|�w=�(�z	��~  b�� �E�AJ�1!0���n�o���>����G���;:`e�n)ֺ՝�,�g�U\�����F�oh�GY�9/3����g���i0Ol[@�kU�k�P��t�<�h�����f���"\�gv�r�9a�6�nx�d���2���'b8}���0��jznV��:�S���ی�s��u�����3�F�.�/[3�[������<OgG`���n,b�.$�VU����C�d�=��www�w�ߖ��9�D���H�Tq��]�Ã��'��ŸJ޻�[��+Ӎn��m��v�CWWW�,������܉��W�Uy��U�iZ�iM0c�$�nI`}ב07j�&��LoL~H�e�Y��D�1Ɓ���������g}����1X^�66d�m�*��V��LoL`{nD���K&��j+i��
�QI�g}����1Xj�L���"�i���Z�"�R8�%��'���$���N7n���xݞ�@-���)H�\J 'E�D���=�`gj�L�����J0�YV��0LDĽ�Qx�/&�$��!���E"T8U0�!τ����Ԛ�G��w6h��\��k探q(:jTC�"�=皬=�~�).��}[�V�OUb!)ӥO�f&;�0=�"`M��0�������{�X�k_�I�7"JFܒ���1Xɒf�[�/���נ{2hI%���]�z6Ͱ�n��U¶�-�>H��g#���k������1�������Լ�́2�����@{�x��fO�3/�=q��[����5n
R����j����;����e* �+1Ŕ�j�D����;��`}ט��8req��2k��v��� E��4"VFVA%V$b0�#�i �J%̦-qE4l�4 GX�#41���	.U a	 ���i6�*�1�E�0��+$Hز1�T;��0p�����*}�v���G8	��0�0$HX4��j�� ��s��i�b���$�# EѣK��$"0�Fʑ�HHM@¹J�-!F���X�@b0X�� "��B�����3���o~0�`a�Q��!�G�B8C'��#$"DbD��$��;�~P���I������}Ǿt	��/�)��"����4*,U��E@(�_�E>W�? '�T:�@��+5�*�]�8'�N��MC�3��6�u�)%�6EYq ��<LDL�oFeo=���P?�"�;��`f<mVBTCEJ������e*�32�� fwM�E��w'﫢&|��y�G.�a ���϶�i�y�۴
v�Q��v�;h������ML-����ݾ���R:`v��
�D%6
�$�v��K�U\��y�ޭ۫���� ҷҒ`�E���c��Ɂ�R:`yl��7s%���yR&4�Q�4H�5{ջ�<���fM�2I�0d��'t�G
DH�AS���T���u�/zՁ��Sc���i�9JJ�<�K`�cv�&�H��_����ӵ.K��ݮ�x�ո����z9�F���-����C�\���kF��v9.���O��`n�D�ݩ0<�K`l���!E'E
F�ܖz����=�ݺ�:����̗��I�[U���R�1/@]��T��ȣ��;�{�@_�j�<���q�:jTC��X~]~݊ �ݚދǠ�g�[�*-l�*���*t�q�{�,��{�5|�ݥ@|�̊$�+d� L!��P���F�L#D�yv���Y"���8դ�;�\��:�⦹k:��v5�8s�8]����H7nmm���8c���5���}cE��0���wlk�a}����p�\j�d�G��t#��u��;t.���΋��jm������nT��C��:���^z{6�\���e��Oc���.�Ur���F�)ۦ7[��qJ+�v��c:���8��1�o/�䲥������|�{�}�����d�Ƹs	u�O\u���<\�.�=v�����U�ɭv�s?�������SP%D8ےt�����k2���w1��|���e�����n�R(��v�t���-�nɌ���UL�$̢~�!�GH<D��I
S̪�;��=�ɣ�&N�q���ݥ@��r5B����?UUr���e��\�07jGL-��"�QJ褡���_�XU�sޭ߫�:����̖�|`T�Q������h�k�۞'���v�^���v��wE�s̀���h���.��07jGL-������UU�y� �i"���dF���n���Y>>
'U��*�!@3)��	�0J�uz?�����c��Ɂ�]0;je���VU�*�I^[ �Ɍ���ꤻ�|��=�`b�ck
j$�N6���7^��Ŵ�z3��N�{�@e�Ʃ��$c�R+��˫�+ޛ����;ט���Q�Sj�/\	WC��\.S=����]���{YͶ,ݵz%�헰K#N����7QW�{�uX��,��/�9�{M����H�
����0�1��r&���gd��H�4[tB�N�JD�ܖy�$�g;�R�N!�,F+C9�rY`��`w1�*(Ɗ��*g��ߕ{�� _�&��|��z ��4qD�N2'Q�Vs�x���g�2�u��^R�5�$�����pY�VW]́��C��歭��/[ u��t'����ӛ����;��u˱ϕ�����0;nD��N��; ��[-�)��rD���%���`}Y캰;��X��{��o�I#h�0=S����0ޘ��)�i��	��pr������%�;�s٩>C�����j�ք$§M��g��T�[��mX�����%B��!`ޘ��2V��;���ꪯ�~����uґ����nwB�t�;b��ݶN�<���`.�;�9�kv��-���z���Tz�fI/��٠3��j(�H��+��eՁ����;�d�3�د�����)�1Rt�SN��X{� �ϾVչ�V���%��%6
�6�,��K=�@|��J����i@c�؍��Rіb�˼�`M�����0&�A�o��u$)�$�Z���g��>3����vS'���`T�k�5$���Y�\pN�m�qu`��ge��̷3�b�7Qq�]�vm���s�N�蕒9�����t�
[ö�ѽ�ν�k�X�۴v���v��϶��\[l�kѯ&]vӖ�[c�h�zEq��r\��qltp�{d�'��:ͳ�s/T5��fͽwb˦;�`���Dh��������*Jd���v\�K%�y{��;�;��n;��8ll�c�GN��hA�ó�:�%={s�:m�V�9�.[�w#Zd�(��~w����7�w�0&�D��u]�W0q���
J�3��X{���K���U��t@`i�7A2�P��̔��4���93���Ҡ6�t�=f��О<$�4�&fn��ޚ�oR�3�8P��h�ȇO�f!]#+,řylT������,�;�x���&�J��H�d�#@�չ���^�L�\�F�u��P����n�s������('c��ܮ����`�XS��=S�����/���.����^��<�UU]_���ljO[�$u`{�ج��7��'�#nI`|�K`z�GL��ߒ�s��'O���2�x<L�Bf(5rh���T�o�`�X,�;z�<���7�<ʠ-�y74foO����>^̺�33*� 1��ے��R���;��ع;n&8�v�Y�v���݀=I^��97�X�
�g�W��7zc �����}���R˨���8D���^�$v��u`j�k���,y�j�TQ��*2I���˫}����|)���|mX1Q51�J `r9L
�L�E�p!��iP5]0E�| x��51���H��e�}�bx�GM�N2'J9V������`I�0	�1�+dt��ڋ،R���
"b�2�&��Qٽ>�g��V.���؞!��)'L���q��4u�<s��(z��ݹ�n�r�]�nq�6��7'NH%#��3��`ew2����c�s� 73e��ݸ�F�!h�,�`J�?�H�t���}�od���)#m6:{�nP��^�b�2�&�L���͚U�Ҡ�H�d�P��Ȝv��K ��%����F��mLY��2.�O�s�}�v�-���N�c�'���g���GL]���1���<H��uqt�qN�	�7)����K>����c��[��exy\�%8�Fx�N�g���e�*��"�3/'Y|���ؠ-�l��)��Rd�����`�d�>ǘ���]^�mz�D��ԡ0t�yl�����T��˺[Ub�xTP)��crX~�R���`mnmՁ��c��U%��,{4����U��]%���0;��`�c}�{u$A��M��`,)����1�Z���Y$�dBBB�(��J�S@iCL!1"i�I#�&��� BBD#.~�V�F��X!.�p|�)��D6%M�B3	�$$FI�X���,�$2&���3��a7��`��"wH�����[�̪�ʏ��j1su8�� ��E ��c�:+�C8Đ�jQ�aB#	�����r�`ʣ�*P�c ��ҟ|=>�!���P]p
� |�H�C��>��x���q2�c�W0�!	M�bA�qϵ����D�A(3����HBq" h~�jd�"��!�d��~H|je���*%&8F1�����{�w�����'~?-�~@$ 6Z��`  -� [V�      \;6Gv�-��@nX-��Õ�v���8��E&��т5=�+�k�5y����]�n�S'cr��'e.V^gl��ڳrsd�Xl�h�u�Y���v����[�G*�.U��M78��*�Ij��td�%x6^�b�3���u�Uڨ�j�����F�v�[r:W��s����2�u�7Q�l>ە�R�[�FB�����E��.cEu�������m�O>[��p�'Lu9�+��{^������7+q��3G�p��[���y�v�e���w&늛hKkK��Qm�XS��se�bA�D�{G �V�(۳' ���M +�����O(��ˀ۳gn���T�a':���w-:�d�[bN��-�ٹ5iB�����tS=�m|�A�Re-�IЧU��Zմ��uف8v���L#���\=��9�f�COl��!�n�66�u��'f8�����][v9;E��a2�wg��ƋK�[x56"d���gv��<sL�FV������%D]<p+��ON�bP,�j�x^�[��W��Z��W��]�]/�GjԒ�P�Eh�xx� �4:�G����ue��֒Ko���B%v����` ˝N��ԫ+ q Rv�6z���NݷM�u]p=����������	��� ����BJ'��B�f ��n�;�1�֍�O,9�𘺏*�����u\(�<�5ʮm�-5���ɷ�buv�6U���[d��l�i�6Ҹû+Q��7U��bv'V4�c9�t�b����'L���A��TX�U^��V�ƺtU��:� �^�[8l� I��g7m���u:��DAj�g��T�{m;/*�/-UmHn��J�����xX��ur[��.4���ٹř�ۮ��T,�R����p��55]v
m��W&�ŕ,shU��q���ٜ���@:&N��ȧ��d�:aA���D�T�(iL���H��`(B"�"�T""D*4@�Ч >C��b)�L(t�T�l��9�c��8�UN�W�Q�E@ىJ�.Q��v�$3ų=�/VC7����unhk�<J�뫶��0� *���{�y#��s���"�mx�o;�::�/�c�x1���M���9��#��V�-N��>� ���b,�=:�����%�ڹڵ)%]�6���͍�l<��n� ܎]=/�5�]׮cN2�b�6b�qm�-�3�' �s[15&rau��n�K�s�Ղ��=r<u�z��qm����>b�nK�<���K5����.3�.�&��#1��7���* ��i��*58����d���b�':`wvA��ʖC��Yy�ay���L	�:`wvA�:d�T�
!�%FD��inn�VfO��`z\��v�*^]�v���!������W76����V{2���a���(܂�#M�T�)1�'���M��1��]ۮ��J�[�#����w�.���R<K��Δ�/l�2�d�+��}�¤�&"X�'��~�M��d�'\.~��.(���e;Ĕ�q,K������p�"x�� (!�C� �M����&=���&�X�%������Kı=�kK�|r��G)�{7��PcN4�hJf�7ı,Ow�٤�Kı;���I��%�b{�צ�q,K������|r��G)�y�����U�4��bX�'{�zi7ı,Ow���n%�bX�{>��n%�bX�ｳI��%�b^I���ؙ���.[s���Kı=�k�I��%�a�H���~�O�X�%��߿l�n%�bX��u��Kı? ����C���l\�W%i��<d�;;v�8v�q�tTF���P�an������#�5�{���D�,N~���I��%�b{���&�X�%���^��Ϣb%�b~��~�O��7���{�~��+����!���q,K��}�Mı,K��4��bX�'��zi7ı,O��z�7�,K�r��s�g&1pd����M&�X�%���^�Mı,K���4��c�
�� �!J+��4�dU\��ı1���I��%�b}�{f�q,K��=��E�	C�/*T�S/�N2s�	@˷���Kı9�?�]&�X�%����4��bX��"{����KıW�"8D˺��J�N�%2�d�'8�{>��n%�bX�ｳI��%�bw�ﮓq,K��}�M&�X�%��z��}v9�ݫ4s{k��,ԛ�8� y��#�k�y��a��u�mv���y���6�p�c�n�q,K��}�Mı,K��}t��bX�'��zh?"�8��W����ᓌ�d�-��&IQ2
fLL�J�_�d�'dflS/��$q,O����I��%�bs�~�Mı,K���i7,Kļ��Ň�33KL\��3I��%�b{�צ�q,K������q, C1��~٤�Kı=�k��n%�bX��u�B���nnnq��i7ı,O��z�7ı,N{�٤�Kı;���I��%��Y�Ox'G`���뜚Mı,K���q=�ۛ0Y��\�g�Mı,K���i7ı,N����n%�bX����Kı>�}��Kı;�jy����L�n�\g���A�^�;��.�϶�@�.^M"G��K���IS��ۉbX�'y�zi7ı,N����n%�bX�{=���X�%��{�5���#��R9[����J$d�Ӆ��X�%���^�M��q,N~Ͽ]&�X�%��߿l�n%�bX��u��O�A�LD�9�߱f�9��	�-�M&�X�%������Kı9�{f�q,+D�Ow��4��bX�'����&�X�%��w��r��&1f11���7ı,N{�٤�Kı;���I��%�bw���&�X�� �'?k߮�q,K��=���IN@L�����_+㔎R9H�g����Kİ����~��}ı,N~Ͽ]&�X�%��{�4��bX�'���k�0O�-��I�����9�f<;u��S��י�Zp6۱O7R��k�8ܝR	�g���l.�9/S�݉^Au����8��Iڶ� ����S� r��lr;��eq������3&��\�nЕ =�v��ŝ�Fӡ���K�vn�����{U�ٲ�I׈.�v�Vqn^��Yƀ�d��r��G�nr�I�PE�����v�v�=���!�}�n�]��� v5���^g�ϵ���ܭ�u����g<kb�f���e�gS�,K�����f�q,K���ﮓq,K���wı,N���n%�bX���.�3H\���nq�d�n%�bX�{=��n%�bX����I��%�bw�צ�q,K��}�M��b�"X���b�藘w���D�1/L�8��N2����n%�bX��u��KK��}�Mı,K�g��Mı,K�{Y�:$�Ӏ�JH���G)�r��צ�q,K��}�Mı,K�g��Mı,K����&�X�%��{X�+o���g8�,���n%�bX�ｳI��%�a�c��߮��%�bs����7ı,O����7ı���2I%�*[���S���z��WZ�!zc�0F��@q�{r�vMk��ۊ���[��g����&��%�bs����Kı>�}��Kı>�{�@�Kı>�}�I��%�b{��6r�m�ȯ���G)�r�隴���SQI�A[S:��Ȝ�b{Y�.�q,K����Mı,K�g޺Mı,K����qXI��G�w���oq�s�ﮓq,K�����&�X"X�'�Ͻt��bX�'��}t��bX�%䞞,����-1r[���7ı,O��l�n%�bX��}��Kı>�{��Kı9���I��%�b}�v�zf��1q1�ۜc&�q,K��3�]&�X�%����}t��bX�'9�z�7ı,O��l�n%��ow���}ں���٨v׶�b�3�ۋ��v�{nݶs��P�n�0:u(�d�K�f�7ı,O����7ı,Ns>��n%�bX�s�٤�Kı9���I��%�b_N{��	����Is���Kı9���I��X�%��{�Mı,K�Ͻt��bX�'��}t��bX�'��c�2K���e��Mı,K���4��bX�'9�z�7��Wh�SB��(8T#V�n��� a��	D�3BE� ����b{9���Kı;����n%�bX���b{5�3)�Ypff�&�q,KB��=��7ı,O����7ı,Ns>��n%�bX�w������G)�r�r�ʂ#C�F��Kı>�{��Kı9���I��%�b}��f�q,K��=��+㔎R9H�y�� �j��M��i�\P71��\�<��#�>|m{9Ͷ,�uu���˃�=��G����'�������oq�����I��%�b}��f�q,K��=��7ı,O����7ı,K�=<Y�1��Zb�9��n%�bX�w�٤� R�$Ns��j	 �w��)"}�{��OD�,O�ۯL�%ɋ���ۜd�n%�bX�罽&�X�%��s�]&�X�%��g޺Mı,K���4��bX�'}�b�_�1qqsf3-�t��bY�V!������7ı,N�?�]&�X�%��{�Mı,!�R@$�1_�=��5�s��Kı=���c9�	��\fK�%�n�q,K��3�]&�X�%��{�Mı,K�g޺Mı,K�羺Mı,K���߻����������G�����{]���`������;�ۧ�~{����>u�u:�Lc�O�X�%��{��&�X�%��3�]&�X�%��s�]�}d�,��ze���N2q�B�bGYŗfnri7ı,O��z�7ı,O����7ı,Ns=��n%�bX�w�٤�ı,N��ǲfY1��cc9�3��&�X�%��s�]&�X�%��g��Mı,K���4��bX�'�Ͻt��bX�%�����L�3�qs����Mı,K��}t��bX�'��i7ı,O��z�7ılO����7ı,K�;<Y鋜�Jb�9��n%�bX�w�٤�Kı>�}��Kı>�{��Kı9���I��%�b{��#q��֩��L��t�ͭ�*�WS�u@)%���\���&kY8׋1�aՓ��ZI�œKĉ���f-�Ny4�,-G=-̽Ót��F"J��0vy�ggL�z�3�n�ṙ1ص�G�s�t�4����㣷'r4�i���,�<��%��U�E��4��=]vt���X�.`5ٷ+Ý�xyy�a��YE#t�j�]7��\����/)��u�=۷w{��u��k]g�tmq���M��ζ�\�N\�wZz��m���.`T--y�q��X��r9�&>ND�,K����I��%�b}���I��%�bs�ﮃ���b%�bs���I��%�b{�����1p\\�g�3t��bX�'��}t��bX�'9���7ı,O��l�n%�bQ��w^�|2���N2�Ӹ���L�\fK�%�n�q,K��s��I��%�b}��f�q,C1����I��%�bs����Kı>���a���1��0fc��n%�bX�w�٤�Kı>�}��Kı>�{��Kı9���I��%�b{����8̦qe�����Mı,K�g޺Mı,K����I�Kı;����n%�bX�w�٤�Kı9��M����û=�m�z�SVC����.�ַ���n�펛G7a-�ۗ��Z�4�3SU�n%�bX�w=��n%�bX��;�i7ı,O��l�n%�bX�s>��������oq���}4u�l�I�t��bX�'1��Mà�EHdH�"�>��	0�Q)DC`�H���|�x�&�8��'�,N�~٤�Kı=���I��%�b}���I���G1Ľ���g鋜�Jb��s�&�X�%��{��&�X�%��3�]&�X�@�"b'=�~�Mı,K��cI��4�R9]Ҳ��B���(�_+㔄��9�~�t��bX�'=�~�Mı,K��}�&�X�%��{�k㔎R9H�f�ŵ#i�$tG��X�%��s�]&�X�%��s�Ɠq,K�����&�X�%��3�]&�X�%��1�OߤͰ��3�)q2+�[���[�<�h�d�s�q�\��Z֭�e�<���������q�IRJ_�ߔ�Y�,N���&�X�%��{�Mı,K�g޺Mı,K�羺Mı�7�����|z��3�~{�7��������&�X�%��3�]&�X�%��s�]&�X�%��s�ƓqUı=����k�fS8�����M&�X�%��3�]&�X�%��s�]&�X�:���������)��+����8ā@��.���
e�d�Y�,4I��p�G	&�L�pU���iӨ�F��SQ~.�\����hjL�i%)}���*��a��b�
��M��T	a2�M�� B�!(@"�ʶ��}XVR:b�a��`�5$ISHH}��432E��� ������tz(,A0��L�5���P*�Bp�Q˔:�U~p�S �|b&bk�q��Kı9��f�q,K��3{�2����s���79��n%�bX�w=��n%�bX��;�i7ı,O��l�n%�`�؟s>��n%�bX������L�39��\��7ı,Nc��4��bX�'��i7ı,O��z�7ı,O����7ı,O�=���39̜��ֺUz�:F��c����8;n�Q��n��㎨��ԕ���7N�pr\M?��X�%��{��&�X�%��3�]&�X�%��s�] ��X�%��s�w���#��R9]Ҳ��B���(�i7ı,O��z�7�$q,N{>�t��bX�'q�~Ɠq,K�����&�X�%��wX���3q�ř�is��&�X�%��s�]&�X�%��s�Ɠq,ElK���4��bX�'�Ͻt��bX�'q�_\g9�33�$@y��_�d�$��e���L��,K���Mı,K�g޺Mı,�Y1K8	�z�Au������Kı>���\_̸�Ř3.1�i7ı,O��l�n%�bX~P ';�߮��%�bs����Kı9�w��n%�bX��=}�qCZ��3�m�i����Gc��z	�q�u�*qt���m�mۙ�zlt�z�]�����%�b}���I��%�b}���I��%�bsﱤ�Kı>�}�I����ow�����Xp�j�MG�w��bX�'��}t��� ����%�}�:Mı,K���Mı,K�g޺M�������b^{��\�&s�����.st��bX�%�}�:Mı,K���4��c�!��������Kı;�k��n%�bX��vx�����qrg�s��K�,O��l�n%�bX�s>��n%�bX��u��Kı/9�gI��%�b}�{X�q�B\��c36g4��bX�'�Ͻt��bX���{���O�X�%�{�~Γq,K�����&�X�%���+�X��iZ8,���k2g79�st�[��f����5#��yɍִ����(�`A,�"�F�_�|��;���O]��:�X�zt��ΛzoBkm�)���]Iӈ�%�oV:���U�6�Kz�K�a���m�ir���rݫ���.#<v8����Wm�c2��l	���$���ǯV�;\S���MѬ�m�(����Ű��m���ݺ �V�:�(��is�2�aq���
�C�������aK��8�j���.^|v!$��x8�ӻ/e���.7aQ��+�j��}ߛ�o%���k�I��%�b^s�Γq,K��;�]ı,K�g޺Mı�r����V�:�c��p�W�)	bX��ﳤ�Kı=��f�q,K������q,K��;�M&�X�%�������2[��ɓ6�Γq,K��;�Mı,K�g޺Mı��;�M&�X�%�y��:Mı,K�;�Of��e3��&3�I��%��������Kı?w��4��bX�%�;��7ı,Os�٧�7���{�����~��-Z�����bX�'��zi7ı,B��t��bX�'��l�n%�bX�s>��n%�bX����9&1e�&sHc8��n�K�m�d�gz-���b��q�7%v��N�[r�R�J����W���#��R9K�͚Mı,K��i7ı,K�=��?*O�b%�b~�}��7ı,G�ӓ���x��*b&f�|2q���c��i7c4y�>:��n'�,K߽��7ı,O����7ı,K�w��n%�bX�v�=�g�%����qq�I��%�b_��gI��%�b{�ﮓq,"�1����&�X�%�����I��%�bw�����Jr��Xk��{��7����È���~�Mı,K����&�X�%��w�4��bX�%���t��bY�G+�6�$M8
7�9H�(�%�;��7ı,Os�٤�Kı/�����Kı=���I��%��{��O��D����cg��Ȯ3N��-�z���v�����>{�uA��1.ns&Lیg:Mı,K��i7ı,K�=��7ı,Os=��~ g�1ı/{���n%�bX���؟�\�2��n�ɤ�Kı/�����?
�q,O�Ͽ]&�X�%�{�~Γq,K��;�M���=��;�ow�ۏ��#i�T�_=ߑ,K������n%�bX��ﳤ�K�1`O���A�� :5q1�~٤�Kı/����nr��G)��f�B�IH�pR+�|%�g����߳��Kı?w߶i7ı,K�=��7ı,Os=��n%�bX��vz��g7-�ɜc9Γq,K��;�Mı,K��{:Mı,K��}t��bX�%�;�_�d�'r�4�e�8DD�(x��At1�O����ѳ�������ns�H��K�9B��\mH����oq����s��gI��%�b{�ﮓq,Kļ�}�&�X�%��w�4��bX�'~����'Jr��Xk��{��7���s=��n�B&"b%�{�~Γq,K���k��n%�bX��{��n'�����q�߯ݾ��nzDm�B��w�Kı/{���n%�bX��u��K��LD�����n%�bX���~�{�{��7����}����F"����7ĳ�1�}��I��%�b^w���7ı,Os=��n%�`}�q�E�T
�!��6��
)����0aH����'ɠ~�L{;�t��bX�'0w���fsi���1��Mı,K��{:Mı,K��{��}ı,K���t��bX�'��zi7ı,O�e��Iy��R0����l0S���磜���9������Q�v�喸���U����w�%�bX���~�Mı,K��t��bX�'��zi7ı,O��z�6r��G)��f�B�IH�pR+�}ı,K�w��n%�bX��u��Kı>�}��Kı=���I��%�b^I���f�����s��Kı=���I��%�b}���I��?�V"b'��߮�q,KĽ��_�d�'{*�A)��g9�Mı,K�g޺Mı,K��}t��bX�%�;��7İ?2�߸�_�d�'omt�LC���\�$�3t��bX�'����7ı,?q���t�D�,K�}��I��%�b}���I��%�bPd�������ww�����Y"��88Х"캩�7�A�NN��c"p�-�i�9l���ݰ�%t�vE�ݷbIgFl�V#"��4rU��6�t��&�9Q��7]bƭ�l�ɮ�\f���.��g9L�u�d۲O�^<>>`ѹ��Ԗ��<"��	�E��[���B�8�A뇀x�r9;<YMۊ�;���js�7��,b�.luJ�&�]��ɛ=��^����ߟ��'�9Uf�6*f��s[s�<8�m�s��϶�q��/'X1��F�������w��7���{�����Γq,K��;�M&�X�%��3�]�UY�LD�,O�Ͽ]&�X�#��wS�GI)�bd%K�D�2�d�'X��u��?*C1��s���n%�bX���~�Mı,K��t��bX�'pN�ǩ$�a�\bd��f�q,K������q,K��3�]&�X�%�y��:Mı,K��4���{��7���q����U�����Ȗ%�b{�ﮓq,Kļ�}�&�X�%��w^�Mı,F�������{��7�������ͺn�RM�>{�ı,K�w��n%�bX��u��Kı>�}��Kı=���I��G)�r����V���1��';]X�:��4u��Ӻ�	�kqi2���;p v��rFg���.qs��7ı,Os���n%�bX�s>��n%�bX��{�ı,K��t��bX�'x�Xk`P�$ڑ��/���G)�r�麴��C�B!�.�j%��w��n%�bX��ﳤ�Kı=���I���2�e'omt�LC���̺&%��X�%�����&�X�%�y��:MıFı=���I��%�b}���M|r��G)�<�5dLiĢ�9|�ı,�01�gI��%�b~��i7ı,O��z�7İ? LEvoz�|2q���e}����Jw��!*m�3�&�X�%��w^�Mı,K�g޺Mı,K�﷤�Kı/9�gI��%�b~v��b�.q.�9e.�i��E�.H���趸�n@q�{r�Mk�k��;��n���l���u�m����bX�';�߮�q,K��;��7ı,K�w��m6	"{��SP@L�њƏ$�̢bf&%�2�g��SQ=ı/9�gI��%�b{�צ�q,K������qPKĳ�����*(H�p�_+㔎R9H�~�}�&�X�%��w^�Mı�"�"+�;�&�o��.�q,K���ﮓq,Kļ���{���.f3��7ı,Os���n%�bX�s=��n%�bX��{��K���,PT�Ls���&�X���������r�0�o����7�ı>�{��Kİ��w^�t�D�,K���&�X�%��=�M&����ow�����s;��U;:��6x��t���\5�[�۶��z��sű�;cSL���pL�7I��%�bs�ﮓq,KĿs�Γq,K���צ�q,K���ﮓq,K��<v�H1(% �QG�9H�#��R�e��T�,K�{^�Mı,K�g��Mı,K��}t���1�����:IN��%K�D�2�d�'<Nw��M&�X�%��3�]&�X�%��g��Mı,K���:Mı,J2�Fj�tH���CĔ�ᓌ�L�'��}t��bX�'9���7ı,K�w��n%�`k��DJ�S���2o����i7ı,{������2�S��1�������oc��4��bX�%�;��7ı,O��zi7ı,O��z�7ı,{�����}�H+�ʚ�!t�h�7)���L����lS:C�Wn�M�[j9�T5�	��Mı,K��t��bX�'��4��bX�'�Ͻt��*},K��cI��%�b^����O���-��s���I��%�b}���I��%�b}���I��%�b}�w��n%�bX��w��n%�bX���ZlRN8�H_+㔎R9H�w�5_+q,K��ﱤ�KBı/�ﳤ�Kı>�u��Kı=���N�5��c��{��7�������4��bX�%���t��bX�'��4��bX�'��}t��bX�';�v�@�VX���w���oq�����gI��%�b}���I��%�b}���I��%�b}�w��n%�bX�*ǌ�l�*���tuD*�Td�A``F��4'�F�� �В��D�-)BI!��0�"�"Ā� �5Z��Ua!	0��	n>&ɖFX�K��	�AI��Gd&(?�o[`5(�
RP�� G��K�'0.7��6�E��W@��h�0_�)�`Ͼ4:b0��h@5˲2 �4ao��@6l���0!��@�� �p���@���S(���\�(�s��p5?k�.ͤaܘ9��P��	���p��#�VҦ�I�P��C`�9�Ҡ�Z��6��o|�����K�JP������X��7d!�ʘj�����=�s�wo���ʶ�����[�  [@"�  ~��  �b���H��ce�[d���z��(3(q Nc�r�3�(b�dK�Wul�`9��1ڹ�M'�o'=����DW@5�j��Wb�Lq�qȼ��ɯX4*9�ݓڜ���tDa�v�cv'a���*����j�-�c���.Q����I-���^Q�ٖk3Z�n�W�e�f�;njT��sN��T�97h�r���Ks���5E.`���kg�/6�<ի'j�箑�q���r�@�u��g��N�t�W1�7H8�h��{`ǰF��]�-�] �ۣ���ӗ�g�vW#��1 �k(6��[X�8���*������e%��۳Ʊ;��(��:���>�AM�g����`l�s�a���GdsE�M��	��m�m�ʊM�e�g�ڢ@�g2�v�6�	3�=<!6�.˖9��<tw�	+���v�ɴ�U��aʶ��7�x�i�Y۷��L�^]��9gڹ	�u��a�^&�M��lsB�-��մ�V����pVz�`�3<M�Z�
N����$x�������9�]!׹��N�f9��`�앇�n�mus&n���7W�=��<Y�vA]���7^�ٹ���Vݹn�����Cu@ܴ�����;v>|2�n�hM�	o����hՖ���c>i/2��K��جi�8�"�[I�t ��A��s$���mV�b�N��kf %��@�R��8=tx�r���ϛ���[VƩD6}�^CD����ِ^V�v�Y-]+�괂e���s�V{[7Cj�L�gn����C����.�؃:�-E8ƞ#�[��U�BvRZ�Yƅ�����5�*��T�*���wd�I� l�vE�
]��4S� �9@�{$��;�n'��@�qb�;��7��i�^��k�r�.�)��.���MP*�\�֦��VY��«���Ԑ�	d��bg8�rf`x<GI�D�(| O�U*��z�Cjt���@��P2!͟pN���ͼ���UV�\�:�
	�5F�-j�h�4e��L��[v�gv&;hz�.vճr����fIKq��Z�b�c���x�;m��t(�U�&N.�S6�#oc��w63�65�g��y�s�����iA+��叹�|��us�l9�Ü�yۖ�δ��;
U�y⩺^u�[N��uk��nM
����h�hg!�kvV���	)9�h5�aw��w����r�_v�J�Di��l�Nt�T;�>k����r����+�s���1ӫ����=�n̸̙��t��X�%�~��gI��%�b}���I��%�b}�w��n%�bX��w��n%�bX�ē�1�I1�f�bf�c9�n%�bX�s=��n%�bX�c��4��bX�%���t��bX�'��i7�,W1���{���"H��	�����_�d�'\f�S/�X�%�~罝&�X�Xb&"s���I��%�bw����Kı/~�����Q,�������{��7����t��bX�'��i7ı,Ns=��n%�`��9�cI��%�b^I���n),��s1��I��%�b}��f�q,K��3�]&�X�%��9�cI��%�b_��gI��%�c߯��o���Ѡ'�=�E��r�\v.�za���&h�G�J۝l;ʧV��J�n.q�I��%�bs�ﮓq,K��ﱤ�Kı/�����Kģ/^oʙ|2q���e��9�@�1�8��n%�bX�c��4���k���O�|"j%�q��gI��%�b~���4��bX�ew9�L�rM�N2��ނH�_%���q��Kı/;��t��bX�'��i7ı,Ns=��n%�bX�c��4��bX�'���}�ܘ��Lɜˋ��I��%��H���|i7ı,Nc���&�X�%��9�cI��%�����w߳��Kı?@�9�"�x�Hy�L�8��N2�ﱤ�Kı>�;�i7ı,K�;��7ı,O��l�n%�bX��^���Q$&P��rJj%�y�/������*�ۘm�é��f:6��۷f�l�m3���7�{͊ �����)r�ɽ�7��~��RRR(�tI�}�d�33&gsכJ�=y�@|����p�ZmR�T �29,�6��>�Xr�xA�O1=֨*o�?o�Nwݖw�U�	I5###�a���]�l`j���oL`{z:`I0B�`��ĩ�rX.����}�>�ͺ���,�3$Rq�R�&JmԨ-��c�;��ړ�'i�����]v�+vL����w���h�Q5)&� w۲���˫ �}���w����ir8�5�&�������wO��oO��{d�@{)�$�I�IV��%�}�d��+��H�e��f�X��s����H���}�,�ݖ��]XGs�r�J��/�c�a�j('))n@L��{2hI�%���|�f� }�d���P�:��D$MԤ2-���[c���0[���\q�l�Π��s��ej�E�y�oGL���oL`�d�3��ڬ�JI��}�\�32N�'J ���~��\�&fH��!l �c�S��#�;�4���h�LJ�Ǽؠ=j/&!:X�e%hŘ0I1�����t��酁�d�r8�5�$���@s&L�"�c�=�:P�y47�������ߢ��UU]l�f(�s9�
�k���r=q��!�ݻVݽ��Odu��W5v��9.7/n��[��6���ݮ�Ê]:3�C�1�ok�v�`��K�8^Mx�v���������g�8�(S�'v�F��5�:ٜs���Զ��{�p�v�v	1�����A���B�c�;�|޹s���rr��;��nѭv�=�c��6�ύ�l�,m�_����ﻺ������@Gi��A��tU���@�c������׻q�u�*quʻ��<{m���9�J�`j��;ܘX��{�u`y��7!���ra_��~32M��@fwR�-�y����QD��#q�8Xw6X�e������0q�J^+T �.^&h{2�o�Ƞ=�(5.fI�/����66��RMH�"r�.���2Ӧ07dt��8��)+Bg�%v�qN�n�OJq����0�����+Wb���nl<񛰸�k�7T�?6�����0N��ݑ�����_D���)�2P�y5�ĳc3beɒ���]X������a`}����N�*�9%��za`yw���\K=�K �f���x��ND)PI���8�����|0	�1���@l�KM����G#�=�L,ܮUR�fπ������c��#���У!��nk[���s��\��$ʚ�Ovx��t2Wm���ȉ�$�5"����`��K������od{��/ݫ�#*���`E�-���6�cݯY t�R22HX��v���jp�O*H��AAq S�`��� �� N���̛$�[��w:P�"q�$wx�q8�w� �ײXg�U�-~�vk3Xt�)(��6�cӣ�[����`l�%ftKX�4,����H���w*�y8���}��.�p�l��v���#r1[8���GL���;{!�y�T��L��ND��4�`b��򪸑�ɥ�o�vXg������4�la��l��0	�&0=::`E�-�{Ƣ�9N8F�dp��r���-��4�6��w�@��
D$��&�V��2�ISZP�	�b^""�#+3�0"���� �^�`nx�W)����q7Cq4�*D�C��۳�vv��M��v�i�7�:� %����[f�jFFG+�5{5����d�>�eՁ���c�	60�#��`{��0	���0"ޖ���I����&ܤ��HX��e��{.�]�;�����=1���fcӣ�[����}�/�����m3�P��'PjJ�1w�����RIߎw:�o�wF��]�d�*��wv��������-�EUtt��+��v,�3G%��-v3�1���t�n�!�`ո�6�csn����D[Fn�1@	��
);JN�Qϵӡ���e�au��U����X�Ҕl�]e]��5�u)�8�0��sI�ޒ#�]��쪘�ͣ�:N]l����{S�\���5�z�d���Flwm�����\+m�'6��r��V��X.M�9�\�ó�Kϓjd���z���P�K�D<�<L6�:��`�d��������>qӹ�g�u�nn��F��m��������3����]X��v�3�$�8�������oGL���=��0
��#���	NK��.�]�;�} �]1�6�K?LWIxe��9�b�b���k�y^M��7�@n2��R0I6�q8�u��z1����-�l�9��eb�e'LӺm��<..�J�s�p��)���}��7''\9����;n�Э����o��~���09o,}{Ɂ��^^+��9���s�&��{5�D�D ��@F HF+�v���L�y3B����E��y^MmUq#P��mBB���,^�v��&6�c��@l�KWx]݅�y����D�&�L`{{ ����`��J(���n:�E`��������=��0<���R�����]�m�ı�r����:�G2���]�;������=Yۍ��r��|�~?�[������j��ĕЃ/�3[������,�酁�f�F	'O�A��>�^= }������u�ۦg�����e0�I"�$3 HC �!>�8@p�a����K��>2�1#0I��	�"�$\w ��#t!�BB{Ȓ�	�O��8$a5�@�7`�p�M1�����M9��ڦ)ϡt1�je�u�&��8/$8j�Tِ3�\�L.�;��.B�C�2A�X���,�iGQ�_�&�`
���f�'ei��8�6noB6F���3��8�a#�g��@~t�@H��a��;1�|+"i>d�r�6�&pS;��&�h*� ̩]��Fi4�@t
�N(��t"��dC`&�����~@P�� ��j�p N��\�lE�4T{�^c��e�����E�
���r���Ǡ�i�4�'JבA���'��j�;�5�H�n9��K��a`E�-���z1��U��WJ�gmip�]n�c���(O/���M�}ǉ��m�&�����d]�s��6���?�܊�E���^N�f��ד����pm�r������>��,�酁���{T���ԕ�'$q�����`{{ ��z[ ���_x�R18�n�cQK��a`b��M���Rg�ﲹ�F��C�ংP1D>������'��S�N��2HX��v�}��>��,�酁����4��)��Q�N����$vv�s�P��5���۶��yŰ96��:�A�ԌN�����}�,�=�����mW�5{5�토*J�(Q5���d��$wٷV�f� ���{�U$wrj!Dq��r�%��>t��z[ ���6�c���U)�R�4�a��U-~�v�f� �ײXo)w�zX�oi�$����`ޘ�=����t��zcRL����Hr��L�\�櫣�ӵ�Θ�h[�E9��Y:%%��8����\r`��.�']�J^����z��,�zܔX��:s���Q�ˣnXȇ6T<�U��a;<nQ�Gn-�2�m#�����b�gn�R��ƴ�.��H���t�2���'Wț���XG�6z;"y�6{[q[��.���2���$�LX�Ʒj�M�O+�W��Z3�n�*�w7�I%72g��1s�e5�V�N��wm��;1�8����6سv�b��{C�(A�Aȣ�$� =��e��}0"ޖ�=�1�W��Eywwuye�*�ގ��U$|�}lz}���K��U$o�JS�RN��29V�O��{zc �:c���u�P̰I]_��/.����0C�0=�X~�Z�����P%c�(��K �:c���-�l���t�����#K����c���u�2��F��>�0u��x�Om���X-a���f0=�0"ޖ�=�1�z1��tx�UJr��IV.��+�J�S��@&@@�5&3�gRI��vXw�u`gZ�bm��@�#����0C�0=�0"ޖ��蒸��A�GI%�}��Xw�u`b����K ��x)�m�NSdE�0=�0>�������0T������������Yqz,V�n.5fL���b�\oI=�n��C�M�O�l;����/�/+�E��`ޘ�=S�0=�L,y�,$`�t�$N7�}�d`����09oKߒ'_���<��<�<�� ynl�z�
-re��(l��$.S���BI42d����f� o�f��/)��F�q4T�$�>��}��>�X՞�`}��ʩNB��A��ב@o(�ޟ Z��>���2?�����Ӳq�ʴ�z��<<+�Q�*���7n8u<D<G<�����B��m4��ޘ��'L`{{ ��-���k nn
9I,���`}�L,.��}�d����� �(����07�|09oK`ޘ��'L`M�)N<I:G�!`yw����%�7gy��L��(��`0) � �D4�)�UN���X�0�R0I:|�'��>�X��'oO���‷��P�&|�uA�G�c�\���s�`��s!퓴��6�\.K����Ɏ_f�t����	6xG��`{{ ��/��^@oO���͵F�$N8� )%��}0�<�y��&��̼��\��F�ô��"��IP����&�fg9��@w�4�=�Ie�n$�Q8I#�oL`y�0=��a�R���`N�@���@�K�g�X���^��y�@z�h�a$	��I����MU�p�]<�g�ʫ��J��v��v�t[	���kj�ڒw����<�3��f�[p�1��b�G�Y�DqQ/n2�<�v��uB �����]��^��⸟ۏ;{�o���bU���� qn.�źZ�񧞞�#Ny�!���W��h��̴�%�5�uguP�t�%-�xWhQvy��h,�u�+7m�c�q������%�ns�Av�A��l@f��b}��1&s1.q�����t�C�:��[�>��� �;���+l�ԍ��<#
DQ(���NN����������0<��Ag�+�^ff[���L`y�07z:�UI��]H�Cm$N7�w۲��̼�?���m*�b���̀�)e����:cgGL[����,��j:������)�`w/)P������{�@y��"���c�����mY�����=��604�c�O]ی�^n�Wm��8�f�unp����˾��l��յ%�6tt�޺K�bm���D�$��=��s�ӕO������B$G�T��Cc�v�9=|sXԇ�r����c�;�aj �RP�"f���fE�fR���;���P���}��H���ʍ)N;�̺�5l��7d���-�;�2ʸ��e�,�`j�-�nɌ[R[veՁ�<bj�Bt��L�R��R:j�G'v6�ӶюGn��m��v+�>�a��k�����u�=#����H�n?�;��`uv����.���;�+1��F��I`jڒ��05l��=�cӣJ�J���Jq����;��gz���:a$s�0���UF��2Y����_tP�E�ô��"�]ayyL[%�l��յ%����ٿU��:K(��q%��I�}��`jڒ��05l����"�}v.�����N����9��!�W�h�����J�䞎-���|��a譔�V����`n�t�ղ[ �Ɍ��{����ʍ)N;��]_�$y{u�}�,��c�=�#)�IЂL�e05l��=�cVԖ�����f�4�RD�q�o+��~�~��1�wE�^R��k���v�V�L�3��d%$r�:C���|��k���>(�P�q�,��c�7z:`j�-��d���Veb˼�\=1\6�a�)sŕ�;"K��5����s���dsƐ�D�ӑ�r6�L��;�˦����K`jڒ�.����-HS��U������I^�v��u��e��9�U$yQ�SmĔq�◙l]���յ%�7dt�ղ[��ʵ(N'�ڡ��7��^~��`^�Ҡ<�̊L��/v({�漺���4�9,�2����z{u�Y�2O��Ƥ��EW�h���DEW����@DU�"��@_� "*��QPT������"��"� *X�,�"��B�`���"�R�
�U�, ",D ��A�"��B���P�"Ă"�"�� ���"� ���H�,",��"� ��"��@ ���"��,R���",",�, ���"Ċ"�H�"���"Ƞ B�(� �@"��",�*D�"� ��AR �A H",@P�*EH",D�"��X",R �D ���,A�@DU� ����EW�"�P_�EW� "*��U� ��� DU�"�� "*� "*��1AY&SY��̌Y�hP��3'� a{���  �      h  � @���   � |�*�R�J��hhʹ$��**� ��E$�R�UH@JP�� B E
 ��w�    8�@

  P���zۤJR�s�N���@z{��:o`A��'g��47`t����C��:�  ���x�� w{�6z�9�/u�w� ���EE־Z�޷���٪9o{���  �ϠE�h
�խ ux��k�O����כIw��Uk��u�{�(S��ztw�O=[�kا{��s�W
�+�Gy�p 0�juO��_f��&� ��<��`���·�}�A�������G;;]gA ��@ P ��J�� t�>��}�gV� qy��^��Ӿ�73�1zr�zy<�g�}}"����й��  �vOz�s��-���@��Cs��{�{<OA�a�r=:y�  ��t�� ��-� ��A�á���sh;u �}��;Z�y�C�Þ׬�x����7a� !�{���-�Q�w7��:S��C�����^�eI� ـv����r{۠@ ��  � ��ʶπv��5s���7w��� >���
ng@��@YJt� jחo)M4ܰ)KX   i��r��l�M��ѓ���:h��B��`�wpJX���R�;�� 2�R�YJQ�w{�R�  |D�&��R��� ѐO��6�h0#LOb�T'��� �Oi��lUJ�40�Ѫ�m)J� h ����$����mW*���O���g���c�I$�\s%r8���P(
���@Up��� �*�����tV �"�����	LE�Ԯ2�L�����
`ʚdH9��@��,�B/ �8�.6���t�	q�� t��O�@�2�e���(K�aF��.�a��iX8B�b��a&f�s�*�#���b�h A�@,��[�����Dr����R1	_��!G��^
��R��P�zV5�2H0.�7��5˖8(�),R	a�)�X�e!�)����r}��э@��~�ܻ�'�82)��y�)�,���b|s\��o>;&w��ƌ�:�.��$l*�+
H9 �,*:1Lg�0�7.�@�jEb�N|fg�o]�7�1�sx�1N���
<�i�\!�a$���HH�HYE�d"�"4H���XC!!	�fsvP�.�o���"+L)�����~�GP��d�VB��!��7���ß���K7϶ާ��ϜWG}��m�(�R�诹�R���L�_f�1��`ˬ�X&3��jh��jK��L�Lgf���|�n�� ��c�LR�N���/�~	.�ۄ��L,`0c ��1���	�HR)Vx��.�L�0bkBVD�|�$k$�����������L�rgs�iʽk�G���.K���B�hV2%�B�������7���i~8��3�gd�C�f�>q�:'D�dXg�b��n�e6�Ƅ�\8�Ŏ�02;���c��f�S�41	 Ӏ@�����XEcXݛ4d��-�J��B$�%10����`��x&&��fFǆ�*B	B��"B�(���`ո)��@%���dXS@�������
��H��o�ܐ�1�G���Z`�H��	`#��P�vfr�?v�&&XW-I1���gZ>����;��E>tB�_�k��mJ��.��Ą(�������X��"� 5�y��qd1��7Nh�&�dF,��l���#$	$a�Ɯ�Ѽ�N��e)��P���ri�$�E�*�A�HK��Ē"�k��Fm�jsY�)��#p�n�ְ�&ͱ�!dM�J��،�T�_���A�$�Ѩ��sD8�HXYh!Y��9&K�@�Hb��B8R@�Ŷ�3&�*p�B$P�3s��s��9�J��.P��+5��Xd��uO��q��wlxD+�WVLc�ֈc2˖�I�8��>��JO����0�Ė���I�+ȟa��du�)�A�@��6`�saXSD`i�$�p�#H0�e�P�0d X0D�)�Hi
�ă9��N�� ����)-�:F'Ƙ�F�k���F��6©!0�ZB�_}� ҄��f$IRO��>��8���%�(F�T�[4�sZn�bp�
I+��HU�u�9ᢨB�"F
b���@�i	X3
�i��͆l�7�3�L�����cL1�����K3�b�{Ϸ�І�%��ad��K��8��:� Jc<��3s\�M$6%�ψ�� �bȌ �&���8"\c����s/a�(�`� &,)F Q$!�FB	%� �"�P�X$bЀ��
�}��6g�^����u��¦�@*HBAH�1F)!b�-1��A$j`4��H�X1�9�2J�I0�8L�,Z!	�0�$Hd�$F��"���	�$�&�)GE�pePÓI�}/4`�L�4JE�(A+P�0��X�H��C%�x�>H��C26����`X\q4�4q�5�]��JH0\�t��֤�2��!�w0�2�e�����K��%��HB�B�а�V%HQ����\��C�sL8������7gզ3t�c%1�����h.跅3���7�J���������V[n�u�����s�E�)��1ْ����W�)�~5�y&��}�o/�	!0c�$�8���(D*K��r�1����J<6�9��(K��ai�$.vL���1�]m���	L\�:ISѓD
�1�\��:�k���{HC_F7)�XDٜ�RV]g�>��u/9�.������C����Q�p(�}�S�7V%��ˮj�`M��n*gH��,����f�!�7�k�vj�Y�XLS_}��6s���%>ӣY8l�э��h_�3��\:+x����a��&~��xN!��7ϣ�#��H�
J����%���O<��I�K�%���:����~|����O���!q�'�n<�>y��ya�%���qe
|����%���=f%�������O�^��3	XIr�L[��a�S_AJ� `b�b��B�J0�n�]�2J� �1"S��W�FHP��DÙ���I�2+h}B4��)�1Ϋq�5pH�}�7��_�qI3�!7�3�c�+�1�e���p�pc�Nr7Ѱ�ٰ	&3��6oX�!�w�INc�)0\��>�xlas���۱�6��(�8P������g:�_��?Z�����:�����gKw�Ý�����}��Z\���/�6g%r�+s��7Fn�>���@���N2���L��O�qݴ�t�����HGo�0�(�����)F�2B1��dH�aH0�8H� F3He��H&S*�"�ə�.q�y���]HK��0�,,#5���MƐ �0HB��A(#H$si����%!deeHRI�!I����`B!��`b4�B�#�����#8�0#@�I��$�a�9��JL��rݕ���
�ȹ
�4�� P"$���2�8�|a.^��D���1�lΜw|����gs�7����L.`�0f�NP��C"h ��$pe,�P�,
T�)c�f��t�V2`Vj�z͑�f6�IS�+.f1���B�
B�c&w��Ze�(}�Rb�$�ajB�H� ��.
KpI�F�����@���@,�BR)1�1r}��	VR���!;J�j�$CrJF�{�uK�bg�s�s?M�t�����(��U#/�ΝgR�.YHi
d	d�+�\�gc9����$0q5R6�ɤ�L�;�#3L,�H�-��.�n��.	�LkD��R`Y# ��5+�Ip�LBư"�4��.3�"4`B2-�$�	ag��.�8�B�_�����%Y.�ki+u��s).��I"�R��1�(�$.4!s����К�3��`|O�����O�?�er����F�
Bȼ��3��1�t�8[�3����ǘEy�z���G���~^%/Ӝ����~9�k�NL����{m7��..����~��$�B�n��Z�	�
+)��	�c�HζT�Ra+�I83R�2B�r��͚~�HR�#}]j�!	�%�iӆF�s��F�X;k��K��[�\|nSTq����~�R}B���^0���.8g��]c;IR֧7��K����nw�u��КM$�NN��a����u'.6� @�R@0�o�o6���֣H^C۲�z+�,2�HgV�9�$ٜ}kd+�m�6�+�7<���C��R) L�Hl�2d.9���~p�+)r�g���c_;5�JK�b�gZ�讳�XYip`jR�1�И֫
�&�s/��e�m��|�ێC��)
	�h��&�����ð��G��H���-
�F� �U����z�-�5	B�ВR��e%�;�LU�Z��`Ah�*���%��K���H�cRHq>]0���F�D,c ���7�r'0c�@A`@���Ӂz2%Z!!d1VV$k�aBq$���gf��M"�]��M&�0k�#��9�F!!!�m�F��Ʋ���$)�kZ��!e0�e��\̗Q�)���0�IS�@�Bd%�'q�aL6B};��?2�������#6�K!�,��;G�}�>����.����c9��n�Mа�0�t��&1���g3�W�M�����N�S�G7�A�H[��b�Z��HT�oD�VK��!a�k�0�k�pD�6��5�*Bo::���d��
T�I���,L�I,R��m^�a�u��Аb����X֘Ί|�L�ѹLA�艞��X`H1bĉ$ BNJŬJw���sَ|o7�]�Ɖ��K�L��ҙIqu=�Ld�t�!pc&���4�R��d��.��bkX��ak���tO^�_}��K�;�/����  m� @    ���`  ' 8 [@                    	$ �                                 ��    ��  � H   o�     d��ۃj�-��m�,���(�U�P �kj(��2�Ji��Vx盔��bI�Kh�޹w�Ѵ���$���&E�i�c��	����6��*
�Wks��]���1�mf��b�EuT�v릫�f+����V��)�P�&���2bh��4(�QmU�&�<��7����/&��UR^��q$��e�����F��v���l3�d���۲� 5���@U���U*��$�`�` �x�B�X]��y���v�s��r�3n�K���"���4����U$�&�I6 �6���m���� $����p��6ؐ �mH �` �[[kn$8���Ӏ��it��M)���X��ڡ�= jGm��ݶ��,�+I��*� -�Y�ګ��+m���}/�[m�յ��]@mPJ��JK.�H  p�^�m�-�l� �'i$�����O+m.�b�*��5A�m��k%��p6���}���UWJ�PR���ݮ/3m�� m�%�($ 	   ��� �v˦���6Z���-�m{J�5�-ɶ�%�!�-]N�VڕjKv�"7nj�H6�[m�l Tݲ6m���VWf�p�c�� Ol�A���#\evU���/<�p�_UW�v���(��=SGY�wm��a�Y���T��P�ZĪ�R�P�d[������h��.Ͱe
�:ڡ]a�ĺ*��l�ȣ������.�ma.^5Ip1���B��Zr�buK8��-I��n�	����Gq����Aӷn�:\1��X��1�&��6a[WL��;z;�	�T�f���l�f���X  l�PT��a��Z�0�;m�[r`�WV�[*ި�s�V
�3��4Q�n�^Z���ٝ�"W�lzU�i�it�mH�W$L�+�)�{�wY��X&!��2j�m�❠��9�H�Nnܝm1�;��J���7BEGd��K�fc	�geH��X#��m�F�N9R�ɵmr�W(�t�S`Y-ۍ��E ���m�0m
�2��C�!��
���g��8ݤ��	Ѷ��� pO	�U��[e%�tT�l� �[N۷Z��z��a^�W��]k����U��L@@PU*����Ö 6�[N/Z �m�Hm�����E��jX����uma�*鍆.��{5U��u���L(l�*i�@�1�U�Bۊ���vV��gj׶�Ln��#0V��0R:������Έ۴/U�ua۶3hw2\��i�sQ�F�� ��bݮ2����ʣ�E[p��+ƸN '[PH 6�	�ԃ[:1�v� �	-��l͵)��$%��5���XRÖ���l,sy���I[F��8�Usp�lԪQl�U+��;s�X��)W�Ɯk����QF��J�.�×�hT� ���UܨJ�mU7j�@^�v��x�A�/-m��[J�S�>�~_�P��j�m��O/'�	�m���V�Z�  ٮ��\rt!v�6�.^zɮն�
�V7jt� [v�m�-3��J��m��P�K����l���_���T��&�f�Z��J�A�6��2��X�msj�e���UU*��R�˽v(�$i6�`���`ڧM�$@�� 1}�����;*�UWU*����L�YMي)wkG*�wE8� Im8d��bݶ�m���M���qd�	-���W���n�
�`�]���J�İ\{ \gt�`��A�i:�*k�ɸ�0�j���chzZ���3gh%��9��t=\x�Z�P��zU�������R�	�㷌<����jڜ�e�uٺ'9Y��`�FLOQ�гm�"���+W8�w]@=�OUmV�@1^��k"��uQ�fu�	)]MQ�T��]n�Pyn��dѫm*S)0��[�@8��m�[%m&�+��ؑ��ƮUt!�������ں�^Uj\:�� �6�v������M���`[%�ր�h״�h-�p�m{md��H6�l�l�m�ڶ�A��Lؽ+lYfA �6�$�<�I�vƮi[&�p� I -�k�h �k��pp�m���f�j�[Ul�t��k6�4[hnBI��w6�ZL�$�l ��Hګm�H K��p�^��$gJ\ m	 �m�ؽh�b��`����@�m���8���)yf� <�,�d`	-��6���ޛ]$��̀�v�m��`p	�[��-��i$[}�u�bH    �8 pn�fU�Bj��T
�V^[��EP� �
KUWG5QlaS�����%��k`+j�l����֯�$�$�p,� ��*�^Wvxi�	؋�U����h���(�e��l�6��ʫs�媭�.��V��p�y�۲ꚛ�*\s�h
��Ű�r!�64ݣ[���@�4�ۑ&<�;Um�sS��v#�Μ{]T���iz�����m�)2���W�q�����q�#5p����ڨ�z��Z��N2+��n�X��۶��ր�%�mm�Rv�����Z���U�@p<+eg4�G�Y@6��7l�L v���mmR�����;8�UU+.�[r�*����HXt�	�%�6�9�m�a8yP�+��ft+Ul��q�f���LNۘ�۰��8m�mNʲ�t����Y8K{[[d��� ���%�S�����] q�f�m���X
�Z��m��h,0�J�Y3K�[(hkeY�v�T�6�(�
\5*�A�b����K�r�.��s���M�n p�[l6�ާ8A�K��[[m���lm��t� H�[v۰�  �kN8)x����)TU������ulY-�ݫm���y�л*�Uj�X&�ݶu�%��!���I�*�PM\[P�+���򪪭UUUh[n0g���pp�jLHKu�m�L)n�V�h�dF�-�9J8	*�t��X�z� �`�t����V�6�A*Ե���iK�T,e��O��b�t�
��Rt@;I���v[mڮ�eZ�
���Jˌm�7<��J�l7R������n�(��O4��Uf���VI`;jڲ67#[���v��am�6�����٪�����]��;v*X K( kXA��q���6�`-��X��VM��U����M�m�m�K:��h�c\읤�������`-�[�4\��Lq�YF���D�ݴ� ��l�m*��� 6�-�ݵ����\�k[h�l��JW�2�īV�mUWT��rH	�P嫪�%Z �oY�m�j�	J��8�i�e���h�> ��$�����3uآ�k*��H穵T�\�6��̇lUPJ�lm��6���b��[�̃n�m� qU*�V�2�+=���vU��  mK@�0�z��֤�$ 8 ����  �h;�	�� �.�kn K(�%�	m�i 9��m�m�nuZ�:����� -�Y@q��`hN�l mJ�Z�����l�l�C�����$�}!�8P�YKm�̖H�;` $I��k�큶Ɛ�+R:*���^j�]�8���jD�ɭ6�u������ X`�a����m�nݗ��(
��P*U�H�`�[O,�@�C������.�X����n��K)6ܲ�����Zݺ��^ ����L�6���n�m�[@l ��[V\��&�r@HR���Ѷ�[���p5�yI6�h�۴�ưR�`��텫��u��L]�Mfv$-���;aA��-��Ci$� �� v��z�h9$� m6`Z淭�,Zl�ջ�� 6�ӡC`m��ͮ��Z@H*��,qUR�em:�$tه6�h�`m���j�x&R$z:�`Iê�`-�Z��m�[M�n�I�i6���m mp �� �:�*6�����>�z��['P�I��n�  	�l���Վm�f�m��iol�m8[h
�Ge��R^W��9�r�ض�  ��y��ٵ��7e�
[h   ڶ�6� ��ۭր[iՐI���lq�����`�*L�` 
�vUT9iVU�vP�A��l�` m��h �m�! ��6� �� 1�$t�m�<��m�d�3e�:�� (@  ��[v�յ cZ8�e���K��m�  ��6�  $�"�6�U�L���;��.����m��?��u^i7[N
m��ܭ,�cm�u���b��`m���A�v�4U�p� m�i6�m�h�3ԫU����\�!5�%��j�2-��Tף� ���[Nm&-�n���8�Z���j�+L��ȓ]V�h��29\�Z��I��999�ri'��O!�v�����)�O�p��:1"Ċ 	 N{B���
��8/d  �i������D0� �A���QˀG��m"�t����(��| }�Tx�TL�Qأ�M���-V��A#�Sq,pkF,B��H � �Zd^�E�&��#�`t��`x�·(�P�=S�&��d'b�@�S�k�T�QD�C:O��d��"�"qz��'#�ʙ������*|:>"t 2
�A�$�x�.� � dp�O�8�^ B1 0 +��b+�R� @�u08�Dx�U*UJ�iG@�W"`Ȁ�j����Dt�'�D�P�; 4���!:`	��Gc�E`�x�b
EU:(�`�+�������P5�	�*/EB�L�
��Q���b"�@��|��p�D> C��YU�D: � �"�(4���5�A$!� ��"ā �!B��H�dEc��|�a�� ��9�R}��=@�/@Q5�6.$d��! �"$�Ȑ�D"��2��" ����T2��N#���A�~P��NDB�dUaEB@! �BE��`@`���T���B��X�"�4���
'ȇu��P*�e��!�r]�(�L(=����B?�U��� ����V D-F�b�B�Z�����m�m��t�n    .��      ڶ�m����; �"p^.�n���i��ċ8Kg�����BH�Q����'S�m��L�G5��']�l�5&��
@J��WT4$��WB�Ӻ)72���W$YDx��w9��2�r���L�R�)b�at�p� =�0Y�4�,=�(lH���Wˮ8;1��\v���񦓦ΒW�4��)��3h��*�n�YC�e�Zܼ�&�=5ЎokdN3X:ƥ�ΰ�H9�����*���nA�	q�ڀ�8��ݧiI�1tf1N7J��1�����0�Ŋ�FU����ӆ�p@�!v����2�A���i:<c�je|���ĺ�^�a�탚�Q1�!��vUY'��q�ey�"n6�zC�D� 磮�+��v��Z�A���nК��Is�@��/����/)�pO6͞M��!�֠I^۱Y�bq��Y'9�C]F�ؐm��ƃ�èqbU5q��M��;c�Ӯ�i�/<�Ņ�r��L7gE�
�h��W�( ^̵��gF1D�pl�Q�=v9�yn�v<d彤޸�[t�b�eǕG��7d�hlا�s&S��۶��Ld+M٫�[�����W��*���A��켷�oi�s�n:ݸ��y@��;1����8�m#���v5�g��ӱ�� ;:�6(6��*k����t���vG�n3hv�C ��ل�v����b��д��|���+l����)q��h'���5�ȗ�Yv����]�d�r*���mG�ɨY���Pz��9[��Q��˰(����y��*$�3��5�p�7A�$	��bmnM��%��x��wM#�z�^�2��6��{&췭Χtf��15�]T�X�Q�e�U�p��6�����5��������vH��2�B�X�掌E@Kc��Hm�M\��˃T�^�*��@Z��/t<���CF\�f��K�6�;!��rO����w��.�A]<Q@�
mä7Eo�T������|��*��
s�/�^u1UUUT�bl�K�UYs�g���׸�m`n�Jkm�^,И�f��Vu�.mav�Yn �݌��s�n�t��Z�.(��-�ۭ]��-�ui��v��=����8�md�� ��mΥ	�@K����q��Gc���� �(�P�+�Mm`�4Y��m�,�1
l�]�u%+���,밎�۵�d�s��2c8�&s#U��2 �����1ʽ�}�;gp��g)�]ۇvL�P����y�s%-�l�A��Y�@���Ɂ$D�9�e5�NK�.��蘉bX�{�ޓq,Kļ/�qL_�Ŧ3��MD�,K���<D�K���j%�bX�{�ޓq,Kơ�*�Xr��G)��A4%n�t��Y��7I��%�bvc��MD�,K}�w��Kı;9�MD�,K9RL�g+㔎R9H�ME)�c�ɋ���5ı,M��ޓq,K���ta5ı,N���n�q,K��^�|�9H�#��T��Q7m�M7VS6�:Mı,K��ф�Kı;�빺Mı,K���j%�bS�����|r��G)�܉
��V&�maGs���-�iI���LEѺ��t
�m�-#�SY���#�kF���}���ŉ��]��n%�bX���nQ,K��{��7ı,N�wFQ,K^N�~;F+n43ƻ)�'w���K���ja�SF^��:���&w���7ı,N��FQ,K��{���7ı,O�v\SXe!6����^B���<:��%�bX���&�X�%���]��n%�bX���nQ,K����K��=Gk[��O�Jt�Jt���t�B8���'��{7I��%�bzc��MD�,K}�{t��bX�%�����.��fs7O��N�����t��bX�'f9ۄ�Kı7���I��%�bvs�0��bX�'����H:�X�vv]�ˈ[1���v�6���I���ʜ��ۀ�0،�Ŗ��9�O�X�%����5ı,M�=��n%�bX���&�X�%�I25���R9H�#�5L�¬m��&.s���Kı7���I��%�bvs�0��bX�'{�w7I��%�bvc��MD�.*b%��wV��8�snn3��3t��bX�'�}�	��%�bw��s�&�X���T7L `� T�uP33��j%�bX��{ۤ�K�S���f���Z���<:S�8�;��Ɠq,K���;p��bX�'��;t��bX�'f9ۄ�K�B�w�����X�i�Ƣ��N�!y��T/b�V	Kذ	�ذ	/c�-�s�����D4��٩��e��aW1% �դKq��<�n=gN�c�i�U�V��w�<�	/b�$���	/b�$��Kվ�I�k �\3��r���\�^�\��;/b��`������+J��`G�$��Uq.���{���;4N	�&�;�˴6��$�� �\� �\0:��U�UȄѠGB|&z+��c��u$�9(�O�,v�e+M��}.E�I��ư	/b�=\�*�D��*bhu������}P�َ�R�v�;k��t#B:(W�)i��5be]*j����Ik ��/Ur�A�_������+C��M�M[f I%�Kذ�Ȱ	/b�>�Jcum��uv��v��^ŀ}.E�I{ I%�t�EX�%Ce]�m`z��\]�{׀{�<�I-�^ŀM�U)`Z��wi��k��W8��z��{�<����ӿ�;�:OI�=<�V*��s���gjQ�^��z}��w+u[E���v��w���������]gq\�j�5..����B�n��k'5��[bu(��BU���x����f������T`ܺc
 ^6��V̶�Hx��{p�=[&�F{pn�qv��3���랸���a���ǎ;&�d�ٰN��9��� .7b�y4-�dױa���0-���I$wA)��J�6m�O�&����c>V���X5�s 3�I�s������]�U�� ����Kذ���	5� ��8'I�wi�x��`)%�k� I%�M���*ݲ줮ݵ�|���l� �Kx�ذ	����V�L��N���~�qOL���o �{�^ }P�q]��ڻltն`�[�$�� �I/ ��,���9�p���&���{O8B�ۜv�$�ܱ0�^9Э�'�'�������3��M�`�? ��{���Ix���UW�{޷�w��X��T1�U�V��^Wkª���r�2�P��{��w1�gSRI����I{7UT��j�ݤ;w�I�$��	/b�>RK��!
��Ĭm��Ur����x��,�$�f�`�'bCe��e��n���,ݿ{�����	$��=��>�.��١5c1u5�ɶ��04瑮\!�v�����E���c�0�l�i�������Io �{;z��n�i2��;�w�l��) ���x��,�$��T%�Wi+��ںj�0I-�^Ń�UEr�	B5�X��|'���u�I7�ذ����[m����ݼKذ���	/b�	$��}+E^4%Ce]�m`)%�^ŀIo ��,�tR�wQU�۱1[E�wLL\i��Ҡ�fԛ��|�㟎�q3t�H����ū|v����O\��	$��l�� �I/ 7�D���&�Ĭ�� I%�e�X��X�ذ���"�7ulwv۷�l�� ��"�6^ŀv[�7����,M�e+M����w_��	�X7e�9ʪN�Uʉ�*�p������I9�9I��Iqc*�SWm`5� �r��'����,�܋ >ؕ��T�۶���4!��nM�l=��0.�n�{�p�0��ځ�Qb;.O���vˡ�f M�o �{�nE�I���j;�m�Ut��Э��$�� ��"�$� �����B���*�+k ��"�$� ���%�X�ҪU�]�R�M[X��v[�$�� ��"��"��E��ؕ[l�&��x��s��;��,Mp�9Uӕ{�m�m�۩	�W/gOe�.-'[�� ��U�`�l�#��M�a�kl����w:jk��F9��n���!�)$�V#XNs�9��Ě�8�W�e[#���S0�Xo痯��"d{v1[�����f	�0f�Kj���N�\�J�ۭ���E�.����b���;Do���GqfCk��A��|&���5�,LWc���Dӳ�T�3��a1m�d��P��3v�c�,��f�㱂!4�pGj�A�r�9���%�77n�ı�Lm���i���������{�}ۑ`^ŀM���	�TYO��&Ӳ����>�Ȱ	5� �{�^ŀw���V�`ڧWV���$�m�w��%�\��;��,.�"A�ZvZj�l�&��x��`v�X��}�v���m��]�1+n�	/b�>�Ȱ	5� �{�?�����E��R��m���\��i��>z��{�).n۫N�XF���G4`֋U�V��nE�I������s��|�޹�waU꼫V�Hwi5m`k�փ�q�#�������"�>�Ȱ{DH��QWwJҫm�7e�Kذ�r,Mp�;4w�"�e�˻�ݼKذ�r,Mp�	�-�����-&��J�m`v�X�^�� zO[�$�� �s��U��.�6�t��cr̸%��e�8�����9E���g�N�@�CnQzS�V�WM�uuj����v[�$�� ��"�"�$e�e����� ���%�Xݹ&�g��H��k��[t�]+|t+v�z��nK��ʼ����C(@��IUzh~��Y�{�΃����~H��C���:&���R8dLʱLHpu��!\��n# I$:�@��(R�6�0fI'> DS�A(��G:&�`d����"�\�D��	>3�!���oY��M�+���c		I�.1�Fu:�bߓ� Q�c.�$�﮴ˡ4I!��R�8��z���|�2� ��RWqK6���.�C�F�3�x&�5�l7u�!p�Cjp:�	�H���A�Wx��g9�f@O��
 ��F��@�&��T ~4�j#�q1$!���`)��;��|7�l�(��A�w�k�B��`�`�`�~�}��A�lll}��}nfKa�����w��g޺w{=�Ѓ� � � � �w��t �66
��������pA�rNp����默3�.�'V�}�y`���=o�=�Xݹ��W�����[��3r� s,�)\
]N�[��|i�ݴ�.x�н�x�+�h��?{߭�/b�>�ȿs��<���ii�p	����>���|�$�i���,z� M�o=�URD���Yi7n�V�k �߼���`ݖ���`��X�N�T����X�s�RI�s�Τ��9۩2y|���� � m
�08�Pl��><��sq�}u$��l�s����ˡ�� M�o ���<��wo�X����|����q��Gh�Q����=TD0i��J��Ւ�H�d���&�7dD��t�]+|t"��7ױ`ۑ`/b�	�ǀoMJx�	�ʻJ��7�"�$�� &�%�X���ʴ�Ո�����	5� &�%�X��X��*�E[�V�[l�	�ǀI{��&�`�q���v� �wlm�^ŀz�k���{���	�ǀ}�U]���H��t�uU)�c�D�UٸH8���sA��r4:���5.J_N)�GX��%ҳ�"v�m�V����6�C��gv�D���5�F����K�0��c���q��;]�훣�6�n�'���q(g�8c�I��=V�#�>���Z���l*Q�`�S(!��s�ѽGƙ�8�Xz���.�A�}����������,�eqfn.n13��_)�T|�7��I~�.����;j���C��$��bF豅�(�Uq�݉�^�Ih����� I���c�$�� �oU�m*tڧWV���� M6<e�X��X]�D�l��-�V�o &���,{r, ٱ�wSQ�V�5WJ�����`ۑ`5� &��4QU�T$Sc*�+k ��ŀ~�+�\����V�<f������qf���M�q(����7 ��A�a�/�����f�L:�z�Y��ϏI��f��Eݤ�k�'�����/b��s��m�, �J���U��iX�0$��;�d�Vd$T؈�k�͗�`��`k�{���$w|���$��c��m�}�� ���QʤI�� =[<�	�TYO����i��6`q{\��$������"�>����VҧM�wV���wc� J�ǀwnE�N�ŀ~��+��D�tx�8�&Wd� �N��M!�A5
]$��Y�����r
k7]��U5pd�r� =[<��Ȱ	�ذ�p�=�,�n��I�J���e�� �{ݎ!���Ij�-P�M��mc7RNw�ԓ�w=����&�#C��C��B��P:�ئvr���x{r,f�R�*ҷV"��i��wc� Hlx��e�X��EE+�RwJұ�`�ǀ{��g��t~�~X���W+��XR�Ҿ��ّ��l/!(��-`��mx]�Y����N�8U!J��O+_
�m�P0��g�� �{�u��Uϐ�O<o���|.�j�LH��Kس��W*������<���*��=��5m*�mS��m�v?*lx{��K��� ��y`[@��m�;e�Vف�-���:�}�g�RN��ԟ
��)@ ��6A)j�� EQ��P��y5$��s��&3��3�x�m�w\0s��_ݏ� J��z�����m	7�!�!��]D�aaHܭ�)�(Jm%��L�1���%�ܒ���j��m�Zn��?~�~X�� �6?Ur�Aݏ�=<�i6X��I���u�?r�W9Uv���<g�� ��,�s�H;(� ��$�iX�0���}�p���U%�\��;���>�N	�I[b�wt�x�R���{�<����Uʯ�\��_������)�NջN���X��`����=������ԓw�5$��(<P��s2N��ӭ��Hd�S��hOf\�,�H��ݐ�Xó��7;�v�4��z5���;<����K�nz��Rac�j�B�;ήOe�y'6a�v[����s��5<c�ݎX��9yOv㝶{��<Tr�[A�eۚ�'f�E0�:�l�׫�N����ٻRDF2�<Z9��5�ˉǉ�&����C~}��8�x��leGB5�2N���~��N���O�h�e�Ao�H*䋹V1l0��t�;I��Ԛ-���@f�'�Ru�2E#uj�^߼�gRIJ�5�$��W�s���/����Z{~2�:��-����u�$��?�{�s��=�}���u�������h��*� wg���%#q,I%��C�IJ���������P�S�U���o}�i�$�fxϒIJ�5�!}�>��I-�T(��Wn��ա�ŉ$���>�$�Q���_wg���%#q,I%.j�B������ �jZJ�e�1����|�	^�i�6��YMCS��� <�>'I$��ϫ�JF�X�K��C�K�'��-��C)����;����ry!.�0�Jdi��7�hL��)���y��ն�s������{��ӓl�����s�ve�;��W�$�{��^�UݯW��Ē]�{�����<�ɐ�)1�:�rm�����ݶ�ϳum�s�7�o�?
g������oeO�Z�7G9;��<|�@ܟrO}��������� ���þ�S�}��_F�h����uqĥ���]trtV�nBBNt��%n�nw�k�����j������<_���E��lK����$�w�举�)�����<ϔ���N}"������?�Ē[�}_}�]�S�x����,�eE�@�_};��������@" ��TlQX�b"�`����L�=��ov��s�: ���Xy.50Gd�^�_�xx�JO{����nIv9� o�03�KZ�;1� ���;�|�^����$�����J-���$�ר����L!3v�ix{A�uP�aq��fF���t�Rݛ�B7�J�oK�`�)�]�Il�e,I%��_|�Ql�����#�=���`y��92E#�6a�	v9�$�[/)�I-�>��I.�̥��������A����'}�z{��= �y�s�ϧ$�E|�}�: <����߇�utMHg���z�M������y�{Eն߻���v�߾ l5�	���4D�A:#�??������>���8w�Kb�3��� ��y�:/�ʪ�S�߿-Ԓ��~���$�fC�K��'�
l���VNNݮ��
�08,���6��G�]��\�j�0_�9^�m�P5ūCV�u$���~_|�QIyOIṅ��rI���|�/@��}O�Ʀ)�c7{����3��c����ov��z�/@������'9�?oG�03�h�Zm�II�}_|�]������Ur����_|�^^�1�I.�Z�
�K�IK�d��Q�	������m�����<<��9'�rNE�߾�;��f~��!4R:`̽ �>xw���g߾����}�߶ov��;�V�t�>U!��k�я'�iiM���@�� M�R�m���@��|����z�Y ɡ�S	��� �x,a�9�¸��?2�)�q�Ne>;r�#+)߭��h�B(LQ����$�X#śA>`�ː�0�8X�$#	� ���J���q�jN9�&�G�dF�a1��L8s��It%˛$)��Sm��C���Iy�>7F$��}p8� nU� |G�"�!�i�����U�`�L����;���HI��20����{�{�?/�-���kx    �V�     j�qm-��NL�t��3u0gi��Eձ��ç���+[e����R��J$�#�erۈ�)�
$6����F�yj1S,R�^�3E)��;�)\�v��\�v.;XnC�g����8n8��hclRj��)�V�/�WT�fa��?�=��#Ip�5����
�K11�6J�Ch��UΡ��8Pٖ	�f��m.���F�̨Fݲ����ѯ`�ν;u��Ԗ�1.������ �t�0�)la�sp�L-@�!�k���x�Qgf%�\#��7KZĴ��-&���jv�M�D-WnQ����uٔ�s�Uѧ�M4Nv	f\��7�(�A-�2��*�D�z�Ν;��.��u"��:x�Έȝm�r�X�[����V�\h�K��5��<�K��x�r�[�,�],y�l��wmѷPcl�%�ېk.	K�2�M�jl�Qg�(�7J�U�K<F�4kjˇ<��od��[8��q�LV�5l�}ˁ|�ˀPcqU[�ۊ��M�']�C��#*��Sav��R�`��nݏ`��s�tΨ5Д#����pN^0��{�P����"s��`�&;t��m]Ͱ1�kyN�]����v�C��,��\I�������Y�6Y0�n��-3�2�9!2�)
�]XKX�G]F�F���фئ&����䮴bʫ:�c4���p��J���T�2ݍ�G75;u��!�$O'm:����h�l�bZR�X��W#�Ayxe.dt���@P#M�\�m
�j0\L���9��+�Ll�qZڇ@茎d��xֲ3(��h�:s��l�����Ge���*F`����˩ƹ���2֖Y�q���vÝ �Ht�նR��6���/_"�M�s�t�t5W!#�]�8�Z���vڭ���o+eq�b��\Ie���6��-{�BG*�fSY�mW9En��G�4�C���V��`5�pC��])�?�*��h�G��S�@ ��0�|��z�������0 �v�+J���\��kg�wI���X�B�N+c� �Q.��.�6E���Q�,����b���f��߭�S����-��S[J�5у5).\芖cDF��r�&��x�̖㎆1�s��5�{���b89pd�P>M�b棈����[�W���ͱ��i�2m&qQƶE�����Se��u��F�јJ��5��)$��G��''��98�vûM�ƅ�9��)mHf�)U 6X�r+�T�&�!t�l6�I9�[�l���7G9?|���� ~���� ������w��}����ut�Xg�lx�KvO�￹\��Wj{��1$���~_|�Ql�<�s������%���AMNg+;����K����}��rM���1�I)=��Iwy YI[�j�V��F$�U����=���%�=�x�KvO�{��1���.���<O[�$�2�5m}�IE��$��\�r���]�Il�z�@������Hy1��0���;kX��Ҩ�cY��M��<�Z�
�hL����t�6:�i�+��-{ <�޽���]ۙKIv9��?s�ʭ֒���� �|{o����He����y�:�'a�wD���Z,F)��s��dO
9�w���{�-S�ǉ$�fC���r�ԕo֓e�L�1��޾�w����j��N]ܞ�|�[/�KI)F�U�Zv˧n��䗹�U�O}cĒR{<}�Iww�C�>���Ӝ������`���蚐�E�� ��y{��I?x��;�����$�6e�Iwvp����pG<e���(g�]q��a)�,t5v31pUK�BQ?I��yo_5
[�\��������X�Kc�}�IfX�s����u���~��݀{Ϭ�S�&�3��>xw�#�b�w��έ���צ�m�s�u����y����Xh�&����/��֯V�y��{�<]��`+��:Ǵ] z���`���u�s�շ�(��}��ߦ�m��?h����罻�s�#��������V �f�[g�$�V�M$��6d��I#}�CĒ?y�^^� �?<Y�3��K��5�F�]�}]�띉�wm�ӝ�c=�wj���/���u|����8鍘v y��}�_�<�BIl�s���Ke�)bI%�<��+t�v˧n���;&!窪�Ҟ�xϒKc�#Ilr/��r�whؚ��)[㤛MbI)�g��I.똌=����y`�{�}�)%�Ut��k���0?W�UU�����O����;6e���9��$B"֍X	 DB.(�HXP$iD��� ����`^�(��i�ګ����`�"�?W�W+�����:���0��+ �֔�M��E�e��ۭ�u+�!�X���?r}�01�v&e�����I%��,4eJ�j���߲�v8`wfW���U���� ��<&�Zm��v�ـn���UUUvl�ߖ?_�� �d�g��\H����I�IZ�*Vـwc�v\�r�T�w��`y��;ڍDݫ��q�Z��r�K|��n�،v8`z��ݙ� =DD<�ӱ�[.��k ��b0��s�U{߾�t����}�>Nd�I���}��ܬUUTW���ۄǴ��l�5�6�4B��2Ԙ3����d���F$ ���ߑ����)��{`��{V��/�X�ZM�!ˇ��;=P1��s�<��@=��ct��:�f�xW���Jvŀ:a�IP�D���橣��ZL�AO/Dbu�t=�X�lu-�7o`n�N����t���;��{X�.E�{��b���3h^}:10\���N����N��\m�kb�kg�[ɸ�6]�<:6��W;��8�!�{�nM�ߤ��̋4&�
_m�������eȽ_ 鱗��z�\2Ђ�k���0��eȰ�̳ ݎ�$uo!E��:n��C��}~��>�2�=Ĥ��wc�uw��E+�BwJ�wm`z�w��Y�I�� ��e`z���� ��T�[c�;v��7c��Uʪ�͟�v���,�g����kl/��F��fW0uQl���n������3��X5�@�\��ͪ,mi:-[+l�ｕ�v\� �ٖz��	<�`���nՍSv��]��>�;ۭ("�T��{�Ϲ�MI>�s� ��eg�W9����]��W��m��X�ӷm`��e��p���%�����{�ն����:(�����վ�<��v{+ ���?r��{�l�7��I.hAM��v��ٕ�~�����;�� �0�n
��i�T�[@�tQ��&��qY�J�O���^�p,���f�{>9��;��M䵋���ng�����x�fY�l��r����mz���?Cm.��7�=�������;��t�c߿?��߲��"�r���$uyO	�V���WI[��{���vea|�PEr"��D��H�@U*B�E��ʈ}�7�'�����'Ǉ�|X�\f�e�[��䓇��}�jI�c޺�w��5'��&=���MI<�|��R.8鍙շ������rr�vg��	�?ݓ+ �U�_����߬@9n�n2���;^b)19�CFQ,1�Vkn`-��F1��������߀}��F�8`vL���r���~0���:-X�.y�Xx�}}<��:Zs�ѩ'}��jI����_�������ZSmr�v�g�e`#��U%ݏ�`�~0�g%)'M���hj�`{�J{�� ���0��Ur�U�ڈ�vpG(���5�tԓ�:"������]$ճ �����}ݙX��~�*��j%G���]:�wu���#m۷��9�;<��&�uh]ɳ.�,�cX�w�.��˶Q2���~����?�e`#�����~� ����I�tZ�*�l�>�Y�H���n��:�������9''�I����|.5]+��]��'���w��{��JO?w���	A���c�aV��f��Rݙ�0Oy�vL��8`۷-�6��J��&��#�=\����|������¨9��I-���u�T<�;&M���I��.{M'Q���;*F�N�-�v����.jme�X�2ǝfm��R	z�0ֹ�әA����V�ٜ�u��u^�x9�����T����Y�ȧ���ӧB��λ�68ݼ+F��ƋLn�y���4lv-�T�8y��f"�A��l�=9���p�u�n���[��i�cj�	V�K6�L8��U��99�'9��m	7z!�!360����YH�Z.��vܬ�<��pt����ܜ�Մ��9��������oc�����{� ݵ�E��t��]�����3�\���~?�@{߿<}=�������"������]$ճ ��� 7dx~�W�Oe`�>ޭ��߷���1Kc3z��N@�{� �Oe`���W+�9ʿO�~0���?�5��5�S+����������g����� 7dx�b6躖�bb`�H�b-�SAص�n�Wm��t�: ��%:�v�]X�]����}����#�W*����V z�T=z+Bl�����޾�}�=$�:C�F�5Z�*�\E;A�+��׀OOe`��=�s��$����n�*�|t�f'���vl���Us��Lc����ԓ����RM�-��1�KM��v۬�fV�r,e�X�s��qI�}X�UR�Uۦ����n�ˑ`�Us���<�O{+ ٳ+ �y����)�CX6��V�HI;u�6�>@��k|�n�5�I�s����{�N������ZWI;��z��&V�fW�s���ܓ���[����=�Ce�[4m`�e`6e`�"�6^ş���S�����_��Ò��3�o�{�S�'��{u0l �1K ���˗z�"�D�3��2b|�U*����t�v�B<7�LT�����tI�$�
���!S�Y�2�D�ݩ3�18c�D�$c,d4B#!!#>n�l	B�'����80đ)�i$RTC���$�4MŀG,��M���h��c�DB/��:.����lL�B����i���J�`��4�0���@L*�T�ʘT>>�~ �A2 Q��@��_�D6�0(�܎���t~C�����+�v���6Oe`�*KjՎ��;�]���r��{��X�s� �L�M�X�Di.鶂��uv�KذUr��{�W�{��X�"�?Wg�5��
�`���R����y-Q��=\v �	5�ٓ0t��$���sb��v���]���`l��>�"���~�rI������V�����6ԄT�ʳ�6e`\� �{$�Y�W9�$M�U,�����]�����_����j~��&1����5$��g�ԓ�,m����t��kܮUW�X��e`�g�Rl����]�ԓ��.$�]�e��16�	$��=�W*�=3��{��,Kذ���K�Ɏ����u���dj,�G��:��hf@�"����wwt�y�KZl�3���?�%Ȱ	/b�r�\����e`ڳ޷J���;�wB�u�Ir,Kذ	$��$ٕ��s��$�z�=wM�v�$�޹�n����\�W���w��, ���Sn�*M��X���ʮr��������� �\� ��,��I,*�QM���X��{�'��}w$���]I7�wF���@@�`C�s*�PC	�0�rZ��}$�0�i�톝3k�m(�����z:̸8��F{Fe��u��ݬT�G1Bgka	p%���ny�i��7L��{V��iVh�hMfx0гe��b��i�J��k̑2�W/hʐ��2��i|֚��7G]���v<�r�N���Ζ�
qI���)�;3���A�W����t`��;%�v��ٽdטf�Chƣnuٶ�'>�w$�w�ہ9bje�0�n��]u�`�]��W��u��آ�t��q����7۠>3t�Z���� ����0�\0��}*R8���]�WI;�����RGd~0	<�`m�Yꪤ���䚫��n$;f��v8a�9\�W{�?������;�e:�t�I]�l�$���Kذ=��3��ǭ�wn��;�[f���������`k� lԬ�(wj۱�kE�oF6N;U��z|�x�II����l;E�xT����+Ce�'�{�����~�����vG� =��7lct�R���c9��o��f�`@8	u�Ϊ�2 c�y�}�g�RN{��ԓ��"�>ݔ�|T�\�ݳ �\0�\0�W��y`���":Q��[eڰ��0;^�ٞ��,�ތ')I���*�~�J�R�I�f%�Xۮ��}��wb)b�K�f�u`k5���,49z�.XNu��{=76�.H�ƶ��gt	6�p�DS�;#�I�ۮ��{�<��+�N��i��؁6`k���%�Xۮ�${ы�ݎӻ�wN�X�f��w��ԓ��;uAL�J�hUF��Q�����R����W����~0	��`�۵d���-�I[0	/b�>�p�$�UqvL��_��6�������>�p�=\�W�=�|d~0	/b�/���~�ƅ>-`i�ص�B�MFQbm���������%ف�*�l�(�fkbYtZ��$�Xۮ��~���W+���� ��xI~�iX]�V� �G�s��H��y`G� �fV�j"�'ڥt��k ��,w\0�W9\Kޞ��;������H�v�,tVJf�7R~�
8����RO߽�F���;۩2֊��ELN纺�s��u�����+�*I� �fV��s�����{�<��p�>ة��Q+um�.�*��mF��	���l�[&�]�c=�wj�������3�����t.�������}�b�7u��s� �����%��yX�Ae�I]��I{{�U��ʻ=�?���~�um���_Nr}�ͭ����V(�h<�6��y�0��X��X��X�eZXR�tmr�ݳ��.�������n�Ł�����_���C�/ȶ�J���X��X���	'��$�{��DC�c� 0A�DZ�`D�R"���a�Z·m�6�g6]�.5�� y�Z�,����� �.1Ml�֪	��/7N���b��8�Um���n���E�\��p�*tc��Z��m��1]^Tm�qmWe�(�WKt�u����s�9�yۍ/G��n�n����\l<BX�Y�+�N��bR���(���ŕ!��Y�Eab^{..ח���0�M��� � ��NI=��S�y��Ϋ�j8ׅ�h��
�Vụ̈́�֡�@��ɍf��=~w}�k�|�)��,�	��~X�̬�&V���
wi��E:T�k �ٕ������w��,v�,�ڋ)�WM4��%n���X�8`��`�2���Ne���;�Wn��p�7ob�7ve`z�U�r�}�}X�]�y1���n�V�v�,wfV��x�z��?�����"���/<k��<sA�6�th��"�r��l�k�USiӫ��v6��I=��}#���s����<�	��iaJ����wyɩ&���kl`Ⱥ�BB�D�� ����&�5�g��r,wfV�@Q]��Yh�i� �Gv�,=II=��w�~0�D�$媻���M[0�ذݙX�8`K�`)���v�,tS�M6�ݙX�8`K�`��`?�em��q��V \��-�s�b���6�3�;O\ >�`��:�m�H�+���P�����X��X�̬�!u��V;�N骵m���X��X�̬�0n���V�5V�%v��{��+r��W
�8W��$'�x.�q��jI���, ��l�n�N�]'˱��ݙX�8`K�`yH�6z�,)R���i]� �G���{����=���f�{�-��$�f$R�z�α�cV���CoiA��œ���gǭG=���U���>v��n�ŀw�� �G�F�!8�]�J�'v��{���0��X�lh)ݫum:T�k �c��~�%�~��$��vC��M�LJ�[f�+��{^��s�������q�)�:o@�
�B*U�Uj�	��|�|�;�����>����a�WF�r�������\�?{��	??�;<����M�]�g��n�h��y����6�|����q���	�i�@�mcp+F�n�]��E�/ �c�;=�s����� W|����n�*W˶����&�'�C���?����=��I��w�D�괫J���������Ň�s�������?��[B��躱�l��UKu�,�O^�c��r��}��o��BO֩ݔ��wm`�e�v8`H�w��`s���
�0B	Ge� l޵���a�8/4&`�C��ʉ�"���Ć�&��r��s�;��M}���֐��^�4�$��pb1,E��'�`�Y! ;�o�MBqiB@ddZK�	)�)����&2I$3�_��b��hekI���D��M�� Ԏ�Bp`�E$%�5�>�R[b�p��_���o"ci���4����L�$��q�d!	�C����'�?�[j
���Њ�   -�      m�a"�[����(�WRI�ŵ�(�d�ΣY$��u�t�:k�n��j��^X\A1Ʀ�^l�荇��A�p�`���udV)cR��Ó�6�:ҩq����K��6���=2���0�΍��@�h
�7Bf7%���';�Ya5rcl仫��eB�Ɣ�Ũ���f�4h�K)%+ۦ���y��!v7�Z.�t�(�I�x�T��
��\K�Qa%���Uu�.-�`l�>�8qVw<˗�)r38��ĵ�C�O�E�a�`t�qø�r9����E�^A�n۬��&p���4��`n�t���#�| �u/<T�u!/.�**�V!B��m�i��9�;y3�d��iI�m�jV��Sx��O-����q׶��b|F����͔-��a]r9zɩ�j}v�ѬÁ�eB�����Ś2�1 �a6�%���-j��ֺ�J�d��@u�\�T������SR\���v��W��l��n�:�3Ve��.��WnjV;i�Gms�u�z�Z�1�h��x�4i����h�N��`�@�ld�������aM��a�=�:���1���,�W�u��W���;\U9��t;ʁ�9�5TmBw9yiQ��U�MA��(�,��|u<z���Sm�Q����XA��X�j6��n����C����j3(�\�;�%�`@Ҙ$�b��9�:5����6MZLb�m���u/F�V%���G��K�e���]�U"�� y�C[]�j뺓#鱎V���������j����RM]����LެgE��lK�V���@msݫ��p��F��j��Q�kP����Z')v�M`�f9�u�vy��kۤ@��9"��Α�bNc%�%��Up,JJ����<��6���j�7!���:X6�N�d�2C��&��˛Uml�\hm�ٯf7du%X�v�U[X୍�{���"8Q��E��D2� �R
pP� 4�M��A����P2m*؜��~c{����ݵ�,�1]��h�N�J��V����,o4���� ��M�u����aF�}�֞;��Q�ժP�lV6�E�;>��{M��ױ�rd�l��4[<�)��n��V6ۣ�n��n07jr��%�ǅ�G�}�^{DG�j��\��l��&���m�]IY�G\�ݹSb��t�h�9�@�i.�MB���ԛ��[��{��v����E��RV%ݷf'sێ�44��5�Zn�ff��K�w�>x��b�FX+����� �G�����v����x�x��۫LV���l�>�� �ob�ݏ�o�>^���>����O��n��tI�� ���`�ǀ}��}#� C�eE`�@�n�]��䤞xw������ Wb��[�N��[i��}��}#���ŀ���I�$���m��a͍��!e�l�ѭY�q�:�CO5#��]�)-~�f	�!��S�+�t���0��, ���r�_ ����=[j��v�Ut]X5l�;�س@�@�O��&���RN���ԓ}�{5�m7�J�'�T��WI;�����v8a�����?��,�%�
N�-�E] m�ܪ���x�;�?{{�r���y����mؙv���l�>�e`�*�\��I�}��mn)�q��͏b�Q�-�D���3�6 ��y۞�L�>Ѡ苌Q%�̂�v�ѳ\� �ob�ݏ ����+�9U]��߿e`�'����ۢ��.��ݏ?P��Ϲ��jI����}�9ۯ�6�}����lh/����;�~0��XU F����8��q��I'9���>�}�ki�Њ���<�I��^�����I~��wc�>�p�%v�-��]V7X{{�R�y�w����+ �ةQwv�%um+��t��,�kn3�.�̴ls�w���z�V�&��R�Iڥt��k 7v<���&V��ŀ�����n�`����0��X{{�v^~H��Ci�e�n�� �����U%����� �JT�Se�j�]���9�[�y`I��>�p��5H�Ev��L���[Q$IHI[�������1�{M�;�C�g&Jb�˶�[���0��X{{�9���B_v��5�Pd���Z,D�]k*�a5�Q A;s-�x��]<"Pޙ�+⶛������>�e`��X��x�eZH��,���1]� �I�����F��,>�8�Rz�v�-�PWc�ՃV� �ob�5n��>�p�>�e`�m!�Hwt��wm`�e�v8`I2���, �M�����ݢ�Pۼ���&V߱��I9y��RL/ ��� @����v��򪪪��X 
�@�pKf�ѹ��ka��i9^`�����D�0��#��.���Z!Z���e��,MS(����0Փ.��X-Ƥ�Q�3�}�қoj�<����fJ`��ݸ�5�E��8��W�=���#;�r��UøV�k"���e������L�+v���{K�i�,�<[�5�ˋ�Ӯ'#��9h`g3l�GGq��V���NI��Ǿ3�6⍱t��N6��:p7���c\���{4#`l�S]JP��2	�]wm�{&V��ŀ��c�ߞGK�c�h:&6gV����ïy'8$��;�~0�p�r���H=F�+��Iӥj��[X$��>�pü�]����� +�V���и]��}�L����� 7v<{��%j���.��ـ}#���ŀ������>}�BZM��75Vmj8�xp��t��;l�o���z����dn���.uWu`�g�n���ݏ ��e~�|����o����Hwt��wm`��u�~�D��Ը�tjI��=��}��Y��A�J
��r��4��� ���X�8`��X��x�-:t�i���u�}#���ŀjݗ�}�2���tJt�;�N骵m�{{�v^�d��>�� >����	��6�K���ݦ�pޟf��M�&��J۵����vR���.�N}����ɕ�}#��*�A�s� ;E�g��� ��[{��Χ_I _�}}��s� ջ/=\���*��O~�B����.����7����;�ذ9_�꣇*U�)F��( bT"X��Q ��e!�P�~��׀ow�X��[J�����0?Uqn��O<�ɕ�}#��F�R��wJ�'v� n�x���{�������ŀM�T��b��t����&^�|
�痮���{��`^�Vmp�t.6#j0)�պ�3C.������������U_ $�x��N���ʻM��۬�3�W9č۞X$�շ��<�u�I&���GK�SWh:$��0	/ߖ n�xݎ�8`�v�K�$�ҵIX��r�)'����jI��=���C�1HDb�^#��g���S��n2���ZJ�j��>�Ȱ�����ߎ�%�������Ы`�;.�wwb*�c�Q3�kf���r1�;$�ݷ=N�vJ�:�܀�T��ƒ����w�"�5l��}ۑ`���P�v>]V[0�\0[%��Ȱ�៪���F�%�]���M[0��x{r,<�����~����-Qw9wv��t]��;ۑ`�� �nE��Us�\�� �^�t�]���v���ˑ`�~�?~]�߿^�܋ ���J+�Q\�1HP �ĉ�0BƢ@?  �SX0C���$f  �dk�k�e��;)eأ����&ڵb�gX�� ٔ�S6T�0�	a�M`��Km[\!�S�v��\��z9�ϗl�n�5w78�-+�@!
[j�h0��8�t��Q�o]�y0��n�/M�qɧ��(�ع^��v���e�jҕ�C�.0�W�]��#���nj�FfZ�X�v��y�ɧ5+y�%�g�훎����6�'99�'	�$��?�_�,4�V�ua�nN��:�l�6���u��Sp�n����l���7Aں6k���E�j�/ �ob����� �l�^�cC��RUj��5l���7o�X����܋ 7���V�SlN��6���܋ ����[%��*�j��v��V��0���[%���X����)]��EՂM� }�ղ^�܋ ��/ ��
�+�c��+p�0.�v�xD��7k���^~��ė��t&�ŌаP�)
��uOz���XV�x����E�k��ml�;�>o}�}��?��d$��o*�Us��U���׷�v<�d��I��=ف6�0.��շ���;ݏ ��/ ��"�$�N��wwm�Um�x��xV�x{r,r�m�z�Q��/[-�B.��:�K�=\�*�[��_���� �s��߽
COH��з�.h˪�lE�v,�wU��t��/`�6���k~4t��4��6��@��~Xv�X���UU|�T�� ��U��e�\*��Xv�Y� ����{׀w�"�%-F�*Wc�Ձm� �dxݑ�9����x'�!�$��F D�h���X�#H�������6衂�#1!  B,#!L��5P�	@�B�����P�n��6eQ�R���H0��,X\p�H�0BX"�`�ljF @H�$� ��
(����GP Ñ6�.�$��0R�.m!i)�(A��B�
�1�H(��U�(��94��Xh��B	eXI�60�P�2ahT�)
H
Q�B4 B+hD�ƒ��,���P"Q(����% 4R3A����E����+�[��!E> �3�~>���(8����a�p�̴l�����F�u�
��/�U
8��M|
��M�)��v��T�2�t��˹��>�Ȱ�mP�-�mR�C�o�R���s� �nE�vG�t�,V+�i&��6���X��Uw�� n�� ݹ��&R�H�M�]u���9�����RG,��ާ�����݂��PQ3l�`\g'V��<|�[N�G�n�����<�z?5t�]�V�ն`we��Uq"K�X�����H%Z��m%h*v��y��;ۑ`G �dx�U���؝��l��*�u�� ���`I���u'TCH@� P�T"�)⊲#��6�����RN�Θ��e�qUۦRv��8`{���� ��e`���Q�U�~e���X��ɴ�$B"be�F��/��?fx�b�qnN��{<v����c�M|��3�������>�0�&V�0�mRN	�mR�C�o ݎ��$w}�}�� ;ݏ?�UIa(�ZW�4����V��������s�č��I~��7u���ZM�۶����ǀn܋�+�Ur�{3��~����P�t�]�V�ն`{���R?y|���$�w��ԓ�k�D�AN�)"����F	!Q,���'���9V�UU�tf�{N.�ӌn��&i��;�phy��im�ֹl7�1��g�]���iP���r��x�x�^o<�Z�M��[*�ɪ���;��=���P��w&��*[���̭Xm�b0��T�l8`궳3˼�T��{�W4l0W�7n�"³���Pu�gU����5tE����1k��s&\n%��h��'��tzt�I���qKv0�!5�\�t�f�a�5��\�3zݹ3���(tc�����' K��[j�h*vށ��~X{{�?W���K�V��e����m`v�,�8`����ȳ��9U_��Uɵ��~���f�&�iL�[|���մ��<?W+�l�y`۞X�ՠ�.�u`]X5l���s�T�vy�/�Xݽ� ���6�'�ۺWHwm�ۑ`����V���t	���`{��_�_7�fJ��+U�Сm"����&6%tj[���4n˺��v15��^��e�0�0����������~0	#K���b��wv�0���RrP�!.)��C
t9Y��9����g�� �G� ��� ��ut�]�V���0����ᇪ�.}�� %j�*;�t4��o���w���;#��U%�<���/5m�6��*i� ��e`���x�vy��"�7n*��VT��g�5�9F�od�.%��G�i��.������4�Q�i�L��c�J���}a��ǀn܋ ��2���D�һYEՀ�0���Ȱ�{�3�F���/e+�n�]$+k ��ԓ�w=��>f�@�j%�R�U6�p�&�ŀt�*��LB�Wv]��g�����wnE���JI�0{�/+tRM��n�� �G��+c���I��0r��^���q��&YM�1�[�RaL�S�H���G���L���Ѳ��#�o��}�s�-rr��z�~X�`��}#� J�ڸ�t�5N����n�ݹ���r, �V�e��m7N�;l�;��`lp�ԗe�� �~��>�ʱ���*�|bM��0�互}�w�Rmi�b�4�(��%�0q+))	E�~U9�g��W��cY�ԓe������ueV6`mȰ�Ȱ��Xv8`�9�r���J�WJ�]][-�I���A��&�Kl5���muź3�svWE97	�c���WI
����,�{ݎ�+� �y`a(�*��1
�]ح��{ݎ�r,�r,���W'�~��)����`ڶ�=���m��~��{� ���,d
�C�tһn�U�l�>ۑ`ۑ`�ذ�p�	Z���j�*��Xv�Xv�]I>�s٩&����I� VF,$:�{m�ꪪ��M�����i��@z#y�lvk&@�`��ٍȨm�M�:ŸH�![��mpv.���[j��`�����v���m���:�J��6\���8 M�=��U'@�ngu�n�73��+�ֶ̜�s�8.Mnm�\���Ly����D3�4VW�n!ec
����ՙ�0�-J�&]
�%2��k+��Q�������a�%��-)�\Q��ihr�.�{Q����8�����n�z��w���bn��iSvց�_���p�>ۑ`ۑ`��J���˥o�I��wc��܋ �܋ ��ş���DD"�WV�`�������wnE����˞X�?��!+��+��m`z�U\�W��ߖ=���;�� �nE�i�q*��b���[Xv�,�0��Xv�X�B�u��um�O'���}�%ǯ"s�sΔ���g���mڶ^= ����`���m|�?�r,�r,�{�PL���b��*�o3RM���E_�ؚ��q��� �� ��l�ۦ��Ңն��Ȱ��X{�K}�� �y`�Z�VӷM�M�*n���-�y`�?�r,Q�r,v*R����*�|bM��8`mȰۑ`�ذ�{����b�����[�B�S!�.�Q���}�֐gm�5a��,��G�;<�m��~��7nE�n��0��!K�7t����n܋ ���8`K�`�6���b���[X�`����V�]�UUu\���!�b�S(�A�AGB�6��)�@��C��sX��m�� �1B��`��n���ʥ��� ��Xv�X��X�@�67V+n��Vـ}��{�Og�ˠI~���p�Q���i$��e�)��AbP�uu�^o�=h�ݒV�pa��`��Ң�l�;�"�;�ذ�p�r�A����~�cv��T�Ҧ����?UU$l��w|�`ۑu�''�=�=�uVnf6�[y��}�p��s�Ķ_����, �(6�����
�l�>�`ۑ`v��Rlveݰ�C�Q1�Cc��R��� ��׮��ҺI�fݹ�ob�;�� ���M��JU�����/cs�Lp�4�E�љ�H�;	n�`^�:��&Ғ���5aLM�2um���,�0���9ʪ�����z��$�1U�ݵ�~��g����� �܋ ���g�W+�ޠ~t�-[�J�[fݏ�ݹ�ob�;�� %�t�5N�+fݹ�ob�;���r�W*�{�� x���m:��7t��k ���`��}�rjI�1��I=���C� C�%X�va	3
�	,b��%��9�qz"�8iIk?d�c\��C�-���"��h_���42�H�T4:͇zԧ����@�1�2 �"H�XTLq#2���dHaE�u �����$*�3 HH, 1$9�8���o1�E�T�c��!!&~C�!E��79#�jM@�"��g[J2̦H=�1H'�!�ؘ���\2��!$&Ϝ�FHB@� D�@!H��l�p	��b�`E���F2�T��@:��!})�@Ѷ	0�cXM7J���9�"5"|}�쳟
p�2 �A��>��)�h'��0�8cO���`&r/�X"��~�m��9�rH�@   �      -6-�m:a��nК��!C"��emB8�֩%	Has�I��r�[�M���[l��v�x��iU@�#5.x�&J��]� �*�cj 1�j-�G�oP=��H(Z����r"�Ł1��<���-` %$��:�V�kR�V�Mp͋A�@�)��ܲ��Q�	-c�����%)-¦3�h�������v��˷q�
h�+��i���91�6��n��<�#���]tr�W۝t��'W�Ȇ�#b-�b�9wXV�utdY�8� �]v�7>`5�ú��\瓮S����P)�p�gP�ɹ�r�4����m��
��X�Nz��%ƅ��&������ч�6z;�%�Vh�(үUN�U"b�A�:/5��i�*��!�{��!�
�� �Gcu-�e�Ƹ�Y�7n�n�i;RK׶��E�׫��Z9���������*�狍s���r�˞�f7g0��T��8M��Q�[pS��$ĄFݗh���k�j	�4y��]e�
p�f����[���I�&�Mq`��m��b昣�R�#��=�q��O]�-vK���7Xs��\�ѴԵ��z��u�Cu�:�ծn�6� �XjNg�I�c�U�Gu����fY�/���i��πîxz �jp��m`0�Co�/������]�Qt��6��(��-�ͳu���m&w[C`]�*�@�ʸ��6"$4mmiH����%��i�9s�]�c����V���UÕFMb��"լ��n�u�T6{)�@����*˳Uj��F뒐$�g4`��p-����[v��:�U�Wʙ�Q�̐�����Z33v]دmWBv-�!�s÷f��k���jdn��ճ������4�7SO�u�>�mU�F�Uf�
Bm�4d��@WJ���K@uT��};�W�H��m���$Y��YH�ҭ)u����v�ڬ�+�����J�� <AaD�?W����'8��/ʎ�(
�H � ��@��A" 
�	�4����*h��������?�������m����ɲ��'V^7K�=�n�������乳�R��sj��Q��B<��tc���8����N�2���WuC�'\���Y�����6@��-�QکAe�.-�f�A�S�Y6/ ���lj����YK�GE�噣R�:��뮸1ڤ)ٜf��v�Xp�r$����������V��GZ�@�R��CF��'I<��4'�Ts�pLi���e3��jɴ{��<l��v�VL�mZ�yBsj犮��j����r/r�Aݹ�D@%y][��T$ـ}�p�;�"�>��Xv8g�����5�:v��5l�6_���k�ݎݎ��Eݩe!Z��������t�� ��� ��� �܋ �֥մ
�ab�I�� �����r,��vEM*%�����ދ�)�	�f�� gJ3n��t��c=�wj0�n���y����-��>������"�>�{��|�g�� �Ig�WM��I�q��'��{u����UPô�gr�c���o��f������ԐCg��m�Vڦ�6��;��,�ݎv�,T�K/�����M��۳+ ��Ł�)����=�WI�M�l�>ݙX�Uls��&���>��{������+�c��{>V��'��c^�]6r����a9�aJʏ%GP�y��������h\ۭ߯���7��`lp��+� ���Ԕ���׸�+Uwbm`�\0�8`n̬�{~�RG��մ
�ab�I�� ���}�2��\9\��NG �D�5UA)�s����#��h-:o�[�J�[fꪪ]��V���5�����/}��� z�z�ū���:T[V� ��ŀoMp�>��}�2��ąWmQ�<t��ny�&,F��,0�P��p�[s��P�C0�D�'v���*����b���H�`lp�>ݙ_��.y`����u|Uv��&����9Uʮ$vOe`.y`��,�U��%m��J��)�j��0���{�/b�>��wu$�1J�t�B�n���Y$���ԓ|�{5'¸����f����^�*�.�SiZ�.�m`��,�۳+ ��ŀ}��)U�{���Ć]���<q��U	�h'm�n��pgݖ�H�gR�<I<��Lg��>�~�0��+ ����s���n�<�	���V*\��nS�>}����I:��<������\�) �IW�j�IZ�J�j�`.y`��,?W).�?d�V t��%V�un黥M��=\SI�0�?۳+�9\[��=R%뵉��*�|b� �c���{f��;�$�ӝΤ�2?5_:q+���ܬUUWWf�C#�ݦM�jI�!*� �/k6Z��#�a�!GCp��z�s���YU��ӹ5�53��.���"�7Y{]���	�l�AyѻOG�73O/����j�<s���3�N��c��8sێ������<�g��Ǳ�h���P��]+\<����m]	-I]ű�n%:b�K Zm#D�mђ��pf�C	tc^T+fm��wB&�@m�%�&�[5�N9ݞh.Mt�=��`~��e(��LRZّ��K�BM���e`�p���r��A��� ڕ)Rg��t�B�n��`����8`n̬ ��iR��%6����m����z�T�d�V�?�Ժ��S��ZT�f���ɕ�wu�ܪ��ٞ0	��N�b�M�m[f�d��?��&x������ܮW9ͺ�BV�`��d�fۥ&kV\j!\��,e7*��+F`5K9W�4!t���.��s>�?k��}���W>A����M��.Y�Pvg�Oﯧ���I�H�B�P��S<�w5$���V�ٕ�J����M��lg�`lp�>�Xz��=��ml~0�څ�J��)��$ـ}6e`ݙX�u� �c�ښ
���ӧh��u�wve`�rV����~0�̬���K��fŨ�
�\-���Zނ����1n83�r\.�2�q��x���������p�>��}6e`ݙX�9h`*v�b�J�l�>�ឮ$w��X��k��lІUۦح�e�Vـ}6e`ݙX:���r����1"T��AH��Z�}UU�����w�p�	F�\E�`��J�j�`~�W�{��%l~0�p�>�2��v$�؝[�n�5n���ݎ�fVݓ+ ��UwJ�򢔅ج8he�ˈV�@��̷DoYze��R�:}�b���
�9�Aṯ����|�?ݓ+ �ɕ�v���d.RT�QV��&��ɕ�^���'�遵���;���\H�MI�j�Ӵ]	�u�o�{+ �w\0�Ȱ�&�I&�p�$�K�1LLb\�ԞD_��}��RN��]I7�wF��v(q�Hν	�,�=�z���=�����c�X�Ҧ�0�Ȱ�̬�&V�߯��������)��O�L��Vmk��X-t!����z�޻�Enښ
@DPر?��`��cV��m6�@�����wd��6�������l�y`���ȵlT�Qm[��0��ݹ�ٕ��6W�V�uv��5n�	R?v�X�Ixv8`�R����|T��v��c����z��p��JT�� ������ꊶ�	�X�IxvL�ku� �܋ �*�Ԗ�s m��	&���'쏟ڐ(\5�]D��e Xbͥq\J�
�yfK-�ɬ!jY��A�N1r�gYL�HUv���"�Y�rԖ˗I��r,u���v5���;eqL��LvA�H@�S0m@���C!lk�z�<���Z�a�7d
1���=�c�t������]p�m��.��.�HM��j������٨�R�yt�y$��{{섮��G68�����\�ԃ6�c��l�y�܏6g34�&aB˛�A�з.�}���mn�`ۑr����^���kޥ˲��"�R��M���p�;�"�>RK�;�eg�${�~�0Hv:�U�Cl�6_�������Kg���J�<��!��+�WL�i������X��ŀwnE���q��j�*.ݻ�;�e`�r�^�~]z�~X�Ix�u+)Q.���]�whi��c.��[������ ������j����"ۥvՎ��X��ŀwnE�|���wd��%n�/[l)S�L�V�}�w�Y�$��jȎ��	�	 Q���
�S��v��a�n��Ơ{g�����?W9ĉ-W�SE'TU�pN��:��^ݓ+W�.y`/�X��T�]ݰ�EЕ�x��s�W=��k �z��`ۑ`-���ݥeu*˵Jұ7Xkob�;�"�>[%��2��[q�^���c���'���=�%�u��\6{.��m3k� 9 ����N�u�t�T�ZT[k�O_�� �l��wd��;[{�VRt�j�]2���>[%��2���ŀwnE���8�z�J�"հMS�E�n���ԓ��n�66�%Q�!���4
���H�e���&M�0j0&.5�� �E�@�RT�5���0�`��L����\e6�"��m�`�X�`� RCa����L��!n�p��B��������> ɼJ$C)�[E�*XL� �R��I�#�r4�be�L.$"Q��\$2k�)���-5�/Ѓ	� �*�e ��`������0hАI1�02!�t�E�#�����Z� h
'��E��jE:���P�
|��T���w�.����x�퐵m�WmU�@� �m�X�r,��9T�L�z���n�;t�5m`mȰ�8`�p�;[{���p�$/�I۶������we��n.zG����|w�.�����ݷѺέ�QV��;k�o�?������s�ϐv_��	^��{.��v]	�����UT��.y`��,��nҫd�.�+H��`��� �r,?s�Ivy��==�n�2��
�tZUiQm���^��Xg��l�I��� P! H���W0����7ae'Jƭ��.�m���ʪ�\��߻]W�ߖ6�X���m2%vjWf[q*\��B�2��ܤٌ�a��j�-Je.��dm��6�l�Xkob�&܋ �c����q�et�6gRg�O����_����~�u$�g�ԓ��tk�*-��������R��L�V��~��>�ᇫ��R^��V�.y`ک*�g
��	�X�0	�e`��� �r,zJJ�˻�EݗBm� �&V�<;���I��޺�o��f��U(�u	�!Г�^����!�� �*��T<�r�/j���A]�c��4�n�+GZP��p��r�m8��ۍ�x���N8έl��F#`1��\�]�i�
�lG;��˦4b�󦈸�VhpZL�[=���]���Sp5�ɧ��"y����g�luŰ�S�&3���=�6�MR��7:��F��1��rA̮�p�lb��*�^�������L\����@xk�i|!����b`�f����x�9��
V蚞+��FEȂ�\ݕ�t,9��&31u�[�����~�`�ذ�8|�����= {�*M���*-��wob�>��}�e`��� ��):V5n��vӶ��8`l�Xz�ڗ<�O?(�Wj�&�Ң�ف�\�R����j\��&��;�@��իe[�[����`c���l�X�}��By,v̰k����^xQìbv:<�k�;$�ݷU�-�Vy֔����Vʦ��lp�>��M�+���s� 6rP���V�T&���ᨎई7���������|s���&�`m*S.��v]
�f6L�ku���r�����w�~0�&!)������&��(� 1����~����>��M�+ ��X��X�ҡ�`c���l�<�}��x����t�\�jŖ��۲9��2�[����uT���+��d�fSod��U��V5n��v��|g��l�Xku��Ur��O?=JR��Bj�*-��l�Yꪮq"T����� �G�+��~�W.�����M�i[)ݠj�`�y�0	���=\����
�@i!0/ �oz���'��hԒn�wx1]5E]�g�0=U�/Og����M�+ ��p��4�ƸU�U	� �G�+������~0	�� ����)U��k�e$ �Ћ("����W���w��hV0��cu����uۆV�v]��t���+ ��p�&��0��E��jqZ�iX��ku�?s������?{��`���`c�~�s��=�C@�[��V�� ���}#���K���*\��6B*�v+�WL�N�0=�����~�ko���i���Q�*��V�@4i���s]�5��$����Iݴ&�Ң�l�&��r�Ts��=<�`H�|��B��)6�*vn��8�4�ڻ;j��$SS]1������r
j��q�E�H�A�|�����	�� �Glp�&�w��TUۦq�k �0�p�&�ku� �wyj]&5­��M��8`c����U���/ߖ�ߟ� �MTKƮ�uwe�m���nָ`c���qw���^��J��.�+J�l�;��`���߾�t���0	�� �I��n��o�?g+UWc`֩�Eښe,ԚG@a�#�N#�ݶ�s��|��Sr��b	($�Dq[!�rlcV	�j���4�����ӵ��j�z[!��݊KGnu�c �qA<]��Eщ+J�Q��Xaj��dz9/JM����]�SacT\���22�K��F�)���
�B��!Fj��;v.K��ڬ��V{m���Tv�/\�'O9�1�Մ�u���l�v؞�|xő���Og�ۍ�F����(�E� �Tv��U�ڀ}���`H�wc��s���|�as� ��x���cV�鉶��>��=�W*������~���ȰJ[R�v�I�t���`��wKذ�Ȱ�p��l�+t��n�4ـwKذ�p�>���g���E����*��)���;�� �Gv8`��,Vބ���un��L镅�A8XqP/ӿ���=���
*{q�S�&;k��O��Q�U��y��7c��/b��|�}�� �z*�iۢ��m� ݎ+���Vap�Հ}��}#�UUU$jQe%i{�j��b�`U�,�0�\�K���l��v��Q���b�T��X�l�x�;�?v8`z����'�<�(�Sv�鉻l�>�� ��v�b�;�� �W9�]H#�دab��n��g�5�U�{m��v�q���F��c�X<�'�I�h3�jT�%��t	���n��Xv8}_ ���;ݲX��t[)�@�f�W���� �8`�ឮUW=藮�]5E'eYJ��5{޼�0�����TU � )�XZ0,���0�^ŀumm&5E[gJ��>�� ݎ�^Ł���UU~�s�sy�_|um�}��ۭ�˴�]�oV���~�*��<�W���>�� ��%�p�2��L�Y�[jV�[�x�{>��c�^w3���p��V糸��8m�n��XT���p�7d��;5N��B��Rb)շ���7_rs���y��$���ڽ�?s�T�%x���b��t��ݷx}�� ݓ+ ݫذ�%�U�K��n��J�f�U/{�lԓ�1�]I>��q�?"�������}�zjI;��;&1�8�������f��:���}#��&V;q]ҲP���n�T�-4�u�-]��vc�`6�F&]/��Q;��l�t�v錫�`RK�>�� ݓ)� ~Ğ��MI;|x��K��C��B�x�\0�2��0�%��e����.˶�0�2��0�*�T��{׀w�����J�JҜ�Jұ[0�0�%�Mp�7c�٪e��.�ZUj�0�%�Mp�7c���� r�UVU!�~]�!�Wa	D�A>Mܩ�0 ��s���X�k���p�B�� ��H�R��fk)�&�q6a9��j$�M|��(�fŊY"���"=�@� ��&Y��*�h�s�!#� t���o�m�L�.�	<�@�$0&(�"V0�O�kAL��h*Z��U&!�$X��� ��h�lD$HqJ!*R��!�6�3IH+��<��I�qb!8�PÆ	6§����\�\a�C�ab����1������h��!	�bE��� E�0��O�[R��(   �`     �l9 �N�kYS�\���\@rц	�4�x��\p�	1��;Fyݠ;��3Ic��:���I�Q��Vׅ�)b���A��h�,��n�碮��bi4=�0��6���
��J[�@��ie���ZRB �~7�۾�a6kk�
� /B�vxvk�eF��ɇ��;=dۡ�i�B��:j����P�MYm�.�a�z�v�u�d:S�¶7M�|n��a�W��˳\�|Ŷѧ�ٱ���a��.��]�g\�ur7)��&�W+V�uuʓ9=]%k�r�#7m\�c���]�W@�cnv�Rpeׄ�(wm���Jtڠ` ږ��TT���	���x���*���ʇ=�$�4ƍd8�]ړ�u6xz�� ���~o�����&��tG����q���`g�����4��s�;�^7f���ч�F����9Ø�ۍ�P9.6E��������٤�A4�*�-[����ì���4�$Bv�v�.
�h�VuZ�\�<���60��\/W����Gb��]v��]@3Ok9�t<r���4�\����}d&�J�����l�gHT��\�
]��$-�Y�`�����#v[�,fÜ�n�X�6���l�,OP:ﾾ7���K��7O�]��N����Q��m>;X��ۭ�hL]A�>���Ip+��,��-���t�f�(ʆ�
c�6du��*���	��w=+ʭ������6��:�v"u����5 -v�-�E�Eu�l��U�1��6�:�
��C�݆�S�� ��<*�mKəX;Y��K�VGe	���[EP[i�1���'L�n�;Į�93�
]���1à)[���T8}��>~����e�-`�Jղ<5�Je5XW���^V�[�d�#m�N�<�U���ɲ�D��iV�Ce��F�3������	X[��^j뗷]�	�4�yU�b!�z�����C���n���0�m�ߟw�{��{��i�@�
��&��(�G���Qw�b��g|��!'�O��U�UUpG2��d#-��n;9��&s�v���ƒ��JҚ�\<<�sa�p��=���重��C<r����/Hk����r��&��|�q�����[��8aՁ�:jk��FRK�X�3T`D�%����g9u��LJ:��-��ڸ��WV�&���ٻgMtu��q�<&���ԕ��ֱ����������X֋�w����|c��VmkJk͕*��ڸ�j���=n!S=�����[o�{������l�J���w ���0��n��uI/ �f�Wv��CT�Qcl�7c��Z�v\� �G�r�	��^��Wm;�i� ���v\��Us�w�~0	<�`jR��TUۦ2�ـv\� �Gv8`~�R�� �*Q~T���\i+k �k��Og�����r,T�QwJ�<��K�kt1��f�n���>�q�m'y��,Ʒ4��av�.��ceS�>���eȰ��`�ݥe]���b�[�q��'9ɞ�s��*rW9]���L�}�`��v8g�q#}���$��ZUj�0��� �k��0�0ڂ�)]*l�J���w��s������� ��?������I~�߿o ��=��F�XaS�7c�����$����X��L���J.BL�m���\�,�.�l!Í=�V[��>Ø���X�.��g�q,K��{5��Kı9�{��n%�bX�{���~X��1ı=���4��bX�'�޷�1�b��!�g0���f�q,K��=�cI�~D�"b%������Kı=���4��bX�'{ٯM&�~�LD�;�.��̱S�L�;���/!y?}�_^�q,K��}�M&�X�S�@�t8q>���f&�~�ɭ�&�X�%��?~�4��bX�'���M�0v��O:|:S�:Jt��k�I��%�bw����n%�bX�ǽ�i7ı,O��z�7ı,K�Η�1<Yqf-ĸ��n%�bX��f�4��bX��[�߿cI�Kı9���t��bX�'{�zi7ı-��xS���r�ٚ,!���y.;�.z᳑ ��;4 ��`�]|�t1�ZW2�g�.fs4��bX�'=�z�7ı,O��z�7ı,N����n%�bX��f�4��bX�'zz{f0\��d�e��st��bX�'�Ͻt���#���b{ߵ�i7ı,N��_��q,K���]&�X�%�㹝'��E�Y�o�>)ҝ)��y���X�%���k�I��(�%��g޺Mı,K�g޺Mı,K��q?W���T�å:S�:}��^�Mı,K�Ͻt��bX�'�Ͻt��bX��)jA��a�}�}�M&�X�%����c����!�g0���f�q,K���]&�X�%�#�3�]&�X�%���^�Mı,K��צ�q,K��=�10bn�`�	�<#q�+c`��h16�L��(��ʗ\�c��K�2�N d듻�^K������q,K��}�M&�X�%���k�I��%�bs����q,ay����{�{�-��rwy�ı;�k�I�~�"b%��zk��n%�bX���߮�q,K������qD,KĿ�qcŗb�K��&�X�%��{�f�q,K���]&�X�T!��������Kı=���4��bX�'}=�I�Krg�8�i)��Mı,K�Ͻt��bX�'{�z�7ı,N����n%�bX���l�n%�bX���\M��s3q���7��n%�bX��}��KİT�}�M&�X�%��x��&�X�%��g޺Mı,K銜埧� ����sq7\Ɣ*t��u��Wl�`��`�sq���L��d6�9�!�����Ntub!��r�݀N�t∂���d�ۤwn�n�� \�D�C��v�B�)�v6�$��ΨŽ4�5��+�J��ȵ�i:�V��z�>�.�kc�Y��l����f��5I��x�D�E�\��U�av��랶/i�K���Avl�؉�u_�����%��vm
=����0�['F��<�1��#�띟c=�����#T��t��jڑ�ʧ���%�b{����Kı9�٤�Kı9���I��%�bw����s�:S�:_~���������O�X�%��x��&��D�"b%������7ı,O{?�]&�X�%���^�M��	���b~���c���d)�d��i��Mı,K�����n%�bX��}��Kı;�k�I��%�bs�=�I��%�bs:Lz��Hg9�m���n%�bX��}��Kı;�k�I��%�bs�=�I��%��"b'k���Kı?�O�|ڰv��[�O�Jt�Jt���~<Mı,K���Mı,K�ｍ&�X�%��{^�Mı,K�=a=�N��U�S`TT�e�C���;k���9&���s���yz�	�p�I��%�bw����n%�bX��}�i7ı,N����n%�bX���Ο��N����������\��W6i7ı,Nc��4���<'�j%��k^�Mı,K��}t��bX�'}�n�&�X�%�ޞ��ٌ37)�s��8�n%�bX��u��Kı;���I��?��"b'�~��4��bX�'q���i7ı,OϬ��f���&�rwy�Y!y<��ۤ�Kı;�{vi7ı,Nc��4��bX�'}�zi7ı,K�>�~� ݰ�7Ο��N�����]&�X�%���s���i>�bX�'{_��q,K��s�]&�X�0�����˦�v�,�KZ�LM��cd�c��k����]�)7m�d�l·�T��U׎�2ffc��n%�bX�ǽ�i7ı,Ns���n%�bX��}�7ı,Nw��.�q?*b%��~<L~���L�f��4��bX�'{�_��q,K��s�]&�X�%���^��n%�bX�ǽ�i7ı,O�=��`��*y��ҝ)ҝ=����:|8�,K���K���*�'0P�Pd+$Dn5A�X�"�6b&�c�~Ɠq,K������Kı/�;+�1|b\Y�L\fi7İ���Kı9�{��n%�bX����K��3=���4��bX�'�O��!�.L���q���s�]&�X�%��{�Ɠq,K��=�M&�X�%����4��bX�';�{I��%�bs���'�Iq��*ՙ텐��4q��ڝg8ݭCˌ���;�o!�|�y&���Wy��ҜX�'9�zi7ı,N��٤�Kı9��غMı,K����&�Yҝ)����C��E`�K3��å�bX�ｳI�~8���'}�~��n%�bX���߱��Kı9�k�L�t�Jt�K��{���@v�vg�n%�bX��u�]&�X�%��=�cI��)bX����Kı;��g\��B�������ۻ��l�I��%��T b'3���i7ı,N���M&�X�%����4��bX�#  �dI�m���0�P7Ț���I��%�b}�&?S2S9��l�3�&�X�%��{^�Mı,K��i7ı,Nw��.�q,K������Kı?">��?bͶ���B2�sv���t���g������h aղ��V�Mן�4<���66��'"X�%������&�X�%���^��n%�bX�c��4��bX�'9�zi7ı,K���bK����Zc8ɤ�Kı9��غMı,K�{�Ɠq,K��=�M&�X�%����4���1����_�2[�&ns�c81��I��%�bs�~Ɠq,K��=�M&�X�%����4��bX�';�{I��%�b{��Ll����JLۜg9Ɠq,K��=�M&�X�%����4��bX�';�{I��%��	����߱��Kı?Ϭ����̹�
c8�f�q,K��{�Mı,K���Kı>ǽ�i7ı,Ns���n%�bX���$�A�<黺n�Ǿ���UUUv� �ښr0�W\�w0l@)u�ZF�ȡ5!�:�Gg7Y�RN�r�9qn٭�N+�����O��a5�������`mȬ�r�(�֙x��lOb�7�,��۪�yE�r{c�˹����	��s�jq�Ga.h̵�:�����,,LҘ֦3��p�%�N|Fysa�,�Mc�v���X�T4gӜ������[QaLck�;��m�i#R`�tv�35��+5�0�AMAӛV�����M��'א���/'�~��I��%�b}�{zMı,K���4��bX�'{�l�n%�bX���ݷv+���\��B���������?�q,N���M&�X�%��{��&�X�%���^��n%�bY�{<���Fkbl�rwy�^B��=�M&�X�%����4��bX�';�{I��%�b}�{zMı,K����4>L��66ʞt�t�Jt��}�I��%�bs�ױt��bX�'�����K��LD�o��n%�b��<��Jk�i��W3�N�!y�bs�ױt��bX�'�����Kı9���I��%�bs���&�X�%:'����Yw�gnp�UVܾݻ=.�Kɐ�6|��j����q� �-�\�+��W_��N����ߞ��N��޾�D$���5�,K���Kı;�ަ6B��JI1�c:Mı,K���4��0� Ą")� ��� b�A`0@� ��UO�����%���ݚMı,K���Kı>�}�i7�*b%���|_��l��g-듻�^B���}�f�q,K��{�b�7ı,O��{Mı,K���4��bX�%�8y=�bd�qSfu���/!y���5�]&�X�%��=�cI��%�bs�צ�q,K�1���&�X�%���O��جxG<Sgrwy�^B������Kİy�k�I��%�bw���&�X�%���^��n%�bY����I�Y�^2�tLAYI��%X�7F8��<w��[�)F�D��)-WM(�h�-�3f1�m>�bX�'{�_��q,K��{�Mı,K���Kı>ǽ�i7ı,Os��Lf3ff&11�g9�Mı,K��i7ı,Nw��.�q,K������Kı9�k�I��%�b_�vS��3.,Ÿ��f�q,K��{�b�7ı,K�w��n%�}۠$���
;u���	�mS�����<S!�ԟ��Z#�pָ�Ĩ��p��~>H�B@B�%D�x"�S!�81�L�W�jp���G)����P�����s|`hG���2z��u�A\�6)��;����
{�(mza8��I����ζ�Gt�-y݈ �)��4@�A�lE���ĈW�Hv�IzE��	 ��(D��ϭ@��'	�}��T3��`���4
�'����I�*pB:U4P8�kцH��@ۦ}�e_�#���MH�
�$��E�@��($�(�^��]�@M��&t�A�USHPQ��: ��r�0���]x*�D�'u�ri7ı,N����n%�bS����~��T-Ι]|���N���1����n%�bX���~�Mı,K��4��bX�P���{�t��!y�^O|����l�ٌ�+�n%�bX����Kı^����n%�bX��u�]&�X�%�}���å:S�:~��⟶��L�L�����;�����-���.@��#�<�!)��j.���L�\��B������zi7ı,N���.�q,Kľ�}���LD�,N�Ͽ]&�X�0���s�~�bd�qk�����/!xX��u�]&�X�%�}��:Mı,K��}t��bX�'��zi7�LNMy��ޟm�uX��x��:���,K�����n%�bX��{��Kı=���I��%�bw�ױt��N��N����/�2�X�F/�>,K�绯M&�X�%��w^�Mı,K���K��9��@�d �T���\�S��o�{��t��bX�'���Lf2fY�b�9�f�q,K����M&�X�%�=�u�]&�X�%�}��:Mı,K��4��bX�'�;�����������m��힑��7��} �a�s�]�O:Q`�4m�6�����S�O�ı=�k�.�q,Kľ�}�&�X�%��w^��蘉bX��{_����/!y���(-��Ι\i7ı,K�w��n���&"X���~�Mı,K��k��n%�bX��u�]&�~ �LD�=���ve���L�\�ns��7ı,N���M&�X�%��w^�Mı,K���Kı/��gI��%�bx�u�1q�g��2S79��n%�g�X������Kı=�k�.�q,KĽ�}�&�X�bs�צ�q,Kľ��O���7)�O�Jt�Jt��|�����%�b^��Γq,K��=�M&�X�%��w^�Mı,K
��$��%��w���UUU\l�cGGM��l�p%�j�m�p�(��oRx��뎲�eϷn����z�f��ӯ��l���l/k�&�o;:i)p&� m��������,��e���	Y�zz��d�3��f�n>�������.M	e&�E���]x�K�u�u�-�ϊ�ju�I�$���ٽEsX�_���O�&�hg��8m+Wы�S���y9ܓ�����M�B&����-�kÈ��2Ҷ�۳eh�I$��-t]���i�d�e�n1�^��X�%����:Mı,K���4��bX�'}�zi7ı,Nw��.�q,KĿx�/���3��d��s��Kı9�k�I���bX��u��Kı9��غMı,K���t���qS,O��?I�x�əf11�g9�Mı,K߽��I��%�bs�ױt��c��"b%��~Γq,K��k��n%�bX��OZc�m�&-1��i7ı,Nw>�Ɠq,KĽ�}�&�X�%��g޺Mı,@�;���I��%�b{���2PYTS:m�u���/!y�y&�X�%��g޺Mı,K��4��bX�'}�_cI��%�bt�l�O������-�gl�k͕'j��<Y=zԫ��S=��Ѳ۫a�h����8�?x�Kı9���I��%�bw�צ�q,K����i7ı,N���5���/!y����^�K]3f��SI��%�bw�צ�pߺ#� UL�UJ���'�,L�?_���Kı=�w��n%�bX��}뮟��N��}���G�5�nS��Kı;���Mı,K��}�&�X�%��g޺Mı,K��:�����������nu	��(#�&�X�%��{�Ɠq,K���]&�X�%��w^�Mı,K�ϯ���Kı/�:K�g9)L�f��4��bX�'=�z�7ı,��4��bX�'}�_cI��%�bwﱤ�Kı? �������_��vC���vL��|�mpp�>�1ɵ��*�0���4�4f�J8��~t�:S�8�=���4��bX�'}�_cI��%�bwﱤ�Kı9���I��%���=�=	�����2��N�!y
�'}�_cI��%�bwﱤ�Kı9���I��%�bw�צ�q:��^B�~����%�k��l;�N�ı;�w��n%�bX��}��K/�$ 00P��8�h�G��8T((���'�w\�Mı,K�3��Mı,K�_I�y[�D(�듻�^B��=�z�7ı,N����n%�bX��=t��bX�'q��Mı,K9=�����k`�١1�u���/!y��u��Kİ��C�����>�bX�'��߱��Kı9���I�������������2�a(�m�(�6�4L��ԉc&�Qa�ݺ��Z�;+]n��uGj�o\��B����{�G�\�ı,K��}�&�X�%��g޺Mı,K��4��bX�'����7fKLs��\�&�X�%��{�Ɠq,K���]&�X�%��w^�Mı,K�����pı/�:C�+E���;�N�!y�^O޾�i7ı,N����n%�bX���}t��bX�'q��Mı,K��=�wn�a]�2u���/!y��u��n%�bX����]&�X�%��{�Ɠq,K�p��."`�m@V�ECb
��*/�b&1��t��bX�%��Jc�-�	�Lg9�Mı,K������Kİ�Og��cI�Kı9�?�]&�X�%��g��Mı,K�~��N}�>&5`���`m���ml\3
MZ���@�!�K�o[n�	��Ŝ��>�bX�'��߱��Kı>�}��Kı;���A�'�1ı=���b�7ı,O߽��fY���g��s��I��%�b{����q,K���]&�X�%��{^��n%�bX�ǻ�i7����'�����\bZf�0�I�c7I��%�b{���i7ı,O{��.�q,�1�����n%�bX���߮�q,Kľ��OH�\��e�rwy�^B�{�{��n%�bX�ǻ�i7ı,Os>��n%�`~b'�{��q,K������XC<Sgrwy�^B�y��cI��%�b��}��Kı;���I��%�b{�ױt��bX�'��y�{�s��S�w�X�������]���z$T3k��!<z�y�� �N�"��+Ŵ�n�w'��2lqx����m�U��Tq���=g����订v凷
[oE0�3p��';=�\z�+�����ƍ ����	�.��[�9�[��Kp�y8S���n���v9��6���7��F�o2�F`��-��qN�z;X�2qs�9�fY�hbZ4��;KH���r(/PCʧ�@z�_���1���X*1>ys��`a�v�@{v	�������P�e��Y���"��ݝ�'���bX���~�Mı,K��}t��bX�'��{A�B},K����듻�^B��������E�+��'I��%�bw�צ�q,K����b�7ı,N���4��bX�'��z��ݓ����/!���&67���˙��Kı=�kغMı,K��}�&�X������߮�q,K���k��n%�bX��eצqm�2g8�fp\�8�Mı,K��}�&�X�%��g޺Mı,K��4��bX�'��{I��%�b{���̳��%Ͳ�9Ɠq,K��3�]&�X�%���u��Kı=�kغMı,K��}�&�X�%��g�=g&"�
�٭��r��D��W��ð���i�A�݋Z��k�@�m�������u�bX���~�Mı,K������Kı;�w��~�D�K�����t����/!y���|GJ+SmS-듸�%�b{�ױt��> �#��p+��� ���0&X�m	0��w�'��]Ɠq,K������n%�bX��u��Kı>�m��s�ْ�s��gI��%�bwﱤ�Kı=���I��-�bw�צ�q,K����b�7ı,O��ǩ��3��fLc8�n%�bX��}��Kı;���I��%�b{�ױt��bX�'q��Mı,K�v&6K��g���n�q,K�ﻯM&�X�%��{^��n%�bX�ǻ�i7ı,Os>��n%�bX���?YOؘ�ft��6S�w���-vyF ���#Q�[��̵�;]q	�MMs)��&V���y�ı?~��غMı,K��}�&�X�%��g޺Mı,K��4��g!y���)�q�3;7h+��;��%�bwﱤ�Kı=���I��%�bw�צ�q,K�ｯf�7^B���|�'q�-ڈQ]�'w��bX��}��Kı;���I��=0!�*�&p$��������&�X�%��{�Ɠq,K�Og���clÄ́%�'\��B����w^�Mı,K������Kı;�w��n%�`~����߮�q,B����}7�t��6�2޹;���,N���n�q,K��=�cI��%�b{����q,K���]&�X����s��>���ͤZ�$#�2�5n�	�s\β����\��n۪ɹn�l[�(T-cC<k���^B������u�q,K��3�]&�X�%��w^�Mı,K������Kı>ǎ�zGD�-lm��rwy�^B�{���I�~�&"X����4��bX�'�~���&�X�%��{�Ɠq,K���,�]ܢ��q��N�!y�^O=�i7ı,N���n�q,	D�Oc��cI��%�b~�~�Mı,B���i�j{.�&s:�����H ��O~��ٺMı,K�����n%�bX��}��K��hcB���\sP��5����W�)�r�ʛ�BV�N�.��s���Kı;�w��n%�bX�罽&�X�%��w�4��bX�'}�{7I��%�b}�]ZK�bc3)s�(	�ogr�͎��Xz��� ܔyT4SX2�J��x�)�@U�t�t�Jt�O�}��7ı,N��٤�Kı;�kٺ��&"X�'��߱��Kı�O=�>1� �!.�N�!y�^N��٤�Kı;�kٺMı,K��}�&�X�%�����7�*b0���s�+���M��'w����b~��_�t��bX�'q��Mı,K�{��n%�bX��}�I��%�/'�����043ƻ)�'w����1��{��n%�bX�������bX�'��l�n%�`~��������wy�^B�y�Ч��4�Dl�2u�q,K�������bX��~��	 �'�߿c)�$�w��n��I���>� /��P_��(
���PZ����W� �*��@U����PDP Ab�
B T A`	T �E�T �@�E`�P��B0DX���aT �	 DB	T"@	E�@�AP�@AP� cT! T ��DB�b�BE`,BP�E a@� �*��A@U�
��V��*�P_���W���*��U�((
��A@U~A@Uъ
�2��;�tx;^�����y�:�������J�
�         PD*��+  0�{*��[i�MƱ�M3a0��ܭ	��=5#���G� xf\���[��5�޻�lz�4�Oh�[�������͛G� x%���ִR9d�ֵ�:���ͳg��6���I+2o8 <ٗ�ӝ���w4�+ZGM�z�ܺ(��J�mi��u�ٶ֏` �f[ٶ��f�[�l�+X�;b�;��Ǘ]�W�G���[i�  >�d��J�        �ԥSQ��L`�B)��Th�$�� & �L	��ت��=B       SP���bhi�#�$�i�jOO=&������N�w��g���� D��*��@(
�r�'�O��i������X?h`�@�\5 �DL��7��&bv;��>D D�-���U'��'���F{�Nc�͋J������K_	���F@�)���E7���I(���$%�F�A��,ہ�� ��d�A�C�RB�C@7c�j���1f�8�V!s.ar�%�d�1��@�����)�)%�4ƣA_�|4_�l!F�V6B��E���w�(Kୋ���		���h,����L�*�(`�Ĥ�8kl1���)!A�F�)N̄�ѰPP
��$�$��L!���TŹ�2��B+E�I?W����R�mI �ń(��E�h��N����Ѩ�$HS�# ��V�k[��D�d���[8�������Uf!Q���C���XtI!$g��[�h3S)�iа�-��[�,�D�� �vQj!k�)�ƫI���b��g
�n�P	�4R<�pN��uVU��A�h"�(_&*�t,�EB,f:�Ų��-��W�9�#��i��5c
@�PPJ��]�҈��
�� �H�� E�������OILn��,F�B��Q��A�	��XQ(`�	1B����db��-P��R� �D�0ڂ�����>��8\,�0z�Ё����������x                                  	%��  ��;                                                                             �`                                                                            ��                                                                             T;                                                                             `                                  DY�ŬYV����[��݌�E����v� �n�m�u��-�����́!h	 ۻ@� ��D��2������`[n�@nړ-��F��  ���d�[h�I@Hڶ�Ҁ[h -����t�-�����Ԁ IfU�2HId� ��I n�   ��-l�栻ke��[���	�v���U!��cJۓ-a4�)�R�P*��km�i��4��ݪꪩv��m��3! �z� ��f�������-jU�� ��HMUU*�UT�j`�vG��UR� [j]�k$ ��m�ܪ�m �d�&n�6�f̔Hm�m�  -���Ի4=��ݖ�յ�em���z���a���� U-Ԥ�c�vpƦ� �
W���iV���  �@�f&�ƥ` n�n��W��e� !0sv�[Kr"֔�T���@U �7��lO\�)>$N�M۵T�/mP�n&���[�d�@Y�S[��W�+$�E��[V��nȶ��m�:��UJ�m@Ep�-�ګ���5@ �l��.��n��`5�TmW��#l��e2r�V�J��uR��F镚��� ݒ	5����Ɨ����b�P*�.�<���U��ThQ��Ll�<���-�����{ʪ��^�4[�U D�ְ� ������s֗ޑ��t�vP�t. ��6�Pn��b��q�E¯s���0F�l0�t(^��Ў�UCh]r퉮irh�2�d�bS����.��()p` �v��9��+t�CXp��b&�ʮM�<9��0��)�t�~зL�D��Tx�fÂ�4��#�
U��=� $Y'ڸ��juU��m$EQ.���/���     �am               ��              m               ��              m      m����[d��s �::��C�eenm�k�=��6��6mňv4k�LF���p�`t]9q�����Hk��vwa��p�'7m�'�˙��J�QN�g\)gB[�vWF$����uc�-^��E���v�ns�䊗�UKܵ�^������AA�8��������z�������Zְ  [h  [h  [h  [hT�u�Z�q�M�.\�:l9��k��]���z�J����\�`_�7c�P���w�7�f���.}�w��Ӳ�s����QS9���{�'���}��|��  3LK$�f�Y�����_��n����46������̫˵OXJd�m���9\�O~�|   �<}>�^3>(�>n�L�+2�.��Mr�}��������UM�.M���T��$	��3���fu��3�r;  ���]St��7T� ��5�D% �;�
�Za���`��]R�B;��e\��� ������H<�g�J�A�A�)���d@|�z'N��d��"���wX  �n�7l�-�-����R"9H:� �8��kUYQ��F@22��ખs ��󔃨�Y��UZҀ:H��H9� � �t�l�V��9B�1�A��3�}�fu:���@`             �&Fݜ�;t��g��vκ����u�.��K�d�V_ْe^�  ���.����3�w�Ν�n�u�A�<ԩ�r�o�A�) �@1*��;  ���dd�g�:���� �2���K
�� �1���dd� }�{�w` ��J��ief۾u��� �d�̀b�P7T� �����P�� � �t�mk�*�i�r�uy�A֨GS�U�p��n �4#���H<�U�j�<� ��_}:���g^m�  �U�[Jݪ�N����wY �@20A���ZՄr��!���T�����ܖ�U�uq�F"p{��oٿ�a �2����D���  ���dd^������� �SU�d
�-�����Y�"�d#�kv�Dx�F@22��ʍ� �2�d��$ImbU��:� �4����4Aڐy��V�a��N�9�=uH>�3����  Iخ�l�VSt@1c  ���w�:@=̀f2�d ������F@9��b  ���7T��{� �@=̀d`�Mn²��o ���뜝fu��>Ƞ             �f�6�k�m�؜{q�F\�dY��q2�mˋ�λ�:ɬv  ��nCdKRy�g_}:����0�� �@1*��;  ���dd�g�:���� �2���K
�� �1���dds=�:@=̀f2�d ���������,B�%�
�-��g\��3��H:�҈DM�o�u�UkL ��,�)�n �ԃ�Ў�7����:�ՙ��Uͤ����3�T�ʬ��o��  6C4��Kqm�l���ݬ��*��\����	�����d��Q�Qj�	b�$(�C��B%ޯ]K}��4c)����삸H'HC�M~j���ݛ7xH�︪��U�(E]Ay�WZ����y�~  e\۸�-z��*��|R��� �G{�z�jݷU�z�U�(E^r�U�W]���V���Њ����"��B*�x�uV�`E^r�3���޳�����f�'ݹ�<��>   5bf˞����s|���&Kuyv�y��Kv��᬴�O�.�j��'�׾�����              +sfؕq�N�7m睬游n<��|�6�w��b�2�s?���/}� 	�-�!d�ke��w��<�8��L����ׯA�K+߈�N{x#v�ݚ���[��~s�9�}�� l4���>>��PJd�_w���5��w"����k}�i�e��u��r����y�r}-����<�:�ß�� �bm�e�-M�w����<�>���{�~������&m P���/�n�{���s{�3y\�O~�|  ��Б��o�׾���y��9����صL�����߳��Iׯ��5���?f˟}��|���� v��|����}3���̫˵OXJd�m���K���2��e���fq�7U�}�>�              �\��u�K���ϖ�><sѮ�d6��c�i[��+6_.gh�  &�7l�.��[?~~��/o?��d�ns�-��3%��vjwS'��;>����̼���?   U#"]�۰�ə�Y55%��LMIw3�Z�[9�;���}�l���}���x  V�pf��﯏�����~����ڳ��n�I�I6I$}���Q�w߿o|�f�^s����@ �k#��o8s�|�O���s�����fR��n�o��̗S�y�NV�JF�@�����~  6m���Jd�^}}��x�� 7wQ"7��(�6"D7{�Ί7 7�XΚ�L�ݍ��g��d���: G��	$��;Z�,8��A��`� urd�����{�      ]�h                                                         ?�v           .\��r�P"�B� �/R��Q٥ge�'�Ƈ�8�ٵX8��:qQ�^��s�8.�Hq'| �iD��f�;C�X�0�斝ۂ�5����KWgR�E$��m��t��V0�=aIY]�h�Z�p]f̋��λ]!d��2٨�\���﷿���"v��:Uv�ܗݵ�����^���           ����j� ��o�����\W��1νO6m@�����w�` $3b��m�1����)��8��Z��d7v��~�	Hn� vky��M�o������-� )��~�;�  ��lD���^*�My׽��~-��~q�dD|��S)�d�s��̕��~�w>�}�6��{�~��  �	������PJCwN���%2s/*��<�/�`D7U�j��|��es'�]w��  ���--[bZ�=�N�z�Y��wt"}kx��@-Ѩ�W�EU����Q�iC��(W�")�'�S%Gr Db�Fb����ǽ�{� *���O��β��܍�#�w>�����5G���U�>�i ��-������r1R��N�h�-�f���3%P�!�hd	���n�   ?�;         d��7Cv\��5�c�m�Z��U��t�+٫�s��P  ]ٟ	Rez}3�Uz��3EyGk��=���`�fkGPy�@�RfF5��3�}ѻK�3�w3#?,���� �yG�fsz���<  BHjB�ʵw����1�����S�2<Fk舏������q��Fb���̙YJC��;�R(w(�Y����G�  DS,���S�	L��f�f(�=��#CN�(j���-�MQ�l; Y8ek{�����0���Vs�9�T��"����V{��$�>BFw������ �l�,�k6ݝ��sִ@f!Y}�fL�.҆���
w��P�Q��<cW����B�ha�B��H��Ƴ���48�ڋ�>_=�  �П�e�N��"|�u�c�7�Q���ԃ1g�"8,.�}*}�Q�"�Geg�̕C�E���^��R���}�'���>�wwx        �;    �̘����$]�cy7kv�:�7nlWx�ݛ���;��� m�������z��	Hc�e��.�ʖ�*N�P�mF�݅y�,��ܡ�i�G�"�Ch~n�;��ҍ�Q�*�~�:�s�z  i��@��̯J�Fbj1�A����T;�A�����0bf�r�$�3��֕gdU!��P�Q��%"��(�Cu�d{*XJd�m DfL2Q;����  JR2?ffemw����Gr�}�P�k(�Ѥz�f!��A��e�=H�� V�!A1DKniB�!2�*�pB76�H��Mv�Jʅ)�f���vĪ�>j���O��*��#uG9:�<�  7mM��t����2T�"�C���/s�	H���2��Q�M�p%2Tf!v�Ad6�Y�¼���C�� ���P~�6��5v|��2<�'\��>  ��-��mU��w3x�s1S)�:�#��$g��pUI��g�fF.d�����fF$f�{�t0w35��b@*�%����            ��*�T���^���[zW���� �>���s���fu�N� �n�J��7T��cu����_tN���Ρ��1E��(�фz���mF��o�f!#yX���k1	�{��݀ ����j�m�;Ͼ�b���̖Rtb�[��cu���
��dc���m��&5D7Y�Hϼ��v��u�dbMwwwww`*ۖlD���N���u�L��rމ���1��B%s�fF3X�(4*3�g�*��w3�w3#2^m�/\���93��{�  Y�%�
͗;Ͼ�s��}:���y��&dcu����.蝵���C��ՓSWf!x̌i ���-�����}:���/` ����TX�UZt���k1	���Rx;��!�w(m\N߁�*a�T��3{+x%#s3X�f![uuI��f!#<A�o]u�vt             �Rٮ��Y5��bq�����힍k;m�rٲV_s:�v  ]:���U�v��v��=��ά���1�dbF}�z&�w3x�s1��*W�1
�G�n��3%P�QDnιɇ��  .�Y���ޟ2Vz	J38D!��x%"�r��K��c���m��&dcu������/���X>��C��ՓSWf!x���ru}��  ��e7!#�Ui���1��B%s�fF3Y�LP�=d��(�@
�w(�����̕# Eچ�mG���R(n��Cuu��rw�  YZ�v��V�L���1	�]�;ks:�s23�&���B���rމ��~��k��Ada5�T�E�"�a�ڌ��  ���54ZͷgcuE���Чo�̕0��j�Q���mw�)7Te�=����(|�C1C#F��3�2���F��&8!z/5�F���AM3��W9��nu������     lZ                                                                     r�lْL���6�+G���%`���A+�gzn^a�m����� 5q��Jc��	��aB���r�{B�k�j��=q��pk�Q��A�	ю ����N�;4��v2\KmUA�]�z��%�xa5s��K����)p�����}����w>�]y�~뮳�]g]~ϳ���>��              �jYv���h��v�Lu�i���G]t����MP T۴��wZw�N���Qچb��{��=Hn���,�vT�>���	�g�
�<�����̌�v^���s�rg9:�߹�  �g�U�n�w��{��w��{�s���J~�m(��C#1F��1zM�F�ՓSWf!x̌HϹoD��o�\��N  ����%�*�N���f!#>�{��Os�$�Gr����fJ��*��"!^!��n����r1��B���21��Cd���~   %)�����Ρ�̌깩���fF$gܷ�ks7�w3Ԯbj�|@^����x���o|Rx>��C���6�  ݕ�%u�J��n��4^3#3s=��=��c���m��&dcu����.����Ρ�̌����:���93��w�<��@�P             '#�.�	Og���Y���1��X秛g�V��~�}��  "r�b6���>�uxǹ��J�:�21��BG�C�{ઓ�����FF*J	��B�21#73ݒ\�>�u�&}�뛖�m`�!��[��rg�N���N����r)`�h�	�dgVMM]���21#>�X;��c���J�'Ňf��u����  ��+7L�(*��w3�w3#2XUIы�Y���Y �w��C�FZQ  Ȉ���^�&w�n������,����9�3�  Z��f�J�V��1�dbF}�z&�w3x�s1'�EJ�f!V��P�=d��#�b�@�o�dݰ����fF$f߽�  Jn�.�VICs3X�f![uuI��f!#>��Gt�w3�w3#:�jj��/���-�������(  �B "� �      m�     �#.]��4oML�+��e�̃��6j.��nS�  �VKk.�ݷj�ӧg�c5�!#=��T��q�db�K
�:1�dbF}����`�fc��+n�n�3#��$fOo]� �����6V����gP�fFud��ي��fF23�[�5����;��D�bt���k1	���Rx;��u��g�c@̗�wwwww`��l�d�+6ݗ�w;�u�$f�w��;���s1
ۨ�L���z����E��em�niLb�����,ZT��P�H$
�PE*̫�H@�I"F��H�+`�
X�2$Y���P�N�cb.�$H$�� �Wwg��f�OD��u�dgVMM]���21#5�t���� C5���v���>�t�f�#	�QR����Ck�Gu��̕C�Eܣ1eg��*GEچ�Ȉ?ʎ{~��;���s1	e������m]�V~���Inν�g�Hdf(�=�W�����#�Ck�C7�Q����CN����hw(�!��Ad2�ڝ;>���$f�/�>���Z           �*���=�Qƭ�̆�.t�|�lv1n���I�oٟ�y�~  i�ݺ��ts.�*��{���21s%�T��c3�_D���/s�	H���2���DߧS%� ��b�Cj7n�hn��?~�{�˾��  -M��%&g�z0�R�ϠHmG|s�F�r� ?�ƇR�#I��R��U��,��n��3%P�QDn�Ŵ)��3%L2*�f,�'_���  ��	�F�U��`�fk=��+n�n�3#��$g�w��u2A�}��gMM_��(�C�����e�:�Gr�F�  ,JnjF#ml�dc5��H�^{ઓ���!�̌\�aU'F!�̌H���
�x;���s��>A��A�V��>�n���/�� �JIh�D�.m��}�23�&���B���H�w3V�s<�J�'Ňf���{=�U'���C����Hs=.�`           UUUSl��/� ]�>�P�_/S��2Eͣp�t�  	%n�f閝XUI������*���fk��~�	L��]��Y��{�/I��I��1�g�gVMM]���21#3���  �˗WQ��oy�����"W1:vdzAZوHϽ�ઓ���!�̌\�aU'F!�̌I:s�~�l�>�u�&}�����  .A F�VInιɞy:��9���,����ά���1�P ���z��[�5����;��D����93�'\��'_{��  ��'Uf�ëuaU'���C����*cv��Y �w�&eP�Q�� �PȜ����P�j0��"  C�_{��g�w���u���N�ɜ��  -Z�%؉[+f�sq����uq��9�hw(�!��DM;*W��*�23k��̕CuE��@-�N߁�N���fF$e�^ a6PB� �i���[
Xv
�.�l,"$,�Ռ"I��a@��5�s:I����y�s�}��}�      -i@                                                                    ���-P�L��V9�ib�t�4����ڝ�#uw�^i�[��u�Ƨ������W(s;;&� ̛d�tU� ]-'F��:�V�8�4�6suI�*��<�Lg���7%��h�kl��)��6&��H�vm��: *���c����6�?v�������            UI�k#�
�b�tr�mq^ vZ��F�[�����  ��A.�P����hn�!��a)���.�a�����&�r�#�Fb�5�Q���Q#3�[�5����;��=R������E�ʃ��o}}��{�t����
�<��$�%�C���T�aU'F!x̌H���
�x=��c�����w}�-�׾����79��9��� Kh���~�������~�:�s�����o
>�2=J3�_A��e��>�A�K���\����O1��!��{�����*��~~3�w3#{Q�ڭUUS��\�o���|�_;.dU(o�$6����L�ˠ�!���A�Д�P�j�;�1zM�u�,~�3k}Wg�^3#N����  �ѹ��6�hn��!��@24�^�ЫQ�f&F��2U�Gr��=��d��"�Fb��{�L��2��Q�|NS��             ,�J[�͌�ֱp��ƶ��]��%�*;<Y$��-  �m�2�S����Rg�cu����_p��`�gP�Q���e�}��=H|[A���
4;�z��C��4�^�ЫQ�f(� w���  �jXͲ0Zʹ��(�������� l""D��Q���:�
d��Q��ܡ�2����ϼ��1	�������1��׾̻�  � ٬WJ��Wf!x̌H�|��ks7�w3�\��ّ��	�Q	��r�Os8�s21w����3���t�  3D��`ڵ���}��c���m��&dz�������פ��Qdw(�Qf��>���V��=�L��z&�w3x�s1V�]]��� �����#ml��93�'\�A,{��o|���������̖Rtb��Č��p������w3����vu�L���79����|�             d�:�'�1��ݶ5�zB-�V�L3Yc%���vw�  U,�#"]��|Ϲ:�Gs�y���5v|��21#=�މ��=K�ܡ���zB�F��]>6��>�u���N���9� $���˫N�ՅT��c21#73�*���+��V E��s�9�3zuf���RfF7Y�HϢ��,����ϛ�<٧\�w:�&s��}�  
H��0Xlo��������������ӳ#��$g��r�Os8��Yq#�lj	r�1�=�hq�P�ҁ���7��c�o�/�f�N���fF$f�w
�x;���s1
�p   �%�
�-&dcu����.����Ρ�̌�ɩ���fF$gܷ�k��Q�c
^B%�S�gc��$g�{�wv $3d:�6�m�;Ͼ�v�s21s%�T��u�y�y�A%��ª��fk|�B���21��BF}p��`�gP�fF,��U���ݴP           UUU8靥%XU6oi\�qs<F�͞�����6`  ʻ�DJ�V��1�dbF}�z&�w3x�s1��N���f!#>�{�Rx;��;��Ls�3m�z��}μ��rt}�����`K����}��L���7+n�n�3#�	��f!#>��Gt�w3��_|ϼ�Y�M]�!x̌H�|����>�t�g�N��9��  ��Ui���UZt���k3�Ǽ�v�ʨ�˄@"��Pڸ�i��3%L2*������3*��釈w(dM�2Kvu�L���79��9��� ��]�J�Z�iзt�w3�w3#:�,��F�V��X �s�F�r��>���J�'Ňf���%J>���ݝ��N�����90��  WWIURaU��XUIшf3#3s=��,��c;���P7T����>�Cj5���hw(�7P��m�Gއ��u�L�'O�y�             vd�ݺ4���r�Ge��������5�V�$��-  MիWv���n�P��w3x�s��J�M;*W���x��ڍ��3%P�g�fF.d�����fF$f�{�����\�g�N���N�  ��T�R��WUa��̌n���E�#�X;��5�r?� ��&�ϐ�g�bb���P�Q�Cu�ɧeJ�6�Z뛜��ϻ��  b�WY�c.��Rx;��;�B!s%�T��c21#73������@��!R�����.�a���]��4;�a�3��`  �l1%ŗmlӨ��21#>�#x;��c���!y,��+��j�5�\�U�F�"�~��Rt|�c21#?{�.������Y-[0�V�K���N��Ͼf![uuI��f!#>�����w3�fFud��1�dbF}�xF�w3x�s1	K��RZP6G;�)�`�I$1Ɉ����b�1�ff\�u�Y���?~      �]�                                   �`                                7
ݳ�Z�@���e��+	"i2KI]u�N� ꝗj�j��"���iWFv������ev�k�{S��=�FfoQ1؞ :ѱ�ҭ�h�	h�uW�L�5˛F:M�@Bٳo�(�~]/=v�a��-O]V����JZ��^���~.�4,�4h�aQ�Sz���+���            
����5[uѻ�]�݂wTnyqr��Z���V۴�( i����[+���g�$g�g�Ω��g�fF.d�fJ��*��@-�ڏ:�	H�ܣ-��7/�̒ݝs�<�u��ru}�߀ �MFD%fٽ��N���ӮFud��1V�f�Y�����O����(�!ܣ�}�T���/2,nc��~������{�}:�'\�  i݅WVj�:�VRtb���T=�sۼ�C�}C�;�2'=,%?yL6�c�~BF~�?�M`�f!�̌�ɩ��\�w:�&s��}�y�  ,СIݧiզ�w3x�s1��N����ϐ����:����C����ªN�C1�����	�����;��Us� �m%�]@��ң1
�Fb��[��47W�P�;+�z0�R��j7��hw(�!��B%S�fF7Y�H͂=ޝwwwb�            *�����^���m����+�J۫�1tu�N��]w��k�` ���V��e���q�db�%�T����}�Y �w�
�C�FR�0�~�	L��f���\}�SX;��w3#7R��  YWv�l�����x̌HϹoD����+��D�bt��]���Q�Z�L��(���z��6�/\���u�yz�ٞ�:?}�  V�Ո�.w�}:�s>�u�n�n�3#��$g�pT��b��U���,���f!x̌HϹoD�y�ӧs>�u���^� �ںV��UV�;21��BF}���T�w3�w3#�,*���3����ખ�$��k|ő�	�)�{uuI�93�'\��'^�׾���  �0���իn�*kG�3��df,���q�z�f!���9̣C�G��F9�ӳ#��$g��>uOs8�s21���}߀              l��6Ė]�k��˺���bg@ݍVXԓ%nϳ3o}�  5b�:�����*�����1#73�T�w31��bn�uI��f!#>��A�hn��7P�j��x/C#ԣ1g9:����   ��Ij��Z9�;��9*��;2?Q ���g�{��g�:����C����aU7F!�̌H���T�w31��b��  m��V�.լ��3#��$g�pT��b���Xњ�k���M)�8GU��4���`2n�Hd�$��Cx�@�G0�w��I�m,�@�EࡓL��`<Q:g,A��j;��hw(�!���"!��eJu�<�u��ru����  1[�,*N��U;uOs8�s21{�ªn�C1�����
�`�fc���@�RfF3Y�x�'��}�SX=��>�u�L��<  ��nO)*G���0�R��Q�s�F�r�R��"U1:vdcu�����>uO���oo>ͶNv�<�s'���             ,ݒR�n�;n��Nv�Ą�I/Gk����{��*� 7md���E��n��{f�p%2s*��ͭ`�-�w{��Z�9����������;��  M]]+ñn�U�NLɻ�q�~�À�����Y^̻���fKw�����O9ߜ���gW�}�  *h�Xwwua��ݽۿE�k�R�M�r�jkޫ$'Ă`�_��^���ٓw�����}�ϼ�  �f�uV[�
���&�m���^�߽�+�n�Mc:�k�ʫZoy��1p"�Ep����{�v��w߾�gY�>�<�  �f�66V��������͖{�}�ޗΩ���$wI[sછ�\����n��}��3//`4P             �&Xm���X��N;m��&���)�;bՇtݤ-�C|	� �7�  �D�K��[�*�ڧ�%2[���e��}�v�ӳ7�k�|���e��}��>�>�  $�lWV���-����<���6�9�
 ��H�7�r��
�{�~�������;�y;��rKw�|��<���  YWv�Ս�����y�o~��}����9EJ̪��#3_�Z�M����y�m�s�9矏��  �[V��������v�v���n�I�7^{��-�w{��Z���G hfM?6o�׾�<��` %��=�%&g�J̪˷�Ūe7���=u��N���߷��-ߛ�S��9�x�?h�_�$$����$ D����C���i @R��+'jԟJ�,� ""�QPI�J%~��nH"�(��ȥD *
����Q�P������j�� >0/����~=�����R�׹R����_<.@�Y*�|d�W�� D�A�[��j�
{A ?B D�����)�����������9�!�� 4~��C������<����x�	з�[���Ϭ�|~��f����O�70  
�Q8����DKDP��@BXC>��d*:�n�c�w��eO��D D��RB�n��}�a�~ ����<��������q�������P���\>c����<��r-��-���������������=���� :`{+��>!	��#�Z������ �"y�@O�x~ ��`��zUP�Q����Fȡ�,��;��;�M�){ϙ�Ȣ%!g$F��C�n�d�>!
R�% D���a���>�R +�A�:1�`>b 4�09d��sj������J D��T>?x�A ;������P��p�ϸ�w�Ñ�xXg�(� T�y>�y��lǠ�&��ϰ� ���ިk�wwJ=�=�����l��=E� }���� ?�����,w��w�`���ɹE�?:_s4�����!�@��Dw�3���H�
�Y��