BZh91AY&SY�L3�� _�pp��b� ����a` �P        @  �        9  �  D�IR�P PH � ��
�)"�)B�(

%T   E   "��  @�@���� � {�ZUf��k�+�ť;� (w�ť��뗓O[�n���)@���\ZR��  9���y�
���;�=P�0u��@������*�#{�4 b;��  P *�
HU(ZaT={{�}�|]�S�R�iW�� W|�W����mm����MK� �S'������nT�eO>� �+6�j���/��JŔ�� ������ri�˕zr�m�� ��*�� �H���
y����st�\��������P=�X�����i��L�uo�� ��N]��O�ϯ�o�x�W��yһ��ziɪVN�n,�[�ޯe� �{�t��j����wԫ����AD�(U �,X ��3���w���[�+�u+�@��_nL�NN��<��{o0��}� ��J�|s=�:�/]�Ӷ�}����J}*ͼ��^;���μ�y֟x��=����\�}k�-=��7J���P��@ ��*�̀ �}T�ۆnL�z�.Ӿ�T�xU��|���Ů�9���}�O����_-s���ם��  n�ɥ_s��ڼ� w����֥ɯmw��}}��v���(��e˾���/{�����w]��     P���e6ҩJ��S	��ѣ# F�24"���T�P �#  '�UJ��M@ h    "{JQ?T�@4� Ɉ�d ��S�UJUC i�  )	3U%LЃM=�h=M3S�����W�z�o�������u��k��AUá���
���TUT�¢���������AUo�`�����r��
����t*���������I�YG�5���9�[��|�	NLY	F�)�l�7����.byN~!(<r�r��s_�=
/�4o/���%&%�7k� �����ǱN	Ic�,p�<�h0��j͘�t���7��g#��i�Qfb~4ţs�0O����G\Y�I^������#��Q�?����|r<�7xp��x?�Uyf�_z36>߲��L�|�it�i���MI�d���N��,wύV��iލV�F����ȃ4���o^����[���y��py�ằ���NӖ���>S�����l�����X4�����:9����f�g<7���3�W�;{�"J��^LED\Q�ܵ>�ۓ�j�>�^p���$$���8}��6T�	By`&�pٮf�#z����,��;�h�R!(�l�%���X��/5̝f0�K4n���S��p܆R��X:��c��� ����FXbE�����7��>k=C1������7hoMh?Vp̃[�5�k3E��k4c�̸K\�Q�NG���O��t~�m7�h����k3�Y�a�+���u���f����NRjl�G'5��q�'��q}����5�&�p�J0��K�k5����|���y�Y�y����k�`?/��	@~2B2�͜��尝f�8c�F���p�F��~۷���'���h��(�#�q���(J����.BP��c�?n���<ggN�ѷ����Cp��泈V�Թ	���%8�����Q��%����Fd�Ѽ�x�	F�q&��9��9K��#�Ƶ&o���E�Ra>kD�Q�<��̖Ȩ��ћ8�X�D��fÛ���tn�5	O�BP�&�|*C�b�7�f���o\#t%/!���zƍV��퇅^��<�e��I�`���P�d'��eS���,�m���	_��5x�F��	�bi7q��%���}�s������6Ѱ�<�1ѩĊ���D8TJ	�	�t�dG�`�d%	By	��%	BR��2!2�&Bd&�)y���|ϯ��O�����������X�`�Z�?X^�{����ub�a͉BP�	T	�)��nBP���%	��$�(MBP�����/�i�o4�RPy.QTN�� �a�𩭚)9&&�/$0�
��6H����pʚ5��ߢϵ�������Fy�NK#�	�x�P�`�~3�����ЙhjR�qͿ.I�oX�}~wY�<��� ��`�J����F��޲)��]BP�bE��Dd�&���<y����ddm#Y~#�j\����yA�㪃$�dՖ&�_sF�L�Σ2�#��gTS�����r��f�$� ¦8y��a�C��?�dC�ꊲ�l�>iʎ���r��0�p�}�`�\q��4d��kn��F�֟jq�<�Q~=��,�h�����-��4`9^��rU��Px��2O��6aE���l��l�I��&;5	A�~�8	��K�MM	Pp,��AY8�&De�S�:7�y壛ɏ��oD!� �$�>ާӨN@h�x&�<��F2�>�C�dZ�K�`G�`�%	K�'��� ƌ��?��*����5�^��$}^�98q<�\�f���e���y�mߙa��9g�w`[5���&Z��8ލ.�I��D��z_5o4��}uI���y	BPe��#/�~�
��I�d%���}��2N'��(tm8��ZM�m�m�璮U��L"T$�>��Y��w*~�q������p�א�O0O$�d��A�_�a��<�y�q�9��q9�4٭\��9��O��B�X�:�C-7��&g�dE�<H
��7s�����3ۚ�"4~m[v��f���o<���۹��.;u�~�m���8�F�P�l�翼�g���K��~5��#!+`Y8Ay�	Bn|$�L�%	@a�!����6�RI�4Bn��9j]:�\�� 7	�L��(J���e�9T�21��M�P�&�(J��(NBR��d�faj��\���Q��;5�ky$�L�4��M>p´�r㖒4}���A��<Ǒ�Ց�ӫZF�Q%�%5���"�,�Z��6n��<���kXBP����d%	BV����Ǒ���a!yi��z[��π5P�	�A&��'!�Zw�a��F���^؄�&X��4��\ѥ7fs,�������&�:�̍1�����zI�G�x%��kr1���h��(�1呭�� 绀�!5:\�q?&���5�I�a�V��OJl5�\0�F����W^��{�Cu����;�]����s|9�9h�s��Q���!��>�,�$��y�3[��M�33Z Յ�5ZY1�Z
%�����J��(J��J�7syfk�k�����o�̼&�+�d%	q|r\k��NF�!�������{�5�����$	/��hr��y�Q�g# �m�gp���O3#��r��(O!(K�+���;��j�2�m4j�{d����Y�����aʢ�����V�v|{��,��16��&�2�OX�A��JG��(J��A���(|י�����Y����~K��F�_kD}�����Й8�	X�BP�Ƃmǅ�Z8���*kQ�$�jM9I�Y� ��,�̃vE�<�n��Ya�I��l�����!ɦ
���#3����ƣ%�rv@D55k2��9	BP�P�kI�j<Z���Y�n��2�,��V�e\$˕%�h��$y�����ѩ�4��\(+#+,��4n��x���(NA��0&�1��JK!<��,�M����d%	BRp-�s0J��(J��(K�k0J��d�>~�Ô����k�y�}��F��g�}�P���.99I�A�J��`�%	BQ�2��)12Y�P�������Y	��3�LhJX�BR�bd'���!��A�;�ᓇ��~a�i����T�?�M�#�f'�e��5��
P�c����:<�Q���%u���492%���Z�G���2����K�����~����a��%	BP5	�M�MƬ��J]98u8m5	@}�B;�FF}�V�##Z5hp9�2L�$3 6f��լ����_����S�������e��P~�m�����5���Y��ÄQ�rrrؔ���J��"م&����eh(���fJB$�k'd����kN;<�`F�[-fa�؆F����7�0/5�|'<���P�����s���Q���vk'�����DOύ`j�!�2p�x�
��&Z��"�3\�a�5�e������3 �P����%D�	BP��FN�_w������kXa&���Pa����B^>>���0nՒNG�_�5�nL��čjݣ��#�A�dh��x{�n+��P��5q�xo�{�l�G��(�u���5��c�9$kg�x�}>��>_<�g6�����f~���3��MɾNox���;��>�y������0?&���e��Ԇe��c��A�py�&���!�\�c-�U�@f���s���x��F�<��f'ɑ�dd��P�����M;���(J��H{��%��~N�=2 �K�3�#~�n�4��{璥�����FT��A<"y��%�Ͻw9�J*y�W�R�TA�r�SW?w��B�3��xil�w�Ʉ�9�6���4a��{�o�~	�c��~��v�f�Y��Nj�$�3čBS�9b�޳���|N:mO�w�7��4����Fo��x�ݭ����a�?o���eZ6��g�sN�Zیfi�Aj54r�*k�=��F��MZ���lLa�՚p�%	BR�%	BP�%	BP�%)BP�%	BP�%	BR�%	BP�%	BP�%�J��(J!(J��(J��(JC܄�)�u�>�BP�%	BP�%?.C��`�%	BP��>��J0��!�%��,�u��Y�dQ���f�6l�[����9��	Y��`l�Z-s{���sZ0("3�6oͅ��?kZ�a���)�2�W��+�2p��%I�r��(�WP�%	C��~���w���w����}�o~��ߜ �   �           
P     ��   m��J-�Ͷ           ���  |����HH      �      
P                   ��  �            �P           @        �R�  ZÜ�[V��m��&�6B�6�q�  �� N!�	�9%P�^��kmV��jZ�`6�N�tݬ���$�� m�      }W��U@R�i	���U���IN�S%PSm��`  ����� m � 6�h����M�Z���� 	2�����  ���a�yk��]4#N� ���  	 p   �  3���Vmy�.�M����yk �"O�}%�]�����@UU�.��@Krcm��k�m���I�mH	nm�m���-��m   �@U[T�Z��U<�,�F����������=i�c���D�$�k;P ~��  jMA�UTv;J��Ð���p��m;���oM����`6UU�`ؗe���Z�	e`� -�V� m�mR��S�q/0R�UP6� p	ۭg�i@m�� ���-p��-j�21d��P��C�A� ඖ�Uٹeu����, �dh� v�-hZl6�`$�Km��  -�$��].��6�U\   p  �6�徧[BG:�m ��l H	�`�n͵�$U�   8u��6�@�8 �-�H �[A�6�8Wl$m�Cn�׮�l  �J��m  m�ݲKooH[�  � ��kn����P�Ku
���	�$     N���gm�  h����,�����Z�$kX ��@�`M� 	N�$����[@6�bC��Z��jX��v����*��Y�f���vs�.������&�� ��m��K@ [�m�89l�k�Y@����� �lݱz�x$ 8۷aą���  5�m�Ѵ��MWJ��	-�ն�� B@ J � �M�l  V��h [q$�v ls�m��  @+h�
��)kj��]�Zl�  �am�m�kn�p۶� m�p 6Ͱm -��� �v֭i6m�}��&�.� ��Y@-�i0 p$8-�om���im	 ��n� ����  ְi2��Ԁ   �   ��B�i�0�   �����(�6ض��i6�    p���m�       @�6͙{[�%V�2d�)^���r�m�+�PlkX I�Ԇ� ��l+��m�j��(�� H�m�®�T�x�^P �Ul���I���@	'�[���t�� -�?@� 6�� [Ԑ[f�  ��     ���Y.�v�mmL��` ְv��m� �@m����U��v����V50T��Hh6�|/[�     H     9�k�e�     � ll8  ��@-�l6݀D���]�]��l [@��[A�I�l� .�Bi%�� �       $    H-��z� ImN�Ch�)�N}l��Ի-�Mk �n m��6�m �l�,0� �� 9U@T�٧j�.H*SXh �
q5U\�-T�U�R���nx@�X@pU�-���v���'H�` nNɦ�am�ll�����hZ�m��j��V����W[mJK*�c� �u�h�#UR�-W@����ďAq� U-��
��B���],�mm�l��ݹU���`*��
V�!�U�7J�6��M�hj��� hkR0pm�UUU[J:U�Tj-��mf[u:�v�[M�l  m���/T���M(��R��[J�
�R�V�V�T��� B���G�}� [�+m�d�kh���p  n�ۀݴ�m����m���*
@�d���L��"�/�}�� ��mH�ں¬��eU�%��Sj�m�ժ6�8  I�� 8 $m��         ��v�Cqi�ye��L�KKN�v�����9�����hq����Ij�cIKu�Ȼ�M��m��8�I�d.Qz�K5ض��ٶ l m&���C���n� t��.�Kchm�=!�M��ҕp[E(��3%I$ -�۶�X��um!�S��&��ě[)�����l [oZo[�I�@ s�� � ��I�  ��4IO$I m�lpʻ���{M�[@ Yc��5�f�M�p���
�T �khW���>�} ݳ����[t�V���U���}��+(p�UU�m���5�    �JP IH�e����RK�� �k5��ٛa 
R�5����aV^��R����m [@��$a"魸-��0ăF� j��U��MRV〓�m��ͺM��f�u(	�N��mnl    �            �M��� �ڶ	�$��HI�$8�	2��-W���V�v�tٶ�	    ��pڥ\Xpf��ammn����Y��l �p�A��m[:mpp�i��/�e_����VI�TIz�    �-�Em� 6�%�1Ĝ]e�e՛   mY�g+b.�\-��uu@P
D�W([*Ԫm�`6<��JlU�t����DI���"�u@=��%s��TdX6��H��# -�5��  �� Z ���B;`��\[Mk[[l-�   :���3�I� l   9���-�e��[��v�mSf�Z��[I ^��H ��Y�m���O������t�*T&UX�i�e�mTڽ�H	 oY-��۶�J����b��*U�h   8$�ڧfۤ��Cm����ְH7'[�b�[9!�� JIp�h[#msm��z��n�w��3k��bB�m��'�}���Z�    �` 8 ΀�]�i,6�SF��kX^��l��H6C���M��n��     $��F�m�չ��=��gm��зt�ע��liH�N]�m�  -�۲(:M��Y�6ݍ�d -��X��       �j۶m��@�v 4R�%�v�p�:�ȶX�m����d $  �{XknYC� i�q��$�m� �m��� �Ę�d� $�6��p���ll�m pm� I  A�/E�  IŴ��   p   8     )�6�M�$�*ڪ^%��A��
��V�[V�Y�I��$� [@   �Ͷ-�m��mݻc�	  m�$8���n[m���ԫ*� RE+UU) 3���H�r)]�]nċnٶ��M�`   ��  	m��Ӈ�   jջ�V��4��VU�h	vP�V�S�� X`��%6��ؐ6��[B�;K�` 6��H$   l    6�    �>        � 6�9��-��W��wH��$umuP6��(K� �   m �K-�B՗�8�0�f�UP-��ﱶ>��W 6��Ժ -��� ��m5Wm[l ��8�ie 5�4۳fȶݰ p    $H �   R�2��� �  �M�p  �$� m��n�T�l   	-�m�KmhHm�� �۴�]6��Im��   $�z�@l  䍚m' hm��j� ��K�l H   m @ 	  �]6		   ڵ�(H  dM(rmpo���<-�$ �p u�P�`�8	@I%��hl�`[@:�I]��:��pX�@��
kp  ����k��ַm� o5�� �.����c{cn����i�On�l�Finz�۪����ڀ��ʩ-A�jP3��h���tm� �h�]&�c"�Tx�S*Аm��$�[E� 6Z�$R4�g-�[cj� *@6�6��`Nn�$m�G�{��UW���*
����K��������������M���
��8��e� ���n���L ?�B! 
�h��)�`!�C�Q����.��PT	#� N!�O�M���~S��6꞊�� VD��)�UN!�_��b2L@��	� qC` lS� }�OA<���"IJSB��B�	��$B�3L��P�	M!RԤ�
D�,��B
�+T2B��(| ���B�PP�߄|�"B1�8��A���P�A<@E�&�-�?��O�*�A�p|T?&i"���^���l@P�*����F�	���!GB ��V����O��>�SQҮ�^ ��t*B�<@x��~P��L�z ~�M��� UW���������?�p��$�!Adh� ��ĦQ���ww{����_m���i�  m�( �ǀ      �     � 2��lM�ۍ�GM��Y�M��l �͜Y�9`�%�)��k�An��km�լr.�6�b쁘x�j!�5��h�]9�,��t�v�L�6j�R�\�g�vc���[�N:�p�;k�+T����⍗/S[AvOJ��w	���-`){Yv��ϳ-V3�l L"��۠�$���F۲Gk�����G�
ꒀ�v�\��hH�%�.��Z�MB�e�-�!Y�S;�Rl6إs�:��lIzՆ vU^�N�Q�K�/ ��(�YR��9n7!�&m�����q'3U�ju�LK�I�mUe۠j��L��VgF�����	��ŖF��ݧ��A�,.v�7-��,!m�n������qˬ	�;jnNq7S����۞���d5�1ٔ		� ��t��3�o �&*��JNc<�>6��� �X*���%ƃ� qq'2�d��D�tC�d9���m�9�rW!n�6�VF�mZ���i[��<U��N�-.�ã\]�Y�Ĭ�1����|�ݳ�s[*�vQ�yp�n��3m� ��^xP��U(�%�͹�hc�� પ�كZ�U���ѭ��WFX�e�gpL���cTp�;+*��&�#%)�M'b�L�h��Y��#b��9�Z�]�v]cNŁĒ�Uڴ� �j���*@�ت�C��r&9�eiX%L�뙤�Ki\�C�UR�U�癳��ޮ�܋]S�T��s�܇KԱ5*�\QUK;�������k�-�@m���m�d,�t�ԩ����Ɩ
�Ld�������si���S�Lu*�$$s��lq4�#�Ͱ%X +�P�b�Y�
�u,<�tE++�U�;A;��Q��eX�7k�V�*��)�@ݔ���������ʴ �DO���PЪ� ;@C�|��f��zެ�Uk{��*�T���]����x]���p��c�\��6JSΆv�9Յe�v�s�1��T�T�Eۅ��)Pv3`
��db�q���.��ΎL�������vM���rB�z:��q�u�1݆��cj�Ӵpr7貸�y܂�\]�&��w�]��c�k�ld���^t�	�n�l:�m�##u��3v�v�\�����{��ݩ�9s۶��G����wv�a��+�	�v�g��$!�$�4�H�������ޙ`w���9r��7�"�Q3wuT�RO;���Z�D$��!D���P��8�ݜ���i=��3��M���� ��# %x\�0��ytMX�\�5V`	r���^ �,��ﾁr�`�@�"誋.�������^ �,�rY\�0?���e����Ŭx�����뭜X��9�Z.��=-����en{5�Ն�b�j� ��# \�.Y �+�=���A�LkM���s����6�菢,�ő�\� �%��
�(�IpT�Q4v`\�0rW�w��g �lӀ{����ǒB|6nL��^�K# \��,�}!��A0NN�n�8�}�o�� �r���^��UaW��\�Uݳ�a;\�a����4�ql�+��2h7JN�S���6���n9�'��3�o�i�=ܲ0rW�o%��t��]�M�U?MU���F .J�Id`���}�f�=�5��#�P��� �o��^}��9h�$"��"�B c
�@����(`���}�I]� ��d`�J˪.�j������RY�h�;�d`\� ��cl6}�Lo���7}4���# �x��0�J:QUD�D�M���6T�O$���ƻ���b6����<j�^zvY=���d��k"8vk~l$�F %��Id`	u� H���(Lk7&pw�8ww��7}4�����;�2kƤPCF��jK# K�D}�w,� K���4���6�x�s8列���9U����V���uS�D��w~� ���18E�n���8 �+�5%��%֌��G�0�Q.�lyn ���g^53c8Sk���g�c�p���m/���;󻻮���r���n�w�ӼRY]hqD}�	'����;�X�����8ww��7}4�;�d`\� �WU��.��*������F��# �x��0t^X��blpX��3�}�g���p.W�jK# K�F �%U�VMܑrPQUw\�0��ƀ�yw�p�]�����K0�#X��?!4�v��@
ڵ�4Eb,��Pן/[f�KPt�^烵"���k���6�dۗd��XL;\mu��vrAk]S�'���6#Mm���8�[(=�3u]��<0��M]�qp�	��įPw=d�Yr�����b���s6{rV��b5��R����=l7h�"��vg���b�M�@�tF���"tg@=�����<��j�MD�km���o6�᭸�'�J�B�e���TYN����k���8ɻ;5;_�d`	r��r��� K�F��#X�M�ci'�ng ���8�����d`�d`��iE�w ]E�M]� ��F �,�y,�.YG|t\**�˫&l��� K�F ��F �,��ܲ0ˠ�w7TE�VASUq�/%��%�# ]�# K�F�#�v�C�9�w�9���ӛ�����#��cKt7I���8�덜9����.��/=UD�Uq�6�F�֌.Y��8�~A����C�������ӏ::"�V�# �K# K�F �%U�e�ܐTPQUV`	r��5%��%�#�{ޚp��L�ؤL���I�RY\�0�`	r��=<�(���_IPMD�U� �,����h���jK# ��	Q5�ˋ�.��=0vn���DN���a��c�#ö۪[Z��̑�L<��8�� ���8�Y\�?���(_).QeՓ6A����J�(�Jd~n� �:T{�Ӏ��fȣq4��b���n�8W�{�H"��)�>A��[�� ���8��x�}��oM���d`�d`	r��5%��
H(�E�ԕd��U\`�h�呀jK��7}�� g�%����j"5 0P��%�[��qsH,��n�Gk�V蜧0b����R	��1�p���g ���8﷙�=��\���&�jEL0`�RY\�0��8 �+�2r�I��	�M����py�W 7}��wwy�����$bp<��U�
s;�h�}�/3)PuD,"3���b^�� �ߵ5��#�P�K� K���d`	r��W)�=��e��n�֮]<[�����'6�pP�V8�n7V��;M �M�/0n�+j�c�M]]� ��F �,�ur� K����M���#Ǒ1$�����r�}�F�9�Ӽy,� _�QH���*Ɋ��� ]\� �x�Y^�g ���$$S �4���`���呀wW)�7�"-TT�͑4PU�����呀wW)�/����~Y�>w�w[���kY�  �Β�����_�������m��^n;k�+��ݻa��8���d����A���a��!2�g'd4Dfh�Ƶ޽�3�D�L�g�;"�uj$�E��b�M��2Yi�����l@:.	�K��^3H�\h"u�=j���z�t��'���!%�\��v���OD�v�I6Zfz�3�>�魢7�q�^z�\���N1w{�+m�� KwZ��pT`�Y�qa�nI�N�sù��6[u=�1Cn@�q84�Ong�?���3�{��p�d`�d`��QwDՄPY7w��8\�0�0�dpg��&k�G���p�o3�oٔ�؈IB�o*�1� }�B��{U7EM�sUq�/%��%�# ]\��n�y��ىc[>dx�&$���5r��}�5i΀�y�Y��۾��r�&�3S�٥���[:3�:����g��Q�{]{;W�y`��q�.�S�%�# ^K# K�F�7_"�ML�Lkqp�o3��y�}�]���`ܲ0��p���wudM�wq�/%��%�# ]\� ���8�=�[��kx6�p�,�ur�.Y�Y���QwD��5d��B�r�}}���<��L��Z��(�H��1@�%�՚̭ٹc�E��M����1n�Gk�v�g�-��� ���Ӹ���B\�!w�g�]*����
�nj�!j吗+�]�Y	v��~�Ğ��Ѝ�LI79��ٙ����'��?��$�U~�hO?b8$`A�������)�����B�	&ͣ���b(�(h�%���	.(X�``f`*Tc9ed�.d�fZ�#R����CM�T�@C�㔙�`�&I�����8`f0B�S�J!�j�a���D{h��)b�)Y�	�R/=K;��4c悆���a+9� �4IP��2\�Y�AA����� � mF
LSP$�
)j㉙��J�,���������Ȩ~D�T����DD?9��<�a>@C��=���AZR������җ_s�����l�o0֭kg�T({��w��)���AiJN����� %)���R��3�m��MH$Ǝ}���9�g�>JS���8(Ҕ��߻��Q)N���┥~���G�JS��>�?��>�����m���Li�m��:E횶��sI�t�kgUqZ�'���'n���)JO���8>JR=����)J�����)Jw�w��)?}ڌ��o[3nf�Z��>JR�����?�"���w���R��;���)H�/뷙�O�����u1;�4�L���z��)J�����)Jw�w��);��w��)���R�����/�k5���l��9�p|��;߻ÊR���߻��R��~�)BHtP� 
B��"���H2!(�(��y����>JR��H�w��f����Xk5��JR!y��QdB�	�>��x�(��d������1�H� fFے@x��'�{[cђ�䓯�T�ڸSZWp<�^t��h��k|�R�����)J�����)Jw�w�R������%)K����>$bq,lng>��3��������{�y�)JO{�{��R��~�}��`g���v)ԂLh�s��E)N���R�������)���R����������K��赽�q��F���JR����{��R��~�n)JP��~��JS���┥'��ˆ+"n)>JdRNg�>��ݔ��JP��~��JS���┥'��o3�}��ٹ���{�d�m86�l  �r^7k���h�0��������ʽug�����s�˚�۞vu��9x��(cwlMT���15�:��uK�����A'	��$c�-G �EĻN��ə�=1��h�Z�v��&8�y(�fI����fF{*�ݓ�\�ns�ŧ��W:�5�?��_��')q�LZd��	 #��X��8b�6 ݱ��-ig��#Y�uWAA�v��.�8�/�s�M�;&��v�ngʶ�6�1Ɠ��Sp��`}�}���>JR�����)JOw���)Jw�o��)>=}˽�����l��7�p|��;߻ÊR���w���)Jw�o��(}�����)w�;���Y�o7��o5��R�������JS��}��)C���%)N���┠}���X���#y����O����wۊR�>��{��R��~�)JR~�����)u�3���4k[�֭ow�(}�����)���R�������JS����)JR}﹭e��"T�Iӥ�ԫ��tNnz;rMh���\m�8��q���>>���+�M�W8>JR�����)JO߻��|��;�}�┥����|��?z]��E��[�h�޶qJR�����#Ҕ���$2��Cr�����)JP���;��R��~�)��)>Z�;�Oy�<��.���(�!B��٨�����{����O���\����v�Y�!d����\�	��vx��f��(}�����)����R�������JS����)JR|z{fw��[ۛ���f�����{��qJR�����%)N�_w8�)C���%#��m���1����$��dL�^o!6�VÙ�6�۰�������6��n�o5��R�������JS����)JP����JS��}��)I���Z�-�F��7���>JR���qJR��}�x>JR�����)JO߻��|��.���ݶ�Fky��o{�)JP����JS��}��?�/��~x�s�������u�s�R��i��v)�6�$Ǝ)'9�t����~�nKJR~�����)���)JP����JS�K��h��{۽����D �A�t�Ȅ	-P��ݞ)JP������JS���qJR�sn�Lr,�E�&<E���C���"^�n:7�\��*�:]�I�����N{j��޷����{��8�)C���%)N����)JO߻��|��>����]5�Z5�zх�o8�)C���%)N����)JO߻��|��;�}�┥'ǧ�g{k5���ٻ�o���)Jw�o��)?~�{��R��u�s�R�>��{��R�������yo{�7���)JR~�����)�����(}�߻��R����*b�~�n)JRy�~3+]6��y�7���>JR���qJR��}��%)N���┥'����|��/�s�Z՚�k�$��z�ŕ#Sٞk���ƽ�ez�^��:�{k�ׁ�v!˛vW���{���}���|��;߷ۊR��~�{��R��u�s�R��_wY��{͛�k[35k9o|��JS��}��)I����%)N�_w8�)C�������K��h��{۽�[��)JRy����JS����)JP��w��)����R�����:Y��o{��F����)���)JP��~��JS���qJR����x>JR�w_F�]5�k-���[��R�>�߻��R��{��R����{����{��8�)^��~����M+]��  ��О{UeM��q�
��r�66�la^W��:�6��R��]���a;br�N��a�v�"DH�q�\��4h��]�N�ے�gTc%SV��*���4z�GY���K���A�D�#m���$�a���	���U͸|�elq���ۍ��*�\�T�`��x�秘&��;9:��0��K�c\s��.�nd9���^-�z�kp��Ϋ����p�ڷ�*��wn���|O�������M�;UJ>"D-���!/|ۥBR����K.JP��������p���I$�dnC�}���g�[x�Ű�	I�y�5�!��{J,��;���)>��3+]6�a��o5��|��;�}�┥����|��;߷ۊR����{��R����ֳ5ط�Z��5�z�qJR��{�x>JR��wۊR����{��R��u�s�}���f�Z�ȦDӘ&5�9�g��;߷ۊR����{��R��u�s�R�>������2�}���?�ִ�J6��;�"�#1�E�c�'��c,���obY�Ҭ���7Q��N݄���"B���QdB����A�G�ۡ�R��{��R�����v���7��[s4oz��>JR����!�:��ϻ��|��;���)=����JR>���t�����v�h����(}����JS���qJ�H�3wiE�"�7f�D ���H���va��n�f��p|��?w���)JOy�J,�A�9�j!��BI(���p|��/�H����[ݣ[�c�kg�)=����JSߵ�s�R�>�߻��R���{ÊR����s;�5w[��t��5�q�6�x�h[6��W76�0On�6�և.z��6.���N'�5�{�{ݥ=�_w8�)C��������R����{�����w�35ص�Y��5�o8�)C�����C%OwiTB����ҋ"D,|nj!�`}�mj�"�N`��>9ǟt��>�{ÊR����{��C��0Ԧ���8�)I�߻��R��������n7�4kz��)JOw���)J}�w��)JO}��������xqJR��O��gw��ozۙ�{����R����n)JR{�w��|��>�{ÊR����{��R���t��n�7���.�l��\IӉn�q�V;=���T�vss��kC��J����xح���{�'��~��JS���8�)I����%)O���8�)I���g{��oFn�ټ�9�sC�)�{�R����{������{�R��������)J�f�D9�D�F��}��`}��m��)J}�w��)JO}��������xqJR����WM�-kވ�k{��)J}�w��)JO}��������xqJ6ĐH�I5	(�������� �a,���,����
DEd���"<��w�p|��.�����ŭj�[��o8�)I������)J}����)=��{��R����s�R��>�3�u��z�o.��n� ;Pq6�����7�u��v�4&�D�)�k����.�nÑ�7�{�{�J}����)=�����)�{��(�)I�s����JS����{�7F�o[8�)I����#��D%$B{�J�D ��:��,�A�����`}���eT`��τ�)'1�R��~�)JR~�;�t>H�"��U�!,y�J,�A�^J��v��Z�n�,��)JR~�;�t>JR��{ÊR����{��R�����ݵQ"B�XLw�Wd��̕ڭ���{��┥'�{��|��;����)?}�}�%)M���X�$2b<2��`�f5}��.��ٚ)]�V��0��4�%1�4�YIJC��F! esv���20�
B	*	d`⒁�!`����P��Q�&`�:I���A	��%!$�Q�E�N9�PK�bZi��$i]� �H�^�y�TJg�Z�٫������d�5�A䁩"�id.#���.50^X�ᑙ,��w�t=�FD�Sx�'��)f%���U��-���P�JU0��6��p%��@A(>)�hR�0���c��A����h�k@�	�b ����8`&C�<����zd�~���-u�    m� ��E� ��       8    ��N�Ѵ�l㤜���.�+UU[m`u�ke��3����8H���i*�4��V����i��ݍ��E8�fNՕX��h
�[��� �n�2����E� \�C��	Q8�XY�mN�:TO�/_=��R�t\8�f�X��ʹ�S��^�vx�\�5m��=*�B���8^�h�6��+Hbx8����̴�m	W-Rv�W�Q��u���VU��Zݤ�[;-]�rV���R�2vp������u2�d�U�4om����,��[��ok��z��Lp���U����Ӵ� fγ���@��tvݵ�s�H���M���j�X>�u�[˫Y�ŵ�M�R� H��$��[.��#�:
��ה�X�Kz��iЉ�"��HuT��L���[n�J��s�D�Kn�V8�4�s�^nK�u��{!ns�$��{rg�24�ĺD��0ת۴��H�U��E�ے�l&�xnN/)��WG9M�Yq����J�T�p�nݺ��ܹt�����ݵ��ڪ���H;:�GgI��k��~��eLe���M�6� �&��v��	�H�U*����[�	���^9Pm���<�r�W5��@ݕA۴���L����^'3��X�:*�#�v]�5[\���I	7Ab�٫�bG-��qlYy�Sv0Eե�%5]�շBF�;[m������ŠZm;:
�Wn���h3�o��M&b͵B.%T21�U���t��!qOO<dZ��TH-�9�ݴ��.ҷj�������$PRGv��i�m6���$  m��ݦҀԨ3��0��M��W6@���s�}R���:���7v[�m��Cnz�j�����.���४�UV7`��+s��@���nB���%��J�<��]��D�9g�k�8;D���hpӶmSڧ�|�{��{����.�1����� �T��<�{�������������[mt� F����]\i��Wc<%ƭ��v���tZ�m�T�6WgkoV�`b�{;D�C��&��(�P}k�q�IJ�uV�W���Rt���R�����ӯӰ��>p9�݂�xD܂�Vk�4��[��x�'bK��9Ͷ��1��Dem�I�ś�`�F8܍M��$��A�Wi�<F����=���W�S�����΋u��n;���3�&�эݚj�&��Ђ��.�v�\ù���۸y#9qGUr��w���o37��7�kg�JR����8>JR��{ÊR��������~�xqJR���ܮ��Zֲވ����|��;�{À@$�'��k��%)MoiTB���n�Y�!�&x�ֵa�Ʋ�l┥'ﻯ���)߾�)JR{����JS���8�}���kV�ȚsƘ�8��}��~��8�)I����%)N��xqJR�������R���v�3F�o{ѭ�h޷��R����{��R���)JR~����>JR����┥'����?v��-�k�U���Dg�y���8�r��b�*H�ԈLr���l������>JR�����)JO�g~��PD'��TB���n�YK��/��n"$�����]����}�a�f�$�!*�"kW}�}�W߽�|���V̙�	��L�]]]��꫖���7��l�<��: ��\�r�,�Hpo��@����ٶl5%:�i@n��F���������>v�ܭ9�o# �M��p�v��`��=��ښ9�fjݛl@�����:W���8�uk�]��g�8��$ݘ�,f��y�otճ �kV�ȚsƘ�8t�y���݁�:��fS/R�2f#M���K��.H*�������jق�}�{ﳜ����t�y���X��n9�M]��	���{��h	����>M�U���F71dO	���� ��y��m�@��\�=[�JB)"K�m�,��$j[�����N^��K����"Q�>R#�"N?�	�$I�m�����:nprX� jN�������&�0���	�s�{��hl� ��X\�6���I;�/���{��h+f��� p%AT�	�&˒*K��ܖ3@i[0���~�3Oj�mj�	1F9�cLo�4�ـo�{�>�� �r�hnM�/�!���m���դ�[mv]�/l���<�́��a�+�"�$.-c�T�7Uf�M������3@|���f�	YnO��9�@�{W ��c4�ـo�{�zZ�%�wEU���D�us�wr�h+f�m���\�"ؓ�IL�b�w:��p������;�{���ue]�%md� ﭽ����=����]����_ǲ'�0pr1"R}�w^���_ߧ������t  ���U����"��J�t�b���*�tFpk).�ռ�׃v�������V�Y�lQqp�X�u�lʀ+��9ձqv�v�����X(t�Pt;5#ì�x�v���U�]�"�UZu�I"r�y�3C�-��=�
��x5����N���bW��ڙ͘h�:yݤ]D��=��2�`皵�m���okn�ʘ�ݻ������s8|9��U���e��ɑ�"x�t+q�[:{s�ǚ#NK
f4p��: �'��Dxa$������=����3������wn�5l��o'�9Ӳ.I��h{1ڽ�5��@}��v�6�V֭y$� ,l��t��;�{�>�� �i�h�K0��. ���0�otԜ���Ɓ}����Ta#R|'���z�'8w7��>V��m�㛪�%��[g`ץ���9�M��X�ɵO]��ֻs�����2�V�.���j�����4�� ��{�>�� |t�lIǈ�����t�)�fg����y���~�s@{��j�%29�B��9�	������0w�߷@}I����h�)�6�TTI�6�I'z����{�=�e�����X�/����(��x���{�����e���{�~���'8�*��ETM8�� �:��N!-�-��Ց�u��s(c^9q)���L��5�<�d��6cns:�e8|��Γ�����<�K0��.�����9Ҁ��w{	(�'��f�����@�l� �UYnO��9�@�� ���4��T�`������a&xqp{��:�e(�m݆Ϸ�f��2Q�ٞw�N��٘����+f�m��I����hzѼ�LPs��"�"&�"�-[��gs����n��m��n.�ßZ:�v�l5���T��ݘ���Γ�������8�ʊ�>�#�	$�@�^Հwr{��0�otS3N���l�"�n�p�Oc@\�F�m�����U��t����9�J���mP{wn����5�|���}����T�D�q�#	�ɜ����t��ܞƀ�<�Bj��5d\Ĳ����{iA�a�h�:w�:�y�H����;p΍��#�V����S~~m���9�;�=�ry�������e�E�]@W8rx�ry��ށ����_�؛�2%�>�����=ͽ�<�9�;��hZ�pNd��I�I���m�@�^��=�@�m�p�5eD�mᄒn��I�ܞ3@\�F�m{��?�ȚU��&  7k����Wn�����@s�R]��:���V�v����>�3ݯ��ܦ��S���/�'[�7m�I���Cu����j�u���Ƥ�գ�����5֞�3Z�z�:��c���5PrF��Z�6M�7�v�+��"G.��j�v3�9�nklquX�$�n�5r�p �[�=26%:�!�6�c�s�����s=�{����r�̮�?��q�l�a�Uڞuu�gi 8�k���J��:�:P)�"�g�b�LTM����o�����=ͽ�<�5�*�n�I�c�6\�]we8�ot:np�i΁�Y�%�7up������Λ��Zs��g ��U�#q�I<jG;�?V���ӝ I;�7�{�zZ��v[cd�'�$��{�6��o���[{�?W�p��Ͼ�v��x��SF���3.I���n��:V��pva�m�����D�l�O"X��q~ ��N�[{�?W�p{f��*��:���n<\��/ͻ�㒧����@^>�� ��8ەarO�6���I;�?W�p�i΀.N�����*��u�'��R�ٵt}�p��ށ�� �Q�d&��irqtrw�o&�@�� �+Nt<�V����\��n�Ga陇	��(ET��&����nznoa��:�k�����V)���{`}�v��u�����BJ#����w?��%��H�!?�����e8�Zs�.O# �M��nje�uEE\M�D�]��Zs�.O#��#�Ȏ��@�0��$�Z4�f�P�`���+�e�HY`&�D �I`S�po8���,�H�_l�� � :@$%	a&Y%�IV`�P�ZH�.��$O��Kc�~`$����&Q�q |/�@ �~�AT���@�����Ci��@�;}��@�YN���lNF̈yD���'��o&�@�V�ܭ���u�9R&�A9������e(��nl�:T��&_%pS���ʝ�s[��h��t�X�Hq>�MGk6����6��Ц5��021�xa$����� �'��'��{�{��*��u7WU1Q7W8�<f��<�ܛ���NV�uئ��iNp����=ɽ�<ճ �'��9��d�AH�O�����?{m�@�^��?{o)��9�-��� �eZ	\jG1$�jJ��<�9�=��4��`������<~�h[�:�JC�Aqu��L�k�v.8s;�3�����s��nKB�L�#�]������0rot:Npz��Ȝ�ŉ<�Q��@�m�p��{�?W�p���t
��pQ����I��ܛ�Γ�ܞ3@\�3�[sP\�G�Iށ����{��h���;�{��&i�3d���us�{��h���;�{�~��r��d%"�Tu)�BZV@�� _�?�����՛�k; ?�ﾣfJ�Α�w�f(�Ӊ|FN#]q$˦���Zâ�q7z��[k#Y��l\��{.(�C[��F�u��nu>y�ݍ�v��n�ν��!��\D�v�qϣ�B��d(�Nѻ6��܇c;3�gv�����[���v���ї���	��:��sW]X���0)ۚ�x���Mў��W��N��=�w{�����~��,J\i-��"���6�ِێ
�8�Q�j�I�mtOg9��#��Wծ�5�˲O�f𿇑�w&�@�� �o�sQ4�D�q�> )&pz����ڸ�o)�7�y����A+�H�K�IW��'8sx�rysot6TҲ&�Qc�I ���:�o3�{����ڸ�CQdNF�ĞI��@I<�����78sx���q<RF4A�B3�rI�]n��E�z픹�r�4������P��l5SwM\`ͽ�<��;��h	'��w7\�G�Iށ��W�(J>J�Q�n�,�:T�ۻ h�q;q��ɋ�����@�����������F�L&9�`U�a�蔞E�����\X�X���N$Hԉ��I3�{�����0��I�`jd%��9����7i�PnÁ��3������F|��&�m���)&E)�HɈ5#�������4���;�{�y��]��L�vD�3v`��4���;�{�y�N�P�Y���'�B���7v��^����/t�
�~Q7��wەn����c�	�$pRc���=���nـw7����5
A��UPAww���`��4$� �����K@�%�#,�m�L��L�,-퓞t4v�^DS^�n�b�q��nF�xdq�9�[�twl��������F퐘Lr��wY��$��ͽ�<ݳ �o�~���� �a>o�I8�m�@�l���3@N�z��aWsS3�M�^��� �o�'x�8�=7e���2���1��A�� ���hI�����`ÝS�J�P5ۜf�e:5��\�m���/V���n��!�M��+MLv�7�~l'xsot�ـw6�4-A87 ۀ�8��޶��[��޶�:n��6�j�`c��,0�M�V������xsot�V�����$ԇ ���΀[�pz�ށn�p
��Ba1��������O# �m�ڶ`ͽ�$��w�}��ߏȓ�&�H  M��X���5U�֌a�uk���k���}؁o9�y��s��s�8��nkVC0/l m/!��'Y	�V��g��؛2Nõ��pn�*��ՍR��s;t��RSYн��1��O ��'RnNʜ[bİݳ�wtv�úQ�k`�9���ĖX9�i��U�Bn��3� ܳ#���2�[sB����oD��m�d):�gUF��Th�$�m���M����Xt�����˩l,*�����]"�h�Vi����{����vy�P�nՀ��g ��5PU�8�K'�H�z�)_�%2fn�u�*�m݁���<�c�<xҐ�����-�����ށn�p�sP�$�8,O��s@m<��7��l�=ͽ�K@X�ۘۀ�A����{�-�N��v��Ҡ6!7����I9��vy�bRy��kŵ��:դn�Ad�6���.K
f;Y4dY1d�01�yG'��Y�psoc@m<��7� �s*)���@oV��f�r������ >��'9]��������p
��k�<&I�
��� i;�;�{�>v����tۨ��A��?��p{m�@|�soc@N�z��E]]D�j);�/���{���@����=�oz�Z� ��"�$�r8�I.�۝uٝ�>�n��z{\5�7��#�^�g&D�1L�7��.�[{��o3�{����p�sP��$�$'�Ĝ�t��`ͽ�Rs�w6�4-����2I1��ng �����j��Ŀz��:�ڸ��ŗ$�7�a�s�`?s�y�2�~�9�ԡB��=�� ���+��D�&O�#��~��S�_=��{��ށ|��w�U#Lcx?���q��nzIKp�$[<^��hQ��X������h|��c�6��:��8y7��NpsX����L�e]ԗ�T7s�w�{�>V���3@�{W ��(Z�q%��);�/�� �5���u�w�{�y��i�i��F�2H��]�:^���m�V�nSa����Z��g*󻚅a$�xD)��m|߶���p޻�t?m��5��I�;�i�G�vs���<�NnR὏n�[lqx�W֎�	 ���$��H�|߶����汚�N�����ส��#��n�~�9�S'�]i`l��P��@.T��dR<2c�.��yM�'Xy7��Np='*w5�;��� �{TXjP�y�y@g����ڸ�]�:�QQĤ�����w�{�>V�roc@s����ݚ׉KD�}�`��_*
�4%-�~�iBPɂ���6����p�	��Sn�х�H�@�P�D	@�0L%`U\�q�%<�/�k9�PV))3̨IL�(R$$��j�G ��+~��"�h�<#
"��l�f�BD'O ���%��N���5�g��%�i��yr�������Po�dJblC`_�D�E)F��
�lT���lh,j��ʌ !�s(*�r�A��c��f�о���`���?I�*���IjٙefLEc�3D ���h� mj������k[��   ��� $�G@ְ     0     v�]^q��[�`*�mxs* -�Md���6��m��;�jV�=vP���Ʃ� -
�8{]�:�vsq�K�
�X�l�ə:;�7R���Kog5����i��8��\��x�^�>7"���8����`�j��WU/c���x���sk`3�FTxv�rl�<I�kpɐ��yͶ��Jg�����N�{p�
�(g[0�R�6�uE�KׂU�vmSQ�I� \�7\�:��hc�TJ�9Nۥ��ګ[32�� I�e��l�"Y��Y`�*�<e!b�d�@,�"I��t�ܯ%�i�ul���vhLY�*ݰlP6�:�@��%�Y�;t�����k*��` �m��9�m�j�y7mΤ��7]E.c;��ہ�V�8���JM�m@�n�u������KOBt����f^l#�I)�m�cnA�ݱ��Eq!��Wr���J�c��Z�y��"�R/��^� �K'�^C�n�W������)�q�3�
[J�muUN3�Z����X-ѧH��(�kBY�`��U"櫶����r�T�]��.WBɶ�$tCf�'B` UT��vv�D�"�*���Wom��&�WUS���s����p�[3���eZN�#��Ƕ�m<⪜�2����"���+g��9�)g�[���g�\��taj�nL�`Ms�!n���)��4�UP�]U��5V�:ٽ$�D�P�]T�չu��*��,�=��7m�6h�x:ٮ��D1�\K�Zp�KJ��U@�iw��EZ�$�PZ�F:�R1n�)Z�����H�P�x㦲5bY[nݶċi   6ݵ%V׭�ʓ ��Im�ݙ0j��� ��$u��Tr���9�OT�<��m�T�u(��T��	��� mmI�Ӓ�n*tlQD�˗˘�[��r��§��g�����k97H�bF��n��^Z���e��P"m� H���4'ϻ��������{�7W�V1d˳P ђ����ܭ�Unͨ#K͹�w1����n46��q�3��5��tR9z��s�n���p��kX�Cm��i`��YM+���l��v�Ob���lueQ�c�ە�[u��;�V�OY�⪞���n{g��ܩd*Z�<�2D
��󺝐�W\���ΐJ��8��&X��6��Lb��"�
���ŗ�ׅ���ӯ��3uʭ�d�Ӵl9�k�n���;m��u��R�㧝Ւvs�.q�0Q�8�F5��[o3�o���@�v�����:4���I�QTI5q�.M�hRu�y��@|�F��'r)"�D�Nw:[��4��M�`�{��wwWe��T�]��`i��<���&�4JN�NL8��**��.��@�O# \���<�9�<�{�~�#�rʪs�߉��卆L5�����w�=�N�xC�{+�ub�:rh����Q��.\7~m��lh��`i��'��9�9UT�$��Ng@�{W/ٙ��̙�Y	
������(�7j�DDD)�o�?�ĦG!2|�$�\��������&�4Ԝ��0n���䒾��{v	N�(�vՀ��s@|���ێ�'r44��� �m���'8�ot�ـ.�UD�K�M�m�aqsms�#e��od3���[pnèmܑnG����NB'!���xt�h}�݀��s���{5֖�`od��$�I"�����_l� �뼧@�{W ��Յ�>"Ȱ�9;�'��{��i}[v�������[/�H�%1�9��������:�O������������Q7e���Pw�h�9�;ɽ�'��~��S�jU�r45"fF�\����5���ڍm<k��]yns������T�����%"����ށ|�\����ڸaCk��M<QIހ�����3@j������"d��i?�9����8�����.������{wn����@{�0�5ޜ�E�����7�h�9�;ͽ�;f����2}�s3��v���-��1�	$ƞYws�w�{�.v���f�Γ���3���R��!�4C#MA2�@�Y�"���HԊ�Y��|#9��n1;�p��	s�]^̕Qsw~�~���w5��9�s�{��� �^;�S&0�	��C�{�i��$�d��٠3ۻvy�T����^)	�6��:�ڸ�[{�7��8�w���mk�H�'ɂ���;ͽ�7��w5��9�s�o�2�׉�0C��������]�,>c��6�����(����鉥k��` v�X�m=Z�|���Si6�\�㴊k���.3�����<�8Z-�v����Hժ��*넄�u���IJ�u-�|�l�jܴn5/�X��Ҥk�x�;�
-g�Tjt��ri��\�UQHd���Y-�:{��8�,�Y�y[�9�u�;n��9�u�Rvɉ���O<���6����&���	����qλNg�]�t{��{��ͻc�Ƹ��7^�t�·Iv��3�B5fn�u�Sp���s�V���7I��G�5q�$�3@�I��m��h���=���ّD��S�:�ڹ��ٓ&{wn�y�J���)� ����.s�'&�$��{��ށ������^ݔ�9�s�%Ц
�
����j� �%��w5��9�s�km�4��U��U�EU� �X�9�s�jm���/ߪ4��n3rdM�8���Gn8s1�D۳sB�cY=��mq~}fy�����PT��:NpM��7��#>�Π�o?�����q)1��>LII8������9%��9�s��P�IV]���E�����X��ڸv�ށ�qѤ�F��������9%���� ����y�ۉ;�2C"�%1)��ڸv�ށ}o3�{wyN�|7cNc��X1c[��kRfq�k�Xko=��$���{��.A'��ș���NI��I"��oz�y$��T���)��q73UUޡs��n�~n�j�S&6�K_�xۻ�
"T�{�l����.t��U������9�a.��^Q^t���[���������1c`Ԝ���� ����y$���'K�<�2)�bJE�;�oz�������ڸwRpN���ǐæ��)���;.I݃N- ��s$v�Wn:�1�a�hp�F<bs���g ۷��^��-�{�?n:4���Ә�h9Ϊ�t�ԡL���h׻v�t�T(P�G�T�5s���<�����`k�٠���~n� �:e���!��'�D�I"�����8���(HJ2��������QԛnL1��z��� n�e:׵p۷��K@����a�UN����`��;�bMsv�.u�X��<���ũhbncf�11�����:׵pM=�7����:��..&*����@j��SOt��`�c7�}��ٟ${�/�\I�q�O�R.��_���F�
!)�x�K_�!\��� !��D�z������:�c�P�B��^�`y�iɞj���y�U5Uq�%��5I������r���J�=�����՛�f����� 4ڤ�^U˗Z�v@j�g���4��$ln�Uz8��nvW�m8�������"Y��7����| ���&s�gf�3<K{z}�fͲc�*Q�ɰ���^ݜ.�n5�EW���8�1��J������lk3&�4S�4�Y�˹�q[u��=v nNf ��6½�N�Vx.i�a��M�ve]����Rz�&��z��~�V���V��h
�� �ӗͼ�;��e�`����Jg=��nnj��p���Q�7y�ho��Ҥ﷔��L�q'R|䋀v��@|�F �,f��'8qФqvMɆ9�@����7}��@����v����bnb�11��.X��Npm=�7���)��E2b��rs�@����v��_[����S�~��
5c�R0�n�a6��k+p��z^L��5l��w@��V���9��Rc��|ؒ�p۷���Tg���	%�=��!j{�9ӻ�5F��5�<����9���Ks�yRs�ki���d�7155tQPW\��T��A������������94�(�;à]z� ����y\����)�D��Ϝ�p��ށ}o3�{}��@����E~l�4܂��(����3c�D�usH\9R��S�,)��a�~o���"2&��n9΁}o3�{}��@����m�@7k�����1�bcs8<t��JT���h�^݀��* �ǵ:���,l'8t�j�w����}�==bB���v�s�M(Vk%��@�a��UHH���)��Y��BQ�8R��;�lG �x"@)ȴ����즂Y���)
	! C�@�B�@��(�I��D�=<U�=XU �A�
侄�{o�T�������Q'z����Q37s�i��7��6�3@i�\�����BA&����y��׽��5�������9H�{�*�{j0��WX�v\���6�sk�r�a�GȽ Y3�5�yA��.X��Np�{������q2��9"��‧xt�j�����8�yN��L�pm9�|��M������T��	ǳP�LDM7&s�/��pv��Uߵ�s��G��N �*`HqJ{�����ʯ��nֵ�Zb��
*�0��hRs�&���t�IDG��9�y<8s�v;ؔL�T����ɴ�t�n������q�C�Q� ������s�����1���rs��?��ˀ[���_[����:�G�d��Ĕ� M7�@>o# M<f��'8�
Z�$����;�/��p�yN�uڸݷ�ێ��TX�rx�0��hSs�&������0��J��rD�lp����\�!B���߾��T<t�bKx����YSk�� 5�:�tv�nӪ�N�l�v�k���F���rX�<��Qֹ�x7�:��cm�^��(�ӂ`�79�̯	��͍pv̸+eA��9��g�4�a���ؖ��S��s�LŪ�]��X�,m�����Q���
�;���D��:�,/-EKd�Fc�w:��L��)q�^�ڐ��U�x�ףC��z8����w�{��sڲ���`�x�c��S��t;��f���K<c��i��k�򾶴;���>�v~����.�p��~�&�0��h���6�q;��IɆ8��@ݷ��1�X|nhx���S	Hno7��G�$������s��]��m�{�.����ښ��2)����'8t��� M7�M�`	���<�h�b�&5��ē��m�{�>����o)�.�W ����"�$�����O];�#��mgn19wV��D�<�iӳ�F�La�$m�	c��ӝ�m�p�yN�uڸݷ���HuE����QU3Wi�5}}�����ɽ�m�p��J�s�!��B����� M7�}@4�F �x�Kt�8�'jA�q��6��m�p�yN����uڸ��n'rbi9pE����yi�4���M��yeZ6�3\S�/��>R$�XX$2���l:u�p��{/]vrrƍ�Y[�ۜ�bcs8�yN�uڸ�o~���v�g /����#�<ors�@y��o��t���,��|�h�b�&5��ē��[���]��ù�V��N�uڸaM��A��xT���M�`	'���� �m��u�:�x����i9�wo)�.�>����@lB�I/�t��O�l�<]ۣa�F�َ6�l�q��mx�èm�-x_kC��5��7M&W�����k���cn��Ҡ=��N`�8�7ԍO��p�m�L������t���6�q;����st���9'��np6���w#jc�L������]�������.*D(���a%�ʀ-=����a�Np�]��G������0��h0�;�&�/h���ls�V�;b���F��^�rN���c,�N���9�Ĳc�)&5��ē��{������t��t�ĈJ�k���y=�Q9����@�o3�n��:�\�<n��)P�I���3*I�Bx���4��Kt���n%\�b�%�<P��uڸ���]��������S�j��)�MH�����7�m�`��h�s�Gw���~?"mr[d� itv�7�����n��.ט�pV�ɝ���^�����z��urGg�-�J�����Ks��Q'mےx�V�Yj��v�#S���vr;O�N�q��w��4�qY��q<.��CU$n[qͰ.E�ɮWc�e�4K�WGcn�ܚ�v�W��+m�Ҭc�D����;=Z7>b�ф����gRj֣m���{��im�t�6[�M�N�h#�ծ�ms�.���]��x�`�Ӻ3�<]�����}��& m9&/������p��S�Z�\��{��yr2b��LNe��L��s@|�n�(I n���L Lkrs�@�ڸ�ݛ
ν�Tǵ���ew��y=\���3���P�	D�^�������S�]{W ��)���R`����t��`��hRs�y��@��n��~�Ŗ񭽚�n1h�]I�Ͱ��ۍ�����ڱ��=�wt�������US5q�.O�5I� �7�{y����)"X�#�>����_�jR��8�n��ݥ@?c�X-�#cr<p$�����ށn�g ���t^��6�q;�6��!w�a�	(Qۻj�&��i`fs��oz�^\����<�m�����J}{4�ݻ��*�ڊej
7(�F�"R��\^��n�Ƌv�%�sړM�mD�9�mt�}j>��{=uU�a�%M� �7�6�0��:��$1���ƒN.}�����6�0��4���7�1:��i�>x�s���g ���t�{�fq�0#\t D2.�(b��|C1@4$�sT`1�6�(�?��9�?�?�.���oz�ti:�x��1�&j� |�3@J���ot6�0�+1�ƚ"��������I(�ok�=����:e���s��n:h��Ń�֭��Y:�t�l5��3 >�m緑݋�I��6�2e��j�@?f;�>mҠ���,�c�n{7��jI1������k�X��4�1���=��ruO`\]��s��~{ZX��4
G�1݁�����u4���E�99àfs�<�vͺTQ�)(Q	�}��d�r�t6��ȈLI������{�y���sO�%I�����e�N�󷣬[L�Ö!2u�ѓ���Xjۊ��+�qգY�K��RF�/>9�݁�n�玙`fs�BJ ��J��ӈǏ��뷔�39�h�n��t�BP�9�j9�H�4��xt׵p�������=v��i�q��F��a�<ۻ��*�2�Q�39�h���n�f�$ǐnw�~��8�:e���s@g�w`~ȵ~�	H��ST�$00W�1�Ƣ���BhjX&RB �H�YB"�U8T�rִ�	��g�ӡ)���� �b,%�0pd � �����RG���
�(K(B@�	$��: 0\Y!Y��S�fT�U�m�@��]�g�~���Ձ⃄!�y��7�o[`    ��  �����k   0        *��w	+z�=��1���F*j��y�bp ������X�pE�eg3QsU!hU�T��\FB�,�H��d�Hz;U�n��OF��8��oa�1-v�Ds�Q�
q�̓k�8R1tp5�;n˃(1���(lpm�̭z0�zL�(g��r#κ�X��m;R���$`]1$)4[��t�q���ݟP� �T��R,mtU<�[WK�Q*UWf�.�c��p�\�f���ml1Ԩ�4���)� $@ꚪ��%�͝@K,�Wr�eM��%��b"���8īJlJ��n���<<�&��S�[m�[@F�\�$K,M��.�#m�� UB��R;�c�Q�nnIֹٹd�N�mk�RfX*xM���m'Ol5[����B�C���,���v�6�5W[;u�x���ڀY.����������m<-=��Zݭ�V�lv�=�[jg9d�ñ"tm+�lK�T���ֵE��o=kB�`�P�-ڵ6��"U�4��e^ɩ(0u�-je��yڕ�8fƝ}o(�kY!y�:4$q:T+r�R��Px;��  b%M;]ӡv��V��:sV�yǮQ��Z�u�g��i�u <�{OEc�<G�7��MS���ښ�x6v�L�ch�Dz2�@��w4�Y�e�%Uogf6-X�L
���3�ʵU[����5Ҳ�Uz�2��½d��G$-餒ܡ�U�ڤ��/n1�\�B;M�PPw@�2�V�9IV�U�Z�
���q�LUU��5<쪨� q�m��c�&�F��,[�l�I5�Slq�ݶċi   6ݻl�fܛ[f$�5��}q�`*��켔���R�V��C�.�S�<�n���z�=l*�e���� ��V���6ݮ��qL���jx"��#�|j���Y��] z���횯<V��kF������E��H����?�i�EL0 ����?��������՛�kVI� !srV�ޱ�����V�K�$l�8�3W6;gXh�<mQ�wM�X7-NE�Vi��n\Y�p<`�N�ql�\�={<�y��.��5�H�f��:�#A�����϶�uL��n5s�ӷi�F�A�m���<=��\v޺��1Y�N7p�seu���F�nx�����D��0�Y�1��G���g7L�;#�ww���8�4a��J�Ӻ�l��6%ӹ�ᇲ���O+���ccS���s?����:g1��m�(�J���J�<�c�$V,#0YNp��j��oz��8��S���}���Hd��ě����6�@m���x��np���r{��Bg��9�݇���Tk���o�����n���2������cǈng ���t]��o�������n�`��RdBd� M�[��`����onE9�������i�L�h�o��{�?|%̎bR4�@O�:���7���ۥ�.C5�i`zwtGy�I�t�xku�o9W������iF$���)�N��@?<�X񹨄�myb���mI&<�s��y���S�Z�\��ހmY����"��p��|nh����6�* ����+��<jNp��W ����[o3�]��tn�
5c�S!0���`-�b�Þ�2�RK�Ĳf�yc�J��C�}��s�R15�IH������0��h�s�o�BuU7SQq3W�U��yI�4��<����ʉ+Ti�F'���;�x��74(�ꈔ�B��w�f|���v�8��J��i�0o	�}��-�s@}���ۥA�����,N�#���'H��ݽ���p��S�Z��v���1�i��u���!��h�rq:���Puϸw4k�K
f;XMߝ�8LL�&A��I�s�ݔ�ݴ��c�IE�y��`ej�j��J�.@��� Ԟ3@n���'�{y�� �2�hV0���XԜ��-�� �I��y��0o&��LI�����~��ށn�p�WC�ٙ��|��J��a��ڍ0�O�W{�6���m΀�'8$���k|�9�RD�_<�&���ՋnM�u�m^��9��7.�»��
�8
$y�cTL�v`��:t���{�h�� ݻ�X8���Lg@��\�
d��݁���x���>��y&)'�@P$��{woz�)��>�>�g�ݛw�f�m������9+��W�;v�S��J�ݛ�c�G�2��V\N�S� ڐ��-]TDBIn����۰β���D%2��Pr�C	=~�?��萛]   �1Ɨ��p���+,�d�u%�_}��|���Ū-��;����q��21����Kv-4m�:�f�{�Fw�@�RZ��1�N����f�lkv#S�j�a�3�7[pt>z�L�g�,r�WR�v1�l��'�wŐ�i��$df4Y���r�xH�v��L���tp��de�jv�[lЮ��<m�qn��͓��)v�=��v�R_�C��!��'�˧Ef9c]-�xu�z:�ܻմ����I~||F>��vz:���`
��8$���fG��m΁��9��<M44�qpn��@�e8v�W@�ڸ}��[iE"��*��@m�0N۝#npI^�ʉ,�&�!� ��j��s�rI���6�|�]�tO:�.�r�S`7�����߾wg��;�Z���o����F�A����\E����7=n�����m���9�v^��;bL2I0�d#ƠI ����vS�wl�g��-{W ������6�I�;vy�V�(�D
!(����ݛw��@{3�9MO��J���*���5;nt�9��#�Otճ��򸕒$�<�$s���Z���'�jـjv���������M44�qpn��@����p햮�u�\���pq)$��P���:N]�ʹ�u��/��메���]n*	�ls�܎��G&�19;�/�� ��j�^��=���ʉ,�&�!jC�^>�7�DDLD���hm��Ϭ�6�.+�'�����^��=��症?���/�	�T|�]���p�z��~Wn$�I2
@�,�����`��:T���q�r}#Y$����@���햮�we8�oz����ŗQO>�*
�Έ8A�O�vj8�t���]��4h\��ϳ����0S�$ c��l�h+f �ot�ـ�r�5p6�ȲG98�ݔ�Ͼ�����_YN��W?�ϳ�H��Hcs �h���(��v��(��̀�:��eT����"c	��?�ϳ3�bJ�֔����3����HP�	�@\��'7�󿼫�홇��kC$IjC�]���.� �m�@~}e��(���uO�:w�8ORgv��y�][um�܇9�{cǎ��z���Z�w����s ��y>N/�[���m���S�]���?+��L��73�]���_YNv�W@���Ͼ��3 ����rd#y$�����`;nt�� i�� ����%>H$ bs8�-]�e8m��HP�(��t�#�̹�C����������ym��'��;e��ngۖ�I(<M�I$�I�o$�[����U۪��8G�k�#��1���Ҝqmʭ�v�lk'n8��E�ۙ��u��W�!0b�eq���Uj�ڦ9��u�:۟3�m��BX���2�����n���6m�$5S�'M�ܮ�1�
�+���i�r9Uy�1�����s]w&)W��J΢g�2V��l)gX;=����3�q�s։�v{��{�����q9�S�Gl=����%��r�\��jN�&uu���6],����u�Lr,N}m�����{��?����m���ϳ�΁}���;쪕�5$�%E5{�>O# m�s�>o# v�ށ�Q%���2D��&�8�W6�t�"�Cm��c�@f4��8���0}�]�o3�[m�@�����j�Wn$�I2
4�.uP����%J[�mP��ٰ/��p~V� 7Œ<k�bI�Y�]6�h#&B�Y:�x�M��
狨���L�L�Lq�;�.��pl�t�y��oz�f�w"k 19�+�����~l�$%S ��$!�!���&5&
1�^��h@�����������O1ҭS ��S�xO9��\�;]��77iP���y�� ��s`cg+��D�M!I3��g�[m�@����-���/��p�*�m�7&�<SW�I�`�nt��`��@��n��~�Ŗ�5ݫS	��sqm�cqiV�6�c�ۜ����Վ&8������}ΰ��$ә�-���.����{�.����.+�0����qt�Ҡm݀�To�͐���vHLb�P��-���]��Ù3OE �d��? H�'N��/��	I!�i���'F���$Y�f@� 3Z�� ?�X<���3H:��c0he��^(���x�? �@��������������.���Jn7�2&�p������0ݷ:M�`@�otv���O�	0�ۙ�-���+n� �n�ۥ@j�0i�y='���5�6�.�������bu�nX�VU�B���'��qa2/܆I��M��ȟ9�����@6ۻ�t���60l�ub�6�HRL��{�.����j�m�p�*�m�I&!�$�zM�`�nt���m��d̦�<���uO�'�T�N��������-�����{�m7��Nd��
���o# I'�M�`ݺ�����q��,�E�1���u��΂m;������#Kݯ�W[sM�3:pH"����j� I'�M�`ݷ:�y�iM����D�$Ƅ�z�iV̟n�vl{����v����:�>H$�ng ���.�������� ]2�&�Q���"|�@i��$��7��kv��	�e>,��Sm
I�wv��gٙ�ٟ�vՁ��wf�x�*#�PB��!�A �82�44J	���ʘ#5߻��ҥ�I� ��ޡ�6��Y��z�@M�YX{e��6�D�dn���Zp1v���=o@ j���o��ak���-*�)&+��Wc��PO�m}��;5�nglg��팺�δ�f��n��*t�Y��0����/d�y-e��ӑ}W���8��Q��=���z�t�I���؞9m���jNk/[ly�GJ��45u�K)`8k�}���w��w{���������6?9��Cs�{Z�H'�:\���M�kg�ۉ����;Z+rк�.JI1�rn�������W@�o3�n���ʉ,�&�&i��ݷ:M�`	$�@i�������g@����7woz`_[���Z��v�H
DĢ *��I����[��@i��2���ǌ��I�	����8m�΀�yI=�=l�$�ʲ~��j�N�w/kl˻!��g��űΞWՋb#y29���	0Ɯ� ���O# I'��l��jJ�ԓs:ӽ�s��*��w�4 pXP�F�	 X
T	 �����{�rv�[��@]N�cqdQ%1��$���{�.�N�}�D.G9��wf�׮�~NY/�&{��IQEL���4��m΀�yKoz�D�[mC"�5!�/�-ZM�`$�@i�0	��d�\Y]��`p��՗h-q8s�;r)�5v6v����%��4p7���c�3�ݺlp�}6��P3�Y�E�o���`y_�2II�J"s8��ށ}e8�e��]��ϰJn7��1C�\�y۰>��>�6	D%HID�`�����{����s�H$�*j����:M�`$�@i�0�P�Z_E�|�@�o3�	(O3XY@?�[�[s!5��ܖ[�ݶ���b�z/�9!�ZtI�m��v���t-Z@�Yc��Uߛmm��Y@?�[��t���d�Ĥ��''z�)ϳ� ���t�y����@�#-��уĪn���s�4�F �Ot�ـ[w`��'���>�33.��r�����ʻ�wە�*� I��HQ�>@7ߵ��*�ߺ����{��t'�T��v�$�F�֖�z�l��P�%���8q�q�vCN��ϖj�h�;/6�<M�����g%�3�����{���/�-�-\�o�6;f ��9�O# M�� �á�d����8�6��wo3�]����)��]CEhY_I�|���:T7���@���:g@�:��ȢJcC�8ݷ��`	���O# �B�K�����C�Г���S��g�fm�)�.��p�oz��>�2�f� �M,r MF���6��U�\���LRh�4�۱W$"����;�E�G//gB5![.vK�u���6һc<eJ�
3�ۊ�'�s�h�,�e��؍�ga7Ru��NTi�h^ɑ�M��9�'8�lQ�=��nSq��l���t�#t�{��}����E��M\s�^g�	v��؝��20c�un�ne4f��5DK�����w������{����ަ#1�c�N�f���;rm�;mJug7\�$�r@�)��s@��a�F��m������*7v�t��52�s�'���:J���`<�J�"!(7v��0��hi��vw�LWi��7��&�3@i<��M��7b�1Ȝ�@����6�X1ҠP�P�x��9O��ت����J��4�I�`	��@����?]Z>H፷~R|�HƤJIbk�zK������H�\n��֌�Iq�z6��w?1�$�U?\�wy���yi��7���}��}�m��t�n,�$�c(���4�뉒y��4�I�p��TU1)�<m	9ށ}o3�c�L�(ID�t�x���bo�3��D�s��uP~(���^��,oip�oz����ۉX8����5�h'��&����0��h_Q�VcpJ8�1 �Ș�HH�ݢ%q��n�ϭT�ݸ��9�痭������p��n~�I�XL����m�@�o3�m��\��� ��qكpmE"����utg���1�@c���J"w�3Qr��4I��3�m��t��xr�$VRAI6	뙟g�G�v��m����P�V���Q����1�@c���ǎ�BQ�a�o)�=��Ȳ2 &1��� �ot���O�&�F ���m�*������]���m� ^�u\s�آ�G1Ψ��F�<���<g��t���O�&�F �ot��-�9)�ccs8ݼ�L�3��M<�4��	���.N&]�tM}]Y13[���yi��O# O��~�zF�ou���͖���"*1�w`c�J�ǎ�a�R��Q͗����R���� ��ND�zݼ� �x�4�0�{�t�Q5SD����;�ը�背��|�pi�6��|�m��@��!D����7x�cs8ݼ��玕���(��3�Ҡ𱡪��F��a$��뷙�6���y�n�S�o�+"��K"�}�1�w`g��@�D$��2���������bR&�x�I9ށ����O�sO# M7�H ����.
����0��h���M����U��G>�����p�l�Lo-,h,,d�� ��5��F�<Qx��ՙ'.xa����~H�+��FI}$_9{��=XU�	D� �A1���`b����CP�@�$喖��3�#1�1�@bZu�s2I�Ў����bu�Ê���*H>���k�#o��?�?#n�LH0��Lp �%G�=�g�֛l � ( ,�G��       �    몢Ţ9�ųJ��m�N�����-�N�]�k�E�ng��.�+1PUU� �z�ݜ�84m�x�GS];F�L�j��7U�"v$4W�z�[b[�IX�<i&M��]����D�ź"��঱b��R��R�wjg*��x�]�G�t;�����5�kt���:��ZE�7Y�e{Nt���7f��mб�6zm�.�,tV�x�z�V�U�*y���5y��u����
�衵M�!�5;!gCC�j���S�o_
��c���ɔyH�F4�N&�D���j4osnUiH@����'��)SJLl��0?�~��ҥ���l�ᥝ�HƤ�����U�T����žp�"����-��gA�^@6LFӛ)fM<յn���;U�ʾ���m�`x�fX9�I�u��̷Z��Ƹn�펣y|y�e vM����t�r��3r���
��2�$�]dVh���j��vu�v��Ԗ#{��ڌkv�'�ƙrɐ	uIT�iv�c�J8�F�n�� Y�VS���kem ��۩ݞ���.�Pr�t�t�݆�  ;A�o:ۣv�ih��L��3�#6����U�p]��j/XP		ԥ��py�C�s�3^�����	��׭n��)Q*�b6��wm�l#�qB�Hn��v����!Xc�{gHJ�U[L�;�#�@յV�/a��r9U�yV�m��*����R��W=��=���loZ�����/8ŗd�j�ZU��&^@)=u�j�����T�58�+=���KV��\�m[�$��k�T����  ۵�f�l���UB8'���,��ݣ�|�b�U���YvT&�@�^i��<���u�r�λ��IZT ]��yV�����q�b��&��]R�.l"�輝��2�F+*�u�,��h�kY��޵����f���O <Q�= ~EN "���?�t*~;����O�Q��>�mt�  �ιە��W]�հ/b��)�F����۠ܽ��v��u���Ä�8㭓���pv�8�P�*�̬���3Ƅ�r@P��ݞ!0x�e�C�=��gC*eݸ�8F����5:�l��w8�ͷ���R��lsR��c��:�����S�0Ul������Lש��t.���q�O^=pmڷ��[;~�{������c�?V];�����|�,t.�pq��]�pn�.��-�O����w������*⦾����������F �ot��8ݼ�@�v�>dd�""`�� ����HJ"&G���������J�g�}�i���$�`؜�@�[�@?��,؈������݁��Z�s!��'�ě��/�@����/�]��(~n� <�9.xL��&;�w��,��P	(�o~�״��^S�|�����Ȏ00�x�v�:��c�����q�KZ��ݸ"w9���-������	���*��@����i�`��:�y������H�!�i$��@~n�~(j(I�B����ZX�Ҡ�ިI(S&I��w��9�\��p�:�����o*�1݀�:TǊe��xO#��t�3ˢ�TD�u��o�����?'��<� ������.fl*�0�=�O# ~O�7���?~kv9�H��Y�I�cY��qj2��h�[�]�6{��Xr��k<�˄$�`؜�@�o3�_�yN�n�g>����ށ���̆7&&c�ۙ�?'��O# |����0���eLt}w��i�`�{��F$� C%��N�9�s�K�������Ec�Y�(�I�w��TD(!B����״��:g@�o3�w��1)�<X�9;�O# ~O�6�F �'���O��g�=[���J��c=Xu�ey틹(Ş|�:���W��'��u����E�M�.j� ~O�6�F �'�i�`��[\�	�v;Γ<�,�ҭ�7۰7^Ҡ��ͱ���c�vfzW������@��3@m<��M�`7I"��9އ�������{ZX�A�P�MDB��X����2ܘ��ng �������v��v�8~�Qģj4�f�5;��g�;n��T��b-�.d���Y�����s�h�Xb�B)'8tv�8������&�3@�r:+.b����(���0�{�6�F �x�������������1�	��vS M<f��yi��9T���u-ǍbnC�m��tv�8ݷ�ݼ����bO���'��t�,x�X�@c�L�*"P�������[   ٻ��6T��j;)יCU�(�쳸��mHy98�,ۛ��f�P{.";�jnD�r�E�r�A��5r��u�&c���x��E��x�q�t�C�y]�D��z�Ѕ���iz�Nt�'-k�5]`@W} F͇`��6�],-�G�;���g��խ�3[��g�)"	�%�ݞ��-���VkE��33[��v�n�U��
K��|����2���刔�T7k�[�Va����6�����*t�h<�$�Ns��{}�vx�P��,��pM7�7I"�Ȝ�@�o3�i�4���MD��wEUܕ1Q5Uq�&�3@m<�4����p}�TJ<kS!�I9àZ�F �ot���O�w9��I�(�!�3�m�{�-���v�ݼ�۩�7RbȜǆB��'N����&��|s[	Y�pd"��']�lr6�x�hNw�m���v�n�g ۶��{Z��4�ā��s��ǎ������G8=�Ҡ���v�8�V�O��p_$�àmO# M7�i�`	���<� ��d�舅��v���y�n�S�m����n7pn�E��9ހ�yi�4���M��cq�q����s�t,�غ瞐��^-��֬<����O
kAc��xy��rѓ�Z��4�i�`	����O# 7�Y�D���dRNp�v�8���	���&�3@�R:2쉻���'���z�x���ң/a(J$�irYK$���9���lhO�F �!:���J�
	�������{i�`�=�9T��v1H�@��s8��{�n�g �����y�sۭ�$�E&D!'�
p���`�\N����0Mɧn6�ܥ��w�	s���}E�Ns:ݼ���y�Oc@�l��.����.�j�0|��	���/4�4����(7q�9"�Ȝ�@۷���{} �y>Ot�%�����*b���� ^i�h	���s��K~){#�0�W���ޜ��6���@)�ȉ'3�{v�8��݁�7J�Ϟ;V��n����vr�#�I-uNW^����'%�9\<��d��,��	kv���P��w��|�tݡSk�~O��M�`�=��y�ͭ�F�0Nw�~�y�]�΁������ށ�u�C��ŉaUW�Oc@�F}�ϓ�ɼ�}�+q�'��<���tn�g ���@�o# ^i�h��+"諿��fn�j�0|��M�`�=��xr���F�6`��4R�e���ޞ���ߟ�߸�V�Y& 
�y��5�1��2u�z^9#j�l�'������ȽN#��-�9,�Qk�:XN`��:ȕȜb��+p 3֑���[\��v[s���ܬ��Wlq�@ݴ2�u`:��|���IN�;��n:i��+��t]e�/1����`"�7�"�F�\v�6ۃ���a��G���.����xg]��a�^C��ݭ�J[�Ωü���8g,�V�xkV�����=�:�O]d�����[qh�c�;�����՝�����,��P?��������tn�g �����xY�#�Ʊ�ۊ�Ϟ;W�
d�����۰>��TDF|�\�D� S!�Ng@���p�ot&�0ܞƀ�H�˲&�����J������<���r{���������� x����Ҡ�"�����*���������9�(
�HǑ����FH���4���y����#�N��S�y�4��EUUƁܞF˖F�K0\�(̒qO<��x�1��mX�ү�!G&YD�S{���U�w�*�����g�|��̌r}IF�s8�7�i�`�=�4�0|0�����,��v�8���:ݼ�z���xY�#�Ʊ�m����j��P�c�J�y���J�=�V���MX@�<��$L�%$��]�ˮ�8�{i0g�[k���j�z�����EIwyi�`������>�{�ި��9hܙ�/�[ހ�:T�2�o*�	D!�c��C���ݼ�m�:�������~���'X��I#0&Ia�2���,#(�i���X��@�Q�)�� IHH��{����!a�$̂F	Yd"x�0HмՎӊh<	��1I%�"He!��b$��$���*e%#$�h �������r�����b	��@��( ��IRACX�T�R��$���Z-�d������Ph�D�XD�-d5M4�~z"s/���J��C�e�hQ�a�2c�����2@�Ɛ��K���/��o�.���|Ae�L��Ap�UL����E=���� ���*��U?[�~p�_~���ʽ�]&x��xt%�<�:�?I�=�,״��=�O# Ԥ�ʺ&������ytX�@	BI?f:��J�e�:��o�pII�(��J7$UJ^\L��v��u�w87m�sm�y�kC����>�$�I��n�ށn�g ۷����p�h7q��G$�9���@c�L��J�Ǎ��
F���������$ۙ�/���s�[���=}��ݼ���y�D� ��<]�iX�@{3��Ҡ��4�DM_���t���g$18b�$!�3�{s��(~n�x۵`<�J���fߜ���g^�Y�S�iZ�r��:��aXRm���,�Q��;v7R旌񳉫��y��ƀ�y$���Li;�X�6$��ݶ�:}�g��*٘��~n�j��Q2krKӗD��T]E�w��~o�F�'�����m�t�ʎdc����I73�{3��Ҡ/v�6""b"������o�d��&D�z����mڰc�@{3��Dz3v�ނmt� V#ur�l����-:YJW8�8�U�o�גպ�9�b���szfvˍB�A@Zn��;OY�nr��#;נU)�.�E۞��Of�S4d-f�ob�&�;(^��</�ul�k��vjH�I=�unuG
n3��عK���'�b�;<5˻+6PX�Uюd$e�jme�[0���ꍅN-۸�ۃ��T��_��X�9�w��1�;�%gatD����c\K%u��`;xn��Li$�6�O��<��I������:I�`�{�>o# S�P����$��Y7W�h'�� �ot��`m�΁����'<lܙ�1���~n��!D)���j����~kb��CF����8�nƀ�yG�m��9S"�i�E��TL�\`	��4���m���8}Eq<U�dl��"0M�	���\���ɻ[�b���۱��;Zi�>ևDb��6�ʋ�����O# M���l���:�eG21��pJ$���6�|�����	� ���� ��{���g �L�v�H�p*n��@|�$�ƀ�y����1�}���i9�ݽ΀�y����� �}P��D��H]eM��F��y�jm���0n��t/��AF9�� 0m�F��T�&ќ]��`��h�4W��g_�ܿ}�ї4X�#C`��΁��w�_YN�ݽ΁wo3�w�S-lR7�hs��y$�ƀ�y�����ʙ�'c �'�73�{wos�]����)H��m݀��*��N5��+*.�*�c@i<�Sot��`��3�o��G21��q%M�����"!�yw<�w,�����\��vN�h�vzuŨ�#Ag^e�,�/��KgQ�.(�ks�euM6�M����0�y�Y���	;��c!&<K"M����3�o����m�@�����*�mL���$��4���5��@|�F��# �j5��bp���8m����g*��{Õ�����~�Pyx����xͭ�F� М�@�����!6�U��*��v��c��~�Ş��wi�L!��V^��X�zxzю,���[���\�O3�H��0������F ��F �ot��`u
�q��<���s�]����{�>o# I,�#�ȅ&E�Ud]'y3�uP���~n���mҠc�p��d������v�8fe*3�J�R���߬����oc�7qq35Uq�$�F|�,�$��v�8ٝ�>����Px��  -�6�ے��U�ے��2�d�2ɴ�[a�y,�vca뱣v6��	�*�t��j��U^i���*�m�v�Y7n��H�+�n#�+k\�x��dm�"N�lb�a��d�v�c:2^��"6�,��-k�O8Ķ��8n`�i�k��nB�H9U���[�3�ŗ�ؑu%F�jN`�����$�;]`�.�r��������{�����wقRC�&ئ���9՝���C=�uC���5�>�����;]�����ر�)�~��c�{J���w`7��∅r�iP�Ec|X�`�������@�o3�4�F �,����@�n������#����@<n��%-�@]����jb�9&��M��k��呀.I��y�$�tMY]E��W��6�F D}�y�6�3�]���7����9�H�B�ƞU���j��\\��7h���3E���bA��%ϊs��21��dDi73�o�oz�y��t�Qr�@nja���p�y=������������Cd0�DEBQޏҠ3��T{1݁����}	&LKm��m�p�o3�����v��[���*�˪��Y�U��6�F �'�i�`7��{��[O���!�3�o�oz�y������p�
�N��"s��h
�-p���8��q7"���Af|;���,M>��b��q�H�!�Ntv�0���呀.I�Ҝ�%;�����*	���o# K�F �'��y���[G1� ���tv��_{����W�*+hɐ�u�����mmҠ7��T{ �K�9�Ӽ.K����r_�@m<��l��n�� ������$i�a ��@�nF Ӷ`	r��M.&�+�ێC�Z��5֮��s��=\p��Nt�K��J�ւ���{-����5�'"�`�� K�F �ot�����+�Y$�\���+���x�V�%2n������F �Z0yH�������*��9ު�n��ңR�/Y@7��#���ӽ�9"8�݆�D�	n��@<}e��A֒I�	Db_g?����@��4��nH|����V�.Yi��O# Q�U;&[��1����G�玂�\;8��݌�̀�'k]���K�[q��mHWm�������o*�n��Ҥ�${;��[��21��pJs8�oz�y�=���R�Q&榎oN�{<�z"��tߟ�rY\�0�{�nٍ���I2bX�ng>Ͼ��n�8g�� �7v�)z�� 4�t'Db�҂���g@۷��%�o��]��^��~ܫ����0?�UU�� ���������b� �y�sq� E�P@����q��
��֏���X����������W����o�������ؿ��}����������P�U_�����=?���?�?�*������DUB� |/���'����������UU�o����%�/���t�˨����~���_���K���U��?s��]T�F$T�		D�I@�Q  �	D� �H$%$TE$ �q�(�P PҢP�B!J4B R҅0���(HH�2H$�(������0��H$ 0�"H��2C �	���H2 ���0��*�# @��2(��
�!$# ���! ���,�0�2��1� A�(�J20,�! �2�)�Ȥ�($�
� � � (J0� ��,"! �
B0�����H2�#B4#�%"4���� ��
� �
)(�(J0� H ��*�(� �� ���(��� (�2� J�����B
�J2
��
 ��"$#(B$�	�2�	B4 4 A( ��H0�#�£(*���� ���@�0��*@�� @�
I���$�JJ��H�, @��(��(��
J J(
�9�f��������@EUX�?��{���=������?���?�������a������#��������k�����O�����;�����UW� ����8G���QUW�����ͨ���[+�����s��ʟ��NR#��G��o��BP�"!Z���?�� ������ᑿ����r?����F �����Ԃ*���������z~��?���g��/�j��6����y��������g��D���������{� ����s��\?�� ������+�?d�W������e5����� �s2}pg�    *    
   �    @�  � ��P   @    � EIT��(�DT   ���� �@   S   F  UU QP�(i�S������Z��u�s���{�@��']5�}=Ž+qeWܐΔ���8�|  Σ�:}���� ���{pq��;Q�  -�m�Ӗ���Ҭ^�[� > P*T 
)@� >�b�E9�t�����)N6R��� t���AK,�J;�)E.X)��� ��(M�,�� ��QLM)@���JR�h��w2��M�Ҕ�p��R��4��٦��M4i���� ��QA@ � 6  ���
�����G�.�����G���ruK:���&��Z������R�� W}���w|[Է� =��m�Wcs��{�/�A�-�{g�_<��99�Mo �|
PR@ "� �j�����o)��[׍�9U�P��K��S=��i����u/��r�-���ͫ���ݚ�]�^��GyK�Zr�����nm֗� Z������z�{<��N�-˻m����)@� 
�6 ϊ���V�ϋ��kٜ��� �����nn���ɯMŮ�����/���g�|�x�y��{<}�}� 7�'�k��ק�'�on��鳼 }�����������/v�u;9q�� �JT @����ʤ�@ 4 ���R�dT4  ��T�EPd21����)��R�  �!JSH���㿏���?��s����3��>��k�PU~��AWB�(�qW��T_�"���QU=��bHB/U �b�E?��t� ?�1
��l�A�)����8c淚޵��@����
��@��Q�G@D!�!���āB5�aH�"A�<#pYpc\A�4���59��Ƥ��y�������)�0�"�h!��y7�!�b�9/���Ku�����A�D���+++
@��XJ��$�����#�R8tl�)�IsFУ�Bxxri�dM0��F�p��n54�8��N�I��	$�)��%4�<tnG�/9ɥ�"� �C��i��Ƙ`�8'%H��p�@�X� Ĉ@E�A�%HB�^���A
!��{T��I��(���ֳg<<6�! i6*��� P�[�������HB+�)@� b��CDݷ{��{�$)���y��e1�.fg	o�]@"C�#O0��q�qЋ��
�y�y��2��<�p�x� D��)��@�� qӠ��8IB8�Hj��,8j���4�*J\�Ӳ�xŉ���R!qZvi!L5���bA"�0�H��y���$k�������煙�$�	C��`�X!T���ȭp.�=�<��0J�a��ǌ㢛�8�Hi �+�%0� F$aq�F: B�s�_���b��8#7�"�4B�ONo��3��jf��<v|�9��͜٭;���N���
O���Pq�s��|�z,v��W7�tB}�{c � E(��!,�:'d�@J`qU�����	r��Z°�I�z<>��$�l�H@�42�2F"�D��w� HR0���4���h�\t���]Sa��8n����ÒMf�T���o��o�\4�6f́y�h!Y�5
ᤅT�bVV,X�b@�E`H���D�{�m8�I$�$�d�אHjxK0�m0��.�у�i��BHQ4臜w�� ����`�l�������EsF1f��_8<P��w�� �YM���L~PXz�i���!ϧ��=x���&:~t�$
,@�E�E+��
!�0	l$Mo\ܻٛ�{%��Y�xa4#P�H\HS\aLHF��&|�aM����ތ6q#	�<�.h�Ii���9��u�z��U!Z��<��\���a�05��IpѶ�OY������l���*K�}���(�����H���.����3��㽞����ZB!��c��p6�O��!L_`W\�ܸH����� �_WD Eb�
�F��F�8�O~��xhhԟ\)��~M�DCK�~xH�p4�) �-0���)O���0�<|U��1*A"C	��H(�B	S��p���`���*2��	a1މK�	�٥ѣV	&�*�$Aas���q��a���x������	L��14�;�N�2X�7��[��AHcR�h�ɪ��j�!#���41BD(c.a����L+����#�k�Cf�@�-+���^�P]��!tv���:f�&��C���������s&��/0��eѾaJ��kd�y�0�RJR�8F�V4�1�.���HHGǒ�,i|y$.�a��@��0���2)��D�MxW� �)CJ��5B�Mb�)�R���g�L������N/�cX��D�F$ �!`4�*AH�h�*	�h���o	1!4pM�
Ƙ�6���A�x0(�:M�c�܌�l�5�g"m S�p6������!�6p����"L4l��@7$K����k��@6�p#c4�C[��u��F@���r	P��𰤎 D�@�
1V��� 8��Lt])�ۯ7w�}��9�p��_- bq�-M�F�|8DXڦ��"�sG7w�p���D�j`��|<������B!\4����x�q�V%�C�y�}B�@�8��JD�D<�a�=M`�$`!��w+�WA!$HĄ@�d
B����m���d�Cxy�����]h	sU�1`�@�Cc�2�5_=ôA)�n�`�P<�/��`S����S�#L(n�%4�j����8�JW�t޹�y�ȁƲ�6�v������S��!3BA0 �B����&j�aG5	$��! �X�BH�$ D�@�
� @#a�<!�HɁ$���Wf��r,���"�$���(j�F��8BfjSfH<�D�S)���$2�	���
�ȑ�k7iԆ�.H$$���6L.�.��H°�L&5ke!%�@�@]���8o���P���|�=ߜ�w^y��No1�Ĉ4�8H�
�bb_E"�X�x�ݱZ>/4F@�)!"F�2!08�`@�m������sXh��ԗt����# 1Fc��`�H@1�7���a]��<L!S�T�@�H� A�F�������L]�p`P�ѳ�����$� ���F��y�&�c�<�L4l�H0�pM���)���M9��s��7�L�����6m��x�k��s�`p�ɭ�ژ<<�
�Z���� �#sR;��vA ���0�ā"�¾�]ģ�ВD�CS���/�!��`����(x!@�6xF^��R$cY�@��ԉ`l���
f�I���l� rӳ�j�XI%`�`N;�!f, F��I!%i�Jf���ܚ�G��;Bd�$#V)$���	ŋ$H�H�ъt)��$��v��1�������z�)"�U�6�Q�O��i�H @=s���,�w� zy �J&�J"�HI%*V�C� VI��M��,��+�bH�%��<�	�$�s�k{O�о1��F�)u���f^kܸ��x�ǀH�(FC��L��v�8�'�q��Gk�%�S���:@H4@,���&�(��"YK-�%�sp�l��:7Cc���9)�+�#HGNߓ!�"�cP��F^I�L.�q����%�&&�(hӦ6BY��`a��!bd
8�FK���&$H1���9�tܔ<6sY�^	���c�A����B�����S�����BBP��v�	$)�<��7��<�tq�|&�h_�6E��� �<�E�h��1�4Xe��9��u�kZ  ���             �       -�                                  � $                           ������ �l$n�H:�		m������` �"��#m���^���` �۪����Fj��h6�kvP6[�ж��  �i   ���n�-�iW��6�� Hg�V�M�� 1oT���o�5u�2�-��� ���2՜l��5^�ޠ K.� ۱��� 	 H �j�7In=!���6�v�m� �n�mm&9m   �[I&�Z�[׆٫I��6ֲJ!:m��*���s[9Jݪ�(�$�a��6�&- ��p�`!�d������`  �n-��궪�d;d)T8��F�M��nݤ�pl�  d�Öq�� �s��|�����v��m�-���[Co��| �_i��N^�� �[s#�	�Ԁ�!� 5Mw� T����J\U@UWQ��U]����-���H��K�z��8i�iu�Pit�l�@t��d����n��� mSf�$ ��I��MKhN�ܴ�)�H-�f�!�m�At[*�M�l$ ۶p�7ll-�۶���$�܃��OY'Qm��H�I���^�&�n�
��_e��LV�*��V�AO0�۪�ŵ�&�p���q�rݴe�� ��ʇK�7l�N�*�v]�:)�� �kh�snͰָ[@ h� m� :�2L��@6� R�� �� ����}� m�@9&�P  �t�  n�kI�NtA�ŵ"@$���i��  \���À�-�� pH8[e�m'`8�+�< [m�	 $Ku�,$�ۅ � p�˷`�ط�0q%�Z�-�B� �6�[N�c�� �6��m��G$�l�P�& �`�[���@$m �v�m�6��m�u��6ۭ���N� �6ؐ n� ]6�ԍ��L��UUuRˬP!<�pH �:Ge�m�8o9l�+m���`�!	.�۱ �J	6ؐ*]�` $[[ml�e�:l@���n�OL� H	[G��`m[f�[l�6ۀ��t�[@����  t�$��
^�5moUJ�**�   $ 8 6� ��� 	OK5ŷ����H   $Htݰ[\��0�i��lhm�8       FۯK`	 �6�9�m&�  �f� ��` 8�'l�k:̀ -�  i�l4u�h8  ��     �6�    �b�n8H9w��>׶�ж� [@���%�6�        h  ���~�6� 8HH��� 	 � �H�\� 	$�A�mt�Ke�    �AcM�`  �$     �2E`[B@ �� ��ޚ�o��   ��d�n�[ yar��P�v�K$����lm� �n� ��� [Kh$m�I  �OM�l�-��P ,�:[r/B���N \�3����  ��@ n�����    [m�˦ͫ`E�$  hp 6� m�n�4�i-.��Nfj�v8����H��yYX$��'U��� �E5�-cm.��N��V�T���mR�'I,��6��;m-� ~O��m��vҮa�ks6���������h���h�m;[s$�h �5v��jۜH� � vٺ�`I�v� 8/[֛v��r@r�`6[J	�Gk��C��ݬ��  ���� �Ӵ���4NSS�Mt��)m�   d�#�q �sc��I�ӟ>�N��|,k{n�`��7+UO,�fې��n��^gF��\*2aـ�m
D��HUR�Un��Jؐ��V���L�ڃaUQ����9�[pX��Q��L�h[@ .���mY� mR��v����gv!,�ԫJ�T�v�l��
m��% �kZY@��"��V�[T�5R [`�I�m�
Ak��-US�0dMcC�^U�L�i`���t�kn� 6�H���vݰ ڶ 9m 6�7�����D�*��M�oNn��l���,�����i6���*wB�<|&�v�\sKQh� $�   �V�[n�m�� �   ��n  f�$`ړ\ m�  !�k=�� � �m��m�� �  �Uoju¬RV���U�6� [v�6��m�2���ěI�	 vհHJp���m�&���@  l� VӠ p  ��@Hm�mm��BC���8mt�	 �N�l � �l��,��5P �-���eP�m��6� H�mmn $���$-�6݁� l	#�h  86�6�.처^;k{� �\M��lfd�8Z�)!Ր��jOT��v�Yy׭��uէ,�&9���:9;^9U��)�I��%�f�P�mz��`݂��U��A���wD�UUS���x�Ǝ�>UHN�m/-vh Xa��� UU��UT���!��mm�R˵��E�[@nղ����j��o�}���9#��Z���  [@ ݶ-��p  m�  �:�$�t �M��WhhlsZ��4��l�n8� h6�    {m�`��Hlp �ii�M�ii7H�&�6ܛPv�u�  8$'m�[@�`��  � H ��@          ���,�m�mm�p�� ��[~�ci6��D����[Am�mmŴ; �v�nle�3i  a�[����J�]�m�H�E�h( p  � $ � �     mZγ#m�8m�:�C�m@   ۶�    �mĂI6�n��QƳ\  8       �k����si6���*�U[ T����Uv��I-� H 6�Yg$� @�g��z�    m� 	 ��-��U�&՝���`��l�	�}���ր5��9m��� ���ݰ M�f��Ԇ� mm�r�   ;m�l  � �0    �n6��m�-�@m�#�+�*����T�F�        ��B�:�j� ��m&Ä���H�$���� -� �n�v�Y%  :M,���l��� ��M���ko`  �m��h����u�ں��A��m���nlְ�  H[@ �|����UaWev�UJ���*�˳��vYH���j�̐�((
������5\9evMW*�\[�I�t�  �@�@ �L�M6k��� $ �H6�e�J�q�C�jP��n�P+k��6�E�U��m�����n}(�A��7b�j�C֦8(1f���j�geMM];�Լ��A��vmN�-˶�C�k�������x�,��*�ACU*c��j�ٶۀ���H������Ӣ��6݀��0��6�� ���� �EkŻa��\��� �X` #!�ͪU���eZ�IiK#Q�U��XKt�[R �  p*λM� m�Jͭ̀p�&�   	�!m  �$
]���6�]��U@Tm�:�z��  �   m���"�m  �Ep	  ,4�m��[p� E�m��ܴ[Am�m� �e���8�P  Hh մ ��  m���!��l۰H Zv�h  ݵ�  	����@  
P�m� �L`   f��	1Ā %�����    -����m� �$��6ہlp$�[s��m�m�   �8-�$��  �m� 	ZIm�l��B���[dX`m��  �j�ζ�Cm��m�6� ����H��  m�]�6���� ���	*i6y�m�������m�+i6�m��k�[��g�@��=�e��F�  !�SI-��l2v�������	VBi^iV��Vy_��� [A�8�t��lp ���w���{����w��ya 	d���v�?�W�/@�v���Aڬ ����E9�!��@�"hҢ�OOpQ|��(o�NFM�L#�

�t(�x��DChb��J�o�%A4�#ϑ@�@N �� ���W�_�� {�=T�TJ?#Tg�z(<M)��y
�FԠ�[@�8���@ iU<G��@� 	"$�ABE��H1`��U�EH*��| &T�/��Q0給�PB�z��:=C���T(�����O��3c��6�	F  �"��R,@���A8z(���=�� "x���*�}@��&ͯ� |��������b��SA�Ep�t
�A0>Et�@P�t�/�
�qWj<�� �/�$AVͿѶ� @       �     -�%\֌���4��n�`ʭUs7=�v�Vv{[�$�\�*�{Dr�sl�6Χ��N�Ɔ̭�h�V5�3��7cKAJm���c����=��ӶyN�b}����m�ۋY����{;AݔA8�ǲ��`��[��z���dWO��K�Z�U�]��HR�U2m7C.i��
��ont2��퐀r�muJ�[*�e����9݋ �4�ŭ���[C�ܢ���6mM���l��1���&����R��Ke"i��!���e��Yez���8y�
����$ڶu��J�J�3-UT[*�v�FM��$Ak]�Hu��lM+y���\��\�B㇣�IX�Z�\��u\	�f�� ����=UÂ�5��*���7�x��7%�ɨ�������pn�㊧��:+��UkZ�`\����8e��cԉͭN��^Ȯñank��$d�����+���%�����@j�/m������;e��N1�@��D����K+��Ԝkp���n���)WҪ�7�j�T᱀����e@S�S��U^�ۉ�v�qA���C�ݻm�i6ۄ	��%���Ma�One�
���ҳΟ\\h�vmR���s��]d{��ct�  �o6��7mnRc&���&@�iV�`	bI4��F��m�n���-�:����n�NTȵc R�mf���mHmJ�B���Y��Z�Nv�4��;�M� ���.�p6��)ʎ84��p��a a	L�T�S�n۳�-���P�������e^�s�^��t1&���<P�1��s[6�@�ܪ�A7�ohS���5[5m@�v�t 
��-jvV5D"@X�P�a���mpW<����P�[v��˷$t[��*��ջI2�3ʬ�2/m������n	X! �=b�0ݪ�m�ֳ5�SZ�kYl�J���W�����Qq �K��R ��{�˿� 6��gT�M��O^\�s�,�;E�C
�]��Nɂ5����k;�`9�b.�ٴT�]�FZ�1O��p����n��\�t����gL����x����n�ɵq��sm��H[�G7Hi',zYND꽺����U&�g��I��N� t�h�C��q	؞ϳ�.4�m�W^�M��yW\u���$�lv���{�V��섺� b&�i��,4C0�*n9�ܯ>q�.7w/��06=���wg�";<��'����d�u��O:;<��D�j�-aB	�ܘ�S�z��o��(
T��2i�OV�$�{1�'�=��AH��Y2FӋ@�gJh+k�>]k�;�U�w�����x�0Dk/4@z䘀��1 �9h�n��ו�6�I)2F��=�ֽ��Z�:S@�[^�����1�n)�d�qL�=/gq��&�qn���2��w7N�!Ղs1�#��D�0��)����ݝ)�|��@�u�@�wx��ӭe�u���y���($�!R�D�*x��ۿ��
���Ϫ��U#swu{��$��Ɉ��@s��@{��Ց8�	2!�H��Z���h��M�mzs��q7&%�7�������Δ�>Vנ|�נ}���LM<�4A�D�,9�%��`��-���@�v]��-n�X:�Iv�6n�E$ɒ6�Z�:S@�[^���^�����T�F4'��F�8h�& =nL@7�Z�=�ߪ�=r8ۘ,�i8��<�k�;�U�Ы	
.��E	b�^z{��������H���a1�R=�r����& =nL@t�W�19�m���@�gJh+k�>^�vI���Y'j�P���t(�"����y8���ط)[;%b��V����ֳ�� ��!�"s#��y~���.��Ϫ�=�Қs��ɉĠI�jG�|�נw>�@�gJh+k�;�u�#q�G0�Ǡw>�@�O`���1�rbҜ1V��{ �L����=�Қ����Z�:
�4
�Q*���^�rw?j�/~R��OL��|���rb�r���Ht�&nޗ���[�Y��=����C�y�ܮ�݈�ᇀ�u2�$Mc�6t�I�������1�'�~�d��{,h�������d����H���a1�R=��Z�:�h+k�>]k�=]�G,Bs ۼ�ʹ:qR�$��Ɉ��@�� �'2&��Nf���ֽ��Z�:�hٍՓ�H���Ԏ�<^�vIڪ�&j�'�3l\�����6� �+ �H�w绻�w������@��������8��dӷ^k%���1��u0.�F��r\��������rv���7<�۩���{\9wj�8���KE�P��κ�]�I^P����s!����!W����Ʈɶ�c���%u�h�	q���d;j87�R��YP�Y���=Cwe�]��-�'3Xo[���Aͩo)�vy��|��R���=j@����z9��qenE�^�o$N^G=�@��g��u�{q�.6�f��������2~�:qR�I�[���v!R)!HA#i�d��{,_�UT������<���@�v��T�F<I�$��Rf��mz����j�;���z��9�,�i8��>Vנ7�Z�qR�I��,�ͳ&9�Ǌ8��j�;��4+k�>Vנ~����b��ؠ����dm�u���X1]����#�x���,���3ňNdi�"�r�Ɓ�mz�����h��$1Ĥ"hH�!��,�wʪ�:�
� byn�>��Zvt��m��Y18��b��z�I�����@z㘀o(vL����'������z_�@�,�h+��+k�=s����G1,�Fӊ�>���d�]{��I���d�y�Z,�:� cXL&���Dxun����g=�v�k�ΧA��͜�nǍ�����s�y����'�z��ֽ���ݝ)�^�G��$NH��Z���bE�?\��|�W�֢G�Ls	�����=�ҚO�E>S�PM��u��rO/�}��s��Tq��72$�iHh��M�z��ֽ��� �EIq)�2�D�9�[���Ξ� �������u�^���å��k����Fzܤp�B��헉�V\�љ�f�y����1 ������ ;�`��NF(�8��Jo��`ɦ�=[��ř��
�A#��႑G1,�#m�@�,�h+��.����;�]dc�<b���''@�s]�z�u�'���d� +3�������>��{����Y 8�����Ɉ�`��͂�����~�vHNł���R9���Ր�l)��=��g��2�=�ݶp�c�cSƝq��w���`��͂�������*8�#�m��4w���z�ֽ�Қz���Nf�YvY� =}& =}& ;��͒���Ց4�7�z�ִs� 9�`������9[�y���(���{�4w��ֽ$�����}$�������   ety�:�0�3�3��/%����S6�����&]��u�)f�v]sK&����>��u:��-�n#�:���8�I,���q̒-�y��ܶ��C����.w)��HI���vy�x��d�'�h	�m�\�à��C����p�WȚ�x۵��:ٻ9-�θ-��p��+��\Tt�GU�l�4j,�%���v��zч���.�����q����ɶ"����Nٛ_D�eL�t�J��8�J�9�c�n��O�|�k�>^�����W\M<�(�!�@�������c���͂ �swr9#L��I�����@�Ϫ��fg�%֓�yu���j$qDd��˽�@{��@sf���1��1��$x#�m�Z��M��_��<���}��h��$q&)�=�V�&��}���&�s��+�q������IoH`I�$1Ĥ"i$�!�|���/Z�����Ħ�k�e"i��$vI��c���)�οb�ZJh/uz���#I�5��ff�ݎZ�6_9�_I��i����bX�FӋ@�q)�|���/Z�����%ު��i��1BQ���K����Z (��}�Iy���$�|=xyĒ�*��f��Dc@=��+��.-��m�ۭO]�>���Ųn.-۲��
�U��fA[?BIy�ߟ�$���ޤ��gm>�$��Q�I%�j$qE'21�R?�I/7ջ�B�if�<�Iyd��$��8�J��I��F�mGԒ]�_��W��}~Tx(E���b��1
���"f��f���6Iڃ�]o��6Gှ���� �F�,�Q���H�+j�Id�D���h-�Nk�;$	��"B@� ��I �	R,�%Q��(�$��A@�"�� @�"Ą�# �RBH2�6,A�u�;ԪE� 0�$F�d��TFQ���*�����$Ba$�!A��C �p�!�v A�lxF0�*��� J�B���>࠯��pQ��"t�T<@�@t��*�0�T��8i=P(�4v��s>�����m�g���3Y��q)M$QNq%ڧ痥�I.��{U޴���n���a���K�{�w�L�ԓf�� >����������I/x�89Ē����$�©�է���5%�+q=�#���Ѡ�]�;v볓˄\��X��j��b�������$�q������G�$�}k��뒛(H�<���z�K��ps�B�Pm�,�]������$�[�7��������0M�D�ϾI.V~������K��oRIw~ϾI#���Fǒ�&�������Kٞ���m��=���m�5�)�A]���֤�_^C�BNdcĤ|�^O�z�K������%�ҵ�$�}�u$��O�r:�M%�Г;��۳������!"�ۉ�{����7Ҫ(�z�J�������ZԒ_>����`�'����Y��q)"M��Re��Iyd��-(6��u�%��[� q��a���]��A�=m'q�c����]y��͠�^o5�I%ʪ�����Ir����6Ҷadiȓ������$��%���$�/���m���$������Iu�[(H�<���v���a���K�&������u�%�Z��]� ��[�Bd�I#o�,��tZ铦��Mg�OF�'���պ��p����n.��+�,vUh�Z�<U��G���b'��l����y6���2l@Wcɫg�j��\��X��틆���v9���y��OS��x�nɶ��Wl;R��q4gS���2�i�.��1�����G2,��4�\WP�=NW���QÅ�C+��Q.k�B m�Ր�j������|�~��t8Y�9-�q�-k�z�x��ɸ�����6�kt/]y�N��!�(tn!�w������?��K�7^��%�Z���9��I͸���fA[??�P�������kZ8�K0��s�.�痥�I%����(��H6<JG�߳k���ԒV��]�Iyd��%� o�7_8�K^�G�171��JF����m+K���I.V~������KϥkRI.�
Hc�Im!
C�K˥������KϥkRIw���2�U`�+�I�E���rqM�^'��5�e��61s�,�>.6��:\�H23:l՟������} u�cV�K�>�?�(Uw�%�K��Y�o��`H�K?_@o���7����A�bP*+��~�}�<�Iud��$�f>s@� Il;n((H�<���Z�K�]�}�Iyt�Ԓ_;k����ZԐ�rU?��&҂X�bp����ZԒ_;k����G�$��m>�$����4ђQ�։%󶿾I/>��I%��Z�����s� ������.,��.)������/(s��>x�n�=3�=�=�Bb����أH�ԃc�|�^}+Z�K�����%�ҏRIyޯ�IWة#����m%#Z�K�uo�K˥���_�$��J֤�^�
Hc�Im$���%���I.��>q :�$�<|Aj ��7��컶������r����������V~���r��k����ZԒ]ӫ|�^](�$�ߗo�ސ`H�C?_@o��� ����߼�\��=I%�z��I.v;���v�Z��srom��\�ny��΍��,� Zt�걝LX�1�zUd��K�uo�K˥���_�$��J֤���T�Ƙ�H'�M�����G�fcm/;���Iy��jI.�տ�I#ֽQEh�0j!��$��W��%�ҵ�$��V��$��Q�I%�R�(��H6У��KϥkRIwN���Iuzav�� T�>��|�I-z��nUpR| ??/���� }����x_Iu��%��ZI-6�:N�&�l��;�J��\��w5���V.����ys��vjw,k��{Z�05� �~��K����$��W��%�ҵ�$��V��$�y^:�N4㌎H=I%�z��I/>��I%�:���%�ҏRI}��N$�mG0����%�ҵ�$��V��?�m�t�Ԓ^w����
�P�ı<���Z�K�uo�K˥���_�$��J֤���T�Ƙ���țN7��%�ҏRIyޯ�KϥkRIwN���IyUw$	$�H��I?�1]��DL��y��,.6;6�+��:p�]g`�[t�����%��;v���.-��� �ۑ�<0��9�j\U�e!�Eu�k�y��:��ٺ��\6Sa�]�m�4s�`��y�tokjB@�vˋrK�Q���.���!�ݪ���i�\�7[�\t�/`��m;뜭�C�x�ń5cu�۱��E��/<�ؿ�����/_���т�m]:�e�8Põ'���[v�X�A�r\Ŵrk�ұ��s�p~I%_����%�ҵ�$���o�B�*��bK�&�i$�3uQC�HQ���%�ҵ�$��V��$��Q�I/;���I*�$x#�&���I%�:���%�ҏRIyޯ�KϥkRI/[�$?�bm$����Iyt�Ԓ^w�����Z�/b����U�lN	���<�W�z��@6�e�=�`����+7�6���m�)D=t�۷�ӓ�� N@���i��,f7��X9��ȇJLQ8������-�{\s0w4���q ى��O��_k���� Rd��hu������$^���5�`�DdM��>�JhW��>^��޵�(�?�0�Cn\s�s��h?U}�W�_8����H�5�dQ�=��@��Z�>�JhW��>�qD\PpX��r�t4qּQ�\u�5��9�f�ָ�<�ϋ��)���{5��I%�H6���{�i�{\s�sID7O�L�M�����t����H���z�_�@��Z�*�m'⌎HhO/����r��ٹ�S� *�f{�}�@��)�}��L�q����@��m��@{����L� �#�cdM���ҵ�}��<�W�|���Y�u� �LS�G[�ۮt���vAg�ݼ�`-.����<y�k
e9�1bx�2&ۍh{�4+��/uzwJց�Z�Ex����D\sU���1 ���@{�� }��EkȦ,QǠ|����+Z��M��zob���9��a����̴��q�ATUz���7����4�JF����ɓ�s��h�ɤ@p�cn�k������m�S��N�����8��m���Z^e'M���9�_9��̿�_}��9�� =�h�&b.&��D�O}��U
H���h�?���\|XABG�țn=��k@��)����K����]=��S�i��16�k@�=��9�_9�?}_W�$_���~z�j,O���Cn������$�ޘՒy�L6I�@��UH"��#r���Dhı� $U��H�=+n
kj @�+�b�mIjI#,c)-�,��!�4�R�fr @D"��.BBC¦#ZT�C0��%�HD>C1�� ��!��a�HE�͂ŉ��FH:0c���1Hb&��H1P��c�j�& Z�$$A*���(,4<H D�B!0�B,RA# '3Sh0�#���`D"�q	 ��L@�	�4�p`d�B$�	 x�]h���0B�B)�׿6�kX  p �`      ���    �PtE^^6��iΦ@q�6�55Y����dv�02��@�Pn����VZ%�Iӻ\�l���{Q����/<H��=\n̼4�t9c�AZ.��7s�X��b��G)�i�;Z�:�X���Eݠۧ�W� cdu����)̮Y��$��d{�K��孪�"�l�֏Hv�M�Śjԅyny��Y���s�{r�TF霬�T��e��Y6Cm�^ݵ��L��`��&���m�c �a#�MUm*1J��l��T��m�Si6 J�[�n��U4K��`*�.Qj�Ij�ݷ%�l�i�l ��%�t,T��u��q�����E��̧S	e�r2U�[�&�VyV�)�#tR�eYV��V��\1��pt����]���K���vw2��\��r��ɛ5Hc]�ٕ�G2Q���ΰ��"m��;��4q�bN�{cN�,� �j�3���VuѹK�,�/i��E���� bvi2!'[FlW��� 7K�֬�����1q8����im�9��]J����sulٔ�{b�v���Ve@u�	�P���f{��;��	ۓ�$�4:Ki6/4���ErI�.�ڃ�^v�UR�*q����_S3uӤU��\�j��m��t[L	��mT VFĝ��K�0m�:6�R��T�UU�����%�ꪡ�6(�r�9$�Y��[��ɔ�5C�Hx����V�*�G����vf�A�UjP�/=�5UU�aI�%8Z44��R���݄k|���Vҡ�e���IW�%��U"7.�.�:�b�:Ĵ�/-�T���^!�U��j-��(�j��%�C�f�q�<�fțK�ۨ�.�T�avyn��Dm�<뫥��6C:#��z�`�e�f�ʮՓZmv�FX=�nx)U�kl[��W�J�n�@/D�뛲�g�r����tR���ԯ.���e�lѠ��"!�S��� �lPE� zl�{�w�����_��H �`7Me�ۋ�'�JO$zͲ3����-�q8�����]m�g����C�>|.ͷ]�P�d5��]r!��F�#�T�bY�,N��Cų=���m�D��k�8��6�X�#!;����-�!��I�tmM��#��OR�fi�*KՖ6%�6:U�3l�u�=Lgl]�\�֎e\�s��Us�p8L�M�m�����ww�ܧ�����;b�k�ݍJ�����wk�^�cQ��	ɺ�	ywlsLjb �2)�q��~���t���z� ��RG�$��ljG�s{2���Y�s��@;��b��b �(��2'�i%#Z��M��z~���K˯�[g�
�+�m��Q��f��� =|� {2���>煤i2!���q�/uz1��@{���� 鼙Zm�Y���X�J=uΚ7o\v݆:N������yN���n{p]`�Uk�y����~~~S-�{\s�s�UY�Y�~r�np˚�f��5s35�iȖ%�by����rN
� B0A�	B*~*�P!6�i�7��?w�m9ı,N���6��bX�'�}���r'�L��,O���9u����5&����M�"X�%��~���r%�bX�g�w6��c�2&D�_o�v��bX�hw�zn�h#A��T�(�eCWE.�Y��Kı<�~�m9ı,O��}˴�Kı<���m9İ?"̉��w�m9ı,K��K�kX�N�e��᠍h#C3/Z��bX�'���ͧ"X�%��w��ӑ,K��=����Kı/�}�kY/c����b�O\Zû��6�`���a��h��5�ST��#tBv��n�[M~�r%�bX�{��6��bX�'�߻�ND�,K�������}���%��w5t8h#A������e���/Z��r%�bX��~�m9ı,O3߻�ND�,K��r�9ı,O=���p�����h{a?})�����.�k6��bX�'��fӑ,K���ܻND��u �$���@,M������r%�bX��߻�ND#A����)�!0�It8hX� �'�}���r%�bX�{��6��bX�'��{�ND�,�lO=�e45C}��v��J��b��9�i7�}#�g�fӱ,K��߻ͧ"X�%������r%�c��}��|�� b���b���[v�M�6�Z�7[t���C""RB%��^�!�Ԛ�2�ӑ,K��>�siȖ%�by���ӑ,K�����m9��F�}���p�F�4��3J�E�.�]�Zͧ"X�%��w�ND�,Kߏ�ٴ�Kı<���m9ı,O3��6��bX�%�~/f��-�5���k5��Kı=��}�ND�,K�~�fӑ,~!�2'���6��bX�'���m9ı,K�zN�j��-��
Ct8h#A�����,K���ͧ"X�%��w�ND�,@E����}�ͧ"YA�׃X;e��l����AD�,O3��6��bX�'���ͧ"X�%������r%�bX�{��6��oq�������d�vK�.���7k�c.�q��;m�ac�p�km��f��L�\M5��t8h#A���k��bX�'�o�iȖ%�by����|șı=�w���Kı=��aL��E�nGt8h#A���fӐ� G"dK﻿�iȖ%�b{���6��bX�'��{�ND�,Dho�O��4����7C��4K�~�fӑ,K��>�siȖ%�by����r%�bX��k�ݧ"X��F����$H��	��7C��4K���ͧ"X�%��{��ӑ,K���_v�9ı,O}�}�ND�����T�(�e@d%#�4�ı<�{��r%�bX|�~����r%�bX����6��bX�'��{�ND�,K=@�?�>�|�p  ev�.�o-��w����g��Y`*�Łغ�H��
�gpp�,PM$j�wJ5lN��q\�l��Jwf��;&�S����$���j]�6�Nj�<0`�vA��v���ݐ�'nv��^V��ۭt�Es��v��� ���P-�F)^�յ�<�^kP�I3���,cs�/E���[��`�n^�:�$�+��s���w �0�u�2S��em��WK��q����|:{q�8�����.��t���Sۀ.�\��{��bX�'��m9ı,O}�}�ND�,K���ͧ"X�%��{����A�F���t�C18Ke����r%�bX����6���TH�L�b}����9ı,Os�߳iȖ%�e�m�4��hk�ץDQp��5��jm9ı,O}�ݻND�,K���ͧ"X���=���m9��F�����p�F�4��	݊ά�\�us5�]�"X�%��{��ӑ,K��ӻ��r%�bX����6��bX�'���ݧ"X�%��u>�K�G
,8[r;��A�F�|6���,K�~�fӑ,K���}۴�Kı<�{��r%�bX���ɝ.V�(7<klOkSα�b1H��ݓq]��o�|�������`#��47f��B�^Zq<�bX�'�w�ӑ,K���}۴�Kı<�{��z�șı=�oM�᠍h#C��k�$a��0�˚�ND�,K�u�nӐ����MD�5�����Kı<���6��bX�'���ͧ"ʙ�[�|�(�e@d%��4��h�>��6��bX�'���fӑ,K��߷ٴ�Kı<ϻ��r%�bX�������n�k.d˚ͧ"X�%������r%�bX����6��bX�'��{�ND�,�"{��~ͧ"X�PF�߾�!����
Ct8h#AD�=���m9ı,?"�u�߳i�Kı=ϻ�6��bX�'�o�h᠍h#C�DDiehA		��KdG���[k���umqe��CB�*�y���X��O,*"�D��$7C��4����ͧ"X�%��{�siȖ%�b{���6��bX�'���ͧ"X�%��ڛ��,:3*�K?=�[�oq���}��w6���#�2%��N���r%�bX�����ND�,K���ͧ"X��F���YL��E�m�t8h#AD�=��}�ND�,K�~�fӑ,x�>�-5Q=Ϸ��r%�bX��n���A�F�棩��b�<356��bX�'���ͧ"X�%��}��ӑ,K��=����K���ȟt�?M�"X�%������ճP�&jMj̹���Kı<ϻ��r%�bX�g�w6��bX�'�o�iȈ�F�4;�7C��4��`�z�e��ɃZ�$��������w#�GnLY�t��J,\��N��UTҺ:�}��Kı<�~�m9ı,O�>�fӑ,K��߷ٴ�Kı<����8h#A�[��!�����R;ND�,K�O�ٴ�Kı<���m9ı,O3�w6��bX�'��{�C��4����t�C11e���m9ı,O}�}�ND�,K���ͧ"X�%��{��ӑ,K�����4��hk�ץDBp��@�6��bY�D�_��6��bX�'���ٴ�Kı>��}�ND�,@�~~r'y��&ӑ,K�}	�a�3p��)�᠍hX�g��m9ı,O�>�fӑ,K��߷ٴ�Kı<����r%�b�� Ud���-DKNY�5LJ����v�ԮC;�q�ϛs1�6�a���]m�Vp�(� m��C��4�����4X�%��o�iȖ%�by�����Kı<�{��r%�bX�Ͼ���5��F]�a����Kı=���m9ı,O3�w6��bX�'��{�ND�,K�O�ٴ�Kı<���洑e�˄ȋN��A�F�^滣�,K��=�siȖ%�b}���6��bX�'���ͧ"X�%�~�����8�#b���{��7�������r%�bX�z}�ͧ"X�%��o�iȖ%�by�����Kı/{�;`���(�-8�h#A���r%�bX����6��bX�'��{�ND�,K���ͧ"X�%��]�������� lm+:�Ăq1����u�9;D6(�;qBY�#-��c8ح�<�4�#��r��lV���t喺8-�7n�F[u���p��vv� 5���M�N������KG�Cp�>�A�X:�D8�vЕ�`�9{i�Q6Q�w.xy⹷�����a8 2:!���K��ؕ��gq�s�t<��X�����Y��i�ˍ/#{����|��6ў��c:�N*�؃�P��v0�C\/gn��9��˺!;E���Z�ND�,KϿo��r%�bX�g��m9ı,O3��6��bX�'�2���F�45�kҢ!8TI���jm9ı,O3��6��bX�'��{�ND�,K�O�ٴ�KĦ�����p�F�4��	͆�E��k55��m9ı,O3��6��bX�'��o�iȖ%�b{����r%�b����t8h#A��Û)�$���fӑ,K�����m9ı,O}�}�ND�,K���ͧ"X�%��{��ӑ,K��w���sWXh�F��fjm9ı,O}�}�ND�,K���ͧ"X�%��{��ӑ,K�����m9ı,O�wG{��Z��m��#!D��ݧ���C�'���،��m۪�<��95�t9�2���Q��׻�%�bX��߿fӑ,K��=�siȖ%�b{���6��bX�'���ͧh#A3uQBʂ(�NGtr%�bX�g��m9(�*0�P��Ati�K��gw�m9ı,O~��M�"X�%��{��ӑ,��h-�Gc��PD�E��ᠢX�'��o�iȖ%�b{����r%�bX�g~�m9ı,O3��6���h#Awt2�L@�i �7C��ı=���m9ı,O3��6��bX�'���ͧ"X�%�����rPF�4���*"�Ę�$7C�,K��=�siȖ%�by�����Kı=��}�ND�,K�~�fӆ�4��y�aq���2�!B͡�^۲qF/ �rCͮz�T^�j6cq�.6��[4cj8dq��F�4:���9ı,O}>�fӑ,K��߷ٰ�<��,K�����r%�bX��;�,�d�"ā�#�4��h{���6��bX�'���ͧ"X�%��{��ӑ,K��=����Kı������p���u/-�{�����{��{��6��bX�'��{�ND��z�b�>$|!X��2F.݊	{�h �< ����b< �"�e!BD!)!a	�)�IiB�)'�2>#P4� Ȱ�(`,�Č ���GX`�a������Q"U�� 	 �ĊU��WZA��a��!�*&��-Q�/�{�A=POD�V�ѣg�)ӱ2&��{�ND�,Kߏ�ٴ�Kı=��/�$[@��2"ӆ�p�F�4���{�ND�,K����ӑ,K�����m9ı,O=�}�ND�,K�3Z28���P%$wC��4��3߻�ND�,K�O�ٴ�Kı<���m9ı,O3��6��bX�=����|7�O1����m���8����v�7g����x�9�Ynp\]�ۜW,�.��ND�,K�O�ٴ�Kı<���m9ı,O3�w6��bX�'���ͧ"X�%�|�I٭C5n5�e�֦ӑ,K��߷ٴ�Kı<����r%�bX�g�w6��bSAᗦ�p�F�4���*"�n��֌ֵ6��bX�'�߻�ND�,K����ӑ,K�����m9��F�}���p�F�4��	͆Ĺf�]]M]k6��bX�'���ͧ"X�%������r%�bX�{��6��bX"x�Ow���ND�,K�tql0�d�"ā��4��hg����r%�bX�{��6��bX�'���6��bX�'���ͧ"X�%��ߟ��kax:��N��/m���Wv�F�2m�&��[���%ƱS��bz�\�]�"X�%��o�iȖ%�by��siȖ%�by����r%�bX�}��]�F�4=���I4"�sSiȖ%�by��siȖ%�by����r%�bX�}��iȖ%�b;�7C��4���f�dqE*4K�k6��bX�'���ͧ"X�%���o;v��bX�'���ͧ"X�%4:���h#Awأ$��L0˭fӑ,K?������9ı,O~��M�"X�%��w��ӑ,K��=����Kı/��;5�f��F��K���r%�bX�{��6��bX��>��f�Ȗ%�b{�w�m9ı,O~�y۴�Kı1 �������i��馭��IKv�M���=e�t�n��#���'d˦qm;��=n�;7lu�Om�>۳۵v�9K�V�S!)��חF�{X�D��5���ؗ6�eE���h.}��,��nz��Bص�ZТ;��]7*�Jm�8i^MV�`){��n㑃n5�'Wesu�s�d�
\7�tµn4s��ʑ:ާh�ڿ�w��wY���k��;6ݮ��@��l��a�W��c6��8v�f� ����،Ґ]W5OS�%�b}���m9ı,O3߻�ND�,K��v�9ı,O=�zn�h#A�l,�
aƔpǚͧ"X�%��{�siȖ%�b}����ӑ,K��߷ٴ�Kı<�n���A�F��[1�$� y���r%�bX�}�����Kı<���m9ı,O3��6��bX�'_�]�᠍h#C_��r�D�����m9ı,O=�}�ND�,K���ͧ"X�%��{�siȖ%�b3&=wC��4��{4�CM˄�˚�ND�,K���ͧ"X�%��{�siȖ%�b|}��v��bX������F�4;���K���E�sn�H��l�����9�W71m�����קpP�&�"�.��)�����{�K����ӑ,K���_v�9ı,O=�}�^D�,K��{�ND��F����(��E0Z����b|}��v����PVE�i��%����&ӑ,K��?~��ND�,K����ӑ,KĿwA��q& �E9t8h#A���m9ı,O3��m9ı,O3߻�ND�,K��ͧ"X�%�������)��m������wv�7�;��7�O/�w6$�H�����pBhi��e�4��hn@sa�T5��Y���fӑ,K��=�siȖ%�b|}�y��Kı=���m9ı,O3��m9ı,K����5�nd�y�:�����Q�O,��9<4]k��짜OOT����:u�֊�,��z�Z~��{�D�,N���m9ı,O}�}�ND�,K��{�ND�,K���ͧ"]�7��������a��.���{����bX����6��bX�'���6��bX�'��{�ND�,K��ͧ"SA��K�1$�M���4�4,K��;��ӑ,K��=�siȖ14D�!!���ț��ٴ�Kı>����r%�b#AwsZ28�����wC��4���=�siȖ%�b|}��6��bX�'���ͧ"X�%��w�ͧ"X�%�{ߋ�]a��՗	�5�ND�,K��ٴ�Kı=���m9ı,O3��m9ı,O3��6��b�oq����S����箸���ӡ{��d�g#�p������9�[�N���NGa�Xe����r%�bX����6��bX�'���6��bX�'��{�ND�,Kߏ�ٴ�Kı;���˫3Z̺�F��5�M�"X�%��}��ӑ,K��=�siȖ%�b{���6��bX�'���ͧ"X�%���'��3J�Q���p�F�4����t8Rı,O~>�fӑ,K��߷ٴ�Kı<ϻ��r%�bX��S��Z��Z֬0֌�ֳiȖ%�Ł�>��~�ND�,K﻿�iȖ%�by�����K���������6�[�oq���?���kOAu/-�x�Kı=���m9ı,O3�w6��bX�'��{�ND�,K�O�ٺ4��h{6ވd-4�P2�H8�\\]���GUv��²8�n���3�ۗhĵh*sZ8sl���{�����{�����m9ı,O3��6��bX�'ޟo�iȖ%�b{����r%�bX��jE�(YP(�#�4��hu���ӑ,K�����m9ı,O}�}�ND�,K���ͧ"X�%�wp-22J)AL�wC��4���>�fӑ,K��߷ٴ�Kı<����r%�bX�g��m9ı,B��:d"�0�!Hn�h#A�߷ٴ�Kı<�{��r%�bX�g��m9ı,O}>�fӑ,K��5�Q#j%�9!�4�����ͧ"X�%��{��ӑ,K�����m9ı,O}�}�ND�,z�w�w����w������?�� {=��Ψx�a�ܦ��d��f9�ɛk�c�u�Zأs��0�f���Y�V11��f�%��s\k���n*�Yd��-j�=��D\Of�v���Y��q���[�6F�iQ��.ri����Tg����z��s@��=
��֍��uvv���!,g`y�c��;q����F��Y퀺mx9"3�����N��,b@�v�]�{���w{��׋f�5&��v��Ogݯ�k�ݜᵍ�e�E�E��h۶�΋�YX.��f����oq���?g����r%�bX�z}�ͧ"X�%��o�iȖ%�by����r%�b���o�����7=\�?=�[�oq�X�z}�ͧ!�T��2%������Kı=ϻ�6��bX�'���ͧ!�{��7����w�Xbz�ym����ı,O=�}�ND�,K����ӑ,K��=����Kı<��}�Noq����������@"��|�r%�b؞g�w6��bX�'���ͧ"X�%�����r%�`�'�����᠍h#Awڑz�TJ)��9ı,O3߻�ND�,K�O�ٴ�Kı<���m9ı,O3߻�ND�,K��y�Z֦�)��%�e�2N��^��x4cc/:9��J��zʡ�wn.gw�wo�o�;cb�����{��ı=���M�"X�%��o�iȖ%�by����"X�%��{�siȈ�F�4��!f�1��
Ct8h�,K�~�fӐ�~RA��WO"r%����fӑ,K��>���r%�bX�z}�ͧ ��bX�ώ�d����f�=�[�oq���}������Kı<�~�m9ı,O=>�fӑ,K��߷ٴ�Kı;��Օ��lT��}oq���{��}��w6��bX�'��o�iȖ%�by����r%�b���{�siȖ%�bfm�RE�DCێ�p�F�4��O�ٴ�Kİ�1�����yı,Os��ͧ"X�%��{�siȖ{��7������۩�OD�'��α�cF�s�y��T2HE���ڛ�4lD�=�{ݏ���S�1�F�p��F�4;콛ND�,K����ӑ,K��=����Kı<��}�ND�,K�~�~� ���|�}oq������}��r"!bX�%�߻��"X�%�����r%�bX�{��6���X��F��"��,��wC��4X�'���ͧ"X�%�����r%�"+�*�4C��O���m9ı,O3߻�ND�,K��Yۭd��tjۆeֵ��K��<��}�ND�,K�~�fӑ,K��=����K�� �ș�����"X�%�~��~��p�.H]jm9ı,O=�}�ND�,K���ͧ"X�%�|���iȖ%�b{���6��bX�'�MXt�^�SF�I�e�r���Eۮ�B�7k� I��#��Y���8ܱ���{��>]6cI��G8n�h#A{��ND�,K��{��"X�%������r%�bX����6��bX�'{���ZX.�F�O�w���oq����{��!�@b��L�bw�w�m9ı,O���M�"X�%��w�ͧ"SA���'d��$��$	�%��bX�'�o�iȖ%�b{����r%��bX�g{��r%�bX��{�m��7���{����5�'������,K�=���m9ı,O3��m9ı,K��bXT��)�~T��"gM�ɴ�K�F�{4�CM6��(SN��A�by��siȖ%�b*�{�m9ı,O�>�fӑ,K��߷ٴ�K������߿��F��(ջZ^��s�f�;��tv�Ş����vb6)G��f(�`����4��h.�v]D�,Kٴ�Kı=���lEyı,O3��6��bX�%�~GT���PB�	�%�᠍h#C�>�fӐ�@W"dK﻿�iȖ%�b{���6��bX�%���[ND�T3A~����c��$��᠊X�'�w�ӑ,K��>�siȖ"��b_=�u��Kı>�}�ͧ7���{���;�����v�|�r%�g�T��=�~ͧ"X�%�}���m9ı,O��o�iȖ%���{/M�᠍h#Cr��Ġ�k.j]f�iȖ%�b_=�u��Kı>�}�ͧ"X�%��o�iȖ%�by�w���Kı>_�&��S�<ـ�D�b��&��@�D�ʒRBR0�4�(@�����~f�O��$�P8�5��)�@�A��`G!�AJȸ�H�5T�4	'4m ���IAH�� *E���B2J7�\�t��yU
H��!Ŋ�J�#�lx f(s����!H�P
B,��B�F I�@�.h! �M	$&�4�0�������w]����;���l   l      6�    �j	�e�T���9�c�z���vX`����˻q/K��`�Yhl� V����vye�j����s{d�Z�S���;��!h���7V���mlڶq�f+"��pY��6G,��6�1�;�۞�r�f5� ��ɓ*I+��29ђ��:]��q�^[��Ki:p&39���[GA���_�����1qrK�g��ic����h�ƨ��0RVwJ����6%�B3	"���mc�׷<A�`� �A�F��l�]�YI�
�*��l�ҫ�-UU���/0G��Wl�[j�L�V�KUgq��d��:V���B��][H�m�o���-�
9&@]NuB �M�c#!�����n���^F����ݞg������+$뎪�/l��D����hq6��*u۔t-�����nY�ؓ`�#��V&��u�ga� ��:c8`�a<��!��e�%^�(�9v�f�a��(^F|8̼͢�e);7<JD�:�e%U���g���5u[�D�]��s� ��A��$7Dl�2�ū;��r�l
��W��y�H�5N� �BԠJ6�)2m���l;s�F��-��.�n�Tl�k���8��Y��H<%�m��ʅ*���ʙL�hتD��ȝ�T��� I�lIڹ��3�V�Z�ݸD� 2�UD�n�mj-2���]�UT��T�����as�j�H7n3T�J���n�M��*��ɽ��;4�UW&ң��ݕ���(n͖�7`(BZڪ����[m�V�:FkR�@F�ȃ�pݳ��ݫ��Gjw����jWTJ�y�0��%���j���G+S=���K��"EI낪#&Fhɷ/��UM=��X
�! -��tmu�+��:kj�Jһ0[�lmdK�ڪW3��mgnB�hl�;��j�V2��u�*��!�Ъ�k�\Y�9�lK�X�Y�f[��]XddD`(
�x;U(��GH/��SG�ww����k_А��nbK��v�d\v��/fw��m�M��:�vcu�p��e���uz�؏�ۑg<�pa��$(מ�h���<��������X�R�9�\v���Wl��NG;��@��Ӹ��u;/;g�8��Nz�kn��Ě9�������9�����8jr�mz��W p�IE<V�ݳԹ��u���A��a�g�N����vn���Y5�5����=�s���'���s�8;]�7n�1��Y.��xz�����V��@�3֋��ki�Kı<��}�ND�,K�~�fӑ,K��>�sbȖ%�by�����Kı;��'sF�j�-ѭ\���ND�,K�~�fӑ,K��>�siȖ%�b_=�u��Kı>�}�ͧ �bX�'��ٜ�շ2�[��2�f�ӑ,K��;��ӑ,Kľ{��iȖ%�b{��}�ND�,K�~�fӑ,Kľ{�f^�j���I�.��ND�,T,K��bX�'�O�ٴ�Kı=���m9ı��;��ӑ,KĽ�#�FIE(!I�Ԓ�p�F�4��o�iȖ%�by����r%�bX�g{��r%�bX��~�bX�'�G����� LB�d��D�KU�[�nskG�r'5��k����Q8Xퟝ�gO�;I%0�%Hn�Mh#AͿ��ᠢX�'���6��bX�%�߻��"X�%�����m9ı,N��s�Yn�(�d
8n�h#A{���6"z����C�9Ļ�}�ӑ,K�����6��bX�'���ͧ"~L��,O��?~ՙ��tkZ�fj[�fӑ,Kľ����r%�bX��>�fӑ,Rı<���m9ı,�׻��p�F�4���N�fIkE��kiȖ%����>��?M�"X�%������Kı<�����Kű/���m9ı,N�d�h��\�E�5��3SiȖ%�by����r%�bX�g{��r%�bX��~�Mh#C�r���F�41�c�"��� Ě���y1�D{m��v�.-a��t$���]և5W(N�+o���F�4�׻��p�F�4�͜$�M?
���fύ�O��?CP�	�3q {��1��@z䘀%�T�����C�ԓ@�)�}��EL`�@Wbfr��ٹ$�߾�䓹�ᑢA��h��6O�*�R���:�~����9�`� �d7.��A��4�����4qҚ��M�W`����q��H���L����s�vG�ú�Ty�h�z��f���#��%#���h�4�Қ�����y$�ǒbmɠs��{�I������UU��ug�2'y1)�&7�g�@�[^���?�=���:�~4{��D���Qō6�|��@>�Y�{���衸 �؊mD���߿M�'���&~�Px(`�@>�Y�{���>�Jh+k�>�qDX<q(��NKmM�5u��Ų�x{릻^�����*��3�fǸ������C�ԓ�:����{�I�����n���Ja�JpY'���zG�w]�O}�,��u��
vWH�q)Lo��>RL@�5����p�� 9�� #�-�i�L�������4�빡<�'E
]{�쓙���$̒"ݫ���t����& s��&/�	�~��"�d��Ԛր���t�D��\�KuF�DXm!4�:=97\�e2&����6�Rbȓ�۵�p5�hLu� �y��<��o���{s��tW8����g�5�;���닚�ۃ��<[���H�vx�v��h�5���O)]�l<F�*2\;yA�m Q�&�79��&�/`���<��t�;��Z읁S��]��p��m��ln*�f��Y�fL����G����3��|qv�']k^��������6h�d�v�Λ��v����n���y��'w��<Y��y�d��
��ѿ�����[H���X�n���'���d�x{,Y'���z(I�j	��Px(`�@������sO%�t�|��@;�g3 �Ǎ��~����ۧ=H�7����1��1 t�ᑠLN�h�I�}0�'hu������;���{����ɂ���5nܺ�cEqɎ�^�v�gG
]��8܅���L�D����h+k�>^�������?����&��y�w��� =|�,�����n�T��{����$[�a�F��H��&6�z�?*@{���b��b7w1T�<����&h{�4�Z����ݝw4{��D���Qō6����1�������R��t�~;=�NӂU�6�<���;�ݵ�^9�۞�.w�ݛ�l��[e��NZ,�-����@z��@s� =�`���19�d�H�00ڑ�'���
#�d�d���vI����+��;�����19�_��h.��?�UX�
���K��d��fX�I��dm8��d��9�ֽ��@�g�œ�UU�e�N�v&��1�-/wq��1�N*@{���nb6ߝ����hT2\Z+��n����;�X��c�5�;uӲ��]JY����:6K�H�Tn�ݬ���ҧ�Hs� =m��=a���~��/�'y1)�7�L�>�JY'���d�.��y����P��9��{"Clm(���p�9~��z�ֽ�λ��Қ����
	@��vI��c�O<=�,���a�P��@P��^;$��/!"�����N*@~n/ǀ럿b��b �9S����箹g\]uv��q����l�8�Of���6T��^��ԝ�6�e��R���� =}&~��*~T�??<�N%"Y��h.��/Z��e�$���o�*�	 st���0d�(Tq�'�ۮ�=��X��@
K�g�@�=��Yrd�2Lm��?�ܩ�Ԁno��rb��bNJ�H��<����&h�Jh���|$�{u�'��I�eQ�w��$�U��&
��ml�\o{p�B�絨y��ݹ ���]m�]:t sklpP�q{r��%�P!�1��<\�]��qT���*O7��N���=�rD���ڧ����ʺ*22s�48�/@�kRg�mɲX-��m�AA�۩xE��f�.MJ�r˴�냳�m����1��qȝ�Vr�0=&�px�-e�ۀ�v���m��>|~u�&\����F�\�QcpOUm����d���`�n۳�F��ȋ!�6�qcm�x_���>^����X�q�d�d�����b
�E@Zq�'�����*�9�b�>�M6I��W�����a�JF4ґ������[���u!��m�e��^m 9���rb����Z_�f�~.~y�6�JD�1�9��Ɉ[��*@sqR �.U��N�6�m�vn�N��Ok��뵅:��n�vrr�(@��zh�o��uv�|�,i�<N>z�u�'�>�Iｖ>*����נ~��a�F��$FL�n=�빫*�E~��@پ��7$����䜾������K��8������u��Y'�َ��PK�7]�sm�$����E��6�qciɚ˭z˭zx�a�v���/M�O�ga2&
qjGd�/f;$�B��a���O�6Œ|�נ[��$XbqG��7$H�u��{;�p kc�u�����hWɵ������>F�BS�Li�#�K?��4�Z��Z��-$x��pC`)�{�L7𪪡�P��ϖ��O���N�4��卦E���9��߾��9}����|�j��1!�*�P�L3�ȑ��E� i�$HC-��A��`�H�e�@�	BCS��VS2\ �n:P�P�
�X��DV�B*P#Q �V'��,��,"��`%R�f
'���P 1!�l�@�t ���P=D7T����(��⾚��޾��y��lܓ�f�q&Lq;'@�^n���Ɓ��M�mz�adjI�4a2ێ�=���d�T({2������|�נ}�`����'%�M�{]�u��5`OgvM��v���~�m��!H��ӔJL�'p��bp��~4�������>ÓM�}���DhmF���p�>Vנ|�נ{��О���  	�iL�&F�N�*=�\��ǰ@s{�I���/!"�
�JGd�P�K�r��3߾�f䜿}�n@v`@V?�"�Q
bEHmF
�ӝ����~�I��m	�)���I�[�ǰ@~����u��m���ۮ�v����kW{t.�Xv���@��pn�u���;N�=�w{ᮟ�A��u�a��p�����rb��})�ya։��L#�o��.��� H�M6I�d�d�,�vI��H�p��a&&�z��M�Қ~�T���d��ݖI�y)�D�Q����p�?/f^�$�n�I�%���b�]�h���$M��Ҍ�i�h�& 95�{7�@}U����� �ۮt��-��9R��Ɏ�̄[1aѤ��{N�e�t癹]Y�I�k��7���m"S�5�)�k����skI���kv�^/91T�:od7Vq���3�f�cZ�U�5�`넌3��7;kf@ vm�@�Bu�tm˸�0�nn��tR�*3��sx;�ⲩ����`%���Z��z-RL#,�z 
·nDM��L����/np��k���۝��bm�F���%�j.�����v>|ß��v��V� ���ڀ������ ���0�%1Li�I4��M�ҖI��c�I罒��(U}UB��'�>���D�6����߿O�|�W�wY�}�Jh{+�i3"�X�Ƥ4��(U.��vI���d�x�a�O=��ya։��L#�oq�.�����_t"�x�\s�ɡ�E5�g���u��v�v�Ծ�"���۫X'���ԧ3���ROT�\-?6�_������ =m�@Nw{ۼ�L��y�L7 �,V�UWg���@-����)�}�ܑ&<mF���O{�x��vv�U��&���� ����'�8�0rG�zۘ�����?}�}U}���@�	���P(e'�y���?
���/���>]�����\PdX7Yñ�uXru���tr��W":���ф�a.&G?��	/��M�4��4'�=��<^�?���"s�&�$��צ4���,hcR��z˺���0�'���{UA#�n��q&L�&�Y���� S� ����� %�#Q�"a&&�z�?�^�-���@�^�@�wW�_rR�$�`�o�@��U�|�W�|���;���~�
�3�%6"4�q�����{.6�6۲�^��b�rt0̆7&������D�<mF�I��9�����@�c���Z�Q1܊q�`�@�wW���"�;�h��Z��z��j�bSƞ$��;����}V����=���@>촑����m$ёŠ}Ϫ�>W��>]��w����ʰh�z�`��g.v�Z����i3	LI�8���[s���9hnd�7 �s�qy�ܯD�����
윗%�u�����-��/�y�a�X^��3�m�~~~�1>�~�d�y��D�nk�N��vF�D�������}V��>�@�^�@�wW����z�1���X�P������
�� 'V9h7-n�U�X�Q��'��^���@���hs�ޢc��cNcS$z˜���Z���9�U�}�U}�_����H �`7d&j��UR�<�.wc�Ê9wg:��î�'m�۰5���d(��N��H��lV�v]9e�z�,��F[[A��cÇ�S:'F�V��uΜUY����.%繸-�m���6�49�g7m+GD���X�;�=S<���َ���EnѽR����٧��3;(���\n���V63���8�8Nq�Lc՛څ[�����z��F��ΉN��nK]�)8���X#\<�젦��Ǭ''n��p�bu���O����*$�w������Z��z˺� ���G��8D�I�#�@��U�|�W�|���>��Z^��L�Ec�-�z���^��K�w��=]��,;�&���RA7�8�?/;=�w��>��h+��م���H�2)�r=�U�}�)�|�W�|�נ|����?䉑�7�!������Ōnrm������NW��t$O�e�}r�0D���:���>W��>]k�>��Z������Q��93@�㘺��η <�r��T�::�;�A�RL��.��p��?�/fm�$�nk�I�q&�i��6�����l�h'�H\s�& �-$x���M$�"8�u����z�Z��}V�{�����r`����tRv��;�U�r���1��	��;�m��=�7�Ċ,hcnf��^��ֽ�U�{���<�n6�I̬��@u�1�c���"��8�zadiBH�L�n=�U��{��74��lVC֠UbHRA"-E`�Z�J�h( hPvb��;$�n|쓝�S�8��!���~ٻ�d���vI��@����>�cPCj1��$I��c�N�*�n��I���$�ٖ,�k�	�a(�y#P�BcbT6�ܗk�l��;f݉���gvϖ��:�$�t�E�� :ۘ����"��Uzï�����&�C扊bm$��>�r*@z㘀�rb����_��W��D�I��������z�?ٙ�r��=�w��..��_�j&$���$�g��'�َ�<�~�d���_	T �,T ���~��z���&�����7�8�+k�>��ZwJh+���μ�&���R��Lܓ���ۭ��Sǰ��pm; ���s�;h8��d�T����E�	=��U�}��I��c�
��r����?w��D�Q�K&8�7��9h_I�\���_����~[�Ǎ��bqh�~������JhϪ��I�q�<jdd¤����(׹��=��U�}��VO�f/?�����5�3&@m�#�>f9h��=q�@z䘀U�}_U��#�AMr�UĨoZWI BB]���
�ib$(q�H�R�Q`0p�M��c	��E Z��C �a�� а�i&�S��SA$"��M��.!: "�M�
BB�A��$j�gOt���=���$~?f�  	        6�    zܹ.���v���1ҧ 4UU%nM�Uǝ�k(@��d��>��drV���.y4������٣��).;�=����;T��
��Χ7`�j������v - lb2W6�*�.��D"�U��cK��l[Qi��1ی�K���kF���%X���6�@p88�@�y������)��P��t���Ɲ�L�eRT6q�ڙ:�BN�h"i�btL<q��ݎ�ؐ�74띮`k��iz�ӛx^(%T������ú�e��M��+�;J��J�N�-��Mt� �]Y��3m��T��lֲ@UFڕZ�F��a��V1!`��p=�6���� �����,�����N2ݷ����b�Y����g��9�KL��D8��N� ��de ��}�`"j��m��)j�
4�S��7
��8J�Xn�e{����j�R��;��.�5�t�!@��mmJ�M�-ѵ�G,9y���j��'@��@M%�H�!�90�ݠ���T�&�HȽO2�չ��T���Р-QT��f���UJ��s�܉�mH�ƺ[���.����A�@9����c���/O*�&En��Q/(R��7��2l�;=�`ݸ8 ��ն�xݝ�t���H�N4�+I����m��H�hpӪNЌ�UUgt!�<�ϰr�΁�+�Z�A[;��)�ՑZ��wim��[J�Sm�u�OZ�I�F`���g�6�nS��vCn��ףR����Htձ���ԗb�m���N2s�`����mnU6��z��Fơ��<����nI��p�2�=����p�b���q]l�4�9H���0
�Ya��[<�>����ѹ]�k���'K$��[�A�*�Ga"��ڪW=t��Ǖ����c�g�yU�@K*۱:Z�G0S)�<Z�W
ZVKn\5��[l�ў(�")��j<@6m@OC^.� �
�����=��&���(���k��MjMkZֵ�fcUNM���ဓ�#����:�ڮ1rY�9�sϞ���u�͝V-E�JJ����m�z�tvݬ�&�v7j��`�ٖ�r��Bm��%#��[.�م;Mǭ�^E���u���<:�J���{b����ƭ���8��B��:��b��%1h�L���y��gk��.yn�5ٴ��wWX%uj�z�B�m��M��A��r�ઘ�V9;y��g\=ut�����q��;��B�ٸ��2۞�w힭O��6"8��v��z��m�����i{�O������L�˒Z��[sf9h<��着���D��RA7�8�V�z�f��;V��^�oL,�G�D��49#���4��Z��z�>�����S�"N(�%���}m�b��b ��srV��^uvrX9��ы��X��u�w��i���-��1�*y���$�s�Nt������ s��<�5��- wK�OQ���
�;$�w�/�] �F1 ��H$#a	H�d @�X��~��ж)�x�=q�@��.iC1"d��7&�}�Y�}�j�>W��{���-$x���$�X��=�%�=q�@�j�]�S��?[�~g�#I1���^�{�f�w���>�hʮ,u`&�2�YqS��*qu�/:�{m* <dP�/�v��o��q��cq���Xӏ�9u����f����@�^�@��F��"�#3wq >�5��-�b��b�I��?$�	d��ɠ{���_��7*���$$*�xfc^]~z{-���8�m�3��ʹ�9���@��A��UP?m��I��&����jI�Nnj }Nj�$��9�	&����0[<vh�U)z�^��xK��s�g�����&��w������3�ݍ���.��'<3e�y瘬�Ş�� W>Y��z��ďA��r<rhs�h+��]��{:��$~]���GcLrE�y~�����^����M���� q���q�N=˺�$�t{%�y瘬�ڪ�(|�޻$����I2F
d���{:���z�uz�c,do$��X������$��m��r{;���B����O���$Az��x��`�/5�������ͷҽ^���_�3�쿦��-�<Cj1�ڎ��{�3�#����^��i'�Ɇ��l�}���q�Z�D`.H쓋w�d��d�� �sf�$�nk�I��a�1"d����C��%{/�{6i�O{��
����$�G�U�MH�ɠ}�S@�^�@��@�t{%�o�lUP m�f�L�I$�鬴�ZM�흓�V�{4�̩"�g%���<�ܽu���z�ZX��6����;h��n�:G��Y�/X�:��8�M�b�Sv޶��Yxc�,U�ϱy.ðnm7>�Cs䞒LZ�p��n9�wl�O��[�d6�m���.!�ю�uh"���|�� �*Y��׷��9��1�|��n^�Q��a�۪2�tc��!����qѭ����z�kc;-�;Z��k>sv�7ih��Y�n^��&��"�I��
3��4�����~��z�uz���T8��=�d� s5[����6����� ����$��9�	zadj8H�L�c�= �gY�}�qY�).��vI���d�dJE ���ɠ}�ՠ|�W�y{��������쿦��4��J&7���c�O��י������<��+'}�w���h�hLγ�-�y��G��ps�n��͛F�NЏV�͓�ԉY$�qa���_9��9�v9�U��9~���w���ĉ�1���@;��R������Oրv��@zۘ�<�CcŐs	0mH�ɠ}Ϫ�>W��������_�@/e�4
����/sm�b��b }NjݎZ�;� �I��M�N=��@���ي�_��=��Z��z.�܊b�^,�b�\Ŏ������ l�\u�w���%��N�ݹ�Q٬���I?��9�v9h\s�s�6�{�����rY'�~�U
 $z�5�'�_�@�r�4��lj<q�6��O{�x��vlJ�T*��P����@��~4�s,�LD�97�s�5��-�b �p�0F$O鍴�z��4����z���@�"⃂qc7������=@���\��I��`}K�;^.�&HH�d�LR7&���U�|�W�|���{��*�sʢ0#�-ʹ�9��v�h�5��o睊#��n$�)4��?.���w���}V��z��0�5$��#�=�ٙ�^��h�-��z*0U>F�8 �����nI���I�I���4�����vI���$����:*�
��\&"[GLaY�2g�t;m����ױ����Նd�#z�)$��Y�.X��~߿���s�5�{�xM2���ڳt��@z��@����]��אՆő�16��@;����q�@z��@u!��u�F(�ԎI�}��<�W�|���z٠U��Da��%!�y^����I�s� 
�ﾪ�[�H �`76t����4��݀�n�ļJs��nN���ʺsț2��R�4���<�q\�8�\�$J����&ԧ6��'n�����F�~|�'�a�ó����V�A��zG��꺰6�V��d�WeDN���6��;jۉ�Ͳ��i�]t�˰#��l8�$8n��NxY�F�%6�]��n+;>�X;=�J\�/M�{ki��)v���w~{���g`F۞s��]Ek��{m�Aul����6^�7%�����Y9zלl1��;U��g���� >�P� :㘀�mcNLr!L�c�= �[4��s@�^���@��$I�& 87$@y����������n^���DlRf��z���@;���u��S�Q5�LD�97�s�5�qR�9�WN#~��B�W�Q�j(�;����vTCC��0�s�m�nLM�&Jݝ�N�37�5�qR�9�_9��J�x��1F6�rM�u�՟����	U"X(�$� ��,�g��'���d���K���:�1�Qbp"��������/uz޶h{����7a&D�4��>^���5�qR�9������6��v�wq >�P� :㘀�{��>Y�u�bO�D��5��D�����ɰ����);8��3����onm�+P1\n�f�����8������ �l�=�J�`�8�j&�&hW�@z��@����H����^�MLD�9#�>]��z٣����ً0� >��bT�������\P"���O��"B��X`B*�� �)
��(����Ɂ��\�&�,(@�J�(�M,�m��㳜D��B ��.)z6�n���o]+�(��W��"�>\A� =Qǉ�O�
 (_��ٹ'���^CV3Fd��N= �[47 :㘀��1�6�f�^����mH���s@�^���@;���:�װ�a(��D�`�Kں�c�`�r��Q�n3.W�[u�I��OZ.^�D�E1	9������uz޶mUPD�3lY'���F�L�My����1 >�Pn*@u�1 ���4��ȉ�LnG��f��u��<�W�|���/�)IqI���N�
w3x,�幮�<^�;'����gKf��T�6	�㉢6)3@�b�d������7 ;�ŃŲv#�R[�k����;�n�gvy�s&���l7oe�^`Y�TJt��j�*����t���qR<r�Ge���!Jp�q�$�s%褏s6Ő�]���uz��[�1�F�jL�����㖀��1 N�P�GG�Na"���^}V���@/����s@�uD��$Țʹ���t���qR<r��
��(�I�|kRkZֵ�j۠v�S�C;Es�gI��N�֍٥t�Z�nz谊K;q!ץ4�k�h	ݵ����`�&wNM2�]�)�w#�!�MW����D�8�q���kr]ʱ��U��k�&K@�	ۛ�K6i�lm�<v�6ލv��z��i�����$ݕ�9Q���m��e���������69�ٰ��k&{��lqԎ�����+[�m��M���\�ՙs_�i����&�b]t��w��x>K��`Œ��WPv���i5r������0�iˣ]25~������<�T�����;����mɄ��4���y�Z�u�}l�;����<$q�(ғ4��@nj �&�<�T�:;����<jb$��@>�@/����s@��� ��5a�3�s4���5���r��� 
����m�Z����9�������=G���oC'j�s{s�b�d�x�3����o����H��@zۘ�'9�	}�nD�2"�N$�_�\@`
�0���@>�f�{����n$�L��[��9ט��s��g� �3lY'|��w<:�i�9L���Z}� #qRv9h	�%��e�y��	�h��h�U�_;V�_[4���B6��GƦdX[[������'�l��kjƍ�-�9,L����/��O	m�I����h�ՠ�π �'s6ŒO��b0��LREd���W�@ )"w۲�;��,��~�
H�n"��E��f�n+$���[�}�l��S�U$@qG;��������}]U8�Cdm6�rM� #�-;$�:M@;��n��	�RpY'<���?P麸I;��d���Œ~4j��PD�"#r�dz��uOkĻ��oe����L�������,��c	" �I��@�_����@/����h��nD�Ƞ-�d��̗�I��I�y��9�j�;�)Z�r)�d�f�{��<r��& 'H� �^̽�/(q��Q� �~
�m���>[���9��I P�СT '��I=�,r4�Q�����<^�vI�U �w���e���^}V��}\����<lX�x�T�]/gq�a6���.8����� đPpk���{��D���!Jpґ�ݱd���y�^}V���^��uT�Ősi7yy�Hn*@G�Z���� *�Y�5�R�BNf�y�Zˮ;?T+�*����Y'7~�d�"}�F�L$Ț��>]k�/���=�w4Ϫ�;�r4�	�	n=�̱d�� W�7���ǚ�����d����ww�_���� 6�5��.���mӳu��ɫ��_�mjz�m�(���H[uY#u�//7ca8���$��LOm�V�nՉ�6����T*�a.��Qq�m3�^�Vq���h�M�p]Z�cq�b�r�2��t2e�<;%��Wm����n��pH���g��A�VԽ�6�u�g�\�����i�����Ц�1��0Aۈ曷l���[�)�4�Tv���2fˬ�ZѬ�-�՞���	5��t��p���擶��U�w��]bH�����K-�����f��������/>�@�u�@��s@�U+Q�<$q�TiH,��~��U =Y�쓾ݼ�=�w4וr4�A���"�-���� 9��9h��ɧŕ{�m�{���"�7 #���B�]y���gt���i6���@sqR<r��& 'H��q��`�1 0C��X�&.�v�s���Ĵ\���z^H��ٹ�x�ͯE$)e�m #�-�rbt��UW�W���4 �� �I��&Š|��N��T�t�=�R�~T���yC�ndD�4ۏ@��s@�u�����ٙ�~��Z�����S���q�d�*�ٛ�d�ǚ�����d��]��T�F���УJL�/>�@��1:EHn*@y�ܙ�{w�hLt�l�O{s�8^/m�.웯*3f׀0�v��7W���{��|�c]�.tU�/���� 'H���]^����Ga�O�*���3.�q ��h�j�c�d�/f;�B��G���q�!rFSi��O�6Œs�ج� �@@3�췠_[��U�]#k�LBNf�^9h[��T���_UU�?z�t[�n$�Lq���>]k�/���=�w4Ϫ�9un�X�X�����qZ�z�^�o% �waq�g�͖���6v:��vX97 ��n=�����s@����ֽ�tu�7	0��n8,��{,^� ($wj�OVn�$�r�h�j4'��&�Rf�y�Z�Ɉ	�*@sqR ��f�^U�nF)"�tU
��u�'}�b�=��œ��UAP ��3U�Nw/a����6�2�w�T���x�>]k�.W��qAĒn,�8�rB���j�Pڻa��	��}��;���j���9�4�M73@�u��/>�@�u���"w۶,���1�R�ͤx�=nL@N�R����q'��0n-�ֽ���:
��6Œwj�O���B�p������� 9��9h_Z�����na?�8�s4w]�<r��& 'H��g�WԺ�>����1C�x��(������
Cϑ�L��f h�O���S@�@� �H�a�d �-�����7 ��B0#A(dhB�$ְF�(6"P@�.��+b� @�
\01Va��2)$��C, ��P�h��@�@�BSFA!,Yp%1J�yv�D��+
뻻���^����� @       �     n�:fX[V��g9�T�pf�UJ*�z��c���B�w'�wj�z�فۏ���uj�p(>�<��M)���p�[gd���I�j��P�֌�q�����3u;b#�[�$��l,b�g[�a��K�R.�nC����ɻc�槑��7���V�m�h�[[l�p7W&�xz�%�j��󐗧˵�\������R"A��e�=��d��7fz�&���M�t&�9�5�6v�;]�1��yR&+����U,|�k|N>���Ӓ�)�N�m�M���v�%�bYN�i�]�(:N�T�d\� Hm��okB�6� 	�� U�V��n��=p��Q�!q�<�r�K��CR� g@�-۩��*��#��gMd]�T������t�6���8҂a���8�Xٚ�d�5Y˪�E*��j� �ePJX��/�������Gc�6�gg���Ȥ��-u	Ç�{S�g��ݑ����!��nu���F�8�Q�N�-�]t쪭z�_�����8�m�8�m�R��ƲumPUGk'I�Ͷm[e�06�91>�>J�iw���c����k��[l�������	m� �]���^��n �]5F�
������	��R��;��n�M�$�uq��:� UWU�C�+/<�YMQ����9��6$�k�%]l�T� ݤ���v[@iWbP�,�Jȓ-�j���HۖT8�'�$6�����6Ͱ'+�uv�D{]�'m2�e)���J��"n��U^V5nm�۝�]Cm�ʴ����R��#��%����q�s
�ӋsJ]9��+�F��ݧ
��)���@��L�@r5�жӎ=� �,�쫫�b{g�.��]�T8�7R�;S�)eq�٤Ȫ�KQM�pX�ͼ\S��u�{* �*���ldQ���%`Ŵ��:����	\J��u�ֵ�d ^�!��!��p
P
�����V��~�������   etݝ4E��ud�z�O3��-ШNs=g7!�PYغێӞf�)')"�=:*��Cq�2���mJd�c��x�t�ɉј�%��%���H6��Wg�-�p*�$ud^�4b�i#�Y�v�e�9x�'��8�sp�X:؍�$`�:ѮbK���W�?�x��� �s*vx�ˎ9��{B���G����A�55�����������6ѳ��\*k���V�v�������{+��nh�,n�t����F��{�����>|I0��#Rg�;���h+k�:���;��h�����
@���h+��� G76Œs3lY'������B��6N}���4Q
`M��N��X�O��g�UUIf��d���vI�3�\a9�cM$ۙ�wu��:��@�u�I�UPno�u`צ6��C#�i �9h����x	�~T���_���jx6[n<�]]u�/m�$���+�8��^#���u��u�8�1��s�ўٛh[�8���H1�@6��q����c��n=�]�������^
�B�����$��+$�{1�'�=,N%"�	�1�#��{��h_U�|�נu빠w���ОH4(ҐY?UUC�T��ߕ�|�}�����[ʹ�9F�RE�}nL@8�7 �-��{d�򓝧�B'�0�����[s�
�s���*�'Wn�g\�l��7:�B��qR���c����W݀���� �?��G��s#bm&����s@����ֽ�]�����$$x!\ѹ'�g�]�9}����1� � �H"2! 0B,!�
�BYP�hz�n���h�Z�'�$ȇ�qh�����o�;$����$���I�?b�N��A�721�i��׮�����Nk�VI��c�O�<b�tГ2%�Q/^���N�{�r��N¾��ᅹ��۱I��?��v)�I�����������Z˭z^��z�Z����HƔ��>��W�P�I��vI�ͱd�o*�m�
d�QI���1 ㊑��]�?*@O�?Z ��2i��P3m)��,��$�3lY'���ɵUUDUv�
�y-�'�g0����dlM�ۙ�{��h�̿��������w4�]�FLC���$��章N�ns%۔EGA��Nώ�v�����G	HE	9�W�h.��z�h�=j �K&F<��<^�w�I��I�fزO������k�n̌pcn=���4'��X��T�k�VI���d�w�dR%"�	�1�#��{��h_U�|�נu빠w��q<O�bDiI�c�+$�Uכ�����Iｖ,�*���{��w����������nÑ��N�S<����ƶ�����m؎���������:ؖQ��a9�F�/l��
5���e��+����b�㇑�v����H��ػ�f�w|�[�^q���4�2b�6q��&�3��3Ś�{�'����'nf��1���¹�ɷ*Qvm'G�յ�'3ֻ���sۗ'+t���`nN�5����a���{�ۻ��39;\���+Ԗ�[q�m���;�n	΅�m��d�a$�}���^*��j�4��.����׮��빠u}V�z�a�#&71����z�o���H�nh󿖁��^��e���L�	��s4w]����Z��w4
���4��s4��@zܘ�q�H?}��?z�`�~�F�X�21��Z˭z^�������Zr���64�2(�9��.����{[v6�mȦ��ؼr��3�M�m�z���7�LN$6������=�w4���>]k�;ܫܑ)�O�I$�$����U������>[���>�e��T���x$��&h_U�zܘ�q�Hn*@;�����W�FD�REd�כ��9�4�'��X�O��ޢ�a�#&71����zQ��H1�@zܘ�+���Y�^tm���P�WK��܏I��;/1��Þ,��i�ͻ2M�4HH��&I�4�r���$��Y'�ُ@D���d�Y��q�Y!$�h_U�|�נu�M��s@��D�cq(ǃqh/f;$�=0�"��@(�@� �@�A� b�D3��6>]}����?�h�� �����U���� ��� �9h[���� �Ra?�I$�4w]����Z��)�}�:��D�73����:����q�vv�Ȇ��[c��!�v(i����SGC�<�F���󿖁��^�ץ4w]� ���6�AI������=nL@8�n*@9�- �������i��z^��;�e�;A,ך��՛��<�s�Y��I6�hW�h.��K���?�2W�٠Uif8�,��r�c����1 ㊐�T�����{��9��:�0���z�Ɗ;^%�汸�u6��63�
�.=���c�������φ���6�2�;����@8�7 �/@�ǜ�A8���q�z�h�T�s$��Ɉ���Z^��ѵ�I�{�e�$�b��).��vI�߿nh�m'���$F���uv��ֽ����]o�@?~�����
L$IE$Z˭z^�����}�ج��U�T DU/W�Bd�IJ�T�L���t��=������
s8���p��Kz�::ێZP)[F����c�4lw<[m�
��kz���O��][���ƻ )�u��llp[c ���;�x6`;b��A6��/k<r���Y3Z��ۧ�z����j�9yx�q���u��]a��� ;)g]D,����0]�e}p5v5��OAV���{m�ksT�kF�ə�� �� ��o5�s���Ɏ"♒z:^����pe����ts���]Y�p��c���k��pS�����R���d����1�	A"B6�m�d���b�($s^�OVn�$�3,_�@PH��;�B$1J.��i?g�ր��1 䊐�T���D�h�"E�|�נu�s@�u���b����@�W� �M�J�ێ�>��I��Pٛ��Nk�Z˭z��1�Jbm��5�����{�ۛ���^�d�]4���>��K[�+�9�1wU9)�O�I$������-��Pwv���(�i<M`�I3d���}wEP�E���Ъ�\�;$�3,Y'��X�� PH��[$m�&$��-������hWj�z��񈘤x��@�b�7 �-�rb��WI��F�M�,��{,Y'EB�f��'������hˍ.(<��$�ga�N:�z�i����-d�Z�9vܼ3��,���#�"�I��:�V���^�����빠}�=n(��"�xf�=}& �R��H2K_���31#�<��A8��&�����͒y�l����`�UF�Q0�T}@�*1X�"��пzJK�#4+�� !|o��YWd>!�+�	���)��Q���Oht�M���Q'���� 1S@)���"����A]AX�"U�� E�B�F$�B�ߔF���%@����˺���{)�O�I$�'�UR�f�Y'5�$�{1�'ٙb�>�J8�O�L����h�ʠ*����I�ݱd���b�<���ȢK�k&	�e��s��np���7a�;u��6��؀��D�^N5�T�Bڬ�I?s�}��,���,|8��{��'=���1�O��m��=WqY'����| (�|��A4�"6�m��-����:�V����@�n�^�^F�B@pI	��:�V����rO~�훓� w�ЄX��
 �B���d�;�Mj(�Ȭ����d��PU����O��b�>ǟ�ͷ�����N8��>J�H�^�of�υ��.8�Hv`��"�+���q�u�н6���@9"�s��d����נwr�rD�Ra2�I3@���_�@�����?�VI�ϾvI�fX�O:��6��<�F)3@��Z�ֽ�����s@-�d��PRa"J(�Os�}��,���,Y?T>���_�+$�ϊg�h�`R�JGd�H����%�=}& ?��~���  7M���*�k�f5sn6��D�S�Hg\z�n����<s�Z:�ͺ��㘪���,ݧ����nҽ�t��D
�s5�|�i"�Z��͵��Z�n�u�yh� �g�ͬ�oM�A:�C�vָ�3�#���}��~��<��������r��Nz��6%���jұqJ���۶l��_;�k�<J���ú�U�]�HQ�:&�}��q��#|�ͅ7�H�;p��:MڬP����	�}N5FҗQ�3���@V�͏O�ʐd������rEH:�l!��RE8,��y�� � �W�]�swlY'��X�O�
&�ME��VI��c�O�2ş�B�^�m�$�ߖ��ǜ�A8��&����i'��X�O��+'�*�_�]�{�uX�)�O�I$��빠uv���^�����{�sȉ���R<�n����'X]��]�c:���gI[�����άͤ�$��L�:�V����@�n��u��y;"m)0�%ql��Ͼ��_PD�E�B/@����{ʐ�ʐd��B�}����yW{��rEH� �-���@�e��&�fH�M�h�UH2K@z�L@9"�K��XC!.�N$�b�N��_�_	9���@�u��<���G�p11���l�FI{m�3Z� �+у���x�D�xu헉�[�M�48D<�@�u�@�e4w]���h���'r`�0��@96o`�s$��ɋ�U}�Z=i�nH��L'��$�[?W��r�(`��b���_f���IG�y&�'��h.��l���Δ�y;"m)�%qY'�َ�:(Uݽ<$�M4�ՠ}�,�j6�PJE�iԣ��;�f���U�k�s�.����pf��è�k�dq$�)���h��M��h.��W-x�6�2F�nC@�O`�s$��Ɉ&�~�����ø5i��a��
I!�Nk�VI��W�u���:S@���f(��1���3v��& �:{ꪪ��Z Px ��<�s�]����w �Mɂ��7���h�@�4o>=$��x����;���h���R��^x�/m��c��9I8#g)�l�$��zRv��D�:<�d@s��@9�Z����`�}/h�bx$��NWj�>]kПfL6I����UUA�~�S�D�1)0�%qh���@�e4�b]r�Ɓ?ߖ�z�����O��M��=�̒�~�������� ��.0�m)R4�r$����~ U 3f��'�7]�}��,��*��B��S�H �`7;gK�Ϋn�x���շ]����.4�cg]�սz�\�r��:�h�)攼m6#���Y��W)�5�)N�9��'�1[t[�%K	�J����Q��z��$��8���b�i��mX�O�t�Estv�5X����	,�$ʻq[]���v-�'r��ٻ\P��Y�ݗ����Ł�浵�%ե�BY�A�ɬ�Lܔ֫5'A�8'{����$坛��ێ�a�9v1�O��Y8�]j����3�-�7I=m\����lAHl��y��<^�vI�fX����u�?�����n&��Z�Ɉ$T��O`�s$��}��U}We������0P�F��?[?�=0��UP�=�d���vI燰�0��O�6�4vt��|�Z˭z��;�J�hx�y&�bp�3�1Y'� ��7_	;�4�'��l������rXb1
�%��R�cv���y�9���k����oO[���¨m7-:	(��@�u�@�Қ�:S@�v� ��:��/�a1�R=�Ji���ؔP@����d���}7$�;V���^��r�ǉ��H�iHl��L6Iμ�gE
]Y�쓹����F�B@pI,R�h�& #{:{UӒ�3w3��r-�ֽ�Jh��M�ڴ�Ue"x؅2F���fi`�v�lX3ŷ�M!۱q���ə$��jY34��Gtٻ'r`�0���?ߟ���=�Қ�h.��vu6R) �L������K@zܘ����R�1���I�#X�4�j�>]~����<"0��A@��# �A!$�P�AB�E@A $��; _�1Ez(���vnI���ܒs�m�6����-�ֽ�Jh�za� Ao��I��
E*���YW{����:{���#��Y&H����1�$�ɕ��wG�U�q��Y�G/>�۱/���{��ϙ�8m�d�&���u�?�h.���U���F�B@pI,R��W�
�H�f�N��VI$�!֥���	2!��Z˭z��i�@T��d�d���VI���aN&�	E��d說�T)���+$损vIh.�������ň:p�Z^��Y2FӋ@�gJh�ՠ|�נ^}V��X� �"�؛�ƦamѨ��ĽM�)�&)ڀ[�n�Z���CO @�s��I�#X�4�j�>]k�/>���U�Nh��I�ھ�6�I)QEVI��c�����y��>��M�s�1^�I����&�08%#�O���9�� 'd����1�*C5�mJ���qY?  ^����;纬����d� @-ɚ��w�1�R�I �6Iμ�d�����I�za'�kٹ'�EAU�؊����AU�����DT_􂠪��W�B*
��EU����X*@��
���  �B�*�* *�� *
���ET��@ �D *@`*U��B"� F� 
�EB� P��DE��X
�H
� X
�*�EH
�A`*@����A"*`*`*����QAA��W��*
��PUz"���W�
���T_�"����W���*��EAU��T_T_�����)�����(l�8( ���0���           ��       �  �T��!Q*�B�*(�(
P����
Q@� JH�T���	 �  ��   ��*  Hf�E���g���,�q�^^��Ϧ���(���C��O�ɮ�"�h^� �w�������O�v��<�P��o���냦>�{�(^�=�ٯ�wS��m�^{�W��'�Ux �� $��*�()C6P ���W�׽��n���=j� �t��M��s���� Ε�;��}��� �'����=��( }�wާ��_Zrj��}�+�x xS;�zW��U.MTY[E��< PU@
 F6 {�.3�e\�� m`H� l[fh:v M��	�iF�� � 6 ҉�   ٚR���;( 2��" v � �� ���
t� Q� �@ � 
 �T ��"�� G>�k�w�W�� ]�N[�_m�׳{�t���=)� ܯg9���z���>��yw�|SO�J�u�r�W[��z��i}��{���Yn-϶�M$�w}+� �|D��IP���
��Kc�{�=�ӓS����g ��r���7���U��g�K�|�>��.Ov>��|  ھ}�y�{:5� �S'�>�C�NM.���t� �{��yw�=^v�O&�g>�R�   =!M��J� hS� eT�� E?��4T�� �Ob�Jm�R�  U?�	S�T�J� h ���l�Jji )�'������/�����?�5��w���u��@��C5� Up @UO� 
*�� (��� ��T����?��������!
��u�5�H�$:B CL�-JSP�"��B%�Eb�4aZƁ��ل2f2�CY�����h�$�%� �CA
�i�]K�@� D���DH@�`@�Hu�Y����-4M�ɄQ3W���AG���EEL
�/�n�`3>eYK%�t���5bA��Ɖ�a�ֳp�P4�kQtog#u�Ȝћf��j!��@��m�3zI�P������a��5���L�3[��&���M&L�"he����J�0�hČ�J�3G�^~����޻��0��X�@�D����?~�!'�Y� A#T���c�1 āB$a��c#�y�ɲ�RB�#��Z�q ��%�R�!MW���! ��H\޳������
W�H�|E-zN$��K���]f���[��m��
�)�!FM$J
1�B(!��WR�	��Ѱ�50�h"B��0�R�+n�f]$Zl
�biNɉ��ӆn���T�ҟ'�"Q�GKĪ8���ф�^HQ��B�I�$C�*JX�hĀ��m��B5��Ѕ.�˭��T�2���}϶�
B0#!��!P֍r�g�H�'��2M�@�,jD)
aB$�c5x}�f���� �X@�1�Ʋ��Z������4���X�Z��V֘�t@(i���D���8����}��־e4B "���$V&�}��Z�
D��0*��>�D�E�T4���?m 4l��6�x��)�� l�����HF��!3sqN?�0`B�p��s�g�$+�7�䌒�WLClx�(kp��u����*D�!!7XHGo5�0�H$w9����9�?�bos��#l�G��7y�?1hhɸ����t�n�WXϹ P8�F+%�Z�������8@6JI)��d#SA��)���b$I �`nN"��<4��8h��g� �X�6��U��"E0H%�H�F � ,�]i:�l?�?����c��D*&�$P #�A�?*EJ�q6!�\]��bAk���j@���a�|�O�]bkg��"44㳇��ц��?��:q۷�����)t���ߍ�%͘c��d��If�a����.�P�`O��ą�X�!B$*h�0ڲ�L��*F	�^��Ѩ[����$�+�/�B�n�$�����-�,
��
��X��f�e���rn��n_��Q�A�������1L# 6g~Ϸ2+������߂@���&�]c2�͒��8���A���B��4����H�bSI����H��FSZ����$H?��R_�͇>m۔���$�XhH�I��71�XΈ!C���O��������Ec����p��#1�
1 @F��bĤ@�A�(E���D�� S�Sf����h�/��?0ы�P���Hl8~�oG�Y���o�����p`Gg�]@�,)f�3F���vA�$���3��o`1�s_��n���FS\e�2�I!tc��P5���n�x��ĉЂ�ae?s���~�B�_r��p��h�Ku�ow�s�х����ħ�#�@�$"A?+�āMf͝@��Y���ђ����!���1c0�H�Ɯ�M`l(*M0�0,n�J��!��(F�Ra�;�!.��.���!M�,c�o���.�A#�K
�#ZjL�-������y�����rB-Ng���������35���V\�N�4����4/$R"tf��^Z�b��gSJ�,1
�B���5�Zj@j��ѹJ�/��)�|ֻ5��2t�����X��T�ea`$�D �l�2�1�3R�B��_����.��	���%4�°���#+(J��C���,�&ka���ޠD�5�i$+��7�٭��C+�"T����3DH�����kW!��	�Y����X$"f=�j���g�$�?]L᱒<!]�,,����
�J1J�#�DB"��U��{=�qٯ;����k;�^�%5�HB]�?k7�5�̟��Mf��74a�:���?d"�F-4a��BJi�� Ņ� VY�Mkf�6�K����!�
k]�'��`m�h��Z� �xJ���Ytļ#u.oV�"kC�?!��B@�A��+ �������n�X� L�~����	!�O��ī�~bB��E�bB�h��Yw��&����˛������k9��^M�s���[�u�
H���/8Ye���j�6;#2%M��7�ٲ2Pф7����7?k7x�߇�0�,�lW�(�����G��;t|t�3��˰☟"mH�BT!��6d��Ą����O��C�Bi�6P� �H���D���c�F^98m$��oe�L�71(�Z���E ;Hac��06�Lv,��ad©B;��JI���H쐉!(kS@�����F!F�7�rM��Y5�%��f��|F���q����I4L98�mٲ1�SN8��`M8ZKK�4`�X4t�)�ٿ����B����g��8���q��!����?$B��o7hi�b�!�I�� V�n~͘q�qv��H8�#�%pq۱0!�N8oq�l�Į��/	��٧����ۜ7(b�(C�!�"@��ٲ��4�) �6`q"SFÉ��٣�Ԍ#dю͒��L��M i�"P˸]����h��`mLaI �Ƹ�(�͡�;ջ>��ʒ�cl�u,u+-lH���1�@�cH0,�(0d% ��BB,ClB��~$��\7)�0�6�b&���_�5�g�i�6��2���m �5H�A��n����b @�
�@�1Z�F�W���l�%!e��m�@��#E��ҏ�E� ��
��%g
jSa@���B�j@`&�$^��!�&�a��ַ�H�b��pM0$����s�+�@ٴ�]�5�0�a�������%�3Fmv�F����m٩e�3�6R2+�c-���H	,�@b��_�K!��g9�$,
���a
,hŉ,� �B��C���"H$�e
��c�	��4�HA�d$,$u��nx8�xr\ٸ�Q�X��0ѨU)�i�����#ta�h�t��o"]`CFCa
i!]'E@d�_d:�?}��Z)������l���D�X'�#G���PИ�A�21/�~��@              ��                                    � �                    � �            �A�                            �     l              [@6�  h�Í�`�d�pvY&U� �  ���ڐ  H 8 -�խ�i �Wafr�l� �YV�]��vٲ�u��m�   � �[@ �`��D�i�>��[BY����X��-�9P����VX6���ڀ���f�x�k6���j��U]��Xs�*�VV�u/]T��@���V�����e�r鱵���W`�$m� 	m��x�[p[@ [U� uK�R����*��p'=-<�*0[uL����6ڀU�j���l4צ�f�:F�  � m�m'2���m��`  ���w���  �[NsZͶ�^ �8�]dw/$k��ƘL��b��0�[T]Uqd�We@6e[I�mi��l6	mČ  4��Tյ$v6�M��-��5��-j�X�Il��&m�)  v�f�e'f�	�( 	���aF����N�&A�S�t Ġ�8�UK�*\둵-UR�P!��� �UUʷ�E����Hn�]��b���8$\�  �����wg�ys���]�si6 ����`v�U��+�NJ�C]kl�l��P�ō�a$������m��H��m6kv�H� 3l�;o25�$�-�e�v�\��mHW)m�h-�m�@m� U;�Gv@y���uV�Um��`K/� ��E�ڶ  ���m�	 mM�]�ӧ����А-4�� ��P�I���m�:�9���n� p$ 8��,����k,��vَ
ڪ�U��$��6I�m��V���h�R���H�#L��*��J�8yV�6�U�	�,-�	 ݮ�-�������xW�<�W]�ګ�d��t�4�l��M�-��km���   �h�L 	+�A6!!�8`����. =�䞆�m�m� ���tЉ0 9:H�m����z���fXD�RP⪪              h�I� ��  n�H��l-��V���6�88�5��l%�� lh+LIۀj�m�l6�i�JWvm���^��u-\ H��lJ�6�Kۃ�m��T����/Q��&ݤ� �[����M<�8  �uE6$	�-�s�U�ck��m &�	;m��z����[� uR�!�G=�aBUں���輴�z���m���-�ڐ۶[[lź�nѴNe�@6؃qm�^�#&��p�`��'�[/Ut��`-G��m�`  $Hpt֮l$$�[v�pn�  K)�V�q��֤ VV�@;� \�@4u��lm�&��GH[V�GA�6����5�m�-��vm��ާi5�%�� �$�]��!���88��l�V-�,���T[�-��si�`�Ml��-�R-���CX�@m�In��m�܋Xq!�	 	 6� 8u++Uv1���sJ�Pq���&  �.�  �H��Ŧ�6l p�M�jN i2�� H  ۶ŵi�u��a���V�U+̪�*�Q*��F[N ��   [F�8 $�7m�V�  ^���sz�t���I��L  m�      -��O@�m���D��À H        M+i6�
�}澨    ���i ��S-��� �	m� m���   �oDw�۪�ÆT(���Ί � 3k�Ԏm��     �b�[@ �H    ͷ6�my9:�p@ �kD��d`%>;Zw�m���^���[A�zJ[\v�X%T���FH,�wNQ�M3�Y%� �˰    K(�HIm [@p[Iem�v�$     2m�I���כ       �f�n�"EK7,UU]J�+���� �`�,�6�m� �m�ioT�d�t��dͶ� S,UT�/�n�`cYv�  �a���mzݎ���@��f6 @l�'lȬb�{v	�O�w8� h �  �  nݧL�`lt�#r�(e�����	�/��d8   �oPmH �i�l$� VǾ�%���N��uc��u�8)V�T�@�ba �kh� �  m�m@        6�-�  ��} :l��� �mm� ڶ�4���f��k`�ӌ�I$l崶��  $ݶ   �  �cm���O�m im]Բ\ &ٶ�` �ֶ�m�-�!mm�L��t�l�&�Am��l�I m�F�m���m���8 j�`�c�ezꀥ���\�K��3d���bޤ��m��z����fV��[� ��I�h �I%/m�G^�.�p ꪁ 
�������    $ $ H6��d[��[����k�H[Bں�6�����ζ�e��   �m�m�%�  b����뛧�n�E�j�8+��ͲK3�Iʹ�-UUUp�N��ۈ���1WJ����r�5m&�;k{�d��[@n��	v��'Y��U��$ �[p �c]�p`�ћ`  H5� ����ٶ$ C�tݧIr�� p$UF���a��	�l m�6�c��K�m&H n�.Km�	6P2�m�++UUP���q��    m�I4���{M��v    �^����z�,��6��[�Ò� �n�nÀ   � 	6��hi��m��-� A��$  �3     �d� l�i�褁Ā    	 ���  n�f� ��
��V��b�aY��%� �3��8�����8�hm�����p5��z�mr��eenVU�e��� �l�v��hz��m��z�`'��@l��@�۶/]�[l sm�#�l�` 8[m�e�lpv�^�m&ֵ�  �v� �$ev����*�۠����  �nkm���g^�2�U��(��  �&� $$��|�g���)V�A�பꡛl��8$z��e�UUU!��yB�YVEF�� m&�[I,T�],P:4+!5U�]&�|V�ڱ[��4Z ���Hzմ	e�mkl����������J�,���m� [^.�m2\��Iҗ`�p    kC`ͷ^�-6ۋ�Z ����&�[\  �
U�����U'���� e=5�� q�ȷ�"@<�"jB��P�K�/At��ی�5l�U] �᪠*��_Ӯ��(v��m� $5�� �V�   � �    =A&�[�    6�ݤ�l  ��`���lm�Ե��Ā �m�t��h /Z �mjٶ��K�]6݉[@ �ki;` �Pm�m���*���(/]2l�l9j�l���<�	�)-+�l8     pp��l��N��   md���m��h�+�m*ܗK�l�  ��m��kdkh�   �  ;i+i �nYB�[AJ �����U��R�N���1�=>W���QV�����Fh��z!�+f�e��  햁�m  -��������� H���}�-��m&�m�� ��       H�HՆ�  ��  	$�޸ H�q�`     r@  �6�V   �PHi3l  8 6� ��  �  m�    �6@h�U��m8m������mI�l��6ͻ]������ �3�� $-��ӳY9��x2sK'\��� NRte�$8Ͷ�z���&[I��m���[@e����	 N��m�k��L��n݀mf��Y!�p�m� ��I�m�x-���I3mmd0p����  mږ� �[{l ����m @����ŶJJ�jj��G)+mUp�Cm�x��wwy��y�w�����®�W�� ���|���(�
��D�(��C�� �+ �$X �(�� $1�+ -~U^< ��S ؉�� D@�^(�"#�)��������j�% �� ����U������R"��Q6
���"^
��`���| ~G� _�$�Y"u�"�����_�UC���@D���E�	c,�$Q�!�?.�zP�A@�����D8tv��Z" '�� � �B����4s�� ��#�E�� ��PB�XA��Q��P:��j,W@�`�UlQ�b� ,���Z"��$X��A��C E ���D�@�U.��%#6��/���@_ȁ�~�(tN� 
*�Q�q_� �"TX��I�3]���� 6�      M��`  �@ ��    @  B�����&�v֜�ld�ꩲңUTj�\�V6V���Q"ܰ��6�+�p�	�*��U[U�6[pW]�1ԸȈ��I;�p,�b���m�Ċd�t�<*�om�X͡X�3��S���EJrS�X��R^�����,�u�3�rnJC�+�12�Q�c,n�mu�N�ъe۷2�Y�Z��Okj�ѻRg� 
��Ԁ  ;m��4�V�e� �V.yG�h���+ɨ�m�����b;0�0.E�J\Lo&-k]s���`���*�.���-�.���,zy(�8@mm��x�U��sjz9����*fg��<%�J���,Qʍ�T��ͳE �,�l�`�S���5��KN4ʩ=��҃��U���n8B^z���E�Þ�z�UV�<���Z������;>D��1J�`6�n6ֻX]
q�s����ڦ\��v[�y�I�KX�ݗ��m����m�̃l�\�5���i!��������ۙ6�5%��9�΍%N��b#M�4�P������2k'6��J&�T_]��LOH{\tv̭�&˫�;V�njT����q���3��uO���c:�KJ�R�!�6
j��4�*��/
�]�:���šn�zd޻tL����]ۭ��Xۼ�0��N���;�k-uX�g:k��J��pn;4M�Gd���Q;:��*�аy�,�J���n޻e8��3�ԭ��*�UR��F��:6k�R����ib'e8�5��=����ź��)< r�ĕ[K��<A���݋R�u�͵�Nl�^���-�d�.�l�*�lЎ1K� sR��mU�JAv������FH=rg��xz�d8H����Ԫۖ���+���\���DY�\����h����>UW��b� S��D�8� mT�|����'�~����!7X�ӕv%r�pS켌����b�f���EnwI	��f���ј�mG<hn jUM�+�Ў�
m���ų��)m�I�I����֓�2dl�UC�����u�;Og�M�qX���X�YDw���3]�<\��k92DP�<ΎI�k��ގNziN�y�D2+�Y�e���ܐT�zP׻�����{�V��Epa�vs�v�.ܛ���q�<`�v�dxݰ�`@�p�^U�^��Uw^���`�j��v��13 5����R�Uv�u
����蘙�F��0y��^���Q�Jc���Ɣ�Š~���^�@��W�[�ՠr�f89��&H�R��h^��z:�;?�?��{��u�c��M�#�"�Wx.r�	�X��`G/ ??v�o?��k��<D��y���;��P����ӓE��]��JA����q�H�z:�޲���h^��T��s"b#i��@��)�����HB �X 	�bb��d��D�o��<������<�E#�ѱȆ��f���@���@��)�{���ʉ0Shn94/uz�Z�YM ��4�á���H�&�z�Z��{�̳ :9x.r�Q�IK�8��JDx�s���'kt:��A��0������,k������ө����oK� tr�\�`;�����AH�$j) ��4/uz�Z�YMY���ؑ�݌��%$#��Wuw�y{]`��X\MDL��19���3�E�)�m�ִ��q�8�q�H�z:�޲���h^��T��s"b#i��@��)��f���@���@�1^��5�����vy��8�c	/�K��Л`�D��ŵ>�w{��V�r^�4e�@����9X��,z\0uY�,�)�DF��@��W�[�ՠoK� tr��ϒ���v�u�UwX��,z\0_}��䎎^˝z^(ޥ!#�)�@��)�I��w7$�}�nO�	�t���� u�{5��'���ə���$j) ��4/uz�Z�v��ffV�$�8�P\\XE\��K=;�#mt�����2���'/���9�at���y�wso}h���)��'��������5�}�l�1? 7�^ >�J���lq�����uh�e4׬�<����,vF9�i��qŠoK� tr�\�`;��ey�)18�n3�3��4��h�uh���=�E��UB��EU���Z��=�+��{�����~�nI�W�!�Y���"F"EB�+WH�hj���lA��4��6�5�X��� l �aۧi����k�rJ�Gs+I���d������v��� �4䵩�1ɓ���;i%��\a�m���a=���u��rM�ۤ�v�'��gv�
��\����/	I�p�]PlJ[m���XX,���ԩ��<Tjݔ-�.ren����$N��ѣ���J�*!��q[ҝp��l����	#�_8�#��m��VC[g%�����x6�B��v�un#��$r���(W<nY嵶���Y��Z9tk�WŲ���A��Q�������6K� tr����uq`2X��t]�ut��U����&f% �}x���z:�+l�	 �qI�5j���^ �8�	�X�p�:۱�)0$�<�)�s�z:���h,Ľz� ������rD�Z�Z�e4׬�;�U�}����c�sȇ��"It��.���a�n=�0m.����L%�Z�@^�G0�"6�N8�ﾟ��hϪ�-���/:�I�����Cp�I��w7�� �b*��kۻ�}��@�l���uQbWB����&����ގ������hx�%&
���.�j��L�DB�y\�}���^�@�}V�ת��%22BGR7���M��現�OkoGV���IO���'L�ژ�I�����q֫R�':2�P��st� f�,Z��	 ��I�5��z��s�z:���hm�Ȕ�H�I�]���gD�DL$w;�Xuw, ��4�$��q�8�ܑ7�oG۹'{���hA((�)�C��s�l�-}V����dc�F�M'Z�ՠ�f�k�h�uh��H���dlrcR- ��4]�@���@�ڴz��D�JL)n�6j�{8����b���M՗7m�]",�QbGB����&�k�h�uh�V�z�����J�y$H�I�oGV�k�h�Y�Z�_>���w�������V�B�>m����h�Y�Z�Z�Z��c��RH��#�C�K��M��-ݺkLDz6b"j&&"/]���)ZR`I"y$R94��h�uh���^�@��J�q9��1�9?��y���x�E�X�,i�g�a2A�n��8i6n��\�S#r68�ܑ7�>����?[)��f��������27���ӕk ��f~���y����7�M`r]H���dlr!�h�Y�w>�@���@�l���,B��Q�����;�U�[�ՠ~�S@=z���E���H�"�-ގ������ְ����"��  m� �����z�+��vupZ7b�;a�6ܗ�Ji�2�9.�#;6��N�-�RMy�a��gn
���͎^�n��2�v|v�m`ۜn�n��z�+��k�|��un:��*�K[Y����.�yv�����n�]���S��Q�;q�Q0X��������(�3A����;�,���v��f��gBt��8gR:�x�|����O�����غBt���������]�R�i�6�h�&�^�d�2��aG��X�ѫSR7�����@=z���Z�Z��c��RH���C@=z���Z�Z�e5$u��Q)0$�<�)�s�z:��ffb_|��h}~���V�rF��&��$wQ`T� :9x�"��c�1̍�"i��@�ڴ�?�������X{t� �iT�$�
���q�N�Iֹ4r>Pm����"��E�$&qd�[Ѻ5�S�Yͦ;R�$�?>M�j�-���-v��TX��ɚ�53Z��k3rN�]��b� �X�S(on���� y��թJ�y$H�I�oGV�k�h�Y�Z�Z�^7��&HH�JF��-v� ��4]�@���@��p�
I��qh�Y�}����u�/��w\�鵀tDD�ǻ��K�act���s.��z;m��0��p��IYx���Ԭ΂j]3Xt�w
c�uw,��k n�X���I;#hq��"n-ގ��33?�>������4]�@�yc�1̍�"i��@�ڴ޶i칙���1�dD"��큀�Cj�T.��: <��,WD�J� &�~�]beTց�J)HU띨B�([!RFe�0.��C����ȉS�	XԀ�H���!BAP�dd�I
���UFČ`]o�أ��]�SG�H��C�!�(�X�$_�Q�)���l<��8�U������r���5�)l���ˬ5�i���a��w'A��wٹ'��z�Qyd�;�X}30�uw,Y]Q]e�WEަyw�f�O{^�ߕ�ｚ��� [�k޻�O�����'���Y����e�˱$�mmj|��\�6�m�R2�cv��7'AX�	#�l=Pi4T~����]~X��ܾ �}xt��]��>���yHթ�e��o�_�O���鄃u���ܰ�k:5wu�YW�E&8�Z�~��ՠ_tui�K��-���`I"y$QI4鵀?m�Xt���ٙ���LN��M*�F�Q�*?������䕰�1c�r&��/�:�e������,��I����K�^��ㄪv(]�uq�W`,O[�R::n;La�9bA���9#��"&�n8��j�{��-v��GV�W���FF�&5"�z٠Z�Z�j�=èŖE��$nM�j���XGu�/�7{�:ba#_+R�E�$]"�ݬ艘��|uw,:b"R7{� ���3�o�*�Z�h�.��+��XLD.��X��}���X.o+� DD�Ǜ뻿���]����U�z�c(�8�U��S�y^���u�y����ƃe���gF�1ؕwI��.�/:�:R�ᓗhp\�a�ni���t
h�5g���fkF�,�/kfN�T��!�&����m� Ү�$]�]�'^6�kDi�eΤ�\�iȜ�ۗvG��iL�:�tg��1�G�lM�1{#As�� �]خ���H�g������|�+�%χ]slu0��q`�۝�n�g�`
��X���mz�;55
vde��O�??^�>Wj�/tuh�V��׮4I�$��E$�-v��GV�k�h�l�ܒ�F,q��"n-�GV�k�h�l�-v����dc��D�c�-�j�z٠Z�Z�R'1����LjE���@�ڴ�Z�ՠZ鈹<q-t*7�[��:�r������D�>��a4�Pe݇cq�JS�Z��n�Xݺk n�_Ș����׀k�E��}���"�-�GV�ff<�$b+",��\��k޻�N��p-v��?���#�~xި����Ɠ�ŀwWr�{]��k o^Y�y7f8ԍI"�p�- �z��j�-��-v����$��D��E$�-v�޻�j�׬�'�ܖߒy�tv-t�s�%q�_)nS����9y�n)����np]p§38V��T�f��qh��h�V�~�f�k�hW�;#�M����-v� �z��j�-��*�u"s����ƤZ����ե����}�3&f.&"~��K�,����}��!C��Q�#$�ɠZ�Z�v�ՠ~W��=�E��\O&H(��h��0�����_�ϫ n�X���ڄ�ݛB�R9D�:E&���-���t��:����[�;�/,BF�L�NHh�V��^�@�ڴz�4+l���!$�#�@��W�Z�Z�v�ՠwr��D�H�9"R=�j�-��-v��^�~䕰r6��&��;�.t��>O]`l��LTL��Ż���^X�s#x��bRa�Z�Z�z��j�;�.�Q��<S���A�q���kd��r��y�wnT^�Tb�,���m��(���?ߵ�IR,�� ��X�L<�.�j6�dq��]�@�t�h�V��^�@�X���y2AF���@�t�h�V��^�@�ڴ�^7�&�)�hq�4]�@��W�Z�Z{��@��ƤjH90�Šj�V%H���J�`�8 0 �ÔV�lpZ�v;3i�-����Ҝ��7n�[s�s�-h��%l��u�u
Ӷ�N�Z:��ۃo$ln6�w)��v�v��΍���k�vwc���v�mp�a�k��ƛe*3/�ɪm���6�9�1���o)�Okt[$�F��N���'j�r�jCS:�2�f�+�x��w�k�q�oe�+���G8������"~{�����������ٻu��Gh*I��];d#�^ܕ���e'g^��{�f�5�;[LY�@�wi]��~�_�,}���>n���Py}~z�I}`�m8'$MŠw�83�"&=�|`\���ְ'���dolJL4��h��hϪ�;�.\.�Nbp269Uf lr��ŀ>w<`w���]&��� ���v�~�$�:��� ���[�$���X�Kd�n����x�Kd�l�g��$Αb��6r��\{��x��v�O1Ht3���U�`�Oc�=t�Mv�RI���$�ɐ�I#���$��_������~��K��ə�> ^w���#�TZ~ǃ�Y��Lݶ�ݗ���IwIq-�g��6�n�G�� ��5���$z�MI%�:�ߗ�ۮϱ�I%�ߏߒK�+�D8�'�B+��$�v��I'N�bI-�!���������������l��U�P���N��RĒ[&Cu$��ĒMۇ��������r�R�-s�XK�l��F�3s�y�u�h��S	x�����������F�6�I�~I%�v��$��)1$�v��I'N�bI)M'W~��E�V�U�|�G���&f��n�/�I*��Ԓ_��~��^��"�FԔ]�U��$���I:w=K{�{���3ĕ^y���<헉$���)4T_��t�Wv�RWﾦ�'�Ē]&Cu$�YI�$��U��IW��z�2b���"�Ա$�ɐ�I#���$�v��I.}.5�$�Z	-��b�8�d����*�:6�A7ZV��N�5Ӑ��sujLp�6S&jf%: O��m�#�m�����I'N�bI-�!��N��Wh�I��E!5$�t�~�٘�\�\kIt�Ԓ:\/I(�RYV����ʮ�UZ�I'N�bI-�!��GK�Ԓ]Ӫ��$�����i�"����X�Kd�n����x�I�qn����!f2�P(�"1  HA#$`��ү�(�h @���;ة�*gsY��ݶ�ϒ�E&7����p��$�YI�$��o*-Ԓt�z�$��2�%��R�Ѱ�c&!���;=9`��1D:�նӛ��0���c�$��T�^$�n�[�$���,I%�d7RH�p�I%����Ez�t+�Z����N����333UI{�8��7��Ē[��}�$���=2"BG$sԒ_��}�Iv�ĺ}wm�r��t$���:89r
L!$���$z�MI%�z��$��ۊX�興���w�}�I:k�r!�$�<ndRRIwN������$���g�$��l�K'�,���%@�%R%
�
�� ����t��Bg�IUӦR(P.�@8��!�2K3J:�E��H�0 D��� Q����O�r����0�hAYsbA��ӌ�Z����8B��7��E�F*B��
���0ִе�J�p�a� Čc!5j��4�!%�R!HU�44D.���D�<u_���c CB'���c1 �u#@�ŀ@ F�b�cӈ�i�#�H f�.�� !D^$M�Z*��H�0��� A� ��2E�'�t��?~�}          $��6ހ  6�`       @h  HSU0����nۭgZ��H��UUF����me˲q9��knA�]{=J�a3@�mEq�8n�@�
��l�;�v��R� ��p��d�2�2Ȃܦ3m3�p��F�V����v��eI�wIV����P�K�+�4#�d'�+�rDȸ.
�[�X":s��l��8!����8B�)'nʓ%���W/.e�ۋ�&����gH5`��L�%�M��\M��Km�  [��Fĭ.�&�Q%z�Ǉ8zv�T��(A ���>אsF[E ���Usn$��#u��8��i�ZP��z����t�]n:�ĥ#��i��D��R��ضNh��	�l�(U)����M�-�dp��m�9e��V�U�l��: 	zm���l�F�^VVq�^T8ی��-U���hw����6�s��q-�V�]���ut�m ��q���yׯ����G;ny	��ŮL��t�ܚ���[n�
M�{7���x�;x�vj��U�U�	vZ��pCN�8*�Y�'ӁRݻ{�[8��E�g���v4A��8P|���vs�TR=�pT�J��V�a���Xݹ�+�r�
���&b�7����4�dJː��*]S6�L��XI���i���}��I��6��MU�L�.�e9��N�UB�n]v�&敳=���D�:�죰���(٘*�w9g�Xq�5�����ۑ�>���<��l��֧/F�n���獶��|����q��<Yrv�۠�Rɛl�{���dݰ lQP���ܷDk��xs�vD�&\5��i#6%��u�F���uؔ�p�\PJE����P�s���f^Wd���UP��TCb��k�����F �U�X
��Yö�#�1n�q�a1ֶ�s7g��9�o���!�ŗ{Gf��(�AF䠥\3.9)K�Zd ��� h8���Gh<C�ڂ'�|�������ϗ��  6��jw������d��Y��V�ٸ�hKv�絜 ���$rr-v�ꆎX�������]�;�{ff�]n8��nկm$b��K���c���\�Dm^�]<�E�z��
=�,;
)�No
��ٺQ�g��M8B�ungn������@�+��HCvY��u�-V8�f�FF	�G����v�:خ����vy��\�����{(\�Wi�-�wϟ>k��n�ƭ�8�:�8݈�9��
^Z�՚��U���<NH���IU���$�[���$���jI.��~��B���r6�E'�Ē[&Cu$�K��$�v��I&�������E&7����p��$���X�Kv���_�"j��}bI/wg|�^��"�FԌ�7"Ԓ]Ӫ��$ӹ�$�ɐ�I%��I%�i�,�y21F��H�~I.].RI~�i��K��X�I�qn��L��tW��]!8�#�N:�i�v��e��v�F{Um�h�2��0���5jd�ݟ�ɐ�I%��I$ݸ�RI�s�bI/>����G ��H~��K�X���@"$	�Hf���;��[o���RI~�i����͵[���C�I"x�ڻ��$����RI�s�bI-�!��K�X�$����(�A9"n/ߒKVۂ�$���>�$���X�虘�o?~�����s���s�]��� ?$�n�#���$�v��I'N�bI/�����@�7^���v�\�Ș��������������HBK��ZE,�8ҪҪ�u$��ĒMۋu$�;����w��}����� �~����%��-��$���I:w=KIl�Ԓ:gfo�*kZ���z�z�f��Y����[ou��m��w��_�QCjeɝΓRIw�U��IW��f��mne,I%�d7RH�p�I$ݸ�RS�> ?�����f��WkUo���YV�K���Ԓi��X�Kd�n��R��Q��;>�s.��tvۭ�a�#�����<soj%X��T�i%�"6�Z.�bI&�ź�GT�W�$�L��I'��c� ~������6�����=�I-�!��I���$�v��I!^X�Ĝ���7�L�jI/��?~I$��X�I�qn���=�I)LC���U���vn��n�I$ݸ�RH꞊�%�{�{�Kd�n������.�%)�- ���~�����K�	l�ԒMܵ�$���'�/D$���n��Q:�k�ks�ۣBm�[d2�
�˶F��j/c�=t�MqQ������$�ɐ�I$��X�I�qn��MB���DHH�D��jI/��?~�?�i[>�RI[/��䒫��Ԓ^}j��(Zt@�_V�?�m���ϗ��Ԫ�)5$��v��$�n�\�(�Iz��]�ĒMۋu$�wQ^$��2�$�t�jI%N�l$Q�$x��7�IDI%�d7RI7r�$�n�?? ;�������w�}�}����`*���_b9ؕ��&A�L�p=$枌u�Ͷ���vc[1���ۚ���	�F�幔s&�5���oc��m�����wQ�>�p/�:�k<l�"��L�6�Ր�<Q�at�\������r�Fsl�N��0k(U�H�q�
�L�]�t�ݿ��Ϙs�|�ڽ�{)�]���'�n��&�Y�!�b��	��m�<���{��9��I�]մ�i���)QR�mvN$Zݪ�Б͓��s�$E9���Ή\�_�������?%�n�$�ݽk���{Ԓ��^$��b�ի�tU�>�$��Y�35T�v�}�Irw\� ��f�U�(r(�mH�#p�;�U�r�h���=�)�~�]�,�y21F��H��Ix�p�9�� �8�[*��dD��Dd�ɠ~�S@�t������կ@��6��c�/�ɓ�Wga�v�`���j膹�PPљd�r�n����c��I"Ra	$4wJhϪ�;�Z���h�n�Q�'�ݫ� ݭkL��)���C�V� ��f��ft�D�AÅ�eں�]�.��qh���~�S@�t����� ��;&7$ldQ�ґ����=�l�7kZ�鈄��u`����XU�]�T%v`ݶ`:������ ��S@/S`��<Q�� <s����)4�S��x9�vT�ϡ�&�� v��yhv9�5R2H�4s��V��YM�Қ�k���&F(�1I�ޤ�gL��G�_�|`�ְ��<��$$j#N=�YM�Қ<����;1�o��9r�h]j��$RH��G#�@�t���ڴ�V�7��w�߷ߧͷ���}h�5P��[ r�X�RV �H�n���o?����˺��.�q�o)�\˃8��#/G&��\0��ܙmp֢{��Zy�^��ڴwJh]�@-8vLn8؈�m�#�:�V���M��h�z\#�#��FF��$Z��4�ՠ{�*��ՠ{�@X�#Q�#$��C������W��]�>�r��I�u���*��O���{8�7�t�9
�]"�]��=�i�]6����m`1>��C��n��.fŔEe�F٬u����R�V��7;�k�s��+N4��]CU��V��w,�;f��X�m5�{�O�E$���N-�����ڴwEV��ڴ^櫑8�I"�U]�� i�X7j,eH��p��
�H��H�N(�z���@�R,z\0�����߮�]�uEU+Xʑ`��4ܬ�?��I��|� 0 Bn�h����5ձ�c�^O�t�E����i��G;]n��E�����L�Jv	x��tQ ��T����
a�F�mnyk7J�[m9��-i�Iq��N���Ke�P��RY�:��=
��qeN�mt����&'nYG'O(�[jf�\qs��=O�_�����L��vۇo=Y�7�D���e�6�8�nJ�}�>�}���ߕ���p�x����$�9(Sp�l���ܩ�����iE�M8�,�5jcdD�p�)�r�@�tUh�ՠ{�@X�#Q�#$��@��X7j,uH��p�9ҟ�&)�4L�Ǡ{�*��j�?z�hwW�����L����8��'T� ޗ&�`ݨ��'�I"�AI�N'���S@���۶�����~����oK�����7mvSARON��َѺ�GQ#(\�������̮��Ut���yh��m�����sv��:;��.�]��L�kYu�.�[�~�콻�)�B/�����UK� ��]%`��rL�8�Ej-�ڴ޲�]���ս�"�G� ؘ+� ����t�V��0�PYq��d��h�k�=ϕz�Jh�e4���U2H��`�"��-���Y|�����n��=j+E���ӯ+�d�i�"LSh�#�@�>���l�=�l�����͊��\�5�#z�Jh���9zנ{�V������I ����߻���}w��ٴG�}� u�D�e���X���"Q�cd�M�Hlp?0_�� �F�Db�&f�1�Hȉ?�TKaqx������Xb�@�a!, �B���@a�2p�AV �I𫠿
��C��@`��T���D�!QW���] �j�=@֕ m\@?"�V����k?k�5��>��ٸ�̲D�1Ix܊C@��^��|��=zS@��)�����0�G�'��|��=zS@��)�r��~m����������~�i�`�g�Z�V��W�����E]��Ś�Ղ���K$��DQ���}gƁ��V��ֽ����"�G� ؘ)f��X]%`T�XGp�5�c�#q�##IŠr��@��o@��ʑ`ԟ��Ez����뺺�5�uX��0�6�>������-z�8O.)��	"$���!�l� �IX�%V���y�7*�E��F��Q��7"�WXӒ#$v�k�r���i�j��영)�.�*E�5�V �IU�tw�:$�8�RF�6���9zנuv��z�����V�^B�(Ȝ�)n� r���:;���X]%`�n�"q���r7��b��h����9zנuv��UDZ8���P+� ��k �u������ �~���6�|���ňHE �����o��s33333&c  l;B�WP�Y��x��mъ�e�y��2��^:�ZM���LěHf����6v�tooF�]l��-�:�珛|~[6�ivb����A�5�ˉ����e'�6 �éNK&ݪyR��7��<Fɵ����۷U�6�s]�8.�n�4��(�vkq��N�\X�z�+�b��B���YV�FB6u8쉻p&Gb-?�w{������?2���a�g����f�X<<��M��՗V�Mef����Բ��>m����k ����tw��X�'�^��(�2G�Ws�@��M�v���z�O.)��	&Hܚ��`�"��+ ����?t%z��H)0�4yڴ^��w;4^��/:�!F)#Ocqht��D�K�:;��R,I~?]���7$��/��q�v�{�;�M�݌�0Z��l[�9�����mu�����m��M�W�� ��w$�$i6�Q�4^�ٟ����?�'�fc0�ŀyou`nӼ э�8�1������;V��ֽ��f��Қ�b;�7R24�X�t�`D�K�;���6��S�YP�b��D�z]��ץ4yڴ^����.UL`�)��N����'S����:��A��ۛ�X�r�r�y�)�4L��4^��=�j�9zנU���;=J�c�I ��Uf�R,�q`7R���^u��H�)#OcqhϪН�}���(iM$H��@b�3����h�+a"���"�9-`7R����^ �8�g7rL���q��Q94��hz٠w>�@��Y�Z�mQ�����f8;a.b�x&hp�pr��[ҳ�q�k��le���D��bSi�Hhz٠w>�@��Y�~�S@�T��5R�R���q`4��%� I4�;��P�b��D�R-�]f��\0���7N, ��*��֋��qv���{�8��׀nֵ��b0����y�َ�Sf���W�G"�A]�Uf >���ŀGI��6IM�6��&'��LA(��I�tvۨ���a.��c�H�K�����&!��x�iɠw>�@��W�~�S@;�� ��UܑFD�A7�y�+ �. �K�� luS�~�nb$�H�N=���޶hϪ�/5��p���bQi�Hh�E�7N,:NV�\0"�Y\Q
26F��@�}V�W.�@�]�ܓ���n������ffff �  .�uX�k{4��GI�M�:4u���gm׊S<��F-�l��5c�]��.�jW�jMͻv�c�=[�;[�~u����+F9��k���n�m�m��gLj䋴�^����C.��:��UT���p�z�;qt�v�s狍Z�^�'l��bRZ2�3֧f;cU�+<���\qsdM՘����3ɹ��
�D��3KF�N��aXQ��w{7� �%c.���{]��^�pp���]���.�v]�Wd�[���}����Ě�Q�m��/߯ n�X��Xt��6B�
a2BF��7&���M�g�Gs��Z��@��ٿ�$v_��=�I&jE�w?�Z�ՠuuW�Z�Zs�tr<RF�6����?�}���>���m`tL/u�, �4%�]c�I�n-����j�?Wj�-v�����_f?��!A�1cZ0<��$��Y6ڵ�E����n�.ră_��3oxA�Vb��ܓ��_d�_7ϗ n�]1��˫ ��>*��+Df���k2nI���n���(����w���u�� ۶gDL�F��WYt(��N-��-����)�}�l�=��CEE¸���)]��������;���>�`tL�B��y����L���D�=�)��""#����wWr�=��� պU$�/Fz�u�F��p���@st�Z�]�F�:X��&���7:�ww�۷�����	N���;���ՠ{�V�l���}��BG�H���R�տfg�$k��Xw_���33	��.踞89$PMŠuw��l��3�?�����MDDD������� ku� 7��I	#J(�G#zff/����;z���u��"bbV�}U�r䃸����uT��� ��� �3��W�uw���)��"ǈx�G!&�x�U-k��cr�{p��b�aI��\��VWq�������{�ǰ�Q��H�?���}[�-���e4q�*"��.��mju��"b?DDDEQ���Ɓ��?ƁWuz�w�2d��".�� ���v�:f""��V����;=J���RH)0�fLB��q�ro� �֧X
&&n""$�����nbqӶ`��2�˺E�ڨ��Wf ���&bc]����|`z�h�	*��0�bƟ�Ǌ%1I�<5�����y8kx�6^��Ln�T�nL�F�<Ƥ�A���|��/�����S���w�����_�m������"������?D�舘��_��`�w��=����fbG���Ħ"6������ ku��&&�O��޾0�U���B�.����0?DD���o� �O��=y�"%n�q�{G6�E�
dl$��=ϫz�]�޲���{�� �?"� q�$�F�7�#e��X�#R�����'4���E,����@B�Մ#�MJ�)-U���"�lTO�0��~"� o��Oҁ �*�@H�D��I�Z[al+�$H��!�E(iH�Y[�AQ��E � Ac�J�Wp�$V1$R0"1$l� ��mZ���3��	�,`)FZ��RS7�}��o��         ��   m�        m  �MgY�o7�u�&��J�gI$��Y�z����&�v3q�m�(OR�ks�bB,��Yw87SX����+m]h�Wn���ic���I�£gB�;sӰ�B�Y�dJvғ�
6�V�n���m����S`�Mu���[t�����F�c���6�붮���j��1�{�d����\i�#�lz��&�Wt�,�!G&h%Z��b�餓  ��[]q�28�U\�:>��=6���5qvp5�9
g3m��Sn-9��Y�7s��q�i'0<���i�n.�G]%�صv�l���[InN��,��5�6�e2��Z���n :���Q<�9B���z��d��UUW<��U�����=<����UA75����]6�(N���6�C4�t�X.�4R��A��T`�7 �9�Y�ct�Q��hxj�z7E��Qv�j�#v���Innd��d�*�:�Ls�� m����j�q�V��I�JU����C@�T��@���B��s;v�bĥ�.ǹ6*m*��ѭ٪�F%ۃ�xG$���t�Ts؍�ވ�g�e�B�4S��r�T�[viOn0H�n��E�Nj���t����-�.��$�.�u���JU�^s.�*ͨ�N1����S�%�g�(a]v\.�#��1R����s4�P��R����n�s�w# ��Yz�7um�t-V;l!GA7L�	A+)u=͍*��]���)���U�n���U�ࠠ��ۊ���S����9�e
�m�sո�D�r�t��3M��u-[S�*�]!�6�˺d
��pͻm&�;��X`
&�يZ�V�s.i��yչ�6�mr��[3�x���+��>g�[;v�@�)�.�-2�`��,qʖ�GK ��˻Zh�.K�U��� A�>M� M
#�`�16	�Ƞf}������̶�[@��l�z#B�_5�7:�����G,��Z�u�{`e-iN��;�� �N6��
CWM�4`����7������î�0뵻q���A�y�Z0�%Ktj6��s��=�&�W�e��ho$��gn��)9gK��5m]�˚W#�]�Ы����6�v�*.���e�^KC�<��kl�>�ir��Z����C�y�
l�/��jҒQYDV�F٬u��0�;���1�"닡n���w������2BFF���ۚ�e4^n�ff>A����s���*�]݊��*���.]%`��XGw7����H��?�!#D�&܊C@����׮��YM �F��7�5�zg�b�w�����{�SC���U��= ����$$�(��EwwK ��{ ����n�,6�������x���؝v" ɭ�^6W�;���Ԣ��V:���i�|�ܔ�F�s<���4^��׮����c���Dl�#p�9{���D#���t����֧3[��`�~��7vٟ�ff!#�9.9p+�$��/?��@�빧�1+l��*�z�w�2d��&8�z수�����w�����Oo�� y�_G"�AI��Rf��Қ�_wW�5�]x���wA%tQ�.���8�������ͣњ0�����k�+�`��45�v�'�O�����I��u����r%�bX�{���@�蚉bX����6��bX�%���՟�˚��j�f�M\�m9ı,N��kٴ�Kı>�}�iȖ%�bw���"X�%��}�ki�6%�b_{�׌�33-����˚�fӑ,K�����"X�%����6��c��T����2&�w_{��r%�bX��}�fӑ,K���v���ї3Zѭk�"X�
@�O{�ߍ�"X�%��w��[ND�,K����m9ı,O��p�r%�bX�za<kژj噭L�5�m9ı,N��{[ND�,K����m9ı,O��p�r%�bX��}�iȖ%�b~��5�=s2�f�SV�l��ۆ1�t�ר�97!H�4$��+�l[�F��Ě�������%�bw_{^ͧ"X�%����ND�,K��m9ı,N��{[ND�,K��{���ə�a����r%�bX�{���ı;���ӑ,K������Kı/�{ٴ�O�T5SQ,Ov[�5ɬ˙�.a$��6��bX�'���ND�,K����ӑ,KĿ��fӑ,K�����"X�%���~�k535ffeֵ�s&ӑ,K������Kı/�{ٴ�Kı>�}�iȖ%���H�qq�O{���ND�,K�����̋%Id���{��7��/�{ٴ�Kı>�}�iȖ%�bw�ߦӑ,K������Kı���{���ߝ�?��njZfk�̍�qu�
��{��09U�);Y�ڰ7U���/ή�̶fffd˙�O�,K�����m9ı,N����r%�bX�������bX�%��{6��bX�'��D�����Y�֍kXm9ı,N����r�!�MD�=��kiȖ%�b_����iȖ%�b}���ӑ,K���	�٫��Y���Lֲm9ı,N��{[ND�,K����ND�ı>�}�iȖ%�bw�ߦӑ,K����6x����I�&k5��Kı/�{ٴ�Kı>�}�iȖ%�bw�ߦӑ,K������Kı?jw��<\0̙�&ff�6��bX�'��m9ı,N����r%�bX�������bX�%��{6��bX�$��1Q'��ffffffd��f  m��S�M��k[�V�:��ɰg��3��Ea��޶����fs�FE�m��l�t��5s�F��]f�N,��k�K��n��q��N2�U��tVNbson�jtQ�l��L7Bͭ�BL��Y�o5`�g�c<�I,p��m�"V��Ok^�omTe�jĝ�9$�%��]]���q^��V�c�C���,�ZG� ~E��eٮK�D�v�8�ۜ�Ĉ�ˤ�3q���ʵ��R`+��{Y�EV+��]���oq�X�'����r%�bX�������bX�%��{6�@�Q,K������<�<�<�<�����`]�s��Kı;���m9�B:���%����6��bX�'���iȖ%�bw��6�� X�%�{�M_kY�˭f�fj����ӑ,KĿ��fӑ,K�����"X�b؝�}��$�uoud�L�z�UEUREUU��0�$}�w�6��bX�'�{��r%�bX�������bX�'����ӑ,K���v���ї3Zѭk�"X�%����6��bX� w_{��r%�bX�k�{[ND�,K�w�6���oq����ߊ}��av���	Icaf��r+��=a�:�xII��u�B��Q��f�4j�6��bX�'u����"X�%�������Kı>�}�a�
�D�K������Kı>��62Ma��3$�f���bX�'����Ӑ�dK�����"X�%���ߦӑ,K������Kı?}������d�ї3Y��"X�%����ND�,K��ߦӑ,K������Kı>������bX�'Ot����e�̗0��5�iȖ%�b~����r%�bX��{�m9ı,O��}��"X�%�ｿM�"X�%������S�5P��[��{��7���w��ӑ,K��_w��r%�bX�����r%�bX����6��bX�{��~vP��){ܒ���/��q�v�:{'�/+r��D����vŽ3�ư�V1Y�3W&�f���X�%��w���r%�bX�����r%�bX����6��bX�'���[ND�,K��ּf��n\�kYf�5��Kı=����?�T#���b}���M�"X�%���{�[ND�,K�}�kiȟ��ꦢX��������\iUk|�~oq���������ӑ,K����kiȖ?���C����7��s[ND�,K�����ND�,K��gOf��fkSF�d�r%�bX��{�m9ı,O��}��"X�%�ｿM�"X��MD�����ND�,K�����.k�I�&k5��Kı>������bX����6��bX�'ｿM�"X�%��w��ӑ,K��_B�Yl�-�'���w[Z�m�.�:q�4��7n�E� �R�^��N��\�����<�ı=����Kı?}��m9ı,Ok�����bX�'����ӑ,K�����.e�̗0��5�iȖ%�b~����r�uQ,O�{���r%�bX��}���"X�%�ｿM��7�����;�ow����S�5P�љ6��bX�'����m9ı,O��}��"X�%�ｿM�"X�%���|��{�7���{��>�����D�RY���r%�`؟k��[ND�,K�{~�ND�,K��ߦӑ,Kq?���7"s����r%�bX���kq��F�����u�u�u�w��ﾛND�,K��ߦӑ,K����kiȖ%�b}���m9ı,O}��}ڀk�\3��	s#�3K���˸խ�X�͂��7R�e������z.4���ɴ�Kı?}��m9ı,Ok�����bX�'����ӑ,K����&>&0��Lkk$Q�J╢��̛ND�,K��}��"X�%���ﵴ�Kı=����Kı?}��m9�&�j%��O�l�.k�I�&k5��Kı;���[ND�,K�{~�ND��Hj&�}���M�"X�%���{�[ND�,K��{�].fL�s5��r%�`؞����r%�bX����6��bX�'���[ND�,�&�w;��m9ı,O�)��K�s3%�$��d�r%�bX����6��bX����{�[O�,K����m9ı,O}��m9ı,N�y�y����t���m�6�*�Z��Ć�u�C�;)�J;��rX�mk��|sOlvm��ۄu��()l��N6�wh��̡�8�>�ݰ�5)��8h*t覵�q�lĹ"�u�p�C��]�VN8U�h���zum�b�x�z�.�c��;f�Z�5p:�s���6�ݰ�n$��灳fʊC7h��^)��.u�\׋%��v<!������+e�]x�n��;Wa�۶�)^�{ ��f�c-����X��m5)����j�2~ND�,K�^�����bX�'����ӑ,K���ߦӑ,K������Kı/����fk5sY����5s5��Kı>�������uQ,O��o�m9ı,O�����Kı=����r-�bX����0���r�f��ff���bX�'���6��bX�'ｿM�"X�%��w��ӑ,K��_w��r%�bX�׉�ښ�2�fkZ5�a��Kı?}��m9ı,N��{[ND�,K�}�kiȖ%�X�{���Kı>��Ox��]e��M��iȖ%�bw_{��r%�bX�k��[ND�,K�w�6��bX�'ｿM�"X�%�����C�骵 �g=�ۖ��\O&x�۹�n�s7;�i�^]�/�y}�'��W;8�5��r%�bX�k��[ND�,K�w�6��bX�'ｿM��3�MD�,Ok����r%�bX�w/����a�34fe�fӑ,K�����!W���������bk�ߦӑ,K������r%�bX��}��r%�bX��J{\�2�f[��ə�m9ı,O���m9ı,N��{[ND�Vı/��ٴ�Kı>�}�iȆ��ow߱��gS�XY�[��{�K������Kı/��ٴ�Kı>�}�iȖ%�)b}���i�����oq���O�4�E���9ı,K���m9ı,?����ߍ��%�bw����r%�bX�������bX�%����׉��\��b�Q��]�M�/mn�B������9bA�|��;�6���6q�|��Y�X�'��m9ı,O���m9ı,N��{[ND�,K�｛ND�,K��;��SWF\,�kF��6��bX�'���6���@�MD�=��kiȖ%�b_����ND�,K�w�6��bX�'}0��&fYfkSF�d�r%�bX�������bX�%��{6��cE�qH�#`�X����d!(��XlCF)7u�DP�R)]�W�8���Ut���&����@�7�сF	a%�%"�X�0%�)!�Q�`F� @�R� DX�#u
��
��k®U� �� @�4CP���H��c� %A����uN�"A#IUaE4k��>آ�8:EC����P��t|�E�D?��W�C����br'����ӑ,K���ߦӑ,K����6x�a�35&d���ӑ,KP�/��ٴ�Kı>�}�iȖ%�b}���iȖ%�bw_{��r%�bX����B��p�2fh�ˬͧ"X�%����ND�,K� }�M��%�b{]���ӑ,KĿ��fӑ,K����kV�$Ɇ����ɣ3�P{t��WoQ7Js2̹mWutM���nu�ә)B�,����Sγγγ����~�ND�,K����ӑ,KĿ��f��Kı>�}�iȖ%�g�����3��<Ί�=ߛ�oq��N��{[ND�,K�｛ND�,K�w�6��bX�'���6���X���~���ٙV
"�O�w���bX���{[ND�,K�w�6��bX�'���6��bX�'u����"X���}���z��U5�~{�7��,A[�w�6��bX�'���6��bX�'u����"X��P]�A熓v&��{[ND�,K��B�)U�⋪�������D�&1��ӑ,K������Kı?k�����bX�'��m9ı,O�{�����g�<g�&�㞭شXX���/S%�`Rs�n��b)��;aߝ����|�$���,�jkW2m?D�,K�������bX�'�w��ӑ,K�����"X�%��{�M�"X�%����vz�0��5&jL�kiȖ%�b~�}�m9ı>�}�iȖ%�b}���iȖ%�bw_{��r%�bX����B��p�2fh�e�kiȖ%�b}���ӑ,K���ߦӑ,lK����ӑ,K������r%�bX��H{\�2�%��d��6��bY�Q;�s�m9ı,Ok����r%�bX���{[ND�,K�w�6��bX��}��Fu=5���[��{��7�����ӑ,K��Ec�{��[O�,K�����m9ı,O��p�r=g�g�g����w�����Ŵ*��_	��+�t时9e��1wS�rZ�m����kM�+-;[g]a��JL99�Ũ9�\�ɂ3ّGv#sp�bknt�6gF�������c��KfX�.�q�m�w�����lE�[,m=m��C�hۙG�<����
�O<��=i'Sۋ]pAX��:nd��r��&��sNP�<y���n��Gg�����wf�o?;]������aںǮ�7A���wi����^�8������G�o�2�j��S�����{��7�����~'"X�%����ND�,K���6��bX�'u����"X�%�}��ٛUA-i�����7���{��~�vӑ,K�����"X�%��}�kiȖ%�b~�;��O�T"��<�q����o��F�Ε�n�����%�b}�p�r%�bX�������c�D�O����ND�,K�����Kı>��Ox��]e��M��iȖ%�X�������bX�'ﳾ�ND�,K�w�6��bX�'��c�a�DǴs��]��.�\WY'"X�%����ӑ,K�E>�}�iȖ%�b}�o�iȖ%�bw_{��r%�bX�}�Mj�5���-.d�$�T"�tˮ;Ln�5pa�����wT	�.��\�F�닮�OU|�~oq���>�}�iȖ%�b}�o�iȖ%�bw_{��r%�bX�w=��Kı/��ї2�Y��e�30�r%�bX�w���rq@P���j%��}�kiȖ%�b}�{�iȖ%�b}���iȖ%�b{�}�5�L��tk5�Y�iȖ%�bw_{��r%�bX�w=��KU�,O���m9ı,O���m9ı,K�zOf�Y�kD����nf���bX�'��z�9ı,O���m9ı,O���m9ıE����ӑ,KĿ��{&�SX��������7���{����O��D�,K��}����ı,O�{���r%�bX�w=��Kı/{�g��*�m���m���Ml����k��*:�^�4㮈��NF':��f]�"X�%��}�M�"X�%��w��ӑ,K����]�"X�%��޻ND�,K�L$����,�jkWY�iȖ%�b{]ﵴ�Kı>�{�iȖ%�b{���ӑ,K���ߦӐBı,O�<��˙&��Ԛ�f�[ND�,K��v��bX�'��z�9��j&�k�ߦӑ,K����kiȖ%�b}���Ip�2fh�̺˴�K��g�v��bX�'���6��bX�'���[ND�,騝����ӑ,KĿ��!��.eֳ%��s.e�r%�bX�w���r%�bX��{�m9ı,O����r%�bX��=��Kı?�S�߻��;�m��j��n
���t\�q�qru�6����h����֯nhnn�f�k2m>�bX�'�����[ND�,K��v��bX�'��z�9ı,O���m9ı,K�'�Y�ֵ�ffj�3[ND�,K��v���%�b{���ӑ,K���ߦӑ,K����kiȟ�j%�~����k&f�%˙��f�e�r%�bX������Kı>���K,K��}��"X�%��s޻ND�,K��;��SWYsSS3Zֳ2�9ı,O���m9ı,Ok�����bX�'��z�9İ ��Xx�U��8��Q?����iȖ%�bw鄝��3��.�j�2m9ı,Ow��ӑ,K����]�"X�%��޻ND�,K�}�M�"X�%���-���L���u�e�v����F�g`�:�7�,����{\�r:n�gڶ+e�b鯞���7���'����9ı,O}���r%�bX��}��@�Q,K����ӑ,K�������3&f��˙v��bX�'��z�9ı,K���m9ı,Ow��ӑ,K����]�"Ab��H��H{D֬�&�5�kpI���fĐI�}�M�$OD���]�"X�%��޻ND�,K�e���S3Ffe�5��\��r%�bX��}ͧ"X�%��s��ND�,K�g�v��bX�b_���iȖ%�b_}�>�ʽ��گ����7���{�߷ߧ��Kı=�{�iȖ%�b_��fӑ,K��{�m9ı,M(b��w�w￟�� �  &ݻ*l�15\텷�������}v֒���{��Mq$��	Uʯ�Ύ4n�����+1�<\C�&��S@W[Tm����Z����x�qs�z�uU���u<��qq
�3���;\O\u�ٳ���pg�����Js�&�	�<Z�f�Ӯ���kf;qx�$0������$�6\�h㍶�ݖ6Į]b�si�[���k26��:� ��N{��*�a�2�6�������*��ɚ�m>�bX�'����r%�bX��{ٴ�Kı=����r%�bY1�ϫ&>&0��Lut�u���E浭fe�r%�bX��{ٴ�Kı=����r%�bX�k�����bX�'��z�9Kı;�]�_I���Y�Fj�3iȖ%�b{]ﵴ�Kı>׻�m9��D��������Kı/����ND�,K��3~��I�35&����ӑ,K?�"�j's����r%�bX������Kı/�{ٴ�Kı=����r%�bX�vz���\0̙�5�u��ӑ,K����]�"X�%�~��ͧ"X�%��w��ӑ,K��_{��r%�bY��}��>s���n������H˷[jc���c�\k*��n�W!B<�=��%v�E�WXL̷2�]�"X�%�~��ͧ"X�%��w��ӑ,K��_{��r%�bX��=��Kı=ܽ��jfh�̷F�Z˙�ND�,K��}��!Ј)���bw]�5��Kı=�{�iȖ%�b_���iȖ%�b_߻~��U�WI`���{��7��������"X�%��޻ND��!���{����r%�bX�������Kı����~��Ҩؔ���Sγγ���`j'�w��v��bX�%���iȖ%�b{]ﵴ�Kı>�������{��7�������#b�����ı,K���m9ı,?�!�������X�%��w��[ND�,K�w~�ND�,KﳳZ����.���u��3/F�^υ×�C���%0=�m��^�ع�m[U�<SW�w���oq�ߺ���ӑ,K��_{��r%�bX�{���r%�bX����r%�bX���f�2MfLԗ	��m9ı,O�����"6%�b}���iȖ%�b_���iȖ%�bw_{��r%�bX�vz���\0̙�5�u��ӑ,K���ߦӑ,KĿ}�fӑ,`��`�@R�EH�ȩ�O�"$�
A1DP��I"{^��[ND�,K�����r%�bX���h˙uu���ff�m9ı,O��z�9ı,N��{[ND�,K�}�kiȖ%�b}�����{��7��￱��f'���6��ND�,K����ӑ,K��B(�;�����%�bw����ND�,K�޻ND�,K��ɭ[�Z�s'c�1:��"ۺ��e|�����VS�:ۚZ�Ӫ8�Va^�t�
~{�7���x�>������bX�'���6��bX�'�g�v��%�bX�������b�oq�}>��j������~oq�X�'���6��bX�'�g�v��bX�'u����"X�%�������K7����߯\���R�������%�b}�{�iȖ%�bw_{��r%�bX�k�{[ND�,K�w~�ND�,K�L$�����,ˣZ��v��bX�%���m9ı,O�����"X�%����M�"X���pq7����v��bX�'������	�ɚ�䙬ͧ"X�%�������Kı>�w��Kı>�=��Kı/~��iȖ%�bw]�����D&�J�u�V���ҝ�A䛵�C� �TV��]Z�h\�ӑ,K���ߦӑ,K�����ӑ,KĽ��ͪ�"X�%�������Kı/~!�s.����nY�ɴ�Kı>�=��Kı/~��iȖ%�b}���m9ı,O���m9Vı,Ow/}u�˚3Y���k&f]�"X�%�{���ND�,K��}v��bX�'���6��bX�'��v��bX�%�d��e��sX\��s3iȖ%���Q;����9ı,N�{�iȖ%�b~�{�iȖ%��X��{ٴ�Kı/�_k?l��R�#=ߛ�oq�������6��bX�'��v��bX�%���m9ı,O����r%�bX�oI �0�Z<>��	6�CA��!k��`:5���1# C-+���XT��PСBQ,��6��B"IH[Q!�4 ���X24HAЭ����+�|.�� @�H��OX?j󹙙�����       ��   m��       @�UUA\��:��U��U�M�x�v��T�T�;�7M�f�-(����%	%�0��!\v��Rqv�ʽ;Z�l::�{;V�!uz;]s1s��Ӹ�m�!ض�*'N�>͕����yؓ���9$���6R4��ť�#=qš�Gq$����QD�7U�gk�Ύ��m�y���a6SDz��Ɖ��Ɖ�؝q�N��l3���Y����N�t ��nn���ki]�[i����  �˦�k�sj��X:=��5���V�l�D��eL�;GU����eF�Þ6�d��$۳�v�$����<�uv�ui) �y�������n�6D&�&�2s�-��X��mUAԱ:�ʆ$��!�����1��ۯ[Y;X����L���6��:V�0�d0	6�mk/,ۤ�;N��ɑa���T��e��H���r��P.��yۀa(- Y�kb����rfJ�P+<���{RnT��Y�xxL�ʆ�Z������Z�.��4RJ�MHh8�1�Fi�u�MVʅ�G.y�x��qShr�s�i�誊�Pζ�s�L�D�73������0��!�͔X@�wA��.�m��J[�p!�͗3.^$��H�����U�୵4lUC�4���A�!ӛ+�d,7�۲qm�n�S(��I@eų�[ v9]�{;M$�t�5;��OJtWQ�6M�=f\�ml��n��)�Y��YUW�
��f��j�=���"�']�Mۤ�e�eX:���k�Z���J�
���ӳ]��\&��Թ�@�le�YV�vz�LGNѲN�;qk�k�Nu]HNu��mI*��uQK��sp�ˤ .ݴP[v�ej���MF�M�̭�*Ӳ�mE#M؃�(m�:�ɏ���5�L6ݸS�vf�[�#=<<v�g�6���+ ��n�Slg��w ~J���&�O�E��� *G��S�GD�U	ݠUZ N�ߞ�� 0 �Ôb�G�]�<��t��M�p���phϝT���vg2h�<:��Tάi!�g�=�sZqn_.�um��œ^�"��:D��I���Y��:�ɮ.9s69Y1�خ0�Q)Y{�4WH��u��dQ<`�Vi�N���v足g:�+���1�nL��bl\)g���{��lݖ귳�/�oTp��`w&y�֨}��9Knn�Ө�ۄ����m&<rn]�o[�i�CsٺL�*=<�H�k�Kk5��Ȗ%�b}��ӑ,KĽ��ͧ"X�%��s���R(~���%���o�m9ı,O��{�L��\֦]��˴�Kı/~��iȖ%�b}��ӑ,K���ߦӑ,K�����Ӑı,O�N���w]�@�.��c�a�Dƻ}v��bX�'���6��bX�'��v��bX�%���m9ı,O�=avx�a��4\��e�r%�bX�{���r%�bX�����r%�bX��{ٴ�K�lO����r%�bX��I;�.e��3-�3Y6��bX�'��v��bX�%��{6��bX�'����9ı,O���m9ı,�~�~��]z{6�v�f�:;v�g6���.�]nڌ�l7n53�sv������ѾC�Fk2��a32�9ı,K���m9ı,O����r%�bX�w���
$�Q,K�g���r%�bX����`R�"�����7���{�߹�]�!����~@L6���%���ɴ�Kı=����r%�bX��}��rbX�%��|k�5�ֵ�35��W2�9ı,O���m9ı,O����r%�bX��}��r%�bX�w=��Kı;�����̳L�k&f�m9ı,O����r%�bX��}��r%�bX�w=��K�U,O���m9ı,O�0���33W5��E��˴�Kı/��ٴ�Kı>�{�iȖ%�b}���iȖ%�b}���ӑ,K��{���ė�k`�V���x����[�^�q=�z�\r�M�c��]��gGK��ww_c�l���i*.=O�,K�����9ı,O���m9ı,O����r%�bX��}��r%�bX�vz�z�.fe�35��ND�,K��~�ND�,K��v��bX�%��{6��bX�'��z�9ı/}�Ohˬ���fe�3Y6��bX�'��z�9ı,K���m9����HQJE"@dd��CB��]��ȝ�}��Kı?w���r%�bX���n����32]�a32�9ı,O��}��"X�%��s޻ND�,K��ߦӑ,K�D!������ӑ,KĿzj��$��13�������ow�������bX�'ｿM�"X�%��s޻ND�,K�}�kiȖ%�b_�-�{���]-Vu�IL�t^�!�(A6�L�^�aw,N����A�YX�j)]����D�&����5�r�<���D�LG�5�r�58ꎺT�.�.ꬻ�0u"�9s��s��.�{��G|<�I28��ԑh���uH��p�9ԋ �։�w�ʠWJ�� �R,z\0u"���{�s=4��V��E�Ю..�]B���X��`�E�r�+ ��(ʠ���۫y""p�-�nш����Ez�X�0wd�8�7;l�1.U΂Ռ0�6�/k��뮉���{z��>GT�qG�H'�9��h^������`޾0�6��DLEPo�)UW�]]�\ZB����߫ ��ه艉J���r����+���#�90���{{8��r�<���;�LLE;���U����8��&��G��Z艉��}_��V��� ����&IY�����"�������  6���K$�O3� ;]��[e��6޻d����n9��֝[*N���Mbu�v�N���lF���cS�����$ݱ%{]����]����m��U�l�&�*��gkȓ��k6��*h�y#a�b1h�;�y뉃t��ֹx�t�N�\jm�ޭ�e��>�� Б�W<<����F�01��!	l�!fr����{ Լ�P{���t�3g����9Mu�m�=�����Rs�i# �L%�o$�Tt���h�ڋ�<�~���Λ_Ȉ���=��u��ϱ8A�Hr=��z��h�j�9u�@�a�.)�$�<R$��=]�@�;V�fffbU_�z/��@:�u�qF�)"S"�h�j�=w�y=u��3��r�9�|�P�D�H�Š�f��3������|h�j��T1��L1)��U�ںǙ�۠�e8��U�^������-�
�m��̍(������`�m~�����ϯ =�tWYT��f�3Y��f�$���۸�
�����__���z��玸��I�uUe�Y�o���kw�虉�KW>z���@�<BIm�LmI�tr�Q��T� }R,�G��¨����U������33����/?�Z��h��kTx<s�
B	�U�0���۝��^y��g\�:�Mqu��'�D�2d�G�D�z��4�h�hW����N(��$J����7�����"f"���x_��=��ZG�:�P�D�H�ŲI��w7$�{�u���? �Od��L}�vY���k =�)US��ګ���]�鈉��ϫ {�r�7���^�@?T�;�l��&G�>�E�>� tr�Q������ѮF5[LBI��d2k!�,���#�1I��X�����{�ĳ�Wm+�FE��z�������ZQ�Z8�l���"�^�g�311Tj�V޳��V��fb"%#�Q�L��Lr�����|���Zyڴ׬�=�_苊d�"�H�]`tDG蘙���?,�~���]�8����V QX(�$n�z|X)nb�%2FE�w�E���r��Ȱ������|w'�i��.c
k-h	�:��랸֍Q����N�����AI��=���|3�~0Zi'�H�����������Zyڴ�ᦝpM�9�%�@�k �;�7���=w�12�{���cj6)#�a$z���;�ՠ�f��z��\:����FZ�7���=w�y=u��)�a�@��F�i�ڒ- ��4+���
��h�=k�$�Iim �u��m�Wl����gj.-������^$yyi�Y�.�e�n�NDv8�2�!-���ٽ��\��n:ݵ�L��[���`ү��Xr���>V�4�ݫu����ʲ�6&�O<� �����"3�U�j�lv�����ڹ:�<�<oc#[���!���<]�r!u�랞��8hg���*P�&�q�&J��d���'"��Z���n���l��t��$�^F�T��{[x��<�����.��Fn4"^GLa���\=sYv9���߫���v5�o���&&g����5�����ɒ<l�=�aV��v� ��4+����
E���L������ y�?��"f"���������Q�N�(I"O$�#�@=z^�9X�dX�`s)R�V*�.�.ҵwx��X阘��3<��~^�~���]�7pU$��)TRJ\�zk���� ;�f.^���P�!��G\�u�'�1���0�=��U�w��@=z���z*�u�8ҟ�e�f\2�I��w�t�2�T�"#�¨sb(��!���s��'׽����U����H��F�lrB5$Z���'���8k �Sk ��Ip�T\U�T
*���Ḓ�}X���h�j�^�@�eG�E�2d��8��;��Zyڴ׬�^�M������=��.�`��K��N��u���=':�ď
�Mғ�
'�w����>X���RD�E2/�^|�׬�^�@�;�h��$y�y$�Z����^ ����T�?=��䃺�4�yP�c��I���h�s�r���XT�$ ������.�W4"� �Hh4\�iB$P�R0!`��h2�;)  c�`T�"VT%ւ�*�E��kJ�m���"�a�"� E(��4$M1�ЅHRQe`ѕ"�!pփIhM	;4�
���e֗����!�/ L QWh�?�b i8�0�ADĈ��&bc�[� 5�x��N.�mF�$rd�M��U�w��@=z���?���@��G�$q�1�7$Sְ�"��^ tr��=�}���_�O�]X8�d�f�l=���	��ڂ����L�$�sY��d�������Wv� �}x���8k�""c�O�9��� }�\~�Qt]��E]]�G/ }S�`�E����?�.)�$$x��&��w*�;�է����h}~�}�u��F�)"S"����&bbS��X����]�8���s?��:L�@�iru�<�A<�d�k <��з�_�=��X��X�`�W"�Ģ��L��l�cLZa�\��/;��:�s���λf���vn�g�dFz�c��I���M��U�w��@=z� �y;�1�4)#p�I�w�ʷ��y�����4׬�9Uì�ƣ#rE2-��Z��h�Y�w�ʴ��$i���!$�@=\� ����z,]H�d�����Wb�QWWx��xLLDK����'��޻�O����'T���QtDO������   �5tWN�Ux2�J�N�/h����#Y�d���s=Z6��R���6�N�]d��)z�����D<�Sn�����V��I�&����!bdhN�;[۫3C�6�&� ����hRs6-k/k�qJ��jy2ǘm�6�ζ�M]6�΍���Ǳ�+��y�ol�qv�2̓,�<��/J���w{mD��\�,�%'r��s&kZBԥ�׫[��t�t���H<�n�F��uEl���"b�2BG�rps�*�?s�h�Y��@/�ΰR(��$Je���]H����ܼ�OE�_4�:�G �I!Z��h���;��Z�v� ��`ۏ"�ߪ�uwx���T�X��`G&�~�N�c���NI4�V���X���n^ ��T�Q~Wq��'n�.Wm�����n3u�t�0Z��nI3�$yt�gS!y���>m�?���� ����z,��-f�3Y�&feܒ~�����,E}⃛��k��u"�9��.�5 �,qɠ�@�;�i�����K������4\�����L������OE�k� tr�����gX)nb�%2)�h�ڴ׬�*�^��w*�*�6����?����9.
1��'6���LfF�m:��3��Ͳ�D�$y�y$�qh�Y�U����t�L��9�r��u�UuE�9��4
�׿fff$^g�@���Z��h���H�8<�D�wX��5�=�����莉���#�M��|�Up�$q�1�7$Sְ�E��'%`�z,��:��8��$�h�Y�Uּ}N�<鵀t��Ou���H5hj�.I�6�e�������={��:k`�`��зFƢ�Ű٘�k�m�~����z,�H����s�G։�~�!#Ƈ#�;��Z��h�Y�r�^�_a�`�Q��H�ȦE�zԋ :9xNJ�T�X��U(��r	�$qh|�}~�W�t�ܒ6 J<[{����$��,q�Qd�d��@��z����o���s��z� =�IlE8/��"u�II���;��P�m�6��#g�f�]����u9̘�n�?6����V�yڴ׬�*�^�ʮd�4�2F�dZ��h�Y�r�^��w*�=��$i��rb�- ��x�n�鈉I�tr�7��`�`��q&	�&�˭zyܫ@�v� ��4vTD\S&HH�� �S������/�7�^�[�d����_��� ej緈Wa�C{Gj�DOm���X'��E6[<��m�d��x6L��EOFq��K�vþ	��q�n���Y��i��e��OmݚEb��mY�=�0��fEnh:{*����m!u�+��jt��!u�n��;-�5=���%�(�����7D�s���7/<Z��/<�Z-�g<Q�ٶ��p/F�Y/�wc��w4�TA?�����޷5�s2\!�bH�,9���I��:�֫�&�g%[�l��r�k�;��������~�����z��.���r��K���#�Uwuk <��&&R}Հ=��X��h�qǒ5"sd�M����=ҤX����T���ؤ��$�@�;�h�ՠ�f�ٙ����|�
�T2G0s6�dZ��h�Y�r�^��w*��tx��d�L��'��ME8�7	/2��L$g��Fۊ�N�d{Q����I���wk <���[�}N虙��|��hZ�0_yQ&	�&���Y�^Cu=� �R, �������$$x��zyܫ@�v�>��鈄��׀4�� ��v+.�\*�W�-`&&V��, �}x�n��\�@��5a!��&H��^� i�XꞋ �R, ��"��k��L��;�5�8�O+�[�ƛ8tvH��u�a�V���w��,��;SvmMހ?��xꞋ }R-��:J���$cj6)#p�I�{ϰ�{��X��x��bR���.�ી���U��ܰ�]��&b �H�h	�E֧��srN}����>��dj9	1I�z����h�p�L�'�ܰt� \
��Չ�8��^�@�;�h�j�^�@��Z(���2A�()#d���z�h�n�k�[\u��)�Za.mѽ���$#x��&��w*�;�ՠ�f�z��}�u������L�dZy���ba �}x����8k ~��\�nA<�d�- ��4׬�;��Zyڴ�X8�`Ԙ�$�����Ky��k������D��f'�ff*�_^ {����*��
��rI�w�ʴ�h�Y��f�^�C�sd���G ۆLC/]d!�8$���\<�z&�-�+]3C:gH�Wv�-`�m`���=w�ffc�����/��� آ�BLRE��^ tr��= ��X:S��8�L�M ��4�V�fg��%y�����4vT.)0����*� }S�`�E�� �����
2b�%2)�h�ڴ׮nI?}�srO�k�n�w@"!�E!JA����,$��4�FԅeHT�HQ�X��"�#!&��F��Ё4�*X4b�����)� J@*�! @
���	RT�C`�D4����4B�RX�Y��A*�������u�l��x��cXW�K���(Lی�2�ǋ
B�(�*
�R�9M)Gi Q����ҡ*��Me��gٙ���      �� ۶�l   �i        �-�  ��ajɯm�hm��r�)��t���"5+�����[7okT����]2�.-� �y#���K��l��.��J3�e�/�e9%�A	_�����������zݮs��GD��d�kl��L`6Iy]]�:��R�;:u��.�����9��pᴑuZ�d�f8��x��K;���P �k�J���&L�v��4 �c"�vd8�@���U�  86�t�ݧM���x:��uh����k�3p�<B���-Py�*�Dv$��]xw<S�-��:2�E/M6�R��F��Y�L����u:{D���l�s֦��S�\�G�Έ��76�5]����2Ÿ!n�u��ג��E���M5������e��M�M��P-��Z�MUHFf�����'���a�Kq2[U+��5E� ��q����-�v���$�+��n�L���͝��������ዄ��WiC	$��K4��gn�n� �ݖ�����d�%����P�����̆�&MT[^�B�#C�vT�.FgM#L�% \a�q���SU{]�sV%�A7)-G.�;vh�X�ӽ�B�Y6Iz��×MÑ�d,\�h�&ٶ��uURz2 �M+�m����[Pu�Z��@�M\�cG]�l��UL�L�����$j�'	����%%�i�Mt��)(\�yՒԭ�q����Pgk�fӚhbI�d��[h^��tE2OJ-c��X���,0�.ƥ�U�j�(%[�v*5.4λ�j�Z���Vie���k�.K�XvՇ�uJ�j�iV����c�$���j�8�N��[��5�@ �'W]U��9��
y���08��><��*��'M������nԓ��\�s>�n܄[5 ��ʄ[���g�q6Q�'#�"5�jM[�� ? ��](èQ�(��T/��C�)�꿅 ��i�����ffff`� m�{_4�D�rn�w�k�k���k+c&�^�s�;E�+��v�n��۪i	��Mt�G��s�5��4�l�W@W�Ck�c��mm�5�n�lg�&5,�sv����-΅b�T�5�ޮUrl��4�9�E%�עB3lث��F#qm�90`�/1���ٸ��1�j7F.^�F�mP3�l4�ਙ���]��rK�a�!�����wx~l��wb��9�Y�GV';����C�����]k����=� $Z��w��~:me�=U��ր>���ۮ��8k �i����Ơ���E#�@=�f������ć��� ��z�:&?LD�Por��H��lQ���@��������O�LDL�F���o� ����wW�rdS"�?s�h�Y��C�����O��_�#�A<QE!"$�@<���b!k} ��9`m6�yا�]��л-�k�����n4;i��&7+gFM��.����wb�zbb������>��u"��^�[ve�EE]]��p�t��1�3�13?�'������x��y�&&bR;`��+*�*�Ҹ�qk �Z��h���;��ZG�\�U]�����X3�f���׀����r��;V�^����w�ܼ�OE�k� tr�6��˚g;n���<x������tsb��u��I�җZ�겒�e�$�yܫ@��ՠ�gٟ�o�@���̑�jb#nL�dZ�v� ��h���/�ʴ�hH'�+We�.�`�w��w���&d���*$����[�M��9��۸��Ĩ'��D�����ff������?:����k ��$�
�d��8��/�ʴ��Z{��wY�z��2̌O24�HӉd����a�0�9�'V�+�d[K)��\����>h����JdS"������ �u��V�Q�W#��O$�	V����)�׀v�G,�ր^����M �u��8k�	y�r�o� >ݪqweR��]]U�ww��bfev�G,λ� wﻛ�(lT`�jk��nI�ߴ�$s��ۓ"�����@�/��~ �~��V��|6�M�
H�'t�6f�����LUJ�˝4�Mؒj�M���"@�O#Q�I�H��Y��f�|�U�w��@�5sA<�"�]�� y��1��]�:�Z{���$w��?��)�$$x��&��]���X~���H���[��;�g]��L�dZ�v� ��h���/�ʴ
�����O.�ີ�u��ak}�]��|�}�o;�Ӽ������� A�� �O$���^���ԋ�N�i�z]�l	=����O��Ҽ�Gl݈�Ю��|��J�Bz�u�8/K��	!�0���5	�X���݂��\�ml\��*�4�����lE�����+�����7\`i�^�=�Þ��;]��3[Tq�����Ĉ��ɞ^6{�Rt��tf��Lt��fnI���۶�͗iԏ�6͜k��? �P���w5�vjM�9�9���ѓᗷͶ�ƭ�^S�Kѧ������j٩�y�2�S�\��$�����Ꞌ �R, ���iOT���q��D�h��[�?�=_�- �ߦ�{����u�Ȧ"6�dZ� F��7/ �S�`W� \��r"H�Vנ�@��U��/Y��@�?����"`9#�n^ �OE�k� Ԓ����c�����8,���u��=�F4"����yu7�F�l�:���]N�-���O,��T�X�`I+ :9xO�e]E]ZW�-`�mg�L��I1?�����Հ�~�]8k k�G�X܂y$�Z+k�^�@��U�w��@/u���II��9%������ �Sk �۬ ��q�7c�7$�@��U�w��@�mz��h_��2d���;�K�r�F�̯�ϓxo[�bSREg��L���#���Fܙȴ�h���z����~���`����*��u!&)"�9[^�z��Wr���Z�w1,��G��z����n�7NB ��m8����=��5�� ��:$L���wQUuw��a>��X��X���^�@��:��#q)�L�@}R,�%`G/ r���5FU�$�n̓U�cm�N���Ϧ �� �iKl٣,�$�~��}���%�]Z��u����5ӆ��6��X88����I�4׬�:��h�j��� �R������E����5�o���BC�����@�պ�b��ܓ#���v� �����������""H �&	� *�g��N��;�w�.[�4��x��@:�4]k�:��ht��?DD��_�������-URog�6�ۍQ�\tg<p��z�㪀�Wd���������h'F����|�����ܫ@�v� �l�=����HF�n�*z,�H��/ i�X�g]��L�dZ��hu��JM>��7�����]YeUت$s���f�˭z��V���Z{�RH�$�I&�˭z�8k �� n�x�蘞�����D!Y���=�ٙ�����` m�d`ɻn�h��n�zƛg���e�Sv9���.�\�#��9(-cI�M�I���q�n���mR�\{/]lM�p):0t��V�8��'�ڭ/i��5���g	P4����a�s�EÓk&5�l��n�Okt[k:66��{[�aw��X��9!��uj�qq�og�^"'�����7ϔp���^in��!u�(�W��$��-��OŹ�B'\���!�:�s<���j��N�b�]p��X�-d.k,�fY5W�������� ��X ܗ����.���26�ȦE�w���$����׀yӆ���D$>�GqvU"���x��@-���f���U�w��@�5sA88�44���h��X��X�""}�x���E��..˪����]8k �10����ﾚ��h+�Jȣ9��Q��H��'ktug��v��8%.����X�Qtk��L��ƦE2/�r�@wt�w8��r�;�t� ��y$��]�'��s{@X�U] �&"�<���ӆ��6��f"a#���5��H��h}~�Wr���Z�٠��:��lQ��D�h]ʴ�h[f�z��.��H��Fӊ)�h�j�>�Ɉ���� �}x�p� =b)�QT1N����#!��$�ps����	��q���խY;F�"��$v��I?>Ix������"�9Ҟ�'�FƤ�@=z���V��v� ���LLLJF���E��..˪�����tr�7���j�" J̑�0V�1@#�澊9�"C@J�R$H�W&�E#4�ss�X	P��@�%"0�RP�BH�P�cX!�	m��m"B$0V���J�1A�'��p @�!Dt���uu����T"N��s�
�R)
��ì�#�H	��Ĺ�A�3�q1�.�G���@
|00 E*�Hv �)i �1����S�$�FD��$�v@�$H�`��Aֺ��mUx��Gb�Q�;O�Oá���Tv���U� �`�c�6"�AQb�q,���f��z��.�L��ƦE2-�fd'�ܰ�u����5ӆ��kRD�!H�Z�٠��3��wׯ�WG,}M� ��$Ʀ�pr\k�fSۥ#h���p�n�Rvu!�u�at�۝1uV�n���=�O����~�`�m~���^ {��]ER��n4I&�|�U�w��@/u���o��3?�>_T�dn1Ldm8���y����f�z���V�բ�(�Qa$#�R- ��h�Y���������
H� (
���'ʂ~w_���I�j���Y2�e��]����?D�Om�r��ܰ�Y�{�EY���FH4$��/#sÖu�[ƛ�ʳ�%��]��@�u���N�,'�$#x�rh��Zyڴ�Y��f��Ë��S#$q��L�@�Sk:&% ���y�����33ؑ�:���J)	2G0�- �ߦ�z���V��v�����5�"y#N94׬�/�ʴ�h}�����w������������,��/�ʴWj��f�˭z��<��;�����  m�m����a����,�ƭx���$�%�%�<W]U�����Z�]��ځ�,m���n���xj+h�ۜ�鬀Aъ�BeFخ���ڥx��F��\�u�h�gX��s�ؙ�<��sm�Sș��7�ե��۷5ڮB�M�.x���]��T3g�fخ����n9��3����Z3[��������{v��w����~�ܼݫ����X^��ˬ�>�It{���Z����Չ�mHΖqs���X�_�, {��Z�`���<�Ej �LjE������ؑS���9`t��=��@�%VZ�&�#�@�ֽ�ܫ@�v� ��h�u� �L���܏@�w*�<鵀u�D'O���3��)^FH�S"����Z{��9u�@�w*�?z�J6_�9�71�1&���z��8�W/\��뮛
c�LC���|�	5��ȔRd����~�.����Z��h���Q(�y�qɹ'���[�?�S�#��+� ���̺���7��`�w�18�ER��8�bR=�ܫ@�v� ��h�נUy:�m�SN(�E�t� F��9+ �S�`��PN$� �ƤZ{��>���?�}���h�ՠ{���d"Q�K#-�yMt<�N�� �I�݁�kG=(\hJNG5�cjf
bO$F�#�@�ֽ�ܫ@�v� ��h�j�
�y2B7�r=�ܫ@�v� ��4]k߿�>�)��L��ƦE2-�|�$�߻��.�6����_��nC�>ʴ\�ND���$p�- �r����>��n�G&*�V�R<��H��<���^�g���ƀz���`�T�����+j�+g�rkX3��9�{��)z�Q�G57J]\�g ڍ�8�bR=��U�~���^�@��W�r��q7 �26�QOZ�7�� :9x.r��=~|��y~"���D7 ��@��W�w�ʴ޲����+�y!:*���\�`�z,z\0���y 1 t t�̀����;�4{��PO&HF�nG�w�ʴ��~����ǀ��x�����
��[��t����0��\���J�2��ў���IiaÊv�f�t�d�.�z\0���r�+ }S�`5*pr%��#QHh�Y�y{��;��Z�YM��#��ڜR<��]���_V��a�"a/o_����T;�lQ�����r�����z��f.}~z_8ۖ*�.�QWqk ��ـ~�\�_�j���/�ʴ������]�I$�In���U�v�&ӥ� �:UC��Z�k��(�$x)�+pZb���U���6T�%��;\����P��mΥ�`}h��N:�^367Yp5�;.��nխ��5��n�E�6Z8�/ �S���
�QNѵė,���i�n��Hյv�G����6N]n�㵟tp���j��u�dr]vZ�$�ٸ��V��'d�Z�������ִ\�2墇�)�DҨ���rkW�Mkn't��K\���>B:-��ۛk3��qd��n�8�\�A1f��{�׀y{]`���������կ��	��1F�#�@��W�_;�`y�0����G�)8�p*���꠪����9`y�0�3���������z��#�L�dZ�[� F�����'T�XMH�ʸ�Rd�E!������ϯ��s�>Z�YM��m+����H�D���|m����Z���5ړpIYM����Pn�d�NA��E#ȞHӎO�r���/�ʰ��ɘ���^ >\��*��
���j[���;�];w� ��"(h`I �XP�Rp���V{� <ۼ��� i�S����F�����S@/u����u��s�>Z�yԊD�2H9�� ���9s��N���p�9�s�Ɏb�G&���@�w*�7�� #r�\yx^S�Z�)U֝�2�5���=�F6���6Ag�^�M��':a���Y� X
��캨*���;k���.��r�+ ���įԯ�D�5"����S@/u�����ܫ@�����J)	2F����srO�����ȉ�`A�� � <B� ۮkg�ܓ����@�k֢p�9#y#N94/uz�8k ��ف�e.o� u%]eR��n1)�|�U�~����f���@�|6�L��%��P�a��j0�B�̭���cp�o%P���c�u�.răG����L��r�#i�L���ƀ^�4/uz�V��u"�<�� ��Uf =�y�e#V����9`y�4sW0YqI���C�ɠy{����XtLJ^޾0���>��	0�0̗4]k3[����������'����$��w7%��D| n�޷$��|7�Lq��8ԊdZ�YM ��h^���r���iY	�����`�F-�1�K'V�ힶk<� P�/V,����5�[K��N5R{$�??>=���u�?S��bL��O�5���߿~���rF�F�rh^������s�9`޾0�Έ�����RU�U+�(�q�H����-����^�4/uzT��s#x��c�"��fL����q��^��u��&�� �<�I�����D7 ��4�v}�k������&��}7$� _��
*��������� U� QU��EW��EW��T@?� !P�@@�B�T P�P��EP������T"�0B@T$@T$DE�	T$BDDXAb@T"�T �#P��P��P��Ab�����B�P��E�P�B"0����DX��
�B )E���T 
�(�Q
��B#E��T"B+E�EB @T"�P�DX�@T"�AbP��E��P�E�@T"� �T #E��B �Q�B ��E� ��E���T *�DX�� �P�E�� @T $D���� U� U� QU߀] 
*� U� QU��EW� _� U� QU�@���EW���e5��ƞ`j3�� �s2}p��4�(      @  �   �     ���@A��(U

� �P �� P 
  (���B�PT� RTR�)ER� PX   � � ��   >�|�-�nW�7<��Ӿ�ͽ��}�
;�ڞ[�r�>����-�ow��ڷ>���^��wZg{�| �#DX�  :��淪^�sɥ��ҟp��z�S��;�q7y�_��Up ǉ	 @$LmB�;�7��s����Y_N;)�{� =��{�8�CwZ� ���	/`b ;�2}=^}�K�.O]/y�ﳼY]��z��= ��_mqjU�s�[����-Q����R@�  �@F@ >���ϰ;�{s-�n.�W}����W��S��uŝV�n�� s�+����>�x m^-{����j� ��y�����������s��V]� ��qn�s������z��u�^��B�� 
PP(H� g��m�����|�{��� D j(� $�@ 'a���::  b ��  �3� @ 6� 	  ��:s   ����tvt ;� :2���(   �*&6��� �   ���N����W�j��}��m:��[��}��G�J���η�{�|  �ǻ��y4��� �/�'��O=�{���5�n Nz�۟n���>6w�W��zw�wԫ�  =F�ة*M@� 5O�L�JT   D��PjT   D�*��R*�!����T�А�JR�  "�!�I!2�☔-IG�?������t������u��_o�%	@*�e��AWET�@AW�A_� ��DU8��Ocga#Y�BH�3�D�H��_����ѷ�M,��<�of��$с<�CQ��`j���T!�Ur\�Ϸ�����	 0�<�������C�A"�HX,i�"� �X$H�	���<��tYƇ���x�"H!#�A!(z�D���ٹkV�5�®���������$���r2j����MH2F1�̲�m(�&������o�6���<̘:D�J��_?{�ŧ��[�<}V�bjc$��ɬ���
o��!����)&X8�!0�=���=7��7��>Jl���=��=�3�o���P�K ��ӆ>�`D�d���c A�F$,���O5Ӊ��F%8�6�����h�f�4�4�mۈ���p۵�]I�v���@�i0�#SxI�fdP|]R�s����� �/VN];����p��:|C���adX[ML14@�$���j	M���)���CY=�>c�0��K!���3�q8$CZ�l��l�aHP4�f�# �ӎ���P�I]�9�n<���^>��+�I(fqq�MbMK
j�H�����$�Y�B2%�+��oT��nқ#X�]�n]B�j]���[�l���,&��)&�4�k���A��PX�!L<tb�0��	iH Đ�!#�A�20�]BHR� @�Y%�2]3%$	`�4�Z���fH��̬`ȹJI	Yml)k�b� ��;�0	"#����y�NB�
��(�`�iA� "�Wa^?�
�f��y��]�aN;6L���#��ܒ�hqv$1`�g�-���ѷz$u��@�ĩ��!e�Z�xY�<|�2�Xׄn�C[�KMa��3S˿3|�q �Fk|.sz��@i���H]k)<��^\]o���6��k�
0�,��(�I�FF�,l�B:�i���4:`h @p�6�!�<%Ma���0���5w�NyE��9��ѷ��%���p}ChlB4ц�`O}��)|�N-�XaB#H�R�R:H��OtB��N p�abB#2�	���!�(EEl�`�F$ h�x����T����Yђ�hCh�
C�(B��bƚ'��D�t�0��WA�r���a�D ��c��r]$�m'"R%�CHn<M������S�$CA6� bD��3<��$8M��FD�uGo�c��vl���8��ka��� HMjc����!t�<"qcF`f�/8ƺ6���:!�I�qNIbn	��������B T$c�	���a
ID�D.�o$ޗDo,����
;P�F��Ġi XO<�NkY�9��A$-B���"�||�48Ca$��0��	!�8s��9$+�Ns��� R0���!��7^cXK�e�.��yT���xRR$��HR���ܰ�R�3V��R�V���,Iu]h�/� o{VkW�U;��~ʁ)S�_+, �����X�A�$,i*F$+0�
@
! ��ax&I B�$�ѳ�Y@�A�����04���3�W���;q}]�(:RA"� @�j*iqB
E����	].;8xl�a��y�St��޵���xpRDӃF�cA"�4Ji.����*�p6/�l#]of� �4``�vZ��n�9�7������7��avK&�T�7R��4��]ae.�����
�d��XR�HńCg.�]!�ėF]Ɇ�<��rY�	t�*B�M�
J�H@������l#M8��`c�V�bm�4aCd#�ƢhR%4��E����āMaw1��)��0H�HЍCK���	
iX]No^$����c�"Ky�g��zx� Ąj@����|`�4i"�:b:p6'F�0�9�$9��{���$5<�9��n�bSy��fIKp�*FƆ�4aXQ��)�SA�D�D��q��	�@�XX�h�no|��=#m%a�D�	tK��kCBB�`B�HaCF��n�P�W%��w���]!R*���g�JѨ�� �F B��ܙ����i��	�Q
B�b��˩	B����v1c���xÜRS m����B@���6��(ˢ�Ca��P��ٴ|ԆG�<y��ɸqx��]`l�F Vn<�974:U��b�@��&�s�=��x�Hj��`�bB�"�P�(���D 1�'�pN!�)
q���x�}X�aB	�$V&:4��h$.�IN8��]#��4�Y4h��D��0��CN��A(uF��=tjChK�_�p�0�)BZ�Hf���P��������!�5�Y�$��h����������e4d/�>yh�,hR��������D�,=R#�sFMCq,�K��,
�:LH��c���#]&!�"P�$hh4kI.����e�t\�	�#��^hF���@#�]]��0��i�N$+k.�8A(�2��)���HQ%.��ֲp�,�0�5�2�.��6ˣX��JlaM1�7�5��p�5�|�$ѕ�]k ��+�����@(�A��}�W׷��j���ERN��E7T�$�Cv�]�%/��?9��&	��:׬�WL�%��x�"@$H�Y��+��8pFta����tl�#��4�1����ȒB����p �!�
D�
A�.&;�y.�]�}<R�&O4iq �HӌVO�6�!��ю�6�Z�1�P��N�hh�g��4c����$ PҘ6p��!]8�>���`a�a�#]8��ˑ$�j`a��ƚW;F%8��aMf���]��)��kg�#CN(ā��@b������p8p6p��,��!��������0��@�V-a�Z浳ÑѦ�L�"Sdi��3�y*F��'���`����M���A�<4L�%��.o<�/��F�I	0�
i��� SEp�H,Y����2֯����pk�4�(s7����۬��f��$��U����]�H�ƭz�$�<��T9T�~X�!D�H�V1b��r��d=SBxh� ��@bT�B-.�o^�y��]a.oDߙ��B��BD}P�E����*:�H�A��D)���|� ������4��B0!�!t˦]d.ss���H���b�5�����%4ozeҒ�2� 4��$`H���%'��L�)�5�Syf���3Y˼IN$5�r�&oD75�O$��Q�8�B	M<b�a!	#�x�RK��M��*:�Z5/78f�5�$�=9�8<.��14D!��W���;"W�
���޳�@��Ԧ�l������rhܤܸRS�l%�!��hlxx���$ۦ$cH�%��f��k�0ћ6<X�Y���ڞČZS�P�u�y��0����=ӯcn�]�_zzϿ_��� �@�      ���       � m     �               �                           hq"۶�r�Y`[uuN��V[�6ٲ��I-N�� 6�`9`ٵ�m&�q����,����[A [\���o[�^�� ���G6�6ıwl��
�UUP�t  U���
�-E�'�����KZL  c�ۗ��m'��m�&�V��8;e��p��-�6�M�Cm�M�lmk7Z�X��F�Z5怪U�UW��M������2	����;5W6��g7n�j�L�UR����U�e$�N�x	m���!r�+���iU�\  貑\I�l     @� h f�      �� ���V A�Z�k�ݶ mmff�^n��jV"�M&�0�@3��-�e�i]��\���k�c"d��T�Ie�`�s[Pz�Q�s�v���vT+E�ԵR��W.Y]��j��P-�[%y5���m�\���E ���nC HA� 5�i0 ��m#m5i���9m!�k6�����۶[C� 2�[@�)B����W� Cj��i��&��H��ݪ9�-UP*�B����|�	v�"�a$k�I-q*�EԭBn]�r�b0ۂ9��Kb]#��C��*�vf�V�e��B��4��� [@u�mh H�   � $)D� ���    �        �            �������h�q��7ϟ7|�����%r�zݚ���Z 9!`ݦ4�9& c�NJ�(g�2�Tz���
-$��[W�@l��m q�ҙ���-�  r8ŵ�kn����k�l������US�n5�QRC��"[�m�I��l$n�;y"�8*�U�(;*�R��ZŦ� [%�Y�[J��v��-�c��ᴛ����l   |��m�� ��hyj�.l�V�J�ʐlN�m�l�����$ m\���fͫ��v����Jමm�]���`μ I ���m'M�:۶lWXcj��2�J�UT[@m�ei���uu��<���ƥY*5M&熶ۑ�@UU�k��c7Y,�m� -����N���e��jv�  m� @Hmٴ�n       l��$�`6��a��@ � 8E ��'�o  $ln� [m�Ԁ6�  �mn     ��I�@�	$a$� ��` �~���`%� ��T��H8p��l �mn��m@�\ѫ���j�l�� mm@)+:Zr��uP� ~�����L�5Ur��eX籁�j���V���H�`6�   [@Im  p$5�[e�6��&��ʷv��/h8��� ��l�-�5�n�^��GW7��I:	�j�قi`0�>U��-� 8  �-  ,;7h��:/�I��ͻI�6� &�p� -� ��4�O�|Hz�L[\ �H�� �9�8 Ya�Ul֤�gN�����@�lyi�	  � m� � �f�F��=&��-�h	8-����K�V:lksN��檥e�.�^9�  5Ͳt�$}%-��[v�-��{ �h�r�%d했�s��n��U�V���CUcm�Z�-����$	l� 8 ��^6u�V�)��d�^X /D���hY�#mV�� l�����v���$����N�,��k� YKh�$�ր ����-u���k��Xa �n��( h۵��+k���]J2	 � m��� �Z̀r���ݵ���6���M��lm:�8�C� -�m�ޭ�F˵J��UJK)/*�c4�V��/[��m��k $'A����jK�:��   �[p�c�h []6̀[@�Ze���oav��sl�X`�6���ZI�h�i�b@i��`�^/Pm��$���� �v�5��D�	6�:@�� Zn� ���ڶ�@� -��Am�nݶ�  �n� [@�3`H�a!m  ��ڢݵ�� m�(@kj�eA��e�f��j l��	lh    se궶��p�[L�a�߮�۾��8 m�         6�p  6�&  -��j�9��$)@m�@   Hi�p�l[@  ���-� �߾�ko͝u��g	 	$������Ŵ  � �r����'[@ �%�m�U͋h[��89��n:R�-� m�  �������k�-�h���]�!���� mt��g8�2�ZW8A���K�z��@6�-�&̾� �!m�*�6ٶ�߽��6���  ]�*�*�UUk�n�*-� -�V�8 ��e���]�Z�e��}��hy�v��܀��0��u�j���u[WF֭��nղ� �i-�n�Hm�  	e ��l�p [D��kp �[����`N� 8��*��j����@���� ��6۰ $G-��m���[s��    ����֮i78 m w �����9   mm�  )%-��*ޘ����6�!$� H�  �e�� ��k-�Jڀ�L�$ �h 6� �B��%.۶�@ ~��i[o��� 	/6�M�in�[A��$�kj��D �eؕ�9��j��I�i�:�vR�z�Yˬ�6�Η-� 2z��ݑj����$NӖ�r@�BWvz����V�Uy�������.�k�H�%  m���g��Wb��瀣q�['!��7��T�C5��a���]t�t��j�V!YV�mPn�6����:Jt �vzS2U�T�g��;P�lm��T���ڶE�`	)@k�X��%�^8�mk&��=���n� K(I�lp-�ͿP���kd�>�am:�!d�v-��6�l�v m��z' t�&m&�ŀHX`�   l&^Z��5VyP�5UJ�-�Iy�!ƖT�Im "�VW�f�RZ���m�J� �`�@K�UUWU*�R����*3W�� �!�N6��yn��J�V���n�IzU����.�H[@H �� a��4�mm��K�]�5���G%�%4I@����[]������6ۃa@  6�m �����kh$��X���%I��� �v�f��������!^U���ݻ`�)��A#m�6ض� $M�   �����$B����a�-�m��[y!g�2�z��KX   ��m�km%�r@�p����f[D�;i6-�m��nA��}�χ� j�C�l�&\jڪ��L�� �cm����t�\ $6�#l� *Q���t *�T��;(P l��(�`�N�`8��lZ`�X%P*����Z7ϟ)��(-�m�B�4S�� �m��m�y�p��4�l��u��Ry�m�j�����@����^�  H:� �����m��n�8�٠
+����B��T��y �]��m� $ڤۀ�h	 � $�l۶%6v��0�@�mR�*�A�T1I�l��*����8U��mkr� �Mf�U���۶�[@ $���6�]@mt�/2�"���-�ms���k�ݶ�Ͼ�ﭒ�6�[�@^X-'c pU�*�U -�6ۛnnY([4�ͬ�KnpR� ����� �m�IÉTs�;@T��n1�V t^Y&���r���V�j���J�SUU ��{m�m��Mj�t��U��e�zմ I�-UT�m�US��l�]m8  �B@m��kh�Zu��0     � � >�|��          $         �cm�  T�6݇1z��F�;` �[Y�ͪ�0�Ͷ`  �  � )�ڶ�   @ �P    ��m/V)c� m p/ �m7k\�z�����'-�K�UUc��v��<� m��W I���&��l $ �:m�Y��]kV�А[T��� mmm���h�:][$7]&@6�'6��L׭I�A�t l��m��v��`
���?Q��ղ�l�gd��۷R,W+�e�  $8�[��n�f�m+]�$��᭑�[Y-6�`�	S3��^k������w�R���?�x ����+��Wm(@j4U�Sbx��H����(z��D'���#"�E
�����)@t
+J��S�L �� �^iS�j��4( �!�� ^(!�����Wj+��TO<(��h���(��UM*���C�%G� ��x�mD<��mB�)06 ����� 
�@�,�P��>>�h~b
i�/� pA�*+�`�'����GN�HB$���p}�>@��_���@����� �G�D�A<�X�)�&��>P!�� �����P�b��A�X� ��DD�� +�pA>@��`��6(�������}@��DH!X���PG�}=P^TS��AM�G���H�:"j�������(�ӊ��<>�G��^��"@O�"�Oڿ�m�6���   m�\    �kxF��ʵ�gl�=tn����g���uĪ���]V�!e�-���e|JA�8]�s�� �`m� t��m]�v�a%E�z�k�eu��L�r�*�n�pBTFP@��.��35�y���v�;y6$�J�d�i�{7@��X����R� 5UUC���=�K��x볭�ͧ�����}sv�n6냇O��� � �3tl�S��F��`�q�,a�x�{\f9�`6��	���iu�;Tt�(�]i�V�2A	�{l�7*�p5�rD�F�a��*�mҤWj:�lO1�d���vL�8��D�!��BZNN����׷=)M84uK�����u���]� D�j�kK�ۑ/5�hN��E���n)0����h{������/	��.`M���9ޛn��f͋rn�6!^h䮘Yn�hV[P��j��=�ݬ���]Q�����M�����N�x��Z�sX�2k@�A�׭p/��ݍ:���l��t�1F�ܭ[��7��W�V70MRDV��6�z��P���j���n`قVqt��h�؛���֚\�J��Nɻ<����H-6�B� I��v�ِ�[!�o;v��ll�6�ݎz�e� �@��s6����:EOl�wcu��n��y E�]��C�F�j��+�Kd��[ZR�-GN�7-��]r�ͱe�zւ�!۳������ͣe�,����3dېf۶�U$ݘm�+��V�n�m��v�Ƀs�uCԹ;5F��A�\R�(�me��r�"F0%�S��`,s�.��˲�@w%�L�n�WV��ې��Sm��V�]d��6�[2�c�.PR���е5��nt;'
�9�v�T,����   ��ۨ�6��n�pm�kS+�N�x�,Hm���;�#�(1<�1Ȇ{k�Ѧ�g�G\p2����WY�p_ފ�N�-" ?�P? D�
��Uv>���ww�w�~?[��j���X7Y��񭄻]]30�PIQ��Ö�5�9eت��`˶�]��7'֦�wI�,v�㣲��X��T�z9�ƪ]���\� 6�]����nSp�[qe�L�uq��E��) �l�v7VE��ctO[��;a��-��8�0C���	��q�j6���ce�۫���:S��t���ŹC3҇g����w���{��s��ۗ)�D9x�69�er��l���ܹ^_&э�i�����9����9������P����V ��ҪD岊�钦i��V��%	(ȅ�Q�]�`fonh=n�Ώ���6F��$�-u�Lލ0"�`{nJ`��O�/�Y�]�07z4���i��V�~��تv���XdR%��*�.����뒘�{oÿ�}7Ի�'VZI���D�p�>�����X�\r&��6��d��[�5��ŕ��ے��J`n�i�K������"dj9�|�[�P8�V� T��lQ�
�!D/x�o�X�6Ձ��vl��,(ȲI)Z{빠\��0=�%0'\���%�y�x�V�0���L�F�ے��J`n�i�e�YQ�H1�����v��|��B��F�t�0=�$X�Yf�͎��8ꓦ;c���iK5���W<p���n�p��`n݃���t��S6ӮJ`n�i�H��rS �Eu�
DI�qh��s��h�h�ճ3�~�H�lŎ��D��$M���[�j��ջ6(J$ID!BIC���A��(I��[�`g�mX�&+j$�$�)�I�:�Z�h�`E�4����)^Qk
ˬ��`N�)��Ѧ]#Lm�L���8$��4,��&FI��9��{<�LS��FܪZ�F��Hj2�lb�{ނ:����$����-��s@��w4uڴ�j�=mk6~jd1d�j93@��i��)�:��F��)EDD�$r(�3@�]�@�v�'���.��s@�m��9������Y#����ݛ�͵`j��V�D1J��4�%N�z�<�fv�I>��:�#r(�LmŠw����[��s��`nV���P��8�S1.i�sT��p��mٙ�hx�zqe'Y�y�wk/%��[�}��1c��H�d�Ȝ΁�}�4uݛr�g�K���VqZO1T��r^b�ŕ��ے��J`n�i�����i���c�y�E�_;Sw�L�F�ے��R����2��,UY���U��Ɂ���r��ڴ[Z͟��Y$�L�5f��"^��?�]�`{ٶ�FH$�@����"F�	~P�e]
肐 "��"�`�b��!*�����[��@����k��ٌvn�դ��X���'lI��s)�n�r�S���t`�㮑��֨������v1	���;�_�>`×���=�}v3Zy�Ӯ5��P��L�����ogD�W�i]D^�T��I�x7O6�'g\Z46��kri��*m8�2o���)t�F40�c��qm���]d�
l'Bm��MZ޶
�p���&i�&����sy����=7��p���2�$M�5�V��{v�k�u�vAy�B.�(�����6�ń�f�Ȅ�}!�^ڰ9|�xO�q�7F܋@�v������3zՁ�{�Xz�f�=�NI�6�++Yw������H��rSk�h혱��H�d�Ȝ���u0=�%06\����U��ɁиT�5QLJdRf�λV���Z{빠{=n��ZC+_6�0ID�[9�]��'��鎰s܊��A�6�˝�M��1��X�&AF��p|��h�L]#Lm�L�)\+/*�e�k5�˹'�{�������*,)o]�6������ݤ�L�ڕn�Y$�L�._]��v��ڴ��s@=��"�7�9�$�4:""'����ή�=��V,ݵ`}Gn�l�ő1ȴ�j�>���Y��^�gZ�>�ǹfd�PT-�Cj���t&���:��#�εuBݬ�²W�#�X�!�e�I���?�&.����˒��+�f^��sM�5`b��W�BIL����?�Z{빠w��1��i91)�f�s�}�ܓϵ��s�: ��
��8P��}���gZ��iEl9M�k
ˬ��`l�)��Ѧ.��:�Z�Վ�q,���G!�w��05oF�ے�.J`!uR��ڣ������;2V�v˻6sj��Hz_l5\s���m�~���Y;���nz��]�S�Lm�Ll�07z4�7z��Eo"�7&H�h�h��=��V��m_%	(�=�/��*��k*�2�߳�����V�i��V�w�/"��F␙$Rfo�����+V�Z�>�ǹ�%��������_s�rO}�
k�3Y)3�y�x���Lm�Ll�07z4Ϳ��޹�']�������tFk������PV��k��d�q�ۧ<��]�b�$.b�ŕ��ے�ِ`n�i��z�hw�e�E�!��)���M�Qq	U�֬[�j��ջ6��U@ʬ��W��Y��07z4�ս`s�ՠs�S@���K�s!�$�nG1��z4��ܔ��̃�*����=�,���Ȥ�ɒ9�:�Z;f���j���m��DGDB��Ҫ��US��{9�n1���x�B�� 0�m��L��:���ks^K���麼��cxʚ�m��\Cvq�=�FiC`�cr�͜�;'G�l��nq���'=P㈬��i^lrͮ�:�V�n]{�K�a�ѧ;`M��˞��OCk.���ū.J�e��� Ο�'E�����7H�wE�f��H�m˦"jۓ���5<��<�X�{��Q{ ��OD�&��q�-�M:p�)��S�b�Ӣ�=I�;�N�����	��<jF�&�]��{Ѧ����rS �Eu�ʼ3Y�f�09oF�뒘��י�혲�$pXI�'�h�zڰ>�ݛ?D%>�|X�֬��'a�D�NI�̊L�9�j�9})�w�4��`�
�)^Qk
���s`}���9B���|�޵`}��6���y�wVF�c�m�ۉ�<�q	{O(;k�mDEr��p	ʹ^Z�ef`������i��)���M�ֳg�̆<�)&h��ڱD%�QJ�$�(��ٰ>�zX���{�Yq5�I�$s4u�L	�%3>�*�ލ0"�`{ee�O�q��L���|�Z{빠\���:�Z�་�)�E2cḿ�fڰ:.[�������ݛ�%�6ºU*��JeәmST�<�ڜ�nK3m�Z���.m���]�=k�<DK	2D�Ng �/�nh;l�/����٨;�]��tV�J4��ȤV��]�B��2v�t��֬Y�k@3���H��Jb�M�ڴ���7=�qI �� iq���#H&��D�$��j��3fn4�V�r$d�H1�Ќ�9jR�j,X@�S���+�$X��W �P� �  e�D4�h��Gh��`BA�)X�#�/���(�Ĩ��kK$�"� i�h�RT�0u!�@ ��   1C�G�!G�N��(�AR������'��~Q<�}=`��j�i3T߾��(��$�{���OgJ�C%�$�I���͇���o|�I���gA�y�{��B��k�]�6{��n
i��l�7N��r��W�
&C����&{k�l��\��C��{����ˣ��&Sl�B����&ӊ��&��]tu�v��$��9c�4jNr۪�T���	(��ߝ��I%����37�Y�)�[�j�䒟p���t�)�i�Զ�����!~�
���֬���f��{�������ퟜ�曗,��6�Jw{������/�=���IL��t��Ԯ���P�nk���k�9ou�脦C����B�}��#�C�@ Db�� !< �	��o8o�!l����d��sWY�kXe�7$�#|���I=���HfoZ��$�V��T��l��6+4���0�'�7:�BI�={C�s8��R���ͯ�����g�N*�?��po�����`}��/��֬�P�Ogs�gJ�C%�$�I��
����foZ���<��Հ{;�D%�mwM��$�y�9Tঘ�6��5`v�Z��IL���1$�|�(����37�_BQ!�ޕJG#bm�UUM��	{t�mwM��$�s7�X�ֹD%􇸮�8:
nZuE76DDOk�3z�(��ou��)�>�?�2"7���J��m�SӞ�y{v��P���sS���ّ��7lr�%�Nq�Y��V��e�7/C�kg�v��ը��t⨲�Z�q�qZ�2�&;\҄�lWF�v��U�Τ�z���ӌu��EK��,vR��{AN�0ݬ����q���T�^�`�ipF$���
��<p�u��giؚצ���³���u�m�&,��R��{��w}�����m�Ų�b��+��������t�ڒ�]����{52�7Ny0�n;�Emr��o��?Ͽ��;{�r�􇲻�B�O(�o�l�jWCcs(m74��W�d��`{+�z���6BS���3��y��̺�m���j��=��6�wOB��37�X|���,�(�')�)2]K���!L���6f��IG��֬.">Q��߾Z�|���pC�&5#�C�ħ3{�`owZ�Q􇲻��ޮ���M�?q�?�XkcnkOb�T���û>��k�s�]v�]s�L0�ԕr������nz�e�5a�BS���=��6t$�w��� ���g��I�����2��S.fkSZ�7$�/��{y�@i�D�Z,B����~�w$� }��9$�����Q�'�@̞����4��jMf\QḾ�+�龈�
d�޵`owZ脳�w���u~q�9�27��ѦI`{nJ`t�)��1R�HH�d�Ȝ�����v��ڴ��s@���u�3Md�r5�p�#Vmu�0$-ńn�ά�-�E��s/���
C�F���$��v����ލ07�4���R���U�Yy���L�w�L�0=�%09j�`��q��ӎ{빠w��f焊�>��8��g5Ϯ�{�},�ʕ�E4�T7S.��%
$��LV�lt�07z4�$�J�FF�)#crf�λV�����������s@�w4v֐���"dnLO����nJ�ɭ�#ja[��g�9��-Η�
۲����1����Z=e4��s@�w4uڴ��8������ލ=�䪊�0=�%0=� ��lŗ!�a&H����;�]��v����{빠sâ�ƢQ�$˵���ے��`n�i��I-Q�|�(��_yX��br�����e�S�2I%����{�4��ݫ@;O�>�B��,q�dd&.Ύ�Lg��\�ۅ[\+K��dv�-f�����H�ci��Y�w޻�:�Z-��<���2�#J9��i��)��2��0	�)_�fF�H��4uڴ[)���3�})�s޻�2�p� �$�lr-�d��`wti��)��/��Ȥ�8�4�Қ�빠s�ՠr�M���xے4��I��f��^�TV;8��]u9�n�V�)��W-=u���un��pd�g��,�i�8��G5-����WA�dhcfgG\�ka��`W$h��]�:ђT;N�����K3c*na�(Ҋ��[)�&�D8�f@v��f6idݻm�N0Q��(�oMmk5�S��d�� ݎ��#�c����,�7<e�0��֦������ �^y��.h�n]OB�F�ó�n��f�(pmsӎ��k]���G�
�8J������O�������ޭٰ>�z~I�J>���Ł�W`��9&7�I�:�[�~����߾|X���33mX���X��5LU�Yy�����d�`z�K`�c�A&29�������ղ[	�_}[S ���S^(cd�(�4{�s@��@岚{�M ���K$1ƙ��Ӎ��]���q5E{s��Vwj7<�nڣ�N��H��4uڴ[)�w���=�]��]�?Đl�B69��e/�BK^��r=o�}�j��ջ7��g�Ď���8�܉��)������jΈJg�]�`{��`{�ԭL�A�AȤ4{�s@�]�@岚~��޻�w��_A�5q���D��ܔ����d�`w]/���٠ڶ"s �����h�����8T�]��<���������w�tu��e�^exِ`n�A��Ѧ��Z�V;�"8 �Ldr{�M�J!L��֬ewM��[�`d�T�b)�*���t�`n�ڰ>�n͞�
#���V�;��ǥ�}���Ԅ��7&hn~����j�9]�@�})�[n�̮��H6H�F�"�-�)��})�$�0=�%0�t�_�Ҟ�l=u�c��LN�F:n�eX��h�!	s�K�n�k�KI.�̛�M����L	$i��)�%�Lي�P�āȠ�-�w7~��#�v��ڴ�����rD�N87�3�rSK���ҘH� ]�a�d&8b�G"�-v��~�rO��훓����(a
A �b@ 1"@ @`��#��"@�AH$# �6�@��ń�IeV#A���!��w��$��]"DpA"��-�~�@��~�n�λV�k�h^�
�$�#q�\�t�)��͖J�q�F%r9���-\�2Q���̆6HҒE�[n�λU��[��!%�eoM�{w�T:��:*�Vޭپ��"d��3+zlm��9�ۃ�I���Z�vlz�f�Ir�U=�j��Wt�-�YQ�86�p�@�_��-�s@�ջ6�$���M���J���̅70rG�m��:�Z�ՠw��l�@������4!+!6��|���\��K�0H�	#��@��� v�Z��M����Ռ�}R��!!$(|Ł�g�&�ā�1`�!הM	 �D�X@�_3P A;�Q�4a$`� � "#�����B��] Ěh0�1	B�ST�UHX`��dX"F$p �"�4	��#RQ#$GHB��֥�`��1`B)$�sl�B,�"���%V
E��!a��`nA�`YJR��(��'8CP�d�t@4�EX1�t��������:{�����o�  m�   �����  E;ev�g��mQ��ݛ�=O:%��3�EӐ��^Y��U/���,��� �]Kk�2�e��v�  [BA�Jmm�sm#�V�Iu]Xљ|��UҮƬcYz�mHí��ݞ�X�5+�4·<�ݎ��ܷn�J�s�7@�����6�[�ۀ��p�n֒��-��=bH��˶�r�wP=.�):x��S��	nѮD-��� x���pcy^������d��7]`F�ۄ#�'��iڸ����j�+m[[kn�o%�&����햨-j�S�\�ҳ��FKrLôv�vv1�ݕC���/),��Fx.�t��z��E��<F�貱�[`ظ�;hbuʻJ�*X���<u����;k�tV��MO	�%�ɞb��Z��� ����^z�����E4�gu�ngu�v�q��)�;T��u-Q�J��W��^&�nѝyY��j����ƙ	�uc 2�o�n۔��g&�bIm�6׭����x�)��ۛ+���Z5[ڪ����̽m��ў�������oag����8�L+�vi]0�ήQ�Vr��n����v�x�l�rٝ�dgtRD��OX�ct���mAą$��D��ƓZ�I"v�2D������+n+B��ָ��AX�8Uc�;$��1�&l=��Qv덠U���z�%�����	]�N����b�,��Em:��2U��Vc:6h�'gCƁ����3�ا]"<r��d��[�5��������52��]��v��J�Y�q�
��av7b ye�`V�V�L��N8 ���͡���tܑ�qR�ǥ�3D��lc�nq-b�گ)l[j��f�l��"Y���`�]v��V�T�R�y��;eU�\'E�x�4����Am�@   $.Z-�j��n�� !#rAoN�X�N��� �\�� T?�7τ���[r�At��\g)��u�4j�P: &�莢���`��D�Ǌ	��>t`�T6|95�{��ffd����yο�w�_+ۜ:I��iͺ�N�!�ภle�({u�8Z��S[�'G$��z��ӝ3ѱqۮ1����ݛ��9�D�<`6�TsĶ��kgM���c�qYdq�D�'#;�W[i.-ޯC��%�;LI4[��[�N��)��� �۬7S���,�Yu�R�P[l�����r�}�i%�XA�����a��K���˽����]O/]�������iF�Lmq�y��mΑ��݌�ko�9�̀��A��i��I3�{���	.J`n�J`I#Ln�ɂ�Xb�)u.��v�f�}TfV��wu��v� ���	�qh�͛wv՜�%>�������̩��cd�)$Z��hVנZ�Z��Z�z��$k	$�nL�=�%0'�)rSv�SI`����u=\�����e��N�<Ni�S����;�9np��7C���>�a�n���`IrSv�SI`{nJ`{ŕdF8��#�q���[���߸�$D	r�C'��X>� ��w�S&�*��*U7,��9�;��06��Ⱦ�*I�뒘��Qaj%q���L�:��@-�h�Xt%�������1�b�N];`IrS���4�ڒ[����o����,c��؉���N�O�#���*k���R)�8����*^Vq���ٰ̭7wmX�ݮ\�A�]�`}�k�9���Q8�[w4�v��ݛ2�f�"&M��r���m�Tڰ2{���ݛ5rP���dBJ<��wVzl��V�5�*�5C�WYy���rSw��4�UmȠ�eY�86��(�Zz�@5}��0=.J`t�)��؋�j��Xbbn9cK�8�kR]j3���f�̷V�S�D������p\sz��,�[����߿�rS��L��0'_���i�y$��s�ՠz�V���S@��s@3��,2(Lp��E�s��`n�A��UU�`{nJ`{�,���PqL�5"�;�Jh���λ�ܜF��;J�!g���p9mk�9���(�4��s@�]�@睫@�)�^��ZNdra"
I6Ks��g ݓi���V�K�ܜݬ�I�M�un�K�����������\�������+�4��&"�30Os"�E�s�տg�[>4[���;V��U+Ȍ��6I0mȴ���0=�%0=�%07f*W>�qb�"����;�]��v��v�����=�E� 8(�R&�I3@�V��
=��lfm�ٛj��Q� Y��B�z=����Z�ffffP[,���t//�k�h��NV��a�H;�Qvwk��]K)<t�q�ų�g�N��ƷUay���͕Vݷ]2h1��4up6��-� 7B5*<n�J��k�ϗ=q��2�]�\���՜�u�xg�ᅼ�jM�&��9�v���n����楞*n�h��ܡkr2q;1zؖ�]��Z���B�=������U����{��q���j�̳B���7���;�d$�3נwV��OE.�����9X�!	��QȾ����Z}빠{3mB��C�]�`{zS�S#�������=����(P�L��V����R\��s�%]�c�2�Q����$��^g8�K���+���ٵs�%�wCRIu�b��2C�H7&s�$��RIs���$��wCRIw޼�q$�v��� �8�E��I.zZ�Ē���jI.�י�$��=I%�nBnc�`�z� ���'u�f��O@��۶&I�9����3Ѻ�������wCRIw޼�q$�]��߳���f��$��"�ŋ�D�jI.�י�}�PLPD˖���5�m��;��[nf݅�D%	UT���W&�e:���9&s�$���=I%�KW8�^��I%�z�9Ē3����1�j9#Ԓ\��s�%�]�Ԓ]��3�I}���~�}��]�,cJ'����'"�K޻��$��~��o���$���G�$��j�I/�7靏��ۚ�S�f��KY�܉Ũ��s�XӚ�ٍD�ӦuxP�ݛ�˩W#��$��^g8�K���$�=-\�I{�t5$�]�,�$1�$�rg8�K���������g�.q$��t5$�}���Igl���	�G$z�K���r�}���M�������޾�xs�$����I.z��"2G�I0mȹĒ���jI.�י�$��=I}��g���w�8�Vȃ��E,r(9��$��^g8�K���$�=v��I{�t5$�׿��M�7�N����텹Vmu�u�Apݬ%f �r�\��!#���]vlȔM�g8�K���$�=v��I{�t5$�}���Hκ�XR!�j9#Ԓ\��s�31����K���s�$��RI.z�wQ<�FAIq$���K���s�$��RIs�i�$��fU؊i�i7UT�0��䒈�����-����5�m����9�oTC�4��
+���\���{�ʨt6*m�ES��$��=I%g�մ�K޻��$���/���興��
���Z�JL�UI�b�L38����3lЍ�k=���ubr
�0Vݗ�#���<rB(䏉$�~ߎq$���K���s�$��RIs=v�h�I<�nE�$��wCRIw޼�q$�]��I.zZ�Ē���,X�P�8�K���s�$��RIs���$��wCRI{��.Li�y$��$�����m�RIW�_8�^��I%�o3�I#:�Y`H�Q�$�RIy�_8�^��I%�o3�I$�l��K�߿oٿ���ݶ U�9^��h�:�
D�]S�&��^-:� �5�>��Qu����3o�v/�WkMq�I#Qc��v����n��\�Vn�Nf�';8�͞$\����P܆%�͒*s\���v���@�&��c��i3��9��6��[�a�WL�u����;N6�&�<u��&�;M�䛟��i�[�y�L�Yrj��jK�In�k}?!�G�y���e�zg[�Du�t���U˝q�V�4v�*�e��a�#�R�4�q��RK���jI/[y��I%�dԒK���$��Rɿ�2�H�r8�K��g9�߳i.�&��W��q$���K϶ŏ�d�9$�nL�I.�&��^��q$���K��g8�K�W��9x�Y��I%�l�K޻��$�m�s�$��RIs-��$pI�p��I{�t5$����q$�]��I%�l�K�33�7쭴��>N<��Ln�ܸ�]y�!���=rt�-�$j7
c�Mf�>���\�!#�9#�RI}���s�$��RI.�g8�^��I%�O��h�(Z+�? ��������?{ނB!BBLs5]�_}33��as33����Hκ�XR!�j9#Ԓ]v��$��wCRI{��9Ē]vǩ$�/�.6�dpr2I|�K��3�y�ԒV��9Ē]vǩ$��I*��?d1<����$��y��I.�cԒ]v��$��wCRI/v�X�ƖHc��nUe���8�e��tEQ^�磲��v���(��+4�s�ՙ�V��� �?~Τ�붾q$��~�����J߾�s�$�����D�9!G$z�K���Ē���jI/z�g8�K������6��.ٍ#�O#�q�%�]�Ԓ^���r�ڎ���cB%bD����bJ4��W�QE����	$f�)A��OT�*	�P�1 �����!5� B�@�<<�A��40@�I���!��"����Ő�H$X0�@M��_	��,bFH���)[Z���A_D��� ����N*|��6�!�� ���z�����M��ǂ��D$���R��v���ffr�6��fgwoPL�G,�(GI%�[��Iu���붾q$���Kޞ;�p��R&�Rg8�K���$�]��%�]�M�m�߾��[oED���gMj�m��ڻ8�w9��q��b�X+o�kBF�;<����'V�Q�q$�� �����K޻��$��y�333�i%�lz�K��K�������$��wCRI{��9Ē]vǩ$��I*��?��F�r�����s�$��RIv�W8�^��I%}=\X�Lr
9"mɜ�I.�cԒ]���$��wCR� 4������r�o�g�&���tk$"��RIv�W8�^��I%�[���f�{��?�R8�y&?�&s����&a��Q<�ηS��[��\
F��V{�l��'�������h�����4�j�;}*�(�ŒEㆁ�#LvL`l�)��2���ÄO�7"�4��h�զ���?b]��-���9�u��)!�4�aӜ�����Ł��j�=��`r�B�j7���ȜZ{e4���������������BJ�X$b��*H�$	Q�@H����D�P=����zАu�&���]Z�v����i"{RYQ�!�����a�4���є�����S��Ҡ��2���vqy��jt�]�nn�Qb6�m�8ݧ�2�C�k���-N��)��Bbu.�mv�����V��vC���.a�ݭx���iv���	r������n�;QvŴO?��g�����v'v���Z�MX	C.�dɣ�+no����}�Ӷ�1���杔2��!˻6[5�Z��r�oI�T�N[��D�Sm�/���i�nɌl�07fA��v�����rDۓ4��o~���s �ݙ�F�Ζ���ʫWy����1����07z4�7d�3�W��O#���;�)�n�i�nɌl�06vJXf^R�y��^^ލ0�1����;�d�7���Iǂ�%l\�v�m�F�nt��62;z���9�j���ͤ�r)3@;�f���M���{빠s:�X�)�䢊I�s�Y��� .�z���y���y��ٸ{l�9���[��H�Ԏ{rލ0�1����J?���$m���]�܀�@�_�9��@�_���A)$Q�3@;�1����07z4��_\�ve�yQv;XI%��RB�d'4ܒ���h���n�l^�{>�a�:j���̃vd�`�c�fKWC�<R!�!�w�S@�}w4��h��;}*�qǋ�G	���rI�}��Ep,A'@IJ��IG�9ϋ�ץ��V����D�r)3@;�f���M���{빠s:�X�)�䢊I�s�A��2�`�cr,�VE~�wVF�n݈:�n��n*#��.^Mt;=DƮ�
�ݒ`�IM�m�vA��#L�L`ñW.�S?m)#JHh���4��h���=�k��A)$Q�3@;d���L��`n�� ���A<i�G$��{����;�uXC����Q���Y�iT��2���E��Sgd�`�c�rS6�>���ι��17��s�I̫���d�m������J�[a�ͻ\�l󛣅���f^ލ0�1��)��%4��e�<jD܊L��٠{nJ`ñw�L-�t�#*��䢊I�s�ՠw�S@�}w4��h�Y(2'�H��R-���ލ0�1��)�+��L��0m)#Q�h��w���v��}�M�: @Ҩw���hֵ�&ffP���<{>���d�ohWg8�q<&�&�ce�S1E�&��#{g"Iב�u�7n�w*k�l&�����l��D:6�k��Z�N���Ÿ� &��G,�vhq֝V�jVю@��]�u1��ᮮ�v�]�-��ۂ����'�Y n4Y@�yݎ`�Sqn�ɑ�4�y�t.!ͻ9����|���C"�=�.��v� ��Wh��ʽo��޽��!>f`kj!51K�v�s���v����nG�R�!��r�&4�JH������F�� }}�4uڴ��h��v����&��t�6��[��&L�|X�֬��z3�W�ԉ�)�h��7z4�7d�Ԓ�;"�j�e�N��L��
w{�V���N�Շ(��}��}>L��F��29&h}��N�Ձ�k���ݵ`~QԲvzol[�+fa$M�{��N0�s�K�g���ժ!���N�n��;��z铟���7�"o ������ץ���k�G�gs�;�Y>D�dR!�G���M�?g�_�""�DG�*�w��`������_�bG�љ��HA���G!�[�ۚ��4�k�;�)�U�b��2dm�uM���3������ץ�,�����f�{�����m'y�@���X�"!gm���֬=����{o�*����+����9�R�Z��٪a�ᥳ���=���/a���ww�+�ɹ(W"&���ύ޷s@=�f��mzo�ŏ��Ǒ�(ㆁ�[��~��L��s�2{��{^�Т�;���25�9�8�h���@궽?~��K�
"��>ץ���j��z��V��S&�L�r۰����3�f��
&s;����O��42�ܕLt�����`~J"7{�_ fw;�����0V ���	�
�@���\�զ��"ֳlY�L��4�������Ff�ĄJH�r߾���٠u[^���M��?�d�4�7&X����Q	~���Tl�������`f[����0r��M�rM���{^�tDDL��Z���`|��iT�����[��S�Q��ξ,��[�O<��ܑUB��B.�G�������.,x��<��I4{vՁ�DB����=�V��K�^Ͳ���Yi&!˷
\i"��� \7G	YՎg�4�(��I��[6����� ��]���ڰ=�ztBI}!�ݹ�w<��ȓPN~J(��U���%�DBUF����;�~�`��Тd�U��dL��"�q����@��ܳ�(�&gs�2{���҅Wc&�m̺�X~�I)���Xgs�=;�V�""s:��:s�ʨ��eM6��6�vL`mI-��2�`O�/!#!H�5�~X�x�F@��&�fb`7Z4R��A�"ŀ���@�$�`��2(��@ڂn!�#�v��#E�:.� �HkZ��� ���ta�D`_�<F%<Ri��}���*H�}�U�HFI�� 0`+� @���"�P�� 4�$V� �$c�>䱅m���P
�% YJR�o�����8�`  �   -�m     I����5۴��3٧�1�j_U]l;e���q���@���;X��Ӳܼ �٫.��t��E���m���\$�R0һ5���m�O!�&a;���n��IG#����m��7Hd6ֱ@=��m��u�ԝ�Ą��q�,n�0�$��$�[v�E[G[@i-�m� ��gn��h"��vc�
qn��Ns�[ce��giV.�@k)���U��;	�u��Bc��q�[�fݨ���Zk8 Dklv�XV`�����1.R�ۨ9�M��n۰6݆@$-<
��&NP�غ�k�휦͹Hl&�b�8�ʣՃq��0Ep�㗀l6���$A�sM��vm�d�Zñ4i�T��W82��Uy�l,s�ո�y�:�bu� r݈iD�)���[p�g6yz��B��9�v��2�� �`&�#��tjk��3�䣮�ۄz8^��f�m`�:���AN�kT̼�E1�=!�KT�nIK UR���G=,ne˱wU\�[m�[a�ƫʴz��#ʒ���8�t��C킅�Ӟ�)��
�l��1L�v�wP+t�d�H���n�0�h��I�͙1�S�r��n��-�Pq��5+\ K���t���nvNc���t$�\��g$�v�%'AE���/
gP��\�8M�-����u�;9��y
3�#]]T� �R�����T�9�I%rd7a��nZi���s�=�a�(v3�<e��6Gf�ڝs������P.Ied�\ݵ�V��^UZ�
o`��X�W��c�}���+��*a6 I�ܶK����I���ώ)sWml]�����R��C�	z�뎌!-�L؞��=6� �����9��	:�T87�yu�-�JWO["�t]6��  m��U�3A�m�C6�rޮ�`&�q��A��,��Ҡ�\�:B�8�d�<�۱�m��yR�Ɗ�ҷ{����T4*��@ ���t�oJ)�����B��������wwz�/��j��1�nX8��\��([T� ��wL�[��Ƅ�K��M���(��m2�Nl�Ql�;���]�v������l6�BkWtv�ʖ�wM�V[x��T�l��%竱�����hLs�:Z�U=�JiV���b;Gm'U��t�n�mXk&͉#nrݞ����6D�Y�յ�%����`x������c<�؃�<3バ�fu�3nez\]���l��p��f���k=�z��������������|���ݙ�N&�9'���w�S@����!B�@��v�s�U"�nj���sT큻2�`�cjIo��*��Y�,x��<S$RG߾���٠s�S@�l���zQd�E27��Sn���9����s�����a�s7�f����c� ���䢊I�s�S@���`{ٶ���v��7��s?��X���k�Mv��8�ܹ�y�ն�B&&�KΔ�G���h�x�ͩ��!�����͵`��>��,���UL�t:l�=��W���Q�(��	\t%
:!%a�]��s�����}
!L�;��T:eS���6�3��{^�~���Ł��j�73eT��ʪ��5I�n��B����Ł�ϋ����������@�{��ƌjD��rL� ���� ݓِ`��~�����uv������]y�&ў��N���2��5��I��3�n��ۙP^ލ0�1��+���w��0=l�X�H7������٠s�ՠw�S@�}w7�#�����Aɉ���˙��y�s�rO<�>������R*��#�Q�%�{w�j�3ۮ��rSҥ9�)�ܕR幰�J'3��3~���٠s�ՠU��?Me�^`���� ݓے�� ͷ����p=��Ԗ��j���i��ۆ銵^=]疗����X`�ݘ�Y�2�/ ݓے�� ���� ��Xу�m���G$�9�j���|X�֬�ۮ�$�B�<��R�1�lN$�h���@�}w4�#�ﾚ|��h��<r<h����@��mX��]���vlJ%	��BP�����Ī��d�)�M�j�5l���ܔ�ݙ�F���}�߿N��PR�6�m��&.�2��k�E��9[@�.0<����g7hk��YX�3<���Lِ`n�i�j�3@9|�Ѭ�Œd�d�-����섔~QF�~�`���`}�ݛgT埉6�q��h��w;l���J&}��6v�,̙[b(i�N�n����]���vln=,:!DB�z�����,h��6�pO&9&�νٰ=���=��V�ۮ���З�D{�ww�����yZ���`�=���cN�;l�Y�s�\��ژ��ݖ�n��v�rՇ��
����Ć��ljy�!�N�����I�)�����U4l���+��u�tcbѶm���f�:	�Ԃ]r�6d
H�-��XK��2�mSe��u,l���{&�9,,elNaz2�đ�wF6�qMø����a�i.����n]n:g��~P|�3˙�.�FkS{p�l&zڤ�=�=5��&��BL��s�j��;l�,�1�lN$�t��Ɓ���h��_BP��ewM��\�R�6�������j�BQ!�;����;�)���3�G���"����I�˿~���L߾��p�7di�嶤�j��TҚ�	)�������;�w4��f�v�c�Y�$��ۛ�ץ��#3���,�vӻ��[c��8�'%0��x�l����$-��C��4����D��Z������]e��0[&0=RK�$�_�[�?����,��L�q�#�L��]�$�O�wj�����33m_L�n��F�m�ƞLrM��z{e4{�s@;��h��^4cR&؜J*�V������޵`�5�N�Ձ��q0�'&4HB4��=�]� �{�hVנr�V��\��k&)�@�é���v��]�L�АM��,���n=�Fym�n&����EwͶ���߷͏T���%0;�4�ߺ��,YW���L��n��kvo�I)��]�`n�Z�Y��"�2�*��s4�SM�N�9�=��6fm�9D%Q	e�|�I}
!I��݁�ٰ6qeJ�c*�s2���`��0=.Ja�$�]�}��>���0s#MG$�)3@=��K���%0;�4�ڄW*�V��-rj�`��H�cu��	�7R��S��� N�6	�/i�x��.Y����%0I1��Ѧ˺cvd�hƤM�H�$�h-�~���m�s@�oۚ+�o߿�/����rbDc�n���֬Y�j��kvl�ݚ��!��(�ĜnE&h|�[�3@�Wt�ۺ�?)�
�+Q�������3�N<R����ڴ�L`wti�˺4���J�g��
��-��O]�q��O7.�@�b�U5i瞢cWf�T��<�Ffc��~}�����Ѧ.�����:�L��0���˼��`wti�˺4���)�z�7����}�Y���B1I#qI�[�j��kvl�I%3���`n�Z�mYq9����s"�4?�~�|�
��Vfm��%�o|��}J�U.&ؤC�H�
�k�?�~������Z�>�ݛ��W:�T��mʳ�ƹ�O[5����sS�cIl�QˬsdJ(v�gV���Z�zv���)CZ�@��q��cl�^וb;\e.����h�bęS�,9���G:��� ���v嵶!����^*�vM
b�l����U�M�5Յvܔ��OJ��4��a�a���\���B�ƺLS�1�c9�ݴE�a-�`��4�;�n��{��˶O�^���17�tsv�ͻU&�N�{zV筗���N��>]^з.ң�����������;�)���q��|�[>H��&�'�I��͵�%2fs�����=��W�BG߫�>���!�<���=�Ɓ��-��#LS�L����u�W�f,������-��#LS�L?}�]�}��>��g��!Ғ<qǠ{ޭ05N�0=.J`ul����J�Yf��D<Q�'k3�1y�n�l4s��	�F�Ӭ�\���_��w>��{}$�F�(/���֬��f����~JK���Z�Y�!�167ndRf���M��"*h!Ћ�Z���5���nh�빠w�W�ԉ�jDLt��>ݫ�ݵgB�P�qv��1���;�.6qǉ�ܚ{n偋3mX�n͇D$�L�������J�ܹ�S4ꛖՁ�3mX�"Fc=�����mXJ򜭙��eS�7F��c��twf��Q�i'�ݴ���Eҗj������ww���g|��<V�z���o����[ �Ɍ�05oF�%+�4憛���� �ۮ���IBJ���ۚ�����mz�<�:a!ҍ�6۰33mX^͵g�<��(�"""���ňE! �#��� �Hā F#�,t��T�! E�� `���9P=CD	�T����ă������(�yK
@ѽ�Jđ��b�H�U߬������i(d�� Ō0�H����%���	 �@bA0��T�4MJB��
>) �<U� S@ x��_@�S�@�� zq�9���]���@���z`�A�I"�L�����D�����>��,��V�l��4�&��M̊L�8��@�����?,��~<w~�`y{6Ձ�n��UU5XM$���]Dh�o![v�5{z�즵�;��ʹ�m��y7%�F��������X���/f�䒈_Hz{���|�8�Ě�G����;����>�ݫ�k��B�
d���%CceR���̬�����LT��ِ`wtf䓏�٩�.SY��Ff�ܝ@�]�V��fm��+��
1(b�@��Ǽ��y�$<��fD��	$Z;e4����ٶ�z�f��Q;��%�&fB��S�J�F����e�Z���]����g:��:�=�߿~��4ֱ鄄�F�:���05oF��%0=� ��%Ҷ"�eQ-�-��/fھ�J�3+�l���w��h{V_Ɏbln4�țV�[�`}�zY�
"g3�Ձ�7�4�J���7�H��ȴv�h���ٶ�:""���6g>U@�]6�j\��L�=��V�Q�7�_�]�`}�zX
#Ud�:UT۪��{���u�ne6qmB�L���";pS��w5-�wu��U�6���9sqqhw[�ӭ�Y1vq1:��Ӷ��:6۪�6�<��G.�^ۺۢ���P\q�ة]��ݟ.z�5�]5��s[p�����ݹ�=bx��R�B.ۡ��q�vظ^̸� S�5Wnu�eg���	��[����VM�;<YS��`�,8��7n�V�ꙓZ���f��H�tuVδAp�%�PgO#��i�$rO����ٙ�wR�A<MƤRg �~���7nJ`{fA��#L�mqdW����R���x��%0=� �ݑ��������PCZ�������Me�4
�9�3?Ł�nڳ��,޵`fWt��eJ��ʢ[m�6X~�J)���Ɂ˧��%0=� ��%Ҷ"�e*���m��ٶ��P�f>�����@�m����E�!�i�֤:��Θ�t�GgAU�mg�Jsg�5հ�\��<<�ׇ7�E�+�m��������2�`jލ06vJWB/2�֮��3Y�rNy�}7��W�@w�@9��}��}��nh�h��aZ�L���������#L[Ѧ~�䒪Z}���;�J��L�	�n5"�4[Ѧ��Ll�0��_Ww��L���ϱ�Qc�bO$s4�ڴv�07di��z4�=��)�G�2�E�Q�pZR�3�j͓c�Jm˹�<�ͱ�Au.x#a�'?"8��dX�c�.�}>4�vՁ���_�">�̮�;hڕ\!���32�0`n��V�i��rS�������k�9�xԎ)$��O�07fA�|���̃vF�앱4SSTU:�����:'3���ϋ�ݵa�8�{�`gk�U")��UT���̦�d�`jލ0=.J{o���~��K�h���U���.���3F�3�4�8��R��1:577W��.�2rbQE��>������]��ڴv�h�T���F�FH���ٶ��L����]�`ffڿ�d2*�g��!�ły#��w���@�v�?DD����V�Z��nʦ�r��j�]fK���4���a�}��Q�;� 6��}�y7$��OZ���EZ{n����e�~�p{��r�V�w�r��8���4um�p�]-�����y�q��R��]��+��Y!��5#�I3@�{�s@�l�������В�Pn��j�;�J�E5USW�Wx��vd�%07di�˳m_�:��;k�T�����&��`{���`n�,V�4��� ��qUʫʒbQE#�h��޻�{e4>���ߧ�-�υ�!��H���˺4�ݙ��L�`g�.�ww~������j��c�۶��ٳ�`��m4J���Lp�u�$Ӕ�Mm3�ex�mu��!�r��cmTg��uFְv��9gl��]����5l�#�9��WM��1�:�ÑIl�B�F3��=����T�`p�K���+�'�#�9�������c��.��{ؘ����7];=�.��=�S��vy+\L�1�d�Ӄ{=����{����|��ڴ�:�g�:�6';O=�-m�E�pv,U�1�:0�n������|N�qc��G3�_}>4Wj�;�`r�0�IJ�Y��+1X+����rSvF���Lِ�_}T}YZ���EZ��ۚ���V~�����Ł��3wjUX��R)�r�já%�!%\��yX�����v���s@=��Lsi��s%f&�IlK���`r�0��{>>��3��n9�^cPv.�h�u�3��BOF���k��[��{���ɻL��
ŗ�^_���ݑ�.��uڴ�q:'$���)�@�mܿGBJ����X���ٰ3wmJy�i��d�L�=����8��@�v��������Yq�A�<�V�ID~P�^��V~�ߦ���mX��s@3ǭX�2,qI�"�M�ڬ�~K�w�/˻�� �n�w]I'�{n��Fr�L��q�eܐ�5�5�*�ɞ��
��M���N�M�l��09wF��1��rS�mJ��sH���m�fھ�!���uwM���j�36V��MUT��6Kj�7ۮ��+vl��ϡDJ�(6�.��  0D�ARB*�E�TO@������rO����Ҭh�9��N
'$�<��0;��06�K`v�Up����Ku,�鹰3۶�В��G.��^�}?��ڴwхx�LiQ&�n�<\�n��]��=�6N�l��1��ۋ�[vd�<�R4�"�4g�w4�=,��g�_HnwZ����\��8�O$s4��Wj�=�w4Y�j�L��{�ST�U9�nlg>,��?BQ
goZ�3�zl�X�:a!�H�nC@�m��;����O>׿]��W�PM  ~[�~��_��Ǧ$O"�I3@�w�s@�})��l�0=P�
ŕuYJ-\�`����ul�9��^&�z4�n'�l1ׇ7.V��+�m��_ݛ�k���n��J}!�7�X��q��7�ȉ���v�h���mX�ͫ�
S'er��i�کn�
�/�ߚ`jލ06�K`{fi`ffڕI�[�����Շ脔)ś�+:���������%
w;�V��U��D��<���;_��9�)`g�mX^͵`B[Ȋ��>����$P��YtK�$��$�%�İچ���Dj�$�R��@��a�1(@>6�v#�.��[@􊆂��!��im@��Cb� "a�L""��*�` Ia%(%
H0 �B4�޾���ޝ===��>q��      �6�    In���m�6���w9�ki4�le���U^���4�G���흶^�FH졉�(�PK A�&�j�I�f$�L�W�M���.▤����;�Q�����nV���ڲ#�Y]P �í��[n�MF��K<E��_��6����m��
ۛ]+gm[��kn *9-Wt8FҚjƞu c)���Ҏ�1�\��a�eV�H���+UHp��y�Y�2f!�W��$�K�Ss�vsXkZ\Ӓt�n�Am�1&��|�����X�r�T��ӡ��86�ɺw&Z�K�.M�r�p�IY�m0�<KX���m�gq�ܝUɭpݍڬ5�R.+v�1���W�,g���W��9%4x�\��k�\���z�R�U/�vsp��pT�]���N�N�z�':{h1fu
F�؞ݪ@����s���F�mV�m�8zM.���e(6[=��[kq��f��q��<J$vQh�]&`R��T�\p�P2��W����YQ.�4;vYu2�qnX(ڍ��QK=[>��MM���J�+8�q:�L��[r�@�V���FtɌε-N��n;R��Yݬ�-�,�`knX�K/Iҗ�n������z]����G9�!:��j�쬶5���A��0Nڎ6�a�K�0nܼ��Ĭp���ড়f�i:���b�5v���h�'N���m#Nrʙ�m�j�P*"@�l5۰�gM@B6��C�m�C�iH�5m;�Հ6�"��mW@驶x�yuڡؚ���ܨN�u�xհ!5����vc7kݖ�lN�m�^�z�N��o`�c��!�YuIg3�C��	!�R�����X��a5oB�q�%F� ������q[GF(f�� m�@�67j:�0��pl�U����
��n���f��Iֹ���I�����s�]!�V���Q�1U�C2�WV�x��N
�P>P��@� ��	 > M(�؀mU(�I�@�‟*�� ؈<UҢP`�r�EAК������}Ks35nk33&��)��G�Õ�M�L͈l�m;5
I����W���Z�zL�A�p���Id�qw&��.:t�qr�	�89uvlۃl�khܑą�]5����[mҝv�����l�N��ܦ�q�{9�vp�X3�mv����n:d�v0��$v�������k�ê�㗞k>|��ϵ�c-����Y.�:$����OЁ�峓��dѓ2j�k:AD��m��ض��5k:�c7�)+�g���٣֤X�"C����$^�����۹�u{6��~JK������<��W����̻��4�ս`l��k��!%&wuJ��sH���m��O�06vA��l�0�J~Lsr(�E&h���9�)�{۶�9$�N,��X��QP:j�U7&+����oF���L	�%0;�p�&&L�LqG10s"M$�I�2tIZ t�l��m�1jW#�Wi��=�{����]�bR5��>�}��w;빠s�S��fq}���=oۋB)��H�nI��l�A��,�lA
 �ϫ�Ł��K�͵��2���\���/-U���������d�`nw�s@3�mX�8!��0jH�v�,��V��mXtDNWwU�ӫjU|E	��H܆��[��w;빠u[^���M����@�!, �J
����ӝ�Z��{��z�uu��K$�Q��zlֱ���Ȣ�L��_�4�k�9�)�{��h{V_ɒ���YY���$��d�4�ս~���ϖ4a��#�=��|l��~�f�~	 J��A�T�$��������V���z�����N5�{��h���h픰��B��B��������֥Rc�ʥM�fe�`jލ0=� ��̃w�Z�w�G�L��2"4т����!f�K�3v�;�m;]Q��r��w��}�ל[�SY�0�0䓁��fӑ,K����iȖ%�b{������Ț�bX�w��"X�%�NϿ~���K5�X���˴�Kı<����r%�bX�}���r%�bX����ND�,K��{v���%�bw_j��3-Ʉ�˙�fM�"X�%�����"X�%������Kı=�w�iȖ%�by��nӑ,K��Ba�tMf\���iȖ%�b|}�xm9ı,O=��6��bX�'����9İ:��%A2'���m9ı�{���mͩp��]������,O=��6��bX�'����9ı,O}��6��bX�'��w�ӑ,C{���~���t�\a4�W=u�U��df��N8�Z��\"��m����ƴffI��̻ND�,K��{v��bX�'�w�6��bX�'��w��D�,K��{v��bX�'��}.�u��.�ܗ3Y�iȖ%�b}�{�i�~��j%�ӽ��iȖ%�b{����ND�,K��{v����&�j%��{��M2�Mh�fI���iȖ%�bt�p�r%�bX�{��m9��D�Og��iȖ%�b}�p�r%�bX������2ܚ��0��ND�,���O~���iȖ%�b{�?~�ND�,K�~��"X��'��w�ӑ,Kħ�����Y,�]f�\ɴ�Kı<�w�iȖ%�a�R?}��O"X�%�ӽ��iȖ%�b{��nӑ,K����
����t��=>�?/���.����j�7+�=�nTЬN����Z��tnC2�8�v��i��۶��H����ݲ�g��3�;뵷4�r�Vԛۻ6�8Ρ�lE��]/-��Ԙ�#f;��]#kI�9eG!�Zێ<��5΀�s�`7�im��6�]#���G="�)˻tv�\򳭵ñx
d��7`���<���{�Ѕ@NפȪ��$ɦt��������c<�7 l�-�V�))e�ö�G\�T�I��U�4e�F�xrL�rd��u���_��,K�������Kı>>��6��bX�'��}� ND�,K��{v��bX�'��uMrˢk2��fND�,K���iȖ%�by�wٴ�Kı<�w�iȖ%�b{����Kı/�v�sY2�V�Y����iȖ%�by�wٴ�Kı<�w�iȖ*�b{����Kı>>��6��bX�'��ԝfkh�fI��s&ӑ,K���ݧ"X�%��w�ӑ,K������r%�bby�wٴ�Kı=;��]3Z�Rk2乚̻ND�,K�~��"X�%��=;��O"X�%��߷�m9ı,O;���r%�bX�׽�&L��uLɭe˖fn9r��4RHl��t�K���%�B��Z9*��FL��Z5��ff��r%�bX�}�ND�,K�{�ͧ"X�%��s��Uyı,O}��6��bX�%����֮5�SY�0�0�r%�bX�{��m9��x�����q7���~�v��bX�'���ND�,Kύ����$)!I
V��*i�JsN�-\ɴ�Kı<�>��r%�bX���xm9��,O>>��"X�%���fӑ,K���֛�3-ɒfeֳWYv��bX�'���ND�,KϏ��iȖ%�by�wٴ�Kı<�>��r%�bX�w��5�L3.��˗5�m9ı,O>>��"X�%� y�wٴ�Kı<�>��r%�bX���xm9ı,K����h�չ�����-����8G�n�a��g�Jsg��V��[
#��uG^�B��Z��r%�bX�{��m9ı,O>ϻv��bX�'���ND�,KϏ��iȖ%�by�}I�f�։���&\ɴ�Kı<�>��r��
j&�X�}��6��bX�'�;��ӑ,K����iȖ%�bt���t�k5I�˒�k2�9ı,O}��6��bX�'�w�ӑ,`�Č\@~A} �'A��K���M�"X�%��s�nӑ,K����&��s&�k5���a��K�D,O>>�6��bX�'��}�ND�,Kϳ�ݧ"X�%��w�ӑ,Kľ�w]���&�T�hɅ��r%�bX�{��m9ı,O>ϻv��bX�'���ND�,KϏ�ͧ"X�%�}����.��4]q�1��K8��^�spyE���Gb�ʬ�]!߮��w�&};8�e�:k��i�Kı=�w��r%�bX�}���r%�bX�|}�m9ı,O{���r%�bX�w�M��2��5�uu�s.ӑ,K�����Ӑ�Dh�/j�p�P�Bή�H"B�3Zn'�@T�K��֟�	�eԚֳ̺5�ӑ,K���siȖ%�b{��nӑ,K�����iȖ%�b}�{�iȖ%�b_��:�˖�kY���36��bY�P���'߷���r%�bX�����iȖ%�b}�{�iȖ%��z(� ����Mt�<6��bX�'�gԝfkh˘\̙�v��bX�'���6��bX�'�w�6��bX�'�w�ӑ,K����ݧ"X�%��_}���S3.OC�v���񛳧+6�H��cNӎ��U�f"3�m�Y\s�]���s�Ϻ�M���J��'�,K��~��Kı>���6��bX�'��{��"X�%��{�ͧ"X�%��{�Y4d˙.��XL��ND�,K�iȖ%�b{����r%�bX�w���r%�bX�}���r�X�%�|��]���&�T�hɅ�6��bX�'��{��"X�%��{�ͧ"X�%�����"X�%!b�����$)!I
V��*i�JsY�Mf�5��Kı<����r%�bX�}���r%�bX����ND�,D��]�u��Kı;�֛�ɓ$�e��\�M�"X�%�����"X�%������Kı<�;۴�Kı<����r%�bX�����s\�UU���胳��񐶙�ti�uNX^�6ND����[4r*;2�Q.�&�+�s�:�>�dn2�.�ܗN0된��-����oS�-<>�c�R�2r�P��X����tm����pݦN{%Vm�Rm��C���ܽ/�۵۬�;'���� �k��nS3�j�컮/Rqks�)��59�k-�ܭg�.�	�zrv �ے0��{�����C�m�M��u3�u��GM�HK�LtԵ��s�JgO�4S��)
����v��f����ؖ%�b|{��6��bX�'��{v��bX�'��}�W�,K��߻�iȖ%�b_}�:�˗Z�Z̷0�fND�,K��{v��bX�'��}�ND�,K��ND�,K�7�W����$/c�G@骤:e6�f]�"X�%���fӑ,K�����ӑ,Uı==��6��bX�'����9ı,ON��٦�Y�Mf\�&k&ӑ,K�����ӑ,K������r%�bX��;۴�Kı<����r%�bX�w��FL���k5���a��Kı==��6��bX��@� ���]��,K�����6��bX�'�w�6��bX�'~���C]��h��k<�ܹ���,b)Z�ķW����c�4an�6�r�gY���%�6��bX�'����9ı,O=��6��bX�'�w�6��bX�'��w�ӑ,Kį���,�]f�.��˴�Kı<����rڨ�Ih�� �h���J�/� ؛�bk���"X�%��߻�iȖ%�by�wٴ�O�ꦢX��;O�f�dԚ̺�˚ɴ�Kı>���m9ı,OO~��"X�%��s��ND�,K�{�ͧ"X�%��{�S��ɓRk2���"X�*-������Kı<����r%�bX�{��m9ı,O}��6��bX�%=���s.]j�Y�.��iȖ%�by�wٴ�Kı<����r%�bX���xm9ı,OO~��"X�%?b�ď"q�l�0A��1��,��wSv�M�'v)x3pr�]Z�{�ދ����5�Y�3Yv��bX�'��}�ND�,K�~��"X�%������Kı<�;۴�Kı=;��f��f����.�k&ӑ,K��߻�iȖ%�bz{�xm9ı,O=���9ı,O=��6��%�b{���FL���k5������Kı==��6��bX�'��{v��c��8$4h�j:*@* �/���LҮ	-
"������$X��YHłԀQHF5RR$FVP�t�0H�-�t(h@��X1`�`�"�8�Ib�h
V!YYv�WKhE���eap��Û�l4A�HA!+)���e`��	H���ee&�WD�2�՗:�-H���x�!�Z�>V��� v���pDM����@CJ"p��:X����o��Kı/{��ӑ,Kľv}��N�S(�Hmڸ_��$)!{u�r%�bX�{��m9ı,K�w6��bX6'��w�ӑ,KĿO��5�2٬��B�e�r%�bX�{��m9ı,K�w6��bX�'��w�ӑ,K����nӑ,K����?����9�ӭ�srJ�Av�v��AC:�uAÞT�V��v��/g�D�b�.e�yı,K����ND�,K���iȖ%�by�w�a�E yQ,K�����r%�bX��m7���&���55����Kı>>��6��bX�'��{v��bX�'����9ı,K�w6��bX�%>���s.]j�fd�5u�ӑ,K����nӑ,K���ݧ"X�%�}���ӑ,K������r%�bX�{�Ru��5�.�\ə��ND�,� ��Oo���Kı/�w�m9ı,O����"X��!�OQ��}�s�iȖ%�b|{��f��f����.�Y�iȖ%�b{����Kı>>��6��bX�'��{v��bX�'����9=���ow��ߏo�c�1pL���s�� �]v�ŉ�wH���#(���\�^�F�2e̷WY�&fk�"X�%������Kı<�;۴�Kı<�w�iȖ%�b{����Kı/���f���k-5rL�k0�r%�bX�����&�X���߮ӑ,K��~��Kı>>��6��bX�%=���re�Yu�����kiȖ%�by��nӑ,K�����ӑ,K������r%�bX�{���r%�bX��}N��r3&��.e�r%�bX���xm9ı,O����"X�%���ݧ"X�%��s��ND�,Kﾴ�Y�2h��3Z��ND�,K���iȖ%�a�@B>��߮�Ȗ%�b{�?~�ND�,K�~��"X�%�� ��U�`@��w�w���;��v�kX���nv�5���fr�H��Ůev��M�2I�&s�=�bt�����;���]�7!�ɍ�����8v�vDun��6��m�����F�sn�l�b��vr,��X��d�u�<`��J�(��\pV�7J�ru�Z�Y�۳s��1�#�a�����\"{!���nm�׶�;Vx��c8�IջX3Z/�h��: ��l乓Z��E�k�#l��8V�T.j�N&�z4��V�F#C�c�B�VF���{��%������r%�bX�w;۴�Kı=����r%�bX�}�ND�,K�s�N�5��3Z�s&f��9ı,O;���r%�bX���xm9ı,O����"X�%����iȖ%�bzw���7Z�S3Yr]f�.ӑ,K�����ӑ,K������r%�bX���bX�'����9ı,N����s-��k	���iȖ%�b|}�xm9ı,O=���9ı,O;���r%�bX���xm9ı,K�gu٭a���M\�0��6��bX�'��{v��bX�'����9ı,O}��6��bX�'��w�ӑ,K��V���2S&d��ja�E��ɺ��[W��Y�#{N|-��H�ڻW[���d�f��5	f�2�9ı,O;���r%�bX���xm9ı,O����"X�%���ݧ"X�%�ߧ���fB�d��e̻ND�,K�~��!P�D���M:��,O����"X�%����u��Kı<�w�iȖ%�bw��T�3Xdԙ�5sY�ӑ,K������r%�bX���c�Xj&�{�?~�ND�,K����ӑ,Kħ�v�ne�uf�2]��iȖ%�b{����r%�bX�w;۴�Kı>����Kı>>��6��bX�'��ԝfk54f���f\�m9ı,O;���r%�bX�}���r%�bX�}�ND�,K�w��ӑ,K����������(]B�m۵�� t�����\�L��9vn�3�d�b�4|�~D�,K��ND�,K���iȖ%�b{����~UByQ,K�����r%�bX��~��&:�2�]fd���6��bX�'��w�Ӑ�(D�K�~��[ND�,K�����r%�bX�}���r%�bX����Z�S5���&a5�m9ı,Ou��[ND�,K��{v��c�S��9�5���m9ı,O�����JB���wxM�̔�l���|B��%��s��ND�,K��ND�,K���iȖ%�b{����r%�bX��}N�0�\̚�̹�iȖ%�b}�{�iȖ%�`�}�xm9ı,O=���9ı,O;���r%�bX����K����.�R�d̚$,��z�4�����;�����ǥ�D9�WM���n��YZn��7���{����{��ӑ,K����nӑ,K���ݧ"X�%��w�ӑ,Kħ�v�ne�uus2\5u�ӑ,K����nӐlK���ݧ"X�%��w�ӑ,K������r%�bX�{�Ru����sY5�35�iȖ%�by��nӑ,K��߻�iȖ%�b|}�xm9ı,O=���9ı,ON��٦�Y�fk.K��e�r%�g��������Kı:w��m9ı,K��m9İ=<*�D�����nӑ,K����
c�3-�ֳ,��a��Kı>>��6��bX��:��߳i�Kı=���]�"X�%��w�ӑ,K��G�}���tՖ�udPش��6���	\=Q����-p���a���s|ߝ��~?3Y�j䙄�a��%�bX�����"X�%��s��ND�,KϾ��"X�%������Kı/�}�fd�f��5	�k3[ND�,K��{v��bX�'�}�ND�,K���iȖ%�by���bX�'~�S�fL23&��.e�r%�bX�}�xm9ı,O����"X� j&�{������bX�'�����Kı=��M���&��˚�f��r%�bX�}�ND�,K�}�u��Kı<�w�iȖ%�by����Kı)�ݧ[�r�]\̗]a��Kı<��w[ND�,K��{v��bX�'�}�ND�,K���iȖ%�g���{�=��������O+V�U#=P�vo:n�^y�]Vz��
�닮sPv�R�W���[%�:;F��A�֨ ��ܵ��	��p������`!���6�0tq]���q�9'qy)�S��@Gf�ۯQb:�\�ڮc=���sV�B6�<ب�S�0��1�[\qugm:�H��Ōk�^-�4;O&���H��[H0���Us��C���4c�S� D��]nٚ�ְ��$���]Da��mR	�����;l!k����W���i�{L牲ܴ��w������Ͽ�iȖ%�by����Kı>>��6��bX�'����iȖ%�bz����f���f��k5�v��bX�'�}�NE�,K���iȖ%�by���bX�'����9ı,O}��)�d̗SZ̳35�ӑ,K������r%�bX�kﻭ�"X�%��s��ND�,KϾ��$)!I
HY�_�C�2�T��W�,K��_}�m9ı,O;���r%�bX�}�xm9İQ�>>��6��bX�%���]ɖ�e�j�3[ND�,K��{v��bX�'�}�ND�,K���iȖ%�by���bX�%��gԚ�L���%34aӪ�!��y��t��*��i�֪�v�-fƜ�o�9:��)~�~���u��=�}�xm9ı,O����"X�%����؃Ȗ%�by��nӑ,K��߭7�k��Y�Z�f��r%�bX�}�NB!�C�x�&�X������Kı;�~��r%�bX�}�xm9ı,J}�i���e�us2\5u�ӑ,K���ͧ"X�%��s��ND�Q,KϾ��"X�%�������$)!I��Q�:tT������ND�,�(5�����9ı,O{��6��bX�'��w�ӑ,K�����ND�,K���ηZ�S3SS3&�.ӑ,K��߻�iȖ%�b|}�xm9ı,O=�y��Kı<�w�iȖ%�bw^�������+,E�nT8V��奖vB�XK�c{s�W�DW�}����Ϻ��-��A����=�%�b|}�xm9ı,O=�y��Kı<�w�a� �$��wpI,�өt�Rs@�)�j(A�>�q;ı<�w�iȖ%�b{����Kı>>��6��%�bX��{w&[5�Y�K�33iȖ%�by��nӑ,K��߻�iȖ>(!�R*1D�>(� �p�<�ӿs�ӑ,Kľ��siȖ%�bw��7�L�d.fM]f\˴�Kı=����r%�bX�}�ND�,K��{�ND�,U�<�w�iȖ%�b}�֛�5�MY�5��a��Kı>>��6��bX�%���6��bX�'����9ı,O}��6��bX�������28)8l[rXE�It�u$��t�d�ې���r1��Ru�L\���.��iȖ%�b_=�siȖ%�by��nӑ,K��߻�iȖ%�b|}�xm9ı,O=ϩ:��jj��L�jf�6��bX�'����9Kı=����r%�bX�}�ND�,K��{�ND�,K���ηZ�L̚��5�v��bX�'���ND�,K���iȖ%�b_=�siȖ%�by��nӑ,K����\33WV�3R�]a��K�[���iȖ%�b_=�siȖ%�by��nӑ,K��T�Ck������j��$)!I�����Rs@�)�iȖ%�b_=�siȖ%�by��nӑ,K��߻�iȖ%�b|}�xm9ı,O~~��kW���̶L�,\�a3q,���z����7<ݱ��@Mų�ōfL�k.�P��s36��bX�'����9ı,O}��6��bX�'��w��yı,K��m9ı,N���5�L�d.fM\�f]�"X�%��w�ӑ,K������r%�bX��{��r%�bX�w;۴�Kı7ve_AM2�M˪n��_��$)!i����Kı/�����Kı<�w�iȖ%�b{����Kı)�ݧK�5�����p��ND�,K��{�ND�,K��{v��bX�'���ND�,K���iȖ%!I��Q�:tT����黅�
HS���ݧ"X�%��w�ӑ,K������r%�bX��{��r%�bX�!�H�#`@�U�z��£7=�Gn�!H4�
,
0
,(Ʃ(��E�JU�0`�H8	�_5�<Sˮ!�I��t	�L�
�V� z�Ŕ h`��*�ƩK@��� �e��#t��%B"@!�Ul
,X��H�+Ѧ�@�@#��F%*H�"B���iE"���]d2Ձ*��{������       ٵ�    ݐK��٬�f��ͭ�{c��n��.Em���1�l��@"t�9��t T�wi�۲Χ��m[�HH�6��'Uһ^g=+�l�h�l��Kv��h�`N<������\�˵:s���W�lq;��I{t/�Hŷԑ;��
b$q-Ʀ���Y@j���g�j�v�m�Z��8���68�s�	��U��8N$إ����VV�����6ݎ$���^�cW�b6���z�uO.ݐ���p�j���j�+Nʤ��-\��-��U��V�,�W��)r���t���r p�-C�ɕ 689���Ю�\��n�9�(��d���ئ��m��p���%��ܲ����-g�Z�U���A�K˫vV�n�F�����S�5�n��U=�u��5�B�%��:�p:7vܫvm˖�˽r��%��8YbI7^!�nsNĜc[�5X�{�D�=G�9���.�HJu8���D�U��v�
�Wvm����/�f�8�H�!=@*�U+���g�U�V�x�S�nޮ۰��%97�&$Uf
�lV����pءBіUV�P�G%Eu-�%+������Kp#��l�5�݅N�r�gs7@.������3�ukZB{u�vݩuaS{m[\�8�nH�{<vږϳ�Wv[����v��U��sC�l�y,�3m���[2��{Z�L�rɺK��Al�9��%���`Ii�$��]]q���*COT�G����VE쮚URLf:��W`,�sL��0qc�q�D�nN\H��*�;(lhN�ҳF�'��cj4��I���{�>{�7Ov��2�m+qX�a7մ��n�{r:�Ύ�#�pn�G	:ഀw�nO�K;o��YЏIt/iy��#�ݻn];V���\��`ٷi  m� H&ʚ�֛Z�m�N�l ��&�r޷����Y�8�3B]�mP�)Mr:��8� ��t���IrۣV��V�Z�\�˥W��*����=U~�C�< "5����������ۻ���M~�7m� �v���8'���D���KֳL�4�6)��3��[�b�7K�ڼ��Yº�=n:�mn6�ɤa��N���u�9xv����Ӽ�74\��Uu��ҍ���dy9����9�����=,�m�M��zc�k-�bxIN�q�0񛒸����fP��Y]��.:)�ka6M�^��kTMd��h��zd�����{��}������2uϴS��]��n<�ˋ��t,m�CL�p�)R�fҸ�������o��֍d32jk2�2�;ı,O����"X�%������Kı/�����Kı<�w�iȖ%�b{�vS�I����Y��2��"X�%������?�GQ5ľ���m9ı,Og��iȖ%�b{����O�D�MD�>�?o�ֱ�j�e�3	��iȖ%�b_~��6��bX�'����9�� ��MD�����Kı:w��m9ı,J{�a�t�Me�j�s36��bX�'����9ı,O}��6��bX�'��w�ӑ,K�/�����Kı;����a��!s2j�2�9ı,O}��6��bX����xm<�bX�%��߳iȖ%�by��nӑ,Kľ��N�XM\�S;7/12΁E�驜����Ο8h���GB���A���g�D�������K������r%�bX��{��r%�bX�w;۴�Kı=����r%�bX���ݦ.k-˫���a��Kı/�����?
����yQ,M}��ӑ,K���~��Kı==�xm9�:���=������i��6Y�_=ߛ�oq����߷�m9ı,O}��6��bX�'����"X�%�|��ͧ"X�%���}g]h�C3&�dˬ�ND�,��Q>���6��bX�'�߿p�r%�bX��{��r%�bX����m9ı,O}��t�33WV�f��.��r%�bX����6��bX�%���6��bX�'��}�ND�,K߾��"Y�7���~��g�� ��fU��
��hn�ʵ��[k���[^�<h��a�\6[ͫ�S5��k0�r%�bX�ϻ��r%�bX����m9ı,O~��6��bX�'����"X�%�O��5��)���B\.ffӑ,K����iȖ%�b{����Kı==�xm9ı,K���m9ı,N�>��	���ɫ����ND�,K߾��"X�%���{�iȖ=��!�+- <@�C�'�/����r%�bX����m9ı,O����k�&�.[��ӑ,K?Q>>���iȖ%�b_{��m9ı,O;���r%�bX���xm9ı,K�����5���ɢ�Xm9ı,K���m9ı,?,}��߮�Ȗ%�b}����Kı>>��6��bX�%��>���:��z];v6᱑.)e�ݩ��ڌT������N�#����al�3Y�ND�,K��{v��bX�'�}�ND�,K���iȖ%�b_>�siȖ%�bz��Y�Z��fd֮f��v��bX�'�}�NC� �MD�:w��m9ı,K�~ͧ"X�%��s��ND�,K�{��2L��չ�����6��bX�'��w�ӑ,Kľ}��ӑ,[���ݧ"X�%���w�ӑ,K�����ֱ�j���k$�Z�6��bY�A������fӑ,K���~�v��bX�'�}�ND�, x
��tz<�'�3ND�,K�����%5�Y�K����r%�bX�w;۴�KĒ#7{�p��5n�� ��;r�I3�m��Y�nH6D�x���X�,DvSe�-�*��p[�飓�����`r�0t����)��K�n
i����mX�6��J�os�;���w޻���K~Y ���5MX���mn͟�"��޵`\����~X_�q4F�$drh��`oti�˺4�=�c~��'�vE�A�#r-����?��s8���@�l������g�g����nI$�ID�ei4��'V� Ł&��:LH���]%�Np�V�u�Wc�X�ol'/]��nը�j���O��l�8wl�ݎ�s�c�ۓN]�=T�V����ʤ�V��J�E �a�Լ��ϟ>o��0ݬ��R�<=v�ۋ98�Y��#m۷.m��#
<ڤ����k������t끠靦2�u��[�2�l��D���Mf�޵)���0W'72g��A���{7%��wH�c�灐C���d��k#�u�L�蘭����L�&0=.J`oti������Q27crf�s���;���z��09wF�킻�
W�yb+ff0=.J`oti�˺4�=�cwU(�]b�VfW�Y������ti�w��C�ߧ�-���l�9�a$S109wF��L`z\�����k�����$rZ���*�#J)@�.j�N&�t ��칌�����+��*���7zc���F���Z<�����h��Hڒh�տ��ߔB؄�����Z�9w~�`�k�=�E��"� ڑ���۹�{=빠��9]�@��F�RF8G���O�L�~���Ll�06Q����dn��� �}f���Ll�09wF�U�
\��)a�]3r�S�����u�S�$:^Ӟ�a�-�Y����C"���0RM�ڴv�V,͵����ߝ���e~�T�LSY���Ve0=�4���`�1��rS{��y�x��fa�Y����L�y�f��@���(|��J��DDz��ޛ�޵`3el����Z���?L�o;�]�`}��V,˹�s����&��$��M�ڴ�09wF��L`nȝ �W�0�LM��u͡j�QI�]f�މ���sE��/<�Ƥ�?�I��dP�MH܋�zߚ`r�0t����)��2�,2�I�$c�s4g�w4��h�ՠw޻�ie���6F�LnL��u�mn͝9�֬[�j�{D�2,qH�#�h�ՠw޻��nڰ(D$�})$�ZP:�٠[R˸4�C��8���s@ś����v��f���BK�	��w��Y4&�CQѴ�gW^vz�{S�Gr,v��ktR�th��;��{�}����97A�׀�߿Z��u��ݛٛj�3ޫ* �$��� 筚k���`r�`yu�"|e�]w�r�7`{kvlfm�9%3�{�X�女��~E�ۉH�MH܋@�w4]#L�&06\��ݙA0YY�VVfaxe�`r�`�1������7$��O��@ b}��Z��!5S�k��V��ma`
�z�X����[977%�*NSC�we9f��".�4dh0��t1Y1�\���W&�� ]zw6΍ؓtcu)L�z x%,n�lӱ�l�lZ�*l�<�.�f��Ȟ��#J*�������������k���k��'o*&����P-��3ְGZ[��xn��ό��>����!fj�)u��!.��ֵ��ʮ�:������x���H~f�Qz���VE���q6�����=��c�D��a�����w��yƢdn�$����@�v�����=��s@3ݦ;�R3�$���f��ɛ�j�ս֬��w��d�|����1ő��D��=oۚ���h=l�;]�@�����s �&ڰ1f� �7]��ٰ�
'7{�`o�>D�#$��ۙ���@��g>����V,ݵ`5�n�L��\c=$���]Da��de�MZ���rm��k�w=p� ۲�k�a�KQM~m�e� ��4��݋ �c�m�'�ys2�٬ˬ˹'�����EpB!��Q򈄐�Y��`�������%�#�� ��1I ������ 筚k�h����YF�梍�w���10t���rS{�L]n�g�Lv8�f�I4�j�:"!,���j��V�n� �$�A��5�gaӫng�sɰ����k�*��i��L�d�v&KU���{	6.S{�L]#L�&06\���#Y���A�$"RL�=��s@9�f��ٰ=����J"d<n��"r�%P�������mn͟o�D
!ģJ�[д�#FI2x "v�Eh|�ORh�#�#p��ŲBBE�� "F		0���"�Vb�H0H*�(A`�F�	�D�jB��c
���*����F�,�BF��Ѣ1��$�B�
KA��"�dB�C]0B�)����AI$C*�B#�"2�
��bĀB�R�D_S��RP�!�T`)FiSN�+9��y`@���a
��i2�BKQ��� ��@���B� �0$R�H+�M�}.�CB�օ>�Q�@�,F0�`B�����7-qd%2VR{tp��g9�b	�D_<A^ -_@Z��̈�/� h
��+�+��!I�(��j���аb <IDC��]�V�ڰ>YY(�:�]K��В���>�3w�X�vրs�������7�4�"r-�͵`~�Z��������ݛg۲���ZK���;e��d�lI�6B�N��i�ix,DDu0���qU�L��F��L`l�)��Ѧ�J7?5l���䙠��@�v�ٻj�ś����
P.�¯�NU9r�tKm���~�ٻj�ś��޶h;V:SX��-��r�ś��ٺ�?D ���	(�D�T�
o��}��s��T�3Xd�3�i�`b��V䒜�����6�n�{��OY!�4ĤkI�=���-i�۵��9ͪ۔�۟*�nVCTtn��$�Ĝ� ﭚk�h������h�?,/�8أP�H��=��7��L��V��`���D%�#���>���ȚC�9���ۚ���h}l�;]�@�l@��I�F�d��Y�j�=�������t(Q���߼�]\U~��.�uL)�-� �n��[�`{7mX�vՁ�DDF�~}�����@K��%��5���N�"�IW���M-5t9�P�$m��ȋ�7h�Qr%�m�Rj9�5۷\c����;Wl��z�i3�l��j�[�"�<���WJf��\n4t�҂F��U٢AГ�[�I^�{�2���-�+����ql�ZbM��c�N\�Ҭ�q�N�������W)n�ccfLmk����۳�A]g]{Y�e��{����w~;�-���l����u�\��q,�6���X9��Q�0�����@M��[�nkts{TKm����ٻj�ś��ٺ�v���(����@�����Hս֬���[�`f�ԫpSL�m�3M�nڰ=��6��)�����4��VDAH"2HLI��7�J`l�)��#L?���Ɂ�\�}��6F�I$qh�ՠw��h�[��w�ՠ���2~"��O�;��Rr#6J�:�LF�1�E�Y"��\]]=&!9�Ɖ"r-��s@�z���v��ڴ����D����0ܓ�߾ٿ�|� ���	%�\��/��M��]�`}��Vs��w�Q(�n���s��h��`{z4���4��
�)^VV|e�^e06\����i�ˤi���9ڱ�$iE�H
8��9�]���/�s8|��@�v� �"��-���sr��ә����ML�Âl���wX{e!X� )���gj�wͷ�~���뒘.J`oti�x�+0Dd�����s�ՠv�V��z�h�[��bGr����l���H��=�w�rO=�훟�v�<`��((S��j��Ձ�Y�`|�Y&�*���D�Z}빠{=n��;V���Z{bE"LRL�L�=��Ձ�/kή�=���ݔ�-�v� g�W0���� ��P��i��{9��8�tam���[��]����u�L�%�7�4���4�lw ��9�F��hVנw޻����h�oؐw�,�dJ&��$$��I��.������KZ͟�2$�JI�s���<�[$���1�<��`DQ# |G����k�g�����S��I��Jf��>�ݛ�_�o���|�~i�ˤi�oQȵR�e����vf��l���F�z��sŋ���G7͵��������dl��G���M����;����9�j�9�~E�ԊH�D������V�i��)���U����R$�#��4g�ۚ<�͟��3��Ł��j��z��ةs.��b/Vb`{�J`{fA��Ѧ����� ��o�����E�s�R��	,���b��V�[�`4��%����?g����`�N��vغ{g�[L�k��3��Ц�ʗQZ�n��[&�a/S�y;��N�tq�7U��l��$mț�SKz��c{�IӺ�`��m�NJV�~q�|�#�׶ϗu�m֨���p���`����H�k 1��u��N����J�N֎�Y�����ZЌ�G�-�N�,яP-��j�=�t$h���jK��K4a&�Y�W�T�p_D�����O5ɫ��SXj������Y9�뜺+v^9zKf"+���P�&��$G!�;�������;W������@��͟�2$�JI�[Ѧ���d����U{�gآR
"I�3@�|�v�,���n��oZ�>YY(�:�՘ffe�0=� ����V�i��V�Θ?"�q�H�D�8h����b���{k�l��K��[3Ji\���+���3ř2���rY�gt��^V�]�����NR�+#;�^͵`}��6�n��J#���VgΏ�cQ(Ғ`�E&h�k�߳6)�B�J�h�b��/��I|��v���F���L=�cw ��Hb�G"�/��@�uY�DL���V����>����S��*�0.�/)��Ѧ]#Lu�LN��=�[͟�2$�JI�����<�Z/�4��s@�U��m5KBZXM�R�a�9
�䪤�n�J��k�=l�`�ٿ��s��+���~��~�뒘�`E�4������#���IZ�h���s��h�h��/�$�0�ӓ`{3mX�vՒ��脔TAD$�D�����C���-���؂�"�&(�N�`E�4��\���rS���O�L_:?��D�JI����s�ՠ_;i��Ѧ]#L	��.V|��-f���q�ٜ�0tj�0�q!�={L^�n���٣��{���n_�c��X�h��~���07�4���i��)�n�L2�\��	��́�͵���{�X��Z�h���?dI��4
�vՁ�V����{k�l��V �6�-̙�s3&�kZ�ru�
�����`~���lfm�
�
bIDRQ�DX��Ձ�k%�T:����́:��F�t�0=�%0=�|0�-�.	��]f�9[���HD���K�M�nN^i������V=�9�e�Cٛj�՛����g��$�A����-��?��H�lL�f�s��o�~����t���6�6��Q
d�+I�*Q%$�L�L�;_�-�ڴ��s@��w4;�cw ��L��G"��	(J{_t��֬Y�j��(�c�Z�|�����I)Z{빠>Q�{��mp��Vd��BP�DD�AU�ʠ ���AU��
��PU����AW�����F*A`	E�0Ab#E�!E�P��Q�DX��DX(Q
�E�A`1*(#E�DX�)E��b��DX" E���`��bE��dQ0IE�DX�B
 Q
P�Q"�DX �B
�DX�A`�AP�$ ��E�� T  1DX�DXB0DXD@DYT!E���_��*��AU� ��A^

��U� ����_� ���AW��!b��# ����e5�׻��fRݘ� �s2}p<� �        P        ��  �  �P*��(���AAB�E(P
  R���Q@� ��   (�TQ�  ��@P� � Y `z" �`QA: ް ��� w/���]��w>�ݞ�w׼�}�9��{�yO9�|  �|���y<T����/>ޗ�^��ܫ��^�7�
 ����uTɪwWǻ���� >� B@  P�
'�R��v��&�b�_}��C��b�w��N�x�:��� gJ�3].;��1��}*�Ы�x ���۪�rʪŪ��n�\� ʪŪ�žﻯ^v�Ye��( �� {�>��{��m\�WW��^��(n�Ӝ�S��S�r�[ż+��9���ε95� �>��U�������@y�V��s�yn��ܯ��_p���	���VM|�s۾Y�n�_��(@ �� �� �������7He�Z}��W��
zT�j�>��3ɨ�Z����[�+'���}�|6�-����w��P[})��)�����G���7+����ﵧ����\���&��� ��PUP��%EH�3 ;�/v{�N�����&�{ϰ �ft � � � � [ " l     l  �   -` "(3�� ���D @    4�6ҥ*  S�#S5R�4� <z�T�4��  D�*�#�*��db41O�BSmT�R ` "�)��*zD�'�l(O�O�Y�y��3�s�e����N��qݽ_֑PUt�"���TEO�PU�"����
��DQT����F��t��j�o[�����~�?�*E�F��A��D��?H���>�u����HO��8@�hG��T8�a$H@)���͙��V�SFݱ!�B$

2�!�@��F1S�������RF$M���th��Y @ WP�.��sP�j���rjD4䐆�Y�V&�X��-X��"0 �!�vH<t@�,�$�c$�t`l��B0�,I,���FM������o���$��Հ^�v�CB~ޯ߿g�х�og	�|h��V�ē�)��x��,��Lt��p:�H�H�F?�l��cMY���jߋ%!XI �t\��~��|)��v�> �X6O�X�1g�B~?a�?0�Ӣ&��8����t$J�!��Q���ɾ~9�i5����}�>7j�Md�o�߸������τ�oy��樂0�¬H�:HV��Eх#JB�B[�����6B�P�!D�4��!�t�!��Dc.�6}��B���ɭ:a�߿r��d)����Ͽf��)�tF�5�f�K�� ��`$X��a!��4�(pxl�(B�
�����q	GBc��rCD���8�4�bGd9��H��0�����9d80)
p!t�b�N)��a��)�n'�XRh�l8l# #ta����S��Ji"��T�5tA����.�XSa�Zblɚ鐺�w\��u�e���ZjB��d�	�ӈqaM)))�@ػ0fkfJh`U��l6ĊĈ[����C5��)3P&�.h��2�0!T�c����K�2o`��%5���4�����bB��AF  S�>WN"=�[J@��8���f�%	+���Wi��,Ն0+���MI�J�0v$����+�H���2G6RBIMol*��c+���$ HP#aI�i�T�DO�٬�r�oA�h��CFi��H@�A���I������#lu�&��H�4͙m�k���l��V9��,�(d��h��U�I`��u!���B������� ВZu`GY�BF%����C!\N������&R�4��W�tF�;BFn	X�R!A�1�l�$RM8n4B�?#�4Z��%�8a�!��"V�a��6F�$!$��PіX�#
!�`�J.�$�Mc,� �$�L�����IcHE5$Z2E(HF�!	�C.�~��ԉu�g6m?F#K$A&f�6��ZT�H&В�0֩�o�7� ; Dd �H���%BF�BB$���ei$	m��I s��$��𐀜d!�@�B��H4c���F�B0$B�!FH�4~@����T�a���rc��O�@��	���~��Bb~��� ,#CI!"A��C$�:��a ̥ �2@��1[	+��������H�	!���j� 6�p�k.���X#C��mB5юؤ#CI���A+!��"����X��Q0-�ta"F�HF�X&�Cђl"B�0܏p$ɣ7�8V$k��$�5�N�+���|�6CK����H�4f�Cc�6k/���npk]\���Y7Nr��_�u������q��%a␪�W�\�!�$ԖC�v<vȐl&�n;(#M���H�$ �4�l��,#t�!tŉ��ma#CKCCi�1��ťt���� :�����s���9���\
�r�g��N$T�jD	�Y�e��[�!t�Ɖ�#!E�A
��qH$BD�a��!�k��!�?&�8��|���G�l��D �R��~	�1��v�'#�dh����D����bSFǀ@��k�����"PÒ��r�9Cf��Ӵ��p#d[BXj��D��~�����
���^o�ѽ��n������s���]8l�F����/�Z�Ѡ벑�`���QީÄ�,�p�su0ĊEH�`5��Ms�ă]8�< �@
���RS6�˼6Ja�c]8�	�L&m?l��l
 B�t`K�YM&1��v�l�͒�l�	
�sd�<d5)�hi�C)��E�b.�y��o	d��l"���b(� �i D"��F�B�D���!c#@�B4XT�`PM&B��Ml��$$��H�"�I!C$HŅ)���9
L6mH4ю�$i ���$
p&����|$�dK&V�Y�O�N�]I��K�5B�1x���a>�����9"�3h��~�il��"�
�A�Cm8S���`l�CH� ����0H(��A�	��Ѱ�l5ӵ�&�%tὐ���@�f��x�Z�H�"�04�jh��p�@٠�D�w6nP�,�&�����4�d
��!�-��aD��*9M酐7��B�n�8�#����F%]0)��L"kS0��Q#`��d�]dij��3�!�!#2Y�3D�[�Z�\�|�����H� �TM��)��';�����u �48�ĊQb�@ �`�5�W�F[�>����j��P" Pb�36��|h��!O�7�;6����� � �AHAR��F�ԃT�T`���@� �b�FH`�BKH"GBAJb�J@B"D"����E��0 h�$a!�]1�8I+�&.��	�@�Z�d���L
���h���²щ"DcbD"BH- �eR!L)���(S���0(� q�w
hH��ɚ��4�� "R4"�X�����$4��D(djŋ�q�R�6�X%4`GlB+ ����	H�`p��c����,����q#FR�`B�7�dY���s|+ā�ԃ1w$���5�]��?_�7������D� ��#X�@��EB�Bi dV�#�]6��B��)$��^��WH���&��*�o�!���l"
p
qbH�>&#3Of,�`�bߪ�dm�$�@   �>                                                                      -�$                 ��                                                            ��         �j�m-�T\�J��K�6��� ��I�5� o@� 6ٴ�]6    -�/�۶��m��� �٥����8!m[[l�0(  ���`�  p[@  $  ��  �`[���z�8m6�  �q�� m����]68 p:N 	��*�R�-��m��6Z ��$��n����mH��n[Rp�lf�[@k�:	05�-��$�      ��>�    �i�  iͦ�� ;m�6�� ګj�e\=��U[U �2$5�l��)�H4PAKN��ت�TB�E�۱��[@�;Em��ڱz�G    A�Td%�*��,�*�V���9��t��6�/]�n�  �` 9:8l��F�57Z��� mӡ��7f�6  �%�ڑ���m� ��۰�X��I�ip 9ö�Vɛ �my��moP   s�BKi"�'�U��R�T���@	]�o[N�H [@�i  	 A��v��m6���e٪��jU�@5M�YЄ�v0�@-�Tp*�a�   pM� �j���ZZ�j�����>�߄��m���*��+�U\l� z�淳k�gKr�*�ƅiyj���FR�&Am  -�m�� �`���M�WH�ӢZ�]���[@۫n�c,��`   vۯJ�kZBV|���MrUW@��7k�Ͳۖ�&�r۸    m������l`MR�aYYZ�c`U�U�>>�V����@_RU*���n�bY$�L�U*�l(<T	 =�pp٫ҧ��`�54ki�@�*Yc#���V�Pg�I�e�@�w:^���Ԯt�e�N l  ����E�m�n�m,(A[$6[,�m*�U��h�ZNt�h���@[b��[���e��/�xm�IVݳ�Ŵ�(���h	Ѷ��`� ���l�@�Y�:��$ ۶����	��L[v��� n�u� 	�]J�6�	�(���*UUUM�eZ�հ 6��r�%���6ީ��PHmB8�UԂ���d@���8d�mm ְ�h����V�X��T5�Kh�$�-�^����G /[\$#�Ϊ�GHq�ꚬ�T��U1���Z���U`���;/�_}	+l�� U,q*��YNj���
�:���V�ԯ<ʭ2�[Rafv8���2,�]�� 8����8�g6�h�m 8$�K]�A� ��Zl��-���)˫MBF� ��h�*�CԨW:%L�;+U	5� ��f��Ϛ�  @m�:�     ���6��l  � #�� -�*�]�H j�����Y`��@    7m��B@  A����M� |:I��෮���d���mq۶��y��!qe{b�q $�ld�l�\��%nm�]�$[m�N[����4� �k��[U[����  ��d� $�t�n��&j����nZ�|�T�J���8�*�I���kl t���^ֺ��[r� g��]6� �fʵ*کX)U٫���6��Ӆ�m�iX�l ��68�z�G���|��}T#�ަ�Җ�u���Ͷ�6� 6֭��u������Vض�/PHI�ٳv� 2� Ry�V�55+�ev�p6�6` �� ���6��L�`m�Hתڵ���  ��m�k#�\p-��H-� n�˛ni�����'��8�` �ܒ� r� m[ ��m�� 4�KͶ��j�z��U����  �m �h	�m���pmsm�NkXݖ� p n���\�  I �� $� m� @8� m�09 I  ��m�`Hhm�0�_����` $ �`  l@�Ãm�m�l���[n�   ��Ԡ[Cm�$   8 �i�m��(m�E ���i$�\�具9m �7m� � -���k� �HV�ޠ6�"�ݶݭ�4	�ݭ�*�P�]�
�
�
�͌h#]&�[�	'M�E�xݜ��FE�vݪ��UVV��]&���ګHȑ&�z��X%]��kv���:�M�M���[�	$6� UT�*�Vҭ� �v�����h������om� �[�[D��6�]R R��*�l	�U*�6��k�]�� ��#�^kk��VUU55@%��I\�jU���#�U�� ���M�3���[sI���u�̼ʪ0P�w3���j�Vm&#j�h�mʒ�8mW�[��@6���N���@  _������Q��V���ؕ2s��Y*�B�� -�ց��m $�p$-�t�涀�	E�Sv�B�
U�
���h��1�֛-`�	 8  � k���i6�h��ѥ6�q�`l86�۴� m���-�m�[����J-d�m�  ����β��d���Ͷ8�����Q��׵�ᶺI� �6n�R$m�   6�cn��I��f�
U��'f�r��D�) *�UUR�U-2շ 6͸ $  �j��Im�.F-�����M@�S�m6[q"t��.ٶؐ   ���V�h��r� ���:���NQ6��t�plm��  8 �`�$ Ie����sr��6� @�� 6n�����mH   	�l	Mjۙ $��A�l%��ˇE���[V�$���   [@$�ճ�p�m�`�� 2[d��t��W-�`I�y���}����  ԀH �p    �m� :��*�S�sƋ��ԥ�� 6�  H H���m� h     ��� �`      �F��	h  M۷��m�� m�,]� � l�� m        $ [@ [@f�m��� A 6�ޑo\�+UA�T��j�c]P UUP��v�N�d��N�h s#�V6nղCZ� �N��-�i�`�2�6�m����0v�V l �  $	�v���#[l�j m��m�   �Ā   $  6���֭E��� ���pմ����[@ H�`E���-�#Y&Ț`� K(���   r�H  m�� ���5� ;l�Yt�E{�  �p  ���Hu�B���f�@h �� mvÀ�v�l  �Z�p�[Z,�۶��.     l   h�p�H$	:�l�E�� 8�mm8H8�� [@       �� �j  � m�Ƚ��g	���(�� -�	   ���m�n�v�հ	mm �RZ����ـ�UBl]��m $  �  [@	�k~��7��ݱƚ͒ 8�  '>��E��`�K-���������m��m�H���v�n�$��(r������� ִ��"ڷ�����ƚ����:]�
yX9�Gmc�+g�g���8��-�)u�'/��^�GJ`��]�B��֪�z�N�@HO]mz����jAr�ڞ�����n\�@2�*�{vy��F�$��:۶ͤ�5u�ڑnM"(���+�*UUW<���,uZ��v��%�Ā,0�ӭ� �>5�Ll����հ   &� %YV�U�^U��i	��   [@ Vڶ�8�K��x���.�6� -�Ei��m����l ��  M���m�6���V��EW������dP[\    lp �kM�nͰ�6�q�ml��e�3333-���TEM�( �@C���� �Q0
AE�.E�DA�W���E� ` yUP�b`�X���E��Y"��h(R
�R1�HQT҆�D��AC�Oʅ 
~P�('Ȼ��������E����4�� t*~@���Gm A* +�~>D>0@� �AG𮄐F� �,�$QB���(��E@#�P�P �v��\���Q1�� Ѐ@� �ED`� ^��:TGj~>�f�E>?"~Q9,{�M��Pꠎ��@D���Q(���@�C��WBH��~�(�� 8����*
����"�b��1=�{�ߏƵ��    ��        ��`  kX           l lKYt˒�����[�2�d�e�S*���-ysg�r뗉z�۰F��
v�$�(90ݬ�hE��;l\i0��Z����+��c��m�Ӳ<PQ7+�,A��+�Ɲ�Be�iV8@.� Y��t�K6gX��*�3��T��n;N�ʀ��*��e\/�9õ��W\���P��v݊R��1	u�]-�]%$��r:�h;��J+�<����Ck M�U-KU�M*�[�5�^�*O5��[�'g����&�^�{�\�t;�lm!@�d\M.��KV��[8��j�6���������i����HpK7Y4�
h�u�t�/Y�W%6 �ͳr�7iW��� y�9�x�Ѱ����t4Q)-n�b�b��ζ9&'Hd�%�-.4��+vUv���/m��������	���9q�4���Y$ ݙZq�N�Lܡ��Y�Y��.֛��c�ܐs��	ܡ�&���t�3�/m�M�W��]!�0Z[l�sD�_(N0t��n��1�Ž�62vev��Ӻlf57=�J\M��rK[�!�k�W���� �l�����T��k5�H��hn�%�p+r�`����)d�1�ڦ]��/ewm�\�.;]UuJ�9�%훓i�6IP,���m%Msh��E�m�rѵ�N�mڶ6��e�ʲdz�!j�X�@W��p���E��NܝGS��pT�ƩY� J��va��m�4:6^�k������R�*�<���Jv�:�ZU��"�WM�ت�]��yv������c��Cin�*�[m�SR�e\s�a��%��0���[v�N7[q�v�-���/eS�z�:܀S� ��;�9
�Y��k���[`0����6[I$�Cfy'j�0�$�8
vN�r���Q?�����iQD؇�w���3333333.�ҭUUUJc���	�ml�n��i��͖�J�ўzbW����/3�	�c��f�v��+�[��]�lۓI�$�i�),㦢�-=����Y�ẕ�N�ͷgS�kJ���]n��]#�����mʜf�ۦ�c�p�V픏F��h�\З��������χsQp��2u�ڙT��ެ��I8�7	:���u���w=��zu�8���(��v{ "�^�����7'n8܆�(�K!n���Ѫp?Gy��7��s �	"o����A>��������MD�,O�w��r%�bX�x�e�ոL�f�nkY�7ı,K��w6��� �	���b}۞�7ı,O�w��r%�bX���̉��%�b^-��A5Sj��U]Wy����$'�u�&�X�%���w�ND�,K��]ʛ�bX�%�ﻛND�,K����Yu5p�˭e��7ı,N~���r%�bX��w2&�X�%�y���ӑ,K��;*n%�b����~~8�	��������oq����7ı,K���6��bX�'�vT�Kı?}��iȖ%�g�����!�*<��]7Dkn6�uS�gR�J1�3��D@1�۴�Zt]�jk2�fD�Kı/���r%�bX����Sq,K���{ͧ"X�%�~7ı,O��p��uf\-�ZԳZ��r%�bX���D�"�O��U"dK_w|�ND�,K���D�Kı/���r%�bX?h�{e�L3	�Z�Z�Sq,K���wٴ�Kı/ﻙq,KĿ��siȖ%�bw��dMı,K�w�L&�p�Mh�s&ӑ,KĽ���7ı,K���6��bX�'��["n%�bX����6��bX�������2cK[����oq���ͧ"X�%����l���%�b~����r%�bX�ﻙq,q؏����ͷAd��q�]6r��6�R�s���b�x�� �ɮ�t�kWkYMf����r%�bX���l���%�b~����r%�bX�ﻙq,KĿ��siȖ%�`���s,���R�ֲ]k��bX�'﻾ͧ"X�%�~���7ı,K���6��bX�'��["n�ؖ%�{���)Bs0FJ�{���oq������dMı,K���ͧ"X�N#`" �P~GFD�O��l���%�b}߷ٴ�KǍ�?��.��s@��}���,K���6��bX�'��["n%�bX����6��bX�%���D�Kı>���֬˄�j��5�ͧ"X�%����ț�bX�'﻾ͧ"X�%�~���7ı,K���6��b]�7���ݿ;���VQ��f+��a��Gg\\X�cf�"�Md1Fժ2>����iq�.Ja�M�˘D�Kı>���Kı/�w2&�X�%�}��ӑ,K����dMı,K�w��	�\5�Z2�ɴ�Kı/�w2&�X�%�}��ӑ,K����dMı,K���fӑ,K���T�����]��]U�RB������ND�,K�{��7����wٴ�Kı/�w2&�X�%�x}gN�K�[����ֵ��ND�,K�{��7ı,O�w}�ND�,K��s"n%�`{�⊧�z#̉�~�3iȖ%�`��w^�.���u�]k��bX�'��ND�,K��s"n%�bX����m9ı,O��D�Kı<������೉&ȺҢ:y+1�u뎕��d��m�M�k�>��wwr�����:�a�k��%�b^�ّ7ı,K���6��bX�'��[ xȚ�bX�w���Kı/��ֵ�j��,�55�n�"n%�bX����m9ı,O��D�Kı?}���r%�bX�ﻙq,K��﷪^�Փ0�]K5�ͧ"X�%����ț�bX�'��ND�,K�}��Mı,K���ͧ"X�%���׶\��0՚�˘D�K�TlO�w�6��bX�'������bX�%��{�ND�,K�{��7ı-��������s4]k�u�@���o�Qq�$D
!V];���    ivw3 �Y}Z�ݻ>z�n�Z��퍵B�\�iB�>��v�񗶶3<�]�t�1�8���7R:�oe�뭓uXS��a�hӭm�� N��c!&k9플Z�:�ۯ.{f�ykO��R�LM��c��������6�08j Ḧ���	��cc&.y����<gGG��7\��/��ܶ^Ѣ��m�6��۰��dݴ����&��\��E�*m���7Z
�s<�x�I��8ț����M��X��_$�!/�6u�`�;	���5b��Uwx�x��&��X����u�ʇ;�jb��s4t�09t��7�cd��.X�l����bN.�����=kŁ*"Q?{_� =�5UN����EL��-�zt��0;z:`r�-�~�~w�ߪ�<�&;%��M�Q�5���;3�ݶ���b����ͥ�wLRqr�.Ū�&��{��׋ ��� >{f��/�b�$��j)3@�u��dB�	$DUk�����6�d����H>�[�	��LpL���9u�@6I��:`wL�հ�E�Wib.��ʫ�ID�>��7��`��`�נg$�X	��7E$�@�o*I-����l�u�������W8H5���p!�'a�#16��5��ۋ��u��m7��'d�ke���w������Il�L`l�� ������ۘL���9u�g�$���7��`�l�i;C�.nɚ
��殰�]�m��R�Q�"	�0 �t�%߽�lܓ�����q�E0S̊I�z۹�wu��9u�@>���\�"$L��������˭z��h��hgq+��0jc��Y2`�,��3,mQ��ڤ�ղs����#�+�%T�,�*��BUk1e��<�ȓ��*�����@��4���$�S	pn= ��vA����)�����F	��7E#�@��s@�빠r�^�}m�ʇ;�jb��7!�J!)������ >m��		DD+zS@>����ۈS#s4
�W�[f�oJh�w4�^��%ɋ%n�'\Wl��e��K�2s��8#gV�F靍�c����:���t3��zI�	; �����l�F]Ish�EP�n� om��%
�UCo�`=ΰ���iIând�v���Y�����ˤ��&06H�{=�f)��Lpo"Nf�˭z}l�=m��X�u�4���8�iL$q���@/���)�^빠Uz�$�>U�@u�wٙ��������ml  i���в\���l9!�4���F�*��n��K���eے�b��Mas�b��[��Zٸ�͚3OdػX�7��,Y�Ȉv�Ss��_�.��F�d�W%/jR��f�4;+67\�dE]oY텶�\��l!�uٳ]/&'���l���-�'9O=c�@k��=;��:;];��Ҽ��N|H�J��GM*��]Fet�`�Ӈ���a�b��y����v�p��f�1G�3�S�"q��?����h��h^�@/����I��S(�p�'tt��t�6L`I�����M�%2G3@��z}l������&{��s}� 5�t\ݓ4T�Cq���@��4�w4
�W�wv��&
!���-�M�%����:y�`�w�	�f]]YAGn"]�v���n�Z��ʘ�r�.�*l"�N3��=�PA�묄�컪������L]%�	�cd���ʙK(x)��I��9u�~������٠u빠^빠}�n�ěJa#�D�l��$tė���.��mLvm)�Œ<�@��s@���h�נwY�|�T��Nuk �u��9(��t���7׀y�� �Q	z�wUU]ڛ��J���A3�i�+���nMsP�X���z_$S:�j�X�MH����_ߞ�}�f��n�>����QH$�'IǠ���#����.��݅[��"LCdrM����빧���?#A�@	$RX,b�bI "
�
�b�a"D�A�F0�H��$CT���d��Q"@O�PC�SrBD�@ ©���*�ۭ��H�"���@���KZQ�*�!(����"�$B*+ "*z %Ѐ�D�D���P�&� �|����TЏ�U���_��*j�'��� � �_�����r6667���lA�,llt�x�չl�0��33�<����6?��p؃� � � � �]���UNA�����}�yAll~���b �`�`�`�zw���M��Z6(��k6lA�lll{���؃Ȉ�`�`�`�w�͈<���6?{���A�A�A�A�����@9-�F��o���MC�V��b	�����V�QV����v��<�����j��q3�.��?�������o������	(���|��Xr����r���	$��l]A5S6��U����{��� ?ʢkS�{�f�B�_krC���K�N�5�J��&欲���)�}��>N�u|���6�`���l�l�)�I�.�������9�������`0BD�#�`(>�ٜ7$����s&\�]�Y�%yl������2^� 3�.rH
2A��)�96��nRJ�On����4()�nM͵W"�]��]J�0Q�$�@���hu��9u�@=�f��c˔�D�$��~�[�s�<��â�r�� 5�����C{���g[��h�M�V��ʻ0/�VtDBS!���%	-���y���ďe��X�M�0���y����f.���7��`k�`:Ӭ����)�LJ,��rh��hu��9u����h�?�3��,�d�I$�I6   `�λ�Im�X����qÒ��//��N9k��v�Ɍ낭i1�˨�T�$diN�\q�t�ڱpU+o��z���
 ��W&
]Y����BBZ[	�����:�fn�n��4藎�9��5��@�h��F����U{���kjd�<��nk6��=�<.gVԸ3�M7W)l-�cOgu�=2���pZS/g�T=��
j^c/7*Z�c���8��+ݮ�ЈFJ���X�jng�z����\�@=�f��n�u��n6D6H�i'�.[ ���:`{�A�mr�v(�mb�ۏ@=�f��n��YM�]z����$H��$�@��s@����k�� �u�ݎ�"Q(�0lD�f��YM�]z��4[w4�R�ۏ1HrE>�ܶҪ%4�V���|�~�k��:�g���Li�L&2@l �>����z��x�x��$��}|`M�Q73U3h������� �뼴��$�)"P����Phd�����?~�~4]r����_��&(�b�ɠw�ߝ0=� ��ҥ�����'`,l��D��hu��9u����h��h^�&�dCd�6���.�-�{zcd���`v�����r�^�l��=]�`�ΪvyJ��.�VG4n(X�V�^�"y:h�ʺ�3䮲��L`l������J�@��䮒6��Q�I4[w4oGL]*[ �����1,K)]�h��`{^,gZu�����@��hz�h��0�<�CǑ'���}T��S�7�06H�7����.�D���)$�����?dow|���,gZu�}��*���SY���!�;���t3����s!��bk�^���FF�?��Ɖ�<���h��hz:`r�R�ޘ�򜒹����Rĳ�SoGO�UU$r�N�޳@��s@=�kI���$iH�h�T�7�06H�7���˱آ�m���<�@/����������*�P ���=��:�FM�ItM�SJ��`m��&"^��|.�^�}n��gJ��4�o�(�E�Ɲ�j���q���7l8j,�i�TckDD"Q)�L#��^���ҥ�&��'d��eE�s'3@��W�_[��[Қ�۬Q	�L$�dJdz�x��مDD%2���Ӭ��C�&(�H73@��4�)�U{+�/u��>W�N�X��%�N�l	�:`I�����!� /Z  Tڶ�y ��:m��3�9�%���ZIK���,�{F��_�ﱸP%�m��`��͡�m��Ol��Ԑ���5���h�x���٫�.�Х��Q�.C���7S��<����2�ݮh�\�0zs�:���iET	�8%��fS,���uGy���CɌ=�6��;J��jo8�;n�n��%u�mR��jꝽ���(HpY��Mx��f2�-tX���u�!n_@sȱ��
�%�eїQ���:y����X{l��)(I}A��- ����E�m��ĞG�}m��آ�;��6� ��u�{vY3m�1)�<�L�-�M�]���^�}n��c�H�Jb��"��'tt��uK`M��UUU)/ �>�[L'1��$�h^���]0$�wGLоJ^|U�%#98�\3G1�a����z烣���<�����EƎ-��b�LJa#�D�G�_[��[ҚW���g!��j�ʫX{l�
��˧ذ�k��}�s~���Ą�$݀�J	U���X������}� �w� }�J�mF�$�rL�*�����`��DB���, �D򮹊dm3�����)�_u��*���첶����'?�Lvnj�s1�mF���Ki�p�-<f�h:��d�h�J`��h���}�s@��W�_u��>�TR%���1H�0�x���:y����,��`���	��46D����^�_k�{l��ŀykQ7$Д�)$���٠[ҚW���eUF�i�b��$�=dt�����J��&��u\�ww��ɶΏg��B�/]�Fb�g��:{b�`�ǀnm���Ђ��.�:�e��'tt��ҥ�	�cd����[M��Cd��I�.�^�_[4[w4�w4��d"���LJ�-�M�$t�����J����T��#`��h��h��'�����]�F0�Q ��F�"�*�E ���"DcC�j��}��ŀ?Q�qs73jn�4IwV�	�09t�l	�06H����l.�.� ���vͷ�2�TE����r:6Nvړz��ﱻ.���m�����ج�u���9|���x�6�~ID}!�����D,h�E#q)���w7�D%2owb�;_b�6u�X�9wUS55%���ՓV�6�`��a�!)������nh+�7`<l�,��uk ~׋ �֝`��`r�S�������i��l�2I3@��+����<�ŀ?kŀZ���$(J�V�����E�v�0�����$���0�	k`�V��:1j���$� ��Ą���C�J���1HB,P��`�EH�Y�1.
�tS� � b���FaT��1"E�H�XX&�A,�"�4�E! �*B$GB�.$Ą*�EP�� 4Ҏ�0�X��A�`��E�% ���h�:�d$ �`X,H�$�!@ЊA`D���#����     m�        'l  m�             �^�lm��25C����ȅ#\��J�����z��e�E1ٻv�s������A:l��4ڝ���!w�5q��[Ag3;��s^�Hpkv����|i���!l����SjI�b��v{`�֋U@Q@Og<�԰fM5����6j�v�݋��a�ʦt4��@�Wk����@��:v���9ʎ0�5:@͵E�[5D��<:bwIX��H�����!Y@������u<�P�++�:����y�nҳ���gX��ez�[���u�P��*����R.�c=P�V75Z�L�l��,I�id�$�E�ð���7�L��嗊p�C�mյZ#�C�[7&Zc*#P���6xw����ZSsh�ssϡH�vkY���;Eu���r��6�	1rD�6[\�SzN�Y�)y���͎�49� JKJ�Ma��vڭ�Uㅊj����vU�E���+jx'v�؉�;\5�(�݃�6�mm��G&��B7N���!s�,F�嬙�X�V�����QW�9��љ]��6�yE��ڥ����f��BU�&�G,��G�Ap\��X��cW]cnRMY)�m3����a������P�O�e�@�-�L��}�%ɍ�����]���ꫩ�1Nh�z\��$��玬��U���T��<���*�R�UPr���崪y@�$0h�3c�i&��\ <QK�J�Wl�Q��n\]7sR���m�nk�-u.d�D
�T��J9r̪���Ʈ�l����kh��q�I@U+k;iy/[�ԗ�l�*d�E�0��Y��P�b��gӞ$bm�+����#G;6���i�utq�m[tl)*���˱v�ңU(�r�����;B�C�_|��\˖��UB*ڠb<�� C��o�"m�� /7��� h  ��r9�aq����^qϮӫv�=rd{T�:H�l�f�{M<�q���o�7/&	�v��ș����`�o777n��m��tNV-m÷�ŌZ���^�V�`&:��u�;�6�]k{:.�6��B��[� h�I��#��ې$:X˰�Sz&ݦ���i9�ƝV�r����`�Ѳ�z�w���vK�*��'\*k��Btm.͋�#�i�͝Z"���7�̽�\���!Db1ɉ<���~���z۹�_u��9u���ˣ��Ħx2�$t�����J������2��(���&"G3@�빠r�R�z:`l�� �Բ%�X,��v`�)�˥K`M�遲GL	��V�X�0�F�S#�/��`l��oGL]*[e_L��/.8��z�gv �H��K��r^m�����e6jŔ�eF�6����:`M��˥K`M���]�aj��J��ʫX��YP�	~I$�JP��B$���/�V ������׊��j!�H�$� �α����GLwGL��]����"O$��Қz���빠�l�;�%d�F(����h�:`{�:`*L`M�� ��J^]�9��xMӋ�Lv��4ř�su:�W�rű����R����!p�57|ʓdt��� ݩu"`�S$�'3@=r٠_[��n�� {�r�=ΜSs*iZ.n�U+��;{�`���ˢt�(��� w���h{*��6���wH�;�����Jtu�yjK�0��0Y"nf������w���;���*�kmǃR5bid�`�=��Zk>MsP��i�2OK�'Th5�ٴ��j!�H��4�-��w4�w4�S@;�]�0�#�D�^ct���:`N����{�c�h�#I���;���/YM ��f�z�����I�18	�̼��`*L`N����\���{+�
A��C@=r٠N���GL	� �:��)ywTR���T��i�ʌ�-=�:����v�~���S�>mYE�����E<�W�m�����0;�t��2eI���]�V�"#����;���/YM ��f�z����]��ɂ�I�h�A�l�1�:GL�0ur�X�Q�)�n����������hrK��b1ȓ�&��#�t��&A�l�1�P�A�E���J}�{ك� ��  ��,��,�	�KsAb��q�۶<�(��Q�$A��i�&�Zr��vH��Z���},��Y)vئ�7 l�z(�+��][���j�%���v������Nlr�I.�ٖ��sq�v[�����;�r]q�R9����O+��f�n�Θ���������۲p���u�y3���%�n��.��4]�w��n(%\i�'>ڵ����m�IXi���\�]i�Ev%�76�k�m[I�ή�Oi�[e��߿b�<ݳ <�w�!/��ŀ{�ʏ�I�18	����=l��zT�����GLueB��������t���:`l�M��qV�by0�G��@�s@�s@������e���h�R)��w[��z�M ��f��n��e��rd���li�bS%�R�5
[��k�0��aŞ{.���B�v��6LBH73@����������� ���I�5�"��i��$�*���`��`nٜ�JR�?4L��r$�ɠ[����n��e4�-��Tl��#�1��nf��n��e4�-����}��:%��4�7�����`��.���ذ��`�����"9�77:��#�%5��m�����(�<-��&�U�����=��e�5� �]׀n�� �o����;v\��0�s0֌�ܓ�ݛ�PF��݋ ��� <�w�l�9wUS55!jn�����,��8	@y�� �����.��d��p�-} �1�'GL��`���&&���IŠ�h���=zS@��Z쵥�,@�dȤf)%N ��ΪvL���@;��l��^�#�	�2df!ȓ�&�o]�ץ4_U��h{�'���S�yL��0$���vԘ������E"M)��&)��k����޻��Jh������ 6]]��tBP��z�� �}� ��f�.����rN��z�ita��a��������0$���vԘ���w~�~~�m˔;l��/=6���vV�l�o<U�M��b�k��<[]�Z��|`ֹ��n����>^�`,l�,�����k����޻��Jhݜ�L��d��%x�mI�	::`l�K�ԕ´L��r$�ɠ[�s@����0ړޔ�����7���Jh��@;�l�/�����I'����!� .�   4��ͮ���%��N��&M���-�+k&�kmW���:q#'��W��c�@:�-�m�`�q�]�M˙޽2+Z���:iĘ̰��s�%�r�kӤ��&6����I䮸9^.�Ʈ�����f884�i���!d��;O؈��:�]���H�N�ju:��=�7#Y-Oh솆i*�j�g����
�ҋ�9���{�����_C�t�m�Y^,i�E�+1�`��.�������m=y�X��X-.!1H�4ߝ�����޻��Jh��FL
c�6G$Z��1�'GL��`I}~��h�SdȔ��&�o]�ץ4_U��h\�YHl"�F�h��`I} �1�'GL-��&!&$�Z�� �e�@��,�m��I���~�R�l�u6J��/�� ���,ZV^�Ξgk���"�Ç�

dQ&Fɉ�5?�q|{?~��w4^��-}V�uEaZ&L���tJ���x��K����� �Ӏ��4��Ɋ!�S��h^�0$���v�L`I��e�1&����C@��Z�γ@�����M ��d��9�drE���tt���K��|��컅3��Z6�����up�]rtsvW����7��X���d�c�4/s�7���f �k���_H=T�t�
�����LJD�s4�Jh��@�c��Jh^uD<l�J��L՘ε��U�p�Ę�*��H��Dd3��D`�������a�G��$M!,�`��T7 �V@"�R0�� ��X�H��� b$H< ��
5(X�* � �(�uC�lQ4�� ��*���:؆����7$�~���Z*�#d�ڍO�Z{U�w�S@�����}V�qk
� F`ԑ<�-�Қץ4���>� �Q���UWUE]���]*��ų!�*�cn:�Q�W^�˥�3K1Hʵ��k1�nC�=��Ɓ�}V����h���=_
��4�7�)��e�Lھ��'GLN�06��S��������j�-빠w[��Z�����L7�7�D����t��_D��edi�uh��mbl&%"r9�u�����6Uș�I�JJ�2����H��Cs�']��E�d��5��OA�-x�8{6��y2@n(�������䒵�-I%��E�$���i$���{�$.�KL��j5?�pZ�K�%��Jۺ�K�߳�J�(�$���´L��)y_|�V��Ԓ]���|�V�E�$�rZ��$��K�chl�7�I%�'��I)/ �I-��/y$����$�����4�7�$��>�$���i$�VH�䒒6$�t��y$���: $X�X�	��O�~A� $  *��-��$�홈�݄ڱ�6�ͻm�HpF�v�k��Ӑ��i���g׮���g[;�͘}�=�;��n%э�Y[�]��n�z0щU�2�u��%ʉC˵)�.s�-۰`]j	K#��l�Kqڙ]6A�ݰ���(s����: ���j�f�=D��&�{rb�(����
;�'P���Y�[!�j��E�?7w����P��\���Y�;Z�7j����t:㓝�v5���>����bH�����]�6G$I%�/�}�I[wCRIw[�}�IZ����;��Ҙ,n"%$o��$���i$���{�%%�I%�����$w���������jI.�=^�IIy�Il��{�%$lI/?:�6L����䒵�-I%�Y"��JH�4�]�z����yۍL@�����j�䒶����䒵�-I%^^��$��E]�����M���B֌�npse�nܱͼ�����6���d��iH����䒶�I%�'��I)/ �I-��/y$��d�1�6
b��I%�o�����ٟve���M$�md��I)#`�IzsK,L��Cx��L�䒵�-I%���$���i$���{�$iu%��.������+��KV�I[wCRI{�su$���jI/������cq)��^�II�K�OW��R^A4�[2Z��$��lm���mb���d�sa�B�5r�:��h<���x��Xm-by �#�@Ԓ]���|�V�E�$�VH�䒒6$��������(_ffy^�IIy�Il��{�%$lI.�~ϾI!{�i�<�jF� RRIl��{�%$lN���U_��x�$�>�$��pԒKܗ4�dɑ�ҐY���I.��4�]�z��[#���ْ���%_GrL��L�7RIwI���Il��Ked��I.��4��?��?����S�Q�g�!���n��8W,[�e^wSO n�s�\�]�ffW��Kdx4�[+$^�IwF�RIw[�}�IZ2`�S�?�8ƒKed��I.��4�]�z��[#�RI}���6���H�I�$�u�$�t��y$���i$�VH��6������A(G$��/�7o��ϾI%߿<I-��/y$����9F�����s�!�d�I!ϾI%�v�K�%��I.��4�]�z�䒊�wwy�W�oN�]���!�鶁�p����\	��ƈ��8�k �!��k���� ?�Y"��K�6$�t��y$���i$��.iVɓ#��E��%�wCRIwI���Il��Ked��I)|�Ve6���n������^�a�$�VH��I%��(bV�U�"�Y���$��$�����]ѰԒ]���|�G����<�0O9�I%��E�$�tlI.�=^�I-����n���ww������ ~���� �^Z�Y0�NO7<��%�VqغԈ�p@�K���9uM�ĝS�m�ӱкD��u�:"u��Y��\��7�v#[b�-j�OH�X��<��4t�)V[�9��v�3��va����*��+u�Ý{k��t���lJ��vM��R��������n���4�p��2n�)�奮�rs�4	���Be۶�<\f]QՕ���fK������]��+�XN9�]u*��r���H�IܒV��I%�o���$�G�I%��E�$�[P���J�0K���i$���{�$�G�I%��E�$�u�I%��b�D<l�/�$#���$�G�I%��E�$�tlI.�=^�$�z���c�5��jI/\��y$��`�IwI���Il��Io%�*�2dc�$_|�]�t5$�u��y$���i$�Vt^�I
��U߿%��yy���y�Gd���ۧ��^��Þ%�76��+jۥQn�Q��-���S�~�{�$�G�I%�����K�=I%�NfX&���i�$�>�$��x;�������K�d���K�6$�m�g�$���&1���CRIzVt^�IwF������$��$���150x�DJD�8��$���jI.�=^�I-���_ƫ��N~^�I�����by �#�@Ԓ]�~ϾI/����>���y$����=�I%6����J��g;�fI5L�4u����%����ywZ������︾ё5���^V�I.����IwJp��K�6$��~ϾI!^���0��E#r�K��g�rQ	UT�ف�33����陟Sy[��{��@����]9�"uo��-�}�ɻm�����.*/�9�~���vԻ�6�|�K�ܑ�"0S��j��
�{���fv������ֱ�}3?����ƭ��MI%�O��S����e{�%�#�����}'���u$�?:`m�s@��n<i�2b�9�,p��@D��Sm�ˮx���e�둊Ag�������N��-��V��.��w���׋ ��s@�wW�}���68Ȕ���`n�Y�Q�DB��߱`=߫ �y)�}��]j7��"!1�3@��s@�w]a�(�o��y�ŀ})��\�5%�E���Z��IDϛ��5�0�^,
��
&b�o �USAt���nn��kV���o�_��nh��h���� M�L�Rf��1�&VuS�g7g�Y�Y{q`6
��t�H#J6L���md���u��=��hۮ�$��C_+� 7�+����&n
�����{[Ŝ�S!����_��s@��+,HiLn&�B9����V�:Dϛ�X>�X�KZ��H�Uh�Auw��w�g��X�x�?BJg���[ݔMM������Wu�0=�0;�t�=�1��VvnI����P҉���(E Ȥ��h��]-���B)&-;�����T:�T���h%w���bA${�o�J����Hh���KJq
.�b&QB)�p��"	��-D"���F$v���8��@������I;w�{����     m�        'l  ��             ��/bW�A��j�ڶ7"�ŝ���hV�e��W8�iݗ��5s��.�k��d���n^�Nۤ����X08xۍ>�[q�)M�6b���\mCn2v�[k�
���!6��պ�m����H䝉�*n�S!Ý�=�q*.����M�(��;���( �����tUuĴ�1��V�p�MrW.�BM�*��Ns��&M��[N��(�n�;m.�!���{6�@]��� Ea�5j[I�p�J�!N!���+�<�����'@�CN��'gq�0U*ҫ8�M�ػ�6�{9��ԫj�ѷUA�ʵYv z�ݍ�豯P$rA�2��[S��[n�O��C�m\�,�m[�acd�nE͵��P	�i[ti
Ó���ձ��-�H�ڷk������Yg;Ky���盘��(93��b��|���Q�y��52�E�d2�H6+vP��4v��	^R�Fb�!ՙ�8���0�f�(���6#;v�����J�yz����yv	�/=if�ST�� n;�}�C[.���R��zt�e]MoS2c�Nn.�,q+W[S#�)�����Eg�.�75u�'8
8U�#L R�q������Fц�u�![(����8.��@��l\v���USJP���Sq�s;-�Uvu��v�+�V��-��Mmě �]%l٪�C�ڨ z���8۴郝�HR���o*�vѷJ� =�m�pUU^U�-��U�.壝��/F�W������h@T�U*�*Ҭ�Mj<�OS�UR�2��uq��کs��+j^d�ڠ#v�d��ĬY�a÷m5O&����cse����e���;۵W����؍�S��9vـ��U�S�ļ�7IUC6��fx�;;��]nv�ʪdtUT��0�����Hp�(`���S�(���P��
/���1� K(  ��a����q�<���l�����X�ӷpbȜm�Vm�q���
6K��+.�Q����P�P�m��rK=-�h��G%��]�!�|Ƶ6N.ΌO�;���`�7<�Ɇ�JX���Rs��[nm�����7Z�M�XA�l��������>�r9�/[n��Ԋ�Fl<(�s^��dx�{;$��*�Q��us�]9�q1�5ȷ����<V��d��v�_��v���/-�]i�w�����X��x�VΈ���ŀzSS4@�BG3@����=nJhn�X�x��d�������-U]�sV��W���ŀn�� �u��Z݉F�1�#k$4����s@���h뒚��D�0�E�bY��ޑ����zVA�����������Ͽ@���<��"�,�E�5�e�u�e�۞���n��!��ڈ�T8Xq����Z��/+�l��07�d�w4��\d��9��ɚ��پ�iC�|��K��ٹ'߻ݛ�׋9BQ2y7gISh�
�u7sUY�d�遽#���������O*n�UZ�j�Uwk�(�}�,�~t�ޕ�`{�:`yW\X�V�ʿ�Yy���tt�ޕ�`{�:`oI��{���Z_�!��J'��"�jim$,�RvcZ�w@\���8{a`�Tv�����B�yL�Y����}����uK�~�6�1��!�{�:`oH���遽+ �6t�*F��3q�&h�w4�������Q�!*Vk�|`�ذ�)t�*f�U�ME�Z�䒉�}���|`n������y�0x)�`��rf��+ ��tt��#�t�06�?nvsά�l�R�i#B�1F9n�;Y�s�w%[7��q�<7V�ػ<�t��f�:`l���dҲ��.�5��Y2�4[w4�)�{�Jh��h ��TCM1�D�̦t�07�d$t�ޑ���4�	�&8�2
C@�\��=kŀ{[Ł*9(QQ�}� k�|���H�8)�������u��7Z�`	z�>�����A5v�I�ڊj+[.�ve�&�h˗^^�=4�n����q�L��0���b�>�~���{����rS@�[��}�+u�)��UB��X��3�I)��W����n�|�r	���	�$s4�Y����0=�0=[a҅0x�̍H���u��=m��>�]��䦁�{)u��71d�L�L�6H�����+ ���t�����{�=���G�� z�  271�5��۬�{8�;v.�m���5�u��˳��ՎE9C:���v ��t�s��]5ym̻K`ۊ���8�cm֛Ӱ��vp�	$<^�܎�uu Sbn8sv�{O)�zD5�lQ�/<t��l�aGe�1��s�,���1ikX�:M��͎�e�nG�Σ-�t���3̀�nnܽ��'���O}}*�[`:�a�zN�Vf.h��g�|Z�pÎ�c6�����n��b2&�����Z��ҲoGL��h�Ǔk �rh�%3�"d��ŀowb�����3�]U6H�8)��빠z۹��1#�\�䦀{��m4�&���t�=:c�VA����r�CJcq6̒C@�{��;�Jh{���n���V�p�%&@�h�6��;Uzp㝞z��K��Y����뫉j�J����|���kŀ{[��!(_Hzu�`��Z�Jm]M�UV`���t��#����t����kq�nbɐ�$��z۹�|����%4��s@�yVW#hɏ �Y���ޖ�`{z:`l���ܱ$�cɍE�@�)�}�����^�V^��)��mt/^k���YhZ�8XQ�(��`.��t�6)�"I̍��1��!�}�[��ҲgL3�e�Ъ�䛵�{[Ŝ�!L��}X|���kŝ	L�t����*f�U�ME�Z�=:��֭�L$��|�!%�����h�w4���&1�O��u�n�l�>��X�x�9BJ}[�Z��������7���s@�[��|�k�=�%4����i�^#vW�jy�+3W4��tR/fŰ�9��$dj7��2d&I&h�]0<�K`oJ�07z:`y]s.쩩�Y4M��>�7Y�Dɯ��n�ŀ{[Ŝ���:D�D��-T�ī̶O՟��GL�0<�K`�m�Q6H�8����s@�^�ܓ���[��AB* %P���?����0���II����ˤ����{��]�������C�V�v,p�VtLj9��!^��z����N�+.2,+����Il�Y�GL�0&�ī&)���$z�䦁�빠wW� �u��J(����C�T�M�����v`�b�7[Ň%�ϥ�V����<������5hV��Wv���`N�X�V����:�|�H��H��FLy�I�˭z��Mۯ��,�IBIwe������݀��  �ۭ�2uJ��8�n<�cn��y�5�u٠���� {&礕�m�nvx�Iw޺pvۙq�5n� kts(7ny9�5�X�l,y��nb{M���k�������q�/Y,%�BʰPj E�k�wn��:����4�ӷ H&�ri{5�w.���tkb���,�t=�<�p�ǋ��COd�5q?���~�V�6�n��	�nm���uV�Mʚ�[z�n9.�E8�k �, �Lq�䜓�_~���=�w4�w4�h��W$M�c�%2C@��ŝ#}ذϺ�6���ڹ!#�mĔ��w[��u�@��)�{��hW�:І���m���`$��YI0;�t��0���&����rS@�k�t���0	[֔�
�ZY�dH�J�5W��r�����ݝ�ΰ�L�Z[x�����7�����7[ŀ}����J#��W��W&YJjЭYj��`���؄�bIjK�7LN��{���u���e�B�J�U7k �u��<ڶa�S>o�`����Uy��(
a1��5&h�[0�^,u�X���� 7�UrQ6H�8���빠w[��}�w4[��{:����3ǄD�.&=�I��Zi�y��z�Yd^x�vw6�k�m[t���Sp�a Fcn$�π�����빠zܔ�>��O+�iLn&�����ş�(S&�+� �}� ޷s@�0���&̊L�=nN��9��ٹ��J�O���"p��j�?h�v2���J�P�FY@��H�, �D]�|�X�bbDf��ё ��D��SHD� ��]FRЁ	BH� � �		�Bu�)�dHI�����P��$��t��ɤA �B`H1VE���I�.�H�X))��EP&��4*�$d Cjh��0`B$H%�$ ��Č#�� S�$ �ցٱ�1�0ͬ*2��CFE"E����VTF��-H��T
|:@�E��

	���6�x�� �Q���llo{s@��w4����s<S#R'u�0=�07�t��tt�ޕ�`|����)MZ�-Uݬ��,�G���k�|`n�X�ʪ�)]UU����$�&9��T(Qy4�2���k���]�ϭ*��dGli�&<q8)3@���hҲwGL�0"�uwV�,�*�/���`oJ�0=�07�t��u���\Cl�#p�Z��q�ӣ����J���l]0A�#1�Rf�׮��e4���%D���R���@6��3'�;}٠{�'��4�7lD�,u�0j����,^�XB�����~}�a[���w\�H3u��"5ESm�k���[����a�GY�Z��UuֻX��&���������n�׮��e4�<.9�)�����=lt��������_D��mB!��9�L��$��]��빠}�%4���w��J4dǌ�L�=�0=ҲwGLt�Yj��m�nT�ݬ�jـ~������k}� �u��:$���뻻Wwv ���  -��m�T�X��)IK6\�B��=Tp�[,v�'�0�ư���ڴ:�3�VדB�V�����83X��N�1�7)k�k[��{'C*�R%�ۣ�GK�r��{Y0;Q��з<����3<C�7=PJ��[͌%�EX�hۛ�(k��v�^u����Q�/e�%�jz�L]�.T+�����>C�MH�WV�]r&Va�l9�MR��}>�Lű^_n�d�Dcl�#s	��~��=�w4����\��U�	f;�IfS{������VA����:?�Q���� �mT��Ғ��`����+ ��tt����6���Q�ګ&j�.��D���07ذn�� �h�g���1��25&5��x������}׀}�[0���[v3�����D�PU�7�N5l��c\�s�kѼJt���i�&�y��e07�:`�czVA��GLsNʛ*jEj�VU����6"�P$��W*}8���^,��vZ��Lj,�hq�Z���~J���4�ߦ�x�Tel�#s	���<�ŀk׋ 7[�S��q�����	3q%&h�w4�٠{�Jh�w4�t�)2H�X���U,v�Vk�mk�ônz��n���1f�F�I6��b��M<D�f��ֽ�U� �o}!���S9Qh�mU�]���l�Y��:`j�^�}�{.\s<S#R&�C@�[��oH�KWGl�Y�q𺻹V]�ݬ�}�,e�V�jـ{���h�5�2c�G&hZ�`֭���X��X�"�~!��u�;�������ZA���8�����7WF�t.YJ�}� ��M�v�"�,��?V~�:`oH遫���Q��0�q�Jd���s����`/��kV� �Z)�at*������{[ŀzu�áL��|`~��>�J�-Ƣi��I3@��� ��l�=���؊�
 P��"�O�  �o��rN~�槍L&K�d�QwWu�{Z�`�Z��_���ֽ�%\���bQ���洱�e��ۇ]X�͑Ð��3u�����9��=7=Jm]M��+� ��� ��� =����(����]��ɹ�Ur���X��X���֭��x�b9$���yL�SR)RUMR����=���{�ۚ�s@����#�Lx�*�� �jـn�� �oBJ&w�� 4;�]T]�WV�m]��x��w4�٠zܔ�;��d�H �l   �2ɳ�*�ָ�\��s�y�`��x���N�|z�Qy-p��v虵��֖Gk��>�t�ˮ@��5k���u:�e��]��N��4\�X��[I�N�c����Xj7..<��c���V.�w$kӪ�O�bc`t.ݙ�6{v1[u�IdA����d��5�5J��H[m�N�-�ٌ�CZ�$�����8o|ֵ�ֵ�$���X�4" aJ�����N�
E��p�A�cP����qo��Q�v���+�ݷ����l�%d�:`z\W.��cQ4�Q�3@=m���M��X�x���;�ڮTZ(�Ws4���� ��|`����S-�b��������6�Bm]M��+��Q�!Ww��Xw�ذ7l�<ڶ`�G&YX�0�	I�u�����=nJh��h��l@5� ���ngn;mΎ\��[�7e����͎�l�9�J3w����Pi��x�y�����h�%4�w4�w4
���� F(��� �jٜ���ŀ7݋ �v� �\���F9 ����������h�%4Ǻ�m0�%
��I�X�D(_�U߻�� �~����S@�s@���xS�����07l�?BQ�����ǀ����e4�z����1��H���R^�ڢ��s�G\!�vv�-�n�kq�۶��v�2<Dng�_�'�@���hzS@���h���q����7��k����2>w���ŀk�l�<�ʍ��Ʉ�H��hzS@���i����C6AO��P�������iP��M*#�%�����_� ?ou�i�S6Rj,8��@���h{%4��4�)�Uܞ:H�0��D�s4�Z� ��/Т����?>���7� ����*��D��U����+Z��Zçsv���#q��e��cI�YͣH� �us��w�?m� �����C�;�h���#i����iɠ_t��#�ھ��n���j]�*�+WK3/�GL	�}?}�RGu�4�g�@����LPS$I�J'3@~U�p��x��0=	bQ	TB�С��x еt�S!6���]\�ޘ����j�&���*��ݵ�^ŭ�,��T�2=j��}�����U�ݬ��ˮ�Z�n� ~�f }�� ~U�z"!} n������Ġ�Q`���n����s�����ٝ'N��+��F(����- �����4�u��A�ղ0�r@�Z�ϵ��������?B���[��:�_�	1�܍94��>�\X�s�{]��Q�QJT0 �(�*���R��
B�.�& H|�G[F*@1�#AYB�H��4CA 2 b��X,A�.Ņ�%$D�3w��fffff   �         I��   m�             �7r7ky�7��UU��rJc]&h��.� 6�Lj]��`^Ul��mPӧu�9R���0�B��l�oUӗ�{v�9ظ�\�*�MLn�m�eA7ayKd�!��㶐IIcx�����S�R��BL�̰=���*�؎{[rmT����b`�g� ����*�%eQ���K�*v���8B�[�2�T9�^۶��s���zj�n��gi��� K�(�>��-�P2��ԨIڈ��s+%�U�����uv͗����\����Tb����d��[u�[Jd@c�͹��7jI3����WشN�$�GI��]�T��qtݍ�]��#�N�/6����v,�nM�X��r3q��e��m�2����*6�tiom\��Q�m9�S�[[.��-����N��� <�x����mv0������X�=��J������PL���C�ݕ^,�ٚ(��U�H���n鮧D��N3%J���2�r���̮P6v<��<\�����ɓ.��\��]��[6�Z��*�g�O����Ks��gg(��^��qlrO+��u�C(��َ�eZ�8�˞�*���d��m�h]��iN��=���=P�N����m��Q/Q�a#�vl6X���p��< 6N;A���̮n��iUW�u:y8��i2� 	�/i��ؕ˴HMUP ��@  z��N�ɉf����,�݊ʰ]��Ke"��v�	(��ٛ/RMmu�1����N��m���9���MPc�sgbZ�yZy^�	V�jm� Ul�T��e]��n-ڶ�UW��U�TƶB���$��1�2`d�����<̻mm��ʹ����1�[��8䖬t�[I��t������tq)-K�W.��v��T�F-�l�W<��d%�:��S�gp��������www�P� Z(h >PG�?<Ҥv ��6 �hTB(���;]�ow���33333332@  M%ѫ�nt<�6Є =^�;�1X��Q�a+��9��h��>]����Ë��;ڴ��5����۫�����\	ri�Vɭg:�x�N�R���Y��gau���c�;�󢶛��e�5n�Mn�e��v�l�c<�h���nj��6�{;{rc\�2�nU8�{�c��-��Az�wql.���{��{���g��8L�Վd
9{[��n��N��t�Pٲ�8X��u7)�T�prQ�1Lj&�,�8P;��h��� }�w�
����9�:*��6�I�#s4�}V�{�f�}Қ�or�!�k�Tک	�u7Wt��pz~���0=�0&��L��C���	��
I�_t��}�@�Ǯp:���� �.�S6T�ܢ��Jf�`ޘ��W�0ޘ�������V�U�ۆ7�R�uq.�&�����g]<�q�t�&��}�;�b�s�$ڑ���- �����?ٙ���s@)����F9 L�- ����HxZ�Y �d�"QH�P���D%)BJh�w� ��^�f�����H����@���h���;j�&�J]�ը�x�H�y{��;��� ������q�w9�:*��6��iU�]��W�0�1����&0	]	����nV����S�aFj*�;Iy����|s�ܐ ���5qWK���u�%ɱt�',x��^��f |ۼ^�f�YQ�lq��H�$�:���{��^�f {��tL�NZ�⤫��Z&��wu��[0��^P��_%���f�}Қ�9a��
a1�7$z^�M ��4�)��W߿= ����da�S$4׬�:���˺���M�uik1dc�U��闌��Ziسst�Բ�^8�vs�5�)g� q�6c1�$�-�� ���V��K�Ϻ�:����b��M<RG�uz�����h�����q�����r6�Y�&0$� ��h�\ncX)�%$�$4�h���{u��H��S/U� ���ʢ�L���Mޔ�wY�[�)�u�@�u���m��&4/��'e��QQSE��f�/`�e���hT�.��ز<�	�@�>�@�c��~�C��Ҝ�w\��-R����� �*�9�d<�� �;� =��?B�r���L#�S#�@/~�4�Ji�$�M�׀=T�p�l���.�Uڙ���>�`���7ʵ���+߿M�4�? �1���8h���?DB�U����^��f.�
����sٙ�������fe�x�` ��^4�Y�n��K�<��Tˑ.��@kk������"�3�<��.7����lu�
�����nn5�	�n�Ù���ͤgV0�DAXg�jg�ظѳ�dF��'���s�9�k{:6�kj���&�Ŭ�n�ӹ��i��n(���I�&��nΧ#63��t��$#��e�sjz����q�÷"�����}��v��+q��,�`
{�F�*-۫k�|��r�ݕ�����Z�r�y1���������Z�l�>{l�(Q��wV j;�QV�Q6�%#X�Z�l�>�)�y[^��/uz��TljbɌ�E$�>�Jh�����|�_V =� ��YHy� �N����>�@;��BJ}�8�=(�]�!6�T��d���>S�u�"){����=w�_e�-bQ��rLo!��l��]v9nG��^�P/Om`M$�;����.��9!2)�w���v� ��?ٙ�q��@=�/��@�f7#�h:nsQ�"%B��׀5/�`�٠w4�(��'�z���s������uwN���K��Q)�%1�$�v>�@;����Z�]� �r��K2D�f7�o���D)�w_�o>ŀn��8ߛ?����� ��۹'WZ�8n&5�Ӎ[+��8��mٽvh�x����%�\�1fc ��::`wU�L�L`��T�����wx��Y�(��DUʻ��?߯ >m����n�)�Ly�9�v>�@;��&�>( ���s���3rOw�ـQtEU�ͫ���D%2�����x��X�s�-Z拰�f7#�h�٠z���;��Z޶h�eILm�������c���9j�`:m��v)�����n���LmN���w{����h(��#��;����wc��l���@��&��S$JeUk �U�s�ТU@���=�׀{�d�g�$anT9��H�������x�n�=x��Z� ���eMMʵE����$��BJ�~�x�߱`����B�P�T�w��*4<�8d&1I4׬�;�k� �7x�n������L�L�98��{��{�@336�-a��=���z���������{��t�n��ػu�Y
���;�w���w�6� �׋ 8.��F�H)�Š�f�}[� ��x�s�
L��jz�.�1�ܘ��@=���z���;��Z޶h�.E���$rh���7Uk� �7x�!B��w^�bk��S$JcjI4�}V�w����h�w4f[,�L�I$�	e   :��5��P>���m�Ԥ7]�A��{m{mY���+`�[&���OA�E�����ma���xa��q�`b2����mG(]$���l��!<ƻ$���/&�p08�nj{k��%]&]Ԅ�v9�q�qg�ѡ�t'k�%S{�t&tv��jd�<����Z[��v��r}��]�.p���ϫ���v�������_|78����a:���AT��%sv�vNp���3���u�A���19��H�����߿M ��x��_�!%�j�N�x�2ʚ�ő�"�I�[f���s@���hz٠�v�Ǔ��)&�z�uV�â"!L�{� =�׀}#���Ly��h��� ��h�٠�� �_��M�Ȕ�W8 ���ȅ�!(U��~� ~��x�>�@��ۍ�Q)LS"��[\��4��$8y�E��Z�&�s̻PF3���4�l��f�ݏ���f���X���G&�wﻛ�]+@("��v(PDK�I/�1�}8��x �w�����U�Z���w3j�j�`ʻ� �� �٠^빠��q9��R�3&�p?DBS=�׀�׀=׋ mSk@�{�����,��RM �٠^빠[�ՠ���}cm�l!n3um �Q��S74�u��uwn]8��с�4��=�}�龛��J���?O�~t���D�&ɌI1��DDѓA����[�ՠ�� ����Ŝ�L�����jK�j���� v�^ 6���	��Z�PA��Ԛ�Y�pX�#��t0��z(@����(�V ȂE/�Ut��A4���� #� �3>�}7$�Mw�@=�έ�DF3���4�f��m� mSs�Тg��x�pN1F7��NM�]��v� ��h����?V���&9�'1$غ�a��QM����P˲��n]����ݴ���Q)�%1�����c���_[4�o�_ȏP~��� ��UZ�S6����x��1�I&0'tt���D��{8.ljb�̃�M �٠{�)�[�ՠz٠�v��0P�rQ7w��N��0�>� ����Ľn��D�؈� <�Ȝ4꾉�{d��&07{ ��S���W�׳ЯV�n��k\�q)X��s�����0��[=�K	�-�o�l��=$��d������Dc1�ܓ@>��������[�~4�٠z�pP�ba�^cw��� �Ɍ�L`{�!���"S���ݝ)�z٠[f�{��}�ЎcX���R����� 舅������rO��@�"��
��x8 �@  �F\�l���ӵd,�n99[,u�O+�y�\9�����wێ�v:r�ܔ���|���9���k��v�)Ӭ�Ibӌ��ڲI6��Ӵ��ւ��L���At��݃r�a�W��m�2=�zpy�g���*��om;; k�]�24����Sl�t<��>&�Y2��+A���<��]��[�I�u�.��ML��s5��TS��x��%]"[�g�j)u7Df�s/YB�������wx�q�n��VD�Ɍ�E$�����{�)�wgJh޶h}��lq��I�rM�]�uvA�M�����	1�A����wgJh��@>���]� �W��J19�ZvL`�cwGL꾉�z�t�1DF3���4�l�/u��;��Z}l��ܕk�K$Y$�.Mn'n�!��ֺ�Iy鰪��m���N3F��v�AF(���94�w4�}V�_[4�l�>�#����"S�HnI�ƾ���CJ0��"�@J��	�c �Ɍ�0WT��J�'28E�E��f�}m�����o���w��=�๰i��&2DI1�zI��} �I��-�1�������ݏ���٠[f���u���Ba�saۧ3�շet�4��+`�Z��K�^��B"$Dm)��,q��;��Z�[4�l�=�w4��_��m(���m]\����DB��wu��b�;��Z�vul�"1�܌NI�w���?}�vnq�"@?����h�٠z�pP�5�d�F�GL꾉�{���&0=;��1D�H��F�h��� �����h��;��&�L72&݈����ʌ�U@v��o���c�!v^wJ���M��X�2LSs!�X�^ ������������W�06���k)Vc!$�@>����s@���h�l����1��
&1�4w]��U�u�@>����I[J�J�Uuk��RڷӀ}׀6�r|"<Aڥ�=TG}���`<���m(��jdqh�l�?��(Q>���o�`�������Qp�	&�%��y�'X٣����-����7':3ZZ��p/�����Nw-v+��=�׀{u��7Uk� �[�Ί� �5��M��s@���h�l���@���&(���ڗv��Z� >��IDL����5�����ܓĜ�D�)�}�� ���0;��&��!�j�T�T]�ww�6� ��������}��ff}gY$�I$�I$   M��y��.!���:��ێNzM��n*pi�Tg��<���L>�s�6_�k�77��#�YB:��7�i5��m�e���In�հъ�h��<S]��C���k[ j:��똫r�7nӔ��2��Sb�+&*;d��5�npf�Ҙ�[P7ݛ;���y��nC��>vۋ�,z�7n���uNx4��1�&��P��7�ֵ���:���u�v�8�Z��t �g�O^.��i���hT����&\�Ź����OΘ�} �I��L`yBRT�U3j��U]Z�<���~JJd<���w~�4w]� �+�SQ�1�V+�`�1�nɌKd����D��nL�@=�f��׋ �7X�J"gϺ������Bx̉ɠwu��=�ֽ ��4޶h\�X�sMd��18�d�.�-:q#�_��}����I�:ܛW<�W4a1D�H��Ԓg�v.����l�y���(��A�ذ�k�U��3j�q^|+�`�c�$rc{��ҝ^���R�`�Q�BI&�w���^,9(P�e�]Ӏ}׀[��eQWA6*�����P�R��ܩ����@=m�˱%]�M�cD�yL� ���1����6��;���e5!Z�uIR;��lˎt����6�Wi=����C�ﻻ���`���1��$_ {���@-�4>AquP�T*�Dc1�0RM �mX�� ڭs�n��P�Q2{��� �(�قrh���n>�s�P���&�C��Mw?f��f��Ia���"S�I��Z� >�w��P�B�7�, �~����L�q��Z�l�z�����}V�����X�#4:ݻ��y�)�73�\���dՂ�\�ݛ�f��ù�&1�A��	��Iɠ�������� �h��,bbQe]U����,脡D�ܩ��}׀��.ė;�JcD#��[��0�1�I�$t�%j'�b�&誻�V��p:"Q2�u�s��<�Ł�P�BIGDB��V�p��dQ���dRM ���-�M�}V�[�h\����$O#l29�!Y0�Nk���v)��k��n%�v3f�ƻI�DĦ	����)�[���z��$�G�s���|��&�fH���n��� ���z�ޔ�as�&�&(�1H��w��9(��3���S��5m*64L'�$�z�ޔ�-�j�z� ���X�651(����)�[�ՠ�4�f�!y�
q]p�]�}�J!�d$�"���Q?/Ȑ"`Ń#(�DhA A"@�%JD�j�Y�+�]+(B�R�� '��"�~�4�p������ Z�8�`�"@a�D$!	���J��D��b��5�M&��1��R���XE	�ѣ2�����4��I#�THu*�0���Ca��p�i���Ā��H���o��3330   �         ��   �`            R�aT�Q��V��B��BȜӄЭMS*��ɤ��X�B�t�ό )����j��ꪮU�W��f(��-�8{i�u���U�$]P�.����cvrb��Uei���;眝�;N�,E2W��=93^1��aV�s�5��=�=��r�m8��%is���W3�	u�$�����3{j��8g<c��J�6�N}����&wV�FE.���56�u:��
vm�*�%A��k�l��� ,5j��CJ�rk0��]ˑ����@P��dl�z�v�M�@;�53h�m�k��0b��ȵ+�N���m��H{v��"۠+�D�B�>�u�]#���Cg�UuRJ\�#&���Q}��k��LC�h��U���\�]�WOd贂�Y��V�յΓ	4t���O��k��@�k�n]����5�3Į���� �W��`�L�%jvڷj��,F���@^\S�������r��d{lEvlZ؝�S c���8�zK�YÃ �3l�(����q�=��(��p���i^��bn��e)���q���)K���^v:(�SY$��H[r�U�;vZt�Xݢ�U�;S;�s�E.�6e�8��m�2�T�b(+�Rٜ�-/i.�N�G��Z��A��M)�,u ��U˶�h���� /�!��E�h]6�F�k 6Z'v'Y.����l�Pz�:Y�m�Pb@{eT8�.Cc�U ����$�-��h�[���\�q�k� �n6�Z�U����vW�ëm��c"�6;�L�͌@%Nwk����ovBm��� �ڀx�K��k9�t[��㝤�b�X�z8(�����Y��v�<���v�]�>���~x6��Z[�,
N����q���T�7S��6��V۶x�U]e5�3Y��W4[sE��Dx�J��¡( lTM��i�>=�w����{���~� �6�  �e��P��m�˘=��s�tN���@���Vأq�v���5Þ� W2�Ҁk1��t�o���o����Hb��g�l��+���r�kq�Od�s7ۆ���0��6�'1+P��ȷ[��H�&%���h����+���k�ٕ^'gn�,�l;���5����� �������-CS��r�-ՙ�O*Ѿs5�jYm�Ѣ�F%�Dlr3he�OGY�+:��������ﻻ����?NT.Mc���m�����}�[l�m��S@.y��J2��eZ���ۼ�$��!��xw_j����(IL��>�.nK��UwE]]�wu��l��DL�*� �~�4^�<�)�L�NM��4�78�n�?%
"g��x�/����m]������7Uk��P�����~��h�)�vs䫀�1&9:X�Ѷ��Ce�U%���x�vNq���7=/n:�aE0��&�&(�18��l��Y�wt�����h�J��Mu����ܒs�w7EN*��;�� �S���w���	)��S,�*��
Ф��~4�>�@>�� ����ė;�51b�a4?B���泿N o��x��x�m��Q��H�Q��"dqhz٠^�@��M����*�um��H�MɻVwNJ��j\,�Ll��3���E��3���"eh�`�dQ���brM ����x��s��{���t���S��I�w[��w��Z�l��Y�}x�0�� �8ܙ�w��n��{�������a���EI��r}��7$�����<����S5j�u6��p?B��g{�c ���0;�t�����!�i�a?��)&�}z����{U����������)�mHiDfj�zy����nq�!��3�g��N����cX650Pƅ$����������� �����J��51b�1ILھ��N��L`N�� �V�5#iF7!�2H���@>�f�z������P��Dc1�Uwx��x��`�Z�R��(�QP�(��u���H���͢�7w�=o�U�s����$)��y�,KĿ��fӑ,K��G��}����- N.OEǰ�v�i�Ƭ�a��ca�9�O<�ٵy'H�tuJ�n���{�,K���w�iȖ%�b^��ͧ"X�%�{�ͧ"X�%����ND�,K�N�z�a4[�0˩�Yv��bX�%�}��r��Q5Ŀ{�6��bX�'���m9ı,N����r%�bX���OY̚��	���33iȖ%�b_��iȖ%�b}�{�ӑ,�����{��9ı,K�fӑ,KĿ|[�=�5����Ys3iȖ%�b}�{�ӑ,K����]�"X�%�{�{6��bX�%���6��bX�'�x��^�.���i��m9ı,N����r%�bX7���iȖ%�b_��iȖ%�b}�{�ӑ,K�҈�}�~��3 t�  ���aª�h㫞��,�je������q'�m�8�:�ܝF�V��{t�GZ����!q(ף:�^�
bm����n�nr02]k�\ZY)�Ů�����,N�Ǡ̫I���2p��ֻj��n����ͼ��g�'�x��M�5U�`����+n�L�G����f��s�5\9z����hY��3YnHK5�jja&��T��T$7�U��Ƨ^�:"�v�=wkbbMq*u��n]8ь����v�ִ؝!�~Nı,K�����r%�bX�����r%�bX�{���Kı;�>���
HRB���E��tP���ffӑ,KĿ��fӑlK�����"X�%�߳��ND�,K���m9ı,O�����I&\-�kD˙�ND�,K�{�6��bX�'~���9ı,K��ٴ�Kı/���/�RB���ٝb-M�j�(�fND�,K�g}v��bX�%�}��r%�bX�����r%�`؟{���Kı/��g��E��	��u�iȖ%�b^��ͧ"X�%�{�ͧ"X�%����ND�,K���
HRB������]UL� ���O4��x��US��
�kǅ�)�t�W��q���MYP�^a������{��2_��iȖ%�b}�{�ӑ,K����]�"X�%�{�{6��bX�%��^��I�M\%�j˙�ND�,K�w�6������C"dK���˴�Kı/����ND�,K��}�ND�,K��m]M\)r�Is�"X�%�߳��ND�,K���m9ı,K���m9ı,O��p�r%�bX������kV榵�	33.ӑ,KĽ｛ND�,K��}�ND�,K�{�6��bX�'~���9ı,K�{o��r���5��Mk36��bX�%���6��bX�'���m9ı,N����r%�bX����iȖ%�bS�ݷ�֝I��ӭX[u�rX�m�(Ea����s���!��ۛ��^5]qsʡm�{E_{���oq���}�{�ӑ,K����]�"X�%�{�{6��bX�%���6��bX�'��o�	��p̚.�k0�r%�bX��;��Kı/{�fӑ,KĿ��fӑ,K�����"X�%�~'{=u0�-�L�ˬ�ND�,K���m9ı,K���m9���DGX*PA�$�:Tٸ������ND�,K���iȖ%�b~>{�˗ZոLu�Y��ND�,��}�ND�,K���m9ı,N����r%�bX����iȖ%�b_���Od����\������Kı=�{�ӑ,K����]�"X�%�}�{6��bX�%�}��r%�bX��{����6�͎�vzsQձ�����l�ʖ�tV�-��/=�BmmU8r\q�s�"X�%���v��bX�%�}��r%�bX����iȖ%�b{���"X�%�};��nf�njk3)&fe�r%�bX����iȖ%�b_w�ͧ"X�%����6��bX�'����r%�bX��I�kS.5,5��K���r%�bX����iȖ%�b~��iȖ	bX��{�iȖ%�b_w�ͧ"X�%����[<jٗp��f����Kı=���ӑ,K��s޻ND�,K��}�ND�,N`
`(�D�w�ͧ"X�%��ޛ�Bar\3&��]fND�,K��z�9ı,K��ٴ�Kı/��fӑ,K��}�ND�,K���{������a[�d��垚9�ӕ)�����v��|��;�6wJ���L��;�������h�Xe�&fe�}ı,K����6��bX�%���m9ı,N����r%�bX��w�iȖ%�bt��N\�֭�a��Y��ND�,K��{6��bX�'��p�r%�bX��w�iȖ%�b_}�fӑ,KĿ�%�Ԛ���ܦ����r%�bX�}��m9ı,Ow;��KKĿ���iȖ%�b_}�fӑ,K���[}��K���.[��̛ND�,K����9ı,K��{6��bX�%���m9ı,O���6��bX�%�痢��չ��fBL�˴�Kı/���r%�bX����iȖ%�b}���iȖ%�b{��]�"X�%�S����{��_����p 	   �l��ݯ��7�ED��N�r%hN�]�ݣ�=��m�=M�5��N����7�C�R���h6�q�ڀ��\�Y�ꌕg��hKr��j�˪�����.���X����:���W�ؾ�y �@�݅�#�Mi�f;�ۚ�f�t=�0���1:��f��qD����נ��!�Xҹ�3؃����~���.�j������P���Vtӱ�h��-��ɝNs�LBQͷg��b]Z��w���oq����{ٴ�Kı>���ӑ,K��s޻ND�,K���ͧ"X�%���wg�ճ.᫢�k3iȖ%�b}�}ͧ"X�%���v��bX�%����ND�,K���m9Fı,O��߲��5f�����Kı=���ӑ,KĿ���iȖ%�b_w�ͧ"X�%��{�m9ı,K�׾���an��3Ff��9ı,K���m9ı,K��ٴ�Kı>�}ͧ"X��5�����ND�,K����˗ZոL52k33iȖ%�b_w�ͧ"X�%��{�m9ı,Ow=��Kı/��ٴ�K�7�{���v���*����3؉ĺl�3���i��cq1dx�Dmi[�0N���r��j�g�I��؛�H'~�{v$�H<����OD�,K��ٴ�Kı?ze��5.���n��fӑ,K��s޻NC� �ʀ�@q�Mı.��fӑ,KĽ｛ND�,K﻿M� �6%�b^ώ�ۗ5.jkY��32�9ı,K��{6��bX�%���6��bX�'���6��bX�'~���9ı,K����je��u�����r%�bX�����r%�bX�w���r%�bX��=��Kı/��ٴ�Kı?{�vx��e��5t\����Kı>�w��Kİ����r%�bX��}��r%�bX��wٴ�KĻ��~w�߲�]C6�2���p#T��닋�������/&�Zv�Kt��+�5f�ֲq?D�,K�����Kı/��ٴ�Kı/��iȖ%�b}�w��Kı/�o��L&�L���̻ND�,K���ͧ"X�%�~�}�ND�,K��~�ND�,K�g�v��(%�b|u��L�֭�a��Y��ND�,K���6��bX�'��p�r%�����-�(�F���C��M�]�]��7�1�d)1$���!
�B��
@�J��0�
E��� ���CQ�MX�
�X)
�k�T"%# %�L`��14�$$B��"0D�,!� �@�"�
���b��4GBD����>	�j��!�T�DRBa ��d	1b� ��!�c
��K@�K��F2��`���8*P@�
� �
b� qP E��� P8��O�n'>��v��bX�%���6��bX�%��ޚ�I��[�˚�fӑ,K��}�ND�,K�g�v��bX�%�}��r%�bX��wٴ�Kı?k��{3R�j�K��0�r%�bX�w���r%�bX }�{6��bX�%��{6��bX�'��p�r%�bX���j�j�浭k�LȔ��l٣+0�]�[e�5��dB���
Z1�|<�c��(NZ݂��������ou�}��r%�bX��}��r%�bX�{���Kı>�w��Kı/���_kS.5k�f[��ND�,K�｛ND�,K�{�6��bX�'���6��bX�%�}��r  X�%��wz�xճ.᫢��ͧ"X�%����ND�,K��~�ND�,K���m9ı,K���m9ı,O����h�.�]ܹ�ӑ,K���ߦӑ,KĽ｛ND�,K�｛ND�,��dN����Kı/���ja0�d�fd�r%�bX����iȖ%�b7�}��r%�bX�{���Kı>�w��Kı>���kZ����*u�m�1k:���n�-���hʛl���7��G�z��
���U������ŉw�ͧ"X�%����ND�,K��~�ND�,K���m9ı,K���}�5�\5�e5sZ��r%�bX�{���Q[ı>�w��Kı/{�fӑ,KĿ��fӑ?����=�����ݿ��p�����Kı;�o�m9ı,K��ٴ�Kı/��ٴ�Kı>���iȖ%�b^Ϗz˙�[���d%��6��bX�%�}��r%�bX��}��r%�bX�{���K��T"�j'}�M�"X�%�{;�K��L�\ծ��nfm9ı,K���m9ı,O��p�r%�bX�w���r%�bX����iȖ%�b����33330 ��  k6_"�f�;����|b�9FܖY��{H�t��C�'����VwK�����lz!�z�s۴�t�m�X ct\H]�p�b�up�J������2c��g����y�3�WG%�m�c��@�]�ɛ���md�v�nps�v�;i�`���T��m�5*E.7��S�h�䞜n�����`�۷��	���mv�:������U��{`��8�
I�0�5���9�U��qv;�5q��d�jZ�5�h�.G��������,O�����Kı>�w��Kı/{�fӑ,KĿ��fӑ,K����^ue�p̓Z�ܹ�ӑ,K���ߦӑQ�,K���m9ı,K���m9ı,O��p�r%�bX��w�50�-�Y.I32m9ı,K��ٴ�Kı/��ٴ�K�j&�w����ӑ,K�ｿ��Kı?��˭j�&]f����r%�bX��}��r%�bX�{���Kı>�w��K�FĽ｛ND�,K�}z_jMkW�f�\ֳ6��bX�'���m9ı,O���m9ı,K��ٴ�Kı/��ٴ�oq��������쫰R��7 �0���D�zţ�����l�Q�9ZK^�C3R�j�K��-ְ�r%�bX�w���r%�bX����iȖ%�b_���iȖ%�b}�{�ӑ,KĽ���3Z�55��Ks2m9ı,K��ٴ�<� _ �N� ���X�%�~��ND�,K��m9ı,O���m9ı,K����ֵ2蹫]k2���r%�bX��}��r%�bX��w��Kı>�w��Kı/��fӑ,K����[<jٗpֵ.\��r%�bX��w��Kı=�{�ӑ,Kľ�}�ND�,K���m9ı,O����V\��4h�3Y6��bX�'��p�r%�bX�}��6��bX�%�}��r%�bX�����r%�bX�>�ߛ��s���C�o:5,mQc��XS7h�aݩ7l��.��Ø����si�,6��bX�%�{��r%�bX����iȖ%�b{�o�iȖ%�b{���"X�%�ӽ���u�[�ˬә��ND�,K���m9ı,O}��m9ı,Ow���Kı/��fӐı,K��t������Y�W5�ͧ"X�%����ND�,K���m9�b��b��q7�}��r%�bX����iȖ%�b~פ]M\)r�Y-�ND�,K���m9ı,K߽��r%�bX����iȖ%�b}�{�ӑ,KĽ��z˗5.jk3)s�"X�%�{�{6��bX�(_w�ͧ"X�%����ND�,K���m9ı,Oh�}�fI;�1�5����g%e���ڜdl���n��>��9�z����zPܴfӑ,Kľ｛ND�,K�{�6��bX�'�w�6��bX�%�}��r%�bX�}��֬˅�kZ�˙�ND�,K���m9ı,O��m9ı,K��ٴ�Kı/~�i�bX�'��z�.K�d�4\��6��bX�'�w�6��bX�%�}��r%�bX��wٴ�Kı=�{�ӑ,KĿ��fE�k%ɚְ�r%�bX����iȖ%�b^��fӑ,K��}�ND�,�P4���\�>�}�iȖ%�b~>���˭j�&]f����r%�bX��wٴ�Kİ�b�����6��X�%�����m9ı,K�wٴ�K�����~���*�,u�+�h���'����c/O1W\<��/Pq�8x�\vi�r�5ӥ֮Z���fm9ı,O}��m9ı,O��m9ı,K��ٴ�Kı/~�iȖ%�b~׉�f����R�ֲ�fM�"X�%�����"X�%�}��6��bX�%���m9ı,O��z�9Kı/~/��'5��}��oq��������ӑ,KĽ��ͧ"X�%�ｿM�"X�%�����"X�%�~����]J�_{���oq�������m9ı,O}��m9ı,O��m9İ?�������iȖ%�bw�ީ�j̸[���r�fӑ,K���ߦӑ,K�����"X�%�}��6��bX�%���6��bY����w��������� ����I,�gk��uΦ�r���:	n܆ձ�큮ɔW�K��.����إ(��R�:��օ�Vlm88��1p��:�^�t�K�m�*qp�c\B�<�׭��Sd��5a�ʩyЖ4�\8��mm���s�y�r�������Y���k2Ny��q �vݓ�g��غ����9�Νҫ7�����e��O"�8^j�k$�Ԛ�v�u�"��n;����j�`eۑ2A����k_q^���b�][<���w���d�>���6��bX�%���m9ı,K���6�O�5ı>�]�"X�%�z{�_ĘMᬙ�-̛ND�,K���6��bX�%��}�ND�,K�{~�ND�,K��ߦӐ�,K�{=yr�Z�	�Y�336��bX�%��}�ND�,K�{~�ND��Xj&�}�o�m9ı,K��fӑ,KĿ���ڒ�W�f�\ֳ6��bX�'���6��bX�'﻿M�"X�%�}��6��bX�%��}�ND�,K��N�5e��.��k2m9ı,O�w~�ND�,KK��ٴ�Kı/���r%�bRog����$/R��UWH���]v0v}��vWUCQ�y5�X��ݬ2OC��i�����'5��������,K��ٴ�Kı/���r%�bX����� O�5ı>��6���oq�����W�:.�3���2X�%�}�fӐ�L���� �9��s��ND�,K��~�ND�,K��}�ND�,K���K�Z�.�j\����Kı=����Kı?w=��KKľ�}�ND�,K���6��bX�'����.Ja�M5�u�iȖ%�b~�{�iȖ%�b_w�ͧ"X�%�~�}�ND�,K�{~�ND�,K�w��&E�k&hə�iȖ%�b_w�ͧ"X�%�~�}�ND�,K�{~�ND�,K�s޻ND�,K���o���p�4�an�͕��}���VGm�y��;G)ۇ�������Z��
he��ͧ"X�%�~�}�ND�,K�s޻ND�,K��ߦӑ,KĿw�ͧ"X�%�=�ǵ%֮Z���fm9ı,O}��m9ı,O�w~�ND�,K���m9ı,K���6��bX�'�zN�2˩��.]k-��iȖ%�b~����r%�bX��{ٴ�K	���,c� ċ"F$Ī���@�!�"~�u��fӑ,K������K=���~�~���	�Gik}��oqı/~��iȖ%�b_�wٴ�Kı=���ӑ,K�Bj'��?���oq���������zPܴ|��bX�%��}�ND�,K��m9ı,O�w~�ND�,K��{6��bX�%?w��Y��L̺34�5�[�to6�r�Vz9�2��
0U�smM����~��ݪ�>�4\+���w�{��7�����6��bX�'﻿M�"X�%�}���ND�,K���ͧ"X�%���|�˒�fF�f�Xm9ı,O�w~�NC�:���%����m9ı,K�}��ND�,K��m9ı,K��{$�Mᬙ�-̛ND�,K��{6��bX�%��}�ND��Xj&�{��6��bX�'����ӑ,K����e�ոL�f�3Z��r%�b�X����m9ı,Ow���Kı?}��m9İ(��P@�Ț�����r%�bX���ڒ�W�f�f�����Kı=���ӑ,K���}ͧ"X�%�}���ND�,K���ͧ"X�%������Vܺ��óۧ-��D)�h|ܝYR�M�#���g\��[5r\q[�a��Kı?}�siȖ%�b_w�ͧ"X�%�}�f��Kı=�{�ӑ,K���{ڗ3Z�55��fj�6��bX�%�}��r%�bX����m9ı,O���6��bX�'��m9�U5Ľ﮵����F]Y55�n�6��bX�%���ͧ"X�%����6��bX�'��m9ı,K���r%�bX��w5/�j̸[���r�fӑ,KlOw���Kı?}�siȖ%�b_w�ͧ"X��	5_w�ٴ�Kı>�������ֳW0�r%�bX��ﹴ�Kİ�F���lI�?}�bn	 ���ٱ$D�T_�T_��W��V��*��"��������qW�T��T"�� T T"�$���B* �@(�T"�P��P � F*� P�DX@	T$P�@@� T AP��P��Q"P��T" 0B*#T"�P�*�B� T (1DX(�B
$AP�P�AP�P D�P��� T ,AP�$P�$AP��P�$T��P�AP��P��T��T  �B ��"���򂠪��
���V��*�T_�APU�AU�tW�T�h(���
����*
��*
���(+$�k=��>�A��� ��������[Ϫ��3�.�R��)@ZeS�������h��w� �IJP�� H�UJ� )� P AT�|@����ƀ �(|�#���t=Z3��.�li�{�{�E�������     0 Ї}��<�؝C۵�
>��Q��U���͸7�A��gT��P�P��5���8Ύ��<��t�hz}��xWѦ�d���
H�l�v��i�]�rpPPP���GF|/��t��T�]�}�놄�=���x� }���<�B�����B��]j,�џTgG/�Ϩ�hh4;tW
�MC��x�
��x�opt4��=n�p�i�Vz5����ѭa��_GO��]qD     0��%) �14d1F&M d���R��P       =��RO����ɓL�CѓM�i��)"��F� dڌ4� $A2�&�dLI�<��y&���G��i�
��$O*�C ��L1h�O`>��S����?8)��d~q�Wઢ SK�_z
(�U��́�&��_��Y���b��?����9��H�)�U������a����>��c`K>���ñ�꾼c�J�}7�����{�z��� ��o�6� ܃=��؀/b�=�.�
���`pf���cz��`�p b��b���b(#؊��=�m�p1��{��5@��]ߴr��ٜ�Wwx3Y���Y��{����w}�s�o9�s:s{������www���������]��9ywy���w��}�{����7wn���9�33.��s����f�����f�333.����wv�3L���[�7wwwwf�����{����������f,�����y�ײ�����������+./��V��������V�ML_�S�0e(��~iy��'��!=A%�9ة
i�ШL�ͅ�Y�o5�2�z�JIM)�GM"�M<�3�#|OM��/�E{��zx�*�1��ʶm�_�ׯ�}&���[#!U�f�g�f�J��g� FG�ol�4n�g���V�'F$3$��rar�cKf33�������й�w=uۥ�If�)IobЌbB4YsV2ZzC���\YG�O��N쫎8Ӎ8M1V�� ��N�t��ѨR���ׅZ��>�>�ŵ�[R�;�!�#p�ml�ֶ�m2ؑb��6-\�B���[(�D�"��m�mL�>Ɛ�laK
U�̚v��2h����Idi��Mɔ��A���� �H8(��Z��sZ�\���a(�*�2b�ZJ�
2h٬��
/!�&��m#I`�.�jB��u{H��*�	VY*�x2hؐ�����4�^q�f��I
!�=	t��u�����a`�C�f	#V1�%fMf�E�c4�"�(�$�d�ƖQ��r/[N���zNZ�$�vpz|z��N8�<ox�\ˢK��`'�Ŷ0)�����23��q�tယ��f��?+����*�l�F	�C������
���C�),h-���j��(�Q�Nݚ!�)�c�)��M�`�XU�!�8�w���4h۰�(l�~/<�o3���N;x֍8y�@a�<@[ø8ou�W�D�%�xof��H4�"����d#Yi�M`�( �����r(G.�0���F�F�w�e��E��q����ř5�xΝ�cX)�4��p�
�	�a$�+��ٳ9��f4��,aNA&T3�1��̼����S@BD!Z�i1�c��E�]d�yH�]J���W�<"�r	��>�b�aCV������XMf��ӣ�]��:5�Zք�}q���V��&�zz��<IgC��B;x瞚N:��^�[.WW�S�IΝ�����7�޴�4KU⌚V[��,1(
0�"�2�,s���Bc>	<5AZe�@���E��,��!l�y��]��̆O&�M#H[�Ć���m5��G{hD�c-JX�!K*�&�g�����!F���;Hו���泬]ya��
ƛ�!=h�Z��O��&*�C�����(����;KcZ��wէCUE�O���{#G�PF�9���F���`;Vv�x6N�h���:��S�%�<ӗ<"���i�[��Q
HTÒ����Z2�(qV�(뵻��:u9�W&\�:�-��K���\�4�ȋ8�,%��\W�צ�HY����������P�oz�{�!�i�{!.9Әy���!>�Q>���-�[�Ni���p�w�÷(_���$ݭ�}{�7��׹��qş'�C���?^���G!���5*�.���thՅ�]�m! �x	Yh���.�Ϥ����z�E���]����ر�����<��%�l�a��B0�ʰ��a�.$�//�@�@�:��v��{�����ۇZ�6�WGH�N��}��H��zo�޳t�,:w�}oY�X�q��9�dF[�G�M�m�g���ɚhV��5Ȯu�u�������^*���g���Q�hlԙn�㥥��N4q�hHp�n�����d;o���:;<��B��ta2��,p��$h����*�ăI[�J�+SFL9�JM��(��A�Cs(,� 2\gu�^^�ك�� Q��^!��΍Dh��MXb�t°b��xte
U^2h�0`�dp�d�
4l�[�Y[ɥ�������eN���e�jͪ��R���G���#�R?v�������6��[��x���r꣯�f����=��1-[�؉��&��\�w��I�ƌ>����Q-Co�� ��im-Jo�p{�����+`퐗�ק�?��=8����>�{�5��,��j:�������V�$�H      ��    h      ��H�� l �`              �=                                                 +4�9��!�<��L�;����{t�`8�NƎ-�ݱmu�X` �m�[�3Yn����� AU6UJ��K�R����b�VՍN��xp$;������6ۃm��n4��MU���(��J�'�-Soꇮ��` l  � p��M+ ����v=`Uj�Wvc�$[M�m,�l� � 8 � �6ؗ�y;U�@$�O m���F�Kn���H�v\�m[M�@ �	lm��ٶ��̭��M�W�g2M�*���ns�$ ��hڠ�4�TJ�����m��@���m�E�	�����m��/�i2N�Ӫ@�nn�]���M�9�BV�R[n(
��U�3�v���i(;������HU+ۧG7m���;�:����h�����t�UH� �6�v�m�`����B�6�� ��ֻ6��6�� n�-�� ��l$.�\m���d�mS���l��8qm � ��=  .ˀU�8jxSD��
���;m�-5�޸-��m����I�m  [m�ۀٶ �`  �p�Imp�kp ���[s���Vؐ ��8H'm��	[AoP-���	� m�8�$ -�� l[m���u��f��H ��6�� I�$h
���� ��<�����4�  ,�e��mU*�R����7� u��ݼ�K$�MI�i���lHl �r۝Ey�ʲ�W/^�j�V��=�4���ۭp��f5v��e�i��������Ԅ��ۄ��   -�  �f�I�� �m� � Y�엥.� �Y���=�v��B@ !�� !�͖KT�bڐ�tV�Bޠ����N�u��(WU8c4�`G���{P�ᶽ-�9  
T��7l7Pڐ%���] ��h��b�$� h 6�   $[E��η`�66U�i����6ۆ�Yvu� ��rՍ�UP8qYR�mf����
kt�N� !��UU�iP�#�)��;.����l$ 8  :	�: -cj
=��M�X�$c�����5V��[���l�^`[A&@mpm�Cm�� �m�Im   &��9��6I����v�sm���u�o2$䲁������ ��5�m�����[���([Cm�ʐMUm6�6 ���l�z�m�Im헭�u�HԠ s��Z��h��� 9'8�5Ѷ�Y���1�m���T�Ғ�	.�UJɀ���ݴ����k`6�[;UT8�V��e��*u[���G*�P p�!� ����Sd
�8*�jڦհt�� *�Jc-Um��ݶ�-6<s�Iu���մ���ru� m��C��N�8�sUR�n��l[T[f+b� ��  l�o 6ӳV|(U�X��R�>6�   :���m�[J��@� �Rm� 8a��� �]��gM,�+  ���  ^��yt�����	 �$�h&Fs��`l�     8ktm�[D� H  H  [E�H�   -�  m��t��=w������-�i�Ŵ� [I��l��U�*���$���5�d�˴��-�l �Qm������6�$Ӝ��ݵ��V�l -�d�`8-��m� m�m� ��^��l �`$�	�lh:-�  [@  hH   ��` 4P �� 	�� �  �mm�    '%( 	 �6�-6K��  ���I2�Ӭ�dq������W��P ^�\�u� �Yg �Q����vV:���� ���-����T�(�m[���;]���Ͱ  '@u�i,���m� k  f��ib޸%]�PVӈ�j��n�6�����	�m�$6��U)*�:L�7J�H
�I� ���6��A d|Z�}�H�k�^�ޅ��g;X�(�ϛ�/��U�����p����{7;rtK,�W����� �����0���W)A�?���6�=���±�e�T�q�r�J[�*W,qQ,��K��6�BV��[V[
�� ���E~@��TOaE�<@����W`t�Љ�t�PT��
��P<p�%��Qp�P hD4��o�[PS/����i�b(P�;Aҥe2+�C���, T��lD��H�- <�ZPO4�"o��q_8&S�B,A��Dh���^*����$%��͕����&�؉�C��~6���i��-�8\(j�@"P"&��BԵv��'�0��R;w�����2*�������r*�����򪪪��*���������*��dUUU2<����������*���������*�*�������*�i4�I$�H�M����P  ��� �s�}�jM��{�����{;�>X߾~%�Cl�ƙ�y˻�Xh{�z��6��}����#�7�]#�w>�|�d�|�UU�e@ ڶl�  l         zt�nYd��A�õd�g�����l�T�N<JQ��n�T��Mj�nݥaq�ͱ(�V�;��jB�J�3��m��c�eݝ5NG��C�
۬*gn��h�ex���k��sr)��1�t����ce��B��U��v��a��nQ.k�����p���n�.t�%-sv[tY��f�0���e-�i^<�l[Vp;N���tx�E�9��zP��@GkX��^�D�N3��V�Sevum�.���ʹt<xޮrv��!�D���5L�gd�l� %��@�UX;K���sę���^;-��Gm����	e�(	`̭%V3m%�mAU�lk�c)ۇ��U��j�h����e6�s m��D�����]�68��M�x̤��]AӺ׻��>�Om��Rj:k���:�Э��ԧt��j���yU��:���������UX�J掄K�≲�Y-��py�ɚ'�����+Eʼ�wd��"�!�:��i�L|�C ��:I>���������ͼ��ʪ��g��ѳR��b4���\��3L�Z�q�C���sŮM�W%˃Pb�j�^�k��dNO<ggk7`Ih�ԫ��Çy���K=�֛�̓�s�ki��߼@OY�ݻ��c��--��Sk)6�كj4��m��n���8��h}x��UDfu�ieޑl���냼��X�e�=�c
-Uݰ;ޱdv]NtX��N��m��u����2R�B�{b��}u�	�l�q���".0P�(��x��[�Ne�)[/w�?;���W}b�v��24#kB��΅�G�zf�C1���O��}Vz����&��\T��b�ë��{L8���[b��]����l��Ho1�k��:��W{��bG�4�6�L��Ѱ�юClh�@���7v�۫ +�6F��bD�)Z�t8i]�.�]��J�f��� 8�۫�u��ElƫWlo�uw�V@r�j3#J=�u��:�J�����x���V�lԮ6�F��D� �P8�Q�ݺ�v�ݰ/gw�aD��,�����LY���������fu՚�akdٚv����)B���j�a���%��]ܮ�nػ6�
�p����D�n�^�Ł�L����`�f([�ꧾ1/������(ن�vƹ�J��N$Gu�|Q�Q��˷\�;*�=K�G�a@�)G\�u�J�~M���1��y�^0UU�ȧ"TV8���{`�ZB �����^�I�N!��s����E gm7[!�w wK�5�wZ�+�kdc`@j�n�yכ:Ƴ�ssЛ��!fRn6(Z�:R��=�j���y�m��U�E�����A����12�b��i�q��tDn�S��\?�]Ɋ�����w��/�^X/ /p��I����^s��������;jf!�!�8t�*�V*�s�X.�-s�j<�,�o�f�S�b��^@[�uB��Ub��of�Q� 0�U����`����L琪���L\�rL�Ya7+��J�͒t���\�K��̨�]�y`����,�p�\�ˬX/9�`� ���)�$��Ö����PS���pK�b� ����k ��,��q�癩w&*zX&�z�7������+:�b�c*<�-�G���K1�
�#��4�m7)D␈�-\KM� ��|�����N��r�wk�Z�9��|�*`��1R��@@�"c~Z�;��{���/u�����j:�����4!�
������^�fF���}�ߛ�����Q��+1r��y`���r�xs���'/ɉXi�Y7d!�x��T̹x�����^Aysz�s��n�q�癩w$Ā��mGz݂���^E= �@�zV�$��� ��l�7`����X.7����X��<�]�^_,S)�x�����]�[�0b�LVQyuz�A'9,�ݨ�[�bYw9�sO,R��zpzz�6q��l�U��P�s�UU�V@��u^�fF�3UB��0�C��0^�w;���"jV�U��.]b�y�,p�ʵs��ȤѪ�0UbLU��7�Q�8X;��;���U�y��rb�.��Q޷`������7�|��[=�$Q� ����vԦf3�,(`��u�9(�[M���]	k��U��I���ޗ��3�^��Mh�Vl&��A�M+]�0#/]5]� Ն�����|gu���{B{qh��˛�v��(ESz����&.�+*<�,�7,����~rLb�b�u9˰]�^_-G���>np�1��YE�E��XQ�9`���G<��p��]�@^k�����y�� �����W����^Ty�Z��ߞXW�S�uB�����$$������5�(���T�����\8�ł眰]�Z�,39�X/77�\��d��;R�/{�sV�yjr g��<�˹1P]��[�j#��`� /1³�&.Uc*<��ȋ\�b)7�$1��5��^s��\��K��g&��ۘX(D�l�k�b�16��\Ǹ�`���N��N�w�{`��)Q3�n�b�.� .����5����{�{���b�yQ�9`���pT3�>�c�|�����{޵�~�������:>���V�R����kd���[����-�ġ�����@ifb��.Zn>�b٣%�1K1�ڱ��"U��@Bx{��)��(��@� u�X��� 7�	�'TS��1���:�t� �"��n��I?}ԣ1������p!���
�7��`���mE{��;0Uɥsy�8��v�qBcx{�SpC�勁$A!L�S+e2�L�S?;o�>��؟��%���g�ج�M�\�W@g��'@�t�S)��e2L�S+e2�L�S)�e2�FS>�|�S)��d�L�S)��e2�L�)��e2�L�S)�_}�e2�L���e2�L�)��e2�L�S)�e2�L��>~;��e2�&S)��e2�L�S$�e2�[)��e2��2�L�S)��e2�&S)��e2�L�S$�e2�L��=}U�\����e2�&S)��e2�L�S$�el�S)���L�{��l�S)���L�S)�e2�L�S)��e2L�S)������l�S)��2�L�S)��e2�-��e2�L�S)��|q��e2�L�S)��2�[)��e2�L�I��e2�׿}��e2�L�)���Gɹ2�L�V�2�L�S)��e2�z���.��;q�:x�e2�L�V��L�I��e2�L�S)��2�E52����}��L�S$�e2�L�S)��d�L�S)��e2�L�㌦S)��e2�L�I���L�S)��e2L�S)�ξ|�S)��d�L�S)��e2�[%��L�S)��e2������)��e2�L�S)�el�S)��e2�L�)�$�H&tp�b�1ZВ	 �
�-��e2�L�S)��2�L�S)��e2��2�L�S)��e2�&S)��e2�L�S$��L�S:���l�S)��2�L�S)���L�I��e2�L�S)��~����e2�L�S)�SKmL�S)��e2������Ǽe�L��e2�[;��}��L�S)���L�S)��e2�L�S)���L��	�yٓ1w�Ȓ	 �	 �2�L�S)��e2�L�S)��e2�L�z�|�S+e2�L�S)��e2�L�S)��e1"�!B ��QW�娫�2w��t������� 2�YuP��Z�sv�\�8���:�2�S)��e2�L�S)��e2�L�S)��e3߿}��e2�L��L�S)��e2�L�S)��e2�L�Q����)��e2�)��e2�L�S)��e2�[)��e2��e2�L�S)��e2�L�S)��e2�L�S)��g^���)��e2�L�S)��e2�L�S)���I�I�Lל�V�ʬ^EL�S+e2�L�S)��e2�L�S)��e2�L�{���L�S)��e2�L�S+e2�D�yo��#���{�V�0V$�c*v!"v ��h����{�Z&�{��$�y�{ G��b8�̠� �+:�b�dG�흊��؃�Ё�U�0�*ih�婭H$�I$�H ��n/3���1��t��O���C�rt��qU�ܴz�-��ېm�nl��0���N��Ѵ�e�,�#R!U�ֲ�hE�gR#;RXH.x��zww�<����Y`J�K�f��(������f�k>��'s��s
b y}v�{��.3�N�I��ʏ .u�Q�9`�k�L/w��{�Q�u`�(w���[�{����X�Q�{`��¸��P^���.'��V�ʬ���w{�Q���*���h6�d1d�J�#L��F�5�ڪ;6��ʃ_wN�$Z֭;;��{��S׮ڎ����Ud������z���_3�j>���@�ǱZܓUX�bTJ�l��b�">�/{@��v�1U��V���ȉ /{J=�l��V*L`�VTy1K�V�G���Z�7����6Ό��É��)B��c�IlA�DWmU
��dP�#���f�򻻬��Q�]y�� �;(����;U��r�ł����}���P�wh��ڕ=�H\�:��P����@x�a�P���lü|e��R��ֶ�(��0Ռ>|�m�Ee����!��jF �' p)	1�F�f:�X��^&D7x��@���c�������F Qj����f:��7��@�n^�bo��1���Pc�x�Ơq����ηޱ����$۳H4�l�AA�3�#q�ta5�]sDL1�����:k1�uÛ�Q�Qha͠x<�\�u7|m6Q�6��:�3�`5�h�dĤ:v�}�ÜU��K8$JR�:��8j��u�5�����y$  �2imKS[�i�yԱ��q��W���	P�۫rSQ65�Ke�#.`��er�8���-�Hh4��+��.
ͨ,�9�-Y`�
�5q��,�K�^����7�ٷ��~I�$�S��tW]G7[2T��E�ۍ�`@ٮ����{�0)E�g�9�>�.�3�k|�3j��@�u��a�cY�q�4=��� ;�B5��=�JJ:��8j�a�ƈ���(�D����έή��:�������G5ڕ�vwV�v����#I��$f!�o��1���#���Cwo�� �=� �yS��	�D���2��>������F Qhws�gWlWM��� �FL5�������\�>�sǽ�B�%EG[�[�������$�c&hg1���,�ڦy�I�)I*��xP�vk�C���o�f3سZ��Ut*�}=�����q��Ft�bg���c�1�n#���hfc���Yó�����tnEl�b+t����6ܜ�",H�
&*�fN�k1p�c����D Qh`5������kv �FsL�5�:�fA���b���C3o���|=:�1	e���bng@cy�l�x�4�uܷ��Y�����?~�~���[��4n�������b7rE��4,ֶ�ݺ��R���eWk������W�Gc�ơ��c���Y����7����$fd5��«���9�á�(���Ms�fc��c���w쟵�;�9�k������޾�: ��"���v�$|�b��m��8Ȏ*q��.\.9�����UƜ��_zpI�gy�����8\gf�e뭶��Ŷ��d�T�i $V�Ci��Bꨚ0Hq���,�����\ѝgK��8��Z�-�G�cY��s�bqYr]{IĽ���'�\�j�й׾��I}��{7a@  ?=��             ���s5�^�a։��� hl��3
�B@;T��K[q����9[[�mN�m�[g��qɝCg���Qdn�&�۠�G9�\%DX"���m��<�ڠûer��F�Ih�!�7]���&Jk| }1�k��4�m�:���
PZ63hT!E��p�vxL�Z�ۙ��36�mn�	ҒP��� d+T@93��W�(]�+� ���Ϯ-��B6��3,l
E�v%�Ӫ���^�X��P����V��r��b�pmⰧ1�v1��� ��t�FUt1V��l.�m+.�yh�d]�l7��oP\�Nv37%v�f�ޒڮ��=u:[���F���^camEI��we �i�dح�����j�\]�6段I�qz�қ�W-�C�-�0�k	I����R%���u7UV
j�+���Ӯ�Tm����_�p1)�J�yV y�m(H�V����#^+`��T���� h>W��C�W�(����Tf��&+ŀ :�N�����R6��h8�:�u����p��a�!È�!�qt��@��[�������D�%فD�uv��݉�O\��Zn&���v�e�����g��a�:��,��7t�K��V��챕�&6t�\������O}�,����@s�M��;�� G�Z2�h�f:��@�T�.ѐ�Ҏ��8�G�P�b�5�`^���3�4���6A���6������e����^����G����Z��h����]� �6��Ie�"�����uu��b���&N�1�h
��36_� #{�>�C���<�3ַ�!22"���5�:�fA� �p��#�54;�:����:Fg�9���a�n�����q��E#!��j��f!32Vo��Fb*9�d��uwo���;e����!��1��r��~�����{�c��*hz��{��f�n!:;b��s���uΝ��bR

'� �ʂ1d&$ƣp��(�,5�.�����a�;���@f/\�w�aK8��E������`�Z9��!�b2�
:��8@�C�tPU��g9yq}�����S�c3n�:Ƭ�",��M��yV���������OL�Q�>#�C�ۭ�ރ��lEFhs3'� ��o�y�"&�p���h]ۯkwg@��X�k|C3La9y����F3�۫�ud�|w۾��4���} � ]m�����[coG2�6[i68�e[���Q�g����v�-����n7������zܗr=l���%��bے�%FSe�$�K��q�w��}׽��g[V��X��tbح�$9!)6c�3$QX���Pr���{���6ے���T(��!�y׶w��(��ha �l]�s1־�V������
����:BD���Ywpa1�3�p���D�� ��
�0$�(�tf�)������:k���f:޷vpC-�#��Ub�
�w�{�u3�U ����Q�!7�7��{���5T4w��"�Vz���zŚ�uf N�����1���c�B��{Vy��mp@ۍ"m� ��nvz嚩k�)o���w�'�ԣ3s3%k�|��:�>��{�c�:4�����v_�? �T7��|�?�cZr!'__θC31�P��32V��6!����q�u��	��y�u�N��J`4�m��$CWhM��ݱ�Mf�Fd�-fd����	��Vc2�Q�ݺ��vƍ���2���5��wl|:(U��*����S�3"m��@����%k�����*�O{�J%$�!��<ݹ�j�ng��B&[��w�u���}�q��q:�fAMf!����7��-�5�!w��fc��fL��k1	����VjC�Xr"$��u����5m�.�
f�  s��o4i.Ӝ,�
\��Ӂ��ib`��̗�a�n�nN�;-�ll�j�b9��5�4C,�\<�����Q��'/6�c:�eb��5�=��l�I��e�ú�ƽ�����Cm�����9v����&B�SUf��.��ݺ���M���fc�����;���_m��w+ޖb��؉��N�Ws �t�b�c��^�:W��[a��2T*]=v�� �i�"0��u�Z�����67�0`�.LG��p�P#�� ���Y��SY�̑��ƈ�z��]���ِ��i���5��f:�m^!J!5Vkh]۫�cz
����%��X���a�A!a�7�����+L׼���^���U
�ׇ��DPC��y׮�V�A��D�q���\#�'/z��k]�����������{�����$���nKZH�R�r�Z�O���Z\ֶ�����4�>�_=e�ӄZqc�I��v��l�}u�{	]�-9.[��SC\ܹiɬ�.\�D"H�ԓ�ɭl�CYm+DP�0a�<���M��J�Q�(Q2D;�@9��>�����c�D2�uG���.���0��U�Z�v���ַb$d�?�5�1Ù�����x���i! -Q
�lT�X�Nn�ٕ�Ar fǽ�Y˱+Ƴ}Y��ch���fd�#�:�f�Û�&B��^�Xk[���3����\i���{�lklt��Ο�}�E�����޾|�ޑA�=���5v���5nHHA6������K�!0�uwn�j�x�c����0��vF���`fg� ����C\㬼u��f��.Df�VfA��[�5�A�]�!�����c  ��b�>��| @4.�
��U Gf��~���@ sg]l����U������=�P��d��I�\�����3(cO^��ػ��^�8�q����������d�ɮRӠ1�<�g��W+h�e6��lp�ִ�?zI�C���z���dP��H/���v���Gg�U��HRP9��oh{��wa�I׻�6P�5�!�m׽�W�R��pE*���]�]Y��8%�q�QJ���I��31ֵw��EŪ�[�1�����k�zⅳ+:�;jb^ؽ7Y�q�TQ� ��
#1��Eݺ�R]�1!r#4.��|�U�͋�:�qs�T�Mg����l|O��] {ˇ3f��	����8k�C1UQ������ei�C{ۯ{άҠ�V�0�A�!@��"����Zj�V�.Qk�/���Y�>�b0��wy+���fJ��:�1@�Z٭m~ �5ڪ8<1D�	� �#7�չ֬�fp���k1	����Vk��݉�2&���o���k"	���� �	V���s��
�-F�-F�3<5w��f?|��d)����Ad�W�u���ƛ+H����|¾��^5�'[<	Db(�{�`w�u�~ �^%�.{ð1FJ��놖cv��>��7��J�(�n�h�+A1#1�܈ģ'�Æ�8�f:� �s�$d�Y�Mm�ݺ�O�V$.Df�ݺ�z��]��m�*ڍ�ݺ��h}3%f�o��"��5�鋻uzߐ��ժH�%���<mӻ��;��y��鵽��F Fyr�c���m��p�wl&��xspW@�̳l�:^8���m��,�
"�'�o_�y̰���X`�5����;vݞ��FL�\���͕��+�v��=N��6~�t���mB�|�c@�u�m�)vi��QvD��λ�����������F�f��P(�2����/��8k1x22ab%*��p��v�Z�mDLP8�V|F��f1�3�s�$d�5����Wv�i�.�d(HC)@�AC1��4���W6��9�}e�;���r�VUI9�C��d1��������: �����ww�D��[����R�C��Z��u}�,~}�I���� �!��׽�%�Kf��%�C3a�(
����*��d�Z(y8�JD���ᆚ����X���$��4.�R�1�f!wn���؆)N-U��@
#|(fc��y� .>uA!��+4s��w�Ow�"=T's�Y��&���4=TP��+�n��b��m(����UB���35	7�MWj_�{b��:�c]H�RU��YU���;��J���RZ�| �D���9�!&��$�~˸�ei��B��*��U!�!'ﾐ�|Q$����qs35�M��<�M�!NI/X2EE;�O@(fkZ2NJ�Nʓ�*�X"�Vz�zĒg��E��p�O��K��s2Bv�3�_��a���2����L�*�#@Ѯ���kq�x��No�։9�:(UUi%�N���3$&s�'��P��s$$��d��
V֖q��"m��I��!$��`U >(���bEm��d)E�� ( ��$�I��	�T��BI��fD�%-�>>h�sr}�HI8Q%՞f�O��/���y����<��7燚2�T$@�v�XؔT��r@'b��1�<i�P�m�����Ѭ�s��9�9���9ɪ&I&�i�Z�y�r���g����pԲ�k���C{Հ{�ѽ��w�����}  l Hh            ��u�]z��f�eȬ�aLp�n�{.�q�
P���(e)r�-.-�!��b%���&n��d	w �6���\�c&h�1�hxۋ��	��(*���ӬY�0)c
�R���^�����gI%���X;Ycc�ƙ6�t�{
3�7K����$`nx�;�h�*���x�e� ��Rٗj�T6g]�6j�T2ܱŔL^��,T��#N;	�dث��F�ob
c��w0Fi��FR`�����/�]�5�h�B�\�j����<��Mcv�����BK6*¹1�ƍ%�l�A���	���H=��9���g�|�cO0������-���+;������@L�9mu�bm�I�n��*WGE��.�-��9�ki���XX8��p��KZ��r��I�6��d��0	 ��C�Z�F-r�˵�,,�՟A�V� mu���S��q��&�.2���������h_�$]hT%+�]	◼�B�%/�KB�)~�N��X��"*P��>(�AQ-Dr��
?�����u@{��l�O>��wy���p  5�gl�Ae����m�EԊ"HP�vd�gnbv�F���VW�%]��&z	c1�G!��ú�L�cd��:񶹃q�7-�i)����}�T�gn0Qs[v>��ē�H�+n��2�f��U��Tъ��ӻ�>>R�F� ���P;��	'P �8Q&f�p��o�D�d��gMp�NfI��	��p��q=N�'es2BK��h��c�Ј�H�D� XY'[䄜̐� ��Z����Fd�âNfHI�{!$���P?/���o�&�ص���8�sfi�X̿���Ϩ��U~-�̐�vQ$�D�̜�'3�O����=cRI�^�	�q�J�I�RO^��}�wZ$��c�ȓeiql�O7Ǻ>��w:��P8����>��/��F��>4�p8]�2�`�u�C��l�̉���v�����������B(L���fg� 7��y�	���d�W�Mm��uv��g41r񊘏{�3���+�[��
���U�����mMw�+��fk ���QD�Q�ӷ\<#3���������,m/�vͦt2�H7=�@L������MD�%i�5�l1�y�ګ3Gh�F��o���Y�
@٘�D����]�5wn�{j!'Wj�s�|Њ5�B	�_ola����b`Őf����ػ��!v��
��ޔ��$j�%��b���<݃����}A-kB2�F~��]{ʰӠ7�&H��=�~��� �^*�5�y�~ێ�Q%uv�dxP�@/g�>��{��5+Ku��lfc�T�Xu��J�Dk3�a�_��
׊�W�x  2uݧd���6�m�V�!!fP�%C[PI�h�Q�H[�M�bٗ�`��;Au�E���8G3� ���ŉ��1ўRX��=1�,��M�e�Ճ�R�'���;�������\e3Ak�[]-HF\��8�UI=��L��{�uΡg��P{�u��#P��{�ª���c3��&����3c�k|wF�Vb��e�YUTf1�c��da��7��be)����� ��a��c4d��B �h�g�B1��%Gd�U��i�Vb�G��3¨��y׻���Q���_�s�UT4c
��A�:ĝl�%����u��XxF�`|b����%]��]�x��#P8�qV�fcv�[�\��bTn"ډ		��"X�J���]X�,�}߅Mm����Cb���ˑk3 1{��B5�^=�@U�G�FCJh{�~��߀�: �@��1� ��(��H<}�P�f��P��J�;��F���|kz����T���ܤ�1��QE܍�kj�vڬb��̵��~~~i��:��5�,=�1h]���C��^��L�#P8�f*�����u��r�EA�Ykl]����@�sX�P9��-�� >�˽W���p�h�Ѷ�ap��a���
�jǴ4Jr��431�Ua�31��W�(��:�U��.�v�Fs�������x����#ﾕ��8t��DGf1;���C�B��5s����C3w�f���A������F  K�7;D�ln�%�8�7�\ ���#c�!'��v�݊3�'q5�k��X��ڣ���.��I��3p�X����8����&)Uk�������bjw�I��_M|)-��F���nq5e�i�\-�ԏJ!��9��5~ޡ9�낸o�eA�?
 ���u��GZ� P9��1�����#>����4.��:�7� <4��=ZW�E��b�����ݺ��g���I�@��n�VJ]���˘73~�'�����j"�|�yV��'���lB/o�&F��~��@�d}�]w��ג�&��}z/c���3%]��U@�5����(�P8�f!���1�P� ��[�u`2	��5�
���|�����<��kd/p�P��bq<P��k���v���B���Q����1�s��Y�s�Lf6�л���U�
��s3pg�1D�Q�mV�㪪�	����[��9�s���{�����uPy�-uW��qR�PJ)�E5j���e*2B��(���e�M2�W:�Vg)���V�'-Ħ��[��(����Ӿ��tU'6s�s9����E���Ȣ�H�[Y��������D�RL5R�i���M-�֟��>`�S�K),<���ĥ�B2���=���%'�w��>|Х)u��e$��aY/IlI��� ?U0Ep>�O��
��E ��'�3�g�s����Ӝ/R�Z>H)>r�g��ǵ�6s���I��5���h�UB����Kʼi�������
"m������ZI�`^nzH����UY�B�31��"���L�E+3��jݱwo*�Pn�{�B�3C`�3n�����#Tf1������6P�t'�o5�F3m��G:��]�i�A0�-( )��,�w<�Uv�*�e�;�wW_xkm�M=J�U�H��.���|��8�+Ku��*�O7�=�:�A��{	0�5wls|�@��9��ޗ��]b�w���)�:�Q��!��(�����?P �^������~�42���`��I$�I$h��`2:M��w��A\fҔ�n�-�]�a��Chɦ˫=m���nX7,u�u�m�C��i��*�ۅo\�2�݃^��z)�#n�-qIi���k���yu&C3�t�7[�2� �,�;��@ 5�	�!N�ʳ�Z���
f!�g QĤ$�fd�<�u��¨
�@㥼�1��P�_��	��G�e���Q%c¨
>���;��^���\i����^��{����1�,T[�k��1�t��&�l� �I�Dz	0�5��w��
Vb��|1ޗ��]b�O9����[���W�#��'��2��[#(@��A����[�d*4,5���c.�P��k9�D�$���c��ܮ�4�������	�:��+;��]�
T�B$
8�f9oB��s��� ��Y��Q%��\5��.��U����q���;�޷���W~
�yF���a�GhQ����:]f!�����S\=���Z�ڬ�bi�0�F�m&�G]�"3۶���@F��2Ԭ�[5����rV�}�2�6pP ��g1�b�w�r#I�G���9α� i{�a&�kX�f6�֏��5]�������\^�ڳ�֚��(�FG_|���������;0��=F샵X�F��]����Z.0t�^5�m�O�}?Q��o�$�q6}�H7κ����D�	����\�5�ۮ����5*�V�]������#!P��S[b��]��]�*���;��_w�   �.ݼ�.�.�밨v�Լչ��7\tS��T.�h{cvF˰��åm3��T�hU�^��w�cEvb�t��n���Gvx尩�5��#�Z�Yp�X{SϬ�.e
M�����ny���4�RI��f�뎲�4ﻴc1��оۧκ�Wv�sef�))&�J�G��y�{γ{���4�Qn�kz������ě-Fk3���1U�O�շF)�U+Y��R��0X-L��%@�p��ݺ�UY��u;�1$%��f/�i���ǽ�Z������55�.��5����b�P^1�{r��^4����ciM�{#�Uf�ޟ>�O��~o�n��sb=���tl]Z\e+�������}��fc���w�Ɗ�[�>(�|xw��Y��wW���x����:ݞỰ� �� +��U�X9��q��=�u�n����t�� �F���?z����y��������b�I�e�:�@F�^u&�ؑ�ۑ�L��]��8ĻyB��oYȌq&!��c{� Ø��  ��s��ciM{ί�ء@�31�^˼%DJ2:�\#��1���W*����h�]���)��5�o�{<뙌o�O�^7<�ݻ8�����r ��%D$�&ˈ�f=��:�ʡA��h�<H���̂�Xk3*� ���H$�Y�vBk3��o|�c1�f�� k|~>��� �������Uʬ@�{fu�y�;��~���p��3���I�_�߻����G{����{�jM�I HK%UI%@�'�.�4�0'��4-m-�6�λі�C*D����Pb^�*N��ä���4�i4:'9�g��̸�#��-d9�q�-��g1b��,L-%��0�K� ĢSP,�汼�6UP�wD��e�:D���E���߀ � �            ��۸�1��Y8��Úٟg��Q��
RzK����j�r�*��n�ηm`
��iU�-[�����*��M�Y��YgCu]�N��2	�.Z�g�Cn�e-�t��P�U�^" F��]�v�:���(tL�q��He�CQ�W<�UT�A���-T��݅� �O\��ͪ�.�L5:
Ly�HAB�����Ve�J4˒.֗Y�
dV@Z9W�sĎ+�s��mY��q�Un�aM�]#��dU�6�%�`�6�I�D��&��5n�g+-+���M������h�'KF��w+�r��:@76�Pbp��@�f7ZgV�L�^��c4n��u�"�o)nr���F��c`"�5��T���W�`��\�v�ȍ�S�l�`��$�[�qY���lU:A�Uy����N*7Mմj��5X�zkl��h�5
ت壬�J���m���9\]
�a�3�,���tb��i�/��,@<�@x
"+��[)M�i��Og���߱  >~7��{>;u����G;��t�9��e�v1�V��d3	q�����5tlN­�qnѰA���u�sϮ�N��И��<��!2�G$%�`cY}Pz[����~��$��|�.��M����Uֱ!����D�Q7F3Q������
� ( ���7�<[pю��[5wl]�� ������H�n�Y�����!�>"�qa��7�1�v�P�8j�G��9Z��Uf�v�啴�NӅ#)���2ݦ�fq���SF1%F�f!���cv�o}�c*f���8����36�y��y�$�5��7�:�Uf�ޭ�l%4.��;�����cCX�ZSR�p���f:������I�h�Bi����M�e�J9���[�V�F�s|c����D��a(�]��Q�z�Ҟ���މ��VNrr�<�p��*�i(�		!���Ts��o=�c0(�]�٫�~��@}^��\�s��ThY�o�fc��,
�!��
4�����3�is��G6�����WD���1�o�l�z����<ֹ��1��SC~wTGmV���u���+Q�V`U����y�{ν����P������31��v��������m�}��7�Wj��������4j»�.�B��	4�0Im��1���f0;ݺÀ��8k7x$��[,��cfO�iw��DT{tMMm���{ҽ�$ץ�PF����]���� �-b1��V/'{�}�彏{�=�>A�UO����^��E  ��Ԑ�v��ݭ`]���-��{r�A��3��ټ��:
���6�u��{�}�z�W=�maK��7 ���;n�W��"s
��n8]�+�8��MmN��=�n�xqG.N�1����m�:�1Q���r�9N����V�}��P�9��9���+K9^5��{γȆm������s|c���*�]Ɂ���C��*�V�9�X���(�f*٫�wlp�d]��
L�p�J6�2��K .�F��wß|����f!�o 1�P�f?�w��a���F3Jk�3��U!����5�xZp$�u��\�1�fd�����(in�l��y�=�>��9�)�(����A����h�Ί��°b5�����ҫ5˖�1��33$�{u���n�F$
)]�[ ���2���
 vjz��H�/��	@��ؠp���f1g�����d�ن�1��P�����<j���	�bi$`�]mR��X2���'N�R=(��������VG�fc��'��
MGY�x*��f?
]C��x%	+An�5���߾�W1Fi�����h �z�g<徽Q�܁$b� ���H�7���E���xݪ���,V�Ǒ���{]������B�vۆ(�
 AВP�[5��ffJ���R��V�\��뙏��T���M�k~��{ʬҾ��MFҚv�UdePfH5���)5f*�U���g]}^���v����$�I$�fq�N�������v����rm�^�Ӛ�uƉ�A(�\A��v�֓`���S�cQ������[g��r���ȣƶ�A���d�
�\΢v45�gs'�O�@�K���5�4FF�NE?���Ei�����A��h ��Fm����f1���f:�]�`o�Ƣ���]�ʡ@�b��`f��H`1J�U�Ȼ�.���n��dI@f��V
�7�����CXu���#!�%$��M�r��]pzy�1�DfI�F�ݱ�u��p�4���Q���ݿ�uC�=*`�s��R3�^���1*���1���~���͟����%ilz���\���f Ƚ=��1��9�:��w�����і���Ů!v���DSRC8*�7����Ɩ�f:�x�[��v$f��v�5wn�v�5yj�I@f�M�e듒I��;���y�O<��<�~4B2����H�22n>G�b uX�lJu��t�Qt����\ˁ�4B�	V�B��wz�* ҄�(5�K��YhN��sNk�PB��Ii�� ��<F%�%դ��%X��8&OF�6(TCG��� ��A��.�ިNkq��LC]�����Fg2�k3|Q5Q�fc�uU�8��*��|�Lm�X��el&��˘6�4m�Z���u�*ޕff
�=Z�{��>aFJ��|F�k�N��f��L�]��vsa�����E��P�^>v�|�������V���j���QZ~M����Ӽ�ϯ��uv�R����f0�2VƬ�`P�����Dn��RMo��e�J3Ud	���uz���#2D�CY�Ʒ�Y�U�A�]�Q���ݰ�:��j�؜]�Ђ#��B3�3�����aFJ��|��P�p}�]{�{�B}I!ӻ�wI��}��UUUUUUtav"2Ļl���@��m�D��K��@7���9��2�
kY�F����2�p�-�ol������F�d���ѕ%�xg���e���iܖӹ�{�BS�p�E�&`��ciA0�FS�I"�GL ������B�5��/l��Z��c��&񁙌�tD�)Y�c���33%s9�rD�3C����X����BLڌ�p��bo��F%Xk�=��B Ѩ��T��m�ǲ4IQ�����[�uU��۩k�Z�"�uv��ECYT س�'�ǯ��_���+Ku�[���+K�����)�Q��9�:�Uf�m��dQh]ۮ�U��w �J�oʲڴ�lR���k0���3�W-V�]�P����s=k�0f�Ϗ�
(��{�u�5�[��b�vƷ���ڠ(��||i�7�q$���y��	*��cí�xZ�"�u��;5��]���
;��a��|�F���u�؆��A~sAFJ��x���>��f ���"�&��s|uv��}��ɑE�wn�՜XxQ�{ j�(`��>>�4=�;��᪔B�:T��r�3�ԅ2R�@ַ�.�Դ!^ˈE	U)N:x��λ!�&�p�wlk|uv����0�()�wn��,�wA��w��"-GZ�6kꪠ}�?{ν���oM6�> o[h�c����S�/����*��`~����˼�~` ]۪c�����v��PVu�kv�d���R��骔�i4�siB�j��D�3h[�i�:0���{��On9��C�^hy�:�M�MJ�Ҫ׭��nU,�i�������N�W�N%��W(W�鎎�KQ24�.2cQX��λ�> ]�ww�ʉ�����dxNc�j�uHShYklffJ�Bf��$�5��k|b�0᧚��%43�UY��b����?%��앶�����.�&HL�%!j�Q�ڭ��3���{���i�-׋�1���{n��df�L��fc�]f*�0�^�J-hfc�uVݰ5{�0�]�٫�b��^�m����uiڸv�AeL�h�eJf5K�}߇>�������/{��b.�o��hYҹ�0U⪫��{g�r�L�uB7�ԚcX���b���^5B�9��f����oO���o�{�u�����U٥�b˝ۚM��Xb$b���E0L�e�o��в헶Lj-�uޡd��f���b������ݺ֮�T�8KkB���v��~�� 
~���fH����y�o����>"t�1"d)��e�v�Cp]�z�V�a%�s�t!��T����!I7%]�٫�b��^�s.&�kOu��k|c�����S#Ww�;κ���F��Oh��Z��Uda��.�v�_����9���y~y����6|`IB0:��"ڍ�wa��L戀e H�@D{�T�ʲy�0�*�/P�Ŷ�Y���`�O����   -���           jM�������=�i�6�5�ڗ�%�z�#Ř
6�*�6uZp��B�۩��[�;$,/n*Ѷ^v��\.�+�3����l,���py���1��n{8I��{8�U����ǭ���T��A�ك!ˋ�:P�Nh�ب�a�M1a��bŊ�B�v
$65e{if�9Q��hRaDX�<v�����R�*���>P/H@�kj���)v�Y�Q�ukV)<�f�s��T�\�Et\l��2�m(�g�wTnS`n�c8�-��Fq@ZCc=���U:��˕��Z2��`vٱ�#��[s:�!Ş�� P��=���ͺ�6y.P���IvDۡ�� ��$�C	����MRݴv�-�RC�}_BZ�`�κ�ij�9y��\�6v��m�KG)W�@UHHqR�-��ԸsD���U�Qn����3V���E`���U`v��u����ɰ15c]��hY�%'t����N�Ћނ� �A"	��"о p4(���z������k�0 Y5ҭ��؛k�!�X��GV9�wL���n�B��ӉrD<�#"�0�-�+^�b���6;6��;��V��޹�ъ�kg���R��뀶"����*]=:J��vK��V�,S���[����B\�q�r!��O�l�=l}���s��jB�����ػ�Wk���!jH����5�1�  qf-���xb.4�׏���j���%��jB�**�C�<�k����]V�A���h�QD��MBLfBh�)&I�3���j�Z]�G�[���߰�kX�V]b������4��զ��A�� �xc�7�f:�P�v��ݙ!����8@��fJ֮�T�1Ւ@��v��+Vv��36^��,�����3��HԆ�@]��D]�daf�Eƒ�x�Cv��w��
	�Ǝb5�ؠ�@a�~w�쀃�����+K�����f Ƚ�"�&}����Wa#��̎3!aFY�	.�v�AN �1�je�6��K-�uΡ��`^�̐�b�v��PAy�=�1�yֵ�t�"�� M틻uv����!��^��f1����y��T(�;���{[�آ24���ۮu5㙒�9���H�a@cp�!��-�Ճl]_+�B��������'�g��fc����ai=���T!9���|�A���q�$�2��|{# B��c��n-�h���Y]��E�jCJ��8@Wl]ۯ�pP�@w�  [�t��Y��pc�Il�쒛y1��/5P\Y��켶�(��pk���t�͔�� n�iܛ�\�3s�M�v�<�F��r����.H�d�Q�8v.��S~Ν	$�Ƚ8]��/0�dGRM��&ጃ QNl�{c3X�������]��q�Fe��	T%�<����'\��@WlC}���&���n`6@s��Y�����I�aolfc����;m!��e�	@���	{��r᪬�0mw||�Os|uw�,�nX{�ƌл��n�����~c�f��0�k-��v�]���E�d��wlX&��wm��#N5vƷ�J��!�{{m��A�PT��4H���Y����fd�ݱ�F�c7|
8�b&����M�.�^��\1��[@[�_���PR� ��5���՘�w�TL �cw���lL@d��a����]�X��,^�v�q"�.$���]�����.e��̽3����]� .�v�o2ʀ�Z�4��31��Xح�|q�����]��hy����m��u���5���@z��T���4u�I5�lp��ػ�*�Vy�6�L n$�p�BZ[e��粳9��=�3mC�}O���}�������2�"ى 9�z<\u��֏���)��3C2�w�vpc��,������c�����Z��Ld�Z@Z�.�]��~�_wn��gu��|K�   v�u��KpT)Vb�K{-�Q�r���=N3>3�Oj��9Yj�J��������l���%���X�6AI\��� �&���&����@A:� �vpp�]���{��ӧ�$����3�c��j����ڟ�N����>���;�1����w@�M㈸�e�p�^J��`��=�
C����;��c3f�s����������>2����[��������a�0��d�%],��k�Ͷ}���f��0�AHI������b��uz=�LL�]����� LB���1��J��fC2��[cٙ9���)N�g�]� >�V�.&��v��@�n�uvQ, �RXf@Ɓ�@�u[w
�_�\�Z��GY��z�y�fc���wі��{@Z�c3]��E��0v���Ɩ���Z��;��Z�����<�w���#�,@�[[U�r�n'/������!9�i���;��͝�%��7�p�4['5�� �m̄�`�F�eD"�J��X#
YD�*�}4�3�2e�<�q�DpA�Ҵ	����H���i�m��f�͵���SIcjz��-�#�7�58е�Lj-p�B���j���<@~�W�y	����c�v�ݼ#[#2�b@�l��6���+�;m�E��`b@��������Fe���c�F�����n�-���_9�"�)M�sޕ۷^4�ޕ݃Mc�]�G;�=J�V
�#Y�{�~��*��u�K[c3]��l
���#q�!$��L��<����Y8��&#[�,s|u��Vj�=�c*=�a���՚wz�T����J9[�`�d�c�-��b2d
-V[���f1���7��qH�0ֳ�����u��UGw������"�  �rb��$݃]�F.׎�$�v�k.�9�t��n��٣�[��ݮ��$[�L�Z�\���pLs������r���D�s��sve8)�̵ƆF)tc��ߒwtq�yt��<f3v�ՙہ�1��F㈸�nl{�u������ի�2D�Q�ݿ�O1��u����i4΋���3��γ:�"�ȋd�@����w��1���=�cJ=�u�u� +�!7v�&[NBl9�HR��l)�b�c�׿??7���j��\���Ld�KB��� 
U\�5@V����u��4/����v��8�ڻ� ;֭�\eG��:�ۇx�y�b΃!�����c�v�ݿ�(w��E��(���P�1���1F#q��Mj4�zO��ol~����2����[ ������0V������^�����O�V� �} ׈	���o| ���zݑ�M�v�j�2d
-4��ݱ�2���"c���Z��v9X8z0���f$fHY�f1�q��X���-D\eG�wo=���h��5��$-%f[ +�.����e��OA=� -����`�Q� �1ZҀc�՚�9q�JV���q��X���m�d,)�Mȫ�p�{��V@"��q3B�߈��0�B�u��P�Ù܂�#��j�2`�E�d���w�2Y�cCyȌ����a~;�]f[@y�ِ�ʏB��s�udv�y�w̟^��0 KYs\X�!����ӣk�]��F�P�W��mnwc�֮�ۖvwc���-��zR4�G��;I��Y398��6-���J<�i�d��~i�T��-��!�wwԝ�Ot�;O{���{D��a��[�SF�13�ك��/@Y���u{��q���{@[����B/���	�j�o���Ś��`��&4f�f4G{�A��77+\�P��]�� c��+�y��p$����"�Dֹ�7�l�/S�'j���ǳ2Ve���"���Hֳ�<m�Ǜc3��g6dD�w<F��^?
�#C_/p�\M8�=�:�n�x��bb�	J<#3t��c3^�s�l='��K{,a�Uw��?[}��2�%.��������H�
H�`�kw�s|u����[���L�wo��XifjV��"����r�� �B@*�S� hQU�.��^�2d
-U�Z�vœ}{;WȢ24ۆ�v�w���n��f�m=8=qnX�����ƐƢ�I!��ʁ��c������%��`�����u�J틻�^�r2�zE쑀���fc��X�_9L@�{g�yo{��p3`���2����E����ޱ�<�;el�n%BB����\���
,]�#)Y�놱�x 4=�:�s��2��*��c3fu�ys����6a=���z���="-ڌ��SB��s�uf����0H�m<#3�R�S�{�u�p�?�*JߟR�����r����~_��@��(DT�s_���֮�N���9��"�b"H
 Ȋ��((
��UdQ	lٹa���Vښ��#)+�Μ�מ9���"�%��UK5}��T��}s�Dڭmjuy��4I*��+&�lYf�[0�&1�L��ח63uMfV��͛VM
���VH� �-] ��E� Q��ͤ�mM�TR���k-�739`ֳj+K6�#a��nC�ł�Y�PE��qj��
p��`���-Q��o�ly��**��( H=����O���g�� �|=Z)����
�Lz��
%���ZDu��� "'��?iA�L3���L���^l�c��gч����(������=��D����܊� "���j�2����~����	�O����>7��{����?a�HF+�bO�
� s�������i
�4���������?tt���Q����9�ݸ�AD���\	&�������]zc�I&4"*R��DT� �Y�lh����jfᴁ�3m,)�e1�3Lf�3jm���AM���Z��R��ն51�3�lr�e`���Z�����l�1[m��������m[��6�3��m[j�,V
�)m(ځL�3V̭���c2��m,Q�+�&K2��B[���
aFژ�XfVm��j2��)��B��Rڔe���$��H)����LצS�<��?���������(�顐�
%�?����g����a�v�6��a����ڤ�������`�U�JO��_��r���~�z������ӕ~ϣ�!�����a?�'؟�ק�����
� w�Q! |�����O�}g�~��jq���}������ ��������A�*�>M�����,�-O�>� �>H���?��@
HB�?U�oS�A&`f��
":4.��-��cv��0�a�@� (�?�Ҿ������>`����=�E?��?���������?)�5S�����t��� ?AI�����<p
� ~"�����>�U�a�����y����~�����4Փ,p~��F.;�1>�1���9���8��ӗ#`� >��8}�U(����
�_�w���x�ADJ'��р��� �����H�D ���m����@O��y����T@���V��uq�j���p�}�?���� q������"�(Ha1jـ