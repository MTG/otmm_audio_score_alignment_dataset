BZh91AY&SY���H��_�px���� ����ay�     7�� 	� 	P*B�)  6j �]�
*��T�P
�P(��@��AUT
T*! � Q��@ Q@%���Q (  �A�P(  UP T% )G     ���hh  J@ |�S3�˖\�q���p ��	y� 4���x �� =�Һi� N�T�t:ks5Aӟa�)��B� �+�N����U�t ����   {� 
   @r :�S��ޥ�U�J�ru+������Y�J�j��k�s��=� 3�Y�ԫ�__ n�*ŕ^ t�d��ɮZrʩ�T�� n�2�*ū�]�����t�x� |�P
  B�F �K�˾��m:ӓU���,��._-sj�d�Z���N\��� �w�_q��Ҽ�\ �W3G[�^ڻ� �U�}��m*�5]n-J��@;�S&�Z�9��T��ʪ� �  (�� �ڥ;��My��Ҫ�5]���*Y�RŽ[���秕ͥS  �T�wەy���76�VmJ�����Ҭ[�\��W}n�_;y���� h�R�S&�j�J�yr��z �   ��
b ޅb�i\ں�si]��w ��ҹ���^m>-94u�M*����J��]^�N�  ��Թ�>�J� ����vK�]eɥ��ҹ���S-�S�W����ruK�            ?Rb��R�H�      �4��$�bh2i��@ 14 E?����� �Ɉ0�i�d���U)#I��� &     D�	&ʒ�Q�      � JPSD�L�@&hdڌڟ�?����������������}{���� 
�����
��PT��
���@\��U�ە`�����S�s�U�����*� Qu 	�	B"��!D��!�$?�U�E@�T�P@��>��_�~�A~��AW�>�P�G�QS�T� ~�Q>�G�O�A>��`�PS >�_�@>� �ES�O�~�P�DC�P�G�C�����'Ы����(}=��D�_�~�PHB��	H?w��J��{ r>��� �S��>��_�{���$���/��!��*~�?J�_��>�?B4�~��~��~��z��C���NK��"@�"}#��C�_��G��_�P<�9
n�(@�_�>��D>�9 }(u}*� @�'p�J}+�����JH�B�����!��H}/�һ��D��O�����Z��O��Ч� ���)���S�*��$҃�!���?J� @{#���҇Ї��Ы�	�}?@"� }���>��G�C�S�_��O �i_�O�~�>�>�>�_��S�C��ZC�C�O�>�>�>�C���>�<�>��CP?B�B}�_�>����>��O�~�>�>��_�S���G�~��U>��;�~���G�S�!��}!���r��O����	��ԟB}*}�+�Ҫ�
#�
	�!��/�('Ђ�J����9u��hf���]�5�,������d�����>���t��O�}��_|���N�T�$W}̾:|������wwvJR�Ɩ�)J�8�Ӫt��e;Q[WP�w.�V�RT�[�QvufD��T�>;nfE���Z�7�%��%	o�02L!(JY�j�`)��1�(JY�;`�M�5� �p2d�I�Ydh�!7�8HfBj(����5:7c���E�}�~�d90E�c����p5�jqrLk-�gg�����F�;/9�1���c!�kX8Fo]i����׆���I�����(JP�˧v!���a�N�;5fF��x�睚���Г�6����A�F�g4jpևPD{a1��.�2p��8c��]l��3h6mٜ�ё&�;��g�Ӥԇ(cElk	��%)I���A���	̼������/,b�E��iD踜�btZ�R�������������d���=N����ʞ��#��Fʜ]�kDZ��MA�Y8Apɷc5��1�����ky�LNc���n�a��s����ݗ.7n��/rm.M��w���ڭ%*I�h�Q�zs�\�uî��up��&d�w��gx�d`8�&�`E�\��;���2t�y�q�r����8l* ^�L$�u��we�ǆ�浬�=���(tk{�"1�8�JL�R�ba���,δnM@et�=Hf�c��tw&��21�X�����l�obQ�v�99�cNP�Q�� �[�&5'~�g|�V%�^F���h,�8�� ����,g�}�;��xC�z�g��!S�)��j�Az=x'�r.�ڧN�J��\��Ws��Y��!]�K��"��
��]tl�7���z@�S��3�u���x�{h�#]���dD���嫫n��Ș��� �	Bu	Bs0J�&���5r
�t�w��dq�XD��i�Ga۫�w�F���0:NC��w��`�7=�ad;��z�q9�a�ph�Q"*�W��ƦZ�f�>��9����9���1܆d��e���͡	��Ȕ�]��y1�oI��q�>b:_�,�U�MR���E�v�'ftoÛ'�z�h5D�d�!�'���p�����xNç�J��BP�%	Bs049/0v.�}��w�w��v��Y�m�T�vKU��7T��a��bd��3\둔Œp<�h�<�9���k�sp�cS�`]Bw	�'R&Bw���՚n�����J�$OΘ�jZ������|��������+�'xʰ�1��F�(L��)�<��:�wN1!�8����X�'Tl�um��"�Ћ<�
�y!9��X�բ'o���Lc!(b��׺�9	���'Qóy��\4[���T2��-wޑ�:7,���Vc;��3+�]D0�����]Z�ѓ��L���wK�N/ 6nC���잨<k�n��3�Q�N��!)�����"���sQ`f�K1c �Y&�!(1��z����d�#��˜#}�0�q�5��7�#�0�A�JO�\ΰ�k,p��hb�m���h�f�5�yb	XD�kF�܄�4�9ٚ�^o���EbA�r&����CE:,0�N�C9�hN�3Iy�k�uޤ��OԸ��;�a��i�6�DF�Xh����o�����`ua����z�2\r1�kk�F����OF7�dh.Z�`f����O��7��/Ᵹ'o�ި��2����	٨"V�b�y��b�"�yǆ�8��bh�.U�H%>�	@J��\�d`����Dp�Y�;�{]�_���i�;xf+8F:��f�|-k|�h�F���N0gDRwf݆�\�����^������S��5G(;�<Ԙ���x'!%�qtÖ�NN��5�.BPf�����npĝ@�BPOdR�٫F���³BP����R�I��\$O�fή���@��7;u��Y��P��Y�z6����$�d��h8��4�&8Xhհހ4�٪N��K�켌7�r0�u��uӉ�5�������%�<5�k,���wꄶp�2����'^Ys�S���]y�!	%	D�U<�1S�N�.�c�����uެ�|��Z�44�3�O"d�:ۋ�'P�'P���T�a����;z<��c�3#�r��FN.N0{9<}�]��nN��;� �%�㙓��p��tu��f�]�BRK��\0���l�J5p7�<s^�e�/<��^g:`��q�"��S��$P��P���LYrBP��Q��d%P`PQ9��k���hᢽmh0sI�=2p�"BJd^�`��#C���n	A�r��4�M���N#0J��A��uY�6�fPf:ޫ9���xuΌ|R:�d���<������d�e�Y�`i�(���Y�P�;��:�5��BZ��`6�Qh!Mhs�Û�D�����e�A�0�޳G(9�!+I�N�:��Ԧ"�X[w��Y�[/-	�10��E��o��.yg)E|ã���O��Vv�uCw'�����c��k��j�#QBpm�.9	Ocޠ8Q��i˲��k�v�ǫ��s��u��	X:u&�棼y���5��6t���6A%�f�����p��\����xGCC9����u���냑ݮ$��2qw	@p��i�&2M�K�Z4tm�b�F����.��	��!�!�˪lyU1�}<c��N��#8v�pc;�5dm�j�Ώ'�xgn��fs��u�u�������o��y��z� ݭ�Z���8Ƥ1�gH'wnx�i���K!����N��F��B^�s�lѾBqNy���_S��gr{�V4�dM{5!�vÖ!�d'��	(��I;rq�# ��}�y�ф�׶���qٳכ����:7ͧ,4�S��֝�eB�Vg�C^���f�i�u&:M�������r�r�DYkQqt� 8!�;�C��yscW�����o=mOf�XU�cY�Z�ɚ�[���4:�d�q���5�(Jt;��EҎ�/2���~�-�MSM���?5T�˜T�'Q�}��挲ʝ�U�������0(�p����Z1+��s��q����*�g�cY�F��c�Z�F�1��������T	Hk'� �B�}�v�ۤ�j��������w�!8���&,/����fI����9�.��=��ۧn�=�4C��G]������e%�]����ݒ��
��X�9�BV,a�6�hؕ�lw,��V^,8��j.R��B�BW-�ۨp:��d�%�0J׺�I����&{���Z���L�q�پ�Ѱ�M���j�j8��J� 0�JLc0N����^���Ĝ�d&I��&<�+|L1�;�հ�Ņ㶲0��ƍ��\�4w&1��e��;�:<MKө12ˎ@3P2�<���P���N$���k�����u�y=�6�p������%z�ç�<�`�(	�@@wb.�g�����&ԛk�0�l5������5[����q�͜Nb�MA��f�.BP��d��	BR���ō�!�p���#r�wb�ղtF2j�z:疅p�u���m%g{�!�5���+*%�����htD`Pt�Qxl�jq뛼�d��]Ov�8�w�{��]�M�R��瞤��2p1,߱��G�{��:��5gF��7���P��t���Ԙ����Hw�	NY	p�4fEW���t߮�O����Y�$㮞�sG���du���v�VE�Y�F"�5+���PF�:c6n�D���&u.���u�������N����]9t�4��N���O���\󣬟��p�P����.X�a�է�K��7Bs0Mð��t�sN�خj3�6�e���Y������E�==�O�ݳ���,�d'���u�錃E99��'�`�=]����,��A9i�ַ·��뉚Tꚢ�j�f���E�nb�w�?�:�N��ݝl�C2LN�0�qqɌ���w��y�]L�FۭEn�:�pJ1�'TA�k��s��ر4�����4�Ӫ����5']��!5�.�5	��fpu&Hg���P���'P؇�����d�0�����-�!(��F�!���`h4w!��{!�z��g!���DU	�p���(N��l5cg�u����`�t1��JэQ�1e4�da�u��oy�3�ը��D�aw�w٣w�۪��8;\�����̓,�n��Q��߸'V
�>;�R��X_ts^�A������BV&���I��$��%��F[0����h�Z�9f���{%��Q���oQ��(�<�Fff����%��l9Dd�rU�^�ms=��0�3;`ja�$g��$��Ԙ�fNUdL�r	��YFp�g`u�Ç^����)�8�ă 1a�8���'��+8�îu�2W�J:�.���N�b�靻����:�Nu�;_��l~=N�;����7Hv��<w�}���d|��I���7}�.;*�����5�s���b�}�}��8�]:�;]�՝-�SP��)����]}{�߻�}_.��w���G�� �`�   �<�v�   :$ ��@��   #�  �-   �]m    t� ��Sl 8�$��`�� �	d   )@�y�5*W-X�]��@�k���K����P5���&�5��UV��2 R��ڒ��6q��m�q;(q�V��4��@ ��m�mz�&y��v:�Y[E*����	�kiI���i�*ԫ�w�<�� !MU�S�&y��j#t�d���ӌ4$��R0:m�[u�WY�(2Kr��"�7j�e`=z�n�*xÂ�IgP�]��.��M��`y���zA6@|�=����T���ʹ�N��� �pUJ�*��i$Ԡ�t�M1\$�D����;=v�ٹ�k�U�F����8��vʬn8���R�Gk�m]���YE�ud�3Y@ۄ��Z΃���$�5�Ȧ�Hs���Mv¤��/^�u㭒��96��V��i����{ 9g��s����A 4P�	t�n[@	ym�v_bD���6�˸u�[�ۀ-�I9ɥ`  m�o6�I�a��M�$���$�   n���k�Ŧ��e!����ڕ� ̷,�    m{ 8ej�jc�P@,6r�X��(*��- ��ŲʵSN�
�T9�ݰ��p��%�%���m 8HP��S\SV��  ��+��[qď�v�������$l d	����UW6��i*�^�4���g�݅`ڭ�ʇh�X�	{leƎP���e%�ƶ�Nh� �@ۚ��b�n	�H �\  m����:X�[@�$9��m 	u�RN[@H��c�6믓�v[@>�@m�� �lXe�)p��C� ��s[@�  ,16���m o��i5ln�v�Am$n{.ݒ���`�V�؆J&��b�6� ��1�g6HF���%Z�T{�	  �`7m����[A��'P  ;h�,�ު�U�nͮ��s ����W��H�x�5Tkj��av��n��VͶC�����0mm���l��t6�`���IÃ�6���5� .ٍ�6ٴ�� ��=�[��R@mR��[U/'Y٨H�L` m����D3F�n�0H[D�"BI	$ ��Ŵj�$�$�-�p��8� ��m   �  k��m � Hf��Y�l [[li1m�� �[Ku��ڶ�-�   Ͷ �ۯ\��  �� l� ��6�m�  ᢭��kk�$ 覨 �(U_�|�z6� �� I�I�� �:�  6�� 9�t�e��R�*�6���[�yG����N���m�-˨�	yj�\� ����r�l�Pm����H��-��٥Xi6�[Kց!m��g$`m��<f�z�Z6�n��#pfIg ��/+��6��X�����$6�ͫ`��eX
�	�����W��M�[%�GY#E7e����X8�B�.�-�=�m� j�-M�YG�HoI���mm�%� U�����Z�UPe�T�ەZڮ����t� n�[@4ݨ$���g X:�2h-�$浭��d��-�8�   �Im5�[RH��E���l &̣�� d-�m� 6�8 �c���z�li��   �`-�H   z�m�w[���$ Ӧ����` ��F��i m���5��qL�@   l�kp���� Z����m$���\m� �)��^Z�}��w�|w݀w�H���` ���I���]0��& �t�f��8	i6��E���GҮQ��u��)-T�	3�� !m㭲H��(�nĀ$��Ŵm� gKz�v�[t� *��iOKC�
���
,�z�'�R�m��n�H5��q Hm�] m��5�Z��5�Fٵ����h� �m��s$��՛cd���ݜpm�mt5P� �`��:`:���$����s���@Νa�����m-���h[v  .�Im�[��d[�k�4P[vӌ?}�}�}t��V�	�e�j��� �ާ  [D��Ia���8 H�P���Gd���luT�KT�q�d	V�{`'8���u��M��%\g2�ꪭSPN�8�i%꧞\Q�$Ud���'(�����UU�z�-�v��C�l v��&�@k5I��Pe��tT�f�^eUmRf���c5��N�p���6,�Y���d6jU�.���&�ȲIu���m�6�0 9Ҵ��ݛn 
���GZV`�^hs�j�m��e���lK,�5��\��[@  �[pX-�����V8>�� �{;�Nݦ�T�̒d�V�6�	a[ :I6�I��駕n�H�ʪ�6{���<�үSI��Ai�@[Tq�xP'ej�(��������cw1�1RQl7<[�*�jU����*�� J�B��X��ۦ��i�RAR�(n�Fu�-��0��UX���WU�,��ܨN�UU+���ŵ�v�m�$4P    .�mv�F�a������ �sm�vu�I��l9  �l��� �`�� ���m7[{ 0p��h��c���E  A�� lm�DQk@	$�`9m�bt�q�i&i6H�	�\5�-�*��U����鵶FB�:�6��@��m"Z		����[w9��pbdc]� �[@[I   m��qm�!��m9"Am8j� ����O��-�� �a��Ͷl2H ���Bu�R9ٛa�y�̀�iͶm��M��$�   Cm��am  � 	�=m:�ހ N�� 	 $m�-�6���H����m��b@	r��J���t�h�!��  @ݶI�m� M6 ��v^GV`J�]UURUU�R�J���.ԪpPR�(6�Au�,S��WD����Z�6�3lp�qK�� ��)�X.��[�ڷ4R'ggn�ɣn�9���݃i2��ͤ��@X�I)"��e�$ �v��O6���k����pԀ6 6���vC)hm̰��6�U.� �;T�-Ү��U*�����r��&C(J�pUV��VV��� 
��4�:�@-��`V��m�yw"�˦��p6��]��sLUqU�II��[v42�Pq�B�0N5�]v��zme�y���Y�H���yӹ�Uj�\��
�����rG6ذ�EB����
��M�p�[@8a��$sm� 	��� ���\e�/C� �l����\pm[`�I3��  m�  m&�m���;Mpg4��B�����|u׷��] �k~=���ަ�H���m�m� HԝzԀ   l[@ �h-�	 v�  6�`n��`�@     8m����` �A����m�`m� �M�)<�R�>^j�m��       � A�$$m��K�it�r�[F�Z� -�e�%�WM��� �\�` � �m�6���ӀH$ �e�6� 6Z �-�@ �   !�R�u��[m� pԴ�ۀH6�   m���  �   6Z �` զ� i� [@�=   v���-� �Z�Hf� m� v�R����I@[2����6 ڐ���M�-��T�J�V�)v��*��m�ɒ�m  �����W`$�:%Rp6� lڴ������$2$��Ra�ڽ0m�m p  e�M�L�v[�m�5���m؀m3Y��N���c���[@m[B@�skj�n�6�m�U�lm�p    ���g ���n�m�`��6�vY6��كc�S[�6���F���@;Z!��l�m�UP�R� �;2��ص��d� H	���uUHHUJ��{Y E֩�ʷDi�Wge��lp��Z[�x9��ٳe-P�|�����<�-p�Z�Vзu��p	�5�ֽ.�66� )V�� yZ�e`B�[@� $ �    BM�� ��l�m�C��9�m���F��6���� sm�	 �ۭ`   �6�  �ζ:^�5��[@�h[A��9�l       �h ��}�k}�l *F�2 @ �lm�� �m� m����$q��UJ�UUJ�[mm   8z  6إn�k[���UJ������9�\�ɀ�-�Kj@ 6��d6�@*�UyW�s-�UN�׶� 8  �h�    ��	gh�I������<�����ἠ�����l �������h��"��,�"�����,�*s2�2��*�?Y��"*,�s�����}�"0�0� p�����o���U�DDDDDDDDUDDDDDDDDEUEEUUUUUUUUEUUUUUUUUUUUUUURR%P%	E���RU�!@�f@��S���������ڧ���I�H��� ��=��6��vpE�`t� �� ؗB ���	(! �� 
=�J��  z�ҩ*��	)�!b
i�7��7�����)У�"8*�t��&t���誌��m�@6�����^��������[CH��t�k�'�)�{�#�� �Q4���({:� ^��;GA�E{W�  	��A�%�}$ ��@��]� ����h��x����b(�h |��ACb��L�6I� ;p�"�!�㊽ w�|O:z�8x� =U��!��qz��T|A��:�b�b$�=���=�S��A����F��`�y �6���~�b���i�qUd;�z�@�C�DSf�\�F�=�v=	 �h҉���r9�A�S�A�1Gz��;W��У�E�<�T�A ���{�UEUUUUUUUQUUUQUUUUU@                        UU����@W�.��j�#��������_���?��k{�o���{��������$���AEB���(T��%402�D�+JГB4���o>�F��k��(��WbT�њ6D���;r�j�nJfr�����^�e�v�{�H�$��h[Lڶh�Rs�H�.Z��=�:�����R6gj�V��^bٙ6�-�v��6lգ�봵){[)��HӦ^Z�*���9� %��;j��DN��8+h���u76�Qu�m�K�^+m���n��]s�Sk��8�����&�8��DȄ�m���?�=}��s�h8�lշS�oXvX�:�F��{��)�A$�bp���*�I]t3��f��;l��P�f��X�3�;	i-��a��<F��<��ku ��[�H[5�#m$��i���\ ��A4��+��3�"Ƥ��e:+�f{n�M�����~w��~~�s���$6W�iG��C���4�D�gv㓴`E�r:�2��9�-��3Oe*��5ZV�`F%��5�<�l,�֪��mqR�5�Ѷі���	Z�˰��n���ο�d������GZ-R���l�V0�z�A�mX����_4����Y�8�M�#p5U��e᠞RP4� Kks��\\9V���& �,M-�����n�h�Ej�e�J��l�۠��j�kG>tHU��	��E��Y;��oc[���i����6<g�ѲcQ�������`x)U��۬�5�먖��(,n�����q,�MUI�k$�gk�ƍ�9���^ZڝA�Ȇ��Kuis5$��i�c�:���l3����}۷�	���s�3�8�K�8�4��8��zy���J�.����=�#�\^^���9'����l�k�ӡ�m���Z�
���_m�GOL������!t�m:IkUq�/��4��Ҳ��viU��[+e@kyض�h�kX�VUBeU���P;k�����i\m�p!��59T�C��l�"�����h��y���fN����wC�N�j��m����<�spHһ ˡ��`
�j����M�t�$ݯ6$8��jꪪ���q��@@J��V��42;��n���eWo6Ռ@T K��(|�/��I�������@���+�^��0O��A~���	莎f�^����߄���ɗWj�ud�L���u���>��J�;\��tTsl�ѝ���n�)>n.�i6타C��m��a��ݭ�(qF{����ee:��5��2�q��t���F�6M�4�ۨkq����ض)�rj�T['�r�N�O<m�.��+[�
���r��j���9�9�	�;��Wo8�!ݒ=�FV[���*:�]��w���2�<"�l�ێ|�TOs�vݗ�60��9�y�����e�nù��]��1%��8���ybK��Չ-~6�6X�H�G �C^}ݼ�(�(E.��Ձ�ɥ����V�P�`�%	ے9r�%�n�.怜Iw��1%��u��Ҍ�(��$���`}��X��B^}ݼH)s۸bK{�m��n%$n+�{.�/���d¬���~`g<�6�c�q�4�(<&��66�^�yܫ ^,c{�Քz{gurl�b��=ĸ˒�q%���ė=��%o�=�����K��n��q�,c��Kė7w�#J��HK,[3��jr�y����e����c��QF5�M�M�AN��`}�1X���/f;��u`w�$*Y�F�N8�{�f$���y��n������Ik񷱲�$�r9�Iw��x����É.��U��{.�W����@��	Dr1�FQ��Y�v��n���	�H�;�q���/=�v�J���	� ��X�˫�y�����bK��kĒ焗�[�I ��bK��׉/{ۆ$����H����^��X�)ӂ�$��=�eՁ߽0��S0��.�FĔ�S��eB �Z�R�E*��w�bK۳V$�wF�V�i�B'$��.w�V$���bK��Ո=����A���6,�IӨ�JB���pė;�7�{pė}�V$��O�e�p�`h:g����˶���&^:�>�X۔���}`��nU��!ە��<��ڌ�T�wUŁ�m"��I\X���^4���DIȰ���9�{p��3�����oce�H���%r;�n���n��{dU��𝚭��ܗrL;��Fw۸{��]*�*��AL@���@t�Q4�Z���U��ÎY$�w g}��7v@�}�Û�ꪪ�=��'�����b�&��v%ս��Ÿ�hw �.<����/>�NǓ�n^7==;�`�����I:�ϷU�$�Dp�57p��hv}-�e�;�K���ۇ7vw��=�l�.��Rս!nr��n�ｸ{���{r��Z�A��ո��ｸw���{p�`{|�L~4��wra�{`|���;�};�n��q	G	W }!B����A�C H`X)��Ҍ��j�^޿���l���5@�7N�b��w4��kX�Z�'B��@J��d��l��py���$
��k��h���X�5�q+�.��y���
��N��՞ևpn��B�t"���[v�۶�u�M����P�6Z����eW��҇m���l��p��N��Va6����e냥�R�F��..`�ݦza�Ã] nz��2pA;�Z�i�{���T����:��g�+��c�����C��,	D�Jn�n;�����;惞:�hm����~Þ݁�����G=��;�Gݹ.�w���(G=����w��=�$�z���,�A���{pｰ3����m���^H{�ډƤ��Q`�U�߸���9�A���+ۣV���l�N��g����m����;�l8������~�!r�\R۲��������[b���v�/���]�!nd��#����]P�M�9'�����7��;���KUޒ�5n4�r*�}�ͩ@�v����H�)���iP(;H��p��Vo�i��KQ7q7s���#���;��U��Zm�l�����RJ�{�}�߯�]��pｰ7�^��cQ)m�%��[��ꯨ�~߸{w��M��ڐִ��=���Jh�ȩ��=�@��=��ۮݮ)^m[�ŧ�6��OQ]��w�{p�{`w�����u������q�ԑ��wv [7���>����������֒%�m\�\����᫾�
���46��TV��&a��nQ�-F�zԉ�Cq���j���n���o}���6���#��-ƕ�r��-�{��ww]��g��cP�VGm��j)-$�h�r��ۄ���ku�W	�|k�����;�s�N�dIɆ���������ۇ�My`���QHJ�w���W9F�����6��{%o(���P��D F��'.��6�o}�n��#����%���\r�$���߽�a���s��"��TQ��T�wo:4xw��\n5$w0���Y����~�\�|����p���4�M{n�@�Wv��$�2F��X8���j��=sJ��t�N���ӑ�*��f]f/k�{�ܭ�l7�M]�P�Ke�hrL7^����R(��gvo�}��#��ܭ���#��-��r�{��7}�3���u�]f��ך��V�K"NL9��3����~�\�}���K�����ܻq��3���۷���Û��Ue � *�ڥ�*T���q�H�W:�mG1��F=���[g�u���Ůo3��Qɺ�b㍐Ps��#���ٵ��1�
Q gEb���8� �����\�;���b)���_/�u�L��g˻���0��2�@�.mrq�]�ԻpU��I�z8��!�.e�(��x�j &�'+2gN�R8'/1�[�6C��(� �m�ɮ�S�\���)�mQ�ʻ+L��R��+$wY7�6���qp���=o6���5���k[H�w6�����wۇ4ݕk=��;�%���\r�R�%s��Û����W���F�
�K.�N5$ra�݁�ww?*��-ߥw~߰�����[E�n��p=���G=���n��uh�.���r��MI2��l�����o�;��{��]��p���gV4��n+n� 
XC�*n�;E���3����ud8_~�~�4�ev;7")$��wp|�������w^����Z?�D��ȓ������>8+T t�H�D����}��������yx��܍\w-�$n@�{w+˾ۮ{��9��|x�N�
(���w0������l{۸s�KK4��I ��u�{w���o����<�����;�@���-"�[F�1��k-���ǉ�[^�7[{��:;m.�wVݛ�S�N7<����5���~����p�����7�l�;5�"ܷr��s�)j��u߽�<9��|#��W�_�5n47jI��o�\�n�����>��_�^�-�n���m��)�DG@�����?�Jl0�.odc�^No�j�����l�'zzxt8�R�o!��Ț���52��Lu�D�c���SJ������P��]�`p��./A�T�� ��5���kfM4HFf�&�,ݰ�{��*!@н�GL�<PtD1�0�	tj���h"�L���ֵ���k �0G{� ��}��w��h�5L�~����
���ԯ��")�Q�?!*�=_�� �"]9�@��`׿t��8~���%=�~�)JL���uΜ�(9VWf�4o`�B��*{��\R���������)O?}���({�߾��A��8�����ָ�)C���fe�����{Ѿ��s�ԥ���ÊP4����pz��=�=�\R����o���)J~  ���24�~�����޳Ւ���7h۶�us�')�r��֎6�h.��+��AFe�)��{���I�~���R���=�\F����߾��)Jw��p�4�'��{����v�z���oZ��JS��ߵ�? 3�4>}����)O?}���);�߾��%)߅_>�ky���Vkz�4�~����)N�����);�߾��)J}�{���)I߾a�����֣y�[�9�s�ԥ)���ÀҔ����pz��=�=�\R���`�J)$�,01�H��]���|�^o��pz��>�?����q�ݭo7�o�R�=���pz��$'�=�Ww~�*�T7�*���j���MTB�8Žw][�fx���0�k����A�q%/Wv7+�ӛ\0��}���{����<��qJR��}>��ԥ)����J+��ۮt�(9�3U7�M�SR�9�޸�)@w�}�R��{�8�)I��{��JS�4{�qOᘥ��H�� MT�H�]$��Ӝ��+�o�p�);�߾��!��O�׿g�h}���+�����5���nF�;q�j��)JRw�}��R���{�qJR���~����{�)I�ǿfk_��R"5r9uΕ\r��5]W�����=JR�y���'�����)O�z���_gz;?FtkF�,���F,٪�,=����U6޵���M�iG�L�ٳ7-��v6�sF�K�Rn��T6{M����o����ڽs*L�S��6:�v�u���xǭ��N��N��H*7�۳U@��s(�����+q�N���m�#�����7`���uhu��D�<�^�� J�/l���Z�˲��nZ7_fq�V���[��ϻ�u�m��m3��n㞵�n{F�E5�Z��֍rlu�jݗq���չ������ַ�┥�?��=JR>}�}ÊR��{��pz��;3Ͼ���P���}r"��S��¸���<�߸qJR��}��/R��y��k�R�	��}��JS���VZ>�n5��k{����R�?{��pz��;�>�\R���Ͼ��ԥ)��ÊR��y�XR��j"����9�r�^�wĥ(~����)Jy�p┥'������Ps�f�Zӭ�l#q�JR��~��R���{�)JP������R��<��qJR�����fK��]Z-��i�-���u>��q7�ȅ��b���wN	����� m}��u������ԥ)ߞ�ÊR��{��pz��;�=�\��)C��߿pz��?g��~��n5qێK�.eP�P��w�q�~��O�|���o?:���!�}����)N���S�b��z{�3_��ݺ޳7����R���}��┥�����?FJy�߸p:F\��W��߮�Ӝ��+�l�S���N'$�wJRk���Jw�p�4������)K�=�|R�����/�D]�7"��&a\UBA]���U	U?{��pz�����~��(z�ﾺ�Nr����6�.6�c��pi
PP���'�;�b �=���g��wW�a8+�g����5��z��)JO����^b�)y�~��(~�߾��Jw�p┠r��q-��n$�:Qˮt��Up��~���JP���}��R��߾��"yA�����:r���H����7��Z���)K�}��JS�=����(�����x)���O�����)K�Oo�R�=|{��^�Z��ݽ�����)ߞ�ÊR��{��pz��.����JR��>��SBUG��o��!q����2�J�J����=JP�X3�~��JR'�~���R���~��)JO ����n�`��E9�\��69��n�tvwl���V�M�C�N�h�[������y�)J]���┥�}��JS�=��)JO>��=JR��E�����o5�{��5��R�����pz�iN���N��JO>��pz��;�=�\D���߽�_D�ĉh�E�2fUqU�~��)JRy�}����=��\R���߾��ԥ){��a�xF�f�k{����R*Ry�}��R���{�qJR��>��R���Q:��P(*�b�h`V�dA�e�8���_C�"����U	U	Q�y{��q���Z�a\T��~�߳�R���}���)N���n┥'�{���)O�������\��d:g���2Xb�k<��C[mG�8ۯR���v�l<�����?<�b���vo[�)JP���߸=JP=���8�)I�����R��<��qJR��}��Vh2�!K�˺�Nr�����u/�����~��ԥ)y��o�R�>���r�ҹ��+w�H��Q81�*��%'�{���)K�=�|R�ҹ/�����ԥ)��~��)JN�<�3_[�kv�z������=JP�~����)C��}��R���~��)ZO���=JR�x�:qG�$�rK�(9�
��wmz��?�}��)JR{��߸=JR���o�R�������4e���~�,���/!۪ʑ��� ,�:������3gI".{^;Zu���*���)��g�]���yd̼]r�'�)[ey��y�E:�&�'1n�C��+�n���\]x�݀p�5��ܶ��q���si�b��"dx6�cc:��ݮ�GAz���3���4�L�8i9��θ�Y��[Z��IGs�,��q�WW�u.�x�[��M��w���c�nN{���}�w;��ݹ1�&Wnۗn��=!�A�TaI����J�eFTR�����<U�%3�s�ÊP4n~�߾��)J^y���4�}���)Os�#�W�N�nַ��[8�)I��������$�����~��({���R���f�]s�U��o��[���J�F�pz%+�L����)JP��}���)N���R����~��ԥ&����TR�7B"��7%��sssn��JS�}���)<�߾��)AKw��ʡ*�"����%h���L�]���)Jw�p┥'�����(�}�|R���~��}��R���ߎj�O���a�[��dy5�[=�6��ڜ���%�]��c&wm����e��x�)>�߾��)J^���┥/�}���JS�����);���5��V��R۹q�¸����~߯ ��h+
���`hW4�փ����~������ԥ)��}ÊP4׷7n�ҫ��Vx�:c�����|���Ͼ��ԥ)���ÊS�U=�5'����pz��>�~��)JRw��c_D�KDp����WRUG~߰�JR��>��R���k߳�P��!��߿pz��/ǥ}~�k	ޭ�����g�)<�߾��)Jzy�~�'�����=JR����8���no\s���)�*����PQn����:�-��l]�[Q�ݞc'�6nt��o{��)J{�{����C�}��JS�����)<�߾��#JG{���*n���!D�r����g�v�+� �Jy���8�)I��~��)*�_��2�J�B+�����
��"��7�o��)N���R����~��ԇ�=��7�?�ùMf�޸�(��W�W\ϗ9A�Rܥ��&�j6܎���R����~��ԥ)�y��┥�}���(<�ϵ�)Hu'~�j���$�ˮt�(*��ٮ����}����9)���ÊP4��n�Ӝ��+ۥFҧ=��QSl�\�q�B.{]���k.Nɺ�z��p����ٸ�tơ��#�r����r�ۻuΊR����8�)C�����JR��~�T%T%G�{F��2��efff�H���~��)JO���=JR��{���)K��}��R�½��k	ޣz����g�)>�߾��)J^�����fC�}���)N���W�);��s>�����ލdZ����R���߷�)J���=@ҝ���8�	�4�$��$��J��� ��!bI$�H	)@�Z�ifX	�J���`	$H �(�g>��T?�g��T%T-^����e�b�V�����)C�}��JS�����)>�߾��)J{�{���)Iн���?��5��C�F�۟k�WccvӷT��5�uu=V{V�/\��������֞��k|��)Jw��p┥<�߾�{��~�~�\⌹)K���~��)K[�W�I	�(���|�9A�������Hd���ߵ�)J�����J�����);���fk[�n�oZ�����J�'��ߵ�(���=H~Us
S��~8qJR���~���Q ����喭�����J�H�|�︽I�rS�����):�߾��)A�%�^��\R������_�{��ַ��|wÜ�=JP���ߺ8�)I�{��JS����qJR�����R�Ds����ַ˴URT��x�k�G���(�%���#)�O`
R ���a�4�䗚��a�ʜ2"��ՌE&�A�HS��� ���� "�(�$(bR����Y �i��3B�R�����Za�B����X`�)�*��H�BA�Im"::ܦ)w�r��9<t�2�M:1�%GF���3BQl6�K�)RP�ҁPT9� �2�-KB@QR�Y��$�2Xj�b�Bd���O ���^�uo�L���ń���<m1k���rPE-	B0�Ħ�`b�.���]H�Z�8�LV�n[,�Z9؝A3քp6F*'�d�LT��$��"f>۽�h�� ՊN��P@�C1$�
U2��8CDBHI��0J��K RK3!!�΄��ũu�ޓ�8�,�����z�$�߇�	�d�AD32%AhM�+B�P�QY��J�e5*i�d+�"9ʠ�����T���o
]�J���}�ۙ�=\u|.~��k���,k,�R�k�����n#N�
Vێ{2��kt�m��ƾ29Syv�Y:ys� �qՁJ��hN�ʛ	����t�������s�ts���:0���1�:��"��h�>z����c.��Ru�wT����)^M�d����^\�q��x��F�!���y�c����;��.�˻=]���a���r�gr�dv�[�m���/A���Y��������g("�O�up`���G���«�q�U۝β�hq�(mE�H�]t����#��%��vU��U�54�ZZ�68���+�]�ڨ�'����l��Bl9�Qg�]�n��i��z��&�3Nj�Mhth�������3J�G=�PAv�q��5�Z�b�U%C�����RvB�c5$��q-H���X(��U�6�"�S�
�L:���ݹ3]�����`z�.#� ����<k�t$Mmm<�<�خ���}aÌ���&래vG�۴lC�!��I�\�]���pv`��I�:<���[���a�\4�J��)�%�s��e콬�1���Ƿfi;a��1�����e��i[-3��M�����&U��9�a��wM0Kf���><��q5U5Q�h��L5C�ŤvM$���H�yT-�tC\�>�ʝ-I-ˑr�Ue{;��6Gi��m��z�����6.��.�8��䃪�.��
�yx� �f�p�9m��#�ٺ�(=����k��6�2+i�'-MU*�� ���
etZU�s�B�m`���kf�쪩�K��	�+6���[#*�;������J�nS�T
��YZ�V��Ѭ��W�@�S+ܛ�cv������W�9.pݶ'�����|l��*�����휾�ԓ']=im]S�ۋ��98�m��9�T��9zb��Z����nګ�,��H�9&�k���A��L�mk[�\v�JK),���tP�<�� R����E<=��5��u�v)ڧ�0�D�zC
(yÊ��Tﺻ���s�m5��nDW[P�p7�00��E������ú�Z:Zё#��G�)K��7�6n�7'e�g�Z�B�F۞��X��o4[?|��\X��b�h?>���>��v�#��m紬�,i��m��E���z;.�p9Z5�n8�n��1�c�A�Z^�-���/a�k�S�N� ')��h;����ngpm�ܶeSU͢�n5�G]�¤�t�YP�.��z1P�����}��5�k�mœk�+�u[�/.�ם�(����خݨ�-=�nP��y{n]��z�k[�����JR��������R��<��qJR�����R��}��8�<��o��z9JEJ�
��9�p��߷�?���JP�����JS������f���J��%F"�(#]�� ��N��wz9?y?f ���~�+�~��H?~�T�Ժ�6��@�?\X�<��}� _jw��ʙHoTUmI9Vwٽ����>�m���sn�̣x�4�m7H%y�v{��q
=��6�Fd�3�Sħz�K���f�RG�8����]�g�;�
�sn��{�3��R���"���vW�ߟ}���l�� ��`���]U]0��
�9ޭ��������8����ܪH6���?Q#��"�%�˞���q`|�<��}������$v�:*B&Ԁ�a���oz/f�O��`z#����E������5T��Q<;U�)�O���9��Ł��ozk��,T�*��&2JI����p�i��hIF���U����3�9�w~w\f8�n:m*$�Q8�^��҃�ͺ���r"9G�C��� ���'���GQ�ws�}��WUԏ�/{҃�]���͝���lHM�MSm�$�Xy�f �S�\��Fr9�Y�r��X۟���^��)6�#��UR}Oݺ�k~��B[w$�'i;�>\+&�1�E%H�������`eW(��u\X����}�} �>�DpF���5�=�;z�H����M`ݝ��S���fpmʎR��G4H�;ww:ۛu`cI� �S�r!$� ���=N����G�����^�v�����>�۫�>�N%��$BDaMIސ
u>� i�N��X�<�s�����Ң@�������Ӡ�����ߺ꿁�x��a�fbA�iu&ݠ�����k�]w�,�� b��;n\�ۛ.��7�|��v�~�}�r��R��q(A7�n�2Ru�۶{n�v�t��\&�Z'���]��]��Bn&��ڒ4���{w�Z�m�y�5�J�͖����r&����f��s`}����$����7�x��jQ���RRjE})�s5��X&�`.�6��$pv�]��k��˻��3�����ـ|���A���_@�PSͤ�>HF��~�� �Dk���5u?w�N���pV���uZ3=ӭ ݆o���q��K�%l��͑��[\��I!����i�Hɛ��sBK�,k�n,�2� �.�0�6޹�Z�8eK���E���AW����(��K�9�x�I���A.�J�s="y��7B
G��H���z�mh y^ub��k�c���LS���>��8vs��1���)icS�q�3R�+IU���n�y�n����R7�#r%%��FQ�&#�m��]�M�]�VX�g��;v�Խl�Z�:v� �`s&Ӆ���
K�1vJ��� ^�6�����w����Hk��� ��U��鴪(�(�=�7_qH$�Vk�������5I29r�GQ;��@=��`}Y���y���u�
�Ɛ�`�M����`|�y�}�nl��7����{`G`��qIއ���V��+��{�w@���>M��qD'��ńD�r3�����M�m�mעSp����v85�X��{s��h�w'
�����"��R+��{����&�/�5u��
��v�lNF��wo����U��E�Us�����*~��7{�M�ou>���""dj����m�R�A�%�{~�@�������_@=��`o*�Ґ,�J$D�]�Uf������� n�V^�߿}�7�76�E�V��}Ͼ�Ci��5�y�}�nl������m+im��;��pGX�=��7X,��ڍ���cv�q@���O[;֐�9#��ܹ��C�~m�z��:�lىdcbi��T�>���W9�r��5�ޛoW��d>�U`/�A�Pv��A��⓽�{��|�������X�����o�VT�&SP�JmH�
���6�j�O0��ȃ}O�`8�t��N(ؤ�@����l�;��ށ���`{��V�Ur�fV%Lth��@=���p��X�wnC˵�X7�3m�t�oW&�E%!A(�ʍ���~����>ך����� ���`f�q-�N(���N��� �|���=��X�s{�7U��M�QDR#��-{�ljUg�}�~��7�~� �rL���FT�������W��������һ�^����x:�UG��|��ʼ֐��))��qFܒ���f��|�5�%� ߵU����x�z;҈ ���05���n�L��t.N��Rq�F���͍�z4�v^tRA�M�/���W���l��`������y�� �dL���r; ��c�}��ٽ��6X[�V�D��R�v�}i�G�Մ�<���s��L�S�l��}�;^(2	c(#*7P����f��m/f��[��=�,��d��	К��W�]�ջ��>�K�}��uW�;@�����יoF���zNs���F���K�ɻ��q��9랃������]�3F�ݬɺ�E�g�)۷dwm���|A�p��n۵�'g�|�.�c��.�v���[��݁��N�5�92/WlP���Ѵ5��Ju�(�[N��Z�ڼ����VN�U��m)ՠ
ӝ�`���M5�7V{Ncq��&U,�eҽ�f���;���;�lԲ1�G�)��a�(�뇮��t�;���F��:����F�Bݻm[�� z��^g@SX$�P��*�#����g�`��X��ok�j�k�>_/ A��QSW��p�V�O0:�l��o��q�n��m7"�I%����z��]�ջ��;�d�;�e��r6�ڢ��0�O�Kk��%V�_R����3J+�բ&SP�J�G�@�X|�j��y�	7V���yL�~�)ۓ����3�Χ�7�m�7nz^�au�n�v�8,����<��:�!n���/C�'j���I����XiU��@B���(�	�,(�����U��U��r#����S�Հ{�U\��%W߻�=��+�J$BDt&��@>�l�
�̖iŊ��nX���@=庨CqF�ERE�U�iU�g�U��o0�w6X/�!#5�22��]+����j�8�n��S��%�x��v/�!�zz�uV�ٌy5�Ӱ.�����Pݨ
�H��l����;�:`5��NX �U`?{����N� r�������ۻ,���ߣI��29�w�|���).ئO��X	�� >�Q�t�r\��K绷�%���X=��wv���*�%i%Iv�D.؀���"߲,ZL���8YG'�u)���;��M��i�iuPPy)ڡAS��:�)�ؓ��:4;NQk��n��h-&���h|����ց���i�3[Mh�!��:D�E�lz\T��y�q��ӷa���=���8(t"#� s���@�}D�GI��O�G�v�a����b> l<9�N"�[�:�^�vx�u��}�Uy���\�Њ�H�6E*>�B*_{t�}���y�V�c�=�A,dJ���A�;U`$��2gw�̀`��g�U��PP����\�JdV�BH�T��-����>{�\�6�) ��Fv����	���j
H�C���5fc�������@=庨CqF"(�(�5fgl�2>J��y�F�S����Dة��;�!\} �۲�3kwo���VfM��1~~���Hǎ'M�$������y�n�9�4�a�#�Mr����`fר���N(����s��#���@�`�U`$��Ϟ�d_a۞���v�.��[�<��{�ƛA�m�{F*m��mV�7ny�����J?6y���*��y�> ���
�"�F�Sq)RvH����37w��<�`V��v�/�PU�"n�uPw�U�&�� �z��靟7� �S�ߵV�ĤR���mIށ_y��K�����K��w� ��W	;�Q�DqG��s������e�-_�~몼�^������b��hVQ�hLpЋ���1��(�X���3����)��+� ���.�]�`2F����E���k5��oc\�8(j��a�OW;��[��Fuv��kj��xN�x��v}E�U)&�g��4#u��]Z���x㔎6/��═"�0���O=gP�6�Qcab��8؊���g�ͦH�hv��-�F�����p�e�X]��ђ�
!=�H��(c)�N��vZ�,�2��sm�����۶c��ݞ�@��SL[�]����}��������9�!Σs]�=�β��`u�������Ӌ����ζ��2�� ЉlT�ʊ�j���~��M��7z��@�� k�#��W{�jE�Kw۽�s��皬[���{%ď�^�vF�!�9NI��5u9��g�G"8H}�Հ����>��EeG����NRjE$s%�dϒ���^�y�F�S���2��Lu��r>�}��`�nn�@��j�
���`}�$�ۜ	J���J�k�ృ�]�ç�=u�(�j�o[Ϟ��(���� ���B7%������Y���ᏕV߳%���U��R9BDm+{�]U�����>��4 ���{_�+�lߵW�!��o0#�n�Gk��R"��+幎�;��YA������U����RT�ʊ�j��}I{5�nn�F��x@�-g���3�#�܃i�Ԓ]����y�+=���>�,��̣x� OiF�AE��{��ue��1'QƔy��yY����շW(���ir����#��=纬ԏ<�`��,nn��Q�V6���U!(I��|ҫ�UXA�7���������)���.\��{vX�ߺ���#�b1 ��+��*H@�a
�J'����ߖ���V�ے���F�R�ƝBG%��M� ҧS`4����U`|��jzԎpUH�w�y{5�+�̖߳%�������
ćT��ԉ�c�;q�3Ãlp�ۘWVn�]e����W�\�:�G
nTcEE��} ���`�X��{ӮbI��퀧Y�"_�g�������`ڝX�y�}:�l�,(�4�Y���N�$�����0u:�f$��J�>J��#aˠNH�E�w���V<���=�vU�b�U��g9�\O�����QSiB'8�����ݝ���,(���z��]��ԍ��
�J"*NJ�՛�;a�:�mV=����]�b�^��ٽ��{�~��]A�d�%��nO�>��=�[����k���_,��=@�F��:�����o0��>����Z]� ϵK� }���=jI%6����������`\��� M�����w�+��TQ�K5UR�y��;��X���C˜熞l�<�����I�MTT˛��ڝXA���}�)���Ҫ����zQ)%	U^���>��/���`L5����h�)��mu��ٶ�]0q��G&���9��Y�k�X�]�(;x�xxAk3����v�<;���ۮ�V���Evۉ�A�\s���:j�,Ȼ�;�2�k];�Wq��<�Թ�:��⛘����;s���0����~9>�qێNԧ �kv+�t!�1OUeޝ�YBf�j�b�]]�K)�!qeU�@U��o�{�����|=����L-�5��	������;m�om�^��-��n�Z,�Ʊu������!���[*ᴓU���� �u>�S?KK���UXh�hR8�E�����]�����)ϛ�}�Ձ�M���@G� *�M�B))G`|�1�~�J�=��ށ��k�2�ܠ6��2BGnG�9�����֛����a���ۮ��P3Q���Q�P�I`{�n��|����̖߳%���#��T��m/N1o�b���L�m��[,��ud\��v��LEv��NEUjԄ����D������">iU�gڪ�ȈZo0[�
oj1����n; �s%���_�k��ܮG�s����YV~�߳ �u>�DD���i'%5QS��N�}�͖�7{��M��/ۮ��4�Y�n��ٮ�XG#��7�ө���ZQ��\;��Xz���B��Hr(�s����`{��7� �S����&� �D7�^����=�x�hꝳ�m�n�ե�%ƴ��Ν�Z:힌���_����o��^�4Iڮ�KK��j�5�� ��u>�_nPmF��Jr��} �0�u�@�y�ө���Z]���@u�Dr'P�$��n��|�������AI,Q2Dz�u��{�\�f�>���V�	!IP�I�� ~߯k�wo��}�� ��������¿3�M*�q�-�r�s�gڪ��y�}:�l���Wb��]�V�zK��"��:ݻv7v���2��cm�R������M�?�X���W~ �S�Zo0�S����`-�c�i�J9,nn����*�#�7�<�n� ��ج(����B��H�G#��/f�幎��P��.����zޠ3n�t�mH!��8.�}��i����G��FA��p""))A{÷���
>���5�++��A�r�!#��#�P}��XQ����^~���~������`}?
`��.9�tk�l�\2�sca�tq���<�]���xN��`õ������G�ozĬ]�@������`l��ȋ ϵU��sTfԄs�P���@�{5�+���;;2gڪ�i����LHG�<#�����J&�r����ȥ�� �R�� �m���jv~kF�͂NH(:e��ҏDDDĦ�V��� �u>�G"���y�B�YM��܊%��^ozө���Z��j�DE+��|��T������D���p8"O ���y0ޝ�: �!${;�1�7�;�&S��| מW@&�q1�$��3�g�0�tdʣ�O�J<���[C.��
�v(j)��_A�H�*A� � e�{���H�o0�!׻��1���a�5�t0�*���8�vjnwXf�N�
Jy��w.�:��Û-���H�D�oH���,,���%&$u,B$@�� ĩ�/�$�s\�)��fiO���|z�<�g��J�
m��9!BP��Zr
#\Q�{�4@�P|ΐ4bU$�Z�ۣU.]J/Owwn�Rg�}j�����.���G�}/��Kֆ,��l�覽Y�f�Z.ܲx[I�s^M�5��MAm(�aJ�j%�N��s@�;Nƺ�&��i�nwU9�g��=��v9ۦE��JI�tP��;����h(;96��m���9�5�ԝ{�$�:Nݵ6y��㮻�x�:;{���Ĉ]��u���\O�-� ^g�����T��*ӝ�{{FʩsL�ڦ�0��:���g����Y皪�6�oCj�a��ӳ  ��U΂�������)�/4+�Ky�IsXa h���Z�7gp�԰pq ��lp+��wE�[� m=i�u
��=����)�S�v4;�[�[�qlzۮR�\���M7�+r�'@�`��R�J �n-�l�jjIֳ`������R�Qm��2�rBnp�V�)�ZX�%�=�D�a-t�s.�Ê�C��ɒ�qPp/���.͝۞yCN�R��SN�"���B����)�E&j���kM�T[s��q����%���́r��ݣ�W�lt�0b�V�e.֗A����۳����M��R�N(z���8ڷ�[u��݌�H���og��A5Y�:ve�- �Vܰ�+m�+�wi�w�;sFY%o6� �GSJ�URe�V	w9�qa6��%6�Ry���e[zN	�G8�5&��^R�n����d�y�2M�l8�����$�+�6�tV�F{0=r�n�֝�Y�<B�9���S�����/'Z	�={T��N����M�KvZ0Q5�W:�'��eJ�P���Z�j�������h����(��4�n��U �r�,i3��TRԇ0T��K�֛�m��I�EQ�,5L��r��=l[m�C�vN9]ٔ]�'B�+8��7c�\����1=�K�r�P�)۱��9�ν��jc���:�V����N��m�lA�4l� �����4�*�5� 誕em�fg�y��vu� R�5���w�]��n;owøz��j�i�<�����C�����q�4�:� x�}��ا�@��Z�'�ך����w//!����R�8��\c���Z���"On�.ƴpGKe�����J55gt�m��Λm�öۭ��Z�H rͧ	m�-���U@���#Sۉ��uu�n���Q�gnq� �'n$�5��nP6�0۴`��=�4kF��mǋ:N$�XA;^΃�l�nпt�����mI�AZ�ٗ�[���s��tp�NȲM����N���~M��;�ۀ����I����>3k�Ɋы����;��E�v�gd�L񦊻U��ey���Z�d�j�[O0���+6�7M"H!��-�; �ڪ�m<�>�O��n��E���˪� }�Ձ����S�e���K)�&:�	$�	{w7��~xck��m�Iw�قK���''Cc����V��;���,n����U\��~�%N2Sd�����'Ss;;�jN�=��b!Ən�V�ꗵ�ݕ�:bd���MQ�Q��1~��`����ͼ�r9�GA.�M�r!
=Љ�	�UMY��e�溪�Ͼ�?����}a�����r(��~���;�OӀ=]��ɑ��n�Pm7"�I%��ߟ���|��j�<�1�~̖g�RڎF�$$R���JT�6)m��3�QV&So:ޠ7m�i��MH�,�v�"	ϵU��o0��������g�'?�l��9��7�n�y}��.�ݷ.�s��:h)۠��U��c�		}�@>�l�m���9�#�}�!l�&\2%%BI%��7w��<�`yfc���@}���mH)8!�i9;�>����^g�����:C�2�x�ݯ~�,�f�z��M�D�D#j�qX~�p�-��ڝXM��>ާ6�?V�[�'!"N�����͖����}皬(���`w+�aNA��Q�U����b簙�a{]v����U6c͏�|��3@�ʊ��Q(�������y���L�@}��`n�~K�)"T)]�f��9�6R]��UX6�=�{(��&�
9I���u�~�V>s�ș������M�>n�Ӳ�)�Gۑ�
>�l�777��<�e�c���k�@z�G^�����+���%�ȔJ��K�i���9�6V��}��Ds�����߿���\t�F�,�um�N9C���YMh�b�����֍ܙ��Z{���6��=��j�W_�ʙ�Z�`n��i�UV�7�m(F1G���~��r""y!��V��� �z����v��C��v���e���ސ�R>��VV{����N	��q(�777��<�`yg�����,(��j[�ܥA!"��ށ��j���}���y���9�"��Ds�������_�7��y�ap�8ԗ6^*Nݺ���� "<�%�t��2��V;uIפ�c�ˬ�s�4�c��ĮЙ�%I^;vk��srV�Ԣ5�M�s!��3�`����s��qE�7�4u�:=���-ȕx�f���L� TՒ<�n1rksWU���m�ZeA@�5�_-Ü��X��B1���%(��-��;b�8x"���d�:nr��ܪ�8Au�|8���ECc����s��v۶h� nm� f�q�mZ�m�g�e1�H&�V�ٮ�;��X�s{���r> 5u�lB���t�E�Ee]U`ڝ_���<�����M�j�Vr�����(KQ(:�	$�����K�����Sk}�K���Iw�0�.Ӻcm��IP}��$��퟇K�ߥ�����@+u�S{PCi�6��v���"#�3�U`4�̙���s`z�[��le:$
d�n�Jr�K����n�^�n5Z��v��y�l�ߗjɋ��p�๻� }�Ձ������܎s�Ȉ�_�]��4���&��ģ������r"=ϹȈ�r�>�&�0��l:������U �����J@���8��K��`=]��L�UX�y�}�T���(E �#��*�yo��~�Kss{��v׷h6ܨ6�ˮ�`ڝY��DG����6S�l����s�e�8�9H$������\v�j7DGG ���'cs7����\e�^�ȑ&:�	$�����/f� �fNr�;�d��=��ʐRq����J]No��s���~��Ϲ2k��2C���f}U\\����R��ƕ5�`��L�л�f/�ty���Ev��4)�����}ށ�<���}��n�NBD:.f��7�uaM��5u9���G�w]��4��9$J(�%$�@~M��#��	̈́)���X
5A���?�U�Ĺ��Y�Q�V#�1���юz��q�z΍��V��\�mZ�[� �����Iv�3uU�@�o0� ʔ������f;�\���X��� �*eǹ�7�w���{Tv������ i��@|�2����`}�V_dI��BI%����uW~���^{��c��"F�<ZQ3j��Q�T{�~���E��=�Kd"Rq&nN��&�%�fd�}�����y��0�z�r*�.�>3�pweK=�����8l�1�'����p��F�q�%�N; �fK
iw��`4�Ȍ�M����w]D�pOj�];��� |����`JO��)c���*���ʤn�-�RH��%������`JO�z""eKo���Vg��[IJ�		���
�Ut��5�
[}��aU��9��{�\ ���iB)9���&;�(�r���ڰ����`JO���G�r�7��_����#Rܣ�-�%��^�;mrMېs+���'6vMc�۶���3Odg�r����#�&��'���62�z�ܛd�&�GaP������v��ӟc�FJ�k[aw�3$vOGg��(�e��n[�vE�+;d�S>�:�v^څ�:��9�����b�vCK�����5��x!eLn�*y�X���z���Y\�Z�jݽm�o[�7�|�:�����vߟ��K{uċ<UЬ��[��p<���v�pc��q�g��c��voer�ճ���u=���u����`JO�Ȉ�6Vc�;�Y|i�&:��rK�77w��N���l7U\s� }���.��I��nN��͖yfc�?W8����?o�߻�
�Xl���i��j&�X).�f���`���N��~t:6����c��v��f�s~�������1����%�|�;�w-൚�oW-๗�x0l�ݶ�\�<d.Cj��F=b��+����8~e�����߿���`�:�6R]�""#$�uah?����G%��K��L��@r	�� ���  ;��s��ɪ}�֪�&�g�5��g���6(�������w]�;�d������N���l#������ܺ���:�ja |��GJ���3�[t�Ȕh����s{�f}���e`
Z}��U`{EpS�=�����n�w��{nLq�}۔�S	t�Fε�㶒݄m�]㻷T\�JN6�1�/�|����4Z�`����y�T�ĦI�M7Q�rXY�vp��.�����@>��`wG�C�m'r��Z�� |����a��Dq�|����U[��}��}��}���D�Q2�"�5-1QLg���ΐ&3a�l�i)�I�£���]I��rd��`Z:��9����o	:�˚�fm�� ���52�10D�ݔ�MK�<|Sf7!�m C������P@Ah��i���	�]�RC&,E�������F��\�:⚚ ��F��P:h���sG��X=
T�Q,#�s�����{���P�F/ IR�
�F��P� D����L��I�=��Wo+��ێ�$=�m����p17a�14�)�!��\(���,ݚ�j�TFaѣA�0��"0�h�hѯ����G��O�?��aT���`�lU�ꢒ�@�x�y�Uڏ��^@q�D��g~s\����u�3�B�q�ۉ9II.���W8r���~�e�v��Z�`������L�
D��';�>Y����R���(N�&�`����. +�ET�JX��E���m�eB���Ou<[��wY����[����9��Rr;
�v�{%�����:�3]��*Ц�F��r����]X4� �R}� ժ����eJ��D�D�G$�777� �3e�����`��Xz�]Q�)8�	&��@�>��`�d���,?��vy�"����!�CN���������!��Q5rX�UXn��i����`~�r9�n�z���T2z��{ ֺ�k��k����R�o�Z64)�ub{?�*.�x.�� /z��i���۞��U`w<E��"�8'# ���曽��P})>�Z��3uU�� q3ؚ���I�s�.���Z��x��!s�ـn�oz�@eJ{��R	���r�%��� Z'K$=֞aS1�G>]Nlg�3h��F����} �3e����G=�?}��/ݰ�]�?G�s�����۟�q�q�����T�
曞n��XE����:nk%ta�C��7m!k�m���1���
�eɶ�����v��R��k;=���U˔]���<p��&̎�w��rSr���Y� �܏�FwSWg��yq�.�&�R���u�ӜN�-<��vź��hŗ=rz�앂��j؝v����:|��5�>�R`4�f���ۊi^C�+����P5O{�����>{׻��۱��\s��i:�b�>��8w/\���}[X24�����B��z���{����������MEUU`~��� �S퀥j�b�K��Tl�JN5Bs��]�
V��#���:�=�?fz""91��rC��(�RT�4�����չ��;�Uc��{�ـ9Oݰ���`��Ok�TUD���p�Dp�?U��O0:�b�Ş�`{�X��F�NGNKu���DDDB��l+WlUp�¹��j!�dQ�
R*|EE����U�\\����.��v웣��wcd.���Eښ���o�����UX@�O:Ux�2�l)�E���՞����?4�-����#�n�(�Wq��&�`
u>�A�Pt�*��j�������0ӫ6����:�l�g���{UaJS���J��KĿy�0)�����9�3R��>��uF�D��T&������՞��-Uam<� Z�h�t��J�{�N�{�+Yι�aNx;lD8���Dv:��q��:9y�&� �%I#�IF�V{�b�Vm<�9)��`b;���#�HIJ�+��R<�e���oz/f�{��{�F$M�$q!8��y�މ�����.8?���c�|�e���~I�5!J(�$Rw~A�՛n�+Wl��i� �EC�:�Rr;{�w=����@���`s�\�Vf
��m�MS��sN'Z}����v��[�ݑ6���N����un^.��HI"�r�������[�ށ�ٮ�՞�g>����*%B���ƞa��$�)�l+Wb�1{%��Uq#�[��/�)8�$��z�~��j�"9�U��L� jQFԕ$��� Q8�<��c��Y^���u�z�����H=7�b���	�W0�n�����Z��)EZ�x�N�9��w�)��`9Z��&?���SPs��SwH����И9�m�O��ݦ{6�+[�}��a�#�k@ة�j��?f �S�D1j��A�� }��������B�QB8��J^����� Ū��y���Gb9΋�u���`&����`��
=�=���f�/n�F��H�9"S�-�*g��X	�y�	'V쾭]��<��:*1T�H�3w7� �͖����*�?�*9��{Î�+�ٓ����q[7B])@�Jv��Y�Z������:)��'L��7]�Y�]Q{=8�ݜ�v��2�pl=nۣ�m���3X��y�5A���VZ��0���@��L���r4���t�2;v�,�"��j����-GQ��xЦȦ��*�Pt.�hg�ĉ��T�6N��'Sfwn	��e��7N�8s��lJ��f�m&G4��1�G�����~{ߝk�ɼ!s�\�U,���;��F7;����ĺɞœ���<��אOUq�ȟ�I9$�$����r�R�v�岻V&�� ��8��Ԉ��H��a�Y�v��K7s{��l��*��3?/�(I"�U����zj�M��zdi��KO�@n���D��Ĕ��j�\+�~���S�l+Wl5)�V��냵D8��qIށ�ٮ����o�}�n���{t��|4�������"���ݳ�G�n&�p���v�.��FN�[6�{��;m�uڂ�T9 �#��=��;��`f�oz�͖۔�ҕ!�v� �uq�3���
9|��l��y����,Y�v}@𤰢�1T�I$�i������L�Z}��u`}�Ǧ�{7���0ݭo��� 8�g���|�#�O��UX�)� 5<G\Uv!�Dn;
5g�����
�9�_nl����@S�b6���#�v*���3[l�5��ˠ���C՘���.����jȔ뤔�K�FJ���Z���ۛ,����V/f�V{��э,�MĜ�$��o�{Ҫ�U@g�e��=��;��e��KR{Cs�M28���{�o�}������ ;d]h �0&����U�!� ؒ�bJ������?����B		T~�����:Ϣ9��}�]~u`n���T8�k�v���j���>�O��N��F ��]�����9"r'ۖ������r&"""!����S�n r�v���|yc�5(�EMB$�9H#���6���ƪ:䎋��\�skx���/l;�ݺ�QEUU`	�y�)��`9Z�Ȉ�9��K�>ݤj�SuMRT��z/c���纻e̘�U��6�3܎DL��Ə�HC"���u`~[��
;����r"""W�y�)��`dI�9&h*��������#�ͺ�-6�� 念���~Ca�� �E�"�3^���IkI�D�I��I�aF~���)>�V��$��6�$w��˲�A<�C�s8������"h�������'��M���Q')�9�R_@ř��r�v�1%W�DD �O0P*W�Tt�Wn �v�1%Vp��f���(���@���E.�� >mՀ�O0��R��L��]������Jq'"��[�����V�~��V����'�ȟ�u`/{�9����T�M��Y�����`Q�fK6�`̏�1K��B�TURI/�����U��fX�Y�5�I�YU�wٴoሚ۴C�Ԇj��8`wpPѰ4�!�i!�/Jo�v	�m�.��O"{;،=1� ��t����B�`iԸ�!�'�N@�Y�r,Z��8,�bP��SQ+fp�+Y���ec��f�h(gR�Á�FAI��)��,R �(
��(�	�)����Z=��C#0�H8�R�cT%;:��;W"��# �	�Ĥ�!η��`�%d��t�0�JQ��CF�FF���xO�n}��|��x��0On��X�[d���N����յ�m$7kp]r݁^��&9��r�PA5�3n�q�y]v�&�6j��(+k]!����2�j��ő�����+��l��v� m�+�Yt�[(7C��UP����)WV-ha�^ջԎ�p�]Nܻ��8�&[B�#n��7݅5���r�e�);m�2�'k�Y�h-Xp��m�㞽N�8�6�<�*��uܐ.��a݁tl�� !��t�+�m�vh�V��lf�.�3�ƒ#�X�5T�6���C�-)��c]zm>T��K������+��r�^3v��L;�m���Jq[m�!��3�Ju�(�z�P'/��Tm���XA`���*��ʅM�Ь�c/@��j���\: eZ�m��L�R�vxv��fՊD�UԦF<Qc�R�v^wh^�"�	�K�t��:Y��ŷ 'qy�x�Y�;"cl���ކ�r/,�&��.n�q�挮pU=h�@�O�h��
�>X�M��,v�f]�5�ƽ��id�,�'{]f���zw��ӌ�m���l�vW�F�:n-Wl�Yi�
��4�b�̅'d@��^��;4��%aԛA�΃�@ꪓ'��I�W'@�mk8�jm��l�ګmg1����j��r�A�vKEC=�y���U�1���zi���òMQ�d����nGv� �.�ޮ�j���a��ɲ�@Tc{�]�˝�nv&�n-��R�9��&	�ʻT���q���n+5k�U������h e�!�qZ�j/[VBx}����V�A�d�	-tP��ҵ!�m*�Ԥ��UV�UR�mN�+��Z���:y�e�S<j����s�rET���4.�: We�ـj���u�ή��`��L���zT5M����A'@q�1��8��Pn�*�U@Bed��WM#�݉5��)Vٷb��i`b���jU�M��h��@�mf�{J�c TTo�z����eW�:vP<���zCrTN"(����M���}wУ�?�{�������� ��ظJu�v-���7�m�?I����M��so9m�3�ewa���J\i�;�۱�[*ǌ�SB\ї��ڸ�i�sϒ�dL�/2�o˧�M��y��:�Z��<�ͳK�V0�Su�^�vll���9�9��+�7X5��i��b˵�/`z@pGj]�b�	�n��te5���=��+@��힧�Ss��gt�g[��|s<�۴����;�/|��w�w�ng*��b7��7j�8<�'9Ì?"sLs�&{Z՗�c�uJ��2JiF�� |������̖wsz���u{�}�\*;�3�ϫ񙽕���b���o�`&��Ko����\��IcI�D�I��MԖ��� �I��2�� �7V��3��P�L�);��\��U,{����nk���J�<ra���P
b�S5$j��ڮ�V��jUgfSi����`~yZ~����
��Q��BuP��h�n0�h���m�ծƱ<b��u�jݕ��f�]%EU=۫�|��p�`����N�}@��ޔ0e*���~��s�\�: U�?:6�ߟ�1F���x�>�2]��j�-j�"���nw�y�Y �j�jU`&�� {0�P�F2Jj6�5g��}�,<�^oz��`U��,��	JJvu� �7V��G!���|Tț�X~�v�Vצ��u�5�PrE*\R�=v;o=�m�άJ<ҦՉ��]��]��WI9��8�rt��w���`j�c{�}���3��R�"L�);�J]XV��-U`&���Ȕ��D�(jHTrKV{�wْ��_H� $��@2JQI@�4X�.�A�E3��|�G7k+Ӿ� �N�j L*J��T�T�.��ȅ3�n��y����~[���Ғ҈5J�B)%���� ԝXR]�Ԫ���=� 翧Hh�k�'&={n���s�(ҳ�m��㶢b�_9t�\-�ȩ.:��k�nH9�]�ԫ��#$��f yLx�RB)�)�ے�4��`�d�3ww�(fl�:��k�48(��� |���m��ț�X��ly�����n%$q(�3����IՀ1%����vb#�B��Dv��e��A����3���R(&I���6] �%��u*�m�F�㽋�7Gmj��(v�;�ޡvn�� OZR�ۈ�δ�`ўמ;l��#v�[���߱%��6R�������V5 '=*�*��9u}� �7W�Dď��� ~� �$�~����Q!L�� WH�������{ل��Y�s��r&|�u��ݖ߶��ŭ.EJ�N�=�L��V��� ϒ��"_��w��~0���H���#�X�˶��DD��� ��{0u:�?E�'���1�0�'���?��ֶ�͖�h�%18��D�e�f��֞N�]����P$^	��f�g��h�۸��z<��x�$xxNs�lsέ�o;���tpɳ>��ӱ�cu�Ok�c#�D��V�rkt��4m[�ۦ��8s�C����ڨ�"��9<l���n��}�/m�IƁ��� �6�7Tk`L6���4M�9�¯)ˈ�H�^��1��\�����jƚi���{����E��V���:��v6��
��=���;pt���y�;���?%���RN�������U��O0*S���]�7{33�TI�9I�,���@=���՞�`�d�=��)m�8���w���N����"$>MՁ�����4��DP9!M�,^����}�������95'V�����U5]���� kN�M��ԝX
w[�?Ẉ1�'J��IJ�J!D���ct��8���5��'h1��q��	s�������	�TQSUX���`)>�
w_yvI]�d�����.-b**K�	��,�w�G��G."#��9�zi�� ��>^}�o�1=j7I��Q��:��k� �J�"#�|��e'�K��2��#� �R�@>��`w���@���t��m��I$�"Q(��ģ��ϓy�s��#e'�g��`�U������c��z9�C[�9�W�Z�d	�!kur���s����s=1 gv�wf�ŗS3U����큓���3R�>�� � a�PP(jHA���{5��s�G2���ʻ��ߺ�+��ߵ��9��m[_�Q8��F�r�@=����;�{�_w����'}��#�Q�`��G66?M���?{�l���uP�2G$Ĩ������q$���ė�]�\��}�,sv�%ŬE@@)��`������`�U��ky�}����^uˮ��t�ܹ+q��D:^�gI*���rt��ۆ���S�@/.>���{������jd�j&�nK�ٮ�;��`w�n����`bՔ��iI�$Z��a��4PSK�߳KۿLmw�s�;�Fd���RG�T�>�m~�@�ٛ,�f� �%���iKx��Ҧg���Drb9�M���C�l5*���"���s�}�f�2 ex	BRB��XY�v�fK�;��� ԝX舎s��#���`��v=�������],3�ܝ�q�u�!�۝����t=z^�+�ʫn��wȜRG*5w-����X�30Rup}+_l��ޠ��R������z�͖�r�Հwْ��UPn�Ը�Ш�I$4���ӫ�� #��Ԫ��	��@i�CdD�&�:���,��; �J�ى����s��u:�>�쨝j�NBT��:�-��ݖ�7{�<�5�-�v�OW9\�޳i5RTt��Υ�r���J�u�-�/7#;5��ݬJ�vL]���	]3�e͝�)��ۣF��۵��\��@�sO=����2��R��
s�<ջ��n�Υ���]^q�A{Na{\���xm۲������1�����m+�z��+e��	t��˞e�a�#Kvq�s.'�`���t�s@lhY�Ȭ���qF&+�뻽��w�~߾��ڃ�ٳOZ��ǋ�s�������v�b��Y��|q�}����3�jT i�k��~������ �I���Z]�s��3�V��B�JJ�eJjN�
���`|�1�jU`k��g�#��L�����UQ�Uv�����`�U�#��DJ�~΁�w���i�"qI�]�} �7V��`��큒�큜DT6�2�J�RKۙ����Us��k���u�}�,���� J��DuDɹ�[�ld6\m�.�������$Ҟs�\4�J��⍪q���w��͖KK���X�y��!������vԵ��ė۶g���*���mA��|(| xyY�}`{W�`jN��DG92�{��{	�SQF�ӏ��ߥ��������Z�o�t���=�X��&�NGnKG9�'��:�2Z]��9?&做�R��"G)���s���͖��]�Ԫ�֓�������⧫��n�������{v��jx�V�杸�����T ��E8%$*9%�չ��3R�ZO0Ru`}�8���j���r����n�8��y���廮�s�
���0�5N�1T�E$�7u<͙	IՕ7�G�j�*�$��/hJ��hx��C�fČѳF��t.��O˴,�Wo#�� �hxkj����%q]�+�]��t�it�D��$�ִ��b��i��c�&��p�p �f�{�w{ҧh��8*�� }���J��xK�TqM����8��9��s�>���G3�K_v�=�����kb�F��Q�ހ{3e����`�d��9G������+v�q4�##nK"^_n� ���t����X�e��U����T�T��"JC��r��V��mr4up��kg��s��}������t��{=�� k������ 5'^���r�y~����$�"MD܊$ܖ�dg�$~�g��l3R���#���VʊD鉒�'z�͖�u��G Ԫ�Ԟ`�L����L�Qڪ��s�+���u2&���Kف�O�~�9�f��r��������H�k�]���u`~�Go��o�`l��`w�K.��@D(r*j!5�$�d�o=v�q�v(ǎ�_Y��ݲ��6��=X��Sګ 7Ry���e�����U��n�ŭ�R�J����fl��£� ���l��U�n����!��*H&�Ԥ�q�[���̖�=���@�fk�
�+����Mʦ��R>��p�7V�O0��l;3�o��i%�����ě����7�(?W+�ȅ�~�p>��as9�U`~���Ds�R*>�"{��HAxp 6��M��SB�
Vc��?��=+��]�.��÷\Z5;�:'���ugm��vz]�9�Kn6�=u�1k<��u$�'K�'e�Г8�*�\�����P��˜��ͦ�iz���판cn�/]��h�rʂ�Mt�F�p���y��pO�����̝s��Wd�\�{v��%�]d	��;#r���������J����nݲi��=�[{cGlUn�+.��r�Q�����w�� �
ȸ]��1�Dӎ7.�DFgvgkn�׷o!��l��N���GY�u��v�m�y�������_���[���fK�*��������j�
q5$!$v��l3���I�������[�RG"r%ۖ���e��fozs�U\���k�<�u�A�Pf�:�QRQSګ�"uC~� R��`l�o�߳%���o�[ ��I�Iށ����9�s��۫ ϒ�$�F l˗������s�{h�n�(�s�Βr�;'1e�{u�Yp��Q��P��Y�۫ ϒ�$�{���)Oݰ��W��7I�Ƈ����+I�v_���_$F%Z 
	��	aCJdDp��>Ȉ���	i�0�7� i�>�I,FH��Gn)`}��]�
R}��9�{�=�U�}�Հ��[�ahi2s�˜��Ue<������3��ӭ��x�H�3UEUۀ�������*�3Ry�y{5�R3y����*Q)�$�Ou�i�v����Lm�ծ��8�����n��������	#�9ܗ:��e������O��r9���V�����b��D�j��{3�ȉ�J~�y��`�����+��y��ű��Q�ށ�{���U��}�_���A]���\����X����T���#��Nj$��k�-�V|�X	$� i� �+Ե�i'87D-�'@77e�G"#�Rw�5���n��N���;��"k�����=ty�u�'���d�$�L�D�[\e{`ƫK�0-~l4߳ k�̀4�XԪ�H�\�`�i����z��Nꫜ�k6Ӽ m:����`�K���Of����6 �u �*��� k��$�}�z}L�\��y�d�_�P:���U���f
In�͇�|�9���q2dt!YL@�FHA�
�"�h�����|���e���R!�P!���3?w�UUV����p ����VO�Q'�I���}$��:�ɺv��!�I��s�Vp���z{�ڜ��v
��\��;l��#�P�_�n=�`	7V �*�>�$�2d����LM�jRt��;��:�^̖ٙ���u� �k�l�49���-�'@N��O0�r99�<��M�d}��������HGnK>��ހ�[� i����MՀ��9~�����vzw�v� k�����Dy�Հ?�ʽ��u�_ó��f�`L��V��AϏ{���m�Y���*Y��^�&Rkם����	d'K��T�[kK�V�=n�l6�s��h#���he�ӓN�=\]2pvy۶��h�N���R�5�V�E�4]�6V��@4vm��6��y��;n��u�p��I��j�gCg�x���n�!|�l�#l�M�軛'hr�v������c��#f�m��ۆ�#Z1��V�ڹ.���5��g�o[w[������hF���'~v�ՓP�2;�d�v�g���%8qѽiN�ck�;�j����v�\��+n�s٪���M�4�XԪ�[��a �wU������H�NEے�@77e�fV�y�=�s`[�T�Dw�"PJ9.��{7��w]�F�vX����t[*:�N��N���l�u`�U�#��y�g��S����RH�>J��� ��%���oz�{�����9�1H�$�:ή����ӷl���pt��#���=ti���|�J������mI:���,��{�<�u�*���vX�нK!��$ܖ����+���\�?%g�;��D������2X��kؕ)*E�U��o� ���� n�V�S��)�D�iI'$��ʤ�?~�`�V�W�}�N�y`k��#�9nK� �ݖ>�f����w]�n{e���K�Ƹ�*u���R�H����zM��@��q�7$��8-�넹��m�~{��ݷ�Zc�qR�"rX���z��>Hǻ>��=���o�Ϗ�b"IT��� R���U`y*��y�9�W �.��D6�H9v���e^w���>�FFR!1Y%X �G�@<D��@m����<����{+խ�N���D+jJ��Ձ����?.����#��r!��Xxh�-�NA�p�;��f��>���*w�h�7�i�{�9<=����P�]�X�8��]�q�.�ՠ��7�mչU��y5bާQe>>$�->����ߕ"�9-O0���'RB
G`Q�͖UUUr��oʑ`}����O���vj��{U9uWX�L�1jy�l��`V�2�����#BR�ÕU�s�d-O0��ljua�?Dr">��G#�Q�H�Fk���_w��h�5�FhĪR�N�-�w�l���d�Çsٽ��5�{TS%6Jr�u˚���8�f��c;t�u�-q������xO�8�q��$j��R8�<�d�,}��<�#������CQ����c���B�o�uXN�`b�� �m��[,�2BB6��,�f��l��a��s� �u`n�E���멚���Ȥ�Rw�yn���`{�0�;��ށ�Eb[t�II'�$�X��`bI���������G�j�*�$�J=\���D#�$[pA�A)�B�i�P/��������.	xx�o��w%!�p56 b���hD�'�)�0�����c$\���h�L���;�0v�k ���4l����j��� ��Nv;�X�i �f^��i�-Z�8����pC�ڀm�T)�8#�ż��u��z�f�f��2��ߚ��=���2TuZ�����B����i�b�4�\�i�����&{e�R�5V��I�]�*�6�X���%�-�]������ʾ݋8�
�N��L\p��nql��6��i��
5ۃ���a���ζ��[��s��j�2��tH�q֚i����;�7+�-On]��mz쵶Ԛ��+a�K�=��Cq�ez�T���ӰqnH�\H]�-����+M8�;t�h�I�
5�o���|�܅� p&ų�IK֫v5�ۀ82k]�ֺ��Ҙ�۬�m��a��Z֋Y�F�=�O�^�9�te��ѕ�;�d/:g�:Jr�=ۀ��غݵ���g.*��)�'�t�Q��1щqa��bZ�I)ʴF	��F�U8�!���8�zpRv���vr؍)!�( �	M'i��r�I�#�h}�f�C�ΈD���BѮ��x9�g��U�W������� Dp���l��ۄ5!����v�vP�jU �=�W�n!�%��q��pc
��3��дnw,�2����rv��6xˬM힠�)!�Ր��P��\{['G9�7n�-/=$��N�ɖ-��x(9�������^���;$�I�l���UQ֣$�H V!6|�u.���kj���/b�C�PX�"�:��sp�d��V�Rړ!!��.1���A���cp��>��{��Y�x�q��'�v�9x7�%q��^�\�g���.�V'DE���i�)ݸj���k�`�s[ut�}��� ��'���{9��`��$n����Xu���I% ʒץ�an����-�e�m[  �[��V�z+�͛��],�����J�ݍ7+�U�s�>�t����5DN�q��V�ɲO0R=n6���b�K��齮L���1�3��pWK����@�� q[ ���tջj�2Y� Xe6-Mym\��l0R��Y�0��I�s.v�-e��ݱT��p��~G״v"�w��"&
� M'�$���ר�`���]"/��DL<���?��&3i�)�#�Xiy�v��,��]�^���tbӮ�W\l�=�� bʘ�N&�U�F�&�O��VW�r���`8��o�� �Nh��9
�k���f�%�"�a�{weݸ�Ֆ�m̵��8v(5���Ѳ�9��� q5�+����eٹ�ޓ��yK���bu֛9iV\�aY��O�]Փ\��o	��O!�"�՘����w{��~�ߜ��'<~vg����>�}��
���x�n�'>}v�@:��r��������pv���p�4}}�����_�O0��l$��Y@�K����ns3{��ܮu�'��l�X��n"#�s�Ȑ����=�&J�(;�U��{ݰ��=�s���N�`|��`=�@�w�RWN�b�j��p �:�6uJ,Z�`�#�[����=l�l�M�
ڒtͦX���?}�
}�w܈���N�jvlIn��E�c�u��we9ۂ� ��f��.C���m݌�t�ե-`c ���0��������T�k^ĩ8)�I��B/=�w�+�W�Tp�_�G���f��o�u���r���?����UW)#4+R�t2�����g���T�=3�o3 k��l�nV�iH�RC�%΁\�fl���{7��w]�g�e��e�,n�"Q%!]��ũ����-N��H�=Uʭ�n��9���4�H���j�)����6�7I=�^{:;c�J��qe8E�b(:����~��`S��U���｛ހn.ָ�Ƣ�.� �ڿr�m�2�OW� ��ŀG9��=l���)��Jڒt͚X�g�u¾B��A�1L1h��q�9\�R_�Oŀ~��,�eA�w�E=���#��A�O�`ޯz&M��,͚X��=�T����
L�5�e��G#���VN�`b���;�8����(���*�D�Ƅ
{�q�cbk���t���vï�q�}��iJ���� i��7U"�ũ���,��7i4�N)!ے�@�٥��G�?f ���`@�:�>J*:�bh���A]��ũ��;�Ð	�5`{�0�7ڵ��t�QTE
����U���{��0��uR,?EsTs��r9a($��%=  �@ܮUb_}�� ���Ҝj7Mҥ(rE`S�#uR,Z�`@k���dP���x��x`l��խ��h87�:..�Q��Oc:ݞ/K{+v���6~�#r�8>&����}�*O0}nlju`}�I,�)#d�6A'�����r����zl��L�T���l멘�*���
N�k��`��g�UUy�{4�>������Z��QR'�-N��V��<�5���>PA�6��N)!ے�@37e�s�����}�r���~�*��� va��?Y�������}t�y�ў#�G�{N�.J����y�[��N��3�9S�L��$��p�۶ݲ� l���®#���f�5խ�xC����Jt��nŠ���C)�b���`�[�\�a5][x:j��rs\�'n����o������G>��x葻]�kX����@/\�����)m�Y�_b����\n�x�e��^ݤ�6j�Oh�̳������uT���-.�Q�(r*Q!5�x;X.�{Tte�1��[`f��y�ݲ����-TT�B)%����~;�=�uX}�!U�%�n�K�����,�˱T��	�U}�/wޛ��Հn�V-O0*�|����IFP�RrE`��`�U`b�� �����h랸���;]&nf��&��ũ���͇� �I�����4����(F�#M�`w=���z8�^��O�`�U��{�w����b�+�n�����9nyq�s]c:s�7!�7Z,��g#��i�b�Qe>>$�Wϭ̀-N�u*�1jy�2�]�n�Ē�o�?b�?E
�����G9���䜈��W���?~�e���r���(����JD��.tw��`b�� �m���V�@WISخ�J"!�Õ��;��	n��f� ��%���Z��`����$�@�������>Ԫ�ũ��'5t�`�ح\b����;(;���Zά�[�<Eǲ�Zsbe.&���IFRQ
9�g�e�}�V��[��`���-\L��ӌJҒt3^�sٽ�݆� �f��Iy�qB��$ܖ}�ߺ�>��g/��@�)!т��?��	�0a�0R(R�`��� !�85��_�:�"����`{�t{�JI�H�'zr�7f� �:�5*E��$� P��;�&�DmHD�,���`{2a`w���@Ż�Xs��i��QR�$n�䦩�m=uیm��tu���g��{2����ջ+��z�"�R�JD�r\��4�;�b��-�����,���Db��B���Ev�>Kـl��`�Ձ��E����=L)D�B����@���`�l�9\�}�X�3{�
�*�oZ�����%��=��`}�X�3{��A�)�,c1Frs _+��+���[�~���N���v�����$� �M��6u`s�ʛ�jt���dj(�D��9J�R�u��۶�o2��fM��q�����0������K�$NIPj�,f���,�v�͖�Ʌ���bU*9"�I��@���`	'Vک(I�zdP��z�#�DmHA��ݟ��d�ª���?w�{�>�(�n�ґ8��l�5:e����WS��=)�dXT��H�-N�(�,���ކ�ٷ6��,�H�2?C��#��G�i���_�Wz�&��GC%������V�};4� �A/6��sۛV���*�[S���K��Q��=��q�ج��ݲ�F뛦s�3�ٶI��RN1}���g`��?��σ��v>����Zp�nx��PV8Sq6�:t�ǂ�#�#�� �e,��ݧHK�qϷC�N��K���G���T#b'WsQD�;s��Iz�
�"�c������m�-
=9Ր�/���ǻ���A�
(�}�7V6�9�D��.�n�nۗݹܥq�Wp���^��L�x��=��HR���������f�X�L,�3{���7�F�ڦ��+>K�S����&O��Ys?CoفR�77�DDp��z�{Q:Lj$��ٳK�fozP{j�=�۫�i$�eEN�	�Qa�Ds������6�X5���`g٣ؕJ�I$�Rw�f<s`�s����X�"�ϒy�dzw���r~�{uŨz�/Ѭ�c]�x]�ȝ��q�ڹε1�3����ܡպ�;JV��|n�� ��<X��]����Xez��MH�R@Q��@�6i�U{��  z{ U<<���߾몽Ǻ�{6����\�s���iR#5�NS]*���߳ �Jl��,�0�6��KS�'�HR����Y���;�)'�OـS����]�WlR	�q�K�߱�IEݚ�%��w�
3j�>FVkek�R ����Y�=ۘ��1�m���G��v�#ϨŶ�����0��G)A�h����n�,�3{�3j�>�mՁ�4�3!$M�@M�`gڜ�vdr�큺���>n�q���ĪS�G!$B��f�>Iy;�>�֭��iv��I$�!(� �@R{�t�$�Ap��65Քr�*�� �����H��"*&�b�jH��c�)�O{p����68QY��"^�tvo>њ!�=a��l��䔓f8Kw�4E4�$��jʍX]�x�QD��������C`QD@Vda���4�T��3rr*(��0�v��l#Xj¨	�,��C}q���1�9�Na�$����!PZM��[��h"-jצ��U�[�dG�͡jM��;�f��oF��f�ѱ��v�O��h`L>×�F�BP�w8�a��L� �:tj�2@�b��d���,0c��К����5���a��� ��1	���6�:Tty@:�T}T�� � �[G	��1��u�v'	�כ��_w�ߺ�|���Z�u(��9��/f��Xn�,�����/�\�����FW��MH��J�UY|�2���Ds>�����`}��XE��b�Y(�"!
(���^���-�.�]�<��g���Ǘ�n\e�<[h�US�,�S�JO�ڝǢ2C�������蔟!JRr.�13i��w%J>��=�HyO=��j6F�)Dn;5,�����d�:��e��@�5��p�jo`��c�%M�����jy�������������\�(�Z

*�!����"f fbD�_��Nr����\H�i$y��b��	�����2 �G��`}��Xĭ�?˕��c���iks�<��|�8�$g7]��gi�g����Nl���Y��;�
�������`}��nH|��`}���x�D�"�DmHBH���ug9�[H�>�S���]�G"#�ɓȂm~E5"�I��t~���>�ٵޞ��<�f��u`fz��t�A@�.�a������ �e����Ň�9��v��?o�K�tJN�)
�''z����Ł�R,���O�G=|��w~'���}���:�m\%�Ȧ�3�Yy�˷WD��"���Ԫ5O:گm��Y�E˻98�$D�n�cM�ûs���BP�&�^M@ֱc-<V�g���d���b���.�!-�����;��m�]��Ѹ�c��uUϷ��"��8��n�F�D�Ҽk�Fcglgl�T㭃���`-�&�����h����14n�΍������U��6�n�i�����z�|���9�Eob��Ugl���1���ϧ�ݢW�n��e�Ny<�������|�O���2bT�wW�˫��Y��5� Ӥ�R�w]�٥�������}�3[��7{32)TvJ��m�X��}�s�-{�^/��?0�>ݚX�4{�(�I"�RRw�d��`}��Y���U�}����T�{KTU(��9���n��L,��oz,�v�Ue���Ohq�T�Ln:;35om��|v*�<��� :u�q����۷i�8ԑ�H%'k�}�4�+ｚ��1fk�=��Ձ��B��:p �I���~{�]BQ�DG���S� w�S����q`bT��?/z'�Ш;Ĥ*D��|�����۷Vs&~K���ހW�\����IDSD����۷%H�3�O0)>�k�޺;=���������,�S�JO��ͺV��S)���P�!%>϶�d9Cp������A����cnw_��$���w��%��$�P�X�o��^�v�ͺ���a`f�b\��9"�!Iހ�S���q`b�E��jy�(��Z��DmHBH���u`w=0��V�`��S�`�1��i�	�{�^:������7(�b��I��t�)�}�� �S���q`-ؒivc��
&����X�����>������酁g�~�q��#i�9y�s�M��x1��2F��W<u��j�q���r>!�P��$i���j��`}�ݺ�;��X}����\��uJS%(�v����ɋi�O0:�l����t��S�n��ۓK��ٽ���j���g��V�i%F<����*tX�����O���Ň���\�r9c%R�x>"'�޳��ܫ��bUR'!$��5-Y����u`w=0�>�ٽ���)�hڎ:���ĵܣq�>��,� ���(Ch�oL���9P�8��DmHBH���u`w=0�>�ٽ��6;�QFeLR7�)���>j�d�jy�)��`}��_�s)픩Ԩ(D�`{3w�L~�}ٹu`}��X��KS	C�n:����0:�l�w�i۩� }��٭FҔĉJ'��n�X�oەw���U{�{��ʿ��WX!XIYE��A?���֭k����f$��0�+d��b���Ϸ�:{i`���v��8����i�+c�W=4o2�܆��g��,n��v��֓<�%��{SW[S�	�ڜO��v���Y������[t�]���9e3D{e�3�9��t��rvx���q��9�����i3�q�j���4mOGlg�.sX��O0���K��Lӝ,0V�I�=�׎&��b�gP&����Z޿�D%�&Ο;h��a������}���;f����F'���$@�S�S���:�w�p;��ݾ����k�|-��n����� S����7q`}���<��$�P�����ޤ�^�vٻu`w=0� �j�I�J��D�UTUx���`|����s�ɟ��X�����(R�(�QRRG`}��-�XjO0:�l� Jґ�$��t�&�`}���@���f��6�����s�a�o`� �(r*(�	�6,�Ǳ`�8������z�f���m��t�䎥HP$�à{3w�b�on �7q�r9��	j�`y��>�`�;�{ֵ���^�}�C������#Ӽ�}��=q`}��`}�ـ9侭j:jR)DR;�ݺ����{7� �ۮ�7=F��i6�O���Z�Xn���o��rv�Ζɤ�yI5Bp�
B�����@���e��n�X��sv�)�I-qD�0moPu�X�vW8���6��9q�X-mm�]k�N.�D���D�9Iށ�ۮ��7n��>�L,ff��g��J��R�ڐ�Oj��w۴�wS�o[�좌�6���JJJ�tnM,{ٹ���Dd�B�"#y�Q�����{^���hsP�B'�;���{~�-�s`|۸�>[H���;Pw�Ҋ��G;�3�ugP{f�Xg������H��&��"7JR���չ�N6�l�R�MF���I��wϨ�>O�w|����]���{�۫�������ށ�ۮ�7=Eֲ9��R�n�kT����o�B����W���7qpkI*1�$0Rr��>��{�1{u����K���Ձ�ɥ�����J�q��Pv�0=�9Ș��>�{� k��,�׷+?��$C�½�����U]�|Y���%	�$Q�`Wۻu`}��X��{�1{u��[U�֕m N'j����=i�ݺ�F��<\����hԡ>3�۵n��Z�
QG	%(�k�#ۓK���~�/n��UU���X��1�܍�J��T���g��DLD����}��`}��^�q#���K�(|JB��G;�5g����`|��`j�� #�<��}�$�ҥ(�Ga\��n�Xg���oz,ou�3=Ekz��T�D�рkT�}�F����zh�H�������� ���QTW�����G��W�|޹s{� �JR)#"Ѕ(��S%Z@
UD�F�P(iUJD��J XY�J�&B�iB�E�R�DZ)V ZZE�F�V�A(XU%ThE
A�A)@� �QB�T�A��%Q�P�
F� ��h��� �
R)I�d"R�@Ќ�@�P�H�҃H�* ҪR��*f�h60��(4��P�(�!BH
Ш̊�JT��rQr�� ����Z��Q�Z�
�h�JQj�%URaF�QZE
A$QH�A�T
iR����ZE�Z" Z

EV�JQB��W U��QF�AJPD�B���B�
T
A@��
�F �8��a���h�
�����������������������T�o�/��A�#��A�S�@c�1A��������P��q������������������/�QA�����Q����'������ U��H 
�������4�?���}P�������� �H�� *�������?�q4�s�ǣ����AB���?���I@��ID�Q�@�%�FI �Q�HQ!VI	Q d�H!D�Q%�`�"DH�R��`T`��	I�"� �
Th� iB�)$QI�&�P��
Z��)	%��b� ���B�(	�!���V�e	��BP� d��	U� �`I �%eI	BB���BBI�%(	B�)B�(A"P�	B@��$BDO�pC F�@�%Q� P�Bd	@�!�%�"P��
D"�B!�$F@�	BD%��!XBd	��"E�@�BB	a I	B�$F��F��V�XB $(R�%a%%	�a�Q�e$�A�� aP�!V� � Q! P�E% ` E�a �%�%P�Q��
��h	Q�%R�R� X Q��UP I@FQ�%DBE�@ YEF`YP�`RA�	BHVQ�%�B�deQ�YF$! `X@�TdY @�a	BU�Q�F X@aQ!X��!	�	F�$ �!�dXB% �	�aQ��QB�	 �`R�aFP�		FHF`B �dH@��i	H@��@�&B	�%R�$%@�edB��	U�	HF�aTeDR�$D�	Q�	�	 F��h�I@�BaG?�m�?��7��EEiB�'��y��O�<N�8�����W������?��i�������S�� 
���������7�C�U���
����O=�_� U�����j 
��Xh���sO:�@���r
���q������?��/���U�?���������*����M���8 ��?� ��S�B��O�Ξ��������:�ao������8�^ �*�:*?���d��f�h�:�Ϗ��}�u�� �*������QC�����｀�*����a����9����?����
�2��S4��	������9�>��� �P�J*!"�� *�T $����I iTQR W��(���� P   @  R�P             @  *� �   aQEEQUB�����T�����Jwk�z��)T<,z�uq�}�D������輀��u����� j�h�ﾸ�\�#��[Շ{�� �z��j�RAΩc{��^cvk�C�Ͼ}ʟ ���"�@�UB���H��ȥ������a)E4���%)J;�R������Z�(�@ Z!� @
Q�  @ D :$P��@�@�J �JP4P`�=좀BR�H�(����  TR(�� I�Y
I`iOLE{�ϳ���}����ި�ݻ�U�oK�޷J����+ {�\O��w�u�j�7S�}��ۇ�(�{�k���_O�WC�1|��r��<FO]�x�{������}o�����>>%T����U($�B�QD���b�l\Z|�s���޼�pUU{�,��/��>�>�ۼǥw 7	Y>�3_x �^6.�}�Ε{��F��6ﻓ����x�/3��{�D��<V&��|�x�}�}n�� xz�JU*B��D��/<K����Wcrjr��9��'־�S�=z^6�{��5޷�=w�G�π��b�7� ����xOYV�UU.OvCK=Ο}��j�� �o��w}�#v��'��   5?HT��T��!����5�%T�@h2d1Ǫ�E=OI   D�*���*��db41?�%�)J� h ���ʔ���A�"w���������������pΏs��u��A^����UҠ�*�������AX
��PT�"��>����I���1���k�p��<\Hэ6�i$T�j6 ��HB�.BIB�!��#�%�S�0p�L�fs�	��IC�R9"1D�p	(~�8b?��PbD��R@�56�$�;�6m��Ed+I!$r>W?0��OF�"B	�ԃX:�B�E5���%>o�G��ӫ�"�
��<�j��P�*�ŗ��\�,�$��	�U���j3O�,J�ʕB��1%$5ٵ�fn29y��*E�Da.����%!B$�Jd*E� d�0�a�j.�Ĵ�2"�Q��U
q��Q-9��~�F��/�׌l��Q�~�5�[�0��!j�4o�R�h�A�%0�0��\�ٌp٦��Tڀ��dD�Hb�l��R��uT(�cp��;Y3AB�s�V4/b�7	�����4� ���$B-I����~��\��l��?'H�'-d�1H�bivg&�VYbE��9�ֱ�
kAS�� �����1�
�����E���D��w�\��H�q�m���J i��y�L˿�O���0���77�HK���14�"�j��6�2,���;s׾{��=����>�Ϸ)n&�L$����,��yq�D�S�X��
ז!,2e�KT����[!$�046�F0�fWA,�i`0�ٝ��i��@���!��"Ę��MM̯+J���Ц�.�a�'�;g�`F������ٯĽ�5��lt�$(@�0 `��>˽�hc����CJ$�~u6��sy>�DO���)6_ۆ��c�F�!p�������*��=�ȫ�#96��{�%D��ū�b8�;
SclT��Y;��J)rI)PY-	�^dM1@kz%i�����X]�(�F!��
�(F��i�XV]O�I�sH��v�"Ɵ��f@�P�n�k�
|0'd%�)T��0�U;�vj��[U4L�L*BN�M8�{u�JLF�%bB���dM4E'T�]<5��ʻ%G�%��{��)���M�wR"|�'�ע���/�L嫒B�=s�P�p̒�d01�X��� �kX֬-)J��X�$%`e����-�1��w��.c��� ���b�Ń%A�F �� @����L��d�)�6H� �`Ƙ�D���"C)�H:�>�	�������?�ٽ7M.��!i&�3[�&�ԐӄBƄ)�.���Z��+����UE\(B�j�LqLKSM�ƏfuVm��<IJB�֓���)����R�+M}�Hu�
u4�b@`��5�to���d
��"�.SU�	oj�ۗ��{��T�k�
M����B�ZH'��G��	K�A��dvdn$8H��P���LM#$���FH��5H���B�������FIE�!\�/Y:�q����ϐ-�&s3�υ�~�`A��ŅX~���]�"4�(Sib ��U������zqFCjM�lT�Jdv��4o���9�+�S
�I�]Qb���1+��8&�vO]��k�}!�?2@� �GI �̮�$d�jQ�g6�&�.��K/
P��]ϣ>�a"XY�+��3��H��|X�'�2l�Դ��O�đJ?%�v���&�S4fȔ�8��l�e!LbCI�g?a��H��C��'��1(a�g�@�c�i�?��;vp�HP�7��ae.�%���Ww4K��i�!HS0!RC�
�"��5j����&�"`�B+��`�)����Al ,FU�W	�u{M�!(�QW>�D!E�l���Z�B������?r�PY�k���
�
��c��E�B��џas��8IO���\h@�,	8���R2eЇe�-��BLP�!
9��j F&���?$
�)�&��Rm*#y��I
(��W����JCI ���
䁠�CO�a	I�J8��6O��6�	r%�p�)�v�M� B�	"DM$.�� �	s\�!��~�����͛atoI��$*�9����ƠF��.���6����`|O�\t���(f�����1��
��*AǿHl�	��a��#B��jS5
c�m�9�I�%$r0 �6B!ǐ�o�pu��1c��S�]t���n��n�rB�h��UV�yfZ�X�T�L�j�1Yu��5�Zj�X�Ӈ:�L5�H�v�~�9����m�0�k����J�rd�&��Ƅ�s�R�����h��TD�t��Iq]����X���7 #~��.�;Yx��$i�0��1�r�laXԁ�r��\ՅP�k	���g�n&���ڲ���2���?����k&R5L�5Ϫ�ǥ���	G�����_	3N���"IXBXd �p`�`�� c�O���bi�B�Wr7�$�)0i �ĸ��s�����n�_�[���{ϻ�}�'�=���ݎN��<=��'a;=n����'c�y�ۏw�wq��k�1�{�:�nɑ!.$���l�{�T�jF��RS4��KM����
7_?�l?!�ጃ.aH1B-�\�
e	�ԅd�;��0����q:�zXB7���@h�X�a��5]���,U�x�=��F��T*��K�.��{����H׊��G9|�=c��ni4l�0�O�'���?w�>��[Ԧ�m���B�&�g9���V#v����X�4�GF͟��HS�������a��`5�y��4;�����qM�:+�`F	� S5���s�&�&�5��v�mrU(�D�esn�n��j��m�0,*+��k�i
E�$�³+e#B[���`�4�axoZԲ0ه:Wf��M�!Z誟A�y+��~b�P��"���M�m	�F�*��>T�#��2L\M;����6�D�M���� AJ	��
�I��L�����=t0�@���&a�0����R��FY �����	a� ��ܿ�$�2A���Kahă!!�"8�?>v��~~yrߢ��&����uap$��4X��8jĒbd+!���6Z�����7���Iݏ���n��Ǔ��Em�|��<�x����{������{wV��m�tP����!(���!�W@F"�"�c?$Dk���1+M~�aSfR.Q��q.2�Ʊ�*@���.�h!`��"B"~	_۽�{4�i��8Y��j|O���A� "0�/	�WT��sG>�k�R����WN�q @�$����L�\a�d
C��s{f���$V�٨���_��F�bDj�6f�������w�P��V�B	��p�&�6Ư?	�2�K"�َ�~����U[�!��8�9�a�I���f��Jf��@���M� $%2�(�{_��0���KBP�a��)"Y@�R,B8�La`B#��*@`ēZ����77����J�D-�r��G���^��;K��T��)��XSGnk{	��t8�㠅��0�߭�ngə�d��.���%�h&�1I�eLi!���HnX�u%Z�DNZD��
��!pֈTČ�+�4�P�MS�T�S��Z{�5�G��ў3�w0�3�q7�dǠ�9�J�KCCr E"�D�aV!@(�q%��!�S��aRT��D����1�$"6!t_ߍ�'��
@�������vT�IH@˩+`a�:6�@�?ۢa,���� \��:�\�>J��5�BA�a@��(�*V4�8P���)R�RP���"�H�BW_����0�H&F�(�(@���+��djĒI��Ē������[��ǞJVSA.Jb��j\%�[
�����h#m��    p   	�  �  �       �`  N�� $�m�      �h�` �`         �6�   $    h H        p6�     Z�[:7"�Km��a�Y�^K`���`v�Lm&�$H��֐�f$Im�ۮJ����}�i6�f�p�I$���t�e� -�!�lH ��` �b۲еnͤ��ܖ�x �9m^�f�H6�vۜm�RiM�x�j����	�0sm����Ir���m�����m�6�ճ�m���$��r	'J  #*�2��*���e<�
ҭ�9���eRڳL��I���C6�s�l�,6�md��i0��Ul��R��ʫ�h]6$�M�SV��X�Y,��b�m��/^���3�y=e��沌����ۉ��e�o=V8瞜֭�n0������E�O=��E�Q��C��xm�K%�6��l�G�D�2B:���YZ͝�-�.������\Ֆ69�ہ�P%��������]�/����Ω
W�����i;vid�I���4����-�芃`L�3��Y�ͻ}��~��]j��(d�t0Ē�w6u��B�cZ�k���m豥�#6rD�E��I�U�5t�\�"m��{]t�;H�b@m�^��m�#��V�kqa�KH#e���en�&��+[�mF�-Q��^�ݶ#��V�:$^'v����2�5d��va�ո)�t�3m�Im �`qm2tZ m��9�h  m�khj��ko`  [����;b��7k&I !m'B� ��#��W#������\ʽjt鹤[NH��kl��i3mm����u�8jCi;f���S��8�L�1�ڰGYV��Hl�96��h���,k�1���/R@ ��6�$p[A��k���8v��g�� 	��sf��u6���4[�hxl�m��릶��ͳn���ݵ��Mz���@�� @@�>6��-n i0E����ln�I�  t%� m�#m��!t���@�v�jM���m�r�B@ �`�ճ���� 6[Mo;/Q�lh-��ˋd�k��Y1�mi��l�	,��Y@�`[R  m[@��qm�`  H���:� m�H�v�km��ؗ8���A۞��d�Ե�D��-�kdd�&�R�nj� m�Է[�'����CZ헪@��I�6� 	 	h����-��I��kM���p6ݲ-��l��Ѷ�$��0z�m��۱�`  \��6�O�O������%H��['] 6����.�k-�4U��A��.��6�s�q�7m�,0�l��- t�;k��ZM9����F�14�j-ڹ�� �9mI!e�*�-��v�IɌ5Nԯ�K��rA�L��2�䜷��I�g]Wn��v��D��gQgMѪ�]�Y�����KX�h��/i2u�4t�M�h�m�Ûm�v�]-�M&  ���Hu�[m�� N�rY@�^�հ[Ku�� f�Z��n t�  Znm����ŷnu��m��h��l	�zۻn85Mm��F�IŦ�6� m� 	 ���l8��P � 6�oKv ��&�EH[Kd���.��d���m�)4�m'd ��Z8 �hڐC�۰p��5�a�� ��l m�5��f�Hc�Im�v	�ܶ�ͫd����6��H�`�{�[v�  ��k�@�M͸�q[nql�R�©�睅����kn�� ��>�[�d���$�Ɓ:�e@���b�X[e� ���Kn�	gP$�N��l-��6F�K���MC�m����{{bY�4R���v���U�x���:m�������W��p��w6��j��]�0c8f�0n��jB.�u� �j̲5��  k�s�����x ���}�P�`�ִƐm�	m�J���Kh �  �}~��ۦ�L[xn�8	d�m�    p�d���J��A{M�ku��m��mHG;mmͶ -� ۶m�`��l��q���Ci$C �l z�	 ��  [.��l-�I6�  $m�l�gj���� 6�`�߾�m p[Im�  n�d�!�ٶn��qoP zٵ�  �rA�m�m����m7m&�b[[ie�>�גּ��&�8���h6�m��m&�Hm$��.�-���QmpH6�mm��l���t��ͫgI��@h�m$� I����[�����ƗK����  �l�������pm��-��-�` [M��� ���� �K N$�6�kl�5��t�m���I�,�M��HH$i0 ��-�!VP�hkWM�[A��t�@H-��5�I@��ډ�P����\ }���� ��[��+ji�L&8�/%݀ 	����n�V�N�n٪M�%���  	�Ͷ=��� * ^U�v��t�T9�nVœ(�N� q�Іcg�1XYw��ظה{x�]�Dî:��ɶ��`���3��v���[J�U�y�NnZ����X� �vÒH	4^���g���؀      �ݶvYYk[�l�$��r� 	M����  �[]mlJ'f[M,Y�	e ���$�onl9m8���f���h� ��Z 8     ��i0 6�,��m�8l  m��m�m�d[A��  Hm��l�9 � pR���l 	6�[�L�ۭ`�l�M�P�� 6ض�-��m�	��N�   �  p  �p���i�� �ۅ�@kXl�!Ā ^�[A�I�m��Ͼ��<  �l�  �    ��$q �`-�$�km��5n�� C��J�  �l�mm��u�Y�	��e m�m�f�z鰐   6�  p��   m� [v�km�۰     ��)   ��  @$  k��  M�$  mk��v�m9��}���   ����Im �` �ͻ`[AkM�l�N����      ~� L��m�  /^p��۳�  ȶɶ�� k�M[Pݥ\ 6�ͷju�@��i�$�	9n�$�hk}%�kRb�u�-�  6� 8`snݺ�I�K��&��\sd��'B�l��E��k;]JIm��u�i3^��E�l�]��J����&��s�r.��N�Wil�Ua!!��m�m��d�� [V�i� lrF�  �6�V�� �l��6݌�     ]6ݳl�`�רiۭfհ@��ސ  I�6� n�O�$h�#�t� m� pi4�6��6��ݻb��p[Ki��`   f�  �  �)��m�,�mn�hl� -���,զ@6� u���}�����qi�m���.I-��(v��[Kz�m����@-6   |����ӧ q�l�c��m�v����ޭ+1֛Hm6ݜ��m�  ��ͮ�i���C��m6�X 8-���nH��[N�km�e��cm�&� �.��l�ۛT�L�2  �t�Y1���e �7]��p$Kj�m��^v?�o�2+��e�2�m� �,IS��גMٶF�2�d���l��ͷ�'�~9�4Ν:g�E��Ν:m�m*A�M����ܵ�6�m�8�ܦ��:�f�I6Ѧvt��o��-�I��&Zq��m[K�&ݷk��n)@ �D�c^���ж��ڶ��m m n�&���}������i1���ݶ-� ���l  �	�\�f�m��m m  !� l qV��6�mm�M�`���ݱ�`	  �n��e�I/N���sMP�h�$�m�X�W`[c���9V�t� ���Z��6�G-��$'M�I�&�7Md�h-�2R{J�t����f�N�3�si:W&]6  m:��m�!�����L[@ �Ͷ�cm�=��m:f�n䚦����m�l�f�A�5��l� �cj�Y�*��l9ђ���J���vF����֝-���᱙W�f��֖��ۡ�v���յl �[M9%  -��t� K�mt ��  �: )�K( ���붥m��`�i m��������' 8�����6�@m�i�	V4�m� E)�� Àm��q��m��E    �زҸm� m�6��e����i6�mF��קN��mmf�kZ�n���kM++b۝8�� �5M@�V�m��X` ��   k4�-�m�4�U��L8[M��m�4�n�ٶ�M�$ֵ��sC@I��h�8-������F6ړZ�%3D������b1'����6tp�(b��,~]�����"�?"~X��Q~>qS���FȀU�qD���\@�P7�����~W�#�xpSN�@؀B)��
��b��%* @SX�&�1 �Fr��ٟ�>H�,H�B?�T��C|�/A���� �:��*��%���? |���&"��p�P��/�A��('N��~d	�U���P�*~g���@
ǀ�1�4���H�c�B�
��Z���������P�=!� �#����:QhN
q�?���uC� ��`��TS��^������?(è�u��C@��8
\P8Z���$? ?�+Z"'�P��&Z�����AS�p�;�:p /�@�u M�P�� D��~t$&����`�0�D����*J����&����JPCPg_��~�窦�`a�8h#�^�ϕT�41����"�BA�z}�C��]k�D,4��@`@D`���QS��A]��S_�! O��%PH�0j% 
H�b�V(�`Ƌ�b� �j,��������?.�m��F�-��v��ׁ��'@m� �m��5Ty�d�fK��a��6	�ejS�V�9�Q�H�V��Ǘ��Xa�b��O)ѱY�[�3�v"!T�V���Վ�˭��M(ڪ�9ֳoK�$�v��4�3Wc�_W$#��V�v��#��mݥn�t��K���c�i�[�Y�,��Ӧm�f={E���\�@T�u������r��Ҵ�nʰƳne�"�)w,[�5�v�6�Y4VzG[���z0��m���Yx�a�ݓm�6�C��u�ͤ�u�[i�dzZ/	J�E�*� S�AA�6��^�-�r$3�n���-��aYN����*e�e�쩦�ې�hq�@�m]<tYnT��E'BI YL�:SJ�����9C]�⣭�̺.�GnJ�
-T�r��v��b���d���ܹ���F�H��N��q�/nn탶�N����`��p��M&���q4�	��6u�p�ܸ�Ayj��v^��L�I�8$�&�nkm�I[\�pՐ²�x%�����g������ӻ]a3q�[tvF��GA�]/n�B���̑v��{p���}�ٰ6�%�'�,�6�{Z�kkM�Y!�/[ �c��1jY"{j��"��f��kp���RU/6[ �m��n�����֒��n-��$���)᤺fזi��md9��8m��im�-�A��u�I��M��Z��cê�F-HxN����{O&1���.s��2���`��Ůp5�Έ�+)�%m6�pK�R��6�v�C�0�b���H�W�tnX��]�t��9Yd�n��lhY��ZK��їk���g�v���ʚ��*\��2��Z�&�=��:�b�'�n�66��i�T�:ֲfv���m������l9�[Ƃ��^֠��r.��v]���(-�t�q���gv6@�jjNh��LYu�]2wk��"DY ��E�т�h�Kgq�;��U���*�2�����m�z����������{�t�i�L�q�Db!"?�l7�sH�
��6(���a��z ��ߤ:[.i�S�v�d�;v]Dp�頧��k�t��^�I�D$ޗ�s�bS�Ta.��x�M��-�=O-���	�ҽ��:!u\�#��\���s�c�hL�!��s�������ۜB�N5����@��F��㇃��f����t��������:���s�=p.���r�Ͷl�i��g[��ѢJ痮V��������^�y�o�쉑�97	�w�ܼ�9^=�����c1����"�wu��;����/z�����ˉ��<� �v��\��6���5�m`I��y�+��7�A�C9!�[e4
��5���X�^�T�uYcL��m8h{��۹�{zSB�-��-v�R(�F9�����-�s@�v�I._�V��6��]M8�n�K�X�ռ�l#[�ם����u�q��������dc�"�rs��w�����|h�M����w4����R��L�`wuqt�+�Դ|Ԫ&�ۻ&7�����Vv�pc��f_��RC@��@���57ݗ����������C��+]�]`I�56we�n��u�%`\|~i�\m��L��{zS@��0���I1`�&��(QR�O���ݹv�D]�i҂=���+���h��\�='j:Lp�C#�"�	!�[e4^��m��=�)�v^���"c��uf��wv���XӷIt�9[AG�69�����-�sI?w�vnpleA�@-�#1����W�@��z{qJ�����(��=�)�^v��������X�My&&�^v���������4
�P¤��� �eΓ>)�n^��R6[�m5���xcO����ܼ���ٴ5Q�m�?���͋��hޔ�/;V��<�4�X�I����i+���y�mY�5$��}�����o�� ~~�߻����Y�3<�$�ғRI^��<_g���ϚԒ__��<�$�T�i���b����J���6ܮܧ���d��~m�4'�1���ߕ���nkv�{�̏Ȑ�@�&؜^x�U��jI+��������n�o~�{y�m����59�Kǵ�<��'\�#��z�:s�F�M	֢L��n�D�䓡c]�N�[6��]f�6�ٻ�~��d����������m�K��I%s�ſ"AH�2	0�g�$�zRjI+���%_J֤��o���K�.�ǚ�8�LM�jI+���%_J֥�o���g�$���RIZ.6�߾��V������~}O���߿���	�&����W�$��d1����O ����m��O������s�fi�m�o޼��>�r��m�;0�R���J� �*9�WJV 4 P0i��EH�@b�$Q"�E7&����LDҍLLT ?I�˩�>����\�3 �Bl�M:J��m�޽��6T�ՒTY�-�����t��Zm��%�N�;E�-�[�6ۦНΰ�8ѭ���3�n]Ѷ�#��n��y�=��!�[K�J�iz]�gVt��flv��U���.$ܫiX)ZE��7��v�A��/*���_J��M��D��<^\b�[I�l�����<N���^�b��2ڵ/%r��v�23��m��.ۋc�]�ƭ�8P��c���:���y6Gg��$Iٮ���9eְ�~� 7߷�| ;�j�Ē��kRI{z��x�^�S4���dB�$&���e��?�a����ϚԒ]����Ē/JMI%}���ȒB��Ĝ^x�U��jI/o_3�H�)5$�{-^x�U�p�#��1��.�<�*$�Br}����H�ω�$��j�Ē��kRI+���$�bq�273�H�)5$�{-\��>�r��o�����w�.��� ���Zz�u鮽�yK���2�V�N���v�1C{;l��g��v�=F[?��ou���r�r�6��v~Z�8���z��X >���~չ�!j�����~�� |�B�= �k���}�r�_�G�$��j�Ē����[M��
H�kRI{z��x�Ut�Ԅ.�Z��$��ZԒWۛ��q�# ���<I}��qV��+m�������v�<m�����x�^�S4��b��M,�A�I.�Z�~m��۹�_�m�f�_�6�}�V6�ꟽ���ŝ�çl��g�5�d��Yˑ�(��᲎�:���yz� �8^$��Ē��kRI{z��x�Ut�Ԓ]�y�IWaq)HlQ�hN7�&��������UOv���s���~m�U%? ���ßނ��B�n�� ��~(���ܮ���Z�KL�+���NT�z֤����y�I{��<�L ��RbԒ]�y�IWekRI{z��x�V�����~��V��6��?? ?W���$��|�<I+]�Z�K���<I.c��?^�0f��:��]=�����W�Rq�u��V�xS�×Qȹ�Uu��Ԓ^޾g�$���-I%��W�$�vV�$����&ЮH�173�J�ݗ~\̷�k޼��3��ݶ����9�*��>��q&�p�j�� ~�o�O�J�kz�K����Ē��ũ$��V�~F��.�������_����������ݗvހ�8PV�I�����^���%밸���lQ�hN7�$��|�<I/��}�/I^�|��$�w�~ ���?w�Ź�}���e���Khk]]9/*,N����� y��!rm�̯:JYK�������������O��յ�I%���y���0x�Q0��$QkVn�oߵ�����
MkWٚ�V6�����~m�*bx�o�#X�K�>VHE�/<I*ݭ�I/om<�$�wp� ������u�y��U�*�I%���y�IZ��Ԓ^t�y�IV�oRIw�717�\��bng�$���-I%�KW�$�n��$�����ĒY������������^ܹ�g,Rn�l�U�%��]�O�*/J�K��z����ӥ�u�v8�F�5����`8�0����=�W��OϢ�[k����v��r�n�S0�E���w�;]����ptixu�B9��W�X�`�M��.�t��n,;\�nd���d3�8�t'�eD7�on�qɮ"�Rr�ɴ�g;q2�Iۛ�۫Z�+��M���|����|M��/nz���'������n�Xx�:�O��`�E�=��a`�1�M�N�7j�rI/~����J�kz�K���y�IZ��Ԓ^S�M/"�$؜^x�U�[Ԓ^�_3�J��z�KΖ�<I*�*JD�6(�47Ԓ^�_3�J��z����l���%��$��n&�#N#��G!�%WJ=I%�KW�$�}+Z���[�g�$��]���D�<�eU����v��1�\�9�3J��o�o��%_J֤��N�^�1�<"jk�N�M��e�4\�S����qՀ��(Ǳ6g��͸�բ������~�����g���m���o��۹��ͷץ���r�R���_��߿���}��wn�
A�bB*F�l�4��M���g��,�Q�$��j�Ē�����nnbm
�䌃s<�$�K�Ԓ^t�y�IUҏRI^���Ē�ҽ�a�&1�c�#RI^��<I*�Q�I+���x�W��jI+yV�<�0s؜^x�Ut�Ԓ^�-�<�$�K�Ԓ��]��-�� �z{9�[5�IXMi5���S�Y㋘ŧ��<���j�x�#���r�:�4j!���K���g�$��u�J��y�IUҏRI.��n��ֲ�D�h�-��k��~U��}�{לm�r��m�V�ߗ�ͷ�m��,e���Wn��1�����~m�v��.%��4z�Ҹ�
��D5���*)>��*�6ij~`e�OŨ8X��(��H��FBC�T?A=� �����c�>IC�9A������5�\�������*>O�p�8���F��HZ��c	�HIEx�������8����^�vF�:�[��	�S��) �F�#���}kB5!SK�S��}��p:��
p��h<8M
���
�G��3�	T�%W��l�~�ÑUM uP�ۥ5�ɮ}�����Z�Y:�����E�yz�Nɋ ����7�$���x{��6?�M�n5��w4}}V�;R<�ۆ�qqq'�57)R�R/��^�c���a͸�#��ە�>��5�<@�3P�ǘ�B��l��9�y���/;V���M�����u���,��Ъ��;R<ԓg��� ٻ� ���[�͟}��l؁ �6'��}>4��h����h�
�ph�OpШ�w4��Z�j�D?�Jڨ� �u*|�ݦ�^�M�A�̒90rf���~��ݵŁ����Ub�����e���uv��������r]l�������ݥ���lU�%�$\Ț��'����@����z���}V�iVjŋ����E�yzS@�n�޾�@��[���ƞ7􉵍ƣQ�@ٻ� ���x�H��K��*�%1P��`�Nf�ﯪ�/;V��S@�n����_��bɌm�@���홧�6n���'jk�;�.'�ww�<������H+�ff�3��\v�½��5�fJԓ&���U2�-�Sv��PG��]�v�q]�A�w.RK�N����]Y��B3���x�)����W|����۪,������Kː��=���cp]�A+:2ێՊݞl`v�K��c7�<�e�Uܡ�;s�`�.eF��N�n_g�I$2�EEn�i
��{;s)�l���ڧ/Q\M�����{��>s���-[u��󄃱v�ְ;~o��?<��\��s�n��9-ù ��6�p���:�>4��h����h�
��n!$�������@��Z��M �ki;�&�$�I�s4}}V�yڴ���{�O����Z	ᨁ�$MH�9ڴ���ޘd�0��ǀ~�h����0��I$Z��M�]n�xs�-�v����+fHҎbQdQ=h��f�	�W@ls;����gd�G2=���w���Oa ���j8x[>4}}V��jG��s��_��U�z�?�t�D�d�E�	ST�_&��>�woL���縕Q��W.�V��b��� ߿~���ş�JP�Jg{���?x��ߖ���W�f�	 �	��h{e4�S@���h[f�}��9?��$�6�u�����@:�4/Jhgp�+P�cȱ)��n3�}ck7(&������CYn�xL����I�nV��H���5!��޾�@:�4=��[)�yŠ��8��Z�٠yzS@�e4��Z��:�I��nM�Қ[)����B�Oªb�s_g}Z�[4oC�7�7�\0�]� ;$�q���`�3iS�vݻC]��T� �K����'���.�ޚ��U�?*UI�zM�x絢��Q�`{kgd���Vyݤ�A�;Qӯq�Y\wLMZ��������� ��p�;%�R���n�Wf���`�`�*��������7޿��< ��R�9ě7�f���ʫcn��� �����#�W9�s��n���O� ���䑷d�r~�ؒ�����������ZM+jƘ�(��"�`�1�R:�N�$ҿ�i(���`w�|(�(-�ՖS�x�%����i�	�z`��Z�����G?(ӑ(��zf��y.��-�-�;OJdN,���:v��r3������pŐ$	����hzS@��j��f���A�N�A2H���3�y*�J�� o�׀}�H�x�=���ƾ$Ą�4���@:��57����&�� ��%J�bj�LUuoSsf�����;;p���I���=7�J����aTWx�T� �8��7����I^�����'>�A���&w�X�ܭV���ܺ��#�<�6�l.0�ƈ��]�GKu���p��pE`ɹ�i�^6e�hƘ�<'^nTv�F��T8����i�.�W<oHgj��bN�^v��N�']���NvP���Uَ*�v7�P�d�UJ����썵�Nk�19G.����K6�7%������:k�$�}�5�N���iQ-��0�su�U����}�{���|���n�q��1��[cqK����7On�����z]�Dl�;n���|��gˮI6'��O�@��j��ϳ��}ki}�F�ds#�G�]��Ē\�)�S7�����<�\08��Q' ԋ@:�4=��y��z`�Mx�F����Z��	ܚ��V���h����+��M���ǉ��54�S@�����n�������N*�Mt[��]��Ď�ڻ,v�<=W���ٵ��愃���uw�y>lGɆ�����w�m���M���<Y���� �JI���X�u]���(X�"�P�p��KA)��M���7$��׍�_U�~H���x�l@�D6I�}ݽ0�p���򪒷� 7����
��c�5��n~W��@�s^ vIx�9���y��Y^Uun��uj���Y�}�v<ޭ���^��:�M�{*x,��,l��X����^����Iǖ�޺�D�s�;Z������հ��kuue����<��޿�~wv�7oOs��}ښ��֭�ut�0�V�� ��e��\����������������$u��ǉ��A<��ԓ@�{^��s�}۹���  "'2g�������U�FR���.�c��x���5�����v^�9��`����I��&1�28���@��/�6�7oL�����&�V]'c���vղ��Q���9\�GnN�f-�������mBw���$e�k�m���xgn�G���wo �l�M�!��&���:�M��${�Mݼ ������mjwv�]��];�0�wk ;$�<��Q&���������rպ��t�]`j�swo ;ٷ�vK��W�6�BI��*H(b� E!��+F�H@�c��B��!
i7i6��=U�́��	�2,x�B%nM �޳@�2���x���h[f���[����f1Z�#�,t���#HNq��/m;�Y@1ٵ��N3Þ��H�3�-�rU������`�� vI~\�_Po� �W�<���91�I�]�}���o�@;��@�e7�H�Z��1&1�2;x7v��ݗ����*�޿eo�}�[l@�D6I�����hv��?}]���swo ���Ww|�]�N����.�}&i�n���>�ܐM��,#��@ ��H@�Dd�? ob1"	�0D�k�*���|���O�9!6!B+�"$XD!$H�FH"D��D�X1���
��aH��P�_���}���s��Ο���Ơp"�2	n�!�	0 ��bFH!�5 �'�!� j4���a+.���uv��"A8��D7�Ha� ŉA�E�����C�_<�Iy C/���F»�aX]+V�Y ���IbL�x���F00X)���0F�3�
��]�]�N���r5D�b��� �6:���c
����H]�/v�h����y�PX
v�	�G�mf��`�6� ��m�dֶ���ӭ����Μ�k�t�Kv�m�[7Y[%L����Rnۢk������&��t.Q8*+ڐ[iF������]�]��t;:޽y/Xi{2�����d�#K��k��b���U�2m��Ӥ�nE���6��r,�=q�\�^�=f^��\��ѯ���sMa�U7��k���.3L�z�)���Bi[�u����m$�����IdKe�tֻp՛�-��(�j�l���v�zM����p�T�P�z�V� 1�1���Y�r�|�'�7|ƾt�&W��lI']�����7.��9�vs���v�&�%�)�"��ŀM%B+�Q�glAu�Pq�qT�q��[u��6������]�ɕP�:�3]��l6_�����.�Rly8'���(���5�8���&M�$�ɶ�\���BMgI�\/D�ս"��m�f{(\�W�-h�66.s]��II�Z-ܜ#Y6]6�7St���0i��`;k��F�KV��^�M.��N7�3���k�ۍGWam����mNW;	hEjTH�F�Y����/�d��!∡6�j���7lMӕ�Ј�[Yͤ��N�+U�mu*�Ş���e�ݹ:m����2`��925:�6��$��M 4��e���K�7@n�7��ᓎ�iYP��nl���m$�۴�.� ��L�;YK��q�n�N�v-�g.ӯ'jV���<Β�ڰ���6�i�4��m��[N$l�n��<?0��P�Hɦ`Rබٷ���N�l�gFuĻRc�Wf���ۊx�f�0$v3�U[f��y^��t�N�`���]w�%c�QG�n�vI��ܝ.��Y��Ɓ�j�-��t�m�M�N��\�j�\����t��Gj�,�!��k�vˉ��[�lxH0�-ꨕM���gm�Yd�����kl�M�ҁi�^40x�I�e@�W�'$ф���Af鬺J��r�c]�扫oY��5�٩�^���|i�p ��C����x���0>��? @N��C�c�����g.��lm���E�r���Ӕ�x�+�6�N΀:RjWq���n�t�&�h��[ɴˬ�"ȤYb���U���s�g�g�!�t���m��!ٮp�u����\�r�g��dYpv�R��x�KX��h�j�t�yU�D�B��p��쉻8�oZ3׳a�f����.�n��Z$:��'[���ْ�y��e7]�s��}��7�N��P:����w�w����wp�_�c*�r>�ǘ�G�k:t�!�u�nTU�^[�q��c�-���9�9�����n54�ύ �l�<��hl���Z�o�9�D�p����I��S^7oO�L�g8��4�w���oq���N����ڴ
-m9ı,O��}v��bX�'}��m9��Q"}�o�m9ı,K����l�A#�&D�,O{�na����ոjk2�j�9ı,Oo�m9ı,O���6��bX�%��m9İlO��}v��bX�'�l��x�r�h��Z��r%�bX����m9ı,[�{��r%�bX�����9ı,N����r%�bX�|Y;�m���ô=fS���l���k֮���S���,I9j�������C�`q���d+|ND�,K������bX�'�뾻ND�,K���6��2%�b}�o�m9ı,O�{�%9�%.Yufd��kiȖ%�b~���9���R*@Ah���Z�*Y�K���6��bX�'���m9ı,K�{��r'�"dK�����^|�����w���oq������Kı?w���r%�%�{�{[ND�,K�u�]�"X�%�~�������n��6�����{���7��{�M�"X�%�{�{[ND�,K�u�]�"X��0C"{����iȖ*�k~��&PyҨ�SEML�mxj�K������bX� �����9ı,N����r%�bX����m9�q���}�����P����2=vn3�]#plѮ�v����69۰�:݈��
��ww�;|~s�j�(��������ow����v��bX�'}��m9ı,O���6��"X�%�������bY�7��ߦ�����Xzԅ=ߛ�oq�ｿM� �X�%���ߦӑ,KĽ����"X�%����ӑ?�ۻ��{��7����`�<��Þ`�i��Kı>���6��bX�%��m9ơ��1���2&D��߮ӑ,K�ｿM�"X�!�����;�뜦A�{�7�����b��3�����r%�bX�{^��ND�,K���6��bX+b~�~��ik4u
&�&Bj��R	"sﻤ�E�#;{�ͧ�X�%����6��bX�%��m9�q���?���}�l;���g-'tM����b� �<u���^1��6��9o�����5^��V��.j�9ı,N����r%�bX��ͧ"X�%�{�{[ND�,K��{6����2%������sZՓ2��k.�SiȖ%�b{���N@,KĽ����"X�%�}�{[ND�,K���6��X�%����8h���]Lֶ��bX�%��m9ı,K����r%�bX�����Kı=�{�ND�,K�z�y�f *������k�P5���~�V׆X�%�����M�"X�%�����r%�`x~�@b Gj�0��1U �H1`��Qj!k�ڦ �%��H���'����|�~oq�������7̽����=�Z�r%�bX�����Kİ� {��i�%�bX������r%�bX���ٴ�Kı/�BY�3	�4j�=�ƪy,wsc����mzNr����d��[�ǟ`>v~r6�|�~oq���=���iȖ%�b^���ӑ,K��w�ͧ"X�%��{~�ND�,K=�����ۋ�Shg��{��7��{��[NA�,K��{6��bX�'}��m9ı,Og}��r%�bY���{��{�68LF]��{�7���{����ٴ�Kı;���iȖ%�b{;�fӑ,KĽ�}��"X�%�������m��� 8�����{��"w�ߦӑ,K��w�ͧ"X�%�{��[ND�,K���]�"X�%�����eh6��&�=ߛ�oq��'s��6��bX��3������Kı>�׿�ӑ,K�﻿M�"X�%��D;��\��lԗRB�m5�\��*ѸI$�neF�Iy��.�G3؇����)�q��u���8�j��+�k���;sV_7>�GLJ�y��
Z�.ik�ַ;Z��yލ��H��/=�r���v�2��Q�m0)�C��|l�	�n�c�ӳ'H���6ݧ��������{q��)Ǒ�*��&�$�N�j�u��Mٹ�����Īi�����rO:ZZ������=\��E����Y�WZ�n:�vfnõ��ղsu��Tܝm�[0�.G�z�nh������7���{������"X�%����ӑ,K�﻿M��n�Q,K��fӑ,K�����;|Ź{mV:F�����7�ı?{]��r��"dK�����r%�bX����6��bX�%��m97���{���o�{}c0��a���̖%�bw�ߦӑ,K��}�fӑ,K��;�fӑ,K����i��7���{���}>�?y��{�2X�%����ͧ"X�%��w�ͧ"X�%��=�fӑ,K���ߦӑ,K�������]fY5sY��Kı>��ٴ�Kİ��W��{�6�D�,K�����r%�bX�ϻ��r%�bX�=җfId%�]Ml]=[s�\Xy3Y������c�d��[<'nvٰ�/�WXz���
=���7���{�����m9ı,O���m9ı,N���m9ı,O���m9ı,N�]�7�@p���w���oq���߿>ͧ!����&�X��sٴ�Kı;�{ٴ�Kı?g���r'���{�Os����m��id6R�&�ND�,K��fӑ,K��;�fӑ,K����iȖ%�b}�o�iȖ%�bw��.pѬ�Fjf��fӑ,K>��.w�ͧ"X�%����ӑ,K���ߦӑ,KȞ�}��ND�,K��ԛ���f0֍SF�5v��bX�'�k��ND�,K��ߦӑ,K��}�fӑ,KƷk��k�P5P5�Q�� U*��&��i�_7���\N�*�4�u����`�̏i��㞘�.� ��w���ou���o�iȖ%�bw>�iȖ%�b}����Kı?�}v��bX�߼�}>�?y|�~oq���b_�{��r��G"dK�׿�ӑ,K��u��fӑ,K������Kı?���̟з$-Յ�53Z��Kı;�{��9ı,O��}��r%����k��m�L���o�iȖ%�b_�����Kı>��{�68��F�=ߛ�oq��ow��~��m9ı,O�{~�ND�,K��}�ND�,�U(U2'{��M�"]�7������w��yz������,K��ߦӑ,K����m9ı,O�w~�ND�,K��k6��bX�'��w�Yy��P֦C[�I|u�>��V�K�����k�e�u�Y�3ۤ�[5�4�e.)�Ϳ=���7���{�_{�6��bX�'�뾻ND�,K��k6/"X�%���ߦӑ,K����.pѪf�֩.k6��bX�'�뾻NA,K���w�ͧ"X�%���ߦӑ,K��;�fӐKı=��6g��ch�5�����Kı>�]��iȖ%�b~�w��K�,O���m9ı,O��}v��bX������cB�P?=ߛ�oq?��{��iȖ%�bw=���r%�bX�����9İ:��v?"���O{}���r%�bX�1��͟���{�7���{�����߯�w"X�%����ӑ,K���ﵛND�,K�{�M�"X�%��w������/<��wn��6���z��˴v{:���zps�K�0��5���/������n�Y��ı,O��]�"X�%�ߵ�k6��bX�'��~��,K��>�iȖ%�b}��[�5d��]Y�e֮ӑ,K���ﵛN@,K�����iȖ%�b}�wٴ�Kı?w]��r-�bX��z��C�E��f��ND�,K�{�M�"X�%��}�fӑ,�a�2'�׿�ӑ,K��u��fӑ,K��=�K�ե3.���Y��M�"X�%��}�fӑ,K���w�iȖ%�bw�w�ͧ"X�%���ߦӑ,K������N5Lњ�&f�iȖ%�b~���Kı;�w�]�"X�%���ߦӑ,K��>�iȖ%�bq6pg���o�����w)�ȽJ�t�S���D��[�:�\L��G��5�Ȇ��Z3� X(��%���NNPr�c���`SX��A筄��rq��{v�Z��e�s9_/..�B�c����9/H1qn�BQ�\��[����f�G�.���ǎEN�@l�
�I���$�J��Qrۺ'M�_$9���-�u�R�^��:�Ϋ��J�1Zw�{��w�����n��6�xu`���g�j�9�7-�#{c������ד��g���qw�L���kW3WiȖ%�b{����ӑ,K�����iȖ%�b}�wٵ�KıY��E����Ϻ�ꒉ�&d�5nf�v��bX�'��~�NA�,K��}�ND�,K�u�]�"X�%���ߵv��bX�'����I�2ܷZ�-����Kı>��ٴ�Kı?w]��r%�bX�}��WiȖ%�b~�w��Kı?{���K���决Zͧ"X�%����ӑ,K����ڻND�,K�{�M�"X��C"w^��m9ı,N����岖aufe�5v��bX�'�w~��r%�bX�w���r%�bX�����r%�bX���z�9ı,O����;���!��9��8�+����:�=�
���y]�ܖvڕ�k�-������sZ�O�,KĽ�����Kı/�ﵴ�Kı?w^��<�bX�'�w~��r%�bX���=fh�Lˢ�h�sZ�ӑ,K��;�fӐ�wBtk��TRu
�! 1h�w��?D�7�^��r%�bX�����ӑ,KĿw��ӑFı,O}�I�$�T���.k6��bX�'��޻ND�,K﻿j�9���Dȗ������bX�'s��ͧ"]�7��￿�|w��>:�Z���w��,K��~��r%�bX������Kı>�wٴ�K�����NOq�������������V���D�,K������bX� ���iȖ%�b}���iȖ%�b}��ڻND�,K��H_	̓՗Z�z���u\0\�sr�:��둹�N��l�(K9+���ͻ束�2eF�{�7���{��g���r%�bX�g���r%�bX�w�����P`�dKľ�������{��7�������M���4��~d�,K����ND�,K��~��r%�bX������Kı>�{ٴ��x��{�����ߢ��0nx���~x�Kı?w���ӑ,KĽｭ�"X�<}ć�?�s�6eM
��@��(� �ȓZY��]hM�4z�l�� ������U`�\~eb/�>	s?��?ځ0M`�5��@��RD�jY"��STр0D"��?K"j2ͅ ��
C1�+ �	[�w8����U?n��~jqH?���H���H�:��M�e��~5���QB�"��9�� �b�]lv�^�b���`�U:�4�Wf� 'Ȉ��'�t����l8�S�~��f��m9ı,N���r%�bX���z�֚�%�5.kWiȖ%�bw���ӑ,K��=�fӑ,K��{�ͧ"X�%���ߵv��bX�'�}��f�L��L��˭]�"X�%��{�ͧ"X�%�w=�fӑ,K����ڻND����2'����v��bX�'�A�ݎ��h�8|0p͝O]���tf��1��G�늲���-�oOm��y�ݮ�:����g�K��"{_��ٴ�Kı;�o�.ӑ,K���]�"X�%����]�"X�%��v���ja�5�jj\�fӑ,K���߲�9ı,N����r%�bX�g���r%�bX��{ٴ�Kı;�n��k3Ym�SY.f��9ı,N����r%�bX�g���r%�bX��{ٴ�Kı;�w�ND�,K�O��2e�ՙm�M�"X�%��{�ͧ"X�%��k޻ND�,K�w~˴�K��2��;�o�iȖ%�b~�w��&e����f��kiȖ%�bw���ӑ,K���߲�9ı,N�^��r%�bX��{��r%�bX��>�ݎ��ʗt�f�ʜ=n��mr�;SUx�팃�FJ��\,Y�r0`�FS.�v��bX�'}�rͧ"X�%��k޻ND�,K������bX�'}�z�9ı,Ow]=fkMsIdɚ�Y��Kı;�{�iȖ%�b^���ӑ,K���]�"X�%��wܳiȖ%�b|g�=fj�ɚ&]]\���r%�bX������Kı;�{�iȖ%�bw��,�r%�bX�����Kı=�O��4j�њ�&�Z�r%�bX�����Kı;��̛ND�,K�׽v��bX�%��m9ı,O{��L���Z&��fj�9ı,N��s&ӑ,K��@c���]��%�bg���m9ı,N�^��r%�bX���  �x���8�aP�&"V�1@�B�����dWw����{���q��ܛŞ�֑��ƽ�r ��fq�92N�3��ђ[���C��4���^�m�t��n|���Mơ����3�͑�%&<��W��7)�ҽ6�$J�&�Z��{i���M�nEr����Kk\�UX�=��e����xt6���l8�P������g�P���m�{]�J�N;s۬��ە�����+i5�u2���w��w�|1���M.����s ��=�j�a{;����;W;�.3Þ��n,TN���Z���%�b}�]�"X�%�����ND�,K�׽v��bX�'����iȖ%�b~3�_�e�,֬�s5v��bX�'���m9��DȖ'}���9ı,O������Kı;�{�iȖ%�b~�^����Kuar�5��ND�,K�׽v��bX�'��~��r%����2&D�����ӑ,K������ӑ,K���߿T������|�~oq������w�]�"X�%��k޻ND�,K����ND�,K�׽v���S"]������+ϗ���*>{�7���{�������r%�bX�g���r%�bX�����Kı?w���ӑ,K�������2��#��[��{:m��Z�n#&�XN��pc�H\�g3��x�12�f���v��bX�'��{6��bX�'}�z�9ı,O������Kı;�{�iȖ%�b~�����4j�њ�Թ��r%�bX�����(��|5󀉷q9�����]�"X�%���z�9ı,O���m9ı,O}x���h���u��"X�%���ߵv��bX�'}�z�9ı,O���m9ı,N���ӛ�oq���}�~n>�8]e)��D�,�@�;�{I�$�}}�fĐI���M�$OD���ڻND�,C{���C�x��G9������7�������ND�,K�����Kı?w���ӑ,K���]�"X�!��Ϸm�~��H�;Cvc���|xۧ��AªC�6�5������@ɋ�N���8�Z\�j�i�%�bX�����ӑ,K����ڻND�,K�׽v��bX�'��{6��bX�'����s��r˫3ֵ��Kı?w���ӑ,K���]�"X�%��{�ͧ"X�%��{��r%�bX��z�֜3,Ԇ�k5��r%�bX�����Kı>�{ٴ�K"��� �T֍ı3���ӑ,K���k6���{��7����;�T��:"(���Kı>�{ٴ�Kı;�o�iȖ%�b~��fӑ,K���]�"X�%���.BpѪkFjkR�iȖ%�bw�ߦӑ,K���w�ͧ"X�%��k޻ND�,K�k޻�~oq����w�}��~��H�ؼ�a���J���v+LĲv��Ļ\�ۇ	��Hg�e��ɩ�մ9~{���oq���o�k6��bX�'}�z�9ı,O��z�yı,N����r%�bX�=���赇�R*~{�7���{�������Kı>����Kı;�o�a��L�bX�{^��m9ı.�]�x�v��l8X�����{��"}�{�iȖ%�bw�ߦӑ,ı?w]��iȖ%�bw���ӑ,K��}����j�2�5��ND�,�H9�����ND�,K�k��ͧ"X�%��k޻ND�,|@�sq;����Kı>�o�ۜ�[�]Y�f�SiȖ%�b~��fӑ,K���]�"X�%����]�"X�%��{~�ND�,Ky=�Irq�}�5�]�%��ぼ���<u��wdG��/d9b.��<�Fvji�����{��2w���ӑ,K�����ӑ,K�ｿM���L�bX�{^��m9�7��������T���;V�>{�7��,K�k޻NC�#�2%�����M�"X�%�����fӑ,K���]�'����Os���~���m��G76�ciȖ%�b{���iȖ%�b~��fӑ,K���]�"X�%����=ߛ�oq���}�������@�uv��bX6'���m9ı,N�^��r%�bX�{^��r%�`<��������r%�bX����t�뙩�̸jk.����r%�bX�����Kİ�����v��X�%���]�"X�%���ﵛND�,K�ت�	ŀ��8h잙��}f���z�#GO nT�������tZ![�\ܠi�k��l���~v�hn+m��ݬ�#���W���v�݌9��K��Bz �m�8�nŠ.��^�KE�'	�n���ѥ����{I1v�C�/n��J�)�ے2rl��h]����%s�d�7.��9UڽVv����=S{��C:�!Ws���;� �.���\�浴Is��5jc��w�����vM��<���ݞ��λW^/m�v�1��q��9Z����9ڷ���������Å������oq�w����r%�bX�����Kı?w]��iȖ%�bw���ӑ,K��}����j�2�5��ND�,K���6���,"dK�k��ͧ"X�%���]�"X�%����]� &��ow���~�?b3�j�=ߛ�bX�'���m9ı,N�^��r%�bX�{^��r%�`"{����i�����ow߷��)^�x��54��Ȗ%�'}��m9ı,O��z�9ı,N����r%�`A0�����8�L�g8��Z�hn�&�5���r%�bX�{^��r%�bX�����Kı?w]��iȖ%�bw�ߦӑ,K����R�WS3:VNk�i���r�e�����.���s���I��"%T�������Ό��nm@��w��,K���6��bX�'���m9ı,N����<�bX�'��{6���oq�������9;j���{�2X�%���ﵛNC��B0Ck�.�D�K���6��bX�'s��m9ı,N����rX�%�����w�s�֒*~{�7���{����6��bX�'��{6��bX�'}��m9ı,O��}��r%�bX����x��	�5.KsSiȖ%�'��{6��bX�'}��m9ı,O��}��r%�b؝����Kı?{~���-5�̲Mf�ӑ,K�ｿM�"X�%��,~������ı,Oo�m9ı,O��z�9=���ow߿��ۻ�P=b��t:�����ٸ��v�/Z��<��q
-�w%���������皷�w���oq����ߟc�D�,K���6��bX�'�׽v��bX�'}��m9ı,N���̛�抏����7���{�~���|NA,K��=�fӑ,K�ｿM�"X�%���ߵv��X�%���Ӿ����ڵ6�����{��7�����iȖ%�bw�ߦӑ,z��b RB>U��D�Ok{���r%�bX���ߦӑ,K��g���TѣT������r%�g��2'����6��bX�'����v��bX�'}��m9İ?�I�;�����r%�bX�ݝ�3�y6��g#o����7���{���ߵv��bX��{~�ND�,K����ND�,K���6��bX�'��};}x�Pv��Z�:}�ٲ���l6S\R�;��k�d{OG�x��N���SZ��kWiȖ%�bw���ӑ,K��=�fӑ,K�ｿM�"X�%���ߵv��bX�'�>��&ze�)��-���r%�bX�g���r� ��,Oo�m9ı,O���j�9ı,N�^��r%�bX����BB]��fY5sY��Kı;�o�iȖ%�b~�w�]�"X�12&D�����ӑ,K��fӑ,K�w���}\~�g<վ{�7���{�-���ߵv��bX�'}�z�9ı,O���m9İ61�Ah�$ ��(19~�O�&~�y�{�7���{������֛����r%�bX�����Kİ��	�f��Kı=�����KģY�T[^����]�D_�*�D�qrq���z���%@�/]aSC!�ך�=K7��x���{q���h���{��"X�g���r%�bX�����Kı?w����9ı,N�^��r%��{���s����:룛�:c��{��%��{~�NAlK����ڻND�,K�׽v��bX�'�׽v����r{��7�����r'��۫���|�Ȗ%�b}�o�WiȖ%�bw���ӑ,Vı>����Kı;�{���{��7���������W���r%�g�"�Ȟ�����r%�bX������r%�bX�����K��?w���ӑ,K�����I��s%3V�5��ND�,K�k޻ND�,K�׽v��bX�'��~��r%�bX�����Kı:�8���"��$@�P���@4W ]ŌQ=ĉBj� ֔$$������\��5�߶=:BE�ȸ�2�:�D|�����`@6J���mҖ#�(�@5Q*V1ΜD�<D�"D�����*l U�>@�;�����S� ����\�'ˣ��X8�u���M�b�$����*� �H"t0�2A�U�|��	&��^;c6B<��	^6b?"�R�Hă'��T6�4_��]���.�-�� $h�kk� ж�۰�YqѪ�!&�%M��mm�K�(-�m��TK��5n%���&��J9��9:�E;��/g��� �;V���5��d�ˌ����)t�nE�.�VC�*i���69�ŝ�J6�v�2�v�[eɥ��l��M;^{(�^��%�`�E$Z��,՝v��'[=�YܠNM(���r���}K��5��Fi7K�V7/R).�g.֙u̅�[7e�/Hix-�<��ڝ;���ʴ�*��rg�!�sPV-��>Ϭ���t�9��IF�t���"υ�l�x^ݬI�6ܰ�Nٱ/.FN"�Wk�l4��:�C'FC�#[��m�9�a룢]n{N"v��zn�z4ƞ: �+e���=��[�U�`ڋ莨ݳ�f�L�]�n�u����`�T�'�rs+\8����e���x�,�P���u�X^�u�h��y��e_Y�+�g����LV��t3�nF.����{O-�l�*��.`=5F���KPݹ���$a3i(����k �v�u�i�-�����V�ۧ\�K�=%�&��t�8�׮�^�8�y67�Z�:���I�U��:�\m<��g�U��&��xV�v�v݀U3��:F�e(Hm���.juɵY�Fp��nؐ�Vɵ��R�!Z�m���%��׫�6��$� ���i$�&NT�	�\&I�k$K����z��K��D�B�Ĵ؞;Y�۷��M̗/�꫙жN�R���(6�s6�C��#]d��ML-�m����6�mAӳ�T;Y��EeWr/��현{Oű9m�k��t@�^�&�>ɤ�sȭ<{r;�'�W�s+-����z�2jvڸ��@�q�lI�m��d��@��{P��tU��;�nr���p9��`ke�(��-Y�oY��t�Nޞ���Mz�V͈lh0a�����0��n��&U��*�������<6�t�Y��H�֦�me�ce70\\�	ڸ������s��D��z���N�UN�@۠"}t�U8<�a�'����T�[o4jܲ��
ٙ"�g7#�v½�	6�K�v�H�YVf���אrۤ���v����w�g���q�OnV�ݶ��v�p1�/)=�{b�v]{m����ٛ)@���x|�S���ϣ��`n읃�<�n �$6�5gi9�]�,Z���8y�Uܺ����=5���PMm�����C��)�h����-�����3n�jޗ�W-[\u�e���笧n��`y�GH�n˴v����b����DD�t��ْ�t�+�Md̲Mf���,K���{�iȖ%�b~�w�]�"X�%��k޻䟢dK������ӑ,K�����,��[��Vd�5�M�"X�%���ߵv��bX�'}�z�9ı,O��z�9ı,N�^��r'�2&D�=�x��k/\\F�*>{�7���{�������绑,K�����ӑ,K���]�"X�%���ߵv��bX�'��i�g��:"(�����{��7����ϻ�r�ș������ӑ,K������ӑ,K���]�"X�%��Ϧ�VZ�YV��ٜ_�&q3��So}v��bX�'��~��r%�bX�����Kı>����Kı?������8���<M�T.�G\u���T	�=�7�p�Y;i�;�ņ#rv9�������S&fj�?D�,K�{ڻND�,K�׽v��bX�'���6�$�"X�'����v��bX�'���wO鬖����������ow��������B�,��т�>J _�{�_}?}�k�/�QB�} �lX�N7Z}���:�V��t�h]�@��)��bPx�����'6�^����ʑ�y�w4�7�~Z!&�Qx܋@�X��������oLJ��N�v�w�ՇWl�ҥ�u��N��G\p�q��p�u�wm�v83۪�M&(�I?_���<�.�#�����/m�ڏQWv�2�v���>��ٻ[� �I�Z�ՠy��ʈ�d�c����=�`{v��Ȥ�JC����	��KZ�o��,�,݅\�*�QAv�(��x��6��[� �K��k�h-Q~�M�c�E#�hT� �wsO�n���?w�-���B�{|{�{q�õ�w�u!v[��S����v[����ռ�u9�Eofȸ���>��IR<�{rޯ�7ku�woD��cULv`T�7�6}%�v�^���I6N��7���l��U��>���%H��s�⪞���?�����;�er9�dj<k"�-s�=��xwoLJ��W9�s~j�����gQ�D￵����'�����1�I�h�)�Z�Z�ۖ�	*G�{�\�T���~-�4�իĺU9 �K˹��;<���On�l�<��[��g5y%Ƴ1�v�
��e��z��y�,Z�ՠ{l����%Ƥoh�����~�n[�.q%�.$�T{��<>M�z�`ݽ0�v�-U��MU��wWo �jG�}%�s�\I7��� ���z����Ѧ��	��@�����������M�ɴ�q���X�O�#ID������YM�}c�3z��3���%�kI!:~��Z����{��n�.73��Ů��'*��:m�t����v�laÁ���#�6��u�ٮ��{MnӘ]�u��Z�c2�s5p,9���`�tpt�V8`����+��ln���n��v���-��;�L�йE�
; �%���i9��Ax��	�`��-jț��NĎu�<��%h8�<��l�͹�d�D��N�<�wS�ƎS[�Wuv�6.���|����w{��;�?�.��mm�ba�[��r�v��%�\�v�C�k�����k�҂k�	!�^w��z�hIp�K�I$�������W�tݔʻ����ˆ{��I����ٷ����u�����f�G���5EZ)	4���{�SO~K�u��e0����T��BeQa�$�vd0�Ϛ�=�)�{�S@��%Ɖ6h��Uf�ݹO ԗ������e4���9#l�1�!<=��r�^�gc1up�Kl�:D�iu���{Z�.&�A��h���=�)�{�S��$��8���o���~Ez��5V���UoW	4��
�I%	��7��r��e�=�$���Ϳtډ@)��?��zV����e4��h^ISD$�
	1�Hh/q%Ro�S�7}~0�.�\0�e�9�ƣƇ�Hց�e4�fu���ݽ0���x�Q�0vn�98�vi}��:1��s��G�k�h���=��$`�q'\3�:���M�6��߷���.�v�?s��vm�|�t55v�
j�B��,ޮ/�i�n�_LY�����?0�oL��q%�Q=��RwmU�-�C�0	=~��}ڑ��9G-T5	���{~�uq`n�q`jފ�''x��8�q�����}��-�|hv\0=���m<�����ꕎ����ˆ��M�������;*G�o�����w�dׇh�ϰ��1��Բ��m�'eG<wK6Pc�B91b`Vݶē�9X�v~nޘ�K��ʑ�%���>4~�/��X($ǎHh�ek?�qs��mn�M�0�p����POG�tݔ�Wwt��{� �YM���<�,Z��T8�8�Yn�����IV������ �;r݇7�@ԦjM��$�S���X�t"j�Z(�E��ـvK��/$�������y���E:��;�wJ4��qw4���Y�ge+�g�3�W�м8�j$�$ǉō�D������b�;*G�Nˆ�s�_�M�� �k�Tjq7����G"�:�V�z�hl��v��\K����:���W���R���][�=��d�a����{o �[� ��� t��bف�㛹����xeH�<����x�T�ڱ	�
4��I��Š}��K����?��׼��\0�s�7�x�n�~��ls��g��-�ۑ2�@jG[U����8�Ө�F/kac*�r�Ɖѓs�Lj�d�wl�;��v�z$zL�z�1	�n��b�<d�'��o{tn��mOFl6S�[tpg��4]���z@ܼuj�P�؆��Rʙu��vv�\�4����\�;��ϳ�q����F��/��Ù�R�tj��s��Y4��q��C7j�[k�Y�w�}��{�����������w���v9�Or:���;d���vtu��f�9�vs���L�鄦o��&�*�0�w�;g�,ޮ?6�k�=�Ϣ�/̧�qb�F8E�@��y�M�0�^��>�#�s���l�\>�$Ƀ$���o��@����qq.���l�� �t��:����-�!ՙ��l���wku����Ĺ�&�Zm��un�UR������=�ՠ^��u��<�,Zޙ������N�\����`;��k��f وv9ʔvO,�9�S�o��������"��n8�����;�����b�=�ՠy�����`�4�)���5iE-T�1KBP�$D0X~DJ;:�T�_��mn�v\3�&϶6�c�hv7CWwf���xҤxyq$�ߧƁo��@=��b�~Q�&�"�<�R<v\0�\0=�ys���zށ���bq��8�
5"�/YM˜�Rni��^��>�#�"�liȲ�]�G"�Վ��V���W��ZeV�v$ݴ�Kz�'5j���_�ww8���η���9�o��@���h�j�/[��{x�7x�L"o�yzX��߿&wku�7q{��I���b�][��2)$�@����z��;3=XfQ:���@�0
:7Sv�J�����0�� $�ե��'���J�Q�f�� P�:?� ��*������ǕB'��ʴ��{�I��	��]��(���{R$�$�bp@�Bi#���1�$b�C0I$Mq���a?L������@z�JmJ~C���"�?
� �q6C����U +�x| �sC�ҩ��|���3og���Šx��WF�5�7v�U���W���`�~0ӷ-�޻���L Q�ыF	��/�p�=��.s��޷��������V��=��۹6SY8�'����ݻ�z���|���z��r��҅��$q��=]������O�1`I1y$�0���@:����?(�C�I�}빿���gww������o<��dڌ�V�dk�6��߾��/�)�y�-��s@����2cP��D�h|�J>޿�7�����޵`�tĚ[�nS�����M�9��t�n�d�D�	�@�h޻�I1`��ǀ{�K�Xn�!U��ݡ�W&;%��X�H�*���lh���ct�;X4:W�#����w�۝�v'�Q��~��4��hz��βŠz�Qv���[uV��1f�s��l��5�M���~��y&���� wM�i��AJ�͞�,oWTY���J#7��`M�ŀ}ލ�hRi�7E]����Mͷ�}ٸ��1`o<�\\Uٛ���!�H���ME$Z��Z�6�}���7�������Г[�؞��pc~���.�xq\V�C��؈]�a�Ų�}M�rWcC�;E]9�<�q��9N:z�C�c����F�^ܛvn�y�Wtizm#��dۘ���v96�m�s�x,��-�֠v�M�d̒ɥ���Wr�ZC�҇v�������(L��vyݐ�m����V��x����m3`C���m�^��t��TЋ&$wi륶�������C<�Ζ�w�x��-՞��qr������>�^mt��v�*��[5�3^zQ��{���>|�dc�s'b���ov��>�H��.[�_�vV��=��>��L��&(p�=�j�=�.��Y>�{�rN���ߕU�DW2w�/ʕU��Wh�T:�x�_��v�x�������5���*6��n�;.��ݼs��9�6��M�� ��#�=�,Z��`��bd��-�f,x����{���{o ��#�?Cx�������[��]��zZ��#I&Sy��������Y&��)���t�Wj��me*�`v�xݗ-�v�~\��l�X��)��&�b�&9$�@���o��<��J��X�� �s��]��}���;V�[S�I�Llr;�xݗ���8�en��o���rc�8�
Q�@��恛=�`guuE�ɶ�7��1G/�ΦLj ���y������/ ��ۚ�w4y��b�p&%$18�sAG\u�۵]��Y@�.z"۬��v5�c�&4��48�$�&	ȴm�-�z�hvb�\��v���ث]U7lt��I$Z����-빠y��m�<��6u�IAZS�l�n���X��V�w���PД(���7�Հ{$� �S��ULN���?�s^���x�1`y$�f�X݉����;m�Uwv���o ߻��~vn,����K�r.�ҫ��e
�:�Uvu��9S��[$'�n���!n�ؗrkgE�կ���}��G��(ԑz_��4z�hz�����}}��6�x(F��`vb��gݩ� ݩ����Ş�I���ռ�V��i�c���}ښ�	+�<=��ݛ� ݛ� ��v�$�,x��@��Šy�S@��擠t��3DM�!.�`�5p���S�<�/o;���<}>�3�3-՗wuV����{�[�/�vT׀I�t��
|{�=r��L0��j\2�7Y�/D�ft�=�w=���Y���<ì�ӳdP�e]ӻ?�7�k��Wbz�����_� �ր*�;)5T��`v�%v'�~�`vbȒ�r�����m�����@���{s@��|�����"9<Hnb�?v\0�LXݮǁ�NK���g�,x��������}V��;�,oW4�T$�Ѽ�����S��t/4���mmt�Od�HIn��xZ�ڼݳS/E��[B,�Vh�R���3��s����0����D��m͋nz�v��'�ku�L#�]�����zs�psH ��8k�i�<���/I�'L�%=:��Y�����DKʅ����wmìv�p	�<���]V@�qG��Z8�z�v�@=�k��Y6�K;K���0�ַDC���n.����|�������v��1cO9j����;��v�اS�q�糳�O1��b�s�&Lj#M̠{]�hϮ-β��������8�,�"M	ȴ����YM�n��k�縼��:��/:e[)U����O ���`�����}�5�T�����B�*tX��;�R�9]���h����;�\Z�e4��``�%�C��{Ϫ�;�\Z�e4-���ʁeX�Hي���y܏�i�Ɣ������bV� ��K�}��>����|��mF��$�x���@󬦁�s@��U��[�I27<i��ޮ/Pkv�m:���Z�3����uǠ^�B8�9x8Fㆁ��k������U`M�0ɩӶjh�n������7�j�
�����5��V���~�b�$��J���U�U]�����q$��$�;����;�{�k����Ǯ��vUi�y뛡7>r�V.�ݚz�7NZ�ck�o��WJ񧞄�1Q7?�o�����<��h��]����`��T�ݺwf�I�=��.q����<W�c�<�)�y��S�ō��Ұ3gz,��Se5i$��?�jj@�Pc��!T��>���7��4"C�SC��
�w����4��J��И�-�uǠy�S@�۹�^���������<�#s�m����wͷ����{�����{}~0��*�/��I$��Ӵ��j�����HӤ�rό����;R;e�V����i��$%6�26a�3��X�\X���m%���� �=�j�ա�V��N��;.�<���j�fޘ�&,�.q6wwL�O�����@�߱����عė�wq`6��>�t�T��n�TBH����S@�۹�^����� �r V ���+��|��=��`�x� �MHhY1`��u��V;.�}��ӿ{�=�p��c|m��Ӥ�creL�Ǥ�eo����pkW[�.K<r����m�m�G;`����%��7f��$���6��5E+�� �Kkf��ͽ0	;1`���9��Cv���wʹŉ4�=����-빠^��W�=�����D�`������7��6m�G;`j��o�x�:����+V�mZvX�`��G;�lޮ,��V�V��CmS^L#�Hl��Ɓ�~����d�²��O�!A�-����Ke4�2"��~CBD��$ӈF(C𸹎hТ�F(4��Z@	����<A	�h	�;D&�9�F��WK���H�Phh�N��(�["�jHA�|Px�ZC����fg�d-�鱶ͻ`��I�����m�z��6݀�6���vY�;JXӒ�L�G�ڕt;08�n��-�،�H�䶕Px��6�+���h�V�].U�j��;v�����:In��J�^�I:�$��w]���)ݨ6ے�YVn�ڹ[.�$�jV厈⎻.�$@��%�e���am�� �tON\�����f8;	���EN��GD��wċiݲt4������u�m��#�90s�c4�pd4U�0H4Hl-�cu�<<��'g�����H3�K7X�6R����i�6�[O #v��*c��uӱ��ct�.�%�.������-�l�p�+E���p��J�0�Z�ծ��ֶ�6h7�D'�̝"�����X2W�n��:	�\N���C.x[g=gѣy�7/8��rb8���={u[��"PupgMΏ��.ZF�Y.U�tn�%��֐¶�vK�����6��
t�ͤ��h�l�i��fǗ:@�g�ֹ9�8N��7��R9� 	�n�����nH�����-v��-ó���\K�fp�e^��/#u�ћZfL�������;�w#����WB�3t�]�\Mke�wg���-�E�.�t�/E�ar�d�N��) ��8�h[[l��).�5^вRl��nؐIk-�䤗�K��meKy����s^�Hm��˹rAmi6��L�,�7m��GL�D��[��9�d����9�lpl��\%v;+�q%u�̗iۃ4[�a����U�6]��A�6��^cMJ���8�dJ%^��<�N5�
��)W�.�h���#mr{`D�Dƕm�4��A�6�]���;���ݳ��M��G�.�vϟ��vxj3&��X�kf�Z�kn��T�=���%���ƺ3��N�L�=�ˀ��
G��#l=a'��\KT�:W0g��'c@]pt귒M{V�J�U�6e�����5Ыm\8k�٫�,W:_S��I2��]2k�ѭ��"��#7Ii�H/����O�lqi�Q�������_�?"�"�k$D� v~4�!+ށߟ������s�&�g�i���޽[���+	^������,.�K�:�۲�q7dל�m��tv��A���z�í�/:�)�˷f���0ю7�X݆��vy��=��q�`�w��t��s��t�r˗0e��!��ՙmt��a��vL������ڌj9ڀ�x4�Q�E0�v�P9����sg�|t��ay�d��	�.��ҝ����w}���䩣F��얍:vr�׭y��Q���hB���{vM�h_8s)�O$;�^�l��`�#�$���s��������}s��&���B8����ՠIً ��9ث7��g�Amj��"qŠ}��s@�e4
�\z�j�;޻��)��xch����\\Of���� ���IV�ߖm_&�D�cI!�Uz��=Ų�_�7f��'e� �)�(T-�v�n2�j��W��<���v�,��9�wlnƁ���wv���>Z����7?����'f,v\=��~a�f��'~�d�D��P���o]��?c�3�I'�ݥ���ե����l����3�����j��N�U�woL;��k�h���=��񱨱��"o�Uz��/;V�o]��b��������Ơ��9�=���.$��ߗ�n�� �v*�7�wc�E�M[WeH+�םq�"i�NF`Wf5��Tv�����r��?������Eݺ�����;.s�V;R-����G�6�M��/YM9ث ��'f,�� ��M�tQJ���5��X�H�qs�q.E��$�8`}�K���$MD� D� �7@t��5h���VoW�G(�*�U��&��V���8������׀n�ŀI.���z��U�I�~WWwAEƁIp�-빠[e4
�\z�S@�ȏy&	�D����]�)lI��	e�+�T��i
{sG�����]5j���Z��ޘs�V$�y$�0ݛ� ݅Ҫ)�T�UۺM՘s�Vof�ޘ��X���d��Q���PI�)�=ﾟ�qa�.s��ݽ0{5V���(*"��"jC@���m��*��z\ӴܷI��oR�H�R�-���[e4
�\z�S@���ͷ����w��Rm��n�5�f�2Ο��N�7��9���2�$��ͺ,�Kv�vj�Uwg�5��X��Iً���n��G��[V튮�M]Suj�	%� ��ŀI.\�U��s��Uz��l
*郻�uf��b�=�����\�8�n=�� ��� �
��t�V��n����w4�#٪�	*G���[��� ���UA^4v�uf�;`��Kv�_�&�ŀI.I�|BP}���)�zMJ��ԍ�4�۬���"/\䱋^ۗEK��������y1O����ֵ�s�XD�iۀˉ1��n1�Z-���[]<n��!��73�Wo.뗛t2�U�<��L��w]n6x�M�^8�	+�l��k�[f���a"E��,�+�$���d�#�id�7q�Ȇu�$���0�"j��]l�mۮu�N\����rY�����]�f�.�����w��:��ۛh�v�������)�{s�"]��\��.���r�C�G#� �DN5���c����vvb�$��/�#٪��趂�X� �N8��w4l����ǠZ�Z�ٔ�%0y�173@�ns�V��׀n�ŀw�q��j��R��0�b��M�+u��q`y��� �^��nت��!USnc�/;V�o]����*�q���w󿿸>=���{q�ӻ7c��m�}X^�î������L뻍���5�P�вM3X;�n��vn,v\0�b�s����@����JD�dj�s4�Sm&4�7�)Mĝ�����tX�ִx��r&�NW�=v�xyy$����,���w�t�8��%!Ǡ^v�޻��)�Uz��<Y�W�����H�qhvb�7�\�ٹ��5��X�H��ݿ�~�{q�e�笣�W���E3!1��u^N.n|���g�@�n��ܡ����)�Uz��/;V�o]���J�CY�I���fb��%Ī�m{� ��ذ	�p�:�W#K��lm�1���@���m0&�P�O����C�W9¶���7U`�[�Wtt���woˉ$��f�Xͽ0�b��hQ���<X�M��/YM���yڴz�h�5q,]��5���f���y������(����wc@�vp,}����v-<�>��@�p����z�j�-빠^��{�Q��%����c�/;V��1��ɿ}J����� ��5��z�(wx6AH�qh��ۚ�)�U�q���@�לa�LX��F6�ho��8��o�x�<��V;R<	�s�7��k�ww=�`nit"&!TIH�I�z��/;V�}빠^����w{������l}97���c$�#���J��I2X麻F3&s[��#��"�����{��-ŭ�,rF�����?��_z�h���g�>]~Ǡ^�/�`9m)N-��s@�e4
��@��y�.$�>�V���i�e�Uk ����*��=�h޻��G��U�~�@N^�Ǡ^v���V�=��`���0ڶ�n���Rc�/;V�}빠^��^�Ǡ=��w�{�ۀ?n�`M�vm<b�$s�۵ۦ�j����u�$ݻY����I�W^;Xh�֬���A� sٽ�=ȓ�sK�m�W.��pjge���b�Zw.�Ӂ-���e���n��)�Q�ط�8Yb�n��y�8	g��]�n�fm�Cn?��n~�w��,��lh���/i5ĝ]��u�#Ϯ�zr�1�&���CL�q.��3vC�۳[�o2�W9��8��;�{������'����9����s<�=Q	w��y[���8�ژ�G��/�����<M�R'^��]����*�q�.s���en���Н��!լv\0�"�v�x옳��..6IoD:m[���Wwf�n��'jG��s���.r���b�=��;ԫsǒ(���Nc�/;V�z�����*�q��;� $���uo ����{�$�����<��U�^v� �ӕĂ<O�Hɘ�x��Mx���ېn(�l�x���ي��gn��8��Bs4��hu���ՠ^�s@���<j�kț�8hwzf����NC
�?��E@���\������I��	�p�$��d���:6�Ɲ;V[�O �[� ��{6��&��x�Β�qS��۫�x�s�������=�_�J�<�j�<�2��(���$�hˆ����	*G�w�b�<��E���q�J�,G�N,��^y���7R�x��7<���a���X�{����{�!���Z�ՠw[��^���v*�Ʊ�<1�$�h����n,v\0�We�o8�'vۭWm��m��i�h~�s@�e4X\��c��kX,�\���<�քؑ���� �u*����!�١�$�Z
�,�-Cx~�Nh��!w��,�@�&�j@��[��N<��9k��a��4��JbAb�7���yt�ĺF1w�TƐp��3`~��|���R��ۇ�0x�3vXXDa�Х�)��]�j5���C��_�#�����N�{aPih0�!�O�( �G�&���~�������?}S`gu|_�gȚ��ő�HLI��/�O��_X��p��f��n��U��W
�vМ4=}c�:�M޷s@�e4�����}�P�˧��帄�crng)�m�.�fc�9�dG 67��x��byz���;V���~nޘݓ�.�y,��W��z/���cOd��޷s@�e4=}c�=�)�y�L@xbhs4z�h{�ŧߓ��� ��ŞM�ٮ��t��CeEUM��TX�WŁ��j��H���@��܃����f����֭5J��B��uv��.y�%7���7�� ��n[��A��t�W�ݻ�`m�;�ęM�d��;I.�ǜ�K�8�v �$h$�����޷s@�����,Z�e4.��ő�HLJ�`v\3�\�;6�o ����>옳ؑ��x�?���HF����Y�Zu��=�w4m��-(�����N��wuv�=�'&�f�,�.����/O�خ4�<q)�4zLX���ٹ��>�M��'e� �H�A_�?�1PƉ�� ���w��{�߻p�߾v�O(�>��a�^.��3Ҙx��p�a�9Ry_�\,o1�S���W����S	7Eٷ�,���H��xE�n,l�ڎZ��l�o�͕D���[�����h�ST�	�SwDˬ�Y٫L�ɬ�D�\>���;X� �]&��m:lU�:*��؞I�s$K��':�;W �g=��Μ��0h�ݸF撞y둫�b���$A��"y1B��d�)�JM3Z����~tp|�u�q���:n�]c$�=�'nwX5j��b�7t�T����o�~0�We���$�������X�:M[�!���<��M�e4=�s@�s@���IX���'�e0�I�K��ɻ� ���0���ǆIM&�4=�s@�s@�ӥ4m��:���cY1�I�`옰��;�?��� �K�����2t���u�f�cp�(ݟUu����9g�q�=������ѧ��8wf�A��,�����w���������X�h�R�t�[���	���f��:�M;�Q���nh�}_��Z�3I�у�����&'!�{l���n�߸�ě�+u�ݽ0�-A�E;�*�2��^K���}�4���>��{l���=_�idLHc�$4�Z��hl���e4s�S����loW:�Q�j�Ugr��y(��9�{'gmۛ�9/�����Bs�GegWO�ښ���0�.I../�$�|ց��_c�L1���"jE�u�L�$���ݽ0	6����Ǜ个�����jڡ��m�ـl���;+�����Q�DO肔���!lm7��L��X~��X�T��=0�p�"LI�@����=���:�����M�QG�����D�-���)�4��ޘev'�y$���ӳ�UݣW`��[5Ő���m2UƑ�B���[I�m��tv�
v��އ���t�^~��@�l����Š{_U�~�Z�t�wHULe]�~��s�F����վxgn����+-�j&$1��߱h_U�u�M�Jh.�)$m0R5��)��~\K�\��o����vv။�$�%��)b�`�#P+�4Oi voȁ�6<�߽.䟻�_c�L24��5"�:�����/�~<���ZW�h;�X��2LJ����ez�G,��q�ы���;&�=��ۉZ/�Ձ&��1���<�gƁ��-���)�w�G��U`�r$Ĝ4��h��hzS@�l���)Ʋ�����"�Z��xgny$�^\��m��7�� ��~���<O$Rc�-�JhzS@����6����Ң�B�c*��;;p�<�6�G�{6������夤I�N�#�B��D���d1�<�4)�F���tv�����vzضW,�\��'T��"ZZ&�M+ؕx�l�ی����o�k<n��[�=b���5�D��Hй��]�'\�Y��7d�uG�l���z��K�Ut��mm�5�����������3r�ǰ�t�]�^)�1X6l��+���U�K�i�컝��f����S�bC��:c{����w^������l]����H�e���z]oRY/i�����污�;�H���C����꘮���J���?�[���-��_��/M\_�n�� �ɣ���P;�i�P���#�����Tn�ذ{o��v��ą��LY	IH�#�;���-�M��ŠUz�ˀ��J�d���ޔ�=��ZW��/UI���7�L��b)v��h�n-�����h����=��Oݭ��8��M���������H�!����!ݲYŜpp�����p�I��
�W�w[��[ҟfx��}�@�S�͋�kh�8�q���o��.���f[��S�#���l��kD+�U�N�۫X�oL�R'����&�&�,��i]S�1�R��0<�v� �&��ɋ��__��@�߅$Jc#X�b�Z]�X{&,}.һ�j��A�}(��nz:��ێi�
ݕz��׈�U��Κۚ����ۧF��﻾�}~�đשe���n�ذ	��`J����}���g���&H	��-� v�������y.6n�2ӤU���۠ufݩ��#���x�p�!��P �@�
�H���Ȣ�<Q	�{����w�|hJFز��X��$Wc��s���LX�\0=�y$��{7��:��Uʝ:t��WX{&f�}�����Wuz�;a�͎D�q�f���ɣ)	���nў����W>NG�g�@�n���a0�6߿����=���
���;���<�^���"������]��.y..%Ty����{>��l�MݗE]�N���>V���w4��=���}�\��$x�$�C�3�g�V������_t�aO���4����g1$����_�ެ�J���:��d����e4k�-����w�m�?����~�&
��3a-p��S���{n���D��K8w)��T�8�:-\=�vx9bN���W�^��n�߿g8���z`M.����]v�ŠU�W�w[��޳@����<^��b��M5q���;����Y��q.7ݩ��5�m`����uB��Вs4�Y�{_Qh{k�=��h[^���"6���$�s�-9�X�LX'e�~�/��\��#>�����#av�H���H�"��XաdJZʈ��qE�8�^��T����F)�����e�]�RA�`n�A�#�y� �Àh
@�R,�i���F��� ��I�j�	Mq���"|�M9����s�~����?Z�d	�����?�+�`WO��"Ȃ � ����w��;�����������@�f� $�����շ���'@�� �6�鰖f�-$y���-���A^�X��c9����,뤉�[34�U6n��8�&�c3WC�ac��]E��e�x5�/,�i�<:�$�r��f����l��DY���hv���i29��,���u"�Mď;',����ݘD�)� ;S���7`�M�"����!�M�t�t�7�DV]z���m6�Տ�ƜrJ���;Z2�ő��M�wç�M�;J�˛B	���kv�����mq��q��R�C��B�5�׭�H]�Xm���[q@���&�r�7R#l�A��,�^t�K�̈ǧM��;=����T��+��;s�3�e�l�ms�w[z��e��/vMm���d��n�ܯ���7iCi��Hv����+�(2�0�d�V\ӡ�c�c��:a�m���Z,m�s�U:Ӭ�M�n���nl�����ˆ�[��.�|l�U�G^��Ƶ�Xζtͤn�(�m�rҬnr;;���v��]���'n�wl�`�td��@\=��>=����K+��� r�<08z\�n����kկi�uҔ�z��z��m�3dH�h$h�Yl��Y�l��{]e3,���T����,t+U\�V�B�Z��� �n@.�ˬ�	�#�I��m��Ke$�Z�����I�bU�$ڦ��gh��u��!z��m��sE-�H-g&���G��K�m�V��Q��Rm��Rqg si!۶-^�m�.�)O,�86N���ԩj�k��Wki&��Cmx�H�Y-��u��m��M��L�m�hC�j�"�L��ph�*%���훲g��u����;�J1��F�1�&��Y�c���lnn�R7����m��Z�j�n�U�I���� �z�\��<0��&���8�3����[=�Kd��5F�m�K%&�/WJ ��Ȅ�7]��� �y+;���9EU#�Y4in�S�e��'s�:�b�n�*iZ��b#�--���J��66�$[N��.[�ۣR�j$QN�+�E_� ��("�4��1AH�^:D(q���ҝ D���򿆁��j Ҫa��P?��/nSvXl�O2�z���b��^�<ܓ��a���E�}f��������-�R�\I� 9�:��1�-���ǁ�#��L�m�$]:u�NE��6ь�u��v�D�7f��nm���`_j6����p�ƻ+)����� vrm͇nājxk:�ph8t��6��� 
��7�W����:ݙN��[Z�n8yGh8�؎t��]�~����{����?;c��O����a�H]GE�H�ۋ��sQ�ಂ���zȵ͙�����ϣ�L�lR�W=�n�[�hϨ���a`2G�A��m��	;p�;�����^\UG�^�����VZj�7V�{o���`��Is��{6���,N�-:UtӠ���4��ZW��=��hfb������gѤq�E �
�e`K���~v^������4x̟���N��u;���s=�9�J%�v�v�R�:�["ɬ[���U5[��Ȉ���@�۹�_l�����@����JU.�whC��X�\1���=C��٣��b��޳��rO_��ܓ�&,��8�l�f�4��Sm�J���-w�hwW�{m��/�S@��#��`��b�Z~���w�}��_l�����@������IH�#�=��h����ˆ�U����������ŝ�l�[�L��kŁiW[m�2�smki��<�b�s�g3���Iݦ��'nd��9�[�~a6ύ���Ok"PI�@���Ēl�&�6^��\3Sf���gѤq�(��ߞ�ץ4�O�5G��C� ��ߵ��'��x����	�*t�Ӳ�������sfi�n�� ���`���?J]�Q��B0*��$�� Ԓ��ٚ��|��=�Jh.r
0�R6�(']Ywu[��*��B�˹��NC�ѧ�.���&�Y�?��ǒHhz\4
�W�u�Mޔ�*�� ��n�Z0�ef�q&��z`���$�h��H�D�$�����'ny���O ׳k �⤶�2�Wn�]�Wf�����fi�G��X��w7&�C� ��@�,� �El?��D)�y?�s�X�za�w��*�i�U�v��9{n=���ޔ�-�M祊���M�$�L�vŎ͝����nԵ�*��p�oS��WH����3��d�*�^���Mޔ��ܚ���خ4�MA��@����bG�Y� N��#���~���:�]R�Wf'n�د�M�ٵ�M��@��z���$1�׮M���zS@��4
��FF3 ��ۙ4
�W�_��x�Y�'����$�!�P�X�d�l��>u����Jɏ��|7ɝ)��DOK�=T�9��z`��rk�%�
�dڐJm^�g9gKa)ӯNC��1n�5���ɸ����d�[mݤ��h��.�ۉi��v3���=�<�FNb1�����u7{۴�s��j�h��B������{6���{r�8x�aĞ;�4�Fܼ-��k[]�3��u�ک=i;K�2��γ�n�!35T�*����=I7���'�R�s�zڮ�_Y��8�F�̇0�ܵ����Q���t�gJ�f�hk֖��~�?�����`gb��ı�s��?��Oa��Ɔ�H�919����rh^�@�қ�G�_���8�&D�' �_�h^�@�Қ���/�lt� q�"�&�U����`Wc�Ը��U��+�:�xN���M5$N=�Jh��@:�ɠUz� ��YE���&�����h�q��\�n9Y�"[��zCdiܭlY4t�o'H'6��4�����@:�ɠU��u�M�k՘��F�!�$����WM�I��\�벣��3�Jh[T��fA���2h�%`��a���/L �5^ߥ�mH�D�bR!��?���Ɓ���@:�ɠx�����X����&',�>vV�9�U�����;;p�?~����Y����\��ٽ��/^-]��=m�3����g<��WQ�x�\<�óiLNG�z��<^���)����XU7ՀzҪ�v�0�����x��@�Қ�ޯ@:�ɠz�)��Wi���Ǡu�M��W�~�����gs|��DƄ0�]$�J�n����*�:7~��+F(��T�:`Uف��]�X6j���J��3L�ݬi;�M4����� u�@�{k�:�������<젯;�]��V�)��I�S�j���x�#������𝝷nl9,d���ݞ��U�<��|��)�z����\���8�c�ĤC��zS�9u�����@�{k�/�:�,hid�c�N����e`gb�<�>��6_Ɓ{��k�'#�����o�X��`f�qa)�j�Hc����V�2�m�a
Z�KRI��ɰ=ƕ2�8��B��&j\�@�{k�=��=^�z�e�@�����}ߦx>�h���f&����D����Y�v��b˔۝ƍ��������&�M4�����������W�^��x���s�`	Ս�Вs4W�^�zˆ���נ^�s@���f(��X�q��zˆ���ק߳1/��nh���]�E#I�,�bX�Z0��+ ������=��=����b��'
DI�z��#7�����X��6�_Y�����}�;���ɻ�%��x#�:�ϙ���6�^��]lyx]�V�b��.�pi1GJ:�]a͐.D#�V�v���;�[�����
��\��l��j^�����dܘ��:��D���$�4�m-��1cٙc�ʦK�h�m/Y�Vd[F�mX��kf�B�,�-�J�v��2sFH�UF�3�fz8�ܢAjw<$��K���۲F*�TN��7\�v�b��xS��/�����_�.���CZ j�빽\/��\��NrPyv+S�8�ɗ�qkgH�d1�1`�Lrs8W����/Yp�<^����h��1�Ʊ0v[���	�q��>}ݬf�,��eg���l&�T�=-�7Vʫ��`>��;&,��e`��0���S��n����U����n�X_f�;.#S���XҖ��tU*�mլ��e`I.l��~����'dŀZ�8����?�Q���ӻL��˷Z���
g���������|�H����c��ڎ�L�q>#X�4�>���a ��s�;�d�����RN4��%�9�����7�@j�� �̓���ݮǀNˈ�%��q*�۶�mݰU��v˻���b�>��;.�x�W�w�5��n����}V�zˆ��^����ަ�x�"�܋@�e�@�3?g���	����]� ��Uh�wk]�	G=q���蔎�s���a�qĽۘqgF4��5�bN6�Ra�x�W�u�s@�U�^��{��1<j�LM�ND��/[��<��h��h>�Vj�l�iA ��u@��uk Ξ�,ޮE��P[��B�4�ܛ�q�8�d����B'�4����`0!~�[���2IH�XHI���B<'�#)߿�"��8�����0&�����I1������4���9�6B@.��7���0d�`���b�# ~���M��H��h ��{ �a�<xp�q9��	��_nYӌ8�b�6d�J�+0��`h�`���E��b~���D��d������B�j��$H�@���"J@��S���}�~V��'H��+I+䎗ȶ�X��b. ��#�2�d���+$� �=�H���� ���gԐ��H�5v � ć�@��=O���f����)�?*�aT tY�s�
i�� ��'" HL�� Gm�&�ߟʦ/^����˯��ߘvo�`l�Ɠ��t�N�U����s�f� �ɵ�Nɋx���5�{5�U�:hj�P�n�����=�s���~�S^�ˈ�>�(���HOV��I�۝��Dx�c�h�Y�,D�&�N6g�N���$R$�A��IH�#�=��h�]� �e�{���X�U��
T�p�I9�����ˆ���@�I�7��9�ٻ4�T��h��-�v�~�a�wY�{m��<��h��o�PI9�� ���n��,����ܝ?HHaV�J� #$�IH"b`H�Z�A1�����2(�2>7ZE�, ��Pҡ��?�d�}��4�����dq94m������ˆ�y�f����q��q��ɨwl�u�pY�$f׈�����v+��	��'#�s>J]s�l:Sn��߀��� �e�`��{��ww��~]��I��Gͷ���~�����pm���xww����R��8��٥�]F�$�s �ߦ��s@�U�wYp�;�+q mD4���bI�w,�S^�ˈ���|*���~Qē��yϪ�;��h��^���#����4���v})Թ"o&�]�j�lW�Mt�J����:l����d��5����ͬkd�}pUÛr��l��ȓ��n+'lXǓ[m���v��dV��F嫯b7Y��nCv3F���ng�2b鵇/[%��,:Z��vR��؟}lg]��;��Y����&u�t��������e{e�=T>qۗ����%Zr'��ܪ��Y��J�:�������߾������ ?�@�nF��&װ���6V��9��X�uӮ�/!�q�	1�dX2(����/�g���y�f�m����� �(���H$9����^�m��z���.�~H���	��	Ȝz��,�Wc�S{�z��k ��<���l�9�z���.��z��hu�fb���NI"�-��x�W�[n�޾�@�;�`�y���ڸt훐&:�[U�eW+Ԭ��Mq��\x�.�n˖�wc��+i�4��m��;��h�p�/tW"r ��$�c��۹�������!���?~��~�ޣ ��e`ފ���H�*��L����l�h+��۹�w�K�"��DcR-�.��z��hs��Ϗ��o�F�9� �[��-�s@�_U�[e�v�}�����N���L<>4j{6�p7��^�8z��0qVwp���z˒0�H'"q��}��޾�@�ˆ��^��\y�O.&�M�'3@�_U�[e�@�^�@��͹��^���E�&��E�[e�@�^�Oq��3D��qz�9��N��n,��׀u}!U�X�c���i�4��m��;��h�p�/tW"���IH�%`I� ��������`��V��������ད�1̢�Y��)��[k�o7 f�m�r�.2L�צ���"؋���hz���.�ޯ@������6D��ԋ@��U�x���	;1`}]�W?0"�h�Om�SX�M�Z�������=��Z����_�65P�� ��Ǡ[�r��N�Xӫ��M1�])4ږ�-�p�U57����t󞌙p�r��C�X﫱���ů�>ͬN���e��>g�F�ő7�$Ļ��q�YL��:}������X�8������
,14ܒ/ ��s�x���z�hz����M� X�16ۙ����X����Wc�$���R�$��	#�28	&���>����y����j-xϳk �*r�e�&X���y��l�h/z��w4{�\x�D��R-�.�7����`{'z,
m���4�k����v�ۭ�v�9���mL��wX�1��gf�۷M��q�|s���B]����ۜ��Kn݇�gqi�r���دe��i��\u�^���6;4��9熺�N��YB1ͣ��}��ݸ�ۦg�V4F�mcG�sA�o:<��E30��\�ӳ7
X�m��Ňn�\����:�;H�=��{A���ܹ�>�y� ���Y�3�l�ģ9�3�ܜL9�Ζ�������A�' �?d�.eֳS2kti��W�d�l�,�H$�ƫ7�m:����>W	����DcƜ���I��|��z��hz���.����M��)#q�}�ۚ���@�ˆ�����<��8�1���b	��<��Z��0ԓ>ͬww��+-'u�E�&��E�[e�@�{��۹�{����7�X�d�m�0�<����Ձ�;�`wur,�M'������j��ں���vު�N���K�e�Yk����+���r݈�i�U�U]~ww���x��7�����o ��?�H�7�,JD'3@���n��5�!��	 ��"��nh�T�ʥ傶�?~�_�`�~���h�;�Ǖ�	H�"�-��{�h۹�y�����Ɲ"�p��$�@<���-�s@���h�p�=���cWi6AG�@����_U�[e�@<�٠���;~��{=����|;�9�rz���%��8��5�w�t���;V���vs�	�������l�h��4m��<�׳1G��b�ӒH�l�h��4m��=��Ze��,@��bs3H�guX�֬��i,Bm�@�Nƀ��D8������I����p/���"F)�Orh۹�{��l�h��4.:�&�ą"��{��l�h��4m��<�eY�
&�<�#�jbqz��n����F��l<���u�iMF�F�m=�zvБ�ԋ@�ˆ�y�@����_U�LWˌ�RL4�m���e��=��Z�\4}yLlj�M$�
8ܚ��h���<J�7 ��f����i����	����M(ݮ�,���E�{;��m�-CKSisi;#�Ձ��Mˊ�T�-�.���w4}}Wͷ���v/;�]����N^g�*۵vʶ�M�=����GWnxN�{fÒܾKp��8���&�Na�{l�-�s@���h�p�;�n9&E�S&$�&��-�s~�����׀n��0�ݗ����W�]�w�c ��hu��\4��h۹�w���Xq䉧�~[�����k �LX�� ���Ҝ�U���]�?�+ {�.s�ww�����MI>�>��I�����U��U�EUj("��H������*��EU�A� �T!B1T#B�T"0T"��BT"B(T" AP����T"�B"�P��T"�T#BAP�	BDT$�@@�P�AP�B	B#P�AP�B$@T �P��P��UAP�	P�T!P�B0T ��@T"$	B"EP�P�AP�E�EBDED$ !E�DBAP�P�EB,�,�B,U��BB�T"AP�BB,��P�)B
�B
�EBB!P�@T$T� @��������� ������*�EUj("��U��PEW��A_�EU�U��PEW�"�*��A_��PVI��|!�AP��` �����[��       �         P�   >�x  } P� � *�RE   	 �@Q"(U��B   
 ��  	@`   ��P   �T]獵'��ɮ{;�[��}�io �*Y�l���ק�U����[� ����ͫ�s5�{^&.�ˡ^�� �¬[�K��F�sn{u*� �J�����\��ͩ�]�۫�o�  �T� (
 �,����'ݽm�uJũ{9=+�� ��z��mj��:�s�G���W��N� g��r���+�  �=[ru����&���� ����{���ݪ�9{o�k� ��    H�UV0(�JVm��e�� 
)(tt 2 h)@�� �  f R�     �  � D O@�� :n� �   �� q�J� �@U,0  	 =�������X��@�ո��^���ֻ��V�:U����m�o�v�Ź�O-�ɮ����w���O���;�׮�wm������ 4�}K�+�ˮ���m�f��)� �| P )J �R�}�+b�\�>���s��������R��{���ݼ��k׭�ʫ�=}�.���y�x yyoV��=��� w*b޴���W;K��OR��O{��������8��m˒�    ��7��J� h�H�mJR�  D��Rd�   =��I���1 �?�%�)J@  �h��)�@G�z�������4�����g��}>��b���J�
�����UPUqEO�������TX����������i�-$���q$�FI9��+.�f;05kI�`l�F��8oP�&�kZ����F��7_֢y����g0=N1�{s@�B��@�Aa35��x�>c�������ߜ$�2l�!t�<�'$�)CC�����6ƺ7#�6s �h6�(�$B1 �><��O��<���7�a=du!��
�A�]04n<�Ј@p�	�� �td���H���*h�!'9�a��$�)N� �HJ:6��(��Wi
q�х,aL6B��$�2!�Z��].le4B�z�ńa�t���3z���z�7>ގdu9�=SA����B�*�l"I�{�B@8
:S4�Sn�C��<`ň E�!$��0`�;��8�+*AZ1�H��a')��ٱ���B6F5"�t���$�40,��DMjHK�8R��c���kD3A.o�2qٳN�l�:�J�����ѐ� ��p �A�A��i�<1�BGG��3f��!	C�#d48m���4�
h�44,�j��������#�2XJ�`@��l�Ұ
&��}����Դ��`�"�H�V@�d���v��$����p�����3!N�$n�Co�D�CB���$`D��-)SA�HH>!�P�
	��ᧂE�#�B��uY[I%1��2І�nݴ�M�;YK��i�^]�XP�����j�I1���a!H�H��tTrBH�����rGqK ���椉�����4� q 2 	P��|v{��HRg���g��T��0"Ut��C��`į�����zH��Ct
}��n0a�.�XB��3u�P*@�0��xSAD��D �]$�.��g
x"lb%WF0*i@1�L���y|xqĐBW@�b�0�Ab�XMD-Sd`S�!$t��E� T�><&���1%4`�"M�	�! 4�l�1�M<6�>�|0���AR�XD
c)� 8�%X(T 5=�����F��ћ������&p"�|�v�~᨞_�0�ˡ�c<����`��i	��	��8I����OI�n��NM�Đ�Y�@�i�"� �U��_z�&��"B"R- �x���8�>>I �F(8�&ӏ�`�(Pӎ�'|����nG�	(k�7�t�I�Mnn0X�L�]I�{���0���@#�B��@�U4�"k^�N#*B�HP�E�!B	f��V�F�q4�I_4�Q��"B!C�0��~����`���jb�}���FMc��@�
ƺk�d7#,�����A�
i�`@������0�k���C>���|L�� @O�-@�Mnp�9�<�,ss8x�y^x��`���#�ӡ�4h&�f��%�
%��BH����P�"h�R���f��]���� `B%H1D��N:�M�SXBY�7��g��i`U�6��lױ�rY�p�~ ��r&�`@<|OIa�wm�%Eٛ �!d�X�%���"F+���l�1����ؐ�����?�~�d���lp���,B� FBᰇ�<��O ��1Z2EH��!u$K�MJi��.h��'��I�2Fyt:�d�*,�AR��i��.�Ǆ�
J0�a�WL!���d�:�Cp!�R�y7�՚u�2��P�� ��SX��,k
:�w͜%�+5�f��0𚄤^a)q"ՉOH��E8��A���C�2��фə��)%,�<�����5t�G4y��!�f�t@���ys�n�.���t��E�$w�4��f�]��i�`k�0�	���%xOOtB�F��Z0H!�b6d�H�7���6R*����� %!��*����T� �U`��9��	��F���!��%4C7�wYZ<�5�]�i�01�J���(��F)"F��/��ֶ���xp��!�B���44���L�Nl.��mK�]!@`D�T�ɀ��m�'&��_Ns�I��IYYp�$ ���۱�t���9xO#�l�aH^x<%'!Q�f�O��I�����=�m�1���|8��]a<ֶi��҉�@"@'��M����=���,Gф��sP�ᰄ	u��u��9���
�	)��t�8{��ᄐw&�Cc�ǎ����5����8�9�)��i��� P�x����=��kЅN݁���aCFx�]����WC¸m6��<�5���N����͛!��ڛ�7ɬ�"|��{'�#SB#%4��7�'�EN|��5�d2�HI�)�X1�ӣXEta�
hI$4�_R0"�NF8�
�(�)'9<�����RGD!����~2@���5�&�!���8c��l���Fʐ��{[Z��0�T�yMA�6\��M��,3FK��.��f�90̼�BkWӄ9NSlt�$�7]�ͤ+5���H�#�"�d�(D�hAJ� �I�F# E�d���dp�%��n�����'0��D���	)8_�˯������$~���<,�1����Q���ɷ|�!!#$����M%��Xx������,ӊ�b��79�Yr�� �yōB@"Xy�4���\�}����q^1Һ�_V>����ѢhĔԅ����_�7��/�f�`B�g3W٬"���9��FY�f��![*�i��	�2�)	
WC��Ps{�3�c�K��KsYÄl)�x���6�u��4�e��*F����XQѢ#�HG	F4��7i�"ɹs�hDR��G����4������P���\߷ܥ5ϟSN���n8_�WLn��K����#ur�Pв��`LH�Jw���<00CJ2&Hi)"�0�����$H�� �lVAbj$O�ߎ#�8z�:9��E�F���j�����磾Ml�$Lb�	�F_�Yu�s@s�J �`2H�7��~��(�	�,�E�=v>?$X��syK����g9x�u��<y���o{8
1��o��Mk��v�X���2�%/�_�xo�<����H1!���=۩��6�)����K�]�ϼ���zz�g�u���B�B��F	c=�o�CD&;9��H��B�`���6l�0�f�$�!u��a�0�6nJϵ9��&���s�������'б=9
�aV$!#��~!>�MX���<k<��y���9��rя��F���׳Sӊb@,X�����CI���˖4�B辔��	j�B"�
��F%q�M��Ů��;9u�ME1�!R�Қ�h9�%Ӹ�!%���Cr20BpĦ�h�I)�x2A��x��P4�q���>������� $-�     �[@    [@     @l       � m�  �   ��            �pm�8      �  	�  �  p � �c�   �  p   �M�-� ��m��  [CX�uͅ�����"̨�k5�m�e� ۖ���o��  [[l    �$�M���܌U�=���(��<���n�H�mj�ma���I[m&�n�ж�X`s�/��ڰshV��en^ݚU 
�Xi���k��$�q�a����-��jUP����[�n���G85���~�w��>�sK/�'D/Y7^�f�=��[cR�9ه���k�������m��CƳ��m�s<R���c�Z��Yy��r�ns��aŵ6�PlS��: lT��!��l� l�T�ҙq�\t�V8��4�nm-��Ij��d�r����;T��:�*J��rmAүu]=�L��Z^z�����P�e�^������i�������G 6͒�D��n��ۚ�j�t,�%lGRHt�8Z�@-��ڪ��%:]�)�"���X� 6˔^v������m�KQ��B%���l�n׮��  �p��m��/�m� l��� �8  ��[R 8;m�m�pX���5���x6�Ԇ�;t�K$�u�T�u�p.� -+f�[p�8G	l;C l�� ��n�YRp<��UR�p�@U�7
�mvH��m���b�v�   n�  8 !l��m�l�j��cacdՆ���� �!\�n�~)~�|Hk�X ��� H�8�['LZ�[R�$6�˄s�� �v	k[��6Z�t��� ԆN�������u�͛I� �z�@H�baڪM�޶Ӏ sm���U�,���m����}���.��` $�d���,��$�oH%�"j7m���l����5]G@�0��J� ��m��k�u�����/�]Tls��+�r�`�l �h,�e��n�Z����\Y}:���4�η�^)�\EBEnqN�gn�A�٨l�\����qۦ�$b@,3��H+H	7@Uvԫ�g`��M6í����^�l^�lH   �V �.j���n
�,n^k�t�4�V��v���[@9��2	 Im�"�  �W&���Cn*���Tm�,��  ��,l�wm�@ � )V� m��l�Fw�FҮ �}��� 	8	:N�ٶ6��` [K��qmm� �-���   �c]��L$>�}� �d�$at�ݰ�I�M&jC�� ��v��m��i�i p�-���m�    8 �'G$��� 	@� ��       �   ���   m�m�  �;m�ͫ`8 -�  @�`   8:[���@m�E��� -����M��i6 H�ֽg���6�m-� Am  �X���6��`l   R��ܪ�ت��`@5 �YEV�ʵԠ)��   �   ]��^ăm��A���t�l�m��­��Z2<�T�t  *�[zMo$�9E�`���m5Rp$�v�T�S�d����܉l��k��"Y�s�b֊n��q��8m�Z�j ��&��ŧRɈ1\.�@U��+�ٻkv���    ��Z���m[���� v�a�6� �  6Z؛`mۦ�f@�$<�v�M��x  tZ7mf` ��Jm��Ӏ�z��$N���m�� H� ��� �m��ٶ��B@��zʝy�V�����-�   ��n�Y��\�` �%I�]�  �N ��lZӉ$��m�[%m��v����۰lX��$	 �g	-�kz巅�h4�L� E��5pm�j� k�f�u&�m�j�`�6���h '@H  Uյ�Y�
����ʤ���t�eZ��y@m�E-�sm�� �]�lv۷� q�HnA������4�]� �mdE�]�հ6��  3o\ �!^�m'-]6��v��ٻm�amkv���6X:�-Tnn�SQۭd��  �l�ۄݮ 墛 ����llz)�WV�P�.��م�Z��Z�y����%]S];�K%��M�m� ��JZGk�b¾���mƊ�vÂG-���8kZ��
쪠�@� j<�*vniU��UP��9P��@J�'D����jgZ:�I�cm=0 F��smYj��2=�����F|���A�U6������&țq�B�0q�y�ٺ�+e�jۇ ��lS�p���ʻ�WUU���j�l�]6m�m���mmUm�f���̝E8���U�j��K��6b�yiY�����I�5[������pp�f�l�4R	5����y��m�ݤ� �)[��U����Y5�-�m�M����i��	p  �$-�4ڃ`�cD��m6��Ԭ�/lt��ԯ3j�lkV�Y)��� p� ���@-� �e��V�   $�m�   �l[Am����H7Y� ���� �Tu���&�d[@�^�m��`  p	^knW�����t�.` ��c�N> kE����m�������lmy��[Il  n�&��m�    
��ʵt�5U]t-�[v�-�^Wl ��h�m������vZ��ۢ�  ���@ �l�� 6�m� �i88�`�m���m�&�U�@@]t�tji��t��T@U�#�k��۵l�o���& � �m&o���EH�:�6˭�@KhF���lp�낖]�� ��Lv*��ضyVK#l�*���WJ��UU�n���`8�@MV�5�y$m(���꟪���M"+�ɚȯ5U���!�O/5�+����T�[����$p$�M&���)d)l]�  m�l��l�rmp��޶@  H ^���  `H��F�l�  m� ѵ���m��Em� 8$	ѷV�$�9�E�}���m� �� 6^)h8   u�          6ͰG]60�s�  ��  H�m�[  �m��` +��
�lj��n�  [@  �   B@L�@ [@lͶ�ڻ6�m�5Wa8�H�    	@9m6���mᢶ�H	-����--6  ��fٶ:������g�ͻ`I�H���V-���,�Kh [@���m����|    �2H  M+[R8����S�5[R����U�`� �n�[@H�kh�]�*۶��6�9�VԎm�^�Y;l� ݳvi&�$ ��kl�r@9 M-�lH@�g      m��l $[Ki֛  �۶�q!"BӪ�"�^W@Y]ڪ�]�$�SMv���VZm�@�m�J�,q��� m����  �kgJ� �g�m�� �\   '6��Gkkn� R���5��bB-�lʶ��;m�mQKm�� �:6��:تt*��j^�j�r�ת�Qkd(�9٪�nڥ�*�V3���+9V-��H�5�Ü�Ý��di"i{9 6Ȳ��$�Wi7bNސ6��� �e�I,ԚSl�8l�����f� �^� m-�Hm�9�� �p]Wv� ����(���  �m� 6�n@  JV���p�I    m�� l   Khm[  I&ձ [���Հm� �'1�Ͷ�N����`q�m�6�[@�6�l��� ��`[�	@ m:fm�[ ��`   �   ��v�   �3�d �u�� �  ��6�     �H2)$Ҷ�l��:M�l 6� �am�� � �:Ւ��5J�[J�eᗚ�-l+Ϋ��0qTڸ� ɵ�`6��Ͱ ��   [[l�  ڵ��m���&9��� @�I�UJ�,v1�Z��������B���_[\�ۓ��UX�s�I;5mI�U! ��W*�+j� �.�l� �l  $<h� Ŵ��!�   m� 8         ��mm�m � �kY�3$�f�EL?"�@P�1��c�O����ʜTE�.����g:q*8(T4��Gd|@x���QR(8���H��H�"�� ��D� ��c���q �,��>~ � "+����� q ���;8�Nz�P=�>�N*z*�l���D�@N:<�D<1��!P���O��
z�@�8z�}4K�1�z�8 8�����pS��Oh�������AX# HF@�E�W��6��b�I��#���P'�||��`A�*kʂGa�mt��T ��#�����C�>��A=� 
�U������.�����O�������	�P���~1	�3�[S��K�6�
�`!�8�D�h ��<@҂?}�`*���l�4_X��z�!�f�=uS�z<TW�� a��xK�� !S�����SPH�$H��b{��uUWj?�S� 1@b D"2�b�E"�V��Zj����`���l�$��  Ik��m�YE���HHcD�3ѵ�&,Lku�$ەݶ-�hL3�JY-�a�8'��S�����Qp�J�����R��$��qY;!�V�q�x�j��M �k\r�GZR�nY'aj��m��n���d�r���$���N�ɮ�GZ��rLͨ8s2\������Ct�ӂΨ;a| l:t�!�����le��vK�>=Gg�������Q�	^�yB�m�ܕ(5hd�&�����@�<kMe�FwX^[sM��m��i�\����*լ)�m�=�&� ͯ5��=��y���A���4�pX����U�8��v3�
�V(h=�7\/	"�1N�ӨsJÜ鞶�����SŁq�d�^�K�:�N�T֕UWB�t�*V�,��n���t됻,���aSɌ�f�\gR�m�vj�v"_mS�� ���g�/(��,T=Qs��U���ȼv}`ӫQ�T��HHn�=��Wbsl�1�[g�v�.4��9)��ʶ�^�9y煶��̝`�k���;]��T��E���)f%"049����/Hp� 'i�Z'��jG6ݡ�Rb1�-d�.ͰM@U\���J�)[%.���iۮݺ����i���Lqe�R{ɫ�ym�v�s�l�lgͻm� *ڱ�7k���jv�.:���L��vwh7-��ȼ@��i΄��l�m=Wdgm�6P����U�J�R�+�vJ��u�ڬʲ�lY2n1�%[]�U#��C�n��"��� ���[eB�����l��l�ѸĤ� hB I�R�s�g��zLV�@K5*�CT��/B�<H�w!ӡ��W/m�N+�����3�l̙���[��ԼK��@�@6P���e��4�UW@����U�hTVF����m�r��U]T�e�j�j�{`��=x��*��g��Tٞj@
V�p� ���l����m��m�����̹2a��Qꇨ���T邊�V�$�#�QȰC� �pG����EO�����/y˶i���\*j`��:��,�ӱt�on����88	���KA��C^�Yf���$u�-��$N�v�l�n�X�ʗ�l��©�hYRD�2��o��Uu����07u��v+���Ucq�ەn�.v��]v��s���s�i�!h��l�0�\�)���u�o$v2D�:�`ͼ��.f���X�f]PSn(���%ܺ�����Y<�=��ܜ�&��q�'q��~m�c���`�����/'�޸���V��i��Wo��0'������l��&���^,�
�P����:`M�t�9$�e˸Qw�+�R���Lݔ遽��rI�M����ŲL# ��2G2f����`�c�c�ꯔ�)��e�Փ$pn@cNf�ym������s@�빠x�?�+�1��1�q�]���yv����='�۬�֌�ks`�.,�JI�	8�(�������\��;��h���=��ps�s�pJLܓ�=�ٰ"��}M�QH���U��t�'d�$��6�%��fa�x�e�+)���� �ٌ�%�{Θu�74{�I����ƌ�L�	ݘ���we:`n�t��n.�O�QA4������e��s@�빠޳@�?b�|�I�2('��F�%�%��٨=l]ʗ���"��ΓA\�1�ճѓ(ہ��4�Ŋ93�=����w]� �z��n���-�a�qĬ������L{��:`rl�Z��Ѭs$q�ә��Y�s�ٹP�BH���(�F�TH��b'�Q�%�P��
>��ߖ,~׋ �Geɉ	8�(��������74����ùbnb$2H%&h�)�wc��ٌI0=U�o����G���"^펩0�ca�|��X�D�yc��#wN]�'L�\V������{-�뫓++�I<�ovc�GLM���|�Q�a�ёI���������74�A���QEi^c�GLM��-ݎ��f0=�W��X�Q����yz�������'�{�nO���U
�H-h����B���f�ｗy�L��]e�V^^VSwc��ٌI095�XDB�����5vM�蹹�k˳-�;k���j�8�Z������زqc�,��˕��̑�@CNg�_����s@���^��A�ذ���z�L�5ujm�1��#�&�t����ovc���u51$�4/\��;v:`ݘ��� �mi���.�*�VS�vr��f09$t��ٛ���n��0��%�I����%ww����ŀn�ŀ~Q	'	C��$*�Dj��*�  ��"+�"D�h����D,@ 4x������m]�oT���b�p7��������V��F*^]�ld67�u��6���n2<#��N�Mal���J� ��Mک.b�,<���K$���!�k�����)}�Г�s�v:3�R1٪�q��6�����lf�Z̞M�������R��۔��aj���%[�DkB�V�8G���㆑�v��C��Y�aŖ0RpZB��_Nv0�NL�v�Ʊ�׎���x��p�=q����V���,ϒ�$E���?=�LM�遻�� ���e�u>-�$i��G&h^���ٟ�-�nh���<��h�)d�1��0q��`n�t�7�1��#�$��&ףX�H��i����~��޿M}��� �[�9L�}������,E��`rH�� 遻�� �z���
#�?�C�1��#�x�m��7f��#v�����X��Y.�\��%��f��Y��;�xt����ovg��߾�s@=�~y��$�3@��~ٸ���Q'j�|�IC��]UZ���{Θ��H��.n��8Ĳ)3@;޳@�۹�ym74�A����5Yj�z���`w��遻�� �������I�8�M(��<���߲��tv{$���Ԩ����˘����M׭�lh=�yA�oku�@rgGlu�)v*_�) ����(��	�.����4�l�<�����Ѭs$�d�V�n�� 7�w�	)���� �����uz���VL(�"rh�{�nIϾ�lܢ� )���C����-�Ǡ���=�,�,O�d˵y���t��ݖ�7�1�rl��~�5�RA9�#�3@��W��Y�^�@��nh�)\#�w5�n�(�8��j���-�=m���J��PZ�b�g�7s[oTmD��~ w�1�rl�$������2�ˬJ�,U��^c �ُ���I��:`E���Y�bG|��>��7i���c���L]�l{�&�`N�K F(�q6HL���������׀�����D%P�R����ך��dn~q�$q�{�h���<���/z� �Q[1�Y#Pu����գ�7=��`|O���瓳�\�E˂��ں8hd�Ғ`�G&Iӓ�~�M�i��r������=��:����Ff�5���'>���ኤR(���v\�Հ�׀�w��5�*�$I̘�8ɚ.����4�l�<�ss@��sm�D��z�ٌI096S�
�殺���Bǈ���C"m94-����b�6w]`������&b©O��v�6�3�\�*�F�]�F�yN�m�.��Sp��z�{Y(�@�%��Iu��K�"96h'uH�vh����v�qkn�/i��j�*��أ���g���`�Hތ����lh�"�U�k���@!vn�I�so�"����&��73��p��Z_ݨr蔟Xlf�P�	Gs�!&ݺx�&�'L�*:/�Ms��] ���w���|#�WOjݗ\��&Ä���N܍�E��I�;v&�t��l�׃��{]��������e���`rH��E��2��&��2f�˺� �z��n��뛚���g�29�q�$q�wf09$t��}Iw�����Q>�Y0Y��iɠy��h[�s@�wW��f���uŉ�x��D�� ��x���m7���׀~��`�`^�ԁl���i(�����z���p�hptp����Ks'�=[:�AV�U*�V��u� }�� ����Q�C��}��Z�V��6��9�G�}��!E�� �HJ���7��`�r�h���)ac���"e�c{#�6Tt��-�n��kU���4�BC�RL�<�.��^�wu�{n�央`F(�q6v����u�rI.���=�ŀ6�ŀrP�J����T����uw6]$}����:�������'*�IgVMI�
��&2dS �H����|����ۗs@�^�@��VI��nLr8�� ߛŝ�N�]� ��Հ9m��p�'\X�'�)&
L�-�w4W��kv��c�.��bg�c��c�"f�Qv���P�r*�Ax�K ��M�D�`��S�% "���Cb��(6B�0L���ѝ�><ڟ(��}�x�]�x4���4c� Q
���@ V���VHiEb/����
�_����Q
�m�$����b��SԢ�|�o����*'�j�����?f~m��_���	$I̟��1��.�r��U��JI�����J_��i/�w����r�{���,�d���5�jKwfs���K���$�}��q$�H�����{��{�~���l;o��-g�Ystn����rc�p �lv�c�����mOe�į*�v�3�I/_��ƒK�}���$���[K�v��g8���z�%V�.��D�357m�����9�@?9�~��v�MkW�w�s���w���<֭�w���6��kY��Ԛ�ɇ9m��{��wm���\���RK��;I.IW8�]�-��ɑHcS�s��]�Y�%]��J�Ͼ�p�-�}FD`D�H XՍ�q~���<.����:Q�N7#�ry�IWn�RIw���J�w���ܷRK����'Xb�"'�sk���VU��vB����\s��G�8�խ��l��q�O��#5$�q$���4�R���J\�ƒJV��3�$�'2~mBy�IZ��ԒUޯ�J�u��I[i<�$�x�͘�<���nbԒUޯ�J�u��I[i<�$�wqjI+�ԳlY ���2�Ē�#���RHg8�w~���i$�_���%կ�o䘜��<$f��Ī���_��3=�ا���S3�����T��{_�p���?xO��~�1�Mk5���v���4��l��lٗs1�ۨl
C���Dy����z �	'cV�Ol�3��N��H���3f���:��v
}f�Qg���\�r��]��ݚ�\x��Cns�ne�����/o`ayø�^i�sջ(Z 1�o���R�nC����\���6������b�{r���kE�^�!u�.��d���7��^F�IF��n3v���w=�9kp��ۗ����Y�ݖ�r"�7��I�ۚ��� ?����� �d��$�R:��II*g8�]R[-U�QL��Q�jI*��J�w��Vܳ�J�u�K�u�5��7&9 �~x�U[��$���x�V˨ԒU�_�$���q=d��E$�I�RI)%L�JL�$��%�%�����߻.xd�
B~�d�x�V˨ԒR��$�R:��II*g8�]�L+~;�;3��	Ku����ɎE'�W��۴>�8m��V�{4Nx.�#�5F!c4�R��$�R:��Il�3���K��4jI+���YF���9�$�V��������\��ޝ�r�{Z�K����ߛk�_<��1I0@�̱��Sޯg8�R\t�^������~���W��~󱤒����
J�嬼WaRL��J�w���m~x�U۬ԒK��<�$�v��C`�ǩ$���$�܎ƒIl�3�I-R:�������ZL]\�ѧ�7:<�vصŪ�7h:_:vC�㣎^%-ˉ�7KLrA���$�۬ԒK��<�$�[��$�;k�Ē���OY�E$�HƒIl�3�I-R:��KnI|�Im�٩$�w�˞#��'��S$�Ē�n�ݶ�u��k��M���J&b	���~͓��Y�$���x�V�J��4��!
9�RIs��<I.v�5$��r�<I.V�=I%ߺ��C#�ё��^e�%�#����UU\���ޤ�^�Ԓ\��K�~��6��dDO�f4!�[2^}H��(���Շ'8{(���d�vz2b���L0�$g�$����y�Ir�q�I.v��%��f����R�7�$��&I�%��ǩ$��_�$�;u��Iu�g���?6�?�z4́$�2G1�I*����%��f��g���ڿ}�O<I*��q�I/*��s�ܘ�ay��$��}Us=�X�I)�W��I-R3[��K $T0�hP�u3߼﷜�߾�r]oS%�آ�`�f��^��<�$��_�y�Ē[~��q$��v4�_��کK֫����c��[���W��P;��;;\Wk��:/m��2K8.���{�wӌ��uq���o���}RK�6_8�[r;=�r�$�����I{�I}�21�2F�(�=I%�_�ffI���󱤒^���s�%�GV�Io�K��y23m��%��f��]��<�$�[��$���~x�^֫��1�
��fX�I-쩜�Ij�մ�]���Ē�n�RIy�j�ı��q'�I2O8�Z�um$���O_z�R��cI$��,�Ē3��V��jl�����Yx�JZ�GR��U��3������#��i�Aa��tk�� �n zV���;k�d$�t��[���t�k�	���07&6��T�l%cxx��vr�q2���ra��A�]��j�g ]�(��Ꞷ�u���m4���(��m�`�Cse���e���v;m��Y�5#X?��eM��p�hJ��4�w��{��g��up�X��:��2ε��=�wM���]���2ш��篻w�����-Yvu7?�����_��ۑ��I-쩟���Q{έ������&��k�r����?>w߾�{���}_}wjo���$�^�i$�se�%ߥ��M�b�I����Iw�,�Ē�c�i$�se�%�#������\*բH�jd�x�\��z�K�z�<I.v�5$��nY�%kĮl�'�X�B^U��]���Ēۑ��Ise8s�%��ǩ$��n��I7�Lx�܊c3����5�2\u�w��shxk��ݮ�\��[Ō��#FFcM���$�۬Ԓ]�ͧ�$�+w���ޯ�K��y��xI0@�.fjn�o�}���<>��A��ʫ����:�N:��J_v_8�[r;I/:�R�7�$�2/<I.V�[I%ۛ/�^����_��h&�&T��c#���Ȥ4}v���^���[09BQ?s�0���eji]U�^e�x������?����ݫ@��K;u��s��'�q�[�n�l�e�3����c+
�.��~}���^X��`�~��)�yzS@��j�O9�Հ}�`�jK�UE�� ��ٞQ	B^UCu�N��Հ}�V�铺�_f��y�j)�}��9{�ᰡ%�1\(P�B]8�+�`��w�+���h��i����ο=گ���fD�ou`�=K ����!aK3-����0=�G��{����R���PQ�A�
�=C�s�o�����-m�� �xr'�jO<~�}|Pq�,�WFfU��;�;&05we��7nO���?����$�`�R��ʪH�ݖ����097 ��B�71����bNM��^�ｒ���4�m������xآ�`�z�j�`��0��.ދ��H��,0�Ȅ"HHH�F({
BC��@	 E���s����>��a���7v��U�� ߛ�`v��n�`uM�����0;�Z[Mg���R�],H7=)v�]���n��u��J�d�u���s4ҳ� �ٌ����YUUq�y�����ȻWR+�UUU���u��IuP��<0&�Θwf09"�O뻬Y�P*�����m���,:DlU�M���y�U"X���q'��8h�0͘��-������`j���X�ԒcoH�h��h�����0�m�-�H! �	FA��4h>�Z���$l��� ��Y!)�V0ӲCf��D�țA��t')�L���H,0JGy�$$b$A��BFA`ČII� BE��$b�"F.�CA_O"F4���b�#�YQ����cHF1 �Xb�FB޳������� B!��&͒"ă�� �B�pX�Hh;�`�b1�[(�%j�D��� F"�"0��@�E�E�!$H�H�2		�#$`��'�b,`�A!F1a���FA�X%d!��I2>14�i��(<�2��R�Xő��d����?p�B�������  D5£��r��g-0LME�aB��"E�!�lŐb�p!��H�$�P�c���"��H1"D�$ �D�`A�zm�.f� xxo�jQ 5�B1F"@����rC�@-�R��ڶ�l�m��K\ۂڝ������Y#�	-"
I���Z��;p��U8�2;[mָ�
��:l���2;s[��{s�- �X���ܻ�3�cY�|�Zx����zi�(�;�2&�����l8y`iƉ�jۮٲ���/�rP7lv��K�	ͱ���6�E����jکl�v���m�r�"�nEyʐ3��G&�m��n[�h� �i�O<�*���kk�1���.9�>l6��v)�\.õ�F�6vg!Y���p��T�a�84IWYm� 'B�h��c��@gD�Uur�(�N���q��Qk�v�v�,:j��%*��籕�J�JN��k��X����&IʠsΖ9eۜv�R�%�G<�kδp&��LFv�G"�<@�J1����G/;�mX��Wm���\l5*����H���p�N��6E������m�J���UjU��WC���a3��Q\ŁQ�2m���;hyܩ��g)l�]�_F#t��7@�ß����t���2C��mS�v��u8^�݂�8�-T�,D����63�#Q����mf#���Tl^Nno*5AMV��R�I��t%��씥�7&mۛ[zۨ�Di��ST��f`�njr.	Ѻ%@lǃ� PiƛY�g$�W �'k.ڳ!E�yq�0'UһK�S^k��Uy݂R��^5��O����V�eɌ��od��U�m����K(�n���4P���*Ի;K*n: UVՁ�'U�/<R&��&�[UV�+ ���;]PH�\XP-J�O��CBu5���g`\旴gc�a�*ˋ��MaL�vݕ��D;��Ϊr�$K-o<�ic=V;3��:�,�rjT��:�Z�ں����Y���/�4�h*�Uv]��}O�!�*�i�e�ڳl۶p:��hݥv�nT��mW�Yƴ�,Æ��g�n�[c���Z��pdm� ��lJ�t�x(x�����x� >��_TO@�"�!���Q�
��_�܄��ٳ�9�4�==}MΆ��z�q�h�F!�;��&�{�Y�ڌV4�;��ӻh; R�PW�'�א����m��Ud�'wp\�m! ��n��tWgs�2��F���<h�G��јA�����5��g8�N��Ӥ�(�Q�	�+k3���F������#ԙ:�1*;a��-��1I�{Cnmw<���]1e����{����z:��Q��﫵�����m���k7�=��mtq.ۛj�	�n����6ߧ����	5d�0:��`s���]SwH���ٶg�BS#��X���=W��<�ߺ���nI'"R��, {���S;<���o�K�}q/�di<�rF����[��=W��:��;�w4��U=�&F����rh���yJh^���f������?�ݦ��5nˮB�g��c��{s�6��۫��1���er�yk�����H���4/Jh�@��W�yl�D�cQ�"
D�w��j�߿~`�j�
" �SI�C�QQ
�/u� �u��fٟ~�Ď_|��F������ �ߣ�l��Y�GLib��Y�8�NM�z��)M��sC�%3���Gq=�]MJ�.��7u�lՐ`odt�&��T�l��?��Е�ˮL�ۋ&��\X̬oN��8����]�����4t[����}�ۑ�t�]��{݋ ��z��BK�}A��?����K�6F��'$i�9�{��S&�>��� ߛŞ�Q��'�Ydh��m7&�W���@��SOs�?f$LgG���}� ;�^ ޺YWjn�`�M�]�z"=
��?�`}�X �]�y�~o��{���"X��ܑ"p�7�`�����׀kٶ`����.�&���1r�Ӵ�d2��<딸�k����v��Y0�
����O�<�4�E�Z�����]��m��C����{B�nG&E�9$�$���Y������v�ŀu�t��w�U&��5#�h�Ɓ׮�$}o�@/��y��u�r	d�)��ߖ s}x ޻��.&&!%�"�"@ſw���>����kI��4�� ��h�f�ה��o]��V5������#jg�Ft�C����� �����T�Sغ簆�a(d� �6��@-�4��4z�h�@��������d��G$�6j�?RG�<�zOc �f09&E�,X8ԑ"p�-빠�� ���:��=^�F��$bx2K�`vc �f06j�0$����.�dxӒH�NM ���>�~�8�s�X �]��U�}	t)Q�Ͻ�}��w���~���C�n�85��.^��_%�T�fΗ=�L�Ë�C{b�s���:�ٝH3fwt�\z̼�c����bէ�غ�k�Y���b����s�YL���qgl���V����pjqez������m��x=���:�ݍ�(�ٺ@�v_�>��t*���lW-87�s�݉�ƑA�N{;U�q5����'9D{hɵ��w{�w���������C1�I¨�X��v�����I��:��=�{C��[���8��X�"�p��|h�������@�}x����Tݕ*�n��x��L�7׀�^�f٠y���6�A9#LQ���f�u�4��4�w4Υ��A�B,�7&�u�4��4�w4�Y�[k������d��)$�:��:����f�u�4�iborI�H�9sŷ�v�]O[���g�nrg*����z�[�Ȋ�X�$��{6�m��o�@/u�}�4��4W���29���iw7f =�x�_�	J�	$� ���x�fـ?�ٝ
�2m�}�rc�ӒH�NM ����;ڥ4��4���=���F��̎De�c{A�;���y.�{�
�F�xԃY$�C@�zS@��I=� ��c{A�߶*%�/�=�8�|s�7lcd�r�,�`��s�q�l�][���'cģ$M<�rF��C@;�� �ٌ��	��06��,ªn�ʪ��� k��J!)��� �����f����nLr~2c��`lՐ`N�A���k*���&s�@��T�5��0r'�ј �]��]�t%
_9�0�u�X��r1<�C@/u�}�4{6�����!ms����M]̗E�*�<f��G�n��j�gMcn�d���:8�d�64�rE&)�9$�$���M�)M�Қ{��=���F��̎DG$�:��/�)��� ��������G�8��R��4�Y�޳@��S@�%Y�4�WwSD�Z��3����׀kٶ`(ĢP��܅	Em~f�=YbR4��,m7&�_z��)M�Қ{��>Ͼ�?�rL�B#C�Z
�RL'9��z�v3���a��틴g3�^��$�&1�RI��Ɓ}�M ��h���<�U"X���$Ƀq^	��0ݘ�96c{A���tk�G$�Ȥ4���/Y�%����7� ���@y57je4�4��@<�f���)�w�)��f���h��4�6dr"9&����?�ـ�� �� �Id%~��^��.٦�\�ĢM�.5Ş�z%�G<��m{�7G=��[-����:M���`М���[��i�ٳ���YN�'c�N���}���,VU�Iy؇�۶��[�p�I�Ͳ\mi�;%Ѱ�����[�ݗ�n��q����GO"�:���l��g�'sIմ٬�l/ ��5˲�yݍc����tH��h�9ŞK��D�y ��a�O�"�-����=K9gs֗�Ck�l\%ϵ���<F6��\���m�i�D`k[<<ݴ<F�g���ͷ����`�1�N���,��))c���'$i��4����Y�w�Jhޔ�.qU�$J�X�nM �ٌ�Y����`rIl12Lra�%$�{T��}�M ��4?����@���D�cR8�Ƀx�����`�1��� ��3���>�Rc���2H�?�7�ݏsغm�mGk����ju�zx������>�����]-1f ���&�`mvd��h�
��LNI#I94��ne�߫꭯����	7 �6l�~��F��̎D)$�=�s@�zSO≓_u����ڃe�*nU]qk+3)��܃ �Ɍ�f0����S��߾ľز!���j) �B]Z���>ŀ?�ـln�#�����5i�7G�5�a�v
y�/0�Wm�]�y���y{�w�����Qk����Հ}�^,^�_ġB�_P�������T��]�Z�&�� �V�X�r�&0"��~�#��yf%Jřx���]����[�%b[�DD~���L1�z��*D�[|��)��`]r�n'��_M�x!�&��4�� [�i]E@M�b�c5��#3�����0���SqKa�遨C
/��10Q�+�|���� ��U㜂��'��` �O"�y��@@�胈����U*!�}_���*p�*�>;������t����-}yy��YwB3/)����c/O[�"t�ٱ��h
��&
'$����+��u����b����<�P���\��4���p��4�6�y�㝫dn��n^���XT�q:�]{g����i�m���N�6:`�1���[�A�3�b��G���s@;�f���^��Z�4=��ز!���b�f�od���l��I�[��y���c�(H�#ȱ�ܚW�h��s@��sC�˛��۳o$�&?<%�&vD遳c���l��0=���~v�����\N��b۴bn������t�MȊz�r�"u����(8�)�k�Y\��t���-�ݽ��ݑ:`z��F�8�do8�h�����`wdN��09��[���]�f`��;� ��ȝ0;�:`onE�y��D�ّȠ�4>]~�y��y�{r&vd�Q�k^Yj�Ww6���XBKv������O=��rJ��OU��V�1H
AGH�ZTtUh�2$ �D��n���t �)(:(�"��ϳZɘM[�$lg��l�ݼ\n���KȆ��J1Q��Aw=�ۧH����m'i���r�i�pƺ�M�s�.�@:���Mѫ���/��/��=���i��u�9�������;q���v�HR�7Y�V;l��jlf0j�{a�ؐ�.ىY����\G�n~�>,����"��vb�=�q�1iu5#�{P�5�7*���V^[�S����w{���m��M����+��#]6LW���v�P��f���u��vs��n���*:3�fGKw�o����`wfA��؝0;�:`mt�lņbP�"�&��=�)��?$s�4z���]�@�n�1�pra����ۮq`kx��(K���׽8z�Ӏy�U"X��$R0♠u빠y�npu�p9N������Suwwj��E��09ۑ0=S�<��y:`l빠�Q[U��Ld���_���&�[v����7<�v�6�m;b�͵A�'l �p�nI&	���>4oU��u����A�?�Z����X�Ll��X�����8�Ӆ���.�$�/B_|{~�,��|��)�w���5��7�f�Lv�L�}IOL���{��MĮő�N8�#s4=ϟ]��_���<�&@��^�f��q~zE	�y��+�L��L��&�Lm�}���s��)��i���#���Wl�^y�lv��v{OW��de��`�(o����n^b�(�����/�o�����t��܋��W_����|��"�� �f���t���-��ݖ��:~�H�ٍ~����cRf��|�W�^��~� 0�X"P��X� �P�AqT�.����ܓ������I�LM�$Ĝz�ޯ@�VA���釾[~����/;K�l��Ez��4�{�}�x/��@<�f����QHMi��m(5�Xa�n��P��v6����y'[f�VWkDQ1HۊC@���h���ζ}� ��S�@��K�"�q�D�h[�ߩ ���������L	��H�"P#Ȳ4���[4=�SN��� =���ZR�Uv�qJfn���k���>�b������<R+,�:�Yk��q��Nwc����{8��c�� ��>$�����,4��w�v�흊�u��\��n��	��m�NnM,�z���Ԥ�^�Vepo���&09ز�c�o �[	�i�$�9&�y�~���}=� �}� 7��:!L�9��S6U*��J��0;�^t��v:`�1�r���
6=DlR6�s4>���Or�S޶ɳz��݉�`l�%�!�D�0�f���^�����_��<�띛�{�lܒ�=���DTO"�D�ݝ�ə�d�e�f�&:.a�8���&ݕ��nٻ^��DX���j;t�	���uH�]g�1��v�$)�;�iSC�.Ʒd�1v�c�XY8��.�����M�-�wV�:�Ә�*]�OV�y:��r',�C����]jt�����}G�ix#�vyC�۫Plk��%�hs^�u�خ��Z�k��qX�3]3�u\nr�+͋���z��{�w�w��s��;�2fw`����V���cW�qmr����ş8:����.0����g���2<!1����@��R�{�s@�u�@��ن&890���Qɠy�ͳ?�B�J����l��X���:g��|������0N)��|h[%��f09�YveZ�2�.���J��09BIO��� 5����6�B^P�V��x��	��+�5SUw$m����4=�)�y�S@�u���������h�L��R�=Wm�pk��pUƸ��v.��m�5�p���{�./�A�l�q&���U>4:�h{]�DG�[��9�⨬�ꉻUW9�rN{�}7�@FE*��7�3ܘ�;ݘ��b�?W��D����ĕ����+����M���wvc��:`sl��綷�P�QD�h}����׀}�=� ��ف�DL�����B�����*�������/�K��ǀ��h��hu,M�NI�	� r�ɣ��ˣM��X�V3b���N؜9�ݖ�r����d�G�cPsd�'��ߧ� �Ɍ���Q��veZ�2�]ک�J��0~n�&C[��>ޞŠy�S~���;��-�16��H��`�׀~�ͳ�(��B!EDG�X?l��=�h��+�Q7��nL�Wx�O��ߖ�u��w����+o�@���lǸ�8��C@�L��W�o�� �{�Y>��@�7`��Si^,��q��s�] ��9��x���6Kd�?{��j���fa�	��0ݘ��b�09&A��n����e\]+�u3wx�����*�_��`�_� ߛ����Uu��ɈRM�j��<�SO�"��M ��4}g;�51Lr �Rf�DO��� =� ��xDB�	,��%`�����'ʡ�٫���Uz�k!�H)��$4��h߳=�޿����,��ӳ��SWs%�p-��v�����ݱ���wCv6��=�-���Gܹ͂�.�&b�����������:`Ṅ����c}�^v,Wj�\�\�Uw�~��Ş^QTy��`?z���%�NmqTQ��우UUsV�޾0~n�򉓛��>ޞŀ^��͑�̉ƣqI�ٟ�����='����0�K������ي�F�~�"�I&�^�4=��h�)�$�Ͼ�� �OU�"��*�,�&"Ĉ����y�R|�@�a �dG�x��C1b0��<$9���&�(�UM+�H)���7^�њC�`��J��'��k@LЈ�j)P!�K����z�#8� �H1�P��<ւ�@X0MA� �Ϫ��!1����׾�p�����ư="�";-V��GJ�����<SC��w��`�"�T�q�=aB1H�<P}|XB/��vն����	 ��Jj�m�� Zv������j�[I�W;*�1cUu�	@�*�E��VG��W�ug;���㢉0B�tۃq�������(�\�c�����
x;�f��nob� �g��ӌ��h8u�'����*�
��e-���	 `U�(�ڸ�g�6[-�f�xऴ��9�lf�&�[;�;���
^�����T�VM��tvm���b�s��ێ�vڨB{�v��u�صq>��@_l��c���&�kv�����ۓv�ŭ�8�t�V]�॥ �퉪� ��-l��-[KT�����]�J�����UƝX��+*��;�v*��T:u��9Pcc��K������הv�͊���l����z�dhg>��������I�iK	͎����^�ܑ͎�N��%\
ڼ�n�Jm���{l46��i,�lڪ8���N�ͳ�� �nzbjr�U!��`q�0lٰm��&S�2�&xب��o;��6{"�����9M�ccmfv�(9v��S�v�K�ir��*�j�3���A�wbk�St�S΍��9y�x.@���MJ�]���X'�6�&��ۮ��W8�rl�:��^4����hE�SUV=�r�:yb�%@�`W:��rH�Pj�K�U�<-�#[u�۵��gZ��r�y[T��nԒ���B�HOSm�⺯;-�`ѻ{z'Q�UR�ԫJ��S��H��n2�*��\�;*NM�t��!*�b�`�����US���) �vtn�ꚤ�&^2��gI�!��QRJ�p�̬��;&v�ֶvU]��Z����QPM=]�5.8�v�u��2����@�N��L�ٵڹ����u$�� P��[�Hm�lMM� ���m�8,�;lm��W/�l�@i
�Y`��vawޛ��A��u͙Ӭ�0�&^��3=�Vە��q�q�V;mf`��Y��UD]'�'��5[��)H���&�|�t*��N m`/H&C�@�"z
�>�>�����5�@険����sc����f;5� �lkA��n_Z윖����5�۩'q�a;`�i���]2��=I��#�h����3\&.�����N$�rq��3ƍӫ�E]��d��;Czv^�D�9��k�t�z�f^1۷�,�ܨ<��1
vP�g:&x�nHe�nvG�H��8�NQ��t�6�֘1مGMm��1�v~���WF�P�:�APq��Eǌk��C�<;����$G&���$H4�œ��)'�����0���I�`uz�������e4��h�@�ڮ��f5��$r&��!��1�vl�;t��̃�AK[�b�8��$�ؗ}~����s@�l��ߒ���@�����k8��5y�v(遽���f�`~���naR�Y�<�o0���@S:�ִ[�k�|���u���n�v�#N�@��˝sVX*��^W ����7�c �ٌv(�@͑�̉ƣqI �m����h��AM�%�b]w�ͧ"X�%�罽��Kı>����r'�5SQ,O~��Z�33T�4e,���r%�bX�����ND�,K�{{�iȖ�b}�wٴ�Kı/�����Kı<���&K�-��p��fӑ,K?5߿_�ND�,K�~���Kı/�����Kı/~����Kı<����ɬ.�2Mk.��r%�bX�����r%�bXhX��{��yı,K߾�m9ı,O=���"X�%�~��IܗV�uv�:�}�t9n���9�]6�;E����vm�v:q��z��k�
]��O�߉�,K��{�ND�,K�߻�ND�,K�{{�a�'�5ı;����O��Y��g����d�����̠��r%�bX�����r%�bX�w��ND�,K�{�ͧ"X�%�{�{�NA�,K�ߥ�53WTѬ�̳WY�ND�,K��{�iȖ%�b}�wٴ�K?�о�v��xdMĿ��ٴ�Kı/��m9ı$�ͮ*�?*����UWsV�����D�߹�m9ı,K��߳iȖ%�b_{�siȖ%�by߯xm9��{��������j���[�w�x�,K���6��bX���w6��bX�'����ӑ,K����i��7���{���ߧߣ��c�ѹէ�p��n����,��Ρ�؝��\��\�S2�1�2�ffm9ı,K�~�m9ı,O;���"X�%����fב,KĽ��ͧ"X�%��w�2\2�]�[s3iȖ%�by߯xm9ı,O���6��bX�%��m9ı,K�~�m9�j��X��w���rܓ52�F�.��r%�bX����M�"X�%�{�{�ND�� A�MD�~���r%�bX�����iȖ%��{������Ϊ�'.�}��oq��K���6��bX�%��w6��bX�'����ӑ,K1�b?��!��C��N���ӑ,K���d���&b������7���{������Kı<�׼6��bX�'��}�ND�,K���6��bX�'�^�����7���=k7�f�ZrNca���O�ݒ������٘���w��yx�t��k.�,��f�Ȗ%�b{���ӑ,K����iȖ%�b^���ӑ,Kľ���ӑ,K�����MN���,32�̛ND�,K�{�ͧ!�j&�X��߿fӑ,KĿ}��m9ı,O;��fӑ,K������y��,U��7���{��;�{�ND�,K��{�ND�ı<��}�ND�,K�{�ͧ"X�%�罷rvf\�a��33iȖ%�b_}�siȖ%�by�n�6��bX�'��}�ND�,lK���m9ı,O=��ɒ�Mh�CsY�ND�,K��wٴ�Kı=����r%�bX������Kı/�����Kı �A;QT'twZ..�C'X��E��l�_V�\f�O$c���u�ɥ'-�6�vAD����ݷFR��Vv�v蛶T�$dKv���f�uG'nJ�]p������Zk�����
}V.p��!��wX�l���ט�I�-V4��.:����n�ѷ%:��)�2Gm�؂���ݸ�����N��ӧ'�]�q�)d֣�-�d�\]��BT��j�~�����������-��W	��f��[���z�u������N�\�N��-�&�rqڝZ7<�[�w�ı,O����r%�bX������Kı/�����E<���%��s�B�B��������LU��]YwU3Y��Kı/}�si�~ �&�X��~ͧ"X�%������ND�,K�{�m9Kı=��/u�L��Ys32�ffӑ,Kľ���ӑ,K��M�m9Ƌ����pI���ͩ �'����au�m�&�� =��~���r%�bX����iȖ%�b^���ӑ,Kľ���ӑ,K�����C\5�ɬ�L̸fM�"X�%����6��bX� _��siȖ%�b_{�siȖ%�bw��m9ı,O}�-�u�5�L�e��U��;7a�5�j�u�<'\n��c�۵�a#m痫�5�p�ˬ��k.k6��bX�%��m9ı,K�~�m9ı,N��͇�R'�5ı;����r%�bX������f\�a��33iȖ%�b_{�si�m�M2&D�;���r%�bX�{���r%�bX������Vı,O=���e�,��)-����Kı;���6��bX�'���6��bX�%��m9ı,K�~�m9ı,O5>�f�d̳��3&ӑ,K�>����Kı/}�siȖ%�b_{�siȖ%�bw��m9ı,O=Ϯ��9���k&f�3Xm9ı,K�{��r%�bX�����r%�bX���}�ND�,K�{�ND�,K��l��3Y�����H����׎6wL7vr9��zض���q[�Y�[��f*�j�{���7���x�~���r%�bX���}�ND�,K�{�ND�,K��{�ND�,K���jf���e5�f��6��bX�'���fӐ�"�uQ,N����"X���MD�����r%�bX�����N��"�TB�k�P��*�˻�Y�iȖ%�bw���6��bX�%���6��c���:ODޝObr%����ND�,K�zo��r%�bX�}�ޜ��Ӭ��\ֲ�d�r%�`ؗ�{��r%�bX�����r%�bX���}�ND�,Q;��~�ND�,K߻n��3.S0�Y����Kı/�����Kı=���6��bX�'���6��bX�%���6��bY�7���X����4���˒�V�q��ǭ��v;bŇm�����X.
�Ec�&Hh��fӑ,K�����r%�bX�{���r%�bX��{���%�bX�����r%�bX�j}��Rəf�.a�6��bX�'���6���:���%�߿fӑ,KĿ~���r%�bX���}�ND�)5Q,O���=���RK�����7���{����m9ı,K�~�m9ı,O{�ͧ"X�%����fӑ,K����m���L�T_{���oq��d����ӑ,K�����r%�bX�{��m9İ?P�Q�Dx�$M���ND�,K�z_���]SZ�k2�]fm9ı,O{�ͧ"X�%��߿s��yı,K߿~ͧ"X�%�}��ͧ"X�%��ѝ.d�+��*��ӕ�k5�Ӻ�Н�9{x��X��]F�8I�N�2^rR��w�{��X�'��}�ND�,K��{�ND�,K�߻�9ı,O{�ͧ"X�%������f��d˙�e�ɴ�Kı/�����Kı=�~�bX�'���fӑ,K����iȟ������'�vݓ��.f��e,���r%�bX�k�kiȖ%�b{ߍ�m9���Q5�~���Kı/~��6��bX�'���2�J\�2CD�3[ND�, �=���6��bX�'��}�ND�,K��{�ND�,�$�O��kiȖ%�b{��ߦ�d̳2e���fM�"X�%����fӑ,K�[���m9ı,Ou߻��"X�%��~7ٴ�Kı?!��w�����\�HN�PZ�tganLW�s����t3F9gg�ڽ\4��]��l�F�Kۇ�Ưj�XMp������۶�1��s��u������)�1��V�:�ϊ!�khK���(DW&�5nwF�<���m�y�J���u6�-1@��q��2U��ͳ�AZ�F�l�!xvJ��;I�����l7���̤�n���}������{����}�=�L�M����\�;gb�^��.ks���0�,z�§\F.������fj�32|�D�,K����ӑ,K��]���r%�bX���}�yı,O���6��bX�'���u9fj�Ys32�ffӑ,K��]���r%�bX���}�ND�,K�{�ͧ"X�%�~��ͧ" ؖ%�����53WTֲ�̹��f���bX�'���fӑ,K����iȖ%�g��߿f�Ȗ%�b}�����"X�%����f�f�,�!�2��iȖ%�b}�wٴ�Kı/�����Kı=�~�bX*؞��}�ND�,K��-���]:ɗ3Z˙�iȖ%�b_��siȖ%�b{���m9ı,O{�ͧ"X�%����fӑ,KG��~��>q��	`�����!�
�n���Y:@8��]�f{]����wu�v��+Q�2�ffm9ı,Ou߻��"X�%��~7ٴ�Kı>����~yQ,K��߳iȖ%�b{�pɗ&[sD���m9ı,O{�ͧ!�*� RQ>�x�@�	�@�yq,O>��6��bX�%��w6��bX�'����ӑ?j��X��w��Y3,�2CE�5�ӑ,K��߷�m9ı,K���m9��,Ou߻��"X�%��~;�iȖ%�by��=��uV�%�o����7���{��{��r%�bX��w[ND�,K��w�ӑ,K����iȖ%�b{��ۿ]�5K	UW�����oq���w[ND�,Kʩ�t���%�bX����M�"X�%�~��ͧ"X���~���?�b�iֹG:�b�Vݱcl��8J&���v9�=�:-�n]��/����fCY���fkiȖ%�b{ߎ��r%�bX�{��m9ı,O��{��"X�%����iȖ%�b|zI��s5s5u!�RS0�r%�bX�}��m9�D�K����m9ı,O����m9ı,O{��ND�,K�����f��d˙�e�ɴ�Kı>׽�bX�'��{��"X�v�@!����ڦ͊MxqD�b��<�m�7E� ��ҍ `h$C_b:|��oD#4hH_���A4�U>$ �mX���Щ(14��H%5U��ڏ.�`4l�f�$�SR�&�*���@�����me�Z���G�� H*p�|<4����� �� ("�@�D�\ڞ�>�J"�5؛�g�6��bX�'~��6��bX�'�ϭ�;s�h����ӑ,K?	Q>�߿kiȖ%�b}����ӑ,K����iȖ%�b}�{�m9ı,O=��2L˖��2MI-�kiȖ%�b{�gxm9ı,?# �s��yı,N��ߵ��Kı=�{�m9ı,x����~��5t�m�\�[����jם˼���7;���e�^���r��d�E�m{E�Ma��Kı>����r%�bX�k��[ND�,K�w����Kı=���6��bX�'���]���3S35L֦fM�"X�%����u��Kı=�{�m9ı,O}���"X�%����fӑı=��;�9���]\�̗Y��r%�bX���bX�'��w�ӑ,K����iȖ%�b}�{�m9ı,O��/y����fCY���k5��K��{;�iȖ%�b}�wٴ�Kı>׽�bX>�T
 A����Or%�;��r%�bX�=$�f���f������iȖ%�bw��fӑ,K��^���r%�bX��w���Kı=���6��bX�'���]p��v��)m��.�Aq��,q�v�c�ppA��t��pJ������}H��Rř6�D�,K����m9ı,K�����Kı=���6��bX�'{��m9ı,O}�]�ٙf�u�
���ӑ,KĽ��ͧ �bX�'��w�ӑ,K����fӑ,K��^���r%�bX�{�x�L&4e!��Y�ND�,K�{;�iȖ%�bw��iȖ�b}�{�m9ı,K߻��r%�bX�j}��Rəfc��&��r%�bX�����r%�bX�k��[ND�,K���6��bX"��｝��Kı=�;twP��̙��f�32m9ı,K���m9ı,?*u���f�Ȗ%�b}����ӑ,K����fӑ,K��w~�ߩ߻ߎ����Z�g&��c<�s�n<kv����+ڮ�Y�0FvnЫ���	z����3��T&v�/zh���8uC۶'Yl�J��jt�.���r�(�퉤7d��u����A�Xm�+�lm��칼�WA�v�%kƪ����q�v���r����&���C���1�L��	��A�qq��&�M3V9�:m�y9eD����&�~{������o�ݟ��k\�XNHם={m�W�,nޞvcr0��86�e�����n�;}R�:��\�ͧ�,KĿ���6��bX�'����ӑ,K����fӑ,KĿ{��ӑ,K���������fd5��nk3iȖ%�b{�gxm9ı,N���m?>T�KĽ����r%�bX��~ͧ"~ 	���bt����f�\��˖ۘm9ı,O����iȖ%�b_��siȖ?����w���r%�bX�~���ӑ,K���Rޜ��Ӭ�s5���6��bX��~��ͧ"X�%�{�{�ND�,K��w�ӑ,K����fӑ,K��ߥܝ��jGZ0����ND�,K���6��bX� �����"X�%�߻�ͧ"X�%�~��ͧ7���{�����~�̡Uюi^N�ц۞�V����o[C�#��"K���JC��HoV3$��)2K.�6��bX�'����"X�%�߻�ͧ"X�%�~��͇�yQ,K���ٴ�Kı=����T�.I�蹆d�r%�bX�����rSH&�� �MD�/�w��r%�bX�߻��r%�bX��پͧ"X�%�߾ޮ��U��32�32m9ı,K���m9ı,K߻��r%��bX��پͧ"X�%�߻�ͧ"X�%��~'um�fkYu.�5335��Kı/~�siȖ%�b{�f�6��bX�'~��6��bX؟k��[ND�,K���jf����k5r��fӑ,K�����m9ı,N���m9ı,O��{��"X�%�{�{�ND�,K�}
nt�K��8�ȍ�m��c��=`�/��ݻm:4#n.�xx�,�D;tX3o����"X�'~��6��bX�'����ӑ,KĽ��͂�%�bX��پͧ"X�%��~��9���Y35��s2m9ı,O��{��"X�%�{�{�ND�,K�{7ٴ�Kı;�wٴ�A�,K�~�s�̰�kRaK���r%�bX��w���Kı=��}�ND��`��Ѹ���w}�ND�,K��{��"X�%��w�d�2��2MIe�fӑ,K,N��ͧ"X�%�߻�ͧ"X�%��{��iȖ%��&�k�~ͧ"X�%���߮�f\�1њ�2m9ı,N���m9ı,N���[ND�,K���6��bX�'~��fӑ,K��(!��;��:]]��^ӈ{Yݣx,�m���@�c8���wk�����?�s�V;�'��[�&fM��,K��k��涜�bX�%���m9ı,N��ͧ"X�%����B�B�������	�wuW4M]�.ffӑ,KĽ��ͧ �%�bw��m9ı,N���m9ı,K�{��r'�5SQ,N��sS5f�fCY���6��bX�'�����Kı;�wٴ�K�,K�{��r%�bX���siȖ%�b}�'N뙗.]e̗Fd�r%�bX��wٴ�Kı/}�siȖ%�b^��ͧ"X�P�s���u�8 y�O��ߓiȖ%�b{��[��\�nL�f�\�ND�,K����r%�bX�{��6��bX�'~��fӑ,K��{�ND�,K�Ƿ}��5�Kutᬜ�\<���1��s�c���YN8K4�.5�#^ L�e��F��f�iȖ%�b^��ͧ"X�%�߾7ٴ�Kı;�����D�&�X�'�~�ӑ,K�����fj˚&I�,ֳ6��bX�'~��fӑ,K��{�ND�,K����r%�bX������H/���'��߮�dԚ4SWF�7�Ow{(@�'�w!x�=��!~ı,N��ͧ"X�%����S�52k&kX���a��Kı;���ӑ,KĽ���ӑ,K����r%�`���~��"X�%���vkZ��2��Y���ͧ"X�%�{��ͧ"X�%��~7ٴ�Kı;�{�iȖ%�bw߻ͧ"X�%��(�o��y˳T�������t�ٲWX �q3p���ݨ��z�qu����n�𛖖 U(�a�	ed)IpE�l\[��5�OX�+vѶ ��,����:x���RΖ�H�	ζk��s�w��r�-�u��n�}�&lAp�&ݏ�� ���;������.��	��r�m��)���Eg!m�p��m�ڗ ��;n��i~����m�\/}����0�]�{:u�]����ݛ�uX\�^���@'d�X���{�^/�&u[�$�ͧ�,K�����r%�bX�����Kı/}����Kı/{��ӑ,K����;�f\�u!�2]�iȖ%�bw���"X�%�{�{�ND�,K���m9ı,N��ͧ %�bX������\�nk.[�5�ӑ,KĽ��ͧ"X�%�{��6��c���j'�����Kı?~���ӑ,K��^����5#tL-���ND�,��DMD��߿fӑ,K��ޛ�6��bX�'{��m9ı,K�{��r%�bX�{�xᚺ�SaA%U�B�B����ͬ�!r%�bX��{�iȖ%�b^���ӑ,KĽ�{�ND�,KﳷZ���*X���]��g���{I'F[��"�'���]�E�I����;����i�2m9ı,N����r%�bX������Kı/{��ӑ,K�����r%�bX�;��;��L�5�urfd�r%�bX������<6��"X���3iȖ%�bwߍ�m9ı,N����Kı=��˭Yy�lɆ�5�33iȖ%�b^��siȖ%�bw��m9���Q5�߿p�r%�bX��߿fӑ,K��������532�sWY���K�D�ޜ�6��bX�'���ӑ,KĽ��ͧ"X�%�{��ͧ"X�%����s2��js%љ6��bX�'}��6��bX��F��}��m<�bX�%��fӑ,K�����r%�bX�{&[�u��3Ym��r
͙;\�1�f��+��зn�uϷOc;�5��p�����1U��7���{����ͧ"X�%�{��ͧ"X�%�߾7ٴ�Kı;����r%�bX���ۣZ�XP�&��ͧ"X�%�{��ͧ �6%�bw��m9ı,N���6��bX�%��m9ı,O=��s&��sD�5%���ND�,K�|o�iȖ%�bw�ٴ�K^
��@�T"�H�0tb���(� ��SL�J�
�@
����
z��O�,L�y��fӑ,KĽ��ٴ�Kı<�oou2��ԸjL�3&ӑ,K?!Q?~���iȖ%�b_�~��ND�,K���m9ı,N��ͧ"X�%�ӿnS��Әf���L̛ND�,K���6��bX��D  .�~��6�D�,K�zo��r%�bX��wٴ�C{��7�{�w���{����b��Du�s�}�睸��sp�`F�F�u���m[�Yp��fkP�k5����ND�,K���m9ı,N��ͧ"X�%���}�D9ı,K�{��r%�bX�|^�S5f�fCY�����r%�bX���}�ND�,K���6��bX�%��m9ı,K�����O�j��X�|t��k���ˎ\�tk�"X�%������ND�,K���6��b���b^��ͧ"X�%�߾;�iȖ%�b{��[ә�Z2ffe�s2m9ı,N���[ND�,K���m9ı,N���ND�,	�q���G��݈�ȟ�~���Kı=���u�5ln��3Y�iȖ%�b^��ͧ"X�%��~;�iȖ%�bw��fӑ,K����nӑ,K����?<��������Md�^���0n��v㶞$M�s��cab�Y�f/ΖkY�ND�,K��w�ӑ,K��{�ͧ"X�%����ݠ�"X�%�{��6��bX�'����f\��W%�3&ӑ,K��{�ͧ"X�%����ݧ"X�%�{��6��bX�'���fӑQ�,K�~ܦ��\�Z�:�32m9ı,O����9ı,K�����Kı=���6��bX�'{��m9ı,O{�e���e�
mU�ws����'���^��y�%�b}���M�"X�%���}�ND�,�>�;۴�Kı>>���jꙙf�[s3iȖ%�b{ߍ�m9ı,N����r%�bX�{���r%�bX���siȖ%�ba�o�GJ�0z�
����ד`��[9�jȋEtWsJF�YF�' �P�h�&�S�8TL4�ʢD��P��m�P8�$���, Ra�!
#ثD�@J����Z�H�h��
����6�����ڏ��_O|Q8���&���$�_��:zN�L���M�nÇm[��BE��`  �K\������AFյEq�� b�X�Y&�V�+��6K�@�U/-��s�ǥ��#�]�I��vk�	lvts��j�G���эgO�HN��O%.KOB��\��1����oR���u��[Q��[5��R�#�P.=�۴k���4��6�'	px��I�����u��mN�v�>�B�r��<��:��N�Qo�X��K{D���@���e�-8u������{YjM�8���k��cl[���nm�������^�X :�a��t��r�ݻ�Aāuѹ��e�m냰�@x�k36� � � 9�c�V:øf������\:[����'i����4��,�Bz��lg)݃J�� �Z�Z�wY�UJ�r�8VV�L����N��8a�R��	���!<m=bEi�-#��s�շ�K:�d���h�W'Hk�]��Xظ��ef2�>��p�g�l�ݲ[ؔxz.Vo�M�[�[��L�ڑ��8@��탧Rg<���3��.Q�-��v�kHa�v����2��vy�����e�.̕Z�Kl9����(�6�6'Kнk�H�]��r6���O60&*Z�PUQ�+���-�A��m�v��>�)�ۮ���#1scK<#א:<�V GF�)�`��RGB�ƒ���8����V�2E�u�i�˲�]J�R���q��J �٫[@���쬛�Q@�R��Ֆ,c��p��-I��Yr@9�N)!ƫ���&,8������#)-URq12���Ynַ	ֻ&UҲԵ��WIp�g������L�[hi釦�F� �<����vX6:�tnԋ��U悖
�vUUA�B2۴�m�l��[�I@R�U]�@/,���lZlh�i׭^���n�m�	�[U]�{�ղ������nѩ�KÜ�v	f� �jMY��_��� �Ev����6<�J�� ��A�U3D6
G�爪|"h���}T8�>��}�30�2:�j�.���7^Mۍ׮�ƼA6�`��N4N�ts�B`�2���s�;<q�{vq!�C�d&]��\��tj�ͩ^{]�☠��Ը�<.�뤒2���W�ݗ�5A��O�7Yͤx�cj,DX�����ɛ=��Y�JK,���-Ýi���-�&/A拎;`�큲�Q�M��n�N�`
7D������=���}�DV�2 �mr�Nւ�|��v{,�9×���n�}��8wU���-��\�3Y.���Kı<���m9ı,O����9ı,K�����#<���%��m9ı,O����s.�d���r�d�r%�bX�{���r%�bX���siȖ%�b{ߎ��r%�bX��wٴ�ı,Ou����w�:ԘS5�v��bX�%�{��r%�bX���}�ND�,K���6��bX�'��{v��bX�'���9�2ܺѬ���Z��r%�g�����6��bX�'�߷�m9ı,O��{��"X�!b^��ͧ"X�%���^�Y�&f��Rk0̛ND�,K���6��bX�'�gݻND�,K���m9ı,O;�}�ND�,K��ݤ��ѣY���4e��k���]�	ؖ��&51��Ӹ��e���<]����ܦ��\�Z�:�32m<�bX�'{��v��bX�%�{��r%�bX�w��6�g�5ı?~���iȖ!���~���d�]�̻T}��oq�X�%�{��r�~��|E <�"y����6��bX�'��o�iȖ%�b}�}۴�ı>=�^��kSS3!���nfm9ı,O;�}�ND�,K���6��bX�'�gݻND�,K���m9ı,O>>'Mk���fdɚ�p̛ND�,K���6��bX�'�gݻND�,K���m9İlO;�}�ND�,KޟRޚ�]hə����ɴ�Kı>�>��r%�bX~D#�߿~ͧ�,K�����ӑ,K��{�ͧ"X�%��K��>3���N%���p���#O�om���qn��ݧ�OV�䛠fL.�zv��s/Ȗ%�b_߿~ͧ"X�%��zo�iȖ%�bw��fӑ,KϾ�����H8�7�`���/�%L�m�LI1�"(��*1awS6�.�]�w_��8\%�J���r 0H�H�GQM0 t���!�Ϲ�ٹ'<��h/Ac�/�bn~J����~��}g n��V�%���� �z}eL�<b��6E��4-�M�w4]��w?ι19#$Ɩ6���]���5�^�*�M�#���.ǷGj6-˿W����Y$1ƢJI���O��w4��>�P�H�׀|�G,�����,�2C@����uzm�@�ܔ����U�}� �2H�(G3@�[��ۼ=	B���|`�ذ��$����bĤzm�@�ܔ�-�VIl$���}߳��k�WWAuJlk7&�}�)�[n�y�Zm��m�w��~V�j�"ʘ�rj��ݫ���F�xz��ܜq�]ճl�g��ckZ�1��$4m��/>�@-�}��w�>4�����n~���/>�|�d;�� ��_m��K�Cu�^U7wt��Sj軫� ����?=V�<�J!)���X�}X�[2򋩩Wv*��������5�`�ذ��8	(�����7�#�.ɫ��,��m]�m��=
m��;�� 5l�%=R�4h���ˬ��m�d˔����.g9��:����BEc�kH�I��.ʗ�⎷��T��l9�gj�
�0�4!cMWK�;�ΐf�H���4�[\�nx�#q�g�T��] []d�6�鞮�.'9��v��|�K�+��U)볍�oj�["ln��m�j1�GT��<<����ƻdk:��{ni���s�uk��؇����z���{��ϻ���<���mƦݙ�D�%9�$�ڮ�y8 ��l�&� ���%2H7��#�	!�}g�ɌIY�q����ձ
��դ}��@-�h[���S@��M�z��A�onM�rS@m�0�m���xɺ�%6H��L��-��wJh���?w,� ���U�X��j�.l�� �܃ �L`��0$��l�ݿ?sa�X�.*�����0z�[8�u��,nNn(n���s�MN���̾ {��0ISL������=�R�X�o$�8�II4�r�?b��JeB@۶`[u��x�v6D�$�#�9�h�M��0�
d�� ��u�5��Z˲�*�$����� �٠[�h�M��!6W�#�a1a4�f��DB���_�;���7vـ|��SC�c�n׭��ebn�������<nWg���-����޺l��Y;k탒T�� ��܃ �L`j7ad��˺.�LUڻ�v��BP�^Q	(UGuw� =�z��i� ��%S��?E	!�w>�@-�h�s�f0�M'�($�
�u
"mS���Aϳ�{�O����r9#Sˠ����(��S=�׀w.��l�;�U�y��]b���5RM �J���d�e�	$�{�R����n3nq��[W	�v�g͸��xNz�۶�`�Yi��}�w�����k��46���fp{�ၫv[ �L`��0:�ʙk.ʥW7sJl�� ��]gˢ!DEPwuX��^�Z_�)���d���4��D@��@-��h����)�r���<��� �Do)��C�Сz!(QU����=�_�g�u��B?\3�K�h�z���##x�931�$�05n�`I�IQ��W���?���.��j�,7I����ͷ�����..Mh\��?���q�w{������!���P������^�h[�s@�e4�rw����L��G�[��i���f���:"%2}r���D�Ij(�rh��}��^��s���@�N���'"p�vM���=v�v�� =�x�)���3@�g�>ml�x�<P�/y� =�x������?DDB��[���9Awf;=4�5�|�U�J�&� ꣁ�w�;��SlN_X;s��$a�uV��:,Z�w,ҋ&(Ϥ�7h�u���V��#d��Z:��I;XvvC���Vw����e��.v�ؽYv#���[۸�C�2��8�{J������+�]�aT��v�q"c�)��f�O��W��ƛL;f�n�;&i�]n*���Qy:�r�n�q��w�������p�`F�"r<���g�(��)� �/a�6<��!�r�:���].6�&�����9�^��x��x�	/�u��z���� �x��RM��w4	�05we�	�1�>��5/ X\ں�E]���v�b�6w]aТ=	B�=���7�^ŀ5���W5qT]6e�05n�`�1��*:`N�t�:�+$i"~S#"�����?�fg�Q}���y��`;��9�B��6^��q���g�N�>�{qe�n�u+ۜ�^����B�n�8��$k�����0'v:`jݖ�'vckh��yWWB��*�� kŔ�+�!$	 ��� �����4J���D*����� �}x�e�=�ɼ�s���7�)��h[���Y����vx�l�Wuv�կ�+F ���DD%3������ kŀj���<��2C&E��B�h{I쎘����1�������V~�Rĳ���n�:�!p����u�mfެ�*=jK�0�?�������h�]/�p����6�&ɳ��m��9h����s49�Z��4۪ـo��g(J&A�s�U]�S7j��� >�׀~�V�-\5!l�0�8��c"�`d����8�� �١+�Q���SI5�b@a��$�4IH%�!%��c���kDu�.����c$�MT2`l`7�D('��)@��*; >��|
�'���q}P@8�T� O�"�>�>ٹ'+�;9+�(7�C�6���q`��X�s�Тg�}x4��N8� ��3@�z�hs���hwe��?�?}��8'#�$�CB�F*E�GT�3��<��[Am�h�n��u�;]�+�,��"m��<P�g�{]�h���?n����$����ŀ9}%UO��
�є����96c��07�0<��h{ҙ!�"��X(�����`��XtB��������HƜ͗6��J��v�=���� �����]��
>P�]�`ovM+��T�j��˫X�s�yDO����k���빠��lǅ��2
%y����ԛsٯ<�ƫ7�d{*�=;�7g�Dp��d��)�9�j8� ���@�.�}빠yϪ�<�䮴��Ij(ӻ���x���DU}�X�w� �f�{�N8��71��/�)�sobg�H��c�W�0%IR�[�uE�sTU�v`yBQ?;}8�����w4�Jh�y�[�!�������<�%��~_��w��k\䓊O�P��E��y���T�ty�	5�!�`��q/A��-tn
+8��6�y#��F6�ۧF�I��m�˿������Ɯ�T�g��u2�'�W���j媓r�
6n��OP� 	˰{1�)x��cM=�x4��@����2K�k�Q��Qa4�䞭u:#.���:�6�MԎ��p�A�
�ZQ�5մ�ݻu�Xv2p[R�ų$N]U��ewNٚ�Y��5fk_�` ��9a4�WS�򲴆Fx�^���;u�']�xptr�7V3�&�x��'�����,c�$������l�?mk��B���k��6O����"�o92L�/�)�yϪ��Y�y�w4�۩�r<S'�wf�k\��]��%
&~o�`��4���ҟ��6��C����~�d�����09��GiawYW77SWw�~�x�%��ל~��ƀ_z���-{�, �CM7�.mt�N��gN��e�� ���۶�x�{5�)���4�	�3#q����Қ�Қ}�?������}�|�{l��<pr�s�s鹉 XT? GH*(��׀}��`�`I��UR�AeIsd՘ ��x�׋BP���>4m����@�'��X"����$�*����}~0۶� �������"�o�$�����0	ݘ�9�1�ov���Ƭ���'n.t�v-�E�`"#�ǧqʕv�%Ḍ=saC���{ݺo���<N���_���� �� ?n��(P���ش��QFҟ��6���_z��3����;_b�?n�3�	L�4�{��)?7i�4�~���4��������P '�Df�@O�����M4����=��cn"���/1�;�7rwf0n�`-Į8F8B6(73@�S@��~̞�����X�^,Ѱǒ��t�����춺��q�;���;fE��m�|���v-�[@q����Q�X�4E���~�7c�����09��a�+
�YR�.���^,�����4
����#�~���#Ȥi��$��{fx`ow ���-�ɱ�Wdj��؊����˻0:!y%
�������$����rDH�툡U  E6�E"34��b����DUs�� >O�nJ����j�EMـEݖ��UU�Or��g��r�_?�r�i��3�5fcWl�ܓ\OJ�؍��9���X�Źw������t��������������0"�Ǡ{��cnőȚs4�]���M�z���s@.[���6���L�Uk ߶ـ~u�p�B�䒪�w�LO~t��;�]ڗV�X����佉�ɱ�{���l~ٞ0��r�i]*�]M]`��X/Ds�|��_���u�)�� �(A	$		  �}��^r�&a&d.[0[��s���7���I���w%ƅ�eggn�L�]��n�֔��õ\p2�D��o�8D\Y�lP��'���o��ŵ�w9�yc`A���隄��W&��m�{ll]���/I.�݃�uc㭹�@���)1����,��-I71��	Ǚt�B��T��=\�5�ir�zج�x��>̻'��RE�%�LҀu�pS�5�]�Lպ��.V�v�rF���a�`�����s���3��[Mզ��I��u��?�����{��lM��]�����-b���a�����A�ꤎ�O[�y��빠=�D9Q����4�ln�L��Ln��ԣ�D��A��nG�y�w4����t��߳����;���8�#�#�4�07�09��`qM����t����<�G��(�jx"z	|�vc�X����G����� M̒���ut�Y������08��`sv:�}\A6y�QՍ��ƿ(�"�p�<W���y���]��빠w�)�y�JB)�dO-P���M���:g����3� �ߦ��;��7	 �b�L��?f/������ ��V��� �}�J9�87$X�#��w�)�����s@�۹�}��#���#iLsm����v0z�\��/Dycry��;tv;Vr���ݙ�$��MDbsҐ��￦��lt�����wn�#��^x,J���8�RI�{�d����<��4�Y���IL��]u]�wr��榭`��7$���sJ���� � �H��iL^�(�:
���@��nhθ��1HL��Pnf��vـu��u���B�P�y���Q~bl�x��DPN{��9�0'dt���A�ٲ�v�ff	5�ppL1��bV��gx�w0�]��nҜn�5�Y#��R
��RM��������7f0:�����3�\�M������z"�J�ޮ����M�빠_z�y&289$X�%�09��0	�1����;#�+��殬��݅MUف�B�3����b�����DBQ�"!%У(:��@��K�dhƟ�$M)$�/u��'dt���7f06|��P������H����O]\�m��J'��>.�GC:D��ō�2HIG"i��/��h�l���<���}A��b�.���1IL ���e4�Y�^빠_m��=�{�I׍b ��C ��Xr�J���ŀv��y�Jd�"����
I�^빠_m��/�S@/u���L1��C���Y������vdݘ�����xx!�⚉�T��lր����"ED)���  x�_��T���+*/��@	�R�|/�
PCK!<"/�5T�������П!i����ht 2*�?x� ���G����Q�Ta ���j� ��e@e�u�F� ��T�x�^��=�������m�e��m   ��ぶ�e��dQ! v�X3"�{h9�hf��e6[\�M�u�@c��r�X�M�ɳbl�S��wEG]��e��P�`5΃a�J�-��λ=Xk�q@�X8���^�8���w3��Z�b�g[u�ܤ��	5Pt��k�b
��Md���ݫd�:�Ik�Nl���#;��ه��eە��pK����<�V�n�l�vM�z��%Ѷ�{2�e��hu���hw$�TME�����2t�dg�=����a�nwA�G�O�[�Z�ɴ�B�t������Fے�����w"��+���$�� m�ڴn�֌�U�ͦ����9�� �7�?�Ͼ��Z���vK�΂�
����Z�%��s����yݲ����rn��o:v�%���=vq5J��-����F~�{,��a�5T���lF��;VِH��-�ٰO�e��9�4l݁cev6uFt����׃�m�ax)[<.D��H��!Q�ua��l���\��r�2;�K ��%���=�:!�லVۈ��m����\V
%kVv�NM�M˥�@8��`�*�^��liۨ��c�̖l�\�vf��4��m�u�7"�dq{u[Iäᴡ�"��j���J�g�"�)�؍RwJ�/49̝9e��Ke�9�:�V'EںYN�:.�Kz�9��DIA�kj�RKa��'�b�m���ۡ�q@�q�౐kj�v�Zv���si"��@�Z�㇖[q�����c}�-F�����2Um��I�b
��uյ��a�m��q[;��IP�UU���y�i3�sr��'`&(j�+Wv�7\�Ny}[��moU8S���:$�Y0�2;nٵP@Tj����z�Ŕ-[��9iy�+�S��'`ۋ���	�JKU�T�I��>;�,��:(r�n��9�R�PU�x��(�z۳)�u��'Ap)��+,�m�S�� ���<�S�p<9Ӣ���4��O��_�>DB����&��T�U�|e�,��cb&Bٷ	/;���km�5����V�wO`�.�P�0��l]i٣�~�_۶����Ot��g�M�n��73ujۇN��vͶ��s�f�[z�t��rf�ȕ��]v�ˆG��/]�"\pZӮ�V��N;��B:n�U|��cl���z����)�n1��;'��צ��/V	b�S����[���&�\�-��s�QD9����&ٹ�$u-;r�t��t�K5uݝ�-�HZ�grg[�_wώ?�{��濟W:l��.�h~� �]�u������ڢqƔF)��4�Y�����2s}� ��ŀ7�r��B�To.��Qu"���������=��,��,<�B��޾0���?i�m�%ݕWWsSV��x��ـu������y�~ϗͩ1I�D(73@����O>��s�]	/���`��~���z����Tm����Y�ؓ��Mێ1�4�:�X��'.;k&���`d��0&��&�L}��j�WeR�E��Wxz�a	b�kb!$\D(�Y'w�ŀowb���z!(Q2}&�UUWr]��)��X?y�M���1�&�L	��̫.����������Т���� =������/[��=�D�(�RI��6L`I��l��� ���*Fv��<�&A	�Ƀl��}�6zGٻ-ԯnruz��0=�\Vѵ�ne܏��&� {� ��Xz�z#�P�z��ا�$���4�h�������;� 9�^ ޼Y� �9ꩻSwr+��l���w>ŀ[�6"���"����L�J]R4�D<�����i��v/�V�Ve���"!z"���^�w�`[ŀ7�s@�ޔ��NM޻��(���~��, z��:�ST�~8O'igp::���p�v�n��@��O�K�nn�rGd���?}ۑJ5tv⪸���&�Ll���c�ݍ<��F���&h������ ����>����^�s@.{j��Q�
����[��x���݋ ��ŀy��]dhƟ�$M(���������`��`�ŀBQ(!$��
B���9�*��S�}�ܓ�ϋ��� ����3@�n�o]� �l�-빠y�W�8�$�1���a�Ҏ��hTIƖh�D�۞덴�݉��xw'RI�����h�����޻��w4Q�&�v1~"D��`��:D���ϻ ޼Y�2{�|d�L�������>����^�Q3�݋ 9�^�P��uE�E�)$������h�f�{��{���3#QH�x�$��e4)����� ��XBS+���ߜ�٦�f���bN�4�dR%�ɓV��$ĝҙ�dJ�z^/k����o����%�G�ŧ=��T�R\ҝ����tp�h�5 ;l�u��U�;s۰k��y�rIv��uɲ����l���F�9^wA�[jW۝�ZBk9{mn��E�hm+��v�1��(Wq��6��4�⓶�h7n�t՘��ܣ:N6��L��SZ5�0��$���J����e����<�u$���^�۶+��6����h�ɹ�=#�u�͒w�T�]��x�x�����h�~���R��F�i��DҎM�{RJd�݋ ��� �x�5:�h�E�Țs4��h�)�r���]� ���I�q&H���ـl�� {��%�
���� ��&��,!�N'3@�mz$t����iF�������8���V�޹Nͺ��oX:{�5pvn��R�9�	�yE�iǠ^빠u�s@�۹�r���e�`�r8�G��������7T�V�
�Pާ�߱`>�V �^,SדJ�e��c$��[�s@�mz�w4��h�mQ5q%�dƓs4>�����[ޞt��#��09��Gi`�y	�)�H�z�hm��-빠r����kؤqN6�y��r�]�	���:��u������oG�����N(��e4s���4�hm��/��h���<�}A��b�˽34����h�*�0'dt��$�ݎ�$t��;���Q`"q9�+k�/u��p���$d�R�
1@Z"P��!��w�7$�]����Y!2b�E�iǡ���}o�L	�y�vGLRK`ol��)c�E2<1I&hm��/��h��@��s@<���q̑5������å�I���q��8sOmm:�\F�eC��ݺf��2܃Ll�g�}�}��r���]����s�TMEIb�1�w���$�ݎ�$t��c�79+��<��Ƥz�w4��a�"&{{�`{���ju�SsV��QH�s4��h���9[^���0�dYIH�Q )�fKz���gT��)	�s�h�ŀl�� o^,[x�(J6�;�ҍٞ�v^���l��8�Ə%��hq��<�:��-ma�{�����G�;m�h���>�� o^,[x����<�_U�dɊ<2Cӏ@������޻�+k�=���%$���ݬ[x���áDD˞���nh����2���6I3@���e�Xz�`z%�w�����#�$L��nf����z�hm��׋ ��!B8X�N�Wwh.Ȫ��0;�2�X6ܸ����b�Ÿ��6ӹ�;ַG��Z��bF���G`;;&Ghx���t�5�	��\�[s�z�#�<m��q)e#\[v[$�X�si�)���g�pUF����D�/��e*˚9$\�#���%���
�c!�Գ.�j�F[Us�����_qq�n�r)\�#X�r��MY��X�@J�I�al����A@�*���,�
�ӫ�g��9�����1�]�Mj2�+n�3��d�c�-�n���Z�.
x����0$�遪Iltڏ[Q9�C"�4�hm����f$}��s s�Հ7�y(��S!�>��VM�j�WVUZ�;�b�6[u�7�����{ɶ�Ȁ <������ٟ�����,[x�z�`�ծU��jn��XUM]`���=�$���3�/�������U��'$Ȣz��ؤ�i�ۧ�ۓb�tZ�lN��'�=G��fhQG�����g�u� �u��u`��kdN�fY�+�T�fa�'�{���D� ��Ċ��"��"*p��ϯ>�X�ŀkoyG�%	*�����*�%M�TTݘO���?=x�m��;ޔ�<�䮍A��D8�5#�<�06H遽܃T���Tyweթ������X��`	��? ׽�`w�:`O�lWMe���|�2z"i�y�ɜv�i���{t[x�P`��s� �l�AHLmLN��=��h��@��w4��h{ͷ\# ��b�Ș�����遲GLK�?W�}�G�����D(�ɐN=����ݛ�����!FXE�y�"ͤ(X����H��D}�ͺ<K��D!Q�,�$�j�A�FP��c	0�!�<RX��,-2:�H���	
�ϡ�0��&%,HI@�&�= H��2"�
m������Sm�&���hFb1"\�4���@ ����.�}}��b���<����_c�� �m"ؐ,��BBb0�O=f��d��=���|�R]oݾ�L-�j�`B224����!��"@��� <@ �R�? !�`OP�DXm,H�@mA ��ʡ�\ )�7ﵿ.��}�[ފ�0Ĥi��,nI���_����>��e�X��ߖ��2�t+&�䢨���~t��P�:���o�4��h#�����F$s�iٚK;k�����d:���ܝv/n����������1<S&6I�^�h�w4���%�C���>i��6UM+-U����`n�t��#�%Ș�1��G�IU/�S6]Z������X��t��[ �&07v:`��+�JBdjbpnf�ⶽ �l�;��i9��=HF5�R�H8 �vg�>����<�(ڱdxa������ �(��~_��݋ �-��>k��V��s����sv�βrkku��j�r�8�x�E�D�mz�T:�1ml�y�ݎ�dt��[ �&0ۗHB������*��� ��Y�^�
����X��� �׋=
"&O���raND19&h�����f���s@�n���.!�x�Ln)(���xo�`[ŁС%�J�������g�n6�2Lq6��@�빀=o�[u�[�אA ����O��T��"[��k��on,tw`u�m:-��S�v�n3�3��qϤǭڵ�}�����#=��i݂�;;EU�c]gp�s���a3]:ٮ�kLr��`e��tч��pvm`��ը�<��۶�F2�1��/�\[^��{ N(�1��jg!@z3t���Ig�Zy� ֳ��<�����.�ͮ���rEal��]����������n+��1�FȆ��n͓ͻڜ�s�a�QLj���9�M�z([��o����08���&Ɍݎ��
��������x��ă���[~��/u��/���# ��b���vL`wv:g����'�0:��l�r��F��Q����s@��s@��-�佾�0=��E�e�V��+��`M��Ų[ ��ݎ����oϲ��ծ'�癗�8lv��M�١z����@tv��G�}�Ǟ2�Ok�a`r�̮�=�`�c���n�L��ɍH'�d����ٽ����� �����`�2o�9�rO�����ֽ��JQ��l�2Dҏ1����7c��lvL`P�(G19�(F�h��h.���٠{�w4���%2L"���`ql�������6O:`M��������~���\��w�Qĺ�W=0nĞ uی�Ɠ�γ�&�J:{m�]�_ =��0;�0&�t��ob`{�J9�	ɠy�페[%�	�1������Q@+�K(�*j����,�\�j���" P��V��e(0{����,�̦���'"��4}}V�_m��۹�^빠u�l��sS&1�\����<�{_���w{�ծp(T��e��H�A	�ڟ�0��������spܽ����'���tb��n�
̸�6-ZYy�vGL	�0;�ؘ왠�+J�n~�������'d�;#�꤂OW�]bYY�bʻ�^Sv� ��쎘v�h�(�udXCɋ#qh�٠~��X���q��+�Q���(!8�S�{�}�ܓ�=�[Ԏ6��J"	'&���h�����;��h[f�޵Zo�+pQ��&"unˮA�a®ۮ���ZM�y�v�1��˴��d�Iǉ�b�䙠m����@:�4=�s@��e�&�C2<�`w��0�c���d�����Ln@jd�8����M�m�g��y�v���Բ�*��1bYy�vGL	$t��oba��{e>ϚP�cs�p���-�s@���p�� ��x�� !(@��J��=����;��j眠����yn���#�n��L��Z�o�wb�5�E���9�W&-IQ�8`�x�N��
�wX2ZQ�끲�v��l㴳d�YҼ�,����eb�$�K���;]��RAw^jΒ�.��p'�'[�=Xp�>$�7^��(��[Ym� �
�s�`���݊Zpvs��σ��q�s��%�l<p9�����>�ve�[k�Gwww�(!��m��$��o.f�S-֦)�z���si��^�q��lB`��6����Y��Gr�<��&Ln4�P;��h������%�C�� ���Mt���JҬ���$�쎘$t��ob�H�=`�j$� �rh��nh�Ň���wi�����>t����blX�I&hm��;��h^�@����=�6G�dq&G$��z� ��}���b�5�ŀz""�7��7]��Wh����b�=�5�rq��y��2򼤚62nnMt�p.a��kd�������^��ŀko�I~�z���߼��(BV�^f096:}�xE�! �$�
�@��l����h�� �8�ZR+�W�e��H遽܃?����~�nhu�	����9�{��&096:`n����˵qV*�B�W� ��07dt��zS@�U�0i�RA7 ć�n�����Y� ��x�Ƈ��j٥^��ۄ�"|�Z����+XZY��;��L�07�)��f��uن7M�)$�vGL��L�L`rlt���)l��'"$�4��Z�i�%�DBՐ���)���b�;�b�>z�cL��5 1��{m���恻#��M����%y+�P��fQ���`rlt�ݑ�{{ ���o���;Y�&]�\�땎{=������N�c�wl]��oj��w.�}���u��
���x,��'�遽��vI�M���r�y$���f�������}�c��t�ݑ��՗j�H��%\ݬ ��x�
�}��zύ���&҃n)&�(P�^I$�}��`��,~�f�IF��"!�J3f^����Ub��R���L�07��`�c�f�y�abo$q�25(f��l�W��[���]���67"����NT컊�ӡ7d�L�;ޔ�m�@��������%�w{ �ެ*h�wv������w����>�ذ�b�7�x��J9>K�1!'��j94~�nh�w4���ym��+Q�������MZ��$���~X�ذ�n�=>�~�4߳�O ��Nb��d��� �I%�w_�ou��Ջ �DD(*��UPU�*�*��UPUj�����T_򪠪��UAU�@�+��T$P$P�AP�BBBP��P��B�T )P��B(��EBB	P�dBD	P��EB ��P�@T"EB*0 0DX��T"EB	P��T �aP�P�P�P��`1�@T"�@T""��Q 	P� @T  �b*@T"@T"�E��	P��bDT"@T DXP�$B DX�P�1DX�B A`$EB"�bP�#E��@T"��"��T  �E���Q$B0DX�E��BQAdV
�
𪠪���
�*�UAUꪂ�UT^
�
��PUҪ���T_򪠪��UW�UPU|UPU�b��L��z��h�п � ���zλ ����hG�  h}     � 4h  ր   ��  � UDR P(	 ��� B�B@J@ (T�� �    (�� ��H�  I��(  P� 3`{�e����ް����mFMz݁� 0%�{����}��}�{�)��a�6���e{��7w���ѐrdB�  @ �Q�
�m�HzM� �Cv��7p �$��9 '��H|pp`2����� $� �d x8� (�@3P)�I�dzL�{ � ��h� ��=<��`=�A�@{ N� $2����	�s}N@���  ��EG�� 8	=�� 9 ـ � A�  l � � 0  l  �,����� p���0  6 �
 ��@@ $ ����   ��� <�H	��݁�p ���:�zrڀ��I��a��a�a��.|�ϸ�pOn��{�N@�����y@� ��� (CBM4��2bjj~�ͪz���G��h�l�RT`     Њ~=U(DP �    "{J�� h   � ��e'�J�4      M��P �    �~���ѽ-S��K�9�<�����"������*��*"���@DG��PDj������0� �������P��2 "21�t3�}�Tތ
Å>�*�]g	�Kކ�)�3� T���S�D���!7����"���(
�ݹ�K�a��%	v�f�M�L0����)��F(Ρ
��Q"T���\��D��CN�`xC���vq���Ӵ�M5�h۱�]f�M]]iܸ&��;^C�Y�a�H2�i\�Fr����G�o�1"AJ]�	��\B%uu��&���7���-&�%��޼0#�
��Ǐ�<��q|���D*k�:Ę˰�	�9O0����]��!XR#cR�LI�֬�xK�<HHB�E�,�,�t`WLײNk��Y��L4Cq
��<yM�=5��ˣn׏�jh�o<��4�0��l��F�:�f�0�m�Ґ��� i!t5�fa.h���ذ��\�/^�m�+hy!R F%e�<�2�3̾�R x0�
0�ji�H�caM;�yMo�m1/���bHV$SD���{��Y��� Fp\8w��3�������C��wX��A=��)�u�.8���t�h!e��^,äfx#�֘a3���=�e�51Դ�B�H��y�s�wx'�"Xz�a�{M%0}�R,]��b�4�Y��P�"jYo5�����H� `2�D�A�@a�Zy��NBeZ����W6�jCg�1(0�H���y���.�fҘi=�0��8p}�%=�a��4E�.�=)� x����BYv��5��$���,)�������{�tnH����6�s$�{7�������X�L���f�t�y�́)�<�Hc�|T�!aR�f理F�1��
B��+� �X�H�F0"�<|_d���!��!+��M�䌐� SC�ԉq# Ё����@�L��b��xƣ��i�1$��Mnp������1�))��;�~�BD5�:!�0���{說]"iLM�|7��Y�X�D
F�Fd9	+�`� �tB�|֌e7���oy��;]f����<̛H�4�M���޹�|H&	�% �K�U��O&�K5*j�.�A�&�X�2R���i#��k��@������Fw��"$H!F��CǄ:�w�}	,H��:��4�p���v͒�>��g�>�6t�����q<�c<Ӂ��o<�\�A�l�����ǗX1��X4M�1ؐ+��7����O�g5��F^rf��&7A�!YVB���!a�����ד3 ��
B�K3|��tt���V\��+
K�]2뻾L/=f��͓|��.�!)6���]��!���_|�/7	42��B�)1qvN�T�GYMEҺ�>u}�)�̪��,=�]��o���T8��l;p'p�0߾�7��L(�"X�p�`���sl=��#Ä*H���$!�� q���Gcs��c�(B]0�v�n�4 @�y�� h G�Pt	�*@*@�(��D�q���#5c���0$�o����`በb���WS�M�P$4��!t;"�4���!B$"R,`8ƱX�F�R�&�R`,CQ)P9<�|a�nB�j,����G��(0���BO<O9�i��2b�0����GF���i��:���>=���1ڷ��R|K����H��[$E�@
��nj2l�Ѕ"UH5�댦�b�#[�z&�c�`V7Z�dߛ�M��i��y����]bѠ��q��v� ��]G��+��a��1�6�,����d.��֧4]�����S�O=���PH�"El�aR1`Ab@��
F��
	t]i������.��2���%�HZB�+(K�k�`'q� Ny����@8܌�$H�$�4f�� ��!X��F,D�Y$y���[����[ap�4#5�5�3�6�%�/y� �Gm:�c��F)�fMf�BBIf�&�"�$8�mLc�(�h��WA���= Ma��AU���AL6����K�h�+�]4&��:%L���H�
,a
P���u�Π{�\�<�*�FJ#@�
JxB�h�%	XV��.��7��'�/�̇o����K����kxЏ� \h�������K<3ܳd��ܦ�ҕ�7�&��b��Pp]PcRiPmր�y%�*�Ĕa@d�pd�M����3��.�����%R-pe�8oQ�� +���4�&Î�%]fp'6n�O@i�dI�!T4a�Ʀ��[p��i����L�7��{�y6MM\It�}�f B��+/l��j)���� U"0a��aR\f��4°����
R�HjSR��CI�e��`���Y�CF5)�2@�����$y�	bD`�N$B*A����/���E��.�Ê�����w�ԗbE �����V R0I ��0��,|�'��, t��D�%XS��@,��!���P�Mf;
y����)�J)��0jĴ׆��4008
�p�`֚�fc�u�g�xj&'�.�- 1���B�I&�\��9�b]WLB���r7Fj�������C���)�7�(�!����	��k���l�&��-��C@)�D�*h�e���>^++� J��+�����o�)�I�
so5�@e�P�
jU�5!`R1e��
BB1#�O �0|}IFP�	HIYtamx>���,,��4+�H �����y�hnQ<r��!.�|6��$;Vk�.`J� @���R�����^�����x½�	���K�i�:�ks��J��n��!q0�c1��$V���4����kf$c�4�`�)��s7�-x� �C�@ؼf�-,)an�����(��0��E�
�C�*�`�1�Gq�)\-qET$>�4:C|+ۯO3��3���~=�~��W�>@                   ��      	      ��   ~�zm� 88��m   m� $ l  �� �� �  �p�          >�                                                                         p�,��n1�U��mRv��TpK��	m�[B�sdP�yU.��������h�)8��+��\g;vvj6�qm��+�t�a����u`�
��:X��{����qDʬp�σ�k)�:^i`��v��iÎmN-�L~>w|i�nȵʗ�U�y[�F���ML�4�g�u�e&v�vKx�ȉy��ce,�p]�D���հ}��l�l����m�D �Xؠ��P�]�MiקK����o-�6 �6�N�    � 
��V��j��w7*��[6�Mn[UJ��l0�:{4����
f檂�5ۂC�m�5R,�6�[��yڥZ5�N԰W6�*��P�*�J6��ML�$ -�l�Rf�b����@	 ���M'0[m� �Vܶ�p�ao���[��ɪٍrC׳�}��6�m�˭�      �@qm��8�e�H�$m�xж�p  ��{ﾽ�l 6�-�k�B`*�j��+[:�m�ѷ8�d��]. [m+b�kl  8�g�G�-�әi6r�$�)%llC�[@ [Kh[F� �kia�� �6��
��S��fi����P-�`����  -�� m	 m�'M�[[UI�A#i6p �8�#�H�.��H4���	��86Z-�m�  �U��u[��ݰ[��hGm1����X	V��[��f]��@Ye]#�T6�kq\ �M��mm���j�`-�  $�h��i�ԃm]%\�` �[q#�   �[@m�� �v��Z�s��m�-� ���v�� �mm�P��e���j�l� 4jz<�6���`��ku��c����c�t� M� 6�:H;l۵.m0�� U*�@[+;Al[@ i2�H�l8���[#$�e�����n@�!Q�[vSl�����f�Uj�� [KhHn�,��s����ZRg�
��V��� 6����oI��N�lT^!js5uԙ��[�`��   �M�Jݭ��piv���6�] �Z݃����ڠ��snx.��s���Ksdˊ����m���i-Ƨt��N�v�+k��e{L�+rJ�9�P�*�]mTZ�����(�p�UU�, ��Piʙ 	���2P#�#m�f�h�a�   8�  �*m"��m9�Z�Z�n�`)V�l�v��l����«UJ��vQ��� [�$H6��6�طyz�5����6�YR� l�]���d�Rg��UuUpM�^�m����d�$R���`�hZ-M�A�����,2�H�m�`R�R�8���UR�*�J����VҼ����]WA�r�V��n�mr@n׭   � �ch� �����m �"��l�`  �m$�� -� [Vq��к8�'N$�0-��s����{_,���(�T�A�Ռ�\ù�V��W������)��K�HÈ  �` 6�uԬ���6�մ��.B�hluΞ�Eq]lv�5�ɵ�ًkdɲ��M�   I�����u������кi1�lH��I�X$�#$C� � �nl�\��Ö�J���x` �^�$�����V�i�I6�2h�[l $��     k3��ݫi�2p�-�W[vͶ��u� �/K4V�m�  r鵒��.�	� t,�Ѷ��� m�- �۳�m[[v�k1�@mU]U!=@���[I ��q �p 8�Mk[Kh4PH���äm h<�i��פ[m��{����$������"M��]�,���m��Cl�� [H0���hIg�%���m�ݶ�[zŠ��I|{�����&ٶ	\a�Wf�j��W������$�@[V���Z��e@eW���V�2Ʌ*v��s`$  4Q�ۛ\6Ͱ�B�sŷq]R���N'��C�����Z���%��^{g�U���a��( �[t��N�@�-��t�\�`�l 	 [W�H�q�Ŷ@�"��i[�U��s�:��T��/[.FB���Ӣ����5Pҧ\����u��|�Ф�37:;P����N�:H'y�6�쭛�St�nx���]J�UX��0[06�T�m�z�zK��� 8j$�k*�H ��&۰��M��%s���͵�Ė��$pm��: � ۫v�`�U]����� ��6�۝h  ��}���׭ �pM0$ u�s#m�@�   ��� Imd 	 ��V�6ٶ�� ��F۰rt����� �8� Yc[� [@�h-�l     �l [@      ��d� �J   6�kX �`  m�!#[D��IJ���� $l����� M��\   m�m�bN m� �Ԁ  p[\����l   [I 5�     $ z��Qm ^�[�=�若8�e�@ @��� m���8q�m�   -�   �-�l�����M�`8  H4k�ф�2;6�`  @    ��v�     m�O��@p�v�ʹ�@ [@  8 ��L�-���m�	  [@  -�        -���  I&�  ��n����`2U�Px���V�Ē   H�@8��� 8  ��lt�S���CM��d%]۠:tm��]6��� u�������o}Ǵܛ	�hֳ���l�[:\�4lp�vkh���p�di5��i6HT���+e[.�5.�]+@-���;h��1��Zm.h�  CZ�2m���.�H  �[��� m  n�kRI�T��f�f� ����͙� $� �m�  -���%;#����mw:�m�m�  �ݷ �[d	6�2ԙ"���a s� �t5�K� �pI�m۲@I:���� $�h�fڃU[[�V�쬪AO06ٮ�嶕'��m-E�q� ��qJ�����j�wml�HÀqz�m�Σ,�&f� -��;�d��v��Ӏ.ڶ  6��RڥZ]�d�-�@AE�U IT8�+h)��/Z۶�6�]��<k�����U궫��Bʻ�9Cm�/]m�k�i6�    m�8r��%�6�[@ �6�c� p���kH  6�  �۶�M��9�p�Z6�  :�$Tme��  $6Z`�kZ��Ar�a��·��ܩ@�P+t�ls��LlP[Az���	 [N �j�-  $�l �d��K�8��xw�x�";������~�P���̊f���8W�Gp���:�h����:��,AR�QD=th 4�t�̀x��рp��)�Pb�b����9�@�q C�C�T�/�l�~�G� ���A��!�_�t ���q6��8"D = b ��� i\�EV$�� w�P����@UD��E�`��OG@
�T�C"�C`꩓���#�/^�C`���v�x�!衈����C�UB��Q�-9�S`�@�_QG�tA��5P_�h��x)�����[R-]���i"�� z(��
y�lW^��I�)�=*k���T�@\���aTʎh �j��ȒO��^g	"l �5 �X
���#R*X"QP $B
�UX�y�w~>�gO~�    ��"��pI��m���`             K"ե&YT-�9{Wn�f��h��>���#<���ـ�Z�ԕ1�-�b�ǝ�n%�T�:-���mn0��ێ�iT��@������;vq/2���NKcj)T�n������mNb�6+��j��jP�RsT�� �0�wY��V4�-�dƋC/=j���'���"�p��O`Υ@J;!�ql�u�h�G��v���1D"�Tp�!nvD;6�6���Pt�l�\Rh���흫���m�J^��JE�!µJ� ��Q�ʻ)u�9�c;"e�U�f
��/M6ސ�\�;(�����ўD��ts��d���EZ�2*&����N��9�C��g���oQ2���Bڹ1ҽ�j��Q6;�a�4�t;7(�l�'���d��Y��%e[�؍����X��ȹЯu��:;m�6�d��tƊ�f�X5J�`3;hݺ���p�r�lKȭ��Lx�*n�8D�D�k/m$�Y<q0:li�P!�<�-mN������lV�pr�AnyvӀ���������m�V�
��c`|�F�<��N�ݹ�:�[{���)�ķ�a�9��u�0�5R�[-@PxY�mYdV��e� jH��x�vGN�T��WV�9�y���y�� �[9����چ�)�+*bF�N٩��B��#
���E����wlm��F�����F�0���C�IӅ��Ge㌆*]%UD��$FǠ@�{jl۫��Б;;��܍�'SQ�����}��s_��� (	�;8�x&��5��8p=�@=Q�;���h�g,浀 �xi7E k�7�pCm��+;ͱL@��7�11�l0�X	�sX�^@�pˢ��P8�ݭmgb7�jq�݊DO�#�����k=ttr�6�9�r��V�P�v�݀�[��t���sqJ��vL��:���pC��nH�����׍<Tܱ�La��!���K�R�kMֵItH�����#�x6��� ���`��y�FY�?k1j���Cz��ڢ�E�Xlj�$�$�2����pܯho}�׾����Yc��Ih}p���oLf�94H��x2�����Cy�4�ɡ��[�.��k�v�yȀ�G4>�is�>�ǟ�x�	Z�(g%��:���w4�����n��hS���������wx�+��h�is�7Ѡ�%�1����ֳg=��x�Hl�iH@c�.D=>hw�h�]�J(�����hָ��6��?��:_ƻ�m�Ye�h�G���G4y�4��/�X+J젊8���;��>C}gTqn�m����F}��X���v��tW�ɺ� 욋1b�6����)ZZ<�\����D��-�aC1�"���G��Z��C�Wi]���z�`��`��p�8��>�����.� V =��w.|��4�ܼG+2�C3�;��>C}��f<�ZA me��э�9v�9zi9Υ������z�H��ņ���%b�1Z5��C|���<��%�k3-̴	ţ�2�t�<�\�/���H�As�wI���͡���zHNBm%c�R��y�4��7��^I�*c��\�������|kS- �°�5�D7�3^�C놾�*�o�U��t�D*0�:�4U�PS���.�h�b���{D�A�Q8���ܢJ����_]��g\4��8q�b'
x�+�C놗6��h#���+2�C/��.m���G��BQD��]�+F�Ȇ���9����[v�2�^bD�Z=�{�����߸y��s�|� ��%Itx����""Q���i4hX"U�V�BJQ���j�5S@��M0t��r-�����������F�  H���Wj����<k�ogV�/K&�݌.gh	��UK�V�����&�� u�#��ɮ�월� �3wce���8��g��n���zz�G=3�۵Ҷ����v1m\ٮ�m�;)�mV�;PS�'RY�J��f�'�Ǭ]b����Mֹ�Ol�1���c���(�F�x�WG"<�Cj�m���Yͷ4mqm�CNS%9N9
"��}{���V����4��Zi+���ţ����4=�Dw�h��0�@$QC1�����;����C�+)]�
� k��x?�y�4�����(Y�X
��9���ϐ�F��wl��{��bw ��%�I�U�v��|Qʻ��$V��fRYhe���p���o�C�B�o���w|J(�K�b�kdiP5AuU�\[HrMw>.�K2�e�J�ţ�"�9����!����bI("�%_E���:_Ɠ|��������J�
Ѵ�h�k�U�G���@w|�~����Zk�fwb�6[#�Cag�ۗq���5 [J%B1��!*%�܊�Ǉ.�7D�{��.͡wy��+����~����u^׎Lˋ�]�G8��h�%w�h�Fh�5v���t�x�+2��Xo��&������	E+���ĭ������?u�mN���b�ǵێՆ�wl��+����9�80R+	Yx��qh����p�o��|N5��F�����o��l���Z����?I*
T*G:�+�&e��v3]���3Y�H�E�kdhk�q���ݙ�S�R�F�Ө�/2<��vm��X�G��i�&�u�M��k�h��"*>UI���T�|q�C�Y�l�e���u�Ĳ��"F M���#M�4{�o�����\�W��Ie�7�G��� (0UP&�����@7��<��%��B�1Z5#hk�mɣ�p��v�+	Yx���4zH��rh�k��/�Ʋ�H�A�nM�w>Cg4����o^G�-�  v�muBTc��3\���'sK�����kRQ���&�V:rc@j�2i��C�7��:�+����c&r4ƣ@n��v�<���튴:n^6�͂u��3��c��	�ms�vō�=h�+#�"u��kuJ�rn���[_��}�2T��W˪8��[Q�^�FW������.���z������1��� Osz�8��v��vi�Չ�8J@�J�F�����|����ɢ7�a�8�h�8�7��<ܚ=�{���6��f,	ţ����G����q��b�,1����k��9�5�&yY��W�G��� q��� <��Gq�$B3,�e���N��n{uV�]l��6�Tj���s60e��\�n45�;�ܟP�����d���u���kg>��d �T���*	�A��@	��놛|�K�q���6PEf%tܓGu�M�!�ۺ���M��U�h�X�{�o����nM��,�U��b5$hk��rh�k�\\\�5]f���Q�m�0j*(o�Q���c0��8�wk$ݩ:��d���nF���+���͚;�m�=C!"n�XY���(P-�Ƥm�����U���-d�͞y{}����E<�� B�� ��
�ֲ�c$%1�CFPȨu�� /�J�"�M�rP<E���"衉ᡰ�Q��ᄑ�� 0"D��R!1�HB1��`F##�a�ZM�;#1�# !���b�A%#pw�f�-䮔Cp$l(�Sʣk*�<�q��Jfq�Ԃo��g@�Q���IT�x=�$�/q@,l@���Zg�v����7!(�I��hӍ�����G���\̑�V^$��f�?��&��6��P� 1v�D�o
�e�
̑�r5h���vz�}+\��%G%v:�RcV-��O�����!�z�6�YV�������o��F���ߝ�>J���"������ho����[����$�f�G�D7&�;�H��)�#PD�������0�}ߦb��X��������r47݀.>���D��N�`)<�cT���}_c�V�4���	JFJ|m9N��ϕ�i�̸���%nI��r�+X��ĭq�7͠9ɽ_eiϬ��6ӒW}��z%��{���}�z_լI+)��9&�;���!��=	�K,�F�Ib��p���.������{�TB �z�d�M��5��  Nk�Gl��f;`���9�>!َ�t�S�t	�{Hɞ�p@���n��0Q�6'�$���7ں¦2l��c���͔{�Ͱ�A����9��8��uqY�h�sq���~�|��k��*�n��R�g�fF��X���'�-ON�ݬ(���窊���q��y���w�ԕdפ��f7��>I3������b���'+�͘��A�hEa�j}�!�m��4y�4���(�'�t�nM����������X������o�ލ�	#��1Y�����o�ލ�ɡ��	Ei`��V�9͠9�4>�y����t�DJT���JT� )�@3n�v�n�lv�S��H��K�;;uQӒW+�z%y��_ei�$�B�܊�XH�9TH)#�sM���~�7Ѡ'�.ie�h�)ZZ<���}G��Cj�r}����,���T�Y�#NF���7&�;��}e�1f ��qh�H�������7ʼ��7n��Ku����7Xn�`f�ۍ��7'-v���7��0!�]�+��ɣ�ˮo��F���b9Y��A^-.]s|��47&���*�*��w��t�ho�T�W��_
�@ 5�Ohg���m���Yx��Ś=�!�nM.]s|���/-bX��D$�5�ɣ��>�r4;�����N�Q���T�$D��*��s���kb.��l9:��T���BWh��Pr��Y��c|���f�rh�"Ù���+1fZ��5�t�jI��<\���QGfa�1f ��qh��|i�&� �>��4;��aC���i" � �>�G��o�!]���h�	����9�ݟf�k�(���Z<\����G��m�6�%��+��M7�}�}��Uˏ�Ϊ�b��r�p&�qu����w���T�Rt�%s��ދ�fD�3�߭a��_�{�GN:rJ㏫��ĳ3w����o���%���+��	,@6���双���� >�.�K,�Wj�ZZ>��W7w"��������^�?:tۜh���]I �MI��<\�[�%����M��  �w%S\�pe�A��u�~��:1�;V�j���糺WsB��n��=�$�f�a��׹�N�l�Ҫ���^�^ۓ`�٦��s*{b���n�V��Xa��A�5v�%�3b�Ҝ..��㇉ɢ�vL{\�:qV�e�\s��V�c� �7YU,@-����ww��{��}zE�[���["gg)�/*wFw��};��6�+����|��Ea8����@6�����D�����P���f�]�@6���
�*��ԑ��������mIT��HS�Vo���sK���3�ՙU�%A8�'NR��{b�֕��:����>�06JrJb#��kJ��:��Nfe���2�QJP1���GK��c�7X��B���ޒ�L�$u�MI{����ض�/ �}��;��}���᯽�f��*չu�3g=�O}L�	GNa�	R��;��Xr��:���M�Ɖc���7�� ��I1��y���hbn(F.��ؠy�]-� ̸�|�YQ9TS�Q��37z�����7r(�Ƞn��^��*��I���8 �%�Gl�{st>(U�t^�S���[� �]�z@=�����w�����jT�Rt�t܊y%Ĺ�T^�P�oW@���\����������I�oF����	U@Un�ψ�� ���GRB�6�@���t�� ̸�ێ���QR:%J�NG@��ˊ }��{�]��������M'\+�s`q
`���J��=�%s�4�R�AR�NpD�1àn�P�� ����c��ʔb"���8�{�w���2ސˊ����5�����}3w��e� � �� �nRU>IRA��[���0�$��$�0&��R$R+H2� �
M(��!
��c���t�Y�G���P�� �� ����c��]a]���	��l%Î�n;U�������WS�����#��j�Jb#] �� ��:����h3r(� �H�8��C��g���*��� �Ƞ׎��x#�GA�.�x�f\P�� �����4l��#U*Aàn�P�� �����Ho(��B�����y�]�� ̸����Kx�R���e)`B���Đ�.�LHO���h?�x�\*Q����"$$X4=�hZeHHA�z��ŉ$P�ZA=���y&	!%�"�H�bC��D�!I���b0 ����+E�I��
��I�L��R���\�C<��{ݦ&�		b�t�0���!�0`B,Pc,��#I ��8����,��_6ߔ�  m� H�Iڵ�z��  ��              ׮�rɚ[����o[ �8iVGk� ��]�OU ع��9aN�n�v�t6�ܧ[+ԯ4��^��Wn4܅�7�h��ϛa"9���v�*��U��֕qv��:�ʐ=� 1E$̀�*�a梪�U�t��R��%U�B��K���F�lRgn^�R�.6CL�-.S��Z�WRl�uv�:ʧ:z�O�S���,` ��X.��<�;i\[	�+q֪��>^��p�d]�'r>8��x0�������� -$%,n����2lqj��]�WQ�����d��'F�nH���pxZ����r�eP�9%���Z�Bu��S�����s��m�ӵ��r��}��z��vQ�K6�m]3�E�4餕�J�&:t�T��	�gGYp��=�b�� �si�\b�K��׭r@��:�����*in=�J\ܳg���*�{[i����t� �x�8l������3��c={u����k�Y�����k�����1<�;�B�WV�6
�U2Fv�t�[�iV�z *�)v�z` wm��s9�U֥�`�<� �[q�عa�av�����<��DP�=K�Ғ�ڦ���1m��R�M�6� &� �8� �R����e�n1˳5sm��eكn�݄H.�\�t.���"�Ft /T��*�Wj�Cɹt� O5B�;V����W<p���mp�St�N�S��kYX��^�ȼ��إh������Cm�(ʲ�Iy�˻��c��O����F�G���w��]��٘�9
�r�( �\��Z�y��_~�����#m�  �.��Sqq,�]��;�c�r��^F�c�f�K@����JGK�aj�m;D���:lӍۭ�6v���ed��b�t��9*ל]�0���ɏWg���r蝭۞^8����+�."�i��h%V��WB���c���xx�l>\Ɖ�t�uRϦ���{������]�����v�&ۅSt�q�V}H��M�.{��l�]i)��j)*�r�q���z����q@�\��eIT�$I���I����Ƞg�����2��*���UMʇ@�Ƞ�8ys�r�3���7_��;Azd�������@7|�y�]1����[�� �d��H!�}3���=�<t܊ ]�$�?~��_^9ӷW-��p���|�nq9�p�%�.�FW���
��#T��E���2�~~�g���{}��NrR�QG���J�$.	Iz�fk�f{z�c�?q%�ʣ�ښꈥH������8י���V��@3r(�;�q5�E9M���[��ˠn�ˊ�q/$��� ����%S�U$��f?�ˋw:��� ��ut����u�T��nSX��n;����[4w<�1NP:f9����&��So��Sr���� .��.��_�?$������5OA�NIL��] ����37z�k� ̸���..6g힩*B�A�����]	��ɲ�� �~Q.w��$��>�Ձx#�F�9$]���O}���ؠ������<��(��:�)�J�1�W7�'W��]ﺺ�� +��UF:n��B�S~��a�8�lN�Qn��$��\Oj��~O�����ӳw�`��]�ut��˝��ȧ�q���j))���7{��^= � ���ܪ>�i�%>F��8�k� ̸��� ������So��ے���{�� /u�.��]\�]H\PF�b�@�KP}�U# �`�PI� 4��Ϧ~ �z����*5�����ߗ�^�ˊ��ULP)���.���*P�f�|��W�z���g&p�#.�b�o�^n�t�� ���ێ����Q#T��E�>Ǥ�Tf�P����:��V�479)T���@�Ƞ�8׹��2ސ�Q0�S�)�����^gW@�z@/.(�;��j))���/7z��g����@�8K�Kם��Ur���Ŵ  	nۧ�2��k�nN:�Tv��S��4$�:;u�e݌".�h4���"5n����[R�t��*D@��6�Otd���Ϛ��#�p�&��Є�w[�/��ͷ�|��dȕ����p�8��9��tQ�ɩ�Y�6����.3v,6��>��u���tL�d]��	��=�ڤYN����gelP�����������Z��k�@3.(w�������tU���T9U)�w"��Pfk�f{z�c� �S �$�QQ��fk�]�utǤ3"�^��d�r �M��ޮ���fdP�\k�5$U%*Q�"��HY���޸��W@�Օ�:AQq�� dAN�{�ls�]�\�;��8�v�f(��ގ�QG���@�p�ޮ���}yD�)
������ⴺ�\�>�\��$��%��� (v{��10��)���nﺺf� �Ƞ޸kVa%>8�)�S��f= � �����?|�����㊡*�3�f�P����oHW��+����6�{\�aϻ�YY�"[4�IzQ��L�¤)9%9%'UQ��f�}w�]-� �Ƞ�#���H!���oW}�r��~ � �c�z��CREJJ�$r.���^dPk�D�/q�>����m����8�*(��3v(y����t=�.%Z�� ��SP��J�.�g��>�ή��{P̊�ī3�N��j1�n�k�Y��y 9��Eېݯ���tu��g%��4�7}��2�jy�@�p֬�P|q�S�S��e^��"���]�W@�Y���8�J�:�� �� ��z�Vm@;e��rS�S(��I%�����I.ܴOUX]^ 
�)��wn:��T��7�33z�Vm@32(w��q}���)��&���8�c�q����R�Nrtm6M�6svT�Rr�r/���T/"�~p����nn�6:qB!�QànlP������H׊�!F&�B��.�fk�_ם]<�9U��@76(�;�q��87n>������ �Ƞ޸ի0��ds�$)���h����'�b$��h�H�P����6����  �����G��x.���(&z�h�*�N�
��"盞iL��;(�8s����념kK�Ҷ�cu�����K<��o�M�Շk�����4�+׋J�H�f�q5C��g`ێ���B�0��v�a�-��ٮ+`]�ss��u��9�y�U/3�L��4�w���|?v+��afݽ_��w�.�1��,]�l�r�q3���3� #��NTU	TGVx�����^= ap�I�RuQ���p�3��^= �E �n:U��r� ���^�W@�z@3� }z�Xf!�DӔ(�tǤ>Ƞ׮��Y~ߗ@��E��C����@������H��1�~����^�Ћ���:��ctgr�6�w��::�0�R���A�_ f��/�ή�x�@2�(��S�rJ�7n>���f�P7�Z
�B+F(�*�/�{M/]e����-$��m��T]~[���#��!N.���@2�(~��fo� ���](/?*m9QT%GL���Ƞ��WC�IVl� �L�HӒRuQ��/=˜�^o��3_�^E �]B�QJP&S��X2c�Ɗ#�μ.�7�#6n{tk�J�=���'X)J�����utǤ/"��9�~K�����~��p�4�
8�]�� y�ؠ��W|��=����dD����P�"�R�����}8:Ӕ$)����3Ap�:�o�CP��#6g�	�� i��" ����L�� �!C<��J&�X�"E0 �!2!#�t����XD�$�H$ �yY���� �
��(b!�h��SH��Q ����<S 6
�H��c�R��_Et��gPA�A 6&ϐ�g7���=�]�!���A���U"���^utǤ/"�_����!M�T���Ѥ�y
$�h"O� �?�B�>Wo����u�I��m�
k\6Y���z9�.��\Wk��o򮮩�Jl���
qX���e�P��^]���ut�+|�iʊ��t΁��@>��^�tǤ�>�&�R4䔝Tmt�E ��:�jUY��sb�}�q�IJ��������H^E�׽P�3�DԕPr�]�� �Ƞ^� ��z���������uE��,r͇j���ܳ'4m�N��Ϣ��PTQ����Rsb�}y�����HהgxE
IT�E�/6(�y��/���;�GQʂ��qt�ޮ�x�e�P�b�}KVa%6A��8�����@>��^�t��j��**R�:�� ��$���t��W@�~�$��z�B$"Uj�X"�H�T�_w���2�{x�m�  �/m9" ��k���y.iS�X�n�V��5���8\�������v1pU�@�s�t��P �Qtǒ-Jm�v��$�����*ݥZ��sV��
��ύ��MZt���61VNN�:�6�Ҭ�4�:��H;\�d����E������$��of̻�SY�uM�oW%�B6^8�n2�����22�u������x˺� 4�nF���UV�ؠ��W@�~ y��I9R
��@������Qx�nlP��2����	����H�k���C�\�UW��/=��=��Sr
T��@�ؠU�@/�tǤ��3�$��R.�u�P���� �Ƞ/��?m�v����G&���9���v�ųTU������R#����㎣��2�i�/����^��Z�F�8I �:��E�.%Ƹ�͊�~��s�@�g�mʊ��t΁��@>�ʀ_�4��Hp��nF���U]U�F�s�u����e�Tl�� ���@�ɧ@�z@2�(��~}��]mk0���exy��3�]�Ѥ���-�]�r�U!�D�	#p��H�E �ސ��:�Y���"����@>���sN�x�}�Fw���GT���H�s�s�K�@�j��1@
�y��N� �=��e��	�T�@�ɧ@�z@2�(��}Vj�!)�4ۃ���H^E �ސ��3k{*U*�6��m�pP�+���:�3����`�vm/:�)�sb�}o�sN�x�w���jIuQ��/���:��w�@>ێ��7"�F��t�&��� �Ƞ[����#d��H�:��w�@>��A.q*��Ӡm�n��*����@>̊۹�@��Z��@*:�������T��M؍Ō���e�������n@��8ڧ@�ؠ��t����flP��q�$���uN.����@�z@2�(ױO%T]/-���NH��t��y�@>�E ��i�>ǵZ�i�"��t݊��P���Vl� ���nD㔝UF��b�}w0�[�y�@8��O�HK�.�E��ۮfZS2�̶�`  �&�K�eh�v�`j�Yɖ��n��	.�IJ-n,:M�	*l=�D��5��]R7��qIn����
�ث�:;n5���b�ȗ��Y�Q��9�5��M�#�t�!' D��>�����V�:�n��Z���cu<��XK�!��ӊ��,i:�	��zd�n��������~���.��^ln�$��r#�v�7�y�*���v��I��u���X��}oH�E �ȠXf!�6H�$�à}oI�qq/ɳ}���@>����Q�6Q�)�%J�HHt���e�P�玁�� �gS��ƤrD�].W��P̚t����s��Ǿ������$���m��/2~:��^dP�� Y��d�����n�y5z�c�jW�K��e�u�c,x��$�o뻗�ސ��rENB����E �y��̞:��^r4�E�3�f��W�U��>�P�'ݐ��T}�oj:r�r����@�z(�s��?̊��t��"�F��]s�Vn��@�~ ��J��� �i���#��9@����������ߺ���u�T�uJ�J��xG �v���<���Am��j�
k2[��}�|�.�v�:C�7ފ�dP�玁�= �3���q�8�n.�{�Or��ɧ@�~ �ڣ-�nG$�S��f���/�H8������UY�@>���Z�Jj9"�!��U�<@3v(��~J�3�ˠ^��#NTQ�Q�:n� ��7��^g���� ʻ���뭽���s��{�s+ә���.+�f���Lٮ?���G���)�):��|o��}w�]���^dP��O9 �5Ck�^f�w�_��پ���@G��(��1�GA$r.�x�^dP�\���P��W@�i�T��$M�(�}�$�{�2I�<�f�WU@���R�CA�u��I=��ݖێ�+�qt͊���y�����y�@���S�$r�T霠��i��g<��=s�=v1�g��yv.����ے�n�m��~�.�x�^d^I$�Ay�R��!)�4�N.�x�O..U���@=y�]���/_��iʊ5*:g@�ؠ^E��W������,��lr�r����C��8�7�Tsw��^??s��3�~��S�NH*�P���ޮ�x�}w�ؠ����Ƅ�L�P�H�X`��H�@$H�F�����ώ� Ha&0JjB@ͱ��V�PpA�}yD,P)�XH��H@�
���@�m�����	M!�&�)�0�Ћ �_� Hj�0��%�MC��	��CkjDdFT�U�!4k@=�Ԋ#�	�ޑ5�>���  � �	��m�h�ŽN	 m               �v���2�Cl�����S=v�fV5������.v4X�.
ڸ�{e�˫!naGtZ�Y�V����Z�#�hwY�ţ�b.��v��SgCJ�v�i�Yb�vV ���x�-ڕ�#3�T6�̶���U̓;cI<��c&6�t�u�����!/<���-;S���l��^�͜�&�Q�cl<�#��q밊u�Gu���<�)��z�^�Wu�q�ݹ"���)���ػq�:+8��+uW��%а���
�ZiYU�ۭhܓ4�@vnE�չ=�٠����u;Ȳu���,ƫKjh�{s�zX�A�qfM��xm c"�Z�l�#���UQt,=��p��'YM{Jһ8"\av9�ծy��q�K�0�.Om{k97d]��f�+IV���[��Rl���'9�d5+�lm^'�9C���.�����*SbW)h�������n��V{\�+�WZ:۫��ed�l�3lfW��9@�K#R�l�
$�C���*�UG:
�U��R8:� @B9��h�tʴCd��;k-É&�R��z�$5�l��/X�k��%����i�V��mU*ʴ�UUU�g��8x�M��K������U��,��Ss�Rݻ\� ��ׂz��4ȼ�f7R���u��RKi3h�U�VBd�I�b��ڇ�}�ݮ�Ƚ
t.��u��_���#�� ���U�H`f��l*����5;r���:�đI�Y^'q�kO�M�����@N��T1C� 4��"�耉��~}�om��h  ��7,2�Mn�;;I	fi�f�2�J�hӸ��3WUuH�G;%ֆ��,粗;%�b}�m�.6r1��lv�s�n���t�5��9�v��ɣ0��sڝ\V��GNlK�m�<��k &��q;= ��bev�V�إc�j�Η�:ȇ�aP��Օ�[��'B6yD���<�7=�;Av�tE�kt��c������='P�qJU*I�g������/.�{wz���^���m��"�}yo3��^= j�ʪ�ʄq��]�b�e�utǤ븠�q�IPN�uN.����|�k� ��(W��}K�t��Ԓqt����P�b�m�ut�X��]���O�?m�dy��gT�1�8l��������O�vt��r��J��`o��Ƞ�3������p�;r�q�UQ���a�<I�H��X>+����i�7��E?U� �N���������@�z@/2(ױ@6��C��q:U$n�� �Ƞ^��^g|to��MS�)T�Aàf�P���W@��Ӡ^= _U]d�d�fƇ�戼&`NG��N^�N�wf:9���$&��*Jr�n.�y�@>��tǧ�.�f�P��q�$�'R:�@���^= ��ؠ��0��ԉĎ�y�(�͠���<X���R�k6(}s��=+[�H�"�3�f�P�"�}w4��Hl�2ʑƝUF��� ��3�|k� �Ƞ�
�E)@�LMЪ6���I��] 8���Hn�\v燷%c�qL���ؼɧ@�z@/2/%��E �i��%D�t�H�:��<�Q��@/=�㿹ʠ��uꦛ��H����E ��(j����������f<+8��NTM���f��^dӠ^?�g�&I��6QD_�[���I>�^��&⎓�S��^d�tǤ�"�}{�I,�b�(��7+��m����Wn=tr���m��į���>��Zsԑ7!`o��y�@>��@>��t�����2E*:g@�ا���$�a�� ������ 햱��J�ƝUF��� ��a�˜K�Y��7b�}�X:��ATj��@���^= �%���W��z��%4�t�H�:�� �Ƞ^� ��i�"�sW�쑵�`6ےI$ ��B��]z�cq��@Y�1�����k��y^�3�Q mc�8n�R��s �k��O,�7Z��.�*����iɲG#�v�-6q�bh8�P�S6IK��<c;q���eE�+1K�r�A�:*�cƜ��j�m��Wr�A�����fG��I9�8��?����{�����]i��r�����v�.��y�����<��@��Վӫ~@�z(ב@>��?q%�.$����?�Է�M�Jr�n.�y�)���r��ɧ@�~ �Կ.qqs��_��Ru ��GT���O�@�zB�*�`}{��[e14�T���K�U�� ��_�Ay�(�O�@�=��IQH�GL����8��ޮ�y��@�~ wXW`�j�&U�l��h݀u<[.����v����OI�s`Jg�}����wX>��tǧ�s����%��� ��zJ�U���/2~;���q%Ĥ3_�u� ���K���i�S�i�)T��t��x��}~���Ӡ���SN)
Dd�C�qV�x�^lP�玁x�@3���*'!�/6(�q,����@/����>ۮ�;<��>��|���qv�m(���5vz��H�Iԃ�@�ɧ@�z@/\]���P�yn��'�D܇@�~'�%Tf�!�r���w��<w��s�I�<���F���J���=�� ^E��y
s�(�L���o�v�X�N�H�N���U���M:����f� �5��pU���/2x���g����}~�~X��+kp�ֳQ�����8�S��;�N$����<Q5#U�RF��/�Ǆ�ؼ�Ay��@=�~eSU�"2C�f�S�IU��'��x�O�UF�ڭN�	ʎG@��P�����^dP��9T:�� 8��f���%���O6�'�@`?U
�
� n9�}KU�	�Qț��Y� ��Y���3=��f7�R���\��p��1�QB�]pk["n�;��ĥ��ں��1�U�@�ؠy���9ľ���T�1oe7*GuQ��3=�y��2�jw�O��_����7��y��pc�P���~��Y� �Ƞ�I遲PK��ZKO�*�UǾ�n� ��P?s�J�3�ˠ�?M8�)I+�f�Pq~�K�[��|n���Y���\K���]f�T�4���  ko]Ⱦk�g*�r�V�3qQ.&M��2�n�į�ȥk6W�NT�Y���!LJ��q6�����;=��Qf��5;Dw)Q�pA�pM��y��>��M���96��Kj`zM��U�vy�����c2v�,�lqnL�Ph��[�k2Mk'������&I."��g{9�p;v1ͥ8�=�V�H��B�6����L��,��@>�ή����˜I.�f�P��d�m�p���/3�]��D�mI�/�
�Ϭ|���G"m��6�� �Ƞ�ĳ?ut��W@�{Hڄ����@�ؠ�I�tѤ�
W2}h��X��1ZN4�5�3=���Y� �Ƞ�
�g"���(N��"F��c�a�i�<Cnȵ1��#�Iqr����t�������ef��"�]�P֯)�35���{}��)�I�� �A�)���B����A�k��=���ӿ�P~�?M8�*����7ފw�C��UW�?k}Pőb��&:d�qt�E ��a�2�j���$���(c��TH�H.�y���?$�8�﫠f�P�E ,��Y*8�)�����(%Ɓ����V�B�C,x��5C��M��T��Qț��=^�P̊w�(�sN��0�#pNFQt݊{�UFf� ���eg��-c�5RJm:��t͊��æ'����25! F|Mro�z*�a ���q=H����U�m��B$%ed���p�vT�OC04���5��l�h�a&Ča��ꮐ6� ڦɽ�"~3���{��]/��D8 ��/�UB*���@@��U�e���.4'�_2�S�:NECk����{�}���~��E �����E#�(�I�@�ͨ�.~���/��ފ���t��:��bv�v��EݑP�ӻ�onot��=l��n��Z�D�N��)%t݊y�@>��{���k=P���U8�i�����~�/2i�6�� �ȧ�.Uo?5PtEU �.����@ʽ��E �Ƞ���IQ�E������y�\�"O|�D� P@\ ��{~��A�85R��f�P̊��Ӡe^���u��=P8T���-g �63ӧֵ֎uZxZ4�Lأ]���_Y�a��Ձ�ߢ�}w0�W������u)�9:k�^dӾ��6�� �ؠ�~k18�(�I�@ʽ��E$�8����'���ص4Ӏ��QI+��q*�{���@>��:��%�V��P�"��q��S���3��8�W��>k=P̜�}���;�~��wط�<�m ���a*P���+k�W��Q�6K��md2��n:�>����9Ŗ��1ۜ2�r��]���4JrZ�H�.�h��aa.�ו4�I��=����[���ř��x.�pg��Ӯ��b�[]��x�<j�sŲh��j����欏L��sv,6�W�<��ݩ���ܑp����B9��Km���E[�GG�..s�N����(*�Q|����2�jy�@/r(i}��JqH�H���W� �ȿ.v�=�@/2x9��%ēf����jN85R��{������W���7�G)�uU�~I.s��ߺ��4�W������u)�ۅJk�^dӠy$��k�W@�ؠ��^uFભ�ȡ�-�]˸��С����Ymn�!@;sH�2"q�Q����{P̊{�~�]����{=�M8
)U��lA>�T���P+���&tP���@32*���t�����빇Oq.s��k=P݊�����('R����{P̊�\���@>��j��RrG���~�������ߺ��X��(ǜۙ���XG|�ZVM��;8l#npq3���Fv�����Du��E �Ƞ]������Y�}�-}��9N����@�lP��e^��"���UFy��Nn)������W�����@/r(�X�U8�(�I���s��=P݊~Ƞ����{=<����QI+�f�P̊��Ӡe^���߷���z�n��hKIo�'c�	�jx@wF&(�J~\��ӭӜn�d�qX��(�s���y�@>��4A����Qt̚w�UF�z����O�qUJ�#T�"p�"nC�mg�w�C�J�?lP�'��x���ӎ��G]3b�^dP��:���$���X	��`@!@p�/z�'�0=W�S�):�����%�gt���@.�(�q+��Ҷ*��2�CUEH�fG���e�֦y��㵃�:2vG-@ۆ���o��g���{P���s�>a��o��aj��àe_�]�P܊۹�qs����k�I�Tۨ�~�v��}?�^�2�ۜ��d�H�n� ��àe^�%Y�� �~���*T�E5�>̞:�m@/2$��$���E��i�L�h���  K�7l�=d�n�F�nh���8ajV��1"pX%�LpI�i�r�ڑ��[���[n������^<�rn�M�m��Yv��#<֯5;��ٹ.�����Ka��E��:-$���%�ɢ,�>���pcܘ���B�@�^�R��]di>���[���]��:ݖ<	���of��\�9��K��ܱ�Jk̿���V��Q\�T�`m{� �Ƞ_��v�i�>��БF�tT�:���Ƞ]�:�mO.Ua�v6��JN��]7�@>��t��ʬ��P݊w鐩*GM�Tk����Ǿ�ߎ���� �Ƞ_��Y��D��*H�:�m@/2(ױ@>��t��V�"�rm�Y�Elv�-[n��i��`2Sۚ����{���-NFQ��}�^E ��<t�ڀ]�s��n���^lS�qO.%ޙ��N����ב@>��2T*�Ȋk�}y4�Y��\��ؠ���^�����U8wj�..s�I���n�(��(n��}m�"�85R��flP�K��Ĺ��|��g�]g�~��Ҿ����j�8���h��dl�iΣ��#�`�t��=WI�:���UF� ��v�a�.�� �Ƞ{2:p�ASp
��}�4�丒UFV��� �����T�TM�zɹ'��ܒ{�d�O����DП�G�����5�k$�}�}7$��4CS��E$����@����6��0���n���������+���y��I�4֖�^��i%�~{�ߞ���ۮȹ��=�<ٷx��Cu�ք��O#*�r6T���#�����}��]ۖ�-�>�UU@m���"O�w����N:�QN+=S*�̊w�@.�i��.*��b<�E�U(����y?$��8��2~:������m�u �UF�g��]�àef�Bu"`@"�#��d���6:p�ASp�5�32x�Y� �Ƞ{�b���%*r������ۻ/&'����/�L%<��,����luv#E�$Ko�2�j��@.�/%�s�����{}<����"�W@�ؠy��+6����3riM���S��qt�E ���@��T3"�]���NF�t�
k��$�w{�mo���@�˜\{��P����N:�"�:V~-|���D�{�:I� �P��<"V�
4�꾞��Q^$!��X��4R���!H��� �t�<"4��IH��R�^+� "E�i �ň�^({<6(b�P*(xn�6��� ��2t�}��   ��$H�bAËz� �               'Z��"ҫ]:�e�����
:���q8=��l�u\Y�-�5t!�V����Pb�j�V&�����]��d�������큋p]�˃e�X�kKU$9�U�7B4�T�u���,*��p��V5!�jF��˒�S��7%X/�(�˚�s�b�j��2��T!�\�9��B�$ޤr�(�)���4Vx�����@����;�E^W���Jtoo$mʵYn��oA��i��l�����:2� m;M��+�iiYq`�����g�θ�L�S����
���[�[����^]U�9���W  ASQ�lq��f]�:3�u;:�:ν�:��4�rreۭ�y�ٲ�O�j�Z����vb�g��-k���sl����� ���"���M׹�,�M'����uq��ē�k&GV�8����l�c'
x0ɨ�˺�@��-�n�g�3�V�M�ӭp��bI��vn���͎�u�yN�=�1Ŭ��창�A�3m���uIW���"s=��U��%j�Y�@�)d�&�ćQ��gX��`%�)V�fl�N�ɶj5�Y���t��nٶ�J�U�Z�5��逥%�U��eZ����<��T�m����sƬY��Z�B;@ca�n8�X���� �eئ�uڜ�[2K�(��*��iT]���l��.��V̳���Jv�I'���"§�����wm��-�{�vB�A+UV�����j����.����(T �D���!�AF��b���>3�A�K��G�:�=^ )Q_��bP=�sz�fkZ�0�RM��  ����Wn+rT����xG�6��d�Ig�[^t�ڊs���ka���su��1�,��d��sԶc���H چ�`�/�sr�9J�%�v�:\�a��TŵHn�WY8]!�Z�(�V�ƕ-s��ڋm��ǭ�Ã6�=�ӵe.9&���l�Eٍ�<�����{c������:D����A��;WN`'I�7b�]�P����Ŀ%�[W�T��v��)�8�Tk�f~���0�Y� �2)�.r���68��P��Dk�fl��2�j�dP��z��EJ%Dӎ%t?qV��@>݉��E�K��?mt{��MNFQ��۱@.�(�=��Y� W�x�R�����ɳ�u����iK/pvf-�&닛=3�����M��1�N7�n�(�fut��~\K�n� ����NF��*.�w�MT*�z�r�'� �=����ԯ��JqJ��G@��T��@.��:�ב�Eq�FG]�ؠy�z�\�{�}foj:��9��]3�@?.q+�ߗ�mo��dP����Ƞ�ƣ����\'d�5�fUx�	�vLu�<�=L�9nܷn��}}}�Ѥ�nZ$��'��B����hYO~�;�\�3SF�Y5�m9ı,N�\Mı,K��f&�X�%��l��Kı<�߸m9ı,O��ύh�1�VᙗiȖ%�b{��17ı,O}��Mı�m >�AJ SA+��M��J!K��M��~}�iȖ%�bw^�q7ı,N��xZkX�3W�6��bY�05�f&�X�%����ӑ,Kľ���7İ?#Q=����bX�'{�����5K5��.ND�,K�{��ӑ,Kľ���7ı,O;ݘ��bX�'=�f&�X�%�}�}orsY�-n�Mn���q��FLUk�5t�����[���)�\�iȖ%�b_~�X��bX�'���Mı,K�����MD�,O}��ND�,K���_��0ֲj�Z�r%�bX����Mı,K��f&�X�%����iȖ%�b_~�X��bX�'<���5s.��֭�ND�,K���q,K���{�iȖ?�j&�^���Mı,K߾ى��%�bs��֭۬�Y�f�.ND�,K�{��ӑ,Kľ���7ı,O;ݘ��bX'�g"o3�&�X�%�ϲ����uf�u���Kı/�}�Mı,K��f&�X�%��~ى��%�b_<���r%8�⣊���D*�8'�q�"�<�&����7��zݝn6ŰًQղ�\�R���oqı=�혛�bX�'=��Mı,K��fӑ,Kľ���7ı,N����kX�3W�6��bX�'��f&�X�%�|���ӑ,Kľ���7ı,O;ݘ���T5SQ,N�;[%�Z]]fItm9ı,K���6��bX�%�﵉��?�Uj&�{��17ı,O;�f&�X�%���&e�s5��36��bX�%�����Kı9����Kı9��17İ?MD׾��m9ı,O{���L�k&�u��"X�%���l��Kİ�"�p��Kı/���m9ı,K�﵉��%�bi}��]k]�s,l�nfff` ��I�N;,t��[��u�ʭ�Յ����L��#�#O[���7�I&z垯c�cs)�퀗,���
�ڧ�b�u���6.gI�s��=�[��mb�n���=d������gg���%��6�n8]�+V�x�u�qs�]��bӗ[��vE�IlнL��"�������Ҽ��m�Y���u�3��$��V���7�Lf��jZ�P��{�y,K���vbn%�bX��=�m9ı,K��kq,K��ى��%�bs���W5.�k4ˆӑ,Kľ�߳iȖ%�b^���7ı,O;ݘ��bX�'�}�q?�T�K��Ο�MS���r%�bX��ߵ���%�by����Kı=���Mı,K��fӑ,K���|���I#}��⣊�*8���7ı,O|��Mı,K��fӑ,KĽ��bn%�bX��ݝ�SX�5���ND�,K���q,Kľy�siȖ%�b^���7ı,O;ݘ��bX�'�y�ِ�3ks۪���T�A�O�5�n{=���u���K���kYItq<�bX�%�~��ND�,K�﵉��%�by���7ı,N{��Mı,K�<=���Xe��j]fm9ı,K��kp��]�D�%��}�q,K�����Kı/�{�m9ı,O{��|Lֲ̄j�Z�r%�bX����Mı,K�;�q,ľy�ٴ�Kı/~�X��bX�'<��W��5��Mj�Ѵ�Kı<��17ı,O<�{v��bX�%�﵉��%�by����Kı9��kY�sR��ˆӑ,K�����iȖ%�`��}�Mı,K���q,K��϶bn%�bX�����k%�$��5!s7#�:8���<mb��e��1V�V 8�ni5��:sZɴ�Kı/~�X��bX�'=�f&�X�%��l��Kı>���m9ı,O�������C[���m9ı,O;ݘ���bX�'�wf&�X�%����iȖ%�b^���7ı,O|��.�&��kW�6��bX�'}�f&�X�%��}�fӑ,` ��#E�A�Ӱ8n%�u����Kı<�혛�bX�'�緥��!��f�p�r%�`�6'����r%�bX��}�Mı,K���q,K��l��Kı9��g�̺�.f�%�m9ı,K��kq,K�����Kı9��17ı,O����r%�bX���zK�mױ�ܶ���n�i�K����F�FE���֋���������T�Cpu���gTqQŞ��Mı,K��f&�X�%���{ͧ"X�%�}��bn%�bX��{�^j��e�5�sFӑ,K��l�� D�;���A'~�X��H���&D�~���'���Mk5.jܙYp�r%�bX����6��bX�%��kq,K�����Kı=�혛�bX�'�e��.f�Z]K���r%�g����~�&�X�%��{�q,K����17İ �#:�Ț�yɴ�Kı>��e���!����ֶ��bX�'���Mı,K�;�q,K���wٴ�Kı/~�X��bX�'����_��WWRn�y-���'��[���g�����~;��{�Z�X�5���O"X�%��l��Kı;���r%�bX�����Ț�bX�w�17ı,N�;��%ѓ%����Kı?w��m9ı,K߾�&�X�%��}ى��%�b{��17Bı,Nh���ɬ2�k2\ɴ�Kı/~�X��bX�'=�f&�X�%��l��Kı<�>��r%�bX��w~�32Zɫ�]kiȖ%�by��17ı,O|��Mı,K�3�ݧ"X� ��{����Kı<�{�^j�ֲ�5�sFӑ,K��l��Kı<�;۴�Kı/~�X��bX�';ݘ��bX�'�.��v�fZkS-l�h  �݌,3��;\7%."��g$��8#U��t�S���S���{x���h,\�-��nn�V�mӉ���2�ڹ�n�xuc#o��?m��M���=ch詞퐈�u�ù�C=���8,�"/N6�B�s+��v��zv��'��٧���]q,C7&����b��n7��c�q�΃g���عoz�ɡ㵕��tw�k����7v#��%�bX�w?~�ND�,K�﵉��%�bs�ـ!��%�b{��17ı,O~�=:\�\�����]�"X�%�{����Kı9����Kı=�혛�bX�'�gݻND�MT�K�������!����ֶ��bX�'��l��Kı=�17��D�&�j'���ӑ,KĿ~��Mı,K�{�ˣF��kW�6��bX�'}��q,K����nӑ,KĽ��bn%�bX��vbn%�bX�k�~&�%����Kı=�>��9ı,,5�����Kı<�혛�bX�'�~ى��%�bz{��k�a-֭.wd��v`�焮5��ny.ɞ悜:�\Z�tSvj�9ı,K߾�&�X�%���f&�X�%��l��Kı<�>��r%�bX��߲K�5���eֶ��bX�'�}�p�Q5�;�!׊%���&�����bX�'{�v�9ı,K߾�&�~U5���ߵy��Z˔֭�ND�,K��ى��%�by�w�iȖ%�b^��X��bX�';ݘ��bX�'=�e�Y��R�`K�ӑ,K �=�>��9ı,K߾�&�X�%���f&�X�%��l��Kı=�,��s5rYu3-̻ND�,K�﵉��%�bs�ى��%�b{��17ı,O<ϻv��bX�'~0��2f�%��ʑm.�̇K#wg9Q�l]�ݍ\��}tF>�{������f�����ӑ,K���bn%�bX��ݘ��bX�'�gݻND�,K�﵉��%�bw��lѣX�5���ND�,K���q,K����nӑ,KĽ��bn%�bX��vbn
�bX�k�~&�%����Kı=�>��9ı,K߾�&�X�C�t!��2@���Bh��A`�\�"�ϴ��Dp���B�����[l<4WMmia@��>
A��5 �i$B+H�8�}��	|y�|]oH:�H�Z�[��1��b����F�b�075aC� @�.�N����T(CJ{<���"��϶�_~���>��*>2 +�&lC�؜��}ى��%�b}��17�Q�G�^�������|qQ�BX��}�Mı,K���Mı,K�>ى��%�'�gݻND�,K�ÿjNj�d��.���Kı<�혛�bX�'�wf&�X�%��o�iȖ%�b^���7ı,O���Ǯ
P6�N��R�@�	�W)ź��v�\=��`�ΒmJ�] JIe��V�����q���>�혛�bX�'�w}�ND�,K������G�5ı<�혛�bX�'��ٯ���jXXm9ı,O}���ӑ,KĽ��bn%�bX��vbn%�bX����Mı,K�-U#*�IQü_TqQ�Go��Mı,K���Mı,K�>ى��%�by����r%�bX�w鿦��a�����ӑ,K?D�����bX�'}�f&�X�%�矷ٴ�K��L�C[��~��Mı,K�3�ѣX�.��ND�,K��ى��%�by�wٴ�Kı/~�X��bX�';ݘ��bX�=������m���-��p��A۸���]�� �ӊ����.�����{��oq��'�g~�ND�,K�﵉��%�bs����Kı=�혛�bX�+�(��#q�#��/�*8�⣊�﵉��%�bs����Kı=�혛�bX�'�g��ND�,K�߾$桚�j�2涜�bX�'�wf&�X�%��ى��%�by�{۴�Kı/~�X��bX�'=���\���h���a��Kı;��17ı,O{���9ı,K߾�&�X�%[y�8�qQ�GW����4�q#Xm9ı,N����9ı,?1�߿k�,K������Kı=���Mı,K�3c��&4��Ģ!rpO:�IRUE(�`  ��\����Vӫ��v�ŗam�B�a��V��n�vX�6l�[��6ctvs:�ֆ0�:��v��j�.�i{Y��q��t��-���t��^�8����vk����z�+Pl��'���N��$U.�XF�uv�^M�[��]�^����̓�#���������/���0��[rn;���gvx���N����R8�3�zᐳ�Uu�iؖ%�b_�}�Mı,K�{�q,K����17ı,Ou���ӑ,K���M�5us	fffk[ND�,K�{�q,K��ى��%�b{���bX�%����ND�,K�s�Y�F��]\��ND�,Kϻ�q,K��]�u��K �,K���6��bX�'���Mı,K�wޙd�efjf��ND�,K��ﵴ�Kı/�w��r%�bX�w�17ı,N���Mı,K���8:��Ȝ���㊎*8����fӑ,K���f&�X�%��=ى��%�b{���lyı,O{����t]�����u�> �ZWWNt��,/eՠ-�{i�,��������oq��w�17ı,O|�f&�X�%���u��yQ,K�}�5��Kı�w�h�K0e��ChxгB�4#�17U
�P�� M��K�w}�ӑ,K��^�����bX�'���Mı,K��I�5.�&��r%�bX���}��"X�%������r%�� �5Q?}��Mı,K��f&�X�%��^�{%�jܚ�Yr�f���bX%��_w�m9ı,O�ݘ��bX�'�{�q,K�c����TqQ�����H�"	S35��Kı>�vbn%�bX����Mı,K�}��iȖ%�b}����/�*8�⣊�-��(GHm�q�#{��'�l�;���n���韽�����<��	���iȖ%�bw����Kı=�{�m9ı,O��~���Ț�bX���f&�X�%������fe.]\�k�"X�%��w���r�H�&�X������r%�bX��}�plK���vbn'�5Q,O5'{?���[��Z��ӑ,K����~�ӑ,K������K�_�T*!��"n&���Mı,K�}���r%�bX����C��kY�rL�kiȖ%�b}�vbn%�bX��ݘ��bX�'����iȖ%�b}���m9ı,N���j̚��h���a��Kı/��7ı,_u�{��"X�%���ߵ��Kı>��17ı,O�k���m��=u�g�˟���
b���+�V�8z;K7�5�j̸�����~w���{���?�ߵ��Kı>�{����bX�'�wf&�X�%�y���Kı>׳��u���k.��5��Kı>�{����`ؖ'�wf&�X�%�y���Kı=׿w[ND�,Kﾛ�j���$˙���"X�%���ى��%�b^{�7ı,Ou���ӑ,K��]���r%�bX�}���jM`L53&��r%�g�Tbj&���bn%�bX��{����bX�'�w�kiȖ%���A�1K	 �0] �"&�D�_l��Kı;��ٖ]a��̓0�r%�bX��{����bX�'���kiȖ%�b}��17ı,Ny��Mı,K�<��ẉ��kv瞷���9y�?�?}Zۍ]!�Wt�hH����RD�*�"m���TqQ�G�����bX�'�}�q,K���vbn%�bX����v��bX�'�C�j�3Z�[�\�m9ı,O��f&�X�%�����Kı=���6��bX�'��ﵴ�Kı;�o�ՙ5��ѭj�4m9ı,O}��Mı,K�=�fӑ,��&�~�~�ӑ,K���혛�bX�'}����ɩu�5�ӑ,K�����Kı>׿}��"X�%��~ى��%�����ቸ�%�b~�g~��5,.˩�d�r%�bX����kiȖ%�b}߶bn%�bX�y��Mı,K�=��iȖ%�b{��_߳�~��Jk�l  ������_V7KͲ�6��v�\�a��#�m�Ζ]�2 ���u|��f��i�=�`��<W���#����ɵӥ�Ew$��2a�����PG"��s��TP�H�۪ۑ"m3����'��t��\�N�A`��A$V���v�u��{-�G{�}�]����w��q�{Oh2v7��ݛ�q�[8wm��3��"Wn.5sY��v%�bX�����Mı,K�=ى��%�b{��&ӑ,K��^�����bX�'���.���fMa��Kı=��17�:���'}���ND�,K�������bX�'��f&�X�%��3�ٖ]a��љ�iȖ%�bw���iȖ%�b_>���r%�bX�w혛�bX�'�wf&�X�%��^��fh��-�a5��ND�,K���fӑ,K���l��Kı<�17İ4�D�����r%�bX����sP�k5n�fӑ,K���l��Kı<�17ı,O|�~�ND�,K���fӑ,K�/{z�"�"���8≺
mD���NgNIP-:�u�g�3L�R�=������b{��17ı,O|�{v��bX�%��͏"X�%��~ى��%�e�g&a�p�F�!�<hY�f�����r	����MD�<�ﹴ�Kı>�혛�bX�'�wf&�X�%�����.�P�ᬺ�Yv��bX�'�}�6��bX�'��f&�X�%��ى��%�b{��m9ı,O����WW22]k6��bX�'��f&�X�%��ى��%�b{��m9İ75����ND�,K߾޾�F��˫���iȖ%�bw߶bn%�bX����6��bX�'���m9ı,O���Mı,K��{{����:�=��ӄ8��]���R�&[�GY��L.��n3Xm9ı,N���6��bX�'���m9ı,O�����$O|� �	��{�W$�Y�5�6$�H�����O�X�'{ݘ��bX�'�wf&�X�%��{�NAlK���w�C��kY�r���r%�bX��vbn%�bX�yݘ��c��T((T�D@�P�U����E���O���6��bX�%���6��bX�'�w�^j��e����ND�,K�~ى��%�bw���"X�%��k�߿f�Ȗ%��u�ቸ�%�bw�;5��.MK��6��bX�'���"X�%�|��fӑ,K��ى��%�b{�vbn%�bX�����Kl'���Ӯ9{Y�v��	V�9&��M�m�H����Bˆ��kY6��bX�%��ͧ"X�%��~ى��%�by�vbn%�bX�����ND�,K�7����!��f\�ͧ"X�%��~ى�~ ��j%��~ى��%�bw����r%�bX����6��bX�'�wz�].�fMa��Kı;��17ı,O|�}�ND�,K�߾ͧ"X�%��~ى��%�by�ӦXe�Y�m9İ�;�w��r%�bX�����r%�bX�w혛�bX��XC�L�O��17ı,OMt��W$�Y��ɴ�Kı/{���r%�bX�w혛�bX�P��T4гB�m��I%�w��%V6;���p^����[�`��A�T�ӯ,҇7�㪊�I�7v(]� ������\�=����=��v7	%F�:q����@.�a����7v(��x�Pe9�T]3&� �ݝ<��W����fb)�P�')�p�{vt݊�q@.�i�71M:�
��$�wb�e�P�U���@7����ēE#�j���U},!'�����J�u�]x�@}P�JR����2#*�
o�fsI����$   � (�� 
@D8�Bc9}L7��#UX(�&�)&(� N�9���I    ��$H�b@z�  -�              s\�Y��:��`�٭���q/f���ـ�5��n������n�Ĺ,2D����lK�T��*��'jM�����"V�C�r���8K�U8*�[�)rB�9�v�(�mW{lp�ҋT�v	��pML�S*r�)��n�r*�&�}��JVI���-Je��5\=��:9y�a��SM�,{�@nҺ�#;������1��ѵ�"�)#t�
} mɹVe�V��Bt-��7[ulk[���'
�����jI���zj�,K�
y�7FA�����Y�ڸ퇚�3:l���+v-�gs`�Vj���ܫP����@]���q�h��;���<<ٳ�ԵT�K�
ې�
�S$]�+ct�UUIr�!�I�2b�|7+m�^�L�h�0,���=g�ͷQi��F�]��v:���O��Ghʂ���R�Fyش���'�6qm�5kW/@m��ɨ�V�����mc���i���g��n$�7\��]�0��4�T)(r�T[�yj����c gC��e[���%j�.�m�Z۳+W�v�WWJ��fY^��U��l�f������Ca�q�UF����o+UUUʵ{ ���R��1m@UP4ڒ�"N�WI72���r�c7���V.y@������C:i8��$�vˤ."=DL��6��L�S%ts��v\o�����Z;UUm�����ӫn�h�r�Nq]�Q�.�$jy-�M��s�g��-UAvii��2�d&���7&�';�wf�ɺ�fN����߼�j��%��)":)��� `lQ�A	꠹�v�T���3��o2ҙ0,�h  z��n5[4��,.x'���7W`ݢ��o�������kP�VkQ��9u�$���v�oc�Ul�F@�q3�<m��lډ�1���vb�
�OZΛv糵��e�c��=��糹)ŀ6�V�9CiU0�nx�\��hm�:�<�z�lHqv6Vn������{ޘ?�����m��:B�whe8�T�
9�8]/�Vl�4~;�1���k�(qh��@.�a���:�� ������R�&�E�32i����7v(]�?�~�l�Z��P*���à�����?s�s���Ƞ�<tZ��ID�I�7v(]� ���@3wg@���G�Tiӧ���fgt�}�Oq}A�z(�Տݍ;p�������3�R��ќ-���<8�ݘܻ�ҕQRTm�NrUE�32x�nl���< Vf"�e
�r���}����U�$��q$�g���]� w<w��UG��:�
2�)�:���� ���nl�^��i��Q��@�ސ��t�͝wb�_�]a(n(�1�C�fdӠnl���< +e��AU�\9�9q��"�m�z^��a�֦�qy��ͩ�낢)ànl��H~x{����?���ݔ�����I:c�~�\�>�����~��2�{QƤ�t�N��~~ ��t���s�y�N���@>��Tm�Np:ٓ�@.�g@�z@;����B����à{��~�K�[��@�z@;w<}��9����umV��%�X�'`���A4#C�ݍ\���9VY/m�����O������ ��Ӡ{��}{�����
��rm�=ė��ݞ:���tǤ�Yk 7u$���@�2i����3��� �W�p$�J*�")ɹ?
"��~�7$�u��'�׳$�	"��
AD�s��|7mn�Rrpn����2ސ�� ��ut/vt�M��mS"��\I$�K�e#,�'$v�9�1Ş* ����Z��6ސ�gW@2�g@�z@>�Y�7EAӉ���︒��zt���< ��1�T�#��{��]�!��ʭ���n�tf�A�D(�R7$�oH|��ws:���:^��mөª(��@�z@:�Ѥ��E���hUm �A���}m�om��[l  n��\WQ0�;�խ�G��1s�W-".6�:�S�も��ځշ�����|ܽ=�%�Y��+r� n�@�v;r'D]�<���c��v��!><˱�U[Vs��d��"Om���;h�����fF��
:�X]ێ�r�D��rc�j�pѰ�lSv��{����ｻ��n��M�{p;�؞��`=X.5����t竕����8��S�'�������L���>�������*��{BJt���(�] ���@�ސ�� ��utś�L���&ܝ�z@;�v�{��}��c�G*Rtܨt�� �ٝ] �ݝq%W�����#
����@���] �ݝ�z@;��� �9 T�UQ<���S�gvϩ�ƒ�!Րc��x���gq�"�w�{��}�Hq� �۝]wI�l�
!ԍ�:�����9�%TV< �s��{��^n��T�NQD�:��w�ή�����}�HVZx�8��%I*��>�ޮ�����}�Hm� �W�p$�J*�"���Y���g���< ����3�W`�GPR�^KgZ��!�Vi�Xmi�4t�iz�Y,��R�j���>Ǥ��w�ί%��7Ϡ^o��"�T��P�[�߳:��澁�= n�!T�Np:I�I�I2����ª���2����B�8s��\�q�@>�� �e�P7�ER�$]ՙ��}�Hm� �۝]wM���hP�>��= �d�nut��} �]f��@�EGN����x�v�=�v����ۉ���G=3��Ѕ�N��t�� �ٝ]j�_���~ Y��ۊJ�	T:����W����}���IC"��*�.���f�|�}w��(���F�df�#�J���c�ߝ�����\�=@�	H0�
J�@�޷!w�뮠ܩI�r��>���fut��}�z@<�8�}�UJ��"��rg6�u�񗙐�np��k�4�-\ٮ+M��������澁�= �� �ˬ�n7\��BH��澁�= �� �۝]wM���h�L�9@����w�ή��y��^n��S��TdMà}o~���W��\�^���jm�!R��t����6�5��� ���W�K���d���$�l  x���]6qJ�(<���o.�X���q۲�<�H��7Od�6.�C��(F�v��*[:���i������3��Q���@�t���Ȼ��W��3���ܗ!Ee�����]�S�j%-���ۮ۬�S�{S��U��5��3�3E˗Y�z@AM�#�9�j�Q<�ƷAv��x�
�9�����c�3�H�[��'N�8zE*"��*�,��y��� ���~������|�N"QN>��= �� �۝]j�_@��]u��)R��2�(~���W����f1Tt9N�䪋�}{�]j�_@��?qU�u@=[���뒈BH���_@������s��u{�}�{��n�m��Ŋ�c�����voZ
���{\g���Pq:u�29$vy�{�P��e}��Z�:u^�2&��.��:�(�A "iD� �����.�u���=Tmn3U7N����/=�{��}�H�\P�|�T���Ȉ��W����}�� �۝]q����7Q9Dq��琢O��"N�=I��f�Kw"B{����q;g�9謧=���F�g3�5�����q�II�r��.�(~���W����f:�N:���*.����t��}�z@>����Y@�n�EI@����>Ǥ3 ���w��@����g���`6��YM���f�z��H��#5D"���!��wӡ$���y�)R`0"�BB@���E(k#�Ya���0bP��vF2@5�֙�K=Қ]4}��I�%�DѰ��#B,R`�Q� �*�o��#�\�����p��B�tʬJ$�lHw��n�"��m�m�,N��h0��px$�k�ClR,BA @"B\`�d3K�b�0�@%��H��� '� �!�@!�S~�-�E����Ch
i��{Dz �/��@2�:������g"drH���W���"�w�gW@�f�����C�Ȉ�Mà^dP����6�u��� ;�WY �G	+�(�*`������=��i]�Gkɮvt��in�I����z�y�:��^\P�|�	PS������>Ǥ��w�ή�s�%T{�v��N���9:�� ����������>����II�b�t��Aw���I�"�~���$TH@�#$P�X	!d��P���	DRA0X�H�$5(E�`�@ @"�In"{�K��~ ��q��9
��}~ޮ�^n΁�= ���ʥP<��.�]Y�6��nƀ	V�9&��.��]�YaѴ�u�(BH�y�:��^\P��W@6�z�:��b���}oI�$��܊��z��{_|��J��l<�'S����@�lP��W@��oW�Zs���!��9
������}Բ�������C��t
�8P�Ă�@w��=�y�����0��?���V.��VUݠ  n��/����r��y�$<<�L��9�l�O�����;T�[���!�䓲��+�.6aN9��n�8���۶F��w71��:���B����۷bk�Ŷ�nW�J.��[C�/�Y��&śۥ���U�X(�t���ңM�I#�k2��NĜ1�3S3	�@�\�%�Hc,��eu����w�%�I�]�۱\��4�X�ז�PC�K�#x���k�����;�Mne��W�+y�Ѯ����rh�\5��yk1,9��Z=@w��=�y�����
�%tPE+H�G��?46s@l�r�����KG��?46s@w��&��~�~��ٝۛ��:�Z9��AY�(����v�����RQQ:�����9{{r�%d�=�o>��A�J�h�q�%�� :
�P�7����<߾��p��p�w�x����=�{[_��� >�Ͼ�W�vq��Z;����ǌ׼���\Xm�+y�Ѯ�kx�{�N��ӞK�s+J�)@�P�E��pEZ��GnD�VxI��F��$v0S+<�t�?�������;����K��Ŋ蠊X�׼���p׵�6_;����/-a�k��k���	��� @k��k_9�7�]�T��(f#]����{�M놷�`� ��"�Y�=@|;���^W�}�ȭ}E�� ���MJn�m��ݛ<@Uoi�v7f��FRK����x�Y���.w{��&�u�^�hl怌9�1^U�Z����{������sG���VXŊ�^b�j9�� ����p״��³
+2�&�g;�p=��{��^�@�*��B��@"�C��ǀ��tPE+H��놟6��h������H�����SX��ɧ���\N���\t�>�#<܉;����9�Ɵ6��� ���7����T��(f#QȆ�h����kpDNb.���h������G"þ+8���A^ 7��u�O�Cg4�8���8�XRZ=�>m����
*��J�fwVUݤ�I�D��eRS)�&�-V�;f�p�.Fpݚ����[ry���ٔp6�\����ys���R��V�ԪE؝ga�km�r�u֨���yܰ\h�v2�7�'���v�4mDV��y��b�O)��p�Ӎ�]
��+q�s�H�{C�T�d5��$۳�Ϋ�v0Ո����pI99̆Y5�&�!���M�7Uj����M���y�tV�k�cQ����V�}��|���G��i��fVe�N-� 74{�|�/�<+��)Z@>nh�\5�������1a�b��pכho�@w74H�]��H�b5�D7͠;��<�~Is��WY�"��T�7B#����=�p�����i��{st4V��8�����?_��盚<���D8�R����$
�<�߷�C���+RЁ �0"��e �"T��ƷdC}�@0��3���B��G��O�C}�sG��K(�����h�r!�m �����i=���(�8��Z=� 74>�i�hzp��%ĭ�ͻs�;��K���+/����5��3�ř�ʺ)�H���|�Ѡ=$1e���VX���>|��h�M<0^�!�a�j8��mU��EP��*�*���4>�k{�31�%i+���D���>mà(����$
����>m����q�%����:%��8�Vi�)�z�Ȳܣ�B%n���X��-aX�>�i�hoF�|���(��c/�j9�m �����^�{���BXm8�yȀ|����͡�|q�8����E%_����'�#��>m(P�@ :����M��VY�C놟6��h���u�H#d�h0���݀9�����Mq�gѦ;����sf(E����0�8�I�����xG��31�1$�֏?�����Dw�͡��w����wx�)#O��\4�����CiW�
���y�4�����&�u̖QG+y�Ѩ�Bh�W�#�zic�x��2BHs�	����C������A޽���!��?|(c�G}�a{�H �y"
�*����; ���"� ��PQ,DQ�@�X@ZR����P�_ک�`
�#� ^��?�������r���լ�C���T����fKX�CR�R؈�"?4�K��:C�w��">�.
�����	CO��w}*v��M�n:�ψ��*�^���qY)�Wr�~��kH��{����[c�s{�hr�`~][u���E�AD	 J��"�� ���� ���,",AF�T��@ �� ��A�"��"�E�"� �"�B�b���"�  ��b��  ���,( ���",�"�����4*�"�(�",�� "",�* �
�"�����b
�V�H
A�^{��&�e/
ֽVp������
�#���M��������M�a��Cבo��3�?����*������~i�é�<��(�0C���"����<��{���7��n�EGWxo�w�O_Ǖ��Q�1H=b���I�PD~g�����(��@衛��2.Ay���a@UF�leʔ�&��"4�4r	I�5 i��NC��R��,���q��Mj��#��:���o���oy{R���iI�g7�)�q���<J*("=��}��PDv��}���<.~;5N�b�-
���P�#Iӽ��P��Q����AۭNi�9�d���9sfm��2�i`���dm �G�`v<J�Sf뀨"<���*q�G^cDۆP��BwQ�K���w$S�		�D	0