BZh91AY&SY������߀`x����0����a?         b*HB�US`�(����T��"��IPJ��!$�)U(D�
CJ���@"�*AH������	 Q� AB��BU@
��H�(�$� ��  �P	.     �3��    ( v 4��1!�@� }� D7�-p :��wπ P��t�
���7b����)�Ψ�8��mN&�V� >�^<(ng@'g6��N'G>�t{� BE  � 3�G����d�lv{���<�=����OxK��c�ngG��o�@9Ҭ���6�縯  ��c�>�F6��m�Zy�^-+�q2�8 zy��9o'��n�ݼ۔�y��-x >}@P 
�
 ��mޱחO69��3��m��F�����;�疞����6yOx y<��-�r��������,�y�v�W ��[��-���{�8{���U3�v��뾚��8����� ��E (
%"�� ��Yڹk�<�ƻn{.�����w���|os�Ξ��� ��E��`�b� �糗��p t�5z���=ܯwx�S� 8{��a�Ǽ�R����  ��
�P���8� |K��^js�}yx�{7>��
S����{�C��>����	�X zp5��`�7  ��Ÿ�u7 
`u�ϑ���f��w��Ox Q��w<����s���G�           ��i�6*R�L�� �2&�0��	))�11 �  �=U*�# 0   	���U*LB��      ���1RT�      )�QR
zS���h52z�F�ɦ�����'�������O����퇷�����u��*�^��@PU� ���UU��(��*���"
��r�Du���:�Q]���4	�!r���H����:��	�!?�����G����%�0���=�9�_%�b���7��$9 rP{�y
rS��$HrD�P�s�
���� �)� �����D~J+�AH��Uy�P9rH��D9*��@!܂���F��P;�W�"���@�%P9*!=� �J��Dy">ʫ�y �!䢾H��U�*�䪇%B��y �P���9�%䢡�1�r^I�NHr���OeNH���S����� �W�S��!�C�^H��9jC��%9��)�@�%C%y�' ^\���#���<�aL�NBr@��Hr��P��@���!B<�y+�9�9�C�$9���K�9�<�9RjGR�B�����'$9#�B��^K�ےr�y)���0C�]�$NG �$y�!�NA��^k9���C����%�G�%�' y)�^H/.@� =�!�!쇰Ȟ��'�S�H<�9�C�r�<�9">�r2@��S�!NBrC�^@'!Hҏ!B�����^H��NB�9(rD��9!���$9 �yrE��P䜐�%C�<�9&�Ԯ�9!�NBr;�rC�'.����J�9/$9=�r��w���N@rG���@�<��{�$7��9��!y/$众�9%y ��:�9$䔏$��S���b���G�<��S� ��9!� 9ry	�C����G�!9�H����!�@��$9!���J���H� NHr���!��B!y$9�d��9#��	��9(�J���r�9$NJr�<�9 r9�9#\������T�����܇!�rJ#��'�''���
^JrNB��9r'$9�yu#�NH��������{�P�䜔�/ A��H�B�:�9'$9$9 <�9�@�yr�$�!|�}� �w��������9%y%<�䜕�' y�y<�y�@�=KԨu'RP<��n �����<��'�������v����!�����ٴ��%�8��Ӡ5�A�-h���]&���M�Bх��Ѥ��Z]4j���h�h����%�t��cZtf��fP��:WC�J3Z GB�'��ȧ��}+5�/҂ ����3ӫwC�"ϱ�W�X��T�ZS�cASS8p��jo�f,�I�����J�1zH'�v��g�����xu��O#s���������{�F̌[.�ï:�:;è�{�h�:',[�h#]4���elv෭kGM�@��I8yh�P`�6�th���Ը�
R2��x��<�/���C�����;�:5��U�syu�u�ͣ�@a�[��xu��7����A�0	�r]�:d�BP�H2RZ�΋Ub�6��!R1`����=q�sx��2��AҐֶq��H�9�qҷ�ID��u�o�S�r�A8��G�o�bj�T2�3���m�<�ǰ��C�c��a�F����di � �'�y�V�:��˧�7`z����a�16�&0r�M�C�hw���!�A�oy��[�=�y�YŇMk\^{ѳbI�J�f���~G�ghe����>=�c�f�*��8"��4���	3S[4a���S�\:�� ��k!�s�z�ݜ�8E� x�3�JP�&BP�C�!����`�C!)1<��3A'Rp��g������*�(<'�� ё�P�Ƙ�q�,����=�Kv`i��޴3��[�OV[��X��	=�Iթe������I��u�=p�	n��ֵ+�fP����֚��k��n�qk��ܐ�����&]�\[S��5�b�J��D����F��7�3��wO[�>�;�����L���A
�@�u�����Z�z':6�5�NN�w�,4^2hθ�#':T9�^�Vx��ٙ�7aC���������4\f��DI���6!4�z�g�=���8�-èֵ41��zԗ�<����ç����Qt��Ċ�DP��%D��37fK�F�I��@u��=�h�3cy�⒐�FND$�9	BRΡĥ��Z4��Y��X�Y�F���ֲR'q�����팞�یow�7�p
y( D�fꏙ���8�NΝ���2��|�3|}4i\f�r�r�%E���w���ZlO�#DdB':	ʇ,���7��k#��CQ�d�NK��Q�:�f:�5��ˤ��A��h=5��%ٮ�tu7����ן=Cv��P�&��a���I8PFu�uf��Y�!��Pl6�%N:r�ц��J�!l��_!0\P�7��J(��,9�M8n`ې��D�1��e�
o��8*U4$��6g	�2Y�f��Znr���ש�B�V�A8a�ĭL�Bj:X;��p�3]������`��I����2>I.��K5���ؚE�XT�6�EDI����e5��8�w�{1�
����j��!���ѳA�!�/q��=����'}	Og�	No����|�;4�'�|c4n>�h�7��W�I�*�U����y6�J��m�§/:!��ɑ��BPx#��9�@��tjRL֯7="�L(�|x�D;�.�;��i��d�#[��F	k�;�/jh��M�,���	��i��]�N�띙�hȡc�.��T2eD+ާwޝ1G�a����6�D�s*�A�d���5�k0sۙP�p��'���r���&i�:q�v&��ըu��5�K6�%�������M�n4v6�l���u u< u�OZ4hh��|��t�:3V�a��������&��Y��ͦ.dLuf�zl��ޮBRw���}zb	BP���(J�؄ق���Rv<���a��U*n�J���rŌ�\�tΠ�X�c��,�r�4�������{�^�nâcV%9�L�8��FR�Xp�D9q1�Mo��;5��؁�CHh��]#K�<�J�R�Z`�AMc�sh�si��s\N`���4bl@���N#q�zЇY��*��:�Z�ش���-���6�Ėj�z�����TL8�ה���j�q�	�O&!����Q�CĆqą9�2Z!VR��XU��Q��4;5�l��Xuf���xTnw��9���v���$,r��)�j��4�Z`�$�ì�'IZ�KF��&�s��2#�%�y��W%�7	���)�6j�5���͞GP`�Ә'ʇ2�N��G4��3�"��TצU��Z�X��T@��gX���F��]��A�a�j2�t:���#Y���irBTSf���K�*9�$W5��ڂ���鬪���p(ҙ��p��Ŵ@�t��@h����bd�Q��Yfo25&�����26tA�4�a��u��w}zw��a&6	ʣ
cC��Ȧ]�ؒ��<c�Ew�c�F0kY���SPT�FF&b`Y%��6a�a��P�і8�P�%!�' 0�L�n�Y����y�A��M���`�����[8�ɳ}��Q:naP��;;�o��'tS�u@a�n��<Ovg�{�Y��� �!�24N��۴n���W�Z��Mf��K�Y�j�5�����r$q"�(JX32���%�==��a���'�����8FA���@n21�*B�t�bM����`U	X�������C6�������d�h�9Zֆr0�s�FN,2Dt��F��)��8��/#�\�֥Vf���D��eu�Zc'Xj���S�5��ӻqbgN�;���kB��T:%�j�E��JS|�Xބ��k�o�bgWS���b(�A!P͉��ә8e;�3&1���Z�F ���xA-c�z���!�zg5��,92{?W�F��ł�6Uf�C�Q�F	f�M�o�jԺ���mhŉ-��&�v��\�~5�{����U����Ʃ՚D�daqcFo�{6��F-��W�`䘙����.��4l��&GJJg��"2p�5�O�O�X�#0H£���f �7;�9�;A�;换�����
�f���)��7z���9���m>vqs:�����(��s|�7F���br�f��t��:�w;�Ɠ�	<L̂4�:l�(���� �ө������J�JOuto4vx|=��g��kaʉ�����lX�|��`��d��Xk��>k�����{���euu�{���2�$n�};�P�.H|�Ǒ�����&m�	�A3k0O2Vw�j�s\Nf����M�]
i�.����A�`�аh�s��(�Xe>%�F�4Sf�2	pt&8a:Mh-���FHCK9��W�bo1�`�Q��Y18�U�3��m�h,�4�j��њ�:z��2�12� 0�sၨH��{r}�l����n*���d�Pc�E�ߛ�2bQ���Zˬ4 f7sK���}n��:�h�+�k���LL���CƄ��'�=�u	@wd%{�J�J�ёF&k�2Cyb`jO`�4Ud��K�d����r�Xt����V5(�kKL�4kDȇ���*&��T���J=*�p�t�Re�������3zxL�)a-ѼC=Zj��	t�j5l�s��5oC���ϙ��!�BtNkQ���k��vuN�3.�2�A����n��4�l:'Z�������i�u^���dѷ�cD/5���r'�5�f�N�O���E筝�KzZK��3��H�(�٨3ZMj'n���u�Gf^!���M�F�֜�i�5�g��K�'�i�oW|;ӻe��zrk|�tq�{�b�:L���'��2L������+��u�Y��-T��q��:hЎoo�,h�,Ʒ�����)��"ز�����U{�I���5�Jv]��,3N������0HADc�4̃�,t�1��9�@�:�i��D�U�������Gr䥋�BS�|����ީ���G;����)91*Q�9K�HOkF��	]�ތ[G��aթ12q�,��8䍓[׸��˚pō<�(�x7X�`�%`F�I�]kF���v$̥[�ŕ���JDSD���I��#d�Z��F�oC��S����4��l3	jH*LL��ֺ,��#��M���s1�h�E�0F�Z�F{�J��|�4N��іڄ�sddi�Gít�T>�A��dL������{��x�6L�DBĳ�a툌+��^����"!O8SSokYՄ|Ŋ�nG���޻�[4]��:t����.��"1�h�\s�;����u&F��va���1�FF��2L�rt����.�<����X^o�󑳏t�8""@��Fh�w�Ƿ!(�N.F�İqT�������&&qk�*���:
[e�F�m��u����s�E�-�Sf9�dQKDHP�$H�k��7	I�a�����$՚��X�L���<>kz�"����μta�n�4Q�W~oJs}���ޯe4���lֶ�~�{؍�f�cN�p�F��h�u��܄�Ѡ�Vt�Gf�ƧY��XtY��X��:#
�,�f�՚�]f���0h�E��NA�-"��E�H����&(��e�ūuZ�G���%�z;�>ۓ�����N��Y�"dD$X� �*��u����G��h�e�X��c�9E#*�M����iԈ�xi�/�:����]�3��&���F����J ƌ�6�)7�m#K*i�˔� 5J�N ��o͕r���Y��@����"�L9$N��5k����f�J,Sj{[X��ĩ-���5n;dɐ0�����S�M�+�sG^6��1��/�����yb9�d������P]�r�]u����6� tP���u���n�������^�]�����ݘP��!���ZwmW2�l��S�	Ŷ���ldK�vE�� ;���շb��l�o�Zi$�d^
Ĳu�Cu�0��|�����o�y�/~|֧�m���m�����-� .�   ���8�6�[@���$   �  �  h m@E� � -�/       $��    X` [@mְ�m,1����!èڷ�/^�leu�z���R\��Α�Zm�	-��i��ǜ $5� ��8l����$�m�릜��m�A��>�@�h0
�@*��  �0 ��А� ��l�J$;"Y@�   [I�` l��$9&�6�m��۶�H�  m#T���t�q�À8۳f�� � $tv�S�m��ke�l HF�XF��AV�oNە�M�IW�V�8�������[ �SFҮ��≕��*ڶ��\ �}��[��|t-V�e���\,ۧW!�צ�p2	i���[@E�I�Z� $ �[v���e��`4W-�ko�6��@�9.�Ա�l���ȶ��۶qm�Ε�Ӭ��saͶ��l�5P�Z�٠��+�a�M����jc�9��M���j�U�� �mU*��Uu*�T[AN�g;Z�6�p	  m� � �`  z����ڛm�N�Ů��Ā   m�}��񭭮YF�A��6kj�Z^ۖ�k6zmY�����-�@m��P %�V�h۫�	Ug�U���ܯ��V�j���h�HK�*�eZꪨk`ݫ`�4IzC�}�qL���Α%������mn��%s�p;���m��y�u������=�+ �MU���N�W�T��7J�n1��3|Xp���BFٖ����bL�e�����ܮS�UUki3!t�U[@������]����{N��4���yt��g�`������r�*�8���]ݶn�l��Sm�� I�����a�[ԃ���-�u��Y3]��'q��*ڮ�2��7F���.�#���5��0W��z���̧F��m3�� A�m&�Y-댔����J����i��$�v�j��;`��e$��bE�T��m�Z��p �e���f��Zi��,�UU��*��.U@��.�-�� m�#�(��
Id��m��sM�۶��M��8AoPpI l   4�}���^� *�jU��3�y]�s��9#t�i0޻-H۶� ��VÆ�H�Ŵ4�my����  5�l  ��� po0  -�h�!����a��  m��`�����lͮl�Rո%�jmn ����(�HS��UT;�(��0�KPu[@7m��Hn�]6 � 8��@l���ېǇ&�$x�4�h�l8�  B�^lji��X�	>-� N�k    6�  �m�M���u�$6�F�c [Fճ�$�m�tI@l� l�[�5��uHJ��U*�*��]�| Imz�\�m$rK��'(h�6�  m ml�T�f���Ḱt@Z�K�� [zR�픑��G[d֛`5lۯ.m��`�$ɮ�UU, K�-pj�W���X�T���K����m`�� �;�#3�s��W���UQ�[͹�6+�(Hj��qŜL��&�OX�y�ks���#bW	{e���� �vH�E�U  ;+�囶����`�
��إiy��Ÿ�i�	 ��� �:D��m$��HR�@�R�l�`    ��]&���F\-6$   �l�        @      �  (�G���6ك)ŽRu%2��d5�� ,�6휑 m 2��vϮ�}�ݶ [�-����l�n�ei�v-!PH;�۫=d�8]�C]P��+�vq.�ͫ���v��
囕k��֐�Xj��Le��z�ZU����� 6�� r@�/�6f��͝�l5�����m��m{�cE;m�4��вT�OI5�n�i:�)D���k�UU���t'���9��uؚtu��u�,�ۓ�ݶ�h��[�S���m�ӵ�� 	8 ݲ�Һ�xv6S�b���U@ m7fݳ   IxM�ڐ$��;$��   K,�E���-��j@\. �<�r�.ֲۨ���ۢhԒ.m������=a�g,S����YX y)�mt1��6�(:ړ��f��L�,<mvn��r���ݝ�k���M�y��pvw%Hp���h�$a�SS�]�E�l�5����/F��	zN�rrt�q�6�4��T@���vm��H�HH�Ӷ� ְ6�&�-$�,qJ�g���.�bZ��J�-e��Zڥ`��8�Ue�A�a�֭�޶�*��Jxd(�PCb�-���դ��Y�n����SnU���p ā� �M���L���n8�p$����p���l��tݤۭ�6�@���� ji�\���pmwA��i�Z� �����N�m�ר�m��M��8$�n�t�� �����ڮml��Z�Y��		{ �WMUP#d��u��m� m����ZŃQ�UpQ2�p�: H8 ͻ���ݗ�m� m�s�[Xm]�����` �R��+v 6�d����N��K#m��lۭ�v�(���j��>v@���m&�I�[� ���՛Lg �u������)��vv�n�h��������@8ݎU��v�\r����lh�� [^�6�ٶ�Z���
�� mzD�v�p�ۦ���Hl��` R:ʹ�U�m�r lUe@�l�sn��+[.���=��׎%����k�6�&��I5�P	�ʠ��ep]7e����^��k6�8Ht�:ޠ9 ����� �^I&�Am�I 	z��>]�ۓj�Zp^X�$8�I��#E�#m��"�ʫ-�u�*yXsN�P�� 6������l I6�5R�ĉ#m� �vݰN���lH�Wv��BcXF�r�H�mm��h �{n�	$w�o�8�n�v:�r�]mT�g��*��`A��[�mkV5` ^� 6퍶���jд�kV������i79�m�ٶ IĀ �H���h	8 .��m�v���[B��m�$����A��Z�j��^ j�ı�*�nӪ�*����m�  䔲8I��v�mo-�m��V��P�s7:����j.�3m���X�]��;:�`��z�rD��� ��Im   ���p�   v�6�h�` �m�Kk� $�D�/Z	          =jF��Sqڭ�lm��n   $��l��3m�� �I3n�ж��Iz�q��mmXe��� - m�"��v�l     �>   �   p�  ��^�i]����<��U���m���mU���5[�K,�dR�j���n��*�6'Y'^ ���In��q��.��U*��LY9:k�bY��#m���k�%���׺����4^�g��T]t�ݻ��u��f��P�I&X� 9��8�V�m�6���+�pO@�m�Ӳ�L���-&�Ēɺ�s.����/@���!M����H�m	c�4��5(7gK������zp��'�vM��ڕ{j��VIj��U�e�YV�=��i���7���Ɇs�)
[;��׉����[t���V�Ͷ)V�xl Ѳ�m�lZ.J� �[R&հ      h-�A�����~�e9���g�k:����/@ݒU�Y�$n�Z��t�9"�ַlA�ӑ=	�u�v�%�@qю,��uɔq����ܕP��&4ްtV
�U��d�%e&P�����P
�F�����R���cmT�˅q�x���vj��b�v�ZU6�_5U@Si�z--��tK5�  6� &��� ��m��E��q!mx��6��:@ �� �ٺ�d6�n�S�0��v:I:9� ��M���j�l���]WT��2HM��mP�P�6ٶ�]���a�m�6�W���VB�Ua!z�ѝdi/M@v�L[@ �-lO����N  f��;l �� g��}���   m�Xkk��u��-�-剸�Nš�	�S]� �m�ݴ�K�p \�a�qm�q[`1��[��t�;v3� l�L�eZ���+�s��5h �Ct�mn zݶ;[m` s&�[A '5���]�������q.ʮЩ�  �:� m����>�'UUdR����Wc&�9�n�r�]�(+m��xy����aZ�ƷXg����eѣFo%V�+��u ���Yx��v�R�R�YU�����#�� ��� @�n�������%�m� f��m@.!�I�
��CC���km���5��� �< @U]�>�lP��������tEa�;Hk)+��''�j�c�F��%#���0��s��1��M��a�ESH�X�RnSZ10�1R�ffU!��aX��.c�a�a������@@tv ��00 4�04�Ƞ�_�����C����c�5�BT�b)���;�A!����h( ���`�謁L �,'^�t�
zG��Dӷ_Qv���l�P���~'B)��I�r2c�_H�WPj��*w�/�H�m����*|zUD�)�"T�8��|@C�N��G �����=T���₾�"(h@;P� �DCb �(|Cb>
����O�L��TC�w� =<6�����l�ʎ�OS���Q{��} A�#҂G� B�ZONН���"iG�S�} C�> ��:@_0���T�A�iT\A�	8`�� �����}�@) K (�
�(Rv��
�24�b�,�fC����3!D�ID!!���H$&��C�a��%
��T�
t(vz'�P�<BR���E5$�'B�� �:� ���U=� �Snb8���D�,1�J!4
- ��l�	Ҩz��0�)�Q%��Y�e!,�$I+�mt!��B�v�� A�(mEĵ�T6����
�<܎L�I3	$�$�0�L�I3ܫ�r������EUUUUUUUUʂ����������*��������������������������ۻ+�p��ʾ�]�٘a����L����_�k���?������������Z֭��MkZ���Zִ�v��o�oo��������t1����)"���-Jdd!�k0���8��yx�ƕ��m�q�`�۹��zO�6@�����^��{������\�-�[E(��l��$�䀂ۄ��ܳ������kWH���ȵT欰�iU�\�ګ�V��d��sqsc�J�x�l@ �<�b�P�p"��xs*QU��6QC�r�ו�UUT�QvE�T�jP��6�۴� �h���{����Fmg���xgs��r���s�-�i�F���:�G�ni5u�s�:i3��t�:�/=Q�&ڕv�X�秮m�u��g f��[�k���J;s�CΔ
��H���A�ʶսצ�r�#VS��z���Z�N���`9k��yL\4�6�1�����7g"�j����4���fpB/P��m\���E9��ٺNy���-y��l�78�)m,qq�&�����Ed6���T6�U����x<ͫ�0���d�l�q�oh��W8�V6t-v��;Y{�q�k;�O��,bj�ՇOZ����Ьά�\i��t�R�n�g��s�)���)�M8��Z�:��^z�ۃ���#Ѯ�*�<Lvl�+�c�.!��i�����b5H[h�Sy���b\��j���rh��6���.ʩ��íH�"4uT`�@;�v݋����[��Ҋ�n�9^��Cs�7���mPm	�k\v,��s�\1��ېI;Z�UP\k�l)���bMs&[]l9T��r��^=F�xbؤ�Y��Vx�3nʱTL��a&�h ��K�Z�� ��,k�5R�@U�cAݹn L#r�lPq���\=�gC�ӻG,ᶢ	u����hM#�rv_[N�͆��U9��H�'�ĵUT�Ϙ�%�K���v��ֻ]�9�A@����y�ؼ��v{^��Ф;t
��U���Y��b��l`��0Fd��c��W^@�D�m��{�a�#1��=Upq��rq,��=]%�`�e�i�aó�˞��@.�U6d'������z�Z��'�������}�Т���^�~"��������C�U�
��lX�%�K��')��V-��t��yu�m�InCk:&�e�qFm�ג��{bMg�a���0��	m�`#s��8�l$s��nԴӮnr�n3��.��\ʣ�qf^����vg�.xW��,�Pu�\xc��.�/[\��Vb�x�Ev��Ur�"�QEv�X�S�ozK2p,��ˬu������!��"糗fڟ�fn��k6X�b	���:��웇��p��Ç�=��nN���n{=���/{vG��t�	���y������{�nO���}�s���+������us�_h�}����{�hk|�x�T�]�N]�C|=ۛ�;C~淋�8yDy�$J*����qw��E�mT_�\E�f� p�kUɯ.���w�Ѿ{��ݧ��`x?��ߧ?�:���v�s'8�l�w�7h���I�v;���q����Gd�z2�r�Ͻ��7�z����{�hk�G�^�跭E����ݿWk�	tF��Ti4)�E�b��$��R�I�L�֐4��h��jd��͂�� i��{3~���}���Ϟ�G��=
됑Ѫܖ��s��h}��}���ﾴ9Ӊ�%��mA1�u9�:�}룝��w���w�mDV�T%uP�;�h�=��s{�h|�o�������G��l��ۍF���#�����kjy/�ݮ㐘�v�wo]Z�� �g;��9������;�k����"��!��(o���s���}｣|���#���L�+T�֕�G{�o���� \~��ݧ7�N����
�ꖆ��{A�zy���v��;C^�k��j�&�$�Ѿzy\�b�;�q}����θ��$�u�^� ����n��;�籛wc��uv9�gv�̹�\w���}=�����n�����7�v���{F���������7�wG9�T�|����C]�nk���j���(�����z닏ޡ�s�7�v��αg�kjX�%Ѿ{�wϴ����>RD ��T�t�
*>�����$l��y�%��ˇ;��{�J�}��p���'���d�E^�9w��;��όN�u[t�l�j�kõ\J&XV�V�\�9�����{F��S�3g}��]�<��JR�D�o�z��=��;M�u5��۵��$�Ѿ{��};s[�ho���{�R=
됊T�q۟`f.��S��o���7�z�Μ^q�OJ��u���|a�s�������<��g��Յh�C�a �&)w�t�+J��*H��bܢp��܍����إZ��]6�6�������c.�m�a�e���ܜ��c���-��U���Z��^����y���秾�}�F�.䵹�V�.xݛ��I�=sv�7��kNnH��2�z��Y�K�1�l&ms���m ���`��ۑ7i��n�s�R^��n@��5�;��s�fۜO;!�;��(�YjCE{=�/ZX�jx__eݝ�� t�cN~~�|��x�z�;i��*B�(s���F��\9�v��;C��|Ŗ�څ�1�tk|��������;��߽�����t�V�k���M�w�Ѿ{�9�1��:�b�+Z�M��s���|��߻Ms�}M�%)qX��K7���7���;��[�i�p��{���.q��lA���Db��F���5�xl��\tW6��=����S�q�k����m}��K�g�����L�/����V�Uأ�R���U��i�k�������@BD�AH� Æ�
H�P�gz�{}���ϓ�9�i��N	�n�󾡾w��]��;�v�̝��++J7Kk�>0\��G=���w�W7�v�����-���e�jK�|��ό��{��;��O���v�c����^xRO�'�t�q���!n��R�U�y��t\��K9�{��s���Ξ������#�����)JV��G9�S`}��9ߧ��;�Ӝ�'S��+K�&���w�ѾzxX�<gs*��7�v�f���I�ŭ&�'n����9�v��;C|｢��R=9d�)RU�*��ݦ������h�=<����~�M)��{�|vK�I�M[�cɠ6�c��[�|ᛄ���v�́^']�u�}��;��}�|���{ަ�̝��++B))es���� ;��g~�����{�s��-�dJ��9ߧ�9�v�s������x���κHA�UmY�s���ݧ�|�Ӧ��:L1
_P�7���ca2a�.C������#�3z��z|���i��(�}�����%�BI�[t#y��q�d���i��:��a.�X�:,,�V�)NP�;�h�篫Ȼ�z��{C[�BA��*[��l�]�ǌ��ﾡ�w���gF���(��U��=s{�n%�w�Ѿzyg7�/��*6�Q+u��}C\｣|���w���̓�̮Iq���}�秐s�~����=�fb>"��2�f�QAE��*2@8 0>���)e=���~7}�����x�����Pډ��/�lH��V�Oc�s�:�x9��ng[�wX|I��-���`�h�����e�%vr��(�V�8]�ۤ�h7�{������	����;��<�ӵ�<=\���g��&s�᳒#���i(�syj�[bش�Ǯ���M��^ks�Í�*cr�U���N����y�{��w�^2}��lZ��v���,�������3�^݌]�&�ћmqH��-�q+,uYxo�O�s��������h<p�y�l�ʉ#jV�Y������yﯴo���9�1��:�b���$����:���h�=<���]5Ίu�,��br�F�}��g���=No���� $L�Q������������h�\��Dܢ�F�)N��%z�b��h;r��8#c�\K$F���nf��%b����s���uʃ����=�O���q|G}��Q+tw��rt$���v`��繣����{����S��%IH�	l�����\�g�w��9������%R�%e��]��N{�ѭ��9�����y��$y�9�z��{p���h�|�|a��0���q|C���]8�GZ�1��m]��θ\�6��.�ơ9�>��kl{��V��au͌ջ=ﾡ���Z9��<�=�w|��U��M
\E�n�G�r�A����F��P�8��8""f���]������J>�/����ꪪ*�.�ꪊ�����SEU�o{����?� x�e��� ԇݚ4���X���},]vA��6��������%4[cMF�����88Ƴ����ҏ�GaG@X��������z��vڗ�����1S:\b��K,��U�4�M�Z�]�숈�pZm`��[�z�]�!�b�λ���:�w�4@�]�GR���P]w�a v$��dh�:ւH{�F�)�gDdN�iِl}k��𪗈��>�(x�Q�S�� v���J:��$��+�>���t��t�� ����� �uB�sơ�>�����hOy���Mc2M��h�D��Ľ$��2~}������9��4�'�{��d��䘼�����HҔ<���k4g�l��e��L�]m{��yＺ���h�'Ϝ������s�t�	��즡&��2��O�����	�L���b'�V�η��vv���Z�{H�����z�a;l"VQH;e8���a�����3�JS�5�3�(Z|�Oߌ<��0d۝ԩ�L�og�3�f`S+[�{��~s^�:���>���J{���J��=�·�~������8ߞ&�D;�<��L�n~�,�J|��z:��Ϝ����R�����ј�`���ʺ9cp��Zv�>y�W�N}��oJR��>s�އ�qL��k�gJP�V�nX@� �l��;�D�}�ݏP4��}3sz���޷Fo35���)<���·�O3 ����'����/�}��O��ͩ��=�o����xkm@6G<u�������F��Y��GE8�aΝ�<m��]��v?��L����:R����{��R����T��3 e�ou&��2�cxr�I�&���d�{��MB�q4�ٷL�`eﷺ�X́�f�k�2�vd	�q����<��)�M�2S�y���)JO�=���!�2Sz7��p��d	�6���d�>�0�3�z٭����L��d�>s����R���}��)JP����)A�_y�;:T�{���4�K����/I�I������Ҕ�(`|��폞���R�~ﮔ�)>|��:�)O˗���A��;���=ۿ���
tGX29U3lg��7W)�ˉ[�M�r�n��wj�6�F�4�NyLv�`�n��J5%u��9�pUt���m���kq[0&��g$Y'�1�9���3�s�,negm=���Ɍ�ۈ×&�n�4N��u��x�x����N��t�l]�Ƚ�F�٥��֮�3ӻc���d�m�-kkv���{.�h[[M�v���<a���N-�,�Z����a��z���s�s�����H�z�9��6;'<n�g9�ֲ�f��R�������)O�����)JO<���I��R���s�)J%�=�?~U�+n��j[L���=��T��f@����Mhf@̳�zb��)B'g��ǩ>Ò�|���zַ��z�Y��5��)J�>����)J{��t�?`2O����cԥ)��s��)&Y�h�Bp5J���&f�X̃�=��}Δ�(|�scԥ)��}��@L�q���ԚĘ�s�ʉ%�$[՚�t�)Cߜ�ǩJC����~���Jd�'�߾��{��=���R��_ɿ?�痿���|��fŎ]sm�8�9zhq�"qͶ�ֱqö���ۃ�˾�3u���u��)J}�>�t�)I���p�)����A�� �.�(~�����0k0�/���iYI	l��Ĥ�=�C�~\�_�����S����)JR}��4=JP�O�{�gJs�)�������*%�rI%K��k�3-��:R�����4=H~��)�u�tt�3 e���&��2���qk���!�{΁��I���iz��=��tt�)I��y���J��=��>�JR�7��g�ĸ��N�����3 fY�ގ���&G���~���)J{�\��)JR{y�t=JR�|�zsEݲ޵kFݸ�f���8�=�#:f�!k���c�b�l��I]U�q[�7�%�%�~���|�2S�k�gC�I���I��R���tt�)I�>�4hʾ�7�aD��k�&���s^�\3��i����J'ߜ�GJR��{��t=���s¢`��ǐ"�zI��->}懩JS����wO ψv�H�A���ĖU)"B���H��ZNpsπ|�]��·��2�#��2��	�Ql˻��EDT&��	�,�L��2���'�M���0�J�r��t=JBM��6)�N�
&bU3 f@��z�(��y��߳�)JU�{��^�)O�=���)JO�_Ey��f�oyj�V,�fr��;C�w�U�Ͷ�e�5���Kې��8?���_�ލ�El=}���x�9�_�gJR���|懩H����z:҆JRyϼ���)Js>�2~淫Z5�c���)JOo>sC�}�⦥[�ԩ�2^����X́&����2�5�%�=�?�VV�)ky�B�gr�9��F�S%)<���C܇�!ܜ��}΁�)9{�JSߝ��WQ\�Ȝ���>A�cF}��I�f@̳���2X}��n�d�@��}�������y�J2_op�Bp9KK��Q34�Ę���s�Ҕ�`y|���=�R���tt�)o�>�á�R�����d~0q�t\��mW��t��.���w���2ǳ�q���ݸ�\���N�:�̝�ixŶ\Q���y)>�����JS��}��JR��~~��~���rSߺ����(~{�3>��GH;�;�TT�k�3,�ץL�n��;&�)=����r������7ҙ)K�����,?�1�Ý�ڮ�%e�B[)Ҕ�'�~��C�)��3�)��R}���R��9��GJR����9��mr7h�W.���0k������0HN_=���R����z:R��'���Mc2e��S����(�v��/L�)I��=��)H}�`�~�t�)I���O�r���9�]JR~=Wp��#B�Lï�k~���;kض�N����,�3���m�֎k-����;��P�V�R�������8݌�� r�M���%pq���0JcǮ5'[6 &�Us%�A��J�w��<5T:y���Ǘ ���mu\��;Rrh�8]v��̘��kWӤ[=���M��mZ�q�N�!�1�^m����]җh�֑��7.���w8s�F��D�:M�]������u�H�',�����^y<k��Ky��v��y�6�;��! ��[����J�j�ei�R
f�l3���=ߺ�3 f@���ڡ������Ғᙜf@ˌ̈́�3 fY�S1/'x��r"U3 d�����Mb�&q�gF�)JRr����(�{�GJr 2R��}�����l��X[޷��)J{�\�gIܹ)@'������������JR��>��Cܥ)�>��u2<��w�%�&n�'dɚ\g��R!�N{��g@Ҕ�<��:�(?B��y�ۥ)J>��֭}6f�u��Cܥ)��s��-`9d��Ͻ���ϼ�ۥ)JOo9�%�~}<�|I#���bm[j2�>�z��T�b��s�R@������\���w����}[�V��Z5��oJR��9��z^�)O��|�R����縟a�)O~s�́6��M���t�f^"&^Z^&�X�)��@}>��_R@0��f���*]�]�U,#�w��4�����4� �P�� :�N:�R`(����JN����ԥ)��G@Ҕ�{��t=��E�NgӆG�5��4kZ�[�)9�>��JS���t�<�)�=���JS����Ҕ>I�y��8vJ���������k�~m��T́�,�[Ԛ�d�ۓ�3 L�g|w}���>�'�X�Cv�RSY�������{��>�L~���(_���t=JR�<�ގ��)=��k�˻c��b^��h�
��8��{-�cIͽ4�	r>���RYZњ��F�I*B��]ܥ)��JZ�2N�s�R��Ϟ���)I��=�Cܥ)�>��ֶf�Vn�hַ��}�%)<��t=GԐ2Ϝ�GJR��=�Ͻr��Ϛ����HϖΟ7�F�_)T)�tA�R���)J>s�t=Ó�~	P�B	���h;:���_���)JN^{�Cԥ)ﾶ�ݸռ���k[�Δ�i>|��:�)O~k�eҙ)C߼�cԥ(����z:��#x}��U*���uQ�%ћ��=�^�:R��2�s��R��~{{�Ҕ�'Ϝ��r�|�p����Ή�s�9��rz��;Jy�.:ݹ���D�d��=����q]���t�Q�#��JR���cԥ)߿=��JR���{Ε;��=Ϟ�[�����}�T��㣎��Zf�`��w�}�X)I��=�C�)�=���JR��}��f�bY�=��,r��q1�)�)JO�=�3��R�����t>ɒ�>s~�z��;��)JRyϑ�F\�6a��������JS�{�5Ҕ<�!�\���)Jw��z:R��u���MJ0ia�Eh��#�P�w�I�f@̻VC�J���0��t�)C�=�c���=�;zR����8}�{��d�g��.��)>
����cHTc<q�F�OU�j݇G��$����3�ٻ�oo�>�ܪ�'�n����ǸS�yεt�)I��·�JS���5Ҕ�|�ݯP�L��ߍ�UQ��ҫi��i�a���f�aJ{��5Ҕ�|����)J|��z:R����#�v��f��m�}r�����JR�=��v=JR�<�ގ���2��m&�2����LC�1*(9;�۳@g�h(vf݇2fL�����r�߁Ö�Jp�qt�p�)goq��c��P�d�[�7�o�r׿�wwUUU7owwUUUwV]�UU}��32�9�y�:���h�� �|�M+��h�0I���F����՚g�2ϗz�����X� .�C{F_7w���E�ac�8��b�d5�f���p�Qk� �Hp�Y�Չ�MZ�(#}�`	l�т���^�Č:R�>G�s{R>;S�Xcwn�68Xb�F=h�05�:��!L�kf)��9�zC��'������$,��׿3�z�� �{ 4�h�G�a�jRJ������q=�;m����s��
F$=ɉ	$e�̳y�SA�*���2��X��c�X@���M��R�$i�m����������a�QƮ�'I;J�i�vs��ʃUQ( �$i��V�q�藞����n����Ws���=:g[�v2E:���6�.�;����\��ĥ�ꁣ�N1�n���
��K���J��"�΄�'D}��w��+�!���%Ut
r�/v�ҽ;�궙%I��+��Bj�S�� MK)1�n�;i'5.���26�ٍzi���;$�7V���7mv�HGZ��)�l;�h�4�-�㍸S%]R���vS<�����(M�1����J	4���l �"Z����ں��e7;v�}#0�[��X�"躍[K�m֔^U��y�Z���C2v#��uImʽ>HЍ�P.��9�BD����PX����ka�l m��m �9�;M�4�n��v$�F�e�1x��#�#ϴZ��3�m]���z3Z�uc�=�Y���4�m蠖Kg� �hMq��A���k��]�����)���a��k��,F��V̆z�����·Ͷ�۾��4%��;��;)��=iQ�^Ӷ�;d���m2� J v'=Q����t�yg��읽�c2 T���ݢ���tp�U�i�]�xG�u�8ﱵ�R���{v8��c؞ڐ�#՗�q��ڊ�:�	���lp��+ɹ6K�bХ�K���s����;*���'���K�.҆�����ͣ���#'lSê���1ݝ�ݥjS���U�����`�N]�ﴔmZ�e�mt��u�)m ��S$Şy��K˥�mn�(P��j�;�k�8z�1��%��\q\�'=Z�\]�wZ�Y�[(��]�L�ت6� ��U.��Ī:��`ͪĜ{�]����m�$=N��ӷnݱ��j�a�C]S�S[]	�8��Z��˚�e�h��5[�pƫь�iG�p:&M�����v쨽v�(^Y[H'm�� �jV㞸:N��gHR�)-T�PslŊ�`(�� }�����A:~l8 ��`��ق���@�U� ��3���ҵc��18Gb�*9.4l]i�B������%���v%[l�7�9��X�fU�r�l�t�����;�������r�f7V�6���y9��sR���V����pK��[j�!�-�3n)gP����2Kۍ�g����.��O	���(���jMt�r���{9��%���FћZ�nɸ�g��������R�Y#�ᙘ������D�ay��#�gӅ�ބku�՘Aq�s#5��������Z襡�b)��_����bKoM ^v�<nԕi����!8P���w�	f���k�=�QA�w��܎)7� �Q��^��|�ڦ�[罣K���~��Vdo= 33_�5;�w}�pQ_D|K�`fwTT���`^c�`��s>�����L�L�v�]��=ʂ�u��ڊ#7~�WC�1h���X�z�q�s���[i��{fxF�c�z3m�(�-�ym�D�w�{���O�����u��ب�3�z�.��}�.I�&u����uU�=�} ]!�	H��PI�d�O��R�/{v�z3^��u��*S�8�r݁�ި�H�޻��;ʀ;�][�kRږBM�9�q*���ݻ��b�7wf��d̝}���vC���(Ré�����Fr������ڊ3�����;�b5���ۥ^޲����vۉ�{3�Ex5�=���-��������ix-���|�>[�4��ɠ=�ݾL��!|�7��?)R���3)���.���y�|Fwu���T���(���33�m|�
BR�4?gw{�f���"��j J�n����U|�=�*����̼����̝�$�{'y���4��ȫw�ɒI?�n��V�G�ءdlM�Z�Isݕ%Q��M�&(�޻�;ʀ��:F�1��V�!p3�g�.����<�ϗa�lp�����7f(���ҭYZR*5iڮ�_?�b��ݻ}���I� d���MjB܁Ωr������J�۠3;x�I�fF��۹4�ّL���դ��'�PKn���T��tG���"���v�&K|�h���1��y����&O�����>wE����u���p�#"�i5�I��iQ/P;��]�U^}9�*R��s2�	�t����h���vw� {�z�oB���r)C���P��3/=Z��s��gA��(6X8"}n��nz3�`G���W����
ۤ��߾��3gyP����P�렃���_K%�D<L����v�3^��L&Ny����`��3�ͻBd}X�m�raD:$ڠ��@�����ݻ�`f�‽����dp�Զ�����頃ݻ�`f�� /;]��9�)�H��b&&&h���`rI!�n�yϼ�U]����W�.݃23b�g�����$�crV�e�I�\gh[�we�u\K�mS�nX%��yv���.��Ŏ$��Y�f�ܘv�*�U�{Fu��˻k��a�Y���ʫhx��\9�[�����;q�区�T�,�����˾�cg���\Bc.��Q�S�R`�0��\Gm)`vY[�i|�;:��%�����KM��[7Q�����-��!�Obx�eZ�[��sa��[ӌV�"r�"��$��n;��>0����S�,�����-�n�94�C���̾�?��* ��t{���i'v�]�ڵp�&!<�!�<����nMrL�?C���3}��`fFk�2fd3��,��#�b"T�(���wt�{sn���z �ܕD;�Ӓ�>N%&[t۽v��*�����@|\n��4��nS�r���݀ff����Ή���wI�=�ͻ�~{�߯���2q�	��e��;���w��<m��]:8��]k^-m��ݟ��{�2��BM� ��ty���@�w�菬7y���z�I)�J[��=�7��w�q A�T�z������װ��̛��2d��9��y�x��N�,CļD� 3�z���zL��@��@y�7��HrT'O(D��"bn�Lّ��{��@��@�}������R�9��B�0����u���3�z���TB��9�3������=�O�v��X��0�ӌ\q�Ͷɝ<p䓨Qh&�Rprj��])uM��;��۽v@n����D�}�6���.e�� ����;Ш�uВ��u���tCr��mC�j]����{�4~I<�IK�H2dy�[32_2���ߦ���v�>�N}�С̥ �j� /�] ^溂73K��ɒL�;�@{۰���1/(q7T��i��@�ޫrw� _{�I/�f{�5�U,�\�45j)'Qn��=�>{'�m[v̼j�����W�L�g���BR�Ӗ�������T�ݘ���@{�J:aBpC�Q(r�����z@��܌��S@{ۛv��u
F���nH��� _v� ��tfv���;ʀ/ѽ���s2�(sI�;ws�3;z�7��E�D*���T1�Q�詀 x���hꯙ�tM6�S�@�ۊ3��͠ݝ�@n����;�d�ɖo.�C�<D�k;3
�ű{f���m��N�d��-�.�/)׷!1١8�C��)8,J�~���P�k�nk�33��WGB>�p�06����� _v� �nà3;z��|P�ى�hr9%4?���� ��t�F��������n�s;2��R�!�岑go]��ϊ ��t��@{��ġp�2\��=������t��qC_,�޻�"P̴f�.��N򇉁L����:�'�w�';U䉩�z]����V0�Yٖr��l,�q�����c;�*�Y��[�͜X��9�`��VÖ�p���'����QNLZ���MSE;i�iZ-�:t�9�`ި�k�;����'����X}4�L���D�Vnj�|]������8�[����sn��g���D�ڇE�gŻgd��]������������M�Fہë:ۧF���*]�qϻ��N�ǘy3��Of�>�tu ��R��{�� f�3����=����F�
bfy̒��D�����@fnm��(�r�rk����y�EL�<)�D�3-��߮�������{3]��:"zRpBm8`�݁��� ^�M }�d�rfL����<��8��JJS,����tyfl���vٳ���97$�wo<C�J�)�����u�-gq��$_je��N�+(��q[��QIR���,o7�-�K����B�7�����|$���@f�9��p(�ȕ.�����{�I:d����|�hG��	B@<�ڤ�&`��X�!&	*!'�SHih����b�`PcUD�T�(PL�3@@|,M�-mR�X������ff�"*����I��=���}����qH<�6k��2?�IB��aD'y��`}�:�^�rl�9��٢w�~��;#y(��X����$ɗ*�w/w&����T}��`2L�͝(��BS3�d�Ά������G��G�w�����/;]�^In�~3�`�U�wijghz����	&��@CIA;�4iD�Y^��j�5m.:Z�J73�w���Δ~ܟ̒HfI5���ؠ;1�(�w�<�<̱17`g�t����>{"��s6�vfI�~\Ώ�R�8�ܕi$���]$���M/���e�;�Ye��UUTݽ��UUU�YwuUTW?~�^���}�y�ݒHD�@PA0T,3DTDB@�|S�X���Gk!ƅҘ�A� {��b���h�0�Nw��-�����t��쌋'D�H����5�δ�6�Ll���c�NdXGfވ(�� I%�J�iBe-���i �g��n��:�"�Ў���������aCP^A������V0Xlf�S��@�)��t:ш[�:�������%�Z��� n5���ˠ�`�b�e��kdb�����v�4V�3��v�hAko�� ��bx�!��? �E1�(iQv�:C�<<T|^(��Qv���8 �
h�?*����D�~* ?"����w�_s|���^'�jc�8pܤ�Ȣ�6��3;���y]��ϊ ���X�y̱D�\4�)6���޻#�ϊ���@c�}4��=�O��+ �eN�T�+�[-ۧ��x�wR�[U9�r��d�]v���~9��w�1���˫��%@��i�f�@ٽv�o%��9L�Բ�/�΅	nN��޻����	L%�eK�h�����A��� ����$�g;:xT����ϼتfeʉ!(�n� ���`nsℑ~�䐔�P��٠;�\���wD�Kv�>( "/ݮ(ۚ�vo]�׽�~w���o�`�y4a�$�t'q�n��Js��[.=�9#<��-�����w�7|맒T$�\��΀=���~���,�|P�َ�G	�I�]Kn�3M�@{�z��|P����jrɒcJM�@{�z��|PD���jY9���ã�����݇&L�s����ݤ��=�@_{6���wTТG�%D"^%nM�!?�5�_;z����:Pc�I�fF3ww�~?��6��5�l����QPlq�vi�b����DlP�J�t�NM���C��Û��ո����w�mp:VM��T�=ϛZ{b&^�t���4*GL�nSӦ;u͸��8�]lv����~Sf��=}�|���`��fβ�5hj\r' �<ah|�W�͹}z�;m�.��d�ӷcRb��q�6!�V��+Y�z��+v��(�C��'y��kqk�\kۘ���]����:�]u�q�{N�/]k����v]����}�S�	������79�@��@o�풛���bD��a��{�z���|�J������" ;6: ��8P�N���w>* =��G�����36hvo]��zc8�	D�w�I)�P����5��޻#�o>(nGD��Cr�s)Źm�f�: �>�voU���Ҫ��{����ԭC�*�7=�\�[���s*�6^&��=ury#�f�"l��SW�o����m�nΔ ��)�����(|{V�%5�@ܻ�;9�J?�DMW�(���� `Lբ#J�h����%���hϾؠ>�f݈>�4r�(Պ�I]��[K��WI/>��i�3" �f�݁�ϊ۱�*P�L�p�T��|�3&InN��o�n���0J �-�������Ϣհq�RtMIe���w�9�@b�٠+g3f���������'�i�����s� ��-��s���pAɬ%׶�<,�1hͶ�w����������L&ӈ8u`{��@�k�n�}�f
�ϻ���Kϧ���t�GTJ;@y{�hY�% =��Vw>*>�� /r:Bx!��əqN[v���|�;�?�PR�!DIH���Bz�	|�2�z�@o�h�)|y�"�X�.e��ػ�����jA���?�'I%���@g��ĸ�;�H�Цe݁�ϊ���k�-f����뽷������E:�瞌�c���^y�=m��ʛ��rnͶ����Y ���x͸�x�W1*��4�{���6hvw_��fe��=/@{1r���!�Jm����鿾�;w����� {ݮ��g�%70�����M��뱥�Ө�fH�ܕ@y��&hn:Ԉ}O.&c�m��Gۜ�� ��5�f����蜄� ��$��$
B ���"Rd�Y);��`k�jq�	S
;�D��v�i��� �ގ�;����ؕūS��.9أJa��uos�>��a�m��ع�B;��=�z��q];?mb�*e�`Fl�*=��vo>?��AK3�;;�rrɒ�iB%�T�guؓ(��Ҁ/�ɠ>�|Ȯ2N�9q.:!�aK����;zx���٠=��
����3�䢢ba̸��PKĔɒ���X����{v��������ÔD;��O�LZz��`/ln�k���37�;��ޞ(ｻ��f�BR���
4%#R'd�T�a�!��!����Ih�tf�sy��7��v�O\lT���I���zͨM�k�e{g�Ƹ��~7C�V4R�n7Om볃��i.r����y�A�U�mt>:��[�
P2��9j�&Â�֍��������v���M�]n��Н�=��Uk�i��r#��2��n<�7+v�t�N(F�-M��T���]ӫ;��V��Z4sV�m�m�ӭ����cٺ��{sX^ۊ[�3?��n'mN).6�tm�����I�;���t��(�mv::� ����{��/��JnaJ����)�P^�����|P�����Tw�: ���L9c�m݁���z��3;2I(2�U����mX�L���YŰKL(xt��X����;�(v�]��ϊ)+܏�S�RG\tݒݤ�0茶zIo}�v�gG�$ɒ2fg=��oC�I�2B�(D�j����vY�TE {�΀̝�@f�[
Q�E32ᅶ禓��/lp�-<�a�z19�	88#���ջ+��tD}(�PЉ�
	p�\�ϊ _}�@}����30�ݻ�f��P�oZ٭��kwU^y������R$@�S�S��Z��������sgQL�̀������D������{cu��nݟ��w��SP��4��{$�U䅩�N'k�Y�`���}�{7�,9,ͧ@DD}�Nj�;p�zN���=��K�}�7�7g�P�;��#;a.rL�3	�%Z#B��m=u�y �N��ͧ��nԞ�#���w�ك��F�t�n4;%��K���I#���@_gu����B�'�L��*"U�D́�F��&H�nڰ=��js��摆%ޯy��C���;+�K�|�;�>s��/�`fBR��bC2�� C$A�`�F���LIV	���Q����ݮ�����5�����ō����P4��DDfvңϳ6hz7^�~��w��w6�uY!YGH��i$���t�0vw�I۽`goTP���9�i)I�i4c��m�6�9wN�8�nۆ�cY��F��]�����R�J��oNG*B������=ʾ�w����*(���Z���j*&fG�D��[w�$��$���@ftЃ�1�}�.��@M��3���H��:?G�G��"=���ݻ�`|��8���0��<�L�L� d���T��@^�݇���) �# ��Җ�t��k$�~L��"�R�(�O���<�$<*�"f���u�L�'I$��Ž_��J�>C�{6h��1�J�2���q�m\��lgM���o,����n������ݤ��LL�&�I,�.�Km]�]��`{ٴ�{v�2L����u�p�=���J:ˉ��]�J>��lс��%Ͻ�@+�f={�۾L�L陙9�8��B��2;
i$��~�Io��zK0$��f݈=���/>��w׈x������rL�>��=>�޻ۛJ�ff%�w�t�ﻋƭ�lU��P��3������@g�u*A��=�7��zֵ�kF��kZֵ�hֵ�kZ��yϾ����7��y�LF7Rҳ�f &)�e�`F����&�!#[���tvw���j|[�7�s�Q�`���zE��H������6F�1�����1�&��I�$6�Am$�aB��^2m�����J	 z�)&I�"�j5�{N��:��f����Q��d����&juc��:�gn�0ز�1��|N�F��,�3�oI�z��eu�VfAf8e�S�fbd{��(�H���̂�*>V�t�d6��8R���� ��t�m�׮����tQ�	����N�.�2AIuH]���Ӫfu�@[�a��Q�a80Bf�/).�hEN�s2���ٜ9�ۘ��1�/1:Ke�lݚ����`N@w�Nq,�E��3���"������$��SM&���aKg+��@�֓R�Zh�:	*�:/D�3��$��l�+f���z^9��h�&GR��n�'P�c^����s��.�G<�lJ�Bܐ�P�
�K���=���7�-ǡ傀��b&�R��lE�l���}�g!���KS�ֱ�J�L�a�Y�ښUu�cUB����˻&N��%�*�W I,+��⻭�rf�u^x�k��x8�[zf�k&Η���5	��/�:8��/X��ݶ 6�t�h6�E�64�3j�kt�͙"1���n�+��7�a�<��Ip�g�	e�^�;���ms�qgj�@j
�UÈ�����y^�֋r"��9�볈�m��֜݉	���'hw,��0씋�.��{;�,h�y� ����]۶۫��&ͰP�+>'K��嗢���h������,��H��tԙ�Dpp��A��l�������܆���EƳ�2g*��+^�2�ݡf������=6*�cX,�:�Y#������a��.����u�(�rl��i�$�0�F4���j5�xs)@�z���n�rZ��k��.��b�) �ӷ]�vm�kF����6��� 6ض�*����5X�5�s�g�p�l"<����zh�u�Xf�;4/C���I'�����'��)�t73�q��L��i*����͵]��y:+[�f�{�>+�y��X6�;��N��b������»n*����˪2g՛��ɍ�"F�/-�q������p:mb�$��.΍�[��-��^�!�dxx�F:�N+�	��ꗝ��T%�ZwdW��8�Ie8�/�_��4PQI_�B�J����`�:~��}�m~�����|GS��S� '��H>��j �
�U���<JD���}��k3Z��[1��d<]��v���g��X%RÛ�f�{���a^ۜ�Y��Lc�^�0ar�J9�n�����R�s���V)1� 2�o�/[1H���9�+%�U�ۇ�����ז�7ny�,�Ǫ6����-l�bE�j�uc/a�Ӷ���}��֠3\��c7;e6���p��۪�l�)��e�xk-w)?��0ݻ[#�Ilv++��)GN��۷���S��,l��,r��n��E�`֚*oP�'c'.���TP��*ޝ��t��+d�'�;������t�;�e��=��T�;�����H�ꨬY�cK���{n�X�eܯi.v}�/�����ޜ�@fCeL2���KmPx�">^��vf�ECH��9PG���T��pЂSP�˻3z����9P��T�w]���������r�}uu� ��K��v��7'
��e�ݓ^�Ōd�qA��"٘Ҫ����D�.(Y�1@^Nh�����}��Ԩ2f��:!��y�%=8�P�ֻ���y����	��ʘ� �n���v ��������eKȠ������}��`{w�(>�><��5I�jt�Q!tJq0��9wdfoTP^Θ��k��>��;��ű�Y�T�nb�Zi%���$��o��t@_gu���7M@���[D��|�>Zx�]��9O�I�ŝ��v�2Vy
��<8N	M9��˂ܹ�=��� ���>�m7�Mi�8y��a�`6e�&H����z��obI{;����������Z�hD���L	7v��Ύ���|��?�C�،��M��16�ׇ}:��}�v��Z�)yyr!C�J�I1��٢�6������n�E��2�I�2���j����TPD_v�X����������m��LhB��W���<��������#��{��,�t�������&^F�Q)�Xwo+�>��T�ټ��ۯ��ȍ�NI���n���J��������ۿ�fd��~Z�n�S��&"eP�Ί��҃�_������Q@f�.�W!��rLJ.bbÓ��k�)����=��J���}EN���<�>�!��*
�$%X`	����*��`�;} 4 ��uk�z꯾�!қ�K�%
%6P��u�����9��zT��#M5Ht����gg��[,�1[���ԧH��͢����ض�=��M�-�zU��v#�]m%�{� ��&��N��۰�7��ZZ"a��nr���k�耼ǥ��}�i.{�M�7���q���jJ>'���o�x�=��v&�6� _ۓ@f���L�8�	�2��4�=��y����ǥ��p�Bq3�e��~�33iPɟ�v��nN��7n�w���h1'BHX$!�2�Ӻ2m`�-�:ce��n$���s�gE��g�ys���
��uz��ٻ&^�Y"6�n0:��c\]9x�v[�7$xLٱ�6����p�0l�a�9���C�mNQ^�4p��������N�*y=q��an�����	P�)Y�m9�:E�G�n"���x��um[a��m��on����n�6�ƶn�n#{]rl`���$�Q�cfg��3�0�����Ű��7h��<n�ӌiG��筐'Zق�	�N]ۓ=x�:��M�M* ���y����K��L��77�j(��!+��nF�[M�w��}�vy�2v� _ۓ\��$�����K!K�$�Se���]���H�/DD33�ޕ%�E�M$����rbsT}�}�ڊ�ۙ�t�9���b޻8㾯�%��)�Iˊ �f�@3$��G����۰>��T��C��=�f�&v�.7�䞮�\q��!�a:�=sg�:{Vn�RR$T[$���t�[5n��\�=�>�f݀���T�& ��&��y���ʩjj�Gk�K�w�o�N01�b��"i�\�ގ��;�ϻ���¿3&&p�x��ߔ�tI2��7�ߪ* =����ǥ���F���A�x��2�932d�I9��>� =���3�wE���7#�%r̷#��n����">�f�X��K���뤖�ԫ��ev�)er��Q���n�^x<�Ħ��A҆�N뎺.Ǟ75�];Jp��i"l�=ٽv�z��/ݽQ������f���NX@��3vٛJ�$�3�}�٠>̝E�{6�$����8��(���	�bU�|��u|�<���u_���-$��D	!�
!�2 ̀R�M��ɒ�O���߻iP�툈��2�"j�US`}��x���7�m�fڰ䙓�n�P����4��G�<DI@_{6�d�!goZ�>gE�<����y��V4�[]b%i9��c�=�>|\/�$�D	�sN����b7;���ܦ�K�;z�����>�Nꯀ���.?Ə����J�i����ކ�[��T������)��11<̷$�)��b�̌נ>�fݟѝ��ԩ �Y����`ٖ�e8cI�Z����޻}����"���<���[��1 L�CA � ;=�}�:����/�i�'aq1Gn��|��j-q��'t��|P���`_�퓄�Ԧ�1õ�=]�Ɠ/<��)�f� /'b�7��]cS(�/�W),���� ��6�o���%�cҀ�f�;7�(ln��ʞS)Á��\Ӱ;5�@{�z��3��� ��%W&vs7ڙ��T�yDDĊ��f���͵`{rh�N"��=����"g�ݐ��)���Жv�(9�'�f��?-g(%;L��C�˔nM\�{2��3����5�P��<Q~�)"�~����w�����-�;<$Nj���b��4��WJ�V6-��tX]�]�y���۝�ۭ*��&T��� �zAݎ�'m����:�b����h����+�4�ƀ��Ŗ���]n�u�l��Ļ��T{uv�@ε�f�TI�c�u�#���5ٓ2�*�t{cj�S����g��m.-�F����]��Ϧ�����y�v��r�-W#�9Um�[ep��� f��c0��7�H�VK$(��/n˫;�vx�Y��v��]��.�όZ���e�ٰ�-�e�4۰?d�r�=ٽvJ^������t�h��3,�I��\* �}�W�̙��oT��f��{"GP{?#��4�È7v�uE _�]���A�7���8�%�%&�S�'O1*�����u4z3^��fm�f�Ł�aҦeO)��he�uC�;'yP�[�`voR(����;�|�9r[]x7g\m��̼���:N�h=s�Þ���J�Ņ��e۞�/EW�u�vUiP�޺��� ��@V�+K�f4
�%�!< w��}�J�$�S0%�@#��U�u�}U��ҚP{�z�?�#��|��'�I'.U /��4}���ڰ7ٴ��ؙ	���ĢeŴ۰;5�T�7n���Ҡ�C&s�v�=���lDI9*@�b^�����v ��&�޵~w������ȥ~Nf\�s��p�vCf=c�<���9���L^��vO�w��49�a�(n�v�"�/ݮ������i����1o?5(�rfD|����G��sTP�o]�ٽQ@_�)R���p��p�:vd�-$)�}��q��>����ѽ�{ֵ�kT�������UUUUS�o�ٟffo{��R:r`�1!�!�	"�(	�"BZX��@�s$��3����hG4i5f� �j�^���Gf����q(4��S��顬	YC8^D���A�rs�i, ����/Y��H���^vĦ�Юc`�u�A&�i~bddP`�È�� ��f��dK]xi�<�b`d�6�fZ$�ȉ�&b#��a��5�)� ݁;3fh3��Δ3�u�]7����@��`�W�ZS��)	�]�����c���I>[І��y�3�C,$"t����?������6YVkY�@���ݶ�>�lb��u���¤Z�1j4�4�t�5�i9��+rf����hlf���8V�]kZ��i��q9$֭��a�4솛���a�a�4a�`A�����:�����0��	���EI F$�e�&T$�>�?�Si���"�A��4��S�懊�v���T=D���b�,��D���Usߟw�^�s�Vܪ���Gk�_�3Ł���~��z� _۳@g��z�s�=���Iwt�!�n��fҠL�_۳@g��T�;��1$gJ64�����m�qlf7i뗧�x]2�u8��>Ӷ��<n�ۋ�G�$p�̥ ��
 �wC�7Ӛ���Ͷfd��m5l�h��Ȧ&`"%E��X}�\�{ݽv�z�o�}4�Ďux�^��F�QUezŝ����oTP�Ѥ��ͅ@fg%�[J��&���mf ��F���{����{�W�3�+��d%���" (��{WhlGb}�ն~9.�����B��K(^�2sU�޻3����D�:r���]X���˺v��w��j�5��ݛv��s�>%�%��=X��r;��X�wWi.��"�{����޸��7f��ϒ{2�*Z^�y���f݌�&<����nE�Fc��s�3����x���z�-��N̒`ϡ{�����|X�mPJu0C�fU$��glP��z��۰�왙voZ�C����C�r��i��;gyP�޻�v� -���@/�'f�,&e�iu��==d�	h^���26�,Y����ų��$+����\j�B����b}��i�/�����۩X�c���٦�NU�yV��裣�ɒ���9��3���ݻq1g;��]�)�u�$8^4�
�Q�hi�x��<2�����̍]m�%�.Ŏf��\<�lN�v�[u	a.�����\�9	M�c'n]���u��yf㫱4���'n��݋vݻ,�k������S�����<�������|�x���䴢I�z�Y�v{smX#�{���ܨ�3R�4��?�	M݁��Q@Z����j)�;���>`fc^��7�4[Tn�6We�K�wD��f=�3�n�]���E;߰}xxx׈yiRZy��Nɒm�ފٝ���ꍴ�����O[��50I11@}�j۰&f[����vh|�M$����5���ꄱ�!����]���l�i�c��j�"m�����۵��������%D��;��(����r��I�p���<�jq��%:�!�y���W~���P9�H)�J)�(�$
�
B��&���+5����۰7w^�Px�.��jˉDL��M͇!gt���3$���[�$�n��yL,x���Z\y���̙�ً��w�R�3v(d�ϙ�@{��}D�w	�- �<������~I7ѽ�`c�lQN�{?u��>���\�e���O��T:ۗF�q�8ca�ۆܖ��qϋ+��N���j�(iˊ��M[�4�;�#�7{�(�)�S��p��S`b�ؠ��ڰ37i��7b�f�}�bce�eKK�D3�3n��sv���!$�&C/����<E5�[�@|���B}R�@�x��Ksv�o��@c�2(?'�gw�>-N7(%:�D�2��vh���;����Ҡ>������l7T;姱�����ĹӔ�����Ll]i���{���u�;o��ɖ�n�ս�@{3���� ��t���n�8��@{3�쏾�� �ݚ��dW2I��v��.<�y�,��6���J�/7T�Ƀ��dP����3�K����N	n�9�q@{�4ތǠ>��۰�%�$��I~d���2b\@�jrUC  � ?JjD- &``�h|�3%��=4���DDr��T�nn�Š͞�@g�z��ou�K����}Ue$Zn�EՎK�zۺ�<�����b�vu-��}ﲿz#�m����n	�����`nnҠ�7e�P��z�s�^֡B}R�@�y��77iPٻ4z3���ͻ�$���V��C�L� ��΅	g�%0/=�v@{7��(�4�p9L��q6���{����3��( ���#t�s����͉6ڠ=��vwuE��@|��}Ϊ� �$�
I���c�l��7P���vyK��9٨�48^Kg�N�Jf�n�g�8��Ǳ�[m�"�!�a�0IذI�'c�tl��v3�j�uѮN�	�N�T��8wV3BQj(�vd3���Lk�c��MǮ9͂�;�����b��vm�d�8�*��=UQɬj���H���U�N��R�2�e2[!�7�ֺ����ڜ�h���}�]'�t�$i�䧢��+X��q�y,�\���ݚ�}�\�ݮߞ�?Ȓ]LB���q�j����P#��ؠ=���fo]����}-�m�72����1f�В���#7�������"#���T��wy�������3nn�7{�y+yD����Z��4L;���zd�?���`��@|���;���{~�&̂a
$�.�w���zhl��;����݅�nH�ֆ .#q�*o/��`�Aȸ�.z�R[l˱%H���CY�"�
!Yn���{��X���o]�n�: ���J��ܸ�4������|pY��2d����Mo]ߝòzh�3^��6��2ɑ?��m74�w]��s��3;��z(<��{�-	rE1܂M��A���#OoM廳P�i�`^��w����J�݁��ȡ!?�vh�;��37f��/����ߵ��7hT8��8׍6zyp=8�3	�n��
8�Uص�a���UbK�k�~�sS����/s��{�֤/N�^�qY����YDK+�H[�~�{@$��A˱�9���tFo�D��pC�u<M�fl��flY�'�d%i�o�J�	1A�!!d��d���ғ2O���_v���S��)t)�@����̓������r�/3�]�+;y���sX�Y
KEĽ���ס����۝�_ goM�9�(�0��T4ܐL���v�1r��]���{nr�H��w<u����%�k�*G*D�p	�.j ���@f�:rs�}@g�uP��z5e��G,n�;y�H�N��;���3���dÙ����$�LJwO14z7���Jݚ�/s�]�n�:^�3�e��3T���T@^�u� goo���vH>`�AFfJ⋩0̀R��0��a&bB��H�K���`��������5�p�j`%6������@o�yP��T��\�2��ψ\�n�-��Y�>]�y���38'BA֩շg���w{����0��
D������Akq�z�Fc�d��۷`-N6�%Ц �����*3ӫf��������:��|%*�U	.M����gܪ �����@o�yP�&��"	i@�1/A�d�����`�Ҩ�H�s�2Ig�u����Ȓ]L(�R�n������:h�/s��w��(���_�˻�����UUUUUUJ�������~̬��c[2�t�S[' ��"#�c�;��:�&���4gQ�h��u
��4���zl�-i�z��޺;����x&���rMk#0��>fw�gzȝ�:�&�2�C������|>5�֍bunã���D�.��6��b�[ �q9
XhR���P% F�`�$�&eL@����#_t>�������a����]�{��1:ذ6j�Hto�٘l}�$�S�2��Blٿ��C�4�I��{Sr���Hkz4b=������ ^�z���B���Ф�3�z�pi��P2j��"�|��� ����/~>k�l.�׃�X�F�I���|;(c7;wfU>��4_#q����G=͞�έ[�fnw����#��w=��vOy�L���x�񽽝�{���'�!���WR���t�!i��[A:uUuJ��XD4����V���T,&�0���^���[U�PU0 �-�Z��Ɲ�2�6�\^�=m��!Ϊ
��*�Qn����5�+(f]q�"��n���'�pԫP\m+Xj
��R�k�n���LGTn��"D=�f1Ld��N�-Wg6��DK^�1��[����d��N�%�d�9d�l�2�ƶ��^�uΌ��V㴷d�Y��-����9r����[Rtd�4�m���gX�������ݙ�qW2ԡ��n �wXg�������wEu+<�ڤ%�WGݴʛ&-6`*Vq���p��I�F��n�\g43���]F�U��J4��Nrj�#[3E;m��䜶�4��` #��[A��K+7\ڠ#�]�fŞ�����P�.L���j�/Zv��1˦�U��9��L������=�u��ZRb�[������8��sk�bL�:����q�v�l+�͗�����mv#ocm��ٴ�q��,��ڒ
�;��8�n�2�h ��g���F�:��'Pg�,���"n`z.:t��'���(�hk(V�`�[V������+��ruY`��';�l�Ƙ�焽$rv�1��v�;]��섋[��|'mq-�K,�nJ�����nT^���'��VM4MDݔ�X�t�R1�iD.��n�˰���'%u$�մ�-j���۶Z�k�צ` r)V�6W�	�3��� *��[B/n�5�$ӭ!�^$r�:�t;jv�^�ר��Ź��W�q4��������,���x�	�׮t�Ľs�<�s�RZ8K���E���N{Y����i�:���m�l��I&�n���͌�7F{zM[,W��M�J�4�kC'��{[�����AӦR'm��Q�)6j�mX�#$�٤��$�<j�����kk�`�݊�]������q#+�i��g<uR�ݭ�Q������v���ӯ��N��@8=��O�� �	�UPpC�q=a�����{��N��iV��M6S�������y���ͳ��.٧Ì���X�V�}��^^W���rft�aH^x��;��#����֬��\躧=��>�'Q��-�`��f-��^v�]�V�˝˱�G[�m���Χjۖŷd�X���zl�{o��i3�D�C����s������<Q.�{ru�˚D�I��w=mq�n��46����b�޻��x�c3��c*�\��Ƴ�r���9;7m�7=�q��v5�'z3��7�����L�ԼD��9�z+����@^{���2fd����T��rw؇�瘖�0M�<:�p��A*�;��@{w�(��*>��߇:�������ڠ��;���ޥ@gњ�}�H��m-�P��P�e݁۽Q@N��+���=�� �t"88js�m����*%ߓ6zw^���u���T$�%���J��:x��]��q�	���{�;z�vA`���mw=wW��Qҋ��jhI�d�\���#r;��������\��7Ѽ�۪T�Kw.$��%�w�������J�{z�0y���ј�{q�F��r� ��$���� o�yP5�{��W�{�`n�#����.��q@oњ���Ǡ/=�j�^��T ��^`��8��\�����jI{��В�d�n.�}��T�7�D\����:��x�c��n�o;m��n�;WJWn,z�vzB9O�e��p�j`%6�{;���ި�7ӫ�����#��0��
D�*]���@o�xQ@o�uP������59�LI���.���׺�����J��66JH��]iRq�#4�@�V����b��*=�(�@�0�B����{��>��= >��ۛJ��$�.�ߕ�1�e2&D�pܵA�n�w�ͥ@gљ���n��<�������W.����0�p�l�X��gubs�"3����K�ջ+",m2��F�_���v�E��嶃r^��/qw]���;��a�I�!CI����U�>H��,�������a#���)��]�71Op�n��@g��|���]M@w�y���s�D�2��N%�o��z�����y�y�W�D��꨺｝���K�҅
]�D;�݁��J����@n�Z��w]��x��ljn��Ѳ���n��m��G��G�t\k���1�;�"(�#J�e*�E����$���7h;��@U��{�{��(�ؙ���2be�ڗ6v�(�.�;���Imw�C_��Ͼ,>rX8���D̔{;������9�����B�ϊ�n��19p"I��;��P"�sb����A��ə�����3$��s�T˒�3)݅/2�}ͅ@/g�a@{�n����T�jI��m\┻]��]�l��:��&��\c/cU��n9������]i�q���w7.��P|P��̇iv���k$Eo49�w4�(�8�{=�*t;L��b�㧬�S��n��q���uв�rv�E�nx�g�qr�-�l���R�S�ڤ�a�1f����/SI��5m��:7P�nvݝN�ݮn2Sq�qٰ0�]F�R7��ꒊ�:�?2�g4��g��&,�Ķ�۞{7m�i������Ef^ZTMC�UE�ߺ��������ޚ٫�=s
\��`�2�3��vnm*�sb��zp��$��/j]_�0Ҙ�J_�����<�h�zP��ȍ�}��_�R�6��==�(�zP��]���L��!o@ԧ)�1)�w4��|P��]���J��7^��$�=�d�K��v��t�k�qqj�'N�/Nn!ܶ�q�\U�,�x���m8XW%��;��m%������������O.&���j�;��O(�râ��݁��J���&I��d��3&I)d�6)O��|���(��۰3�\��n��CI��3�ܨ�zP��]�ݽQ@^p�����?�L;��t����PA~��;���==ʀ���L֔�S��,�=�;��(���T۸��/;�&T�.e��NC�Y��zW��cɝ��4�� L:^w./&�HQ2@�D�j
�8ܻ�K���$����D�=(�w]�z6��h�m�@g��P�zU��w��;��(̅���8&&\rԖv���>{�xyl�k���S�L�IQdc�)%�$ �(��U�C<�����Ԗ�O瞒G9���%��R�c��$��n݁��J��7^��̏N�m܄��J��P�n���e@��@^�Ҁ����t��.%��!�ݻZڱ�g[Y5�q���݇oq\ ��n��Jq�Fӄj��������]���$���= �ou����
9���ĵu)�+�S���Bxݪ7z�����$�}��<�.�0��D��wu���=ϊ�^Dt�3���P�)w`Fn�I���@Z�L?����	�qTC�wί3����'���ykx)m��39�@b�L�� 3w��K��wɸ�D�p�R[#C�����v���!�܅�f�.@
H�X�vx�d���˂U���ܘy�v��E���y���e2e'J�@{��vn�TP��Q@j�L��S�J&[P�M�X���������۰=�B*Z��M�Bi��3�ܨ�պ�y�v@n�TTy���4ӆvU6.����v������l���3$�#����ʇx�r%�׶5�LV�U=i �Z8ݮ^R`*y�ƍ<�:r�:]C��xn%�,�xMȈ�sZ�<��vwCg���W�l�Z0Y����Nӟ�-�����s���sumY����/8�Lm��;w]\h�-�����
����{7-סZ_=����r�Z����p���������c��8׳�kz�V�
�M�gY��
`y�`5Z���RJ�M�og<�J���q���3u��u�J�,���g�}�����R�)�� �C\����?����L�-v����yw&�3b?LM(�R�v$�w�"����@j�L_�m�舄���S��p8H<'��������옙Ж{?t]��ߪ(̅��JM8P�\8j寬]Ɂ��������*w�2�$����h��n�国j���y�|ǐ=���:#mu��-�v�X������h]f�	n��og���
��*��-mQ7n�������*V�`z��va�Њc�F�Zv�Io��s5�fn�{���a/��j�&I$�{˟��p�e]CN)X������7n�Fn�������@g�|&kJSS%�=��`f�EE@Ӽ�[��qy��J&�)K�7z��/�z�S^�.۸�D-;�~Ndd���� �܍7O�u��n�\km�����OW3����5��V��춛Is���I/?y��{+j��ި�����Cp�Jlm[�`r��~ݻsz���|P큚�S&Rp�!J�@{3���ߴiQ{|9�֞���kZִ��j�Zֵ�Zֵ�Uo��ٕ����2�H`L'pI�wg@�fd�8dÍ��௑��g��=6�ttt���c���"�������^i,3�:����A 7�u�υ@����͔���0�v!�f��:1Sq��Nk�W��Yy t!7iu�e�it�IṑC�<I@:�A�牳L�uPLUu�HtA	�231u V���>9������1S3�B=*�����#�i�t�Q홐z&P�T�:VI$t��G��<�a��*!H� v�ڀ{ �~�Y��*J������t��q0?{5�I����)��K�wTT�.|P�S��۰23��J��8I�MD��P���1���ۗ`ffҠ?36���2DB���x�Cd,r�ɞ�6���vy��鼻x�n�b׮WjB�tvH�Q���'Ɨ����ٗ`fg*\�2�����f�$k����D�=��v�����T���P�S�=�~&�)�eR%݁��Q@^s�[�4n�`�B>�։C���H��L��o_���.�������At|�4P���x���E�����1�M�	�2������I�����3w�P���X����},9\hl/8+DM�i�{w��vp��[Z;ێ��)��͹�-
hP�ݸD�f�]���QP�=+�L��I�nP�s.�����G�����y_{�v��-PR�/*T��eP|�{j�Ϙ�rd���ͻf�R�/�d���u������۰3w�(	����%^��U; �LJ�T���`f�TP�z��uo�a~�)0
�N�Du �mI��LRP�$1@��\�Ӛ��j_W�S�:�ٛ,���n��ox��k�qٌe�-b:��y��:vl�C)&\;s]��]/lI���=�l�$�8��ձڭؖ7<��:�v6���F�p�m�3XJ��H"�-3��1�4������p�]�1�0l�Y���ݗq<�1�_|珄b*��Rڢ���fKn�y�o*p7�\S��{�kb���Nj�t�h�q��M�o�?|%�N�7V�6c m�R����[��=�2�j�e�ܚ�֙��g�o1v���U�����?��b�L�ͻV|���#��n[s@^sҀ��L�3b��|P���}.p}.Iw-X��0/s6��|P�ڨ
��Tk�<��2$'����$�|����[�<P���9w&_��Ѥ�7���S.����P��T욥���۽���~�o�9��{*qr2dŞ8�kK�S�^��ד��+�:3��;�<길-�'��
p=��=���@��2/�d̛���T��������!�iN])i�}ן�o���L��go]�v~���>��T��P�h܄JR�%�ݛ�`{3iQ�I���v��1�^@�_y��T�Jr$9�.�:#�߮* �O�Tl�U%��ﷴ���>>J*1��iM _��P���ٷ`f����:I��[����Tq�cv�C;�&���c�`ѻJx�o6�ru�f���n+�-i�1���3I�Ao�n��ͥ�32�}��zo�k�<�20����;�ͻ�L�(H������c�Vl��脏ٛ�I�y�C�D�w��f�R�/�ŏG��ȑ#�bf��	M-�ʧf��/3z�A�>��e<�"�qD&�m�^������۰��q@{�d%��2��\�	Ұ7�� o�����fӔ��BI�3T(�bb��lp�nسc��ݵ���:�:�q\c61c�Fǜ����V�#rF7V��{���͛��/Ӻ��сwϧ��1)�P�HOv�6�s2O����z64�G}���Y&N�3�.%;�w��(d�*3gIh?{ٷ`nk�T��ԢSĂ��'��9'Ν���ޫ�̹�tuG�PN�QþV��H�`�2�{���$o�xoN�QGr�X�ٛ�`f�TP�zE�:0���_�c���r����z�*�����{;1��9؞Ѹ-����vO���h�+�p\Jߏ�5��q@nkҀ͝�v�6����E7	�P����cҀ͝�ͻ7z����m5(��!�j�64�3>�]��$��7z���Ҁ��ښ�F�bP�&P�@o�]��n�E~��uAə��ΝNZ-֋yi�0;LC�����T$̻6��3cI�~|��u~��8�2�!+e `�`�R=}��ټ�fl��n�-f!1��&(�Z\���dK��>Bѯx�ؤ�5��9�#�ĳ��a���ɖ�	�ᝬ�+M�=z�O[o�~�������x��칅Ͷ=���y3����3���",�kɬ�v�����v���bp��(��a��+ř`��t����݊Ҧz띻or�vNzs�2q��s��D+��7�gl�u�{:�6�ni�����Ag��Yؗ��N�[q����y��Q�vy�l�W�Nv��|q�g\3+���~��@y�@�����/���*�1?rO.B�y�Dܖ������`F��Eٯ�ٛ�Ӕ�%?�&�T���7w�(�|Q�M�ȝ��	�I8DĻ�7w�(�|P�Sr������N��n( ����u02��v��E��#\91�9P��R� m��]t�q����X��|��c��<��Fn���};�\iT�X����ۻ7z��;6x��:�θ��!��Y����_����3.\���z��� {=�2w3��h��X�ds3-݁�ߪ(��T����a�aKg~P�	p)���P����Ȑ=��۰�fd�wz�>����0�NH��s`�, ��m����7ћ
(ff�n�)x�x�w�Q����+����ݼ�՘�-��m �j[�ح�c��N[R�	q"p��́����7vx�;'ydZ7T�.�ȝ��	�I��w`�,mf��;e����8��B�CJ4@��@w�z o��w�Q�ol 
!A\fL꙾I������]�}��@��GUJ+�US�iwt�/�ݻ�A���r_Ч~T��R��0�$U {����f�;Ӽ��3vX��w��"nZ��rU���DՅs��ɝ��q�6xnf�u�!�;��z��I�tڥw`�à;�ܨ7%�A��m�����	�e-��+�f��,
��˰��5�����<�'�&�;�$}�e�ft��n��>�F��9j\�	�eR�� ���I�~�}�ߚ��M).d�U�GtH��F"dwe�ؔ3v���P�� n�2��v�Ҧ[5���H� �Y^�5�Qױg�=�9yn۞:;N��FT��c%,e+���%�'�=$��dH��Y|�̒����@}�G~z~��W�P�U4������������4��MHjnL)I����s҃{�����<�S���y8s2��50�f]�{w�ޝ�,���=�w yo�?��P�n��N���Ś��/ݷ`���w�ٱ��UNn���X۪�����ە߷_��ι߁�-W	C�`:
>9�XRQ�΃��(lx:�`���t���X�V3��׿>[%[�]��:�5�_l�5,�Ὶ��ȏ���8�E$DI,�('A�z<Q�8�T�lh`�b�E(�4%	B�f!�5Q��3I�AT���A3� b �M4r%فM��BH�^�J�h������:-�$D�'p��Б$F�-�2�b3!b��e�fH�����i�M�娔v��lTF�CJ�	�)��M���bd=��ݖbw���2�������H�"H&+AMPLjA�APE=eEfh����%.v�rCJ6Z����LɁ�F��f�kZ"e`�,�0�vLֱ�Ɖ톯:S�`a���dȰH��mE�|{�G��7����!o�{��cg��;p{��m�X��{B�`��P
9m�@����������v+�j� A�*Ak������m5��4ʖ\��&on�Et�^�\���	���������Y��0����1ױ��e
�ۘ��	�9��8n� �UU{	T&c��k�^l�lT��$�}!��,�A���b���rj�WYˡ��1+g��,gѶx�sWv5nL�7;(��P�p$�κ�Y��$h�Aiڙ$��ȝ��o�,����N3��s�C�$ͱ��%�\�zG*�]e��l.����8d��G	��0���K6C�%uU.��S[��h�6����A=�$�Z�`%W�Px�D�˳�V�ts�7M�=�q�t��-c�]�W���6�;��+��.7NE��3[2��& 6�Kp-�5K�Ks'jm|IQ��t�:�<�1:[��=�J�KF#v[��ʧB�ݹ��>^�l�ƒ�5�rBrI�ڌ�7I�r�F!�Nq���;�[�9ˮ6��Q��������=�Pr���Wg��t�ӸuZM<x��ۍ��� Kc]�`���������N��h9�g��M.v�.F��ͭ�9ueICtD�/[#��X�$�s�DٟF0Ivݞ�n<��9��i�U�n6���χ��a�À���X��$ѝ<4em��:g*Tz�b}*�l�b�!�Z}M\q�vͶ��w��l�o���|�V\�f��TW�4Yj��<]m� X5����>��;���>�6� ���*FM�'a�����-�mm����u���Eg����:�fi_|�7��e�Ybx'<���Ϙ���M�p�a���U�;M}��s�0=[f�vݬ��ty]y��N�X���3r�nHa���GAZ��Q�i��W/*��,�K�\I�p쩺���������$��/��HCtk���u�En^�.�D�WN�6ܮ����͢Gs�)R���b皖:k��q<�������������H�9�0B �� g�8?RA:<��Ch|�P/� y�����mד�ԶD�^��0%�lZ��@����:�-�]����[]5��˞:���5�!q���[u���i�<\�i7(�:q%6^�v�qbh����α���>эk��"���#�"b{*+�gL^��3�p$�S���(d��ツK��"Qق��w[l%�=U�5�l�c��l���m�|}ݢ�H�Ds���m�[����w��`���p�7�3嵃z�<�һ�G���:ۚT�"�x��pgm�+x���Ñ���׀���L ������:�;ʀ�dlLӖ��)'08j��f��ٻ4��@y�ǟ虓3;��آ5;˃̰�P<����h�3^�I$���y@g���F��S1�����*�U"�v݀{{�{�ʓ�2W��3TՁ�:&Ͻ����7��ؠxȌO*�ÖZ��[�xM���zY'S^����u��s�f��[�5�ʣ��9�Q���n����߿o{H7;�~��@F�ML�g���iL֤u�H���K����y�����	s��������>y�{�u��;��k:q~�R��'Q13H��B�02����7;�ZI��|ژO�>��{v1�@����٠���;�@{4:i�R�i'#�&���a���7;�� w�p��g&}�j�JRs��B�Wm��-�.�[�q���"iS����&��DII+nĥ���'*��K���F��@,���I2���b�m��ΩL�)R��S@��{^�����@�{��tfv��ܒfh�L�(�9k��LB)�9.US��u�}�e��sQ!�8�JC�!"B�L�l�d����M������y�"E;.aL)I��s?��s�:�=ʀՙ�@{���p�.Hs$�l� �͚�z{�>�g<�����8{���pZ���n7%M����s��K��n��]2p�'�5`�͟nz��	q���	�>�`j�N �{��sy���u)������qO`k��d�N�{��`��tz{�P~�٤�,���!�����`��@vOr�fĩ/�ޒy�b��IJA�l{ؗ�;�7�P�����$?Z��$��I'ei32^>��W���>��S1
T���u vOr��Kٲ��{:�ټ������u�������h��p��5����n������.�sHG$ړ��&��+��>��i��+ ��`e�6�ټ� ��@n�MY#��m�Y4��{﷿�chY��@vG.z{"@���Tˑ�xw��� �ٳH|��s$�&w=���{:��a8�i�DC�Q334��=�6��������y��Gt@��'�䈛�VK#zX��w �٠7Ѻ��_f����!;��w+�7P��.u����n�cA�!ы�Y;r�5�鉡v�K0���r8�G+	�ݵ�0Cv�ќ�\'i��`J˹ú��q�ƆUO���]�p���L�m:�R���I9�Eɚ�]b�8pk�N�.�y�� �K��c`�m��m�S����tt�; ����0�eU��u��t�{d����mm�Z�vE��m��nz�:�u)�Oo�.�[njG\T�%x�\V�7\���s����wC.��n�p�{�J+h�N+E)�Q�'�K�=����ټ�
�{��3rX��3�'$�,)��7`{6k��'s��@͉��e�d�kc��.�2�J�<LMޝ�4���a�{;}� ��t���>s*�_9*�XoK1%~ݻ �ٳA�&d�?zw���4rb6%D�%D�4o��]�{7�@��T���-w�q�:FQ��x���1�'$�vtuc�Y����\-ó�r�H�	�[��g��͘�̒L�� �o:���t�oK}��`A����T7˅�tzw�������J����3��v >�l�i��f,<( ����b@���v/��=��t������Фn	r���f(�~�grq@w�yP����zh�a)��ln����	�=���嚘���&��0�¤����gOn8懳�]A�G���1���N
ܔd!����۠7�ܪ�E�$����_8��4܍O�O�$�AJ�V@<�8��ٛ�`��@o��P�8�$��$Ă�I����;��s�����"iF
 YO� �z�־��uW=��[\�3��*��:�R9w���}t��&�Ѓ�F�{�;~������0�D̷Azw���AW��~H���K����KmMJQ�B��,��3,'Ԟ���N��l����I<��z�y�q;N]��	E�=���$
�f]�}���2��w�1@f�.�H��jRp�%���v��tzw�ZFL��
����$���؄�������Tg�F^g]�� �HG?	۠3'yP�щ*�λ�������%	B�����~��y���D
�B�UU
�3�}����ݚ��ء33%�߯�㗒Q�,y����l��7mg;����9��yL�n�Ή��:4���fsܝ)�`{w�]�go:�w��=����ݩ����6�&[� ��:Ġů��3�2�W��w�䃻���%�Z��n����h3�,
���������Hb�����̹���`W��unٻ4̙$��wl�S�Y����n%9�1#�9�����`7�h-͊���;��B�`�YC��e����wF�lOS��a��4�n��lR�Q��Q.�v�S��mB�u�_c3�9r��[�-�Ŭ�Ë�:x�)i�l�㭫n7Y&���2y�\�vas7����^�^!�s���.�όz�j�q�+��U��NF+�n���Q+曎F5���;��ufN9v���'d��s�5l;�ţ�uE,��3n1�@M�4��&����}��ͧ*��Kqm�ݝ���w`l�wz��';g9�u��]��p�*	��Ha*Y�#C�-� g�:�w�����sH�q�`oG;�P6�	D6�oM�c�^v݀vw:3�t.�S�bi�C�n��35�X����gs�1{�b����2I��a)L���wu�f�<�:hK��*K|�}�r�XJ�F����m}��t�Κ�� ����_l��·z�!mv4v�Q�=m�s��(-��˗lɃ���-��n5�bj;/W�m��0.��ٕ@��@v�w$k"ޣ]��뺾|�f���~�2J�*PO��y�w��}�|����%��~p��`��y��'�n��\�H=��~� ��΀��t{a����RC[��#�r�����1vt��8`z�������� i�t/wM�ͨt����ۼ�8��)�&eÆ��C�����my����v���e���Ǚs�>�nz���?K���N��V�`U���gs�����'
`'S)�)Nb��ou�gs�1{zhzp`{��jK"\�1(C�v��� Ź�h��_��UT�۫�kR�n��kN�n���������HXR�I�P�d�'�M��sy�&���
��c�7�v�HQE5t�Z��(�m
�����N�p(	��7�:�;	�w�4�4L�QUBP]�`����7�f����5�S�S��	�;�2�i�k��W}�,ٛ���͗��H�P�!kJ���J��6a�.�J�Ҕ�Iu�E+��T9��vi�M��Ȧ'y��c@w���jD~K�J��쭙R��fR�4@i$7&��'H�Ol�'zqԉA�%wD&�΢n�}"P�0�'{�M���fB��t]�����ȥ�D2��v���c������l��`z��$6����B�&F���G����;A_��C���rX��{�� ş/�G4���n]����g���T�H}�ʰ�����@vj�
^\D@��f,z0p{7n�;;��s�����7�M!YM�W'[v�Yٗ�p3�]S�7l�Lt�����,R7���O�2P��v�ݚϞ��2J�=��@���4JS��� �[�����^Κޜ�ۿʥ~�/�(��	L�4۠-v��ޜ�g�v@�΀��h�*O�Ĕ��T��j`W�7�����s}W��Ύk�:X�A+H�82:q0KBI0F�cJ��|t@�H ƺ����V��?��*��&�2�(�mI@{���`Aۻ4����G��ZK�9l��4��8�n�����G;�)�zM�<l�ܧCXi�\u��Qs�UWg���?����{�l��Bz<s58��v݁��v���;��)-�m���M~c��� }�� ��S@{q��K�)����������ݻ ��t-��`-�'���̐J���2ooz�?~�΀Ź�h����z:tI�	��H)n�;���s����ĵ���{K��L���f��?]�����Q�Rg1U�Q�7m�N�v��/DY����q�}�ݻ�fګB�{^�n�E�(�l`�^ ���y2tL�]V��u�uJ�e� ,P<=�vR);=�6��vz磜mV�8�9k������*��Qi�<�P9x��W�k��-�ǜL�F��6@Muͺl�	���5a��YiI�G ��Woo $F�Hrgz5�=<�d���=�+�M�D%ʓ�!r�cu;1Z���Kbx��h�t�+����;�m\���״�������4{0+��M����X��t�R�̟S �U6����f��v�1nM}�F�q2�D��(o~�vݼ�^ޚ=80=���8m�L�~C�v�v�t/oM~�AW��`bߗ�҇3*"e�3@y�͊�%��(�;n�?v���2D�)��ʘ���.}x*zt����Ynݸ4����^T��GӗsDӦ���:0*�v��y�A��ĪA{�m
Id��&\�%~{�w���x	�
L�	�K>�}�����^��}�=80+ޏӢM@L7 9%Jn��y����V��88�3��
�ȋCr�J�n�ՙ�A�<* ���v��*��f��%l����ұ��:3��ou�{����夗�0y}'�1��mU�H����'�ݞ��q�����u��8f��M�������qr힤Q(M�x����� ��tzw���!��gݪ\1)nT�݀wo: ���@g���;n�-�}��(s-D�"&f��њ���52mC2B$����|@A��u����U��o�;67���h�bIWMX�:1�W��`�ΰ@�;ʀ��6�$�RM�)@�P�n݁�3$���`c�z(A��xb�8r��К��|2D�͖ݗf�7*�ݓ;O�F�; Hx�v�n(�^�R�� wo:%B���31�@_�;�����AQ)�PA*[�1{zb��c�{��ݼ�1f�<LT�sBL��S��75���۲R;��@����@f'
`'\�)L��(��n�7sf�>f��$��ffa�aD	Q� ��T6�xT���������R۽����t^Ot�y8033:�L�G94��hz�v��sk����[����{q)�.�u���x��&xj�m������l_��=��v���@���H�L9 ��&���^ǥ^���f�;��'�����}�}��Fݪ+�H=$�������tz{�~��B�IK�&!��@x���:~��z9s�������vth��*	m��R�ޝ�@_�_�n� Y���G� ����}�������j��$͋�жm��c����6�.1'�յ�ђ0���͏FP�Tlms�ܘp�/(�Vyr�˧s��z%6^�	�j���gg�k��y����O @T=<;G��f�<c]V�gmH��EhNɋt����Q��	�p��-+��͍��{4�'Wk;��Й��ػbu��Y�n6��k�ݛkF:�bQoY�ֳ0��� �l!������H���QXۤG�˽u�lm�ˮݮ��v�.Zgnmu����g�M��hO���;'�������o:�;ʀ�bBs))��%"e��� ��tzw�~�Aw�T�#Jf�Kw`�΀���P������5f�}�؇2�ʁKtJ]���=��������@_�t�8S#�bbH�uJ��l�ϼ�)�}�K}��&d���Q3*f�jY۞��I1���u�Y�pkǑc�����훲s�l�
X��A0�!�����__f��v-�������Y�$��\��J]=���:�4	��� ��� {�'�GWB���&�L�:P�����g��p�ٟ��z5#�#�a���@ԧQط����~ί��z����L4��I5 Ԫ�Q��q���Q�՜��#6eL)�ĉ�$�:�}��{����o/�۔�{��D�N��!2���Ɯv�mՎ�&��\I`t7�A�����y�;j�^(D�_{����g��ێ2��_^����l�$UȘܯG���g7�ӻ�~�G>��k9��D_'"�D�z��w�\���h�3����Px��� ����Y������||�R�P�Yb�[����s�}������qɞ�.ԓ��@�
]DgguGb�__�g��TG��2(_���-�mZ�{%�86.ǉs`v�5s�C�F�q)M͒�
"��hE!lhU˳߾��o��9�����{ﵜ�x�߬$z�ɭ$�w�S��}����磿{����$Q�:&F'	�Q����;{����l���s��&eӢTK����̑���lΎ,F{ҳ�F�&��-���g��6��a��:�P)qQ����{���3���̍�͒�g��P��ݧ�;����9�{Q���j����Y�EU�!""����B*���}�S{���ۛ���kY�%�y�i)�D��eɈ�_}��̓3;{�FgO�}�K�b~ԓPK��6I2�������"�1��gS^�w5�����/2W�&d�Gu'��*���7^�|ڶ���""��1I{��P�䗽��7��C�%/������?�QU��� _���a��E@�[�ZQF$P����  ����kZҁ"��Ԋ 8 H���Y�+@2(`�"
� �2 2� ��vJ#�P � �E�UTABi@	@D��i@�����AD �"	Q �DLh�T� fPF!%UJ^�D	Q{;$�5�"j������@� ���5�������Q?Ԫ)��A��U?�"������?��"*�J*�J*�J*�H��"����R*)b�����������������������������������������������*��"�"�"�"�b�"�"�������*�������������*�����h��(��(��:O�J��QH�� ���?������_�������?��? {���_��A�U�����5�����TD���������������G� (���?�?�� �Gn �����?�C��� �� �~���3���}�#��P�U_���=���n��O_���w�=?��[�ߍg����_��I��g��C��Z������/���\PAaHBDR ��FHA �Q`�FTID%D��   �D�TJI�RaD�H	&H �R%D�TID�R�EFAITIBTIRTH�R!D�Q&H`��TH	!BTIQ %D�P�RPRIHX@)
B$(	$"%$��d!Q! A		D ��	d IITIT$!RBA !  		BBFBBBBBd$�%�&!"B$ ��! 	������@���Y��
�)��& 
 ��iB������@�YH		UBP$ XId	��
@�I��	��H!��
P�f�%�� ��� IT!IBP �%a!T�$��IU��BU!!���%`!I��	$HQe	@ITXBQ ���! a$��RBEIH	T� RP�	I�B@ $�P�BB��$A		BEIA �$THB ITa	��B H�dHD�$B�%I�IBB�����?��� ��"J�$���! B0���$0�J""�!(R�"P���@2� �	 @�B�H(B @��@����*H������0����
$!�!��(B���,!#@�02�$(Є0,�(�	0�$J2��I�(@�	! !*�� � @�H���H�$J�
"���o����'��w�=i�� 
҂!3������G��ҁ�E�����D���֎���l�~x�O�C���U���?�*"
��g���@ ��_���w�����U�j�����'���* ���y��u�AW�~�GG��+�{�?�PD3r"���?���5�p�����=�<TDl��W����eDAW��> ������: �����DAW��������?Ġ�_�����M����?��_�{?��6-�������g(G��h`L��j�����|*5�O�֝	�g�͈�A ����<�?���� Q_�����A���]�|Dr���O����a�?ÿ3�
�2�ϢN�@,"�����9�>���  ��/�  ��2 (Q'@ 
�  � � ���R��JT(�@ TJAQ	E ��TI"�R�E(P
H�QD����T(QR(B�!P�   Ā�U *� Q1�
x&�����_{� =���oT�z�qs�qk����U�}��5� �^-�bﳪ{�zs�2��]�>^����Wζ���>z�����x��W&���Ӏ �  �@ "�M
Q E }1 � C� �D
 � f �� �� 9� b H�@  �A� �k �� f   )� @
� ;;� �� �      Ef`���{��KŧMqis}���Mo= ���>�v�6��;�{���u� >�s������R�k� Z����w��������/������W��z_3���>��+�qs�޽�Ϻ�Ϋ���z�|    (� �B�� h���y����k�۶�<�=n Ft��geqgɸ�:�YJ�����v.\Y� ��MS�� ���]5���f��t��͗��>���K��mqe���i�q�:��  P  U QX� s�����=�z��I95N� WNMS����ם�f�up �=�,^p��� g6�������{�J�w}���u�^�ܯ6�޴� :S��� d�     OPSm*R�  EO�CSeJ�   <z�RD�F Ob�PiJ� h?�%3ԩJ@  �h�ʔ� ��w�������������I���G��w���
�B�� *�(����� *��@U�AU�������K����!O��M��9��'�"]&;x��l�f;
ͱ��s���~`FIMF��Ħl��ۻ��5������o���,�j jYϮ~?� U�`VD�t�?g	�i�B_�=�I�K3� ~�Hj���0$>�l��K���O��
i�f���ofB���&%:���X�C�����Ygvt�)~���~g΂,��F"GP:#��N�Yut�>`R@4X�t&��5D�X_��&}?[�2�` ����b��������4`m8q�@�4a��<(~�M4�|�p�Hd�DӉ���l.׌.���{�`K��P�!O���No�a��!n@�
I�+��I,�7�ۗ_Z�����HBCC!��!D��-K�J���UyU��o��٠�~bȡMX�D�@�E�k�ջ3����,�B�~�|	$!@�n|z�5)+�*I����^���f��>�#MHb!J��(U��5�D$B%YW�j0����z�.��rg&c�9�utI)(K�R��wI�����]�i�����Bg��~?qSp0!��*B��, ��,!�����c�ё��ԁR�D����!�aR��`P�%�q�ϋp��{v:8v�r�����%��Ժ���d�tZJ�Kk��B�R����-�&��~���y H!�$d��0�F��$X��
P F!bP��B��HE�!!FF*�d���5$���!�i���b�!�Ͼ~�皺��x���xr���&di��jz}�p��֦�Nf,cg�����K��������ݎ�z%cbH�3Y��	u����݁J2�Ժ+��4�k��7Fl��CG�P�feu�s��j��]��ƻgՅ)B�������O��  � A60��H�$
s���g'!C�)��`@�
!4䡁�!����l�������#M@&�b���tH���or�����#t�/BP�41 ��aϾ���%.�Yw��hv�{�ȩ*~S�1Wk��p�N/H3|�4
:>&��.�)�h�~�2� �� E�!VaX�
ju.o��1iI)�9�k{'�$c���6n7X�!]$i��cL�3F�o�f`��$Jm5��%8sG	�����~���0588�EF��|��F�����2���L9͌���u���	�	�;4CZ	`]��˭���D˗g!y)�u7�a֖�������+Ư/b-	R��)Jy0bF j~p��LF@H�au���7����s
�h�4D*�&���I�ˆ�e7�a��{�b�c(ٔ5�Z5yX��[�իT�JՉ�L�����z)eΗXU�yVU�.�wJ��[�u��Y����7���}��Q�E�i�Ѕ#YP 0wi��a�j�?s3>�s���8��B��4f�����n͜��?i�4~uU�.�bB�3۟ʒ!(!Q4҄�+%��ߤ�^{�Q�ą* P�*:\v�ǁ��t�m�p�®�6l�o�����4r]�\�7�	 M��č?�xs�%�i;��oz��fo��SZ���L���P�D޸��#j��dUY^�)y!8� I	
���2R1���FHIR-1#4R�Sc��7���!"@��B��B�{�����u�4�~�$�5��F���X�X%%��,+�6���Ek�RM
ĠiL�s�����6��ԃ]��c��Ѿ~B�$��Ʀ�1� R4C&��th�\�QaHFY5���c���FoF?sA#d!Oپg6)�����˓�"D�!~�p.�ؐ����H+��8!M^e�{�8o��F�!BĀ�!(�l)CBXMkn:6}��-��ɹ)5��a�SC�B��hM�A�?h�r0�3Xo��;�v�Y��Ǐ�I��k��CB�B1z	)H���(^Ċ�/��C�8R�~1�H���>�.��1�c�D��)�02A2Aat��J�+;޷\?@�
|�$���H��%T*����5yQ?g�g���~Jr�������
j�"o YyTQ��j��Q$&�}>e�&���l�MJA&f��f����7�ws!�>_�ۯ��p��뫃��q��N��af�]C�0aXY!H�!H2@�HЎ��E�b��
���ptmx�̺�~+į���	WJ���~��.�k7��;l��u`�|��]k0�g4� B5��?�z��'6[�?�!���k�?~7�SXc��0%��ԁMo��0�k7�ߡ�B#R!||P!da����5�������BV������3��!MZϗ�!MZ��˼�~�������n~9��9~�FcXXX�]\��~�����gۚћa��r�B,(Ƅ���^7W�Vϥ��`V	]4˽}���o9��/�T��5L��?|$�Flt���H��j��̩�c������!5��D�!! ���Ddb5B�~?~�0 P�F	V A��āB:0��Ƅ�Xl�	�����J]�O�ĂPӈI
H��'u�P1:�#~�m���$"��A���%�쌉
Ɛ�D#,a!J���&�}j)z}�}�z�Ǖ,��\�6@� c bF�����H$R�ϗ�I\U�<$/|/-��d�B�R�l�H�j���>c��@��l�~Yu����٫���ύ���E�����#�7�N$h��p���?'�␒˽�9:�\qb�"@�!����B�1 GdX��$!�6��X�H0!��D��1i�6#4ua	
�0�f3A:C��MhS�.�GֽU1U��U���^��CN1 �ֿ~�M��H�R�h1�9�]dְ����'+�]j;�|14�k�N�`�%6�F3�Ym5!�Ԥ������O�};��!�.�.�0�'~?N:� �9�ۣY.�M&�]a,^�o�0�����`Px�H�4c� F�0�`��3fmNI)u�xq�;�5�dg$)K�
�@�`B��4ĳXnI��L Q���ݚ�SL�Ѡ�_�u~Mg��6t�R~4u�s�o��
h�b�ћ8p&��Y����i`��i��E��O�?f���������h�|���|��h*0^�DS&��"���հ�*ZJ#uP5g�a��;�>�.t��!]0����V6p?@��	I#X�T&'�F��}�����;8��#��B����BK��rN8��0l���|4ћ8"J�K
Ku�f��� ���Ǚ��R��iǋM��ܺӛ;�1޵��77��?J��p���
B��l�<� �l��R!z�*A��9F��WY��k�8FL�[�˾��:	���G�60�r�D� �Ur�3¡LJB=�9�ٯQ7T��.� �$,
�aI�f�?���!M������hea�n�$��ψ}�|˨~��?,B,!���"�.���]$,�KԤ�l,�ZL4GF�U�!M1�(M\�cû��Gd��֪�,/�Q�O�� �9
	��++}])-��n]�u�^����\��2��&�XI���c+����}��E�?���5�HV�1ΝM%v221�Ý��1^�`hx��%!B��H��y�'5GN@���	%�	-#]�8��MM�o�(K.�)H[�g�5�����ґ�c)��l��A�6l����}�d�����&�!�D5��.�����������;N�d�]ރ��I����O�>�ͬ$R���#a$��ep�SA�(@�k(h��Fʐ��LRHP�Fl�ԔiH@�cԗF�1�X���
D�JQ�V^}�n���Ŧ��dK(B���k���P�:j@�B�2ĥ t!B,&@��ٝ�p��0۴�t	�0��f��(��d#É�773X��ߚ62������o���rU�H���m���~�,U��e!,�u��!0R]B�kXInk��ߥ�N6Cg�Di��7��|�M�.�~#���p�?B�`č!v���hБ��r�$�u�p���JQ)%��B�$�տ�����.�F%ؒ����k2S��|�8�
�1+
���h#��B1�l���M��f6���S%%��g���7)�����I&�FƬV2�3>?h��
h��d Q��.ptLSdJr]`J��3c
i�m�ٛ��6-!M1�JB�͚��$�"�J�i@UbDlh�1�\�Z,��+e�����7�&~dټ��r�9�p�&�˭6�pə���+,7ot^���N�{�y��~�  8  ��  �g   �`     p    $� p      	e  ?�|    m -��          ]�r�I3���Y�8r�v	�ݥ��������h� ���$�l  6ۜ;m�g���u�ҵ6�aWEPn���ݕ�Ѱ/����kH�A�A ��v0h!U*���� �jU�XZq�V�mHR�U s�[wm� 	6�UUlu�6:$M2�l %K6m�p$N�l�kX8we�۵�� m�$6� Ӎ�6��U�wKX�Tq)[E� �G�i�6S\�mx)��m�m��R����Yn��e��HWKʨl[*i���m�/	���s<m���e�\��OWl�Z�@��:�74y�����!�O �+<Hz�[��\;n� ���j���� � $�`)VUBju�9v�����P�%��ܠ5մ6�h��Z�`Жku�J�]*�h9��U[�qS��l kbro]m6�h(���m�M� 6�]����m�v�lݑ����� ���|s�O����U�Pte�U���`7m�$m�ƻfݻ	���m�t��`mv� � �A�-�)�y$44�[WWTl�a0
�YU@�%��U4��mR���ŵo]�Ͱ8D��j��	�(��>�|�Sv�td�4*�@P ��I�ښl�}���m���ж�I��۲@�� �KM� E�m�d��.̷\�q4� ��m����J���g���( $H�m�tZܸ�f�6Iz��K(n��kX6Z�8ݶ6���m����ڶ$6��H� 5V	�\m��  I���հ����:��`��&�0�`��z�B@t@R��F{@��ݵMe�ۦ�ӝ�ڥ��xT.�A�S; �mWR�F��jyP��UΜ�J�C����.����"Z��"xvY%(,�s�� �E�:����p=�Ѷ�n����g=Iö���������r�����s(�PQ.8��]�"�I���g �Qm�� ��Ѷ��i�j�*���Xh)9�yM��5�@T��pI��l���m��m�٪��&U���{p7d����vJ�d ۈ'j�֠��
�[�a<˔Uiv@6:ۥ�	Vغ��H܀�X��$�K-���7��Kn�p�Kbt�iH �E;&�9dA��A�J��=�
�� ��&��6��iH��m]br �EU!����UQ��L��������ҙ)�,C���hX�# �I��{��[V�X$ m>�I�I7E"���e75me��*�૥ZS���&�ݪtU*�UT�@v0��<�ʫ���|>����^��K��F��z��h����H�.+��Mjj���u:Um���-�	�Uvy�ڶ��UW*���8�%y,5�mY�ie� H $:� 嵶܉�t���)vv��Z�V��l�Z@�Ic�rԓn�^��@sr�T��*�on��A�{�ZDT�͵\sm�m������k���@��u� 99��b�V�瀨3�eZ
[��6�D�����m��6�r[��knl 4P	 �ݛn&EK�mv�uK����$s�;i��Hm�[d�^-�kh�psm�v������ 	m� 	�H6�/]�*Yv -����    ��    �H   	e�6���[hI�Ž@�H��[n��ЖT*��8$�� H�v�� %��p��� mm�si�� j]�
������)�ۦ� �`�URZ嫩V��˄^j����v�ěJ�T��mT��  �$l��"����ﵻm�ku�k�&żrKV��ٶ��p :N H[A%���C���u� �i��$n�\Fx�m/=������?[���n��s�nΖX�(;znKn�g�ZG�s�z�2q�Gd��GQ��+,�*�H�lcu(g+ma#.v�v��a:��.y�O�t�8�n��t hP#&v�u��Ԕ�� $l|9��4�YjBk�C^6$�-���p����  � [D���*�B7���us�v�eT��UWl�05�$�j�ky���Cwm�� l�K�� ��C��:�Y�.J�j�6綥T��z���kմ��gP��n��@�� �UG��BP����en�PZ���m"m��m���ۀ֭]Sz� ֣H��Uy�&Ce�q���z�ۨ	 m�m[��Ҷ�sn�
��j�S��+8��C�$ �  ���i;H�   ��N��;�&�X�V�A��@5�zk9{B�-cm��%H���e	 ��޼�5����W-vF H�t�8 s#�$� ����(��qȍr�U�^m��$I��N����V� 6�ñ���c�C5kp[rr�m��:lr�]�F�U�KUuJJ@�'YBĺ���m�Kmm�h>9σm�8jY%�Z��gDmZ,�8)\ં�2~����v���n�U�e��t��))��UZtvi�[pw^^���ut�6�րpJ����l��U*�[7`#���D�T�\�q@@��jh+u�p �<��qv8���5W \�a�mJ�@*׫I������m�( ��U�Q���m�ul��azА   l�	�v�i����,#��D��`�����PV�����T�Ka�[\d[Nm&� ���� ��.�$�Z�t���� 	m�"Z 6��!�U[Ug�U��q�cC��T�K���I��i;n7F��-�m��(m� �  �`�j���$ ��NHV���h E�� �kn�c8�l�Ā	�n�Pm�  (U��VQ�怩x��vJȻl6����CbD�$���   [@   �o�  ,1�� � �l�D	�lR%qUuQ�p ڑ#m���p�m�gm6�H�����l�`3���%� p�6�2��UR�sT��K*�V	T	V
Z� ���� $E�������N[�:ޒ�%���`�_�}��[T�v��U�ej���b@6�5�vڧlpD'	l5UUF�M$`�@v�FU���J�V��
ҷ+P��*
5A6ҝ*��WUT�*׭-�z�V�m�[A�E�B�`�孻\��vMɛ��⺑�}d�t��rkR�0_}�}}ڣ�2<��Zٴ�	g�   &�i	Hu+5Ҭn+����Td��Uf��UZ��n��Y�)'�3a��;9���6^�$�Ӫ+MH����ܐm�P�E�����X�G�	V���Z�����X*v�ly4�P�` ���u��l�O�J��	��
�X���YX�T�-� �i��ų�R!�q:MY����lz^r){:bYv�6ӳ@v�֊-�Sg\�T��w�UH)�J�*���R�p���*��[�dܑ�m$�jh�ޣm���	$�]v �H�I6  2	,
�++V�UWp6U^��4���i��-��-T����b���K����[%n��v��[@��]ol,5�p  YVӀ.�F�    ��y���\�W- Rt�e��i����UV\u��9Wm�h�m׳m���6��9�+�BC:d��,�6�d��-�KͪM�p9�3�� �H�C�֭�f5�6Uj�	��]5+� [WSe�W��a�8K8타 6�[p	8� Er�l�R[@$d�f��tڭ$��C��Sͱ�Z��[��~�'��ig;m�� [@ l�lm��@�-�d�6�[t�	/T����v^@yV�V�g� �m�$ۤ���T 5����.T8��U�:�eY�TpQ��� 6�����m�t ��m��V��  Ȑk��I����v�j55���ʵ�I �sm������[os�vi6?A���  �m��Cm�m�V�+`� ݶ *��t�m�n�ʶ����M�Ä���*AR m���`�ֹ!;k$�����f�  @p�  9!   � 8�U�@y���U6��#"�]�`A    �v:Cg���lH  2v�]'2gJu� p @   ��� w��ܡ·�UU�J�gjg����dȒ��ZM��⍺8(�	P*����YZ�>�/,�d{i+T۵Mr�m   	7E  ܍�M����۳`��A���|6;*�r�n�sZ�UV�2+�89��BU��bRZ�� �gϗ ��I�2q;*�j6z��1p�<��7I�[Rԁ6.uMGs��PJ�T �`  �����k��     ����[��    p			            ��ͶI���8�v� ��     v�  !m�f�[Rp  k����H �����������QAM���@?қ ��<������ �S8(�����@ � ?���t&#Q:i"��0�0��"�P���	�ںj�� ~ �!�MhA�"�Ep@�; b0�Q � �O� ��? �"0@4W������P���=E�*���/C� 1��U�c^���P�D��H=LQ�S��v~S`�� 	����OȇB�(�~(�� ��� �E��v�� T�N, �
�z��@M�PD�@&��A:�$@~� |�@Z?�IG�^X��>7 �b(tQz)�T #X�S�R�>B� ��I"DdB)J��bR RB+,V2҄�J!*A
)&���Dy�N��@��EdV!A�M���
���E$���hJ*�h�"������U��أ� 8.�~Q���	`��! ������ ��O�������p�P�8R$V$_ˀ��� j)�@
��QP��Ѥ:��?#�|��� *�Q�'��< $�Ѐ�H�
A-J�Z@@@�EQ�3�;�ֵ�ֵjݶZ@2$ Xm�kj@�`��GL�-m���X���Y�!i.}z��l�h�ڳ�����l��V ��^��;�ڝ�=7qOI.�tꎷ�&��*[Ѯ��+2٬�eUj��9XA�eͱ��<�pCg��G��FqɊ{HZì	
eSa�ㄣ%n5U��l��r�Ө�5��4s�D+Wl���p�m�c��n�b�h8�J�Vz��ݳu�����x�go_M��� �F����cp;�ۣAr0�e�nV����ѺAr]��c�i�;9��Hp�=���ы�Ԗ{:���)�k���6�5� �d�������x-J���dk���WD�:t�t�I"f�#���Kg\Bmұ��89�U^��:�_5��l��[XƯN֓�v����:r�1�-J�U���)�ð����`�n*P�S-�0�;s=Jd��t���z��	�U,`u�
Q=5��tKN��l{�pƞ6֙���j�1]��Ѵ�Z۳cJ���U8_8��(u�ؐ�R�ˠ�-����;ID=jh]�*l�:.�l��"NWK�/[-oH䪭��.J�]�1��%Um��c�6�h�ts%����/=Wg���6�P9j�V��|;��/(�d�8�j�6ĺn4Z6��������\�`@�+�-�MeX6l��gn^stNr��)�Dz�;Yҧ\M���նy���jYk�Cn�,�=�wAi��[�Ɂ�Mb�:�۝��vs2��' �Z6-cs�l�%��^�b�C��R��kl�/:��
�D╠��+I&ɤ+v���Қ��;Tr�&�X�p���:r��h)�5g���� w7g�-�,H<=.6���ړ3UJ���a�,�zf%�L㲲�\����6Գ���텙��#6��u :7k;`�y]ua�6G��볤�^e �
Fw;fZT�l	<�'	w<Z- �msPn�$ ��;U�m�cvt06���}��� �?� s��UD �+�P?����)����Wj�q�
uG뜓Z�sV�3Z���L��7 �[Eq#�R�U����n7V�z���wU�`ۛ�.�#rs�G��v��m��y +v���"�Y�x��x�+T)m,�qy)��wj$���q.��۞`�j�/'V]�A�gA� ��/n�:测\3��.�Jj���n��6sr�k�#��5��pO#��f�p���h�vC�i많��]ܲf�f�����J7{���c��e�/n��x;l�<;�9���=����Ww���Ě�Ƃ%]���Iqvb�$�9�����߳3�i/;�ԒW��O��j<����I�ܚ�Iw�ϾI*��RIq�_�$�s��k���,ds&��]��J��cԒ\v���$[w&����E󍑌I�mr}�I+acԒ\v���$[w&��]��K��=���q%�d�RIq�_�$�mܚ�Iw�ϾI*�+z�K���fg|j��50X8a_��c�(`����+h��N��K��X�д�ѹ�.�l���
&�q�${�ܚ�Iw�ϾI*�+z�K����$�j�-	 7��brd�m����8t:`?�:!BA[V
�[`$VT��� Mi`���$@�,d ՕH�TӥI�qZ��@�#�([s[��kv�y����m��w�RI\�h�ǍL�xԎO�I*�+z�K����{��m���&��V���H�{��qcxۉ��ޤ�㽯�H��MI$��g�$�v�I%�t���ƣɑ��$�mܚ�Iw�ϾI*�+z�K����I/fff~����I�j�[m�g��Od^-��r��u�r56�ݓ���ΓQk���{9�v9�#���BI+�z}�IWa[Ԓ\w���I�ɩ$�:Q/�DcsA�|�U�V�$��|�E�ܚ�Iw�Ͼ����k��������doRIu����J���3v�_� 1E�fe��O�I*�+z�K���2)��ƒ�?�I"۹5$��-�|�U�V�$��|�\��K��1���5$��-�|�U�V�$��|�E�rj �;�}�6i�+/�#s�c�VGf���&���#�Y��n��XF�����K��<jG'�$�v�I%�{_�$�mܚ�Iw�ϾI#(;A�m�ӄdORB㽯�H��MI$��g�$�v�I%�t���6��q����J�7I$��g�/f6��7�$��|��$����X,�N8�$�jI%�[>�[{��m�����9m�|�1b(� +�|"��é���7m��x�Ѩ�bR4��O�I*�+z�K����I+l�5$��-�|�K�*�[2Ƈ�v�q닃�m�N�MH�����^:u�t
N�c�s���,�`�ݴ�~ \|���I[f�$�9l����4����@���Й��H0�������&�<�\�_I�1ʻ�F���������@y么_I�ܦ�r�+�X��<q��#�Cً�z��[��@6���@L �6�i�QG�|�k�=����������>�r� �J�"T)�*�P"A���H�@�#�{�|	�ww7�����Z��aIG`�ۆ��׷F���6쥮����Z|�3m�s�@Vk(%���B��;�r�q뫰kn�5�O#��jZ�����:�q&�������Z5�IJO���67l�����F��^����� Jԡ\��I�:vWm=�K��ڮވ��;���g�무S.�G�Sl�oN���G��>�r��nz��1ӳz���<u7�K�]���T��^wGglj�������k;�ҹR�oJf����r�=v��瀒o� �Py.b���p�Q�?ɧ$XC@>��~�����@��@�{)�^R��2�w/wwPy.b����� }�f���Tm�"LP!�6�����@����hu�^�W-"�ӐmI��vS@>���:��6w]`�-U�\I*�ʻ�6�S�·�ts�&Kv�=Op�m�cnۊ0�t���ƹ��"�1<
G�9�zhq�^�{��(_H=w�����*��iL�MZ�f�����|�PX�k�LP\$@B� t@�����}4_Jhܶh}�4�"�y�������;���@�5�ʫ�..�����n<��$��fff\q| }�vK��;��q/`��'"XE!�r٠{?~�vyy���M�즁y�A\2G"�~ˌ��DV���#�!c��3؇����l���F�������irM�X��s�h�e4�[4gKab�a�.jnp��yВ���0��x�v��*�n4�QLi�&�ܓ@�;)��5߿~̾�r�rj��(�L��#��}�f��,Uh9�4�/r���NbsȰ�ɠ{�\���=� �I�_��sn�=yW��:�r�=N�;k��y�	Š��y��,�G��n����y"~�w9��`�=�jݒ� %_)�������jJ��}���IBS!���]=X�k����7N��L�	'"X5!��4��@9�٠w���9�T�ܑ���b�9&���X�k�}��ix��$
&E䦖'	B��u� kú�L�-M�[�{���@}_ ��ڀ�d��������{p�Օ^�ǯsk�7b��聍o	�q�`�Ү��c�{lk��xt\�a�37u ���M@{�\���>ZkB0��jid�՘����
��_؀�j�� ::��ʻͤ�9�a�@������y�M ��� ��q�#X�6�i�QG��5 ���M@�M@J�$0ō��qc�9&��vS@>�@>�;��O߾�nI�1> �U��d����nӧ3fj$7���<K���S>�xvR�;y]��cQYn !����ʶ��z�֬t��밂�6T�v�֫�I��7]m,�FL��߻��j�7g�]�-���ctm�qڻcc]���]����9�s�Xq��e�Oc��iu6�9v��R�I��=5�Ls˽F4�]n�q��v[1G�-���H:7�4d��vn	��
w������i�u۞ݨ�YF�����4�
����ۃu�3��;t���%d�πh;%o�������	���@>{t%���Ӓ1��@9ʬ�9��h�e4�[4gGSYI	�#�QH��{�@�5 wK����	Ħ$�F�ܐ�;��hܶht���@z��WB6���(/n������Q>�:�u��m��������ݼ�t�6����G���r���jc��`�N��.�{v۠ݮ�灌�J�Uw�y��{m��m�
�;�M ��{qoq��M��vn�%��� %l:�֪����� >sP�P��
����ͺ�ٻ��� t��=�^�;�)�}���HI��K�4�[�K�s� {t%���Ӓ1��@9�\�9��h�e4�7xDD(�O���55T��S���e��%�b[ӥ�3�J�ǱO ��Ghh�� ِ�&(F�8���;�<h�e4�[4����jlN
`���.���7�l�P�C��x��׀{v٠}�기�)�� �p��lГ������{gA�C�8�q�s< \0�~n����ep�X�XK �6+�"1"{�]�I��+��h�>3Z(&�L�i���>�U�_T}�Z����`yd ~�2��^�j�!�,!���~��F#Lh�J�O�}����h�]����7G^>��W���wd�(��� :�C���`��)1JŌF?�b�㮜q%`fb�c�h3��Ƹ�;HPh-{+,'Gd>��^��)!$Bm�}�Б���^DI��g�l���iur	���Q~�S��G�
b�?l$"� �@z|�=�6�D9Sh��V!�S��~0�ـk��qR����M��y��;��@6��`���k�ޚӾ�4� �6�MH���`�m����;��@}UWį���{N�2]�Z,:�5��U�KjZ��t�n��3uX($:ugnTFc�UI��M@�f�_�`�߄g|O!'�C�,���l�rڼ۶�wm��!L�{�*j��
���ܣswP}������ {���ѕ�I	�#�!&��.۾0��������
��(�"%O�Q�%�(�}���?�TM\��ի�����}���P�ou|�� �H�q7��LrF82F�4,ۧ�c���������xYu�^�rGD����_��S&'�H��/�4�R��짳>A{g��瞱�R$�)�	Uw�y��L���=w� }��v~H:w�ƜDbp#ME&��g�}��9D���x�]t�O���m9"��Ib���@9}�s�:�=�m�s�'����!ȖHh������ ��W����/���}m�^n^k��X�MGmxڭG
��y�tq����sŭt�6̜�bys����GQ�y<v4c�iݵ�g=�ջu�
����o��t����T&�ӑ�Z���Ӟ������su�v\��n��/Dbk�"+K%+m���m�mZ���-Ū�ͱ��6�m�wP<t�n���x�D���!�����t�#��5�s.��n�k5���� Xu�N��������[ю�;�O�}��<�d��:v���=��i��k�����v���U�6T�ٶ�Q���w���@����;��h��3�X�Q�a"o�$qh�d�� yɨ�rZ\��ݥ0Ndm�I��m�/c�@�{)�}����bS&)�H�rj�ܖ���vIh1XФJLS�4��ՠ���������s��@���Il'Ƣi���us���k�[s���� Pr��u���a���n8��Nn(��>��v� {u�B����n� �;�QUUUWw*�]��>�79�BIlR
�w�n�Ӝ�orJɫY|T�3JI+v���@O� �ܖ��Rݒ���Rl$���Q���@�{Z�����75 �7.��m���v�6�r*@{�K@��}��ޤX{�q$G?(b�L0!~�#'iN�:�Rɝ�s0.����ծs�":u��iN�Ȋ��>�~��w�h�c�@���he기܊d�0Ȕ�Š�l��"�����nhqڷ����
D��0���@���}�w4Y��B����*)�LGI(�DMUe]��s�Š�l�:�hӈqH��F���@yȩ��- ssP��h.��6�IL	&h�h߿;���w_��o��v*����wZ�n3a��N: �0r盅�#�e�퓏C���9����v�͐��:c������P�̴����%�:B#3,��i8��7&���V��n��;g =��?B��F�]u+���d�AswS�y�b�=�np脢&Mo� ��t��M	�LȊ��4=��w��X���ݷS������T�;��{/��a�ɒa�)�@9�٠{v�N��� ����?DB^����4�L�P����`�ev�qh��$v�u�v���;�8.s���}���t��\�>��h$T���- 9&���L�⑉��E#Zm��8�Z�l�9��ց��h�r'$K]լަ� 5�x~Jg[���wb�>�t�i	�$�KZ�l�9��h$T���-�=��	{fW*�Uw�{v�N�������n�~��O����)��(,$`		����w�ݿ���y���9���z�;�J��Vcd��¾������X�qK�y�%�x���Y��`I�˒q�ͮu9�,��0m�5Z�]����\�CK�Q�1���6��)x�:�x�`��=�`i4��W��8cn����� ���Y���xSƧnx
ۡ^s�D��!n��ݹ2�aJ�7�Z���n:�&b&�ݧ8���x�kX��zP�-��֥�j�5%m�[8��b��ˎQ�c��k����Bv΋=�������&D��N5�9�����v� �{��;l�Z��BpSs"�9�ަ�9L����w�8��g(I��a�I�#�"R'�_{�@��Ӝ:"���X��� �-��RJwv�)
��]�"?(I*��\����X�M�$�P�_w^ �{��-U��VUsws�ko�%	n�t� ��h�e�@��8�rF���ƈa����:�MQM9;�����v�G�V ݕ\@~{����7G�I�ܑ,�s>�������u{?|�����;Ф��&ě$TԹ�rI�{��PB�)A5PB1���)���	CX�)E�s@����2*�����Y��ק ��b�>�gL��ܦ��!�ő`��@���v۹��D~J�_��`~���L�Йv]���V��m�$�R�6I5 �܋@�^�МĜȣRG3@��S@��'����uӀ9m��>�h*�� �<�8'gu�ƈ���#k�t�3r�x�^z�=�]����-��o�P��h	rL@{��:��d�ueE!Z���wn��%
d����9�Om�@��X��p#qJ���� ��نGD(H��(M.P�B?%���^��뮜���H�������J�n��(S��� ;�� �ۧ:���y��zz���ؓd�c� 6�����������yPEq�9#q�`61!d�c$�ݥ�`��BL�&�<�ۧ�8zQ��	��{�>���|FbqdX&��Z���U�����������s�g��$$0PYR=�n��M}|`wu��-�t����lN
`��iE$zo�� �٠w�Z�
��@���3P<x�D�Us��x�Ku�9m�J�؈Bj���p�Uf�=��'�;sSVS���xdĜ�:�^����y�k���[l�;Ǌ��0X���"K�epǒ��ڬ2��|����v�V����86+'3������[^�λV�[l�9�Z��G�IƜ����y%�	$�<$��& m\Bx��"X���m�:�^�U���i��؏��]M�yD18�,�Z��r%�bX�w'���"X�%��{��ӑ,K����]�"X��u_���ٴ�Kı<L�ڇ�̚�	r[����r%�bX�׽�m9ı,?�}����ı,K�����ND�,K������Kı"\��x���Xh�({!! $���F�%�3�a��ċ(ix�!5�
��~�Z�4&�E�*�քp��R�S�������E۽:���'�)�-F4%`P�`B�� ~���ԢP��q5
hL`Db@`E�E��]leCP�@Ә����S���|UF'���ߖ[�Y-Ms4,!4�+��,c�\&e#��40�>t4�K��_�?������8�'c�'��P��)*GO�wN� �7��/���kY���v�h��"@ŵ m��h�ą�1C�W+G���F5 ��M�pI�jx$<��Lg7lvԨ�P��dmWg:z�� �w]���f�l�{lܓ�Sҝ�fW��<�r�.�ԇ
ͷ9���[�9ݧ�&ݶ8���/4���ӈv�;nv�D��a�)�DVp�6�)�'����G}�A���ֶ8v�!fD�9U+�ծ����Qm��3<� ���8m��ە.�{��^j�;c����;��!K��d�㎮�@.�FSWZ���7
�`x6����u�nv�&K[z�ö�����Jsv�>�np�)y[� ����4����D4��As�8���x���ic�Gm��7*Ux���gc����L�hz�S��' `[@�ht�M�*'mv���cc�ʠ�[=���`]{X�gmq��ϝ�3�v8;yKNe���E3X��n�u��!{jv8�m��V���3���{/!g���n��In�u�ث}����i����[=f��V�nL�9�k�MU�q���]���7k��Nm5���&���q�^����^
�Uv��Z{=��|��n��_lq �8�ͳ��l���x�sL���`���l9�8���=�*�j�k��Dm���m�@T�r�/K�F_QU*N��*ݵQ���Y;X��M�Zj,�M�9J��� ۖuj�V;u�4^f��ݸx���0:mdx���vn���7���d45��8aӶa����:��)�z_3��-�wB���/)�Ĥ�-U�V�n(�(g<�m���p���g��hث�n:�+=o6.ݲBH��6^3�kX�N׶8�H�����ݤQ�[����nn]щ�tA�W�F	�N*�ui��6m��X�X��)H��a��+�`�6�R�QgM�Lv ��ۜfF(+E7����i��ݦ�Ѣ��k�\Η)�O�GRk��s����k��ƑН�ނ�%�5��P��G ��B��f�5U��ѭf�k-�  �7�6 � �pS_��N����'� &�-n�9	���K� ,�A0N�M�Ka�Ɨ�m �<˹;r�N���p�.���.���Fy��`��4xv;m�GC���+�I�P�m��uՀ�t٘W$b�soR�a Ū�]�Z�Q��d۳�>Őۡ�m��U�CO=v�a���e��s͵���'^n��8��8���)�'�ۮ�&��r��V�m�&^�A�.�v�uIh��d�f����b�5�o!n��j9���Ѭ0�9�3���kxL�[�;b�k���l�n5�B�f�h,EO�����{��'�����Kı/��fӑ,K���=�lyı,Ok�����bX�'�'�NKf�ɩr]e�]�"X�%�}�{6��bX�'���kiȖ%�b{^����Kı>�{�iȖ%�b{�z����dӢd��3iȖ%�b}ܞ����bX�'��{[ND����j'}���iȖ%�b_�����s{��7����������+a���?x�Kı=�{��r%�bX�w=��Kı/��fӑ,K�����o����{��7�������dY'��Jv��bX�'{���r%�bX����iȖ%�b}������bX�'��{[ND�,K�|z�묚%�$�a�jiӇN��qBW<v�g[pgfi�ԗ��y}�f	�h֦e��k.ӑ,Kľ���ND�,K�篵��Kı=�{��?D�K������9ı,O�=�u�I���S).����Kı>�z�[NB�qQ`�@l��X�"n%��{����Kı=���ӑ,Kľ���ND�U5���3���2k$%�nk.kiȖ%�bk���[ND�,K��z�9ı,K�{ٴ�Kı>�z�[ND�,x������(=7#Ac5_{�[�oq���s޻ND�,K���m9ı,N�=�kiȖ%���M{���6��bX�'����NKf�&�T�.��.ӑ,KĽ���ND�,K�s�����bX�%���r%�bX��{�iȖ%�b{^���!�\�&Jk5n��o=�`^��łW��a�GCr��۠�{}ۻ�Ք�k&���fm9ı,N�=�kiȖ%�b^��ͧ"X�%���v� �O�5ı/����iȗ{��7������9��l�����߭�ı,K�{ٴ�A�,K��z�9ı,K�{ٴ�Kı;ܾ������bX��������f�f����ͧ"X�%��s޻ND�,K���m9ơ����"j's/���"X�%�{�{6��bX�'{'f��h�4k3TԺͧ"X�
�D׿���iȖ%�b{�����Kı/}�fӑ,K!A,O�u�����T��J���r���Ē	"}��q7�F}��6��bX�'�����Kı/}�fӑ,C{���~�{s���n1i���-���<6p[-�-]c�*��v�j�;�w{���\�73SY!.K����ӑ,KĽ���ND�,K����r%�bX����j
r%�bX��_{[ND�,K������f�U�������{��2}���NE �,K���m9ı,N����ӑ,KĽ���NDı,O�Ox�,�ԙp�.�36��bX�%���r%�bX��/���"X"ؖ%���r%�bX�w��ӑ,K��ݗvM�k&���fm9ĳ�����������bX�%����m9ı,O��siȖ%���F$���P���!@b�|,TG���%�����r<oq����������+e�-���D�,K���m9ı,Q���]�"X�%�{�{6��bX�'������Kı/��OkSY��3P�j�0�E<;����+�8�`�7-��d �Jc��Y ����o��dY*�?{�[�oq��O����r%�bX����iȖ%�b~�O{[�Kı;�{��r%�bX�읛/��hѬ�SS3.ӑ,KĽ���NC�@����'������"X�%��kiȖ%�b}��ӑı?zwz�ѯ�����K�fm9ı,O���kiȖ%�bw^����K,K��}v��bX�%���r%�bX�=3�T�̚�	L�535��K������"X�%��s��ND�,K���m9İ�y��Y����$/WwMT�YV����]\��ӑ,K����]�"X�%��{���6��X�%������ӑ,K���kiȖ%�blh�����t�2HL5�f&j�&�[��u��#���d��ԣ�J��nݧ8�0h�����r�رL�s��q�a�l/ ݩl1�#�ϩ0�g
�v�ѻGc%����j�>9Pe�t���;����ood��cۓ��pӧڤ�^sNC��Ap�i�v�-qv^�%l=:�v��s9D����Ƿ��8\[vnURq�痉�d��FG��@���Z��V�{���wｚ�8б&]F�ƍ�;R��z�@�x��Z����.����k������ݻ}�Ԛ�R�˙v��bX�%����6��bX�'~��kiȖ%�bw^����蚉bX��{��9ı,Ow���YO묺i-�fӑ,K���}�m9�#���b{_����r%�bX��{��9ı,K�{ٴ�ı�{��������+e�-���oq��K�����"X�%��s��ND�KĽ���ND�,K�e����K7�����ߟ��%]#��w�{���lO����r%�bX����iȖ%�bw�����bX-��{��ӑ,K��d0hѬ�K���iȖ%�b^��ͧ"X�%���W�nki�%�bX��������bX�'����9ı,O����R{Y�乽W��;<x��v��Yh.ӓP��d��8{Wa-k�u�8�{��'ʮ����Gak�w�{��7����kiȖ%�bw^����Kı>�w�b�"X�%�{�{6��bX�'OL�����I%3S535��Kı>�{�i�h�Q�Q1Aı,O����r%�bX��}��r%�bX�����ӑ?�b ����7������A�v*���}��oq��%��g��ӑ,KĿw�ͧ"X��%���=�m9ı,O����r%�bX�x��I�kRk5K��5��ND�,��{6��bX�'���kiȖ%�b}���ӑ,K BĿw�ͧ"X�%��ޗvj�z�]:!����r%�bX��_{[ND�,K��v��bX�%���m9ı,K�}��r%�bX���ѫn�h��j�42��v:���u�)u�=g��F�@)�� �t�4=���௲s;��cK�G����X�%��s޻ND�,K��{6��bX�%���m�Kı:w=��Kı?h�ޖMMk5s0�tY�˴�Kı/���iȫbX�%���m9ı,N��z�9ı,O����r*ؖ%���a�CDѣYa�35���Kı/���iȖ%�bt�{�iȖ8��
�(� $#�����ڃ����s޻ND�,K��{6��bX�'�L���OjkZ�W)��Z��r%�`�bt�{�iȖ%�b}���ӑ,KĿ{�ͧ"X���D�Mw��ͧ"X�%�����kO�̚�%���f]�"X�%����]�"X�%�#~���ND�,K���6��bX�'N�v��bI
H_���G�򫛪.˲BB
�L\\�m���]AF3�'E*���۵�V6��k�M�"\ְ�.��x��X�%�{����ND�,K���6��bX�'N�v���bX�'��v��bX�'�=|Rp՚5���Mf�6��bX�%���m9Rı,N��z�9ı,O��z�9ı,K����r%�b}��ݓE=Mf�Cu���Kı:w=��Kı?w=��K,K��{6��bX�%���m9ı.�_�����h%��w�{��7����]�"X�%�~���ND�,K���6��bX��q(�lMD�����r%�bX�{~P���Q�f��߭�7���{����iȖ%�b_��fӑ,K�����ӑ,K�����ӑ,K������~~�s��D��ۄ�1v�3�����vf8cQ�ݰtV��Y�w6߮�m�]�{/Mf��35���ı,K�{�6��bX�'N�v��bX�'��v�"X�%�~���ND�,K���ֵ=��MY���ͧ"X�%�ӹ�]� �%�b~�{�iȖ%�b_��fӑ,KĿw�ͧ"uQ,O]˩g��Md����̻ND�,K�g���r%�bX��{ٴ�K�,K�{��r%�bX�;���r%�bX�k��ԗ5p�f�JMkY�iȖ%�b_��fӑ,KĿw�ͧ"X�%�ӹ�]�"X�%����]�"X�%��O_�5f�f�rSY�ͧ"X�%�~�}�ND�,K�s޻ND�,K�s޻ND�,K��{6��bX�&�m�A,A�?84���c�c�!ћƯ�L����9y|r󥼗N�u�ԤvܞBwM�s��V��.؝�׮'�X�]]HIrt<�aU\�d��4�Cn�G�m��`�]λb��i�m���nd�6۩�糣5�F�a��a���۰cX�k�V�M��&-����m��Q)&��<m��Tg�gcu۹�q'679���n�v�7�	b��O	���ߞ�w������f-P�=��Q�6�ݛ��ի�V�-�2�cuÎnyMFᰙ1���v달�'"X�%������Kı?w=��Kı/���kȖ%�b]o�!|B�����{�eUئ쩻��љ�v��bX�'��v��X�%�~���ND�,K���6��bX�'N�v��bX�'{�}�M9s3Y�fjMf]�"X�%�~���ND�,K���6��`ؖ'N�v��bX�'��v��bX�'�!�_h�Ѭ�5�Yu���K�,K�{��r%�bX���v��bX�'��v��bX��D�Mw��ͧ"X�%��kZ�ښ�ѫ�2��36��bX�'��]�"X�%����]�"X�%�~�}�ND�,K���ͧ"X�%��ݾ՟�M�u����웎�"�p�v]jԋ��
�t�{u�Qƛg�!,s���c��iȖ%�b~�;��Kı/��iȖ%�b_�wٴ9ı,O�s޻ND�,K���u%�\%��%.��˴�Kı/��i�|����B �1�	#�"�WKR��L�DH��� � �	i8�����0)�ʆ"|�%�b]sٴ�Kı<g�ӑ,K���w�iȍ�bX�t��I�WE�Z\���fӑ,KĿ��iȖ%�b~;���r%��AuQ>�{��9ı,K�{�6��bX�'�z]�4S��i�0ֵ���Kı?�z�9ı,O����9ı,K�{��r%�`��}�fӑ,K���{���n+3,�T}��oq������_�˴�Kİ���6��bX�%����ND�,K����ӑ,K��]����ԕ��q�[s��M�wX��Vnn0q=X}=�Gvؔ�k�N!�w��믨��SYfh�̻ND�,K���6��bX�%����ND�,K������X 蚉bX��{��9ı,O�He���Ѭ��Me�fӑ,KĿ���iȖ%�b~;���r%�bX�}���r%�bX���ٴ�O�b�j#���9����*d���5}��oq�X�'ǳ���9ı,O����9����F$���im�ŁF.��&�d
0��������*�*Ȥ��	��R�����4�*�Z i���f��r��*Ml��.����@(�!`@��{p��kR�H�!�C�)��~,
��la@��5t@�d���/�a���tDx"p��bVq?0B����л�aUH1""�aB���E��l"��Ɛ��� ���1i�<C�hO�C`~sL1�(�@��RQ(E����Z��+�4"�mE�QЊTG��| 	�
'��(�� m(���U�v"�(<�"X�|�ٴ�Kı/~�iȖ%�b~墳�˖k$��Ffe�r%�b�����]�"X�%�~�}�ND�,K���ͧ"X�%���{�iȖ%�b{^�������Y0���e�r%�bX���ٴ�Kİ[��{6��bX�'��]�"X�%����]�"X�%��]�&�fML35fh���ry��W-�DWE���D\c���J�9��LBt=I������)��ͧ"X�%�}�fӑ,K��w=��Kı?}���3�MD�,K�{�6��bX�'{�.�)�Mf�CkY�ND�,K����ӑ,K���w�iȖ%�b_��fӑ,KĿ��iȶ%�b~??���^�>�~����{�����]�"X�%�~�}�ND��a���~￳iȖ%�b|{?��ӑ,K������c�35��.��e�r%�bX���ٴ�Kı/���r%�bX���v��bX ��'��Ӑ�!I
HRB�
�k��5E]e]�fӑ,K��ﵴ�Kİ�z�9ı,O}���r%�bX���ٴ�Kı?�����-�4h�u�Jkv�(p]�Y쩱��q��X$ۃu���n�L�]�GO�~r�㣒��w�{��7�����v��bX�'����9ı,K�{��r%�bX�������bX�'���h���Y����33.ӑ,K����]�"X�%�~�}�ND�,K����ӑ,K��w=��Kı?w;캒氚4f�Z̻ND�,K���6��bX�'��}��"X�%���{�iȖ%�b{��ӑ,K�����NZ&��䦮�6��bY�Q?����ӑ,K������ӑ,K����]�"X�%�~�}�ND�,K����)OS3M!�kY��"X�%�����Kİ�P������?D�,K���ͧ"X�%��}�kiȖ%�bl?��I����[�"�,i�z�5IG�<���¹ć0�;,���l��{���ǩK����9x�õ�>��_��m���z��0ɧFؚ�2�ѵ���ix�q$OI�cC�;j)��t=���ds�0��2���<h(r�$��,�F���9��k=�[�n5�������z�˥�tC]�N��h��y��>u�釪yksV���� �&��&Zs\ɢ�WW]����v^�>�mǛ4���7Nr#����yx�>���}���qZ�e����,K��?����r%�bX���ٴ�Kı=���m9ı,O�}�M�"X�%��gg�)�\��f\�.�.ӑ,KĿw�ͧ"X�%��}�kiȖ%�b~;��m9ı,O}���r-�bX��$ç���SY�\�ˬͧ"X�%��}�kiȖ%�b~;��m9��U`�����]�"X�%�{�fӑ,K��k��׍kR��S)����r%�bX���~�ND�,K�g}v��bX�%���m9İ����ӑ,K���Sz5=�,�BR]�ɴ�Kı=�w�iȖ%�`����m9ı,Ok��[ND�,K��o�iȖ%�bx��Բ�y۟�\�۹�@t3ss�͢�-��6��۶,v��/\��[vy����}��oq��%�~�}�ND�,K����ӑ,K��w���)Ȗ%�b{��ӑ,K�����',։r�䦮�6��bX�'��}��!@���V$ʉ*H T�` '8(%�bh����ӑ,K����z�9ı,K�{��r%�bX����rRz��i��fӑ,K��w���r%�bX��;��K�,K�{��r%�bX����ӑ,K����hֽ!fd�k.�Z�fM�"X�@  %��\, P�o� P������
�?w���r%�bX��v{2����feˢ�2�9ı,K�{��r%�bX����ӑ,K���o�iȖ%�b{��ӑ,KĿO��]Md�Omst���ѝ8t�ψ��C��=��-�0���:v׉ܽ��{���n��w�xxm�0���Kı?���m9ı,O���6��bX�'����yı,K�{��r%�bX��{��f�kR��\��5�ND�,K�}�M�"X�%�ﳾ�ND�,K���6��bX�'�ﹴ�Aı?w�ލOe�5���Y�ɴ�Kı=�w�iȖ%�b_��fӑ,x�$��D���@���@DE�)"X��w�m9ı,N����r%�bX���j�IskRf�ֳ.ӑ,K�����"X�%��}�kiȖ%�b~���K�����ӑ,K�����'�Yi�.���"X�%��}�kiȖ%�b/��~�ND�,K����ND�,K���6��d)!I	����]Ab(��*�E%uC����l8�rv6o0�e��b�r����������ѐ�2Mk5��Kı?w���r%�bX�����r%�bX�w���b蚉bX��}���"X�%������fL�e�f\̛ND�,K����NEı;���ӑ,K��ﵴ�Kı;���iȖ%�b{����c�35��.��e�r%�bX��}�iȖ%�bw_w��r%��bw�ߦӑ,K����ӑ,K���e�5�h�-˒��"X� ؝������bX�'}��m9ı,O����9İ1<��,��dOg}�iȖ%�b|k��f�Mj�W����m9ı,N����r%�bX�~�w�iȖ%�bw���"X�%��}�kiȖ%�b{_[=MEySo�&7��;�Mm�g�'Vz�]c�� {�7b�����>�;�۱؊ɴ�Kı?{;��Kı;���ӑ,K��ﵰ���j%�b{���6��bX�'�����k0ֵ&a�k2�9ı,N����?�b#���b{]�����bX�'����iȖ%�b~�w�iȟ�PD�K����$�.�Me�h���6��bX�'��kiȖ%�bw���"X�%����]�"X�%��w�6��bX�'��6R�\�!�kY��"X�(%��w�6��bX�'�g}v��bX�'}�p�r%�` �'~��6��bX�'}����2f�.�2��r%�bX�����r%�bX"{���ı,Ow���ND�,K��m9ı,O��UD����7J�E^�nW5󐙙u�f�W0�rR�3عЀq�A	u�z{s�7���yR��uY��|�Gk�^2�nk=�T�n�7R�ѹ�����ͥ��H�V�]�5NƇ���/�R�sc�9�R��E�ǭ��Nxg��4�qTW��Q�N��;9I���t�NG&9�Ý\�GP�v��1\/.��q
�	���cB�7N)v���b^Z�v�7�D�̘p�5�sVٙ��jL&Uúi�^kT��K�ٳ������Lk$ߝ�w{��>*D�®��w��Y��bw����Kı;�w��Kı;���ӑ,K����ӑ,K���0�]h��Y-˒��"X�%�߻�M�!��CQ5�����m9ı,O����iȖ%�bw��� �%�b~5�{34K4�ᚦ�Y�iȖ%�bw���"X�%����]�"X�%��w�6��bX�'~��6��bX�'���sS^�usD��sXm9İB����ӑ,K���ND�,K�w~�ND�,�"(�{��ߍ�"X�%������&k]I�B�Z̻ND�,K��m9ı,N���m9ı,N����Kı?{;��Kı/�u�~!�mWN���l�Ż/,��޶y��<u8�^��K�ےd�}]v���w����m�+ã�f���"X�%�߻�M�"X�%��w�6��bX�'�g}vȱ�5ı=���ND�,K���f���̥!�Z�M�"X�%��w�6��E � $���]�%�bwپ]�"X�%��{�6��bX�'~��6��)bX�'}��$�2f�.�2��r%�bX�����r%�bX��}�iȖ?ʰ�MD�}���Kı=���ND�,K���d[X����{�[�oq��ۻ��r{��ߍ�"X�%����iȖ%�bw���"X��]D��~��ND�,K�����&�ufan\�Xm9ı,N���m9ı,?�X���ߍ��%�b}����ND�,K��m9ı,Ok�-횾˩��2\2�n�y��n�h��s�Lu�ݜ=���3��Lq���������Y�W�5�̛ND�,K��m9ı,O����9ı,N����Kı;�w��Kı=��.�Mz����.k�"X�%����]� �bX�'}�p�r%�bX�����r%�bX��}�i�!bX�'{�^jٚ�TјB�Z̻ND�,K��m9ı,N���m9�jP�@� �H�#*F"�  �� '���8H��o����"X�%����iȖ%�bw���N�.�S-���6��bX!bw���iȖ%�bw���"X�%����]�"X��Q=����ӑ,K��稜l�?�fh�2kZɴ�Kı;���ӑ,K�_����9ı,N����Kı;�8�_��$)!s}J���L�wWU%sv�M��y�[���a㵎R1vu�p)�@:��������|�wm�Ia�Vw����,K����ND�,K��m9ı,N���l?�蚉bX�����"�oq�������[X����{�[ŉbX��}�i�#]D�K����ӑ,K�����m9ı,O����9��MD�:x�{�d�.��.Meְ�r%�bX���6��bX�'}�p�r%��X�'�g}v��bX�'}�p�r%�bX��w��f��ᚦ�Y�iȖ%��X��}�iȖ%�b~�w�iȖ%�bw���"X��8
 1�(]X������H�y�M�"X�%��i�kW�%ֳE-˚�iȖ%�b~�w�iȖ%�a��O{���ı,Ow���ND�,K��m9ı,O�e!��u���Fa	2�=t�=��]]V3���Ö�%��f^��n0ŀ��4f�ֳ.ӑ,K���ND�,K�w~�ND�,K��l@�,K����ӑ,K�什	̙�%��j٩��iȖ%�bw���i�
bX�'}�p�r%�bX�����r%�bX��}�iȟ�(�����$�����J�UfB��$%���p�r%�bX�����r%��%��w�6��bX�'~��6��bX�'}�^,�2f�.�2��r%�g��@�O�����Kı=���ND�,K�w~�ND�,U[��m9ı,O{;=�rL�3Z�˗Vk2�9ı,N����Kı;�w��Kı;���ӑ,K����ӑ,K���'��@�hi�M�4�?-wv0�A�!5��	�XSk�hq�4B�J�Z[㈆��$8���WQ�B{,4�ka��f�(�)*ȀPX� �SiA�A�ǜ����Bi8	�_ı�~��F���޶��Q�H��p�۲n��4�S�i*"r%�"Л�j`-����on�?����R�UO;�  qmH��"��q},��ķ #��Z��7�4��2`M�к�l��cqp�ʙ��&l�)ae�!�"у�W�CF^�|%<�x�qo.�l���`s4v���i ;F@3����^�Z��\ҫ#� <����4��mz��g�Rls��q���9F�nU��\�x��mo)e�9ĩ�յ�^prir�u��;��̸m�}a)�kB����'��Bm]-��;e))������}�;I�����x5Ó���i{-!�r�m�X:M@�ݶݴ���Pʎ6��7J��VL <��4��G�Ӓ�x�g��}׉0��3�m����n��$@����9�*�UC��%b6�STT��r�H�H����ܔ�y5ع�0=�h��\j �ـx���'x�ݶ˛u�q���,�E�����������R����:��mq킬m��%L�.���	�Ɇ�&��y�̄츅q=�
�SU�����#�)�`�ct���5�q��NУ����� V�b&h�� �����у�E{2m��s[/�y�mc����fkd�7;C::p`��F�qD�VƮ���k�nK���n�(���m�zr�J�1UC�"��M
��QuJ�ec���[�)Yn{Bb���؍�{DAd��oc[/Y]q�/<�l����U��|���Zm�)�瞎�Zɘ�5e�$�(�Gl�q:��)����֖�f�ш%}̆ҧZ��yGt���3Θnp+6�vpjƳ6�^rn��x;tt�V�qtbg�,�K�mx{,��l�
H���T��{xɎ�X[��c[��u<���Kی3XP��m ���3A��D�M��f��{ -�9�i��K��j@�l��v�mQ00�
�q�k�iy���s��H�:-�NnϮa�v�a��w����-�j�)��  Z�X��#3<����{�}����{ݤ D�*u?*~�	����\T��D_�ǽ�{߷����BI��p㜱�Zܑ<�$݂��$�ר�K+�읩v2���E�yg�4�
Z�,=�m�.�85�\fr�۳$����R�嶬+J�]�Kja�Ƽ�)k�\�݌ur+ν����z��fw��8���O1`�Ɨ!&�=�N֎ɍ��U����pq��6��Ʀ�PR9���v^:�A�s�9gZ쮺�\v�uສ�	�g�{��y��o����:�tʣ��GE��ST���K�pd7n�^
ph�76ߞ�{���z�;r.��5�Z�iȖ%�b}���iȖ%�bw���"X�%����]���5ı=���ND�,K�^����f:�f���d�r%�bX��}�iȖ%�b~�w�iȖ%�bw���"X�%�߻�M�"�X�%�淪-l�Ĝx�(������$s��h��H�`�q�H72�w{�Yy[�)�����	)|��=w��^,�ߗ=/��|{���`�5��4�m��>�|��N�^,��e�j�]*��PX�exӝ���axmgKy�Jkf:�3,?���n��fh�0��>��Xε��^/о�z���<O؄HG"rE���V���aJ��)��#$}�� m������E� �nH�m�"�;{w4��0䒙|��Ӏ{B��r�4�&(8���w���;{w4��Z�߱__}�1Zߢ��?525�9^�X(��[��ϱ`�`���m�-�:}���Uժ�&)֊^�8:��n���uٶtT�g�@m&���x)���|�\����7�l���Q	z����s@��։(��b�ȴ^�X�m���Xε�tDDɽ��e�V���]�U���� �׋�4����
��tT�DW�|� �o ����T&�˥HVUU�
"[}��=��p�x���4���!Ȝ��f��}�@����|�|`��`hm�w6�lO&�79��m�ǚcLv�{,����)��"�`#�� :Z�z�,Ī}���ߖ�� �׋��t�pЩt�ƛ$�s4��M�f$[}��q���>m�������[��S%�M��Wuv`�ŀ}��p����wb�<���/*X(��X�)s4?�r��O���nIϾ����GKрT  <}��(Mh�!�&fb�,"���rJ#ߢ���,~�$��Eһ��s7m�"�������/������곮����n��[Уnҍ�ݳ�tf�<sS��ɻYW�w����v2.�s3v�9��T��c���.�yԱD3.(G�����sz!)��O� ��ŀ}�`��J��D�r&�$��>ՠr۹�����<h�ۚ+�c�G�(�iH�$T��=�� ��U����:���Ɠ�1dq�3@����?�~�������6�`�DD'1~4�.@�Ʀ�k<M�uNv��7K̻�\��͹��9vN*$��-�/T��;Q7d��Ј�܎��Cpt�P$̲c�Z���p�9�D���]���v|��q��Pmp��:��c���I��7\���7sة�:��Ũ��v�,�G�xn��t���G�dG�������p�&^:�8����+�����%��ɉ��͗���::X{���{��}�߯���pl��ѭ�\��\�Ĵm�ո��9�v�zv�Sre�sKEć%�t]��{�`��X�x�(_�G�7�_�S�bQ��H�(G3@��k�>m��>�l�7u��IDL���$��EһB�����݋ �]�DL�V�u��얪�T��(�V�����R���I ;��^�Bj�]*B���0�x��J#i��������M�<]���!cnL��:��^Ί<9�Ő�����R�^�:m�n3<��1Js���nD���qw��[w4�e=�33>Am���Y�L��8�m�L����{�b�V �@m���� �kŀzw]g脣�P����9W�,�ݫ���ͤ���� ۊ�m�@}m��>�kv)�1L�dRCC�1(K�Eww�,�w��>m��>�l�*Yj�mā(G3@��k�=�3���|�_�X���$Цj*+/g���̓��+�y�qo.-p�]�v���ܙ�y���!F�s	!1~I9���s@��3 �׋��Ce�����wV���U�]��>�l��$�)��ذ����x��Q�*��fK
�t��!]UU�w~ŀzw]a򈈡(��� D���#"B$"i�J�B�����`�ʥNФ�#�6�&hy�4�l�>���������f��Y�L��8�m��ɠ�j��E��$�*@���ԙx��j�۷g\i�hY޻����T)����OnL<�lg\q�Ҝ�ۣ\�q�W-U���;� �׋ 7�������)ު�L&4��Ȥ�����hy�4�l�>���${�Ko� ӆ,J�@ϵ zI�G�@6���x\�HL_��C�s���9�<h���ܝW���j�ؐ(D{�D�/D%9�>��˓�Z&�]\�m����I>�x9��I5�����N,�tv�Y��n�=Bw\�Sq�v����ON����y�f �ζ��{v�fh�m�H�=$߽a�M�@_z&�D�r&��� �;f�}m�ײ�{۹�H���G332�su w�}�G�@6� �ɠs8Ļ���I�#rI4=��=w� ��X��x�S=�׀yI�5�6�i525�I��s@������������s�gf����Dʬ ���8=n֦�KsÑΕ3]S��t�F��^�ܞ).��\r=Ƙ��gk<r�E�5ƍX�j��Su�+���ָ�$�%��l�#�P����M�z5��g��m�h���%V�.�:�c1�,�I��\sFȈv4�Q�b��i׳$E��:��s��k͞nQ�Eu�ɧ'wH�5��7T��"紮c��9�s��L32a�5���9�[��ʮ�z����z~�߳�"�O��n ��9Mr��tApQ�vܔd{
;�
�ny �WCN�(G3�����f������=}��s��X\	 �~C�M ��~Q
��w��}� 7��?(�<�x7s#��$�=g��۸�9��},���Q�[��nff�G �j |���_}����� d�G"m5&hy�4��{����J2e�^��eFY*Dn����ju��̊[��Ml]�6�"ժ�������}G=a��W����\�P�`��qR |�'ao��SFa)�Z��ܓ��;7�H0Y����P�3&��nI=��7$��l��b=S���725�I��� 7���!L��^�w��������cě�= �;f�s��@��3�_��[}��`����h��S0ww��w�~JB�<��=/��}�h/SM+�	��x�L?<x
���-��&��qDv�Kmr�p�.�,��o�����}���0p1L�I>��Ɓ��@;���� ��@��0g��$�m�`N�Y�%	L�-�`-�`k�`�+,s2Cj4��@��k�8��u���3�on�An�1�f����7CY�$hkaW�%���Sl�FńGL�W�% �3K���@����#�@)������ܿ}�A	kB�iP�����BBoj98RH�t����ȁ��wP�lCa��ic��q�� E�XP�;G5�چ��l��P��)� L6�V��]�{��GF��	�q ��O�k��6hJ] i��U>O� BB$� �E@!d a	�SN+�!�DC�O�0~P��Q6��h0�7>����:��@��,���F�a$z���d/�!%N��V���ӭ���u�^1.�bǒ`�!���l�����	z�u|�wN��u�}�j��&��5�o��c�ݞ�;�\v�Ԫ�p�����ڸ9J:��Y��ۋ��:*߭����V�M���u�BQ�}|`nf6���cě�=�ڴ���`Kn��(P�OwuJ
ʴ]ݩ�ŗ�hI��<�T���1�Z�F*��U���d*��9B���}��==�X�Z�/"!D H!(B� E�1��� ��%
�BP���x�T͈���]�wwv��& <��@��7 ?���ē�1(���Q�&$�#s\՝�^�9l�[Pl�a ��*^�wwww�?d~bHbmF�q����h{�4�۹�|��@��Y"�"�F�bR- ��y�IL�o�`���s��~H�X�=14�$�dM�&��}���?D$���Ӏϯ ��w6�&5"�ԙ���1/z�h��h������`�3uA�b*�T�oowPx�	�����j��
D�B����zd��k532ܗ 	ŕ�XhqQ�[;�	����ȏcz��ݧ����Nc�p�Z�A8*�*��OC9۲��3m( m�v,/,Ƹ�l^x��;Tu�:za�	���d)�lA�����V�sڊ��[0�m�u�Ju':uF��dY��� n�nz� /[Ot���;q�R��X3`\��Z�W�.�5��`�3�%姃�?���޻����;L���]�k�u����N{5�q����mru�75M�קsۏ�wg�ٮkX\�I1/���z�hu�HG5�Z�r���Ѻmm�f�<�T�$sPx�	��(�*#�O��\���ˣ0�L����߻��mk�?$��;�^��k�UH��Q�94?�~���1r����׀}��`z� �M�sr��n�ʪ�&n� �xD(�K����z�hu����x�j
D�
��z��5�g��mΉQс�n����8�L��!6E1��)Ӓhw�s@-��s����׀9�����j�53+��nI;߻�Ҍ� (��@	���C�D��k]�'���p>�n���Q��7x��I�}׮p�w�(Jϛ�X����Ђ�-M��&	&�p?$�%3���7ذ��X�J�����"q]�-XM�s!Ww�}��`�#����t�p��ȵP�8��L�~lı�`+l����t����:��`�l���r�4aݙ2'�d2)��|��@���h{��D}!���\��BK�MT�M�n <��@��7 =rL_W����|��E)�cm�)�[}4�^,%JG�۬�s�2g��c��i�4=��1r�}���}�ڴ?���hyx~�bDƣ%�Tݬ�m��y����׀}��4^�/Ἅ��##�cIbɂ˘�nצ�-*',N��7�n�F�D����{��˷ը�Ҳ��778�}�� ۚ��qR�mz�W�5�r`�N- �{fr��O7ذOwV�ֹ��#��e5&9�DH�@���>Vק����r���M��
2�O$�dR��`Kn���� n�Dy%
�'��ґ�4��B�.��H	�b�lgu훒w�f���"A6�I����V�����m��[���mz�f,�U|G�a�, ��>�^�\��tv+`L�gQ��s1'',QP�"��m�%"���}����m߾A�s�U�1�R	�&�<�T���1�Z m�]���_��yb�@<�7�/{�@��� �9٠}�]��ԣad0n�&㕀}��pw]�n�X�'��Հw�h�Suv��I�� ��xۯ��� �k\��X��%�ЙR�k͑�]5��Ƙ����dzv�
���1�K�-u�v�+xQ�Mɝ�ä���C�z`���S�Ѧ�\q<�s p(�]�YKy٨�)���k�b��;������c�4W0�'AkE�uͳ��㹴��^�i��-�Ջ�p �����L�:I=�BgCi�tv��\�l<m�{<`Y����E47meMi��.^ڨ�i�']��{ݺ&�&l�qg�c��㞝�i������^Ͷ;�Ūڎ�"c���M�$ړ�F�H��^�ۚ�Ɉ<r�nj�^�`J��ݭ+ov�i�b�� ۚ��qR�~H�<�Q&�i7��6�<�T���1 ��{�Xm�V�j������ES��x�~ŀ}:�`u�� ���ы��M�&��qR����9h�������f��D�[�����&nڞ�K��/��7�k����)�2��_��=��'Q��`�}�<r�75������wb*�T�j������|����*Q���SAO���,��� l�5�r���Z������i��.+�=��-��F�Rc�ډI4?B��}��=/����� {u���؊��]���ݬ��� ��#{;���~��׋ ��j{���W
׮�����\��;�,�η��;6�\yN�פ�ǣ���	��������9ɨ7 :ܘ�nl��0��G1��ԋ@9�f�g�H�Ɓ�}�}�ڴ�,��$�9���М���ܓ������@" ���E�  ��E���{���ܒ~�߯ �r���J�UUj�b�����R�}� :d��95��n�r��؊�)�����s�r����߿_�����qvנ}{X�kx�`LS{C�[Ձ�S;HAד��7b��c���{��n��� rc�@_��@9�f��{w4.�����9]��*��i5&'��������׋?(�6_u`t�p���?bE�P���7�d2)��u_z������2k�u�,�wAIɊQ4�I���-z��4s�f�La#�����!	
��2B,"�u�T�V�R0�Pu�0GNxE�w�y����H��H�4��8��M@w8��������̼�,�dq*N�4z��:j��h��5��3�4E�&TIW�\����c��lVk��u�,ӭ������(��@��x�{�<Lm��/�I�mz˖� {[��׋:J&Mnf�R�T�1bM����y�-�O�.��s@���@���f8�LX�9��?b]���7_b�6u����%������ŎF8d��rh�n���^�����6� ��B�*��I,XB��.�����%>�6��~�oZ6�c�7���H⁹2\�,�Zg?r�*�#At�qN)����:2P.���l�f��#��3$?a��S� @�)B��d�CB'�5�$R����8ŃcČH$J�UM���pC{�o&�A��	���m��
*k(�k�0�?+�HqNI�
D��L̩����g�%�cR	޴�茐IÊl�w6!�vE���(K
�b��:.�FI�/
p�S����ӧ�����}�m�[�mv�l� 8�������{8��Y#i��X-�,�c�����+�� �S�.ŧ<�2ۃ8LH�<Cd��#]O:���=ړօ�u�n�l���:9 `ې�W\ӈݺS��"��Q;=D�G&���#�Q��@%� ����%6��� �h�TH� �������m�­��t�沏;�;/��ȝ(ή��t��Iѝ$.��u�Sl�m����=L�UmԪ�d� *;�%xM8[��ts�tn�G�v�0�׌�]�,)��[F��nƣ��)i��7�;d+Q��3��;�m!�j��8���v��Sl�[f�a�,[j�!�u22�d��Hv�Ji��)mɮ���yZU�U��-th�B\��DaA(S;z��x����Y9�v���t�V��f�պ������E�{[�7�:ڤ�Иy�v7uؗ�H�a,��[���k$�p�l�L�^ݹ��m+�v5���t��h��p�p�Vm�+ѩ�׶���{f˽:�dR"]s)R	n�Վv�;�9�XVP*7m�'��/Rݻd|[���&�Ϊ��ָp�s��;j)kh����9q���S���NsJ�B��I����/*��U:��%Z��C'.�P��S���Щ+��M��B�l�2lCÎ�pHf��S�F����\-^k�c����5�Ck�nόCŭ��ۘ焪�ͭԥ�mt$�x�����1�9!�qR���E�4�MΕfy�&�vc�m��5ۚ�{`�Z`�=Nz�e� �Μ�\��շslR�l�K���CȗG`����M�u7$�8^��$�.���f%�A۶)m���k�Q\m��7Z�8�F4g�<<����-[�,N䶀v�i���5JH1�ڒk4ӵ"�֮T�8W�5ȇ8ɹ<�x޺q��«y:�'*hn�m�'U9m�j�VsZα �A/^�t  Q�{j�������PM����&���.��mE�Ȇ� �|� )���T���W��P���U�?M//��'�#խ���ъ���k�rrhpv�g��b:۸��A:ջS�;[\8z�.�a�	@F�2{;��oEYLCю&�1��Kcg#��K�\�����fyUb3��+6"��1��,����p��%۸��
�M��e]�ӵ���@������u��!{ \gŁ��۬p���ݹƺ���Xdon�vI�3f_T�j�fO׻��{������?x�� U��$E��U���D=vLbw�d8��i��Ӵ�%蜩�ɝ�7')7k �}����� y����$���������8��-z��4s��W-{���}�ע���16��= ﯦ��vS@��@��ՠ����[1b�OjI�>{�����j�WHG�ɍ�1�Ȝ4�Z��z_/�7�^��f�Dm	ҢJ*���-��/;�����3�5�mx9�vVL�2�C�D��b�6��ŎE�8bě�?����^��7�l�K�;�Xq�)
�Uujԩ&��p�]��'P��;w���^��}�@�H��c�9�����*@;�1�Z ��=��0@�7�����:�k�>��h/l�;�����$dX�m(WXε���>��z������������t�Ƭł�<>�W5�9n�mnn#m�v���[-
<[�GSay�W{��;��� t����V�w��u��b� �&�@�;w4�&�=1�@u�����^�dժ,W7k >�w�|�\�/D/�:`$X!!bEEdY"B�
@C����ց{n��tQ��bƜ1bJG&��D%
}��p�}X�^,��B���M�=�l��1bR-���@|��P����̿۟��U�����켷<Dz��Oj#�N�m��5������%�c�9��jH��s@�qR���s�wZ+2�\��j���ŝ	(���l���9{w4ޓ,�k$i��NL�;ɰ@u󘏮���H|� �ܹ����#�&�i�@��k�;{w4�n����w�t8?wYɹ$����SU�)�'zon��-��;{)�qs����<���#q�?ɺk�5��>:m�v=�':p�v�m�=��N���1�[���@m9��E&|;�nh���8��������Q��4��)��>�_9��*@{�T��������6FI1���h]�zon���.w���/��Uz�MH�seT��`���>z�`�ف�	(�_o����@A�7��	��}{ c��9�G 
�(��~�ں��s۞ˬ'.X�,�'c�_w�S�qHn��-8��:K������L�s��,A֑�ݓ��.kd�u6t#��"iT\ƴ� � �cVt�Y�n؆��Ѻw��k���'Ѯ�veC��J5Ny�ڻƝh�;�y5g�ӳ#;hq��ci{u�^C�6]�DB�U�j{3n���WS9Ȧ�ol�uʇ'E��{���~���ju� [�F�"nv�뉣�]����3�
�gT�6yt��H�]��o���`|�=T��qRɹson�v�sp��ݴ ��@z8�����[���tX���H'����9��HG c��9�	e7+r������J�ݤ�����@��׷s@�:�ljǍ8�	B9�x�� o���׋ ����9(���G�󍛱ym���\c���U׌�ynI��:3Y[͒�p�srX���7N�6���6
?[s�@z8��R�9h	q��*U��������Y�h��"��\BQ	J��v��מŀnֹ�n٠^�d��%����>��r�75��Fmf6�.�r�.��7i ����@z8��n��T$28H�ؘ�Z���G <�T�}�Zɵ��t��sn 5C��W\q�v����f�n��X�m��a4q�S:02�]���*�m�����"���njY\�nP�7L�E&h[w4�ڴ��/n��tDljǍ�,�s4�k���O����K��Ѐ!+�@6(�EM"�^��ٹ'��=7!�J��	&<X�'�w��@����>�S@��@��J����*�wPT������5����?����޽q�,q�4���,ړ�r\�Jn��R�g�y��9�ڳ\����Ht� d��;��G ;zLxՂ�$mD����تۊ���G <��~����t�ݩi�����/n��,���ت��:đ���&�@��ٹ'>�vnI�~�۹8= W�gu��M�/i��q2��y�� �ۖ�<��G #wp��ݧ��wOl�8��3�<Yn44�cZ3^�V��]�5��Ɨ3<-��rǷ- y���*��a�� '�X�\�I� m����/n��{w4��V�WjU5"�#����*@y�� �ۖ�=�j�  ��c�1c���>�n��ت���4^���y�j�E�D�e��n�Ƿ- {��G =�,�.g��{1� ��I2G�H�Ѻ�,i7u��V����;fz7R��\�.���K�q����q�۵���GmŶD�fT��}M[�#="�v�D�$�f\�I�u�y�{���.�a'�r�u�@Î�̼�����}VG(`�t[	��Պ8��W�Ǝ�c�6�n�ޞr�m��=��\�=�������ٲ�b�uLYW�b�pg=WTܵ��n���x1#A)�ܹ�a�75��M�����rm�	�n��î]�0�=�H�u"nv5F(9�I�86&Ӎh;}4�n恾׋�G���N wuQ<2+SV���^�=T�|��fZ �sWٟ�<����n8�q��/o�4[+Zy#������nh�DFƬxۂ�'��r�Z��l�>�;^��ҬF�"rcňq� ����<��_��� �v�p�v���Xb]���:�N9�͘�`�V�5pWh{&N�M��"lsA	B3dl��r*@u��6e�t���ޔH;.�U�)U7V�O��2 ��D����)%	 ]�� ������:!(����ʧ���sd�SaWu�?�߲��M@yȩ�6캷5���$ЛN5��@�-��9�)�s�V�޶��x�x���q�@>�R�l͗h�M@Hg�����v�ѱ�jx;f�B݇jU^��õ�`^�].ʞ����{,��6��`��l�@�jt���b��	8�4�*Z�[4�w4r�h�jo�H��&j�g =�� ~o��ZJ=�!��*h��$��,Ҕ�&�bYBt�f*�`S�/!��"�C��������1��!NWa�␋(�+(h��b54X�h�\�(Ɗq!��)P0b��J��dR1*�~	�� lsB��dH� �f~h@&�7.� #"��8j럿~��w���T��)
Ⴡ5�]k��5�g�[�A>L�:�a"_��L��	Xhf��q��it�8H�@8;Q]~>6&���t*h
h"mQ����`#��*"�V�$�1	��5�f�v�p�ԪjFӎcNrI�^[��s�S@�����@�z�	&83����se� �P�T�~w{���n?���4ۤ��m/Wiͻy���R�qٺ�hZ�;f��w=�����X��I�A�����Z�[4�w=����留�k��I"6�Z�[7�������x�/l�h�m���9���@�v�����- �-�QK\xG�q���;��䒅;��`��L ����	HB�(P���t����݊���L��ـ=o$�:BS���^��9�)�[��I�<a��M��s`�j.�byc6x�)�g6�v3vڤ���K��Ȝ�r#@9�f�x�Z9e4�*ZU�U5#i�1��������&Oo_>���{\�;ެ���I�#X�nE�}�)�=v�p��M�׀v�t��&�]�1d�1��p�/l�h9�4��hr�h�X�cX��CB��K@;���Iht� �.�
���  �F�CC4��j 8A֑�B��N�M�j�f:ֲ��`)���a.��������ld���;nwTtpvډ�FLѸ}=���<��q�n���\V��d���v'��3�q���\��f�m[�$$��h'��Y�O+[��,��oNӓ�J���n�a	�vK����эQ�N䓶t�o�r���U=p�z:�n��m����w0�z�\Z���vyڝ,߾����"�Аs��]B���	Y������Cqڵ�FTI].��[�c��&��Nz��}�)�w�T���QK\xF���r-�6�˴��=2K@w2�l,�6�JE!�w�T����ڴ�e4^��#T�9$ܙ������׀{��p����U�UDӎcn&9$�9]�@����{aV�}�٠Uڱ��?�'n�J/ ��{u�\]��U�⎈��T<�A��	�I�#X��"�>�n恺�s�{]�D$�������OALY#Lj8�����n,��?<�Y����sڀ�Z��on�&��XۈhX�"���4Wj���?~Ĺ����C�@��	���<��u7w��	K}�`�ذ7ng >���umQ�`��8�C@����I�� {���@u��~��,/FYy�7	�=���e����ta�d6�G���7>IM!��ۂ�(���r�fp�k�|휡(���,��O�H���	7���7��?~�ċ�|`�ذ7c���N��'*���$��LnI�[��@����_a��7����"�:5�1$�B�\B�u�8����ʰ�j��Z��*���k���������S@�u��<Y �j8����f }�w�n�f����:"���_�+���ܚ�v7n��l��n/<��'���Nչ�hE��;4��ñ�٧�9ϵ �� =�*@t��@K�I���<�8�RM�����ؑ�}� ��|`��yСDɮ�:��-�nGBHh����rS@>�l�;�)�w�!��,�9�ħ{�q��׀n�f��j�Xj�D�P5�4�b�=���l�-��jr' �ć��;f��� =�*@IX�<̰s2�K�8���=�{bݗ�j4'�ڻF��H�ӬM�r=��9�И3	&I��y18�ܓ@�����H	)���@G.�,%n�������n�s��S� s�������V	���Q�&h��0�k�9(Q=���=��`S烱��p�8h�����>��X�(�������UjKEU�������ـr�������I9����<RR�BE��Zy=n�f�����8��k��N�{:�5���
��R�=f�%�;��׿�}��|R^tf��7Eu��Y�ȓ�k�^�U�r�l�F��e-�b�8�����Aۍ��C�h &D��P��t�=On���ܠ��'��؃nܷY�76����O1s��v&��Y�<��sX�s��7)٧�x��I�^�ch�������.��޺��ǻ�߾���n�v�i.�����Ḏq#�y�� ���ȩ��ۀ�a�@v��%���
����f��߿����0�k����|`�,���1��QG3@�;)�q�@H�s��2�V
�v�j������ {���`��8�%=��Wh��G����4{)�z��@IO`�=�j9u�a+7v��.��st@z��@IO`�<�����;nW�[r4�$�1G���� �əը27l9:K[2kj���nnu��y�ˊ����Q�Ǡ[�����4{)�|���g��k"�������x�(����0Kn���3�X��|��c���sqɠ{�x�=q�@IO`�9�V��̢����Ywf��u�6�ـ�w��#���]�w�K#g��pX%����`�]�� �x%/fw��M�/ki77n���ɹG^79�a���UM��t��\�:w=�Ӊ�V�c�z�> ��x{l���_H5����,�&FFɍ��$�x�@���M ��h�.9&Llŗsv`�� mm����P"D (|BUEؘ�nM}�����9��{��`���)��4s��s�����5��K�{u���4��G ���=��/�=��[�S@�^,�s#Pc�1�
b��O\q{�����-vnh���Kʅ�8�es"r�s��7�h�V�^v��v� ��r�����RH�	�@����Z ��$�-}WgO���<M�`�Mɠ{���@/;f�k�h�l�-�������uf ?k��np�]�r�|)?g��{���U�.8FFɍ�Ȥ��%�	�jJ�9�@:�����sV��ϓ		�n��'�;^�ùe���Tݵ�vi���1��W\����p�]��l��w�"/�;����o��Ʀ�,S#rh���٠Z�Zy�4��	�QG��4��)�^v��j��=��{������X݄X��&�rMܒ��5&b ��L�SCx&����@/;f�n;V�^w��'{���Iӈ�bӛ$$>+	�JȐ�K��� H!��K| Q>�,f�I#����"&(�hX��T>�:�[��XpB@7
YhnU��D���ZWL@�M@�k�S *�Ӥ
�aXFk%U8�G��j������	Qm���U�ڲ���c���` ����SJ�Jİ���ݽݽ�����VU�U<�Bڶ�8[\�6��g��)qh�Wh�5S�D����0K�a���h��RT�a���7&������ecl��ۮۨ{ks�n1�pt�u<[;�c�N'GQ���[ um�U<��\�n�I�l�r�WO��#��.N�@��:g��R�#�Fl��Ypl�&�pᖸ�(jT1�)�c���SO+]AuQ����T��v��F�@mch8���۱���rv\F�7ҕ�KE�.���A��Ӻ��On��mvv�9Zd�h6bMdv�֫�In��
�yd��d���o��z��g�1�1tC[�fwfT��B��L��]pr�:�W�Ɲ��A`���..�6�^&t����BQ9K�V��ݻN@ *���� �Z5�=&MF����K��<�(ⵒ\�.�mקI�Clc���Mv�zv�NK�ܩY�ѣ3��q��+���!�]�Y��UV69c�L�cF���홻v(]l8d�l��n�NwlF�g����[
��H�T��B�;W �9`(=��Æ`S���+�I�asô���Վ{�zy5c�����F��l"=�9]ٳ��5��Q�Ut��vQ%�6�3�n^@�ދv6��"li�̡��Uu&�)�1�3jt���,�Wi\�
�cN��j��+�Ő�9jz`چ�ħ����3��lkU8��:@�t����0��H��p6�Ec�\v馒��M4rb.Dӛ5u�6t�-�	
O\-WN�]7�M�Hǝc<�I�l�ƃ.��Wt�ɞQ�UP�cB6B'��Rt���l����x��[��@]Y�ǜI��iKu��x9�NZ�Y��c"�`�ƽ=jB�/k�7'H�Humxq�v��1*2����[�zin�H�b���`.�q���V�K9哬�ʳ1�
�9���Qn�C��r����q���Wf���w�&�݉�zsu�/39��zB�d:!�m�;lk�N� �#T
�^V�<#�b�� ��	�Oˀ�D Q���V���DG����)���p8	�ʨl�w�{�����R-��v��K�v���jQ^����y^݌o/;����]����K��e��k�.�	��G=��I�1���^M���*Sv�q�"��]Vk�91�r�l�U�nW��m���F�0m�e4L�k�'�z��Z�[���_q���`ڐ�:��Ox����F���ue�֝D��%��Ų@��]f	����Ųpl�n�r�]v(��~��>��?Yz����lq�a�f�a��ss�Eф놽��
u�ڣQ=�:is3���	7%��ڴ�h�V�^v��*���2,)�^v�������T���Jd��%r�.��-U\�swxuwN ?k�:!DBI{������/j�
�8�LxŋwwP�5%d��'9�I5��k�X���pŊdnM�v�ّ<�������� /��sWs���O�Y9�1��͢�h�.��s�Q���g6�lrF�~�!�B<M����H��٠�4�٠[�ՠ}��1���f��]\�k3rI����(H�"#p���U@����78 ��΄�1"���x��������M�v� ��h������8�7$�rh�h�@-�h{3�^���=��H���"Ȧ8hrj nM@ɨ��W&J6+&���㫬����sۮ���2��=�%��Q�y:�Ӣt��U_l�� =n�6��	B�_H�� ����N9�ᄒM ��o�?$or�0�u���΅24�e��m��R������0�w���A! �tD(��)%DJ"��z�����S��qE&���G�{l�^٠����)�}���4�Q8��G*� <���<�����8 ���>����YO「Xd��L�L%�ʹ qxz7`�;8:�2���e��t��V����@ɨҶ95 tsP�h�lqǉ�bBMɠw�%7��DD�s� �}x ���>l�Re�pna�dS4�٠��@/m�yrS@�Z��(���L�I��D����}׀o��`|�%��P�"�!JK"yE|����l%�57j���ܚ{l�;˒�{l�^٠qt��[X��dN<cX����{Nz�l�W(v��ZI��ٮ:y�N۷���U�K���ddnM��)��� ��{l�9����QG���O$x���rQ	L����}׀|�l�>R�[�(�Bk#�M �{f�^�4�D$�L���0�u�N����*��94�٠}i)�u[^�s��@����8�hI�4���ܓ75 9&�.VuԺ���^l�3�N3�f�:�U�s�+�q�U��3�Rs�NL���e�0� ;�W���,v�]�v�p�^E-�ܬ��Z�s�u{q���N�Ԡ��G���g���g��U�F5v�;g8j�X��Wg�+�{��5�����g���],]8m�۶�E�z��s�c2nx�sϷn\��cFݧ@cu���C�ۂ�۝b�^V��\s_����w�w���;���:���
�����^[�8:O0T+ma,"���i�ǮLI���m����}� nj rM@zM�h\��#�&�iI�s������ޚ=輴�k�~H��D,��xa���?���ۖ��b ��9��^�Ʀ���$���V��u� {u�(�2���R�+�����hln5��{^�s��@;�f���U��Z'�EHs�ɂ]@鳚5��_;E��v�mv�TIG]qfm�/8rbQ8�#������w�S@�ت��٠s+:V�'�n8�	���و���Q4k˜� {����4w�F�d�,m�P$��>�V����%2y�������]Q���8��'k@/{f��{)�^YM�ek@�5dr$�L�I�y������fZ }&�:�]d���-��zx�iS��Ή˫ a����s�cآ9'&芒�v�f��Z�����ٖ�I�UW�:M�@w-�=ōL'�9���րw�j��T���ɦuy��UWWS��� �vـ�!	(�
PD/B��)a4���5�u8�.��&A(�B����즁�۹�}lUhy+�zh���6�<x�q��f� :8��6��j���@a\�	cSSX��b���q�VաM\��0mۑ�d�/���U�ƞuZ�Q6"���w.p|���x�G������^oTȠ�"F'�@;�u��H�*@zM�h��ᗷ�G����4w�s@��s@��ՠ��@����q�1ǆF����X�s�u��x��0��+\��̄�U~X^�ՊUM��Փfn�m 'M�h75��H	�*Fߞ���������մ��d�1\�Sl���:�5źw=]\����mv`���u]��&�Cbq�� ���;۹�^[��^X��;�Q[	D�X$��9��9�H	2��9�_~�Wdf+�<N8�L�=���֭zy�4�w4w�F��i�&�`ԷX ���m���	B���M���[E��4�Ȓq��l�9�w���׀4��f��*+��q��\vv�4!>����>�lx��=P��hAw���:�.���aƺ��n']���m]�^,��Ƀvz�Q�㥀��ک����ڹukGg4�K��v�`��c-s�í��)�I�^�
���@�9ݸ� >n/H\C'�/'�Ӯ�藄9�)ݴ��H��묛���9��F���r�́����ͱV-����[��3Z�5� :	�2e9��B��[�gv��v^�jv���u�@�nK��m�&(���K]�ٍ	��hHt���~~�?>�9�@J�%�	�j�^�ur���E�4�h+�h�l�-�s@�[q�(��xԒM��- F�$�R �&�:��0��4ӑ�"qh׶h۹��@�]�@��E�	D�%�4	$T�9�	S$���6��Y���,Q۷�w�;��=O��u\��\��;--���v���6��c6��K	�{r�ǳU�}���� �<�mR��y5%U��SJl����t��DD%�B��B���P�x� ��f o��֪�Ǒdn(�bN- �-��S@9�٠\�ՠuZ��$d� �LnI�[e4����Z�s���9|���1ǆF�� �5�ܺ���ou��� ���mUQ�V�g`��F:.�:��<�u��7]J�7Yr^��xnn�]�C�5�:np�7xm���@�}x�w���4�DbȜZ�-���h9�4�ڴ�TV��$G1��sWxm��{]��q	�5|���ifTO���T����:,l�:T^ t�d�)j�"B����8M
�(��"R-���F�ύ����)�	D��x c���A� D�a���^�'y��꤀�1�I��6w��,{�B@�
ĪB|��?vBN�����!uU%�%e!	v���Mp�8�
�%P��Ν� N����b����T\� �t޿X)&��"5!HX������~����w�j�#�p#!>?m�S��솳k	~�B&�e|/f�8��#��@�T9U���D8#�*���D(�-P��A�@H�YD@�H�_����P�Ӣ�� |ۼ|VӚ�M�������$�)��� �+�p��:����s|NR�����)<QI�\�ՠ^٠[e4��j]TlBh�F`)� �/��C�x�痦��x�Z��l�meu�c�s��$��q6�lV�j� >z� m�0}��!(�߾A�����U��$d�22&9$�v� �k���� ���S'���b�JL��2� ���U[4��4�)�_��{��`��Ǌ]]�\�x��x�l��$�)B�IQh�� ����h	*�h
)�$���7$�^���CY+NEH#�@>��@��hy�4
�l�=��Y|�I�m��p�뎹ގ���q5�<�u� �;���v�;q;0�-�"I71��m����4�����K���xiN�jQ*��j��*j� ��y�BI)�����wu�l��y�-n9$q�1�rh:��M@G6�5��e��ܫR$(dBqh-�@�l��w���v���YXH�2ddLqɠw�`��P�%��j�y��׳����|}���xۓ��ð�c�8+k�C�VәE��&M���'X����6#P��-i�]<¹�z_%ڇq��=UV�m����fRB�tma�X�Ks���<�v-����uo]c�\���:�\�d���c^�P��1�x��p�r�3dYn9{v����&-�)l���ݓ������,rk&m�f�{/fѻm�*�g'E���w�ߝ��N��4��:�� !6	���n�]Op��M�<n��v�r���Ƙ{HWK۴Ym��~~o^ ��s�m��9��tor�T��<lq�I�\�h-�@�����7߿bE�n��c�D�Ȟ� }��#� ܚ���K@:�v�f$G1�2b�I�^�M �m�λV�r�4����	�6�q~��rjS�- t�P͂�\��k �E�	C�6Ǔ��лl��V,ra��'ۍu:�r��q[��[Jك7cp���@Fd���Z��@�4�Ui��H���qh�տ~S�D� D**�A�6n� 6�%<���.��f�Ln$�n-��h{l�;�ڴWj�>�S��ȟ� �p��٠v�ՠr�V�m��.p��Ʀ��ɠw+�hWj�;l��n��$��[=�X���&���nNyg̛�ۛG1	�ճ����=�gk�������8��&�D��y��@�����]�@�*[����MI�7wv�M����	S$��Ih��ѠX�&�q~����נ\���m�!��z��PM�fg�-~��;�{s@����8���w��O��IhI :ۘ�������IC&$��>�h������/��o� յ�p)ݦ�.��W�G�q��E�:Zgm�e�7�́u��,���x��4v�j�t,�������H�� 1�@y䖀���]\��x$�f���נw��Z�v��۹�\�nn,J`�8�cqǠ6c����-�"�[s��FXc��rF�PN-�ՠ}�w4��w[��@X(0��!� ()Dt���Y��w$�~�i����[[��h9 =m�@6c�����h���Ĭ�$�,2G��u����tiC���;`��ۃu�gk3��e�ά�]g�36��Kݤ����r�x����9}��ݧ��&�j�����:� �k\�kx��u�tD(Jd�����Ģ�(dBqh��hv�H�l�- ���Vi����M�"�����}�{}4�_j�>��hv���Gb������h����s�|�ŀz"!X�IF�������^nk��I{^�S:�.�n{��Ԭ�l=�m������^^�ZI.#�'�ɱť�&ff�m�\��T��gu������p�5�G��[����;H2�e���������mč��(�D���˲� F`����]��Pu�u[�m�:t� v��և�1۵>g�;m�=�����k�8�{ۄz��C�[W+���{���w{������n>Jq���y�i^��9�x��h�6�;���<�\�{�v�n�{f��ˊ<jI&���hWڴ����v��W����maz���t���5*ۘ�up�����2d�Š^[���l�..����V�s�����/�I��9�	V���9h	�*@Nd-f�5!�b	$��.�=I%����J��]�l���������!4�a���/Հ,UЪ��kq&�=��X���8𣴱g�&,Ԙ"�v?���|��$�n�jI%�v�f~�K���5$�~�,�8Lq�O"n9�$�{wCOٵ�E۔�H#F �T��.P�B;��[o>���-���5ۛ���;W�$�-S�Gb����ԒK��}�IU�ꚒK�v��I.����Y�<J`�8�Ƥr}�IU�ꚒK�v��I.��]��Ib�A܍A�nF�Dn)�$�/lߒK��pԒK��}�IW��z�IS�h�);KIg� DXw\�gW�}��Ψy�%�@J!sWةN6��N�O\S_��
�M�RI.����%_c��I.;kߒK��J4	�!�����$�{l�䒫��5$����Iw�t5$��J/�m�'#G'�$�]���$���]&�� Њâ�.���{�i$����K��G�4%IC�ME5$����Iw�t5$��m�|�E�UMI%�mǉ�Lq�R&�q��Iw�t5$��m�|�E�UMI%�m|�_�����S���s�gP�4��i����vkvL8:�5W=�@u�]v�u��qfgm���|�I[�O�I"�*���㶿�I.����Y�<J`�8�Ƥr}�I�U5$����Iw�t5$��m�|�K;���xۉ��5Ԓ\v���%�˨ԒK��}�IU�ꚒK��ۍ�ln5L�H��%�ٙ��;w�#U�����r�{~�v��F@	B()b�$TI���{�r�jgf�?�n(�E jI%��>�$��uMI%�m|�]캍I%�sA��E�=�r4���z6M��h�Q!�2 nܼ�v��s���L�Z�N6��~�?����$���K��Q�߿|�I[�O�I+|�{#I(�J�SRIq�_�{3?fcm[=�ԒJ�z}�IU�ꚒK���c�ƤB�4���K��Q�$�{l�䒫��5$����Ir�0X�$��� �%����o�>�$��~�RIq�_�$�z��ԒW9�?��S��5#��J��cԒS߳;���z�Uze�m����r��_��_�AW�aV� *�� ���Ȃ�����H�����
���H��B�*��
�b�A �@H*�� E��  �DH*AF
�A��D��X*��*
��� �@H�
� �� �������� �F*�`*��
�X***V*�@`�@ �DA �AE��B
�P
�E"�@
���`�D
�@`�A
�P��H*Q �EX**`�D *"�@ �D��
�*��H�� �F� �F
�*��@��
�
�� �E �@R*�@�
�A�� *��� �H� *
��"�
�
�X*��T �E ��@ `�@ H*����
� *F
���@*R�`�E
�  �@X��`�E ��AP��P��AA"**@X
�PP��@ *�
�H
�*E��DB"�*
�F� �@"�X
� 
� B���DUH*P�@ *E`*�D`*Q"@T��������"
��_�
��_����
�� *�� ���Ȃ��B
��� *��_��PVI��C�H �	�` �����_w���5� $  ���
 ,�` �r t      ��  >��((UP+f@�	P�}ۈ�R����Cf�tb%*��+�*�� �J�v ����(P�	 R��    	� �  ��kǰ�� �{����rx�Us�(�R+'����]j�wEz���z���U����ז'��  <�.{��`G����;S�=�>��}��z����n��4�wS����OO�a� }�� >�   Y�A���^�	�}���v�{tx�����Ԇ���y�W��T�u�t���<��n� �g��À b����Ϯ|�����]5z���aN8�7[��`{ͧ!�;���hp�� }�C@�� ��zl���L@ <���R�6P ��y��OA�� ��: s��4Qu���@�� w���c@ ���R�{�@���or��(�n�(M ��`�()K,�����J���@�Y�� p  w�S��� x@�[opR�s��;.Z���靽R��	�=�۶��\Ý���Ɔ���i�s��v� {��zs�� z<:7wz{��ݏ6�w��y�/�>۾���!Ȧ�v� ����(  4}: sǸ ���w3��ŧ!��rn���=7��t��!�`鹁�����4}��6=�� �	��a�`zo�_`��t�̓������ �nͯ0w�w�vN��A�   ��"6�%J&@ ���R��b	����U*J��U4  ���UޕJ�  ���R�ڊ�  �A1J���OMN"���8����,���gq��q����@^�q�TUȈ�*��TU�!PW���*�AN��@����H�ą� B��ae
o���l1ɰ@��/�9{v������nl	�ݼv8�
%��P�$�I#BXK�j�Y��k�� }�a��q��`DM�Iq���o������D�B��.2����7��`���h�r|0��c�}s���Co�(J���0.�r�t�䄦!\2��n�@ѣ�e75�@N��p�d"D�"����Ӷ٘�ǗFrX�Y�')�&_$�Jg�o�����8b&L�.Sq0�J5O�k��P���|��}����+�C�9t�۫>����'WH�⨯��# �6��)$��B\��8p3L5��3D��!L�1�LbFx�Y���y$�5���1�E
�>�%�h��٠���9������ �)�a�����.�&���&H�b�0�U%�b��hP��2I	 ���Se�-r,@�E+�d�&):Ӽ}��d`�"EpD��Xi��.	Lo�H#a���|u�� ���466�g��.���@h����4i�>��r����yW��v��:yw���U��BN�>R�������>0��:�1��ts��Ȓ�ֱ̳���B�9$��`��O���B%9�g���>�0ˍc��� Ŕ�?6Nc��ɢ�;- g�*!$L|ﻘ�>�����w�	���%�"�q�K����
C�r��L]0(c.�#�0dӸ��4�fG&�fMn���2:"Cn�4��H,*�MHP��R�c.�\1����s�h����9��5��Lsr�v���.>53��>aC];XBɭ�$��901�fK��D�¤1�a��r$3
m�	�O��skx����9�9�xrF�$�XF�0n4cd#cC�$�"i���a��!��ِ��M=MָL�,��e)�[��8��
Ƈ�.a$�R�䅟=��Hi�sB�)��K�S:љ�:8�Nd��P���a�CK%�Âd���{+��Ro�ί�ĹƸ�3
B�F� @�B8>�P�Ŭd�LMq��L�� %�.C&��
ă���A��.�1��X�XBZF�%���I H�%RP�%RT��%`B��r[B����r�6�^_a4�t.���3,)<��������OFg��4�fbF� E�\�k$eR��BXK��9e0a�	\g5��&�qX��H�@�d`HB$!$�j�O���$�CN�G����	��s�O�B>2h�uѬ��)��4�����ђ.�'���.v}w���5��!B+
��)%%�1&�7��;�`Llxd���6�a0X�H!�[�I!�)G��	���L�^rs��s�K,��F�$<�da�ޏ���(H�B��>3ώ�j�Mkiri�7��a@���HRHY%�&�φ4pd��썀�5�H��$��@�'7����Z���B�C%�}��M��q�bg2k)�B&�-�����c{��gG�H��P�F%�R�HH�0~8sn�1RH0"A�h�D��Zd�H�d1�Rl�%e΋�Ԅ4��R]k��CxK	�Y�I�\�XK�\��r���)�6�x�(�NWu�K�)��h�	C��޾s��-3�n]1�K��I��-��$�	BZ�����xbrF�,��a�%�<�%���d&��r�r��]�k�6o�'�MC���F^�~��M�3�ߵ�x�q�k�L�(R C�19�:�B�)�^=�Ri�bU�@��\�Y�[8k7V��H�������HXXȰT�BYrkr�2k�A.3���~���S5���C[�ۆ͟oY&;�"c/�Lii��ć02A�e��3��8��0$5�Ns7>ZsA���fB4da�e�l�9m��]E������ΦL�o�����]f�:H��"�)�!)��P�9�]��ξ&��9���kن\K�Ћ!!aHY�S�:��s�3��t:�훝�2`��ǎ.�ܦ���	!$a�� ĉE�@�����.(C4��1�Lfl��a�}���ɑ�#L�d�BX�ZDkWmY$ąk�5��Ÿ&�]�.MF.)9	I7��g	XHrCj�-!���Y�B��5#*k_&q5�iݹ��9	4�F�&�y��$G��3L$�2HB4�%�IJ�a�!un4K�E%i^kX�&�}ʿ�v���k�\����+�Ru�.NgWf�\U;�9����Qx�0��̪����3��oӵ!q�R d�w�˽`ԛ�ɼ�7v_���u��_C�HI3�ƘBalZ`�ˎ��e�q�m�ą�)#��1�|Q�	0���0X�p�гN.�H�
`!K���4F�%�4�j�F4k_u�XP��HX�$0c,,�+����LB�ro�N��{�5���m�>4FBB�r�bR���J:62��MM��	�Bf�#'�V0��w)!w�+/��w�r����[~w�8s{�>YL�ن�kc�N�v`�0햘��1�o?}�!i����s}�K�Lo:���!�F$�s�\��3:�!��
4p�H�v�������~��\��!ec�HД�X�H�DR�2^� B�k��`�a$HS5��c�� F`�������MD%���a���d� ��U8d!����pd��cy��I!%5��M}�P ѥ6� �a�c[Loyƶd�w��Z�0�b$@cE�P�}��cO��sNsTx��H�$h�"�*�+"XC1��S���W)�hۭ�Y�j�����`HH/8V�#"��B22���a�"@�@��S:�}�H`�i����N�*I0,i�HF�h���έ��Y�I��gDz�vƸL�E`�Ĭ���#L-kH�e2')��Mgw{�B��aP�aa$c��p�(8c !bE�K���T��d[���E�H@#p��HҜ#FXF�F�i������(�
s����8�`� 4^.����P�41������c_7�k�2kF��m2M��%Q�
b�u��7>�t�	u��|H��1s���o��~��3Yno�|�*�Ö1�!
��"�0�B��
�8l:�4u�	��t�$ �6$2B��$���$,�� @��(|20��n���N>֔��"I$���C�� ��ζ`ѽ�8�M�5�~���I �#%�2�d�I��4h��F�5���HƱ ��
E.	pB�@�_����)񟏈�!L95���k�k���g,�ɭcP&
������Y!m�q5�����L��i.7�n��k�h٣��61ZY��CA,�L��27��K��Y���!X�d"�1�%�\�c��� j��+�����W&n�̡�8f�kd�a�>��78����g�\�œ�|f�%f�`ocr��5�\|m�B��2�H#R0g$��)�¸2�<;
b2��%�ε�Q�Nk�~>Zg�)��bGk	 Ʋ��	��,��,%c!r�gO�O�Od)�,�(JFJE�R�B��
���	3��l+3�a��m��Ƴ�����%�}�$�8}*� ��7�(GζK�O�4#Na��.2h�&e1�CF� ��$ � � �`�ӦЖÐ4;#SE��h�1˞}f��pff�O���O�H���X[���R f@�c$"��8�4d�`b��a2��>ќ�h3K�i"B0�,2iə��I�K�k�`!HЅ8HP�3�}��>�Mѩ�C&Lˌg!�̚�X4���w��Q]��_w��M][�|�:(�n�L��`4�(I.^��2������e%����	n.��p�`A}�w����^w)W~���s�.�EQ
<�$HIIqܲ��N���p�4`�Md�A��U�B�Υѩ�u���o[{�BHfva�;��B���aHR�"��!JI
ՊR@��Be`W� D ��A���0B4�BK#����4k)�%�4i��ư�35����w\&�ⱄ���&Vp��S��IJB0� B��	`F���Z�}���i�LщLo�b�@�;C"D��3�s%��Ll%�a SX\6|����HCA
���ѓ ���MjH��4��.CG��L�ܸ.�4S2h`!fl����2w��1�t(���%X�81 ��l���.9�.!&5���G��a~
�`���cZѳ�ۍ���}�nH_�oD!X��Q6A�aLആ#aV5#!���eIRRT��b�r�:���a HYI����3�s�]! �m%�Y� y�va.��S��]ӏ����Z     l �m    	 �\   m��� �  6�     @$�     ��h MSb�5��:���AA� ����l�M�˲�Q���[k�$�h���۰��y�7�W3� %[skj�l��]Y�h�h X�` 6��6�Oٶkn� ��PR�T��e᧭//&ųr�E�m�j�,lt���/�l�9�@� 8���	� 
�%e�(���1�Um��6��lXa'-�m��;Nu,FLÀm[�/A�5�K���M�6Zm l �     m���,��,���m 	$-�j{i�j��I]�Ѹ��n^]�^����v��t�`�^�{GY�q�X
U�ӻp��.15]<�1(!]��BG�+c$QWT��4i�U��E�Wem��d�%�I�v�m	&����2a�t�Uyi�
���۶ۉ��]� �[�vp-��e��
��xOp���[WCT��P�X ��nBK�kJ[�a%� -�B�n	,][m� �K�>��>�� �@z�j ]C��0�k��h��V�md̀�����~��<sL��lj���p�"F�CeP
�R�<��, $H��^�p��l-�ݶ 6�vp�� m��[''Ss��[ov� �C��E�f�pkn��p-�A�����.k�=����m�5�uU�J�@J��-�S��ge����ض���1�]k�T6��o0rq<��t[q�������u@FEv.��(� F4������8uY���R�J�0[V��ե��Kt6%��>9�}�@),򡫉(�ڪ]b���v쌖�@)�:�c.f��ɸ���5�J�F��kj�Vf����[���V��5.0��)��n۰���H�>/Z��-�դ���p��9�c�*�HJǜˢރ�q�       ���aĀ  �bR� i� �m&[\з�X֭��������@ -�[RH"@6�e*u��*���UY��V����UV�#;
T��   � ��MȬ�2����[R  kRi}�}�}m�Ŵ�����õ��!:녎��V��Ij�À �]U
�J�Uq*�mm���-�ٶ �H[kF� ԒK�.�a��ge�U���,� �j$!�ye��ݵ,q�!ϛ@��oc\�X�vԆw5�AUFB�A��B�Ŭ��+�C�Zl%� q�7n���]l�-Sv�[)�$��ku��(
6�& �mp�eM��sH0�i6�*��@]���ݺPAej�eڪ����6����R��y�ĵU@�i��I�m�j�i����Z`##�VҨ9�Z���0�jh6*������e.8���c����:y�Gj��L�9�v�Hm����ޒ�6��H�����U�
�\3%K�VQ�t��H�f�%��l	$ e��Ą�l=&՛j�	�R V� ��E��d����^����
� \�mr�b�8��m�ɘ��=���C��d6X�.��MȜZ��Y^��p^�`���m�����3�*�)�v�,�RS�kV1��;;%��� mT6����^���\v�U�mk��6���`p� �&׫�ä%9V�9�����;.��m���vT

���j��OUR�H��t�t��f����Utt�mP��Jm�$�cZ;���m��Pz,�Wm�U�q/+M��l�	  pݻkjN�H��!��M,� [Iμ6 �;K��H���ҳj�H-W���Ts�3��8�����j6���ڶ�����l�w]�l4�a!�JZM*Ú��+]��"����@6�vͶ� ��f��()j�P"�$��yT �L]�UuU�倨Z�j�T������ � m���ݰh��8�̌ �#mw)m�M��    [���m�   �` $m���Ĭ�*�J�U[T�R��,����-J�D��PE��[[@;i6�� �@��4�9�δ�����Z@m��H�	 $��m�Ǎ��m�  $y���  m4ڀ�i��Ę6���0����;Z�J.o�I���Jb�2��kF+q�4��z�I���t�1��T�6y-��g@p�l�A���-5����� 2%��K!z�-i����N��� �[m��/�Y:j-� %����YN����Wm���+����e����hGR�V��km�G�ts�-6[M���m[@ �&�퍶Xs[�L�*�MuR�AR���vE��^���휑�^�%�m��`[d��
� H�� �  -�Y/q!�hl  [[ls�`Q�4���`m��` h ��](����;nJ����IK^0G=�+��*q�'5mm��$7m�i�Β0 *��!&X)	"Y�dK/�F���p=�UP!]�Z�lK��}��)���  m[m��ӛf�-�n� jEj��N:7h�R�*ʵ[Kv�)S�iI4�n��h�am���Hӝm�  � �	uqOw@ ��W��6*yS�_k�륋H��k�q�yM��Z�x���j��j�I	5{i�m�z�W*����g��:)��v��c���j���>
kڶ��	m�l,K�5��+ͻ�SX;g��Q�fGe$+l��(�X�m� m��%�^����pɷ=�K-�d-5-�颏;-@�=�=����Z�eg+��� ��[�M���6��V\�m�� :��^��f�(� m�nNh�&s��4IN�V�W ��M�W��b�[l2 e��p�	  �M�����H���ɵti��sv׮��m� 6�6�C���im 
Z*��UR��S�8`{s`��n�H y��m�� $m�	)T
�J�n�8Dk.�mI-�lx� 25A�T���m*�P&�mJ��bǂ����T6�d<䪨wl����lv�^�Џoe���+���Ry�2����#UUP�ʗ��lښ�1 �t�2��g�؛-���ZU�(�v�Z��j��6� ��٦���ZUUUT����*WK5�3{V���d  $[o����I��#�� �l�m�j�6�������m�� K�ϒw�mA�����vºv�
�ҥ�i�ٶ�@n܇n��`B۴�с v��`,3\�l[M�T�8�h��
UVT6�Ֆ���,�v ��n [m�*va��Ҥ�#Z� D��v�  ��v�a������V�mm%�`P�)����m[���t����`A���ͅx:��R�5@T�%c]���<�}�;)XV0�{XvT9iW��������*�.��t� ��ߍw�ޓ\ʰ�[AY3؛v9�u�&3�iѵ�,����jHu��U�
qmWn]���厭�ڦ3��EE�#s�vۑT�n�3�-�)2p6�&�    �`�m6�n�L�ݢ� Vl�IW6�@ U�mٶ $   5�          ��l    �� � �`   a�   6�]m� 6ؑ�� ����o`�cvٶE ���K5H�VF �m�  ��     �A��m� 2 �ImD��l�y8Z���P��*�[O8�f�d5���d�X;j�&�{$x�mͭ�B@p�^���i��[�}z�3����nV���:YRkH��&�ym�m�Z����s$�YF����U�[m&�^� ��&r���]��\ ��\�:�
�6����j�@�aݠ 
&��xRN������@9�6�@A��B�x��l�AJ�hN��nX-�G/l�쀤�̳�n�[x��kVv�^֛ $X֪k;U�mm�pI(��K��޾��(ym:WC��UUP�U�iVBg;G^+��n+�  87^�7r�Ŷ�u��Sk�E�n�l��b�<�UV�]{�H=/:����� �m�p6� []a�Iڶ8�a��I'` �`�z�� ׌Z$u�d��]X�sV��ݢR�b�+�@�@[��f�t蓝  dH����q� m��m��e�kכ�E��h�m��f�zѶ� QP
�m���iv^��I(�	��!&����[;f��m��4� 7Z�>�o�{/�mKZ�	p�����6�b�Rsj�N��['U�  �K*t��� �mץ]#�Re� E�V�f�Ӗ��qR��R�WW(+�K+mJ��U@u*�����-sFP[n�v����bƖ� ��m�[m�m3+m��Im=m�N���E��5�t�s�m6��j��M���jMm�]/8��!��-+m���� 	�  m  ��m�tŵ;m��� ��j�m!AԐN�-[�6N-'H�3Y��$��Mn�)w]���u��V�����.2-�
A� nj��'\�v�'hy���=%*��ٻl���w��������T�GH
Q
�ȧ�!�G�@�'ʙHej�U�L��+�x��p��:)�2H"Ev�T5��hpC�_�r�� +�
UG'@��@��Di�P�Ca� �A��H ��Q8�h04�P0A�ЁŠD��!"�E)PMi�.��� zC��"��x!�w��M�q(!�껣�N�`ChAF ���xa8&G��ȃ�
�AC�&@���h |��R *=PC睊��\!<� AP�T4��S����B}HE@È�p���� $I)�����(�|��~T>F 	�u��H�U�u�!$>b�hc  d�C�DS'D_�z����T�^�z�L�P6EC�� �( S DW�
��S���R�� � ���6U6 N�T$1�IR5RBh�KD,bŒ)�D�t.(��AHDI�SbQ:�G�$�XvD~x"��VD*�Q��� � EX��� =T4��E6�&&�i���L�TȜ�"��  N�ʟ Q�t0�=��^qѝ*�BE��"+  H��X�"DX���+�D>^�2&�tb�"�2"��������d6�P|{�����:�b�� ЭZ�   ��P(9ε�s9�lE-����my�-5e�gn�F9��h��Ƣ�i`�ncۣ1X���݂T����:]Z�U�,s�4۶ځ�.�'<�.z]�T�˶��'9�e2�6��Ϩ&�n
�r誫��!�d�5�.����I�vM�e�uL�V��9݌4���Y]g=��{c��=Df�2qng�A�.�N�P��뗣W<���<]
�)���vyQ������*�����![8Z$�a�	i
G@H��.�ֶ��:0Je�N�R��K��:%G���β���{-�ks��tE��r��x`�ΧZ���nL�i��z��;v\ȯ&������&];�F��j�E����PpP	���sp���!�l]�*�r�b9�5M�<&�]X�X���t��˝l�fu�iܛ)��P�u�6i��T���������b!�MU&�L����e�9��S"ʹv��A�،̑Ԏ,"�kua�8=�.��mƊa;	�
M��g,�w�^�u/6�r��v̤˔0a��Tx�eb��
�t�J�p��Z	q�p�Ԯq��#v�[�܁�0���S���b��4�==tn�]h6�c�.AnZ	�vF�y�-�\���mrt �5[I��[6�y܋J�'3���D�,t0s,W��D��#��(�����!���m�Fa닀�E�ٝ����uu��S��
�.���ͺ�U�vx<���T���몓��j�U�c����a	�-�nQH�&=9��B��I�ȱ�[D�u��)j�VUT���k�m��` ( �M�����X^��f� �F� �%.�u���kɡƭ:�S��PݺS����K�;�m-nm�u�f�H1�Q9k�ځ��djL���6��]+�)�Oa�佮l�/<�64nv)��ws9m@���=��K�E�h���0�����s"�q��-��l"�U��o^ jj�uG����in�Gn�=��ޔ�*�L�~S��:] 9�
�D>~mv)�/�E��GB�z&P��1^q�'4�h^u�6��3U��8�ֵ;�ꎉ۰6`�%j{#b�6�D�Lq��8��u�S��v��!�^���v�X/H�|`m�͌b-�4��ҩ�;rgo�#l�6��ˁم,Y���,=<�(�)Ճc;���{t�.Z����ɔ��@v���^c�&^j��-qhC��=�q���A���k�۰���3�����ӌ�f� �࣡ʎ5�b�[�,��{y��83���W�1��;{/d\<p�ɻ;/�����]��E� n�8�����_}�Oe`޶�g�Кm�?�ݼ ���}Il��$���8�ǀȨ�B���:j�ww�j�ǀn���8�ǀqI7lmԺ�- ����2�)��RG�j�ǀj�ԇ-	��Wwn�wX��)#�5wc�7ve`��ﾨ��o������v�t���6�kM</��u�/��J�۫��M��{]TS��v]Zj���{� �ݏ �ٕ�qM� ��X��Zai;��r���[@*�^�	��@��-H%�A�d��+R8�9`L��2�`
 �U��1������6<�H�H:tĨ��颊�v�ݙX���|�W��E�� ����Q6����WwX��)#�5wc�7ve`%��%�M�򻵀qI����+ �{�$�����{��ر0��q��S�j��S9�OV��b�μq�pڴ�^Z����.�MRwk�E�� ����9ŀs\� ��6�]I���Wv��̬��X5Ȱ]����}I�EKꅌ]Ur9������>{����v?�,Z�,T��۾��o��I>�JJ����[������{���ٕ�r=� ��X�h��շk �ݏ ����9ŀs^ŀ�wvl%��.#h6ݪ!x�G\��B��$Z��V]�@
�+��j�Y�
�v�n̬��X5�XǱ`��5J&ۺ��������X5�XǱ`ݙXf�Cd�Bi�WO�wk 潋 ��,=_}IvOe`�y`U؀��%wE:j�v��b�M�ѩ';�v�N '���P�D�E"�c
56��\	��>̼0u�m׮�$��@
�`ݙXǱ`ױ`ŀzh{�J��8�`���v��7<ʡ	�?����Ǩ�N8{]Z@�l(Gl[RU6����~~��kذ�b�_}\A�=��I.���,�G5�r����=���{8�]ۘ�I%��.q$��ˎ���"�V݋Il���I.��F$�����߳�x �n�j�1e�ݮq%�����q�Jz�8�]�pX�?u���@?�bfS
��$�^��$���헞IO\��K�}՚�ۑ�v�5�����BQb�#"Z�H"6>2^�Ű��vl�d���Fl�PĬg�ݮ"A5��<ٹ�L�t�D3�q�Pw:y3�pFXHz�c�<�@v�6�X��$���aZ̵����8�U�5��W]&��UJ��n��vlKt)'6;Q�2����i��p��b�&�&��'nŶ �)Ʒ��(-h��?����\2��Qٸ	�����Dsۨ�mC�o4_�n��������z�SO'U�N��=O#���s���K��K��Q.�Xm�7N���{8�]ۘ�I%��.q$���,��+j@�x ~�������m��~�1$���.q$��q,I%6��u,$��T	��K�s�$�\��I.�� �{��@?����\��%��96��}��������ߞ�_ ��w�e�H��)�.��KIl�8�]ۘ�I%��\�H���?vy�2CeS67FX�\��-Z��qӝ۱q����Z�lXz3�d��>�O���֢d= ;��Ǿ�~{�| ?u�O�9?�������b�K�b��n�m�s=՚��؄8R�1�QK � �$62i�a" � g��\տo;����{n����z{����:����*[M�.$���ys�%ݻ�bI-�"�K�s� w��6�X�al=���rG�3�bI)���8�]ۘ�I%��\�H	����Yh�����������g��$���ys�%ݻ�bI.�G���ܱ���R��\���ѤnEg	�V�3�Ĥ�B�����(iQ%�Nq$��1�KeȹĒ��ı$-�"����U�ڭ�vn�< ?u�W9�m���,I%=~��K��RĒ]��{Y���r����=���罻�ۑ�&^�l�3�躶�߳��} �;���5��C��^���%�s)bI-�"�K�wĒJHѹ�:���S�@?�n� �{��$�u�$��r.q$�wB���]�e�S�U�ۢ|�^��[:�R�A�"AP�#��0l��1
�f-�����^��ԒĒ[.E�$�ݹkI)�Rz�`j��T������9�m��?|{�޿'����I'6�?t��o�Qe֤���?|{�����$�ˑs�%��I.T����`Ո��'����~�'�~~������umޢAY�!��^4�C;��{����IsX�+��� ��s�%ﾭ��K�$�\��IwnZĭ�;��/l��rL���ft�L���*����T�S���}+�(ݢ����豸��� ���< ?�?�{����x {��v��y�^�9@��M�$�����~��������I%����$�vއ����]�^����L���떱$�6d9Ē��ı$�v�.q$���B�e�m&ʞ ������$�����$��ܵ�$�7Dܻ����}����< ?�?�{���q�m��uٽ�m 8��I��<�H�焚O<���8�4f���q�-������w;���,U�4�j��L�-�S.���F�P�r��rƔx���6��d<B�5^n�^�nJ��lz3�^�kM��mm���odөshM�:�\h���⳸66%�����KѻK�m�#�B��O�$�6ާ���� o8�.a6,���&ͷ&ŕ È����3�V�8]٩3�ߤ���l�a3m�P��n3Ѻ����:��<���T��c9�h�I���/��kY(��R!�ߞ�����]�������� ۰���ڰ�Z�	��Ik��$��̇8�[�`�����@?���1ș]���I%͙q$�;�Ŀ}T��s˜I%�;��_ӽ�,3R,e�o��~�,I%ݹ8�K\��$�vd9Ē��W��P0kS�����O} �rq����$�g��8�[�bI.��J4}�`^^�N��:��.�[��9X�y��"�펋�݆2%[�]�T�v��*{���oIsfC�I-���}_WIl�ys���/�X��]����v���[#E#!�h ����Gf�Mf��%ն�w=�����Ψ���v�J7��}��W���]ۑs�$��oIwfC�I%[�T+�iP��IwnE�$��%�I%ݙq$�;�ĒZ�)`]	5
{��w�� ���;}��s�x ~{��@>����W�/�7
%[-6��D@�����.WA�U�V-�9a� ��*���9+�v]���y���Kc�,I%ݹ8�K\��$�)�IN�G5�������Ϲ�m��_�9ĒQ���$�vd9�}T�[��~uc�IZL-4�X��,��Xv�ꪭ���aMʑ��.	�9)�@麚C��+M�t�󷁢*�9P3�"˄�HQ��e]|fɜ�*�#!j@/����cU��'t�N2��O��@�t�E��
(� �.ŋIk8|N��_���s@8��;�k����:�kBS#� 	8+���4��h������!\K�LF,i���/D��4{
�&��(aS��D��V0(T���2��Hi�Nsn��.1cP0�����b�x	���%�v%#0�A/�.±���(@���8�EL�: �-H�B!P��g9�IA2�Q�$���p)�2�6)�&�*�O�ҩ�#�q��D �f� b� �T8(qU�� U4��M��	�D8�b���P�W���9z`�"�5�4��]�XuȰ�`�"��-��,I5H���
��Xv\0�`�"�;�E�{諾=����ګyS;�G"�q��m�KU�[<%�����\0�=F��g%��E��w{� �r,��^�������� �^��T��e�Bv��b��T���� �s� �{��M��(��~�.���hWk ��,G�aꤶ?y`�<����t��r&Wb�[�98}��]I9�{�RN��Ԙ7��@����ʭ�DL15�S�O��������=����XL�Ȳ�o ��w��r�}�������~:���`�K 楯N{r��9�yȃ�Zޫ�{LWK4�2�5av��d�T[����ï��X v�e�6?�XuȰf��;�E�DB6�M��Uv�`�"�RA==x��,cس�K��G���hJݬ �����XǱ`�"�wDܻB�e�E����`=� � I��	[�T'`�J��`=� �_}[/�\ ��� ���;H��:������f�2a��cL�E�D�u��!ck����[y�hy�!Y^�5�䁟1��~v7�E���9ŵ��\�;=�M�<v�N�Zō��	5������E�N����$��6�RxM�s��]p��<�T�m�-˝c:�n�y#&�R����6Mv-s@:6��+CF�=.ND���[[sy��p(Ff��=����9���FG�-l�SW3Je�}^l�\au]#��ջ7�����q z���ӝv���BVZ�+��O9�l���X�b�9�n*Wv�v�;�m��	6^�r,G�`�"�8�RE��\�f�^���o �w������ w���'��tEJ�`\�G�`�"�	6^�r,"��h�+`�Z�0�`�I=|c���.�L���v���n�[w>�خCrѲ���g���y��|V�]7<S�S����+I+���+v�we��"�9%��}_}�q��, ���]�X2�J�ݼ��Y*������]�9|0�`[�窪�#�"��Bv��7o ����7\� �ݏ �)v����.���v7f�r,�v<�lx6\0�+�E�V�ݶ��`[��Sc�9%� ޹�9ϴ��m�K-+JKi��:]�	��`Y�*LC3@��nQһ[l��T4��-u�WI���5{�x$�`�E�j���'��tEmv&��]�>w�N��X�ذ�#�"!h��
�1��uȰ[��}�r�����61�a+��K�`p*P�	���Li�E������I7�p�;�5J$����
��XV�xT���p�7\� $Z�ی�-$����:�� ��U}7��H��uM� ��W^Ƽ��Qv]���Szy�����z��"r��JӞ�R{c+#n�uPM��%v5iRwo�M���7�E�uM���5zy��b���-$%e��n�z�Yꤍ^�x�O<{.��N�ߝ�J�vU��<��>���Sc��UU_RS}~0	��Xڒ��v��ut��x������ �����Ԛ�>)D�J��s@y9�� ��'��wm6.�n����T��� �9�uM� ���W�ޞ����vNn��-����5��7� n��v+q�f5sD-(�������V�,.�����v=� ��.7o�D���R�k �{~��6E���o����7\� &���qЬZ+�XT���K��}�奔G���<��� ���GFU
�jҤ������z�	��X���=_-~�x�X��z�!�j�n� ޹������cRI���ԓ�$�#H�@��I���5;�cW8ɂLf�e������cr�vns�{P�L[qLk�"�����F�9P�kL�)�m=f,-���e��Jf� �V�v"�eZ��w[:��0
���n-f�wnAqQ�5ܑm��G;Mc��y#��u�o����6�Ǧ�q�n]wlz-����]q -��s��@(�A�M #�ړ��<ٲ�s����[n.�I����z�礇&��O����}�{a�U�����VKTv�x�v�\_����ۨ�|p���ɡ�~w���2�s[\�l�@�}�7 ������_����&�y`�)껢�ڷe��j��Sc��_��l7��׀z?ߖ�v<��_RGj3�]ݴ� �i�x�{׀s\�W�_%�x�<�B'�jt*�%k���I�y�o~����<��� �ݏ�UW�UIw�����j��+�����`�c�=U�W�V��> w����"�8��Q�)XXS�� �횽�hZ82���K�L�
0�����f9~䜒M�!�񀔵)��o�y�$��w\��}���I�J�1�k^��Cgym���|��BK9�y(��4Ae� :�r-2椑S��Tab��&�c]O�A�f��v�I�㾺�}y��^TR=Z�R�ة.�[wx��,u�X~������U7�~x��~��[q�T�D��<��I��ǖ��~�yhrIx��[/�XcJz�諻��t�v�������U=����	����7w������.�1]�J2�(����F
�b��f�K#�.�L�J�B���x�<ܻ�i��Wm;���޼��X��}�=-�w﷖��֟b��PP����"��U_��=��� �߿< ���W�%��/!+���	�`9償^w����R"� #kE&O���W�Qf����	��� &���r�[i��+�X������< ���;�E����%�,R��y���������^諭���.�xV����oxy|5�ᢘ���4�3k9�U��p��;b��kw*kqe�,>�$�i���v;N�l~��5nǀul��U�}�^��kΛ�vZV�Rn���,�ԑ�{� ;�z��g���Ɣ�XE[��]Wpo~�� ��z��-���j�� �d��.�]��� sd���,��,	UN��Q�W6A9��)�r��:���z��h��	]�X�+��9ݸ`��襁\��[<��%��ж�f�jU����Α[ۦ&�lv9�Y��ϛ;�]����l��-���F�Ѷ���u�Xv< ��~���WXl��0���&��m�ZI+v�.�xݒ�wnuȰ�\cQ���������/ �v����s�ߖ�{��;���^�e
*We�~�����N<��`���~���W�7��������ʹQ��ng ��{��?I$���Ϸ=��}����2����*��UU��]�ɐ��`"�p� d���rvq!�kF��|̄A���!��$(R,��3+H13���Aý��s �/!m�B��h>4J:ka�7):o� ®9.��3d)me�`K�S3��$Y��,Br����4ʆ�l/��h�cK��ZY� ct��S���9�2k	����.tH���P��4� � ��$ơm{�	C�I
ʤ(BRK7�XrG����~�m�l��IF�[Kh�!�T�
��6���	T�en��&˂@ ���d[j[m��
��hݸ&HcRK���m�6�QH5G�J;��[N��X�s�`�f�r�h��ۍ�Y2O~k�?e���lӋl��<Q�uUO��^�l�3(vH������G��#����9lݴ��quQs�v���:�m�q�f'���[Z��L� ve���� �2���Z�UҫB���kH2�G��*��ȪYh��+v���Ce�E�҈i1�2�b�	[�%��� �ʼ���R)��JZ'��nׄD�����i�U�y���-��^���v�n�����\�(\��n;~-�}����q�M+�Ɣ�l��g���f yu�v�Z��7�*6جY��4�4��6��4<���&KjmU�ᆪ���P)b	�Ygd�
�cr�64N+2�V;SWf�� �������Ih.�&�L+�.)ٝ���6��LD�밃�W9MJ�j�'nm@@7@J���зNń�\ �݄����2<�*J�Q�C��uq����˼۱ԼeTwl+����K�zPuX�E�U#����^U�˹��<�Jn�������S+i䵩"ƍ�������w*˳$���p#�؞��K-��[���5�<��qˆ�����:�댫�Q���a�聈!ևf��ۮ�FD+q�[FhvPY^�Uۭ���Y�/�m�{&YcU���y�+�[�1��q`���s��7��Wl�����ݴ��m�� �m��m�f��
]�o���?|}��]*�m�����|��\\�Wv�(�Ӵ�d��CW-k;t���.ۇ������U
�����'4,;(J�:��"m0m��t�k֪���I�l��u��<�8��h����]�z�;s��2])�����:2�d�\k��䳃Vw2�ZVf��pl]*�S\uB��uNyd�j,�b[��9����1�d�R�`Q��z \��Ct(���~6���"4@���������ɹ'/$��N����!��v\s��հ,���c���|f]I���s2�5VR6*��r�j�L�U�$˜�dr���<Z0����F��q�]\�S��C{�S���8���xmg�U7<F���a��@�z���ț�rko�@�Aj흒��ش]��P�S8��qR�N^(8"úE��ۨݯW:l� ��Vn��xnp�������{��{�����ݏ�n[ns�kh�,��(ջ#k��9O֟�A��q��~B�,"���)���~��~� ��z��ٕ� �����Vv6]�;X͒��}U_��߽�+ �~���b�$�/4RG�Wi5Jһ�z{+ ���oߟ�, �~�x;��T�utZZn��e�,y�, ��x͙X"Z�Դ���i%n��ŀ�/ ٳ+ �ݏ 4��T�kn�͢h�h�4"f���[-�WM�	�h$Ң9Wl:ׁ����ym���\f̬�v?�}��A<� {hP�yK(V����{�{��y7�C�	<��YTP�+Q��^s�ԓ�c�<��w��r�~w�L�
�\���<��b�l��ov�s�-�XE[��]Wp�������=��0=��W�\�x�#�vv6]�;X͒���0���G�`�{m�q �f�h6�,�hm2Gqwb�2��\���6����-��p�fv$�1H��+��7�p�:�c�9�ﾯ����z��7K����hm]�V�y��;�<��޼��������伆��J�m�V���~���%ᵿ*e	QA< �s��jI����|s�S�>[�T���?O$���y&�����7޿�ջ׾�������m���,��)]��|�ވ�y�m��|� sd����tKi]�k6�5»3��<s=��m5ں��\n0s�e�Pt����sy��g "��f�m�'��{ sd�W�U\A�/�մ�ذ�S#4���=����y-��^�/�ջz�� �G����M��]�;X��^�ۆ��KT�xc�X F"Ҷ��Ww����C�{��5$���cRM��ԟ�1T�<V&[�F"��
�@t_�T?����gRN��Lt~���@%j��:�c�=_v\��g�x7n�r��]���1p���c(�ܭKl����y���8�=ő�<PK��Gm��9w�����x͒�n�=��\A�O<jKm�0|�&�G-��{ן��O�y6=���p��� 潋=�RG��B��Ұ�v+n� �� �ݏUR]�y`�z��n7Nݤ�]�[)�f�k���;��엁��3���{���23K�����o ���O�����?Ĝ���jI��;�I E��B :	���i?�v��p"Ĵ����\�-����F0�"<s2�f��v����ά�܋	����
�+X��+f�#��H�6��kf��|uS2��4�pb�|4*\�jAài3kV���Z�ˑ&����r��92f��*I�Nu�s�X�U�X�8��{L[-�u�04#^�5�5�\iz�����=ҧnQ�Tli��2�ܪʬT��rI�������=���1yyȃ�D�Yi1�k�͡td5�-�S���aQnH/߻�5�v��S��'k@?~���9�p�:���_}�~��7�ߖ ~�~M�4~B���v+��9�p���}�F�O<��, ��y��;R_ʅ���J�ـj���9�b���D�z������jNZlh��[�x��%�, ��^�&V����� ��k�/䝍X�wk 7�^�����_o�߻]/���ױ`^�[�C�Ɉ2��j�/b]WH�ә+�\��9-&��.�\�E��r�<��a.��J�� ���lx�ؽU�'=-���ϖ���}��@E�u�����wȻ����| �w8߮���{�ԓ}�tk� �T�';1~��nfM4���~￯ =��^d򾯒��W�� v#e�J��m�؝�W����S}��;�{+ ���y���}�x���u	������U��e`Sc�7^ŀ�/ �Ʌߌ�8^؜�v��r���΄�$�cv�\�3�vxX̣cؕ�rr�6��[�-I[���<�ױ`�K�UUq}=���~V�h�I+wo ޽�? �1�=�߳�'?{��I>��q� ���Zmy�����n�`�z�M�ji�B"�� "$@��K���W�Z��x��� �b����ؕ��}��K���`��x��X��y��<�M��ߞ����K\��%���:�#�=�UT۞\ ��� �ٓ�~����v�m�
��s��a��3T�ͬ�5��m�q�am��	���@�-�3
�v;����\���K�96e~�靖5o���D�]�݊�]�;X��yꪪ���{+ վ��7�b�߾�ɰ~���CS�+��.^��߹8Wdx{�, ��� �����`�դ�%n��W�^�� ��, �d��1T�CG��^����j@�PO¶$�RJ����b��K�9$��:�#�?}�W�V��Mӧah�/q!Sذ�;e՚w"�lX���<#��ˑѭ���瓜]�0>[�T��� I����e`]�����$s� ��y��m[H�ĭ���eg����5o��	���K���ߪ���{����[�����eZ��)���7�b��~����;�ߞ�￹8��_zL�
�6�9��ꪥ6� n�׀rl��:�#�Dl����[C��'k ;�/ ��|���nI��{�s�s�RMF S�?r~;��b�+�Z�\���w
	%��1��J7S[�؛�n��'v�ͦ[HFW7lQ�l0V�L�l"��A�
���-��r�F�n� ���̽I�^�n��v��P炔fǂ���ý��.l��vV��i�z^,��K�������R�]�;jVq[+/4͓8��$��|Kd�hbO&ݴވs;����7�=���017�?O�8�����v.�Ս�� �c��bzm�&P����O+�922ܐ�+��Nc�4&/�10L�/��}��XWdx��^��� 7}��;%����7ui I+��:�#�}�ԑ5�, ��� �ٕ�ԐO
i�[hj�$���5�, �d�?}�%�Oe`��xzm��a	ؕ��v�=UT��x}=��uvG��着�}�?L��~�_����N�!݉[��96e`��׾��\���K�?}���u����c�`]�0�o��ؿ�)/9 U��.ֱf��лl�QͷU�q��������X����Ww��Xtjx�tP�ұ�Nݼz�,����PQ��UmW�Z.V� ��" ��$�!E�! H ��ȄE�&B$��B! f0I��B44��gDHA��GGU��^Xgv�	��������_$�'��Wv+hv[������2����~�瀞�~��G�� &ĝ&
�.�4�؝��&V����,}_WԖ�xd����;�iJ����꯾������z�M�X�iTt��8�AP�F�3��tvGKT*lɁZ ��e�.k_Ͻ���~��^�L�cU��\���K�96e~���}��_}]a���yX�����+n�`{%��2�����س�Wߪ����?F/���]��!݉[��7��e`]���V���;�����a:\oJ�R�
����8`�5"1b�q.���J�ayr�&`�Ik�S@)����`�M!�|��tR7r�p��	��CL�U��ac�&(VHq8@�A�3dj�(J;�Ʀf���p�7����#�7D��'˝W�ɴִ&%T9���I ��$�!CHc1�u�M�K�MhV Aa96�3	F�""������XH�R1'�ً.kZR��b����$�+�p�W�?(aB(��:.����&EM�PMeh%�*��M��D�@G �G
F�	��
��Z�t�])�ؾ����m�u`��x�lun��ݰ�U������-{�<k�X��x&̬��S�(wiX�'n��{ﾥ��_ 鱗�����������R�lsnZ��n�[/`ٹJl,��hz4]�s�������I�N]��z~�x&̬�l���W�a��������_Ŭn�h������uM� ޽� ��z�;���c�	%wX��x��X~����7�~�����X"�n��n�+J�V��z�۞XV�� �ٕ��UT��}�^��<v+Q��'bV"���8�#�=]��+�j��o^ŀ~���y�|�Y ����l.���8%�m��#8��=b���ⴙ�R_�sk��㛥�\��=���XWv<z�/}\Aվ��$��4��]4텲�]��ݏ ޽� �� �ٕ��H�J���V7I���&��qvG���.�{+ ճ� 9�{ն�WS#������&���ۀ{�߲���x��X:D�:Q%ujҧV���fV���UK������qvG�~��E}VmT�K<鴨whh��hz����rnV�Y�GD�S�H�w;W7(����$ۮ��ձ����ſ����j��l�ݶ�l��p��ˠ,t��:Z���1�ܮD�TI5��";vJ����ޜ���In�'�H�K�P�t\6���KAQ�L�µ�d2�(�T,�0ix5ڛ��y0v��#5�m�iX�8[��DE������ss�:
v32�Kn�����
��mG=��O60�Ωql_�P�2#�0l����.�Ҩ�B�V|�������Xdx&̬ ��7JZ�B�m+v��س�U$uo���{+ ��Ǟ��H݊�ט_»��E���uo��M�XU}_U~���{��=�,kQ|�� T;�V���2���x��X��]{�<O[�N��]6햭U���:������m�.վ��>w��p{Ѝ��e�cb)����]u���GK���+v:�+Fw87�@?aJ�Qы��髷l����	�y`]���e~��� �s� 7Ȟ�I]ح���n���T��V��Ĕ�%  �@�P�":�{�~ѩ'���X�ذthJ$��ZT�ӷ�rI��w�b��UW�RR9�uo��~y�n��@�g��>���~{�$s� ��	��_}�.I8� ����ۤ�i[Vݬ��,��<�Lf޽� 9�8��l��)mHɴp�֘&�V"�j�Z�-[,�sJ��I��C�k��YjQ�~�}��pI1���=_}_}\A��<ח���h;�ݼ�Lf�������N��Ϲ�$���՚3l�.ݳ �_���,UU�W�Q_U�H� 8�D�*.�AS�}���W�ǀo��f��[PUt�۶һ�n��9ױ`RG�rl�`z���z���m��/�(
�����Ӳ<��}�Oq�G<�u�Xv��͖&eY��:6�0��������\���Ͳ��0mPP3+�� �mrD��I1�Wv<��/�}�諭�S��o�7I�`��iJݳ ��Ǟ�����<�����&3 !5҃�I�Ҷ��X�`]�����/{��`�y���GE���%b�ݘ�}������ ����f޽��Wʏ�H@@dA�u�w:�ԓ���TWc@���n�$���U���.����8�#�$��t47�eS7B��k������Am���6��7n0u�+r8����k�qڎm�5�s��{}�݀Nˆ�����=�{�um)��]%v��7v�	�p�}������l�?~x�߿c0��y꯫䂧��]���V�馮��}�lٌ�:�������5�ŗ��9�h����Y��3 ճ� �ۆ磌�}������ ��7I�`���@�N��:������znI�罍I;�wY��a�D��ꪑ��`�"�@N+��e��ffˇ6r[Q�2'�S���K�2p9�s�tD�rvx��1'V�yх"���(�.^�;���6�h�#��C^N����k��۳��M�.v��H�'Z����n�JZ�Q��v������X����w��6z�I�c�8.�c���5�p�3�A�h�:ٸ$��շF�TJ�̖�!��)4�*�ы��(��8�롶�\�.��bj��>�'��7�!�|�ɘ���nH��8���sh�Kfl�h.8�}/;O\�#мN�~w�����ٞA!3�`�����<n̳ ��ǀm)���J��An���<�����W�|��{�Y�E=����3�U�|��ח��b@��]�;v�l�Y�uwc�9ݸ`/�{���S���kZ�8D�ﱩ'��}5$���Ƥ�
?�Fo����8����K��kV]�p�ۆ w�^;�,�;�"�T[ױ��v9���<�ַ���]Vm��a�AX;Ya2,"%�����w<&�c��5vpw޼wfY�w�E�꯫��UUO�����}m�_�A�Lۗ�;�;��q �H��|(��3m�,�� �d��}_}IK��O�ի` �v`��X;�?}U�$n�׀{g�� �j�n��m[v�?}�W˻3� n�׀N��0=U�Rݿy`��΋�+����0�����U{g�g �~��9ݸ`A꣡� ˢ���tcX�0��WI�u����Xtl;S�s_��v>���V:�6�� ��e�Wdx;� �d������1��TDr�-���{��s�we���z�	ݙf{�;�׼R�MZ�i'bn���~0��������W�b�B �F�TR����x^�}��I;{�� +u;Bwi[�鶮���%��^��0���?}U�R���OKI�*^���ZN�wx�̳ ��Uk�y����x��-_ū�,�ۦ�듍��ܜ�1^��!v��a�l�nMk�S����,��CX�� ����j�y���0�e�ve��j�n��m+v�v\3�}_��l'�~����,�5vG�m)���
�䘂ݘٲ�	�2�?W߾�瀞�<g��|����ӂ�!,�2�oܓ���{��jI��{�o��Ra6�e��)S$�1��D�!� ��л޿������v֪��� �_UU~�ꯪ�{���O��x�ܵ�;}-������dvH���mB@ggbP�gv��WT�l�������*�N����9ݸ`f��'v�}�}���o���G��	ݥn��ڻ0�e���_}U�6~��ְ)���9ݸg�'�y-;���l>�nn��>����Wdx~����K�/� o�� ����*q�������杖{�<�/� w�^ﾪ��^ٞ���Ct�걱�%n���� ;�/ �ۗu$����RH���t�y�a$�t�#T�X� �a��"��&���89GD��hM��Jcxa��&E��<;�-8 i^}78ؓx1��i����O�p-IO�ARI���&s���c���/C��L��$Ѡ�F3/¦B�Ӹї!pjF,��p�����k��Ju��+(@�T�G�h>2ӦE�B4 @7o��lm� p��[Kk�Hl�`'l�$�m��$ �S�Q�E$ll1J�R [��:p���ض�@R9l)0�@{�1TRU�xp���-���Z�uRa"�� 2-�Nc�)�b�����ˁ���v7KC[[҆L]�l΅�L IH�'f�� D��ggN�hNpq���զ�^�c����O73�l��X.Ӛk����F�3��H�9��`m۵�x�����3�T&�����5�%�!9 �p�m.� WpD�!�&�mԺ�4XA�t���<�rY��x�K�ȦA�mCL�
a��v��2BA�-Ӗ��DA�8��*[�eUe3W�f�3�kۂ�h�vfd9t�cy��j�k�JV���x����#<dH�my�܅�,�j\�T�ny�⭲Y=1�͈R��`9ʚ;v��X����	� 23UR-*�R��FĽ��ykn�k�n�p�&"�+ҭAN���T�B[�hLm��q��z8��F}:(����h��jA(����#n݀���V�8�Uӝ�-�֐�BuN��]��ݗkU�E�6�������T��`�e�<W<t�v$�vy�8Z��woL)ч�]&����5��@ 6b.bF��K�'F�Ng��MUQ�����z �4��E��EkI�t�.��6C�&3˂��;R(CB�m�V3��caS.���@K���"�v��[K�"����6̈́��
�qn�jZ��N�d�R��9�noCSPA�V�<!.�sJ�ZS���rU�5*�:���   �n�q�t�E�&-����Yzڣ)+����S��5/G'@+��p=�s�t�"h#3;;�3��91;�ò�����-�p%�f��T�pLEgB�����^��9��E���f��'Z����%��]<�ct��t���!�rkv��yFW�u^�:���(Y8���)7���R�h֖t6�=nK��OVq���ǻ�ϓ�D��\�b^����H�x�S��
��	���(+]����v�͚B��LL����W!<�Ck�h�أ�X.�r��a�V��^�[*ڴ0�3n%��d؞���V��q,�k��bWh@��=�k��9b�Q�1Q8�X�i��� �v�� ���y2�t� �{��v�%����bp�k5����tv�8��N�fU�48�:��%��@P�U�X*�ˋs'']p�GK�k"qisZ�x^t��5V'��9ɱS�3[f��t@T<W
�cL�n��u<�Z�z��-1=V�W�I眏8��_-�'��z�	ݹk ����_W����g��{�}���R�c*�;/ ﾽo �]���`nǟ�������6O޵�X�cuF�r���%<��~���s���X�%��=�M&�X�%��w�Ɠq,K��;�f�7ı,O�f��0a°3]�y���/!g9!y?�wϯ��ı,K��}�&�X�%��w^��n%�`%��s�Ɠq,Kħ{g��L��i�����/!y�~��>&�X�%���^��n%�bX��=�i7ı,O��zi7ı,O��;��M	h��JL�Ktr_"����� XXKu��ˣ���E�х
1�'�[�:�9*�̹�s��%�bX���~��n%�bX��=�i7ı,O��zh?>���%�{�߳��Kı=�iŲc�$�&,��\�7I��%�bw����!�A&r(TA�LD�9�k�I��%�b^{�Γq,K��{�f�7�8���%���1���0�%����Ɠq,K��k��n%�bX��ﳤ�K�,Ow��n�q,K��9�cI��%�btǻ&=�e�9m̲g�Mı,K���t��bX�'��{7I��%�bw����K�lO��zi7ı,O���a��e�2\���s��Kı=��ٺMı,K�9�cI��%�b}���I��%�b^{�Γq,K���}q7Z9����+<�jݱ�b۵v\[v8�n�L8T�����1��YX�j"*�r{y�^B�q�{Mı,K�w^�Mı,K���t�B�1ı?w�����ay�^O�D�?�	�p��e�r{Rı,O��zi7�q,K����&�X�%������&�X�%��s�ƹ=�H^B����~�%2�t�Y��Kı/=�gI��%�b{�׳t��c�Hń��:04W�F�n'q�{Mı,K��4��b[�^N���O����Z9|������1�}�ٺMı,K����I��%�b}���I��%�b^w�Γw����/'w�`�}4qhK�<��Kı>�}��Kı��zi7ı,K����n%�bX��u��r{y�^B�k����KH<�]�vا�tvt����d�ѱ�kΗ�����s��1��Dv��'�����/'����7ı,K����n%�bX��u��)��%�b}���I��%�btǻn�J�Ե����^B�����:M�,K��{�f�7ı,O��z�7ı,O��zi7� b�#��w��n
Є`����'�����b~���7I��%�b}���I��?����������Kı/}���n!y�^O�w��+D\��'���bX�w>��n%�bX�s���n%�bX��ﳤ�K��/��B*p�0��*>2&2��(� ��+��c���PO؟��s7I��%�b~�_d�13�g9��2\g7I��%�b}�k�I��%�b^w�Γq,K��{�f�7ı,O��z�7ı,O������q���F�Fݦ��U��Cd�f�y�$͉'���ƍ�(]��>�2P�M1��O�X�%�{�~Γq,K��;�f�7ı,O��z�7ı,O��}|�����������f�[Qk���7ı,Os��n�p��LD�9���4��bX�';�~�Mı,K��t��bX�'y�8�1��1d���st��bX�'���4��bX�'��4��b�%�y��:Mı,K���Kı/'zc0c�eĳ779�s4��bX�'��4��bX�%�;��7ı,Os��n�q,K,O��zi7ı,O�dǰL�\�ɜfi7ı,K�w��n%�bX~U#�����'�,K��k��n%�bX�s���n%�bX�_����xY�>�}��tf��eU��j�.��n3�����@�MfѴ�\.��g�V��l�!�'��兮��� ��[q�r�� �3���A�[���*���m�Dj�ӥ�]�yc+A�8B���'j� ��z�lM7\x��ձ��K�p޷\c���l�9�K�2�c2��ayX���,$&�IsE��6 ��n#B�h2���23fXE�8��A8<�����a��LL��C�-����\�<��'W�Z�[�X8�ώ��M�I�1t�V�#�W/���!y�^O�w��7ı,O��zi7ı,O��zh?>���%�{�~Γq,K�w����tYX�j";>r{y�^B���צ�p�D�K���M&�X�%�{�~Γq,K��;�oI������c�O'�����fò�܁rs���,K���M&�X�%�y��:Mı�ű=��MA$C�{�4��H���$�Ÿ�0K�e5�W�/9�gI��%�b{��7��Kı9��f�q,K���צ�q,K���)Ϧmu��/���B����~ﱽ&�X�%�*����&�X�%��;�M&�X�%�~｝&�X�%<���9o�xE��+_�:��lۓ�$H���[�׍k��=�r���;d�;+�&�X�%����4��bX�'��4��bX�%�;��7ı,Os�����bX�%���.�aq,���3��Mı,K�w^�MÈ��́t��6&�X�9ﳤ�Kı9��ٺMı,K�{�4���b!���b~1��c�	�˜��Y3��&�X�%�{�~Γq,K��;�f�7ı,O��l�n%�bX�s���n%�bX��<{�s-)�8�q��9�n%�g�AH��������n%�bX����4��bX�'��4��bX�%�;��7ı,Nsڞ����j"*�r{y�^B�~��{<���,K��צ�q,KĽ�}�&�X�%���^��n%�bX��d'��i뗗.��5�]p`l���]�Ekc�ⶹ����} ��Ո��+�]@V	�i�Kı9���4��bX�'1�{Mı,K��wı,Nw��y���/!y�w�}�hetXe��n%�bX������?�T�&"X���~��n%�bX�����&�X�%��=�M&�~����'���)�
�2ە��䧒�Jy?}�����Kı9��f�q,x	� �)b� � 2
��ȧ��(�S���O��4��bX�%����&�X�%���MĦ=�.I�%�.s���K��9��f�q,K���צ�q,KĽ罝&�X��	�������n%�bX����\1�̸�f���4��bX�'���4��bX�{�{:Mı,K���Kı9��f�q,K���=�Lٌ��˹]���;Dm�q�&�ur��5�c7$y�!��s�aE�jZ�����/Ľ罝&�X�%���^��n%�bX��}�K��%�b}�k�I��r�����ۂ�!�9|���,K���Kı9��f�q,K���צ�q,KĽ罝&�~�k�ǒ�N���v��W+y��ı,N���Mı,K�{^�Mı,K���t��bX�'��{7I��/!y�߾�0�Tʀ��8n%�bX�s���n%�bX������Kı=��ٺMı,��� RV+ 1)�L SH��D�������^B����o�i��.3��&�X�%�{�{:Mı,K����o�n��%�bw���4��bX�'9�zi7ı,O��Lc�r˜ܚ]��Lcm���2S�0N�2	u!��WV��7
V"⑨��-�_9=���"X��u��&�X�%��{�4��bX�'9�zi7ı,K����n%�^B�}7zCRo��.�L*y���*X�%���7ı,Ns���n%�bX������Kı;��ٺM��<��c�O%���Mt��%��J���Kı;���4��bX�%�=��7��1=�k�n�q,KĽ����n%�bX�1��2Ys��JL�3I��%�b^��Γq,K��{�f�7ı,K�w��n%�`~Y������Mı,K������ZS&q���s��Kı;��ٺMı,K�w��gI�Kı;���4��bX�%�=��7ı,O��E@�?DT�|[���ɇ� �L���n�3V\��u�v�Kn���b)��� �S�-ęl�:��Ӭ���lJ �W�V8цv�,�k��t�Y�K��YQf����^��Q-��R�v���ͪ��ʽEMٶ�ҧU���Ɲ�*�l��@�mG����Z7L��ÇzR®#��u�jmxMc{[a�c
�2�
�9�����a�PQ>����Ґ]:Ѫ�v�x�����B��R�U��3
�M�v�V��P�˪.����%�b_����7ı,Ns���n%�bX�����7ı,N���o���B��������	�nT�eΓq,K��=�M&��D�"b%�}�߳��Kı=�k�n�q,K�C��|�������>�o�i��Ɍg9�Mı,K���:Mı,K���Kı/�ﳤ�Kı9�k�I��%�b{��,��nl�1l��l��t��bX�'{�{7I��%�b_��gI��%�bs�צ�q,KĿw�Γq,K��;4�Sԙ�)m1��8�n%�bX�����n%�bX����Kı/�ﳤ�Kı;���Ɠq,K��;�g���ma52-6��#u���S��6����#V��^Ӻ>�}2�<����15��q,K��=�M&�X�%�~�}�&�X�%���^��n%�bX�w�٦{y�^B�w�~�}���%�[�ı,K���:Mà�!H���:
<Qv�GJ�_�f%���׳t��bX�'��l�n%�bX����O�*b%��w���sm)�8�qq��I��%�b{����&�X�%��{�MıK��=�M&�X�%�~�}�&�X�%��wS�3�&q�g39�s���Kı>�}�I��%�bs�צ�q,KĿw�Γq,K�LD���ٺMı,K��Ҙ�r�.6s<����������>�r{xX�%���9�~Γ�%�b{����&�X�%��{�Mı,K�9���x,n�+\�h�͈xܳ��s�����n�t�/����{��[bY���s���%�bX�����7ı,N���n�q,K������g�1ı;���4��bX�'���,�雛GRܥ2����/!y���ϓ�Ol�X�%��{�Mı,K���4��bX�%���t��bX�'�٧����IKi����7ı,O��l�n%�bX����K�2hD�,Ȯ��p.�7��>�\�� ��3��@� ����p
��[��0c;VD.�!�!��/���(:R(:�� "D�o)4eE2Nf�� �vL�m$�њG���@��s	𦒹T�B#�?F�ˀ˰�)����c,І���GB�G�K�嵎 D��S��M�CS ����x�p9j:b���M�ܐ&cqv*`B����lv9T��P�!�P$ �G�
�@>|�@ �Q1��$t�uW#��>z����D�x�ND�޾Γq,K��=�f�7�B����m1����Z�g���K��q����I��%�b^{߳��Kı;��ٺMı,K���4��bX�'^g�Ǳ�ie�KHL�3I��%�b^w�Γq,K�W���Kı>ｳI��%�bs�צ�q,K��3/i�[��K�^-����kgR�cs�W��X�V�m0ٗe��ᖄ��a�����B�����^��n%�bX�w�٤�Kı9�k�B���%�b{����K������_���g$�Eʞr{y
�%����4��bX�'9�zi7ı,Oc��4��bX�'}�o3I��y�^O��xo�6eʕSag��Ա,K���4��bX�'��{Mı,K������Kı=�{f�w����/!ߨ||�gQ�,2��ObX�*�'��{Mı,K������Kı=�{f�q,K��"D#� � b�aH�aШ|�i�
�j'�ν4��bX�'��b�zf�˜K&3���8�n%�bX�����&�X�%����4��bX�'��zi7ı,Oc��4��bX�'���LI�q�6��y��̀us)씙 +3�4�j&e�2�b'����j�kI�*�@!��9=��%�b{���&�X�%��{^�Mı,K�ｍ&�X�%��w���n0���/!��t�M7͇+p.g���%�b{�צ�p ,K��;�cI��%�bw���4��bX�'��l�n'��LD�<w>.?b��\䴄�s4��bX�'�{��i7ı,N���f�q,��}�Mı,K��4��bX�'9�OV�9��ɜd�.3�&�X�~���߾4��bX�'�~��I��%�b{�צ�q,K��;�cI��%�bs�����dɌ�4�fnd�ɤ�Kı=�{f�q,K��1����4�D�,K�=��4��bX�'}��Mı,K�>�
 ~80ŀU��ߦs3f3�3���mR�Z��0���=Wg5�T��Ώ��R1�.�NŃe�[qH�.�Ό�+��9V�6��]	��Y�sSΕ��-��vQ�#��N��h�pNAt�.��Fڬ�qA�y狵���A��m�U�K��ż��7Nt�&���X�m]@=�8h
8;ckV!�1��:�b�#�۳)�O/ ��n��;��bp�+L�&3���Dt�c`2I7�c4��fV��M3��K��5	�+���a�O�P����u����&�-�R�l,���ı,N��4��bX�'��{Mı,K�ﱳI��%�b{���&�!y�^C��}�e3��ΆV���Kı=����n%�bX��}��Mı,K���i7ı,Os���n'�D�	���b~�LS��͗8���qq�i7ı,O~��l�n%�bX�ｳI��?�a��������Kı?c߿cI��%�b{�t�<S9&in1�I��%�)b{���&�X�%��w^�Mı,K�ｍ&�X�%��w�٤�Kı/;{���Ofa�K��&�q,K��;�M&�X�%�	�w�Ɠq,K���l�n%�bX�ｳI��%�bs���3YQe.�9��4F�n�Y/-y�#�S���N�cI���d���Й�f�q,K��;�cI��%�bw��6i7ı,Ow�٠�(Ϣb%�b~��i7ı,N����\g6ҙs����q��Kı;��4����*H��!��B*9T����LD�7�{f�q,K��{�M&�X�%��w�ǜ��B���������U&j4vM&�X�%��{�4��bX�'��zi7��,Oc��4��bX�'~������^B������1���q3��Mı,�
$D����4��bX�'�~��Mı,K�ﱳI��%�b{���&�X�%�y�o���gWi�3�y���/!y���﷜�ı,K�G�~�Ɠ�%�b~����&�X�%��s�]&�X�%�|r��# �[L)1�e�����k��yHK�BSR�pڪ��=[.�;��ru��C���s�i7ı,Os��f�q,K����Mı,K�羺7ı,Oc��4��bX�'�;�)�&rL����n%�bX����I��%�b}���I��%�b{����Kı=�{y�M�Bı,K�opc1�Y��ĸ�ɤ�Kı>�{��Kı=�{��n%� ��XPW�j'��o3I��%�b{���&�X�������& 1-vg���B�X�X�ǽ�i7ı,Os��f�q,K����Mı,K���4��^B����O�2���&y���,K������Kİ��~���I�Kı9�~٤�Kı=�{��n%�bX��w�����c&s&Ie-B1��ɮr��
�s��<}�n�[�f{c��<�[�*٢��9���S�bX����4��bX�'��i7ı,Oc��4��bX�'��o3I��0�����;���b����<�����b}��f�p,K��=�cI��%�b{���4��bX�'��l�n{�=�Os���?�?o��s:^g���7ı,O����4��bX�'��o3I�� ��b{���&�X�%��{���Oo!y�^O�{q>����ss�i7ı,O{��f�q,K����M&�X�%����Mı,��_���(�F-~6>v����c���I��%�b{��8)OY3�`���3���Kı=��zMı,K�w�4��bX�'���Mı,K�﷙��Kı?�Ξ����fL��9���{i<t���p>[t���l�y�L�΢�<��3�%�q���,K���~٤�Kı=�w��n%�bX������D�K���߷��Kı<w?�?�!�7�fy���/!y����Ɠq,K����f�7ı,O{�ޓq,K�����&�Eb`�'y���Ҙ�,��SPI�}�f�I�>�;��D�O��l�n%�bX������Kı;�j���dɜ�4�����9�Mı,K�﷤�Kı>ｳI��%�b^��Γq,KB��}�f�7ı,O��c�1�&1�9�nf3�&�X�%��}�Mı,K���t��bX�'��{7I��%�bs�����bX�&�������O���O��.��E�GZ�����Y�櫧r6B)��r)BY�cpM֦�^ ��3Ȱm�h�t���]�e��,�;�W�v���2��kaMs��Q��aC#�wZ�^9h8-�=j�)���p�ې��9�]�q�f�^N�8�GN�̘Dc=FK�G����b��u���\���rF�`�g�\vM�:9��v��zޝ���x���t��01V����I���������F�M̝��񁡳<v�fx�%ښ�z��e��tO��'�x�L��3�E�rv�����?~�Ϝ��%�b{�׳t��bX�'=�zi7ı,O��l�n%�bX��}�OL�\.�_9=���/!y>��|�rn%�bX��u��Kı>ｳI��%�b^��ΓqA�,K�ӂ���9&i3��Mı,K��4��bX�'���i7��C1���gI��%�b~�}�8�n%�bX�o�ʹ�����9=���/��'��';��Ɠq,Kľ����n%�bX����&�X�%��w^�M�/!y�}/��g��k�<���,K���t��bX�'��{7I��%�bs�צ�q,K�����&�!y�^N�߽�&f�P1�ًP�����1]���+,�Б�[g�V�.��}�wy>���##�a��'�����/'��ϳt��bX�'=�zi7ı,O��l�n%�bX������Kı;�h����Rh�O9=���/!y?}�zi7�$�"t �@0i�`�1����f�q,Kľ罝&�X�%���^��n%�bX�w��>����EQ�7�Oo!y�^O����I��%�b^��Γq, C1����t��bX�'{_��q,K�~��w̤�M�7"�9=���/�9�+���~Γq,K��{?�]&�X�%��{�Ɠq,K��}�Mı��/'��'ֺV�[r�+�'���bX�;�zi7ı,?
D���cI�Kı?{��Mı,K���t��bX�'�������2fL�Pm2�X&X�4
�k�+��fvy5ҫ:�"q�v�9[��hB%�.�r��^B����~��i7ı,Ow�٤�Kı/y�gI��%�bx���Kķ���y�����w���B������4���bX������Kı<w�٤�Kı9�w��n%�o!y;7�K��6�3RZ��9=���,K�{��n%�bX�;�l�n%��D�D�E���E�"$&u@tF�DǺ�0�O�~�w�i7ı,N���i7y�^B�w}�����r���K��#?���I��%�bw��Mı,K���i7ı,K��|����/!y�߾�����Rh�%�2i7ı,Nc��4��bX�� ��~���%�bX����:Mı,K�}�Mı,K����3:3i��3(�F1�)vj�yf�I�y�.��q���șh��̈́Ռ6���r{xX�%����4��bX�%�=��7ı,Oｍ*��bX�'1��g�����/'��w�3�hȳ��bX�%�=��7���LD�?����n%�bX���~Ɠq,K��}�M���b�"X��g�-?L�3�c��s�&�X�%��ǿ~Ɠq,K��;�cI��(X�'��l�n%�bX��{��n%�bX�p���3�R���8�n%�bX��{�i7ı,Ow�٤�Kı/�����K��� � �� @��)0� X�P���0b$��)�B��P�	����O��Ɠq,K��9���A�����y���/!y��~���&�X�%�~���&�X�%������Kı;����n%�bX���gh�+�˹^�n^.�\c\uk� Y���FX[e+rn�h����fE��n�4��bX�%���t��bX�'�w�Ɠq,K��;�cJ��bX�';߽�r{y�^B�w}��2�����t��bX�'�;�cI��%�bwﱤ�Kı9��f�q,KĿ�}��'�rB����~���+�M�1��Mı,K��}�&�X�%����4��bX�%���t��bX�'�;�cI��%�b{��=
bd�q�9�nm�q��K��@�N�߾4��bX�%��߳��Kı>1�{Mı,�1���cI��%�bw��ߖ�M�5��9=���/!y���7ı,O�w�Ɠq,K��;�cI��%�bs���&�X�%���øLN!���J2�܃&g�1�1�c$����u�"�@eXE�c�'M�T��C�T:O�ekXM�o��X��68*��131& ����Y#|�̢��;0\��ɩ�N�@3>z�NQ�|� !�k{�C`#�Ml)��\��b��$!,��7������c��@�H�4cxw�U%u�q�wǨ�Z��؈�t�XE���������b, ��3�x"`"��l	 � H���Čc�m]@���#y� �L��X:>���Y�̈́CxrE3'�HD��"@�x��7�m��-H[\rA���P����F���	 X)T��U�"��kvk�-u�^Vɜ3Hr)sX0l�2a�Z��l��I�
X��e�n�퀲dG��59�l�����Ur����S�v�C�4��Sde�5� m6͕�Aڵ��`0�.z]�Z�lvm1�GI��U�2�u���rj]Ƨn.�fe�s�]�-�u����)џ#;��͘J���]آ�)cXN�Z	CrGg�: $G�/#U�%4��mIvD�4�ܦT�O� ύ$�<���1>�9� Îx]�q�;Y�Ӧη���rgdq�ΪB�uuY̪�K\*���]���tc9���ݢk��b��bl�4!km��d&��W�eBCAÓPū=��5x�J����\�.�{Wm$�-�8<j�� ��̫H����	���T
)�c`�֗P(O����P!GQc�ej�>�B�d+5%�; ��QBsڥl��y��ɬ�
�+jڷnu�5�5Ւi�d��/����ȶ�d�R�k\��Y!�Su�%=��K��GJ5���*1K����s���.nw��na�sΝ�µ�q�Z�9c���/��)l\�1kr����P�b�@1�S���uf&�r��F'VJ�,��*<�/2&�4���s��-������N75��yK���l6@A�
���Z"Y��4d.�-а�.u	ZV��5��nX�h��Y@=�8`�n�X	�͵��:�V�.q��g�����UZ�9�K�YGU*ͫ`[@m�l�,3kŠnF�̲��� ��j˻5F��n�2���X-D�sr��+�<��Җ��k+��3�n�O:mA�$z��v,�5!Z
��y7T��ۢ�6��Bg �뱶�73��'�[B�ri�F���0Vݜk�$��7j�J]E�u<[����u �^-�
�;\�ض@�eX��^m�L,�W����S���n0���{��u�!� �0 &] ��t!���
v�u 2�T��P"�TD�� �D~��'��U9�7˜\�ɌK�
X�6�F���r����
J�GA������}\�y� �0��1d��qg�a�t���E�G�8�zV�n�]�R�3j瘇�E�v+ۮ���:�;��q:m*��f`��B�)��P�9ݮt厳tv�!�\�ˣ@;Y�����h��e�77Dsع�t�����A��xqx����	vq4Sl�!P|Yf���3G�:p����Yr�\fb�I;V0 �i������{3�ՙűŀ�(M3*ш�#SB:�nɕ~�����/!xp�{�i7ı,N��4��bX�';�l�~H��1ı/?~��&�X�%��~�pa��3�R���8�n%�bX��{�i7ı,O��l�n%�bX��{��n%�bX�ｍ&�$/!y��}�m���b���]�'�,K��{�Mı,K��{:Mı,K�ﱤ�Kı;����{y�^B�vo�.�8�P�I\fy�q,K?@�Ls����n%�bX�1�߱��Kı;����n%�`';�{<�����������e��2l�I��%�b|c��4��bX��>Ͻ�O�X�%��{��&�X�%�~���&�X�%��P�]_`���9��:����qd��:�5�e0�6�Fn�ŻYsr���8r��el�`͗s��y,K�����I��%�bs���&�X�%�~����},K�=����䧒�Jy?~~�ĳe�j]���Kı9��f���|k���X������v<�F�Jzn�hVYwu���x)l� ջ�ٕ�Mq�P��U��nӻ��9Kdx����̬%�{׀l�:t�Ȼ�RK�Wo ջ���Or��{׀r���n߽j���h���������q�e�2s!�y4:q�����i�?��ϛi����n����w��ܜ ��Rݏ�qRy�����n����m�� ��Rݏ ջ�}�'?Ii���ݕ��.n^�/{�jI��w�5��)c5�r+q���$3*��DW �l�����' ?��^����X�[4X]6��~�����ry���X�%�{�<�~����ۀ~���ĳ
a��nw ����I/ �-��[���}x�F3m��Ef�����ܰ�ҩI�:�*�;�X�.S�e��_ϰ��v:�S�]p��� �-��[�������1��4e��ʾ[}����}�s����;'���K��I=h��A�Wt:I}i��"�� ��� 9$���G�uM��NU�m��N��ݾ�I&���RM���5'E��~(��U^���=޼R����MГ����� ��R��v<��uӤݣZ�Q����*��XM�Ca��2�mf:�]M�s]������;���G�jݏ ��� 9$���;b���h�f˸��{���i�_� ���9Kdy꯫�������R����U���߿_� >w�x~�O"]���E'�޴�ˡU۶��[� 9$���e`�c��U}_-�>��~�M�R�*� �=�����|�_� ��	�EeU.w��ƴҞ��s�KMv��b���Ӽ,p�q���s��u�I��\=�@ڧ]8�����Gs�N���+cf]�-�q+�2:�2K���=��`�!#l�nz
���ծ�z'�&xX��T��;����;u��=v��!��q�7�pα�S����r��m^xh8��GD�C۱AǨ9n��e������0�|vqh�*�Q���Jmfb��NI�/�6�G��ˆЍ�E��5L�nF@-�.���52PMH�.�-`��)�������ݸ`$��r�fV�7��9V��"�I;��sv��^��2�[��磌�Kޡ��MГ����� ���9[&V�E'��_�g����h2*\ܼ������}��;�p��]��x�ּ����n����+��5nǀsv��^�ݸd��<Oj�Ԭ�9��V1�G&Ɨ5�BƆ,d����)�<�v�D��Em�447i]���p�~0)#�9Z�.������[�Q�*�Q���{�C_+E[�z�����VU�U|�/�#�`v�N�r:"�H��w ��G� ���w�{��`^��ݧ
'��I6�� ջ&�0)#�'ap�:���*ն�Zi'v�	6�z���>��~0[��j"�$�.ݸS4.c��Ű�T՘���.��˙W�M�v����f�6�r��/{��'ap�5nǀI�fډ��iQuWt�ڻx�.䈤��=�~0������{b��gB,3�8����w��f�L�^Q���(PD�_�芝C�U0�'����x��/�#�
T��Cv��M;�����3���� ��� ��:Ғ˥Vڶ�e���:�ǀN��j� �nR-��E��R�YOi���ù�F�ɮ��-�)�r��8v����1�[��k`�sj��}�?N��<M�`Sc�;��C��]��&�v`�#ͯ}�g��`j���7����_$uvn��V�i�[��6~�V�6<d.������s��܃ٜ�I?I$�}���ߦMI'>�s�>$%J׵�J��NI�O������wb�,�H\0{%�d��:�ǀ~��?��}�K,�,��J���.n7VR�CG��?�$y�M]фL�i�K���wsD|t�Jݺ*�l�4���� �&V�6<H\0	�R���]�7wx�2����B��/=I���Q�*�We����w �z=8���	�e`�S)���'i]��$�� 7�^6L�W�-~�xv��=��M���엀M�+ ��� گ���}���I ~ۥBܼ�J-�\pe�9ɐ�6��F,�n{�Eە��	�n.qd@��:�]y�f;kblĖMՌ`�3���{r�v�p�DuF�ű�.�F�َm�=�q�Ɋ���n+�C�"�拳 �������
�r�q�`y<=�Êr��[��γ�`��Tm�&�=������9��Ś	��鲛������.I5���2f�
�P:�@+��wǪ�˟%����>xWʱHlA�G�E�6n(X���`��^+��r�w�9=�kذخ�W��W�`~��� �/����� �6g ���v+� N�x�Y�����;�L�)P�鯮��'���	�/%'�y<���ߏ-���#���,YQ�	�/ ����&�� �u\0�\)SwMخ���vL��}���sˀI�~0vK�'Z)��V�F�)n�� �fb�r�qt,�D���#��qi�s�Tfѫ��]�p�����\0vK�7d��;6�S_]�Z��v[�=���ϓ䄞vxy��`X���	����Q�� ?{�w?s:�s���I>��q�Ȋ�wi��Ѓ�+�	&�� ��^�&V�6<v+�޸��)b�Э&�n�ߟ���k ���<v+� od�R�D�i7BN�AcwXT��خ����2��S�{��w�P����;����U�F�α]�Mۛ�v -%������,�-]���_� 7�^�&V�6<�+QGM+��kT�����=�{��?����WG��hn�v����$��:�ǃ���Ϫ�sj���T 5�E�߀YzǟP�:0 L�@�u ���a��b�� �����6l!�C!�G�֝�_o���mvm#�H��%i�
ع���a��0.��8��F���Q\:�H0�S"	FV3k.�:
��L��d�FAB1f���BY(3gƂ	RTaP�	T��3�]4&>��h8` �N����0)�D��>E�U�b�tLtz�)B�A�.����Ԓs��u$��),�n�]�Юӻ��lxv+� od�d�Xf��k뻫MP$�+�xv+� od�d�XT���s�w}�@�ik�Rfc����cq�2ps������Z�v<E��N�8l�=��C�$���	'� �&V�$~�����߿�����q����Ҷ�\� ٳ+?W�^����~0we��ԡ�m7BN�E��)#�9�ذ��$������dE*.ꋦ��]��}_|��X$���p��gުر2�'DR�o��5$�s}n�:v��WtZ���/ ���L��:��<�=� ����-ձ�&��i�u��մ�p�4-h��V�7�_��l(Z�rPs56J�����޿N���x4{ n��ik%����m
�[� �<�U�}_$vy`�׀rm� �1���V�|Rv�ݼ�=� 7v^�����~0�{� ;����	"ݬ�O^�K�ql� �b�:�7JX��������p�?W�U�=��;<����j�*�H ��j��HTn3�(R�� Р�<�Ο'e<��s46A��X�����:y
<���ƍ�Ʉ�%��0�*7b�ț�i�%��7n�{p�����^������7[�~���7v�Ʋ-�Z�ɶj�5ׅ�$:��%n���u�f�s+�^�����.6c�Y�،�/&�.��6�@��ų��X�W	E�s�v2�a^Jy]���-pK(v��}s�A�b׃&�<�����v���#�f��.4��!�9&��}���������L�U�(k����z@X��qm]>���n���I�&��xfE���٠u{|�h�, ���nU5��C����]��=� ;�/ �ۆŲ<f�QX�ӷn����ݬ ���n��i�����t��56�[A���<�^�g��{� �b����9֖�]�]�Юջ0-����\���׀rm� ݖ�q�(m��T�LdT�����v�s�W<ŸՈ����YX���J�&qb:5��Uw ���������p�U�}���S�x���t ��՘%�g��O���P]#v��IT��H�h�,��ct����ZM���ɷ�dxz��<�d��({J[���'e�ڻ0=��W��ߞ��, �v^ɷ*�C"��骻Wo �b��e��p�8�#����We%Wuvb0V�SV-�n��Q�`;/C���m�E��xw�r��.l"�������M�`]��������s� ��~)S���EP�[}��Ϲ9�8��߷�vy`]�������ؒ�?]�]��&+� �=����X~�j�*���B����yv�t��ؼ���>}��8��gy�ѢBl����.y`[<�M�`]���J��:�t$�v�.�x磌���ul��9�ذ�Wջ3�UZb��S���֠�t��r���X:)�c��bF��B�z����ciT���5]�ｿv<�=� ��ǀl��)n�n�;-�� ��Ǟ��}_6o��� �=���p����T�g���eMS�wx`��ݏ �ۆ s�/ ���ښh����7���'�'�۞�����`;��+)���Ti}T�L��0��PL�y�&>��/}�%�SSh�m��������ݞ��9�qwc�DG/�\*[��s���Zn�s�؛���*�D�� T�*l�?��� O����p8���;�׀sG�`]��M�`���X�����s��|���������m� 9ݗ��P'��ӡ$[��qwc�96�ﾯ�����Tٳ߯ �ߖ޸��)V����ݧv�M�`;��h�,��˯g�=C�����	�hm]����}������׿_�����jI��=��p�"�0�D�L(}���eC�K�[��Ŷ z�ٞ�];� H��!jhe�m*�70S�5�5��]l��qu`9Rܔk1R<��LC. %�������6�ZU�h����9מ��!�6�ٖޝ��I�d�a�f��	�����s�z�뗋�e�+���e�9(��w9��(,��/�h��cp�؅����%Sr��p���0�.��2�$��rN�rr�������׋aYZX���Ebk������鱂e�ls�0�ɶ�Y�i��|��W�{��Xv<�n���� ;�׀OtO���,�vO-���������~0��x4{�k�*������v�M�`]��h�,�� s�-q]'V��hLwf�ݏ �b�8���{��L�n��N�ut�QN�wo �b�8����p�8����bvR��W�-S�j�E��`�mZ��RB��r���u���.:p��A'V�I�`]��M�`]��U�vy`�n�����7i�x&�3k~���UU]��#�;"�8���ﾤ�����@ݖ��ـul��9�ذ�_%ճ� ���5Wu�QWM|���~��]��,�g�ɷ}U�.��x����t�۷E]�hn��ݏ �ۆ�ݏ �b�=_UV��J���J�|Sv��cJ�MYpG,d�V�]��M��Y@�����SMb������|����|�ߺ{=-�w�m����͢.ء��V�3��X6K�;�p�}���x�:v�.�������?y`6Kԟ
H�\�i
b��)*�aB�\�s�k=��r�Ƥ	��:O���BH�k 9�^�ˆ��,�U���3��o���~b�N�b���;�p�?}_W�\����� 9$��cDi6U۫t"�&٬��,v	`�p�*6]�rT����|1�W`bm����v��7e��v`�b�9�ذ�K�96�ޢ�N�.��wk �b��U|�w��������~�yi߻���M3��i�x��޼�n�ذh�,�{.�Uuv:j���+���_}K��� ��,�1��I?���C��_.�xǲ������n�v�Bc�0ױ`��X�%��p�ꐲ�wVha����C���/]2=��q�m��t��V�r:5�[I�p�ƙ�����7�|�� rIx&�=_UU~�ꮰ���, ���?R���$�v��K�����y`��X#Ԇ�(���blWwx&�0ױa�������޼`����`ݖ��ـn�� �b�I/ �ۆ Wz�D$*vQt��X4{ rIx&�2I�c���|c�'��#�,a��F[~1%p��b�e|)S��(V��z���t��P�GT���L�@�FP��`pN.�r���$�F�F���"EBD��r*��"VK}��P�Ȱ�"���5]i% R����:!��2�!p�`W	�Le� �Iq��9�vU9E(줆9���^`@�c���D�\eL�"�H�2���1�L*4@jU�b�~�D3\�d�L��h�n6J�"F�#2��Fc�y"�p�����ɾݾ|�e*BA��0��n��%˽R�-&��
L�@V��ݶ��I�[	�nFʵ8���v�H���lR��)�)C��6�C�f��MA(T�m�c3
�I��b݆,!�C�-��Mِ�ve�
D(
����[��e��ȸ�Es��.�a�:�6�s���4%�g�RM<��������ӥ�M;NgK8]����n���I�N1<O��U]�I���V�I�uѽ
��7l��N���t.�0b�*�5�U�������5��W����ah�ۛ'`7f͂U�&6�eW&x��'Cj����-ƃ�LC��n��+�K�,	�[ @gR76�v\�&��d��:���
�M�p1��f"�gt<{d�ٵ�B��X��ƻL۵k��q�1]��	��z1�M��r\Ҭ�PrK]J�UHL�������2��4]����L�d�l̝��\+.��؞��Ē=Κ��
�Nwvn� ��u�^��	<m:����rb� ���5UJ��t�f�eWfH�����Ҽ�<��ۄm�CFH��s�p�HK����*�X�m�bV�#츷]�X�NyP3rkv��:��F��⇎�	�8̀�)����Z쒕���� b6�Ϣ$@p
���6���D�q��9{h��.���Vm'`<�\c�]3��m�E-��zx�ue5#@%�U0cǕI`�8��v���8�K%����7P�`Ո�h^ �tb��\����c�������ʹ�L��� Ul��*��� �-UR��U*��*Ԭ��k�ۦ�������֗BE�m�UO[ݲ�r@ul<K=����5[M�r�T�RhKﹾy~F��,��-dW�\7��Z$�3�p=;�$/�aEW!�V���9��M
�6�dk+��#\�0��<.:�C���m���V�*mt�-ۍ]nk�j]�h�!*2�]�c�c @؃)K4vq�k)�5��1�I9=�''����"�@b|�� cQT�!�P;�
�	g�����g���D��#!��dҹ��ͰŹ&�M�k����N�v���;ey׌Aչ�����Z��C�E�x���d2�����n5��5=i�_̼o�fyc����U�f�y��ѓ�ӵ;`�.T��;.,y��#m���mh���-8Ci7Nq�qnv6z��e�l�t��m=�yup�l`�f�6ę�ʛ5��]ŗn۪�z�epCZ:�X���g9,�s�s�*{���b� 8ICV]l�olg��B���[g�tn��/n/c���g|�癷E]�hn�@?~���M�`�b�>zo{x��^��i���V�W�|�0ױ`��X�%���_W�����bK��WM�n�HLwf�����X~����#�޼��� �d1���˥j�v�v�h�, ��x&�0?UR�'�H�=Iտ��n� sd���}_w�<pRy���X�g�;��,����r���w46v�X���fǳͬ�����u<��[M��/)��wx&�0���h�, ��x��'t6�݅�j��:�cª��a	�(5��:ؘG�8T��7g�1��$�{:�o��f��l��<y�N�.�����vy`6K�96�unǀlz��t�۷E;Cv�?}Iv{׀w��`[��~�����������c34�*Ъ����unǀsG�`6K�6K��L�MCۛ4v6�2�3F��٫�q�n�/%ĸJ�4��[�g�`뗵B�s[��c�9�ذ�%�����WXo�_� �߷��h�,m�g[��>zo{y��<��v{׀w��`[����H�$y�����H�k ;=��96����ĩ�Q�F
Vb�"�0�R��..��U4�9��c�7��X5�Ct���E�M����R�x�5I�sG�`6K�6i8;����.�Wfջ���� ;=��96�n�2�wm]�Ү_n� ��B���k��p��R�br�nn�$������Y���W|��߷ 9�^ɷ�v<f�Q��;v�ahn� sd��_Wԑ�K�j����M�o ���ܒ�fi�+B��96�unǇꤻ<��޼ �RQʺn��M�LWf����Z����vc���M�Τ���Q".j� H�����mֹ��I9�of1Պ��E;i;x4{��v{��;�~0���RJ������L�ɚ&���|�a��V�gӢjY8.OF�f6ͣM
�T��sx����;��v<�=� �M�Dv�h�I�]���p����|��O<�s� 9�^~��'�(O���ݍ�� �'��Ň��ꯩ#�޼��� +�QT@�S����j����X͒�M�`[��6ڎ��v��N��ݬ ��x&�0���h�,$�.����|�'oq���2LɌ�3,��m�nz�Dq�L���.�����>:�B��� [{`�=v^��tu�r��q״� �q��pvU�y΄�Fӵu�4������hFP�@P*�q�<J��ɶ9玄a
Dɷc��)�*A1l��lp`�u\oY��L���r� B�PזN�x�e�-�I�N�	+�ͺ�n"pK�ODGm;	uW'y�s��s����˼ܮ��b�(+�Nn}vx+�%�Q�y�5�t�������}��P��&%�fmhU~�����_}��ֶ< ��xΤ��t�v������v<���Ƨ� v{׀rm�=��RG�/MՎ��E;i;x`� sd��nV�x�H�t ��+(I�`6K�96�unǁ꯾������{��7�ɍ�_���X���ɷ�v<����/ ���|�6����M�, �b��v�@��<׎��b��eSh:,1��ڻ*-�)v`[�� sd��._���:P!�X���-��~�<�HNW�ڪ�ٗ�rm� �ݏ ٶF�;�j�v$��l��se����j�� ��`�:��N��Uwv�]��.V�x7U� 9�^ NƔ�WM�wiPخ��v<����/ �u�j�e�
�̫�8#ֲ�g�yB�M4Yq3�qj�u�p͢h�l&u���ק >l��rK�����{ߞ���t ��E�$��0�%���unǀsu\0k���)m1�blWwx$�f��^s����H�NJ?'8X�,`�J���g]�w5$7}/ �hN`�M��ڻ0���wmŀ�/�UU.�g� ��G�!%I�]Z����s�n, ��x6\0����浲7V���;I]c������D��z�M=���y�&����r�{O[pg:��۳x����;צջ�����o� �?:�ӫ�MU��wx$�g��#T�xd���/ 9�-q]'E�mPخ��v<����/ �wT1��UwE�)�I���|�"���^�/�R#��$�b��$-�(௝|���[�m}�f{#�"�ֆ�H�P�J��l��rK�ջ����|�}�ϱ%��6��$us$���\㣞��]����=�9�E
���N��>��vۡ�blWw}~��ջ��p�l��vA8;bnƆ�ـunǀsu\0�%��៪�
�Tx�T��կ��xdW� 9�^�.��� �'���$�8��ʵAi'f sd��\0���?}_}U����Ӏ{�}�K4њj��*��\0���wU� 9�^+���0�%�7�ϛD�U��:�֩n�.s�ajA��O�A*n�O���S��f8�&]�v }�v.���Q��6�Jm��7=%��أ�3�����K����a�n�Z��b�GG 챶�p��(�gEjk�a�bzݛN�3�i�v1vǢ�@Q��U�2mb�[Uj �LV3�0�m[�ؙAӞNV�4B;t{V��獮e8��76g�9�I��{��$�������-P�j�ጣ�Y�G6�6]��t,�l'���\Չ��Ɍ	jն������� sd��.�cX��TS����s��͒�l�`[���F�t�%'J��ـ�/ �ˆջ�����/��Yz�it�U^�{=�0Ry��K�޼dV��]�17Vݬ�v<�U� 9�^:�XV��ڦ�R���	�P�!ȼt�U��|�,�u�l�i��]�k��L�D�[e�)|�w�?��?���5n���׀w^�T�4�,���jI7��:ِ"�	 �!H+�|)�
�s��yu$���� ��{���-=��,��Y��+B��'������l�f sd�F��]65e�.�]�XV�x6G���/ ��X�cX��,������#��l��lr,�v<H�͇)�¤ˆ��j�^#k�Vh�]��  ��,K*��=F �D��y���ݲ�X͒��E�unǀsdyXw�F+�:,M��� ��XV�x6G���/ �I`�.Ƙ��aN��ջ͑�a6��U�V%_}Uڵ��eP�֢�a��|�`e�HlM#��ٳ�F�p$ �ҙ	�8A�!$D!N�N���i2#J�&"R34�'C)¬X���r?c�8IR�\�r@��l2h#M�jO�v���(k
�*�+D��#TIw����c;�عHm �rD��Q�ס(«	m�8��&�t�ϳ�hHJ�n��ˀ"3S��o�S8|a@�@9�}X���X�*��%���i��&�>��LB`�)Q��ҟ^Qܢ�
�$d1AX�P�lK�`n�EI@#j��vRa�01��р���D8�T~U
 ��A ����\����S5�a�Gq	�IEE	�? 2���@����,�&^�xӥ�B���ݼ}��K�����^�H�=��U-ry���0k���v�ـ�/ �$xV�x6L� �H�p�[u\��i9 ^d�v���'&��N۴Ňh��z�B]�����%�F�_lj�<�v<�&Yﾯ�����޼�i)���e�������:�c�9�e�͒�d���#�"�ub����m'o ���V sd��dxV�x��t�	c�L���� sd��w��n��^s�Ԟ^ Sjng(1�01dS(� H�@���J���)T�F$f�H0��A��1��'ow�y��N�b���&�� �ݏ ��#�l��z��ѯ&4�]+CL15���ZL�hĢ��x�� &Bwk��.��n�DP��d�7������dx͒�U��q��X��x���.��wo ��#�}_W�Ig�x��XV�y�H�~��1��`���v��g�xױ`[��vK���}�ꅚj��*��y�������"�x��F��]:l�՗V��xdxd���e��G�?�U}��	^N�:SJաۻ����֖���eݐ�.Ԩ���-���]���m6��Y��3/5�9k�@	�rV�;n���F�/��G�4��2�Ѹ�2˃ fbW3^㇣s����N����Oe�hȂ�����e�/<8ٮ��;{����پ���iU�^�b��[�-ȎG'O^�sȗư�m���������*������9'���5�e3sa3tlV3�z�%Ғ��r[q6V^Mn�#��Lnz�h�($3���o���������dxv< ���HK�eۻ� �v^ղ<���ݗy��H���T�ҿ�E��+��5Oy�]���U|�V�]����K�v4�ݍn��]��.��9ݙXV�����D!	�]������r�wfVŲ<��ٱ墊����
�2k3�1��u�߭�@�B*�r��(;B[��ˍk�������{��dxv<����Z�R�W,f�+f�8��{���	!<�d�	
J��2hC[�wZ�5$��x;�+ ��-�Ӧ�-Yui���qwc�8�\��ٕ�qI�!1Պ���%m'o ��r�wfV�$xv< ���HD]�E�wx;�+ �<��ź��_����񮮖,���r��t�,n5���q�^l��*�����.�[Cy8�7����wu�:��<��ź���̬�+Bp�bnƊ�v�.�x뗀s�2�)#�
�!�'av/��x���s�2��u��X"2[�f"�*o���uw���i*L�ڰ��-�wx;�+ ��ݏ �ղ��[eꅌ�l�g �{�w �<�����|�)��9ݙXͺT�;�Cnl����\H�n�B��蛣5qZ'Up�Ѝ�+����a�n�����w �ղ�wfV�6<`Bc��������V��9ݙX��.�x%GN��t�Ai]�����8�ǀqwc�8�l����T�4�����)��]��-[/$��F@��@! ���# B! t
9F�ލ@ٶ�NcLM��V�� s�/ �ղ�wfV�6<����M[e����2[xof�B��:6=��F��hېkn�Q�/mX%�iJ\��c+�>zo{x��X���W���'�~��X�L,,C�X;�+ � s�/ ��t��I8�Ӥ>[H�6�M�yC��� ;ݗ��K�s� ���XzҾ�f��cu]��<����߯ ����ɕ�qM� ����N豉X7w�sG�`�X���ٝI6�p�"�pU�.!���f�6���ϓDOe�e�x1�2r1֔Iaf�FͤM!4�kX���	�c�c���L6sq׬��aJ�a-��=q��1����V�rM�ע�S����z�5�	l]�K�vD�W�ݮ��bv��+�;�߿��w���<�{l������m��۝8�m@l��������^����GRY�nғH:5��w�1�n���g9��� �r��MK�Z}N9�8v�'K��%��o`�cgp�W<����q'lt\����::iK`�e� V���+ � w�/ �b�8�>j������)��{��h�,��+ �-��WlM6�h�wo ;ݗ�sG�a������XW�� W5Q�!;�Sj��h�,��+ � w�/ �����bL,,C�X;&V�6< �v^�Ŗߤ�''�d�y�~����kE�t"��[�,���3Ff[V7F(%?s��.��Zk��v���Wn�j��< �v^Ώb��ϔ?�����{����4Z�cs�jI>��β�i�B<�b�23F�\����6�MTΧ;1�]����8�#�6B�;��	����,��+ �� ;ݗ�j:t����颀.�`�Xdx���ŀqv|�"1���(C���8�#��e���,��+{�����ͱu�S�B\�wS�	���e��y-�O�.��a^zH �X��4U����K�9��X{&V�� W"�	$;���wx:=� �d��8�#��K�$���bL,,M]���+ �����|���5ₔZ�BI�g�ԓb�^�l��+ʮ�s8���� w�/ �Z��vL��il�t��e�.�;v���x:�ǀs�e`]���ꪭ�K��P&Ю��N��cm-&3cL4�uth/d�ؓ��Ve\�f��gn�t�X'w�;�O<��+ �� ;ݗ�`���R������9�2��RGV�� ;�׀s�lx:������tP����8�#�vK�9ֶ<�ٕ�l��l�hM6��wo�W�T�w޼����;ݙXHmb\20��BТ�,
Uh�}��:���D"HvMSJ��u�� �d��8�#�vK�'~�u�F#�R���RVR�Í�)��v�m�6%[��h��΃����Ÿ@n���ٕ�qvG�����5l��?:|�j�U�s<��w�Ϲ�$�w޼V�<�ٕ�H�i{�wE;,�eէn� w}��:����̬��<B�\uc�tX�����_-{<�	'��.���K�	�t�Q)]�Ej���2���������fI����I?
�*�� U�"�*�� Uh���@_�E U�* ���PES��*X
���D * **��H
�R���@"*`�D��B���A��@ *`*X
���H
�T� U`*X��H
�D *
���B� *��� ",�* �F"�
�`���"�����DH��T ����A"��H
� ��Q��E���X�,PH
�H
�Q�,H
�
�Qb�� ��D�",A"*P *A ��T"*P *�"���EF(�H
�U ��A��DX",��AH�,E��AH",P��A���@b��B��"��,��"��"�  ��PW�@_�E U|* ��PWb(���@_�* ��qPW��@_�� ��H�
�Ƞ
���PVI��]�ڃX�6` �����]��>��@  zt:ѣ�    ���(     6��TUU R	T*� (��A" PB��P�%R� �T�QTEB�D 
�(��� �    � �  � 0��|�w���^�>޽����sy�}�S=}�ž^�x��-�5��t�� n�ͻ4��׀ ��d��:p��Ӷd� ԛ��t�׮]ũ\��oc������G�z P(�� �QI�4 �)��j��νj�59�}�"���b�l��w/m\�u/}�!��@u=9o���Z� ���et�ˀӽ=+���S�K�O�X�x {�Y���}�����������u*���
( �EU� �W�n��S��n�헞�W����{����sof�����<��ۥ^� �;�n[��x�� W��w�Ϫ�x�O|���y�{�w��[ͻW��OJ�>����6�y^7�y׍�ż���� >|P(� UP&1��������@l��� `��� ��S@A�q� �z�@��A�   ���� 0T`P� �`  ��   ��4�  @�  2��
� $Pa 0:��P1o���[���zˏ���w��qgc����y�&YO\} S=K���k� }���K���� 힤�|���w��x�N=���}�{�_so-�y��70޷n�  ��7��J� h�Q��T�@  O���G�24dتT�(� ?BSd�* �"�)��AD 4x�ȟ�����9������Z�����{���H�
�C2�芀��"*��U��*���
�DES���!�%�0�����Ha$ ~M*4�@��rY�
h8��\��\����(Vz��e��`{=���|]FJ�u�8�B�fa2Fp��E���0a�P�$!M5ӽ�zn]���
~�$!� �1H�q�|p*F�F�<#"�y
j�ьf��6[7.����g��|�@ HAz�]�+M,H:HHH#H0� HVXRHR)r�	��*U��[�Y>�cƗ(��C����#R0%���i.F�Ϲ�����1���vn�3G%��0����C8������jA�����c�(K>p��!�U����ݱ�B.���s���f�����'4n�zW���P��t%�B�#}��O���nH~`C���~? �ώk�ঌ��0�ؔBP�P�P�!t`fǇ#��n	 �a'�4�HB&B�A@�*�.�2�Ұ
�)
�B�u����.�`B��t��������}��������w<s�}HAm�I��MɌ���v���*�J,�����~vhr�Z�4�r�}ffB\�����5� É�`l%��m�?�64�0#ď90�Yk����}���aMB H�D)��x�#��T���b�-����B���?3S_�WA�'IHG�ޝ~E���*�u�PbBƙ
��˯�	n����'댋>���a���a.���#�����^��q�����]`atdi�Gf���N�Hr"H�Ҭ`F��U+�HӃ"����Sz��`B�$4U0P�HB.�3�ٸ���dJJ2¨�[�+MɈϚ�HH�>t-�y_!���"3*��"����[��l�}�`:�Ĩ�S@�(.�HGJ@� :LR$H�H��� ����RB 4�V#X6-�H��	��$�H]<�9���'d>2- ҄b2C����
h�B"��As9�L���!R�]Jk	���\޾\�4�'��RB�.��7�hnt��8�z��O��?Wl4�0�,��-�.�4s�?�0���@��!O�5 �FB�&˽��L��A�$
�$�X�?F��}'4f�s/㌌5�j�k
�� +$ꁷs��ʄJ�$P�c��qH�N.ג2B�q6p�P��u�ܛ#�D��Č��0�r���CR�	]p� ˬ�B,P���k��<W��W��щ�#^?*>���6kM���;��.�M�)����Ǚ�v���R�)
�F�.:���yJ�>$�:���I��3N��d"IB��ĩ�*k[H�$���%њӾk�W\y�g�M������,~�a��M���h�h�B@ü9 ��4A�����YI+�N�I�}��F@���� F-�ѭgIrC5YM��n�!��R�_����W���Ԣ:vq5'�v���n�
�0����Ȑ����0 ��`ID�K$)��Y��4��5�P�eJh�)T�
j	�J�Mf� _jER_��@�5�BRH1!)KB@�FR�]��u�F�2ShB�+IHK3$�5�B��LJg��<d�ݏ��c������A-�%��e��.�P�:)�,Y�c�HA,���ebY`R� BH�1�2R	dԺ#����e��i������!l%!%aa/?]��4d���� &�B64#CZៈRf0�,�]�)`���)$B	!F!5� P(i��D�")�20�XV$,�d8\!�����H!���Y��kn�R�1!]m7����bD�F�*B��,$dȚ4��?����Ċ���6��dj@����d5H}�>n�v��A+.�u��!c!ֿA����)
�*A�i
�
�!��/sM��aԁFH��#H���aNIܑ�P�7!)�F�L+�ь���HN$)�����v�pHV0͜�S��
�0�9�A��ß�p��?p�T܆ߒ�a����53��[��$Î��\�����0�� !�/T�O�����6�$L4�,V�"�o�`HN���'�@� Ʊ����>�]��d���hE�����̟�	?K����8�a�$p�~�i�����3_�HA�G@��٧]l�M(|h��5b	H�]�c�����B�CF�1x=?D��SD��F� �!x���CI�
k-������%H�.�P�@�hHCH�aM~������B�a�C|���k�4��
k8J0��xJh��d��ͻ"YH��F�M�BB�"��JF^��l!��0��
�.��Za D$�I�nrRt%&�X��#XO������#	)�]l����q���@��	})U�w���#䉿����;;����5��Rǻ��N�Q���1"��4��N�iN�I�e�{6�:M�0�� ��T����dv1�i��)HāIIJjD�}r.}4b�Nsꫮp�N]�E҇J�����e���! I��Wd)��&��٭���k
�|�����R	O߈]d	.�]2��Μ��bB���2�����)�4H�4f�����SD�oz����~��	M�5 �8vI���=;�.���0�CdHq ��]�YMc����O�]��KF�ΧM���J.�(U�(i��7�vj苩B�"@�! �Y$�	&?~��s�^��w�n�F�����k|�^�ߞ]Ng�b�$��0�>��d2*T�4��)��@��X�?e�@�6�a��c�%�5����h�6�@�a�b�DBFd��t�Y�H�D.�7t$5�I���Lu��F�t�D�ds���,�Ąd
g�w�;�y~?sf)�U4F,ji���k�S�53��٬1���MCL͙to������X��E�B���޸B��Ѻh��Bo)���?�iu�ӯ^�ުƘQW���S����cv^~2��Xغs._�ꐏٿ�����HCa�Q�! A�Ha0`A�H\ַ4r�$��[ �HA��
��h�If�J�!�dJ�,�]$���bv�hHWP���X WfňA�ё�2��|�	F�pa�1"�@��|o�]f����Sg�7>	�I,�ִ�?k��S�a�֡&���"CP�����;�;�]Ḗt��L���̚,1���hBY��!XV�6!������Br���t��d�/!Bc7��?��)����6H�HR%�$R0b@�
1
E! @$(1����F0`h�B#B �`
T"�B&�dMm� ��A)���"S1i��bT���sf�?~�m�0�H�1�@�(�FE�	%.���b�t��R��j�0��T�U��UYG�VQ�-њ������f�8qg04���HQ�V���,�F<w�|��횔�ct�]��������a�1�$F.+�SD
��u5�c?}���$HVt�"�H�vŤ������Ju0٩Bp�O�&�+f�Vp�K�4n��p�!��!r��Z��,���.���dް7%t0��2�������tˣ���`�?MȰa�!RP�>!��tˡ�"ĕ͛��#��d�XI������>üӠ�����ɳ�N��މ�(��;���uR�O/S�o���{�X��W�������!������
�A��b���f�����쟾>����ˇ'B6C6���"]a�ax~�F�c�8�)�f.[������|~��A��bbp6�J0��f�]o\�O��[wB$$�n�%�p �Sq�)��� ����F)*��E�J�R�@�I�a5��i��~H�A�G��'̶f(f?�j|���Y?�&ͧN��
�`�!����ct��?��\��]�B�S�):�K��r���:�vZ�ݐ	9M�?3�0���LF+,R$4��I�3r�9��w��X��g�}�>��j�es�P�K_G}�e:�K��e8vr�c�0���J�+�K}����0���!D
�ZA �:	b@�WZ�5Hƶ�(D�3�|���wF�$5�k0�ٌlZ�)��0��q�]f�ʛ��B���NpT)
Z��q��I�Y�T���	s7�ɩ�\YdR4Yﴭy��+:�[B[��I%wi$� H  � 8   6�  �C� � �   �     H  6� <       $[@  @ ��  �`      <��KR��]U �JKʁ�@�����Y`m��ց�RR�J��Y{�5k�\[I	���d�:�����?���πpKL��4U�@�A��Mmm�m�����5 -��Mh�4�ِ8	;e��*�.����K5]+*Ͱh�zv�I 6�@UUuU*�
�*��R�@�m��Ѷ�l�j�е�35T�gk;)����޶���� �ԓBתt�.ݳ�,�� *�䪎6A��V���Z�..l��|����t����Ɠ�j��"�8�Z��*���2�����;mvF�윱�t��Il2�_\P-�̺�d���	
m�KvL�|�[��vn�V�J�UX�! �V�I���r�X׬�6��m�����Y�[C�r 	q��0(l��v���P��v�6�m[� -� -�6Z�����WP
�Ѵ����-U�uU*�m�	 m��$��m#��R�	�Z����36��ڐ 9�
���uK6�A��V����	ym�V 
;up�mO%��]+U��e��V�[4�2��#���� ��6� 2'jgs�)�eUX
���W ����F�E�iXl�R5N���Kڞx���5� ���헫r��
NINnF����[�|���3Z�� m��œlK������p�&nͫf�A  �kk^���������p� 6�5&F6�$$�p I[��iu%� ��[@  �	-�
^�kjCm�� ���p��it�4��@,0�m���h�` �  �Mm���mHm�F� I�@�l�M����V���bBh��6*����n�v�(���h�m@�`�A׎��ͤZ��xԪ��UUUR�SV�:-��,-�	��9�l۷n$�l[V*B�v9���Okv�����*2�ə�|LO��p�:jݩ��v�\�7P�y�.��q��u��Q����6
�.,��mT]6��	��HrMֲޠֳ���I^��dy�UKd �sV�U)Ҹ-���]鬓�����Sv� �����d!�B΀-�� Ԩ��ƥ�.ݫn]bl��n���ŷJ��_orq�,`ë��gE*�����e�[gm�l�U�1�1s�2�mT�H
Ɛ;T���KP�S��(�r��5�+������*Ԅ�R�fU�$�\� 8 h6�8    �ޤ�m�z�lH   �� 5�6�v��	��� UT���D˲jj���cm6�jG  m�{[R���[#t��rJ�� -��*ER�8�6����h4iT��K[pT��]�]���lm�G��i]�d����F*��*]�i���үREn��(-�mp�I�F�k h e��m�jٲ�WA­. �)we�����^j��e��N�T
T�`ŴqM�m��8;m�$��) kk5  �\       I' 6�P�U�  v�U��s[�ۖ�� �\�	,; )v�[�� �1��   I,��㭠r޲"�%�P ݶ&��� u�moZ^YUv%m �P�FJ m�m]+`�`���[l�߾��qs�k��޹k��c�z������L	9�1��(�nR����O���$sm&�u�p�QmH-�}���z��Ҥ�qc�ݰ�6��Б��gd6��f�� ��6� M���m���n��@mmJ저U*ԫ�[l��l�t�m�p�"[�N�  m���kd��η3Z�[V�m'��zf9t�i0lh����S�c�	���9��l݅�H j�!�t�m��l�Bi��}wq�n�(6Q�	Iú�m��[�S�*��t��'A��0��i-s1�cS���!�l�� ��F�E���ݔ=4A��NI`ŵu)E�@+�s��J���Ugps�K%��kE��:FTn����v��M��ic��� �i��u$[T��9�vŴo��W� m�rۚY#]:j������)�Yl�8�ݰ ��9ma�%���3��@m�F�Ib���[�e�m��d��fĉӋj�]����-� 
5î�$����i�r팅�@3�n���  6�t�i�Λ��e�wmb�m�	��2M,6�k�8���	��-� j�l��&UXJѻ��Զ�j�ٴ�۝e-���a��ڨ
��VѴ�R���y*\�\ � fj� ��e.roU n]��䖩x��i���5I9�;m���P6�i �Q���KD;�Wm��p��  [���m�mH�}��6퍫m����f��f   �`�ao"5��q�)�5�֚��W�A�Z@� ���U�-����Wf��
�X�Y��&�%�%�Y��c��&�X��$6ضCieri�%�6�[F��[Y-�  hHm}�� �U� �ZU۩f�g��0�X�,ڬb*Ut�lW�
�g[�!���5�Էյ ������K@mpm�m��M��mېm$َ9Ŵ Hm��݇ ��l����X��v�eݠ*�*� ۶��H�a�HyJ��Oi�魎������v�U㋤�'4��bZ��E��B�s�4�S�A�@�!��s\�r��v�i�����0ul�vݜ�Vu��&@8�JK��)d&�� �R��U:�[S��U��2��T:	нKn���hd/}�J�jz�j���BZ�ө��em��x��-�@��  >>���82R�f�kL�M�h ��t��� �@ ��   -��[B��Ą��`]�9��TqKUR�5���  A��v@�[p   4����8�m� �7m��%ؖ�M
�,
v\UPS��8,-�#u�!5T�*��N,5�l��-6�J6�� @m� � $WVg[@   4���׭  �m����m���@m��r��P�fܡ�UTq֒��m���f�vs-�*�*ܰU/e�`�ީ�� mZD��H� # k�F�$r���pm�$l6�U*�@V�@�uR� 8��t��d���#\�e�I��   F���B�Y%tr��T��U햱�����$]6�im �[@�#m����n   � ��      �� �      H���{�6� �i6ݝUT������z�U������	VVTr�*��6�&�k��m[ ��lh�A��-�@�����kn$�쭚lM� nӱ���\�I��GgL��Ҷ�nls�m�-�r�cj�!$�sIkHmʪ��R�ԫSq�7FP����|��=mSnR�*�mV��U���l�u[]7:N�f���@g�Q��[��<���WN���j�g4�ctԫPgn̶n��e[j�^݃k6��ki�  [x��`    oR�  $[G�m�[@��H ��?}���d�h� [@ �   ���-�m $�l6� ��8طZ�d[I�i1Ŵmm���      h  		e @  H6� Zl      ���lH�m���m��JN������H��q�ܐ[Kj�X  *�tRt�UmYp»�������Jfݓ��rWr���'��c0*�8m����ݴh1<D��P���a�-�y�[p6��Am m����i   ��K5�    -�D��ܙ5�� ��	n����bmq��h2��}�K�HI"@8mɮ�-�  ���%����=S��ݖ�f�m���h�D�C��ܼ�l�Sz�� ��I�mٴ�� [@�*�Ot�g����
N.���nE�m��Mm���KΥ	$:M�i �mn�� ���Vy{s�5F�]���׵�#sӠ9mm��	�8�������}��ڶ�ۆ�S]� u�`bր�媪Ç+3�R�UU����)r{#@V�� �S/]Ve�  �mփm&����u�    �i�ɵ�u,� ݩ���6�L�p  ���ɰ   �n�Q�;aU��]�z���`8��b�zf��YE۴��^7���Wm887Mt�X��Ht�@��}l�n���+���U�#�J�&g/3+T��T]km��v�    A��	� 	��   � �V�%�G���[B@�H$h �`�ːۤ�am����}�s�f�`d6׭��v�  � �WJK+���Ud���� ��i��E�˻���{���+���R�@�(@� ���G�����!�������D�ӕ� A�"�C}h;v�**�T2�Ө!����1��v��#�W����8� Q���	��)�U�C�Q$`��V!�9�(`�� 7��A@G��xtS�
8���N�� :	� �| iQ�7��V�?	Dz
�?"u*~A��T�ӟP
T�(�Ȓ w��|�`��=��x$I) 	���|=��t
"=���D@�w�k ~C��t�:�� A�uD4�8
QD������j�:~]���C��"	�pz��A"�Q�b�0)8 ���'�������)�
� ��R�"��l DM���ژ?@�! ��"��@�����l`�@ �U�@��bD��AO�
�P`��v��D$A�J������T� ,��`?	�� ����P�b��A��+*�(�p�H�D�=tA�)�2�I� � *� �* ��*,������*��?�W��"!ŵ �iR��� ����b"B i 4bw{�{�����m���hq �@d8�h�lm���UUV˱���@�d$�l�����Z�]n}�R�l�s���*H�*U��6*�Z�5��G��k��q����\	�J�J���8#XƻB	�4�U�p��*vi�e�ZȒ��m+�Hў�l�v�˚7<ݵS��oRѮp��8�H���7`�Wb�Wc���M�rԤ�����3f�c(3���m��t�WNS�.96��6[�Qz{z���7aݺ�᱗c���P�asc:c*�Y�*���,Z,U�,��� .R��ܽY�	��v�	��t�-T+Gdi����DA��'i��շ n�v�<�^���S��$0,B,��;k�L��tj��RF�!�U���l���ө�ͨ7g2(, v��vN��<��.�u�N�VQ��^ږ���YU#��V��%8vxX!ִ�ebkn�qyt�q9P;�ѷC�.�#X�vG�mZ�t
�ء�a������R���ZbZ ܭgR�o#���/��6\�v�T�N�\�;s�(�q�؞U��vLz*��0��� ����;ӱ�	Jm��/r�,�L�(��\A(<�S���)e�n�0vx�{E����.+�5�tf��6�v�w7�����n���jz�kFA{D�t�⚡[lqM�-��j7�c�2�S�[eV��Z�iH��i�"�<fp�5v�
�ȧ�������x톨
�ii�U�@�ehl[@��kCmg��E8D�,[u��sm��s��X8AB���u�۴�����y���۵�`&Y6ݣh��%q�*�*H�*�#�i��e%�W-UF�ݵK���B�b�VNT-��=7�Vn�Uvۨ v]8�N�X1��A����m��A.vV��]�7�=J�\��T��\�-V���2V[)��ȣ����*� W]99ʺV����W(��Q5���Y���2I�a��h̺_� �Sʟ�ᯐ@�~6� � ������z�w�|�����D" �G�ܹ�!�CV�̙�̪����*{]buGvCgX.y��[�GB챺�m':7���=7Qt3�˵��Eu�R#��)���D.�O2AnX��P۩��Jw��D��-��F%ܫ�1� ��Q&��F�z�݇�X�c���;\Z�\,����n��tl�{f�8�-�^(�ܰv��.�3�:y6{5�|���.)tt�w{�������ޞ�ȯ��;��1�+������vv���x��2��:n�I�<���٥��rT�����D~�>�׀s����eZ-Z�Mح*`oH遰��oH�dt�;a>�Yk�Ai,ISa�� ޑ0&���GLL��e��ċ���*`H�dt��GL�GLmE���TeZ*��$��#�m��>f�X �w�r�
9>�E)(��X��ٍo&-�<@r��3���ZZ��fh�jQ!Ϗ7%�������~~OΘ���l����K��e5���Y�7$���voc�C�Bt�M4JFѬP) %lKR�aUq�J4MQ
5(����!t��F��f� T�:J�LU�~�&��Ɂ�#�d�̻��X�]լ 7x��XtD�7ذ�=�`f:�bR�'Q))%��ͺ�'tt���0	�&�.^*Yj�R����L	�06u�Ll��?}ݛ�xS��ޞ���kY�̹M[\�`�g���[�{lwf�i������ѣ3�`��%@����D���^����7��V�mՁ���I��S�H)(���M�0'tt����oA��U�Z3t��z�(����I`{w�V�X=���	
�N�1`����~�Yk��V31SwGL	�Ll��;��R��u�/�V,T���t�&Șz:`N��������R��-����=#�^9�S���\�]e��r������,h��:��/%X���������wGL	�GL�[�$��:��II,�mՁ���w� �"`I�.Z�.��*�&칻X�x��<Xy)������ՀgV�i$�6N*j'$�s���w�?����$�!�B�	�5(�Њ� �y/}���������"I�*�7���kŀ=׋ {�ŀt$�\�u�m	K�=z�x�������ɳˇ�n�lva��M��U�,�t�z����_ͷk�X�x��<\�G������|���SV�,��X�x���� &Șz:`�	u(,WX���b�L	�Q� �"`M��;����IH��
��*�ԗ�ޖ�}u`nf�Xܭ��3n���c�*�3wx�^,�B�o�/�v�ذ��srG��n����$ !P�#��ɚ���.e���خ���uJ�ݡ�^���1e�n�	��ok��q�ES?pt��N��e"8G#6�+�9�#�����K���vj%����9����d+���9�p�ؑ-��c-I�w����ڋ�l��q�r�t�-�<�m��v�6�[s�6n���{SUR�[��Żn3�y� �Ԁ�@�%�޷E9����7�v����ܝ��݋�@ڦn䌜�i-;v�I�����Wn��,��=��b�.����,�h�苆��R�
B)+�=�z����mՀ}������X�j6�N�jR�rJ�ڞ,�Q!�w^�����^l����H��`n�7����0'q0;L�&�HVD����t(J~��� m�,�<X��� ����S��9L#mʰ33n��G� ?6� ��x����h�R!O��vۉ����v0��\�q֓�[ 6���(�aeUM�Y���Z9������?7�, �ۼ����~�m�, o��I)%"7S��`n쾇�U{�L���B��A���0!GB��y?j~�7�rN��nI��mՁ��I8�*�$�P���ݺ`wtt��ꎘ���&T�j�2�V�Ws7k�$�[}�`Z�X����ͺ���m$�6�⦢rE�n��`�S�w_�>�ذ�x�7��K����Sq{n{x��ѥyz;�x�[tf����l5����3P̛�'�̤��"`ztt�������Rbn��14��ۛu~�D���Xl�0�n��}:���NS#mʰ33n��&�Np�W9M�&�0:�|}
�1�U�0;z�����������	���Y���IRC ��0=::`wv�Xܩ����mJ�DdcnJ�v��Q��*�6啎:����X��&Ymٹ9��t����J�
I`}��VfmՁ�Ȗ�=$L	2��TY�*Ut^%sv��x��BJ&G�Μ ��� ��۫�r��H=���$�4�㦢rJ�3�?[ ��0=�:`wtt���Ex�e��ņ^b�I�#�w<X��J!"��s�6�ڤ]T�X^]���0?I?z�tG�`n�3���%(�EI�*:
��<'\��u�}b�m��nkv��<�il�����Iy��`�f*`wtt���K`�&�GL��@B�̤�b�L�D�������,w^, �Y,E+�U��I![ ��0=::`wtt���5X��t����J�
I`}::`wtt���K`dL	2��TY�*Ut^%v�0'tt���K`{�ܓ���7$��@�J%H0B=���_�Z\v���CRN�7v���8x:9^)Y쎹�nY�\�-�3�x�uζ�+�n��n�i��t��ը]��V��AuN��5a-g>t;,�2�M���a�u#�<�/l��T��`N�'���k��7�)�v���[[<tZ�0�ۤw�Έ	Z�y7Z,`^�rqɥ�x{*Զ��{ds����d9��7ct�q���/�%Τ������w�|}Ϟ��QѕmK���� W#���k���vLe�+n�lt�v�ʚ��^$�@�?"[ �"`ztt�����y�8�E:���I�E`��`}�0'tt���K`I\�P���@���ӣ���ll����S-��fb�%����:`v�%�	�&�P`K���+��K�9VfCU��{=��������u`��R$���H��J�S�6�J�/.����8����u�3Ȑe����ʖ-ٱl��$+`�&�P`wtu�����+V��Br7JD�P����vn4�SZ@��B�| ���L�D��"`I�&Z��2�*�-%i!������-�zH�n�,z�mt�D㤢rJ�32�����[����tW��aYI+����B��"`zd����� ���
[Ȳg�W]ڵw2%6˹�[K��r���o[��6���s9�a{no8�8㱷R:#t@�14���?yX��VfCU�}��������|BLr��� �׋9BS#nΜ ��� ���H՞��TLu'r��Kwl�����;5�?��(cG�t~8!C��Q�0%����]&s���q��'���ь�>�[���C�?OĹu�ΐ�@�	�K@Sk6ߴK�Ǻ�a��Ng��5s5�5����h���PBoZ��5��D6�����!T���J���XT����q ���	����������яR7XkY�a��td֑	��qR��E&ׂ;hl @�D�N�����it�O�\4� }�ӭ��-=E4�4��T�D��6!���@h��֣A ���_�>U���WHr�Dz��X
���w;��[j�ۅ��_f���U$"��ՓGi$�ٺ��$���KIz����Ǘ����u�.g$�AՆO�������$�ͺ��K3,���$��c��^����L��͈aON���N���)nz�<ɮ:s������ۆ�!�K�B��Eޤ���i$��kW�$��͋��ͤ���/�I%�[@�6��ID�-$�w-j��[�b��_l�_|�F��K�w*�����s�G�� ~�^��I}�u}�I�u-$�w-j��6�k�1�DS�ȭ%�o��y}�I�f������rۍSR���B�CJV��D7�o�˻m�?,�� ��9q}�I�u-$������s���1$��O�ZI/�av�_<���!VW����u��<�Ი]�ź?���O˯e'=\�y�X���hs���� ����~�ϒInM��Iw�z}�I�u-$���h�D�I��$��ح$�{��}�I�u-$�{�j��ݕ56�bQґ*��ZI.�w���76�ZI.�l���$��b��[��Z��iJ�$RW�$���R�Iw�f��I%�6+I%���_|�K�[@�6:ڧJ4�-$�{�j���s����I%��}_|�F��KI%۬�U�����k�> �M��lY$ǆ��ve\�.2S^Wh习����y�����v��=�f�:'�����:���:2G�_F�3=A��y��=��a�ۮ м��z���-,��;��n�U�\�X�^�k1��t���k:7tʈF��f��7Y� ����q�s2����-=�mM�P���ˇ�v���v�Eٷ�v�ws1�-��׊ӛ�2V�Q���<��sZ�ѣZ�i��Bk���[{l7C�c����QD�e�����㡥*1�H�1&���K2z+I%���_|�F��KI%�횾�$���B1�DS�ȭ$�{��}�I�u-$�{�j��Kwd��_s��F�@$�A�+�]ݒGI����d�뻲H�;��ݓ���$�s��!I��RB�Iw�f��I#wn����w~��I%��I$�4U��ȤIT���H�۩i$��߫�If���Iwf-|�]�j���I}��u�r:mr3��3��q��c[t+��G9��E�*�A�j�� �?����-����&���}{��Uߵm���KI%����R�C�Q ��J��Y�h{UT���ڋ�g�wvl������=^��ʦ�0kh��^�t�MII%�����$�ݺ��K�����$�f�-$�ݿ?%*sG8"��� o���� 7d�{�ww�4;��ܜL����TW`Ӣ)��%KI%�����$�6�i$�ً_�$��۩i$�u]�KbLdmpƷ��Q��Д;]#���(��fh��S*�����%H$!�>�$�f�-$��p���$wv�ZI.�/O�I$��4�"LU'N9I%��5��Iݺ��K����Ifm��I-
�D�7|�Gwn����r����S��,2�"�R��Z�*��] �b��U)5S�l�<�uJ|�n�i$����I-�SSm)IGJD�Q$�i$�ܽ>�$�n�-$��1k��3v�ZI.��=jP��T@'$���Y�p��^�g＿<Ē=��Դ�]�^�|�_��z�yz�����r
�:�l�q���o�����v�6��3sуc��᫠N��(�RC�$������$�ݺ��K�����ZIo�p��Y�ލ�#JH�I(��$�ݺ���W$�n��|�K߿\-$��1k��s�ʪm���Jl`J�18�i$�6�}�I-ݸn� *j������-����M�m����r���BH}�K��r��{�T��]�����m��w�v߂��"�:)�}��|�}�s�{9�m��c�3-Ԧb�ԕ-$��3[����{�|�K����H�۩i$�r��O�=M1zF	��S�'�u���f�S��s�<n˯��O8�~��w�������vl۪���� �����.�/O�I#7n��m%�M^|�^�Sɶ����"U(�B�Iw�z}����D{��i$������$�n�/ʹ�޺~b�r�I$��$���Դ�_lů����/~�p��[����$���P'M�C��i�*ZK��׫��Io�p��_d�_|�Fn�KI%����$c�I)"E�$��ۅ����������H���RҶ��}{�r�,b����"c�H���������]�n2�6�j�{M�eу��Dܓ�2`���Z��.��4�%�ݮNs�Dr��|.�<�O���oA�<n݊�Kն����v��n���ȹ����y,m�̰���6�G=��@t����gP�p��n����)rv��v��F��\%�@K��<s]'��dv�j�6��g���ӷ� n�m�cn��%�Ij�me�/�{����;���ևmg��[��;-{	-�p`,�<%rm��l�	V8Jv���}�˓u��rFjI.�����$f�Դ�_vb���ZK_�l��]�W���(��BB8��$�ݺ���Wꪒ%�<�?�I/?߭��K왫�\�6г�9��&*��IR�Iw&�?�I,{��K���o�7��H�z�ZI%���BIME�!z<�D__�򬙙���O��L��+�g�Q��'ٚy��%�u<�m�I�R%P$��m��gݼ��B��᜶��_v{[�#�Ձ���xĜ�$&�duf�nŴW`�j˸kO�`rWe�e�e�����w��r��R���	��_ g������~oDG��>��R�M)�\�殮fnI����[��G�$��!Q~FU�&�%R�dGHod4���Z�B�Q,@�SB�	,����$�G(�/�v,�]Ӏ��~��F���܍�TƉv��X�s��#�T?w� �]>� ׆��$J�1IV�ݛ�`���>�Ů�Է=���2��;��	Q�]�W8��u�z#�����ذ�Y��̪z4�i֨�TL(J0��Y���ƣ8��np�l�=�t�6��*/���v�q��MG��^-v{�u`g^j�+� Ş�ͦ���u	$E5v{�k<�G�*�uޜ��� ��9u��&O�����$�"F�����+���	�$�Ġ��G�Q�����`?{��Mm)E�H�r+UW9K{� �i�V�����IO��� zT��t�t�n8����`z��Y������+�������#���Ӌ�����u�e\��\&�0N�˙�]6���v���U5-�nFڂ��$Q��}u`}�uXٛ=\�c��`�x�li)J*b�IV��U����`w���#��ڟLu�`*�hX$����1���3�07�K`�wТD��N4�q���n����Vq�����J���O���`f�"�I'���2�kj�Rh�*���*R�`{dt���-���-���3�����q[�F���7Omj�\׃�����oe�t���N�Gu�ܜ�n0���Ҧ�Il��l����H���Mm)E5 �	��Vs&�{�s�0=�%�7L�A���K>ʵ������H���-���cǩ�j
25M(�?.��X��+�������̚��3ǈ�ƒ���(��`}�uX�9X�|���k[�s�{�rL*mP���4��P�D	�?�˓[�Mt8ji~]�_�\a���?@����2�?D EHo���ָ�h���5����4�D���2	4|t$M|=�lj
���%���J}���l�.Gz$e����c
ц�L�C�§Ä31DЩ�t/�����W�"@�0�	Bc��|�Ĝ�I�Ӂ'��'u�b�g4pt)υ���Ԕ��7�������@�
�j�
����ĀH.����{UUPr���+\ ���m�5v�����]&'��s��h��C�w&pT/5<Du4<����e�dv�efc�c�T�ʲ8�ͳpn5e0�,��A�|�l�N���	�.���U�8�l=dҘTv�b����-�	����X����NC`8�p��/M[����[j����0:6:� lV�/)���d�*S���LO%��3�/lV�Euj�q�����a98�W.j�;4�uQmm��4M�ʺ6tA�Lͼ�uu��i���6�+kX�U��V�<�A�\$j%6�m�b��ƶ�)�f6cT����.�A4��� �9E�Kt�%+*�xjXv�`W�)�)II(��X[W
�N�`6ő!��'[r�jٖ	��"�(k���YY71�ͷb(E݋�1�[���hM�t�I���� ���,���'N��H��kK�t\ʹ�������ucKm�\'�:�պ;4�A�ʸs�5ɸ�.�$���]���7m��E�e��p*��lp��#�2�u���m�2�m��ɎaZ��$kDGN��֛
5�Z���:Ǔ��R�����v�i����訮3�m]��h���q�??n�}�פ�3��"iz��p��n6��ʳ��8ۥy+�cpvNL�m�)Uz
��i
Y��r��:��68W�Y�b�U*��C�2�v�H\��&�kݫ`e�m�ۀ���'�Y��q5M�a���>�݌F��:��]�n���oR�=���izokR��rV�	$p`��Wj�i�2��;�aV���V��Tv�6��L�Rt�U�m��:�Dٜs)��Wr�0U;%�Z�6���G��`B����V�d�6��v�ڥb�@'�7.�UL�<���;���:PZ�m������� hMMO$L�`�e��u$�ś�;\�a��`vڲL�����ƌ��q2��s0S"ޢ�B �|�=AH��_º@?{��wq��z��ZԀq����M���A<��[Νθ[)�٧,t��0�o:��^�Y���K�5�xf!0�35���mGs���VM������vC9���ݵ���]Vv�%� .^^nyλ+�n�'k�Z�Z��u�O	퓑;��U�Gd�{�LT�J��L����[X7^��'vڠ�v���\�u~�Q����'n�y� ���)rf�O������՝�����;�����n,�sۣ����iYw��t�Μ#��u�)v�l�ա`���'�`n�L��GLǚ��̭8H�IƐ�V�y���07���7���
ݕ�YR�WLrD5#vٻu`wj��8�k�+�����z�o`��$j�JJ�;����������H�%\���h�r+��U��^kvۻu`wj�1v��F�#"Pk��n��1x����M[�tU�UM�@[U�O[�^Λh��)��^kvۻu`wj�W�7vx�7�&�m�r�)SD��nI���721`�1H�HX�	B�_Ȋ�]>����?}Z��+����D�M%)ELR9*��?~��s�DL���� ��b�>��N�:	J(FG��K6o���{����XP�<�>���ttxE��L�qSDq�u�`z������|���w������j�VVUy5�mv�%�Q2�GtR��g�K��<�6ݹ�9���}�=��nc�!���u`wj�:�5��s��W�WXf�~n��S��o�J�H���Wk �k\�%&�}X�O����,�~��l�~���R��$`8ۑX���ܓ���u�Δ2QP(�ϳ�ٰ;�|��#t:m���%#���q/%
!V��U`�{�ֹ���"�ow���&�D�DF��mX(Q�޹�:}8�]V���������Cz����㩓����حg����Mq�y�&�����p}��
�5�*b�I_�����y����5�r����u`g2�^j�"�Vr��rQ'�O���v,�s�
d4��x��M�8�%"�;�|݁���Y�
g]>��}8 ��Z��!QWw%M�V�z*�{�,�w� ݭs���  �FB5!�@M�8�A|=W����ߵ����z�o�&S�F�D����U��Ϳ�{���mՁ��V���ȵxmK�ON7eݮ�r��yg�OX��d�r������{���/�]��.�W�m��~���&�_���I�06E�Bt�~MTE���^kw���_�����^ >�^ ��frQ2|�u�UT��(�D�� �o��w3e���l�`w�� �qiN�	J.4�p��L�}x7|`��uX������T�*@�,�����l�<�!z5��O�y��`��x�!""AU��/)��t���9D(l��Dz���eG��\���:�{�-�
�n@�:�y�̷`ڶ���u��&��(su�`�g�ŵݴ(hZUr8f�ւ�˫��l<g;�5p�^�:�� Ijh���A�$���w�"n]sڭ{�����Jr�]�'d�,�H�6�[.�܆^�m�1���k���c�rkIŲ��VƵ�${���~w�����5I��m��6��p <���i��}�&���ݦCCۥüO����^�vc���S7s�{������ـ��Խ���Ӏ	��KʑB����M���l�(Q2k��9���?|�\�L��u$ߢL`H�B' �{���ɥ��̧�V��Ł����R����2MU]�tO7�`��N �v�Q3��������7��@$Q�X�<�`y$�
<����5�׀?�ـ~ҡ��@Qr�;۳� �A;��답����v���ӺnW�,�g7	����ww�o��7iSiWw?��w� ~����l�I~��O|�����t�JQq�#�����,��?.�G��75�g�'Z�Ӏ?�ٞJ!B�D%F�//T�*@��#�G`~�OŁ���V{��r��l�`ug����iC��Rq���ÒIN�Ӏv�� �?7X�IW�~�Xf�ԩ��tSq6R�XܚX��yA��Y���e�V\��=����\����;�!nڝ״1�+ͩ��OW�w����;jN�6�m������l�>�V�脿Hv�� o�7�U8ܨ��#m�`ori~��Ḩ�V�g����~�RGwct'M7��Xr]]`��N ��fB� �� �dB$S����Nsw�{[��`w�M�#�F�*U$V���ל`N�V ��u���m_�+ ��_��T��TĔ���w^��}_��T�pz�`Q�N,����:�a�nq��$�4�s��٫��*�@tZ'���'Y�E�Ӝ��Y��2� �V���8�x������^
�C��Rq�#���i��9ʙ>ŀ=�Ӏl�u���.��*�S��㉲����o���w]���%���`fS�+2����(S	��v�9D�[�X�}X��8�%�BuSb�xN{?{�rN��5�	5�2�+�����:c�gK`t�����?W9UU[X�_'%	�8
!��Aa��fֱ[��I�y�u�,<�=i��k����N��q*�8������`f��X.�U|�W�����6�4��F�$E`f��_��:��v�o���G���ă��^�M��TĔ����V���3���pϱ`�Z��?�ЊB�V�0:�L`{L�l�0>]�v��iC��Rq�)��G���:`z�L`od��π��Fݺ��]Qu ���mS�u�s��$�@�[=��[[3�s�@֌ⶶ��fMu���rd^�\(9mD�Z�euv4�J{l��b6����U������b�E9����cdr�����hp�r&��l�&;P������;v�hˡ���pu��v�،��ذ�q����x� ��\]ۊ^�Ψ��6���/��9콌^z�L���~�{������`{
-�xC�n�d,�f��/d���mm�2pN��=�]��l�fqG:~t������-��3��=�p�ZE�Tj9V˻���=�`{L�l�0;���V�-!ee`����=�`}��?%��]XY�v�#T'MSؕ@mH�=ŘM�1�b�?O�������=��7���QCJ9Ҥ�H�ܚX�^o��o��X��U��մX(��T)7����m��Ն���n-�xJ��\ݶ�	Z)یJQ)�t�S#����k�3^j�>��s���|`C�%��,,VZ���nI�u�n��(���T�^*�Q��X�Ba ��a	�c	FDP����H@$HF@�M&�Q��c t@��8f�БCbY*��] �A��7�5��'�w?˹��I����jND�"�7J}8��a�ꭗެ�]����J�6�U�N��VnM,�͖k�V�qf�Vpz4׈�J�V\՘��� �	$��O�7J�7&�٪�nS)')9��R8��6ƄӀ���+�������字��Bq �߽���}�)��(�t�'$���+���5�В�P�K������Q5C�(mH��{���ɥ�w�� �Z�=
=
*��^��P��n쩦$��=���`w6Y+y_.r�+�t�mN���9L�e�&ƍ���vi�T?1X�ؙ� ;j0�WHBQ%M�C��]�B.�� �Q#�1r���N
n�;�;3�G q ����"����5bC���?�c� �4�җt)р<�|�4�%�X�re�
���&��ҸB�(B�������IH�hj� ���6�o�6.��3o �d�m�;ɠ���iSN�Cp��Xgh��Tv�G�ثM���@Gg N���(����O���`Q���G���R�J9B��r�vp�N ީh�T˧(���,=ʤ���`o��X��[�(06��
�|R�|�!$��\�����>w� ~�]���S�CI��iUD��9@�B�tN5�gu�\��Ҹ��#/�?�Ͼ�۳%z]��6Wzp{l��k�G���p1m*z�P��N��VnM,���5��j�>���֑2�9V\՘��w�k�s�$�z�����=���`fl����R%�D����}-��d����;諾U���`oD��ġ@�jE`w��VnM,�͖k�V��+��4ƜQ5K�]���\����M�a��o����1�j��ڤ7�QR�؛dq|�g� ��3��7L��u\�х�b�.��,C ��3��7L���ٞ�>L���V���\�� ��N�����/��t�Հ	���;�Rr&)���R��+}�Ł�3]���U�}�)P�iE
���E`k�f�:����}8�Ss�BQ��ww��ww����7Wt��;m�z �FM��.Rx8[���v��˸m��];Ykpv��$���kNY�N���?}��　,���� ��vɦXy^�sa��t:um��
�n��pe�aw[qָî{3���WZ��Ѹs�n�p 	b�g��^R�}�V��pɽ<o6�ݶԅ�
M��ض��]�ɮҞo[������B�j��
�����&�ˆjkZ30�n����t���m��Ń1�n^1f'R@�v�ݜ�ڮ�Bj��CR���~��,כlC$�NP`wEY��Pf W����vk�W��{�`o�x�5w5߫�͍P����@�jE`w��,^�0�BJ!yEW��� �Wzp�e��DR����#���ɥ������y����RV���Zq	�D�uf ��u�t%	��O�>�N��K����el��D�N��Օŝ�e8�:;�5�Hp����ޜ�6=g����*G�P�,`tΖ��2K`t��Ur��[�v^��x�(!5'#i�a>�ٝ�٠\�/�+aT�*��IAE�����_��ٹ�=���uX۬T�i�
���ڹ�5�f����(�S/��p�s�`v�V!5[R��P���kܪ�*"��M��������5�!N���3vS^�(iԢJd�vn�,�Ū��٥��s]��]���6'N�!�^�kś!�ł��u-�l%�O8z�g=l���UUQj�N����������[�`/]tBI/����9���$c�bqE`f���Ź���٥��ص_�����{Խi$��Br����X�}X۶�-\A" @�6�+2B$X����
�!t(�������;_b���\4"�,�,X���lW-����TB�\��4�8]6I57quUV`�s�t(K���~�>���f -��W���\6�nu3��HN��k66	=0�k��y�ݬ��I�f؋t��f� ����6^��>ݶyB�B��?E�X^�A5_��@5*5���Jɭ�޹��?kx��mT�)��S#��̚X݋U��*�.�u`j���܍P�	�J��09B�{�=8ϻ���@���Mmm� �I%�ͪ�
�&�np��,�$�s���|`݋U��2�қQ!��qA�K�Bc���G���n�b� Xn�uq�y�&��ﻻ��r�HM&�I�bJI_ o����d��ߝ˟/�>�XC��\�Eڹ���>ݶg(��*���}8��� 5��^����9/H�/MMM�]UU���W���GL�D����0U�RQB�q46���r��.��X���n�0<���~�>��]dԯYD�*m]Mլ ׮�D$�Z�q�I���z�Iϻݛ�PG�"4"�E � ʁ@ , �@#W�ǻ�ݿ���u�Hn�igt�	1*���ڎ�Ml�D��Z�i��Ԇ��:;��[�ū<g�	^*�x4].ɺ�p��o�m��Yy8q�hg�qBf0�[TFz�����16\I�Y:Q8�3�L���a�;?�Wܛ��uLVp��9�.خuA��q��vx��K.��&�F�۶�]7�VU ��aZ�+]gd69�v�B���0�e%�.��k���_�x�����=��2��g�6C!���ƭc���e)m��v�ܠ����U9j��{��Ӕ�Ԧ�%S#i�<g�������GL�D���E���P+��� ��f��P������ 9�������\�*����"R���W�������"`l��Z���m�6��T�)%Xz�U�U%��y���0<�$��IB�~�� �w�*2(VEڹ���� ���0��&0T,Ř^d��������ӄ��ۧ5��v�����?<3�L�I�Bd���*�\�s��(��&�:o�~0�x�~n���D(��=�~0?y��F%*7�Ӆ��ݺ�r�J(q� ~w�w{�nI�����9�ͳ9(I)�SNɩ]b��U6���X �����0����|`_b�>̔�ԦөC�#i�,?W+�K��K��0�^,�IL�}xn�QJ���@rXf������ss}�|��K �se��G�[D�(�M�M7)�R��5�o<Z�7�ݎ�m�\5�y^zZ^�c;c�����D��R�����ԇ�no��7"`��
��;��B�/Ꙛ�X�]�(Jd>�׀=���7�x��Q2}��D�Z�"�\�]���7$��fvn @"$B0"�
�$�cTX�"a"��b�B �����]Հo���7��8�ą���������ŀ���u�� ��^�J(Tn&�8Xf�Ձ�%�������-���.�f�𞕑R^�a�+b�d�9��b�M��Vz/]2p���~�����l'}gܗN+��	�~L{�`v�A���{�e�F1ԡ���$��͗��U���q�{�~0�{ k�x{u(�ST��V�3Wx�sl�?kx��I(�>�����V��(FH�jBâ$����`�׀n���U90� -M#��@�1L@)�! υ�Lw�v�rN��ow��AV\�*���X�]�P�#Д$����:{��ݺ�3��$�$�V���t��U��=<DI{'i{,Iڢ�Vn�mF���U�9(�U5��͖��f�[�Т"~�>� ����nR���NK;���ʮUW;��� |����y�Q
�����jf��uE�QV`>�X�]��
$�L���7<OV�B�[�5*1]�%
e���o� ߙl��(J��w���ݔת1����$���GL�D���}*�D�҅����XE�3Sĺ����3Oߍ�e_�E��h.J�e!!b�O���\HG�I9N(U��l�n��� ����������z��b��*�17���c �$C����.� ���\�4�Ģ��Q;��Cd
����)D���ݍ>(ހ�!�����
��r�*]�����"JH5��m� $ q i�YY]���L��qУm�cRW�)�"q�p�4PZ�EuN�.(lvҫj<���8��i �\q��A�ؠ�V;n t�cU$u�ul���P�&���v�T��g2�+P=�v��K���[6�W\�v]�3=[L��uv7D���9nc` z�W#��f��N�iͶ���Ĳj�I%�パWn�(
M�2gWiP�V��=��y!n��]�I��XgsţZ��#!i�l�[`�1<+ֹ5v2����6��v���7che%�kHT�#j�LM+]���Hԝ���[��`wlo$l����q��v�w�� :q�6暬i�L]++Ae�0�L��
���]���݁g[6�[�nX��c<��zɮ�A��nA�:�z��
���V٘���EN�wA�=��DV�wb�8��=J�7M����@wR��#^v�U��U�����^��t�vqM��{e�cK�^;v��j��m�V퀭a:!;p���r͊C�25�%��w�[�5���alͷ-�l2�����2PuB����H��F�u+uӍ���a{�^ܳU�ہ�v���a��' vNSa��wK�����Q�q����l*�h6�����q�n�U���B�O�D,,e�.��@R�ETq��R��+�*ɐ��@pӝ�,��T�	&�U��l5[u+�����6��l� fض���@-3n�F�ɕ��[�JjA�;��U��n���n�����d)ꓓ�X�oj�\�;��7k�Ihr��&�c6�m[AL�X �U�YV�ڃ�-6.��uң���G�&����x��.�9���o n�^p�^М��@b���O�K��� ]��m�;F�%n�M�q�r9�/�[���k�YĚ�+LҼ���SI��;ېf��e6\u����A�Y)���w5+��T&��bj���Y���(��2k35l.H��m���u�� 	ѡ������T? =PS� 3��(����w��M�d;5�zki�LB^�Gj��'vU�7M�N�ܭ�IvP�w=b8۰�;k�g�j":��ܭΝl�`�^{ln�pvn!��۵S� K���n6�`�k�N��5q���g���F��8�������F$�m�9y��^Cy�'q��[M �eK�q���T �m�@9�{wc��Ԝє��nݶyt3���Pl���{�w}����uMT�'!u���� ��<�1z���	А�1��٦������>����7>�
��>�/���� �z��(^��K�}�����ߪ�J"��4��o��� }�� ߙl�P�L��E�j&SCrU����`��`{��0=�:`z}	[�P�>YYk��)�o� ����oB�R�ߋ �s�^r�%�rXf������(0{��0���d����d�k�w����/fܩΏHH��[Rp���fﴵ�U�n�\bQB�d`����b�5� >�w�Q�A�� �'e&��R��`gviUv��*�+�'�%�� o�� ����>�ҥ�e7R�Q��$,��,�I���U%�����Ow`�t�{ �(P/`n�A��#�lPa���䟕���TiHڐBi�B��wn��{����^�̶`�e�1XH��y|�[��4�*���؀��+������z���1�e$�#@�Jj�n8Xݚ`m��̶z"<��{�� �G�O��T �Y@�d��݂�H��3�4�s�o6��nR����������v�."���Y*@�� �Mu�;�gf����l��*��#b,=\��z�`�|`�s�?��`�lUR�� 6�V`�l�:#������,ݚX��6�2��7%6&�#�E�gN�\=w*�ǆ�;��#���0�\H��EK
�@],�����A�7�n���;z��9�%������M��� ilΉ��������l�EUr�=�}V�Q6��l��=�O��0�Q3������ m�.L��)�i��a���������߾3�ry@80 !b51�M(�O�R���E�h1X#��D8��w����'�Ǻf�B�WH.��v��f ۶`�l�=�"�$�������^�X7��nv�O]��-gz:�����(-D��2������M�T�rB�p��Ɤwf�	�A�$P`��ѐ-Z`���v`�fz<������=�_���C�6��T�5*Q,��,ݳ�����wu�|�Jt]
�t���E��A���K���`w�����H�(R�p��`�J;�8�o_nـR�x���w32�af��e̹�&�q :��)g� ��&��T�^�<�K���K#�С�n6�v��Z�.��؎���v��^(.
��HmG����3�q�l�r+`�Mƣd�S��e�{9_d���Ұj���j_4�����źv���/$9�y7<;��)]�۠L��팅r;m�UY�d��3=�).�\Wg�����v���#m�T��b2T����s�_��÷�Sln&�B�>�m�����������ޞKnhȳ1�j��q�D�ґ� �q�N��������m�<��B��=ܯ��zI�˹
��R�j����ٞ�2wu�sj��v��D(J*����`ȴZ�Awf�z�`u[0�"e�e��v���4S6�UU
f�I%�V3 o��ؠ��$���]R�Z`�U*��v��$�������T��3L{!I(țn�b��GA�O=f�_��Lq%��a�������7g=v�)t��tZ.��������yG�(���~��?~��n �5�����;7�DX������'w�� {���M�z"!/B���](T�^���`M�Uf��~0nـ?��`f����3h��)R	'��a�J%�
���� �zpt��u^�f�ޡ�hu*QJ7,�f��_t����kv��eH抪���wG<k<n�����֒C������2V�ɝ��&�#G	�������{�������l��K}X�iqUYH�]]�$���u[3ДB��u�}-�`ݳ9%���򒗔��sJ��]�{�� �;��q�"!
2#�*@U٪���	B�~��|`�V�Z+b�j�dWE���%?S}X�0۪ف��R�z�X�^��n �5q�`kv��|��? ����ֹ���?��d����mP�����OU�Z|%�-<�8#��9�ghN���5u�#,`�U� ���s�~�}����x.�D�����p�3vi`}�5X�4�>̩����Q�!�hu*QV�!��'�`t�o
�A������
��3�Ic�P`{����>�s�rbA�8�����i(<{���$�������MC5���V`�U� ��w����l�z�{4�
��d∌�6�T��9#Uaڠ]nY�r/uh	3�SȐ��g�uAӌ��!^RIe�C�P`z��0:E�zû�<X��8�Dp�>[��nـ~�V�[�g��*�ϺZ�Q��JH�F�q���~,�*i`f����fk�7*)���IP������0�0Ӻ��
���X���i�ӐBq9N۳L��[}ޯ���~0۪ـ~�J!�J�H(�"�k�W�.e��+͵[qA�F	��xC�jaeCۨ�]��m[ڡ���\��>��݌N˶뫄����k��P�����nL>$��n�vS�$��nm�<f2n�l�f]�e���n+{5maWbcZ��A�붺w`Ҩ�cn�'��.�'9^��q�U`bO	I��������P>:�����ö��O<�&{�ۣ�A�Re�� �a�7��8 u
 ͓8]~��r��ݦ�y���S#�n:��w�͞��Κsn4�x��m� z�Ϳ6�������l�?n�g���|`4�D�������[�g�%'ͫ� }�Ł����I��^(w�䨓p`l���A�����[ ����R�Z�$�]$0:E���\�tOͬ� {�{E�, ��б��0:gK`{��9A���:�A815�(��4(� �a�A��ճm�����Ԫ�կ�v�O�w/]��F�r|��eM,ܚXّ0	��E`eD�T��ĭ���P���'�i�@�i��<��'}����� �Z�<�����niF����r�,��Ws]�������Vs�<X��z�IԩE(�v`O�� �M��歘��BU����]�"�ԑt���t�����~�_�V����]�
��vy[��C�Z�]���N�����7i�:h�<�i����^}���N��?������0��s�Q�A�wN }Ʊ:^�(D�I�7f���UI�|������v��n�l�ItZ.��>������6"�QIe
1Z����7
���4����a	�kI���	�]�A�����?OƵ���;�EM�!�(�f�E�k[V�?%	;Y!�m�4�J���M#�G��I��D�٣�oC����8�O� �!���~t @w���`���+���br�B)#)U
�ZK�*�HU%ѩ�Wl1\�H���"X�ð�3��D�0^����a���'�T�DD,		 DV�#�$Q�$�Ez�@M��"3�pH�� �A���A��� ��"~��J�{�K�E�De'R�#Q�r�Т!/(Q
���N���`ݳ �^j�7*)���IPI0n+�l�=�
";���������~�ԁJ��m.�F�1��5�����v���ip�+e䣗�;յg,�q�U��l�?N�]7=	(_�>m_���߁҉6JTR�������&G��p�W����y(��O�O�+�Pr>9#�7�|��*i`f��`|������(w�䨒qXz�IO��q�>�Ӏ~�����B��X+����F �����A����ܒw��R���&L�BI]$0:gK`z��0:gK`{����wƅ��^i5Pt�j�uP��W&�`�۟=���cu��BQ:z�ڛ���{����В*I�J��b��;5��ʚX�5XZ,�#)8	�ӎ<]k���>m_�}8��u���${�)��R"L����O��8yD$�~�����p�l�6��'��a��[�VV���/BJ"��~�{�u^
��5E�B�����?N��'���j��O���w$��H�O�lΖ���Ԯ�.-������utc�Yܴ�r�������D�Vs��.x�k)Iv���7N�]q�ڠ�{��8�Y�mq�����nSgl�ywa�h����5�N��煐c�x�����L��ٝ<���.cc�jM��n-����KQ�`{2�ݺ�y''I۝8�C޵�����l�#]�����n˶Jg��۵ R\��L���D����E�ˬ�Z2�'6��F��A�7LHgƺ�D��f������ʪ�9T�_%D#�>��{�`{��3��=}���Q�]�t�*Wy�`{��3��=}�:ٞP�G�%T�U5A�e�5e�ܫ� �WzpӺ�$�_;� ��|`]��r�$Tpq����\�W^�����`ֹ�>�N�]
�!"5q�`n����s�ʮ����yff�)j3i�)9$�Ts��.����y�2�d�h��l �����9�U]���C�7%JP�,�ji`n����w�
��|`i�X����,�ˬ5�rN�_v�)�W�@���N�����}�s`{6x�>ͩ����=CQRl���(����]��a�DB���0�}X�KZS�j�	]*���BI)�y���|`~�X��L����q���9*$�,�ji`~��כ��	'����҉F}�D�,���YwZ�W�Xe�/aR<�'\�:D�i�J�������1�M��B'	$U!��|�36��m��I~���_[˪����b�U�X�;�&�(0=%(0:�5ߪ�I�-�����n)%��;� �ڶaj.��IB��۝v��͖��E:knNP��D%?w,� s�� 7u���ŀ~�͠�Q ��$�Jp�1w5��-����/��R�ӮP:�x���Ra`��{���"�3㋱��mf���z�Fjps?UU6�v���ڔ��� n論��IJ��w�]�?�+�+�Wuw�~{lΈ����|`u�`fl���H�6���`Ҩ�Di�X�W�����Д����;]��i��j��IHX���36X��vnO����<��0`�P �A i�X
�	� �O��*��>�ܓ�|wZ�ə�U�jj���=�8�o+�����`~��P{�LIJL�n�Ө��Fu�p��i�/a��Z�v��!�`�8��!�t��5$�f��ji`j�k�ʯ����=�ʊ`�ɹ8!J�l���wD����}��}J^�A8��|M����}��w�;���͉�j�jR��bK��	��~��?c}��8_%EETnG%�������5X?k� {����P(IBS�7WA۝�n�Fڷ��l��C��\����BM���[isd6�	]l=�`�=v�݇KҮ!=ki���; N�퍛�����X�f��D�nU3i`��6�f+Bܜ�s8�T^�y��l�\:V�#�K�t�Wnr�u�����v�c������h���MJ�ټ]}��sz�a�u�vv��qg����۳{t��q�]���7�~��v�xĀX5������>-nu��Lj{
�ڷ:chj�/���t!TQFH��@��=l��wD����딭`$!^!,V�lvt�;�`{�A���j�ߩ�����EG�V��^�vه��oYӀ9�Հ}��]�p(�n)%��������1w5��l�7�)���I�
�b%�:��0	�Ӕ�ֶ�q��
B��'�n�h��V�ŷ[t�u���&E��lՌ�q��o�����$�`��K����	�X��8������73e�� C���~��ӟs=7$������J��V�T��V%�0=9A��v9�Ц\���o� ����$�sst]�U�	z�����/�X ��`zr� �u�V���e��hV���]`�{������� ����~�곺R%���s�6��r��ֹ���,�n9�MGf����n�x��֫�ݕ��ĳ�������b%�:���1Vf��ҍ�N)%�����q#��yX�|�s6X�U��N)Ĉ�N�a�����c�ʢ���A��J��� Ȃhn� ro�
!/FY]���z�`�5��j�໻����D%�_V s}x�(0&�K`N�2,�3WEZ��� ��Ѿ��>��zp���;������ge;��Y�Ձ��h����:���RsU�8�%i,��G���^�6ޞe�0=9A�6"[�zg���`~��`w�U�z�*U��p�7�W����_V s}x��䒙��W7H�A�RE"�5f���l��r��}�Ł��<��Uʄ�C�����N�����-���V]}Ema��$ !a$�j���B$�"� �5T�Dc�z$\| �����nI�}�5,�V�V+I0=9A�6"[�{]�nf�V�։�ۈ�6�R����u�]�974Jv�v��<%�9i�9�L�z��J)���s�М,�������`u�BJ~����v�y�Z�*�RKb{�rL`zr����U${}뒛�P�)QJ1H�^�������{��:U[�R�����=���8�r�0���yW_���69/I�S*U��T��U�IJ��������������H&�S����2���v�k>����%����،1$h�HJp���"�8�����|����� ���~�_�6����y�(�k�s05� ��q��8�zD֜4��m��'?��
 �xUc?|�#��B	���_�D�m��4�`�P�����#�^`�#��6��޴f��~����		 ��FE2(�ܦ�Y05���Z~�j�~"?|�1"B0���l�|q�?k��`�X��è	��p�>>�	�M9O��@�
��g6E#�Vu��m�߃m����@H��m�$�m��m z�F!{	X�9Ѷ3F�7o\�[�m��X��Btn��Z��U�P���N��)�%�D4\�t��ڧ#F��Mn��C8�� `O6ܶ��#�P%],)m4�a
�C��������c]r���v�>n�iݮM�z:0���S^M�8\�vR[ɖ��U�T�6�L%����5���� 0�c<q�7S��\��:���s���{l�����8�B*ZƐř�;l��4g�G��c%�tS�^�,��I��.��)� �K��J�؊�y�/����S�L��r��^����ɴ��
�{F�8N��E���.�� �H�r��ni�2�M����v4K��h��S�Q�� �&�8��oi��ι�ǝq�Ҳ�d�sۚ��K,��O,@�mM�\f����h�S�c�M��3����e���\:�Nx1�>�,Z1�ƺ�	��cm֫��M�^���P�4�U��@4
C�a���n���:��s�u��n6�R�(�n7��u�m��n�x#i�]nG��635:(s+N���8��9x�ے�1
�ь��T�=��lc�v�˶���=\�Z�SHV���.}�ؑr��N�J�&�[ u����[���"K{3ceV!ZC��۞n�u�a�t���D��Ě9h,�YH�(�hj���L�r��[3��
[!-J�TZmm�՛��u��x}e��
�C';/]]�˲��u<�F7�On����7U�g,m5����sb��:f�rKL��Krȸ-)IiU	��'fUZU�Cv�:��lIw�Q&n ��<��Ӻ���K�{BCf[@��d�̷�m���FOz���y\.x1u4��V�=��gR�v�Ip�������\<��ŭM,�/#L\�n�c6�S����:�W ��Ja�M3Ue�R��` kJ�S�^�Md'C��MN�J_������z���ÿ�1@��"~O�?
:,O�E�'�^h ���O��}����3	2��kF���ђ]��m�ⲳ����9fy��O�<�\Vv:y��;q�.��oY�M��4N5�$X�D�I�sv�Td�����Wm	��-���-�g!řo:���ԅ�쓜�^�p,ny`3e��;�����㚼^�A���4v�q=��ppAP��ۻtѼ�n�؎yF�j���Wj�zȡ�7o-��w`-�y5��fݫk*G*���{�����s��x�X���W%�v�vD����ЪC���Lqɸ
\4�n��[�ʚ��"��REH`�u��u���<�$��G��W� ��=9j�H�X*�K}&0=9A��R����U�����}DbJt�q�Ԏ�����>m[0��8ηXt���s��t7��4�3j�:�L`zE�.V<*�+1}k�I��l���A��)A����ww��o��_�K��i��S���<�ZܞO&dޒ_',iƲ�n?���𥳐N��J�w_ ����?=�`kV�(� �_Vѣ�"�h,T����?=�x9+�Лʺ�q,N�f�6��bX�'��{[ND�,K��v��bX�'��7�ir�kW2�Y6��bX�'��M�"X�%��}�kiȖ%�b}���ӑ,K�����iȖ%�b^���̦kVfe�fM�"X�%��}�kiȖ%�b}���ӑ,K�����iȖ%�b}���r%�bX���z���&�S��m9ı,O����r%�bX(�~��?���Kı;���iȖ%�HN��d/�)!I
HM�D�~���Xd�z�9��Q�<����"��kns�<��Ԩ�՟����8�\�,�4}��oq��K���M�"X�%��|o�iȖ%�bw_w��r%�bX�w=��Kı=��!�5�us\�5��ND�,K��ߦӑ,K��ﵴ�Kı>�{�iȖ%�b~�w���r�4��ʔ���$�T��9HK��ﵴ�Kı>�{�iȖ?�� �=
0�b��J�P)V�B-�M .� :B�?D�_�o�iȖ%�b}���r%�bX����Z�R]I���K���"X�*D���v��bX�'�����r%�bX�w��6��bX��D�w���r%�bX��g����a&CD�̻ND�,K��ߦӑ,K���7��Kı>������bX�'��z�9ı,O��ad��L�u�.���63&�v^+��]�y��sA�d���5��N�� �(�I��/���G)�r�}W�ӑ,K��_w��r%�bX�w=��'蚉bX�w��iȖ%�b_�ȕ9F�$QT��9H�#��V<ﵴ�?��&�X��]�"X�%����6��bX�'��M� ؖ%���/�0ɬ1�k50���ӑ,K����]�"X�%���o�iȖ?�5Q;���iȖ%�bw^�����bX�'tw�&jY�5��5�v��bX�'��~�ND�,K��s�iȖ%�b}���m9İ?|0�xT ~�{���m9ı,Ow=HjMz]\�4j�&ӑ,K������r%�bX�k��[ND�,K�ｭ�"X�%���o�iȖ%�bt�;�=��nژ��0�1�ǘ���ݶ;�v��7K`�/7Iz]Wgh�˺"����bX�'����ӑ,K���kiȖ%�b~����r%�bX�{۞�ND�,K����kW,�Z�X\Թ��r%�bX��}�m9ı,O�{~�ND�,K���ӑ,K��_w��r'��MD�<�{�/�2.����"X�%���o�m9ı,O{۾�ND����������Kı?����m9ı,O�������um��k&ӑ,K������Kı>�=��Kı=����r%�`
�5�����r%�bX�����2�Y��j��ɬ�v��bX�'�g�v��bX����=�����%�bw����ND�,K�=�M�"X�%��8Ow~��Z�ݶ6kQۓH����<��KB��]:���T��69ca]�
�ck:6�s����r��#�o5m`�z7�c�+m��� u�ͺ%G8]�svI6I\HF��M���#h�bjݚ#V��q�&��p\��;f�\1�@S�r��d�<�N�V�8晧B ���M���re�Y6t!������[\͸�g�u��v4��=U��.`\�ݚ��߽���t�}O)nREK/u�����=bP��ۈ՝�|�\^�^��ó��L����5��e�;ı,O�}����"X�%����M�"X�%��zo�iȖ%�HOo�r����$.�>E�%XR��f�����"X�%����M�"X�%��zo�iȖ%�bw���ӑ,K����kiȟ�]T�K���HjM[����n�m9ı,O������Kı;�{�iȖ�b{]����Kı=�w��Kı>�e�I���ˢf��2��r%�bX��;��Kı;���ӑ,K���ߦӑ,K��}���Kı;�{���r�u���f�s.ӑ,K��޻ND�,K�w~�ND�,K���ӑ,K����]�"X�%���������,Л�ky%i�4P�y���Pύ[�W`�Zl�'d��r���^����3/�Kı?���M�"X�%��g�]�"X�%��w~�D�,K��z�9ı,O_]�[K�j[���M�"X�%��g�]�!���B��4"�8��'���v��bX�'����9ı,O}��m9ı,Kޝ��Zfd3Z�33Y�.ӑ,K���ߦӑ,K��޻ND�lK�w~�ND�,K���ND�,K��/��2k$&�Xk5�iȖ%�bw��]�"X�%�﻿M�"X�%��g�]�"X�%�﻿M�R9H�#����8�n:�8��Ȗ%�b{���iȖ%�bw���iȖ%�b{���iȖ%�bw��]����{��7����ߟ�E�E���74�g�ò	��]�vj��x�
�#���kWGEHh��]L�5&��iȖ%�bw���iȖ%�b{��ӑ,K��޻ND�,K�w~�ND�,K��?y�!Ӧ-�������{��7����ӐBı,N�=��Kı=�w��Kı;����Kĳ���}%6�mJBjE|��R9H�(��{�iȖ%�b{���iȖ0/ >V#�ƣ XD�U���R
�� N
~>�bfl��ND�,K���]�"X�%����6q�0�Pњ�˴�K�lO}�siȖ%�bw����r%�bX��;��Kı;���ӑ,K��}w}m.Y�.�k3iȖ%�bw�=�m9ı,O}���r%�bX�{=��Kı=�}ͧ"X�%�~��d���3/�ݴt���+��Xe-�d�y�p����%�U�8�������w5�|�9��6k2��v��X�%������r%�bX�{=��Kı=�}ͧ"X�%�ޞߦӑ,K��K�L��		����iȖ%�b}���Ӑ�D�=�}��$�w���hH����;��/�L*!I	׽>�ՕW$����w5�iȖ%�bw���r%�bX����m9ı,O}���r%�bX�{=��Kı=��!�k��f4��5���K��j'�s�m9ı,O�翮ӑ,K����]�"X�TlH_�8�!�|�����iȖ%�b{ޗƯ,3S5�	��FfM�"X�%�ﳾ�ND�,K�g�v��bX�'���6��bX�'z{~/���G)�r�wW�"S�GND�p�=��x�v���B.\�Q�b���z�\4�_}�w}\2��2柽���7���'��z�9ı,O}��m9ı,N���6�?D�K���}���"X�%�׳���I�����f]�"X�%�﻿M�"X�%���~��r%�bX�������bX�'}��m9,K��}w}-&Y�5��Y6��bX�'~��6��bX�'���[ND�,K�w~�ND�,K�{~�ND�,K���Zk2��Y�̛̺ND�,K��}��"X�%����M�"X�%�ｿM�"X�bw�o�iȖ%�b{��\�5�M\&35��Kı>�w��Kı=����Kı=���iȖ%�b{]ﵴ�Kı: zo�'�ӹ&R�ֶ[&j��T�:5�5]��*E�/\qI6|�̪�J�h+�ݸ)�^�:$Ԝ��gk�-�e܊�B�̼R��rQ����ճV�z���N9ѽ���鍙z秒qZ�y��.�..�紤�1������<����xJ���n��C���M���	��)����bM����v�z�u�5]Jڭ�-�PD>����M����;v���1n��������l��%�y�vs�ծ��q,�T�����D�?�����r%�bX��w��Kı=������~���%������NHRB������R+�wj��U��%�b{�ߦӑ,K����kiȖ%�b{��]�"X�%�ｿM�"
�j%����/�5���e�ffk3&ӑ,K��׽���"X�%��g}v��c��D�O��o�m9ı,O��o�m9ı,N���au���k,��jff���bX�'����r%�bX�����r%�bX��w��Kı=����r%�bX�~��ya�m�Pњ�e�r%�bX�����r%�bX����m9ı,Ok�����bX�'���m9ı,Oy�۫��kзGґ�ݮPãZ�9:ou��b��s�6�9�=ג,�;)��7���{���w��Kı=����r%�bX��w��Kı=����Kĳ��+|ȕ9F�Q�_+㔎R9HOw;��:xL����E�؜�bk����Kı=����Kı=���iȟ� j��X���/��.U]�6�UufB�B�����vx�9ı,O}��m9ı,O{���r%�bX�����r%�bX���bN1R��Q9�|r��EW��m��r%�bX��w��Kı=�w��Kı=���iȖ%�b{��CD׳5�.k-�6��bX�'���m9ı,N�;��Kı=���iȖ%�bw���"X�%���g\��p�.���{o=���s�=�ng�]�&���n'�-q�1��r8����:b�ff�2m?D�,K�����Kı=���iȖ%�bw���"X�%��w~�ND�,K�s���35�sYe�ֵs.ӑ,K����M�"X�%��w�6��bX�'���m9ı,N�;��Kı<���r�2�f��5s&ӑ,K���ND�,K���6��cѼB}�
~� �#�l5�������/�'��+`.�g?De�5U�6	#�
H��:�O�4�}.����?}�O��I��>Q?:s|i.�@�:�0Y�u6�I����J�0.�  B"C�06�E��7�?�>E���0�||`��[#I��I]9�$Ȧ��o�؁�
�|����?�0E~�!V3��݀���'�*~`�
�: ��bx�ND���]�"X�%��w�6��bX�'����i�RkZ�k�"X�%��w~�ND�,K����9ı,O{���K��;���ӑ,Kħ~;�I��jfk5�̛ND�,K����9ı,O{���Kı=���ӑ,K����M�"X�%����������;����:�nu=lu���<�7n9�4�ʫuΝ&t�uu�N�t&�5.e�~�bX�'����m9ı,O{���Kı=���a��O�5ı?����iȖ%�b{G��0֋�ԥ�k4e�d�r%�bX��}�j�/D*!I�����$)!{�ޝ�"X�%��w~�ND�,K��R&���M8\�[�m9ı,O{���r%�bX��w�iȖ%�b{�ߦӑ,K�����"X�%��z_\��L�\&ff�2m9ĳ����o��iȖ%�b{�iȖ%�bw���ӑ,K�wV�)�� ��k�9�6��bX�'����Z�՗5�[L���iȖ%�b{�ߦӑ,K��c�����ı,O��o�m9ı,O����9ı,O�d�_��;)�枹�Xx9���Y��	o;Y��{%�kS�l��9��n4��;���iȖ%�bw���ӑ,K����M�"X�%����]�"X�%��w�6��bX�'���7�i�RkW.a��Kı=���i�*$uQ,O����iȖ%�b{��ӑ,K�=y�B�B����+�>��ʺ�����6��bX�'�g}v��bX�'��p�r%��	D�Ow���ND�,K�����ND�,K�x��̆�$���f�̻ND�,K��m9ı,N���m9ı,O}��m9ı,O����9ı,O�w��kE�沙u�6��bX�'~��6��bX�����?���Kı>��]�"X�%��w�6��bX�'"�$ 3�B�P� ��4ւ�T��%2'~�5�R��f�f�F���4�Ӻ�����Gc6�Y�p�Ν]���5�S�7[u���e�;���K���4��u@�@����f�n�4E�X�7Ir�cEA�����mR���=�»I��n��#��z���sK�;,��;c��i�l�t���U
r�Rۺ�j��.�I r�-j�5�Í���6��K��Mj�q']�SQ#���y���՟�V5^J̹���>�����/g{u�"N��s��L�'����dɧ��Z���Kı=���M�"X�%����]�"X�%��w�6��bX�'~��6��bX�'��|MrCa�Ѭ��fd�r%�bX�����r%�bX��w��Kı;�w��Kı=���iȖ%�b}����q1��J>�7���{����w��Kı;�w��Kı=���iȖ%�b~�w�iȖ%�b{ӳ�)��e����̛ND�,��D�}���Kı?�����Kı?{;��Kı=���iȖ%�b~>�~��2�I�\�ɴ�Kı=���iȖ%�b~�w�iȖ%�b{��]�"X�%�߻�M�"X�{��?���푸�����[���x�կ�tdi���Ҁ�8��Ɯ���4]�t�5��̛ND�,K����ND�,K����9ı,N���l?�'蚉bX�����ӑ,K�����3!��!50��s.ӑ,K����]�!��^<D������iȖ%�b{���iȖ%�b~�w�iȖ%�b}�=���0��˔��˴�Kı;�w��Kı;����K���j'�����Kı?����m9ı,O����2dӅ�I�d�r%�g��D����6��bX�'�����Kı=�{�iȖ%�bw���iȖ%�b~��|MrC5��F�2�3&ӑ,K����ӑ,K����]�"X�%�߻�ND�,K!sy�B�B�����>�����J���c�y�*{n���{�>�7���r&Ճ���pԸ��t%{���oq����޻ND�,K�w�6��bX�'���l?�~���%���{��9ı,N�OO��fL����Z˴�Kı;�}�i�
�D�K�����r%�bX�g��ӑ,K�������O��MD�>����[d�f�֮\�iȖ%�b{���ND�,K����ND���F21_��IhW�(�D��_�涜�bX�'����6��bX�%>���!u��fk2�̛ND�,K����ND�,K����ӑ,K�����"X�%���~�ND�,K�x��̆�#50�5ne�r%�bX�������bX�'~��6��bX�'���m9ı,O����9ı,O�����R�R�~�ua&Md"M�mǋZ9A�Uϗv���h�&y�p�b�+�y������0��˔�\��~�bX�'���M�"X�%���ߦӑ,K����ӑ,KĿ��fӑ,K�����/�2�p��5��ND�,K�{�M�!�,uQ,O����iȖ%�b_����r%�bX�����r'򚩨�'zK�5��9�5�ˬ̛ND�,K�����r%�bX��{��r%�bX�����r%�bX����m9ı,O���FfkR�e��\̻ND�,�������r%�bX���6��bX�'��~�ND�,mS��(D) ����_~�������9ı,N�z{E8Y��Uֳ5��Kı;�w��Kı?w���r%�bX�����r%�bX����[ND��G+kw��%"��R$I(�Ԩq�A�\�W=��s��o����6�&J�2	Ɨ�z5�m2�I�\����ı,O���M�"X�%����]�"X�%��]ﵴ�Kı;�w��Kı)ߧ��!u����j�̛ND�,K����ND�,K���kiȖ%�bw���iȖ%�b~�w��Kı=��h�d5����K�v��bX�'�w��ӑ,K���ߦӑ, �5Q>���6��bX�'�����Kı>��j�\�e�\���r%�bX�����Kı?w���r%�bX�����r%�`*MD�=��m9ı,N�?�CD��̚����a��Kı?w���r%�bX"���~��O�,K��^�����bX�'~�m9ı,J���T�T��%����h�e]lW\s��1�����H1�X��	ʷ�ƺ��+O��ƽ�Óӛ��cI�:���]:鼱��!���s�p1��4�n��M9�q5�=91뛓m[�vM8��t��9��7	]glD��㰆7[rcm��қcm�⸇s�pi�ʼۺ���@R�v�k�� ���.֒����Z���Ⱦ0[tb6��q���v��If�5���^|��x��"9-r-��y�u��x��K۳6�nG��p�k`�n1$n��<L5o��{��ı=�3�z�9ı,O��}��"X�%�߻��+?D�K������s{��7�������c=�1�Q���,K������r%�bX�����Kı?w���r%�bX�����r%�bX�zv{E8Y�%���Y��r%�bX�����Kı?w���r%�bX�����r%�bX����[ND�,K�y���ē,Ԛ�˘m9ı,O���6��bX�'�g}v��bX�'�w��ӑ,K�����"X�%�O�=�I��k3Y�fd�r%�bX�����r%�bX����[ND�,K�w�6��bX�'��~�ND�,K�zSz%ֵ�5rE.�4Zms�Wg�Y2s�c�k���ղ�h�Ԝ�zn���ְ&�5.e�r%�bX����[ND�,K�w�6��bX�'��~�ND�,K����ND�,K�a�[��2CYr�.f���bX�'~�m9�SdNDȖ&�ﹴ�Kı>�w�iȖ%�b~׻�m9�T�K���CD�ֳ2����a��Kı=�siȖ%�b~�w�iȖ%�b~׻�m9ı,N��p�r%�g)�׍�}�a$nI|��R9H�b~����Kı?k�����bX�'{�p�r%�`�D�}��iȖr��G+O~�tH��!R���(�%��^ﵴ�Kı;���ӑ,K����6��bX�'�{~�ND�,K�@������j����kN�59ųn�uS[�\vv{&���\HC��3t����^,�LMWZ���Kı=�p�r%�bX����ӑ,K���o�a� �$����&��	�y��'�&Y�5��0ؒ	"}���n'�X�'�{~�ND�,K����ND�,K��m9ı,J~��jH]e335r\�m9ı,O���6��bX�'�g}v��c�:��� 	
�P���D���C�^'�����Kı?{���r%�bX��m��ְ&�55��ND�,K����ND�,K��m9ı,N���m9ı,O���6��bX�'�ú�^�fk,5�)ff]�"X�%����6��bX���}���ı,O����6��bX�'�g}v��bX�'����ￕ����Dniap��s��'f{X�Y���e�[nN�BU��v��apֳ�"X�%�߻�M�"X�%���ߦӑ,K���o�iȖ%�bw���ӑ,K��vx�3S4k�ՙ��f�m9ı,O���6��bX�'�{~�ND�,K�w�6��bX�!n�q���0��$.���JE�IW�m�Ks&ӑ,K����6��bX�'{�p�r%�bX�}��m9ı,O���6��bX�'ݝ��Nd&&��Y�iȖ%�bw���"X�%���ߦӑ,K���o�iȖ%���R$?���9^����Kı:���'�&Y�5�30�r%�bX����m9ı,O���6��bX�'~��6��bX�'~�m9ı,K������WR�I�Xd.���u�Σm�Q��^��d�q8%�::���ff�\�˴�Kı?{���r%�bX�����r%�bX�����@g蚉bX�g��ӑ,K�����S5��!���K�v��bX�'~��6��bX�'{�p�r%�bX�����r%�bX�����r%�bX���������\��s&ӑ,K��{�ND�,K����ND�,K��޻ND�,K�w~�ND�,K��S��]j�ap��6��bX�'�g}v��bX�'�g�v��bX�'~��6��bX�'{�p�r%�bX����5sF�%ճ3.\˴�Kı?{=��Kı;�w��Kı;���ӑ,K����ӑ,K��CP���B�	��"D���A"���H��*�
K	�8���=�*��kD?�	A3 �~�؁��։�5�>6� h`T�`E� FcA_���"͊�(7d4	�SB���"�b#P1�'�=��?O�Z+ߢ�7�]��"H�J�
���C��¤W��ā�h1"� m�!JmC�Y4t��|�� !����kZ����EhА� $�6��~��'�u�t��%�� �Z��<#�%����+Z�N�CvH��d�����Y)a���ˁ�.�v���:r�닒8�p�@��(v꧈na;
BR܎�sS��������;<�a��*v�&��v6�7��utq�#pO*k\�v�#�����jU�[�o�[@�.]vŅ��h�y���Ͳ�ҵs=���b��Hs��N\:瓝c8;�йU�%�ڵ��x@1Gf�n�=������c��Q��x�u���a�����V��q Pnbk�ݵfyX�mfA���d�N�j�^x�@������;�"؍�����@�  �I�Ó>�V"e��(�� �6��Ë�`�sќ��$�gN���:�|�V���[��Hy�4��Om9b�<�ݶ��
8��h����z�in��u�|c���\񝇜@j�z,��"(l�6t�``�#V��]��d�z�;;d|�mv���`(��u�J��\gg�X�ꉇ����=E� ��,����/ϵ����U�Q��b|���k��Z��*_��8����A��1�cfB��J�*[��C�;	��`e5��ف�x}B��	+�eS�&}�c\E��9��)�tmg��n�2���"�m�An�m3X��9�m*�Umҗ(Z���\�r����zn`�M̏i�6�"�`�O�NN�{F�6�Z6�����ji�T���l��I22�V�:P��S�̧9����g&�:�Su;is�Ǧ+�ו�鍳ٔ8�&����h-�UeZU���Hf��~RYU\0�-UR�U�a�cLn�f�*aڮ��=�.�E8[mڪ�{ERtnt�geLC]!$q�X�w\���9�s��d�,�u�;D���v<o\��P�]��	��&Ű�/T+�<�;B[Nď=UJ>ԁqF��:���I۵�����v��@����H�6���ֵ���sY1 ~D�!�sb���" Dj�3D>|�~@X��?!���Q��6 &wf[�4jRˬ�k-�*X�M��xZ�
G\�鋙�L��ٻv�짛nѥ��7�n���Ƹ��՝�0�{^���(,\:�:�H���lTs���ҵ�c����!Drr]�3<�g�K@�u��d69���3�n+��0��m[~�0wo��RUۻ7;��{j��:X�c��捈/m� ]5�v�ӷ<�s���m9�9Δ6���f�;�߷����!6�1�8L���t�W%�m��yS%P<��e������3Q�ڰٖ�d���D�,K����m9ı,O��m9ı,O����9ı,O����9ı,N�w�D8Y�%��f\�m9ı,O��m9ı,O����9ı,O����9ı,N���[ND�  ����'���Y���AUu7k!~!I
HRB�_zr"X�%����]�"X�*!D�Ok���ӑ,K������Kı)��4B�)��j��̻ND�,K�s��ND�,K����ӑ,K�����ӑ,K����ӑ,K����_I��0ɫ��K�v��bX�'u�}��"X�%��~���O�,K���=�v��bX�'��}v��bX�<w�\lV�Bx��Q�n�n�z�4sΕt�p:;��ז�:�.Nv3���!�e5���ӑ,K�����ӑ,K����ӑ,K����ӑ,K��k��_�RB������h����%�MfND�,K����NCA`$`"��]�P(+�2%��s~�ND�,K�w��ӑ,K�����ӑ?�]T�K��O㚳Z5�]j�̹s.ӑ,K������Kı;���m9ı,O��m9ıRB��q����$)!ky�E �&���,�3.ӑ,K��ﵴ�Kı?w���Kı?{���r%�`,�O��]�"X�%�����<,Ʉ��3.f���bX�'��~�ND�,K���M�"X�%����]�"X�%��}�kiȖ%�bw�ΓZ���vS����Ƀj�.��A��RԼ�%7�+�bQy�ۓ]�6��6�����%�b~�w��Kı?w;��G-�z!(��C{�� /�|�
j�]��Z��vt���'�`l��0="�����G����T\��F)��w�ܓ�}ݛ�������(D(!��DBK1��� �[Ӏk����V,3(V#��wGLH���j��6X�V���j2�F4�����V�?_�7����tt�����v{���"�x��;g;�;s�%�vlk��3��2ѫ��ci:�zL��
lHI*`{���oD��tt���t��<؇DQ'$J�B�+ ����UI)�����ŀ~��8z:S��Qw�]a�&�������:[ ����?$��hjB䠪���D(I���nI��w�rI��w7"�m��.��]�_VnU�V��i�I�RIMET���K`މ�������l����Y�B=(,cyB�Z��.�T�}����۝��"m�sv�KMn�N�N%lw�`{z:`{dt���K`Hea��S����Xw6��U�RGs޺�;�|��͖cժ�4ڌ�������~��X�\�Д$�d�}xf����M6���JJ6)	,�$���07z:`{b�vtVe
��$+�촕�މ����o(Xu��n�>"4�	C������k�]9zx�h[hڞejۄ�G�XŜ=�w%8	&�z�Pt��$�$Ԝ�l��Y6�c���f�	أ`���DKr8ЩWWph�Y�CWM{d�	�Vn�u��'��g2�z�J�lu�df�Wu�R��%�L�r;�B��6�n� ��k��\{nɋM�璑���{qἳn.{V����?��mo�A�'
��%��e4][ֵQ9�q.��ؾB�γ��f1�;]�훀u���Dt�)�%LTҒX��Ձ�ɥ���-�M���K�����`�g�d�k�p���}� Cn������e��Cے[ ��07z:`M�_v\$R��
���loD����7�~������y{���u���)*$b �{�u`M��$�7�`u��ee����D��f\Ve9�.s��A/j��miq�:�8bƕ��F���J�ߟ���ܒ�މ���� �q�yw��҉�j8Xu�\��[\�͖ٛu`ori`wlC��c����%� ?���u�Ô)��|`���;��W��ՠ�
���Ll���������0=U�u��V
�Ŗ�0;yA���Ӣ`{dt�7��/n�u��rƷ[���A˞6rm�^k���m�ˆ]�����<���籣�������� ��ގ�}�	�~^ּ)*q�QN������0;yA����W0�X���n� ���X���)�Z�%B�0�DloX�ל�����N��srO�z�Jm8��NB9V�&��ɥ�ose��soŀwǏR�6�J$(��!���7�`{yA�7�R�V�[��):t��(M"B�mu����*u�ǈ�p�ZBNx�����#Fz'��6�3މ����P�UU��<X�y���E�LRK������ၽ�ztL}>�W*̵�ŗ�`v���Ӣ`{yA�q�RVQV��J�eZH`{yA�ztLo(0�||}�}���'M����j����(�' �se��ri`gri`}ܚX�����&4�ͧH
iSz�ŭ�
)��#���N��8tqs�1˫��T#b��*$iTjI�͞,�(0=���=:&vL��2�`��HI�P`{yA�ztLo(_��wO�m��R5,����0=������tUx�g׉�٘��=:&������}�$���8�gR�����3*������P`{yA�ztL�ߖ\�Wm��4�ڐ:X��ѣv4�7(�i���E��÷5�5�اq�r�c���yȜN��iC��t����Ɂ#���Wv$�Zz�b�v�)l���XL��N����r�!Nc��l�]�W0��OhҶ{DuKvg��Xx;n!��؂�)4#��F��$n��ZvY��t]�&<Zsaݡ����+�ZZ����dRj�=�������{����ߝgLj�u����/u1�)ũӋ��{�[�Ӟ^&J.�Zr�i}�qq�u��� ����`{yA�ztLo(0$���u��e��C��Ӣ`}ܚXܚX�I��.6J#���ztLo(0;yA����Vؔ�B�F�F���ɥ��ɥ��ria������~~R�l��J��C���P`����������8������1�un���Y�8�6<���C܏::�Fg��liθЎ��v�Z�x� }���������e&����,�͖��T) ()	�ڈ�����rL̚Xw&��$n��J�)E(K�SI�����o(0N���2��iSQ��8XܚXw&�7�`{yA�@�L�u��bʴ���� ��0=�����l8��]���/,�;�N�ָz�NxLq���x��δh�<�][�N
M]v�P�&�LtP`M��t��L��R��K.��`{��o(0;�5X�6X�V�M6���$RA�7������+�Wާ�*�Y����!�~���ٝC�M��JKMP�iͽC�������	5��;�BSG�!�C�����;�#�s@���n#Ј��$�m)"���+�Ƹ�ً�6�uA	�X@!��x��?|~8h? ~���R,�� lw�MN|M_γF�nwzX�h��g��J�Ą�*	 ��HA�\C�Ibm �8��"U��[��~�۬��s�4�%�y���+��&����H�������p��
�����>T������#��H2I"��B H�$���� @�uX��� >t*�1d(S$�G�6�;�>{l��cRD�%"%n8X{�UK6o��{7���6iaꪥ���`f���㏉�.�V�&�LtP`M��t����~ߖ1Z�J�|��s�b�U���<��Rۮz6�"�v9
��GG��<D������f ��f�ֹ�Q�@{7���3�JR�)��4�N�X�Z� �x�v��2t�wP����:�`f����`}�4�3sn�[����R�"�z� ��ـk׋b.�&%�)
$N�QHEt��(U(2�M)��)
���k@a�Us����V�<ؔ�B�F�F��vIl�07������P߿�����yV�l���w[\����1�u,��c��6ն�d�TЕttF�WV���į�?OΘ����ꪯXl�yX�ǩ4ҜpQƜ�`wj�%
!L�s��>u�8z�g(�2kwқ�>' �!�"���Xc�VnmՁ�y���tTTԩ�Ъ��9/�B���N ��,�s����;��wM�MJ�R&�3sn���,76XǺ��V�[�BF�@%Ĭ�ܾ�M-�l�8��B����^guõ�,dx�6,�V{n�kF	�[r�z�p�35��v��@��;��a6�	��*L)i�m=�������(��L\M��b屵����(��P�M�9܆�kf�P���vyd�t">1]���݂�W�BAvC�Ʈn;`z��ƾ�qݞ�p���g��].�at��P��s��:�J�)�#j�I�Q��].��	�=:o#^k[��t��]��_�M�7}�Srq�B��6 �͖q�76��ո1k���5(�nӢ`wd�����dP���Wf��bR�
�U�X��VnmՁ�(0��u�U���QE�%l�07�� ��07�K`�oiN8%#nJ�;�4���`f=�`f��X�4z�N0q�A�-�흷��m�b<["l�$�.�M��`ku�K��i$�ԏ�ȒB�,76XǺ��07��v�u�V��2����'��ݡ��BH?"��'u��ܓ�{�� �͖y�n�餩�PJ��܎�"� ��0;�K`z�뒮��bU��1*`l��D���-��#�4�̵�,_e�H�C ގ��np��X��0P�Ki��[��$�۞��mTg76�YݻQm����u��K#��nNv3g��ڐ뒗��?~��"� ޑ0:g\�I%I`��Bĭ��#��P`��`w����'$rCrO�w;7$���sr�� ��"��'
&!,��%�+���X�mڦ�|nD��!`��`w�;�07���e�B
³I0>�np�Q	k������ �[��~y�ǳ��V�q�V9�[i��D@�MX�u6[���u/@W.Q�a޼ι��u�%���:`oE�"`od���g�*7%28)*��٥�w$L	�%�7�t�&������
���;$����^���J�J�Uv�`N�-��;�rN���ܘ)�$"ED$���P"��B0 ���,z��\�T�e�]��+`oH�:(0�vIl�Ձ��Ăd�x��]�mc�s�&��E���VB띌��m��ůTכU]�����~��x�ny~��݋ ާ֦���J�����;$��]�9(�S'�ā�$��`�UDݦ響[zGL	�A�oH���k��"f�Յ�us��%:��,�_� �n�q��[��"*nNݥL	�A�oH��K`oH����ww�~��}��\�g�:�"������O\�[���BM=v�i^�eCe'�m����ĵcRupu��]ϫh�'_���[}��(h�*�2�x]��Ͷ���.$���ŷ��Z��F�y�,�D�D�V�m�N�=�9^��Qf������o8��E2���ۃ����N����[�mt˶�x�Ӏغv�	��\�z���[���$�����ȁ@A�	��w,�.\��a.���$cs��(���1`�Kq�skm���H2�v���j�$�6�*�à���7�`oH�:(0&�t�.� ��K
Uv�`N�-��#���7�L׏S�j2R�NE`w7n�͐`�&��;a>�e���ZKT���:(07�t���I��$�&�,��,͚`kx��ـy$���3=A]t�Pޑ-ny�Xy=T�:���ݴp��홌��v��s�R�� h�c�e6)'�{}<`kx���пH�� 66Qt�k�&\ɹ'�ݛ��6����Q5�!��H�i@2"4h�JTB�*I}��]� 7u� ��,��n�����8F��`nl��3$L	�A��GL�2�`�#3]+�0� �"`oH�:(07��ZJ2P�uR��X��;�:`N�zD�����ĒVl�İ��<̠�u6J�/��{xv�; t�&�4�����ԥ*S�H��X�۫r(0� �"`��Z2��}�-%�*`N�zD�'H��:`w^l�㎐�I!
) �n� ߻���O`X�Q 4q �3����M�J�WR��`��¯I0	�&��� ޑ0�~酪��HZĘ�:`N�	}&0��`|��"�7C	C�
�^�`�>y��+�z}�����D���rg��q�h�I}k.Ҧ��7�Lt���#��	�b�J���J��D�'H�$t��r�eݪ�Wa���E���d���� �ݖkǩʃ�J��R%$��UW'{���9�������S1�
YTs��]��� �t�(45)
H�T��t��:(06H������K�+ױͻ>u��6I�e����q�g�b�������ێF�fx�`ۂh��� z�ͼ]
!~���e�ܺd9d�t�U��f���ٜ�!DL��ذ��Y�kw�2��Aw���0:~����0�{�K �8n�����8�JJ��+������:~��b�zGLY!w(RJCndNU�w7e��\�{�;�2I��_�nI�����������
�*��"�*�U��TW�EP_��P_��IE�BDYE�PDBEU@T$QAab0DX$ DT �"�b�QE�E`DX$Q0DX�DX�D@�U��UU���QP_�TWH�
��UU��TW��P_�E@U�UU��TW���*��P_��PVI��J��� sd` �����]+�4�   �(�  �(� ��� 
N�
� P  �(H	   )E()UA�PB�%(��E	R�FP( 	*�  )B�   �
� U!p    X@@	d ):R�bh���������{� ޔ�۳S��Թ�M\ZSۀ �*d�g��x  {ǝ^��� �Խͪt�ח����{<�^�� �zOUL������� �   
F�9h �`N��I[D_s۾�� ;K�mZ�i����Ի��Ҭ }�r����*���  ���{���zν�� 9}�>����[Ϸ=����y��|[�[� t��֜��η�;ͻy�Sͼڥ{�>    D(({ }��Ϸz���_Zrz��o���S\ z3ԫ6��95�+�n�����7� {ޚr{��ם�� Z��ڼm�����Ƞ�O_Yr|�W����]�ӯ�j�^�� y����Խ^n_=��wK۽���W���@� q�@v׺�s}J��������sn�p �l9r{�������^mɥX tn�m�����嗀{�;v�]���^< ��W���꫗']}<�{m� =/O�ũ]�s���mK��J� }���  ���	��-�Ju� � �6R����r��,���.��@�  4�: � ���)Jb   � �R�� Ҙ��M(�=�t&� 
l�)F&�)L�@M)@bh  z�����   ���ڙ�JR   ���R�hd`	����T��UC#����J�iR�  �A1JT�M=C1LJ��_�����E�����S33)�㶡����HEQWg�*��ES�������*���TU����~??��!g����M1 ��@A�����6��ɢ�v���}�����-3�B윗%�v��
m��(aѷ�>SCFߜ'�8�5���aq�oS)
�����������ԾJ�ƾ��ㄹ�N#L0�$P�8ɧ�$�ī�`_���ZH�}����:�^��%IB$�����!e�IM��\d��~��̳[3&t�Z��1s��'�|'�e�3f>�y����r��2@����s3;$M)9�h$.���I�i��Ü�	�ܼv?�|�U����UT��Ȩ�IT�&25e?1�!�3dֵ��'HR D�Ĉ]!�"�0)�Xܙ4F63�{L��c
as�F݌.2�0ټ��%�#pe��q�LI�5s�������3�\`%1��k�%q,�!Cd0ք�p�[���
�)q�NI��J H���Ib�0� E!	$qL`�B�7���ֱ���\K���R��\S�5�.u�H2딓?0�ve����]��_��@�@� ���4'��lK
�0���!j(La�cD�uJ��)$0F��Y�$"BVIB2#	 ���HT� #Jd%��Dp3 @��!rI)�De�LE%��pg$i, ,h��,�ٳ.�Q�9ِ�$a!Nl�q5��[�D�ӟ��4�
�-H}�,+�$	0�IB��(Lѓ0�!���G�]Gdٵ��3N��@�2�v��}��v��
��
˭&�:�aLBȐ���;�>�uw��dҐ�B��轹�B$�c�������!BY4�ゆ7�J}��QN	�~i5�Ā)8C:;&����N�E��˙I����#�B4afF$a�R8��`aH�HŔ�$If"\�'��M���u�k_�`, ��4F�҅�\6}�A �h b�D�B ����ɽt��Q\����.g!5*ŋ*�[�3�o?c����th5���a!B�q�m�9�!R�×��Y$��%�HC(Q���
}�i������b�pNUy}�H���uX|�J`ɍ$XE���4n\$���p��`�,Ü�"g3�Jͼ>�20B�� K���pJ�]��&5��>� F���o��O���;�\�u
J�c;ޱ	�|H���'�y1���Z�����#�6q��-R���S!F$T"�)#�H�H�D�
�8�de��bi�HT$A�dIHB)H�l��-a��X,2B$c�c�GV�2Nl�9��0o.���&�a�rB�2�@���ɣ{��,��vprł!xu�]�w��~�4ԁ!"1����t01 @���!#F,H�Jcy�.3���86��D)��C� �;0����Mp+;�޹rC�+��䆵����of,�ѣz8� �0p���zƄ)�����2�51���p`������h�ތ��2|��X�.ز5��`�D�Û�%�+a]B�n���P5ް�4ae�&������3���5��jW3!
�v���L�Ή\F�a��$"0�rd���ZL����ɋ�g:8nF����˖��"��z}ڄ҈I�HJ1B�``!��	��}��sfy��c���~��܀D��?j��F��&1��r1�]u�ǋ3�S�7Y��թ邥��v屄pe�5��8gym�s�,R �.p�Z虆���(�L��d�Ȅr��o�HK��ktap�#.S!��\�_20'9�8�9�e�d��b�'��~��FF9�������.��3�y���B6�xh�sZ0�X�ޡF ��I"��_���B�cX:�8;�&O����)�#`1��!Ja�$
RLX�P�
�d�η(o{7�MF�1�Q2�_���*�;��Y|k��^�f�E_����R���ͻ$�Ce������E��I���ڐ��o'�IM0��ξ��ƓI�2}7��h�>�	�w��Ø9~fA��B�M
�:�jdjd�GF0t��b$Va���X1�H�
c&Y�<�6j�$vF�!1�G���hH	#X�b0t�d����X��[#�Y7��d���?$i�:6|`>j9�2g6����a�\1��f��q��kntl$���n\c8�Ż�c!M�\�X��ƍ�t��4gf��$.8u���1�@��8���p�bSa�@���Q�	�I+B�8uM�g�B\�z���cB�
B��D-Ӹ����7.�0cZ��5
�ܳ ��HKK�[�N�Yyc&�$�?_�P����u���ʒa�G��
�������Y>�c�ۦ������� �4 0�R$,R9tE���5H���aZc!
`�I��,�0Je���� �!)��X1�$��3a����� !�)�q(đa#X� P����|�ɩqs�Ra�����5Ñ4}L�1(�.�K�����ɽ��ia(@R�EQ��"��M4�	w������S8!Lcp+,B:��>��P��Ln��G]�����(H���L�ɒ]��392n��B4p�`@��)�1)
hb�N'1~�	MI� �X��O�	����`ِ�}�K�a�:H@Ʈ��u3 �; b4��H$!"�b�cd��!�^��n'�h�1����pı`��>bD�	����Da'��L_�P6��H�e�0g�$$$$ȑ
H��I�Y�kI
��+ �a\�P+#.u��֋�w����	q�$� i @ƍ��	�Yq�����vi��X�p�e�B�sd�~0|||0�
E����Z�ㆎK�̜�7�0XȄ�	�)�H���y..����%`C�	 `��	L�\h,q��y�pS]N�]��Ϲ��X\k��>�f�l����!S	0��H`�p��$*`B�
`˔���\3�s.}�	4?�?���5�gX�p���1l	�0�
��$H��+@�C1)5��ˬ��n�>���z�״�wy�ga�b� VH�Lf�#\�kE9�k�ɂi�$!L�0�!q��H}1f��x!l�� 11�Y ��d
Ȓ:��S�q������O��k���6��7i���aH�4`�!��|�iX��څ_7J����;�3���5q#%H�C�]]��~s�ϿCy�1�X�~�}u�$��9����3��D6D�rj�&%��ύ�ĊWS���.�`&�D�	\��8��\g'�#�1
TU9G��XΘЗC������BH��J�cR4����j�M@�����@�+�1	Il�B)��Z"r���Gn	8�hU�i��KH@����h�H�R�
T�B�
RF��"Ҥ(Q�+-�de�eŁ#�I�a��r�I��!!	HcF$`D�$H�I!#4B�H�� ĉ�B,��B�jR0��#a�G ����BhdHS�q��m�+Ja��ԛ�:�c�)
B�t���]w��Muڋ�,j�5��k��.,6f�6d�>4M��"�%RH��d���{ο$*��B�"�H��6�dX�}74k0�䎵��e��?
ssc�a��B��`A�:�!��q�2I��3�x~�0�۰�ʑ�	!�����!
�l�I���}rm��;*��թI!�[��� K@�����*B|P���L2��IB�ĮP�2$"�a�\9%0�%���5��U���4�qR��;t�U�1�gY I�0a$b���B�ͥHC���3;�2�J#��7�����q9s���0�"��A��b�f��l��;�)40���L�e�,��2�a�$X�HD�@��P�"�X0H�#RQ�T:HAd�H�0!*AX��#	��d	A�!8\!"F�$�'�ܓ���,� j߳�f��S�!�h�F}���e�s�B�)
B�ư�E��c{�~ַ�w��i�#"E�1�##�D&��s���e%C�&�H�]�{o�~� �       -�m�      [d   �� t� � �@�kh     -  lm�   � m� [@ L�ν$����$  m�pm��� t�-��-��LJKUT�*��PJO[`j��x\̳q:��v��V�xw$╫kk��&�m�h4P��)���J��m�5����N�d���m�Z$�8��m	b틦�[T9f�����h m��-[B�m6�d�H�g8eֶ�6�mBK�k@8p��88,���ŷe�r�[T�� p��N�̘��lm��z�$^'JmZ��||t���	 q�J�$I �m�FջkY mm m���x6w3V, 5l�AP*ҭUJ�*��E�6� Z�y�lڵ�&�pt��۶�[n� 4P�n��6/�U�>ј8  ��hI#m׭l� M�6�`v�m�@�H.�r�m��M�6lm탆��p�� �U[@l�V�[R�A���up�R�HN���n mb]6!�̶J�Y���l�����ۭ���UڪL�U]UU�3�<�:A���S`�ꭺ���@R	�����mUR���!��Y�
��"YVP�T�fʪ��Q�I,n�X �$(�A�ʡ��W+ss�Ƹ���;�Nm��l�h�A��P��qm઎s��
��5�<��Ö���W��e�n�Z���BUiU	]���t@Fl�uۇ���9��sk�8駮����T{4hx������M���%Rަ�j��ƽ� ٶ  -�   J 5�    ���   @[Kj�۲�   ���Ͷ�@m�� ���]t�L��ҕ�WJ��\L�Ѳ��ۛLn%�p�a�Z�   �UP��Ԛr9-��VW Hlm��rIl���ѐ[dֵ����g?�� ֶ�$	 J2=UT��*�UtP Ku��4PY-6�t��lm��p�Svk�[= Y��4X�f�6�b�lJ�M���H 6�h��l!��6��[��e�5�kR Ά۶�(�k[��D� IU@uT���/ �@U� I�r[��My6�ǖ���"�6�i��fyjud��ʆ�V�����6�׃6C8�ca�r�עc�s�tl�ӫ��*�ڰ�lF��FIm�m���Ԁ �ZI��p:E�v�۶�;v��� 8  YУm�h�-��۶� rl�½��Tp����,�nÂ�i7'��|��8u7U+�Tu�/-ژ��ZlM��e���e+S�*�:�)y����ݪ���
��u �2c-<�@5R��l����ˬr��[@��ٛ��WfTUj��V���:psc�&I�I-�"�D��m�fE�d�^B��]���K�H囪��
�E���Wm[� 8 �j�uEU��*�($�)�޸I��&��%�H-�  lvj�Yղ�Uu[R���5���t�m����m#�i��\2u��HvƅCv('ꜙj�F`:���q5)@s��s��t�d%��UJ�Pm��z�\B�A@Hv�oi����M/i�3P�`'Y� I�V�H�՛�`m���[bi���Z�m����Cm�kSm���ʭ����� �Xk�R�Eڄ�M���VӤ	 m�ڀ�� BjU��W���!2����UUT�-��-�޶�����۫`m��xm��h��]6���`�P-�n��� 6� ֈ���m%F��Z�8-�H   �> r� -���Q6�m��SnU�<ٲ��Mƍ�ӎ�R۞�Mv��B�[*ÖUR�@*�*�P��
c��Zm]�m�lY�$m$�qmq"�[Z�4IACj��6���pOJ�vp�m� �m� ��h ��m�Y.$: yPu7mmUR�s��;n Xg   ��r��$�h�6�m�$^�`I([v�:��ʶ�v�sj��vsE$$�������:����V���i7 �����u�445�F�:��yb��OZ�m��^l�sl�'j�pdk���RpsU]��I��Q�ņ$��%��m{���� �cl6H����{�*UI��N]n dֳI�n	E���6H �z9&�%-��Kz�8� l:I�Ր*�����e�*�T�9$�e %�� �m���Y.cU[Uy�'9$��`�$N�m4�`���m��k@6�m�l ��@WWA�U esU@[]i�y���> l�����lI $�-�j��� Ml�o� 	$6��FY���]��Uy[7a&�9l�u�	����yp��VS�j��I-��h  >$��~�&�Pݷi�ӣ��gb����e�:|���U�m�k��f��:���i�úsΘ�r�R��[]!@6����׻�}�H��^�J��m��\�T+��Ppl+D[j��R�����3�`�2�Kl��������嬅A�9N�Z�`ڀ�vGJ��5B�)� [s#i��			:����UJ�ɺ��*u�lH� ���-�z�p$�^� m�  �E�oOmr�8��' ��j��sb�,0�%��cqv�%� �H�I���!R�*1UJ�ԫU��]�a�		�#^�mm�    �  6̀��� VԒ�n,jܺ��l  �@o��� �۬�U�z�r@ 	($lr� �H m�8]6 8�`p���   ]6�C`~���Ί���%���Y�ԋh� ��I�%�m%���v� .�Mt��m    ����%v@�]�,��Z����'Z�����h -��m[gIѶl���m([��^�4�&�fI�IUTi▹�-ҙ)V;rN�Ԡ[@pB��Wg*�k���X�x���=�r�ޖ^Wq��l��R��uJ�+�5C��l�{N��������Hph�m���6������A��j���e�    �    [m� 8 m@   � d�6�q,�;v��\�a�l���8$m&���	���mpp�Y��           ����@ $k6�m�$ְ  p9"�  [@  ㍴�m�q�t�6����`m&��c�L�x��$!z�sB�u�=�x�mV�n�YC'+��ҡ=���J�s�wX�V� +j�#[B�H��g����/m�@��#v�l�8 M��Xk��  ��ͥ� �f�Hֵ� �&۱�ڑ�t�E�#rkw �c��s`	j�Ul�  �  t���ַ[I7mٶ�l��i;�im +F�.�ۀ[C<]�C��['P-�[�p��gV�A�� ���s�I!mm��]Wm�9h�E �g�[�ѯ^ܼ��%T9٭�ں�	 ��@}>/�-��@ H۶M��v��.�U�����v� -�m�psm�HuQ���� �Ұ'Ko�-�;;HJ\ �   ��V⭕eLvj��l<��+ ���L�������)�eU�aV
:�B�킐%��5P�qI��C�d�m�Zղt�ΐ٫vX,v�@�]���v�k���x粍UJ�$���n���Щ�-��.�t��;m�	��wm�c�8
�-�˦�����iy��i4�Ӭ�D��T�v�[N    -��k5�m�k&�i'�: 7k��m[A����m�$  [A m��on)e����`�2M��H�i   ��[@h�/�ۃi�0md�rޠH��8$m�z����%�6  6Ͱ	 ͑vm���l-� $E�   	�"@ H p     �U�I      &�[`  6�[0U�#n
^]�L*�)-�*ѶŴ�"4P �%6�m�$H��	 �@� ���� 7N&�[&v��$ ���   �@���_i�[d���4v�/cl�h  ��&�� <�I�D��dl�.�I�F��L��Z�SUP���1z�p�t���{ &F�������l\ �l5@<�$ �t�+p֛2������NvUj�����6
Y�E�N��yzx�J 6��Khn�Wm/J   � z�  ��ݬ����C�['1��[l h�` n�[A�� �Hl�  �l   ,7$���v۲r�	&�/Zm�[�R��A���fZ �hi�V��5�%�h�-U�TܰZ����P6�t����P�	K+UUp ��K�MvL`� ��  �$[N[FC�$���d��O&�&ʽUn�����e�m�c�Zq��4-�kE;R�&(+����à6̓���|��zs�h�6�N�E�G��w{������"(�h@�����pЃ�U��&�����U~UX��O��(^�"�"�H 0���t4:�>G �` ��׽4��AM(������dX m ���A�	�� �|u�"0)(@���P�������:G��+�D���8(Dz0��;V��a�Q0 <�A�;~R(��ҢA2)� "w,	BE���y�E$*����~:�Sc�")���D"�$#B��T2� ���%��N�D]&�Ĺ�� ���E*�(��:�h8���*�]�"�v"��(� ۀ�A��@6�~�"��:�A0d ���P�dp
������`bZ����´�a)��$C*�ɠr*� ���Sh� �dvL��΄�JX@*� ���/0�bBA(�!�
D�|�mM��L�	��L��F
�R ���t��AB�˅@ɡa� � �E�H r �"�)��F��t�h8�1(����&D�����ǉ�`EQWH����
�"�AhaF
U"�TH	{�8�9m�N9 zѶ��� �UX :���1U��mr�Q�t�^\gZ(��Gn{��`��li��8�ʹ��L�*��l�`�Ӫ�U#�%�(9��e8���L9��dt�ja�I��dI9�^��vz��g.=���tr+���Zp��K�>;$v��!V��[s�5�	�m��K�ݝh�ۂM�l��^%YgU[s��e���C�f&���+�r bcE)NM ��a�Ãb��z-�0.;6�At�B����5.`��a��N�絍je�S�9�&�CQn�I�T�r�{Q���y�{z����v
Mؤ`gq�; ����čI�����4�4R��$�t��ґ�ZݶB	��T�[9 x{sUJD�gL!T�%H{=�,���^.�9�C�
�i�!�!�չϺ2̫R�k"�]�楎��Wd���s�����-{];�Jk9�Ʈ9کh�p:�r.�M�m0S�E�Km�N��k��YE�v��,����A�&�ܢ�d����=�KZ�v�p�`�Hmqٴ�nwn��G5�(6�{���H&d�n�HmD!y��N.1�6u��S���=���ڭ�n�7@Rpr��ݚ54�ʷ�Vң�:ݡYyhz�*�vMr�(�B9g8nԜI��۞e,':�vV��q�I���D�m�5^׬���e�qu]�v  GJ�2�L�ڦ����.�L�Z,q�P)@�Wn 9j���l-��ՑM�� ��u�i�e������/<%�3qͮWM��v�2�H7!��Xł�ۓ���@c��k�nl�÷�bͭ��һ�pA7�#�j�-��֕K�	@�"��y�)c��H)pq`��f���K�fj�Ѷ �E�m�w����I�p��
�9�$9�k[�)tK�1��1�ې\[\R]���6�
��^��jWZ84�-�Lװ��&�
�ѫM�;l�i�vW��k�Ń��U�j�F ���=n*��DgI����~EAү���p)�خ� ?#�l���G�4�6=���绻���+��h��Σ�xL��[+��es�u�!�޳�&�glW2v8�2��ݎ��yKny���m�8t�����&.��NUye�v�Uz�\by<�F��>���ym�������m�
#���.�95]�S�w#ez��xVx�Ha�qGع�r�'�B��Y��<�O fv��\.��:<��M�c�IJ��3ɛ2c8�p�i�m�j����ɷ=�9����EA ��wa�.9�����:�:�ֵ�5��;�$�H��2��H''9����=,K�﷜_�&q3��]�'�q��E�N�ݶ��X�%����I�z8���'���	��%�bs�����bX�%�q��a��&q3����d��)-n	��Mı,K��ф�Kı>�;�&�X�%�{��15ı,Nni�_�&q3�����Q9����W]�0��bX�'��w��Kı/y��&�X�%����I��%�bvs��L�g8�n��n��T�X��n%�bX���sQ,K���u٤�Kı;9�MD�,K���n%�bX�;�fc�3`��U���n�/V��mǒm<H.�ہ���B8�X)�6y�(�:9���[�����,N���4��bX�'g;�	��%�b}�wzMı,K���bj%�N&q}�S���ʭ%Pi�L��q3��bvs�0���E��RJ�X���JɄ� 3�)L�S#�5��V%%!��\�+(�S
aU�
�E����K}�~�Mı,K���bj%�bX�>�4��bX�%���)$)�%3�f[���j%�bX�w<��n%�bX���sQ,}D�N���4��bX�'�}�	��%�bs�1�Lkn�UJ���㉜L�g��,K���u٤�Kı;9�MD�,K�睺Mı,K�s�sqkr��jrZqa��&q3����3��Kı;;�MD�,K�睺Mı,K���bj%�bX�U^ߟNݟ�v�	Zۙ���/9�մ�&3�n�$�]���+������D���4��rm>�bX�'���	��%�b}��I��%�b^���MD�,K����&�X�%��Y��s3��9ssq��MD�,K�睺Mı,K���bj%�bX�>�vi7ı,N��FQ<"b�"X��}<c��rc3���7I��%�b_{��MD�,K����&�X��T��K1;�MD�,K�g��Mı,�g˷Y#��
դ��qa��'���{�I��%�bvw�0��bX�'��;t��bX�%�{���K�L�����Z!ʡ����q2�����T+!I
HRB��9������,�#����-+%�68jKv�s������|RY�jz+[]�%@&���e#���׀���:��ŀo۸�����ݏ�J���ݖ�Ւ4���i���)���rZ�\���ڜ��_n��?w��7�M�����;�m�섪
Kc�v�0;$i���)�n�߾�%Է� `�TZ���W)�/.q.}�'�X�u�D��«yX��`d��`�-��$i��#L.�{�����Y �[�H�\sr��c\���F����31N�y�P�q�3�Y���<�+�Wu�	'���$i��#^_%����<�f���ºW���F��4��͔�7v[3UE�lv!ʡ������>��0������X�{�H�NPjYB�S&���`j�`vH�V�F���ӕ:�����ps��9��ߗ�wwmXy�X
�B$��0�C�JS�b�D��E AB1rB���a�qkC��w㕱�E�շl݂���k������:�,��a�Xմ5@Utp:�vz,��N����l�u�Uٺ�9'�O$��Ms�f��	d����p95����.;�G��Ƣ7Yr�r�b�.�g�ch�	�Հ���챸y�� y�:;{�nм�^����y�-�s��Co9���l�a�tݳ�:\=]���(��=M�/D�GێD3kF����=���Nֱm�u�'��n×��KX��2�*'*v���}��4�ɷ����.]p�T���ʰ��ş��g}�� ww� ��w��:��e�R��KV�n7e�5d�0;�4�7kW �;-REb���M�w� ��{������L����$�a]��v�Ւ4����&�n�`{�.{��O0RQȣ�r1е21z\v���in��^���4➭�ێ��˵���9�s��8��]'��&�n���v�W}�X��I"1�-���ڰ�����*F(n V �	�i}���w-�li�ݑ��X�9J���Z��7e�5d�0;�5�}��`'����NT�Q�p=�%Qo�����4�ɷ������p�uAIl|,� ���X�}���w}p��q`i���+�+���M�tV��3�+3�M��"�ŗ��k\i`)[c�[,��QVIj�>��07e�5d�0;�4���W8TU|�U4r�(�p��>^�DD��nڰ:�q`on�Wgxےl��ՑG-����vF�_g�}�%������}����V"ڰ��ŀdۃ ��lY#L͜�8�T�v��YUwi��n7e�5d�0?wwި�\�x	�t��Ic�Q�l�dۜ&�Ao#��A�Y����^������V��g@6O[VH��.�p�>]۪2�j'*v��W۸������:��X��Xs/a(�����A�Kk�eX��� �{t��ݸW۸��u��6�-"�U�r�M�0ݖ�Ւ4ÿ|�_���|�K�\_��� ��� �;-Q��a|��f����v\6���������QtnK�s�1�^�۳�^.��mlE�0��h�aI����ݰ5d�0;���ɷ����Sَ&��V"ڰ�ۦ{�����l�����f�s�C�\�E.W,��X�ɷ����F��t�;ݲ7ѫ��l� }���5d�0;���ɷ-�(��+\��]�W.��F��p`dۃ ���RM�\
�b��(E�J
\K�B�����Z�R+�3]�B������ͫ6[@ڲ�Wek]�O-U����Ip�!��4i�����A��kS��Ogv#�=uЄ֝؝c]�c]98:��<A���91������=��6I2]�v�ax�,���^y�k8���[��K@��jݟMj�;�n��&׀���p�m���v���e�N��r�!�4�f��^۷�w�x�{�w_X�{.� ؑ��e��ltuZ��iґ)��U'ӝq7!�r�e��N]�|_-h���ɷ����n,�����YUR��%0��L ��lY#L�06���_.�+��_�7e�5d�0;����{t�:�:�q��Z��(� ��cL�02m��f�f��u�W	`KEb-� �ݺ`�s�������W۸���Z��;��#��*�sŧ]J;G"�s�v�k� H�y�㍛�VDVԵG(ݔ�>��0��n���/%�%����� ����6�J��9�f���s���j��4)�HIddDD%ޝ]�`>�`u�`w��-qX
�j�[�u?�f��t�>��0��n��n��; ����W|`we���n7e�5VI���Sl���Q�J`on��q���=n���V�P�Fo$j��ۜ�9��9ƍ�Ә�zm�l8^g�M���K�u$�$����'3զ�[cd��5VI�vF�6��ռԊ��e��Dܶ�O�ٞ\�g���`����ny&��S�����+j�����&��J��ۜI4�P$>�0f�!1�Lc8�$i�IIRR|]�B�c�
b�{R�W<���.%B2!�È�p@(�j�(�.�� E��H!�v�'�5#���5a��R%#�f�d��J.H�T����"����?`�0�`�3��	Q�ZZ�}p9��Ype#���M�.���1���y�B0�%XF>v��ٖ�p��`!�vXw=�C`�9͙ț�.9��bcE��fQR @	�H&���Fw�	�������*����$I�-�H��E���h||?8p-Sy}�:p+�ڝ���w��*�D"*��mE���3���] �@��}����t �6667�=��A�lll~�}�co3�`�q�.q��w{��Ѓ� � � � ���΄�����罝;�������hA�liĸ�o��)᪢U:������]o�ͻV^q��N�������.�k�5�5�+Wnӿ��s�ma��A)}vL�]��}q\�}��~��쑦M�0ݖ�ߤ�Y�*�×w\]��#L�p`�-�u}�s�s����Һ���FIj�7��0͖�Ւ���H�w�W#z�-Q�b�����ۀu}�Lw�5&��T�L���`bL\ľ�K�3�0.Τ8ےk+�7-���W�S����~n���������e6u������3czx�JW�m�f��[��ۥŝ���,d�ԋ�l�02m��M���\�vIȬ"�:������ 7�[VK�l�07e��qT)Z�V���,`d����`dۃ��ו��S�[-�:�ۦ���&���ߤ�_+���U���.�I`y/�������5f�0�֔g�[�F���.�����Uq��[=Vn�6��7.���2RQ9����΅����'XW�|�>|��Ʋ�)�m�ϱ��9�kg��Euv�K�]�H�݉^���&�+tu^[v���
8i�gmf�)�Zmv65c]�.u͓���a���q$�L5�{s�;oj��jU�j���^k��\]v��ʁ]M/rfa}��M�	݌"�����2G[7�s���,S9��%���ʟbg���3�<mH�׮�O'��nN� *��-#�5$r���]0�ݸW�t�>��X_N���j�K��vK`j�p`eI8�ɷ]��n9��Y��[�u}�L绱��nvK`fj���WWG*�Wh�X�ʒq��nvK`j�p`��$"����l�>��0���>��i`v[u`cTNL�
dҞ���u�ۜ���v�+�_��q�����yOf����CU��tj��N�e? n�� ���X��y(J���X�پ#��Eb�ڭ��_m��8�ge�V7�Xc|����n�I���p�喘_��}��a���z���� ��m�6�-#���r���%�5d�02��`���V�e�5-,� w�� ��n��wf���w{Y5J+K$��XZ���n1y�G�K�U�c�����D:ƈ�sg���r9\���i�[�u}�L绳 �{t��v�}���P�V�E��'6��7d���7�$�dVT�P����� ;�۩��P��PF�@9��4���"�ȨdO�7����u�ޘ{�"z5`r�U���ow�Y������g5ޖn�4��ʬEU�m� ��n��9�����|��ŀf7�ы2�U2VԪ��u�v��m�m���v�;2Ȇ;Z]��r���&�ܱQ����'�-9e��o����2m��f�~K�o��<J-s����UUMrl��/ފ�{�r����ݛ�<�����~E���t����w�.�2͈J��[�`f�i�j��7#����Lr�qs�W}�,u�6^q�	$�D��IRP��F�������I�t��4`�1�J�j$��f��=�nx�������0丗uxy9���t%D����9�۵�׫&A]v�1�%���z�������U�T�R�_�;�0�����~aݞ��7I�H����T�S ;����F�y����f���2�2?�+�2�'Uu[m�5w���f����~�x���,I�3�5(*h���`f�J`dۃ �l������ʧ���ܥ$�����L�ʱ��5?sŁ�k��P�B'��[iO�91;l�%�&���b�aG�6�;�ܔs��cIs�vo5
dg�h��'��yP��p�N���GZ��NJ�u��m�:���wGFG�m	u�/�Nx	Gh���m8�g�ƞ(.�t���1�7���]ƍ�+��Dnn^�*8�c�8e��&��9Vɩ�g��;﵍О*�x͝(G�`+�W�u��J���Z���HET���K���tN�*�:�r�ٌ�uc^|n�Z����C]�PE��R��3������;-Q�b���������n���~_�w�|`g����X�jy5�X.���Q�F:�M����`����9���S�(�%RUJT�r�́לe�
L�Ǽ��w��׮6݊����Wk��K��\\���~�,��.�sa��DD�8�l��$O�UD�u[)�u�ݘ�8��j����>��<��G��������7�WE��#�g����j׫��q���s�>�k9�ė�f�i��l���շ��o��������u�$��{;���6ޥ�|X� ��ն����m���TB�yj��Ȧ������
�D�A.��e3�G\���>]y_���3�K�m�c��7�m��C=�$�ow[x����ܥ$���~m��_m�}ݟ�?��/䕷�����}����6�޺��-Q�mE��ߒRm��~��z������_�Ϳs���~������"�ؘN�O���>�)�����}���6�}/�����wg�ͷ���h*�G��S� �i�5�=v�7.^�+��s���r-�6�w���o�ﴉ3���U%�~m��}�?~m��]6��}ݞ\������ئ6�{�?8�v*�Aڣ���6��.�?��$��������m�?b��o�ۚ~��s�H�I�H�U����eն�c��7�m��;������!򮳬���M��{�g�x�o�;�Wn�'UvY��oˉ �:k۳V�~���o��{n��U�9�o���oR��,s��Ie�[Y����uٽ�o��u�[�m��;�ov��wEմ>�7�����3=st��B��S;v�S%H;�[�H��$���<fv��{�|@��3Q�]$��}�m�m�x�o��vg�����3˟�m����6����~vZ��v��Q�m��۳��)#��f6�ﯼ�} }�� �����aa;?_�o�m������m��u�m������m��6 P%NUJ�r�m��{w�m���mն�c��7�l`(h2`D���L'2f��$�#�~ٲ�u4�/��5�٫m��N�ln�Yh;Q\�������x�o��{=��;���+����m��6��W���n۱m�ڻUP]�(:Tǜ&�F��	�M\���{�l�\�\]@���Oߛo�m������m��tx�o����[�D���?~m����1���w_�ͷ�e���gwg���G�z�H"�$�ح��m����������x�m�����m��7��}�x��e�Ie$���~m��n�����ݿ�6��Sq<m��⓻������k���e�:WhWfmն��w����/:g�.������m�s9�ۗ]W$�� M�WP�>��fpFH��v�0&���h�\媙"659 �`HhH�P�eX� ;�\e�rdN3C�h�	�5������0	���v�̬1��}���|w 4@����r0.2����>P`��� �
��!#'�΃�nh�f�04��@9!M
]|nGgۆ��8�}��c��c`�0�mw�J���8>8^s�5�jw�!��w0�f�܏S��RV<p�ŋ�G3�$qs��*���.��[vڭ�@$� hI� ;m��A����(�椧�e5?��'��'��$9U��Y�
SH�R�����}�����`�U�8ҵN�[9��-���ԪӔU�oHH�[Mi0�mmW]���ڄ�:��1N;�2��y�1B��k�}{OF��� ɉ��ŉ�����̭J��@*ԇMO+UK��&A3�e�h�g�Y@�8�u��%��n��������I����Ҡ��hɷ�B=a�`c��gnK��������K�m���3#���H�ͧ	��cY�h�z �6�n^ �wfAȡ"���8;:Ȫ���z��+]j����t���\u�ݰ�q�z��v�N��e�h(��h�Ma�v[�ZZj�X��gnɬ�2ΌI�h t���:u͝@.ރfy�kn�^E5De̲K�uT�&�&6�Q�'mgs�:��4[;E�l���k��bYU�mN�!;�h#c�%�9�g��P�������/h�:��Y�aե�v�y�t�G[�8䈥e�#�%���LX�ha��mɑ���q�x�Iu:r8�\�Zځ��5d�Fũ���e�6�=�r\$�`�'�kE�\u��JO4��f�e�[H��� �受]��*1�m�T��T���c�c���-\��էM�����sw5�#l��h��n�<Fg]I��  =$�ΪW4�H�qu��*7B����)�e����c	U۵�R�j1rK��U�Q��f����Qe@K-�%�7i4�a�v���,H,���;6Q��9����9�'�i�5 !(�W"�H�,��31Շ��1*��z�q��+��J��+�0��U����v`�X�e\a�mv� m�]�SV�NW�55WF����@�t��
)nVwn;d��6f�۴dg���!�-m���[Nkԭ���R2fn��W�zĺ��C���WDGk��xG����Ԏ��ƀ����U]��C�0����	�*�� �T��
?"u@}���������u]����٦$沷:
��o�ݪ�IV�v�*�NFy%���kt�Ԏ�O��hS�.n���5�Fσí��z�0�sp)��J�-�k��7 �ƍ����v�c[�9�۶X�꭛C��u�HnmlV����+h�q�蜜���gG�T:�̛��kF�r!�{;��#����6����:we��eZ:�[��<<�w}w������Iex��ܩA�"!X�
ԅ�u���U(<c�ܜ�GI@�X]9ٷK�z��9\i�m�6ߺ��<m������m��u�m������m��v *GT��Q9S��m��.Iv_m��z���uM���m�e��T��ߛo�ˣ��ow�~~䓺��<m������������T���m��ݿ�6��Sq<m��{��������ޮ��Q�[�Dꮩe��6��Sq<m��{������������ߛm�V���k�$�z�ݛ=N�kѫ�4��3,Ln.�ntU�y��Kh��햩�� ~M��ߛo�ۭ�m��ݾ�����Om��Ǌz�-�K)#�������y��*)>* }��ﾶ��w;ݖ���3m�����˜�?M*q��j���+��m�{}~m����1�����ߛo�ˣ��t��9)-�;\��m����껌��{7�?~m��.�~\II=�z���}�=�#�XR�����{7v~���w3��m�������Ϻ�����o���֫!�@���t�v����}���pn�V�㭫�*��فک-��6�ݷ[��o��~m� ��9�����;ݶ��o닉u)�`����o{�s�>�\m����������y���mo�����]nU)��ns��l���ն��w���
�
��L(yUC�ֱ��ն�����v[�t�Ƌ r�H�.6����\�V�{���v��c?�ն��{��v�>P�;�f >���>r��J�a����?��m�Is���wo�6���x�m���? }�#I��l�yʳX�f܅����;�*r�z��ܜϙW�Ц�?{����[�	��B��G�������m�u].6�}���9Ͼ�����=�㲶�v�忿6����y�%�$m������������wo���IIv�C���)iT��m���_ߛo�ۭ�~I)#����m�꾯m�N��D���q��{���﷿���m��߳��m��{��o���b8KJ�����BI�`"�>�U�����￯��o�_��eS��%x���ʲ)�����;��LJ�ev\fXغq�#�tռ{Y[���m���n���7
�tɻId�����C�vMy\.�|���di�����K���lI��dE�9m�[L{��?�%��Fmo��=��,�g{	L�͒x�zWl�YI	-X�7� 7��$�ڶ��=��,{ҧ�e�ж�s�L=�W��l�_��a��s����㲶퍻d����0�sн��W@ͭ����`Tr(B��8�l�����-�) �.���T�v��Ys UW`d�0bć:��N8!��:w/Ol�^�ܺ�6����V��<�	�V�q�E�-��m�� �<��%�ql�s��8�y���&h<�	Ǆ�\u� |����;��#=�Ϝ� 9���Z8�6�ۉ�UBk�]��/$5����T��'��s۞��KU�Hӭ��jK�K�\�����J���vwF���uy�	��K�M�Tݲ1B���K�;6���s��ֹ�������͔�2IĻA�O4����"���9mX����%�s��}�["�i��#L�aUʦQk�Z*��L$��07di����`~}ݒ�Q*��WT���'����7�j��+�j�3����;��ЎPʮR�qX�ڰ<�/D(ͽ������,v��k�H|�MpT���q�ɻ�<>g����;�����u�q#���"��\\�yX�I��d��9]�~��f>Xb�kb%Hu��`kg���+���+�� �۷"Ii�%Ĺ�
"6!$��K�ܵ`f��`}��o�#������{˿?w���0�J�U�m��֬�v�Ԕ%=t�l��XuMP�9c�v�'*������� 맳`�|���B��[��7�J2Eb%j�`�;� ;�v�������ŀn�\h���%Q�P��EP�'/�fQ�4(���b�+e`T������w�&Q��G
�*VJ� ������������_�}�|�?o�c��Ex+�Wwv���~K�Tg��`f�z���ny.q��J{ԶA �RU�O��hԓc���: �$`�,�H�"��6�x �f{�gRN�Ǳ`��:��]�KeU�p<��8�l��,�j��D%�P��w� ���S���+���+�� ����6G[7��{��>�c��F�5K�����
Fbܦo���!Q�9]�䢹tFηM�s�>k-�*�����[6Հf7���9�$��7w�Z�P��%��V���`{�s���;��l��Vك�{#��L��+(;x� ��|������$��t�, ����7��ۏ�W��%x�)���`u�mX��,/��	G�S�@<�Y�u$�����\�9�W�]_9˴���`�-����`g{���.q$�G�5#db�G$�� o��n3=�	ݠI�c:]��8mՆ�R�[]���)]� �R��}��p�N��>�w�0�t�,��:����+����v��se?U'�`d��`�-��j�Ƕ9]�ЮJ���ŀ~�MŇ�>�z�vo��4���[kn��r�i��d���=��l�ow��j��R:�R����wq0=�s��6O4���`_X���`�����غ�<��$8-��Zs�+��l�5�p�F�M���;\����a�鬻�s l�j��aKQ�OC�`]�I�xu]>rKeۛ���&��wZJsۭ��v��u�p�5�α]�6ؒ��AY�o4\��(�Fz}dކsۊ��e���.�c[=�(H�-���ii�Zsi¤;M7o.qe��GT��N9j�Z[��I~��y��Z��BL\�v6��nݭ���8^��xڒ�Ds�Z�WB�ܖ �dV��9m_�{���`f�i���4����M���p�Z*��Lݍ0;�F���?};� ��u�,H�vIj�?n��vF��l�nƘ�I,��c��e-X����?};� ���X��I��{��;�۪?J퐶P���0;��Lݍ0;�F��`~��������e.Z�T-��zqo=�bKq{�'IڶU;��Ŕ�+\fL�xJF)���뜺�'�`wt�0;�4��s����GB�[q�9eX���Y�,E�H	�$E�� ��A�`@z�Δ)�
�	�
+f���d ȎMQL�XT��$�	$a��! �@ �c1a�$ ��c�HŁ �HHH���B�I		0g���������'�������Td\�縕�|%TR����`��ׇ�����`n�ŀ��a�U��ڤ���͔�����������'������1�UyP�W�}�w�2A����L�6Sg%r]r���3֮��a���a��E!��=�ٙ���Z�yq%�30���eu���~�g4�>�v��X��	/B���XI�{��DX܎W,�����X���;Vه~�Q�J*�ݙ�*һd-�!e� ��<ﻸ��r�< �A��H;R�BA��]��#��"ɐ�D!i��̻ �	 a� apHE�@��"�	�����i�@Π%r�X�!���da>��!�ZY`SA���"��g:�;IJ�a��PSj;c�a�!  �$�#
C��Jb�@�1 :P��!� @��p�&:C�	�@�ff�\ �����6`9��ŋ"Ā%O��4&L�`E	��T��}���ځC ����ځ�>V�|�/��)�t?:CB����� l]
L���Z�����s[�V�\SR�v�*-���{�'��,����?}�� ����iw�ж��v�Z`np`{��{��d��0;�`qs�����Ea��v6��g	n��Ԟ�f[�r�y^'τ���v��gg��u��ݾ��i��UU��1�Xec��㵱�[�, �|��"��n�%�`�;� �li���������x��:��D�r��`wڰ>�v��B�%U�}� 刺�ߦ�����t�Ձ�$�S6y�w�)��$��s6>���dE���r�j�?}�ŀ{�s��3g�`wv4�����{�w\�@32����\��[�[/=�GM*"���^��1�Df�րy&)tQ�5�[o������li��������V��/�wWj�݇+��`w64���i�����gu��K�����㰲ʰ��i�����͔��li��\���k�\���*���a/V=�U��[�>�n,�{t��7`�dV�ڤ���s`z=��]7y�����X �
`B>�C�L�l�����xn'��kq@콂z'�ѱ��t�����)<ݡ���]/%v1b�w�1�5Ι[����9�Z;Qm�d�|Y:9��
���l�XPζ��9�lp9;:C���1�8��:��=�m���ٲ�jG�`������nX�\�":��Ϭ�cyc/1Ӈ�;h+��e[kl�̥'wT	2=��1�ۮe�f�L����*ǈ!l��Y�s��?����+�~C����ae����!ndLy�`��[�/8��a۷�?l����T��tsΕ��]@?{�ѦwcL�Ƙ�l���Km����WI-X{�ŞI���`z{� ��wy&�K��Nȋ[�J�)�qXǶ��76~��B�(�Ǿŀ{��ŀoz�T�+�B�BZ��IL�Ƙ�a�f�u07b���v�[@�������=�-������ŀ~ٺ��}nNm*�ns�A��\a5�=�T��]���nv4m���p˰V�K��[J��,������?}ݵ`|�ԡ/�;�mXj���'��\��.1�c&����Ѭ8i*�~�X(� 	���sJ��~�o�����Lݍ0�"w�|%�ImX훯 ��w�9�q���,��`�F�	QX:���ulBJ"��ˀ6�Ձ�s���D(S����;�|Y]n��y]$�`�w�����S���������+�t�R �rC��n�j	n`z�q�b�b��\kqS�n������|}ٷBݬU�'���������%�I�`zkRzWlVZ�j�?l�x������p��Ş�I6}�UH�����B�Uɰ;�mXf>Yi
	� �֥��5�L(�P�}�?�Հ�f��㊞#����U��v���� ��u�{�{}�`j����U���n߻`{�z�������`ei_�n�m\$l�������-�\��2�&�6�p�[$��^HzT4�sL����76�� ���(��k�Z�7����qJ���^�{��ˍ������,��׀}�ݲY[���Wg9v���`nli��*��=�`g���;͛��kr&�Pv�.=����'�ǽu$�y���#�" BF
�o�n��7��͕��Pm�i���)����I=l͍0>�?&^���Q��F:�F�	�.�R�렜���\l���iݠB�����˾r�ƙ���+9ˮ���i�n��ƿv��Oy����#������ʰ����""=��׾�`g�ޛ���$�Y���?uY,(�l����,��)�ٱ����t��"����Wj���/�_*�_�L��Lݍ0����K�{}���;�����	��VNM���j��In�����Vt�ܐ �5Ah U��D`��>�Jv�ˌIs�\g79�`��m��c�!Tvk��[�z�P:K����Y�*�N[�Q\�8��@�:�-�*�2�\1�u��glN݊�SMi�.ڶ�8�[b�����;���V�<�.!s��9��s����������O����PYe���ޓ�uP��2�$Uh�V�x'�5+3liQ� ����Yf'YA��n����㳞����IU���f68����A�W�����jV�_o/[{���v�5��Y�΃�������Iq�Jܱ��Ij�=��ذ��ŀn�׀~��,�ٺ���"jT�����j�!B�DDDU�{�`g�֬��Y��s�6{�S��%v�[A�-L{��0;64��F��`L�jG6[,U[P�%x�9������=����;VIB�BJ�z���9��b-��Kl� ��ŀ}��,vn��wq`޻�ڧ+@�9m��]��=a�s��U7iSm��8ް��m<�<[����v5��,,�q�ʿ��b�7f��cv��G�P����j�ͩ��3����%�s�RM������)��6;q��Ƙ�~���UG����UX;i�}��,�����qs������ذ��V�+r�:��W8�<�%/��omX<v�5BI����}͛�숵�J��X������==��2{�0764��j�?!���m\s2n؍�������������,�Op�N������b��l+]�3��0;�4����7cL�V�se��U�
Y*�?wwy.6owذ���{��ˍ����%����-�+��x�Ձ��j�P��
�K�(�ZU*FA�T�V#HB�������Z5$�}��s�VA��8�dr��q>����>���nՇ�%�ߕ��R�䩞R�ª�U��`vli���{�]l�L�w���,�f�![",���*1��[n�7f��N\���9��t�f Hj'��?��H|]L�V����]�}��L͍03vb�7��,��1�]nX�U�Ij�qڿȅ�QT=�Z�<�֬��V���Nȋ[����Հ}��,~���脪�}�V��Հ��N)|+���\��W8�5(��ǿ+�vՀ���ɀ����$�B(E ����Q&��g��'��ɌY��Ȫ��[%X����?�8�����?����=�Z�qڰ:�]RI�
�ۉ#Qn7��^|�*:'#�Js��m�Y�nsFBђ�X�mm���*�7��,��Հ��֥	B�C�vՁ��*��R;*q��r���qg�9�ě=��,�vՀ����D(Jd�zrT�)rJ�v�m� �}|`���丸�����Xw}� ��{xHEU`���B��w����;�Շ��I)��x�7�钺�r�:������� ���d�0;6��߾�WBB��/ʔ)��P�BR�%ZZ��H�V�"e  6m@r
��ShB�2���'�ʻGiI";N?;w�8��)�κ�D�G�.��XB8¡�O�ۀe6 �"`��C�s�2�.9�%h�$BI��ק��o�"C;'�C�h`�A�jd���=�~��I����	 � ����ioVٶ۴��KPa扒��L��gi���m�-M�-�Q���s�YMNa�,��r�y�*�!X7�(Af�*�,�p[�1� I!���P�ܯ1��j�y�y6�ɊjNؽ�zI���f�M&3��λw\�����v���1�{:�by��X*�A�ET�SR^�]�;,�Vѐ�6X�mkdjxT6v���c�[$P]�np�R�6��tl���zԈ:���9s�s�=��X����3��-�km���q�-��y��3�cA�A/91��@�t��# �C\�t�7������[*���0:�4�9�/[�����tK�}trR��ʓr��#Ue�,=�a�ے$�w���S�UU+;F��ʠ�S�����6�:�v cْsMȁP���˚U�3��}�<�H:�z��Ѯ�m��.η����$ s\*k��dܲ��Yrv�6ٝ�1[HX2�b���C79���"nmE�T��-��	פ��l�6���+�ۖ��Vh�9<��+n�5"a�s�H�'(F�R�M���a��P�uQE.��/e��%����cV\�YL��I���m�!US��&%.��ru�(�qh���԰�v����nY��qu]��l�k�V��$Z����"� -����eQ�@�gA��*Щ�.|N9��	6��*2r5Y�n�;���t=2��v췣(!K�v�t �y�I]%�0�����Fܝa	ke`���OY4�C��jv���+���u��5���b`�8�����rL��XG&�gCr�D�m�U:C:�X�iܶ�2�1��+5��N�.Kb��� 6
D�P	��vGr�U]nmni�<��s�� ���)���̇6w]Gb3cx,�)V�54�٥`�a��흩	H���-��X*�$�y�Nlmq��+v-����x�c�oe�2�`�,��LKs�8:
����L�����M�Dz��6�'�
4*!
�EEj����%���F��u�$�-�%�� AQ�8�v��[8�e�Y�&Fr��\g�V�;d�Y��73��mĸz���o7eu9���y���p[Hu�-��<��Ym���[���m��歸L!�]HFր����Wv��Vl>�K ,�U��a��e1���c�ᦢXD��[v����	����R��4�^L͍Fdۧ��W�S����Bƛ�>�����_Or��ҕ2�x���n��jn����e)��HWN��n�~�{�ǫ��%�W$T�j���X��L�����G�(��{w֬{�g�|�\�.R�(&���d�0;6������Ɵ�|����:�d��Ȫ��Z�0�z�ݍ0764��.	�.}w�.�N;\�����x�7��X��Lq.'��<`���kը�G[q�0764��.͸0&������;�,t!S��܀nK����H���۶s�ԒtZ����D�K���ʿ}"Jܰ�ݪ��]�����ۃn�?}�	��`�7��B*�T�����>]Bq��(�$�zw���|XomX��uowq��"u[����L;�՛	L�o4�;��X �jyT�\p��r���{۾x��� ���`.q�wߖ��n����ح��r�d�0<�K=���<�s�)��=�O���)s]�R��/�P[s�8N�6�$LW���İj��g���u]��p�>y�X1ڰ3��}�y%�?_� ����-��kn;\�����3��l��<�/aL��r�����H�n9V���n���Ԑ��b��W#�9d���߾�3�L{�ŀ}�}�V;e����^�N�́�|��o8�K�=�^�ψ𐊪��e� ���`��`�w^�;� ׻�B��"���TT$�m���x�7.�]��-`;\���}�F�b��R'U�;)�n��w�`����0���=��nƊXB:��0�0&�e03v���.�I|��=�c�/),���nYL�7� ���,��U��x�7��M��'��J|��Wv����p`L���IL?}��G�j��
�I ����!$W�� m �����ԓ���L��m���-r��wݛ��7�Sd�0?%��D{�j�|9W�YZީ���I�y�kΒ�h��ΝGW��@1x���k+Q�T����|�����7y%06K�$�03lE�\�9�y\D�rl�no�!z*�����~��`ٺ����UV+%x7�Xmڳbe�ǹ�ń��S���D�;)�}�����x{7^�8�����o���[GSn�`l������.�4���ż\�s�+kI�rZ��D��r�L������:K��{{ThZ}�l
=����-�n�5���pᇴ��h�> ��e8�\�ӑ��t�=Gjٻ\{w �i	a�����N{m�c�%�c���n5���n�Z5�z�9��S����+A����d�w-�V��=h�/G\5;=\\qy�ݚ����-gNݸ�<�,Yfط:'Tt.�d�{�ߟ{�~������M��fpe��.s'l%����V{rZ΢kru/k<Y�����8:岵-��}���;�t�>��_��%��O��y�#'��Em�RK67�_�Jd�ݵ`=�ٰ3)��K��$���/�2�S���Y\���޵`c��Ϣ&s)��,�R��*�iIB&�b������̧�`cwL��ŀ}��Dc�F�N�!�^�Ḿ�%�oO��ݵ`c����ުӆ�@�7U�[$��H�y��S�m�m�[�a�W�^���/b��<�v������[v�t��B���D$�A�^�x���R�\��:���`�w~���R�脢"��uϦ�yX����ٯ��Uq���1����!��Y��ۜ�}^������`u�j�x���,�YP9\��s����\��<}�x�:۵`c������jJ|��*��T����L���~_��Oy�����zܜ�URq2�$u��ѸK��v��#�t�-�Ń��wS�G��O\�Z�6W)�n�q`ٺ���~K������d�j;*���r�v��!(��g^Հ�y���;W��8��R����Q�S��rՀ?���I9��R#������(�P�*��(\]Q}޾i`f7j�xk֣�)U�@���=����m�wwq`%�����>��v�VDգ�3�+��,(�{���{Vf<X��Q�(�nXۊ�8ۑ����;v�1a�B�ƥ�[�h�n�/M��}�	;u|(�Z��X�쑦���wc^��{����B�r��*	,�`}�W�P�F�ڰ;��,�v��2wt�q�ֹV�+� ��b�?n�0ۻ� ��v`j�^�Uk���XK�a�������ݵ`d�:��cD�Vڒ�N�F��X��5$���mǵ��	m9i�~��X�9��ż��t�������d�B����ti v�L�:�L�c���W��X��7[6�>z��tu�e�;h�-X_{� ��j���3c����iSe*�j�p.�͍0;%���#L}������O��r�VDՅ�J��~��2F�[���`I�͖s��dM�L>����{���n���\�{�� �|�P����J�ImVNc�TyC{��<Xu�V�'Q"���KU�D�%�}%?q���xv��p/F�l�Y(�%8WS�\��E�6�d
{)�%���-��yE�hp�qvR�8M�n#������g���Incv�Օ�t6jɅ����8�]X�q���uv)�Pٴ;��Wu�Ms�{`m`��<�*��v;�jl�/�v����p�W�ݜ<f۲�5�O�+<��-:�;R�Fz횫v�1��c`��e�DM��h��ߣ}�/�g���l�ۜ�c<��֎�Գ�
�`��w[�,����K�5�T��]�쑦d�0;�5���J���>��g�*��h�HKV�v��Q
d�nڰ��`w�~�2k�T���tv�G[NZ`�{����>��,��� �Ӻ���F�N�"�V��8�͑�M�0�U���`lR����� [f�wq`ow�wq`n� ���Y �+�J� ;�1`!�5���c=[�����ջ=���ՃA�`���1d�!)edMXXݫ�7��ذ��� ��v`ww�����Q��f�5$���t:�P�� ���]P�TCeO~u`<ݵ`u��2{��S^N�]%A$��_}�}�v��P�s^ڰ1�ڰ>m�SJ�\���ݪ����6F�64�͑����➻��0�V&J���+%�`x�X��F=ߗ�9�ڰ;�ڰ;��ꭡ;d[l�� Jꀫ������Q\iv��g�t��-�����~ '��s�uEW-t��L������h7��X�=�Fd�v�m�`n��"S#{��׶���XŒ'"�UX�l�;��X��Ň��O($�E L�Q�Gq �F��Q��A�@�W"� Be�2�A]���L��5� Έ��(@4�v���O�� %m���0CW��	�	3��t(�FO��@ �v���5�@���@�>�;�_ ��n+��ga�L�:2`�N��f�a�P�0L
�v��")#)�
A9TE�p ��1v.��EI�
+��q�x��D2��( @γ��F���w�ԇS�v5)edMXR;V����9��V��j���u`f7j�n�8�V(�uW%Xۻ� ���K��=_�]w޵`u�`by'
�L���R���u=�b6�.�&;m��yBF�5��۔�^�EU5S�V���Հu��0��V^;Z�P����VwuZ�U��WWv������0;64��#L���<�8��>��<�*���+�Z`g��`d���l�vF�%�ڏk��0+�`{��8���� ��}�I9��F�� �@�	H �H  a�
|���]�c�5$�ӽ1m�3-ŗ˾R���`v�g�4��li���� ��xfH�z@�*�B�T���M۷j����(���lvne-\͐JZ���?����O&Y"�UX�,������ ��w����??�� �nƥ,*��
Gj�>�;W��!)�7vՁ�ǵ`f7j�I6{�Oޕ�
�0�V�0�����f�3��/�T��L�~��j��l�YP9-���N���b�>�q���(�~�����4��ɚ8�v������0?/�͏�@�{�07~�q�&ǭ>���$;iq&�)qV�f�9�jWvml�p��"�q�r�8ۑc���Z���^�4��n�8U^4�*�n8����<`�t,R�M�����ͰM�]�\�`��c�::�:eڱt༽�I}M�=kjy�؅�n��3�d�h��A�yEև/f2��n�qҖq�t�kl��^�#��:��'���Ƈ��D���Y�uʝ���jK�s9�˟�*��A7+��e#��m�N/>wJꗋ+�cE����,�̛��w��\�X�*�K+�+�U�7�|`n�,���?����,�������� W,`d��k6q��#L��3�q.s�q%�!��򍼔nR�D[�+%���n՞�3�|���ݵ`w�w�"�UX�,��K�s�w����~$i��͜`j������Z�|,�]�sn%��%����V�L��ŀ~v!���7k��!�Xz�t񱱺��rF[2z.&�ń�Z�gqR�!Y�ݦ����??�� �wq.s��}ݾ0�����V���s�RM߹�k	�@�A��
�a
� �_�S�*99���P;�|`n�,��N)md*����X�ڰ>�q�jP�D�n���� ��U��U�W]a\���q$���,��V��ua�P�)ow�`o}cmG�����`n�,���sg��$��`w6��ȴ��˺UJ���,6�!��A����sqvs�3�s���;P�3%X�ꍻ(ܥ��[j�??�� �nՁ�s��B�_Hf�ڰ'QsK�V�U�"�v�ݑ�sn�4�?}ݹ�..6j﯇
�*��
Gj�'��}5$���L��##�Q����v���� �Q��,hVA�����Q�����,��Xz�<�{�̼k����r[V ~�v�$i����0;�(�A�r��5�Q5���w���A���ݮ"b��3nLM�L<j�����b���B�jl����{�`fm���#L�I�d�"�U�,����m��v��fｋ ��ޘ�wf%��o�m��%�8 Mp�ݵ`}=n��9;�Vc���ꍼ��j�֋mX����'{��RO��{5'W�&؈�QX��
-DbU�ҫT�A�GO�� ?�}u`����"��r�`�v�Q1ޟ��Հ}��`zֺ�)�C�<OS����a��^ڌ�ɝ�ָ��re���:Z�)m��aTMXV;o�;ݾ0�ڰ>��Z�=���r����}')��%U�Lw�� ��ݘ�ݶ{�e��yDs��Tʉ��5T�����sy`nf���64��Ț�)md*���v� ����t�7{��=�?�}�}�U�#��+�����f�li���8�$�l
��	 $A,T
A��N[�v[��fg8�m���
��-�މ;:plt�z/#sS\/5q�8��MS�F!}�]�|4!֬����e��s�Ӛ�U�JS��L
[���#���/%m�WA�WS�/q��C\U�����*��v�{[�Kq<�jeZA�|!>�ny�F7\.d��	�j�Lf��e�b[<��n�N�	��������ma���{��_����7S�Y�z�펥���x��a��e�h�;q�:��8e�u���?$mG1�[#������ ?}�pw�p��� ���H1�r��[m�k$� �e�36���cO����{�����"-� ?���p����߽�ŀw޸~6�u�a`5ad�s��T������֬�� o6�����)!��`��Xܒ��-���t��ʺ,�1;>n�:������^mXm�j���46��9̶�D/s���X�q�*%�~ ����	6[3n	64�ɱ5\\���V��nـn�qgRIb�R�X�N߆�y�k$����U��]�WAwʻL͸0$��?}U�������j9��� ��\�Q^�����~�X�`w��Xw	�1�r��R�V��ݘ�K�%���W@Ǽ�`7�Ձ�P�V4]Tj�7m�YBƹx�<g�C���[A��Xs��牎��Rn�8c�J�,��?���� �m��&Ƙ����J�|���|)]ݦsn��=��l��7{���M�����Tv��wF��s�Ԣ��b8�
��)�h�B�S,�8���IB�$������K�&�ɩVTKj��\�o���o�`w�Lw�� �{��$��J����n �;V��	���{��VӍՀ����?�zݳ�gү$;��A�=��E��g�ۭ�/M�t�f�Ş�K���|����ۃM�0;['=�]�����=�X�D�����	�Lw�� �q���j��g~�������$����KmX��� �������}ݾ0{}� ߵ�׎)(�DYn �;Vs8��v�9�! �A�4E.����"� G��IU�s�}����;���배j��ݦn�li�nIl	64�0�~y�~N��R��Ҷ���4�{ggu�ugiz!��F�M��{M"�S��\��li�nIl	65�Iv�}/��W����;L�[V w�ۀ7�Ձלe��;W�%27�3j���R�bYn�o�`on��w w�ۀ~�*���mn��;V�(S��Ku� η�B����X�X�G<�-��r��w w���o��8�T��BJ8�A�ʮwKM��v`�a%!&���C	�}w�ٜh�[�j�.0b`��s`���x�#�V)<ʉ�'C p��b��*�����@֘�f���2a�d���.Q���d��T1���B/����@�H	 ��cP�C�E9.5�#��;�/̈�|*a ���N�]�~Wt!S���qC������HoÃx��� >I��x�QV��9N*n�{�{���{�+��&�[ 8� u�� %�H[Ԭ��٩��l�a�lM����6���!�X	���K�\++u$�h�����M�s�a֛+��E4��'[��5%���m�&�\�`��0L��s0t  �ۋ�牶�c�S1ӡ���UЅ:1�Pr7V��C7]@i�쀹�s�6Ͱ������Q�X�d��cW0�2!�������κ�b�r:�"tn��"��bQ�Lb��,�E����p۵�Y�c������pmM�%!��g((�ͼ�ɠ��8���9���w*d݈�ǙH\�b��g&5����(�-�01�5lb`�%�[<�kr؞nݤ�FLf9�Q���e���:������D3��.6��؝k`��/W Ct����8�B��;'\J�m�dꁷ*�$p����3���0� ��ڊ3�K�nS%�7Vky����V��*>�%�����C�I�6�C�8��y�4JuvO2u�t۬�$7(�a�����! �h�E�흮�;�q�U������u�b�Y.�������+\Q@.ɔ$'nt�eMk;�]�'k6�8$z�e�2�+��i�*��8XeQ�ۛUڮ�1���AU��m��+��m�t��qF������r�Snw-W=��1)�j�[R�lU]l�r]d�&�\ vSS*� L�mݘ�峎Ix��+tEqҐeq����s=1��p��G����kv�m��n�oE�N�����b;v6�5��GTkg[K	��{'gti�a�&۬<��8ٝ�����:Sl�c#�퐫u���fV�AgCy�f8�zIUM����%����qoIn�Vp�܌��UjU55Tl��.�q�=2T�Ƨ���x��;m�*��gA����b��:���\������^�aъi|�m�y�v��"S#Gj�����@3���n݋q��0�P*���Q5F��+JI����e� D
"l*���u�`P4�] < ��(".H 9"�C�@BT{�q���u��m���z2��uc�����<ni����]!��JP�\��K��M9ynY�Ŷ��tWnE�q	���j�WT$ǃ����̓���q�r��f��-�z9��j�'�h�iݨ�0k�S�Y5�NJ^sjbݫG=m��κ��9���z��]��q�Ŝ�e���Uk�e�jg��Xj8J�
㎖S�S�s�9�.*K���zGgUͱќXK:��!gR�٫��h����,�]�ΐ�,�YY-΂p �1��o��8�D(K��{�ذ��m��)(�E\� ����:��j�3���D%#�<��T�aTj��ڰ�o�w�� ;���7{���&�FհduXݦ���XǼ��j�ДOuޖ`�����c��[V w���?������|��o�b":�K��
�ʨ�48�.�k9�Lk���kkh'!\l���Z�[n���Z�@�UT�X���?�����ٷ���ݠ&�[=�וr�R[I#,�Հ~��3��s��~K�w���`ݖ��cO�Q'��Q��ˢ*�cޞi�nl��`~��0�wci�����j���l	64��ۃW�=�����:����\�s�x�X��׵��q`~��˟x�g�����-�c:�v�|cm�]s�_췐���ݍ���=��=�HWq�X>WX[W�u�{�`��X߻� ����;���l��l*�I|`I�����li�ڛ8��F輝���c��[V ow� �����l��f�H�$��B��r�
����0��VUc�U\3�\o�ԓ��tjIÛ��	%UJ��N�p?�.s����ߖ�׵`7�Ն��z�^��{��Յ%��2��X�ـn�q`~��w�� ���e!�l��Ȥw�u�C��'�B�ͶWm�2���:�8��[���L����9$���� w���7{���0��}0龃EX�C�V�U�gq��B��u���j�o���������"�ۀ{��X�ه���ذ{��w��ۏaQe�����f�0$�� �l��M}����K�\��~X���-�6�Q�Z��]�&Ƙse�$����9�~]�.�Ex�i�Q
��r�2W�\�d����OqCPv����n^�/d��7\^��$�s����;�-�&Ƙ���ݠ���`}�/<MI*�U)N�p��0��u`7�Հ}�|�(Q	/%Tg�qyL����FY�׾���w�I���� ��ذ��8���VF�9�X�`u�X�a�"!/En��<|{�6�±ʇh��� ��� �$��>�{6x�X|�LB68����F��ڼO6�'�)��GFQt8zVu�����zU�V�F{D؇8ݻ]v�\�V�l���"5WU�G��S�ܵ�tWi�.��qŬ�N9�㮨�g��"���p���M���s�v�p�[*�j�0�����p��v�Ӓ7\ca��kMū�w\��PkK��|��;���^&�m�r���R.��UH� R0!(�..o&*��̓��3l6��9z�� Z�?fW\�5 �"�,�'I^�3����kb[mp�Ms���Vec��v�"�sv����r?2�
���`l�w�� ��v`��g��M��{��cj�Aʭ�W�{��X_۳�����,���}�]�4-q�J�%�`n�&Ƙ9��li���)�\�-Z�Y�AW|`I��T���`u��0�ė>��x����ٻѬk��nwJ��^RƊ�9�S���|�M�9ꜰ���FY��~�Lw�� ��vs�{}� �f��c�+nF譸�5$�y�hCLH@v��TG���]鵓�`wv4�ʒq��lG*�c��[mX_wf��Ň�����������XV�5�RP*r2�0	64�ʒq��#L���	���r=eՕ��`=ݘ����/�k�z`ow���P�7����2���������{tj�m��v��Re�>-\n3[,��j �V�l�;��,��� �{�����嫷���H핑�x��n�aDɚ�Ձ���`g[�`}ޭx��UT�R&ـ}��X�w��ѡ񩤠Ā�~*(�E��,D�*s���ذ}����j�%�%��2¹�a����`fnڰ2{����X{:���6�v��q`wf�۸��{� ޭD�)d���sh�qǖ�h�֬]��F<�垛c�v������+&(�y
��v�Kj��w��̑��%�3$i�BQN��j#�X���}��?/s�\�;����ŀ��˜K���uѷ&���ee��`���3$i�f�l�`o�}�6ڕʤRKp=��s�M���N����I���I�E#*�8��(�]�Z��&Μ��l��-��.�U��`�[2F�l��̑��z�E��[�dU[]��HJNA;��ۇ��7�1\�^�LKT<f{o�{���|>q�*��R�������`�ݸ�n����p�-�T���$e��`l��̑��%�3$i�䒪=�Gl~%m��$� �}� >���>�w }�ۀw����:�`ݢ��V�l��̑��%��K�����ywǑ�+jq:��[n�۸�6K`fH�`�[ _}�۠UT9;%��ut6u�v.Tbn������단^�J�칔э$�c�v�bCl���O=q�ۚ�q�W��\���7Ub��%������S����Ȧ�D[����qD8��1�x����kZ	0�c�֗��G��nEm�d� ��r��A�����W�����w8oi�1��o2�MUs��m��1�t�r�\�6[�ni�d�(r��@
)�������gK@�n`�l�2�	ƴ���on5���>d��uu�,�u�����=�`fH�`�_�|��|�p&�b�<�y�R6Ԩ��:I-�>�u4�2Il�`�[���"�Scl��v�V w���>�w_ː���{�~�`cl�T�k��qW*\�]�3$i�n�l�L$����ڵIaI-rFXKV w�� ���(M�˫�}�X�v�Ƈt���!����hguz'����6�2��n�kW�:Muƈ�M�0
�-|�}�Ț`�[2F�l���"����v��E%�� ���7��� ����4�
}�����I&��X�j��$�&MY���9�)U|\��`n��0�-�J�w�M0���?j;X�z
�Օ�ڰ?��o��[w�M0�-��#LÛ�g*��k�r�,�9v�̑4�3d�d�`�ݸ�I}z9�qG`8F���<n�V��[
ĳ'gL���^:N�F�%g=���*�ʰl-����U_ o����#L6K`fH�`l����\�tZ喩s��`fH� ͒��&�n��qq6{�����,�@��� �}��I���S%] �&t�18�p�e%!J*��`�)�!Xu�u��	5�SF��H�Bf��BXᑦ1�]E�H8��R����� 0L���g�
�c;�&�P>a�aMoa(@�(	�bP2�?$ �6m��q�7WN3�HE	�A4B��e�D�M�� 5ɿ�&RS�i6�P�x��r|��>I�G�6�����~@)3Jiq�iIPe4�S*)O� uM�Q꫑D��+B;�]�T�"�p��N�%�W����s=Τ���Ѡ7��H��+nF�%��n�X��,��V��{��5N�꧊�誻9v�0�[2F����[V�D(�X�uQ��
�&�9À����n�g�79ؠ۝�M�s���Gl��wYF8���T�Im����, �wn�q�^I~(����,�7�L��%s�WUv�we��U�ɦ�z��1`|N�6�*��J[m�>���`we����7��d�����UuN�-�ݵU���ĸ��w� ���0$�9��J&�$}+|N��]�{'� ����E��㮦����ۦ�/%Y��t��Ձ��:�;ړ�u&ݱ�<B�#�Ѹ��ډrݻVV޸pr�ս]h�0�N�z�C2�\M�`;�[3bi���8��K�g6����+nF�v�ﻫ$��?����r���x��/�&�d�uU\S��������\��t�ˍ�n����b�:�n��+k U-R[p?��f��`���36&�f�`v#n�nkU�+��`�n��$�����'9�gRM���jI����0���`S� \"8L��J�4�Tic�S�Y�LLvf[qQn7By�n�V`���7OZS�J:�;�*�ڿ��|�7�0LQ���h:c�/^H�k�n����^,n�{)��ͮt��OkWW��Gc�tԎ�>�c��m�q���ٳ�kNf�Js��7r^&����J-���p �q<v�k�Y�Ovn+���㸺�`�mp��tI)��M�F2������5��ǽ��~b����8dT�*aP�Z�8۵�)K��ʑ�%�2��#�m̒ɬl�T$�R�n��{V, ����?}�O����� �#j��m�"��U�����p`�-���4��(�V�%u5� ���0�۷7��, �w� ߺ���`�6Ê��0�|�������<�`�-��ۦ��d���n�[m�>���0͖��K� �Il��9�Eߞ�l��pMrW)��v�)������g]�sa��W�V��nZ�m����[�.�%�$�_}�������8���d�Im�?}�L�q/�q%Ԕ��6�s��&�f�`v#n�d�*�VW[��??�f��Ջs�l�w� ���0�ӯU#n"�uK��Q�o|����,�����u`wQڵ�cv���j� >��p�K���q���4��h�K.��P�⋈�s�<��7>D�#�6����Rz�r��2��E��䮦���������,���D} f=偸�T�`�6�'e0��ٞ��I6w���3������P��Q�j�D��L����p�,X��ۇW?�s���P$!$)K!wT$�w��� ���������)-U`�wn��� �Il����):⻺8]�\�ݰ;�`~_Vo�}6y4�>���?��%��Oz)!�6���I�ϲ>�q����_췲|k����Y��9�lz��\j�Յ��|����ﻫ }�ۀ~��� ��:�R6�/T�����V�пP���`c�Z�2z�_�I�|�U�ݍ�+edr�V�m�w64���8��lM07vU5��嫾I,��%0<���~X��� ������������z�`ܼ��RN|r���`�6�9j�:�ݘ�]0��Lﻸ�٣�R,MG]w+�]m�=9ɵ��3l�m�p�)���9L3�Ė ��+nF譶��wV,��сٱ��I��)��Z��*��wv�02li�ٱ��I�����պ�8�+!\v�-X����:��Y�
""e��j��{j��K�Js�V���]�v�Y'�L�a�$����� ����#n"�uK�X�jՁ��5���;�mX=n�NB�R�-���Əb[�f�uĝ&��Dm�h�Ik��mX�C�8�b��J�58q����X݂������g���6{q�v�@s7�CPu�YP�$0�������\rڵ��&��r`��F���֑�/.�Y�ګjl�,�;!��ַv�uȭ)T���AɎz�������5�|�	b���m��̨
�ڎ�T;�:�1�����P��X���ʗ=��F�'����ܯC���]�*9l��е ��x�d�u�/+���[+%���������j���u�P���j�VofmR�Um�YS�ڰ����5�ݘ�n,~���7���N�cl#��Vl��i�3cL�038N(�zJۑ�+m� ��[� ߻���ۦ o�ۀ~�ձc����)"�L	�`we��L�l�#L�w��ݿ"=���1��bm��#�����v��{^"#�G7Mv�,m�<qq6��J�����~͖��R4����~Q�6��M��RJ`�ݹ��8������H�I`dۃ���2�x�m�T�I%��{ذ��� �{t���p�V�m ���F���3cL�p`6[|�ʦ�{�������y[c�*�vՀ}��`���u7j�y�Ձ�"kR�M!UV�Q�S�0��\����c<Kؗ%�ƺ��R5���$�t�lM�������`n)`M��]���,�������#tV�f�w�P;�צ������?|jj�N��F�� �9��I>�3٩�j2�B�!
Ti�z���w�w�Ѩ�����)Y
啹)�}��`��X�ݫI)��K�D���J�T�r�9��-������~on�Ͻ�8��kH�$�Q8�-����`����:�:kw7[d���r�{h�v�m9��j��9v��R4���M�0��p�t��[��VHյ`�p`dۃ ����F���\U&�luҩ��>��0~���-�X��L�W]Z�,em���	�[7Ti�7n<�O�$� d�SÑ�}�njI��=������Www�n��n��p`J�&�����c��t��
렧&��^�ѭX�)��G�r\����Bټ=uá��O8)�\�g`}������Q���/�XW����qJT�Y[��v\�N03uF�v��ȶ�UNk�TڪU$� o۷ ��[� ���~��0����q��$� ��`Mۃ�.d������2�Y+#�Z��n���� ���Τ�s�tjI�	��Y@��,@��H*��
�L�mQ���3 ��B-�|$^T��xŲ��$�ҁ�"9�DK"y���S8y�]��>z���<��XE�7�ji��E'�&,����K*����H2�d$�&0!� �H�H/@����1O����0(@#H�8IH��1�#$Ō�l��"FB*�)
8T6��w<1�c�hp����m�@��*���U�9}����-��ڙ�T�Fe.�}�n�Tb�d�E@�acb^ح�bl�a��Nl�:�d&���(M�L��+&	� ��� 	l�U�F�^�KK5���n�0�u�!�t�UƎ�W0�c�vZB��z�X�p�,�L���K��K�Xͪi7\ ljں��ȠF�vz;BUF���(��Ckvo*�y{U� .	��ʑ�+�GZu����$�f8�v]Vu�ڱ�&tu�5�����m���v�֜&sRkPPh�;�(ڀS��۳��=��\��f��q����>هl�l�� Qr۝Q�۰�Gp�{1/���^�x�(��f���b�ӹ۳�ˡi�M��c���Z��I�P�Zr�cn�X�n���[j�gr*��+�scU.@Lʚ�L���b�e�m��v�C���m˘���yM�]9awg����=��w��G�1�Kx r�s���>er"�H�.�8X�����E1��`Ԟ�P��.
�=�ŵ��j�9.���P�M���n&���z���v1c��G��%���Pt���mz�'G8; @�M�2�v�R�uV��9�����v�tAu�T ˲�T�݌<Je6�wQ�j�c;�Q��0����ٵk�����ֶ�:�)���������6��P%Z9�Riz��z 
��x�ʑ2���#�ϊo�C���1�%�U�m���\�U=,�͝u�&�UX�5�A�L�U�v�8��r� ��*��K�kU�=�r[*Ϋ�}��Wh|9�6�z��n����;v�C��9ą��,m�&ƫF'�I��<FjIT����̐�U��6�s�%kP!�Y�����R��Z��+x�ji�!�\��	$4W��!�Z��:$-�.���:��}%�kN�8�$u��;\���
tUK��--D��&yUek*m[���k+�d�M�9�r�kJ�ā$v��7* Q7u����e%�� |.
�U��t#UD��D8D
 |���<�"��ʁ�R�\X��p��ht���l,I��ϗj@]ڴg�&ٳ9��庋��cR�ѮN.�xt.�Z�v�۝x�\�lk�3��G&��C���ti�Z8���;"�A�{rn�']�N��:�G;�o*R���F�f3�M���;+��r%6Q���<���묀݇Qͩ��c��'�9/�A�f:�a��nSu�²0;�µts���$x�7Y���c���������7ϟ@nzЎ�u�f�w4m�PN1�vxl���d"b�ļ���<fv���ulu��W)�?{�L ߷n�z���� ޮ��8X2��`;)��[7Ti�7n�?�$�J����F��X����p�b�7��Y�	%3׼��77y`w��e��<�
�es��0&���ݗ2K`}ޭŀ~[��R���X7i�~��0<��l���y�͸0&r����nq6�蹂��l�<�2�m�'�9����]��@N�:��m�m�}��7Ti�3n�p`w9RÔ�U4:���`�V�Ƹ���5�&�?)�
 �~�gϦ���٠5��3�..&Ϲ�*�vB�Y+#�]����p`J�8���`d�uD��m��XB�`�n���� �z��~���m����vV��9cVI���n���w��mu���U�T���9U�	��
�MH!P�q�kV�uԽ���źx��)m� �z����?�q3��_{���~B},K�����n%��&q{Q���8:������)�_�&%�b{�צ�p��D�K����I��%�b_����7ı,Np��i7�b�"X�?~����L�ى���[��Mı,K����I��%�b_s�Γq,r��zE!_A*���I�i�򮏢}y?}�I��%�b~�l�n%�bX��۫.1�Zd�2c%�34��bX�%�;��7ı,Np��i7ı,Os�٤�Kı9�k�I��%�b}��{7�).L��1��7ı,Np��i7ı,?w߾4�D�,K����I��%�b_s�Γq,K��'�`�1���XTX�G;�U����hN�Q�6����o%�q+)�=���]���U�Mı,K��i7ı,Ns���n%�bX��ﳤ�Kı9����/�8���.�S����t���4��bX�'9�zi7ʨG1Ŀ����n%�bX�����&�X�%��w�4��bX�'�;�O��K3��l�8�f�q,Kľ�}�&�X�%����&�X�%��w�4��bX�'9�zi7ı,Ns3�K�ܘ�-�1��9�n%�g�  b'z~���Kı?w߶i7ı,Ns���n%�`g��B��z��N}�z�㉜L�g���E*���F�ri7ı,Os�٤�Kı9�k�I��%�b_s�Γq,K��{f�q,K�����ݹ����ŸɺWf���۲�����l���� ��皎8���$Er�B�`ܫ8�L�g8��g��q,Kľ�}�&�X�%����&�X�%����4��bX�'xk�9=UF��9)�_�&q3��O�����?(1�LD�;���Mı,K���f�q,K��=�M&�X�)�_-��u��U4:�RKs����&%����&�X�%����4��c�TB�����~�Mı,K����ҿL�g8������b�P��j�n%�bX��}�I��%�bs�צ�q,Kľ罝&�X�%����q~8���&qwڞ(��V�륄���n%�bX����Kı/��gI��%�bs���I��%�b{���_�&q3��M~_hݞ�JK)���N֨������-X���m���Z�x�$��v�-3���1�k��
�.��ȡ��ۍ<=��M\�n����g u�[6�4�k�v3�\�ճ'mGX^�x�ٍ�v�7��aN����HL��Ǫx��K��&�	�^�\����ڎ�v�|n.�\��a���-՗����R����,0!���a������tw���㻎����,J���<H���F�#1ǵpu&�Y[z���F%�VS0��YI
�L���J}�Ӊ�L�g���gI��%�bs�}�I��%�b{���&�X�%��=�M&�X�%����h~�K���s����&q3�8w�4���"b%�����I��%�bs���i7ı,K�{��n%�b�ŽZ�~q:������j�/�8�K��i7ı,O��zi7ı,K�w��n%�bX���l�n%��&q|����䣰er��Vq~8��bX�s���n%�bX��ﳤ�Kı9þ٤�K���!1�}��8�L�g8��7��F�Q��NJi7ı,K�w��n%�bX�rw�4��bX�'��l�n%�bX�s��_�&q3��OOj����#nX�p��RSb-W�@�{\=nu�7la�7��g=�˫k�6⩢��$�8�L�g8���l�n%�bX��}�I��%�b}�k�I��%�b_w�Γq,K���7����B����q3��L��}�M¯���Lı3�ksI��%�b_w�Γq,K����٤�Fq3��[�(��V�륄-�8�,K��=�M&�X�%�}�{:Mı��1���l�n%�bX�����+���&q3�wqz�Q��6��Sq,Kľ｝&�X�%��'��I��%�b{���&�X�%��{^����g8�����1�YJ���K%Γq,K����٤�Kı=�{f�q,K��=�M&�X�%�}�z�㉜L�g���K�&��	��!�fK/^K��Pr��8m�']��h]\�mͺUq"�+`�j�/�8���/w�٤�Kı9�k�I��%�b_w�Γq,K����٤�Kı8{޴��6d�7&1�I��%�bs�צ�q,Kľ｝&�X�%��'��I��%�b{���&�X�%�[��D�ѵTj�S�����g8�������Kı>���i7��H��@�:�������٤�Kı;�k�I��%�b}ɟ{77�)2c8-�s��Kı>���i7ı,Ow�٤�Kı9�k�I��%��f"c��~Γq,K���Oh?�p�U���g㉜L�g������bX�'9�z�7ı,K����n%�bX�r{�4��bX�'��>~ݮYy؍��,W���9��]���g��7;�M�r�,۶pK���-9��M&�X�%��g޺Mı,K���t��bX�'ܞ���'�1ı?{��Mı,K�ϧ☗%��n,�&n3t��bX�%�}��7�q,Nv~��I��%�b~���4��bX�'1�{Mı,K���Ŷ�9�Ɍ����3�&�X�%���{f�q,K��}�Mı,K�Ͻt��bX�%�}��7ı,O�v���2g�K��bg94��bX�'��l�n%�bX��}��Kı/��gI��%��4}�Z�Q
��D尿�I��%�bp�i7n&l�fn2Lc&�q,K���]&�X�%�}�{:Mı,K����&�X�%����4��bX�'�����3��d�k@њ�;s��ki%_��E�Gc���3�Vs��zػ)!�'\ܔ}����ou�b_����:Mı,K����&�X�%����4��bX�'=�z�7�3��_.�z:�n*�*�&����bX�';=�Mı,K���i7ı,N{>��n%�bX������O�|P�g������p�U���gㅉbX�����&�X�%��g޺Mı,K���t��bX�';=�M�&q3��]�7�&畲X�ij�/�,K���]&�X�%�}�{:Mı,K����&�X��	�����Ɠq,K�����q���7�$��Mı,K���t��bX�';=�Mı,K���i7ı,N{>��n%�bX��,?E�����8D�yڌ%ʗm�9x��瓈�t��u�W]�Ye�M-��zL3r���:Z˂3����"�ʹ�v�v���+T��7O�;���D���vY{.q`�MC��F8��Yg�-#���t;uB�ru�/qA���@OGN�����9���y��zŲ^�}8�Lz��ݷ"@
�\�&3�a�#6Sd�L1��p� m?~�w����{���~��=��r\UU��=[���瞎2M��*nݹa9�av�<M��%�a�n���9�z%�bX����٤�Kı=�{zMı,K�g޺Mı,K����/�8���/����
� ;DI���n%�bX�ｽ&�X�%����]&�X�%�}�{:Mı,K����&�X�%��O{��6d�7&1�&�X�%����]&�X�%�}�{:Mı,K����&�X�%�����n%�bX��ۢ�_b�&)�1s���K����L~����n%�bX����Mı,K�����Kı>�}��Kı>�Ͻ���n�͘�s��7ı,Nvw�4��bX�'��oI��%�b}���I��%�H[Ov��)!I
HD$��N�.�ZЫ���sew��#�p	m�ܽV:��%x�+�)Pr²�±Wj!	j���q{��SPI�q��	"y��5�,K����&�X�%���]R�x�K-!m�/�8���/�}�_���V*1R,� H��W���'���Mı,K����&�X�%����4��bX�'y���:�rr���q3��L�~�z��,K��g}�I��%�b{���&�X�%��=�cI��%�bs����?[
���K%����g8���7ߖp�Kı=�{f�q,K������Kı/��gI��%�bw�/���j;D'mY���g8�����-&�X�%��s�Ɠq,Kľ｝&�X�%�Þ��&�X�%����q�~�'ݛ����V�ns�����#��@׊I���O@j�M�&���\hn˓i�Kı;����&�X�%�}�{:Mı,K�=�Mı,K���i7ı,Ox��./�s�b�1�9�f�q,Kľ｝&�X�%�Ӟ��&�X�%����4��bX�'=��8�L�g8�]��u��U4U,V�9�n%�bX�9�zi7ı,Ow�٤�K����,�E�sE���(d�Ѡ��	�I@b���`C���če�z�	̥����iMT��J���GI�s��"�=���&�P��z4�4������ٳ	ܟw�!�	���U}
��y�a�I�X��	>B`��eR*Gﲵ��`�)���$$$b`2i3��N��*��P�Bs�b�,�&�hFl��]�|h���Ё.0�a�.�7�.���s/?�lHA�	`  �ك�Δ ���P9ӘHƙ����f�Dj��p�`����x�9@2�G�^���M*`'RiQB�`�x��"�q�t�*��09
|��D�L{���n%�bX�c��4��bX�'_zh�������I�\�3I��%��@������Ɠq,K���k��n%�bX������K��"LD����4��bX�'O~�M9?��V�ij�/�8���.�s�I��%�b_w�Γq,K���k�I��%�b{���&�X�%��翼[�O���[n
g�Ӎs��a�����Sg��V$��u�3�$���(L��1���Kı/��gI��%�bt���Kı=�{f�� 3蘉bX���~�Mı,K���ql���L��%�1�c9�n%�bX�9�zi7ı,Ow�٤�Kı9���I��%�b_w�Γq?8���'{��ě�&2f���!s��&�X�%��߿l�n%�bX��u��Kı/��gI��%�bt���Kı/==�Rj*�\�v՜_�&q3��]����Kı/��gI��%�bt���K���@�#���#�$Q�BEG�E�H!1��A���"k����Kı>�?h��-3�d�L��Mı,K���t��bX�'N{^�Mı,K���i7ı,N{���n%�bX�����`�M�o�G��ӪIďm��GC[���vN7.n^�>֣{��\v��
��D�,K�k��n%�bX����I��%�bs�צ��>���%�}�߳��Kı<~��O�%�nrLB��Mı,K���i7���LD�;���4��bX�%��~Γq,K���k�I���T�K���&�'��dVڳ����&q3����I��%�b^��Γq,K�����I��%�bs���&�X�%��{���:��������g?���L{߿gI��%�b~�{_��q,K���Mı,K��4��bX���i�6?[
���Ke����g8X���zi7ı,N{�٤�Kı=���I��%�b^��Γq,K8����G7O�|����v*F��H�i۔�$�wN�t�%�wA�6n�l����Mgv�wO&0�j��u�R�c��u��;m틞��VR�[�z+���m��%v��Ñ.��؜���[qBe��8�����cf�\/OWr��e�ezu�sC����{gY�3>�]�Lr0;enލ�3 Y.���,�����Awk3h���E�ʴDϝ��+�������}w�|�ۖ�<9EMuq��O8�G\j�v���ɜBY��\M+�yv����n�9�.q���ı,O���٤�Kı9���I��%�b^��Γq,K���k�I��%�b^��$�0d�7��3�I��%�bs�צ�q,Kľ���&�X�%�Ӟצ�q,K����M��)���b~�Oڒ��)�L�ɜ�3I��%�b_߿~Γq,K���k�I��%�b{���&�X�%��w^�Mı,K�N��1F�����nq~8���&qj��p�Kı=�{f�q,K�绯M&�X�%�}�{:Mı,K��tz9!S���q~8���&q{}��I��%�bs�צ�q,Kľ｝&�X�%�Ӟצ�q,K��'��T�I�M�tѷDm� 62s�u�����mb����v��\�0�ь�94��bX�'=�zi7ı,K�{��n%�bX�9�zi7ı,N��٤�Kı=������s���&	1�fi7ı,K�{��n^*@�"�#'��M;���'��_M&�X�%��{�4��bX���<g㉜L�g�O8��*�L��q��7ı,N���4��bX�'}�l�n%�bX��u��Kı/}�gI��%�bs�/�&�I���9�.q���Kı;�{f�q,K�绯M&�X�%�{�{:Mı,K�=�M&�X�%�x{޴�����g9��M&�X�%��w^�Mı,K���t��bX�'N{^�Mı,K���i7ı,Oȉ�j��[k��cx�ez�h�g��'d�<c�����N>�.��Qw[�vC�뛩�׻�%�bX�߿~Γq,K���k�I��%�bw���&�X�%��w^�O�8���/��<��nPh�X���ı,K�=�M&�X�%��{�4��bX�'=�zi7ı,K�{��㉜L�g�����LVʜ��&�X�%��{�4��bX�'=�zi7����)��'AB"lTCF�j%���gI��%�bx��~�W㉜L�gw��ByY\u�喬Mı,K��4��bX�%���7ı,N���4��bX�'}�l�/�8���/z��N�e��I,�n%�bX������Kİ�������4�D�,K߿~٤�KĒk�.�)!I
H[��d&�GP�ø.��v�}u<)��{jC���t7A�����4�FX��I�5������,N���4��bX�'��l�n%�bX��u��Kı/��gI��#8����~�����v�N�g㉉bX��}�I��%�bs�צ�q,Kľ罝&�X�%�Ӟצ�q,Kļ=�ZI
`�s1���94��bX�'=�zi7ı,K�{��n%�bX�9�zi7ı,Ow�٤�S8���/y�8�V5T��L��qX�%�}�{:Mı,K�=�M&�X�%����4��bX�@T�*D!�����G�}����n%�bX��c36�fJL��s��7ı,N���4��bX�'��l�n%�bX��u��Kı/��gI��%�bs�0c	���
�.s�ju���db"H9&�N���X�g��Q.��Mø�i7ı,Ow�٤�Kı9���I��%�b_s�Γq,K���k�q~8���&qw|�(�'������ri7ı,N{���n%�bX�c��4��bX�'N{^�Mı,K��i7�*b%���O�1.K�g%��6�8��n%�bX���߱��Kı:s���n%��b&"{���I��%�bw���i7ı,O���C�3fi�8��q�i7ı,N���4��bX�'{�l�n%�bX��u��Kı>�}��Kı9Ζ���fs3L\���f�q,K��{�Mı,K��4��bX�'�Ͻt��bX�'N{^�Mı,K�u 
�H��H�9�-��&c��D�Qm16Q���7�2�����ӎ���n6-����m��x�c<@�h^unפ�jN�`���:���;�3���.�j�^l�mU�c=�Ɓ���u�\�
�we큶8S.�eY��<&���Y���Պ���#:�8|�(��{+���y[ݸ���s�+��]r�c�$*��,9�z�W �;�"m�ska�X���*�p :A0M`1m�Vd��T+�k���Ø�9�۟;��]��)=�5q��:�E&6�MES��Z�����+�����4��bX�'�Ͻt��bX�'N{^�Mı,K��i7�3��[�؇�n�UJ���/�8�K�g޺Mı,K�=�M&�X�%����4��bX�'=�zi7�3��]�sɩF�CN�`ݯ8�LK���k�I��%�bw���&�X�%��w^�Mı,K�{�Ɠq)��&qj�<^�HT�l��;)�_�%�bw���&�X�%��g��Mı,K�{�Ɠq,K���k�I���&q3���x���VVJ*떬��ı,N{���n%�bX�c��4��bX�'N{^�Mı,K��i7ı,O��ڳ�~�L�8�&&1$VNq�q�8�Pv�eݫ-w\;X��\ܦe���u�i�<���������ow1���i7ı,N���4��bX�'{�l�~},K����I��%�L���)�µ*�r�3����'���k�I�k�0��h`1�U,�d	RɂB�6�'�,Oߵ͚Mı,K��k�I��%�b}�{��n%�bX������J�- Ӳ����g8���}�I��%�bs�צ�q,K������Kı:s���n%�bS��Oz4j*�%�r՜_�&q3��绯M&�X�%��=�cI��%�bt���Kı;��f�q,K�-�~c���H*�V�g㉜L�>ǽ�i7ı,N���4��bX�'{�l�n%�bX��u��KǍ�?7�� ��ܽ�5��[��r=h5�B�p>��V��q�	D�t�i1%�[L�9��8�n%�bX�9�zi7ı,N��٤�Kı9���I��%�b}���I��%�bw���f��,3�d���34��bX�'{�l�n%�bX��u��Kı>�}��Kı:s���n%�bX�s޷fbKed���j�/�8���.�s�q~8X�%��=�cI��=u"B��D���}f��M&�X�%����4��bX�'��_Ź&q����s�fi7ı,O��{Mı,K�=�M&�X�%����4��bX�'=�zi7ı,NϬ�./��L�1��8�n%�bX�9�zi7ı,N��٤�Kı9���I��%�bs����Kı?���ع�1rs��;�*�AY�3v���
�#gp4�!�a�m��猝�Sƭ��M���{ŉbX����4��bX�'=�zi7ı,Nc��4��bX�'N{^�M�&q3��O�{ѠQT�mM�Vq~�bX�'=�zi7ı,Nc��4��bX�'N{^�Mı,K���i?L�g8����ͺAU*�S8�D�,K����&�X�%�Ӟצ�q,K��}�Mı,K��4��&q3��_v��,+r��R�v���K�� @�O���I��%�b{߿l�n%�bX��{��K��|w�J�H�*�Ic�-0�>D֢{���i7ı,O�h�nq���9�K�\�3I��%�bw���&�X�%��w��n%�bX�ǽ�i7ı,N���4��bX�'NtװfB/[�Sۢ��r�{v���7��On����Q�1�.yui�6芻��%�bX��}�&�X�%��{�Ɠq,K���k�A��D�K���~������&q3�����F�,�I�۝&�X�%��{�Ɠp�1�LD�<w��M&�X�%��~��I��%�bs�����bX�'g�c��&i����q�i7ı,N���4��bX�'{�l�n%�bX��}�&�X�%��{�Ɠq,K��:_�3��Lc&%.q���K��=�߾4��bX�'{����bX�'1�{Mı,K�=�M&�X�%�y��b�B�2S9�Kq��Mı,K�﷤�Kİ�~J�?�~Ƅ�I�~�j	 ��{�BH$��U��*�eATU�pEQV�*���PU�"����E_�(�  DX
*���TU�pEQW�*��Uh"���ATU������U�"���E_��*�J
��������PVI��N�h�@��@���Y�l���6��*�(�m5� �>�1��eP�
    TY�6dx>��$��P��h�h��Ņ%P �P �J�E� ��wOh�  #�����Vl�Ƕw��j��[2g�ׁxg,� { �� P0 :_p��nÝ0�j�:Η�˳/v;������ z�o�!�NF�m��44ѡ�R����
���%�+Z��顫SJ�\�95�t�P���H���
�d-������N��hi�����_{;�������{�|���C�R��F�=�7����(r���t<���械�[:h(]N��(n⋆���!�x=�����| � m��r«�ӗv;���Z�{�aO�ΌZ��+�M4kBXr馝5��HB��!EL���%J�      �z�U        ��T���P# ѣL�M4�2h5?F�C)J�`20	� �d�H�J�CS	&����j2 L�@T�"&�ROT�SSԙ��<Q��A������������?�?�?��_�=�\R�� "�M,?�芈�aTV�͇�����n���t�w�W�;�淘ZS���9g�����|F�-�63a-�G��OW��:}�<���V^�tN��W����Q�	?���ID��?������[js��V0�E� RE
LB��i��;|%Y�ʐa0a"��8k����ZA�
b%$$`3J��1�/e"V"��(�5t��	�׊�i��_	̓˼e$��i2�8�5E=9����͎��dM#�h���v��s����+��\�F40#d��F���w�s1D�����BD��haV�)�o{��+�g5�[�ec6V��˲�Ư�Hq��$��P�g�gD2t1����FHRVgY2r]� �B�S�j�Tɫ���l#R�A�������g�fx�W��+9al�Ωf��PJ=k	���sM3���]��AD"$E�8�2��0��H�!B^.4X�5��L*�QV�c�[JcU��gX�M�2�x|jy�-Y[�N%9���1)�g����$"�2Xc; c��S���n.�,�E�gG��˴�����V��M��ϖ��D��a�ZE��3�h˨�̋x'i�,-�t���*�U�e�ٓF��!��Na��Ƌ�b�&y��ː�)�h���,f:�.gm��S}]���ջ��A�+f/:тV�#��r�%4uP�X�]d����OR���2�Bi.��Å���	L�(�y���֔"�hEl���Ex|�t�'^'�v�Mi�mj�B5f�l�5Ҫc:�F\�8$��R�&MCc�T��;�nAaNp+Yrp�0kl��F�l��Ljl�ɻ��qJ.Xe`�p���m"��Y
�s�u3��-�9�P�7Xڼ8pt����r�ed�zh�MJ�lC	aLR��A�$h��d�(�I���ޘS*�g�0f.u����s��]y����Y͓��i�b�M,[�mf(�A�Q��Z�q�Ua�J�e%���WcB@�Qa,-�O��>����:�S��fш���p���m���[�WG[���,z��!���{��}�����<?y�ϥ�K�;�4��Z�բ�X��������~����|��xd�wMav�w�A�)d)�!D��T�tJ5P��x�bX	"s9*��]W/vr��㋾CWx3��y�]� !`�I��9n-ŷ��&��g-�ӄr�9��h�q8։Ģ�#p�cCwD*�a�Z�눛�m{�XB�k,f��TY1U�Lp&��(���ԹL�RN;\,�&�������-c�޹��r�:ˤ�h��kM-����'6ˎt��%�Rދ42��y��&��e5�U�B�L�/�S32���w�;983k���xo�?_ĺ~�B��4�3�Vb�jV����C��W���
������;a�bb��g˳�U��1A
j�eB%�Yd�l�t�.f��[�	f)�&��\H=�&��M~HX7�HXwX�;�vi ��k~�Wvd�aN�m�i���ahk�k��Vw�gn�_�.��<7�M��FV��0��.�Z��!%��O���X��3�S�btVP��S�k�Cq�GB?��~[v _�����+���eΗP�b�k�,�;/gB�V��f|٧zA�w�wD�Gw��'{ޏ~G������~KteAYХX��W)&39���7`',�S���p,{4e��=!��G��O��E��n��4���U���O�z ?.ԿHXM�]*К5>|zq�ߌ��O�43ie�E�h�P�����ܒ54!,�0B��R9�s:=�4��̋JѺ74#�"�������>t���Y1�s�a�x����0���[o��Bk., �Xfe�ۜ�t�����<��^�7�c�2K��Kt��Y��	a/f��U.��;z����|������Πs���,�k�M�I��u�!�M�T�;Y��;K;4�C/N4�{2�������ý�w-�.���ѻ�c��_ӳ�M�~��s1�n���y���S�߃�U��a��~w�����gz��;��{{;�R�a-�w����yq��;�{����Yl�9�厉�~Bȧe�xM4���pr�&%�a�g�AQ&,f�v�&�/eYot��S�6i���=���%�3�h[>Jw�3yy~'u����(�wK>���-n�P�~�r~����f��'m���e	�z!t��7w@�X���(����/.�:A)f��Xv�{���Y�<Ӥt�C�zq��=9��JΙ����Zpd�C9�rI��c�̀C]Ӑ.l����:b7�y����|�,&�9�K��:[ww;�<�h�l��!���Xv�W�zK�w^[������^�t۷����p�s�,�'I��SRJ@�L�)�Ft��{�p��[ٙ^�z��p\�ִS-��l��^35Ul�� ����wb�̊�E�v��e]�+�٭�{śģEj=���䩧r�W9�#�I���}���;^���[�*$:�eQ*B;	�h�7�p�Q�@�(��@䌌���!3[Խ��J�n�i�3��@������3�f�Z���P�(�ۣ��WIzXp�P�*��{�~���N�8k��%�,�Ж���L@��!�i5wxIc%e��K�����x��kE�f��v��je_IbgY�����E��{~
�r�j�2�$/8�XM�sE��r�,  O'�tpVJo��N��C/��a���B��UH�}}�e�`G�A�y�.���ސ��K��T�k�d�߹��ޥC�)��ɴ�oX�UY�e�otjr�W��1Zɘ\�̕��o��F��1����DxJ~��^6�*���@@�GC�ʪ�)�ΑU���3�~�}���yRC;�����S���5�B��I�����j�H��x����窪#�_��4�2Q�X����ߟ�~2~FO�ٿ��c�1UX�               Y@       � �  �86ؽ�p�x�M�`�;����Y��;'Ԛu��QT���8T"۪�NxS�b�N��������ۖ����g�(�&���46����HCK�a�jqUGef�Օb��@��rOn���*�,pK�4vr^��ݫu�����Bϑ�]]]�z��l� �'�P��'=�8w-�r')aHk�@���"}m6�B@.�T���Um���Z�eZ���`�ꀫjP �G>x���S��D�X'�W<�������[����*ع�  �v��6�m���p���v����N�>>|�����_9�So�/k�n����G�n���tM�d� q�6�m�$ &�4lt�+��d
��^y%�M908X��)Ѳ��He_@Z����f�ҵmT�Ǭ����ʫ@O�\���K-�3��5؄ք	t� ��)��MB�%� �R�퓜K�\�Ћ7hv����X.��i����S�v�g�^�l��v]Y�k����`�t�Ϋ�;8���P�SLJ�+�F;s��WFPZ0ʤ1-p:����c�#�-���nq�R3l��S��ٓ
��Xܓ��[���\����8]1����bC��]cvx�p[kb�-bc��a8�Xl�YǍ�ƺc
j���3�!v)�NB�B#���'�*����Ҳ��{v�N:����v̈��f�� �#I�n�n�`�>9W���Bm��i�%�����k�����q����|�|�*�b�����R)Ϥ�`Wk�%E^�<��^hĻMR0�X�	���Ѥ732q]iҥ��q��\{u�s`5�'Sr��J^G<�L��Cf�>�1u�5�捴r�f����SR����⪑�v��+�� vu�.F9)�Re2�uM4������z6۸��F��

m��VCF)�͊�3�v.��B2Օ��31���)@����T���N]���m��4卞7K�݃���7 +�X ���PUJf� �h���+u��'g�Рɋ@�R�p��-3��@Iz���댑˛�f�ˉ�@��2�^�/Y���%;�%�9�����q�S����kh@հ [x  ���v�����l�` �m�u��m�ڲ� ���3n;5<27+�+�D�cb��v�]�r��*�KR��j��vn��3�M���:�`�Z���r�J�B"bԃmm�e*�JUP8@!���h6˰����[lm�6�8x c0�̅Ŷ�8�VA��h)��V��p����U�hGm���3��j$�����z�<��s�e;�˛uӦ�c\��X�3Ki�-���̽y��p�:w\6��W���S�9���vg�0�;>���@'Y\��^k�uBu�nR��DL��\���m��0k�v	���;q��L�2K5�c�؆�҂�mE�����׽��ݍ��m)B;eP6�S� H</��[��k�Mk���l�&�m�L 	���e� m�� �t��6���-��5J�p���ܫ�v�+0 ���    �m}�:m�n� l�mmuWUU�j�*��L��I�yŭ
�}s��Ek� ݰ�`��e��W+=Q�Cm��5� ΋;�����yugq�jϠtf��V�g�]�Z�u�ϚکV������r!�5C����pp�!5*�R��%q�x��U���7@p�/]�^6�c���n0 ��j�]����6d���nM��  ��5���$my���U�k:g%���p-�hp:�:[vH �n]���m��ݬ�I��wko6� ��"��6ŷ��  N�S�ݲKh �f՛v�gK:Q��-�В�m��@-�N���� -��͵�sm�M�Y��fZH$��5�m����n�I  ��`l :�L����*W�w�J�ʵUmr�>iU�8jj�B�6݀�۶<v�ojO�g{�θy%QC�P.�Gl1��ѵ�u �b���aݕh͒�}R�h�Hp�m�V` I;m����d�-am  m��$M����:-����`$�	�  WIL [m�n��F�ҜM�ݰ�a��m#I�i�l�dx����H o�z�l�0 �n�����0mpt��X�Ͷ R���mp�bj���l�P
�t�"�7.� ��7R�����Yc�L4��
ࢮ��0��o�|�1��x��r��I �
�av�$��.Hj���r�3m�@��;@pW*���U�#��a�kX����m���%VT!��\  m�� I�ăn��v�Hl�d0�[o\ hր  �� ��"�`]6�c� � 6�l��U�v�iV�	`���l�   [@�m�8H�X6��m 'n� �vM��J��Y����Jɣj�F�a��	����l�0��lKzq;^�7Ik$ RJ��ukz����z�k�p �R�!3i7 9�f�nqcS6���8�u�-�.�!��k�i08[D� -�m����pl �)%u,gK�0a�+v�"��Т(�H�t��(�(dPO�ʏ�u��0/��9D�J~@�D(F�W` �2]
��jȩ�fE�Y�#-��pw�Hd4��[� ��hN��hi��$��Cj#NȤ0�@�I��P��bu�Y�B'R���H$�:����d*��r1!L��v	΅��9� ���`�� 6`yba��FtН@G�D�SeB�m�F*:1F
EF�o-޲o�A��l�J
�ڇiИR(u8��8��\��S�)Ch�� SB���n���#�E�a8�&P2+��u,E��&�c!�
�"�A�
؂@iAN��S���6��]�*H ��!�%A����\+ܚp pU
]�a]�fA�g�px6�! ��!4m,2��U��m�`-�$BI��MHE�]E*�[�f����N&����Z���`WKb)�j�8`FB����t0Ev)��#��f�6J��i����������י��3���-�D�H��sf�FygLxx�:��Ϡ3a!_�L����I���,3��,󐜐''r99,�~|UQ\���l �!�u�2k�͓K�a ��<vxXB�ꖚ�2�,
e�����u�Ӥ�J�܆��n��]���um����\��L�E!mنnt͠$�;%�!�j�8�b:햀5u�\=�c�\p�p�60��w*@�M�5�6�t�nzT;���9;I��vM0��X��%KX�q1\�l7����=bz� �]����������5a�}���\s�tL���ѭ6q���UR���k��q+�(���a���yY������\6�8�,[P7T���˷n��bƚtl��6�y�,�ѭ`�>�\�M#��Dl,��J��g�*��R�6�Us�]]9N^\gB�##�kQ�i���`�:�sl[�*��\S�A^�F���1�S�v�G��m�-u�`*ãx6^׳I�K%�qs
l6�ͮ�gD�ʜݚv���]��܄�+�V�ܝ�P�+VN6�9|���H fI�\�&]rnw*+(UY�ab]����کEV��x딤�"�	��q�=�����]I�r�;M���@Z��A>��|	�Dz���e&�)<�D6�E`�&P(�toļ^%Y���'0�u��!t6�����z�үQցwe�'Lv���9��T���@R�\8��3bRn(ۀpJ�VB��ݎ��*��9��q*�Y�&�y:��c<����*�P��Ch\cZ�%�g
���a��6�C��55T�����,z#���$
��05��Ī��>B��wu��yt$u��:|#>���FD'+�;M+�I�#=�dB�fA�U^V.�p�#�B�fH����� ~ŝ ��f��� �V�,�]e�%�������w>yNs�]�1VV
ɾ��2D( 
�&#H,,���`�HY�F�v���qn=O{G�pKtۧwM�#=�4V��g�U���U�|>�s��1{U�^��Uh�|�;��b?&,{uuWw`R���UU�5�Q��AZ.�6����d&�G�Y���u���4��&d�����c�t�����qL �����ca0�2!|�2F{� ��VHϳ�{ȉWn�A5i��S\�Z�1i��X���ڵI�wt���ȉ�`�Qd·b��'1��{�ڏu5S�d�T��ԣ���}��'� O.����M>H�'�� ��"d��!�GbP��(�jv�Wb� �l`�@"$���y��/�ib�S1���r��G�,1�3n	�v-�^��~�Ⱥ�(㽴�=�X���]�e�U�Q �:�&H�'� M�TX-0݇�A��y�Ob � ��]���wulC�N���P/�J8��<���U+�Ld��y�QϽ`���F���y�I�����MDդ��-B\������I��/k�����뫣�l]�k�с5#Tv�m��n��4�s�i�)�Z*z��j�.���I'd�6e�Zj̇ ����R�b���F(�lnk��i�ˋ�J��~:�>+OSt�ME�g;������_��q�X/��X.�@�ē���V�	$`�PzF9�wQ �8�]��ؤ�&H�'��&DH7#�Mv�w*���y ���k ��`��Ll&�@"$s�d�y�ਘKV��S�tP�t�M����V���t<�ʏy���`��'�"��J>=�x%YW��_{��6 ��8qF(�%j�}�Q�ujqH���W<]Ub�s�{�g����q��_]pɚ���'�R�����>�\bI���+yQ�;h>#���u���Gǵzd�J�ʗZ�ְ��(5��dTť�i�m�wT���ȉr0/:k�˹Ux%d}�]n����2F	<���a�$2"A�:�=
:�#�]��t�fn�b�]༨w��'��<�dD��j�L'b�L��O1 L��g# ��v:
��A#d5�uF����Ц�U+�I+v��9�"A�����wr}w8d���P(CZ݂��֣���̝��/��;5�N{̐y[@"$�$��J�X/{�Q���i� 3�hG�sv������������A��d�f��R�Um�к�N�9�94��D;���K�Ɋ���(�:�^�������N��\��yQ�;`��-G3����h�+	ػ`$d��� � �F<�R��U[�W�Aʔ9��g# �#$8�O��pɊ+ޥ�V�z�s;i��
�T7�������Y1uE��Pn� �Q��ۃG[����;���-��{I��5�ઽ�nr�:��(2�_`C���q�v��xk�d����&��g���;)�6���� eە�)�Cf����<�:v��1�����ȶ
2%�ŷ7M�-�wJ�j��_	d`��$T�	��qT�I]�&2FH<��	��X����n�\ ��=�H3��L��O;1��wI L��{ΰ	�0	�@�ʩ�Ӧ�>�`�� �D2"A�|�nӵA]�	�]�3���0����]D�x�U����\�{��V*{^�]wu^�%I���d~� ډ���
�iF����j:Ϗ��pɊ����GYՂ�ް\��o+�b�V���=��'� L��}��t��T���ȉr0	��y�����]+�3Y�y��E�Qn¢��5���ٖ����퓇��y�d�yٍ�úHd@"�����`��)� kړ�1W.�^T}�X.��EOАo'@b�$#��X1TPX� ����L�H-"����-D,h�h��R�!Ůn�aØ�s������)Ԥ�G]�t�'��8��9���ֲ%+���%ZM�8����bI#)*�Uoy�?��x!�w�I�	�	���ʎѳhh؊E�m2 atAihx��� |@L�Y��iG�4k��i�L����&DH3��F�T	 ��H$�H$�k��_�tL^.cϖS)��d�L�S)��e2�L�)��e2�L�S)�����e2�L�S)��2�L�S)��e2�&V�e2���]2�L�S$�e2�L�S)��d�L�S)��e2�L���n�L�S)��e2�L�)��e2�L�S)�e2�L�{���L�S)�e2�L�S)��e2L�S)��e2�L�^=�?�pV��g��WE�
J�J[-��lt��	���L�S)��d�L�S)��e2�L�)��e3߾�e2�L�I��e2�L�S)��2�L�S)��e2����l�S)��e2�L�I��e2�L�S)��2�L�S=���l�S+e2L�S)��e2�L�I��e2�L�S)��>�t�e2�L�S)��d�L�S)��e2� ��H$�H$�c=������ƴe2�L�I��e2�L�S)��2�L�S)��e2����n�L�S)���L�S$�e2�L�S)��d�L�S)��~{��e2�&S)��e2�L�S$�e2�L�S)��g�}:e2�L�S)��e2L�S)��e2�L�I��e2���]2�L�S$�e2�G��92�L�S$�e2�L�S)��g�7S�ʪ�*U�A$A$A$e2�L�)��e2�L�S)�e2�L�}}}w�)��e2L�S)��e2�L�I��e2�L�S)��>�t�e2�L�S)��d�L��e2�L�S)�e2�L�}}u�)��e2L�S)��e2�L�I��e2�L�S)��~}���e2�L�S)��2�L�S)��e2�&S	 �	�nz�X*�V�$�H$��I��e2�L�S)��6)��e2�L�S)�����e2�L�S)��2�L�S)��e2�&S)��gǮ�e2�L�I��e2�L�S)��2�L�S)��e2����n�L�S)��e2�L�)��e1 �	 �Bc�O�rOn�v٩��e2�L����L�S)��e2�L�S)��e2�L�S)��e2�o�z�:]�e2�L�S)��e2�L�S)��e2�L�S)��g��]2�L�S)��e2�L�S)��e2�L�I�*��~��y���Ns�^������7�(�e��\�E�a��p���סލ��_^YL�S)��e2�L�S)��e2�L�S)��e2��߾�e2�L�S)��e2�L�S)��e2�L�S)��gǯ��e2�L�S)��e2�L�S)��e2�L�S)��g�}t�e2��S)��e2�L�S)��e2�L�S)��g�}t�e2�L�S)��e2�L�S)��e2�L�S)�ϟ7�|x�t��w���e2�L�S)��e2�L�S)��e����pC<�z�1�݉����/�tL^.c(;�/ �9H��=����`Ew�U\0b�XH	�R��GL�����h���j�g*�b��,C���|��֜H	��B� �� ���	G��������P�mN�$�lA0"��M��uۇ��\qƪQQ'X��^��ِN��*�܈�1Q�3������6�*L�ǚ��Gzu�N����`^��k]';Rn�W<�Aݵm#ףeV,=X{!#$��'%�&�~L�VjhńK�XJ���:3�G��b�bUV1UV!�`��r�s�)>�R%��݂�۞���]��o��ReB
{۴L)�������VY0���(�{�ҰS���aX9��ړ�1v]༡� ����;i�`�}H��}�Q���%�w��������#���`��R��}��8rN|��ǘ.�G3m��`��� �L����3��i�o��P�">��>@B*}��p�<��UWL����(M$(�s��}j9���D�K�<�+W�A�� ��#�2A�;D���w�-�I]�-� ��`��$s�wP�Q'w���-�n�\ �C~�]�"AO{v�ź�}�ߏ� 1망g�X��WNqk��y
��t��쇾��v��>��G>�4�^ԛ�����YQ��`u &��AϫIz��Ol��w��+8}�Y���!�� �`_����7���}F{��5����-n�_Fk>���;���RIxpUճ��̳��+��Đs|��һ�4)Q�ra�mh:�\���*���t�^���Ϥx@�|� P�LT�U-�i]�����5  Wb?|�M}�< �}����J��U�ߩ�2%�I�z�{ײ��K�VI� 	=�5���z̀'������ϵ':b����}߬p!�w	�S�VP�!���^l��@UT��e�V��[T-���p[a�l�����������=���]5j�_�����{�wu�f���W�B��8O{�> �2����ե!���%\�V2i>���H�u�n��m-��m�Rc��`r� ����n��HӯN~��P蕺��t����v:S��'2��'Q(c�o"9zm��8s��
�m���s��g<��F�'�%zn�gsc#�.샕r��XS�n;C:f��ge��0_(��p:�����{#����jX��V�A���ʺʗ��tg3�۽����s~����kס� ���(�5�r�UY&z��Zݾ��`�^���o����:Iٶs��]��47i����]�x1��$��O{�k�iF{�X�� '��Q�𧻓���W��G�A����;��$
�V1��V�Ûs3ˉ����.'[x�%c*��Y(�1E��V�f��}�l�5�q�;��W/���h�H!����P¡�S�À8lp"�|͟j�Ͼ�T�c>���uI�n��w|,o5����a7a.B���� �ر[���w��VpV_z���8����t���꺆�Vh��笨ڱ�fN�RI �Z�N닂��|��s�N�����r鰝��wu��G���yCs���ĺ�b�2{��u��"b�H�󏹋~��c_�كr�0�>����� �o�SkԛWW���t��,w��}��~]�ة5v��vh�A���ť���n����wP�ڛ��vv����/u�##���$�U��:̑�Dy&*��vH�s�v!e�I���ʩ.�	ػg�2y�Ȅ�g;]P��-a�(�!)X���,��[T�wMض��u|�C܌��	`���ّ���EةR�v��=�y�b2!s��ն�����u��;�{��fa7a.j=�.Fd�%���N��dpZ�D�a&]�XL���\xݓD����Lbf
��cF $nIew�p���l! O������v�K�>� �K�K��>��eĖ�d�1��3�6�:��|�1�c�m���m�����L�㓛�ʏ�V�v��R�;Kk!���aH�\u�sБ2�E�`����a��ĵ<Kfض+	W������-�=V���g�1tq�Y0q��{���ψ�Fݔ��ѧ��i��J9�t��7n5���5�Ǎ9T�[�na7F	W�.���!����D��e)�^CL��Dp*;;W4&R��BZ�V ���><aq������$�]s�f����}�!m�L9Z�Ar��6�1�G���G� +l���6�p��WیK)͠�����f�Pf�X��[�f�
�cYB1�n��QZ��c]����X����\FiV��k�u��m
1N����t�o�`@�H�Dp�Ų�E�v��I�vM��G,�9�C5���nU���*66�5C]���+c�[z�nwi �P����\���m�U�s�O����8ڕ�Jl��Llܒ#Mq�\�i�W)u�\��4y�(�uˡ5Kyw7F�yU^��ڇ�jz��MX��sJ��Fi��Y�[
����{h�Pr��w]�fJ�*��0�������9N�P���NXVm�gm��: x6x'�-S:@mڥ�����%�Ǐƴ���h�����l�`S�-A�UؗDel�5n�.\R�eZ�Xӹ��=sf.���j�'��V�LE���B�9��S�v�8�.͡�U??�k�u:B�ړk-b*��r��Â���@�)�gE�\�Q��ub��L��B�]==i�Ӥ����B��rk=��LUi��>��@��j;��*��M���ْ3�C@��9�����j�۫������̑���S~[V�� �:��،|��%*�[s5tf�M���L�M\�k�d�{>����߷>DdB�K�m;T��6 c�Gu�Cf�Fźv����@�$`r�2�L;���s�fHƂH�G�;��i��>����<�ȇ��Z�ݫ���&:�Ӯ��l�֗�[a%lS���v.ْ3�FM$X#{����Ъ»u|9������+�=�]��u��S��g:��{'f<����:����ҵ|� �~᛬��9�H_|�wmն��L�� +���y�7<�>�K�׎ZEH�a�i][����7�$����d%��G���^�������;����k��wu�j�44sk���>��s��;�ފ��6�v���FD:>" �E +�d	�8U��@>5�����}�K�W�����0��@��TߟK*���eJ2�ܪ��2R�+
nU/���|�&����P;ߊ������\�_9�J��~���KO�x�}�Ҁ��{��d.�y�|�p����~��׻G��}������y�Ş��t�*��*��AD��*�woI�U�,Ca����s\�114�pt�+��lv:뒋f�և�;��ݷX_�8Y�ݞ[��P�H��vsDp�ѹ�e�t[��Eq�n˺��g�6���0fV���ikN��X��)pY�㒰�l7i�{��ć�|��h�9'Ab�t��P�˸ZGv6f?���(�n �vy~Ef�]�<����������{��߾�
�w@>�p҄�w��<P;��/��|�v�ҁ��P=�� ���=��T�N�����(�. ���#T\��F��f Κ20,nM�J,�.���x�?\�y w���|��8̷t�^O��E�I�RN{Xē^�1�B�C��tJ̖�Ҁ��ﾨ�.������C�{�P>��@>�p� ���+6Q��<PN}�p���Ϟy���
6U�9�]j�O�����˸(1��v����ˀ>��<�@�K�������@{�@��T� ��}R���&��bI�s���4:4:��\�zP���v�]�?{�|�p�y/}��{G��~������y���r{��-��.�.K�	`�t�M;��q.�x
�%� =(���}P�\����7M�������(�. �t<���]�<�� ���
��@�g��4s���� �P<|Pڍ_�\���x	����&��U�������Ҁs�~d}�@<�p�I$�����WF�7,4�E�#�3X�����x�V��=����� ����_:.���x����@��@�矯v�3-����J���x�����L4���@��@��/�������fc�y�������<(�$g��{�L��7af�h�Wkw�SN�`�L���j{Ys�r��v�q�̚6�VY���^�"���3Sq�hXFƒ�4aG���.�I�m6l�� j�P�)�ʵ���Ħ����rzK�|���ǌ��	�XAN;7/� �Ӈj�yn�������0�@��@?_����y�����<_�KO��[���'{�� ?�_������`��n+S�y��������Nr�J�K�E�!w@��T��<(>(����YlMt�1c7J���d��i�S7v77�G����`�����}�@=?~�\W	od�ұ�EX��!J�`�e��K;*�����c���J�j���ZE����V����UZIU���RJ�*�M
����e��J�� "�;S�wU_O�ꪦ'U]\��Nl�t>��|��O��I9����� ���9�1w@������0�y�s���ޠ}��\;�{y��r�0���������6nU%�����b�jۢ��B�Ӓr����=�O��@�������rs�v���߁�O�Z��>{��������s���K��ְ^�ﾨNW%�:Y�Lg��L�(�����gV�)ɑ	�AY2��`S( `��T b���er`����x��ǌqΔͩո��G\��:�lJ�ef�j���:AZ�֣IE����[78�!ű5���B$�E:��B֜+;﮺�$��+H�Z���.ha�R��`@L�qQ�(S�P�
U�v&��
lM(d� 88Q�P8�R$��)A��ӯ \;@��ܝ�$�y�I;��׻G�����n �P7����x|�lZ�@<(�~}�@��To� =��[�e��2�g%�L6���)i.��9r�v�0��}�@���{���rq�}��~z_���Gt����\�ˀ|�}�r����{���/@=���n?�!-����}wU\�*��E�K�Z
���߿����	�O\~yJ߷Zҵʪ�uU�'9UU�:���uU�����z�����6K��\a�qu����YѺ�_�y����\�����ﾨ���ݣ��w@=���n���/����/��-����꟎Sﾨ�\����v�0ס�'�������z�߮ ��p��c����|�@�������� �(|����?�d2˔FsKm��8	��^����+Y�L�T��2�̢E�]+51���Õo(��lK����49T��I�]/oF�ܱ�Gk�3� ��:�&m�l1f\�bY��ܨ[f�[��Re?���y�8�	��Sc�6,5��N�f�KS�zL��T�ݘҮ����>��z�|���}���#ݛ~ y��С߿�����뼖���+�Vԭ�}�@����$��c�ۀ?\����-Ղ�������<�=���z���|��8̷t�.�r��P;��}P~ϥ��~:/KZ]h�Rq��0�aD�לE���%� ���?>�<���v���ϓ���l�^���WP�l������|���{�bH~�p����~Ŗ�w@����Ǽ���n����~�e4��t?O R���RI�U�=�6��k��$���_�O��Ϳ <����羨��������F�ݮE��,$8se*f�D��9�r]�ݻ�R�RM��ē\�1$��x1RM��I�Ox�n��}�� ����\���V�b�b�;	>UUn�UU�N�.�"H�W����<	�_��$������ص�o@?\����4؝Ub�m��S\�����V��� �ˀ>{p_�&��+�J�1��Yn�F:�/�8	�Ef�;�}�� ����_�?�'g&����y���
�w@���rZ\}�@���>����;ܴ�� �����-����{|0}���ڕ�Ӎo��$��q�&�e��E��XEu�q��C�ӥ��^���d���� }���y���1��E�΂�����2+�$o�{�|�8̷|�t�>�}��99�}�@=>�|ص�N�~���->}��}�����s���l�=���k�?{�������<���b鲎�Od����'+��^���%k��$�Ӝ��䫇t���9�s���P>{���T%�&��+^�9���K��U�U�ñ����6���`y�͘è;"��<;�&W*5v�r���&���7�H�n�:Ξ� ��^˰�/m9�X��`�j�^��-����\�EEp�d�M7�9�s���ݵl\�cWff4h3��z��4R����.���'�������;�����P>��!]���o@�����(s��1$�}.I5�ZqP*��'���n��~����`��|�@��ߎ�f[��I9|ޘ��ﾬ�(�TV���Ē}=��\�\���$��ߟT�x�}����z��tz���]N..e�9�O��䜓��ߑ�ن����>�P>�O��rI'p�� ��_"�e�>�8�h���x�W.I7ڹ&{�c�s�Z{~�������>}���uU�.�w����j��ߓ���꫿}wU�H"_S����+q4��z����r}����� |��;Oy���2��ѲqZ�t�e!�h�\_�rJ��Κ������o� |��;��~�wh�2��?_�9h}�p=�@����=>�|خ�$��\�:�12mX@$"�b��/�SS�g�z�.I�2wf*��zܿ�����(o� �������(���y?o��}P>|�޷fX(�D�@W;Gr�4����Z���^���5��/�ꪻ��W7nꫲY�Ŀ7���_��GHc=����>z�w�I�&�Ҵ}��3�Y����j�JՊ� �m�{n�E0.�4���һ���cs���m����4 ĐW�9��w��sߟ'�풵�l�h�ո�[Y�[�0�]����|��<�1���n�����i��SG7��Pf��w�[�W�C?l��c.�n���� 43�{���uֺ�iګc�I�g<�7X��I�}���ވ9v^4��s�ٟz�w����g���1��kHK|~ D-�X0a(�S����c�>�^�����;:���.h�%���c㮘Vf�1l-��I�Q �UV;"W�;�n�V��4�-,�"�$-�id��8�Vp�ܒUQj���jEijT�+iR�t|[ώI$!�Ú,�i����~}�x�����LB4gZ�����2��(����NS�f�|�M��UU�� -�^5�����^ԝ�wf'���2�t�|���ĝ�]�ܫ+U�˷�0�]` ��v��y�j[!a�`��xpmƇ���k�f�3�e�&����B�D��7'��L�gu�6��jx�8L�vMs�6�(J�z��`���Kq��&�Z��f	B\�X�yK����k�1�F�̖�G����Q���+��h;���z�ӴۛP���X��	�9��v畸�������kD���qP��EUg`UVB��f�V�م��9���M�a�^y<pE'Aŭ/��!�c��T�YZ��a��:�a۠M�v#4��^2J�vuX���"�Օ�s��E���w�,rk��犄��Y�Y����ܘہF0���Yz��Q� ��m�f�e��c#��C=
�8��T�Xڃ��q	��Z�w7�4<-/�0�,��AH��3�
��v��k��d��鱐�cf�9���e2�G9c"�e�P+ʪ�{n�]G)���[�-6�Ucsa�<1��=uюWV��o�4]��iP6���^Ut=7����]�`�"�6��h�&QA�/ �ΐ��i�3��]��K��L�Kf�qSc	��׳;�S���R�kv��5d�vҚ�;���#���O/nK�b���Y��(��78+u2279x;>�f�V�rr�V"Rxz�mʕa�߾I�uo~:�d�3���������#�k�{����>(T��c���o��'��#��ߪRT�+�Ͼg��=��G��[��m�mX�ϷY�#��9#2W|��+uV��B��s�su�Ed�2�Z�-0݊h���3����X~���l���v��`T��(f]+�jh�y�\���f�?'�}g��{��A;����Z�꛷V�n�.���su�o���Ŀ�����G���߾g7X�V��6�Ҵsu�f3��k5�tz�j�_n���6�G����,+e�4�R]j��׭y�&U^��.�����m���3H���<�ʑ�V�pmJ<�1r3��Y]�^�n�*>�b���p���u���Q��V:�a���7l�YC�w�ެu����ul��|�G��^�<�
�j�v��'嶸m�ծ����ò~��|�y�}_Q�q����P��9����i]�G7^��r���zn~J0�d�㒪��M��뜿���ܫl[j�&su������X$U�uH��P-��L�!3>�y�}��t��Z���w���;}	��%c��:�re�k��e(Yu���G�ct��9��t~}ǻ�J�7:&:����_dzhg�9��u�hśI:�vճ��{�h��;���w�7��vþ��<�1��>��s�o��bV)߽g�s�w�[�S���DG�r{=�c���Y��7X�T����<]�f�m����X3�d5t��Ȇ-�Ph�,�{i�@zۋ
�g	�.6i4 �]�cV��-�vp���<�+�I��if��s�U��ۭ��YN����'�s��iк�ؠ��v.A�nW@�Z^6t�V*�ϵ������� Ͼc�{�i�ub�����<��H�'�@!���[�a�\;�<�=��=��P�����I�u����{�ܘ1ջ���d���w�s�Y�3Z$�~jLJ��D�Vc�	,q��<B�^������T���}��qI��@���gk?S}>/^4���D@�҆Ǣ�Z8/�c7�G� �I]σM˴���>��f3߾g�]ESMX����ID��n�ߐ�\��&dV��ՊL�	�G��su��I�K��-]�m���ZW�mЎ�Gctt�\\�|2#��#��c+�����i� 	��9����?��A[�N����o��S�J�``�ʑ2}�q�ǇkSB��V��
���yn�� s���~���;a�Oڏ�Gs�9���u�ss��e����U�n!���9-m¶�o>����s�zE��{�գ��V*�3u����#�����Zb�V)33Y�#��9#2Wk�j����g�N��1�Y�N��*���\��-0݆�������gq����G':�3��+a�0�1`WA�[k���2���n|��sϪ���SB��V�Mg1H��� |ܯ~��~�w���<�1�3��F���J���������"��=�Ӓ��c&��|'Ǆ��_�N~�Ρ����$�?�>�5��3a3S����ø:��b���gF���P���^5b;h�Lm%r;<��f܃�V5ҝs�W.��j^l0�ͷG|��@��J'`Ӥx7WpnP
��R2V�B�%���� �� !��of%�(�v��1f�ӯLiq��0Ujջ����V)3��s�ρ���f�B7J��v/��s�su�ev�^�n�H�u��3��f#s�VՇwO��3��3�S��:��h$�U��Fs��\����I�f���uA��a���1Қ3��LW6�SK�nϓ����#��/��_#I�]�um��imRҵ���j����|��f�k��u�Hg'���ujꯃ7Y�|���G{�ovҫmX��泘�������p���50�ե��G�'~�g}�s߾����{k�d6�̤]���:�ӌ�����x>h��vG7X��;��G��kή�'t�;����g|���Z�$�U��v���!�!�L P�`Wy��SL�Q��lb����ZM���9���#f#AlP;m&P�A�9��KXd�*�5I|�D��#1Lق����m$��D�	)!�	E7wm�!��C8Q.�ɜ�:F�J���XHK!�`�F����V���Ϋ�����"�2H�t��x+�!���N"������GLҌ���g����J�_�9�Ə��
�����������c�����Ƃ=�;���<�]Z[�b�ۻB��*h+slt6�%˛s!�����_dg��3�P����iU��Rg��s���	���۫K�u�1{�̌v�Q`��vC@��s<��ҁ�XT+�B���?m}��M]XN��w�g}�g|���<��sKqֹ�0Vݚ���fy�+ۂW7�O���>b8w;���ߴ��1r3�uR��4W8����y�}�;���i62ګ�h�F/1� V�Y�#v5h�j�¾���}fz3������|�ޕ��VڱI�{�s����?i獳1���6�*�SjAu��vt&1�2:MXT2]���D�$�<#`LO5Z�P��nN�՚�������9�xq]Yq��e�F�j��6��m8ƶs�0#�r���6�i�w��z�{��{ǼW2؋�4MiM(L�)V��Ns.�~]�	r�)�v������q���fF;\�`�a�#���3#3ā�$��x}Wj��|��s<�(}�y�Ɗ�F��7n����B��>�7����uR��4W8�����$�N������]�a�m7lyK�.�.���]�@6�4�+b���db��> g5pjӒ�cc&��GV#H,�"��1�em�5(96zo'�ۡ�3������ګmXI���q��wX��vw���;�p�Q�������Vj^�a���� ;�Y�k=�n��/��H�3���&P�n˥b[b8�#��ɻ>���߿�>x�9�����ݻLﵰ(f#���;���>�t��7�x��@��7��8"�YmUҴ{#�321��j<�գ�»�3u�g��F�c�Bc��R����j��6_W[��������Մ�٬�#{��H��|�L7a].Do��$fdEeeV���i�b��W����<ލ�uv�;��^���-���o��@H�`���|)��;�ݜ&��wd�������nF.F{�]�;vұJ�w_�]5w˚���Cz�;��ߠ�8*���F��_�?�
�c�ԓ�&�մ{������^�tV���
�n����"��{��mU��$��g1��'�Y���+K�D_q���<��&������<E��Ci�r����#jۚ�ՖӒ���;a�k��\��0k�CЁ���ר@��V�k-�ͥ�0Z[0F������1�v�L����L�Z�u���%����hm�J�P�=��98s�݅���4]�;t���@�2sX��=8v���i���g���G�*R�ua;����y�����K5['wi��g1���χ:�~��N�/��,���g���g��9�)7�Һ��$b����f#'��"oZ�:����ڜ�g�Ы�I][a
l]!nþ��{��E�ǹږ�[j�L��  G@=#��G��^y�;�<�V��"/��< ]�f�3�[�V�vG��^c2y���pJX.�'t�;#9�31#A����w���k`�%�kZ)���%��i����+w=��Ͽo7��r3�uR��E;������^�2y�Es��k-�um���D!4H��tD�К�ž�7�{f����@�vϤgq�Ǹ;-*�Մ��3�����7?|����f&�p�K�x�,�K�aH��-��f��۞yK�1r3'�ਖ਼V�vG�8�{���3�M�N�j��|��{��"�cݥږ�	��fH�b2�� 誠GFT$HE�ڝ���T��;��������̞f�2�]��V{Q�s��ʬ��c<'I]Z�HRnեumH���� ���T�)v�vFs�fb.F=��iU�v)3$g1##>��^n��ip|n�y�/u�[����z���4�7X�ݽ�-��Ʈ;4 u�&�!�ϷC3�!�Q���Μ� �)�_dA���lc�WD.(h"�b,�\8f���!���X1H0	G$pT��܆��I	¹���ZԶ���,��\�<���!)K
[d-�XJ@�%�R�2\���jU˜����[�ZZT�ˉV����\\Q���Z�.,��s�����rsJիRI%k-+���[��K�Nq,J�Jty
u�vt�*��jd���O�� ��d ����A-�l"���.&��Nv�>�k�n�n�'�X������NZ�"�8[��Ub��Ys�M!ʭ��;9]�.�X�g]C!.���G,h���t���I��@c�[(��p�mm�D)�R90ir)k��`�R��y�/�YX����#aCV0�;2�i��nً7d�u��;�!��U����aq���r�1��<+pۅ�]��+�-�Q��YPN6�GB�4ޓ�!ʬ升	[�\��U�����a^C��Xļ6���P����[c�v�5�	�GM��9�z�Ѥ��m�d-S��d�2q�Am1�D� �SJ�;W3Ĵ;��� ��@�^�O=\:��l�0�n�eێ�Yz�,�����ܧ"����-�3j;b��V�l	��K�)��.'��Ӣ��I9w6رn)V��A�q�.4���s�cT+�2�X�@�DMhɈB�3�T�7"{B�r��q�v�qu���8%�igecT����`ؕxu)�t�	N[VC����L��sɮY������j4�n@�ucWGlD]6��[��$������L��I~*���ڇ@��3+N�N�	j�iEa�O���'�rrY�yy�AC04������l��7F���dv�B؂����\�A2,��
l\��j�Ї�N`n_Whʙ¸�c�����^x��7;�Uɋd�t8����%�;��i��G��UuW��n�Db#��Z1Z�5�]�nB���Eۍ[^Gd�[v�%VZ�mRwOg��y���A P��&R�z�;�L��sr1r3�u%��j����wQ}�/u�<�9M�i][G�1}�d�*b7�R�-�w���y����
�Ǣ���ZWM;�H�cs�F�����(#�
�N�&wu��^�#>�ؼ�+��i�$i� 1�F3��o��ՙWa�#���d�3���I�>$�f��f"�cݥ�qФ��fHƀ�׏��������[ty]���-]mLfQ�LZ����3����wQ}�/u�<�9N��WV��_q�<��]�Pe0݇|����	=Q@�� a@� h��ǽg2k��������sr1����3ez�aXv��_q���<����Ӧ[��n�]�v]�Ӻ�Ѳ��ta�rܤy#�̞fb<�1`��;����y��� E{+q�I�V�$g:���g:����|u}?D_q��g�@		�TL�ݙ���]�bb��g1�<��<��ꅻV,6݇J���8�m�4m̆t]d7a���{�΢�bpvZUm���3������H$��OF�v�ú��1{���lE�Wa�#���2y�$�+|�y���.�'t�;��{��E��'''��k]�m,u�ʹ�sH����KcX���!����ce�s�sh����6iGa�cVfn����l2nYZ��r�WK��w��h�Qͺ���c�<��UNV�t�u����������^�P⚫���5�3��`d�Xh4�U���s{�\���K_��[���\ о��g'���+��M�6�մ{���3��f")��;�����\�N�J���I�#9����@�����C9ò�jͰ�q���ZiP�t�BU�L����y�}b�\ �<��Y��7a�y#�:$Y $�,���Ɍ�G�*,v��������\�N�[��ӵV̑��\�\������ڮ__N�/���<���>ߪM6̪421�6�I�Z���������	�ͤ=���g���E�ES�w���y������+�L��AQ A�P��4*&R	j+��Y�z�p�y��ip�E����ܥ�N۰�<��H<�Y��f"�W�X.��6��J��10����P����.�b��;�|���������떛;Ul�P�.F.F}�������W�5�c����o�Rk;�h�F9�̞d�&�$�@�.�yڊ���$g=�{r1c�+hU�l]�i�t��Ӻ���� ��+�`����F{����{���:����1���]JY��ӱIH�;���{���a�������b	�F'k�ئ�ճ$g������ ���%��n����A��$�m�m���k��Pэe*]�[����o|�v�l�,Qt	\nu�"���hջt��k��[�i�y��U�C��:]l.�S\�5#!t����<6��ȭXz�5{���{�rC��$#E�W@���^�wcZ��Q��B�:�h����w㿑}�?w�2y��I:�N�Z<��f3'��_� (_kV�S�w���}�8(f�{�oGvҥn�RbMj��r1��{<�ë\>�����<��E+���c
�V쁅��lBWt���-7jݦ�;	#���2y����umXwt�;#�8 �6��\�@ �]ю�[a;��wu��,�*�X�ܮ���|�wQ}�/u�<��Sle��[G�1y���f#��W��t�L������#g���%um�M1t�v�f�9�3������iR�WT��3�E���fA�^l+�e�)�n��p<{Cb66��
X���J�}��4�x�d����샣)�
Os���5duT�!3sZ�Q���$�a���/��}�R�B����7�+	Dd���H�鱯,���vb.���IE��L�:��˜�)��UJJҠ�k�
K��8�<D� Ϳ3��X��;t�$�=��2y�����ڰ���vF}�31#�ކ��q�zellQ��ʶ6� �������wul��Eɤ���<���C���w�>_
�c�|��ũ����Z=��f3'����ES	�w����H��ΒA��Q<{�oD��J�X���Ƒ^�7��Kw
�%�4 �Ջ����WE�J��j�v���:��"/���̞b�,x��vG�=�����3��9��V-�V��vF}�=$P�#{�ok��렝�[;���\�\���K��};��n�g����+���! �~R�����ѽfek��v���Uu�uu�==����n��6\q�:52ڭ�ȚM�׉9�˰��䬜��h3Q
fGL���Kc#V\��s����X�{/\�h�p�ItT[z�)yo�wa�[mm�E�q�lU���F]��K���p��?}��~�}���E�ES�;�� M/3ȋ���Զ�[��L�΢�b�fA�^l+�p|En�y�/u��1u<N�;	#���2y����J��v��uV.0�neVwZ��'���]n·O��3�y��H�C��o��O]����HJ�܌\�nv���E�������]��wc7ũ����Z�5߾c��;�g������w��3��n|��y���ߞAȸl]j[p5��i59�6Rr�4����̑��.M $�����aծj� ����;�r�Z����v)#��9�cA�F�	"�sQ�7�JŻ
�>�g��=���]t�t��fH�q#��$��&���B��]���#��ka�j���������;�/��>��<��Tt1��+G�?���;����B�5h�5Wa_n���;����T����R���+wY�"�Xf@�j��6ð���/��$g�?i�ϟm�١e�qamuS#�5W�!�P/�NrNv�ݹ�e${#�3'��G����]�+t�=�Ͻ�yr1��]ݵa�v��3�CA$�W���|З�?�}>��c�X��݌�SC�N�Z<�c@#�����u{Lb1h ݞ�Nf[X����k�N�V��+�k�zC�FE�Z�t�]�!�6ͼe�ʗ-L�*W6�U��ʻ�@�v�j���\v���`�ê�|y@�vM��⳦��{]JZ�n7F+{C ��o`k���B7�5ۂ��]�9[r�eaҪbՋ���+�>�����ȹ��T�j�X�̑��.F9#2g�a�uk���c�3'���'n��H�F9�fO3؏9;)X�a[���3�y��\�s�]+��Z�y�%Sh듎�-PH6*�[M;��V��fH�q#���T��G/��O�s���83я���7ѩ��N�Z>�c;�Ɍ΢��SUwt�&Fs���o5��V�۫�Vw|�uq��Β�}���wH�Z��X�g�g3��;m�n�������r��.�u�t�$��c��y#3���vU�n���&Fy�;�$Q.�<&@|��{�o�v�n��=���3�� ��9�о����������g�1ɋ.��XM�i�j�y�-�ǖ������њ��um��s�Σ|��S	�|#<���Fv19�����&{#9�gc����v��g�����|,
#	�� z�غ��+�N�H���y���7<�y�����a�R^f�S.Θ�U�k'�=�E���}dg��3�O�>��}�]ݫػg�|���GsX�k=�h_�~�]_N�s���Y��`��+V�=�c<���o�+�e ���23�y��gc� p�$�6�X%��2�Ē��H �0PU�j̻Qtd�Z���xZ�:yK6|sw.\Ԭ�%kV�h����g�H��4Z"�MZ�H�������R��D�����)�v���J��ʭ-.-�	xYa-�K��m�XS�5imk$��K㮺���:�Ѝ������s"k*a�v��$*%���Q���1'� 	 h  �����	Z��A�\���s�凑�Ľm�{�a�k���G@�@$
�w6���]��Up�(��mgOH�U+����I�?"��v���k��j�\����u���v�݋�"���=��	ؓX�c�3�{n���&�s��'����Q��.!�OG�[��ˍj��.�� ���m��(ڄ�nَ�Լg��/o���΁ii»B;(�
� E�Y��j$V�!�Z�N'��e�#WF�q�ף0f�xő�������FxƻVC�ܷ��gv�9���s��q����Us�m�qD&S������a*x�����NF�(�n�Mq,�9�ŃML���e��؝�?�#X۴�8�H*[6��U�;=q�L)����'���!dA�k�ݫUu�N�%���i��;1�u���HJ�qs���������Z��y\v��'r�<��\ӏ(Z�����M04�0�V���V���G�rC����^�a�M���ī�MpURe��:�3�8^B{Ll<ݰ��̋;�aU�5���ͣ��eוq+]�e��g=�?Bs�w��:T��)!��iM���tt:)�P�6D�/ NIg'��~�|��2�,pGث���\���n�ݧ��zt.����Ɂ�`���F��h�rZ#u���C&w=�ThG�xG�ì�1��H�]..�L���37
�+;�l<簄�Vƚ�ңsl����=��KZ��:ns=�ݝ�����ˋt���+<�g:��9�{�mӷUWÑ�1;�� �\��~Wn��H�k�1�I��g�����X��[����{�3ȏ$bw�˻L7b�#<�\�N�{�?p<�P��B�ӥs9����ګb¦-�M�hW�<�xgȾ�w�d�7�)7�յh�G@���|$l�:�5]UlH+	�OF}�3ȋ���ĭӷWT���"�bv3 �ۧn�������<��ԝ*oB�;��1�9F|�%���lzzV�]�v)#��q�=�g��{�Z�[t����k� 4$��Q{��V�=�v�U������򎉲7�(��"@X l4�}g��q�ҿzg/}�/���Y���`��;Vգ��{=g}�s��{�o϶ـs�.H�U���ɸ/k<䎄6��8�~w�����".F';�vۺ�̑��|��wG�y:V�Z�ȋ�1;��]
�x��;�����3<���@"�1�8L��Y�;Ϸ'�b�V.^Os������y��O��ɭښ��lsmrq��E��sī�L���d��r1;�T��|�w��_@4/�c����1}�I�Bյh�F3�ƐH�c=�yuU�2�V��k>���E����V��wT��3�E���g�g>}��=C\�CjGb\�Ҹ�M$'
�	]�b�FNz��6�A�\sф�}�]tu��c�mm�SQ��k��nq��s�6�\`�l�^h�&3,8�&ԚE�s��6�Qo�	�q�S印��WAc1u�	yI�9��Va�aH#tWX�WXg�}�7�̞b���Sn��G�1��2y�Dy�کbӥn�HϽ�{r19�vի	�ճ$g���� ���<�_A�S����/1�n�'���+n�U[t����;-�]�;b�����T��ݡjڴy#�fO3؏.�(2�V���	(n�>�/u��v��m���3�E��$fA�/7J�\>����1tjfSL;���{��3���y|}?N��'f8��(�w]�b�7v�&бv-:VHϳ��-7P�w]��a;��wu��2!r3|���񧾧{�d�H��`K���~�;ޱ�M<bյh�B��d�i5��yU�G��i�f�>���FD}|p]�B�3�2�]]g���N�ٵt��ҷm�b�2F{�ɠ�C�gtf��5f���#2F.�L�mӺHȅ���G���#��X\��o��pW��A/أ��Oc�b��g���NF}�(W�Z��رj�sճڬl+�k8pPp��ʧ�}>�s�k2F;SO�mZ2!�u�#<���%U�i�OF}�3Ȍ�K�m[j�2Fy�ȇđ��;�66�ۡk�5<��Y��;���^�WGj.�V��/L��٣q���(�i��ݣ{T�:���y�����o0/dF�n�X�tP�צj���[�L����[=
���G9y0왎�O���b7)�����;�R��w���s�Ce> Z��JH�b��y�p9�Kt�o=������g�r*�ӥapOF}�g��8�V�v.ْ3�FD'#7ȩ}�>p;������Y�12��xūjё��<�{���w�c�ּ���U�Jf��liD�.��?�~?A��y����Jݶ��&d�I=`��7���Mћt�е��G���Y�1ty4�wI�:̑���=�U�ӥapo����u�.�j�Wyz�.\��Y�:��\�*��m0Ӻv�v.ْ3�FM1��x;�R��R�}>��7�̑�����1X��=�ά�ywJ�YajdL��Y�{�GDs�%�L9�(d��7J9P�����J�1�l����s.�Ǉ5�jR�YM-.t��;�\JԬ�i+RV�U-)�Z��V�$�$SU++VV��f������I$T���a-�V���4��+6�c
��*+D���+Er�6�}��9�P\�5�E�6�ۄj=�h!3�s�!�g&\2���$@��}�*a\��WȖ�)D�@��i"�d]F���; �Ҁ��9�9]�˪�����$l�2F9[Cպ�7�ջm��L����"����V�t<�ʽZ�Zi��٧l;I��N�\R�q	���	7u����I�-Q�s�fH�*V�C��X5�t�.�ϳ�r���N�)���-�{ff��ѓ
��!IJ��Ft�S n�D$��,@�Y�D�E�G�}��w߉]1ڗx�z�����Y�1��\��N�a'aPQu�-7S����Zvū�tdC��2F9R�.�(2�V�� �$c��wP��nڶ��&d���	�̃��0�е��+ڎy泻����T�wI�:̑�DV�C�>���l�mX�`�n3������q�aT�Ex�qj<�=c.��[;��)'s՘��=�#;kl�N��8��\�B�R�p�H����t�8��ŋ���c�>P]+쵴�x�z�M��0�<@�஬J���N�*æ�]�����pK��3�V��g��FD'.J�a�l��#"�� P��/oԩ7a�L��>����U�O�mZ2!�u�#<���A����'�>���FD!�}5JҶ�V���E����藓m�Vں�̑�b2!9���A[��}�.��)��4k4{���F���L;���s�fH�"<�U��J�����<�"2!+�rZ��ض̑�b2!9�	�Yv-��\�9N���uZ�z6`3�v^5o�t����#���~fH����Vգ"�Y�3ȏ.��H+O�z3�y�������
� o����(;��Aܬv����3���	�τ��R
�\9�A�7��:���hy�V����v$t�
Fش����a�$dC��2Fy�"���:V�g��y�	U:;t��b�2Fy�Ȅ�fw�Y6�V�]��Q�Cy�mT�"���ʊ��՞7˪��Z���;γ$g�qw*���Qk��FM�{I�zI�
l]%N��g��<�ȃ����m�RfH�1��@$P�Y��V�����fH��&6�!�[�w����G���)�t�.	�ϳ��#"  �����Z�s	q����ʳpc�	�]h�v�\#�۶�K���g�g��86���TR	 R�܃B�i��zڬ<�r��=�Z8v2 �m;��
�+L��^��4�{��Y]7]O�:t9f��U��8 KW�9�¯X�Œ�D�G R�����e�N�ғ�J�V�ض���#���fw�jJ��w��G1�$b]T�ūjё���G�B�IS��=���"2!w#v��3$g���NF~ ��o���P�UT�s�,-�E� [ڊ�W_����϶{�w$��N�A0�2/�c� ��>�&�D��E]bߵ�s�9��5�x����wџg��FD �}I&�ض̑�b2!9��K%j��b�ڎb�fH�D�Uen��x,
mn��R[��wH��;�jڴdC��2Fy�Њ��������b2!s��ն݊�{�ۭ�q3�U^
L�Tsڷ�����]R����B�fHș�H&�FD/�fH�b<�%qU����Uj�b��lB��\���(j�<X\#>�3،�NT밓T��$g���\���K%j��b�j9�^�2F!��K�����>������g$gN*�Z�v�uש�t�3u�{��#">�����.�
�6��k��v���Uv-ڻmؤ̑��2i$1��wFmUEb��i  (g���;����	�t���Y�3؏9vS�°�2F}�g����uM���$bi\�>����x���$�$�䌒HIT9�� f���-��,����γ`��h�T�?O��FN���j ���՘�l�m��K3ln,3n�g���6��c6S ���.�����$ d�����(��!��� �X�'��_�Z����_����[�O����s���s�����8��i��O��eK~6hÞ(��s������(�~�l~�f��|���9�M�����������𗿷��__m��������~�??�M;ۛ�9�&>����{���~�_��������g��ڤd6Q�������O���iQ Ö̓Vl�l�l������hg�l6�`�4��Ff�
EQ�*�H 
�D�Q���4GOҸB�m��2��#����� ���Mį�����_��U�����~�������w���0���yi��������C�����������R�*�����,���F�������������쪠�����>����k_������z���[c�C��36������ӿ��~�އ�9�c����������3�����0͇z��O�G߿s��L��p�,4�ز��a �t�m��Ɯ����FT�?����~��
��`���#�xO����g����඿�����y��P���_�~!G��?�����|q�Uo�ϕ���?y�����������������?�������)Da��~��H�����@�?�n5���𪠠S�'�0������r����9��T�n>7�B6���GG�u��n}߇����~���+�0���P�'a�_����HO�ҿɄ@�P�����)��� 